BZh91AY&SY�I��_�@q���"� ����bC=�           <0��j���(%����H
��%hj�kZfj�D@Ѡf�l�MT�m���-���� *E(�*02��kI
�+$��T�����2�[m��@�b�Fѩ,��k-��ִ��i��+A�J��ٖڀ��,J����m�����.�6�=�f�U����6�ckk�Cv���k5\ݖ�0V���gv�R���mcV�Ř��V�k��R��3m�j�cUDb���j� rv�Ph�� �ҤP ��5|��l��✠� �v��H]k���N��i��J�.�r�.�k����l9�F�n��ӻe��q�:+��	*��M�i�&�f*�7�J� ��޴( W����h$=�{��Q�Kދ�����/i����yJS�(����� �w��(�G=�EWZ�;� 
����QիKVF�e�V���RJP y����(J�r�}|t)J����^ڀ�Ե�㺼 <i�q�wU�[�9�B�<x�UE
P��{���
*K��� = {�o� �_{�M�2ٕV�l��6�+�J�8π��d����@U}�k�^�( �;�Ƞ����M�l����mZ [�Ϸx�zj�����۩T�9�R �����ʊ�Ay^*cj��)T	+f|�T��oo���L>��m {�=T�6�U��׵{�{m�&�{�JP�my��Us����J��yJ�AJ�K�=
����i�j�f�k]t�6Mf|�����T��7�
wK��*�U*���{�@Ҵ��w��B��������(�� !�{ǢJ��Y�Gl q�w�:�JTE��kSe@�Z�-x>�\��� g��h����tt���� �+��Ø w� r��E �s����@�U�Z�3h�Ԡь+[o ����C��à ��p���K�@��� ����p��� ��w օ�^�����J��[e&�5�Xg�UP=�=��Q@��x� Q� ��� �N�x :6�� ��4s��C��ŻJ�t=� �+�fѭ�ə��KfEO}JR��w�t�]ZV  mGp�(6���zW�` һ�4wc�� E� �n 4o   T�R�'C �J� j`�R���@  � E=��R��C&�FL 0&&& jz1
J���h   �O��%J����10 L�0Fz�$M�R����ɓ&�4���j3IJF�����ڠhh�����G�U���X'�ȟ������i�Ѐ7:���x|��7�~o�\=��{��W��DX��"�� *�����
@xx	�������u�T�QV�*I$��i U�*8� ���������Jb�-�lK`�٦%�)�lb[�6Ŷ�`�LKb[ؖ��%�-��[����-�lb[�[��%�-�l`[�Ķ���Ķ�lcؖĶ%�-�0�%�4��%�m�l`[٦�)�l`��Ķ�LK`SؖĶ%�-�l`[�FĶ�-�lKb[ؖĶ4�ؖ��ض���-�l
e�m���m�l`[�6�L�1-�lb��6���,`�ؖĶ�-�lK`[�L`�Lb[�6���-��[��Ķ%�-�lK`�-�cl#ؖ���-�lKb[�Ŷ�m�lK`���0�%�-�l`��6����6�-�i��ؖ��-�L`[�����%�-�l`[�����%�-��-��1-�lKb[�6���-�l
e�-��%�-�lKb[ؖ��m1-�lK`��6Ķ�m���Lm�LK`[ؖĶ6Ķ��`S����-�lm�lm�cl`[���%���-�l4��-1�6�ت[Kb�l@m�鈶�R��[`	lm����*��ت[ �ت[`�lm�lm����
��[`l@m���Q� 6�ؠ�c-��Q�6�ت[ blUm��b��؊[K`�l-���T�*��ت[`����"�[bl-����
��R�"F�m���A� 6�F� �b�lE-���A�
[cK`�l@m���A� 6�ب�b�b!l `�l@m��� �����T-������R�
[Kb�lU-�%�� ��تi�%����آ[K`	l-�[H�؂�K`
[ب�`#lm��[` [ب�b#lAm��c`#l b�lPm���A� 6�Vجb��Q�(6� � ��F؈�M0[`�S[b#lDm���A�"��؈��(��� 6�� �Kb)lTm���1�*��F�
�blTm�-�b��`#lEm���Q� 6�F؍�D�m���U�
6�@�*��i���A�
:`lTm����6�V؀�LU-�1A�
��Fؠ�`�lm�i��i�[ �l[`�#����-�lb[�Ķi��)�lKb[ؖ���4�`S���%�-�l`[�Ķ��%�-�lb[�S-�lM0-�l`[���%�-��lclK`[ؖŶ�-�l4��0-�l`��Ķ�-��lK`����%�-���Kb[ؖ���-�lK����-�lKb[ؖĶSb[Lb[ؖ��%�-�clJb[�Ķ�-�lt�ؔĶ%�-�lK`[ؖĶF�-�l`�٦%�)�l#b[����-�lKb[�hm���-�lK`[���-�Lb[�Ķ�-��m�e�-�lm�lKclKb[��2ؔ���m�lKcl`[��-�lKb[ؖĶ�-�����)Q߾� � 1���י�f�����L�"���7wJ-e�i��x��rT�0e��ٷ�����N�oD͎�̳��"�R���9y��ɫ]0뽌Gx�J�1G2�c�ja�u²e�[�C-��遝ڍf'f�l��'!��TN���ݣikrVң�*�򔟒sr����VZ�.���z�,��@Щ�H˵TУ�+Z�ͯA6�q���V��GH�oʂx��k-�́�ȃ�wI�ư�eW�ixw
�M�0���ŕ{���?� ��p�6�co[����˘��/E�J�k�r/�Z�v�%�೚�mܞ,1���u=�;�7n�un��e����K���DcT`�Bv٘�n�ɲV=:r�r�5��-��wm���ȑ#�)͓w�xccpiU��Cm�̪6Q�Y���Ҷ��k�K.��G�\R#�m�[v�{"5�r72��n]⫘Bj����+Y��8ΜśY�eݺ�k�k(Ė�yz��6N���-����;FlA
�Kwi�AV�����Y+�t��Qҧ���r�Ʋ��ź��9�)�7z�H�L�U����3e�qi2���b��]�k��op`)�L�T7�˙4�9"ݧ�����UyZv'�nn�F�W5'6�"N��3�AW.^P%�if�f֪�f��`��1�3q��ec���0�ӨXW��9��ل7[0�,�Gl	�yFk��4^T�ln^L���3[�V���U�Ki���amKj���z���ڻ�aSB-{K��3#���U�պ^�{s"Wxtnش"b�u�n�h�yU�4V�7n�f�}��p4�
�4e$#[�s-�r��x�v�i*��� HQ�A+c
�LJ��D�=�Em+W�E�VT���%/V��m
�����T����M��@������^�cM2�Y��nfJ"��?{IT�'1%��M�1Y������N� �
R�Ń�9���Ꞹ��l�ө{w[
�3N9����u
W�|�+콵m��l���m9�ӕU����7{�X�ji�Z^%�b���^�!���s&EG0M�V��h�n����<��f�x���x�S݆534�P�Y����W�n-����p�2�_���z��Y�#5J݁	wS�	����d�r�e��m�F�VPv��-6�cbf��{0棊�t�kS2aPk6Az3d�j��{эk�V�xE�V�y��V�';���]d6rS�
#I��'�H7jF��j�Y�ff�]l"ˌbj�={GT z��Ú�Q���?AS��<��j=��j�i몳[,f�f=O�7��r�h���؄���^��.�%�Kŋ	�X� ��-���BE�J4Ÿe��]�uì�4sqM:�3TCԮ�.��Å�$ :��Av�D�xj��y��T���%e ���4�.��.SoXyE��4��<)غ��ա�ۨ����{�\�D[��4l�{V3sX�U0Hܿ�8���=K��]x0-m˪�d�i��R�-�״�%�e�Q��Ʉi��հ�au���Y�Ȼ����ȿaW��u�ҥ%:��&\6�W��0)Ti	�I��'��&UbVn0�H�&CUvZB��V�f�D�V�B+�
̽W�e���ԚC]��ӎ��i��/v��xa�ѽQ��l�#N�.�6���t�{�TpӴ�j��I���
%r����uT0b&��r�c�u�i�u*[e1OS�LV@B�f�&�H�S�%C6�{q櫫Yg!�dx�]Y��仅�yU�v���R"ޒ�Za�직�O������H�We���3A�a�-i�Ǯ�Au��`�
���h]lX1��>Ɛ�9��ǀ�\��(c5�e�ɴնU��3-������K����z(�L�C7�� �F����F���4�tIY�.�YN婘���V7+'q�	*V.����X6�z�`�l!�]nZrAܑ�&Q�h�4�ٴ�	f�y��1Yh��4���ͦ-�̨"����pƖ&�9b�����4����Kkm�ud=��U7Z$�L,���ƭ���c�4䱡#���,���������{k*�lm�FYO���K�Ek�-�*��M[լj�kt�x�h�OK@b̭rI��ֳ��R�2�(U<[6�`l�n�˧�l]j�;ȴH�J=���&՜ʢU�F�&q��{�ǂͩ����ؽ�7��JMYBDz��Ǒi&�甞4�T��D,0�k��5��^�X�v3|�巛7P�$\�)�݋b�S4��u�d7�bY���(f՗*�Zckeh�t��9Z\tIzrjY֩=��N��-��:If��+�J�<�0�z+]1�F&:���&F$�����si�y�RtU��E��%է��kad����Qh�,3T4B�2˙����hV��x��4�;��g$�!�'/�,�J���h��m�2c��	�6;4�mH7sD�2��vQ�V6�V�8�o�����1�Z�a�U�Aaiu�Jb��Q��e�f���uH�8�ֹKV�<�<v����w�F!�D���ٝxt�u�Ʌ��wX�1��� ��g��ksV1��U�*��ۙ�H���T�[��7����a8��Sc(2mG�<W���m	s�'�PD���jy]Z�콹��{3]��x2s�0�+w5��X78m�fԻ�X����d�ek7Y�,Ր3s7ש�l�ۡ���2b�K�h�ԯ#<�4J�\%�[I�;w$2$�I�9^�^$�V�T:��&���=Ï^�Ǝ��kU��zI��f�E�6cL��m%S2�����%3�zܫ0����y2-V�-d�*f�v�V��V�-���/0B�R4ՇFQ%�q��n�@�gU�:�@K˱{����ۛ(;��	Lt�(uUk/څ��-��j��n8��M�iĻķv�����@�ݧ���o)`�vfU���-e��,��Lf��u�e�ZU��a��U���lY��r�J���!�$=���z����C��~,��a+^�Ҳe�▴_ኲ�Z8�4ݧ�?�M�omu��E�F�bʹ�iWxޫz��RƝ����t&��ر��1挕{Z2���u̭pVI�����VmVػ$�Hn9U0*ÚU�T����%^��n�{����UI[y0��:���Rxi��+[�X0�PZ1i7�T�k	6�~-"��Z�����h�d��w4�wxIb�L���iE6��IcQ��S3tT�fޣGZAe�r��E���i ��\��j�
�"�V���d��ӌ�q�~R��LkhbM^=AR�a`���Q�6k��׸�#]ޭ"B����-�XfLY��5��֣1��KA@��*�'����B�1�J��P%�F���wQ#��<��p22IgvPY.]���h#&�U��.֯�ٰ��uI��#����J��c�IWwdׅ	�Ś�:����<����S��zn�o�ZFVR4�iʼ+,"^��J4��L�����Id��aǹ��Yj(3jG�&�W��e��%;V�Gq�˙�݃H��X�7a�Y���^�ia�N�+�HͺО�.��Iq��5��7�j�e;�4bM�VSVK���ם�-��z� .O��eU�ۖ�$�9iT���17�ia;c.�Jb�A���M��ʸ�[��p)xU����֙c5��\���	��VʹYD�F%DSƕ�ZSں��Ո:���QH�j[���/Tz�]Z�ǧHo\]:kZN�O��u�.���t-^�^�f�óL��8�f#{CT������:M#�ܻ�Dm1�.T�;�����jŷ�ʃc%�E�c,����n�/^}j΁�Sa��gm�t{ ��aὔ���
��ܼ��XZxn�����#���Tu�,��m�R䵍�f��uY�U�z-�]jє�h��,�L��m�ZM�%��'3n�X����[Cu�3a�Tl��fjN���ZNnA1�!z����h��c.n1��
nM�{$V�a���1��n��3(�N԰K�fԨ�2���@��w=f�OC��n(�B�H�:�9��V%W�-=b�=`����tUГX����9k[���ے����GB4����`�rD63"��ġ�#���	�lX�ɒm�[��[zr�����`cPWOl���`�r��W���ݘ��q����Q��wm�X��8�T����ncbm�6jL�&V1f��µ���%V.��Z2�Hڂ6w*e\��=�u��ao4mj�iL��rJQ��3qə�*�n�S?���n�F
����� V�Y	l�v֬r2mUfL%�&qhǸ�sa�n��pP#z6���J�KrͫV��T��N�U6�;�z��Q��8.�ԼB�`��smAukhhsfݢ�[��J�^�Hb�ĸ��[�i��8Fr��Ѱ�jT����7V��Q��s��Fv�$4��Z2�2��ӳQ�J�nfk��QP�u���i��N��V	���8�U�|�^��V�^�8�R˂Rr�P6�r���~e`b4�#SsU�[�pT����-��	�ޘkӱ)�y�m�v��!�]f����Ow�޺�c+�,�T�FZ��53v�QYw�,m���{d4]1R���]��ڪ���e^�y0:9��l�T��p޺�'h��a�)���F�{��)��nO�sf��!��n�K�)��Af��qM
�!c35��̖�b4ju��K/מ�����6��f���5��5��nlZB��#ä`S4�,i5I���;�ư���`YU���z��[�/(�(J�iF%$MVb�[7mI�zm2�&w*�ot9��(nnC!G���=�DaK^�Y���E,Yi�T�Z��7s��`�Y�iJ��Ẃ���Ï$R���Y&ek1R�#��6��YL;���	{��YH��q=�F��Y����q�g���50��X����Yufr��"UV�.�BBk���X�����(�t���u[QM�q��Į�t3�����F�)툜��v���F�{zh����ӎ�^���,Z���N��m��]�n�ܶd�L����J��E�ͷy.�c�Sv�m��S�"s7)C[DnK�C0A����З�l�Ƭ&rϷYTq
��+T�h��ک-�^�p�͟^k	8j�]���ɕ-���*��d�.]���i���e���ꠊgY)�i�P�h�X�1��e+F�Kpa*H�T�����^���x.�M,���k�n�V,7&�v�vUAU�e����c�5��6�׭C%VG�ԅU�H��۵�d�3W1�Rvs&J�1�'V�c�+%Gq�m���ԭ5�f����U���o)�U���zLaI1�{�F˰�r�%���e�����m�YVFV+3$tC�u�4�
9��u<�v��Rf��sE�4T���ʔ�1Qh��A�[NmJ�٧SR�]��h���J����9Y���72�]�m�� �-Yƞ+R��F��na�!�U;ģ���4e�.b�x�r���.9��`��ݤ�kJ�]�b!�Ema(\�3(��N���mKQ���:d�X�e�[a=Ri?MK���0�
�%7rdXT�{�k����n<�P�2��NJ�ݼX[Sb��yA��r'+1�u�If`�2��֜�;m�UDpQ��{���qQXbi�b�2�X �,N�En��r��^	y�e�v���2�7k�SRʽ��bd���Ų��,��K��.��I��,	$	^��g�01diܦ��W���F��A��+4�7);��T���ۼ#^Z.��z��N����u�p=l�"U��:�u��v� ]ԧ[����x�B[�Z��+L��E�S�4�-�()�	�k)�P�SɸK#O9h^���ʶY��$<�N��T)^G/ó�nMz�Z+���>:)�_m*�&�m�]��D&:��G��]+}�����z%찘d	���������ҷ	���{p�X��Eob�Y8�<�Gr�m����A�Sѓ�x2 CtD;���A��\mo*6,�6<A�,���oȵ-VZ�(B�����v�P�ɛI_E؏*ԟj�֤ҵ��<��*�Àڳذ�#ޮMcjj���p�� kض!d-�S�qQ쨉��]Oj�`���Hc�$3x� �(qˬ1�W�(����(�%���'�����>�D G~��hzKi-V��T�(�$HX��ܹ��m� `d;������u� U���a��A��Sfj��12�o`�z�h����R־�9�F����@J[4""	�[31�8[�K�tD�������i�ͥ����'ݶ��n)����p:�Eu�k�4˛Փ�V)�@�+Q�,�C���j�Ѝ�5�ʾC��+�-�V�T�F����*M��|��406���@ �k;�z���U�9f�L �)W���˄�o�Y�Z �����M`;��NG�AJ��Z��s�غ��Q@sA齃j�؞�&��|-��ӄp]�à�h{�V�sF!� ��4.�����`�	 h�  lt�ܼvˀ��57N#��K���Q`8ZM*�K�buGCπ!�Ђ[��ø�q;5��Y*�.����5�G���t��ijV�Eg&����#�70A�=�����䭕�D����ގ��J���6�n�7�h��������K��ը���$��:6���<1�m��)���l��4�an��d�'�f��|��������3�h��۬@_)�)�KַUV����=Y�:KR}9�t�����<��D���  ��3FX/���%=� �w����8@q.�; Z&����!	,��p�v�:�i5�ZI#i>U�,��YiRۑÉ�����H /E�4 
2̫O7�  p@�/Cޣp&A�ۧ��gW������ߛ�� ���J���`ߓK������9�ï���/.�rNS�+��z��.תE|L��Q���-ۼ�1�[I��I��K����Q0&vtͥ�6���X�������O;��9ճ�st'oի��x�[c��t��/v<�"�P&�]�Юק#��hhЩ��XU��cٺ���KKe	7Sk��ڹ^����:*��ݸ���:W6����MY%��'cUt#V���h\�c�.v
ɂQ�r��|�mok�	˼s�_'�U���;ƝA;�ǭǺ\�����M�M��'\��n���ɾ�2�W� #t�T��H]�:e(-�Ȭ��zT�̋UJI��i��N]�ގ���k��{k[�oH1�����L�GO"�������o��,�q[���d2�C5z�Bw��1��% Ո7~RI-�K;�\��7.e��.��)��=l�#zsL⦈�f�N��dB]��r�ҥ�q�L%+Х�v:�}+8�sVr�n#���.����V��\[�a�=3x�a��빵s��yz��%Λ/Տ�>FCj<�	�-�q>�9]�`\�h��hM<ѻ���l]X�6Ȗ���,v�l�f��M'N%�0�[Y_`�\�qf���A-9����	իTk,qs�']I��u靼k�L��,�6|����D�ɾw�B�q�9�J�e1*I�̛����cȱ+j�BZ�f<�\�j��(�4L�a�|�mZ��ヨ��6�s�v~%nt=�e�U�A�3���OPպ�Q���"%�yK-��B�͹�JyS��\���ZU����6���'��B��{"�ݝ��eZͬ�k5ż҆���E�� 6�)z��oU�٦��͒��M2���Zt�g{�o�a�������\��5���h�'�����n���۫|�K��o+p����DQ*�^���=uGF�ٯ��h�;ʛ��/N�|^M�
���|���t!܆��܃�L42�4���Z�׸�=��l�q�~ײɸ��o!UB��X�Η��u٩�q)��c8�GC��f�vK�`+��ltX�۰��]�Yꗚ�Cb�KN"�\
�a#��O��ם��gX�z�mR��8�b�F�9��u<���龳�9��,�z�����I�ҙUZ]X�4V�.�֓���;&���oz���m�,��٫���x��Wr��C��p��l�
;!�����ֺ�p`�v�����n�o��.�Ӑ�Ak���76��ow]7#�xk�U�4�8<|��N��9�[���+ш�v�3��2��8�1�pX�wZ�Hϥ�̳X�Z�f����.�F��q-+��ݐ뙸�ZwO�j'S��xi*a�#�2^)=���^gm�I��r������4�������v�_o��m^�w��+u��4r�X���of-bQ3������zmw�^%�:Ž�x�lu�J`�|��ѯ"O4�-3���3�#�3���7���|�N��x�4��ܵ4mjW	z�&t�ӏt�W挥���o���24)�C���.���y؇4�'�.wUX�̰��YGz�
!W%�k��Z�E�]6��Q쥌���[��cu��;Aj���X��n���68��:���/r˥��<���iYF�_wF۾��y|�v.������,gnk]ԥќ�����ۑ��h96�|S�R��ɂ���ɼB�h�0Uwi�.�X�8y�]��rJ0<�,úZVe1r�FZ�ȧc�x�52���;U�b�Y�KY*��9��S�Ք�M�9�72s7��Q�����U؝�#�Zs�o�5�Gi�>3[�H憷��!�*��*�̫Ͷm�g@��2�>�ɈL7Fo-̕6�u�{�72l�u�c
���Rԛ��:\Ѭ���TcV<-�vla̵�gv�i�=[�ʥOo��n4"ȍ�D}qbk4w#Աءzb�)1���7�Q�׀]��@'q����a8:l�v�˱��C�[�P�r���E�'������O$'f�G;��w5;��-Um�c��)��,T�l9��A{�/&ݑ�]ӧ�y�.����أ�o�ڥ�]^%g�{�c�sX�}R����df7�Vq̧��M�#����d�w)ȟwrk�ȧU�m�xKB.%�(��˼�`��m�l�-6�t�˺Yf�%u�[�9�lvi��B�H�F�R|��p}�$�0��W>A^M�jʣlu#/zoc��e֑�]��6ȼȉ	�,��|���3G����O}�QQ���*�&�G�&�
��R$�h��f�U�Q��k@zt���X��Оj�|)��~�1�f\7QFr�����z��;%��vS�yZѡ�ܷї�"*�2Qٱa��Ca-��5(��R�2���J�3�����ꦱX�x#��M����	�}�E��5�dSt3�[]&�̚!_}A��xvp��:���֞d(Z't�&�U)�R�7;Ry���i{��c/�s���ne��n�J3.4�ѷ�X*<>�����Y�W]ʕ�!�T67 F�q��V.�fP[�\��y.��8��&+�8�[�0�װR[�%�K��p#u;�Z��N��0ڈ'n�����L֋�,�8MV�1��:�X���>��2�8VX��F��ɷ�)�zou�8VX��ё�`�sB��ugf9h�%7��ӷ�[�j�����3!`��]
w�h�5|��V�YR�X������L�K��sm�&�^���&��/*�"k�%cz�d�������C~�v�,aU�qú�ɨ��\sD�f�x����+�gdBo;B��t����zފw
�N�1.O�7T��8�)��
��jm`Ƀ���y8=/u�>�B�"�Q����q7L��;�$���]�=��R���5Ǟ�®;���@w���FZ)���a� ��[}玒�0��Y#�I�ku\����T�ż���ʝt:]�[/2�EZ6�;��ݤ4a��q� �������vN1$�r�Ҝ���7sg3��0l���k[Η���ج&���W��*p���^4&K5��''s)�V�*r�j*|�M�"�d+��}��\6�{�mC�D�����F�p(�s3$9`��j�9�{�:q*U�V^��iZ���ՙ��7��'���)�۵�SYܲ����3j��/�wf]������xcmz�釺؊a���V��6L��.�֏jЅ��=Z�YGu�9c0wI#��,t���� �I�^�ն��<`��Rܙg�v񱣜sMByr(����Y>Kc6���:�NBis��+qY���eP,FR�a%�1��:ם?q��U�q�\r��-�*+���əML�3R@]���U��W�(\ܔ�[j����̬��e�X���F��mP狙xe!��k�z��f�rY��u���dA(:3�>��SE�n'eI�����]����~%�s�x輺㨚Τ̎�۱x��w+he#�؊({�Eb�,W�:-���އ(�H�B�c��=��N�%(֥p1o���;h3�K�ݝ�i�AK�@��vP�`�V D��p]��//u��G�c�}�Y��CrfX؞��CLXv5��,��7��+V�![�!�[$��	�0�v{Y�>V���-�NUCqچȷ�W�B'����B��܃{[��t(X2P�����%ŹW]PuAR�2��;[{]�/5����}h��V^Y)���w�.차,�a���kb1��.K�h�G�K�՘��p�Ku5�o��μ�J�ekL5�:�Ge+Y&�Q��n@�_�}���w�E�_�3� �w��	��,�]���3Y�=��z�3@�#����N�^�훦:� ����ȴ�T��I�V�^Z�� ����	b���!ͭ
�$�TR�>�z ��}.�N����.�P�[��"e*��u<��Ⱥ�eپ��;�Ho���j�s	��H�Z���9kB��n���E�>�py/06� f�y�RUn�bo�t�	���0���@��K��I�`�'��Ac-X2����P���9���l�b���Z�\쬗ǩ��d��$�6��K��Z�]^��XaׂVҺ��R(�$�T�8jA�}c��Z������|����w��{ȩi@t�.�N�Q�[��Õy�+e�R�>�z�����1ڤbzu��5B�K������W�zfgD,t��.�fśy�=���5�sxp��`��L��J��0�CD��J�S:⌛kaX�I/z�3��b���o�%�:M;�w�a��]N��Y�ub�N����汌���T��d��Q��Ya�uh%�33*w�C��)�'�&����XIY��k6���;��5�n.��=���`G���F��2D���ו�jw�5�ˮ��gf�;c�\��b���n�>�Ƶ6ȅ���v���G
S,�ޅe�B괽�WX��y�TAL��v���f��V-b�G��*�+	r�cF��"�`l�������n����k��{��
Po;��0ͺ��^	��+w
����U�w�r��]�+A�c�$Ո���xy�H�� �TRMy��)&��t�fˣ�e��&Q��u�S3���)��:��9���6��z��פ�YG���7r�Tvk��N�|���l,jG6��͌����5im�����V(�.���Hɜ�MAlC�c��H�'|�h電}�g>b�	Z��.�������ܒ7�L��P���v�U+M�Ä{�J���W���#H�w}�P�S��cޮ�ꩅ⢁�h���/��4Ι�g`�)���U�&�]9�fMY/�����U�+oE���8; a��8�e�OS+L�va}���L�cN�d�:�Oh;z1�5p�to[ab��E��K3p�N5���gr��0vf� 3W�[|N�%Jc޷�%��Ҫ����rs�V���Q�Z�m*}b}���n2�f�ؚ���K��n�\d�ф���~�%�Qv��R+�=���ց��6���u�g����{�a�YZ@x[�%��,WVa�T���;���e���+p���qT�k6���γ���Ѷ�>���uZg���^Ԯ.��{���!)7WC;��Fn��Q�,��l��^	���g�t�(�ֲα�j
�|',H+�[˰8Z�"TGDm6��17�f�qBy��y��ݬJa�7�SћR�X��3S����1�}Q�F�*F�LX��v(���2�N� �Mt]MUǯ `"ӛq��7֧�Y�u���w0ëVcuAib�ǃt�m�%`Wg OsCR�rD��o�1.5�t�5y�ўPG�V��ɧ8�MG2o|��e����W܆�w׶��/�$g$:���J>mV7��GIE�7#ʻ'�Z��i�L���uҢ��M	(�ٜw��զ��v73�(VgcZ��G$�_v�vp�]<ڹ�b�=on�̬؞ɶîf�8ա�u�ݫ���o�"�/e�44�ȹ�T��t���"�ֺŵ��*�f���Պ)�X�f�@��Ns�`�5���6V���pƻB��\M�>�'5U�9�`A�#�\�MR�eN�f�\C�k��Q[om,�y�e�-�R�͝+`)�����[���<��e�`=�5|Hj��ZS6J¤Gi�V�w�yv(*���:���|�Ait���&?�՜ ǀ��bMW���Ǉ��r�c��W*::W	NF��h��+O@��%E��5�]�x�Q�{#{�O<M�'7b�i:~��Wm�h��L>�*�Z��鹓�b�h�7���U�*syy	� ��͙���z6����y��b���� y����sU�/WS��;ò����-��8&y-Aׅ�\��%�>5��f�g���8]�����#Zp���`��kxGy����nb۽���<N����ָ��ح�wmX�����ƕ�չ��:K�)�@��̛�O������[N�����3��yB�	7r���vxI��T�5���Sz���
&I��{��OV����2��՜�#O,xz�z��U`t�H�h���}�.Pᢺ�)���r����~֪�NK��dA�;Ysr�����d�1�?x� 1���1��nj�wz�d�4��y;�=���T;�!'��v��@�\֍��*-Un��[�3u�<�z^���5R75 H���Q�;����^F᪠'�D�52�PU�ה! �4Me#g�2ܯ ��]��yr��B�'�=�Ym��ή`y:>	.�V߽�@�uª2Dl��5�#���C�û��,�ө���fsy�K�&��O%k4H)؊��b?��!Y�9z���B�(�v�(��Q��^ԕ�7���&��صuPM��(�`Eה��B	�V����tU֓q]J��K�s��`T��=�>0uu�d}=������DPG����u�(����!?gߧ�����������_�#����c��5�C��7�Ղ��)��n1k�yM��v�d�Y�֑�Y�蔸���b�Ë^U�77�������;j�nQ����9c�1�-[H>�x<�^3䨚�lI��V:��]��D��6Uu�/z�b-�T#���br��s�������-SP�j�F��@] ]���-�ai|�}�@z�HF�Y���f��5>zJ�и�u*�$�k��,�||�a9�f�SID��T�.wp�����r�oV�`g�A5٧/sO��6yb�A�QG4�ҷ��dr�`Sn^��ާq������Q��&Q�.1��1��!�ƋU���舭�6,u��Ֆ�.BnY�`M���!EA�u�ܼU�F�3I�#���(��x����Z��sJ�Yw���r���S�7��"W���>v�P�Fv"]�Ś�a��=�K�t=��Γ(�:�udii�,�L�{zt��/l�׊��F�βd��l��N��Zpl]����b��İ�_XKh��ׂL�ZY�V��5��>V"���-5|��j��T�x��ռ6��r9�U�9���^��1̸K�A&<*��(h:]m��Ll�u��d�G���k�Џ:��j�S��^�!�9 �NYE��b���q��h�y	˪fƆFL[B��~��t��8��8�n8�6�8��8ӎ8�8��i�q�v��8�8�8�8�ݻ�v�ێ8���8�8���8�8��q�q�q�qƜq�q�n8�8�8��8�8�8�8��q��q�qێ4�8��9�fy��/��c9Ae���v[���Tn�Z��H����]¨�io9��6G���K2m�toQ�E*��ԷY�����Y����/�-r|�]���yvح��/��Y�&����D�Ǖ�W��v���%vڵڙCgB֋�6c��}���*�&�T����E�y��zoFp$�郱7�]�`��}�(8�5�5����sE_U��G�Q�W8�J����4A*ɜ��o7L���� �*�F�����\��;'{C[6�Y�
��c���d̝��i�72ݹG��<��1��7�ڝ[MV;�Ek�W����wr�Ĥ��]ԨEH]t2=.ky.�'�.��kç��B��ޱ.�e΁��V���IyW"�t�;�^hݹ���f,w{q
�.�Ao�:�j߲5KIn8��"U�g�Qagm[N����dO@Φi�G��;�y(^q[�",K4<�l�t5�|�9@V�.���/k�o֨,�3�����ฃ1������b�t��.���Y��5n���y�(�&8 L�ӵW�EcC}y0�e��#�����e����t�I�k��ݰ.�U�x8N�K1��y6��c:«��Ye��䤆��2sk�}�>�w�y� �W�_<���cǏqǎ1ێ4�8�>�㎜q�q��q�q�q�q��i�q�v�4�8�;v�nݸ�;pq�q�q�q�q�pq�q�\q�N8�6�8��8ӎ8�8��i�q�v�q�q�x��8�8�8�;����2�;ƆLq��N@�i�a}�qGt���.Ы#�0��-ϻ����0�1�y�/^�}��\N�������.C;546U��eCV�JKk�q�,Ȗ�;y!�e�i,���nҊ<
�^���+�]���q��2u޻�S��1�I�%r�)�+�Z甸t���'n�~��]3�C�TM�➵i;F��"����w��j��V�`�s(j��ۓO^sÉ����U,`7�Q�dr�t6�뚝P��Z�~�v�,�����N�-��#��0K�8��$q�Q�s�ݻ�ҭ�n��,�������;��<@�0_)Qĩ|��Q�6_\)m'@�z,�H���)L>ۻ7z+bݰyw.�o�8��F(�Q���#Kɝ���=��Fm�w�*��8ę4.ӵ��L�[dVX��r"�kzG�!y�AXs!�k�6�7�tz��s��GL���9��b�,sD�7tގ��la���[M��ya���S�z�v8��2x!\%)g�'V��;���W��v��ʺV����J�����/m�宧:��<	|!O�æG�2���A���s�޴
)R�p���u�bJ�A�u��-$�ȝ�mvR�-��n�8�8�8��8�8���8�8��8�>8��8��q�q�q�q��q�Ǐ;v۷q��q�N8�8��4�8�;q�8�8�8�q�q��qӎ8�>8�6�8�n8�>8�:q�q��q�q�qێ8ӎ:ג��%s�9T���0;۔���Vv���C�m�ɭ�0U+�kz�MqR�νw�6�����`f���Ldީ�j��'*��ύ�A�M#��!C�Mh���9vNM��T�P�\w�l��m�"P�r�+��н�+q��[W�<[�"��
��f�B�8�����tE�#F��p��5�������>�B���Å��v���򿍴@v�-����*V��%�r�YT�"vĢ�Q��i��v��8�-N�Q�G
8��НƯ��7�HC�ҍ����y��˻.*���U��r�� {Hj�Q�=��ݣP3���0��]>I)ߖ�=�{Rb�q�˛�n�J�m�N��̝{6�S��z���f��y��q����5<�r�[v:��CN<o�����UUOF�w�0\;w��q`�p꺗�g^�C����fط�5����f`Ȧ���T����X��a�c�4�(M�ԦeKW�����<�r�2�z�iS=y�����WH]\��N18j�y�3��ԯ^"�2t����g1=�tˬ���ێ�2`�\���)*U{H�w�'uAn����/�=jѳ�r�QJ(��� �"�%ٛEg��9���s���t���n�08��]2�$��@���Q8��;VN���<���_�U��m�����i�q�v�q�q�x��8�8�8�8��q�q�q�n8ӷi�q�n<x��Ǐ���:q�q��q��q�m�q��q�q�qۃ�8�8�c�8�8�i�q�}q�8�8��8�n8�6�8����w����}� StY]�Q���=��xw��hZ�������:�5���d5�4��dݔ�*-�'`��U��uM�9�H�%������]����N��1��u�\&� ��9�UԾwF�V8m��
�p��޶;�t;���'L�x������ޜ������x5�y(Cv�
�״�[����'�c��)mv�_*â�fQ�ظ(c�n�T�e`"�`Ν%]�k[N�=�I�M�g�J'c�R֟���CE��!T��)�iKo�,C�Z��� {ݛ�au�\�b��|�|�cޱO^�pW9���u�W$d��]8�3ػf�յ-��G�KM��U���c  �O�˺�R�B�5�Y��l�_e�	o��[6��z@�q�NP��n�6���ڤE�ƃj�MG,��e�<If�~0'���(e�f$�Xv���i�n2�ڪ��;�թDRE����q�tH��풢9zvj�W�=��Ma��1�X°X�Q��M�GF�ʪ�˗TiK�*�:��h�2�jV�.���D����<q���*��H^������}�L��a%�9�1�s�_�������kh��K��3���Z�{ co�^<y��tZ�UR�?vE��5�E�� G��,��Zs�q���))�Qo�����2ⶨ�.n�1 _�1ZZ����LmˬE3�`c��ޣ��)+޼����r�,�]wc��C�(&�R����Q�9���9���S�O\g��\�]A��r�a\�?+�vƖ�V:G�9�˙���D�`u��:l��ۍ�d\5��O�&c|���ʾ#y26��bb��D�=��r��R1��2��RĠ���z�t;�u�>��3���뵐����p��X����)��ZX�II��A�k�5vl���-�jyqe�UQp�Cs	٫�2zە��PG��1�tp��G#�u���	�1��L��)`Yb�&�8�5Z�t�p�N�b�,���d�c	�co��d'G��Ty��{�A�q.�ګ�(�)ú��k+��̝��<�Q�+�z�V�&�Ψ����n�^=���:$JY�>ՙ�c�8G|�&c�=��n�3a��Eݎ����]��:�vD���lZfw����:H9h���,�7Kw��P��w�s�{K��ۭ+�`��wZ�\���+U��]�̗Zr�Ymi�@�ޒv��Wu`\�1�G�&���ٍd���>��T�}�UŹ�;ot0q=�����9ЍX�̆���x�/8" [o�S8�ӼE?z�U1jv���-�8�N�2�?�=��Z���M�mc���(�\���x��uʈY)����Nsj��{
��$}7/���B�e��L�f��8��Q3w��v��>$���8��ZL��b�r��aUp��3t�9�N�ne^�4^�'7)X�I%��5@�'��;��=�t�7�^��*�^"���۳�N�a����Y�o�/31*\�!36�ܮ�%V�Q��Ù��jX��IUY#��/�i�V��'��	3]�c�N�(�T�t����Z���3�ʰ�<������ٽu�����-*ђ�9�,'��"1�fuS����þ�k��7H�坛�]�9%\n�G��WUU/um���*<�s`�j�[�^y&C�$��,Y3���F�����9FQ�`|=��s٨̐�E�sip׫�u��fշw�biJ�k���BU�z�Ĕ�R�u���:=)!�vB�R*�����UDűԷz94<7Mj��=T���-V�ֱeT{�h�l���C���݁�.�6��n�I6wI�dLv�n��4be�z�6Vj��W�"��i0*#:f����q%��Kn6a�.�g:�;f1 P�����m����$��5td�BbN���^wj��#u�f�Cq�{ΝL����3GGݕz3:�������j*�Qw����YB�c7�3zy�g7-��$S�ʱ�
ĲV(����%�v��b�t��B�=����m7}@m���kB�*nA����[s�i\�z�3�xV-c���<��+��^�H]�Hn[��mAƁ$1�n��/R��F�ͬ��D���T�JB�f1fj9r���٥ �`Ç5ӫ��iu8��\'&K���"5��Q�@�Jݺ��:G����j�ݗq`��p!�i�s��Bۜp���j')c麯��t
�vPW1-v�)�ǋs3X����_<l�Ho>��;/����J�B�X���:J�kظ(Aa!U�e1��vj�]�P��A�]ݴ�Rz9fMk���zf��Qձ����͒���v<�Pr�z6���z�^�uz,.,.u2H��Y�.��҄s�+v�&U����8)�|�s��A���Pf0Q���ƹθx��c`7L!:Y�K�2���sK���t}-w"�꼟5�+b�"G�!Z;uI�dބ��y��#E����U���\��o1�sq���Mf��[=���Ѵ��1�ԽJ��$Ǒ�j��اd=���ug7��:��k���SX7�t����c�o�������'6�(�=mq��N�QY����̼�`�y�`�G��oeaŤdg�^���&r-ᆮUV����4)�Yٵ/�$�:c�N%��$������-���~܋�Ǆ]Q�%2�u�!E�goN�[gw���R����o���i�g2��q���x�,�}�r-��J�}y�&����1�8��]��d+Ne1����AV��I�h�SH�ҴCwoX�pi�^Uv�+��U�O+RZ��,V��k��2f٤VV��q���g��7�C�;�91oU�ӯ-K���!�B�e�Hp�>�L���RV�r�;Oz��K�c6�j"j.���r��I�nf�نq��*\c1D�*\C闎2Պ�g��n��;Y18�+������%���au+��R�rufcΝ�g����ʗA�8�ӥby�{w;f�I�u�S�݅p��ע�=�hm�N�K�����UI�\HCv��αw��۠;۽4��^V	�sFx��n�欰kr��%.+�˵!J���;I�F/����K�sT����],�%��0���E��N�e7-fM|orF�t��e�F���+�ֆ�r�/B♇�Slb쫥���.nn4��x�okS"t��gٌZ�
�ĳn�́[)�PO3�]���B2l�UϵrS�wp��������v��kZ���j'E�ݗ��*�sj)��Y��U<99t�h���m9m;����C`���{P�;.S3��ۺ���.�gV��1[q�`�x"�::m8�����SO�̺{�kj��/c\��҆�����Oq�6u)|2l�w�K��v�Ŗ�c{]�g=b��v�ʫF�q��t:Zz7�+��TM��f��e������`�{�ٯi��/r���h�܁s̠󦅴�='5���5ȥWǥi��$l�'n�:�<�Yӯ
	����(:����e��]N�xd�.�0�zG�:i��j���:�c����<I-�-U�z]g"th��R�SBY�X5s��|i���#��*�Z��-ɮ��Cn�f��Qԑ�����tʮ��{�q�[bzj��+^j�a�<rv�l�f*i`�ì���6���˖�����)��SMH��`�;1��6cT�^�#�m�GY�
l@���tgإv��'2p���Zi%.Zm	�;��)jҷ-��[i��]�Sh4��q�n�f�y�ŰQ��9�o��[��Ψ�2m�A��7u����Ř�v����j��:P'U��Y��q�A�9�/�z^� �m��*�-�vm��0�#I���u���QYm�^b����b{�F��4�f�����
�)�O�߷�r�?_��P_Ր�����~���?�E����W��Ouʿ/��>kʞkZ�T1�e�UP��RH "Ӓ�TZWT?�hO�	Z �b�ԁ6�A���JA ����R��j��S���%$&JeZ�E��7B���~�Bah!)�̄%23����mU1MÔ���pF >l�CT�D4�@��4`�	�	��P
LH,���7F��&6dfNЊB`Q�8'�m���#1�¦�D�%�U"�څ �BQW�>���㾉�`�v/sx��yK�9k7ʉѕ�=�����|C�z6�Kh�'"�Z�Jֻ�LS+��ֻ��..��s��4�r>���*>�Ϊ��:�"H��*�	���� ��z"�����i���Ʊ7&۝6��0��O��cXj����k��k����iV�#S8s��WX���rR�r*2�'8�ԨR�}�te{\�k3$�ڻX�g2�% շ��(cW�
�u���ykZ���+��^R�^�?�Z�g+a�vL/ �b�6V�hT����Z��%U�G��J�ou�&�}�-�/'^r�K͚�YyS�Y��	�r]����I}R�6�6d�vJ�dA{��$�0�m��V�,:�\�l��u���j�%�N��Jҝ�(�����u�{s�kC=1Qװǖu[MV�݅�Y�����hr�I���a�}�UAG����3E�[0Y�m|y��m�X+��q���8(�V�'�h����8���k�[�]o.�e�z� d���iɫ7�`o&Ҿg�dzl�o!9�f�ÃP��n�}&��]�K�|ݲN�f>ն�@����A���ۣ�sC�M��ڲ�C%������g^.|�W�j"%CA�%
T��P$�q��D�'
�e&_�QL$"HQ��/)���	���-�m��� a-��d�ai�Qp��ʒ�4AF	0Ēg���-���\d��ۀ�Ll��FS��#l"(�@`�"A��	ċ��*FL6ZD���,�A2��KD�Ɣl��bE�a��ܑ�.�jS�i�P/�A2���j""RdM4SB~��Xi�?)"M2I'�	*��/��G�e�؎~2&��Aa�L1��M�
jDG�10Y��mOж
d�1�V�f�"�eH4���-��DB����ޱNQ�B���d��ۅ���U$ф�O�~seI�Դ���H��$�Q�A��I�[�d4!`�J��h6Y�@DR�D�L�A00� �@�fH!R�q �a'n~��A�H��@W�	 �Đ�
E�	��FBP���]�����q��nݻv�۷c�1��BB1��_�q"1�'u��$��r�R�W�������~��v�۷n88�a#!I!$!�c�`L3$Ԑ#$�$���q��v�۷n�pq�z�d
��BQZ����O;�s�]�߮���`��w]���mvRQ�㭺]q˧R��3#�wu��sksD�tRB2T�_^�x��nݻv�ǣ�C_'�4���UE���wv���1F�ns㖫��m�[�\�m��-�rwb��ˆ�\蹹�W,U��m�v�W���k�\���ns]�M�^MD�]�5r5;���\�5s�Ιu�]t���#����|�˱˹���r빎�1��]::��;�wn�ץt#� ��c�]�u�K��u�٠�r���i/��r���v̒hƁ��۳;�����&�ܚTK����K��C
d� �nRCI���L�$ʈ�I�����n���\^;�BWUR51ֹZ�f�������]���YR������J.�h�v%�ߺ�F��<6�7��[�N��`�>;��2d��}�Iy�͹Ļ[�3�����Q��7C����EZe���ч1ŰL��%P!
)��I�#$O�"�?��B��AO�\b2ciD�*B�,��$Ԧ� �		?�2c.�B�?�4횫��y{�;s8�b*�Ss^,n�񾼽;m4��7���Z�lU��;b�g��暭R����E�[�E���~�Ԯ獬��^���?w
|�ʋ�sj��)�{�y�y��v�
�ܷ�:�_���K����B>��[�L.��7߆�݂hq  �4�z\ܷM�/��y�7_l�1��q����A/x@�}c5}����ٜ�C�P	n5�]{��{�%�S�;�f�5K�^�l/,��fz����4=�i	���pRJf���龮^�`�|��fל�<��|�����*�x��=ɧOJ����:�hy����<�n��+Y�g���M�\�e�!K���۵�}��o���L����y��ݷ�yP�}Uy���p������V��C=��]I����ɟ�~�9�76���qOr[�{��(
y�I4�ҹ/3��SwJ^_ߙ�?9h}�OٸIsZ��i�=W�vfͲ�f���u�W��zyf��w�gm�Q�m�\�+��-�pML>����\S��o�$�t����[�>���Q�%��b�GFm%�ff}�Hz��h7}�roST�F����S��C=���`/��u���_b�.[`���W�}�2t>�6����ݓ�Ȁ�y���o5ە�t=s�n�m�@�l=�'��~���������\VxN���<���IS>���� ES=�+�7���42�?K������.U����蟲��t�/A��C���n�v�sz�{��٫��X��:8Uq�}�>��	��I��q>2�m�y�N��+��	��:�G�F^�z�LwO��w��� ɸ�c��z����k�+u��~��)t�T
M�@فG+͜8wqޓz��$1�ݽ@M͓BL�����}Y�|��=�v�5u媟1�JkW��v�3s��h��ˬI琉��,-�}���wu:�^�Y���`�zӱ�	������IＪ�����a�'�G���jCA=�g��7c{�y}7�w��8�\��ȭW����!NބW9eS������("d��*���42	L�x�����-֋�Ww1>�֐�/0Ny[�M��5m�j)u}�qM�jk�;����y~�������Df����h��Gj�e����7��y����_oL��J�#^����{�o�ds_�:�����������:�K�<5�����8-vOC���{ӵ���n��+ܾoD��b�Ł'�M��F�](t��k����	�|P����p��S�����;�S��>מ/Β�.�Z�v�zT�4�U浪2DQf�V�}k�u�~x��,�M����A�Ve���0�J�Uly��{���S��ϣ0���b;��r=�ˉk�	���~�]&��W�5��>s2J�u��Tuozs}�z���.�b����@*��d�d��ث���4��8��rz�,F�*=�w�n�O,kc��Pt��'�v�Pe�í2�}s[��\?={^��|,I�o�f�^c����i��ߗ�X���w.B�xT����4����j����ȥ&q��ZAm�w�Ab�����V�a-j���o��R#%Y�����G��5O�N�[��0�gLx�.e����;X����:{�	�g'Х�7��cl�2�;��퓬�>�#Y�7�5�ňz�:��~���ݐ�5s>f�S��xz`�i"I��k}�r���f�s�o��3y�y{�f#��:2���L��Ӫ���o��K�{�B�t����n۷�tL��@2c�S�F]9���u({}���h�	^ª�.}I��ǯ���oGm8r4����j�ͱ�	��CU>�M�;��i�zsX�oh	�g��7�!>�9潂z���H��ʅ!W�WU�+�������k�zd�Y�W�5<�z�k���8n���Z���*��o�ޫ_y����}W��6À���^(���t�Ǩ��'#��}���>�l2�#���{�/�;�|f�͗�d܋���f7�iz�-�Uy^E����5�M�w�֜�=.w�ޡ��,ؓ���v��n��$���3x��]44� V�]ST�J���(k._����1��'���W���lm�8��~���=����*M7a�&Ў]o,�D��&>!�3�t�+�x��d�/���Sf���q7:P���>��m�|�:�l|.�H�G�k72�iz�0w\�i��'!���+%�n�Y,�����\7Y{�'�����y^�,v�^�*������"�)��*�RΒq�f�|��ޣ��Y�ðNb�����`�я�W[�#X�h\�y=>���eH�Tu���g���k���s�}��!�����$���}U95��Mpʶ�#b^CP�#ގ�t'j�~�?o����	/+<���@L���>]���^���D6&xz�I}���=���}�=Ԗ ��o��L�����:MGng���ՒY�D�v�a�������<�|}��O������Q�ە����S�����\G\���z�	ا�$��7�oZ�1�|���X��Z=]<��
�]�ӗ��a�i#'m��ϱ�sz��n��	�x�h�D����%��s��}-�����<F�d��x{�f�TQq�^=�w�[��t���r���HL���{h72t\�co�f^]� �4�WS��+'e��X�^wb��r�t�qb���vmv����^-<�dx�BAoe+S�ɹt��I���R���Π�#ܙDV����[%v,^X
��o6RْoR϶yv3�/_�p�{Ꞑל��~�0� 絖�u]������_V���u�>�yf�s��5��5<ٯs�{3�3�ݍI����~��$ �;��h���w�Σ���]z�B�Ok�ל��}Z���rdS�~�jƽ���i���o�.���l'�͛�g�txm Ƀ��t�u=\�UFr���M|���ς�k'��z�}j��E14�C(��sp��xdY���z��a7�k���MeD�ȳTkɫ�\�;�q���O}�}��h�����ا�>��Xz����B�L�>�~åmq��/?��[���F	j�\tF���{���pd1�q�O����b|t썾�3�o��v�퐓�cʺ����f-��0CC����wH�x��A�4���_�o��E�/yɬ�0m\���{2d���YU�i�M���!4����*��=�C[�7�-��60�*��H��:��^���Eg�����:Y
!�k@�oh/��ZѰq+��F�u{��� ��������}4�T�����'�/��ܘE�ˤ���Ż�>4�~t��X�>'
�:T���}��)�O?i����u��_�̡�����F�3O��o�{S�'���O9��OOn��O�x��T��wf���X9�O�c,�z�0��ʤϽ�g�'������W�����.ۖU�=��bl������P����-9��z��t�fث�J�U���|:�d�
�����xmߖ�<Z�����<���Γ����?pӾ9~��]S�_�l>_y�8s��؋�ؗN�������[�Y�7ڥ?f��oj��K*RwS�訵�}x��O��}�|�����Aj��t�.v�vHl�H�h;'u�\�f3(u�fk'4R��\��jO�SF��N��PWw�Cs_�O�wa���<n6�U��O���:r�мD��չ�zӹ��(�����Ḫ��& ���L� �\�_TL�6]쵎�;7%H��e�]3D�Z4��v�9X2��|�p%��Pc$v�5.��?�]{��SĊ��{ݝ����[1�s6��4'ƾs7��k��;�9�2V3N_��:�ǡ�M�xei��/
�}��v���+�f'>��{�E���x@�p4��i�n�ىd�U�|a�/�&�sˁBe��D�/k3��z��$��a�m	>��4��Uɟi����=[0������49*��u��	��W�|H�>����^>�y�5�������C�uf��	�m^�V47ν䨴����W�|9��������v8��U��'�2M��c�4^٥����ϯ��I7b�&����ּĒ�I��9���=��+1�I�v�́"�px��19 h�����;�u��[���ئ��7��;�t���P	���[���=��¬CT{7�#X:�#N�q����s��|��u�݋PT2�4>{,T���`u�?yo����p�q8;4v�Gۿz{,2�M�b��&
�y�[v�d�.j�3hFgquZ��3DYj��Ivu�Ç:.w9���x���-G�6ovw)� �;��(�YCcsm��Eq�<�d���x�
y׽9si��y�;�i�,"�� ���ч�ƕ�o�{�
��=A�[�ŕ�#�*�`��ŉ�gfkω��2{��;�
�5�q�h�c^�������;��ئ<���,%��n��k|߳~>]_}�=~�<=5����3��lV�NO���&C�0�S��[%�������;
?=������_	��)�Z��?*�~�:��)L�}4�ڪ��=�I��v9�����<+q�q�{��(�}�@@נ�m~L`�V^�c�B�gt�|��l߹�;��́=^��{]P�����O��
��A�^�������S�����>A~�(=Z���������^��g��}��U��X�����<�OO))I�,�]MwE�G�Q6A�O�Cb�2��Tr��:ĕ���u��"�O7���4�1��u;�T�Vk��"*��`�ɫ���Ĺ�aE�}����-�4�g&�M;���P���1"72�	ʩ�C�h(6zx�
\�	����Y��,�7�tx��s!�����vN�nV�j-�՝s���Sȼ[��f��Ou�b�+wZ�ó�uM��z�9>V��^v�ϭ��ų��}mu�@�K9o.�$� jL���a����II�"����'���1+������%T����>�Ǧ�uڗ���@�L�k�Y� �|"��l��6*�k1�;n�0f��>�� װ�4�x�el��s8�6��`瓕;� ^A�����,���}�g�x�{�0�6c�~�Ts��M�dT��w�~b/_�fX^��iI�mM�9�<�ϗ��k�63YB���N�=���~/�����@{O�jsu�@j���jy����x�<gz<��zZ2N�\�����k4���Ў�ٴ�g��~kw��w���&�?K�x�����b�����U���������v�f��6vҩ�\"9�eZ���J�O}\�*�MS�u�#��� ��1떮�::YÆ-^���*_</��~n�L5X٫�F�������>Mq$�Q�5��/,��\�+�i��t�g*gEs
m�Kn��m��cUOn�Ou��$Z(���7Lƶt�c�˗r%}���k�����n�}yBUIcOv4x籈��\��#0pѳ�+O�y��7Ԁ�7pP�S�np��k��t�طNvB�,�5e��/GqQ�v��G��Wv��WF�J���-4a �Cy\
L���i5��:�aXa�b���kh���I�����|24Ҍ��jƌ��H��f5z"�Q[�M�Z)�s(�A�]����8����U�愚�V�"KA��FAi��p�P��^D9��	���Y���\���lӑM4�v+�Ү�C��Lkwی5}g6!77
x��%�]��/nk� ����8�&mgs�h�T�f�O[:7�m��\�Y�;��Q��f����:�,Q��ǵ�Ԕ���8mj��eQ��=�Q�W��ѸV�b�rQs�е.LmܛyNΝ6w0��[�7����ǻpػ�Bގم�6S�j�op���"��=��w��OJ�fS��eZ���3N���^��[Qgk��j%pPh��J��_J�d}wJ�ڛ��2[��sMl�c�F�,S�����v�m�P�,ތ<���J�,���s�p<j㡽k�{ғ��`ϻoޛ��R��y��7�1hkƵ��Յ�;;p�Ɔ�ZD����Y2�P��zk��82ř6ԥ��$��e�w:/A��)�Hi���/��_Ѿ��᣶��k�:=�nV�*��Md�y��R8��x�7�x{���s�w�J�%�NU�֮jj�����5�I�rce('q�	��Ƕȱj��A2�,��gL�^p�꫔�A�E��dU�/k��k �]};�1>�N�r��)�勺��rW8{zM.��q���0D�/*ڒJ�.�Ό�-YV�E�(����l��K6L�s2^�:m���jޤrcΜ/z���������"G�9��n�|⬤)���%���-�goP�����F�f5�\�Q"�	�(H|6����;h�i�nMZq�,U[��8q92�� ]a�q�!o&..|��ŋs>y�u���4�L��ѯuA��ݷ:�k�M��璸ޕ�2e�fH/%�W�)��k���7^z�1�M�͛�V+kb�!i�
�ֻOc���w,f�l��V�2r���Ru�be���}\i,��a���Z�Gi
&��5=�14R��.��t=Z
�߶L|�����ۘ�Z�X�4���.l7;F�� z�-��s_fm���D�٧O3s2谈o���+/_f�&�; �mk�z*h��f�w����w�����B�!��;�1J�v[s�Ԡ4�-)��un����ALJ��]^K~�/ǥ�#I ���|q�nݻv��ׯX��4��Ok�g�\#`2_r1f��o��|�7^<v�۷n޽!$��#!%��X�(�[۔i�$�B4�^�z��Ǐ�v������L^9��u��^���O�F���{���7Ǐ<x�㷯GeRT�$"�w6"�T���+�����:��L������^9��)H,HaDMk�� �
!|qh�bLE�mȈ���dɒ�Ih�c e61���X�2l�l)��H.�V(�Ɋ0�[�E�"�nX��%��@��p�O���-��g���ݤ�ۭ�k!2��Q�!%W:���EjC�K�ȹ�|V��m�-�9Ӑ�i"X�s��c�>p}ד�s���W��{��K(���_Ϩ��]�㾫?�35�ʿ{��Oz~���ѿ���t�beOo��fv2���$��ፃ_z�o&~T�?�b�0��_�����.!Fy�"=�/�5��<a�Ǯ�}t��^��L�hS����?��w��C��}o}琊5�Ga���N��w�7s��4_���x�\�Czo^�=0z�Շ�E�E�'�>��`4.|눔��ӷ�E�Z3�Y9Þٗ��8sL�Հ��zܵ^�@�~�9��U��-l�h(ޑa���ā08 p��23�D�4���dG���`�P�����M�lV��B3�)��۹��t���~�c�3���MP��*��ڹ:����]8�/��d�9�{�H]Z�!t�Z�F܉�Ƹu]�ӝ�F涪�T4�X{��#�s=����N���X}��`�ݒC�i�u�I�.�C�E7�<�Ǟ����!�X�KxT�.=e w;��� &1� `��?L�y��l��/5�]��{<�(~L���,�Ø�J��bj�5m� �@<BԁDA�0�����`4�!L�i�=�B�W�P�s�w�N;9P9�<=�O��o*W�����.���Nv`����.�f��ƒ��MU�+����"T5sY�*�?Z(���_P}��� 4� oa�od��Ŷ�-�]�3+-B��.-<N�:���(E�ڽ;�[� 2-;�MWd��|�ֵ׋�fNv�̓���>��./��ڨ|�/��&��l��~?�������
]7"q�U0%��)���K�h J��w�^���9�"�7�Qcc��};��o¼��!5�<g"^̩�;[��H͌\�q�v��݆g^z�vn����n5�&��c�=>��ڀ��_�;���_��� ���ka{�Z�C���]�����e���>�0�D���A~�,��~ɺO[ɚ�i!�ngo!����O���}Pr�&*��o��Iz&��0�+y�u���kx�ʣV�sB���@g��VV�� '�A�[�?8��X䳟/o�c�]l�y}��n#A�C�;\���*�q��Y}.������:<&Bm�{��x���i������"��M�n�{��~�|�242jK}���Q����W@��R��	 n������_�Ԯ��)7�^i��_+� f t\���3�xw�ɶ5Gƿg@'Y��J��Ɏ�sސ.\������?�3#�S���F�>���!�\/C��9����#Cu�;`�����Z�*��>al��l �\8�;��:Yo�Gg^0���qbo���{��c�U�Gފ��C%�wa�&/�μO�8�pB!S��)~����[lH��E��k���C�i��	ڥlX�)ތޖ�>v:;:�G;I���'cw�)ͬ���+���I:$f[0��~��> K#X�Qk�Wy�ne����%v�2'fU�� �r�5W/[���x�T�?l�GGu���^��gۆ���&��|`;�z"S� �^	D��8���}1��6�F��:��z�-����z����?���識���ٲ7�<�2��$i��qj�]D����� �G��Aj��֮|�o$�kӟ�>]Q�PZ��V�"}tU���2�X]��,���/{û n�݊no&�nW[IM}�֎p��<ʁ	����e��5���<2nӝ�o,bm��ܬ��ड���@p��<U�0�rO<��W�ܢ�
�Ɨ��)��8c���{����;ԷcW�]�ҏ�{���g��4!�Kl.����;-�3� sy0�T�O��~���������U�����1�ɻzQ�Q^�������a�ͭ�alP����O��ƂL�p
r^��TsxH;S��]��i��S���eC��F!��dje��hd
>;��h��Zl�e�����MCy�7��X�LxN�ع8_V���~��޲5ݚ�"�C��撨l�=�&K��?ɼ�\l�=���wZ���X�f1�����!t� �\��vc�s��D� [��-�y�a�Y�j|��t���O]���������gtM;��r�+�b�1.����ٽ���Vv���S`4���9Oir1��0�cwz���y��0��pr��<V��&���Ć�-�������.�Z���;j��P��r�����:ȧ__rCx�����7��{��L� xc3��Fl_@�4��>: i�O�G�3�`J��`�U�+�ҫP {5��t%�Z����n��-�����a>W����\cz�7C�=�,�[��uZ�+.^xi�2�{���!���p�q)���dT�h���amW���z�\���\Q�� [����������>��*a����$cN	��P�^}����G�n��k�xC (,4):�ݶ��\[-�Kj����ވ�0X�1퀚xk��v4(��'�>��&T�����cc��:+fZ9���Fn0o��_)���(�~,~_�_��b��O��5����l����������aOb����b�m���s���~f�$�ϟ|����f̭\I�TLi#I������OC������״ϘΧW'�����ϭ�ë7���R|ac�J.�Þ �4����b�'�:�*7�]M��\��]�.� ��O�eLn�hR����\ca����ʀ���R	i���nĵ�M��II�+������P����Z����9�5��c�yX^�F1��M�ϯ��U�J�%3�񻳌�fe�o/ղ�4�w�����z����-�1G�ˆ��=//0�Y-�� ;{z��M�]uŔK�rb�&�q]�o� �{[�
������K�f	���k]v<���DgN���#����s���������|�浩U�X��<�Uk}�V���;d)�袻��ɇl�柟��W䲆�#W_�?m9��f/XU,��vA@x{5�ޥЭ�ў]������$&Fϊ��^�r�`&�-�	cۗ��44����6bW���	M�k�2=8�8�4�,:�0h���`��9xU����#�%���y&dd���Ovwl!�f�?{���r:��s+M��<m3|�x������O�1D���6Ff�8џW�O�/]q�����xfx�+ "zR{����Ⱦ�a9�K�^$Cy����`$��ky�[��Z�)��*��<�����-���-��B��)�p%��	z���$z��m"w`Ñ�7�?C�å��8Zy�Lu5�%�>7�s��O��bKO�Q�qk=*���Z��;$�w`o�����^>Y��y�%�$cgR�g�����9!׫m�^�(��=������򟝿���+_�&���U	v݅��k����^�Fz��tCmK"K�];�^���N=���"�M0* wv�n�N����7�����o�l��b !8���8
SL���om�: �t�y�gy�:/hF��L�MP>��T����{���[��d;6R�G�ҭ�U������vK܋��P��m��V�3ls��>����|F�����9����N�Q��f�aI��3A�:í�&>����/��z�#)���=_�_ьc�3�{������ה\u=���W�.:wL/�&!Ǌ�L����H�oC%WָH1���q�����{,׶Bw=OMWI��k"s7����TGѯ��h�&�og[MQ'-��"�A��5C�f6�p��O���B�{���q���k�#�u�9~�5׭&v��C0
��N;��u��):�[��^�n�@.!�|�y�����I�����bh���/]u��<���W�O�-�z���_NG;��f���D4R���e�z�F������ü��a�s� ����^?����6��|v�bE��뵭�\� ���m��钜Z���iO�T��zw��Cc5����S�/P���u!o_���z�]�DC�t%�)�"������ܝ��"�O��?�hC��Æ*� W�u��[|G���+��a�-z�d�jg�e'`�4��㳌�_��+���P�e1XU�t�ؼ=��CC�L��C���s&���~��2�=��hV��X� L3s>�ca������ح�xR�<��I\�;�Ы�K�fl��xt��Z��2<⮺��W3X���c!Φ�^~C��]�Un��y�je<�"�ȁ4�nV��d��
W������ssc�Z���tG�� Y��g��G�o�s4��C�}�r���b�=�@�0w�g^*�J�#��8�S���ң|�M�Z�m����o0�MkZ�~�E4�SM4�A���o�i��L��O���l*�w2:9
nTA����U���J�6`7Ud��~��~orٯb���g���Zo�~�-?P�	C����!����/���9�+y�q�$��b��Y}������UQ��M33S�-id���י�"�h�a�5iN�]��8���SSp*ݍ��֯�wPC���̽�B*���BO��g_�����g��[����:�����<�<=O4/Q�� ���h���^��C���xS?����]�hL.;\�!fХaU���AY��c֡C�81��5OS�)��xBz P�]Nzk�E�.(@	������%:��d�j�cK��s"4� �8��M�y��;:q�ۈu,C��@�����Α�
S&������_/a�l=p\��ՋE�xЯ>��\�K�1�0�?T�#�m��,��oX��|��2��Im�r�/{��ճ��1L��g��9�a �ֻg�>�;�G���!:��q|m\�#GF"vw6L�@x��t����,+�<�Y�E�������O.��|v���s��y�z�\���z�Cr���%�\Е#�#���	TXU��9�إZ�A{mi��\;�����>n�
�0އ���z�k��ڻy%�^�݇c(���+`�x�18��M��m��"+q����a�]��nR��$`���CA���4,s�i�Z�WsX�aʀ3���ǩU�Xn��b�/�6hw0��ξ�x��CM4�M4�L�"�#�>�wΝ��>����`�̨0t��T&2�2)7Go6�Ӊ��]�.��%G0�O��7�җ#M/mtc+{w2`0!��r�
��ϔh��T�>0^���.���r59�36"p������P��X-@��^�9�R�f�>���h����߯��<�ݚ�H��O7]�u�x�����=�b�-Ȕ�;7c����5���_�з��yOl���Ɍ�C	�@{�� 6Y���4^Fy�?I�C͜����5:L�?�#��W������*��1�N���z}h�2�Kս5p/|�y�-^��^��W���26�O�������ӪX9�M���B<�xy��Sie�YhY��b�d�W� �Tc�T�k����H�8���u��]�gr+��w�����=���a������HƜM�^��r���	���h&\و���MF��l}�(Wl	�Bqm
�1U��̥e������ l{�?�)���L�P��*�D�{x��UY�z�ARXP��{���{g]�����L����(L�s����Z�T���(\=������X�����%�QImkg�l�)��äꛒ���zcײ���Զ�cWN��$��=��wB���g��o07�!���Ô���}��9C;27�F��K��n�)^��ێ2<|�nZ��%��k����ր�)��@i����  DGյ�m�R��������=��L�7&Js�sıO����.��?E�{�[B�E�p�Χ���b�ruriDy�2l�2ٔ��3h��w�\�,V���Z��k�9	�ZU&~��DS����1�v��M�J�pca������H��7ͥ��C,�[��Pu�%��`YI��Z%����cL/��xN���� �rV3
�0��������q}_�|��<ߏ-D���
�k���XE��݀�?0�:=7���%�P��Dn�0��yRkUN�
u���]gB/r�H�CT@��������� x.�_�GW�4NZ;X�����_���f�����-�4��c�9G��@��e�0@�����x\�)78Ck�}b�=fW����^��[����VR��g�Z��)��*�r��VV ���nJ�;58��@z��33�8?s�}�W��X{����G�gFk��{��_�� A5��o�'�*[r���nNk��5�k�
���OC���?5��ʿE@Z�X�������ݒ��A��&��SN�=�/�}o�����
Y2f��Sz�rf�>3�nu9��9�H�f�Oh�[�u�Yȃ�8]�4�[Q��@��^
ŲJWp���Z�P���9%U.;�[�_n��%�7(hj5)��%�]�]�w4Xz�t�\����W���$Q��E	�i�Q��$@	FE ~�����W�����^`���>�S�}�,�����xPQ��,G��_�,}�}C�%���Z�]�=�.��{絛:�5��|آ��W�:
I��Hb̓��~�6~���3����a�N���[����y��y1�]�V_<VH�ǫz�����y�0<0\Kh(�Xh�E�Gu=�+��E�֑�'4ĲNR�dD�B��s�:�E�F�̩�eP r�Tmr�1���phLd)��1/c�$�*��&��s^f��ƁKo-����1壐��WG��"D?2=Q��
���8��J�|1	��7H���Q],)D��.g
���3�%���}zfly�t�bc�l����m�t[&�6 ĔN��
�ֆ���/{��6�̳v����sL��/avC�|����D#L������s��5Fk1����09tgw�n�	�*��ܼq!�M&5YD1�1���ܣ_7j ?�5K�0���^j�0�Y�k��I�Z����򸁹�w1�G�J�"�J��כ�h������o{��'+�]f4Ad�&K�%R��5\�<���jȲ���gu���R�ݖ�}O�Ul�¨]�&1^�K�m7%�t�m_R��qe>Ūܕ�.��2#�����V�;��T�k)��S�ٖ��9K�,���|tt]��!��')����i�n���#[���ϣsh���뷣%s�3���ո��% ��!�&M��w�h�x��j�]OwH���.���u�y+�z�ܩ�4
�Z�I)R��5[{�����QȒ��ϧJ�k����`����+a4.��YX�e�j��r�Ma\�9�*��C�{�V�5��b[s�w$�m�ib�e��j:�t�'�U5d�"�\7�m�%���(��K�9i� �Il]7����wZ4��9���iF�&�8#y��R�v�UJ��̗MK����w[j�rF�eW\�zx&��������]�r�F,��؆�YvzR��Vؽsjt�v�Oi|[��,_r˕>�DP�.w�"c9H>y	,��5t;�ul�l��N�v��0����qp���\� XQ;�;�h�cf�@�\ �=��V
x��=�ݳ{�q��0��ז��/��{)lw�����K�_V�j�C��=0�4�%e�kP}�v���[�b�����8��O��'GG}-Yկeĸ��o2՛�t�!��%���.A���4ors��Tx�%M7�Uᕷ(v���*<�K�%�=��J�������pU��l��
���n��H���w�~��K�����,u��S/�e�MKa�UJ�L,���\�!���I����P��	pѫ��!:
).V^�M[���yK��i���`�!�kQ�R��=�91�@��`��"��ߖ\�+��w�[J�r����������kX���|�q���vs32��X��Sq!��ܡ�����oTr�d�xf˵m���|s-�/��f⬭��+OoV�<v��f��$���wmiZȭ�����kK.�\׼N,�o>�맢ݬ��8���TB�[���V�<�;oM̷���������6�NJh՚���S��<��MS�����}E;�����x�-QP6���G��5��.�ޙ�lY�YQB�k����"w�P���.�����h\ۅUy��E�ە҅�=��q��[��Χ��Q�65ݳ�;�NIe�-�-��rcDib`X��28q�|1��ثK�#��S�f�0Ruu΢���}�"Z�����}�P���W9Hp΍�hY+�%̊��ӭH���8t��mo[r�s�3/Ua]��crm��]�]��]�˱qU沶Ec6�KrGӮQJ��(ٺ�mbD��m��U&\�Ҵ4<��Z���y��[	��P�$b�Sn]�ۄc�(�DH����PF:m���x��Ǜ�~o��|����(�)d�1��)+�Fd!	 H�q�v��Ǐ<x����BL%H�H��$o�鼑���k���E&���\۷o{�{����׏<x��ׯX�0�H$���X��Hh�FM�F"���)��q�v��Ǐ<x���10�"�Fƒ�j(M�EE!EMX$�	�h��~9� ѭQh��5���b��n���HI�(� �39��"ѧu�C(-3Ra"�0X�,X�ZQ$b"�!F���MAlnm¤�2,D�ɶ��F�6�JJ,nr#��/�D�;�������9� a�b��B(4�Q8�p"\r#?'�����~�.�2^�q�eG�e��s���vZ�v-�f�uSE����8R[�h�ؖʹ����c2J(DF5�6Bp��$ ����"iF�-6�"bD��cRQ8C6_��5#�T�,�M�d���2��5-L�$D,��~���A���$�V�h@)��dU�A@Ud@�^o��������I����V��>9��2��G��cp�i6X���=�-�࿥�Wt�qG���{��N�W��BؿX�6�r���\��-6q?�:��9kj��<�.��E�z})�w�"o�-QM,z�Z�c�U���[�w9��gh�ϦU�d�L�@l|�f�oD���@�S��
��q3K*�Dv<�U���J�e��o�k�+��~���_ٚR����1
����-�����
��qD�'2/�hb�Zz��瀾����w�4D�+�Ǉ���];w��Uo�w1x��h�>�s�;1j	\��Q��y4ʺ����N��mj��.��o`�
5��a�TdT��Z�o�5��	�*`K�F��.�)�ׂ�+7�,|�v�b=��}�~<��<�1 �|��ύ�7�,�kCz�,J�B��ʫ�Sv��<j��[�9	�:�q��O����?N"�z}ИZ�-Ɗt�בޔĹu�{��\�D��_�P��$���ffڶ/m���y�[R�AN�e�Ts��s�V������A�P��L?�U}��y���
r����Uڕ��@�}��:�\���aS2���9��S{���E���L����m�p�-�c�f��Tr����6o��pfC{�����<�ͺ���9�s����e]ܟ���m(� SMZ�۷U��n�[cj�U�	D�~�t�����E���7��dK���%��¼��^z�[�0�p�{m��$��� �}�y�'ڧD�Ὕ>#����y���=�&�[�g�-/#k��W"AU�E������\�U��eg���Ȇvg��ێ���o�OW��7�P�O<Ǟ���^ʂƗ�S�q �>�k%xǡ��y�l��JЏ64�"m׆����\V��E�]<�n�k	�gK��&�uyj��xm{Rdt-��Y���&�, k-�"����qC�Jײ����g�R��g:\��XWL�yZ_r���K���ϒ$�wS�&�/R��ʳ ΘK�)�'����n�U�a����(ǟ|ŋPg��,�#	��/~�q{#&�_S5��~��^j�F&n��,�\�f�~.	���1eyMQ/������Z�_ǰ�U�gr���dR�_�Y#�͡1OꃿX��O�����.4��Oe�wvf�ٌ��1���`j!� �Eך���ס/V��omp���	zJ�!^Dך�%�;���SA'H��U��|�O=�j�̮{�����^웑3�X�E�Uˇ�7ww���|��,8O�t`[˭�Q\B�g����zE]^bݾ��I]
��F��`U�1:�ז��ɒ���m����q�z���Wu�q�{���jkW��?��$P��i�@)�� �YYG��a�yή<a:@��;3GLz>.3�!�|��s�����5���W�gZ�}�2�E<�y<��d�oW[��.�v�ױM������5
��Y`X��A���KFO�n���e��Gw��f��3��/�������J���-�+��3��-P�(�ls�<�`&�צ/7�ZٗZ/Y;u�^�1��%:��Sߕ���v�E^+��
�AJ�b,��O�Y�q����n�ֈ�'�E��moC�^����\���L�@�u�.����\ �s	�\Ymݘ�,����elr���/Dki��ں��.�7���ɽR���LV��9��Z���&�.�ѐ��9օ����S"2=�G7P�	�lȓB�����=^�3	��~�w�ᶰo:�/���@gMsۂ^�e�~���X���^8`|������4���+{�W���&'�z��Ŏı[̭������}�q��T��a|��?� ���#�� C-�7�m�0^�탔Ύw"�͞�I�z� R� Ϫ��ٞ��>�
����$N���N{�k\��'���OA�gx�&X��;O1�e&����ī�7L�y�b��Z�A5Dt�Pl���ɤ߳�f����{H�Ęˊ�i�b��=��r�K�g7Y�OrIYc+��Yy�k���K��=�9�����~ �$T��i�E�)��R�iA
i�Aw�����oo�/���`P�>����,�?�֎���q��۶	�h������'�];@��!�,f}���/���U��-�m�������"����o?\�h�}���u�Ȝ��u���mޢ�ѱ��S�����<t[<5�W��U���r\���4$�CNWX'Ec]y�{B�Iy�_ʢ*htK<x��-���$��O$��8����5n�aw�Y��5>ð���d�A6���nm= �yVS��O�K!�7�qi�?��`�{b.�r�`��b���#�f�
�P������b�d?fͧ�{gM�%ޅ��g�'����v�lX���1^J�g���!� DB�:���jZex2j"K�t�
���[��I{�f �_k�4���v�s7���7]n@�:��Aq�bY ��Ji��F�W�n>753�x����-�wt�=���+@;��D��w�eD��$p�Ly�LK�\T�c@�I����:R�*NOm��c��qp�o�H�`kL8�/��X-��qú�$��7�T3����ւ�e
_n
�F��ewJ�J���`�F�^Й{mnw�q�]�T�T�u�)�HK}|6^m>�}o�	U�BԘ�Vvn>�4't��2����]ң��c��ʜoE�e5�>�[XbJ��'�Qu�j��AO��E�iUi����hP!$A ����%ߺ�W�k��f�����U�h�GP�Ee����a끫�/���^�52k񘳞���M��i�!Q�!����86ۇ/u�\��<5���p�p�S�;��Z��͋�KH柷�^�Dw ����~kÐ����u���5s奛�'�ڱ�e�
�rp�_��y���{�}ʇ�o��+��_�����:����ns�s/e�'J1Ȉ_P�a"�P��Mw��]��;� ���O�`�ʡ~tA��2�)��C�W�uz�"PH|Ȱw���L῅�w<�f�q��O�A�曮�r��!�`:�?�x�z�ԕ�Y�<2�'n�`�pp΄ssL>2/ޱP��r�d��N:�/�L(���q*�:(��E繩�g��)z�4�F�Vf�g`��&��-뚁������/��6�I��*r؍�uz��fC2i	)v�E�s�9��\3��-�������]�N)�!��#F��y����g����(M{zO=x�>}��-7����=������*|�c��X�K�4����S����P�N���5�]齞Z�V�L��i��-�?4����Y��Ϋ����7Q�<����-̺���)c{/��fgx���+Yٞ�/yRԬm�_��RM�Tk��?�/�CĎ+,�I��6mR�bV�r�$�.Pd�mV�օ>��Ngj�OiX���D���Ǘ &�����b�<	$M���ƚd Ji�E���iQD�r�����o_h���Ú�y�=��
�\��r��s�5�zO[�%�����x~�%3�w%!��lN���"�߇�%Oz,9�4�A�����&��Xs�����4<�;���j�>3B�(n��G>w�;�K��=��J�#*acȷ#�	��"w?L]0��|FlLV������ze��)�QO>l�N�0��Шt�zC[PN����+�bE'�����Qy���AVOV�(Ą�g��Qz	q�O�|��O�k�/mp�?^I3�z^���G)�(X�f�ӵ��NKש�9V�}�Lo��\�:���}�'�]�=rs�R�gO��W����=�J���W�םI�fA���rQ{���ơ���qٶ�U8�'4�n�����]�s0��r�%�_e�:�=#��x��&|���k��L��4�gK�˶W��T62�*KH ��B�w^�kǳ�b��^�J���qC�Jׁv�t�%��۟T?�?\��ސ�k�zgVUr��<����6[�D���O��a�R��j���i��:�Ӽ�]j���~~�+�Yy��>�3���H4�2�U�͛z\K�����gUB�vҩ�O6�;�3i��z!��u�k�nv�V�E��4�jW!G\�!���X�wt���Íq��ܞy���<�����H#M4��M*24�"�(�
��� *H(�(=��|M,�n��Z�?Mk�q�F���Qv
��``�+�� �����?�g'�Y��Y��a+a>��>׳�^0�� 3Ȟ��C�&{P��aix|<ƽ�x�
����:�	��<� =�n�
���4U�r���=���~��~q��\O&|t�M��{��C2�p&s�'����c�R�oMV��*�s�U����B�&��m9��ۈV1ň����#z�M^?dv��V�W�i!��1�L���-�r���|rj�3;�7b}P�f��Q��V���� [	�ʛ��ئt^y���qsqI�d��8?&�Eٱ�ջ��r�l�d�Ȕ�+��{�b�Ui�6P7��>g��H�Y]�V�u�q����֐c������	�b�B�"����?S�n�$8�c����4p}1֝~�Y7�𰾖����Y�D�S��(���D�NF��)K��U0����s�ꛏx�GvyvAz�@��Aa�"�y]=�T0�;ȭ�e��P�S�=[�"����.6W5�o2U߅Qp����}�5Ao�6��w�z�d�N�C/num��dJ2E����[�z���X��b�o,�o3�t��}�z��-��ۂq��y���p��w>���UԎ	a̸�i����e���*许2Su���d�\�g/,�@
���M"��MEhڴݺ��U��k\�S �H���� }����w��f��,G?�r!6��y�nt;yI����L����k^�EM5����M�d��d��T҇d�9c�q-���h���cTW�N��x.��[i�F��]|A��m�Vk;��q���vm/x�#9�,��@1.�|�Ћ��� ���f�ﺽ���^3�������(��!��'�/cŖ�NKԼ��Cb�l��tAw]��(հ���l �������ݮ�lS�#u�4�_��׸�4�v�O��O���3OXU�dE_PxU[ݷ]c7�����$~9�">Y-�m�@=������@�ޟg�DKs��ɕH�'�^����~NY|��vm}ʫa砣�J[�H8Py>r�<
Q���]�{W��)xZ���m}��U��e�����tԘ(�O{�"�{��yYBj�7���];B���~�q��Ӛ�*��f(S�a��ao���	�A{�H�)�d�v��lOY��TfW�z��9����
[A�b���2:E$�Y�~���*�Vj��b��L;���a�Yݽ]b�y�/����۸)�d;�c;th&�����7�=n�2���N�
��b�a�9���k�V��&Ϯ���y�م����I�9�&��60�D��]t0�n�{Ɏ=�}�^J�%���w�1��P��h� ����ƚV��� �� xa�8��׭왍U�[��$�w>\Č��e>y�J��j͛���w��}���af�|�."S]�;�A�XbS�[Ӭ(�ǫz���nk��b{+wh�=Э�r�Z~L"X7y�w:�o�����^m�Ԟ�Ji��4*�Q���Y����4��G�`���v�2htϏ>k�@0�q�EA�N���h�.�"���B���Z��Q�W=��}[W"{\?WG�	�d[W�)��5���='��$�4���p:�jMk�;����M�(׸�0�b��|�>���	��'�$Jn������Υ�6.ͫL����e����~/I��G4o(6��J"~�at�>��Q�ׇ_�#��� �m�aF�@�^��G%s�z˄���u�����������!��9#���gn��7[����d@�s�[f7k��zN(���͊S�U23^���f
02�� �^���<�׼ᖇ���y쟋АY�O��r�J�?N���tk,rz==�3�G������/(bks�
��A��C����Зd� Y��/e'[�Xe������]y众�mm?���I�o��tֲ�lZp��j��k^��(�T�N��9�(\�q�Ye儙��t|�������a.Y��m��R���^W@,����Xu�3�mr�N����ҸMM�۹���W�@xxOu\�mT7n���ݻmWn�j�[j5�E��ѵh�A�Xt�hD.��/
=����5"�C�+�<���p�#��&J�5�L����
r��Fm��w@�ޤ�bS�އgma�<��{�<un��S����>ǜ���q7S2˭�7����֢��Ǟ��	��E�4rn�l�={�m�֯PvМ@�Ȧ���I�@N�y�O���-��hcx���a�y�\HdQ�י�[���gO3�Uֶ���b���7\��L<
|�`c��ޘW�}r;��8˝'���)�P��!����e�r}E�D�c�"۪9���=�d��rÞAʇ��*��l����O�[6�uV����cw��&��&����S���qL"�rޱ�Ⱥ�I��ހ�Al�;���&ݮ�(��5�t'$	�rR���)žE0�ȶ�����趔�8�C�C �۱ć���}?,߾d꼑 �5�,/2V9�QzK�
}wʒ�L����y�`W��w�[�xY՘�y��=C���C�S����b����r�v[�;Vm�s�}�����j������_~�J����1+�rn��g��ce*��]�q2^����ʜ���o8��
�n���u�uK%S�-mm
��]�y��\���=Mقm�������4���oqZXM�� oA#u��Wp��st�h���b[��1>���+-ڹ	�k���d��l츘OK���o&�b�n�Y�H�-s'k[6�v�d�7d��0����ԱI�K������v6��C�,���|�Hn��A ݻ��su�ካN�3�l�V������2��J��#I��s����v&U��C۱��N-�;��{��9j�^�.J�i�.�b�p��b�خ�
�w�٪3��9c��Jˋ6���M���R�xn��Q��r�j��ֹe��0ֻ®��$���&��l��9ES���D�]k�ź�Etn:�GtUM�T]F.��N}C������=�KЮ��ǈ��Sqdu}�t�l�s%ackx&��>,u,'����SK�팜���	צv\ۚ�	y`]ǔ[Ds���̍���t�K܂�ӗ,˨t=F�c�nԃ�b�w� 	���W�kia�K��ES��+G&�X��*c��e�� ��K������	�z
�4��#�9e-���b��U�w���4K��Oaw|]��� ����<�iu�wk�a!����x�"�Y�n=5�L��ڽ��j��� ��a*$e.ZJ�n�a9�F%F���g�h{YN�A�O2��٦#Yz�'�y9m>�?�����r��h���Z��۹*�P�=�e�v�G�	"F�m!���w�u'd~�M�7�H�'Q��w�����x�+v��o^���s�5���#	b�h��������i�L`��5����A��ꡭ̓oOh�2P9V3��<PZ��6���v5�nj[v_=7;��O-�eJ.�n�b�}ʊW?����J�'�g'n���k1n�b�j���g����l����,��n������$�"W3��ȭL6�'�x����	
�T��X�.��@�,oj[m��o���$خƤy��5%A���9�٨4�#*�pO�n���%�	�p���J#V���+�N�I����Wt�U��
�gmmpW�!'c32�؎D`%����`��4��2*��^�;�wVr����J>��%���q�,Ì�u��ٰ�o�2��+xtR��j%���y��yuO
��E��t�@��Xb�%����T3
�_<}Z�"�s���ɤM������P�����̓WX�&�r�y��v7Pg<p��G-Z��$fh�:�WmCn���-&PT�"�6*�{C7��T��ە5|@8q-=g��M|��3<�v�GH�J����w��͂��A����ˍ2�eK��c^=��n��\�;)��!��S)�>��_}�MAV5��b�o��d�����6y����ۏ^8��Ǐ<z��I$O}�^��r�b�&��ʕ"H�T���n8��x��Ǐ�z�bȁ! �
� b��o�4ch�BA�d �cm���<x��Ǐ<z�ꝃ#&@R�pbŐ�-ͣDQ������zq��x��Ǐ<x�����D�~+r�ەb*�WM{��b��7��&�h-_k[ڼY4D�nj#j*5cb��n[\�&��V1%R���.m��1%��UQ��4cO;W1rܣZ6�X�^.F���<⢌kM�h�*-]����汷.���We�\��9�Q�a����#Rs�;ҟ��K�k5�J�ʘ�n[�Wr%���RaL��f����-�ꪾ���Z���Zi��F�U
��#"� "�}�k_��?5VT���Lߌ1��:��K���"M4�UvI疫7(����X�\jC�Q�T��1'�^�I��;�&������K�M��.��(��^��I�+,/،�S:�aE�Ĝ��\����_�4��x����ma@8P��`c)dR��<\oF5>1�e�PO���~���Ћ�@�g��� Xʕ]�~�~$�� >'���5W*��Ô��I�|w�wZÙ_C�tM��vE?�zi�3���4��]�m�v�|�}ЪZ�N�MR�}Ba���`; �Z���7< �a���:"X���_Z�N���|�f������)�����О�<�2;섄*��ʇy�;ǣ0{C��z����3��?FZ�xjB�3>��	A����$D_�T������ԋo��W!i*E�efS�n���=�����Z��SW�T*�C���*�	����}*3F��0�4#��LJ]Y�}����A�����u��ǵ����0�8&)���j����#�S�"tv
�L���f�B*�>�Y��6�n�%�3uv+��؀f��}�Ӕ1�8.�z�H]�@-��G�uf��ʒ��xw��r�<�Y�=�s2�Ne�h�LNk��n�v;�y�!��{*n��;qG�ٺǙ+��0gN��=��=��L��u�d�~��	Ѡ�i
�c�v�j6�v��F�`	 $Q�uϦ�}�>�ߟ��6^��[�	��ZhRxW��5tf=z���;J1�k�@���mP�,ݎ�"{#�Q�1�!	-��]p*S��R�w�ɼ�F�3��|wW��uث~Pk���)7)����g�[����1���ƿ��~�W�z�[�x�)�ڢ��H�I�\l�8��3Ӎ��B1�"X�Z��k ��2Xny�^�r�=}%�}�]0�ʥX9�Ҷ͗hQW���2t�r�p�@����_&"�zHx��	�&���4/�;��3��S�*�d�֫��5W+���r��9�|N*|�~Əǎ�z�W���>#M�a�=�L�ӕ���5v��2a� Cе�(C��Ax�T�b
���:��?4ڸV�Naj9#V���$�b���hl|���J�)�z�#-H9��l/�r+�LH��P]��Q�r���3��C��i�f�y�tS*�46��S��[�}bԉ�ny�؏N6���k���>����& ~�\s�'�2�&�������:+�����[�>��ZEZw�Y'�vU����{!�h���W�՜��v�R���^��9�:���=pr�rrS�r��w�qۺ3��<���斻ⓢrID�y�nez�Zq��%n)�fJ���$�����c��<è��v�@�opwͼ����q�v��ȋ G�"F���i����\�+IX�Q�Ed�R@$zM�ߨ�5�eo�w��[̪�x�#}e뷎5��kG4%�����C�gw!��f���S��_*!�/��Cf��+QftNm����}�9��>�J�U~��_F?�\EC��D��"4.9��$��z����o����_m��}�������	&�@��z�ʀ�-31B����Q��X����m�$�P!�1D���}^^8�{�4׏X��A�.�`Z�7��I�l	w�aŶpkj�z����Y�k�=%�-���!5i�1"K�+�XE�p�����E��}�TM�+3�"��|�5`�a�"O!d�ٱټ`P��=��۽�4(W73�C��oDW��[H�QύML����C�G��qt}U�R`��Tf9wLI�q��y[��%D�S��7�I~������ ����kgڿH�{�\(\�$Δm��X)ܞ�q��K��wXD!�\d�w�������e��"���sW�1e���<�l#��L)����\���W�4j2���i�>����x�Ⱦ�h3��$�R9�iy@��	���1l�<�=��#��ah�6i�M�8�f*�;��Di����m*�6���fm������3�N�p����}t,�c�Q"�|2�	��oK�c�[6�t��ȵd�8��o>"�%����v���1l�V=XĻ���}�7�?�@���5 S@4��E��j�F�kM��la�2�L��
fT1ó�[�9�W��P�^�^��cS�:kw�<��[;�e�T;H>�xݘ���)��|��t���|���6\n�5�B�(B���b��T@oc�t��kT&���^f�� �R����Z`����vN��sfZ�F�������=>�pxEϽS	.f�]K�A���AC�����D=�<q�@\��!՟vz��I,����ّ�8�{t@]^J��'�r���C��<3������x~����L���{wf%oc��+A��t�Dħ�q�ni�0{�U���6�����~ю��kn�s��ˍeJ�w�<�k�p�j���Z��^�TB=0ŵ�>uz*�N�.�#q��#��wjX��`~`��ܞ)Ǖ<מiB.(fG,�B��!�^M2��V�d��v��ُ������o�$0 X~O0�oL+�p\SX�'Ƶ���fj������N�3/m��+��c�G���3���DT9���V�b$��#=Λ6�}h|����9��d�	w�ɷ6%�m.�`7�+�Ͼ`�o��Yǂ�B�-�VX�=�����:���mں+�y��Ë*'�Qc�zS&F���x���	�B�y��1d=��.�����z��Y��oPa��YL�ƯkG^�>��N��k~���n��z_������i�*F� ���"�� �����%y�5��'�;]�qmfrq��.E=���J��a	>�6��3���zhe��G;Z��*\O6s��N�R���d�b2@��ȶ�]8މm3��NeN��HQ��f�2����=�*����m<�פ�Ч�!eS�VB򒤥�y��gg�b��d��k�9X����P��*`p���z����۞Ozb�Y��-/������p(��~�yz,�'V��w�Ba٩��q���V{����N�lv/��s�{*��:{�����§�f��u��ޟ2!Iį??��!q�c�o�ӁE�I�b�'���	TX0��j�|=��w/��՝����M�G�yY�9ROP!�lm��M��o�����^3&3yh��y������.2�7���/��!�����^O+��>�v�o�����6�q�L�Ս�i'^c�(j*���{������v���zi/A���k��6ƎԵtL[^D�A����R�<F66�����f��ùߗr7��{����W1eyT��ܑ�O�G������*|����2���ׂB���)�����'Q��?=��`�qf$o�=�na!e�ŗ�}�v)W�h(��v����Q�VΌ.�����MIGH��[���˩�} ��r��]�������v���`U���M�]��Mۭ�7n��v��������_�}���}�_���1��@��Y=����*�@^L�w\JpCO�����kk�0���K̋���;��)ᯞ���P$�����߆�n}ïxzj���]�pyOl�v���\#�&��;�qZg̮2�j��ڡN���}������L:���KT�o�0���ԩQq'���}^Y�:���^͛if���׏݇���\=b�0����"_�j�n�]��y{W	-z`&@+2$���ǳ)3u���B���0<֯�YW��I�SȔ)��f��W�4ڍmr ��M'XSzS�[�U�{gO�	���{�R��'��:-��x%�9��pS��'�gٱ�y�X����r|�ݣ�
�ot�.%���p��/t�Ow0��X�[�.$4������|ފ.�_*�]OK����vz�W�ǣ/SƑڋI��R��-@ܰ������S���n���;��A�䪷��ֱکv�*�B�/�_����a�'�\>ߚ=��|p���?/�0����}?�~gX�9��'.q,l֜烑����CE<3x(0Q�2�Ot�H�n��v*j�T������씞$H$a��D#�2��
���𵿹���]�F V�HHÒ�U�>��;��0t�؞�K9j㎧u��t(v!c��J�cwUJnݻv�Wn�1$D���$
[���z�,Y+3��������[t�?*���V"	'}������"���?֣X�C��b�����z�&���C�,3E���F3�D��LK.�L��YH��L+��V��L]/_�_鄏��@TD�`������9rb�*+�����a�:i�f�g�QLhF�)��]FA3�Ǭ�\v~��'�V5&�������3�*��き���mO�q��FC_,�ռI5�3��>��+�%e5��[�]�Y�ӯ�͟�yT���gOߺ�E�M&8.��A�}���_����������[�|��/~��,��kX�/��WN��$zk��'�l���k�6��1����1���*�Z�B���tc�]�n���郣���(MwO;��sB~�z�ʹKL�P�a�$(M�)=*�v|�ħ���-O�m��z��έ�-��f~�Ȩ�pX��iy�iֽ���O^��sˋ�u%��)�A��:�)�\zdŰ]W>px�Mza1"K�+�XP����lǾ�3's,-�D@�8�μ]��qk�"X^z W_��@SY��܂���t�
SL�q�3
v5N=S0:º�>�w�<#��͉���J�i�W&��!ֵ���0ȳ������.b��/���A�t4]ȟܪ�UK�>�oe}[�!c�	g;�\�B���;Y˹v;6Ԧ�l�3��u�6���u4Y�l�oOd�{�ɿ}�_3�?=Oƚi��i�������I���!"�;���ϥ����1z՟�++�����1�����$&�4]Aǟ(��<a��+�gk+e�ǩ�{:E1��&��ۑ=�p깣� ��t������}3���5�Z�)�Y�/˩����{x�&*ۥ>(��ǌYx|�<�`��(�yȆ�}���"��f���9�A��hׁZe�oa2��LZ~AeK������v����>��V���@�I�;k��Fܓ=P��̄?�D<7��ۗ��Wd�y�fBcEw���>;��# ^��سj��ǿ�T��������"q����vg�e�}�qM2�+���ی8�'k���ҟs�!3��k5�g���o�-H�|}kH5�����z.���.[&�E*~�a��Ygz6xԆ}ū��y-�=z��|نYQ�:h6@�5�V�
���x��a�ʄG��2$Z���'fl��l58�F\Z���0�߉��W�ԫ������T�����C�+~�C�F�OE��J���B���O�������y/.=�3�r���鲿j��b�����_1��>I.�}���(�����wW{:.�<����n��W�+��f�#}�˜�8]���b�^}9�][O&Ǻ'V���V�ҕu)����<��Ozc����v���V�U�S�cbU&ɛ�rM���z?�ƒ�!j�i��hj$Q� �����������X5k�����f�L�_�9�}�۔^���HG�K��i�sͼ�[�c��Kk�k1�����p"Xg�&�-�^D��*ao覥�.4NG-A+��2zc���n�yV0-/V�ߝ����M=?�{?�[���O�7ɶ�Г�X΄�l�z���� s0f�{ȇ�
5���56'NhK����k���\�l~�KO���ƍ�I��&^����h�3n��x� &U内+�\�w'
ꋇ�{g� ��4�22c����"����,�:ݜ�dj!�M� �s.{�N�RS0TC[�ɶ�Шt�zC[u4�`���]VWfQ.���N�9i�T)MǞd��Nt�Р���f�x`����Sn�S�m߹q��(uz�:�5-��ʷ�ڶc���)�V^k�x)q����"o��YǸ�l��J���nS�����%�L"�"8!e���}ʄ^=~a�}I�Sv8�Qw���8ɨ.��z��Y��5p��b��|��F��0���{�65�	�^:��"�_P�����8����S뎆ڻ�����Dn�܎��|�����Q��E˹n����N����0�Vؘ���lD�0Wa[�'lN�ޭe���p�g�q������7��U�pP0���MA�qS�0b���Za����-����J����SL�4�B4T�H{{Ͼ!=>��T³�X��k	/m���F�`�|m|����<��n�hM��k}��ܭ?CE���6+�������ޅ��*;��}���"�U��,K�4PC��&_��9yi��:s��O҅��=9�����3�#"�[�4�ޓ��z����|���P�=�x��T
�0Iy�lp��Q]���E���![�;7'�f��i�½�F/�a�����%�ȡr��I�De-�uy�u�.�8l>'� <���t��۳Q@��v\�w*���ou
B^;2�+νM$�wPʐ�c�҇�@���+�����v)Y�4o�po�E6�J0�3���Õ���\,�Y�!
*�[�n��}��#�G�t�N�eYx`�y�6���ӛ����$�B����aC���+�M���'5�zDͩ�cQ�r�`�1f�����V?s�M�g���y��hO:��r=y�J`.ƙ�L��
O~��(x�x��[Խx�\KA�]��i��Z�{Kt���*|�@��2�n�P���4�gR��7��~���i3͜�43�R��OfG�ua��ή��!���V�Ԥ�9��y��po����$��D�7o;*�F���A[���e]l�n\mj<;�g���Nb���]u�t��7�3�H�I�u��:�)�-ևX���p�=�u��H%�8���\�[�6�LQ�X������������8b�oN�����h�&��:5)���t�l����jʒ���^�4
;(f������r�Nچ�[$�ZcT�.����ڙlu�Q��2,���l��Q�D=�O%v��ש�0�ڃ��F��6�X�^WW�b=�r8�	�2�T)h�y_y�����Jƛ�y��Spe=Էj��4
�p�]u���oD�;��aEQ�,F�zƣ�)U+z�J>���M��W6s��K�����Q�Ʒ-q8�QOl�X�l`��"��h��ʥU-�-��ݝRs�C��֖&�%N��ȡ�'&:�����n��{XIW!��q;O���]/���S�h�,om��+|�Iz$�7wbZ�%ۧz�5� �h���z��}1l5��^���|R"�cY�4.W7Ob��mh����#Y���L�vRW����q+�tR]Y�^
؂4]G���ok�hZx�W�s���8�8��_f�T�4���w����P�'���>��G���}S�qnr��<
WSmG�b6��K&�qQ�^�GޗB{;ڒ�d<��=z�5厔4k[�W?�neqH8=>��zx�=���>C*�򯺻w���n7H`��U�J��r�=����C�E"�`�'ie^}���RY�ie�e {d�S����\�w�T�L$e�¬_!��5 �?�'2vK�����Y�a���a�G]�\Eq5�+�Q6�P��}I�
�cU,����ȳc���vG����PYE�d�X�X��nb�D�Q���PC�[�ٸ'V�OP��䌑Xl1fr��w�b���#�WS��^I�f�f޾q⇵��鼺 sA�L�Y��̆�hX�8w/Gu*��-�I����`
s�1�O�ȭ���8��ޓc�^��I:�ƭ��Ψ����yrF3��b�������He��ޢ:_,Lu��\����֮亂�Cy��,%��݌�իM�z_k�jF�4`2��»����)n��SW6�;��;:���p2�x�<|L��lɳMn�q��i/�iYjsv���#ͫ2��,��LDo�Ovzf?o^v�u"�+����{����Qd9���A�e_Gie��n�=3x�����`���ɐ�¬�b�U��/�TҨ$6ͱm��t�P`�7I�s�j�7�؛7w������66��{W���ٜ�l�VU;OAv�I+�;u$8Z����*���Ny���zTV�E���m�cb�m���͊9��n Tj���^<q����Ǐ<z��bB	9HbSPn#Q�$SW��W1�άk�6�Sz޵��<x��Ǐ<z�����D�FK~wd�����λ���UE@�a*@�m�o�8�ǎ޼x��ǯ^�H&�=�P���\�E�hւ��DL�5P`[�o�8�Ǐ�x������m�;ŮksQsQnsF�������+�����5�nnN�ۜ����_J��-�΍Q�^�m����x׋W��5�lF�:V񫕣Xۚ�o\�sF��sh�QQ�-ʢ�+��coT�#S��r�F;��s���N�X��r�˕���Ѩ���n��(��*B��1�c(\��&�ȃ�E��I�E7�:����i��x:�޽4�Z�u[q����mQq��fi<k���f2���h���wf�,�7�\�-��DY	0�Q@�$&�0�R���.6�5JS�X�\P2��HLa�AM��bJp�4�u?�d�m$���(��5Z�R�5*X���.��KK��k\��J�7�K֦NW���˧E[ۙ����	����ߙw�!�[:}O8�����{�/�D{����89��,Sި�sZ��?*6[ �����]�}���>��Q!]Ǫ�j�.�IM�Y�} ������*�8u��Kz��/y��~����'��x�5�՟�_���Ew�/~����"?��O�&�fT.�3\�����n]�lw�V��={�Z~k*]&�0��K]�Ly�� `�s�֟I��:y�Vҳ:�*5o�ᕬ�.��x�/6a�RZa�F�� �=�s�Z����àC��и�e��y��(���ޡ2%���0��ek�*�O4�@52�l�F���]��;�4�8�ΛA�!�a��)������#���3�7��<���Lz1���9��D`�8��Ŏa����3S�`�p�Ht��^a�������Am�(���*�ɲ"D_�b>����JV	;Y�(N�7��iP9P�{ߧ�?/pT|h]��CI�า@���Qe���6NHl�蔮x<^k��dxg(O�jh�ʡk���'�A}�cQ�]C4�E�>��c��^?|��ۺuN�l���e޴�Ά�����Uz���H����󱪃/���ۢ��k��u�WՕ5����kb�g��Q/�W�HI���]���*<[��[�a�{�7gt@��sin뢶�N��]f���3��,`]�y��o����bF*�,��y�����m9��w<�}W["ovS_��\�	�6�/���[�)�|a�^�i�ﾼ�~�)^�'�A��F�=驎��Z�����Y��FoV'�k�>��e��z���?`C����伈���(z�X�,�͘D��e��WjWO0� �+ߓf�.����C��mp%�������F~�>������+LK$���ɞBP[Ճs.�q���*	�縰��d�FҸ<����?&mG��4t*~�2e�r#)=���3��E�d>DN�*}!��F�mb6�Od\:���`[LW��^��˚�����B&b�Q| �K������w�"�i�p�VQO ����槲��sQ1e���<��a(�T����r:��Y�,Oo����
�.�{���O��L�sNr�m�g�w8��t�,E�V�k3�ǌӦQaC�؅�!����-�zhU�\�B̄�������[�C�e.��^��I����;����ܔ_��d�k�)�7�k�������0:�ƨӨ5�X�-�k�w���m�sM�'�m�ǁ�;��E�30k���M\
~��jY �Y_�z�t/��%)��Ez��,�Y;�g3�G^��;7:��N�s�}N��-;�F����}�[#XE���D�`�|�{[ֵ~g������,c��n���	5�tC6y{�3S~ey� z��p;�+y��͟�؋N_�����5���q�������^�^j����B��~����D)p�"D���!�>UY���K��66%]!��y8����;C���A��NZ��w�4뼼H~gj8"������F��e>�c��P�&/��(w'<������C�U�����տW g�kӃ��g��ٝy34��1�"&z�3�]��_�<����u	�gI/^*>G�h��lO�oe��I)�1�T����f�"Bd5m���K���॔.'� �_o�m,��I��;"�.��vWr�=n���݄}R־c��D�X��,/|�����8a �z�ٽ�'�����R�"-(��{V����N��a%�5���ҳ�c�u���O�����j����1�7qb���-��:v2�7�}0�-��; �,�o��,t�a�jP%W7�5���'�\���m�����|��t�z��x�ަ�gF��Z��r������ߢK��A	Oz���6���	��h�����v�|��#�L:�~6��pUnN�E>�&�rwn��eJ��"˺�]t�|�yk*����8'�;8�8�b���K«쿫�~#0�B��J���N�'o��S��|�`Nۗ�;k�3��Л��FT}�\W�֝�u1�Q������0#0y3��o��'�ٹ��ۃl�����)�@&9�x�'���/QX�����gn���UR��Q~Xh��uႫ���;���v#�-�2�ެ�>mG'��d]`�Y���ΖE�鯰���݌b�}XF��H;_5^L!�Մ��̪���4>��K�s�W�m���n�;�n�Ay;"c��t#]J�C�ީe�.5%<;��|{��`�v6>;ɗ��	��_��8�^�u�^&x�{Q.
��,-gM{�г'�`����~^*�*v�
N@BZ�!?�i�"j"�5�S��ʊ�խ�C�����zV�$�K�B~a�5�־wȎ�6�k�\]C��ި}C�n�w�O�Y�����Er�s�/}��.��	qc�Cs�q`d;O�C���u=<F���� ̀��������c݁>򖉿�����;���!�`O����vfL�*����-k@\���O��Rc��4�E���t����HN/&PLV{��+�g�?~��1�N'��[�*��R���mg��g8ᘉ0%���/R�U�Iǆ����ퟜ�������KX�ۤ�kk2]*�!��P�6���'-���$��]J��W;�"���h��쬹�6z�\��Ku�'Lyv�#;4�Wkv�5���S��nIm,�&ql�+a�<M���\�^��F�*I���Ѫ=�1������z�=����e���.��/��T�]���Mz�����]���6���U4 �|e��g:;쐆�Q�4���M]1p��y�����4���Q��2l�̝��g1�G����q\��틤[V� Ǝe�q������c��W�,��3��WNQn;���;й�;�s��s�2C�o-k�ʄ��,T)=�+���ǫz��7;�7��,�l�ɘ1�j���R��J5��l�tJu~*K��鄪�� ��֎�2���_VM\;���>�^��Jj�m���w���W�?p�Y��?D���%�8I0T?��X�]�������
}w���Y�C6q~o�4�����> ���|�^ѐ~�W?K�ĥ�s]3jv���ɛ6��޼Ku�Ag��z6@w��Іǡ�B�?Ky�lşp�W�t���qg�����r��;fq�O�eAbޠ�? ����OF�^z=>>t�ؕ�J�o���C%��!�#}ÛFrT.�4a��F���*�sז@������-f���j� V��lb��l���/0��6��Ķ*�.����3���u���إ�D��n�]e �^ ���H�s��*�_��zܽu��^��n;��:��a�7%��Û[��w˯E�9�D�s{}�S�ţk�"�E���{��!�JlU���jV�#��]���Z�d�`m�uk}��ϕ6�s�#��b�.�|����?��03~�_�y��;���>Z'��G[����PW:>��[_���<�e)��Ѿ�b��'���v}G��HJΖ)3���9�>�k��J�}����.��E�f{oVJ/�,���ٌWu�<;��9��vf^�Cp@[^�������]a��4��q`_y�},�˾:H:��54$�^71��YZL��c	�TGt$�� ωꆐ�����S��B��0��o��~6�l��lS[4��$����X�^��,��ay}Bk��XO���C���������z���z�<Cq���\�V�q³�e���6�p��Yu`Lz9���е*-x^�:���>��a�6m;ޡy���buG��K�-r-��Z��2�o����."Vt �;,��t/lrOO��n�f�����+�{g/"q����pP2F�"�8���\-�=.�bOnQV�ÞChN�����ټc%o�����,�d�煵FҸ<�'�.����o`_��6�=�0�,��vvV�\8��l羈���SL`�I����@>ɹu}�\[P��j-k%�\�9�U��%(�x'Z�xlwx�,���j�^���N�OT�>�Y'��{Y��{t@[���?���M� ; [��Ǆ0h��Ӷxn]�3}h�B/
T��׏2�k���V�7���v�*�v��H}i�َ��ܶT�����e��y�k��c�0u�����Q~ûvW~7�hpNFÊ���չw\��
6Usj&,�>8o3߶*=��p�ͳK�ّ+��Am����	�զ]�^�2��LZz�ᔎi�R6�M0eT���h����x�v����9!��_��Aq"-���%����������]��	N��+���6cb�%V�5��P��;�c;
 l �ܠkǽ_�W��1��h��{��#=�1�,-6�~�Y��gUO(m��:��v�'�	���|��9�y�h�
�D��H�dR��^�7�;`��0�C��,%y�1����P��{=Z���o��u���2���a�?�u���`�e9�Y��_7����0��fy8�/҈�x:�{o�z��.��^W�$��и�%�ù?�3��A��̢��@��H�>D�;
�&���ݹ��;��\
��Z�rpCɭ脨�`��@���ABi�����v<��oG�(ț�(�K�2;���Hd�;�	���{����ة��{m���4L	���)��x~��~wN��_?z���z%�����ud���Xx�U/���7P��X��	.j���b�H̔���Y̰�L�;Fx�^������a	�YX3/��C����,�}�����~@���_r����0�Y�\�oVw���7��[�AO���r��Ar
����cҍ7��qN�󛓋�$)�b����f������O��Rm�i��x_y�=��o`�'�{���y�Ͷ��,ؚ�7�`�G���Cv8'��%�kY��:�M�T������l|%ĈxǠ�yօR�9��{=���[�H��=f̀l�Z�[�0X��,2)_�W0�z;S���b��И-�}�C��t��2.s;�H�&3�E�p����c����YF���2S���dT0�G�����C*��.��{���*����]�t$Tk��_@�fʤ�<�X�oH���hrh���k�Z����u����᥷��%	�i�)��S	s�e5����؞?�E�[wma��g4郞���K`��|��K����I|��@� �3����˃.xd�~�2'��0�+Zv�
Ǘ�1���;�q�j4��u]��Ɨ��	� �=z�?�����>;ʢ�_W��}:ig>Qռ�'�@m�'���ͧ@q����~tG=�t�UL�����aX����k ��W=�41c&c7�)S��qD���r�������n�3*�� I�Q~Z�lu�(���OcY��/#9���}C7��x�-�Ա���ۋ>��\��9��9g
��]X��f��0コ-��)�\s����%����Ru�=Pwg)�+�Z�]K�gw7��w'+�hdU.�UK�p��%v����\��o5=�J���c0cȺ��e��Z�x�ߵE�q*b+p�30�j&Y	?�_�|��]�O�"v��<�6���ߦ�ؘ�8�sP3 ��+��vmcF��S�͔x3��@Jd�@����ome�����+�x	���j�·�$�{�^s.ǜ�^n����b1D�;5�Wf�x*���)�>�l4?xy��g�j|�����舫VX��ڝ�z��u\�h�.�P�u��8���;3��I����X�GߍW��!��OT�Ȗӫo-�"h�ؘ=����;^Z�� ����=>c댧7C�=�yg���N%[f��bc.�Wu�5��B]�GEH��VuXֽ|��C��=�*6Y㦽Z���|��,�<�i�T��`�%��Lny���q����k �?�O�����VdIu��ŃQ���r[yN�U��Y�xI��馞|gh��i.�-n�*g�C�x(Ɓ1��k�N�.��	��}y14��,��ŧ��������Ɗ傕��@��f:/p�q�F�*���L�璈�|.�)
��؝��V�gE1������q�Z�>SPA�&-7�?~G�����@6�B�XG��
���>;܇��xyV��bwvy��Ȼ�U�{���Ԛ��Zu�x�⟒&�VK�'��{!�'�'G���@'J0�6U�o1`Yh�&�D������̙n���mӒ#�C��"w��yy�D�ng4rG����b��D>fUż���wh�J���Čc ��ﹺ÷}ٸʫ��u�|��N]s<����c��Pw�w�X�z���ܤÛ˲��FVֿua�a�D�hq>�u=/#�Z~k*�a��'�\�GcG�o\;jf�����:�7��|e�H|����?�i�m~��5����q�Q��Q�b�T;���Azw��f6͔Fn���ru���Q��/� C'ݞa��@Z�9/6��[��q��8�3]NF��ql!�+��|W�h�ߝ%_�')A\���oyX�c�mkzy���PA�b������:�θ �@�������� ��kNyTG��&�Z�A.G�����?��9�����xg��!yM7�>�t��6����o��!�K򺒧�ú�:t.?��.�l��V�Flg�1`Ѐ[��C`/��<��P�^Ȗ���cp�U@��/[�/s�?5����O}�.{�8����_�C�4>}ˮ�l6l��{"��r%���wF˪����[�+����Y�|�����ң���*0ņe@%V�� Q���/��uӪ氌N��n�����"�"e���W6��{�g:�B�"��j��4n%��M����������t�&�*]���-��#Ů��'u�F�'�w�t#{� �{&��ܣ{�g��},�v��[{����HW!}�ZS��nT���;��t��J��d��|c:i@�}�#�zGq�HR*�x%��NS�Ri�a0U24�9ݗw��}�N���Xd�c�!m�(1Td 8_r�)ɋb�U�-���}�3B�ݚ�l�5;Ջ�U��m��1�j����^{��
䆭.LԢ�D.x���O�鰢��.��1�1�녲��}�̒��q!�ΗG���ǜ�2���C�DoWu��x|�>���Y�lY��Ӯ�'��ȳX���[��cD�i:���seY��gK򗝕&K[�����˃a���,�/;H�ׅ3�jI�y %J�ەpf���*�lZ���k����1�&]�Q�0(��C�� ԡw8Ѫ�v5xi�e@���w�X��Z��ʘ��v�1�R�U���|�om(��/[�,{hsi�&�i �+-޳nU�+E	}ט�U�4n�/�6(:���Xk07[��}*-K���x1�.>���)���Y�.�礶���;WI�ْ���ک���K��VVf���b��Y3�]ض)1�M�j���n���]0��>�>���+�Mf�(I�8���*z(�jJ!x2Mǟeˡn��x�3Yq�ֳ�֩�/?<�d�9}od��r�����T����W��W4��s%Ś�B��e<�H�a�{Nm\;��eV�g��`�7�lv��>�yL��(.׋wd�w6��&ӝ�q��c�d,�)e�W�7w��F��O���t�F��Gd�D����xR������$�zϻ�j���Xs9�XєR�!�z�ek��%��B����+��ʭ�K`�W��y�,���X.K���o����u�a^��Y[
��Kw{j5��܆���M3Bз��32�ÓtS64D9�\:6�X(V֔����tO��MuFS���zK88
�ԉ÷I�/x۴�����^�n˩pn�njg6h+�b�zƺ���pֻ�绯2++k�'}��nV�Z�v�����xQY��s'���]X�c��)�VN�{���^��Dk���V��A�6XN��5D�8b�h����9�,"݇�r��5��XB��Gc���"�=�J��c��A�]{�_	�곣3�A����x��N�&oF������2�fG)#������>�.\�A���������%��,eZ�6��<(����8��])��i��������d��۟H3'jV����3����9��6ښ��w;sw0�����/��mͬ��I�I�k��D�$BAH��ݸ�׏8��Ǐ�z;���$J�������\�����5z�n8�<z��Ǐ�z��\��k��b��Ƽ^Aj	Pd<���|m�q�ǎ޼x��ׯC��dC�B� �%S%A�$SR��K�H����>8�<x��׏<z��=��$	���WƯ*�U��צ��[�5�v����湭˘�V*���n���kx׍EI�1��\-͊��9�U~�W+cli����m�M�M[�_O$h�����;V1j�W9Z�ܭ}�slj�9Uzk�m�n�ƥuY3kOk5��N���dϹM�c3[V�C�gd�V�꾪��L�}di3���)k�pr$J΁�	�گ}uW��{��?�Ø���l)�1�/�����w��څ��$�##�*1����!5^�A��ܕ��X�C�P��cTK�
�M���eB����(�?�#��l�zBO^���-N˷ISڮ��3��`�T3Qp/u����(���շl�XW�Z��n��?�K�S��s�n�w��W���Qݴ���]�"��]_��LJ2�
n�ܪf팇Tc�9ųT�aji���,U���rn�h�Az���\K>ܞ��U�}��LA�#�I�U�9��yN'�>ǟOkN>5��	�=�����ؤX+=�B9�L �>�\
��-��~��i͐�G4���k�����"���ʌ�@݌�`�wA��`��M�k��O���U�p�ϨUvO�J�!1���|�����<�-�ܪ]k�}�jڰ��}���}�����V��WJ���3խQuثҢh�`c��%���*Bѓ��>�<�s��g猪�?Kha ���ܷ�F|��Qi��5��\GS����֨�'P~�aßYZ������-��w�A�!��9�x��4�����v���F��m3�5>6Z��(
� �ۍl�Vf�Q��W�����ۺAʫZss�ͱ��('���W����4z<�)oQr����pj�ۙXL��)ձћ���]�V��Ŏ1�]��(s��9
ݥ�;h�y��o7�7���V���k�7-�[A�?r��4:��>�c��w��R��V�a�e!u��o8��Zύ�mfu���PF!�o�Yq�?z����4X��}����y�$e����
ʧ�w�#���A�k�p��["]�hq.L_�Qz�˪iNu����5^��r� ��٭���gv�w{3sZx�v���ƭ|5KO��	��ଋV���r�?�f�Z(%�֌|U/=s>�w9��+w���\���v��eC�[:y���~�L9�h��V��)��r���<��J~�tr�jfz��VEc�^�zPO`N@�4WV�׌u����s[��
ȱ_ð�U��%�%����p3f�\�
�C74��kO�bC{�>.mQ�J���({rbU8�v��j�L�'�ٍr񳭚����s���n�-�a�w=���tQ��G���Cv`yvR�Z��Z��]�y(t�G�<{B}N&�R*9�4�@ͅ+�<[@)h]}C�+������̪�~�`�3�yV:w�xaX2�Ƴ�Na���=���2��|�:}>�8�v@J����l�L�A��o<r2R���(%�H_o:��J�PNWd���|-�A�kuq�-�ai��[�e����ڕ� �����l\������tz���)��ho*33N��F��Ʊ'��!N�Ҏs�7Y7ʽ�ZN��c�Pg>�������&f�?�w}Ӳ̙b�K�j�e�:Y�eˊf�uE����(x�9@Ñ:�|����@;�E�xNC.z�-�f|'����pn�VV�vx&��]�\��@�E���,iq�a)��$�/�_w�Rw��{V3�'�}�7g6ئ\�&GOd�h�S[�qTaV��y}R��"��3�*I�<o�wu��A��Yu.ړB�����k�Ln�}"����'�m�]�.�n�H;S�C����]�;�w��jA.ދ`���d8(Ƙ������u��ޥC��Mcܤ��U�yʡ��1�KB�7�2β��W(S!OA��İ����!0g}�6&�{�v������^L&�f|�wZ�Y�|���c����+��1+�r�1���1�g�j|�����y	�����*�.���z�B�O��ߥ@ ���������g�o��'�_��p��kMvIk�B��u��M[H��騚q"Q��\�9�ϡ���~*� ����i|k����N��49��ƃ��o5ѡ!Ip��f�!ĸ�5.��>�Ax�n�חozz�k��"��88�b�U5�+����Mt�cH�]�ljp��J���k�o(��P%�0�gm�F�j�xs��C;$�=T�ؙ�W˾�U�",� "�|^��HP�L�ʾ�b�Q���q����7��T�Btk���VwP9�Y'~fV��9�V�ه%�33�ߥ��A��1o7����>qu�� sF��B{O��l���4��:d&T�B�ܮ�O��H��rnT��{��u}؀�)3��%aE���C��q��G���~�h���z�&��;�S�U��`U���h]��.v� +�F�����f*U���On�!Ųd_}�Ry`h�3�jh�h��� �Q�����h��y����cTS����)��ָ�`�X�L5�C�m9.ύ�ĵ10���h'7*�q�I�.�|�9\��x��[�:�?dy�����!q�㻥�s�_=��������ɛ���/����P������j�o�?����*KM.��^	ı���h/Tʢ��;t�}�vn��~"�<P��WV����$�������4.��F�Cnz�z�w+ �V���r�?��O�'�/�=#��c �zf.y��lT&D�}��;��t��7q;��E3�3+u�p�ݷ�*B�Y5�
���1�]�?4u|`���W�e�yL,oF��yq5vC����r�l��[��Y�ZDy��@vѣ�'����Q�99�~Yߺ����to�a����׽x�2>x[��������-�"�k䋼�GN �=�ۼ�3_���\|�h>7�(�!�RL뜕�-q�_1N�rg.�s6AM�V�	<P���d��%n.|/1�u��]{'�Y�4��)$�CM4Fa��<��z�*&?v�}��~�����w7(oW�Й�}a��bi?�จ�踸7�g�H��mz��UUM��B\�U�����4��%�gA�7�!���5Վy�/V��ɻ�t+�t�0�Z:5��OR�oK;�꺙�vh��W �רˊ�e�䈩�����'/�.�k�!O,�8E{^�d9�ȴ��1�/4�G��B�� C*	M�񿽹0��"��}�ݜ��fv�L���S����pȧ{-�Xt^D\zeE�&�Ϝ."S]^���ζB�d����A�T��!���N�<�n}�"���|��DKw<�^��=�l�B�Yp��pc*eQ1�{z%�r�K(]"PQ���++�+I�H����+s�i��u�ɉ�Z��b�.4 &�Oc�Q	�O��b��*E7P*�m66F��x�F<���7��*��Шכe��Z���C���.u�;�.f�I��&*��"��\�[��/	MC�,Pv�`������B��)f}.D&��Ce��'����[s"�LZ~X�G3(/��x��+��b��ht/��.���|�s�{��f����	r��4v��*ۑ�}P��8,�^���l��>��F�[��^�\�����̽��\�HR{4��aT,�jae�<�;}*
^�w��¼�9�������O���F�Z��������39Ɖ�j����M3�4��Z)��Bp9�	�:m����N�$'����ԛ���_�f>�"-�' {�8-P��I��� �;�[;
dn���n'�"y�8��X��~R""wD?s�l@n0�V��9)�?�#��i�x-!�-�����v�x�ɲ�*��k��,V�^1)��tk{ ��UxA�i�}���wm��p�88d���Z�HB��
Z�}n/^�b�ّ�{%8��i�!�f�g�.CQ{x�Qkf��Kl���FY|<�	���R�������_�{
�[��ٹ��,�����W��Cg���ذ�@w�ү��J���Z��2=W]"s`��M�rbD*��3����U�a�kW>sͼ��;^P{aa�-�{��L��e']D\��(�ևB�����pd��W(1Fh��eC�[:y�x��a�{��za�}�Q�ƴ��@�6�5G/(���a������ZUy���Mz��W��/��O#<x$�yFugW�"wm*�ݕ���#5�U�`1�!v^m]�����x]Y�'j��
�1jt'D�Dmp�Y{��1�8�6��ҹ:�s�����"� �"t(�1�V�HN�El.��gp��3��)ҹr�hJvXz�/^x\��~�4SL�������t���A.���$���) 	���l�O�P��
E?r��Z�H"���rLO��O0�s��~#�dI-�4�a�����z��t�O6�9l�=�2w=�D�E���Z�q�V7�b���C0�0�zh(���|hWޕ.(C�e"�[�_ ��l�Ls�d��,����=�w?a]x-*�D0پ�̄��#1�y����\cÔ�h2������e�xT:��e����6�f�ܝg<����;5��^Ȉ��cE�\�%�wb�S1��ǳr��=�n�yZ¨Y�Q���fV���.5%<;��ǿ;��&��Ň4K�:��a����w�I�d�'c��­�̦�J��kml���E��7&��B�ݵ`�W�X0���&2�R)P��Ϛ���{*	{hO�4��Zԕ��ZQ��܆=S3�3���ft&}�>��ve�RgC���u+�Nf��|iu���Ӻ!yMV#ū�
i���p�	C�%h�a���A���.2}��F�o���������_;/�^�c-��D�e���
�}^�zb���6�c�����]�[�u��/�D�ӹ�D#[*���b�C��>jvS�4'��2VPOe�Y}/o8�evg;��3�ܡ��!U��Z�3Bp��n��<޳eW��1�Sy�ݙ�Wy�����;-z��,htg/:��  `@��^})�����c#Y�f5h.��v[�3蘶��>d^��40�P�?G�
��Z��X%|>bpW�>���h�JJ���8�/LE��{k����կ��W!
Dך}q�髦.}�,�Y�Tf���QC;{����+��(D����eAE�}�q�>��c��؂��d垇gB������}�w(]x��c�8��	w���'�7�7���L��b�)ބ����҇�<�Z�l�����T1U�`�e+6>B���!O�h���D�UG'N��Ѿ�0���YK_`w(���%��5���]�9�C^��ϩ��x[G����L�(g@! �8���[f��W��nsպ���%�{���F�
��_=3=��}ap�����:T�����wFn�uds��I�0q|�Qu��S/}���_��hw�����ε�/���Ԟ��y�]�
^O�l8,i@���ԝ���zg�i����I��L!������h���ƴ��M��tUD���[U�J���i�M�G0P��9;L��:�=�r�y[���]��'���>����.r��V�ĭ-pe��X��mam��,�͎�S��n����S�c ��g<��[�F�N�{�������;��{��bD����ǌz����/Ƶ~����5^Xy�=��N���I�:���l롌�ON���"�����uG}R~[����ڭ��-v*��y�뺃�����l�df�0�pA�w�w��_��s��<APԪ��X쵛S�"�lf�X&@L���<�9nԉ/A��F�fh��4 �C�n�e�KXU�L�^�y�N��g�ǿL�����A�.���B���9�dt��C�4X��a|A|A�I�T��3Ȩ	������_���}6�5�r8ߞA&��
hP��}��޸�g�w����\ΰ@�Н5ÖE��N�8���	��,9L0��8���8Nr�.UT�`�OV�K�y�����)�C��K����ؘ�sȧzw�ԨU����FM�'���]�o2��[,��:+�q�Ks	���1��p*2=3��ǐ�7��k&�(:w�ܫ�G
�y�Sj���RȒ�tc���ޭ����#K����n&�� i��f��b�ү ��a�N6�Oٽ6���
�Y���T�]���S2޼��o��W'\Nne�q�N޹7Da��:MW��DN-Gba�Ք����&�Q͸,s�6�J��4�<���:Ǭ����_�f��f���W7����c����2ɽ� �y)�߂q�LK$�R�d,J4+����Nr��P
V�y����vR�gYu���i"S�S�$T,t�x.�R)�FSSuη��k�:t���.^�B��r��Ԫ���3�P�M,�e���2��[�rzHޥ@$��3)���"���s[���v�t�#H�u���<�+��B=Ȅ�Bc�l��Ay�]���}ŧ�R�f�eX�ʗ�����C#|�x��	�t
�u�a(�v#������|f�n��B���$d�ކ�F�ѧ��y��^�Q������겈���6��P5��7MM_e��I�:"rm�����Ц�St���d���)�j�v�=f�F��6���z�]<v����0�7W���n��vsd6��o$����.�ݾ�a�[B�Wb�-��:	�8�x�]3��<{X����%��2R������B2�@Aԫ'͑F{`��m �\��5}e��H�W�_9��]Q��9ݵf�m�mݳ�s���T�w�^�w��>k������j��÷6�uF${���c\���k�кT�]�xN%!��'r�#�^a���[ʎ_rH�����xd�lP�98;C�����Uy�g��l�4k�-�ڸ��r�t���^n5%&��4\���2��Y�+V�e{��0<��v��o2
��g�FJ��hv���͹x
q�Ŝ]Ȅ�̽���kѻ]n�o��y|��]��t���a=�7����j���}т�.���Kw�,T�T���g2.����RQ:��wlEq�y�H����+�}/��ZZf�gV�7�O�G�n_*�R��`�*�cu�:�;g4X|���M�t�N�Q|v�[[�i>u�d���m���B���[w:U.���T���Wl�rIa�2�n�Řz�;c[.�N)���m�dÈy;�ٝ��f5�%�Xl�)�b��uRyq0���lsU�����z	�WD;��|�+kD��NU���)�����5�b gS��1��2��ۙ��DVN��qEe.Z��ax]cn�av�S_(k	V����cllܙ��rD['t��E^�rU�q�kt�r�!��~�g9�g��>�۰����EoFA��잏�U��noSM>	���t�sa�Ф�]k��xÙa,h�.�3R9�ru��H%-7��X�^p��%� Zk�-��qj/�v�1m��WL�V�c�^����vE����Io)��_3�BuKb��Ns����3�vv<�ڡ��Z�a�e�N��f�a�gS�S1,�'?�YX��%,<S��}�3+t�"6��s�wc��#��I�V8IZ�l�����n�N�v��J��e���8VH��6���5s\/W] (�T��6�v�R�]�4��1�Q׷�h0��}������k��eVR!J	�[�2)��˥�������[K#����$��o�	��y����#�	&1��6�Ƴ��H��ȹB4o;���ZcT��y9%ho�b��ھ����yC�9,ooF�Kr�P���]��/2���B�e�����3_Gb9�ށ��I'#��B��V��!=�{���b�v.i*�P����jCsP}x7��>��������p����H੮��Ϊ`����-���5�Zw7���v���bI�_���`���V��O��eA �h�u��BJC]��.��S�D��!�-c�1��*Z���3���g��9�GIyI*<�27y^Е0c���Y�q�X���?��iKŶ4p�`ƀ��򥱌B_l�� ����54�i�R�n�5���N���7��7��:�mc���bOr����D�H#�e�J*�W����ͣ�| �=�"ςȒ�jIq
����M���Ǐ<x�<x��ׯT������� T
z�n8�<x��Ǐ�z#"�/"�PB��J�S��q�x��ǯ<x��ݏ�i"��X�\�nk^ŃPd#�M��<x�㷯<z�|�{|i��75]
�h���ݶܭ%����<�76�6�J����nm�\�j�M�b"�Ѷ����Z��U��DJ��"�*)��[���Z��mx��颋x����nZ:H�5 AH	(�r%O�.�q��(���n)HXa4	@x֯g.O����u.���xv��5�ۖ�̂���k4>��+�ҥ���5U0M�5h܃���Զv;�%���
�rB�"7��O�K0��FdfG'��d���.2�8�@�d���N �����$A��(�_�D��"(��TI���1�co{�w��m�����~{��5`�^�cN�$R^��	��]�,����2�c!�*�PX4��©^�F�����61�$�{��/C��es����l������o��s¬d@B�y�ѯE\�g35�����1+1��B�kо#��0��:�������$�KE֚xh���)�5>�<�W��6��]� ��W���kjmA��5T��Dj���RlHh��|4V���곉U��A�Tw7�!��)sJ�\�D�9�g�� ɟeu�T�p',_#��	W�+;�j�����9f�Lc��������K�-̜��B��Ȃ
�+��
���U��a�VF�i|}���ŏ=$��6V�U9����eJSPEǅ^��@|y�����Npf�����_�Նg��Y�׶��Kp��m�ງZ����U�f�����}5���s�F���w�)nƺm\q� )�C�?v\����eM�Q����X�v~�n47�n�s�5�GL,��+�9�V�|����M�~(n���Cn8�!�����ᷔX�.�Z���MB�J���A��Ɠv/���+D6��(�����NrLO�1�c�uәyY�
��_g����>��s�^W�h���r�V��Θ����ط�\�v��oP��Ǌ�`� `UH��fwh`�O��e=�I��L��տ�(~��Jy���n�+��4��ET���'����^�S�kR�m���ob�����w\�h�[�;R2���Ag0�"Ӹv����Kpo\�][��n�q��)-�Rn��y�����-��7y�c�
��=p�P��F�w��qW�����O\�5�>ק��(|9�=_O#B_�0ګ��уd��q�"@��Q��@�߮�~�U~�Z���$���Tm��;{�i�}�כ1��۴�V����C�ze��n�8 ��=�ή\Çf��|I�e�u�O���������O^�?PV���
�8���Ѝ�C�jD�����D����S�=V���s�%Y�Wf)�H��w���-0�����ҿzG.u:9��L'�6:�v8�u�KtP���i&>2	����t�0iF*C��P\nnT�����^e-z�y�r���u�ؑ[��n�[*"8��+\��)��b�j���b��������z_7���	��fa?z�1���N��0���G���M3�\,�'�r���-��ս���k�o��PL�n�$�����=}Mv�u��Y|�#Y�Ϸu����J���e��ήH��=��yml��np-�q�O3�1�WL��ڧ�i���J]#mr�8��\�Ɩ��L�/��f�dk+%���ќ:�n�n��T2��&�վ^Z�7�~�v��$�M,.�۹u9�gzc1~�^��*A��i���zC[���!k��ީl�ƞTc�]��#�^��m�uꂽS�����ǧ�j`�{/A裖�|��5��z��*zz鎟6�5�F"j��K���ʻ����T[�,�Z����t�����w�����ᴅ�
��h=5N�,���yⶺ't����x�t�X�'%r{��Ƥb�^eq�\�����>�$��	k�٣��/F��j�7
�h�D�֓��'
`�<X;{�=X�$�79zFD{yӤ��NV�i������J��h�7&�����R>/�*ZZ�Of���=��1��a�w����:m ��.��h�B�=���W&�jz(f������8]	��+5F��xg�F��o/�P����@!;/]�����S��$�=�����(^�R����	��P�N���6]4yH���p�[ X
Z2/�d��cS�!9��êe�5C�^y/M�̭���:x�#�uꃶ ����y��y;u>�y�Oۣ������[�܎Y�Oy%*�.�9w;W
��?3���"�'���:$e�q��
�����[Ȝ�UqTJ*y��݇ۥ�-��ީiZGo�0���HH�������k5`���IX�\i�z�V�6l�h4w6��oJ(����3�Ņp���n�ǧ@��Q����s%��>�{��͹�9ݛY��5�sv5�C"7��uA��aU�Crʲq��{7�n/oM��4
�]���>�\yfǘ.�\r�З�a��+����^��o�t�]I�}�	*P���Od���<z3o6gLӘ�G��3	��T�"�	�@���J j��K�����w.8��a�`Ckw9�K=˻uZw�&b��Z�xd�E����k�%�7Zܻ]F�5��;}��>> �/c"���v���a��*,v��r�'@fb�硼MP�H���e�Ѵ���3@���Vp�d�3V�]!�nD\f����մ����U�; �䍠ی��p�rM�m���9�+ͣ��<��9�թo6�K7v��ȌG1�����8�u[�����Ҁ�����q��^�t{����m1q��G���y#s3(
���)~�������;}2�2�1%KͣV�a챝��.̾�+3�每�$@=��i`�245�Qj�`ѣr�!�U���YaoV��E���^�}@ϒ�$�ג��2t��>K�?0�i?3vf`��{�=�S��QeH�p����:��q�i�D�ܸ�˭޼���f���P�@�0�*��x�������+2h;�V.K�s�!�T��:x����y��9@0�a(�p�b�v��K�=��Qz.c]T����J��rxߐ��J�.i��r�'4�w�n�Fy�e>�By�08
�=�ҥ�7^�R\���ԣyn�F�"+f�7a��¹9�{V�ƻfÝA	h��ئ���+��W^�1/j��f��>���j�����������g+E�b;2P��z�*sr��c�zu�dy%�!��)����~�jY3<����0���Y�\�4.2+e���'1�Pu���XweU���v�G.��2r����Y]^W�������};���送�e*%�v)�ٜ���=�?n��5�K�3"���/^^T�/>�r��\^����k�k&
�uMћ��>�eC�z�V= u��ȋ]�!n��2#��[9�n��%�[gX�`�������qg��k㇧ڲ��R���lzu�%��\�E�bv;{��|�Bg���8U=��W����(���Y\�n��s:��F�ڌ�A��,�@x��t�߆��Q�;�T&���5_A�D�]з�[�x����nuڐ9��ч�?6�3[M+~��n�%/ET�����D��{�<tTk���{�ЀA5t˽㒧=����^��oT��+N�`%�@�"�I�J��$8��[�Rp`�q*ӎ�t/|���lCl\��}����wX�ߕzs[ۗ�e��.��$�;8�MidM�)��`��7u\��������dr[��S$r%	���1�gO|�3];�	�᜗��W�uk��w�yQ���{$[���]1����}u�����8l�2L�>�_�F�� �ui]xnpRn��M��g��Q7z��J{^��4��4�o���a}��iM�`B�YB�ڃ�g��k�ǋ�T���%T#��ȩ�3V�Y�r`+!e��u��MUI��m�/Z|6s���(d���F�)��p��۟&M*"!����u���&�DN��-��3�ا��*���z�{�[���a��觧ۜ|�`�Cڷ�GL���=���G������7w���5�����a������'��P�m��j}��"���/�y�]��%La�ߡ���u�N�.��iL��j����6�O�v��5\Y�x����u�y�K�5�y,��L���w�,��� ������e����߱�ەԩ��MҧΙS3���9M\r]+_���&+>�kR���rՕN��A��x�x�!��
P�DaB�b�]����dR�;w�L�A�v���Z��.�������}�[�xk�v���b0��.��y����g��cǞw�o&kU��5��[�ML.��˴��1�>Xb阧*�o-ʯ7��AVg�A|�݊��zo����6�5h�4��6�����X@�|<網�Ϸ����������s�Td=�P��~�{�z��U,P�5��ƨ%
��J�`���q3Ō9��a�gkw�q�TS쎆pC���x�ܜ�4��H�<c_G��hb�?֪T�^��[Z�<_,З�[y�0�`��7���&������9���CC�<�;�=�h)uٯu�6���-����»m��V�3Z�����g/6�v7I��u8�r�%���Z���( ���mP��u��qT+�)Q���*��z�IJ��A�G��]\+��b	�=�x��غj0�41،��S��٢�l'�&��蒨�k�p��Xߔ3�;��.��v��{PU�9U���Y�D�
,��V�F򎁽��柧�܁2�{ɭ�eR7K�q��3���Ի-���Cz��'-�uX�Spڌ�ެ��H��ų��R]M���H{%֌�2|��A]��c)���S5$��������d'�ڳ>�\�`�1�1�m�i�"eL�Hx������p�L�{3ۜ�7�%|��;�ǘ���=Ξk��Y��,�f;z�c}vl|6��|~ѮV�}+N���K_vn�z㺍E��+��s�d,���gDoLBމE�l����֯u=�t���v< ]�m�o�w�x�h���Y;��z]�nA���B�#cUwK�*S��8RS졠[g�+�Lf��DE΍F��H`�r��"�wJT��[A�N��8NM{T�ѯ)Z0�4����g�;�n״C ������[p+R��$�ٱ͒[�^C�mj3�vLm�/����N0l��W��K��m,�����B�kFmueC�]�UchF_�����񗭤���h،�s�}a0=���W����Uq�fޖ�QN�j6����m�zu�7π�!w����XR��}�9;Ӓz���J�i֋鏘�s��^.��}hf�g�VK�u]j� ���{v��	�]���/���{ɻ�ku���B��s��.��oT]�K����-dDr0�y��N���ɰ�X�$K���`~���������܋~�l9qE)���Vp=➐�Wr�U��jw�uK"�r܄N��@Ӄv�UE���_��{�7�5�'��Ǫd��t�4+�g�Yl�[��}ɜ�a�~�H����W\_�:a�lM\=��an��n�$�清�ܷo�i��l�����% W���]�g��Uǻ�o�3jY���}xI~2����d.��"�3��u����b/�&9<f���ysz^��I_<zM%�Cmt��]��7]���s�j곝[L{=�w���@s�$�||�Wx��V�5�W���}����a���Q�[8����U�V��	�Q���U�Qy�N;�Ģs5�P���V-AEs��ݜ��7���=�|��u}�Zk�%l &��T�L)[�������n�����C*�	�6�������f��Mz�1�����4ޖ�94����뎒����Z_&�E:h#�K[7a�h�k;XNNnF��gY�-p5�����q_n��`���}�B6*�(f�ػ]���6��v;�RW+�� �{$��l�C���V��=.���ps$c���D1m�*˥yg)�EX�;L�=�Yw\qƳX��]��suMkCy�ip���e:�q��r�n�ҙ�/#F��F'��.(D����.��K�ЭHctfU�E�ܚ9�;�<ʻ���z�.$5�t�(�Q5�{�m圥(�yXǇ�^Z��x�)������w�Æi6��ޒ�8�Km�qPVBFd��u�r�e���"f�UՍ����B�C��Uc�k�f�A���'�O@C(X�-�,��7�4���^&�-Ѐ���Z�ޑ%vf[|����*JE
x������_�^�T��Y$�d�3�X%s5�xh�E�>[����*��Vj7[%+g���L�Ә$6�!BG������Gv+385h�訽�T��q�ώ��f���b��3����U��e[ͽ9N���:�n��+�T�<��ZT�i�9�J���qۧ�ћ�3�,�)������&ٷ�Gm�����h�9�v�0��D�v�wg&�܇��,���3jn�IM�������xj�e�L���+��Gp|5��7sl�Vz�wT}	�]�ԗ���q�tf���h�ݮw�����j�jm��{]v�J�5+B���Y^�2��r�䓂L�L��8;�VJ0�^�慱��k�Va$�����S8]e��.~��ɝ��h����~�Ж�����W{��3?��7�,);��v[�;�##}�V�L=Ů�OtH��v[[٦�3���E�X`�'#��YdV�u���CT#�.�sX�;T�T/&n*	�J/���ځ��&TB�_V�j�	�:�C�zotJP1yݙ��J]����n�L�/Z��Ǵ����Ѷ3�u��W4��*�2I���-ff�ӧ�����$ON5�F�������Z
��� ��&�Je>$�r;��<:6�e`�t��0�n-aZi�R8� iu�D�x��#���K��!�2���s+8�le��IM�
�7*�5�8i�|:ژ�i��k�-[*�橁VSr�7��r�^�B��Z�i���AEx�N8[�y�xn�l*
Z'gWF���%j��ɡ��&`J�M����tr]ܛǨ�/�\��;�a9כ�E��Ɏ��pr���ܜ�S��Y��V����o���ᜥ�u������r�r��9A)�]Y�V.���rs�����g%f��7ݥ־p��[��k����N��:4�\����dP�W\�,�t)vՋ��Pk��΁Z89�N��O��}��j��⹻Z���${O������OX�Au�D���y4���ǯ<x��<z��v�j,�\P�� H��D�-�M=z��<x��ǯ<z��E��t�TV�2*UP�t���8��Ǐ�x��ׯb2"ȭG ����#P�R�m��8��Ǐ�x��ײ' d{Dd@��B@��65t�._o��Q���N�sF�6�mʣkƮ\���׮�lZ��+����r�WKr�ʣ������m�5�j+���������`�k��o(�oX���|�����#Qz��|�!1���R'�N�&�v�A�X76y6E��ugN��zV[WU\���מk�=�M�ӏX�c���y��Øx�d���=�3gg������7�Ƭ� Q+O :��ށJ��f��[�H�ɺ�����o�{A�<{Gф��Cp{�l��b���ol��y�S	T;��n�{�����<�-ӵ�O-���w�0 ���_m`��Lz�t�D��c�hk���^N۷ڞ�n�`�{DhJ�/~�z��5��?�Z�e���*�L��McIzam��QO�~��b�U鋉5Ꞻ������L�F�|��HM'�q�ֿ�a^��R.i��R�y���ʢFq7+E�^��={�r�iK��I>�ʲ�>W�u�7!�Rf����)M>ܷ
��x�֭�gD,��X턫�{�t��
l��u2�zx��a������tSٞD�y�"�{�	*�^KxUC���M��r�6��ylɟf]����^V��2h�{ڎK�ŻG;��o��l�&�;��� {扆h��ʙ�2�Nr�b��dB��so�L�E�}���IJ��<wlD��̙�5Q(��o���=�Ӳ������������ȎDگ���~��$��`u��{<��W'����+7_':�]�u�ɦi�v;�"�l?0�1����A(F��/��rh�:�7�/sj:T�d�>5��qx�;�ߑQ�ᵫ�}i�p�5�aܩ���Vh�s��sw���DgOw�\oz`��/>�֓k�ƙ�c_�-�u0[��L��el=�0���x�(�Y���g��H��VzT��+�Wx�#�M�tg��Rlq��42���B�L�����si�'�k���O�s�<��0�e�����tru��;�CÌy��`��u��p~�����;D��%��Ft*�,+��/9������Ő�κ�]yY2��/����݊�1Q��uĽq������[,|����������WY���!��t?`Nwe]I�<VR�tS��%��Dx��j�_���,7]�d�cOn�^����t�����ܣ�y�.;�3?d���wëz�X/�}�1�>���
�!_m湨�`�˴d�g0�$�`i��z�E��bq�MӢt���.���N[��	U��A���$2jj�*M�1�cכ�o��t�|�;�{�O��t�e2.U�Ա5�(uMo
$S�N���i(�H���Q�>x�f�5�(ˎ��I[��l�kt+�����J���w3Ƚ^\ә�H�C�ކ�g�C�uI�#$����&b�V-�ogA%%*�-�U̎��{,�bu�ww#�J������.jE�#C;<#՘����V ���kI�o� 볲'zYhmwvC���O��@G3��<�����s~�%� :����G��޾7v��N�z�u�� �]��f��H���T��2o5��[�D����'����r;;����ˮjb��HE>��\jhd���_H�ٝ��=i���v:��r����z�d���5�O�*�(�L����^��"gdloWq]Kt�JVN��&Pe�%Q����������*2�������ڷ�3�u�$����޷�z�jcӼ���I�5�oT���+'���vSW|D�cF�
�R"EJ�Ær3n��z7s�p�i��sm�g��0�G���vt�b�.��V�Ė	/^�H���ݚ�|$.f���y��k_JvK����d6-މӻB�k=��������]I���|�v<@^za���7j.��Kw�W�n�M,Չ��ٛ�Ѻ�o��ގ�!�l3���0 ʺ�R��o����Q3�Տf����}�l����<L����y�+�����?}oX�Uy���	���>����j%?��׎]j�b�΍��3]ɒ�y�ǈ�71�p�����_�*Y55Y�j��JP���}���:�s�����ҧ��n��:&��z�T"���2�G�7S�=Ǳ�э��W�]E�t���wg�7�"�8A]�T���r�����q7�Z3�|6���l�չ��wc����8,
�Q*���56�mMF���u�Z�^\g��|�>�a�]�-��.�A�g����,�3/��=K=��++�8�Q����|��5��m�j�D4���c�?kj���m�k���s�y�C�j�fAb&��NΦ��9��C��XKj�1i)�f�M]�Ya�1\(��.)s̖�<�$@N�ʈW0��os�3�y�,%�gt���GO�Ӡo�! ����|���l�~c�1�j]w��vM�e=�վ�\��Y�U�Od{�y�A��a��>0���Mq��g�PP�r�]D�+��Ǟh�4
�w�+ˍ�/���]p���}mXvC��Q	H��:����mwW�Ʋ�9�b�V�?t�T~��oQ�����f�)�i]������a���݈���OR����WF���g����Hu�爉X��*����r������Ʋ�'�7�{A䔆V7����V�Գ=���fwZ���"t
>k�[\��3�-��.]g�����^�Wu����z�~�Ǹ���63#!��W�[X2;��Izםk�4��{=�i��)�|IMr�v$33l�b�@ ��B�8�DMI���b�b��m��ٰ�(A�������R���Oa���j�.��`l���`��8�h�ة����ͷ����Z�fc�Z�W�C9R��ޡ�+�����A���x:���uոj���@��2��˗ƙ]P֕��̄��-�ه39���
�9(� �|o#n�e�E�k�.3���L�We�M��L��@�~�������9�':���_���rוu���׶���w��A~�V�r�j��OD�bb��1��I�\�b�B��Țu�����dg� �KU�P��gךԳ��c�;�;yz�<��E����7k��QrL��!{l���.ܙ�B-��MSa��p��j.lO!=�9��Vm��b��x�}�}n�0��A��w{�g[��<��}��˳ˬ��+��"��L^ӝ�w]=�G�a�~�8;��^�},=�E���tK��v�cV���M\u�u�4��n������,9�0�W����Q�:�j�C�l��AUX��U;��V��v�e��w�0;{���装�qݟA��3��p���t��m�r�]�<�OGgr�Ȏ"#!�P�KJ&ax����O�����`��&칍�<]Qf[��!�¤@�]*C��m�t;��q��H:Eh��HX����=S��~�?=�X�q<��N�]ҙm5��O��I�m��{u�\��J�#W�x�����_"�3�����V� ���	��B��X�U�+'˞�]�����J�¬X�����%��v��M%:$v�e$�{��>>>>>>0�K�O�|3Φ#�oӬ�m�Ttq9G!7瘃��k�����{��7< ,�E�oz�Xs�ϻ��r���c3FƆ��j�<ۍ�T3����r��:�b;��8OX2��-�,���v]I��d��u�A�g����O�1z\�B�9\�'�tlb�O]���k�}�F:�_o`���D�s���;�#%�s�!W���
�%F�i~=��v�7R�;hV��i�6�6��2{�;
��Zx���|y�\�w�ޡa�2l�}�A2֒�+~�;��]a��Z��ZI�~����R�uE)�ߠ���y`c���cfI���^���i�����&���u��+u"�������`V7�E���>������z���7x�{�g3�27�L�J�:n^�uQ��F�8�l��-=D����3�����6���KW����0�p���$+���~%��~/�q�����Y����X;q6��>���Z?:T�7�Ʋ�Dꊮ��8�����ء��	�svNY�}�s�Wfp�L!��M"֣tKr��A�A�kso5������f黷n�b9���M�4Ž�.�:�^����������p���߼�6�Q@��E��g��S����[�/�]��2���3ң��B�$DnH���Q�r8u�f�]�c�5]��l�MKm��p����%�5;v�4�)�}3ܕ�gGOx�w����U��3�u�\�f�6������ڔ#��/Α����R64��X���R������������OPc|��7ɤ?b4�G=��s�U|ԛ{9��m�yߴn����	O�|t��g���h-a]���WM���6�lY~E��6�4�P~���K�������.C@y����-�ξ"Z��Zg�yņn�/e!w\�3���|���kݢq�B��ǃ|ïlfv7+&X��:95�XŮ���н�p4��%�H��Rvaŷ�6�so
Z�������&����f��*��:}�g��LT��1wJ~x�?����
K���qog��l�J�F�\Z�f��V�(�U-��g�������/1]u����[���c�W-�*T�����suqR캙�r�f��쁪�f�TɆ�I=��|�:���KzZ��������G�1�g�0oa��D�u�t�ݿ�>�#���x�-�)���\5D����k��b��ن%�i�����\"h�W:3Av�Ɇ[z�<%@��Î4�v�wn?^fH�>I�9��H걅�7���,�u����]��Ec�Ao�tRރ�q���T�Ff�`E���QToj���"僻
��@�
ky�ճ��ziQ������;<�zh'�lj�nݜ8lH^��!�wg�t
1��Ά�pz+�i�9-_{&L5�D�.l��*�_~�\nF��u��Omz ���2s�N`�����_�;k��6֯/�T��g���t+l��3a��`WLn+0��{_�
ܝ���3����tG<n}�{�\��������޷�FH��X�V�{_�ʾS������W���R��-��E��XE7�7ˈ��!J�kj�9�3q-	�і�R��Fu��횲�J�J��;.�o1�L]���0�ϽFȣ��ٓ%+Ww>���i�F��D��u��O���y.b���Af�9�2��·�_d|>�u�Uy	-��`F1���3}�n�vW�τ1B�p���m�/��h��6�j^�_b�MwP������X���`<T��O�g�s�߮�9�xǴ��~��~̌+c.�2��p^%��d4=�����zI�
�����`V��
#�پ�r�u�H�����S����Xꄙ���.�tE�eB p�Ɍ[��ANg{�f��bY�<{n}�n%�5��t*�4�w)N�<.�&Mv�I�½����$V�U�'�"i��~�c�����h�$��e��M�����V[D3:�h�.�E,�6w�-��_H�IU�e�m���S3*K�a��{�0o���ğY~���� N�-�M�s�X���)y.�>�B�C�<- ��x��T�u��:���r$���^�g��T�̱�����m�-c�x�]x�SfX�����ms�\�{��ө���I���9�#�+��u�J4��m�Q�vS��j�vdz޴�ݎ�ޱ������3i�J
x@�3�aT*�n!уZ�]I�\D�2����Jy
�a'��ےP��M�k�I�Z�u�p�:m�ڊ��'���<�)M>��]�q��2�kj��v3esxpɹ��T;T��`d@C#��댃�Т)�h��v�m�wֵ$4N�,l�y����
օP�5���݉qw�1���s״��X-E���e.u��Uu:�U:��EG�OeH���VJ�69�tn.�6�J���jmŝ��Z��D��(�M�ɡ��w��gKJ�;uw(EVi��Sl��$벯vѤ�0ֶ��|��M r��B�+c�p�
ST�5U��@we�0p�bo)i:��CS�˾���m&�g.��m���NL���K;i�;3�v�(U��'a��:�x�F�՛ ��"�/d���Y{UF���.ύt����e�\Z�"��^��㽛[��-��K�U+2��S�p�����ԕNɬ�.��*vݣ����1��)���̽[�]a��j؃U�K�M�'���^k̴�WW�����N��>�L�]�X����	|8�%;R�f�Y�aP����H{��K�fLZ�a��&��xL������t�����V���H�<C�������UA��4RͶ��#�$��B��^�.�?�m�yzw4�%k^��B!f�÷��;tZ���>\~"nر��v?n��N��&i�=[͗kzĒ�+�j�z���CE㼊
����r�Ws�gn��l��R��1C�z��m�A����\sM��v��c����;L�;�����D�o���&�B;jG׵�*�8��>��rt��
B˕��J��b�w��Ht/�t����\��+���n�k����q�3z��̋�C�!������U��.����4�'�2�f����Z�D\�X������|�N�]��N��e���ش�����P�XOhG��v{XV6�7�������cN�sqm)�"-�=�]ʘ�.�4y����҉͔�����Zj��΁� ���崧o��rY���|8�� F��Gw;.p��j\9c�R|��ӽ/k4�W��\�μ�rf��q�R�r�*s��u2�LR�b���>;z��`+^oA���t��*5(���U�'�Tnj��ٳH��ˏ���tc�4Z�u�Ggru�;�Z������9�J\�F16�;���]��ːE���:T`s�b�1%^*9�H7��̽�x�oe:rb��$A��KPZx�#��%k�a����(�.r��5{\0�',�B�3��Τt1~kl��}v���I'U"b��*:ٍsd���?�C	#�� ?E�2�y�#�U')�%��Ǯ޻v�۷o���׭=;�d�s{V���M��#�k$�BD�CO[z���nݻv����4c���k�u|w�ȥD!�=z���nݻv�뷯_���w�6�Z�͹�ݵͨV���z���ݻv���o^�z�*(S�����]5д�/�b�����\M\����3���������(�����^�ws����\wr�RhI$h��a7+�$�L�Ý˘��9sZ_�ǥ�z�W
<rY���IU!b�З.@ �����
}�lP� j�&QS��0[dDl�dh��*Fb�0��M~A���@�FT�L���,8���;��6����^3n�9�[{4u�	�O�A�;ӻ5�:�Ι�kfb��� �K@��NDT$!�H�!��j�(�\���A%'5�
��Z�C���Q�h���1@H_�&A(�R�2	m����ު�kUF�R�E�ue�^=c�M�e}��J��I/���vѧ��|�.�`@��]\�q�e!M\�R�legL�~&B��(�:�.:��l�P�zz̖��7����f�)=�gp�I>����n��@�?c-�a�X��9څ�ל���u� ��D�+;�� �j*S��^�)n�$�FD�#���\wu��Z����J���eՙ��f`ڲ��q���n;c�V9dϸa�܎B[bJ��c��-~�9�(�Τ���x�x���rߝ�Qfw��z��tI-V9��'��A���ã6���%-�+�b�y(�)G�v.ܩ�x|����Qm�e�@xWC�J�rD�i��\[ڜ�:�/��^SY�#����6Fw<ܜy~�nl�<B�UU���)7W�tދa�f�0���GR�+HD�:
:���R.�@,�j9���+9�7vc�(���Qs&�m\Y�h�����q�T^d��.���e`�e���7+��_ۂ�n����L��#9�b%zj����T�ؽ��_�A����m��"��[�d:K��1t�l@�Aq��f�1��c��E{��ߴ�Aѐ\�Q<'"�ٳd��BXȞHU��s�߲G�1���k�ٜ��Ol�2!{�XځB�.���ۼ7�:I��ʕh�i�wМ˹�޷�'K{5쁆�F�~�k��9��
��a��:�v�}�6�To�+�>ݡ��l��_"a�5��F�9T�u˫� �z�$�	�\��c�$����/0s5���gX� �y���=�f>�H*bY�;Օo�o;�	�H�_��;=C4���	>�b�}���'��K��X���ݨ��ٵ8��i�:�������1Բ85s�����]��fۉ�l2L=\�fn��A���6B�&=��(���_�%����u�cMW`���1BJ�c��'�l��{D�c��}�x�Q���	��W��cN�nս|�������?l1�u*6}�{*�m��<݈�y�p��t\6��V���5Cv�o_uQ��TH��v{}�V��+��w��ڑ��ǽ- ���gxa&\IwR���,�|�Y���ڑ���֡�I�J�)W)�-�t.�Wo ϴ��ݰqe�&�����r���vtI*�3+K*q��^u!�$m
�2��#��;f��'syYk�}��������-������k�CF�Rv�3ş�OH��;^0����v�L#_Jfܴ�dHwg�_�}v����
"kǹm�^���0�p��;4{"�Cb �4* X���:�E\�S��;W��H��d[y��U�<�o�A����,�1�%����j������W��z��V)F�hW3^���w{mp�P�\ӽ޻�uz���HAd{SK�t^ޱ~����d�Y�'M�6dЃ���y��%�	�>�e:�j����[��u�	��� s�]|� RS�i�Vn[����-4�d�{*�y��=�U^$O�?�a#�JK�W��Pi��]�}����_���_����2��Oj����Mo4V�*��\u�Y��Q�i�F4F�b����^?Aa��|^$.���mj3�ǞDѴuG7��u�Z��'f��g&Ť���;���:���̾V�ll-.��t�7:r�/�+�U��F-��fk�o��T}�����H$eQ��Gġ�"w��jC�f����W
֞:�E�k�{(V����3v���c2bvY�D�V�{ٜ�7R���1�c����}�gk27���u#��q���0[սQL��5m�==�6�ܑ|�鿹���F7�����l͆�0+�;-7F�4�4��)Kc�RW�`���C������sq����] o�o�3�7��T�V��C	���ch�=:�J���\�������w���c6.�Mp��m{'x���;o�1�ZA�^?��(�D�'�	����;!�L����߬�^�'�0��J�g3�E<*4"�<���2���D��D%NT_e\�yަίC��Y�y~����L������ޫ���*����h���꺫����ٳ3q2����o�;����������F�cf�5�ě�"l�c�w]�m���K��d*�9^��]r�ßV�n�S�w��z�]�")Y�G4�܊�|�i��W,U�^i�<�u21���zl�zQ;;�����~U��̓����.ka�ǖF=t�u!&ƭ{LS|K��c�CxI׸-9�Sn\��h�M��Ģ�a����e)U9�<�c�z�,kj[y�V���#��9Y�ׇ���c�u�'g���_]f�s35�y�c�Ю�R����4�d��_��������wv�Uǒt����]����j��1ëN\y�g�_���O;�=T�@�$)�M��T=�{7���z:	|�z��7D�w��щ9���O��pi�Ǐh<��)�/�tra+7aB��ٻf�@�UU�F������K c���.f�����-��g(	I�1Ƚ{�r��g�"����HFc�[c�\-�&��6�ҝM�ec��UJ;	�Ȏ>�]7��x�b����Wt��x���O��x�U�k7zZ⢨�F���$�V;���>g_����{Ū*WK�y��-�ZϮ�L�r�ʦWףw�_��~�8�S�˚�2V���I�[S�������"?˓G]��92��y�˅wE���~�|݌ҩ����CB ��GZ�v{E(�ٞw�!�,��ť>�{U���e<8��wD;idK^#�.!������;�)wC_]i�"�gv�<T��r����2��Ou[�î���O8]��$5�ݯ���t�ׄC8�u�Umjfu��W#����Ec��zv\��2r��6v���>>>>>>Z���u���ѕ�����lI��O���1�a}��[>�i��R�y��p�7{��qy��ŕ�𮭞U�P�%���Y�u=,���D_Y���uf9/�w^�
j�jM�!(��bm)�� ���m�4��c���	k�"��5n����\uz����-B�6�6�z7�m�E:�v!^=
�����Fo}6����k֢4g7V���1L����3V� �yA��
�(�fSh��О�̫�������V}��T�(��>�{��ipk+��M��!�$��]��|@�P�E4^k֙)X.x�������f>ܦ�����LH���Rf�r}2)�<'Eb����|셞���qL�i���.��3��%C�@�:��u�Oc����ea���v;n��m�����g��b���XQ�Poq�Ql��x�Tvn&���>�v#��{����/��v���Â�����W��^�����d�T\���h�یؼ3�nSޭr*p׼�)�s�[\�iڽ�����d�Owgw��7��?��m)��b!�"3�y��7�g���X���s��ު�rR�1u�������78�reI��G�"����H�^�J�ӽ����o5�[�cT:����*�n������#}C|�CǷ�X����&�1͕��bM�&��s�Gg����C�v�>���\D� Ҩ�A���xt��m�u|lZ�cݰpIS���EF{k�Y�z�E|}����{�A��ټ2"���U�uϚN�D�����(26�;��6��|y�|0>�y"��J�sR����@z��K©��v�kvjwsby[��2f�gyd2�X�S�Y�K������{��w�>\M�QɌ�qB����=7��ȼ--��3=>��n��y��8=�0���j��U^�$ك�����:i�i� z��r]��dV5��SM��6��o�+���0Cp�t�o:�vmz���hB���[�s���!�g�F�I�Kt�Uz�g,U�Jr\��`�0��v�gJ��fp��s��X�4�,�����Z�6���[G�dͨ5IV��~�������ӝ�wo�����f�#��WQN����u>ܷSٛ��$�tN�.�E���|�?�U�׎Wk��q;ɲ�6�C5b��.�K5�2W9�í|>��v��=�N�h�ʴשq�FXN>?D���u���������zx��ipW<=z�1Rj1�/���aecw�]SF��T3�����-���/_��ug�ԍ�4+�`��o���K�{���~�%Mm[����l��h`WbF�&m���kb��tk8eQ3�]�/ՕǺ���6��=�����FF�S�1���lu�l#�q�u)�+�����ݺNA�2l����-=��q���ϣ�<u�@&�P�D�t����gѴ���N|I��mV�=��@�<*4"��tם�空,�Pn����e֞��0NyNMD�>'>??���Pѡ^���f^�k����hv�33�c������N�w8]҅����D��a�}Q+]��U���}z{�.dpd��_.�����r]bsq��8,Vn�ۗ�Y���.�5q��%j�{���������[DΫ��w�9��	N�I��=�K���Y����`�i<�a�Cӑ���m�c�S�;�0_�,�sϾ��n*�C�Y�,�Ul���M�)��UFe���}T�f���|s^�1@{� ��a��𲳻�u'+��x����g=xfٜ��FP�gQ��[���E�\���4~�������k��qJM�5�=�ۺ�sӮ�r�fUL6�m�R/�觝��,""=Th�U��]tZ�&�ϛH����*Ttd4 �/{r0r��@�cL�
�Y��xT�B�D߹ஊ�܉
��*�l�~��`���=�k�R5���9"���:���4�j�w�Z"�Np�3�v����sAW�ݷ�Ŷ jp�p�>���u(�`]8�R�}zl�HjL����*=�"���_��t��������q�9���M�-�Z���6�d}�Ÿ-)ܺ$Q��wt��-^�j8Bb��p^M.rV��l����2g�Bv�<{��z5lf��a�"g���Y�P�5����+�Ƨ�ҝ�;n��V`�ܬX��H�[Bu�{�m.H�v9"��|T��*�S�>d���[ڹnR�j:���ܗ+�'^�/�p)D��1�c���5����^������;�؃�}��ܗ"L�)�b���wl=Uh��j�h#3IX�z��C K]��]�=��T���YͅFZ���rb��4v��J����X��3����7�
�dޥ͓S6Y�����s]�b�2��'{Du�}��ց1�&sf{+��S�tj�~]����q��5�$w%>$qnj�da��u�u����3�v��&7L[m��WoV���e\L����XEw>��Y�t[��fQu6!<���X��ٙ�pl�N�>�u�Mi
I�hu�g����߫����f�~N�>�$|X��=给6L�酁q+

UǼ|Ł��5���9�M��ٵYm���v�����\�W���]��;b�V��c\�FtS�ѨogT��&�����V�j�� H)�:̬���xgbǯ�E.���R�q�7��KYa���nr�g:@����oI�����ۗE;�D�p6Gn��&;�ɖ��P(��·�FB��b�A١_79��[VXq.�>���;8V;ٶ�h���$�@�H��V��`3�N���"t��V��iDVNܳFE�/�]���ٛ%o=e���:�#.b!R���:�
�W>=`{�;���'N��0Sr�L����[�+5[b��$�R�l����#���Wi���e+C�ٺ=��*z�<
ٷ��{��n�V4gl�G�6vq[��݄���7�#qh��k�"��d��n�!p��
�wK�݅w�zR�R����<��޻V�������w�����b�VnU�E1��|�nV���}gcطi,.Mtf�Owrا/Uk=TՎl�K������ ��j����U<�{�IB�!P5��;^��Mw�avQ<����a-�6J�߸��>{D<�[���ǻ܃���űQ�gs6,Y�]��P	�:*��5��cy�ƦV�7pe�k������0��fj��r[{ia!��.�\��p�ӽ{�G��n.ΖA���]^��i�yF�˳ԛ�Q��v�h�͍�JL�
�+m�fMJ�b��T7Ʒzz�B;r0pq��M�87BĲ/�؄��a��b��"��>Ρd�\U�[̳u�RD��e2�Ē7[�^e�,Q��*��T'H�+�0��\[�IO�P��G�U��y^�ɫ�3�:�P}�UD@ͦ�Μ6l�EW7g>�i�/�:*�K�H_��Ģ��vq��,��_��2L�u�L���Į����&�$i��:tp�GXQ|�0j�nv1��"vr�Y�zs4_-jH�&���F[�,Y}��N�V�^��f��Y�ЖhwZ۪I�б�h�ogcg���^�гFI[wF�1�2$�b̦U3�Y�T�J1ݭZ%:S��^���Aqe��]_I*��q8��z��ި,�Q]�Yx,Dل���_dz�,�ZYDf�r��%V����D�-륵�����)���I�ԅ��a����b�2G�;x����H&��u��H�F竁�UFX#�����k�Ν��I��g[W�wi�%*rsx5�f8f�{�o+��b�5��/zif㜭�2�C��gi@�1�掷����P�m�3ah�bE����n����ˑp��+g��{9a�O,�p�>	�0��J��{J�;������(�f��;W�@�BY<�L�uGp�pU�ޞ.&P��l��t��jmN��Ш׊Zy�+�yyB�a�1�R��;����z	{�ӣ*U^ʝ��1��e�56ej$b<��=�V�[��2!*�'.�:G9&���o�L��B0�P}||q�nݻv�۷��|�7�ѣ�]���L�����ۘ�b��w�76A�o^�z�۷nݻv��ׯdZ��G��Q|c��~9zrM��jP�I�y�o��]�v�۷n޽z��$!�L�)�����2�2�H\�$�����7��|�6ݻv�۷o^�z�I$�A�L�`L�)a��CIR|W2DL�d���̌�]!��^"���$�b�$�4��HQH&ú�3ή��WNH,���>��p�3Q��J�qI�]�@�m{�ć�2D��>�nC J��!x�(�0 �dͤ`�P(G+�����!&A�su�ח��FA$	��I-���/mv�+dEV��TȬ�zaq���HQ�W�evϚ[?a��V���݆�p<\�g�n�T��1�`f��{7�jt��U�++��u��5�Q���=��9O:\�J�@�����[�s܎"�)��}�Io9�*���R��=�Cf?z{0Q�L�ˬ�Z��K�(�vc�G��	��y{���EXO�k��NA!����+wgwz��4���!k��7 �Sֺ6�F(�b�|��Y����Վw��.�?]�~]�v�H�������l���w��T[�5_��	�nr��)��+T
�͖���fǺE�.��ب�=:�J��e��s��ƻ�?8�����,^����D�ܽ\�}Gu-�k�K汳3��_����z��U;g�G����>z�	���S�j�S!3�
��|��3��C>�B�C=u�=�L�=b*0��{���!?���}_��n���A�ҫ7u��Ȓ����K��6-��ײ��6aw�B,9�����ޗ^y��ڔ+��
Q%��Í+2co7��<(�\e����Z�v{�'���0���6ͩ�.xv�<��%�CU9b�<����C�38��@�^8:�O��I��@��)�>����o7�����X8��Y��.-��@���mv��Q��p��K�?n�#L���[X1��H V�>��V�!����P�z�zn���*��و���]h�D�"st�/v�R�'��N���xsXY����fg��m���ƱJ+��U�ܰ�g�j�r ʳ&�U@��v"^�4-�F%��XA�
V��5/z���W�{�7BT
o$\��>R>�v�v�~)�sc�Ft2�Ύ�N�Jy�lB�ᢳ�7})G6����K����"�W��ל�/"��ٞv�7��u���c��!S[̽"��i��)�L�n9'&�Dqn��n�~@�N����"��кatz�mj'ԪP�t�'�s�R;��oU�q�w� Z���
yM��~Oo�k�bd�����Ƭlm��7_�n�z�n���+vU�t�����7�Z%�,&�"��K�X{*�aϗD�R[�2H��fˀ<0�Y��0�@��B�q�x���M_Qu��z���@�rk�º�3W�/>��4��� I�,�I�qF%�����������#��yF�Tf���a讷l$Y�z, ( ����@>>>>]�������������U��LCM�hL��i�j���~�'�e+��X��co�[�7�\�cue�tU��z�b�:ND���K��/y���LS����z�f�#nwSg�܅�g��2��[�~�G+�L̒:jp�{)��*�����M]�G��Y
��b2}��:�qV�d6G���g2k9(�7��;��ok��ϗ>>�@h�F��hDy~��tBZ�����z��\/WV�L�ߪ������^�Q�7��-���BS�r#l�1�]�{��w�g���˝�M����H���yF{U��tןn_��������y��3͌��dFC[����ґ���Q�=vջ/Sv�zw����p���Sm�ix�ܺ1�dR�l#�;=)A��bbita{�[5��sw;M�4��!�
90��w�oX]>���K�c�hwo�M�a�Vb�;��Zj3�:n��Y��Ǫ����j�j��ݦ�K~�+m��b����ޕ�?I��ZW^mi"�f��g�l�bk˕g�2z��+�d��9��G�ݭ2����ϯ������3^���lL�����A�=}M��G0pj#�
o������D�Q.A�435�M�b~��S�Y��[�b��:�C�[��hjw��{��.zr�����:��_ ޥ��O���>D	�u�l[1)�,���#Y������:��Wg����(���~;��k�m�\_6e�溏n��;���E� �� ǵP��Ǒ���]�iD�t���͕�Sm��fhdlT��2�1t�ˏWI�����n*�k͌��y���wPG^��P��=0:CnsP�s8A�f�Z�l�eY8��9���-���n��?OSEǟE��4���Gvo�
�z�=X�;�h.__q����5��hf�l����X�I�dS��3ǟ��>����1�6(�4����O�b5����sy7=/Wr�k�׶yEkdz�"@�����pU��0�����=�!+��F�) �a�g敓M��09�߳�W�&��y�K�>�>�
�I�w>�_,���x���sP��9�p�g*Vur�zm�G�󟗙�;�_�;�st�1�c��M��In����6;;_���`|�
��N�����XӋ��U�mC����^���Sdt��
�X%�ἧ�����a
�J	�c�f��ٹ�l�4"XƼӋ���]HAL��0z�W���!꯶�'*�����*�2|P)J�w-,��w#������B8��R��_�W�s=W�p༼_C^�~���q�q]�Ò�Uڎ�u#H��%�L3�܉�uʸ�g�{���OzR[��F���Tuq�"����;v�\�;��Ω��΅��6)�ȬM��8�y�$��{��U塦nظ�2r7X��~HQc��p�ޟD-����du����Z����S����nx��k��V�-�m��#�,@�3�sk����ɛ���L�%�V}�T� ���= �0͐D�8(�m��`���Ѻ)���7GW�?��d�SPͫ�>]y�u��aY\�-1r��%�8P��mj��֪���ں�<J��X�7�R�����Տ#��\u�u�]��4���Z��23pJ�CE��o�ܕ�R���ɩ������o7��7	�rO�v�[n~�^��=�PuzB��C<�=�f� �z��_lAS ��3Kcի�	��˷�`��Gl��;�}!ކ�,�2�Ml���m�������p�Ʋ�����xv��tq�?`���7z���m#+Za��0e2�x*C�q�_ �u�#4��#c�E^oF��?u�<i�]̥y�N�CX1
1..�E�Ϫ�����Kv!õ�����S=�w9�&jx��	��:����W�����UF�Y엎m�U�9ˌLI��p�@����6M��N����\�kx-��A�ݑ�],=4�Z$��ؾ�X�Ưf7�*��>A^�G�g�F#T����OM��ߙ2�F��p�Ί���<���m��ֺ=á$R�0J��T�F�b6e���ImS����k�1d�o~)-�FZD�^A]�JK�O(Tښ�u���ۡjC
��u,��V!�)�2ތ*\�,�8o�cM���;4p����A����*���ku�R���6�0�&ݵi+8�&��f�Wǣ[����;�!�9_ri7S7XnE���u޾m�L�9F��~���������Zȁ�|=cy@���D'G��(Ι�'.:�QӪ�����������5S��hU�s����aH��[<��f�H�w��������'y�N�Ky�x��]%��6K���]U[�����@j��4i�]�y֨i������kIY��m�)B����;co��x�Z���W�访C��������!LՇ�[��L!��0�N���G�w�v��qq�k���ս �V��:��<3���X\Pq�u@��"�l�}W��_��NWM�z���{.M��2�������y��D�U6�Wt�N�O]��b��!��"9�lq� ꧱�·>Y�ʍģ"�������e_5�J}|vޡ���Ԅr�e{�y�	�hا��g;�
�)e�v*�V;&���W���������|,v��/��I�=d�k��`�M��^G���9׻I��b�[��G�a���-�#m��4�ۦ����7�km�}�r�ʹ�vY�/��mhދ�9+�hzo<�6[)<�f�d0iN�ZS�B⋄�bZ��U�L
�v�O��9�-ё\�oCX�c�1���L�;��tU<��gs�Ә.sT���7�8�4��2�c~n�1sL���;P��']�74�Q�Ŧ��d��z���Q˭�y�h-������x�ؑ%��n/��z��?/t+P)g����I��;z#:�����f�c{���S=�>�lf��8K��0�єz�Y-`��S;um�F%Cw��8�g��3�=���[NC��נq�k&�4�lg���&��úx��1�U�ɒ�g�k�1g�AoYl�9)�˾̉|�<[t0�gf��D"f�ѵɰW�t��`з�d���>��.�.�zӶ�魷���)P�b7=b#��nz���g�Meg���*�tea����ƤZ�X�w���9@u�"#�!C�ww$V�D�M/o�p�����Ѽݻ�}֢�̚��oo1}}��R{0+��	|d޴eJ�{)j���:����`�V�E�k��HJ��2�V�.��޻����I���p����R� 2��r����en�IwflUey[�K�9����j�_Zi]�'���:�W{��f]��!���<���z:�G��9�n)���;;��[}�u��f��x��˵Tqp��na���������~�ߞ앨���̺���@�o�/y����kik3u���2�5U78Dw-�iK�$��e�ìI��~���ѧ���q;;�H0.�2ˢg��ZW��=����B�x좺sDûw������ý=*l$G�j{/��eŢdVp2��w�^�{�+�ݎ�q��ɛ��݆����z��g��rU��@�u[x�g� �ȓ��2N����K���*��yR�2�3��~h��7�����Z�'y�T���t����;-��L�Ld=CЃ+:q�{.�ηdq������OZ�K�k�<Q⊧q��.����A���T�X��i-�9E�xZ}�.���گHޒ�at�����	�'o��k���&�������jʳ������n��w��6r�o��Ie��g���m��Cj�nQ}�*;��wm����ۼ�4l���zQ*ꑍ����=�HeR��v��pJX����KGz0��o�S���Uz�d㓽g8��u��$G.�40>4�q4V�.=�EKO1wZn/7����D���3��r�6O�lWF֨͵�]m���ɍ�i�y<�4���R�JV�i�k[A��u��U�:����B���［{��oMLP���Y���"��]O4f)76��{[�c�R7�,�<{���x�䁴۾�h�r�_uA�#k�G:��Y��f�<s�zWW��N׉��ǣ�L��w.�43�Q��6���8`�z��C�S���9���l0ow�=
��w�Ӌw��2�Tq�>
@�q�D�T�(��E����ѡ�2���(^��܀D�^� ���Ӝ�(��GU�I�.7�4Nz�m�#�aVI�~�����Q�tϽ�L}�������s��������Z�r� �_� �����?քA���4h�P@`yj~R%F
	
@b���e�,c6�����YY�Lb��U��b�m��f�5&V�2�+-�ƥVVZ��kLd�Uf��e�1c*�&�[2b�m1c6�Ʀ�,c6�c&3m�1��Y��-��f[ie�ɖ�c&3mfL�2�Ld�V��V�*���VXɕY�ͪ�2f����[Y��[2��R͵��3m�Z��f�Ͷ���2X�k,fem1��k+5LX��cR�Jͫ3Vjm��Ym�56�ʷX�fj��-f5-��mJ��t�Y��,��S6��3k+5R�[++eel��ͱ����YY�+-���Vkef�Vj��l�f�֌���YY[+5ef�Vj�ͬ����l��*ͶVZ���Y�++eeYYm���AG��|�Q ��[j������Z�e��S@ 1D  1��@ 1T@ 0�Ym����R�U�Vm�E ��k@: ���R���VZ�J�V�YV�Vkj�f�T��j 1D��@ 1P�J�Z�Y[U+6�R�"����b
�R�� 
@`	��V��m+-���ҳm�hU Щ�$ ��Bͭ+*Ҳ�������kZ�)��$
�V��ZVjҲ���ZVmiY[]�nեem,Ym�f�Jʴ���Ͷ���HU?�y��������*����` ���\
����������������[�?���?���^�vq�����>��?-�7���� < ��G���_���U|�X@?���������E�T�`�ڇ�  
��������l�W�$�ޛ��?�NX�?�?�~�D��EUH�I�IV�jY��mi6���)���mi����F��5i�m,�SSkJ��,��eZm6��m�5�ڕiikMSV���Tեjkijj�j�i���ٵ�m5iT�J�ڦ��Me��i����KMZj�� �X"EB"�E�U��J�Ym�l��SV���S[&�Vʦ���eY5��VM�����Y5�e�V�md��V�L�*H!"� ����HV�֮V�����cUQ�����E��m��� �����%�������	�����Z�*�EZ�����[�U������?_������o�EV��h?��k����&��'��,?�?x���ĳ����C�C���������NADW�@@��������-`~�ס_@�S���(?�������r������G����� 
��!�߷�~�����I ��o��?���/|�������P@}�������A U��~���hPH�ҽ9�G�(8��A����ˠ� �9�����W��I�����M px������&|��TE��l
��Uj��G?<����?z�b��L�����r�>� � ���fO� �p��{�%@�JH�$�*U 	D�@E)�)(��TUT��"�����*(A(DR�"�Q%H�JIJ��HP� ��ԩJRR����H��R��	T�A(��H ���AUID(R$�����THUI �TQ[��*�$��(IR
J� R�D�@BT� �T�%)DP��*�(�!D�!H�"H�$) ((��*�JT�  b]m�-�_nw6��W6��J�컸�cv��띻cu��ݬui�.�ն�kfT볶�4M�:d.ۢ�t��ڻ�]�*gE5v�v��i�+.b��TB")H�
(�<  �B�C�С���
�:(P�B��C��= P
-�E5K�f�i�6��K�n�U��;�J�3�ۭ[j�ݻ�vp�Gu2��v�lm��������.��Y��$�*
��Q �� k��Mv���4r�Tr+m���]�ʕ�Φ��j�km�k��F��ؕ��,��whu���jڮ�ET1�)�V�ڰ9WP]���4(��TJ�"*��X�!+� {RX 4�PJ�P�f+t�WC1��T�h�`�@gFt���0 �H��
�"��R� 6q� J� 	�z4��ܔ��4nJ���A��U؉��u7]s�t�����t�J��J������h��ƫ
zk�vt� +vn�h -K ������MEP4c]�vwwk��kB�m�(��E"A+�"�" o �=� 4��Q�  �Y� �� Jk�@`��: �[�:U�t����5L  @����� �*�B���  ���t��e�  �  T�`: �Xh��:�  J6�v�c��C� � ��*�DDB�U
�J�)׀ ;�  f� zt�+ (�G  F]�  2` �Ҙt �a`� ��� S�� �h�"� U*�x  n
P=
�# h Z� �C�V�  ;��@4��`( .�@ `t�FCC�]�]�� / E?!1�J�A� �{FRUF@24Ѧ�S�L�2i�  ���R��   ��b�*��  
D�j�@@��s�̀� �$W &fsQ�בA$�x����fɀbfv�hW��xxxx{�Gs!���"+�  
�ܨ���z�"+��Y N��3�o�9�fjO즍��]n�*M[e�t1�!c&���n��&�?7�ŧijR���Q5���IU�;�0`+��H��#�At���e�-��-.�R�
ōV�⢲�On*8��*9����6��iߔ�һ�q�f�m��!�V�J�.Z�����TՊ,�j��˳W�bR����*�`�r�6:�:�zI�qakd3>,X1��,*l(e1�3ka��&�`��X�U `�S�v�����NFѬy�����wRZ��Q`��fR��"/wI�$��3dĩJ�[���5�����F��] �ĉ5v���;@��1O"&���q,l˕�Z��5��
L3Q�P�ڽ�nP�RՑ�p��7f+��̓�Yp7��1h�n�"5�q8���GP�]f���ՠ���0�toD��1+X0��v5(�M�Tpff�4���ӫ���G(�M77S9�EYCi7
��#��$Ւ�ȥ��DT�����-<
�e�h��Υ@�!��Ҋ*�����dn˙vV���(�o����*��N���"�݈V�*m�\B����P0�E�b��*W���&.�^,Զ�-�;������ %l7 l�.�d�i�Ar��z
�(di�=�ĳlM�-G��V�7�V��ˍ;���J��O������X�h7�@�ւ+�u�V ����"Rw1-�b�7Ckf<�a�ӥ�	HY�J��2�2�ό��K���HKwR���VȰ[��x�uv�>4������̂�i�7n�vԼ��ak%k����ja�M]Ԋ�I�����91�����F�9%9���9���J�cjYt�^Pu�UI��D�u��%
ו
8ݢ%حd!�4>��Q�ޓhI�&a7��R�b
��śV����X��{B��6U���r�
�w�T$��r'1u�bQ>{�*�҂��I-^�uwb>K���,2��;Ah3]%��yR�ߘ�x�6�R<6�۸(��I5�&^6�+�l�KXu&aV��sM�s����Fc2�������v��x�ׂʤ4�ܨ�p�=ӕO[(�(l60Ԭ�����TĬ��j֦� �<��T�D�0rС$�ZmH�P�e�KMD1SۗQ�V���[�1�Ĵ�&-�R�k$��kQ�*V��z�d�5��%�Ѷ���v&�!QF��:��#F��e�4!�M�[qFkm`�˧Qd���`u�	�;��~���*'.�b���V�zm7,EM&���\��kJ�$꿂�i:�'�5�>��J'�Y�A��=<V��уt0)1�����]eeVd�M�G
�^F���V=`U�mGm��p�uy-n;�iZ�Vʙm����q:W���Usk0ۢ��ݻ�2� ��A � Fѣ{��t�R�Ҏ唆=Z7mJ0ݪ;��{t�E\��M���
Kd7��-E�Cp�
�7�w�Y]LJ�X;3bo(8���Utl�IVZ�/VUnQ�ׂ%s���+ ��8�*[��u��R�Y�ʹ&�1�06�)���]d-n��I�̭�m��)BY��;
�By1��v՜�-��E��r,#r`uLեH�;�ܵ����Z�Xbp��R�{��D-Q&��XUۥ���sUI�r��&�2R��SY.b�L%��aE9 �ْ�:q����"h��NJ� uc)aMZ���]c���L�۲*l���hHO� �X�G�������k�Z���f%���(SX ` ����۵'S�!u����D��fmj�2���xZ���8-fYneeX�b��Y{���)�����R��0���XV�>w�6�1p��\%h�5ݼ~�Y�NW\0l��L
f�4��ee�L�Y�C��Jڀ�)W���N��#ǅ�{� �A�mꔂtSҭe��|ѻ�5���I�4Z ��O�µlw�:�p���r����+��u�FؚX����z�gi�փb�4�u�"kkr9�W�IF�U%v��ld�l��VC1h����⧀ӥ6�niJ��n�f����* �����L�R�Z��h-Dq�&b��%	����2�j��F2��3��K*��HC�F��B�ђ��3e�U�	����I��[.�K,D~�7�Z�5H5�.X��X�D:����Њ�6�;���KN/��U4)�^��*�����Ÿ� w�,��tZ�F����\hI������Z i���eG�Dl1&e����Hl���.����% �nfu�g6�v��&d�	�̺{��f(*��J�M��8�����Ti��MҲ��\�t�d:*�"B�����o%� ��.V(Yfg�,9gk3�6`�YaA22�Ĩ��6[��Q���\0*[��9���
j���ѣsd�9[L7����&%[I�;�WNDv-����ʄ;s23%6�iyt���gj(���[m�z��Աuek$���H���D�Ӗ]��?���0�X�eئJ��-<la���.��hay14pe�QJ&l��ե@��jy��&PvY�GC�#*��ƁeC۶��.��m�r��D=oo(Z�2ֱu�a�6�*Mы,4��{j���'�Mn|t�f�SD@@��S�#���V��̄�5i퇅���ZZ��Ñ-X�-���osm����u�[������@ҧ֦֢	S�Q�
h:J���C,�kC��(�Vf5F4��oV�B�G9ڻ�IA��u5
�Z&Qؕ��_n�ZWMmn,��R��ZulF�`�5,���nUb(����EL$�]�5���#K"��9w�!�k31�WA�S��/kZ��C�u�����f��2�1�J`�Ɲ=�%k�Wr� ˰K����î��2�ʑQ�Xg+-H�ŵf`��,kF�^�L5�n�S�l�Z؆܊;F��0�Y��4�"�t
d��pIn��&�4���%d�1:m=�'5�:ɰ
�gZ���
B�gk~o ��W/tZ��m6��6�t���o
��g�B�	��C:T��ԭ]7����v�1����Yf�F+dLK.�]���4��*��ur`�/E����!��{$Y�@�q��ܚE��q+��[�]�%�Y��q�uR��`����O�5w9�yb	wҠ&M��mE4E�.hR^�>E^k�L	[S,�;N�!�fj˽[V���z%�f�佻�.ͲuK#��B^�%Vr� 𚗆Uԫ��� (3t��ܱu��:K� :��JmJ���aPn^�l�m�2W}ST�0���vk7X
̆lc/R4!R�-t�P�)r���(Y6�AV����`�y�S�[�|?+�ځ]�r�weϚ��g	hZP�J�;���-�i+���U�L����f�t�l��Mj�I��2����+�tH�cŘ�l��L1	- ѽ%�Z+�) q�z�G�,a5���B�.�'p`эb�w>rK'5j�]F��m�:t�TW��[�un��B��ab�ހ	z��v�[�/5<[b�+Ħ�3*
�mljj#`�!o(vEc��^L3�ҩdg1�e������R]-̭���B���G��uڴ%4���L�N�`gseKŋ0���V\ǔ�Q6�������Vm*JԦ��մ��l=MV>Xr7b�b�i�.�S2Q�Rt`�bA�X�rf�̖2��J�r�ef`ܥ[�b������4ĕ�w�ZT��K�"�j�(�`K�.Lyl%dZ{d���2��̽v�n��m�^�_�uaE��&�+5�b-X������|ս��h
��r��%Z���P2�lǛF���Ũ�-M:��	���� rj�̭�HA�%��s.$��i�&��-�����l�W��R	^-�1Y��jp6���%�:��1��n�����D�F�ԝ7e�Dּoc���`�j�m�a�b�n��J��;����ԠVS��d��/]�0�f�6�6幚"��u4ڎ���e%k,�XZȚ{�|IKp���a����V�gh�XnV}en�kt(��Ы,�L#^@������2i)��jts�Ǆ��
����f�t-��RGF��=B�ݥRl���9E'.�� ��2��Gf�T!B�� ѥ�ͩo	��#�;\>��I*�1��4�N�u%GX����m���,�q��sF
ݻS�MfIS ��Ս,lJ���h���@:юG+r^;n�`��W{V��yPc���!H�ʼ%�5	c�0��xnQ��W-8�c�ӗ�.�0]�wi���m�v5$�i�@����]��Z���\&�M��ů5���v*�����R&ig,H��8�����ۧ��j{y[�Rt�*z�����,l���� ~�Z�*L�b��ҡ�nP'�{���?�yI
@!��j���y����K&��#�Y��y�xo��ҝ͛c5a@eM�@r��<�����9�Mx�{W[DކՓ��:s p��YG=���������,q4�����6���.�b!�B��9E��*��hn��GLES0�k�f� e���Mcf�'�J� �.�:l��h��B�T�:1��S��a��F�c+e5�4���j�8�w�;�'v�d�	�[��4�/̸vK(\���3o]\D9*e�+.m���D�W�#tS��ѤV6��MT��n��|mPQ!^b��x�	�I�uG.Sy��n�apS��3qAPe!�1����恤+�d���
�Í�@;��TL���5h}p�w�U���rP�N��R[Xҥ��[d����d���g.�ҙ�-,X+#�1bh��*�<��d�����b/j�m"D3[-E1!�vl[��o4Д�4�NXe�����f�ڳ�3K��%Xݺ�v]��U�U��e	N��ŠD5mKZ�f��W��mY�-�m��j}0�n��j���F���Z4�E����-d'(��ڕ���b���,][�N�R��a����7�C�+~�������P{�ee�u`́A���H��J��ڔM�N,�/rȨ�,�Z�4+��d�� H�n�5�"�Ed 57{���Ҷ��8��H��C�:VGk��� ��t�Zẛ%�Q���kf"�'35�Y��:�XŪ�
�ט�6ü�e�1�&�P��A5D@%R���ƭvvf[A+kV+�%f�8H�Jm�t�b������!)@�<Bm^V�Fn��Qh:�ֳ�tt�Z5�\X�h杸b�ŏ�z*-�N�gh�j��4=ߝ���!˴u���iN�nh�O3^5e1�n7`�U-[V�`�K1�?aс,�hԮ���@T������9S�r��8�����FQ�z^d�j�i0E���WM�2�]��qXV*��3Me���P�"��6���_��4lK���轗���I��zc��ȝ<�n��Dbv�õ/��}���3u�Eh"�e�����7Q[�Qk�Ht�Ƕ������Wa���H���jS�bR�[�R dɒI����ђ;C(���x�� f��S�`�&Fa1`O֐�K(ZoZ��.X
�)ە4^ҕ�v�En++]�1Z�����{�%� � 6��3U��u�WE8e�^�Y4�V'[[�)�2�˶��;E�S�%�Y�����m���i��Z�
UV�e���Mm5��L��n��n��Zհ�=F&h�V��\�%��p�"�*��"�i�Ż�!�.��C�&�"��k��&����y�,�V���%�㄄�] �&�b4Z6�e���WL�vX�SU&H�Wj�&��kȝ���w�6F���*�0��,��m�[V~(e�fe�$�ؙ��l)1(Fb����FD�A,���nR�&���V�@��cf�d.�B�,e���^��fdt�cwtcрc�%�7(���	-F�n�:�Y�{s$�`��%�*�}�b��{��Yl)�Yx\�n��p��,�Dy�L#�u�7�l���iR�[q:3w͙)a$>V�4%�u�e^�jƹ�e�(��LX�Z_a��T��*�I���JJP�%Ŕ��3A��$J�V���Z s<I��=�TT�Ђ��Y>���H�%	i��6"UY ݑ³f��y@[� �Z����k�K�����i�c?a�[�M,�b��xzj<�����zӽ�����uw@�V��vR�+~��u��ڙ��&6��1w�p�2Sq�O�X�f�!e��]������S�]<���AqY��L�ԇ/.'�F�)SQ[F3�I�9t���۶V@�G����K��T+)�V�4-Ǚ��]�)�ӳBQr*�������<�f!�N��X�0K�@ѭt&R�0�YYW�C.cӊ���X
A��ⷛ�սn���R�-�oO]�6qe�����,��X�qn��b�
%�.�G�nFO(f+jfkZ*R/%&����Q��5�U�Z���U7sm)�ܔ&[�M;j��i�J�i)�9,�+H��j=ո%�/�����2�\��,�[%"�@����̤���P��4VIWp�r�d"WP�ˍ��ٖ��h�H�*S�F��ԎRnk����5M�a=�v��;��p�ӹ/*��n�S�aaAO��8�%��%[*F]��5��t:�L
��S�6�?�M���l��
�4^8�
H(�8���ł�Jz6� nZV�ZB�,֩�.�c��V؃�s^�����lI���zD�T+*��(�j阀��P_=5�Li�+n�H����:�Z�IF����v6LI�R��	|G-�iI_i��/��eNR��+]+�ͱs.�(����p��:�^X}�Q����#��]��oj��V�	]�7I<:s(�F$-W�3�P�_'�;�B'�Y�)s���[bSU�Z��kwl�S5��a�;*Y��X}��xK����coH�}"��PE��>����BP+�˛���Sn����h�!�Kp\��	�2�ca�Y���p�0�^NN�!чYM�h�}H[|��5{�3�(Tk�-�C�!Z�4dE;r�L(᪹/�;S]暒i��Ќvv���p����5Ζ+R�r���(e���`9�]�f]u��+���37�m�i���h�2R�A<�u��pDa��-"����7*���wY�QDj�R"!��ή!�D\5�NV��͘�Pv�����g+r���E���_0�p�r����ۭ�ܮ�aA�N�9�kWfP�F�}$U�9{�4�8���y���v�%!�i�sآa_X�+����i��\x�gcr=9ǝ(k�o��G$��U,ƳhE33*�(22�#��Y}mS�XZ(����-��Uu
�u���Mc6F�����gl�	�������)Br	�x�נ������9>�y��/�孶�ɣ���,��Q��gE�Yγ�:KbHZ��s���/�dy$�o2gX�J3�+��Cm�CH�|��\��v���F�wm��Â:��Vg'�7n�%z�Y"��dIN��Z�ܺіm��sg)�Q&r����J��,���N�'8�Y�f_�����bc��#�@�G{:+�����]�#ɕ��:��pB�ֺ�U����roV�e;���8ZA�qI�(����(B^t�̋{]Z!وE���h�Wuؽ��b���H�u٢��K��b��}�����D�m*�D웩����U��j���{4�C���rQ��(�jP�Vͮ���:U�-흀�4�gb8�u}�d�R�m+�_.A��M��:�,��}s{�l_�������ëDC�Z�H]0�wմtI��]��F\;��ޭ$�e����lUWK*<��̂���(P�39SI��^uC��$Rx�+im�&R��ݭ�p�}|��F.����\&_��^V��*���/�H��K�cp�����
d���C�|���=�S��p��|b�OG_8����2`W��ޠf���V-5:\V��S���f��9��ɤ�˗`��uI�����m�/�b�R:��{�>�����H�3�˹�2fh�_�R���-C�ScHqZ�:������t)�e_m�"����Q� ��wgT��
�N�^��S��Lv��ܮ�9՚�
��UJFyC �7������I!�1e[TAҭ���	��,P�n�x����д1} �-��#EI`uen�&���f��=3��g2�50��2������d:�e��b-�ݔ�ՙj1j���*�u�_Q:��	�}��!{Yӭ��N�]��sD�EI����`��"ڴ#HNY��[DkW/5U��;h��".�N�Q�+~��Yy��5}j"�y&��C[&՝�c���$&��;�R�O"U4����k:�������#iv��W���w�_PnT�s��[�u�S&�45.�t���X����;9-�^�Gw�@���-��Z��=3���LIw�M�芻;P��\:�r]R�%����
��@�
7�lMʾ�e;�5Jn��Luڸv��ȓ�*WV�><z��ûrEƆd/ԣ�S��:hAc�����BV�r�6b�Hέ��@"�k[}V�����ԡ�9]0j%���İD��C���޲ĵm���M������i���|��+���aU:Dﬔ`z������ܽxF#,�5;�:�#9<i�H]���Z���Ctѳd��ajVS�]��N�U�������i��ۄ����U�a���.���5%xY�鍍�S�̚4uwfK �u1u%b����R�lN�L9e�$�&�r�=��Ƿpx��E�JҺ�4-�;!�S�oq�|4�5�a�.ا�s�.\�wsڕ����Pt�y��鸏^��EuXi4��K&�AX�8	񮳬}�p��'f�.��Y�)i��"�tj&����93��/TvF��V���HJ'�VW�k���w����v^��)}#��y��'����4U��Wj���.�ss��Q���n#�+)+�)�x�Q�r��7G����_o-������ҷ���K��"��)p�յϡ^AK>*�E�^���X��O�=]���Jq�����P��j�q���G�7F���٩uԺ(yDk@=���ET͇xQ�6�f��4X���qN�����F*�]�p=u5���Ԧ�V���V:�	nO=;~�Y��|�:�j�f�XJ�a��9 �aY�n�ǯWUe���k^�ԕp[��F��7����[�8����᫑;�D{F=Ͷ��̏��5�^@�����x�>�r��Y0d����lRP�N���7�IX�:�XyѩN�Z9���^^��=���,����9�tk\ɴ�|(˼�����I�)�Ҿ�w�<�#�����ӯ%.�m`C�̭6s%�[������k_1;t3������]�{��ǂ٘�^�7��騊���J>�jū�.�/6��,|��dL�b�Ĝ�`�$�sTwQD���YG%�����em����ե41�%���K���]:f�ޑ%�X�Qn�Y�؀�;�-��e��l�yQN�
69Q��A�>��u�5���d�"�l�Vu�8�����[�&��j.�3�T�z���B>wՂ���ql���=�q�M����2�N�}�J>��
It��#A�>�u�ƈ����9Po)��So)8��M�1}�wu��Hi/+[���B�-���{9_5v+��L�_S��jlrFj��]w�=�cmhs�����*�Q���qT �ˈ�엔����Q��n+��:���aX�)Y-]e�w]���2�s�ٮ5)� �}mu����Q�i�*�ޫ\r�Q��Xg��:q�avln���t]}[��3(�ˋ.��ďB	N������3sS|�;RεK����@puf
YAM-ը�v��<:�j���w"�Ȭ�˶� ]w.r���!6qf���ݖv	:R�<�Z�D=��y����H������yVQ�D�-i߂H��6}2�3�hid���zi'ʯ����FC�v�(�йT�mK2�E]�PV�ou��@���Il�m�1t�P
k��d� ������; �Ym��J�L�6�Is��
��-��M#4���Upd���;a�N`k�Y\w�Q��k��wf1��%n��QyY6\j�J-ZIt�7Y�⊅͔�ւ)���4^L��g.���j�Y���ss�kI&��8�1�q��"����w/z��c:�	�G��al'7���6���Yuƶ,᷍ 3t+E���K�`��[t
«Y�6��:.g�{���0[\��i�4[w�.��l���u�7�.*���:��m&�@�jŊT-N�3�CT�n�r��@VIC�:��u��zk	���/JO��a�i��%�v0wZ�J�E�o�WF�ŧ�Q`�<��\8!B�X|+�}�;H�yib�.M�Fi���&p�|q	s��ؑђd��:;������o�Ы�E��G���*ŝG������@��am���9V�;X梅�ahN��$V�#3&�ݩ.�,�I���^ROu���jb
�Õ�9��+��F�v	�unM�r����*ZZ�?�]�K;뺔;O6��>����`���8��uvZ1�Mu�{J��X�ws�ʾ���Z0=�Z�v-���-�Q�</�/WX٠�Y���s�1��t�����^�A���JAC6d2�4��vun�WL[b��osc:�崩d��y�{��2� �NL�����h�]�"e}���PR�� ���8lWFNAt��SC�[د�fG+��*̘f0`�oR�R-9��k��`-�*]�O2U�}]t�E/S�B�#�^K��8�V�}�~���ީM�p$�f�\ZέS��:�ྋd���9�+3c۟
��u%�����\��)
q�`��3��v���2핌���vw9&R��r�oN�b�����H޿e��vu3-��
�ػ��o'�dXMm=l��^mΰ��ev�E9Z� {�7f�����9���ȇ�һ�{8��[aNz��X��ٓG`�;��q������O:m;O&�˽���k�)J����z�r�V�A��t��kbwC���*�����3dC���aBo=�c���螝��:�^�"�,���7Z�Fd箃��R�q<����oj-f���ZfX9����]#�Չ�;Gt����{W5]�b�jIS�QH+��b�Z=.�Ü�F[�ti��[��x�8���͛��
��Zy0�}��N��v�	:���n��V����S}�u9r\�
$�O=Y�SE��.��4E>0݇�w>����oRx�ڙ,���:��_f&�Ҽu���{�7:��ZV{�]"��JRs�D���Q�f[{C�7N8{�2�vB�'��w���J�ofs+��8m�^�]m��+8L[�w2wb<Z�ܻT�Y�@�s��th8�U�[ͼڈ�H2��果�|�[�d�,��Y�Wp��`�r���$t�=�ƙ�5���V��X ��{N�\Q(��w�/�
۫\,�זd�ZfgN|�Ұ9���vjdh��qZ���e�n�tE�I�X���f�����)=�����������l�T�4�0P�Ùܶd޶���vTtx=ֱI�9j���ُ�ݬ�-_�X9��N�|�Ba����ӏq��(�Q*�������
Z�qz���J��M��	���[֯�ur�0�eھ�l���gv�mFJ����n-�;�맫�fr邅K������6>{��uQ�����)c�d�c�W7rb��.�ߏXUtl��
6��Ģ���Tm�|��f�$�-e�c�LY����i�dT�6Ƕ�vK@�AG���1=4�0@�ra�۽���o� �yb��cFe�ˮ��Zu��wp���U�ǵkb�*�r�4������e)�nl�d�����\6����mZ�Hj�Ҿ��wKL�:�����D��L�e�^6u�ܺ�V�>�݅5L��r10��]���؅�NB�I�5^���2u��W�9��f^��s��I�Z�""�[:{ҍ�+V7�۽T�Eg&ȻM�\��no,�ǜR̒��8�a=ҵfNxtd�_MŬJt��QZ˳]gXᣫzsR�}�1��#5d��p���Vy�0�=�y�p���^R\����5���V��nV=�r�fdS#�*�U�ǻ9�(��Of�Z������Jo�A�*����0*[�*��F�ք�+h��k&�|�]
��S����D�\7u$,�P_�.�^�4:K2c��&\'�|y�Fe6��6��o��q����sh 8|
�ԫ��B7{NN�ɺ@��s�mf
����H<n�G$���մo�삍ջ�\�ki���e=!ͽ�U�����N�X��'B��f��6�܊6[��� ��"���ȡ�v�.�}�;�ذ���75'�T����Z���ѵ�wX�a�Jp��Ϛ�+kǙ*������P\
�Fgf�l|9a8�u���]����1Fє��x��cS}�_5p0� ��H�o�uP������e���T\+n�nE��K�nvn�+p�W��;;3g�khN�-��7�s��=����<i���]ºKt�|�+.�p�y�dd�c�����!	�y�o;���QWr�4��:7Щ&�f����Z+�����qb�/�ĭ�!�x�g�+�P@W����JO��ĭ�]�O��4:�;޷���W9QM�o�������4����w	鮡�aG��mU�3~��3Ro�M�����E:�[�Y�K�I���I^�z[�z�
���/�]G�j��W�T#S���P��VT�
H����l�BU�3����;u��A���^0�nm$�w��)�Vb��+fr9,�Jocx:Yc [��QU2���U��>��RyL5\�r9�A�Ԅ�W��W��5:�[􎷬�aʙV�a[��uq\�*Ց�s3Qܬ|�؅�@�\��㐬�8zm�E��o^��x�
�������+"hB��� EM�7%���B�����Ǩ�9Q:�������Q��H�b)Z���a˵4Y�M��J�鵺�p�;2�7m5�6���q��o#r����U91��¾��n,D_�Ӂ�K8���W<5�,�������[f��P�I��5
	�j�֟5Sk0�w�]J�FS�Ԧ�*���pM�B�n*gx��Z�o8;J�ϱ�ۛ�t$\y�/�mYp|���m�����)� �ٝ�C�s2V�1�n�cţ@�'L+��4�S�#\�^Y�Z��R��'m�d 
C;{��!CP�v�%�.y�o����F�Uv����v����!�
u��d�2������<{����sgf������<=��4�K.c�.!�����t步��U���&nț�0��5u�iJ�1��ҽ���f�pZE�ԁ����}��-�	�"�0�>�l�P�Y�X�\���g0j��]�E�f�%��E.���8RM�r.Y�4���H`�����o�>apt:�[�j�2yK�*$wN�,aܝ��h���!s��B�F�ؙ����%��giJ�ǽZ�!���k�&Hh+5�펧�7q�:����#�c���15�WWn����n��=K|g�?wE]1P��9hNy0J�v�2}�8#�r>������{ʆ#��8��H���սeR�5G����  ����^��f�Z����u��ݏZ��f�!m��g׺2��#&�:}�#��$��CG=	�l	�䗌Xd�neumWb�`�b����L�wB]�`��.��4:#�\c�h3|].��R��	���l`e��*e�K���Y�n�!̆�D�Wq����nB�*d�9�l��S���dF�L�W�&��vΫT�i�B��/}O��֯s�+�*��X]�R��R�t����ܥ��X>+�RS|&���v�EA�r���WQ�+�Nb=���t�<^��|�B�B�hN��b��3 Eӗ��9��ɮeR!���c����Ӷ_.Z���6�4�v_;X�r��t���]v?���k����	����\{�}�^vǨJ�k~{|-IpE��6T�u���,aOF6�9@`��e�c�0�!m�[�ٻH�WݦYDaՃA�_+V{�K��W\C��>��JW:J�(���x��{՗f�ɪ�ef,u�[Ż�ݨp���JҰS�z��E�.h�h��ݦ�N� �4��b�35�ZE��X��uX��%�Ot��H���;���yuik�I�`r[�4��n��
�y�(t���D#����W�?��N�KN��wsʻ�w�W��S%�E�����`��tKɻ�̔����F��v��<'�v[�>9{Z9C�}t���TU��8�L�6��zF������9un�I�4�X�ie8�u�]#�ʓ���(w�F�h�SS{��wRiG��T�U�k�l;����1�nJ��g&=YX�9
V��Yz�	nE:>�0�S��E�Y��ȭg �pJC�vJ��F���Ү���z�W�G�ݥEB�Ԫj-JZ�]8�x�Ӧ�Y���e�����g��I�G0�����N� �OxY��ɼ^I���=wm�)\��Buc7�ұ�W`E���0�7��<�4�0�ٽ�C@���s��Q=
�:<;m�%�4�ut2��kS�Z��&np&u�m�:�r�#]���؆ �(n��t�P��u[�o��sGeb/�K�{ѽ�e>���y���r���XR�#� ��Z�q��BjlJ�v�I�9@�بd�YG^�t���r���
���Gw<�v[诅�����$�\�&G��#W><�F�N���v̚-=͵y5n�W;mVT�Gt:�'u��'d5Q�6е���� 3�oN֒9nS��p���e3�9J��B��o}�+{AV�O��)��`�].����L|����ٖ�KF�i,#w����[�E�@�5����|:
0Eg��8�`�(�����{��K[q��&���aX_�L}6eӣ;PPR�8�L��w`T��uըd��tK�����.�4��f�T��ֺ�R��nY��M�M�� �QC��a��}��X��������w�gn.��:�pfH��� w�E���˘�]j�Uǳ��*��8�w���z��]�'")h�;8E�^f�5Xz��d�ӄ�i�o��ϗiY�L2rV�Ԧ�8��"�.�}F��J�9�63���e��Q֎�T�5V��Xئ���[�W��`�[*�cS;��=U��W*[y}v�ʙW�8�j�2g��'Wu>��J��*�{���m\��jX/@�d7��`����,`:t/F���ms�=���*u�	�w��kRp��Z�Y(�㴞�r(���%(�`�����0q�M!� �gY�R��QwYY�%�b�mVeG�� kT-tL��n�U��-���ѣ(.Cu4�.u_]K���R�{rs��K�����5(�wV:�j�ʔs�N�f��{�c�5�
r
M�n:�g*mM�ع5,"�ڕs ��4x3܂U+#\n�N��tPĝk2����,��mSi~�w/��\����$��*b��P&th}"�p��d�Iˣ�̫�Ǳ�"*�q�ir��&��`޻�ӫ��1!�X�c�*�(�za�Ug��
ķ��
$��L}�e�phu�%WJ�����!���Y��9���t�#B�ahRV��|)��k�c����f�u��KNu�]�V�謬�L���j���Nպ�i-�t��	D!7o*;4���a?!I�8�GX�<Eԁֽ� �T��t��X�D��F���-y�;L�v���gT��^���L�]=8^[�\+�(R�Rk�N���b���V��Y�9Y8��5+�h�. ���ۥyۧ@]\n�0������EV�%z��M�R=&�8;ZA"�_	ɻ6����*\���d���Z㎢���-h���Ź�*���	��ei	[���Q��j;��L��p9��bl�T���p��v��#a[�����5����c��ٷ|�g�[V���{�#o�e·
���'�d�l�9�,b�H�WlR��b�m�HL��9�B=��`�V�)�J����&�G&-�B�;�#�׳r-��Mҏv�u�Mp����Ѐ@�Wq)P�ﶕ�e��Rt�n�_�$4fU�ɦ`<�N� ��|�]F���:�f_�׻��)����u&λ�UW�{%�@���Fɺ7\���sw*V���[[F���bFd�ұPm N�i�x���2X�2+Tr��:o35���?Y2V��������-t2a�n]u[�m��>E����A�T=qڙX%��@�L��bF�ovH�.�����p�*�L6{ot
�]V�^�C��TP��R�8	]!ٔ!W�X��;�Վx��烉ٌ��yHV��|�q�&s�8�L�B-����+V;b�[� ���f��mk	�ܫ��*,�"!Q��F��e��e���wI�	gg8���r��Cu��V�K�A��X�w��Y������T����̦�i��c��쾻-ڱ*¤yQ���F�剦N�q�9���6����\Ե��(��q����{v�躵#�KT�LSg*]Q.S�.ܷ+n��L$hhη�;�ԝ*�+W���ʜ�.[�g&J3�o�
��wpƬ)62<��i�зݼHz7������yK]n\0.�jī�/o6b���lq��q���PΧWb��<�e'Z�X�\�U�"(X�Z0b�B��\��nRXGD�m]�OXu��78qs6qͧ[��-��m>E����\�c�pS!c��HX�{��M�K��<��S��2�V{B��N�$��9�����Ah���=�M�M*�dc�@�"�lnF��VlR����Xr���'@���E#s��:���h�N�n�,:n�Uy{�F��i��՗����O�"\���mU�N;��N�uТ�Q���x����=Yc���|hG�u�ky�Ad ��Cu��*6�i� �R�<mogV[,.�l����L�ѴsN�F�,���m��N;vI�T	��ʹ8��o��;���,��O�S\����WC^�NK��qp�\�����������ܙ��5� ��k,��c:�rIn�-�?:�"���u՛&������/�\���%3BI�X�4m�\���}����n���9���+H{�`��wאۜx����f�ohL�U�����j�.�n���O��]��M4҇F84�mX�h���_j�v��!�����o:V���vr�Qc�[g"	C��YC.�;���u�<0���KMO�U��R
�a.o����}�������`Q���n������S���3�idu
��Vr�d�F�[O:,����mb��U:��gWI*7�cq�*�}��:�BJS��!�X�ra�{�JEV��9� ߨS�鶌�&������פ�r9��[ZAW�)�����"�s[�`=
�[�9P����j{�@V\�I:^Ɠ�[vxt���A�o,�ƚ�T0is��,��2�*�pX5��p]%bh��u����Rd">*H$�g�^t,�g�zm2��AF���6�a�CTմ%�\�+�qҁ��u�G!z�e����呀1]%���%e�ǽu/"԰CAU���9cc[��U�%-V5���ͩ)p��H�`�����oZd+��p���e����Z}�{�6���զ���Iw<����Ws1�u�U�f�� P�mpWb�wƏ`��r���ʾF��ϐ���˨r���7���o���١Z2���cY�;"�hŁ�����e�,�D]�AmPM������l�b�mZ�0r�<5�p���˲jvwi�EYK/1����2ے�kBrճr�N+]� ��S���ݽ����D��-���1�s/]���v@¡+8k]���m�����m�e����2�
T�|'u;y4Z�y���-r�m:;������>8&Κ+{�ږ��fвd��V��3�r�o(8l�:�������x�_P���6���}�,gU��wjyw��3v��P�x��>3N*��D�ƚ�Z�4����"�m�KD�p�E]�|����W{w)q�����)]0�T��u�#������`���1�Xv��˙��V�$8%���[���3��R��Wr�\@�pQۏq�G *�uw7��]s.Ryz�l񩘮�93��ї:΅A�o:��O60�=kev�Ny�V'�]wQ��τW�{��3(ЧΛO*m�Z���B�Փq#C��H{ aJJ껙�<(�h�v�zAܘ���W�Ch��k.Nق��=&�߭�����;���}���\���S-�����k�vw;��,_���d�vx0^cn��6ag:�Ix�k�5�p�p��7���uI�,cf S��q��f,�w��ӫ����7�N.�<��V1��=��M��;�V�A�q�dqT�N��<ِ��`�N�ӏk�� 2��HݑR�R�[���BS�Y�8�э�������{uz;��t4��s�v��˫�!�u�	��s��ow<��L�f�(�fMQ�j0V�	�Z;�1���+xAi�  gH�%$�	�����.��{@r���-P�[L:�U�wh0M�R۫�D$J�7*�h��O������������^�=��̟v�.����íVl���[�Ef���L�2oED�6�̶V@����y7	���f�rvk�[|e��^�!@uҍ�%s6�]�i����>�s�Ԣ6�UCL5BД ���6���WfR�	OB���'��z҇"��Y]��:b%�[O�zX�n��FX�In�)���Xػ��T7МKu�
�Wr��Fu:�,#)!{
�B�ͷW;+���=h�\�w34\�F���y�Q��9��=��%�V�g=���v��pbk6
vPS+^oٽ;9�6�-4��o����Sg*����.,�)c�^��q��`�\�j^��Ն�.�n��tGi�9���$\$�Y�r�ѝk�w?��e�����;F<4��k]e���5���_t��t:�)6�$�Z�4�B��vf��FM���5Yb;,��^�o�5j����ާ��N����C���@��.+=FQ �Q@��ա�Tڿ�9F�spd��T��V�$�[���[��R�Nd~��V��"pr�]H�G���/���7�@�؀J�Rۃ+��X������W�]r��i���� pe�I(�`
^���rT+x��k�^�ҳ�f� UȉKVR4:\"�`J8����wg�ZX9U<|>������t����3��:"��6�i*ר�[���-��he�e��
��NRٿ%��Ɓ}�M�K8s �@�	hs�wϟ�"�����UѺ�Hk	�1ע1��%�P��EBPN	E᧧%�&�BG��]��l��(�q�XnO��2���{oi'lWbJRW�B��^J4��[��ۤb�!o��e�4ږ�������i�("J���r�]�fފ�[Y�'[��D�ň
�}V��;cqś8�P.�$^��W=]Bm���5�mY�Vջm����9�i�1t}�=�j�/x�0;A�݊<��@�=#!d�7��vpZP���k���|�>K��v��}�M��]�,�wW�w�5��4���!*K�roO��
�sue�C��Wa[��A���0��4%�ޚ�L��Q҉�v�1�.�-�]���5�ַ{��ʷ17]����J���fs�vjծgm��WX!��wV��8`������M"�#�	�o+����P��	ɣ���a�˕؛'yVV|h�G��o%�c��8�eq=�U�/��u�� KgjF� +��R]vY	h�q����ew_H�ob7�zwk}�nj�WJ+ˠ�(���N=���7	#��,([6h�ݦƇ-J�^�=n� b���/�1*-� ��5�9�e�7F�0K�N<��W'�d���E؍\�g��B���fB�z�ұuL��j:�Urn�5!�Ep��a�B���M����KA����S��r++I�Ɓː�Q[�q��o1@r\ћ�������x��=ꔌL�Z�n\�V�k�S+�s��>[-e�~O_)�b��F�1S{� t���[%�\�#��,̸mq�W�%2��B7�I�%�A�Qw%b"��Ϋ��zͣ�#��
��*�]Ѡ]��v ��sڶ'���`�4>Mv+�]��φSO�bb���p����+�� ���]�rŪW�����݌�>�	�]������ϻt@�7�1:/t�)�Sŷ����sK�u�Vdf�hw8غy��N���u���<|2;�t�f຋R R��q1Vm��$)�7z Z�a���ξ����w�����B�lE��S����
	X�ُ��:4SY�v��u�*��窚��%W�]i�,p�����T�|���E�o�'X2����������Tl ۑ�O�vt\����q���:��R7r��`��7I�hݚ	O���<<<=�o��1u�X��j�>G��j�nJ�v�N=Ԭ�T�~����v�Lm�}�+i�?�����+:hR�2:u/����r�����qwMP��
s�D���(�m*�t�=���74Ϸ���{� T!�m}R�tf��}�&DԷ��Ʋ��t��)�o�-1mc��p'���'5��ۿ�4)�pSB��p�b�`�G��W_���/p_n.n�>�N����Os�W���w-QǼ�Z◢s�yJ`����vb,b�l	AK{�\�W{���J��������!!
윍N���	.�)����Or�Eg*��t�� ugp!^ ���ڛ���WAO�_q�h;=V��gh�]���V�W�-ngw'��:�u���ov8k�aV�h�����Ҍ�q�9nJ��A���n�����,n��v�-��z^�=���,M�/_�՜��nW^��O$�nV`���V���@�����������O>V%Ŵ+k�3��]V�����(���|;[�ǚ���K��.�Mg��I��D"#&���wv`���RT�:U ����1ل#[�J>V�����d�ˍfFE�kK�W]���Qlؚ��r�w)C�*]W�ؾ�s)�KΠo�v����s�ੜ䵲�1hN��t���k+���N��O+�n�5;�������ν�D�:{[ W���;~c�ޜ�3o� � �@�(P�* �"�i��������"h�����*3*�Y�*�c3"���,�"&�����������3"�*�ʈ�������h������*��1ʪf������
"�����h���Jj�����"")���i���JZB��(��� ��)�f �B���JY *h�&�����&��������JJfJb(l̢fj�b(H��(�"h)�(�)*)����)(*��bH��"b
������)����� )*�&������)�i(bI����(��"��&������i(��������
"�(*������!���� �h���� �� b)*��i*����)�����J������&����(�b
2��)��"��"�������z�w�o�V� �{�#8�<���@�A�D�ŕ.��/Q��xn���nwf�NW;���w�Iز����0\�z�I����x�nqR���L�N���S|�&���K��j�#�ᆛ��R��������f�4%!W�Omy���,��VY�{����*�PWc����LI��\fw�v_q�k�*��y�r��bRQ�
Ъ�\6���K�Z;��c�}~�A�K5/�:��.�:��<o/�r��F�Y���n,�X���`\g��I�uF�5V9�b�វ��e�.��S�)���{iD^��A
��=�;�<�xI�<y�4�C뫲I��ms��^)���t�xb�qY5�N\L��(aXbc(��F���N����/jX�8=*�)[N�nY~��ޤԝ�x�N�?1>'s��it��1�L_	V[��v�!�ѦY���n�Z��|qM���M��^��pnL̙5)M�h߯�k�X���V�?��`lֹK�[׋u���D_@1���9�8�ً�$��΂N�������_4��t���.�I�������)R�"L���=Ģ�W�p�K����W�d��7܈!�/��n�L��3jt�|����9^x*�p�̤����A����
	!��{�솖���z��\-��nw�4}�p�f�mj���M+����J�
��� ��d�N7�e+� ����hj��o�mL��dJ<.��m7�uX{CJ�y���4���7ivY'��]P.s���*P�cb�㚤a�N��Q��c=R��t7���a�3�tA\k���<�� Tyg�;�|)Vߞ'>�����;�:d�x+�]����s��}O��wv���r���~<�
&<A���@:
kk���h�2�l�z*��7�s#L�YEpw]s�m{}!i����MzW�np\�=��z(.�V˗]�sz<&U���o1B�۞��> 
��'��������.�/�Q�~S^ӌ���e��u�C��/V0.��k�F;�V*��jHm�A{�7�$��{�Z����"�~��+wpm���˲XΛ����߸��z�̹���m:����o��h�6Ū�)j]~��Z�pH��4Ѿ𤂽�x�(��Z�l�Y�s}*}���׌����gP�eD�S�m�5S7x.q�fu¯7f��v��|<�넪Ҹ�3���jjt�o���WI�5��7�Y�K�T�Z� ����4s߶��+��C�u�q*�8��}��'A-rB�oI�_!��csu^՚G{�wŊU��=�����{�wq�N�
=c� K�ҝ�6v�R��ާB����=�8N��5A��k�ճ�f�Ąpd�%P�FB&T@9��j{��v-��e�1��;s��N�xA����;F�_Ww���^jvI��i�{&>X�9l�T�o��q�l\K���֯%�
�a�=Bk�6к�׹Ա�~�)!嚮�T��W��#{���Ƶ}rcFmI�����M/j���3e=����W�]W�{���8((=0�\u@��
*��I��k<pJ�3a�P%�51&�4�ݠgT�އ���S����`Ue��]�.��4#����!`T�� �W�ˮ����VЮ�F<�L˾l��'<�{��X�sO�iW������]}x��z61���g�T������@�nLmV^]�=2ݓX9��8#���"�)\E�t��϶4u������m���UA�UEª��3��r(�;J]0G���<�eOG �#��T
�d�;^�1�k��!�����[�9�yz��'ް{yK��5;/�bp�Tv��*¡S*/��Q���@�Ar`_�J�q�T���;k��J:�e�	D�a#�K����Ȟ�^��41UTH�H�φU��N��[h���~�{����i�Vs��U���ԋI<�0�g�l`��6b{���0\�t�ՂN�X��q��>�)R-v�k��g�N����t�i�	�<�Ȼ�]�Ú�u��ט(����,K�G�Œ�����;��򱪳,�ow=��tD+�!s+��t��C�����Ѹ����X�b��L�V��|{%{�J�)�(�ټmy�Wt/�ȅ3Q�P_��~�+n�RҪ�>Fo���UI�A���J���3½���g����R��Ǌv/��[����z�ʂ-^��LS�z�B���X7�-��ÞC��J�^�<5"�[0jM��yz���AD�����`�q�ɔ+���������H�c��|r��Z>��yN(��M7<nJ�}E>���Ys�.5�y;�v��!�䍄��gpU(���@㼅/f�AN��=�:��nz�j���P�Ǭ	.ː=J�&�{ؕ��|'N����L_x]e��������/*֡�c�B�� Wd�(G��#ҧB�b��6p]�z���;KSvI��y" ������4��S�s�lp��g�,]{B���|=�1�s���Z�!��{5���d�(.gfTړ3&�&����%)��Ǿ��V޿x�p~���-L;�,�͹�˓"�70�p.6��>�<յ)��`L;�Q�<��x��ԍ�J�=���+�K�b볲J�:��M�ڋ	f�i���q� �@�]�b��uI�!H�x�aJ��ب˽:Kǆӂ�C�`8� e.����d��{Z7�3V��f��n,�eGT"�ӞIv�<��b��o��䅵���,�:�s�]�}���Ҡ��j`z�q�╾�]И#��uݕz�բ=���5�ݶ�pX�v�\��}]�n}��Jt:���W+�O'�smq�u+h��S;�z��kM�0��&"wz�)�q��ߍty�B�鬗:&F��m��:ǂ��`o�e��R���wlgV��H]�=
����ciC��&g��>�ݙ����D<�hݩ�9���'�~E��⏙�I��;Ռ�5�iۮ����]��9u�wTaJ9���N��0��N#������6DP.éY�E���[�s�~b����=�ϖ�`�D��� -�w��;�u9��1�7v.}�c���
Ш��j�݋���*r��r~ۮ���䡛U3r�䩼���q��F�Ys���t�P���S�f�dn�+�3�׭�.��-Fˎx�]���V����U�;��8^��F�w{�
v\�پΧ�1F�(bs�U�YXc�N����^���Ux!W�C����!D+Le���v5I����U�JТD���9kO`v���ͬ��Gt��Eu�NW��)ӂ@q{�6�c�m�m�]���T�^lֶ��[�&��g-�{j|dU'(��{��:�!bi�/Ek ͤ���ܐ�n'U_|���;�VP�`�[�M�J����Sq�+xM{"�3�˅��@{e~ S�[���O�{��~h���~�g]Ov�o�oҗ�����̙����4o����*yuۄ���+^��D��jj��0#�Ox��/ߗ\�>���	:M��k���)�*��q�t����S�1�}���^���CU._N�G_�Xd��,t�\w�B' ���~p?*�)otw	ڌK����N,W��Jlg��O�:V���8nU92��:�v�������w�6���1�	����x�^:�����Z��hNə��t��N���T0;� U�e��-ϽO�C����Ht�pLx.���p�����qH����vr{F'w��=�;�ӟ��M�]0��z�g��UW�z�'{\:T��-�Ɲt��U��9q�W�R��U�. p�'����n���Wi�8�T{��5�8�j���
O��R�q�N'8���v�>���յ+�y&�%@j��׀��,	��c�1����T��_[��O<㌋�G>*R����T��C'p��:[4@s���׊�f���.�.���m�Mu���[�_�D��nnt5�\ܼ�A�P9]���Nڷc��Q���e�:�}��Sxr:1�	I\�zS�1ޠ�0�����1ZW.�VW�7$����g�<|���n�UZ��.B�w+�1~S�Q�T	�U#ڤx��D;.�*�"9���1Տ�n��#���u��+����p���uu�����}:�l޹�ɍ��K��w�۩����#vB�.�2lNh�P��3Jv'V˭L��:�>�O�g'���yY��������c�Cٰ%���(l]Is'((��g�+�`����7Q��ohQʂ�f�'�b��މ췈��dعIu�V:���xc5^�洯;6o�[�˛�#o(O�w+.c}J���#y�
����Rd\ʌ���U�c���1kk���vm*����:.v���5؃*%˹!�NV���Q�[�\�51%��?&n��y��x��Kdo�+�Kτ��o+�LG\@�H}p�*C������GM���i�3�:L��z���R7=3*�5��xJ��pt�Ѿ����xX��Ƨ����v��!�SKҷګl!���]cq�0}[Ȫ��(�w��ì~��+�J�h�˵y�f������%I�ISs�N�-۫U�%dM;.K���؆���M� <y��:�j���gN�d�Y�h�g7����^�HT\��C`플����#V�춸�^�Փ+ q�:녩��9���EU�%uTv�S*��5�&jl���+w��Tq��z�M\��M� �Q�@�NM��l'{
dMޖ�A\��S��]W@jw���%7s^^
O�T�᨞� �|tR��+s�o��ssjj�{��59	����z$$��<�cD!pT��
�)�h)���̑�Q�ֿ[B���'/����&T���dX�No�M�%&*�p	'��e��8�\r�d>� oGL�����*,1r>�_k�r.�V%.^���=>��S;�P*��"�kb����j����dm���r�Nz2�9�����ve3½��\<%f��G���kTr��v�Ҏʉ���0�lt��q�x�Y��Яi$�=�Nc����b�ҽBxX;���<�8q��"�GM�%a��@B��
�C{���$z��l���6�r������^-$M�o(U3�Ð$V.��Q�.b&c���%_;�<%��+�6O���l<�����}ME�{0�V~��_�:�>�f=bK��B�i�sy#�<�20s��"�ϑ\����d�"�e���cE���C3sR�x��S}�G��
���v̸ھ��U��6��i�9�!�f�h͗���b1*n��v�)��e�|��7�IV����1�˺��7�vZk���������N:ה��f�U��f6	���pf+�{;i�z��:'�Ɋk�qڲ��hgJ��Eˁ�yI��[����u��\��෉%�HFA]�Jn@���sF�`T��WHݓ#�o��D-{%b�������*�Ja�y��ta3�*o�L̛�fB�\�S�T��#*}��"g�[1T��,�"�l��c�K��\��f�+��/�O���7���G��R`�Z����z+����5(�k���Rvp%A�3���6��F���(3a
Ϻ��Β<�j�	K�9@/{s��ZZ�C#:T �x������o��^��5b���J�zI�����\��bk/cnV��w[Wv�����gfR��D�&z<��B���s���l6�Օ8���>�5W/W��~�i�3�#�|t��(vWV�y�l#�R\��Fe��uڪ�$(�q#���$;w �@Sqp���?3+J'�a����g�O�ufz�	[����~ޭB_tv����+
_r��Ȱ��TIq>fc��ѭ٨[.�7����+&NR�����R��8�y>���c�a�o����u9f���)ցS�"�Q�]-�|��uwS�}�\a23N�̏V7׏v���hӌ����=Wns9qe�;J����w��(�r|�L�ĕ�mr��Ƕ�%�α�����Y۴��Z�A3p�/0ΎN��2���X��l^yI���L\6}Ckˌ�����զ%UE�]>��Ζ��s�d=����,3v�����N�E)ffd`\7s�
��I�2��!���&_ָT��u���c��,�^�G����e�j'��Re.���ڲ����l�����]8��O����
���D���]%S�!K����Ϟ�7��[8��E�Y\/��ۮ>�ω�E}����ി���? >�"&H&j�>ٺ��(B��[�;p;��v{Z۸'(�ɛ�Jnh߯�!��@B
�Q�n`�^Y���D�&h���C��W�_ʺ���Z6#;�jEA��=U�!�
�J�G���'q��Pb�?T�8dS��jx�w�T�}=Q�ͬ2Uk����Jq*��r���q��m���[:6Dܦ$��9֯�`*P�c<�<JK��9=ĝ�����
Ds:
pf�{2�g(y�x ���jw_ߞ%s�A��.��f`{��T4Q&6�QRct�Y@�e!�hK�i�E*\@��`S�Ԙ��sy�a�S�!R�Zp3Y�1�Z���]>�08���2mGl��g1c6xE�q*�����q���:E�nUx�ttwEXFZo!6�e�Z�����4$/:��Ww)��Q�eb[�5�WM�Zv�+V��|�C�f�hagC����]C!&��7snq�c!��ιЩ�μ�xK84��V�oyT�xC���i�'-(9�:7lP�պ8mq�A�0���;J�d�������� �d�4��;��Ca��}!����*�seN���
��[F5�q,ΣЧ����R]�@^��^�K,5���lt�ocy[Ҁ4�s�,h.�]c��m����c�B㗔�v����W<Ҳ_j�.v_;y�հ"$ʊ�Jn�]�.���Ws\��a���N��, ���`��g[��3��L�����­L�<�ѽ���{*0\����MAΨ.�x뜖�Kޡ6�g_}4ic�{�ֻ���cD�u�s/��r��D�^��ܴbl���h 5�;�|�^]uOD�T���,��iEJ��XA�*(�NҒV���ԗ�t,�}�\�q���O�t�wl^�����MGX̴�� ������Fg#�OU�|;1Դ#�[7�Rjɘ��j,`WT�U�Z�[���ڄV���kj�Z�li���(D�*�6�L��up���w]�.ǎ�PN]�I��v�>���û��-!��+�����q��s�&���n�����}��d�c���Ұ
Clr���٘�P�ո���n�h���{"�!�����i����6�������x�$�o��*oDɆ�ub��������=���.Qu�[�da���h����|�+�/�|�J��������I)C�rz^1b�&>맚�Smv�9�1Xw8-�;v��7�P�D�p�V+��S�d��A-U6P��:���>Y¦^A�L9�:�N�9�����es��Sz�<;I���*J�� ��Y��=���-�|��+���;�n��r�2�G��-gP���Ӱ��u����-�r���_\�Oc�L�6�ڔhc!��:��.U;�ek�ny�sT�t)q��#sp����ƻ��]�Z�"h�U�wb;F��/ %e,h��zM�`�U�2V�c��X�RS�۲2�(jS��'�����¹ʹ��"������/�-E�ғ6��ud �Yu���ֽ@�f�;���k��6r�s=���CC���ǜ�,�x�Z��*T2�w}A�Q_j�U*�{GqN��G����&;0�pK�[��/{��%!����I$َ.ko�(��h;Y+ƙt����z��㾽�T�;���[�8	�1�S���D:�s��o[̟8���^�R����1��C���1:���!yg�PU��M
���uYS%�H���,AX�g.΃�:�U˦m���zd��8]]�]HH���'*꫺�����
h��f&����(��)���)�"�
�*���"�ji"
����
(���)*�h�b������"��Z*b$��*���
��*�����bbR�����b�(j��� �����R� ���X���
J�)� �V`((J
�J{�ª()������!�hi(H��
���hj!������i�)J���h)�
C,�Z��H���"hbhJ��!* ((
j������
B������a�*j�������b
�������"i"�������(
ZF$i�h� J
j�)iJhj������)JB�(�&��Vzif����!�hg`��z���mIZ}�����/��j�ꎸ�p�.��h���������`̗4��J�_P1�h�L�L}��%Q縚�G�j�~��bӓ��:�7���9m�}��FAְuQܹ��5	}���NJDD!E�'_|���}�ꎬ��UU�����c:n����`���"@�9�!���Q������.f>:�wr;����kzL�._F@u������ֱf!�ۯ�rN��z�C��S�{&��|���%S�r����J��� x��ï��_A#��p<�[�j]K��k���.kCs7�d�\�e�h��?s��`�:����.��^��\�~�OZ��7R��}GPr� ���g�o�s��������%Ǉ�"(}"#�:�\�!��'S����du	T�}�èwHu����<�Q�r��1y�$��������2y�t�~�2���]A��n_cq�R���x,�{!`�ʎ��6;y�6�Ǧ=��L{�7���b�:���>�.������y����m�?BS���}͟��=F�+�kKEѨ5>������?�A���|���5�瘺���I7��?~��������=UDD}��G��7	~��?f��\��:4a�{�=ˑ�X?F���j�����~�.��]��_�L���=�ח���O>�׬��Q��<�A����w�{�~m��lz��s����x���L`�$�C�j��C��jMG�u�w��}���N��%�u��G�����2{�5�pu�=@}<�?y��!C�{��~��	��������"��UȺ��wA�?��xp�#����ʗ~��m<��������;��n���ϐju�y�Z7	O�w:�a�<��*����7pd=o^��F�a���>��$��fҏ��;�g>�N����c�� ( �o޶=W1�/��!���|���6�/P���i;���rO�<��u�.�U/��5s�P�w��������j|��S��u�#�:�#R������n��,#[>z�xs � ��u�y�k�Zr|�s^�r#%������]@e���u	T}.{�}��5	~ù��4�~�%��n;��S���@w�/����!���
��R�{�/��sV�F�)���x�l_C�s.�%.2�汔�v�DE��c���v0LwY��h-i�g��bWt:�p9*��-�{�]Xt����*E��\��{)L��oyv �re������Oby���=Ypu�j��րk�{����hMy��=��>}����?����/wѸJ�u�%�b��d�k�.�9d>����%�����y:�I��=F������Q�vu�����ϱ�����s[�!�G%�@���������wþ�ٮ����rw:�:��;�u }FK���{�C��?�h�����_����d}����`�K�+�����cx�ͧ%��}u;��߻�\׾���OcP�_`u�����:�Pj5r�X���2K0�캀�2;z�p��C$�y�7���{>��ϒ�Q����ד�ܤ|���g��D|X~�s��>�F]絭�~p?C���>G�蹂d��]}����?BS���ܛ��P�fE���Y�K�Zr6k>�����'����]K�Y��%=˝y�:"<#�aG��+�'�<󥙾_}��|��z{���yj|���h�#/%�5�4&��~���u�	������������59.f._F[3�<�����%�=����䚏c�
��4���[(˓�k�v�rޝr#��{&���c�%���c���A�{oN���k����\�GSܹ�?s\���'����N�`���7�V��2��:�q�~��9.NK�>��naV,���V:�VG���q�ď����C�{��s���CS�Π����dj������y'ѩ�o[��2A��\���j5}17�2L�>枣��u�g�l:����H��r��Vv,�jv������;�P���~�������/''r��b�3�^�S�x����z;�݇[�2~�����I��5	]}��9���5z�pPy��w	t~�T-v�7N{�������|Fu���}��z�7��>�F�)�3y��B];��%꧹ro��r^�OQ�PF_��=�?BP��}���~����sk����6|�=�k���o(����|I��4?��p���.��Iw��%��I��w�Q쟜�ѸJ~�d�����BQ��:�I�I��&���k�䟃�:��2{�?[�Ժ��2~��{��d��%�E啟���V/f�5I�uc�k4{�v��]SB�@��줏oe��xgW��%�Oʦ���k/�j�©y�;5�~ʾ��#���7[n_V^&�/��]���m]��Le�S޻Ϯ���T٧
��"��{pIs�8��kimES����6�Uw_9�U�B��[�9�觩r>�w���sHnz�*}���reI�=�nF�P{%g�'�{:�a�GP��~N��z�I�j_�c���2��?s�w�:�$��#��$en�u��xK�� T���_�FI�o{MG/%��~�Π�r��g�lz��9u�Gg1<��ܹ_sGq�.�'�?{��9�^�Uѭ!�y>ڃ#�5�	����~����害��y��=����䛟#RN�S��F�����`�h���sg�~����7���>�C��Ջ����]G��4=GP�G��;�I�x<�P����r��s�}�;�ƥ����Y�K�R����M����?�� �@`�HP�<�n�/Q��L�u���1y{���:�������o��J�:5�7�>�P�a��iy~���j9>k�?�P��G�sO��cP��ϯ��]s3?ws����������[��54�Xw�bn���N�o%�#/���}fHS����K��pgz�R�rkϵ�%9.^�����I�2��`����=��^����|�|͹/�ٵ�h忳}}�!sRF�#P�u�5�O�ܞƤ����� �}����5�h��@}?��ܛ�^˩7?F��r����7��>�=˾i~����7|���ow<;�ˮ��>-��������<N}����b����T�'�V�����d�zkZN�I��5/O��}�Q�5>��p�KEsG�j���5;��#�멊|��}������>19Y;Ϲ��r�j5	Tq��mz��j�ϴ�9.�|���4u���Z��˸�/'�|�y�B�������k�C�S��b�}�Cx���1O�8A� }Gq����nf�׹��y�^�����Bs�oh{j{�I������?BS�~���j=����a��C��y��ְ2�8s�m@n2{��?h:������h��.o2��(��9*J=�l�����$k� >�����؝�};��tX��_�~,Pf���JB���b��F��7ap�ޗi� Ty��&��sv��D*��^7����)�G�{�/uf �m�G�XG��F��zT��o����+��<�Y#��s{��0�#�e��Ӿ��{�qD-cW)�!��n���q�SE��v�^�<���}]D
�� b���O�x]�k�ȧj/Md�ّ�f�.�������ރҼ�G9���j�)�+��H��@��u7r�EX�P�ǎL(�).}���oj=�ש�|M�yp�Ȩ�?�r���҉��v:t�^3)����i�j��DNt��'/���.pl�@��R�½�hz��:����~Z_��=y��E{�_�u�&Ag�����Rj�f<'�m�;�wz}�r��� E�عY�1)+ʀ���i��0z��<��JQ��']{����OCS{y~ސ�A�+���Q|��Br.)NWN��T�Wu�:��F!�I�_C���:g��fsv�E�8*���;.ts�r���K��RD���a,JCS�5�����Ux}�x_�'f>^X���F��w���'e���K�����.Jzu�~&p�c4r���ٕ�>��'��'MEt���H�`�¤��=����$ں���ᜬ�Wn���1��m��]�r�̙�JtM���31��2����,�hl��X(g )�Ǯlq�46mFH�4�76E6j�./,�C���5�1n����Z^R{�b�*fE��$fP#s���s����r.�-f\q�P	%�NZZ{��"�%���z�}�vMn���-���NFwt�a�8j�s�� l	��槟?�]sD��z�J���' x`���v��-�t��{qT��!��8�SV5<}:�r�w��:�XB���o��:�A�Y|����NBB'�H��5
�1u3�WOӝ<�ƹ�S��t�F=�aC�f�eNq��y��H���z����:� �=E���P(뾋�V�{=]�E{7�}#�e��&\�|�[Gt�]����0Q�� .����`�P�1��Lv:ܔa�%����y��O,��+��}\�x!���$� �^^��2$p� v��F�Z�������;�$�d�D��H�Ps��(sJÙ�ݘ���@��@z#����ʦ,�a��#Ԉ���u����7�:�ntAb9%�{�7QiRs59����C���&�SW��ѽ}Sur�֙S�&u�j��!�^]g��Ö���r����Կ/��]��&�1�TQ�]۱�������=}�y^��
P�^�X�]f|�ưp�Fك�������#�AżiJ�.�2C'�aR�Si��Htc=;v��J�F��<��8"��>ύU˷�:Bm4�(�Z�3P�`N+q1171}.��M2�K��d��+5d7*ŭ]ßE��^ʼ�]w4���t�W��X�6ڝb�$?��c?g�`�V;�n�'S���_}�X�X���Jd���`��oe�33�z6�n'vB�����#����ͼ�	o�>�3�܋��|mZ��Fs__�7��z���EWYc���:G|N�~�c����f�%Cc@
/�_N�B�=�W�{��E���Z!0N�����u�VI��ej�U��<�59�[.�f����qD�.cE+򃞔�o`o�j�D�V*��_�S�a�j�����,�����Jbx��Y�3`{��D��9[mg�a���w���ȷW��m��GJ�A�Q^�B��E�k�����C�8��ۍ��V^���\XQ��ڝBͫ�W�}���Q`)32��\i���I-���������i�蒢�����,��:������k�}��VPG����wM/�9��+!�}ӕW[ɹSw`��c��g���V"�MQ��M� >�~��D�ҕWa�֦Iz�9;F�N�@��.'=�T�)�U��{Y���WW�ʑ<���Xc�v�F�"���wQ,-uc`�G����u
!�z#
xg�N��Y�Bަ�8�y3x���Kl�$���3t��F�5cB�ѽ�znhGN��4��βF�k���ܘ軫i]����f�I�%��%BCqV^�'�`����]�{�0�~�&�Ok�����fN������FF�1��k�&4!�O�=��W*�h.��89H��]��tܷ�.vШaULv��/*��6�?����ևNZ"�O%�9^�)���ʊ�Nw7�3/�k��,����~FW%��!�K�Չ=+Ƅp�F⿐����G;Ҹ�H"��&��T�qqM{"���\H�Wl���?5�vP�^�����
1ɕ3!��4�:qmvd�~�����Sʘ�}�LS�ThS�ډ:�i��a`��{Z��i���I��/	��\j�"B�׽y|<&J�q��Ad��ٱa=�Q�\NH�2���ؑ�0B�>�ƻ&K�9�{D�;�U���*���-����|��	f����4�9>���&�����W&rm�8ێ�+��>]!l�F�t|5N#���+�M��뵫ϙ�x��z��"�]��q�*
�ep�����1N�!�j��� vE�b��tb�[kd��܄�:��d�j�#�hi�m��3�$D����+_����\�����C!�S�9���Ò���;�v<;�l-y�$���:*�V�_y������L����̼�JcBΘ�a���)�qج�2�;��O���*I)-��9 ���ݵrT�S.J�{6Wq�.�VE��h�Y��=�����eL�y6�W)��k��{�+xѾ|ͺ�)di�
3�֡����3��Y��gfT�S �շ�+��gpg���K_8�gJ/�/���_�*}^�6��:�#���>���;�}�y��ڕ�� ��Rb5s�C�x�)�t������6.i�r�m��Y�0���$F(�J���+��ހ�r/����O/P��i�ʻ���mD�#�P BGDd�3�U�)T���{�yV��Ε���^����9aK;^zo��m�2��� �T�&#�4B���G���B�t�K�3"0�=u{�q��PJ	�,%��݋�um���D
���C�ҿ�p�̈́pu����Օ��XsɎ��͟aT�K���@��r�>���GA%iӷQS��+�.wR�P��O\כϏ]AW�횢�x G"��[�hz��1��I������J��S9�]�7�A��72X��&��U���,<%��N�0_+=䄼���yP�>���Bnj�p���p���Y���j�w<�`Ӓ��s��b�,��n�Y����~+����*Rz���ķR��I��~�թh�Ƕ�r�İ�?���n�����!�V��� ;�����i�OT��맗D�#�㫦��S^�r�,ټ���V�A��J�U�!+[dog`z�B��3����c�/��o�}MV,�����U_U3��ɽ�D�U0����&�V���tj�~k��x҈��t(Ю�c�
v\ވ����:�[���~�mA�W�y�,1�
�\�i��q;3����Vx�ޛ��w�	�Mۚ�<�ڸCWc\����|^ٌ�Z��ٕ��dW��q$�+���3b#'�3�u\z�z��'k ���%Yn��ۀ�;��vzǟ.ʃ�e�3u)M��3�G&o���K��h�۲&���6�`����
���`ո;Kp�%]Rɉ�)�H���u嘚o�o��x;u�uP�]J���SV5<}:�r�w��:�k�Uk��9Z�Bۧ4�jH%��p�� ��A����&5����zl`k�%%�l�̱��leT����S���
���eu7�Z� �-��u@�灉϶|X� l5g�͜����;��s�X��{�ʮ�q8nWO��
5D�@�'���26�"��v2�JӺޚ�%�)D ࣱu��)�j1耆�O�ϕZ�T��4P�gy�,�k��v���zn�麓
j�����\���j�����
�1ZR�h�<�=ʸa�sx4�z���j��
�e����]B�+}�]�/x\����5�����(�����ލ�Rʳ�!y܅<�y����"�R�q�Z�u�Dz1�)��c�g9$/8���{���+��Rg����S��'�;�&;;�5�J��
� E��Ny]�"`#"rV�S���5��s�;�=[�쮋wE�\�-���XHԊ���L�IP�x
����+c�*�ߤ榳���U�\��: K���'{�K���Ry�#\�L�鈮�r�Fo˫)PU�gr��B����ڳ]�X�k�l7��ja�b�c�������hBou9:�tS�<�B�]���ez��5��L�݀�k>�Tٮ�W�����o�����b������?#�M;v8��Ob�vm�@i{�ޗ��XNd*�ˣ�:QXrn�ŋ�WD���Um��5S9!DC�㍥vF	P�Y�O���^ه�[R;�th�fr@�In�ʳ{z��RSgP�{w�P3�e�"Dg�v\������j��u�{U��v+�)��T�A�&�>���{�`��	`���ڪ|���,���Q�;�TR��2׸p�2.�v�1ٚR�&��T嚘�biA`�\	բ�^�W]i��C<�>��~��hs���}��-N1�\V�A�Ȼ;�3�TI}�������{YW)KY�Og��Yܦ���u�����@nGF�o��sW�卮��0�ւ�vR�x�[[O�$,�S��9� ��#���=u�֔}�"}~�LV�>���f�27�`��n�W3�	b�z�Y`����u,t8_wan�Fkne��t!+�]n�;b�X���������Ś]�S�:�J�i��g>�>�I�YS;	w�3Hތ6�f�n���|��͛׏�0�*P�#\[�6�=�NB3�ò]���CY0���B�5��Rc8",�X�W&�*����X�g&D�����B�ѝ����R&��iU9�I"�vhwT�M�fL�c�Ĭ��aG5��Õh��cŘ]���n��dh/���C�詘WJ%Ċ���z�s�K,]ռ�pJ80*��8���[�P֨tr�$��:�OV4썴��y�[oP�+p�X�C�mu�����;�#�R�K%�CY�LD��o�WT�-4� �uL}�O!溺�lK�[ne4gm�ᙥ��]o|.�v�I2N�kG9B�fMJ�����p�v���hҬ���g@�E%�.���d���:�r�X��Z��d��9VS=o�>�j��0�P* r�	���R-b�Jqgm��Z]N�S!�֖�n���4��ghU,��>�m���R��46�+@B��FƷ�@�Y�!�6���p
�T�e7yZ3W]��������ΛVذn��V���[��,q�qH֨)v�9[��agp��4�+��'vt�P�u��GF��9M[E��P�kp$�9#� �b�x���(�;�7��f����Vg��� ;V��:ʮ�İ3���f�uM�j�S����Uf��nW5f�:L�C
ﳩ����:�7E��j�ċ��84V9�T4��P����ɺǋH���Y�ʌ�m�)��OWa�$�[��ť	{Ϙ�o�˯�S��T�Z)�[�Ұ$��V���Ś���O�Z���K+������k%C�%�fTj�j��pdo��:�`���ϖ���򧯭5a�.��{c.#53ۇSgy��˅ʑ�2��铸���Βh�[�A)v�g)1?[n�Yٷ�m�3t-��<'w&� +p*)�St�0b�;���.f �7bup�:�.+6��v�H���{kd���>��Rɭ���҈,6pm�w�j�#6���k5I�4�A��:����F٨]�@��N`��n�)�Z#�T��8�h�5����W=U��`��1��N��E��De��^�}�(y��s{v!oY��:��{���Z������){�v���G	�Q�JK\U�7���JJ�ncU�3��R����r-�r{�����eݮ��c��N_K5f��]�VnU���	m6��J_X��U�7a�4�>�$;�Ǩ7����

�!�
���(J
)	�*��(�h
B��2*��h���
h*�Z�JJ" �"!�H��((�@�#%Jh
���(�)b$"�
�����bV����*��2C	���F��F��!rQ��(����Z��((i)
�j�2hhC 
r�)
c#!2+ r\��\3��i�@)ZF���h\��")V��L���2JP��
�� j�h �i����(rR�������iiZ���L�3������;�F��^r��v%�)��d�!�Ի#�����C5�8t �wE:���1}ݜ����V���6b�}���m�Ӗ[u[�{��<�
�T���>:I�TV �i�*�U���ѯV���k]l����lҪ����LSr3Ϫ\� ���O�z�H�Q#Dp��"�'.���ܹE�.M=[���Rˊ�]q��n��Ĩ��k&�28O�9UJ� �>`ޙ�и��m���ؤ�X�Dʱ!�+��`T�)�U��������Ɏ�<��JD̨{�q��	hzo��ג�;�PHG��v/Zj����ЦcD!eO�=
l��{n����8�Y=^6���� �R#v�V*T�(p���ordv�&:;��|�gL;�<�v�S�%w��T߸mJ}�Y���\��C�K�Ո�z��
6��qeVq��oXe�Q�ǆ�I����W�{DT.��;(D�>�u�5
�'�E����
�];G�R�y�B�VPZ��l{�f�LPS�Wy1O}Q�^�I�i�1�!W�nѾz���͞�݈{E;�z��6�,��,;�@�6!eR����-?TH��9Z��������͵:�u��qn�2\b�)�fw] ��"�f�r<VU��luHT�����;������m��L�:'eK�RP��-5��U���	�݊wvc8�J���8���Q�]7�R���p{j��|��z���0�l�K̤��c��NGL��������Wqn��$�ޜ�������\�3Ӟ�k`Rf���R�\����v4�:�0���"�k���՚��ѳd��<��b6�[U��U��z�.Dj�����ޖ��J�Y�qyN�wL�Y��ӿ
��A����<'�Ɋt�;(Zc��@c�KϮ^�����\��5�����;44�m[ZX�+6���QZ�"}�>��
��u�\ԍټ��"S�����v�Ʊ�M�Ƴn ��3��y��K,ɕ<��6&�&��K�]ʕ+Vԉ��5�qǏ�L�eS85����r>��!�YDv�<3�e���� ����z5��H�C���P����nt-]��M);8���3S �7��yx�a��t�9����MZք>鸨1��2H�P F��2v��ЩZF=;��w�����y#�+�+���[{+��=���:�������^�j6p}�ʸp=�'�1���GvNbL1��g�̍s6��6�^��w8R#�|t��.��4�Z��ULt�� Q��FQ��E�� ����w�S��J�k���p�z�lf�1u�P��}I]II�qB�E$�	N��<!+��>���~)�V��/�o�#7.z:��7^����H��|󣁍�㴯���%��E%��W2��:A�́�]��������>�o�����#��)�S��G��TDXʐ��J��������hax0=�������ɷ�^4���J��N�����Tlh@���ꚸ�c$F�aԬ>fX�̋W�پ��c�bā�\!B�u��3�� U�$/��n�;/)�a���h�^[��eP,_�Z����ţ�&�WIsc;7=�C�.b˝f�ŕU���)�8�w������}�2)O���͡j�F���Y7*� �߶��6�zy�躝�qo8�'nt�%V����}�Y�8�2���^���8���x���
}P*��'����n߭�2�Z���b�!;�2^Q�g���d��&�����䰷�Tf{vx�=Y�_>�~<$	�k�P=�	�U�MR�#z�mW��������9 m`��{�,��k�m=M�I=~u#� ������Awq�'��NFj���a)ڑ�E=��M����EՏ���	(� ͠��A�u.
��Jj�<}-L��^~�n��epO��)밭�=�}ӟZ��j�P��M��/z�{�4`u��٣F���}1Q[U�V]�.��_:g�]�zV�`4�gRF�)����hذ�Kf�k�����,��v����>��r�l��8�N��n��x.���[�-�6��U�}_W��]����7הv8�N��$?�O�gA���g�*�]9��.=���E����Oc���&�R΅%�S�m��8=�H�t7��� � [5��������؎���FT�ƾT��r�ڥ�*�&�+��p*�~�`��D�$�05c�J�h{�N�5רr/���{B,'� ����F�[e��:6f��y��z��(!��;K$a�Ղ�Z��/L!�evz�����=�2�����
��D��*�W��c��1��+��5N���C�'g^S��wz�w�
��U����H�\��]$��pHب���L�����W��=Iq񡼻h�F;|7�ئbb,A�Xc��l�;ؼK��㛁jO2�`}^U1F�y"(m�="���b�o\	���� F��r��W:��¼���{�c�hZ(Λj�sZ'c��S�ۨ?��Lo�W^?{ku<���� :C��B��^�\,qg@5���^fz_n�T<8x�`3Nv%*|陨�ƾ�7yu��g��[7�}~�+Z�:%\Eo��2�{�euԩM��ga\�fs�C��k1.�Z��0����fc��Fx�^%��[6��ݐ;)nmp��ϻ3zB4��Z�)�V��)j&�p�wv�X��ܷ�jw��m��p�kRh�f���ym��qd�$)0����R3�Y�����^�i�:���ީ[2d(����4R�#�q�ք���=�ڐ����խj�z/k�F'�3��4l<�wӞ�����QK���_�T�ocx����}��S���y{z�	�@p~�%��Kڪ>@h�>�Cc�026xU���<��$+<�Ε��]���y9Q�lJ��51%�^�B��E�k�����g���M☜]
g���w����%����	�qz���΀��O���!E�32�k�3*4]PQ3&�k�u�����d����n��'E��W��Q˅1���'�j���*���%+��U�P�1��KY��b����W�_���x),1M�ә�TFq���z�M\��M� �k��Ω-�W$�~�߸�[�Τ3$.'<��R��Sk"y7��x�;WynY����)�Cx:D��֎u`���r`eJ�q���oD�ij\ȗ^���8��4��:	c����9�˯0Ws�X�ۤ�Gl�.U��6�;=���Z>塣W�+���Q<�\���.[vx�˚�ae���h��r�]�͋��@�����*��͇-��&���LޠSүv�t�F���ڷ6�wڍ,��g5�B ��%}�]o>��eMr�d=�q*��'b Bx�u	 ��U�Z�4���a���s�Т���T�f����T,���o��K�ԥ����r��p��'.&��3Ҳ�S��nv�J�}��J̸	�:��<���l�؋kr�NFPGWl�\�Jթ������iIub�'�= L�]n��S��1�ySX�w��������`���߼jӛ��'	\��VMf��}ӗ#`l^�F�ח�� �㼤C~YT�g���`N�$X��߲�Iȣ03�M�w�0����X��պ��Gx�,>f�VL���EK�s�����܌@��7S��[��������Y��ѳq/c��&#b�|��O��
������n)�ŋM��֏K'O`ӧ�w�E7ݪ
��� 4*
�tW�XxJ~LS�\���ф���/!U�Y�iL�txsOT�9[n�5��d&�����D@4��Z�F���#Ľ���o����/_�Ã��O6�1�\���3���-�ٕ6�3&�0��}�N�5e��\l��-���L�*H���a6��r5�0�sύ�;�}�y[R���w%�B�5cNi�#�gZ�Փ�څ�򔺚�ӛ[7f���:�۷h��V��R��3ck�</l(�nn܁����J>�OI�:�u��o3��{���������$���5[���(h�7]���#e�Q&�i�[�������L�t���Hr\���j���|��.%I��%A�3�f��cy1��r�?_�f�E��f�_YjT�&瘇]S�#O����s���(WaU�������o�w���T�541�1jpf�-G�w�D%�Q>���h_UT�� F�*}��O�x]���{��C�+'3.sPɻ��Dl�e"��I_�P��)�+��Gu*V�E��is�5���%L�Q9��(��8��1����)�W@R���",	�H}]7J�ƙ%i�t1�{��Q6�fUf����r�܌�L`�f/Z�5G������o��%����Tz�guOP�솧g
y����Xo��l�Dc�1J�L7K/0�'Q�Ʃ�m���`[d�wfӭy�#e������yP��6}V��n{U�[��`�<6�(��1S��w�����!Qe4��n���v{�t��U��$��F�5|-X�M_�Η+&�ָ~�\.��y�K��[u�a���Y���;g��~���x�X(b�vp�+�x:q;3�����I�^���N���.��D��;�Y�T�>�,������;>�:�>�ube�F#�fC+-l0��V�^�4x��י��T����{ ـ5�q�9|/�:�ns�v�]!E]���A��)�:�[�z�e.��exY �D�B�Fa}���{��M,'[�6b���QI�wcT����K�1��9jt��]�^ȩ��^ji����M˻ӇOh��2U\��2P�DΜ]4��+�>ݖ����+ϙˋ�7^�V�з����zh�I�L��AS~]v�o�����
���e5n��0p=�<&ӆ#J��O��K�����`	���3Ah��0.��S�H�5z�>��\����[ɭ��y<��d^k36�(~�[ǽ'�� �' ����]�Lj=ӟˏ'Nu*�4;�|�|����U����1�X�1��8v�9�!1X+@U@� ��C��Z����Cԯ*����L]Hߘ���v�;&g+��b���F
9�u	��ctıP����%Er�[\.0����
8��yO�Q�0x��� ��Z�P ��*�}}4��Y�EKD<Rz�W(�.N_\�N{��^Pw��J��m�1*� F��'��Y�0����T�-�2��[�8�����ߧ����]K3�&0���+��Q�<����1fЪ��i�TG���c�b�'�p�eG"�����i`����Fgflq]t�:��+Y�4���֐��c�FL�Yu��J�9�h�0�d�z!ڂ>tx�Gڹڛ^5/-r�G[45�SGWW,[�\R󑼅�c9s��w���UUW�+������@��UW�Z���1��l�{�Y�q����h��r^ݶy��`ajJ���X=NgU�ь��c��چ�����f�|���u����sX7���3��Fۿ}��}��D��
+{�ྜ�e��U3.��U�+�nW�f�i=S�}�/����c�鉉��Ë�vXQ�3Nv'�]55�N��7yu�5�=�4��YnzVr�.�׼ѽ�dצ�l1R�ɐ�#|u�q�]�q�ƾ��0�0�+jFݗʚq���zC۴zU�L�\�d��`廾����� �J��%�s)_�
��c�q/hd�����%�xυ�-4���ti{UJ|��bv��5P����О˔'"�U�ț�̄�:��d�ZY��*4͆�@�8,��+�X(WIkБ����LWA���7#�U*ՋiL���OE �PM`g|��O�쐢���ʿMt@�T�q���3k���9��z絆},ڮ�{��k��>��v�v��k�T��r�Υ����Y�ۊ�*�!�Ɗ�P{Mߡ������w%�x�D�' z C��<��R�;����\� k3݇R=�8An�d_�+���[v��*WTU[玓ν<�nº�ʝ�1��%�U.j�.�N������vF�Ru�:��}��U�� ��>�-�#�Ff�-޴��"p)�{[�6�κ�Z�K���@.zgZ�[q��o�����,�z�ESK��lXMڡ��h+
kSdW~���g��Ъ	���Q�\�;Ь�X�	팙�U��0�]��qǺ9�
۫U:��6#�:�Gj����[��u雇"�:8"��maJ��N
	ѯv�(=6�پh����䐖���V�Av]�V�^�,L�ucm69�����d�ZᶗFQ�]Fb�%��b���|�����K��Ô��rs���z]�{����e�L#���7�Į�콌�.����/l�9�}N�=����;��s����6�ʉ�V��gvju��v䑺������$V>Y&�)��
e�s7vʘ�Sϳ7ӛ֒���6��݅a�78ioP���
�.*�����˜W��#o�����o�T�k�-�2��8�W�QS�C1� �� :�ͮ���=�^�ݢ�BVK�.+��*��`�u�+3�2_J���={��}N��SW\:#ڭ���'eC������vK��d�LӸb).yh	��d0Q�<��z��еKhNR��C�t
[;��4,�(���2�׶H��!�נfE��v+Ѕ[ú�"�<�WY�H�Z�8��;'�}t��f�lQ���}(��˕^�E�y[�:*����x�@�y���Ƃ�DWʍ�R�i�u"��x{:�A��y���A�з��zh�W-s+1̎l������,G� +�D*�_\���f��1c��V�9gū[{��=���V��WG��9K�F�]�C{�q���~�q��AU|�P׭�Bn�l��K�9D�����z�s w��v�����/w{.�q��*�(-A�W��O�����U�9s�g|yS�2_kڶ�b�x��4�%e\wk�-
��9��.Q�.-�!��>�A]4�L�;B�tWb�i/�J�tW+�+No�#��Y3W;��$�]��!�y���X9��lTzoD-�se�h��0Wjx�j���؟I�2��y-�xNU���t�}ݴ��@�K��l�/^��c�/Q��y]ѩݝ;�����`�x�	W,��뜳��!��$���s)�Õ;"Y]Y W����*m�/��2�Y�.���*�Ii�hmۮ��KD\�{���tJ:Ҫ[$�Iup9��r�sr�{�r�y�v@A��屯ssM>���dcFt����=D��>��e�W�3w�:�N�����X���R+���E���
�}7]Z�|��WQJ'i�,u��fR�2l��5.к�J���qCGL#�=�]��Ҟ�&ur�M�ݬ��ή��6��s�,����Cn��y3i]5��9��+�fԝX���u�EWy��B�4v��mq.�w�%´�$�+������J�*�V��?o6��Ѿ�\��n�@�������#p�te��m�&*��÷��� ��L�O���.�霳C�v�s��^gr�v��`�!���H�Pr�K�L�%�)X\�]��^;ΩRp��W+����
@U^J|)�]F�]ŎXw\��cg6�UƓBh�i��|nQ�E
%���ɏ)������4.�h��E�Es:��"Zқ'0]vS��HP[C>r�us��@�'u�1]�c	���9�]@[9���[|���u��ٽ�V��EM옗iݜ��6���#�t"�� P��t�*R�(���\��FN=��fY�f�oS$��L`Z�F���Ke��J�u��-b9}[R�g��r��J�����p�		bi��b/�=Z�ܔlllﮠ&N���=�]�o��)��wMy�^M�o�[�jv�%�V�A�_�AF����y޼���s��o���ݦ�� (�U�()��)���J�*�D�i�(J
$���B�����!
F���(�(�)��)h)B��%B$ZB����A�B����RdZZ
�
@hJV����()@��(��b
iJZ�)h�
A����X���i �)F�JA�Z�)F�)J
F�(R�J+����9WN0 ��Hu+��ܕ��m���2��!uj.��󛗬�/�/CeF:��rU�X�9��T�㟞�����Q��&+{H�
�k]�v�޵�j������WN���"OSuq�oVQFw��GQn�[Me2�J�i����A�p��j�3�=�=.]��%j=tf�h.�SC����0&pi�����V�"k.�hn�z�h�����'�F`�RJŕ8Kg�k�B��t<m���b�f���f�c�l��P��f*WRSŋj�#��4w�ƛ�4)���z�[�27����^*�#�B�Y�����<�T�ӣ�).V��>��חGRq�n4�B�9��ժ�V|�@���+�t##L��2��ˀ��u�+B���
�Iz)M���K��i�P�;<�	�s,�%�����M��~i�\a_�.[f�N���V:��l�B3쎕y�vw�Y��N�ڽ[^�z�%u�8����zY��[�V-�[�P�i�Q\t��J76�,5�-b=������i������W�[b>XkS���^���/h:q>��!�]��`:xv��#��e&y�.X��5���v��=!�;��2����B�X�,���Vs��l��i �\n���W�U�Vv9K����W���,�^�K���Ivpja��'cr�䖈�� �c����y����#f�q�5��]�{��[cK��x��2����o��(�W_"�AD^�ƕv{URw�������F�}Զ6�z�]��JjRY���{wy��VA+��O����כ[�ln¼�2�Օ����#�\���*�~�$�b��OQ����k������w�X��WZCM�deV(�ǩ��������F�D��h��tsZ��l�8;�Ň�g�&�.+ju(ئ
����;�a'���xSL�t�Ti
s,���{�����/�b	�"V*I��R�U����f�ܹ�SdcME�f*��<�Mv	Z�Gl��1
8\)�_,[Jds��mb��3��"�ҷǓ<�q������-x����տ[��i���.M�Ka�]7�܄a&���� ]�%|Q����O]�+N���|��V'XN�����NQv� ��"�ܤS�GS�͸n�xٱ��|��OR�����&o����<Gm�x�Ȓ��[E����v��k�N�ɽx�ߪ����w�����#�o��"r��s�wj��|��@�ǯb�ݑd�xOJ�b	K!��vSK�7��b�oE�V����]Z٘kw��#w�b�o��n�IՊ}�����z�\�m�aㇼe8xT3�(�cƦS�W)�=�b�7F�	|��3�z��s�e�I8���!Tq=��Ă2�A�N��Er��' �f�vB;�I�^��V�	���_S&�����0yI�:\汁�hF���WOv�k��(��[��1�]1s�W�9S��×��x7]~��3�#��@��Gb��i�ĩ�O�o[�{|�Ʃl`I���tu�po6w�ԝ��SD]ӱ��K�g���^�maſaplj㬼UE�����{�zjr7v��Ψ+��[7}[:��ݹyB'�ҭ��@�j	e��Q���.�u�����V�n�(��cj�ظ��\��)[�-atȻ9�7M�a;[�9=i�ꈌњ�nA��Fu��D1(��Y[�H����
ypoQ�l��	���������8N�>=WB5Vp��p{�V�11���2�b��j�kg�}��U�l ]�5��~]�&m�}f'����A���%�΀����56���m2�9L��Zm����A�f�IWRM�2��@�R�4r��Y�嘃'X��`]�k�&�`U�`��H�.��*|U�&�P�y9���Y��'�ꇖh��]/��e�`���5mJ^*"�]�x���Xz���Eء	;�{`u�V��u��7o�\�U�rU8�f+[�F.˚g��������V2s�w��}���He'Oi��'R�3?��k�v�� ��|�\�0w<�f��+	�fM_��s������k�����U:�f��δR;W�N��p�#��\�]	��L$�ɝg��I�MN
	��90�Ge+�T���t-�m&f��1}7M�<��J����6��M�Ɔ�d�Z���wuj�y����0=��A�+�=Y0�
��� �`�	� �F�Y��~�ϒ{�7�+��GM$�ݹ���HӍ1&tҺom://^�Oz�i����$�yςkp7s�}�kP�3%��B�7r���U㊇ �h"eӺ����K��My<�����D��9t𛚾�ݱG_sν�D���L9{N�9�
�5��v���"��X��!v�$p_F���bۧ��4����3/8�}.��R"�\�ݢ0jS2Kn��D��}ZTF��֗maŹ?Z]K�'V�y���j��i�ޠQ��ؙ��x�f�Z�VDVV� ��UMR�g�fT;�X�q8��.#W �����w`�ֶ���nV�.M���;1�/�fKX]��m���#H:�t�m5��0��	��~�w3���I'<ܵ�撤���a�`��,�sx���3��8%aX8��b�y�6afQ�{�e3�WR��,��%���}���=�oLl�*�w�t�S��b�Y�U=�b�4����bڵH�%���gdJq�������_F�Wig��^*�t�B��5��"����F��nJl�H�l��ݝ��k���t�� ܦ�N�Cv�tp_Δ�&G����Xֳyd�\R�2�̠�|��ڶlJ�ws�i���T��K<+�?�u�s7*uI��fp�H5�&�A��[,�iO2u�Tj�_j�A�;���k�r�.t���t�}�L�[�;n�ՅU*���\�t���u�{��S:j'-7�us-�����y�z��z/αҙ򿴎�B���wk9&�����~�Y�R{+4������!����*:mJ�T��Q�9UWvY#�DAvԗ���z�UDbN&�ls�5�����t:s̙U�0>y�r-���twek������뎦���Qw*yK���Ė�m�7~f ���n�{�3���=�#��&�a1yuw[�������#���u���<�X�ݿK5��V^6l��|W���z��9OT�{e�4��>�w��#2���,L\�H%���&G_V�K`ޡ8Y�K,)x�����k�����5T����pq,��"y�:v(�oѬ�Q(�[�i�G7�Z���X��������K�0��w��K�C7�C���9��x���{m�$��(]�n+r){f���r]	a[:�ijk��Q�e���N�N�����̤s��<J�YN����8�⇯�k�H��jԮ�:ڋ�J�cL��U�xoU�M�S�5U�����u:���L�lG|�@D�T�b�*�SY���m>���LW0�fM/���s�9{WF;%ܵ��/
�n���e*�M�}r��؁�//8�&�&X}`6�g�ky��`#���1PұRK�sy��6�sʤm'��Mn%���c�����;e�8BB\,P�X{y��,��WP����T���a��v�Nԧ2י7�|Q-3�����f
���|w�qM,�s{�,ދ��TI��O��T]�3Pz�t�f��n��l$.m�a�=p�>`Q0�9�[�:�u��z�NZnPƏg������ٞ�F�V�ٱΩ!Ws{h���Q,�8�-�XjܑO��R��R{W�[\��]u�{a�$��[k����XM���u��h�3hF��F�Sݗ&��4+����5n���^�B.|��;�'o%Ӻ��w4�I��s��p�3`��ar�3r�
���]�g'-%2�|�Y��Jٖ��]��֩��+��p\\��s��H�KP��a;C����.#)�=E��\�F����U��WsRXݚ����վ2�ja��U�΢�k�Όg{��vXG��b+�U����~���5�����-�&^y�tu�7y9���Lk��26��2��}Q�����b�������$e�UE������<�ܥ����pT�ҍ�J,�+��+�\���jK,6zkO\ĺ���Dʜċ
���_�����	�+(D�lR��Z��p�w�b�&��j��^�*�M3����ߛ]/=f �Ȃ�T�;8�w(hS�fr��_���<�S�ۖ�����osX}a4��+vJ�b	�xj�m�`w��s8�S'o�,��ŵaR{�j���vӶ�;eV�dU/+�pug�o�cC��^���ަ���Ju�n3�z�Nu7���[3���n;J��ڧ�u-x���	
�L�]^{�*i`s��1N�ۮ੘��*�r*��F�;Nx{f���>(tS�L9���Io-�4���Xe{5S|<J�ݿ}��B�kݓ�4J�ck�92�]ۛ�y��<���VR��&"�P����[]�
#�<�8��!�wv,�FL��Ӂ��הr�}�}o��s�=)wG��m�]��U*�B6 t�f��=�C4w�h�3ۗ��4&�UD���N0�:�/!Ъ9J�%J�#��T��5=�V�M�Uv-�*��=2U��e��I8y�x�&0W��6e���̕��Z��}G���.�^?R;Zs|y�IUZaK�lsQ6�`f�z��Є^INi���%��u��s���G_g�m�Z%֭L9���rs����:̧{S�Fiӕ�w]�U�6��|G.���|�fy�5L�"�I0eߨ,��WbQw�s��b����z�-��%ʰ�ܟ�m.��>ys}��b�%O�#(M��q4��v/��J�o��P��Q[���>��۵:�y�bn`����\�,`
�k]�sxH|�N�&Ĭ�ˆ�6��X/a<[���1��O°>�F�9����+i�e���k�嘃zk��ٴ��c��;�Y��sΦ��k<[�<�t��;uk� h��;0��M���2�*܉�6�:j��TE�n��B�)���:ىl(<��S��\��Z�!O�H����}n���i�[
�WU�XƁ�����X73.m�����<6E����c����~�j肯˩!������3��8%aN�@��8�;�fc-�%F�(M�A�!�u)_�YXT�-���t�(�.�.1kU��1'R�Gl�^*�<$A0S4�mZ�tNe%�wM#�K�9��wQ��8�� �_/�B^��p����UWK�q5|���
��6����L�Xz�mݺ�U*�|�@���ޘqQܑ
0��>��!�u�p�ބS%B�O��m��:�V��Y�E�N�O{���Wi�f�ΩO+t��+(���0��N
ON�A�3�����޷9j�s�u�}�b�ڿj��z�%ucq6<���mKjP�j�lb���1Yh�	�K"ٸ�v(���\5m{M���ڣq2�L�l�x*�.�+��u�
~�7}.���K��<��+[�-���cHS�q]��议�#���Fո�γmRy*�m�y[/��]��ύvsU.�H��U������Y�|1�_^�D�Ի������2ź���WƻMNڎI���0&�
[[�X�����p��� �!�V���.1ZA�K�^|S��Ηg9g,u�CGX�����XP�L\�7��+WX7C]�� �EV�L](i�*�4F���S�ڹ2�CGu�:��w�j�����6l+�WY2
<i����l:�!]�H�!5:���k]QX��d9r����t�P�I�������[�}���[#.uN}�0�p�0�q�[�A{5v �^�@u!��U:�`�>1Zy�1�g,g����v�q\H �|���2�EL�v�M9-"�ձn0��|�+���
@���Q�J@*��%��I�!W�7�fؚ�u
Y�Wct:�;SyD�`]�\6��y
lVf,��;����}�xr�w���M6:Ӣ/z�7/�:��-K�g!��uŇx�BvQI�v��D;�- z�H����ɲ]�/*$5�;4����`�(�\w��w��_u�I��-�7�t�U'�K��YǮ�a%���.˛л03�ѻ�٘>����^�JY9W͠�SSW
7�7�����"����A֣�y��,]Ь��*�������o�UYÃƻb��͡�$ی��œH������6unMȑ���R��e��7&1�f���@IN]�.����zm�!cb�ح�7z�	v�5]�����f�UðH�s�����SX������&����J�9	y�h��k���q�3�b�;�E��eGX����Jb�b&�=W�]��):�hE�����ގ+
T�9F�9Lo�1�,ެP���ԫX�`2�)i:�\���ɓE#Bc*wX ������E�}mu�b�hr�w.Mkә�4{L�:�ۤ;���Y�����Ƌ�iG��0�fm��K2���;��B	�F�o|#�#�Ӈa(jw�+�f;�щIo���wv���=�,M�*�gsC/�l��x�EL�S����k�u>"�b�U3s_��
�c�b��ruy]MD��Z�q�[��:���{dͤ�ux�����ĂWc�r���U��hP,4\��2<
�drȁ�{)�4��c쬛�\��oim���9�t��];�G��
�ķ.֗L�,=�a�[�>__q� ���q@7�]��onc7ݹN�"iև�Ԗ��gj&���:=*2�\�����̥�uwp}�wmO���F�m�����
�ճ"�yx��S��xqu5C��ΝQ�M��u�iXM�u	1�l��P}�k�A�y���$(У����3m�=Ǥ�1�@��3���:y���Y��nu����1��1�İWA)��w]�����r��S5p����X�"���:��3 m��:�����n�?���}S��B%R�B�(�(ZR�hi�hJ� �hJP�JZ�*�h(P�J))�(R� )�i�������(��
���JR�((��Dh)��
F�����(
R�
D���hU���JX�i
 "(H�(�"�
h(�eﾗ�z{{��]g��y�)^r);iv�� %)�E�����V2�ҖA��Ȱd�H�v�k7+,�Z=����|��z��זu���G<��xS���I�Rf#3��^��~�|F2*JA���ޭ�m��HM�,���&^3O���6���="t�J����D�K�﷥�{kԢ�\�'
1~��
^.)�8^�kh��\�w]����׌���/-.�o�5�~�@�[�-�����"DB���ՑC�RD�\mI)4�K�f ׄ�#�T�t�V�����M��{"M̜��E�K��	.�g%i�vQb	�>ʺ�fY\�U�M��.����W�ʊ����0���_�O�J��;eZ1
���&Heq�"oU������L_N�Y�aR{�k�;�i�1��N���׊�<�'D�Ʌ���b��vs��>�u�XT��Z�j}���u;SiԵ���f�ٺ�1g:6�u��6� ϣ;ݥ����w��qz��ذ}�7ʽ��~���!�_�����}�4�S��rL^p��tW��Fs�Z�-O�%g�qۚ��(f���b���i��o)�v���I�6��нD���F2��o���Ռ�kI
�uH�,δv�Z�y���B�EO���	نI�A�"�7]^)/��F:���\�kHRÞ�_��~U��Cf��n����B����M�6w�a��9�\�9zx$8�G?8(#�-V:1���m3�z�����tFZ�<�!c,2�I�~��M��<������rE26�Q��R{V��t86ɍ�Ɍ��eRT�0
�x9��Xua6'�[�`�bF������N�o�|���bT��|��{x�q�ژr���vy����g��ܡz�6�9�٥��V�<�bWX����O�o�T�|�4��������̎����Ui��aln��T=w���\�$�/Qc�����hԬ��sop�,s{��kU�͞��ݿJʉ�t�exj��춢����^i�+_Sb���)3�[���Xֺ�^A7+(D�oԂ=�"�����t�c���Z�$��(3�[��i��}������x,�g �<����= ^��U��]�k�����
������]��2��Vd���yD�Sz�R���i���է���uʒqs�9N�FN�t=^�렓�����CM�M{"!����4:��Z����yD����IS���o2>�\��8�ma	_ksG[�������b�Ի(�|*��)��o0>��=�Wܹg��g�;@��"�1�3������]JwRJ�,[V'���<�[�:�6�莸5K���Y��՛%�{�p�LT4��m���R�>S�����L�Tz?h�n8ճ��aݻ�`R���P��!b93Y�]G{�*i	)���F��rnQWGSn����1o��:�:�;~�C}���\�{X�zԉ��d�N��h��G�.��Z��8;���T���F�uץs��5*z𖶸����M��m:�e�H�ZI��Cc�)�A1��s�2�V`;3
z�o�{���~���VW{V׏=xWW��6��M�Y�c��9u�|�d�1�~��~��b���[B��g�w�50�޿,������b�GB����y������r����k��Y�Ҟu�_��)���e�{�v�v7�N��B[�f�W����f�Y�.]�X���W�֞�1�9�\cO+���%ޥ�۞���<���&ҥ�4r�Ks�{N��LE �(�Jdz��I]��-��bWu����\�]��nN:ti*��;���C_���Y�=��b��;>q�,�t��ި/g��uM����֮�}LZ���IQ�yE绤����M:��Z��Wr�ݰ%e����9Q^�-a�7�����o�QrZ�1Sm:���zl>]'/ �����:{�=jo�kb�57<�F�=��(�-���k�s�VMu�q9X�Sѕ�ԮHY���H�z�Ğڕ˥#�g�C{��g�J���bۗXm�B+3�5�R���a#zxL"��+�ebʚKy�a���E���W0��zӹ��Mt,l��ax���iX%<X��.;o�����u����u��եlj��1�|�κ���ix��B^��WJvk���*'�=-JE����I;ϵ3�o\�VT��נpڶ��SԶ��"]q�b�[����id"�+�)%訅6��SQ�
���s}f+�����X��\+�;�HN�3X��Wps~.e�;*��\���ni���{5��t́�^t�:�۶�r�-Jyi��wa��:pp���_��Ng>!Q�%��֪�:� 3�t9��W֩�c�J�,��v���](�Z�>�δ��`Bsjr�M
gFPJ�2���ճ�.�8�G�N��m_��@0�.Hm�a���8
���x��=�Js) ý��u�z:�K���V�sՁ%ucq3���s0X���C�֡�8;�M��4S���lGc�Qݕ��a����usi��Q�
g�<��"^����'����6nو5��7U�ݕ��_r���
���y�6�<r�}]�x�ǵR�c�Eٕ٢o;���6�X�fA�2�q!�X�:�>��4V>Xj��O��[���o^mj��\�\��C������4�!'b���)865(��e�T�OI����0*�斩��p�s��r���/#�����R�� ͈��F�@�[��kUL\_n��YJjV7���Wr��>b��r���ѽ�o@��4�r+��xe�4���+M�G�Q�1�|�I6*�Upm�G_X�[صǬnM*P�[�异�+TA��Ƹ��d�< G�>��z��&��u���X�5���̨���7�����Y� V�)gy��t���g��h*�� [��> K�s9r��ݝ[ܦ+��Є�D�3��t�G�.��b���6�K}}���:����0�氺�i�+l�l�b	�"����x��J�d�Ս���q��T���v���1����햼U����r�{wz62��h�����P�4p:���L-g���E�s�N��T)ѵ^浠ޗ�j빦;˽�&*����ޅ`��9�o\��S�Νp��Fm4�������Z���:�?k��w�G�K�[x9�v����α��#C��6ܽ�ꭾAy�Q�V�}6��4��C�N�gjƭɎ���R�b�\���zU�IĔ����1b�X��l؎����9�;�OM�/M��3�����ǀ�ukXu`&���[~�4S1��qD�����u�>�O{A�'���ݼX}��sa���yV&����*,��R�^}n���괼G�yZԝ�r3+!�x�:5;����U7vU'VG��9��qM��J�OZ3b]N뫷(��dG�]�h���_T�e�wN	�O'�[�c����$!�vE:�r��ͼ&.9���]݋�1�p�prf�.�J�����pVV)qN��x�e2��j-�[��\-���zl��@�y�����\3ն.�J��q	뎗P����ճ=N�����<��N���p�9M�2��d�j��N��oP3�S��{�V�<N-�������O5��Xֺ�^A6%eD�
�yW�!䝨6-@˽�ǯB�6�
�dju�u�4�;/�V�k�ш<%���U�ӎ��P���WL���S��S/RX#�����k�4�aC���>�$d PQ��#��@�rj��N�I/<�mXT��C]����9UTd�������^�t�ɢ������	
�4��+o���*D��we��̔6c32���8��N�
�U��]�x�p��3Ai��䯤gi�w4D��5��)��������M�ۻuaUJ�P��=��\�8�/�F�Od;��.ҍ��c��[�a����x('n�˭aM���z��2��F�0�;}�CD�W��af:E��MY�z.�"�c�d���4'Q���%g
5�����l<^kӯڍ��!�g��ui�/�)7U�v�C�bJ�R�2hNQ�N��ss��q�V����oz��{[�'�x�|��Ἵ��i�W�[Z�Le�Z��������]�˰7VNls��r��ԉ���*W�U]H^��]g�D���d����=y������6��Ma�9�o�6���jI/��5�@~���Dn)[�������K��Z2��([�&�q�{�=�o�yc�ꅺ���Ok�w�O[��-�{�����~>�S��3�eM�g�۽�J�����v��w�j|�V��8{���6ÿ,+����	S�h��S׀']ڱ�y�ض7nVP�P��L���!��L�|����V�VoP�af.K,b��u{��=(?V���� ʳ.���L+Tg�K-��<���Q�m3��P:�u��X�rV��=�K=8����&���\��A�,�IV*Y�R_�RY�c�oq�eF�ʐ��3��mu�/�)Ξ,	X�Ӱ��S�eL%ީe`YS^Kh<{�k�cr��(����ёy`���$���8�%ꆛkcd���o�v+�0�׎h쩨2A���eU��Ʃ�3١e���w��ak���D����,2n]�b�)t�mX�`�jTn�m�ԗJ��R�J�9�!����αF&բ5i�Ӭi�;ꮐ�֕�/[���x���xCJ�INp�a�Q���Ar��)�z���-k�1���v�y/��U#�H80�������EcY��ڞ��b:��M,w�jg�޹��u~
�U��c,%'b�Z��v��'�WI��d�B�N��!��oE��]X�0���fc�o#�e�aL#��>U~��V53����!��Gm������v]��q��V=�r�=�C=��R�Zw֫3��ܕ)NF;�����fFU'zXB�tN��)��cE����n;�ݱK]_�l��ŪF�[f���&J���ÛP�nsG1�v�5��F��Otk�s/�����&��,d�S��Z�i�\�<��u��u@'yK<�F��"�n�3�md��=��]ʎ�]������B��3+!$���>;�}��y����ʁzeٓ�^�w��z�[Q�Ӗt�f�:@��%g<~w����}q�.0���9)`�5�Ӳ�*�h�-�V�w0����K�5qU��J�JN�C}a�C�b���КčnW�b�<�ǵi�����)�.�v!I�*.���#I�Y[b���h:�\�X�*zΧ��D���آ�4���Ӵ	\�(������YQ<n��6#X6#P%�ēz6���IFT�$Z���-W�ˤш=(�O)�e��jĜ&p�.&��r�5d<�)��!M3G�e���Wz��9[	5�Y�e�ZP�=l�:�)�3nxk�&�d�oe�}�r�9M{��j�����!;px_m��V,[V�=�5�ƛzgm;o#�\t'p¼�F�/}8�� �k ��u�X�NB�{S�z�mPקc�]�N�ɬNܝږ9ԫ^J�t�HW�kY��z���9ͻt���<+.vb���.�a.�`*�V��X5ߠt�	��]���x�B��'br0��ebȕ���7��P^A\��T�Dtښ�!���Υ����]�*ً�D��]���=��K���}�&�+����jc����.kz�C��kM��xv*��-�����%�Ʋ�^2Dֱ�����*wϔ����U�^�f�Vlr�ˮ���i[/�f��ʀ���k�Z2���w}�َ�j�2R�j�-�{���sr����go�9��:6��"�I�a[��w]�R���d'Jղ%R�T�����kT4��W�taxS�/X�&���7��u���Oi��0���63V�ҩ�<]y�)�@�T%�ǽ[�^���u�Q�OR0��`�e�%��rkX}=w녀�p���)I�nL���/�C�S�z(Uhȅ�c�����i�*n���y�uƺ�j��;f��������(Պ+8�q:��Q�p	`�dy�e���ʼ��0U�y(�x5E2	,�k�$���:�l�es�ƻ�*	.���և��c-]��1��hI�&]
DV��ۀJ��v�6Cd-�Gy��9�T�ymmdɗ%IB17a��C��>�dQ��ĠDӐ���r�[9�`G�A�D�T�+�t*S,����aV��P)�jP+�2�\6v�YݺA��N��V�⑒O	���5�y� ������i:{�"�em�z���iT2��?��p�q�sM_G���N��z�p���u�w{X��g/MԋP�;�w]A}4Zd�Kzk�y0^�B��cEp�U,V3��������V3�Xr�V񣡲�/�C���u�9�>��Չ�=���u+QL]M��x���\]�g���̀��gQ�6W*�;=ڗ��Skm�����S�la���Ջ�7|��%'�:��B��-u3s��yJk��C5�Akq*o1�zX9.v��Iɕ�g��$�����l*��.����a��P9�n��=�G6�R���%wC*;r�"�jz���2��VG`�|{1[��V4]�Q��ytI�}X�הv$c	����x-��0��l/�Vz+�gC�a��X�P��ћ,�
��c�a��*!��]��0�-�g>�z*�Q�t6��v���*�՘�j�8VR]qc+t�{xXͣ��˯�ڧ,LJ�����#[%Ky�[�nY��*�e,]�#Q�1+n������k�J8��@t7�����'X�>3{5v�@j�r"�)GdƎ��8M]��FP�FZ�>�ҵ����ݾ��|l��+0c�B���v�@ΝC;�apjO �w���V��b��-f���wjmc�����E$�����Ӣ���\QT�,}j�����`m軴@�&�D��:m)*ﺡEh��.-oU��	��],"�˲�M���=z���eve9 n�Cln��$g<�Aw|5n�A���X/���2�������A�i�uc3�a��y��>�gXu�h*Ю�����]�Zf͋.Wu%s�˩]�2l��tt��h���W�3�oWq�%�y�����;���Q�������{��gz�����!h�B�i�(Q))
B�
Z
��J ���R�hJ((% 
E�ɡ$L�2V�2�S �22J2�ʐ��$Jr
ZZW!C!��2%(Zh)R���(Q�3[��;����{��z���#1���m�՝�T�;6�R���:�[͗����;�
��k�A�}�ʹ������_Z@qHt�ԯ_�7VI��ls�B��P��93���d!-�Kō{��赽��ʱ�;Z�O^<%�XZë�lOYu�9Ҭ���nV�(7z�[��=��y����Rݕ�x[W��=Ɵ`�ÛmW7;U1�C���²Y�vN\��mFq��V3cԶ7S�{|����j�/jc7zYSx�T�F���N��������cv�=WY[b��cP�u�<�,a����䱳؃�2�os�O�g�ln�=9�����W���48����텹�E���E��8��cz�k�� �VP��$����bkZ\��ٳ4�덦r5�:����g��%a��K�f �z֊2ka�l�d,��X�j�TJ�����>��k�OJ�+��uoV�p�r�`�I��)Kb��eL%�$�X��R{��k�ϡ�
(��vQ�5o(*�b��%V�-��CV�=C�'���#z�.c\�Ui�sL�����D[+.r��{�'mx#��<�T�|�5՝�`���n�zjSK-��sS*�;�E-��1�Ru�gm
=�E���4)ֹ�����84���Z�����;k�Tw�+�[c����&+�Fv��.oqB+I����\�I̾^*���BB��5���\)�q��&�i��A\�Sk�5��a7��ҙ���#��/��F8�t�Wc���x{�=�a"�9fz�`����VS�3�㙻]�h͵��&�rtԧ���#�;���;�a(�£ܢ�-eߒ��2M�峊[����:�ڽ[G��I]^&�ls\4i�������['TZiU����U��m��=�g�ڬ��_,��ŀ�}�\��gA�53Gu�a.,Vk�ɼ��[ꅿh���|�S��X�=�������مyI3��ꙞFr�V�T�~�N���.��TMϲ�3rg�g�R��u�L��؟V.Y&�y{�t�y{N7�Ҿ�7M��g�$x��"��Y��a��ګ���d�����N�=�,��$o&MT��	��s�o��dN��|Pz���]�NQ�m�]v\��6�϶�AG�d�WqH'���(������3��L��-�#�Xx㭋��y[��s��;Ss��f�	Ae����;��oK�u�{�͎�[<a«UU�>}qf2�I6)і�L�C��[���Ӣ�z*)��$��Ա�)6�S�x	F�T�;Hau%������,��'۔��sz�a��I-[g�+:v��S�}��J�YJ�T����;ۖ�r����Z���*ޘo�>��J�/[�Gl�^*;�ƈi(�4��;��-}ؐޕ��ժGp%���~z�l;��C�v�UH���1�f��fm�A���Y��e�K�����E���g�v`�Ne6�ych^�,$��龫g:�G���N�.)��r�<�Co^�zu�}�+��C�3��k�F�#)���M{����RKB�ЖP��ˮ�vy���hۋU���3b:�v���ڱ�hw=\�XqT^�!ZrZ�`�٣��h*j��v���oǉa��j̯j�.�!�(>�V^��-Y	Ǹ$�39EG7o'T�:��bo]_5���ct����WDX2��k�k��.��cAucn�x�d\��R���	�����K��s��4z���M�g�k��-���O5�n�_�OI�Lk���.b�e�*j�s	^<ݜ�ÛP��7�j���K��g�%� ʕ�fLV1Wm!�Y��ĩ�[����<M3�s�^�咪��ɮ��'�X��뗋�Vz8���D����[�mc冩lbL����U2�J��F�-�Z��W0�7lO`e�em���z��F,	,��������+��UK6b�Q+��9���.[$��;
��<lW�eF1�5
ț�ܽ�����j�-N��<����tsx�[��h��D�n�*�f�%�i�W�]Չ-ug��b��i�i���������14p�Ub�y{�"�uqשuњ��L�:���3n���4�%cy��a�����Ɓk6x,d�"�N`�l� '�\��9�6��;ne7����V_RM�ۢ*�d�P�.�nb��'�=��qڐ������u+��J��L2/[;{�բ#����b�\Xz.��pȩnꭚ��^I��[m�x�|hfY���g;�ce��|Z��;�d=ZjQ[׫�$��3g3Lu5MnL�p��,&ٝ$#�5�>�^��b�qf�]^_U�D�����'���&Yں�LbÐ�b�������]�y���	
���w�X4�of�e�q�Ɯ��a�t��/�>c��~5؁�3YK�pBjD,�*GO'��0z��m�a�D,�����Y�Du`�Εtȃ�z�vwk�n��������~kh�`$n�$�oɱ� �����'=ɞ��
��*T]��N�*ou��ܢ��枼X.�k�Bu�[�`7Q�ه;;��#sϩO7v�V��K���[Y�̾Z�y3O�Sl=�]�j���b��F	�V��=O��v��Q<���eU.�V��5.���yu#}x�X�۾������.E��b��q�.U��O\]J����u6��(���/ƨ�	������k̠�r��qϬ9���*�t��5��e�|�QAk��
��I:�P�;�K��=�3]�dp�y�1��8����䮺���;����jP<�M���7C�D�aG���/+9M��Z�v�(r5
�g2�N��dHc�q��*ө\��^�a���V7R�,oJ2b�wMΌr�X@gR�9_]R��Jʓ��eq[���_�����M��(��n0�Γ��ؒM�*qX��L�P��[��M3��앆�k��i
���ณW8��TE17��v*Q�
�V��G7���a�M>�t6a
���-t�[W�#w7xҤ���<�`#�xL2�T�b���ժOq�k��Ô����I�/f-a�n��%NI1���{�Ҙ[��H�1cjc�c�ݩ����)��R
s_u�W~�ٛç�!HU�+��E"W��n�b��\�$y-�4����Z!��n3��uj�U��#~����r��~�3kޫ�}�쓕H�w�I�9fx�x('n�yU:�A�r39ɽ�X�P�Mv��!]IN�S;W�N��	#U�'=�j,R��m��w/s��Bq�4.��e��ʗ۹�Oj�i珼���Ôvy���H�u��õv�i^odp�Kj��0gq[����*6w�ص�9Ꝿ�b���=���4_a�hپ�!���fu�uz����j��t���P���C�B|N�6���uf��=�y�[��Jn�{�kbc��f�0 ��e�������,����S���7��Z��&�^��G���^N���Zz��הڝ����\Ν�8���:�N��c&훹�}).u��s��/�Q�!P�h�/S��"ʲ��=��xS�Ͼ�?�����n؟�z7WǓ�ӭ"�I&7��R3JvVF1�O�,5E�������8�r��R�=��9�=
�G�Ki�em�D3z��F.K,g�6�״�}�W�[HFW�y��Z�:�dαy����N��؍�sѨE�V�J)����n�Պo����v]G,��k�%]K6)�JDG7��Vl���9���s�b/`�m&s��f�zv��A��2��+,�$���u�ȗ��m]-%Ҙ3,w2ц�>�����z��ax���٩�;�V_=G�>�o=�/|��Cܽ�-b�`;��˵�b��r�Sf+g9Vҷ�m�db�jj�0�
��W^Mt�Q�J��^Ϳ�L�/+x�ǵ�[<�g�"h[�g/s8�sV��k��ݏt��Yu،*�N���NWkL��%�(�Y���mI�1���&�)x(�U�0�^�X���������}b�-f�P:��i �y���E�s����$t3��{��»����� t�O�W<�B'z���a⁪gw��j�z���='K�V����rzGk� r�R�+u:<aX(���Q���̋����������G*B�:mMi]c����Zu}msљ��Mxv���9�e2�s%]^$�o�69��Xf�eOg��M�}��/[��� ������j�fe���ջ��[q��/p����2k|�5��S4�L���-F����{`k[�kI�qs��^Y*��y�Ȼ�^ <�h�6��y����yix�r����a��U39�Z�1J�5���5Y�)N��3ow��a,����ݹy^�U��ۤ�ߵ	�����fV]��0I��$7:���0^�V�t��9���O�F�H3q��͓�*����cB��ˤo�AeF��$���N��;A���]ɧ�B.$�� �n4����4P����Cn頷�V�NTn�v	�h�f�8Tu������6�r<�jUҨ��ỡ���[]]QT����*5vr�.��7��X�3�<sUj<U;i�vw�5���t��kҍ�W�j֫�O"���Iժ�B��ƪg#��-��i���+M�����c�
4�FȔ�ǻ�y��۞�g:K��r��7���5��O�ұ��*-�|�m�J��q��.�*j^U�;$�Հ�=�5�ƛL��: '�*���b���Sg���Mx���K�Y��.:��H������0f\�ڎ�4�r�(`5ӷJ��N���Yt�_ug���~�y�<(>�D�=RV:���ز�{b�|,:�VT��k�XG{S��w��1��W�;���jk��H��ه���B�A;qaV:1�u�RfLɽJ}7��6�x,�e]?Q�����7VN%65�Z9�X��/%@�6&g'xV�u�bT���^֬�z���&�������`
�eG�~qP�O�)��ۓڌz��<�b,���N���ph�]�,[4���k��o��i�YL	-�蹚��t���&�%|%�����b%�Õ���t�bsH-K�luo��T������Lu�/N��G����Gc�S��PT��A�d�FiD�}~��t�n���[W��8���Ñ���=$������ث��$Γy6وь�u]c7�[z�{r�u�TI>�����+������ͪ�e���I��z�����b�9��+g�ig>*���>Fd�	����^�ד�屻bVW�x���j�<�r��h9��Z�X�@�c,��QG����k������lՇ��n��s2����"yL7�B6m3��P��-�&�t^�+�Gaq�����uOR�w��b�A�,�I_�]RS���r�����z�l��@=��S=�~�k<�}T��l��:Ū�0���T�#ĕPf6��
AH�T�eZ�E)T�x�s�7���!��ͳޛ}�B�q:�buL>�l�p��H�/��@�R9FB�}W++�7`��_���;��8�v��L�=�!�8y��uh�s"Y؅qU��!*��EA֠N�r����TfM��w�mX�f���6t�ZE�a+��Ė�/�(R[W�V��n��lv�GZ�(3�X�*���5_ẗS]±�Yڸ⧨̋`ӏ8I�	M��䠨�#VQ�%+�w[��ק�iR�0(AO�����yot�r�`��;�G��6���1�ϷC�(��^.�mq�]u�,mc���QuȾ\��q��n���@b����wsB�]+���)3��ޮD2hP��٤�7Bsed]�A�m�ǫ�C���W����/���u��Z�N�GHj=J�QA�Z �ݧ�i�{R�ۮ=p�wc�t�9��M���-f�P��]���#V����K�+w�g%���RS���{H���v�V͙������qMO��5;k��݆��������\�n�uN����G�ۮ�T�'|�e`�$�:��K"C�FVV#>�f�ʍQ.Kw�nTo�,�G��qՑ�����5����G�x�`�]��k�(&�*{��3���o��i᫬���[$߬���!��9!����-��yx�{+��yx���h=�];_C�c���|n�s8��˫7t��
���/h��Gr(m�������K(R��h��*&"t^*<��(��3�	%:�'�{{Y��P����)qb��u'C$	V�z��.R�>�}�O�Z�4�ޚj\��J�I]�i��ا+N�h�XYwGٟ-=��9r��3/�^o*ڧ���E�S˝�j|U��8��ǔ�>�t��R�����3!U�K4���Ŋ�z�`|&$�W�%���8�;�3bҥ��;�_4��MPv�+�֯L*r������T��R�e��i�[�D�Ø�t����;�
�u
!$q�Zl�^Xg髂�区��a�ٲ}L��]现��n*3�kU�#]�%��Km�KWm�����pW&n�n�m���ըr}Zܫ��j������������vl�ջiz�S�1��Wr�3��/�,R-ߘxlVk!9F���Ƿ�	Mts�o
ח\��>`��]��nm�:t���^v�ؚ��i(�M�w�a��³"w��@L�{�	�������ڄ��Q}B�,��,�xq����YK�C)��Ju�ٯ\$�K2���
s6hLlTI,6�i��Ҷͺ�c:�_��!ڔ�-oI�Z��[Χ�Mki}��j[�szJ͆�t����]G��vu���K�$X�e�.r�q����V�����U�K$`Ť����W��w-BO`�t�./0IC0M�ܡ,��C��Lb͚Vc7Y#S7�|��;�� fY��-&�إJ����7��T�B�/{9G-2��K)�+w�NeRIg��T�	���{�aJ3�����' Wy��yAbH���	��w����MGS��7���VU��ಌ������u�N?���Ytv�x�hb�<�f��`�P>K�)C@P�@R�-*R9R�NI���dQ�d�fBd�P% 9�)�f
�4R��J�д)HdP�Ae�4�E	"e�CF@Rd�RJR%��ҦBe�a)KNNAI�C�#ﾠ>��Iu3A�xa���X�=��$�,m�{�,䜊2UkHN����o��M0���� 0�j0[�r�E�"��}8,��q���Gfք��F9Ͷ�;��&�\;��by��g4G��B�S�}.��?W��	�>�M�-��(uvm��u0�r��>.q�G�Rv�)��ܽ��FMh�ݪ�G��!�j�Gk�Nي�����5y(:�޲�K��ZJ�/�,y��Vǖ7�z�^M{yi�q�5�끛t��!��;ꊉ[Y��S9Y0�s���]z����C�U5O7���02\o[O{�f����U����am:�7V��iXo3�N�)oa��+��ڹ�[���ޟbt�o.���wCo�L�� �X��d�W^�3pQ̚�=>Ji��GTy̓E�:�^^�/DuM<1�N+���j������a��3X}�����}�>P�M���k=��բ�NQ�q��ˌ��^{�C�y\�T�YL���E���H������8��߶SMQǾ�J��pf��<2�5�Q�� &=��q<���SnVC���".�����bf�|ݰJ�c��9Ntd��X&�ٹ�a˙㔤�2�1���<��8�C��j�|��С]Qy�"�5v����*v������r����b��h�;,�,��t7
�.�l�v���bj���D�RA�Mio>OwOeoh[�J�qR�ޚ�%k�o>6���y�X���^�k8d��HA��]&�S{e��]Հ�q"�����'�?��8���kn�z.x�ƾ��ў�WF_��r+fP^�/ck�?n�Nזvә�jϴ�W��n����1ޕ��g	V��'�g@����I)LT��`�g<�=��f�g^�V�_��>ޤ�>����Q���\-���2�O�����ʌ�d_�j=�P5��c��k�X7옸��ܫS�[
����:ZTk���;��wv�/�,����Ч�9����s�C�́���8��P��w��|�C�9Ͷ7>N�I����p�&��u5^�z=�.z:�ܢ�uMJ(�$�m����]Qپ!�ՠ˞%��c�|���fN�u��|;^�'�'�tڸ�����q�W$�iѿ��9WP����P�-���>��,�7���r�Ix�0W�� ���RwlU^u1t�}6vlTJ��WR��>Ĭ���m�U��W����;��7�\>j��DG��L�܁����t0��^�� ܱ�g��立k�D޺^v���BZ�a�n�q���g_������\�%@��n�eƺf��I��Z�fQ�d���V�p<��:-C7e�n��󞯖7�>}8�����~�]S���i^��:]!��i�٤�.�v/�]��/*�0Ckʮ���e�)���Ѩh�K���]oN��SH��X9������0rb��[Cq�Ch���fw9�������R���p�dd�u�=�u>�yk��}�i��u=����w�*��eQ��u�����nfgw頕�+�C����-����^{h�^a*z��帣 >/�����3{�<�{�_��V�^ˡ��N�fax��+�Xn(�O^R Lv.�5��ʁ7��c$^5:�{"*�1��y\;���\=U�{�s�xe���f:\�������n�	����@�:���DN���� >�\ˬ�p�^�}q�׭z�d�$�%�3�R��ޚ�q�J���r�o��ML?��5�i�Tc�	eS>��3��CЧ�}�p��A����e1q[J:|���o ��(\T�B����}�4\B��0y�t�{v�W|Uy�n�^WH��:]�u�=��_9E����p�@E#�3ß�y{)׆�m4{5���c��zMw�=�q}^V']n�xnT�p��ʌ���)Pvy��0��v=��T��5*�.cה�2�˛�s��3x_%����Z4�X�FK�BS��* 54H�0R�
�׆W�^��o��O��9���͌�z�Yԯ��\�O�\����re2uү_�7f�4���Y�Ɉ�E��@�n�Z�&�{�%,�F���"V���u1�s,9�sy����g6J���uÝ2��el��Hʎ.��*ʳ��<�ȓ@c|��6�;}����Z��ϴ�r�`6۽��5�*���I+� 3`'\+҄�T�QP���p�=�9�e�����Y��Z]nM�ܾ%�|\�%�*�	�2F*�:7�$.�{*�BR�r�>��x��]/\d�5��p�]ф��'�9p5��ȭt,��Vm�e��z`�گ*��;���IL\�u����x=J^��Pʎۿ=���_�Si�u���$n'3`��ϺF���FT
�7���J�0���w���xn�y~�7�^;�3�o�*��,:�Y�;^�s#�X�/z�:��SCm�g�{Ϩ���>��s*�z����'����Z?9�Kss�uWoC�zO�*c���+�?�;?�-x��a��UC�;�պ����gq��j�����6[.���p��d})ֳ��yq������d��А'�g�We!����^?���{���Zp\S��o�b�������2���7��#�Uqw��xڼ�gv�|��gk�o\������S+��NB=q�ɠ���؋�+Н&y��yGIᢼ��K�ʔ)�W�ݛڕ� ��΅jQޤ�N�V�6��Y��Y��/-�Kw��f&�f�&�m_BWV��0�r�����7�JY�e���3+{��^��;DRPC�Q 0v�kT���5{�9Ԅ��r\0&(M�����Q����O�H���S�Y�O���RS=�ꥎ^�^�/n�==�ͧ�d�S'������&���q����ft;�P��9�*f]��%�B��)��xs>^YqJ��7�iN�WW��9w[��zf��>�R�=��y�#�a����H�ԝ`%P*��A�3�tk�ѹ��y�y�����ˊ�t���L�=�>nNx�G�M#K�ꄳp��(�5U�T�q��*hVw��إ���9�(W�����ԺH���m�C9�w�m�N_��١j��5�s��:��{�O����Gy�L�愣��`;�h����C�_Yg�\�%x:�DOk¡�}�(��vd��VB����<m=frDwJa�����2��bs��U��B��BJY/��FM9�J�X�oFk�7\#q�*G�|׭ɾ2K�6�
����S9WP��k�cv�jr�/l��d=Gg^Qq��6��4����.CU���M��S��QX^�끊cn�
�����m-/���uX{���yt�ju#9ȹ�{$,�X끓�;���9wW�'ڻ��ع��~p ,�GƯeT� ��К[��k��[q٪�aɡ����%�M,�S��(�%��J>]9��wo�a�r�1i���R�]Xd��Z]5�0�Ev^udl�a����$7��vԕӫ>Ҥy`e��]�s�-�M�E��%�Ql�EU���<�yԽ'���Qy{p�SOrq:���1[������|�a�~rNN~͟��@�==�.�J��|:(�N*}G�d��6���\�ʝ�>����w�c�x�[!Ы��v�����|�G	�6�%�B��Xn)H����W���|��*�ܥx����ͬOv�<s}�ƹKiG̳��rve(��vh�x)�q��H�&C�oOg��y�ӆk�Z:/ܵlӵH5�w��*���ۡދ�$񨒸���F_
#;�޸_R��n�������i|=����Yy�{p�K�,iWZ;�<��$�L��B��}�Q"�ͨ��G���o���ɟݕ1�*v��/M3W��>��YZ}d���θ[��q��Q�P@���ނC����<(?e��r���*|�����n}��*W���k�k���!㸜�wv�,�"��m��s�@ϲ;6g��}�@�� i��P��w��-R
���Bu�N���vIp��+�=��q8\+���ښ�x�H9�>�+K�
Z�3������|AD}���L�M�����Y��N�l,�ʠalRR�DTp'���<��=��n�N�6�i��	yݖ�ٿ]
/�I���X,yl�W���{�-���̭��ͭT�l��J�6���s�u�h���i��Y��&��j!L���s ��HD%x$��G��g�=sw���~���q�D���`���Jf]Nq�W�|VӣqEiʼ�L�MY��V����/�:����8��ɿ�u��r��*�	ݰTͺ�Ϻd����ب�����ϵRʞ|6}��S�>�ᕆ����wu���-�&�7@k���\k��s���c����.)�NY����6�`N"�0���B�2^ο\/w;�1�N)ɷ���t2�]3enF.vx���m_��'� �U̥[�~5/�8N\d�u���C�����Z�s�D=�f��K�w���>�$@��]ݽ]=G��n�� %�e~���x�j��\R�.#) &+�m�U�O�gy����>w��M\�s��#3�_������%q�n��WYg��;og�]Z���ؑ���}��^���C��\�S,y��'�ù��s�['��ω�2�j ��t��9�x��󸐍֫�w����.Jq:����s.��w	��=��Y�-��*7Lʙp��m�n
DΝ�?>�:�[���r9J�,��|�ܲ�S:����*��#�e9�8 ����ǝ�'ƵS	YE]]1r�խY^�n�7^w�:��H��K*�H����I��ԇA��1�����g"N2*�#|��"��Q�痜�+GQ��7B�V�������Zm��-]X�7��:�K���t[F���/c	Ь2�;Y��i��(�[K{:��
�E`
��?�kυ�K�>�頪ֿ1�σ�3ю�;i����`z&jJ�Nk�a�~�=9�h�0�M��J��΁��H�T�~^^�B�'x<��G� �c�-K!�������c����'�V��nT�h���"����_J����w���-����'z�(��4�Rgs�N�i6�Ԍ�whJs2� �D�3�J�F���w��Lͱf�{U��8���b��:H�3�-�s���n�3l�*����uI]6H�H��O�eLy��S�o@��+⧸��|�_vh�W	u�7��Y�s����T'V�
n]kݷ�:�8��o�w�Q��A�*S4.)Oa��Xj7]�!.���Iْ�p1�U{u뫼�c�u����@q�Y'��_�w�+�}��ԥᫌ�2���C����_���}�������`O?����C?uďJW�PY��>�a�2���C�~��Z�8�W�W��.��ϧa����U�[>�憵~����j¿����b��&�0�C����g��c����܍�(j D熌C�+;i�;1�q�.��N�`��)�f,�W^rv6,ͥ�J-�kL��8�%�{�\���R�����o�*�Xy.v[�<�q����p��PL�P�{��q�2�^��_Z0�ֺE�}����2��Ls>��LV�1�\7��9���p�̯��4<�F�a�M_�loh��X_�V�������U5́�N���O.7�^�P�^L���8p��㼷����8YK�_u���N��]�.�����u��R���\n�^Fa�:���������4,��e�@:P�_�!��d�}�� ��]�^��3�Oc�غ��Uޝ�h�?C�ч�m�>��z��>4g����3%�[�/]�kwඪ{0�xxP�5r�3���>�^�S�� �Ӵ�B�Ws(���d �c�����϶}ӹ�c�jq���]\�rR�	v�R�}8���C��G��a1��U)�:������#r���{Z��qFx�>�<��T���|�a��:��wV�'2%�PG��wE�>�>Fn���ts?�z����鯻6�/*v��D9Ͷ�;���'����:��wU?q�K�;$��$�y�п�N���Ͳ�˭�=_Yg��"S��8:�^s��F���w�b�N���R��&e7���<ޜݚU��,�C{�R�j����c�����0gmbrq�U�
/�{�l�7���2���& �����Pީj�<;�vޝ�ѭ�:&���}��ZxR�[n�Q����ښ��K�R|W7����`�9��{���{�\U��ңĐ�~�b�m:7Wd�f�.]w ֖9EM���1�"�saEu�N0����z�S^�&��/�����[Y��QL�\eB��cׯ�����Z�Rwm�qʮ����H)�����J��v���>��Ǘ�z_t*���V���MYl���\?w;�>��&�]1Z�H�j��n��x����+�bMz~Uni��}�{fׂEm`˩xN��ۅ��xcܜW3�LV��<u��3X1�ڎi��"�p���ӈ�c+ᓃd�N���r�P�oUr�*w��9�{��LϮ�V'��o������~K�t���s,�?W�_.+�Xn)H�)1�W���y��
��Ei���鞜�����k�V�)M]xn�BYJ0|Y�S��ٔ�h=��A��8-�C끕A�}~�c�Rv�ev��uMyyӼ��[�����W����ۡދ�$񯤮 ���Q�ƞV��]X��}�v�����.1U1��j���{%��{p�O�ڦ;�+��z4���$�L˾���v��Ԫ۹Z�1T[��J^Ȟ�)�d��[ݳD)�J'����/�-`���C3(��,^����}{�i���sF���-����	ZݾWiY�ڷ�æa�3�-(�1Txk	��y��h�n�����O�+̷�%]rj�<�nXƀ+{xR��]k��֕3rK�pw�N_&v'`����k�7��Q�&s)Ɓ���c�}��!:����S!���V��!�&9l똮pm[��F��[����^c	���f��4��e���M���L&������8k�E����@80��t%N�,�k�܎r���|�U!9)R7w��ܒ�-,�c��t��S�X���}a�Z ���R7�Q�5ϱks.ã�u�Gl�[�D<u����*Ŏ5�*�;�(�;��ͮ�#e���������|̟m�#�m}�yD�w&�u�@R)|%
��%%2�t�u�+��0�ͧ}�˳�n`�3��L7�`�Xj;�������=�2=@vP�ʷ�d���i(����م��b1!� 3��ۏ+qkO*�_i����ݛ]���L�S��osv�i%��Z�Y�E��kf�s�3��i©f���Ѱ�G��0v��_�2Y�l�@�*Ȍ�dR�VJ��=2��RY�10e��e2���zȶ�>�/�7��F�)*3¦(��:�ľ�c����	+�Ճ���M}v�"�p����[0�8�
w��h�!w"zt�� �;������%#bT&@�	�#��j� �v���;/�T��
cN�M|���wv<��h|b�k,�)��ͭܗύ�/�V��!na��FX�{��s��a��:��ͫ��f�rN�@����7�f���,�sF�^n�VN25��ˣc6z�� �vԦ�-��Wˮn�lBъ:\����$���#�{D����I�u���bO��:�p�l��������{�x�Ǎ,�'@!�$
|��uc��/G�\�DX�fVj(�s_ư÷�b��+:�vTgL�V��5 9�"�*U-f-�ˎ����>=�F�,s��j���s	Z�҇sn_a��i�kQ�el�f�cpp�:�N����'��'sk�V��Ͳ�vQ���SozE}ٚ;zM��A3�5NU�����F��)��;_w7[��ň�.�P�#ZT�t�<�6��:t)���eѷb&����,�w'rR�E��Ĺ�F�@���Q�z�L��K8kTv9:�lP��q�L��b��Ӂȹ�TE�6ԗ]X
Q��8�g+�yF�+�vpۘ�����T�Y�Z��M/{�. �� @`�3f�RJ	kΚ3Q���%��&�Ax�%󘫴�S	�[+�����B:���&��3n^]r}h��Z� ��i��;|3kt�s-̮���� ��ә�񙮢y���	aX�	��%�cx�.Kswy��ii�%(�t�Hn��o��\]^���@Ԡ3d�)�t��w��c�����=1��B���Jr*## �0�h���\�$�
%�Ȫ��)j�rʩ��������3�F ))��r@�r�&�(�r��A��(r�2hJ �����"2D�Ţ,�&
F̪s1p���)�L�Zl��)20�h���ʖ��D���2�Ɨ*����!������h���'$�0�����	��d��r,﮻3���/w�Lk:�ԱR��u\-�^ԝ�I�9<�/"WcZ����'�j3�EvA[Pۛr4w+6�'�,F��ۭ�s�x����3�1u.�B��5�S�zK=�����ꅜ]c/�6pJ2c_ 7'Ң��;��z����\Ә��g��D/*�V�_K]�9�a��㸜��E$.f�Ϝ�U��S7�h�8*Y��`�� �@y���
_v;�ǝ5h3�2���������yw؏�Kkn'
�u����"���ζ��Z^xL.��7� �5��f,��נb���>ƃ�t�^p"[s�5ן��̺������4��+iѿ��9J�B�ğ	��O��Η��5��q��G%���6�p�1�^��`��u1��%���f�ϔ�*�j}u�77{�a��N*V���|r7^\?}	+�7�)�&�t�|�P��##�x:S�X��0ڊ�|wC���htq��"����+
��U�.��w|c�bqNM��vۺ����~�W���c�p����za������(�>�����]�!��}���C���Cɞ���ڬ��������g<��^Ώ�s/�0�a�7/��}�@綅A��o�Qh����t��b��I���7������-b��i�]�?���l��3�3%�G�r�Z�m����Q��
�1��ؒ�΄�nQWJ�����.�>��+�v���G_�I�%���/%�0���8t�q��eWj��V��x�Q����m}Z�a�NF����C�
p��aY��
�+�Xn"�d��z���<w��L��f�\ ~Ol��Ȕ*�1��y\;���J��z�]TVO�z�+]r��Tk��2��]\jah��T]@zl�tGr�e�[�L�]Q�ֳ�\=U�xWOO����J�����̞5�R6	��JS�oK[4���5�
���G�ܦ{�E5p��Vq<8���!��r�Uo�\_I����OW��|�н4\B��0zHf9�qS�Z�g�w^��}#���s�=^F�nT�p�UA�q"�.R73ß���P�I��*f��+2E+À�z~��'�a~���lqY\'�v���,�B"*3`�@T�g��ai�Tq�!��T��M#�oc�q�׸z�>;��&�:������:�sh���F��)T���S���M�n!9��_x�A�E�f��|��}�}���C���mށq����B��(\uI]3��:.:�w��o��w�
6�I�|<�F��EB��ܛ���,���/�W�����"���I���Y���>{=�U�_��1�o ��<�vn=����c{�,VWH�.���7=l��@�� �E���/�
��O�3ߟ]gY99䠅��v�-�yB;@�t,vp���ق�w9-Ν0G�K����`	
�K\I���n�X����Ʒ}���T[�!u��.uN{^J�Q��iu�I:2y9p5���̸l�cZ�
�Y�%���T��W�l��ͷ�z�E_�U�i���0]?/�\��Wm߂Ϊ��52Y�ݏ<���9W簢�ɗ�,	ۄ���\e@}u2{ \��9�Ӭ�qEa{��CR>)��)�{egm�{ӗOC���i��3*!�XU�ّ�{=#�}D��|��T)��7s��ꢟ/]�w�ѽS$�ሸ�^������9SϟU1[��7s�>Ϻp9D����Ӈ�Ҽ�5�->�V��U���̞7�{\2��-p�\os�q�ϲgG��Pu��̪oQf�?�|=Qe��tp_Ԥ>��(�U����T�2�!߮7s4dC�,�"=>�j�o;�#�ۦ}|Ou�C� Δ/�|n��z�d�}�� ��]�W���x���4,Ϡz�3���
j�q殸-�U�1p�ۖ}g�=_�ƌ�!u3�fK��렂��P�����u^��nnә��a�	l��o�N�z|���z o�Q�x���1�&�qFR"��	���J�q����^�+&(�ŋ�G Z��nf��Ѕ0�)]�S֒�K7�uu��M����9I�<����'A��M+i����3���
��G�J�kw�O:��
�d����*<Ҭ޻S}ѣek틟)�l����P��K��5��}�y2��O_�3oz+���ި�J�CRZ���!�y�#��wl8��+aH�ԝa�ކ��"�,W���;��@c��7�e��y��)U�yL�=����:��wV�ZuBY�>�_`��������w��>s l����xV���fօ�;Hǜ��G ��&�w���÷'�6v%�eB�x��U(ک#�ā�9t��)�s���ٶB����r��:��r�K x��	�t�cxf��u�5�K��*�M:72B��b��[N��]�XP}�D!�ǬJ�=�з����R���_���	ǮC^�&㌒�������}E3�t'Et�؁�%���]t���S�c�sUto��m;`i~�f������`6���A}����c�}�D�D�23az^�����s���:ɷ�LV�R3a�>����x���Զ�P��է7����lY����1�/	�q������]&_�o'���{T�o����9�
������g�/�q̓���{��	r�W�O���N\d�+�n��^��T�Y8���Н���Z��G���7Z�|��>�e�\��߮���_�T=��v�?[��kh�]�7��E:�m�������p���_��h�3�:]k��T)6��՗�3l�T�fP��b���xc�|��]5�e������٩�Cx�>��^����1G�����@$�^T?p��՚�x]���@L{��#.c}�ێ�����y�9A�{�
���.lf�t,kn��ω�0�j�B�3�"���U��͠���묧����"u����ا��Qn�k�;�qW\��x�ą��z��d���7�g=��ʝsFG�j/���聮�����Yy�	��ڦ8����y�J&ed�o�����}�.������1WP��Nb�Ur>��k����K+O��G^uB��̬��2����O3]��_�(޷�t�P@�_�$9�h���L�s��X*�+��k��5��ۄt�u���k�>��}^��:�ю�YRʀ-2�@)(���@(mDv;�ǝ5h)���D����ɧ�{��w<�;���D���QN!Tԣq�@]_	D�u�n(�/<&G7ױ��/3���V���n2kZ�sĵ�s�p۬�y�*�UT�o����#L�Vӣx8=�������O�Lr-o
�|�ܛ��p/�� k�^:�
��S�%���6�'3M';F/�oB2�&	CD�54���Q;9d�[}xL݈�}������d���e���Eߕh���k��Ǡ���E��$�oeDx���C����l�u���׽x-�Zj� L,Y�	e� ��h��+i�ۃ�u��8�����Y�1��'#���W
�������ח�+�>E2d��M��t0��R��T^��O��b:�*R���6EOa�qK)�����:�p�����'��9}~�
:�T�`:����!�����aPϷ�'���.��b���(�>���#=w������n�@^���Us33�7��B�^��5��1\V��O�u��}$�˃0��Na�u�p�;��|�d�7_��ؕ�Xb�=^����fUx	S�>��A�N�����S��Y�^5�B��UaLk�ڟ/a���x��n�%G9�m�0�wY<�ULc��O+�{�_�rOt\�ʎ�T�`���Y��;���'�+Cx��N�U�����p:1Hʹ�Y�+�O�3|���rO��0ќ�\�x>U:�e�u����L�rJ錈�#���f�^�B�rˣ��3ފj��S\j*���|I{mj������G�_I�� �(_�=\.�_)�/MV����|!��Bvj*�7"te�w9��8�N�hSl���(�#ĕFt	�{�\�n*g�?//`�=5��q�@l*����%����:����wR�N��y�eL�&����6��.u��+\���,�����G	�P&^A=$�R��qdn;,Vkz���fH�R�o=,I�x�������mY!�u�Xɒ����fR�wK�͝�G%m�I�]Y����ݜk;o4���{�I�ϵ���+��N���ܩf�9Q��R��g�R���F�ʟj'o_�Q���on*���p��q:���Hˈwv�'3.v 54H���Z�g�z=x+��`������*�&���P��N�>�3�-��;Xn��U�j�UIB��;��Ó��M���)��d��%LU�KӃ &v#�EBK�����,���K�63��F7�]���m��oQ!�z���L��4=.u�N{_�+n�!%�TcRN̕=��޷t��oO�9F����2*P�5�r{��}bw�
����5FJ]�~{'�E���*Q�_��9;����)�E8㟢����*>�̞�0��Na�.s�(�/{�썜/&]g�~]=��+���UON'!�P�*�����~�P��Q'(�fL*Z�p���i��8\QzN�g=[HluU-'�r�9�>�b�я}���d��N�:M�Ƕ<�s5ݛ�����s��W���d�*�>�~�3��O*l�|�\o{����a�����&�����)�85���(�H��b�o;n���ÖM!�����C�v�����w_4
)��FU�=��Uݮ�=֊���9��*�v�ޗR֪ҙ�.�:^7�R#*-��0�R��o��Yw(j�"�]m�]�낁[�u�����R�0$�M���c�<K��#�%%�]��My����ʠws�f�S���f�����y�5��a�/~����(������fP�:P������!��Mъ�	��	}��;Tjf����<�S��I�u<qU�1m��g�g��0��҇����uR�,ĜH�~�B��Ϻ}��T﷏h�p�	����-���!������s�tʔo�x�����ty^qSK7���,���ɜ{E�Ύg��.*�+xZ%����zm�T�N���g$�@�>�=��a�#V#'+�|�=uL���ӹ��
��)�g��rp��R=�;�F��]�����G[վ]��bh��0�L��9���V�͝	�֔�;��Þ���
d$��/iE�]c[�?ȶ~���I8�+[h?�"?l���d8�@Cg��Y{�h!j?]�����{M�Kr�E���^~��@���*�Tӣq�$.�;f+�[N���5�S��*�&�w�`�[����F���\$����,~�F��T'�׭ɾ2K�gn����S���)��$ʉ!�wi^���zo��A�ui�́.��B���Y�:d�������Q��R%�4c��Y<��}]�(�I���~�.���-9Z���Iq&QJ�v��H�*O!�tgsb;�}CJZ��1����3S�prnN�r[���i)16�� \���������_���yly%WF�� �:`a}�\>p+�x��
OC�G�W�w�s٬m[��ef��az}�ᯯ/������r��]1[���T}3s�nUS��3����㈃���p2p;��!�/	Ã�߯/n��i�G'���S���	�6K����M�gWG���BS�ư�;ȜY)/��1`��������x����B�OD���/k91���X���`|3�O�O��3�/f�W����(O��@{є����s�����;�[��]U�N�~��[sʝxn�C{\/��폍�6Ot*�e���)�o�����9J�5�{��80&��o��}�뛚�(>uZ��|-5�C�sĞ5%q}.��z��vۊ-��2gV� �]?C�,��ۄ�}�Lv��⇦k�^�7��#���?���N������T/~�.�M~}�z��s�J�D>�����s�y�kʀ�K��ǝg��/}�,�>�Џ��q@����iLI<��/*�JUp��K]�"�N�P��<� /o��� �Y�$X���O���/��e����y�ɚ�y�;1�Y� �Y�b��w��;٢�ӎzs���l�S��C����ՙ������mM�����Tz�ū�AG�٥2!WN)JU��m=.�&wb(�x�(]�3����#���s��[�K* ��� _�g�Mx6��c�<�y*���~ӓ�s6Q��h=�VƧ;��<w��ݻ��SR��T	D�u�d-/�<�j��0���_�*�ֽ�-q�����=�\K�s�۟����W�S����A#H|��Fю�nG� ���E�Eqʿ��Q���P��]nM�n���\)�1;�
��S;��s��u ��yK�Y]/���KU���>���a�חВ��yJdɸ�7@kBd]����J�Ѡt^!�7�,��cӲ��p6|��ᔲ���Xk:�p��V���rN'�1"�x_��Z���p'��]���f��I��zau��
K��Jp����g���<0vi�����J���c�$�վ���6w��3���u��}$��3��Y�ze��"61<��5�fzͯ{���πS�C�uS�Е>r��y��k����T=�
p��aY���y� �Ѝ��~գ�eb�."��{% 3���E�:�B�c�e?N�w�'���z�+'�?��mj蒉�'����1�׍�Rw��hK�2�C�ڥ�����MC���*U�K#+ih����Gmk���{ܭ�ʔD�D'�M�cYC*C���� ��bH��2fѓ�{����V��f�W0�>�`��x�� Va>�Sv����7geM$Ș�ݻ�Uv�G,����']�e�BU��'w
�V�X�9S��a�p)��GYGQ"D���2�k��iG,4��^����+:�#���F�IH�w�F7кp�Cn�ŝ����'�r"5<���Q�	�,�+�єI�*�����Ш�R�ɖ)�"=�D�o)^ꃑ��f�/�D�v�Wm�sf��M���mv�яua�nm+�v񨇞]��\��V��p\d��-�^K�6�;��}I�nji���c&�2��lX��"И2��_b�c�gYV����� ���%G}}{{Os�F�p�"Rt��80���ʵH�X��Մ�ĐL��FP#�2�d[���L�
�t&y��m{�z��B�	�-I'=�@ht��r�`�z�Act�v��F�1���|��LwB�S�m�t��ܹ+aΦ�i����j*�d��Ve V�xu)��f7�u!3*�խ�2�WCL��:�l+U�\����kC�ή���[��hj�'H���t�J��Z��-+P�n���V�J�T2-Oy꣯�v�S|<�ܫ,Z�.8�m�ҕ-v\�Vw71�ڽR�c絽��B��㽷Y����ϛu�X����	m"U�P�n���Y/����	.��_U��n wG"���lj�Xi�bZ����lr��L�Қ�[�hf�tǦ�ڹ�=YQA0Q�wr�xR�t؝aG3�R�i;v�i�1��е�\7�$��;�����g;;0 �1$��y����c�o��g(�V.�yb
� �][��ԅrw\91CRWѷ}��j�_]��6���e+O:Ҩv���8b���HF\������ov��)��2� �˥�+7��T^��^8l�9�i�E|1�-�Y[u/4�����#K�����H7�LՌ��'l{H��Y����[Q�63G.\u,�R�+�s²&�ƫ,�;�m�3FDz巗�]j���t���'���[r��u�\e�+��f;�gb����nN��
�5���|{7]!����e�7�N��怺#WX;7h����+���@�:�^�ۣ����s`gX0Gc:�֪]G���a!ڽ{��J=�i��3��VQ7P0αSX��i�uo^A�|ɫ`�iY�T3�No���6�tڶЩ���Ȗ�{�[6񼙽j���ar͙ɺ���G��ۻ��v�:�h�n����3���:
�)Zl�G����.ۖzV�vH�2����n��V�r�H�b���eJ$�x�[^��3K�Q��>�y`�7��+��ZS��$�p�wu��D4e�C��DT��e�4FMRQAEd9RQM�4�IVX�`9�EE�SIFYDC0�FTĔ�Y9DFa�.fa�AQ4�U�%Q�aQ31f&�ALQY�RS1�DLXc�4Q0�QDKTD�ULQD�LEEAUA0ALY�EDUADTASQ1�3ADF`eDUES�5RIUA2TTUVX�$UTE�TUQPCEUNf2UD�EE$5D5ELEET�T3I�UUMEQQ%U%E,DT�UM$D�KQQSTEQQEQM6YE���`���N��>R��/V.���M���l5��_PZ�(��LNď!$.M������'s���Z�P��ku�&lA�>���~�t����;�uL�����p:1H�w*�]d[�L�E>����o�T0j��#�2�{(�wm��8+	'\�_	�
�����)���2�\�Վ�G�ܦz�ǈ3������G<\o�"���F��x`�	=<3�|���AR�lx{f�w}�/�ӑ;�o(5��>tۄ���^fo�Q�G�(��$T)����������^�C��z(?���Ki���x�<��:u�nT�����* O�أ�n:�kw�;�<��1�ʊ*]�S���Bu�I���e��B�:�r�����G��c>�uw���1�E��p�UA����a.N�,���Nv�mށp��Rۃ�A�_}�=����v��o
u&���6H	�
�T�82gc�EB��ܛn_ϋ�d�{3���B��0۱S���ذ���{^�F�H]4=�Y�S��W+}�脗UQ����5@C��¹y��]|̞��3XU�Q�ש��|.a��'|b�v^}J^��1WC8U��|{�E����&�����¡��ي}��$ ��V��`}qxOy���[�7w*b�,9q�#�;$����YD��o�c���8vѥ���A�]sq��i6Vݭ�2u��oeN`�cF��w7�j��)7-�K�9[J�]�� �`���������Wt.<�3p��'n#���޸ʁP��2z��-��a\S��g��mߕTf*�^}��\y䚶�
������2��9��U�[-��s�z����$�|����~�Q��u�����ϭ�V�q���7��Y��C�UKI�,k)�S�Ǿ�m��N\w a�Y���x�s/ƎN�L��	�ƼT	��j��T�2�%:�y?Tf�1F���(�IUz��n����}�({�p�(_�L��tpJ!��F*���|����]�m�	^���^�����j�{��3W���[u��g��Y�=@Δ.�_���xռ����_���j����}7�f��v�=��b�	�g��=
o�kknY�Ğ�3��B�{��7�w�M�{�~�{��C���;�C���U�z%����C��c���=��rG���w4��ޘ��[s�Șw���=��B�n8�F{����ye�\*V���-N��C�o:��^�'��ƬG�[}�>��YI�]�
j��9.N0=�����Fx�>����+�(�3�y�8z�;����cg�^.�[\��m$P���D�J��Z�����J\���x0���|��1]p�{d"7���.�(�����7\���V
+��L6�e͛�)�a�u�d�*۔�gPo�s�/,j�D5�ohI��Lw��Y���{V�)�FF*��=I�̛ˋ����$������0��<*ӽ�Z�IQsm�<w��k��F��>�5��x�=�_�m�����
fe��!u�`s��S�����!?a�C��ީz�M�8�n�>.q��zB~wj��$��v����Q]�X$W�̱��J�i�:�����!�]ȸIS%�9`k�7��\
�k���q�_��Q2���o����3~��]g;��9Y1�9�-���N@R�N�_����p*9׌�(�h���*{ݺrś��������A⹝�Z9��*��ie^������%<�b������P=^0V=�2����F�q�5Dj �xta��+��]J�p�a�j//n��xcܜW~�����cA������|�}��+�7�|�a��>�l���2p+��Q�<쌔מ���ɟ1�>���1�����ԯY�'4�vk����u�Ў�qaz��(]zk�쬀d@����B��Br�kx�\yVN�~��SnVS���Oƶ돾�>'���/��a�_|Њ��ɯ�ۏ�+�Q��"L�3��c炐���(�9����7�eȵ-%�èk�����׎o�@�s	؅{lx�cڒoffQ���'mk�� �^ސ���>��]�՜%E�p�K�l�R_��v����t�����/D�Zs��xTD��w�ڞ�U����g�T�@�@v)�敺A�|��1މ^�	���sĞ)�^[\*1�w�{�o'�)�Ηr�_�e�tz#p������%����>�;T�zW���zn'�_7]��𨸯Wy�V�)�q:>�RJSR��/M#X�?}%���(�{�At �t������
�\.g�^8%�Ut������$�NU�𮞭���w
d��4��f���#�Z�q8�[�K7
��� Y���P��	� ݙ�^���7����C��cq:�&�㸜6���\*��o����H&><�h�	�s�j�J����~�J~�̮Y�Y�10�}پ!�ՠ˞%�p"m�X����V����$�>L?O��ɚO.��^�k����\�m���ʸʎF�xT.]NKjt
P���'T���UA_AZ(y�v�k�\mک��Nl����U�Jg(�^9�.J��yJdɸM��|�5z��1ZN��N{����P�+z����厍6T����+�#:�p���w?X}�P侑�?M�I�ua׹e@��F��}�;ޠjWvY;�e5���k��*oV���7a�����p^�7�yu�:�
�z����]f.��#�}���m�������Q`����1f�C�μ����t�5x��[���s����J��`Z�4��U{Ą9p��~�T�Q��z�a�7���=0��e`WR�ฤ������Z�����i����?]��9�Gu.�z���f���c��7	�.�_O�=�9��^�1��+�u�s�I���{!���o� &�+�����>J�9�>�zs^����8Ne���֘6P���VF���1�_��|���7G�=yHغ�Ȟȕ}
��}9�y\;���C�['��R}�]�3#r�=�[�U9&�vA�t��E���u@�@TGr�e�[�L�}O�3wӽY>�&��a�ϵY��[9E���z��C���EL����R9J�,��0��.�ۃ��y�]Qv7ttݮ���N�����7���5ă�g@��BOO��_)�/M^f�Ѧ�+�:uɭhX��(y�:��j��Sl�聹R��ĕPg@���H�����>���2��̽qX�fm��P*N�5����a��|w���8�L��" r�3���r��lUw{P�}�ׄ��]�n*�.�B���q:��<u#U!I�˚�{���qﻓ�<����EХ7V�f��K$2�`�#%䮣ðV.ōu�>�A3ae[Kp ˯�F�Ŗr�bZ�s�4TT%��ݗ��K^M�y���Z�snlAvn��IR������Z�7N�fj�~���%�o�a}�P�_Z����-9%�����$dbQd{�P�����. ��O��T=�W���٢alrv��9�il��v������m*�A��Bq�c�i��T�-T�� �n�T����=٢�Z]nM�r��m,�N[\n&�;���{���*����-W�Ѹ�F�J�f��N{a^9���UU�2�\LfGo�,�vd�r�k�U�Y���NOx\��;�+��J/Ʒ�%�?z\3 �z�V5]<���+�=��п'A̦X���Xn5�T�S'��,��U�po�,]�ړ���qGt��c�b//և�ުz}��fnU�[>Nhm���y�s�[p#�q/�o��}�����ô�>U
�O��E�8o
f�׶����i>�T�3�U1[�{����t������d϶]�Ƨ×����s��W���2x��*������*k� �>g~�-�����lj��'�R���/��by�����x[�%��_��)�ܦ՞t$�*<|�zv����b�0����~���7x�^5�\}���peT:P�/�W���+�v˕���cli�VI�ˉJ{�e��]g�Sb������m�E�Q����ps>eug<!�w���V0$2.���	���{ڳ�d���y�ڊ��n��݄�E�S��P%��T�Dv�Ǔ�]������I)�j΋����-n2X����b�Vg{�r3�s��v�{��3ވ�\���16��I�3��B�_6�e=�}��˝sE�N~��t^��߇��l���Ӵ�D�W�R��3.*�]�Aء9Z)迍� �,!zj��e3$��U�TWOS�mIjw�h���L�l'v��pJ��/!�~7�x�v�{��) j���L�2��3�i�y��\*W�}
g�-�㧆̗��3�U���^���1W����V�_*�,�(#���d%P(NxW�Zj;6�/B�i�p�ig�����G���.w	�I�N\C��hZ��F�H]p$�Ϧ�����c������/�VγSJQ����d&��2��(��J�5�I��U©�G�!v��1R��k��2�;;y�'=;�WO���-�!���rR�p�F��W�ǮWNN}�I|Nt"e���f޵�����8s�]��y��^=���Utn<� ��;`ih�=P7�ʍ�G���p���̽�������m0C�~���V�1����5�]��O�����LV��W�{��㑧�Y7�=�dc�*�3�A�d�RK��E����r�Y[x��V3���
�{�6�JyA�픵�0ւ���G_V�"����Hk;im��ފm���yb�{��;�!Қ�q��eV�w���&�N�+z��J#�٧���=����@$Ly�c��cs���򷨃ƾ>�:�Nq�z�ˈ�XN���^^�/}SOdw�Bn+U�S&�ۜ��l;Û3³����O��>�?9''.&�8���]?���%���9VZ�ܧ{��oz���p}U��=�zϾNi����(������2���?p��՚���<߽�|�I94�p�y<���"�?@�mʗ63�{\/ۮ>�>'�����:UU�,�2�o�xVn���7N@]p2�1ށ����ssYn�k���^��ۡЄ=��ܷG������[�I6\��Fr���eq�������ᮟ��Y~_=�O�Җ6oá�pd\�Cr�^���z���U���B�qS)L]K�G��H�%O��,�{��s�i���;<|f�����g��I�-�X���������<DҘ����м�AV�٘����y=��k��V��z�;�����0�T�p��ʌ���)* ���T!�q��Y�_�ۼy!�9�Ї��V���m��	�i7��q8]S���Tԣ�@]�@��9�U�ڨ>��O��}zo�:8�)�a�w����'}Ϭa�K��[���N7��wxQ5��V�6�Af4�~�O{�_�s�/vI���op��p���e�	ث��!�����|׭u)Y$ *���t˵b�Aݝ$��|��OVf�r7;0�r�5�qQ�����h����<�W����&�|����D�ͺ�.y�*�US��m� �/�po��u�M��{��,����ѐ�ϽP���¡\G.�&�u��L��^lL�ڱCަn�8u�4�����WN��/k\EJg*s��߉��=J��k���L���rO��jxz:'��:=���L�\.��56��r�F�*{�YLU�J�_Fu��f�ڣ�V���ɱ�=����y�F�rnJ�;7t2���b�}$��0�2p)/�éN�N�pߞ{�vǲ6wd?r�趆�J��R��c��_�f���c��7	�.�|�H̸3��)�r�n�]��7B>v-lz�D�.��9qH1^{h{���>J�9����5�`�~ˡ��8Nb��NsVtf:{3x�,ղ��;�7���Xn�d���������ȕB�cNBy\;����"w�y�.����=��"���P��_WUŁR�8���u�4�E�]�2�''w���NE��d��9δv�Ǔ�-��V������2�T	�
I}1��#�W��~T-�]���qy<�&
Cݿ�
߮3�E��k���Ng$^ܺ��N�'�����[޻O!�샎k=ͧ��l�A��vdXm�����h��
��)���\mr��:�'���suҚ/��H�cf⵵�b�FvH�]�ر�mB��Z5s�A޹7,R�>��@Vw�G(�GE:��z����e��T���|P����uR�M��ZEc��˚��ep�s��B���:����{��e��ϸ�'����g1{���̫��3Y��d�B����s<9���P�I��G=��\<���;w7�##���s;5]1T-�ˌ�QZ����f���[��*�R�pG���|�Fq���e��B���b����͋yJ��$a�<��eנL-5ٵ
�;H���KG��f�lL���U^�=?���F~�U{�\mUIc���;H#��=��`)���EBK���B���g�����?q8YS���U�*�f.��$��j�}*u�G|f�<�{�	�b}>�����n�1���1i'd\7.�B5�N��\�9�W�v�T��������ϧEb�4�[��~{��wt.<�3',�Q6s�q���\��sES�5�6�s�R���M���?Uh�~����{E�h��OO���37*­�}	��~��}.<�{��Ǚ?K�Q�tm�ڜfn`g>����(J��;��V�l|WQ��������.�u���S�$���OE3FH��o:4��bn_u����*ZR>�]�:�)z�=�����z�T]�*q�T�f��J�s���8i�]��r�oo#�������W
rmC�&�(��4g]���ľ��$�3;�|'KjJ�VT�35!�Ѵb�"C3fN��W���ʢ$E!�o���+��\�0�v�u|�Y���h�s4&�N�z%��i�ᬳB�r��;�#P�4FT�ۙ�Ί5�;�ѳ.�g<�{�$�5Vvv�ǉ���3I/s'L��]�n�Z��D�7�3/r���>���L�vw�t�Y7+ϋ��Vl��`�o�"���Y�-��ë)�Aj�ff��M�V���"VSf��ֹz��i�+�c��Ca���z��W��=�cv�#G�뒶9ݯ�E�]\�m,¡\�V�gr6,bT3>@�����m���n��w|12�w|0�	FQ�Q�K��vR{�mgVʲ@[�T{����w\y���x�quof��5yb�w�dRZzSnIV(�G���"J5;]++]�ݐ��v�ëZŜ��X�yq-0� 3 ��p��޻��u�M�����l���&.@���I����4��cGi��Y]���.U�q4ma�*�\��2�%q��ip�#n8����a�h�t�q�;O3j��Xm����oL��-��9u7�ݮ�u:��v^����:x�;�F�
:��J��93"m֌\%�ki�[V�@��֔��<��;���xM�;Y�ӵ�����I��v�7�e5��녣ɥ��ua��7���]��Z;��Ȯ��S���Â��S�n�Zp#;�pv֎�*��5���C1���Nm��Րj�-��j�L��
FD�YYE��.����xM��kS�Zu��Y������D}/;L:�fe��`\�����#�1.�*\��,a{�9�0��/k1�Inr�S5r����j�W]��N�C�[��u �qz�o�^�H%��n#�]���zX���>V�dF���KX�������/Q���a�w��_1�
(м(�ΞX��1�vq��4l�wZ#I]�w��t�.�&uM��w�ڹsr��]o;D,v��+7�gZV�}���)�����{Nv�sX�Bc���G'�JՑ�(MΛ(�&JCO^��V�˕�to���̗�����:u�rZ����� �L����T�k+d�7n�}�ݎ���@z\�ڭ�
��g�K�Z�Xkof�	*[��%T��Y�d�s�г�;�v�Eͦ�w.������d�p�3�6�0
Q��҃G.2����1�Y�>S���v��M�Q���
�iaZ�;�6�9���S�:n��ۥ,��@s���J�h����l;�녖�+��ئA�>��/��Ϟ �O�ʻ�������(��*�����h�"�(�	/l)�&ifb���a�������l̂i�*��&��(""����&j(j��
Jb�
�&h(�#$ʨ��$�j�������*)���*���(bH�h�(*����"h�2J�*��$�"b&"��h��j*�3J���
��*���"�
*�(��"����)�����"*��2�
,���1ɬ�32���������)��1�� �(�0(�&&(���("
���*(�
�32&���������*�&�"����"����(��*�h����J(���"�#,�"*��h�(�#,�%�!����J���&������&����**� �d����J׾���,���N����M�r+��h�ͫt��^bfc�+�{�u�i��%��ٮ�/]�g�*,��Q{���4,��]�1�}��x>6s*ש�����j3׷��UOO"Ʋ��1Zy
	�Zy몲y�W�OGw>�e�LW�钧��Ui�̑��LF���<g�}��U��df�]���n��S��Η�ʯگ�v#�'�TC��Қ��	D>��9� Q=˳����vצ��q�w���i��;�����u��l��TWt
�O��~㿅w����XN�e�m����m��}:�
��n؟Bt�^��pz��kknE��NјZ}���a��u�Մ��$ޗ�Qc���/@����-�/��CۈN�|}��W�nT�VX��if�F슌]�|��X1����;�<���3��0f;:�>��������s�V9����2���v����ku��G�q�H��I�#�
��������ˊ��J�ZS����w��^I���7̣ͭ��iNpK7
�nU��tM�=��qօ)H�O�6緾5Rx�5��#�U��?���|��廻f��*��n#�� H��🂈���{򮰝b�Զ�f���V�Q&�!6\�,wfI*�]k��͈?��G5wUF5��b�c�]�PU�\b�;�te�v���im�Hr]Q֧����,�2:�.��]d���G2oWJ�r��e��tBּ8����A�:`��sp��
��u�\��~�����C����}�s��n���QY
���X��y��x眝�\��t\Q}�Xt-��"+{]ȴ�2_���B7�?\
��nM���}ۉ�Vd��D�,���j���gިXw_���]��Xsp��4�#4=�}�4��R�c�N�hsy�8�^���a��"�f���xW�Ge��z;�ޟ}��Oex�=[މ��Qs;9�}z�O8J�d�c����<_��k���*���dk�N���חP��[�>�L�C�#�78�?��W3�LV�����4�~RNN_�?�P��Qo��Et�'z����v*}~��{{_�>���uS��c<��=����c�]G���f�K�ùw#:��ǥ䍫�n�CՎ��>�2��w���|�Ъ�=�n�7Ky<<�*����{W{��DH���e�p޺�(�.�C�uL�t���eC@�@w)�敺A�C��pׯ�������<[���'ؑ��㡎.t�Ƥ�4faTI�����}�L/@�QK$������R�JϬ�1�Q�}�Gf)����Hu�v���uɭ��;�¨)�FEW�A�#����W�O$�s�޳���Ug���Qn�P�4��r�L6t�[�F���le�\'�hҝ�yY�)�ev�uI��ʴ�D5�V��7��oT�MW�{:����] �1N��$�D΁!�B��g�T}2�x������v�ꆼ��r<�Þ��5�r��y�|.��%��2���(�"*�΁?@��h���T�2���g0�f\.���n�����,t������*��F�ʖo�P@�Fc`$@�u�
	g�/�w�[[4���ވ�R��{�8��N�I���pۻ���5(�qTiު���������㱀���T �O`L=���_ܚ�<�u��p"nu�\:��UV�M(�nf�/�zF1n��$���F��>������	���P��r[s��C�e@�ֻ�9����s���I��n��NH�gv?��N��=��~��s�S�N�[�ڴ�:+��2sz@�p�G�]MW���|b�:}CU��#�lJ}��}��r�u
���3�V�O�mB}��G��Rz�vỡ��a�ē�2am��
�����N��qC=�FR�:�ٓMΎ��߃ާޏ|��f�M#Y��+M�~˯|�@j�~럜��s�sV��R���J+/��m�Č��NG��Z�����8���󍴅��f��ho��v��;�:]oZ��kJ~��*?b4����ĜM�31ab���\{,F%����y��CY����bS�QO��Ѹ+:�)و��F��ve<�I.s{���Ѕ9>�(�<�B�����x���_��w���~�V�ԕ���?~2]�~���&�飯�e��kQ�1�~'g�����><�ULc�ϡ<��+'�Wh1���I��ޮ��|r�%\)�<2����Pgj:�����7\�6���>���`��Q���ۄ�8����-��5[G���8�(w�L�WS/�/�R��g��O�K"��qf-���P/OE#��uGM��j{L�辒`�(\T�pfMB|��5�r���o^��s�/�4�j�<�,{�B9˪2����O㤞���fǏTU>u��M��0����qS,rV�����R�ײY�y\'�n���H����°t���1q�f6 �HzS7F��7qV�w�yNS㸝Fq�x�F٣2w�^%i�3��W�:��K��$a�=��O"��	����jN�,�a\_���'�Qw}���{��{��.!-��3l�B��(\uI]6H0�=��d���
����H��x%F�����7�T�;��	�����6�)8�^��'n��v�wO��	&�lq�x3�V�^>�cs)L]&���qu�7ej��t�������g��I��d�Z���S1,]-mR=z�:�v�F�l*�o�}ڸ媀�3:p����l�C>d����Rul�7.�GL���k�����
Rn�ok���2U��m��ގw��*��]ыI;!��c�Rt<@�k���}Q��vX\�����#+�U�O��ԧ���ǧq߃�wt.<�3p��6��W�ƸʁMz�Ogz�����u�׷�oiB�pF�J�x����\0Wח��/����yVl�ddO?>����.q�I:��KR*�6\�JI<��ps*�W����c���^�}�T��,k5�G�n�ΏS����6J�f�b�]�'��=�T#go��З8�W���Q�H�w�nM��ӫQp}�����F��Ȁ�c)��n+��*�j�KE�#�"U�GF�3�|���r�[xy�$HFz:U�-Dk�y;�_n��`{�T�2�)��u����}�ft��'&�m��2.v���7}����f����2h>��p}؝�>��2���AU�b�[r/�:I������-�\u����W�K3���ёÒ��A�߃�[>P����v��U�O�2�~�d��4�A	&�}���v�K��ʔᔪ��)�9,7�h�}�a�5��*�:��.`���рjR����L^�obJ� ]�]_K]�j؊n���ca�PE'�V�.v�u)ҹ��n�ڲ:�����f��B�3GP�/��\�g%,��F�K��rw����I0# ��Q��qS,s>^�3�m��jq|��zEO_٢_�Tw�΂�K�o��Q��V)�:���q�E���;�.*�+��30X�]�ۋ�+�w(�s���NX�G�!�Z7�s�Y�qU2��*�Y�8ak�ۻ|��\�ОӶ�{�9�ǾNw	�m�Y?I?'�m��=΂P=�SN��:��j�;ѳ��qߊ`Ø�e�׼��=_Yg��"m��@��󸫅SN�����b��<�'=��n���}��7E<��������w"�%L��偯��x
�O� �>��x�
��柊˵9�m�.�sM��������}Wꅇu��K����)a��v���y	�إ�����V}p+��'�Hzs�஝f���xW�Ge��{����u�R��mə�KGGv02Ni�8�+���d��>�����t�_�+	Ã��o2!�NF�=�~��<��q�;����u��(V?߮%��f���>�lL�P1`uH����������!�Y�w�o�L�힚�3���R�x��Dmp�s�+-^z���8�ܠ� ��zkG.=��9�J=�;��S����Û�$[Ĺ󷺡3�c6��oQ��g�H�J��<�9(������"JL���Ev{��wy>������nX^[�C��N�ru��sL�f��1q��t/�A ���唻��u�kO�l��#�7���ٟE��(�+�A���r�h��n�7O����5�\|}�͎�{����r�*vM�=f��F����R�\�c�b�*#�W75�[����m�k[.=��dE�n;���۠�sĞ5W��¨�2����o�����
Y%�C�Й�ܐ�h>��ۣ�ç֣��·Lw�W���.���<	=_L�T)'�c*�r*̣[8O����z���l��:՗�%���=����>e88%�t�U�$t�4J`�{�rX@z<���F�k̿e.��9��ʰU�V�5���#\G�\��ه�R�*�:o=���>W���]��v}�k�Q��E�K��>u�9:�&�x�'��qV�Գ�1<�:r�޳�=��@��}�A;��[��!��<�լ�g���`7�Ȋ^��~���fQ���#�{�VL���F�� !��=Ei���a3Q�*����n�׏�QΨ��~��e��3C�=C,޵�}Nu�X�ur���՜��7#��~W~\}��z��vK���;��vH�¶�XB&�'�t���W"�W1��12mr����MAf����r�f��D3M+�����(t�]{��\�
bY�}��I���6&$�Ռ�:�����r��~�B���:����+�i�蕴�]K�p/�&^0���粠\.��;:����L�܁���Z�x�����O��cg¥Oa��N�VN���M�y�V�WJ�ƴ����kwtb��R��p'69��#�ē�2ald�Nfq��s�����J���NG�h�'L���doS�G�k��nM�[��+M��]x�I'%��%�-<�U�yGn��ӎ�|�+��O��Np������C�uR��	S�>��A�O��`\7���7[$��ݾ�ٵ#�'0�!�a�Ez���O\e c�ceUs!L��=���Ǯ.hvz���l����WзՓ%���o
��~�6z�.�r��OC�����1���C��/w�O�o�UBg��'q����\cU�xz�'�\���3�\EL����H].kۥ��x�ɭ{� �>�S�+�]7)���z
���Xe��Aރ,u<PR��PG@��+o{���*t�*�9�Y��vǇ��t�{�t��C����(��R�� �N_��<�WO�ʝ�QE��idU�^���3�O4r�׬i�v�1�Rݯ+�>U��K��V2�لŸ�1���*��+x6	ٖx[�'[�u�.fs��Ѩ��0
0���Q�6�3�R��n���R�t#��YI��i�Cc���ݙG�f32��u���vP�S9S<9+W�CU'x=�BZ;致Yۇ��p��۸r���}��ئkm���.5 ' R**f���*�.�G�r�ϓ�3��f�U�*2M~���;�˿XZ=ն�c�]��f\� �*H�?�DJ�A����|��nN���V�ꉉ"�[���y�9�����$�F[��j�UT�/�J鿉ds�%ic��/�k#�g��\#7g�yi��q��}�|K>��+�x晡�����\yo��nr7ylZn�����+��㳙:��9L�.��.���vY�r�k���z�dC^�&�fa��S2fW��{��9�m���Ұ�䡕��1脕��<�3p��5�Q$9��՝bek��^�񥲉��b�[�^k}nd�sˈ�0�)�a�+�F�/*��uz}��fo�aV˖�**'&���Y���s��=r/zI=����̨W�z��+	�a�j3׶�����yC�1�NfE�铔�w��y�x^��+}�}�;�Q����/�Á{��V��A�Ǫ�Ufr����Gߏ0���N��1U���F��K3U��N���f��^@�'�<i8�;%���r+K6����"��+��"���'P���NP*G�]nn�=��q�nT�=���j�y�C�SÛ�lL�� �W�oW(9p���,�]�3���=��T׭�?���1��Nf=�U�S��L�b8rR^_�#����"�����g�pbnpp���A����0=�i��O����x�5�\zω�({��ʨ�Dўw���:��	�:\S��\@ɠ����b��+�2�N�=
}��3w�SAJ��A��bN�Q�s35���S2�� rYR�[�C�-��=�:�����޿z�ew���w��O��I�1�$��We
�R�#�ꨞΦ�C�-N��mU�	=ba��j��Gii:C}���i���@���wT��#tg�g��.+]yTΪ�xN�z�'q�}E�yN"��.�����eú�W��ͨ#���6��{�1���\{
�s@�o{��%���֎�Ν�c�sm��紛x�'/�wlиUU(�Au@�6����nvꔛ�v�Y�p
^��	Ӽ}qٶC�N�C�_Yd3�N�6�2����M1_|{,���܍\�S�����n�����g��u@�Ʌ
w0ۣ2ׄ:���ݝW𨈊�ڢ"+�(�"+��\TDE��"+�_�TDE��"+��_�TDE�Q�B���ʈ��*""��DDW��""��Q�j����DE��"+�����j��������)����Io��9,����������0�>��T��" ($(�T���@$�P��J@%�� ���J�Q$���UH i��� 4${qB$I%	A%U"*�EJ�*JH��AJIB��H` �E��-�*�D4�fCFT��֩Ъ)�RA� �DB����� N� 
���(�ws2����Qm�E�CX� ��HUu�EUlb�jV�%Zb�JR�3b�UQP�q��ـf ���ڀ�2�,���AFF�HTI$���6�X����Y�M��0��(�`f�҆Zѥ4TT�"7 � �Dj3% ��E6�֔� �QEh��ЛeR���. 79J*ʢlȪ*U3�D��!h���Z2$0B�U(8h7H����*��B��
�P�4�X#$R� �\��KX�L�l�Z��R�T��R�d-�UET� � ���Q�`�f�A��إk%V�AHJ@*
L*RJ� �hd� i���
R��i� 14ɣC0"�2�0��&&�S�x�Ѧ�x��A�~%*�~��      4�ɓF�� �0F`i"4*I����=&O(   [��{����K+Z�ZӅm�R����%u�Um���$h����`d X����Af	g���b*���3��� ���>R?K�?�!�E(�H�(��C�O�C �40	�d
����]�����.>��k�En�-�&gY�'���ڇ��'�^����o�y�(R�"����i���M<�֊ OeؕkHKH�(n0���K-i�+V�0^����J��g�yx�YV�ng."���e��/l�([HZ���p7�6�i��j���hd����š��٘�̉��x4m���^V�-mu!����~�;R"�52�c��r+Ҵe+�y��I[	��i;���|�=[���)�ծ�\�ǜ�8�_k�8�`]-�ڞ��SPx�!R]-�eS.i�F�4uV��rZ�jS͔e�HޭM<�)�P��ϔ�9��h�n�)z�$.���q�C��Wp�.�g��vX'��j�Ir;{wU�Q`��"�B����J�m
I�$l'�Z�����8F��܏e�X�;�4�L��nh��������
�PJ��Q��Ek�<�w�X��|��W­h�QidbH��x嗙��=���oz�#�hm6�2�CtJy��5V��5PDN�[�˯��^�Rٺ�
л�����O^�N	b�c�J`����r�T�E�u�"Ud�4�ۙrj
��8Į�]���V8[�M=���]�GlѺۑ�7{Nn�Dh��ɦ@wR���z��*�S���:��G>��.��y�����Հ1'���e$qv��9�<h�.�K���\2�-��,os��L+Ae f6-��Uը�m��ѧ�e�N�D��UQ	U���R*�kj��%Tk4��Xg+��EDY�*�5��нŢ�'l�Xh��j�n�m�ȃ�ѭ;x;S2��f������ӓj��Flb�ɡ:AH��;Y���t���٘��r9Z��Aaf��&�f�5H@uc�Fn�oB/̠�r�.�]�,�m�D�t��nk�"@��Y�5iY�w�\�" кu��q�o��R����/�n�K�f�-\.�"�G \���.�`��{ɝU�(�Igj��DX�n�0P%�E�;�Z(�@��ᬭ;,G�J��*m�R�gB��2��N]���#�T6]a`*�v��h�Va˹v���-MĪ%&;Վ�uY��e8�,SH�Y���+5+�Ci^�rX_R<I���PN�پ�o����6Bc,��e=ա��v���j��&LB#�X�Y�*�Pb�=���|�Nl۬7Ŕ�!��S?c&ZZU`�I^�0�i�NjI�*��c�f�Lݕ�^�J��d]=@gRѽ��ћ�,iSY���:�0�9q0�9�S��MSM]�ߪ��{�Sf=/�-4bb&[�,Xb�b�v����:��ɛqӊC
�5|F0�k:@U��)qWx1�|1��4h�&b�8�e]���\���v�v�u,�GܥVHG�v��NƼ�
E�显g*�]lr��Y�mz��2��f8lXɱ۟bYYZƞ�=`;��r� Ǩf:8:�c�ƟfՃ��k�p��ݹ�ܻ�4����tV=�x�<���%���:;uXu_V���V�.L���opX�w���bc��i�͡T2�*22�,�0!�Z�����\���j�&�H������^R׭&�4�弨�2��	8Ob[I"+�;]�(^м��Y�a��3��pA�s��i��Ç�F��:T��/XZ0�FɵH�r*.-2?��(7H^Kt��sX�ci��@Լ�T̍�����N�^S�x����l��eY-�v����^�k���<Z�۠��� |� �k��f��3AŦ��볔�]!� 1�K�N�i$�T;�Bk�i��u�_M����|�_N��!Y���X�xl�95�WkP.�S5�6�]�̽��[
�٫9���3g.A�5咔t�9{&����lH�K�`��m�V��9�y+�m�+�tH)�łո~��be�q����n� ���!CK5�mՂ�ba�����j+��#���H3��$�D�o�=�	&e����O��rk�m��&��r�;whIi�W�ua)V'�b��{���t��z�m��-��r��j�pf��э�XY��˙C �33r�4���eق�kFf:8��B�:۴r�[���XY��h�����0>=a�sC����.B�-�3E4�C�� ˼��E3��� �����u2�fM�ݥw�)�NiCB�^��UR��p�G%��gR�s��ͤ��kq������/�!fV��wGb�ݳ�3���-q�Ѵ^����ػ#��x����U*9Qa"�k���C�5��ތm�6�;�î�\������6���J����$�`�q�U��wLڼb㓞�k��t������U� Ba�2F�(C��J�1g�%����݅��4��
�{m�)*�X�;(�WWkF���%n�u0�SA�Aƪ�ػ�+kT[[�m�w*]\SSh5��I@c��!+p�(v.]�eUZ�z�V����~׋��93V[y�2�9\���f��|o)$��z���Љ���y�ɽ.�G7)��ɲy���� ��H�"�t���UR��%��vU;��A�5f���3è���W�D��H\�.�m�v�nnۣjb�j�I'}F�:�gu�p&)��X�}������\�b2�mX;�^V�N�A���=)�4�#��l1(�(b{n�<��h:hr�i��e]�cJYőx*�����3(қ���ca���8-�{H�����d�Ǜ�Y��wA@��ٴ�e������a�L����a��N7�A齍bm�4���d��mk�����M(�n�RZ�ٰj�,E��0L�n�gPw��6f��J�V�̷r֑�r�n��	r��JH�X�e�a����W�����}��9��b�t�8��+}�"/b$=�^PG��yϰk,� cκg��)�Z��q��Y�Ԏ]���_�W%��/a�ɻ9g�|�k�w�L[�4pR���$F��Z̴-�@�ʨ��u�n:;�e,���G�x H`����r*�[���(���%"p�R� �K&�]��%fՆdx0����h���Zbc�N��Y�P�c*ԪM���e��UF���Y�R�h��ځ^Ժv�Jݍ��ȤEMܗLJX��ଙ���śTD�%�ʶn���4
5�u�ͭ����^h�ڠ�m`P��k��V<���@!�tv�䱓n�c���q��Ő�Z��:EU˗a��@��X��U�KF��}dvM���9*��=��$�M��&�r�Z�*a�h˻[��!V+�N�of���)"�1���$욓R*AdKJ���tՍ����E��X�a�3��O�za�);�$Ae��wM�j@�7�Fg<u(�����������w������~xf��w�8����,�/��.�ǵ�#G����#�e��]W]-Q��3�M<���F���;�-�U�y_��h�ХR5�$7��0�%rM�(��W&��c9�c]�E٠kTX�<���P�kME�6���Cz�����k�9�}�=������]�Sf���,�.Z������8V<�׸v�ï7Hm�i�eu!�qoV��`�m��K3�*��,\�	L��)����'*�n�Z�j�O{DDob�&��W�̽�:�g5��P{����8���eqWm:�V��"��ӊ��^�<�f�}t�\��v�ڙ0��(�D%y��Ou��9XΩ��CL/h�*>�#�r��э�Ղƭc�7�t��/����\�A�eL� ���[ ���9�P7V�u��m���F��m�"�∂V--g}��+�4��;]S��]c�7�IX��* ��i6�=�8v��W���ޢhC}(u�x��*rRK��Yz;3� �p5gD=)�����g���j-l��[F�*��rpEQ/��t��Lz٣�3v���X>wc��R�����\�o<�q�}[8���)e�KM��kCnDM˻�Ë{h�[�[�d\萚�7��u����iP�8��\��ӷ����<�I^�	��sԆ�lV���nS��M�*�U�z��-�Ń0i�EnNֺBnE@�JsU��$�	](����fp�W6���w�v��2�,��d��_8VNj.ڬ;s3+��㲜r􌛴��atks���;Nf�wJ-�O&�M}�C��j�ݨ�-!���כE�5�9c��5��5ϻ�G�f��t���q��o2Ɂ"���g$&u#f�FH��R���C�����N��U�ﳥؠ�KX��Oi�t�\!t;>����*�Ӽ�&��P}����Sx�}��t��g9��Rf��5&La�������o%�sח�K�,����f�eb�bAH�GH�v]N:I铅Zy�ơ����:�S!QVRu���)�­�=�a��Lu��"��d��Y�vP�O�S���Gn
���x�{��(�u�a01KF�;v�+$�ᡓⲾ��:9G�e�����-fͮ�"����\
�XCH���T�`*��6*�זuU������]7��o{�r�'TL�7rūƽC�qi�-�"�eq�Չr�L,�C(�5c�����U�0t�m

p�����j�N=�gr�7����"��g+��5:�3��]�׉��(�.��Fe��/d�ݬ��
m.2c��[�]
=��V�p2í=4����.ޔ㏠#G@xtҰuvCʺamfh��P@��<I_<��}8������7+����}O5�`Oe�T�<�ni�k����.��Y��ي��W�M�u���M�u�ǅ�ڣ�kn�WG�X�"���E���MX�~\�Ѕ3$�^օ�עu��'c�
v�&���u��Ƭ�5.2gt�-�6��7L�q,��8uA��E����T9i��l��Z�b��M�ܲ�v��}+MY�S)�aZڻ�bQ���T��j`Д:Va��fem%Y/���K�v%�~�m5{�L.7��"��H�{�Cr����`ծi��^���/-�(���)�m��)3�ϯ����d�{$Z1��$DlGfl�L��MgN�$g�O<��{�le<����Ge����adLѳOν�]$��������=*x�@�BV��W�j˳;#A�DG�u�-�8lz�
�_b��g,�fL6I��)�W7���
 �'���Μ&dg���T����w\[x���M�u�	�ݜ���i&;+r( i�!�ɤE{��5:�g:�f>�O�BY�rf�c�+�l�ʗ.���Q�v�ikI�J�ں�H�Tͧ_Z{z�):�\@Jp<�J�Yz���T���I<I�cn�/pweR[O�;l�ݬv)��ȘG�+z�Q�K*DVf</�%�v�y�_
�X�q�[�ۏ�A��e9r����F�l��[V3:�k�ޑʴ�T�%T��u��v��IR�-�i[�y6�1/A�hR/h�qf��g.��GU���n��k/�Wr�w�)A�u.�c�M�ٕ�|��n^�7���BU�׹�[�6�n6J�&�]����� O5%Ŕ���ޡc�#�������:N�"���3�倀�eβ&LQ X1]��8��0�p������;�B�g	��|����J���Vnv��/���Rh���9�b���x�F�ͻ�[:�yk�k0�;��@�퓕�ԽY.�1����2o2�L�tS���$hs{�}}��U�#��yPi(V��܂[�*�fh��W�f�[�y�Q��2Օ���'�ٷX	08�ʵ����h"�pӇ�Y�{;I��
U6x�2w�{�όڱ�1X�pԔT��s/�h䕥��Ff*p�f�A"�cb\�+	�ypf�ͨ���κ�$7��X<��:�w<U/�d��j�V9t����JŴ��
�2V��7��y�)����8�Ε.V]xD.��c;��d��Rj�u��i:��
�X�MP�6�ѳ��]�lZ��Ք��r�nړꛭF�C��e�s��,a�'�,=�.�w���',}�.sw�I��JGp�:�gr�uY�'.8&��%�\�ӌQ����J����.D$�6K�I$�I$�$�I$� ���%X�I$�RJ���R�Kr�2�:���n�g�^* rU��;�p�)9=iÎdE���/6u����XcP�5�hj��}��,˻�RG wSD�ucLؤ����
��܇p��d(Ζorc���
�)�G(?���9�"X8��{� �会"�_C��Ӆ�����,�d��ٛ2��S�FK���/Z��A�#5�A;�lN����l�0h�l�9Ň����E�uh�ۓ�Yd����*���g�Uf9�c��e�Y��P�L�gN�+5�K�|���a�j���-��"�!��&T�+���带K���fF��y7e-�ْ���9�®
t��6c�g]��+D�H)��N_#�<\�����M�����j+Ë2�jFn��oV�,�'�0������9.�]�<c�m�����T�,�=؄ڗ!bT�
f�dⱒ��űe�7�H��y0��yw�k92��Ƚ9Ja����m�Қ���L�yw3H�-ˮ��י�S�7�)嬮�5��P0H)d�Q*�1Q�&��C�%�
�'��3�����'�����������;�7�oF�|Ŗ���'*�I�.�"�e��d�ƻ
Ã�Z�r�h���Y�7��Nż��^JT��rTٝ�UG-h/�8��M�F�-�]]͛:���X.�Eu�y1>H�JՃv�l̝��CP���\����m[�+xFIݕ�n��T�/T]Dn�Hݜ*����Sr��YM^���I��{}�K�������BZ1]s��V��{��R�������a�kZ��rҵ�"�Z�~��vQE�X-cڙ{��,+�l����������_1vU�̫7��\�&��Qӗݦ+|�n�Y�`��A�B��x�Ud��Y/��;i�/��
�8���gJ��܂�����{��c*�\",Vn��R�0��ָn"��MZ�YU����"�x��3��Ambٝ��hY ��c���@��Ku�&���%�z�ڣ��m�r�Q�	��N��g�:��x��u�i�����R�&E�B��RK|������a�8nT��P܁��˔�`��}�����$�{��;�r��B4�/ 
%3����d���Ơ77��@B�a�n�^�%ZINս�ګR�֝�	�\0�t��+_+̋�ʔ�WAt�����;E[��v%����ԩ�n��R�{.�#�j�B�e�͈�V�4w�l.d4����ˣ���|�-���A�ג��n@y�vwk4��vF��\���:�b�vm����J}oyj�o��l�ߜ��TS��h�j�{z��vo�����T���[�F�u��xI���F����2��T`�Գ�L�(���V�	WI^�#��'��0g	�\�Z'�
�>Q,���u`bݍ��� J��H�^jV�7���sf  �x�ϣFp%Ź,�o�hΧH8.X�zv�fp��S�ڂ��Z"����o5PѣL�	���Y��i&�j5+�[�b���Me�z���/T�q������ٔB5k���h��&���t��7�n�I�f�~wBFU[��3��1��Mt����Os3
A���.ъb�h*(�7�L��HU�]��S�����S,;�r�T��m4�R��X����N�c�N�h]����[�v�td���AΧ5����u%�ڗ�"_�*d�p؍J�ۯ%sB�B�;�)�swq�
�oogњ�gwzF��̜N|��*���:K�Ju`Ik�Ɯe>��sk]h���AЌ���Smo\�yn��8T��D�LD��V�$�l��;8gf�Y�TwvF�� �Okub����ٺp�l�Tt�{!Gvﰊ�$H�:�R��},�Tw,���u�հu}FvU�0r����?p�ғ#|橨dn�<�4`7�XR�j43�38�}��\�F���q��o[ͮ���'�HV�1r�u[r�)�K������+��l�Op����ڨ��ء�q�`"Х��$ѹ�r�u��z�e70i3G��쵴O��;n�>�t��Ѡ�z"k�٦.�,�&���[{���בh��tI/�0~�wG�7�WgX+��a��m}�<P��W"y���"�l9�q�*�ԗ+rU�F���>����]�9>�t�����u��l�ޮ2�	v��y�U�y�&�����j�d"�w^.��݆������k���s�:2��s����	+�/f�����j��i$*�_@B?9��]�������B�\��*��Qޝ�w�fbb���2�of���]BOh0[�����9;�CT�U���f��#��l�a6�Fq�I��)v��x>��Cy��MZ�PZ,�X64�NDX2�Fg�)ё5�ծ�\*˘����l٢WA٪���|����by���Nv�������3g���rZ�Ǯ�.3�L3,���E;�u,�̸�J@�tpL�p�n���vnp�X���:'|�r���r�x�X��%����æ-��m]��F�4�C_QIelQԬ�WZ�'���`�ƕ�g������mcu���1hE�etN�-��QB�Yܱ��C��q���#*��
F���NaNP<�;�ݩMS{~�w56ky��R�L��ur�&�����x��� �7ZG�#����r)3����Y�x$
հ�����Z
1cv6�pQ0��f�.���!���u�n��y��wNvɬұ�QR��i�8$&�KEt�)g��������(�ʼ�-C2�=�]T�
Aa���έ��GdVӅ+��!�G7j,O��*��+���T�w�+�X�W�55Zu����EV0����ʮ=6���J����jn�"�*���2JW��Q��SH�r�Ҭv�Q������:�v0������FF7�(��L�Q�v���B��&�r򻈃�c�<:��a��m�u)�N��S7`�;D��y�^4�v.����z�=�zk-Kh�]���"-(p�e���Ԝ��+��y�a�w�ҍ��0D�����)1��9n�wN�38}d�Tn�>�JC���D��2���q���)9��aW$�\���{�ץ:��l����a�&|�e��X��-���Yv�VUȍ�+:sJ������jʤ��\v�����-r���%����w��������fS
��-_`ֶ�~9ӹno��j,��]�|�,�5�=ɢb�,S�m�&vwa�3��[�@�MÁ�s��̕{B�E��r��E�2Aw��ѱ�.�j���.�<��WBlq�\}��S���*�U�,�7�v2v蜾TI��Ü�8��pUr��ձM�yc8@J��f�5�+1�Ei��Y�q��KfX�O9C%�����ڝrso���0��纯>k����PFҷ�|r�l&��t�4�;�ŵHV�������y�����Q���î���˖�Y����v��:�2��HBΫ�V��2��\헚ʜK���V�6�j{�Н���|0dN��[*}iu�ڈAZV��@��99��uY#y��j%ݴM,=yj91��9v��Ý�h��ͬ,lTt����#~ׂ�V��l���#r!C0�v�ҋ,��}c�f��CYYW�K�+j�*�����;��A�b_�WJ��FZ�T׆�,s���U��(���Dq�ؓ�x���kV3�m�����̅�cr]��`�y��q�mW]�&�z�hrMoo+X[�1V�ߛ��:�[��ߚ��!	 �XE��0��S�?�%]�>;����ds��^M�(-
c0)�f���l4�bE��Q�9��嵭m��x�oZ/9;�F\��8:q���v�'��	y��fh�;�]#v�RS0����Js)��t�ן^7K+:o]������ ˲��;T��s���즉�Xʷ_k���ż�L�����	 O_��U���VX���)�:�>|z���w-���&��h.i��in��,�;�Z�$�jN�u��X��b�d�;��r�����=�e������i��NI#%����޷�8�MzMț=�`):R��T�{����WM�P�Z�˗�<���;�U�P�eGܨ�ڧ��5-�����DIPīа�6˔��i�"�a�j�jU�*ތ��&
��k*�Q)m1�2��-[��Z"1/Z���e�+bKne#���T��Q���TU�I�QbƖ���5p��B��#hZ٤+���YJ�j"�1�ԵLZ*�Lq�&:�X[�q"���U��Zm��"�ɬl�d̪*5Te��m�m+D�,Ć���*�)�()�0kb�PXT1�\a���0XE�kJ�;�f��*���;��W?�L��Q���f1��kք�/�����&W!M�$��n�`��������%U�ݻz#�3��W���\��6֩�ZTw��6��v��@���}JKr���#]���I�x5��{R�b��Yw�����0KE�|Uڬrٷ�%꺽lp2���6ު���A��1�JF�zd�˫a�Gu�TR�Fs8���*�1�ԉ����M^j^�j�!����0�{mN�yd끬�W ��U�lnK{�&�{3/}Q>}����S�s-�=W���b��dP����R̵�V5phT��v�){#זЩ׳���ؖʽ5�� ����w�z�SJ����4bc\��K9H���-��y.�;�7c�G툺#.��X��?fn����:��Y��sBY�ڇr5\=��_P�R�']����}:�c�g7�_����[�h�����|�kD��e\|��d�,jIIidZ��͠)s���y���%V�(<C�V�oQ���w����a��:nw�\Bo0�\��U�(M
�o�C ��ʏ��������5��K�w�3ӥ>;�v؉�2�m�M�^�9"�U�+x8�nS���W���2��S�VS� [�4����ͥy���{b��j�����6r/%���h:�-�J�Y����R٨ٿ����')�m�*������W>ڝ�8�ߧUR���%����ê�OH�}r���RtE֏�c�<YY\�1�e��u��S�sL"k���|j�˘Y6FaKy=�\��e�	���}i�K2v���=S=kpW��ǰ�qҪk�:n?��i$X���&u��g.��W^� ˻�m7WݑԆō�7�cn�uj��e]�R\TR�ķ�[3��6��+2z�fx��`E.ꄚ�'m2�q�4����8x%/��5y$N<T�@��5�:zv�ƛ~���O����L&�:��2���""#1>�A�qO�ͽѷUv���\����i-F\c�'j��8���{J����N�Fξ��;f�>�k��͚�i�:	�J��-��6t�^l^��c+;{��cb��6�z5�k���"�����R�a^u��B�y�"��[��zlUm���dIU���%���q�ɰC~��5o���E�W<���D���c��$њj8�ߵ�
E�)�n[{��{�4���7;�F�<�k��"O:睙L�CϔF.��y[ϋ��=��O9��z_��n��6ܨ�Mj�:T
{�͹����˧GU���gB�RYRkM䖪|8O�[��MC�	�qi:��?#E�m_���ss̫��;�k�����yi���<Rށ�;����G��إ�r7��:����*?p���h�#���pż�tk��emHs��q��&B�T��CZr�trZ�n&�r_d�~�ϬI��U˰P �Dd&�竹k�*�k:ĉ�74��+~[��\��G�mr�9`{��.�ЮYG���(��<��j���dѫ�ؠa�s��E6���������>�,�=�+=����ki4�Z������ϑP�Qa�!=��@�䷑���2	�8��qJ�z���Vמ �p�Qj3�dY�S�^����f��p�M�w�L�¯�������<S%��{�{'^����[�a���1rƃy�֥[��
�W��㒡"��{i�Z��OiW�"D�$w�ǧ��I�GW�k���a˭�W:�D�@��/��3� �K�4޵�25�H�B�C�'NF�:���ӥ�'�[�I�މ���t���+�<�.���>��T���t�R�T��J!Ҕw��E���e��+� ���&����7��zO�z`9�n@Z{4d5t��g����gpu-ķB9^�7V���Qݺ۵��=�E��>���ck�ְ�+���"�D�-�e�ٳ\�Yp�����URPe��:	w�y��T�$[Eg'���!�S|��Y�+iF����t��6󖷵9�/6\�)�ŵ}WD1��hwj7_NtH�F���!c�Ŀ7չ�y��ʋ�a���%�Q�~s�c�����|�Z��Z7�����zM��u�g름m��%�G�=�S��ө��ge�=��s5��K|8u���vۣ�����b����0�����'��r_C9>�NyF�e���]/pG[C$ѣ��|~:_	[\�dqt�
�i'��3�s�T�֪Y;�FdnU�ܑ��8	;Q��[�x�᱘}��� t3�>ӧ�nw�.�h�f�5�kc�҄)�O�z��vlէ��L�WÅN�o��cDg;�޺	���h�Fgci���ꙥV��@�^i�|E��/^�3i�lV�M�l]�O��s���:2�7�a���Y��:�)�yH�5����,�&�՗ј*>�ݤ����f��P5�G+BYHzM3m�M zb��;��gv�B��Ք53�)e�L盿+~0P��z�-J���pj�Z'u��r�����;�	�ԑI�x�a!f����+�\[S>�c�c�-�ˆV#���Tc���ݘ�!��������T��/ݞj�)9�4��AJ���(fT�#��F���^�]jyN�<u�Ӓ����c'n���v�Qֵ��6KS��_pu�Q��ӯ��)�z��ȟB���vqe`���D�L����ӭ͹<zk��N7�%==3��K��;d[<?^~�Q��H��0�p�~� ~U����Ux{MMŴKT�J�@��d�m��Fe!�Z:�vw�J�Hu��V��;��E�����fu9;�pu�C�Vs���t��8���4����/$��i���MPp�����s�3�oY��R����J.�˸z�V�ˌR�T��^�!��Lb�YWT[�D:M>2�p�/��;9F���D�b��ⶨ�v/�����;�
N��9���»oX��ľ�c�kF�]
�f�cL\��P�����eg�3v�&C���5�Աu�w�a�r����zv�;v2k_5�0��*�'3�:דL�7�O���#i%�hά��[����1���"��в&�)h���u���F1��y�hG_��9�C��żj1�2s� ʹ��V�5�:���!�x��������<��0��Q�]��c��J���i�,K�����o+v����C�:d��N»t�Ll�V�c���[pYx1\9t�w��o��X�J��|tQ|��{_&H�����/� Pr����2|��CI��
ٍ��xԂ�0�9b�՜�TT]n����t��Ai�;��-�hv�lQ�3GC������T���Y�Q��%���p�Ҍ�䌗$rJ	�ob��ڒnD]�O�aV�y.Y�����8Q�*�h뭣�d�x�1��o�@έTe`��,QC�L(�2i��Ye@�F&�Z�EuL\ma�D��.!���;q2ҤPPR�UR(�Z.�&2b)*[@XM��
��Lc��E�ua��B��d�T*��%T�JͰS1Q4�W,��i�db�04�N0��+ �r�1
�ʢ�*Ѕ2�@�(�+%Vc����t��.���U
�� xL�߾?(��;�5�y լ��NC�~�� ����M���:�p+���s�@p�4�5KK��"�ͼ���5�-�:~�������B�ٺg~l�%�3���R������G�gq��a�b���W���c��GۘTf��Vj�V���F�#(�y��x�%�H�V��1�w�q�y�4�ye��tx~6��j�Q
����I�f�
Gs<K��+޶�1φ
oA��'���Ɔ@yTN�L�ݮ��D��%T��}"x�:��jn��߀�^u�M�o��<$k��Q_W-�:��
7ίG%d�$���>��t3���T(���@gZ�\f ������탫��d�U�8��R6�Lҗ7��o-Yz��ą�%���0{�k҇{�
*l��m������s*7����V�ïl�x��"b%��S>A>�~Q�����R���m^N��P��<�}�l�JD�xW�I+�wI��W��	�W#-DQ5�w��Q[����%��%��q���|�lf�9w�~�~S/��sv'��ڢ2C��]�f�p�j6��u%Fmb�j|U�K�^������qLk�a����q��1�O�J��sf�9����Æ%)��)�?
s�Ⱥ��M�DdV���1�C�픚�5�'TmpM��0qݐ�'�u��cytŨ�!�.|��!�ML��#HW�2�����&���k�����<��)�̅l��f���
R<G�o�r�\�u�9�By`z�H����s	a�x�`�m!�I�&2Cya�`z�x�<����[�.ߵ�W�^��� �K\ʤ&�XZ��d|zk̫7��|�Y���|oK(���-�J���P�K��B
Ҋ���)~�� \�O�B��Cz�I�Ї�'l�BJ����t�$��o5�������f��!R2@����P�0�$�k�$�Rq�g��'�v�tá$��������^��OXVm$+�<d=d�	���=M���<Bq4{a<f�jr�r�q	�{�9�~�I�$8�
�Їɦ$RbE���|�6���$�u�<<�|�>�<d�!�,�����4����'v
@�>H��C�RC�OP�@�]�����]�;I8���{�����;I�	4����x�;a�P�J�� z���̹�}��2O|�!�(q��{@<d��q��$1��O���01�<J}CL��z�wֽ���!�!��IYP�$4��`zyHz�g)'��%B��;�v�Vi1g�<��7��Hc!��=H�I�i�:��uOXC�
@<d�(A�yG���Ҿ��'mo'�Txx\ <z�g���!P���C�5���v�P�3x�v�x��x���������:q�.�R��s-�]�����Vl3{�����]M��w^�X�V�	�N�I�c�'+vr>�q����!�!�~:I��v�t��*@�����C�s�@���3]S��5z��{�y�M$��8��Ho��@1$���I�+e��!�&��=}���<#ۋ�įY������2wN�<I5;�N$��I��N�	�m���/�2L5��������﮻	�O�H0�tæq���X$�2v�:d'�턬
�6�ɻ�]}�����}�d��t=`,�'�8�kt��=��@ά�a���6�Đ��2�2T{��s3��������d����!� o�!�'�kvC��a��!�x�i'���æI�y�}o<޼�<$=<d6��l
�m'��,��e��@Ϩq��C[�g�l�����	޻����N����y���n��G�� ����!�g�!�3V�q��ϼ{®G��=]��ֵ{�)��O@+&Ϭ���a'l�v�LЇ�� ̰�@��vu�o�f��~�0>IĊHm=a<@����d8����P'v�q$�'i�>W������C.n���_�tP�#R<��:A�,��D������+5
:�h��>�Q�)Z׼*M����As��Ǌ�x	{��0=���z`\�x��d�$�M��=`x�xι@<I��>X
I�'Hu�9�y�5���4��	8�3&��t'̆�=a��Cl�!�Cg�
����L��Bs�o���z�������'l� `�t��N2uI큌���� Xv�
vn�!�`,3y��W���<랐Rz��H{ߘ��C'hC�I1�d��|�v��B��b0�'��o�7ۯ��)����@ (���{�Jɝ�!Y:I�$�	�	�)�4�8�|�w������{���ܲ��z�Y�X$��L��h��Iq�x� \{����������9��!�yd�К:���H�=a���'�8�x��I�t�`s���ɜ߻��{ ��H6��IS�!�f��$�Y!z��0����	�N�$��$:�k������\'l%gJ��!�5��&�|�1'l>Bvn�<C=��I��C��$�'|���k�w�$����$필�d<d����a����!�&��v�_RCӾ���v}�뫮s�������~�۵���*P�8�Z�6bѴ�~��bVz�b��׆���p���5	g$l��˒)~
�٭���i�s��&���)$�!�I�I'I�,��e��@�!�Y��ïpNx�ȎP���C�뾞�xe����i�佘Vy��'�enӊ���.v p�O#c�t�L���B��˃�tÖ�qZ
��Rh��]�v�V��}��û��h�H����niK���T�ZXՂy�e����f�3��Ѱ�w�M!�P�5֧���X�Z�,��F���Ov�*L㐶lx�B����f�e =��������q���)O���%^�G��^�p��r���:���ص5=���5�)W�����O5��=�����[h�['�����5u`������o��?��J7�ٷ៥V�\��:��>��������۬5����BT(��Q]�v��������I�"5�ρ\p��畫��x���h[ՏU9�tv�˰y��\iR�h���P�v����*j��.6�\T��[Y̾+�/�&"AMj:�״�x���ԥ��5�v��{^��IHOo{K뷇��T��y�}�>J��X��ȏ���߻��Kxa�|kk��9����W�5H�nu�KJ:R��{���]O뾑�����}�{A�be�� {E�]mH�'eq����=7����ދd28�;�V��ֹ��1�׹[�p51˖ S�1���������p�:�,�R�X������N)�vC�Գ��%`���F���c��gs�Vkʀ4*Fx#�!9\Z>�]x+"�1&�_u+�]��]��Q̂�Q�F����|�D��(�`.vbs�O�t�n�m��=��a�V��#ʔz�z��FX.M��O1at�7�!�H�!5��"�燽�x)׺�?�mfX��
dA=�g�� [���b��%�w>�yl��W��6���o���]L��������~��̄Cs�����N�g䳊�Ԑ��j��=�Ȑ��dK'\���\�OT�:����٢�mi�E�� ��_��Q��\s׻�ǘ,1N��Os+w�N1c��2�[YGW��,��o�E��G�鬣�AV����n6��������v]dy�v���p��<R��z� �:�*��x���bap��MwX�2gf	���T��ٲ�)���IZ����Ύ�h��h:�u���p�w�p*Bgk�:į4v�A�*о�Z��&h@�F��X/k;�q[�X����J�F�����1L�z_M��G\U�����t�h���5�4�=�fl��1���u�`K|4���ٮåƮ�����\k��0�bХ彺��q��˻�	Eḽ2<xc6\��Z��.7�]���KF@%��4sc�ͩЬ��:r�z��W�9�
�|E���nFR��M��w��Vc5uqP�.�Z͆��4pVR پ�x�͊ݫQ{?��σ���1����f����N�Ub�GcM�k���>��^�k��m��+���+K�2��#�V�0�}Z.��}��!�ڳDf�����a:����gu�Q9�b��t��X/���Kx�Ǜ�e� 4ٲ���R�FCe�SU��;GA���bs���4�m���w�9�^V�ǍN��W�����%<2�ܷOs�k�i-w]PG���%�x7e���W���br�[#QB������ �@M�4+S�[N��K������������t�}�4W��"d�H!H5%�R(�nI��:/��
�TNN�;{�+��Δ���x���c��}������T8ԟ!b�b��)h�E�dY��i����$1H�!�V�1�I+X,aD`M2cr�(��B�ղKl"��P�CHh6�b��Һ�f&�DE�UB"*cT���b�Ȉ�d��RT!�b�H� V	mV9�H*�,HbT�őA�±`�X�,\k%`��H�(��ŐTJ�I�LIF
*���:���"w�̍
pQ�o����ӓ\,HMbD�K����x �������[�vf�U�#Z§�}�D�f�}޽�
��xK��{:�_��.������c�@�)�����%�L�U����T��,;��s%)Od�ͣ3O+��^<�H��h��w��M�c�pa���b�2���a^mrtŮ������u�z0�b�h�=Y}Ȓ��Rb_<��Y
h�
WR�WN3��o��ThK�wM��5��ף^�A\ş�ެ�~�/�tR��B;��ռ$�g�i`���{�:��Y{ӯ��y�n�J6֕hE�����	�{��p��~��Z3��+y�w7<��K����-99��i�w8Foa����fk�¡�y\/Lt���U��;�;*�8�z/hx½�ߩ��e�A#&�o �>�;�;�]V ~<ai���=���e4��*���gtS��X\Lǘ$$��7�h�<�v];/�'`<�k�r+�zY�Co�n�Fomkڛ�ÏB�8 ��z�U���ڗ�q��A5�=0b�TgY�)r�H@��,�d��45͞��|+Rx�l��pf	���.k�E%��  �V������t'�;rʻ���X5B�T�6�b�k;��+:�0#��N����<�G4G�=��)h�\�A{�_1�,"b��7��1H�h�����+�48���c��x$���+��OKR8s<I��9Ůj�̘jMu[ދ�8����m F��>���n�hf�J�3�u��W���kї���;}�M�zu���ԣ�ۢ//�L�H�<n����c����K�41*�tΥ��1/\�d�15�����0�6#4��쑼�¹�{�)%�W!l&����{�D��zU���moW�{m��ڕr�}��*����3��Y) �F�� �m�jFmi�@�|���:������G�>�<�g��=�½��'����}}�y%g�~�SX.ߎE��2;I��q����y�<���.×�%����hdLV4���p_��x$w��/%䜐�������ܣ6z��Y�˶l�X������r�i��{����O����} �û�᧱زLt��Ӳ��C��k]�/�^b�"/E/}�x{��Kǩ,�����60àO�a��9e�r�CB�x�\�ohlë��ɐ��a������xA�
��[��hU�Z��V�o����ߢ��� �3��c���B�϶��0�Dn<�ba{��7�fDc�ҝ{e.��MC딓]���7�]�����YMF�W���D�/k~��!�ݝS��?.P�#y���VP���]z�W��o�\��#\�P!��u��Gܐ�8�F�Z��L�q��3U��C�P�Jt�C.u�\����t�B�#į�� ��e�z����Z���V~l>�l�2��o��N�!3�c��Е���/D�e�r��<����2sY�r��yֺ�B��O�Oy ����xv�e����C���E�����╎������ָ�=U.�or��03V( �7��5�+�O�����3�z{�$��	�/3 ���f����G��$���K)j�>���*���V���/5'�����Y#z�M� yyQ�eZ|xQ�Ή�ƻ�+R�ЬZ]�j�J+Q(E�RD��=�{��wݟnu3[~�د�Чs(у�d,#��� ����|��K�ˮ����@�h���q^d^w"T��4$�u.Q4/kp޳5����Kl��f佴y��Л/ʥ�����I�^F|�P��9��s{k�!%��*x@�:��65U���">�年��Wr��a��|�0��f���-޳Q��:�U��U���rY�˔;���%{��U�C&��P��f�7����o��Vw�w>�<�mn��<�Y��{�ּN��6v��4\�࣎I��x��ZW�MI�[ދ��y]	
U=��Np!�����#M١< �����S�v�\�ױҧ�_T�uM�������9�Ǝv4��{z��6�����WJ�[���K�ؚ2�q�G4e���/w�J�|�ӢA�g��Zko;��⦝�S�{0f�خKx�r3����wQ��x��R߼�>l��cY]{�TQ�ـ��R��w5�U��p�Lw���^ڨ*�2���'F��8:�9\/��]��!�$V
��	(#��R������בB�>V_eN~Y熬�E���$�WR��-����i���9��j�u��#y��y�>�V���M�[o47V�1��;G��7%���w7ʲ��+���3�4�&S?3k�<�y�!\�g�j��W)�k&C�1�������u�Vp���muu��O�.�>�Ԉ��pٳn�i�b�+�tFs;���GO��VA�*VG�q�����v�N�;�#:Ywf��z8#���#F;��N�Q�Z;5gZ%!�%��}W�Âpr�D�$�H�����g>{�@��d��,P^~xC���~2��]�/<��=���٣��8׹}�Y����,4$�M�������l��dQ塚)�O�fɍ�t���k�E��>�Q�=V��hx��[�:l1���f���:�"6դ(�����N�>(������V�݇ǈ�g�W2q����!�@욑�2%����gݳ�"Dle:�Ԉ��	�_t++[�Q��ϒ�o,��]���L� ���/_���U�?<�3�8i/��_B(�a�U�f^���7�	���L#���� ��A��>�>�����e�b4�͞�Bz{Q��|�[�k7{�Zޫ�2�P�цas[T�e���u��Ru�c�u�if5х�/�� dY�S+����4~2�l���a���{:!y��j��l��v'��z&���m[̲j������0�-ͲU�#�\�ν'O ����Zju�`�X�޿t�55���dD$�����:e,���8rE�N��d�u��{��9cm�K�oM������SN�V�ݷ}���c��QRR]^Emjn!\dR�=棙�t�o6w��B�<˝>�k]>�J���&�#�P
��y4��h����W}M��h�q��mꇙ��l��l`�Kbե�AԶ��ת�>^����Н���kJ�*fd��t�]�G��Ԅe�ٕt0i��L��$�w�V	������E��,�wmJ�3��Φ�8���,�d��v����5�1A;�\��*�
7��6��I�ŗg���L�Ʀat����h��!����Y�����3#�y�)È�;t�XY�݊��=L�����]�m,ݾ�.��3
��`c����B�b����5�;�Ż"J�%ꢘ[�p2���[��rm���ط8�>X�Xb��q.Q(�D�"c�d�#M�$�l6�1���Fd����]�Cn4��f���7���c��gL>CZ��ő`�
H��XV
AE�UH)-�*�j
��R��2EPPPU ���J��d�,���"�YR
EDd�Bi(�

��
`��c Ua�$� R

EQLM$1"����QH,YH)J"�����~�	'Ͳ�f�{7�������P̤Qҗ�=� x�5��>�_P�΢~��b��)����$�V����~FȲ/G��c�7�WJ��w��r�.CK �~n�i��[���3/G����LUI�K*m{k����	�ߝ���:���]���p��������9�t��b�P�v��,vR���H�Q���x�_7��c���?Q�ԕT�Z�^��~�+��gH�5�q��L�q���.��3�@H�Fn=�T7$�raZr��i�i�nՑf���!��-xh���5��kוh^���!D���$f��>�Ǐ�͡��r?D:�~�4�΅���o 
��S�&2uה7��,S! ]��e嬇R<9VE�8�Ed�D�K	]�F�(�+�x{�]��W.>R�W��Q0
�

�p�Q�3���e=40Z�b/�1x�&~ô��g����;8�	cS��`�5�K�Y�^c�O.��q�Z��'\��:��:E^4��
��Ǘ��ux���T�;�ۯ����

�8D�~3�C�����L�>�ͧ@�,8A��"b�~Ve&\P��]n=��>�D�_q���3�E��VBm��I��*uޱZ���x�.��1x���C�FK���<��^
"�E���դ+���o&E.o]gb8~�V]�>�����t�<���Ǯ/!t�u��f�A)���fVlpgs��Si��\-��u��,��О������p\ �[�G�P�:�%/��+���}7"��P4*:">��܂���1�X{*�Wl�XFj�����6ř�<x��ӹ!��{ݑ}��!SV}:O�()�dB�^Y}��i��?x�����:E�4�?U���i��:$�g�q����a�#H�d��b��{6����r��a���"G���G|����Ş��N�t�����V�GR>4)a�[��>�1қ{y���!ld�h!���l�<U�|��S�h!˞���C�P�_u�:����t�+��=y�m^!�I�2B���F�8n/�����˞�'Nѽ�ʷɃ0�h�9�U���]䮒|Wr��l��-��[c����u*�(��+:6x�_xC��{�횋�_H���u�㼑��$h�_�0�lq��|5p�gH���Cp߭l����!G�O�j��E�����I*�g!^g=��Y��,�1��b�0�-}]#t!�t��'&����^׷f�D{^l��a���HL���1���/E>��,�_	hx��O�m^��W�(�0���D3ֆz���B��kM���5�[�N�s�Bf�Х-ʌ*.l�7��b�Õ��O^�jv~d�#�k��5g7X'N�g����g!�Y0�#M�5��쁩=�6��x֧�!0���󗪖l|�{k��^��ϭz�eGg����ػ���{�
��WMŪb*J�(�$�H�� S��o/�D���=���M(5���'�!�09	h�7�Q=#��P���"�D�d�������cwvފ �vGF���$l�_#X���\��uך��Y�K��N�k�N�b'O��f�<�I��fn��K��+hp���1^C��'�#���n��xI�<~Er�*v`�<r�>�1h!�OU���J�˴<G��<Y�YE[�R�7{�R�L�J��G<��c�!{O�6A��W�dU���������_p�~3�����d,X��ܭ�{lϼG5܍!����a�/�*#چj��/�1��X�{S�Ӿײ��o���`W�O@-]��<��v-�o�HxgI{ϖ9�I�7�+͊�%p�G5��K�x{����Lp�l	�R�F���A/���x��)Q�"`td\ ���㺀�l[����5+V��ޗƵka��dY�g��k��#�#��[��{r���s-�S�!�%���$g��rؒ���{~�����C8t�6}ό�2������89�YhxT���9[3o]�L��[��|s�jn�Η/�����V�Ƶ$/Q��kX#�~��;sP�KVY��>"�I�)/ˈ;;�+s�d��>T��GyY��x�k�)1�J�bi�{��ڼ> ���;AC��T����;��n��Q�S�>[���F�����óm\���V]W-�6�em'2r��̦Z����4�����]ڋ���~��]{`�ݲO\���y:�q�7v��g
c�A�/�<\zs��yцa,��U\��KK��> KT�����@?&F����ۺl�,�]�j����~�熇��x����X(�-B	{�ư��c��5��Idh�y��K��=�'��!�Pط!F��gs�qk�^ה0�l��Ȣ!�Udde�M��~�8Ta�׏�� -VsV��m��F����}�T�ğt�jΌ2����q2{n��d�?	�pa�x��#
��QA�*{S|�_�JNW鼇�s��h�aB����}��f�	U�\�'y0��:���-��v�&�
�~�0�R��&��ȥ���S�Ih���r��m|�$/)a��܃��unm_�t��!���Hv� NL���b!����=y�0��J�c�Uy_>"��*й�b�}w7�i��3ӄ�2B_^k���V��b�ya�C�,��y�8G�bӟ.��n��R��(=�M_\C��v���i#�ۧ�e���x�8D#N�ii�->8-x�b���[��՗�38p�g�mp�!O�i�Z�0�yo.�/�/g�؄��,�\�� �E����蛫W�޷�{P�N�k���PGH��|,�����W{wj���S��ck]l*��;��	��t�:�=�tX���@��m%���OV��쏃CQSe^�E���h�	[����⾵jʑ#d\}���a�7���ۮ�k9!�G�$��v�զώ}�h!�7��i���)k�̄�ǲ,L� ��qQ�ܶ�L�1�ohWZ�k�p�����4Ѳ;Q9v@ԉ��V$=u~�c��D#_/k���d�DY��� ��Y�=��J��#��{�?M�őRȆ��1n˼��Tl�A�=?=�iZ�$�1[��3'V��<l��@��{�"(ȉ�f<�� Áf��e"�tk����B��B�hmy�����vm�f=h���J��4��!�S�ӟ��]�s��k�`}������j*_YT�瀈�=YkܗX՘�v���/�a�#��zse��N�z��7?}T�Uw�W@F����i�/��M2oƳ�/9��᭙H
��S�A���4P�
_[�q�z��8l�g�^�*0=�������1-��8��Dk9Laㆅ�~X�������������FX�"|�j���3�s_���<���=X��G�E�6m '-�֛��oC ���˒!�Lc�}�Tl�@���\x�X]~��^���C��|���!�_](��<����߲��Ծl�/VΞ-��\x���A�ʳ~�J��E%@�t��b�yi����u/��> s=�@����iwi��*�Kz�M�V8�6�f�m;b�wVMu�Э�S6�5ˏ3��JZQX�gqs��u�!u�.�I��v��Sm�I���*4��oK9R�m�'P��5|�t���ZNu�]Ԣ'[����A<�)gF��$wĦ*9�Tw����&�v�Ktœy��U��sS{v�[$Ȉ�,&�]���	X��F�lEuΚ�3�lr��p���np� l����&��aN��p���8�������dY��+�����M�p����sg7f��n���y�[6�@���.%w��b����&�A�$��;.9J�/� �n[=|����[{��{���n{�Kq���2̐gd'�r��qa֐k1��7lH�3ȋ��Bǥ�c5�G�ӽ�0�f�f�L���#��uoMS$��e�w�;C�`�E�ܢ0-�1LW�K���^ j<��V��i,t�����]���뫁������宆��W��L����mfuێSX��Ab���!s�n�ld��V��MD�[��$�j�Euk���т����ht6+����Ƿ��Vy:�&$A3�vS��
���șU�S�:�]m	���6M,��!kc�1(�R4�rI03%�#�&ےo��{�v�
a�j^�|ޕ2�s~v��<��׏<�g��,P
��IR
EPbőuh
�Ȣ�)J��c��&+���Y+X
��B֓H��6��XQ�acj,�5��TĨVAkE�bTQd*�e�K�&$�
v�)3v��&&&*+j˫���ۣ��x�����nV�u8�nw	㼆MrI$�or�k����jʡ�G�.#�����yt�X�J��4���'~��C�6l�[ E�/J���R��GT��z�dv���a�#M������=��R�&�ϫ�:�zFǎrWdV �$_�����߶��Nr��z�{�F׺|�k"`�	۶��!�f�2�(r�Q�GB�f��j��l�T�gc��Y ���@PԘ6r��W���6k<zF�չH��4a����t�����?R����U���y���;i��#�P�E��'�}��4cy��炀`VO\��@��rQ���0����b����O�װ~r3����Z:��\4��jO��s�fo�pMꗘn��(�>jh;7z�o��Y�r�nO��}y��w��i�3�E�!Y����Ȣ�?JIN׎���#1Z���e>8w��ç���%_��GE�xy-0�<���������rC:�sH㤥G����_���HĩE���e��	w�l_�.G9:=vb�]���~�1Zy��"���%���Fp�G�6`#�t�%��c�^!�����ɍ��b�(���V������#؝!� K�3��/����-\�IUپ�o��Z�p��nG@� ���QU1��y��ƾ���Ɵ���9p�gH���� yix���f` owc���m�u#���h��(��wW�t�kwwҼme׫���g%+Ɇ�ӕّ^	�lxx�)~xz1�ԣ�d1�H����B��Fl� çh���W [�
,yB���N�$%O�i�lV��s��^.�v�"ȇq����v��L�~���~T�4����6�٢;ˎ�a�覯��:���:��O7��#慹p�>,�Ü��!�Cn��ǹ��gR���6a��WwW2�����v;7^�s� �E$(��(���"��B�6s����>z�$bpEf���YO�e���g���Y9�DkC�_��u��FbKZ���f��4h�5>��q��������C��:�	uS>(H��\�O'8��ף� Sn�S���=j�2=s��6�������w_����Ǳ��F�"gԮsz1!W�į��T�^���ň�������-.��͜1/���3ӛ���s�cU�w&��DO��8�'I�\��۸*׎?R\3X��Q
?P�1^B����{rZ�O0�D�H ~F���S�Rr�<;�=��5m_dc�*��SP�+P����ƙBǇ�,��wSj�H
�ڠ�1��!{L3F�>���5<����U醭it������ִ���,A��$O{}���%��:C5h�8ߖ�(y|�Q6��f_���=�-/�(���#`e�9P��ge�M��>���H�|E�����;�����u\>;l��c}�J�]�;�m(�⏢�}�"�ۖ�.��n�T �(�i�"U�$�.B,����	o7[��׾B\f�_sv+6l�?�0����{�^�x�}G��R�EG��oʍ�@�v}�6&GWc�g�>]�B�ϨC�<aA �P��h�9�Q#o+?w�-C��_`��⍑�R��{Cg��=d�W��[��q�q�v�k;��������s�,۱f��wb�\
�34����i:gVrYC!>#	���t�6D?$���ּd�j�����a�;)�oH~\^�,rk��0���;�a���� �j��}x�Ώ�#k�|�k"�Y�̼��ls��8Ȩ�T+�B�Y,9
n��m��jd[S�ӎ8h�7�K�9��CDT�v��c�\�e��d�IYA�<+��U�hs�k����͊`��YYȤ���S����@�3>�ddt�G�f��PΠvzi��6�)�)����\y޽.k�)�Ń�n�It��K�=�k�O�ô�P�a��9�p�ؾ������_�B��^ �^�Q�ia���S�JʯJ�6(��i�S�_��͜�YQ������}lrꌃhOy�txcZx�����-ͮ�,�,���餟�H���ւ.eiǛ{��Y�p��yXa�f�9H��\s��|�k;)��*��=�a���8j��-Hx��^���Ԝ�Β�ql1k�<t�!�Q"ȬTY�ś5�,I��+�u�g�(��)�v�M��z�"�6J���3H��WGL}����ggQ<����2 �Fvh�Iո�E�����>و5�#'���L��H���l��ܫ����"ʵ�d@�<���^2G�5�#=�����gM�#��<8Q���E_��\k��Ny�e�s�r>��%��e[b����c��p�mm磱�y7����ᘀg��;G�9i�6���F�S"׽Y�9��`V�:w�?j�$R��+�u5Q��u�qqG�.����s�i�Q@����mެ�h��<'=4F�?35�<с��2p����s�!2UHUj�8p琲!����cM8nu�w�4��g���ǖr�V�������U�We����hM�<�͞U��3��@k����D�4�[xD�tH!�:��u��L���b��I:�K�#^��r-O�U
ʠc���g.�vVcFOja��O2[�yb����qF�6G-d�Ȥ=�{s2��}�=�R��X�G��1��f2El��FM�V��Ҙ��ii����o���/�=�u혨�Z��Ab����C���G��^ٜr��
��"��a�=�`� מ�#����{��e�'ƈ�Z|p�I|�
��D%/��	\�w�-�����"U ��#����u5��e��E�Ca���S�<B�4�/�����"��ˈ��vh��E��j�3<�,m?�Կo'��
<��>`�Wr�g�ml\^T���؊㪇�>��$�^K�U��Z���j�5[H��H��/�V=b�G��t|~�j�[�l�v�T��w�wx��
A�b_���"5V��0��W�1���C1��-���X}a��3Z��x�
S�w�ݧC-}dg��(�����n6[�M�y�ݿWO�!QfHJ\Y��uB�t���Ԇ}�����E�G�C��<�,"�E��/x�Y�w�v1FZ~@����(��ӧ�P�g�9���`��� ]:�˟��=3ɖñ��X����"|~/��]��q��<�s��3}}h����?x�_C��Y�`���^$�u!��;�7Žyq���QʶkO�̱S��=�Q�T{�[�Vv���Awn3�,���^���A.����E��X���ʬ��߽T0�8G�ߑ��6�4���|E�T�+^�[�a�����p!eE$
��;C���N�.�;ˍYd���~���S�~7L�2�jM�1]y,!�"�]!��!�!C���1WY���b��6u&B"����?U�HAX��P�ޙY�u�ڀz���h��LQ��T����g���o�����,�����4|��p��u�z�����#*��C�谋�� ��*�<{�^��jddl�`߲�:��11��߅m�b�f��W�=gH����.a�׆�=֗姢�X������0i^_��$9��Tb5��N顾��\na�s/a��iC�S���DP��(������X��W7Yf�U���;4�ʱ9Z#��N n�8#F�m����k �6`4'v�/�,Ә�Y������;'N�Sp�W�.�S�e��ORx�SŨ�$�Yn�57�n�m	ϑ;�{:��b�gN��(�Fl���n���w٦��噉jŕ�k����el�7�u���2i�F�DbI
0�+��-Y90,s�ō�.q8W����K&e1�Fk���^�lݔ(�;��os�>�׊dǻ��sX��`��r[��P��2�9��,W�g}¤��Y�U���.�.�m*Ze��u�2Q1�#͛�^�2����7H]��o{��u�`l��Z��������U�9�M�V����gih6n�N)v��O&�}J�n!A�����QsF�f#q�}#wu�BQ�b�ť+ ���؈������֛�r#�k�K-Yt3�iN]��Ŋ� ,7�}�h$8:�s>��sd�#f�<ϑW��	����`�v�DѴ�f6*��<ʦrq��)#�jJ�*�ׂ�f)�vw��9��:3�WY��m��s{���M��4��&�2rÕ��<:#" ʧ�|a�q�8�Q��Q�$�$�v�1�\nI3�b��V�QtSY���oK�3igJ�[��!ho.�}�ỷ�yG� ����WLkISl�1��0&[&2�nP̻C2�V�U���X�f0�m���*��b\�X���˃��X,�ɴ*jЮ����q20m����H�kq��
�9@ik"��4Y����@D1����̢Ԯ�Uq��m�(�"�11��d�x�g��KJߓV_]8�m���X60.�g���d�I�UNy��g���E#*t�\\ZC�w��=fُ���1��x���R��#U�P��ȭ!��_�%{�׏�2�y.B��ӧ�r�a|Rԇ���o�Fxb�p�<~�Z|FP:�Fh��>���_<F�-�<�5�qz�1�����t�����[��d(���8�hs�|��D����VN,��mϬ�4���g�.!<�8B�1渄�I������GOԗ�>�w �������yw;��'�q֚��!�h���>99��i9W���x�a��Z��Zx�"v�HL���:��������W��8��fg{oAYc��ZՎ,�[��/�M]E��S�6�k8�+, ����������^Ө���p/$�',?Y�W>��$�]��jUo�S�<&0�)���y�:]���-�O���!����T'�"�fǱ��8���z�0x�_0͛k��_b	y��B�raqÂX��ϯG@&_��dȷ=Ȉ�
 ;1��<S����Y�1��*d��sQ] �J7�`���Qw�͕~�h���c���#��������A�6ܝj���ϱ?`>#ǎ�ü����ǙW/�׶������iq��{]�wJ�ۣ��5�OZ*/f�`�
4{��|o�k����u��JԸT@��\̥�x	����rv��d��n�b��	BJ٭e�+e.��/,��Z�\v�=%mc�o�^&$Q/��"��oFG�1�J��b`mM@�������>�g.�=e3�CЮ�3�8I�Y�Hx�?~�zt�߶��i��]�(b�C�0�)�!jY[2fI�x{_o(10+d���3����:��pr}�`����3�X�kV�K�?������9���Π�z�����S>s�S�1c(t(����5�m�y�Y��B���:F�`#HMV�uq��Y�۱P��bZ���wL ��"ֶm (����U���i8zkK��DQ�g��ꭾ�7��锆�~:�X�LB�KB��a;���W�m�uK�7�D��m��͘�q���O��v%�����=-�y�k�T�ݪ4��r���'��Ֆ��l�L�C(lU��M��}
<aD�?I����{k}���6���3"�_c�L�dTr�+�́�K��O_	J D��%^C��b�EJ��we�O�b~���:k�F����UW�y�����E#�O��H�g�lNC��I]UR��遵9 �����
�0�C��2��P�}(�E�wW�x�{�F����}禝d��4�^#�I���1��!w�0��7�=�����цaG����Fj��W�T�pM��9���r�_HN�*6�?z��.k񔆂}����y^Q���Onܝ�2�c�'<���WOoD�3�k���D��΄�Qs39���ё8
V�W���K��s�s�Z�K�y"�;�H��B��U�e�I������d;[A}��Gifi>����$B	L1ˎ�ON�+�4����9���^�أ���d��v�4@��kK���d��jM�^��j�X#��1Κb\\ZCB�{��
T�C>�S����;ڷ�7�e3򳔫�ײ��}��Ằ�E9	MҠT�=q�=B|�����=k�����5�O��Y!�h���=��6+<aP�N=aK�N��`"�S�y1Q�Y�p�\��4f�p���T�8Md����nܢjz�t]��0E�Wb�j҈魫
ڎ�*�3�T��oX�xi�=:�R�t\Xӊ��(M-K�K��=ǭo������?�����ᘙ�?!�X�1�3�_�c7�꼇,�PӜ��Ak�"ʴ4�T�{%�u���XI_R�GgH�Ƅ"��'�7;)5��_Z�������gN�B���VA�G:�g]��GIj��B�j<��g]\�Zf�"�mu9Q�G�vD��0�rj�ؕ�oׯ�wH�����)�ㅛ6s��N2i>]�C}C���ޙ�E9�&6\�b1���F�fp3C%	�QA*!� ��Y9H��k}Z4��=2�'N����7���#M �`��B�e��Wջ�+�R���
��.��.c3RW�����7�}�S-Zٱ{k�L��p]���ԟxxD��y�@f #�z�}S�F�j��c&����N�V}���_B]�:/tĸ�B�0����Z���<�#��ib ���2�X�K�� ɝ]�=፜$�ZdB(��ߵ�t��Ukn�'�i埼|1��L�ǩiDmM@�#m�\�Dk��SǓ����g)ȟ��"P��)hS��6�g��4E�t}�a�F��9#H��L�#��ޯ@מQ��3�. 8�.�N��=s�G/)ar�Q�"<���*,>��_>>���9��������Y	�i�:�g�f��8@�}A���zS�f�XUm�{ �Ӥ[�dk�b��cS]��幙��(��Sb�$3���q�ģ��������}��?_7n���:k�(�X|Ѝ`,�>ݒ�X��]��s��k�:A����`a�����OK;~��3�����C���o6=��6A�vn���W����yY�o�?C �A�(�;�;+����z&��!����ea����8��BǓ:�<t�k�(�� ���~����=�Y��o��؉����P��/��5WUc�쪃��,�[�q�έa�GK�����j9�o�u�I?�Hiz��'Uy����d#�'"�;����G���ZV��<x�ŎB�K�hN.��ks;\lܜ���_�;�o�p�8>�b���hq��a�-��Lټ��3uI�(�"�~����u���g��b�����ި��� �X�[�v�o�ha���VBm�E�\�;�3~Ax׳���p�P��1��
�ᴙ�,j���k���&J���wk����͛"���NM~,N��<���Y�ZX?R�����D;�Q}V��$��u$�_z!��(d ��*���0���H�n�e�6ǋ�o�\�6���6�
`��Ϳ5��!F�L���{V���ƴ�g���EY��C��;0j����:i'�E���[���޶0�X�Gǈ���g���q�`���~Zw�;�N�N��4sӮWZ>m���GU��s�gIxw&E[�wj�� +��C��wb&iJuKy)}���u�d����(��j������Th��y���<���:9}��������8�t��p�����hZ'�P�P`�P`'(�爦���(� �d1���m_��Dڬ�k}{�Ď�����:n@�>�ÅC�p��*�]�z����CK�4p�iQ"ʶ����{B����������i#�9C8D0�懔L��޻�}��p�C�ba���iç|��c\�6��|<�]���q�"
^�',,�;-�M]2s�0�cǭفnEt�쐜�Ӛ�<ր�<��V�F�&
�b��tv���#4�EX�)���>!�dZu-]�Yj���j,����Gm��ݴ/��}�k+NJ*�6�҉�=ˤ�
�m�Y�ot���'�v'un#�`c����/78���1M��`��:��,��D*�(�oV�F�B�A&����We�<���8Wa��ޗtq$C�"��c-缍5[��kR���hȤo8����L�ENv^�3�����i��۾mn�^�)�������(&{,8������A�X]��2��_� ׇ�:�_o2�Iz�V:S� �g����kl b!�]�	k_p��H�p��r��f�6�	������������;��s��]��֕eT�'�����@_ZN��}b�
&6�e��u��N�٤ѕn&wsnl�ǺѺ�B}*<�-�:���νEh,�3C�҃�;M�����O��&�ˬ����;�e!�ӧ����|�Fm��=��oun��I��I)*��	��Ў���^��[�-*��W0���	���2ml;�v�}|Ό̖b<]F�j;&�雃��w=��m�Ԯ�hK{����V ɗ�s��V� �o�=/:j����4�:}��N�:%F;]쫑�m���:[��0����H�L�N(�g�/)%�/��U��&�C\S��M:ݮ����;�gk�_#.�s�h��v��-
�Z���*��1�AJ�Ɉ��v�(k)�f0k���E�L�1m�6�Km�kZ����3"eK��T11bF�Aq�ra2��X��nc�����1A�\��W2�vS([dV�V�e�[IPP��Wm��C�ۍ�C3m��5u�[f&�0unj�4�5��T�(�4�J�[kݵsv;����`~Z�zu�s�繬�{��ZQ�ݲ����رJ�4�O�����J��:�̋�z��`]�ˈ1�Q����I��[��6�t�P�6t�/�$BX~Y�N&�c�g�\l�+6G��X7XScN�&�:�Px�{{��s#"�s��Јp`�5 �S��4�}s�Y����c���#|�彈#��f����U�+��!�4i�~��ϸC��Bޣ�\Nĥ���:_]+����0D |�4�
"�j�}d��n�6|2�l��b�!r�!��@�u8�O{2� r��y�A���Q��0"�Y;�n�m�vv�ھ�!s��O�p�a�^�^�4W�Ȁ�vNm+�b�8����rqz�p�v�;7ɥ��vY܍��i�o}���Ȱ$2J�6�����mc���k��(q��A)%��wZ��N�@�q��xz=I�"�`���t���c��EV�b�{��7�&����?�o��A�U���6>?5��x^�o�e�����P1�P!z�aY�<7Y45�%x�u�i:G����c�����c�(����O��fxl��g����Q��f�7e-�F�_[*��塊Š�{����O<`��B�mv�ȁoP�9�s��ֈ�8L��l(]�k��ڃ�1��' 5<u6��\��r.+��{��?��������{==bG>)ܮY�u���20��3ON=O�*4=w��ҕ�����/w�$ �����x=�u���ċkͲG�^d�ʚ��|�O)�Sg�fC����\�y��eq;E�U[�B���ek���i���zv�-�1�����1����dd{��$wq2Q�:���|���ּҧ�OG�=�k"ڏ��ܵ{�,���i!}i�K����8rf^s�,n��nG��n�/WfȯJ]Y�HW����E���[׳+"�����U���LD�h��`���^ռh�����F"�f��Os��2�iu79>�o��X��z�L��ވ}Z���HT�n-�C]�yx_y;|�Zp��,����t`NC�}���O�lRdS�<�ݓ��r5���4�����ٞ��,�B�,��h�l�F�8�`\:ur��Okfj�=rBG3u��{g��rFN�l9��h�^�T����)p�9����
-'=��7��ʖ~-k���^{<L��C�Ԏ=�ۂ�Z��#�ԫq6��W�7����I
��-;�֭�/��B�px����tQ<��au�H�k�a���j5�=��ߒH\7���yLך}�W�(_��.p�茎�C���33�W5�Hkc���?;�<��̷�ok׳�]���Q���b����Nk�z6�>6�Փ���'K����F��d��^hװ�s'wwj�^�)!t�a���J����*�]:c.�U]V=�d9:�k��F��S�%��N۷\�]�= � k[���>1�ŽDEa�ȥ����>�t��W����%���{L��d=N7c�g^v;�J[1��H�r4[A��W�vB�=>�;B&�nj��y5�aU���m��u�Kvx���?OwvL��f1+TOR0�iJ�^nr�¹�$F,><f�c��by��A�0f��ﺴ��r�33����l�]�b�>�J0_�t���M��{7�уo@��V�ڼ�nb��,n#�1��*u;��2�S�k�3�Y���0�lt,Ђ���Y�蕐�BJ H�n~���<�bb��ƯklX�W}�E����gr�t��Gm@��.fg�3N��he�z�G���x�� ����"܆��yF���ޙ�EƉTs͌*�;|}��_��	7p��)Tz��0
��gs9��z3K7}[��,q3S+x�ۈ*�k���F;�5Nk��0��}��,��c�d�f��n�j�{R����ƒƲ�q]�i	���4v�D:��MTl��z}\s��� /w!d�1ס�Fn���KU,��\�B,��%| ��T�u��߳����"��6oO\�fRl\:V���)�L��ns�}9VV�8E��!�)���C>��L������V	�x�	͑ԇ��,����Gn�k�u��k�����굕��F��P��^ֹ�O�!2�o��'�C�Ymy?�S4R�)vs������4��#U��������R�D��!���8B_6;Vlxr�P���˾4�썃w���˗��7ڄc�Msr�ͩȣo�,��J��J��Y�Jy�����{�e<֐�t}r�ƶև�ų@��$I�S�<E��{�;�yQ�i����J5<SePohl�ʚ�&I��i:ܻ�F�O�g�˂�)A#!k�M��XzZյ�hK⏲�U���s���~�Ju�8&�>>B��������wg!H΄�t9�>���,�Bd������{����`=so��Y3u��tZ=.��iٸ�� ���̫D������T%++UJ2v��4��[ׇ%k��d�ې뱲�:䃵P���NTub$�r~�����O�����W��+�����g����)�c4����uy����!jޜ>a�YU^�Lװ�	��yko���.\���8<ήW�6�@��s΁�)E�tj����+��� �������Ģgкɸiz|�������'�l[��=���T�J����9lwWc�ۧxq�:ҧo'y���ݸ��ׯd9��G�1�K�`$���b��HXb�xŊ��S����`w���AgM>��{G�bj�����b����#ۭ��	WwJ+�a;�l���5#t�)�f�1���+���T��!����`Ǧ�ɘ��vQ׭���(^��=�%�[Xi;�7������P�.*u���u�s��i��X�r*ۘ���������@�g4�k�ZŴ��UV�k���V�u�-6�$yr#��i@�9r���`=�.`u�$|`�l�	l;�L���ۺ�̗�%�d�}�:��o.��cN��fݕ�j{o�9�"psfm��b��僞a���r䌡G�=���d��\A��^l5�
V��9��]�s��}I_&�`<�M\���n��D��Și4Nʮ��]��۱r��d�z��u%[��`�Η��*j�ޒн=�!8�:�Z*�Σ*=lbA㽧S�.�}�w�)o#��L��1����;:��_V��d<��CD�U�"Ep}J�J7��>�9�v7�ay]yM�;���!ۉF�s����a�t��E��ᬔ[��b�Y2��r ���|5�����Hs����'�Sjq7w���r_���Cr�K:����]Ֆ(���W¯�T��2Q����t0i��5"!o�����J(\�H�RG$!Fd�n6TRK�7�W.���et2p]�!3��/�J��M�� %Bsޒ��U�!��
ܹ��Y�cl�L�V�5�ZєM:�]#�+"�S1¤�ŭE�4̋�a�h�at�]888�i��
�uh�����:��!�SPB��[����	1,ֵ0Ѽ�4�e����Ɔ0�a����u��浚�X�n�1J�PPP�Tf*�nbШ#���)i1�����`¢���r�*�6�k�LݓK���s;���V����e��x���V���X��#���xxC�/��~������2:�s�|�tB��M�7����z�9 �Ϊt�<
�Ԇy����0����:���iX�t�3�:nk��O�.��&�gճ�(3>��ݶU�r-��/�$�vՕw��ٵug^=WI�
GM���{FG���N�[:؛�<��U�A��u�qj��O�{���jcN�D�;�A���W�b�Ӆռ���^9"Ҁ�qz{�9���C�W�Qg\G�(�n�'�A���%��:�)=�1���d�������E��T�D*ZBS��Ow���*�z�FۧJ��މ�̌5:��Eh+E�37f�{;1x	�¤S簿@�z�g�=� �� �����{O��-���w�zn|!��V��vn�v�Wk��^ݱ5��1�% ��Qu]�k�S��']��fȭ77��=���!ܧ*�7ݶ�x�/���d����5t��0�YǞb"s1�lN���[q��hQ�[bnh��s��0����&�o$9���d�ӍTwυ�m9p�Vbq����'a�c�Ǎ3�ߎ���m.O���NW���lϟK3�6���w�E�7+]�,�.0�q_˾��(��y/*{���ex	��A���*����C�̞��xY�H�P](�y<�Ļ�ߵ�Ψ�Uғҙ]��5�W��d�G���𧻓(�ɖ�{�KE�V��J��F���r��v�Dq�=�k�2U�����WQ!R�˧/Sh(�����	�x\�9���t��G)cgAeorY6�/LJo��ՈA+v#q
V�2�D^S�X�FV��q%޴�QӤ]qc=�j�tN+3�'`�7�<#.���;E���!���>i�^�Hb\�����~�Py���K�a�{���l��}����>�mm{
Z'���h�c#~���ݿy��xxVI3��m1���rI����p�7�]a�{i���n���y~�}4�DSW�-�k��LQR�Z��B��P�;oމmݍ����?bN_�S����IԂd ��.+5��bC_
���U��(��+m�����/�5������8R����Նp�uV�^7$_5Z<��B���a9c���t�eRa��w���o�dg�fA�&f���ִcTe�nS��c×�&�*ߢY����m'��9��{��E���S���v#dȱ4��C/陓8$���f��Q�3�i J�T�n{|F�ǚʹ��V�e�C$��s��f'�PpJ�ֽ�Q�	�������s�u���V�Q�z��{h�n�^�ړVu�QP���#�W��#�'}Nn��Kh�k��7z_��zH}9 sh|j���kw�|��=��ϵ�D��ʢ{�~T��Ml��u�V��g�5�u�$�Sض�<|S��E��<Ud��g���ww���1ىTS=�
��E�[� �Ex��Fل^d�z�n�C9�TN3�w2��{��>!tmf�c���-W36�g�w���`��J�8��x
�77�ػ����.���0;|L��*��ޤ�\��\�A����V�冒�T���jIR %�;8V��Ã[����iq�OV��G>W��s��J�+��䙣��M�F��!�u�N��M#{��N�s�#�?Q�nH�z��Pm�-�n��ce`V)ˋ��R����|&pN�x�f�eul�>0LfNwmn޼%$��A�2b����s��^㉌�E�nA��k��Cz`^����S����l_�'�����x��7z��X,Uk�m�tu=��"�7�g_DY��_":���m�e�`���X�k�>�H��.޻�e)8ʹ��+w�۬	0k;�s���q����;�jS�=6(��t1���\=M^ڞ;��TY��B=���)���D=<�:vl��sy��Q/*|i��T��4z����o�r�N{U�lȈ��;��a2��玌��x�늑���ދi��+��U�����s�,���]o�~W��;1HZ5��K+Gk�U�Ҙׯ�VO1M���R�od�6w�L&���X6Ŗ{q��զ@�u������(H@�׍�r�f�o�[6<r�KMG#�@m{���c=j�V�����Ț���;�N�lw	j�ľqb!��ǟ)l&$��֋<yg,F=*)g�r���W�+Am�8�D^Ծ�.q�k���}MH�d>)UgC�xz�;��꛶��"��v�tV6H�*d-��n�8�8�f��+��ܹ���L��B����g�W�jܬ�߹��P@רu���G_2���\kv3e���0�[�W#A���{�:�>֦��r�j/��x��mM��4�;���A0�ɥ�ȶ��Z�wd|��*�H�-�ɠM����(x��CͿ,î�.�!a�E�^yFej*�Q	�����o��o��zMiK���qzDJ>�&,dp���Z;�m��"kKGȪ�=�K������,�E�EG��'��H�U�Op��b�fM{�j���'zUG���zn�D�����=Bb������A�/z��%�8��pS��!����t�D�9�5�:^�^G�)t���J��]�i�ò ;A{��� r%]	F�ImK+vʡeH���c��ʃ,ܡ��������T��A�:bk��Nk3$bb��닽�����f��s���~�rZk�� �/�뚞6ŉgv�p�TMb߻��%��&�s��!g����;���|%'�@^��n�&k+PE->Z���i�=0�5����Z���l'�tջy5��-��,U�ly��c����f�w��P���VFs:x�Rj���v�!�_<ph�]�u(��"pE�]�聣�c+�E[�Q̜D3&0cݭ�w�\qf�=��`zr��o$�Oe�l�_���B���/(g�˵�V)��1Oj����`ͧ� L���ҏ-��������]�:�o��f].[��8�[v������c1�Y�1Xw���Ln��.�ei�5'f(U�9���������Yy
O/���C�; Ѯ3R�:L�����$Bm��f���](���
�?�p�ݝ+X�\%��S���@�t��N�1��r]��C��ݥ�%��AKك_.�;��
��=�r�n;�˶ME��4��-���Y���Q��˜͍��.k��n�q�z��Vg�|���)ޕ��[6w9Hj�r2T��Q�.C�7��6����I��=wR����S������͔p`��{�G�����ʪ�
2,6ʕ[KU.`��-�kh���|�:"�dPY��Qm����h�`�Y�Y`�v��j �+R�J4��h���˻M*Q��S#6�V�B�h�%mJ�&#vʢ�D�K�m\lѪa�3XQ���(���ae�V�6Ҩ��A��}�2�)����Θ��5��E�Qx�Σ̹ү��F�f�$�~3Ԙ�s��X�V22B�W{W����g������>(�}�\�t-3�kzЊo�7x#��yJ�5�+/����mp��%�;F�N5����%?`��%�V��a��l��:��k�5�üէ+���g�:�k��r����L[ګ����\�f�p�Y||��L��2o7��*���e=��c4��u��a��S��ˉy�E3�Tٙ&\U�*��(�d��3x��ӳ��`��)wj3�4��P	��.ŵx�ʟ'.�&��.�,\�m�BW�GΧ!	��[
9�1ѷϹ�X��帕��p����ǫ5�y�3#o�*��h}9�ƻ;^lʞ'M��E� ��kI�5�Z�4��3�n�6�t��%���P|�r��$l)�YR���� ��I���۔�єO^�|��*�ؽ�e�n��B�#�a.JSܣ��
��m"+�R�2�1� ���߹_th���ٯ���w���)#��|��үvŌ3��jʣ�Q��w�M�n
 �cb	�sG8�(-����IfU�[e�S8u~O
ZWLB����>�R�W����P9��4����2�$[����/��*$��9���w*�"jw$O'��jE�fld���yDu�7I�]��s�.C)�;���h�f^�5�ι�d��{�^[�&4_&�)�Ʉ��*(q�]�\5������T��a�A
��v�N���P��.��Y����$���dH���}�ܑ�X��ȋ�Ѷ	��zˏ\�]?r���r�Osλ��WS�.��Ok!c�>�3�)L��Ǔ;0ʚcz[*�4�ru΁�)T1�Db�[ۥ��v>j6{��YC��.��A��B�z�n�'s�7zF�Y5��kyu�<Od��W���z��-Y�,/]�+Pv�ps]\�]��5V+��O�KLЩ�E�{Uq�u5�W�����r2�$O��=x��K�2���/ø�c�oj�>�qƑcWP�7V����Y�[�ׅ�����aY%��O�9��(\�S���9��T���&J�gx���\��kϮ�V�Xx�ʦ�emv�N(����23�'a+��$m7)��9k�̮5;�@�i�I&vug�ŧ}nx�b��X�SIX���K��.-�����3��v�yq���l˦�l��Gt�B�=�#4��:<����Ш�N9"эje-�cг��o��y/<�n1P����=��f��4��F+�Ӂw�ҷγ���k���+MP�K���y&W�eڻ��4ϵğ<B*z�L��Q���5[5�{y��I*��+jyW�=)+xJ�q��L�|6�znG�U�nH�����z�.��k��������ba	�}��^�ǯ��留�ŢjNk�ԫ�Zhl{"M*��sZ����Me���ROHJJuc�����V����gM�w��Mv��g��{����%Ա ����ñ�(+ʝo�n���z��M���oi�<Tq:4�z:�rx��u=W�<��(
e��~�=������L�}#[�|�E�k�vl@91�sO_oe̐>9刵��Y�3���:t��D��X�����l�ݏm�n��u�\�4\�࣎I;'�po�ꇠ��V��� z���\������Y�6a0d�l���_)u;S�=�h��B��p#����/����Hl�
�{$ZVs�/;5��K>˾��g,V����͕7I��w{NC��x�~�a`���ml�P�}��{��)���Hm;TsFy��w�	O�#�gͦ���j�b���<�ج�!v�������b�U�[��;Q�K��q1�k�1E��wfv���[��\��@��`bE�*7��26�vژg��r���3<���H�r���I[u��-�\
уb��5�-~܉����>���3��Z���C�Bʱ��v���`�f�{���jq����1N��!�gf�̔{�:�sq�loP"-��s^g��#�"��6�F��+>ы8T��	��uw��,���r�M���A��o�ZKۮ\UR0�c���%��
x�׵9ͭ�h�	�R5�-j����\�A�n �l:��GlR�Ƶ��l���C��i����7��,��{�<�/ڥ� �ߦ�k�����e�KV$��q͏��jp�Cn��J��:[ӥ9�*�5�/�_�XP�u?	%7�9W��g/Z�m�vo��Ө��ם|�Ӝ؆n�\��Oea/�q�MmČ�fZ�}�7���=�7�:4�+���Z���3����x9vvq��njvb"��]c<����N.P��؂ء�r������0|������-cM�.�En����������\�����u�[����э>[�]B&Tǲ���jm�`s��&��,����v}��6gWИ��v=�S�W��v���u�A\�'L΢���֨�֧y�tݷw���'���r�����۫�3JǑ�o+�2xS�� p�G~��|��ڜ�ygF�U�}��%���J����������f�S�q�U�p���<��~��Q~w�p7N�'~�P��$F�_vGh5�U�ɑao{�*��	�&��9}K�"�^�l�WN*��oD��]p�d:���e1����̾"���I��b�G�2�<����e�����ן@�71໴yj���u� �Y}|����Y�6�1PY{ͺ�)շ��bp_i)q5bS k��Mn'L�vgt�,��
fG��H*�]�)�)�����b�E���m�L�3-�8���%���u�S+-�`���<�R�z��1Z���k�L|����&�����]�EK\DN%V���4�ifG�\8��0�9u{ڙ/�[Wc3�n�k������j�'cǓ�в%5S�vhK ��=4�_q�j���a�F�5N�y�B'�X�ר>�:���J��Ƭ�Wʴ\U�4g�c�)}����]��Z��.��j��;�dj�q��[Ň��
E����c�eY�l�mMΰ�4v�K�3ait���xcv�/��Fmpc�ɇ�4�CH��D����*��T�I�\��+zl<�fB��c��q6���\���UD�=Rʡ�{]̹�D��Ȅ�7}��pCE<N��t�)o3� ڴ�7��u��u1�	��p&_'��fn����-]M����:\�dRlƜ�FK�6�J&A�&Ԓ�4���۱�6�}5���S�q�D3�Y��k��Q����8�j�i0�#���2�(��u����.[�eaX-lF�r�0a�.[FeK[i�����E6���U��3KeX��«�i������ĥ6㈱lRTt�"���0F]Ң�EmJ�EB��ѵ��i�jۦY��n�c��jZ��[GC��%J�l�i��EV�����֫KiQ���13,�UFbU���n�ZU��T�)R�*2ĵ����kmm�)mZ�z�[5�Uyk<�-(՘��%R��7u�ȋ�J��'/''W�'$8���é_�{��}�u���b�(cu^�M��/i.�:��y�,N�=�`���/d^W2���UA��WM�kr�*�8�e��r=p��m���込ݘ<ݸ#���c��r����S�3���=q�YSL�'��d�}z65�n+GX�#�](Ǆ����|��z|�}���җX�yW�O W<]�S�6�e�-����L�#�|у���l�Z�}���y�km5�\ ��3S��s��,m�j���7,d[�����k|�x\��d��O��[�#�lל��8��6�����{q������I5���a�(�i����Pnl�V�[Tp����,x5G����Hn���2���r��n\N<N����&Ź��=)���S����M�=��O7St��;c��t��4p����xO,�t��Y�m��{nꅽ�}1u�x�WJXcek��(G^��ھ����i���\��f�Sۙ�s� nz/Y�+&m�x_L��q�X�6�+����}I���v;�7��M��
8�M���ɻ��Q������W/k�\�a���˖�����/�}�e�h�����qU���W��F���)���@�Gi��mB��Ey�9zR�u_&����3���+����X��	��'�q	���{���+��'�Lk�ǹ�{�qe�^[��Mf����k�T9;+�L����nA�֖���0N5���|U^�=�aMB}j]�����	?#�~d��^�2��u��&�9����rB��b�za��c	��8k��[Z�#�W��#��r3ͯS�b�v..��X:D�4�NX��b�����S�OE<S�'X}x&GX��)���Ǜ��^pfV�LQU윦)eڄ���/�]ǭ5���Ճ���W�Z޴���j��i�9��+��m>[K�i�3xօa,986�pMTm��>صT4}-^e�������N��a{���9ʼ�u����3^ܤ/�Ѵ�����~��}G�����D$Z�ݿ:�ys�yYJ�Z7@�Iҷ�9]�ó9�-k�L�5Cf�\jQ�r5y8	���h{+yn?8ܴ���Z�،k�������N����g^J���hʉ�[��Oۀ�#���'&x��{#r\��ڷ���.:!��LYn����l44mo�Rtk��~u��m�w�\lo�A��۾�+>U��t����]�ж�2�ݮ��۵��د�ς�a�7����4��[V�{Wj��#���o^��X�4�l�랏L���t��[��M#��3��F����h}3��^�݌X��HN�"�4g^�PmH�p�⒦�s�7�m��9p5d2,x�8�gx7E�WK2�i&�?r�L���H���,���d�3τٸ��x��fƍ5�٤�f��1
�n{�J��}b�N+T�٧���CvS��+�<C�k�iu��h�1�vml��3'��>l+B�ң��o�i�Z�y�f[�[k!ŀD-��H!~~��X��q�0<#J{��U�^�M��9y7 Qi�3��'uQaL�3Xy�^��sH��+�eٰ�/�KV�����pƝ�3���4��>���9Y�&��X����𞝾��Wy[�y��dJT��R��=�7zCǭz�~������(i�Y��Jw/ܑ��\�CGS��A���\�S]��3ZU򉷅>ըg�W�|����+�hH��Ry8�"��C/�e�^�Ok��b�V��9�
%��ye��}Ņ�3��3���u�N|��vg!��+6�/����O����m�=�l|mڿi Z�*�.ZQBM{�mH1���ƅ���l�='�:��)�Y��:c����^	E�w����{\���o~�׍2[h��ǁV�-n��&��20M(鴷��<.�� N>48"FMY7R��=t�_�	=7��M��j�^����0��;N���<z�#]��0�p*+���&���m�!���gz��Tu���)�:�O�[҅�}-��]*��VC�in�s���;G�p�氍Ee����4θ6gia������*��io�.�N.�.K�gf���V�7kz^*x��C�{��e�m�\���{�Z�m�];9)��wl���ү�(���$�}��яD-بzX�鴜>/,�Or����A��[�}�29���B�7S�F��Z��˸ìl�9��e�*�Y<���]f��ǘ��["1n��t�fqg�i|&�^O�Կ<a(z�P�ltq?q���ٛ$�#��++��C�����u��]{�MrF����Ү�g�<��*]��8������U<�����ֽ���cy�<B�.8`]-��5{�RA��7.�+��S1Sg����ܰJ�/�B/9L��w7W�d��ELv�sS�sW:n�
�2�^)"n=�X��}.�Uu>([5�G�d��&z�y��a�U���WOk���ܫ0�X Kf�g��p�C� @������U�M.=h�݂=thz���m����6a$��}��ֽv�,wGX�7�-}��rV��밁����x,�^�[�B�]�@��u�y2/�������:�m���~-4X�gj�X�yG�S�αz����g�V3y�����Q��� >��x$��J�UX������	1�����w	!�DP �I��AC�)����u�����z��?A��h��עz�&���H�I	 D$��:�Y	��ٚ��fN��'E����"v���C������R���7��~��?<�! ~�"�OhOq��ʞX�L�� �d� �U�@�z���!�(p���g;�;�2g�ÁJN��-�N�L({�{�h;Ԫ(�W�tğW�^ �-��~�j��/��H���䛿�Y�������>�<�H��0��	��th �8�(��Jz��0��""ې��?�d0�?a��А�`Ju���B �C��ى!�Z���gRH
l�i��BD6��EB
�ft ~T%!	 �8~��{/^���1��v"jB&���&I'��T�͒�(l?�P��
hy�i`��C,�,1:�ErZ�R�����tC0i��Y�:���	D���<yɼh��	��J`;� ?�����G��vN-�
��e�a���-:�D��
dT�'�NZ!��eKG���r&:���A=��u�Ю�aň����]�z� �*�״9z�`Zl>������0��2��\�������e�� 	�E@_�x�����0�(���0xP�h�����BC�6�Ht~Y!$�I�t爂�������?(�� $�d�d�;$?Q�é6����}�ì�I@@��=���!�N��~�	1%�<����3�+�qTQ@]L��o:����"({b�!��5�u0>g��&��D���6���1&
i���d�>'T#3�=X'V����#>�إ����g��HDPy��6�`Gp��!�g�%�j"��^�y�\����0/� �;��1s�����u	�@pC�2	����`Leퟐ�N��;/1��Zh����o�Ƿ�]4�o5e2��eU@Y��&�*�rKwnH�e.5�	q�Б��2�xD&�I�-�Ym��� H;Ƃ��M� *�`¾� &n�/�S|x=�m�G,�y.��5�q�!�R�T)'#}��2���ԇ��������4��G�_�.�p�!e+�