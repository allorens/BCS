BZh91AY&SYP���ޚ_�py����߰����  a5^�@�Và  ���   v4   [d*;��DER��J�UGY�
����H( (� 9��J��ۀPH� � ��Y � �@
���!   Zx3R@)S����/��Ot�9�|^K�wr��g!��5�����o��On�  ����3���ʕ�y�}	i��>�u{�=��{ޚ�{�V�Ϡ�����u��ga��p �� |{8����I}�۾����=�w����}��}�8u��Ǜy/g��{���� ���� z
.�X�x�i��`{���|:3}�<y${���vi�}���6��}�={t  �Ϧ���@�{����lP�o#לwů=7n��;��Zy���>��)\ 	 a�\��v���{���ϭz;0��L:�9�o^��=lt����z�C�P������=�N��w#ݎA����.\�p[�vH���w���+ﻅ��UX��{(ϩ��<m<����`e�y�o�m틶�f绛��:�Gz J����*�T=�i�b���t��������;]�{�Mtv������w �L�Cv��}�x:�5�c��������	���v�v�:@        �         � ��~�Cz�*�CM��� 	����"J�	�  Ɂ `� �'�T���        ��@��A� @h� F  �D��L!�&Jx�M)�����b�<)�x�*(BoR�R�#L&21��?3�O�$�R�"BH����4~�ݦ��A )��ɖ����(�TD�   ���J ?w�4�^/������������#���NO��k�������	$�ʪ(�~��p�QU	%��(I��bX���R?�G[� �;�v?���!����������n3O�����#�J��=��ޛ���-쮉k)8^�_W��D��H��WM�0�벾~Y[4i�"mԤLnW0�����R�4ܤN?DEԬ(��%|��R&��[�JD���/L���M�Z����R'1]�Z���=�ˏÈ���~�Bqʮ����j�rVd�D�:j�NI���U�#؝9��N�Uӥ�Ç*ljlԈԳ�ڧ'Ȗ̕+D���CH�T��J ���MW��}7b[�H�|��1��W�Xo&�1&NQ7!z��;�E��Ӓlj'<��G}�B9��N�檓d���d�7"58nDrtMu��5֪���ؔ)"`�J�5�1�~Nd�����N�w��d����bv����/�.	�o���=Οqu-��Ăe�}R~�1�b0{��:'��-IH��Iz$��Q=�f��W�'��:��$��K�'��m�Wz�]�ʬ�$��w3s���r6o����z��bj�&E0�����0X�K��7�&���7���2,8q���A)�/K)�{B�6-[�CĤ�a�&rxT'��7�tL116f��[���É�5�־��oQ����4��&ө�:��o�h�	'�B�uaf�d���IdtI�#d��8�b=,�$!϶I2��Y��zfvG}:r�M��2�w ������J��9Å�GJxW,�,��J�R��&�������g�d6�������-�a��%�&DN������,K�VA�N��X�Y]:eM�u���J�����DN2DG$�A�Dy��R�h��M��+�r%~��Q�%|�Ț�"<����J���U���"q�H�r�h����M��Tt���̕��e�?`��JD{��O��"i�H�~���Xlu�_?=����Vķ��6���벾�������9���1�a��e|���h��D۩H�ܢ�,o��|Ԥ��"q�".�a��%|��R&��[�JD���/L�!���"i�Nc+��~�o�C���N�+D��nI��"k�Q(���ݲ�~�ʪs%fNdN���t䛹�U��N�O$�\:_[.K�jDjY�Drp��Q�2�O�$6H �粒��_o�5_W��:#ɲ�{)`������Jç2^KI���%H7��9��$��NyUcu\:;�Rhs��Ԯ������d��H�N�����W]4u�r%};�jVe�~ì��vH9!ϑ��IG{5�q�J̝�bv�����/�.	�' �"���=�����[R~�?T��V��q,�K2��Iz$�^Ĩ�ԧ���RPOp�P���$��^�>�^ӷ�\Z�i�Y&Iq��f�{'FG%�n k�w�9�?x��<=�n��������D��}��s�d'H�A+H����4<�w��sͦ�ѵ:��,��R��9�{>�N���Q�Q5
�R&�'��4&}g	/�I�:��h��:Y�䉷d��d捸Na����/���
�Q"D��f$�����[N0ǤxgnI�@�œ
oF�'gv�!ü��r�m2	��'{�/BQ�vm�8�:�Dr\��ٳ�܅�-!l��q�:�������$��,�Lu&%�ܛ¡�nKК�&�ol�ћ웆��i�x�B�K
�IҍІ�C�<5��P�J5F�%%�1(��Ϸ$�$��%D�ԶG{%u%�'�;��߸$L3t&�	(�J6�'-��|�L�r&�!&2g�#�D�d��:2��d�x'Q7$�H�(�'[�$4u�#�$E?"�L'�,����H��#Z'MԈ���eB"oi�N�8�Y��H�󄱲}�"&��l�!�RN��D�&|�*�"Rs2D�Z�h7I1�d:Z%	�K쐡�l�7�)K�%��"k�)�P��h�	Q"&�"?q"a��J��:i�t� �*�DJ�DJ�D�Vj�M�&t��5��/E	��-"tvazF�"b'�ԛ�%�פ�A86h�"'>��pt@�a�Ii�G)8&�ȗ�E�e$��L���	�LxD����՚5I	�&�1!�~��"lEܔlM�c�E(�%ĉ�N�G�M��	�"%��&�"I�2�42#��G'DÝ	0��9s���JuR���ɳEȍ�w���^���TKK�"������DD�f�O��(�4YU�"oc��ɿ�n5>�*!��lL�8��鲷0�"=j$Ƨ�'�.��O��iģ�ԇ{�l��:��'�Uʹ��1�x˝&r3�l��@����}���=���X�d���H��";�4nϻ��D�8n�S�<{s��}g��<o=�8MD���S�Ȕ�a�;�c[���QD�ڛdٻ�nl���ѽ�k~fy{���VqOY �艘��L6:$Dyu0�BU�4%�O�bh�}#ʔ%�".�a3� ʨ��"ijQ�F���&�r"�#9S�Fڛ �|���Q;bϓ��5��"hY�f��ު"a�f�4�4�6C#S�7ș�ȕ�ԡډ��-$�tF�"2t���_":�DE�D��*"&d١���N�P��Q�TN���ݓE�%�uQ�T��N[Sd}eT��'ls�fMԲ��y���ډ��TD�Z� ��ؔ[��#��N���t�5(�C'Ȏj���(FeDK�'xԲ3e2�ѯ���,��#�TG�����0j`��T��H�&w�1$�VK(���h�P�(��Sd�NaBSu4h��Yu��K���rkBu(��(�0�D좮|���Q_%�T��H?l�G5!��GR3U,�&N��*Qߓ��܉�Fن�vU�!��(MrY�N'�Y&��}��ѭ�&�u)6iʖp�u"ژ�����k�3���T�b��A�؛uUҸ#yQ�0v�D{��L�jl��*ڕ�����8{;���خ����@����%�7��e�d��;�E�h+�#�Z�3˂�L3�3���SX�j3ی��=؞kX{�o�M�i�)L�3�3�2�t�t��ʹh:���g���w���{�l�c�`�C�c�f���p3�=��g*3�>��J�gHtIڪ�Ot�=��W!�S�tx�/I��9F͏d^��6w�{���)�2R�=/Y��b,{0ە���$���ɜ�����f%�;�_Gq��F��E"s��s�z4h{�d�7�up6�|��}4���:��6���l��:�xѡ�_C~eP6���"���t�&����Q���=����{�U9��cS3
�ܩZ����T�ʩ�N�n �K�V0�Db<Ƈ�-{��wu3#RdJdƦRD�y$��Dy6��h��M��+�r%~��Q9{�_'>D�5)�DN�Ա)ܤN�E�*�${)gYҎ�J�D�g�%lѬ�"mԤLnV}>Ϛ����?k%M��7�iRW��]-5*��*e3��;����XI>3U$$��ܯΓ���j��e;,jy�M�6��E<B�q�Bd�HCo���q�V�q-Vo��U��ۏ�I(��.c�g*-��%����	B#|*g��I�Ǧ�5���;6���5�z���I���*+|0�I,���d�puu���t��8������O��m��0���J�nS�sE�����l���7��:���U_F-�ͬ�[�Q�i<��'�_��x��k����ES�����(nxko�Sg$��le����cY���ҹ^ww�Q��ÃG��͒F{q�w����q�l]&�ɲ�R�Y\���U]��C%)�*l�a��.��]��jx&�	��PZt��;�{�B.�������K�z@Yl%����S$s[d�����q2I����9�f^,;���Q����I8<��r�K$�Ihz��VE��d;n��Gǝ7��-3V@pcΚ\}��4E\'d �|hR�Xk8���'Y�o2�L�ڢ�"-�XM:���� ��yϻɕr�N�~#<�>�n[i�l����ٵ�V1��5�������ޠM☖�A���囒Ia����m� �D�����4����a~��OO���6���w�_$�82������.ǭ�� �.16�g����Q$�6�[���0���50 ��[�5���f&��F��v�${\���=�s�gi0�����_H��!я�M�p��D�wp�  �f(M��;ޖ�S��oF9��Z��Z}ߥ!�>D�q�C�� �DJ��]��|+�` l����d� ���&(p`E� �<3� l\l��oh��c���RN�0l`l��ӲM�3:C{���l (�3o~�e{�  3d84����jr'�4  N�oMc��g9������@bߦ����o���Ն)���$�s��){�h\��P�gB���)��0��J�Z������;Ř�>\���<��l��� 3��N����Z�����筙�<t�=���{�9�Ž�wFG!Me�g3���l���S(��m����:����YLL��"�zhsW��i�@On,w�O<���+���I�{��7� Ğ���J�'b\{�+`{��n>,*I�Ʒ\�'��C�2 ��ut��/���*0��t�]�pJ�o�wx�lg�}O����-ݾ���h��~�OI0�~|� ��_i���/kv���>�H�\٘[�Q�,�Dg�dݽ�����(9��p/&�ɋ�WO��8cF�IQ��wc�v�2���{����O�Z��}��p���|��QB����zq�W�^�#:@ݑ��~$ԙ�l�nea��z����ej��7�d�T�æf�.���������}���%ި}b绻9�R�G�!���,K��[��oR�&h1g�r�<$��cH�8p��N��#�=G:�G�����;�{�N�l�F�7�bw9�U�;�p��I$�x����ÞԂWnOH&���m4|a�����=<�ǌ(@^���G��g����k����	!Nv��� GFH>�J��wd�r�y�&:�={����f��L� =o0���<�P�8ۍ��K�s#%�VG�wk�l�����jd�@��==�p��
*q��{��Pĉ,�kw�M�6lf�1���-�C]�Rz���]O83[0:0�OR襒� lѺM�RMJ3E��ϟ=���_=@  �}�Ťu,��n��o4�D��%�m2���	$�[���I( #���  ��iM�����4M�@)��gL[:0c���wp!�<h����f�A��ɫe��1����g�#]>)&��R�=>�S�w;��:@��v/fڋ$�u���q��l�z)�}o�����2v9	��Á��{�s�k�#T�R��a��i'���M(�}���Y*�Ie�&�SB܀0� )ɋ|�-.VI�l�Q��)[Z�Y{ךqHt�3e�6��$�a�.�kG�ea��<�);o':^�w[k=л�Ѳwr�z��_H�9S�O�a��͟���p����)I�Z�=���sNyVO��m/�Ϗa������^����8�(��9�u������$�ޜ.��$�	Neu��noZ�K��k(�w���Z�+OI5k�]0��=��8Q;$�J�e���y�i/�� �   <x�)�� t`G��tęWuaX���4�Zv��O�k�XL�I'��Yk�ֹ�vBc��K��  ���޸|t���f��k���mR;����֟f��) ��u6
?$��� � ��!��  
0 >���8@�d    �I����L��w>(å}�ϲ��$٧e�r�Oj@ 48=s��6bg�� �/$|���� ���O�2|ّ�5}r��$�u��x�c'�4P 8h۾)�I�H  ��3c80  �8��
A�U��] N�s�㳺� 5$>|(l{��4φ|0s;��=�p��!��ަ(]Y�Ǵ�SJ:R׆g�:}�l�_�E!�u����(�45[����.�� 7�.y�J*��髮{͜0��Y^���8L��i��GP��E��A�����7�H>zN��
0G�������]���$60=�w�<�9@9d���������g�͋=�|3C��u|�	����u�okL �d6>������&N�xJX��!e]l�[z�ӧ�.=��g�v,bd핵��{�R pl$��36P֤(ߤ6= ���M8wo^h�~�pe����z���xs���]\�ѰI�e�z�M� �"I&b�Fv�{Y9��K7T�p�Ϗ;:�ɬS�	ݚ"B������$�iӥ���N��	ͣ��a����,�81�j����=��k�Y�� x�~+B_y�u�<6#ˮg��rБ�&��D�E`���^5<3]l� ��v�v��D �ɽ�����:�,��[1n�(�ET\+ݴgs׮n	��oNaǕw�S��o�? �w�+�<p��8�,�k�*u��oNLIw���!�L`���3�����>�5'�k����H{��^ A�tQ�j��9fU
�va
7��ϻ��(���`+��R�T���m�I&�E/v���C����F0 ��e����b͓��)���r켚��gJ N��Ƨ[wV���Ig'`����[��k$�tn#�f�9|�2ñ����g*����6i˙�N�0)Y�����"zI��8�e�{�\|���G����
e/�d��.F���m��:��'��(�K�.�I������b�,Ƈ�}|d�wNN��� ���sÕ,���zO�����?�	���(���~_����D��NP������D��$�?�0O�Y*������V7(���DaF��!F�L�����-"�Q�[�TF���(f3!kP��a`2H�j�$�)�<�  �%1@��AKdCu'H�*�k�6J���.�6 ��&��KM*f���RH�"4��D�mW.C��1C0v0nĨ��vm	m	]6 �)n���	Ը��o�����Z!�23@(愖��T"�-	ԉ�p�b���CR&,�ƓB�\*��z$�u�xŤD�f���6�7q7���QD�*"E2��?�����nW�ĸ�[��Tz�ci
'�eִ�&Zƞ*$��*�b��2LihQ�k95����R��j�g
%���U�lI���JTЅ��	<1BeMQ0@ˑ1Q���iT!�43��s��(�`X�	)Q��@$\���� �S����(��j�M���KKKKG�V���` �"�&�@A/�(�%��1!i}w�#hAv��D��EŘ��@l��*kV��^\�cTj���J�1Wb�:!��+�q
�yUN�O\�ťy��s�@��AT��fGr�+��Ȣ�o#Tm≰R���
s�e�[��H*)	���>:�v���qu�Z�ɊJF#j�jAZq��s%h��(!&*�N,r-�\��
h�ؤ�6�\���TLs��I�<<p��Z@���n9eٵj�KחC�ҵ)��pm�!��k��n����d�z�Equ�ף�g���L��E39�Y"��r�y	;����.���v)�P�hCP�j�ud�����j���s�)�/d�@	gi�9�vl���0�&5�%��D�^��+��4L�
�#�#�wb�����b�B��r�=�;�k�=��Q%K���ِ�|��f�<b�!�Z�9���f\5�5�T����8�I��ٸ$�����cu��{U*�.��	qwp���Rvqu$u17�Ej� �!��1�RN�Z�+�P���2��<x�-���������q�GZ�����Y�xI�D���(;��8�*�ԁ���3��UP��t�C՝
�W����?�dr�����O��g���2PV�J�������v�����uw��{�����UW�������V�t��UmUګj��[Uv�ګ�]*�*�⴪�v�ګ�UUq���ZUU�Ҫ�V�[Uv�*��UU�Ҫ�V�t��UU�*��t�ګ�]*�UU�*��mcS�鿾�u��[,[B��Y!K*�%��%R��%[,�V$�l�%T��U�-uM�&�JX)"2	QT��HFH�  B}U_} }��W{�TUUTUUTUUq���ZUW��Ҫ�]*��t��Ҫ�V�Wj���U⮕W�Ҫ�EUUEU�Tڪ����1U^+�]*�*��*��iU�WjҪ�EUW���]*��mZUW���ҵT�;�p��Bȶ[J��*�b�-�ګ-H�`[-U��*���:�T�ʴ��-�mKm�P�Ƭ�jZ�h��5j�Z"�mT�����	@$!>�+�w:��U⮕W�UqUUU\b������J��EUUEU^�*��mU^+�V�]��Ux�*��iU^�UUĊ��ƕWj��*�Պ�����]*���ZUW������ը�ڸ�b���j�U�.d�2H,���%	�Ij�JZ5I�嚲[��l��Y!�RA%%����|�=���ʭ���mU�WjҪ�X���Uqb��,UUŊ���UW���*���Uڭ���mUv�j��[UҪ�ZUW���զ�^q[UҪ�b���Ux��[Uv��U��U\EUx��t���+UK��9`�;*�� D��h�".�+��l�QՉ�'(Ղصb�P������	"-E�
��j"�@
��AB�PR���ȈTV���d1j � �����D�TV@{�ߙ����j��I"���?��?���~�������'��(�#�0�#�&�'M��d(AA A �"P�&����8$�"bM�A(DM��0D�bt��,�!b ���4CB&�Љ��pN��0�RtD�:&	�0DDã�h��B&�,興���&��'�m%��NGJ8��6"tDM(A�Ȉ&`��p؛8Bı,���(J# ��t�!a�M"Q��N�:Y�b'N�<���g���K�rB�Wd$�s��=�q�Kg۶��0�]G���nZ��^��z8�m�e�8�I�~��q���}����8}�&�W��ۮ��y��t�����bw�rs��Y{;w)��8(��}�}��dہ���k�nV�ƝZˁ���y�{}�[`NP�[)��4v��b�Mo7	�v��<tu��9��p�|�[X�����>��k��1Z�Ƽ����o�}�5�S1�n�Jp�ڝ��ɔ�m���krG<��֧+se�Ec;�s�� ~����8�\96HDɸ�v��n��݇��[k=��BYUqV�?��-��a���c��^zw0�X�ɻYCs;<�[�v8q��Z�p���?s��Ӻ�8L$��6�� <�k[c��~�8C7��HU�t��9�]`��@��e��gq'5���;��eV睬��yn��k�
�Y���V�v��o\�}����z�#V�ӌ�A�k�tnkX뛮�@����b!Q�.�
��R�8�--���:�����j@F���_W���qP��o6��?��k��ɷ���;����}
�΍���gp�M�S�ꇍ`Ks���45��1r���!-9�t�bE��cqV�i�^9'��4 �n[��R�L��;(u�\�����d�lɹG>�ܬ���v~�~޺�셳���	�yd��Nv���a��"�-�s�<*Kk�ښ�ѱt,>i�&�RRN�K�G�	��:��p�Y]<�a�-��讲'����n}�m�]h�ZY��Æ�	�A�k�	�>��(�{E7��J�� �k������[�`�
`%la�T�8���MG�\s�=���6R�"��JT6�U��t�(�,r���'��l�����+��pR#Ȍ�*�n���7}ҏ|���mŻbú�<�Gn�c�/�{v9j����mk��u�K�=�����n.:��#�nMv�x3x�ܠ��c8V&�� q�[a�f�p�ņ�g'U��[�qN��W\�s�e��Χmr»VWu��@�[m��g<Oi�g�"�U��}�]�ڄR�&ƙ*d��(�
\ͥ��\\��|�5
��b�wg����x���V�;�G�>	u����v�Tnu�1�[/cH�ѻ:�+������[�-а��� X��#u��u�`�����+��t�ċm-��U:�q��'�K�䛶x�w ��8^��5ܝ������q�� ����j;�_���Mӎ,g<i0� ��
g�v�n7]�[�/(��y�N��	�؋��#�Cd��cF��m��\����<�{F��ݷnݸƺ�Ůz�I����q�x���:$B��p=s��[�Mqv�[Gc���klUOs��.޼��6�ږ��۟[�Y.�X���)�q�:+���k��xx�@l�ܣ=��������^��J ���l�۟&X'�`�ۧ�����S�y'��x������;��ǭ�r���s�v1s^ӷ�n�ڷ7\y�v{ �6�T�-����u��A��;�Lwǎ8ﰉ��g�<#F�t�줺�^��w"]<��{g��
oi��_����~>�sn�wY��	h��G=�����py+ȕnێ�N[c�On��5�[�B K�};}|F�yؕ�G]�`�Ͱ������
!6�l�9��L���ony�.X�r��.���0�b�������0���;f�_�;}�Q�6'�\�.f:������׳?��A������ffg�UUq��������{�+���QUU�*�����﷽�ȮffyEUW�߃��7���33=����[�}��?}�t��4!e��	�,O	��%]^Mqyu�As�R* mQ���W�&���pB(�D*ډ�6�pA�B�a�[��m[G��zE)b �qD��*�����]��ld�ō�M�G��n�W���n�}�!�6���Ĕ��I�U���ֶ�A5�#$6��܀���X��2��Fq�r�mȻ��\-�֮�pI�k�1v��\u��0���\���.x�� �NvE#t�\��#mP;��;Z	kr���������qt�5��lw[�Eӽ�gl=�Gf�x�2�c��v4�̦ϕRD�;t>��J(
��\jƣR6�
�=x�n:|��Vȼ��6��>������b,�����c%��^�s1&�2�#a�p'��;c�lyw��O�dp� 	���Ğ4�o4|�m��m�����1\\ż�m[�r�<Κl����C&_���B�hٓ<:Z1�Ru6�I�p��t% ^Z4����kG��ͯ�{��L����E�h�$!I�I��L�w�B�e�3�/FT���
� ���Z`�E����,.I6��6`�f��!e�:h��<pDL��������s�N��6-�� Ǚ�4 GN�Ѥ��&Np�9�4���z}�:�I�$�yo't�R90bp۬I2b9!f�TSdd㣄t�g��	^"�����5{��D]q�!bp�V�u4[�����#��`gE5�N��q"i;�����!�QSR�����q����J㍽mۏ�	�0K0J:&9S��+_j�jI$��Rf���za6_��0��̔V̴u=VJ���'�l�B��p�:iaY�,T���nt�3\�n�nQ�+���x3ͤ��9�=T��|5��pgᛒ�N���%6�l�1�gd�U���pt�h�u��HJ���XuX�e�^OX���kj(�U4*��f��t��D�,�(�jYS>�CL ���v���w8��]O@����oQ�|�K�����&R��MX��1d���[����m>�S�2o=�k��k1wR�YԳX�d�OSX=�u,���2xu��CQ�4îp��q8��Nl�sK6�2l��>6s�g�8�O_��i�'(��h٣����D�tx!�átBK:d�u'�cq�m٤	jm�|5�,�P�� �Ab�FCOA&�|�  sx���B,m��H#2'I�	 �����v�n��q�s����<��w5�[c�m��޾۵2�N-��?s��n.*ΐ�X�֬��n��c9��nA7Ga,����L��ƽ&�M��&�OsU%U��ӹ��Af����hpop8x��4�m��2�xtb	�� 3z�IF��0 G�|	��e�_�G>��;9^*\+���{̖�pG�o�K8kTMLU\�r��41�%�;��V�4*)a��ǋ踼Tz�5�ҫe
J5�ᇎ�8Q,ѳG�"`�'�a���{�z�^��y���[/j�����_h���Y�+�����^�¦/I$;�)ia�������8��FgW1\Z̀	ŵZ�Z�ޚ����P�K�ޮ�@*�i�g�'a�&rQYzp�lѽi��{�s�����1�|��Z���5���x�9��[&��6zHy6d���}�ٱ6B�`g�!#�l񜟙=mӦ�i\q�6������&	��en��%h�kEUU�I$4�)4��i��ZZD՚K�NN����A��rl�AA���xE[�nP��H�6�v�n�fX׺���7w1M�xA|!�:Q��n�ϪU;<�ۄ�rM���L��4����g���9ݽ�u*����L��g8t����ĕz��IT�6䲓'�dɣ�K0(�d�,��"`�'�g�n}��n� �P���y�3��wŜ\@h�S�aq�I�-���6;=dp��#iLЯ� ��C��N�x&�ąl-4�J�$�l<p�$�d�'L� T�ۢ�Y�N���n��*�E�i0�6zy����Sex��r�\`��O6��}h����<c\�&���9JH����̖x0Q,��GKǎ��`����t�
)���i��aP+Aa(�WN�%���!"�G�H��k��Sda�+n�J��2�Z�����޴��l a�n�vA�����(��=s�Jl幻$�]���Ga�����+u=��Q��m��^Cn}8O	w~ǐ���k�3�Ǎ����N�Q�i�X�ZJb�b�k^m�K6��\�p��9l�Rd�Ú�,�)ts<���� �>`CК0 Ƴ2���UTV���2WSa��OY���&=ʪ�Rm2F�K��B���ϟ�yVB-�c���׈��ch�iq%["�D�1ɡᓎ?g�k�UZ�:��t�g
!e�8hK:"pDL�tL;`���d�I�x^����R������a��|̪�ɒ�u��p��lѓ��I�"h�i�nN�h��<� �ü�1���]��X.�F��F`�#T���Y�G���}u$��f������P�(%�W5�-���3o�[�)��<IN�%�p/��u8T0�'���O�(�O�ո��.=i�ڷ�4�].�ƫlݕ���5mY�U�bՙl�U�_�+mG�4|���m>W��|�����׋��۷�i~9�|\m�\\f��o5���_�����6�ϵ~k�5������c֘��{c]�����i\Օ�Y�j�Z�+�5W-��1Z^���b�N6�ح�+���v��_��+�.�?1�=i��q�L_ˊ��b�.�_��7�mb�ƚm�c]x������q�M+�b醘�Lv�+5����L����S������]1�+�m٬\]:k��5�[�.+�5��ok��������mb�����zƷmǭ1��-ƻ_]�c��t���..Պڱ�[���\�R�*�5�U���^*��+�qv��V8�����q�8c�_���o�m���ƻ_?S�>��Αj����款��2�t�#���{��,c;�*��nE�x��g���u���FR�n���=��=��"�p����x�l���;�-������̨3��7�[�
�]��7�]���M�y5�?�'��7�f��37ϰ��%��:굷\_�.|}�o�w�G�ff~����1WO����{��L����{*��*����w~�əy����O*�����]߯3+33��g�=�yWW^>�p�G
��!�f��:Y�ǎ��xO<'��Wh�h5TUQUEUN%41!�2��O�Sr��4i���=�$y*r�}K�.S�-{����*|�<d:1y$�O�/�Vrp�Ӓ�/�C5�g���sx%���4)��I�_�������X�Kѻ��v�qB)'A���@`�RD��p@뢇Im�H>7��a��\	 �)��ͅ�rQ��i>%�� �`�}UV���FZ0�P�6Q�~��+�'#��߻��f❬W�8�*t~~c����t鳦��a��0�L�<xOݡ�:�J�L��ft{I�I �xp�R|A�4
3$6a �E�9ԒB�`u�H�9!�!������
��/���L����a�����Z���	��u`%q�B˕�S���*�%_-���%T�`�krJ8�R���'R���H!������0r@�0rj��Z��d�_�h�dڲ1�����D<A����7Ϸ�o��8Q�eOc���cQ����ɨyO�S�E�}n'x�r��\{_K��LH v�W��ZRv�����Ϳ)��J��ox���;"&	�p����������j�M��C��1�PeV�.`�>:�v&GF5nC�Ҋ�I��#�6�m6�hH˼fؐ⍼���I����ǯV�ᇅ�[�=t�{�Y9^v�\���=n�a���!��ޞz� �(�=�n~�h06�W���A�n1����X�&�%�)���HK>0@a)J!���R�Wt���8B��6�ObΕ�W���Ҟ�8���p�8|FD�VR��R��C�rA>ć�J�Xq
8Ѵ�n�9��ZÉe��e�H h�k�x��fx}uR{Yٌ�uGT�T���n;����Z����lnO�m���l�*��9�&���z�wO�&�JJ2YHB�aQ�����w&�ꗘ��lJ�,���v���6�����-Ԓ���!#��AOؒ�Q"t�3�<Y�l�͚:h�b'���`�:A0�q�kU&��9�3tUQUEUL(���@8D�mQV�m+��=�n�)��PX��X�C�J8�JS�2fIg�4A8��B��yezb�9�
rH�<��C	�l�e���{P�>}nJ!�TvHZ= c}7$��bJ6�z�����F�K:��lk�).H2U*�KK���x�!mc7�Ü�ʷ8�d%���3
!��"��S��HM�: l���D�e a����]UMi�nW�t4����ً��S��QX(���3$Ot�kd4���7=W8ۊtqҺt�4~/�<~8"&�ä����Z�6�m6�hX�Ц#���AE'ͻ� �吭W� g�R�䇽�����6Ro� �@�!	Ci�sܕU*��"ZXs&[GdsK��wF+M�ąHy�Q�"	$�E�@� w�?4�Ɠ�?[m�e<S��&�捕�%6�a�:�,y�0�K���0۲��Ezy���u�륶��E5�Pĩ�mS�T�Xq^E<S��hUd�JQ�8��D��d��?�-_?1���t�6��:��z��DN �E�o5��V�i���uQy� ����=�w��N<b��oޔ������_����w�	hj���QUEUT4CI� ���G8�4�d�\��ݯ"�=�8�(�=He��[VKBA�	�w�p(�#�3�C2�?_=W�U /����Oa۪M�t>�g �O��&�oD
C9i>ܔa�T|y��.H:!5
�R@��ZC�iJy0���#�X�����1}N;0���y䣩���gx�����$0�	���Q�H�֚h��&�3�9�_R�a��vGJ�I�m<=�<X�yZ*��D1D�UТ
 �3|i��W��O:WN�z��:c��0DN �s����]fP2�8m!����$�-aRЁ*`���m�)X4��`�xi��C��~}p\��Q�r�W6�ߦ�K4~h$�H$�"��)��HȈm۶�ut�퇚�]E��cQV�q��N��h���v�X��8�Gn\�a�9�I��P�d����>���cs.���y�j�Y.����$8�H}����gx���m�t���d(5�}�;��|�x���?6�%X�=�Rm>(x��Q��R�Ӹ-5��9�$�	!C�I'šI�#��:�UΙ0ZRC��ҧj���!��Qn�B�T!i ��;�=ӅU`�p��I��s�_l~�Y
ߥ+�ʭ��[��So\��N��9�w��<��d=���s�w�w��꼲���:ڔ�Y<q��cb�)Q����'�`�+5��s�{wK�-�e�Sf�R�D�m��&��m:Xr+8�;*֓%F���B�����4X�0d�L�lО6x�pDL�H&'d�P��I���9������$�H$�<N���GNHc_68!����}{ܫ���CiX���a�d��Zu�0m�YF���j2HQh:}��	�x���yLp�r�Ž��yw|3|W8��tko]��3jF.�#����u�ҔCx��b�:@�����Z�B����J��K��eќ��t>�i6ٌHV&�VosA��Z]�e�!Դ��D0��k��;4�1���Ңla��0C�gJ���9r��e�SD?6h��Y�6h�F	���"`��:A0�d����z�VoA�QUEUT4A��"t�{�98��B}&�8hl���ѷ��`��Č\?l��|�����4X�!A����{>�V��m����`���
y���"�p:��V�*`~�������*�ĭw����g����6�+��5��T�1cSv�Od���E�a H�������Lm3�D�Sg�I};ܓ�6u/��c��_�����i:Y��Z2U���d���!��6B��4}��d6l��G����pDL4x!��_�ļ��:������}K��*~��	 �@�����w/'�:���@�I$!]2��d0����0�`�]Y+)u�3���0\���H�V�;�W���2X���-Fw��0@�Y��r�v�́Z#�r��$�L$��<6`tB�ot`/ra>0���)u�o$��m�)<k.��;����֍������|C�ܓ)�Ru$L���'k�Ѱ�<��-#Nħ�l�q��p�}着2�`��ƞ�_K�!Ғ~4f��pJ�OHx�qq�LxӶ5ںV���ێ�V�mŪ±j�՞+�|Vԭ��暟,ھY�����:_��ƺ_��隳����q�3W��q}c��5�X�.6�[�b�Ʊq���q�_1���>k�c���-^}-�Kk�±j��b���k�b�_>t���|�K����_������X���q_��mq�S���q��/���b�ƽ_�ΗUqq����7���X�����<kJ�V4���q�;cLx�cYm�}cLW�n�+4�MN���c]+�m;ZƱzݺ�5����c�X�.���+�����b�}cLz�ǭ~x�/��Ʀ:k�Mc\\]�j�qƌ>MB>F�����*����qf/����f/k��7<v�R58W+���O�釾�����Q���	+�g�~��Ż�e$^���'kSVɈe�^��!duY��#N��ǭ�	?����C{�>��w�{ۦ��r���a'2�Bb�c�鷫���6l����в륬h�'��U����
m���%��bCvg"%��Pz��є�����#�|�(�ؽ��}�{f��/_��)=X�N7���^z�s{�owo�U��S;��R�:��J�K�؟c�t��� ���/����t&�<�pW���˅����m���Hjf��w���F$J֡L(�`��
����[�>}�d��Ft��nBp,s������7�9�llNy�׻{�0F���z@WR��oP��!G��L����ff6lE0\�r$ծ����㯮w\��sy�_��s3<�����{ˈ�����2�33���W��{��"��]߯3+33=�O��{�����]߯33Y����}�{��33yӶ�v�xqҺt���1�8"&�ӢC
/��}���j���c���1��L��p$�g���;��&8�O��"�:���n@�x���=�m���Ĥ'6�[.\��lgI^%zlv�m�F�[�k��>�ID�m$�R=pUUA���l�#]������v�]n�hs�W���d(�Ї&�3<7F�|��u���p���y�kw�
{h7\b�}qEӲ�!�9�V�=�c)v�þT�{�S������"�����?`����u�z7[q�/�����[\q�ֲSg��XK�W4�Mژ����9<��	\�c���<Yn(�'�
!ִ�,Q6��vV;Xp�o��>{�l=���_&:oct<u�v�1r�)�#V�*�=Y�i:��1�XЫ(7��6�Q�V��)�Ѱ;���	�f�G��m8��h�8��7j�g�*�!7�TНm��&���؛x�^9~:~OM�NԄ�!��y6��y���[Y�vۭ5�b��Uq(�G9$�&SD{ԭ96:!�/SG+^�n�m�O���	(2��cfw��9h��4�8����
ou��Q��,�����I��?:C�.����!�ri�`0c�F�YI�솽��������rǜ[ԭ��qhW�w��|�?E���Mt���@����c6x�FL?�rP� S���z���ey��N�n�۵N�:WM�?:~6x��0DN�{|����|怜�CR/wb������(���0;��)�ƴ�]J��K]$�cf�t�P���<�l��8L^�i��a0��m���w*+��Ha�~�L��M^��( e�L-�Y�<���>1�O���b%Iр��ķ�q!�A����g�g�^^E�f�,��*���d�ʁeW7wu�m89N�!�oW�'��0C�Р�y6`��I
ѥ�#�"����8J2t�!�zJ�`2���Uu�m����o�5��|οx�x���:!�f���6~?D��!�~��1��T��1�Xп�_��I�&pc{2�l�09��snJ#׍^UHSY�F.Op��׾'{��4�v�N~����x(���F���c
��NB]0�Qn2t����������K��n��oy���?s���d�~��\�FQ[�Y�h����pp3����8���?vUT19A�`�X��(;�L/�Z%�!I9��!2��EQ���R_�j���B�k���~���ǻ	$龧O�S�o��v��qҺt���?:z��L�D���u5eV�D�\�ʀ�1�c4fm9���_w'�����с�(``�~Kp���| �6i=&��R�$p�o��6;\����05��e�b�Χ6;!fuAaM�����ID||a�5'!D0@����ݺv��Gƒ;t;!�<�-i�Id1�0�2�r�;p��͎�b$xi7���zJ�<BhvC~J
���0�m��}B��0�P���Pv�B�6�㼓C��y�&�6@�Y>L>J�	U�ҹ��<z��ON4�N�coD���p���"t����׳utX�qk_޷`B���udS[��VEt/nn��p"{8���I��J���Ɲ��}���1���?����n��ȏ3چ3�;N�t6�۶v��\��<l��tsO�l�c��n�<v^+s�����Z"�� �E�M�_����ק�:oo}�wvoT�ݫ^v�ǘ=�� �o;�^�c�!5G�iA	ު�7��6�%ВXZi�tx�|�pƟ0,�#a�5�	:L|O&�惸1TInrq�|t˃�;��T��UwS�$��`,
Ja��t�v���M�0d�S��*�A�l��^��Vk�q�2QK���"p�g�!� ��� Ly�Y"İ���Y*4n4iȬKQE'�<�=�3�X���� x�!f��#A�������ב���=t�i�N�6���Ο>8xD�:tHg���|�ܾw����U���t�D�u��v��//oϮ�3�z3M.��8�u/Ovt�}R|sSS����wi%Knn3֗����ͭ�j�'��]��2���A{���NO{˧h����=�f��6�#ߵ�Wz�G>���杛өgV�#
tZ��z��o���N�<��;���P�����
(��(����f���dt�La(�Cg�)3����$t�Ox�g�'��x$S��g*IZ0JO�������f8F6�v�$2���UVR�%��ֶb�k��N=v�#����w���RG�J��%�^�Y���G������?M{��N��n{�aՇ�ܧi�s8B��_�3���}W�d�(��|�8�kiF���U�|Ơ�)�٦��>w��F�iY&	bQw����L�x��������l���_��s&���c�Iٷiǎ?6�M����"'N�?UUWr{R��d+����cēB]��k���Ae�-�(���D��߽!8a>8bL�Gާ*z��wR����rjϘ��
$;e��'��	�ƀx%� h��pnB�$�c8�0%�S�"������s�!v��[�\k�e_k�*���1,��LfB�"p��B/Σ���m�-��\4[1��_>�mUێ�_�_{}o�_��C�sp��j�e����1ƒ��6h��@���I��G6�^~�I�T'�i4�~?=q?q��v�����;cצ�ӢC��kC|&���UG��{>�R�J�*D����	4�̝J0>���p�SN��=c�f�b�m�<:3�����N�dO@��>$���%��U"��R�3奼�_b^'̄�kf��Pl��%������EUTs���e�|}I�8}�Z�@Ӱ��i�{4ϯ����_2T�焣	��n�1��^@QY��>)�d8�u�$1�"q0Z4Q�M�Zd4��ᗹ$$������$KѺɇ;&�$$٦$�h�Xh��L��Y���a0y!�.�W6�x��i����>t��<&�ӢCל1�Y	�u�M�[#�L�D�w�rf�%������1�]�޶nw��ұ��j6�!���ƭQ9�cۓ�:1�c�CGR'�k%���jZ�u$�d�L��>1�}=�沸�8�ezSl눻�Z���n�)���r�6��I����7%aLg��5��$�RU\���$����'���pYE�&[��*��Z*�w�:�|��p�%�N�;!4`��%�6�e(��rBK[:���N�G�&rd�k��{>:m�t��(�#GR�^���m۷&':0���-�f�Ǧ��M�(��<Y��ŧ�%�Z1UP���_H2�p��8|j��]K%^�vI�ew��G[+�R|W�كmD�����	*���ٍ��RA��7���1X��`+0��9JrC�&�<@0h:�B/nBI#4c	f�<Y�CE���p����p��0DN./!uq��k����$��"�c�*F����Q���d(�e)Ex�����SIN	GxQz-��@�g�|��G�F�i���m��6�K���\��N�&M����Rl�&Rr�";0�p��&ra6`,���Zn���*��_%���(�p�v��L��ĀĘ���f(C"�(I�U��AUJ�oOe���+	�,�G�h�i����(񇅦WI�%����:�E����"�t�YZӵ.ߌ%�8�{�N�=0Ѧ����X6�����j��x���k�Ǻ��}\V=i�[�lk�t�\�ܶV-�Yl�V��V-\Z��t����[v�|�W�|���q�S��:|ӥq~~i�z��c].7���Ʊ]1��V:��M�qk�j��������W5o���Zg���v��k��Պ²�_4�j�,�j��_+�i~Y��_8���+�⹋�,ǍL_�q+�~cm��=V��(�'�(�x��D�I0�/�\\a���cU�X���|�./��i~W�4�[|�+5���ˏ�b�x�����1X�:i��z�v�]+O�t��1x�������׫����p�ƱvƱq�I���x���G���Q��'jD驎���N./j�ڱ��m��K��WW�q�W�m�q��t�kK�1x�^./jŜc_�����t�0����[�3}���s~��DF��C�α�=�#��`�t�[��ظ�
�#on��K�i��f�Z�׬o�1A/�m�-�N#���[��
�mM��_͘���登��N����N�a�m�:-����CM��k�3u���˫U��c#�:.�9��.g�W��-D����v���fg��V�W������߯33Y����U{�����߯33Y����Uz��z�Z��32�3�ڮ�W�ΩӶ�O��8�ǎ<c�1�������������s�>ٱ�cēS� 	�u&��x���'UZx�5N4a�������5�䷉L1��6���|l�ti�&��^$�I��G|QQ$:U	����n~�7���&�_��p���dy ��y��bko��MO����!�YB`��H�'س�=��V�Oa�t�.��/IG�!Ip��Bd�HG�y�o�jູ��!L!?�6�m���������:񤿹UQ>2d��Yv�W RHQÅ�4Z|�8l�c��d,�,�f���<xL�O!u~�6��F�V���7�5����1�Xњ�4jkl|X�����.)���T$Hh�B�ZZ�>���y�1(��>>���m߶ж�.� ]�r����'3��Q��Y���Ν��m,�(t`��(���N�3��D\h3�C��r:���r�d���f�-9���H[��Hc2��
"a��>+Z�8l�D��ل��Ӱ��#����w�0�3�JK�0�Ld�\�����8�X�<6���,�?�<&�ӢC�NjH�횇CTkb�-+��>�Yo����4�K6B�Qv%=X��Up�]�DsI�mQ9h��6�o1�����'
��y�7eu64$�ď=�եϳ�r�gİvy����k%��4v��ݺa�GG{qH\Ddd�$(�h7��d�~�$�h�2�<<�RQ�8��1А�~0&�ZWͥ�d��!xM���LO�GnۚH��������I�蕷�a��tm8i5��Q��t��&9�0��@�`�����ϐ^⊇��*3dݟ9O;�
>̒u�a������:��2W+�;L��9'�;UU(�f�L��5��n��T3�E�jH��08��>��v��]�7YJ�30]/N��?pA��`x1����g��"K��+2�o>������i-�9���{��O8����;m�=v�㧏0DN�o$	BU~�r��A�	Q<``��� �0ైH���B0 �p�'�1=5���{�F�i��R�YO��ӃEg�d�3ΐ�I��S%�7)��=�>r��-�tkĳI���䐘8�4���f��r��x�O/���!/;��2���K�:�04Ӆ�S�`����W��O�>2��0z�e�����$�(�M��'�ġً7ZL�Mv�6�A��ph#�'��>Og���f��$r��N5bB!M2�M�<�\#�<=�'� ��6�M���h7iX�XY��k��k�q+�K�@t���,�&eJ!Zu���O(6�O�'��<m�n��o_<c�xD��!����=z�z�u�2��*�����J{�ɒ���sD��bq��y��$۪�56\�!�4f���/LI$��A����$���>%>�w������e�h��h]�}�uq�;-��M�"j�0D�&�N�rߞ6`���ˍe�&y����朜�r�r{<���S�(�i����)�p�x@�x�-5��!�A��O��/�9s��)8�~K4�&��K��!�hᇎ?<x�N�g7��cseќ���O�Q�NR����V��.~.:g�Q��b	 �	.q0��d��Ř;���L������A9���������Q�oj:dM���HۿY�nd�"�.�߹@#���#�-0�<��-�}�V�J�l�Ա���U��:[�����i�J�A��
-��L�۞���Ze�t���^%dzi�m3��.>J��t*�����b�#��d/FR�F/�)�g�<:C�v��j��lgNOU��6p���?6��<c�Ϟ1�~cׯ=W�?q�tޖ͈�
ш���L�����Z佷ݏ,ǜ�����k�t��["b4�U}z�H$�K�CFV���-��b�4h�RKIb�֘�3R���P�j��hQY��*y����s�w��i���΁j��tZE�u���n�˂c�͍���O&��. D��@N�5����f��O�ړ0�D)�d��!�� �� ��#��i���Ɛɤ��N4�;��y�cA�䆰<�>1��]!6da�v���&.�u�q9�p|�a���8ތ�<.I��%�m#³��}e'�NL�v8j�'IU�_��/ؼ���t�c��B���\�)}P�c�m���ǘw˂�x0~ }���k�ۚ��r�Ӄ�Ӈ箏��N1���z���c��x��:��2;՝�?=�׌V_��I�Is�0)8�><���$$�M�=3
��y2�N&'�J���XAٿ�
*�U��s_TI��f���m)9�	�<LSG��̞�2t�F�mN		;G%������%#��>���c�]�	�I�Ѕ�1��ً�Nl�f���Ui�<�y6x2g��4UUB��M�,rs��R|u�ᑆaI����0q,&�NRD���M�-�m�=t?=�����p�m��p�gMp���㧏�'N�+����N�ۚ6����m6�o1����|��q1'І2�a�R|�Kofi<a�}*���Q%��SRL;�GM�2�c��zM����fq1��⬐��9>�«�C�Չ�`�/��-��)ă�u�d���s:_:�ܩW�&kC���Z����l��F64{!�Q�|��X�
O&��Iɗ�%���ΐ�M��
L��y�S��ц�m�8�������x��'N�D�|��w�ꊪ*�����������S��㓮S��'�hzs�֦ÊB�U��I�1���Y��
�
1u3�HC����~ُS����'��h���m��L[�0�;ć����}��5�ǉZ�3�䌜|��G���^�D4���I�y������N7�Ke�!$�%�O&���a�Yd,rw���&-��G^/y���Κ�����}�q}cLf���<k�q����p�,²[X�X�Z���X�ZWK>Z��k���j�O���N>i����4�x�V�/M��X�K��\\~k����\q�m���:k��n�W�i�ո��<�]ۍv����XVK��b�aX�X�X�V[���x�oMNb�:\].;i���X�ˊ��������oͽ|��5��b�>kO��gˏZzƱ}c��/��aq�b�7�������b��ƪⱦ�V�����~c�lWk�5=^1��;cN1�K�ҽt�/J��k��b������|��;kK�x������q���X��Y����c^1���o��q{^�4��ⶬ]�i�q���4����kV�km�q����M��b����X���6v�J�8OW�TJ��pٙ�\�:�50+W���k�Ru��g�b`��1u��v;�a��[r�$H�	��T�H�=��\X�^������3�f�F2ֱ|�w�n�&��9hw�ז�L�������(�E�"	�1DY2L5�4�s&RU}�~�;M�� ���<9q���
��&#$Q��4�Y�[[ľ��6m����6���9��$��n�*$�T;]��@I�-x���������6N�w%ڦ��)r�����6�c���iZ�ws��n�B�Bk�M�4�m��Uۨ3��US���y��Bb{u��؏� s�q�����s�'n�F�հq�S�$�����?f��,�:�������{33����U��}����32�3�ڮ�W������32�3�ڮ�W��]߯333y������b��d(�tm��q�x��ǌc��׏;�q~r`����d8F��8�]�*�Y����a�;Z"n9x���𚇷\tv܎���� ��:�.=��a�˱����u�������[��'f�V��TQ:��S�E��X��kc2N������\rw���M�ヂ�����n���Kmd�jw�]���j<wc#قڥ�n�.�O$à��T��w�|�8G�}n���r�R@@ʤL
²��H��	�mݢ��[�q��v�Y�cv0��z�ˑ���<�gx˲�k��쓌h}��uێ���h���d���3��0��/����pGg�����r��]��g�GGgq���^+(��v�S���N$!²
���i @$r EO���i��y�=����^�kN9�h�����G^y�R�S�;n�4T�+ԧ�N�sϋ�9�=�;�B;�U�n�3�����/A��vH�X�w�[S"���˷3td$B�l�4k�E��g�f�`ϓdp����_dxu)�d��I����lh��$O����N6�1��K<5'��wR�T��O>�����q��kR#f̘,l�5��r�NH�!3�ee;�!&1>/fL3��q4w��e�j���֤��ְVef�n
��S���9�o�Q��:t�N0� �h��f/J��ٷiǎ;m���ǌc�4
޾������I�8�K��-.&�(tu2a�3�U���2�L�<=��2����)M���i��9~�3$�*��J0����u�BCN��L�p��+��ڑcQ}�}?*�XE�\>�u�k�8�0��,�BQX��7#�/{K�����9�'�80���һ�'!Բ�	�	c��IgN\��$y�%tC|�j��v�0�&͛~ٷn�!��af(��c�;|ǌc��׏'�-��9��2��!L���m��m�4�]Z�:�C�t58�ڒ}�H|�N}�c�?c��ʾT'Ɠ'����I��9h%�<�H�����kUuUS���vO�'^��d��ʁ�8��4ۦ���{8�X����m�u*���Ä���1�%K��e���Ni��Io�O�$������'�G�Hq8X���n���ܜ�N1^�?q[q�x�뷏�O<'�N����
*��QUEUT��n�h�m8v�ᆞL0{��W�Q��z��q=����0Y�%і7p�E����f<����;�L�N�9r�w��}�ɫ����|�o%6��ٔ�q9�nP����ߝyO�'Z;�	�i��iG3��d��������V|�Y3�䆽P�'.�Τd>t}UU_&���:�{{������m��(��i����1۷��1�z�=x��z���D�4!�<��㔅�Pō��X�Jnf˲�� ���*�d0�d򲺋b(X���ieO���|�m6�o1�b�:���A�[Kcp�� ���a�p�:���ha�n�N���Q��j��n������v��I��m���#Nc���<��R�2Y������26�Q�G�T��z�5��)��/��.�B���WWF/�E�x��/+t��:In_����C�M��J�h��Ã�pʜ0Ğ��U�e�n��;u
�r;��ǘ��h����՗w�ܽ�8<4{�L�=lßI�dtS@HQ�����������IG�����f�>^�?I�{8Y|�g&HuBGЯXp�ʳ��13*O%���`bd���Uk5����>��Ӯ��#���V�ڷ�����+����������Â��Ǆ����sv�Z����<sWI�gx����k�� �vzog��/u�W<��?y����*�隷�<`(tm�y,�	��	͸��.K2���!�|)r���I	)�{�1������ŤsC��zi:�t�I'`���%��8h�����|A�Δ�j�@����*�,QZ�8ԏs��L�^��T�(��<�g�G��tۧ+ÆK˔���O������r�a>)4����C[�B�GN���m�W��q\qӎ�:'	㧏Ǆ�Ӥɬ�F�Ԑ8oZ>V��M��X��b�EK9�UQ���M�[��&WYLa����6�ٶ�,�NN�������iUqs�	Ժ#��D���n��v������0��B�ɣ�K`��}ZçgO��*�T�E�O^��I��燰�>M0��%N�9'��ᢇex���O9~̇�$>4��Ҷ�����>�
���9>������o�6�y�G�����8��~|���c�1�Ǐ*����MkMkMkI�;7%2�x�����e�tӷ%�{��TX/|q�6��d@g;#�i�5�g2��1�F��O���^&Z%{�X���:0�5��BUJ�e��Q��]L�E2V<z}3_U�9��$�f��m��Ϙp�d�(��Ra�Z���v���<Jʞ>ˤ�tӇ��cO�>L�I2y0x�8��q�#e}��=�Ǎ��3���M��q\qۏ�c;x��Ǭc׏5��Z�����9���F0*�Ϭ@�$�q�Z�+#�p,&#��,�e���Úw���c�f�ú�H$�HqH�,�a��Ƕ�	]Om�av�� qv����:�U=s��g�ŷ;����]�=vu��t�q4GmB�����m�v��{{ޛ��8��^�'S	�#��:CN�-!9$\�RN%�O�dѣ�:x�<�s�Ii�=:L&�:7����+��!�_�M�\I��a"A�%���Op�)���`ї�ɇ�����o`��>��{���i�Za,��B��5�Ƒ�F9>��E�J������6�)�4Q�g�%����,��26D<�)>�Ԫ�!!��zjt��O8ڸӎ;qۏ�>v���Ǐ	��t��wD�S/��WtVsE˺'M�TUQUCG���a<}��[���>-J e1�-���&J!���n?'��>�9$5�.�T�
~����-�Ҁ�g�o.BByRq2x�ò��5��y�FK-�4���5�G�ܩ�wM�^
����Ij�B"�E%��o!�������k��Xu4��5��XHx�N�&X��z�����eB�8O�t6f�)m��`�|Q�:p��a���`���8lM�P� �;zzzm��V4�6���c��4AAB"'DN�D�"X��L:'���A(ADJ+�%��,D١�tL�tN��&	âaB&�8&8hABhD��ba���	��D�C=c�8�lq�1���SׯZz��"k$�M�܈�䈘"&���8&�%�f��%	OZW���g��U�Ͱƚclm��6x���8lN��4'�vz�y���`�O5�%cP�>n7��<��`�ѝ>�z%|�Zy��>�ṫg�v=}�gN�w�P�at̤�m��N�{��7dͷ;2�3����C��l��7l]%.���C�3��b��d�I�{�R����G*�i9)����)k|ӻ�w�{zAEk^�<PE���R��fW��|%�=�Vkϥ6'�K�v,\d�ҥŰ2R��[�X��\S�n�W�W�m�o��]]��~Է'V�sd�Ɨc����r�%@R��ָN���W��"�����#�b��衼�z�usuwHެ�5M"�9v8��B�,���1��=ꐇ�ٯ8!D�,���3V���<�V������{Qz0H�����|�Q,�����]̾��Ϡ�Y�wK��3���l0@��A�v�u���U]�Y��i�wm�n���p�^���f���o���E���q !��FX'��{}@��\���>=~��CN2�CZ�矟
��ֈ��V�\�V�~9���/_� �\�N��0FPq�����U�<�ǂ�Y��\�3�oz��S�n�����:���(C�O.���yw��F�^� �CRJׄ��$�w��WQ'�����Nv�c_f|��u��z���e��1;�,�u�U�Q�q�p�3��9��������g�j���V���~�fff�=�UmUڴ�~���337��Z�j�ե��ߵ�����{J���V��ç
,��j�N<t��1�1�Ǭc׍��D�;EUTUP�G���:��Za��V���l~3F�1,,ル�:q�Vx�<�:��:��{��|΍�9᳉" ������11,g���H$w��qUqzi\���L���6��@�J&�Oi4�S��c����P�*�Q�l� ф����ϒӾ&�É�^��FO7����w�*����-�Nt�~L�8Q�!��a�:q�<|Ǐ<c��z��~ �O���w��&
�E�X��N������d�k��I]$�8D�|���w����V�㑥d�iݍV+�㣻��	,��$����*��$�L����S-���Q�/���F�8h�%�G����h������HѴ�0�u1G�u�e�*�ɳeg��U#!���,�e�ߜ	���l�L��xф�ߺo}�;��I�X6u��{g����WG�hxCǡ)+$�o{�*B�����zwRI$�-�����Q��IF貏z���Ɯz��������c�|��������Y��^/^���&�t{43bх�uh�7v��2�ƁfD��d"�0�	��*1�dR6LL�S�#��ȭ�wp��X�I6�mc]��FU`�)AX�$�Cn���n;\r&g���V����u���zx���s�.+Dݮ!듻n��\�ܜ`��0��} T�?)�)�������I�>��<(�4}�_�W=�g�p��� �O�KI������PELTf�6��%�cUG;�����H��@p�[Cw����d�A�̺�h���9sE�},�8�SibC�@p���ēe�F��9�K�R�l�Ĵ��>H/���eT�#D��EW�?�(����9M���W��X�㦓�4�2C�J>"-��|&\��a���%0,�
0a��,�<t�㧏Ǆ�Ӳz���'�H6�I�X�m6�m&�Q���q)c!��7'=�پ����!�)�Q�m���$
7��0�]ӈ��-��cMO��~w�<�o�����;���f�����|Za�rXy��^�q{4�~��BF���.�$d��%���L�l�'X��(�M󌬄7DDAoG��9��גdۦ�f�1�U^6�Jw���O�>��DhɂQ�4��޻�����m�
Jy�J#E=��,8n�6p$�P��Q���n�x���Ɯxۧ�<~|��揇�����xh���Z�ww�z�z�K筰�<
(x��6��H$�H$�B�l���m(��3��ɕ÷46u��MOb�R��!W��ss�ɬ�n�W��`�Q�F��&�`�����x�'�ҍ�hl���w��.d��HIi�����x�A.�����b��90vk�2��m�N�4T�$�HGS+=��r?h���,8�������Ӑx�L|Pd�J3�I���`�)֋죗%]\���{��G=%�	��-�`��!�j�N:m��=|���c��^7�!��Z�ͽ��kݷP�"�����$9zp,C�ւH$�H6�u��ּW�d���+&�N�v�������ί��#O�.M@܁(`���J2!�
l6�)����;xa2�-)���=x�O2��e��n�UΒy��ΔKJo����I;i3=g���Б�����;'�#&>Jzٔ(4[I��ߓ�7�k��m�
�������hߔi�o�'Z
3~d0x����	��m�8Ӷ��^�'���4�n�6�4��;q��珞<c��zѠ�/�a�{t�ŷ�Ŏ�L�i!��"'
AKX&�S���ӱ�֠�#�bj1X>j���4�M��I����8�F���NG\ܽ����}���B
3^�m#V��ݮ6��'}��/���
��cq��ۇ��~M�<rD�FT<
�U;QF�-�7���=â#�\��2��l��`,P=��+Wi<|�93O�L��Y�I�f_$���e|���I���.x�U�̚���m�fR���Ifニ���M�I!&���A��Wai�IЧD8�3�	��V�Ur�RYe��V_kA��'�N&�l�N�cIE�����F�H$_���NY�V+řrq��8�)��f�Z8H��Uv������m<vq�q�����O�O�N�<xO�O��ڧ]����RO�H���Zm��m�Єԙ��|���!����fꪊ�\�IŅ,�O�0]7����Rt��}&��!g}��n�&̤|Go�K9d�gɌ�MѺ�Қ�d�>h6��1�g7���n@�Β�(�������t�J?}�9�����g߲�\�w+se�Xܣx��6L�S䇂�U?.�(���]'O��x|��!�Dl����/�`e>L��`B:xr�!'�}c��:��m۷�qÍ��8��O�1����1�z�=x��;�˦�Q0n7�5̘�x�H$�H;�s�J"E���c�0Sq�;~��m&���![Ή	�����d�/]�>�W7����x��I&k^����:��<UT�~O5�U_�{��E�V��c2ffJ��᥷��A��<@�vԪ�@v�<��+a*��A��YA�?&�2�ON�S�����Ĥ��g�	����0���%���}�j���*��L�>J(0|y7:�h��qÍ��8�N�|����N�<xO�G(����9TBUQF�kɶ�i��i4fОs��[��q�[˒�?K1��e�~�4�G��W @�vVg�Gۚ֓��/%��7(�L����G�=�?py��I�%|���Y����82Q����b`��S��'�߮6�_a��lq~�=���g"���9+��g����e2h�d�2t�\&�fύ:�Z[�x���sɆ��Lu54ұ���v����H��xM��E � ��hұ�1�6�1x�cj��艡0Ht��DK�&	�0zM�6h�A �"QG�4%������:'DL�a��H�:'M�"A,DD���6��4"X��0J�`�o\c1�o[V�cz��ׄ�0�@�N	���""t��8'�%�BP�%	Ddd�d,(A(�4&�M����g8x�0�����7�߬���3���R�&��?&���(��5EGM|m��Ϛ�I%�"��$���ɹ����MM�;��2��fm����,���CVF:g�G��F��I�"��=L����O4<���W�m�5���o�l����ϲU4�t�뀊�Vň���l�D9�'ڇ�=��`��G~�O��F_}$���׽�_g^�y�5=5��c��s5+�B}l̑#��A-F�^�S����Bgw��m�̂+�1�ްB��_j(�� ��7^w�j;���.��D2��}hi"E�M�8H�C
|E�ek�x���c?I��߬��TP�����M�m"��+��LU	�)J�#�t�=f��A��6	c$zf�<u�A�;�o]���޷]�ffsiU�Wj���������g��Uڭ�Kw�_�3339���Wj�����~�����{�U]�ڮ�p�e,,�(����,��ǌx�c�1�ǎ��盺���v�7�[@F�_]��׫OI�u�n6�(<'&�9�I\�m��bV,�����/Nݱɜt��r�c�u(\#u�ݻW�5-�qu���ܾ�s��u�Mٶ��6w&�,�֨�P���;*4�L'��o6��ĥ�]c��5�g�+��T������:籹��Q�w�:�6�<k3=k���h�m�l�ݪncl�{6oCC��uz��mr<��
�wU����Ӵ{�݇y�K^My��e�v�.�'��n�&5���]Qrv���������N��S�۷dyv9vi�c���� y+x!�*�/d9U�i�O&��+r]e�,�Z�D�H���^ߩ�sm6�kKb1��T�V9#��$�tݸ�[#kn\ۚ�V�krnDE�튖�gpnW��۷;KT��'/����\[���-v2۶��������d��)$�r�� ���4�g��Q���f�(�.�I	�ʄ%Um��a��E4�{g�'�Co\ٲ=Nт.H1���{5�'�a�Ӣ����H?��G}�	Z�|L�'R�c��yL$���e�i<q�U��$ta�B�]/�E�������kB4��[���D2�����f8�zr`�`ҙ$ߓ�a�F
J��z�G�e���[����w<v���M�8ڸӏ[t�f��O�N�<xO�N��;]�mԃ��A$@!�����Q���!�%��6`��K2u����Mp�>�O_��5�F��#���J:q)4���e�p��G3G�]�|�Y[��T� Nt�#�8����./mV�x���-��׋�QY,�+%��w���)�x�'k'�!�6Xa-)4�.g�\/��d�ǓX�7dL�Q�N�3�|�!����L�)���4l��Ɯv��n1��v��1�����cRT��4�0�f5��A$A$QI�g�6V��<�M'O���-;���3C+��8��Mi�飯��)�E�Q���T��U�˻���y�x��~o����l��MH��y�B�$�!k�_�"��/�9�>��HHL'tG�#w�,��I�z���Oa��iI�#<e�<Y��}7���L�$��͘a�̹����]��L�$)���ӱ�f"]'�C��Z�7���?4�7G��+���z����Lp�j�N:m�?=:~8x�Ǆ��8tr��~�Y�����6�m6�i��U..~>\ͯشZ1A�������N�w/R�6���#
~�܋�W�fŝ�ɟu$>!�RCˇt��NK,(�L&>>�p�Z%�>�4�6�v|PY�qe�D�$�Ag��j\��W�ƍ��;*��N��:t�d&)r��.�&�=!^�P�`|x��QG�����(vE�ܟB�L�1��0�p�i���%-e`�F�Wq�nݸ�����c�1뷀�!k��!�*���gh��S��N`
�<\iT�M���QR�7"%i��g��	 �	 ט+J&�Q�Ka���T�dM�v�kf��fum)Yw<[��:�an�X�������ѓ�>x���cT�uۍȘ�g���}��ބ7M��6��nc�0fs\��e<d�Zi���$<Rt���0x�"|k�fg�|E醎����<|�pɔ����,ǚ=���"a!��Px��UZ��*�ʻ��.2oS^���$']��6M¡�\^2�22�p�El���H�r�b�!Ǵ�!�i��%8>�|r�[F�u,��7��q�b���ʕ
�'�n��emY`�
�h_��G���^�$(��CAK0i�x�R_v��[W�#��om㧭>p�j�N=m�n޾c�Θ��=c�xΆ��A7��F;��{�w7���E�N�3z�nHb�< ��z��z_�;Ϊ��O�6�m6�h����Z�I$��:���Q��:_-<�p��e pى$���D�4�-��	Z,�VJ p����o&O�G�a�%�H>�i�N9߫Fߊ;�f�^�(v���w)񒍐�O�L��.-�3��9?&�d�Y~71�t����[L;ԭ��d�M@�M�%Zq��D<Yg�\��'�}$����-!�%!���o�%�H����n�,����ʪ��V�D�N��c���Ǎ?;8ڸӏv۷��<c�1�Xǯ��&�t��z(鋢���*�(�GQ������I��UB��<�4Y����K\n�=�K�	kd1�j�K�W&7m�L!��p�GXg�%mz$k��ƗW4�O�l�N)[�ޕY�d���%�D��l�l�����l�\��H6B��$4}K��9%W~�4F��ӥ�A�$;��Zr@��w�3=��UK3;�8G��c�~���[b����M�����[\�ʎ���y�x57�kR������UZ�x�S�S&�'�id:���JܔB:P�1�G��k?|�j�����a�F1�O8ڸӏͿ6��^>c��1���������]o[r���f���Som4#B��x*0 I���#8�0����F` F#���oi��ϗ<�m6�m&�<ME� 1LW�iuFu:�p���{;)7E�C�~��V.gF\qڭ�c��l�8˝�d�N;O��Xw�2a��.HM|Zx�βS��N�L\�I$܂��$��I�_�"�!VbB��T��Wm�<ے	��I&����u�J�F��~��~�
)�nӤ�!�A��̦Kv�r|[��/�Z܄���P}I��oX��6�4��޶����1��Ǆ��:aSu�sWA��@�2��
)$��$Rɭ9_]����a��K��fv;U���؊D�'ƛi��i5�h;�YƉ'3z�M�˄/FEt.�4ц���}���^ݻp���w[D�7s���q
IR!����o�W�c�w����5�Y�룾4e>�.�a��ԧi���s_J�/o���HGF1f�&ķF�:|Pt�L��&q��%IU��|���=|}`l���!��`4@��n�&S�����C�LCw3TPw9M'Ǜ�(!�[�M��G\�6�1�����W��u��9Rl�[��bQ���Gb;^���M���5A��!+'�^0<�<q�ڍN8���!���Wqᣆ��:~<a�Ǆ��:a�2��6��(��痶1�Xe�>�%EUTu��vRW[Z����S�?Xt˦�&R�t96���������M�6�k��M5Hi��!�V�kia�|v˺�Qwv_�M�?�ݒ��T�,;��>�y����0~#�3!ޔk�I�ѣ�BU|�>�n	�;�v���~6B4*��x��$���Rg2Pm�Q�0|l��?<x�DL6p؛4P�zzzzzz±UX��c,�e�x ��""&	҄ ��6"'N	�"'M��!�E � ���,�"hM�8pN��a����:'DD��D��:l��b"'D�0���$4&�K�&	�p���ĳGOQ���ǋ,���`�:hA �"'M��8"`��ӧ��6X�i�BP�%	D�:C�	D,(A(J4$6lD�ӆ�8"`�(����u><�a�>�O�i��ҹ�I��3I��!��^@\�\D����T�bF(l�a��E��v3Ӿx�L�;���n�L�|����\4b�h}i�L���=����OI��HZ4��s���O9�\�K���0'�LP��#���z����?dt�ޑ�W:��,���>�s3:��Wj�����~������Ԫ�U�]7w�zffffwޥUx��t�޽陙���z�U�Uo�:h��c���r�x�ǌc�1����zl�o
�TUQUA��4�6�ge!3F&�ٖ���M,��
�!�YpD�i�L��l����GX(��d���ٲ��������J��������Ҟ��C->t��3f����󿏞e+d��[�H[�4^J)8@ɶ���N���\&�x�J�k?}�'9P�:|��.S��_i��G$:i�N��'��l0Yҳo6�5�|m�o����?;c�|<4tR5Z"��0�=
 �	QUHb�*�p�ɔؚ"}��a���He�̟<�_�:C�'�j�u{Z�G3��̻�z�c�c76����`�(��t���R�κ䑙L�M�K0��'ک1zN�����4N;CD9�ΘO�䠳2HHd��`x�6��Py�|��7������݄c�<R����	���֌=Lg.9$K`>�}��|{�=��{<h�!��`��f���?0���x�0k��>���U�ф��,Ǌ��,z�Z1M<�!��"��Vn�tO���}�+����5��n/sjy>�$�H$�<I�"7}�Ts��x]Nxr%D�k,<�=g9�v�ɱ{�r�0UL���,��e��4ԈDi����A��k<��%�r�=�%9�uD�є�4�k��B&Ru�V6RW�9ӧQ>L��o>8��8����%���l(����|f���e;Ԙi(������SzM80�g��us�Ι��=��]�TY����̉wF����;T�M[O/���r��A�"�ۈ�b�����?gI9�>,�I�n{Gy�F�	
��w��h���YW'	�:~?<x��O	��t�9)ܺ�QF��T#�����*��}�>H�K [��\�qlUt�+�z�\�l���el˔�앴>ɣ	څh�w=	�iܼL%�i4�u�R�''M�1�^��B������^�x�L�VX���~�X�u�B9VZ$��g�!�l�z��I�:,p�N%��d2�<�a>`y��	$�z~$!�h�i5Cf��	*QK�[H���k��8ڸ�-鷭�������?1��x�0��j����r%*����dONe4߉�I���;-*��A�i�ܕ��ɴ����|X�g@=�DV�m�ɽ��ڔ�����szdי�K:]�d}���s9��`��L�}��[>p��d!6ߌ���L�0�m�_�8Re<�>O�|a6�N����.B��4�=I�FӉ&S���䲍�rh0Y�6���?1��?1���^?:�����ƌ�t�XUУuB��n���o�>{_�ﮞY�M۞)���c~9�����-5����;N]pM��հ�,P�^����۞a��ZϏX�qw���N���&�ϫdWj*��NRpyM���q�>ܫn}�x��F��=�*�����m�O�A�5�'��;xp���4QF�8wz�w���UD90|/�d�Awcen�N�w4��n��fRu6�:s�Fe�Ԓ3N��&Gf$�O�/�m�-�Ax�\$��I8`�L���O�t�W�>1�̯Olї��$fSGά0T�r�,q�"�X�-����xW�o�0�IгD,�����0L����lz�=x�~�G����^kE"j�� )�a�y>�)9��f���6pV�b��Bƚ��%o�H��͟+֛i��iD��m��n��񺵵����u�����u���i�1�즷.kP���x<c9���b&LxPR`��U���y�}�#fT;�����X�#Me�����e�~$��ro&���l4�鿥�WDi0�p�$#rI!d��[K�yܐ͐�1��(�4e�a���������d~H��!��2\����
4|}ӯǎ�Ot�2��F�i���}Xܗ��*<�I��j��A�I&�!��}�J%fvCM���IKd���LP`�έg{ ZK�,�s�.��i��~O�裥bL�W�6���?1��?1���^.����NMi��Q�M��M��̶�6{&��~�猳�|��_NL�[>>�Ӈ�i�̐�G�$�jݮ�RKX��R���)�
���_�
~*��ʽ=��%���H����@��Q4�h	ʣ��a8�a�I!$oe��4x᳎���.|Q�Ȼ�ȼ��Z���L\W�S�{+��{UUw$��$�4�O>+��4Bʹ:h�F`�<x��	��t�&����T�z<_(�����	H@"�zU%q<Z|c��4*����ڭ�|�W�� ��/ꘆ/�@Ǐ��}d<|I!4�����%���8�_��y-C�4�����*6�9,yc��LĚ��Q�,�S��L��V�Fz�s��#��ܱ�ٷ\l��>�dW3�b��`Ʈim/D�����f�}%��BB�'wɟ��O7i�tL��k��vu��8���Ƹ��x�����x��	��t�� y�{W�D��x�QUEUTQI;&��u�l4������^^8վ�Y-[d�j��m��[U�0���5��
��8�q��>O��!�zBBBBI�!�˳I�DLd�CI�IM&ր�x�Fpٓ��4��^�g�hz�2�t0;�OZSi�������C{��^�uUUP��F$O%��[mיm�dӦ޲5_�L�Um=-��5]~(�i,
ƾ��|l���bx����x��F�٢�A������+�1�]��N,����0N �D��""p؛f�AALE4"X�6"pN	�	��:��&	�`�I�"h�6P�0��"""'J��B%����'��M�f� �"&��ׯX�;~i�1X�8���~$0DD鳢pNX�hM	BP�A�N�C�,(A(J�f�M8p�Â&	�y��p����7�Bѧ3�U�T���Θ��t��q�"SFM7 �� ��e���AA5��G}�Ş��˳���>T�O�K�֪����E�V�?�oU�EA��A@�'r���'���!~zzr`A�&�ZE��XDD�[hJ��7�f���P֦�K[3��O{��G{{��F���U�nør��'^�2Ó�9�����d�t�D���4�
����om��H����jtus�c*9�1�h�rA����v=r�.c�%bqD���bC(��H�E����) �H�6݂M�Q�UP��dXҢ��j�,�0�������U�)*������\|u���LP=qx�]Lh�9�	��Gb%�˪^.mm���U�;��Z?�_�?����ff~��U^+�V���陙����UW��U����fffg��U^+�V�o{߶ffff{=Uz��ߎ4t�ae��4t�����~c=c�~��i�+-��3|n;��v���f��=[b���ԃ�HՌ?E�44U�ͭu�b��6M(�������m��ې�]<7?�v����9x�5�烧�r�8��]j��Ȏ�����
:�i� {��q�l�*K^H��%k�Z��Ni
�"ε�x��{k���vc�c��8�P
�#j�Ppqi1I����|���[�ծ����9���I��z��M�{��vQ��3<����9�m�v.��?}�3��[��;���U�;4��)7~wO��\\3\����.[����睉]n���pЌ�[�Co��%��'�����)�Gr���!�.ήш3m=3Q��rM)*��dK��4�@p���9�~�m:YWz���f�۵S/8Ĝ��ۛ�D.wW��;q��.�x:s�њ�����r �P�)5TD2�<(g\��4�<�Q��������Hl>W�4wGw'���HϏ/N%
$~�I�I/��یp�0|�Hmն|�|�q�Mi���S���t[��j���ӯ����!G،�%�}�m��D�ǟ���N����y+7��ޱeWN%<�e;I��M��M�(���P�!�$�v̟4Y��J㍱�8���׏���;z�=quN��2i�)�S>!�M��b��z��x�%�`v��L�I,��xgd�S�����F���;�fS�I���L�<�$�m���J)�jC��'��qE1k̶�{r������9�et�e@����8�_�U�Л
3���M��'�II&�a����>��x1�X��G��Ա�u<c��i\q�m�q��=x�?1�ޱ�^??)[M�uR�Ё�1��1<�6c)����*I'I��qV����ό-��6�ӻ|�'	$2�>Z���L���a��S�z����dŧ?F�6��ź���W0L���N�<��I�Ν��zy���>.��b�
��pi3��`x�!�̈́n����@��X��v�s��П���O��=l<D�y0����u4�\%Z�}N"e��p�E�,�`�0Y�GK��6'�	�>ɽX�1�J��ѨU�n�uh@�FqS�.�LM&JZn0�	�%xb�$��LH�������'2A	Ȳv�j�}�>���|��6~��x��~�}�vM�:G��%���N��/h�Q�Q${�>�>���|;/q��-2U�̥>��)��6�8,�b��NU{�&84����h��ǧD��%�x`�o	�-��u����R��Hg�x�$zH�5$���K�m�O'�m���Wm�o�a���?0��bx�0ɝ��}�SUDM�8e6/��Ղb��P�kW��{��)� �݋XJ���d�j鉎5��Lt���b�5Y��Ë-�tgyܼ���ktq�듍�3������n��9��wK�Ucڳ([^QX�+��*Q6��u�ջ�����/-��ɓ@Xi��Ǩ2�vI7D�������|��O�*��J��O��9����U�T���a9�6�9��t��0u������?q�Ժ����z�ku��$�:t-��&��:�Ǡ1 �2��Ը�ب��g�̗t��	*����B�e�gHy6h�v}ϟ�X��zj�#��ֻq��8�Y���tD���x�<xN�l�>ˑ���s����d�S[<��-'2�B<(e�����s�!�2��4���M����A �����W����Uw��d��ϓ�/�æ穣��)�.6�������\�:���	*�6�:��]���y��N'��H��5�#�jvV���"����{6f���5�Ҥ�(9(�<բ�snA7���ǽ����j4�dc��]8��������6�掘!ԣ!��2H�}ᄼc�ޜi\q���8��󷯘��:Ǆ�a2WQ���H�����_ǄK-�e4�=ʕA��Oϝ����xj5F>8�do�Ɍ�w1�	�2���􆀉0�e��?E,�cg�٣bZ��b�k9�[�%f��I��O)�����T����q�9��k䧩���g~���fo�MRx8�>NHd�i�.a䅽8O��CUP���h~�z>N'=ɢ͖t0R��n�x��ϝ�c��OXǯ��b�5O�BB@�Fz�)M9-�YۧI�A\�:�s�h�/WRYg#����$ ��?�q(��F/����y4e8LIF��a��5Χ�ܶb�q����t�w��Gᢂ	��?4i��'�5�W�]U\�%G&'�u:i���O����O}_�6� uȝ6;KrPp�Ύ4�8���8��ޱ��c��`�����pB���0��i�[-�#���h�d��ʝhql�.&�j�]"(�n
�l@�STӛ�ۺ��6@\7m�Ť
������Ts�	�Og�����p�?nP�kWe�`��.Q4N�2E:�o���m���u��KO��N�8t������т��%�^Oc�t|�\i�da������W9x�.R�,"m�I�Ng��
6����}��?s�ϟ�>%k��a�S6u2d�@���B6�;�~ t��[a�l��I�Ť��4�����c�OO�:~��t��m�i\q��ߜx���c���1����us}m�1ʵjӦG�Ա���'oUU�$M�a��;0`�t�W�]Y�p�m���ɳ��?;qe�ƍ�W_&�xk�U��a�m���y?$���X#Ҧ;��
��9�Z�q�@�=��w ��->0[�����_��ʹ�,:P{��x�
0����:"`��	��i�6�0�������X�m�t�N1ӌmX~z�^��0N ��"&�N�&�'M��6h�(AAB4Ȗ&�M���t�0�H�tD�:&	�0DD��:p�e�"""'JL���'rDD��ĳbpM�(�"CGr'DK8P�$�D8"'�<a��p��E�,��BP�%���N�A��	BP�$f�N�8lٱ�
�L��c���%�w��c���ܛ��yo_���C�#��`�����nG�C��h���7���^>���HpkƵ��{��ry�������/��A/��j�g|�McS�B�ӽ�ckq�S���tu"��p4+���M�]��ٙ�碪�V�[��|ffff{Ȫ�եV��������*��iU����fffg����ZUo�:h���!e�:h�gO8x��,O���4kTV�p����VGl�mk�콾��#��������!�dN��_��GϨ1�ŔE�޺�Ji�Y�]"�� �rb�Ӑ�c�(���Ѵɗ�$�I���0U[�ޤ�Bp&�Q����O���Y�&�;
��M�*�2u�Ƀ���.T�|��nSa�l���I�Q�Ӷ�z�Ӎ+�6�8����1�g�	��t��+zޫ9$�@�h��`Ӑ�&ܧL�h�Zk2(��q8>�62w>�;��Z��'�fL��/5'ɳ!�	��ak��{��So�ftn��ӈl��=S����N��~����>�Q*�&%@�m,�'\�ܟ2Y��D0a���q��c�������W k<���h�:K$�-T֐+Z�m�����B�"�%WI!�a2P����������'$Y%�nʺ�R�` $5Phj���6��qӯl��ݐ+�U]�Aͮ���"=�ܹ5��=c���RF�Y8'�C�;<q�z&e�G3����F���q6�Z�-g�3���~�ϗ�d�7%He��6y�N|`��(��I�{G���).N'R��[ \ĸ����4D��d�J�w��D�y8�{�p����{I�	��!��I���}��[�ʋ0�%A<�^b`��'�I�Ҳ�fن���7r_��|hѓxq�q�ߛv�ǯ]��~c����!��oI$��[4�L?y龜����cf���S⎽�	��v`��Q�'΂w)5�Թֵs�ZE����ŦӤ�O8�6����@�뛈"#R�'ُ$�d��8����o#Ῑ�$�0����n��W������gOY6�f��}�'_��럭�Ŝ}2�^4��o4�8�񣥘'㇄�	�g��+#��!����UsRI$6�<lO��ғ�Л8t�=J|��p�����UD٣e���O��-kɴ�����E�I�A��uR�~�bJ�;���CӜ⨖��'\U{��<�֗�T�:�.�u�R{�D>ɣM�-���U��/eO�a�_/���lw��ML	�Qt�}��-�$�G��K0��h�g[vq�q��6�ǯ�]�z��1�|<;͹G����ܴ��ύ;�����BK�7u�k�{ϙ$�C_��R��I:i���B�鄣�9�eRTK<3E������I��W�N����>�!��������⪷�6i-!�ohH��ζt޶���&\}ߟ=&�B����4v;J��˃~Kk]�_�M�p�!�۠����:�dm�n�m�gWm�n�t�㇄�	�g�±��-����6��5��X��S1,�Sk�Ƿ�:�8jj�хYD�Jk���Z }� 
k{ڒ �Ȭ%`��Ȥ���<TG���\]Y⚽q������ݢ�=z�[���ܝ����I�moc�����\P�t�FކZ��Qj�ゾ��z����|r��u铯^a��g�oL8�����p1t�$	!F8vc'��g��4���링�>:U�'��r�^�/㘨u2�(�s0�FB��ѫy��h���P�2��}�v�e[�&%V˒Qp�sT+�%�9����{��l�;���T|wgN�gMR��o~q�z�^=c���?<5���=l�c� o�ܩ�y�0orl�$h�Ri8�&l�q7�]H]���t�Y��d��N�Ni��'��ܐ��D6x�`�m�5�Y�K�⪪�ʫ�l��M$<|�揹|�
��M�s]j�DB�6�)j�ɛ�x����./�b��{AW�\_�U�˷߂;.1��桔��^LV!G(�����4��+�6�ߜ|��=x��z>t|:7�uy�����PH!:�s$�C�{���M']��$��<���|����`ټ�F�GJ/����������������]̸ג��q� A,'���y���n]8fׯ5���=|�Q��&&��̧��h��9�{�J;�POO}��mɤ��i2wq���<t<�6d�f�+�6�1��o��z�=co�~h�}�4ܛ��ʻ�@ ���\����pi�n	�#1�u4ssp�IWwb+����}�o�mΉ'�mO��ۣ}�	[�N�T%h�m�l�YǍ��a�P��\�M2l(�4p����sRT6ݼ8k�É�G���f�å98l�q;GN�y'�ۣ��J��!�I���4�L�<d��O���/�Ē�Z�o�[m��m�PI��ܟ������?�����?[,��� �����ԆC3�����:-��F�"ERB�%T%���Җ*�Ub�RU,R�U��T*�U��X��*�)UU,UP�X�UR�UIT�J�R�U
���X�T�K�U"�*�Ke*���V��X�UPX��R�U*����,UR�b��U,UR�b��UX�UR�Y*J�b���)U%Sz�*���UB�UU,�T,�R�*�e*��U*�R�K�b�R�R�*E�P�,�U)U,�*)Ue,�R�UKUT�B�,R�,�T��R�UBʕK�*&�*�����X�U,�J�(�J�*�*U,R�J������)b�R�R���VU��B�*��UT,T��TK)ޒ7EQe�T,�b�T�E���T��RʅT��K*������)b�UJ(U*�*R�b�R�U����J�ʅT��E�*��U"ʕK*�b�*�B�,�T��J�)�b�RʅT��T,�T��TiDԩT��P��R���Qb�YI-*%�Ie,�ZIe%�Ib��Dm�),JK�����)*JK�%��F�%���J�K��Y�QIQIaIQ��6�K)?۩%�J��RT����9�o�j�JUU�H��H�RYIe%JK
J),��������m)*RQIb��J���RQIb�U#E%�%��RQIi*RQIdRX�JF�J��),�K)(��IE%JJQ�#IIJJ��),),),��IE%����),��)*)*)*),JJ�J�IE%���K$��������RX�J��QIJJRYIdRP��RY�)(���XT�T(�(�E
,P�Ȣ��T�X�X(�EB�P��E���������EB��
,E(�QP��*E��P�H�P�H�b*Y"�%JJ��"�T�R��**QR�R�R�J��QRĩIR��IR�K$T�*T�(T��,�R�J�*T��`�P�P�EJ��,��J��)*XT�**EEJ��,�,*R���T�,��b�EK**TT��QR�JJ�"��T��b�EK)*X�`�QR,T��eJ��S0`�`� AZ1��T�J��T��,�IR��(�eK"�*J�IR��QR��T��eK�(�d�R�TT�R��T��EJ��EK*QR**Y**QR�J*X�(�QR��EJ*Y%J*TT��%J*Y%J*E%J*TT�*TT��EJ*X�(�(�QRȩQR��T��(�"�EJ�J��EK�EK
��,�H�)*RT��EK%K"�IR�JEQ��EKJ*X�QR�JJ�H�RT��XT�T�)(T�J�
��,EJ�H�T�R�T�R�J�K$R�K�H�
R)P�B�)b�
X��H�J�Y�R�JJT)IK�)%*)RR�����JQK������Rĥ%(��R���J�E%,)IK�JTR��
Y)QH�)IK$�E*JXR��
TR�"ĥ�R�Y)d)E*R�(�J5F��)QJ��JP��J�RR��d��R������JJX)QK!H�)B�)JQJR�*JY"�%"�,�R�R���R�*��R(R�,JX)RR�K$R�)�R*�KJ�*�E,�J�)�R(R�K	J�,E*��R�R��B�
T����%(���E)��)QJJT���J�,�J��RR��)JT��K"���J�H�)d���%*)aK�%,)B�QJ��%,)QK)JYJR�����X��J�Y)QJ�Y)%,R�X�E,R��IK�H�JJQJ)QK����E"��JQJ�����JTR��R(�E(��Y���K�)R��)R�)dR�(���R(����RȥIK����TR�*)e(�E,���%U�DjR�����K"�R��)JY�J�YJ�X��JJEE(���JY)b�R�Y��b�7�X�QTX�U�B�ER�%QTX�QTKUIb�I*�QTU)TNi�eK(�*�(�E�U)TUQT���e%R�T,��TX��T�U*��*��eU*�)UT,R��b�T(�)UT�J��b�UR�U
���U,R�J��UU,R��I���%�ٯ�O�R��Jv?�O�~� �"�� *(,`���%~I?G���y�������_��i����p?�_���?O����W��_��~o�G,�C�Ҍ�?�?-./�_��f�"������k������h�	�?���2����;����?������}��������QG��k��Q@�� J����~C���_����!������B��_��q���~��?�C���!���?�U ��B��O��_�	 i+��B��j�?w��p�-���ɵ��Ĥ��:o�1i�k��[��O����j~x?]�S̲B@?�m��h�JE (�Q�S0E@-��E��� Z�l$I�D�PI�R�Y�*-i��������Y��}������G�?�`$"Z*�A-B(�DEX�$���I [�'�w���[�q�1���R����?h?�=���� ���?�?���\������ T ����%����[�r��������^�G���~��!�J���~��M�a������a"��?C�@��ο'�������6��#�������������|W�~���鳧�C����DU 0O�*�(�����V+�'�7�f�]���C�������p�V�96�R����҂
9r���>%����ϑ��I$�������A�L�����)�B���JJ!��)��Dƃ�A�t�46F�`���b�8�v<�� �I��ߧ�_�W�F~�/4�� �2'���)��������?����߀�"�ҟ��-�����~��t��'������?�ܐS��!���?�����ø�� ~g��jO�Z���g��򪢀�������A��������/�c��,�����'�jWBZ�����-:t)��$េ�V��`3i���~@���>����p�A��}�*������#���DpB5�'�01�iC`:�;�~����>S�I�HV�`+ 6O�?�4)�~����������g�]�S����9O�xڈ
?�~i����?����������)��+�������O~�������)�����