BZh91AY&SY�e����߀py����߰����a��E� @zt      wv4 3      �4    @h P � �  ���`G�w >�   �q��]�ﻞ��QZۻv�w{��tWt:���3�mݟ}�����t9{pz��6]�m�lv�^�y����)v{��h���;��%�/b� �`:����Y�n�Zvޞ��zp�����۷�<{�u�k֯��w�3�sC�y��ۻy�����c�R�3��WY��n���>�Ut��{�{�׼:��z)ݎ�w{������|    xCW����]wf�t�-�ѳݣ�;��;�熽�Ά۽��o :��A��o:�����κ��/w=z1ۣ������l{�ݻ�^�N��  ��-���OO{���v����wg�l��^ Z�׺�>��۽�W8�o�|/}���y�����s)�{��{���{����Um��{�v�k��   1�{y��w�N�:{�ǽ�p��z7����L{oC}������ug{��{�r��g��چ�0�4��܊�=� (   J� J��@��P 5 � 
               ڀ�~�7�R�� �M0!�`M4i�dda)�P��@'��F��Q#��� �     '��)6�*4�@     H���SjaT���OhbI�MzFb�j@��R��#�2h0��?/�R	B�~��h��� By!�����$�&�D?�	��FD��/����s&5$U+�_���������q����O���c"�BmRu$I �Q����3-����Bq)'�%*1�e��h�"+�E���*9`�O�_������?��������Y[�:O�nWǌﲶh��D}r�C[��#�D�N���P�B�R�4�R'_�%���vW���D׵+�m�M���2�>�&�"s����ߥ�zW����~��u)�ʳC����R�4�R'_�"�U���Z����H���pM������7�W��H�})����9ٱ�����Uh���$�)�#��u]�eP���Rܫ�ۉ�xk�9�g��ܪ7�=�,yuIҏu������656jK�'&�����eh�x8Hp�A*>�"�6QL��*�%��؛}*ň�l���D�w*��ץ�jj�h��w��]�~��858'^�K;�n��ly�T#d�c�O�<u�~��A�Ò'u��%��U]j���A�_���W���>�e���܃r��}����sݍ�U�{^��o�|O�|o�7��p�7S�V����[����n<�ָ�kk�Pu���+�Fs����sqÕ�E寅�^*�K|�Q��u�WV��eU�rn;���^����zrMɩ+��=�})gNy���֥T���Cq9ǲ�=��Z�gN\N�N�I�B���:�N+����{�lܛ�7Sr<���5�}>�OU���Q5jM��5\'S�h�d���I�Ȟ����K�'��d�zOhK���l��lM��.�M�����D�Msd�]�������X�l�e�%=4_�9�ϴB	6��N���~��5��}�K����ݓ�op��|���w�����种�ІȔ��y ��ܞO>����Iv�<G�	�#$�C̓��d�Н�&�l��w�ѭ�K���a�&Sd�����	�(k�}��r}���C�y!�	+��$��4�6V�%�<=�p~�)�$K��n�-!ϒ��u�g�I�J���y�%���nG�Ic��"�l&�{��	gO%���:>8wBQԇ��K)�:,�~��'vO��"%�"x}�P��=a���(~�DN�"'���|�%"{iC�G�JtK8q�>FB"Mt��D�bI�lJ�DJDF���=��N�?tN"%�
�"GD��D��{�K7f��Bw�,�L'�N�&�"'z�ZN�'['NvO��I����"%u"%):h����DF�?iX�Oi"Y�� ���҄KM�?"D��.$��%��):$D�d��Ĉ��D�$��x����u�DS��I�i�:�;������h�R&��"HX���:G��4$�	m����'�!�N�"#b�i�8'-%���-<j�����(G����u:WgNvt�D��㳵::�,߄jY�l�C�A�Nh{��6xu,M�F5,槎�p�ħU(��w��F����M�hw>N�P�Ћ ���#�s��<q��5Z��p���+��m:�O'���ޏN�m�U��:l�/�<T��yQ�Wb6����K�¶z�j#���<pu<]�]O옜��٦a��Na����ޛ�9Ȝ�S��:w�O������\�o�:jl�$5����NNNq9�UG��TO��G^���lAg��Z��I/CQ4i�@A��n�'M������3�#*�&�5UA9=S�uU�#"tt����E�D��G�Q;b:9��Ʒ��#���"t�AUv�&֥	���S��Y��K<;��Һ��Igd��I�����U���R��Z� ��:i�J�����"oMJ ��#�TD_T�u%�SDO�U,��v�'���j|��U�ͭJ�jp�s��U5�b3u;����5(�'Ȏ�Q}R�e�D�ڜ �|���.�ɳGH�">�DV�{��ki]I�5:r��ۃ�k�n�;�n�ϑ���B��|w�h�iJ;B7(�	C�C�C�M	�����%����ӣޕB>�>#^��ȍ5,��=S�w�M�Ϡ����w6k�ϑ���^�8�5$#�܏C��C8�;�v6��=�D<qM��TG�rK7�ڞ�D�O�F��J�N��[��J�ݵ6'Tῼh�p��ѩ��Ό�Ր�V3���%�*�Cx���N�{q�c��=�{���}�V�x���1b<�gs\л<��M���Y[��{��x��Dn�{��6K6K,�r��{ڏ�����Sʕr{�W>��4H�=�]��}u �����J�jx����_F�Qg45/^*��Ur�I�8��W�ǒ������ҧ���R->5�T�ġ�Y�}��^.k��ӓrN�����7��9;�ޥ�\��$wꦇ��{vf�욑9Q����xOSS�,�5;S��7ٽ2OUC����=U8k�vNI��{��n�A�M��U{R[�U�_5�j�����y׾���»���9�� ;$yj��c~����ړ�SS�4r���MvNzMĩiQ�O�'d�|����uQ���#qe��,��d���u��%��'��������l�<q���6X���q��$�}ϝ�:%�͎����.��W��}Ƣ'��DD�>�c���� ��R'���}�c�W��ep��&�N�DNܓd��D�����8:ԯ�#Q(��K��'H#�$��T�G������+biܤN����UV��W�����Y���������S��ʡ�������%7��|��ի�߫��ℋ/P?]�~�g+􍫤4�B(��Ac�y�Y�d(q����B�i��ۜ�8C1��=�xe)1�#H_,�h�3��O^挣� ��]�JCA��������8�� `�7��8ӣ�� �B>$���"�iG�-�H38� �#!�N������!A�n�h�3� ���������_!��1?�i/[�3�0����^B�C4�(��qnk�M�4�BN�#D"�B(�����d� ���(B.���)��RJ������1w��ゐ(�?�������:qƔe�C|���!�	��*ؿ�>�4҈B)G���h!� �G��4�qA�l.�c A~܄� {���)�@y�QD1�D"Er���v{�M
d!��ܧ��ΆƆ ��zi�dy��PE4�~���xz�<!?�BE�*ۢPes�8#M!��8ќH�3L� �E)��8�'�8n��A��W#xR�� j�SkbJ��BB~Q�Q���)�#���z!���Q��A�)򘦱��4�yM���Rѐ� �"�h�(�h�C�\�l8�ER���C#d*��ʍ(h�iL��oOC�2�e��c8��.MI�=A���!A�!o�=��)���1���Zxh"��Ǥ��i�d
12���1!?B�#ӽӷ��n�nNNh�}��|���BO�D��ISx�L{4�Z��V?��b�G�<;�4AÓ��~���͓�/����$E�N��E�%��'�d����"��<���D_�<K�y4}I�-ix�n��J�?W7Xƈ��K��K�ry�{����-7�E�O<6�_)����ϓE�d�~O�����|{��?����RF�y�!7êI���qt��=��<��K=��H��~^opH�GM�ٞmZ1�T*��F6���$?��V_����W�z��*.\��DoLy�D�޶2�8Ģj�Jr���)G;��_/T��!��:캳�Q��fXr�tZt���&�Ak�8]���Vt�x<v��E�8��"L�}�龺��G�DE�"w��{��eN��)�&��3v��}=��'�����Ʀ�p��z�k=�{��ײض�t~#�t�,�`���g�Ῐ����'���ݧ�y��TF��[1C�ĳ�����7����g�Y+*��&Na��S,�b���ѿ��C~����c�iٕ^\�K��Hnl-y��yY{=�{�";x}�_�6n�i-�p{�owl�
ՙ��1
�{���d����5����M�p��,�^�/ql8�C^�#�S�>���(_���A�ƙ����&��W����ϯ�|w9X�}��r�}1t-G�yg�BBVo�9���������^w���,e�������}��i�����W#ݤ�m�t��t����N�OMT���'���\�D�kDC��>+�p����G)�<����P��Ek%��(}s���?P���]b�Kމ��O��t~7�(�{=�wM)׍���cka��<���7�ѽ����j��VNGv���
Ѫ���$z�wA���F���������nyǛ�I��̻�7P��1��9s�H#���ɣlo�ٻ���Hu#��K�۹��;��v����R�sŧ{I4�IQ献��~<s�N�_i%=�?w+����,��i�W�Z}�m�!*�|����>;�>��K���Rύ����/����o��Mh�N8��C�bV��>�}�����1���u�=.�#��Bx��5�x�E�b���/�<�c6�/r���o��I�dc�Hyb�����V>G���g�w�(͈q���)��{O<dw� �$��7Y�H��˼oY��;$;�u�����i�y��)��B���߅�^�6O�_��o�9援��t��~�Q�����j�]�\%������9�����#��'��>��4���]̾�ąt��ǒ�b���x�\Oa}��/J�����M�x��V3�!��<�ɞFO�S_������s�I�'�=eh�Y��ë�c�s�Ʃ"=�Rn/yxuv�	�G	ԋ�:;�Y����<��G	�7s���=&��Ty�-D�|������ֆ�y�l�NM�ea�;��q�L�{�z=���	���<��^����e�]��}�WI/G��J����j}^uN�7N�{�*��J��Y['�7ᇕ��ZU�MQyК˺N� �Čo�tr~�[��S�N�k��m��mG�y�Z����[e��Ӆ�)m�,���z���\ƅ�<zN���^?2y��p��s���ד�#�������݆�7��n��[F�ٓ��M�}��Qc=�GMk:*jSÓ/B<���O<ch�(�]�W�/]+��I�ϼ>������D���!D/����pqD1��̩��4�h�}��`��q���$���!,��(�O����T����d����7�~��?W�ש��W��u?#���	�ޒ7���G�,Ą%�r�
%RU~�?�}�!$��a�1�i��6�D�AP��C�Sȍ��o��H�[��׫��E�׻R�q��6�5k���_Y>�3|ؒ!�g����9r�F�[ڣ�O���M�M_lė�άm�;���'�q��S����<�.�)�/x�c��~����^���Y��ڮ�y�ӻ��?^�y�x�/�=�ۤQ���xy+l_����:�����b��$�֟xʏ���}Ig8����Ȗ[:�IT�5��k�-u��)Q(�����U�δ5��8�V-M!
:�{s5mx��Z���.���v�jIK^�'a��,�d����K̷��^ʂ�W�j���wiFR�J)�$#��k�b�x�%��W����߻H�%�_	��{�.��9���y���"=l=D����<^GuN-��ID�!c�[k^�������}��!�d�G�[դ]s�u�M'ϑ[���^����Y�K�7�O\$�,q��_��f�����'���.�=��n���!#�t���X����>����_I9�9�l61���̝\Icit����=���f�����aVr-�v̈���<rN��[�!O!�-(�kcJ{��u�Z�uius��)Y<�W�>�2��f.���/|���������M.���F�G��F��d�->�&VX�J1��-���ܻ�k��	7V�D��g�I(�d ��Uh�h��s��%��Zٲ���Uvq\����Q;�p�N�Grk��MS�8��I�QR����'PՅJ�P�h�%��6�IL��1X�Ic-K�4�6-z���ۃJ[]n�+��'E+Uڣ����E���"��V�o��[T���[F�h����F�#�ޛ�n��nͪ49V9iR�\��Yi�%���G��Ge��iD���R"��܃W$��lN�,i��+�E�A6��F�q"��]lRY�R8�Q�6�$F숍���j��dQ�I]��S�����$űb�$���&)X��'\�Ȳ\D��/8�K��${[I7%i��)n'�{7�ϙ�3J�^
Q(Վ1C��,WZ�R���bv�*�8���lS��=ka����W�wh��Jl��ɣ%|�r�T�h�.	K,�2�NW�g5sNA�M�r.��p�4ّT�b���լ�����H��B$��dKd�Í�4X�u֪����+v�".�Ò�����Y&H�n���M7-Ier	
�e�Bbw-r8�Sv�Q$���bjD5i���@}-�Ƿ�C�:�&9��NGQ$ IBښR�Q��iTԙ"Q�~{�֦"&������Bj� Pb_n:�~�ʣ��p���D⃂j�+���t4M���b+J�F[e��M�ZhJ��;R؉"{Io���8�Ѭ~}�y�O�ez�V����������h�㌲�U�rj/��W"ђ�ǕW~��>���B��G���+,�7�$��BGv�p��!K�4�7�#��@�u��F֨�ύ}�F��1�����ɤM�M
4OwR�S�ފ�%w�{o)"n.m�H�RցD���o��Ŗʭ!_��1MI̬����Q�}2|�b�i7TK5�6�RvKV��DLԶM���-�֢��Uy�.�G֍���D��{K枺{M ��Ywe-�Q�q�f�N�v��6}9s����7�HNi�Ȋ�#{�6֭�'%,�Z�\�������Dm$�%/�ԗ���~{;R/��K{��XЕ���튴�eQDܑ���E�wD�����'����|�����C����}�(��{�='߁��D�O�.����)�����O������!���������_ňH�Q(�ş��g����{�������ZUWȪ��������U[bҪ�t��UҪ�Wj�U^�UU�iU_*�Uz�*��iU_+J��U�եU[���]�UV֖EN���{��U$��	�QD$@���-l�F֤YZB��q�*�j���5^���}k�U��W��UҪ�ZUW�Umb��������lU|��U��t��U^*�Ux��Wj�]��Uv��ZU[n�t���*��t�*��Yb�����5>���	H�P*���"�Kb�����h�b���O��n�@@�����_v�J��ZUU�Ҫ�Wj��^*�Ux��UꮕW�UmUUU�U^E^*��iUW�J��ZUU�Ҫ�WJ�U^���WkU����گQdU�{����-D�!$Da�dډJ��Kc`f����O��ffb�*��*��*���U_-*��t��UҪ�Wj��^*�Uz�UV�UU�*��*��**��������Uګ�UW��WJ��U^*�]4��描�(�e踐ږb�63����%�nH�^\����[r\�#m�o]��cF��V�Ur���FY�2�X\�j(-���r�x]-j�"U�&WVj�� ʊ��)1]6�2��l�=���~��N��j��B)������U���P��?g�Ȯ��~�����L�'�K,O���!�A�4&��B'N�tM��lK<"X�%��,DD��D�D�bpDDN ��BxD��D�blM�� �����B�B"pDKIb'M�lM��BhJ!�BA6	���"&���h�Bh��t�DD���Q>9{����_	�ن՘)��!p����*�~(�
ɉ�҈��JD�E�4"oHJ\�!�DF,�i
�"A�Q��A(����&8"`�,p�u��QH<�.��.3�D\���Dq���am�E�B�Tet�Pe�-��5"D.�#�J8��dU%�?Qݛ���E���1Y�,�щI���4�4DJI������'-�V�G��q@�Bi#(�(��	��V%c�:������Y
�!�4�,F!���!�M�*&=���@ҺL-\*�uLM�b�Cqh�f��/��F�4Lf�B�ZɎ!DL�)���d~��p�4~�hn�Y�zfq���K�H�AW�j+G��NQƬ�!DԶ��^���-L��J���j%-�(&�Ԯ�dqXK\D�0�W�%�mlm�q��w"�M�!��I���[R����*BE�y$��q�C���cEmLc�Iw^�l�ԭYRM��B����yI��Q�j����R����y��~L֋6R��cP�޴l�V���9���r�z���*����g����w��f���*�9�|�{��a���������{��f*����g��}�����6Y��l�:`�bX��ͼ:Cd4x�"�!FǓDR�ʨ�pd��Bq;#(,�1Q�eTl�2:.(1���b�§X���j�Rʱ�Dڳ%Ww"N$�S�)�V�Htln��L�In`1���D4�!��Ȅ�-�`���C*�4l�����!\
qc
��>�Udˤ�Cc������d)�
vٿ�o!�Ӂؘ8�n�"MC�Tr���Zg�����1��A�A:J��"��PԸ�I<�.]�3Ly�i�S�>��w�t��F���g�â"X�t�Ӂ¹�YV��I$���o�y[4:~lt�p�2�|FM�UK�0����UN�'=	���gA�x��v:`|6lp�����UK�J���:ݮ��3[<*V�¶VU�:FA���i�.�Ӆ�`��Gǉ�����LX��/S��q�)�6'�舖%��,m	�IH2�	GTԒI#�=&zɊ�4h�l���ˑ��$�JNSA��l��ѽ�.æ�̨��ɘf�jU���X�r��V�8����4ĆƛI���%��%039��<4m�ɿ�d6<q�>.N��#��$�}r�~d$8�|؜x|CF�4&�0æ�%��,=��U�$��AA�X�.Gd3��V�4��~8�#K#l��%�3�!
(��8��$�ѣ����ʅ�cfP���p�;u�I�ý��v��r��V�K>M�f����s���H�[�e��rIэN���G�6t���bX��^=p�De2&J8� ��T�"ˏM�$�U5̫Ж�pD�4iM%��B�BQ�,W+,#C#i�we�1��:�ńX�nb,)r���C�A����h���b���+Br��Z���E�J�+Q�$�c���\���-{k��Ic�H3U�6T��D$�HȲ��G��X�Pm{���v�LE��tXh#L+�7f3&t3� ��F���!2���Iw*��0�d/���i��2t�%��I����pԖ��d:���v���e���!m���,����;"U�����LYI��&�r`�#c�2Ybh�:"%�bxK�.}��I!a�ǃ����f�rITt�RV�ƍꘛv�Hl::nۗ6`���ْLJ�}w�n�gI4�٠���d$#84f߶;�ƃ�(�<�!���	��[a�6�XU��8��;%j!B��f7<��⸫���W���ʧ�m����ó$$,����;������GMl�tDK��i�l�H�E^ԒIq���r[f�A�����2Cu(�]6��x�xs�ĩ�ێ-t��_sSF�"�k%X���6K ~3�}���pl�����m��p����X��ni�a�C�z��<��i��c!�<[s�b��샑���fc1���֮AS?v��J��i�i��^BܗNr�F�t٣6%��,K�_Ƴ;�{m��^W̵��9��xv�Z�%j�S+¸��#]$D�!E�ܫ�7)�0D��BI��.B:2���7��8IQ�a�ˤ���hYX{�'R).�IeB������������D�J=���C=�!I��
����ɑ��q�>>>�� �4l��fY�,K�zf|��=*��"(�$,Gt��4FJtIH����&6d��e����6J�6�?ȓ7�وD�iZ�ݢ�Ķc��Z$А�h���$z��#�-���Kmˉ����X�x��$�aH ���m�GcF*�BO}���9����
6t�䄧$�h��qN}��1�z��G�IUM8a�lㆋI��%�^�����:M����\t!��XSXt��Yd�ȂII$���m<~l�6��
+\�h$J�0��:hM�btDK��	�I\�I!�!BU����-�j`��ox��M�:<����X���{$�S�r��%v�Hm��Zt��8��(06SM��(b�aѢ+&$ʩI^GeV%G��L�Kx�˒�!ń���F�g�:o�\����v�Ys_\�շq�el��Ғ�Yc��<����
�a,ʓ��`�au'L+�9:;�.�˸���'�]Ļ�ܫ�ex��b�\]���یq]/�8��nN/��x�'���}U�
(Å���J0�0J0�0�aXDY<a�TL&�_��~?���O��8|=%��C�:#�tzL^+��{g�?4��?+������gÄ���a.N���	�t��gǌ��x��v�^�����t�L2�V&T��k�QG	�jL쉓�K��:K'KdI���*�r���d�]�K�wq����+���Lv��q�+igY0����=�='O�鳥���(��n���ŝ8y���^��~>���]lۋ�~N/{�~�f��Ԍb�r���E�g]�ײ���oS=��k��9���~����]����32ffffc�b����332f+��ᙙ���s33&b��ᙙ���}�}�x��<l���0æ%�bxK0�9�]�UTJ���t�F����Ԓ��F
e�$i ~e�r@x��Уl^��bu�v|IV�X�yP����'j~ol�X�?mȲ���M(z�������r��d��#³*|U���&J9^ҍ�m�|1���6Z��[�p�$����ے�015���|��\�,iz�4���<6Ӧ�.�d[bh���t�&���ի&Gϭ�U�h6VK'��W�&9-�5+凱~i_�t۶�m���=x���o\8�[L⪫�����W�\8H�`0m%#����
db� c����LAl�ẸF��������~-_��ݸ6�4Ŕ�+G�T��[M�hB9#��$����}V�%`y�������Jc�����L
��2'u�zd}+�9)?J0��>S��I�J�>z�lZ�L��(L���!ы0����6x��ؘa�ı<%�Lz���i�l{�#J��#yTPh�&�#��K���7$n�J�B���D�kpKa�6V�ԓ�AAj		2�#�񿟕w��$kyd�&8�!*�U��VE���c�(܆���UUQeBxh����hM%ESwnf��RѢ
�������Mh�ȸ����<��L44�a<�̖}H��qn�̇J��K%K#1m�Ɍ,�=,{�\{(2Üh��v�$�6��@���t@��L8q�l�kͦ�%U٠4�1�eH�h~rG�`�C)#.#FB	�>|Wh�I(��], �.DId�.$E!Y.��#oYO�}�$�6@���e1�����vR�ʲ��G�TU�^1��6�n�z��ێ>z���ӆ�W���˳'UTJB�P�m��bpP'�LC�T<`� xb�21o�21K(���;���+u(4��Z!���a�nj*�WS3�M��0�T�U��	rT�� f��{f�	��N�|@x���'M�&��,m�#�y���-�:Oĥ��|��:!)ä68 c4ܶTݖ��۰i��b<Ċ,K��(#�W�����W���+��c�:C�E�۶P��RӛOSo������Z���t�1V���C����M�m���:p�ÇN��۪>�����#�z�$�4���;� �0�"�ҹ*c�b��X�LTt�������I�WvJ�i�J6|c�Z��L�����!�I#�Qe�"��r�D2��oCi���0����A��
r��4�ں�?J�Xon�I�L��;�jsz�&Xt��UB'k��*�_��|0�A:m̩ZJv?vm�VXz�:WK#�J�O
����W��o��n*�}X�OR�@�B%+�������̔p�f��������O�`�"'��HI&UeUR��Ji%Cf�;.����0�z���U:)�W��K�� � b)�|p�0k$>�mL�n�vieHV�3I��fc1e`x����\�¾)ܯ�79mmՓ[e��&�fL|��a��h���a⻔vS�$�p�zW�n6W��Դ|����j�ħt�����T�����YcSX�;LmFK���ⶮ��U]�k�����C$SLB4�z՘}�}��'��e�tO�O�X��ӆ�U{<�A!ub3+ �	^���Fj1�AM��ِ��G�[%*���)���=��m �Q���$5�&ni��*�LM�5�	��J&9$k�6��J�۶���Z+T���z^4]���M{���W���!=hj�f�^qY�f�Y HҎ�0��r�ӓ�|5ό��'��GU�V��y4�(ڭJSM-�\*���9�q� �a����yd�,N��iq�I����{m\�:RYR�eubi]�;9Z�m�`z�0䌱,�;�&�q	���IPM�LTL�ùa�]%O�b�%Na�V���[�ڵ{j}:�<cq��6~?,æab"xKu͚z���![>�aaҶ&�_k� �ОA�M����$	�rIn@��V��=[��ҭ��pϖv�G�ddt`�L	�?n���c���'~z�0u�-��頫vd)�>?�L���=A�]�><XB�X��l�8��d��`�A~m�q�D �CТ�0c��I�ِ�8A�i�ێ=g Cf�,�g�Θ'L0��D�5EJ*�7�/����^�s�04WN��nJ �Ǖ[�Y���,00|�����!�%f�?&̔2�.����Rl�|Xw�,�2�0���Q�+�ٍ�����a�nB���[��D6\��˶�΁��9�>$vt����6�%�9qNކGl,�f��!;&c%L �:;2;6ɷZˀɒY��6'��a����,,���O��UUX$
�-�ݳu���`A`O3��8�h����HHېpC;02B�5��!��L<�=�Cl!�2�[qc�Cj�!�NNL:�ڿ{�M&����;J�g�sZɳ���]�8g��s���-U[kj�ˣ�э�iO�iC�o_���HI'Z�D3�kX��	��h�!R�	)��N=�>:>��4M�O[J�<~3o��>]>g�g�L(�	���jaXN�V��$�`��n1ی�[]/�9-���n2��Y�����v��b�\]���m�N+���Y�'��q���"t��(�epM%}�I�Ya
�	�$��l¡0�C8����x�^/�2�f/���V'*V�x�!�L(I��\W��3�^����/���_�X������\^/���~^;f/	��хa0�XaXA&$�Q��tN�a�0�'��|6C���g�̛����1U�՜Z�/K�����q\Y��^��W���g�1�mt�V��g��x�^N������˨�bB0����l�eD �8�B(ƈ1�!���zU�z�i�7�� 1�ܤ!F�(���TQ~B���37M4� �� ��6Z�!0!	�C00�!���S!�d��?f�t��E�;�vw�+��n��æ�F���[�[XE���=�z������v�MG�ˬ���ն��D���z�zx/2��iCc�ؙ&XFX��b,X�'~GV�&�g)��11"i
�Q��(h�4w(�h����φ�r�6RR�Y��rb)�h����@�ȩ��GD1!�J/��lkg���h�~�it�q:L#/��W�Ąj��4Q��YM�r��i2b�FI�(�p�H���q�\�1�A��x�bf��܆�B���<�#��5�����"d*b��^rMz����>���m��V���.OgNse�!��$U:����Cm��(ċ���q�D�#j�VU��&�,ll_�ޱ-��DWT$cR�im��v�Yec�4�8�6mJ��X�¸%m�L�Պ��q9$n�B����ywr�Y�xi�nݪ5��,��6����+m�r"P�*��U���OƧ=.1����-O�M$8䷖����U�Tvj�7��3��w߻��g�U�2�39��s���̬U_,s3;�s���̬U_,W3��9�fffR��X���;b�i�n�mێ�q�8�����L@���<�4D����:m*�"���D\�(�m���k4�}�<��Wu8YV�.�D-�#�X+D��V����	�{<�5hF��5e�r%5편��l���˗-�Tg���&���M܄��+q&��U���Y�֪"[f����!��Q*A%�[�JJɊ6�m<�j㛆����1�2�4������ԜM��Gi�;~L2v�q�\���b���=�cv�KW<8�I���m�.��'���ǋv�}>��z�W���d�	A�'Y��p>����e�g#Th`�h[�l��R��'��i�N�tr/�\i��eo��tw����s��K��ܡ�MV xs�:�~�I:Ϗ ���6t��ǌ0��D��eN�v�UZ@�T9RUX)�vڞ�'��I�Gs����˭5����⏾���	L��'C������:@�����k&�~�ϒ���ͧ&N����O��~�F�p�E8�m�vWKM�||�N�1����B���I$i�e�dl,����=h0}����J�kao�!a���A;�/g�!��fΛ6Y�L?0�0D��]�|k5�*��$�N�ރEg�q��(��l���ʢBV��'4��|���=[M�?NN��P��ʭ�`����FzZb-K�U�s��Q%��F�#���P�u>����F��t������ڝl�ӳDES�Zh6@�y�V��BB1���G:v�j����4�ܶN����'�<j�:
>�'���r4x�~{;����f�ٳ���a��"xKx��5'n����ЉH}��*�l�������]�00,aA�͹P#�!�3Sk6mx��
Cq�Ttp9|4"�4l�<�tB��Ue\v8�̸2���=Du>z�k�H���tpӥ��!��������Ɯr�N�apx(N�_���M1��$-޽��t��]E���~��,���=��A䣤�����2`��&>:~0�����Xs��Ї!�	@���SJSQMP�&,)Jɍe)���c!r�eXA�R��EE%O���5�L�D#:1A�2\K�)X�p2]�~9�d�.d_f��d,DԺ��n*Wv�nk��A)�Ƕ�UtC�m��x3M*5�C�x)��S)�,��FG��̛z��Tσ�[u��������uXe WF�m��ځ�!K��J�ޝ������h,�^9m��x����r9��y>����M=q<9��;<Ty�c5R��V��:x��K��b4��H1���,p�)p����Z₋� ��{����|a��A�����Gmh�q��C�Λ,�g����O	a���� =�UV��)��փ�|6���$&���p���8qۊ�Of6:uޕ!ZG�w��s��Ke��i�r�:���鰠Ֆ1���0���G��D�4``�A�r<6QpŘ�1��.���n�k��x!,�#�%ǉ쩎�8u��U>��|V��=woð(����wF�f�:RW�/i���//&n�y<6��N�N��w&6��m���0���0�0�<%�M�֝M��q�|���$�I��IR�X:�8��i��ٶy���>�C	ADZw��[�X[�{#!����Ev6%��L���ef��\���H$.w-� �w�\f�>�Q�y�pS=�<-Ξ-�Z�rv�n�,'��r��3�Nؿ\��[�3IVd5`Q�,���6�"r��Y2�����3��ʛ*l�Ě�IA���e���v�?'�gN3*�W��eba��C09��j�Xw��I��!��<x���N�Ǐ�&a�,=ϴI�,e��2��UUhH04V�]`th,����$����}�d7c��We`$OM�"5х���ф.�XP��Kc�UnZ��)
�.�B1[��5U�%Ӧ������4�|9wփ���C���}!�n6�W#\! p�M!��xV���3��z�3���܄���$��M��m�]���58�3I����7��ΫC٩�G����~�*��&Fz�n�X�r�5�x��C��1�l,*&�CC��6h؛?	���<~0�0�X{T���H&%�b%�����!�q�.7n+���f����Q��r���+C���QiW?���%ƽTy++G6IF�kC|l)M(��g�������bD�uM����N$��Z�(�V�A\,x7��h�Kb���m���b4�!$Ȓ���A��RG��B��Am�˰����1����?=���7�M�N��.'#�@P����]�ߟ�J,mJ���UF�A:~|9�p�t�6g��f��*��oc:ӷ��=s��zS?z~=eGйM!��9(�I��Jp���1����}�;>
���m�o�f��춞w�Mc6��*vڽx�o�z��o�q��:zt�C�A�ܒ�K�Q�����Пn���u��R��zCIM4��AЁ�[�[�x�g��q�r:�L0Ӹ�V���sf�,2T�Y��6�{�����p={n���*���I6�.�����G����A��7"d�E���	.�6e$����l$�[v�	��3μ��iЛ^��r00D�����d�!�y�Z"�x���E�6Hd�}=R��F����"L&	FzJ���&����K��t��8rz]�U�iX�Y�ڸ�&�c�:^+|\q\_q|^+��\_����l��"C	dL+l��	�aՐ�6aP�aXMV���^/��*�q�i\Wg���p��a2H�S$�}��W�p���4M�2	:C��N��/����_�>k��:c��������a0�0�I�\ºjI�p�t٩&a:K썓��t��Ή�.K�N���<�.�]ļ�ǉ��qgqz~c՟����,��V�	�ta��O�rt�ΏI�c���h��=�����}�X�5���\do�Q�!��.H�K�Ω�(�z<@mxzW�,�<�*=^/Dj=z����C1�5�Z&`�f-��*���N��7d�JI���}N�Y q�3`r���B��}��\�^�<I�|@�gq���UW�s��9���*�劼��9����J�Պ�Ü�333*�U�y�(�N�:p���p��`�a��,9���CUUF��ꪫBT<�O@�*L�V��¸A��L�����Xx>]岼�Fi�ǅ�48!������l�.��)>�-��bh��I�$�Ɩ鵶YZ��zu��co��k�������%�K��\��`C#I� �)���$��vT;&]���̄�r\��m8t�o�#F�#?Kj�q=�ں���o�{e�᳧�d�f��<l�����ӧN:t�鰻�$Ɨ9�UV��kf�we�[���Y����64ių�; |6�ezi�!!ər�IR�T���**�jI�{G�WJ��VR9���lf����ϺIgr'��ԙv��8����{;6���{����'F%|h��eU�{V
4a
�â��=>��C��Q�|��A�����h��F�C�`q�e���i2�-)ޞ+�M;v���ߟ��~q��8����N�v�jecs]:d�ҩ�ҋd%x��Z\z�D�Õ��ۇe� �F��i����$���#���P��� �j�D1H�"��{��Z�J��u�J�Sƞ1�{
%6�cIlǚ�"���6�m�G&s,O�I�Y$1ud.�d:i��{��$�$��rIL��b٨9r�i����>M�~-]�NKk����=������n����'��
0�Sࡇ�fFϘ�g͵���˖��:9;�u��G��}h��0�hm\��3AeSg,�!M0�{K*ܼ&Kb����\�J���S�:$!a�6��VI���"$�U�m;t���o��qǮ8�\|y�7���u�;��z� �3"���+f\A«2��V��bB���E/4cpd�nѐ�j�V����EtַSco ��*�P	� �k�UUhL���·�8χ��H7��r�lr8��qga� \�B��44.	u�v�6���e���m�ڐa.�2�\Te��R�"\�ō���7Kq�����H�h��M���rdHJ%!�`�kR�2A��rز	p�HԱ-�.��$��$.*]KBT!#�l�섴H�]�q�	�.ۄK�.��(�\j�&Za%��X�l�KdBHLQ$�Ɣ�PK��`Аbr�M�R#��X�#�T�[�M���BS)��H{HSiíV�q媶էf��,�b=p��������sn{)\��v�K%_�`�,��>ӅQL�f�#� �~f�ಘ����9,x����J�c��`|y Q�'Yo�N�J�,,���CfBA������
!�6x��:Y�����g�:l���I��}UUhM�=cQ���Ed�1�a�$r>`Q�|���htG��g�Ϳ��Äg���m#�����,tp����WH0Є���r�M�?r�֨;]�ћ��(�e2���㦝|�0��+�VV�EQ��U��	Gm��5Xt<
"	s���p��������;J0�F�4G����hx6�9#!�'F���Zx�Ý�:CE�E�a����Y�af	Q=L�T�ԫ�B����В���H%t��#�̿�6��
nܶ�l����p�Z����q;�4YU�ݙ&��Q!��4��`���1���I��s"�p��ݕV��٠��<�)xg[��|��h�d���,�`塁P(�d᳹,�ga�sK���c�&��-�hǇʺ��~N<4|�;�mN���:䐪����4���x<yn�ݏ=#�����E�:xN��ǌ0��0�0O�F�c(���!7�B��(Y
�yZB�ň�F��I~D^���Ȳ҄%i�G	挍!�b?q*.���2Q�(��1�#>D�sRmZ�bM8%^[��L��r9�F�B�c��̮uUm�Dh�+C7e*�*���6�U\�1V�O�:�O���ݹO�!h�>#�4?���p'.v�!���9r��m���t���1���8k�U(!Ka���e?SԈr.�u���Y2���͈�!J�
�C�ݕ���:7hxp���i��!�cTv�"�R6J�� �,����X9��*�4⟾���'�|?cF\��(~rrby�ߟKf��n��M8ӏv'��`�a�`�Fh��7EoD���.��UV��ӵ4U��@�U�f�m�t�8Q$��*�0�3���C���J��=(��B�PM.&�ˈ�	�	�?����%�x9)��(��$|�d<BM�!P!Q�a��2a^<�g�ϒ�a���lht�``p�cDB/ш"GT�L��0�0���H?u��!�����L���Jl�����#N�Í9�|��t��F'D��`�a�M�9D��C�E%s�UV���X�t�V��i>!�FTKv��x(0�!��
/C��#OJ#'8e�I2&N���`/�
�����<C*.�,dJ1��9v�9l�C�w�0�r;+p��F�}�$�p�~J�3��I)�m!PԢ�W}���с�gŐ�B�`ۑ��Z|���%6�bΆC�"m4�q����j�=:�c���!�f�ƄO����a�a�YfD.�HFڪ�Bz	^�te2�.� �m��H�?/�g�u�^�꺪��[�+FQ	�|5�f�	C	ONHuL���a�]�YWG5M��òI��a��D鐠�^17::r�
\<UU��>v����O�.ߍ2�۸.O����k�T�����zN	�ΏƇ	���a"t�FR`�wĮɅuf�K¸W
��-W
����U�+J�c��/K7����g��q|^+�z����J,���"aVO���h��`��ROd0"aXMa+	�J���q}Wkū�q��l���/�a0�RL'Ʌ$:a_a;&l�+���x�&/�q�+n3����:<0zN��:=dzC��zts�V$J�	�ae}�a8a]8Q��:x5gG	�Y:X�6=,��'rܓ�OYzĽb{'��/[�˵����|Y�j���|�ƥV�ì�E�I���\~/���6o�N�����
m L�p�-Y]�47#(�A
Q	��C#�H"�B� ʄ�)e(��i���Lx�2C�K���B(9^;��A(���"BEr!I�)�G��P�!�RE&�iS4pf�p�s�d67�"�4��Bb��F$�&��yTW`��+�!J<e�TQ\�H���o��o-��on�w4z1-�I����+p�@�x�JCE��4n��v�5�.#T�3EJ5jǔ����rn�1�(�sݢ��IH5�ٚ*V=`��F�A\�Q�#'�J9�"6��{
$���TJ�Ws��w4��EJ���)#���9�q2��<�kQ1A�e�^�Pbi��4�1̹��c �J�IG��T�]6���j��#X�l�J�2�+h����A=%����(����i=�f���V<yP!�T��>�r-8Z��T}M��۾����ɀ!�o��&�ڢp���"ɾ-�ol��k^��TU@�r�[]�F�M�icr�CQ�Wd�nƩ`�	�ZvA"V9ED���lI�[[�)]����)Z�*�-V�"[r�w�z�������~Y��71%kJ8��k��1���n��B���B�4�m(�2�'&4�rȕ�Z��h�w(��آ���G��!*�U��RL��X��%+�UZkcf��a-e��(�ܟG+o��$s+���(����s[�P#�����9��J��i^s9�ffff�W�Ҽ��s�����U괯9��33336��ZW�8Q�4t��0�0��0��5�6#�V2�g��(�dD&$Ѣ��U�XR�HJ�	��)����
Cn�X�Acb4c��R�>�Q.q�ui��;j�;H��kI/Z�d��Yt�=�UUZNV6pB	����hNB�k�2�E��%4{Z�	D��``�N�La$�� Y�;�eʻ2��Й8}-�8=%||��$I�����$O�ZRs�>z�ۣ�BI$�p�8z4{)��m���z�i���1?�'�16�4�D�����B(1D<���\r-��ʅ�"�h��S)��0���ӆ��`�Ӻ.ǣp����,�M�BagO���`�&6l��w⪫BY*A��f�WG��.����=%J����ۇo�P��*q���C�w���X�.�>i�{�l����$p�`�M���24$,�n�Xb���<���l��b��T[�i�u�d�Ӧ8�$�������u9]:��aɆܘ�;d�0t���re��nry��U[Sh�C����
!�e�,���G���:p�çM��NHv^OUTTX����	4Qʫ]�t���E������5R��$!#C��t�q����N��xl��g�&�+�)��]�Q3\�ڻZeK!x��~�|��|,�h�,8`���d���-�Ĳ�-�'�َ�S�\��A��;�.����*X|gg	׼�Gdj�����M???8r<�B�ÇB�0z�a��X�o����<�ĥc�x���a���`�x�,���Z4K���UUPMHH^�8B)�Y���pi���D	���MZ`@��[:C�E<�42�QdK`���f*�!$�<�*�W�8�m?m�uX���D�f-6�ba�N�~���1;��iv�J�;��.b�X�Ž��I��[���|�:|�u�hrj�UN	0�rӐ��k���,r��.̖Kt��1�i�O�=x����q��<:tٰ�,F˳�ҳf���&X:!ȑ2Ddb��SP�lDڂ��
A�����F,Y9U��L���6ϙ.-ho`�xVm�ǔ��Y�V��z�OT'��$Q��bF�k�ʢֆ�lmD�89a�n-T{�m<������m�gp��P�vI
8�m�2)s!JG.nxcϡ�gƐ<#�`�%U9���ӷ��ӑ�Ѵ��\[g�nzl�]�m�V8O�XlÉga���>�܎������?i�0��>�$�+,c֨4`2����Ce�����[�O�����nh�\\�n�dU�O\�t�q4��e��̙<����?N�[Uj��c��Ӧ�4���~<a�	��0��N�Z�5UUUUAFt2�x�}��BQ��[T�%=lޟ���e�K^��<m�<l�OK���x�>_�pO���N��ö�����x�*��Q�:��eb��y��I'�%�����mWctD��+jt���?�s�l~�?=��)�m�m�M�14���Z
u�k!m�6���=2��|�~z9x�x4YD4h���>2tOǌ0�0��,�25�I Q�ʥUPO�@�J���aR�Ugn��}бm���4��}�R�
j:bS:}a���<x���5+�у7I�W��4�ͻH[hܛ�:SѩO�R�S0����$|�u@*���s����R^E�2��R3 Ռ�1�L�F����������$9Ƥ��V��%Upu��:�ī��!�DI���N�}�oó��B���9<x��|Y�㟉�0����2O�SUUUJ�p��}���e�Ks�4��(v��a�4��t�y*-;q�9�eB������"�?�j�,j3ehE�n�L�NN�y��o����G!�t�$�IY08��CN�������h��G$a�E1c��O��ƀ�ҟx�G<C���e���?c����k9:|�8�}�r�'%��紷���X��	�X4l�,�0N�a�0L0K,��p���g�, �51������b
J��T&��Wp�Si4��4���R��]��\�ci�iaA�����4o��lH�),��lu��"+Su�˖	��J��F�m����v1�-y]��%�<�nY���-6q��=h!��t;w+h:p���e,�$��O�V���2~�ӳ��_9_*�f*Q��t;�Pa��LZ ۑ�맰3�h�_8v,c����#��mĐ�=�6e��<8���|ǣ��ׅ�4����}��06_&s� �0���C�K; Z�8�d�d�S��!�jp���M�I����ݶ<�n2Q�E�,�g�x��,��BMS�a㊪����p��9%BH�*�AMq��6A����A��C�`d�Cm�dق��%QR����1�>����\�4��Aƞ<>��b�Dv��[�8��g��!���n=�������15��"��J��\�=K;����,2~ګ�7,���O0�������T�����9t�!N�5���K8,��a�:"X�Μ8' � �X��B�bhM��:'D�ı,ı,KıĲ�<lCb"hDD���B�Dٱ�"Yb,�pDؚblК �"&�DO'�"A6"'DK�ObpМ6�f�ؔ%�J "A
؉�4"p��<!��l�x��0�?������wq�ȿm��8^{2!���p��6U����m�׎i�߾y�����(ƿ.��%��_���;O����WM�&�/��{�ٻ�����ֹ��Ux�+�o9����ͪ�V��7��ffff�^*�y�o9�����U⮗���(��G�0æ0�Ŗc}���UUUUT��$c�8``������G�d�
l�-�X��)��U0��CЂQA�c0ӆ?0r��|����!<�e�,��!Kr�F��J+��L��l�[(�r62+I�u����J�2�=1f�3ۘn#DtǏB�ٲ�Q��U�]a���9�dd}�3չp0?Xؙ7C���$a!J��l�%!��	E�>S�6[@���n*�~$��c叜�4`���h�0�`�`�,��9�UP���,�\UUPF�*�+�$�Th�s���L�ǅYkKO~q�Z����q�U�5ȫpD �6ܺ�+��������Mr�x4G^����2[-���p0!Ѥ������|oMW���w?h���rF���S�<�A�
J��!*�a�X����ǩR�r��m��4�~v���&'K,�9�BY�p�61B�(Њ�B�d#(HcoV5��\v����At��o�����7:˞L�<ӫF�yF�(��x̨���q5X��j��P�N��R�gK�w��C6]��|��ꪪ�h��Z\-��T1�b������	g{��.G�Jٮs=�gE���>p:`���:���9i���CA��1���Shlh6F�-t�!L������E4�-�������(m�������3K���u9*z�b<vv�]4ƕ��e�±�u�H����H����cA��s�h-�|Ph�=}�|��*�σ/N(��Ζp��G�>>>:t���fͅ����e4y�ʲ��HI�ja�����g^���#�϶6����b+�2�ߥSF��C5�j���4;쑒6|�¡�(��CX���|��-�r���-�j&�����3s�����Rd`Q����q�l>2�|0)�t02���`Q���16��'�p۳VnD��,���βXd�U�ߚ(#��G����]��ߡ'���P�d���z	i����E�	�vp=�p���Bh��0L0N�6Jٷ˻���nkV����_���6C,x?!!$$lLym~l>>�a��9$�C�ܩV4�j�'Iǆ߲ؽ��q1;Х<��G#M4�8^��TM��=݉�u�D�4�B��Rh�tė+���I��D�g/���I#!��<\���JD�̌v=pHI	1��n�l���-'MCI�.�V����yz��I���4���bS'p�=L'���۩�Wo��O�q��o��>q��N�4lٞ�/�u�qUUA2��c����%Qw�Au�jt��:$3L�h��e���< ����D��z՗Y��lo�h�ѹ	(i�Dy#cg�0�``��a̐�hx$CAc��F�ql N��|�;a�M��f,�9:[JUWH��#m�a0h�2m�ۀۀ��m�X�|C6Y�͟4~:"a�a�p��}�I&�}E} G��
11��tҐ�b+P�DC���^ݻP�{�F+'`5P��A�q9Q
S��\����gA����(�E���Uȟ���ղQ�KZtc
�vݺ���%+heJ�;��1;��N����m�eӑ�8��1���NI`�V&�$�"��CUZq˼R�EH��r�T�K�^i������X�~��q��(%S��vVZ{�_�!ۉ�d�Z=g̕
[>o���ßy�h�Y��N-4GC�#M<z6:�w����u�G͝<��m��m4h�$�N��B�,��T�݈�h���y"eI���^8}[ԨC��HQ8'�Ee~pÃ烷�χd4Q�h���tâ&&',�[�UU�t�yXl,4x��>-�D�*�WtK.6��������n�������K�2<���sۼ3��X����`u���SA��~xdv�U���t�<5>^����Ǯ+�����K4���k-"Չ�"!TJRG�ρ�xgä`tlܐ�#n��Y��ہ��$//���`���+%_�pD���r�=M��I餬t�o|�����v�ÇN:p�f͞MgL22�*��AI�>��nQ��>hlx0q���<�O9\/�fz{݋�	h�y&Ӟ��qJ�~xⷭ�Mִ�
��B�]�!��x�t��,6ivI,wǣ���r=�l|�I�u�������S���e����������&&��񸭳+8�M_C��(�#�ٓh���<'O�DD�0�6Yf��2CW\6�ޯ=�UUPh�W_a�������ųz��m4q�}O%=dۥ�X�l�e!�9�x4���I����-�dm�j�KmK����M����,�d�F�m2�p�{d����1����g� |Lȓ��!2:=�1�HI�#�ˆ��J�C���&D�9r? lx9�G�N�P�:Y&\Nh4z�`�����o��m��������o�=|D�,���p�B � �"Q@�&�؛8%��xO	g���bX�ň�"%��
 �"P���Ƅ ��bxD�B"Y�bhM��Bh�2DD؈��Ƅ�H"&Έ�,DN��8&�$M�6lN	BQ:H'Ȑ��AN쉱��Y�6h��B�q�q�Ʊ��i�m4�4q�i�B��J�1dZRB���R�2����ضѬ�VT򐆴,�@�!���KZZ,�F���k�FR�Q8
�k!F��l.�ʋ�̓gFw����*�B�Ar���Ðb�}�D��[��5LLif������A��,F�7��r��*V=�
���$ǐg�f��_���R������Ѷz��,B���T��Q��1L��'Ð������h鐅L����$�%�n�tܪ���B�K�}�MA�B�-�ǝ�O� �*���U�6 �+dE1����Į4��o�)'-��z��^1\x�S8�A��
2"-g�S��1��k�'�L4(�CJ~�X��@�e5/׿]"9.l��O��������<�W�z�qk$�Jt�naཾw��99��\vTϼ�~���ʦ&�%�հk]py
#��ܲR*��iG�kPJ�H�IamP���%Ԥk]+I
Ԕ���"Cu��Z�br��j�wY[rldCy�Y6=IU*v��(1H�q�G�e�2#�RE[��TK$�t��rX҂YP��v7.������B�W�r]��mQ���u��{t���\R,l�M�Z�QUZ��p���ϳ��*�WK�sy�������t��7������*�WK�sy�������t��Ҋ:t��GDN��0L0M�_�7��a2��H1�2"�r����J��&WU�j�]�D2�B�2��iD�HA�ಷ�)IUq��*��u�ȝ��n'dQ��w���V�yW����	f �\!cuv6�b��WK�4h�-��-��ocr��9h2W�q�d-�ё����r8�Àɮ�q�*��t���ޒ����G��V�����JR�+�>�6zJ��TSEi�
i��;�V�6[X��d!+�x��"�t|�O��g�,Ha��R(��nH�����/�D�f��~0��0L0M�,�^�UT�	�n�Z����`C�$��2#A����0��t�>[l_�i�W�b���~6v�4>:Y���]U��������е�oBX�/�9q�,��%�%�d�:ꍕ�X�
�3�{\��i�!���<�m���:�t�C�^�v0�jv(�F̖t���:`�,�G�'v^��F�疪���PkҴm$u^I8Wͺ����<L>{���E8�~l��΋��4l7:c�>�^��M9+ǎ�v��YHB�´lh�V4�IL��'���y�q���ߏ/'��~�~?~_՘�f2�A�0<�#,2x#A�o=�&�G���׆)�t�3=Ծ�)k���%O���Z��Q$	�ّh7���gs��z�Ov���;~|��Ν:p��u~p�k8�����8Sa�����K��g��OX�X��d�s#q�NB
3�\�g%:�ck��&�l���&�%4���4٭���g�*�����Λ*�A��fٱӐ���A�����ʪ�=�t>,hho#����q��ܿ?/�P��W��+f�nl���><x���4�N�8�xD�0�<h���B�C���)��EȌxC\P�^���f�T��#����<�c묹�m�D�w�ę1�ɪ�m��
o�;5��AÐ�~��8O�5cuJ�IF����=�bM"7Y(����H�4l��5��UUT�ˍ�R��,Ilb��1�d	
��)2����d
;�Y�x!	l��gc��<��댁��I�:�v�0����p������}��t��jP�;����I��5�FBV��&$��dD�q��%UeՄ�#O��0�C�cca�������Gpᣦ�0æ	��çK6s�Ês��ܫ1��UUT(�ч��� d�d,6�A�]lx04�
'���#������h�G�����Um�y�m8����h}�2|m4�ݖxĽ�^39Nxp�b�I�r��A,M�^&ݖ�>NC��0ҝ'�Z�8�)����>�LևA���h�%�x!:�H6=blx��FJ,ᣆ��~:`�,L0O,�XT+���b���B����Ve�pv��x�����*�69��>y���d�F�`(�B`��D��x�,�D%�P����U���a��"JVD�%*xW��*�l��N��j�5�
�*1`��Db�ı���1&�q�D!��zi���tlb$�
T)P��v��rD���յ�YSbyXҪ(�XY`�[F����.DQ�t�����8��eiZ�+y�C@�1	$��LM�J�eq"���DC窵V�UH��%�1cI�bC5�؄���Ȕ�<��0i�jH%���As4����D�h�je�bȒ�O�v�),uՒF��iW��!���Ȉ��V�U�YZD�r��*�mc!?���tq<���>l��4u;4���M.%�B���2��8�)��?��4x鳧N<|t�g
C�j�a�y�a��"0���bA�YCP\@�Lj�\BI���.��6�)�RN�-C}����Z5��t���]-�X��l-��5Dʓ.��d7d֐�@��<UUPJ�%oʕ$�����:f�$i�|��2(��'7Q!e���D�&7-���S��nYc��ya�������O���n=zZ�:��I���d����ƃ!�9� H�M[mя7�i�f<��<��W����|�튵��i11=J����f�L:`�,L0O,�B�}�(�cXA���J��4b�`�X����T[pL�㒉�Hx0�VM8D@�I�ج!g=3pb��y ���P�ʖR-Lո�$��MjT����nr�j���m��2���m�̅��1VL���tM���n_M�����h��٧}��p��I���������q�á�ym�W'�'�;T�njm89� �\9�h,�]�HG(�hv��Y�����4t���nCI	:T��(��Oqb�,��>6b��ۤ��U��>���bh�G��DO�'����W��!y��Fd��UU�n�HwfC���L�/�2��a����M�M����(e4>�`��ǹ�J�~��Ul1��4@�Ё	�+����m�>��\��0]zv7(�,��2��W�Xc	%1��7�|�]CN2'����WgGM˹��:R��t�*̸�6{;�'[�oX���|��n8�`�a�%�(��4P� � ��P�dЛ8'N�ӥ�I�<%�b"X�%�bX��%��J!b&�DО6hA(M��$,N��6&�6hMD�"lDDnD�B�舜6"tD�,N��6&�2i%	�g��	�	�����G�N��Y��lن��8�n8��or��o+���9N8�p�Hz[Si�d���n���3mG�*)�ٻ�z� ?G�*t��p�{�Z��̗aPF��w��SU�;y��$݉喒ڴ-�-���{mZ��ř��kF�֊׵^����Y��lz�x�0�w�����I�9���߿x��s33��U��s������Ϋ�Wo9�o33333:��]��9������|����(���GM:"xD�0�<h�K�����ge<ҥ��5�B����g��.ce��Q*����$$2˰�x4Q�Hl��r����%�Йs&½Oq)KZEhIxgN3r�x6�|�pk�!��J��v���4?oנE~�~�3A֣d�:�'�ö������3�0�o�m8{74��5o�8�Ǐ��>x��g��=,��=�y�ar׾⪪��~�L3zm�p:�G#L,(���� ~JQ5"x���X��	E#I��LHys�&~�sz=^��<]2��p����C���xl$$�w�:~^����>;9��_�xv�Aڿ��l�	]�4Y����	���?��Ӿ�
�Q�ː�F1�<G���Xk ���l�Rc�!�Ei(�+ �!JVA2���(�'��:2�d5�"���e�����w�&ye+��2�!q�*�YdMISlc�s$IId�c-CĨ���m��a��H0G3�-�\��S�u2�Q�l4�n�r���!����?����:���-UO%�❥4�eC�8�eJ��x���`h6�CЕMm�Cn��Ck Ӏ˒,������(�?:�a��<T�Q��]Yo��h�P�t��vV��=��0��0����c�:�	U#d�,d�,Bn(�)�r;���0�|�ˁɣ5*!��0�[��hOtD��ba�x�fW<��g�qUUC���3��*�= Be#��\tl:��F�ua���VϬD�v�J,f���	d&'^&+�˕���8� �$��9�Ye^�n]�=�������G�:M:u�oC �x�$;*Q����n�E��7e���hMcD���k����!�3���-����V�?����۠�A��Un?*՞����:�֞4�����ǄKƋ3йm���UUUUT�N�G
�R�e��$F\���,M��4i�c����2T��>����|u��J}��{�Ҷ�K���k�!&�*VĬ�X�1eCNS�n�|<t0x�^=c�������҆۾�g�T�ڃ�i�(���9�6>�vQ��[���86z�x�J#���_`ாM4V���'��<"X��Ƌ7�hR�,�#�qUUA��᠌1M?~�獛�Odَs��M��J��icU�ݖY�
����p����:�	��tj�CA�>���у�Z�v�78��ޟ&�g-�O���Uh�|���d��qC�#�y)�����'�1�[�4���~:"xD�0�<h��a�@�
І4�Z��c(�F|iPݥ�Z�:��K-�2�M�55��Ȋ��N&1�&~�u�+����Ba�&mG8=�� �K*�b�����N4j �";�*��r� ȘĔ$�&JKj�F\��i�S٩/��Զb~<7ـ���s�|¡^
p�Ph=E�.8FD�C�aaa���65�&�B�c�m�܍)����J%?S���CN�;~$��{<*)�xg%�%B,3v�m-�v1cQ��LC����u�ѳg�\�,��GǍ8zp᳇�N�n�E�j���a_tw��gXߨ$���i�|w�۶�lDW��v�<����+�&�G�Z��vφσPܪ#P�Ue�'\��g�6}Z>�C�C�`�)���C���3(v<��!#<�g×��<�U��a^�����'�6{��x���Bh��?	��8zY�M���}���]���Бҭ��g�n�{����:��oN�J�O��t���Cn����8 N²�A�DD)]�Ve�9�Z~�I!�i+�U�VW���.�<0v�i�Q*�YYvt�|z2%n��h�a���i��^��8Y�U[;>���0������F�M!g���۶mv��޸����Ӈ�>:p��g{!ꢙ�UU�
v�~�t�2>�O�c�a!2�8j��3��o�.�x���R���BL*�����d|5!$'�?.���$&������� d4�C�ի�\(<am�l1���8�Z�(�tg�S��]�1ſ���Ww~�t(�tx6BC�=؜(�e~0؈��,O�a�!�
(���AA(M6'��<&�Ǆ�%�"X�%��,DD��x��B&�6"""'� �"P�����tM�g�f�D�"<���B�DM�"tD�,N��6&�	��&���f�!ҒQ@���B"t�<%�<hM�Q��C�a�|痧-�m��1)LcL鶗LAR�#-C�B�m4Ҽۈ�!�tB�!�ʊh��cd�244A@f�e��
SP].�!�!F�)����eE,E�Q�Eu�M1�&������M�D�YM �����+�*ʙf^L��(�GiE��h�݈IG�����P�ϻ���_*lKF�eC��D�zU��'�W��en!1�z�Y�Et��u�#JBQ��U|�WI��db+�1LE�$v�Ԅaaȁ
���<���f����Q|t=�<��f�#(���x)��Փ���Y�d��%P��d#"/І��(�
k$"V
bS�n�Rȡr���c��-�Eq:2<�Z$�G��+P�!B�EL�*��=�x�c�ו�r��um���w{��UƱ$�\����?"��9��۷�<9}ɬ����P�O8����P��iQ;YQG�֫#R5ۻƦڇ��"��Ȑ�"��T��,�ؕ�I�R5bJ*��A��ɒ+<�G���v$�[1��b��+�j�E�:�-���L��i	���%������#�D��yn�Ɣ��jĖ1dDo�8Ԅ����G�v�x�����RS��&���3�3T�� ��d�C�����33<����9͹������Wo9�m������-*�y�snfffffyiUy�
<h�Ə<a�L�/_8��=-q����+����)"�B*?�M7�Yt��	)(���֑�,�DT�B	��Wn��M%��Ad������R�1�dVV'*r�E���풱���:Ĩ��x��#j����=�^ؖB��r�\.��c&�y=����ɳ�u����O\�c��<Ķ�Cnfp�B��YO�!>�r�x��$$�����d<�*ĉ>�����s��6;'�	��\�I
Y$>r��CO�z�4?u�4���Wi�3�VWk�	�ϋ6a�?0O�"`�(����j�����T�@�X�=|��x8|d��Y�];r3��X���F;g��v�2"�ݢm΃c��׍�FG����0�{;U�)�����7��7'�`��q,RM���16P����-�L6�&[r-���G��F�4h�F?	�O�xD�����W���쩭I$�49�q)�=-�|���'�������N_�4Y�u4�`�n-mY�0�ϥ����GNǏ8���Tj�B��#T4�V�dT�"V�"j�Զ�C%�C���>Ӄfʪ�C�aO=�C��]��L!'���0BD8�x�5A��n�*`�%��)6��f��h�4~4x��:"xD�:p��qڽ�9ɭI$�8��:!�\�c�ۀ�a�2Bu���!��&C�eA���X���4���SU�X�!���!����������ܚ?[Uj��Y�a�f�?;b{�n�I�J8���8i��JL�ͯӥSP*S���t5�$�v8�[dĐ�Z�!�@��<h���	��M�=!��(�=���Y��`B�!�2�W,��������(�q��),d'ɋu�Ld�i�PŨc�)-���*SGU����� Y��554LګD��bu�W�CJu��rX���&<�dv&�i$�oM#8�7IuE���HBht�C��Ç�!nB�x���!���쪄�Q]�4�������V�����z�M��xvx��Td��=p��a�C�r��x~�I��
%&&�$<:�'F<Jv�6~N9*�Ǯ�|�fΖY���b%�x����kP���$�	�����)	�*U��۵��x�l�EW��p��ِ���Hv���f㐋p�¸��~��({���Bxs�,1Dd<<�C��Yr8�Pl�L�⩪(�,�1����wSC�G�r�\���z�wx�)��3��g�����J2�8QG<Y�g�<"X�f!f�}&ꉹ$�@���a
m��!!8t���G����U�jHJ�S��o�+�JC+��7�p&���e��f@t�5n��R-t��f�|�w�佸v:���~(���
��{��j�����E�ǂB�������i�Q��$J�E#\�"u��G�4�7�d����`���	��l��&�����Lfá>���&�0؉���O�"Y���I�HLmRY2I$�==�B�Lɞ�;g�SNd��Ae�L��ڝu��'�c3�P���y��LUp��Ƹ�t�L�\�Tr�^�!	&���)���À��8,��wnN�!���ԥw�BI������������e�d�0�!E�t����4x鳧N:p�0[��|-��!
���
�"��u�!-�ٻD�+#�"Ȭ*!Yy��&�L��wM)����6o�D�q9e�"&=꣍6�Ӱm�d�\hđtqe���cS.����I$��8<c�%		��JD,���!%P����d|XW1��5U�1���<p>�����J|3�óa���#a�|}�?N�$����Z��	ƨ�h#�}��S��=S
�b��jZ���R�<T��K"MD�V@r������|��x�N�ބ��4�6hᣦΞ0���K0�j��H��!&s�˰��a{*�!���u�����巉�K�Y�$��(k�&��gH�*Q4����[$�q�+G�6QD���ʳ�{�:�ʈX��>�s������gu�nUwW�6���z��Chh6<v:ӭ�zt3��}9
�+)�vrn|h����G~1�=;(�����K�æ6`````` �M	�L��4pD�x��O	�,Kı,Kı�	�(�b""X� �hJ4"'�"'���b'Ԛ �$8""X�(A�H�ܜı:t��f��JBQ���H �>Ђ��D��"xN(MP���0�	�[=����=����o�_{�w��k/'8�����Œ|�C�*C��7_h��M��Ҍ/�IWU�~N>���ԓ���=��ꉮ���[�9�����Uy�s�\����̶*�9�s��������U�9�qs33332ت��:Q�GM6tD���K0�<t��֤�H	�n�;.���+���GC�����c�AӬ3�BI$����nB=�Y^ƍ�x��L���X��Bܭ���q�-*�X4~WO:�=ǡ�(%U�t�k�l><�o��̘��!�ٓ�O�?��W˭���A���{���M4a�?��'�K,�d8`ԏ�D1�$�Gxm��Ox���r�+���⮐�K0A_H�6H�m���eI��V;Q�jeB�BàӜ������F�)��QD	P�<�Y�}��s8������Ϛ�RBFI��<�O�ۧ��H�t-�x�>	���]�J�v�0٢�	��t�<"X�z��^�]�#M9V+�D���GmU�U""��J"��rH�!��H�h-F��KT��Cs��k R�f(-s0�$��m������`5�PJ+�
�2¥"%
��4#�I$���pYr�[	�� �&$�Idv�-��IS&g��=��=3��7'�4<<vb���E�:��d���{Ǻ��n�N��$�o�l8;��)��A�ߝ�-�!T�U7ק\�9�8������$�2<���1'��E"�v"�!��+c%ߡ��0�jh��$Z���,���4Y��'DO�"Y�+���I$���/��̎�E��4<�p�S��>z��$�a#'���x����x$ѽ�ZB�둻��BI`d#���X�b�U�ǄM	d\޻�԰�%�?�2C0�o,-�`>_��N���4)�dy4+d	,���^��]�Q�m�25��T򵽕Ҿ����N��=~�m۰����|�;�O��ߎ��m�M����]�	��K0���rI�kEI$�$�I�����%�ŘgCF�.6p��$�*�i�������:v�|�{������Rc�"�cTe'Z�U'��Y���;�YMv�b{G��.*+u
�]�����5`\������Ú��}�1�zO��a��v|=|->,�E�0t�����b%���7�U�P/.I$�v�7��X����z{�R��6���Cz�������+�I�r�L�I���R��%�<xi�B��f��}�p�4ēТXӗ�����[���GY�[
���sq���2�)�4|����T��T}����Qӆ�ц�:~�%���~OO�>8��Ld�HQd�O�4���B9p� �ewX�GD6��c�>UB��~Lh�hI�B ��G�0�~çx6��DG����$!(D��R�,�ER��Q�F7F���$�7�3`��A!q!P��*�2��dg���L�SD���y�+��C��v��CA�Za����G,�{$6l��q�P�-�1ƃ'�6�8,�24te����H��M�F�B�
�����ǣf�Ͱx�:៦�8a�Ə<X�?�<"X��Y�Nr�]LVd�Ip8!��)ɭ�6�e�t?��FI#$$BY�˜KN@�������m��E5Thy� �����]9��l�[�nB9��H�X��<LY�����_}MRUd���)��=�	3צ��vD�����d�������<"X�Η�����(����I$��[����!A����0C~ QWfx������n�8����Q�?�b��Ȣ݊\�Rb�$��Ĩ�e�$,��ǆ���ᲊ�v<lp�$>��!!�\���l韞��#�a�#�٧n9X�eYl�t�,�nYﯳ��4p�f�0��#r%��08t�$�5x�ԒI�X?���8��O�C\�����Y���b)�5��ܭCB�45Q
�TuöI:x2m�]o�>��=�$!<3ɓ�rt8�wN|BITptC$$�KCA�>w�$��$�O�|(|d��y�L�\W���I���Ύ�^�4=nW���m����4YG��HU�C���G�T��1?�������0%�4ѺQ@�s@K����������o ���j���Z�,�*R�2��d�Y2�Yd�i,�S--)�)e2ee��d�2ee�ɔ�e2��e2�L�VY2e,�S-,�L��)��L�K)�)������ɔ�d�YY�)e2e,�Y��dɓ&Ve,�S%��̖S&Rɕ�,�L��)��S/<ܖSd�efS%�ɔ�e�Rɓ)d�e��ɔ�d�Y^:�YL�L�RʦYJe����JY�e)��ٔ��JRZe,���̬��,���ҐʘQU(��Y5C
YfY�e�e)Il�iK,�Ief���e+%�L�J�L�S%+%�S*����2��ie���ie��ۙe���*�R��)e�,�4��̥,Җ[2�SI+,�*R�)V,�L����YK2�-���fYKQfR�̥,�)Y�R�Ye�JZSK,�iK,��-�Ye�T�%�l�)d�e2�-t��L�*��,�e����-�e��U2�T���Yf��Y,�Tʔ�[2̩Kd�&W�eK"���R��R��RaEJ*(����T���
,)��J,(�������*QIE�c�ژ�X�թ)�M�0T�T�Ȣ�)(�����T��0QJ(��)E(�QJ,S�����R��*QdQE�X`���Ģ�XQIE���XQaLRd�Ģ
,(�EE%QL�IEETQQE(�QIETX�I�QIE(�(��Ģ���,�TS�J)EIE%QEY%%IU)��KJZRԥ����+)��������RR����4�ȗY9I���Jk)��R�%(R�R�R����E(����JE,��
S)���MJ����iJ�[J[)YYe5���)B������)*�R�J%,E(��JP�$�B��R�R�K!J�J�,�R�J%%��B�H���"�JQ)d��J�K,�V�mJm��RҚҖҕ��Җ��)l��+)��e5��VjR��YMe*��Sl�ԥ�D[̫��ڔ��e-Jm)������Vm)iMR�R�J�k)����ҳl����ZRԦ���Z��Sl�ԥ�-)�����-)e,�VjSR��[)l���Rȧ��
�K�E,��E,JP��K$�
TS5Jm�*��)��$�E(RQ)d)a)I)Q)d)D�B�"�"��R�J�J�K!K!J�(��%*E%�JQ)R)dJQ)D�I)K)m��Y���)VR���R�)����me*��e6����)�)�R��,)b)(R�R������,JR)RR�H���)jRԦ�L�*�P��IB�������Rĥ�J�EiK)�R���-���Қ�VVm)e2�jR��R���ee,��K)YJ�jR��Sl�ԥ�ԥ�,���)e-����,�e+)P�J�RR�*)�XJU)iM��KJYMJl��e�����jSYL��YKJ͔�*R��J�R�)�J�����������5������)�R��6��"������E))RR�ԥJR���SR��ZRҖR����%%E,)QJ)QJ���)QK
JR�R��VR�YJR�,��K
����R��(�,eH�d`Ĥ��PT�����QJJ�T�bԲ�*YT��TʖT��VYZ+d�*���Y(��)CZ�SxI�C))��S*e,��2�U2��R�eL�R�S)���S)J�TʖTҚU,�RS*YL��JT�iRʙS+2�eL���eS*YS*eK*�S)J�SeK5���S*YS)�,�eL�JeL�YL��,�Tʥ�2�T�L�U,�L�)��e�e2R�ɔ�d��Y��2�e��L���e���d��M��-]��?�)���H~�M=hZSAHv��^�Uj�ͭZ�kjڢ@3��������	����������C���)��O������~����~�?t����� �����5�����03���JtG_���%����rd��L?���W���h��g)�_�5�N����'����������QU��O�����?���_��r��A��D��QW���w�(���ُ��C�?h���C@�Z�)w�0��Q��� �������r���XJ���QT����(��?i�� �D��̀X�Fi������3�����p��lܝ����%%'����E�F�f�èi�?�N���O+��O{����yΑ ���?�����_����T@�cu�HA�DڠL�"0LfI"�X#%��T��B�*��0vӯ��@lp�E������6d�����ni��  ��s�s��t>�!P!I�T��J�AaK(�&RL�RBI��

�������Zl?�| "?��-xM�����?���H���� "<j����'��P����O���O�P�� Dg�������N:��(���~�gC��_�4o�Jq��o�@ �w����``��=@?y����L�����	�*`���>H}�������!���~��?���TU����#:���V�+�a�ӧ]�����J��4*��e�ʊ�?���)�a��,S��2����X�?�������?�����V
Y���P" �r�~�	>� �$���,�KH 
�J����l ��0�ar1,�2?�?��&�"B=SHs?����`��N)�㒄����	�#�UPG@��=RC�?����'��q**�� ��d_��X�&���AO�N-C����?��?_��~��x���K� )����.�~�����	����t����䈵��Ҍ�X�����x�����EP��p��W��A��̿b��F(�Q�1DcF(����#F(���1Db���#"4F(�Q�4Db���#F(�Q�1F#F(�Q�1Db���#F��FѢ1�1DhŌQ1��TQ�F(��4Q�����b�ƍh����(�Dh��F�F(�Db1F#�ъ(��(�c1DTEDmQ�E���F(�E������QEQ�F�4h�F4Th�4h��(�F�X��Fƍ6(Ѣ�c�1�cƊ(��Q��1�Dj6#QQ�lh�Q�EEETQb��"�1�QF���(�j(�E(��b�(�1EcQ�Q�(�F,QEQF(��(���EQF�X��F�(��EE�6�Tb���*5���lQ�(���61�F1�4b�14Q�lcb��lcc"��QF�1b�h�ŌEE�cQ�,h����,b(�Q��F#F��F"�E�1b1b(�"�E�1b1b"�E�Db4Q����Db#�(Ɗ1b1F"�E��E�1b�1b(�b(�Q��"1��cDDQ���E��Db�E�1�b(�Q��Q�1��(��b(�(�X�1��E�(ш��EF,c�b(�cE��F�b4b1�1#F�b1�#�4h�F##��F���h�F�Ѣ1#EDb4F�������5�QQ��4Dh���6�b1��F�#b4Z4h�����lEDh�F�X�1����#DF"4F�Dh�(��4Db#DF�Ѣ#"4Dh��F��"1�F�Dh��F��Dh���#DF���"4Dh���#DF"4Dh�"4Dh���#DF��"4Dh�"4Dh���#DF��"4Dh��Q�#DF��"4Dh���1�Ѣ1#Db�h�EF�TE�4E�4Q�������Ѣ4TF�4F�lF�4F(ъ1F��#Q�4F-�-�4Qb��F���lh�14F�h�F��,h�Dh�F�E#bѱc�hѢ4h�b�#F�#EF��4X�F��4hѱ�F�h�F�hѱ�61��E�hѣ��h�1��bƈ�11�X�cF�hƋ1��cc�b�h�4cEhƌh�b�ѣDE(�F4cF,F4b4cE�4hƋ4h�E4h�DcFƍQ�h�Q�cb1�(��Q���ŌQ�1"1Dh��X�#�(�E�#b��Dh�Q�#�Q�1DF#F(�QDb1DF#DF",Q���#F(�mo��k�oo�������?�"'_�������ǳ���������������ƣ�����6�b��������W�����H7��A?y�����S�H���	O�2��2���L�*���~j�J���)�E�Q�����Rڸ���Ӡ�O���������4��2%i����8;E�����G��B�	��1���q,�ô
Q����? �N��	���&���?�R�����@�����?����?��$�?�()#����w����)�#-��