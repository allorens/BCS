BZh91AY&SY"���ֆ_�`q���b� ����bB^�    ��O��I��T@�J�a�MTڲ hʀ�*���Zj�JѣmL��PI���1�PP	i��!T+M+l��:�`Y���Dֵ[a�m����۱�lZ�ֶjֵj�`�5`�v�fʭki+(I&�Z]�P:�LU�jڦ�TiI+2�i���|κڵj�f�a����Y�i6٦��[i5X��d�+3 ����Y�"d��ƩVV�mE���ml��h)kV�+d�V5�������lw%�F�5���  ����j�v���@(j b�ӶY��:ý�*����պ�z:$=U�����W�4�z�k��o]��/m;��6lme���KmJ�Q�  |�A��S�]ҩ(
���ޔJ��뷛y묥%v��U�m�����^�.*R�N���=K�][.���T��ҥ���=*�vԪ�uyR�^��k-��-�lԚ��1��SW�  }�{����i�^t�t��B{�K���ꄥ^�[���t��wTn�%R�]ޞtz���F�u���7��J�*kk�w'��$
{���*�i
{�L���ֶ�L�f��  w��J�>z���]�uI[�gx*��vԷ{x�ڽ����u)B�+��;�Jtҥ=޵窏Ym�[m��{�Ul�\��z�����s޷zT���y{��mM-i����d���i{�  zn�}5JSMg����iJ��l}��^�Y^:��ҥJ�.�תR�������z��*/��8�*�J�N��
�*�/n\lԧ�.t�R�)����6��-[2UmU�Z��  {ꄾ�;m����v��Twz׽JUYM�Q�N���S�W��[o{�w�T��X��f��)�IS{̮�!{���3��J�mp;zHT�w��͕l�fL�fV��	4m   ����v2��p;�B��c�]ޔR���[�[j�J�����T���׍J�(oG�yu�$�U�^���L��s׏=*���K���'��ͪ�Z�Z�hֲV��  O�R���ZS+�����렷�x���%{�\@=]��7oO{�8=��F����
/`s��@ =�����2I�f�UL�R;�  �|���Y���{�����t�1���j+�W�q�t���^���U�y���7{��%U��-�T�ȫVЭk5�0��  �{����������^���ztw�8�����ZW���@Z�� h[�{ލHy�N��Z��O=QA/�     �*R��	�2b`�M4�S�4�)ITd�F2 i��i�B)�15)*���     ?�hIU5@h �   ���&
�*3 ɀ  &	�T�ީ	�=����Fh44�1??��q�?�����
�5�砮�)/c�˜��2�4�ñ��_>�>��~�W߾=��@W�A@EO�@U��_�8���������@X?�UU���*�>T�2��+��������_����=J{2��́�_��C�2�2�0��H2�0�2��__�W��_i__��@�d�W�W�OP>0�2���!�+�+��2�2C�� ����<d� ��<d|a|d|e|a|`_��̯�/���+�+�x����0} |dC��D�H�hP�J(y ��*��"@�y ��	��� �J��)䀧��B�y*!䊇��J(}%<��� By !� '�"H(y"��
���0J@���@ y	���
H�y �䨇�
@��(ЪB"y ��� �B�y #�Ĉy()��>�|��S�O!@�(�� ���@ � )�(���?�>B�(�@�y )� ����H
y��"'�
�B��C�Q_%@zES�TO <�<��'������'�'��ġ��W��C�C�����>��"R'�!�(|�0�̡��	��O$O%�<�<�<�<�<�=������S��!����ɯ�+&���sC��ؙ�R0|��Yb�<9T��!8�{Y�4l�Fú����~�|�E������/ͽPLw%��64�T��O(=*�^2us`g	���w����v�og4�n�����olD�{�a��c7H�RK)b�E��(L˭�;��8�e�^�R��ą�
��U�)�ϱ��e�VܴF�*E�E-��Z����3�WV����ؤQ�n�D�N�Ȟ�դd{�����JOs�A����n4�Ai�vT]��^�qN'M6Ί�$c�tW��m@�71EC3R dKn颔j
?^}B���`V�Ti��s�@�^��D��B5j�1�M"�v�1�:+|�\�O"��[��dAֶ�B:P��tkq��4�VГjk#�n���6b��ə�At���L,c��2}f��M���Ev��O��y��!��j�x-�sC����û����Z��k5���ؠ����#N�{�ʪI'M����7n��&�a�M�{A���2F�7wFt��j+g'�g�f��Z�z�P)V�0K��ˈ���]O~��o!v�i�q&ǝ�f��9;�6
.�b?��s��'ux#��r�W���怛���}��Kt�ʁv���s��Z�������}��w��d&�!{��ˡy��:��j�ֶZ��KS�+����Vm��ǓY퓵5@��W2�����T
k����|y�v�nuۚӝ&�/x�=l{�#]��	�,�NR�[��Тn�*>�����=�+_-
j�5�Vل�1d���7w5�b��ɍ���u�{u�'pߌ�Y��[G7 ��q�oN�>�w6ȅ����li�?s�\}#�U������x�ٛ�;D:���]�ݑ�����e���xfB�R��ШRۉL����~sxW2�q���{����<]�@|����ub�]��h�"�DNpL繨��b��*�چ��Iv����a�nM��D6uu�2L�n^ɜ^�q�"�^�!wo!�K*ƙǯ�8]�b�[O^I�w��sU���k��i��Nd�%��$EB,9�c�=D�l�Q�ѿ�m��"�\B�O7$�jH\ȩ[v��!:�+9@n�T���;��z�+m�h�wH�%�Xޑì�_h �9�M�"�z��<: Q�(�����u޲�ZX������u���q��Sn'3F�`�ؐa�)�-0@oo{����HR�x^�Z��9�����VWV;��n\t�*�
���m&s-�,rTF�d�;$�b�7f�֑�u��p�2dJ-{��a�7/
iT�{�QY�VP���2-�-��۹T
q���q�>�Mc��A��Ⴌ,����e���of�5c�����%BQ��GHajc�#��,����k��h[Zis��WW�A�s�ӝ��H����tr#3��ĽG4��4|��T��*s��(�c�xbC+ٳ��WG*X��#�\Xˡ-����T�Ω�����>1���$	�������-��KH!�׸�&����v"�rv&����V%��2����N:qP�af#�bIeS
�ˤ�E��˦�j�2���If����sO|h��(Kr�Չ+Cj�j��� Ul�M����<�F��Ȱe���V	��Bgv���V޻-j�Hĩ�vv�����©0Vb��V�M@���*�Ɯ�:���ϭXR���TP�;9S�!������B�9S;	Gby�k�����\���uc�T��/��v��\�8f>�:j�(�c�Ol�ǣ��Ŭa�^^͸�G5��n
�RĮ��A=YX�2���Y!0��Qgw	�Qܑ@��{M��n��Es�X��&ȥrlcw@c_Ϊ����)�JC:�f��/Ȁ_4Wi�U�\��1{�h��,��'J �	�ã��.�ו�O�Vy�q=�f�Me��:4�qh���wr]l�PKG�^�.eN�Ĺpkq�#���,�N]��n���Ⴎ�F7�J��D����v� r��	�=T���ӫ�qؚ��,#��6�����9v@��m�
�4�9�ܼ�r<�4l��2:��hZ6<z�1�
i}C����>�V�``�	����	}/R�"2��S�p3��f��[�U���(fBE^搝�o+�!a	���&������'ۗ<xN�(��{���l��y&��&�9�z�f��v�M��4D��ǩqN+V�e���n�6�9�k�0կY��S�K������R��ZTt�6::Ε`Y��`#����3w1�Os�c�"����(�SA��;��$GFl�i;�$z�S���oν�����	�xR��u��9��������v�v���&��;K�ֲ�dZz���b�T�]0�(����P������՘C[�����F7N)��m{�0�z4~r�ڄ�h���GS!H�
M��yC�k1�tTL�w�ia��<��.�F��zLcv��ܝЛ�j��^Q��V�l ���?�'�/5Uü�xӥճ�C��.�
�5�Sދ\',�ծ%3]miF��k^9�����2��/g-.�9NX���qV^�,�{J�j�1�SV�x���Rb�~h���)ef�ջ��Z&B�n� *��L�d`�q�X&���bnf,ݬxSR4�{uka�J'��D����{V�&"	c��_=Z�G/^S[�D<Y�Vrz�`ȑ��@5��������i��M���(Kү-�Չ�OwV�4�]o���iR�i+�wHV&m^�,�qnf��p���ר��$m�`"#��w�ږ���x,���	f�4�[�L����<am���I1�����X�ٯVP!M�Ã@75	d�$C4�KP��'K^R썞�rӔ��Q�h����F��E*VS�o�ͫ3eu�k��饍�)��awq(�7:�r� Usq���͍#Y��nMY�!u;K]�%��.lQ�ƍK����X����d���=�D�4BU"6��V�V�r%-<�Wk5�=� 4�	*ʩ�f+�7`!��-�Yv�0Î�F�v��Ul���Zw2���8v��ZV�R2���4ͬ��<,�h�q�Gɋ��X罈,����f�Z75��BF�]��D �UL�@�T#v�ͭ�0���UV���Q0�u��<������c�Dj�S+u4�b�0E��7�����4��=u(��-S��N�Uj�ɬ��������8"Ot��򔌤�d��$�_Z�6��*ΈK�F+�)�	fC�ze�n�2�T�QJ.��b�뮣j��gɏ�tc7x�7<[�l�Ǣ�9
�I<�X����mI��Q�I9�9�j�H��k�bv;�Z{�
���&U���4�E���v-,�*���6�� l�v>�c%��N؞wr5��N��I$s�ܫ�7
�G��f@�5T�ϩ:��0�j=���{����'Y,�+`7@����w%��qʞ��T���A�	�g�Rݵ")�.�	R��Ζ�+���1��4�sڞ�؀`�OKs���{5G�^sժ͍�y�e�Dp)�c�9Z��щD�O=Wk���F���}�qn�\k�=��m1S�po%��*�X��j��(�x.j/d�p���ٵbZE31_M�ٸ��{x���$$��p�A���t�5*LԦ�C4л�� � 42�Wp����x��ȯ��*�����e<z>괼��<3�;Ə����7��(�s[�d��:N!�u��SKh�Z2���d���ndj����s1���䂘��ܕ���1R��z��7�4�c��A
��/�]�*�b�.�;�ũ�o!�!�^�ÂmeE�5Ҙ���	a'Y3.n�wR��q���"��\+��k	��q}�C:ed.�q�9@�wtz�pG%ƍ��
j��(A�Z���7�E�������S�]`��K �j��`o��t�X�T��sX�.�ѹ0��"��٬#��8g�����]�h��4�/��m֥Y-������vE�Z�Z�|]�J��']���Fm�1�ktc�J'�Yd��1t6n©���VM��C�*R\��!�^8�Q��>�i�v�o0��"�Î��*�����4��ѥ�!_��uj�yV�kQx��4
�6�qat�;٭Z��uoL#f����`�za�5�%�q�%p�9�����o�!R���ZUǭx1��^�_`\��(Qy�h+I�v����OM���l|[�'w��L��O5;7AD����os,��Ae�C�f�Kҧ��v��W Vn�i�A0�4s������b�v1o�/N��n��*&pfH�#��I�:9
�*�FL�s{^X�� �;u/�E�^����+sv�yFs�|vw4� gWG��
�4Q�爱�����<X�t��d�E	��%R	��m9�ҽ�F��F���t�)���itt�g���
�v�+��Ƴ�L�U�Z�M#��Ojӡ��W2L[���x�9
�G(�R�$�U�c q���Z@�S��Z̆�;gQ)��y���v�]R�9ҷ��y�ħ!�}�^��:TZv�%l�Y��V�-�aY⨜WϹ]i�����M�ð��J�������#����&ɗu�ABJ�W�5ɰ3'L����TQ-�:�rp-�ɠ)��)4��7�L�3�2�3[���Y@7M��)n(0��k$��uԅ$n���#�a�\z�b�o^��>$0�"
Uu���X�f-���j��u�t.��0��D,K>���;��غ���&$�)�O����Z��x��j�G�q�&_�ǝs%��ZC�.�����}�a-���V��:���;7�sǨ��3v[�fg措Z�Xx��&�m^�4�+�$�f���4�;�ֺP�zKS$��v�#���]7���c�cq�gs�0}�pDSם��
��04㤃�9��K�t��f�	�y��2�x3^N��Of�xe�.טg�Z�d���v��rT�!��`'���q'�'�ba��93��v����t��&e�X�>�f��~2��1u���D`ln�#E����\Ȏ�̛7��Z����:�t_���f���Dq�"`���|�`;;6scH<w�\�y�����hhY�=+S�-�b�J	/
;���bR��n4��"*m����)v<��'7u}�t�oy��n?��ͧ4��-�F;�X��g"]UwZ%{	U�tǫ�etPu�� ��c�i�$�p6j���Dǯ�p�3����#�c������NObF�dgY�D����x�]�ϾHb�ZۨÎG�*����U����/���q0~0�Z�\��2ytL��57Ghq!�^X�r�5��z@kOd�V˅�2�Ջ:A�vh-���xWk괐��G�P�7�#WZu�gɫ	E~��~Y�^�`K,�B&hK�֬{gDܼ� r	��t�ҺD̼̚����&0�{N�pm��8�.��1"'fj(*�}�+tX�t$�u�/w[���lΧP�ʢ��1����qܱh�A�`L�2�M�܌	�H蹺�-�r��SN�Y��V�kݘ�I p�B�I�x�܎�˓��t�Et!��������vl�Ƹ#����W\��u��ه�N����"0XA�}�U�ᯏjy��]r�r槺�⛃�Q�ap��	q�Cق�Y��CՋwH�cU�	IpM���������Ǟ%.�M˸��3�u�][�1���E[zW��H���S�Gv��m�jU}�t��ќ�
�hʙ��L�F�]�r���`3	Ѹ�Ɛ�OY[��&��p$��V�jq=�Uc��8e�z��W&Y�S��0KwkZ�3ʙN��j��CI�L������ϡ�|x7B;���������35�ɹRx0o5�o 		p�֚�Y.��L+k0��^�[����Xn��fu�٣Yd�2H���+�6�3e�6�&����s7Q�c����.-x��gN[ٍ̓��껷6u�s���,���{n�!��aY�LAݏ�W�4��^ ��5p}�PU��rǛX=��˫�+v�]�Za!�PZ5�m�׈���͆ܵ�8��i����]<�C���'�[��n���>.e�w�Q�f��"��YT�ot-�6��?��;�ѧFol2w3$��t+��WbX�[F[g�� �P٠�/(�`+�Q�"��G#�Z���	�� �˚59�F-�H|�%�a4�y�Jn�#-�'* �nв�P̫Z�`Y�f�d�,y���־�Et��a�� x�'��$�n�X���UҦ�չ!ۣ�#�6�E�����Vޡc�S���s�@��Υ�dY%�䄃�X�t2�M��'���݃�KD;a� �ݢ� �wI���8G�����8�_/ ����m)F�c^RT߷L;)?V�7�H{<�;���Ow �Fc�fŢ�X5Ø�ݝV.�N�ŷ+$���S�6�ݚ/Tȴ�J� Y��@c��j��m[�WJ)�Zͥ��c�MAg/UXx��VޢG��a�f���dݽw����b�d��B��a�R�o�1<��,|�)��pֹ�^��yQ��r����򉩆�.�$�ys�µ�H��(U���lWwI�I��c��{����}�J��w1PC�ZR�r�f*�9��2�C&p�1v6�;R�R7a����Ф)�Z�� ��-WMyk7e�j�"�&�"�a�5�
�M��:z�EM���k1D��0�f�A�����9l�qq-1.�h�wq����|����%��}��~��v�7�3��m;y��Lg���.7�V���nɔ�[���hަ���V!yӉ��\{���8͢�;t��Sw����K�P>�z\���}d��V��ȱW����Gi�k��'+�P�}�/iË�OE:��57+&uZ�U�R�m�jﮉ�kx�Y���ֳ��i�|{J��~ݾg�o��4OR�hlTV��6u<I����1���4�/�s�m>�rNc�t`��KV��q�,����Vu̖�:�_w)����z.г�CW��et�:2���u�d]I%A�1��ˆ�W�Ó����{-����R�̹ܰ���9�A9uغN�4*#0m0ܽ�C vmWhz���ioM�e ���b�6�{��Z�9aK�Cۙ�Vx��.�6�Z엑�u(��`U��dW��wv4�#.�	�m�I�[���}��{�Y$�]R��΢�gRs���5k�}�ѫ��9��b���n�v^ڥ5]�V�H���={,i�}`��Y:H H7������}HD��w3�=0�H{����t��[;�6�jsÐ)�g�^��e!z�p�����b��u;ft90��j㖩�Ad`#����>�Y]��`zu�[��m�;6\��sV�I[�)8�c�u�+r�E��[&�Ji��V�Kt0���B�f���dhL�!��G��s�v����Ѥ�]X���Q��/�-�;͓�e_����Y�w�9,ce�J��)f��>���u��ՙWg����%�6S�=�b�;�a��x��l�E��*	��J˔j�V�s�t+N�yGE�{�!Q�o5����n��j#oN��˪�U
�4�O;�ؔ��or�p�C�_R������9.���sd��Om��:���o ~��p��7Eb��4��Yy-g�hK�,V���;J�j�/)��uJ#A��Z�L�!ޜW2�8�1Gκ��,�M%�jU�
�#J͖�J�>��U��o�ۍ�sD_eg<rO��m��7G�_���<4Rkt�Ji�P	��?[n]<n(h"�XkR��w�������ڝ�9����x�5YYĹ�ip9�}���0��{��׏�"�p�͒.&�ؕM�WKn��9���gP-*4�^q��C�n�5ph��xr}�`�ms+y��郪��C�A��c���&:���gq�X�� |h�.]6PZm:ǻaQ�ޑQ̨nb
�w���e�@ܖ��A��+n��/���Tx+'��R�G��ަʛ��#ݺ�9�g7_/�/Ӑ,��9pY�p�9�bF�~�<�m�xUt�.hM_����VS�Ef�v#�{��[2Е�����v��l�i�pn퇝rј�S�ҋ�>K(�H�r�pZ����������_�X�Da�Y��aC�F����.D�:2v���m�a��X@��F��m�)"�az/Xiu#ZyG���n����63�)�{�7���
M�Qpo�Y�ï{F�ϴ]�VY{WNg;�)tPn�����9�@^'�a=�,ޞ��dt���e��b���1\�ʏ铖C���ۙ˳����Js'$�v�c�/ΥH;��wdv�mf+k�b��.�*�%�U�C���b�ʫs^�"�nc�e�2U����E��`�� ��\����3�'���D��i��4~�ge	���*ss��Fit��*>��d%;rz-�	�]v�����v]���+߮?5z��[�X�6߫��l(�B�emZ�=7���N�j��|��خ��$��[(��Zۢiؚ#��c��&t����������ݶ�z�oKQ�я�V��Ѷ2���q���0�:c�E,��N�ޔ�� Z�orIR��-;N,vf��LG�d����9.�j�}�Tm����.xB�Fy���;����/{</�a�\O(w0o��_/�*�`,!�,b�������i�G6��r���!�\M���7ѻ�YHZ�Z֎�kOkb|���o�zu���Q};E��u���e�B�L���P�ik�Jy��W@��M�oL��\x���<����`��`�_�_(��|��Nr��G��:�|Qw���dI�����y+ܙy��t���O��U+A�nB�j��Ɓ�\��������3�JݦD�D1(ͺS)P�{��n�JL�Ï)8(�W�0Y�e_h�㩶J���/Q<>�읝��ux��̪ʳ`�h,Jm=g�g+��> <޽4�1o�;Vwy��6�e��.�:#2d��MԱ�by�(�Zc��*��Nrك����͝q�ފk�#.Jy��\h�Ve�x���|���q�y邱��4��/Mu������U�y��(�+I�l��Cj�7%5�k7�Sy4��OV�y�KE�u�[��,�!v3�<X	�X�'�����3X\��C��3ϳ��L~��R�3C�3O��mҭ�]u�R��h���淥7<��@�䦯��>����r4;S�pv�i}�i
�B�0���<7�{;�@�W�i��Dp��T932��T�V��
��*jt!������*{�|0%4e�o���!Z�,,��ݢ{�S牜��=������{i	�+7te�*ָ@󒑋��I�y�X;a�W�lG���vN�|t�H��W���@���S���ΣAr��j�5���E5v
��ioG�b�ii8�Xi5��:3M�X�@�o]��7%�x��5!;�M�7ؽ�/��$�mC��-�)eSo38SKM�Y��lΛN�2�ݲ�DP��v���xf9�A�D��j��pZ���+��c�%�ڣ.�=��g9覱f��[\('Y�sUo (����e�cX3�E���zfq��J9V��YL�k�ԥ��rܮy���[���c�|��}].�&�᭱X���<�X��Ez����K�i��aA7z'��PoI��f�<8zc(M)dY�,�Ҡ�Æj�$}[�� �+�	6V3z�wT��:u�׆��'Srd�t�y���xR��@�V�]�3c���A��';6��ո��i�K�2+���5c�zy��n��w��?du(]�^zY
7ېl�&+Ց}�������b���A+	kje_�-ŖI��4�v2�6[�5].�8T����[K$�`�p�|�WS�cޥ@C������t�Jۭ�:�TM ��@u��S��T����E4+0��C'Yn���{,�q�d��Ga�%�:��&s���@2��I��M٤�F��j�VQ�W&O���M�HF��)Ĩ W� �ok���a�i�熙�l�]�O��}���^��x�@%ﻆ]{�O1��C���Snh]̖VA���Y�{&�׀3��y��W�F��R]-��A�/�0deM�j+�h�Ҡ1^aNZ�X����2����6��8�*:ӭ
 �[4ھi�PD�����7�� .jc,ws9�u�]�2�1�1�0�@�����E�[�K5�:�4���&�q��l?��R�Z�i�f�2��5��3�`=Lo�|���<�1�}��'�yFr�1n3}=Y�r'F/	���w��+�9tLWsv0�1qYvW;��Nf+bpT�f�B2�E-�$��vC�b��\Ub4�+qQM�|�;q����O`�ˀ�u��pG�n�=�F��BY���{G8�4Mք��t*����g��J�.�
g"���,k�H<H3��ߟ~���i�4{���_s � �li̮Ջ&�a���0i�8	���;y����t��ʯ��5�+ ѫF[�I�{ۧS|N�S�V6�ۜ4�0A2���uu�b�W�idۘ��-�*��4���H����ZyNu�Ԟ�g�ý��S���bM�;W�J��Pq�}��vǐWh��@֌	Q�8k�&E�3ۧw5d��o.H���+���<e�����nv��"�]�7\��K�1��ظ
�-y�V�����ȕ�auB�!�9��c��R2���Q�sԀ���,���HhH+&�}F����w:НA*$}�%m'�p�]���2i�t��v(y!@�{�g`�U:�WTٟN�<��쎎Ꜯ-,cF�x�J��YY���jӽ��7�1k g�dx��޼Y��g/���A�a��ޚ�/&�R}l��ne�̲Vë�f�X۷FaN,6 �Vq�,�4�R|���y��F� NV��X��O+7���T{�_I�֧�5��wP0��W�t��[ۉ��x���%z��$bW���<Jb���(;J�F{���V^�0,�Ƀ��(|��L^�@���[��J�k`�8�]5�������,�`㽢��&�z��oo	L��X�g��;T2X�:��<�.���9�)��"�8�����z�!��]���t�f��Q��(d9�5�B�R6�����m)�a�{�j����u�2ܫo�������`������O|��<בSՓ�{y�{'�^=���;{���*�]ʡ]N��f���6ڜ�R��r���ns�>�0��w_5�t�v�e���dQ�}��L���#yI�9�^�3��7E�p]�Ȯ��r���n���N���JGޞ���6�f�i�2�(:�)d�h�e�Q*��N�^3T����7aޅ�6��Q�K��&�].�m־Ո���ľA񩱌���Ш."��
س�,:���!�[ɪ��	�K㤳�ͣ,�N1w.�^ɜ�]�t�)KJU; �Xg3R7A@�4�J�\ :�'(X�Y�V�@���,�J�6	]��SO�ݮL���p���S�5iS����Nf1�ZT$kr�v�������б�b�&��8u��>��Y"�.i�"p�굕�ś�!q5�/Tf6j1�wR�WP������]�,Ԡ����fb�N��6[0fv��54�����L�|��}NOk�����-Z�{/^��+�]sT����dֺ
��v�?�w_gPO,���F�C�(I�l�N�|Z���+aM�Qd~�����=y���	����f�����P4wU��5p1�;��]
����K@�æ��^oض���]�.��d�Iႊ��u͜�cW[YW���vsZ��dǆA�5^�.�٥0b��܂����%����2�<�ڬ[q���c��M��!y�i\�'����io��'ʵ�2��@{*��ʀN'J�ʔ9�'�Ő�\��oZ�'�	�+jr]��Ҭ����،眓ߦy/e4�ݜ�9,ă>��g�K����/�$�xj^�9� �mq%���\ĺ�P�����O4n��)��/#(lo�L�a�Ɔ#�0n��䆷*��>�����_7b��L�����F8�z��Ǵ��Cפ^k�v�*�;t"0vJ;7���ͧα�w&A�a��H���),?�1T����gVV�CqRƶ�*My�<߲�}!k-��6�e[�
��d%��G%�Z0m�<f�\�@�Z9sR^�X��^��@��M>����
ew'*��B���vSiU,����]�W<����i�͒�;H�.\^u� \+l�^f��1�ǵvV.Ó���Wk��Y�	�J�U��d��{�����d:���N�g��B��+Ē�o-B�<���yLaD�/.ma�V^���WneEG�Ht��]>���$r��6��A�E�7�J��-���y`�kz�T�Xe	9GƸK
�	R|�3�㹅��P�Lޘ�e�����1j�+�-��b��7t��Ntx�j�t�e����)N��]�uٶ��Cf�9>ߥ
���W5GS�=���=��H�K�_���ձ�4�6y�ٌ��k���v�=��{Ãya���:m������}RS!	Z;�,ջ�V˷|bS�W,��,&�TC\��n�*Ԧ��Y�mgJ�3���ޮ��\�1YM���0]�`�j
Id�kB��t��;[���N�HdV��5i[V�Ѻ��!+�� ��R6m�镄�1>�R
^a:��m]Ǔ��O{)] ��{|E7Q�r�h)�Hb^��Hn���y�
�Tk |�p�#w��D�bBd֑�݇tPF��� yH$2���"��+�����z�Z�'�w.Z���9�i9c]\Wơ��n��VΔ�.���4�һ0d⋫�$���s������}:������	E}�\�{n5�R�U�g��~��׎�vf�4��R�浌��y��b=0�}ۅa���ۀ�0��]%��a�#��Q��jx+5��w��XIpB��F�\#�;�{=۶ר�d�!"#�n,w�k"�E�i+\UM���1EA��	�$��ĭ��p��9d�}���#�;��OXK	��|ǻ����7-��WLzCɝ���z1��q�+d4g1�e�Nv�j�DX��W"� �fX�B��mīqhΔ�+�xt�3a2���en�"*�4�ocE�J����Z���+MM��S�eK�ވ��d��Fd��J�VF�=�F!�p-�����T�=E�0>��2n�����jv�F������PSTɪ�9�B��B���r����b ��C=��خ9"���LsV�+�ZF(���˦�LAs����U�ݜl�:�����6n�٦WHݩ��9�E���z�=*b9���/b�1��=��0����#���Ӭ �I�E߱�*Ɵ��4z�úvBw;�Y�RL��v����|�������^�Rjg{�ӳ���[��S�u��p,ݶVS����2b�!u��.�K7x�d��9(i0;��{(���c�D��Ww��K��`�O�'��\�ɪ>c:3ԍ����ZJ�=9MEūj�-���Ezhy�z|��r�=�޾�{�i� f���`|�n'�E���i
V-4�.�i#vU"�F�T���7AQ� �E�.�w���o⪠����?���� ??d}���}�?����
�g�������wn�n�s��{>�w�����6J���:�mo�ɯ4��!Wn�,�Z�����9"������l*h�N`W���-�]I���S[x��y�IéVxD{�N-3��Cxj��]��|SF�ٌûb�OIo�T+Vk+^z�/tmQ�[ļ�/Q7�g*���q�Rʁ�m�)��1�'���i x��[��j׽����ಫI��C흯�M�P��h�Ւ՜iu��������P9|#��W��>��,hk��<�w��^fbө�w	*5��ЩV�e!�u'��:(�pwZ�8�G�����\�v��ͨ�nJ��{�,�ƒ�"�>���d���q�o}Lc=�	V�um��/	j�,ʺ����%��$���0zvF%O(K^ ����N�D\�ڦ�:�Ӈ��,I��ӄ0{�����&#m9Ha�uۦ��1k4�}8C��X��nջ��`�\��ľzƁ�hQ���᳢Jm]�X��.��mފL�d%�θ��蕕�qLӒ��"ۺ|m��	@<��N�_@`ԃ|�r{�.6v;��)�-c�O�ӂ{zh�f^YD�����r�7ƥr��:�VVMC'u�(��ask-\��oA��ј��<�q����Mǥb��6�~�ۛ��T���9%ۻ�;�9�
Nc�.�&�<��\�F�{W)�=\U��)'�Ƨ�݋��dWޙA�Y��)��7n�<��o �:w����y�[�=�`���S}���4:�N�p�,�9:�D�qo��7I(��I�/�^28:,mγR�J�#��F��,�)��Q���TK������Ğ��./�����*��8����W�,	f�{��x��i�K��C3���C5t׃���U���p�p���a?jW�h�IY闳�rS��9x��N�U�͔�tN��	���<�����7���8.��#'.<�L|�)e�]6�X��r4����0Q��Y�(�^m��}4�|�Q�ʍ��Wi�s��n���)r#Q����1ʋ6����ͭ5�s�4]�h�m��c���,n5v�z�u�'�R̴CZ�--Ii=��'�olǏ5�3��-��mh5���{����˲�+�o�N//%Z�:��^x%IֶݮkF�kz��b��_x�{|v�������B>�)��B:��;��s��V�AZ.�ǵ����f*�]Y�>&j��b��0�oR	�][bI��vPr��0N֫��ԡ�J�S9 ��X��j`S�3���}��ќ��� ���y�k6�Bd��-��לk������LeM��O+P6"��Q��M_e �Z/,b�5q�9�k�M��Ξ��-x�(*f�a.3�۪��R̨AG6� r��|y=�����hiW���;����rN�]�f-ᾄ�v 3�Q}��r��k��8��;C�X��РIu��$�I�F��Mc��v�~�P���'��E�{���T�,i��*�:û��QL�l�q���=��F�Y����)^}��$��'�p�BAu}�!���X�nVu2��a燚d�OP�ʖ�+,7S+���Ȩ&1�G���4�L�2�;��)�E�C��7s��x	W�o��<U!�8�^y�n1�̻Cx`!k��X�$$z벵��Za�'v��bf�䶻�+9�DJZ�sK���`q�e�:�Wz��̬ �=J�ͤҼ��^!��R�@
�� ��}\���s7��	�h�dmy �>��]��J!�:9����Y�,c�i��ٯ]�O�O8���:�ވ��2	��7v�xL�9غ]��&U��gT�9J�ͺ�Ȅ�34���>*�a4�*n���Vt�������Z��d�Ջ+-N���c{}e�N�v�U�lu7B\�y�(�ZD�P؇S��kWpu�5�ǉ���擰��'��zL��+oM=5�Ǖ ���ؿ�'���`�{���7�"[	�K����:�3�H����>�x�Ӛ=���!�=3:��F:;��ښL�ۙ�r�mq���]���������6�s�V�/�3��˜k��ټ5F�ݢ�A�v�>j������՝b��,��,��;LkP�DNj�������@�<�����
�39M�vŵםg��*��b��#�SՉ���r�YR��m��5)z��D�f�`��KYM�6AYΔr�����
��� �a�^Z��1g�~��O�9O7�z��W:�p�����̾[�9�ز�H��<�F��s�eD�_Patԥ����m=7�����[�
w	��v�a[/*��g06�]+ڜ�EE�=��m��G�ZsH�O�*���t�τ�i	&��1��*g��;SA8����4��x���Ge��ȃ�`x��:�rg+�x��Ɠ�};!�e@yl��rCM�"���ֈ�(Y�ː��(��79t�D)'ջ.���2s3��[�|2&��%�j>�����wYf�/hԕ
�{��#�\�y�+���X�g8z�Pܱ�� <��t�{t������C�{T^(I����.�ۜ��G�ޅ{7�.��0�xgS���i������<(}w��{=_-���'v����k���r����ⲩ�6�V-�$ɻ��c�,ȧgq%���uS�o`z���u�"]7���z$p((����B���bG ܷz�J-��i٥GPa�\Ne��d)3h�����y�"{w<��I$*�����tj"qQ��Qr���vG1�xt�B�o��s�j;λ���e��eqj���z��#�Q�,�� Y�=0�!���{�z]$���D��_[����=�>��c���@�No�d}�;$��p�h�g��{�a����3����C:��S�
=�|rr�N!b�^�>��?��^�}��W�zZ��N���̴�%���[���7f����rꤰɻ��xS�� Bn�C+zˢ�a���lt���g)=���X�ы�Nس���Dz��wթ�I]��e���r:���!d�9JFx��є���ͦ�4�-�^�31�J�P���-�W`glD�0��䛸z��Dђ����}�*'R�5@�M�e�t5riU���=8�U�1�3�h��e��my�+;,�B����`V��ے1]���T7;��{;�="�u��0�:n����8c�Q��w���X�G|NyQ.Z��X����n�+Ĭm;}\4�,8-l�Ժ�L�r���KR���%�t�O7	ֺ=��Ӥ��7�`�QJxg�>�w|��TvM5���F@wE�ͫ���[:sPP@����Z�P�X6!F��yV�+$���2g��O���r,r񙥘;�odb�(!-z:�|zr긖����f_�n��h�VΖ}�W3x����TX�R<��/��Z|F�5��Ü��rn��Lui���@��${�c<:�Y8D�}Y�-���YNdZN��띭$����eh{ucce����T0w�� 9�^�N~�����{o��^���XVK�b�@�m
��lf��tn�%[lU�B�i���A�dŨ��ն!�o{����&�kĲ�{��U��<=/��sd��{�x��h�`�zS��7�.�m1[y-%-�ѷ�aO+3(��c�t�%�+/l���!tO"k�M�	|0��%���&�]�J*�{q9&i���J�yeN �gY ;y��Y���$�ǫ`TF�t�9}�ۡvfSc_��/��*�1":�7#�
=�x
�5}�m��Mj� `	Tۛa�ij�i���!��q���Fh�6�U��k8���-�#����4i�I���J9��f
�wRԛn�҆�S��J$�������*q��/�\���G6Ψ�1G��\5P�b���b�P�GMD&k*��������"�YȻ�I���WV�[�O�m��8��Z 0���+L٨��I1X�z�h�5�Fmp�t�N�>v���{���
5�cy#i��Q��o-��>}�'�^���mg�<D빹��F���TB�z��j�q���k�LuZ;!�Q*��w�xл��5�+h�Wa�yv��+!�S�:����2m'�\)n�u5gj��d-��c6;B׍��Bzy�LKz��f�h䜜(�q͆�1��ŏ�ٶ0��y�w�q���w�y�bX�ݺ�$|��zb$@����w.�h�w�S��������֊��(�i���)�{ʕ��pڼ�x��t�¶��Cy���ug�Vb�46�4�V�n�M����W@{h'�Hߞc/z��������9���L1�r���]q�0,�g)"d<}�t�6�J�a16^�O�`1�'0�E���D�ܒ�>�״�Ńlc��̙���[}ڸ���7�M�f�@�KA�>I�M�d}�q�Ջ��La�Yð.�A��`8��+�T�+3�虵�I;���Ԣ�4%ms�on��{[�g+	���q�%��V����\u�Ȧy�n�K�2k������$�*����5gr�`��7LX�Q��!f���e�9!5=Շ���nr_"���RJ�n�YN���+�hڜkkN;e�M��s���r*8�,	r��ѐ�vF��w����\�V���۰GK��y��6��-��]�k�]X�u��*���u�d�����E}֪��<g0�o�����s���Kr����jfR��Ûom�6�?N���m��&�\�E�N5y�\�Y�G����
�����Y�PX�F}�>�t����n���!�g9L���+�Rѝ݌WW�\@8a�E-�e�m4�l�t�t�S�c��y����@��H����Cݪ��o�Q,WO.R������7wv!:��2�ml֨���ls�;z�I�B��hf�)�4n��|���`��N���q.ąj�L:>�j�2�[�F�]8B�9����4[96B1d�5$;kV-ֱ>�7��ly��2�^�e�M���s�]tx�٩o�:����u�mX��] bރ�m�z����ݔ�[��n]�\6�C*�:�Ӛb&B5q��e��LV��綶jy��1���.��=�4k���f�}��'4�h�J]L`�ZR�u;}��soH8�����|VT�~��X�ĦIc���7n=M����7�q�Sq��ne�srD��9j�+��{s��@�!d��8����t�_h��'b��o&G���3����*f�bx�/� ����������z�5C�`��qKHHYjvt �O<P�\��9UyYɹ�øaWc򚳤���b��Ec7�ق/j�y��&��ds��l
�+�é)���v���Z�§B�U�d�ͩ���Bb�F*��������փ�Z4V�[Y�0����&�i,OM�1^Z+����N����l�]��v*"�s�WY��np�tyHH9�zQ0Pز�'��!��;%�7��q���{]���Fqds�R�&?�#�M�1ρW�\�
to�����y������N��T�'�˅ݿ0�w�/P���Tw�7@V�����~�[���̞]����=�rD�{pn0|����<�73��u�C���!*JPL��s�ǧ+ND�\�������H�ȱ�E£ �u���g`��>y���	pnR�P1z"�<u��8�p�2<w�9� X=MU9��F����^��A}�X��w)m3Pu0���SV�&���0%s���f��5�����g	 ��U����i��ۺ��73���J����v���E%s�V-vs���ZP�V6�VE|e3*4�F��.����Emb�lnع�n+�G���>�^wa��{�$X\��5�����☛�'����t.��ky��u*�k���z�!�v���[�,�>��j��{�Td�y�s�F�#u.�h����O7����t�c�����r�E'ef]�48��u3hY����K�鸁�1����+c� ����΋Q�=̮n��Ϙg�x�	\�`�Z��U4</��骔��v2�e�n�<�s\��tR�J�7:�e�f�j�5��r�Z�s��K���Y|p�	C���Y�ZWe�0$3�����<��V:��@	|5��*��к�T97��(n-�����$$]��ɢ�Y��'��V<�YCd�ɰp�=�j"��5��ΩV�?t9|�������Z��8eZ1�}�g5h���ilcc��	���yT�&��a��s ����G ��JС��H>K��n8���]�v�9�e�9ő�7��d�L3�n����i&<f�&�Y������O`�7�E �Q�jf�	��ƕ�Zt�7�MB��2r㹁l��sp;Ib7z���L�T���X�wl�b�����+������G�����C�hQscz����yԷq>�N8�6�a���k�W�����L�gF���x�/RśL��`�)����X�l�|��+�<�+��I�4� �$�y��b-�8-�"��B�(��K�Y��Y��(j��V&T{�0����Ӗރ�2&#�����^ܾ{�<1{g'nݑ����ܳXeu1��N"_n}9"������3��pRS�V1J)�%�5�obYtz��Ъ�δC�Z��p�Y�Ǜ�ٶ�AK����U#Np�h0CX3d��_���,і�5�E	1h)tg�����Ϋ�n=;�׆/K�o�*��Ե�ۍ.j�$e�0$�_*��^�M>�%>)��.m�|��{�(=��%P��>�����@_�w������޿�~���w��O�ݶ�������W�O��m��h�
��@���V��`a��f��uk�a�q� �q�݀����8z-Zyߚzom�t�ҵ�ݜA�=�k�)l]X��NvQ���'d��RP�"t�yj�tK{�m�	�okq��]�	;�����W'(�P�<UK��<v�t�g��&-G*h>���UH�#6��6�%|�Z�E!�;�K���r3y��ʿ?nÞ�H V�cȤ#Ƭ����qMj*W&�V��nZ���������t�p)u�[�ئ���1�Asw:륲�X$�(ܕ&�Mf��ƣ���Qt�����.��7$;+89oK�G@�Eӊ���tj��[��S-\)4���9}����I��$,ٸUeI���Er�j��R�D���?0zh�f	�C�۾���9ճz��z	�R1��}��fH=X�12ga<����`��^�>��2�1�qeej�@��Ԍw��.󽐲�3V���1����y�6�u��-�Mk��@um$Q�*���l��ڔ����1�:n=ۂ�g�J�*hl�5�$���-�ÂЅ��jΩdU��Rژ�Q\+�oR=6�;s:<���bGP4ؤ+
Z��A���q"��X.�w��#7X�'a]��Ƣ��>"u5n��ݒ� b��[�������ۑi��3fk[�:�&	�� !��4�*)'��Q�>�
��Y��q4�AET��Qwc��b��&��
��[X��&�WcTCWmP�n�T��� ���F+c]��jn�KL�T4PLUQ-AD�U4]ۡ�D�֐���*��U�4Ѥ��#�!CM�hu������N��b��A��ǩ:��lj���c6ة&�m�pl���M8�"d(���=:����6�I1l�;h*�U��F1��������Z-kv��we�Bt]�LR�U=j��gV��pnΛc[`���GZb�F�rƌ�0kN�*
.ب�u�Q��"��U����������#�;`��b�"b ��*�((����-&�������&�@��T��������]�j��U3;�ؾ�V��t��3�[������f� ���4)a�Y}���y�R�?n.�N���Ro��IG� 0����2�ج�S���q�W)Cz��6�<��3��n,��$(��%��;�t�{�&�TI��ӕzAy;�������f͸�}���-�aL�&O�4eC��^����5zt�W����$�=j�Dch��;|8�U�g �&|�&�8��W���b{���b�����#��Z҂�g�M��H��bpy/�v�1��VOa��C���%���Ta
�66��o�\�2��W��O��ӛ����;�P�����/rbE��I��OM�J��龛 錹���Fnխ�h�T���7l;���76�S�q����ׁ���w��'��u�s��c�Y�Ux�ZL��y C�1ι���գ	���Ioˇ��^����gݭy�M�2���*/�W���� ��f+I�~�^�8׻G|���Rn;�A�/�ͫ9.��������Rݻ7b˝��mn��`�޵�M�V �~�Tbnq��t�\�aE�ʋ6���tSgY:���5��:��-��TG�r4����pc��k�2:r��[�|���7Ϣ:�;u::-��6vЅ����k�ީo_��A
�/-zme>���5�Mc~N�n��&b~�z��.�oX��=�{�:�v��2��Q��W�J���%� ���R{m�>�=�m٭<z������M�B+�U/N�ے
]�硥����7[���'H=;��(��ǌ�#��r�.!W��~�v�2�j�B�fx����K������M��x���������=��;�6�v��oH�ۉ����~�a�U�}=F��O��z�oug��=��6��;����~$}��7�����~�?6�A��~�tc��.���\�:Vj��W�=��xc���jnBAx#�;;�"G�8b�oğ��C|�J���x�����Yu��ͅ]�뾛;�{'��-�=7�{����)��s{�V�H㫜n=yZǻ�X��>l�=~g=�	����I��ަ������7~�X��@,���Nq)\�tS9���][fj�[����F���܏��=�B�Jmx~�AfQC���HfgYG'j�{���O#���+��YӚ��\�nݱ/�6�����4�;�9Pe�%�s��>K#���&E}G��XTo�%��'9@�u4�����+�\p�m;���UB�1yM�����^x��Oz�{�7�}��"W�y�f��� �o�)��E����6��O���nwK���=��G�+7w��|�W�yR�CY�s��~��uӹt~����~���B��7}=D+n{��o�u���\x<��n�xᬻ��D�k��b��ts�(����<|�:潨���>J��ԯLmOJ�S��#I�CD`�����^�'2�=]V{^A�٢r��}�r��i*��'�w�~��
���7�d�V�=ݯ`��q&@n����vΟI�}�ܷ$ێ�>r"8�=6,OH�n���wf�D��Di�$NF���8�W��v��E�VE��F�KU����/v��ֻi�ȴ����;B���+���E��[y��U��WyB��>��W]�~��T8|���iW.�Jdֶ���\-^�Ù�
�m�3%h��W;�W�����KB��Xb��I�Y�����.h�2��i=y�My�ʱ֯�������l@�:!t�Z��g,'6����?f,��rէ	�Y�ԛFpl�*�X�X��-�~��pT�1[�Xܒ���B�l@.��8,���?0=+�M�s���u9^����O�|�����]�p�-�M���v#��l�H�U�~�yS�P�̜k���Vx����w�n�Ӂ������������������FQ]��~�nN_�C�j��˞ʓ�r���y�Y҄��.׫�P�o�=^ͩ�vuc~�5s=�5���I�c�8�f6is��2��gbͲ�o�lvU	絒��U:�����AɻFұ�<���}�\�k�N��q��� �lu��d�{�c��}{�m��^�5w��@�z$�������^���]1yV�_������熷��}���>��:�/}�tO����s\ύ��s��[l���z@|��X�a���I�~۷^�鵙�3'}A�$>�_�����{uz���'B���UR�W�y����x�a9}�0�T�K.<�Y�.[R��2�Bc�式���P�S��38�0=�3�ő�7�-�&�ީ��s�w�.�ԍ�Ҳ�?�{#�^���;���0I����.a�XH�f
����̱�1��,7S��On�a\ qF��x>��,����E��M����Yx��n�o���O���SV�L�Ƚ~5oi��
C�Ӿ���9e�^u�Ǟ35�� ���lry�����Ё��Q�H'X�+({���Nl��s.���W8�-�+l�sٺ6���tU��P�hG�S�l2����NU��sX�k��Okx�#��t���I�����~/��#�b�a�<��&�'���r���T�1�5���W��}���T�n���.���[g��E.jM�]F�\��M��ҷ�jy�2z�����%��K��{#��q�z�N��N�� �h����S��Q�>p�ɵRg�蔎�:&e{�-;])/Fi�5��w>&���y� ?S\�x�\���K镎�Pk�v�d�3��A{�{dg?�M�Ni3z�m����,�RK6@u�h��X�m�D�2��;O-e�}�݉a5�[6��A�JJ�wa;�a�(.�����j���ԯ"�1�r�#O��wk&������~;"̜�pocoS�K�8>MS��o!rx���}�.`���+���jFl�1)ˢO/�N�nu�s��e6��a&N��K��x��f��]��7I�`�����y��Ԭ�z��sguqh���rf�~~",�\tm��}��7��q�u��[���=�AsԴ�grR�y5{�z4&
����CX7V�EnD����v��9�7}ݑ/��G4U�ٲZ��H�w������?vv�O;�����8:�4�|9�WU���y�yju��9��g���Σ�;��$%j�K.ߣ٪���Ճ:o)��9��7r�5si�����rsU���=����_�W@j�?S���=LO4���&(���1��\[�<��֢h3��l{1f�rv��[�:�ueǌ�&ۨ''��]�=��3E�����c�W����ˮ9'�GOU�3{Y�	�\Y�,6ܼ���?T�^7~�{4�d�>m���gM����,����M�ݦ��{'LȮ#�A<1�CvP���k.�C4gi��c��U������/�#an��C}���xy���ķ�=��j3�l�)�c�y��4����������, ��p�zG\�\j�4���D�;�k~[�� �A2�����oAH�8㬚6�l��1���l�O+Ͼh�ϞٛC����<r�v��gF�F��OS�7�le�=��L�/�Q�H��V2�y�&�!6��'{u�Z�k����z7��"���q�}��s͂�T�qg�R��ڻSl�{~�3f�&�o+���aN�I/�bF��n�p��d���귞ɳ2n�j5+�����Ǵ7�;χ�-��Jϖ1m���s����S�xfR�{V�zT�qs�9r��U����#؋�I'����k���h5�7�����K�a�{��R��������[x�g�� ��;L~T �=�Eg|Ӎ��nܨЌ�x�L
��V����%$�Ye�^�L؎%D�Ͻ�IԢ��\}�d�U���Y`��4���6o_g$����q�d��Y�6��O��ʳ���4�W�({;��=ځU�6�s(��J�CNb��y.b���v	�f; r��<�&_lKWwK�Yj:�i�����mо@��st|f��v�ڳP�\�q�F�4�98��sXjQ�Ӊ����I�^�@n/K��~k�O7�͸9�=�d��:��z��3��Z�0ΫF{]��0��%����
�__�^���w�a�jЏ�_}8<�Wj��Lu��uޫV(CI���9��S�U�[Sq���eb�c�=��ߣ?�߇X�>�`ԯ%���_�RT��m�Jv�Ai��('b��.���v���t��a�u?9�w��]�Uwt=^j�vf��{_O��'TZ�
��1[�Xܒ���D��L9�څt��A������Z�*�{�k��	�7=��rsM��x��7�Ϛ�;�1�wy�p�+E���n��{5/K������Y��ϳ.��̊��z��=�7�<�)yo�֙�>��>��y%A�t�o�w�/9'��9֯G�L��2n����/`5�y���8�ើ�;M�I�`�}}Y����[ǃ����Ĺ3ꩭ�y8W
��ߪ��[�x�����p���ʭd_���9�=ܸ=ۛ-����֟1����˒[�˜j�vVe�� ×�M	D���J���Ս72N��f�e�{ ތ�ʆ\�_H�H^dV(Զ���8*�w���Ī�鬕�a��rS��X������sd֐zI0^I�� ��~.�kV��/ϳ�;��~&5��9�x���36�LU^���;@��6��M�0]��M�����薯kȵ���fޙ�&,���hݺ ��E��{{f������Foe��$;�������|j�m:I<���|��n���eK[��/&��B���O��.z�z�kG}�PK(�8���K�:�� (�Ia��訏@5 ���)�n"�#�6ؐgr�rl�qm��Á�-~�FT�7]�c|ӧlH�t:Cv��>�s}�7Ľ��ʿx�s�$�BT~PI��O��R�"�4 �26����r\1���%?��<|pS���=Ʃ.��R`͏u�٢��y V���%�g�,ꕴ~vQP7�v�z�oUg�����oޯ+�gk�z9u��ǥ��ԩivAЬ}�����g�q3��֮�ĥX�i��q���T5�Br�v��y����x7,�"�#����Y�(}������h�Z7��܈��d�i��Y���x��׸^FR���B��s�o���yk���.���%���|�O �n�@և|U�3L�vL�d��m��'�O���{�M��y�n�� ܟ�#� �V��v'��2v��r��)��� �:]�'W���΄��z��.��|z}��9��X}�7���D&�86n~_ߜ/����|�Y��Y�-,�M8���/v<���������g�i�m��V�{�fi��sְ��kO�/tس�_�l �w����=A���{�7�[�{��ʻ�vo2�o� ��ޘs���+s��g����f���?W�5m.�֨wK�}�ؼ��ϔ�@��|�;�g��vm���=5�L���N�{HS���7{��DN)�њ<r)����c�gً�#Td�ߗ�!��j�O
3�g-��x�Ij�oDqi�3umI]sg}t�*�˥�)����4� 9�G:E��U��o�荿�sjn�������9�<~잹�������l��71:����_�C��g��2j|�.��P�=;������ΩV�!�2�����Q8�-%bL
(0�V�u�O3H�V��)���sx��a`��M�ݏ �6_�K\̴�`I"r�&l�aKA_eN�k���<�զ�x��:��֙�^���5i�����G��iS5Å�`�brO%����j6F%�{z�:�H=��߮����~��o��yR�{E,S�ˑ��l���.n߰�I�l�r�Ƽ�[>�y�S�9|u��I];��o-��N ^P����}}����]��ltmmm]�Eud22�E��`��nn��fK.��ⷺ�ik�%u�1�5�Mn�6��P�s�sB�N����( 1�xw�:.��|U���;���&g�1�`�M�
��{t�o�b�+Q/0���<���4lx��B�� h��3��Sv�p͘�ˆ�Yִ�.x��FZ��FV-��-�'G�q7Vl��*��G���?m�g����&�͈�	G�:vn�@�F�q5�c�W
j��wX��L���>�*[���q�K^ι0�7��8��@W�	��_@fk��C`e�)rj� ����uբtmG�	�U��/x/{��F��W�nǽ�J�c�]^��V/�Mڷ׭̷�h��8��JB�хq}�b9@��fA�ؕ	u���o�Y!Ңb��^v����ᩋ�]�]#\��1����}u��>Ʌ���}�qN�⣃b+3U53�%��$^��ָ���տ�����h5� �3����Ш�P͊ ��V6{�߷���>#5�B[��z�V��!����Fe�=��o_s{Z!
���UZd��0��e��y�����w�z\�Eˎ��/3����T�r �ffvL��~���.�F��O~�X�]�]�`cU��O%�G���1���_������
Vu؁Bg��ΫW����Gn��ƅ����QE`�Kh( ����(��CQ�k�m�TW_U O;*m>�Y�*Ɏ^�CLj��t�`�r#��r���VB�Q��
�H�E���Nܻ=�X��cv/��F�X`�ĝ_ز���)M�*�olu�I>/5��9��#]�2��y�m#Ӊ=��|��^�P��E��{9��4B_��3]�y����n��QH����ޏˑ�||Uo)�z[���MB`��Ԏ˾S�έ���ŚK���9��(lQtͤ�r����O/��=��������vW��200�P�#fgT�;�g\5�$0����3��o.:���ݰ-�X�� ������ד�YS4�+�{}*t�X*�nyj�p�ol7u���rl���j �cܓg+�}�4{ľ���_5��x1�|�/,\�:,	�)�鵅�Rbݼ�Bx��Sm9�ƥ��{,>���&�1��W�6���G���q.�B>Sv0��9��y�z�VW�I�A��{���g�|�|�j"���)�� 1P1D��G]B�;T�[ww���.�'M֢�M��::���tV���[W�Ch�ر���h���(����EU�z�N�z���O���l[��6��u��1]{ZM��{D�:J(��6=�����u���u{q�bk�`�:��^�&*1�I�w�\w�pw���rV�5l���`�z���료�6ɶ��b�Pc�S�w�F��Si�Ǩ��F}O��W�w�h�P�H�����*

��!O���Κ�ѭ�Q0E�������j�"N���A�j�)(S��1��U4�����(+z۰^�h��)�=������CZt��[������^�3A�
N���Ӣj�34:4kE>���Q�@h��H�����T�1%�ݚ4�Z

h��M��t�+���PQ�{ӽ�ڵ�k�;ssL�"���+�Y����k��+�ԐX��^uɝ�"�A��A�P�Q�����xݥ���>8���<5�rF�t��
*S9���m&���ţs���2q�O�eL�jۗ2k���oő��l��/ry���)�3��2��m{��l
�N�������Q?g[��	YX�^eǏy-<��Rj�1��7��u�\���� �c��ݢ��hr�am���|B5���s/�z��<ozU+0ۼ+��_��I������vXțaԵMP�R�ᄇ���ݬ;zf��蚜�����6�{%�Iط������|ǟ9R.�4�e�t<�YW@�����ؚ�fu_s�U��[��x�A�PY�L[�l�m�Z�t�(AC�XMT��Ლ�$`���<����d�=:$2ܽEp���xV�	�N���I�(נ��{��!��fò���,Z,��)�ni��=�!�Գ~tF˲��;�
~R��peR� ���اՉecj�s��n��тf�����|��zD=�@X�Ȫ�&��G2���#�_ny]�ޑ��#����-LJ��c!�.���9WA�hP/��ݱ�����P~'}���&����f�j�͏�A/�C�D��aՇ�����3�Iڣ��lc8qZm%�\Z�.%����[��R�nS�]��-�f�?X�����ˤ�p����+�(��!	�_0iwL���ǡn�R|�sd�&F���o&���r��Y�C�-� �}���w`�����;� �v>�P�$7ﳮYٖ'PTF��Оb�%���lT���T-��n��	Mٸj�zC&2a���a3�ǧ��8�Q/�� S$Q�0�d@z� ;ZGI�U}wv�S�l���(�u��_����z��~Wz$f��p�%}Bp3k�����	�������20��)q��ؾu����u�E8�`Sqi��#��3�~�t�#��b�9^!�5�;��P�q:��/"8� �.�-�IW���`�Zb��R[�)L�4�lc�|�ys�v�]�yL���KJ��!�j�mN #ӽ"��;�?E뤮@8�^ǄGg���1�n�G�I��=�o���o�b�����hְ��tY?3��͈�.ӓ��j9o���"�����MFϹ�CwkaI=��D�����Qj���ɘ�$̱Ӽ�*��TU�U�ޗ̗���a�3�Vz8��ˁ��������`d�Kj#�T�u�4��F-ڕڪ܅�`��./Ş@�ˬo��\�\8e��"��Y"*�ȓ?_d��V��#`V���_��|z� ;��V��v���7e3F���&"6�2�7����Q�Ҳ^kF�Ҋ��^,�o)itҷl�֥l��o��Ry�K��.:u8x]s=E��g��gn�Bڷ�b��ዂ�eeZ̄D��9�����~c��L���T51g��#�<w�F��;B��Un��=�Cp3��W��c�;;���h^$�}��2!w yi=SgJ���N��b�k�oP�S���8GƲ�u������,��qˍvm��0/��7��΃�UA{[ ��}�c�ݒT��T�n33.��v��''�e
��}�S"�f=��+yH	� C\{:s�<�*���3��|��K6w0��ݺ�T�P�R���`QR�vtO6�
�h�ZT��/ld�B㱀�˅27O��sYL��v�u�y�׏J����r��xwli�:��r2U��B���n\t�֪Ө<j�g\��@����!�uu��l]�U)q��Cy5,��a)���2_�IO322��R��j/2�<j��54��h�	zb�������$������ ��-�Pf����y�V�F#�>���tV)�A΄��s_�I��G�(����}8d{�)�]-���W��a���ȵ�82��^]�1�솎P�7�F�]��"�i�d|tS�F�j��^�)�Ȑ��k����)���7���6�Ee�I0a�v���������Hv�v�������b��hO�v�nNws�V��:}�5�7}�1��N���N�/�k��}_5����{�o�(�e�*����+�F`f��b-%�S��f�1��2�P���4,W]B�[���>&&F�=��h*�5{�nY�PQ,��=>��DO�N��.�8�F����k����o���^�X������O��*m�O��gOC�]W�%����N�'�������duġ?z��	
��}�{�<��T��,�eEB���~.h_M$}��DF{��}[��]��.����;��������}�5,a����y]��r�'��ÙW�YB��,�$r
����D������z��Z���K����# �����}5����m�%K7���ni"��z�̈́;i������{�H�U)�J�[UJ>H	=JD.�jj��Ur����R�:�7s�+D��w����s� T�m����:��8,��Qy+א��P}�N�&=E�q�^�$b�j���ڹ�wkt{�2�%�����%:o�n�	U��-�����p_�@�J
���y|�̏=��^^L�#|���(>=v��������4��;�~n��J�o>��v{�]Ѹ��F�˻�gwi�!�z���~2#��N@��g���r��Ӝ�0	u�H�ޱR�
e0�sM��o݄�?��5�e�H��Z=��b=x?e)	�ȏbW�j��W��k�؆���K��~��i��f����\n��q+] �&+h�U�cO֞�Xْ����|�{��7��>B�'�X�J��������w��ă|c"T�	�lh��PS��A^z�BK��	�7���h��F��b޳�։�պ��2��g�]�� e�d#��Nl&M��Y�嚨B��3��a��̟����ܬ~����}��`Z� 
�M9j|�0MV5�`2]�� �鴅�+6�����8�Q�>����0#os�!��̃=��Ǻ����ؘ�?G۳-8	����<��1Z���jU#=[��_�tg`)딊��t�Y��l�=��@,�dP��3P��^�m�Ӟ���2���f*�����x��+c�Wk����7�Ӊ��J`�����m��BE�����d�3ֱL�dpۿ��k�/����Lcx��~���k�f��&�'o�~JPm�l�lt�+�z�U+$���	�_����6Y�}�"�z��+��(����}�O�z}����R{t
�9N^��������5�q�͏�ri��:�|�-7��_O��ꐐ��T�r<z�`o;f�'!��22R�{;93qr�@���xaMK"X��[T�`��k�.�w��Cj��yQNt� B�hfGq��}���n�`�A�4�DSD�%���(掮 �;X+1�d��gk�sM`Ǿ�{z.���v�p����F:�f�2�n��V�y!�@�Մ���Z�jP����\�fEr�Y:֕;�M�;�s�1��sp�Bp����VVG�&Zb9�^<o_��E�{������1I�|]��)�ENc�����z͇�WI��5U�A��[�U�^F����N�v�#�v(����T�����B��V0օOT��<�J.t�y͡Lu5é�^��E��K�G�@��r@;�'����*/�DR}�I��=D��e�w�ɡ�L!E�'r�3R� ���2Kt�Ȅ��h8`&x��P���U-������	�����}�:���w�}�Mj�U{'��w��$�*Ȳ#� l�1��f���X�>���6=�g���z浯����˒�.��4���=g_��B^�n�F����<�Q�N��/�v_{5O�v�����X`Oq��[<О�l�.��k���{g����+�Ģ+%���z�ڽ��������Գ6���B�wl�;�H�~�����Q��?t^٣Jug,���A�I1��Ԍ|�#K�m����;�u۔��(�p���ky��"�4K=�v�
�+�޴9w�,XZW��`�kXE�~�?@\w�TGb����ش���o���7:�5)�� 5<.W\��ld���p���U���3�B�y[��+�E9�6,�A\��^*
L!�pW'R[��^Ԙ�NG5��2��p.rWi�?����JI
)�z2�·-�"|�U��̧����fq-1��V��:����X�j:Ւ�Sz����4HK�����WD��d��}d-~+��퀘�f���;#�8~9�󷶏WC����J֓o����S�vE<P�դڌ���W�c�t�+�!��ϟ���)�M��7�]1��xZ�qM�V�5�j��Y���P�mR%����I@�$�BT��yM5U5�X�;����v8/�Y�Y�|7���"�C�?�h���]����~:l�2�L`��،럸�t�q���;���^D|Vy},p�ν�Ss�!�>�|{^�ؤ�x���R�K�i�Z�TʚS(_oT�=I����|b���(@��U�+�-���5y̪M��H���W�a���70{�S�4x~��4�y������w\*L������q��Kv��!��:s�;�$���e>�\Dw.����W�����o/�V��x�&t�HEfrk����_��1ۄ�T�qO!�����z&��):�s�6���Ԅ�k0��!7G1��R&gfҮ̾���ƅ��ԣT�:�{ٱ�	�U�,*&�%��<-CS>5�wg�7�+��+�U�*eO��k^�ًuo�s�g�j�Vxz_*�_zl3�7���T���d��3�:�C��;��@5��J�z��=S����ܺ�HE�<Ȕ��߳
8�!��&��}Dwp�;��y��m�k�W�*u\��{Y�A}�_��Z��BO{�p_��d��y^�w��\h�BZ}�C|�ȉ�\����8��*T8�Y���#��ZSz�{������qć�}ȃ\P�2`�ncz�*�S���S�����{�1��řk:�q��t���ˉ�/x\̝2/�~�d�.%���o��@}k�l&�1��XʻXr-"f7��SN��ag�Z��5������؄vF0Mꏝ|ըv�oڡ���j��x���Qᙗ��JzL���f@��pY�u�¤n��c��O[�)p�L}���Ig�'}y+)+���\���HdO��f#�g�w
F��KW���y��oG�=�J�_d5k���Ei芒APl�<�� +��4�gk5�,n��ÜjZE�L���A��H�_G����Q �H��l��剉�F��W}N$�X��=*�!�T������Ƽ(Ih��o{÷K�ַ�H���Wҟ��E��}[RڌR��/:<d7L�C�Md׋V����˨�,����𥙓Z��Ji�V*��hK2��ܧ����>�0��, �Q�4��J�^�}�{2�jZu�Re�_��o�Ɛ���O��W�Յ.e�N�m���۷�X^	��]�GӚ=�J��r����u���ĨE~��˜��Ѧ%��62�"}�F���˩/�`���]	B�֙c#��f�׼9F{pn���13b�;�cw�E�<eǐ�%0&!76�SL����L+�2q����!����}׶u�	�����{ݮ�|���inxN�q�t��SM��rq��)���6jt5uΑ��3׍�N��4p���Ɨyz�,�Gj�N�L�~l�~l����F�۔�w��a�Q]��&��$�Yz���NEe���'hE*�;'%�`�g�*YTp��N���yw�ΊՄ�4�b>+q@K�0��M�b�[d^�-mc
UfdrMbӨܝ�9��<(���
���:�-��T#���1`��d ��L�\j1Xф^���\�9�͒ao~ə�>�䨧��_����j&g[#%םZ�O@la;�)�j�5DOS�p�+�y��S;��z.��5�zf��1�}s�lOѻ0R�8��&������l:���3!�#����Z�R4�.�X ��Eσ�E�#"Ʃ�ONb�;	��t��_R��J��;\&ٷe���ץ��͆}���Z�:���g	�G!#��7�ظ�̬���.���R4æ���,��x6h�S�t�j���}��[�j���лN�g���p�y;�Fk�^��]c��'���*.����\u�QM�mᛣ�l����kg~n>���|a�t3Lxmc�ه���/�Ӓ-�0���r��,�$�RW�3�yLK�����a�m����C�ƀ����o'�Ǽ�O�����<`-م�%]?`p&є �.�j&>�܉��i�*�_d�VV#&3��t�=�������r�fע��B�0j�v��7�/j���-�������o�'b��}�ڇ�-�</
͖)�\N�v�Lw��}�ư�z�f�$� {k��FuƿSe4�Xn]�J��O<�P�T��C sEU��Yށ1I�|���6��S|�fUcm=;_,UG��Wr9Ws}������^3��������#�B.(9�I9OI���^�]�9�@��y�hu��A{��MM���%:!n�������<%��g��9]Ӥ�٭#�zO<v���A�%���oI�6�X��Z7����5�L���>�����Y��glgm����Y�x�T@�ɽT�\�����-˷F�oT3�����"�.���G�,ފi1��YC|��$�	����#�S�M���tG�ǠZN�^�D�*ˣ�|>����}������?x�ԕ<���v��CVd͛�J���:J�C:H1_]��>3�v�NX�\��`W�0�AК;Z�����J�e]7ʖF��������U���i�*��]-z�Xu2�h����7��Ǘ�)�'���=�3]EOy�q�[�R�q�r}��j�	�T�{�옋X;��8b�}p{����Yƞh9ya%�OKi#[��Ԟ���v���&CX�P9�t��z�ٷۭ��շe�i��P�2
͏���%*ac�je�[����=�̂[�g-�_A�����7�K+��4"��"�Q0�����Q���Gͮ[eJ���lTD �a55
v����{��3IvOh�(ڛi.�v�,|Y�Xދ�ʷ��uJY����_�y�C
G�/}�W�ҳ}}��_�{��^�<���#c\����]��*DrޥI+�.`fJ��hAÈ� D�M�����+�-d�{�G����_v�4&ܓ8C!�7y�f�T����Ӛ�\j�y�Y�X�/�*ܰnr�s �Y���J����k�\2�� �Od��c�'�<z�7�Yy�iQ�<�hI[�{��_ ��g{ �Z0��ð��6<�����Jt��WwKK;b\�j�����2|�x��௔]������\��.�{�A���Q�hP�u_6�"��A㔴u9�q�(�U�*5vn�a9��"���c#EΏ��\��+�ϙ���[v_N^{�J�l��&Μ���c��):�Ω2=�L�G��������_l��A�?�vm��f�oPmCƯ�F��С"�N�K�3�73KD�qJO{b�1�Le]B{&Z��BG��:�b��'��sx��F)��OG�W��O�=�<���K.E�.�яy9��k�GƯ$�PÛ���O��z7Z���y?�[0�B/&�'|�eI�=$��:r��aV����I�&��r}D�]4�� �8kzY��0Cs��띊t��+ݹsS0��jQ�Q��sq����ʘL���s�[�9��t̚�o��U��^�n �徏�P���-�2��o@}x��9�x�S���N%g[ܣ���[���fjF�����7X3�fʁ��un�墥E�u�L���B9W��ŅX�ծǵ.�sOS�Y� F������\Ħ ���>>��8���s��1\��`�'^���i�xhn�AN쾮a����۶�t7{�b�b�����C\�9w��)u�.��hŏ���ޘ2�����V�.h�(Q:�L�@.�贇}Ϥ���ʧ��T�n�[ׂ�TPMΌd�G����Tf&�#f��w��l/"��:�`ݜ��!�l�8V�ux���4���u��p�5h��Q�R�r��n�{Ev�\�Q�ruқՆ�\�ZCݗ��Sy��_sO�A�y�v����sѲ�>�(�P�ٜ�f�L�������a��2�.m�^)�5:.�K��1�;������VI����0n����ǹ��ݖb��Ka��Rv�;e��tu�'G����LMCzƚJ�f�;��ˈccC��b$ѧ�W��#��".�u@��E�*��>�d��
	���gHEZt�i�)�Ǭj	�4b����cQ�����
5�f�"4���+�i&:IR�PZ*����4BST�����K�����1/�@�T�D$^��)�C�!�tP�HЖɘ@���ioY�CITi�%44�T�^����%��']:����j�V�"���ѡ�v����S��C�()
JI�J�gX�R�PUt��C0SOvQ�{`�TE�4:^�A�JJh+I���6��ıh�D^��LA��(���+������E���!n��A
xn�g�BóR��3�Ɋ��r��8T��P���I�d�lX�+Wf3]�f�ͅ,}�F�H��[+{ܯ���*ޞ?�?Ю {�3����t�vJ��ml�Bz6}C��׵��F�R��;%z�)|jgݗ0��<�%A^Ն~�2��򇙲:�ÃZ�u#"ۏ��Us���<��ֽ�{|��k0�6)�����h��<d���L��5�a�T9�7���<�-�������t	�%]t��M��v��.#Ԅ�~�H�	_HLL.a�b����PM��.~"�UTV�����k��9����r�k r�V��F(J���yP�9���~~9�����ne�_�p_2� �MKW�A!�%	�^��E�IWN�(ͻ�mP��̋�h��f�f,ط�ˡ��1�b�4��hЃ(z�<��h���8Iy�P�h��p�����˅�WՓAx�Y"�"�#[r���ʛa@f�Z��eAv͗�dNr�a-��KL9���Ӊ��܂&�����}�����5rNH��	�:ה��2�hh�ws�o]V_5�҆��Ɉ�SyHO|/*Y����?��m��.S8�nY��j��_���o	����4�ģ��"aI�)ٚ���o���HԤ�@�eH;����|��	�҇	��MF���o��5�o^!�W&j{��@e�����Ԯ�%�, �B]c���\V���|h;xػh�����輣Uf�[�ŶTp��ˡx	�����x�v=�%^�lb�x��2��啲�=���_2C��V�W�'���U�I��o�����S�Fn��1y�h3^�&� BN�<S.~�z>��̋�s��
�^E*>k�b�۱
y�[e��L�Z�'��ೞC��4�P�R���)�gB��~P���F�g�߱cynf�cv�Wo��ܼ~~7��B~7"㚤
Q�.������'k�8G��{�la��Vfd���n�C����Ѫ����!D�-����6Ӹj6�v��{��`%R����3	���6��Z�!����^}+sXM��U.8���d�{ɋ�y^&���q���4�FJ��9���4^a��J$�¸��T�u;3'�:+�����&��̀�|D�d��ܹ�Z27M���ʥ�jn��Z,�B�Y�4�6=��o�fcL���vF0Mꆍ�l�"�1h�S7�u�]�W���KH�t�W6x$:���cp��x��{��~[�)t�pU����p(�����Z����C��Y��qRoi�h��n�c�0S�{�(7�C
�`��3��y��+d����xoj�)˖x����� 5�?,P��e[�7oA�Q\"�X4���n�� 0[k��V�U��=�x�,4{�A.��M'�sT��rM�N"���:�m�L��4�ӓ  ���4���&M���x���ǳ�n�;�����uhr���UZ}�/d򽶯��|"%�[cXO��騳�{����3-�VzWy�>�,7J ��8F)�K���Uk�/����ozQPѫ����K�j�m�4ߵe�1����Z�M�U��|4/����r�b��Vl�P���>2���=f�����o��8��]yW�_�{����y����X�����'�ݕ}I��Ve���)�����ؤ%T�%'�L-�'��>F����vN5�V�"tُ2��L4�&�Je�����ꩢ%wG�=4��C�p�;c�r�flX.حv��ی��E���1��r�]��tüUJn�U[m�c�56���--L����G^J��L��吃���BH��Y7ax{Ƒq~sJ�|�X|;nZ��/yأމ�e���1��J�å�E@��=/��������<1�v*���&(EqU��n��s.wڝ�o�S�V_.�ۯ�d:+�ēؿ�g1�/Hpܛ�}1�z�t��C���᷅��"5c/j��E����gL��P�O�X'6�@Q����]gZl�b�q���¼s�S���B͎/)_��x�& W�nl�uó��L�����g�h]��!dz�QMr�6���cOҞ�O�x�}}�t�ux�$�U�8+UK|�;}�4��)�۽�87�C70\TܜT�ǻ���^����ٙ����1�����G.�k�5�|õ\���ޟL>ft��Gg�d;�-f�Y���jr���k�}9���8\#k�H�8�<�dc��*��e�¸���vKhFֱ|�6&��e�t�;5�*G�}0���zz1>3c���C��F2/�Ҟ.����f����ڴ�]塵�\�ոst��ͣ�(��祘���0�o:���]�`n��9�w�@�t��u0�t���<�b���z�O+������!ڪ-mX�2��}��ӊ�����M���p�-��ίob��[�v����ED�<f��;f*�+⃵੉0��ʹ�f�X�I�x����띎�778��%%U�ʆOG31d��&�2uuO��P��i�g���Y�Τ�9Ⱦv7�oo2U�mB�
��沮�^�*ֱ�eMb�%�m��]�מ[8Զ-� ��"n���©�����Qt�L�y��V�j@�4��_q�������ث��<��H��Nc�1��i���Ou]���)��л���K�^�K��4n��=q�@�Qqa̪:�)���7ɹ^�?����*V��	��5�:w5jVڐ���>��pX>����Q}��>1��{iGѳ��1��K�{e�{[�Ŏ����J��u�0��S'fr�L�dY{��ru���f�)\��tK X�A>f�[�u����|�s7�$z�0H�%�wn��_UUV'݉?M�ݕ����Mc��ǣ����#�c����U�Ta1�^�Je���7��1�wO�l��;(ul �):�*��,YE����0,�|p��_�$�����o�Q�urv��Es�U�t��2v�ze���]bx�E����H��},���VE��Ȅ�}�j���/M%�o��c��`�9�*D����-�z9r�K�FK-�9�E��ᱎ���.�d��'1svg;^3|����_,�r�<�Cw������u[����k�����|����&����ٮ�Ңx>*><�韡�s�)��l���is��dS]!DRP��t�4���]9~�e����@�S����M?��H�צ�.��)�[��wf�ե~(�S�Mm;����,L��RXej�P>j����k�sӵ�L;�PMK�q��+Q�
&o+��y����}�1t���#��ގ3���ai^�b-@Tg<�B��9�Y��-)̭���lҡ���Dx�^�]77q�Af�����v].R�q�\�ԥ�iV��ʛ�0k���{��q�mn_E^�\lJۧE+�D�ʦ��:���q��D��ձ��%r:ؾ�ɷ�{�;�=�DJ�s:0�Eg^l}��%:�.|���(�o�E��� ��Ւ �Zai�{7��ۯ������V{�L��?�N���N8����Xʪ^��A�=6׻�LK��<$�����I;�&��+ʇU��˸zN_��H2�4.��p[r��ϫ*m�j��e�c���_o�e
�|�Nө�xM�U�������Id�<��p�ďEľK�-c�'������8�X�d_o9�p�p�)[�"���+ܶ��5���ڲ���j��m�M��T�A��[�h�ڭb��i"F��yu�#23g��#W3�/���&��b����Q"��]+HI��3P#��Hh=�^�ˌ��K6Vg��$�A���=�(���I�'�e��
�l�f�m�1�O<
�R�TM�=Dwp3"&vM���&�]�T_*\�(���'6c���q�q��oGR�|��8v]�p�����ݦuמ#�*\Bc^p[��q<���N�vlӋ��\�Ƥ�Y,s<�C�2��2��e.��I���s��B�g���!�X[]�l	�� Vl���R�9oT'SK�䜾v���!���s��OoE���b�5sJ��	�\����jsb��LwQoz	:��_WT5������E��i�-j����,�̧��Ө��z)َH���uk/�;���0�m�_{�����cF���<-��}y�G�w:�9s�aî+r�ZO��A����"|�e�3��쇊�g&Z�vL�٪�����.t��>���{� SuW��"b����T���}�]OL��#��\��D�LG5��Ů"�aI�. �>����\�'R-�hmr����P��Z�����z51�솎��&�CF�]�ޓW��ࠞ��>�D���̌?
u(��7�E���)�b���$��;��AK��pU���jn���ɷ��@>)�$Dd�=3Qڽ�eB�Gֹ'�����	p7��EM�i볣k��@�x��v�3�>�k��x|D5Y�O�/�O�fF�&����c�Jm�O]�[!�
�{�����p��oM%���(�i�85��e�{�"��>��8�:d���bS���J�oB+��������}�X�s�+şm��kNy�����)���2��Oފ�ɱSI���yU�`�,��[4˯�k{i#��+��5T�␕R�����6'I�����r�S^�p>[���'3��_<�&XT�.~^�6ڲ��e�U�7��>�r��\0O�7tHPLM���W2K��0z�!�������%:a~*�7vy*��Y'_����^�͚����O��ܻ�I�xo{�k����M����'X;���i#v�����E�~�H{�~}�Y�O�y���*)͠�?��7)���>\�2�feK+99�b�.R�o�yqc����.[R��-��aG40�~�q5�q�1Y{����5}w�C�i�A�ZD�	I�{٘���!Ʋ�@P�T��4��N�_�#�
��w�W�O��\���΋���e��@X�ܔ��m�?�-��jo�~���Qf��`�����]$E��V*�A�O'G^b�RQ�Y�$��.>1�}�l�O�����Li
�g�~F��ߗ��,�����5��*a�p2:	~nYжKj�%���ɉ�� (<�U���;�(���t눟Ƭ�����Q�{��s½����ɜ3Z*��(�`�&=��/�]�7���pXi�)�gU���Ǒ�5�����g݌��"6��Ce���a�6���Ќw�V��5hq�\٤§�@us k�TM-�Α��b�"�� �����N�	WBQ��=�e��r��Q��!��^�� �e�\YQX��g�ibWK�9ݏ
�v�������ж���&l�z3u	�?B&���З����	����|����[�rw�I���M�H5g)d��v��$5���H�{�d)�B��+�c�-E�nC���x��?�7�2�'�/u￟{X�V�!��3^��0Ebf[�7�f]��K���\E���[�t6ܓ�"z�������t��q�;�/F�"��7a��qZ�Z��jq�qЖ�2�Mq�.3aa|#���!/':Xj�U0�ƀ�T=v��򪾯��xm۱4oa�l��M�m�|;�רX*X�=Ѥڟ��$��B"�[�n)Kڧ檒s�H�L�b����=�*s�wΠK,����+*�+�+^����d��Kj�l��w�Ӯ������C@W+1[�܇���'Db�?��=	�E_��M�6:bN=�b�����I�r�M��i7=�{Tjt�f��lИ��|���%K��͞8��K�\X~�K^��/dQiasw���.x���[���dG�(�x�2������:!o��*��mΘgk��[��4pܮ淍Z��TX]3i��H:�ek5��ʛ�_Ph�q�	�)�;y�6E즺��Orir4n�4{ٱFE�uu}�?���W�c�چ6@nv�Ϭ5�κA�4��|���f}��vEr�u�/8��H�����&^�r�4����[�g�hE;�xlc����.����#u���c�{Z �L'�y.K�l_=G@�V�vl8���6=�f��-��
`S:�)�c��:-�2g�+���>]7D�ϊ�V�� B�+��q�ŌZq�$hc�vX��e231�
��[~˭�1/܍�rl}��R)��\�y���������k����ץ^O-�Q�̝|��qJu��,ީ�n�)�����.��&�r̍�
3��s+��7��-7�9��19�$�4%luE��������q�%�6�������o=�t�Q��	l
0�3u-�O�3��j�=��^^3�ӗ�X����� ��Jw�H�ny�՘�+��0m?���������)�mU����Y �sT�!��4���3��,�AW<d��r�ҽ��Z��`0�Z���.�,�E��Ɂ�3xD�5�����m�f3*3J��Y�a5��E@�%��G�T]�{��v��E��C�V]=d���<�%�SP�܎
Z
���jeS�����h�� :	�X�2��-�gݓ]��J�p���	���|n����56�|���>�1���s��S�
���Z/K�-|#F���"MߚhP�h�F��_XX�)��yO�b��0B�>7<9¢Zx�cƯ�"�n�5Ӡ�ͧ;�&�%X\]���,(c�.m�M��P�3��,ψ�DY�c�{����ڵ��!IjfRtTywZ�V�fe��*�M+HI���CޅJ|�j��nj��঺��0����5i2h�3P�Q{��$���1�8
�j�T7A�؉�&9��χ���~__�����G��������B$B���r�s6V# �u�{�4|T�qw�!��Hz�9��Ι����F�bT
pAF*R!KE�R;Y��#�Ձ3|��^���1;�r���W�P��p��=���Q�L��.�z��Κ�*�4E���/�1ˢ��8�W��[��Ԯ�v����Y�R��N��|؅mY���D�%�Ť�G�فE]��ֽ���q�+@O�j��CH��5�U�s��v���qzu�	Y��5h�Y�����
A��ݘ�g���7�᎜fy1�(y�K�.�Q�-^��L&YW���_��o$��Цi(x�0M��x�#	b�U�H�{��nإB��l�7ˀJJ�Q;}դ7mYWf�z���dS0#�yƼ�� �9��r�$n��5�����Y�c��
׮"F�!Ϛ�{f	�;�9���uow�W��ʛ�-�d	��M�[���<�`�ڸo4�9��z>��|oL�����rd	�o�}Ǐ�]�ڵ�}��%�mM��,˘q��+Ei����˃ޑ�����wsl�ޔ���8�Z4�N
�E�������}�N�K�e�ؖ���%�Y]=���������o��׸�M��!�]����.i@��E�
�h
���9�Zݒ���ٮ]��ԍ�ڽ�z�C���i\�%d���k�+%�OL�����s�q_w�u�{��Jj�Ku���Z@_��F%�Vu)��tH7S-R#b�Xn��k	;�˛���Aۣ��j5Z��f���.T������2�T�L1�-t���Z:��;{�i��Ѝ��e��o�v��r���E�n��s.�R+|M��Y�ɭ���7*Y�E�$��ի�h:`�S����ͯ#�������툽������xP�b��g��.��.Q�a�J��oXz�싒��\�&�Ջ�cX��qMy�rJ+�wD��g�l�)K�5�V�C�!=�Op|{�j'��9��j�{��H|R8�b��X�Zj�1v�k���l���ʀ
$L�����h�"B�JͶ�3o�Y�Nw*볇�EEK�oYXN:�5,�'pX�Vv���N�\7�k�"�<�Mў>�m���өb۽?J�Q���"zvr��j�����{���wY ��ხ���$v֢4-v-��|�f� �K�ܼ�]�a�30���C��oS.>A������O���z��v_ �4�<�����r���B�yO>�o��'f�8S|T��yc�;χxg�g�&��p<��OK�a��ʠޭ�����Â��fv���z���)�\�����~W�w&nzx�h(jk��17z2f,ܰD�1l��o^�P��5��4�5�v&�-b���y���l����K�T~l�K�A��=��<���Ӿ��_of��*�"4�A�D����9�"��3[c]tRIKC�M�wX�f��`袀�����((�����=A�ViuKJ�夫mTRm�6�AEh7����(�+����A]&��#�:���u�l��E4[�������EI�h�)[�ZhӪ�
z����G���$HtbJ-�5S�K�jf�r��A%it�"����&
�z��Q�	���mAh4��8�ѣ��:�������7N���;��Ckh�ѶwN��w]E�Z"{b�(�ѭh4�v�Vٻb����!�-�)֓E�:5E:m�44��������&(�A�:褠��v�:zuK�b)ŉجhh�&�i�TU#V�Ɗ4��F�lcb�q'A��h���26�L��GyZ�)_g�����s�g��{ޥt�[[$�xD0����i���^�<��{m�������}�N�[�#�n�� x{޼��2���O��\��"���s�/S
��_��l>b��ǰtO6ג��3���V��������Z\�͢��!>90Ɯׯc�<���*�d4��mO0�����tqk�f��][Gax��IC[9j�e�J�&��g5
Ͻ����K����AmL�5骝��kЮ��E:*
q��K��i�,���x#��A-s�S��\��Y1��q^�{3]-�'!�e�o/jXln$j1��-�T��#��\��sM0���k	�|G�ǉ\��Lܩ���k-Q�k��'��q��>�=�{5��g�"��zt�!���z�4m:�oљ�o�mF���i�|#�2���vC�+��gef��XT��<Lozx��R�j>��e�}��WU,~��",�������pd���7��c8�U�t)�}������pbE�̙�r��m��ؚ���x��:<U)�\5kf�."�j����+i��/2d��.<�:8Ξ�g��W:��;�����?��X��������i"~D����yo����������1�MVp1���l���i����y���P�N9t���6�\P��nu�1-P�VE�9�uT�ٵ�Fr�ԦǺ���oJ����{�$ܫOh_K=:C:܎�%ˇXk��q<�����&�8��L,/nt�U�]�xg�����}UB"��,�~ֶ��HJh���n�,�6���b�}���d���=����|Qy�Юn���\�S��I὾�L��6�J�/ֶi�^*���+2��[���j��R��%o��O��ת�_��F�v�w�H��}����¼L�e�
�d\����՗6��Ȁ��=H�x�Ѷ�f]]ʾ^���Lބja�;�@�z}G�<��V��yN�QU)��%Vڦ�郘?w4�h'I[���B'��w�`,W�ߌ=�F���&�����+͎���x��g�nw���f��x���Ã�r8��԰�*��*�P��BO��+/ F�]8;.��~�Pɡ�g6��]�nv����B\i��	u��R;���6^�r�S#�ل����破��lr��V�����f.҂�\��0��z���;��u��7�����	��� %�M����K����s�&]9e9��f��w*)Ύ��)eyڤ��j ���K�k�6��v=)֕��-��!��O��Gj�S����g����1�~:Dl�{H��Z1�ڃ"&�1y��L4w�J*���g]�?g2]l�;�El���S�";���R�897��t~��ZfVX�*�=��ZC�n��B��t�U��GnG�b�w�gM>�qE���5�Z��qt���&���pWrn�����g�6nS��v�3k�؈��"n������z��Cl[3~xx�����=�KkR�(�&_��Z�q�d�`-|B7Z���)[w�#F�G�w˟jU�iկ��|��nzM�xv�8H��![�(��[h�H	�L����zY�yRѭˎ4MlW�N#*��+��"���%ZTjw�ˤ&��X�T�p�`�\'�Xm&j
��`G=�?D�;WY�+�]ʂ�y�Le�E�4�ίc"�i���l�jk���1}�Z��ҹOإ�}	��
�����f��|��Ԯ:�vXb2�j=�C7j����5����2Y��%�X��[.)���p�+�|�-f�Z�jG�f�U'K�Y"�:i�eԄ^|+*�w��>k�ɥ\K��-�m�kZ�`��	vY�ss�i�[)3�rq�^>�~�;s��(dy2�Y��lw\����)�{[_�;m�9��dEY�`OGT��+��=���|o�v�������Y<��E}���0��,��@����Qjr*��ɝ�͑�u��!�Xα��5��s����DG�x����y\����V����p�)�ʳ�,���E'�*A=,���Y��X�6-�FK�88\�<@+�Y%����R��'4͊��͕2B7� gJ��ZO=�Kgޱu=�)_�>���i�]d��q�
����E�Q󸉾�B[R)[�.ʔ����v{ї�B����/y*ꥦ;c4f�;fk3��d�t�<=��|�����o�8��UA8ko��/=,�i�jU-^*�I�ܶ��[)#�l
���Xkp�+vܵ�7{����_��Е�x�z���fs�R)��ɗ��)������p9�E���zJ�2��UΗ^�`蚎ԑiP<�{������v��Ԏ�4.�T�m������7�,y����ϲ}=ws�\GA�7Z�_G����"��W<%��o^|��f���2���ԹɊ����1^>��_4�ܑ��&������8ZD�7�C���Զ~��r�hm�L��L���$^�To����K�􊎈�B@[�ꄢ��mQ�Q
�S�nW�}�C�>=|��^B�[Nɻv=��S��}]�f��
�MNb���C��x�Xy��)6�2v�Q���ߘ�Rv�}v�V�>n��ۮ����9�i ��g�f��3ol؂����ȷ�ƫ=�|w.WUΟb�z�[n,�h�Wr�9�eS��yHb?��B{�Q�����y~�BOyY(}�*5��%�*�&/[�f��W��Y�ֽZ�k�^u�C1�POTMK��.��#܍�����M�Imo2��a�
�e�yY�nE/�M+�,��L����+/�9t7��(��·��B)�[�g��J`�u��2+c	U�K_Gؒ��\�^��h����hݧX\{8fr�r��H(#r�a�e5��B�sfF����������KM�r��2篇j���	iYr��6���Da�+|�+1<�5~�+/ym]�ѝ;�ɯ�x�v\��v�c�}^Ŵ/m*�C޾�dz�=��~??��Q�x��`�v37_:z�/3�L[�zI�ޜ8g璨��3(�������Yw#w�Tk��i1�9*D�'Y�F�t�����r4�`�=��Ҽ2r�rr{g��j�T7MM�Gd���+��^����{��Py���L�����q3��/�V�
>���'6c��s{1<4��YQw�u�z�R���w%|贡k�R-�Ȅ��c�j�J1Ee��
��B|r�s�^P)��'���D�{umւ�� V������B�`�!�Xb�:*=��f��5^��OU��vf�ML�2�����'X��/���qZ�J�:�Ű+$�^!�-��Q�o3���`D��
4�*�{;��B�n
�,.x*�nj�Q����7 HmxY��h^�l�w��w��5�}̅񑸖�[���z��1��,9�i����k�xLD~}���=�*�a��y�H����B-��7xV\/x�T�u����k��]r�=�l5�"��rn���i
�
=����8�S6en��i�d��3dx����~a��(����aU���溲���tb�w>F
�9}cu�}0�;nV׿���o{� +�;:��>���^�VD�5Y�c�+�6U�<IU)�ICUeJl���;��S%��(�}W!����lV�15��f3�@�]�JӼ��s�j̯U7)H2��=��'r�pc��x�q�H��Mm�+�ʁBj,�_�T��T�ӑ��T�\�W6u�e��-i�@#6׹	��Iv�Q25���V��O|�.9��9��.���]�q��,mEL��aBSE �Al�	m�׾Z�*��ʈ.�(J��/�
�o�|_�渫V��.�ɖB��Q�T�M{��ޕX�J�NVħ�Q���wB�d�:��}O*�^���r+���rTs=���h7[@��,(��˰TҌ
)�]Ͱ�mE�չ�&�5��8Ԯ��P��\�4'KF�!��@Zmn�K:;VbS�UJn�X�K�^��a~�Յ��,3�v.�{�J��%����B6dF�$SX��^lv�};����6̥�_X�b�z��5_:
"��_�G6�
ߛK���������-�Vp�Yc���;��2�L��N��C�%ykʅ?�`��5o�O
k�iB�{��������N���|�]�z�Mo�]OJ��}��WoU�i��y��ދ�,jƳZ����� ��쁆]f�q4e:=���u����8"9Oq1�vh�Eu��1��ɲi��z���"�Y]�fV��Sd0��x-�~��M����Ʈ�!�����J�8��	u���TV(�$�1�
�CYXDv����v�mᕊΎR�HQ�eYҚ���K2:���{��t��L�
�r~�	͐�7|εf��U�KOTN��Tax/���;��͋坏K���?#1�3g4���7��o7�,���묅��qKHI���
A纤B8�T�S�*3K���%���{�jm=��*�3��ߕW�]߹�1�pޘ)a��\�67~�`�`w���/C�ͭ9+K��>�S�A�:cBͫ[���k��e�B��G�R
#�[h�Ji*��?GTi5���a��[�nu��������O��M�Y�����p�g��D��Ӈ��K�8�+0�4�0|#��WY���Iuc����a�{u�\�p������5��6��Cmr�am:��<��OC��߁����Z��ю�	�x����q�0���/z�e\�r��6è)�W����z0�R;�$׀��DG[�o|�̥�'>^�5�KGПi���yԵ��{.��YW@ގ�Z��d��%�-�U�h�!�"�^��i�lI�a_�j���'������li�|M'[W����C�;�L.�{��p��p���P[�
<w<W�ϟ�����Z=�Wh${3�隃V�EOv�nR����s��K��i�b�-�2�M�������3{������<��ʚ�-�褙�1�	x�z8�[)W�Sc��������<��g�;9������6�]̶�"^��5>W9�m`����V�������^3�wA74��xG���B�֯ϝn�E�Gf u�m!�w?r'5P����5�q��s���&
i�Ƴ�ă���t�jfh�}�:I�7zYv�ټ�Z˄TR�����U�KP�
}(��q�����!��]����x�WR�0畮�>(��G��2>�#z`����m	�gc�՟G��^g6XI%M���=mw�^L�����(`��<�/�	y/��D�Ⱦ�B����7P�N�FK-_o���o~�4�y�E~���;�����J;�����,y�фHz�T�Q��]=s��63�L2gO�\1R�� O��Pv<O<��蟾3E����9�ߦ�&�ܴȄ.��)�3d`��顯�թ�D�L\L-/�^�c�h?(��]΁\��p�D�^$`*��"X�C���t.,3��,fzڗ�PZ�i{�[��en���E'hC��
�)9�|Ȕ�.�z��.S��.(��FO�v��/���Tױ�)�5U�R6�`Vߋ���M�4�y']Й�m�M���ywf-��0�����8,A˽�d8�a�@)dL�9�vk�u��maξ�1l8uv���y��^-�=�ӥC�	a�v^�X��즦���@x�xxz�r��J���O�CHw�>),��s��=�m,��X��4���-~+����[ƚV�c;l��7*4�p�^{�2d������_Ӑ*ܳ�5�;��J�[7"���#���^mfv�4Wr�,�7��5w�9�G��_)�^Cǲ�AἪ��� ���E5ϕ�U4��J�\>c���W�Rg�%�[?7��ށ2��_}����M�V*W��i��PЮ�6��V��Ǥׯ�\��(��~�+o��}�>wP�����
�P2�/���򂟢�.�NҞ^Oe?en)��VܔĦƲa2.��>��3�e���+˖)�/��׾1F��.�	�}�Q����[Ms�kgS��I�I��gi6�ҫ�,B���H���^��ޘT6U�,��JkW.�KoQ��WK��A�o�A�2���Q{fRu�tM�.t(�B�v1b�e��8eYۇCvv����a�)Mр֝�"���R��8˽r�L��/����Z�Z�$��
��kVg&c�g��]!/�LniJn�d�n㼤R�P2�@����C�� Rk�#��>�xj���2�����8��mN2{>;nj�b��;t�� P��Ǵ��BL}��9���a0���\�g����#C? �zy���P�:(�d(_h�3���p�3�
��3���['�s|5!�:�����Q���3n�����%����g��}��3������ԗ2���US��~�%�g�H�g�Y��+E0���;90ݬ-��Zl��b���=㞻��V�nq	Cu+4�zy:��qiFs��d�=`�e�Xea�P8Ũ�J��F_x�W���'k^Cr�|���#��z�8�n%&2��]OL��#��\�D�	�ie*'���g֨u�&�%Y���G�NCk���1Z��e�Il{&�F��RX솎�p�Ƈ+��}B�'/�6t�\Gɮ�tW)��d@�]�-��M�HV��P����x��X#uu���p�$A�z0�����w��i�\ߢ=c�֡q5��2�bv�����KV���N_"��j�����"}�I�`�	��r���pn="��/l���Ç��C�����5�k�n�zb�42	Fjw^�s�p��}4�]��im���_�}�,�po���
q��`&�J��F��ג��;P�*�ZW#�W�e��߰*s��=��80@{7w/�O������Eϰy���Z�y�e_�_�������G=��풬ػ	[
?�}���}�/����}$������p�n,HYn��m[�����3��LJ{7c�]�硃�U�X��>���x������d/*�$�ǆ���环cƦ'��{��}�5ˑ�^�9�s���:�Mon�p(���Dl��6ew����2/\�&�u���ڶ.�2�������n��Y�P�'�B��Ɍ�S�1r=�Ow��]hN�7�&����94�����gj����	q�T�f%�o)�C�z��N��n[��1)K��L'�׺N��Q�.��⠰��Pɲe�W:���U�2�'P"u��}{��ݢTȨ����^��<j�8u��Rq3iA�S� y��E7��ݺy8�f=����9tg=*k<�OZ�\�)�]�l��ڋ�n/��|�B�<�uq���I��;eX�I-r��,��CGff�n�2:��p}�S��r���h66��1�>���;���h���Ʊ
��ޣ�T�n=�KMc�q��V�D*�f��NR�-x8��g�sQ�<�v=B�p�S�Q!�t�p�I+�	���s�{��\��F���]��;�=�s|����*ö{�(��Q�բᙉnUKn�y�qW�e�&u�V1�pe
�n
�c8^����7�|�٭��j�ʂK�>�G�efEt�S1m2�/3]HЭ\n�)D��ʂma��vgrڿ�dU��}޴s?)�D��� ^����):-�8�ܱ���ipH͔y�dAt�Ȇv+͘�\�ȍ��)�9>嘎�e��ޒ�F֌t�%�sg*�� Z��&���w��,r�(�T�˚��3N�����Vq�����6������]��!�&ʾsKW�tnR��H�x��ya��`Ҫgm�S
�/`����X�Uѽ^�
(<�}��M�f�o\@��mo�����FlU��)��-��ٽ�1�zx�೷�|yw��=~��վ��^�r����\��:��F��Vf�6o2b��� ��i�o�h��d��iV�3�V��;C'&y�v�������
�q3���0L8ӭ��`Uhs��cp��"wMK|Ԇ�u7Ԣt5��\5�S����ЫfR��ۼ������7$�A&�]	^-ſACfN�d�è�w��0���b�9±�B�nηG�ch�I�2�l��"go�Ȇ;���)gyp��=r�4(�յ�/��ɹ\�U��d�b�c��ވ���h���<�8�#�ސrs��@��}p{���v�T�%&1��u����j9ݺ�;�����I*�!^�g�D�`������x�${��O>=�h+7,���/
��7�����.%tT�$�{}qU���~풛BM�8a�c�:h0�D!{N��X��4�Wn�W�#B��n,U}/�-C%��c���$,;Շ)dށv��tf�[ZS������`�r���(��M�w�R���TX�u���'pK��%�2�����
�^�{�x��9�����[��	S�}����Qv]e��$�̰~�@����qZ�鵎�-��5�����몶�=jb"*��tQ��q�Z�:��K��������km��-�l:�F#Q�����QI[m���l���9��5]�FZ������Z�4kDQm�� ѭ��۱T�n���h��GӣTRPE1��M4�g�m��\@����.��Wctt�M&��킒��kMM�uP�`��gI�m�ۂ�

"4(�
z.�"(��(�.���ƨ;h�:�W`���m���J������K���E5��nӦ�5�c1�
��Q�kQE4�Z5ў{b8�Z(�.�����,�m�Z(:��jƭZƩ�l��qDG�讻�I��j��8���=';ltn�;����Z��V�qU]X����h�N����ݻ]�Eŝ8�4WLX��v;�;-��>���2�?q?�ѳ6{�tk�|���e� ܍�o/��Y��<tcy���9��H{7�≞�nC�~��+5g��|)���;�2@���fg��h �T�Q�<���}~���������8�/��P�ԙ�+�)�gߋ���z��3)��
�d\橶�G�苩-�m�gy�s���KQy(^C�dڷ�B5"�ؤR�^z�<������J��(>��=Z���q������>���s�hg�o����0��R[ބh��_����0o�]��(��u�,�7]#��ɔ���+�Z�G6�R���K����&�_o�;V^#k���'�#�9���<yٓ���T7��s�zpEoFҕ�1^�1M�E���g2�b�$!C8�����ڎ[�o1t
��B��e��n���ׅ*��������=}q��y��5�sN8b64��WxR4��ϺY���*�sy>6;��~��KFW�W��I��xZy�C�.vr�T�\�Z��2V�3��N��A�U�)��CG�U��(���Mg��_	;���oq׽�&��9�`�>�6� l�,.zD5u�O�9֩�-���;_E�{�X�����f�>�] �]��( �m=y�^��
Q�HQ�K1��zY�#R��n�ː�E�1��%O������<Im����M�&ߦ.\܉]W��y�o���y˓�T�Mib:�R���5-m�v<^���E��&����EoT�SwZW	9�����ǝ�^:�&���@�Sx�W���t%�l�'dmND[\Ɖ��{�7���f�� ��{������6�ቛk�Zi���S1�Pmx�j$6�={�O���f��&pX��ݮ*i����R����;~�����l̵{7�;E�/��5[Hy�:z�}M8����~�ɐ������=@���:�5U[�X�^}޲���x�E��[�V{VS��lsm`�l����s���%w�}�R�RUH�1>�D��cx��ʑ�WyX�������V��.�Cm<U��e6�Q(�q�Ƥ;���r�9�(�G�H���j�[@�1'�Cn4F�8��7����V)�t�Noا��D��|l�W"�ސ_٪R��oB7V��|�T1���ڋ=kjr0��)ɞ���׿���B�d�m�s��v=�A�1��)�Ƌ��I���D[�
��q�>W�I೪���T����(�O��ī����u+�lF�7l�;�	��2���1�و{�'���tד:b��3Y�f~�r��O����֗]�bxԇkk�lc��8j�GIqXE]�9�}�Xfs篔�j�L��M%�'0C�F��}�q^@��P�9���J#/�U��R�
+j���9��D���nFlZ8>^�3��g��3��+�	����t�	z�fy�yK�Y:{e.4�hma�KrQsWa�e�uf{�wlc���ΛC�j��h�2CD��u��Mׂq�լ�V��>��]W�W( � P�@����w�!������˹��lvo�Dhf��}^�/<轊ؾz��(]�*�p����ޑs�lW\ps9K)׊��]�8D�⾌�Ĩ����Ȅ2�ȥ<����T�5ю�Е��9k���q#C�#A��Wv^�Ft���&��Hʮ�;w�V�)��u�]�4X'���n��Z�s[C�7>�g�ି7<jϥ2��2w��T4�y�å���1;|f�n"���ה��d��F��ˏ�5�Wf�/��|o��.��@~3jZ@F�z�Ec!>�ic���]&�pS����u�/ݘU����Q��ځ�b��%�R�sW]D��&by�gG����^9E��/tLTo)�B�C�n����^tO���S�{u)>�WɶeK�̕a�{T�k=����C��FQ��ѯ��]]�/ʲU��]^T��2y>�M���/�i�?\����{�:���EgB����~����`Tj��/�&�Q���w�=��f�{ԥ�Z������t��lbɏ:�����^�U!6�y�7n�E�?}}��vh�~���~�Nc����[��]�;Ѹ'D��C	�;:�%�.�a^���jH��'�-��(�@'��G^s�6!�d�9P�QM{ʣ�{�ZQ��6-rH&9*vڮ��xI˪>������D��<�9�\C��M��Z��_ǿ�����m�����1��4��)H�B.�����	'#�k}�s��m��_V�k'��f���8>D�%�5�ٙ#hr�2���b�whƸ���UB�Hq1�p{ЩL.���h�2|��	Se��fRu��s����flX��m^�_�CH�f��3�7��m�Ξ�,*/Q=�h9���<�/!��¸Ԧ)�-��"Z�\�;����^���\q��Ԃ入_+u�-�8���1�5H��+�	��	�Oʝ�[r1̘�#^et�Z�Rae��Kc�FJ�_b�SHQ,E��(��Ha1��k��)���6�v���x�^�#b�R���AzY����.(o
��~�À����	>��;Z��u��[�?�@LƧۨ���E�@����ܺ6)�r¦6faQ@Mn1$�S���-��X�I��[��L���y�,9abZ�ĲN�Q�i�8�&y��s=��zz�H16�sRL�]�gx�O�P�}�X&�GϾk�����*�dH�G&�,����Wቊң/}1P�8�qz.+� ���џ��
Y���c�����v�D�T�qSY%=�Cs��nʗ�y�̻	���S\�lA�F�m�ξW���x8|=�T�B��;�Y�[��i�Ձ��YX)aºW���)%{F�߯i���t�KSn�8������ك��r���81��f��t��3����]\ݛ|#r�Nkr�0�p��y��x#2���g����
Ġ�#@�
����>~~�������6�����86�(H� �� #6�
:Z䙺���o1Q^��p6os$���-p�pom¶�=-j����^�2���Ct��=7�IݨW��;���U��L���z�J��]��a�ˈ`ZPuV��q�ml(Bh ,�[RYB��ݹ"dWT���R�QӚ}�`답�r��,�ȶv������m_�_B�j%K'�,��������B���H��P"M��t��O�[�R�O��*��;�0j�����\)��o÷?{�c����@���ڰ�ӎch�ښ"~�~T����r�4F��l���s�l��<�����;vb�<���.G�����}&�ǌ�k�}����9=����d9aM!ޚ�>��"8�b��V-��O��SU��e�5��лȪI�RS�(�/ͩ������j�ecrS�c��+;'���h�,�;�VAk��n��5�q,�����z�0���7�9ys�]�����^ΊŧT���;.�B�
��d�=��!�x�"!6���[f��kkCW��s�ki��A�ӈ\�kj�pϬ�vb<5�#k�����4y�S�l�e���ΑR^�7�![}���οI����E���R�.Y��MÒ��P�\����`���~������'r���6n�vn]��k� ����@5���|ݏ^�Oh������ �F��F�R�Q�Z����������B�����C��C} ��K�:j��֟F�U���J�r�J��>�b�;�=iQ"L�CLʃø�#��8z�Z̀���P�*�4���D7s�{[uȵ���0���S�S���c�}�IY�çn>�ق�����>L�����b~��t[S�#K�=9&��;��v���ʻ������i�G�.�"�7=��m�E��e|�4�2��+$���"8�^\�b{}��<T ��t�/��{�˷ULռ P�
�H)��Ec��������Wu���n�b������NFsľ2�v��@�ژ3��(����$x���R�0�q��\��L\�za��c�O"��>���^���u׷&��X\��VT�x*6>��M�j���u��4�yЮj9����Ҕ�)>K4������3y沮��0�Z���p\�`�K�bkj�\�ӉO_\�����l���&o� o\|׏��
��D�y�,G��n:��f�������n��Wg��:�Wb�~�Z�S��c�N6��͇eu�y��w{��W���]�4�OOs;X�n����qgr�e̵�LmKէ���d{��䷓�r[�ܻLgɢ�_�q��T-"s��//����Ct)��l���p��^
��]��b�wW��]9=�KhR.W,;��\:�ۄ�9�V	h� 3�ϸ�tytո�S�v.���� ������Z7���7|
�a >���`u5G_<�ZruH�W6��������Uy�1�XUr�i�uJ}Q{,�9��ߝ#�{Ή`]d��K⨵�������T=�(u�r<uV����E�na|�T�����{��
d-�@�8X�8<dO�B0Vt�͗��3�N���l�R6�$�̽�#�� �B�I��a���k+1T(���N)�KOY�/@��iO|]&±e��;F^>��W�a4��;I��ua��^.�bT⏲3dzo��'k���Ko)r���l��XZ*SBz6}C��1����`F�CtK6�:��C+\D�;����qS���a45P��_vH���o:f1w/�X�A��D�^$^I"���nT���^mu���H���o����g��۽x��@�ޡ?-���J�e�n����8Ń0�c���C���)٫�o�|-�����K>͂t�|{���P�"� �Ϋ�7sq�V.�+�LE�U��dx8~9��/��N �c�(Os�m|<:!�V��h�Z��ĩ����,��M�V�(�$��zp�x6��jf�yg�p'*�>�<�b�X����o��YʽR�����)g)�QR����F#�<3;`���Y��ޣ�K8�%��ť�T��O`�	kU�JcD���9;Sh5v�U}������� ��*�ʶ�
Y��t��6�����&����uO�7����3�u�Y�H��r��e���oC��յ~��Vw�� ���%��'3�1O_��O�hD_\�*:޳�r���(eԢ3s�͵d�T�{�A�8��(��KhV�t�g��5 d�{$�4�|�kF�O�c��x��~���DsJmW.W�G=��Ư	�:ה�õ?X�U9�+}�*O��;ja��u1;�x��|�Hl����z����-�4{mV�k��E���O�T�c�^=��7c`cA}xQ7h4��(�BዒaU@��R�!h=�P4�d3H��J��fu~O)�?MHe#7��TuOdf����v��P�y��p�����=�~���)��nߛ��f�����Z�uM}���x�\��&*KA���HH���Ҁ���!>9?	����<��cr��w01���S�\�vd!K�g�ě�Z��&K%�o��+С��L���L$(�;9"���7��}�����ձ���Ĝ��5�TyE��0���+��]*�oݱz��|*)�d�r0j�4JK-fۈ��y�v����m��u'� �f�+�@X�f��GA�{�yy/�J�Nۿ�H��Uzm���ǫ{9���
Fs%jy��3u�S���z�����dɜ+����2ۮ�W>�X��3�FXY|�T֐�kD��B]l��ۑs�,��o�+{�������x3{����q<.�ҹ�3;�?�fs�E7LwQomPģ�Z���32��Lc9x�g��F����v��&�u�LMw@Q��G�>��sL�ОU�F�0��5��\�.n�m%���p�mݺ6_�t�D�d�G&�+T}jh�"�j�G�aP��:{w?P},�F��`��ȡswȴ�t�eų/q�-Nn[��a��Z_�P�<��{�V�_�2���Sݞ��Vf���7:��j=�'O��Hm�BF	�J�����L������RDIp(=!�[�TW�91����C"]:���3��K�Tn���������� G�_M$��DFCF����[�k�U��Γ���9x�^�ˇ��{W=u��vE]�6{W	MH-��P�{խ,Պ�!���"9�j]���2y:�%����U��2J�k�5����l@*�%�L��*���d%6�#��W�za�K�n�{�﫮SQ��%��+�ix���֕H���dWdO�4�܈�]�]=����]鉱�������P1&��Ew?SbG���^���8��?
Z[��q]���Dz�9��`��Ρ�r2�IL�I~U�w~��68�Fޣ1B�]e�z�c��sLQ+��B�[t)s̃�Μ��:]��Y�gJ�P�����C[GhS2��W��R�4�i���ͮ��m�ӂ0'r`,DԮ��lrV�.KZ9��]��V��� <^VgLa-OOw?�u�0���1;�4خ���5����j����ބl��D���XOV��ϳn�$c.:���ޔ\P�U���Oͩ������aT!��hg�g�U#@�k�9������Z��)�Y4��V�?W�[�C��zs���s�]���Y|�R5bI����͈ZUك+�L��Bg��C:a~��m�ɖ��%����%r��mGy(�屐������u�%�ͮ,�=�;Z0�O�b�`.�
>:�T\Yfσ������u?g��-{���k��7Ww���h���ن����p�6,��`(6�T}?	gj�-O(�0��;�e��5��f�b����5�4��i�u���"6���I3-3�[-�^s�!���Z���A�	�C���mi�� �P��3�|�K�FE�S6���8�W�!�L��4ͽ,ך}k�(e�=8�\�I�:��K�a�~�����mۃ��@�O�i�׌�B~hw�1��w.Q��Kld��;Ɓ�L��}g�G�wF,�!���NДټ��[N�i���z}ޯ_��UYv�L�m�ɳ�s|��_��f!�
�'I��\�c�(mnc{�PWru������]�f�Gw��^��C����Y9��KB^ЮRw#a1/��R����l�>��������D��Q��j�\d5.��P�}5��+#Қ��#:��v�r6�aƏVq�"�w�P̈.�f��}[�,���n�/5�L�&N�mX���(��5��)��B��tG;�K�5�� �
Sv�����tqYR�fGήОр<�w��h/?��ԼK�|9Nc-���K±V�<�fOs
Q�y�Ʒ!�qk�������4Eg�T�A�0eͼ�����[��wA~i��Zp헤^�w#��/n�cm{�U&m-f�����!��и���L���@	h���^z���89�E�&��/�)��m 3���:I\6��{p<U��Q��=�b��Q��T'��|�Er4��Z0�e�k�� ��ECݭYa��S��}����0H���oZ[wO~~`..�k�13Dl拠�Z=�ww����D�d����>��,	y�=���WM��͈�Ym�}l:*�r�\�݆�n��F������	��]a��|0?��y�MC�W�"i�sD��N��'�"�Ꞌ~�����-Oj�x%���'�P8�Լ[�Q�N�=Z:�h:�B��or�����_9w�5+��f��T��
hU���������@4F�o����ԨMJ([�i�j@�5��₷��f=튯q�5��Mx<���7�xge�;Y�'CFJ���܏T�Eu#׽��+j$�%&�C�-K�KK���Yos�j������=��o^Qݛ}�<�����fi+���R��Y�l���B08)_?��:��R�z�Co-Y/T"�wrnث��-0��p�=���즠K��,5�cy���������yl	M��]�pُ�qޙ&X�rG\L�%eۼ�Ꝁ��H{y�W�5�n� p�7L�D��Yp�k�IF����n�^�9���&�zN�ge;Eb�c`����͒AMi�r�]̺=`�[��$RQ�˕��}Ap���ʷ��ur��+Y�Ƿ�u'���սR�uG���5�gӓ6M(��J[չ�S�Q�Wa�A�+�H�uR�G4��M]��m�v���}W�`�"�E�{}�E|3���7©_N�!��<;(s#�EE/Be��QJ��s�)����Z�jc5�F���V�A-��wUa]�K�&����tLmॺ�uu!c)�Ǔ{JDE�:�k;d��u�+ɡeu�uo1�|g�X�xi�6A��JY�=�M2�s��*X��2�n�V��^ՠ��Rn�Q����Vޥ,���,�� d�<�{�oK�2]G���Md���9�
����1��]��]�Y��W�O4��3���=����)��|}=��O���b>�ш��i�D�Qgn����]]=q=���몙�mq�g[;Y�TkmX�X�5�QZ�N�(i��TDtj���2tU�:�b��n#m�h;`��Q�mu�ֆ���ѻv5�Pwc����:�Ӷ[k�k��u�ִj�C���1%�u�mg�T%Q��v�gE6�pPŧF�k��6tj�gQ�Uţc3g�����Dm`֊�k8��h���1��۹�YևN����4ŭ֊�&��F�5Z:8�h�+ckQ�荍�1ӭ�[:�:��ݍ���uc�J���fֶMT����<j��ŴkNq��V��]�Qu����[[l����Y�fJ�clE�j����SS�6�t=UDtmgX�"-��[�U�������{��c���Z^~ nDVr�n��
�Q"3Z^b�x��t�z� �a���ߖ��]�ȇ���� ���4�WSI�������Z4�~�N�'��h�]����uD�)�d�Rz77w�wO>��ىE�������R��Hj�G�z��P$�xL��E^^X<έ���M�̥}�c�^Ůl��M2n��l���]�V;�PaK�|�m`��Du;�Ҁ��MV2t,����Sк/�r�.�i�&)9N��Tq�I��7j�����H��/�3\��\E��V�[U0j�����M՛�D�F҄�5����/
R{E���[?~E];.y�1�?�w��?~�ŏ�n���+�#�sf>���W>xM�C(���*�`w�M)��T	z�Ŕ9l�|Yq�]d�w�I��������OźCf�L��V���P�NV���l������^�Q��Tu��M?So��������^�3�!z�W�w�����z_��E5{�ɗͱ9tӄ3j(J��LU-1+�����Kc���9J�$��n�as�G��8�����7�!]զ����%z'�yc*P�9*,6��y�=�>��q��;mx������,XxS�yi�L=��}������W���`�!���X/�d�}vf��f҉h�B�)S�0Nĩ�,\I��רsٛ�����d��vk72�$�&�R�!R�3L��g�\n�(�'4u�SaΓ0 ��bqVl�'�����{u��.&6�޺��� <��ڒ���>	�c4��Ng�čc~�h?R��jJ0|ޢ&�u��^�~�7;nb]u�v@>��T�X�G�H�V9��팠��S�EO��@솵`|��Lr2��Y+�F,�������g</^���P�f�3�k�݆����3�� J��MXR�\Nњ��-_������%zPv�s���">s1㜪��/+�'n1=b�~:�Qz�f5�P�65ѝd���`nzQ[�R�����j-B�u9)<4�k���	0��Ӑ&���I�YU��l:B���uH7a�Q�I@ݏ$���-����-�|�w��Qlah{�Ld���r���BU�m�ޅ�B� ��Ȥ��H��U�)�5��/�W���Y�|Dc-�����|�N��.p��:�jb�x�h�n�d]k�}��+��q�P�/h���'"7��N�dT��d,�/��.�B�(G��i�X��I�n�I�x��'
����I@�������oE�ީ�S�+HI�UC݅Jah=�P4��	���ڎ�ܸ�峛����9^�EYW\^Ib�s"���0�����t�͛��ٞ-�,�3% ��;��o[�}2�E�Eg<L�[3��ǳ��N�#7嚟��=OV�p9��ⷉTuj8ގ왬;'�Υ�12���&"!��]�Y�����
��Q�ؒ��e'��E�0���n5Q%����S�������{��厸s��,3�[ta�=�D-1Q|���A�X���3SyUϚ��;�����:wUs{(c�7#z:���煥[�R����9_CsW�-�����
���k٪ �2yu�<���J\P9j��Fwq��#��|U�b6	
%���O���MF�{����P��A؇\�-��+6�P:U�q�ѩ���q�F�밖c�D؍�N�6|������
��=�OS1���)�P�E�@����Keґ��Hٙ6TϪ,Ll���%d�'YR�j �GɃh�0��o���
ϲG�O�Ε�֨�75��ȗ�&-pMu���*�K�QǕ�B=�|���Γz����0����=����3ɀ\�Yi��_t8g�|��Vx��P�^��Y�)t�l���lT�q�S�T��Uw�o7�SgR�|�M��c�0��BwA�|	IS�k��P�j�Hn�4�crt�fyU6Z����'y�uC��`!5��s��guScc�~Jm�BD�{Uc�yF��[!x�8'�ؾ�MK��֌���+��,���z�}�ٞ#|��Jc�B��5"u���ɫ2�p��R�씶`9���n沗(&kX����^�����c�Ӄ2�V��=XV)��;04�2Ӟ��0a�2��mV��I�x�l]�/� ֳ�-���UUh����ng��9����P�<�.L��["�Զ��K����^+(V=�בQ"񈕧޸���j�r�V�9<��	Q&L�U�mBg�0
i��۝*�����Y4�ZC�{~�]y)�K�uT�R��(s�I���E�M��`�x1�������XCG�[��Ė,e���Z�>J�S�׎y�əc���m�fM���E�@�^C���*,^�+��ǵM��n��uF�n+��x��2K�1)�T���J��fF�Ơ��YP��c��l��̻s]o'��p��dǕ6����y:M"�ÚTS∢���QʹT�~k���?@��p�5<M�l\�W>�b��w��t�Yz���)��],�en�@���W�PK���Gs����aW�`_dV�",�_�~�U����P�&����wM�B�['ת�[^��@�1A(��Q�E\;�Њ�ͮ��vZ���(e�P�Gmo��łsR<�~�T���8}"{��N��O�=�o	�*�-jݲ'"�GY�p���w�4g��P�N��زsXB��Vb�S�)�d���z
��Z\��3Z5�E�@J��ˠ�S���{ؐ��i��61N�Qx�G���^ު�^���4˱{N-w���{2��4�!����t�\b쩁�^T��1�*�ΚU�.���S�j���Xj��j�gN�E�]��6��j�w��� 1�!��Y���.~������Lק�Գ�5x�ms D3ly�!�	�M�75���,UU�߉oc�����C�����s#�|cS�{�dP����uH(�m��2j,M���z��V�<0k���WY��5���3��ހu�7����X�"�[3���iY�Ә�`^=0ޒQ|
�LĘE��w8�pl��;7n�5�&Y�@JHe^�,eS���s�ִns���1�r�'�͘^\-JW�kʘ���U�롹5�:�)�U�,�7x�zɋ2�Kޮ>r��9�8~���E?��-7|a3������P�b��l|]^l�^J��EE&V��=5V�h�v]N�S$1k��r;�d绮l�ݑI3�c��}}�7����A���}~��Nf��Z���B�+�utī{�'%�.�No�l�T�=�*rZ�lo�Շ�FՆȄE�E�W~�<�#�Ha}m��kVC#�*q}*V��TZrpj�z�m�����G�Ν׷F|�}�'j�%��˽@�
k�����W#�	��e}��:N��όj�EP%� ��xd�1ǋnagf���sg��
����_��1�c��{}�'�ZG6��ON;���C�)R6^/Et����44:DiW�TcV)��<K(�u���஥
I�/�.g�9�9�� 
�WsN��r��F=��,�Y�;�fe�Q�Рbw+^"?�=}�a�u�WO�Lԇl���|�6�\v/ZJ��>��r�g:60ܢ�E'�2|�^�)�[���z��C��f�xkC@�mu��Vb�Q�7�1G��Io+�r��Wk�/ETGd*�zcWwli�:�����
�c����,�����j46�Ê�t�X��O�\ A4�et�L5lsju������E}6�tH��L�c8 M$���_z�Yyd%�%�ϗ=��X&q8Ԍ�m�b4����Q��50�� CDWp�G��u�|3Jp�3�i����,�{yN����5s8�i�wJf��`j'��_!�5��=�<���x��Pe�~�?@Zw���;�}?<ش�~S	����/NNdA�>��]-��k�L�Wz(�V�V)�r��b�լC<Q�;忻�~�7]���|w޼���W5��j9�$��k�!� ��g�f��?�Th��yfE��R�%�[�()�Q�ׁ#QG�!�U/B� ��O��CL��*m@�$���&�����q��.
���7�~}�	�����e¬�.��)�#א�����2��D���Q���N@uMʷ]χZ��1�'�xع��y<�d�O�i�=m�+l�f�MJ��� ��WZO{P�/d�7#�f�B���+sF��S�B;�s"t��UUU��7��?��J�\��*�m��B��0�(u�&��u3WoE��Q�ծ�wy2�!�<��׷j�rl,b�gZ����j�l�+*u���M�`a2/kb���н��u���dE�fe����%s#u#�֢��'	tc�S8�ŗ�+��&�[��_q)�$�"����;*OcK�ۉC)�,�
�ƥڣiO�����*R!h=�P42�4�)E�c+3:'�����{���3]w�n��	�s�y)��Vrƙ���nk�b`���5��ar_V����Wx�쩽��A�%I�r�LS⊔˳�Qn��B�煥 *s�Str~������uA������׀�j�<�]g\��v�Bv�ӄxGvΞ��<!����ͭE0��}�����]u̝�3Y�ě�g��r�&as�qm��hU�U)q�=����,��~	N��d�<�[��6���+aX��|ؠ�\A'Vb�C�[�%��=�[��VP��S�q^9�"�4<?�����3�>�E�����XH9֘6�k
M�"@vk=Q'��ѝ8dk����K�Q��5�e�.�yk��N�S8�8�Q_�nͭ*8|��x��{'g��^HYt�ص��\2���r�՝GS�{#��:r�0��[���w7ҵ�u��n���W�M�/h�ejޮ�V�J�;��)��f�j�r���������p[Y'������ކ�yy���c���y�P�v�.��2=�P��i��@�ݺ���D_ޢ����]g��#��\���a��{6�P�âU8�iQ�Ɠ ozx��R��Z���DL�����z���m��hu4�ܡ��7aK�0S�vN�f�BE��Sl�+��5k��6�+Bг*v��]K�>�!�V11�Em��g�]̘4-q֠w=����zo��
>���%��#df��s0��9��� ��h�Ρ[�`�`��7���Z�)��H-�E����7Y�?���]m������#��'&��+�7?|��;͹����(���<��6��(�9�R����ƭ��$�B��=�~�v���u	��ʒ�RUJRz��]��1��{�F��\8���֪�;�m�Ny�*d��*����/��窦����M��T>�)Qb�˶P�	�;f�.�l]��ǫ+[�_��*Ȯ�U��T��t�M݉U�זI�������e�-��-<��&���U�ز�*��u�^�(��������ܟ�$+kP����$�t�c�F�1���u��\�rr��f�hkk	Ñm͝.8m�൰V�"�0�+qə���r��ʽo$�O����Ư_T�oF�
���q�۠�쇛���w�2�S�%v�ru]vgr;1�3dli�A������s1�wj����3ǮDDs�P����ȖR;)\����qW����$�Τw=����q�v�&�0�̋����$�8ňv!�!<"o������i�$�_t��9ZΞ��Q+m&�YN�Tk>�>���Z%�uY ���sO����Kκj��������ʼ� ��b%�gia�ԡ3䫯;Vtζ[%�׌08u!fVl-v��Z�{dFTE�όdGm�z�2Q�Q�F��+3�ϳ�mc���v`��@���n
c��"�j�����fyn*c�
}�i]#	��\��E�>~��a���,E��`�J�7dF�O�)]�S�q;�]�`G�0�!]�iS�+<c3jQ���\D�)�p�F&ޘ�;��R�/.��k�(K���$Ċg�˓��cݟsvn�KWw�y����i��g��g���Ɏ$3�����J� x�o���R����f���O~�yy>�)�LD���v��]��S����.����5��GZ�߱J^�-U(I4����T�����Y4����1�0����w�S���A@x��nl��ᦔް_!G�ξ7��}�â1��%��n�^-�t�Z�=���n��V�^�?pm��̹+�q��,��w�' ��Q�Ke���Ч�U%&ͭ]�P���2!�4��:ܥW�
�D�٤� s�_%/?D��S����>���l<v�r~�F%k��2jdK�Et�����z$����h}�d��:·��{w3�|���D۸U�K���gdu���wE'E�"fӬ��$�����!����6�=�4�lvs��x�۾����m���;�
��\_�ʥ�yE��P�j�c*�L����m4�Z[���d�y��W��8�������f���r��%%���,���2໚A���4#՝�ŝ��P�t	ܠ�gҏ� c��6�'ا�Z�g�_�B0.��GpN��f@b��tMՕnuۗ���'�v?<.�H����}bI�dY���k+1P��l\��B�0ұ�O�Cw���[|��v�6a��t2���=�OW����*�t�7�-s� >|_/6�!��4�#6���ZT�ޘ{�����d�~%Ra�c��:͏E,3Xgm�+������엹��q��ZSpL앥U-3us�JuEFf�m�܅x��2�1��U\��`gO�:㝟X������- �ߒ'̯bFdq�q�d{r�����a�e;�&K�f~��|�߽���%g��S��y��z>L{RY�B���\����\hbw={J�b��׹�f]�A%�pc/��vzƧ�:K��HC��^~âa[+���&��W�-��^@>Ktu:Z��L�'e)}�*ΨX���o��z}-�w�w���u��kL���\�%<���R;����ˠ�4hk���UbW.��4�飈9OV�*Ǧ���ybtvw���f����c�g�/c���o�\�cJ�|z���Ρ��j��	���Z�|Y�nU����2��Q7γ�Q��0=作���ó�1�� �Ӭ���gc��k3�������U�7D$tk��$���V"�S�xr��Y��..gq�y�],Ý�փ�����Wީ��D^�w��u���[��9��f��0�|k;� ��<�G�3���]�S�����œӍ�n�@'t��6>WL��s�+�4�&���>��{%!��*mS4�/�����kI���5����l'�n�F���!�*=k��q�od�\�jh�,l୲��/�jP=���(ij��*�%�=��6(���g�S/!�UY�����+#e+�*�w�o]��10a�vu!њ�-oK4]\���ז��>T�qeTx6d�\�)"Z����9b���R�Kx�Я���|��+���R͍̦�_k��[�D\�-V�I�k�f��-���r�R��|���i?a���݂����J�8Cv��ݐy�f��1D�o�Ý�Y�]7`c+�w8���_u��Ɇ:���:iR���ۻ�D a ��J�c�Ѹ�"�����׀�E�Q�X6<���Psqͦ����`��ч�4�����j�/t/����t�~R�f���{I|�ٖ///��3���A��qhZ
��3���v�{����}D^���t����I����}ݡ�M��y{z0\ZV�g�!][}K7,pJ�*OL�4�q@ʹ��a(Z��=�����%h���b{kƄyp#�[{��]��(i��hRȷn��ӻ8�o6#�A�k����	���H�\��dŽ��8IS�ӈa�ʌ#�m�]&0a{��$01�����sLd��*�
�|
�Yٺ�D���a����y-���8����u.:�8)h@zb5��w�ԩ�,�:HX5�#X���+��9�O�A5z�b�R�ST��.ݕ�:�cB�h�7��S�5x��J6�)�	!Ư��嚛g���v���=`WW0unD���x	�w&i��Q6���K'o�.�<��}i�3��(}���&�:U���!ᆥ��a�]�9�a�r����٤W<j�TkL1���^�M i�|�9���%�4�������#	�:�0�KJ-x&��q5��(����_ᝑ�%	xu��yL�hɆ�6`
��h.{WW�:&s�憰+%ft�n�$���F<��3���йJ�no�,(��Fc�б�V�$�y	��eW7w��x�8�3�w�識}G���7ᛧ ʷV.����뽦���F��nűEU�S�\T�]��Z:;�vնј�C�ٻbѶ1�z7X�Ӌ`�6�vk���V��[gF"�[cSMIn�II�lѫZ��3�"*N��cU�QD��x�����cwb����UR�kkF�ql��5i�Z�M�����֊&5�ki�5��u��mU1�n�NvLMWm�U�v�kA[�3TV��q�j���Uu�1M����(��C�ƣwqf+bۭ'E�A�h�c]�ƻF#h��v긭X��U[j�D�#bgGOb����D[b��c����:��q�ٶ���ڍwq؍w��&�۷[v:{lΫ:����Q����#lE�4F�j�j��v
���w����]����b�uG(֨�QE5�[]�6�*���5D�-Z��gQ���Ul��c��Q�61���h����������<`F��z�KX��m'+�/z%xa��x������2n�{�Ug��-�W�U������W��2� �����?%�!b�ҽ(WT=�/>�y���cߜ�r�,�����y��kq~P^E:L�Un�����|Y;�*��_!S~�q�4��ӛ��4c�尤t��w>��(���"��8�Q�۞��"٧���g�f��8��D�k�{2.�$�rt�ھd6��e1��޷c�⛖��j7�ܽ�A�:������褔��L�%Ki��㮝�C��P�3Li�8X��3�/�f'�2�F��Z�����B�K�/�Ȝ�9V0���O���f�.��=�Օ'"��j!��~���D��)��Y�W9��i�w[�Y���uu[Ý9̮+**z!﷪Y�h�I~?;�ƯK��$�f��W�[l�-o
S$o�A� ��u�b�p��O���ԧ쪩썯\�|�L��U0���T��������!��(�c����{G��%��IՄ�Mǡm)��Vr����"�a�)@7F>k�b�!h9�r6�ak|�U#�C�.��1��Cȥ��3	���9���1<"��y��4L[�H8@oD��{Qɚ��5�7ጀ�n 6�V���,dԯ��2?>���"�1���]w5"ѯV��ݠ�)yy�B�.\��u(�������b�����u/f�Ԛ������k�%�e�X3�d�Ob�;��g�V����)��M����x��N:�?����
�m��O�\��+�������J^>�R�a�,�7\v�}nmvt�9Im�勞L�5�`�O|a��5��/��t�6.�T���[��dw8�Jt�&��q��6�w3z�(9{t��W`��H'A�R�[?K��\��ww�J\Z�}i<���hE�f�i�D\O�K������F�l&��̀�|D0���;b3�
�"�w�"��DO-���J_^�ñ�����H3g����	�Q�F��v��:� �|`���R�A��q��������'6(�C����`+u_ozx��R��ZԾ�[��>R�=N:j��=���_D �j+Wb8�����q�%�˔�Ì���M�iFm�=�}u9}ڥl�{�!<~�����u��j���n/ٱ�p��r��_[��(7Y�t5M$Y�s�}6�}YE��s����^a��<���G?VYӇ�Je�����HM�n��AW��iܬկ�?:r~
�����*����sӾ4�{kf��:����P���jޕX�	]���V�a�ާ��lM95��<O�5��������,N��@cz�bޚ
ۉ�Y�2F��6��`�!S�t�k�-����2f���AV^��ũ9�����%Z��U�B"��wq��)0<Ǖ�Q-�0�/\�>����?�fxVd�a"�ne^����SLz�V���̱v�+Q�Iv)�*�)=J~��UH�Ɔ��t66藅<��Hr�ښ,,tAe�⪘�9�R}�ַkXP����!��R��}�]P�����T��jք8#z�'A��;�;�_���酀UJn�E^7_l�ss�Aq:�e%�FM�E��]ȵ����Z������vi�-�.(�\�����#T�m�+�����[4"4�k�ʣgY���S1�m�)���oU�1�Y4��et���b�W\��A/�m�csC��|�tTF�~2燼�n�+V��B�����x�"!6��ʦ���5Y�[��IU�ݾ�j���q��z{m�Zz��j�&�Bb�k2��5H���(6VY*+�b/�<�
5�2{.��S!�N��K���?#;�hf��vF�HY�!�JO,^�Q�71y3E_:��L�yw)��0�7:� n��EN��v�ϬR��3k�!�f�#��R�'0�L\d�]sWt���Z���[#:(�cYeѥ�##��OA�Xga�X�諰_��6O�����2�ާ�ռIP�x�4��O��"Q�3M\�b^8!�k&C��%L�Lĳ!53�=wad���r쵍)���x�/�i���y���}���펍��r*�eȅ -ܣ)%��r�&�����	�D����zr�]�DV_�*�:��'�c�ᚘ4��F�i�B���Rѭ��"�}��l3�8-�D3UE��:��nU�Nıuޤ�K�e�d�}E{�1�k�S�~�����&/���G���)��S�&��oD���GR�,��OzF����~i�#
���j��ɺq�4⍍�ƳU��,
����1|��J��D����(��~M�)Kڥ��o@�����oR��YG*�1S�Y���gE\���f��k�Ť+�nl�ڦҲN����Γ����K��C��=���>��{OR2O��5�N���&�h.��o�&):/�����"�8(�z���� r]2���cU�r���{N�C�Z�w��:e�k�g�W0��)8��U-|�Qi��"���߉×M�W3Q�Ӻv"�����R��wTJ�y����y\K�_�9����Qf.P1��"�WEUչ���2��z� m��ꑝ��n����L�8h&x߱4z6}U�μ����Sgo3�ɭ2����O��~1f��k�}�1�&U�f>�n��,������ʏ~ψ��vC����!��r��(��&6�rXo��'f�ڲ2��}����ʖ����S���%������0>T��q)-Y��צ�j�����K�����>B�^MGkf��<��^�Yw�Y��=D�I�jN�E�Br�m;R�@y���]�ch����SW�t�z9r�K�FN:���BU6�"nv��t�^+w�L1�箵���(���*qFFt��J��ml�Bz���t	��:�l�����Q(�)�D�޼0��<a�P|ά2FV�S�e��5lW!t{�F1�#!�B��v3�z��-��=���p�=S�+��A�����+y#_G���l�N������N��k���j��u=��k	a(l��Ϛ���.^�<��(^�E�~�0���K`
˟��^�ͯ�D���O�2�ܡ�Q�އ)f�`oz8���ai^�	��
��DET�rw����O+Ok������Bf��Z��������'�B-�@*�����F?���|��<�界Ǔ�}u�����"�ap�>C�~�ˑך���u�y�79� �o��Q�I�-R۟_8���c�m�Ǐ���H����b���^]c�^���K�/)�+�'G*�$��\u��fi{�׵��ܨ��}���]�U�}-p�ν䦝���㏏�_��<��۷���2zL�J�H�٘D��u�ɫ��6� �s�zT���n��s���1q��m\��5��;c�kqU�H��鶭]^k\�/.�+��"�R�ζ`M�%Y�m\�1ƕoJ�4�U{��#�� �c�e��Pa)�����؃7�4N;�֝Ĥ���;���<[�T�9u�ܰ_�׾.�;���Ǻ,�y3��/+�c?k�|A�Ū�<��p>���/b�x�噔7��K�>�qM>|�K�Թ	��^�rz�M_u��^(�ʴ��'c���)�?`J}����1^o>ņ��7F>k�b�c��3&2�Z�eL�]'��z(>L8�&�u�{+a�oGR��iG��y>f^
�5K���Ǎ�3П�L1�5Qx���*��hˊ9j��F"����P�*͢��מi������*�;Q]�B���Ar�q��_q�Xt�T��ޞ/K#��_R��f�0�h��v^D�q�<�,$҅a�W��|�%����[�ڒ�#�Q�ul�*��m�](��}N_o</��n�+T��A[;L,�
�"V}�p{�VUz�3�ͻ��B7�u�d5E^ڟ��E��-+|!?��0M���k����UV��6�Y����OE\��:��*#���z�z�ed�L{J��X�`ozx��Rꬉ)��o�_ ���m�U���z�U��©�V�l��O9���psgf��J���w���z��{.pX5y�4�i�ݾ�6������Mc�4薱5:�f��z\�pK��� ���<̷�:�9%`<���y��M��M�A�ʝ�����ִ��t��v��٪~����~�+A�&\��ʗ�	���ۨA���H�8Uc�sl��d�xd��N��FK��b��թ3�6�Wk�K���[��/2e�3�zq����H��T�e��-QM=6�2v�O7ɛ&�z���d.�{
u�����(iڙ���*���aBS@��-��	tD=$�_��~�{�;��>}����mma�H��'���R+&�Y9Ԯ������x��f/���m��8uĞ���Xު��]BjǕ%ا��RI�|S�O>ƫnJ�K�wTX��m�d$s��GWLJa@2��%Tȹ��m����A�W��S@t��%D�]K�y���,��}���G���^�����`fܶ������E5�e��fv��/�u��]�Ot%z�Ah��4-94v���.ʒ���/�z��d��$�>��أ�2"�%a��ť�������+~�f�M�I����}���:Ur}���=_`��yQ���Wo���rc�Ek�V�V��,��B�B�� 8����S-�/U���X�g�T'���ހ�Y6��50!�[��`+�-u}��O=Uf �h�*�"T2�^�;.f�y:b���{ކP3�P�K����
��5��ջ��ʚ*n�[e�mv��zN�t���ޚ��+7�Sȟ��۩�8W6�	{g~S�����c�H�&�綺�G�!���W>s���ӽ�����3��l�P�d/� (���R!F..8Fx�r��3p�ߘ]����ies�X��*u���y���T(݈� f��wQ�lY9�-옷��)N���+=^aa>vPz��k��Ǒ�UCv>�+kt��ٻ0RӋ⍭��F� ������L8M��5��$@�Z�
��wz2F@�{"�b&�.�]A
S6��L[�L_
f����y�T�@(�r!������u>7^��"kb���͹O�ji]�5C��e���ש����a����9œ��(c�g������{s_���pq���Q��sZX�B�o/,[����_�����H�}%��0�v)J�Bb-BYF�	�-9��7����_��]X�)��d��*k��,�(%�]+�k�[dS�T)pd��s>�Եh���J�$�u��W��P�K�#��f�X�e�,̠ɬ�M�\�v�������xi�GV�`��R��ߴҋ���e�DOt;e��ml���8�LRt_E'7�D���K�=V*k��Q��ԓ;+ւ�54@�����z�W5�Ϧ�u��F��ϗ�֦AΓ4;�h���hv���?^��Q�=۶G7�ny`�@����9[��5۽0�w��Ѯg}�w��!M��,֗n�M�
��ܧR&&��:4�͌��-A@P�3���v&�������yY0[��F���Ǩ��6
���*N��(���lD>p���b��-��Q�ewM�-�P���eP)���} =g��a39Qϳ�4�:�y��w�n�i��Tn��΅�f��hR�PR���W�����F84%>�"��<��ۛ���i�O��O�3v@�0��W+��/�O:c[)#���ȳ+���D��m�Z�U[
�i�z��Ve���S�w�LNQ�VC�Z�>���񞻓����"�NX���S��k��Z�:�4�s�+p.e *̋����ֶ؆R6,I6�k�(�2Gm�������C�|��ٻ�Ǩ�Y�r�8�=s˳-Tm���voCLL8�m��2���4s?���f�夹��6W��cy�@���f}��7��C;~���g�������8Eu��YF�a'��z�%�RC�����$_�i����ӯVB�����E㼞�әsl�d����<I�Ұ�^;�5����Z���J/�.�J۬E/{�J���ܕ�o�;��}��0O-���r?�d_�6�F��;���VwD��>�Mˮ�-9�MąԵ��R�i��*�x>8�=�x��G��̓[�d�\]=�O.�jx��!t�7f;��pI�$YT����mR��%�\e����瞋n�>�����i��15��$d�iSt5c3풵o���t�����)�Rr�O�3j�g�j'O%��J粁㵵SU�q1:gI;澙���:-�]�e\�5��M�t��WC��j��&�Z�n�7��m�q6��O%��m1���!���fBC$Y���d�4�n/)�^Wz|���g�إ3������^t��-�һ:o�'ηM��5/�٤�SW����7�+v�	Z���3Ms�s!����v(/�ޚ���`��sU.�
�H�=e���*�H�	�-����#j�����p�[h}gA�7~�۷rK���t����l������^�Z��w%`9�y���n2'r��*d#9�%=x��oQ�=��T	J2�Y��y{@�g����̷3k�p����v2ˡx��S�Tݸޱ��``r:2ӟ{YQ��;��ZLFZ޽#"=�
V%2�R�@oHœ 9��Tjm.�׆����9�)R<�c��|�z��JZ� �8����n���t�2c]�M�~�����+���%o����P����ŖƩ��\�*I�]�(�S���!��Y��5�eG�� ��{�3�_xP�ކ��<�^�:�}ku���}�0������0`Ī��"�p;��Z/yjR�&��\@�xgRZ�q,�pԓ�μ��^�yQ�Y`�k��n��D����jv�99�%
=�%Ӳ�1��|�ÎN��^��U얂z1a���H.6X���^�j����e��2m�U�?M���'�!�h{�C���`�٥;��'^ǽ�8�80�����)9�V䅃��.����9��SNV�9��^cՂ�f���2����#����('d9��Hir��ǯ`�]W�"�r."��u�`|���Q���3�w~�E��x�G���>�8�j櫍Yͥ�)ۥAA���KC�n�{��M���ȡ�7ϒhC��gD�ۣh�t���k�jk����<3DG���%��t�����A��ua��J�=��J�l�������W1�XZ.�)oM9}��S���7{.�o3 ��M���%B�u.���f͝��gw��b'.��6_�ɢ)y���y� 
`}�ʈ^u�[f�`���Gr���W��^��Q޾&\��8}�wgc��ѣ�`GY���#����C�����b89�J��WE;4����b��3v����ʾ.��
����MX�#/�o���+V����]��`~���Ka���8��	��x�1b&�G���T^���#q���(K�է=�o�Jy�90}��3��5�{��h���z�ęqT�a�3["5��2�79��r�S^�oxAxR
T�^o������g�S�vu��Ý�E�.'j��R��v���ʰM�� �l�=���b�}��$#���V�\�k�ʺ�����8�قbW��n�!��v�(�O`����m���� B��ٵ�X������c���m��*��%K�<w3Zx趄�Ч�y-4���+!��H+T�P��/r��#.���T��9�G�e��T ���}����E�^�b;���v��Kr	L�>Al�ڭ}���FF�{�V��8���e>�U����Jnr���FV -��I���X�6�m7i���
|Z��(��A�&»tS	�L��0g��D�DD�=����w7��o���;��|���}��g`����T� 4n�=Wb.YX�ޘ��Co�ފ]\��.M��$���zh_/r�-uzk�\�����r)�o�ϴ	�;���9J�������μ�RY�j�Zx��n��n՗7��H��v=�~E�
go�~�x�H5�\VV$�����-���Uث��n�g�\TTPP]bN6+clj�눵X�;j"'Uݓ[�jN�p�cUj�k�榞ӻ�Gvn�����]a��N�U���m=v��դ뫶��6�u��ӣv�.�-���Gg6��9�
4m�S��(�Ѫ.-�S��5��UMUkLb�;T�%$D35���=����Df(v1��UE��[�**�ݻI5$�QPQ�luݵ[�n��ŤƬb뺍����Z�Z"����'h��Ӎ�Eu�f�VV��T��P�S]�wt4QӪ"I;b�""f)Ө�X���B#F�)�F;�i�DœS�h�$��:rEի$��Ѻ�5S��kZ(����j*�j��m���{�4Uk6�IF�Q�:뺤��\�Vي�QF�ѵf�*��2����x�6	4�^�JF(����#�����Ӆ��9�e�6C�I/{��e-s�<��+(�o��.��V��x�(�s���W�?^\^Cw�1���c:��.z�g2��nrw��u����O���'�u�h���o�W1�ق�O�5Mp��{�#_�Փrcw)���$�7�����Y��j���M2�s���;�������;s�;#��`���K�e=���-w�;��ѷ��+|�4o4���ǻf�\�f��ILi��B�4�ew4Q37��K�0٬�A���Ħ&������1���H��h8�v����3v�2;I����I���Ǡ}�k�����<�ՓgG(��W�ș6ލ��Rݯz%�:R�r�6���xx�^��K�SZ*�8���I�[Ӭ���QWݤ���Y(��Ve݀�Y�^2�v:�pky|1�q�^���R��ۢ"r��>TaT,\1VI��AҼz��@�.�Q�ߒ�'K��R�f�h\g�<d�My37,xĈ��p�UF.�O��t*��J��DMaVЊ��1��J�#~yx���K�Q{��V��O+J.�;�f�1��^��쨮h��8B'�h*��3���u;�%�T�X�|��X�)Rv����1�a.T�y����g%QT��J�U�nN��!��G{4�ru�)�WA��Km5<�r�p�@����q�^{r��]I\��euW��������=ҙ��?8��pޛ��Ng݄ó\ry�j�hi2��A�s�Y:K�;a��W����%X^�5z�^P�w$��8�f�;%V�9ͽɒx������?,eڱ���_�sC�9R�W�m#;����a��:���09U�o�yFP��z���jc���;����W<�'�әګmfݺ%ϲ��}�-��A;��zEg�=��M2�[;c�^8y��\��a���..ي�1D3�b�l���QrF�E��ĺ�ʇW�Mc�b�� �f��������Эc�K/h�6��hA�>���dj�Cj�E��:�6�d5���ܟ�=U���2�L��j�^j^H��ȋ���O�ky%z��ߚX�J)W�ٓ[�J�6A�V��z��w��h�k{��A�m_T��9�5Z��t�H`��f�^Sr�{���/�'���f+�ٻ�.�T��
�Ѓb���ŮQ��P�#�1�=y��4nޑ>�L����<�����'�L���O�K��2t����9vJ.���Ӗ4r�#bnu�b�d5^`Ȣ�t��J��[-m�G�Z̏<ݽO�#Y��d�-�w�y�!�R��o@��T3�a�(*��v��Ĕf>SWG1�j��"��\�v���M<�m�m\��Z�y��	�������������"Z�-!��nj �W�"񶥖�k�)�}|mi�����ˉ��7�V��i���y�����&�����e���P�r�܈���u��A����mt]Y5�k��u���-�� ^V���l�f��f��n��|.�l=���d�?x��O�c�e`�:�E�ϴ�h7�7����sm�զp��д���$�/pq�a�Qb: �����Sۄ�z�ZIrߔB�'ی��
��UP&�;9kD���a��"$����5܊���^�V�g��kZc��h�\��Lʞ�$H3�8|�>WYmJ�٧�\�����$lڇ'��ۣ�).����Y��Q/U������y����̙b�����8q�;��'�[h��5�^����G5޾û+��q���n����G1�df�s,΂�93�d�j�p�0(ߠ�sX*6	�*��X����6����7�m��i93�;{ܣ�1ۋ@��fE�9ߤ���ay�{ew�U�~B��'=o�ڻVO�і4�l2��x���!F�k�tn����L��6ITvv!����F�t��.�f���}�f�T�3�-����k�uqrc)�a(��@�6�z�g(w�H��i "����֦t��4n4\C�X��9S_�V�ۀDڪ�Z�q��@�<3J��l��m��ډmo�Y�#�������I��}�s}-sU�j[~�ϕ�vT5ęثj�p����1��6o����#��g��3�6��~[ڡ�����	�x�j�s���^3*�e/%':�ε�}T,u#5��,�卲-l�!���2����ܴs��Hu�~׉b� �[ɫ�O~��u/�EH
��^E�9���䙳 b����!Y� A�%�Iז��o9�M�Zw@����G��
�^�y��6	���.��q�|��>�g>�IR�@�9�:��B]�[�]��+%�}4j���N���$��yȸE�>��l���teo.MRz���Vd������*���ڽg��0�@":��X	Ri�$���J�Vsh�y�l�]ӺOw,*�y�殆�u��`J����.�6�*�H�	�-���FԄ	wg� Me�!>nS�!�r]ؙ`v�>�޴�`�螺Z�'��Ta�۲*Nn��v;oI���p��7oH��wJ|s�{;����dc�5e�{7����"�E ��J�i�5n���������2&V�n^��j�|��ڼ��Yq�)�a�N�]-i��7>�X�Vm�me������W^��Jokd���su�]n��Gn�F�&�ė��2�A�t��Yi����=�[d_�2�P�UD@8��/�ռ�u���4�{�jC�.ȆI�N�=w`�ё�M�|ly�^!b4&�)X7U�<�_@e`��$nsM'��mk�TZe��$l6��d5�1�H6n���̇ͼl�%s�BK���p�PsDkht=�[��5+v�(���|Z�2��x~Ț�\C�� -��-Ţ���B�1]�]z>������6�����V>K{ݻ�W�bTb\6�{J��V��
V�խ�8�꺈�\���G�vk���Nl�T;I�X��}w&��t���CR�Ȏ鑷���9��T4��h�Cd�0A�t���<����Z���dC��Fu�j�ϫ��9�_���&���1��7�Y(�N՜[^+2��q�[-�����j�L�{��n�yta�	<�#�z��G	u������Rį�Y��s��~�ys���cv�Z��Y����P�u�i}K���J*V�%Y#f�YV�&/0���ꭝ:j��WA����p[7�;4�H⌎yZm�*�CY5B�'m��Eͽݭ㈥}^RK��u�Y�C���nom9ǧ}��;�oyv���C���T^W��=ryA�oR���v={�z�g����,�i]�}Y�[A6v����*��itZ�˗:f^����{����#�e'�O�tSS�[�?<��X��j��me׾��#;<Z���q;*#{�S��g���m��œ�:��e+aq�
=`V��1Y�v܃�g��l������9xr��?ݸ"����_���]�>�Sê~�>�K�~�om�>�-3g���QQ�V3�Jق�Rq�t���V�jw<�q���=�fŷ�.�o(�̌R}�7�)�dM�H�wj�P�V.uܷz��hG�Y��[^��yԴ��m9ϲ���b��?���z�hk���pӾ�.0qU��}a�X�W�Γ:��XX�+Sst9�'26���X�_@9r�A���gS�Ό:�~��W�a��Ȑ��p�ٟ(��ڱ
���E;8'��g
��S���lL�M|����s0��=�m�9�y����l��r��x��#$i
�S5�L�vS��d��wkJ���ym��\���L�m�1)]��C�ɯYA<�FHJ��ر���� t��m�9o�:͵7��:T܊���|�+�Q�94k�в��@���;A,�*�g��[g4�	�tļ��������8k��m��JEg�TzWu���M����Kͮ���1�&���@�ڡ��&�Ϙ��k�)�}|mi���i-n��c�������Wu{�dh�X�Y&�m7�wn��#Γ5�k�ͫ/V�����yX��t��_~���<���Ґ�9�+�Q{O�9g�t�q`�L���;.����w��$@�#2J	ۓ7~gfq��=�)n��;	Au6���V���5u���[{�&�	��ogˉ�wxr�ovI��s�(���L�RN!�"�'��|�k������Ca�u�'�(=��v�̆��*om�m�Ըܘ\���.��]�ƨ��;/5����ѝ��;o}m�&�b�1�ZUWa1 �B�T���B�Z�\c2��v��-���f���fv8YR"���F#��t�"��f�����y��_�֝�zi���&�[�Mcy��Q�A�5�����~�$���{�pݙi��D)
z�;%_l�JViay��h�b.��:�����wyb���w7k&�c���[\���f���<�<��x��C��5�[T���n��_Y���߲��P�_J�ҟ�zV����L�f�Q��N��7��q7>B*�u�������!"!"�T�t��z��qV�r������U0��o���ZkyLO��/<H�Ҧ���4�Ρe�W�u���_nE���;i~>��ܱԕ}��hפ�Ŵk��Ѓ*�����uGku�X2ϓ���}����L�܅�N%Z�pC0򾂟-�ʾW{��S�
�8���M��7����.�B ;��g���Դ�j�V��oW#��݁����d:�L�{5t'�e���p$�qFp������9�4���Ov�R/��j���a��1���(����V����dl���V]�nO�g�<QF��WP���]͚u��u5�i��Sc-(Z"��Im}�P�>͙3C���%"od�wy_O�+�+IE7�{��-���1�^�<tVS��Ȳm_&��c	���K *7��M^<�DA�kǊ���ӝ�Y�<��h��"��ن�o% q����~l>�\#_�7WS���ԇK�߳�ب���kn>yٳO?s�Ÿ�d,I��W��.�;oگwGw����%N�[m	�f�`��C�LAF����2�8�;V���3�d�>mӑ�=\&Ζ0f,�tϵn>���ͥ�K�[������j��u��r�b�D��^�U��l$^�^�H錑ܱ�>c��o/#���P����Ϸ�k��4w*0^K��KI�'���X71u�3�<ۚ�X��tN�׮���1�҂�v*ק�� Fh�
Y����u��G~�C�����4�}pHe�t��=�bы(ls�FhL���\�\���rw&n���7�����W�y?��&m�;m$�䙒:Cu�-�ql��Zʗ[�-��y�+��5�~��{Ty�Z��q�8��������vLv��x�����������p؊��ѽ#7TH$�!n0�ݽ�*�*�7_p�p��I�vߧ���� �L�:���X�ӛ�"%�:��^u39�f�L�8��S)�l22<�5O��Gu�vʇ��en_�qWrr��x�U��GQY9�q�-�a��ݎSo�ͨh�M�jo���i@�)�7�a��Σ���V+����lNӳY<?Pm��P��3zI�غ�W�P�ɲ)a��h)u�T��l���j�L�>zK"����֑y�U.Gs��Φ��WW�cN��]���~�K���Oi�6f�r��)�0܊�$�馹��s>g�r�g��f�r����Q��>������ff{4rf��A��ac=���<�reI��I�'gyjRD`�B1"��ꡝor�lv�[�J�'8f�[�S��L
���<_cO���f�<{�| �'��6s/m�wH+��l�ҝ__n�5¥�%^V�P�ɬ*2�s���}`luɪ�j�*���m&� Vn�u��Zo,V��V��Ón-R��݈�t}]�V��%�IY*�>�Z��fa�+b{{a��K% ����u��ԁ*�c�+V���y\�z�(Xam�Na�ثbSu![W���א0�_S���.�:W,�9�\�h
C;T�Ib�]J�`��B��.�t�����i�A�t���725D��Gv�Y`-�s�����+��0!K!���M9*�T�!���uY�΄VS<tQuu�K3�ghP!U���v�p���Q���Dڊ����ҩ0����/n5��$1ΔF��h (t�U�=��PkջK2�1��3t��H�4���%$��Fu�{�$.Ux�W[�_f5�D:��x����l�툦`hͲ�L,޾���Ռ�\$���
�2$D/y�������gw�r�����o�7ןn���NL�LO�j����Q���!诳O[�<�׊�IѸ;S�9�W26�]K��T9]37z����4�U��i#NP�[KG��3o!a�ɲ��fj�r� �����xR*2�h�mt������%!��9?1��j�"�M���21����ர��Yu���,��GnS��X�)c��0�
�Å�B�(Iܔ�2����,���,���֫�Fe����xL�B�&�H��̑Cz�k6N74�;�,MV��2�^G����75�k�|��ڬ����12����v#e��!�uY�q���2s��YeP����cw/��6���4�AJ��]�:X^���Ϳy��g�bDSg�H��J�![-���Ub���z�	|;�	�﬎r�pd�[{��sb�ѦﭥJW:ĩ�Bܖjе}�����74J��W�[�;o���u�n�LS6�v|ߟ�Í�6�zs�,r �If����3a��	o*�c�S��2�뢜o����%�B���w��Jz,%�k�3����x�ި��{�nV*�q��]A�aSղ6�w�+���U��Pys����6���
k��yQ.b;(�����[I��7yc�kQ-�]�:!�Y��ϲq���4�5�q��k���`��2%����C	�^7Qb��c�C/jJ����hY�_�mlaymӀJ��bGݧNp_!r�t�A����OH�{�y6=/vRR>F����d�.�N�V𬼅��P�����8D�ʇQP�Tm\�r�B,mw#�S��0_��s|ݑ�����`��*�z��t�^ꡝ�r	�ꌩ�+-_H��C�g7�qjn	q\8T{���U '�����9纒D��\����	�8��KH�ȡ�ë�� �hj����b�fm�Uw$�4Q(l��D�_�$��G:��uZ*趻b+�]�MEtb+mUTT�TE�]5h�V�D�c:(�ض(���lkn��v"6�F�;k��$Ev�qwf"+�u�ڪ6�3���;b����b�"�Vڋh�LT�w:;b�wF�������v*���6�j(����5�mGvz�Dk1=�u��K�3�������DQi�E]g]u�E��s4vb��Wm��uv:��v:{m5TL�RUgK��QUPV�g݊֍b�mӢ�QQ:��-��b�lh6pQMU1ti���%�b�*Ѡ��골�i�v(Ѷ'mu���wqLc3�3C�bmj�j� ���1E����H�"���5��cZ�E�4݃l;5���j�Ѧ��F�kQTAA�ƪ�
*��AQA֨������4�}�ǻ����v�7S_0��uw΅�C�7���`k��Չ}u��#<�IiT9kt�Y»oc�5�W�VԪ��`֮1I��H��뫰�$3w{yI�WῚ�]�*�5I.�����-~�poF��/cc��9�z�jJ^�
�!>���6��
����g�n��-.�bRl��kyV�Y�sG>a����^M��4�r�Ltv4�N�ޗ�r7$>Cq���k&�߭��z��걿/��Qn����P9�}i� &v}ŭ������3{L��V����ٮ,݀�{c��+���?,��=��;"�p
�ռᲷ��J*�t��� q�ę�n��ȼ`0ϱl�㨞,�Li�[ۙN��^䰾�tWO��2��|�qNȼzY��o�d���Btپ���px�U��ƫ�N�x�l�7��*�HsL�l6)w��5�Ǆ V�|�����<�i6�O6[��.]�����.t�r5[4ye#��HxX'rK���C�bm=��B~�G����qV��}E���Fו�H�l�-�y� k��"G-����y]!�_��!/�z�wxyem�����ۤ�z�o[��N<�	�Gv=�sW��u#ޞG�8f�:������/�M�e���>,At�Y��w���L���!Nh�]�]��RT3i��%�/"��5�*S��Վ	,Սg7m�h�����.���5uf�:��t Qs�Ti�����{�e�}���4T��k;�>��s!�����r�UkM���0�ݱ޻��O�y�A�~��S{�r��y4�n�Ž�Z�Аپ������j+E���7c:K���qg�u�4t߰�H�o��ܺ�x���ųN�*���q>�9Q�I����H��&�"�'�+�U����Eoc�q��Â)cƣ.��{A&j�����V�����}�tt��e�.�лh#|hz_����N�w���C�1�f�3x�ܳ���H�*b�����V�1 �(T�8ܬƵK�`k:&�^X�=T���n������0��B�
�x3܊��~����w�o�2�0�D�;�3�����ko0H؃�k%C��9ov�r�R�f����X|��<J�m�zR��{ڡ�k74�ǡY"�w�g���p��g�����:�]m��$�r�0mC�g��^�G�*h��6�B��uI{u�hWZM�(���Wf��M+}��9�qt����;��#�P�b�\|�ӌn�V+3Q��o��A!�WT��:�.�{3����ܧ.>����PK,N�uq�=��P��n>~�R~_�U��r����i�3fCdt6�?�'���N58T�ԎD���QO��ٛ��{�{����c��5"�*2�����vN䐛:�k���Ș�m�g)��kۣk�]�wqnĒ@S�S64��}�����C72���)��<l�Oi;����W��P��7tR�wa���g���0��c4oS<t��sp<�S�g�.i������?jA��턷��;cjoj*E�t�tS�=�t�U�B�j���W�jS��.�����k�ޫM��~�WW�IU�YYA,��N�^2�wzm��؄�'�����n�����)�$���ޠ:!u7B;|m"pj��w���9��w_D��{���&Ǜ]�H�wߨ�nr;r�8�ɨrFCD�畻~%l�g5�9rrc�mOQ���kTS��R�l��#����o��ƑV��C�����j/��EZ��������t����^�N��$����,�����^�^��}�z���{M�	�d79�2٫
e �S�
��7�Ö�uH�׉Vus3\�iO.��⫞��v,V��̌���p�r^P���?.�k%Ϟ#��~�����ݜ�44}a5��K˨�9�7n�$��]�1m��gl� 2�h�4�����f�����O��w�ٷ�s'I��5�M�K{P��ǌ�������~QhY�Ȭ�]S�ϔfz=y:TX'�E�G^�LsNOq� �>�6� ��	{N�'r��r���L5rt�C
��,�r����d�ck�2e��j�=w=��Ek���gt�Ӌ^D2 ,3p}��YO+Fa��z���o���{��y\��)��]l�[�{�WMƍ������UE�k�;��Q&�lIwRcL�gK:�G&�ZSf�׹\��+q�s:k�D7V�%��Dl�R1[4�]��04�9��`��h�뚎q&�<�ζe��ج��5��ouK�j��Ս+6�0�s U���m�߽=:}����Ә�v�&x!0����]}^���_���S�mST�m�n	OE%hVb�Y��������=Me�hKߊ�
����wwu�x����w��D(q�T7YZ\�9���,=/2�ڃ��;�:an�r�Nm�A�A�mn��'�(�')�8qV㫬NtN�M����g���b��(�R�;W�WX.VV<NS��ТD��U�e\ʳ�|��꟞i�"����D�]`�]j*A-�ё�3����E�Y��N�~���!��K�vb[���џ6����ڟ8���L��+#�����=�+~�¯�F�(j�'��`,Q7�]b!�8rfDL�f���m�U�K�KA��+�RW���G�Y@���6�l
�������g���j��H�#��h�v\����t-0�'5�ѹ��ث��j��ӽ�^��[�{k�G�ʃIw,�J��؛6���+��.���Mvbl`�^5�,�e"'[s��+>/�E4ǉ���ݱ�� ��_���FsW���-}&?{����fC$���LY�/)H};>��Y`��Y�X�Fa�0j��f掬.qW��������e�1��Xs����ZF*�mˑ���9��Y�pu-���y���
S'.��1lF�S�Ɏ�gd���NR	*�l�Xp��Cղ��Kxm��xZ*I�����[���D9v�����W{��n�RŌa��}|��6�������y�b~��r��|�.qL���nTQ�7Pe;�!���c�RZ1L��ek�oU���(ᑶF��ME�R�e�ر�!������������s)�|3O�%���orI�i��+�U�#,��.X��<�'D�n�ީ�|ZULi׋�˥��Nb� ��(d b�Rp9�d�[�+6h�tu=3�-��M�e�����7P/R�����wo`������z��K>�OI�93��g���A�!�@cj���{{jV��'�f7�xL�~S��W�ҙw��=�ʲ��eP[ղ�b��MnSO]��M=��,�l^T�W���9i:H�c	e��u5rn��v�͙S\T�YO΃Z�M��!���"=ٚ3y��)#`���K!WVP��@7vk	@�QRկ>�ȋ}���T�ƻw��P^D�m>�ĲKu��H�"t]�5'�U�����r%��_'�n����X	ر���X�/)G�3S[��9|l�sv2�P��I�{���ks�Kz=ʹL�|VFOk�,2�]�ܬ�v(��0�FL��c�c���AR1��k�����r�����nzg���3(Hr։�V���+��k���E��y���䆴e��H�L�������t��KR�&��Hx�͒]�����}��t`5�m͐!o;��O>����R�(��x�q*K%�l�y��/qΐu��W�8��{�̳�ܔ)��Rڦ����G*挱�8�۔F��N���"�!L􄭌���0o4��h>Ok=��|�U�m�øg��
�#0��k$7M wi�1탲����r�Q�.�@}s�.佈��ysl
Ո�m����t���O+�W�f�c2#z����<65���|pَ�j�|�tl^a�ĎI��P�~��s.ߞnI߭{�7u��X�g�����*"���bޯo)��E��{}��Z/��T뼺��)�be���̹�b�^侾LN���آ��ʬ�|��rO���nn��-�|���<[��4�����X���L۹g����wemɑ&|p6��~��]�/e�r��I"��`�zM�'u<��ڋ�!˺k�L)ƛ�Sl4S���w��ηQsF�Y��峹�w�r�9L�hV��(=�X�b��wH��o��&ʏ�T�w�z��̺Yx��u7��`B���-Ԫ��9l��Hk���Q��ށP�qO�:�w�,�{�/�-�u�G����B���*�a���:�,;V]�{D��M��B)��K6_����|ZA�1�����J㩓�Mcr�3u���5N�ŭ��"��6���u�x�n�ZEV�����j��Ϊ�~�qr|�2s.{��"�$%�.���^M=c=ɥ��/~_a�/E�jZq�w�=�����I��%������'{'�-\�7���]Z&��fP�j7~�B�~�wmXKN�M�F�ga�K=*q�R����sýq��UܵnbE�@X�Le�8���N)엨w<����	ڙZ%�5r�f}7����̍�p�4q�2fp1���M��s�u]S���M�.4!���Vl_g�V�����b=�D�>���ߤ�V�X�+/AF'S���"�xK��f�$�_U�c��� ��4b�OJ7���Ԋ
-���#���m��2���꘢W͉@��.ף�u�Y��)����������Ww�-�5$v�3#6;:��d:4ŝ|y�Wd�. 
����C��=�]��G�)�wS}[0*ʠ0gF�j�Sr��d�wʊ��x��g7�qx$?�g�gytf��y��.�NvpZ����ݛ�c�*��A�V7õ�I�B�K5��F�ag�e&��<�*Pu]�=���a*�{6�aQN�b�%�_��h9L���͖��1+ג�����٬��1�eW�&n0��,�J	\�^-���ePgط�i�7[��KC9#��V�z8�[�,��9�<o��������cZ=Mg/�4WW�,�:����v�-�l�x�e���������U��K�2[�쉛O�:f�+n�1�Ґ�b'B�����x�jc����h~$V���������߿b<����یE5�V
wh���,d7WHg��>�n_%SYq�o�a���:+!P�]z;9������K$zIufƩ�:�dy���tH�E/ٓX��[��Tq��D'3`J���}^��en�F�7��p���;�hy2�1e�z�	�aӬ��.EM.]d�H�o�幫,3�2�u7�\kW��3�Y�����&�Ek8>ѪCv�L�3b�}��R:ngZP�������L���qNR�W�r���[A=F�;!�cI��Gm�:�PA�\,΀�w7v�#c�m���p�i�Џ���U�6+���t��<��i�G1F�lȹP��k��f���ƪ��a�Ό�F��S�ϲ:gI�Ƴ�A� {1_m1��"��+��&�<�ie�]�[�;���Oc�n��|�H<��\8%�d�f����^��מ�������X�8�i"�] 잁��]:Tz�g�[�tw��E����j��P�Gkىf�Fwri�Df��
�hF�a�i�.�s�����r^\v������=T�YΠyI�����Q[Pt�ܫA�[k�s��ιr����BzQ��5t�ƮV�B�,�@���Q�b�U�-x���TK�ͣ�r�	[U��sj���1��!r�Y�{=^�4��~^���:�ܐ��ȴھ�R��5"�Q��۬�З�ťN�.�lU�����1V���%Wi�&��/pf�G����� ��$��b��Jh��@-f�rR�7�����<];�v���kk�����ei�	������]��9��9b�~��}0�z��R���ʜ�Z��qV0�7͑�fkN��U�f���rM��g`�ܱ���v�9���Q��qɈu�L��E�e�.\��V%G�%t��@R�v�_9/�P�-�2!��u�2��˸��@ܞS�|��{B,����Y �����=����lޙ�d�Ř	g��Lf��>�v{��w��;Sʖ�ꎖ:�wja��L��Ώ�Z7xѢ�\İ�T]�ŕ+�Y�[k�t�э�K� ׭��m�3Frp[�^�g.�q�(�j�\oi�C�[c"	ը������ ��+�ۉ��@�چY��^. ͏�"��ϵ�]޼���V_7Y�����O=ڹ/$�g��LFy���Ɖ�qɕkV��۬T�,L���Ö�n�o+2Z��E���#
Mͺ ��':ܹ�"�X<�;�������]���D��k9����8��1�2O��:6xXg�K�
�ΌĠ�#��՛��C���s
 �ݎ2�DȊASم�Q>r�<qk��:������/ErQ"���{If��f\� n��S:��m�)�j�����o�)�}�o�.yi��wN�gmv=�;m�zs�z�G�w�C�oP�jF@]������$2�%�J��Dv�U�Y���g��<~��=��w!��7�ϑ4o��)\�`��T�u�SIŵ��<�Q��n�'W �l>���jI����p����;���.��2�-��7��(�)�h�w�����c�q�9����0�9U����X[{�iR����٘�f�ER�R����\2�_�J��4�n�nf�-��
��ނ�0D��������W�yI�|�����?jF�}!xD��	X�u8hl[ �.�%p��M�ݚ�T���wr�Y鯢얪
�b0���]� 6 ���$v�HY���^L�z������i㼄�]ʍ�Q�	���KKE!�S7Q�Tdi���Sӏ\8m�V�R�"�cɳz^af̒����pF1�G�+w��[�����gN0vL��ܻZ����'Q���MuD�aBݯ�+��yM[�ѱ&ټǰ�6*`���JZ�O+\�vr��F�+J�R1��t�`�8�`:(o���`��M�h��i�M-1s��H IM� Ρp1{l��e��h.5?�sW�+Y�7�{� <4���`�e�1V	�o�}���1c��ٹ��Ա���8��@�c,�z��EM��3�os�ʵ����{f�f���J�]du�V�8�w*��k0��ʼe9_ qhw��C�r�դ�n�\�:Ma��ڽ������O?�f�ש�u_��Ω";��M����
-'s�b����d��:)�4��u�T1��F٨���m�v��������h�1L�LET���Ѣ��H�"���� ��<iu���:���.��h��Em�b�A���h��;n�4f���D;�ŉ�[7q�m��i1=/T�GX��j**��(��lh;a��c��E;&���'q�w[1U�j(����%��h�Tݺ��٭:(i�P�bn��m�h�*�Qh�kUD�D�lh$�)n�*"����Q�[�t�&�DQh1Sl���#C�B]8�f�Z�+mq"*g��D[�Cv��5��������!�Ѥ()�{�QF���l�LKQ%4�V�b���V�:�\UvC[j�*��h�DT�8�5k5MF�vt��-�]h��$�I?3�
��,A��ԗ�^o�]җN4�����ւ��zo@J��sQ'3R�Q�/�`��o#�5�-�j\s��y�|N�
�{f?���x�=c>�J�p��U��b�i�`���lc��w�b�aїO���i���"�����&�*�
ﶽ��'��̃U�Gg�����7�W��l�68m��K��$�B�*ʮ���yӛ�Ͳ�7�ur�����~�^JXi�0�t#��]"�tnw5�I��c]=Og{��-�ww���B���9�>��:��m�U�LI�Kf�m8�6\<���mݑ�Ss�O0=��${��������~���3�o_�z��7��%���+��7,�sZ�dw�����!��ڍf0�R����+�.Z򉔶�R��G����T�%Lpw�C�6�m:{�76E��N���,��\�OA�'lvK@��LI�4���b۳ym����^�s#�׸��"����G/L{��p5��q�Ӽ���/��2��Oá<�{N�-G[�M4��'���ݏb})���4WU��4f���O��f$�����k�W��I�{�wX�F��=Wq�Iդ5$3�47G�5���v;�պ{*2�3[6�_��$��>��F�.{��Ym�����g��W�g��	�����*�`��Ż�!ə̮�A]�x�����1�VH~�7����8ʑ]t3)oX����;�v��mvt���� r���ّ�.�q����ɦס]��w�(Vj#Ƽ���V�I�}fQG����P�Z�&[����%n���6���C	v�������5��K ��*��r�7�۸�5ݱ�8�Os^����P�ɲm�5ђy��(�X��4���;���u|�w\��YT�crl�A[dX�����Hߙ�*IԮħf��p�k7;��������s{z���Y��_�Ɏ�+6]�w����"�s�e慄Du�d�/=�ǰ�%�������@k����zbaܶq�Or���s��<�'U�]a�v*m�f����pe�_�����G�9��C�-��x�k��XJ�ٻ��=�XM^|��.*��e���"��ɍ�{7�oPV^i��DM��KU����+�R��Q�;+%���������N[�����x�_-�a����lɣ-��o��ʻ�w�h^ʱ��8#��ĴoUT=W]�l�جƛ���|���ʫ�N���Ֆ��B����|��[M��7u�gw
52ڙ5a�������8��&?�k������TE�����QY_K��b3���'��Z8j}��8VN��$���gʜ�ᆣ�����[wi�8��!��6�7�b���`Ϭ_@�g����7��tm�u���U�	�3�굈(X�4d4���d2/��Y[�'��b6�����ͪx�V���v�M�<c;ˠc6�^`̄�{g>�G��`���V_<B�8�A��̇��z(�l��Y�ǩ��x�}M��V�Zݸ��M�^�&��Wg�)�\�y�Q�Ij/��l`�꓿R��r�$h�7?~lwM��ĩ��;�+lA@U���-�r��T�"0�D��UTFN3��j�eG*96O���Xuߎ�)v=Oy��5�_/#�e�],�!��îU��F`�C���I�I��ޙ}-�.�1o����ߗA�⻆"ߐR��zuu`b��{!�2E;#R���<DS0�4�Օ����ѷ�N<�C���VQ�� �!��X��Q\�7t�H�P�fi܂Í�9t���>��q�$bhm�����JAW�7�*]�a���Ks�gb����;CD�t�ޗ��)�O��*���sd���oU��"�|�lSP�bc�nRwL��Em"�Fk0����5�uƋɵ`�ԕv�%����'���k)B��N��o�|�yT��^Ϸw�� W)O�k��rJ��<̄�kX���Y��NX5ޠ�4}�y�{�{k�����ܩ�L
�[�+�i�?n��ƺ�X����H}t:�1�F���I���?ޘyd٪��L�O1T�s�X62拈s��S��P3�3�>YQ��hd��Y�V��A/�{:�ݝ�ޥ�1}e�������z�t��\�2�|E³��Aj.#n_�v��f�t��T p�Wt�HYd�/%7Pe;��(2�s��{�)�j�	���>�K��!�O_��$6��<,A�[O�2��g^������ݚ�Ѳc���'+\x2�`炄N��b��,-2�|�e#]\� -�mŚm�].���Ҽ���*4�S4�������&ާiި�v�֗!�wN`�K�[�8������R|�?��RY���+W�"��w��h��[�޹��f� �;%^t�U�3φ
_��;�\8Z_u�C�����a/\����)cS�����m�xC�CR��E����ΐ�����Dg=ǲ�Z�T�r=�]����t6�z��WS:�@���Բ�\�C\��?ߐ������Ü<�xVE%��Z�3�^䶶�ȏ+�x�&D]�8�2�H�s]/+"�M���c@T)�K'~�'�䝫*��̢�Y�If�Qq8r�q[gꨄ[�S�$mn,��#La,�Q�����o*�9��q��m��3x��k��^q;L!�7���һ[�I4,�b��k9]=q�f��9'�6u��r�u���A`�*u�u�+���j޲�6fU5�w60�*���˟:m�9>nΘuθ�66Ү�b�N���Wզɖ�Lf�x&U8u��6�w�g1hSd�38kfϔ���Fg�8T.�F�I>��?�P����2ڮS(��sT���$�ov��+ҽ��Ԟ��Mf9�3Wd=\�i�I�䎅k���4�y2DP=����ɵ��1]��&0���LK;��h��mQc=��C՟�,Mvf���.��$�BKVo5d4��v�E`����@�����HW�s��dm�����_�J*V��7k#kM��	�YF@~G�U�'�i~�3�䭌����N��Rc��\�a�/g����Y���lu���r��ei�m�6bIcA��[ͦG�45�ٛ�[|�g�1��7 ��}z���GHby�����E�7wv���CTU�1V�^�m2��i�B�17ʷF����-�����V��~�m칱� wP��c:�S>�8ґ]U�kQ�v���e�j/'�4M��G:f���{V3G����O3�B~���z媗�wKuJ��*Qx�+�l1)�Va@�+�vP''(i�U�J��6��bhY�0#���u\^��q0Ҁ�͛��ef����UY���P9l���g���x�R��]wϻo�<[T{)d�8�O�����@tA��IvH�Sv30�aCr�_�[������,ɾ��x�X���	{�U�6����n��r{DTyxT�׶�ů��ͪ�&1 �wi�cq�Ɣ�S
�(�}(4͵Gsw�r�����J�e������e���,ճ��f��񾎁��>�e�Ѕ�z��d�5��l����ȗ����5L,�PuǴ?�s�W)F��5N1������;e�cY>�S�Ց��M�� �[Ϻ)��r]Q�t�i��.ٝc��:��!�d��_Og�զI%���Z��;Cl�~�;���;� f�=NOkZ�8���u34�s���/\uJ]��ح�G0C-��v��r0g%�ϝ��J�{��Oʭ�{�VXKL�Bۧn}�7���[a۬��|�=�&8ИY���rs��,YA.{6�~]8g3n�5cӊm����#\�J礽��ئ�}J��7:թ�n�5���&��g�_b�~ɉl�w�m��ɘ��L�v�ׄ�w�2 +�}z��IݼM����]�.��֞]`��g���}n���Vf,�Z:���\e�H��m�F$�(�HdrF�C����C��
�����Ӭ�y���1��W�A�l�v�*F(u���WS�od�i�F��3����M=/�Q��}������b�i�I2U�^�K�K�<�{x��9�n����O������X��Fy��V�UZ}Y����hwJ����K��'&pǒ(��G���w45�}�15wB�ǯ2bwQ褐��**f�7$��[������.}>��Y	�Zڹ�"���0�;*��\��F W ^x�Ү/U�L+�č������/���-�j-�kU��Sp��:a]P*߯����D��C=��A��w��ߒ%�c(�x<�C�f��>���Y��`���cN1vm��5sQ�K��3r8ݪVD^2�f�,�<������r��U�UMqx��%YT��{^����q�u�)�pq�4�)g�_:���[��t
�f�^�\N��\� ���C��"��Co��[w��e��#4�\p+O,��j�{:yU��W��yZ_�
�OC�1��s�Ŷ��\?)z�6ު�k�|:ʂ|���C��)���cJ��s2��(�Q�%�}��K����jQccz�w%�P��a����]����,U�̚�z�+
����ߜ�Q%XϏ�s �K�3�Q��ܛ���0�j�j�w�f=X����	�w�Z�̦|똼�^8�arʙ���2�e������U��1-�x��I�q��O��L�35��v1�Y�ᚥ=��'r��������I�g���>g���F���'�"'�3��v�N���G1�8�WQ�;�3������{]�8e���v�,�M�α7�{�}�����K"��y����-- $m<��O��gO�a{u4��ݫ%�B��!��a%�0��푧G:H�R�1�u3Ѥ�I����z�!;2s�'L�&� '9��V�}Wp�7E�����ױ;d���n��jf��m�j#ly� 5*��3u9ts�(3G�P�eI���������	���Lq��Cw�c>�)Gz )����E8	�#�*��X�O3�mop��:���+&|���2�J��/<�[w�r��k��d]*�@�
��2��wO��%x�����TV������V%>ob�~��K����#������ѓ[�@tL�1����$�M���U�X�q��R\pt<QZ������z~||A^��q�f���y�oC��X�J�6�m`Ȭ�-FSam@�yd"�|�b�Yu��˖�e�v<ә�j�(G�7"˫5�*m<�qfV�h\��h�)�I�m������Y$m)N���^����r�lW���K�7$����ebg�{�1;Փƨ�9fsw�S�e}>g�r�����l[�37���⾗Jb�\�׌8�	��g��g��8�����yO:!��}��ؿwO�bt-�-l��AA��Oe�_'k�㳤�d��y�h�)�w��8e�0���+.�>��e�[8��Th�<�h��mⰮd�2��8�Sn{;�ў`7�F0�dl�e&�yfJ�/_Wt��a����k,ya�-/Ҧy*c���-\�u u\?Kfb�3�!�Z j�]t�T4�x���'�m�z���i���u�V�{��]����\`i>"�2?�Q���=����:�A��+�dʻ����u5F*0*>�76}��1�V��0�ڟ��]�~�ף��$�F)SQ�*��)���<td�E��B �c[�=W�������?�?����l� *���������!�r+����=Ã�}���!�ÅbE� �V X�bU� �d�
U�Z@)V��E�@P�DSٕX���J��"�����{���zEVUX P��$U`�  �U�V	UX%U`�U�ԙX!U`�U�  �� 5�U�ª��@ ��H��v@ �H�B J J J�B J B��  A"�
��
��EVX%U`�U�EV	UX$U`�U��U�V	X$U`�U�V	X$U`�V	FQ��Q�Q��A�E�A�F!�b�F!�bQ�F%e�b�F!�bQ�%�=������|_��
��H��Ҩ�3'���������p|}���������������>������E������~�_o������
�����?�AA�_�*�
�����>�������?�>��!�
����@���/�H�~����?��'������b���APVU�UiUZUV�UbUV�U�UYaUd�U��U��U�A��P)*����*Ă�P�&;�X/��~��1TV��h
 �G�������Р��O�=��|~�� @x?L�����}�ׯq?��?�3����~�ܞ���� *��އ�'��߂|@��ܪ *��>���ڈ���?�p�_p 3�����~��������=���p��� *�j��~�� �*���������}����}���}BO������W���������������_��1�`�O������_ ���}>�'��� *�'�L�����@������_�|��j��+��c��AA��?�������a��S��(+$�k0���;0
 ��d��H[{�)"BJ�$T�T���%T)RT��*��	P�B��BH*%T�HET�J���J��"�R@���HR��ԩz���Ѣ�%UE")Q%B�!QI(*��T�$T��U�"T�!B�@��$
k�RUJ��UJ�P�@���T� �QR�;4٩B
J�	JBIURDIR�T�JQQ�P�R$���JJI(zH]b��<  ��t��E��:��tt�-�hi�me2�)U-��CEk �#5�H,�Jʔ*�X��vt]�%��Jh�U�ڔj�"!R��kP%W�  faСB��4=�Ӏ��4�
�8t 
(�np�P���G�U�@͕{�Z`�laZ�WN���`:YԮLԠ4��6��� @�PT�D!  q���Q8j��������Ԧ2�mR��mJⳣ����Wn�M5���i���J�!���JSN�Sw'Z+Mv˔w��u�TR*��DDII�  �x iz�ʮ�SwS�m�g��p&���!vݵ1���m���;��]���i]�즍�v٢ҫe`,N�@�.��B�[%AR���jU ��  �UU �c�u@D�e��LQPՁU(�2A��)Z��W]���
Ʋ�4��(�T��I�  �i�k  ��iF� ��ݡ֫P�Vڢ�1���` 
�5P ��fځCb��% �A@��^  k� *4�@*��*���0j�iB���#j�%�PQ[)` 
�5P �` i`�$�T�Z�R��
U\    :m 4 ��
 �`  A� �VP MV  �V b����V� �J� �����D�   ,p �`  +e�AM��P & � &� = �����k� �C  �6��J��JR��$"�O   ��� � C�j  0
 5� �7*�  ZF  2�  F D�� ���R�Pd21�{FRR�h@��ꞈz� )� ��@ 4 h�JT @�H�2�P  �Jeed�'���Z$�eq���T�ABW�'e�j��U�xx������`������!$ܒ@�BC�a	O�$I?�! BH�$	$$;�}�kW����C/m�t��;�a��	3BEI5㽲2)5�A�]�ƴ��Ef]"Y��Cha�2�H�ťr����B�k/i�\*����N�^�v,�n�N�ۖ1^*�[J�z`fF�J�F8ӏP4��)j�n������|�̑\�#��֭��v�ݻ6	�GII775�f�
�ޤ�1�p�a)�w.|�LgW�H�Vb���dʺ�B\��f��zE��w�m�6�=8�&r�n�1r�
f3X�5Q�RG8� �H�ݤ&QӒ�72SyVuf��P�n�a�l�"Ϊf�S'@�5����B�b.1�n !����1��H07����.�=�2�N��˭v�[��@��7i�ś���y����sV)�*twu�V�l4#�j���1Xf��˧�dL���v���h�UCuyJ��ٛ��,X�Jʨ>�ԭ2�o�i���>��k�Bڟp,��y3~�@���k1;�a,̗E&�ZgkP��$�D�E�Ƞ��!�Qk�[���]* Md��B�9c-���v$��Cg6RQ�`|�-Z��^����֯7[�����3v��.MOW�5S5��,����l�t�P&l���*��Һl�@ ZeČ2^�˫̴��*@�͖�S-�� �1C�V	bTK�,�7Gn5�Z�
��Ȓ��2U�E�ʴ)V�5,�CB*j[Jā
J��f�B^S�����O&!�w�e�Yv��ڶ�� ���a�6�:zV��K\�@ZP���-�T�F��ѻ�k5,R3�;H��B�Ō��YSiJ��	0C�`�l�{I�Rn�f�Z�%��X�#NQ��A�y����n�N��l��6V�t��&K�m>B��z�k01��J�m�q��ʌ5w��u$�l�Mf�]�*�z�M:�̰�q �Ko`s�fÚ4=�ɿ8ށB7�w0���QfJ��`��V�ZZ��)�O�b�&��;���:�] �*�Ig]T�8�S����[ܕ��%h���ޛ�2ÅR�F`����S�$b��������*+�GX�u�a���1`�c�&f^�m�%�ƫ^b��Jb�nV][
����g-�Ө�K0K�f	AT�[ 'EҨ-�f��7R�c7,�[�wl��Un���4�핹�gE�GTiP�(vB�m�Y����L*_Ȫ��7)l��QMJ�*�f��Io�*���+�����C5�\�kV⼔�	�),��e횳�ڌ�T�9�L�x��@j�l凂$	���j����]����rl{,l�2�� 
���3��m��-�̈��ظ��m�Mǵ�[:/6Z&�i�b�w�n&�R��� �V�&\+5Br�te�-u��5�O�al�SVX3�u�#�w��Fd--�(��"�٘P���0T)�X�S)^:����Ee:͛
�v@�[-c���i�ġ�JV��os�4j��^��
yYbZ��]&�¢�i�;��+j�&��L��T�-F2r��*]A[��n�x�y/��ƨ�ևۦ++d5-�dG#��<���1Mɐ�W�=�a���J$��UL%[�3�7Ff�F,P��q��R�J@�t@�חT���XWkQ.�Lb}��;5���U�l�6��al2#N�f��m*�����{rԡ�[�H�R������u�l�J��[��C�di�; lԭt�<yW#;YIf�Z-8('�<4��)�r����t�*�bǬ���C���x��t|����okx�ӆ��v�+���fݥv�4��=�+GE$�%��4E��N�:�P�N�r��e6tnAXp�˦�M���p$���I��Q�Lv�0�Y̗+qẊ+[��D<#CaL䗰զ�!C ��9H�Ma�v����Щ&����e4�H�g�%D(����M�1�v�� ��V�L�#�	fvQ{�헗�A�{6�"ϢP��$��g)+��f��+&��[O-��j�K��ӊ��dV0RD��|3Lzhe'�i�6�.�L=��K����/j�v�$�E�f@�dd��Xt��R�̹�}c2��N�̗n��W�F�H-U��`A�m��m�|V9��D�:�+�qR�u5YymJ�b�Bƒ����!�$��Y���-eMۑ!Lt�D���U��e�j�㡡e�푲,����s�SFT l0i�m�� @`g;�E�͙1+���}�w��B	[�EG��\��C[�4E�Mm^��Ӵx�KQ�J[�50��+l�y�*S-ʎT CHHYr�YV��.�B��qf�V�)Դ��`;ʴ�^@u.�^F��	8���M3q�,��Y�VG�+ʺf�d� �Q��-�j�z�p^�r��6�c��f�Y�sJ�7��1b�7�(�j��A �u[Ԅ�k1kv~�1L4Ȇݍ�*��zи�j]]e���4�o�fm�}J��e�V@A�#˷�Y�h����]mJ�;J]7If�֦�/F���e=qm 5�J�/�ݺ���<�+".(�VV���y��4P�t��wv����:�Ʊ1��5�a5�Ɍ;�͢��7v�k�E^͑ZHi;)n��T�e��<��mLJj�5&n)yA@�)[@hf��A��3�cSzLz�YJ��q:1p��m�^n����v�v*�v3�V"��Ȗ�.1T���;�*�(ݷ�r�R�4^�T����B��Y@Yj�Ȯ�M,���j����O2�)'q)Q+�p�S��x�X�d̋(�1R�$���͗���*���[��`����ze��j���Ӻ6â;(�J06<�f���TU;A�$�����̕���V��(�FS�^ʔ!n�/XőH3c�/��Oe݊v�ݢ�$0,;*Qp=�����i�ɩӵn 's��	������e�)�F����tñ�x7F�v�P�c�ݣ
������)�7Q�%2����݉H*�Q��e�2e��*��N�!hn��sm������B�i:�Ĳ�.R�h��]ټ�;���a&��t��M�r�B]Ĳ�Z��e<WF�;j�m�آ]��9� �if趫B7a��]�B�SS+oRJ�,���z�|n�=[@aˑث���)�,;W�k.�Q�SH�*��I@D�͠�m�5�&�-Z�Yk��2��t1��>�����b<��j%1���84�̩�S�S"��)��C��+ں����cfU���*ƌVwW6�-CX�u7A�Bu��V�N�b�e�IkP튳���e��Nc�{[Q]�(���<���Cw2��Mǎ��M�Ó)G�%�ق[>������ ���b�#wbǒ��/�̡��	�
�%㴦2��(;.àX�E݁�@�5j��#1��8[[��FrT���%>C5��QC6��Gj�5ek�r��el(\�G)އ���0B�Q�C4h;J��� ]̵J�Y�\�R�taՌ�E%��+]�v#z���ś��uՇZ�E<��Z-�[7^*z�R֋�h�s|��4�U�Tv,�ݩ��)P�ϛ���q�U�X�^��2�lڎ�	Jȗu�`nJ��,�f�w���ۑ卦�,�����tg҉�V�n���li,d�y���f
1i`�BS�v��`�Gen��{B�G1�7ߍn��osoF`�!S���n'�r�<*�
��ᎳLoհ[+Z�k��$&2�_I�6�S��T�Z#9�ѥ��ʹ�f��ʒ�{nPˋ �X{������1�dRtvP40�o+bq妴Ѥ��x!�v���P�H+�A��j��	Ol��������f��5Qb����$.f�򃶠/�YF�6�t]��7n�M<����$i5ٍ^1/,Kt�r�������OfS��"0c���v��Y�s$���.���㔵�OL�Z^��Z5䊝�+�FLIS�D��;�U:��� ��A;���$�y�D-�֑�.ƼUi�Z�4��J�pĨ�xօ7�io.�������V+AbE�E�5��Uƞ �ܠ�C]���pS��-С�+�-�i�[4�cXӗ�r�A�(�:f�.P�^����oف�_GK@�ui�h܌ �É���6��j]c��Ka=fh�tYm�*;{�"�9u��4G"���fi�L�B��e�G	�o]��7(1����zF�0�ՀeF�j�m���ߥ����Rٚ��+$S1�
3Q`���F�n�l���t3��a�;�/�6N9v���0���F��2ռ��'x��f�8�֣Xbp�n��h+��*=6*�4[�w�a��c:6n�J*���M�$6���O6���ZeE(��u�-�z�X34b�:4�m�Z�yQǁe-6Bغ1����w�
.oԫjU�m�*̲*�Gcm&
*=�8Ar�+H�b,�V�[n�3��-�f�l�u�fں�R�[IF���M���WE���F�hNj��Yw{�ÇSi:m̸�a�Um��y���2�Jb�Z���3��2�%i��Ө!!��A���n�^#��b�xփZ�������`J3洙�Q���i]��.+mA�ac�y��S���OMC��u\X��ة��U"�Jj��CC�w�ҷYzY��K,M<�Գ(��b�z岮�26RV��n67X����֦����Â�Ѷ^����4�Ӕ��Pnހ���(R#u!I=1^h�Öt��aJ֡)�ʓj,��UU�am�LE=@h*��Ô���7!@m;1�a;��{�-�m�!�e-�Xeo�$�PoZ�����K�B���uV�"�U���G��5{�aS)�W1Ѭ�Z��Yd3v�gYݘ��fFȫ���mHiSi�P ][�������@f�'YM��1�[���L���
�z&�7V�cn�I�{[��Y�t����Sv�ؑ��b:e����d<H��K$��؆]jmJJը�(�
����e\1+¶��N`$}�7-���j2�yQ���qcŦ��)ݪl;f��Y����7�=U5�㣢���h���ZW2,�5�CJQ�:�x�W�%���m"�%MӮμ���n销˒U����Y���Ot�-����t0Rk�ji�#\�X�J��ϯ$0�r��ڀm�%�V$�c*��GB��+LLf���x1INL��� �e־�����톓LV��z��՚sh��V&�j2���%)�F�XD�y���E�Q�u��ٚid�E�1��f�m��(�VmH�+��t]&�Pܣa2F[�("�mR����	``^4�Q�i:�{E����i/]�B��Z�$�������EY��:����(2�l��]m��X����.૊F"�eՐ6�"ۢ3�k&�X�n�q+��u�U��z�(e��hY�r-����(lԋCrD
*U7P0�X�75�!��eH�x�`�$Á!>�U��j��z1d�I�&��MSk+8��3af	d ۥVo\�6Uc��s
��zo��SԡI�Z�-v��V��JymeH��/ U��	��P
��tH
`����8��m�&����;qÀ:�T��[����mQz�@R��F�;Ǎ�cQV�ɬ��w���4�bI�gi��a��n����4m#�̄(��]��WQ��
(����H�NX#,Q�Q��
\$�[��n����"�tv�m���4Ȃo]eSL.!5^�mh	1�nKI��ZU=ZM����0��5��р!x\O(��[X�Kbܽ����3�L�h,�U�L�t���{�4��:t�g0f����{���U���	aU*��	e�B���dWd���H]��`��	2��.ܗv�#M���-�P��1���-�<x�2f?4�4���X�9��t	n��S�Ʈm������Ҭ�[Rf�0c�ƹAX����)Р��.R)��׀=1P�j�̰r�U�N922�s��Ү(�^;�����dk�KkE	�kVRY����%�2իn�s �%1+#�vV<�o+2�
֓F���9�h��n� ^�xl��Gm���b�%�� zTSv�@�{��WO�j�v� �ѡ���Y�H��x*��y6���4j�0���AB�\�M����i��nd��>? ��&#�{Pl��h#ͻy�=����k����J.�(�"aw)ZOM�F��˂:w%]�l��*�`�����.�a�6����4Rе�KJ�w��3t�,ӥYy�M�k]ܛ{�&��F�7i֬ņ�:�ټYPCEit{m�sj�r�-��Ԙ�FZ�Aly�����m
�*�T݀�[o~w(�ճF�Ġ�4d��4r�]��bjǛ�9%YN��*ķ�kn��s(�v�^���X";�����D��Զ�R�W���t��o�ф������ͩ�kq�Z¸�	�eh�)���G�aH/��e�p
FY�����]$�s1�1ܺ�nҥh)������Ǚ�T��SlZ�̽MQ^*@��T��0�mеV��IP�MTZ�[��ĮU�)�e0V������ 	
6�i��ݥ#TM����RU٥f�Kұ��a�F�L��B`˨WZ��o ��n�e<�[��[��QsF�Rb�@-u���e�tЦM�s,��W �VN�e��_cr�l�I��9�3h2d�.�	�V(��m��%��Z9gpK��jr�8�[6Q����e�$�ѭ8%]�o#�cwN���@�d��Xu�bA����U[�x�nܩi��Ea�N�EY�E��I��t�U�,��f�l�� c/�:t��Z�wl��LЋ�����ӷ�����N3��$�Y��+x���;=P8��R����&M��6w�N�}�t�x�]�`I\K��;��Z�YӒ
�+8��y\�T�Ӷ�J3k:���`QM�q���6aT�w*>c]v�U�7��u�u1��>rr�����ۺNhY|ٜ|y�ĕ9��V!IJ��g��wZ�7�!���
�q�ɖ�GU���䙽���!�*5��`{6�������T}��}��#��6��b�w7��ls�Ck��m�h�ld@DzkZt�2v���*s(ݗA�h�Q�^)wEѶȽ9�;��1��19���\�.D;��j+�}4��]M���Ѐ�N��9<�7	릆*���i;��p�")Gn�D�Zn.��`c��j��v�׀ݴ���:q��Y}x�M����w�o��.�S�4����ˌfESK�NՉo���6Z%�}K�v�i�x���k,湮�x���B�{����,:�c��wxօvUn+�3]+e�7[��:�!x\rdɑۂSW�}d>u����T�P�]+�V	\0<�HcP�/J��7sc���޴��]�z2��vƻzHB��������CF�S��uʖ�`|�Ճ�^٩n�I�!���U��fS��+F��V�)N�ͫ�Bum��
�.���2S�
��`�����g!���y�����H�� ��ܝF\F���V*�)[AB����4�PH��W<2.{��;\�Pr`���L�\γI�/]b����vb�׼�k�;Y�^P���Jݡ��V<���97������sNP�7���Юǻ�;w�Q��ʹW��T�ɭ�de�$�-�v���O$ũ:I-�0�U�<|r���Ϡ��L�OF���R��h=qQ�M�O���[zW;��5��+d��
���TX��g$�.h�ٴ�7xE�nʘiNݹ��)t�yJn��<���Fa��d\�0���֭�2�,�qMΧ]+F����Q=����*@������[ g3�D�mMr�=�b�,�1X���x���X��V��o����is*&�����S��s�M{����Szj�w'�\���^rl�$֍�x�
6����![�ȝ܂�ݥv.ƾ=��`Yl�[��n�i ���yo�|�*��}�5��d�v23����;d�)��0��(B����6��|F��k�˖�z��j�K�3k-J�s��ds}��f�O.��сcݳu�p��E�畕������ٽ�9���9�l�ctEֻo���R�
���wU�J ���ǣU��{õ\ֻt�����9���ј�n�.FѤY�(�X	V>�a0vq^��*��Uj_\�'zU�]x�y�����b��lsRb�x�E}]ڦ>f�zč�v�iК�.��LY�d�7X��i��M���1J�U쵪��1;�`Qt��w�1��b?`Ykȑ�z��:��5]�Kkq��;- $32�sL!`Qwjkϸ(DJ����bd�L��7{-��-����l%O�U����DsG`��+�gl�gP�Ƿy��&sއ���G����oXH��v
�S�d�$�q35fa\�Q¸^�"�'6��{��̕��&~���wD��\����B�ts�k��w7-W�]��bX��r�e��u�:�*�7����7G=�`tjѰO6�L	�l����P���6�]_fbY�颣B�^���{Z��(���ΩǧM�Uu�ڴ�|��h�k�5��iˎ��,wH�i]�r����JWd�u*]��t��讗m3�L{1�oq��+Z�G��}�VY�o���1;�oḇ�:�Om,�
t�R�f��2vkFh(Q�ǑҊ
3�d��_*Z��l�U��C/H-vC�\��Y��&��g?�]��c���/�Rv;�y��+�]���:����`D'snh�ܮEow���30���3�(����w�> �l=����,�6���+�:����"�e_=�C��c(�+6����{�7��s�-�=/y]�q�E�z��K�Ճ{(S�Y@�>4�I\99x�ʼ\r
J=m]	wxEw[���j�J���\b�NZh�y<�W�ö����Ju���ѓl��A|�P0�V޵BkyW!�啔����s�$����,q�5���3��\%�y}SgfP�h�"�1��۩-%��D�f�F�t>��&��������]ruf������-�[a]���ˈ��[Pm&�'ǛWR�[�Z�K�r,���z�ipOE�7φ�	1GvV]��a��2���Qֲ���
U�Cf����Z�.l�2�c޻�D��ˀٛ}� e��gJ��\�Y������VF�Q[���U��gT2�>��e�G���oi�[Ҟ�W&��c�7�XhR��+`�H{/ ��-R�b�~D��Ø#o��u�s��-*t'�o��=��:#g0OM�eX���a	�2�p&.�
N7vu�`=\�j:v��[���sY�&�GF�X�{{��[c�y]J���/��F�8(�v��:Q�"�[|r�M�*Z�)�=�1X/�P��t�u(�r��5	�ZОF���u����!��V��Ŧ�G�۪/��qLv��T��4��O��=�)Qj�:���g;�3r�#��ၷ����W���ސj.Dwj3��;s"94���¨_Q�6jҦ>����P�Y8V�����Ȳ���(����C���[M�$U��0N[,)����X��A����}r�gw,-$񡋆;�սr�3{ʆ����]���~Y�}N�2�4�����"Ź$��I^�JZ���We�1�����6Ha�W&���K��,ӛ���|J�P�B�X���ґ�����e����44���c��6�"�1�1�#;���@�E4���҈!(޽T�-Ǹ�=��G:��H9K[���@�������	��sk{��-�wΠ�&� ݝ�b{�Rn�{vjN��#s_ge��=�b�7�ژ��3w�^��MW,������s����qU��7�*k璵��h>gqwJ��,�S](ݲ���0d-u|n�'����W|4�#��Bv^��5ж++7�TGB�qӶN�r��v
+�i��7N�܎��R�����ld#�i1y�tӽ��-��˼�wWc�"���RU���9׬��um��U����j`�::�O���m�ܥ��Q�YHe�LN��V,E�p�e�ɜA����Y�iR��Ԇ��kZִ+3Y-�y�F����ڎ�J����[��=;��g�jkjF�c��AeA2�'�f7��n��K�s{7VS�VC���r�P7 �az1�ķ�z���|�Ɵ�/�9�E*�\o��-���Ao�]-PH�m���Ʋ�����.����c*����zF�[��䤸�ޭ�����:�c���E��=E��YG�|(�A�Mg����f�C��8���J�[]+�V#�7�Yj=�M�5�[zv�+�Nw5]��J}\.���d�һ�;���� �/).�Yx�v�޷j�dh�+�Ծ�qk�5<��K�) u�^�PМ����.~���RZ�uoF�y\+&�;:�F��g�]�%:o��[Ԯ8��Pb*uYƻ5�B�mG{^E���k�Ta2j�{ʄڰ��9��K��&]Jެ�(W#�Q���7/$z"�]�3;��Cn�jxK4���Yn�4Ե},e�r�҇m��˩S�i���&���5��=r�3*.�ښ��69�E]D6v���3�0�I��3�������m�ͪ�ǏU��7y��Y�ʨP�[��N�^�!c� ������e^]1*sj�N��t�,,��sZ�!Zt	�>���	෯*�Ͷ�2:��X�<�ڻ�7+(7چq�8�F�j���,��1��VQ����5�c,\�-�@<��0Vp@B�o8Dt�u)q���gb���7��o���ܤG{M��c÷+�j��wwu��31�OU��*�z[��٥��T��亦c/&pݮ�nwa�z�g
�S��G����h_���Vvљ'A�*�f#z�&���Y�����Q�f�fU�����Oxt�luo�4��V�*qp�)
/U��BwC�i*ߥ˞��TPb�b:�o7Q���浕��4*nOz�ue���ӈ[�9�dIl��jA%��&}4�-U���@,qUz#�\������
N��V��. �Xы���RR�V���j�Q��"�ic���M�q=Yخ�N�����[�b�^�B�|�Z��֊ �����ǘ��,��֮Ӧ�.y��R�jV�B���:VW�i;M��0"�9}n���XvAO�B��+���㥴ᄁ��o����>���Ȯ�!1ZY*���-q�i���X��}���${B�O=Qm
c8b)+��[��9O{�*�*-���)jM���0-�/��K���	n$�m����Z�up�Cp)ǯn,j���)��o)Q�:�+΢�J�tU���|�3k���t(Qw�)Z��z/��d���u}�ѤvQ��Y���vV�����>��Ź ;�����k�\Uǻ8�٫ΙF���$J|�(r��%���b�X����V���8�
+�I�}�s��|hV
`�d��Q�����R���ke����搮�rL_pj�:��{ʍh�ﰒ�$ƯP�p���6�ojR���m%Lh}�i��5��Bn���-�v;py��N��%�se��n�
�؎��WP�*���T闻�ԏ�:�7��y�j�
T��������:r��˽��S�%�Ϧ���H��������rj�x<���Q�:�A���I�òHc����S*d鍜�t:��!�bb�9�1��e�i�'�[����S6�m���70�1\;w^L����ި-sM�/�U[�9B�ք�a��%���Ñ�9��b$�k�yC����Q̻�4Pf�ٜf�Ԭ�3�62�[7"�3;�	�U�("�Y\`8"�F��ob�D!���<O�L�er���:��B����t;/8aU��F��ʷ���9KE
t5ힺ�cU�]�PB+lh2p	����l躶�)���뷊����6�V*_�`*�[�<�ۈ����X��)`%��x:vN��t\����âé�2�I׃x'[��s�6؜��%�;-k�w�ƼND���eM}Dj�o��{�v�e�:%�B���
��oe�R�d�1��Jژ勻įo�t�X�����%pv�$��V���;|%�:�ky�y�4.�8�`����if�K���B'=��c�W�+~[m�u�uc�9�5�G��F�B�]u�����#x�g�Ύuvq�ƘƊ2�������R�|��y�x:��k���A�է5B��cU���7a��l�c���u<GgR%5���;�
I|��\�ҫ�#��^	F�]s�2tYۮ�rwX�N�a|�u��T�����QOb=��>뤬��;V�䫃{^��S���2Pk�t�mG*[=/�1��&��-�b��y�<����s]E����4�����<C�l�����Ά�S��6f�Y�o����O7Q��E�l�(�n%�2(��[A����'.D�-�}����\�#�2�����[ޅ���s�be�[���-�
@�eIp����ֹ	l�:ؘgp��q���]����8��y9m���[��;p�r�N�ݴ��i#x�Vs)��XM��']-�ա=ax�դ!G7��p���P*��n`���	�Ӝ���\� �](�U�c��� ������[�-4(���^�y�*�(���qAA���~�(|mNvssjf�5r3�]:�oH�Q뛕�W]I' �!k���\����
`�9Hغ꺵�'81�	U�h���kS�ˤ��X��'z��C2��R�Ɏ��$��q�s��hep�Ħ����rY�(V�U���A[���K���=�2�����i+u}�b�*�!qO�i�37�򬘅�e`-��tv���Ls�Y+�Wu]���Go�Y�X�H�[�`��g}n�ʷM޲F$��,�J�f�:Ű��;V2�q���օ̞�k0�+�G2w��pO�AKQi 
�,��A��[;�;��ҨN�6Q��7�����d�8sp�f���yPaNł�li�h�S}��)�"�]O�43��gG�+��TU�I�������X�p;@�v�/
V�u�e �1���V��͟G�B�]a��2��Yo�C]�]YSww��p|.��,�7���s�QOr��[|Zƪ���!��*�x:8�Dͣb���LU�;��̰.�o7!��sE�-��q�ݮ�$�9�գy�C9�[�
N��	���ǡn5�RCƬlM�xsP�=��6��E��l5d���=`�Z�T��r���"��ۦt�c�t�����\:crE�ƎCw8���P�4�O4�m�'S���[�x���p�Ky�}i>��;�l>v�e2n��td��gf�GgV��2�CYv������:�D�D���T��St.�����H7����ʜt���Ktyd<���� MV�*�f����6�w4�1,��i{�=�Y[4��ؾ��T�7A��w=Co�[���SU�V$�^������r��RLn���[�� y���j�iP�j@�9�)K�j��|ߓ�{��y�鹚i)8���Zhi��<�ǻն"BI�������!����K9��'-z8[S���76ƌ�r�N��˅s�]fj=ى鈭� �CX�nw:��dj���/z���˾�byy(iX�a��q�3���,\�m�aK�t�ڀ߲��.���c�VAU������ܬ��Swt6p��^��'#mm�ww��������	&����׻�7���Ё5�x2�R�|@�p3�J*��$�uN�p�2�F�7B��L[�n*���5��&�<���%��$r�V�4������j���F�6���NU�H�u#5��NA���8�-�'�[���Mz�z\�1�ɇ��!-�������A�*.�*��w�
�C<yWd[����a�Ceofi�}C���>ڒ�W�&ǁ���|ه����[(�0|�f���3�¬�r�.nj�CT�����X�Y���Mո%�ۘ�o�����Wb��(���^#wW�r���t�8�9C�pՙɒ�^�v�ūz�A�/W&nm��5��x��A'�Ok�X�5�"���M.ʚ�Ub�z�N6lUg��5�0�t)伣�\�E��A���yB�>��nt������
X�r���8��l�a��
:`yO&	��nm����Ӹm��6�ѭ}�����@3ݻ�&b��Q�A"_�^��T/���A�E��v����8�n|�j�R]�7yt�����ӳ6���4�[.�e�MfK1b�5hc���j�U�i�o{��h��J����SFlgzt��U���c����ޑ����ק�4��c��uXC:Cu��Ui�m�[����œ��@潼va�Xl���}�N��9�/�S�s�,#����Y3"ə�xeeIy�V��24����]2�l[�&KG$f%̳��D���n�Y��14�=�A�D]��<]4z�v܍��
�3�b���E.o5� b���#g�����U�A�N��"�x�9��5���0�آ���o5R����Ue���W����u3�?�Z�pP��a����l@�e8*���B�J�*-�: �o��C�-Ot�te̕qT���ߺ)H-p>9 ��ٸ���!m�}�<�����&�b�o��v�PJz�̫&��2#�E�#W#��K��7Sxsu����ꮬQC�J�8��S����_N@[o5�<:�M�X��`���6���Kg�\Ĩ�j|�W�;̀%��X�i�p�3f��wT[��걎����Аwo+)�ϮjC��'ܨ�yΈ2�<' ]������b�>��n�����+�Z);L4�>�s(�`�
uxOme+\2^��:̢�����e0It:��bݵ���JK�{��H;�p��s��\*�5T�5wG2�h[����h��s,�݂�}�ڻ�W5���wG�j�lLs��w��u�tƥ*C��,�1����W%5\��b��y`��'�41�bs�`,a�-�y�:�M�[7���w]i��d��jͼY��&*ZO�h�f�ja�g�]ؓ�����IAΖ�T�l�֠�Lj�V��v�`�a�`m$����*�a�}-�;��5忱�э�Y-����-�Lcv.�QJ�M����v(��]e元lYd$�T��|���"��aF�nC���ޞM�|���t_o	y�\���n�� �-��mRo0�g�szClo���KT	����]��Tݕ��%��=�%�<*�ҥO��@Z'F��%��8�;�jl��=t��Y�j��y�t:R�M���*�T9E�6l�Ҏ�ҟg��ޏ�=��q���i��2R׍�-���G,�y�KU�]�P���[.��u!��V�U᱕�X�t��_6��ZѦd�I!�S+�j�4����Ay	�-��Z��h��;��:�r��k�"�A2�֕�����[ -$��d� {������voaT���
��`����i�Nuz]@�P�9=���Fԗ�o&���+�s�c�W�V�^�OA#xN^p4��u�,e]�̪eH�(ƾe,2��u:+��K��#8b�NN��Z�����W��S��V���E�}u���=FZ� E�5[����;�fb��� _R��pI�w_bYC���I����g9*�s��:��S�/n�M��7���6j�#ovh6 8�\�Ѳ���㬷��[]@r*��!B�s*�\��ˌ'l��S;�G۫%�ӗsue�lVnR��o�V�8h�}� �`���f #��eJ]��\Y�Ot�w�v�`�R�{���⳱ә���t]�8�X�d���er���:&�9�Pј��Q��j](��[{��[�s�:d�&CQ4����m����W�����1G�ەC� rb�W$\�C>H����i�u����=� �K˺�.��kʘ�����ϯ9�;�7h�[)f�i��n��s�Z���e�P�Jh8�����%MS�e�Mم�r�FM%隀}o\�p�N�Q�CV��@4�Z��\������W>QL�a}tv��x
��9�R���6@��ɽU�� �hК��B��3!��n��G�b�ln�����D�P�ガr^DJ�U�4���� �M���G*U��P���yv;)Rޒhݵ�+���ڼ��`�=�3����jI[k����NH־�wg�A��}B�(3�/EK#���\;�8)X�ge���[�ۢ�+�n6֓:���@Iε��-�־�����;h��x�+n=T:���D���rc1�#sl��=��o���Üwu�oN�4��;��ӣޤ��ʚ�'����_u����Y��7�)Ľ��N�����u�^������S�F:	K�m�:���]���=qi=7[ �����J��H� �ef�`]Z�=�̃Bԛ+�jf ���܍];L+1����&���Z1N��į:S��}�� �8�m#�^�5��5Z&w:�Ǒ�]�$;,�d��N\vd��-<ڙ��@��Zr�u�GR2>�@hԀ8"(`鉴r5���v%�Jܐ��7sj�
a�۲k`�E�n� �j�=?=}&�5 �$���UwMUګ&�$k��gmN�4cЀ%w!��:�H�d!��ru��b��%k8��Z4[���44�#Y���0Lq�6�ٷ��}�C��I�w��t������$4l�^�u:�q���w�q�sFc��4l������0z��n�&-n.��lޱ�x����v撟uk�e
6��8f ��q�.��FzGyҫj^����#�8"������;#g>�h�*�vi�$Ko��n�m�+�\Mv��miۛQ�f���a�Y�(hݽt���-�>�v�K���܎��8�,� lCCC����f�	�LJRެ�N���i՗���i��Τ\2���.ʴ�`���.�$����r� W�t��:����-�iq�F:�:�}ղq:�K���.�> ���g/�2���H��{�ܖ����'�^֪/v�e�O�t�7z�N�J�	��jsQ���/�8ʾ�2�����G+�#��&�p�7$B�	�:=�"�۝���G�2���qi�96�tQ��P��{N(�;���d冏�J#�:F]�I�ʷe��(�KR�<�F���o�:Čh�Y�������7UK-��u_P��t^WO��e�t��}b�&����Sd.���՚�]�ŕ��O�l
Od�q�Sy�:��sf���V
�n�>��=��>�����*���<:��б�oa=�x�hb�h=l��Vo�33��Ȭ46��m9Z�QO��f>�;z19�g���X� 3�8Y�
u�:+nn�VD�<ѻ��Q݀ەv�A�l�W#�n�m���A ���+�tr����|��aNt�v�R,�
j��&ŝMc�7+{]L�`Ч�����\{���������U�� ���s��/wMr���W^��!�ó,�b��:p�4��T2�''}e]�$���Eu,pOn]^�y�ӳ�8�	���i#t>P�Ԛ�fu,��2Hó���-�ui��ӫF�����KV��jƃ��@;��LԺ^��&)<WƢè�e�b꺹t&�,�Mn�W����49r�ɐ�3�v��i���󺰊<��[�	}���^터q�˫Ŝ5�%�����]�e�����O�R�0-��匝�+j����1�m6�앏��w]�IWj���q�c(n�}ͫ���_�Yv�z�+���Q��T_Mz��|�2[u.j�����V�9f;��et��������[��/��E}���������Ӄ���K)+��͗Ƒ��vn����O|�v�1]fr�X�����)֊cf��-���Fi�c�V�	��$ew=���O�N��ޙ�=��*V���!�j�ƷZ����64%�C}�6��M�;�f�VtC�f��tc�h�щq�-%�ZXGǻ>4�:�i1�plNǴ\��.�V�3�k��1�˶k�0:�z�����G7i�l�X�>��e�i��0����}�2�Vqae������bY\�8�E�`�WbPͤ�Wλ��,����N"�
�ͪ7�1ܔ�,5ۋivFS���vZ�p���dY��E^
	V]���^<rM$����MI+y����9{�"�:��Y���L��k츌�-T��w�Z�D��\�W4:�{)����ZU��%���^M{ ɠJ:Ƅ�R�+��+ݻ��ěk\!.L��
]��Ԧ�Rsw��`�ғ�^X�5�`��6�qf-÷���=z=�1�n�a���}�i�E�����"�K��W\����t���T5oa�}z�����ܽ��f+H��*蜤��S�t�5%�k��ݮ�Ӝ���(_#���f�9m�yһ��s�i��J}ב�j}Hd�X�/�ʲ���l�w�/�.�^�v�]��T{������*t垏p�7K(s4o�WW{��l I�gl�|����`%�!�����1�0�c�5ޭ�o�Z��à$"�+T"�*5�.s4�4 ���2�yuJ�X:[!p?`�J�MČ�>K�s�X똨W���)�O4� <:�>��u���'�g����Ѵ�N��0�+�`VD3X �� n�Y�e�o�P�jv������&a!eZ���L��R78�{܇X�6�WMuk0K��$���C�CI�W>X�C1��M������SF̠e�F�ƨ������/g��v�����3��ɉn\��'M�5��d:�GgcR�q�g�-�d�{K{��(�.���n�߮U�m ��ut
�ztU���v�vFp�9�n-�pˈu��D��(�Վ=�umUޭ�{W�����ƪ4�b��h�DoJ� ى��|�l��O_V@�bZ�.�V.f�`�7��6���[�tO���ۚ��s$�ޤ�7Z;w4p������tP5�J��9����c)��W�7pnq��S�5_X��*}�+���sX*�ڷD�c�����F�fl�
?eq�{b�;�������-��n
�����l��rF��|h��Vv�4����{�8��/n��5��s�������$�յ#2�^j(��\�ayG�@2������F���neI�j�\��n�=�lHWVXZx�]X�:=�u�`����F�F*�8u]Eg���lV���3@��	+�_3�#-�6w�z�l�V�Q���5Ca�	d��yړ�Sw[�[hU�юK/��4�뉱�'�#�ߏ1�b;wa��N�X�]m�f�X�8NB� 0v����Z�XWw{���r�Ȟ���ʌ�}e�0��꼭�M�x�L�,��=C15�ʄ��f40gnGgr��S��Q낹:MV���E�J��Ü'�v&��͵X-j�fS�w�t�
b@`��u6����Y7Eʙ$7��g��6�i�.Ց�/�w>Jro�r��۴�'g��
�I���2UGx[��@kG0tV�۵�*]ۻ3C%YK��4�XH�r�XO�5$)�8J�;9]�t�M����={��e��V.C�1LxH��[WۓW��������I�G��n���W@4{
��*�T��:w	����[�k���%nv`6.m�Ne.�m��AAeäX�ȁ����98LMH��q���}º�D�uE�37�'rh\MT�<,��r�b�N���b'n�*:���__:��#����Pb��u1�+ �p�MU��]�TLT���_34e���)QYy��pW�`1�n��;l��a���w:�"]Z�V)�b�;���q����q�}�nىǷå=(�i�[�M��]k��.��وu7��G���A�z�3Wnf���Hҳ�+�:�\�S������vrq_LX;gp2�T�Z�ch�z����ͮ57��\�cp_��8��m� ��ڲ��1�x��զ�f,%�|���a���g�zVM�q+��YW����f��P۝If-��
�:�A�vd�ܝ��KF����6�γ���<z��69����3\xm�t3D���ɭJoK&c��jw�bg6�f�9U�Zs�^�y+:���x �R�z���{�(g.f�ʻ[��=Q�����7{�	��͛�Q�7@���޺�n[<�GD`�V�|�f�����=�>�5�A��,�}s��z���Y�dKNs��]v@�����#�ټ�s�LJ�@�2c��C��
��g����m�-	�u�b�(q�>�dib�`�Y{8�p���H�8m!L���e+�TҔ�H�5�y��+̸� �0�)6G.��S��b��3w�s�wP�;���*�v�
������0�q�J�)WR�MT�2�#�����=Lj�s�$�����T<[�A�v��]��K�U��\:���o9�tc��@�q�ϰ���I�o���Pp�m�i�͝����օ����4���m:h]�ŉ�̽���CG`�ض�-%.9,.��H�i-�Z2lљ��	3Wa�Ԛ�z���,^��CH��b�����Bd�ݭ �2�����Q�][.�1��'�`���X�5o]��7v��m���Q�'�z����&��?V\����~���H�:��'�ۼ ���XU�Ud���e�*#�]�zAÂAon�LXwRW�^U�W�z����So6	'kE	�le�.-\�e�^Av�:)��Z�}����S)��
�[9�W�f��=/X9$�<����ӫ��ц�;s���Ґ�b�J
�	q7�3|�
�7����ق����OS�+��k睻;%�m�И,h3���d㫇����nF�Ğ��j�P�%��8���dr�[���C�϶�o��#q��U.������r�S�nS���=���/`tcb���0Eq��D/S���a�sOn�Z�JV���S�R2�.�s�6�T�j3�S*����s�Qθ����Qk;��آ����v�^�R]���x���ע>U8�ˁu�_'����vn�2@(f�1Wr���J����v����p���4�sL�7wӕ1v���	��.5�4U w��@��+Eq���:T���YcRL0�)R����]qVE����x��5u�f�E��w6�%I�^T������^̮/%��Z<�]���2�`f���6Uݾ/%����V�1��r��V�f��3A��$�aJB��B�Jw���Z�t�F�A�ml�9�ݬ��9�7v+9<4>�f��Di�]:�6PX2�A�d�,K�qr�3ҷ�������DEERU����["#*J�(��"��1�AAJ�X���)ZV,*�*�eb�,UPXڡe�QATY�
Kh���Q#mQV*(�UQ[h1Q�V**��("����V�X"���bȢ��(��
1���1�F�
�"0��QALh��P��E�A�T���+X[dX*Ȣ�)aTDE ��-B� �����QcX�Ɖ,TdX)RX�0QT�c*,XE��TU$�R"�QR(�Y�)TT����
���`���Z�YP1�m��)��0F,��H�Ar���
��IP"�¢�d���E��%b��eLs+�11�P+�)b�D�IP*�P�-!X4� |1p�f���`���<��GY[ίa��d�Z�k��g:�o�Y�!f��f�j�{&S�yS�.
�>a�|��.lq�2��JM�w���ۯ��K�Y� ��rj�O�MfF�����fY(TȁnS�n�<��,��Aw,� n���v�(/�p�Q_p�R���ɨޕ��l���".r��s����Zg�q��*����뀬�Wէ�ۅp�A�꥿����5�
�t�v�{�����t/��_.�U�p��g��ɳ� �*J�
Lf��6���؝��N��CD8�U����@Lr���}���_�I�P�*�_�2�=yR���u{t<s��3���n�������7$7y\(o�����������c��%^��r�ݩ���Rz|�Y�]7��lW9�τ�+\����2o�b���w�8��`��(�L��X�e��碾��<r��c��W����]��ءc�����<��XA�-q*�^�{���_-xw�zO�8$ �fP��,�!���0�����3��5Vq��G%O�a��2�ߞLp��k�e���
��\9�GzR���*�Yt����s����]��&�So��4�A[�ﮭ����ʓypΐ��Yt�����A��EJ��h���۰�2�¾WWm�a�Ph鏎#'fR4�-=�L�j֣}��p\�����M;���mpu�[��.�IG9�w`�dX��1�sy��h��d#�n���J�_J�U²u.e�@f�{�Q�!��v�on��V#��jut�
�h�m5_τ�zݼ�2c��e�qzgL����e!�Ō$����66�5�����Yq�E|�ݤu��EE��Kw3"�#��N,��K^e߾j��Վ�B!#��B�+i��%#����TCi\Uê��[���ڤЪ�;[ӷ,�[��ٻ}�M S�~��U�r�g�p�N��	�h*��HK�V��y�#�����s�~qx��rT܁�ڲM7��h4T�ĺ�F�n͋�׊%�mtf�su�u�(`r<�����n~|n%] ��&��{	���B�[3.,GQo;os��}J$S��6M@�t���a�'VK�1_6�DW�v��͂5��v��A���T�ձۅ9��U�a�y0��n��j�����r�Ĥ� f�QBD�c͋͂bS��m΍	�	�$�7�2GY���j�)��.;�l_@�r����C���,OYи��0�F��&�V�}.R�
���<�o�5�l����	���ѿ7���Tþų#5�7�� 7*�[��=Q��@�f6`i�ы9nү��V�kS�ӂ1��МX��dW@�34��i/ ���ԺV`|��L���ܦWEw�Ý4����^U�]Æ����#��������A)Or���gզx���5�� =g���:�Z�B��p�ʥ�z{lk��B4Ɯ�N��p�֥�����ܾp��t���`z".�\����sP���~����n�ԟ+����*�/���:L�;�i�o�o���GqߥM��T�[o��铛�S^��hW���WX֎���[���j%��aq=��Qg�8M�e�Zx@׊��uֳK����NAt,���h�8�c���.���VW({�̭��y5ƹ�CLk�RF�D� �����̭]Q(�}p���8�X����(O�v�徖8�!���vK. ]:JAf!#���+��6��&}y��s���w~��q�ӛ�ё+���H��$G#q�'�U#~M�C�P wb��u �/i��fiً]�u`N�c件t��run��f4G
�ˡ�c� L)D�H�;&&9���`2Yu�˺g�Խں�˴����'hs�T���NeɈ���x �c�e�����9b��RBq=�:k��<�4Ak�+#s�S�4v�*9��9�w`����)��kB��b��'"/�<���:r�Uʼ�W]M�������k
y�Qk��q�ԯ���y|��r���͉_'�Ɋޘ���X��4��"�Z��9t%M���>��k)w!�ݝ4��y�m�6�o���U%�>�:�~ط;&�2P�V������S7�ԏc�;�[9��2���m�� �
������7�Ɠ�Aʗ[Wx{��]�HJ��͛^�B�'j�$��~�P�����h�za��XXH���A�Q[Řx~ԍM�]��u~�w�Ժ�܈�����r(����og�k(�|MXվ-1[�g�%��"���e���5K�T��0�S4�a��7�D��+���J�1�T[\&���q9�n{���V'�iW�a`W�X�T�O>0��͆��v5�Q�9b�@�zj:X5�B��1[�J�����u�>��}Ҏqb�U#���p��A��7�ݵC&�,����F��� �:G�yJ�����>�Ub���D��끬�<~��;!˚�uM蹼�y'xjy���+��p�y\�Z�<���UO�xTǶ��/avL)3�����IIì�&�f����xA�g=7G���U�Ws��IHt��������K�4����j����;sE�t��zf-�s(�ޜy�8�v���k,��ʛ���
�Q<[��މ	�1R�ip6,Y+o����A7;�m�T�no3�1�TiB�Lɔy!'d���a��7ҷ�;n����.w��a��W�xh��'ih)�p}a�NP��5�xm=�b��j@�̇Sm����T�G�1ip��8S�[L+�꿥��xtB{\T湀9�]�L"��-�+�3�s�s)fi
�޲����4+9J��e���L�#a���]�1�沀i5x�{wU�\�b ZQ <4���մoL1��a؄���}V�X��U�H;-F���MghN
 �Q��L1�Pg�6�H�s�#��x�U�e;)��K}��Y�+�;��"��f�Dʉyw���$��Q=r��^�5�s��U�����_o����<��f_l���Ϲ����S��̚����*�/���Y��	��_w�?/-�+�do�\��,�]���������؅}Q�.>nN��١������;wN��J���l7�"b�50������ C_gS�Sԑ7��j�m�����w�{��B��w�Q�O 8*��[p�+�$�w�U�m�NWJ<��ūX�l���g(�Ζ�o���V.�<���99(�c��+���͸�X���h�WV�Ms���4��ӣ��l�9��`oKS� �j�ˎ��p�F�_]+B9�8�W�~�W����w*�����g�C0� g]k�?N��z�OȺ��Im�!�83y�x�b�yoÅ�h_*z��p��3�ί��
�(��=�#�ոy��+�o�Dܣ�4�K�ֺ�o�a����Q�P�o��͐$ ��H/Ƹ�K:�צ5�ȹ0�=3�G�r�Q�\N�x)�W��Q��F�h�w� ���
�K��qN�^�]g.j��v־����C�8�TC����t�pḡ{M�/�ʷ_ð��
%Q�4c�
{o�S���Y�RuJ�5g�[��ȅntPz�����q�f"�ǐ����\� cy�FZ��>c�eCS=&4���m��Yq�^[���A�q����'����v�j��e�^f���(C��g6e#ݢ~b[��:��9b�w[��������f��H�2�����(1��;�0��G�Ͷ��z&�,����v:gp�Ts���o��>�b�.q'"%e��"��8����.u<���
!��S��D:x�7��L
��?�,�<�Y�k���>�W������)�n5 Z�'=��ե)S��m����8��#�r��u+�bY�+�_PZ�ɕ%]E},��]JYZ� �ZvFu�utr�.P679Q�ʁ�(���v��fp��Ac�2��c��u�C,�5�>�?Sg��cmШʄ����n~|n'VX�B]V�'l�k����j�Ҽ�0��n�"�s�a'
���6MGA�(;N��/��)���H�����WDP�>*Y�����r����~�{���a����u��L �%L0�+$�9��Y�J�2�&����BѾW�l�	�΁�{\�^�����A�;z��e9D�YN���trVb�3��ۨ��룅׌�rí�٧D�3�k��y+e�tR�b��<.�|v��ٲ湭�؀Ou�&���{��_p^��O�
��f|�X!�:=
��pJ�J��;juRY��pr���(C�꯲�;`��iP,f���_��(�#�������ǉ�F�鏷�37<��8`w3��v��Q=QAX�h�p�����a�\c)����X��0a;��(A�Fis2����z0�
���E<�;A�ŋ��/�\',m�
l^s��uF��~�-Y��
��:�C�:&�<k��q89��#j#����'P�>yK�U<:�U��^��4o^��{.&q$��E[�����^����5��$õ�X�K����{��pp���M�����Q�ڦ�%mj���*n���Y���2����V��;�λKEVPC�GW�@_f���ٺӻO��Uvѽ�-�����ݛ�{�jyqB�&�XJ@��d��BG�����\n�7��Ź�˶�t��z���|��"�!�_[��V��E��THP K'iQ���y{Mny`����l��_��H�<�l�n���t�n�h���vu�tJ���c�ۼ������2�e�t�:
%�ٓ0*�o�8!��<#��*sr�L���suD�K%Wm�r�[ï)����%9��Yd�E.��X����r�`��ul�j�S�&,y��r�s��lf�8���Wz��v6��;u�o0��yb.�1�;��a�'b�HȆ7'_3'{���wy�^+q�V]�D �<b��7.��n3rB��àn��,+$.=g6���:;#F\���8V�Wx�gL�<\O�7UP��8n=�0���0��ޛ�N�z�T��`���{Ow�fL����*�Rw��&��8{ke������"���Žk�n�#��8|���CO���Ib��.��u9k�b*��:}��\k���wh���r��>�4�
/���{�
��)��3������ݼ�ޡ��T.x{���z�tN\{�YI�q&�lv)c��>%Q���4x^��o���ݩ~�`�+�f8����Nx[w�K|]�K��"uk�M��}�v�V��/&X�{�6�vz�xEU����1QX�t7�J� ���1�Q��9��Q�V	��0��+L�7�F�U��ϑ�+RU�.����8�ȭ��\
�e��k�F�P��F�YT���su�{b��}a���vlL�!:Pa�4gJw����d�\h4.�k�H/��F���I,4rˎ�R�v>��u𜭑[9 ��V�S�x>5�W���5r;i������&��y����ʣ�N�9D1�n#��t�Ϻ�q��Q�l��1Ixe9(9��î��S[�̜B�gf.!.�
��ѩ:H�����B08���;.J₃�
��(խK�n	e¡I�J��l�p��W��MG�cQ��O*5���2lDu�J)�{un�Sy`�p,��l���n�GC���\q����ʚQ�@�qp��Gv�����;����dC�p�����&@Zm�K�h��a���P�$�����:�Jr�7'�Υ5�x�)P� u7�Ȥ���~�"7>�x��5v�C�F���&�:i47S���i��s�
����Ymb�Cd;W�!�T�Jw��>��*a�ֆR@eu�B�T��ifʹs���{fr�)�,K�J��Z7�v;���RV��T�)�k�}���Fu׽VF��6��2�%I�}�������ӖM�����y�|�zD]Jc���)�J���;����-���*�7����V	=yP�"B�y�uйx2M�&�9iW��YН��0�f\wK;��y�x\>��7�{w+�n j
��n��Vwc[=�|���FYN���L��t '���9��
�tk���l8k��S�9*�(��'p��\I�S�W�^�,`�4s��":Xľ�2�b�X5���ϖ�C�wp�_�s:����f+��>Gl�%�A\����ҫ�z��L��,�p�&�m�0�T皊�ʖ�`�jo���1��Dt�K��Hh�_I�1���ʡ��-������ղ���1���"4�/�_=5�P�o�W�@ �'���pS=+�ҹ8��-��+�ǽܳk"�D����ua�,v��2�ߞLp�F��_Ѫ�#ג�dfht!��n�Z�u�Ȅ���7�d��W֪�v�<���Kg3���V���8F���u�oc�� ,���Ѣa�&�2��]dD·Z(\CM_��Oq܂�>��ފz]U����3��`멦�Dm��6�]����lXa���/.�_�M� +�n8�p�H�oU@��-��E�.��qXװ3M��K:ا��C����+]�ق�q�U�S/T�L��4�{i�N��3��gn��5�e�˳
���5�lp;������g�=�yާ6���Ԣ�TYv�s)>�Fԧ�n�BM:��.]��$�v��L���`�����Ȋ͸;�;�����:v<#�u]�MЋ���N�c]�¡�ڦ%�8˦��3�M��(�P�,e9O���u���7Vbg��6dU����i,�w]�,k�ĴM���M�g�h��ѝV{n�V��}���Aٶ���i�i��w�欇qm�_K�j[���E:��Ho�uȲ�vuaa�`bY�Yqg@���7Sj���)��7�y�J�3�%j�.m����o��]��4򷓬8i� Fv)6�qP�%A�lQ�;^e>���"�]�{���6������l����]oZw������5=5�31��ɴ.����S��k+*��Wp�/�/Oo����k Z�P�=�X�8���CN�:����+��U�
�p�\��z�t�pk�p
ݦ��G�n�[YK�ۀ:uXl��1��c��W�Wl,wgc��� H�#ndȇ\Op�k!��Z.�����9׬
�g �K>Q��M>Ig]�R�l�~'�/^A�^$����$wF��Ԣ���	�l���fY5˱m��N����f[�S�Վ�CUv۳��c�O"��κ�[���S^6H^WF@�l��j�n<��E[Ұ<��,k�2�V\�v�
�ڶg\S��'w|]��Hj�I��qÂ��V��6��о��M�j.�6�gV<ۥ`r<����m�3�%\�f�d����c�{X��d���a�`�M���ɻ����6�
_�h� vz�[k��js���F��%��*}s��}K0�Ry}\Ф����	b��_v�]��n�k��ӽ� G�Jl�َ�u��U�:��n"�l��]R��q;φk�M��� @.�#	�Ө
����5��s�J��i��g��4 09�rWN���D�%d��/�h�~��+=践�5��ʓZ�ڵ'�����r��;U���Vi�)���R
����{����M�N�E����9*�3_JY�G&�F���t[˥^�]pq�S'�M:�E���o.�*9��N���hzw/�9���|�/yǣ@�Yuj��;�ĺ��8%�kE�p�ϻ�^�aX]��A�]i{7gL��ݚV�e�Ei��WKt��ˆ��X�nƛ����ޱ�'K���A��"Z:�܉�]¯x�f<���X�O/(�:${n��;�q����ꫴ7�,2�K��7�O���Vc�m,�L�-N�g����A.�-ݍ�	�5��A�d���u1`Qމ�t�:�6�*���O�к]����7��V��uę=K|%b[S�&)���ƺv��k ��b�E{h�3* (�
E��DD2�X��1q!QE�P�dE��"����E�E��E���dE���b�X
G)(��� �YmV
���J�(��ET`���a��0�,F�UPP�,��A��U�"Ȣ�j)" �X�X+*�b��aPcXT��Qd��LLH�E���	X�")(��Ab" ,E�Kl-���U�J��EX
AdX��$X�V�XVȢ"�H(E�(1�Ĭ1*V���l���Q
�$U�T�$�5�!���X���",R((Z��(����(�X��V�`��Pb(*�P+%c��,� .2�X.'�ߟ��Ý��㚕mL�/8X��(���@-v�x���ͭս����2���1�VR���Y�w����4�T����]I��s��+����L�}�|�6�U7l������C`T8�M&��&$ܧ��N!�C���iP��N���H?�>C㟳�g�*��9�:�o��"�eg�z�FMn�מ�Dp���;�Ȥ�
�̗g����L��;��v�Y�,*N2�N��EX
N'��;`VW�z�a�x��ܡ��f!�z��36�U'YEz`0/ɃYS>�����g!/�b!�t��6��?$�O9���I�1�'��<I��������6��6sY<Փ���f q+�%G�ȲbN!{f�)�
��j�{d��>���byf2�ew{�=D!�p�p�Lz\�P1�I��d�P�AV�=M$�����o���x�?v��4�YYǝ�����!�����%�&3S.����>�;d���o60{=oGl��U��J��C�|D}��e�|���`:���m�������i���y3�7i���l�0�i1�H/�{�@D�~f3�s�I��*Og��L11��Y�b�!� �f�/��N=��b�Coc���8�5M��������f՟�T&�5�ԕ�4ɉ�`uCԗ-Cg�d4��W��g;�<���:��s��a^�$y;̓I=eT��y�v(��
�
�C+T�s�ߒ�)��n�~�5��c%q�^��=B��z�Ɉxj��f!�y5��
��l����H/� ���1��Si>B�;C���)8�aX^s1�I�*{>�M�ۜ�|�C��z��y|�צ��;�߽��R�d����Y�J�H]Ͼ��+6���ϐ�P�&>0�T4�|�OS�{��8�󏟬;��f����OP�<=��uC�B#7�DxA|G�ET_��Պ&ݿ_y�����4�a�b��g�/Ԙ�;ܞ$�L���1�T��5�+Y������&2~qY6e1'���L|5� i$���������;[a|Cs۴�P��B��C�e���\�oW��k��&���d��j���{���<gXbc'��"��1=C�~�sĂ�|§y���Av��u�P��RVM�_HbJ�O̙�'��\�7�&$�
Υ�?���,s�g�Y�V��E�M�����v�ͪ;7�����Xϟ�S����fߺ|�v�,��>ۋ(����5s�Api�8���ś|ю��j2++/gAٱ�ە�)&�8Z��T��m�]�B��\u�����O���!�̠z�� �>��:��M��<�Ρ�����9����� x~�m!���O�K�5�3��GP� �{���'�c�W��?$�`O��(�׻��������'�I_��
݇�'��1'��q���ٴ��|����'��a�O�M�̇�q��~g�y�a�&�Xz�<I}������~߼�����3��_̊T�B���/Y>Lgɤٻ6�Ԭ����O_�c��'���^Xl������}�v�Rb���d�Y�����P��'�$����_>���ޣ1{�|���/n���hg�Cĕ�|�5�i ��Ô�N;f$���D��M��8�Z������g�11Ԙϙ�3�����E ����<��=CĂ�����׾�o{4=�:�WO�.R}���1�{�S��>I_����IP�~Iy�膒q
Ι��I�sbO���Vx�s)�����*�5a�4�Pէ��>a\a��g|�ì���>�}��©�b��=��p�ݡ�N����$:�z�g�q8�2u�� �׉3����O�Tߝ�\d�&������6��Rq6Zc
¼��i�j�& q+��冑f�*M��~������7�<�o~��kއ��z�`*��_��3����������SĂ͡�k\I����u�@�*O���{�i���!�����x��Y6�M3��q�LB�kb��Y�}����qQ�s������SOr=�#��1�l7��4o�4�'Z�̕�:�'̞8�o�%I�+���9�Sǌ
ϒwWO7�i �>�h��9I�L���1E'λ�jx�d�@��uy�f��w��~�W5�G_}��m1g�11;�3�8�'�������k���$�!�+4�����M�ԕ�>Om��q
��7�`8�y�u�[�`c>3�ěea׎�s��w�S��>�d;�3���D��">�����%B�^�z�4���nj�H|���8�j��H,�3��z��Ă��Xu�C�����x �f��9�<@�T��|�tx�M����&��]�bl{W��fF^�I��:�sgB��ֲ^�]]޵�42��=s�K��0��Y����ҬKv�,�0�*{{c�!9�����K���S�;���[�@m)Ǥ�rH��#:����;er9�,՘�N�k��i���8�����l*�@�;>���V��O�5��*$�J���&�ed�h��CYd���6eI�/�O��O�
��:�y?P�=M�q��a봝����ϒ����A��?aE����N�����׺����bt;���<@�V��L�=z�������Y�K���d���/?j6��'���Y>k<a��8�O�<q�5�I�+�<C���C�s����s<s�s�����B�d��4��}�i�d���i?{�J�D5��m�<g+R~��M��qgbg��3������$Cgy�P�b��>�v��C�K��u*$����s\�]g�ۭs��^~߿]vLI�*'~����Ru���d����~��n�>z��{�&��J�����ڤ�P<9��O��=a\v��?!�������x�Y�<3�ژ�'�bA��]c�w��g=ծ�W�)��P������"Gވ�&v��������Rx�)����q
�?P�+�
͟�'�+
��>��m%@��˧��VJ�w�C�o�O�����	���}�l�i�]���"�!�$������}�D?0���^$��bAO'��%t����<��1Y<J��z�I��lh|� q+7��a�i�Lz��۴6�U�Cs=��hbAyϾ��Oݱ�����o8���n�=�S��� �<eg�t���u
�2y��j�R~B��%M>�*~�Ʋg��'Ƭ�q�򓎓�WiX�C׬�8�Z�`��qgp��4x�Y�u���a�s�h�鳧M�_u{i�ԧ �<Chx�U;a�N!�I��~C�1Y���6�Ԩ|����2x��T?s_�6�'�N`i�������Cԕ���]'��c8�PѺq�T�B�O}4s�ſ��������vm'��cw����C�bk�u�&�:�N�Hq8� [�
�:ʇ���zw�!�Th��ܞ q*O����1'S�Led���/0Xs�.����IZw��oP�qU�/;�y����8�C�J����4��QeI���O����W��1&!~���d����P�6Ns�$�q1 �;�J���s�1=�Y<J��}�!�����4m�a�K;����}���HW޵�2+k;�H����2�`j�}�$*�_o�Xgo"��Q���rQ'�"ѿ���#��Z�-�"rV'�8#��'e�7x��f�jj4���靵 �M�Akdu҅i<�Q�U��;��Z��ȝ
��Gxc��i�剰e���]����!|�
���U4���57C_Rm@�_����c�Y8�E��g��=�m'P��w�ws��g�������<�iԚ~d�SL<���Cl���N4�Ǿk��k3w�77���q5s2��3���|D|*ȣ��mf��%jn�1��1�&1LH,��O|�ӈb�]M��*u�c+%x��1Y�z}�@�T:ý�x�dğ!^N�'^>�"s\��Ưn��0�o��A��/�>�͡�%ea��������Sv�YU�2UCYa�8��0�<��M`T8���<�u�4�Y�|���C����l1Ru�S��>�6��A ��f��,��Y��E�	��?%gO��S�x���bOL��+
«�'I�*~����*x�$�o�:�q��ʆ�X���'ɼ�V��_i�)�&�|��v�]m�_�{g�Ԫ`x1��E��~�YNY��'�O\I�3��iY=J͜�E$������� y;�h�%eg^$����<CĂ��^y�fRb�G�1�c&}C��@�TY:��iً�� �N<v���(Ƌ��'��|���﹞��`)<�S��>K�Cs��4I_�3t�x}@�u���g;�����U��y����1��{�kl���g��}�<O4�;��!�@���B���!����s�^o~�ּ���o�}�vP�Vt��M u*O����&$�6yt��v����P�:�sxk�%C�-�h�����AgY/ﻢ|ͪO����`I���)��,)���N�T�};J�/c(^k��������q1 �}��Vi'�c<Y1R|ʇ���4�^����c:��8����]��sJw~g�U����D�{
�����צ-���P�&���q<�>"��`���nK��}U��u���g�q�v�C�m�צv/p���ֶ�p�XsW�)��1��6Oqg����>���ſ-F+�j^�y�H�6cm���w��Ы���цҿn�^3�G/;j+&r����m`���V-Fv�t�V�ܚ��@;!��7�e�Mƥc�oGS�_9��ok�7��u����V�Mj������]��3�b���)���b�`D;]��7zX{ݥ'��x1ܡ��\�F2��o��3,�u�3Q�P�q�A���a�޻�4kpj=B	V^ooj�ս\',B�&z%:��;
e3�]��Ѯ1�����_� O��c�LS�j]�t'2����&�'�V��w;��|:Z85��iL�5);�s�7�e6��R����Y��蝢4���E;�!��fO2�~��1
�hb{����t禷|�O9ݩ�
ڝ3WY /U^˺�=9?�}�q��t�����P/ǞВ���JU٬�k&Ji�jk����+;|���ԁ��,J6)J5p
��$k���]��%"��<�Y\�c�Vs�ѝ6g�����ۇ0����`=�� "���zI(m�:��_�(��sQَ�!8���V����l�ՙ��Z[�g���Z=>��\7�I������-=�"v�-���%=�6!���������;Q�7��c7�T��[?6j"U���u$��P%/I�Q��t�L�]6���N�k7jE�a��&�#����VK�S���:�2����� w��쏫/�YT��wZ}b%���u��or�s)w�E�;(� {�[�,p�k#���[[�A�>��m.6]&���]'-fAH؅ꩴ�˺r�k�d�P�p�9N�SB�(u��qU9⾍�ɗR�G��w9���y��o|�~:,�l�G�p����k�U�=�Z
upK&"�����s�����VF�I���F��H@���<��9>X���m����e���h��2ع^ȍ;�o�Af�֫'x֌>�J8|.��5�f��xOT�p�o%kvs c�R�r/��5'���uDk9����h��{�������08}'�8J��k����T�妁�֌�N6ka:�:']!]}��N�7��+�����\C��,�x��[�g)ྒྷ�Wb��gԱ@n7�/���+�+��z;"R��6��?\5-ȹaq�����KK� ���ɀ���te=���@�����1S�Y7�U��<�����0B%f
�t���SWox��s?���\�h�`�ʲW!�U��\ ]�I�'�5Oj��Q^=>�'z%���U�WdAܦ;v�i<�@Q<_M|JAf!#��q��]Ej�@i�t�-�r��Ü�\h_t�J]wNH�F��Jé��	�n��� wb���햻-1Z�i�Jv3|��ϒ�͛�e�4��56u������}>	��/<;%�Rz�W1���O�]�.g�[��|N`�Y��p6C5��%D�E�Uu�ƙ_��K{1t�Ƴ�V��F����>�s�^ұ[71��l���!��N���ur�8Z���CK+���ǌSMJ��ȍ��<J�Ζ�ÕQ��3xz���x�L�ko�Wjlh�wS��\K���bc�')�!����8,5�N����+s�n!��u9�P �����jn���x�$����}�rɉ�]Q"�����hvA��'4ν1z�N2*ljH�S���k�rt`vP��:D���n�vN��m���(C������J���*��N O?v�eߪ��M*�7T�� O9<b�Cr�؞�{\S�@�OeZ�n����o���؜��;j7����K<n'G�KuT8*�G�ש�O�i���6�.���`�;I��}J�[�7���L�S+)�"�E�:xm��Me7œ4bw}�'��r�κA��Eϭ1Z���qʇ9ȍR¿��1o��u��i\H�
QԏN�	N�8��3�f�����*�p�'g��(W�F)�t7�U1 TC�O�]��;�y�T�ЖɡN5e��ea}�%#q& ��U�.���}䭯�X�j50f��_L�G%�k�z��Ux��u�@ɱo�/(.��Mp�U��
N��ɻd��^�A--ujO�M�۬�64�Ӄ�
�Ռ�qQ{=�w�� m?��ǁ�V�d ��jk�3¯s{��3r��0�o�[(ak�y�:�`[;t��`or\��y�47��|
�\���K�UnC�`u����P�
�Aը��S���K<�	Tkx�b>.n
�O"�=�DMվw��+���}_ea��[�Z��0o;���s`V>@-tU����u�{NO`>K�;;�=o�����4�,1 �ߒ}p�9l�!��c�"�����l�+>�@�s��˔\�Mn$�8�/������Kd��J��W
��ct�p}c")�C�;���Šn���-�i���)������uP��!b�B�a\C�MC��x'��M������N�Ǥ5������(�u�C�õ�H���6	ZE�2��o���Rv���c2v��q�%3��88� ���
�L����M�bWNQ�0��KX�n:+8q��p�QÔ6R��"/x��U��#{⅀:��dT'$@�0��A����#�N�z�)������%��ԑvv�u�����͛�R��A����$�v.��BW��3b�y]�rv� HN;)��B�`��'�]wm@o@tu�fa�^�&���5�`�'�מ�=t�n3[s)KI�-�4'�j=����O�,q5ݻ7z�%e,�C�۷��T��c8+�:��A��'ol��pY�s�Yx{���,N���١v��o�����I6�`��x��c�T4N۟.n���a��w��7r��@Z>Gl�6�p�eEa�w��5s�P��1�f���N���hMӂi!n�EN�5��>�ݭ����kE�V��a�V7W���K��*~�DsqrU�c`���eɽ��n��ޫf���^�!���x9r�ߍ�Y]��ȡ���Z��݀�g�q�O[?<+�%�wy���_6#�O�]'�5�փ�Z%�~\Oܪ�w*�I���U�5P�tӊʠ�Ϥ�1��$��ϵ�0��ׇc����e=��$��JĵQ�M�t��Xµ���ߩ�5��t�!za3Q)Շg�MPe"юw�SJ�I��j����H)@N= GT�b�[�q���2C؆���t�pc!�p��&6���g6�k(Wm�';9�S,!]���z�!',�+s��"�΍�W���w İj�Gtn�9Sڝ�[�\H��ݼ�23_T�O?�$;�z�3�}f�&�zv:;HR�[co����!�X��H�����q>���r���L�嚅���H�t��=��F͗璜�r��l����Uc_u�>qO���OOe5Hښ;����m�7�F�*H����@���@��A����"f���X�QB������g�kN|g6,�T�/9b���I؛����#��O���EÚ��������#u��ej��֎V���J�Ѹ1j̭;�f�C�n��&k�*���_[�"�ʞ�q2��0Pp�����5�Uvv�3��d��R;�>,<�����,��\���7tIb �[mr����1���M�#�Tu�n�E[����}��Y�F^�������Ɇ>zzR�α1��l�L2��m�ĉ�ՇI�1���u���:�7���qp��p�	C�r���4��m���W�9{ݹ�
݋��ã ��y?`��{���8��++�k~�cVW �QNk���u&ֵ�z48Ϊ=�s�Έ��� B�`:�#�D�NE��̿n�����<���F#~�p�㧡=)�'�Nx���c��WM|�Ȩ���'Q([79(a�Q����SYz�����]+7����@m�v�6��m}���_�ͭ��v���u��rr��Ge�C�U����!�%����.�ɝs:�ξ�\�q)����׼��&�f�xr���=���u�4z�A[��\�9)�xp�����O#вz���-�5MQ�6��ֱ��G������vn��pm�q�=�Ւ���z����1��b����s��X햇��س6p�w��[U%%le�z��x�)��vh����9Dp�)�J�*��P�εL�e�unr���{�=�RP�8]��<ڝ�w*���IC�6y+ǝر��q�Y��E-ֳ�+��N��>�W8�m��#��[T��*Z����ʋ�d��J-�1�;���"�Y��]Y�����C����Ň1��ٻC[O+;{C�y}`PJ��]^B�s�Q��\�Ԉ����|���-�?���j;��1�w2��=Pխ� ���n�ѳOAF�F�Nb�r�
촇d��4��v��6���8j��[�o�4�9nG{�Ln�����B��pT����$�Yp!,i{����I�XW@�.�)���:�77�$�����{����N&�g	W�d�+��Z)�v)l�,��GN�tUN�����k�N�H�CU�/H[�d�0�_���IhG�Z�X5iK��L:��|��31Iq�����i�܇���(�53�l,os$Z�\;1.3[X��;^�X�rou,JZ����t<;���BP��A���$�� T��!��_n�erX�â=s��W���ѡE.�.uҲ����y�c�����p����b��ty�5��g_r&��W�7ԡ���}���{,�ۆ����k듯(R��߫���u\8��ubG�|��vq�Ԫ�]T�f9���|�_)c��FV$Y��f"���X��`�U�:�����nd6�H�ǰ�LGk��rTw�=M�[w�F�7� *i
�b�z5�ۥ�t��@}���ɺ5r���Yֺ��$ti���l�1u o^�g\9�Cծ�։�HH���#�X�[N�e��K�.���'iu 7���ʽ�6�LX3�>Wu.�8�
��r����6��4�IM��n�5�6R��N���.��kw�s����Np�*�rƘ�ϗ+�F�yOn�^d���ͫ�Y1o��5Y)���nPn��/5a
��ݱ�V%9��y��GK:UT�c�b6�9�0���07�k_gv�`�L'�t�X��ֱη��w^�H#J˂���O/.���e�.!.8�s]u��Z�x�^U]�lf�]�3�-*uls��lL�������_n7.�m;v��]�_2���TCU���k�i�_t�yWY}����l
x�ܦ���t��w�Lg[ I�ՙ|��ѷ�X��FT7uwΕwY1a���u*5��(p�f'o��m��ir�mX����h@�\Am`���Z���9��}�����k+ZY���CV��YG0�{�J�>i�i5Uu�D�2짏yj��1�)hpU����p4;��ƞ��f+�'T���u��::���Q��z�;���Q:��}/�xT�fXLI�,���QT�
ċ�,X�������"bUR�V,U+Q�#U%ekE�V*
Qm�R(�ER
mB�Ш�U �Ȣ��%b�L�UE�E�kRc�EbE+PX�+b�ʑb�QKl�-�E�R�@PR,E�%��+aY`�E"��m%(�0q��H�QT����
�#ңAEU��V�
AdU�e�AJ�,���,Q`��Q+�$ �)RH�"E���Y�QA,�����F� ��E�"ȣ1�(��""�PQaU`�Z�Dd,���1�X��d��G���y�~|����}���;�W%����k�2K6i<�f��=H�Çots�k1YT:��x8��c��d< ����O��h�X������7��Qg>|zr�5;œxa#Qj�ϊ��f.�S���m�r��kF��#1}�3��Ld�9�MVx� "�zL�;��DK�e
�P�6+��=4�2r�ĄArW���.�c�5�+���(�%4N�"��?<@L�o�g7�%����iq}���@���)t�Q��������F�U�-���{G8��n)5�qu���X`����b�!�n�i3p����3�2ɍá�V;�%�Xg9����/p.swx3S9�4Ip�x@�ʾ��&)L1�˞�7�p���K��*Ϛ^�Uf���u�^.�JF�v�[�p	�2����(���UEKe$\��X����(m���d+�8��uIД�Oig��S�bà� �y	�j&V���*���O,F��1m���\�y3i�)��C���hc2!����yv$e�y4�p�7�^c�	�(Ƽ���K�*�+{K�zc�M��g�̶2�,��1uP��(���_L���!Bh��z�xH��Tw�2��M�Pܸ������s�g�mmo^�#���qmd��f@��v�m�A��/D,����rr�ۑ����tg���XGI3;~�}f��YyG8�m�*�'Nt;\#ġM�i�G���0M������v�{QA�a�|��^�����)�&�"{)���Q;p(��q�GU���nɴgbN��+�hÒ��eW΢��yʇ9�R¸�P�W����r��Ƌ��(Χ]p�31�qD��Q� ]�8B���15�ɘb�vPV}��m�*b �q{������jVه
��ryHr�TQ��໌�j
�IWx֣��%|}o$��f��8�[9j~===�P�v+PQ�GC��B���Uw�op���B	I��bu�v1tOlh&���y�����a���;�}%�?^�X^�F5S�8)X��
� ��)+��7I%��$�v�l��g3�=�"���pP�x�%�p��X�v��(EAt���(��9Lt�9-�*ivl9@���ӺzX�Qr�F-l��
xh�\�6ab��祐��t�Cj_*5=��s:�[���@\q�OʏI��=�S]��a_��_�NcQᶻ�\ؼ�4�ѽ���������U��E�T����!����bV�t�a?@`{s-fʭ�7\�Г�cK�:d��3S,��\0D�\Iv:���n::^l�*�9`�72�����)~)�����ҏ08�*����vk��ˎ)�)ջ[8w}�GJ"%�ܬ��R�j�o7�d��l��%u���<��6o��UW�3������	JΏFӫ�a@��V�Q�xV�_�v$as�R}�6�	ڲz ��Я/_K;���p�p&8CL��U����� ;~��Y�rD	�׭��g�nWե�h�Ş.�H/��V���Z�N�L:��[�9�����mu�� ~ä���Ҽ���ǒr�e+�/��EzS�^R���=_w����P��S�ύ�����Bԇ�'"r[�X����.#��j$�Xzc0����B+1S����G>��k�G�s��b�V�Ӥ��s�4Hso}]̆jW��XzkE�U���XV_׼��O�M�߱���JE7�JՏ�b����f"=^�|(J�?��>!���bu��b=gܗ�\6+���!�/Z����59���$	��,}��%C1l����E?tz0_��Ԉ��\,�S:<^u��|xn���y�.���04�$s<��[�<>c�Cۇ��CE|�(�썐��zT�-�NY�~㓶kY����T��UrP�*1L&o���ȀX�7��xc��'L\��ѱ�@*	���f������Q�BY��Ѵ��tu��7��jV���;G*��W@�Z�uҝr��X��� lܷ�]��~o`�gR���.��/�S�(<����:���<��s�"����1<g���0y��pZ�ګ�����6��+.�������u�'��Gt�,��Β�	��#>���?��B=o�>������o"Pa����1W���]C����h�#*J�QH�>FɮL�W�]��]<�1��j붛6r-벘�ܾq�'��`�N�C����>�8�$;�Sz���r�����1�����v���$)S�[r�X|��@�ظW �F!#?Ej`e�W/�|r��\k
��m�K��r���l��3_0�U�c�p�+A�nh�OFC��j2�ᢻ�h��w���ti����u��q�n�r��0��rf��|���f���H��'�bȢ�#��׶����{ҕ �4��T���Hm��j/�X�	�R�]BT��[s�������{ϓʻ�4��i�v̤k4�v�uc�Eሱ�����Nh�8D�J�A�❗��bW���*}�[���A�vG��X��7t5�7~XN��w�����y*���рr�����9�[����X:�#�JK�䥎�̫��������=��v��uĄ�i)D�*���5�>�:�5B�yCU��~43X7�TЫ˾.X�r]X�7,w_Gۓy]`)�y��$�Y��h.m�/�Y�����ǝ�6c�!XٛC4L^t�5з#9t�}�D}�z��w�Fץdh�ґ��ޫ@�'�����20��C�#oo;Pl��l��[��3/��d>�ͻ9����VWT�و�n!s�6���xb��n���_\U��e���	�ޥ�/�=���R�`��8����yT���
c�-t]\��B���� 鍁Nt/��Ww�u��nkW'�K��x˛��xpD����G��官�T-{���It{����2ɸ�	;���~�>
j���C����Z�i�������*�w	��15���.���6���iu�p<,v����J�p0r���4ɪ�:�\ +��=�U(��k��O�p��_!*��<��B�K����P��1p{*QY �����V	�uZ���'c>qt�6y�j���\���\cb�^R�	�D��l�=�����:!�R�`��P!ߏi'�5L7v�l\�6�?x�%V+D�����Nu%�5��.�t�wJ^o+z@�j�p��`֩V��=%S�0z�l@��T$��T��S�)��̝4ƌZ�lC�l���{>>�������#6���CFy�G
��P�j
�]" *��t��;]�*}��rt��i��g�J${���zCb;;׌o��W�C� /GS������B����53���Dk��=�:�yϛ
\Ë���}_U��K�L}��y��
y]yQ��3iT�R�G�k����2�Kᒼ�L�ݦ���.��g".8F���WE"�����9�>���a�Q�l�y��S�<-`R���:B���r �C;m8]lh�N�1p�B�T�n�1���'��1_A(5cnx$>�_e�j��l�Q��mv���� �ʄ���n��u�9X�D�U��8o�ޘC"��]����V�՝t�}Hׄs������>Ժ��RYN��"�l�1���k�hފ�A���ީѶQ|x��P�%�ɡW,V9��9�X��BQث�h?��s�d?"]�&���o'.Ϡm����g:��#½���U��U�^�]�����~�-{0R-:��a�.����*��l��ˋ���F����n�D�&k��P���Y�g�CM��*�llV���q\����n�}�ǟez��G�/9>�eW�`و-M�'�:�ˆ]%��*�F��꥽R�Q��9���#YVz�#�N��p�:���l��U���{Ж,,�X��F�%��	�:����0s]Ov�����t����<�T����Xn�,Q�GA���Is�yݴ�*ڔjG���>���[��C�sk�[z�h�O�m�v��0sR�:OV)޵X��)�E滝Y��Q�cX���6�t��C/��"#�P��9�l�����0�U�e\(5�뇟�l�ن;N2�LT�x�S�7WS�F��'���JP�(X=GP��F��.��H��O_$�#�ARf��C��i�t��v����8]8#n>
�Q@H���Rv�v����e�qF0n%j�b{���Lo�֋���xoX�p�u�:GH#9T�DI��4*
T��y�$�U6�t�-y�}}j�ҫ3��� �1�A�� -=�2�V����fv	��[b���+�-�}�p�ZbtT7�l���<� �ȿ�Ȋ�xf���d�m�}�}�:�����$'���;��vW��h���ʅ����6��D����+$�zwzp�������T,�~�+Ep8l��߮q���CL�wJ�=�����R�U��]�E��+.�p�T�F��_ԏ������F��Ca
����\Z��CO-&z:E�=j�U�e4�$Ѻ���5����d1Fz�0~�R��'\>��U
˫�`W�����K���-�Qé�J
�Ы�E��p�c�լ=X�K5
�
�"�I���6��%�mt��w��:�ӄ�>��g������T�:�̿�fwGȤVz�#v�KgE}k��u k��V7;N��%Ag0K�P�t�8]�x�PƖ���V��e�SHշcl*��jn���G�F���ji�|2pUEO�>��(_�Pc�l�����bV�Y�#�}�M��lWw<��rz�L𼔧e-�VN4����?\g:d�4|S�]m{��v������KF�:�x�ć� �ZQOm՝�oC�[��P����ʡ���U��'o�F���:b7���w��4A2�F��{O�&�<{�c�!��A������p�%c�LK<��v��9L�w�y1�
���sP�o�<bm��%1��4��� +��$�9=<��TC�i���-Q2�ś�C��0�i�t�N9GQ�.���m��Y:�20���M��D�&�Yˬ��n[�W��R�`u�wJ�媪w���i;���o��0�v��=�o�.8�C�7�ӣ�}g�6hw��U��؋��U��B��518n຅�$R�]�!>��r��Ȩ�雅��F!pN��'�g�s�I�������F�b��.*�T&m�V���H��zT��0`�e��J�,�<m�d~���te��r��]Y���ZGv��+��OD�Y�*�Z�k�����t���*��Jf��d��3)H	]b�:��|�>Oqen��:;N�ub��Ϯ��m��oJ�T���b���<2E��kx��5Vg;�99s�e���1�LgK[{Ն���Qd�a�ޮ�/���;�aW��1nHTc��x�Y�
A���OU��n��O���e9*��s����`��$��e#X<�u�*�X��ɌGA�(;��}+.��iӝG���l���iT����w�WDQ�Oa��5�~��ąq���)�=�ًm�C��w(8�����Xb�S8���n��u�tŉ^�<�8dK��X��x{��jQ��������{ԕ|��
Ζ�No[ T�(�naq7�UM@w�!"�듆2��z�<���"\!݇�'��y+e���U~3����;d���:�	��vE5W�5=ѳVmM�:�e���d�to�;�Փ�#�ȋ�¯��0uJ�u��p��������	�l�P����E�,S�؎��T�Z�ĸ�*��v��-���'�(,��ٮ����rpi��Y���k�G0~FZ7d]we-B���iԗ)���g�k�f:Z�7}u��w2�3&��W�
v�zP�=��e��U��Q�0�mB��j	��Q0������=�u�ih�v��i�;ǯ��]0���.5����nl�.�Fj|�)PY�.����mB�:�rR�-t��l�]��D��Vp)s��;mcו����`�|q�n=���\�n���39e�ˁW>�6u��}L��1,�ļ�v�\:
���6n�]b����u:O�)�[@'����'Q��h��u�#B��1���O�p�߶��J��r�a`�����`�\�/s�]pQ���Oԥ�qL���1�਷j�|^�e\�;�W�HF���9��L}s/�Bf�%3����&o�s1�8u@���9��Z����e�E�tGAD��A���Ƽ ;h���wzp�M���.��C�ɞ�ps7�#�� R�N�"
ҩ����-�l�{G������Ɋ�z�+�V��s),������)>W��C�Qc��� ��:L�,�����i��
1���<mml��S�_�P�4���|�SI�*T�9v�U��O`����]�r��������Lu�/�c�ME�Bf�̶1:��9(}���y�[G���vw\���U��9��cpܘB��`w����C�gQ�0���	N�Ħ���U?>�"�(���`����M��(!�J����Qx;2�y�򿳗�g�xS���
��^�n?U$-�PH�쾁3�k�����-��}tI�V��ӓ��c��,���-Vo~[���coZvjs��v�G���]��`�x�Rn�w��>ނ�2��{{��K�c/sn�x,���}���nѦ�V�}����ƧK�e����٢geԂ��Ge�	
�|���vM��5@�C�.u�݌�{٠aϹ�b1ǜ�q:c��j�]ߔX^ߍFR%��#g��v�T�,����w0.*I��hW#j�Q��d�oF�3q;
�fl�^���mJ::r�h<n�J��e+��i��Q��;t��i����58�LYv��:�+�+K�+�v�VRW�>�P� ŵe��ep�U���RS����\�1����zb���.��t���s`�P��N���(Q�|oTʻ���2����15�I��@�f*�=ҁM
[جE�v���b�=���z�Ĳ��xR���Y�g	�+Ǘ��-��ԣvne�NL��>�/u���RZϹ^T��=��[��X^�ٝaB0�<[i ����]q��xE�թ��;9�j��L�(tt��+ �urx`�xb�I|~G�#�p��-Hve����O��H�%n۲��('
��\x2�r}4�7WƂ���t��b�w�+��@�]H��
*����oC�\I���)�ϒwu$cԂ�O�*�X�t��M�e Vn�4���S
�a��v�c��.n�+q���lI�#�*�/r�Ng7�����_e.Ր�;W�sCkYGgʷ�+"�F��ˏU�MpWi��ֱpj����L�i�	�LEF�V�����H#ʂ)]����Ӑ�Bl
�k�L˝P�B e�M�ӋV��"�k&SA�����+�n�,�*�z轓,)�J1� �>k`ۖv䮣@&kj74!�MZ�W�
�Y���}����6�`��]PMz���U���tS��[�����_'�S�Wz��7o7,ܢT�j<sZ����N�>�tN�#آ�)�2��h��ڢd�!�/(f�u�WABXق�*BK�%=G��\�\�����\�!�MZ��.�Z��z\��m]�t�_����]��g-J� ��q����w�De���&�Zo;u�0�>k�rf��z�ϗh�#D���)
�t�2��b�v���4 ��=쿺5�wR�n��j��:�����'sCk#��f��-��'KE��f�+$���Ô�:�.�R�z�w`ܱS!��O[�Vks��g:r��ضD�ebt��w� εr�ܾ�5JG�F��լ����qV��=�y�z� ��t�<�\)GkC�>�v͔͙#����Di�W��c�ڶ
�鬃�XUu���1��/l��w��^�{��o�S�*�1Uc*��mUH,1�Y��"��ZPPF*Ae@TE��m�E�H�m%Im�--H�*�Y �Uq!Q��"�a\�J��*Ȩ�"**�j"�*��Ȫ(�1(�m�E���ڠ��b�ب�Qb+1��H�b+�*J�"E��(����R�E�P��E�*P�eE�
-����-�[kPDr�1*���X�R-@YR����B����P��(
!PQaZ *����#[���EE�l��VTU+"�iRT
��XV*��*�P����)[h���b�1b��F�a�T-�[F�E�I�KIX)+QH��ģ"�H-}W�s�'p��[��/�j��F�Yܠm�F�pS��h�e��;��\O:$�eͩʅ,��WvL�����5�3�330��-�s=����ӟ�%[��q=�b���HBB�氡d�1XPn�Sؚw�M�*�2�c�}�5�T�Q���Pۆ��vC[e��)"�i0��QC���u0��OL���5�q��cB��-v��s1C�c�U��.!�ö	��PJq��J��/{���8���,�"�1]�g>���.r�})��(1Ъ��g�9DF�ܜK�Ln�t�4%�lt��,R0�e�E$;	>�x��@�v��(E�����P^N�Z-�*�* ��7��wB�*P�Q�H>�\�����q���i7�y^̱Sw��^6�s1�����tP9��MOQ�y�ß0���aq�u\��y���m6�=7��ʐu��zy_��4�Z��q�taةV����V�~@�÷��н��D%���u
��i�Q<��N
�n�y�(1@Od�Mㇱ��/2�
�ԃC��[GD!��j��&kE��l�n���(X��dRrD����ď�Tw ~�vv=�S4J�/,v����^�Y���ʙ�W�/'�8R<����J�w��g�ή�\�&��Z�b
0��bY���Ƴ�\��+�ɫ�i��&dB�8�.�}�����Z��R%�R}s(��1�
[z��k����
��2�yX���C���Bl��؉���y
��ӴI{V|��3�t�6�	��X'��E�V���]���ncEB�@F��h� 4\	yu����aw��vSG�ä��+ha�r����W)?�up�zI�V�P����5��Y����[�j���۸y�+2���{M:6�xU��U�J�^?��z�z����f5k��d�X�ٷ�5�q8j�=vܛ#9�Y�k܌[]{Dy��V��*fA���#�,���Obwf@�v���5$\7����-��~�.CU��+�����}���*e��=L]�f�任ap�k�f�jP^GS���(��b���=���;xOʞ����^��v��9���s�uz�agU}�cwYT9�*�e�N��Z�������ˆ/g�5�s�'$c�B����ظ`�7���A�T߀W��aB��0���N�VD;|��W&�Gw�Vs�2p���s�5^�^;- ��� +��Mf���)�9��_9[՘b�vT,�5[M^�S�Vf���Ӹh.��Ut�3퐜e!I��lo̺&�i0o�X��s��+~������c��yo�n��rF���r������<�x���C;E����'��e�-V�[����_7�[[t�M놌JK�Ab}X���Lm��^��I��R���J�w�=�

Z��̵3���0`0r���QK�wK�͍y��m{q�r���.���N��쑲K��Uu���ւ8�b��[\�]ګ�x�/��S���e�	�]��D��4TJdT7L�,��0fb�M�]����%�)�3e�߉H��#_1M�qW�͹[|
�\ ��)��b}�Y�6��NZ�/�l�8����e��K�9�ؕf[Wi�#���\�*�_#f�s��>wW '��5�QU�;|)�"8V����W㗥p�{lRsxg�n��Y�^lP��}1�E��7a�M�t���1D�iD�h#�n�e[����t/�&��C==y;1wWs���[Y}���>�%���ndCW?6�V�=��J����	������z�A餺�����}�0����+��g��(H�k}Z�黙\ukG,+u��9|����㻳��Y�����`6��z�c��u|X�ă�@X#~�U���d�A�%�����f����Z�V�W��tQd|h-�w����E#�}���MĹN����U������
5���B��w�λ��i5S5޿X/<���{U]=%�Ra rtY��\��.nKX�n]��{0N^z	��[�*�(�q3�ն���Le�m>�&v��(JW��J�2�/)��ڇ����ffeo2; �s�d�Ez:pC
��Y�FI������Q�}�u���k�����r�*�}���#.qQ�-A�n�ү�ܜ?1[�~\�9>o�UQW���y�-=탻a��M	͍�JG��5MطM}1���g��1��ǧ*�K4��_Vd���D��D^��u
��n��>��|up�7i�܀CY���&�@
�������������ʸ�̠*"�g�DmDpV�����z%���`h�N���R�K���:*����V��đ�7/�xh����x�\^�.�(�X�}p��X=n�`��)Îz��f��Ei-Q�u����Az*;H	���nJ�C���ь+�]`���P!�q�W�ռ�^�`�nF�q��!�%ˑ��R���o�xX�-����z���C���n���)�yN	�h+s�9�u2�Gl7v@�,�&Zz(����O��(ԢE�~�u���n6�T�p�C4���b�`�Iճ����Py��>_o������u`�]A��מ���n�Y�A^����Iwc]v�U��iaSW���⸨n�s��dn�υ��k��X��e����������&�F�p�&����m�sP+��Jk_^u�޲��a��t�W^�2��$�p���}}�{���������0`:�7k�F-�R[ͪ2�m!
�S*�H\�T[j�k~/.Ĉ� g9<~V��97[J�ƶ7F'l6o�ݨw�K��Lp��ل�7�hdr�,�����T5��4��.�lTL�^Z��A�Se�2��rc���a�N����(yL櫨�T�q֢��'e�����k��Ə\k���Pp���������qx;7��yw��Ù�o�������u�n�`��^���r���ư��b��.�X:��W^�9�u��^�/�0�چ����y����]���]F�L@�R�£al7�ó�5>���F��uIWx��rV��I�ٍ�i~��*�u�
����;���ZTkun|��5_Xn��� �cfN�A��;��kQ�.����6��ETb���D�����o��1̱��U�hf�/2N����`]ȩo��졂�����)��W�9kx��Bi}�� 'M��!��BҺ}-��ؒ���^SR��q���х�K* ���z[B�.T\=Ƨ݈�rс#�(3!���l�ЦNeiX%}[������ ��ǯUz��v~^f����u�\�n�p��������W���葥�A̽!�P�,^W۪KrM�۰�q��%S��C{��U>X�_,�p�e_e�/E�r\�hw��8�W���lIP�%� \�ߘ3  
Uc�
�֦sy���3�F�#EYB�觰AH���Ll�bw�ٰTz��TB�)K.��e�!c�=ʇ8�c:��x�_k�9���1!<@+O\������3���a�F,���tY�we�	�8�e���۔��X�g��tĉ*�$����wW45l�U�ݩ們|���5[F�L!��aZ�և�j��� C�� �o�:Ni�ۻ����}�;"��p���r��u�j7�qvq����K�͛�� �%�z�DIE�W�#��������� Ui�v�¼c�����lx,��
O�Pw�����3���lⳁ掰��2�|��>�n����п��4,��Q��΢��:���X:�61���9�
���*��:�Y3����_�I����sݐ���-�)�m[����Ĳc3-e�ʶS�P�. ���#W �S��3���๾�������!�g�;y��4�x��������V�!�-oкݟ�1:d�1l��;����W���\f��b��O����f�F�e!<�x
ӢLƮ���;��8VJs6�SkoB��cuE��:è��'+ki�7�|@���z�L�6���3��<��U�qUu7��7�wgX�\��w���Rќ�jS����'n��.6�<?}�� ͠�ӻj�4Q:�n='���SX�e�VUG:�Y��N�����|b��ֻ[=�eGV[O�Р��y H�%�n*�z��Wئ7��V<�Ǯ �^u��Z��{L48�c�/M^r��6� ��X��?��Y�F�x!���u�]�X�WI.���p7k�ѿ3��9��WK}��p��q<�<�͔��i1g���t��m]oF+��m.�#�N
�W�A�8� d����3�����$t�3+�T�(��ػ���+�$փ����s~�c��T��ܚ��1�EC�R+�雅YD��psuMR�HOL�o�4(���"	H�?0�uE8uP����h=��@��{1�yWi����o�p��Vr�'�<�,u��5l�q�6�Xm1?K{P����Do^��w��wkSWN�#�]� ���%���RU�v(�S���*!�.[�j�ζ�xD�}�d��ؤ���c_ה��_�Oύʺ�#m��<Nو�4�v�uc�^���yS�r��\�2C|�KnGvb�Cf�Fwe�++V��dÕ�Q��H<��a����c���89D�+Tq����.5�\�|�U��c��	���ŭQ�8&��F�L���; ��Q2;1����A�}�W�}�_OEӞ�QVt���L�,\9
��U"9��� ��<ٔ�iȱ��5�9ӝ��s]�]=����
ct�n��j�ʄ �JXb���r��ĉ�
����s`+��q�0V�f�|���g]'y[�Y����}y1����ӛ��2��mۨCM��ª���G��0��P�L����O��bѿ�%�ڎ��7�ꏃ����<|B���ј�����`�b1�ݞ���X2�#fĥ���Y촳ʧ�����?�=ՠ��$Ϯ{}Юv=T���@���N�f�lfb��Q�������N[j�^u��	���w)�G�Ʋ�M5��#]s��>���^�+�4f^-�U��Nہ�Z��	�4�"�'e>wZˇ�v��*�7�+mB��b�{ꉱkw[wQ�ʉ\�sV�t�X�l���8}����cMӬ:�E�S�]+��5�gO�5��\�K�}k�_�GJ��E�rc�����5���+Q��gn�u��O��1�xqۧ���4Sp�e�4��H�9�5��[�{W��J9���#���JQ+ʡ��ו�l��zS�G�^�^3$8s>c����2�*��.s3!�W5y�yAu���Ø�EN�En���f`O
ȱ{��D^Eb�*�%����	���wڛ�B{�����1�gov�F�?����	S�0Aף��S�[,g?*�%�Dt���;{j�=�uӏ��}9�w�f༎�n�Jc��[��l�:d(��o�k��J�qy˻>�#��:�����LC�r&
�0���H��^����7"�;'��u��3�c�I<NB5%Sj#R�X�Ԇ���y<*j1rr��Úѳ�����=��^mI�����5h\6�X�|qd�4�^�N��@�^�9K���^�Ջu��w��1{��(��SP�ӄ�I�U�yr��U�C�kg���nQ}���9�nr��k�Z�7;YR��6���}��'oEõ���\2�
��V\��`�v��������b�eV=��o��blW���W��r�6�7&��l\�vst���o��;֭P�$)Mz}����aY��lR�>������:6q+84%�7���<�HV���4��1�{�`�Y.�Z��%�t�9�s�fayxX���j����]V)[٫w+�j͝ u}Y#�����'��0�j�+�i_p͑m�#C/�f�T�1a̮�ś�<��7�U�[ōC[���=�P���H�Ȯ�C&Jk� �9��[��K��>q�_|�����E��͌[*�۷M��t����Y��)1W�Wb���k��Eų��!����S�2�lc�m��BT!t(��s0�i�壝�T�J��}����Z�ꗹ���ܯdӤ� ;r� BZ!,����`Mc}VKl�n��u9|�n��n���ܾ^�ҏ����˩���կ$�u(��m�C:��]�ۀ�e�qn�K��S��q������y�O�����-��Ź��2�&���o�++����V�(|�Y|�3iE���q�ռ�ٻ��(7/<��Ṷ~y���k����-����TҞ�����s(zI}��մ:�8
��c���_]yk~�fb3�u��_Q�]J�e�^0���+�<;&Uɼ�Z��u�a|�Ż���՝���8�r�tV֤��<�˛f�r�4��`���j@U��i>{/�C�m�%%����*\{��`�]K]�C'NǽSS�ml����{�-\Zw�ަ���>۔��Ӯ(n�
L<j�`dTp��
�S4ٔ�Z[��̻��fd��r�F)fo�]՝ ���!'�E5�15{c 47��C{��s%��@���4i�N�Z;��O�ܩ Fv��%��ǋ�b�>�*�1�J 5��DͶ��V�0uGԎI�֫v��	h���m��Aj���m�*�/P*mw�����B�N�ӬP�����K����yB�v�V7�%E7�;�7����u�B�A������w7ʣ�j;�wu�ua�oc:ȫ�w�hZ��ݦ��β��_;��k��ŢH�6�΍;�����*9B��K�vsP�yLQG��'�x�c��M��:=����X� ��ICN`�J����&�%Yʯ�7�C^k'59�����ta\�*iʎ����TI�f&�R[�n��T17n�w�h�M�n����[���J�nwQ���p@n�у�
l�v+����	��qwBL�=�e��]����@�z������R�bX_���8�$����o�+c�V�B_Myb²MZ�.o-�ۡ�����e[1���|��T�֝�F�_<.A K�VU���fݱ[�&�4:��i�W��RR���^ ��n���r*�=�;V�����g��|D;֢��ZBFX; 4:lw�0�v���I�v�=�GU�uN��nĘՠ�x��;A���m4��F�(̥��U��*W���v��7o7�]h��u�GHm��]-w�ﺱ�
O���>�ȝ�YX���;�<�к>��{�Rcw�ӛX�Hq7}79�쥹�uv.gR�i0٣3T�ZZ�7n�]�.���J��@ �B��p&�,��;��^�$5��#��L���)pwQ�F���մ��0[�&�Y]1��k5p�%d��?2�B�v�i=��G�!T�X�#�]F�|t��˕�V�����Z���]#�0�`e��l"�n�H����2ie�h�$�X4R�p�a�j�Nw�v���#�Q�`0G[��k7n&�9�Ѝp+w��%m�ꅍ5|����W]�k긴5�t@����}���*��Jf-Q�7��=�ֵd���L��m��bt���6�AG.[H�2�J�	�,��]og!OC��E=�v��qˡ��u"٦�M�[������7�x�AƩQ���ѕ����	�{R�|���8���)WQ�+��&���V�VnX4 )���u���{5��<��η��ZsHW�8��l6��9b�pz�ۥS,_�O�NڱJ H���Gl���V�6sD�u�-Ǹ.��6d��@�7-�80�)p���/t��j�#��a���~����+FChbX���Pƥ�I����J�Q)j��P��W�H��.YY(ԕ� -E�-h�-J$�FjR+-�Ud�R�,Aj���1ơU�B�
�%Z�+Q�X��V�ER,���E
�Y�1�%J��B����VJ0X�TQE*�((1���8��`���¡R�+aRT�XQ�V)!U�1$���+X�Q �"�(9@�1
��R�m�*�B��T���(�+U̸�Q�AjEK[K,m�*�T���#AdmB���ł�dQe�,��J��E�X�B��RmE�*���R�m��Ke`%ZY��+& R�T�l��b�X�"%jP���VT"��������y�^��PK�Ьf��Y�{td����};����{�N���&	K�Y���IɎ���S��L�b�Yo��������ˈ�z�]���:GsJgyܺG�����U�(�[����~<�4�ө�Mm���k#V�{S6�������\x�Ʒô����c>E��s���Ѯ�,�����W��}}'�Sm~�+��i����j������ί�mqkaO;܈�ث�����������GW�)����鬒Ţ{Y�b��}g���gUe���4��-Ϯ�w9����o��3w�<y��C�2��*kU��b��
t�mS�/E��,9��O���:�&�]=������_B�Kt������;�OC�mu�����s�C�˟(毡�]��Щ���m|�L���:�a�*[�˪O�Ef���p��-%��f��:�u�V#��y��7uN�S\�ghlNT��P��`��鯔��Ox+�lӤb�ga9��),��+�V��Q�ֹ���إD
#Py���J������!R�UHEQ�U�{��&E;�eL�!Pb���b*T��5�|�I�����R�bA��k'tP7^�ò��հ��Z��o�j��g�Ʒ9��Vh������o�]�y�-J�*I�Yeb[0�<fN2����vw�5�jb�d-wpf_t�p����P��y�3�k��wN
w����x���N~��/y�VT�m�YZ+Wumai�����5=m?*㩻a1�~+z�-�aO��qc��W��>�ٵ$i/	�Է���]�m���S�n���:@�����J���ޘ�}|�z�s���i_v�����뜅P�;���X�am�V*E}��[Ž=}������W8���3X�au7q����\CX3p`d6����κX��9�_Z�W���r|s�r�h\7��C<)*頰��lQ���Q�K�VZ�m+�ʂ�qM>��<}Oʧ��_S߰+�6��9�"���w+O�Nw���-��or{(��k�u>�~�9"�o0Is��]��j{z�o!_[O��K5����Xڕ�֚�6D�B.K5.�Wb`����Gy�9�b���fq���xʎx�t�`"����B;����[�-xr�7FP���c*�O:��=�������]�Jn�B��*�;O�8�q6bSxR�����r=nr�	ݗ��V(8�������?������i�}��]�[^���s�Ư�MnS}_)X�ݽ��Mљ�ڍ�;S���ݨ�y�EZj�-RvS���=��z�r�6�r<����5B&X�}Q��>|�_أ��o\rm��n8����ϳ��#�Fp^J�=[���5���"\��.k�_�neq�7��I'����U-��=;���y<�%�ϫ�B}p��c�;o�g/w-[Y��-�Bv���4pJ�C>EV��s�ekówR�L�u1;<M� �3�R���\�|��}�8��/#���Bc��F���L�����tg�泻\�>ݜי��er������J��
�<��n\*��a)r�z޵�i����OFb�W����P��i�낮�v�kT躛sۉ֋;�%*�[�kup��M����.arW$z*7��IP�Gbs�@+]�Y�T⬙7��Om�:>����lh�V5Br�\l���Ej�)�w��ˌ�Gm���ݺ��£����Sg,���Έqu��斺8�.�
����.eJ��P/yB���z���i��*�ӗAհJ
�eɏW���ꫛ�U���䮕��u�Ye���;��{~+�ߠ*u
���V}��Jgմ�fy�Se:����y�y��^�kg���+��Sh�mV$7�����B�\w(��ب�kE��Z�-��c2������R �.�s-��ơbwHu�.u���p�=���]���Wc���U�s}��1��ʳ��4�<���7s���ꬸ��m�MnD;}P��"����-
��UѦ�8U�u�AsWq�pb'Z���;U˿��CZˎ|�S��B�M�Uׄ+zs3��LK���ƅ������R�Rc/��#�'ί�B��'p�h�i)5������.����ˣ#5D���
�Mf��Z���Wt^�5�;�7��i\8֪܌g��Al��n�w'����k4-�e=|T�ۗ[΂�qs��;�s����W�8�n��;O�ٳ�F�T�;�u3e���3^3�#�w��B��R�a4��P�-N�)Zu0�Ɠ�R�S�����!�wgLB���m@(L��\Gu�&)��c\uG]��}w]q�2��7x��6���/%=W����m��K�k����٬��G���W�R��}�Os���זfpO�K��o��
���'qnp���/s@�K�&�6���m V��F'��^���}N�P��	�Uf��J8y��<��q���\8L�+r�t�<3���'�	�cKɩxT�j����;B�n�4����@?G!�~�s��ޚR�2��y>�	��^�ɱ�f��s$��Ӯxq�U�g_\::-�.�&{�G/[�������oZJ']R�w.W���Su�9ĆCC�=�>)k����=�]��U~�!'ڛ�F�>�u���g8ל�SB�\����Q�+IT �t���;��A�R������_[ڣ�1.s��ظt�9�Aێ.5��í�l\n2Vk�d念`wC�:�<���E�n�ry_�Ubj��la��g7,^�<�M{x�w��,��;� �\4��iY���T�*�8�h�s$S��Ľ}y�]r��@W� b>�s���z�����҈�v��Gl-4,^�믓v��W�S3�ə`��|��+w~z�����A���Ǯ�(�WR�⬙x�dʵ9ɜ�d�����1q�f�t�a�l
Kdiy*�#��&\}0#u ټ��6ӥ+/�����Q�;��z��g�g,�MC]�����Ձu��zh:~G�s��f+�r������?I2!��Ӷ�oy�j5��.��7��V���9�pun���}{�����z�H�gU-p3tU��֎����i��v���\u�b�	-j��v�&��sj\�]ws�Z���z�uD'�8]&��M�gX����{��)4��TJk��ς��	��.�s��3�s���7o�ܳuk_�����oaߨb(�xB��=�q��������24�jo �ާ<�OOv)����|U�7@bc��r�>��؇28Z}y���!�g�P��-����I�M�}e\:F��Cn�����iqMe��u`A��uJ��T���s�A���Xv�q&�o%.x½�0N��ȶcUe;��=�vFJpu���ꈼ[Q��ME�J��r���n�x�B����)e��s�ڬ"I����J)�\�:��ޡp�]�*b�D�[�F���/�Ӝ3��?V����c)^:�k՘��?nr��+�
y��_M�lttoW2�� 2��ӻ�s�P����)���G���ڝ����)��;¹
�wm[��>z�y�N�����ϻh��9I�`^�C��죎�ު�������|/R恶�{6-�B����o��[4�\���.�|q]����P��s�ʳ�V���ROz�E�ԗ���fyRKhq��<B�B���ù������{���B>1Sm���\'���-��f�]��n}*9��\���>כO:X/4��3���kO�S}P������=u��5��EҪ���wZ��.%D�\�t�������~��oir�>�'i��&7+�����ŉ̋.���K�E�Y�9S����w������P	2m���+"ÈX\�BSa*�3.���n��Yٮ;Q����+�+���)={�S.V��Z!,����\.���AĒ���r���7�q��sNu;�g4u��-؉Hp���sϫ������O
xġ.>�t��hf�����K3*�sz#��֋Ԩ��Q����뢒�Ⅾ�f8�]�`��h�/(�֫��e��.�Gn�i��x���d���x�1�Yϛ��r�r�wA{ˢʷM��7��c��Kk�ep��}UQƛ���]�ٝ�g&���;G6Z�V��S&
�ϔ��E������ؔ�&�d�'�|VWܨeD$����}p���G�k4���T�ܵ��Q���{��3��������`s]	�"*6�T7�:�`��y�m��{�k~=�.�ǵ����u�wlj����\�RoP��=V�+�슰�l�t�>
��G�%�ܭ{w��+�%ߠʌ�%����>�䯇dMOd8T�pϡƼ햬_s���q^��w^W<"SkU.���je^��uz�j3��`؆�k]�챎�����<�^����������9�Z���g:��:�q��s����x���Pﶾ{ùpוAe�
��kUB��v�TO9��Ug�ڕ�څ�m�4ֺzEӤu���S�d�K�P��I{Ƣ%D�Q��Tb��
|�kXt�3����V�YG��j�N�����5�3d���҃��G��^��9�6��Ҧ����^��H�ݗ��i���We
H؛2ғ���5+�����QB^�%�+F���y�7�2�;�!#����4���Ԫ�Z�|�{��n�v���������H�pξ�ވ���u-��T�6�,���c�8�����{�Ncr{tW�>�oZO=�FW.UH�ۖs��p�*�m|]'���t��g�/�^K��+�P��m{��]�-	¾٤�V�w+�q��(t�u]w=ܝ�&��caK@}�h�mI�ֵO9	�ܕ���J~�bc���T���]�;r�͠�eOJ|␗��u�qN�m.�s�ش9��d��.�u�Sw�0=	����hC�CD�Z� ����2�&�����V�ˮm]՜Ŵ$*i��ޢ�]*2��n�1�({���{�W7�����r��bH�}�5��֋��\4���t�P�]|V���
<����{س��׫2?c[�"sD��J�[�G��O^��U�-��л�s��)�i������}�9_Fb�5z�b9Sw�W�ht�۩�z��K��eZT�"�Y��C������-�,x
޲��*�Ū�fM��J�k*n+#xGq�>���2{z���tқZ��[*��Ѻ� �/�ׅ�\���f�75_s94\������|X�Vc�Lm���W����
�jvܴ���%�������U}�|�z��V��>:y���iN��=Me4���qֹ�����蹚hQWj�Vo���9��.�Ys���TA��9��b����OI�C.Q9��=ûy���v��R�zt�ʦ�s$7xyTU���90���ck��s��2��]�W��^�{^j�*�χK{�u
���'{b��Q�:{��	s�s�;#�-4�c����&�5Bꌃ�#]D��PD����w:u�@H8�λ�i󡯲�Zm��n6�cw�в�)\��:�����yO"��%L�\�D_5��t�{4�I����0�7q0��"��hFʫH�;��\Š7��#�]�ޒ����R��_��h��"��C��M;�}�^��G)R�5�a)��ak���J_{ޓ%�\� ͮ3�ҵqꜤoc�9���]�J(𢷨�s\Ji�%��=�.M�wʀ��D����蝐���W'�i֪p�zH��5�e���vUʾ<NE�p܇���tc��=ِ;TM�0F��gc��D��,�\Á��N�r�S�K'�.�Egc���}I����Ձb��殴�Y��zaG�M�<nm��Y�⧐y�yܮq��J�`	b�q)��m^p�2�ӛ:[޵IW8�}��߅����M��${ǹC�j�c�ڢή{�k2Dٝy�v,;���N�UXԃ̺�eѲ��U�a�q�Y-�4Zq�Ok+�xMXڋC�{w3��sL@�\֚��*��"̃i��q�vz����-�pCr`fr����*�;`Eup6��֤$ne� CF�i���L�m;V��I!��w[ܵ���+m�"���N�j�������)�]nQ��i�y�sx+=��4�k�Gfջ��꾷*�|f�
�&���8�<�#6 Ղ��y���V�v��z�^�7��IL[H@*oft9t�Tgrj��� �Rl���Ԣ��<�E���HX��k����q/�7�y}��P]�+r��]����}�8�#���з�SR�q��j�DvP͘�5C��9��9ǥQ��׺�h�)v�8qIv�4�%�)]_m��.�&;�h���gT�����Ӎ�Ո�Z��� R��Q�'R�f2κӷT����bV�����Z��O��x�d�+Fr��h��;FV��z�����k$��8�

��E�K8�m�w���]��]�E���z�×2�<Z�c�
�3�2S�=�#u��������e�_LU���VC�0�J�&fά�} a#I��Gs�Q�BiZƄwS*�R��3En=�ZZ1��ί(umgc,�l�aa`!��s��ʺ�,���'���̥����b���v�춯��m޺W�W3�ZU|�/�ňol��|�S���R,���K�z���G�(�GJg�Ҧ�͕�8��T4���٭�؎���/H�G�m^K�Ά���В$=ͧO� �y<�Qᯢt��!gQ�Oj�p�·;�tt��l�A�^�V���a8��X ��+M]��	�u��]Ar�v�]I��n�̩:'um��*s��8�п�7�{{3sޕ��YKeɼX ��f��t�r[hƩ��ל�;�n��[�[��Yߊᣫ�"M�b���fO��h�F(,�}���6��{�kvه]���ȱ��.:���u���N�/o0ґ#x��l@���V�A��=q!��.��.��=em�&x�xkk���X��&��̘�[�Z ��k�ǫi��Z�{�����t=�y��!�#�xV��A��W*i.c���]���˂���\�yE;j�r^Ku3�,�����Ű+FYN��9��Nb�p ���t�`[�\���Z�۲�����R����5��Q!���Rͨ!5�<kWp��t�ͩB�ӑ(�/�=݋�]�n���'r������}� D||�ʀ�`6�֑f4�Lʠ��[�1D�`���������R��P�*4�D�Qa+KKl�
�Kk�E�Yj�*��6�D��̥Vˈ��bdT5mr�T���F6�X
���X(T**"T��%eV#��kZ0s0��1�(a�"��-�m�QbԬ�T�֊
�RTV��ƍ�YR�E�[iYU�Ҭ����+V1�UTEb �°W2ሡD(�m�����-�"(,�eUV�T҈(�Kh����U�j��E����Ŷ�+iZ�cY
�Ш��ec[%"�laP*T��V�IZ�U����j4��m+*TY���U�AT���P�V��[J�EDF�\�J���X�-e�����A�{���×�����@4j+\9���[-�ͦ&�.�q�y`.;��T�]3T�%0:�d]���/7��\�E��ܦn�舏��hv���?Fo��5o�k�st&8LA[��հ�ciVp87s���ܗ^��\\}�;o�ʎT2�b����z��mdAZ�Ft���
���q���v6�K�)8]��֙�Ţj;�NC߹�Um�=;�Ap���F)�-&��B���(檈��W�kN�z��M^���>��.ԧ�:����ն�,�?+S����B�ϴ�Z�zJz��O��|[��N�o\q�}�1_��J�$�Khq��\w�LuAu/Q4���W�≽���n�IF�T�^~��;܋k���{cwEXڞvq	�y6lEUc3��]=x�g#���Z�b�-^�)�y�EsI�6�}���V�L��ą�6Tfo8���r���U+�n���Xⓕ5����h\b���B�
1�1i��A�5������T����;�kW=��'{ټLx�mS�<v�\b�n��aQ�`J�#>�¬yR�eZt;�ŉϷ�,`��v��x�A��B������,��tz��x]��_s3<M��`���C2����S�G�K��u�u�8�h|їλ�oT������7LwK��4��`o�ӷ�����wmd�{3ޑ�����^�T��:��ZJ{��r���ҁ{S{�]`̍����v�kv�S�6��6�s?�W�k�-neA���r\�9���/'y&;R�q��N\��	h������񆧓];Qr���Nt�w;|�1���z�Bs�cM(��
+z�sr��dEZݔ9��Z�Ѕ���u�ⲡ&���=N��͗��݈���ܬn��뗱�M�C�	�ql}�_b{����tj�觐.�ی���;=��"�os��=������I�|��*��J�0�K�]��o.�l��b�\7̪=�E.!y:},ej�b~})������$ȫZ���κ=���K���u��,��߭�^NNA�E��u]6���V4k.�f��SP�-�ه��M`ʎcr�쯎+�:�1�b�0%DxĪwu����c9�u+�ja�2���&Mu%����V��h`�.�:n�z���(<廗��
�mn@j|sa/z����ǹ@`v���V�P�vc��q`��γ�'�s�p�U��P�ܭ��kx�o��\m=�jΗM.�%��Px�CH�^؄�]Z�y9�bG���p����{;������4c�ߪz��^�x����)���N�H.����@M�V�{�{9'�y��+���q��\�6��r����k�X����^V�SÅuC�a��X�����p{��F����oh8�tU�S8�Yh���;b�k��HiP�:@:��C;��ox��OvA�h{Ұ�������k�x��]�N�M:�`�� ��(P������Px��i�.o�o �4Ҹ	6���Dc[E�upx%�Y#z�\�Nn��D}�bS��[O����>�%p�w,q{N����+�j�2:�H�"��� j��~��L�\����i|�)�c�jw�_�o���F��kTpi��R�|��⻜j~�%k�»w>	�7���Sb�����q��#[�v:9����oPp�^���LJܛO3���I���/��a�P;Ҭ�#Qwu0C[�58�ӻ��D�:�U��co q̭;�k5J�X�*�N%u>�`�f�ܧ��m�n�f��%I�R2����{��Ay���R�ks�̃�H�=N���v�˷Q�b��_�{3%Ϋ�}�Y吭Մ��������O�r�\�!ʰ�q���횋���t�{�F6��!����
��C���F�U�(�w���fŇ.tV%�6��D�si�6���=Gj�w�V.�����/g{�N��8֣\�4���w������^���+o!9��#�O���i����͊k ���D)�!��ʃ��-��ʌ��9��,���ޮf���+���X���Ѡ����9_;���ī��ř᎗R��i��]�f�&�v#�sB��s��.�{�j�vW�U����1ԫ�8��Tζv_v�b;�O_-Ɵ.��N{y?��iP�:[G_��#A}gzw�&���W
n��r���e�֛[N:b�꿗�p�k�ד,�����k}]�������Uj��i�j��v��n��i�p��Aɮ:��c�T��G�{��um
�t,�)��p<&ҕ��]�!d�m2'5�Y�-r�Ht��Z����gerN��#nJY���w���N"s��b�[kw�������꼔͕�r���`T��u��۰�{m����]`VZ�7-�35�sx��(�<�c��_
��h�KU�Íy_[c^�N�Y(�
����kw����~��{�J��b>�������E��eq���S�݅��U-J�prQ����������	LWL-u�f_�Q�
e����[R���;SW;���GJ����Ю��9�&V�J�r����K����p�ƙ��[7\uCv�8IY������a>)�G'�y`�~첾���lr��䘦�C�^�_!�:�#˫�mZO­kW��x{�Q�����:�L�f=]����u�B��Pv��:kt�{J��uE��f�+[�ڵ��]�{k���oyGB�뜄�L��q]X1��G����9�$Gw�N[�T:-�.;Gϊ)ހ���ç��f�io%�q.�{��,�~��k�o>^,or��Ci_o��N)��EW]]vW�o{
�H/w���,����:@�0��<�i�l�ngt��yu"�6��\e��v�8��$z���Syl)
Ҟ�0.���rE1g#��}S�E�E�+9l���O�����u���T�^G�C6T�gcs��Vs���y��S��N���On�~��V^����~j����Z8�߲zWh)���^����ݯwajq�VJ�vu��BM�x�5ſ{y?��\�nOA�7}ƨΗ���a�S띋T�#��5՜n�r�R�cX��ؾo�!Ovf-F�3՜mǝܬNd�w�Pbw���J�%0���jym�G}B����;�!�Ύg���T��ٰ��P�65�J1)p�����t�+{�Ut���������
�����u=�݌+��@�L�̹��NY:c;�Vn��b�N�����I�޶���e9F3��U�	dWI��o*9cw���ĳ�k-ki�SP�S�sG[q��ؘE�[��m�9�e)��V�O�E�~�O!�����I�ʙy̸.���C����k{��j�p-��E��k��-+�j#��c���;G�mZ���d6�ʿK5(M�
���%�6�7HΙ����(�1w��o��7y�ۥ�7D�b��3�ًG(��x���#ru�B֜��N�L�M���ր��tlAYB^qo����={7�Yo2-�\3(�|&�h��9:�ƸS�ϋk�\"Q�С����}ȍ7�!Я_f��*{F���Tim^gT\��Z�k�ܬ3j&6�G��<犚���:�wA֔�
��:�E��ߊ]��7��^���l�"�q�����=W{p��������p����ൕ�wW�hz���G���-qZ���˸�(W/�5.hb�ڄ�.<�e|Zƈ흐�=���:��H����}jr�9ƻ��q��&�[�����]�[cq�hE��鉸�=ʢE`T�˹��Qgd�ĺ]ojlU�����\N�syR)̉������j7-�lnx�=����E�N�+��U�Z�2D�E�V�ԥ�? Y^��͈׼�CJ���d�1:��V���\�W����S�媎�����&�S�5�6�(;0z5Ԩ��-��uq�"�mJx�U��U�o��i=s��.���R���67��u���t�z�����3���K"�mh�&q��Ԯl�S6����VՀ��^�?]ƍ�[�y������R�T��{m�Uk/��V�7}n�뿟wJ�Z.�0v_:���3o-WD���$�gK�Ĳ��erI�{߸�Y�~�����wG�����m�ԧs[���w�M����nR�ܪ�چ�;"H��Y�)��f���.wkZx��]'���5.cE���+��e�	sYW��P�c&ޯ�r�k��.;�;iuC��Uk�u��.o�x�Q������o��ܢ�
+z�-��bV��'��Xɔr��N�$�䋅m�+�:��T�%����	��	���Kk���O��t�P��v���b�2����cSa��쫧p�<�]��.�f�\Vʭ���w�)�G-3�D�w�uOZ����w/B�u�u��!Fs��ޝ�Gl�e��֪�^NVcbj/TJT�:�Z9�<�Jv�|9���U9�ݦ���ۣm�]�q�[�}���5�^���ŷ�����L�n�b��Kj�v��Xr����⪍�oj���\k���� �|�LʵG&��|4K�Wt,��So���r6����_��,��͌�^�p��Z��%ұod�s�r�[��,u���|�T�"u���>�AҦ�Ⱥ�^�î���7��������crKs��)�/��=N��k؝pe�2���/W�H|c�9sh���m���3{H^T4]��m%|n�J2j�7��3N9�so-��q)���~�W!�P�:[�Σ�e�}t�z��I�[��F���'pyӸ�/�����߻��P���
�l��}J��*%8�Pg|�}j�|����\8]���=i�,§+�*c�vtuJ�m��267�%̄�_5|�t·�_4�|;rg��`�} 
5�e|yC�㺳��W@��RȞ��Ϯ����G+��h��s��)�C7��p��t�G9R�CZ!)�k������sl�6g2ƻ�<I�C�N��m�*�b&&
ޯ�'1\G&j*;e;���X��a����~�˯��u�(��O�0����Bۦe����bu�sbRq�9��<�+*9Pʄ���=�*�|�2+�x���{Gw"�!u��[/N�+S}#�f(�ko�_>ᶺ��nL���7��9c�����[�:*ͦ�B�Ȋ��;����np�W2'��bv�'p5Di�̗Yլ�J�W	��z��I}�BccF�+�G�'&q(k#�֚u}2��Y���'���G�GΖ�vP�Cf`�i�S;�V��>Ѳm�|�K����Ƨ�:��Q��=ˎhɵ��7)Ƀ�)���,u-���Xv�|s�����}��K�gWr���Ps��_��߬s�xC��R[�na�r�����*��|�|V-�N��ɬ �Ȏ�j�vҮ����M�\<���}����v��:ym�5N�$�̼���iʫpwc���؛n��y�_K���3*
��ϖPu�.�),�wu"Sپ����#r�����sb���ې�u4��ƥL#����o���B�(V?����z+RϢ�'NW+:�XƱ4��˶71+ɦ�	.�Fd�w<��Ur�A>άs֌�ڋ�Z|��5���=��a�L�v2���47)�Q�o9_�B��Q���.�e⎡�
w�������).����97��w����8�K�ᰕ}.f\ђ%?�n��MY���h��Ő񋪧b%H����;w�
㹟M\��5n�r�-Щ����;�N��:(� e���<k �}Iء�]�c7� nnR8����ѥ�ۑ��=*��rr������=�c�J�u2X�b��
T��XxF��D��c*�0��ݴJ����ԧPӦE�o��e�rz��@��� �y�I�e֫��Y�/s_E|¡Đ�v�������j۰�:ӯ�����Z���婷�.���:X�}��w�7�ٓ��-N�N����L�]��5Jꂧ%f���A�;i;��[���Ԑ�j�p�xNW���p���)d�'&�V��8���s����VLw}Ԁw� ��Y⢺�Yr����w]{�DB�Jv%���QK=v��YT��,��oC3��q^q�D.��K�4�	�^0��"O|��H�����庘�P�C��8�ĝ+;m���Ъr�w�gg���K8tٻخ�*Z�sX줱}v�(F�NT�@���u<�WM�u����|ʂF�f�@�Ǖf�D�>��
e�n��}��V~��3���^0�l3��.L��l������� Y��9��f��!\$�]m��Q�%e���R�捬�R���By����]�������5�hwi�id���<ُ�;�l'��ݣ�އ��m���Pu�f���ż��bؙ08�C-�<wva4w��� {���Ў��m]����ۃ�k-��
��L`;b�ZB�k�)W�k{�@+��,Xc��_�K#�YSnr�f�1���'��G��m�g5T�U՚ky"��ЭE:"��ev_n�u ��[���׏5��8�W��N��}}�Ӯ�:��d^�ױ�
��4u��,\VM�R�����g�Ki�o��=R�I�����b���j��0�b�v|��:wtpR���{�f���V����E��@��}��}�f�a��r���i�BV1Stڣo�Q�=}B�̓\,��q�c�tx;�N�L>��;qb��u>���Z��a F�3W�"�[�!үCmҭףhL�K����;9�쬣bR�+����E0,�1�+)����BT�3�]Ș&�a���:&�ة�V'vANձ��\c�]��-���=�lC+[@u��-E�Ǒ
�Z�(�"��<��0!�}��ʞ����E��$�z�Z����(^�Q�4�Y|�7�Mj��'��*��;.+i��4���G�`Z���eZ��U�o5���m-n�[H�0ǂ�2����õIʤ�J`�A�͹�/ui��uW˾ݥm �ε;��];�Wi�l�sz��C[(7���Y�l���|���N������K�CSUP�;E������CSr�B(7�uV�������s����gG�J㇡�p;8qۘ3j���#SW�"�$�\u�(=x��*�.�7-��]� ���ʖ7�Q��s��p]]b��pѬ�&?�^j�b^�����%#R�1�5�P��dRT�,�(��(���"��E�V(����j��YTT--kkJ+Z����KZł�E��#mD�ĶJ���DQlbZR���h**�H�l�Z��Dmi`�a��j�,Ab���`VEPX8�+*���eb�Ҥ��X�UQTb6�F[dD�ԩPF(�U-,+*
V���)kX�B��*T�f%4�V��Yb�+[lY�U�5�#����fR�ܡF5hT����������������%lˌ���"8�b��T*Uc�a��X�����[%jEưV*������U��UDUU�J¡FT�#1�5�3�̵XZ�b֎-(�2�lVGZ�2�Tb�{�Y�I��넗ݗ9� 4�QХ�\�*L�B�3`�h�v����p�e������+�r|YBb��4+6�*�0����U�a:�u!۹�)
��ÿBX�_�_u&5��NQL��!-�	w8账�8�8� ��32�%�q��<Jj�w�n1u�#�o��f���l�yZ`u�ԙ�s��^���/�Ě���o&jQ�I(\�bŎ��5sA�o^�4���?J��ݿ���"�'N�u��f@ww��b��Uè@LG1�-bVl^gW���f-up����
����I��]s�Wî����Ժ��	�:�
ܣ\�/1U��7RK�r��l:*�*�ɞպ/8K�nS�W�C�p�l�t� +��X}h�^�ϲ�������/�ew������(��SW��m���W��ʎcr�TKBH��7�7%�5�\�i3n�.s�"��Fr�w<�sb��!P���|p����!5aɷ5!\:ͧ�χ��U]�/VJ�W��]q��P�>ؗR��Y�ץ��u���JL2��9��{O ��<�ʾ�.�<@�o��J�k	*-� �YB��b3��,��y��4����n���w&ёf��ԡEJ� Z:ܦKʗ��6m�39�swr�:���,R�ts�>�ɝ|_�w�l� қ2mwjo����+�ƲnMm�gx��B�[8�j�pN䀮x4�|�l.�o�{)�B��p����u����ꕞ�[�3�{��Y�|�Z����:{Ц�M��j��������5�;�)�=ŵ��H8�I�d�T$����K!���Y�y:�u���eni��ኰ���9Ǒq)�*f�+�Me�0��i&��ږ8Ɋt�o2YvQ�u̵ָq�g\׵�����.w|���7���	��h7�����w�j�(p�*���T�"yV����_D��w���q>�p��ʾ�ٻ�Y�㚑��NhV�¯�ؔX���ߨW<�X��iw�PT���ޠt\��u9��K8�[�����}󗐯�@�$����׃�U�j��T>�[���o�e�-/��Z��I�r/S�P�*��X�XZ�3�E�glN�����Ti����V�7T����b�����%ֳ8Z�6��A��&T�ڪ�U��@�d���)i�4;�V�D��Y�7��I�Ir�H��HX�j��\w��[�S�ٚz�e,��$�P����u���W����q8�~Š�ݩ�����WR��y��P�����*���)��������;J]��11=�ꉈJ��mh|7%9�0.�Ӈ�F�,��=������O[7����z�����g(ןs��+����/�i�3$����}R�ypN�+%�8��8s��j-C$��7�<��io����W��|ک�7�c?z+�D�W�lOC7�<����=h�{gF{v��Pk�"N/��z�*�t�[���2L�x˽@����f�!��QP�;�Ք��*N�=�����E����lE�G�@�t* �Q�����!_ǡ��u�Q|�Z��|���{����z�bV�`ĹWXc���6ohh��E��ި�3�Q�e����CM#�\����������]�֌�]�7|q��[R���9�B�>�^��!Cs��~�3����_e���� �^:��a����d�a��Wq9�n$.T���I�w$�S�%cs��/b0��Z&��!`.�����Sn�0,��k��P�[{�xJ�gl�`�55 KrY�d�T瀒S��]kT�z�Ak�}�l�ɝ�u���3��'�=��t�'.U�����U��-e�lP�&>��k״�on;3's2G)O�iN�3�:��U�L"� ��w��j��F�dkbwnu��U8�9eG&r���p&BW�wb~Lp�ڭ��~6��ዽ�sNT�ʾ�d�;emƪP�UCNOb��F����`U�fs�U���o�74o��R�>ab�=���:�����u�C����]���MJ�O��N��&5���s��U��ڦ�/6��{-J#k���w��U$�o��_kjBᶛ��`��6����ު��qK�M����2�e�fvh�Ƣa�4ţ�?c�4����<���:Ƽ?V�]֟>��]9�ˌQ��sڌ�l\(z5�{���t[����Wc�nT�=�m'��*�ej�c\K���E�u�K�W]m�$ا����ߛ�����Y2�oeO(6�%d?-	�_�W^nh�:���0�\L�q`�'@G[�n��l�;���a��u�:�[=KI����<��oE	,�g.hi_]��{i̎�״r�}O�pC�n^�y�r�9,�7�D'U��Di��\K��^��s������Z�}g����j+�5����;CT%�;�K170Z��n���W��������bw����-Rw>y�]u��x�wܰ����ƛ�S|�����L���R���������CZ�"��[���|�ni8}}��n����BU�{"�NfN�lw<>>X��|��G<���q�g�=듍Rq�N��N\��ʘ���*H3uW�p5]�Jj��������Ħ��rx��W�A�3Fw{��1�)k���a��6�A����חfpW�5���g;�\�)��XK=Zweb�Iܞ:k�<o:\��o3�U�i]�+�v\Ӛf1\�vg�[�]��7�� v�5�^@���b9k�4���:���Z��&�6\�X�U�v:���m�������p����`�^��K��b�x'�0�d�	
�w�R�&㕞���V��1κ%�>nd�籲1��ـ[���X��{U�
F����vCj� �_m�Ӷl��J �Z`26�<��xJ��zT�:$J։�Fos���.T��bw¢��T�6�cV.?>�5R�{�ܮ���./��uN��H[���؁wu�%�Z���~�d������zr�7I��7�f'��L,����p���=����`����e��Ց�7�q����vTw_\�U�ʌ��3�tblwΖ�_K�һle�֧VQq��c2�C�H\���YԸ�������W���u�tȡO�����EsI�4q�;������'`>jQ�a���ܡ]�>��3K�^檽�vH�{��P;J�5�δk�d�|jtV7�jٜ�9N2{�z���������5����5�&Pt�
���"���s9��?�ܣѝ���ʭP�K��I�}����:n;J]��"�6����!re��[R�9p�կ�p[��ɥOF�\b����LD��5���S[U�,���e|a)��Ϯ���֪%,��6����N�����]h�v�~h)a]�ǝ%6������W\�TZUlcn/f�^ �"�} B���͹C �t�k�7�H�^�Vo�i�V�r��'-m�N�q�6�;+X��o���M>�C�$wη�\R�)pC
����#'�@�V��8�;�d/��B�YY�Gv9^�mƻTG{හsȮ�Z���ˎ)�rzg���<����r0%Xܪ�\�7p�-ؘE���!nE0enM��r,Ugұ��H�s�{*gV��Bw�WP݀��^�A��Ȝ����r٧Ο�����y�����I�ܞ[ɸ<�z�1�u��bа$9ޣ]�������[y�1��M:���B���CyLc7�*ˆX��r�'��E�����"��2�m�j��^}B���d�~�ڨi�����Or��ZO.�V�R�F����-��<��N����;M�T��bo��~��vZn��{��C3W ��m-�q�9�.��+2l=�vIѵ37W���}<�s��ث���j��g�$���x����8~`̿o�q%�ݸ�`$�8��cڄ��ƚ���mUo�g�ͺ;^7r8��P�Ckm�H�)e��YyVeyq��̇�Y����[}{F��}�s����m�]�A���-�$>i�vu�2���;���z��˦�n�֎�K��Ӈ��u��˷'v�Ҿ{K��!#Urw.�\�9}�"���2Y��9��'�k���w�;<��qַ"5��S�W��l��Nu��5)x�b�㍂��Y����R��O�sV�v�uܓ�<�@R
����^7,oS�כa�z��.d%�3���0�����y�+eX\��'�K�#_m9n����G(Բzf>�\�C|�S�����$��9O�oq����О�W�6~�H�D&ʡe|a)��Yw2�ӊ�Mnf'<��u�]-���Χl�i�;���B�����wp�m�q��v,z���ܜks�.Y�9erg)���=�q�݁yyK[L8������}"���u��vX�x���V6�12�Cb�hŭޛ�հ�%uV�*tmaz�.��UoL�-Qܝ|�,�����N�-=�v�8��;Q�)�X�Ցn�9;~��u���PL�U�ry��4	ё�s���$�o_M�T�,�A߬�}K\2ph���+�u�%�����t�������jf뎟a��b.R�B�Lz�w=��_o`˞
:��3�SF������e䦩�B��9�(�Ė���P=8��R�S�ʤ��8�ک�kk[vUO���f��]�=�4�ۜ��Ǿ/�)ll7������zj!,_u�ʂ����r��U��&����rz�/m��P^�w�絉�Qn��7�����4o\��ButM���-�mĊ��-ħ1s��=��Q+Ÿ́����q^�t鬾�4Aa��8vZ�3Y���3�o��'�"��&/�L^L�>ȭ�����챇}OM�X�r�H���DIv�|P7�}���y�p�g�9Dl�SR|�0���~&�]㻇���C���Q뚾7���ԢN�z+�mzޜ��am�_�6�Ô�{!�f��x��)�@��}�G��u��k��Ï��pY���d�l�O�������;E����2� ףg���A���<�����㳺N��!W�9�k�ه��u�;�0�W�܋^�t|Uht�1b�w��(���(��ڞ��>�� �Zs!u1�k�*�U���zv�����y�TL{�>�ܓ.*.�(�+Q�{���D��ZF��4��V6�I�aU��
�ژ�y١j�"��@Nfm�Y���n�C��Mo*ښ�L��wZ�n�x�)v���E`_ ��\������K��}&s;���[�j�Orӗ¹���Mk��������k�����Z>�ҕ*�8��T�W��l���ŷ>�ǽ�w�\����7�MJ���w{�����z�@w�WO�'����50��xLM5[F���%�d��U�Wy�3G���r7��/�>��@yau�x�P�2���L�޳6��ۅq��������W'�
��T��=��z��BJ���	�Ng���`R9m�{>8MD/I.��nnP��N�i�G�����t���u�n;��jo:|=~�fG�z��D甞5���q����?�z}�������7��*Ů���]�^��K��z]�����n����`'����@�����VEw��+��D{unOv9��f=�{M�����1��ZP���ZoS�;ګ�r�~�"�=����,Ѩ���{
���_h�c��_�_�e�H��:�X;�d��UC�Y[Lf̟�r����bO�z�򝒽����i��^`~�>�����A_�t��v��y�R��Kzd1��%zU��_��G�������������r>���}�|s}/���/��ի�Y�PE^��c������#ё�]�����S���S<%���*�yJ��4��E0��]�տo]�Ӧ=�5p��ƑS^u ��5mi�'v�Mt�Ts����z�I��i�����k"m��ξX�&[�DW6������	�a�z�RkKP7�[�w�=}�j�:V�p��a����a�t�b볓G*EM�h�IC�&�-4�0k���0\�f u}X��{˶�|�W#Xʾ���1�Uǋ������z��\�=ћ����:�f��S0�d�B�
4��ֶ�U���i�"�{v�A�z��q���Ƹ7��5bo�I�0g3x\N�CX�LY�sB��t�Y�S9є��WK�:�Z]������s�`X4X�Z��ד*Y���p�� ݚ�@gK���7'V-�mN�y���-�M�6���:+;�CS][�spq�e���A3��9f���]�R����#�F���_V	ZQ0���"���K ��̣�
�M�8ed��K��_2D�D�^�9Y����(a-=�*}���9�B��
tf��V��V����8�
�p��)?��L���-3Ot��h��p�[��ب���嬔�*�c�3%j!@�N/��ҟqX��n�5����]�:T!.�(�x���Η+����a Fh�G&T�fjs����PN��/,?:���>$ rY�/��[ب���{���D7qb}j�֞�Ѱ�H�ᪧNژƘ��Ut� =���8򺷟�K{�uV��Ψ�{8\�Fh���L�����W�r���O�t�t(l�y���+����l7�k�d������f;�Yj��9�t�Q�
v��Q���]�r��}x�)<�����'\�����AΡ�?���g��n4߸ǊU�\��\ppaP���R����� ��~�%,X֭so;ZX����%�0����΄���,�H��������wNWh*r�b��Y�m��1:Zzl;B�S�������[�&5�EM]f�[ؠ��kx����Q�۬�����h���qa���mtg�����U�|�v�.�r�F&�Q{֠+)r3],Zu�kc+Q�*$�;�)��RPX��;y�4�1r�n�#���]�ÈZ��r��jwSw�mF�xk3�����*gt�V%�\s��^NU�"&Gr�F����AX�QC/��@*��X4�5nu�XM}���3�׃!yu�8QQ�7��N��ެ�v��OLU����.AK�d=6f8��m��֦���,4�'eCԭT�}/%�vm��I�j{�/�)q�	�� ,5��x�����u�q�^��%��Բor���:�?�I�:@n��o���|��[�Ns�	,K�ڙ�����d��)�9��V��"�6�mc5t�/�uh%��>���7E�R郕�z�7	n��6��ÝR�ƣ'lC0�N�J�j��է Q�5���ÂX�K�hٓ��m=��Vd?\�ӝ��uM|�ͻ��,�{Ϸ��TX*�jQPE�)Or⢑�YRŊR�b"�X��,�Lh�F#r�Q�Q����*�QDPQeh,QLJ�#��`�mic*�T�\�+�1��U����hZш���S(ff"�%-1
���UTV*$q,Ee�cFZ��"��5,�����UZ�DXF�FQ�����mj8ʈ���R�e�UcZ�*���--���*����E1TUDF,R�
�*6�EU"ň��#�Ab-�AU�+�("�ȱX1`����T�A��ETJ��E-�-���F-e�ҋj �%h"�����j1�B�Ң�Z����X�Q�F
�,Q����A`#b�H�,DKh�(�E�V�� @�u�Q��L$uJ6&%�`�kh�9E��d��@�W����mnF3듵/s�S���m������ZW��(�TfL|�_������]=�^8��=�=9�����z�7��8�q���Єd����S���п��T�����7�����tB��hz�s�=K�F�_��G���y:2�p��Q2�\Te�l�3��= r�wB�l�q��Y
��x�������s���3�ըw����i]�
���G+=7��ޘ�n�I���K[��O%#BR���<�;��+��i�j�@��}`s7��"��P��\L��jИ�}^�G3���I@��6�_N��>�Ei�s���v�<v�_�~ <��~~����9�,u}~�	���38G��/;#Vkn��-��g�n��y]���<�K�_��I�|T�|8*�����f+��	�oy�>p�O�~n����F��_��s�������>51�j��>���C�$���Gc�Do���d�}%qwt¸�����'G��s����|������\_���'8_C����3�����턤㫰�0�\�1��+ğ#�����X�͚�n��5�L �z�̨�h3`\�����U�{O��3�hа+����6�=s��㝂;�r��yr���Ԡ�~�ݙkϫ޾�,�%�˹Q4����$��z�9���I�̔o���c0���V���1�4OobvZ�}B�ȧ)Ir4����3;po��I�zM��K���(g–��~�4�گ��S���pg�{^A~�^��`֧@w���;��lzt�����E� z3��D�c,�+c������K$�ۙc<�"�Q��k��ܣ�W&[���:�����ϼ��vk�����x�j��F���|3�-���d�t\K��wT�{�y�U{4��ݝ�G��7�øɝ����x��άnC/��;ޗ��;sơ{��-�����G5yΏ97x�<����;qT���e���O�!��ϥz�{ l���|�\{'���{�\n���Y�;ؔ�Q�1���e%����}M�Mo{��yU��u�|0�����
����3�7�����i�G�LqN��+.���C����9_�^��D�a^/q��Gguz6�M�L���kUN�gJg�y	Avo��~�S�� n{�x6ezU���s�3���uv�8��8��Gќ�F��$n�����xW��z2˓�G�f�z��w�k:�Iw��H/h���9��ݜ�3��y����u����(�� 5�)̹(��������u���5DWO*?7:�zڮ�~����/Y>M�Km���q�B���&�a/1��[�3C"����e���r�r��p�XV�A�vT��y��.�O%y��;7 J�1}�Ŷ�=��3/J����L�j�(m�Q�i�����=�+�߾2ɟ���td>Ӹ�7�&�7��N�b����_�@~�T��3��n��Z;��b|I�N�R[.��=��W�b��;&�5Ώv#LjsD�o�hOo��\��Ǟy�uw��b��K��
���;%����5q��a����3��]lxwn牺�Vc�1bO�1�w�J�G�z3�ܣ�ޠJ�ꇅ���+���r�e�ۃ���OA�y�X?�ҿI���u��&��������z���y\5�{�wB�����<o�XZn"vXΕ��Ľ����Ow�qu%��BuZl��v�/؉l��W>�p���n!�8it��|������סZ�)��>����\FMiW��lr3����v�W�Q��g�����7��+���ѽ++�=�[0q_e���xя<�ܩ�z�*�xgK3�7N�/'���>�"����=ӷɶ��4�i�J��/���o��j1�
D�d�`	��S3�ӟV�By��btN(�Q�3H_k�k�]������7�6{b=����2=��Y"T�����W+�8.��MD�����N	�7��)Ϊ� �0��Or��}g��m�ub��߹>����]U椯N�b,`fhm���z�
�qʷr֡�i}yM��ܛ\D+m��X���~[��Jw�:�v##Yr_l.��h%�����:�_��<g����Q�E�K�s�T�����ez��{�������b�+"Pg��j��;�tX^g����߈܊>��gN�$� }
Z>܏u�F�{�=���9��O�㾃����~VԲ��@l�D�7$V�k7��a������e���'�x�>�D<K"���0׊�Ϣ8�������>�
��U�F��<�/��5���ǽj�d>l�\wzX�{�W��zc=;\T��v<��-��l��H>�V_�ĺ��iG�����ꋤLO����x�9��p�y�=�{y�l�:��Y�~Rs܏�v��Ku�5���|�%K�L==��m�/Ǻ�F�]��t^�їܼr��8{}f�_�׍�~�=�M���	!Brx��c�pf���	��GO���^gb�R��oJEYH�>~�^�TY����*%��{ <�J�(����z[� p�g���C����;���Oqh�+:X�罻��~�>�Og�컏g��#�P�D� ��Y9��zW�ޣ�O���N�y�����Zou��g#U0)��!����#Ώ�l���j�2�L'�}�X�����(b�b͘*��uK:inΧ�@�uNק5s��7xID>�K�8q�����o��Z�q�;ܸ��f�p�o�n�fY�G(>�َ��� ��#��IO��z�s��luJ]�M-u���=9{�֋�8�����A�К��^�տ�y��w�D:KGn'i��:P��U��� w���n.�x��À�~�cw�(�u�bg�����>��Ar�0w��qp�N鸒��Ló�em1��m:\�y�~ٞ�Ǽ9�c=��l����]���w�t���-��IJo�,a鿨���w�?Mq����t9�-�Jު�uo���y�^9Ϊ6�������?.�XTG���3��^H�e����r�0��&�������|��U����~9/���;�����L�}g�Wέ[�(���b���`�v�,\p��������*�����7�V��1Y���s���7�{��n�[��V�1J�ҦZ�۸�[��n�Ex� rگQ�%���s��!����.!�;a��T�:��Mǫ8�Oo;��T�ސ6���!���=7>7=q10�EңW�aωh�1��9afmL�S�����x�'��'�f��ur>>�@���o�$g�Q�v�d�QhLLS����z[��2N/_ݹ��gj�W�}�P�~n�/R���N�d{����!�L�*e�F�`��%*���? ~�����L���Mֱ�:�]�mwZ����u>w���˥��Uiɸ2�~=e{�_P�W( q˧u~T�y��7�`�ys���Ł�m��c�Ԑ�9P�1�k�����Y�DL�ټ[�vZ���'�r���)\��������/�Ty�Sq�-���/7�Q�yUx��v�߽[@;�*$��x�3�ˢ:��7^Ag��X~��q�D:������Z>ҝ	��s�����t�yw��2�������_a�7���� w d~�8v��Ă��c�ku�W	v1��A�?I�1嘮&����wzl�]x���ī$>9���[�/��9�4�:��[��E������#�h���̐����}^�]��	���<j	h���C�q�W�U���S'�d�1��m�MzEw���*�=�'|u�7�p�D{������Z�:v�X��K�B����K"i�o��wH�W�w�ٹ�`o��G\k�����8�w�Q�Ty⸸�vQ�k$��n'� =��я;��^�{�U���D\�zb�r9�����~��^���;��n�bF@ݨ�E˧��~]Z���d���M�x�q�T�vJ}:�Í>������1��q�^�s���co#t�}v}�W�|c���5��늦�O#�o�)�{S��#�ҏC�,nի��=}/|E�xާ�vV��VfqU���rq�J�)��vHj�.��F�QT�.�C2w�z'm��p=�� Q��F�%�9���1�m���f�na��lYl�@s�����vS����uVY=)��Ht����]W;�G�s�����5�U�]�Y�|=�-Ͻ�X<�b�t+��!T�����k�'�n�7W��z�*��'1���֜�w��x�G�ޔ���ݟk�4W����/!U ��BSD�H�zhb��˙2;�.T�L��6��=y�cꂊ���\S�RE?J	��D�S��^����a�����.�eV�΃���Gg�s �]/��{��Egޥ~�q/�G�8}�� �Y�oF����
���8O�Nx�WQ�)�tdAs�;���߮6��W���ȣ\�
�]���������Q(���*���}q��bk�$�ا�<�c��t,�]��=�vl��*� �N�uW��5Bzo�P�@��&
�>���}y[�竤�۳��Ѱ3���ν�U�r�ǣ��خ�E��y�p��c�>/E_/IG."e��3���Ss�������8�3]r���:z�&�n�LjN������F��˸|M���p��G�7�Ѡ��W5\�s7����~��ɿ����9����lt{�̢s�}ƾ�g\O�Q��Tl�������
������/��Z�P��VWhöqS4��aNGm�s����\반��=�����M	�t[c�%n<���ҏk�HN�W>�]X�k{�H�v:��ٕ��X)v�9��9K��av�`�J�"-f�d[�
��v�^!�4�.Q����T��4Z+[���r듨���[ο �����X���ҭ~:�t7ӎ�xv|ׯ��N2��ޯ"'ngЀ��d�xs�R}���;��D,�񋇂wMě�CՓZX�w�%�o������!�aG��>��C<7��(3yR���i:�Q��$]Ǖ���}eL�>����4.H�SG�ؒ��č�F<���;�u��ǽ��ðc(����鹨@Wz�<��;֧so&�Uns��r�^�]�$r'�W�ާ�#�,.�~�.b�3�9E�d������k#�£*�׶ug"����\�n׼^lƣQ��<�-������v;Ӣ����pVT����L]������&�����UB�K�p��q>�|�\M7�H��S̸�H���F�x8��ŋ��}�x�}�U�P�0Pʉ���zN}�B���7�ԃϔ����c�>���T��տ���vy�H�Qc��Y�,��\���Qt���)�{H.��!���2w����HK=څyY���u~9v�7�h
���!����f=�~��^3�ߖ54zf~[� ��q�t�B��ez����T��?c�[PQ	�q��""Ku^��ܱO��ׇ�g\�X��Ұ��n�
�q�#���w�r���"N�ݮ.s���s��x�S�)���	}�[ۭ��m���;����^7���l���X ��";��:�������k��=ۦL��^�U���Wϧ1z5��>�+���}���ǹ��7�<�}/.��Q% :��+���"o�y.�9]��l�n|�mh���wO��]/����.=���r��}�U��� YWU_��'s^,����ӟIC*r��?��&tV�?���`Ts�dxg���>�>�8�y���J��e7���k�J���&����i��8r�T{
���q���^HV̯TT8^������#���|�oG���OxTTB�]��>��R��*�:u?,�F?^���x�Q=����`_y;�q���m��v����z����B�2J5�ŝ�������G�/��8�^�̾�z����م⧝�c~����_��]F�K���'QY J�Yu��4W����݆��1`�&PY����e��t�rS����[���z_��|nZ����CQE�˶�����6{�@����9�W���N\�H�#��~�=����hu�i����u�MD�x΄+��,�h�SW��?v;��p� \��ā�����26�_s�ʍ�wK�kVk!x�Z�)&V�z�T�ֱ��-����W.W��Im^1W�zٌ h</��Qz{+#Ҙ�xi]*�gm���Y��â
ˊ���i�v��}�����Âٯ�H���j	l�o�˅�GW˷؅�s
T�ָt���|��R3�������޷������7=s0�EңW�a�%�����P��u�}�ϺJ�z�wz;�-w�B�N�9�H��4t_�����q�̀�k�S��/�=�k.v�3�ri%��-�T{��_���]L�=Z ~RC$�=2��w*��\Iyv�߷>��ޢ&"�V���wNB�zm?����ߎKG%� ���$�� X3(�'�~�dY^z����fP�rG�.}�Eju�9����X��O��.;���S=!O���=y�bd�����#���P��	�2��裭q]��Z�?"�<��J����V<2@��βL^�t��h�s�)Ǘ*�7�c�QQ����_�څ���1W��;�|w{�>�½,gT^�����w�f���<���6�������!{ۘ(g��8*;�t�Ķp�ó��K<��}��2wȾ��+���%(w��V���l��=��Q���`�Iӷ2�x���d7�}:nVWPZ��;�7��]ǁ��ˣ�>E>VG�hf%�M5��mZ���5g.��i\o�r0q"V�J��&����)u�u:G���7��n�r���ȦlCi�;�v�^ֱ�E�:=�qg�H#�{D���!���OLF58�r����Q_�N��B(��1a�F�z7L�N��&�qu'�`Wau!c��Y�ktu#�3y�7C�y�R(}�59H\R�e�/3oF�jN}���o0N��;Dlp��s�R�qz�&���`�VrT9ׁ-��% :�۬9]i>��I�g,��irAUt�'C�sɺ.vd�����7�ط��8��yG/�����:3�Y#�Y6�3W���x�<qB�v���m��� S�4q�J
o8�c�w\��+�-t������Ӣ�ӌ9���"O8*�W1]�H;�2��w4�I��w\�
���0T�Ui��yݬ&�����K!�	x;l8p"b�O2�����C��jzemz�%VS8��t�I�g��2���gؘ؅�v�1�Z�;o�D'v�W=÷J`�)8���Vr�+�u>�*�n�9��t���I-&��D�Q�@��]	Q�kw��ХX����Ⱥ�lV� ش]��sP'{��Wl�xp�v��1�[�mve6�-(���nnE�BU���7��y���NT�Xd���:�}�z��!u��g�7#��2�-g_�ä��Y�F��Kmu)Ѥ5ř��%b�qٝ�e�;gh��Ջ�2��̳$ö�E�0�EH�%F�gn�^'�fw�a�4&�s) 3kX�hd���XslbK	k1.[��̔�q�Wg�e���+B�gS�7��g>�CEgv��ׄ��JT�]����0}5#[�
w��Ԭ�S��ق��rHu�]�>{U�%�n���r�61��dں�A^	�tݹ/��6E�+���!%+��0���m��N����.|�0z�7�ހ�v��OF��k�r��YM�.u��
gE�Yx����n��0���mq�K5eLV��..��΂ȡ}�q��n�pF5��DL�3^�]��Ǐ �WM�9��UfD�V��QeR��t͵�{�ō�uצ �(*���q�=w ����jcYG�վ9���s�v+�]�Qѫ;%�54(�!�_H�`4��I�����G&g�_HW'{�P�J�%`ev����f�zoq���`�
���˨��n``b���r����r
�����n�;0�����6�%v9]e�q�X�.k��	a�R%o.�ڛz��,�h��g]�o&�SfWY�7����>�ܥ]Ozw��)
���)e�Bj�[	|�\��e@�bH#���VdS�{�p⹊?*����;�gm扯�����y����
��#�iV(�K����A���QQ#UeV(�0V*��X�֌���Q��X�[R�TbE��*"�،(�EDb�R�UX���"��QV"��������UUEEPUQ�F�6¨(�
���$Kj�Q�"�+*)X�	���V
(�"�[D*"
��"���������B�T���E�VT��"�h�*�Ub�(�" ���Z�b�"�EX�,D��ZV#�DUelT��*��
��6֫*)F҄`�A�DTPAEX6�V*V#0QQ�QEA�e�D��V
�m�[#iQU�X������"
*�(�E5�PX���E����*Qb�)l�+b�(�ڢ�j*�ED`���T@�P�
(P�(-����=�3mVI������o���o���se���3G�U�#�v�a16�zC�R�;ޛ���jK.�ت�ĸ��p���Ы.=�.jz4��pת:�W���G�V��{��MTT{r����s�0x����TK"�(�9�=�C�o�8�=顜߯����V����kC:W�R#��|��*�i5��YE� w�������K��v]�d8��pC���ZP;:�Jz���CYG���㱪,�^D���z��`MO#�o
e�C۸��)�_158�����=t���pz�z3��Z=��^�]�1�¨�#�@�7�&�"i�D��T�ˮ���k�v��Ƿ?}�pY���#!�[7�����X)��~\���ܟ���7Gn�s]��G+���x�W	�i��F�%qW�i��A3����N�?���E�ו��g=,��5w��*������P���3� ���.��q�7qWV����J7��?q��fq�Bxz�g=�n�@���ԕ��jx�G|pis�;����=�+��-�7�_P��~��iF�fv����)�D�����"����/����}q��bk�$�)��!,c���
���Qf*�1y���\C�	���
8���_#��vљ����z�͡��#λ1o|�`$G�+9u��
�T�R 3�]�GJ�;X�� ܕħS��'�ce�@f�fԾ��:��ep�CR�w,�⥉�
�����Ns�޺]K'8�c�1��o�nY[��m^'Z�'G�=��·�����=�A	��D�>50�~��0���t��ë�U��鵻S����6�Hx?P�9̟�:�{.ǆ����(�̱�fax��(��ղ0��sԝe�X󏢽	W��t�MgT1�߯�>^�-I�:{�[��vw���r���Q��K���dz�3�'�/C��s��>S9�Ը���ϼu�Mǔ�5��:�k��G�.���B�V��~,�a><��y5�\d�PZ�g����~�q��g��F�:=������5`U�	l���,��[��.	�7&��=��ZX��g|v\�����V�����uݼ��;����#�y:l���ˇ�<c�0Oq�+	늨��1��>]s�TWv�ߪ����p&n�}�������Sӟ?:�=��n���9�Lu}�'��K�f$6�ߕ�����[���۳�}��P�n_����ߴ��G\o�Å�)W��
r�/"�;{��z��77���q}V��s���5^������[�Ty�l�O��89��~�C��|'�=�ö����'պ�X����]�nj\���=�jK���7�Φ��<��٦<��ɘq�,�ăb�D{A�C�l����+��\��[�a��R�mA�]�ݳ�g1q�;�o-�b��]�G�,�W�ꮺΛy��IW?(s� gu�y��.�o�=㭪��j���H�~Z�WP���6��m]/ך�3Ş�n�V��|!��w10�]* xu���],{ة
i�+��+W(Y6�yu��K�c��\T��w�!g����_��t���}^ӄ�̧����&g�곒�w�o��y��ǩ�ѿ)`�B��@y��%�OKeMx��'Ƣ�{"�l<�ǖ���-�&,oܼ+E�~����@yau�
�z�I��je��̈���9���G��N�{6=!��������>��-i�N�EG>��9ޠ%���Q'�Tv7��h���	���]ʼ��p�7(;���댝��,q���ǯ����/U(dyI����&n�7q3�|Y��'�m���g��죇�~/	-D�1����ד�����ϺX	׮�y��/õ+�O1����X>���m�D�>�f��,�)qȱ�q~��_�����Y�N�CJ�2�ߩ�|/��2�.���N�]p���P7e�%��eT,5�-{G�y�\�բ����\:�����g\=��1쮋γ.̳޴q,LW��MY�{��6r���pY�)�����e�4[��v���ݵ���OnK�{ɵ�[g�� ���%�E򖔮��E@��U�j�+خk�v�E~�?����g�Uo-���5��z�Z7��G�i��A,Y٭�U�����ӻ�UOC[U�d��}�[P���w�߭���K�}����/Z��mU:����i����T�π���tp52��ury�t�r_�=h�����L�9����q����>�^��I��܆����������]��Rx$o���h{�3쫢���4G���e�ͣ�֍�Y�y��s��ǰ-�f��9\Uz��N��h����Ո��=u�잍\�w�P�jN�3�f�9�p�{������8�ވ���.����,..�d���έ�)c�:�a��w
}>E|�ԁy�����R�G\���d���7�K�N�%�u�%��2��3�ЍG�o�y���OS����0VG�� =�67�2x�"���d�~]�Յ!hy
d������=�C��=�O�D5�P��U�g���9+(�]��<Gf��bK,Pdh�t�;�MW��c��i����x�7>p�b�oμnbj�sf|3�����Y��yn��m,����ŭ'r�����c����R,�8h��u�ړ����6�=��K��C�O��#X˛�!�����eu壑�����;o�ئ�ٮV�-;���xy"f��J�
�J��C�LD�޵,�PE�n����C�Y�l��=U�a	NVE�n�%�������&��=����uQs�U��zMn��jҶ="w�7\��Y����E_�p}#�=�S��}�mX��DWxJ�C�;P�q[���^���7��	s�E%�YIlN�A�}�hK����^�-I�7��˱B���Z;���e����C��y�q�&sT�T�YIjз�/E�!s���̩��:� ������:�J������]r��7�?�!b��ᓯ�~��>��2�+n*����s�@u������N3ݱ�\r7x�+r*U��n�}���<0{�䐴�D��z�Y5��L�/�wL�w���7��;����m�WA��\Ѐ���5��wgڵ\<��l"R=.p��`O�=���ҫn�y��?x��UW��"��yN�D�]�g�ǆj�����έ\n{�g�F��5��"��*�<����}Ǡ�����&^�&�y�/G/~�(t�ՁG��u��×�m��j�B�!��A:x� TN�����.�,n��';PȟB-�n}��#P��q�~�ˏp�#پ�4?W�Ô�^�R�a����&$P�rb~��P	��FP�tL�s��x>Cז��{��h���DU_)��A���^�\j�z!�<�>�z3 �p��ib�:����s�N���y�댰�r{қ�����[���o/9�ެ/�+e�ʬ@��˨��,�%v6�����U��N^��R�c�1�S�[�y>Gۑ�
4�+��j�����.=ÿg�F�g.	�Ȫ�Y� ����' �O�`�z��P�����ә������*����|Nq(�=�9 �b�W�c��u�XXþO,��2�n"O���.�3N{�FFϩq�X��Hyy�_�lG��\�r;�cЕu�L�D�tq�d	s�Q5��ʹ���>&6�����n��c�z0*.cr�������脪��C��r=ҥ�G�H#>LN�'��"�v�k��{A� �/�|/uzwU]�t�⴫��g�O�B�Qf����C����N�P�%%��⪽S��;3"�_�Xtt_`>�_��Bݨw��7�-W�u��{2�2��(�y\5�e�zɳyG>�����9��3��c0�����:��'kf�e�)�������6=:��K32C�5{���VF�.z'=�Q���J<3Ӵ�^MiX|'�t;ӑ�î5����4���Z[`��*��Ӏ�uo+U��:c�¤�>YT�VMib�&w�e��{����=k����Dx�U�ɚwu�Tҭ��#j��3�c�+}�2���S�k-o��,EESbz��l�!+{TxWT���ot�m�U;�`��G��Z��3qVYxw���̮K%���9��K�@_oU����㶒�	�Z2zj����r0��^��H�y�#��T{�����(��`���%�=qUƾ�t���5�QR��z/R��/�:s�mT/\�f5���^�י�\�ruv���{E �be�K	L7MrE����|�e4���y���d������q��K¾�Je����jX�=E�}�aM֒����ngxW�����x)������x)����,�S��JF��㑮}�r�O�j=b��pv@}y=�=;��Qe@̌ rQ^�\�M��w!��+�M��1���uÓ�7<2�;���Z>�zF��z�X\�O=�q�h;�bW��^6�|����Q윊�3 �1�>[؀���s)<T�3�4�wPG�3�(�_s�t���}^�ک����~�6����������a��6P�����i�����fA��DL�*���S$��V���J��]�GfNQ�il�b5M��m��u~9}� ��@�b�~%��gǽ�Lv��|�<���`��60m�m��[&�K��9ϸ�?X�����ٸ���r%��{��~�E���4v����fPĖe���>�v���ql@v�=%D���WW�o�RA�3|���]xK��߸^��]1�p��+N���^$�Jn"S�Ǒ=���m��oT`=��<F;��o	�\�$�uj�F;j��][-��qN�f�w ���Ѽe(�:U���V��Owg����ǟ���$�ϥ�	���V�3�����W��-�TO��8j#��/NI�;q���X��~X�X-��iP��'��=>���µ+��=���s�:<}�4+#�h����B#�#$u�ϴ�м���O)��=>�T�Y�|w�O[��W�$dG�[&��~%e��mh��wM�x|��xgo=��*�f{y���]�Gz��� g����Y���o�l�{W��t����H^d�t���	��ȿ_b]�����u�T?d��}��A3�O;��e��Ǽ_��E�g�|ߵ��z;��ͥz;��cٌ��@+�P�=3�2��
g�k�~9��U�d�-9�/ţ��:�����}5�U⩖>vvkj3�{g�dl�(��ޙ`I��7�������Hy燦��z��o��w9^�<=��]�w�)���\�,�p\�= r��Q���+��Fn9�ca�3:s�eQ����w�^��ؠ��L8�!)�H�{��Q+�a�7;L�neI�����z�껩���@?�'u��{�HbV�s�_O\�T�����f}��\������m� _f�ِ�mc9���/4�gD%:wHK�8ݾ�b�b��%h��Hh�S9�f����X��v���ζwt��GBjv��KEcF�^�[���k.��������q-����p�ԑ~�@��a_�N�_�Y�W �}9G�>�Ȝy����f�ldx
g��Aޯa����m�\Uǫ���k�^�h��e��bU3*�9.EW����z�{�$�a#�ï�Q�i��S/M��7<��|>���]��M�N�|�&��ʶ�yd���J Ǹ��n���=D:�ZdT.u�)������]��+�L��}WE�M��Σ��s\�yNK���I)����{O�EH�Ms�z������u��!"˗E>=뭼�)ǣ�����yYy���5��ǲ� ��*�Ė2��^���L=[:��<�mw�m�����f�������d/U����eءy��x�DL�vQV�T�vok7�ӆϗuG�6�N��zV���{~�N{�̣�����R)�+C���gԺ������ǎ��'9�q6y�.GW��Mmm �@�N�6����F���>j���'s}.��Ez9���F���=2��������<ˉ�U�Ȇ�~�	î��t_�[���+�� X�vbU;\UÃ\4�܉�����3k{�"�6��Њ��Ⱦm:ݘ��=��;؇qOS��������3�^��2�3��s+�s�	�'V�G$��NM5�i���C� H�Y=�ǧYw�d;ە{��mD���ݗ��L~Xḏz��v��F��)̓�,��/&u�r��R�]W����/Uvo�+����!^�S��s�w#�O���q��G�9DlL�R|���EO#�Ik}��9�3w3�*�gJ����^j�Ϗ���dA�z�d{��{�î^Zb��!ĺ5��]r���S�5GP��Խ�i�0�Γ����F���|�|�=����w+û]�~����Dt�}����>qYg<+��l��5>%F�M
)��Z>�}pQx�Et:��s�~��g>�D�Ί~����ŉ���k�]k�=ʺJ�@�ٿ��U
����}�X\w~�~5Į*�Y�9([��s`��������դ���L旟����2�I%��鉅���3�9����;�,l�𩒀~�*7��#\�w�j��c�?L�O�`+��� T9�(�H�OE{m~&���x�OB����w<���j���3���M��ޫ'��Mxڗ�ӑ�:=p*lI�@���뛨}v[�u�����qe^+��or���N�MF�.���o�+�ת�7�:�>s�c�<F�/IG6"+D�}^��od�����m� C'SM֙W3��tX[c������k`R���nu��M>�)`��9^`��c�b= ��:� B��q����4r���������:�>��wY��2����v���v�3��n��e��b(�%V;��pp,hR�4���טK�=]=M�yf�r�w+�k�냶�!�0�*3�
�/qԏ�gW�c��ǂ>֭OΆ�>+�=�J�>8��<�h�K8j�Q��2��sv)��/q2u
�@B�ESR��V6Z�Ŝc
�Ýop)ݧ��%U�����mPaU���*cr���yDԐ����
�D�h�1����E>�9�$��6X{B�T��f�>��6��I��x�I��|:����j�ǼYdV��˒�[��p.����"��i�ȋ�y�,�|tU� %�Λ��^��#8��X[�o�\�{�m��˳\��H�[����0͆�;Ir�;R�QG*��u�ڶM�i���ٜ���&���+�svV���D� �V��Ǚ���Έ8t:ޣnu�@�e��hq����+��Z:(ض(WU��P�\%ud޾&��R��X�}�&M=����d��h�v9�N��q�α��9NS��B�����������ΰ=R��P�\j�X���͖Gs)^�	�&u)�'�P����M�2�rZ�o��8����}4|�X8�_0k%�+mI@v�Y�f����b��`I[���u�ڲv�P\�L�������]�I��(s3=w�"U3����������:�(��U��<�z�F5�ΝN���c��+S8o����u�F7��K�X�A����΃F�\ݵڮ�LNY:�J6�f��<]�WY��I�`� d��y�x�T-t�<)�ۧt8>��l�gi5rsꖸX� oz�;�8�7� �T���s.9�����%�R�|�sa]�Ej9�A�o0y�)�9�7�.��Ѯ�F����tN>�`��=��i�e�
+�LT� ���c{8��XN����a����i
9�"��R��:a�Z�x�࣭�v�K�z�}v5��	 �1v�u�Ø��W{.�<�A1�b����m=��B��[3�:y����9�b�p����l��*x2�+��;�:)	��UٯN�Bd��!�Sjk��Xn<����}b�<ʬl
�$}�p.8�Vh�֚ͧ�kUؽ�rSf {:t��Hw��'��wV$�FK��N� mE[��!�jr���W�Z3݂���)��gB���O��+�`NŰ���HCN|���3�7Y��C�5[)ہT�j�L�{.nw<��1*RT�@�c.�<������Ϙђ= ��]�]֐�Wu��k@x�5W1}}K쭍���x������_}��
IM���耸>���n���rAd7�Q#�I���U	�N>��ux� 0L�1T�K�_S�+Rᵝ�^�U���L� ��������Q@
8��������^���T��׸�xv���(|(P��*��U�X*(�"[H�#Z�U����ň(��QQAm,QX�����V*�DER�Uc
ʢ ���QFV���-(�b��ckU�dE*��ʉd��ETd��
*������1b��#TA���%���#�(�X�EDAT�k`�����X�
0Q�(+"���J �(�EEU��Y+,T
�,EPZ�EF��ث��Db��ն���QQ*,����T(�DF(�H���)�5��(�j�Ub1���DQ���m!`�mDEe�D`�EB�֣mAD�����TEUV*ũF1b0Db�#+��UX�X��Im��(�Q�5���c���UX�JEF#,QV�Ͽ]�>���w�����nϴ*�f&��b�iiV,��ւt��s������OjL@��t��#�YZ��������f�7j����|����=���Oգ��2�����*�F�ȫ�c[��4��~s<��:l�D��eǧ�����c�g>�,��`{Ө�#׆V3�<�pr'pn
�	.�h�^z���Y��5����{�Hc��`S�s�S?\�E�~�5������K�-]���8�>�z���6����
��;%��Ϫ��ɭ,_�3�*|�G��.U�w��&g-'�|w�'�}��x�~�^G��p�������(�X)�/	��*�����j�{�&����O:�S;�g��2+�N�m��[�s�u�=`/z��%���s0}9��\�mVx�{��3$� =[��/%2��wp�r_�ǣ�/
��Je��xpN�[�t�p��w��ã����;� K��2<:)��7��wjģp��Ȭ�^������;��\M�imegw��*��<>V}O;,g�k�� 6h����]
��h���c��C�!W��ޝ�2���#'MH�r59��{�aRg7�4�_��<�{+�Xό�\LL7WJ��V.{񴢯7��]����v򈟮�ȫ�]Q_fð��Bu�N.���ϣ���f�W��# ���s)��cN>��U�n������k�e.�[R
�d+6��PZ�O�Z�����������@kUw�-[�m����aR'�ZcmN3�g:ݜ�K�5�ԦyMi�˻�4�oR)ȿG?[~Wi�7�(���Hw��0*��_s�t���|�>u�z�� 4s=ׇ�=�l���U~9��i���z�q�{2�~���_�@��*�������/�C���o�h�F�3܄����WyMx��v�6 ]�@���X�����<t�D�	ٛu��Dz�/ղk5SG�u�i�~�Q�~�f��@yW^�R�	���f�=zyd�qށ�J�ze�񸛖�fևq�^_n�jm)c��w�4��DW�n}^Z+�;�7:;�gKշp���7��^����v����;��:+M��	��+��31��!{Q�D��5|:}�{��{!c�
򣦽�V*��l��	�7Z;q;P��+�X��X��r_x�NW�������V���W�$g���9�Z;�t���'X9�Ix|��Ǩm���"�	���F򗏄#�Sr=L1�Y��P���Y_�������pu�����H{�n�J���&pj�x{G)B|l�L��fC�U}3��N̄ʞwq����<S+}��<Em���2�~3R�~DS�]J������\z���a>����n�ԛs�^���.t5yݴ*y�oㅍ.y8}g���-R)�>>��n>��eb�u'+)�sr��thU<�]1���,���ĥb��µ�`�G::�o�Ĝ1��1���!%����l�[&�c����ϣd	U|=U0'��\<�L�8��_���.w�9�vː��Lø?g�7��l�_JU}���G�z@�\U0&����J��wDx��̧�j�v�����K�o��@�L��������˿\{>jY��q.��)�H�%���y��b��a���37ӛ}H{t��o��;}h!��.�Wq��#+��=������fCu�"����S�wOzq�x<�Ǿ)Wa�Z/2\_<��u�H�?u ^����~�r.!�5
�r�{�<+��W^u�+/� r5���_A�S�G3���~~��/>�+��\x�� ���k.l�~��r�E�s��7'�,r7����g����wNB�zm?����ߍ�u�z�B�W�Mlu����z���}/(q�I�|T����\M�q��}}K�����φ�2l�*צ:����j���ͥ71BT�7 z���5�,�������n��ͽ����#޷^ڼ%�﷫{o˶�9dU����w�d�/Hu�:�7{V=��E}���I|t�����8���uO/4�ecX.Cz��SX"}]c1��j�t�X�ڕ��T�S$�uV����r�z�a���\A��'��S2�}ק0�0^�K�EX�i9W���r�(^��;�ӗ׷�D<e ��ԯ�)N��l�co�ȵ�����]����Uy��7��v���`����>Rr<��W��bE��8;��$��뿫������ wl,�xY��gя���i�S�9�������9��(��=�κ3�u�F���-�x��1�IGng����c2v�td�\�N�}9���~�Q~�e������BX��^���>T���s��p�R��C�gK��&w���લ~�m�����{����_�ɾ�����Φ����~�;��-����R7���ze�G�XQ�:�&Y�u�V!���j��g�r�ញ���ϸ�y��>Gr=��o�V�6��1�퉔j$����`E��C�R�gwjk���^����Q>���Ƕ���#����z2=�Z<�>]����u4�xl����u����G�
~�i�'�N�M���#]�F�{�=���>hς��W�~���2���'�Z����e�l����n�4*t���h��:��x�Ewνi�~��d�{�9�^���eĜ���J����{r.9�:/ 鹂ëU@3�n���n#���eA�Q93�|�4}GNP�ꑛR�>���Ԏ�s�@,��Z�����ky�ğr�w��~�v�7h��K�
U��y�y=`��+���2��w}�B��:��[8%��0��xd�p��M���\#W������^e��hs���\�- 5��Wwe�����J6=�IG�2��z#��i���A�H�g�pi��:��������a�kz�zu�#}��Lx���=�{�d�>%Q%�Wu�2�Lgez���A�B�3��״��yQ�9�܄�g|�Y:-�U��9�R����������DP���7������KS�aڝ��ݟq��7~-�_�?U�=�n�xo�h�-z�M�׶�ѪW����L��fl&n3v�כ^�q�-W�p�}�����9�px��pj�ɹ=s#�W���V/9�KѾ��8mzJ8K�챗���ʮ;��<�n3��K{=���}^����I��2q{2�fW%��A�M�~d0k��#��O�Ǿ�if��'´�jt;��73�7����k�泆<}�fu'4/�|uͷ�9��}j�P��:E��;��g˪��ɭ,k���{�ə>/�z9t��mvZ��{4��������^d����̮��!�����%V��HvO���n�_��ݶ�����B�g|�>����=N�k�S��μ�z�Ü�p�����wqEMCqU���tVGx���nv����@��~�l�7
����h���G��u����htw�7S�13�pd]BE��X��.�#N�oT��'�͸Eӫ=V�mJ|͕��V������[�Gr��f!���ˡ�ڷvz!Y.���bJq�5qY��t��D�鸚�1]���Je몇�?<���<*<S/��������ܜY�>���{^{3^�^�.ԁ*�΁�n(�4�x)��ՉF�+�`^��ʣ9���n���^���dS�:vϣ�W��xq[R��@l��9_��P\�M��w"Q
)���u5Q1^���������6
�i���]�=�⋓������n��t(�ⰻ���t��0�/-
�s�:^��n�:��ǵ�q��P�~�E����Dg� �Y���������Z���yX��+���1�v�N}3���<<��H�g�U����x� �<���(͍�	`��7Aυ\{N��ͱ�E�&@��	��N���wR5M�~���U~#�@�(.� �;;9���\��VZ���lX��Rx������͆:�3h�Q~��Q����mW���	��~�g���T�l�uv���`<>�ks#�2p��|T��2�x��M�6p>����v�F�JX�%��2�N~���Αy�}7w���j�*Pϼ�����Q�(���/N}'���ׇ�ͭ�����ݹ���~�w��[�e5�_Z�Hr�ܧfC�͌��/���A-��9.{��5�ô�sـ�����@��t9�p/���KTgux�;��Pgf	`ζ���|� �����e���jd���]}/9�vwPx�Kz�k6��3������7�A7�{{èO�����y�c��%�q�t������-�ڇ���3=�uYw���%H�ic8�� j�F�����H�{i�r<�Gw����F�5��	�=C*��jn����й��Y}3ϲ��秨��@����Y���o�k��K��
���%R%�]܃�ݢc�z�Ln�J�u�=c�$���g�B}���mQ��"6d&n"y���^�q����72��\�5}Ȯ..Ͼ�{�ƶ�+#dIU2����7޸w��)�u/�}/�c�'�L����쓛��ѕ��Zsݧѽ-��ǳ�t�3y�,��Q���;�L	���8Pl��مz:cW��=٧:A���yx����y�>G����9�>�r������n%ѣ�+��c2f��h�Vi�m�s'1���'ȶ}���P����1���}@m{�����p��P�Q,m���ޮ��s*Lx�^�����\P��f�|����zP.����j�m{ݝC�{}~�����0�3� �$3���}>��A-�F�����wq��~9��Tl�m�{�j�+De�ek�^W�Y�sZ{�7��]�믖��b݌>�:�:���O�b �Ej�,�q�.+�p)��[}ұ-V�p�|fk��q�W��J��R��nn%C��}xK��b&y���K�_��;�u6뺂��1GC:lCn	v�p���ù]< ?'�C%ʓ�Dχ#s�W֨��=�`?�Ц^�Mzn�>l��}���M(�r���>���)D{�d�gĳFa�F���IE��"�:���Z�ű�ד�Y�={���Bc=���_���%܁����&�d�t�CW��^G+3�<��v=�Ns]����y�\����VK	;���}�mX����;��$>9� ~���G�xO'mN^�3~�~�]��׸����@��[ TCw��ϗ��Rsʈ����P���V�q��T���n$�dvםGx�^��B�x���mV��R�T��C���s�Yf��<}zDʆ�?zV�CkU�����6�Z�:v�ef�e��څў�d�`g���ׯ��}�M���+���7�]윽5YK7c����;�G��Ew߻l�Y$n��8]R�:^���b�]&u��]�?yޯp�Dq�l������{��=�(�Qe���8]S~�����W��P:7+K���R�̅�>��dD������t?9�:��^F�ի��{l��϶&Q���T��-����}S��۹�g!e85�H�Ze�p61s7b8ܽ����m\Q:�u�C9Ҷ�di��<vk4��&>[��5u�A��c��)d�8��]�y�5YO�\Ψ����_.S��=���ٕ��Cr�5O9��WnoA8aٸ�d��swaNM�p���'c߽�ژ~���XϏ?^���l��*���] ũ����<%D�>ST/VhF�b�@�zi�&)z�7�x�ȍw�� �M���'�vDo�����U8��W�
�7-sͭ����,�y���>20�H�%��ϟ<�f���u�H��=
�8(ݬ�֯Y�h��ty���x�Ihr`0��P�.|�`,-9����o�gD�5bS�����z���;^����|�w�G=�]���"�˒����*�&&�Q�tO�vC���v�3��琭����xzXۅ���[2�����I�{ۄ
s�Q5_ja�-�te�[�=���l��n�ѽs�=���m�ud�o�^(���s��=tA��|�c0B�����;ޞarV_�n�6�L<�������7~-��xZ�r#�@�˻�V��-҉����5Z,x[`0Vd��7������A�*/n�Ǟe�b�Qeۍ������i����^��>������p�r��\�M��~���+��v_����&"=���ډ�w�b�G��X�5'^U��ԕ�S��0O+�/��+h.�I��}7M[�Jif�� q�${��,�R��Ծ�@l̵��`N��q�/�����:�������WO8����bw7h;w������Ψ�����Z�K���V�wO�e0��_��x��~������uD��8u�n'҆�N�eV�y>��U��&�9�LM�+̟��������x�<x�=��7�Wp�l��+����?r��}h&�u�\�	d�Ϳy��ۻ|X�9���:}�C^�"5׼H�����l<�{ט�o���#��~=壡���MΧ��|�誆�}�u�*�����1�ׯ�sT��r=��\*�CG��2��]sw�{(`��)�!��b&��Mw��FJ
����K���=>�\-�E]��Z�=�x�M'�X�!aM�p�zr��c�%T�;�tX�����)�c�O���#G��%��T����#*�g�|wNx�5>�~�e@��= r��]
.Z&��c��}�"�QCnguS���S�ox���
����AO2��4���ì>�Ib�Ί�:;�-׫��oՎ��	�-�y/W�8�<�ia{�b�*ۻ^,?t�����Ց��K4���8��A2yg�Ł�w���AW<L?�6��%#���wF��Paj5�p�w��_��0��! BI��!$�XB@���$��! BI�I	O��$I?�B@����	O��$I?ܐ�!$����	'!	KH�y!	O�H�I$'�H�HB@����$��! BI�Є�	'���	'�����)����m����),����������01o�{��DB���\ڠ�*E;2��a����T���]��y ���TJ5m���b�����[4��Jx;5�2I��Z�@��Zm�f�V��(:%�{�(���$E��
�xo^��bرMB��e�kFEf�YT�-)�	UEJ�I�f��]�Cj3j`�m�LPU:�6ҵ�׽     �4����M�A���	�4��$�U�4    �`&F F&&	�bi��J����	�i��&� �S�R��H� h�     $AH4h�'�d��140��Tz<���3>��I��'���w�͊*$$%�I$�����	q����?��A��q�i�V�@�C�� H:hR�!�6"��@vb H���s���O���_o��@I�Zđ7
;�j��5�����fT( c}n�������
����g_+p���'�̓�)��*��
 �/lÁ��0ښ�]�B��6�T̲�n�f�lT)ed��o�h��U�5ŕ�E,��K~Z0��&�Z����i�0h �DY	��L�ji��je3G��V.�"+c�2�q�9o0���=�x��ѫ�An�MnŐ	�A1^Jq�F��9��qŎ���ۻ��&ԥ�X�ƣQ-m�2��ܿ�խb��@��VV���1�����|���(��P"�R�v�ђ���Bi�O�X�0��(���&�ܫ�ֈ0k��qb%b�Orc�Vɠnɺ�B���1��o
��J�^�2�H��0i������k�/U��+�PZou<�SfAї(�f�Pt�!"a�,I�j�[��*�w�)A��iMKg�J.�
��yMDf=��:� k4e=9�+RjR�=9�F��x��������Â���m7!�Ζ*���V����kYNG�P��[@�j �0��%�Mi�l�ءBբ70٢U^n8s0n�M�c��i��[7�xHZ�r��X�;��j��aB��9{�OKՈ��թ�KuG����:����҉��$�/qH-X����9��e*AȰ�(3�n�F��-qQܷz�]4U�3j�x.i�`@��5�Q��! �y>WYlI��'F�"w �F��	fkRص���4>�c4ޥ�D�\w(���a�����0����P)��\;M��z���Tͪ�I(� 8�潡�u�d��=����,�9S���-��1�+sb5j�{jDS4��#@r�agl�V�G@��k)Sx�ޛ;�]�Т8�xr9��G1,$AZ�5нT�YzδN��*ʅ�s-�4v*B���-S\.�[��:�ިI,�P�m�r�o&��K�����<��jm�J��K%�A���F�SXb��gagZo7M)�KtT��
OiM��Ct������
4��w�j�$� :&\���b(�q�dJ�d��LL��[�z���K����y�������u�����ZM��EfI�]KzƣRv\��kr�N|�B׬;�w8��񪨝��C�qtO�����?F����:oym��A��BK;�;���Ƴ/_�J��ݙ�XPWc�D���K�]ٽ�o�Ł�ݼ��8�WV -4_oXQ�p��MQ}[�B��j�wk�QL��&�ƇO�NX�gl����(�ݕ��I٤�R��F.qE{]��ڭ�7Y�)���#)O�_R���ge������`*K�i�]�^W�Vΐ�or�p��+�8��H'ٕ��|�YY�4��<][���wB�K�U��>e��������f��V��R��Y(����[�Ҷ�(�A��m�|�a�;�������v����sk���:	���#����zv^�~˼��T���t·m���=��ZU��Dd��D5O�qD��e��	 ��TC���C�T�'t//{�:�l՘#�y��Uk�7���2�#�7���6��8ۼgr�s���R(uh]ǟ�Vjr�.�0/���y�W*[��H����f�s�Ήπ�7$��̺Ԟ s1!z%������+&�L�c&�pS�{��E�(��gcXա��>�չr���܋XqӘ`�|
IM��79����+zu��	�����A�,����λ�S��H=�y�
��鋑u���V�y�j���XWR�
;]Yh�&���1���i�W���Gbe�=dr��[�.ﭱ�v��>�=rK��.@\�����I��:�.(�Gd���I���b��Y������[���{$�ı��#�lN���k�EYȄ%��
�/B�&�O8^��y�����R�Ahdm"�3�ׂ�+�L�KdUp,u�|Ʉe��v�o*Ǌ�{����Ї�H;�![w��zJ�Mr*R]a��b�v��w���������b]��o����b:�˚��A�F���Z���
��XG'��x����MxXX�q�]�Ҋ�A���
�ņ���TH^��Cw���Zi-�n�eX�+���Ȣ@�+�o/Xf�N�j�� �F��A��o1*^�Ǵp@�}�;��%�6��ӭٳ�e�$�H%�`�:��C$�ն(e�t�x�s��Y��l��M�έ���P��y���!z{2��}��1��mwWv�M�e��X��9K찵�9�;ZK4��K�f	�[Q�5���;�v3�m��"�����TM�ާY��}�ã���3�t��$���f�wi$ �� =����	 ����\�/�4cZ��e2�̣jQkXo�f�����Mq�:��v�*V���J�\z����ZȮ�Ѵ�+�ۅg*p�(V��n�/4�.ے�v��yu��Ns�VS��]ƯQUp��]���0�m�ײ Jv��/6V�m��#���X�'e�]��(��:������;^�Q�WG/9�k����L-\�NU��|�>ֳ�auxn�Z;m���7ݙ�\ꀟ��}@P�͔�`�:�w%@ܼ�v����ш���-�{f�#�)�7V���Yٽ���N鑙��Y�]�c�;�m�J�h�{�q����d�6J�*�[�[�W`g(9��#r��F��+\�ْ>�.d�����R��ϹQŋ���u�h��8�5�M���ܳɝm;��m�L�^�o�����|�-��j�Ы����ͷ:��k��U��\g7��u/��㖎*%͢:s�}x�.�][��݈�{#�p5�4�u^�@s�[�p1��lp�N��I��Zx胮<C9�2<��Z.X���*��4+-
ǿc-m
�v��ܩX\�9�I:k�'[t��:�){y%��ԃ���(vܨ�I(I�,X��+�2-���9Ȅ��Z�.�����]XWr�!sos�|�"6�oJF���AV��	&ȡ����:�Q��={�|;�w�YJ��Θi��`^j��i���hTL7l�sB*�_	m���Z�ޘw1ԍ�8B�����cp>Z��N��WEÖ�u�7�N�+n���Z5�N�m+�q>�#���U��}m�{�n���w�f'���n�p�i2�slfξT��h�i`ia"rt5I��q1��[_^,)�
�j���R���<����iӣ��h��T�t�/6��y�E�c"-�7�Xkyj/��z�e��m�L���v��e���;pH�[�Q���ܱ�Q�u�`�C@X�J٪�K�1�:9�1Em
�ټ�n�XB�ο�2�wu={ף�v�k��Lv���j4�p��k2�Ω��\��:�oܔu���

�V�Y�Hr��p9���uBUk�k��/t�����m�ܓvs!��4�������;�"l�\��{f£����]d� ��@������f�E*�z�Y�]�$	 `�����A)��Xo�p������Ẇ�ڭx��U�v1���3����f1۸���2%@,N��z�kOL�4V[)S�ٻ*��vc�;zjV���gp>���=i�^u�PWW�gPK�K��|��7���i���ؙ���]CSTmBq�k5��o\mY,���s��fZ��{2*���Y�痒�<eԴ��A0�g���	���[f��:�8�P���k`��J�3	V��4�v����X���՝W���U�t��A&"��˗�s5fK{���b�`��u���Se�_�֯cM�t�g���Kb�Z1���v��/z��y@�5˃��t�fz;f��t؂�]��g#n��!��d����^�*Դz�]�]0��Z��%��އi9�k7
&� z���r���L��:-�b����ڗd�[�R��{�s�h�י^��@um��g����BQ��۬�3ѿMC}�4���^r������:�5Ya=O�p��/W��ײ�<^�{��h��V�Xt�{��A���l!rU<`s��9܏=����/!C�}y�@��%vjy��}#O��k+q������AT��Y��e���^�5�wZ��x�j�Ntw�Q)�8��4�{�]��n��j��sY0��Q��<^#�����_d�zI�giݩ&<Ʉ1�??_S��;��y��n��Rz���9�&-&��`o�gz�:�	�w��]�v�j�9-�aם��iS9[V�Y�7��tn�^�A~��^���0S�����T�ܑ$�x���L�:�j����j;@缟���ͧ��z��#3(��3�^'�C±��J=�W-tutnO :�xBN�n�S��W��T���YΗ�ϊ�M�9���k��Cts���r��N��ab�m��c�%�]�y��#]f�2�e��k#N��{�^��_��^VS�@�/?$��*q�~s�����\��l\gKT���mQ��C��g�ـo�Y�ӣ��~w����*�T�۪q�^����㺺��V������EJ٢��)��'���.�K�Kʸ|,��]�s*���9��K��?N�u���ڞ�g*��L��E���*c()Q5�r�Jȇ���
!�;y������q���{�̝ټ���v3�G�c�>�"�F��+���kc)��)���Ww8Sj��_sr�4�WL��8������+!�T7�̙�V�Z|n���4�1�&a(E���m��dd:2 �V�v��Ӧ�w�5M\EE�K�X>j,9x�ˆ� ݀R�e%�kJ��H:6BO�et��]�c̰32�1NfA*�,�C�ԒbI7S1�HU)�^XҶ@��#S0\��,\9j33k��(P�¼H

��(��+,��f�H�]Š^7V�%A�Q��LJ�J��=T���bp��AL�	rBR����b��{�^���F�w�C�W��c�	�1�9NG\��׃C�S��[�Ơ�PJ(߁^m��?�D,��M���CA�[�S�s������v�r�ds��8vfne{������]�5�#�_��f��C�m�:�3�.9��^%�q�z�z>~zA4��|�oӣ���"�ԺbJ�J��a?����y{��j��'j(O}V�I��5.m�$=ݤU�G7+6��<�.���=y�/UG��KEk����[LvOk��J�yeJA�u��^x�e��틜����,+��t���z�xF�>F�H�>Ӟ���J��e:Xfy����k.f�3ɽr�B�T��E���HM�H���V�l2�:idhH�^3i#�D$6��K-1\$e�m���o\�oU|��c6�{���VU#9��$s��`�� -��8��ާ��FZ���iC��Xk�DP�����Z�4�i�l����D��l�i�[i"jD���ا��M�.��A�!i�i"jE1"Z1�F.��$[���� i���)i#M$k���� �B8Җ$t�A,-�D4��$s��hK-M$i���$��ؑ�
b%�c<���C�!#M �`�T�cEoX"o�׵��iT%󒽲tMՔ�-�ͳ~�k=��FH�}Q�����W�Q��������\�\��RY�m�����x6��;�z-����D%�<掻J��X�#Jl��)�Cʅel;���N:����1�ø���vME׍gg�{����ˤ��w��z:�8�c���T�~��Kf<�gY��Ș��r�,�������l&�\wR�m�w��Szo���4���,����OB����cn�㬀^�oi���R$b�0#5�4ʗݭ�yge���"-31óϻ�r}{��R����Oٯ)=����Ix`h/H�b�$�NA��dZKţ`�ޭ��L��c���Bn]k-��I�N�������gTM�ql�}Ի�2�'�߹{WHa�9b�^��J������^
�?����sr\����nZ�����dJכ�e4_b8����D�Wl��s���������u���Fd��qU����uo��_?h:+h�%�n�����P�������S$��_�e��>�7r��A�����EZMP�^G@I��eYT[$K�R_X���[Ǝ�$6��j Պw���ަP��6����F�`���wPF U��༅Fca��iBB�wV�� ��n�f�䣦��M�e�ɄZ�����b�h�����O.�E /� 0bn�n즪t�#���乐/W����P"����lvĶ�v��I'�yW��UFe�#bD1�*���ݩ2��M�2VJC$�Y��L�l��ꪳ����U^�����W��W�|5k5Jݻݳ�=p39j���������f�����#�<����
��~{?2}�V�ɪ�;Gv�o�B����'i��Uf��NWzA��p��ER�E�d�K^�i,�k$H����1.��*3���b��7��|�>늭o�������P=�X��`�o��_������E�+�������*Xo�՟`�c�<SZ{�,���7�Pk҅����i5�sr&��j]�cC�<�G���y���K
R(O��r�_V��� |��zc��C�Za^dl<��#��TW��_q��o/5�i�[��$V,o�C0�-�U������<�m���r�Cڻ&1.*�[�ް��3}3�M���f%����X�S����Q��{ٰtZ(������V�r�����[��];'�e��pɳU���G5��f��q����T._�]p^��O%|C�w
�||[~�ϑ ��8�j^��\[�{�c(�{���¨	w�.jY\jcU��+p��.��r��Z��PG�[3�,J4�;^,�[���`����\�L&��T^V��45�(����z.z_}T�ᾍ~`�b�2זe1+.���,]�����r�[��/ѩHf��Q�^p�G�6/2d[�y(�t@^	"���P)�{�t}��R\����I�iJ���Nbĥ\�*���L����ӻ�v掌�Wf���ӻM��H�/�Z ��c�]�^��\w���}�Jկ{���u�dLy\�Gr�����ff������,5t ��/�_��{�{z29]�2(�o*yA�8Yu0�~�8 �o$���{�tn0�5�WY����s�;{f�DE����I�>�h�[�����V��*�ű���G�mb'c,یþ��~�d�u�)yW��s����[`�fg����L��d'�Iv6�`.Y��>��U�ޖ�ʵ���fS2��Q�mP�����WJT�5�n�wyZXw��c[p<�"��]��*��E7L�t�T�4�0�i�w�3]O�I��.����5w�I�-G8Ƭ��u�sti�r���V��^��S��e������s����U#ir��1W�̂���4<�U�	���!P�@/�b�y����fc���2'��D
*�Z�c�� ��+���E'g*29Ԑ�@� E"���,�E��m��J�=OB3L�5�-��1lŪ	s����Բ,�<�RB���mi�Bʖ֓h,�Nt����Q�hDD;��׻To98R[+o>����_R'��V@%x�]� #W��;m� 9��}s(6<լ�.��W�*���ҫ{ؽ�H�a`�gH@w�W�V�7P�;钶$U&��^��?N5ǻ
,'N�ݍE��0��+ޓ�qוS绸�a)������_�y?]�_�N	a'��f�ʙ��>FrD����x\�;(� hA\�=��Bk����� ���ǝ�͓QNp���0ɓ^�pھ��^��ݡ�t��s�7d��
�v\�ߴ��A����Mӓ��:��r�Ӝ6�O'�n�sn�m	^�/3a�/����Y[gkb4����Q���{�
��c[��A=��!��4=��]�v{4�v�H���~�����U�3D䐻0��~�[�R��5k| fs�^k�B;#.��Ui6=1J�b���q�:��L�k6?lS,�^�{5һ��	9�y�̸u7�8Ŝ��]�k+.�|~��DJ�?�N�����`;���t���r�JS��`A;� 0��Ϣ~<JE�*RH L������u���V�īz硰,k�VE�D�o��~b�N_�m^	fnT�H}��������g��30�S�B�X&6�o�Ӌ((7o=�'w\n�ؤL��o��9,�gI�w�=,�-���@�ayK;��~����No�,vdS���0��F/S�[��{g�����lT����y8$��g�Ϙ̻�̻�=(���0��b`s2�p��(j�jFN�/w/-���L!��4T@�-ˆ6�2�n��յ�K�������������o"z0�Χ��Z�-7���fȰ��6ìA]@[C�}Pڡ�������[f�"�X�n\4��sS��7���0*r�k��ږKR�nxe�h�p�P��6іj������;ia�cgP�=�ы���[�M�����4j2����8�b7�L��:���ﺦ�řx��[{����G��5��T3�Ӷvce�bmC\���`�C
�[�A�cZ�(t���5�a���zĬ5/OMe�#Yl�Ds<��r�5\h�rjV���%l8҆���7ʴL@y��.0�gDR�e2ܵ,�U�-��#S[b�[/R5X�'S	[B�kDHQ��t(;x�T�<�f�,s���A�B��tq��FQ����m� �'M�z��U�}�4T�z���N��K��>�Wq���C1�u�E�K9�2�^S��:&�%O̴�x����a���,R��(��+�Y��R�TOS�H�������WS���̥x�'at땜��M2��[���0%����:����qM�T
��ɛ3���K��sO1t���]�o��5�N��8'qi"K�5d���r����F=�G&z�BkD��h�Rv��#�V����#t:3Zl䴚ʙ�T�$��h�(�F"�FY%EY�W�i�L�"��S�&�fI�&\ґ{��g�o$�J*w>30fŬ1��\���T+d��CC�.u�u�f���Ƕ������sư;�d�:���k���:ěj�b4�;�`S!� §\5��;�mv�	�nL홹E���8f7|�o�ޕDء�O�fX�0�l��B�n�9�]�:�	[���vau�jM-ݏ��0%�\q���KGf�S��a��m��Z���j��[f�%���"w�Q��[E2Z
p�ǚ�氌2����n3�Yj=�;S��q.�*W:G]�a����)��'s9��6�{u�\�w�)�5Yd�O��7��)alQ����: �	����>;�u=xgf��qc}���TP��fp��^*y���X��:x.8���A�KM�D5U�ɗM[Y������f��l8�fYMY�:�4�j�����f�㺺ݖ2�SR�\4�6�LՖ��hl�Ƹ�/5L#,�¦N�q��^3��5��1L|�S>�+§s�4����{jmfn�[u����a�����Dø5,.�'Ch�-��>���e��q��T�O�m���8���Nٗ���튚���H^�Zt�̴�K9��Х��P��0ͳ8�:�R!�2Z�)�He���噘!��d�մm���gP���BR� y8��N��^$���7��L���b>`����`z�l�ƶ�˵�X��6SP�9p���z����j����e�t��tіglY�Q���e��ٶe�Zb�������r�qk,���w���^��[M�ѬV�݉�����-��wP�(P�)i�Z~�=zK��P
�2�կV�!�+w�0 i~`<���s�(0N��:�aƲ�5L�=���aLA#a�y. m6*fY.w�Y�aK�ь�L
r�yz�8Գ-n���skR[X�a��al�Q��҆�n�7Z4Lv�xb���5٩���)��;1��'�f�,����vЭ�e*�Tt�l׺}g|v�s�om*�S��3��4�E���.coL�m�Z�e�ma�����Ι��Æ���q���>2�4�l1[��mᙨ0�i��0�gT�pe��K���z�)���S)��,�)٘GƬt��0����W��W�TU}[�{�m��Όox�BH��-��}1��&�HS�i��]��20��)�qMi�PSV�N5�;�3<�m)j7��k��С�mC'0�p��*v���<5�)kM(eL�֢�:���[�6���2֙fh����|{f�[s�R��s�oO��\�Nƛ���y�{B�4!�I%J�$�R���`�r�yۜK�S�I�i�k3�%�Mt�5�S�)��#W	F�H�%��;�3��t̴K�2�d5l��T��yfh��amCP�C�8$obP���"%l�ὢ�t�z�EM ��+��^n��̧^Iak�%�Qŕex36��X���k��^�H2��#�����J�w���/}vP��h!w�䭍<���؇��)�:���#��}f�Z=���e��/�RA��mjU���v���t�n����-���ZM���ʆ��c)�C��Eؾ_���4��.V#[�k6�r@<Ķ`I���[�+��"�2�ԓ�(��Z����*��n@�%���͚WN�8%^
Uu�\9��Sᣅޒ!A�=V�ZS���3A'CӁ����ES�.�p|'8���n�VŇT��(�9kwr�y��#,e�%�u�H���|��06����e����j�dJԏW>%��m��ݹ'X�4�u�ёMX�ЛP��Uv3����y��r��M�V$��4��fa��P��A �	�������a��N$���0����9��EG���/����Q^�sW���/�;z�SV�*�
Cě�5Y�Z�t5y˚x;·h;�z��iؙ��s�y���k�Ç��Z��UR���?z�����=�"9��� +��!*�B�{}�y{)�/T�����&�2n�A�b5��S3�-�<���#/fo+�,�����5h���ЌFݜ$��N�Zd�Vxg��+����2"��]�@��?=ۿfx��1#�/}���3�8�F�e�f��l����"���~6X�j�%�[{LN��/E�!����`<�9t_��:�ŜZH�m��X��v�)�[�:��3(ԙ�:�:������5������}�cU�yi��
ю}` ��C��ߧf{��+M���s��z��vY^���kxy��}����� �#���e��=���'�;_��I��W:�2�� �x�(�#��y�Z��FoU�K��i����3:�E
�ؓ�3+G�;T�9S�v�|ޓ郩��9��BS���G���̎��$-j�)y?]L8�ŧ�z��kX��>�&�yٚ�v�u�c<�M�3?U}@����?J�@������d	o�.�i���˫�g�O.�T�s*{�����{׻��i::~���q�::/�r.��)c����-�WD�TJ����Uؘ����&TC'F�6$6y�ct��c�y�Ǫ��k���>�"�{���b٫Ӕ�+:�W4�d�������$�Jf�|�͚����ޝ�q����yyՁj�`�W�xX�y����Z1+���g�U�]�/zy�G�پ�W���2����=��/�Y�c�=;��ki� c߽S}�����\b���r���B�c�-)�.��P����C� g�o(|�`ʀw�ɯ�=��;�/zG�dG^����
���]`5~	Ls���ܦ[r�V;�\GL:}����m ��j�]#�>�Y|;;��d���}��Ȟ���)9^�P��w(P���(·up��=Np�Me<�]S���z��m�M�u�kw�Uȯ�+ޒh�%�FB��kF� �a#�C.\NX�[�Q�Y+����7I�+�+(^Js>W�,a�y�bM��	�,��,2����E�n�b)B��0c��S�`�P`��2�s$|MR�TA4@	�U�BB��&5m�һ&��x��t���G�y#;o<][�g0�{Eŭ��f]��k�����f5�)��+�v<&r�}&vn�o��Mv;��I��U�������xNю��/s¹ ��c�)��^7�Џ!��X�ς�!�ܿB;�'�񉹇z��t9�G#��u̚v��@�x=��͹|�m���ݔ^�l��t9��е�#Q���+Ɖ��`J��ho�V�ˇ���X�EW���s�{�\dY��u�q�j&��F�30m���?�Oe�ԇQ�������m�b����^�m�bcޝ\�����@��z3���b�H�n�����R?#O�F�N:�V�y�̅�*qMi��O�ٯ����,r��=7Z�L@Ҳ1̹�����k<շZy�&�7d8���Y����o.�++��f��,R��4_��졀ynN��^���o-��UUUM�K}~��O��6�3o����e����>ǵܸU��ޔ�y��t�B�T$4��6�{��S٧"�޵Tl�N��Y�P��	nx`��ʺ���
�fV}a�:�Ѡd�?%mǜ]��*,����$7¬�w'裕l$�׮�S3;Ο:�&���/3 �涁y���9���ݕ���>z|^���M��h�WDz����-\��K|�/K�~kU'��,��yuHQ��Ocδ�bݬ�{=�~�K����N�֮�¢�ZV�j��0�9�Q�g��/|�nٰ�^A�KZ����1jŗ�����LsZ���CK��k��y`�]��=r_���v	�����D�z����B��w���%Q�#%'�[�Nw���j��u�轧j�5�_��ئ�GǶ��^�2�|�4J�o��<,�L�#��o�"}z���w�ګ�;�cf?don�E;�q#�L�Msck�X��.�9xd�Da9~�/��{�t�i��"װMaR�nv"���T��\U���3rU�D+ޗ+��/�
ܻİ|m��Z�#�VUd�^�jꮘ��f��Z쮭fَ���۰���V[k[�����#�(Ϸ����<��0o��2­G�K�o+S��MYW��O
nԷ[J�N-_oo$[Yy(ታ@<�"b�Ӂ����7.[�E�L���X��τu�i;$У�2B��1yr�H�ڂ!��DB�Lh�Q�v��
R�
�em�V�1 �#R�2���6*C���U��h�X{y�L�䷗�N<����Q#��i��GM�x�25�4��"�w�"]����?�d��wnoP�;�J[�<��~C C�Ȫ��z��ئ�.tr�-nL�X���}ˡ���l{�
ڸ_�v��k��)泫,�LAW墯F��M�wRe���W��س1����T����@Z'3{l&o���#0���g(&4+�w#�i���ԇ�*�T��=D�F�!z�����.������/�A���T�W�M�e�jx�O���ס�x��h�����#$�L�S�W����:�- b�ۢ�����u'��0py(鷼�w$	%�/��)�wsK�m>2�lWc��D+\�D{��Ź��g�Ү�0���O�������Ni�އMB,�@/�k�e[u����x��!F����7��k��S�#O��Eqc�;�fP���m�������[�����������+��ًVsC¦2�[������� {�o���}^�b�6�i��>��s��ua=�{.���=W!~��V��>ׁ��vZ�=�������M�C/M��Ɏ��@J�>
�3X��jM�:jln������u�\aɾ�D{�Bk���F��݃a.�b����)�j�.]�L����6k����r��WԜh��Ww��C�^d��cX�Y`gJ�8F(k��)ׇ��{f��_��Ț&'7���^�޲���ǹ�\p� ���+�Rr�Y6�K+���;��c[N�n	������o^O�����q�5�b������ڬts{D�$�NһV �|~�3a��B�Y-ͷ��v�5����k��M��$�{�>֑׻y-�l�t�q~�f^�1=�]�n+��~b��/we�C@S��ۥ�j���Xƛ/%���'��X>�B���R�zfU�KSi�s��)�{]�k�x�U�V�kɣ�7�R�¯ּ_2�㾡�ĵV���YAfTt��A D�߹i$�z�'�Ӯc43U�B�v0�w`)$�"���u�u>1�C.�4Or�c��h��(0SU�J�9�ڒ����|��!�1Ю��A7/1��Ȼ��
<ˮ.��;�%���xG:L:���J�x���6R8>� ��Nȋ8�+�n���(ا*K��'X���[��\��f`)���4��*8�t�ެv�Ѣ��:�/.�J�rV,�]���0V����y=��ɹs��׏6���l[E2B�#;ry^�Y]N�t�c'���TTu.��ȕkP��|o/Ow����{͞����+���W�Jw;"`���󤭮&y�5msF
`�h["yZ�\a�# ���/Q�ac�Q���Ͳl9�#�=�e��׼�P�T1JmT�1�>`I�Tm9|�o{=~t3��5����{ʛ��eN�yYL��njwY�v�o[^�S�D}�7j�O]<@�y-8����w���G�F��^�b�j��y��1H��7�u���u��*7%פ�)$wo��~w�==x�u%0��U����T��+�$Gk���#-c:���d�Zw�c#�Y9E`2{���_(��s�Cն,z��G@c��e��P�����	�o�Xi�o�Xx�\�;�a����]qf+�/g�MMΩY�@9[D�
�9W �$e�7�"$�̉e7�4���=v�0W�� ���0}o8ʹņLGЬ���g:�*sr���U��/��s�G�tI�2�|BkV�G�S�H{2���VIǬ7��G��d���=��qp�:�N�����������XG�>b�j5���{<�<w��J��y��D�a�6��kv�>��D�ס�&JtJO<��d��4�㙅�4?1~����^!j �ؠ��4y�E��d�8�Ї����!�s�=z=�*�vNd��.h#�0�	��*��쮲1'\�(0a��3�]}�ӱ���_q]��l�x��"߷�g?|�����~��W˽4��8[���+��"��@-ay�h��4�P^�ڳ�j���A�`W�x�U�_u��3j�n�{Hg��}�P�程�W����M\nO:I�EP3��3�]b���ܩ�5�i��M�Q���}r��;�Cy���~�{dv��Q��;Y���	����b*�3�P���b��@y?�fx�l9�{iA*��'�E����pC���ʌ;�ѻ�#l۱�P�^����|�CR�T7F�x^>���P�~꺷�`I���2���اp(REڈVp�-���⨡��n�U0M���Q:��cٽ��:�N�|I���^<6�����t҇��weX�6�\�,H:%�"���!ܭ�$��8�uve\GK���cr�\��.�<����=�5��rΧ�߀N��̔t���^(r�T��Av^�7�Y�\��%q��ݴy�\�f���FQ=G3���������8������nE�K�QJ"L�9u�,��%�2H)�&�HE2��h�&��x�A$�����Fasr�!꺪����z{zz�>�쾷yهC+��o_����TV��*��b�����~�O�w��ŏbp1�N��W�1eX�:��6� �w��*��g���DJ]}�>��9�U�6NW,��,��
�נWz��R8M{&3懙ƶ��tI&����",����vk�~I�_m���;<���K33)f��}8���q�v����y�5��д���H�62��g�]|�-f�,r�r�O��qV��T�U�cG=��7^?e�iR��{&_>~�okn�u��H������z WL�Q��g�}&�1�8:�g�K�&�2��B�'���ȫU۱^񷱇V��@r��4�h�����ޖ���jT��#&�Z�F���E%Wp���]�r:lȊ''�L 7�ʭ�۠	���Z�B�ܶ��$bS��F�si�W��o=��IT�������`����ݗ��]�o:1~Y�6d��<�\c�b<�S'�U�������%+O�+���ӈU��{�}��k�[��L�5Q����+��z�;�
֥��Q�R�&N�/-��b�:ĎK�|��)��c�gM�p��$O5t�2��\K���cp8򱤑���Ku�n�ʅY�mn��ҡ�~��S��h�����(&�ye[G��ç�芅������.5Kô{ܡݘ�,����y�>or�]o�P��l�u�*K�^�z04�-�����N��Vݸ��<M��B��=��T<�]�ڣ�=�v5�<Yvx�'}� ���b���δڽV��i��E�K[2�D����|�*[��cH�0w����{|eseW*�}.�*ֶ�-G9��(mY�t��8t�Nx�c}�3!1z��<��n��>v(�WrnQ���S��j��y�C�)�y��W{�C�3��z<��\���J�V6��z�:������|����ˉ�UW��@wpf>��w��D-�!$*�����!5B��mVϾ�����M ��N�Jɚ��X���óA8]���,�J9��%��$������o��-�~h�<��u���]����I��Z�g�c 3��JLo���I�!�Y�����ގ~'�}���O� 0ȽhBA�A�A���	�BR{����pa�IL���d״���=_��-z��� �����~�|�����4�V)��
A�R0��(1���"������%¨"=��_���a����wW�W�	����_��`�$���V�<(���	$	 ��:	m:m��ؠ�/�2҉���fCȴwt�$���a��3x��<������@~>�ZEw�aЊ������_�
������c�A��@A~�����z;��G��pw��`�?[;���� �d|=^��j���<R�?z�.���=�|}�ϑ����$�$��0i����k��N֍iZԍ��9�|F�P.� �Ai�� !$�����_�G�p����>H|֌��}����BH0;�Ƙ��J��@?�h]�"@�@ƕ�+21/#�0*��O8����3�yZ�%1����o%�Z���� ��o��>;�G�IH|�`�bz�w����?wa~ގx����A����D�=�� �P��zX�G�z����^�Gڏ�A����˱�����I I��/�<_���$��_�C��HA	},1�OJO��G�ߏG�/��w���'p|~�#��`JQ��A�%)~���1_�^��[Ǽ�}�ɿ���MI���}���i$	 �z�2�~�ϟ��G��#C>9ߵ����]�ϫ��>�X����b���b_13��5�|���?Wr��z��z���
���`XWi�BZ��%{�l�;�6����u������H�
��@