BZh91AY&SY��F��S_�`p���"� ����bA^�     =��U�e!���l�P�45�l��TIRKUB��6i5�6�+4����&�-V�U���(4ka� ج6�Y�k)P�U�Q��aB)�Yh�E���[V�BUl��m�[4ٱ��Ujڬ���m���H�ke���Z�V�lm�E4Q���T
i��j�B�d��yB�=�IQ,f�ʹ�V$4kZƉkJ�+MUiѦ��Q�K1�e�5P�(��Қ4��0�V�MaVE�j�cMZ3Y%*Ց�{��=%��٪�  ��XR��5݊6֭����[@[S[���mG]����[m��vk�w�Z��v��uķ�m�M�iv�׽B������ҽ}���V�P��e�Z�i�j��[f<  �_g��R�[�qݺUR���ި�T�G<;��JW<���AUGz�ǥ!JD�����TR�H{�}��Q*�����}*T_f���۽�%�en�ɩ�Ef�l¶�"[lkj  ɾ��)RR���x���i��{�N�U*Sx��RT�R_=������)�}���Q*T��{޻i��h_:��zJ��U>������OZ�7||��BJE��km[Z٥h���
jْ�� w]�|�}��+h9�ojR�(=��|���"J�.�y����_l��
���a�}�ﳪ��z����RE{jY�{�J�QW�n=ǧm"tҼ�jw�)K�J8�U=�2�b�M�̍�  fG���j�U�^�)T��Wq�x�3m���=�JB�*��J�R��7*�Ґ���Tz��5{�;��$�+�z׼�$�E�N�IC����+�+F4�Mi�T�UE�S�  w_}��)��G�*U(�=�{ґ+��{��E*H��^��m�^�V��y�
J�.�����U=4�z��UKٔ�oz=�ZjJ%��=�US����K*I���3U,p  wc�ҕ"[���<�E]�^�Τ�4�M��޻R�;ޭǔ*���^��J���ǻ=�L���<��z5�������� �؆����a��+M�Y�   �>*���z.��*��՗�� �w%��E�\J��8QB%�{�P��1�@�3/s�PPy�\<J��zA�f�ٖ�i1+MUE��  }�����V��^��A@gW�=H��{oyѫX/r^{��^<�'� 3�n�%y޼ =Q�ymހ�Z^��:���=iY�&X�M35m1kRض�  &�}]���z+M^y�y�E*����m�������x��ν��^�Ǻ�
����R�h!在 �    4  50T�T`    O�1JQR�@`� #OɈJUD4 2 h4�A�JJUF 0   !�J��I��  4  !) j�LF�=(���=L���~oď~_�[�C����Z3~kh��K�ws���%{�sugϻ篝x��U }s��1AW�(���r�����_�?.�=?����?�T U����� ����T�t( ���?��x?6P��!��?�/�����=�'�e�	�;`N��A�:`�;a��D�;`OL��(��`���{eN�S�A�}��l
vȽ�l�
v��l�*v�r�l��T�;`�S�T�;`OL�l�� ��=��l)�
v�=�'�{`��T�{e,��"vʝ�q�;eN�C��;`N�S�D����l��;e�C��;aN��D�>2��"v��'l��v�=�'l)�v���3�ȝ�'l��
vʝ�'l!���;a2�l��(vȝ��l��v���'o�v���;dN�S��;eN�C���l	�"vȝ0'l)�v�'l��yg���N0����Q�{`������a�Q�{`^�E���0��l��*#����G�W�PG�D0�v���"=��=�(=����(=��l"�EC�&�@�DG�G�S�S�P�AS�DS�AS�T{d &@�S��QS���A�S�US��"��"��Q��`@|0��P ll��l������A�D�;eOl)�0�'l	�"v��l��
v����l��$ʝ��l�� �ȝ�'l#� zd�;dN�C��{e���<7l)�"v���l��;a�:�M>|r��￐?���b��\(K:��u���[�;O{��4sn����L|�[�E�T ;E�c�6� ��[����J�l@��O^L���(*!^f�O�湮<a���R�l�}�4i����ֻu(%��!��;������l�[u��%L�z�[�imڀ;TV\kU��k�mZ'v���@Ö�u�@ڻf�Ћ��U��)���JIx�I���[ 8����A-�gߩ��,Vr��r̡�[�*齗�ۻu�wWϟn�Pz��>�ά�F�)�H�y�0�j�l��c{1oW:�z���4��w��E��d�v-}*��"��SY���ݦ${�c��6�V��֥xͣ��r:K���(l�ò'�Asm��0<�g+7C/�V��8Sn��f�gM�cћ��ձ47�$�*�V���P�Z���mm=f�$�[��LB�1_���
T�Ѩ����YN�L������E��˧#���9�n��d#	�0�=��k`J1�̺�ɊFo<yyj��b=x�)Qf�����K�Aa�X�>n�m]����e�%G5m�uyJ�$��
�������n�Ls<9�ٓp��uj�B����a����s@�jc�Hǯqie]�N�3M=�5�P�W��5�z����R�F�
t���U��+̭̆��[�W�!��f���
(��0f��1���E=w�էLnfZ�kv?�0����En
��`�b�aK�xj�Жvɨ��wX(�L ������*%[T���۫:6,�ӽ�%]Z�Q��Y�����5yv_��.GH��Ѥ��5,�Z��jk�01IL�`�y��ۃ0��,U޽2:-K*$�ܸ��L�Nn�CJ�L������7��%�1Cn�A��(���p�Ydux��7T��,���*���y�qxB+pi��4�)�(c� 	U�̣y ��/nHD� �ʗ��m��U]iP�#1k4Q���Qg�sl���#kseM�j��֓�PLA-B�2�ö\�%��KKn�� .� n���%�O����途yҙ��w1@j`Ŭ�nXwo&��u���gH�t0ҁ��d���[JK �n|\z&����tt�@�0�{gF��`h���6AݤcV�6a��Չ��E9�u��$�ѵ�cUdT>�-%Ib͙����[x��*o�o��Dn��au���� �����Kq�HՒ��_aˢL�[�A".�$��"�b��<:�;��i��Y��'�Y2�2r��z�Eɲ�Vf�Ui
��Y��5/75L�iV�fn��Fnf��*�1O�(��˂�� ;ś>̋^T�0�7�Ө*���r�lY��l٥ULm(��a`κe̴ȀiN����Z��o-?�VnVo�ӥ��,�P6��c;h��b�'�Ok�H�	�Ƶ��w�r�C����>�t��b���j��j�awu�K-ԹW�EJ�35�Єbl[�:�6��n,%:M��wbW��:o:�VR��҃mu�\4�����|B�pk'G�aC@+r�)gqj+N޳5��&ևqRa<���}�4��f���s|������f+���[�h����ځ
�!Z4S�U"��AWY�[�ѳ���ߋ�`0�K�%Qc�Nl�U�M�0m��hF��,�):�y�jm�42ѤʂfJ�ne����q��$��9���q���p�ɽ��Ҷ�0�4E�x��ʻ��U��4X�S�(S��w�{ ��m��ڶAѬ-�����%ԉ5[r��n����-�t1�����Dmntg�V��lTۡuji`�meA�t�<�1TQ��U��`ts=��#ʹi+ٹ�]���vud�Z�fm����,���(ҕb�m�^l�����IYtq��潦�ʲ�Z2���e�JJB�lUv��2��h�ywH$�ٻi�wM�I�؅vf�5��ⵌ���72飌3v�=:��cS�Yø쪡rـĆ	u(Eq��r2�-��$��Lf��n�.*ܭ��n
q-:�,Ն�b*%Yx��a�w���K��T/7 ùM��:���u�I{�81��ԁ���4-[2���S4���I�5�?Gm���b�e��.���މ��i�gj%e�D��u��a��,����N�jâ��i��KF�[�x�10��WUzUU�����|�gO]�3Rl��}�m2����m��­�	MJ�d�ھ Y}j��!i��޽I���^ج�E��f�[�2�Ky�hӥ��%�CJg&�u�DV�z2�c�7V���B��Q2���!ˣ�Q��X[�Zv�P��A���;[�	�YN�SJ?LYJ�E��H��Da���N��Q�؎����X0����ޡucY����Z(�
Z��'B�%��U�D�S��͖,#T��2��}����cN
K]o�i��R�d�9����7m\q;�N�L?��A)��KuG�Q�?�Z"x�ۤ�]A������Gl�.��Vf?��t����[dVS(�:��f�ܩ���zqɂ�|��R��=	��`az0�+U9��i��,/A��3E�M%��ڦ�0t��`R������.zi�V6���Z��|��IǷ6�3�v���x��$���@��(��b�JV�*p�Ӎ�b�(⫅QаSy!!�)a�3@�Q��Zu�tXu��`B�2��
1�8�u��4JH��1z!����JiW$��*A���L��+2�R6fc"!Fb�w0��xJl�y���;*�H|ޠ�%{��3Y[]�֍CY����J�A�~�WZ�E�n�m�ſ�R.�۸�
V�]���Vb�u��e��w.Kf\�X3)E��[�R&��3 �YaX��	{���ӆ@Q���PTSj�+G�R�͇5��C�,^#Y���Dֵ��=[�X������N�����$��O0k��:����V9kehy�{�4	�)c[Zj�/qˆ�+�J>����H�w��u�t���.�ª�.Ae��v]̼�5j��eg�oZt��;�����yqk�d�R�nm�5��-Ʃ�مa�S"ڐ���r1s.iO���B`d�j��.32i��[rZj�H��k���T�y�з�#�uC��܎Zܗ�l|#���5&dw]�y�C�����X2��:���1���B"��I�1S�X�ĭ�e�Q�K dHY��ί)�(���31���N�{��Ǜ[���[6�Ɲ�ژL��X7E���pkF�KA�V�+r��kӰ���XPR�K$��R:�F֗��w4�V]�Ċ�* v���XwhJW+#Ȥ�
[ts���PH�]^��"��P�Lӭ<��������	�(��\�c�%r9V�0�8��6�T�X2�A��X���wJ	�EH����.����zb̚"��5�+
��[a\�z��0\����KQ��c1�×D�h4w$VN�;�����KɊ�nK��+	ϦKn�e���`h�Z+.Sq�y�f�q���ݰ�P5�������jj��[y,���4eJ�1X����H9���cX��h4��Dd��r�դ}bϖV���D��Zj�K6��۸�U�_'q�t��W2Pp䂯�=��"V���-#�n�8UPJY{x.�ɣd�{j:-�Hl;��~M+�+u��#�o1ޚY�ȷB�MO.��2[z�(�.�Y�����1*�D�ZkVk��D�;�\�L`�K(?Yɰ �:N!l��&fͼ���]ص�0f�bǭ9����T+&��Y�夣P�ܖbl�CMa�ޗ����c�2��a�xa�����q���H�7n���{�@(5T��^븫%�!��
V��M�"���'']�YNlL�C��U ��4틗A�����n���f�Xw@̛���Z�*h/T��dj��f�8��j��F��GM�M��^9�nLP�$����^������QX]��;+3*kh�[*]$c���Zܺ���4���S��Z��E���af�Ew!���.֬t^�.[y[��	��Cb����-�Ԑ��I�2Y���9���2�R�h� �ߒ4�;ƴ���V)>��Wi� ^��v�����SCr��g*�KّM�CF��Do7],%�K�t�����1Q��Y�jBk]�X��K5�.@�+&��5
V��*FF���ʼE�2\Ś��˘B�E�u�є,J�5�j ����(Dr��@ު[��m�����ԾKwCk�Xt���Yg�4���M�D�%F�mn��-�G6�|��V�a�
�$�ΰ8�e'M���h]�4M��g6h&6v���5�������Fe���l̶���hRL�B�m���azYI�IJؠV�U��n�2%��вM�a���g)�Շ�c#vq�J��m�����s6��ȃB�B��8�ذKy��� �
�8Çra�y{�@**
�և��i�{"jï^�d����Zugv��	J�T7c�&�Bn����+F��/bT�2�?��w��Ì%��`]彳Pi�Ú9����O��JgX:5�����$������wfG^�����e���`F��-%�deI��&�ƅ9)�,��G-�t�OQ�-v.�O,��e�w0�fY�]�9Ri��e�/V��)]n�ƳoU;vư��?,�r�4C@H��弶�cr*ecܥ���e=Tm�x��+��^�͐��!aW[nnP��ѦR�b�x.m�3KM-�),F���Z�e�b�����6�*���53"���q�2�%"G�DÌYDi��r�p��0��On/���{B�&\L:�@�:s6��	����n3t����d��C܏FJ�1l��FSgT:�ǭ�l"j�l�Y��ܽ37��5:�7hq��t�V^P�)޴D��ݬ�g�UD��:2U��.�dއSC�"�]\�2c��V1m�I��-]3�-�uX&���a�N�����CP�u,d����J���2e�i�~-���|�z9�4k�oG+��t*U���ۅ�Y�k9R�oѶ�n(j#l�^l�O�f�Hk.�܊Y/D��"�kR	�Ɇ�t����P�2��i*moK�cT�P��ep��yr54U��#���@�����]�������4� k)�Y��[�����&���^-�q��su*gU��F��C��p��Z�zĢ�*˴��#��Ҭ�V��is��	�-Fŭ,�E,:�Fr�FH,*��-U�--`Lܭ��Y���Ö�a�y%Z���ZF�$����[JhY�VT��T��**�t�bG1ae�2�Д*{m��!��71+T��خ�;zHh���#�G�7��{���y`DE�K�a�c3r*1#a���;����l*R��0b���r�^�&�wj���`8v��Om�y3h���W�|��zc[t`��)ۧ��T�0��3n�U�Ia�)Т�dh9�����ɫ�z�<�oZ�[�(+`��R9�6��[t-@��#���)�jPbSܤ��8oŷb�<u�֪����l֣M[.����`�j�n�Z�7������K
\1��%b�>�ɦE��}E��R[��T=�7u��#z��a������,����%�F�7%$Y�W��\���nh�U��D���&��9�w"�Ӣ���+�m����2� 
�� ;������ᭌC��2��qC��
��2�v�`��-uu̬�����\�s]�*36؎��o)����[u���P^:N$�=��Vj{���%H�a627��
pc�S�&dkj�`��X��^kA���[ƍ��O�j�˰ZN�c�v$��Z7g`!k��-�"cP2�SI^��XM̱v� e!��;��G6�'c��o�]��qQ����c��m����*?=C��3n��"A�j�����D �a��f�P�1���K0�5E�N^�t���VTܐghY���yB��6��3�	���Uf�Bb<��B�֡�y7U�/usn��e��44�h��Qi�WcL��Y�n��b5��
�Dm5A���	QԼM��6���CNXC`i����(&%b��4�3VQ���.f�X�o~Q^����X�7�GS�Dml���PI��WZ��qK�t�\n5-���{Den�uɇ��8�_?;</�5l*	^i�oZ�4�4����W�YSr���Xv�qQН؍\��*8l�U��v��n�8cU�.�U�Z�-�	:�1,�BkY&�̥*��Çw)�n���j�j���5��*R�{�l�V��-�J}oj�<�BQ���f-y��H4%�4V�܂��B��3~,�*�˿��8wufਓ�^_��Ws�\���Ӱ�mh�Mӄ%!�5��*t���K��<�O&bR������"Bۚ��y�ˤ�mQ۬V�ʘ�-c0[R �c��ѡ��`:�R�@+�cIU/5�N^�l��t����)�3Vٙ�����Ima-�P�t�XrK�^K۬�������',-X � �{޽A�Cf�˷)�ur����uq�C���#���zN�ѐ�(�<z�[�&�\�Ϭ�/�g�O���.c)ُ��'��q9i8u�Y�Ba<M��^���,��)��l�&e���B9�Pp̮+Q�$��l�:�����J&�[#�Ga�<��(FU�˸�T#hl�7�aH�.�e�ٜN�(;�yNCk*0���)$�p�ue�t�6������=R�F �К^�p�I+�S���ek��a���'���(���t�	0�8N�hÛH"Hm(R"<Za�v0n�+�T���Fa��9�6d���.I'\�(��X��o{sVyβ+�����T��j3���I"Ƞ|l�K��'����z�Hӓ?���{����o���9�vy���?�����_�3z>M���:��z8�&�I�|�y�9j��6!*��-�e�Y|�6ʾ]�J��z9λ%^M��u�I[onIg-�r�2�_k�ń�G�4I�Z�[��5�a��I�b��U�6�'}{�l����̩�.��b���1Qdw,�ˁbN��Li���#��M����}�.�.S]'�#��=A4�"d�hp�v$�����;hn�T#4�]��'p���6_c}�+�ٽ�:.l��L����D��'mS���Q�\����>�4�M��P����G����!th6���2�P��-9)>��}��j|o^jy��k�*�A	��bW��V�;����q��{��2T32�qష�u*z��k���#�^�w���:p�:*�����~{<�\��^j��B+%i�p>�y�%qT�E�2��˩M�X��k��V)�9#0�����\4ś��q7)�+���[�:���']�l��³U�:R�����:�,��X�A41�;�h��A9H�A�[Ne�h�M>U�H�gB�����oq�qlm���HREǼr9��,��f�esU�_#Ü��_N�bh�����w]ά`˙��vIJ.W�R:�����xI�����^�+C��u���NZ���A9�5����A��e��|��iI�3]�	
Tl��6��h�u���
�]��tZ�t�������Y�&���T&����xr�G��mJ��h\�8��JΦ��v�}�R��:s:m���B��*���U��enR�p�F�����3�7(#���Z�H�=X��h�u�d��.�,;ب�P��{)�L]v�`�ٚ1k=3�pU�]5!tdڢQWͺ7��MS�Г5L��=�L��kU�Ʋb߬
�������,�s&|�l�݆�J|Ks��d�n�2R�M����k��
�ٔ��c�[ ��J6���{��WX/+�[����Ůd�f�ՇG'X��f� ��TR�Hwz�T�P��T���FT�W֗&%�,H�[�F����]��jYeq��ZT$[��n��d��)Br���V�v�L�ĕ��Z��QÊ�&��ύiM��y)�A�:μ����C�����Ҷ\�+˵��:�I���3����
�Z@Q�vq���[�Ӽ�äɊt�J:�N�-�F7Q����9D�wӺ9�U�x��Q�V���G�t��Ɣ�ΝwL����h� ��;9r�rsQ��z������wUa�e>�5)�'s.G�N"��5�2�F��X�uY�pe�;�a��8�^��H��u��qT�ɉ�oB���b�d[��y�{	�F�cn�=v����d�}s2�
�զ�hzV1��-y���BM���ꁧe����墛�Ѓ7���x��ڬ��YAȄ%>�X�ˊ֋�%޲vwq͎�l�e2s2��!OPm_�0�^b)���3y!}ٳ��.b��Y,�����s��2��I�ly5t���l.9K��r��-�O	:���0MH�������t������&i�M"L�f����`��P>�+�Ng-�&����$�af�@��uۋSp��\=�CIƕ<�L��0�7*�Qb��Qwp�ݦ\+RR��+S�u��׻�v�R��-�F��-�("��Qfe�.|�����;C��]�t36m���$�l](YS:�@�vP�����k�R��\�۸��{3��w���]3�9�'F��$ƫY0[�]n�U���d3�q��8�Qh�|�u�U�2GC3 ��t�Z�/@�6R�+�ok	�;^ƪm�Je�:�wZR<�]C+)�%�v�{Ɍ�I�e+	��;<�!~G�>�b��i�|���b��ɫ��z��c��Y�؛u�1fm^C��i�}V%�1�ת
G�o0]b9Xt�Q���^_
1>�0���j���w�b�լ	����:�������kԥ\�/F
��<�JHR��8�ZS�""�;��*���h[W��:Wd�Ԡq��!α�w�a/!��[0���(�xڅ޶yQ�U!�É�yp���ة��kɼ)р�{r���4�9ִ�&��*1��Dw�V>Q<œ-�Ky�Ao(k]L--]�FI���R;h��h�$\��Gh&Eޑį�����IiK��%����yP�o��_L43����j�1�d)�+��ٕa뗔�gS�L=���W.ѹX�D��t��\Y�������iT���WR���ԫHe$+.�]�D�%��#B`�F��u�抏����a�kؒ\e�	���Z�`����ﳥ̟qfj����(ۭ�ޝ��v�Ó��7�݋�"�K��Y8r��C�5|��Q�����0@�d�'	���Ϥ�A���m�K!y�q�s!��ܥ�/��)��X���5��Œ�W�<;#���-��Tb,u{��y�)�4Z�5-���ͤ�[c8QQ�4���/ax��&�9*\��ڻҨp�xm@z����"���,�F����n�A-^:v��[�h�L�v��v2��J�e���n�<w�M��w��Z�1e%c���eJ�t���}��~�u.@�� >�D.R�;�u�X�� ��[��Qp��-�@e8�N�#�2С��3��#�T7�:�9.\rl˛[io'��;��n�=��|�t'�U��o�,T�]�Rmv��WN��]h�V��X�WR��ؠɦ��p,���ic���p.��	�,ēʟ8r�W�k��,嫳��j�*8�]�JKkB�[���q푛	�f�p;ˋ��f>v���vQ��s�e���p\��POM�y��ҫ�5j��s�l�{	�[E֕���gLp��m�B�=d�\]6��t�J�2��<!�1�-��S"��C:smo������5g	����L��Y71\䰞���^�O�m����1�ٵ���hX���8�ej��<x��u�'����.�suj�oc��@Xͧ��~:=�AR�b���wM���֙7!�ʁ���u�)�O�+IWN���y�bWC0k�q���MN[�M�t����󶜅���f������`k�;BEw.|��Б��֨�X�rtx�R�΁��t��^����@и����"�ʼ�N�{;��(VR4�ty�1�.������^���������8��N����K.�#��b�²��"s5v �س��]�MXv�I�U��BU��"�5����f��hF��W,O�b[�!Y�C���h=�ݏz��� uP��į1^��%�C���t�Cx�������\�F�S����㥴�\I�S��д9�k	yҁ؀K�4e;�E)������Z*��f�@�o`Ryi������-��G
�W����V8)/����EU�!��v)��W^^ኳ��JuZP���f;��r�@�5N/)��B��.�@�h�P�oL�	��w��n:g�9�����wO�W����m.P 뻖��@T��.�[��ʙn}��Qmu��'r=U�B���m42�κ�QW[�(�ow])�������q�p���Dw\�Z�U����X��\v� �Z2���]��%m�r��dK8͹�AS\��}���O=j�j�{�ҁY�]ӥ��~�<.sS���rѠ!��.����4�^�@�(��r����2����F����8�5"N�Az��#�ε#�lsD4�A�h2��*Ԙ��_��ǧ��j2o���`i��+�erv��uƥNp���Sm
�9�imKƳ/k{)�=�GcM��M�ڦn�5��M��l��Nrb�֏�u�1;��]r��K�})fQa�<���e%F��
t��gj�h%�I����K����H%ɩ�Gf�J�솻q�t'��InK�t�4��hdˡ�!�ܭ�U��U��5>�[p^�#`���Ƕ��AnQD7�OH3%����$[k���p��u��}|�z�m3��Q�ҽ��uz/�i�0�{:V٤�\�5I�g7�\r�핹�V��Zb�n�S5J�Ek�2�!#�4na�V>Ӥ��ՃF�6�T_ E�k�H^�TX�K�ǲAu`*x��\���Y�l٭��[��=w��V��#�N1R�X������t�������'g�'�9��m \s�
ӎ�[�h�@˼��-,XP]5t�c�Ӭ����7�>��̭aѼ�^SMM��8�]]M�#���.}���%�ƭ��@�{3�d��M�1_l\����+Q"syR�m�ǔ����WMΏ1�0+mT�'�� ^܋��L�Dfн�7,Zb)��2�C���f`)�Mcy)���!u�.֙�D"���0�U"�nI�3�#�mN�2�Z]�ݾ�]��Ft�D����B�h�� 7i���H9��˺'��_�Ҧ���늤W"Ռ�Η�j��Aɺb�1h;������{�w݋���u��G�v���U�%���a����fEI�7z�tf�!3�����bH��E���ھ�zOR}�v���]�&�SuwR7���mP:�΋�a���ӡ�����0JÎ�'V�mͼ�Arb�e-���Mjo�e;�(��\
�|#��l�S$�g!�2��R5Ŏ�v^�(-�=O#[wr��zd�ɀ`ٙ����d���IF(m�̾����yϢ���G;
,<������|�D�&8������>9�bp�cn�!�7&�*Ǩn�ƺ�Y�aMX��6����y�m0{���ҁrը�(Qn=�ҳ8F�k��v��Qk�p�}W�.�$�&Yr�uj��yhghN�L@����zX�^�*V_m]ށ�(��ZR�o��E$�e�oA�Vs#*Qٰ����\��6��ѧ����w�{��ۊ�ʊ�Z*;)�{�"^[ͭ��� �i�s&��=7�YI5xe�n'�r���{O��p����n�Gm��bS�˨z��&�Ofs7�&�s�u�C9N����rJp�uhY(um�7���C�xD݄+nBs�;��k
�4YCm�<t��wm� `���F�(���q��mͨ�m<��ܙ��{}���u��R�©p�\����}4l�La�Ƶ�أ�Ÿ�̢���\�������
"��r,3.+�+�ې�R9z�Vo3�1(��r�4�o�0�j�c]:�A��Y���5��w	�~c�7KR��{�m�=%O��4����H,�"1"����+R�$�)+2�^і��+����&��lIGj6m%]}N�L��t�}0fn�A���U��Su�7��n�h��FM�t]J�@�vU���J�I��A�x��P� �>�N`F�����;75h���(�:��Nws��b (�G�G	��nl�r�:޼�a|�n���%lf>�"�S�v�
��D��O������\\�vk{ �B�?q��ͱ�2�C�:�Y�%���WJ�Y�,���'h���헢�1V��J���ԋ������B�gy�h��pݞ�:�W���S���\Ë�w�����L��3r@��
B҆��bʼ%�w�թ,eT�3�R=�IHm\�x�2�u��\��	{%a����nN]�Q²6b�w��1�ָ-���T�c��Χ#o6r�Jk���f�5���vs��U&�K�.�J�8���@��pk�\�(A���r���z=7c�Y��˂�o2+�x�˩&^V�������W��z���n˒��:Q:ۮ����un�;k�tHՇO���2!.�d���fu؏�2��a�a������Jy ��f�m��u������/�Q20r�H1Z̽R�t���ɒ���lY���խ�b�1�N{���YR�@�I(NqR"��R-���6켢D�O�R�vp�^ui׹�A�c���("�Tֆ\���\�d3+� &m�ӳ.��-�x�h](����Q1���������%2��nF�F���R��V6����׮1��jvV^�J���\��E��,v`�n*�V[������3�҆��u���+�vB�f�;��n]tz�'��WԐ�v��Z�f��t����z-� ��m�8���)����kqG���x����[cBFe�lh�����T�"�ST/y�ڔ�ꗲS�[C��̫�s8��]�%u��]I$ŏwЬj��8?�ܦ3�i[]�r����{Yk(���Oe��*����IWԅ4T76ʛ�����ƊY���襳9�JÌ�*u�;@�6�i��.���\��@�1Ӯ�7ժ��������ܥ���`8Ur�3�J�����bj�0�=�5��lc(���2;)�o,��fnA���v3:��PR&�C2A�,��V�\�b�D̔�z��ʾ�.�7Wsy��Ź*�u.]�)v�z��h�|�ֻ���A��X����
<�k6�1b�אK�Ϭ�.̑-+��;��)��YL(��T9b�؜����(��f��������^(E,x`��Q]�v�)��akZ�ю��t{6�q�`y;��D��	��ùR��>�P7�:9B�\nP��ԍ����ion�T�����MTR�.�C����瀄��� ��#[%h#�k�/�e��qY/��)"n�z$��m=���D�ÒT!�9��7���(:0�;��	  �rI8�tqG$��I$��EUTU$k䘇�2�/�nY:���|�=J���u�y)�M��;��z�éSJs��:�|�@P��}I���4���4�6����������y���r�g�i�N�����/y�w���Gw�O�y����QE�_y��á ��{~c��S� ���	A�����}�wG9�����^|~��.�d���_�;9�g|����a�+�6��6�K�G�E�G��VP�S��g�nZ�[;��E;�na�m��Z$�[u����CX>;��wA�+�n�q��~貛��IsI�q��g;}�c�`�1p$�WF50�qJ����P����q�n,fv)�Vu�zkkIꩍ��8W�RI�@���ࠍj͘i�a��T���fҺ��M�P���:�k�M3E��)N|�ۭ�� $�{Gք���D�z9�e��nۢL6P)������+1���n�"���Mfc��R�r�
�,��d8M� xUm	\̾gf�B6� �B��S�Ip�çr����v�̹��h��E^�J���/�y����@u��=����@�1[��V���\jL2V�l��D��+�!Ҧ�Ǫ݅Vwe��d�WIŷ�)2� ��w�\d�3�ٮ�z2��]���3r���=�%| �4��mv�g(�8��sB�[�L
�\�R�� q����j��Ma��+�\>\���;��|��cRx�Le�7󾾡HR�8����:Gd��v�U����ΑJ7]#��R��L�Z"뤝n���Q�ɪ�i�}ܷ��������NMb,`e^�Y��Y�V��Y2vf��4��xsR��-��u5�J��p��	�O((/�=�U�3�AT�������=̥v��Z%^�\e����0K����@�<�\������)�Xۥ��R�[r
�wc^��نh-t��B6�0�t�2�t��l� ��7��(��8�U��*rp���묪�)�YțF:�\n㳷e^j�ܘq�e��+�;t��:��nR�t�S_�Թ�HT�����i��W�unEL��Y�F�gG��`�i�v�.�:�M���oAK9H�S缕�V"U�}���&NΑ˶�V����q:�e�8[G�ȉ������v�k3�5hWn@�Uo7��X&媏�ۆ������EFz���d�Y.���|���wd�V�+�nJ
��[�v�aS�/jb��g2�>��MwK��3�& ���J�1���z�f*=C��˸�i���ԺQ���i�۫x��sH���cV�J�g*%6��U�"��Ս��UR�&em�÷�*R1�o���h�̶kx��r;IKգ��k�������e 5�z�c�+�b�y+�4�[�=k�%]G����;6��D����CoJRX���P���漶��f�DV���McAR\Q�؟f��Y��d�X���Zu����#rB��8Y)��@9��I�nHQ�$} ��,[9Tz��B��n]dA K�=��Vi4�V"��U`�oc�N(����x�O��!�{Z�C����^Yk�6�E�v��"qb���m�*��r���N�]�n T�P��1򇱠6<��k���wp�2���I�lU�UԆ�u9�D^��U����������kB1H�FF�t:��WlӨ�Pй�R�r�[W�L,�Cw��������Iaڶ���r�3g�����t�U�B���EAjG�iVj�pv���"U��Ҹ�4�`&4�������]���6��5
�իp�}�vf�9��f�2 
��e8ު�����=1RM�q\�릚�r����ڌW�h��(A�+��.�v���we��İ�nż�Fդ�����I�lp���Yn��fK�˩*a���<��s�I�v8+���7�[�u�Tf�l5}{4U7jY�R��;��$2��f� 2�"�]wk+G
eu�y;
���܊���(+ή�J����Y�.�˛�J���f\��Y
T�j�2]y^h������wTvh(��e��6uk�|� �%��u�(���n�w+x���ao��>u�Mm[�����]���ch��Ȣo5�W�k/\���#&�"�ͼ�Y毕����ϵ�+dײ�Qv�xdBJ&�k9d�!�j��&�4��K5{�q#�q��dW���l������t��S�Z�n�z LR�]1m�zE
�w#���'1mM0}�l���i@/-7��8�묉��;\�ξ��&v�!Z��#�ȳ�];�wA��  �Kr���c��#.�7vD�8�#7m��w��vg�|5�JVV>�Ks�W]ê�@�%�C|�(;�R��yO����~�H\�)������*u{�T`N����ѓb�q�:�PA��_�5&����{�N��8��(~��	H�ˍ1��go��7��e� �c��IV1��T���5|n^�ۤ)�q�J��j�{RQT�)�$���+�������wQ+��.*�TTc�~u�H^.�Xv�)�guN��I���Jt�}���Jfn��Lq�x��䮎���
�ɵ�U�����.�i8�orx�Y%3X�<o#����VQ����Z�I;�Cr��
�T�����%̸�Γ�r��ky-�2����IL��.�]�d|�]+�	V���-��%ve��i+8m$�"if���*�w���Y(8�WP����$�:���A<��&vP[]t+m�JR�(��7����� �Q`�T�^U��7JH��#�,��~������-*k��I���RK��9�VPŝ-T��� F���r
�^^wmH��q���i�|�ߢ��][7fW=�n���
�(U9�5�|��B�0�|��I�U���s��%�n�뢱Ԅ�x���}�{$<tS���DP9��CM����n�Y�Q�%\�('�u|�M
�3�`�>���^�{�J.좵��!�2���h���+�K%�Ԍ���<8,�V0Չ2SU6���g�u���J�,6����>v�X}%l�Hn�p��iu�(�}[ϙXy%�)��ڣ�]
�c��찦�Y���1f7�C�V�5[�Vq�U��7��5����2�3���/b�|E�Y�ٮ��#HLJ�+����P�ff/��!w3��.�o�R95Lf�؟MO[׌�)ƺ1����=#�%ј�+C."�-h����5᳖�8��hnQ[#�ƭS���t���3�e�%h@Z�!K��z�g��x��y��}t��O��a�W����y#Bq����u52�e,8M���8KQn϶��v~�x�r!�\/U�%��Rt��˵L�����n�.�8�]�c�1�q�0ej�5�y�1e�pV��R��8�dkq�h�᤭R+��nƜD�xay��b%�T�+W=L�*�5v�G��>6�u����^ӼV�6,��x����W�ܙ��Ӽ��M��P��yV`97�nrK0
G6މ�.1<TB 	jmC�h��3p�^�F�#F��v������#u��J���T�
�E��ʾ	9�r?������V����B��;�L�����M)�n�8X\����e��jͺd=��<����g��wE�V�U2
�a�RbW�\�� �+��ۨl�emc��V�hg6%ݍ��P��G�c�v���4���L��shQ�H�����C���1��Ŗ�����6���� �h:�@��(��G��D,hx���4[2�HJ��1�ݚ@���PT����i�,M;خ��ɬ
�vF�B	j���������*+�y�S���n��*.7QF�VqX㭺��%��5��
ݗ+��@ڦ����z�\GT{�'_*{�銔S%~����r��Q�f=YW��j����>
���t�0�oF��J^��7�����g3M�
�J씛��qH^:����U��\CB[\(�J4�����.t;�e����z���F�
\&Kt)0��[ł�E,
��-ߦ'N|��g���7�r�i�4)\:�c�n�3��;���_:,Ɍ���օ�u$lv�Ę�]�2�,s,�ҭ�����zr�s.�*��;Rt�W�d��r�ly�a���*�>�׼�;�71�odF쐆���M�fN���iQ�Q%���xf��9�qfn�V��E9�xu���g!�V���K���\�ȑ��W1�\��"�	��@���x���ĩ��+gs�eG��pb9��)n�8���d�n�c6����D
����Rq�}3M�eŹ�ЂuXē�H����&(�h!����j�U�
����\�h��:R����UVӺ�-,��ui�r�����p�]*ۓ$���H�m\�*�Z哫h���>ut�t	߬e�b�a��6&�Ǒ�Eٮ���n�+���J>Ēma����̩��X/-K�.��*�`A��;�ӛ�yi�(]6e����U�֒ajhS�n�d�m�PS��x��&ލ��u��F�m��q4��g`�`qs=��teX�F����Q�╫gv��x=5�i������kc�ڳ;4q���Mފ�o|u�Z{r�̛�e���r�Ԥ��������J�)W��T���γ �eF˔��{{�2 ��]y�):��ʤP.���6��K����Z:h>��B#���VM5��5��'��:�\�B�&����e�X�R3B�U �ir��o�]$l
�E�*Ev�j�'���'7��s̻ű�� �cV�O��t�<ө�G�rC��K���r�ݯ���^�GJ�*�k�_^Q�b���H�{��F����V��9*X� ���\���o0�-�\�
�\��T��DНM�ar�}����k�)�2���ȳY��b�Լ��}��n�k�Y۱�Y�o�vhf�q���nL�0L�"zh	{���5�8���Ϯ P�ؗ"�.�mnbRu��T��n�ky,;aH��J])۸�=ʗ�vc����9�}{@��Y} ��\�b�z�FU�u���Ӹl�T��|1�{yY�wh#)�)�k�����営����'R�_M�Q1r�ژڎ��[�E��G��qM+Da�5]ב!�I"m�ttvhX��omk�ޔ�KoΙ���КpX��M�v.�]�*�bs�G�T��st�,R��qϢ��k��C[e�ȕ�s[]�=ɲ�=Ꙙ\ERK9tT��
�k!��Miۙ��	�ñ�(Cr��T��J]N��_ݝ����XI9�s��ּ�,ۻ��Q�Gg�/�<'�F��&�}�gi��2�bG����u��1��5��j�m�����4-{3vfhAUAB8�E���|띮�j�;�+����ؖvk���M�&%�;V�[2i�zaJ�O�����֤�X:��Z�|2�)�U���(����I1�*̡��.���r��%�m�q��и�C+7m�����K�B�����E�I���-������4 튦}��V�R�Y�e�yݴCҜ������x�`��h�ݬ�ʝPZ��d'��v�q��j�IX����Y6��/4�G&�5:�2�:�s��3;Y�*�a���2�.��m4��}�-%Y67�J�m�t�>C1�e���9f�U����KR���]];��D��������m�[�Ǒ�r�9W͛�jJ�ӗEr��j�K �0�U�F�Wɢ��n�����5H� ص�-�h�̦�y��)iV��)W0�Q�i��Ze�{�h `�;1�5&�n�u���Θ��Y��'.���Y+�I�o-ԣ�IV�y��q/]u��[|�&�t=*Di��6��$�^��lu�aw&��CG"}z���6��l"T����K,�uG�:��z,�Iۏ�6i��82i��(��:��I��gK��.�Pk6��q$�ஞ9t�0���Ww)�oB�A�q����������ZQ��L�ݙ}G�ƌ���=������]DUǎf�ݦ6��k�K)��x���(��[ʥW��&������#,�N���У[h^���6C�)�i����N�ɻ��{�͡κ�p-T�
�s�q�t�S1_Wu �-�Y��\�\���4�ޜ\Ō��,ƃ����<�RE_;u
G�WF�mͬ��D�"['Uw](���d���#-L;�s���'��*R溯Qj�Ђ��|�	9�̱l��	�����n\Rm�;��U�tF8�^��:5��9�
e�I˺�׵�"8h�ڑm�gjy"��0����Z*�$>�Q;V��y��p�%�X��K+�����w�]N%Hie�:���%0�룚s\�ٵ����ɳ[���k"}H-����ɋ]A�G�66%���7�{x��?]K��YT���'.6��� 76ٺ袮���I�V�ɵ9���K�p���V�`O����Z����eՁ cM��ISu��TǄ֩���6g�,��9ܨ��wxu�w��3Xm�%
�u�;HzS*� z�ڣ1�7`(�5R���H|���S-.�Sَ�E�}��F�rk��%�KӔ4��A��"�B`�(���7;GXt~]7k#�3g=��F��o�/��ǿGWf�����Z��׸����{M$\�g!�t�6�������NݺWm=��U�T��i��k�qm%��g_Q��5:�˥S�qgb{��5�u2��,A.��t�(U��O�С�[R�1����*��4"��Y+�ş��@��1���_h�����&*�%YYQN�"�:�e�CB?
qSx�;r3�̫7K�
������fQ�E&e�uإ��DՉW;��|҆+��ժ󌧽2ҫ�V=��gd�)kM�7���U���!ͧxH��ِ.x-�T ����Q�WٻAq��	r[��4xZĬP��ƥ���g+�!"$���!�|��?9�Vj[/+�ݦҌ5Ӟu�Pp��oHNY͵����`�BS �F�T��Tޘ��X����-Y%,�N����	��$����\��[�X�=<w���W��_���_��"�
��O��x��_ֿ{�~�~��|?���Y�_���~?������z~>_��ߗ��XS�J]�d���tȻ!I�a �t�Q�ILP��I$�*) ��/�$��G��E�����I�Bt���h�@ Xm%�J)�TX�M]*��?==�.�'{��Q�}s����ܟ:��X�ejTiUu��\\
��2q�G�bj=9�f�lŝj����m�w
�^wZ��n]�ӡ��^��.A�Xִ�I�=�$փM�����k&���d��nnƞv��No!�b��؝In,��@����������_bf�!2�t������.�c�,Q]��4E��nh���%T�x	R���k��ާ0�2�3F&� ���[8X�&�2;4�AJK�7�������`��[2Q��ȇn��k���\T�TM�9r�i�@vbκ T��<�vso��*,�=[����-1R�V7)��Q/!�z�.& ����Yٲlr����^����5�8d΋'+�4b��c̋�V�ր�l���va��Dz�u�7/���������ax���8�$���e�}��A!y�S�����~Gӏa��C Br �r#:f�ϲ^8��w͎e��Q�ڌ��E�V󈵊]pϥ�1��U^�4��c�0�n�n鹜�)Ā#Gc�2u���C�(s��|[��R�L���;��n(�9�l_k���<��K�!\~+MA��l�\Id�8:�)�����%Y�͋�+�9)1��	�|�e-�]B��
�AF4����@�Ӥ(/�$�薐 �A���H1N�T ��l��:(B�6����lOB�T��Re)%qBB���L|�`��a��!4�$�P���ڂ\���*Aҧ����4Ci�4�#E�(�4�H�h����M��e�Ф�D��hPc����A���@P4_h��>�4�@Ru�AE:�76��\�
(kX�)
"h)j����.a�1B�!O$���j�$�(Jf5�
(Ji(F���i�������@hm���F�"dJ)�hk��0��tR����K�B�������Ҕ��TN��5H�5KAT-"rD�6)�
(��
�*�������B�hC�)4k�����Z���@�b5� �͞M@�\�j�B�
�5��J�(y&�B��"R"�!�
ZNN��h�)�*!�I���%uj��*��4��E@Ps:���Ѣ���.Z
Z
B傚H��(������I�j��� �#H�TőH|C�0�@O��1�]e5V�a��������="<=#3]�:X]�,����
�&�j��九S���P��2��$[��ӡM���H�&�A��:*�IZ%%����B��:4.�P�UW�z��5�ngһ~�Z�80k���3�� ؞D�M-���u�=��Mg�?�yc��^*�'������@���L<�͞E�m*���߲�n�_GEz���Ωܶ�����ڥ։�KU�=�|v�7v��zwF^[�O���`�%[�Fp���]$#��w}=������g�N�]���X��]�S��GǷ��?)����S���p�k멞RMݠ��΋���@뫼O�����:�D�ݾ��t���p[%��q�\�gu���c��L߮o�����/7=�n�ЋP2����X\��ˊ�1�ɑh��7�cl�<�%��q�ܠk{Y�5�8k2��7��+��(����� T׬�^��W\����OH�́�t�� kj��z��6NG����T�7[�_w��{į�+O[���W�;����ꑟ�s�5!�1g+(-#�Kc�2���E𧼣D��܂�*W��d�w��_�b���)ײ�w������7�h���w­�_�T�{}�����22����`N2���b�� �٣�J��ʐPӸ)Mw��� /`v�r��� &}ٱgg=棡G���w��^��=>~E
^����[~Z��ߑ~�� ���m��w[�)�i��2}T2�υo#ZG���ʮ�9}R����%��=�OL}<�V�{��P��������;F��q�����Kg�5�fO�\�g�⾮��W���^l? �B�S�+��'ǘ򭱔#�R���~��&$m������U^r���
��/���=I�믗����Ǥ�ݡ�>>�D�t��#�v^�ǻ/b^���r�b��5=A���Q!�0i"��V����ƽ��-�¾2]�M}W��k�M��W�.�*��3ϥ��5�L��x|�匿�?�ݘ�Q�a8���9Doi���9q������Li�1�g$�ك�;'${�7�{2�T�������%�D���˓ק(_q�cDϴ9 �[���MJN<���+o����х��x�y�N�|]feL,���ϒ�Κf�ˋ	�f��jf�LhĴk̭�S0TE��_myh�v�����ŧr���.���3;j�r�y|��r�FC���+��n�ӵ��>Mq�:#�9F��9NM��5�Q}3��ٗؓ˥N���/G��dV�u�x���Ƙ��<O,���aC��J��^��,�K�P3�H#`
s��za�w4��f$��v��x��UÏ2��^{"O_�@46�R�7��ee��ןN������*{���lf���L�2�}Gƫ�B/�`tp��j��y�[��ս;�s�~�,]�����9�9�	Z�O�����������qO����i�ԯK��o�=\�B�����jϐ͗z}ٞ��G=�_5��:���5B��K< �]�n���&k��k��E�ͨ�C9>
>�Kɐ��1ʄ�1G���v�]~���K�_���
�}u��uu�-��Z�j��\���)�Ze��+�p�/�z�a�V�f� u��Χ}�m'?z�^��q'�}yc�Fd�4��zh�G�mg/��Br���;߮U�Uw��*�w�='W��+�n�"�	���������mZ���L�X}��Vܝjtd�kͬ���s�["�J!�� HVm�ʕ�8����-u__����X�]���We����%8��v��H�5����k�*�Wm��S��t��}N��ΤvJ���}��׹�u�N��_�5���~��%̇�?_q<ͣz�"������$�&�(o�w��j��wm	����b��=�/��U5w�9��'���^i;Vd�'/M�ʞ����>����`�4����{��=W���|gU"�� 3�Sގvo����y3f��}��K'�}~�X� �YW��(�����p��W������&(�3�8F��}��S}�]y�M�����-�=�W{˟u*�-����e���Bg�:���=�ϴ�T1����t��uV���C���F�����}d��'tq�=o� �PQ[������&�e1�5|V��	�cf��8���q;8�u��;�^'�6U��¯{=o�W����˗5�_�^4�F���.w�E��=���y�2�T����zߎ�=�Q��`�ƪ�i#�+�|�Q���=޷��?Y5s p�u]�}ñ�ﹾ nûmѡ�E8<ǘ���v�����s�3ۗ�O4S{��G-�Ç�s��@�#6I�*��xpv8�v��J������C�� ���g�#6�f�
��;�kO��t�-}�&<���7�X��Bf�}��_��y��GķКʵ�9Q C���C�yuV�׋�-�
�g^��������/G��=�*es�bC�>�n�����M�Q�/���ǳ[�`�4޶�|#��q�^=Lg���Q�t:��&f�����\�V��{Y��,��Č<�W�6����Y�D��My�a�6vu��n�-7{*��7�{��(n�S����y71*�d�y��k��y�՞�a�����j����.:�����2v�_[0�6�]smV�~�Dޤ}y�o�~�~w�ϱ�7`�o2�r����|w�a3C�w=�<UO�UޒӁyQ���vU��>�G�؆���y�35�~��u㱼9�&N�3�(�k�T_T�wj�K6]m{_��R�؊�no&��3mV5sjԠ���Og{J�)�����P)��f�ڇ`ڊ��뮵 yr>�U�J�y"ἷ�eқ4]�7�*11}b;��(�t�c@�oo��z�����\��ߠK�L;�Jػam�n��6p�Ϣ2�d\S5
&�:v�{�w��'����w4q7��@m���m�W��T��~�^Y���/�����׌�}^���=y�`X�ke��{T����G=W��xl�X�y�o#�7�_�t�=S��uLY�])Ա�M%e��{[�"��ֺF���	�e�W�]�ا�ߧ�y�����$�d��L]�f��=�GSR�Ɖ�>r�|�8)�����;|�ո�⽾�!��������*\'v�Ek��u��� ��z<�} @����n�w&�'����W�/�,�v�<�	 ʧVT��e�k�^.�V��f��C�,�u2��"���ߐ{PŔ��u]Oo�|f�2�[�Q_e��׺{�����r�S�ҋQ�.�'��_����]�����眚����K���O]h߼W1*M�__y�o�������h����f$�+��6�+� �z��~7W������&k(e�e�n��Cb�@����L�u�/;�P	�>�@\��,�`,�l�"��w�4��ٹ���(iU������c�����gmD�V�y��'%��<;f��W�W������y�15��];Z�9����9s���~Tw!x{���DX��0v�M�W��U{;��j�yO���uz�H�,~��d9��L��I�d��"�WU�2&�	���T�/r�����h�^��Ri�GL�t�y�|��}�I�q^�	{;-W���+W/W�[4V��ŃaҠ#����[��Oo��d�Y=�D������?]礇���F�P3ʬ����gӚ�~��^�2_	��1�ZI{�}�{�<�m?|��t��]t"�a����[���rC�G��,^�q�O}W	9}i�����0vk�Ҡ<%z,�"޴f���w6&�0�3H�9}�ړ�`0Ǎ�3�dQƭ1��Ʀ�f�lր'�������{[>���>����1���t�/{�~ኼ�*ޔz�E	ϗҌ�+�ɬo����ݏ��~X�]3p�=$�:��h��kʷ�OP��<���R�kַ�'���%��u�tތѐ�[�����e-uKlr���$���[o,�.���+��Z������]/��I^��8q`�\D�8��_f+Lj�i�p1���^S�Ϣa�("�#�b����6�m�q�O���^�r��:�F�!tf�*���]I���=�k���B�lU<���m{�a�7�/�W��y�U���˩��ß$�N?zXc�"�[N��{Cxi#�i�SF*���*�o��:��K>)eNsh�l�"w���xd鋟6���a��TT}�n�9�������*�8gTB��f���M��O�����*���ju��v��&�f�Ρ�s&�u�}�M���:�t��Y���7Y^�T0��/oFuo���y���.x/��6Bo��=G�aVއ~�什&ז�a�y/�if�Q��G�dH�i"���8���@�>���=6Ty��-v=�el��y{=�q��{M�8��KUڢ&Y��_V�>���|߲x����6�ir��C���x�4�D���uC����~s��g��s���^���Ԯ����}��y�dÁ��|jS� ��DB���y�]��ur��3�q�3-�Cɪb2�W`��u��od�2����X�Π�xxL��H2�L <�����eo�b���X���W*��h�_��ѧ�����+W��3�n���M����;ǻ	n�v�0h!�ީD*4�0�i��k
�=~���f����.6���c,�W�z��hY��=�	��k��{���7�U�Yw���\��O5^��|ƿ��>���1����[W��ez��wTiT���F����w����8�i��h��l��2L5�i���u�>φ��q���J���^[Z�����k��>���+T�d�r�Mu*�D�ȯ������	�P��3�"��_]6>��!1DSмs1<X�tv1�NJ{P�YR���L�6���gôuW��͢/����1�B�	�^���y�%f�uHv���@b��^f�ϝ���E�~b�������
�	�Z�nխS�Y5}����j�sQ�{���QHU�=W�:a�lM�"�{����*J��&^���I�)f����9F� ��]��y�G&&���|T���2�#�ksng�ZNR6�*(b�m����5ɠP�tx�xd%V9��*�
�=��4�xBŲ�Is���82Q�.&4�'q୦�W����2��Rj�C�rd��w'%�����݌�Tu���	�f�I��b��{��b/�vuz E�c�'�-<�Ӑ�pu�]��;�=�t糀◇8|<U)�W�[wQ�M��{y����-y�ޒ�I�4��ʿy����|���Z�?>�O9��q�w1eU�v-�r�d�v�t/я=-aO2@o*�=��ۤ�<�x-��1~~߄ȵy��}�)-�1�<ѷë�|��n��_��՗�s���w�ޓ���Mz���)L�f�|{b=6���T#��e*�#О͍b��I�q�y���$�S�zu�~�o���n������hk�N�5�������ߟ��&�j�^�Y�w����ۄ�=^�5�sN����E���}3��U��N�V�׍�2l�ӤQ�3Y.kv���Q�ʙ�&Й��K����ʺ?���~=���۟�������o�����{{|�_>�K4d�\'�<p��̛P��?�)�D�WnI�`�ݚ���L<ވU�S�o��%Y<(╼a=�k�gf��yKsYY�^cka&�}y���bw��I�Z����]o2o+V��K��s�i�Ξ>�zw(�R��V�j�k{�̬�c�d�Ļ�h
�x���D�A��\P�~�8�	��w���n1�0b7K]tu��tg�3�җK���]�E<�ψJ�]���#=M@�ʺ:��l;O��[��p�����e�C���-�]d��ح�"�wF�Z�U�%K�V��6�ۻz��0�cu�$�6w�̝4�T��0�װEH��#;}Jgi���q�v��S�i��f��'_M��H�@M�QT4fcA��H�:NngYt�ZC��T��1y����T[<�hl��Ϭ��������|)l��"� ݸ�GcT��v�@�دgo3%\�1�VnG$�x�!�M��}�:�k�Z�=յ�He]�)2\�P�>dQ���"��]��m�ͥ�;�4�jZI���v�QF�݄ٸ�셮���;��m��ɾJ��aJ��~Ζ��*f46;ZVİ��ԏS52�7�����	C"���vZ��]t�}O���Ξ�,��J$����J��7a�:��G���VѮ������}�
V�]�!}*�K�;t�[��ҝ̮[��n���
Qym)ց���m�!��]6����[���a[�T��u�2sh�ga76R�7O����X}��![�CX��3�k��g
����eM,X��j��%h��4;�q'�q���N�d X������}:�=�/K-8��һ���;\�Z��<��ԣ���	Х�l�V�v��͡R��|���ǚ�W�z^�K�Lq�*�Z.��ߜ��̢&�<����N�)K/'9��jH��NJ�e��8���ms�W�IF�v�X�����,���]��\�3R"v��=w�V�#�֢��ڤ�B��QP��Y�si�-�BKyש�Q3^�+��X�<��.��m��$�0᭲��4|z������Sln;��R7�MZv�fǚ�����S5b��b�J�[�rC���w�,�S������ռ����^�q��c.ܶg.���ܧ�`�ٕt���(V���ާ��������t�U�їLȰ�������:^w!E/˻|+"�aH���k���>ߵ6��^*�X�+���q{7�fs/�B8�<��=�4
D���Z��]��f�1�K������*�D��ہ'*�LZM�X�"�8/�Ju��Ҵ*_'M�Ḵ��lp�Yw��0έ�!wׁ��Z�:]^5ƶ�E�1/��-�^��駮@8�ң֨R�͵��Q���m����j�d�od{+nV�����;)���b�;u� t]r'���NoO!]�4�PPD�]ҽ��]<��xl�SN��-6i5�`��x�ϭP3$O{����v��I����J���^>�"{�hj��))�� J
R�(�W���E4�X4CIJR�UR��JRR�ID����h������bhhh)()�
&ff���&�"R��&��$��M-PQ@SMS3	�T%-5AI@HST�44D45����4�
�&���ݠh�ZZ7��"�������Z5z8p��T�j� #�Jm�L�pƹ���\#�SAƹc�nb,cDT�[b"I�ц"(&6ψ�76�T�j�5V�A0�E�뛑���&�js��ٙ�p��.�b&�� �j�Ilm��Q��:5l[�c�A&-�ź�M�F��*���@�B������ܠwCR����(^�C(z�l�٢��ղ���޵5Ϋcs^�^�G]�y�}c�ldnE+V�?0\�-T:�s#[���w�	ouf��w�������l>����F�u~�]O�DtGhC��D3����v]�x!{��wŭ<x&���$`�T�p��7N��z��,�`A�}+���fv߃l7<4��<�>�U�e����̑	[��B���l��
�C��	ِ�Ts:�i_���/����M���>�	gNqN}���Cd5}��.����j���t]�q���y���o�<�}`q����~�DP�2Rv�ΘfF����]FM7�ǩ�qy���6�:��m��U`�P]�h��_9�b�Ϧ�7b����=Q�f��y�Xv $L��j�%�H��|�kj2�;'-�$���ߗ�������{��_��)?Z��B���*vZ�Z#� Ž��9�̌��N�;��^�g�F����c@d�j5���I�鎣k_J�NN��-V7��7.��n�b���V�U�|�z���3���?�r㙢�y�����)���Y��\����*e[��2��0��q����g��P��~�}A�1��/sЗ>�a��x��p��_��31��������Ǔ�ey'�r�]�g#������no*}�}�J�-�J�4V�����62���m�
����̩X\����MK��<;PZ�J��]�VԻͮ-1#��E]�*f����K�޽W���l1�3Հ��T�em�e�-�M�_|Py���С�l�����wt@�_�����k\l�*W����jKm�t<��ᱼ9�?� Լw=����_�b o������	CU�ʃT�:0���gq,-�j�P-��	ɛ Va��h����O�U����?�W}�5�^J_�?]x^.��a[<|�����s� �'A�J!��v�]p���'n ��z�lo4/�叭�����:��Dw�:���v���j[慦����0C���n`&��S��.�5C�mG|雾��ݥ��E���?��ϗ�9����^�I����^t��`A��2��:���^u����M�����@v���/�xo�Nv˸��n�e�Kz���;�fI`A�n�-�=��C|���4�<k��ȭL��{�H�7����x��[��p��|�L�'���p-Uˀ����(ߦ.ݯ$�b�O��נL����m�0ŝ�M��]G�N������&���oY�Pe� ל�3���Oj�P�&N��$o;@�<ﵬ4���O�dKz��P�V�,��
�R��c��^��ԮD�r�a,Bޒ��Z�xy�</"�#J��Sө
c)_`���G��9;�*^q�v�=%3����"1�u��g;puM��7�{���P��aE�w�� l 5���)v(潧�8�e]-��6)=���yi��"kW0z�#E��]�o��y���E�Ԯ�e������D3o��h��|_���B�x�c�mE'�Ô/o�V�o!��yBt�M�J�\⯙�n�DwO�#�����[]�2��V�j��6[�.|��˔{$��&ᷪ�^��|�}>���F��ƽ��q�4��T><ː˨d���5�����y�F&.�2����䭚9Ô�ؒ�l܍�&of9���/ӍR镽K���5��m���%�u�ʉɮ�Cs,�:�TXR5)�|uR��#y��8<�q�d�Ə;60{U�[<��c�L=��
�a���=��_ۜ�+�ɗiN�E,�3�%l=��V� �G�5 =%>Ss�8��<&���d�%�sb�a2�S0����@��b�J\m�b�t�j;�e���Z���k������OO6�R�q����c�l�a�39/>�\�E2�:v�z�I]cq)1qi��Ĥۨ3��3�2u�$@�� wr��Ɩ`�y�aex�ym��`>��sL���U�F��� D�5c�ޢ#��̳��WX����δ?��Z�>`+I���d�oZa��a�X��>�Y���(���X'Ɂ�}�N�+f]���KZ���oc�X9��K�Ɏ'k�i�k�oF�8�<	�s�C������j`j�������~4�e�Hʖ�l)Ob�YD���Qh���X������Y4V��`�1���Ҿ�V˹;o���`�W�5�=�qGN��X�0b[�Y͎1"���wDp�P�⁳����k�yV�6�c���M�3y;5\�y��\��w`0N�)�� ��KP�TS=� ��M�%
܈�X�LY��A�;1�ݍ���G3�<�)M�w��={�9N�f��'5M���n��	��k6�Qו8+�Vq�}�k��d�o㚪"[�$����"DҐ�P	]xV8I�dÇ]�c_-+�i�z��C����PQ{0M&D�9��>r� �T���i�X�X�R�����j���+!e��D��(#խ�Wr'-eD<�&��#T_�����f��X*�.ż�C	l}䚕�Y�7A��0@Q�M۞J��s�vz���ek��`e�9�fƛ�l�L˜Z
��uH2Fczܽ��!Hd����J�W�㢓�	Lsn�J���I��I��Ƣ��g�l����3%�1��*$p�����;K!8!2��V�γJ�p��Mn����cTsu�c߹��T��Cz�"��9�����:O4���������WD0��#��NB�%�����yI�� ,n<�8�j&�M?���l�:�{W�%��,~�~��t�@*{�3.=پ}�����)n�<�[�
Ƅ�ͪj,[]@�ԋ���z���%�ʀ���R�U��C�5�*�+��o0& �RWNed'm�:7���m��]����̘�������=���wUi9p���q�i�J��:�u3����.���D@����6j@IjYa@�Ť���ʢ���Ɍ�yԻ%�CQ0�HZ��춦Ǳ�&��1ػY���\1��O~xJs�����۲e��SzS>Z�3Lq�����v����Ma�b��i�g#if�PkZkC\a�Սw���C��֯�K��{���mZ�����:��-n��gDԽd���)��#}Hsz��掚>&F6�?E��cL��ze�e�-���
�춽�{e�q��4!�{��uC5*62���De�M��׬�L��<X�>y�:���y당�Y�f����383eg��c�
�������4�T�y�E�.aA�+yE�*�[��FeS�l�~��3�+gb���<r�"��ݠ�����g��16����׀���Z�:&���<�\�<$��~�wK���S�g�RRvl0L��|�b�U��m�08���F5@�\੫�O%������̵j�"y8�r��/z^�]��(M�<�z�<�P����N�bz�54c���5��a�]t}�=���1��/XD��/"�B����)<Q�-��@�����L|�v
²���b��-E]4�.�vҘ��7V�lӗ�eо#o�[�Ƹ�jq���:o �롶�!��e�G�m������ }�5��m7N�w�=�>��F.��J��yN�Ψ����hJo���t%��{u:<���~h��F�=Ov<������R�BR�m�����O8�?I���ӓ��^ժ��mS3!��Erq�US��ӭ,�Ob<٫�0ąA����ب�h��� w%@�0Qa�R}��<՚y�󲷊8��koLgVL����v�t��B��M9�ڏ��(�`̓J�x��·�>3�K���,�1�q(���o�F����\�	����b�	)����zݶ��,x��;O85�3�C3���GF��e�D�L�<�:��?����57����j1Q$Y6�<y`c�4���/n1�rizA�3���S�~��u�&EQ*�; sBs��.���x������w�t� xМ�9���WS���t���$��9n�P�i8��4��2���#C�t��3:��04]���o*q�	�[33b�n�.L���4p�cۻܬ�Fϲ�_���sU���k81����S�"��&K�vFO{��yS(���Z�4$:b�d�c�k��g]��^oq��ة����z���4E�Y˸hA��5+GSě]]��E���g�K������L�\ݳn����/���blk�z� �0+_;Jy��Ӷ�V)2��S֏6�pG�.����ԅf��AM3�7:�L�W�u�lnwwd����}TT>��$��w��ϟ=楘uu����G���]�4�m�3CR�����dV�R����Kry���q��gg�9��:3���i�Ӳ�S���,'L��9G��4����B3d�b�D+1�:�0��Ƽ=\�9��5B!�;9���+��=��O���J������k����z$��%	�F��$ޑ�g���yZTw�"�19�`7͜�ܦ�h[%�HP��f���s<_�cv�xV�a-�[���p]$9��*�����"5�׍�=G���w���XfÅp�M��vj�rk�l�����&uuY�z���ͱKeƢ����C���H���zo�4i��+�g�c��c�ԛ[�Mt᜗�u�X��W�A��y^����^=z���-���dz6�5�¡��\�]C$�\3�yPA����m�����;���v1_�(�<��O�i�����9�Â��JC�<�9��]�!͸#��)5gp�mw�;��9��0�f��:�I�x��;7Qc���ڊ0R��ٝFy��FD#��*��k�Ý!�Κ�Y�/���Z��3���F�=�5�nƎ�+&�F��Y���:3iV�E�8��73	�2���L�#�cQ\��w��%��5t��U+����x����d��e��&N��v���0�pUқ�����Ӂ���h��P�N���c2��/y�G�V�±�6�����n>=γZ��*k�љ+h	Q����u�n.�P*r@ (���^=w�s};<�;=��n�j��!>�zfs/����0�P�*�ӧ�Z��� n�Vr홴+Z���&+5�@�.{�a�;�`�L���&<�^��v��QL�3������% K�P�S:�ٙ��J�g�������8C7b���n"�뵻9)�W���XX����&�J���W���q.ӏUNM�i	t�n�V$�>&�a�3F�gCc�z]�Q�vN�����c���6.Yr�Znp�S��܅s6�F�Ԛ���^zk�1����L^a��3L��<�0�ٕ��ǩ55���h6�+Ko�)�L�YUS��kx�3�k
�n�l��4����zb9�xܷ1�j�e��Tν�O�C?��Fs\Ѯ���9*h�Q��7�P��R5m��;C���X�QTq𹭔�����[;ws�O�Ɲ��>�ui�`K5��[�
y��Ԫ���^�!6��=�[��O0�}ks��T}���}����=�eM�f%�D��(�l<[zJ��l�U���88�k��k��[_V���Z�(z�z�Zk��7�D��5E�"-�z�������{�B�=�N���1�f�Ů|[w߆_�S�=��ߡ�ԺSS2��F�sͤ��h��Ҭ�8v\4���f *ΨQk��e�7SA`$�:4��<��=��H��5a�idd�he�GL��Kc<�aʋ#� ���6�Un�ֲ�r	g��T�K�;���R % �H�P�R��}��]�NJ��$��B�L(#2�nTȹ\��H˜a%E���y�V��|ײ�R���v�ϝ�S+���n�d��׻�Ѧ�=�D��&��� J�m�o��mr��)�2f�l��~�Y�{�Y&�'��E��t_5&��w]��f��4�����~d����8��$��S�v�d��{r^�Wv�0�2^�Ii������W�/�En�2�ތ�aD��ې��V�d=]i��r�"C�l%i�c����/���v�jK$�o_��T�[��[n�2�K�h�+��r\�E�� s%�� ZV�˶����h~�!�qz^y�Pʀ)���<=�=L�S�9YB�bC��5���;�c���5U�oC�����<Mh�tx�q���c���n�Gi�[-׋�<�25���8�,3��z�d>��5�E��7Y ,{N�b���~�c�� !����lu�{���nns��^����w�1�K<�덉�b;���=�N��*��Xw�~�Z��{l3۶���i���O7QBF�9��HoT�K߰�`]ꏋ��Me�hMO��g��܃�Ү�RB���a�u�˔CI{�r"�+jU��P��m���~H>�Os%4t_�"n��W�0A<ܺq[[n����yXz��^f5�Ӧ������E|��&M��3��������� 7��-k�̓8�;ŏ̺`�l.M�%�
a:P�~[��>�X=�6}��6�����!��\[�:�XK��<�7!*Y�4�����ӧ�o�eF��h�v�g��*n��M̨�f".zM�Keb�Z���To>�f�G�_C���jJX|��H�;�-�<%����>p-<���oFpGg�a�t@�����>s�ɦ�KV
���~���3|��%x���g��$�jK��#�R
��ˎi��{�Dz�I�|�Si�l	l�����U���p�i�M� ��,�S5��IA�y��)��5C��G�Q�1�q^~�I>�sU���^���ک�s�Nj�Ô!s
ͽONa�-z�A�f��C�5��+�9��}Kvrf*)�1î4��Ovud��s�*�Khu�ym�KPކ2�FKk���a���P��x�h��g��(MԭMCv����}W��P��.�T*7B�K�M��	(E�[ З�osT�����h��Ʀ��j�B��*E2|R���&��tu�>mM�\���pI���3=����^>^�_�������{���w��������~�Ղ}����L�N|��,��P�˺�\���p���ۻJ�*����Eބ�	Hַ�k;AwC{s]�^�KW�&�۾��ʽŝ�y�l=2��B�(e�:*#I��P疧i5�@�G�Y���ko/+C����/���|���b�I����y)R�P��]���G�Y���s�	�!:�V*d�w�p(�}���	��^C��*Ca��3�V��]K951I��+�r��h���?k�dK#��4�Ι��,C��ԙ�D@�$�rV-��O%��6띞����亝�/�E2���!�&��x��kp�.ē��n�l	ڵz�Kf�:-�י���+%嶻�t��ʕl�{,�c�C)f�ƅ�%K]�e`�V��ԝV��=�B.�ȼ�L,c�:�wo5�]ړi�����͙�j>{ns+rRX��Q�e�zҀϼ��QYV��x����p���h���I*�F��KM6�a*�x�qS8�v)����[y;>�S(;��)���g7b�-������)�ӫϺn3|����zK�a��Si���,7�kp�K��x�6ȴ�Y����٥�jv�{5Yn��/oB��1<S{g�`i�YI�V�񥎒�v��-KR�e�ۙEr*���{ez>>��RZug���Y�Z���K���7s%�)�2e�Z+\��ʣb��
�e�8���6k��­��j�E�2�� ����t�8��,�o-M���h����%|[�:x�\�,Л��#V�
6�^Mr���5P!]Ęǌ�����2��߷��#�ɦ�O�)l���c)�s����C���c:�9�Q���!o����s��yE\q�i����_*[�L�s{��C�s��� D���Ւ��l�Spo �s`���!M���ޘ�k�hX:'�'��_PMv�|��]�8f��N���dN���cQRI��\k���gs�
c�gnL���C�8á2��ό�����_U�,�.��i����R�c��ze�Rn��p&ϕs�9mbã�=��I���m�'e%�@���A���$�/���(@n��2�،4K�Z�2kw�ieB�R�.�y
�V�y����;�rT���gwΘ�����
� l����F>C.YZB�qxs��:G?)�k5-oW*#.�Dq�M
�8y��ĺ[�^�[Q�<ڥ��&��Ցӻ5��;l
����f�wZsM�Qs�60u�h,5��]J��xe�)�R�p�J̬���1֛��R���09t�ͺ|�oQ� �[����̍�=%���[<]��<��*3���V�Q�h+˝vZ��kf�{�qfW+��s���vɼ�]��9�&D���K�$�d�f�/e�ժҘ�)-+a��
U���#�c!nk9�obyghfN����m��ש�2�i�˖��5�-PǈK�P\٭;�A!�/M^6��)�Ws��h���G(=�Iς���c�Sm�s���t~���(�1��4��[kf$љt���h=�r���1$F�'F�CR�����2i66��C�]$G*�����-PRi
��hhy-���vԕ��AAT�TD�CEVh���ZF�f�Z�A���(�h��h����rurR��H�6rm��	JOw$�KN�P�:ɤ��l�J
))��أM	��4�,M��CICD�!@�=@hhb���@bZBbP��J�$+�CC��D�DAE$HQ+@R=Z�F�	���ih���Z
��)��6��]2�<r��:�T ?��B��t�~��/�	�O/
�a�P�ُ�W��x�]
����w�W�~ɺ���1ن.<{&�qDj������@�$�$Xa#>��F*�&�qG�h����c��8u�ʀ�z���w��{;�_I�Q��<$ >�G�g/�l�4���Ά��f%J`��k�խ�=������/�^�"�d;�w}Qʣ��J�4���ts ��|O�@K��+���Dw`��N7F�5Z��f[���/�ɇ�ʂ���s�Ż�0V{�C

� ��8����i���>�V ��6�c�$xD��� �c�	��|�'�6��s�F&�7,�aro`�Y����/+S�0LU�5��ݡ�Zz�e��������]�3�z��Rͼ�X������6���L�E6�Rܬ2R�gnt�Lu�q�gv�mmT������!�+��L��ʀ}�j�z��x_'d]Z��#�47o�t�5S���Z�u/Z�څ��Κ��z�}LK�9(7Y���m��t�I(k�GG��dp��GsemN�w�7�±�#�dZj�WQp�]��k0��j ���Ȝ�ʱ�0�}1-��U/=�ؖBwt���t���DWCB���>s�Ɉգ�ݹ�W	��Y^�Q����v�r��"��D��5�HV�ʶ�L����$v1�޻�B��,�t��CD3C�h��������By� OZ+v�7���hеc�;�җ=��X�u�H��v�S.a�6�zӥ�O�"d8�������F�����)_7�WR
��IF��$����A�5YI�"c��{І'���ZSΐP�����[�9O�5��9>����~� y�  ��y�a/���x;��yD���U�+��'%��K���K��	���G�B� �I'vMU���v�^�p̖�JϦtYE1.R�oR9cnL�LW?0oO��.�s�A4�d�!�rآ��rѮ�z�?b����k������6[�Ic�&XҌ{�B� ���jQ�P��W6�jR���*Bb���O>��'�U�U�,d������֌�b��	�J:6c�C�t�����A��͢y���ߟ��B�,�6.�%R���7�O�ׯ�%񟂯���!]t^f�^�\����%��^>�0fb�obf59���U��,<p��l�Ǧu�F�־Z��� �K��0ϱ�6ꐴǴ����b���Ůg�cbr��w�Ԕv�p��MѸ��,�N/�F��y�|zMIj������^�fDYL{]����L�-�9��1�3Y6>0H9l�1j�kwn�r4��>"55 ��4��6'��^��<�y3�ɞ���){��y��*�߾�YT�^���+�����z�P^��T��"|j�x�x/zۨ0':�dqd��i�aȲ�v��#��"���k/ca<�&�	�e\���ы\��5,<}#�{XG#NGR�����R�n��������F����ՙ�*渄CH���c5�����j�<D;�tTWI&Yt��,V.��4���GVb�9��KTf�Q�b/y���7�{����  2ku�A�E��߄D����e��ni�؊����6�rXí���SH���lL<wDQeƺߥ��,wa�jD��)�;�dB��a�_Ú��U���T��0�M��ɷѼC�,=����n�zB�>&�V>�xm�.�*@��U�H��7>�*���V,rg"����.����W�����zS�������u�FE�@�6��f��i2��V1��U���V\�D�Ù�t��h�.�%2ݯ�t�mWX�99�|�S�kf	���r����	q6���E�v���`�=n��>�V�`��Jn�[u�c�6�/��a����M�Q��J0������F���.Y3Y2�q�\XsH
)�΢��^���`�:�����-�I��&V󁌄��s\�*��0lFg�::r��&(E{��O0_��`Y�j�5v#�D����;h���R0G��%xZjg�=��0�2gK�\�z Z�},�F1�G^��LA�ء��>�j.t 
�9�Z<tcu�r|nSx�)���!n�{�f�`���6mh�l�b��yKQ�2�Zв�MJ����ݨ	 �mw�f^����!j��*gB^�VU�}���q�B)�D���-k�Ӳ_�V��ʓ\��^�;���g�l3{��C��)���}Y�ݨ_q[cqV*; �K����u�/_d*��
RP��B��q�Lr��tZ[���m`�T[�غ4)�94ٮ�#4K���0���5����p.3�:-ʇ�����G��9f�����]8_0c>�g<��BWW�ۂtG ,�t��~�/5&����z�3��N;��<�9�b�ƈ�L�Μj"�*�t�21��t��z%��[�z��
��c%O�t������!�e �/0Ձf}�ЃV�$V�]��6��o��m��΀�i�ul��-m�p��]�h��2Ƀ�=�ɰ�J�p�,���y���گS�U;��:�P0���@�S����fhX��FY�1�ڭ�<��<p97���li4e+8���Ku�Ŏw��U�����:�ʔzCgS�/D�w�⟹�0���*�\���RRv�Θd��>r�[�ۀ^!�)�ꦟg�1
k@L�}sRP�Z�M^� K&�{�dgJ����H�!�rz�cu�N�W&�Nu�O7�7��o)zN�t��4��<����RuσTR~�-�
m��}t���l�b��0 ���kJ��u�����	�}�"�3c�V��<���&��%���:�Y�rk%Ɉ�Tچ�Mv!���ޫ�v�i�k�6�yo��dU9uE�ܑ�kv�^���(	c�vɧ[g������{�Ωrūor,��
�@G)7��V�Z9�q�]�s�Q�C���
�gN�=A&���w�U�Z�1O��X���y�y���=���?X�bP�U�)����.˾y��v"��*e  ������>f���7i�zmz��T��e�q�����v��J��ZjЮ[���_n��C�b���F�^Q��Gp��!��}A*-��Wa�s�0?���٢ܠ(ܻ<,V/K'k$̲F�Xǹ�����l<�;�ma�N�A�/��xy^�zn�n��g1;�F�1T�O8wy��l���T&��
2Yn3�X�N�C����-nB�,U�}���nk�~��n=K�r��=s�OJ��F�B�Ϟ��5�����p4�(�ٶ���S��I�e�|ū�!hЃej��g���0i�Ȧ�R�
!��5MK�ȵ���\Ւ�c�n�L�m!�H��!ٍk�L:��/V�e_S!�W��x��y}$v�|�M��3��u��5G�tJ-���!����YLy1	���v<7��
��ÆF_�$�^[���]N�Xw�M��T�1��Sm�~uH<p"om�g���;��a�D����^�n~T�)[]:8�7H{�pӆ�o.����`���$�6[��O��$��zzqEu�$�9�X{��uu��Q���t���b ��н��q[����=�{������1�Zև�����������xV���}Q����{Y�{��"	���ǥK9y��22���>O[C����p�������}�̋�x{�7��f��̈�@-"�*� �+^� 4���߉#����%�[]8�VD#6����\��!5|�I�PJg� S�������_8���^�;��<"/�X��y�)��R��gB���R7�.�J��ʍ��h�P�W7f�u���NQz�r9���
hZO�{�w��c3�%�G3��Z�6�y��3�&ND��'�Eb�qw�j^;����m�.�q6嚔cEvCn�wPD�9�0�/:�\��*|���/^�����gT[��d�f�N���.5�[I�]����ێ�v"C$`3@)J�钝�6��/_4vԷ{��-%�&Fؘ�&�QO����"n��	r�0�=E𿧵ؿa�5)�|uR���
��?492�=^%�^����fT�(���m	q	����^E���bypɗ�6��X(��c�	�w�gkR��O<'�\X���l:VpC��;-r��j�B�R��v�O�����yX�4͓'�!<��wk�n��(֯"����p0	�+�;m
d1������o&1De
<?�4�8>����3w���m#V�fް�"7��mo�9��e�^n��>4�X�bo%D��g<�{�,���jtE*%�gNj��+>GK��vWn�E��,	wq���2��'��E��0,��c����lwqG��*�S����Ǟ{��ןF��
ZB������� � L�L䡦kP��Oʔ4��f<�,Cf�N�½���aA��y�l&�4���;�P�Ĩ[5�&�a,R�~��cٰ~��x�O.��#��#ڡ���^�dE�ڙ?�"^vϚ��N�]Í�.���{n��j��`�6�ՠ斐+�#�6�p�a@�ײ��.���	�y�0pw���v{i��x��+e�0`S�]�x�>�{� �*m��$��U8u-���͝��v�c��a'�)hgF��C�-F�]۸B�֍F=����y{��BuLs�u��`չ����{�G��2)W+#<�qO�w��T�J��'+� PUcZPb�5�f�k�<գ�ͅ�b��������Su_����Q0@�~P;5�=ҀP�J�k�,Z�c2�Z\�?p�^�^�*�����2s�ni�^*���Y�.�-��ɢ{15D/jP�V]��d!�g/4f3.��Aى�*���2�nTȹ��m��]c
Fd��^4Ruՙ��J�C�޼۫V��]r��0.z�4Y�"5Q��酥R��%x�B���_�xr�ֶ
/K!�^�]Ė�J�Ȱ@�dՎ��N�6+ܳ��M[�t�2�ZҺͩ�eދ�I�~�<^��y�-��0�H~���!y��K�.FD�x([��ӡ^�%���Mwn�F�E��,��d|�(JC1g���*sj-�&�����U	B�#H $H�	H�
�4��^��߯]}7��u��߻�[�Yi�)�9ȱ��gС�7	�Lfs6zN�>��8��Q`V�i�:���$������xK>�:���E�+�I�ֱ=��oo�l���oW� �j�
쳀0�"�*:�sE���ׇ�]�m��E�ԋ�j�W�Ym�g+xo`2���9w)j���:L�Och×�r�5�(�4�p2P���ç-�k\�q��b1��f&29f��%��}x�l�/�g���Y	ydӷZ�:�}����������އU���~�h�h����k�u�	\�ZŬ�~�<m�{��=#Z�GN'�&}��g�>o�MzN˂t<��PhDu�gh�}�F��ɓi�2��N_K<6�{�N�*�cٹl=��g7�Þ����ٕ��a�7%,g�w!\5;��x!KC�i�QD
ݻ�#3iȴ��s�|P��RǇj�wB������O^�}�P�p������������,�KT3^�饍��N��v�JHm�3������e��&�
gF�3���g��Ɵ[{	�q��mR0�5��18n�bWeVѻ�M���YȮ�;����݊�'��ʙ��o0����%K��*�%�.���t	Mb�şZg�q�\�`�{���%aڠ�픤έ�\����0�n�/	mWItM�dD@�̤�r�ff����xJ��P4�H�!K{�y��E"��]������2O`&���J�S|.m�N#5�2��R����\���r��K0�3���m���B���-�#��"��`y��H�����.a�xy8���w�/B*�"�[������d�ժy���	�=�}&�rDKrm
{�'�2׊8�>j�Oִж���h�q��(�j��-Ն�l�s�h��fůT!o".�c<�3��>�a�_��L�Q�X����z�[͛�<��٣V��d�x�z��A�o�C��4�4��#��汐��:���{�F���.1w�V'�� ��Ie�I�˜W`�<�� K��y��yb��i�u�g9S��VD�8�/-.�/L�V��.�<{�E���z�l<�s�}a��c����KA}W;�f1��;�G�Ȭ>��.+��*a��d��.SJ{,��{|����ݶ��+nf�#�Ӥ{��1�ጞ��򜗿m����EW�i�`����*~���\/~̧��i��?d�,ǁ�71mҠ����:)��V�j�)�d�	��e8�H��0�>aía31�jлg觵����n�|k��g�꧐�=ލ01u�v��|J쳛�����O�P�x�U�(U5X)$�V�6����Tɽyo���ͩ�E�W_.\�Ss絪�H�n��V|j���\��w���bA�7Xn��4g�\��Ձ�d*D�J���(��C|������o3�s]>��qS�Ha� �+�@�Z��ԽZ�y�M���t� �������t��Pn��~1�-�Ip@sL�L6&�gǓ����v<7�U�QVɇy��d^�Ȕ��d5^a^޾�7��'y,5�]��aroc�S�fLk��sN���Yg�NB��9�k�7'T/�2��U'B���-�ǀ���@އ ��'��x_(X����1�y;��Lux�W��FP�'^��c�k���.�/c�zK��)٪-���#�2e�l���]d��P���K҆k����M5$�i�<��}�oO0�c��P׶ -�Km���R!�Àԅ�J��˧(�d";Ъfd��q91�x�MC��Ep����<_�$��U3�kN8;���M�9��M���[p��p�E��A��hb��[ǋ��`L�W6���ӏ+�-���M^s2���S�J����P�9�慒�+�S/V�=��<��q�Fj�ɳ�'���4
�\��7j��|����:��u#t7@�5�1`C�=����^^�w��������z}��w�����{�>>�_�F����q���x^b�:�<��t�H�Om��e����n���%r�j��Y}H�6�����+\�Ef���^H��p������g7K�\r��"̩�p��������}�t��gr���`tP⣉F�=�l���|���6�Q��ŗ|:cN)�[�i"�h71;p�X �}[�����͠��B���BV+X�,<�[�:�UuY؏+g��-����׋^ ykc:w�Zq���g-	�͜����N�n�ɘ�$�^�]M=�S75R�-l�&�8�:�긻\�&[��M�J��O)7�2c���[LtΛ\]��=�J�5�Th<���	Y��:5.���[���.M�(�����pѱ��ҝ��}j�^�w���-�ݮ����� �H-�0X$x��d�e�45J��<�;�o_j�-wT�ة�J�F�%ᮣ����뻄^��v���F�Q�����h��tέ����Yr�h0�kxW}����:�a*�n_pO�p͹y[zN��sqHAI�F�R�n���w�5�W+�
�z��{[)�+�����9�n�v��V���� �q����1\n�[����5ֲ��(�m�u��F��Z�:��9B4�XΓ3+�
L�&u]�6�]ic&�wP�:F���YqF&v�tKL�s��ވ�[#\����ɦ�eo6"v��ƺs� ��s�T.٩R��78�l��g-���|h�����]�31lbƝKJ��j-&%��
4�]sV(��ж�MK��	��ܺ{p�+
˳�k��[ys҉������K�}"�=sw%]�3��l��u�-R��:�K�Ze^�ﱍ}�eL���#�����MO�٥f�]�Z�W�}�9or���A�{��bքĺm�)�r���-�].ܻ�ƦG/��Y�])>��5�Oy[E;v�rhW�Af��������'5 ��n
��I�Z+�wV�vrxP<MS�ޣI �H+K��;�&�����z�kM�
�P=N�ᖸð���}}�ى\�O�,}gr�#(ǝz���*�4�r��i�Y��f�l������R�)�Cj�=O��i]�wK ���&w�K�ű�֯�P�Xl-�������}��)�d�7�m6\vFSO�ܳ
�y��c�Ql��U�+T�.ERrq+r�ݠ��`��W��q�B廂��r�y���^�.�}e-�Ӽ��,� {��U��t���fVkh�3k;y�[r�������{cT�opQHF�@���_l�����г��ĥ`N�8�v���p�v������/w&�F��t�-2�4�5�Ɯtd�oq�8��!����^T�s�c��W��{��δ��;�l4�݊85s�(�(������Ö�=>WP`͠5�fFi\��K�k����m�t�~X�AUJ��R�0h�B�d(X9.�����+�
RЉ@�IM' q{�B�EL�r����(j�	���͆��f
͡����y.��A��i���$����`kBrBrdJj*))j�B&6�[%&$�Z �����rR�N��X�iy	�Bօ���	�:Ӥ�4��m���l��u�ât�hKg��:��_5-1+F��E<��i9)ȣAȤ�)����M}C쯣~V���W��\@Y�����K�ɨ����������iχa���%|��,t�]iXl��P�w�:��~���C�b �� �H��(���JJ�]^}�׋�;�������ܾ�sύ	��L���I�x� ���U)�f'����E�f"�pL��֬輸7d�d3����
,��r�S�њb��~m�y��M8�iO0�WO7.��b �����	���	��s^� ��$��, �62	��#�v�֛+6Zwy���p��[��r��wJ�g���q�N1(-^n�X��#K0ax�5�`k�0yd�;�����Zݹ�j?~����}vE�1[yW���F����{�I�mjb��.���Ćw�p04BaDD��2삷��l�ջl�I�nmJ�sW��9�,q�ew��?��y]4=9P��Dib���$�BW.l�!I�/���z��)[#ؓm���SV��M@?tGmP���-؆�7k�u�d�/.���|��0��d���;�>���E�MUNCխ���܆���� ��_�j+9^H����=a�{y����G�2N1�)pgF�yT�o,;3͆6��xy x� ђ�ZZ��9�:�(�8�m�:4Ȯ��#=(�1��d~�k�F����}���=������;�yK8$T�;k[��윈�X��ܰ�x�/�9��~�&iD�����~Џ`ٙ�r���𻏵[ƙԻ��_�s3�h�+ݑ�~�z��z;:��iz2ݼ��Z�=6)2���5�����¼u�>��9���߽ׯ��؅*I����T�B�� �P7���7��6��XP�����Z(T�_��૕��*��c6Ux�p*&�Cc��85���[
��0�dNf�`B�W��馮�,��D��cz�z�Zf��"�h��MQ����m�B���{�Z�u��FG�Y��XP�)��2˟���k֮�����uF+T��F?���i���G����^͗vʘ	�=c��,쇘ܔ�̾y.�Rڔ���ی7#��WwP3Q×�B:�O3�Ч1��C�JC��r,,c�$���&C�q�\XsJ�x��@�:�]B�.}��w�!n�e�KB��*�\�m�bW���.6!�9E���=Xp���A���$B��E:w%֑��,�v)#NW���I��l��y��ԙ�ݺB*!�m˞Ub1�Еhֵ��\%tֶB�*9� �幺Ĺ��^;���cV�v�bt�!Svp�}4y���P�p7��ef���:.w���#5��f�r7Ha�_+S%�n7YZd�\T�'��sP㾻�05v�r(��n=��c(�w���'q��6�ϯ�_^�{�p��A���W�i���Ѷe��ruM�����/���g$�ʘ:�7�5Q�.b��ϰO�e���9�uZP)�v6�./�|��(�Z��̦v���;>Z�e�T���Ҹ;�:�sw��U�0���e�4�>�Iҽ�d=���u�c��
�F�,�1<�~���ן�}��H�R4�R�-4	2$��J��P��*��ȧ����2R 
E*U���H
����Z���W�^;�!g�ܬ\kss�$x�Z���U-ٝ���L\�U��i�mmN�9�)`�Y$Vט�)xr��q��#�Z��3T"+c�p���zG8����P�c�Qf$����M�DmQM���ڛyG4�`��"�T8Pw��Q	P����O�Y�]�<v���*fگ��f�
,6O)f�U���n�=xsӾ�u�>@�Boh���d�B����:��y]�M���k�,��Pݯ�Y�oK���9ח秅tb���l4��eRd��".����.{����f�]L縘{�is��A�M(�M��9T�~K+Z�f(���3�_���P�,;S���.�%ڣ�d&=���l�}4q���I�>QI���Za�����,�{:湜Wz�按]�běT9�zt�2�����#��l��wP�`�����d��3��S���O�5+�OA�n��5��S
��x/J�8ܜ0�L��v���o;o�3�����0�1�QI�q*���:�35Ц>}�krh���.�^�W�yqA&�y����.��+�U3��U�\��U��5���*Zw^���^�.d���|�ͻJ�h�j��cְ���]�y���;"�K3,��kORCa�QM\�y���-wV�B���
V$m��d�7Χ(,�����-��R���}T>��%%L!T�T�RA4�EBU0A@sܦ���ΥR���y<1i��.���jw�c6���7�^�|F�^�T��0�<��<xnLp��7.��OO;��q��^����שyNU��<�;�j�2e��M)��,��� ������{�f	�>&�����T�$�䭂��~c�\,=�T��#�M�U&x���е��x �I���[(+Mt�"��k{1��b,�WU��`��,WB����2��KT�E�;�ui�6��,��c)'֡�i�k�ѽ2���ny&$
@�ƛ��	u�k�ěC�ơ �I�ȱ;z�v��d+���u��a� ��3�:7��S#��Nw�=�`-�ݯQˬ���A`���Fˑ�z�����D��oٮD�wK����\��b���g}�a�TK���
�/�V�7'R+3ʚ��/U'"��ל�1�ʀ*����uh�s�2�q�/Y-�m�B���������<��X�w�\;MD�z�ƿ0����K���0�����񂺲e�X��wT�\�]Q�KԘf�D%9)�ad��P�]��e�0�G¾�gw��P���/^]��d�u�S��V���շJ�i"�z&Y՗��ܳ�̨�Z*�������s����=�Ӎ~y�}�����~с)��6�ݹI���jü[��Y�K]ϯe�o^0�Ls�3W(Z�n���Ǔ(>�9̗x;�1
W3�D�&�'_������	ij
*�h�KnUl�+�����ؾQ�!�e��Ϻ����vh���!�v���C5�,���a�a<(�2�Y�P�ө��p�(����V9�(�چ/!�uy���l*��x>,�-E9�ǫ�d8��h�B��?L�����z����|�-^P�+j5�]ĳ[���(��MIi�	����On���J�H!��l�Ra��+̢����s�R9c`���t�O$�:�R�[]���އ�A��Y╇�:;�z_=���<��`>�i0&a1N@uOö���b�i�+�#.�O���|��q���[�*�<��1J� te:n�������^:ㅛU�8�{�0f��cS���g����_;m� ؏i�@7�^gJ���;0��Y��t�k�<ԢPr��5�`ġ�\�w_A���Z��ϡ��#f�Hk8�I�� ��H�7pט=m���t�D�=a�s�x��5yA�������Q�nj[F����4Fjc��mG�A�)��U�\��|���ix:=Y;.#uU���X,���p���%yJhzv� ��¾�������'���Ԡ'f�sD��n>���&Z��Яg�%i}W�V�н���-m��R�ט��E���-R=���M�%,唥� !S��H�DX���V��2S�b�
/B�:������}K��v5�pL>���4�	$ Lx��Ϟs�η�{��޽uV�b���<tR��?�Ϸ`�{�OY��1�R�MKd�lX�v��h�յ���.YDpF����!���0�vNϯZY=-�vE�UPE��p楬)���]o:�6�k���$)�������^�+�4��ڠ*�z�RF��Tq_�^���bDA���?E���Q_*��g���\��y�2���Q,_ݳ3�+c�8���R�1�-�.=oӕ�(���&۬��ƾ"B�&ԪD��i��Ѧ�R<B$=�H��e��]���m�лg�����i�X�ܥ���x��G��z�Zf��"�h���M#'EN`:�:M���0���@A���5���ռ�7m���l0ə��T5Y��Pxʭ/�N�0���iXv��v-ì��`�1ǁvWѹG���ܪy��qm!fC�ڎ;ِ��{L�so�H�n-B!�Tu91��M�wSl͎��X�g	.�z���|��I��<uG|�f��83�ɵ�q4\��<lFgS���f�kt��uNVDX�+$�i�WE6:v����V�����Lx���\�R*�m;wJ}y��0p��fN���7�o޼k���_��\SpX�V�K��<�սk���I����w7�)�ynKU�ա�cz�]s�TvI��[�6��ȍ���z�����TL�PD�G�����p~��/�3�0�L�@6i:�X��b�\�r{Q���#��=�4���P����[i���L�Iس1=�#���ϪG*kݩ��7X-m`V%R�r�u#�7X�"�Sx�S[� T�$Fi�]u|.��a�=�/�D9qa�������~��KFZ�3N5Z�Ů]����ͪ�F]�Jzv��lg�#�k�v�e���r0֘���������L�Y������W��/�#�+�wMD;k����`VPS����R�����ar��rU
�,�����=�ۆ��w�:L0A���"�<�i0��?S�x�Ak�QV���8.*�xʭ��R�3V�v��l��H"|Sy�[xǰ�6 "���(.;�:g�Ո����4��N�i��_��6�ll�i�((6��,�U4�n�=zw�LS=�Yg��N��ʡxp0a��9j��5WG&���`�]W�*�'�JfNT'}.CgZ��TZk�8�\ĉw��ex��;g����cʝ�J-�k��#�j�Z�΃&6�Y6�+*�_�<�v^S�}��}[��3K�7՛���,�Y�p�v�ڇ��j̘��[P�NiQ���fVn��it�=T�˾Ȭ��PM<w����@�T�X���Sj��/*��ټ�R�V�8ړ+.�G�s/�fo8�W*��m�n��iW�}����Z�ĺݱ8���d<50c�����K�BY��nM«�m�a[F�G�|��xö���ƙ�_OdJ�s�� �����欗=l���T"����,�<�5���X�A�:��8q�E��V�Ӆ�3�u���P��U���NNI���Pp����Z��؇U3�͋�7:��(f#��v�I+����)>�%@���Gp���a �}M�֗2�sJE�Z�Scm�������+h�;V�n5�Ix���>���C��	$ܻ]�
�s
:�I�g�`����O�4'ŵ"y�%H��q� ��i�9��:���M\�*��]M��qֶ��,�ˤ��夑��������˖i�r�{���.���9�z98i�V�h�u��z[o٘��S�>�5M������R kX
fx�r�Z��q��49�A�ɦy�b�u&�i�x�֥T�~�E?����T����(@ �	f��2�'7��O4��z��s����^���4�
k۷���ӽ��(3e�&�튇�["]�`�a��"�uVH���@�ubi�ҹV����$k�*��F�WJ�V0��;uiux˶��v�z�[�[�ئ�7��DE�^qz��:L;G�dj����ʹ�k��\0ڄ��fa����U���R.�-U���(p��0�O�9]�quI{F�{�e��M����0O8�﹆�Wӿ �hf�S�C]��=����p�l�"�?���A� �f�.M���W�S�&��^�cC��|O�3ҘLL[$�1�����k4��Y�g2�۽RGyl���h�+���^���͇���NsZ�w�^P�uʭ����S;��K�]����^�a�6��n�1��V�3]��K��9��/��J����^�7��=f�e��c�LS	�����Gn��\�-�����l����z�Ni�a,�Ӕ_!�
�8���%��M/���
�)�����:V��F��W(�]�-Y\�e��7��h�Gnx)W���7�J�+-�FQ��c��<��r��8ɨz6z���Jl�W��,���5�k��ߵ�.��,Q��h�fEs��Ii�bUr����e�2Ae�5f�<��2S�e�lK�Q�F�`Rzp�ˋ��<%7P��+
۷T$L�J���pϬT��^ה�y��׆L$��ˆ �㚕Ζ��[�M^UES]ţ��!sg{9���G�#�cj(�J�C��!�p���?Zxðї�۹�2K`�3�]��W�0��+��n�tY_DN�t���P�Ք��Wy�b!�.���B%���P:V��C]���<*���0z��s
jF�Zb����nq�]J��7W�m%kDR�ڥ�8v��+�,Xn��1���͉��`�`���+���S} '?1N;���Q�A_�:Ő@���܈��&`�7�>�X��]����LUY��Z�����Z���α.l�/,��@�`1�xcݴt����ԡ�u�ڔծ���u���N��oR'U�Ĥ�Dzyc�+ϱ�{5HZt�S8��q:vF�y��~m�s��_\K&Yԫ�����9�-�|h��Н�-^1B`m;la�jqPf���1�aǘ	��DY^~�2gץؾ��X{n�S����} �����3V���MA�sM;��r�	����#�����$>�Q'�~���_�Y%=��}q9�� Vl�w�W��m.gڊ+hn��4��|�+���Y��"l��N-�R���k�43���>l8y�|;޷�w�A8�ld��z����X��JmE�E��X�B7Náȭ	��dC*[&*��7h#YPn����h�B
��zs���t�*Y�4����k��"�B�q/\��m!�ċ~蛾����n��{�11����L`� �ȟ�Цڻ��uc9U�;��*͋|YQ��^�/w�����x����w����{}�>�w������`��36E�4u�݆�������[J�mQo�KlZ��C^��:M2����h�g�qƓB�й� �����7aM����{�����.3ϝu;�⋱wN���c�p�Zk+-j��N��=F.T�^ٍ��՝V~BF��k��K";M9�Q�\\͔]	і�^�(�O-uy����lh�bc��t��T���<�'\k);���9���}�zbZ_S�� ��]v�ʸyvS�]��:�C�{)wvJ�m��LȮ��X�-�.�8 m'w�k���Ȑ��K!����oA(֨��:�<�|
���b���}cY]�W�E��M�Z��IJ� ݗ�6+��̦�q��.e���R%:g)�<���L����Z�-EM5��	�"�W��#��1��c̏h�!%�P;��ʎ�־���%ݽ:E]��r�����:��^*{����˽�M�l+(�nR{�s��JK�̓��x�� �I�
��,9 �^k������Xpp�=�\�U�"obXB��`��%#-�5͵R��v�^6/n�;��u�e#��R�-��-o�֎
�R&�œ�FwL�57s9�؊[��m4C;cu��@uf���B�EnEm�9Q��#h�o���k=��Lxe�kw�: �P7���0.��K��"�n�����$�ۥO0@-���r���@��fөC��|C��� ʙ���b�y�iJ�G�a;۬�zt���]i�v.�U��L���6H�(EX�`&�jt��ɝp3�vЬ�X�hd��MKG�lu;��d�\��̛!ܽ]ϫ-�T�i7][��R岨s�f�u���%�I��T��XԒ����!4ӚT�[������X[�lɠީ���`�.{��;f�w��[��ƶ��>�(K0T�W-�r��\;p�b���/��*�P`�V�ֹ�yyx����1�(p��%h!�չZ��t����9!!�L�Z֭��%�.e�O�R:�b�������޻�K�8��&��0�����:��i���թ�	���·�Fd���sǪҹ�l�L��t3����p�R=��t�����SsUQ� ����.���t�z
��]ʘ6ZPmh'V�\ƺ�.�4�nVh�׳+l�HM}�<�\׼N0���*⦦���u�%$C�����h�S�b˵hH4�ȴ͊��#8�12�T���,���u5��P�al�r���-�K��Bu:+���^��X�|�4�;��$7:�Gj;ǃ�W$٣)� �ɽ��q�>�S���Ma������c9M��V�)� ��6��,U%|��n��d�m���Ty�8�3��gt��@�yv�sޚ[Gp}5�W4�3�Ӧ�%Z&u�X��Y.u�]�#�1wYZ�1Ia��X�f�Ў)+�}@7ѴUeN��x �7��s����ȤVd]�M��')$��P����Ӊ4;�4QȈ+O�d.e�YZ�i(v؇UCl�
B��� �J�G'24SF�<�'����gN :ے�g�u>$�&��|s��ɭ���"]�m�5͹4�sU%����`�h�P�TU�y3׮x ��Ui��˛�������m�:���ҺtQՉ+��WQ��œT�5�F4��4�&�.��yi���j�M]z��4�=F��#��<G-�Tu�U��E�F�$��Q�� ��E5Ehy<���ι��s&����GS��TPu�������)�th&�9Պ
Jb:��V��
�����}մ2E٢�� Q��v_N���o����O�J�6RY,ZV�wۢ�p�r#��@
Kʹ ���ɛ XV��ݫ���	<C���>���� �i5E��t�$�:��%2�)~!�M��W�R9^G<��yp�@?;9g����f��v�g�Pj��A�x,'��)��US"�<�m���mQr�}^oY�8�a���,*wf�Û��47.�^��=r=Vv��������&�*�]r�-�7-�ι�VǐJ����'_�L�d��, �`%��P�zoc?E�T����eé��6��[S'�m�yR���E'�m�dy�����?&��M
���\t:]cOj�im���8<���}~䇻���YKo>q�sniz��c�H�zA"�O��3�!e�m��?GQq��,�6�V�DF1�2�Ga���ԪZ�@��pgR��GX�E�`+(m��X�ƀ#����9���l7�C�t&��	yNZ�0`�,%x�//�8�bЧZz<;f�X�|38Ca�ή6Ѹ�V��p�����l�v�B���e����GOH�������c��<e�{�d�U���)��	`k�c�!��Ё8+�:��r����jhv�Za����|���Z����֯Gl��œ�bw�Ǩ`�w�:L0A��',�){�Z~��ܴ����f㦍�f:幫dt�8��W_R�c�C���k?'�ʕ��/�ȹ���҈��[�����1�9�a�Ge)r�U���F��Z���>���TQ��UM��aJ�d����N �K��[ú�,g��t(�;�9�ݞ�zk*�w�>�	����t'�<�A�1�z4b�l;O4�Ŝ������,i��1�ɰ�O�g
����R$9�r����wa]Ny�����zöN?���n�N�J����ԩ�=����ɾڊ�*�.a��^`_*�\N`�XE�q�X�</dCK�m׾,�����O7�U�1{U�CVS�9��F!��ENM�>;�MZ��K���`���ن;��Q�)���y�#���[�:�}���!3t��J��]4]U󫎑]��-x��%�bv&d���N9f"8��M��9ǜ�x:ً��E���,Ӻ�|�\���ou�@�n��^�P��#����j�{j���h-��/01r�v.9��5�/�ٞ�0NVҗ��װTE�&����U�5�����v=�^h�SG�jt�1m���`7���w�n�F�3��@�����O1s�)>�(
�Ų9T
k�rVv��=�ʮ�3��FL3՞s�4<�8;L�"��͗�=M�{;��c[(���p��T��ta�.ζA�,hw]�2�g/'6Z�W!-��L�ʄҟ�(��G�=�pVF��k�")v�����-옞��[��=()[հ�%Y��<�Q��K����r�����yM�-�����Z~:8,���Y�V&}*��zC�A;Ye�È�!95���r�I֬C�gi@ξ�xi�S�}��0��)�eӵ��f�؟�����Brr@��[AQ���r�(,?i��S���hڎ�e��Oiz�6��;0s����������F�0l��Z�\��V�Ś�iGD<���!��1��q�F�4�&5{sL�ZoHa�/xHRYY�{�udj���Sfh��*���J}����/�;�����0�fˊ����eqd�CHosZY`l����W[�����+���U@�ꀣ�U��&�ǧq��w���m����)��W)��S:|]�f��y�u��d�A���w�%墮�V;���:�v���X���,��Zf�1��܄�%�^��WY,k�9�	��/���s<�?�b�����Es��x&��9���g�FN�ۅl����Ov=]�^IA�%�;�>��M8̕G&��B�/.�1˕ ��0�����B�cXdz�{��x�uCE�q}t��А�
��;G���)�a�o���"�	��T�0�(Msf����,sj ����VhJ��L���P�z���o��;��.��U�{aӂ�HĜR�_۟nc���b��w�_�z�{F����y�?վκȳ�=����	A��cX�����9V����,�'r�u޳����hM���H-_��H�mX��B��ۂ�܊��a�ֹ�k&�\��54��m�5�>��=����H�~Z������}*<��Z�f�m��k(���G�����q�N���1��-Ø����� _��C@��j��a�d�XE1��)�nH#���q�{.�l^Md\�X��֮gSI;c���&�*��^�b��[�y�2A�I�R��l�r�����F��Y=�����6���v<p"i��������p�gM�4�z��eqv��
Om�}��4��r�1���q`�㯁�Ƀb���(����C#��8��f$N�w*��W�{˚;���\�K������~�����_\�����`p0蓐tÞ?3��NگL�s켲�t�&�N�����M���>�
z�,0�C�زm�nc�1_C��.�k������!0����b�Y��8����y��<�o2jKj�j�7ZS;�D�W_M��a؍
���,�"��L��޴Ñ��=S*\�^$>�灅���k�6�U�9[��D��4Έ��#щ��b�d��_;'g��⦲J{�#ٙ.��
�\C�&�Ԝ��X��z��+����5��%_p���>��3/�YM�mX�@��m��R��]l�ؖ�s�d�WlK�GR�g*�_Ӝ�A����AU}wd<���F`WذԴ�+�ԇi��[����:{1X��
���MZ�#��eUǪl�H K�<�M�j\£9�����Cg��"d����R����P*j,�lX�m�E�QhWd���ل=-τ�?�La��A�Ĵ���X�Q�v:a��ؖ��=�X�����C�`�f��-u��	�}S4�C8�6��8��yۅ�{{�Zl�U;D{����M1�v/S'}MU��uNT`�;ՊC����27f�Z�Ц۹C'�f�u�omx��}�m6�zQw%�����^�R<�t�L�rZa`>;6�civjqǞ�t�1�f[[Pf�1�Q�(�̃|��:b�F�I����PMײ�T0�	�=r,쇘�Va�G�FC����T�97�u�)��j�M�ĶQ��E��S�m-"�Ro9!�p�jM�[l�ek��k���1�^\UrqniQ�G�q�7�F���j7剢��v����|�Z��D��Y��X�[���^�1,�a޸oP�v�W����A.�9;e�n�#{NP�<)�K=�j��&��h+�5��El�]�0�x��VT�l��E�ݎ�R��uQ��c �iZ����/?	��MO�Fg������ƹ{�P�aw����u�5�k����ݤ�+�6^J�T�����Uέ��f3~?X�3ׯ r)��%*���㏷J��:E�O^�U�L�[ڭ ]n%��ۧ�;���BCs`��L�-����U��/�����>),�'�y�MB^Z}�Ckz���th�8.9��h�"��R��ꅷp�9<ՒVz�y�K����9a�:M`f�1�k��9kL5h������f�0�>*���Y�NO^�>H�����n�-��ATם�e�8!�, N�B�ZѺ���ܨ�3c��9�[\"tn���n˙�^�!2j��ޑ�+�f��1k��v��Ö����'�����hx�z�2��S'f�!nnn[��/c�>��>���,a��5��BB�O[hݩ'Ò�7�������%�w6�i_�:ImCP��N�EJ���[a�A�ԺsD�u�1�#�!m�7�8����3�D7&v�����uй�>Tר^�d�EJfנU����%`��rj��ى�`�8ܾK�t�K�-I+I�Sn���Ԛ�L/75#�Ô*��t6Qj���y��\�t�ʖ��8�Sm�r��Ʃ�xiX_'FD��v�fI��<[�O[���EׇTT\�oJ�As�=C(����|��O[��Q&+y�[��GE�'�I��H���ʗ�<��
�=T�cm/��8���C�y�z
�zm��JבR�ڶ9�Rr5��oV��n�T�?"+f��i��n�&t��Ly|
][
�WIs0�wlG�c�-�hr�-s�?���Ip��)�X񃻝�����y"�b�a�w�pdǹ�KuK_�M�'}j��Z�a�M�[���U�`�.َ��
̲,��b�\�+YyFC'Up3E��v�⨳�>��� �Z[C��$[8�Fg:�T�oo;�z�Dc��	q�A��S�&��iv�ҮZʹ�q����]9T�j����&��>��]ɜ�w��\Y%0: �M��g<4'�t+��1@��0e�v\����0ۺ6�1d�4��eD�[#w���������d�c�:�PX{M�aŚ��=U\�& ��2���C��������>=�=�y���҈E�U�  S0��Ä3���5,����
���]vY"�9їCz����k�����ڬ�R�#�>�,��eW��� 1�;ć���bٿQ˳2�\Ñё�9���6��X���59�8�w�<�+�f˂�"�"k_�x��m�uOi�[�[0��4��gh˱�pE�ٵ��Y�D�	�ou���/�����칾QYkl=�.Nd�i����:K�E`���}�v��������Ix7��kB��7��ZS<hl�r��>x�~X�~Zzz�qNn��ںU����N��Y��Jl�;ܧoۅ��x�t��r⧤�]��9�Xҡ��]���է[M�Q���%�wn��e;�<��vyV�s%&w��/��n�N�\1�;D5����k6����^�$��Ƶ�Ə�߽�A�3��>����0��j���(=�3)����9�˖�R�n�+G+���b�#9��G��I/��J��'����l����m�9��6�����~��ԀP�XZX40V�RRq�{ ��E'ԮD��E��t�l�Gdx*���>ͬg��#J�EHꩣ�/�r��Lu+��w������.|O)��m��*sV,�a޼�mO�>�~,���ɽ给�:�Fm�C#�^	�� �y�h6��[w�7��ٛ�$M�����SOY�+l��N�������K�0�|z����A`3B�أ��:!�S~u��N�������q��[[n��[9R�Ψ�vÃ ǊT�a�o�E����1����*��A�)��tI�g��6c�m���ϴX�"6H&Fc9\1�d,9٬":��O�2��MB��*M+Qa�7_Gmx��gc��M��d�v�d:Vp"�ry���e�}w�{Na6/K�R�ç���8���Z�/��E��kv~�&���b��鴩}\��[?-�ie��Jr�q0��e.V���b��8QrMY<�Sr���<| ͏޿mj:'��b��z��>��R�-�������Otud�wr�������4��
r�}�R]�Y,X&����N��;�d]w'1�O���ي���yw<�\�
�-�"	H��J�_so�#u�f~��c��[�I�cp%&)CO,a�b��R���a�N��dY�a��~)�r���j�Θ؜�K�S&=+s?��ac�kS���zD�����9p�햰����d�v۶��0�)��3��V�fr8�g�����]#m�����&��V��|�w�d�d͚��v���mP��lN��2^��T�^�OKx��f�]��u��d��B�u6�/ �s4�'�X��Y4�v�Pa�/����c��^e��ɍj�2��
T)j��g��m���j���>�ڦ���L��6����Sn��`�v�DV���z�B�f��Ћ�jÀ٨<�C�;�خ�bZ�Y�(�&ҪD��cH��/���j�����lk;Y89��������&�v��j��X��ʙ9�٦]x�ۻ�zcZ���ힽ՗s�A-��b�#I�<�MQr`Hts���;k=n�����c�i�,�n������R���^ZУu�(�̘�x�I�|h��.]��e�X�4;ޡ���=�4(�"!H4&���w=^㗤d�J�*i��\�!}!�hT7�&�y-,:~~�R���*{��:¶�I���3fIG5�q3�Xi.sT]�Ҿg ۼh���呴6TV�ff键�r2�7��Z�V���L&����S�1�]BSɜ�xWp�[N���X"�V1:�u(6��>x1��V%b/~dh����˜�)�=q֬����*���	dR�IJ.�|ӇTq�7�Co?Q�/Ɏ����|���n"k�����e��dq��
�d�^Ȗ��a�oOa1B+��N��u���Y�00^�$��X�=c�c�e�1+��
���Wvd�ʇqv�Z� CԮ����
~nY�LO.|ݵ����뛫����ɀ�v)���Lc�5f��\X{{ȑ,���k��*Y�x�Lu^ٶ���'�^�����!���y&�3S��m��Zc�F8��lڃ�^�}��ι�2G.h���������o]?�۲���E�t��yhg�������e\��I=Q�j��r/�4>!�P4����1�ߏH��f4ǛR�3�DVC!�B=̖s6ٽ���{�̉�����Efö���|�������@# *m8z�t�}�NX����y��G���B�n�]~�t(*�s��
�L���U;��w�-�3�4yűՍ!�{������y�}�^�w����{���o�����������P�&�E��r�z&йA�E
'�I k�P{��6.�Wb@���V�.�{�R�FR�;c�V���27/�
ҩ[+)5�G�ŷѴs/{�+/c�\(#�z�1W}���bK��{k��J+.(��$��J,Wi��(VQ:7�8ؽ�u��;gܰ�clm��f�����V��.���ѓr�F{�#(��|b=���Єv�OB8���,N����9raC�����ڋ�$�wa�a�a\��pS�J�	}��D�0�����]���TT�ܕmwG�%�rG����ef�!�0⺶����`���F�T���ĕ8�_Yr�t��b���,_^sh����ԗ��e��8�]��{�ܬN�m��V�[�OI���f��|�eD/�K�"z%kS5y[[qx8Kp�rzkg-&�^�'
�̾�/�6AsQOGos��i-C�tT�v7�m7}�;5c����r����U��շI����$�t�]S#=+jf���,Te����m����ҽ�G�v:�|:eϕ�ܚ�vޜ����J�$�7��^�����G�^��[V�!�ԛ�	�C��Q���i��J���8#�O�m劾�w]1�9of���qsM���]Zʀ��릻�����Q�����Y {�3#��oA1e�Ѽ�y�Q�˚�l9��N���78��Jcl	E����VV���3;2���V�[7��qʂ�l׵��|��ԛ���C�k�����f��dt�}� �D�u���ͬt�x�h�!�s6A��1��5N�Q7:�.bl����r4R�Y���w�*�@q4'�1*Ȉ�V`%�=�uctQAQ���1�'^N�	Qen$/��eA��)��(�0�v���2�/x���q�)|�.�U��&�t�+�Bb䍞k��3�X��I5�'Y@�Qh)�9hCK�Ph�N��ʌ��nR����e�[�	]]�����e�{��ժh�P�{Xoa*ܱ`۳��puk.�U.KvV�՛�o)iXh:�I�pdߢa*7���F�d�3��:�5�J�iNR�8�q�9��,���w۰_8�kv�$����<��Lu�=�N/�����/��d��B����X�!�봜ǹ#�Zir�7Ul�:N�*�
�xu�2�-]M��6*z��?I���ݲ2�65��{:N���U�_G�p��}��V��F� ��;Rk$�]R�wE�U1�9�˘�_gcrf������^�:Uq5�T�ǋM葨����_'K�緕�k�y��>bU�+y:�FT}Y����a��8oDJ��lb�3�a��e�=�6Y�bp��ܡ��Y���9!v�h(�L(:���k�%%�D'K1�lܑ˴��#���N���8�R)n1`��≢��f�+�!Jh�\�ykEƮ�DT��%�D��U�5E/#��F�.N9���5UCE' ,gw�O6M4i�F*���`4Ҝ��'Pb1�lhj��6�7,��@�SZpb�ع�f��J�"�1Z�s'8��b4������(��b�*[�
�\��UEF�b&�g7Dsg�E,̓�RUUTFKQ8�j��(���2QUQD�<��㭺�b�!����z�F��NZђ&�f��Q͉����;b��v�SRm��#lǨ9r�n�s:��9��SU;f�-��1�Q�K�n�UATb�#\�D�D�ՙ���m��Qբ(��*h���lb)���>7W�Ǭ[�ou��@��[1�-�W+o�7�����X�����w�c�4@�taO3o��� ����9+���U�	�J*��cI�:��a�{&%�6=?tO����� ��d�#\W[�����s��$���ڬ��&�b9����W)c�.5]���0�>º�[�S��-�8�Py�;#6�0��Ƌ�q[��"�_E�����&D��˵C%�H���&^�m����>k�꽞x��T�!
ߓ�t��G�s����FO��*�W+��i�x�&Bz���gJ2#w�+@1ZDw.a�P{2yżI쨶�nY���ۤ�k�ek�t��3,���];;2]��mxܵ7+@^�|fWth�7�ݼ��=�	P%���-��9O
k����<jy��T���	Qn�r�3�a��J/��5�0'�����P�Zh�\�=]%'j7!�e�a痟���9��)0n�����e�|c�\�מ�"���&\��Q�n��ٙI�=)�����
	��D�n�[�y`g��a���>�Klp�J�
U�<VP�kz��RU&~�<Ξ���=��:� �[�7Iw��e��BN��of,����T�_U��gEM�N�f��F�Ųl�K�5���V�6��5P�,R�dky��@�-�w2��ܼ�U�z�ܽ����٨7KF☹4Ժ�J�]��M�^�μBƠ�֋�ޤY-�%[0��η�6�,#��b����"�(��2�Z������[i���Ǽv�����q��x����x�֠	���CāL�|��䣧�7շj.d�$�9%�2�6��ݪ�59�;<�6���0�f��1B`��u�#UK��Cf��ݧҍ��
��L�f3�LUd�c �ק�3u��ߌ;Xn婰��ە�*��VI�9�(�{��y3�ɔ���c�uC\�1�&��!�v8����헽sc9=�]]�
ً�劀~ɂ�����^ȰVD�h���0�X���&�7�&E�A;>�l]?M`XF3��ޫ\����/=������%���J�h�y/J�<"<�즪��Y��b.Omk���S�\��Sl3_��_B��/'�W�놌�6tXh�NQ�$v1�&�@3�Np����&��c��>��fZ���X2'�BY��>�Q�%��_�~��t�����#���N�c�;���8��
Ǔ^�Єs�i��U�K�C��Tx� �����窆3S�ۉ�wql��"�+ke�c븦�#$N�/�^�A��d�����'����N��=+�N~�0�-��y�ǥZ�+��<+5wk�4J�%�ʕ�m�枧y��r)�U���y<ҝ�4�ZT�J�'�g�a��ݐ�Rv�W�>�범r�nG���qk(�˨�\۹YՐ��[��Kr��'��^���vt��U���x*�S*-�I.뛮���)iS"�Hf �Q;���>�{>���m�d��I��I*���0�Xf�^A媹�����W3�)ku�������ۅ`��[�,�c>��A41�1�p�=S�o1(laɪK��M{β��<	K)qVmW0����g�?Z2lh��+Õe3+�zط8�aW�D��`\���Y���ۅ�Vu
�p�T�oO'�j;�bPXpZ�ӭ@�ޑ�O��E�
��4d���P,����$�3���e==E�D�V7<��ǩ��3�@�:m.���	l����O!uG aw�0�7����Ɇ	xN8f�Z��^�Ɓ�[�W䛵y����v��������mLq",�;���מ3�G㢭c����"����׍�ʺCT����ؑ����[4%Tc�]2������d�cɍk�v~z���}�d��˲����l����09�iq���^���_=�6�Ħ�4�f����g�B��{��"!�-8����5)���]P�G�m\@�-Gٍ��/�&S^��%�l9>��!i���d-�QYI��"�-ɗ3�<�\u��eT����0�G��YA �8����\bN�:u�6�Sҟ:�A�A-�x�zj?I��⌝���gʏV�ˡJE�uN�m;�.�;>u�^WI�9-����jplМp�M-��y��Nc1��=�V��N?乞��y ��'a_Z�Ԗ�%�i��d�t�75�"mZ�[h���z��UI�@�ڙy1��Z�Uw7U��O��8��!ٍ�ȏ"�a�6�v����윎��q��xn�S�q�N�nm@�Z,�̰L�og��#7n!�k�:��o��S[@���t���@l�@GD��6��۫��2�wt����^F��;M��C&��6�lt��zTA^ˑT&e�X�6]�7eb�Cijج���[6�ш;�<]��a�`��3M�ֺ�9�T)�M`�&R;�"���Q�7�����m�x��;E��r�q~sJ�<��	�X2=��g�ڍ���9�~v�WlS=^�ؘ� ����$��g����e=���y����8�%ӹ.�����E�4ЛseEɼ�5��(��TA�c	������ÃI:/"�;]th�>��E�r�o,\��M�7h曞(�mWUF���%ȨlL�Ml�EP������t�j�pO��.�y��p�tA�1z⪞�ve%�b��װ�!�D��`�I�#���3q�u���V���C����H �jѼj\�
�<,y�])��ƻ*��dT1͔�e�L�`�+r+(U�QIc�bP�G��[[���l�Le��>~�G/K&��T7ڷE
FH]�AX�����o:6 i��S���Z��u��=���Z���j��R��w��e̙���X6v��VsWs2���~��?����cZ������E�t���h!����`��Ed<����щ�_�/�۝}�GO�����]��f��{R�3�DV9@Se푠\��u(gܲ*����p��i쪍�'�8���H�%M�Pn�;�b.�$�ep���&��X$��P�`v�2��L<*SO�	���P��p�>��l��,V�3F��R�j7���[�K|���;Z$���eٍ&�d�g��i�aӉMz�ze������w��g�hW\�*;�c�=�/e�)�g�RRa�gK��U~*���e1Q���Y�:v�o�UX����1��JZ��&��YT6[z�����(;Ia؀�-��i,�D⛸0:���u�_^h-Di�~�����W�@�����5E'�%�R�ǻ�{F�Y#�����[,�D�d�h�'[�߃+Q�$=�./��ײ�ӓ�����
��K���{�*�e+o=?^H����f�Z3��?�Bn=+ ^�|;fr��\"�4��^Ĭv��z�ޘ��_Q��.��㉶��ϕ⭤������O
D����]�䨯V~��Nz���c.����۷$��B��x����S�)m@:X�Ykv���qnϻ������׆��\J�$�0���;��vm�չĞ;ܸ���j��i�qRr�4�P/���/��'X4"/�u��3av��7ۙ���&��jw1��Vj�lOn�Kl�IL��:�j0�9~9�υٲ�� ��nhv�&GBxUD��{$��y�u�u׎���rk�E�V�X�rY�	yos"�{-��3��t�2te�ȣ�������������{h�>v�"�?��]�+��w�"4����oA��'.3�(c�y9��Y3���H�ƫ]!��UU�\c9j����ii��P�nA-�ME�WTH1�z��h�y�z��vϙڼNH�cN��gXe�k�������]]%�s�f�IЉ��Y��?��h޺p(n]\z�I�ҧI��8���/7\/�cl�zq@<b�A+�3�5��ߞ�dga캪�#�j���=�Y�km�3w�]���\�1� �ޘ �k�=���Zyח�"�	�)�^�ű0�nM�R�%���9J���A�=��`��y$��%	��(�3J�=��G���?[O�G�%�p��ύM��=Gd�!\MV"�>�U�,ĕI�PE�\���݂�ټ���;�	|z�fV�*Wb9Y����гR�z��l�:��f��Ӛݍf��Ŋ��H���0.���[97~��7EC�C��I孺z�qqũ��T�C�o7�F� 
�����D��X�q�:eB�R}���m�a���(�莟�?�cPo�+�7���}�;�5�����՚]�Ռ���cX�˞�@��P�*sUY�\Z�V��lQ����:����C���i��@�i:J�����0O����s�lb�u�l���w��j��>!8�+�l�n�\0�l�p�S+��6e�̰슐CE�٪=�(�E�;5N�˵���w���@Ql��<�����&s&9�L)Pu�¼5�a���ki�т��ss��h�[}��e��t1*L(#R�����;k9�F�.�ǎL�Q��C!��7UP|�yX���D�A��!-\�R|�8;q^�j���(�du�@ �Cj��ɤ|�,Ð��?j���W��Dk�P0�����9X�T�q�b�t�j;�e�����r��������n5O-d2�ÓQ�I� ��U�	����)��WYo_�[C�����\Xm���G�t*�\���-��f�l��3���Jq�o#�{Q����7�c�=��Ѩ�L��������׋em�"�j�n����ʲ�
iqׁ�
�ƵӐ�o̓#��=�k��r��l�u�� ���Ƿ�W��x����!'�o�^m�w3n�!S��]��Z�Ҩ�ι7�9�1m(��z��5���f����V�%��G!'2�+���?�8�*~�
;_�s��RΆǱ0��Gje����6�>23�9��d��u:m�:d/fFi��}���wDh��#Չ����{a�ȉT�qUo�g4�V���m}ܣJZ��{���T��;������.3ZF		M�iFi�?C���-��[�:�I'�3.��'v�"��s<)�R�hq����z�E����n����j=}K���_gws���e�q��n�w8���6��=�����k��PL���;��zyۅ���ES��4ҔV�ꃓI���oT^�Aؙ�sȆE�ǔ�ɯ�Цڇr�O�Wו̌������2sG=\�K3��z��ojG2��W[��I�o�#T_����Gp��nv�ֶ�m����v���Fx�z��ɔݸUS.s��۪���P*3&z�=*	�{(�E�u��������9
T����
Cj	H�����Н0�UJn��E��휗פhF�������0!����#���+K����V@�v��2��sJ�>76_��t��X��)���}�}��Q��%	�m�k�8LI{�����u֒R���&?O}�õ=�z�q�n� ���5�9�u)��Ǐ�q�������zh�bB��U%5ݑ��c"���� P���d��5F�=��(sh*�-oz\��C=sp����M�
��K���Y�jN5���8��8���b	u�H�|�ts�m2�0�^s�����㽦�+�SW�Yn�9X���ſ���E
���qŨ���yfӺ�Cr��CQ0��q)��9��v��1`p�v�L3���tPp��%��g�e?zb��ɷϻ���Zj΃���W�7D"6�Pa�]�k���i��5�F�桧7���m͋���9��u�5#Z�)Z��n��LN㵨�;6�'{,3 N�A�3��6�ã84�F�~�^�l~�2;|\���b�]���/F"X �I�:�:4^]���S�������9�V�>�C��PFN��\D�	U���(h��4�d띷���3��M��<���eö���]��V�Ю�!��!g���]kfR�!_K�=7f��h�vc7t�rk8�{.����>e\���M��J'ہ!�PSs����m6�^�)�_�D��v�%,L�"d׹q~����NΛx�/�L|�}�i3kݔN�k�Ƌ�N֘ԉWU�I���:��ufW+���U��W�콮ŏb �
��X��S�[�()l�T!�D�犻8ⳗ�	�e�w���|���;���v�i;��=+7�ǂ���z���EB�	
�/s�-��w-�Ȉ�Y���,��3hm����A�P�Y6�I�����/b!���A�K��ȗ.�
V�sE��u���AU;�/t�kd*��8�7���|�Si��-�U��B�l���zu[9�&r34K��Ǝ��U�`#�삉��P's4���n�c����Q�N��٥V��w8숩U�b�{N{5z���и?�ː�pҰU����Z0�n�R�w��2�F�Q�n�c"�c�ι-��I�*�|@�bh�ӕ�aΰ� ���]gC�Yj3�����n��=�"��:Z�6�Զ�q����j�6�sy��͸v�|�E>��c�n_D�L�J�Oc*_�Z:��_���VIM���;A�/R��MVƤ'��^��sS����yi�^2M�J��o�:z����\���~u]Da֖�s)~go} ���IZ�V���{e.(�zO#W lc�b]"۬��5U�\cAx43�c�p�Ff� �D��$$:?�~Q�9���3ڬw=�ݡ��2���ax ��~����o����~?������{�/������>Zۄ$�ʣ���}{�qa'[��F[��eG��X��ei���*j9�g0���o*e3ۣU�P��PY�r�U��Q����y�uŔ�^,gQ�h�(��pW/l]����˞��%�����pr��[F0[�}�2�p�j�p�7�$��w�]�+幑m��X+E)�t�v��o#D��.{3�	c�RT�)a�$�&���u�{5^\v�\Q	f��m�%�f�%rN�)8Qxq�Z�]���B�PY����L[ \3$5�,��*�-����C�2u����(�٣B�2�-�QK�殃(Z�����2�e��PHX��s�E	n�a�е���'��ԥ�A8���=� �	V�dr�IHx۾�b��NY�\����13��/�q� |0��F�	��w�D�#�ʈ�������]NLu�kJ�%_�f��C�M�e�:BաKRܬ�y����Z�*��ù���l�ջ+]n1�F�%�L�X���*\��W� W	%pj��Lk8����h�i�x&���{nP#��ƭ�If�H$f�/�m�ٰ�gN�Բ�=FU�Q'CZt�;�[���� q'u̪��p�v�
�bw����n�,��P7��[�nI�.eE�0vͮ��V�}sS�����i��C<�t�� Ϋ�,�l������l��J�q��t��s����I�|��f5Op�E��[�risJ�Nk�,D6����h<�[ڬ)����>V���z�+�����J�F��Ǐs����QY'4�xY�sw��(�c��¨V@�u�`}�"��ޥG����N�b@��Z�)f��c �}i �H���nd�n��a���&��o�s"���ǻhN3ws9:Bur�g>v��Uu�8̀֊�]`e9T�$�R[{A:�K�hf��qr�3����Z�Yg	�Ek;Y��t˩C��LvY:�a��`�i���*GHB�ѹY�tl�p�sFLT�s��x!i��۫0��}C+"﵋ʙ�QբSp�¥m����CH��I�j�9��ֱ���3�U�Ϻ� Pj�j�0УH�Z���M�FM�����qH!�}q�T�̅֗yM6�ol����OKy@ls�1�3Pwna=G��mSu�EL��u�F�gv��V^��ħ.-��(7��ʂ���UNl��B�E��\��bŚvA����u��7���H��C��㮊����,4�eс��;�LRVj����Z��gFe��t��-��V1��̙#ƕd���j�A��Е�C5�B��'����SB��P.�XZ�^�lT��R�m�c5"���i#XBl���<�*Gr����B�/l�3��?���bbO�Md�"A��福2*�{�b�󎱐��;,Sm2,�5*�9�F}-�N�����ѹ�ܵ��cc���ng�|������ ��N&g'1�J&��M$TL��MG��DU0Es�c0�LD33L�UE5RSW6i���1�1QEMT��<��IMM��8�
�"��1��D�T�U4l�	���LEU0Lu�Mx���1I��h�D��j���bH�&�"�(��"4b"�l-4[j!��&��MPML�$�D܍U%-SMDI����F��lub�V�LQUld�֢�
��*��(#N�����2�tS��PT�EU&�\뜎Z:�71��R��4DMM�UHQC'&�`��J&"-e�*H�ۜ�MSM$G,FڣjJS�q8SU&�D�,TD�\ث�h���L@QLAEƍ}Y��͵�sr�]c�u�b�L�Pl���߸HF�ћ�<�'e�ng��.�F���&�^d��U�]��`ܭy�)E1̼�`g�K��,S	��L�H%H�L�L$MS-h��b��l��F���e�O$=��h I$�"*�����e5�(�9���,y1	Z�0�xoE\ca��ɲ�b�ˣbwH��u�����H����̱�$��l�_�x�x�&�Vg�Uj�墕���YF�\���Ob��5�6*��t����`ct*���0ݯD��h��c:�*��v�-���N��(���\K/+�dFf��ߵ�nGx���g�.�]�$����}=�t�l�!p�n��}���K7�N�B���LSakо�C����^���6��9;p&����;��y�/'�Fw�+���;NLC7-��5c%�\��ΙW�:y/�P��
�-��[ŭ3��p��寷�g�DvC#�ײ�!�ċr�4���OW5��)�X��s��7��kz����z�"�^=�\��Ҷ���7Ey,}[�h�9��N��4�`9s�ڮ9��$�C�E�X��'�]�gÔ����ǎږ���Um�EMyPvL��K���q���WBD���m͡�.��y���f�T�s����~��~r�f�&40yx{5�e���X����*W&G��"%��2������g&v�R��[�]�8�%i���)�:��/}��Dq�)��KhGP�Ѯ���J�W*��=lG���s��z��`�XȠ��^����4���"W�����Ǘ3��u�ٝ�f���ތ��i��8W�x�]2橀�x¥M�O���\<�g��^9[�ˊ4�X Q���su�5>����V�N���hz5�92��t5�覸w>�zfs~��vq�Y�U)q��]9�S�Z������Q��ԃZ�*2��^�=�W�����&n@0X�/��B��읢ޯRa�cp%&28d�R�K���]��q���2Œ趂��������5ػ\���x7�&��
�]e���ތA�M��V$ǳc��#T���X�@�g�]��*����.2��P��ӗ0��r[��	i�}�5h0ۡ5 ��#ڡ�=�:O��a��_�+���qL�Z�M��q��˅5���]��̗i���=�3$7Y�%)���t��f�y>�=˸2�n6���;`��1pb7u�:��Ю��t���ь���d��`�9�m�>]��96j"OS��Tṡ�د�n�L�w�C�0;��F�2�G?ߒ_	���v�)P�%%�k&���=��?�~���J��Qu9Y8 ��(��)�{�(H���b�	�Z�g���F�H:8E{Q��\���k��)PqcO`��m����z5�{�6�u���w	X3�j�c��I�r�BX�ٺXE#=O�K{Y��ۤU�V��Hc�],�ee���Z��},^g���;Q<y*�	���>N%Ђ�5\����fǯK��jء�ou�5Uۚ.�h��|���C������k Q��V1Ӝ{�fGM�x�5G)���Be��d�k��dOLPhm�T�i�&�f��"���Y��l1�Hv������[!���r�_l��h���zh�a�T�wg�顒Տ�v]H�_K=�.`c�y�ѥ���:R�佋�5D�!�����*�\>2��*���1I��tsu�k�; K=�����k���ާ�魔��Ii�g�,�z����C�;��noFq�Kt�p˸��i��E�9jR֪7��#3iBai����-�).�ꘆ��)-LwR�n[D)Q�M$g��~͞����)��V�T�h�����^;���b�i�/��X�Pm6s�ПcE��i�M|cK���Zr�*�5O��X��.F�0i-@f�:��i~��wAW����	���ы��%I��]�ca��E��ώ=�\�jk��7,���Y�HV���7m\"�j�;���`�p��
0�NCc��#�����׼���{;"ę�/^��~o�N�H��˟o��+��MGխ3B�
+�`w<%<*�k2.��,�!�Y{��YZ��Ph-��D���2}��!my�b����_�ߘ�b����HV�{b�/6su���x�,r*�7�4�!5�#��#���K�.߹���T���E���R8�h������@r� �}��z�a����N�1���@��p[dq�r'U�S�\��ʍ���?.�<cK�`3�ƴ�~~]F�Pږu�����=�6�W+~�峝W�z�c��mLL�u��
R�5��Ơ�a��싇�@@�v����/Bj=�B���)h�nWOWXs�]a����RY�ụ�T�T�f
S��(�dY���쁖"�S_l�nt�h��i���T3�P1a��}��A�H�Y6_��SjW8լ���B�G%^�WY5i�CH���R
���פs9����漧Z�j�O�L�m��訶�|B���*[ʨ�m�70��X���T"�jX�S��O8n�+����dVVn
�9v4��XxB�Ȭ�����dS�0�	�;Ϥd�"���y������*���	%��݋"�^J�/id��YL���l�)Qm�+���0SIC��^ E���(���y�<-�piJ��uK��q^��>�V+{fq�@�K��?!n��h.9����hN�KKSn����_����^ux��,M�c7��;��Hm�$ ���F�gT�7�]����.��'��I-�#�L��Z��U��$�1*N�qa���� �Pam�*ث˗������!���˗����׼�����_��5����B�K$$��2��?k����1�.}����������՞/9䲥 l�,�d^<v��,�ST��گ�-��ׄ��绣��AҨZ*S8��OV�	���1�zg��v��h�J���w�A^zx����%6!�v�v�I��:hP$Χ�2F�5�t�5U�OR�2�svn�y�'j�t��s@wf�g)ݥ�Ș��2<�)�'lX�n�
h�䉫t�y�)��0(B��9C:�@�v)��y1	R�)�����n*�#��!�nYu�u�zZp�>C�n	�l�j`��� �sܧL��5�pȉ�H��nO/)h�mY�����Ոӵs�Ď1���Ĵc4���3�k�=�/��/e��v��-�݌L�o�Oe�����$̦��N�4�sz*m���l�j�wyFm�H��;�_�M맧�6����,����.��B_e����P^fP��\t���lJ�OU�)��3�U/
��nS��(�3�f�.��xռK�&�ى�H�l�ð�?��c���P�v0�&'� =v��77!Q<�.m���\Y�U�)�.�l�� ���r��s엀�Z���2a�
q�
�&�`��X�� ꦞ�z`�N��h��.w-i\��Q�z��/z�r�p�p^E�5��w�0wWPε�6�w7Ƅ�������5w��
w��u��R�Yێ�����򫌖��<��u�K
�/�зR3䍭�x�-^P�Y9U�|w��@�R���O���[I�DJ��^���i����r���s2��t�M1��	O��K,mɜɊ�i��)p�/S���*L�z�v[s��t�E�C��^jJ曓㚔ݪ0^��-˖K��Ri�&������]a���esi���l����׆<��؞��L��6��YFK"�9�-�mm���!�3lv"����ŰA��t'�N+�Ku�{`{qgJ�N/�65=Y��E��Ё-S���:h|L�n�ݼ-�m n��"ذ8��m>K�)ٽ�or�"�Ol����!n�L��W=�'�J�,��,Fj���F�,�� �6е���P�/��Sˋ3Ym%�V�.nr�E���_��h6c����ΆǱ0��e�gV����ǲ�l�\�3�v�&ǆ	#�W��BW������g�߃����pQȥ���}~��m�>��Ow0\n\{Cv��Q���Z}�M>�:��2�z��S<z��|s6���
�^�m���!�z�^�*Dr;��K[}/BY7
�:�)�_K%,j�<�Y��q9�%c0�8ﻂW��:G�[�|�.�g�-ܩ@��h�u&�+���U�5#��?}��[�ߎ��F���v�������\D���w��)�gGb'J���S���yƽ��Ү6x�5�1h��w�&o֬Woٙ R���^�6���Ч�F%y�&�^�=�"�ns�X��z`�v��!l5<��	3M�q�SꙦ��S
�Jh��g{L���h�Lfs ��R�5�\���c���6gL� G�(�A�5��k�.��SM��D{C���ț��R`�˼ڰJVXJ���T1c�
f[��<� �5�in�ٶj��ŝ8�'c�c�{zR� �[K''�ժ+/Fy�"��h3���yo�kY����~�l<���z/
Ľ=ֳ��,{�/[�f���>DM��5�Z4�_j���i3ަ����ƀc']�08+e<Bx}�G�ߩ�f�S�*�֬C��6=w�vnr��/�˨5�N��+�f��voy��ٝ7�x]&����:]x��5�>z|��g�^�~tP�W��-��|(=ǛG�_sq<��Z�ՁԠWdl���gG_ט����/wo���[m�JP4p���j�wϤ�k-�{�ga�O�8�f%R�\!}23�7�D�˪B�"�<�������"���]��2��)RiK�Iܫ�09tʾө�⫥_�9�u_o1���^��xɿ).��T��u�}.e��R�U ���"fa^U�k�O~� l�e�i1&��r��q��-M>��U���N	g{s�!�i�;��&S�#ݚ��E�@���^���:ם3�;�7O{W.�Ȯ��M�gf/��Ik�>�Z���fbU��ws���:p�x��h�];mc�4wFmQ��X�(�#��l��TY*�=��m�X�qO�Z:���vܦ�NZZ��X\5�\�R�	��w�|�k= n�ө�+&*A[�����3��Y#g�x-�U�@�L��(F�Ї���&�q����6�-�3�u����֑dʫ(�
C
z�T�|���-fC�*6Z�봅w��oeeŽz�*�%(˚�R��6�(���Ms"ջƦ՝z�<��Wj�V��-{ 3�3�Ǭ�O��]��ӊ��U�g����	���U�-��6lĮ!���#�2�V�Uȳ=&����3�`o�}�l�]s�� ���}�;��N���T08�F�Q��
����KJ+�jƨqʙ5G0�E-:����Y�J��߻f-T�X�5���e���Jž�n���*V��D%R�_s��ւ�nn�pw�h&H@&y,���N�a�^H�e���P*�=�讄�#�͐F�45�N��x�����&�cmu���۳>k܅����k�b[���/A��>Ӝ:��a�ةw`Z���u���� :Y>F��N�_]P/�Y�'���Ά�v#	㞒�G:-�����r����hlnC,���x��il]:��Ys1���5�Ǣ�]�ΌH2�����~P����3_���M��f]^��:}��sS�R��}�5\���\��˯wtx�Scƭ�'J�&��j�Y���ט�b30���.d�-���]q��V.��.����;X2�d3�υ���\���t���mj���d�;����ϔ�iŔ!Q�^C�0��d�#/�QB��h�]��N9jz�wwv��$+,KW6x�lF�Q r�S��/��`�d���8����^_�'d��g)�k;��KL�2�95h��6(Y�B�O]I҆�(:��J-
,x++�~4����v��G*�i�`&�b�w�6�T�̬���� �w��s�&�
�NNh���Y�7��[Qt	'}n���@�~�]�ɞ|.�3�o"0���B]L�jmL_���k;����p}�9w6���%��WB������+y�"2A��j�h[a�@�H4(!ݺvcފ'F�=�rj��鉉����#�	7Y/o��s�s�ȼ���k�s}�1b+g��Q檆���-R�
.:=�
�ۥ.;��Wm\5ћ��n'f���<l݁��*�T���u[.�!�,;�ᱷ3ʧ�:CK�x�;�t����*�G+��c9��v�Kf����up�zqq����;8f�8�i�t�B� ��H��nN>t�3�5~����D�;��.d����"ۼ��6��wqn���B�t�b��*fu�mW<);��g�w="ޭ�2���ӣ�j����=Պ�]�h��̘5�Q�w7�٬�G�
�ȇ��b�����H���������x�/w����{�~�_��{|=�G�R�ݱKnӋ�k���j\�&^.ک}yC�\�8r�8o����u�7V/�D�T]�^��-�b[�2
 �İh�k6$���[ѩУ+5��2�e�:�lZ�[(5�BD���dY],m
�2�P�םY��r��y1fKH���uoWJ.��d���5��P�sp*@��RB����u�Wa�j� �h�����
��� �FJ������ZB�a�C#-P�!��;ܳg�3*ՊU%1:����/6�6%L�ysd�M�̽��Ε�QݧA=A��x$�k�V麗�X��v\�W/i�[�]f���tR�錒HK�k2�L]��R���r��TYB�n���u;O�|5[��j\R������+]L'�髗J����e��yN)]�8�2�ВD�n�1]E��n�d��=:#�8�`b(�,�ɀ(����{;]�b�6n=���w��QF�o�;��i&B-i�J_&Ź�Ѝ1�6�A����\k�����U�V�@	$,�}��Z���+����=!�����ck���I,�N���C�ڍ<t��{�m�*�+;X����4P;CsbП<ڋnv,��#�&7��qK8io�;�;��w7\C|�o%��N�R�uu�f|nZ
k��{�\�!�ВFrr�����nDPU��w����p7E��C|���8f����5k;�J��e.�&�Ђ��������ɳaz��]�>��ݢ6������ʾ�Uͣc�b4Gj�ļ�5N�Y��]�ӟ�{#�k=&������΢�#��g���*sƎ�l����-:��rg�u���)u�M����WnM#�Y�зu\Ļ�E�B�A^�?L���"��BO#������^��7�Fϩ�)$�nM�`s��ۣ�V�����
c	�������ZbNO6�;���M0/��.^(��U�':ET���ST��p�y 2�S������.���^f}�u9_�ܰ>.{Ǐ&�C���u#T�̢B}�R�Z���k������@ �G+2� ���{a�}F�Nҵ>�Z�v��+,c�$�oZ�n��TJ^V+o�|uwm9���%w��뒯12�p�0�Av�km%[c�]��)�yۤl[h���Y�3j�+��Q|�-Z/&�a��ڝҼ���'[�(�fTV��6��ꓖ�Y$L�]ӏ��\�7efX}�F�x�x�`t1�2�F�͝(^"��í��K�����6�X����.h2��;8�JX����y��y�L���2��|�kE�x�}-GA��Ɗ[|M�t;�h6����W����bsN�"P��R�IήCՊ�`�"
1bw�&T���O��vV�zCtA�ë<5l���wzXդ��T�F5���ga�{���F��L��o�2O8�7��S9&yKY�-����'I=�җ�Á�Ѹ4�ɉ��pgTw������e9����܊E�߿��%��)j�(�"�h)�*:�L�E&ڶ�E���Mu�*�(h)"Z����j����'�4ܳ�^1���
B���i��h��*�Jh�������LEPUAEESCD�QMTMS1T4�D�Q�TPD<�I�t4[���i����#N*��h�hѢ� ��	�)��т!�"J����)�4x�Es:͹�Zt�EAQ����QM������4�N�������DEE1R�TD\Ơ�J�h&���*���D�8�b����*�������E�v��EF�6�4E���

�Ѧ������iѠ�m�	���Z4ն��(�X��� ��h�Z�
� ��-.������hi"*��$UGI����� �&! ����.X�����4h > ����+U�$��Y��_J��׽Xn��]��3��GMM����yW)(�KK=H[7�¬�$���˨��C��9�h���u��V�1��t��� 94�0WO[.��+���e�����,ߌe�;''�� �q��n,1']F��,�c�D1쳝��r_��u�$rqX��ǭ��v��r�Gk�6��WR��L�dZ�!�3��vGf�k�og	h�m0�5�8��:�d�bE]ɺ�R�%�|�At!_L^��sӸw�uܝ"�3�W��u�9�7�	�hb`d��S)��u|��̧��bADB:��b�n��>�b���㎖���t�3��� R�:��2��	��lm5p��e.R����a�����/v9K\7����t��v���H�V_K��]�h�y�4c��6��VeW�c��檀����i�C81k(I�m"n�T�f�&�pU��%+h�Fig�,ɯ>[�7��*� Bx��X�7�1��X�6�_k�����h�=ǰ�tfřNrv�보�\i�׻���.�K�"y*��\�ٻ(���ۨ��x/o9�F�$!J�ʹ.F�v�A�̵Dvvt�θz�5��I+��EX�v 
gE�B�i�J�\�/���b��Ş�2����M5��u�;����g�KM�Y"��.���)�\?�~M�,���6��WR=�~MA��@���H�. ��=5�6�Z�%��CK�mӤ�V�qv���ZhfI�5�:�8��g#9�����ܛFjK�T�ޝ��g�������������:�ѼvH��uw�!sO�����N�6���$_���l����Sf��!��VKm�x��pz��q��K�;�7c�����6x=޽�h���k�)�=�r����U��~}�-�s�nW�����~ń�p���9�@`���p��*�)�.��'9��>���j�TA�"�ǻ{y�w��i���E�W��N�ι/����,3t���B�͟8�h�xs=1Ȫ��;2 �8�c�������G�z��,)^ޥ,i��
�j=�8W�rb�:'jb�{f4胋ԿUߋ�"핵��hj���ֈ\�l��n��.�1p_�Ox�y7�yT����j��98q���k)f�mL�V1=��O�pػ�cFL<����i��Z��,�pQ�&�]�zD�"��%�Ļ�]��[�sx&�c�����$m��T.���mE/Xd�2^����{]$�S�0G)8��B=���D����S2�4�G?�>	2��z�Hٙ���{��"��NP�ʾ�z:Er�S�)d����k2��%Ơ^�J�a21�ؖ�;�wǿ8�{�TLb+(^�UjV׊��)eV[V�F�Y�n�����[�3��M����H\`ZޗΕ��dђk�k
o\^��i�L������*���Mw��/��̗�L3�Ý,i�kv0���r�ٜ8��]��W�'v��}�69z�=�xo;\Mv�{�j�>���)[����ו��Q w_K>2[pF�S�ܢ�hWm����=Z���}�'���j�s�H(�q��d�뭄�.�fk��-gw)Ϣ�3#p_)�va3B�) ��6���0.��~t诿tͧ��E�!e]�*b�LBF:���]Θ�����tu{#����-���nT[ؖul9:l��\��io�����Ƭ�����]�zsuELp��J�T3'|��/��op�.>[�Y�}K-�
�Q�y̚]�l�����m$eBm�m��� ��s�ȣ��TYm_m��-s������7ܚS��}_ynUf�q�a-���>Z��(1=>��hd��ƀ�u�N�B�ۼ�W�US{-�)۶�fOm?w�0���8U�+��ڻzW7�/���|���������L^,��P�V�M�y��0�I�2�`%�磆&�h2U?
�Ř�*��Y[Z�,'�2e�S������e���ܢpf���Ay�Č����x���@�[g�#��Y*�z��m�t)����n�)��^L^+�8W�f:x�쨤.{e���H<�+U�K�X�y��_a���iӓ.3��!���@n4֦�t��лIm�dR9O8h��Q}�n�����_u�]ye=��gb9�8���ұ]��ݾ�׌���u"��_K:���WW���Ui�[-��q�q��ֈ�'D��'��7mfmL�h�.`�=���[Y>�W<��}
N�j���W���,s_O�y�#d�nq:���������г,��M����6��57����>��S�>]ӎ�"��8��e�b�FCm�0�vӍY����$���� R�DKV�3ۿv�
l)p�dvdV'rJ�ʓjJR�:	#���;+^sK����!�5�Z��y����V~4�g�AT�ݿ���r����
�TI�y�of��;���Ur�x��Z�Z���P&�W�R��~��%+�4�������=o���_DK���f�v@�.�oX�PZxg�zV��D�/*�Y�㹌���<��~ġ^�#C�X�����WX���F����h��SL-�n�3�R��7�P�K^�v$V4�3a�8m��oH}P"�9�ə�,���E��i���m�/t�lǗ��Y�f�6Fhj4T�ɇW�n�ug���WH~̝�*���Z�F�'0o憎��\�����s-.�|��}0�Ũ�;#��k���{pr���{�vIk���i��K�3�9�y�Co;�G'!O�_Fn�N���o
yyOOm�M��!U�ý�0��e0��e��N��L�0�W��z��18 ����09*��l�BKZ���X�T�k�-��B�l[ܧ 6b�Y;-oe=6�B��y�������N�ι��a��}�&*�n��*��N��i����w'|�+t�rQ[ ��N�`����R���69&��}�Rˮ�u?_S:-Y�9�n [�^?+k�Ra�#��-��&�AR�>d�z5���N��s׊9)\�iu�x,�}���C����[ain��2��՗����!�ޭ�q>�AH�	��
̪��(-[S禦,�o6��������5��Q�/{<lt%���d����EfB0N����I���Q��̸�@>h�q˻.+�u��v�lrV
��a*��.���}���Vs��>�w��m��?��Ej��lQ����mw�i������R'�%�Bx=����2!�9`S�N!�l.��;�xW�2�*�#JV����ƛڏb�#7�#p.���F������G�"��"�jŝ��)��L�<v�����x,
�Z�Sf��p˳�C�����u�0e��f��a��U3���|Up7�^7�>s۶h�r��?�ZH�^'��o�%�k;:��+�u$�a�E��Y�[��4/栫Y����6I��s(�R��*�zgw��P���V�����`m�&-gj*JU�t�dV��U���9)F�ɛ�^Eַ�[��7�e1��Eu�r��amu!Ֆ�(��oz���U�o�4P��;�q��rb��1E�rKݟ0x	�U:��Y>����kh�"(�ex��[a��t�U�q;�w�����[�����O�	p��1�S��Ll�EK���]�[�ni�]���'��zm��H'ǣr*��ݸp�V(�єv*��7t��7t���q��E�ֻZ�����<W%��Y�ݭ�e칳��Sf-J^GD�FN���f�i���e,�����C#S�v͊���1*�UW�_�v�{����2J��T�Q�x�k7;qa�Y�D$�*�.��:"�R�=\��]�Q7ͪ��+h���U�yTdg|�^�N�>[�aTN��e��۝��y����.�j�놝}�FHtQ
��ئ|ڝ���	 ���V�U���H�q��&V�B1����ˇ";ʠ�$�5�+5
UXO�Y�4�����5�Z����(�W�?�Ʀ�gZU3"���`���v.���	��"��\��o0T�k���o}~��(3�~�/��mbι#���oh.�o�������#}5��xH��,�kh�Ź���7����m�q�[w�>^ۊ�w-z��)],{i���0��"?�JLM���6�M7|���V��\m[]��#Ζ�yΑ�~[�^cy�YP�M�����@��*U�0��ؔ�q��~�5�It����)�<���g/g1L��cQɻ��>��E��9�L�J
�'�:���1����8�_�is9@=���_Z*}��Onf��EeZ�E�P��E�Tj�e(^3�0�g�W�ؠ>������*:8��W�y�I��3�Q��+����.-m1��$�P�Ca�8U�w�!���L-Z�up1�ou����fM�'�Zn%^�FCg�~���UC�z��.m/�Iu�)׿	U)K�O�M�����,?a�Ӱ�U��aK=��Jڌ�>��~��!O�韛hfw6��t�� ��4�m�lyɉF�-���n�獀6��Muׅ��{���r#$�G�����Wq�B�&�aZY�O�9��m@v���@gCh.o���W\E����2�`�\���p�i��]&���D�� ��jjh)�䷢6OR��uڔ7�e&��L ��2�a����Ųf*�+z⌈��ŷ��˹���[~��\���?���U����e���UMm$�۬�.��/���q�Ǹ������W�� �*���X�Ј^��+��J�(Ks��ݦd���^C#�1J�Ui7�
��=�C�ę��扴���"����Q��8�NǞ��{\���6��E*���4�45�O�[���*�&`%R�U�ꎘ�ְ�&o��h��G��
�{k��%ҍf'2]3Kż4��7&KN<@�v|�Z��/TKH�H��a����u�%�5�㈛��5�q��L��Lj{��g��Z��ݲ��ۺ�p�-`nY|���Z >j�����uOn�3>ܽ�s=���F����:��tq�Yd�Z�d3c����%�91�$�-/1�5�z�����>��U��v�H�H�-����	<���W��1�D�FM��&�vؾ\���*'a�K��g��>�+όec���:o|��6��uk�jQ�S �*U��{��׵�I����y2�X��d�h�&�cd�8��4����)�pX�^t-c��t��<^�[R/y۶�����gǜ�N�x=_��}r.L{`�}�o��Ok�3M����ln�.��g-��c�`�O}�����ω�v�7]ߵ�>KOv�F�,&�,�^�n:f2��Y� ��[�"���^��̽��F���U�ѐ�r�	�UY�D�Fgvž9Mm���EdvlB�2�wL�zk_����}��,�I�7�1����H�-K3@=L�����4g%�!���WR�gn.�=�P�}ZE�2+�/ ���Y[~�^�|�x��fXgD �0��\���qQ�&5�l)�%xTZ�Pr��R2ԝ�,��]�ƺ�&ih�h�o���w6���Z�� ���C�q�oJZ�Jӑ�K�(�v�"$�.^ҭQt�0t?�
�{���
�p�5.��U��woK�d�
�����}�����8�H�}�L��_�@�f�E�3�8H�����}^�X��{���w�����}��/7�����5ЭP��k+.����Z�k�3�=���RY�.��L�Ӑ���Md���&]�{�aQ ���c���.�1����K3��#�<��:�d@0%R��e����vQd6���\��]*r�^��-J1U�VhIٚt<�*Ιdu�ONhV�O&�ĐkW[im��r�h��c��j˺�HCt�^�e$u�n"��3��-w:`}5dqlF
�M��d��٤��.�������[E/0���E�W��[�R1�7o8�D�v#�O�V�4�ەldW��|"S8�k��F�m9����L�Й9�1̧"���V΅�&�u;��ޘ��ݐ�K��G�,��:Wm)�ձ�{4�/����Qr����խ�J�;H���n��]c���-&�屾G)@(�.��e������̧x�<�����Ճ��
�/��H��8�k�M�O�q毅�t�}uuv6�OyN��'%`6�*Ű�sWU�O��h�شi��,s
=K4aٙwE��-X����_��� Ӿ]�<u�]�������.#��ͦ']�I�I�d��h�sK�,"li�����j=���5ysF��� `Y+vݚb=�X�q�ϻ��^��P5�$Lg>s"�Vt�v�8sa�UҊ)"ы�,擆�L8�k�
S"�G0̭S�e���n��+�\�S�`�c����U���S۝��w$:���VN���X7��-hj��Ιb�r�F�l�D-��n�j���pn�������u�<��VA�t�L��������r�f3*p� :�QZ�>	�t��ċ���g��R݅����3.VL��
�T�.��8��/:�g*!ֹ#����@����ٛ�5c[}&�|1�J�쒥2ɫLmd�2:��v��v�q-=�
�^�-��eu�ଯ��G����N�.�ш�-������gy��!Es�q!|k���;uqI�bs��������N��B�S�Dw:۶L���B�ݙdݤIiP��ܨ�
�]�ۣ�8V*8�q�C�G:�:�e]g,�P[��(M�;��rci*��Ȯ��������R�S����*Vzy䖹��q}�%�B��{�󗈞b��!�Y�v��x�g^ZƧ}���zYx1�hJٽѤ�7�D(�f9XH�Z�����Р���6��X��1�i>e	cgV���=�g�ux�,��2�����
fU�0��K-9o6˲n 1�{�t���z芃����K�e�6c�`��6�%���˓��$��4�	��ȐxR�]:֯b�뚓�N��r��#�+T�K{[��H;���,+���fe��WJgl]�wf�0����=!'	X�>mKz4\�	�݋pD��_T�7;#�;���V�4��96ۛ����V믶�EE5EIUMQA5QKASPDRD14�%r�E557X��15MDUPTLTPTESCHETC1P��SP��L�/;Q1=lQlhM�5%MUSCKri`�������*R��"(����(* �l�Q)EQF�CL4QMAM)T5EU%�T1H�T�)MUR�-L�U�Uu�IP�+�CDT$MU�7X4��DRMT�4ڊb`��(��&��X��bb�����tTDDT1IE4\Ú�h�I�
J"�Z�iX�(b%��)i���Z(�h>K�j��Pu
�(��d�"�H�j��������72�A��X�Ġ�ݟlQ�τ���RLإ��]�a��fX���[��U�%:���v�Pqݑ�ǖ��mMe�����}x	����+Ih�j��RQ`��B�4Uɠl��-��}_U6�:��FM���ը �4	���
A6��6�
7>����>?,���z�5���u�i�V���p�P:�]�3����C5)U�)	���⯨fpہa�}�Q٩�`��i�s�6���@�_L���#�iB�Wr��V��:�6|�/���{���T��s[��7R�nt3��F�`�@7�f�5q��ũ��E6-��3�O�K��@1&c�ȹQ��hs�ܲz����d��m��u����Ƣh>�b�v�^5�ԧ�/�a��`vG��^���:��r���X<�,���v�N�gHq�ɝ������V��o*�m5���|'�j�=�r�=���{	��R���Ϧ;Z�Ƽ�	w*���p׃v��d�u3ʢ
~ov���SA\�z�N��k��cW"��8K��(=5sO���Y3ڹ�ؘ���+3�6`V�/F�I�1S_���>�^�����PA��:�[�ԧ�'U�OU=�r�>tpͲ�U�����W)m*�+s���C��꿎We�b�Q+e��TD�{m�vK�؝�X�N�(N�������	��W�]-f:�M�ލ�2dC��Ÿu���z�8�s�c�u������קz(�HԲ|ըfHJ���]܍����t-���b_X�;�����v���5��!r��y)tǳ�k�1��Y�M�����V�W8�y��}���-r!!��2h��C�qgBY@ޤ�/�=cq�{�v�8x�\�F��,ȓ�R��S\�!nf����#��.M�v�>��pM��I*�Զ--�ՙ��U��xqn[(��;#yp���4v��9/\lV�h��ޕ�ؤ���s����m1��2Q��m�lA�� 0��4�G�q�m*��b<n�҉&��a���k�N��-����8�/�F(#z�3�:��7r+lb�Lo���xV��#�ō�l�ۮH�X��>�f�{Ey���k%G�8��r��LӔ+p�J��m��>�VZ��3;Ɵ��y�;h恁O�w{=S����s��&�Z��Q���`gOH��!(Y��
��=�oO�'��
A'e
\��|"���to�ޅ y�.��d�t�BX��鉇[Z5ݞ�s��:�MD�ۧ�ml�ӪG��c�
���j�QE�L�2��\��U�P�-�%ܛ�:�y��cr_诀�z|]fi�m�6`і2�0���d���Up$5'���AGN��� o�͋��Y�ø�v��FL��N�(m.�f�����.�5n3��q�d6s�o'�'O�*E�q���Cx���;A�j�{3�"n"�Q��T;s��k�'��'��M��x�%�QY��gM�ẖ�u�V���wp�t�n#�s��oC��8�W3���5���!�('�NI��jtJ�g���j�˛���M��NF���͵�]�צNrK�J�^�����Z����-2�H�8bZ���O���Dwf���v;��_{��{Ae䚭��[I��͸��F�=����W5���i�}v@�|�Q�n��D���$zi��Y��ܷ}ݜ�٪��9�S��ΑڂZ�%�n�T	�U�����i�mׇ�.]�1X��S�`إs�b�b�]�Xu�z��8(7�k����SY��0��Wi���	��3�X�'^�X���9K��[��D뿒�i�n�9h�2d�ł�rzqڼ�Mv�+�J��ÐutT�dԮqC��ϔ����y���]\hZ!�����d-��/,v'h�V_�dϭ\�=/���+[z�Ek��;ѩ�RVwH[{>:���y�t��yܮ���|�d��M�w�I��mv
�@��P��,Yv��Ֆ+Z[l���o0[�ry�3K�w��i���6���[;����K��Q�NN��5��0��Z���wy��l-���L�ԑ��a�Ţr�2�l����&�q�j�����A�a���ͤ;e6EfY��u�kB��t�:�]��?�⸟|s�*!���>SBms񜊤i]D`7|�a�5'���.�3<E�_N���)�dH��D-�E9�y�w8P#�Zj�@��x^���wƧ��U@X�O�b2RǢf�#gX�]��<��*f=,�e��x��C�-�g��|*�*�F�j��ʥ��Vl�Ad�)\oK�{�J�)�^$/?�׮^�&b�b�]�\>��$Gq��-f?�MŐ��/hV���囼\9���fQ�Go�S1��<�yU�V����_�RO���H^w�5C�)ֹ��^����>6k��lj�҅Ҡ�jJK7.��+˛��X�M�4���,�C�fpkd��i��k;Q�ي��W�ݵ� U�=珵�GLQ�EH��KB�䓴�תWr
iA(N.�uS�A/��3��'�E\ݰXYf��C��DjhF�a��,
�3Km)[K'�9�]3�w&��.��OݽT���T<�XVȋ�뀦�v|���f�Pq���5�U�o3D�k'�ד�w��;���ɭW�˙�x�te�N��y�6Gv���K�wH)d�"�V�wk3�`p�]i�����&^Ok<��F�� �(y�T��>\�W�G{r|���hn5K�E�;cGrU��W�u�w�
�]�`V�ש�U��nS����7���+�s��&�j,�9H���M���Vv7��ף;�k��*#�\K�!�������$�# GY��R�w���z	�~�n�Z�-��R���v���2����p�컦;ڞ}a�vcs�}�N�5�*Y�W_C��d5���;;劐�%���~(�/���U�X�}rM��L9E+��kON<>nU�X՛ޒ���̵��P����}��jEN�^��VO"�E^��i�h.�Lg-׫6���.X1�wq��x��b5���CD}���q���M �S��e�hu]1ȩH� b� ���*�*u�|��n;d�[�����z9�Z�J�l�9V�'JO���ڣ�.j��c�je������7r_��h(��!d�l��i����"�����vf?��w�G���I�jOw�.��z	��t�Tɣ�n�e�g��//�+�Ĝ�o�^��x�=�P嚻�oP(�ԭ�U�e�y0|���V\����NM�;�e��`�zǟ��B���:�=S-N";�Gp�xc�#L��^�� �>�uo����c���
j�"�-^SE�Q{�{9��z����J��Ye�9WFV�o�f�{�|��S]�;h���fĵf���(�w$�{�wl��m���KeufGZ���J��Qe�1e�4o5�[���ق9O�zE�3F�)ޕ�ؤ��F��l��%���p�FP��U�4㗺ld����Fkz�����C��ӳzuoD.�KO1�e���K��NmA�(�69�/�vB�vQ�'U�)<�{����Y:�[�i5\�;��v�ȕ�VP�Qؘ����&U܍�隍�&S�X�j�xE!����� �b�^e�������W�r�x�*i���l)�����l���t���REw�g�n/���e�/a�?6��D�������ö溭�s�3�wȬ�u�ߏsX��W���GˏM�'��M����03hv+�Gb5��[:���p�6�up���2p�'VP��\��̓����Z��;0�,�<'r*.��ӓ�� 9J�M ���tӼ�ӎh��c�~w1�O{���i���y����)B:�`%B���dwn�_����j�F�G*u��<�mǈ�7yv7��=5��}p8>�ϢmH��40c��l��9��Z��J�?C���#x�����M�����k
h��z�]�fp$V�"eN,�	=4d����aPٻ��� v���']���އ2�����U���9T3��QFi�M�57XqU-�~���9��~C1^�;�q�/�O�M�C���F��|j�i(���MV�.�;r��-�KQ���iv�Ϙ�l^��T^���zYu��9{_,.m1M+��Z$Ζ���P�M�.k�mY�[�tZ�{����'@�cc���ֆ����� ؖ���;)�d��j���u��j�J��q��.��f�-��c��E��r���\�)<��ӻ	g����M*��w
��?T�Ù���ѓG!�z!�LN�a;�A�Y��G���U#=�d�b�-��1�^�nC{��f�ح�� mHj�D��E�%�n�D�+I��%Pwظ�=�	Ω����$�������w�wY>�[�2u�0�OO��B4��C-���x�YD�y��,��,�lk-2?G��p�l��:�썵���e��۴�M,c<wm$yX�n�Ո�S/0�7=��x�k:�7�ߛj�E��|+���/s�Bc�s{�m�RM����R�v�@�i�;�T��+Y�EW�c�����n���A�/�؝�0h��>i��5���)�d8�T�>�p��_F��n����>sp���}�߯�dw��B�t�)RQ����L[�l)�]+pv�[|*�8f�;tt�Zb̧ͽS�}J�D��|�}R�1ۣW7�T	S*��;fuuvjȵ�,��#��{F�]l��w5����-[��"�����)�9Vnݩqt�ݍ��5���3ܞ�6�� �."����yU���x�|ݖȻ�9�*pe&���by:���r��T�֣��� q���,��<���Њ�f����1��o�5�s�\a4���P)�B�3@=L���!�!���������4@aX�v���x��>��}vi�q��u�'�K$*��v޼r��5S6�4-e(�=�3�stVߨ�Ur{b��uB��R��	��
̦��"wD��3,�`��¨����a�D���� ^{��aՕ�n��X�#�Eq��i����@�V��|�e�)j�`JyJQ����7G���V/����0�-G���ũUr7�2(�g�S7�+U3_`�Z��XU�7B��&VY��CT.������6�6���8��u�L����pT�@5�ɡ��ؖ��!��@�m2f�E��/ի�Y��ޜ�^�د>�}��mZ�&nG	+.�Z�����mw������Н� ��r����;�@������O��yV�_���ˌ2M�T8�R��z)bȒP�.�%q���+�ZE�t���r\��In"���Ǵ�m(WCO��@�I><�fE�mx��Gv����"����L���qN��Ӗ������ݻ8z�&��4E�MT�ﰲK �Ԩ	�WH��nJ�7G)rw`s����I�1�}�[�# ������-3��/�j�;�֬���8��`�qްf�Ϋ��frt�~����y�t�#��	L�Ůtq~�|�swy��n�j�z���Ɏѕ6��
q@��lF|0���Hs��dXWs�#���k����
���ЮV�L[Y&������G- X/?I�m��^еٙ~���S��4�H*١d�KY��T��=�7E>��W s�e�LôE�a9f���U����i�1X�K����Tld�5J�cC��d������d=u]ztǪ&1%�z�R����J,�y��LNCo3sZME�1�l�[Tڥ���j?	����<�^�w�����{|���w����{}��/W�����=�E�1ᑢ��ﲚ����yL��	N)���ڧTFPD�r�o\r[�6:y���f��l�KO;9ȟ<�ś�b4b�x��)$�VƷO{ȝ�j=�Zx.�M�Շszȗ@�vL�|֊%2��林y��'D�5��++���t�)RԤ�*�fi;N�lW0V���������c�7;96��_-�+���%Jwy�㓲Պy�%��R�y�D�t��)���V�s��*��5�k+��짎�d�m�B�I�ÕW�����%W���_���`)\���\�Bٯ��ޖ��W��V]���(d��%�n'R�5ө۶3e�F@V®^w+Rئ6.��t�yu���l!�4���xi���s��m�F�)r���/�*���8��tǍ��{�\�]��G���ާ�+����[+WF����MZU�Vu3vA�#�#�V�u�Q��|�w`'����3i�a-{�K4�#�T�.�Dˈ�;�&hζ�W��r.����z2֭��5r��vԬ��A4�R��[9�Z�T��K�ǆ��/i���k��e�^���W��Y�k�[
 �V��@c����cWR�R�))S͘�S�v{���r���k}eq�}W{}0*Mg\/����̻$��6o��pEv ��+'�I�J`��e�ał��w�"��ͻ'y_e]��gu�0T�����Lv!PJ��$�� �a��\��5��ɮ���+9G��z�>��9���׵�P���,�ߢqv�e�[��͚ڜ�ۡ�:#�]�N����-�a�z�<̬���6�n�b��cv#\!��G���w�|fP�T���if���4�ge����巜ɵW
�ϳ�Z;�W���범�ݙyQ����\r�]J�R8�ܫ�b8�ܔ�K6��c�9IG+�/vU�a��B���n�.��(�T޹�N��2�G���Zy��$��V�.���v·�*�
΢�b�r�cg=����*2�3
�w������˹�u�Y�Z�Xd�P�a�z�r}2�$��!Rp�����yf'94�H�:�]�.��B��g��]3m*V�$^�k�̮��1aǤ�;���MJ5���* ƌh�W��*��)��M�K�ѯ���ە�ٴ��XǏ��Z�a*�r�3��j��;N�'��x	�b�y��}�J�q�;�WP
��4�Eⓝ���&K�r���9*�
�n��%��VXM\%5�[+�m��qbi�q�֜ѧm8��vo�ؼ9�9F���S�"�f�����p�!�J�W���Of��Z�+ȵ�����#i姴Y��L���r@�+ufWq��@�Q��L�N�5#4okiD���v��WΤ�+� �����:g!�J�	��`�4^ l�A4��.s�����N^�{5����7����<eG�G0j꛳4����s��|�Ţ��������j�����(������
!J
"j���H��(��i��)���(�����()�� ��(:��<�
H����=G	��^A��*��.� �u2QY�BP%%P�5AUIT�4�p����"Z9�V�)(h+F��N���]SKKII�QH�4�4MP�ּ�"�����gM4S�i"(i�Mi�*���*ZB��������"K���))h�f���rSM-��4��
s`J	������))i����N�M:JZ())+��ii��0RkM��e�"R�(J
>�|>�"��{��֪�V͵�F�>���}M�ι맃�5�u��ʉ����.E�� �����aT%���i��1����c�a�q�wC�~�h�Go��; �5^+*�l�q��m� ��SK�������XpH��!$xs�z�ys�ʹimr��vE�'Tˌ�j����������%_����JV�V�Ybq�O+i��ܧ|��/F8��`e1�d#T�o�VM���C�q��W>�$F���g]2N{��2�X��k��5rb�s����c�iU5�(�N�/f�Gh;�~L�`�������T88e�"���J��73M�=�M��b����(������= �Sd��l���b�Dv�>`��*�wڛr�Ke�:�:K-UGqЃ<i�{�`8��o3�F]p�i
˼d�:y��NѻG�OG�v	�얏oa4 і2�ý�sW��麢���ٹS�Ԇ�a\R��M؅
&F��8�Z����^�!t�M���.�qA�^Nb�r�O��s��ҥ����M�^�q�\�96^y��`���^��$"����c�v�;͖<�r��:JR>ˢ�S�<g"��wv����/�ڶD�,�}�9�%ף[J� j��y�b��W����_�v�G��0��-�!�����l�7�`��i��<��Sln;��/�I}憦�A�/i��m26�=�15�W7�0�#1�3p���m����#h����]M �Yc�R�jc�ـSe��k����|r��.�dy���-�|-hp�q��ܲ9��8�U�4�Y&\����I+P�E��J������6o&U�N��	�ڴ�ٗ<��:`9B���8d=l���+~)r��������k͸x���UaW+}�:����	l�!�����Hߘ��F{:�v�܌����]��k���T�׵�Eo� ��H�Ⱦ�O\a�w�����aĘP�R�nk��������'k	��iL,�C|�qT�%��_^E-�C���h��N�T������:��]j;�ml��°3����>>+:�}�a{F�S1P:��|h�8��� �2^L8����U���0�/~[Fu�T��yJ��vqU%$x����cC�������T�;���1�&a#��Kk��t��Wo�,�l�1e��2e��*��TΜFRy:���a��V�]����}\���U��`�=}^�/)����D43�t�!?\,]TJ$R�28�����A6l��46�B�g''�1ˋlZ/�xeK�.��\�VdgZ��P�ز7��C2�'C�4��a5V����k	iZ�+�y~V��_N�ӿ��0a��r�0����D�V���4"5���}4s��}�0��|�_ۃ��i��I�6'�b����ݾ��b
�u)�=��|ݖ�Xf,�.z'�Ǻ���A���
�-ٳ�����M�2��6�zc���wX�Pa�S�6�*zy��m���2d��x�Č]��:��5�n@����r���f]��\�C�z!6�َ��g��'%,Үr/�.��Ek�������A�ga|7S#Mq4<�����z�m�
��@�Z���ta�jl�U��g�ZٴJ���j���SRF���zR���zk�	��s�'o�j.�o�1+�,n��g��	��T�ӎ��Ֆ���/J���;��֭;E�g���0�JZ��I]IN����y�7��ڿ�w}��F*���3m�FRVkm,	��9��/�b�kR���)��eS����׽߼_^fq�nf/���Z�5IW�4	��uK��gN�B�h��:�Y^-|���J�u�Y4�;���N�x�SC��R;T�V�2�����첔ƀ�F�ܸ���.�)g:/���P�V/��zA��������`]��֧wx��r�'�4:2�qW�34k�Ƚ�r����wݪ��V��#��^G�7l��mtOYP��VC�u�9��9���l�h�Aj��n��Ԏ�}��j�oI߿OL>�Z�j�&��|�����0��⼣�*rQjh٭�7�Ϡ2M�9:�!�ڽ�ڬ~0-�G�ݛ��ۨ:�����u�X�5�!Zl����f?���@b|��Ƹ�i�ص��mu��p�=:��<�Z6g�����a��=�+�6�U����5ߖ���Ԍ�B>�9�ý���H�4�v^�� ��'�z�f�`�-��粦�]���O?Z�%��9&�nEh�!���i���fOطaT]��%-����sA����#���T�5�����)�nL6�@��>ڜ���X�x������z,������O��j���/�^�^'�Ĺ�����ƹ`s�TW� ��m�m1R&�U}��xb9���z<�ԩ�,7R*� �F���:��e.���s_��\�ET{{��m3��g2+��UC�UƜ�D�$�k�v���ה���02�$-J�)em��R祝@��t4ʟr��Մ�����]d뺅�8C�7[��2rʜ*�IX���3�d�]�3�F$9�^˺�8sL�C�ěM��[�,�{�Me[\� ���|>��q��y,��2r����bZާ�R�2��a-�]y�|ֻ�;�szv*�p�j�=�f]�ϲ�i�z����oB��S�5��6�8�������Ka)�ˍnC��7�<�V$w1vk�V/\�Den��t(0���c<����GI��<56#����9���y�3=�?�r����K
g/���HP\�)+��2�
j�u+��[�T��iZ�tHU+���̼��j��2=J��JYe�)[\ږ��
�2ܫ���X�nk�"�^�m�늞EL��ח�,�#I�z���+��cYs?�bK�8汛���b*t<��>\�6�s)�n�= �Sd��X��W-��y�w\l\q~����q{�r`�r����5�jMT������u��5Z�n"���8�$��NS!�X2Qm�v��|�������ս�hFѐ^C������ݵ�/�5��9��5��&Ԉ�
�����5I�b��X�v�,��-I�:/(�Ti5m��y��cdO��pD�-5��;�_y_=U�'Gm�/��5� �z��ccSj������+�����1FT)�Y��:�fi�� �Z��<�4t5�@�Tמ�K�0r�[u�-�{ӂ����e��y�#�	��*�����^j����⛈�4������}H:��5�ddt
���4���.��U�U�t�=�lP��l�7"�J�+�4w{�q(�	�i�uh�����%�R�+k3��b��kdђ�F�۳*W]J�h���z�3��P�d{*h�)DܘBc��i=Á�}�A�C���-�i�h��w5!	/�q��s�Ϩ"�y@]]������殥M����#��9i�g-���ޛ���k���W:S~����a\Z��d��Ǥb.�6����g�������ϰ�ɂ�}d=��j<9ʘ�����I��k����]�����A��Tzk�]�蠺}i��Z�^V��zD�8q����ټ���<�J��-��mT.v��9 ����u}x1��`B��̴�	�2��y��e���WrV��l�x����Y�Ukpe1�v+�1n��"3�,��v
OU�Ӻ����-�=6��m�ݔ��b1�)n��9�9^�#���t��Ve�_Wv~^��%���l�1��%��scB�����������\w�xt�iק��\�:C�O+���=DP����/6�A���e����q�B.lϠt��Zr�p����'��7w���o����4��ƌ����v����ȼXd��l0w�ֱR�zQ��"M�XĆ"�Ď�_�w���I�"޷Y��N�C���+:bl4k�z���K�ė�ۛ(l^�����q�{���U][��궶0��B��3i�7�\�U�F7͋gD�m����F�}x�x�]�m$#�W9�j�>�������7��(+��\XԭC�A��:�[�IPaVg���ww��͹xE���g�b�Cy
����?�H�l'T�y9��t�ܸŧ�/���n�܏��Z�+�O �v�����iz���S1[M�I�+H;Tg����v�%y�J�����WܝU��҃�8&[��m8/��"�VeP���P[T:��}MrzXd>�BWvlP�yp�,�<$üV^�� ��V��xʤ3��S�Kd_��8&-m�N.��x�h�n�i�	EJ��$�h]�t�X�t�9LY�[�'�}�:��<M�t�P�E�,Q�� �|�;�4�����u�h�Q?S��Ⱥ�:9��uͫ�z�n�79C��w�F���e�W۬��P�`u�YWy͹�,��/��~R"�Ll�UV�zʅ�wZ�y�7��D�vs����^��C�6��s�@��J���F�w%k�멬��	�6�X76��?c�X������kmS����lQ7ӐGJ=D���hQ�j��8Zv �sp���M�~��+:�s��Z-Q�Mu7�_��Ɇ�䢫O"�9��:�6�w;��Lᜯ_d�·�����8�y��j�U��ؤ�2~�{/D�Ƚ����������'���,�ycǺ�9PT����wm�w��Wt�C�����N1茱�a�{��]��HoU`��{�#?:�����ϱ�.��?}�>Zw%�F`v;dNYj�yB��n3�⥯O>���!-X1n������9�\E 7������Z�X"U�yCN�I>`�)S���0�'��Π,�fC�(��!dmA,k��:�N���q�NQ@9��N��j��������nݪ�f��2e8
�{�5�3�e,�"�1rv�HF�ɖ�d�۱S/SwBt�n��륟%�MiD`���������P�+R���8Z�x�˧�wjt4�T9Ĥ��[;����	����q�d�-�&�eVQY�@�x�����Ѹ-�$'xL�9�ޑ|���@�"z�9��++��&:U�ܷao��y����E߫�|�n�@�՛}9�N�,��XXbq����]��]d�ӑ���w�M���s4���S��2&!u��.޳ �������F,�d]YR�e�ZݶI��1�ت8�#���Xr�s�|�ⷻJ�]�Fav���f�8F$�9���������e������\���MpԳ[IF��ݰ�hl{p���N|�so�q�6�Q#��l�Kg̵�]�r�|!�s�^���Cs&c;̙w@��Զ�v*��EA���C��}�m�SYZuNk���`÷�N������۽��~�)�#�^�T-�v���u��٪�%����uI/��\��̺���$v0m��o���#8�v�卹BcGg;VD,����˼�ִc_���E�aN��O�z����;��-i{�8!ߕ�0�v����4�Ttx����)�p܍��/q�U�:�֍��Vv85`������6˅�B�Z3�u��{,͕�U:��D5ճ���A57-ʝW�L�����Љ«=ݱ�d?:79��7X:vCC�F���_6X���>��+�sǏ~~�����~���@]���/�}?���IV�P�*���1���<ϓ��"�V`Y�	�f�`Y�fE�Fd`Y�fE�e�fE�V`YdY�f�FaY�f�`Y	e�fU�eY�fQ�_,!�B�`Y�fU�aY�fA�VB�`Y�fE�dY�f�dY�f &�FdY�fU�F`B &Q�dY�fU�eY�fU�|OfE�`Y�fP&Q�dY�a֘dY�fU�aY�f�VdXy�Ҋs��x�0�ʳ"�2���"̣2,:� s8�@�� !�P�(1!�A �D �E �U �A@�X�D@��T@�@P�@� �Q � � �UVUV̪�@UXe a `@dUa� !�U��p 0��� ª�( C*� ��2��ʪ�� � � ª� C  L�̋2���0,ȳ̫2�ȳ"̣2��#2����0,���*�!̋0,���"�0��� ����0c��@�U
D f��c������Ś��������35~��f���1o������O�n�� *������܂�
��l* *����0�����G�� *������ހ�[����=��0�=������o�� *,!H)J"�*J)(P��"�K �H@����*����� �
�
H �  H0���( J���*���( L��R
���*�P�? Ň�~zEDQ�A(T(�K�>��_����(>���J|���n���
�ۃ���������W����yc�����~�������O�?_���Op� ��"�
��Ň�A�}�PW�?!琔_ @g����|������	�x�ރ�tB�����O��~�PW��!�(_������~z�?@;	?����r� ���O��B���������_�#���?L��w�?��v�>�%�x |������ɀ?xt���ޗ��;_�ET���_ ����������֟�b��L��,�߳ � ���fO� ĉw|�R�"T��UP���������TI)!%
���J�"��J�(TJ�T��J�I)U�H$��)D>�*J�$R��Z�ET����R��%U$��B�R�*�T��PB��Ei�TH*-dU  
�D	BB�)@�
@BUB�RTUP$�(�UJ�E$���*�
�
���Q*�R�!P��5D���UR�����  �Ҫ�,6�S
���ҭZj�[-�-�6UU� iJ���T��-j�i�fJTͦ�m�Y@Q���4m�@l��W�.�6jR�E�  a�P�B�
.�nQ"�-�Ci;�
(hhPP�n��AB�
C�mmFʄ����lia��B���%�m)B�hm%����e��5V�*ԡR(�J���RP�'  �څ����i�*�����U���ڴ[j�f�V�a���5l[U���h[45���[MHY�Z����Z�Tkl55�*�*60�"�� w[`��Zm�6�Uc@٦�6�
�[V[55��ZE��[R�h��b�Bc���j�B�Pj �� �
��P�
�UA� %v��a�����Uh�C)����ک���+P�Vi�U�6�6�(�-����T�� BETJ�J��  -8����`QZ�`Hh2ق��3)�UT�*kY��F�IJ�P��I@J��hd�5U�R�6��PQ��USL�   6��[B�hUZ��m�[k i�E�j���m2� l� P f��  �l�J��U*�U5�p  ��  @٪ �  )�(�  6�`  kh� PV� d`  MS  Z��45UA*R!T�%p   p  ��  & �b0  kL j0  �5� 
  �Ԁ���� ���UU ���"�   �@�Y`@6*  5�  � P��cU� �C  �0 �h&  �P 8)���J&@ �{FRR� 4 ���x���  ���R�  ����@j��` !���H�2�P  �J-yWaL1st(��<�	 V!,͘�a���x}�\�b���>���W�W�j����;��{[j���U������[j����km�M��klڶ���T��?�G,����{��;�(հ��sՔ�c2�e��إ�q�n�Y�������L�Rmm@!�vw2�V!�0��5 �x$Ȗ�-ܻ����m�����ڽ��z�`��uf�(�Z�m,F���X�@�P���@`��W���Yq���`wwԙ��ǔnQ97U-O~�ݧ�
�������L��[�[d��9%^V԰΋k(0�;lt%�el7�g#Y�K(�7�a,c;���/��6󱌴�Ô�73�b�����	�j@�;�wv�ĩ��Gv]�m�Y�k
v�Gu�Բ�%U3Q�؄:m��ki���*m��"� �d�mQ�B���;�⭠�f�Wm�!^=�YrM�]j|b#^å��~�Sb��יo=WQV�� �w�"��赍���Í|0�^*���4����RV�li���&�8]�dܖ!ݨ�8�F晤D�5�@�p�ˣP�m�:n��(�_�֖�c�ϓ;�e�M�l��\4��ͫݎ�X*�+���,fu.�l)*��%Jd��0���Ѷ%�vʫ'w[2�Z�]�e�E�%ܻ��b�m+*��Ċ��.��Mz-�{�	�jU�R��CSF�#m,R�C��A�����sfP6�q^l��`��ӹ��`�G�naGY@�F�����E��n�l�QR�g�vGwq�[[-��B��w�[��Z�#� ����`v4M�⽚,bt.۠�JVð:e
�3/�Ub�n��u�N�6����͢/v��ؾU1�lT�*K�u��[}�,��kD��f��P"�fV[�c�@cV�e�,�tK @Uk����-��[��P��	QE�\O�7"d��cq<�E�o40����0�PeJR����f����eƎK*��
�F��E�lB�[�ňєC��tq� J�"�)�a�Ӹ@�h�b��r�Gj��&��yv�X%Az�F<�c49�˷8�Z��7vR	���KZ�9��\�u{�N:�7�bm��7T���x��.�(#4̚�����;�Ό�1$^Djk�Ii�%J�&-Ϩ�B�4Ъ��z�R���ǆބ�`MGgUh���n��kN]Ǌ-7�),)hזi��6�f��+5X{��/f���i˻�;J^��[[o&�4����k��K&����YR/��I"��D�ƍ�P��A����8)��n�a�7L�� ��U���j��[�BÇ&S�ɮ���V��43�2ҷ�j�#B7�uj02���H% 7]�I��	�c�PmS����[O1�[�R��g2���\�f� @��)l��(�h�*�4�0ٳp�H�	R\v���׈�a3��f+Š��5Ө%�tsѕ��2�� �@�[����
F�)�'�)ܪW�=į��c.�ۻl�	m"p���R�ڵf�rf�jHk7Z9���=	�QˣAX(��l��uDG���ٳl�#۱p�"�ٱ����!'w!X�tv	Pl�'ʙAXʛ��U�.�M���[,�3a{�꭬�'VGCs1��Y:���r��LP;-�Vk�?�j��šA�h�!yH�5���8�e��M��Va�74�K�jcl����l�"˥bTY0��9�ڥW��2`u*�n�4�����HؘYLTN��LY6�[�r��e!X��)��@Б�eQEQ�oi�T�I���Y��^Zfө���(�r���mM�6]��B��*E��9W(�0�����b��iU�m��@m%sN}����`�����f)����RՌ����Ym��HA���я7	��i��B����e뻫����dK�Z�O��=��o� {�4��{`�'���B��
=��`�m�Lz�z7y)���������jR���Snr�٤���`��1Z2���2��c"#[�/5�j}T�Mn��'P�Yr��-�?
��Z�1N�k�:�Y
Ief��4Z��pf�L��M��;��Ѣ�`]$xx�4��rd6�XT�EX�QN��^�E(\p#>�X0VǗ�rdt�\�%��l�A�1;�lAB��GPe���/At��];.�m<����n��O[va����wL.�a�&������WZ��,��R�*�&݀��0b���@��N���MqGSrk
�po�0���)އ�0b�&�4)�mHi�N�Oj�t ��q`��SS�K�36]m]=Ӓ���јsm�'o�'4ܨƐba�Ab+QH��v,9���II-���@f]�.?�a>���g�����-�U �	S�7B��Mb��Ԁ���ǂ]c"=���ǘ��<E�l��2�kkN����紾���
8�vX���y�|�`pMإ0P�d"�0H�,<<�j���^t�3G�v�Fr -��Tqժ����F�d�Չf�����0���v^#2�kZ�d7~iX��HWV��'7 @oU���ҫ&�-d�.]�UvUEvV�BL[��%���(aɻ*�����۠y���d"���4]�,ʽx�s7-V�ַ�JIowC�<���L�S�[�@����F�X@Ӧ=@J� ���	D)e��^��[/�Z��VI��F�%,G~�>�b�&��4�!�VU�,FXxu�=1�6R�����T���Ӗl��fIO[��{Z�P&�ej�N�7&(�K#Q;�u�Q���w���r�|��t�T�j����xZ���;j��wbBU���M���*���'Q.��-W��[�����i  ���҄�K[I�`TMOuL�2��Z��.X/D� �V�:�^�ՊV�{�����gM��d7���MBYP:;C!��
��Y�0��R-�h�����zsQ!��B���aJ�a8���@@YgR�Mv�,G2R�)SM��#/j�jrnm�����P{O)�	���eA1J��Zx�]��
�h�ٷHƊ����t�E��ǀ,�j�6�ye�d���R���\�5�R�����cVXA�yN�iF,Y[e�SB��U7S�(�vm�`�Xf�5����ˁ1a�����Q�/�q��$l�����˔�,����2ʕy05�z�C���.�D&���ø�Ta8`����.���w-iJU��ԯu�0B����CP�C��ӡ��#hw�)k��h�WXB:V�t)���@��c�����ۄ�����š��Aݸ�ˬX��J'�f"�!%*�D4��40S�I�tK�v��X�M��U�ڵ
��n�*���+r�!ch�{�KB�D��PV��b����n��I�\�DY�t����V줮�=7##N���l�W6��r�d7+5V�/\�����HC��S�a ���P��͆lW�wI:zp*ф	RVc2�᫉)������إ�p�4����h91�f�v�.SU���0�I�R�<ڙ36����r�77r������/b&$*J{�]b{��̡Ws3��q� �y5%Nm�����֕��fV�snZ�31�+��X�%2�r�F��[�iM����0�5��;�E!�b9�d���-ʴ.��+�o#g1��ꤲ���\�9I�6�&(��Y��}2�)i���u�&��xYa��1c:K������6.0oXX�2ܧ��7@+01���ՕZszԢ�+mBxHF�HLD�sD[���U�֛8��6ki*� �!1�,�!��2�6e�U������t
�xn�]�3.���Gh0�%3��E����|�%n���B�&$�,31�@�h�zUѿ������p����ø��ѷ�]:��7�=j�U���WZl"o�֋snݚW)K&ՍQ"�б�4�֠J��/E3f��@۔X��+8p=����Awf�r�C%����Y��3%&��:U,g\�DYP6άz�ŗ�bר2�3MM��
���{���o1�Xi��2@4l�Z7_�5 ��ŮF�
`�%��6TweZ�l�Khi�E3�ẖ��ۚt�LKn�lʕ�,�"̘&�wsJ�p�Q�N%�t;wM�PX��D5�jk&h��M�&����&�%���S�7wC )�P[z���%^V1��jۆ�Xť�%`[�� u���{HY&L�� �bȰL��W2�i;SZU��en�+�����)�˙Bd��(}������d�W�ohڵ��f<HR���t2	Y�/p���\�Yemj���)in��ڲS.V�B����5�w����$!"֛��I� wt5�ስ+X���e�XMFU�xI�*�w`I#QD�*�@���ՋRˢM���E�tY��Յ>)��:*�Ь�o�^䂍J9����T¬wV@{L��ג�c�+gQ=���\�vd8��|��h-Z��,Jueґdu#Щiw#.���M�(Z��O@z�)�&�)�TP�Z5c�&���J�n�f��*=rwgP��YJ
���ٕ�uz��k/pQ��2(�C%er��"%rh�q8��j��0	evw7�8>���JAX�N���,�qe����"e��۷�mĔd�r�غn��&fT�$EY!v�Zr������Q��v�&�X2��ӆB=�O纵���ɩ�'�öy�M��Z�j;j��ڏ5i!�͵�ݡ��V�n̈́�$M�N5 ;��s�lޫz�_W^��}"�i8�ek+)�'2`��$*�fe��OkP���/)���(
/z�t�	�F�W���5��Sa|�P�a-M%Z,���FC���
����t2�(*��8☛�_N��3`�/ ��w7���E+�Iѽ�Gm᧗J9��T����i(d
U�@�	oo䰳q0c)7��ϱ&j͉�2nB(=�Y�ܧKs��,�Q�q��Z��%�m&�]ԨV-�d��z�� ��+,�L[�}���u�nݝ����1]6�*X3a˪Fat��S�t��7Mϛ;�AJõ#Y��K���Ɯ���E�v�ckC��Hj��k���"'wX�+4Vh����:Gԩ�A.�dI��3FGP�CF,�Y�	�:o*� ٭b��,,�M�ӻ@<�c���l��{�ӻdAR��$�b0�@��2��4Pf���ɻ�.c	m��h�T��e�ЛN9c��DP�;��+4�-�%)`3GEQ�("VSī1MДVj]�w�J7�v�6p雮�JoN�慗2�+m:��	u�J;��BPȡ���`�������r^�ŭL9[,f#ʐXV%CpN�~��Ԍ�R(���vi^�Ӂn�wb�
	�	�vۼ��h�*�G��j�j���q���f �� ���!a��V��7��75�Oy��i�/L[,k:ш��+��i���*�&Lˀ��u�¼l)61�0�]̆�e�V�i��4b2]�LL֔�jLc6�&���� ��N���qQ۽��^ԁ�
�����]껓^�Ǜ*��,�Y[�����CFn���x��ۡ�c�*��i+Ǫ�Ɯn*�E�<�se�Fcܳ�nL�lIKm,.ҿ� �c9�T�DG�%4�c{�]l|E9,��ZF\4�A-�SR�r�)�yC@ku��+�z���^Rc�X�Z�j,�q�֫Ve�� ��j�e*D ��Z�uՊ���x q�֩�<��$�7t򵋛 �� ��[s)�u09��h)�ʃ�VX�-�:ȅ�%3.(b��:
���`75�_8yuo*�azB����T�"�`��х( �S%�í�Nmf��eKMAk�v�Z�r���I&����sR���D62 �6���f�4n�[��7h�i9z�il;�{�S��>n��(:Ī�'�9E2�ҬCH�VQ�c�62�C��ōqkݳ.�qbͣ�ض��Ɔ��*�rΏ:T�Փbݹ��8��rd̟b�&�nb�I����	(Y��Pj��^�)ajP�F;6(Ֆw�'cu�ҕy0����J]HI�ⶕ��SK��4Ka�P�7t�iIY�Q|&�/U՘q��zCz򂂝�f���V�y�PIBcFT�����Q[p��"��B������S�X1k�C�Uݘ��3%��ވ�/�;Qf���.�ru%�x\�Xl�3o.��2V��ƢJ�uM����T���
j���a�H�^�r��6*Kڕ���I5���1�F��b���T6�;��������U{���Ou�UY��ڰ�ڍ^F������c������si�busl��A=��-���ݛ�4f�)j�`�<6�&����@*�!m��b�X*�.�̭%8�2Y`�$Fd��[ю8�V����QR4��\˖�Y�tQU2�j*T�k�
5������b� �zJ�;3L���
��M���ɕ�A-o.�%6�S]<d	-�yy���)좷mZ�+EJ6YD�M����]�TB�����$qOl)�s\��K-\�e�N���+qR�[�lx&P!ɑv��,SJef�NJ����9��+&�j���ʖ*k�V��e9,IO2*��-S���i
zH��Y�+4��0�+Sׅ��j-%xF
���Y�Aع[������G x�]�ܹ�(�`ؔ�VT�&�J��	ݽ�b�h4��]^ֺN^�dO�	�x��+L
9A`���X�u�*���wQԺH*ְt]��d����Tݧ���ۥ�͍�C���ۙ$��e�%�1��0<vD�N�}br+Ŵk�a}&�8�0�4T��ҦC�جkh�7�lF�Fɺ(�;���k���^� wsyܩ����C"�mqP:��۷�w���RP�K�ܺ1�l]w 0��MX��*=���-n;���a��S8�մ�I*Ƙ�/����� �Kh���iQY��+�x�^�s�f�7�^�e�wF��"1��v�M�g�l�U�m
nvo37��ך뷬X�S|�3�q�"��ͥ`���Y'jKs�Z��;��hcb���T���Wö��fhcU����⃕��#l.,T�
rB��Rz������c^e
�n�7��黅��g#����r-j�k��K*B��
UbK��2m(n���f���z��-���]�C�F�֪Y��,81	�J�ol6�p>��0e��u#��*��)c��d��z�%�X�T�\@X;���ٔj���/wy� ;�[��r� M�3L|�Ͳ���4h��A��T`�ݖ��8"8�h����]����f_��B�X�,���&�u����W͍Ȇլ�t�w.��.#gG��Ƌ7���{�8'U�y
�H�����%|9Ϊ�X�!�w��u!DV]_&����ve���1�s�c��)�]�ʥ&����;��ԕ��h��1�Hq�h��#��y,�UW]���kjn����}�m|L�˭7N�0a�V)et�\��V)����4P}u�t�ǰ�W1�k�#w��%�]�9|�E%�T��۩|^��)]���L���2�g*�=ڨ��S��x���2sgc��p�B_V�|�;c��1��s���0n#[�%��}%vo���@b��.����AЮ�0	z�qmZ�`�+��<����!��6��ջH[�]����u�Y6�ۇ����T����ug#��ݜ�U(pHhd�F�t\u(������ʺְ�Ǉr��v)q����73z��LX��k$�6o` 4��������Aq֮ܥĄ��HP��]���E�Ӳ
Odێ��4��Q��5sE(�Y3V!��W���-���ᎃ+)�8��s��,�љ{�+����{Z|�`毜��́Tuˈ�������j�H2�� %]r��vp����U�K:6r�0�m�#���J$;�HO/y���)�-�;g��|]����M��wxK������Wɹ� ��K�L��Ê���-9���	��,�0��#F��T��qr���)�(��p��\�	"�钛7Wo3���|	��2�EWh�Z��`�vr��g�1�����:U�h��uĹI.�ߓ�x�&T�,ZUh��'*��=g�Q폎X3m���`���Aq12��=bu�͚P����/�Ւx�c^.�"Ɋ�*�=MMc*��x�9���X�Q�<<@\]!\�^�M���S���ޝXݹ�,nʚ���)��!Dr��$X��
Y%pg_b�;N����;��Ld����h]��������IM��p�1]��Qm�6���6�Z�ڧ6+�����t�����f�@��Q6-d����T+��Ŧ`ۂs��ßJcr��R^RIe�H-��ٔ�
��T�1����U�щ��Z��!hv:�ΗB�ela�`��gm���@��+
XC��n�Z=7����ئ��ֆ�ܖ)ۊ��4dɼ_]-Ƙw7�ڔ��AQ�@��{ӣ�Ej��\��NJ��kk��owE�$�p�m�4���pW�F�X��]P�8���I��8�c[�������]�˔��aI�0g)��(���2Ĭ�\��{3v�m�-4���'��B�.�b�؟cEۆU��Q���4�K:ޭ�%h��J����B���$�J� �<�IhGׇV�����M�A�ƴ��k�ݪ�JK�=U�v���
_:�.(l��b�m z���x�)���W��V�ف���ɬ��;��*���!�kao��u2 �q��לC�9{��NR�wO�)�)ٺ�l���"�7 �9���E��w8q	�������b0Y0�^:ɀQU�:���k�ۑ�A�"��jw[Ϟ���Z����.��*�7-Y�Ž��cŜv��.nh�-JE�x�o&�+�N�UR�r��h����,��߱���..�9�n�F�:��A�u��Ҭ�-uSwFtN�{�ܢ�ÛQ��:���Ө���%�e�vAB����(Q��-l�>��,U{5����&*�[�.d�������4��&8��J,���U�ƌ}�藊R7q����λ�X|��/1=����F�谟g��/�}=����)w�ňedS�Gu=�Sӧ:��N҉Jz%k'gp���1&��O'�}ID�;��9q�s,��/d�A�}���o����j��S\�oU�\�yf�������7Z�.
�lM�3z���vS�!�������d�6���Z�3�*�C[]W�V^Ұ�'�z��:�J��r�os��v���L�8��j���c7�G��"���}�����w]WQ�3�0�"��c��R�����"�s�ę�)C�{t]L�;K1�G���(Sk8��R�z�d@��T4Ӗ��R�s�널d�B�V��s��Ӗ�/l�(�wd}�8ՉԖW-+��ó_�8L�{��25:��t�H;���p:q|���籽AV�WY��'�o��p}��!%��-�k;����m�1�e��N��_n�z�	�ҕ��q싻l�h��b�4ţhtx90q�\��7/k{z�/��������/�Ç��m��];s(7)��s;kH�nт�Jᖰv]�'-�z9�?gJ��1.R��������[9�[��K�v�^�7���[�C�,+s)A��Ôɏ��/���A\kQ���ԫ`��%f�v�[	�-
����:���E{5]���B����Xl(r�r���M$S�ҷ`��@�gB�SS���C]MYa����ۉ�i�7du��Pq���y#�W��:i�*䱚��n��]X-55���ϔ.���d�Wh�Tn��(-B�<��war���%0PY��ܠTg�#�WkA��o�}H�^*1G }�TN���ѥ�4+"�
���:b�!nAi����%�V�a�daa��1���9z��8�a���`��A��M;O�Q������6ݧ��x��{�Fb\�M��!���'>Z֥�x݃rSVmrJ�S���:u�*���i��0����^�͵���k+]"��}$��n��#U�JY���)[�����b��Qј�Ցo��kKWm8�P�.�nm7f� :��i�d׳K��\�mB��S�d�>u���o �;��ff����Ȃ�C>|�Iܔ��t�0�N�vJ���}Yٶ:��kȬ�Qc��GY�.���U�k�q�ڈFƈ&�2����gRO��p+"�ڲ^ك�\�B�wF~a�&a����vn�o�Yۺ}���#Ɏ�ti��' 9�g2���8���I�Y�军z;ep�D��5#���K;�L��V)�o�e�7�.�E ��̋Ndrd��]�+��+!������'UЧ]V��y#1�r���\r�a�;^�s5!���њ~'C�h4X��$���'[C%w]>Ӫ������Z�D��Sz�C5<U�cj�7K��^�e�=�/�+i��т���l��[}���C�Dj����&�}��t�i'��%R]]nYT����կe���s���=q�̅V��V$ �u�%�nu�YÚ�,񜳶�@U��ҥR��p���»3o:֮���,�n;�T,��ƠW�v0�<X�g���S��W�b�����#p�o��2����ň�u���kU�o�r��yL]��̦�MS���)�V�ӌ_�R�Z�*�˸w&WYE��I�`�]A��i��tÒ�j�F��=��4.1Y����;�2d:�n��<�V�7Vjw#���n�^S����Qc�=qJDV9�_(�u��唵؝z���9>�CuuE��Z��V9T<��ZD��7��f�Jm+�fu�Z8��I2�AS3O�~��-�����=B�-B�o�����m
�$�W�3H:�K�!HMW�w�Eҗ,�_^�]Z��y�5�E��H��;j�(Q-����"�c3ge��I=(e������en�+�(p�����e%wǬX�%A*���M��H8�F��ϻfd�Y��*��E�k�������`y��A�J�IG`�.�l��]�=pw_|�"m��}�.�=���K���u�W������я9+�:*��gU�{3z���Z}�+�մZ�״d�����dP�F!�R���Xs$+�6��fm� b�{����7�5oD�.o0J�:�tG�������*ڑI��v��N�:+���s&j�kp�Ҷ��Z���d�6��fR���	]�6n.�����vA7{Q���@j���WI)�h!7�>��W�0#t*,�UÁ�.�4p�|� ����1�bڏ�t�ִ���*ܴ$FN�n��L�w�K-���]�x��0���q��}H|Y 0=1Bv^Pd5���JO���K�p�+����zr�ʎCԪW�&;0!��SPt��[��am[�_ye[]���()����.��S���4ܠ)�Ţ��7��I����dȩ���z�A����O�mf��kv�6�����3�z�z��ܔEr_:�M�n.4P��H�i؜�7��9�n���z�\�m�Np�rj��o'r���w<�*V^SSy!Ja܌�sb�E,�:�"Eg:�RӷG����m��o��{%����;��u1��8'�v]<��:��Η-u�A�,�L@��]�IXH�]yf���;q^�ڪh71U�Tr�	�>o�1ٯ:�Q�H��T&m�F�4m����"k(�r�^X��e��д^n�iâ�)��GIDa��ˮ-�w\<��QL�c�Ŭl`�e����﷫/u�:iHYܤc�j�&�@��Hi��w���p\�W!e���6j90o)�;��]Y��܀׹ґ�@[��T򺭭����h�#,�9+)���K8���SW��9��gb|3׾8R��_=�$��+�n��\:��؇7��[j�8[�e*#Y��+�'��L^�g��X���n�]�p�8��[:T
�]�K��C����6�̲�{�s�#n�ݡ+zgt�3[un�q���\ _�mR��1=��M��|�e�[��(��N��|��HJ �ȑ�`�q��P�1��z.���,P
��n�Pn�'lLJ�kju�G�i�uw��Ve2���*Rcb�y�=�$��Y�,�p��T�e7yG��˻��)m�M��W�,>L��!5lPD�;S�o�ڋs�H=w���,�iVia������GC��+(2�1|Y:]��������;#�O*5����b����H.��P�R�gn�(gҩ�)��&*sWv��Et�����\)�=��}�r�-��+���>쮥𫧲`��4�b�����-P�WN�f�J���D��4�I��+�]����i|�앮�h;z��(yr����1i0} w���)V��f;0��+}���ʍ��v�(_8A��u���%�e��˂{:
L�ZwUm�rܧ��F�Y������SyκɊ��J�ՙ�or"G�\J�
���h�39��*��-İY�­�%X 	�@��LTt�B�3y�h57_�^V	L@����d�]�V�:�sTn3f^V�v����l�@�7�����+B�7�� Oٽܪ�ͫ ���V�4\4�s���\2�)�ӐfM=;��8 e�7x��W��fB:�9�GFibN��rZ\�"���Vu!C���W\�]c,��B�f�>�v���*��ԤW�++���P}P7NX\�=��J3M��� F@���#WxCۻ�	�7h�E��1'm�r�.��X�&�`:�Ȟps�X;9�6mEI������er�hO�k5��FG�Lu������5�YEvQ�L��h�k����=�J����̾�b�4����U��Eʃ=WM���3��V�Wҳ��AN���5�8��on���TDc;ө6�D��l�����L��`V�nm��L�v�f��=�Z��r��2��iV��|͛�V�K�:j��=	q���.y��X�^�u�!���H����a}},CY��{	B��u�r_a99j�o �{6���o`�V��)�b�3�p���_(U{�:tw���\���Z������+q6ҽr��Sx�b�[b���ug6KѿL[-c��u�v��$/�,_��H����
��90p��&�St|��2v�)�xq����ђ�R�>���gw���:��u� ��LR��9�������Ѕ�4ݐ:\0��*�9��GΕ���/��z�ɥW+�����j@f��R�Zr��O���zA�.^V�ٍĊم��\���J�T �D��>V��f-�հ�Ҭa��jW,��R��r���]��"�,�n�"���G\O-eu6���o`=rr
�i�J��^l��G+��Z�L��	7h����uc�)d�����N}t�_f\ZL�7u��gV�������6W=�MP���;�ֳ��&���g7I\�c�,��q�����1��g@����?`�����,�兜:�]���du/�]j����k�s�IYu���o��}����(S�2n�ť���p�w�����V)f� �g��w��;��%F�%�-�ʋ:��K<��~¸]+��"M��;b����u]]=��v0+�r�8��;T�y|�(1]���U|o'w=�
��D��dKp�����6���[�qE�}���˝Q)��k�٥���99ΛMM�R1�\&mv� ,��������P���8�
��3p�a���RtC!{o_S��5rݷ�\��}U����}_}_�U��}U�}���ϗ�� yY�ve�����G�,��zԙb�r��p,�K[����!�k�d�`ٔqm
쿍qھ�˲ �NlӘ�=)Q�]�Gir��2�� _+� ����<�^_.���v�$���ef!�o]-���/N�A��\�/z�RFwh� �\�)�=ݚ�Kw9ڈ��M�G@H"���e�$)�G�_m���s�pT��G;�O��ue)�җ�����T�XR�:��E�\(�W҈̐.����m	(�]�Q�{��WhI��^ݫ TyK`_f�o���I׃v*�,!�͖��.�|�
x��΢��rb=�J"���9��S4�N��L��1������Lt+�*�1��)��Z��8���/K�LVT�n���	E�V�08�+s��ͭ�aw�n�C�9F1�Y7U�.p�W��A�ͫ�!��0�XE�٫ڶ����&M�S(��.�vh�G����}+���`��B�zb'FR�1V��J�͎��(nv��L��
�hEV��vb�6u�!L������g0*+k��TF�ym���+ͭư��3����� ���Sw]d
�g2"�p4�]�9t�Y�Lٹ��vd��)n��[���%=F���0j1}�}2\�F�gNL��`"Liڂc��@�n�3$���d��/�x�Ɣ�s�ӽμ"I���y�b�vm�4`�I͕2:F,]�����S�����t�Z����v�x�:rc�\43�kewټ��) /iAι97N9p�g�3�>�w�:c^R��G*E>Ԫ�C�R7d�!��NcbyK��C��Ý�觹IRQ*�8w(��u'��(��{_ok�M�rT9�i�X�M}L�X*��p��K��b�·[�}j�b���t�LJs(^�k��vΚ��x]�&�
��Y���r���n���ڱLp���������N�8/Y���1w�/;�8�V�9 ݻ����
�2�ftvX�2�6��`�A"V�}���͕�u��]�]+�65"�g����m�2)�]\Ŋ���͚A=�8�+U
o=��e�.��E�c�v�b�cz��������M��E��9Go�K��Ͷѐb��x�ά�uq �}��b9{/i��!śzév��bݘ�:U����by�A,lW��e,�x��yG\� q����H�R��Q�.� |�C�푼"��YO�DF��b����&]n���m^��K6Vu�T���{�A���4M��A��2�sP�s�2*oU+ǵ�;-���5w,�⫫݈v��u��P�tlHJ�Z�v�J�7b��kz)�su�[�]<��k$��`�0�! �N�H
T�X*�$n+r�\�e���9Q��� ��L�2��M����,U�N���v&,��x�T	l��Y�3:;��+"���_MJ0�.�)G�ve+���{C�\Ժ.���gW��s�AI`�r����	xVkv0��9G�9���.w�o��J_d�+ޖpӳ�,�� Y�t����"��KE���MEB�p��6�񎹎�vsۃ�$�T�z<�+��D�JT���e��7,�:T�r[g��C����gL�DU�
��Ͷ��8��W�M��x#"UZ�;���js�ݬ�w�n��y�;�1�F���_^(�i�BP鎴��NI�NGB�;����O]=9s{�!:m
�($����I�Twe�r��Qw�\�w�gC��F�U!��Y�"����]�;��H�f�L�h����\o�����D�;�JւM����ڣ�k����wp��[����ܴؓ;%}Dٜ���y(�a;vc�H%!ѫ���l�&]�QJS�o����x�Nrؕ�Q�nVD�l��y�3wdhv����͉v�>纓�@I\7^��{��ɴz���nΓF۫{t�fN�f:%�m٠���������Ӝ~c�\���:�M�ʋ� ���ݫ�:,� �����BP��'qf�B.��9��,܁��2�>x�cx�+
�aS*��G:�E�GX�+qt���ɭ��j�T���]��ꙫh�U҂��$�q�M;�kcF�T�t��m�VkR�'1|���*�B:Q���)h���r�i�����7��5o3�`[Ku���4�n�c�n�\��,�G��V<	I��2�Ve���;CB�������`�G�,t z2_!6�^f�
}�PY�5��6�eK��
���:e�*u���λrks����r�/(�%':rR�j<��n��*hOUp;3H�}U�����n$w9o)��B�����Khi[��ہLr��b�{�w8��O*�?8����>س'�.�D�okn��ܭ�f�X�l���8�ݎ��x���p��M9���57M@�\j��@�C(��,f\��ZWM�Lv�G(�Ilb����e���bE��]�Q&���Tj�ֳZ�Z�ngs�K��(�ٴ���	��_ga c\�v���K��ر%�ו�X\�ȝ�nR�"�oђ��^>v�Um�.�Fu�'ԡ�j퓖|�ڕ|{Sc �Զ�Ô�#T���L�9P����	��mMy��ݛz��MB��4�`LK[�ǣX�h޺���_n���نJE�Z[��[�(s6�ƙ	�E�܇�=�
�@e�}��u�%g���y(ZE�5c�PT�C�[c�לKk�\�}P������D+'3a�6�
|���̡�&Y�n�.�=x���Q#)���w϶���-��"���p�1ӻ�['u��aZ7�c��ímu�D���,"�ƑVhl��4&�č[�����YGq�o�L�t���]��y��N헠s�YQJ��w�d"��hܵ�p�AY�.�t�>�wr��n�Yk:�|�{�Kb@7t������2�q�5�P<8��6}32!��v��٭�$�)a�[��luX��L��/{�W�Kzy�=Z���b8�TW�6��uܦ�_L٪P�.ư���t���jט�%�]uX�V�Sm��|���Q�Y�{|LH�æ��w+ӡO�9�������I�Æ���ܶ�}�����Gg�F��B�.֠��j�Ѥ7_5�.���HU���ת�-:��'OQ�*Z�8��;m����51�k�Ok8usܛ�H�}�H�I��l@>�;��uҶ�D�Дm��}�<��X�.�����v:������PR�ʔ2s�Mu»Y91Whǐ�&r�^k���ӆ�.ݼ����,�kaWA�3#:7��q�S[Y8q��]�j�"ܥ)G�A��+n�}�:� T�_"�6&��PL؁�GT<E���(��E��r���;v���di�i�mgw8s"�nK�Y��.���ED�}x����'{���ibMV�u0��r��Gܩ��.ZR˙>l����ê�o*���	�h�6��[*��.iy����|��U��F����Im�ÝS�]6�9:���˔`=V_u��z,t�BQ��Š*;��[c�u)��K�{��n]�8��L��qT���R�vpTƲ���b�v�B6wX��f�"�wᜳhe�Vڸ��q�[��z�X	e�e���u�(L٠ҫո�Ǌ�c�Y�Kpi�j��%�a�<y�=a�AIˊX�vm��u�*h�+�w5����Mk��a��=��ü.���T��{X�<���; ���s/>���S|z�
�++M\]���5�#E����	M�$���<�a61ut��s3:�N{l�|5�Qcl�͎������'m�K�md9��yV�!72��)����kX�0�]�R�ڂ:�+V�jsS��wO��QmA�-7\�w�.�b��gܪ����tB��L#ҙ����߮��*�M��.;�s�r�f[kVCj���e&���K�eԧ�`���D�p�ݩ����w��n�-�kg��%fI�V+��M����WD;�E��י�-95����*�0M�{�&VZݧN��j��W/�>�Zc$j�9j�.ݫ@T74�ԉ�]b��s��y69����4`�ֹ���M�,d��L�j��Ӷ��cd�4� �pE���ݥ�A���a%s3�|��Z0ʝս
N㨅�l�7���e0Mw3��*('�l��e@�aU�:Ę!YwX����9d'N�:�r]�Wr���Vf�A�ըv^��K�h�w��ob��Kt��(�b̨���4�[|�J�k��O�y*�G��;&����V�򘒬is�+���`���+{:[V@�O]�L�m��i�6���2f}���z�+�
5���ݙ��.�w���yȌ[z��Fu�Lڒ��q]ć7m���>b��a+ކ��U O�^�&�P��@�4eS��IT�}Z]R=�b��u�	dQ�I�7�=�{]:wN��B��rcS��[�z��p�;��cz��r�^�S�7e�+O,K���ձ�8r�$�M��q�N���'{�u��c}u�c�����ޔrl�t;���3�'BjZ���'V���Ӹ:�H�u�fr�UI�d���.Uv-�a&���4e]f̝N��,��j@M��F��Z��8�EggwٸW8S�(mf���� ތ���)�m�˻4\�[;;r����
�{�R@b0��U%��X�k��E+l�s�jŶ�g;��+�p�ԗ K4�L�ۣK��Y�y��o�wR�.]�׏_eJWI�R��2�M����`�&��޼�F�L�q��x��[f�}G'n��hi��Ǡ���v)pH�sD۳.�b��if���7�v�:��h7��GL*Q�K+4;��*���IR
�+:���Ef�	�iы�i�.빩��9�Cr(�م��7$[���ӏ�8`�ݞ\�J����s���;KhV#h���p�9)VY�E�8�D����
D?�	�M-]}�n�T�+�#��(���*S�GM��ڷ��l��&�[2�G{Ǐc�,G�O��X�uд8�0Uo��}�z��7R�y�E2of�'�A{bݧ�k��b��WH������I\�W��T��]�%�9XxJ�A�Xƽ�S�x�wo,U�tR�ݭ!F�L��yw���Mh�r��M��V�:K�ʼ,w:��]�~KG(%L��c9�B�����k.ҔɆn� S��hV�)0n#ՊqiNָ�����D�z��'�i���0�{mS��s�=���j��3�ע�3�kv�U��"�wm��)J������x)X����Җ�"�hU�jp�fK���>ٙ���Ƃ�/�Z��Ij|5õm��Ӯ3*��6��3+[��;�>������І��]���25{E�:��͝��i��k�<�7w���	���:R�`7���-6�,���ݴt��L�O�'���C�r�;�y��Ae��y��Ԓ��_v��"�>
x"GF��.�P�WT0r�=�\���M-�]­��G�ou
F���k{^���,5׍ÖCqɦo���S�Z���j�(��N��Aa���߶\�R���Hr���]^����2�b��ή��̼\T�B��K4ǧf�q�;i���ëiR��N���^hz���]u��#�"��1�����Pc�������g�t�.�@u�.������+�}�E��]䋶���(�/��&��)��;�OV���1��ч\��+�ӻɫ|'m�� ���{�Ӓ�<Tf�F�*�	��E�YZ�q���h��o%b�������*�T��ȴVN���q�wz�������YP˚���<4=�1�]ܝ͈���F������ A�.JM�S���=���*v]�Q6�B�ՑF�M�v��YQ�o����2� ��4!����t��������sMĩ��C�g7�/�P��r��w�v�!����d-&nĆ�Êwe�rȎ�/o�r�cGF3VC�{"��G��+k���;Ov��W���G\�m�}�;j�� �Z�cp^�yۡ1�4��9U�ZGC��]XM�U�d���&͢4.�S��[ l�-ݙ� �y�����gq�[�Q�K�ol����]��빅��NX�%8'�R�l��N�C/�Tډ����Ƕec���N!X�ڡv0Bs�[U2��#�-T�bf�d�U�&Y�����d��xA�A�l2�k�0$nn;�[Z���������s�B�$�G$�
ӏ��u���������˙A��x��).f��G�cOFC��>ێ�	Yx�ӭm���'bgM�����V�Ɩ R�j�%t�q��ۯF��Z�}[r>���Iuf�,��w�Uٙx�L,��D�����Y����5�Hu<g�^ۼa�k�˹�2W!�6�K�U�;��������X���'R��9lD%ֶrve��=\p�ϠIIPӶ#�4zQV��`
8;:��ұ����\�1io�o�[1���v2�9mV���!6�jWjc��*v�ԵӭtX��^S������M�]�C���7��K��J܏���Y�P���9\��J�ǹ�}G��(F�U��J��)�������Ь骻j^] ���3%rl�5�̻͋����i�]���m�JWX�ݽo�=�^�I]"�.�|�76h�������ܭZ�L'dZ��gAxƌ7yqW-�n,J���/ ��=��q�oمҵ��<��+�����i+����]�Ɖ7�Y%�8��U��$�R���n�Y��N�jr\Ĩ����m���̎��QѪ���
�
�J�2F�
^
c獼�ymY��Z�J��t3i܎�;�}�ni��.
Òv��3v��4M��GH,��<��w��<�0����^��9v��ƪ��^���ܵ��+�v�Z��d��W9��v�i�X�_=zM����U��id���3n�jl�W.���<ͦ��\ zHw{��z5%Wf�,�=��L��
��x���kB�5�ﾯ������U(�0'k����/pD P@⮹��2��ގ�k;�7LXI��9f�y��l���wF��'R��m� �)[�������,�$+��X�S�̽����.���������X� b�I7xOu����w[G��Y����3��[�(���y����ɜ[ܨ˅��)l��� ��W]�dtS��RhM����s�5}�{������i.��
�N���ǒ�lB�V0�;�&��\�(���� _m0��y��B�t�V�[��<��Bl�zk]$+�}������o�Ie`���مJ&%��5����k�R�tK�����0D$t����]׹��� T����Ţ��E
]Ƭ����9��$���:��h}Xۈ-+�[K�޲,�7��'� �`X�.ޙX�����2i��mu�0:����O�6�Q��k���sv%��	�H�9���
X�9�Z�{�Et�쥸tgd$Q2��n+��{s��-<��P,�u(#�Xd$#�=E��p�"�{.���ze�N���5,�WuzhQT5�z��ޮ��ׅҲt�YQ�:n�W²Ȩ3���b��))ȷϦ,�����Vx%�*1���W�W�r;�)�wy�,947�!T!.6��mWU�W�Vp=@�hY�c��Y���%�.%7���k�}ϴ�����u�mD��b�a�5�s���H�wqwY���20c*2����$�D	�2I2(�WAi#	b�s�#�
4���R�cF"Y�$R�]�p�#2�2�AW5�ba�ur�3#�b�d�D)I	�	���bwvm�ubs���!�Q4�b#%��ف c �hF�	�1�̃#�Q��%���Q�d��6L�D����Bd�w1A&�
D�l٘,�v�cF	CA��f)�&�&L��'ws���D�0���4QL��I)hM@Db�%��I�1e�&LT��P%Uq��{0��uG[���zB���#W��g��X �XGp3�v�z����YG���OKɭ�2��f�:�}U2TO�uw�t.��s9���0�4V�eY���n�S�s��ָT#(�p�H"�����kOUUj -2=]�Ek��?p˩l�u<����gr� �����h{(�ӿd}��N�1�ǋ��.f~ߑ�I��˓ۆP�1�\��:��S��)Z�0�cܳ�ֶ]�8n`�����y�<�e֟��Z=��\=>5vxz]�����lf��v!boN�5��`oR�a���K��7�^Zo��q�?OU�`]h���Z��9p[�&u�o�M�����E'2=�r�1i�������
��oD�r�+�d�b�^��,@����w�����s�ppv�>;5��K�P6��2��T�_�)5�S���D۵�۠0@�!g�D�j�~ڢ)xo�g���p��x������b���r2���m���8����.`��� ;�H	�w
�eb�0�3�77��OS���j�a�X+D���Xm�l�u�Ƅ'�^|���� O�d�6*w��й�z�VEP���1<��b�HJ��3+��=ղ[��[�纪o��d��%K�Wz�w��|��ˇ�,�.ې�P{|$������zW-є �%.�s��f�ܷÂ]�r��woh݊����Kܛ�:��ˡ�1�UJ;`�����m�x5"�#D?�*��ӿ������Z_�U����B6�D�5d������]��>F� �D��۝��DRs�F�ͫ��=�9��ӸcOc�����)_�Jn����o��P*��ޣ�Xr ���mA�W+�$W�e*܀���űOVm$�ի��H���n��������[O|JGv��&��ܺ�f�Y�h���d5�W�v���; =�z`���Z�K��p`����y �wN@!a3��7{9"�[�f��V�0���*�֔�ț kM�&�-7�t�[$-1�~��*��D��^�e�pq�&���4LuG*ss�ύ©��'�J�Dp�M�h�o`�����]{נ������Cd�0���e��Ԗ'�6�I����?yU�V/_�� $�]�޲��G�>�*g����+�[-W����TX8����m)8Xe:�r�Nbpgtކ��F:hߜvĔn�eqӳ
�U�_�Z��x�y8 ž@:�U�C�|��@}�d�J��iQ���9�2�n9�� ��_x�T��Y���t�c8��]�QU�)���ޞw&˧�����܊;�6�`�WS�{��g�%0r�s�5�
lCT+��v.��Z�bD�����홤�����W�]u�;����G8uh�U3��E�Z٪7ș�wWR��\j
1��!� `�s:c`�/	ŝh��jY�8i����z�W�-訞��kN���d蚭'Db;�|�뽔���k�DEً�������ig�(@�����x���0����/��9l�c4�7���s<{�#��Ҧ�ӻ�o��A�Z���|�II���+��&^�ͩ��
�Sg��zmL������R�R��<��jK�676��j]V�5/H!����i��Dt�-�����]pA���W`�hP�#n)�(��q#jj	��?(��\M��y���!
�}p�9��[i��:D4O{����n����b��E��`�1_K��$x�����hpڢ$K�+:�e�G���~}�R�e�V�"��}�
Þ���������� "��!�io=m�w'͉�E�')��_[�qƈ�_'U8V}����@u\k��5���I�
�ݨ�5��$��xy�a�m]���W�z�G'hqr��/���d�ڝ�MBɧG��W���ͣ@q/�uDr��Q�8��4?L��	�=��.�Ǌւ��^^�M��
z�δ���[v�:��0�ׯ�A��-���:�c��)�z���w���T��w�l�+ɬ��[Cf�n+�é�£���@b~�����Hm�(E����N]�
�<�zP1�]Sf0Ný8ˀ/|E�}�W�b��g��Χ�"��
�}�Ƅ���B�T�)I��z�_D���֢m,��9�<c"	Cp��{\i=���wCVWxN'}{;���@�砧ܻ7sE��M�w��D֚���W�R�>Kì�F�#����)���g���-��:�X�]R��LD��BmMr(���q�Z~�o(�� ��p�r��dЎ����7��gH睎s��CQ�#:_m���,֝'[�-�uҳ���.�G�{|��m'eb�\QD��.kN�ɘC��yc����Q�=1�R�C{|;#�ܣPx�!OF+��B���N,l�rb�:���/��u�2��]��\�];NW��F_�N�|T�;��(<�7wV�[��]�_R�Z�#Ἂ���:�H�=x��3�*j��,,  �j�$F�����W�=�k1�=^sg=m
�\�Z��d :�C_Y�U�B��K������<�4$6g�v6�;ud(Wnvn.���WܣAdw���]��ˣ��`�]�����z��i��Q�5�u�V�҃e�i�����ok�_&�V�8�R���u�c���]N��7iPys��C)D�y�z���b^ JT;-�r��q����q�::��t��{�U_��\�B�S�2eJ+@�ȊwB�*P�Q;|�� �M�5���ڀj��4�T_��F4s1�,o��VӢ�|`�h��Y�U1VwK���Wm$-Ȟ� ^�ʘB��	DcW�,j</����|`�j2�!YRc�;uh-jQ�rw�ٳ�EH�yR�ش�����d��Gt��>VG�D1A���N�8��F�RV㦵�t��%dH��0�@�>��>׌��^����:��5��>�e h�&/
��id���G3� ݊#!c�(��~Cj"��<����ew*��C��x�W3I6ʎz"3sh�k�˙��P$�|�_����c������~+�7N���ؽ���T��e�vJp�f|т�v>�:[ʨ}�N��f�J�
�،�-��wE�W�5zW��)�/���~��{lR�����5�41������r�����<&@�ٔ����Tp���X��	È�w)�)9!<�o������k�<cVsCx�gs���*dZ�t�����ҝD.I2!j��\
��a�yx�R��8����%]�e"�;=ϯi�6B�̤��&�8JZ�\�/T<z�)!Fun�}/�zu����" +yV9�Iw�8��V7.� �m:�c__H�}R�%Ht+V �\�i��"Kêg�,B����g3��>UY9�5zo�d�C����j]��j�z�Z�)p�� �o	�^�����S:<��O���ʇ�7��.���]�n�e	���TR���L1�k¯��.&z�ӷ�b 8h9uM���a(����?٬�j�2K��ׂBe�L�W�{Q��F,oE_� -.�b���.�ڷ�.N�^��}b��nK�6xp��UD;�n�w�h�ϙ6�������+��P��V�,�y.����4	��T�&0i5ǑZ�����D��ϲY�;��a���17�2�LM5�v1�"&_���،�*Gvh���!�R�O3Bږ-�{d
���#���@�}H͗�oQP�/J�t��@�l|b5�E�[O���P���)
�Z��5,�����R����^�X ����FB��q(!`����ĩ�93�y���3g+��[5ٰ���!Qv��ܺa�s6���J���^LƠ�-8jP��rB	��to�:r�; }��a��:�+].��M\�Uw[�kS�_�8�֐:�Sy���a�a�4���hb�OB���fv��AB^�>uxD�x';���Ԅ���W�_`��tls�9-��n��{��:���aL�U��%�ek�Xؼ�ӗ���$8N�t��)����6�wU��A��d�׳-��T*3������K�u�C9ZM���ӹ�-�z�n^���p{궩�}��6N�0?Gl���J�K�2T�Cj���y_;G*A��ݱ�Ѵoq�q�qry;?-��0øɇ�Y�gb�co��3�2VI�,���`�ڬ��}�6q��)X�6����@�U��b����ë=���E�@[󃒮������>�Z��A���{�@Xu[�kB|%�g���nկtSR� P.y���RC�z�	�oԜ> �.�|${~��?t5���)��8- W+������)\�4p���n��N����*~���n1�g��Y���޾�L���
��K�������o|��^�R��`��W�W�h�U����~��>;�m���I��?�܍��Ì�a���D��bPb3J���@��� X��nvdSϡ�A��0\=���r���6����-���k��h*Ch�0�?��RF���@2�q7��[�Q)=�|��C+�]keT%��x2p�F��#5T�y� �Ck����
n�m�dU�	V�X��=y����0�����>�=>1�Z�J���Ch��QT�.��o��<]zѷ0h��Յ�c��]�v�ws{t���Ԟ������gf�%M�m��yp9�S��,=F��svH��ˊ�4�ρ	MA<1R�!#��\�/s�]pQ�h�����I~���0�_z�c�������7�y�C� wb����QR��ՔcY�v�=�jɨ��y�ur7۸��Й�.cDp����[ܹ&U�`���Y�Uc�.��o=�+	�j�!�Xb�pc+�<���9��9J�o�b:S���Y4�gU���I�M��q}&�C����Qa4���Aߗ�ej�zy��Trul�A���d8[�D����;ښC(�Y\�����:��y��<�_^.����J��׃ks�Ŝ@B)�)�����qݹ�y�yg�wWb���m�ѡ��k+�R{�AZ �]Be�g�\f��F��oXT,�97��5��LUVzI]�҇*�z�p�XVv$�Q���+f��/�s�bԚ�#6e󺈨[n���΢�Ϲ�/����-l*���{U~�h,�+7B>j���R�3�k5��K�U��*��r�([P�;s�tN����q78���Ȍ�[-B�̬隮�C��g�k�̈ਃ��b��wSEo���/��H����s��ެEֳlj�`�E��𭕩;��D o�6�e w�a��+�f�p�kY�.@�[�:�;�� �@�dZ��G��=Cen�X뵐��J���� ;7y�B����V.nk&�R+�S��.�b �n�
Z��{�K�a�7��j;���M,�IF��q���*�����1f}7�h�iN=~�ԷG��+tI����M���uhߞ��^�:̅���r��F�y�Ch����ek�Ϸ��	��Q���Zc�&�EO�����萭���E`�uO�xS�EfՋ��������&EE��H9l���Ct�(GC�v�g��QV�Q�l���Kw�b��S������qu܄:9�k�B��F�rv��h*�pk1��K�l�(���y�l#�:���Bc��=D�Y����m0����cQ�m�qR��-�Oa���Kc;��[&/�㘘j��11GC�d�1��Л��*hE|Ύ�	��P]���*�Y�F>���K2$:yV���r$as�R��񙆼3.8�!�5�E'c..u7�Q�ѩ��}v\Fʠ#B ��Qnd@f�?!�yDu}n�M}�itv-D��1���7f���C��5L��i�\zWEorQ�ǝ��:8]T�U-�-�WxB�B��RS�#%L#1��j��`�K**T����o�u�٬����E ���U�5f�w/���vu������6Ƥz�q�Õ�ԩ�7�y(��� 
DS�/-RgK�o���a.���
��龜���'5 4|����HU]��ܲ�V���l�u������fO�N�y�����l��˥����50Q���GKyU�����6��1�yYpv�Z8K�k��p_��Y�QXb���)�͞��uu���CK�"r!>��R�l��u��S��b�E�&8aɄ3貴���*����i��:Ѽ��7����:�3"�A�;E���M!�o��è��u���lW:������j�TE�N�*�'p�ou�nק��+T�X({c�c�~�?�GMϒ�g=W�"٠�otĞM�G([0�sW΋�A=Q��KK�0���X����(h�B�f�TO'��
g�s^�r��l�ݤr
��a3��eCr�H�ɍ�q��]PQ��$	�S�8���`#V����6�8q;�8���7��Q����7�<�e��!���q��Un��f8F��c/�Nii�z�I������*�I0��H�+r#U�I։ͫ��|'��C��G��k^�U�Ϗw!ݷ`�����;yu���\��`y������=a7��>�V����Y2noq`s�a�<6�]r[�#��5i�V��o�fVX�ܙ��6��2�k/��:���JWX�*��E�*���H}�����I��)<W�&%D3�m�v9M|YH٢�u���u@�w2���Z唳V�ٻTS�)i�r�����5�lA;����:ܼV��qpWt3}=���7�^�̽���߂���V��N�P��y��3Fwr|�9p���H���i� 0��V��-��Jߦ��R�:.��-��/�ow��u9tM+E�rk�(��K�v�Y�z���2	d�,��*ꝃ X&���Zlh��P�a\4�����{�j���g4����s��t�v_:��s�-���%���r$�_>�XV��oTs�n���ا����*�[�v֬�e�޳i���:��ӱ�0���K���ӑ�#|�J�
��X���"ф3��[��4�UMO��u�e�����2q�6T���s�����݇����8,�Nun���cn,YҫJ����a�-ݍ��ƥ���HR��3��+u��^Ю9mv�~YL�y������߽z�����c:�
�M<0���Ȓ޻=��/|��	�5H�gv�Lٌ �6�V����O�a���wh�x�n�t�:�j]�ְ�-�ߚ���w�6-�[,,�0x\��k�gr��m�[ۗ�)>�t�8�nMt��Ղ�Y���@�ʎ�:���k:�<�Y-e�ǐ3�C��r.�[L�^5�{�X�}�U��1Pb�7f9�(j�(x>�O$��Ck�/'Z�#tc��{��6����Oo':�f�!�!��j��U�u[6��--�^O��+H���"��V+��JR�F�(N�X���۳&��C���#u�^ǆ�^�����X��'��J.�O8���n��Z��v�
e���ç���3eը��0S��bw%�:]�8L������|�e���Ȥ{]6*λG��HG�k%NZ�����Xl�:ʬ�_ȹ��)�Fԧ���������J�	X7�оo9v��{�a�A	�K�$�]*�Ip"k1T��uթ.��wI_5�����yeʼ�1��f\μ55h$��6�r.�@f� �v#Xjզ�!!X��<�x��n�u�R�XX����w��.�`jt���(���������������N���ɹ�Wo�[pwW	�6�:-��v|7vL�U.�y��F��;5T��	�[V�;$��z����}���sv�,�5)��	C5�Gh��ʦ��wƣ���6U�Mj_Y1�q�!J^�xE���Ѻ�,�f��Ǖ�(�CRj�-�m���uh�ъ�}t;y&c�9��Pc%ܻ��b��N�;�C�-�<z��b�^F���X�����%.ڝSsk_RYr�%SL��u���l��%3/k�������??�w��	���dT(� �b��1��MI(K$6JfA�.����	)$d�
����u#9Ѥ� �.�04������`�ha`1b�JC��(2&�!!&	���%%a3��%� L�(����29�Ɍi$��0ɓE��1�d�H�)&F�����(�5	�%!��22�d���ƒ0Q�D�\�(2m$r�
d�B̢�X��r(��]ݤ���b�,.Q��)��mi�fj"f%���ߏ����;��~��Y�h�b�}�[!��g��$�Z���?�f��{�;�FqK�+ǎ���3��i�r,��M�(���[�����������/�5�y���V���d����o^ux�*9_�������Z=ם7�{_�W�����}W���+�������<��nDD�"."�����1}􈊭��f�%v����{oi=�V0��b#D��o��y����m���5{oM��}�澽=������r���߫ߝ��������Om\����^��������W��_�~���]��kAo�G����Ow�뷎(�����"4F�����y{Q�?�����?��U������~���p�}�~z��ޕ�{��Z��]������W���ܟ���ž+�����F�7���_����h����̲��7�j�MG�C����}���Z�o�^7������W��׿�~�K}W5{���{�u_W��zk����6�^�ss|~n������soz����n���o;����y����ߍ��� ������̼v��j�_�Dp��-��_�ߏ����U��k�~���WŹ�W�;z����������[��-���^�%�������ͽ?ʎW���y��^��^/��<��[�D�b#�D�wgK�icW���-��"�5��}�]{W��꿗����*�_�������6�{���_���z���^���}m��'���⾭����[�^>���}��ޗ+�������0�@��ovU' �ɚkc������y��7���W>��瘮^�����/]o꿛�~�?z�-�/��+����h����J7����{��W��o�r��^��~b��s]���ק�\��r�����o_;o��^;�>}����|j�{��#sT��"Cﻪ`�6�W}�����F����W�:�V�����Ҿ5��o��z����o��??ݯ��^փ{�:�����r���^>5�^+��_�����W�͹�~���護4�3��z�֮]^C}B>" ����=[���޷��߾oţ����o�+�o�/{�Ͼ�����5�����m��m˖��{m������_��~_�׿޿��ߟ�_z����ߟ�����7^����� � @�������皽?���������^/~o��c��^/�~��|����W�\���y_���zW����ּ�nm�w������y���|W���;����o�}�>��T�uC2|�\����˵���K=�,u���rio.*��3\:�Xn�¹�j���ﯝH��T�w%�+��b!K�D�A>e�ui��>v:f`����ns�H�\�!X���9}��u �B5�Ff�Ù4�B�]�0������~�;���$Dp����׮������~�y}m�r�o�_�����o������~5��x�����j������������Z��U��+�}��}W�ѷ����zW��^5{�?������@���a����z�P�}b",G�p�z�_�Ey����W�}����|k���������וzk/{��/��-��>y�����������k�_���{��m�����O���z����h}C�"$G����$[�^��Ϳ����/M�W�͹�y�����r�~ߝW��[��^������Z?�ƾ����ޯ�x������o���}�\{��"(B|����*&�p�[���]ˈb>�B}��f�j1����w�z�ץ�~�>u��=��{�ux���}^G�G/�]|_��x������^|��+�ߘ�k��ۘ���b>�<1LV�g�vG��[��}�{~��M��[��~���zWչ��Z�_?���\�ջ�Ͽ��{[깿<��z�߯�Z�_�����>=*��^7�n\�����v����^�����我�`���B#���Et7iD��I���ϟ���޾���zo�~~�_���Wy���|_�o�{x�5�7���~}��W/K��������oŽ+��Ͻ�K�\���]׍s\���/O�*���{k�or�~���������ϟ����\�w���Dc?}��D }� ���H����^�����}_W�ѽ+������|���W��~�[�\�}�x��x�������_��.m���߭�=��>" ��$D!?W���LL��8�*q?��������h�_��^��^-�_�F߮o����;_�6�<o���m�|W?�|�����������{|m���KG��<���6��[��zW�z�x�����b>�(DD�\�AtrL[s(K-�x�W���UAT��>�)
�L�R�|W���/]��kF�W��޾u�W�O^���潍�no���������_���ץ�+��W���.�ֹo�s�����o�����}��Ž�5����������^/�:����L�Mվ�������]Ro����nW-�{_W��_�s��������^5��{^���_�����~��x�^��������^5�ݯ�[Ҿu�W���߷Ϟ�Ǎ���Qw�#ؚ!d���7c�Z�<��E��G�֯�Kqc�i�Ռ��:�A�A�z�Ǻ�![ʰ��F y`�{���@��1V���9ՠ�b�7ݵy��Ͱ*V,-����r*�O���mp�b���F:Q��gg�*fʂW���m��Ώ�C��">�و���|����������_W?����76�z��|���m��r�o�����sǶ�W�_^/���zZ7����~������ߛ���o��x������;��μ[c�Z�+ˀp���G���D��9�?�~*������M�ϫx�/��בh7�n���~{�������k��_�r�r6�s{k��^���_Ϳ����5��~7����{��_������r���X�w.3�l���}�3>��7�n��~�7����x5%}��y{|oţ�����/Oj�_�|k�����^���^/�~z��x������{^+��~}��ݯ����W����#)��U׫����^�̓R���}��_���=w5�o���6�}�j�����o]�~��+�~�oM�.W�������[�U�}�祿W��_�s���U�_���k����{Z7����r�_�#��w:�����E�^1��k͜�����r���x�o]���(������*��o���K���ž������C�ou���^����������W��W������[r76�����{o��f}���|�A��(4X��2M����?�����~}��\��}�����oK��h�?��[����ƿ=v�~.[���oKO�W����{k�_7������~���+��o�w����zW�G����������*kc̺9s�ts�;{A�=w�r�77�����^��W/�ߞ���5�W=�~��m�������߾[ӛz���o~�x�wηǥ�뽭��޺�_[���_��^9_��o��*0G��}�>�^��D�:�=�e�;ן/�^ւ������_�W�~|��>+�^��������~�Ϟ��~����]���x�E��/�W���뿕{�w�~���~��/���6��׾�7�o��o/޷���^���������\��P��F���X�=/�`� ��W����|�[�~-��]������U�y�����[���U�ϾZ��r��￾����r�o?|�K��o��7u�snʹ����zk����o��������=�}]N1B��F��>">�I���m�ܷ��ޖ�W|�|k�����o��_ן<���������<����/����[�����ޯ�w�p����W��|W���o�w��W�}{k�_|�dw2�mֳ�����_z�ޣ�㮮u��.h�L�+�[�ǟ^��zQA���A�s����3FӨr��m�:�Z,M�3ia�|0��6(A) �����)�'#��kQ��ܗ�n�V\�äv	�d��}U_B�t����^?�c{o絼nb�h7��ί_�oj�W�μ}_y���[�����#o�o����-�o�����߿}���[�~y��6��|j��}��ޟͼ�ס�g�����<c�=��9^��̼o߿������~_�w-��~�z�׍�h��.�+�|W���b�h���~ߝ{_�Z=^��Z��_�xߗ�����k����w���W����������-���}�|[��sQ]���������T{�*(fA&ͮY\�ס�>���K�����_�ss_������ѽ6����^��z��
��v�[��^5��5뷧5r�+�y���}n^�����+����{W�~W�k�o���_����/kG��דZ{cYۼ�8�">B"8G7���������}m����x�5����ޖ�W.U��w߾����W�r�+���nF�s����W<�|W���:�-�ε��{ߝ_^��^�����[m�qإeut�!�=�
��>�'�{������կCo�����7+���k���/��_�x���ߞ�m����-���ߚ��kA����ջη��oWߞW���o?��Z�o;ү���뗽��-�DG{2N�c���OMy��¦�}x��_������w��������n6��^�忺��n���}����o��m�|S�L\j�(�mTW|�5���/!ㅱyK'o��z���jQ����3���#`���@O���ƫ�8F}�F�Ǖb\Xss%U����FmN�{�a��h�j�1�<6��e� +��\�;ȉ�{
u��3.Sl��{|r�^w���Y�y2�s����;���)j�yc5�	ݝ��m�z���@[��'���\��i,`�ws��SY\6�ގ��'��փ̹~k��H���@��2�)�Q�T(�{�
OZ�L�mח\�^�Jq���R����r}�o�jƥ���eش��Ҝ�l�V.��!J���Go�`\%M��n�}��+-F4�gk��Ӳ����q�֮Vs=�Wt�)��:�˛س'eoq=���_U|T]J�zϨ�Ch�٘�r�o���1�q,F#_s�4^�kN�}��A�M�n�Y{�o��T�j<�F�?}ia��o��d�xn!�l�w�y1���p�����H���z;ŧ����N ���K _5��n2x1��w��ρh�|O����Rw�Z��<{Э�j)}(��rK����T�#��H�+Tup���D��m_����Q<��D�sE��Ů5X�p�sn�Y��O���Q9C�7��;��@�{�(��t�pL}'����Ce�tt_^��Lq��.�a9sP��m���tТ��9��T*T�]���塭(�����Q���j��{!��S˩G���(p���ʸa=P���1e-��j=�]Y����xj93_R}L2i'�%m֞XYB��\�+.܆u]z���j!+�D���Β����S�q�6ԫ���J���6z%M�|*d��xr.������{�uXh��ԍ`ƛ��_[�䱲agݲ��J�K̕1M�~����F�kp�ʩA:B�2�]2�\��u�r��BӀ��(Ugc;�}x��3�W�#�9�v�0_ r5:���!��1/#�]�jb��AݬU�ٍm�)�h��}yɋ�zF�VS��m֙��Ӑ����h�)K��.Z";3�D��7yi-z>�#�����jU��~�mo�-�)ӓ��?��5��{�<��:���~�]����w(�[��uZ�C��k_ܫ,���~���3X���J+��SǮ�R�n���tH�A� ��ƴYϻe,tćq�J����gZX��eqӡM��Ӯ��|*�����k�M��{���
��&Έ�0�N�	�V�Tur�AK�E�8r��0�T�cK��>��x��hE��o�kʞ"^���:�/i��o}�����P��(�x���J�ӛS�_R��n>Φ��ܴs.X|r���-gg��m�Y}һ}O\m*���K���i�5�]M�������_ڗ�Lv*�O�馤��s��&��ڥsU� (��JB��b5�O��J�HOj��KO9ysx�ｗ�Rz�\1�w)� X�o.�5'��.��K����Ua�Km4����8�ˮ5{��:�)�#x��\���B��@Kf�

R.Dѓ��]�1O=5yD���9�q�{�;��HJ�:9!�;O��d�D�S]�{��m��vp�ϕ���sMw_H�Z���r�f}�݀8+�^��H��#�y"����s�Zn]EawSvu���L�|{�f-Ί�-�z�MW�B[-�UKo��}�Gв�7��nOUdX{L{pZs>�lմ�&�t6f�:����=�z2WF��.s!�Ѧ�I(bƸ��ޫ�&��0��1cGY���Kϧ����[��ڴ��ʌ��ڣ��[���T��}�=�_e��i>�H;��[��
"���9�Y�[�Kt�fݼ儌����1�;��ԘZK�v(�U���刺�¼�l��t̋�\}�Y,h���ߏ�}a�T	���b��`8`pO��͉�S{\i=�	mf{2Gxk�]>fu�Wts�����\S��a9�Ȭ�����^�j̪�5�?��H�l�U�Oo��5� ������ԥ�U��p���N�#�Di�?SyG�s�L`[SPS���S<��1ʬq�B�&�F)��Pq���8������wJV��>��r���ף�{1�g��ث�(��ү���J�SE�OL+�O�d<YW�t��KmȎ{r�^`��Ę���w�������K�Q�����}�W�q�����X��|7�J�r�c؍�����	S-�����ҲK�qb��P����赖���N�GYu�����Ōg���-n�����Q�R�c[j���wɮ�V��Kx����Ù��3vut����h�s�Գ�V5ox�:�VO�>����6֤Z��kx���h˪}�Fη���hz6���<;������ 9ȅ%��u���8k��̬�.#yWե����3����pwK���YVy!���+���j9�͸�]!�ZU�(<�T4���|4B���έ��E` B'1�����5�Ƕ��o�<COS�������[$u|y)�7*v���-��`��a�ث���h�7��J��.�:<���]2 �v�*a���¸Ư��xtC{\T���o��pp�j���\5J�#[Ӓ�*�:���L;�}Us:������L��k5e�nt=w2*hC�a�� C�ȑ_�0�_Į;L��ձ14���Ƙcu�S��G��~�[�9�'e}4aw�kE�˪��r�������YB���W�1�dh���<���{ȩ�/��Vr�	'��>֨�~��L�,��L�+�pВ}Q5��%�$h��6�us��}���5�t�ۻ��0x���GKyU���æ�da�,���7x�J���qd��1��\y�gjծ��G���swS����uGwC]E������jp��!��3jc5b�c�x�d�D2�LbX��yP=�q���9�kK�Τ�ހ�Y.� ���+lK�q�޵(��w*��*�-#B��J�ۿ�����.{��K�>��蓼`aC�
�	���59�_oc�c"�Bq����'�[
�o�w>pT�"����q�/���0pT�WZ#�uҰB�v���@WLZrB�H��B��j0m�WW�5�/��/~^CU���6@���s���_KUΧ�C /�ϗ��5���ejT3G�N�d���8�j�)��lGX_'��Ip��S:<��O��A�{�s8k��&T^�rfĺ�ˍN��0�n},Fi��(h�ySǴ�`4��u�Ԯ�5��D$,��j�_ѓ,��9���V��ې�qQ�c�w�]PQQ�f�t�c��g�ݒ����>�j��X�k7���p�9�=+}���-�;�ۗ�S�s�ie�����>�����Ɗ�]K�tm�)� �K��ܰ�t`�m_���Un�)��qm��M�6*��<���1�y���|��*WU�b��>&8;���㹄��}jZ�rȠbAo+����"�1��dd'Nn �f����&�~��[ �*�׼��{�����2w��\�=@T�W�[�]xC���>�����G�h��wr-��ŝ\����q���.�D�xge��,��V�Ыm���*պ_Z��Р}�i�z�Y�Չ�z�G����r�c/s��MD��s[ȶ�J�xȻ��U�W�|�j��L�7Ư���T&�Ȭ���Y��n�ޘ ���4�P�ĸh�F
^�����%��]�V$�����Ȁuӟ�L��	�0ɤ\��V��v��P�.Iz���u�y�R�C�����抈}�ؼ�9����Y1���M}*T%���r��C������2�
��7k���W�z��C�(;J�K̕0*���p�\�5Z�",�	0���w�H#\�v$�9>X���t�U�.��N�� ?sz�+F�{o��+6��U=�x���� B�a<�#�JK��X�ʿk��R�C�,���Cf݌��\]���{H �~@=�\0ϻe.�LH>��������qgZC��rQ�ݽ>>�v؊�(��T^��f��.�:d���w��Ty�o*4W\��_k��K&�1�{�N�O!O#Ԍ�vvZY�S�R���n}��y-��"�v��Wɱ�ӓ��*���w/��4_�,BF�(Jo�UQW�M���cZ:R�Lu����T���"����i������\ae��
,�	͹�,[��_�l\�9���\�f�{!dX�j�f�J���T�۳��q�C����v�gc;�ob��$���_�,Xm�t:K�Q��]GԪekxbs3��*f�MZd�@���s0�+���qa}O���I��O����V�f<��;bbx��J^Q�r�dr�;\UHok�z��:�u:WgRчA�E!w��<S�/��F+�Z*r��Y�=גmC�	����s�ݤ�M�رCy�uG;�m�w�%��T�w���zh�C�1�-���2u(��zE��X��!�)����W��`���t�9�Vsz�͠"�*���c��ܡ��IJ��L�S<q�d��>��,�V!�v�X�ƥ|7�a�Au+w��U��G�X�FN���M��i��+�{V�,:r)�_<��R�:�7�2�>���uZ��
�1�?�\���'|�cQG���(r��Er,��-��*�e�&�o���sQ�ծZ�Ta8�u�3�wwdμ ��	�F���gk���,�ݞ��+cX�o�Ʀ��u
Y�R�֚Hev�f��˚kjMX�:PW7d7Y)U�ꤨ-���f�}����.gjD�.���yWYb�
sv�(OL���N���-�Y����*�tH�{��$H��H���f:U��^�8��]1IjC��ZDb�>��4on�o�gl�!9<9�|5�� \={N���7{��	G��v��s�Y���c��H,�z�|��Ǖ���݈N]} �5��ں�Ga���M�l>:tO����.�ֲY�u-Pѝ(q��wf�߃�	�B5[�bJnn��0L��tݵ}Mń���z��������puج�Q�'.z����*ňW9�v���ƹ�sVlr��؝D�b�hɆ����Bs�Ic��.^�3��!��VV�$�m�+�+�_9�J�D�Z���$�W�b�%���5�K"Lt��s4-�ū��Á�G�!P_�(�T.������6��/�w��nu��â���b�}�aI;��X�V�ú)�5�閻��On�/�8t+0ked]mא�+3*$����m:�#�4D�j��Zo����N��[Y�C�ڛ�c�g6�t
_[M�%n���E�XX��lBk������e����㐸ݘ��
��"a$��V��(·�c{�5w�6)����Z�՚��M�m�@�%O�!�{%�԰9ʶhB��s�֮H�da��VWi$�Ȭ�1_t���T��.�L�0;NY���Ĉ.�B��{Y��1��]�׷Zsy��y����|���`�)X�QA�w������7���T3����z���w�ëJ��.�)C�)ܥ(���슋�Ϝ�+�t涷U�e��N�i�f&��i����J��C�jo���*���C��d�bQn�&6��m���[��̘e���e\�ڭ
||  �`�d���$b!� �A)Q���
2l��E3�4�"�Q�`�5D��cc��5bD�A���b���7wd�DX�]ݍ�LE\�X�#9q� c(�"����cE�H�d�h��RI%b.]�v��(�A�M4FL�#20��'7.��$D� cH������DH��c&0��JL�1%A��2m�rBe.LD��)��F��,��4�~?���������ln�3�}}B�{Z�\=�Z���-��܄6V6&ܕ��gt���/�)�U�0 U����`��~�>�>�>��OD7�h�b�����3�>?*/.��� ����kt����������['����gq�]���u���v��1{\���uU�r�����_uK��32��wծ�r��������sC���p�s/��Cu�����bn'���	H1�.~3��l�#j�{֧Q�\%]�v�G#c���'i��"9�F�ؕ����!�7�eqE�Ykm�_7�]�����j��&��gu�gBd3#�d���ܹ�ޝ��Żx�u���Iu4GLL5}DdR�c g���q���B�duÞ�19+i�z�������v��O���*z�����=)G�:��ҧ��W��rꆮ*�9P-r���ܢ�����˲�z��",�P�͚�n���J:��Χ�"��)�S2��n5U\*����/��lȆ*��N�0P�� -Ğ0xf�3��
�P;~��8���m:$����1��]G3|�-��n�Yb,�Wp���8o��&�\Kì��7+ՙ�~�7,k�����U����~t8/eg�O�)5�L�F�����*1��i7�)�DYBȬ��e�7���u:�VԞ��0�Ad=+����,�1�r��k���j|rl+�rT�<�uv.����9B�r�u�!m�('D}���VR���/�Ճ�2w^'��~S*�-�/��L��O
�2�{���gf܍-F��:Kz^z�+G�h�Jދ���x(v���)[���K���s�t��x��*���E�������n���`᧾DfH�U��������@Ĺ�[,@so&��l{�\�K�3&����'ւ�TQ��q�#PV:J�ōg���_V���S&،5xZ��Kv��"(Ƹ��|r5����3~�s��z�ѷ�-N��RA�u�,b��&Δ��L�(4�n�2��~Z�azR1��1ÕZ���@- � �����9.���xv\yǢf��ٕ"���]�(5���A�e��n��r�S�v�|{*QVCcX�����!�R<�͏#�B�1жHꂸ蚎I�f5b�e[�W�9�d�g�9�'/���P�rX�� |�Q�=�
�b��
���AcQ�HA�;�bx�c��J�X�Y�rF���*�I����mR���>&�3��g��������.Hr2��\4	qd�����H��\|㫫�Ų��z����3<���la�8���}I�T�gYcdB�U���kwh8��4�,K�Y�:a�Xɬ�J�µh�6����XX�Nu�X�S�8�M���v4�G[���]��>�����Ԓ���8�SED�U��S��!� ��ȑ_�1� \s~�i�dR�j�����-�qup�\�9�L\'�l��΂� :��d,s"��;+�?!��E�{��	����m���V��5���7I/�ݬ�uͺ� }����ں�9P1�S�N�
DT��o�u��k�����}	�_֌b1Q�Q�m��2`)��P�](p��T �N���VjK�
~1�UE�
X��58���j��`�M��1=��M�.�$qq{n޶�������Z-�u��>��P�8k��ܤ2�c�;o^�nV(�l�G�=��c����?�������<�����ͫ�G��ܞݨ릿��ySqu�t>p���W�dc�;ω�W�`mUwu�{��v��������C̹~�l�y�PHWxva߽��i���Rc+W<h�cmF;�ń,lF<���@!p������S:x(oPgL+8�@[�d�,1��m*���%��l�tb��1���}S�,�d�	wa�ۦ�MBO����;�>���ٲ(ì��h@+i�Ւ.X�=b`<y��KӾ�8�Ɏ*��z`wE䮣9^A���Qf��<)D��Z�gv1�iC�Y4hj��ƞ���M��-��eIL,�h��ў�����`��+��5R����z��+�?��ﾈ����,���Ҡ��|�	f�dU��jw�����_*�Rw�_�3�rV�'0�z��\�Z(T��ż�q!�I�<�͍���K��,��*��x4ӛe�R��>�bw�~�;�0�U�tݼ�3������F~'`%q]F(� �~34`�߭T¨�=<4��|\U,��S��E[�:�)�n�f��j����bX2Q���cͥC݄�6�4�{��@u��i\M�.���.�A��@O.�T#!OI��P�%���v�V�2^�T������r3�`gy���uB��5&�HP���P��9C�q_	�� @Y�zz(�S�j#�m���_�_�W�ɓV���U>�/����sq�6�̽���u	�1�}�����ю�u�-ՎuQxb/�(i1Q��Ԗ6�[vV�8L���{���8��c�t_v�Y�l�zk��8��?,�1�O��g��<�a��5��ucB�`�\�bڪ��r ����o���z��'�v��u�~��j���m��5�Gh�}�3����ܐd>2�F��򢳣�0tJV�P&�ʆ�,�5��kr��v�X���**@��׻Z�z,�N.��|#iSO�]��i��/�����D��3��l�1u��J��rH0�R�XN���gp����pa�W�UW�}v�im�UB��=�f�3j�%4�]7�9L�=�v��,V��0y?7c7���R>�-���c-k����o����ڥ�ێ�l�|s��/��\M�^�[�{`���J NP�]��*�!��-Vh��U�Boʯ��]Y.�ˍR탎[=�"�gR��#*R���|l�iϽ\��tn�Y�6����0����F��G�$-�2��	�ˎ���.+PL>r�;=}A�0ڴq�|�L�����{"��UѭW��t� �h�DT��S����7rw�r��5�����r��2���
\c!���*��eLm�
����Q?(R�'������*oJ	����O�7�0���7u�9��b���R�ρ	H0z6z�L���zs���z�שIT����+r\lw��w����֋�)V�N�$.)���f�p�I�)ډ �����i��χgAU��=�xm24&C1�8jrp�����$��D-�|��ĩ��) W�����u\LҘc�s�b��Q���.�����==5ҼV<��+z����1to4�^�^��6��"��l�7������X�ww(�^U%&��͆��㇏Mn���=�0�<w�v�tf"P�1��̶�ivn[��TL�=��+iVve�i�T%T�)��wCfK�����6qP\2�j�Teu��[�{�興�q�N�*r0�:b7�'wK&�&��G�C�iv�Cj�xfX��d\�f�����iJ��(Q�wUɸiyDj�<������K�rR��e^�>>tI��:��:�����.7-�vi������B��d� ��Ğ1D��g^���s8������4A�˨l�o.�a���b0KUP��9S��]����s�p�P�s�3�-�Ę�u{X��l�F�L�t�vK�{	�r(���q����V��^��QoY��ھ�>6.A��ځ5a�Æ�j߅�LV���o�~�]�{^�g�_����{?x�>p!X����L¾��Fm1_C���H𩸫�Q;<%�^�}+;���uᙓ���,K��є �S�͌���n���]��]�|�AXҮ�t5�蕣}��Fnov*��.1���>���b}���W�|}q}�G����yy1��yJOꔋ�龳z�6���|�&r��#t����9��,,/JF5C��D�6p�=m
�����%o9N�L~����N�@(�^Z�=r.;����w&�@�EA�LK��fd���v�m�����-�zeufp5qh��B���S(]�\�}Q���ʏ9@��mw.��p����~2��<K��o+��Kc��R�ׯlȵ�--}g��UW��ޒϯO?zm$�
/���ڎQg�A	�'��E"�;0��U^u����֕=�첨�Vg�bE�u�u����7�T�*P�Q(4b�l��W_}��F
u��n���]M�Ť���d���QC��A���9���*��͖[����0���MLS�;��_���{̖���۪5�r5��x�V���Ҧpz�'���J����w�{C�<�?��C�KUb���u�s�y�@�p��W$��:n��;\c���uf.�C�V�gn�����[8���҆����i�& ��7rQ���7C�.�G}�^u�N���))���K�͛mP3?hVI%�������r����A�a�^z��X��r��E~)դ4��t�����>f1?[��E.ҭ�]�̫��I�b���_��n k��l$v��6�z�<��:�^5a1�o!�řׂ*��G3ZUj���n�W�P�~��}�M��b5��ӕU��'"9/(z9Ω�갭|��Ti���1��88�[�E�s���p���BX-����[X����9֢Lj�ڄ;6T��j�U���5�b�� .ľ�b[�t��w>c�E���)��aL�Sz��I\bO&=��n��MP�뻇/b��˼n����d��v���v��ވ�#菺��>�)�&�}s�M�g��W��^��K��s�db}��53�
!'ӝ3�^ʸ�[\�XQ%U�c@ծ�}z���;�V����E����u Z,���ɭñڧ�O�qP)�&���WTY�fÁ���ULe�v�湆;s�l��E���t���.%YbWc�)ر@Hd��]�Uh{�
�&Q�/�`���[���r�H�ɍhƶdN�cY�����	��b:vU���
���&�|����NH��sw��-�8�aʹ�+�S��}I�zϫ5v�<�Ҷ*�Y:�2��5"%Z0��=��

ǹ�����R׺ݚT$T�(?������9p��T1�{����#0N�J⫨��*�o1�qj�d�[�Ҋ��W+�Gm�U�8S��О�c `�i	˚���	/.�>ޙ��Ҥ��un9�|�-h�M�U	��9Z
ϝ *�U�\�� ;�������=�.De���aTS�sl�Yߣ�5�'�\9�E�ȕ�Η�>�0V3�!r�����pӠ�JÞW����n�/�ؾ���˽�f%]`����SG�=�4>�m��H�6~<W\��!�ѝ.���H�j31�S�
$BX:���%5��1������K���iR���QU�nR��:�Ds�[g�Uw�<v�	��5�w���sn�K��%�̫\϶������⠽��u�^'��5�n�e��΢��_�Ol��e� K�*}ټ�B�0z�8����#[��Uq����ٟI\v�v�u9�x\;<�ij�C���;��ˈ�c��Xb�S6����@��y�'����lG�v��,u�d卾sh��R�o/wy!��4K~�yJݝ��*�pз�]ʷ	�����܀���[Xh�T��� ���.��@�X\J�q[p�%+���o�]�r!��{r|��y���F�V�h�}��Ժ��X/�����+rg\�ꐌV˯���N�7��=�SmW���ry�_!�[�2[��g��?1[���oi�TU��}嵍h㪐��_-�Ps/:�EdhC)4媮�~p��>;�X|j'��.ۖ~��&>=5[�w��v�"��e/\g��s�w'�蹵xv�!��މ�1m�q
��*9$#Q
B��b5��v�N�&�#`�Cp�L�������Y��^t�Q��Rv(P�C��c��RUcOw=։՝�1�VNp^E�>�������vu��g��sa�o�dr����d\;���}��n��V쳓t�75V'd$V:6!��}���}�}�л϶x��Ia?��/r\Boj����p�KӺ��c��.�E_���n�*m�y�

4@�O�⁫���.�(՞��D��rDj7D�v�D��'U��.��҃о��#���� "��C����f��f&�i3p\ƈ��G��"�ǉ���x��. ���2
�yJ�o�zLҘc�=�/�0�rt���ηO#����W�Y�䊀c�/|�Uk��%']i�<N}%#�7_m�LJ��X���q�'�2_ ����]��.	��*��+w��;H{$G ��� �b9�\���v�Z��,�t��p��XK����
5%�b��CE�f��L �H]r���6h��t���nf��w�,�q�힕�Ve۲��{^)�@j��t'캄�,�c���E��#�UP�8�N��ed9�m��*?l����$B�u��d�l��et�G��N��)�e���gd�S�_ݮ�gwQ{G�ylٕ�@��ꇆ�j��i��Qx;7�k��Z�"��[t%�38`-kEޜ�/C��[�9� ��Y�7�k)9����d�)?�Z���VW�Π�hJ��zewV1:�e�3��K�x�r��[j��,0�-$���3D"�Y�W���K��&�`}��fL+�ر��ظ�7C�ndʼ�mu�o�zH�p�W[�ƺ�k�1�H�̻dCQ�.5nO��;�Z����$��N���`�O��]奡қ~��ڗnw
wT�%���=�۝�ŗζ ֢̀�x{��_1Vs�mm������̭:�8��\���e�N���%���%��d�6��f�|h�Nʦ��K�q�	Xղpv�*�f��<%$(��M��XJ<��I�h��i�ad��'5#��*���ɀ#ڝYt������v��0�T�]�ݐ(��q�J���jE���L&�2J����{�pL�.TN�n��e�}ݤS��vi��m���&��(�9�����i��Xҁ�v���[i\�)hKŌQ�� �qb8�St9)�!@������hw>V�C-/�2Wvл�n�*߂�E9w�=�T��As�z��+^R�z�,O�f��u�e*�Ĕ�T�A�)��N��j܃U�q`�k�N�P�6�j�8��A���m���D�r	� V�|N�V��4���� ��ݻ�6��j���sR�2�����u�x�TU���R��ɵw'!V-�m��\(Ӻ�o^6�].A�F�)̗؅-���v�Qn�֒q���� '�K{Xtt+o��5�Y]EvV���yP��O5|�̝W1���؅�TI]�|�ep"nYj*���t�9X�kj��(�-�uֺ\0���`9ܾ��D�:�ǖ'{����O���-�2����9$yu��d�(:�F.9-�X٫�x��3Pwb����
v�f�g{��I.O��>�Q�t����H�f����N���+F��:�������/�V��r��T�Y��x:��bnM��զm�
�ڽ��oa�h� ��lA��5	�G`e�V/xa:�����S�̓�`fQ��]�O�N�Z7ee����:���ڮ�:b��t�E]AS��:��=i����2���J2Y<����Lʛ�G q��M���̐,-X
����*�p'Fl]k=ݣ�3Kz!D�X��]��`E��c%d�ao��rU!vW���6�:no\�F�*����݋���
TmC��_��m�vAՄAeE]�;��t<�AKv���+,'�`�Gr鹖�p���;�X;PZw��W����v>}�#��}�ռ���fЫ�Zq�>�לG'y�9T��
����,�,��E%��;:�^�#��+"�[�F��Q���#ٕ E� ��|��Y4�[��	J1ݻI˖M���m3RS!,2I�1��庁s�i#0$L�j+����7+�L3 0*&	I2�A�!RPi˃����.r�	���wWE����&��#����3Q�Q��̓��k�r"@&����Y�)(�9�wsN�0TF��gn�;����ݺ��"lV��;����6)Ί�r�awv's�����w`��3ۜH(����U���
�5F���}m����QkN�32���%�r�ziN�����:�M���GN�}���+X��Y<�pWhپ�p[iH��G�G�:M�^@R��c����ry�T�*xh:��W��\"���-*�w��eq}�u2��رT�($Ԯ�1 T[��_ԧ������{r�_قR7b�i0���up�!l�.���)� ʀ&��t��8��9Z��GȧLr���]W�a�ܢt����O
�3���G��zԜ��^M�#��?.&��v���/ґ�u,1Q
�o����;�z2f��`��$	�g��O�����"�
�O�"�!���O0�Wu<R�[��S��q=G��!�$�u#>*P�W��F4X�+���N�0�PV>wyY�؝��O,��%"�٘�L��PӢ�D<���S�h�g��0���aT�:G��ܮ[ԜTș��(o-=�*_���b&ʓb
�s�D�}t<9:�J��`��+�_�]pY�>�O��B+��`�N����#b ������W[]��z�=��V^����f�Cv��P�W�3Z�S�@F�C ��a��
�P�cn�#8�;l�DO����yɻ���h�趴:��2�v���p��%��g�
� �G�>�U�uE�h���&Jj�Hb�36m#'�Sg�ƥJ/8<���e`��6��z�U�vxu�[X���I�'aN+؍��Zx�bi�E&I�VK���g;��}_UUZ�E���v80D���*��#j��MF���H���dVN�E�ڀ���l�eR��EY�[�9�Ι�D��V3,F��A����\�3Q������A�7��\CSYԫ�&�6�������p��gjp�q���=����J5vzU�|�
j�]��;��:�����m���׬Ӻ�y.�1r�������eR5�ڷ\��
�as��wh�Y� ����{�D����䍄���p�hۍyQ�Vj�����-ߍ矎�G�^F�޻9�uv)z�C(g����>O9�2�h��:s�[�����z��� �`�X��+]��Sn�]�;/�8:��w�E��l8�	U1������ϥ��<� �ev�U��({r�<v�?��"~%n*���XJ0ň�Tmr����n[)�8����S(��~��6Fӿy�b��S�
˼�2z��5��eU�)�l�J�z}�t�ф��Ց/5gS���9��/��9��p��u.da7AZ0���T�jr����ܦ�YN��6e��v`�d]�֚�.��3w�.��l��ݎ��W�����v�
���P�$�z�M�2:ɎqǀD:/��C�{R�9X�Pػ2���9�zF��W*^������:�u��f��`훥8�M���G�}�P�n1�I'2xH�w&����{N��� �n�C�������#$��*���	��q�$+������}�5�d��(��Z�λ�'��������d'.j@!���U{\Y�h��GYV��=g~%��
~c�M+����s7�������HS�g��	��y�/���W�Y=�Cg$��8s����*wa!3�@Vw�5�B}PŹ�E�N�'�S�{�e���c�;k@O����q���ӗ��!�#����܁҆�$�/+F&���i䵚�Ѣ�ra�n�ˍ���`<�R�_�x��t�hƛ��UeE��%��̉�}�R��zB�w0Z٢P�]0�t$�G<���9R�p'�ܕ�o�ǿ{N$+�2Wi��k��f�EW;�N�������G^ *����}�mv#g�]�L��_γԎ>��N��`q܄9���t�[��*��Ōٻ��7'0'�ʸa����C�$w ,�޼��`_��3x�U/T4R�-��+;�b�xoϳ�nOo��)@�����X�>�vx31��`В��Bd�y�TD���}J�k*Q��ʊ�E��v�{�|s�/��M:�/�Iru�{ma:��E۵��A�TӹG���\/hF
��49��N���'���$��rW�]��u�?��ꏣ��ޮ�Q}Y胘cGQ#,��-X!��΢vzUZY�R���O�^^v��#:��h�=�﫹�r�d4h�>��뻟��ma�
��K\�9>o�UQW�Q+�+ƴvG�M��l��ו��;aa�G��>;�[���M��[^?mѭ�^ө�� ��� ���uq!ʺ�{�n�P.ے����xJԸX����q4�c�cd�HU}-�&��е@�q�Ֆ��J5�B��沀��imDp���ۇ�"�z
����1pz�QG(��'C�;�&mv�`�C���_Ġ0�}=?L�Qr�����))�����$i�����,b���l�Z�*t���AY�.
��/�v������L�L�ʄ��L-��ӝO�:(B)8U�r�:����'эR��IO�xX;dq�0vȑia��V�3��]�P�R�]9U��o�R�j�|;�R�W���=>Q����ҧ��\���{I�;�AF8��*�@�Cn"�G'V�C�A���P�ٮ�_����D���~� ���t�s�U׍Q*�R6��zw)L 6�S�v�sZw���c�h�U�]�5z�ls`T1u|�F.}�#R��a��ym�Ů�s�����2��auu�Q:���͜�v�U�x٭���OsOw&����r��@ܱ��`�E;qf�-�.I��6qut�\D}��}r�%�jS�W#����Y��_�L`J���:L1O��sr �@�#���I��B��+s�{����m�S{P����N�g�+�'LjUR��c>N��}|4���w#!>�T ��?tL1����D�b��X�k)U���J}{S�~u��O8�4-ך��R��q�]�'�z~m�n�Fɫ�xh���i��U��|E�n��5��U��4�l�����Z���{�x;���y�/�+j{�
���EQ;<%U�^�d�u����������V�O�����-�zbQ���{|;9��1y�R7&,F��&D�[�/u	�coh��,�b�}i}���ER�z��m}[���ڏ��{��\��Aj#�;_�է�]f�8j�Qz�����2�*�����_�v{��s,`�]ֆ�S�S9�:�XS�R�Q_. ����b)T1�Ȭ�ċ�\�\<E�g>!���:���T�']5�����Fv�8/*YY �O�P�����A�\=ƥv"5�ӁY�]��[�t�{뷦��*eN�)����rV�tN�2.�ˆ��~�"���nC˔�ﮎv�vQy�9�D7%WW�gnS�{P���˵΃]����Z�t��A��!(��mJ���4`wM�(��1�VQC�V�5tvT�{S-��SW��<�����������yM��[zct)�c�8GB�Txz�|`��OQ�y�ÅL1q�f���C]�i��|���Pd��|�_�~�|87��K�F'9g蘅h�u� �:`�:\M#]��׷�Z�ղ�>T7��i����1��r���#�"Z�����:U_����ʴT'���{�LR�?IF�V��9G!���5EBI���q� +Ώ ��,�&�mC9��7��!�u~�R���|핂�>�&��.��1��)"2�;�7�j�h�l�݋�_�qNtכKv�� z�g(f�]W��/��X��Q�f>i
[�o�}oˎh`�6'5f�Ɣ��~^�㣢ڠ��R�K�`��Ȼ-j��Mm��)2bT�mN��-ԕ	����t:-�����a�]=h��.������ۥ��;޳'Ou�E��ϓ�p]�0*;����P5ٚ:�Ͱ5z�?m�~]K��-/����z�׹+ۃk�
V;G�8��$�W�oƷC��OMC�+2ig�FAcC�x��Q_m�r-�1�kfj�I^�[cn8^դ���>�	�4f��#.�f�s]NOAud��,D�\<q�i!<b�e�m��ZL�6FL���m/D}�D&7m+.�#犰��Jo�՜u�F�+܎��wt�]�~^y�1��+���x�<��iP�A�ڕ���<��O:��J�F�WP���}�T��ò{�y�b5���0�<�u,���P�a~�Klܙ�\��P*�N�7ڻ��SMl@��N�Q�_D�;�;:L���y�5�NRy��"��Qͥq�n�=-�v:ܫ�l$�u�\��*��/С�kg�RS����ջ��.�PS=A��wj�?'.T��o@O�Xyn�b���t�"���T�H�Wّ��Bi/y�z:ἅM�4yy�kF�>��[Ě��k�^�$[F���[�	��[p���=�QbX�κ��j�5J�n�[�#z���[
è�� �D�m��+��,{c�OK��%�3f��S�9�	8�4�J�Y��%�q������Uf��)�y맅sś+�Ʋ�g4S0��v
t(�d�jﱐ$�$]`�8��3 GF
R�N�1�/M�[Yև*�C9]]n�y�cJ�(���������Ou�|��w�)d�n�Ԫs����F�N%���"��/a��(p>�]I��`-����dtk��_�3��R�[N֋Ǌ(�9?�n�����m�J��k��Ή�
~�dÂ�B�[�k�zvg���K~ұm/y���ή����`�b��'S?Pm�3F�O@F����̪�N)��v�R��>�=�޽��Y�RM��W�c�oQ���iy�ݿ����-���7���o:�^vp*�b7j�Z�r�h����[������E��
��1Z�Y�薦v��ـ/)B��-Fe�w��X�{��?��ʴ���<�ȕ�,O{�I�v+#�D�#����*��Wz����ik.�ݸ���*�]Ef)A"_p�%m��=R��drѝ��.����0�cI���q��wz�H��wY����R��X�F)TK�K�Z疴t��!>�Lv�+�y3&�,�����:�1���ڮGi���zAq�����	ӹ�$��lս����] �̋���Kթ:�Z}�ח�%[�J	
��.v�R����=A��!\�r}�I��hM�6�6�,wu8E)�ԁ8�Nt=����{��s����|?�>�>9v��p���]q���*��	h���'����S[�I���u�W48�UON0�BR��Y錈K��s���>��#M�c�a^�+��LeS���WS�o��!;0��m�A��l&�8��w:��c�|��K�[]�\�%G��I�z��9����_bܐ*I]��Ռ�һ�]��ǝ��-i�x�=�������mC�St�"�E�f5�kF%;��upTl	�w��5Qy�����a>�|���SS���W�R8UoC�J�y��<��q�_����F/i��Q1�Mŵ�`�އ�x�����f����u���X{n+��Ψ�s���12��^�t�;Ǆ� ���f��|�חeG���}�?����\��܋e�W8������{�(��^�gV�[v�*-��*�a���:����A�{g)�囯s��ylY���}��N�+���Pp�a$HӺ�E������}�vew��L�'^F=g����IG�Z͹}�]n:V�䁄�	��y���|r�����u�0c$�Y#X��;��Wq.�{{;��WYE]a�݅<����)���}_SqN�*ϽW�?Rz��Ц�Jw8�<�}����]7�x�3�	�¸Ћw���7Cl�=��9�����ל���G���ȇon� {����ks^5���[/�v�Pz`�k���|�D_+
�>u�������y �6�,�{k(4%c��n��B連z�̄�Zj�h� A���YKv��m*�����ڭ�Ɋt��v�_��	L.����4�6j��Z�)w�/'������}#k����U,�+�=p!v��9�'�n,�ۚ�5��fNۙq�e�n�4�ྦྷl��oaT[������l���:gW_
�Y.DT�0��h2�&���x+ԙڅ�[������z8$#UF�cX�qi����xPe�Q��x:i�X��[IQ�\�Kt.���˗�Me��E����.�;Zc���4�����8�����3mZĆ��Uc�BT�h#o鏗˯��tq���nwTMC��δ�=�sYu
�%�K����6�����wOZljZ���լT�YK�e�����b!�]ɂ���ۺ�f�8��՛�7A��o)�^�]���%�)o��j��`n������+z���5&3�۴��-�ÚǛ,#|ys��$W]�G �g4k`(<$CI#�v,�Z�)nK��PAshZ�j�OOc�r$���C�e�:�5X�Y��	l��ܷ�踃O�:�E�]�%p�G�E)�K]�Ϋ�U��.����)��ݐ]>׳U"[;#ꎝ;r�����:���:�X�>늗k��g3*ܹ;6���;�Sb�ǭXA�Š��JPkQm�����I���d���k�R�����;(ɫ]�LCHeH-T=W#9�K
+{�h�Brk 5gL]�� �cB��7|y8���Ku(�%y�V3��ξ�U��o\����91tٻ�2*�'֩�r�cU��v���뱳�=x݀�&����[�t���老^�ې���Qi�b�F�c��̫��t �j�7�]wM��:��gl�9q&���N�Q/�YF��9���WK{��8-ӊ�qeF�nh�Oz�a�U�n���v�]Ib��w]�����(gjsx�Ik�H'(2Z�IS%;����:H~�(<�o���ܛ˲۽�m�V��욱Ւn� 6�\�Wf�Z;y��#n����:�]x�}�U��8[�7�tT�Kt�;�v�G�6�S�=��.e;��77���#6�����.��t�����5sE:$�{9�gpr�Ш(�w�1F����鼺�WFޒ��`��bʺ���Q�����AA�q�Zb�T螚0�vl�v����#M�*;�:����+�ἡ	�j�.����T�ں�r�m�i��O��R�\xo ��7�Gw֡�`Z�.Zβ{صI�[��:�l��:Cs@kO�I�m��olU�Ǣ�b�������IF ����\"�T*;��)L�K�~4���	���volB�ڻVۨ��͜�<���)��3F��%�S2���򃤥���7GD����1#������4�����&�<��i�۹��|���Ҥz��h�F�b���Pm[�%��� �i�����8��-�ڏjC�G2u��kE�<ݽ"u���*]���T�7�W7�ʕ6�#oE�8��QF�l(��A�ՋC3v���#R�]bi 4�ڴS�&U۶�o��[|v��v���V�8�R QF��'�H��i�/�B3��w�mH.Å�J�n!��W*;�"�x4b����?���iH�gu#�@�K�w�z���&�V=ڵ�z�o���l�#͑�3`���4\���#>��_K�[l�\Yq�훂��cVt��'���shv�"t�6~�y+��M;Y2��9��Qw��[ދ�O0C,*�.�oK��)e��:��~�T.����m˺�B�-��Ewu�9ۄ��� ��W.�X�5�:+���-���ȷ,$n�ܹ�d��Pk����sF܊-�t�� �r#��3��r�鮑��u�6]ۜ��w"ዝ���\��ƺ]�	��DPWL������gv.�$(��+r建6*B��Ԙ�66-ssű�ڋ��&�N�n�ѹnn����;�J拤��t�s���wr�����7;���u�b1t�f[%ˮ뻫�5���Η)wW�]�M�&ܹ�+��]�r�ww��]�������5.���뻱�X ޓ2�TO�]4��� ๻���aW�u|�f�'��k!::��c
��E`5 ��8q��]g2�3��}�g����S���_�I��u\��:���ttV�Ί]�����P�7M��j�QXtK��?s��t���g�wF�Õ��A]�qX�k�^����!�M�����Q�U'�WR溜G�f�ϥ��7��i*��m��sE�gL���w�����P�_n��u�2#��g�x�?Tї^VM�n��G�#B�A����{����[�U*��7��6�gG[R'�A�y��&(�s��7n5���ܕ+Z����O:��J�;D�d"^���`����Mf���e70�����W_��Ʋ�~��*/���N��K�u�2�q.0͊���Ŭz;3�{P�����[_(S?�6��3��vewO"�!'�|�rY���\饐�]��v��u�ʱ�W:8�stc(�ޒ����I�����@\���kGJ�(��q	��3a�)���䎙뫳`�9`t��<�3yr�z�*h�gN4|6��7�_�'�{ꗱW��H)W����ChxE�Q�,z�W.0�AL�oL{w���H���tVE���6T�;Wc���X���aL��0>������@m�}�*�o#|��1'[�bj���m�Nu����Ss���a���z7�Ȯ��-wave�N�!��:���dTH�����[�WnW!��1�liC`��0��+s.y�VTrga�B(����j��g%�uO�e��]�K���*�n2�O'�U_[�m��gV�.�5ϰ Ը��9BL�CP�9y]@����`���/3��s���tV��.�����Y��RT]CRU6��}�)�B8DƸu�[���������J��s/�}��篴��ە2�t'-M�7��p����y�2S��G�G�W��ŵAq�ϴ�U�'��/TvJ��OW������_M�] ���j6}<�f��и��4�n���]��6{c�{����&�W����u�}s��O�Ky%�����죉TY�X���4�e�z*����U=J	'u����襛P�-�g�"�wCs�Ti�u�}MH�_�s�z0�y�3n)X��:�V4ݧO�#gF\#Y��Ĵk�����E�JSh8�R�]�he�W$�Lf��*U��y ��.5*:�6���u�o�:bB�k�k���w�ݪ��J"��Q痺d.�mX=��'����YS����9�R�ʽ���|w�����*oj:V-U^OЪ(z@�e^K�a\��ٶ�J'!���5���I�K�q�����[x��ODP�p�R��6'�V]L��t��?K\*����GM'��M��[��8���Y�:sY�.�fk�آ������%#!*�3�K�}k�\-4��AO����M��oUm�e8%��d�N��N\��	mJ~���	��]�qڛ���S^�(|`�}Yc�rK�/��v���;+etwS��3��Ew.~��Jͅ�Z�(�W�q��|쾦�s=�yI�U�yh��t_ek�0:����K�v(M�����ՙ�VRTr���pʇ�yl;By����.sa�/a$�N3Oo-m��ǎj!v��J��F�Cn\)�w<����Rn�8�����!�@wC�m��.Ҽ�󱔏{g#���SF����j�{��`��͜�j�%\�N�)i���2b�����n�SRj��	D�EW�G6�Ie7z]�X�3Y7������4%eu�'eRo�fTz C��	g+�$:���!����eM�/���Y��ɜ�J����>|���V�kQ�Vp9k� L�we;�f��{ЖY��8��ob�r���^�=������H^�2����^,mW��mOU��=��qM��roo�ɮ<���ԃ���=)�?z���v{��?(6� �y���CY��0ȭl,��I+�j-=N�����m�k�~{�j�wL���V�ӣ�\��i�Y��n���,�J�=���gUmƦ��}�����̉_��ڌ��4�p�q�T���T\N�Qg���h��ժ�Jyv��q���-�L�����h��Pttk*
L?����sgz{:�&; �b�A�'A���v�1-f[��R��BS67��s	p�Me�v3	��������Դ�!ƥO$�9�5��G)��}=;*+�v��r���MV�3����뷭T[H�������򊢧z B�&�D��Z�`�3S���b�[��f,�Y�U��q�/0[�x�伂�sj���ڔv��`���;�;|�B�oGK�vs��S�V���΄�t8��]�=�{�%�ro/�pw�wq�<k��iv �[�9AK�g���"х'��G��
op�ɒ_�S'����2�ri��_Sp͠��R)�oӚQ&�=ήr��;��!�}�������9���V�8��w�z�M<dsҳ�s*�P��v�'�dK�xT�T�kM<3�]r�J�*�Ӯ`��jU�*���]�h�Gkwas�3r���X`������1`=�A1�7�B&Q|�ߪ�w���]0gǝZک�zY�}W��~��¶���.Ԏ��o<l�O��b�\W�I�58�Ϲ��������:/��T'���%foy��nq��^NV8�Q��c��	��mn�k�8�ئ�҃a��M򖹜���\.�8�ss����Db�U�������x�������艊ty�M��;�nA���"��}qո�Q��.yAKd���2����x�7 e�ۈ�ͦ�n�1�T&��:�k���K'�������Ҷ�	������w�4��=��Rյ�������&����+c���QX�e�/r���L9̰]=�i��ǺR�e�K�S��kxGd	�}��
�v;\GKG7��Eq�7�}{|�;y9]$���z�b�/�oM��׀[�GY����J�s��8>\��x	��՗ۇݐ��)��]�u�A郱��TN����UN��n��4r�M�o���Y=�m���4���+n���-ӎ8CHޢiY�zG����z�����V���4����ҿ�ݸz��9n�k�"���5���t^K�;{\؎�.�ن���w�W�6�O��N��Sٷ��[�Aٮ'�����MqLBY_Jk�b�vf_�S��5�}��yW>���V��\�X�a�z㟲ʲ���Wh���ne��8+��g�SūV�qܡ�6f�o6K\��*�zR�<�J=�e���{f���#罷5{��\dҪ��q	Ѻ���&��|VC���'�l�Y}�itM����u��h�-�/1��jV]��Snt%-�B������Mlsy�����È�i��_^gU��נ�Z���n�+Fz�;ѝ'�����WR�0ޡ0�ݚ�+�M*v�RSs �.�}�V�%���}V�"'Z6ם-^� ����F�	������*ܨ-*]j3H���`��,��%�5��O2�VR������q�K�j�,h�ȍ�8r��Ш��^ 2�T�s4u�sueq�;� @�Ӯ;`+� ⺋z��X��]�S�w����r�qtrqLz��>�7�����z����<U�����:�ю�8���s����X�%U��fc�m7��/ �Kj�{��.TB��g�\e����6h�V8\ثm��6��Œ�/�tsk�<tY�����J{2�5%Щ9N0�w<� �x[�m>܊oB�������Y���;'�`v��E.'bV��4�Rw���iM�C�]��O��������F�LP7�N�ۊ �Ŗ:7�%A��W�|�b���p]�����P��s��$	ۻx�5�̘��er���ՈJ`l$Y��
���r7zkz@w+r��s�W�)�%�^����՗3ˊ����P��tk�Sԇ{d�5��E��գ�BQ�)v��AZ��w���k�Ȋ�J讧��6�������]��
CA;��sA_F������Z+�}S%|gq��n�_x0v����J�T��_p95&ֻ���S@0Z�z�<��}���͋��9˷@�]X\GJׂͽ�#�iM���nn[x�.d�ȴ��I�U��q[��0½|�>���o��N�����/aXu��,𢷜�w�$�x��WΧ���^2�Ŋ�y������N�
p�@ŀ������g
\iC�	�/-�ݯ�3��zg9��V*������[W�&�>���V|��=W�9�=�E.�+���w�q>�^^��Wi����
�u���r���z���eDw__����}��Y�SP"�5�"���`W�N�q���JF6��V���t=�\v�)/W=o::���N����ަ�Mk��>����y=~Pj�������)���輮�1����]Po�OuY�X�F�[q�ثm��,���e=��,����7dn4�r3��{�/�U�U��\j��M�4���>uUv���H&(�Kyث����B��=%���P�d�ҵti^�^�.@E�m���@��޽�ݱZz��E�0�3������ѯhL�0婀�pu�!�ھ�VLr�p�\�e\��m�}o�ʘ{s�q�⋻�wg��0hO�+7�S֖�U|���l֥b�q�mk���������+�r]�s�!�x�d�C�jz�WQY����v5�J�I���JԎ%�ͅCw���ӓ��@���>��t[��9��YJ�BScx�p૶8�A[-r}D��O��
b�i��_>���Ɋt�:r�\�jU33W�g�B�L�v]\تܻ��-j��h������z��tM:���y*g�T�D7�,����@SY�W�瀭θ;s#�O���6+�s{ƪ�6��-���I� <�!�J{��0�~��ɨ�O���z�VcM5䒨� oR*5��CFxyT�����KCܯ9�*�V��r�l��k�E�{۬���CB�^i�����
f�+!�Y}��T^buR�C�|��q�塓�ͭ�1���ڮ��qWkp:��;��3h*�+�bi�;�����V�VI��aL�zíJ&#z���Wq��'�*5�ܛ���l(��=՘�{͸7o2����7�\Ħ���2���˻�.��+"��xi���&���1�Y���g��;��$.x��;zᕋ�_������=r�ņ��u=�淪�[�p�ٕ*��C�5ҙy��ᨻwTn�T[/2�M�f��kd��!�k*.��t���B[���j�^ߨ����Z�ޞ�j.ϣ�j:�WW�Ta������#���<r�.�>����3�n��ݾ%�i��7����}�a�e�W���MŴ<m�Oa��,��eV
��»�#�L���Kw�[��k��绋^A¨K�mgP��<�L!o9�����팄ѷY.�i\akouC���웅�uDd�����غۆ�Ue���T������t'δ�š�6�+�'B��뭇t���YCq�� ��N���e��:i=<�Jݷ���d�xk�3O'r$�F�J���@�遰�D��ß���g�;��7����J�m��$�Yf9�w]5	ʕb�0�q���mގm4����pmۮBzf�a�q���uLe���O(���O+�Bs����޻�|�'
�NY����K�XuxV\���P�θ"1��c��C5��e�\�FXp��*�H^���K�<���ήo	5܎�՟-���4;C��[�ȣ�;'�����h��J���K'4�5X������<�7sH�bVl��N
�����͙X�n+�̋.�h�i,B�F&0u^�]�vg8�G�1�{�M%MQ\쬫΍M���C��Is�ro	��i�|��U����G����u.1y�`M"+z�QW�z�����a�����b�'��9ʀ|��rM�9J�Y��ɐ���+w��O+�c�T��(fWu����e�����V�7SM�˛�/tzJW1��e�Qp���+kg
�5�ʳ�>��˿��Y]�p��X��rZѯ��!��Q��W*8����L��r�wm{vC�{�N����.�=Z;[ǷhSn�8�� ]�U����v<�sE�Ʒ�4����a���d��m�vj�*J�}˻�N���E���
V4z�Ț�
$��o(��8E
��RV����3ޝ�?e�9/C�w�H�i��D�eCV��)�g��\�1g�˼K�MC��nU�y*�F�Rw�vf���S+�6kw�ز��5'H՜Qr�f�MP8�g��X:������i�j�]o)�U��\���MNҜsu�ǚE��:x� �6���'����9�4�
9e��f8�yrK鷳�Dr�~�N�|z��$��x�l�Boc7�s���+T�G jw8���g�p�[Z�=�{B����odņ���p^_X���s%e��l���
�g��o��KV��,e���n�¯$�a��T2Cl��e��n)-wdt�qV�Zl�w�j0z�݃r��E5�[�&���Ŵ,�Y�zeuw+iU��QZ�Pj�1]׌8��}��hV:Vñ�V2�9�1��t�@Z�6f���Yf�".]b�uY/������$��q]�R�÷.�Hf��]}��)c:L�`�z�a7�PZ�)�::��R��i�n��USF�4Y��24�Dg�ױV�|���*hJ�=(t&o]��d���`䝴7�W*!l�܇lvi��J�GS��VW
�)!f�c9;���i����:��
�ǌ���[�}���"4�KJV�5y�9�H��
TZX��b�f_/�V�n��-unf����o�S��t����o
��f>fΤk2��N���ս���GE(W5�ܥ �a\k^]M�'ǆշ�ƚ�;�A����𭾻o��ڄu)H�P�n�Z�1.�}Ad٬�[�xr���׃��E!�I��JM6 6d{@8.�»͝��ޖ�+\�eqd8�+�d$�\�*[�J����b����S$�&:�6�cܺĺ�VSY��g�a�'R<ұ)�2C���S�����P�:536{��� ��NU����+ u4�lw��t�j��l�<]{ku�JRNt�ש�Y����ۡ
*�ge�E�70_K��`X7���ց�;g}�=�q�s�6���cWMs������9sn�7.5r����u�s��tW1���&���9\�;�v�V1���ۗK%�sI����9���s��r�V4k��wv�jw7wF�\їu9�m\��#Nq�s���F�!��W+���cd���1�\�w[�7#��u݊�Q��\�n$Tȩ΋r��r�)\��q�$��"��c��\��h4�]�f���AIʹ�̒D]�@��CwWFM�2���78��h��\2(nB�u�vrT�u�%�����7��tN]Ηww\�'w٘)�;u�;��:%���K�]��w\c��ͺ꾰(X��QQ�����`�|�Q�y�;C�M��E��;$\��թ���g�=)N6��9\�Z��v1��ڥ���'���P�u��͌'$����A]P���l�*-�a��W�]L��;��j\��X��5���L�j�p�@sg�b�G�j��� ۙj&�<;�hݫ��r��ԹXʍ:J�����D�<�Q�̖"�RTl�-���f���q�}y����@נ�(ޖ�Iz.5Ƭ��lT�����n�e�.C�&�mOU��E����{�n(۞�>6�1؉X�a��|��r�G��Jx���8��}7~]Kޝz+V6eA��s�SFvm
��KԺz�����6����jJ�m������]�Ԧ���s�*��d5����E��r�mCx�]����ty@}k�[�5�]Д�;ŕq�<�)��7ɭϩ�*��=/���zv��fq�����������mG��*��;��|�KYoGn�6�q�ñe	�Y5Η���;d��Q��e%����!t_.�Ա3�����r�G�����k�P"v�J�Y�Ơ=�Ճ�N`�����Ңa�F;}{�k->V�a�Y�z؍�ۏ��<���<��r?rL�ڝ��2��w/���VfJ��rv�ݚW_Vp�� ��3#YQr�
��kss�"��h�J�b��늢6��V��b�Y��p:�V#����\�@K�DZ����]P��V���I`wW�g)%���!�ڭ�ɏ��4��_%��7���2N��7�W��;�w��=Mz61��J�:k��s�[��e8��V�{��tI;s#U�k�]e�;f��������+�<*�嚾	Z�Ƚh�Z��W����ov������$��6�voi���M}���`����[/��gT}oL��5��%E�G9
�l�R�>L���&p�2��L;�^^OUõEnQ�u��n�k�p�6:��
�&o�5C��x�+jz-�6��H����|���eA�u~�xn*�f<s��F)�>�QCx��5���s��G8��zk��es��E�Q�n��0L��3�;{�5����꾧t-L'���1�Ǘ��];8ͩ  W�rݧ�<�4lu�CS��WV$��G �mo,��d�9�P�xsJ���»�i�ξRc}t�]�Ÿt4D�m��F�-���H���+�+�j���ٌ����a��X�՘�>]2<3&:	9��g*8Ū/{k������ώc��33RN� Z���ʽq9s��uY�X��9�������E,چ�uͱ=Ur7Q�+���/l$ȉno�Xűe򳼯��ʋi���Kmьaf�S�ު'U�o\.���w�ה%�@��}�ݴD�4�{^s�o��HL�c�ݻ��?U'ޑ}^>{]�8��9ڃ�v5Ԩ2��_%�XGi�Ѳ0����Q�F���/��J㔶��Żxֳ-��|!(��,���b�L�y�������<�?�w��z:iv�M$�v�x-|������+����l{-L��8P�ojN$��`�9Sʲ�v���i��u���7q<�yv���^f��-�O�R��!��LW	Z�0�����}�ྦྷl�h��OdE�b���.��8ޱ0�\��~0�~�D�ɨ��n,��������	߫<1bs���u$
��M�\��ˮ�y�"<,:f9��C��T'J�h�v5fw��^�kSzw*^8��2j*:��{X�+���Vl(�g:��5���(�TRpV�x�>���!���3�q��	�[<��KolS�1�˅������l96W�Uu�#yM�z��`8i���}��^Z�2�V��Sn��^�C�U����BWn����}k��k5���2��(%@V�{ʇi�_��Z��eV��fy{�=.��tRxp�V`�ꃖ��7Q����".��<��U.��������g(��v�,MQ��}�J��ˢ��i��"⵾�6h~*�Gm�uu.�����Y��ྷ��ݲU�����Yc�쨂�mO;�Yqո����V�m{j�ʭ�<Ճ��7��oqS��k65���L-�u
��Y�Ji�,�I��A�v�$��UaO-�M-�q��{W��\�=��n9�?K)t㡎MÌ݉��_Pm�k�YoGn�6��SM����k�>b�a�����#Aj�x�
 -��9�Ah�|ْU�xr��7-I���������D==�f����c�Vu�ݖ�	��*�WE�ˀ�m.�:)�m���Jj�vB�md�'2���m�yl�U�k�	K�r�q�N��tj@w �z�w.�u3�_T���k��Wj5}I>�Rҿ�jǌ�\ UH��23_,�k6��nˈ8˯�Cs!*���� .v�t�Ҡ�����D����r�
�	ꍘ�t�2�p����S]0��@]�|S�{/�e��t��}PQ@�g;��g8&�C�:4�Kz�1���c9� 7���v��-�'�R��2�iܨ���'�ؤ�W���WnxY\�9��f�*����O��ro�}��ռ�%G��5Iꆳ�;~Z�lň����b0����y�I^1�K��Ғ���Pv��S�㒻(�����J��A��5W�<��S��J����f2�GS{�RTv[��۾��=�HK� Ls\����n�u�����8��>ߊſ.�T_Pg�v��61'���6�ܖ���^�O �+h.:qC邾�i���"�9HF��\�+�󎱽;32�D��-����Sr�k���ym��� t�L�����TFi�]��un�L�1���@Չ���}�G����D�7���˔�c�z{rx���q(�ξ-���~~����#ws�3$�q��g{����>�ծ�~�Ҟ����|�F�϶����~��߇{�O �4�`Nfɝ��A˃9��JڌqΣe�\jn���mo'��.e�	�M��L��y�{<�Vf��g^(�ؿ-����Pߜ.m6C��G�+��.
ޅ�B�s<R(.~+��K��?U�K#e:�e�)�����jS�Vt����Q�D�ߢw�z��M��~[�o�Ω�N��z�E,�/V�G�6�J�\���we[BC����ٟ[j��*���-8Q�]:�ݮۥS��y�ojzN���FM:F�eP��%1�0~�wU�CA�;��$GPq*���ۿ����i��T|����1��Y��ʞ�ِ�Z��E��NweC����m������r�{����u|��34�ڲ��Ɋ_g��4ŭ��l�V��b{���f�9o�z���<c����+Q0$��D�*�z��ʱr���{,$��^��z�!;݀*�3��Xy�!r�2W6��j�T����+1�,�X��}����]|(�
�*p���K8K��)�8Ky��^�Vyؗj[�w�Ǩp��ko�7��!�"�΃�E	�L� !'2���3J�8��9��~/��-�*f����N{��#+Ui������W,���uo�=/�>�n2���)qOq`!7t��a�sX��׹�����&ԕ��kyN�7^�%��Z�zڸ�7F@mλ΁ĩ�3�����[�שF�'|�s@�΄�K�S���v8X�]]d���\�9����R��NTc�u�ՕQw�}���^,#�i���m����ɘ�5�^2�.ri�Q��Ue��v:�{�8#Ş��z�3��:	[=H��D�ϯ�hO*��m��};C��M��8]1�2e�y=j�`��u�=�#���CJ���hu
�^�D9����v�w.�w3�u�(qgw�!6�K}
����m(;'�]}*��[!��SYwއ�&FS��_6��qj�����3-1�U|�)�����������K� }�Z�켿��m��A�"���R�`����b�-޵|3�3x�p�����{�2�����'��Q:m�,,����]��@��y�)�"c}MqU:�Tn�M�,9br�)���s�#U9t܎i�Mu`nI�����gv>�Qdy��uuf���o~K�^�bs�K�k�1�S��;r���ư��Y��;֢Dt��TN�5Ձs��Ի�A�t�����̹�t�b�n��A���G�5�+�S\;~��m
�͙�ھ���N�0s�����7I�޻ru�}�V 4��1�~�%ndF'�c���6�n�b� .�2d�Ɬ��M�!��଎N�![<(�ɞʶ:b�Oy�1Vj�{H��\7⫥�,���������6�P�LvY}��խ�����������X��<��i�x�o�D%N��)>���S�G�<�gosh��p����`gZ��`f�|�/>�yQ�3X�~ަ��>�~O��$k���12o�a����*��x��Eb�^^����ޭ��;�gfv<���e8dIO:��b�9�ݲ�*
����=�){_y��|�	���;�B6�/�L
�ͭ�h$�u�&G�m���Y w������O઻��{wQ�h���� q�x�[�P�ϳ��I왠��F�O�3��+�����FH���҄wf��7(u�L�{%��%*�6�8̷�����:a�����[�/�����
�r��7+�m?D��kM�Mմ�2)f�x��5���.;��mJ�R���`�m(J�f�SÝgV�,�!�G������i�x���	ݔW��,ыZzӝ�������}N�M-_8�����4�_Y{Z�.˘���J+�0���R��¾����Ԟ�i(��n�qM��S�ܱ��/uC�Ip�8��Y�B�W��u�K�����5;�'�j��Ȥ�7������:(G�T��R���1;��ّ��.���F63rF���w+S��G'iݘH��tZ+��vF'�L��&}ʣ������/�a�&�&՛牐��⪜�	`�'H�
� ��-��v��zͦ�G,���G'T���d8r@��8���,bIXVZK�oV�fI��T�R��Ƭ���p����X��t��$$6�(�s���Q���g���7�l�I��6*Wm�u�:�'0Vp�iPri �ؔ�:� m]�[�[�iV�o�`�,m>��q���Wّ��w�"�0�I�v�i�%d�n�lt�o:�Z�8�|��}e�ޔ��|%F���_B6�N6*Lܯ�V�ظe��j�n�I��V����wʜ����g`*�yVl����W�8XW�S3{+��mժ�F��b:��l���sܩ��i�ܪM
�fzӚ��Ml�17u��>�b�Z�ñs�f�Z�7�Y��З��.Qn&V�Ƚ���j;S�����?&6� ����o�49��w�.���;�q�(S�'Yz�{���U�n���Y�J���H�W������9�ۍd�3�{��]�{�\9�;q�w��;qIu?�����y��\�|��j�w��ik�͞��u��y���W��cNS�z��>�4:1����k����i�����ʹ�u�q@��é�=w�7M�QK�BSc�������Wd]�c'�;J���	�&bQ�l�$GR�!�5;�i����"Ѽ]ˤ��Pcxmi��4�&Ħ*���Ǘ�4%�I�\G7�du'�D���)�M:�d�w���2ƙV7�1�L��ɯO9˞՘������W�<F�w{�o)@ q�|0IF��6�h*���on�ᛝ�U��3l�Ǜ��bf�9��*;X�W8mwV<dQ"�]�5������˷&�B���n��v�]��K�%T�S#`�jVB�)��]�(����Fc�v�s�of_#���x7y�&�V�l�N������)n����͢��fJ2�J�ǎU�l�����e>��A�qjU��L3F�������XÅ�΋�:�¹|�n�H���R��]��Q��ٙOk\���":��@�2�C���';,��pE �Ty�n��DM�$a=��.󂙊.����L�^��'�����|��m�z9Nȇ\�G)p�7�Nb��}=�ڝ�I����E�mƓ��Fz����r����|Cc&�o�t���\ٲ��[�1�Q���g�j��otM�m^Lav-@�o�1��Wn�O���qe���R�4J˜��1���[޹�L���Z�V�r>�D�7hj�\0��Ԝ)Ž-
Ǻh*l�o������hL�$=�S9��<df��f�n�k}�
�"֪eL�ٌ�[I�i>�����[�6���dM&�Z�CyE�\%a��*] �u����A�AP!����(�4R�@;b=��I�e�:%ҷ��%��˃�����dvir�1]m���eeL�J����ac��%d[���}h�x�Q���'P��{�&!�[����wY�ܩ`�n	�i�h쒕-�<�<�����"�,rs���KEN�@ҷ��I��4��Z��xb��{��꺵H�9��ݲ^b�b��0,��:�\�hѨ�e��!�$��X�5z��۫T��.��Գ����F�x�JG&ΧG{��@K��>�X��*`pV���A(S��]�2;����=B���Ӗ	|�{�;�g�C{]7K7��N���X��Pmr��f�A�K*�;�0q�!L]��g�F1ˋ�Q����R����a��}:���f �[���i��jc(�#fк뗕|��
�K�6d�=,��P��r̝C��u�p����mB�;W(��]b�b��ݷu�C��A��GY֯���jJ���5Dvem.7Z$�YÚ�l57��k^8�5��&�N][��u�]�q�<9)��KT��������\��pc��$���|,���v�©m��U �b�V:�GOvI��F3x�a�JԒ�c :�>����@�-�sW]��%��r�2@�o�i ��wJ)�	P)d����z�A.��:�}5-�N��3��\���H��@;s)�,��}�X7;J�Q�]�y��㣵)��id�r�4:S��qwA$�p���N�]؛ܮ�kV:���+��P�?Q �����r�s�������;�dss ������˝ۅ���SA��������黴sA.\4nr���s�䋻�7.P҄S\�E��]2�W1�.Q��wq�wr�����k��e�u���4�	$�f Ww2�� �]�9u��ܷ9��젔�w\��nt$\��u�u���+��.�WY�";�f��;Ew\ܻD�ː��b��1��1)wk�w���]۷+�\�]݉38�wrI�Χ.3r��w:��+��0�L�#���q)��B�%;�@�](�PbQ.\��9��i1�@�\�p�u�w\�(�\b4�wa�R�t�7s\B(��1L��w]��F��p]�\�]�+����˻�n�J�$w������iZ��T�}�w�)�E�i�t�%l��Tbm��^5�$��B���ܻ�|^u��+m�-���ǫ^�;�+J�s#e(W��}��sB��LjOE�:U�v�\@��J�u7Gb�ֻ*A�c.�%}��i/U7z:���"3�vVl�N�M9GzI�}�k՘+u�Q���#Vɧ<���f��*���J�]��N�K[�'`�^��-��}f����w�5P�<�;��E�dh{@���'��YJ{�e{�w�͞��Y��4�ͬs]�J��p�י�}�G-(���obP���9���by���Qx�����ĭ�Ü�����\�S\K���M7^�%��`��ԧ�&F��F�{<��7�R��z�b�ަ��\3�l�k�N���p7+ffP�;z�n���*�y�K����=�(���J*;S��}�5�V �$��
��;�WP�o\LR�꬐��s2���b�^t��k�[Mw^��s�oS^�YJ���Ϟ���i���$(�3�����6=ģDi�g=�G�R��SƢ���8����s�W� �#'.�1���Let�z�	:��J�]�fs|a�"	��{jp�8��˲��Y���5*��N�#@�+Vm>�.(m�N~��e�	�M̿m����^N߃�\36&���t��~�%���;��)s��ou���q�}gyÌ�	����D�>}��%��*���iw:x��﫴v:�:��y����ZO|^R���&�͸���KU�ۨ���q��r�{Py8�+>���햟l]�Ҫ�rH��d1٢��]v�zv94���ๆ�%�56 �t���$MGf�GPR��7�jU�#�]��s��(�ᔚ��hV�S���IB|�'��)ڑ��[W�7���+��wpfX��H�1��˚ͤ��8Z�t]S�e���EtG ܖk|���n��u~6������i���%A*k�g9t��a����¯�TV��֣�݌^=4m�.�y��T>X���L�|ڇ�
m�`KLu�>ܖ+�֕ZbU�g����3t�F:"�y��
W���D����e�+�%�首���pn:;�+Y��@R�t��ĪR�n�ؠ
l����n5�Q�w�F�)M�ȍ�)���r9�bR��Y�WB����F㈽�W���s�:�*oT��M@چ��/&�5j�d¬��e�W%����qZ��Y��[��Xʭ]YNo�~�g;-�
��I�ėov*/p�Y��l�~�h;G�iX��yx���e"ڳ�Zd2�ħ��m��d���>�rz�]�SS}og~Όub�qU� N�M��� 䟯~>1�]�7��7�[چ�g��K|�����n= kz�wN�м��׹�l��n~��̈��P[Ÿ�z�5&��Z[��_��gJ�+�%{��ʋ-UΪ�����6ިt���vS�e�./���l�ĸY�X=BI�c��VV��?{���{�5>��|,Ij�TV�-Oq3���v�GL�25TK��d_5���)=��ҹ��k�u��'|�&���p�N���a��#���s���;���fOpU��q`U�	v����iw�R�֛|��{�j�m`u������|p"��iH�K*��̏��=&����,+�]��궧lE��9Q,t%�!X��w�u��E����T��g;�dV#�fM���EP[`-Wf�Ԇ�r1��I�)�/l`f���\��͟��5�r�}ן���s�u[�8ؖ�$M_S�ޔ��|V�p��O�8�T�}�j7Uц�=F^�Ui�+�r5]�qyQ��'���G<�Ί�s��n�=�ܮ��-��r��Y����n�{���Q	̦���{!U������Ѯ�#@{z]@}�i�E�uE�3l����MIN6 ��sx�j����%�9�c�*Sg�p:�
ܨ<��}x��V�9n�IR���N�Q۝����Go�*+/����b<�Q�o��{��)���m������\�o�в^rz�dCCg��e}ї0V�8�h�t��٢ȃӁ��ͱ:�ć���I��Y�o������ۘ����˩K����$�Ԉ5�龘�Ψ��-�N�Sa[ow"�mD{�a{7�C��;�Y�q9��F���N�h� �4U�W	���"�����|`�@]��V q��39��uj�<�e<O]�ץ��ǐ�%Y�M1G�O{h��>�՜k��tsrj�P�ay�o��EJN��j��PP ���(vj$��86���,���\s�bۓ�8�������:S���'ɮ(�k�f�V�ת�Ӌ��q/9��냳�5���Ug���Rw�K�3:����8�Ʀ�Gb���r�OS}�z�T)�V:��PzNƺ�T���不�2gꭕqqˣ\\З}ܧ�I�m��m������r���R�pOK���k�5��y�����G��oF6�y+|;U�ѓN��NWDKh:nڸ�Օ�m5%rh�uΘ��a󻅭W��4_rP�N��ι:����x���]��S\�yqve������[�^nՂ:ź��7T��c�[j��.˞nw�����[�x��@W0�-�L��KA���{��$����붽,~8u�/����������K�[�tԿ���Trb�P��ˤ����ãѽ6�]\�Y�i�Vx�]��sz0�Dz��渜\�䬬�H!�|w�Y�0(�Բ�,V�u����wV����f�͙:��������+xu�QػV6��}��G|�]�mB�)s)���{�u���G���:e�\.�B|�c��S	\srө*5q��,8R���j���s�\�����<�������_5%W������{��K.X�CN��]������m¼ښV%=a����m��Gs����ov��e[���I��+���R��ࢵۼ�H2�R��5Ցݸ�Ϟ���Ӆ�<��cl�I�A�O �*�G<t��k�Mw^�G}��a����-g�9�����]���i�[)}g��Dֳ�����G����{q���Ϟl�4�����=0W�PkZf\�t�t7�\�"� �;O%�.V���],jk��v��ƹ�(P�츗�~�]�M�;7���_E�;R��>_|�v��ۍRގҵ6�U^�v��M`o�X��Q$��.j�h����m%�ѻ��ј��Swz��q�-V�'n��]���.�5?��zc�V����]�'�>����K�:ža�T�j����&��A���K�tc&���TӒ^-s��m��CtsKں�2qA�\r�`V��ާ���q��������=Q������w�Z�ӱ���\l�#�l֞[0:ڷyT�Ō�{DE�o-47`����\rBf_�1�\��8��V���[��)��ʸ�ф��d-wqv]oz)��]�:ݝ/{��9�%��v���*��eO��h�s�p��i�fM��LY̷��t����l���U���9T���>���h�}�5��S>^�NK�nwU�}���3Pr��C==	���'0-0�{i� L�paWc���A]������a�k����N[njO�Dy�w���^ڱ��99���� u�
�{h��H#ݰ'�n$���N�'��a�O����4��c���2!�w^Rg���3�o�2of�\�E�c��]�(g��N%#���B�x��_ٵZo�,mE� >��=�}��\�x�d������x�T=�:�\7��\/mOϦ|3M�챗[p��+�9n��ޡ3���É� �}���9�W�xq����<�K�q���k$��q�=_U!�vQ���8G�c;:�x�E9Pkۧ4���H^���U����.3����x���7���(�R>�,"�w�a��5�k=m֮��l��3�hl��U�r�!s�f��r�+^�XPR}��Z(��%g�[x���%)�)���Zā7��á��<�	�Mv�=]�۸SŋlG��J��)�z&t[c�4z�=v�yU�ʔ�֗��x��kX��L�,4��BIt�9�T���ŋɝ��6�q����������=�>���C�p�P�+y��p�Z���%|�Y��>5%2��D�ȫ��'���>�O���p�ǽ�si����w��1Ȼ�c��w��>��;K�PO޿������W��Q��[�\x�ag��¸6c-og�X�>�>�x%��C���^VT�� ��<su�P[��}��������zK�ӎ��^���`�zCYq+֑~%e����Q�w _��^�� ٹ�è�T2��#���g�s�f����ȉr���b��[�7Ģ��T��mNK�E�IS�N�}f��r�cв�I�;����qcn!?[>�R�Ldzr��O�@]��\LN��.+��\}��$/��Q�}��x���B�MVѸ�s�ݐ1���:2��o�����&-W���CN�M��yԶ���dP��H�h���>���
��WI�/O��j�87F|7!A��O&��y�;Wv�3��x�1u�r�xd9�DR�IG	c�`ͅ�y�P�6�ǃ�ez�곲a;\%�_G�����fQ��;��������f��.�an$�T����0�̚�&�oVq\�bn��_*đ�~�$��q���&���������5���(�-�ʱ��5L�chYd��h��w�r�C��*Yij7��էy;<9��᜻w}]@~��ٻ���wL��L3�򻇁h��J9q,-7;,e�z�:Qf�B�ϼ�Ac9��t"��Ҋ>x�B�>ΟKm�y�γĨ�9<j7���e:��N��J��6�|.�꯷dy�%{��G�X�9�3ң�Xp���N#��;��b��Ʈx�-�,G�X�w��Qa�>�N�~Ȫc+&��_�3�7��x�t:�׼H����{m֎}�3�=���g���b����*x��=ćd瑱��+�.2gY�c�F�+1��=<���]8|�{ר��m������^��8o�Τ�T��t������S-k�����sΌ�im�g���K�9;K�����_�Uj���w��*�3�w��&���X*��>���q���M�6�}�*�8G����Ig��ҽW��Ȃ�����= r���r '�]d[�~�,�茞�rQ
��BT7���gNu�;#׭�<��t|&��,�V�>�켉��D�� Fo��Q̫:\�����Θ���x?��\�{��q<m��N��(Y�^~��b�Y���t�cl�S2���!u�W���n��Wv5[�GWqIh�D�̨�t���O�䘾{PL#�/Is�����ߋ��qMoY4��P�0(����z�=w������I���E՚(v�Wt�P씓IK+8��V�a�z�,�wq+�0=��;R;q10�WH�����9�-�,y?RG�>�y�Ir��G�@�]���J��=���yT����"e�����E�LM9�A��~.^c=t����W��`l�����'�=�j�G#��v}ր��,����D�L�-�6��!U��O�.��Gc���q^�j����y��/Vٿy��(�UQ��'>gĬ�,r77,%}~��ʲ�tI�H���\&����3_.�_��d{#Ϊ\��Q�~��Ǳ������>�E���]IFdd{�t���7�Wq��}y:+M����0:��#���|�N�O���XX�Ӯ���c�j��<cˠK�Cg6v���{��p�k�7����[X�${�/�C�Q�ldz���>��5�~Om����Z1���ٕ�׵�K��S�]��ny/P�]ϥv?��\�q>��]��h��!��}��e��o�,a鐇��Wp�&w���P�ޙ>ڌ�k��@�>�Wq����w�����\o^�|+<�#ұ �R�UP�QW��0$��W2�]r�K�JSIG�NN�;�X�U�Gol��
M�
R:D�Ԡ0ݎ0<��/��Ѡ~�X��u���&��̙���G����\���[Y,��bOY"[�Ȱqv�T	�2u����;�k}.,4�tTnjYZzX�O�7n
}Geo'��w*��hȐ�� �&U��WZA|��Ƒ�5�0�ȧ=�@��ypXI[����gmK����:�J�qX����0�kP�[ے�<�2�.��;��]D�\�S��o�t��3���xk<����ݑL���,�c�)vg��q�+�y�KZ�u]��
Z_uĵ����Zd8cw�p�W[��	{
$�W�dh��|.��}MnY�8y���[m�Oq�`q���K��`3�T؃gّ���P�te5`+9t���x�i�X�X��+�j�7�N�E-��+�xi2��:���x�*|N�W�LrOM-��ur�i�ۏ��� 1Y�^Sj�i���X�ެ�R	s��VD'�&�vֻ��&>��z�r4�k�ӫ[���Ș�ʞ����_��9|�<���'1m��N�E��v�ƃ\�s�w�����Eu��N[y�L�r��|o�
ث8�[�*�$��;!���B�fK9�&V�9s���e�Ed��i��m��,er n�I�ke�c�@��u�pd�.����aV7�si������\X�i��M	��D6ջ����)c[�H+kV�m��ۗOӨ9q';���ڮ)���!�m�ڥ�P�*�M��=�m�Z}69x�3��1N�u�2���.�DWw�S�D#�����OvJ[���"%�w��尤�̦H��@_�s���sJ�Mk��٭t\�l�v)rh����У��Y�3�gW^m	HSugx]����5����E����rQ�pI@�]9A�{��W��A��@�)��(���q�}�Hr�U�}ہi�*�n�z����}K1筼Nb3'�8����<
ö�m�1��{U�붸!���&��*�W[ 9��,�yŋe=�@��o���PǆՂ2�v�\�7Z�$���~]��ޱnޛ{E^��z!��nI�����wΜ�E�N�j�6/�.�=�gks�{;�<��lܧ��#%n"��*�*왳7�Q�yXx���Ѽp2�X]�x�z��t�o���ͱ��ұ�E-U�F�qꊅ�����}s")hk�&�Te�=�P��n�b
�_T$�F[�����hV���$�s�]�$b�.��QC��{�fJ)|�i-�goP�:����^:�A2J�<:>�gma�\����y��iZ��nsD�#%j��줍��Xޭ���,��]��m N�.V:�f�OWD��0Y��ݪ�jo�i^K-�.#A1�P�[��Z�%i<��v�������{��P�a���wC��\)c�ċķ��ohcᗠ��Z[YZذ��wtXk%]����1^��HHLR�d�R�,]����1��]eк���9��s�d��܊r�sDw�F0�����wS�\��6��	��\�n�9s���4c�!(�wn"N�]ۀ�u�mɉw\�B$"0��ݓJ�ݎu�C�����2��.;�F3�]�M�H%Fӝ��9�wF�wnfA8\9�4�vTJ"�����Q�̌�`��h�"��
wsH�&s]���J@�����I����bbL19w8s���wtJ\���ݔ	���s�βE�W"%9���w	$�D7u�\�"\��;����I2�滺7tr��˧n��̹��q)�;���"��R&sus;�ݻ��t2�qG9ݺS�뻴+��ͮg:��뻸��7�1n�9�w]4n뻣��n�Mp��������"���5ҝ���nа���w��9uN;���39�9pv#������<�&Q��=�3h���S�{��9͒�sm��U�3�(d.��o��w]{NG�/�#��//�5�TYW Od>��+'��3<�@�~��~��)7(y��wDz��h{�3�"=�Wq����u~���d���L�yB�B��`Z��a����+���)&�W���BV߱
���	�x�h�� ��ܕK#uW\!��sp�Al�=��Tb��,9�}��낭�FB��9'�B67WNyQ�n�����u���N�k�zn<�����A}^�G3��"�����-��Q�:>ƕĖտ'�W�[ ;�����r���ñ�TZ�1�}Y�+s1�NC��5�zzӘ}���6��F������3�9����e�P�}*I0��oO�{����ڼ��5A�p��!�.^�����e�n�F'>��q���$Tp}D���]Xo�8T��w�`tM"Fi�D�BY���d�t���\�u1�n�O���\_�΁���}M��/���c�k"l^��� �^�+�|v�v�z�+tøͯq���3W����~�.��EH`j&��� ���2�����	��v�PY��3�WE޾�'���e�uvMu�\gY>�Ij��K{iV��yu��ki�5+ij� (f�����З�1����9U��ss0[R���v�mm_n��J��J���)sb+3��p�FTxg�Q�_a�����^��;G�ݬg~˰���x&��tܪI���纡�f�i�/ǧ�O��d���̽�QRe: {+��Q��M|����+�o�=�"��֘5�=h�f�qJ���c�=���n|�F��>���/���	{���~|kS��@k��:6r����T
P��gN��ɝ�Ʋ�^������{�qس��{خw���J�V?"��=��k�zpL�y,�~���{�݇��}�>��^G��^�\R��{,T��o��b��Ny��a\lL�_I�3,	<����+#j�;�׸�dt��h�ní���a�U���NZ=��W�\�C����!��<z����ax�z�5�V�^uR��;��.�z3�z���7W���O���&Yj�A<s>20�H�ΰ6i����D�@��q�D��!1��I/�x�;�	�Q�^��̹>���L�;.,��v;ަ�Lɿ`���9����B���y��>�^>>��Qϟ��w�ˑP�� mqy��~�cc/o2�ҳ�ћ�c�KF�<l�:�-�]uJ�1}�=��f�����F*8즥7v�܀m��~��|�wL��깔R6#Z�i�"��:JW�Ӏ�D��h��,eee�j:u�(�QL�e�g%&�lt2�t8��bQ��!�ͦ��oe׎��+)���o���Ҵ�#/M�o�����;���t�L�zp��ز�e��csM]�o�Ǿ�%�G#�7P�'�ĵ9EF����
�ۆ����W����)ړ5�+��<$d�j�D��=p=vA��H��#�7P�'p���WI�/O�ڿhA��E_ e�zTs�B��{]�/ސ�R<�4B�xߦX��^7���3k�AЭ?&��o�O�5F����Ϣ��F��r�<�e���T5�w�8o�IG.&XZnvXɤ���d=�=1�_���<�v��P{3�����_�=��w�'iO���+�����^�N�z6�y�j�}�H�Pҧ�#&���X�7�F�n#�X.y�sӈ�<�[�㽪�kۺh�w�4��b{�f=��/M�V�*�3�cc&w��� k��^��}�EE����[���2F��rV_ye��}�F/0JF�O�����~8�X�ɝg	�]��+1�'t�{3�v�/o��_����y�O�'Yhh~�(r�dJ��K	M�5	��ø�)������6w�ՙ[�57r�Py>R-�ޭ�[k6�c��KZR��+]H<�.�t�!Y�^���E��vQM/)m
�����is��Y�z��5��@��*ԫ@�)j��]h�o*&�A�{�A����bt����C�R�/��<���]�{M���g�\����	�]0ǝZ�+"Uy�
�:zd0.�Oo��]]��l�D���w���U����q�G����Ig��F�_�_�� ��e� 6eU�[3���{�$$�	�ڑ⧑7>gq��ھ����*�}{M_��=}�Tb��;G������px��k�j�a+�aȍ�K�x�7~V��D��=�\�3��O=w~�V�٫��fD���Jn| �z�&&���>�i�Z��E�?JGE��ʉ��4�/�qv��G\m_�Ͼ�����{؀�y%`~��N������~
��c9Z_�wxF�q���G`�J�K�Z�gй
B�}5�~�P� �~�d<��'R�;'�AᲪ��]:��s��o���+�O����q�/��vj6��͛���s�UQ�r�������܉�*�u�y��g �d�������2u���^�&�Ko�2<������u���=�3�8S����So�jW'��o�'�S:v|}�Z=y:+M���^���~���:��z'�#:��Gb�XJ�`e��x��;X���.�γ�h0����<����$+�]X�3�ԗe� u�Κ9`Ӿ�P(y^R���W�|^�:�9=� �l,ޫ�u��t���ܸ�l�f���A:#���hQ�&��/�Lox��i��V`�{]C��8v�93���^~�FC{�y5��jv���{��5�����.���"��y�Y73�}�i�8/����Lu�*CA���v~�����>[��5k���~�Eƹ]x�`����Ֆ�����A'�#�����zu���
��m�2���(��L�����UP�w��ĺ����p��g�:}�*��z�7���To�?�����Lz9IG�2@��2���H�>��h�y�����{�6�e�|3jW�K������ޟx�w�>��Fl5�,�]'��-�l�����;�X�ǀ�>�T���W1S�ɿ�Pl�c�#���Ŀ�W���Ea_{�^F������\a��`�a�Y��gT텾��F�i��q.��-�*�OĤx���D>��W	�T��W������a�g��eӁc���I�;�<Vzn�:{�R�W�a�Z>̇�w�x&X�0{ate^�w�c�⇦��D�V�v��/=@1/ٞ�Y���<������Т����?;�P�F��.51_v��h��#Y�Tr7��MϺ׎ep+ެ 5�ˑO*�)9+ôϕ����]?H�P�(Mh��n��~s+j_�]ڞs��#��G�����*������Ӭ��Ɩ�D�ϟ�鋒�k2^�]A��kJ|����Ks;��;KC�6b��v���wv'g'v�<�+՟jԶfn9�5]���:j�#�7���������y���)��{�~W~9�g�v'�@;�:a��J0�:jud(�yT����DǢ�����q�D++L��N��#/Ktf3S�M�_��yND:������r�Ϧz��6 �(ӳQR5�}���IG{麏+��/�I�s��|�q�c�'¾����GU ������Ϲ�����E������;P�y[��׸��={l �t�p����5�ޱ��h�ѽU+����~˱"���5����e����CÞ醣6�J��xcf�k��c.��#�=Ξ�G;@
���`�:_Tz5�\�oEh����3�nvX�
*n4�#����������Efˣ�>}7�}��^��6��C��#p���o}�<nI������!����������}U�Td֕q�;鋍r���X����6��>=Ō���w1[�M�ks���Qp�Q���%#�s���.{ŋɝ~���_u;��x����;���C�N�d��4�@��}��q��m�0�퉔jO�SU0&���%=�ۨO=5�|6&�*�W-?5P�B�Y���]��D���5m�U^�O\�����:j���\������x9hx5�T_c�|4=`b�X+�C\�а�A0�wk��9���ػJv��zT=�tݒ� vf	�� �b��m��§WR��
��h�6GS����,>o�93^>R�uI����;��Xp�b���;!�u5�뚇b��M�^/\^�_c�݋�J}}�C��+�,�7������D�wg���^���/"U\ ܁�7*�4xe��K���ۦu3��t��낍E��&���/ģ���	�W�w"����^|��k��P��K=KdZ�Dc�g�U
�;<�`>Nb�~7�{���~�x�%��N�{r�^��l���݋�vJ�}K�DG3�11�j�Ȋs�:3��Zw!cn���}J�1����1=/�G��t�O�h�����F.����k�Q$4w�&�\ex��j����;�Kkw�t����ʊ��U/�zV���=Bvo�P�� �^��ϐg�;^���+����ǘ��N���3�2;�.��� �@.�}��x_�U,߼�&n�x3�HK�%%�̓6���C��&��@����5{v��h���&oj�D'�~ӻ��Σx�B���\.������N\����2j��b�%3�C�ݜ�v�t/�zX��d?Ms(��q��g\M��gJ���r��:���,~{=����%x�[+�L�ySLT��z�be�o����G�#gtkD�n�d�&!φJ��Mӏ{G
p�ة��Y�]�	XfW��u�c�`����VS9�vY���+H8��G(h�Fvk��)
Y������'Z�<��l,����W;�p=)�ן7d��؋���0�aYӸ,�?�����>*���|��<�~R�#�ry�n#'@�����z!G���?*w;!mɝGv����k\k��`���V�Y5��'|{\����������^R�����J�^_�����9����yHn�*x��=�}%��0�mT��gY�ɘ��闏+������ȑ�f;4�->�/W�������]��{��"zk�,575	��é�$2�7�.�����d^�7�U	�|���������g���.!ի`+�gy���<zz�q�RB�o<2̉��zTg�D� �nm�9��|����~Uk�ٸ��O�G{��7�^\�/dl�������dI�$xG�\��뮅KD�Kgs��B����'�l�G�U��H؈u/�3�G׻�ˍˋ�����pz��,�B~0a*�����O3bʞf��a��tK�G���ӑ7�R�==���g=�O���G{ m�`�r�B�>(���t����� 4s: *c����:ώ`��N��QC�E�O:�r� V{��?m�Hו�DL�x��1>x�7)��O֣��w�^��7Z��ǈ�P����&6�U��vV��<U|)��:��3�L�&q1�JY]CtУf�.%�Pf�I�*�`]YݸTz���K�.G�5�f�I`p'I�.��R�A� �m�8���}K�?
���s\e� 7��@
��EC�T�o���q���.��j=�I����nS�7&��,��>��]J_��f�?Y�{΀�9����T�_/O��O��ɛ|vo!�����XM�ͭy;�5��fj>]/��o2�ާUNc��q�;��{��l{&�cщ8����~��N}'�:vݓ�}q����F����+��#��u���:��j�z'��j�"�#�Օbn=�.#�{MĖ��N�<��qc4�d������:��khM���B��
�Β=���NR����R+�h֋�{Mw�>ë*���ه���2��}�v�z1Шa��=�Ԉ�Y�d�b�g�[�
��m��H_ْQۙcM�Cʕ��''\���G���g�=�_��/�y���?_����~+�"�q�J�;����Vl�)l���&��{�1�z*�o��>jW�Jubq:��}���"=��7�W���@9�L<��8W`���,�C�'ƾ��9�W���^�q��gI��Zϑ�0�U~�� ��<�/����d��]f����V�wW���;�~�ϙ��\i߸���cT�wo��.��k[�[Sv:A��|��6�_�gl98�%�����1��9�7j"C���bI������.UK_ٝJn�R�R�ӌ�9ŋi�J��d�rj7�:��'�uR���ٹ�1H��_������q.��9\UH�%#��x�9��B_n?b7��
��*򍵛��b*��\�;��~�c>=�n=������J�Q^�� ����>�E�/\麊^������#�J�$r=���Y*=��~�js� 6j-M�/9lT���j۬��3k٥��w}a��?%q%�~����/�l �ʈ�uN����X|V.��[]�cO�<�!ў�������;x�*^��f1���}��}$����	ߺ\��0�'�4�}��4}c���7\;��땦EDk����X���������~�t�,|��?x��>����~��+	�G���I|U��CW��]����j5΃5��75'���nl?i�뤼��w�ٲϗ��{!��Tw�J�C�;P�y[��׸�zx��qwO۝��#РH�}����UO�N}ӡTB~��#	�_w�N���[;s��{��@7�b�Y��VGy�+�Ύ�����۰-9�x�5pt뾩��Sǲ&|3L��v���*�;~�*e飙���k�=i�<O�{L�;�ں��2ѣ�K|�ڋ�>�����1Z��k��s0vr�&�Э:U��
hh�T�gVC+ڻi�/z��/g���i6���諹Xg;
�AVWU�j:�7�����%���:RX�;�,���$�$�}�M�qdn�P��ek��]n���Gq�U�<�9�C�*!g�^�<�F�T���Q2��[V�m�.hրN�7��s�;Z���)9}�C����k쇔����T�]%p�^��{w���7!U����#��w��C�Q�6l����\�S2������RLq\�I�\��D��*�bxe��F�#HԷ���,��8i_���fx,Z
�aV��J���@y���(X���ת�Vu�MX�Ι�{����խp���i�ҤvJWM�3!uӀ��������.ߛV\�W���B)θZz��]����<�t�#������&�3�<o0t�e�)H����r��f�.u�X������r��U���V�(�sQ��L�8��V�h�rjTu�/����]t��EbH�&9��T;F>�e>SN��7&�\>�(����#[\i)�<=�K�$��d~_%ٓk]�c6�uL��j�.L��w	�#/��`�g,*�1V\�/��ֻ|��d72����][G0�K�o�n��7�+�(ĺє�f5���[��C����Р�a�G^9Ce>i+�U�v}n<��0y������mi��L�b�[��r�)�-���Y=��{2�om��Lǩ��NV�Uz�8d���>��J��UٍQK��75҉���ԎǪ�'���ӷT��\h���.y��1�t�<9��R�BS(j��Y[�Dk�;���-�՝��i�:��w}{���$�F���Ӭ˽I�^�D�#��1$�PU:��zU���3C��C�9p�	}j�Q+�^�$@1u�5�@_K��6R�Jl��G`��e�ܑ{���v���r���Bn��ȳ+X�i.]���p��T�^��L���o�\���R�ܫVt}��!|�ŗmLn�g}����Z�j\�T�R��J���m3{X�D�����M.7WC,b�s�fL���z�8�O �6E%�c3�2��q3���S�v\�v��<,V�B���j�H{���p����p��q�'�{]�\�F�U��)�T�6�L�R:<�;}ݙ����}�+1�]�����m��՝A���[ݮ��+&�XX��f��CG�b���֎+�
���
�(���m�
dݡW�z��e�L�/jEpl�´�u���X��(���j�1��%���d�ߴ����Y�\:s�*d�nֱA�/��|L�.Z����x�c�YC,���rW����B��d6�t�+գ �BGE�~=�b!�]��tY��u��ԑ'3�������LH3���vpܒ.�� ��!�r��$b���Dc��4H� I�B�]�E3W;���2]��79q(.�!����&N�Ą��`J	%���D�	EJn��v�)��H���H�F�p�L�`h���+�u���E殆���9��&�ؐ�N��i��X ���H�
s�&�;I�I&D;�22�9t�L���.�Y�#��7&)	���E�\1���L��]��L$7v�Y��!�����E�%4Iu�b�LD���A�Hw!�Fwn��Ń��� ��J7:(n]� #:�I�Ewc��Ό2bWN�0R��w2��l�r�lh@�C+�#��a���t�q�uȂB�ݙ��#�����??��<��}+��%t�\u��0�'S�Ex��sh�Y�M�6�7��f�緩��ywr�]����dE�Ql�Ɩ.��H_�nOT?�-\����s�F�_���^�e/z�Q���}�<N�q�eDö���򬙌������S
�&��	�LtF�	��z�ns����{Ǹ��7��z�dd��9���U6`��?B��8JD��=�L=���οJ�s���>��o�Cn���y)<���4��]�g�T|c�"g�D�2�e��T� U�E-���m�$Xp�O9tz����f�U�h=�}�W��ή�`+.�{�!��<z�j
nQ.Z[�t{"^��@��}:m�z�3W��8�M��	aw����^�<VԲ� ���7&*��B��켙�~�Q�Q<M�zuh7<��}pQ����ܿZE��u��:*�n�?L����3�OI9Xf�{`k` �O�`��"��TAr����]/��y����X�v	�%�~������ڊ�U�{Ez��)��h��10�r�ȧ=� �V�ϑ�6�?['ϧ�E��yNz���{c5�뫛�޾������dM<��ND��\�C���1?SU�o\�wB�1��;��Ksg��%D���U{n�]_�EXJ�!HS��jy��^�[���O��g	t��6k�W�]q��ऄ�^M�U1�II�F$֮P�E"֪B����Fg_��;j@��ԃ�x�#>���j�T�|�ǖ8ܖn�ɬbIVh�\�RR�A�&���[(K��n8w��_f���9������v<P�Y/x��g����>���L+��t�Wp�]k�[P�����4?Q�������@yd9˱��#W�J9s,v��f��y1��G\{��h�#��~�]Ǉ���ˏx���_��̲o����̇�'p�8���J�E��d^��[��X}��έ���ٸ��ʗ�z��D��H�[���>���Ӿ��Z�G3�Д�^��(i��ɭ*�|+Mƹ��\.y�o=Z����W�A�����K�}�U�ﲧ�r�;��>YLeFMib�&w��\����,t�ن��}҇
���s�}|H�w:�=F��{/���m�1q�%#q%�=uP�k�WLa:�ب��RY�>���G$-�ףk�=v#u����W���x+u���ϟ����*jK�桁q��9��s�O�f��%�'�F���M4}�uT?������N��W��=���.%*𲲥��b���&k.j/ܑ� VL�Ժ�7��w��m?+�!�l���Y�9�|�?����gW��Ƿ��iˮI1�ҸZ�(���S';�_*�x76����u��j���#ڋ�����B�M��#��ǟ:����W��O��b��W�8���+e�_l�s�i�͈
4m��},�BsqeM/�l�3�f����	��TrS}}�TR���w���9_��e�w%�3�ڹ�9Z���=Z��c(��`׶纼�j����>�[��|:T���h��$�I�%x�8\�}>��	�c}p3��c^����<3rYs��H�ۙ)�9�X �z�&�"�O��@h�lO{�672ES�|��C�>b�%hp�O�\�q@�x� �˂�;�̶v�@pi�yG;߭r�-�<�^�a=L��Vf/eq|{�<j=������s�K�=�ր��,���D�L�-εVD݉;>����:;0�r�CC�z5Q��['G���}	K�pݚ��潓�#�� Q�s1��.I�]vws�]Ɍ������g�Ѽ}7>
�ͭþ3�,i���Ǜ���G�T����<fk��#���=�ҋ�;4-�o�G*p��#���>gNχ���>���Zn6]~�i�<�����u"���j�_��`2���?eX��u1_w�N鸉-��ڇ�>���6kN�zԕZ��6m��['���^Vw����h��z��?3ז��+u]���,�|�ݯ ��z���+��Z~Bҫ�ꢫ����ܻ�X��m']@t!%��gr>�M+��7X�!��ͤ�/]���P��t��Ff
v�.�uo]�㼢��ovї��Y:���TT�FW��R^N�4�t�����2�i^ɼ���JGu�W����@�ޚ���V�]�7|�>{�p�gR�%��0���N��<=W["�No��Z4O�/}�w�泥�&o��w�G?_���_���Fi��w�<��+)���s����"�V�v���H���:83�d_+���>
6�x�����<��w��+�G�}��pٖ����{��R���*�Ϭ���Q؉��U0&*yzM�J��tG�{և��g���zk<1i��,�Yx(���7�x�>�U���T���]��+���x���^/q���o'p�ƣ/*����w75S�$z3y߆{��EoOi����VznD������R��^���oFH%˜�]�o��r}�q{��Q~����)�m ^D{���wB���7sĀپ�'��y�e��]�XӖ}�ws�=�o��MϺ׎A�W�{��f�h��N�����܋,�u�R�������_Q���Ӑ�S�׌�/��^7��������GbN9��l��-5�1;�=��|l�.;st�\g��_\�25���FX���q�Ϧ�M?TZ+6����=S�-�u�b�h��ܕ8U)A���QA�K(���#���'7��nF���G\�!͔]�Iu�u�vj�W!e��[�����d���m3�9"7P�<�U�3�+c)�s���h����yF�'t1���`E� �/��;�
�ѝ��.����"�C��բ��>�ˈ�r�sWC���h��9�+IGz&���/�'äֹ�f�[�������ͩQ��	����TU��܍sk�V=�3� ��@���;q;P�y[�l�Ml��.}�P�5�z9Ep3�e������U/���@���������d���,u�<�S�'�ff{z��4�q^��7����q�lK���V�n`������k�SǶ�A�s��>��<��h�>�:2�+n=q-\�`g��9Ϡu�����N#ݰ�q�����-����]�[�VU�z3�G]/�P�d���J��"���d֗d��b�y�.o�46����7��~)S��.3\�m��%�uX䏣�z�gܨ�VQ)���=uL	���b�&u�vJe�]s�W���7��>U\=�x{��u�z�>ҝb�܇�񅑱2�I�*fXy:,�*o3�7=X�/�n�~�k���V��ۏo��gޫ�*�§P��!���w�&��W���n٬�7��j�ӥ�){	д����#V��ϙ�6s�p�ǽ�F����L���qf�F�Ny�3�vE�� �g$qΰ�0� ��׮�جrt����n�|��,��a�qV�r�X�wA`�U>�#��ӱo@ٖ��yi�Z7����5�۹���vF��o[�:6�[
ᶩ>oz����}��s/x����.v��Lؤ��c� Uy�ws��q�d�)M ԰w���>��}��cg`�qg}��{$����R�����оOd�R��&�����a���~7�g�����[����%>��������s�{]���*��Y~]�"��U: \"�뉉�ꈺD�=�cgԸ�/�����Ҙ�ck�y���VL{]m���D�t~wٟQD���S_�^&&���k���u��v6�y߷����Z��c��3�K��������is>Gnn�����a=��+}���ӷ�r�Q;��>���˱����uR���z����[�<7ӽd;%ٖ;DǕ�j�~ץo�o.����{&=�#6����f�.��{��uRȸ�T/�Ub�8yG\�p�b`M����:{�3�i:X�S����ٸ�Ǻf�0�'����o��<N}ސ�dǷ�-�[c}�[^���8}�	�'���c/&��>�u��M��,�\��Ռ=�׼	�?@��,b�䄱��\~|k?���ò^)�/c&��q�;㬁�=^�ڱ+=���:
%S��{+���f$��^��`]�0�V�׷ľc&�s��;���3$=��5���5B�
�S8���NH;�췝���]f.|CG1��c�;Wgh�$7��.O���N�v��[�5(�����됩�}LE�Y��3���9��=�q�:;�t��w�������/	늨~5�خ�����n��{�s�@R
�q������z�nF�[�o�^G��W��u����2�dĆ;����O�o-�y:�j}��}�_��5����^W���zr#�-��=���v��+�Y�Xҫ�X�gOj��X)�s�P	L�+���_bw�����=�ґ�l���JP����:�)^�T�nB�p�OQ���GdW^��D�d��wQ
ڮ�'�lǫzL�y=O����)��>L��:j�n���W�� 6x��ܩ /e+�2W��w�jF��]��H����D�r>r���l�*���Ċ�S��� �z�&���}���S������qӵ�o���Y���?KgB����NRg�|�ndH���	-�^.���EG�'.�WmT�����um��Éx�ji�Dz];p� {�l���d�{����r�h/�<Ew���W�m�j�Mi��Q�J_n�F�s��7�<�:��9���&v(ӿ�[�1k?�q��s�u�ۅC�),�*���5w�ک�sv���l�1S5�v�Q��\P�)8E���̛��q+ᤇ��u��ɧM�C�J�։�fK�ꜜ16R���r��}t��%(��͞�Qܡm:Y�d����anmhw;�5����ǩ�̏cN�1N��>�T[��]�@��Z>�>����*8j?~��Ӓ|���x~ø}ѓ��޹��׶���~�do�����wY��Coѣ���:�C�o��M��gL_z��3�=�"���I�0:~'9�k�hz��*�b�@[��zH�l�M��~��0s���xa#�{�T<#�<�����C��g1�z;���3���F��d��:�{~n�+�=�8d}��H\fIG}���T�/&�=���Q�X��裁V;�w�L���f��wq����;�z}��~��e�c��*=Jۯi��ތ�Q��H\@+�e�_�L	��øɔ��6�x��N�<���}���ם�-������|��[f*l�t�6�n7�啛 J5= w��������A��S�ֽ�Cڼ&�^��T�![�y��h�a�����w�}�����T�!ĺ5�WU"~�R<M�������	������D��!#�	���%q�u���#�r%x�;�܁��Rc>�0(����+�j�M��]�z��+44���N��//2ԗ�kx,�^�l3K������3҇���e\ֶ'��* ��zo�ꓻ&T�u�G1��m�^7�>�}�*�էޣ2��I��O��讂��ĉA.V�$�-�[�̍:�0h2�b)Ѵ6r��H���w�;�1������Vx�H�_�#�d�[�{$p�׫z|j����2-]�ؙ�9�=*;�%P�.7�@Εd.�f>Mz�n}ּp�+�Y���n�_�G����݉-��_B��O�d�"g��è�TDӞӸ��9�zm7�Y�U�q���~��,q��~���n�� �n��{'�Q�0��c�3�C����s�=��pݛ�k�=��G��/~S�iw;0󺇔�7��T��|J��'���7P��n��ä���A��Qo�1���sC��`�}�W'�����dy�;4��ǳ�v�_w�J�rX�م��+t�;�J�5;�����X+֎��g�{~ W+w�uR�Nw���!>��������q/q˿N�}�9�Nk#|��)�D��bu�6�MƗ��y��i�Σ�")�����T��Э﨧��s\����/?,�ӟ�;eҵ��n�v��x�U��1����U�;��o��b%<�ї�}�e��_W�}۷<U�7	�w��CՓZ^���G9q�걹���N3��j���u��"�ѴmPy&֫z�:3����խ�ώH���tIT$mȺ5{��])Ҵ��Aܾ��'�2�12�_=w��ֆ�k*�<��{�N�+�n��WX��n�R�G;nc�yRGzY|��+&�^9ͻ��]/��˩��vv��_��1�~��~U?|�$�]S�x�d����A�:ʘ�5[����h�>B}�^<2=��;����X�7=�񅑱2�D�"���O"��:�,��a�� ώ����7���>>���p�ǳޯsT�Vq������B�򫏥�(q>���6���أ]�F���d{Y�{�nJ���^�4�ԣ����p�=>��'�HaT��]>��_:@�h�낍D[J�n_�#��%g>�	�������3י޵}wR9�\��@��0{j�|��,-8�:_�E�+��mg��ı�$��o�M�~��0�VK>�L~�"c�T�h�z���^��LӞ�ѐ}+N����T��>Q^6Uϼ���'��U�������
߲�i�ר�r"KG�n���W��jv��\�K�c�����[�k�U�y_�gz���5�q�^�=9�<���\?	`�L�su�}�IS��k1/I�J�#��I�Ҵ���ݚ��}� {��r�xd9�D/A(�GԿ��0�"u�R
���:(����=�|3� ��jeF�Z��ZCZ���h�F�,�p'W�q��K*�&>2�{�i��6��ق!Q:�VS�M�B�22kC��& �(
囦$s{�9��wyO�cÂ�\��_T�j�T��Ymdޏ�F��Z�aVJ3.V�6����N*��z�T0mK�.���	uɋ��yV�V�˼�4HK7���2��i�N�`�C��{�^)4lōC�n�2gV-�[ʥ��I��s�T�K�ǯ{��Ǌ�>#:�Y=��|�]��8�K�mm�S/ �޷I{1ԡeϴ������	���!���]H2&mA5��T���ɊH���f|��Vk���g��L>ĩ.}�)�X;�������y����g:r�ξk7����L�܉�G馊�"�Ҭ[����q�JQ��5q=¶��:��H��c�;���Ш2��E��V��}�%���kl�+g}d�}q\�%�o;l�X�ۭ�вs��7W�,�)p��[�J�[�Y�-`�@L�|y1t5R}3_oJ��ri�/\#�v� kX���nDwg�q�;_gKf`���<=�E^`�ң��g<�����
�:�q�wf�Ǯ^�z��|�1��
(����ii\�t��������5�P64u˝�ⷩe�'/�
8�O�F� �W�^��.��dѧ�9��X+�뫾�!(�ºp����Μ(.ѵΙ�Ĉ@���V1���7�r����TutŔ����x:���.!�o�ٸ}��_�T�����Z��D�E�:k�_*lŕ��9�#Ck�nnn-9��ы���\� �\	�Hj���S6U������\��>]WD�n�.d�Y���#�]U2f�Ե=�f�]X�$1B���� O3֚�ެuš��9��b%;(��
m7��8����z�9|]:@K5ܢ��SH��8c�&�a�Xx�m������l)aU���T[W�e�/DzŐ���U�{J�[w��{��G�,���`���N�guI��{\қ����^Ћ��ˎw�<϶��f+�Y��E`޾������Lƺݟ����r%}�3��Q����@.|+U�B��ԏS�3g%n�,��N���D)x�Ww*:�s⨊�;���jEEy�C�g�]#\i�W �6����S�rU���*���"���k�<9��v��ܾUw��6�6�*
��t����rj*�@��.a��hQ�4k��8�5�|��o)+r�=J��qu�T�G�d[=E�o\y�Bi�$l�I`����0�;�g�6���FD���V�W�q�#����@���e�W>��Cʻ��̶W��M孔P݊X���d2�h�n��(_n+�6�Yh���iK=�s}����ݫ.�d���mZی9}�S�5�5U�A�L�]Aw��$ˤ����/L�d[qee6y��l���guЋ�R���u��ڗu�b��Uʊ�ä�vXz�M�ܽ�ǯ8}B�|(`�Я��5�D��$�w]����$L��\�dSHi	 ��&fiݝȋ��PE�X1IP�웻�İ���M�g8ģ�0�M)D�+�����h�$��K�t#CLFe�˄fE;��
���܄�`a�n&4��h��2�Y"��ID�.�Q#0Z�&��HbA����P���0�ɠK�fd���K3(�3��s���Ba��R��C&i#D"�ra�3�B0C!(�4H��v�$1sv&d��J��&��wLb���F(���C0Ü�(�uv̘�$�$�����2`�H��"J2E�)�w���߮�������/���l�ƃ�!}�ʴ䫕j�M���]�P�>���6���<�i��3�� �pxds@���jms����W�͍㛓y/N���ܸ~7	�nx{�3��g�~�ȸ��>��&�omllo(�P���D�p������u��WMƖ=�7�����d?Ms(�{�ǽ�#��^	�d
�G6��[�8}��V	K�����ZxzZ���e���C��oF���w�O�/;�ǽ[��*��׷<b�	�$;>S,Zɭ,_�3�6�#����}x/C�[�� ���X���{ċ����{~�u���7}�<af	H��ߪ����P�
jcS��y8���U��l���3�#iQ������9���#�������a��a���VI���=��-�d�S蚄��q�W��wp�ry\{���^�l���.Z�+��@��`�^���Q(��r���Q��x�L��X(���'�)���o=��-祕��mO���{x�Ǭϋ_f�= r���@2�;,y�U����^?���5~Oɦiֿߜ{K.
��}�=]���n����^��-�����*5�+�aϋ�㗷��Vk��4VW�S�3�|��kq.HjS���uh�W$Y��oX�WCVws8� �|e���`zRW�sS�w"ط6�z�s6���9P!��k+�2��VXX���P�`r����oQ�5��@59X�ݾ��^
��u���.����v��U�uťaB�~b���	���2��e>�Cj=��0)�5
�Z;q10�r���u�7�Y��B�7��>'����xy�[:�U��G�)�=����$l<�M�s閏w���"�{rw�z�f��0�"И���;���ݟ#P�����~U~9��`yo�t �=�,���1���:|sx�B��'�:;l͎y�B��l�ݗ��rz[�0�9�͛����S�A��,;R|�Yk/y�����E��9RO2��2��qr¿�kC͟	�4���c��dz5��f���F�����W�2e~��+D���*���@���^��>gn'k���N�������k���d�3�r3*�ۛ���^�_\1��w�q��U����oz���-��ڇ���,\��w�ښ�f�B�+�ϻ�]��:�?I���+ӣw�\$(צ�/a���}�Wy8���.�g<�=��MH�_FWTz�1WY�@����F�l�d�k�Ev���#�/��4�EWx��r�;��7kT����P��,,UQ�ɝ��@L����~�i�o��+��\o���+��b����)(���A*��ܤ�����Eb[����jƓ�^��+�J��G/��5�수C5�%-*�Ti�Oe�D�:��Q���n.6�6�@>�m�ٕ9q�:d[�7�K��.�sw;v��#�ڻ��&��jV��w}|u�q�7�mO�~�^�edl�*�� ze��޸xJs�g���7��x���`��6��iGY�D�|_JU~[r�͐%���;�T���yzM�J���tG�k"� i�I�ᕔ���6\P>b����tc૸���S��ǳಥ���ĺ5�S$_Ĥx��	�gW�E�}:�� ˝6�K����C>��1zx�q��#j�~�c3Q�Z5��,����^^j��h��a��� &]���W��#"�_�#��m ^}�#E}�t/����8+��u���-"R�1U=�Q��PWS�G2���C���ȟ+ro��{ư �N�
���ͳ��˽��������73�i0�ڢ'�s�v��=
e鸄�j:��]�ϩ/o��H��u.�/88�#|���� w�~��O�I&ߢn������i�Z��;�6����Fr'gw�� ���j�a��J������7���������j�ͽ�|:K�����3|Gtr�=t�y��O���Q��=7�V<�L�6;�%a#�o:��J�����8������>]/�?��w�0y�l
:����B�w#�T7����۫��_[���x[��S�"�؜�6Bu'7�OM��Zю�0w\�l��8Z��+��p��l�W`wjv�Yԝp�9	������帵Q���s��2V���>�a���]����p5m0*�xkUS��p��bC�loz$���y�2/nh�����s*Ͱ${���,8�c�6�N�x��u�-�`[s��Ʈw�#՗�wZ�j���z�T�p��v��ɖ3M���e�V�,>U=���o��u����j�8�����nBf�0�^_b*<�z9�}<�dN}��p�N���z�VMixN�c��W���+鼍�g��d�������'�d�wM#�}�����ܣa�R7��`O�=���L������/{8�轑�a�W�W�+������x{��q�_��6�����2�D�qSqT��1�7R�שnb��`ק�Ҵ���w��#���^��	\{#ޯ�uv�Vq̇2��B��KK�e=i��g�&�@�]H�	���w~�(g���y�K�F~�_���f�Cf)�xtW���g`S�'��M
�� ov�>���9�i\M���r������C���w�{��X,y
�ꐜʢ���}0Xu��|\�ρai���^y������p������r�y�����mN�Åd*���pXC-l�����Gj[�5�����]�Wp��Rk�顤��ɷZ)�k"���ҭ�L'r&����$������l�-7Nf��;\�ÙWui����-u]N�I�q+qT�s�r���v}g<O�|��>ͺ�_CʧD��\LL/U�&��Ҵ��=Wl��d����N�g�ʈWz�1q����O� ���a��IDܖ��M�>���1Y\�Q5�07|�BŒ�N'�u���7W'�~��ȏK�s�z=TA��H��#�b�X��,ݔǴr�Gz;r{;S�}��}W�W�����~�>+�@���]�S���?��ߣ�n�w�twʼ�;����n3v�כ^�|_5�p�m=����E��P��r<�.���'c���'Ia�Ş����^�(��3��N��a�^Uq�,{�o:X�=��0�[�w{W�x�K�%3:Ч�����R�d8g~@��)~\2R��r��ҭ~�����m��G[�>�s��쒜} g�8�X4�k�,/��\����y^6.K��T�W�5������y�kc��e{8���y�C�׼H��[�"��hW�����b��%#q%�<3p+h�3;T{����ځ>�G6�G�&w��&c��ҳ�jv��o�^G����n�`�`|;*u*�k�3W�[x�������7���q��飮�Nv:@r�`����%%k���pd|3ۉ�
�x����L�%o�hk��c萷��5�yҗJY�O��u��ڹD�BD�,��v�/�{t��e�����2Mon�"���ӱ��SW}��A�"�t���&�\<2ֻ�~9�*~y��xW�-������'&z��H�c/o�,��	z�a�=(�;X��)��Ղ��~W�G����#���uX=� �\������7�_��,��A���^�-q�Ǚ��B׃ޟ<�� Z��� �D��ic��N+�w�a�~�d{`\�>`�jJ��J�X{��ӽIt^��wFy�5~TW�J�w�v�����2=�\����q!���/�G{鉅�kn��`:gt
�X����fO���ں�NF̧��<<�~���D�U��н[l��Z�;�%�zm�/d���^�1l�dǮ�{�<�E�1?S��7��=�L<=�~5����W��t�� /`�B�����x�gG��Ω�7�ς�3cï�͢}~��_iz}F�.��C�1���l����������T��	������x�i7��ˉ�9���և�|g�^�%qc�э�b��7�9'�������y�2�J���ߝ�{!����He�ȓ�v�v�?^mh����L]��M�߱��m"�j����Ƀ��=���\F�^P��*�S�>[���Ycp���=h]a��4.�R��Z�G��)�u�D�#m�ޗ�i�W�a,�Lќ^� ��݀�R[姉����[��^�s��]����J��*e^���y;����^W[]]� ���]hX��:�A_Gz�5�ʱ/�S�6;�'�ܖ���w��F�Q�����պk���}�t{��7�]����?I�?u4N/W���hH����k��{#��c7
���X�r�m��ETv�����:�:��9���vɿ���R�u���'hp�|veS������PGP�%'���}G�⪇�3�����	���w����9��x��"u�pٻG�u/*'U�}	G-���ڔVl�*�g��,��\;�&S���^7N�:��h�����*��>�>ޗ��g�q�j�m�r�϶@�jz@�_�L
<�'rPl�p��?wLl�{���fV2/�}l<��z=]�#�z}��z���Qf:�q.��9\UHNU������Ƨ
cL�3������D%o��E�/y��%q�u���~���+=7"�N�޾x��ɜ�:�zG��DU*1E�xp�#���Zvِ�_���P-��WC����Nc3)�Q�d��@#�z���<�E��P_W���̅0�}��M���x�ep*l���O��6���ct��r�X�ꎆZ4y޻솀I�k�'8ns�z��(Wri��Vvd����H���)mو��]�9��y�:=�qhY�s��A@���lN���§s�΁�1�b-y�I��͊fn�q���H��6�>�� 	�!�+��Ԗ��+ͽ]�V[`�]�#�2�I%�Ҧ��DM9�;��ӊe���p��ܪڃex�R�N��8�I�% *~��O��pf��c�3�C��V��wǻ�o���n���U�n��O���3�j�71q�:S�� z��r������w�n����/�׵N:񍫝y��{;%H-���:�g�t7W'��w>����{�V%� ���Hzr�ܒ�+�S���_(�Xdw�7�]�=f��|灚�����~��:�}'#�@u|��bE�碴qF��swK�mȋ�(�X���^�^)�i�~
�}wf����"���<s�; ��y�b���Gv������-y����ָy�G�Z�+��+:���>��.����'޴_^Y�����U��� �m�����m~�t�2-3��O�q��U�����ʧ��'"ة�۹׺�d��� ������9��x�;q�c��Q���R7.p�`e�x�v��5��O�5���R���vN�A���a������^G���{��U��>1�퉔j$�1Oޯa�70i[���k��ZU���v����7�{�x Jc��ނ�r�yk�0����������W�WXv�Z-��� ���"7u��q���Qs=���u0����� ��ů(�Zs�]v���sQZɐwSu�Ƃз���}�lЌ�ܰ��mP�}�z6{���Ӓc��/K�~��SEyO��<��'��
����W��[&g2Ns�X��5
׽H�¼^�k���Ty�JG��,wd{��j�Wu�D)�����٩��B��x��CsPN���W������M��f�*�/ԑ{�F/�W������1�4S>��k�Ƕ�z<O�� �ӛ�,:�T(��9�����~7B�=���T=#=�R��;DP��O�z�8\���8Z��ȧ�N��G�baz�Ց1�9�w�Oq-�핇�5�M_���������ǣ�Խ3������_CɯQD��Z<ja�tƕ 9����~���K�7�&+�v�izw�K7W'��#�+�s�z�� �^�WrP&�5J$�Ƽ1�GL>��[�:�t��>�꿚��vk����ϼ�u��ݏ��
�:m�ݨ��([F�G��$����v�����ڇy��7��3�P�{��/�<ꥑ��W^����=���@�@G��.��3g��X�/��c.=8\�tޗ��n3��1�\;s�={��GT`43o�s��U�V��h�/H�н��Ch�S��:ډַ�Qɧ>ۣj9����WFQ=��n֍��^�<�&�����d�e���.��]4�\�F��X:���Lð�C�l�@ Yu�u�h�)�/��������{8Mj�捷���K�8��bw�yY�k�	�7>�6�i���Я�
��ָ��+y9�Yb�yE���sﴠ9���:�>~������AG��`���~���n�/��W�v�ƴ�PR�ϷNGL�;�{����.�x��=��؋u��'��C�=����`���*	��\Zѥ��}�c�DO۴�j��Y�f?��ʜC��������F���ק�{�Yhh�xO>���
<��Eʂ8:�D��(%7P���\;�(+�1;�㐫���}ONG�[)�0�	�)�毖g8�b�zƏF��}�,�C�%�w�b�i��8S-c����=���Kp�F{����P�fA9�qi�U��s(� �W^���ܖ<Ξ�X�<�ޛ��ӫ�F�b�^"}�lM�~��g�U����:j/��g���,\-�ϕ*5]Yä�z�S�t�X�3�}�T�ݎ�W�hM�Kv�X��}9�:5dz����Nn��q�O�����	�P��n*������8KGw *�P�$tdK�f�su��7����~{�x����km���ڵ���mm�[o�v�խ�mm�[o����m�뵶�m����V���[mZ�����m����V����m�[o��m�[gͭ�kl��V�ߛkmZ��kmZ���ڵ����ڵ����ڵ�����km�mm�km����m��1AY&SY�|'�~�ـ`P��3'� bG;��*ET���D�H�*�D��)
�EE)Q�*R����"��I���� T��*J�UUѪU� )ITD�H
JPTJUB�jRD���"@�"JH*��($�e�R�H-b��))'��T�JU*R�4�T��UJ)DJ���hB$T%D�QH�)T�@��IU���-eD) �z�(U*�I�:�EHx  �W@��XP*�݇h���l�P�kj�
��mT`�Uhm�SPl�PQj����VPж�	JU @Th�/   ��
�����-SPT���B�����WqF�4h
4h��QE`y��
(��Eyn(��� E gf�(��E�H%H�UJ*#�@  ��k�0l4(Ұ�Um��j�ʪ�F Ѥ�&hj��EI@�����C[J(�"T����#� ���h�X-�����@Jj�X(Y+�U*� 4`�̡@��m�����(�Vڳ@�wJ$�]��J�u��QJ#�  f�e*�(L2��֦��`
P���4M�+I�v�@u���4��k`[
�44����X�X��ҵlXUEJML�J"�UG� �*���wHphP
6���k��3 +M6��j(U5����X4�)j��F�b͵4�U3*�
�2�h�D�*����UD�7�  � i6y�wYմ 1�V��jӧp1J(!d[ec2�ڬ�C#������i�C5wnECVZ�E*����RU"�<   î�-���6�T
5�
��� �
�Sځ�jQCMSkaP�U�*�H�6����@m�5@�ҹ�J41	PTT�<   ��� ##h�m�m���(V�#�G1lҀE`]ض�ڢp��6��� e��4Uh� 5m�&�B�R �*EU�T��R*��  6q�6ְ�!UB���kj�-U5H�j��i0��L� h1�a��N��phZ�i�c��(R�)� ����&eRR��@��a%)H  (�2j42 4 �~%J�4 jm4�USj �d I�	�*���4d�HWBȔN.9RRW�2�������0Ex�ܿxm׹��l��7��B����$�	&d! ����IO�H@�~�$�	#		ۏ;����w��83��E�Ym\�Dn��˭�����`�:��s�a�q�m��s�3A�Z�bZp����wZEm��-;{�� ى,Q� ĭٛw��O
��V3F�_ɜg4�8�m���^ɪ����N�W{l�bۥi���CPfc�W���Fu+b�j�Y!���W2�V�ZI	����w�ϣf7u�A�h<$f��q�P�wi�ӰɏrXz0�Q�� �X�Sn��O��T[VڥH٫D}n���ƚ�æ�AUÛr&�"�^��.�hf$�Nd����J]�k20^4�T2�Tۻ$��(�MJ���հ�ʵ{p=��Sl]<s)TIb�2�ʖ��ؖm������TGB�dY��2Ң�]9F�Pۭˍ�#�iO2��$Oo.���I�Yme�̵���Qi'o(^��W���i�QM��o]�JV���)-�ͩ�p�,� x�Q6�8b�X�f��Q�e�:��R
��U�V��n�y�ޝpKB�Q#����6��*�x&$ـ��ʶ�SN}��Yu�̙���wY�/i\`J�[��-<ћ��!c�-�p4^])*���;T���(�Z�-l.��{Xع����x���ۣ����v�]%P�Y%%�S4�wQB`�rMAyF�W�"Ƈ�tӨ�Y��I�;*2�M��V4��\��ҼV�QҴRxfau��t�m��[@ /i�@��T�ݺ�C�m�K�4@�hӊ+cp�tr�F�Rb���[� �1K����<�Cjҳ��[ɲ�bl��lt�^����;r�=�ؤк��
����W��N+m:+/le;�xr]�␕Y���(�`�����~�J��i���W�E�����i����S*e@��N�r+:Q[f�D2�-�*��U�
u�dRse]�+75�5`y1�7��7MjZʐ�m���kUh���9�c�L��V(!
<uz)���S�i��X�(W]�ͅІ�q�o,�zĥoE! j,�7��mk"���G	4H�HrcZ�bS^̽��p)���Xk`�؟;w�ں�P���Ϥ�eX2�|^H4�
ͣ36���-kJej&Z3I�u$\B�r]��T�"�^<%�H�QSTv˙���R"��ӽ��V~f�v�L
�0Z+I9�ɓ�(-�~t��N	�۽�{�-�2^�q�0"�J�0�^�����,�԰2�]��b�,�/r@�(�#{����B+K19f�ڳM��ZY3����u��¨����q�!��A=�"�T�e�v2���E��q�r�ǯfci�J�;�IY�n�V�כ!b6h,��sp�"hW�b����(%N�K���C�͠�W��l*�5kNT�  cVS�(�y{j���[m�їSgyN�[�Q�̖�`�Y���[w2�6��^m#��	�N����fJ�U�$��?*U���U;�re=e�e��t�V)V�k3A�J��TRk�ɺ�j��q�ĲƔ!��U�[X��槆�#Z�B������Ҧ�E©fC�*��N�wp� �hf�f{�+�g\M�dTi1f��t�oteB�+aY�b(1Aj��@�i�A	�O��`Z���B+�ߓ��u+�n���KoC��G%V��Cu������@%�̻�E�V�li��n
��a��2�;U%�ed	�P��)]�j�ݩN-����j����vc�en��LR��
8�AJ�dHX�̴�ִe\�ney	�j�ƣ��j�Ti\��� B�ǄcGj�4R���m���8qBc"��utqT�A�j�d�@f�+i��(Ќ�Y;C!5�2+3od��T����B����W"ʼ9&V�*�x���`��$�*n�f�ћ�ú��Ԏ��;k*=�x]G�XhY�p�k#AXv�I�<�@� ��,�����5�Ưfdc�{�6�&�=��XњZ7𠍔���"�z��x��n-��&�����d��ʀ�J,rI�����&�������ڍ[�0Y幔n�O�(C"����i�z�u0�q��-ͬ�ub�^�`�{Z�]��S��S�e=ou	�Uٙ�T6C[�� ��ۏe��u�e F��5t	Ƴ�=��3�AB:6�F�D�v�ɶ�ӥ���V��L`V����	�����6q��ܦnC�#Ii�$I �ܺ���Gj�yd�OQ��VeʵU�m��"�q��)E�BzՃX��t��H\�05���7rVE���2��.ʱfR,\�[�pRζ�+J��T��J�Q��sSq0Hۏ*��I�-��cN��u��.�@h��i�Y�y�%[Z!U�udPj��U��^e��.�˙���;U�e��*���	nū�)IDE�z�^Z�G���a�)��ځ��"X��[�n����nIZ���<�gUp�-p��PĎ�9Y`'u��2l$9G%c��]f:g]bMnŧ$YLh�W�xŕ�5�-܁�:Rv�mY��E�w��#0n"�i�B�m;OkY��&m$E\��6Q���캺�K�ۻ���>�)���(�"��Tͼ�C>q�573��6r�3���e�Ѡ��fR���ӗu"�JX��O~�V��`�����f�ٓQ��9��c�v��*��,kb�Lڼ!c��n�Xd!��V,ܦ�1@ KZJ���Y�I6&�`��@���E:��yiMQ��n��M�Zu��F��@��Q1JmnS��f��7�3$fV�!!�dT�J�K2-���b�<�:�-������E��ɬ%L�՛Fh��XЎ9a���,�[��u�XՔ-]V��`1�
��4C�I(�`��F���{`0����	J��QqPՅ=�����f^��`zjS�^�t��*ؠ�J�C02����}�bnؖ%E�ɫ	�ۥZ�,0�# W��we���4�I�|*F@�h�d�Ќf�L�Ո#��v՗[sJ��5��;%�Q�l�
���ۛ�9�pe0sD�hfk�P�V-qV^V�^��2��j�nH@R��1A�(S�a��-����6��S�]:������;i�t�G`U���� 1*7�eEI���!�L\7�.P6V��6�T��Lmn_ђA[��NX��T�V��jV��~Ձ�)e����:;%[y&�/i	Sv�uE7jCY@'X0�/��-Z�m]�F���2�0=�͒�ܨ���!�v����]�O7v�#{�b�H�؍7i,W� �V�Ɏ����	�^�XI-;�Y�m]����d`�YrXIe@�;j'/L�7�T4�V�n�Ĵ�T�Eq��m(���(����,�Vn㰶�1���A��S�q�6'�jK�l�Ov�"]�Q0U޴,,�ۺC2�f��åI �F�V[��h�W��g
^�O":�a�-ԢOH�Ս_n՝i�����"l
5+n!��t�L����'KQa�愶`yyd[�!!e�� ��%�4%#�mê�f�v�,af^�#%5oH�ٹY�kI�]]��L{E�Ɂ�gr����2+.e�GU�hnF�����UflVՁJݝ��/6
�$L|Z��.��V 9u���,�8	W.������]q�m���jX@�Bn��#��,٤�����+�{���.`fP�[b'�CoY����iԡX�F��bX�QT��B��-Ce�tp�f�U�襑 �7�H��#,ԍ̒�0�L�+\@��/k$1�6�����Ȩ����9x�A��i�)����W�����Kմ�:h��j�AV��Y�5��{ Z����^hV溒�)z VMhE$�ƭ *�࢒��Y���U�7XE�C{�ޜ�	�PEum�*�Q����vŌuJr�J�OQ��nQ�^�̘�E	tm� P��kO[ulT��B�F'/e�6�B�Z2a�P[����1LF��LdVV�Ŭ3H��2V#�:�ƍ$,���"2���ۺT�������@'yy��̇E��	��Ge�ّ�O@ū[=Z�n��=���Q�F����CjM˧�(G���^��/)#�2�֐�Kt3}Y0-,InU�>]h2ص�1�t�_�*�`q��f�j'	.�y�E"�4��ry|�����[#�#$S���Av.�Kw����WK����Q�,����ѓn'n��;t-͏v:n�ȓ!�L5J�旜��]Y�ؑt@z��٘ޭ3&]2��t-��a�EJ�4R�F�R�������q��4�n���� <�zr�1Y�6��O�zp�W�ڭcZ�KV�54�x`��
sc@�*�0�t���a�X-�pA�f����K-fꃲ���ֆXu��T��-<���"gĖ�"[��F�1�l�f����&�u�t�1#Df�Ӻ���ri�kAYiԺ�C*L��0t�1�"-֧@�u���7g1UX�wHS�#��������!���ª2�LeD�X�Q�*���ˢ�H��x�J:��EM���<�"v�W�×��r�û4/�,���Zɧ�6V�O(��a'��6r`uy+�����x��QeS0�i��s~��1�j�'�&�ʑ�+�EKn�Zi$Λyg$�.���X�6�7X�̱��4�7�AX��mf`��� 7hzD��V�u�eO��F"c#.9��V�|����Pb5Z����ԕ��k`YŎ���-;��;1f|���o�J�eSr��Q+�r��`�Xe�rK�X�#2�q�5i6�{FDh����=�p	-<M���ڷ�{5��K�6 .`��B�T�YtQ�WN�0X�b�[cݫ�SPEeMvL�s.�41�͒�a\?�;O���(��񄖭��B�[6���훐�47�SMF^D��f!�U��d
�C1�n��^����f��O��Za�Ά��B1嫫ׂmm��wwgk����6����ø�FZǊ���*���K���9!b��Z1�MnGkn,��XW�)+lI��a��{
�Ik�-~�/7�M�ŎRf�Z��գ h�P3*�lnn�Kv�&v�[lXZZid)�c:���W��fT%�u�R��ڲ.��T�K�0fn�����Ï%�m�E�w:T����n�Ln�$B�rEOY[�0b����$�����s$Kw]]#*v�V
�=@c��!%C���ȑ̘d�z��Z�a˳yF
��Me'����36	�c96=��͑�te�ؒ�tÉ��`�I�������%�d�Ƭを� ��wf1z\{
�X�Ŷ1����so4`�ͻċ�:��+t��R���$�Kr��p��U�w\X���@h����jm�-L��r�,qYз3vVVQ�ui)0j��o��bAr�Šb�A(��wt��ö^�� ������K1nl���RM��V`d,Ch�tV�Cm Q�6�=T����p�PTr�����h:��^�V� C˵�2Y�/%K�)k�YjZ��Ӵ�GC��k[(Tvo"5�7W�fk��(�F�	j�A
h��k+2,K�0�*�
��Q\mr'gq�tۼ8�	��}"l�����,��DS� �6aC-F����sB��k���i-�����6���e�R�@�P:n�C����w�
9�-c�oK��{�с��qL�m���{�ڹ����l�F&V�n�d�ܩ�B�M�,%��7��n�	j���5q�N�fI4�Q2��@��a�V̢b��I	V1f�aw@��dR�.V/��ܷ[-[l�`;�Fk�SPї�$*Z��T��b8�mfS�¨
h�$E���2��1m��P�@�S�c/*|��L�V��ʹ.��t��{���ї����0f��}���x��[3'�)h4!¤�kVM��.mX����,V$M�����s0ԬBJ{���wI��ȾO@Tl�ҐCEM�/q�C*)YbE�h��SsLt #~�F�ov����ն���dQ�ؘ���؉7y�{��m�Uf�CR5��k[/u#@`���4�eIj�B1�4U�R�`�+oPt^H���ȭ-�z����T+-�P���<ৎ�a�ս����@vRo\�Y��:$��1��{%���v�6�Y kPL�HSb�M���j�I�G���ҥ�PѶE���:ۍf*
���g�%�D��ۉT��\�e�BL��-*��ǭ���D��Rl4�۶Úb�J�0k�	�LT[v�� ��$�D}g*Q0R�W=;�d[zީeݍ3r�SKe��&�r��!͗-��f�[9���F[�yNH�[W����Be/%�ϳE�7Os05B̻�ĦnD�CG2ه��ʻ*�k���7���P�!nf��U�^�*���ՠ���-�]=E�ˏ.!�+Ve6æu�Lʃ$�V�V�j)D#j�7�аBs�ldѳ-��>��ѵmk�t6Е�#&�o-T�!q:��fd�e�������\���U��4SX��᫖�.�F˄F�Y&�ķM�M�mY���mcn�W�)mf�`]�b�0R8C�Z���5.fh�(���ym�
T�8���NՄ�[�%��1�f���HD-Rf��R)��a.�}�f^Rݢܥ�m:��i<��L��`u�R�F�̳�1�*�z�9�1P7j�C�d��e�&�fe�91O�sh`�eF*��%Kҋ8�NL��r�VÏ0��,�R��*mb̻�-��w4�^�X�q՜��*L4V#�B[5���t�lk˹ETmk�g�v�8ZзN�Z�l�3��$�N����4�!��9	���u�b�53����I��sy�*53�3^_nW&��m.�Ce!�Ѹ^`���C" ��ĺ9�<���J�-���
���,8y`9�2���oY��q�)��;/��	��P�t�2����e�J�ZɈ2��Eʻ�]�����;�gTL�Q3�J��*�[�I�au��`��I����9��s铠�8h��|Z�`�i�cyR��.un��'1����<�z7� ��Y4��P�G�L+�w��C*-ШF���4�Vt��b訜���v��>z�_'�r��ow�G�9lS�1@�l��}e�˕�N�dU�M�� ��A�\Տ��뻰��Yof��d�啈m���]p,�#�u^[M�
 MM��_)2���Ю��
:x%Q�����Ot��s-��Wwb`�V�)��j6'F܈1*�]�d]�N��
�(����sf�i#{��.SJ6`o��29�w��ZN)�O��K�<ǑS5q�ɺ����ޚ��;j��Y}tGI�T�r�� ��k��b�Թ����Wf7˪��Ҹ.D�e�g�cD���9�7�
:��oNL�2�!�n�oY5�[-o�.�Q�:S̺;7��ݝ)&�� :�u.��ŪnN���0:|B�FҖ���ڻYt��ƻ��
Vܜ��L-кl�[z�uN8-�-� >�VMo�n��xAb� jPc��c2%]B��Pܖ1���a�| Fm�����1�XژQ0b���lQ��O%^��E۟eg:��҅.��7��c��,�{��\.�t�#��U��)x�-��m�!�fV�hMA_6{�2�YA��=��"�7���\�]tF��{Ke\���S��r����V*��K��"< ˤ�\���*�͓��=�Qꀼx��k9�!}�̼E�U��[��R�0b�����s�u���Sgi.8zҳRͽW��Uv	Y�rs�*�,��$�+Ih��^Z 7�Gnb]ϹR�̈́�x�A�����u�)��Ԩ��iN��Z���ӈah��)�sp k>a�<�cQ&]������JW�J��٬ZL6�j,�e�$*�B�w2�曱SGU�\H]�w��w�Y��n�;nU���8�f�
53Gu��zIh�:��U�k�]�v�-e�9[�\�r�C�(�m
2�$�7R���WM��!�֩�5��g�̈́�Х�A
�h�B��
��*�
��Huݶ>�9��`O�8��մ���]\�M����$em<f�N����
G	EiZ1��^��G�j�Bws�W�ۭ�]f"�5�hW5�ۣz�F��=���_5��9,�J�i��0�%��u�^��ժ*t?#y�2V�����g$&�aΣ���,���ʳ�c�@n�!\��M�^)�n�w�Z]+\ڤ:�	�*��e:�<[.�����ICL6ȣt��d6�Ȟ�2�j�cD��T(%�*%ʱGl��v3G�R^�56x�5l�=����>�{���'mz��^����{�Д�fֱ՛q��Zy�2���2;n���Y��n4�n3��l���VNR�/hw[BU���r<h���>6�o=@D����{�������`��7QM���:��y.︬8���w�pDqr���ޥֱ�6�o���&����Þ3t ��)���۹��P�yٛk�Ֆ+!zl�r�@�FΝ�����,����;w RΑ>R3�f*�9�p��o�|{2�#=�v/o����oS�s��*\��x�L�DY���]l�\tx�ZƟ>g�D���pm�j[
��������BSq�e^p]f-}��|1 *o=�Y������[��qW�G6�T�J�O����Fy���e��ohI{r�$s�Vc�*7j9[}�־�9R�C����Y/�"R�s�^�7B����
{��wF���vF6*��kW)o7J�\�� �i���U�dŜ���;��%j.�gs��eC%�B�mZ�4�AH�wc**�Y�l���wF1�RE7u��a[u�0���	��/EI��"�f6��.��3�qf�t��5��n�on�U���}��٠p��:�N��Y��2�d��Ej^��q�lVE���ۇ����N��#-]��v���԰]�Rv����S�ww�(���*�I�Em��zg'���gfl���p9���q[�U�L��*��bn�vo�����,ȏ*`���W�X{ �Ǽ�Ǜ�:ä���s9m�=�n ������Voc=��"m�D��*)�u���V�.-��Cb���7;�X�DJ�*����X����e�u0��H����$�6��[t�E ��uh�ۢ�� �"�]bV%�{%�ɯy�G��PK���<x˾k[�X��'�Y{�M��q��V���#Oz��{O��z�IÆ����r�biuM�r��X�a;�A���g2�
�d�EbuaVP*�ӥ[�6x���W���tg9�X��hv]!!�w�����+�+k�k�ɴ{y��3x&�>Hg	seZn�R�W� ���S7v�V��b�tαуä=�Q�]��̪�}�b�ت�[Z:�W�7��}�:����5[^>�u��=��/Cl��#��ش��	]�0�P��Y�v7����`�h]��#(���Q;�n>c��|﷡������q��vx(�
��  0�����Үڳo��i�I�m������������L�iO����qj�̺"E��muΩ��6���M�Դ�E*WP�[�5,������:v} W��w���J���\Z�b��%#�c���X�ܭ���zM+�'Td�@HT�����:��	.�	4�ڸ��N��V�]�����Բ�++e��9FGP��=����)�z���r]�vli�"C��w��`�C|��Ml��J�Qڮ��%�P��>[��>ū|����3U�͞�ԕ���;��C�x
�{7�.Y@r�iB�5�)W��FES�v.���@7'�����}K�h�`��|U���F��h��L-ֳw��gk<L1����Oo�,��1�.�-��.%		�9���*��7�����p�}�o�SR�l�+{KV,d��-l�ziC@�SU�ݐ����BL���I4L���)�����zu^xz/Z�1�<�nXu��fGN�k�T�w����J�g������u8�4GZ�QVfk�.plVl.�WyΌ����S��Τ�o!4�Z�����3B��1⓱H�,�y��崶h�̐+	)��TV����5yl;h\�@�{���a��.'E�N�N���ܷp.ޘ���g!���j�(
 āW�d����*;�u�<�C3�rB�KٱJn�2�R��}���e�{��@����)u�P
S��oR�6^m&4�e�*�Q�ɡn؝�տ�p�̨�͖P�]�؄�4�
�v��D_+�i^��XÐSk��{�c[�gu=��̼�7H٬�# �NbI���p����N�똯I�V�N1��.�I�ơ�O��P��5
��L]��Jo1z�洅g|8�M��ǹ���;��8qq�|�/ùS�r:U�c���B�mĖ�oN���o8���ۘ�,�3�+(!tĪ��#�L��CkmVF���!N`W�Vp+�4�'YL;c��Z�l��f��y��`[N���:�I&�-���t�0�)XPꃦ�P�e�*Ûb��������l�{[ƕ�Cɑդ��ㅩ������k�Y��0ܽ�u����6�&Z�0��tv�rI"�V�7�R٦h/K\l�O�[u��7�Vqq �P{b�`T�3��h�[�_!�!�8�Z���u�5��kQ��_Z�[�b���-Ûz
Xj �NM"�b=O�]�9�����+].Q�x`ySzvq��x�a��h���^��=uKP���oh��܋�$OV!d��O���15�ɬ��8K��{��v�6']�՞A��*V��0��s��Nͬ�AC&[��m����������nI*펕̙�:�c}0�کK2���ս�tV�F"�Y}�t��g��6�	[t���sd�A�xr�0֥��'9a�����PZ�c��)���s��ʺtH�1:�oy���-ԱAˬU�X;z9�F��VЬ�nl��R�!DGn���Չ�0�ܮE\���喴 �.�h^�WQ)���/�l�ŒJfІ��Z�5�mw.�y�Y��Hg�Lu�zv:�r��r�uvn���eڭXzT�Pf�l�*Ω5ͨX��4���B7I�+d�,��դ�ܘ.]1i�ھr��i-�.��h��ׂ�6�oW,��ֺf6�<��e��j��� �G�lo+�:��z
}�Y���{�>ꋄ�{K�D�v��Z������e�c�맳�1ـR�F�[�;�҅-}�4H�þ;Ñ}��]񹧌΅R��_��[�c
���`�.�eh��+��y���[u� �k.>R�O�ٲ����e2{$�Q���1�^��V0f���X�蒵��W�i�
u��ëI[g�?�lc��̲���D��Z���mKrԷ������Q/���L�n�%L��L���C��gg&� h�h%,^a�XT`�����H5�4/��k��F�$���;}���y���S�!��0����_#�4D��[�M>W�JT��}�����D}�ILwv7��U�ټ\��-b�Z���
7N���q�-�Yð�-F�rX��Ƴ젙\���Z�7Os/��Ք�6�o��z�fu�:r�A�&��޸Qz�t8^u�ޤ1��GsW�/GsT��>�z�.zؙ��̬�v�7v$�8m}����ph}I�Un�x��`ѕcV�"�U���Er��3�#Jv��r��u�)t��7ݽ�Wk;\�[��#�J�`�r�l\��"�S��<�6��:��Ij>i"��(��-ݍ���خ!("��߃s��^T��b�-9ǚ��������.�\�V.���u:�4M�Àiˡ��bo���!hP̑�7B$CM�c8��s���2��A��V\�]x^��PGgc�U֩��ҵ���z1�o� �Y�����]��c�޺�Ѥݑ�KCm<O�7�W&�'&9�R�Ҡv�;2�t�@R�����]Λ���֎MÓ\�%bN�nP.��	C2��YL7{a��v���l�!y+Y*u�)�}���5-���sW���Z�z�GD�����uM��Z�v�8Y)���5�՝/C�%��+K���>�4Ň�ԡh���5�e�2���W#}s�����\��8���R������s��M��ĢW�.�2!Jj�/*�QW������e�ծ� ��/��; Ays�[�|��+�E6eu<��1Z��o��"�TAB��~=�B�S�;��3��sF���B)�$y`��=�k,��%L���J�N�����;/qU�mG|(��5��[gv�i��C.$�u%YX�Mr�6�«���ț���-Ei(E��X�!��1cN�sM��c;�h{*va^����Z���Ӡ�F��s��W�\N9m�K_
[ 4��+���.�Ԡ����B{�s��YX#�����7ˁ�hڙ2�E�d�gd�v����2�Q��8��s�fβ0b���s��wwlDAw�R��0�\r����ț�c�}����W;�Vf��c4L��7L�Y�����8�����9�YGud]����8I�KX������t���.��A@R��(AǱ�*�n�����+�s�ȯ�,:Ś_í:�ڰi}�&u˭8._D�q.�q�s��\�'2�Zd�z���Nn��]�waZ#7�VB�^�<�A�;����ar6khWj�y�P%J��P�������Qݦ�^�!��N�H�WہTUa5���"{� 8Ia=�:�R���>}d�ݨ�睫t���̰��͝A9�����Qҩz�lv1��|eA���F�U�S7�*���K�������4bv�5,�̣���yr�h���gT���]h�"Uv�v�i��	�*ʰvQ�S5X[��Ad�9Sv�(>;���Q:|v��� �K�Y>P�JL% +��2�԰� zA����h�b�Ŋ�Z� ��ڻ�{��u�jQ�d�k@P�+��k����i�D��i*;l7�ځ�-��#B��H�7�u�Nvj��,s`�7^L�y���0�Uҫ��g:��9�ӫ��s+Bʍ�Q�l����6����oo�À�"h )�L���o&�j��ݡ)R�A��W����jK�*a�~�JJۇx��R��X�.�]p�{}���I�_8��30�྆��T��A��@��'��]�!�P�=��V�
]�^R�hޕ��ΩqrU�ENl��¯�u|�Z�j(W9[g��\�Vk<����P/v�R���\�i����3R��7+��.g>�#PVM�a�bj]%W8$0L����o�0RǕ�<݇j���Ը�Žv
JJы�մ��8-���[(vp��2D�q�s>V7n�b�'<�,w;�d���əW�*Z.���K7��Pb�����7R��)KL}��ejk�U��_[MLn��9��D�
����&�*��B�m�>��5)L��N�N=Ҵ��ϸfJ:Ryln!O6ʨ�^>��6��l�{XJ�^��U�Lꁲe��\-9X^9A�LooVj��Te�U�p�ݽ�\��}��m�m����
Ԫf�+���"�1�%ũ��Va�Xp_7�}��9t�?ws�}	&�#;�plN�:�G���_g
�p�#+�j�:_Rp�rw\R��锇t���M��$��-�߾���k�r�����! ���H@��`�՞��ʆS�6����L�O;i��G����yĩ�w��!!���NWl�U]}/'_ˢ	q�j����W���\v;(݊)�x��n�D�W���>�Wv�͇b
diۏ]An�b�>����Ԉ� ���S�ӥd3tk9�:�og�9rs�?mlڒ]����#*CL�)U�p}f�Z5�15�r��2m�ۯ��̖�r�/��"B�KE��9@�܇PA���}Zqfۥ��o*�i�Oc�v0���/�@A�2���(UWf����|pgY�·n3����X'KTqՓCo�fu����K!ֳ+f�,8$���Y����Ŭ��q��U����
jV=��1��9�GT�-����La�`;�ZY,�\�����n��S�kYv�Dm���]Q�c�Pз�<u�ГUwF�փ�7v^�ϵlU��,�Ѳ���b�;i��N�=�m��Lt����8�q�`b�M��j7��x�;Q�9�[e�j���ѽx�m�8���v����K���	�S��*�hMV�\�b�m��V����#����v>r�[ڍ,�q�p���V��w����}�����)��Q�2�9cS���d��όYB�+�킐��;;�o�.^!�N '2�(�|��q�e�WO���IR���C����:kq	ss0���Y]1G��և���&�Ov�WP�
��8�c����C	N��wܴ`���X{R9{%�����.�qu%��]z�\��zi�s�-�<b�b�wk�%?���X�i�FW"����ܦ&
�{6��(���Avv��ܧ\+*-�]3�����j��t�X��Ø~}�8^��+Q��Msd.�d�2�^�2���&A������Sϧ��4�H��e�8oe��;�6�]ӽ�L����J�-�t��r��l��+ݬ�ut��M.-%�� �uԤ��@��Z�]�RƸ�|;4��'V��	G���v�4�#!�Y�E��3�:��pWv�ܐ��Dv:���ߝ��w��6CK�qg��mJ��|���t;gusd�{��j;�U���ۃ3���s��+����N���u��T��1�V��B�x�n#���ѻ��t�o3�i���"�I�ԝu���Tܪ�`�Eb�٣p#A���Y�3���*r��Γ)�u]BuF/ZY0,͐p����7�(u���>wݴ�P�&(�u�L
��!�^�7�(����V��v���:��uktj�t��:�U��}�DP���Y ���K �����P��N�G}��m.�?99̮�pX˘�\�r����4�)X%mb��-%ݕ���-#��R���jMhq��Vt幰L��^u�z%:k�¦��Ql�B�S�K��J�r�	{�f`�uu��'K �D:̗�!���4��
�E��)=�U2
�sG���t���x�����+Q���̜.�5��y!V���un�N0m��XVk����5&��u����{�J��*�elt�T��G*B��R:/W7�!x�� R\�Y��o�p�WY��<��E�v��Wۧ��N�w\�|�Ƶ�ve`��S�[iI���hi]�Q��������㗊��|�������1�I1������G�JA	����l{��T�.K\�����'a�`v4�S�J�HX�0w�u�fҵ@�c��5(Z��ggZ��]J�_l��V:�E�l�yV^�7741W[-v&5f��7� 3p]8�!GF��gvWN�����ռ���oX4���&ӷ͘��rP��Ⱦ�l�i�n�D���:k�ǒ��.V"�yM�T=���e�}�5�Y]�S���#������]\� /E�a�\j�W(��'(�tr��0�[ME\)�c�Ak�4������������҂�_E�6�J�����rNY��޼�ġ����v�\sJ�Zu������ي���k5!3>U�qxE6��KUe���:�eo-�I�d5�Ԙ�W_ T�����V�[ZiR>�����7��&�3n+��"�'K`u��l�vR��c�kfPL��\ t{z���˴��R������A+���:i��,�Mw2�r<��j'��:�#٤��7k��o����k(�֥\z���[k��0R�B�־�61���G�G�l�8e[��(���1��N����)��@t�� ���ox.]�FRFjA��ݔ ��ܬ�Ut��i�c���V�V�b��㾍���r�:�C{X�r�Kt�\p�/[��Ff�Z�]���q�Õ �n��d�l�k4��2��y[D��M�y�۩��:�Zj�<�&G%Z���Z�Wav�-W<x��ӱ�;�ghߎ����4��f�@k�vݷ�-�n:���A�1)��E��c�S�R��}�Lo)�>Zl��.��^��we�T�:of��*ܬ���2�v'Ӊ����͏JhN���ޑV$�9ݵg���Oj�1N�B�G�j��9b�+��Fv��陜��]�n�ws�����}��;髨�L�t����:e&�,��TV\p2 i�n��r�wd@34�qb��Oe�h�:]�ʲs���G0*d}ϲ$�=W�M�(1\��㯌Z����S\�"��>G&#m���Y�xr���Wy�{�0Sc�����Xn��
�	�}yWݑr��[�ڧc)�m@�ugo��X��"V9�\CQ�(|�gNw7^�V)	�뭦[��K3�I�`s*뮴Vd�\�:�h���NI$�xܤ�,x�$k��DV�X�;����!��>�#A�m����E�НL��2����� �5nm!�.�G�^�V�YB��B��b���]N�/xY�fD1����r���d�/F�K���]v���.�a�X���ب��}�2�M��*U�kT���[�Ƽ�L\�]��(îV�7�g9����rm�qKʖ�|��G��tʢ,��G8��������ܧ#�{���qn��@4>�c2�>�Q�t�ѐ!��LD�p��i�M;&��f��^�=�F��k.v�x�6-��m���r�O��ھK���V�������=��:а���k���ְ��%�G;	�cisp7�B��.���z���~�b�we�w�ۭ�m���mF���Q�^Sg[̱����e�O�`u��$/�^:�,�;N�&��e��cTټ��iw�ʶ��,j�㼆�)�0S�ה%[=qh�+s�X/q��w�"��h�%k�K$�+�]�� K7��M9�L�d�y���S�+,V���5�/�{�f�^�wKğ�3�6_oZV]1����Y�`�9��J�cy9s���S�OV��ʋՀ췊���:�\�����}��J�ԓ�XpX��z��=�M�c{8'�0�cܡ�:�X��y[p��i�ip9;�*Qӹb�W[��*�E���ï@�c�Rl��R��.k�c�Z=潜��$��5t�`b���R�Mq�{ݹn39d|9)D�'��Q�b�n��+�ݩ�U�<�Tv�7��J���)z� �L�V��%]�S23���}�J|���r�p���f>	%͙�/-P1+r�*�a�Z�ǒٚ��^.���[i��:VW=2�q�x������{r�=I�ۤ5j����j�wl�(U���i�;�;�J�7[L�t8%�����X���'
��g7��r�n�*�#��I�{ugfֈ�HY���sB�
�B���&�[9��[g���=��OKƦ���eZ��o�j+����b�3��g]C4�$�N�nIW�Z<\p!Ijy�vk���]�1��pX�;؍!W�k�:U�����[��M��eϵ#��"����aV����&���Y�����5e&���sKs�%�Uvr��/B���5���3��5:�`:ra�Z�%Y��}G�m��]Z,Nַ�AՉ�O

�+�u>�bS�rԤMam:4jMu���rm r����ݻL3]f�u��%p'"߷���C�N��X��<�����K�ʂ]���Wۧ����ӡ�r�� %�4]ҶY�����[�a�����]�A��(��ޤ���y�Pu�E;�cX�Y�VgG�W}��ؕ˧�F�EAzkY�����)}��5�mQͣkE\Wf�� �4�W>�t�.���J�ga�����v;�w�C=��H(CO���ȥ�oL�H�6C��æ<���YtN !X��/D����͝P��o)*V�&]�3ek��/����"�{���+w��(� ��W��E)+A�B�+����y�։b����푆�[���:8��'moZ�F��u����$�yI�R�W,�����vcגV������l��*\�����i	�Wt.�<�gq%q1&��;O�y(����Qa��07@B�ɷ\ݛ�P��R4�"���Sy����[6]���}�Q�S���8`��m�'��6�'A:�����je܎Q�f�z��Ё�<��c�M���
�5Ĳ�+=D�,sC]n`T�yi�@�1	�bg��\�����=��&=���9��gZ��:��r��uO�ݭ������W�E(��ʜNQ'���u�C��H���o�i��ݵC��t0���e1�6W\uB��f�է���`��Sb
���e]oV����ه#��;����ui"谒ؔѵ���..p��Z�� me%�l��fZP:�!�q�S�4(,���-J�ۄpu�D=� YXC�ː�ѭ�:VgG�^v��l��L�)�wL48oF�8�]'��)qs��;��[�ZO+Q
�}��5X4���]��O3�!��a�$�h���u]qi���]Z]�s�s{C�����б���WH�-NP, -;N��:&���m�}��$nM����M�92ja�9�̼���S�V���b����y�I�uoq^��7{K�������F���֤Tp�ux5a�i�p���-��h���5����T�}n�cd󫥙v0̦M)wf@�r�|x��T�t����-
����-���M���w�tB�J`d%39��_�i�x*p�m
�6�VFP���J3if̡�]�v�S��E��pE���.����&���M�ߥ�b� ��	&f[�u.ʋ#��N�gW6��ܺh��)WtWs�P8��6��w�kmPtK�q�J8<o������u}�]X�3�����Ԡe5Ed�J�]���z���a��I�Y-��	�́\�	|jRUJ��g}t��;\�j�.��.�b�)4�9��dJ������àn�@͗B5�̳����"��p�����4�"}{�nw2d��I�ګ�K+�f�Xb�p�Z�|�X�w�μu��W���;2fe;��r�i��{@�%B'e�%��f�G'�n��&;ᮺ��G�y5����>{u��G����I^���^vf$��:|�R�N��hSq��׽�|.3t�]`��3]}b��"�:�:���ܥ�GV�u5�4�V�+�Pu�F�[�6�}�#�� ���u�o���K��7g��;x��ЪZ8��(:+��(����iЍ$��!��fS���]S2���]mr�Z�-���H8��v���aE�Ej8�,�~�״��l�a������0�:���6\I�{��t�+U�AM������G�e8 ���Xq���V.��Q+�)�\��ʏ�5"��w�i���`_UCxĩ����X�Z�ꑻ�A��죐l�P�Z�rG/�Ļ�ݰ��uaff��2�Ε7���Tm"�n�:�ܧ�9s�]%����[��;O�8�va6���ض�t0ԵO`�` �7���'�(;��Q�{��N;z��0Q���n����_N�U�m�v��M$������a��,�XO(kz8�ܥ��J 2�m�,+�z�����<�W�:�����>$lb��g��(���� h�W(D�J%��]:�o1t�amc��:���;�T��Y�J0˔b8�_U��*�U���!y:c�$���%�M^;�:!wݧm��eڢVPih��7��V�J.�vDWٌ�&�+^]K���i��;s�Y+1;k�.�e.�$$�h�2�e=�)ݽ��)��)���9��g4�ir`}htY���3J�}:GfB�씦3��gkW�u�4IyP�D�|�^�鑗�2�hRN�����88�/*�[A��1�TC��3+jR��P�g���k���*��B3�@��
��}l�$��n�V�m���U�"v�R�Űn�aݹ�Ƶ�r�j�=�Y������AV�to�n�[��<N0�'Al��n�ݬO3�����\����g1�|Ji1�T7k,qBmWtT!w�:�'su���.��k.��ޱ�+�󮊯��B��������2��uA��_D�¬Mݔe�EE�eqͦ�Uڕ�����y��:i\�v��|>�iyӗa����V�4�,����� M"2CE�Gۏ�(�+�5I��ju��rP�ٰI+��z7�1z�t�Z\ �Lm��eVGÅ��Q@[���8m��$�ݸ(V]c{.��q*g��K��f\k�2-|Ue_.�(���oSmd��L_N��"���F��1'�6�|<��\ˡt���5�M��ț�4Lz�68�q�H�-����;v(S��vS��³Yq�G�^��h�R���U�Sgw��S���D�d2nnV�X�+^���//lfQPԀ[d�C]���K��F�eº��� ����Ĺ����5*g��JIÝثw�-Ep~�U}���W�}>�F1+���\L���e_�̓�L�k�I�!=�f�q�=~�`Ć�*?M�V;��}�h��t�U@J@��"l�����}ƌ��(c�
��1�_* U�I[ٳ��Bh5'[�5�V�<�gx)co^��ͧ�]l<-⃱u��p��_c��م�a���+��F�M�������̼b�.�Mݜ+���YC�r�����tt��"v#�z��ӊ��������Y���#����)�����[ͣ�"<��7�e�UXq>�Աv����:�k��;�q�4;�%���GJ�0�3�eaW$Β��S.��[c"�_fHܺVP���	<��pg.��XnHԕ'p�21�E滏*�l��̲E;Z�A�r��)EX�)�M�w��C;()s��ݱ��`�(�/�Yɥ9���k^M�Χ%q���a[�����ݞ���k�Ws�^ 9sf9�])'�V	塂5۫��k[|�Ux)�Pc\c��7�Z�_L[DmQ�9�̘�Se�|�u@��ң@v,�/�M��80H��h��,�ieh�u�2ZS�fy�qfv.է[��Q�E-� ,K�)����m�^-[a���%3��w���{���ۼg��b�e>߭�C�F����\mgR��.��� �μR"�;�c��@�Sjg�e���1:�pK 1�t�-��UY���:�n�\�Ā�lu�yS���NÒ�fW	6���N��nLU4c��Mf%��[(վX�V��9s��w*���v;�n��� >	�*)T
��kA���$YP�ũX(�EDb�*"�j,�$QV�`�VU��J��I"%e@�E-`�����+�(�(�X�"
+QFb�`��b�"�XH���"1T���E�T�PeAe@+��ek�VB�T[eV0H[dPR�E��QDb���l���D�d�
J�kH�E����EX��b��2*Ȱ���F"V�DD*TP�X���F2*��A�UAEAbȢ��c�E���*�QV(�U+�bŊ*�b�QX���lTE�Qc("���UD"���UAQ�T�H�X�E"���(��EQF,DD,bň��Qb�,KIUR�+D"�AH1EB�5%��Ym�Xɵ�u��u���cN��R�*�M����� �H��#/W& (�w�$ڥ��A�յ0�1�wǪ�-'���VY���L�)	��`�6�����������M��lrg�c���EY�����L���np5�<wa��%�����"��(KttT��U~��ђ.��G=�I�&7�aچ��KP���^�y��J���"���W��:ePP�nyh�ᾃ�{�'v�(S��*�.���q�j�{�H�(rj�0'w���CQ3���.�tk�߻��A�j׎|E�b�R�/m�7�LމWvѴ9�	-���­e�v�l�W�����ΰ`��a��Oơ�
�w�r��p����3�U}D�՞���l�����-G�,L^��DbE-՗��%�%g	1#K'�{vCʡ�VƼo%dW�y�}l������(|t����/e�
���J�����L�v�R�����f�M�Z�m��v1q]��j���~ۆ$�����x�ܮ���f�Dp�s漝��]���]��=�h�:�Ϋ�V� 6/�l�N��P�ZpNw�3�o��QTL��L�����g7]�/z������vS�=yڊ�A��r��Z���96g����a��`���A�0�y9#�[�,*#mq2T���V��`��)�H��n��>��>�O���wғ6F��y�u,q�]�)<r��q��Np]�����<a1�_pTpϫ���M���610G
gb�\�a�O�iv�ҧיe�k|��� ��-��W�u�e���9�(�ֳ���<��ݑV���Mc<O/7�׍�No���M�ϔ�2.�v;(V�.TX���1&tT���US�VL���k�<g�+�'�Z0�+1���&��k�D��i.��+��8{�s���C���<��8�)�D�.��,=5�pv̢�SńH����ԭ��A�������#�_z�G�c�8o�={�j2�{��/l{����IP��$�4���g�jA�4�������{y�
6|	" Y�*�L��z�7�vnH�z��ߦJ�>�N�O��I��ir�Z�� �9O��w�؃r�� R��-I4���h���^utu�|R]C	W�kZ}�kKZS٘��ܺ����]Z��1��P��n��j�qD&��E��t4���c�5g�~��z�y�/TE
�l`�!�������)[�w0�TK�j߭2��i�z���\>�Ae'�4U��k�&K�.t�F�ӗL���R6�[�/<v��9��ڣ�c0gw;��,I����ל��gSM;RI[��hj�^�V�;�ɍs�CЖ��X���+��z�)D���w{ێ�Ծ*,��x8Z:VV�Je���8EMtg"�k]$ӛ���lN��n��J�5�eg_ |�f�W{�ۊ|p�|�=�x`�u�,(X2̮$�E~��5�t�b`to�b�%�{��v��yw6O{[MA�����-��-H�֛0s�g}��*8"�X���0H�h��Ic�ۘ��l㹷&+,yb�z�j�_�~u��n�*�.���>���X=>�\͋���ѽ܎�����O�����mڲ�b��ǌ�[Zn�)p��(f��X�����n�hY�(a�)߽����x����p�]X�tW��X'��:�KC�yz����xݷ4�gc�����V_��)�ew �ݪ������he�a��-d��u-*�2λ3�'���vu�9>P���2�C'�7')�L�P�Ԫ���0��0|�u�O�;�S�q�(��=~��Y�i�%D�ز)�Cf}6�����L����2�Q,�OW�.��I�Ӱ�B/P����*�T�I�n��
<��=�yJ��BhvE�u�^��wS�����@��0�x'ZI��.�R��wO:��C�#�R������lb��3�Z��u��=��n���7��S�������H=�[Б:�2�]��ռ���vz��#����|1d��"�d+�[�+��}���[#�L��+�F�Z��v����Z���ֹ=���g!Y���?{����B�2�)�Gܙ�v��<�Ox�lk���� ��/�%.�ѳi��*o0Q�ʘ�d���EC`@�*+M5��q�(2"���A7w~�k�Ѯ�J�,%��[�8"��*j��u[�V�3�Ԣ����UEἹ}�n:���_`g�V��P�|�U�3 7�J��P��;�jݚ� +=^ŕ����{6H6��ٯP�������U��Ȇo�[Y�F�ϵ�ED0��u�,��7�r��W���N�����Q�5ZC���;tՌ]�	���5*�\����m1�����h��y��[o*�o�-��VpK�?t7b눯Z协*�Z��ώ��Ào��X�����W���gԻ���S(�\�k"�����Z&z���D*,��7c��w�U��9s�]��)��j�/"����&�{���K$�5�/����׾���W�Cβ��#.6*�[w4��k��y�ލy�]������oT1;��,G��{WC��g���O�X��N�Gyt��`������<_�V�����TD�k�&�i�?�v�m�+{ެr�����WV�����K�[Jl/R�}lx��+��\�\�}A��@�-�}�->���r��ͫ�]��^5�s�>����9=��������_@#�s���u/�&�`#|%0xߝ4��N���
�#��j���T.��p]7�|_����6����U���zǛ5��y0H�9�����k������s�}۵U3�U�P����y��k��WZ���o�^tA5ф���Ȧg��?S{j��y��y?�in�CB=�G?_WS�2��褛f��(�ypQ����)����%�����1��6�c0H\H�C梻��N���}�M�5׃e���OG^�$�$*x�A�z�,"�wi�6%@�L|=E7ī�2�{�g�`}����J�\��`w=Bö������
�Hrv>�+�h�L�Onϣ��c�K���o��V,���^�[�Ñs�{�ts���8W���+�Z������`7	���]�;�e-=}�7�S5�R���t=��#\�^R�V�Y�"��w���8�RyoU�ߺ�[v4EW�j)�͊`8���Q��,�En��;�(v+}p�'�`�]u�A}Q��6���U�jIM��[�YHv�rܩ|�Nƛ3J�k���%srJ����Z�w��ـ�����n-���']]��Z��>��z�v�Յ��}�y�v����u�@nv��4�W�C�Ro��O.�_z�ޮku���7_v���{\�J�v��'i���V}�狪��[���<�>���۶{�/ß�^��öz�Sw��ÿ�6:Z27����VB�9{e���8ʗ���Qw\��P�:򠬯H�z�K�N{�Ny��R��ީ�֩�����ۮ�z|����Q�U}lm�;|���*9e�ʞ����F�q{�-M������YE�b�������8u�6[S��Ì7���w�p���f�����/T�'��ͬ��g�΢�,�:"�_�j�@�};̸�m�2�ؤ޶����N5�=e�B<�o��yѝ�~�Nؖ��\����Ob��]X�Zxr��<c�j*�Pw��nL�����񳲭ӵ�����`��wt�!��j��0h�	�RX���o�g΀-١�uyٴ�Ψ����͈�p��J�ʥݪ�h���5�;�F�_L����5L�OL�y�l%�}�+c��X7oK9�U��˺o.&b=$|��[��ܳ!�R�+���r���A����<�7�����\ybk�u%���˄j��GQ�I���{�-)nWB%A�|��ْ��΅֟I���;͙��qM�@e�5�n�r����Ү~*�pi��������z��۳�k�{��ez�A�{��q���]xXny�d�N��_.
{֒��=�7��|����}�^��[��4� {��ȽG�/�^yOy��g��M��i�,��c��O�`�;��A�X��A;�g�U��y.{�V�&cn{mH������f�J6�ϟm����k��$�6#9�`��q5Gv�X��:s���ͅ���_ec��=c*K���{$���r���o`5jw9�f��ݞ��9R�4��ҕ��K��;�Q����+f��@��w��s��r�}Rz�/Os{��7EJ[�����q�����}Փg���Uq�=�pTr�u��;�wޏi3{}J>��S:m�A�+��9�_�����_';6��H�����Vq\�"!�T��ء�=�N�h�1�Mk(�����θ�.���
ξ�y���@�Ư�T�9!�����9�K6�/�y�c�l���v�^�m�ɗ:�����䜨T/m�㤍�.�������@�c5��P�:�����oK�5�{�aͦ7Sܯ^��sd����s�h���(\�/�߇�%����y���7��N<:�w��Ȝ�}{���1�A��\�ru��_gO}kk�)OễDs�ק��I�����\}��dSH~iI����t/nl�h�B�(x�{f�wi�ϛ��8��,�r�>�N<҂~]S�����콛�a[�T�R~{ޕ:\�ف�f�?\��e9�/�qPti����KLW�z����;�6X�]���W����K���Ҙ��F9�h;�t2�nƬ�g��N>n3�1}�{��������;�,k�Б�`���>Ϝѳ�-��4�|�|�ˬp���Y��U�w����ݶ�1-_o��*y��aHDS4gs�6��S�hE�mW(�t�L���1`<���jK4]�X�+ٸ8r�&�W� �g<?K����|j�-�w��bt�@�NN#3������:��d�������(fN����wC���j�V�ڪ}N�h���@�p��N���0H���8%������צ�ȏy��uYhp������k�oe��o�!��@���Gj�M�=�^l(=�z���J���^�>��_�q�����Eײ2�����^�ɝ5޶��z�Σ~^C�hn�dg&t����'�����g�����N~��7��&o�u�Z��G������x�󂶪��pv�6i�OJ����~�I�t�J�d܉>]�熺g��r�PV����LZ�_[WNl������*Sc5�Z-߸v������F�����r��|]����Y��9ýZ��[�U'<�)�a�U����Џz<�_W;Q�Y�q�O���4��T��ʹ��̌����NzeOT��0�q��ힻ���w�����c�q�ٟVM����+տ��Xr*H��@��>��f�5���ۣI$�e34��wZ�0�jnaOz`o)��i�x��Cʢ��X�i�ڬn�5nm��Ш ��!C�a��]�,N��ݽ�#�@;���/�3��35�b�+�Cv�׻�t�̽<�(�-��2�����͎A�):poX���'*�_^�I���`}��	�>�{ڨ�o�T�*pރ϶N�Jza��{jx/SeW��v}���.�q���)v]�oW��S�ewp��7[%͊��փ�|W �i_eK���D��A��{�^�z8ws�g���>cv��㥞cޯS}�|�#�I�)��S�s�ϳ��:砮�����ȼ���T��I�?aH4�������v�	O;v��v=yl`�H/X��֛�O�ʰ6���ꇇA�#}�wRR�/Տ��yi����[����ܽ�ݣ~>�������8����,��������ʯ���T�'��Qu)~�?���X}����2���[�����������1�->Rp��T-���o�p���z��T�-8�~�;w�F�����n��I�������1kech[��}�\�|�p=ڙ[���k�o�8
%*�9Ǝ�GD1�[}��i�E��my��յb�v.������^!���T��K�e��c�;��u���J��7E����|��<��yʌ3fWv;Ⱥ�h4�!��C�T{�4#jV@q���ˮ��z�>�y��3 ��� QL��
����c[��c+i�P�l��# i�i,K>G����F-9�1�b��`d�WڅD��Ǘ��e
rl&ݵ��YX;�b�Q�J�7ΐ��3%N���:��[��k��@t��n��]��*��'�����֦�����>��y�f�y�U��:{I�|�p�]t��a�ܔP�!g��}ݿ	�C��04��Y��/�e�Ok���`��qui3 TL��5�����l�G(U�[�k��guq��0�+�
[/y_h1� y	��������Q;�;�T�]
r�h�\"��;fK��f#]v�0>��5��W������}}���ƹon92���)��hKoe--�\]�x����a�754& �e;	4#���d�W02֝Sy1D�3)܋P�v��<����.EИ�s�ޤ\�30�D��;�l����U�2�z%�547�됂b�{c���/�R��
���H�&�����۝P��wL޲��Q�/��+��2έQ|]5e�U�B��YnH��w59Nݧ)���Д�Wg�K�1�,�T�N0đR�*�ӡ S
̉������Rr��ZD�T�����%\������ڬ�l��Թ0�k����}N�W���	��rh9����)�Rv���k�o��8�Z���{J�]���ݺ���t׋$��½�,�hc���,�U/��^J�7r�o�/�kA�&t�ܼ�Agvl��l�zsb�}u�L�u&��<r��l�-��C���:(:�c��n�j��GX�d;�p�ø,ɥ�S��t�K].]�Z˫��T��0˂ʻrR2�pc�m�V�uG(�ᓲK�z��Z�+���r�im�S"�ݳ|0��U:�����3�wʌ�})�G�o������]Ɩ�ٌF�}��޵� ]��o�i�,ǲ9��Cy�{�$���z���F�2UB�v��V9:yAءr�&���â_ex��U�t�*6�Vx�b���Lncmn�x��+9ec���d�vH�H7�0ܶ^ǵ*POn�����q7���_�9iL`���x���wݟY��u�*��"~F�ө�����v�rR[0�ubq�7����v�EU�Z�e[%�n]h�Vw�T�D[Tq�������e��-{>g#lx)�]G6�}(��Y�ђ�#j���-n��@7Gc�K�mɯ�/�5���	fR����)�X%D2�YI���`�fQR+%�X��8�.+��w>r�oC0�,��]:Y��.�h�7��ZӢ��K���g>]gX�u�(�@EDGIb+�$Eb"1AQ�� ����������"�ڢ�DX�EAb0X�XEEV�b��`�A��,��E(��A@R,Q�H�T�$UQ`�
�V$db�PQc��Ŋ��DU$�XT��RT
�EX��`��X�F)Tb�TR***6؊��b���V(�AEQb�TX�V�"�����(�"�R҈Ȫ�E��ȫ���[eH�X��cmQX��EX�-�E��U�J0Z�@`�V1�(*,b�`1TV(**�����z�`�,#X�*PX
,F*Ń"Ȉ�(����"���aX��TUEAdEp�EAb+Y�*�*�%�DVF5��(�0X*�Z���L!X�QA���0�F1A��UEAQAH��((�"�Um� �,�>ǆ�5����˟1��5��+e�!h-���7Y(»g$M�kxWN����Ż\�_v\QܾʶI��ކ-�y>�-;��G�u>[�5u.���GM3)Ӄ@���W����k[Rw����y�=����|F�.�,-}�o(۷C�<�|�z��s����-��N���?59<��3�}��,�6PԝKB������n4��]��'����\es�����lT�~�IJX;�η�?W^<y�Ff�����y��r}�1���|%�ۑ��/qۄU��\�vwz	<�d�^��C��@1����.]�΅��O��k��=��깲Ջ|�����[=!�Ws��x�ж���('��S۳Oja�%�gks�}��K~�����Jy0��'����Aѧc����*�|]_d�/6w9�S���'�7�LKw��qp�����U�Is�wt��v�>V%J�s;�1c_b1�9�q��y�U]�W�<)���>D��β.?aD���o-����~�%z;V$�5�ۮ�AXY�U1�xuj��r�\���Q��/�r������2��NU6�7��_��u��$�=N��,�kʘ�U�[Ȝ���|�yn� ��0��6�_u���OPW\oF��T�׿�U�u�9&<���_�h)�J�g�+�o7.��L,������>7쩫�2}�b��s_Q��H�҉S�Qm*��S�W�d��fw���,��oK�g��{�8��ͽ.�����s>�U[���ۺ�}��<�}�zߌ���b�K���f���g\{]Xp,��R!�_s�#�yph�����Fk6c�o���&�j�9J�0n����]38�{}#���U��.�Ǵzc{I��/ۏ��S��FY���G{��}My���wJ�����}�GK�P�k�򇧁q/;��7_t�<�wuߠw'��S��d:y���b_;v�c�f�z]��sg˹���k�a�ua��5_M!��iI�����z�ʼ��[\}�r��;{�^v`����7�W�~y.���"PcJO˦ǇqE�2�x�S��CFU8��є9�|��Q���g.���>�sf׸�P�F�nP��v��ۨ4m��fR��s��9C�zn/I��T��N{�Sz��aB�wgX�z�p�@*��V�+�_6�-R�����R��B���w��Y����΢�>�﯒���cgy�{�������v�q��w��/h�����!V,�.F	Cq�i��1��9>�=B�U~�~O�J��6>�İgx\sȉ��^=��i_�I�v���PQ����C������<�O�x\ϺxԌK��y㏱%՛t�<�6����u�h\�^������R`��`Ʈp���>�Q�(9��}��ϻ���g2�`(t�,�د�o4eH�xx�2��k���2��/'*O/t�^Q[�䖗=AmS���[��^6��R�6�<0�W��\k~�dP^6=^�}���Խ��;޴[�������1L��@Ů��ݒ��\}c)�<�O��go{��k�豕W�W�����e�VW�V�������A͝~������yyKڵ%3Kݛ;��k}��Vv�&_o�nW�z���[N�Ň��,���H�h�9�ͅ�\γu ����c�X��{�]��@������t��Ovx��g�巼q�̇�8��)���q��^�Se��;��)����=B>� @�����4&��Ap�a���1�g�v���$���=��@���)��ݏ�}�������_�ΰ[q���/;�j�B��A�y��������"��5�:7&������ʘ��^�|�z)��=<�р�����S�2Uo��o�ﭩm�v�gӷ݀>�_?G��KS��>~xf��w�W�����}��<g�s��{q���f�+�'����κ�R�9��u����Iޕ��_w�����?B&׌t/O���ٟ;�L��$��zu{n�-f����v��~��c����ƣf�Zz�?�q aς��'Xq��CL�&P�{�
u��`����� ���[���ݫ7���n����>a4���O`{�'Rx�-C�5�@��3���8�S�v�sX�RW��aĒ�F|Ěa�C�	����?B>����~����ܾ������2m:o�:�T�3��VI��{���`h�0�LZ�wd���6��&��a������<dϽ�:�0���qy���7�r����y���I�8��i�d�=I��0��^��):��$���;��'���r�<dš�{�%d��q�	'Y5�~�>���E��o������!��뷹o|�y��	_���C�l<�&P�ٻ<C,�E�_{�6�ԝE��`�I�ɾ�Ւa���6�C���a���a�Sz����w]�3�n4�Y�\���ߏ�N���A[����s��Q�:��,�:�	Pei��]>�9ǵ�c⾧���\9%�/1aoDwd���{��륌�F���b��7F�r�,79>�,����%1�ح�9���| ��;�ovx����X��g��a��3Bm�y�d�0��q'Y�&�}C,"ɬ�yi8��M��6���l9�$�5����ҬO�������y�ҵ��[ݯÏ�m&���ԓ�;�
ɦ`d1I�>d�8�4&��&u�XO�k��N+$ϛ�:��Y5����������߯�L�r��i�T#\��u���.s����Ͼ�>a�|�xo�=a6̰�9���$�q�CąCl0��u��m�f�2,�Ԛ;d�,'ω=}�����B�S����Z�x��k)��(dݧs��C���׉&���q8��|�,<�{�'��L�a�	�h�`eņ��'a�Ł�'Rg%~��#�_�-�N����}����	d�O�������'S��`u�1�M�d��Rn�>g̙C\�:�q���pVq�|�ŋ'��!�ş$��޺����e�e&�W��<	��W�/���e$�F3���d� u�^$=�7��$����!XMw���2xÌ�ZY�&���z�n}���C��yq�8ϼ�;��{�dʡ|�l�E�LP>@�&f���>d�;�i���<3C�'X�
�x�S_{�u�Nn����4��{�u��0ι�����>���/�\���캬���L��$�E��YN2m��ɫ@���5�s	���	��'�k���+>I�nv��M�����0�	��n��?�����w����y�g��@��y�8���E<��:�d��ਲN!��Y9l&!�qi>jE����l�b�{I�l�a�>瘐�>dW_�M,LIq�����I�?}��}�T��ݸf�&��32z̠y9�!Ԛd�,�l�0����IԚ8X�I^ z�̞�q��M:��!�zo�0�vfy�OKaY��	����ۭN�3�m��]]۩E�i��t�
�\��5�谎5�349n�2�xi�Y9`�m����#|t'@p]����<k�eh��뛹�r�V���v�aA�'�xN����oz߹�� ��*�y������?�P�{�Hu�d�<9���$��;C�m��{�e��Hh�1��&f��2B�a��I���Ri�	ư=?G�>�B����F�Oa��E����a����0���(,�L��}��`u5�c���Vh�pE�u��!�&�`k��VO1l3>�ug�����ߏ�W��pG]�ު.�?{[k�ƼƷ�I�i&��@��Lv��I�o^�M0�!�t�Ri����P�'���$Y:����uI���|��_|?D #�(��o�U!A~��w���� ,
���OY;��}d���6�m�'�ba6���s'��	�x��gRh縓�d�>s2E'S}�Cd}�6qꖮW�S���������d=�@�9a�����VLC�c�L g�O�M0�y�	��g�bq�my�I�:���L2qP=��'����߈*�
�m?��E�~[�O����?=�'�'}�!�&��9��O_��SiXi2��� ,'�M�d� VM�i2�����&�gY'�l���B	}�*>G��-�����Oe�eo�����Y0��M�{i���@�k��9�	�w��6����0z��Y�9�Vd�>��d��3���&��<��6�Y<�+�|ˋ���7��)'̜��'QI<v��N[�;�=a��g������q=N0�a���8���L���~椟:I�<I=L���~���?r��ռ��>�oߛ�)�?�3=g��C�d��p,�ԙw�RO��q�������>@�^��Y0:��<z��OK� ���e���_�}��d�z�<]�5k���{����&x�=N��x��ş$�'U�Hz�������&��>�I���:�ǌ�Ra��w�!�'�y�Y�>w�z����a�ݺÓ�_�5�}���1���?����K������EӇ���&������Z<��"6�"Ω�B�+�m0�����;�@x�����w��ucҫn���X��&�����Q�ܩ5���2ٺ����G>v6�b���1
t8wzl+[S��� <��8oZ��Wǀ��� 8����a��0Vq�|�����(L[>I�N*J��03z�I�ܲ}l'��|�Ǭ����>L��}~:��n��<���=�m�N�޳��a�Ocu��0�%��!�;�
�I�3����Y�M�v�<@��/�ug��?���C?��G6���9�߷�ﺻ��}��ߙ=N��O�'��xw���0�d�����j��d�8�/p�0þҢ�8͇,Rz��@�'���|��~�5�}��:c���o���5�~���`t�~�+�'P��!�=d�}�4�8Χ��!�=d���CL���Xu&Y0���`'�';J�	ě'h�{l&<���u�{��_^�[Z/&y���sw_����#�:~������MK�Bq��PY�'Xu{���3�kI8¦���f�'{�Y6�C���M�a�5��a���{��~�_��P˗=!Ǹ���T���#���;a=Ł�J���`z��):Ì��_Xa�5����Rx�9z�8�Lù�8�I��y�z�h�9���.������W:^�s|���]������q�����|ɯ���|�sS��J�9�!�I�d��&�q!�vx�Y4�$��L$:�Oy���%F?�����(��{�;�����	���N���k!�ϱ*�����!�!���nN�k�)2���jb��<d}��$�7;d�8�d�C,�C�1�~�m��ݫ��;7�v.�~�G����{�䒤�=C���g{g�-���+&�i��� �0�y|J�u�<��d��SM!��<�ēl3~����sX�?�l�N��~��?C����<@�O�d�=� m':���'��g���Y&�����d4}�`m&�0���Rk��Rz��I�6ɦMkx����@�~���m]��B�U����o}�����M���-�e�zł�c�hf����]]��כ���̩�)M�ʛ�Ԯ�Hm��ݗz2k8h�k�M���h�	~�Oy��)�j|r�F�;��h>��� �3�qj��fh��׻F�����  ���p���>�����$���k2q�SvN$�,�򁴜d��!6������u����|������i4釳���Ï�}�+tY�E���7�{���}��ɖ tņ���L�f�m�Y3��q��'��u�~o�Z��w�z��NZy�b�������I�}����Y���h��me��V����H�����
��I��Y0�$<1a�2��8�3H|�,��0�ORd5�I�XO�w�8��`k��0��S��q�����E����;���V���l�:���ﶚa6�~��8ϙ4����$�bɓ=�P�I�5�,�g����d�,5�Cԝdι�a>dɮbN�$��'<�Q]J������3��:�����B���L�N�{��`q4c�>gzì�h3�L�����	�CY�
�'ɬ��0Z|ɴ�E���CԜd��o��UY�Ak�
��ߊ�;Wt��	�XOS��N��>`k�u���<~g�
�}����2xé9l�C�L3���Bz�(s�,���M�����������������~=�����ş{��t����q�'��q<I8�k|�Ǭ���I�|�}��L�x:�2x� xw���i�u����O����D���*�jR�L���u���Ƽ����|�}OB.�=dդ�h�u&�^b���CI���5��'S�sX�d�g�{���I�w��`m�@�<ĜCL�E�e�w����g��o��z�w�bTXM��,��I^�x���{i:��&���`l�����a�>�Y�'���bm���Q��� i�ﲝ�^/�18-_�x��~O�k��<d�,ϵ�q�i2�5���a�!�๲N��,Rz��� z§̘I��2�.�'Xq���d�?��	���#����un׮T{�u�����\��G�87ޜ��T�:*a|h^6/Sibӕu�2�����4we�\�]�ӷ25�c����X��H<׹N��"����yYqg>0`W�Z��[�R�"[���3ھ���$j&n�]�݆t�z�lO��!�c;�:o�{￞2O�T��8���	�yy̆�=E�ĝI�L5f��}�\Y'�9�i'5�@�%zɐ͇J��d�2a�/���m׺5���^���o����:��]�8�Rv}`m�z���:�T�2w���u5/p2m��@��ݲd��8ۆ���ņS��bL�f3�{��g\��y�����L3�w�Bh�<a�O�Ğ}�
e��]{�):��q*IY��p2nК;��al��5>�<`V��ۄ������ޞt������5�=�/����(e�I�N�l'��&|����y�Hu	�vx�Y8�&�߹��N��.�RM��o�͒a��������0m��L�����5��z۟�����|? �����4~��e���3l�a��f��d�瘝d�a�3�:Ρ5��L�qMw�<Iĝjxs�	�����l��1��y�t�������x��ƺ�|8�!������Ԟ:Cü�@�$��L0�s�f�4�3�ЛL�3�w!���qY&o�'Qd�3��2r���/C�ߊ�Ȓ2���^������/��l5�q0�=d<�pz�m�a���Xm�s��CIP��u�C�6Che�\��=I�]ĜE����{������=�y�\�ކ[�w���Zc�C���Ϳ$�!���C��L��}�d��,5��<a=M�I�<HgC,�E��,Y:��=���N�w��޻��=��{�1��tY&t�}̜�I��'�9lNy�VN�x�O;�Hu��h�����O�u'��3�L!�wa>L�jg�+:�>Mbœ�x�ɞ߾��k��|��w���>�4ɴXt1Hm'�3��)'��O��|��'Xx�!�hVe�}�pB���1�>d�7c u�2a�|�`��0ü��.7{�	�����h��[t��/�t�4�)p�^e������k�·�g����s��%3o�c�SY��0����v��ÔVD�VM��¶�q^�OH�K	�κ(���r�če��܆�5�����;�$;Ok� ��n�ų�,����| ��\%�~����?������P�-���'Qa�P>@�&��$�2l�pM?0�f3d����yAa4�S��u�Nyz��4��>����~�.��~���ٻ�|�������-$��oE�u����Y8ɶN�"��N03�1	���z�q<�'�>I�nwX=d�g���?_�u�k{�],��>~~ku��>�@�bN��L"���u�d;�
�$�E��a<S�I�R[d��2��'5�	�l�a�������K�o��cox�����3��O>�&�L!�t�3l�!��&�fP9���&Qg{�Hu�(w�\$�I��Y7i%x��?2xf���G�{�=tw���Jo�9R~}����ŝd����ć�O��d�B���q��|��2ɵHk��:�l�E��C�0�'3�sd�a��)5n���o�~X��0�˿O���N~��_�,�N�ɶ�<�d��!�z�(u���2u=�1�I�+4s��uI�Gl>d�,��
��&-�O������Mn�^���~��V�����d鲁��'�� z���Lrì�޽Ěa�Ci��(u���`��Y8���"���h|�$�<��'��^���^۞>�췯v ���� ~��a�7�'̟"��<a��6�m��,8�x���$�8�o4��u�I�,���Q���):�g^�y�>b�ǽ�:Xߜ#度�~�`3��/�CHa�,6{�@X�ܾ8Ba����m�L8�L�O�L��'&�יĝC�M���'�s��s�k�������5n}��{&�q�h�>�a6����qj�aw�}d<>��=a�i>� ,'�M�d��3Y6ͤ�g��a�L�w��hvM󇚳�f�G��b��+�Т����%���h[�H*I�V}.�}=������A�=�����
�sjh��]ɧ�κ��/����բ�%H�)�0t���5��=�<�Ռ��U��^��ZΥFr6@��!�ߓ�O^g)m���yb�z�D��Kᛧ@�R��-N̡wWe��ڶ�wuӬ��f.�D� ����װޅ7I�t:�3�S�����()c_�̑]b|Q-����h�x-�ٷ�~�k�׺���w3��Hp��:p�$�M��s�:8::w2��uC0>#��B-aQ=�1c�WL�ܖ�vQ]Y�w�zu��G)�M���w���"��A
LOV���Z�(З�4�T�-π�i$%>66��g��m�u�[�_L��B��Wh��
�R	·u�0ќ]d�!�J�;� �꘣߄ʬ��{�:����X� �d�e.�c`<����dX�-[���X�r�j���=@�n�j������T�Z��OZd2�:�u��a����$0�1dZ���t� "L���h����[�Ժ�.A=:�YC��f����.�.�yI��t��e�ȫumCFv��1k��gA�GJ@_Y]���̕�;x���cXֹr�N�#�^��%� �}��r�7��k)Pls�N��Wd5�bO�ud֮s�"�b�9`;=;�r��Ԝ�f��Wa[S"���MG{k.�u�Ck�T�`8�2��x�f-&�^�� ���"XU��p1���n�_#�a�w"]�rXJ�p�xMɩ��n����D��tI�͛9��(kN��&�Pҿ�M�)8ܔ2�.os��ݺ<�ukս���&N��t]�^X2�2d�՜��sZ�p�v����0g&s��s.�l��n�=�ށ���X���U-f���D�tP��tֽ��Ԝ���.�g��g-��-V�+jk��[Wy|�1�<��F\闆:t7��3ϕ�.��高��h[��,Ru��]ά�+1�v�`�\�M�nY�F��5�qe�k.n���N1��#��q�VX����d4���������d�w�+��Т����@�fnS7�$���%���D�gp�8)P��P���A�7�b��3�v1ZI�ʵ�%��l�9o^�=�B����[t��9gP,<M�7�n����<��s��2,J�st4d�39����dI%��|N@g�ڂ@e �ǑǢ��
�c���!"
���
h�����C��� ��u���_p�Ωm���Q�v��LU�KDT����T�2��ӵr��T�X��$���3%�+
l�������m����7JJ��^�$���A�]C/+u��f<����p+��FSH0��i�1T։z_��ﶌ�{�����(��c8�?g��7������un`�C,T,�]<qH���k@�Eɍ�)YP�N朌d���xކ1��i�5��*��,DTAUATQ�b�X*�Q
�E�
b�UUQ�"��TFDH+`�TOZ�c�*���V#��PTcUF*D�a0+R�T��)��b*� ,"�*�8����Ȣ�T**�UT�,�Qb*�
"���ł����,J�X�"1b�Q�1cm�����
��(1E1Q�F#�EV �
���DUQb��"$UQUQX�U""�	(�J�*&�TUE
�ATF2�QQF1b�A"(��el`��h�,�QAp�VV�"�5�
��0F���`�T1�UU�[lF҈�(�(a)����Yqn,"�@�4)�{�:��!�v���j�b2Wu'3Q	I�U�ש�R���a�Ci��ڴ�S�U�������kz{�Լ��G���}��|�y�H����E$���$�'��h3�䞲q���a4���l>̈́��;��~By��'����!�Xx�4�n�&Xu��~�����}ݞ[2��{��S�O�9r�z��0�0;�p)&�2k�'Ȥ���';lL���8��3�Hq���3��q��'{��OY2�����z� T_"��C���q���y�����{��i��7�Z�E�L���(|�,�3��3Hz�,��I�M�'Z�|�v`r�9�����o^�2`u*z��G��&Xy������s篏���ƽ߿=�d�3(tϘ��d�&�E��<HVq&8�<��=I�M^�XO�79d��'ٞbN���S��+'��G�_|!�����S9��Y���};�<M���~���~~.uOŵB~/�!�w��s���ht�ߔ>��%��ַ���Yޭ|��΍P�y�i���wWiǆ�6��_S��w/v��zm����{}�z9rg���}*�z<�n��2*�C�4����yh^��s��_�l��un�c�����$�h���� �.3�Y�Da��7y�4�3X�����:��X�ǳ���>�ޅ&!n���S;S�4����T�5��c�Ui��MU~����}�V��6%13�3ڲv�Y��&��#�m�J�|�}�̌mG�\��'-Mb�齏����MG������p�v��h��Z�V�l��2k����]��I�}�J>�Eje����w�]a���՚��x�D��Bx�G��� M���ji��������>�	y�K���|;�?|�y�L����Z}F�^O�=-��:}OB�]�M�ⷳ=�W8��6�=�nq�h9^SÅk��+q��o�Z��jhJ���s}�=މfo�y�S��F���c7u���<���X�s�C�-��[�O;r��m�cý��5�k��i���׃`9C����>S���7 ������Z����Lg�+��ϛ��~�KйK�:����]߮�����v�>��u�]��W���:򘥞p�l�7.>z��M��]�����5��ۺ�x�T;��e/T�]U���r�6h=��.�U�A���i�z�J���I���]�ʿ�B��Cr��1al�lu[��	�y�R��ڝ={�]�Os���#����}��9/ ����@�1k\�=s=»���_7�8z��/��`{	9��NS>=ʃ���CC #�xG&�-*A���Mm���0��t}�!]I�����F$��ϔ
��Kuc_Qꋯt����g�Q��iU�iI�Jwg���y�oW��W�V�mj�c���]��mͱ^����Qe�����.�`Y]*�.�5���_h{�"����yi�?����t��'{]_���B�=+��o&	���;��Ii�����Yu`Ҫy����~!A���C�������ϝ���;�S�\�����G���w��KS���ܮ�SW])]���\{�_vUn0��B�f��r�g7���f眪���ˍ�z3���;j�4�;�W&s�^�ig(�6:T���G�n߼��m�%?L2�:L����Ӿ�kL�L�6���,9G���w�����q�\����[��3�/�����Ε'D�޽���/5�O>T.[�eI��bH����b3���u�{�+֥buΚ/={햢�{��>N������r��S=���~Nӣ��c�{ǳ�r�t�,�{����|���c�&y1������6��tq�N{�o}O�f�ɝ�E���>�5����L{='ފ^�;ôNbS��l
5e� �_<��_R��z�����D�Fk�m��͑SSE�O�N�ݬ�T��,.�m�Yw�����Q�S:�:������Ec��jڊ��tD�ҥ�O46�#��n��Mt�;G���c,���eqH�dή�?}U����{+'�ߏ�gt�k�ld~O�_?��}�V��ĜΌ5|.���^+�96���Eo�tz	ǽ�䰞�`��Y�6�7�+8�t$�[���Uzϩ�מA���=~l��$p��8\n�F��{���''b��ɬ�m�
�:�kҮWǵzc�K�(woc���Ï.y{{��!�Ro�C��0=�w<F�/�~���x+�XNm���-��^���d����m�3D���Y�!��r���OY�	��A�A��ا�H��y}t�{�e���l��^_u�nESHu�W�������~���y�����w7���}�<u�8J�\�����_��T5,1�|����U��m�߃�gy�z�u�׾s1�eʞ���Q�!a�T~}U3�M��ٜ���0�"�����c�T��6%1,��Gig��5�;ݶ����Y�8n�TB{�7��U0桅�|��y�<�8y�Ɛ>�la��R��n]��7'ق�~:g��6{�:U�";e���U�ё���Co�B��o6��7�V��.j�[zU�3�SUj�V��TP��vg����������~�T}�H?|����`-�]sU����=ަ5��1�5�t���S������ٝ��s}S��Ԭk�aYD����G=�]���v��,��\�8���>ٶ�7�o��e[�X���o>ʢyi�y_]4�b�]��'���ά���� ~�=��&�d���{��(%�qg�������'gjn2��}m13͋�l�>��Ď��{ݞ����C�y�.:SK�����{��}��Z�n0����͜��1k��Nͬ��mV�L�<��-��gT{�ߏ��s��uP�6�������='���@�|��s��G{��n���PS/�����;<.�.��%�~.�/��^�L�w�yO��ow��N�;��������+�'ŃOzw��mo�zv/<�އ���T��?E9L=�����ބs�S�[��|=�si\��7�{q�ۦV�C�@Jؑ{�(�������[!�
_TT{��O�N�>�h��f�q�m�-�<șY�Oc���T�Qʛ�� Z86���ٕÙ���{z+�a�e>=����u�t�犯w7ՂǱ���� pH�9O��a�{�x��gyε���r仌§�tg:�K���e��{�#_߯_L�?�r�����y��~s$ͱ�/iܪ��y�ú}����̱Y�G��I�K6��X�/�v`�#zI~9�aS�4�ީѶ�!7p�'C��Zfz��G���tK��g/��D� ��s3�5r���t����;��F���pZ^�v���>;��g؏m�E(�w�N�~a�zBk���N��#C�T��_
�j��E\�y�yN���FgvAקս��.�{�bW�N�:�r|�W<G�ro֘C��K��Wr+fZc���?K��OG��]=��<5�UE��v�I*\[��mE�}��+Dz���u�[��o�ݨ�E<"�2ëK�[cѧ�K}R[[N���7�k�W'^S��^��w��=�2�|K�E:��(�u�̪�W���-���lR�t���Rua��J̇pP�Ȩ������"����;�F�0�9@KxW�ȴ�򼛆݇��w|�V�؅9�»��/r��;.��'D0�{�7�-`؇	 �P(��t#�9�?�W�W�|���H{���d��G����Ю�b���L���ېv�6eK�T�}%���ss�r�S#�������/�F�*6���*}[&�����޻��os�x��8�x�V7W�B���0�zk����3dȺ�����K~����}ҬNw2)��=�i窂W��z2�{��[5��^�<.WZ��ӹ7٭�*~�/$��^�ky;��e��3z{_f���$0�6y��:�����&�y��a��z�����?h���HP�	�:i_'z���O�ݷ����{���{�O���w�VA�ތ�:i£cL�[s3���Q�E��I�]'Q��zI�uտA���1;�.�,	 ��|*s��ަbȦ�:�&�߽'���{/�K�,7	����F��:C���}�K��n=}k�J
�&�ѡ�@��YXȆY"A~+N�lC.�ٻ뜤 ˧1��ʭ�z��[�� ���¬��C��[>O����G[� ����2��'F<Ա�u�˫5��Y�c��}�om�%d�`$��j ��VC��{�XS%%:Wf\*+<h��ot�9֣�ܦq�0yo{X-b�>���.�'s�k��,����=9Xڕ��3��)����ɸz3����C+._e�ƶo������Rw��S�a<������'W�{�J��k���gWJo��-�z��fT�"�2��x��O-���:�]�3U���ʺSOzs���	�)���t��N^޶��rv&6I/s�+��N���Gg�������T�bN{9���S�;���,X$~vW�E7w�yM�)ל|��}^�l>���@]��rI/�<���+']$�̑,��ݻ��V�ע����q��g@~3&#�y��L9\�ki���L���w��]�}�u�L@�W�+���=1�m<�hoۏv��pϬ�t����{eX��<,�A`��PL���~�׹9�G'y�9��7���ܼ�Sr��A�����gj8����{Ww�U��l]�����>i�{Of�����j-�#�|�!xB�ʳa�h3Kzr���V���k��K�y���[�H����co7�XDUƂ��w���B��ʣm���t�g��| 	M������ï}3��+�Guvݡc�T&��%��d��(p��R�f��1J9��[SfL���ү�$���<�B�v�8jXcJ�M�b[ard�md�X�B��9m�fħ�$�y
��K2��.�������½����L�eVIbY�x;���İgx%�~��\<�}�������ԗ!�Z�C({�<�H˙��ōb����-�����wˮ�Ȱl��=W�\������zPg���<��{Q�x\7���r�	��L-�E���~��~�"y�z�e��R�U'[{�Џ[J������y�Z%{���ڱ���3�{�^��޷������#�S��mo��w��pW�����~�e��ny�v�8w�͹�ړ�����v�{nez���p{������n_ε��6��
��E���өv!��'Sa!^s@�77�[��&�:P�u9��8�ۄͮ����t��1O�)J�9�h��0����Y��pG��/N�S�$��ںs�3\�K�߻~�z����p�W*͑t�������e�%�2W�_U}Ö��폷οW�m�+�~�WU��Nl�ْnM�.]e'���?!��ݺ�>���g��j�:U�Lΰ��|������o�X���ڀ�����e|Uﹸ{k�Yu�P3{������*�����Ņξ�\�{Nd:$��g���x�Ngg	�a�T��z,�SǊ��L0�z������|�g-����]���M�ͩ/���w���㵠OG��<wO�T�|�z��{�j���ɯi'Π�Ԏ�׽��xK��d����7*����=9���lY��u+�]=�1б�vξw�)�K8ʪL���l�P��r߯1�A\����v8x����P^�/i����벻��6;�w_�|*��
�#a�T9�����*�v��nW��0C��d��y�os[��o��w��q��{jV>�}��<QM�<�q�&�.|է�ՆƇ��n��+��8�� �M�s,���%J��wJ8qw	�r���WK�ɰ�K���R���gd �UL��`Y���q/���ӆh}rmc5`.��J���K��49�]tÓ{z�I�KM)�o)��!orh����H>��raXr��:�47�*�3��d`b�]b������M�;����I��lF�r��N�fL�Ŗ�Mz���S��dj[��Z��q=�g��n����֏R�nb��8���j���t�η�3.Ky����@~S�;kd�6���#A�>fՇ �y.�N]��y�/��*�Zb�EXv�[�:жuȪQ�y�V��;h�ۤʩX�CR�j��[�i�b�
�i桸��mX�j.���;3��b�j_=��Κ*�����)2�"�9פ�өe�-&�gwEptn�&�^`3s�]���m�[Kvd"j���/�^7�Z�t�.����|U�"�rZ�9�a�Ogt��t7c��4�%&��m�ټBK6�iD_�k�t���w��<kXT*�M�d�;���J���o��ѽ�r�\�M��<���ٴ�)�E�&����ۂ����@�fw+�i��c�*�Hn�z��c�		�ۿ����(�8���$3,�-h3��>-qUt�O� i�����*��՚n�ޯ�S8�\��Qֻx��W{� m2�ޔ^�Y]�Kg���j[sOq�3CV�)_}9��;��C���?u.A����z;�HW�f6�m{�R�WwVr�+O^W���͎�Z%�J�V+�{zC�cJ V(��r����W+�Z�dfŗ���{f�9-2V����+b�\뷬�ϙӐ���1r�Y�5	�//l+��j����ә�o�b�H��N9���勻mT5�p����b�&�&����2�ۤ-��vU;綶��d�D�2W$���T`�]x)�ĝd��'T-�|���Y4�d�.L0�]6�F\����a�1��T�C�� \���N;q���B�nWn��7m��q{�uh]R��m:K�hR�h&���l�U^�A;�k-���\.i'^�u{�FͼS 䑋 w���u��Z9�Gp��ơa�]��E���o�P{�퍯_ʑ�h"-c��Xls����R�b)���;�C���ݪm�me�����h:(^a	'v`[y��U{tݻ�[B-���sX�N���+h�Z��.���Mq$�&�DtU��Xj`� �:F�����X(Pw��8�+�J$"X���%�Z��i�#w�s$������^
o?"���jc +6�]Z�D�(�Z�X���Q\ҵ-j*",R,dKj��1��(��H�En.&,(����������0��(��a��Z
 �1LZ��,UfX�DKe#J�EB�E�F�cPQ*����DDEP`��+`QcX�(��R�R�QkEk
Ԋ�B�*�V��kUA��J�Q���R���[b��b" ���Z��l�j%ZR���m�����*�f�F�R�m��Y[J�h��Ym��ڠ�֊*�ahTcTFڍe�X���m�,QF1AIZ"�F�ģA��Q��ZQeeX�((���h�Z�Z�"�fҵj*��E������R��(�b����*Z�T���Qi[j�[�{����IA��#�>9Ҷ���mp͗Y����������̺�rnW&b�[wϳ=��4k�ꄛ��{)y_����lu���W�ӭ�޼�����J|7�y�W��zb�i�\N9�&���{��ݜ���N��žwS��>��cc�Ov���d��ϕx]���w;X'pu�jǟ����b�|��Q^�x��Z�^ϗ�x;�6ʾ�/�z[����U�g>U��3�b��ziά+�{��^S���U����Nw��O57��s��=��3�a��z���7� �7�x=n��t��us]/=� ׆ߵq�=��^����S��6���a��o�o� �!����}�#A�hpd.����{&	��=�3��>n�
����.u�V�;����6vU��rڅ�lzc���cث쓟��5KuOr�f+,Zr���m�kÕ C�;�l��\T<�w'fn�ب?G�ռ�֥�,ֶ���n/y�oZ��C��A���������Ns=�{g@e���	N۵c��{����b�.=���e��nnVU��.&+�!ǻR��[*l�C�y��Ͻx|}Z��ϔ\A��^s��|�ڕuժ�\��ǡ�fc��G�Uxz#�urή'��1)7*\�l}���y!kt|f��:R̋2��f�p�H�F.����za�}O��U���J��.��� �|�}���G��W�w�kw��<s,d�x��0��?q�^݃��/}���N�	\ެ�ss�>uyr;�*e��N�Zz���|�e�5�O��T����4��D�n3r���I�[�S�u�w
�V��=K2v����>��BS�%K�����o�ģ;�h�9p�م��u{��պ�{��E=�yZ��~�'hL:}^Ͻ�����T"�/5�����J��9	��~�<�{}��"~��^=][�uN�t~-����x�����2�Pھ�S�-��_��n/y����
�QG���� �(�_�yv�v�>���&t�I��i�{�z�Ne�t�o�=��yx⫛ʂ�bN�qs�3�M��s��9Ag��Z,aR��8|<'�],�J���^�N�'��7�Ǥں�7��W�����>�_�����p�YC\j^��Q�9�6��]�o���&����!8<ءe��	�g�.��'ZĨ�b3�^��"�z$��Q�ω͵j�t�[�����D�3i�%��-���������%ݼ+ߖ֋^�-��n�6i�T�53�<wR�V�]���Jׯ�I�ӣջﲣυ7�gV�پɣ����=.�ӝص6�/�mt���c��������`=ʃ��CB=�-s�k�X����.tZ1ok���]���E���:�Ē��r�4�A�����]�T�Zqp8�R��΄�y�w����b���˦�r*�C�Ɣ~�+]#{�\����ُ;��Z��p~��6`�~����C@vӅ1�euOvN��e^w��>U��)˰d���o��w�)�a��`G<���N�<�^<�g�x;���ȫ�_��.�2�$���}�jpq���Y�,��{�<�=�F�l�T�\�nyF����.`���7�R���ՙ��;���>z:�}�m�G�8:yNq�˷�+��𺝨ݴ��+u�h_#�ي�ҕ��{)I�1]FQ�s:�!wSך���6����vX�/M:�:� �jn̬�(1�[�r���ˈde�Ṟ٠ݶ��{9�t�澮mE�y+�Je���9��t`̘�3Vk8���&��\���}�US�'��y"e���y���%묰$�7���U�@�<9_vz�
��V� ���(N,{��ݚ�C�Wy��j�n���ײA�?K�;��=w����I��:���ʽ�'�����ٕ��yLW��Ŋ��S��;��ͱ��߾��8����is������Y�#�5�S����m)����o?�f��7Gu��L���"k�=K��笽���iI�꯭��-��l��ON��.����������}=��Ub��y��'u�qW���]LX[+냪�ZIR��Y72����;�N	oy�6��8_hCB �����k/z'[�ou���:+�#�-����򇧇��Ҽ=�왵���<$�ܹ��}��>�sL�����Ĺ�N���_gOK}��YS#��κxd[%h\��L��ޞ�{�xB����z]�yн�3�y�Վt���-挴�	=����G*�>ַ��M;�1�&�;��W�>�/���=w�l��**�֪�́���8ďZ��{��]��^>tn�]0G�#��o���86� ���?�n5kh,l�&�Q�^Ϋ�
aNm.�Bڲs/
��L��� �����Pu*XŻmvJټs�|>��1���E�o}�C��ʆ�%1�|��'�}�d��흙��V�]	�'��9*�|���7^�P�\Q�az+L�z�_������m����}S���o�{���1/�;��s��wEL���g�A��_m�gg�����>{�X�	��bX.=8���*u�/���ĭil�>.L��/���[���T�;���bW�N���el�j���6�ޙ���q;��|5"ym��e1c�vA��(z;V'�NU�5���Sn����Fzsz�,��zಳ�����b�z0�n�g�5�0��v�/Va^8������[��mk�����řZ=�}K�]�^&��r�H���et��9�k�d�LS9����L՛�������s�������9ޞ�����U���P�#סz���_v����|�'B�:sQ}�᳹q���nzCV��X+��kq�c+ށ�]I�\�8Wf��J����1\*aޫ�{e��p�ws��\�I;;}qT����kjD�V�#���9�#�����^��q�����0������Z��&�;��y��*�=Z�Ŧ=��Wu-�OfVc�l�o��]���  >���[y��~����l�.��kӟM��*{�WP����Ցp�靛���ox/��+���������{}'<�NP_��n9��{�٭��ӎ���/1ؔ���a������+��������S��YN��sݹ���;<C���6zX��ۏ>w�;��^��ꉉN�>���y���vꆇ"�4�ƜO�C��1ݬ�V8��̼���[�^�Ǻ��>}��/�/�&f��W���b�(҅��M@�
� ��Jz�K�z�V���vu�;Jc�>i3�b����)aL��9MT��CF��n��
����]���\>�1=��Ux�(V�#)B����&��\H���xGH�s1�2�{/����3��r�S����¾S*�yq�*Zm��FE�w
��vL��`��'��Z�|=)���vG���#�U�S��s�b`��tTsV�����G�o�lxz�U�#}v��^�4�熓�~R�ZsX��P9m�!ycu�|�Xʸm�+W�	�k:�<z�
���B����J����3��7]�� �s�Htgh�}{˝ּ�q�B9w�Q��g�_U}�T����{��P�<���=���	��Uy�������d=5�.�βү
o�CF��{�[�{g=`�k55(38l���zu�*�l1���x4�|�d=m`x����.��y��K�+��U�������u[�X�8-�K���8;5�ڠT��*��!���(�Syg���;2���U��� �7�J��ڄ��\d)�f]M����5{�OE\��-]�r�Y��vOv6�}����P���@r����Wj$�mC����[3*n>R��`�����y����n훵��J�c��4GR`إ�XP�ZL�,�N4�H]TV{Ӽ��$�����l�ʋ�j��K2ꎄ)u��о��/92�&����j�^��8��3���C���F��;=�IVjB횹ց��\+I6��j*�j�7;�k�m�`��0sOΤ�_���y�B��,e�]*�h��)��r[U�2W��|�V(��l{��u����O������q,w��N�?{�R��.���n��q[��`\VF��Ư?v��Ӿ�`�H�x-�V��|����z�W<_	��'}W���w�wՙ�J��s�Qk��3�}��5�ݏ�y·w+��i��#δ��DV�	.L�'i�4��.ɳ�+Y�s��wV�o]5�M�����MU�����~��VG�݅W����N��X.Wϊа���@�k��ʱ-�,���V�ս�c�&�_�m���N�V'|�Z�N�@_�CqV�v��0:���yʝ�u�l��n�������Ӡ�h�$�:�jݚ�9��W{hԖ+�D������)�_w�ww��y���6X&X���~K>�ՄOx�W�Z#�i���V2�p�9�y���e̓�f��p�yn�Y����)�W�fQ�9jW�^l�Q����خOv��e1٥P	_�=���t��N}�ǌ��@��ZDݏ�K�M���gD�
1���w�\O��y˗����M�a�ׂU[^����0`��r�a�$w�|6[�@��>��@ʬ�:�toZ/Dc�\u�Hb�v�~�p����1]:!z]�1/_T1`���j�A�`[F���:�Y��y���h�[J��i�� ��[v!G�x�V�%� �M(z��Φ�����Փ�i���&2�
��C�=�����o.��\|n�\ ��U�C����D��ޛ��2(���`��k�om�]��B�*������(��,�y A���1����B��u`C�:���H��
탍��O47:�����++7�ܤ�nf����:��S���L�5��0��aN��:]3ח�Ҵ��8�q5���u������|O9��%�(g:�_��[>�(2�?nO)�� ��o>�bf�����z(��y�#vֱ�;~^�<I0Tf�ϐܕsi�^����oU��J�B�z�R��S6�Yj�MN���x���f�w
4x�t�l��-G�GD���|p�C�ܹ}��N�<�zN�{;_z�J>"��&�^X8�yxH?W������lȬ��W���ɗ�{uG[��{����[9a
0�8E	`::P�On�e����!��S���n�N��]�^S�w�8���wڰ���4,<�h���W��J�L�_ٹ"@���h)w����?Z�>"�I�����!ņ����wj�8���Լ&�����H���{�����FN�g>�;țF��S�# �����^(�~*�e�Kw~��u�/f�yݾ��dQ���F�<�po�⏝��i=���;5,�����댩�\���􆓷���&m�jP�+"��^�i����c��7�J�6(���H�7��|L����ں2��w�>ɮ?a[����s��a�1E`^c����z��C�R[����r�����&L��P�b�]u
��-�e0�
+T̝�����>���Fc�0�d�m&�=�ᣙ�*�X��p�u��l�.��T����|)������r]y����lW�=oq}]���̬�6�&'��8)	<��]BY����By��V���k��<���;�p6�1�K���=�7���"�Ku��gC�[0DUёn����s�2Q��\�<�R�x��&y�9��~#���k�Fׯko��nu�'�%~U壊�z.��.�Q�]@F��U4:/Oy8+gOq�;���b^x���N�vc���rm����L:�|��Uif�
f�Q#���V��~��fX����M����ș��Vu�KfԷ�4��9C҅p'��=U��L�M)��0��0����e���#��]][-l�H��ȟ���M�ʳ��2!�@�$N����5㓱[3�jV5%�8D�V��ۦ�������S���ќ���|\WJ`��'a��A�qYU]�gs�"�[^	������׼7v��By�:h󕉲��/�xld��� �_0���qVgr��yk����{_D��c�/�����K��xJ����3��y/M�/�WH�=����3*�h���&e�~�O5�e�/.D1E^h��;��l�K���ܒR<�+�1��{kk�"�{�{v�;rubaK"���P@��`{�h7u��o6�_q[����B�0���/��DX:�N����ȹ����xF�g��F�����3v��� iǜ��y�}�ش��'	�|.�x�*b�rom���EG�8�M��l�w�C�t&9��<����ެ�Ҍ�C32k�8Y]v�����#n[�}��-ϡ����P�t{��Ci�q���v�/sٺg�1�.���(dr<���:���ϰ�|�(�Js���o7y9�iÙ �/�j�XT����;�> ���p*U��>ss�\��Èu(���%m��C��N�_5;��+���&�Өb��w�!�U���}Ý�6���/7|����j����C2�m�j�0S�U)��;�hV�-��9 u���pz�er�ZAX�L���]�n�[��}j�Z�(ѫ��.,c�k^Y�~D�Z2����T/kSڕ���qH+$f���ZyL�@�7����Ɨcm���8�A�E/�tsp����{�в� ��e*
����Fܹ�Vv���Ǯs���w�l	�,��\I�85��kO<��l�\8���73�5]|����=FVK�����8�h��1lo��&G̍Rkh��٬�T�e��$G�+��6��f�Xw1br�x;��k5�� c�iXX�p�\S7`;cXyo�q��\Gǀ���o��(05`������C�9��n��.�1�[3^��7�v��`����ە��.����K���l����E�ȣ����R�&=D<�"�~ڡ��m�Ptd�[�n�Y�/"��[S0��&�OOQ����TV^�Q��o�:�W����I�K[R=��6F8M�^On��,_t)A���.���s���sWm����Q�AG��)|�6��zn��+��f�V[����G�6�u�J�Cz�Ҷ���e�\4��h�5�S@ĤJ�\E��y����Jj¨��'K�.���=Z$Ux^d:��nf��(A��,Xٖ��ڴ���v�m7�]�|�(+:��w]�o�ϣ��<�qK��#O��B0�]jH[Lm-ӄF�s����F�b�Yq���.cE�^��,e�+����W_^r�b�Z�a,��pK�]V����
����V��b��n�޴�l�nn�6L���M��u�O�b��l�8>P��H�\�g`�X-�p���=�U�]	+5��u�o)N����]�M;[�1Ώ!jVP��34���V9)j�<���#\�G5p%w�26+Lw��ӷx$�]u���	N�9���:��\η:�le"Z�7��T�Ơ;�u�^LH�0�r��5�U��{}�,f��tp�*vR�Y���Cw[#�.�ip�	N]�]]W����m�UJ2��h���ڥE����e"*��V2ب؋Z[~�Ub�mUV��R�ҥ��kk*[T��ŃJX����iXQ-�KJT��+��J���K�V#Q�"��¶�Tb�JQ���bZ[eU�me�����TDjQ��f)�VVV�kF��)UjX�R���j�ZԵ�Z���iib�-�+hڢ��[Am�*�jԥ��EFUF���(Բխ�Z��PQAD��e1��Z�m(�jZ����kZ�Q+Uj6�Z(%-J�mAE����F��U(,Z�֥"��e2Դ�F)X,��-mj[)j�ѥT(ŬX7	p҈�U�R�QQ�D��F�DiYh*ţ[[F�D���b�Җ�e�*���մ�Q�/�����ń1�v=����'1��.楥�"��ڝLTT���V�����E�vrp;�E��dWU��;}��������������O���v���ыm3��M��s/H��]�������x������z�p��}�c]�\QR�I�bU��wY7q"�F0L ��5~�Z@���rp��H[�����hV��_��u���Yz|(��9�|,{������d�����#Ǻ��=zI����<�+}�W�!���	�.��%Z����g�o�JG����ƶnt)ogX��K%��x����G�0ץ���W+8�d=t�x��U�h74M��/��{���*�~�����e췊�N����Ţ��?��4����dZ�g�c��p=aݕ�����}N�^*����}o�ȹ�8';�/l�i��2�?m�>��E��ީ�}�z�9¸��P�P�_=�2�{-�﫦`P�굶}.�u���in�_1�]��^W3�x-���R6τX�?��z%W(���%a�.Jf<'տo<��Y���7�]�^�����(�C�7>�C���++����L��+�rr�]��T���W��2t�ϱ=>�^tVϠ��Ҫ��b���T^F�T&��lxg'���eޫ*���}B�_&8��:�f㳼�8F6Uv��.�-�o�@�먨�n��<�B�78n!a���E]��UP����[P"y��孑m-z�9Wյ4�����c��WϜi���Jc-��>f�ᲅ�s�3�WR��=\j� �����z�U��l����Բ��rS֯�xl��=ӯ�%�P:f�u�a��>Kĕ��c�$Zz9^�u��k^���r�ߞ[j�3��3ԅ�6X�Yn\�J��^�K�W+�S�2��]�I}�%-x6�(�a��;9���<��tcw�2��Q�&T�aD�3�6����og����u(٭0K�T�4�E���q?mf,%��[�3��*����׆�����8e;������+U|+K6+�Ea\���,�Tw�\������8�t�ROI�����]	Ơ}�^	��'^�����[�k=�/7¯�D�[^��<�'BK8&,h�ٲɗ(0a�:��Fkƕ�R��r�f�n69n+t<�-�r;��#�vޘ%��C�z�Cv�b��s�b��R3�%��x��f������ă^���z���Iþ��s�|0O���b�ՄA��3c���Kk�Z�9 5�|}2*�WD�U�:�&I��h����!M�.��&d�&�4}�GvcᅆAG6e0�$��﹢̾2e�L:���9���t���5��p��e�f�24P���ʈBCWS�P�Y�c�;2�h�V亖8�.ѕi��C{z������Ow��x���a��=�v*��c:^��`�mC}�Є��2N�Y���[IS�s�M~�����i�Whe�U�t��k #Ԩ\�9}��J���I��[�/?��ۼ������K�s�:���9��vz����^�2�6�ˇ�Н�{��vrͬ�=��oګ�����f1R�~����I�!�
�G��P+��}V�c}�s�ͺ��f
��ҙ��"���ϓ�����Z���K�~Y�����s���D��:�D�6�C�!2U����Xr�`;��ϥT!<�u,������rm�p)��>��x��ŀ�0��v/�����~�8`�^�?���9�!!��^��TZ�rʾv+�c�y�0���v�A���'ZZX�p5���8��[��fz߈�S�d���{�}cE��v_j�h��ȧ���GJOo�}N����|�5�}컹�{��v߼�srٙ�������ߜ�4,<��(������]j�b�=ݎi������x��h��A^��*�[pw��7�l�u*�u�b��E��>�gI�*t-ֶ5��b�.��|8�u�������\`�l �qݼ��w���n��A���.f��S ��,�:D�0dťs�b�ӱ�]��H�m��d�<���)��T��e��bUłoY#09a�U� �^Ѓ��yx���4�!�M�/ȃMZkw��lw��`��C6œ��ǡ=�}��,��A�A%�F,L1ޜ�C^4�؅��{4We�Vw9)_²7~��G%�:7�p�7b�Y�Gh��e�{c�Z�S��>��2<��.N(�\
5��\lr��3ꡞVÆ�X�Ֆ3��3�����ϥ7��J�3���.�v�Q��(I������l6�n��U���E�YC��mSț�|a\{�y����U+k��g�_oϼ|��4���,�������A�K�Lݫ�#UeƷ�O.�/�g�fx�D�M���-z�x��C�i�9߈�Vk~l߮p����0�\)��a���|xk�ٗ�����p�htS�-�s�z�O�B�hJ�h���{�k�QE�C����^�]Vx%��d+�r�xa������~��+����4�Je���<�[�}�B����nP�4�`ꔖ�y�yq6)����D| ܪ�D̸�yL��h�<�t��Z����2��&x[��`��N�]���з������·��P��cl7ծ��T��K&f�7�KϜƫ�>eȃf��f0b����]]�tJ�^�t�&�έ�P��76֔���e�vS���)����lU�1ʮFG�����ͯ�Jkv�aC�B�	=���iq}R���[>"��zoO1��$�]ϵ�ݤg���ںS�	�1�1 �}x��'`r�ܮ�l.V���Lj1/�W\(�ڶ���W�����S%Y�҄*��@��`��/m:'���pP�]�ozoz��z�8ڑd��^���˕W�4	.���zl`ylՉ@҇ �Z褡��:������ᘓ�	@�Y����ֻ����c������^���4GI������<�[�7���Fm��,�2��!E�˲���Ƣ��	�+0�:mӾ��c��f<�xX3����t�:* ½SP�-,��/o�0ȳ��V_�)b^�SGi��6����p�,��q$[f�+�D�5`��b�~Y����-����?\��Ǟ�漙�j���:��6_B��O�ʠY���-,JV�����J"�5��>=����Ow�ά^_vR�m?o�izk�}~A��Y�C�EP��S¡��n�-�F �"�U�ʻ��nN/��c��H4\a�jm+��
�δ��\�{]�ieY̱q������:����o���!tdY��3�me(��orCݩ�vl�5��9)�Fm[���th,<�r_0�f�:�T��dv�o�����Oywy�����7�T#B���j������7¯�W�X{5��C�MV�Ǐ�6��Ϥ|�Oy��<Fx*3��߮�ٱ�W��{�Z[+��3�����������i�+6[ъM��%����-`�z�ǅq��q'�1*�0ɻ^Oe�{{������s���t�&Q�L���4k��u<�:�ˉ�]Ѥ���G��~��r�l4�{B�oo�3�:��O}�t�DK>�#��-���4�n�'��v�h���I"ym��A�;���w� C:����ׇC����4ʩ����
��U����������k����$�9���d����P�!��g��l����n�*Ϝ�h�vj�Ƿ��Y}7��Á�g�nn8���B��<Ƶ�o�L���� 㭵[��:nܧ�{��V ��i���U)�j|_��>�*/ǥb��}�ρ�w�Nu�O��X��rM�U���lϚ�7L���i�T�V�n��V.PU~��'U�A~ўd��*�ض����v&�a�#�4�6β�k��H��k�[���ŰHш�;8)����o�M�&��:�����/�����C~K{2�Z�C�����^�N�9D��ҵQ=��5u���S�%�O�7�8�_��Lx��}ks$��<J��9�~�f`9����A��OEy٫������)(V��P��75�b�SVѴ�zɗ(0a�:���J����9��u2�����G��d՛�܄���r�s�r*�fU{����J#(w�a=�z E�~�H �~��ó��8�ۊ��Io[���\�{���a[v���
�=q��k�237�˼��_nN{�|r��C'��h�+�U���/Nz�~چ�!&۬2�^`����7��L["�Oz���9��^��Y��U]'��G>2�Z*��`c%0o�Lĝ,�/�[�t�㕓�ٌ�]������Io˭{d�7���U���
;Kǁ��3C��/!���d�n^6�p�+������LfeK���޳7��~âCM��+�N_�)�{�<�8q�Ⱥ�����\�C�S-�rxV�ȵ�a��:����Ӕ���93|/��(���m��O-: ����4�=6;9ԋ��*�7���/
>�Y.x:������[� �o9�Vd�w*)!EVݸ*��a:g��u�x:��[��+rmƶF�l�<�y�����+}����ؐ^���J[Ӫ(���y+@�]���t�E�xDg�b�F��g.Q�ܾ`�U��2sZ%{=[��os? ���w���lU/ݦ�`�>N�şL�c�"t�.�#�����y˾�1�o�K}�ӭ�ݿf(GRm:��i:�Ɨ,L<�$�����i(_���[x��#'�ӝvN�:o��j�?X�
���_8E	a�ԅS���g�T>G>�|-�9Kgz{]���8���\�׼댹w<�Ƭ�2�CC�L(���(;�c�k��I�sIU�=Ǉ�L����� }D��������w��./W�y����ա3��k׬����wH+{|�6q/%�۾4v�;�Wr4��O���f�iu<�i��wĸ�y���{���s��VE(�o[4ld�gqTQ�
�O�Q"���g�uvg��K�����X�lFrP�OB�썯	�L���_��м]����<I-�YJ��g93җ�K��f�4����� 
�<"�FY�7�8)Vc��
�7�v��4�S����R���sק��ce�Y�C����,��ѓ|�(?�'�>f��|�r��q��`l���ee�Q�ไgx�7l�N�.d��X�L��Fj���wfr�S+X�(pvΪZa�+�W.�*Ww���L�V���
F��ф�t�y�����y���P�<2q�����:�8��Uɺ�b��SLv��Y�?��}��{�W�wp`ם3���k-�3<֜��#ڬ�lޞϝ^8����M�8u�>����{^�[���T.o6ǫ�W�htS.[0�=y���2:�
���jmռ筴h� O��U�2��9#�2���A��&e����$3ں5I�#{�7û�t4��$K�������c�v%�6��ܯ!N�i֋�(=�^3���;���.;���iM`]]J�!ءZ	=�
���휩X�&>���R�/�7���Tw��u"t�3 ���p9/� Ȯ��z��4�k���+]�=U��I^;~����L4�2e{P����}&x��p�/	�xlD![6�#%���drVV��^�ժ>6U�|�8�͌�����K��x	U~C�d�}�S�G����C�>W�[u疷�βv>�/>й$A2�A�Z���}gj����I���w�UT�j�
�e^��s�{�-\�[4lu��q���
�(��J76
Zy�f�8\@ʆ�@͚�$����6�ش��UϟU�;u��x���#yp���6�gX%s��x�$jE�k�z��9��G�],�� ث�D�i�������u,�~�-JN��Ô�tҼ��+�K �(�a�ݗ&fc}RGĬ�-����`��u�o�`�ϫ�5y��r���P���<���YY�Q*�C|�0U�L�W�����h;V6�"�RR)VD�����O�u�����"�H��������LtylF�6��ӥ�>��z���ODh)�<�z<�e�9�Ř3��/��QϢ㤺�*������t���d=�gLG��=?���{�Aۿ��෦$�P�W���;g'K�u�!1x��҆Yi_�X}��}3����C�(�#�7L��T/���^�=;<p��i��w����d�\��з��;�t�f��x�����r�"|;1�����W�V�C3C�\gq{�L��իp�;�c2�u��?(R6τYP��㨓ͨbO���u�ܪ���^���(�l�^
���ߌ�]�B�
��nP���#ip7Kbȸ�������M�Q�7�K�
r�׃
7=B����L��1ښ
eW҉f�,!_-�����v��'��Wbf�?{o�]JY����Y�u�`�h{����g���٨3]:�0��8�R����P�~:��9�d�j����ws�n�Y���1�^7ײ��"��s_n>���@��꒙tU��s`,����k2�Z�W��.��3��\[]R�nڼ}Â#�TQ������ew:tf��t�TY4�J�! �\�,���j[�#J�x���؊���۬D�.u��
�4����V0N�%�X+�H��M�P�ڝ]�Q�#;�l�Y��%��c������mct���U����'���&=�{!�����|O`�n�Y&�!���h��p���w;���s3���h꜁i�ǐ(Àǅ�/4��8fV��#{0h`�p��}��P��R��f�IT;t:[� zhS��H��5�����L���z��b���Y`���O:��6&+	2P�ɝK�a[9�+�£����I��J�9AY���[Xwe,N�=taLY�6��e��5}�&&��<t�\���@��)�[ٝ�1����l��`%��e���wu�[����kr�˖��An�Վ619��a�)�o�V���r�J��`�b9�N�G6љf�r:G��є٭h=j�D\љ�ӏ���T�����-ʚ�[f�ƽ�8tn{)�ь�����?L�O�PJ�&�[�x�l>�ː��![�ݜiZl|�j��+4�9r�[�Mp��C�e4�y6���C������0�N���"޴Pq��;x�M���u[��4rS;�3pЭ�%�δ�1�x�2��J���ެ�<wi��N��S�c��f8me�K.���TfY=��=�ZH6��ح��56�Z�}PVSB��DpɇI���p龤��9����5�+�Uvn��n��v+w}yX�3�&�px�h!�<�|״��V�0�"�Jr���w[yS�����/�N�VTޜs[�tz�w�B�]�b�TW��H��ۏ;�,�)H�����H!�����n¯�<�w��n
�S��λ�t�[Zͤw@/L{[�.��m��1.�6dQ�gsG�U����<��8���y��5eeH���"h���j�C����M8�k�U�c�Tv��`���������� �s)|�\�m�O�@d@w��%QZR�}8���t�4��n�8t��2�;�Q��ΡV"��=u��[�pu�6􅫇8pr�h�1��W$������Æ��{A�p|ĩ];C���d�gi�����2�/� �Q���Y���Z����'������[T'IEn�,%.��Wָ;��ڴ^S���ok����-���B��J�����zt�_j���TZ��
��N�k�OW85��i�?gd��HZ&}���Ֆ��mB�?B�	4�*ɭT�68Ԓ65�ąjs��ioBG�q12�ժUT�i��1�Icˑ*o4jt�Kyұ;�̣����,6�J�R�:���5Uʱeu��Z�������ͽ�%�����j2��
^���Q�c�Վn]w�(��y'.:�t%�t��4j���=��$)4V�P݊ᴯgd�;Ӯ�t{kUu�9Q��U���F�,�_�-Ҩ4���ڥ�4�Qj�F5�ԵkWX�J��U��[[kiB�؈Ҋ[F�j����Z�ʖ�
TUZ �P���j*-�cYV�mV��TkQ0�KJZ��-�DEU(�j��Q�&
)m�h*�F��J*�K(�R�E[j�R�V6�V�m�*��QF�KA��)[j�YDm�-��bcf-�e[VѲ�[F��
V�m���Z�mR�"*����*�*-�Pim[F��F���*4)j��ƶ��Qj��)�X$c0Z[+ZZ����PF��U
�4e*5*-��RҖ���Z%�V��e
�Z�S�D�ڨ؍jUJ�h����X����[iV5+KZR��[h�F2��Z������m,� ~��D��E�ݯU�/wFF�Z锳94����:�9�����*{�l����:�(ww!���t���+�ys7<�o&99���~���K�4Q�,�qN凯3=���5��@�/en�[2�����-z�O�ݯ���f|�PЁjJ&Z��[\G�OJ��UĻ�װ�h>Ţ&�]����c��_���`� y]��<�)_���z�i����0�}_%q<A��։{�t=W���x�=����a{��4k^	����K��|_�ʊ�n�~�C��L�-��w����>���Ρe_�]�f+���}�Mҡ�vj�Ϻ�m���p���XG���K53���y<�������Xȸ�)�k�e�A��g��	��a�������q�Z�Ol�:�G%iLw�q_j[,��
&�C�ո��;+�d�o�9y+�3^>��ӧJ���V.�q�v.���C�n+��3�z�Ú�a�ޑ�����Ժp����s�<���ٟjz����h#��yZXa��/N]0o�mC^؄���>ꧫ���i����}N����پ.-�dRJ����4S���P�:�{'[��^~�BX�JY���5r�v�<G`�e$T��ժs��vn@���l7d��>�}*D ���f�#����I�M]/+���Z�\� ���b��vYJ�����O
��z�ls��ǧ�X�\y���ݯ�TExѡ�v�����<%k������[,�� �o���g����L�	/��׾%񺆰�X��P��R�C�D#�-wc{7nx�W6=��u�}=��*^��G���tw-`�j����9����~���g(v=�

ZE�� [(w�3�=4�OT,�S�n��+{0[�iw�^&��ϟ��,^(զBP��4�.҇r��"�`}�3z����^������w�ןo���������6\	kL^��P�J����}�&�t�؈j�~�/�f�Fwv��������D$Ĥ���3A:��-Ca�_�ՄyK�W/�gqݬ�}�[Pv����ߣ��~��t�"�p��(P���>�y̛	�Ь^qȝןU�%���z�\e�w<������zlg�{Z�_u(>���9�.�j�]]�l~Y��V�F���B�U�܉���K�a������J�d5n���ԳT��T�{D��܌�^�R-����O��7����Qs�6�r�JN$1ޘ!�AW]�/w_gA�-�eC�I����{m'�F��=f���}`�{3�M��X��)�>A�+��9|��l��V;�E[�v��ew���]����PS�X7�E
S%,��k�N�<�.���I��Vb�X9p�ٙ�V	t1N4�[�M��~֩l��XҲ����We��v(Ss��bk-qK�}��3�N���}n���e�E�_
A�=-�7�=���*�c��Ήo��6��I�_[���a�o��,T|6
E}�	�i�5�*�X�����B�S��?f:�<�Ϲ�U]5�tk��l� �ݕd��v����o�vK�L���_f;�;���ul.I����}O.�^S1e2̱��,�v<x����W����)Z����-�z�9��GJ�G�[���<��\��Cw�Z����ӟNw�3Ұ��ٿ�\�W�^�Ku����㻺B6<�<>�j���1��(��q+i觮��?;g�BAJk��N]ǑI����>�۸X=�¶�����7�AB�$o�WqV;iE��N<�Lk��vm옻���q����u9^���B�����
�,↙����� ��w7�u��|W�s��ڝiM`��Y��mR����>Z�9��X<ge��x'z��;k��v\>#���]���\��$UJ0z���X����(#A�s��#�ݡ�}��(�x�^��X�\^�m��^�Ό]h��(\�I�c�J�u��7A�Q�IXD;��S���"��%�l�y�nlٳ.���3�4w0�R��]8ɳz�Iؠ���˖���E�B�w�&�G�7��.��%Y��x	��^�Ao:M�o7����l���a?Y�*$��Xf�v܋�:ֽ/��U~BIw���zlu���Oz�Kb������RP4�o�ԑ������x-����P� 冔�dO)�d�-��^x^��{/����Y�y*jY���mN�∡H��Ͱ����M��G�������y�;�v�kу���t�QV:T��|W�eV�j�]t3^�UP��'��ܾ�r>��q����(�Vx`��C�WE�5���0���ϐþ3�e���Fl��	���#ɶƐ�������;&^�x����h����\��U�J�=	��=�H��s�	�V�z�~���8/�觃��,k�<��oW�`1�8GC��#nw�lj�س�ցÌ�5���¢^�PWP�Q`���K��u�^L-y0<�'��|_N|̼��}[��l�^���&�c޿����+����>0���il���r���V����j[�:���b��wK�;εu9#��퉜E=�[C�u���e �p�D6�ou��^���ͣy�Ф�t#����ʻ�Z���f�:����v�A�#3v���򛶮������vQ��Շ�ޕ�7���\�i��6�T��]�v�&ݯ��EM���(�η��_V$}J���b��:�5�[u�W%�+Q��+�}��+noӶ_�=z���e��(Шz���(a�R�s�[EW��X2�du�θ��$�k�E8�l����L�n��)�J��^P�V�b[c���RW���ǁ�$8�P~�|Y��Ȳ_+�^�,&{o�v�Ol��eއ#�j�f�w�o���Р$��%�_�i7S&�ڞ�=Cݒg��,e�wT���r_�ښ�'z�Fy�e������R�����Ii�c�R)��yy}�]��(�H7�5�?[9H�W����yO��KC����J/k����_*
�|���J��Ǭv����ڞ�p���NEG��u@�wPӢ�?p�-Gſ-
��}�fb�����}��,�ҋ?S3Bʹv�����|:T�aٻ �sh1�c�5���!#��ݛ�f�_���X�y���qguS�&_҃
u�,�׍+�ﯰc��a��VMM{:�Ԡ9`�[��c�{
C)�e�Z��Y��C��C�i�	7�c�J�~�kC/*;���\(^�ee$���coo���t���Q�#�����Gk���mgdxWj�a�x�>ޛ�#�rN��WP'�;�٢:L6�	ӫ�ǥ���3;$hp�G,��߃�Oƥ�؇��q0á�l���g/%������*k25�f�?m���O�^�k�1}_vW��,3~���9�P�acv<dZ�^P�Nf{'��ϽuQj|m������Z�9�̈́h��������T�����&�I9I���㛹�R����|��ͤi{��S�;�������U�t��k>#ԫ��ץt{9ч�e��������c�C�`��f/\�c�[;����׆�|o.��bT!�y1��Ͷy�ak!�� �gV�cN����q��ҕ�����b3�pz�p�~��E0���i��m@K�"_�;Y�E0�.:ǝ���}=�B�*s�.d�kw1\��m&J��b���Z<%���
V��7�#���a�2X�%s��"��^�����I�┓sP啤W@hrT�z��A0h'Zb�i�o�(�����;y��2Sli����v�|�99�(��c�b�Z�ꔮi��p4u����9���n�I���VG����9��6�s�A޽�ZE=	Os�#���<�C��gqQp2I�s2Z�m ڝnK�kō"�����]j|��]�������$�(Xibj�U�v�n���:��[�bF�נ\벪��k/7�s�BʹFc��jiūh9�����<��hܮ2s�� (���CP���En����q�|;�X��v_W[�,,7"��J��B����g��M�������ƻ���>Υ�B�{�p{|d��^�Ƭ�2�x�ז�Z����n^Y�����wB�w�(z�]Ta��v�C��Ł�.�sY󗓖	u��qx��d�L�u�����S�H���
���6�R�/m�637���Qs�6�r�JN#~�����R�k������`�ٯN�(�;�x!�F�l�h���gqTQ�P.��������y��"l�a>v��s$�AH�k�Cc�LW�(o�x+��>�H�r|��{���ň���e7]�
ܾ҄~�z�|@=Y�3����(`��	i�t����dr��cՏmY`�׾�bY֯����~^�V���1���Zڧ���^b�]�uWI$�c�{w��ՌL���`��@l_���[�ߌ��֝��;U���zM5��vA/�������oK��¬��m\S�Zn���7��:ǩ¯�E}s�>��4�Yj{=�X�X�W!��s�gB�C��^3��͠�׼�{�B��Wx֞��"�e���l��L]DM�`b��a.�%�W�܋.��\�W��9�ɩoZV��\�B�XTu��m�ړ�}��#5��u�>��������Ih�r��9#�6W�{H�:���=��#C߿)��ܢ���4�ꛛ��Wr�"��]��K,����tp~K�R��{]��DNY����z�u�Orx�+mt}2���a�Wr���J���,P��]��Z�q��D�;���2wo�GݳG��Q?J��8�σ��7�[��狼�0��a��A96�N���!�O�^,�P%�X.��]Y>�/Z�ǻ�g�X�.b�����(B��
�g��LP�W�ɼz���3B$/�>�̿����rE�n�kޛa��U^*>�40x��͹����{9Ni�7c��A�(m��M{gm���-�Ν��<�B�+U��c�;_*�8uV>�OU�u�n��j�U��������3�Dl��:Os�!�TTlX�e����*�nZ�`1U���S*��VZd'띷��3S\��ϟJ����P��>
�9�0���eq$FU�^(��U	�Ѿ��{�1�Mz$��[W��b����θ�^\7.����j�Z��*�\k�|�|b���g�v�)���O��gu!���Ϲ(���-U��<E�㇩>�{]��YQ���M��r��ػ��=�M��^�Sw)��G��	����Pw4{/��ެe�|5��|C�\�%�[MNn���Xư�)�ك;&X�z�4Y+�@��������ï��=����zub��߫q����V؄X�ݰp_��A�C�X�o���D���w懜X�ܽ$��߹�ٽ]shح��=u��d�t��A����;,>�n�GU�ֳϏIk���G��+uh�|+�L�OŬX'���0�R�y*`{jo��c�,�mo�OV?r��U5Ǥ��cW�|=��[>�ؾP�F���҆N���#B�׼9�b�ۮ�	o�~Kܙ��x4�L�2ߓ��.�D�v�Xt:��CMԘ:�YQ�yߥ����)��iqݕ��ơßM�l'�ڙjWR��隹D��/�K-��$�݀�o݆��h6�(\��/�gZȦ��D�O��y�\BWd�_U��i)��kY�^�gQ�Z���u��.,�(3�5�J���W��i��Xi�[��$���9ӭ��ػR��w��h��*%ꕥ��mu3`�<��1k:����W�Gf� �-u��q���u٣�����(hd�_1*DѲz��o'[���U,�I���Ԥ��
w�e�p]g�u�a�C�E푻%&u�>����53������A�y��mW	���ğdŦ>���n$��x��+�D!��uu�,���{6ؖ|:b���T���>eW5\�ӄS6 \�
����r���+7����M��Ӷ<�'��Y��A��k�O��!;�j�vj��&kR��Й�nN�����kq״��3~GU����ơew��0����Q>$�P�vjģ!֟���t�{gH�����U���t�Γ��x�CK�nk��^�`JmN�%���*q�2���{���s��שcܾ��V�b-�m,�ǒ�!�T!߻�q1�vW�F�q�3=y�r�=����1�⵲q�˖lB�{T�j���gO��P���>�"	�ޒnqg��{�_M��>�wU�ǝ4��ŋg=D����,��ݏ�+V�P��a�]�g<��#=x�%���N��0��o�[�[��W}�V�)?�
|e
�C̏p1CG���[�eُ2�:x��6��[�m�<7+WC���=fS�d�RvkF:�U�{��`q9����Աou]/o��� �M+yC�rيW���km@=;}{�_)CR�Ǻ����h�8��x���8�e�a���L�t�v(m��e�o�r
.��n��Bp}�t��{2��-����g�!
������c�n�[�D6Zn�Q̅�x*f���Y�(7��zrbe���8w8b�0p���|�{��0�b�f�d"K�Ҵmb�˛J�wbɝ�L��R�m8�!j9��Ih��&��\�g�Y����]�]�
ofr�5c���4ؼuz���yn(,�3 [���Y����|���7{�pKrK�Ԕ�J'i�
�o�պ�?h��֭��H6Ed��p��ę�L���C�������!r��Ey{t���A�muwn<�8GR=�,��|�-�E�S�j���� ��>�K�5��B��W����s`u�E��F�wN6۫���7Z͏�o<��d���E۶�u@ɏ:���b�Xtҥ��H�Rh�P:޼�s�;��/Z�Ӭ�8��򷤖l:�]�q�7�uՊoo}�v�B��LUϧr�m>�8H�"�jf��M���3P늆ܼ,L�eu����ռ[[�մ��
'�Yv!��|Xp4ws7��7ܷ6rk/(�s����7�� �Q[ �V�^,���кO�?�����8��&6 ޵��4�ӳmhIu���|;f�
%��63���`�i4��PV�LE�g`����wvVV!���LQ��_l���Qs���P�X�%�We�\���mN�J��wkj���o'J�}��ۋǙ1d7G�Sґ��X͕u�x��id+	��i}VJ��*s�8�<\�Vq�\{]9�]gm!Щ���.A-��Q[�Ǥ��&�ۇ������ȫ\��J�=,�WN�2���!}1�/���̱´�ّ�DV���	[���w��|zH&"�6l�W��1;�9(�B��P�}�[���eG�K�.�j���M��c��S�����,�&�\ݫ�i�"�C(dAض�+!&���`�f#6m�U�Y��D�f�I4!�j4��LJQ$�ƞȠA&1�u�����`����j���f=ܼ�5�ͧ�B {q��smy�ww����﨎�N2W��]�1�1T�ǖ� �{ ��ڮ�Rnn��܀S
��V���"�og67R\�q��M��~Թ`@ǒ��0�w=@�*�4��TNܱ�Z`;(䂬�*ƕ�޹��3ӻim-��>%姇	{P2��ۨ��6%h�cd���I=�3\6`�YS�Ln|1N�2å�d��H*Wk�o�j	�[�]Z�QC�ko]��$-�okh��+��RNŐu�Ʃ���@��n"��xNN��HZ��Šb#(l�J�&�i�-�,O���ԕ�KV�Qi�J5�2Һ' �!�C�L�;i�B�n�ۦ�J�{M��vn�7B+��O�A*3rU�+pٻ讍�W%l5��3��竲���,��B�*���F��)iml��T�Z�F��Ѩ�J%h�]��bԥ��mի-XZ�kK[AR�Z�ZQR�*��(�X��m-h����V�-�mD��QejҡV��5j�IKK[F�-R���YG	UV��R���Ul��(�������E,W�
�KiB�V-+F��*0�e���X�b�(-�
%l*�QK��`Â��T�ģ���e����b����ckB�[E�Ɨ.,mk�ap�6��b6TTm��V��1[+m�W�(��R4eR�m�1���m��h��Q�Z�1�"�-[V�B��U��b��
±Kl��
	YQ���V�Ʋ��Q*Um����.)F�im%�����*UKj�V�VT���m
�F�jV,�QѵŦ-�e����[h��0R��+F��Kآ%eJ�YKEF�"?G��/[��u����=�׺��$�f�]����'��nN�O�G�x�3=|��b�k��������7��;K��d��V'ܪv�tQ�c�]za{��2r��Q�W}��f� �C���߹����3�Tl!��X�<ic	��0�>x!�m#������o{w}x�o\5w-E�((|�i�WeQS�A�X{H��ٝ3ɔ��T�M3��T��Oū^���^��B�X�V����
���i�T�8�F����˾����3��OL[�`�xL�g��ŦhBk�Z��b��:e��:�6}xVֶ������z�xdu�s���s͸_��:lzK�V�C�H�,GJ�yl�
JN�k��{u�n�uq��K��,�!�������ƥ�ՒU�ܯ�К�ȶ�)�{��8]��R�"��KI��u�U�g� ;r!�W�H�冺U�P�K���ѯu ��Z�����X�VI�?6Y�1c��a>oL���<��f����7�m��&�Wc�q��9�jz���k�X���^�}�T>ଆE���y�l�*�`�J��Nߟ��:�矉~
l�E ���d�l�d��$č,����#hL�ez+K�A����a;c4��v*,A�+�w�5���o5tF]<�/�[>6�a��:�	�u��T�]�V�Ťq�F��6�#E�f�d�!8��h�+�W'S4d7YZ��n�铇Vs���ww���e���Y���6]��r˂+���*v8/�Z�Ivk�a�޲��E�{��o�`dv<Qسʋ��޿�j��O��b�Q�nrցSײۈl$���ժS����!���Vs��eâ��o�)����|8�S���
��j�y�{&�����B�MY�ۙ8?v����͇K������c���)¸�\.c0����=���'tS�^�qiW����Q�_����A�b�mYa.0�O�H��ʹK�̬.Ozq�W��"�jBu�z.	6��
48����;>�[�Qc�Uqf�]���x���9��^��Ǽ�[{�R؅�5�4�O	�(؋��=w*k�'N��adK��h4�(؆���x����<��	����=�|r�dS�e��0N5����6�o��*�@t��?c��؞M��~�:r�~ߨ��X��`c�g+�"��	����C�%�-�Mvϱzz^���6k�$�7_wlo����,D0���������f�g�x��d���;?X}e
H�5vg�7���֭���ݬo-�W�zԠ9�썸r}}�Ɋ噈�7�bh (��;�vb�U���/9������z��!^Jcʳ����^�L�W��{��J8��<��׵V-�OX�K���j��3�Xwîufݵ�rp��Y_1)n�|�r#�Q�ꋴ�Ѯ;^��(҆�RM{
�)���[i�Z_���Wrc��z����#X��X��w�����C&\4e�|��S*��K�Ȅ'��ۗ���K�&���U�9>�o�*S �`=#�U���.���'Q�}�xg�� ��6�ǝ�B�Jg9Yf���V`Ϲ�2�u�WEFk(����tՂ>]�gW��{mH��\=���)��ʸ�,�"�Zl��왲��0��S�y�3���<6磝��7�c����gu����β[u�M^I�~>�C��-�8Ω���4��d�1�n�w�f��������<�ŋ!���e�<�0g޸,X��`�-.��wn�W/mM����н�f��:�}Ь��|���x�cE\Vmi��w�����J���	xv��޾�~�I�:��V�f\W�k=W*���6��#,M����3���y�x�?r�Z޾�O�u��<�m3���2�3M��i�˵����ζ|�T�X&W���s7����Ks͎OK�YR��b���t��[��p]«Sᛝ��Q�Ow�:�/;)7�Ki ,w��<�W�f��urV�v��F��W&�4��I�p���k ���50�Gs����9�|�GA�w�Zk����(���!�^R�+P_ZL�Y�i�3��kk�3��_R~�5�郢�Ooa=7��r;�O������eEC��K��v:��.�^N��D������6��5~f��j�Z.�N��O5�ԃ*��]<u<����g�6WV[����c������O������3���q͈$���L�:S6v���2,ګ��r�oC�O�wŹ��i��/�f
.ԵcC���EC`@���p[�Mx�x�H�l�Kǩ���,U����	�X�2�[�3z��bN�P|8W$�ƨd�/�g]/&/���X�c�긳�T8�,��0���u�CN����;��k������X+�\����y�B���6�w
*Ħ&ubI��]~�2!�rxs�˚�O�҂��)u�4=�����]��x�U�u�ܽi��`�<|Q9�S֕eT�u,��ƣ�/%m����%b�-��V1�v�`���&Z~��T>�Ud�1��i6�z�Y�V�1Ή!���ڙ�9H�����X�X�l�ovoRʻ�ɷ*2�Z����p���v�l�Nk�%�c�+�Y�}�]g������S���7x����c�`9�ʅ
w} ��bJ��`��,�űA罍���
�{��{�H�������
��|�������`�}z̈́k�3��}w��+�(t�uKza��>�Ѽ�{���gD�^�I�����}�޺������GP��q]-"ڝdM<M�j�a�K#Y��������=�k��X%[�f%��p���,t�g}:d��o�+M]�l��}�T��Vukޗo��Eݼ2���PfR�Vmw���Kg���/�;]ҳU�4-���j�Gk�w^g�r��a�ؐ�a�O�b:)Sb�.:�󶕇����B�5�8��'/|��x�o��1s�����NW�N��箌Lؠ��0x�3#�S�c�¼f;����ʑ��ϭ�~�&_]�ެ���Q��Ԭ|����A:�L�x��.F�1�;%K���^v����e�'4Kt��(��[�b�0�BuJSHA����֖�){�>��fS~<���Ǿ����v�����n�R���$����Z��SH�&���S&�r{����](AY��`N�̕�Z�9���^���2U_��x��9�Xt4P��%;Yؘ�c�l��{8e�V�zsi�m���C5P�t�R�ZP�ۊε��q:��ʴ�ܡ:�Q1xޗ�h_C`�-����[(��JNF��ξ�]��-�%mҌ�rS]f����wY6�[5(C{]�C�s0fK�����70�������6����W�Eƈ�GJ��WP�aۑ����iܰ�J��Jئ�o$���ؖ��ղdܰ�{yXE����,����Β�|�pB�G�VW��څ��Нs�����������C�1ރ�C^4��biߕ���P����y�l�{�{X���u/NN���x���
�ҲIu����H�k�C|��C<���g�x6��?K�q�O;uQ�N�kqQc~Z|a�>�ce�
�҆G��u�҉U��,v�x���=th!��z9Ԕ�����h��=�@�	I��U�kz�N�fv�W���3��H��{������O1����<��	OaZ'����s��8ˇµ�o�S��x�u��_�\����X��dO}�V���=��Cz^|:���qO���!��0F�NM�/^u��R5@Y{w��<�^;z���z2��Sܪ�>��	U�.�X��RZ<�-��]�m�����Ftr\W��PR��u�2�y�b->V�R Ⱥ�����f�Q��}f������W��Ouwq��n��f�aB$h#���VWb���&U6��&��k�)wZ:��Ԥîg�Q�]����g:�g�[}:p�h���������,Tyg`=����,Mv��G$�q9�����R$-���2αſ�WI�S��Z�l���r��q��L�2���1���Dę��.�@{;:����̛u,��7�K�r�cS�e��'g�u�`=�����"�SW��d꺛DQ��]{<�m��*� ��
'�ѝv��qC�%�BS�lKĨ}=.b�㕔Q������}�.�Hok��;͔Af�a,�uT���ٹ"ر�KŚ�}]=�Yݛ�۩��b��w�	�fu���ᱟL�j R��0�$�G� ��3i�
���9�pY�c]�y�i�d�Ϝ��/%߁��u5Pσˆ��,����Q-(��H�>�r�Y����^5^g�?���A����Ԡ��DD�\�Ip�;_�\1k���=��/5��>��*���Xp�qgøU�0vL��`��2Hv��؉]ϪU�;�$\�����A��|�KE�A�B��Bҙ�q�f8`�Q~�і����Q��Fx�+s��y�vkB�f0
�\ZX�+LzUj�W~u����x�P������Uc��O5�:�����|��͟T�X���(
�걵L��r���K�˒ߒ��x1}KF�W{�hЂ˷�l��Z�{�u�OE���p���ñ�[9�b������w<��o{n�r�&x�X�2oS�=�AR����������ZU��剿?cTg�����է8l�C�A�Y]5�����	�[�:�5� HnC�������#W���K��v�������;�P�#�E�[Zrz�M�aq�+j�u���t}��yx��bd��z��U4�b_O���W��m��}c�}X�R���U����;�y��p�9�M'z��[�c�z�c3շ9O-�Exj��ӕ3���y}��oxP��h6)z,�q�t�g6W��T6{�̈́��S-J�R�b�}yvkt
��;�����Ȃ� 4cHeUGh0l��T;­�$Ͼk"�T>��XN;)�ʇk�����;{���|%3S_�Ht@�N��a.,�A�T���[��y��|eK�.u{��X���F��gKF�g:��ˡ]t<���T0K�+KY�E������䗉3�ڇp���g���x�Y[��Yg��+��ECb�*V�js�ޮ�[WU�Ԟ��_y���!�acO�����l��[�97�e�� m�CN����cV�n�cO���y��2�h;Q^6' Q{�ic�π�)�%D��s���4��1���i1K�%��]�7h۫�"�R���I�E<1����{k�p��%����ӻ�:�k��/��k�'�@�q�HqMm�y]�`�,v�&�}8� ܽ��ԨkP��+k�s�r�2̮>"�Ęf홖��:���˛��ʾp��g��&*�KN'O��<�Ȇ�k>�jk���A��|6�ƜIŻ���^q>���"֎��m
ݝ�Vm�ؕU���$tc6��|y�*ï_�^}A�&����J�{U��pV-�eC^|��v�`�]ˆ��,vlW�|��8�p3Ҵ�:X�X�k�K����#�̈́h�V��w�Ӹ�J�Wdy%������yU�%��{m�)Y��n��6;��&N����]`��=`h��Ž�b�:�,[�yɘG���P���Ԙ;����V�CK�'N�wӭ�u�������[D������gs��Ez���3�R�Vm}r�<s�t��P�02ٖ*_�g�Jݬ����^���wjyǐ�T.��<��m\."��(q�*5��o;ε��o��h�7�/+}����pq���r�|��r�L�eZ��G2_�R�K��M �(��A�Y��֌U�pT�.fKn}�+��i�;͚�֘�ػ$#���R��h
�lg��u�]�w姪K������3�k^mX����okp�X.�+���I-A��wX��nb�.�-�b�o_r�*X�[��v/<�s�ґ�u�r�a�,���:�������i�3s�������e�rS��gxύ�z��o�v�t��(ؚ�{�0�B�uJW�y�ewP�k[��w/�6�y���I��R��ua�P�+!��>���IXt�ސ^j�L�`�ڡҡ�A���wWO?>���$ ��1q�����Z�>��r�=�g���BEG���:�A�i�4'��ݜ�6ѽ�S:�4u����%-]^��f|v�C�UEϨ����\'��w.|z��'���[�_�N�A�2�i:�xv�3��<]�j^X�!u2>����A��Nӹ2�nLɽ�v��š6P�Vb�ׁ�xҷbiߕÃ���g6T4o�9.�^������{�L�=W��D�	�҉�XW%�����r���T<y�d�mo��!�W���BPf���j��>0����3U�Wx��-��{.�C�[����Z��o�$rd�����pR��\���W���[��k��g�2��Aa�U����N]��Vk�C,vtn�����y�zD&\�0�:���,�c�y��~�:�-�̢U:%ު��w�r�(���r��\t�O���27/JV�q�e��5���3.��.�=��[��ks
� I
�{�w}�M��j��b����q�p]2��K���uD�ܰ@R�W;�'$J�B��a�ۼ�3s(�u�G*�򏩼�M���t7�����քff��,��N����LVͬ6淎��:ziZ��Nlrg7Ǻ f �X���WwufLM����#�.����n"#��Z_Wh�3�Լ^��u5�Q��{�Ў�9�_`"��Z�_ћj�,4�>Iu�f�Z�#{k�`�Ǯ'Ca���0�t�.7�h
�P��T
��v�:,���]� m�V�F'�Xi�GV��7���7��s�`1T�:�K����@���[�T���%�� �v�꧷sB�~��QӤN��u/ H�$�_2YW�`�t��;ή�p֮y�7���so��َ��
��`�ә�xJ�ͼJ�5o&��/��p�W"�2.�i�mwKϤJ���!��Xr�
���ݐT�ɥT�y�%��:��['0eq�[��ܭ�{
j߱q)�"���03[P'�7��l}��rouG`��2hPӘ��MsTa��p��n�e���P�y���j�ϱ����g:�����-,��PՔ���s��6��;��߃�86sF'��<Q��u҄}��&)�\���f��RjX}�5�������Ig�v�:醱�f\(Z��{E��-Q�r��Y�-�	n���N�ct�@�n��K��ڗI���h7o�ڎ��+�qG�%�q�A��Y;��1�:- ���ܭ��8�P�β�����p=����m��c�CIp�sOS����a��e���P�B[��������6�)�����	���귶�3�g�] �jܷ�W]��h��e:���Vj[#����z1X�v�Mb�J5�<G�l��U�+Xͺ� �)�T`]����'Q|��Ð\����V)LO�������p��h�]���]ֱ�x9մn�>�����G{ݚ�Lgm��H0����.!3f]�WS�J���`X��7�B����Vc.��:�i�1e��M̡�c�{��#/o'L�yI�Z���D^���^!�5�Ὣ`Z�Y�p�v�rXx,�̥#��/�en1.7B���,�-9��,��<��ܷ��p�F�����d��gj�V��5�%�׺�A���w��T�Y#�Ò����X� 9b�*SσT�SM֐��U�h;�⌑Z�
}wI�_�4U�]n�ѽ�oMLȚ-*Z�����;�t-��g-�tX4�X�*2]Q��Y�.R5�A4�cQ=�Ud�Xj�PhVfE�v�날�T\�.�.s�7:�CiX�����UH*�Q�+
���@�+PR������PU*Q��m���U��,-i�\YqQ����m+
 ���[J*�-�JԩmDYY-�b2�Q���V��,�b��JT�R�[jVDcZ����KcU��*���"�%�6��A@�kicYE*Z���l�YZ�mb1Tš�Tb���[`�X--R1�[eaV
(��DR,mb��"1E�E�Ej�F���QRT��J��
%�R���UF2(1��Ŕ�b�F"�X�8aQm�e1b�0P��*+VTDJ�، �����V�@VҊ�8j**�����TX��1`�QX�V$�b�m�1*UX(�U�Q�1UY"*���V,XĔaQKaZ�mU��iX����+�`H)AFi.��i��5j��7xass;V �N�\���v��9��Q囗��Ϸ륖��~��9�c�	�]��ɝI���#)��3#O��̓%��{A{�o"����֨�GzT��m��������:D��и�m~������i�k��8OS��Z���C}4�7����?\�gv�1�)sgNy��2�����b�Ӂ�~V+j��Wo �<�K:}@�ݏ�_2F�+�iL�.T#L�S���\��O�!��t7?+��,^��3,^�/zd]~~��:�L��D��0�oM<S�t�6"��O}w*k�:t��"'̭�S�F^ztϟ�$�h8ußW��ה�����b����s!u�e�U���]��z��u��q�=�
]����7��?h"�R���%�_��l�W2�{�u��I���P��+8Z�^���'�ؠ�w��:��m�Y�D�>�&fa]a��nE1{�t�Й�*�n�%ړ�a�~�7K��^���oh���\�iCa��&�<C;KT�f�'�m�ꅖ�绺v^��}�5��y04�]x��]�����:%��p0�T�U��؜:�sY�/l��	�b�@}�t��W�o�Ė�2���E���QB�Ob|=woe�Չ��I���{��k1B��E'�n��S�K�O^��K
�*�n�U���"��t)b�]:+������J�6�Z�gg��z@Yw%H�u)\K���j;�E-65�l��c>w�)�K�4a�*��R��7p����c��ϓ��T�7ԕ��袞9�7w
��s�e�X2��đq��(�s�t׹�[)��J���L��~BcR��++xo��]2Y�R�C���>�
�b�q�@h���o�ב���.J����#�m��X������n]�G����_��A���w����*�^�՞y
��y��f���փ��!�kT���kԫd����o=pth���T�����:�;7�y]gkѲ�xV
�YI����X�\s	
J����f6)�h�0r��m2M׫�i{�t��}<7��W��m�Ϭv|��Rey�m9M��þƺ��������z��w�]��r٘l�F�,�&L�+�����i���?7�<6P���J���yq����7L�	^��;��b��A\^��c��j륐���Q,��*��+��6G5r�w��$�}��N5�W��3݄U[rśSWC�P��_��;'���;�7|��K"5t��j��r=+�4���zO��)���D��C�/o���D����nf�5tz�Z�sH�e�;�Ζ����;�yǂ�Q�w�dcf.��a��ܱ]5rg�,ol"&���-u���2�����:�M���]H2���v��u�����ض盬ֺ|��K�Ԅ�B�m�x���.3�P�rUR����W��|d�ؚ���=�V�C~���y}��T�4�^36���t<���|�KX'�-Hu?3T�����nI,��~5�|��!�XYϺ�=�ze�ޛ��T�!�]CU������Qk�����
�E4�ؾ���Ư6�7�u[Y�*�P��Sh2��9������=�r��wٝ� z��	��'[+P����\�+/o"Bk�mS ޘ�ˤ ���k7�ן9�|�wfm:{mY.�B����W�����=mX�Wo�_�/"7�b�����"���Se=����}Zɛ����g!W��#
;%}�^�J4�!���S�]x�z����3�]���F���4/|֐ƺ�ଛl�X��ֶ�h�l"�K/���nڻ93��G���Y����/N}��������Kk��o�~�}����qUx[�΄���wrۏE���۫!=ޡ,0����3���t����FW��ot{}%�m�]/D���i�LN�u*Эq3ÍI�扐�-�f�뢮�yk��;�6�YV���wt�#ɍ�b�7�Wr�����'�-7]ϗL0��T9)��Й;:��i��v�2JZ��������W��(��bX/w����i��o!4��ۛ���=4��0:f��4�Ab�]�W�X�a��֬�Fܨ�7�98d�fz��V�7��y�鑆޾���ܵ�B�����m\	#��q��;iJt��P���'3�^zͳ~��(aϫ��qJ�W��`\�9Ap5�u������#��{��e*��5�i�=��7*xW�ͨ�\Χ�P`�u�{�US�J�zz�����LP׺§�z��3�����O�QO=��?��]�ʺ%�ӵ��cN��.��=���6��+�E	y=��y����@��q�`N��.��VC�w�b�y��ώIw�m���	5ޞ�X�ţ�㓧9-]z���Z9ء� E�7�ʆ�u-B�K�s��2]痯��}�G|�Q��ǖ��+ڷ⽨�QCDK�(JZ��i���"�qc�$Z��Z�*�����u��>�����yB񰋮��?���)�����:x� �G��ʝ.痢�wu����Brp���ڑ��shV���Q�߫j��^ӥNQv�����^7]}�j���2	um|{C����B7'���]���;#�5�F�����[�˕��^=���wT�x�Oz�����!Z����Y��ȡ�7��h���8�e����|�����y�HO�d����	`���f�iX�(�~5D?,�K-t����;��*4�]o��7�Ǝ�� �����6�9҉1A{�/���򤯠�i�%�]�ܾ����������!|��5x���"�7�e�O�0`�d��3S��������DmU���lZ�m�*l��
^Ս{�Z*O*�[>�P��x�x��c�<�%����^�o�ޞ<KmW^ߟ-h�7�zR�Gk�y�����]�~�P��_��;��D�?s������rӟN�4��M���u^7[W��� ��pם��l�zwp��盤�ÞZ���Ô��D�hg����1yi�¿+�e����#����b:G5�w:w�m�'Q#��̫{J/E�˩��Btڳ�tAn��B�>F'��
�߼�F���ex%c��\Jivm<m�+~RJE���<�w*��ӥn8�T��½�q-���"�+����@s���ݳ�+��p���j��vy���ػ>�V��J�N��7N槲��Uӑ��.�u�a�Zך7���T��y����>�����|�
�|������S&k��\�+���F�'U�v�4�2ĖP����=�m�r��AN���7�$��P���âƍ�[8%y����+f����c��K�pn�����],X��-z�.j��9�,�r�ʥ{^ғZ�C�k�q�/On<�ÁŦ�@�/��*��@�l"~g�V$���3yٹ"�'Ӡ�>�ڝސ����x�N̳^�^��(��&hT�/��e�V%J��t�A��TOS޻�+���yf�S{�5���L�u�����jj��,ݳ�"ǐ�̲
�:yӉX��ذ^U�n��wY7�eX��	�P�6#�r���T���ԶJ]n�=���{���hX�%�5m�B��ư������|��XP�`��"sؕ�wϧ��eK��C��զ�U݆WJ���Bj��K��mX��R/�ك9�29��=?�l��f�3ɝI�����d���A�~Ō�U��4%�L
�Ӣ�z�y&�JV���+���kDrƙ�u;^��5��� ���eٹ��G?�����";��g�2��/x1'�h7^�.x=��z�����=��S+)?K	諧��tbu��b��nK�u���M-�ۼok�ƲIt�M��u`�9��J�H{�y�C!�.Wҷ0m.�z��n�ңo75����d;��K�����
��r1
tou'�!g�K"�ԡ���M}�^�?)�ɂ�"JWQ���,��Rۇ���'Fr�ܒ�Ԟܽд�r�8�I��eil�_S3����qy���54��[ROd;�w<���q:WjE�-՛�g
�D��1'˖�ʛ���)�h5��ڤ�������S�g>�J^�c��0���-��
�c��8+e�(4xOW��g'�����wG&��{f���>�"Y۪,!K�0~��ʱ�N�&s]z+бD����3�{�����9��EOog��*[5<]�S���	֒l%���A� ��Ey�zl��;3��c�e�:����i	=,e��ة���l��C_@�*�L�ϴ*��-v6��Ϸ8{fS�"���Z����,����^36���3��LV0<��XP�7cv^��y�Ǳ%kƵO��9��̓�MBş<�����>2�����!��c�nߔ���s���YEP��t�����'J�(</�ܥ�8�2�]�e3�rJR�^�W���vf�zá�<, ��]sץjt���b�V3o"7�-��mE��3*UP�k���0�$��h|���yn霃�&n�X�Z��ht�˥\����8���;S԰߱����˼oԩz�7���,:S�7�ٚ\�6��]�*�(���5=��"�o���ɦF(���i�$k�|��x�'�r1��R���C�+{����f.'3+�3ғ���HuYo9.�-�o`���:�c{���j�-xxR�m�r�mSV1�[ך}�V�7Y�Ǔ�����ڶ����[����X�׏�e���Ez��6<�q[Ǘ:����f���2O.�3���>�"�c�`��d�`��v�Q൯�h\�ګw�Ĺ�}'RR.��_��wשv�X:��y�����	>x��c��N�׶V��T	�Y�)��r���[z���h�j�q��K���Ͻt��m3��)XD6ݲkU�7�ψ��Q}�\dOW��O��r�����Rvi�n�":����X��<ly�Jε��7�yu6�UOf�ڝ[�էdY�6�ף�m���iX}[WG���C��
���J�Sϱ�$��\p2�t�r\��Μ~��0��z|��Ghc����Pc���᧥���F)@Gr��j�1��X���hJ�����v�l�x��sy�W�{��oal�v��>P����휥g�wOnX��~�75��/|a��8T��s���=F�OW��2��NǁvkH���)=�Xl
\�iZox(y���0�^��� �����	�\^�Z-`=#<��]oo]5�Ɲ��t���ms�<v�V�1�/w�������<)�Aui����/:���;�'b�څ�g����g�O6�#�k}O�y7�k��pD��#�B�P�{|�|�q�2���KP���c�.,���U����I��
he��/M�ylՀ��%���B]֮�WL��ۑ�ڸ��[X�L{�v�y�F淂�ިL��}�qxұ'��[A�1c�XO�<|g����j���=�Wۼ���f၉V�N�h[r�J�b���2����N��������k}°���%���_���'��ƍ�Og*)���p.h��t�`QvX�&6
G�s7{�,��K1��%�hvU�q�+"�7�e�Z|a�9�2�]��I}�{{nh�=��N@O.���w�>|��w=��v��g)�<m�'*��C�*�1�1��,�2j�/A�0ٺ��boZ��ozV��{�_V��Pj���q�#����E,Y�n��n�R�[�zǲ���Y�.g��5�s�#'��ٽ.V�b��b~>�ks��Cֺg5"�i�%����_����zP�(|d�U��N��D�����9��W%w��� ��|JqOar/�&wyX��&��R��s\�����
H%������NJ}p�Ut�����Ci�S�)���p���d���x5���[ۭ�^>�# u8�:y���0�=xτL����7�>ZX5�¶����4R�m"��\^����w/ԥV�(��ꌧ����2�y�bН6��E����7�Y�:����-N{�/�
ug�}U��vʉ����[�O��*79�諹S^s���\w2��nt���_o��:x�b�h5�O��3�L�0�S�ˇ�gӍa���үk؜�^=&{�;�BA�pf	꼜���F�}b 쾃@�҅b[9Y>%�B���vv�����t�Lg��R�l�zJ�B!
��m��D�>�fX��->���zWvOGs�}�}ͨ"س&{�U_��&gZ���62e�Q�,$����$x>��ۿ����0�(��9�����3�K%׈��~rΪB��%��[^Y���M���}�or��C~�-U|*R4s�7�O;{	Ȅ,���0�Ô�QW���٦���v��ˑ�[��Fa���^L��>7���ŝ¬�Ή�,����{D�WK�v!�[�xٍ:���|�$�iBmd�]�m"���y#��wB��at.��wBmYt>U������+��BJ��	{[׎��»Y�g����m����N��u\|�]u�Չ�GRʱ�{���B��1�9��h��΍iÓ�؎ ��>ܨ5�s���6d4�Vp�_r�p��d[@l�M.�QlA)��^�	��xn��ĥ,�!,�;y�D���#3����9�o��n���r�Ǫ���z�Ֆ���[�b��Ǎ^�v鬕�K!�{�뭈 �[0�m�[��˼]�"YDiܝ7�W�\� �c����cC�sp1 ΋��:��� u��IuM�Ւ΂�	�n�G��ͥNnQ�ֆ�B���ډؕ�wl�b#� ����:���J��1d�����,��f�U�(�'M�:��H���ZEv�,:��Kʛժ�{QC����V�1�*�	����P-j�yt�Ļ�!YZ�4�B�ݵ�f*��罅Z������yo$Ţ�� �J
zs��Rj�X�z�.��[�15h��'�2�f�
���;5}����*T�WL��$'���Eb�O2>�n��y�,kJR�79n�N�D��ʺk2��E'�`EBz�
 @��2|-�XyΊ�n.j�f�a���*�H�Ԯ�$�PIu���+���zΊ��3.�=��[=NT3����e\#��u6�i��|�K��L��{�Ш`]��_s�
Ϭi���r)�D*Z��ǒI�ȱt��.���oɾ��]
�Z���9�oqh-֋�4mS�nb����f���1ň� ¾{�2<��U�r��_4��Ǌ�*��G���u��4.*���w�7.��ѣ�>2�A"���K4�=�&F�Ɣә�F�T�1�]�.�3�Q�ʕ���GtR8�$�z�V ]0�L䊶�^C,u(��Lt�!�.�ٝ��˟M�đ)[G�����諔^`�FKA� �˸��C��:��K��Ơ�pb��Vc=����S�4q��=��ѴZAE{Y���@��}L�m���%'ǉ��u
E��9��$��\�u�E��3S(AAͳgS[5ؖV$��@%Y��36��ά:�R�+�&$^���']w�.} ����V�̺a�-���\C�˴�3w��2�Ы߻O�zʫ�2V!g{這��Z�.<.��԰�*���
X��i��e?�����U�E<�YL�U�O�V@����,�w�
!�𝷍Q���K\܂$�5�5;YD+GqӢ����ުmj+f��8N�I�]�����n��[��aFY)�����a�ҽ�2��g'�ְ��]B˨N[���T�c&�Sk*,�Q�"*0X�UkE�#+kQ��,�+��b�V�TU""V�+QV�TTR�b���*���F(�T�PDQT��TQ��
��,Q++T�2�GP��%�AQ�b*�*�"��*TQ�KJ�m��@D%j��(��*$R�V6�Q�H��H�`�B�
�X�KX(Ȋ�d*��F*���b�EF
Aeh�PUX"	K"�TFҤkjh��b�)*6�,Z�X�X����b���U�AdP�
5+���b�VVUEQd�iAH����(�[eB���DETQEQE(��+)E���B���J�[R�Um+*,+�UaR��m�V1�UDR���1�J��"���a��-H�%[km�P��!P��VDT��J��QEF
6�"�[jV
�ʅQ�m`�"��6���V�n�#�Rm�"+i+�Z�VC'��9�}��w�I��C��w��a:��E��}���hJ�8X������,மB���w��Գ�;k�j=1���]q�m�M6 ��Z�w�G��}�<[�l�[��D�Q�{����.౼�|�G%�<���a�7��-���yF�_�z���U+Y#<r�βU[u�K�1Q�g{�Lŏ��o����W��b�ǝce�Tsӯy{�<��ΔN�=tV���x���jzQ�[o�rg�'�����y����=����b`�����P�#�����h��*8xqrWoo^@��:��f�
�y*`{jlW�Kez�3%t��9_�����fݗ�1���~�L��iWz��FV���f��+����O+n�hY�._����}/��\�������y�/M>����>�N��e��(a��`�-� \tt�g��S���p��fu:]'��=y7	��:��@�5<u�W˨0I_���N�&F�u~��nN��y�[�Pl�l��,=��uƤ/���5�i:d�K�λt:�F�ݏ�?[|���lyoΦ��kϣ�R��c-c�x��pќB�D�qo#�
c�8��]pVV�>�+��ݘ�7�
��I`̸����e5G�N�BEse1C�J2�S�8�]��
��;���raz�[�i0�eI����2bz*�w2^2]ѭ:��K���2>�N�Z`��u
���`���b����'|�X�j>�6W v,�2X�V�u'P�J.�}��\�=^c��(�#���Du[_��E�	C��ST�~�=�<�=�/LU=���zR�c�D^۞\ya�{��2:�-J�kME�����L��'r�R��XCzI�v�oSo[�	�7����0z隱�j���a>�>+�B��c����q���'/_XFBe;G�t�s�7�㛵�}}�.P� s_�>a:���LU���o�t����Q�k+xLw�߽-j=��!���Z�7h�%7�~J2���P�r����k0��c]�s�0��_{<�f?NY�=\+�[��y͈z�vVŲ
G~3���W�sïJ4f!��[�]��{X����|�����L��=n�����`}ZD9���x+>���ٳ�?V]5���A8�-�g�����f���¦���x;�x%[^�c�P����	8�ޙ�ά{=-�R;�ܤ��//ѧ��s�[��o�pS���m{�E���s���dC��^�Nw<k+_�9-y�y���Y�o����)�++ԝ�k����u
����9q9svy�J�h���a� y-Z�Df�3���0�cEή�����5���Ա*E+����s{�f>a���e4q�9��3�1��d�k�G���4�����/#�s��Jz�lCas�XyMz��\�V?t��V��������:*Z,5����GE6�e�,gmvڒ���f=~4=>��W��L�&a�M��+�[�l۹j&P<�N���/�k��N�M}..�<���U�Fh=Bc��}\�+g:�7�o�*�WX��s9ޡ�����y��5�B�g��Y�0�gE+<[�r����F���ؼ2Ѕ��W�:M�5�;9��M��^�B@�|�ii`	�8�s�x�ñy��/Ҡ��>L�|-��^�}��nvI�Zo��mB/���+�}|�N��P����z��1����j[�Er}v����Y�6��>%�.��P���{V��M[�x}8c��L���L~���2�/4H��`k�z��z�w��_I����g�Ŏ'	�v��~M��ˁ���SS��!ʦ儕��`��Gz�!�V�Q�~WgU��ͺޝѺ���DdY��|h��7.}W�nɸ�H�4 W�����h�9,ɮ1v�<�%a�Ԋ����p�C��^VΒ�h�������i��\/��#۵�@/($��i�:)ܖ�&AD@��kK�Jv�Ѧ��ʾ��U�9%��E+�:��a���[w�u��@T�y���x^�o7��<��}�	��/v�%Rˡ8�O)�2[��|��0^�&X�vB6�Nk��ޫX;y�n[��;�������E/LU-?�{VE�kH���x�"��,��a�����|�e*�����Ę���W��;�8�.z�[���-����UZ�~��e�]�1�9U��p�Q��\&���ji�������9���gC�����_f;ӥx�Z����y�O4`��zW2���E�1�pS�ae��X۩k�bw��;�vTK������Yu�lmy.E�|p4H�M��#1�:�3y��Z�W�)do�q��V�w3���>�[�b�Y�.,��v�T��͡���=4�I��ç�;��}����}��U��ꔬ�Ȗ(V�_%�P����휫����#^��轙�;�29y�-��ooh�t�ya�t�|z�վ"õ���סX\�uS:+�"�m
�	�gz��P�Y�&�m�5����|�)I���/d���J��m�Y�!ϸ�	3�o�x)/'h�\�����]�k�=�3_1�
9�����Z&�`]�*յsږ������}su�n�uAƜENx�{�������g6�^��}��Rb�^a�\5w+�[��`Z�;5�'�v!�F)��M>����6*����Fݳ�:�}о����=��Z�	�i�OPg�U�$y�jO�c�B�J�7�	�����ۯ�F�����y�O�����O�ӱf �`i`��L2���u5PǗ��x��d��������OLб�ʮ(��6r(n�/;����*��ň"	#�P�1�������n��gZ�pU3l,�㚵]2�[V|a���U�3��<J��yPv���s�]�Ɓ�W�!�WExtJ���ul�ɾ-e7�["t�4�q	%]g,��N���*�z�Y�:Y.ƹ�ʏ�%{��������'��C��W�w�L��cPz��Ov�:�,�W�Zq5���6S�GG�^��3�N�����=tV���>��L�n,�>�ީ$z�|�A�t�����Bu������>��+5��g&Kz~�]u�j<�!�<{f"�N]v���
R��z��é�Z,c�׶�')il��\f|�7��Z��5��W�nL98�ގ�d}ѧ]�T���2Z=�������l�;W=K�s����Y��sm�MzwnMCU�[Y�'-��є�3�~ er�Y:�W�btf>1�W��Y.��wu��P��O6+ȹ���m�RR��c
��.���ЮaC׍=8�w;�現���[��os&������[}[B�)u��:�Z2]L��u����!�P�/��讈f�j�D���}`�Q\f��NCH��ۈ�s�gs�"=�]�8���4�I�b��yq�t�gbȜ�x>{CI��{��v����^z�k8`�={��)]JO��j��X�Z�������c�z{³��X�N�aO÷�%�a�P�]�Q`|j~�"{z�-���5ӭ�-x�\�}�������?��7�ΰ��uMO�ן(�Ԇ|$�t�<�����f��>)�s�n+A�;��G)W��<JVW��(���;jj�ק���4�B_�h�����1XV��k�|������K��� \�R��X.W3�D�S:��Y�y-��Ky�ӓ3��Gզ�4^�|�cӝk�x`S渄t�_�����ԙ��Q]��Nc�����ܥ�9�G��<���[�⟮�;��:>$�PӢ��%ab��d3����z|>�G��{\��kk�H��q����r�'�����0��u�,�+�ICWTa�M�u����H�xU�#b;���Ru�C>�]�s�����-3����x�ϳ���׆j�)�,�=\���I_v�$M��9�gl��ތ����%�OmXK�:�3���&oD&�׹���sÂ�NՌe`9v[&=�蕹G5r����uՕ TE3����W٠qE��T�n�Tޚ�9� �F;]%��5c_�m��uK�����Fv��2q�~�2��� <�Z6�͊��)��}O/�
7뢆�[���]����P����I��x�����U�׭�n��ϑm��l����-u���=J�:=�l,ī6���N����^�*c�]�m��Lg����Y����>|�����X�xJGYuC�V*�p#���ٍ�&��zd�^~�\�yi�{&33ꗤx��������7�\7H���m\."w����e���tn����
�{�$�f�
��7O�|�}��j�&��A@A�#~|5�8�l�e��*�]��#���a�[�E�S��V�I���u#{̩/E;���9���9�(.�1�;�;�pR����-�G�0q���;��y�Jy���ww=o%���}�=ha5��Pw�6���-,�w�����p�]4�����w��ʯWN�6gϝ櫵@����P�({�{|�k���R�!l�{0CC5^$ì�>W2����)�X����_����!�١�Da��X���V�5�7���/[�ھ-�Mz1Aa�rV��Nӻ�O��To���صJ���:�U�S��H���t�$"�޺�S����Z���R����M(�m��~�i��|Yt��}%Y�]�Xu��>W�!�ם5�S�xlKC�� ��u6�	"�`�"�{����D������	�^��>4��5�9������@�s�N�7�vz�^hezwƍ�ˇ�W ���m�	+��>.L�}��x�t!D����'j�[���r�^�-gA�=����`f峃sِ�u��X:Q"�b����J�⧕�C���.N0}RV�	.<���\5�y+"��Y`��虽[�*]%��|rv�U������	$����֕��ݭ���dTt��C8,�xm'�}WL����z?G�\�o��zKx�҆�׾Y�֟p�o���e����3n��f�tר9�϶��wݠ�E�ؿm����=��o;/��>�v��k�򵻝�Z��>��7�ɏT8�u�
a���y�}\��>���0zKx.b��{���^�$�p�Vջ�A(���תWU�	i��Z{%;ΚZ�3Ҽ"�<��w��j���)�J�!�k.�6���_x�K�����"��>�I+�*i��X��}�>__܍*�Å>�)�rE^s�2��yg}q3ԫu�;+ly-r�2�^�äM��ϰ�:�o�����]�ݴ *$�8�x ��g=�d%�	�(oz!Rq�{�ۖi
��ƺ��]-LuD�pu<����i�
���}~ވ]�շ����=%=;{LY��
��X��,�uu+D�B�	w�>��o�wl����]3�j]lg�eOw�qt\�L�a�x��]'��58�z��B]���ћ�uܭRe$�j��DHdw73�ݫ�y�!���d��V&�gؽ���B(V�6�,���>��k6F��O�>:��^�'���g9zP��3rE�խ{�78%U��fu� �/�.�(P��b���u�̚�*������Ԡ���X(C)\چǂ�O��1���%�/,˼u5P>���^�x�*�J���3�т
�j�∪���-��wY7q2�u��3�=S�Ä�x�lcٝ����w""���_0߄��0��3��8՘j-�U�8}U�.��(���u�8.��U[���9 Uga��;?`(i쥴r����=�|�DvN��y�y<Pj�g��L���Q�J�P'Y�U[��'��C��tڡ�.�A�mU�s����+�Qo(!�{`�wfcӭtQ�
߻�4zЏ���ʟbj]�up]a�P`2�V��f�g>��A�*�kE���|����4%
������9���Qղ�q�D����ռ.���8>v��s�Ó�����]u��<���A�:�-⣞��5���c����?OQU���&f�����t�S����.8=pX���+�K����D�x��׼����=�����A՛����~o��.m]ui��.�ٱ�W�P��P�u�^���L��x0��l��->��D�v���{ʸ�[K*m���h��T*�9ޭ�'k�=J�^����B�D���������ʳ���d��2�`��\.� ���&�جd���I��n�`���696�Oj��@6g>�g��L�+i6]3W��Y�GB����,or=~�f���n����ܚ\`�]z,�i�q�Dp���5�T�jx�f��ց���/�o���gƖT�{!�O�]{	0%�ڔ�7�L��<u"|���<�!6
kCN�13ז�n�K��Y8A��^{�WsR�FhM$֘�i�f�S6kJ��^=|�<v/�hX�0Q��%3����?s�{qX��6��̊��\�}R��U�Pf�,�r��r�����9�e��Н�$<�"��H�Y����Xg'ÔXQ�j1��m��٢�+�T,Y��
���ZI�$��z�GD���vNTs��6�y"�v��	s�d�D�4��Gz���y��_G�]�s(,�wl����<�u#�Vh=��q�G��Yi�ƞm-��Ֆ{�E��rV��
Gf�����評�kG��ηjq�uWu���*#��Y���r�.�݁of��8��TA�+e���o��},�/��i���Z7��C��a[F�˹�F;����L��p[���`ʰ�:��k����y��S&�;3w�w���k+�}�ܧT�"!�N	�9QF��Ί��Ns��_W}�Z��\�u�TgVM۹��2xѠx�O�"$���[9̳�'w:�x��lP����8������z2�c����3��ji*��c��Ɉ���a̔�ھ�:�B��+/$3��K$���˅1�����*;���wi��Ef-G�ol��g�M�eQ�<)�RDmа{'�M�p��01WH)�<��y�i�'V��X9������\\�62s��H���l�0�e�0ֹ%)�bz���9j#t�!���0:�g�J�MC��p�d���tμ*���n����յ�#L+u��W��/B�V�Y���)�	�9P�x�y�%J��m���¡<����k��m�ǘ�1s�W�(퇝6�Ҙi���KhՕW+y+.�;�ԝmc�|w:)L=�s�Ͻ��5��}�ê*�u�mYg'=8WK��g ��#R�����E_Ah캓2��l��؍��ea��Y��Zx��}u�;.;#l
28�^I,m�z���n�C��V+]b0:��8`�A˕�������z�;�����x�s4vF*��(ۤ�2LZ2��v�hc�DO����ښ��X&7���8Tt�2�U.+i�;���ϛ��eZs���wW�m%�1R��H���9�F����껴���1�ζm����K#�.r����ڨ�PC4
���
����&Y�F��� u�rm��+�4)�#ot8���q3�x!�W)�i��G�!�'�X	����8�f.�١�u���{�n��5}��ʺ���-:ۧ�R�)��x��9_S����9I��S�r�(/��*oί��+�¸�$�x��b��a�������|x�L=�3����=��j�]x�`��j״�<j�]Cm���MoI*c�Hn�ZQ�M�=�,F�:���]���v�PU�Ă�5�lgVώ�YZe'�N����a�1#���[k9lkhڠk�P���W	�r�B��2��vΦ�c:�!z�.�
¯+���	M��Q�+���C�&������u|���W�~ڜ����/!�m9X��Ԕ�}�:�l��X�Z+�I2�)gvg��d����ke�'s!hu|�s�g��S��2��I�TsK�V�:��X�(���V,Q`,�hT-("AE�E��F�jQUE��B��ҡKm����)�,QQ[j"��EEX�U���DQ��B���**��U0m�+b�EX�Qd��-�1�l,X����Z�DUV,X��@R�X�,J�V�.,�-�b�Ȫ*�iV*1DYPciA�VUAEX�IX�`�cXQ�+Q-����H��J0�Q(�Ң��H���Q"��H���� *(lQPX(�E��iB�\%`�8%m%H�B(��
�1҉�,X���DJ�%�m���Q@bT��ۇ�Ƞ���X���
)X)l����T�Y\7P*�k�I�[aF�Kb!mj�Z��H�kaXVg��5�����C�ή����n�v�Ɂ$6�����P������
D��:�7����fk�M�nb�<u;o�����٘��^��f�*n�jA٫�䙭J'r��mw�궳��h��\-25���VO>%��e¥S���(|H|ׂu�'^�*�KN'O�t�/=A��m��p;��k'�FF�SF�\��yP�XQ�3\�U�mN�%Xi'#�#.�S[��:�-G����ɯK�MTC=T!�^����(�l��~�[��h{gJ@}@'��{��D���7��U���%�n�{=r�݀�ϫH��3Ӫ�9�9,��~�c���X�Kk���ݫ:=%`��YB��A�7c��ߞ	r>�>���n� 'r���Ń�U�NMm=1g�9$�w�����C���#�zƊ����ma�W%��&�i��_gLOD{~�㪺���[;�����}�_�k��^��]j�`��j�X�Յ�<z�e�k��u�CŜ��L�0S�#�#�/uT5mQ������.�4��T��Ց��c]~}�L�CM�C���V��>��Y�Nv!1n�o�3u)D�Y�f��9]x�[�I�k��!���J��-l�����О�u��b�=��G���!������Y�<`�aE�Vp�R4@�h�3!г�@������~#x�� �Vkݓ/A�NC�*�Vv�v�-�5��u^�;�sk�v���GIJ��##�{Z�K�H���J'(��;�,�q�ύV��Ʃ��C��Mˢ�ծf�d^uL�	���v����;+g{x�C�`kL���h)Lŀ�0��v�
Vx�t�Fı�K���i���fZ¼ߞN�s��ƣ��.`�~�3ԯ�Pv��N���'P�N����k�M�t��]���v��l��Y���+yL݅�Y4��b�!_S{ #�Y?_�ֶ�����.��k|�0t�k�����.�V�ܯ�aCDKtt�,]j�y{:͜�LS�Q����cxס�����5�[r�]��z��gAϜ�Vd5n�Ze��X��������ߺ�ƺ��Vco��7-��*�ϟQ�-�a%r1bg�;�rC^4��E�p���X罵��#>o{�g����`�~B�V���m�;���)���9gߤb�C,g�x��{�ow����3Vؑ�!�z�I����C��6�E2����\k���N`Tk"��݋��w'�q^��nl�!Xn�J{{�]+���J��g)9��O����w�#"�N�N[�\;"�=�ɻ�簟/,��y�JϬ$��
�m�N�N�p���lo(%"x v)���qi�,���G���Ն���<'�c*-����s$��k3/��K��E'0oVJ�]u�ܦs���|z\�)kf����ΨGw�ղ�M�k��`ە~�-w���~����n���w���3������q��s�>whMF�͜�ǝ�EϪ�"��L�T-S�2|��8'����_��s���t���kzW%{�I�=]qLw�r^��mK�8�=Na��E��3K�{����.��i�Zr�8����I�P�r��:b�����n��\�Gbl�~�g�B!����+(���	fWv�9���n�\�w!P���-�e���r��*SI��C6�x��/�!_�Q���z���:t��ƽ}��%���ȗ�
��K��+�:1ݲ���I��e�[�����bۍ�:D�B��2���"�Lj�S��Xg�`N�
ϒ櫞 ���;�]I����{^����Y{�J�ș��z���ǻ�g�M�b�*�	2�5J �L"G��W^��	���vSU�^;������ֽ��}��fm�?K�c&\5�T'����紦��%d~}�
^>R��e�ڵ6���/��0�JR�&�w�]R�y���^i� ۖ�8��:�`p�r��Kv�޺Gk���gd��]�4"7����4���V�^=�;lK.T�F���S3��i�s�W����m����Z�%�k9���N@��f�t������ǹ�$7��6l����/e>���L-GrZ�\6���KA�r!|6��$8�O�Xg���]���Oolykz_j���Y/�v�b�t<oR9EX�R��7p�^m%���g�O�Lx/�&eѥ~�n���| ޲Ye�4��H�������qU��,�]��R�|}5Z��R�_��O7*�������LA�s�e���Q�%3�`yCX�d�������Md-��/���� ��Z��zX���a�~۸�z(<l���|�5���;6g��߷�T�G׾hǃ��u���"Z��[����.2ߩ���A�b����۱�D�3�o^�YVmG�Z|��)mz��ts�Y�%�]�c�9G��%ykM.��3�5#���܅���$��s}�B�u�;O��+Y����~P�F����L	Ւ�ڳ���~��Zu�#{��>��C=�m�PE�mpj�b�v6R�P!Z�Ph��z���~Xq�C�K�>u;1��^3�+�`|j9��f�Oo�3���S�L��%�����(.�� ���8���~R֘�����)N;V����s�l�F���;�ֺU6
��C7u��� v�{0�+g�f��:���T��.y����ᨽ|y}��˭͜�Tx�kX��  �w���ۚ$���0�[��68����z�m�RH��)SgV�&�B��)�v5T��<�EsMC���"$�y蚔�L����̿2��L>'�����Z��h��>N�&��,)H3u3�?�<���y�y�B��kS�n����M��C:}�>��
��~�}����dY��͝�5O�����w���fz�>Vt��Ӕ�{!��c۱Fn;8�`B%A�*�D��i��\�9��adSP��W����K&7����x��N4��T�!�;�jݚ��jL��Ԣ��׾Ͱ�/��<�������Ӌ�@�L���S��>�o�2ѫ��Br7�\�Y]{�OT��&b����<8�H�=3xV��q`�jg��"�JL�ļ#5�J��az��8��I>�`�S}���w�)��`�}v�'9��e�^�VCռ��=�`�^J2��֭����u�ܜ�G�f@��Z=ֳ]5c]�ߟ�yT
��}�ǌ���
��W�zO6���}���̼d؂ϫz��i�K+�����k�;���<v<���c�^}^5�sˣ�3�D���|*I�7��`X�|t\Ͳ�ڋNe�Cwޞh�w����+�Mv�!���\�s\��j�,jy[WF����"�g����m�@�������4���Q:Ԫv���d�^'y*I�pX2pL68�����t߻���x7�&N���[^#�[��Oţ��*�_?y�[]A��m�{������C:�^Aī84ӶC�>�u�'k�d�7���AW�,V݈pR�DcWw����{�V�7�������wL0k���P����R����Nw1AaB��ˌ&���4;�Э���_���lP�˅󦖏��vh��5S{>	�r��3l���:�w�|�_�b�
	�yi��\e��#��|l<Bc�i�^��9�E��-f�;5��S�~���!d����=p���u� ��r��E/~yo�v�t�2�Z��]�.N��eO<[w���`���X2�gS�sH��1\�KKu�����2ϴg��K�L��#�g��6�n��K�\���0�&��h�����%�'\s�of߷���Y�G)���77�N��՘�n�Ü��{4�U~Zd
΃���B�[5(h�҄"M� �71�\׻=���}�Z�K^/0�q�xm\O�"����J���ꏛ����_�'��f�gH���^:J�Z9_ozq+�<m�H=��9{��*˛"�g������{�%79[�����.����(\�!�`��v�qs���(�D.�M�}6�@9h;.gM�������'K�n��xWV��u�M��܅�a��{'S�2��O>�=fVu9a�l|���a>t��!1��긳�gϜ����u�{W{��/�p�y��$pҟm�FW�3�
�dQ��pѰ3r���\S��6�8:Q"b+����)��^5�}�A�>n�J��,�9��zY=`.��"�D֗�qvf7Ԭ���'Y��뻞u���e���s�#.N�Hg����{��j��ެ��Y���f:Ŗ��W�L�>q�����POU�ﭘ�L���o`�{i[�9k@�^;R�������'^:ߨ�ΧO��o��������#�u�~�e�w�s�\\|9�`dw�x:���Z�8��2���<$�^~��^��.��1C��P�u����s�>w��6ឿm�w�1:�c���?|�:'QvZ�Ǫ|��=KC�@�+��Xы"Ϣf�^�݌����{�7�Y��;��ȡ���
~Mjc�%�����E����A��i;b�s��ޭz�;[:<�jtUܩ�ӥ�Y��Z������wl�daOn1^��&mFFN霝B���1Y��	��5����#%�00֒�FT�yQ��C9p�K{Y����u��ɣݲ�y��3�n��v:B��t��h���1��mA-x9h]B�Q`��T6�R�Y�KWʃSqc�����D>���Κ[���D&����.��B���0X�-A��>��a�A��O`�e�cc���w�����ܦ�3b�dP�<w�K��&z�͗�xd���J��hjD�_rYDZP��$�[�$@l�i33���ܑl�k^�Ϝ��C�]��?K�u���|���[/��D2)&�wr��@��`�^��<C;K�*���b�O Zv,��`i`�^"[�;[�f�z7�=�/���v����dˆ��U�af��UqDU:F�ȡ��y�d�F�飃1xrT�'G�X�Mtj��YBq� ^�y�0߄�3�%���xPϵ�ᴩ�yt�Oc|�<�tH�[�n՞:Y2�,\I�f����J���Lto�b���5!��Φ=]��mn=o6�1��S�yS������0`�d��e�TpE�R���y�����r��>=s�>����ۋ�i)��z�2=�L�P�Px:�6[�Gӫڸ�-8n���{V{���W<nɳ�v��Ő�����?ߩӼU���h>5�Qq�8�8��^)�rc�mn�UA��X�yb+Ǳ���+B�k<�¶Ձ����X��ʫ+i4P�'�I�I�J�΍�X+WAήL뮫��;#��b��(ஜ�mà�ڗ[����I���N��Un���|�M�R�/�m�Ck��gN|�M.#�:n���+[�)?�łz�:���0ͨI^\[+wr��򡂽��y��<�SA�Wj�{O19~��fS�n��*��}ⴡ��hN^'�0�t{݇s]w�ό<��c��<-�3>��9A=i�=J�c��?rL���w}C������b��n�L���iP�ٵ�2��rdŴ�=]I�a�:����p�[�O7�@sy�˸�5+�e���N5�G�S���J��O ]�K������p.�tm�Ns�1��Šhϸ(|���a..��A���0�/��ϳ���v��V
�>�:�~�7��?�]ǲ��k6��EC@�U�J��|i�f�S6ښ��׼��K+F��A�zH1l�r�T��]�jƼ��Xp���\��M5�r��|�(XY�_���OBk+[pn����ڀy�e�ޛ)k�������h���3wԢ��ƻC�k�,J^;�U^������1\SB��:��*�3L�:E�6Ԥ�n�5	����e��߯��)Enฦ�����s8Ljוg!��s�m6��6=��oM�V��3\����Ӷ9Oe��`�?r�4q=�02;EՄZ=]�n�ب˙t����w�jT� �[U���;�-O;5T�y��釄0�Z�$���xo��x�<�V�U�B�̙臼�Eڍ)��_yר ���~�"�xx}m$,o�m�\���ˢ�.�S��^;�
�W�8un&=�����-3��~�F�гk�=um{�����;�v� d5����리e��c>���*�[�������a��*y�͍a�$G�;lT��g���������Fy[�w����٥��i�_��^��/Z�+	��q_����L�^/6;����Zؼw2�#�zƊ���)��/���YGS�̔m�;��骯ܳ� :�=~�U�W�C�6�˭o9|r]a�
�B�n�1Mx+)����Wz���8�P�#h\��e4��'��Ϫ^��������7����ۮ!�Q^ٯ�Y����� ���R�*ء�8P�󶕽4ϧ�bf΄<��q��s�N���s��p�MqϨ.��Uq�Q#��|h2%���ir�^}� v�/��p{=�ȳ��4�������)�V���\Ύ	�z",`������W�}_U}�����$����$��B�XH@� IO���$��$�	'���$��B��@�$��H@�$�	'`IJ��$�$ I?xB���$ I?xB���$ I?�B��H@�l	!I��(+$�k.`E���B �������+�`y*�T*��(J�ED�E@B�� �IDR�����x�U��%HTْ� [j�j�
�"����T$!�aJ
 f7�:���FUHT�R*�ET�UUI	J�	P��U*��P�@���TT+� �pD(,��@ڶѪu��W]��9�VA	��֔[4��U��*��%WX$"W  �����q�d-��JU�f̢F��t��k)���n�	��n��9k�)m�mm��;M�a��Tmf�D�� ۊp r�    9�t
   ;��   u� �ke)Ws�T�%�m�V6u��ʬ�j6�T�@QU� 6�f�Rҷr��k(��ݥT��MeVm`�Kuݤ��e�ۭu��̝vX�"��*��T�;��*��Z����-6�ՙ#�:�´mShm���MQ�������P�D� NtH�h�Y 	h�Ri�U����M@6�J��8�
)��,�@IA�$ �f�)���(M`Q`��[6���[���
M�0(�d�m`�f�Pl�V��aRمR�ʡle(U� ;��4�V�h�����J&�����& T��l�"�� ��i"Ҳ�,�а�D�K@�1k	$*ѤP�}��   &%J@210 ` &Oh�JR� `�4 &�4h`F�����@4   4  S��*U�L��dѐɂd���A4���L�=C#A���R	4�1%*�R 4�@ i�&6����â�4�h��K�h�`1������DTY���S#������ dF��
#� 
�QO��*���?o͏�������T �@�`0� 
*�� �B1VDT�r�	��*���=���*�m�Biig\0լL>����$�Ds���y��������ն��_�"��զh�)iOr�ࣵ�mH�h�a,����usm&�?]<�Tځ8*�G3'u�5�(ޔb�Z�Ż*ނɬH\�3v�&�=iQu�-�k4�Ԋ�rB�7%[�a;����,Z���cT:�8��Ea�xY�:b�wL�B8�S��T��F ��yPL�i��v�P{��zt�ehգ!Y*i��܄C���wz�xr]3�u�l��Kf��r�u3&��z����R�����.�<q�t5�&Z�hͩwu�������=ϓP���Y�Ų
��Jh��i	7+vI�3nJ��@���-ޛ
��+~����J�Iۏ3uu��^[M=�����F��u�PaԾ���ai��nYUl�����#����Zo!ܢ���m\zr��V�0��+3\��2�x�u��ʐP�v��&-^1y�V(���0��i1�d3��V-[IF��1���RK&bF䘓��[��'���"˸��)�-Gq�Wf�@,���G�+]*ջi�vkR�^�\$ \�Wp��]]Zh����ie����dM�(��2�%mazf�n���V�VZ����P�x��j:EX�n\*��ə5�7f2�czU\�H������0�}w�n��[t2�TL2�V���T�ق�2��-,n*w�2�Svi��8�^P� �ب!���n��v�v�y+\��Bӣ@��*�$؛/�V]K0�S���T)�����vh�JL�;l��
���:�3F�i�Dvٗ�`CbN'��Ifb�,&�X��"[��RQFM���-;�-�k@�ՃV�ׅi�c�èm(c��F���T�{�J�*�]����.��o��@���y4ν�.S����E��6$���Y[���=�pmS5��v�"�n\����V�U�u�NEX��aL�ME�J��7�]5��F`�����N�����p	i��X��3u]l�y� �XY ����+%j�5���CiY�Kژnh�%ܭ�7�8�H��FN�Ǝ����ݺ6L�*9����ʊU��ښ�6��Q5y���c���%o#�ja�	�O6
[6����dz+p�O^���"֫IU��^�AEp����yZl�Hj�mY0X�sA�Tf'DmS�,�/B��cAv�r�	�m�cp\�!��]'�
�������� ���rз5���]7�j�͵H�{-Ł�s�O#q�b�xC�j�;FJ��H@on�n���Z,���%JԆU���f��R�oF�]K���*�82<�4��yuE+Hސ�}��tSOj�6��AP�b��׹"�d;ٌm�0b.J2^^QY�n�UUIy`جX�U*\��TLԓ�E�Š�YY�FȝQ�6���pi=�d��[���P*���4}/�W�XS�M��Җ�t!��6�Yν�:Tx�1-���䙕���;9�P;��-���DM�!9���3�3k#�d*cs\����;���FR
g/F^��]iRv���͐�.=�j�B�V*ۦhV<N�Æ�6/˶�O��oS���m�' �� ܢ[�ݍ�*[W��u�	Dɠ+�dԽ�?�'��p,��V�v�=��`9�W���L�.��ٻb3)!�+*&m��*<�c]Z�Wɍmˏob�F��CiLSvŸ�dN��U����r�����pS���n3���*e˱rk�EeC���mt��-Ӥ�
�qÆ��ta��KkRQP��ŴM�����O�9��ˡ�bԆ檋qdN��Q�UQ��έU��!iĲ#�3oCx�qBm��S-�3kT��k)=�U*؍�v#
�E*���Q�%�80hm\���h�E�ն�5=T-ٻO������ʴƥQ9����J�����Q�)��m�Rl�q	KB�3.���r�6��^���c;(���Tr�T�䥰�I�n%4���z+I�2�[J���V.��-w��Qu�Z"G���kkHG�,�F�I˗X��~T�}��C٧��ʲ+S2�m:��Ե�J�`��R��C3�����,��V�ê
�փ5��H�,��W���hr��O%��[���)�1ix-��*v2f�'4ϒ��Xo\��O�������]VGn-������b�K�[�^l�䩹E꒩���=LZ{+,���<�#Ph+e�V
����v��� ��[An��������ֻڑȕ�Æ:��6����W���%2�g�i"��� �ĭl��Tڶp�+',ͫ���V�RK7l��d:�GUT�i�d��{�d�1К�ٱJ+hR	Qi�U�j��peV�%1z��qn��e6��%�ĵ1�UJW��Ue��h�%N5*F��w���E��bጰI�1B�%ZR�N�hPK�j֪&��:@� ��j��ٷc$.�q�)Q�e-�pQ܎Xc
�Vj�wE^��47�<��=l�$��3NY�YV�hǧ$Y)����!ض��ژ������1]��I�w�c�'^�mT�NE�V�H��e3��gjT��ʎ�����X�j�i���³3^�ޢ�Y5��
����[�SX�f*�2��
c6�`2H��2nR�U؊���Y�B�(J��vMȮ������K�2f���횣1Aɣ	��؁��ɈՋu"J�If��5Rص#�n�4]��p2��V&#ztۆ�c��-�P�4�4u���ZHŎ��.�r�����LWum�N&n�R���f�%`٘[�X��tVk2�r�Ltej�2���Zw]V�j�mJ"�ު56���L�Xb;UF�%M[%�;�������CeX���t�F����ńHjk�ǉ�E�8 �*��̆�i9��ͫ�"��OQd����Ub&T�*�arT�.���-��՝�Z����i�5��{���(�n�i'��r�h�j��{jZ���i�*&�N1�k���*�2�	k(?����X���/�x�)V�r��(
Z����F+�hDsL�uʭ�2��T�5M9��en��(Tڱ�6��O�u*=��N��%����b�cs%n嚔]M(��y��͒�+?n)�(JX�c���j]���mAi\���,�8��c��R���RHBљ�⒗A%m���ͫ��t��j�k1��Na���� ��:H��N#Kbm���.�k�ry`Ҳ�� F[z]���¦�D�n	��m�ڛr���"6��l�3]�ujZ�y���b��W[�\^��`l�h:�W5�T�������e$U�̲.eC���ܕ)�ϋ*KUYs	P�Ә��F��øc���t��-�2�e�T�r�,f��^X�^=�U���-KR�?��E�j�����l�f�4ݨBv,(ҫ�EG+���r8�5����{$�X*m[1��)�Ec��;I��#.�B��E�T��r�c�x��n��Ly(�B�Q6�mAK�E�c_Cc �+T����#R�vڬ���j&QU/\�R�^Y����1�㩠����NU*�w��X�K�2���h�1lm�H�>�3)1�`���Tfm5�H&�nVn�r���j��7f��Y��een^RV�`�UK- a�%+Dm]���J��Ua�lk�ou��I5]^�C7CN�Wa�KZSԖ)2�lߓ�/u�#RӐ�78v�*��������L�sB�L7�ϊ�a��/mL��Pp,3EhX�D.���2�MJ��Vታ�i��/)����L�PX���� *Fn��v-
Uw�	���1��9KA �)��f�גn�2b��(�y�bÚ� ���ۍ�!���9�]jN�m�M'��n���ն/�Vͪ�2�R�D��ZaN弬ʪ)�9$����{Y�t���vub� i��s`�a^T�A֪ui�]��+x�V�Y[+�MB�i;���9l����
S�/v�ZMQ�G�?��|w��?���9�}����I$��I%(D�I%. ��Q�$�)B$�I)A$�IJ$�IJ	$�JP�$�JPI$�R�I$�R�I$��"I$��I$��I$���I$��I$��I%(F%,+��l�.J��T	����J�ʋ�50+�:WX]����ʜ*���'�W�_n��`NȀ�8����Z�vo��3gP�ox1�����)U٣�Ǟ�l�p.g�7]�t��%�}��s�0a�u�S��S��K��F��&��:Ʈw��M��܋d�V7��#ip��+z;df_N\1�!G��r��Oe�h��ӷ}ӣ���ޔ���ӻ��Ʋ.ra��*��u6�H}R�	�8���9ޗ��,�l��Y5wfS�ޒ���3�8�yo6��g�[��I �c����˨��W>kx��}*�kKJ6���+�lFr��eRkk �q������vk�ZIeL싛WM�%�'�qE�j/���Z������W�k��;��L�<&��¶�u��Ky��U��3¤��͗�)+�*�d�2��{q��ExmVC�$AC�<8 ��F���i�<k8�n��tqaҘ�e���`�a<��|���u1TnE���.�vj/��?8*���Np"m��+<�Ѱ�2v��4
qu@��3�gA#+/��[�BK0�L��s�0d7
�ɿ+��;4�Ǹ�O�"�[�V��(��εu�i;3����)fn�%����u2ZtO`��^kj�.�:<����m�#���	�'Z(�tE�5;:��Qc^�{V���Gۖ�tQLf�ԭ٪eJ�=�y\�����ъ��wɊZjȣ�.����R̖ c��C8)6�=�NV�
�]v��R>�;�DU��3��ˁ%��)e��q���il	I���.ts����_m���;��_	�ei�CwM +v�q�� ��q�/s�y܈K�V��`e'�W3��q3�B^ww!���G
���%D
�2��e]g���$�Bĭ�����ozf����d"��4�Uwʓ�s���IJ�+zVo �Tj��v�U�)�p4&G�=��Z�"�Q�c!V��Gϒ#Z�U�>.U�ݙ�R���I�3���B��u��1�u:t��uL�����맭Iʻ2���sO],Msj��Yݫ�%����7��y�8`��|/r	ʠ�2]oK`e�Pfj^*�̗U��,��q%ܹH���TY�i*�.���!�305:�b�n����������-�m���V
�*�u���A�y;tW
뾮Ū�7�S�4�����C�r�%��-9�!,;T7��E	�RP�i\�Yx�@�*1���&�7\�	�������4��F��Y�.�3��f*�{�Wg��i.�;�O��I��*�מ�y��u�J�K�'M�D�r��4i�n���9|�N��]˄J(����^k�}���َ�O��]����Pus�xi����G-Y��m��N�v���Kva��ͤV����$�F�d�넎���#ƍ������}�lʻ=
*�ڵ�����UgV	v�Icx�>;؄�ɝQR3n�Gk�>���ö0\��nh�4���=oupob3d�q�}E���^�`a��Tt�W&�AWѢ8��K���\�����K�P���س��Y�3��ǭ��k2�Ю�)�g@k�t�l�ԙ�k#(t�r!�p������JΡ�̇)��q�Xq�u��RQ��;o6�� ��k)�㶾��p�o^�����=�y�]��.�z�b����C�Wc�8-j��1���r൸�W��-�n3ݛ[ �v7����3
�XU:�Q���q�n��u�����e��s���t��}JW��	0�Ƽ���R��Ӽ�Y�N�uc��+�ʈ�~��{B��Yǵ���.�V��e�p�����]�J���ce�bBF75�����1V�I�.���u��)��08;ޥ�J�5�A5�����t5�E)�/
&HI2��r��՜
�D`���ڽ��omfKw@u�˞)�w���>�G%i���K��k�w2[��R����.E���]�m'r�--9���Kn��X���U1\�fb��7D���Z�;�g���"�6��]Q�c��)n�V��Y�:U�9{!O�Z �N��Sb��U��>ם��U�5��p��Nd[sC5�&m�E��s�ݦ��<������Ӏh���;V	2��{׋���
� [���ۏ�Gr�ƞ9��\�]���P�2��E�쬎���S����}�:�%Y��;��%�@�ո���Z;jiRG{�v���;�Vy�.�6vG��s�,��3�VoC�L��;%uq	��ݫƍ�.����v��&�.U�R7��
�zҬ�5�%�[1����� �36qd���Mʑ�y{;�,Qm�5՚%ȫ�e�PmC���K�I?�v^�zY5p�UN�'oN�wE������i��m���%ѥtT�Qt���]��!�j��қ6�[<=pE��F��u�Y�YyyYe�S��Ӯ�pJ��JM�ܮh:�4���X�P@��M��_7�]/��F��-䗟L�zD@���++�kLe�V��fw ` h=T�Ga�*��I��/�'m�̑�B�c|�9�S�4�N۹��p��sUl�U���/^�Ŭ��AyO1��ai�Sw5�Riu���Od�2^��kA�J��^]��q|r��w趤sj�]���dzc5���L5_t۶�(ǴU^�K��bL����$&����S�\��U���k��OE#=�D4��z����.ᕒ-7`�ٿM�!gn)P��+t����J4>2���4�sᩛ%�t%є+z���cGj1*���<zv�В�N�������V{;�呄��-k��;��g����r��~�q�Cu ]�$](w�����o-}:�vG!�G�͋���
^�ˈp���S̎ﲍ
���L�q[�V𹸰XL�+��.�SY<�w��Ԧu���4���R��2���d�v�ޙW[mX�RZ��W!��w�u;�* Pѓ�r�W=4�$��%=�_r�����W��r%g0q0���(���q���hq@�n�\�Ʋь��.��iШ���J���q�v�E��3�J�_G��%����$�՝�l��U`��c�p�Y�EM�$2#6*���3)�r@�ͩ{�7)�PҮ,W%����d�A�r�NZފT�op�� "V%<':�HP�s�9��d���,Kjg�u��^]ȹװߡgc{�o4�'>�]fn�J|�+�g���\�D�EV���f���ua]d���2�JI˱�.��w	U�O��Z�������utcuUb�Kr�M�'M:9�؊a�#����o�*�M<93Bu��K]��=G���Tk�H¥����AaJw\�e�؅\S��}7sC�����pNp\"�y(�l�����5���XK�wi�
�&���Yx�F��RwSr*�^��.�Ǩ9��|����F`�Y�Z�n3��	t�E�����*zkw���]gΊn�`��L�4��.�X�O��m�]�V���r|z��������F��r�S ܽ��`�8��;YQ�vy�*]v;8L}���u͋t��c)�|��PO�M��k/z�N��Av��1�J����O�0�7���"�|1�C�#ˤ�Y��>7�]�\�d���{k�9{�� �Y��˥)OTSj�F�� �r���<u��o�1�D�El��גr<�,����Gn�ɼb��t�B��$�<�&�tN�{��%���H@+9\ތ��T��jڽ��Q�-��)X �x�%:�B�$��RZ���)Z��T�ҍ)E-�Y�Q�S]s��W�$�"I$��I$����%�&H%%1&�A!w�| �޽���Jך��ml�(NU�>r�M����&#���Wv��=8�ޥx&��Est&�<���"S���sb�R����GJ�q@���w4����%˗uv�ϧ#�N�{�PSj滔�I�Æ�չY�J�x�ac�1�c<�c�1�w���s�l�Fs;d��(�a �i�Ȫ����0w�� ���x�/p٪I���<on�c��C��^��*Hmr��f���]F���� e_#z'��gx��|q�6 �9�/+��`+K-�'�%��ݽi�p�
��3C����-	f5��y��p��Hb"��r�tx�vr������m���;B*5D�Ǫ�N�r�4.䳔{ꎮ�+�F��Zi���У��ʇ!��o�3��ʫ���n��b�-�fL4�U�]l���4��|�滬��)㾪ۅ�}�M�|{l��w�p�/�U}���T&�BiS�F�s��vY������:m�UD̅�꬇]�v�����n�W)-��+  ���0�з�����)��%�O�����6%�z�]b�S�j�;/^��Җ`׆�s�K^],�wO�in�4%�vÄ�W-�V�+�`^���KN�����u)&gII��ٝeKKO_
y���gN�ͩf3�c6�kMSn�g㹩)����j�n���c���pXd��g���7]S�TN�fN��)G%�w+�"�k�������r��m��UBj�eH��L�}A?�]�m��K��W	�ni��ЌoL�|�S��'������6�ڠE�	c�F��SWQp�->ov�*L�)��u����
�Ɏ��g�i�|�QM�׺��`%ҝ���(,Y��n%�x�g畕�9iopV}��V��zk�om��<E�ݜ9��q�m幛.����bo"��I�XϨ�U�m�VX8IK"���FUө����V�NW]��c[�D�et�D���J�A[��q{Y:��/.�|�L�jw�yh�F�6N�K�|�b�+9�5��e�қ\��y��f$Y�5��	�5��{pP���P�����W*�{�0�Pd"`��&l.SQ}}yG�����5V#�tM2�Y�~�	h�b�(VX���תV��q���3R���9�X�.2����-���L5�iK�ZC:5wN�PܽV�U��/�5�u�K�C[c���T����
�۬"N��2�8so^K���pC;x��;.;�7rA&d�PKz�g^��7";i��ho�RL?��d��*I���;*Po��VV�%�Ѻ�4�Ъ�g\�v�y6��j�S���C�#܍��r$[df�����ƤM����}�X2�'��*�4w�=0�\)v�[2�iK��/�5B��jz*_[淝J�©XOa��J<B�(�
�E��g��x��Vu�X��}�
�u��W��4��E��Mďt跠�G���,��� ���]�ٖ1�"ڮ�N�jd�N�)��B����λu�փXv�f��r딮�wmNb&��K��!gJ��{��ܣ{4�ĸ
ڴ��?oO��CGq�)�2]tb�����Q�۱�+H9/t��>0v���fc�����-���$:�klg4�	Z	F �a��뺕�p]��U��6�4CΓB`�qS[$4�$uv�[��A��im,��c��ӳr,����V��u���3��Ar}���f�,[ˬ@�sEp��g
��w<���fmatc�����E�H�ŏT���N�oG�Ջۭ�`�����Ѷȭ��E�}v�ͤiK�%��*�{qJ&�%92�����F����w�6��`�����O�.WQ�NA�NT�Mң�����aK�巔>�T�:#!����K�����rk���ѹX��^J���6��[��)�Ub��ȼ e�ͬ����7��X�MQ=(�� 0@���5���.��rv�tS.e0��7Zĝu�}��D
�N��iuV�G��7!�\�ۮ�Ն�h�n\�Е3ꛛF�ĭ �[��Qb����`YDՅ�9e���][y2��o�圣.1: ��������B�66\��a�,άn���۹�`놗mV�NVe�t�.B��E�kphË_I����]o�N�1�A�eN���q<�.��nh�xDp-��a��;�Y��=��e� b�ަ��
V��֜�+_Y�9r�u��}7�e7{h(�
�膻��F��Y��u�Jc�`�O5sA�o���2�5b�}�WT"bJ���}ʯ�3DqL�	e�$�8���b�����{�-���Fv��p�����Q_w:-�
.�3ewvR������''e����E��bb{Y�J��t�o�v)Z��J��*J|P�rd ���a��+�Y�U���ED�����3fN�S��5�E:�9Uκ7�7�p�sr�9Ԧ(�B��2M�[t�&�Χ.�2�E��Ol �ꙙ���)�H�V+n��@��X���_�X��(�UR��uUaݫ@9�h$�պ�9�_;]|vD����3y���d�'�c�]i�ʻ(��kǀ�oZ݁..ܚ�vAu���z �x�Eyca��F�«��v���\j�()���d�ٱ�ު�C*TD�$V!��vf@�v6s�o�H���C�%ZzE�Z�$��V�h��=���oiwHe�¢�b%��%3c�@�h�����me��ѹ]IA�ۡZ�,�i�XS�uݦ���[!��儾�u��������j�͒a�Xv�8��T��WP��Ek5�ß
���:��%}UO��yp�1�̓rNRu:Ⱥ�Q�W�
RUd�`�|��C�Z���{t��9dv�9v÷�u�嵽Z_�R��g��2iWϳ�90�ɭVJV�u�g�\�����od�Kg#q��*���Gx��4_ �@��n0u�<���	������u��e>b &��W)u[�&Js��n��-t��:�hfn)Xw^�@����[݌��|,b�sH��:�u\��'�lf۲2S��X�yEU������I��q*y�[���ԛ�^��D�{�N�L��3W�����B�%��cBu("�V3z�)Ӎ������u����� ��)�}��1mn��MBн�z�0��&::R:*�ϸ7��̯�v`*��X�xj��kBUΥl��J�+����;����*o_v��3Z3c����ۧ#�Mj!�4*r5�Qe�O�cu��Hq��V]��P�:����7e�uݛ%��;���ޫ�jj�З����0�IR{K(��$��w�H��t�k�HfU���p���1,��k���:�:f�Y���ێ�'�u�3������$���^ne�]%73V5m�ܹ�}׵#�c�p���e"gKw�xu��d�px��e��{R�s6��ޤrb�U�k���4̳��80V�%4a� ����=n�P��j�3+2	CfT�p�IGE+ᚻ���gv��#�fu�w�̝#��I�W�v�hlBe܆����֫�e+ÖRuFywG��ݓ)����d�E�T�o*v���q��!.��)�Љ�Vn�֯E���]���u�� ��:�s\��>K��3-wv��@*�h%'h¡�gM��U�"s���ݛBLժ}�l�Fʩ�l��L�og�
u��b�ܶ��uUQV��[��h�:�Q��Ml��J�c�\9#O��xO�+-�;M}|j��v��Zz31]RT���G�k�*_&,�w�)�ѷM�FƯ�0N��U�?\���Zߓ�e�V+w��6H1��n�^ކ�Y�P�����KHڐ3۽^󧰐��'�v��vFn����n�ج�陜��=�ȃ
��RA�%��;B����\�^�Qv� �<܈-�:���Zқ�34���*�����V��-�Te��:��z�n�JA��!f�E��.B�)�Z��w�	��uG��.�t��{&�K
T��KA�3�E7�'^'N�;ׁ��,������O����Vִrɶsm��Y�m���Y�37H��df�]M��]7���)�M�͹�Uh�o$n��se��*���:�jќ)J׃���fbY��Ýgv=�.����n��M5��n�8�
�E]�I1�OR��L!2��5�������J����֟�!�o�)�'�BH@E���d�onC�$��F������;���w��}}���܃��r����Ӽʵ	�ޜ�Y"h��Ht*�P/�Z�Q�6�d��Xi��4���� �m�طK�m)=g5규5Pi�ctU�(��l�c��4���ݑgp%R��lT-0Pt@9�J�U\�|�֮��E���M7ƶN3����>�6�)�gn�R�@��W]xe��]ukq㮹�]��g;sYݹ:$/l>��+v�Cu�5r*�^�X}<�nn*k�[�'��Nf:&�о� >��oa+;y��Nu5�Z�a� "����ҹW؁�ALz:������#w��;��Կ��ϙ̇���:��4��*�y5cE��)ib:x��j.ǘ&VC��1��1uc�j�g}s���Zc��M��rӍ^������@	��/��8�$Xw
�c�p+�h��Y�VZ�݇'U�J� �_E!�J ޕ��u����}����&�iV��+�1�)~��Uıְ�Xζ3�,QQEb�T��j�aW�GVk �b��ɍr�Pؕ^��'"Dv��F	�M�-�0*����AW&+��Kj)�2�n
����X��_R�+G���(*�ѣR�J�bZU�Y�:�,DYET~K�E�+%Cn(����Q�"�
�VbQ�nebe;�!b�
�Q�b��	�$Q��	U���ji
j ��+R(VUD�*��8E�J�%�>[�lE���y����[XUM?]d40Qa�T��*��D���:��9��T�Ѱ>�e�/ff�Q3/sK&�ͮ����&UF�k���-�3K���6�d�IX/f 8pk�S�O:Aյ�O����Nۮ�)�|T�ǳ�:�+-#��_��}�_�����gT!d꼠�qx�q 4�A�a�۪��"U���l��C
��6�iE�p���~�G]�s[���
�ܕ���pz6�w��G�a�J���L�x.��4��iTE�6����vX\�u�a�*y`���E0�(���+j2��;�q2�d���Z`D��T)u/
T�=�&J����x�ŵ�6�R�[�ԼB���*���wE�v�?�̺�v~��A��� ��N���^�Y�d5���JǛg�A��̚b���������E�������e}����\�*���Ē�g��bot�$`7�r8r�.Є�G�$��̜�hw.l����y�Nj�D\
�k
�hnݾ���$並�(W�\d��$u�#h��+"�*��}<���Eeb���^�M��M�+q����k ���>:g4Q��.��u�zE�i��s8�+�.6N���"�r�����Ye՞w�]�y-0��J1];�k����+u�[��f�6��Y�3P��.'���K�_>��g`�%g{�o:�5Ɓ��%�S���Ǻu��hy�꺬P�/Ơ������HC>ZH;��Wm���ړ��N��䞬Pn��Ҏ���4d�u�]9��Yۜ*�'O>F�I{<{|��X��]Ƣ���;^ŧS{B21�H���jNXi^�m!|�n��v�r��xM�TMg3���Ϊ��y�+%�r���]ݵneXYU���1�Wk[�YLt�gEY\�HS�%�;;�u
����,�&�5!�Z�Dh!d�X�+.{��^�|���5�3{|2IB�BL^�')��˩�ʐ�um{���˭�#���ފ[�Q��X��W�/y@��wrn�^��i`��=Z��B�_��5���ᕝ��=�����YQn�:sy'";#��קX�ڐ������Y|���	�Y�����:�4��+�ѭ���Vn����L�-1���?%�c֞UX�e�Ѷ�u�S��;�`\m��Û���;��9Ǔيo*B9}ON9��U�᝙Օ�L�{���h����\���wv|�l˕�QOz`������9�rr�`r;$l93/��z8��;�RQ�Y#��]�4�٬p��Ho!�4nU
hm�$VV�ZW�$�c2i��O$��QId�����O\���1iU�� ���ë w1i��ڽ<�;�8���rivL�jJOۺ��vC[���uyƦu
m=[�2 S�v]'�N�<�b���D_7{�[6��s\&e�M�u:�L�R:9�9R��0�X���)kM��ꊸK�֠6�	u�L׉*L�T���r����C=�!�i��i���G�ּ^��u��u����V�@]mpw�zᯱi�!fMcv���4���M�l��#M�Շ�r�_!|���1E�a�gvzTu/����> �p�k��.�#�\��S�NE毐|��ȑ����ix�C}*aF#Ny
6�.���Z$ȃ-Rw�Ө�*�7&F�Fz�|�HY�B�</�iW�}X��q}�9_��>�iC��6`i��8�_��}�{�v�>te���S>�L���.�Z@�.O�*�z��Yǵ3��?M�1~u���-�t�|�Nχ\�g�bG�{r���������5vY��t�G�\�Y�zu���2uC���v`A�:^C��Wd�
vg;�1eW��ok�*�G���n�b���Q�Nzd��ĩR�9T	t��t ���Ny�z�?x�$c�w��C�Y?w�;Z�^�Z�3�a��?,��"�1��v�������U��o�:%��U9�ǈöS6FZ�	G�=�/��n�������({M�{Nf��s�/ɷG��1Q����e��I���P��Ɵ����3�&e�v �|$��%{����MY�9]0Dl��F@�UCY~*�!��z�V{�d/[*/��ȱ���b�˘�nS<����m�ZW\�>�&����<��ݎjϝ&��z�ݛzÓ��W�"`A�f�B��&vbbt�m�/��)K�]��rw�� �^1��ܨ�Y���y��ƔrHFv�ǳ��Q�����Y��T
��poiF}P�D��tz˻M_V�E(V�]�j�NEƂ�����5j��Rz�b��4�*�0FE�3�9-�\�O3̎
��*)��^P�R��4z�d�u.+�z�}M�=�U-�.�ߧή��1�5�����^��-p3��S�]�������?m��\f}�0>[�b���B�NL1]>�ۋ��A�)����/�\w�[��-~�ͥDP�U�R��[t(5�h�`��(Ow{���=�\b���w]�b��r��n��C.�h�k|�c��vn��,e/���cظ_1g�q'��W�з�Ҩt�M�)��Ə�w4��|�5� n��h*4Ke�_�\���x�G���!,��p��7������C��١cy��j�b:��p'G�Vt�u��X��^����
�I�n�zu%C�u!ʶ���F��r��]����ð�X]��A�t:�ނZ��G�si3�5�QL�/���M޵��7W1g��ۖ7㩟Txg�i��0�y̴LF:��Fx���6������3����iQp���6t�]sft��{��K>�^�3��Y^�.�
��r�u��_HQ�N�-'���P�5FS��u����n��e+���d>{�d�Mcؽ�Hx(��}��R�8]G������y���r����!��#%�Gc/�"|�D\�;2�`�;�kn{��^>:t"����^A��w>8�3���|�m��Z�5��_�ۨ`0�G�t�X�f�~����(+�
.���Z�G�!������"�8o����E��	�����k�,�E�c���N�;-�����`��oC��
ݥ��
�1Z�96y`��L�h�]ٕ��B��k}���f���3����,� @�cOS�m��׶�}/��Ւ�:�f��0�(��U�B���o��P�g�%���OR��r�|xj'�'�w?��{U��ޗٞ��Z���h�a����
��Xb�P���\��󼟖�O�������Y�1[~Ҷ� B�ŝUj�yU/���5�����W8tϺ���	ى��]���c�im^j�<G�W�Lq��ih�Zn"k>V|~�����s���z�~�Q�����9�����������C��銹Fϫ�!�M�N��a��}��Q,�V��ω�ɶ��U�)D�T���:D��y/"ف<�!�;�+���(L]�>���v���쩄1Hav��K�|]�����_Q��ֈ��8]vAWJI7{t,��x\4�5���GG��[.�}���΀���a]I�H�7xZ��w߾�@m.��׿p���lЭ~`R�t-�u.�}O�~�%�>V���T�*�,�FL?NH�ӤC�[�����s��^k�å�a���_�����.�����#2�`LL��7��@���"}ʏm	���?q�l$=�s�y�_RZ~�|G�F#ӆ/8n��Ӑ�(;�952�e�C���B|:�U����Rf#f�a'�OMC��밄�Y?p�QY�W�Na�]0ל#�׸���qeb|�{&`ı��<*4�!�AF��ݐ�HiuJ���9.PG!�É��;0vʓ>��P&�Miý-���u<|��
��!AO�bo�l��{���˶��S��d���?
r���[�Y{�f��qci�����ݑtU�ܻ��k8�צ�ʹLX'r�:�-ޣ��Cz�Z��`��.�*J���=��и{*���/(U�ι��v��F��\�6&`ڱ/��V��yY��y��+F�b��t�E6�L��t��|oC�v��՛�jt��#�!�Vǹ\�kz�J�L��r�l;�k��pʐ|l�yoŊ������+���HҖ�^A�s�D\9�Bn��==t��X%��N�:��nu�����
@�wU8�grN����ǖ����)C�ZTs+q7�Ho^qI����I�n[.����LD��&��_,Ir��=�(>���!j�b��<F�jaZH*��$܃KR�tH�?T��,�����vn��˸�����ꭄ�*�n��{��쇽�4�w�l��b�޴�v�ƴp�r.�9v��X�f�ǷQ͒3���_���3��m��m�z[����,���N��c�0����'o�i����ZM./;�ܼW�ዬ�6����j�؛���㐍�gm�ȶgc��u��b��j��/XU�_m%;��A�2Z�nH���E�]ԳWIi�XS���t�dV8��#�
�n�6+��r!��s��L��GMqam]`rӄV�3�L*-Ǎ�|�k�f!8n"i�T>�}��$F��Q�8�k�n��mA���j��F�A��l�,�2�{{O������]$w�	Nխ)=��7m(�yx�	wN��B��mؗ��R��1>���2�c�x���sI�v6�=�Bneʤɓ[����>�v�.�ۍ�n�m��x�k�w��~�{���2h8�Aբ+�1Qg�Ċe*������1�j#�����L`��v�iX��Ab#L�U�
�jQ
2�QV
c3�Y��Q4�9h*���r�b�r�Z��l֨����x�-TEb*��T��1*8���Tb��(�����c��+`�����%YƸ�AB���A"�TBڱ�lb�dEXi����<�̖V�5B��1m�+�
]2��>�g���WNac�ƬQTETĤUV�浙љ�MeM�(�T)B������a�x�y�h(�Z;h��ynZ��U5J�����et��1�nn��ޟs�u�T�q��3h�Y��;/���k[\l�5����əH���I��)�@�i�~���T�=)�@����ޯ�� ����C{�|��\B�B�k◍����\=�����Q�B���}}����#dOҦ9��S�ǟ�z�{�у����o>�hO-��f]�M/�w���,TS��[c󳺀��m����%��U[����Hq\��r�c�ب��|��t���#��8�I��)��^+��)�&`p�lȇ�nK�
�|�Xyb�̟9����o�������\�SS)�l��~�[�f����,W��b��O���A���3�mN�e��}]�s ���>����ρ�n+�t�H��!���0�v���Y�����yk�@i1�ӄ�����$����aA�a�K+uٽ�¶����	ޑF�q	6cP��z��x�2�X�c�]����i�я�i樺\Ś�)5�s�c��u�f%�k����ޮ1c-������
�n����\��ܺ:��z�G���(��*�ӺX>�L������i	����VDn��O��c'�3���[/i�_LWR��"��T~2h`�;�f����C�>��y0�z;9kƌ���n&yv�[S%�{��^����Y�+�Y�A�������Q������^��/'_ӑ0����TT`���D�*���-�W�a���3*�k��,��r��ځ���uϺO^�k|�,���ʵt�ύ��c�$W���.�
��r��r��93ߪ��y�S��¥���Y��h���)��t�z.�,�����9�G�S�>����߶���8i�5��������M�����_�T��s�t�p�r��T�������݄�5�N���3�B��I���a��7h���rg{�2��C�z"#�h@��<+�P��&\L�F�ݔ'����d�D�U��'���.��'�O�q�Ӡ�Vi���S9�8���;�e��S��/��8��ͿEȨ��4I8��o�ϕn������E�
B^֪��STH5N�ȨS�@��1��:|\_�F��N��v����È�j�Y71A�zW�y_���4B�D$uL��%Ә䚙Bk�N��T���U3��r���(�_!�U7�>"��U���綧��������Y�gT	�y=�~�q�q=�s��ndM
�m��sV����9q��A,��?\\&ml7/�2���k�zY��m�R�@leL����ʺ̝)?)���i�%x����,��J�
k�M�F䔯e]�.S:��� WEP�2Uڤ"̣��w��Li�3+�f��B���=�#����T�O�[+"�
�r�rÄ)�죇ME�1��ݫ�5�wz�.O��5��0!{�Y��Þ�i��R��T���?z)^�!,���ي�q2:�ȟ7P��N%����$	�}����)J������ g���2eLGde!����=6OR��C�<Wyѽ\x�܇t� K|�"͖���e,��ŉ��-׺xm��T�Sm\E�w��vJӹ���CG��v���x�6֝�s�:�4�3$��Y���8���X��G�x�0�t�t�};�(<��,�l�kqfb�z`O����2$z���J�#Σ� >a�v�(0�u������L(��@Q�	������~��I��]ׄ�H�5��ʣN*��q�F��ۚn�K����������%����PY҆c������qZ��4���k<����w ]	ͳ@��ۯ��䱗'-����~��ͫ�̧��`�20�,�َ��{{�\_u���������ӏ��6�Cq�E7����l{;:y)��7N��m�=m]J��Hk�:"�|J�t��^�bl�}��VaT����!R�E�3����r��'��<M+94���3MԖ�O��bR�Zp�j�߄��f{b�+��!y44�tFӱ"&�Pz���ـŹɁ0�l�#l�
X�F/)�k����.��ט�)��L��u�dI��f:��Mg	�h75k����
��NN�����;"`ɘ!Nt���Z����g�H4ϡ�(yq1��m}�i�H���������`�-��II����� ��UUӏE�q\�J5�Uq����^�<�T�FJdm�.b�]��V�JG�c9���v�ax�^���G���e�U_|��N�����+6mغv���O?5Y��o�&�����R<���}Hǅ��?��������¯H#�8pܿVL�ʛ��y��
�4@A#�'1ƹ}RE趞
����0��{����$�s�9H$2��- ��۝�ؙ�ťcj"�J�DU��2z"k�L�H�6�5F	�M�mLT���W���7O����%Jf|z�\,��a�l����5t�l��=b��_Z���*b��Æ$�1�t(3F�����S�%㼨�Լp��!�Įf�NN�*�e�qsB��˘STWm�*�C�O�t�7F\�W��E�Uk��k��y36>?q�4���HL�!�ٺ/���_@�fT ��K��;76F'���;z�TL3ۓ�g,	�v��:r�xR�R�۶���9V�9�K�s}�u���q����W<��d 
����d�Щ
�: ��7vsc�5@!gӵ�񺺿{�\G�+E)��A�b�Y]�]K7��%����{37K#�K��CZq���E��:����w1V�3!7���)���1�nbza��W��'.��JD�bK��m�M�gYf��(���q2]��H�5Q��s�9c0p=8řS�bs���<|t�:E�_1�����D��߽��v;1ٜ��~ӹ�g|�z
Ц��5spS�R[��@9u��yu*��u��Ʌ0�D����	]O�j�x�GI�(>�5�|~���t<�i_B8�%�M荫�6�`�F�W�S�l�U\����o��D��Ƣ{5��*��j�4G��u��vP�H<��X�iҮ�>���pQ(%&bɂ�@b��{n��:o�|z���3&[UY�5�}�K�LٚP��B��w%�͡�dvһBۗ��� ! 7�����ٽ������a�6�!�U7�>7���K�������%4^�񜞡�Q�VF����n��t7�U�*�g\-�.��|�jҟ�p霸��4AB�C~�]Ϳk�v����W��3�r�~B�ij��-�)X}X�?nZ���{3ѶI�/�l�
���b�f�ܻ�)'���箅��(�T|�X�q���Nʆ/�LnÎ��?�!�<�iQj�������Jݡ���n�rw��w �j�_�Fڍ�*
��p��N�����{���S-]J�u��Ɣ�STI���q2]Gps8��f�t��$��m.��2�zT�CU���#b`�G`9�f���{!6����z�S1*�kJ�ȥG7N7z�K�O
�6GWS�V$�wWˬ�7YL�����qX 
BA��s��~��x�������{�R�0�֝�s�R�,��9+����źs�U��\�����fјS����h�"$>|��>ph�ϝ�"��`���oN�AtW#��x��81��\t��rMs�	��ؚ�&b2FeĹikudm7Pm�τ���´栱Y��0�I�u̧�^�ov"z��>;���tv'���q��m���"�P�]Fؘ�4�^L:�n^�
��!]yDT}��]�
w(*���"��h�*0���ƅ�'1(./��LZ�y��Bש&{������ώ���|0�!�&�k��Fzݩ4#]I�W ǵ�l�1ǈU�Yn?�\cBÎ�{�����{����j��d��cJ[D�HU���T�r��Q��P�t���͙�7K�3�#��D̬��N��9N�9.J;����H)�sS�w##x���'�$RY ) ��@RE �, �(��Eb2���;�Vں�Ŋ���E��u�R���U�j�NO�O\��"�be��� c�>����}]&`ͺ�$�L��Wo�͋�3'8�E�~��~U�ϯꎍ�u��I"�Q�*B�"`�s���W�V�#%�����LM;�˘rf9���zkäV�b�ٝz������p�~�����9���ԯ+U|��Z�G���pѤ=V����O�xQ��y�����,����=����j�����|�"�e|v��S�Lj�`���s�����K�wuF����\�E��^��Z���~����HA���!�Vt��"�e��[��m2�O����d����i;��F'�q�����?Lz=�~g��X�M,Ȳ�<��e��sq�T�t^���u��Bĝb9C*s;[���Ss�ue7]��C(
�/y�ޛ�O����]�ZR�_hRC�`�-S��.��������P꒓�X��k5US�i��9`/������q����Mf�ɦ��3c\�Z�t2�r#U��A�������M���/������7l�ʯ1C��C�Dy���3��v�A��m
����B!��n58��Mu.�f�;#Z�]Y@�8�ۺ���$�}��1)�V�uZ�����;�eFl�aw�1u��h�G]M�Wn��/��[��k��ͽ9v���9ͥ���ij���ɨ��(���aV�*��7��z�$�v^$�g:gu�ف\�� I
����hХwu�d(x�]V�e])��0�ʌIۣ[�W��37G�8F�V��Gֹ%k�V�%k�*�n���Xv���N̘��v�=YT' /�P��"7T���!�$ϲ��~�QđN�UA��k�5��V����$�\<s��*xj�k�/h;��~{p������.K�%� SM�RWC�I�	e�9�f�j-{�.Iv��"��L�ǎ1��v�W����N#�)=Δ��-��"U���_��@]S�m�h�� �,�]zz��I�p4�aq�9]xT����|�n�C��7��f��C�ޣ��L-��X���b��d��:������g�j��r�8.�C�vÃ�F���*n=&�ht'MM��{��]��D�m�0=�G��hPM��mvs�#u�aUd�qJ�;��Fs,uX9{+��r�V�
T���+��[n�Hԉ�M�y�R��R�K�*۵�!��X/�H�p�KQWȥ������|�UTD8�m�_殓Qg�/������TE�������uj���j*el��PSt�(���Eb�"�U���]Z���)r����ˬ��*�Ƃ��Ac4�A����*r�����F*	�
,�Т��*�*+R�Eb**�QQTm�r����ә*��D3Y�ET�y�*��Q�"��TUGv�*F�UL���1Kh�JTb��0QV,�+�V �Tեh0R���m��QAX���Vq���T�V"�����\�TF+�b�g3�Q�る���O.�"*�(��ģUf��U{i��(�:��j�Z�WM�>Z��2���Pw�I!�5�w������c,t�����6en�g�6jut�{��!%H����d����G��
�| ~�_G�(p��V;;�5���4��c�,Z���s5`�fT_��a�~\����p���ӣ����ݧ<��0��KX 
�3�^�^p�ʘS
c��gj���e�<#L^����㇍Z�=��;�:�#���?I�<����_y�x���W����ڧP�Ad���βc�� ��2b�s�$Mv�Cԗ�C���|¡ԗ�+"ͲVq<����3�������ϒ�AH,� �l
�h-f�*Ag��v�'�
,��R�$�1�a����q��/��+4�S�c�w�~�ټ��o���I����Xz²~eM�V|ɭk QVϙ*A~C̰^0+3�gi
�_M�L�y@Qg��c����$�7�����k�y����T����c>Ob�P�P<JÉ�1 �8��)+����ϙ+:�b�?0�1 �8�^0+<���\Ø���c��>�P����<��>�J�� ����4�A}g�Rk�N�I=�PĂϐSC�
)/(x��
2����0�{�H)-�d�
(������ｹ�/������`�ԕ�&���q�C�/�7�g+<���QH)<=�����+�a����]���Rk(b�R����;��P��ْ'<3�\����p����޺�wX"}��Gf�b��6�.��RGS�@޼�!��Y9R��ԗi���#;t�$����b����G��r-�=��l�f0�H(>���:�Y6�Rm
�2o
AI�B�uϰq�a����g�=L@UR���_SL���Xz�����w�s���7�z���*J�ɼ�(�0+���Ԛ��a���n |��OXb{��@�+�
�Y<?Y��RVaܤu���|�>����~��k�=@Qf�*A@�?S�
�\AaS���Ɍ������H����J�A}�`g�O��=�I����X��v���~���w���)8�H)�����XbAd���|�PXz¤y�LCI+�6�V���5�!Y�������(�q��?5#w����׼��y�q�
È}��$���m����{�1 �I�c0�2����2��HVi��'P�ο�1��Vk�w������9�s�����
�g�d��bAH.w�YHT8�a��*O�Vc'r���H,�1�P���Ì+'��JΧ�/3��|����}����P:�?�l4�X~a_���1��H,����2b�<��I���]���
�'��aS�����|�^3�E ��3����|���\;����۶J�����ya�P���=��M{f$�
�ݤ�>Cg,���~��x�P5��a� ���z������{���|�'�:¡�K�!Y��M3l*~���kYL�H/�
î��
�X��q�����P8��T��N�Oz¤/��eϾ�����o�u���+6¢��Vi6�
M��1Ӵa��O��rɈ
*�HT�������+����B��%f2}�D����P-���hy�H�u�{uj�%���]�:ŌM��Yǘj�������خ��!�if��uԵ�l���ζ�jܘ�H��FV,޼��������%jNy��R���
Av�nɥa�
���Y�x�
%a�
�Y�Lv�%a��!��Ϙ}�i�d�"d�c���1����,�G�F�{�1��1�N�~7t�Y�J��
��Ǭ�Mn�}`^Xs�H)7���H,4¤�
��*Az��Bg�ٻ���߿_�R��C�&v��I��2{�I�;�'�'��'Y:���:08�m� pw��h�����}��s1��2�=1���bAt����xÌ*���O�Y�O'��
M�Y���H)5~��_�1���4�S�
�O�1 �7��{~?:����%B���7t°��*~@��N�IR&��Β
C^�u�0���Y����<H(?{���
�L>���=����{��{��.ؤ��r�0�Ag��!����(��J�Z���v�$�aS�sT4�YĚ-�l
�SA��TP��L}`_�:�o?n��w������AHr��*Ag>�b�V�
A�&��0�������E�XT�eH(x����8µ�$�R�.����<�<�����'2��嘐X����g�����S:}f$&��R��<f�q�a�+'YY�2�AI����9��ץ��{�߯��|�Y�mz���8��1 �̚��ed��f@R
I^�+ԋ+���8v� �L��AH,6��$O_�o�w����?O��*��� �m+���4�P1*u�~�1 �b��AaR<�rM3*N!Y�J��Ԃ�@�U��=C��禍���g����ф�U�j�rP�u�T�v�w��qǘ��T�x���f��%ԥϸ�kq[�6�s��﷓�-��]i���iU�3)��Dx)ۏ	�Dϔ�_̕���풢���1�X{�~g�E�Ae@S�H)>B��l��^��>��0�J�YY+白����~}����Ϥ����C�i1 ��4!��P�m%���4��*}hm%H,��$����|�Ԃ���a�cr�E �:�����Ͻ����i ��&٦aY�vLd���f��4����И�*Ap�Y
��? b��bC����g*�w��/�".~�DT���C�ϔ\o�2����9��<ayd�R+'��� ��S�N��X{�~@���Ă������YXbc�*OPĂ�yt�� ������y�ϼ��`c=d�q
�?2VN���&�}`VaS���*AgS�1�%E��*Az�S��_�'��Aaܰ�q���{�������s�~��hW�R�Ϭ�0�
�hT��$�ˤ�W\�1 ����ӶaԬP�L`o��m���*v��
�Xs�/�>�5����}��mH.$�Vi�Z���0��0�c<��H,<g
���I>f0�
�?X��+;�& (����+�I���{��Ͼ����ι�w�~���>IY�%d���U�� ������u��n�I�a�~�E!�� |Ԃ�����U�_P�A@������<�~���u�'Xb���OL:¡��LH/X��CL8°4�z�Y�J��&"ϙ*
E ��<՚x��<a�S�
�SOY1���Ù�)�޼�|���~�R�O��
A~`]o������{�&3�T��LE ��i1 �ч�c0�xj�6��iE�P��R
y��ۡv��T*z��z���=��e)��Z΅W�R�Zr����[1$��X=V�G�ǣ���ɞ�j�U���IX�ݗ��1�&��`��{[EC���������;��i??0*Ϯ�i�/�OO,�6�Y�
���R
k���i �CϬ4���x� ��8��E ����M$�ԝf0��9�s}�>����N��v�2iE>B�+'��8�?2~tÌ*AO���|�Xy�b*�Y0���R9��a���H,���=;���]޷��}���{�E�`|Ԃ�Z�U��M��AI�ө�~OXb���X|»�`bA~f��M0�
��Y��%gRyn (���7{���~�_�s�y�?���S���>�+'ᘞ�T���4�_Y*,�%H/�k ��gi��'�i ����u����PĂ�����}����ϻ�{���qa��,H,۫I�
,7O;n^������ɓw��C��S{{������%��1�b����iޠ%Ց��,\d���vn���3g��_A�O�Usu�C>�K�.*x����'�Ԝ<p���^��+�7JzaOL\�u옚��#=���o+~ʃy^��Y蔫�{�xpgL�>:h�"�K��S��A��$��Ade�O���YZ���s�9_��tΔh]q�O0�s�k�p��z�Wd���WV��E�+{S8<�*�v^��*���v�vՆ�y��u��|�in�,tN9φ��d�C6Ɗ3�[wF�_�{��z;��d҆
�"M���t���K�B���K�Y����XWj�q�bhc~󘰄s�@�G�,>�9�&�P�Ke3ҶD�S����(�e�(��u%�˃ݞ�ȼE:&~����~>3-�ψ����Ӡ�GTNߤXN�-�y&���u!ӑ1�{� +��[~�����>�X��e$m|�qq`���K����������������_�Tt쉨�"fs���O�f�W��[�u9͜���E�g�����#�9v��N�>��8�O���'		E���^Ė{&Ѩw��D2�����t�L���ØvP�r��g��3{����Ͻ��J����nszd]��V�\�huݹs,^Sޓr>�%�F���Z�� ����%��'cc���ɑ����¯�����G�ir=�S����u"&�:���e�ڸ2f�\�R����즶}G��To�����ƭ�
��JYD�οk�U�=�F�v|B<C0�MEm^�BlT_���oj���{A�b�fbd�ӵe3��f��sN����X4g�+˪2Z�;�~�ً���=P��ٝJ�a	�{��ęw�αLx���"�9W����`��(�����a=�.w�����5�g��Q�U
`�8�JxTb�.��N<�j���ova��|��q}�5_su2�Q}�5�aa���f�?��{�:ZFӳ.}�'�7}��U�����To�;a���??�i�S�>#���G185VF��Dļ|}���:ТTT��F�u5�#�˅�rv�Յ!�6����T�}H^��Z���Z��\N4S��}_}_4�NuJ;o �Š��q-i-ag�+�lC��7wo��?���$ӆ�\�n�AN�Pw�}��7֝��Ѫ���Y�`Y��w<�
Ʋ~���;�&��H�6�ⓤ���ȼΉ����ܣ��j�U�B��/�~�w��
��P�/��"yC��A�p!C���菶TiY|���}z	�4�Ч����;4c��ƭ<ĥ����rU�,�G����fr¹}U�/�y�ձ�dY��Ԏ��M�bܼ�SW�\	S�㦲��Wnjc��O
x@Q���ܹ�=�5�<F�vG��Z�v�ˡ��Ug^.�l�����X���D�@�b��W�\�p���gt�����[�iyVKM5�1Qx��U��7-Y���8�C6�ư��"��;�iҬ���g��eA�EgkF�gM ���r��O��G��I%�/�ȑ0�tm{F�*��*REy���ř�YZ�ro����i��h|3�}�w��35�M=O�L輸�D��\0,���.`ĉ�l�x�����|C�w��~;�ۺ�<��o�,v�P�����־�E��}+�|�Z�۪/soj,vp+�gg���j&��VD��������6��r�!�L`QF
Zs�zF��$�x,ɐ��H�%��%c�]WLX������3ŏ!�VKN�7ɧ�_z�6��6G*�$���6|��]�b�p,����g�pӶ��8��Y����u�s��X�1]�AA��-���º����J�(K�S9�.\��=G��Do����x�^1j��9�s���h5�����}�.b��۩R[�;s��UZ�+�JV�㩸;Sb`����6n��ѫ���TI3� �Tr'.���]<9���R��^��"r�^�+<�PJ��nkcMZ�}I��m	�^f��\����z`�u8��lGJ��L��w1�/�^�Q�hw�+��� ��^ͅ�Z���i�@��t����[�V t�U⁴OM*y$Q�,��󲍜K���~ӕ������!�;;�w���)!J���2�[�t���r:-g�Tx'��9+���P�z����?<�a�
�ǕCE '�����]�'��n.c'�)s��O*S*\�*&:.3�hP���X|����t��Jo£f!H��.\�~�ͭi�Di�R> �/�-.!��2����2:�W��VMK,	��fi|2�%�Z��	#��Fľ�PP潲.��D�b4:5653��-M�&�S����=_V�q,�����i��MUoT%+�W݁�E֞ZBB���i��UR�[5�-j����R"Ş��M��9�c�`	��#2[l˚�z���D*>kr��6� 8i��Y�|	霆Jo�"ku�u��R
�HtW�Bh��t�s(Ao�Q�C�kz�iwyq��M��DSK\�Y��[�0��6��^[���f�Ő���ܫ�w.�E��j/F)���*�Eb�Ǽ���\V���jQs9��)NXy2��Y;R�79_^F6���}T��W��xk��r���[Ûbe6f���?@E��%�J�c�+ak���9�E���|�13,��+۔�A�e�4�1,{�ϲ����G�y���ͨ9-]�(�ea��ę�kt��m1�9�K�����(M���7��wV����;{��g�Wb���m��[y��|��Ѻ�Ĳ��]���k��o ��ST�A���;fauS:Z|��l�Av�6͋�0����nNE Y���ǡ�n�n��6�L�S��H`:�i�}yp�w�2u;b��f�\[I��E.�ֲ�v�uy.f�t.�1Y��t6�:I>L��R[��۩�J���S$��c1i)��w,λ]���U3Hd�ȧ�{��B��+1u&�v�������K��su��b�zh�sqb��2gL���������DZ�J^|h��9T��3n���z�|��<�c+j��ַS�U�����Z#O���H].S���]��uV�]|�;��F+�t�Yu�	|sFT���w�ʃ��TrWpe��8����um ����`����e���&�^+-4
8���7��}UNk1�����Y�3�,?3�ar���b��5���EF'P�+1���DR����֖�Qݘj�,��n#�UST�8��ҋ3ª��[y�Es�kKk���+��Z#;�0]�x�EPWƊ�J�Ȗ�X���,ZE[Jr��y��[�����E�Z��"�""�jɞ�I`�ax�,�Q�`�F(��ƌQ�f6՞һ�8*�/�1��:�*�i�q��>%�M:��*�,��ch�[h��Kj��J��Qc�ۦ�4M%,)�@H%�Ι�BV�#���>����=t�e�2.���[dS���ή��2W������	�HbLM�n�;�"�1����ME������u�vѩ�Z&O��&�� �?�:B�DTpܑ{5$@�u�4��T��L�~_��b��A��n�
۵�{���1Ib��p�O*�!�s�%��*_�������_cЋy���0&�=�d���Cn�ג�2f���&޸P'�]�M��a	C���|�"�\C�3ku{νY��ÅR�f����0��
��}�v$��(Y�W��S�m\�k�Y�2&�4X�q�����ܗ�龛�a�����x��B8\_&����uLMw4�gݕ
zy���B������@�O>��ڠ�p���������;��0�Bwf��4����b�i�W��Z��_%Q�����Ǚ�����vnE��J}�W9�ጅڌt�����DA�<Ч鄲���@.���
6Fr��k��r[��oi�k���\]Qꌺ����lH�rr��LdJT���R��*����/ܮ!�F@�)#����!�0�kN�"��P�����ȋ30�i����1Q1�����)ի��l�/-+��mש}�掿�o\�߸ľ�n3�SY߸[u�����i�,�b��+��"��i��Wj��X��q�g��1������8C��R����>�qeݗw������vu���b��4<�#f�Ş����a�8;�Z��q����ۯ�R��7h!�금di0�w��C�����וͫ������b��#��C�3�1ݗQ��3#mD��P�>�T�%��J�.1�'^i�n'���	.WE�Ժ�E��r.�ad��9�L��J�Hn�:����X�X���*㷔h������e�;h!��c��S?n\�a}3�n�qmx�wM���3�8����2���[��c�X���9K��X� dGB6�-��*ߝTa^Y���+�^.]^�=G�{KRlqTbr|'p\<V$O�W�����!�J�z݃�2zg���n!��9��
C|��Rآ�Y����څ�Փt�fKq���Nz`_�I�yItg�ss�������Iq_��y��־��=3���±Q�?ZXY�V�T�����Y�zB#j��w��Q�|~����~�z6�&;��hpW���	�FpF_K��~�n�Q=�VD���Z�ڪ�̵� �GUG�<t�@�
.;�xFόUK�+��Y΅k�����D.�����/z�s��V�I�6�kG+�4��><l��&�TXzn�^B�F�t��7�����il>�37��p�	b��ì��m��)�����{�!߼�y̽}u����5-�mR������*B%C�G��_X��k�n9:T�D�h�#_?��y�b�WW0z��_��#�;���׺��잜�����}0#��>d�����boj:D��P�g!B����,<�M��ޅ�
�vT�l��RgY�I�c�*aL)�:9�J�oK;��C:��Μ4x����ߩ��7JzaOLM���=��r�^(��/���"�ssʼ�����b�b�w�7U}�Q�<��8DK�4��?��k�/��b�7j���:�����6��<u�g�}wl:�'�>�#ϲ�߾c�����?��f�D^+��f��`6�pu�{�*�e�+�#�nX�zVڢ�-�\����	hK1 ���R4�8�C�Z;�������� �owM���Dz8^˟d���ԙR'g��EmLꈹ���o)o��6�I\���������秌�xo��J\�19�,���m8�r2.�3��E��PU)"���|��YӞ��	�����!�i�I�ʵ�FYC;��t�YU+�ޤGj�z��/W�El��/�9��������>���L�s��dx���o 4�0��S����޽�6�5�*GQ���L�5�	g�I����$:�-Ŝ��D����Q�����0�0��jG5i�X������.�����?�70%���Nè��W�cK��}�=ZUU��K�S��t�8{��vb��YWrk�.vc�/��&]F�7���{=��܋����w�8��j4:����I�w���Wլ�:+p��Ut��YY}�WfŶ���-t ������'�$�����AIZ+��ZC�E1����������+��|����ۇ�"�~N�~0b4$��{�s��yC��/Շ�?�c|pȾTM������Ƹ��!Q��G����{@�f�n�������Ǥ�C��P�S��
!���C�Q��W���k��1s��/�y����a,�'�0�=�R�_Y���͒�;ԋž�4��>�Υ��+W5�Դ�+^�&wg���k������dx!����;P�3zm I���>f��N�v�:q>�uM	tn������I��^6�|�^����Z|`��4�i�\~�_-&�-繱+��n\��6������y7���`���=�.�q�5��0)g/�=���׵�h&ƪ1�5&\�0�!b7q�D̤	����r-�J����tj��Ͼ���m�oi���L�<Z��Ϟ�L��5z'����*U��P�1���g���!L�P�`�t�d5�<D0��@8��NNG>��1:�0v�]K��ʘ��5�1Y�Z�ƈ�<ę��{�ڭ�J`�#�Y�v��=��5aO_�~r<�_FuÞX�Qad,�ɏ(T'�+ԕ�g���+M�Mex��-����84�T���tC�xf!ǈ�TY��n�1���Z-��7d'F��Ê���^]5f��)���
�
ޭ�qL��T�ӧ��t#|���I���v�r�8q�hd4�/h�0����疜ϭ��O�+�9�*�P{��|2�0q#{�Z��Բ]c��/��G��y�e��h�o��r�V`;UO��3ux�_O�W���V�{Q��Nd+7�e]�[י[E?�W�$��9Cu����+`�}�i�8,8h���,��%z�w�	���1q��b�W�y��:TK�^��wv�MA�86�y87�1mκs2;<W/�{�l��]giҩS���.C�U�8��Fȇ�z�0���$	�Vd8|9c�^�K�q}^ʥ1~wX�mWvB*����"�X�%���b��,9_a�p��f����?���7������᷿^�83�G6dXg��ͪT��M���Ϩ���U�/�U�T�Y��1�X%�Ȩ�+T�9>�{}^�e���!�L�k���=
�Le>C[Ke����}�iv�_l*�5��n���� ����tj��UߖtF�I���w���&��7Z
�K�u�N��4�;I���(?��n�������U���P�t��C@�ud�EY f���K��D t�+"��>ꏏЇ��D0��%,� ,f02�����<��1�'6���"D�z*���Ĭ�!߫�LVR'pJ)��iBw�]KWK��b�V����W�T�^4�/z�N���#U����!��Y5�*�!Ȇ�>9i"%�{�|�#�kR�=>��~�D�.�Eע�Q0��� C��B�ٔ��Tl�O\;2�u	�Ԉ)q>�ޕ}��|��4p�������B��:�t�KBOG��y���5���7�ܽ�O2����<�r�U7�}ު|�F���4�_e���8cK���.�������w�Q����P����4�*y��a�RP�X=M�hؾg<Vn��[�*ܗk8�o"��~����s+�ˠyZ	��<-zt;Z��2V��i��WU�6�Yw}�e=͔WܣΒ�66I�8Eu3���{���S=99$ј�R�3(Mx%~��j/��Ś��>M<�ɩ��1�~��1T��N`�s%��L�-��{��:�g���q�Y���d����;q���:_���w��p���L`Q%�07'�x���s�L���w_�{����+ʊc�N@��Vx�k��GbDRu��3�{}}�������;�Zl��,�Iң~3�Mq�8����ʗ.T��Z+ܫ�|.6mН��lV�tLc`]�m&����\����L�s�2��u��>w�Em?��2�x�_�/���P�l{���4G�(�A�����|(߼a}��W�W�\�F�A-��F��<s|��>���p��������e�h��{k8����]��� ��ݓ�Z%�3�&�f\8yu���&�ՒJ;�8A5$�t^X!��1[�i1ܮ�./��\��W\�|�(d�n]�Q�������"�n4�-�s�uz˶��d��5�Z���]˲�M���6���xR�t�Xr�)����!7K~c-���is�s�,��W��C�8�kG�d$�	ԡ�C[B]v�ˬDe�:9��b�*��:9P��Ǩ���zR[{��*���Ѧ��l3K����i�}�L����m��W-��7Z�=�T���w�ov�F_s�CK�!�����x
-l��p�� ���+��.�u\��"���ۧK��\��l��)>r�k2\Z{�>�R�*k,?��e	�өr0 D��r��]{\N2�����t�ΙF��1��8P:�BM��m��O/f�0R�չyEq�lb��r�qfL��k��25��S2���t�>\���!'
�r�Wc�7i�Lvݤ�Ȩ$�:�Awl;�r;�Gq��R$�Yb���5�\s\����EX�khx��:��ގ������ʉ���e�G��q.ߊ��5�l�ҭh��s>��"�ӵܮE]�v�7;^4y��y��rC�7|�o���WokZel��VA`<�9Z8�<4ܽJv*ى�]ac�pVns"� �lJf��0Z�+Ī=�}����'�/:�Y��N���\�7�gZx���Ly�uI%�Mh�
�i>ڽ�mGS����S/k/���x��F��0O^�O+�.��w]+j䚌̎����m����:u��M=�uwL������֚��>Jإ�a�,V�Q]R�k+TV[,���C��ۈcUm)���QFDL��LLpH�1��a�U\�����*Q�-�s,����3<ȵ��T�0U[e/�'��k7J�N!\�T��b���bǔ�ҡ�j���dְ幫�)h>����y�f����Eq��1L���}���5�Ĭ�kE�.Y��]{�����GM�i\��kd1�r��]*Q--��p����UX�.c�(�����];��k�N;ܴ�8�$m�b���K���Y���֮��(=�yEw��F�#��<��H43�ǯk$�؞�i���/�&�)�#�F���>ci��c��C4m�w����~�`w�cMl�I�3�I�{�O���eVK��;��H�F��b���_����6�Ei��g��K�Wj��˘g��{CY�b\]@�>�ܨ��:5Tτ�x������,`H��Q;Xi2.kF���?hh8�f��?9��͵h�h�<
5�1[�CHk�%jy
&)�)͋�6��θ�j�/�C���
-9��4���hu
�ٍ�a���Ψ/lD��3B|�xQ��Յj����lW�3_�>�5i��p��v�>�j��}t �c�u��O}q�w%E>���������ٓ~�.���"���%�����o�T������:�M�4���qJ�%A��Y��F�=��#�v�̤Wވ�'	/�~+�^/ȅ�#�׏Ư�k��8�������^�Oٞ�ه�г�UR���ܨ��N
��::��u=�Iڔh�/���飄Y��#����u�X�pw���ɜ�Ow���I㽨=n��3Ӥ��cώ�a���ʏ����rB��!�V��k}���pz�@�3�gb���A8��E��r��Tf60�Leҗ��Edl����'��n/Nצ�gk8MO�ÿ9�0���熫�����!�p7�cr�[f�����m  �iw���.?Y�g�O;��F`��!vvq��j�2�
����̪�31B���Q!W^L�BTj�ςVz��c�X촙�'��:���N��62EY���
ʉI��B��ﳗ��Js{L�q�qĶW.��ht7�b�au�q�Zl�l|�e5z�Mܳ�="�����i����ȇ6�u�n�
��h� b�_}m�{lŕ��\à���.4�_�}maR�8d[9�[88�Y�rY�1N��o[�b��QK!�Bj��S�����0�ܫ�ȳʍ�\h� ��ƻp�v����V��W��*^^ﻹ�Ȅt[�lC�w�Q�}9J{ _���j�V�����;�ۺV��+��)Nͭ��}�͠��Ed9
��+�F8�y�{"zuӞ�>��&;n��I�YP�;�t��#�F=i�,�Y���9�U�>:�ZV�y����n%���R8*���">�YZ���C�W��^0CT���^�U���S��2��H��nr9�z5_� �*����	�g4��+����]@/�hj�Dx���fe��~w��
�X�d,��K9���c����fn�'���DLk�޸^�{ZR�2T]źVZ�ܚ��QZ���3=�=B�D�=?�)�����P�˨�Y.-�����$�]���O�ܙ2�+�����U�l�y-_`"���bwB�u�w��6z��i�^g1���ҭQ×f�F�� �'N��c��Dژ�^���Uǯ�$LWv`�tI�d���"{��^.�<�?�W�����d�zWK�����!�e&s����C�h�ק�t:u�==ם%��\NS�6ϛ�:��~ѷ�wN�=��{�Y�n%ވj͂2���K*��Tȏ�w����Ηe![ζ�x�!G�#�}�
զ�$��1�񂕜U�_F[��(�Ll���!X*.��2�	��-�|{��{eq�3^�=���'-NQ�YU#�zv(0e�����>�����2�o-��\gGE[�,3�(VB�Xz9��=Y+\��n�
���ٞ�����iuw��Δ��3n���g,��77�Fs+��{��p|bg��~ׄ$�uU(�����ECv':���/%a�T|/���/o'�u�&�I�:��8��zS��E!���;��l����x1�wbbQ�z��мC�5�nB{��/k�]9�G^�tq�{�f�����}�������q�9�wJ�9��oC�F�u�RM����i�ˢ`���	�8�9m�1ԊP�����I��Тw�{��>>����!��t/��0�����?��Ąw��/��{8T�쵭q9���g0�;[��:y������j����r���{{��f�K3='�����E�VRi�I�:�!�3k�A���ق�G�<�H�X����8��fuՌ�zp��Է��拾5�;o�:�1��BOR�ඥ�`�[�ن��C5�2�.v�r���cy8��1�v^,A	�l�؀��/X�uf�a��!����=c��FTap���-��f�.��\`�l_
�9�Q��[�X������)��g��v����>U�wo��8��-�".�md����՞[��$�y��������׎ߖ	)�#zv2���I^���;MkX�E�ޭ$�S��(��7�p���[{��)�B��K����Ԏo|B`A�F��1�F�^t�c�9����xi)��4
^���;J�\��\ќ��]�����$�ח��߹I�Ֆd��up�%�M�6
�Qd���F�eX��n�_��x�]DpP)\�(8��x�M��M�N�<>��,�^�\27D$s/�-D�Ѓ�f��^�f�.A��1�5�E��(<�[�#LH9bҢf�T[ࣹ�_XS���q�[;��G]��*�y��b�gB�uzo�U��1�r����Uge�{ev�t����s�Γ�<�Rki�[D��
p�kr*j������ab����Q���mF8a��Իi�C�k�+�FP}Slb*�t�MU���ލ�vc�q���Z��3�~��'I*��(�k�,�=�n�_ʮ��UϢ�+޻=L���x��Jy����.�s2�=�'C�s^6�vW��/�T��g���7��\��G�[��5�n��F���1p{VR����&@KN�b�%VQԷ��=��VU�}�cN�ғ~p'@����/B����J�u�Pfz���m��6*�*�"COC0� �pP��m�3h�I;�⑷X��b�B|MĐ���:Fr,f��sUbɬ�W�R�9o��իU�	"W�Gn:7��{��<}�K���nP�[5T���sG�7��:�I��B��5,���M̢��2r�O]���X0����_Dz7������&���J��L(�K�]�fx�W����)ޛ�z���;s���}}<�x9��rW؈�]�&C��_�;���06�W�����ލ�����楫ٞ���7C�R�j�	�͐��Ͻ1��<ƽ��u;`�ԅ����WҦ�;��O�8�{[��w*0l�k��[:�T�h���^ErdN� ���B��W�.�(����Z�����,:���vjI�W��9�����Tvm�Ef�{�����u���f��X�U��X��=���\�7��4�5w�wb=�'Gp��wENc�6�Oz`[V�{�*K�|gk{%��x����=(̌_��L�̷����_kyZM&�1]��Y�� �߻p��f:��zY�[�Y�=�r!���S-m�ȼ*�n4��&B��>��No_W�TvD�#w-&y����i�C���KPN�f+=�90��=<��	zU��R2'kH�uxf��Hdٽ�z�D�L2$�<���^v�z�=̰0�U��3]�Qzq�����uspOD�ǡ�@^;��bEU���μ
��v!\_��/}+��$�g�Qub�V	]I����b��)����9���c��kQ������ؒ�يsn��N��n�󾬣�M�#{i�A�N�t��J��(�/o7�I|��wfٳY�/R)��L���B����EU�㹁ب��֗��Wyn��i�V�+m��Wo�Å闧*RK�#<
���f�v���JW#{�|{��!D��eZ��ٵF���/�\�R�K�:�U�ٽ-�,�Z�FnI����8%]����<w��*u�c᥎����� K�uh���ﯰ��HI�F+�.�+Js��-�OT��i)�dް�]�Z.`޲r���w[�I!�&��MEw�]4�&����]`��.u;�����Ѹ�v}DWf�+uŮv 4�ks6�GT;7�p�#�}�U�B"o���%�E�����*��|!����nЈ4{>ڮ���IZ䕮I]iB�����o�f�'�^,�j��p���g;V�1�M��Q��Q����6����FY���Wb�V
��G3rD�-I�����t��]Mٔ��X�k~��j]�L��¯�ckb�Oj�f�V�/T;��x����\�W��\���E;��o2�9���if�R��!|���:{շ�E��t���W��*���'_$d�$��]�hQ)�}�K�t�0b��Q����:k��u�j��3���@5Pc<��ܔ�8�`�tr����u\��x�$�v�}t��)L�S�����;D��K�:kD��W+�*v�����u-s z^���[=����<��g ��'}�4���wo��S�ݙ��˪*:��J���A�*�;���z�w.���2PE:�C9w5�k�ݽ��p\]1Ȏ��[��1IY�W��+�xeu�
G�(��+���im��5����'�q�U-�uk�iUp1-��*��V��L��*P`Դ����ܕp��J������k)TDZSi��]]9m�E*e�#�T��u���)��Ab��\���j�!�(���pKk���R�)mua���QZ�{�b�R���PP�TQ���ė�g��-����, �{ˆ�]��M^kd<��s������ct���+�{���ە��+"v3z��ؑUU ʯޏ{�=���?B���p�^�Њ�����e\�8���Ǻ��{DP����|�
�u���|2:p�K0�gu����5�Ƹ�uZ��W��V��f�ct}P�NG^�)�|{2-[�6���މ����kr����5�/����zV�3����ƚq���/(+��1��҅J��n��Ad�E("xbs����h�By$�Q���p�CJH5}��*��s�7��M�`7��]�g�#j���N07v�,�2��m�y�j�8�i�e��gW*��nwQ��+We�BS��K�{9�+���9Hb�Xb@;A�Ί����v�kD��{)V"���^y�J��a���ol[�dnFօO/��d&�:�x�y-����rȘF����l�3��6�����ݸcs6v�WL�%����9�[����|i�`�hТ��9�HzB�ⲹ��XR�-�oL­�]N֊n� �g��Ȓ�WlL�1��%on�l�5����w��7B��w����5�б���}�z�`�.^��=�N4�F�g>ԫdZ'�s�
�X��Dtoa36p���5��[����uG��8f�qN\���w;i^�g)c��;�B�w߃��J�Uln}���5��pm+�k�*_d$l�K�Lu^��w�$���PP�(U�P�g�7-��c;2�LlK��Uq.buL�)��1M糦o�	õ��q���f2�ڔO\sq<3Q�ku0�wy�k���f�.�K3���"��Β�;v{xMZ�IB!��r�"j	������n��y�7���U���*�ڿ�]5�����gG^h�X\I�N^l²[\�̫oD���x*G�j���y��༏��6�P��.��]u�������7W��Qo8�I�Q�5uz*h�͜A2Y������Μ�A�w��V�F��.�K"w�Ov3�k��y�W}�ϾIF�r'�~1��(�2�����Q텆ί�hl��;kఃf`��`�ʡƕ��:z1G�<=�K02�Pb�����XÖ��g�Ό�u٭5EC'_nh�amؑ��n¿=7�f^���;	@B��d��x�oh��0����V"�Bf�ң�V�xC�S3�^xFU�p�vJ3�1�r�-=�+#����^E�k5�0���Q"sN���O.itH75��4/���H�f�H�<BS��
h��rt��:������ĭ�Z�����]j��uB�OZK;F����Q;�Gs�{p:/O>��>����5-+�W����t�b��c���Z'GBd��@#ħ�+�:�kV_�z�"Mb���Eeʜ[��wK^���~�]W~Ŷ��-T��䊒ٳA�pƓƜP��K�!3�=�*V@�i�Oq��ӸI��\"]��P���-n�������D�{�zDja��t�Zop�9���M�V����q�rmb��N�j���o:��S3*�:��h#�)��]ъ��θe\�Iy >���Ok���f'!މ23�.=t���.� �2�8��{s���}3j��q�.���)D̈�ɵ<����vy��\+�ۂ��&H����W\�->�c��4[��٘�)��grơ�n蘕�T��f*���?{� T��y�F�_{�F�F���U^��Ql�e1"
���@��N�;Ԅv��c�3$��&
���gO*ӹ}7���Z�2B���k�b���[H�K
�(��8�u�����Y��DM��%R*m�|6\v̻�v��UU�u2Fo;o=��)%�5�s�z2<�ڐ��Y=@)0��An��p�G<�Z��*�e������nas"5��C��SK�d���G�9"�Ϲx���*b�S�(	�ڲz���p[�[��]�U#�^.�ź.mZ�Y7�ta��|����FJx�� ��٫�8�çc�鹼Xȧ-��7s���������Nºu�U��.#���щ���N�h)��{�iW�ȹ,����-�ۂ�K!��8�,�i���5:ꌃ��`Z���p7��0���m���
�w����.��4��6�X�8\h��w�k2L�o�ɽ�Pa�Q�PH��j�����/6H�`��>�V����!\�b��m˼l�{����Z��)�����[N�x&e{�y9~7�^o�ʉ෨�&U:FS;�����ok����W��}a��k{(�$��e�8��/G�I�����̫nxT�uv�^��NRJ�%����S�zI@���"�w��G��=A,����W�7�
4D�����TP]A ����y�Nj�DX�k,���M�+Gl�=	��S�a�S�����Z��/M�ւ�Wy������߭i�q?L��]�����ǎ����]�Syݷ�6�Nc�O����("'b�4G���݉ށ���Z0La�:Vҳ�����w�I󝧽A
Ö]�g�R+(d�s[�	���hʗ�IYS>�l��w��M�û��Dk�y֡_v1܄�fۮ����Q�|�]��}���A��5/2�n@�n昸�D1[=�[��/34bm��h�7��ܷGZ[D���-�.Msj�#������=Ƥ��X���I$ ����8�O�C�f�����z u��{�A)���X��tKɛ���ȃ�o�
u��[��Uһ��b�s�Ig�����U�LL��8\���iָ)�B��cN�V��V�	��S/o,2�B*�A�z�#�'۞���1��"�`�껌z��H���*����.��*�p*��ס���O9��z5no��R�o�mvMXT�DT�b�3Vn�����w�{׼��P�W��H��Zy��
�Y�FMa��o*x�᫥j��Y�2VN�X��ut��7��7'IWS��j㺳���L�N&�/�y=NN�����7�/m[\2:p�B�4o_�;��5�V��{5��V�a���ֻ�T%cr^�|�\I�i+�]���7oL��(y�(�ӱ�0:���N��w��j+4/0t$�G+$g��]A����m��w�8��h�1(�WV$�'9�2�Y�Hp�2i�0��J;^J�=�12��i뚻�s��� gp��&�5OTk��QH��}�&�7`ě(k�����4�܆��a/��}axS�%U��W����u����w{��V�e[<�_l� V,юgj�2���l^k#H��I�nϢ��g>�fVҰmІ�,D�a��orvYicw`�\z���ȕ��ט++R���NBwK-�֫޴o����s�K}���R��ҝe����spN�͕�A�ȞZ'�ت�GU��kո8�(�=ټp|s'p�pi���U���4c���Q�oy�İ�ʕ����P=) ���+�1��%�O�9�Gr�C��WWt��_7yB�U�{���W:��M:�%�q�(�!����.A>y��5G2n�ܪܙ�ޣ_iM�V]8�;��Uk3d�Ud-!���e4���B?A�nۗ1!��9�}ԫK�ҰE��Y��Hu�2.�S\��)^[�;�EuH��3`���5�"����m��8�$��Ʋ�߈]g5R�0ΒIm�{����K{3��/k�˪�Vx˵To���C\�2��I���1O��2§�SR��X=��Rյ���cV:툆{96��\
bW���9�[�r)���*���{T*��p6�3B���*ӱ��l=�tͽ���J�[#�eR��sYkC��i����qSM������>,jz;ep��ᆄ6-o+��Q�g.齋�L�6XsN����/����4f��[��r�s
�Wz������x49j��2ʻs�F�w/K9g��پ2��;O��=�gup.�&��������Z;g��Wu0ƻfl���xtW����s9�]wTUT�ʕ���:a�F��l<z[Df��M�+4]��U�B����
TY�]y�M�֭z�f
�F����-E#i�+}n,��lc&�|�����-Vb/R��Q5˾P���:��E��`�s1C��;�����ejÏ�⪲*�+#n�"�am��)�]��/��F'�=ʢ���(�=B��WĠ��*v�F0QQj�Zbf[�����䜳N�Q�W�_mP� �3W%VNG�q#2Ş��g)�R��Pt�B-2�%���+z���S�W�M��Y�� W؍煛;$���ې�����M;�;i�g6�
�8%���އ�����΋pW\j
���F��1�4�fU�۶�<���}j��=���f��/�RE�H�d��=�m���Sl(k��d⋄���b��B˃�s_#و~XK	�^��%�*�b�bh=I�k�Gq�#{�d�#h���sT�JpK�~Q�U<F�n
T6�n쎗���BU�!�E�rTwS���M_]�gv�9ڂͼ�(��ہ���iw52f�`JF=�r�M�ic�۝5'W���;5��������wI�&�����7�%}����e���{�2#wٍ&��R���6S�ݸ��p�٫�l��gt�(�ݬ>�p"sf�v��ỢM;N�bb���4�[��O=�3�� @܋pi7�wg5@�W�bx>�l1Gry����߼����0e�,U5�R�W,&�9WO��J�証O�8;�GUhT�C��+�4c�3_dЎ{*�h�x���P(;��ޓ�0F՗,pX�CZ:B����(!A�0v*Y�a.��c�_�����e'i�~ݙ�42kƗV΂�JV�J鲬��i���E����b]���Jr��.�f�Θ&��:vg�~�Bd���}3G��������g\�e��aQM]:�v�Yіj;6�+T,�������_Rs9ӫM�Yt��B�T&����+�_V��To���1���P;b��`��n'b��::�^h�o�#���<�8L>���y�aT��ȝ�w��;��+��b� (��$= ߦ����Ƨ��Vf:���ޕp�(��.A�{���cc��]��.���q��6g�dvV2�Z�T�C���{���)l�6���7�]��E�/R�΢	�=ܓu(��G(�"0����/niͫ��բ�����&V�9���N��X���J�VaޱyEO���<�S�����c6p*ٛq�����K�(
���4p�%��Z�-�C�c$־�mWR�}�(�=�xV���k	C��i��lE�O�p�U��u�#2 p��=yM�q�X����9��(2��>;�8�# �[b���ʫ�+Ֆ�	�RF�d�ō��PBJ�*5]��y.X�oN��wB=[�[��m�zj8�'��Dt+��Ve&��㝰�o�Ko�цP(N���wN��Q%�g�;FJݣW�G\<��r�U䱃�[��ϸX��u5�i�-Z�����v]¯�U��J��PfR?{���+������2R/�0�rJ�@E�7�"��i�=�P��l��^�)Gq8p'�B�y�;`O��;u��Mfmꦫ��4���@ۜ%��Ղ�Lh��2o[
�9����_��;$�����	�ZD^� \��e��;�	�{�v��a�br�����b�P�B3�[�=Ywے
��m.���I��j�^2o�5�93�=3�t���� ���Y�z{Y�oM��\wK��볚�΋c���e"�ȹ,��e
��3-O5<)��ƅ�\��ķ��2=��<J��!Y2��͍�iXj����ED�4���IW��ڵ�ι���;���WP�g##x��Cmч��o���cH$Q�Gu���ȓ}YA�iі���J�s��3�rӨ�ZϤ}�}*0w��-W�pR��ܳ�C��$�m$����Q�vPX���4�Z6%3����B6��Dn�eBM���we��-���;��8��\;"k��whmL��:�o)�1[L�;���M"�m��\-��yk�I3�v,�zɋ�[�Ύ	T��ޘ�y�%>�[�����ZzYS�_{OM^�����>']�c�	��v.�.�h	��[V���8a5Y�/�2c2z��WkI��^[�gT����pN�N���r���%���r��ۖ��������yz��+�)rOܙ�	�3r�U��K�=�:c�޶ԏ��4s�i5��X%>�Q�)K�c/���C䂶cU��N���V��߅�˅��9�Q�r��;!7��&v���XN���S���pa8��@�V՛���;5����WƺbE'�nBЯc�oY�7N�u��SLSg���F���ۡX�z�]GܫzR=;R�����ܮ��jZ/D�Wo����'5ڍ[	��nH=��݋m�N^Y�w(E���y��/աi�GX���o�	c�v�]�pj��e]� ��Ð�z��H63�z�5K
��u�1\����uc�ښ���N��غA�Հ���6�B?@�����pPD�K��n4ʶ_f@ա&9F���HJ���I�����ד[����(8<BC[�F.��>�k��Fn���`���z�'@)YD<�ٴ)����^o�_�'�.��{�ĪO���LRya��h�嬍�()�������'���gOq�e���O�C�o�;/�`O�q���[O��ΚWJ@�w?m��xtm˓���\��+�4�t�Y�����B/+7VEU��2;�i�J7n���YH��F�f��;���W�!7�]��Y�: r��׉t[']#8����$��>	^��j�L^�	�0xn��:��ox��(�[j�E����1q)�{��q���ߗB�j:��$e��ZvDu��
X.wra�|���+��F�'&�bY^uX�G@̜-<��Sp���zq=� �/R!/hf�E��R��)�fy�Z�׳x�1�'�JK;g��a��jy�,���}d�4��%�
`m�V��T��n��{V��E�b���f�{����cy;5��u!�[S\��Zs,/��7Ɗx�;��q�Qv�q�W^D�5z,�4�5d�gePZvT���n�)s�����;(W	3iڜ@�3..�%@v��㽗.Q?z J)l���*/%��"�+Ȧ�����>)��ݙp4��z�G��iqF�Ha�E?7���o
�u�E����O^έ�a�~�I�dR]d\�k��̧�E�v'���EqJ�Q{��,nѾ|݄�ե��D�nJ�A�g/w!��r�u��,�<z�nȊa�8���g�L,U�B��Eg���	�����S���4.f;��#j3)�»��M>�$����q�\��@��9c�������
�Z<F]���g�(�+����t�7�Q�%����ظ����z��w�p�tc���q��,�T,�%E�z�]m^J�O89[�Hh�l˱�����s��-�������D=y����Q���s �xsy�T�>w��\H�<ܺou�e?�㬝;z]�x�&Mr\�2�GV+�l�7 ڪY&�x��LI*p�J.lJ���kݒ�BU3j����xN��d�.��t��u34t�y���b��w���lm��kZU�;���=��������޴�t�8V��/\���,��6n��+ڗ�)Y�#���=yUۧv�A�ȸ��t	e�}(��)ix�!��o��ޚ��ԦoHʩ�\��M�����ð���wѧ�j��#y��Q�x����yq5/�+#�k2�l�d��Z��g�9cB�*�>6G
m_^�� yx�#����\IZ䕮IZ�=�B�t˼�x��i<�JR�M�K����Ng*��v���%P[ݏa��͵��4�p:ȧS�Ar����8�6��*��w4����wQwܹpL�h<��v4KW�/&D����؝�*^�B�QP�+��-��o8����S�D�P�e\U��lq��D��][��h!��qEμe]�;Z���o��CX'J�0Kn:�p��n��_L&:ō�s�#���8�]]��9�`D��ޝOn�i����!Cj�v�4e��ŀ�����̴���_u�TJ�%�s5r�ɶ69��9��G4:�չ2\�E	X�+�/��2;+.����,FOG�k�)gŝFG�_���}G�/�>z�cV���["�U�E-&������Y���JY
c��Ae��H��P(�Ӥ�����N��&f�$�rT����]�2�%KR+;�v�
۷�4���k7� �0X*�R��ʌE�|�ԸR�\�,q�0|}LD֗y�(��/����Z���)����=OG�f��{֗2�Kh�Q�*�f\MZ.%@V ���D���n����fBn�X�-�UO-"ŌAER9m�Q֊�1�k2+�bVc�����)�m�
�)���̸��dp�1�iE�Zx���X�McVUX�EM4}�<h<��ŌDF�V���(��[��j��yIX�]�k:*4���J��L���a�ɗ1�u�0�M��x����D�3;��=�ې_<C��"㣜�<����0ΤZ?oe�r�R��K�N�㘸�<��2sKx9ۮ�N;�ȓP��6$�r`;�Q��d�y��/��k�@�CDl�;�XYM�嵯��U�U�}�����5��=���#y�z��7S�������j�]��1�X_�(AW(~�w&���}T��l�甠cJD�0j%>�}����AP\�����:�8�'{`��[�|���N��>�����f�v>�@��3"��{�����%�ճ�`�)q�-��I�}�r�y�B]��C�����G%7�b���V�ڛ�����f����}�RZ�}���!5��?vK�0��Q>�f(��a���x:�mĩEm�3��p�Z��PX@���r:�E�����o�+��)�"�r�!=�Lw�A�ACэ��"{�Rw��E����.I(�L��%�d٧���c�q�<�q�0�t͑��pz��i}�_eF��R?Ki�SO*�T�f3`���l��X�[�V;�9g��Y3"��� jS�KB�/2�<�/��;R��cH�y
�,�Б�<.�U�Z����s*�r.�tf���4ZJ��.�RS�^It��6��n���W>ʱM�55L�̵H  9����MѽU���#��JWp�����S�Y��E�C���G�=��t�T#��.j�㭊��#��C��=�0���.=�qL]"�(�V�	�L���A�@�Y�5dd+���U�A��z��i/S"0�อrt`K���Z
�enR�m^(���a�[(�ue`�;���]��v���(�"��,��ލx� �fc�F[ƯrQXٓ�+�LvԼ�������`�fMCI��aei���)��R'��쩅7~�7��w���d�
����/�\���k!�5k�+�u@��Q'\֘�����yH+{���+�e�X�v��,�7�4�����;�.�S,P������l�8�Y�������7C���O�&κ�b�0�W���ٸ.��tR��B��������k
�j��2�ˁf���G���C���?z»����Z��y�S������O�Y���Y8�-�V��O��Z4��;5e�8���pZ�z�f5�z�]��!J<~�E�hW�,����Э$w���b�7�z���E%�\�	Tx���Q�H�=#j1(��:J��U��S0�ͬ8(��-Y��7N5Ā�2���û���ɕ}�a�Uͮ=��<q�v�ӯ0^aT��m��˔��x���;3S}�+z�����ڭ����SXJG�{��G��|����j���DN��kQ���_[��>J���'ݢ�C��Z�a�go!�a���=ht�`�pF��-���9�C�UM���v��k���`��m�m$�FtO���P=]b�*&X��i^N8��iVO-=Mx�t�.ְ�wV[�AoLb��Q\��Pxm��lm�}���=J�|���}���Yg{|q���y��w���8V��'��)ۓ0����[χ�br�%i���{6��p�h�_nʰ'-�����Y��F�i&�X斫](ة��@���w5�ɽ��H�m�&���ܗY�'ge^�s#e�ڳ�9?M�`��0쐴f��w�UU ���x��	��W�-[�����.�}��2�F�w6��l�o�}[�!�|i����	��n�o�z�]�C�c�kF	Ç�W�}� �]��\nC����d5V4dYZ:�"���;T�\t2oѱ��[Ό�'.C'�9ޡ�S)@��#��J8�_.�&a�������Bȕ�#"f;B�W�N��*�p/������Kk�nH��f�zo5C��-��Ma�QW�R|��u����w�P9�I<����x�	[����kl6(�]5��S�\<N�|3�NS�^N�H�r�qI��|�C��X�V���8��D{��_T�ɿ�6y���	�:I��H�x0+1(���G9�*t�X�t���a���h�So���\Auq���w7۔��3�ï5�� ���F��msY�{��Kל�Ƨ,���lZ(��D:FO�ܧ��T4�/����C=ʣO��ᓸ���V���26苆]�hI��sU�����D�Hɒ�^�{7�<��n�y������1�3�:ӄ��wo:m�#�]2B�QXr�v�{�^!�)K_��gRW���aVJf*d�7�
�$y�7OM�-���T�;��*��KA�u)���]��4���k�R�+o���2��=�6���˘���5:5{�Q�^R�e7��m��qPhFTXN�b%�A�"5vc�6ÎVW�@��)ctm��ɤ���c3����{�y�}*u��W��a�vl�JN��~r��ߧ�IhSZ�I��.�t�.NijY�a�K+Pd�;)r����x.wv��q���z=7L�E���mD���io�*쏝m���X���Δ�OO�S��kie�n�YY0�\hR;�0n��g����C/0M���L�ޓc�׉�Lί}�j���dT�����!�Yaˣ���;�*]��*���u@�Rv�f�6J�6T��\�.��pnv���������ν��*>��S)�{�O�o)��E�[I	�?b���}&���$��
,�oaE$z��}W�	Y�\X�����1���"����u�z�G�pҌJ7Y=�0H.0��&�o[Og3*cpf��޸�jFD�7p�o��%�"!_:�=t���]�`ᦀ��p�^^�#EΗP�(\�_H'|#[��~b�&�D^������ReǕkglKPȧ���/}�#�iJ�ܵ!�j$%=9�TkWD�F:��MrӐ�2k�)!+�*����E%��Cv��R�T"\wt՟���_�ZK˼��o�\�Z�P�{�ǘ��)Ώh!�7Q�+:UJ348��$��u^L����Ă�w�����:��uj/v�_y�P%�Զ������LN���xFk����cHu�����U�-�[W��^�E^��u�_�s}\ftb�Q@kH=Q"/s��o�s;ڡa w���~�p-��(HG]���H�����|��n�Fֵ�8�e�����[��ޚ�|�"/j��Zրm ���	ڰX$�+:�[�y��!w�b�|�8Z���a �0]o[�u�12�*��QyŝY����f��TX���'���'M�Fc}V�#�1.9�v�;�]}��+6�t�բ�@�����ﮕ��t�`;lFM��*�@\��[O![��,y@I�R�V+�y�m�H5L�j�CUp<xV6;n["��Pȟm' ˧�՟o\�H��t��T�Ժ.Lƞ=�vW+X�Hfj�U�$���K9�����O�=�+�O��"*RQL���t��X�2p�@	�~��W�X���F\�Q-�z�!��w^��#R�N���7�"�e��>ҝlc�2���:�4n��S�����"�]��D�0�GB�օel�Q�xs��H�z����3>��8V�1��DW%�v�Ǭ�`gN��k�,AM�z�-���TŨq.���հ'��dG��q���-іۥ�ݵ��mp�/��t2k��,�\M�r�0kT٫�$�)j���h��j�5����l��ō�셳nc�r�M]e���B��۫��$�?%���31]8Y<��������8��Rv�vZ��.����������₺[(p��i�2
�kjӑ���VbHa	�8��ݼ��4���r�1̲��*ݟ��Y��\���T��PQ����9�^�޺x��iTU��G.���[���Hz=��i��ۨ�����xH��v���ot��o/y_^ȉ�� ����]����gW	��c*�Y�kJ�F�1�j�c�;���[�,b����9mev8*�wcU�c����g��i̾�l*���n0�yά $���ێX�N��V�1!�k3N]�URi�Ŷ;z�+(��͡V�:��T�S��b��Ż8�6�Ǹ���oÙ&J�W��yXre���Zֈ%b*��X��'m��,�i5kZ*1m�*EE��U��Qwj�U2�b*����͵D8�����1b( ��Tv�FڌE����y���K���TV���*6����=qDAX�Tuh�ߗ"#�EQVg���a�5�K���و����DQ��At�ڪ�Yi�1r�Sv�h�Eb1J�.�5E
�W���j1	�
�4T��=J���}h�Q�����R��}�QQn�"3)R*���4g�c�5DY�*����Eb*���U���UPX�	�C���{�E�=ћ�ɉ��q:"k��zv�9o�s&oY��p�����}�%!�N�c� ��H���ɕz�	<n��1q���(ʋL����j�t��i�`N����TMgg�õ�;
_�ş��o�#�k�3���-7�;�.���_l]�Iz5�H[;DT@ܒWn��k��x�*8es&�Q�u-�9�s5��CI`�-��6�'�6�.��*�7*7D���3�E��B�jԱ��2�5hNVEӀ�c��K��G�s�QA��N����<���Ѡ�8�D�����s]�/��#sE�]t�2�HQ���b� A�е�Y-+4MhbgL`�=�<��Y��R����Hk�x��VE�R�6�D�f������}��7<�������M�v���N�x���e���b��0����tM����67�5������U�2 �c�+S�]=�[��֍�]�*/t�4��_gsb��9P8�<\��Ը�|ֱ�h�D�㧽H��#*�U��1��0%���T60OA�Ɠ�=#W'�E� 8ꤏC�U��Yr{V]/R��[Y����9�M rz�`�q�q=h�V��Ǹ�Xy�&]w�g2l�w��	Tu:�Rfi)W2xEn&�XzH��F]�kT_Tu*�\7.Te�O/X��nm��;yk�5֡�ˮ�.���DaWw�������*����\��rŐ��B\�Y.\ry���U��C��v�9��üQoi>;|��ɥ��gy�^%�~�?O)��'9�:j�v  �m���׫X
���n9� s*�P��m5�Ι$��wꗞǞ��������$z�;Q�'�D�yj���5�qLl�"�0KW��:�C�C��i��E���]�|�"웫++�`t^��*��o�M��{삓��ݍh��S�G,�h�[r�k�U�D.�v�'Ku��S�P��/�u��L{:�*eV�y�1���9^и��6j���s��k7)MѠ�]Ggg+�P|����,�W[��Ve��@ ���������)�����
P�������&g�ow����Ԃ�T*��ܑ~5�waF�J�r-�D�6���.1� ���b%n��N�b�.ͤ�9D�r����jj��\��6��s�����w�8$t٨��e�\�["���w"���q��'�2��kmrLSW�T�g��q�C���C3Ku������f�?�޴"�.,6��w���y���]��
�>��	������a[�틄�f
����,o���{Tꡝ��8�̗�x���2�>ԥe��C,�ݩ�[Y\c��goc{;&��%�E�:.��U����w} ���|�#$E�x��Ond�uk�y��M���,:�?e ���{����Kl�KOnk����D��)�{3�w��YU�G)۰8fE�9j�)F�㝪0��������]	2)h��%��J��	�WW]MS灅Rٞt�9К���nK�t�a� :�U����d��P!�0�3����n�k�/'����q��s�`��F�[���M'P�J1��$����'��<)^LR���9�{Q�|�z�vi<����E���F��FgNE�L�c	�7���N'=nq�֌���E\b�)� op��p�VzWTǪb��a�{'$cf{�</f�y��5�3`��CWf�]G�9;[v4�4X�qQ{�#B�m��Mxy�x��v��{ՌU�R���8fѾބ�\�tQ�m���P�n����z9͝V�qt�<_2����~t�/���4�я���#�n5`di�;հ.�'��p{�5d�2��ǽoFqCtK%�Xd(t�CJ�ve�a�j�B�k����<��D��f,T�#B5�V#f�ͫ�iE�2;D�����:��o!fe̢[�&��&���*I(-r7>�1��l��䧔���ƻt�����VZi�9��n�!���(h@�̽��ꪉ���_��9��Lq����嵵��s��Y͊O:�yK��l@�X,P����뚭qS��R�ewX]A]9nC�ʹ�2��&����+�=��pb��	f�����{��6��>�sx������-���Ѹ��=�/�+��ͨ�в�������5��?F}Niz{�Ƃ9C�������6����3J㻁���f�E�f���n�ڣx�)曙�G���$���ˠ����&�H-7���(�J�s��Q�L1]A^�aS`J��#3�]]�]�㮜�k=�6�e��4wWC}Z�ٻta��.�M)K��̚Տ�lbf�WB�̢~�$�RQ�}#Un�T2/�ŵ�6�$(ʟJ�T;X=�K���:d�P�kN��&L��9�v��P��ё���01e�w]�{�����;�;�.v��+����kHTz:�J%hf�*它k��i��vog�H,��',B�T	�"�q"+�.-2ݮ���_g
ǵm�x���4�r��\�y����t�U��D�Z6/\�X�J�z�S6{<y���3ܳ���{9��<u������ ���T�6�_���&?#�����c4�WaWR�U�J��0E�f��Z�p�c�U1M�\낰t�I@k����ip�N�����e��co�{��;`]�ߪ9s�K��y�������U����^����?6~��h�f�ٽB�m�5vw����X��AĈ�wC�����d������%�e�u�3o�`ȍ�����963vs��p�dd�C�Ol�i,�'�-��{Q�b�}�.�����Q/����a9f�4��Ad�_lV��W����R���s/Y���������6)�(�Q,	ڸ�!R�(<�*�`:|�W�qju�ub�Y�*�ÌLU^�^��ᔎT�N7��'-	w��^w��C�/,K�"H���޹�Cru$.�C.�j[��'�����';�{5-�w�cu�b�n�w�����ɺ/�R���o��̔�aE,WW�]������XTڷ*�����i0l�)�e�X"l]u&v��p����ȉ� m��R�.ZB@��hEAu�Yh2��,�<PK�E��ڽ��5fZ��j�Tp*G����k%Cs�ӎ��ա�@]���9��<�M�]���v*%����b^;�t�$[����{!:-מ��v�8�p����=��\M��
F�!�f5j���o�a(�#"��6�\mk]+�<f����&x%���ou�;X���ݴ�]��̜I��gm^kZ�+�WUD�uV�鹼8��ڒ��2�CA�t�*��I"�A�fS�Z��Om�|�R�&k��i��\.%g�9w�*&����Xs%i9��J6T���2D��|���p��nz�{6��wH�Z.\9Ƶ`��&��1i��H��UMѡTE����ɳ��sೌ���*oqBQ&�Wi435)6����2��k3Kf��Ŵ~p횓��Ԣ��J��6��'�ᡛъ���a�r]�d��j����Y��A$L�r��ȏjqu���u��K��]31Λ!ǒ8�*v�dt7]�jY����S6P6�^kr�qQ�wn����5�^nv�;m��2tX����mS�+���i���(�4%�v�kiQ��W�rF��1�e�_߻Y3ar�:f�3�ڱ�����H�rٛ�R���ƾ�����6�m��z#�[��a��E�MxmLV��ܱ��V� �	�;�9]c��@�����j��]�2�mJ�vn�b�kT7To)t��1�N����H������"��W��8�ݕv�<��V� H��G�ZN�[emm�R�7��CV�����Ց5��e3$��V�f'��O���!�k���9�Ꙇ�R���i8h�0�Ʀ�C:nͳ�G�	�ݽV�ق�C�uuN��g=9��X{ㇹVQyA��v��s�˺��xm��v5��3�N���%~�,v�����^����2���M�R�vcC3_1lS
s)��W�hԿ���>uGF�Mm���aݼ���+y�l6�xB��o[a�Қ������{��.��������E|��%N�F/"�B����A��
#�h�j�4�TV"nܥ<�3���L�UF*)O,���O-�ˊ[<CPL�PAU�Tb"��2�9s	U|CUb��b�%H�cZEG-MZ�� �*"1dTU�
1Q� ����ł���
�(�)j����
�]Z�n��1Ae�Kq2[EP�2�QOm�"ª,X-kE�Tm�QƸ�1X����ਨ�X�M9l�[J�M��DZ�#�j,TDc���TĠ��G-A�c0�4檔aU�Q����d�-�	��W-�=�JW�ʕ����kN��=f%�b��i1=[˥+���&��j���g~��/o��o^��t2bj�=�{���.�V�]
Mr��Bڽ��p-)�����Nyt��bta6�����|GTUؽ�5�/@�q�5z{���{�����.��Cb�A�m�9�*Χ�X"���]q��h�4g�T
��oJ�EF'\�x�t�2	�@秢�_��x�l��Hw�u昚�kl\%PL���Î�08+�N	��e�i����\�ф� 3}oJ�c�g/[�b�g�62�|����6t��صkn�}���d%�m�/R�N5.�S&ůs{`�d��-R�ׇm��t;�laX��
��������?i]|D��8��ee+��;Ć˰�b��dn1��fz�r�����vV��7�=�J6�Z�uP�U�r,��S���Rx{E5��QN�2)��`��iߟ�7}���A�L�ʿ=��3;Ќs����춍3����ϻ/I���"a�%�څx@n��<��lp,�����pv�qc�L���p�͛8:U�H)�aA@.&��L��W��7�y(���:��%G���NAA�/�ۺ�m�6��N�Rh�]wpf��c\�^*�bz�}=��>cQC:/]��(�9Q!74��K�i��e�4���E{3_eGF<Pkbt�3{U6�UY�3�C��ش��9`	�;d�RZ�wvA���0dY����p�^O�}�1������1�.��ź��\�z��z����X���яY��+��!�7�ҽ��+�ʅ��e#P(����`Yz�<�����2�ݸ�B�ċIaZ��+j\���Q}����+���GVr9Ͻ3@��V��ಳ��:Ǽ����[�3"k����tOսt���6+(���:��	G&H ώ�dl��zu��ev S��i,�e��b���(̲�T]ٰ��: 9a:�PnK���9r��rT�Gy:������-7N�ef��j^�v�f�7:^ԤQW����'�)������)��G2v,r�"w���3y�!\▽n���&�S�ǟG[h PQ�4�d�]�+!���r�F���r9�5,���Α�
D]�Igl����7�I�y��>���wR��B���v\/����k��`�%��nk�3:]��;��=l��|g�g�׃�&��P�t��M=��M�cj5f����"Mi-��J�oB$�r��鉼Z�-P��3n=�{2��k���N��'u�+<|�7��y��9�\�Jt��	2=_P(�f1OgE/�3�r���k�w��Wz�A�k<o:�:X/��y�(���wx{�Os��֣W����ǂ[_hˍ?fC�C"U_�`X�@	�4���x��<��9�\�](t�sD����-1c:�ш�f4����|��,-����8��(��@ax������A�`�?K�j��*��U���Vj˴�]�%l���9ӢD�Ν���-���j!� E�v�e�]���&�{����G6�^���,
�֌y�Z����ٞ�N�Hr�(�2��e�8�u�����%�v䴂�"��P����W���2Ε�w�9��]�UƮUқ��ٵ�-a���{X��r�S��Ϡ���+x~�Pr���(o]�ԻXwX[��Q@@�<��l��A	�l��	����R��,9=nm��͇�u n_d�{�x��eXp��W{�~�K�]�ގX6�\g+�G�qyׁ��r�����Q���%%Y���X��T)����=��Bn8�8����1N��O+"�wn6�'����Ν��tn�����������Gg8�-:��/�_ 4;G�w��٧��j\e����^
�:����P���\��ePXa���z��]s�A��������Pҋ�7��0>�:�`�b����v_.yS:��� ���W�ֻu���m������julˁ>�i�}�,�i�x�)��ЏO5s0IW�p����f���$�s�����)w�Y(y(����z%�p�� �#,�4�]��v�)֭溻p��Bc���K��%��(PP��`w^���u�Ln䤟l�D�!Ņ�aG�~c���b�l#��:�R�]�2��}��s+����k[��U��ŝ�Y�E�{����w�v8MF0N^��6	��oV��Hׅ"I��8B��$�xp�M�:Z�P[W�8[eq�hT���6�Bdmw#g�k�mtcs�
l;j*@�5>����a��F�6��9�	p�����{���q���Ž�X�����\"�fB�C*�*�6�fJ_G���+�߮/�TT_����������|:Oϐ:Vu5�/U�u����n�Ʋ��M'?~/�^P�~}n���  �V�h������i��;��5�#�Ou'\��ѣ�[��h����M�py�U3@����|��-:� b-T6m(1sGzhtpۘ%-�nz�QL+�'/9`=�R����}G����x�@�J�B��Ṭ<:��p+.tܰ�N�U�[�7m(r�C�^'�����ˇ���sYVĖ���3m$�5Ѽ�k��U΍�?]N����7�hb��ӊ��+6Xw@K�-^3{�E*�
;��%A�%k�=\���Q�Cd�Ϯ)����p{�,�~F��q��&���]G����q=�C��n)Nj���zRz�,�����f7��*�)nn����61l�;櫚�i<i�a�X��x1��YA^�<v�6�R����
L3���D��D2-�-�@ֈ1��g��3�˧xY�j*0rN<��\kʛ��n�x-i,V� ��:6�\N܀A�5�z+�v8�C\�ԎY|���eѩ*�<�ѮG��~��c=��j�M.]t��+�YY6�:�h*�e��������V6��~������4ηe�f�՗��-8�rүi�E=��	-���N�&���4°��=�yZ��&� ?Gٿ��/�z�Ԝ�q2�Y�q�lY"�D�#	�� �<�T��l.�ͬr��̘Ep���"�s,-ɾ����$"���Bl$�E�Z�c�A�-U���=$�^>G֝o�X�6��)��,�����`��g2��1 ��E��`�D���%m�k�����q���
q/�M���Y�\z����9AVz�ޚM�՝�� ڱ�أ��w�Z��U�t�Ph\�B��v9B����-"��Dh1h�Y�X������&""#�&EPT
D��B�*��%�U@Ѭ��D]�&Xf�����%o�jzT����j-��3R����!QI A���$	"�!���C�)u�[l�62�����!@��1�(�w�xg}����:f��.��C��Jˊ�_��C+Θh_="0o	X�@�Qg+d�,�PT�5|,�ק�XC�@E@�B�*�Q�IZf��+�8�q�����'��?]t��@����=[�����
���s����D�y[�B�k%�h�w@�#4��j@��V�3�K��p9�x���6W��m�/4� ~��
����Ts���K�E*���U'�
f�b"��%	���iN�[ɳ@����AP5��Ŀ4�ہ����|�H}���*>��f����E|�g�2y�?
F^-�95�2*��[��T�E�������Co҅����m��K K�>�����_���DY7����n۲���_˯��r7Ȩ*ר��1�Ǥb���d�8�$�U����G`��f(������E}�LJ��j�y�2,	�a�.~4EP.6�" ��hЍ��0;# E<)<6$������5�ޙ��}�԰Old!gRQ�O ���)�E�W	���
��@��v���8���_3��F׷ha=O�X���������6���'w_ �Yc�t�B7���N��H��'�C�nJ|xk2
��y(�*A��m��ރ�$����	�*�����a����������ԛS[��٩/dȆ��$�s��@Qi��d�G��L���2g��#���P��Po-���dT���X3���H���R��H6������:�˪�����y%���7@��"��0nA�o��ˏV��x�r@\+����#v�b�B�S��R��a@=!đ{t֎�ܟ�.�p�!�5Q