BZh91AY&SY�^�
�d߀`q����� ?���bH��  ��"����m��4VH١Q
�H��K�B�(�%6e#5e"�Cl*)��
��m� ��a�R�J��"kk6.�TEٍ���+ZI&�Zf�V��RVږ��Z٭�0�V�L�fBA�T�m��6�jH٦E���"�T��I֦țmih��9�2�6k*����VT�j����1�����m��i��0�,f��ֲ�i&��4V�mcR��J�P5�jm���Zٶ��Զ)f�M�iw7"B�R�   st���+Aٕ]��j(P�GMsj͗u�W=�OU{6��n���:ٖ�v�u��mZU���i]f��]W��:{1vW����Q��M)�XR�[26�ʯ�  w}N�A��.s�@�`#�� 7[� �9��<=��A��מ�QѠo/k�t� 4���>��x��(�{�}>��(:�w�Y�f�j���͚Zė�   �{�� ������4�Ư8ްhh'����k�x����1���T=E��<F�=�{�O<� ��<5��⻅h(=җ���Fm�R���R>   ����:��������J�
Y�k�R�puC����)Р�V��=5�7����=������!�� @=�W� �Kz�-�Pٵ����)V��7�  ��v�-ϵw�h��oxݍ ��= �z��P
+�����WZPҚ�z�� �=Wp  3�� N٩��IR�`�(h�   k� �{�������ӽ;�-�h;��=� ��y�@����w{���^��oy@P��\�]:�w�n��raN�ۡ{��kmF�l�����ֳ!lо   �� �w*�t2��j�� t�OgO<� mwW��x ��;^^ �{ޯy���G��=iC�=���� ��q^h�Z�Z)���kEPhž   �Pw��>���n��:`Ae� 9u� �5��q@:�۪�Aꗼ�� �תq�z:�s%*UU�m�kU�-��D��   c�`>�}�P���:4 �:ۀPQ���P �Sh��� =��@���=�`Ae�IV���B�5Z��m�5�   1��@Ϋ@��;��W��� '�^(P���;��� ��� ��� 4:��HH�T  �=���J� @  � E=��R�U� 4 ����S�!)T�� @h  5O��J�h      ��RJ�U6P��h4����&%L�I�M�&�����bw��&_o�/�����񘬸���|��=�\�ɷ��^�����ϠI �	9�� H$� �A �?A�I���D$�>������G����`�F��H�I��w�r�pwq�����"q�r<�I����|�
0�%� �<t<wB BМ'	������ BЀ��qЁ�' �C�' C��C����B C�' C�=��t<	�����pC��'wC�t=�BBC�"pC�� Bwt!�	�Bw qC����qМq�'#�wq��C��=��<pBw�wwBpp���pq	���'Bwq�	����C��pC�r<  q�w�'pC��qw�q�C�wB��C� wwC��	����q�Ѐ B��pC���p�t<pp��  ���	��C�t!�wt'wBwt'wB�r=���wBwt<wBЇt<wC��	�C�r$ 'wBqМt'q	�BqЁ� �@� K�������_�~�~��'\�ޔ���7y�Y��������2Y���mv2�e'ͳ�uu`Qa���Cn��3-5�U�V��ꝶ�Օo/@b%a���Hv�)`z�\��p8��ԁU�G.*�mܠ��Z��N� ��Pz�dB�,"{%\�i`*�Ue�o0��I���aaPۼ�����QѮ1BD�m�6�$��8F�y�27V<"�d���ӫ1�zi�%E���h�+fA�Sk*�J#�$��E��ŕf׹��ldP�k*�a�[��Z!��P���\-a��Mm�;D\,�(Сi^��U8a���g&i�;J�Fi�C����Gg��q\��h�N�v$�;��9����y3,�ʸ�[���D㻫�;/M���zl��K٭���.�bOD���[w�^��Z�v�n)�e T�?%E��j�*h;b��DdI懏a�P'�l]ؗ fL[���f�0X3�����a~sT���mK[��^�&vQ��cB���؀���#�X��E�\U���!kl�A�C8<�ܤ��0FWՙi��ʭ��3$Kc�4�ĭ\�[�*�/Dz��/(jgi�$�a�t��E�k�)��<yUL�/0=1�=݊Y�H�t�ߜ���²8��f�U��m����4PJ���Mf:�C2L��t:Ȥ�]M�V���i�w�6ʶγ�:��B
w��%n,���ڡ@Ȳ���&ss �`�d�/5��QfX���ӵ[	�Źv��.̌f����`�b��i��9<�v�tY��څa��r��L���������$����d�۱p�a�e����D��!����Bf�u��7%�P8(Q�̑K�h�튥���Ѹ�V)������[��Q�ke@�.��(3���Ѧ*OeT�bՂ]n!��d�tY�+7A�-b�1�L���%A{�,�����)̏h=�0��(��P���#.�� B���=zl�CXcp����q^<:[VPH�j�+12o�
�������W���^�6\ەn�%�U�v�3(Vշ6=�W
�K�Y�M�/s��.b��^�d�[`�AӴA�[���aG�,E/]KMJ�k6��Ƭ9����t������Ȩ�y�5m�)<��f���S(�Q�k	���V!{�.CLj�$�6�l�rm�S�F��e��� M7N�1�F~kVipapf&��*���2���J�������Bܽam�Q�dj��xU�Ɓ�kA�h�R�w{{e�W��������;m�A�wmhg(��<�m��゘?3��2jͷZ�ۊ �yR�%3m��ԛN�l����h���X��^:�)��w.!�����DIBU�j-Hշ��OU�u�����Uc�� ۄ1�At�n�F�r�T���"Um����-�&֜�ٴ�^��h*`n�cDg��h�ș�y�d�B"l����=YX�R:K²�ôc��`���J sV��R�67W/AIQP����D%%��ڡy>�h��f�ڶ3Z8�i0қ�xo��r�E�%��R�Re�I:h<�����nS9�mK6*kd�.\�v�a�$���`�Ap �6�2��nS�����
��z٭�*�-D�*�;�f��c�AK�xq���a�Cf�A�+/SF];2�.���h�����Y���"ƭ1% �T,Q�E�E6����@���r`hl5G�p���Y�u`�]X:w���"�%�/N���[�j�Vkn�2�#�ݕniY�[�i���V�Bcm��-�:�'-5Q��	Z1+��e�.چ��P�r� �E �M�A�B��)�]�iݡ��Z�Iϫw\�m�f�vL.mX�;j9t5P�^;��`�t�$li�Z0@��
ib��lX�W�
Ԧ�~H��R@�֮�$U��R	���KOQ�d!�ē�f�l����8��w� $k#��ʅI{R���YH�EKdB݌�q�;�ܐ^��=�E]<H+ec[�_b�]�����Q;E�!{D��n�1�)�g^O�&`�*����&�O�n�&r���}�Z��Є�U��&5q�X�S�yToc�6�
4Y�[r���[��y"���0�v}�EX��jO��`����AԵ��UDm-�z;�xһ[���"�}��N«�Q�Ze"�m��l��G���Z�������&��m�U�qT�4.Q�;F-3�����D��eŭ`(��f�㡙�c (U�[��ѽ���p��q,pMʳ��/��SIi�憪�4�z�-2���n�U�6���ڳ�h����(�^ݬ��Nn��j��YB2���)wx�B�=��bC���v���jl������?A�w`�h����ͭ�Y�&�� �.�v�n�툮*X����	��!w��:Me�,���b#3e��������J�P���ܳI��� �a�>��qm��I�T��$��
��cܹy,���zi�ZDe
��X2 1�5�5�F�x	�Y([6�C�KoT�&��F��*2��Я܌1�v�J��)�0�i���%�QV�m:T�A�f��KL��Od�#M�Ri���F�Ō����5�h�1��ɺ�bPn�5�M,v��*j�6���
Xr���y�J-�e�]m-Di�rk=�ܼ+mP,�q���+����
�$��S��M⤊��%���-\�5�2��� �qmh�CL;zDm肶����[�j�v�7��l�WZ���������6�FZX2���Ef�m��1Gw�
:�wP�n7b�o, �������U;hH���-��Feu���ҁ������Z�K�E7�Sj�G)�u�hNI2�1��p��u���Nވ�e:�J��9*/LN �4A��0��"��G)k��L��յ������+N1,QGU(Ԣ�G;m���� N�k$�*ң)Ӕ��b�ڼ�:�$�8�C��Ma.V��a�]�<�b�(lR��j�q�3.���mn,y Im华8M\&ƍ#�	zʊ�덼'h�nT���h�Ӯ��T����DM���:X�@��D�N%{��t�S&���D�L{�v��ǭ����P�~"��GL$�q+�[�M=��u�JK�a���3C��#��h[@�.#���<��X���N�E�	Y,���Y{���Zps�oFn3��MڦE����.��)t\Nw�o7���-�(R�J�C4ܦFځ���;��X�xb���,�l�����ۘ��y�d�n�Et�mQ,�ڕv�0�kL�u6a�6�;4�Q�W�y�rm�A�e����ɻ�4�>�f�����ǃwK,lϓy/t��ᗺ�s뭓tw6'vS�е���D�&i�����E(V��R�c���nZEe�kt+̹�i�Yw�#52"���r'C$��꼚�0���.�k�ּ:G�chP׍<��1[J� p�p�KF-�0�d] ��k�g��q�
{Y��:ķr�H��o�[�4��6��^�u��K��>�s{`́�W���?�qJ���u�%��Kt�v��$GYu"� �)�1�F���o5���sf|4Y��4^������٘p�su�TM�P��C��XT�75�2�Rmh�v���d��r��׮�cHa�K�X��k7
��^�R��RP�VV�yaR-�w[7�)��ߐtq���i25��ͼ��매mA��oIqe-�%[8ƜN��UcJ]�v"�fE�7Y��ԖY;WVҪ����2ä�V*]�.�&i�oU�b܊��D�ͱ�V���HѬ[Q�e���uy��.�G�Pl[SM/�܎n����B�j��J-�����M
w{�����U6����!kaEj;GpK�dX�dS#8f�xJ��fi/7-�X�����-��/D˖%]�G�M�R��hy*D^\kq��U��Q�vm�� :�˄:kۖI�w�H��'��Ku#�z�+5�*��=��˰��UsU
l�ȝTd�lf1ј�nl4��K����x^붦C�	���9��`�����n����M�3��Sq�a){V�dĞֹ5�6��Q\��m-_#W��/�˽ׁ������b:��K��L݌���%�v�*���,}��E�SF���=�n�Tt�ˋ+��8�gi��e�F�R�A�D�cq�ᒯ&Ua�qnjGE=����N^���#s3+�mE,�#M3c�r�X�u�
�%�v�AU�K��p������CQ�J����&U
D���d�U,�9v��5��#\r�M�)�:C������f������!\����V#r5��t�r�Į�#���&����Z�ܚ�ġisJ����M��7���P^F��5zu�@	s����ub6-ֵ3&d��g%KҮ�Ս���3F�XB��N���fl�أx�*2�l�9s�{�h�rf��ҤZ	�'6�mm^v��%6D�CSv*l�mL�Q��Jэ���]ZW1-�P,���9��;���E"�̃d�Ա5ޛ���ݭ�K^Um�#9��e�3-\ժ��#��U�̸"�5��dא�+Mn�
w`��?�7�L�M^乳u���Ƀ
WwB���-�j+h�{�^��L��7�t�GD@Y�ifP�,�;[���U��+c�v��(�{�HE�`ӽ��H��*�ٶP�1���jĪY{%�����<8�KB�i� �փ�����zOZʴ��b���"�,܂�:YR�23E&�㕂���2�|5�5����n���H��o0ndv��!�����Zݚ���a��n�2�^F�$f�M3n�vw\&;�A&*�,ݭ*w�̃i^�y[B��"�4��nC�`��v���ʝ�%��n��1��KW�Zޣ���n��Ѥk1��k+yY�]�t��+>cF�/����.���⌂�\[��И�nY�c��֊y	�f�w-�p2�I0i�����=k����'�.�@����I`�s5i��v�t�&�0� ���j�*��wF�q&��'�L��m���턪iXF�6A��m��7KP�#A<Ҭ޹N毜��Cr�n�c��b!㩣bshmɆiDe�Li^���x�&K������j��!Q!�+�
=�ޣ$%��2�A9���MC�f�#N̈́晐���]����3be;4��v�N��Bt��F���h\�Ԗ�i8Z����Y�Ȏ��l6(�6���T�`�f�|�X�9���㥙�&n1+j�Z#{)46��Yd�z�u [V���is��M#x�_W�,��P�sj��,=�A�kl�7����Y{��wL�y��Q��̔�@��v�V���I0~�hD	Hj{����	y�t�iu�fH��ekI�u�_fݥD8\�����wƩ���2l��Ѝ�N�Өŕ
�3 `�-=a&+N)e�p��>,]�e�����vp��ĥ9��n%i�i*ǳ4���-�Vs\K�Iyu��k~Z0bs*�ͧb��3vaρ����`�qS�6yM=�*]᱊��++q�M�eޛ@���X�#���2�K�ê�k ��]k/L;+D��Wm��g)ʚ;��Ȓ��x���,;{6��(i��*kb�R�@J�̠������	`�<���`Ya�ƅ�q�˶E�����fʛ�F�&MM�u���pӐ�pmi�T(�d�2RE�1����r����6m^J�r�w]ܤH�Q-hde�6n�m��#Pi��R�Lǒ�z�v��/y�!�I�"��CU��ԁ�6Ϊ�%t�QoUe���է(=tLM�&��b$�ʵ�`���.nGk]:�e�upF���k��v�c�웂�*�0�pf��t5�l͙
y1mH �(��+X[��� -��+q��bY�Յ��)U�ĺp�a�(�S�l����tn��l8F��V6�P��ٻ��}{�;��qx��{O�qޜb�P�v�@�ͳG.���+m3��%�KdԠ���m�F��&�l%t�66Y�n+ݘj�%�ۋ�Oޱ����NǗv6m��/�i�JI
V����T4	t�D��э=�)�֨C�/w6����V��֙���)�U�n�/	�Y�VQ��5�DVV,�Cs4V�Lhʴ\���!��.L���4)S����-;˽�*����`�H*�mU��]�9�b�e�1[M�Y�ڸ �n�k�R��o(�j޲^���ƄT� Ъ��Y-豓)�z��
�D�ֶ1y����0
�v�c��Q�Kan��Ha�W�h[T�
���Q�B�:ϴBha��B]�bٛ�aX4���,#Ot�YE��k�u�	dX��I�E �2o�^��s��x�6(�.����9N�Rh�
-�P�K�X��u�%0ig+j���T�ڰsf��a9����u��ޚ��)a�v��ّ^]�F��	NKlO�7��ݕt��-��M�iVjxɽ��ޣ�,b�B�7(�Y�[̂��J7ʬ�n
�76��Л�(�:�[�T�:Rj��kp=�B�f�py�z�H�ʴ^��A��x�:���l���,��t�-/&B"�D^�5u&[��E�n#�r������J#[�ݔ�&>.�bo�1�V��r�9��&���7]Ǐ%iՇn���N�*���K
�BB�+x�oa��)gta�e�Qy%��٨�Ջ3H���-A�.�-_��ܳ��<6���DV�޷O{w�rwK�Cy�<�ek�����)���F��d�R݃h�ٻ�E�Yd���y��en�Я w)�oBlS����D�k-�o'D��	Ք@0�7G�+ۤ���'Imh�q;R`�иF=%�(�P���"���WR�s�j����ˇ���.�1�T4�9�ؽ�X)U�!�f���a��(y�݆��XO#o�E!�Wqj��P����7�'�ٿ���_g���׾}Ƹ�H����T|u�/���)��um�;���<fZ�[&�Yb�@�`�#�&|��2V5ݻ���ɪ��*$�j��1a�v#w�֝\�4���Q|il�������-������e/`��Z�H^^J����d�c��rJo������"F�̈́m��=��z�͔�#�9�*nŝr�]L��Pf�,S^�K;"�"MV�J�U�Gyn��DZOO׳���P�{�el�a���W��2iSQf�A�Í���w�szpC�&Qg�7�d��Y���B²�Y3^����v3�d�|��z��+K�0�綉�b�,���tz��L�!�5���ïp1��zTn�)e�,YKK�0�`jw����r�#�����h��l�Z��_f^�7v%��
��r�r��X��k��}��B2��wRSn\sej�e�;&�/�lّ�"�@X�9s`����}x�e�+7��5�]�6P�<Ɇ�ώզ�a�=
���|�wH�,�C�-ݑY��	�c���ڲ��3���w��q�bq�-�5r�s��O��.����&�uF�9��L=�\��*�^���y�_[W��Φ��(7	D�y��dhu��]ʰ�س�n�낏b�2Y�m�1�okE�E�oE���T�R\bo8�	��8:趯Hҏ=/yV���zF�p�U���gZs��i�u׍�nT����P��,���]�l��u��Uי�h��%qC2��4�����6�j΢�иC{dzU�m�5�c}�Ck�����Vp��xIYfs#4ݖ���j�iT��w79���ޠl�����b�&�}N*�b�{�e��گ��+M�͕�`U�a����:�g3��9���%H"{��`�J���u�/Ev�9��|]��`V�Al�m�il�Cz\d�*G2�ζ-�DFɸ��
��9`I,F�C�N[r=ԵI�j����[c��[Y�ӕ��ԯ��g���+1.�nf;O)���e���*h5��{do&���n����o\����t�6���l��r����K��Q8]��31�J�k�7�ߜ��}�u�nF��h��q�%G��v��_E3�='^_*Ő�v�=Q�R�f�ը�漵 ��fN�V��9��ÖpC�jV(��G�DkLXY��Q���n�n� â�U��n_,�Meb��M 8ˀ���+�L*��[G6v���Ts_gP�q�]e^�0���h}u.�I&������n��/����5���k��I���@U���u����B/��̓]�{�Yv�Z�"'CX�>�����;�C;�2�%��]�H�][�p���qU���ƪ-���ۀ7.�q�oC�Hh¦GO�k�+�:挙.q�F�M��FF�Z�27}W��ntN.�t��os��+��5d�y&�P'Wd��-�ׇ�}��[`ƺ�����ə�]yڊj�<���ID�&��p�����o2o.�De��F#�W�ܙ�y���Rx���ZL(,p��<j�a\x
��n��(�*�cn������X��1nc;P����_T��[�{���J���v���r�AI#]'}�2�'S��2�z.�6��Ǖ$	N3��{B��ޭ\��c'��X�������*Q�2��3!�K��X�B���E���y��x���m1����%�דSY���8,�kl�;sv����k������r�C����gM���d�Kmr*܎q������q5�ft���]�'G�Y��`�ysZ�&�^�qЦ�9�CR��v��sۼ�v��e)-�V��m5&�c�ְ���Z�i�{�ғ�[���"<L�=h�C�7Z�vMԳr�%]H�+3���%�g�;:h�7��x��2�y�Bf:���;Mq�҅<��.��oX@�E۳��;�*�x��w��lN�Z���:���eY�4A�*�����t9	3��
����pTǖ������.GN�]�sLj#`�����Y[:XY��'�j��u���Z1ef��x+��̹=���Q�g]qU�S���ێ�����lu���.]AC%����k˫��n�׮�Y�FP�7�IȞ
��63{UM/�K�����f����#�њ�ѽ~pn���^��l��N7�g���k�\Vo{AzH�Cd��d+�zN�~��5/4�5�l[`s�HGf-9.���|�r�E��T�îSyN �G��ߜ7l�}Yq�;//��[����w.'N&�r$Ҏ�Zb�!QU�+�vy]�W%�T��ގ�0��J�nE�֦�*F�Z�[���{z�kYY��A,�'�ge���[i�2��'�X��{�VT�z�RU�0%���ڎp:�&�
��9� ۏ]g+x�.�I뮾[P���̽�{��juŲ	e�r�e��{�^\n�~f�C�	47��/*�C�n
���ir]�.�}
+n1�����Va`B�p42QE��y�k�r�����)tʫ�d@r��8��BÚ�9��w��<Q����P�o0ý�8�٩�e��hE"�}5,���5��p%�,N��ܽ��z�'k��SL�a�����
��6��l�X0@��5I*vT���f�relźs��m�*��vM�ಓJ�K��D�f��hU)c[�M\�'��rި��r����`fHoI]��خ����y����a�a]SG���^JY"�ι�NR�q�p�"���{Mv.���Ԭ�7!�������cd�o.�6Zxm�*3�3MN��syh�!�gL7]V�@�'f�M��l�ʼA�Lƴ�c\}[��1ݙ�^��a��{H�S�7���{.��&�=�[���tw��n�l�:ު i��F�q+�7���5b�:4U�O�*��:�q�2�ѻD�-���49�ʅgR]�ѸcÃ
jJ�WF�kf�6˝�>�V�빬��i���b�}
��cx�7~�4YR�=�*�*�o�/+O'Nr\t��i�#l�>(�y�R�Qv���T�O��Ar��xi��n���weԍ����Tu�N��Xq�!PQZ@fa}�ErY�*�Aި�'�_*��n�<�ˣX2G5�0�$V���o-J��U+	R�ᥨs;ޙ���O4C/,�$�K8ev��ǐ�N=�9��-����QW)@� �CT� �s�
r�4�n�����'
grM�������u܏�E��S�raldBmNO��y�^'�!d�+��G�e�=Z���2s�����l˹���gL�;�]ynQ�K�Q��٧s��Ԑ�$��nض��s��񿅎ۨ��7kFس\���6q2\	+���_�y�a�V�X:�oP�8�m�N��WyNC����7Ok�	��14��J#��'H�������t����^�ƫM���UN�6�ȡ.���or�֦����p�wSL�t�h�֞�u��x��� Y/5�J�a����rPԳ���8yU����w';�#�PB��(Ed˥C��WgJO��J�%�i�;��@ņ�r�3�x���m	H=z���7���u�Ks%�]n���"�XR0�,�����b�N���z�;s���%������y���'c��sL�g��X��b���-$�j�����*vp4�]ɾ�z��1٧Liœ��N�N�j��yd�J�ތ!]�vm��٫�[�7�a�M�w'z�|g\�-�¯�۝�eZ�ݮ��{nw͗۲��4��z�z�ᛷrV�T_�9�����ֱ�.b�0���2������%`�,!c2����y�ջ���.��3�^|1@勈�����)���e����e"�f&�`��K��r⫥,�N���.t�du�u��r�5�nݭ�5����!��(`���ct��}����p�^6̺qL��/b���|����:da�!���VJF�1u1^<W��3V7�c����
��w,*�e�qg�f|�7O�MMW"���V��:rQ��PT�s������i"S��X���\�1���ĉ]�]��6��F�=�\f��߸꾮Z������,�m7���I��gu�����6�r^8�P�+��0��6!׳��6��`�W�3VK�*��=M%�|�[�OB���Ѭ���b��{L4b8)� �I��W�b���l��ǟ]<�1��u*�0Mٱ5���l_)9>/t>�B"�̥�&i�{����{f늁�ŠR�+js�	��E�A�}hH�c��n��ιg�I���׭���gq�r@��ޢ�X�֭D*��`j�F9��+s;`&v�T{l�*�RI�(� ���J�غ^N�	.h�bҫ��[\%\@�^�5�LvWI��}i�����GS�6�y�v�n�Û$����l6E��I9�A���z���.�f���ũ[޺�p�R�3�'Sl�T�,Ud3��.�pDN�i����4_nY�Z�k�8i�1���v�U�����Q'�����`�}s��s�+U��qs�7�c!6wn�����r���r��5���(Cw��oثfl�j��1P�f|��(L|W
N�ZR=�7%�H��L��i^�W�u�ki�X�=0�r���\Z,�k6Bo�z��޳�}8P2�"��\�ԛ̽��l�zL,gb,�lY��s��4�R�S�;5_X����N�xK�gY�Ykӹ�7V ���0�P��0�bN��޻[�����QɇiԆef�����.໮m]٪��V�W��kgl&pL�o����� �G]Y�]%�7n����� �F�y�!ޠ���`h�]+���G%�=�6Kr�Dh�<��%��	gi'vj���Ҏ�j�j�i���&Y�/J�*������kE�X�W���1u�a��b��l	m��L�c��ٷY_;~"(=n�I�-'���Wj�]�zJ�3�J!�`s0h`�ۗ#`��z�okw6�H�i���d씋���G���La1\�-OZ�O:��"�t��9��g�9��B)����!m!�Ւ�߅��\�eXؠ�݉�~q�NY�x���%�wV�!��]�ˋ���}�2�yu,��f��r�d[ڇ�e�E��#ڔ���m�X�V*���v�P�%ec����Nx؍s�[vp�n���6Q����.�&meq��͡e�2�YY�9�lT�9�fL�\��&9��_Ʌ{N�:q�c"�Ѻ� Jh��*͖�ul�tR⾖��=� m-�q�dlw�1�oV[��]w}�^�t�Xd[����m�)n�5x*3��-n���S{]�������&Kn��T����ҳ[u�vy���디��k���wA�Lu:���Õ�;��w��C���Յ�NlȨq�l�ۮ����W����g>��&y��B�*ߚ3)ޢ,����v�{pm�O�R�Q�b����h^��Cyrs�u�"�s_�shzK���ޫ}���)JlE��J�}���^L�1�BnTMx��I�dv*ib[t�R���8�R�zP���Zw+1���Ti��>l
į�q�,XbO$K�� 72�.:"�;R�#p� �1许@YH��l���[�Rmԃ�}٘�w\09W2BM��.�kq��VhGu���`��k�R�B]��2�x������nmi���&�U7���ט�I5:o_F�Tn�}qvl�gxe�=�T=l�';�RT���!�+�xks���o;3F�o��L�7�x]�ݵl8y��X+:V��q���fm��O�GG��h���Ô� .��=	���xvI.��ij���i{UY_.�Q�tL��ue:U֓@]��
[K @�N���v^�|�[z�:�8�e�d������ۗF�������
:�]}�ٍ��]I�h��bPX*/�e��HXv����Cd4��J��ͬ�'=Ȅ{��7��%\�;�k�nWm `��Bp�I��9�X ��X�k{qN�V.���7�o}è��`�J�VK�3oA�1���Lk!N)�k`%y��9��b��r��)����.8��Ӿ�%�gQ���4+�U�����!8�n#�hԴ�'�e+���kmrz�x���Ӡ�sr�iv>�	{Yr�]�E���A�G��Ehx�:ʰ1��gT�f�O�]��z�6#����	c���aQ���W2`�����8��.L��[��-�9���.e��ޏ��]�U�8�M\5�[5c_+%ňM+!�[��W��o��1�׭�> �b��K���8q�Rw�z���E/�WJu�9�	�Ԟ�R���B�Sa��y�[F�q�A�0��:��2�<�+JJ�vlkgJ�e��u��\����۫��IS^����GqN헜g+9Mr��9�ɽ>��̗܂v��D��DM��O�pdm�}iv�w\1ӥ3)9.��j�t�q.�U��I�*h�j��g>�X��ܱ����E
x[�ܸs���*����W��E���<,I�1�E>3*�Q�a��4��O0�ۍ�{qb�9(su.Z���O�*rΛ sS�Y�����j/`Wg�Hކ�m�N��shܦ[���:q�^��d���\v�wҊ�2k�4Z�Β�2�f��T%(s��nQ�+�+o�E*x��+mb�Cq�$q���$��M�˷�D���d)]��Nl��tg*K��V\�B�Y��ԻW!Oj�qv����5�N:�\PI۾��x�=��XZ\��tT�	ɰ����prJxD�3uMՄnQ�m��Ԯ{alY7��r\�(β]�F
�#:��Lj��s�{��;������JM���#��N��q��q��؋7���PǽThݻ�S�Z+�.зi�I]O)��dD&�����m q3"��Yޙx���D؟'N4"�5E�6Q���R�%�D�d�Wx�	�(n�d���UD��P�Q�0ڔ�G���� H ~�����	   ���O� �H$	?���?����������G�?��'�V��!2�f���*��U�\2��os
�n��.)�ZJ�{V���ֆoEJ<ĭᚳ��gICGv:	�K���j63�T�b�fUi��&u��֩,�*9W����rV�hә|�-;9������oy��{�ک����p��<Y�q5w{n�S�Zv�9�EYI���I�`�Gp�lƲ�!ϾZ�@ѵݳ-}f�k:��V�=C���}zhI�M���t��,�u`�qL��e۠h���wה }0*��f�
� ��̆��+�od�h���u�4�Q|j��gT8�U���4A5'��n��f�`��AE���f�z��֧_P���E���%nK� ���b�%�˖�e��& �RPw�)j�2loYL�.n��j�����
�Y�\��g8��[HS&�`��+�4̊�O���j� jԄ*�Z|LN���\�Y�,�`:&���c�+%�hd\^�k�ꑻ Qw�Nm�]�+[˨q+��`׊�����$̥���2f���6�B���Y��n�d��H�b��ov���tT���%�|j��he,=
ItrU����JgUd���WQ�}Y���Y �[k�P�Q6�v����x��M�9-��MU�6��/yP�M�t��v�C�wS�ā�����@1,�ZJQ�Z�eml�D7�+/���̱qv�|00�,X���88p�Ç8Ç0�8p��8p�C�p�Ç0p��8p���N]BGW�M��u҇B"������*k�@91e��vpC����ɔ���i�:�87b���3����7nM��G��zỀ��u��nL��ŵC^�X�>Z򰽤ž�V+Mf͔�.1oM�m�h�rZ�%j(������gH�Ы�'��.�WA��]��eٹAA��v�:�x���.�
���w��[��`����\w��\��Fⷓ԰��P��DS�,%	����Z����q�g~��S\�̇�Ř��� �2J���J��aMtu��Sw�6Uᓛwuݭ����+aޥ���5ϬT��f)vB�s@Ûq�5�ѭ�ݱ�٘6C,�v�'p��ľ�#9�J����3�l&rb����]x΢"��moK�7*uti�v�2�޼gfYBRTf�2sv�]$&�Or�����E>���yp�g��I[��S�$Q��U*�o��X؍U�iF��srL��.��m�v^pt�w^��;6�LkͪY[u ���oO����̓�d�V.���?�:�����4DE�w(���&�T4�`O��&Sb�31 1�,�+�v�bZ����,�Xѡ�7����U����P��镇��vn��a��b�wu,ŘR�e��ͥ�-����<��K�7�5A�Q��S����S��d|/T�&�����kgdOqac��/���y�pZpJ����©�d��:�8= #�8h�c�p�Ç8p�Å8!���8p�Ç0p��8p�Æ�Ç8pǌڝ������hZ����Hl��`�yr�(V�C�$
�M�4�5�[G(K4vP[ib�F�F���(��N�a���i�?Agj��eօ�E�����L�F���	*�{#�J��{�VnȻݸ
�^C�hE,����ӫ)�\��nZ�:\NEv�4l��c8����:�q�6�ͫ�ɪ�jq�O!o/{��N�,>�k�>aٙK����.�r�k#����{�4-;nő�o��5$
�Q�O��靚k41Sasa�eH��yBq��u��ǆ�>b�J�4���8|�l&������e��&N-��^f�����^��A��m�<Z�D;'%�Ϊ���J���^������\A�MśBܺ�G�egq�g��t,� +���޸m[�����Lc��C�0���awTQ�uW�95E��i��\y�����6i�g2��f������ɣf��Be���;�:.�{��WƧ)�X�0�]�X�a�� \�ٔ	����{�\z[�9�Y����%`���[%��E��hF3f��b���Zs�#�x���\3����B@����5�B��r���j��.1x�h��7��K��n��i��M�|��`P�]��v�b �7l����h8�f�/��<����|kc�/��t8���-]�j2�q S�D}Poh<:1���ۛ���My}:�ph��h�c/���h"�إd�Y�m�(�@�W\,WB�&��t�Z�ԭ��+*}X�hӓ��TG.	T9��oWG��4�X(,���n��˼�E3�Zh�'LI�]<ԇ[Yw�u\�������Qqk����D(�G9sV��jt�n�� yҚ|�tGM��2ّ���f������<A��%��w�٠�t�D��G>DVsu�^�a��3�̷e�w[�C�8��&Ή�;�­��me(�����4��!چ6���9�9f��%(gL��J�T$�1ɴ9�s1��ڽw����;�.���,�[���Rh�W�.��gk9R��`��n���6ygR��I�(r�� �O$�������;zscA������+\6S"(����@�o�P��z#��Vvi��Ӑ��m1�pXƥMS,��{y�)B��Ϋ���g�����*�i˛W���!h�X����5I�`Ʃ\�I�j[2�#W-n��++��70zR��F���+�W)��eN�]�hJ����wP�R��L	6]>�Wphα�ʈt*NS�"oR�F��Dl��ݙ\�졄<sVF�[�p�~5��u8�ʋ���K��O-Sxʾ�{�u�3�@�׃��*g�Y���qc���k�'�e�C;��:N�+q�N����)T�*(m�)����}:
��f�j���+;sZ�=�Xe��� *�m��v��`5�y�^�$ۆ�����m�f�U+k�vQM�k�ԭ��:-(�V��]�%�2�s�?�t�Ш��8�rt"���p`&�pd�e,"�we�����G]�I���aݠj��B"�*D�ڳ����l=+_X��򝸓gi��k��X�;o	��}L��z�=�i��^}��*Rb뉗�ujdg9���D���JY�F�<ݮ�ɓx���wʛ��4���M�ڼD#4�H�smUj�Kֳ�k$�Zv�r�YQHr����y�Fh��B�H���pKޡMg,;�Z'�=����Y�+]�gCY��mqK����W�=�Kh%��w�n�K +�#�:�b��?qF����۷YwvEp�y�"�U��hcS�
Y�D��k�R;���;}�v�\���eeWTy�,�E��B��;֙�{��F�N��]ڲbz�dO��2�{�Y%�]�w�ǄN�\0�'FEh�w\��@<HuL>r潲��E�O:n؋or�TF������=;K;���i5Q­��dN�Yן.��.*�oQ��60�h�=��-��/�d��0@�Ww��Wt�JF����z`�j0��\I�.�md�gweD�W����3��MXk��.�Cp��I���	�V�i7:�M�{��x��Y���3�*��\¾�H�*K���GN�D���q��c�;XWr8U�;N��Ԟ����H)�ޓ.�cD�F�f�ҭ�:��t�,ީ1]�y��	�U��ǥB�T����yQ�bL�Mpw���;[i�<V���͢8�ce�u�Sk��fч����ψ��C����Ю��w���͚��F,��-:����tf}[��G7S(g4tb$B:e&T�s��4D��S(���C�hQƮ3ْ�.$�Q˗�zw4C�xV9v��i���ٚ����4M��&ڌ����=g:�Y��W��z��O['']�̃v����ux&Ivjf$���b�=9��eB\���SJ�Y�e]��k��v��xQ�LV���S+�ݶ�ׄ7���=s�!���Jr��ܙ]�71�.V%B���e�m��X)mDG*1
��:sg��]��Q�4�.�*�%��-
C����a.�&�#����
�����I�x�h�9V�􉫸/6����Y�n�@�J������L����K���?�G�MF��$��:U]L����蹈��%ch��A�ظ�s��L���� m=��o�y���n�x�C���	��֤�E��R��Ѷ�˘�8�Vӧ�� ��c�h���%6w�Y�dcB3�L.�nӝR��y����-ȡ�F���iy�v��hV��j���Czy�]�]��A����Ǭ�/�[�C\���|>���9�GQ������&7���K�λ_Zi��e��7ٹO�L�ުS�ݛ�*�].����Y�w�et�xI +++q��_^��r��O	}f�ٶ�r�:
��](^0��ba�C;��2�yc'Yݼt��Fc�*�R�W#}X�e�3/��(��W��/F��i����a�XON�kц��GN���%ɖM�(�]�ɫ
��YZ��t���Y9�*p�r���\	��K<l�&=ʎ��'hoA�[���^miJٗ/r^�F��V�`LP�b��d}�݊� ��F��p� Lh�7����=g� AE̑V�gvm�-:�@F^wj졫��&<`�ՄڮW���r�+#�Q)u�6��,\�&��h��w�Җ�gw5��/x���<�h�(h�Ь�P����Ϙ�a�e�3% ������ �S;�ՍC�L�9����0V0�*;���dp�i�]\r�:��\�n�ִYMҷ5�����v����ڧ�1ڹx��ؑ�R��*�_s�P;j��@���D��ٹ@�N�K/zڪ����|~w���>�v��[	EXt�sz��"��3eq�ottvs捘-ʗ�D}�:AQ6�.3�6xa7}[y�/*J��n|
�:c8�oIʠ�kzv�4��݆͗@�2��FY�2!N�C.g6�E��������l�f+�/���%�J�=.�,`��H�`ʈ��c>f�=�v��B��bvvH��2�5rk���Z�XOx��$�/R�တ�:��iغs �J�/c&1l��h�.���h4ݩ�Z���N���O�d�;�gb�`��ïI�5�7�����jh����o�齦�(�tz�e�.g>�m81S~t e�⫝��2r�*�\*@r���ǜ<
��Ę]�����s��J�:��ox���P��~զ+�o_�Mvu778���0��{�Q�Z*�ӎ�@�u�S0+�E�,�5���L���ƟQ�u��;�	�o�m�c3��j��^��5�EU�T�t{S�&
��%b�{|O:�*�yA�`��Щ���d�č��:mp �ʭ<0�̗���ә�$s�b��G���ى�8�λ�7>��F���ZCk&|���`e�:U؄t[��X�,ٴCBY��VԂ��u�C���M��\�VV�+Qcl��ݦ�D(�;2g!h��)�N��ǐ�EIM�s�������n�����ŰI0��˕vq2�n�v��0N�����WAvJ�³9E,å�!�]�(��os塛%���*�9�e�&:�9��=���ާ�K����]LZb���z�e�g {^�נ�Y�Y��w��MX��Wf=��a�u��:�t�����{��r�!�S��'��MM.�p���)��k����o$��}}0��F{���0�s�6�WR[v��&�['S9�ٴ�	+Xx�O���ҷIQ���m���	Ye���7�_��Mh䐚9I���ѡ]Î�ho<A(m�U,0sE�-CÕ�Y:�*����4m	���}Y4�����c0;꜖X�9�Y]��Z����l�(��ρv0;���X�6�ev�����Ȉ�"�V�[¦�X�V{`���ˈ�Z+��nN��w��k��)�� 5}.��;"o-K�c2��w?�[��(y<�L8����w��N��b����(�*h�]KP�A����	e�mحk#�4��.Wd��&�tl^�&,r-�]V�ф���ܧ�mN���� =d�8�}1�]�^J2�!{��
��f�Ih�u�P�P���N�f��d�;�MլZ.��v^�*^*��
3z]\���huy�W1��R�E�i֫t�A���0"8ܼ#�/U��I����ufQ�],��Fu%\͕Av���a���^�J�k��9�vNt�;�_�o*F��'$�ג���m����7S���q���,E5+t'|�6)#N�_]'���e��aG���/(���ȕ��\ׁ�Ӕ{��;�K%�u;8�,���3�b�-�[b�c�Wc2�l5K-��bDջ����R����E=J��e�X�1K�qD͋5"���]cy3ˮ�=��[W)�hF�X���25r֥�6�F���c;�&�93G�;[��J�N�A�� tw����	�a�Od2fX]ScKf�Ճ�}�KO=�)��L���K�ښ�X�>ul$0l�I��@�ɻҴ��ɣ%f+t��A�Uz��6~����n���	�q�
���D��ދN�����.X�.��=[���ޔ~�y�C(T�ͤ.��:��&�����c_vk<Q7���/eA:�p�iM=ʄl���]A+ٹ��<��G�7��N�՛Wn��Iiz[="���UToQ��N֩�}7euNy��5e=C ����8���H��rq(�;G�4�s3��s��;i���%�e�ңJ���K�E��MԘ-�]��e�ك\Z�.���G{
��h-r����*��˱pcp*Ћ�s8vk�̳�i��e�}��nQ��Wi�'��2�,���VNٿl6��W�˸�f���9�z����^����X�7$��2���������.mn��N��}���Q���Ǔo:u��wkj�V�R�
p���6�u�-��I���틅��;�E�{��G�.G��JC�u�N�]V(����r�R�|*9�c,ڛ[A]��ɱ=w{:�>������~$ ?����~��?���?�������C;�9���A��������c��BU�s�ٻ����gt�����5��ue�Z�_Mw&�����ġo8�g���g_�2��\����\xS3uVfty����W��(�4m�Uo��!��2g{������}afb�Akk�������wueE�|������R����+�g�S[�Jj�z�4#���t�uV�x5���2�@]#��[�ga�t]}a΀�)�\܏F������Z���� �7j�h�.غ}�T�[�ζ�ɗW�N�3���̺���ɏ��,,��|�^ŕxi��lꗄ�0����!�2Mݵz(5��tK8�#��sc���e��#w��/ �Y@J���Ly[���e�[w�.r�ؖ��z(�4�LCn (�h]*]�O58�\h�[,���gۃq�7*�-8��7���;�,�Bdu:�x�P��w���x?	cS��@��b���k\*���x������u�q%����e���5��Qӕ�S.�Y��}a�_J��*⭐uh�*�����*�u��8�a���Bα���e�R��Vfӽ�C5�,q�{�.f�y���|ը�4H�+���9��b�e�v����}Z3&�)�r�9VE3���fq����j��c�0�=ռ'1qUK�vNv��d��x�g�=���K���:�7cٱ�M�(�Ƥ�m{�5��ǟ_;�Ģ��Hɓh�7�ȥ�����R�,�2m©��ZRD��QI�b[Ǐ��|~?t�D�=4�����%�R����D��񼴬�D�I�u�35w����������
Ƞ�3\���JY}07P�J=]�Ŷ*��a����p�s%��Ǵ��w��_<�
�S\\���rhe旕�Ae�[��ah����$zzz�"Z�
*���j���ELMJ�(򢰔�(���^��^�p�.S����%��Q��\��޹���"2���a��Y���S��+'BU��ȼ�ΰ"��e�����,�����״�=2�m�������zg�m�**��"ȤW���D������В��+�>v骪�e6��'�ׇd"�94J�"g=��y�Ǟ7#A
�4��J2���M Hd|A���(�\���w�8N���%�Ґv��e+Y�kb��x ��8j�9R��촦����Fɩ}�Nh�h��-[V�P[��7�q��"?k�'�5s��7�/f��	�{k[�\�/�3��柷����X�J�u%=��۞��g:됱Ԅy����{�u���7����7���E�L{�m�3��r���kU���p:���z���.�ԶQ��m����q�F�N줳������d�h���B� �׆_�̀�.�11��^�����_�~A����6�P�9=���꩹�٩`��A{N���� Q2~:��iJ���Q��|��]���Id�'���熡��OH|�~Q_|�]y^�5��|��$�״�=�Ql��>�7���+}�\7�7��I���)O��-$`�Uu��j4�Oi�o���#�u=&�z�t5@��=�ſ@�U�����xq|;���ָ��ڙ�M�emS���ӓ�zsV�۹��=L"����*5��0믞�e��-�;$X����NV��馲ˬ���r�-s��,Y]K�b��֪���e�u�z��%�T���}N�uYS��+���Y��;�.Sq��C���݂�j���C)ou�|��U�;.�r1W��P�'ޠ|��,:�����5�j���ћ���{x���/l�+����4�eTTc5s�l�X/�����^{��#,���=��ڼ0.m�#){�<�?I�Q��VW�F�O[h�ޠzO�3��6��4����7W�C����^�^�-�P;=���5��R϶lϦ0���=k���J�UČ�4n��S�bbm�otzsFi�������l�Rz���V|��K�&��vq�W�8xn����Uk�f�]v��"�B+0�S'w�*.S�g�*i�_9c���}U�z��3�	�W��k{�г�c�z*��}�=�SP�o=<v��/o�E���{=Q}g��y]O��R������5�\�Ǟ��>�=�3�==��W�<~wB�m�Ի�/��=Gύ�����w*^�]�t3�OW�s�l�^O�jN�����#}4j�YYLM��>�M����Mqm�u���8�D�A��+o
*�{�k��_��aXw��ԕ��!z�]��c��\���H	J�cc_H�u�Y�ۦ�;�SRwwA���=�9묛FS�Z�@�w��h�hcn�uN��Z��&�Ruѯ֪i��S?s�6/��xj�����'�����B6�+�#�x���e�N=�ϵ{릭�@F�/~k�v/L5�^�y�3U�\Q�U,�Pz�/=�q"�2=�4o2��"���~U	��N�oމf��%��^��o�V��YT�%�61pe��5}�fP��i�h��o��_-��^;�+,i'9`���8���h��{�^ԛS*��?�;�^�L���>�W�>�D��{{&��Q���G�_ܡmS�E/|:��1aS��`k �ᵩD��=\}C:=��T��t���~�����= ȫcMM��L.F�{cE�;�wʸ�@�7�7<�籷]�(��oW�}�%�ߊbǳ�ʿ�w�1�����T�&��!�~�ME���O{Ծ}������_������-�+`��/+g�G��C���{>X��1{��Y�{��kZZ�ܴ1�<���ɥ��\<fU��/~�Y�!�j��h:}{{2�0aWc�ޱ�-�ۍm�S9'vu��9p�XX�T�w+��tʹ7x���g"�XF�[q�O2�ʍV���a��o�������7�W4čf%v�C��)��:{٘^��Z떵S�{��§\[ώ�tU��N�/w#ԡ��:��{��:��*�_u%k�J¥T�yCjʯ��k�r	׳�x��y��[NR�ez�/D�vЍI_K�R�r���ۖV^�&�zj��O�M�~�^uչA�Ŏ�_\��7���^��g����������	��ֹDQ�E0�ђx-��]�K���ؽ���~����[��a��v[�԰_$	�+��ml���l�G�z�Uj^uҹ������)�޿�h��'ok����]g�w���bcȄ6ͰE�#�}�of��ŰO�����>�W^��2�@��L���3�z��qWr�0z�]'�X��Y���S����^[Z׫LU�^V�Y��[|���.������AV�ʮ�-��������g�\I�3�6�^��N{!��}�ilD�F]\�m���c�J�^�Hz�ob";ݱ�ք � �	��k��v���K����Yf��q]���.Kv�X�y������$��D@�t����u�x}��{׈`3�fa=#�(n ���셲�8u�!�\;v�q����.���]��l����^E�X�T�Z��׽�m��WN�L�~����fW��հƍ�I2��l/S�������}I�����7WĊ���f�[3�O˪a~P���u잣[�J~UZX�u+��S⌞��'�U zC��)��þnY�}��g��{}G�VV��y���lWTm{���.{��hdĺHx��_�G4�߼��z�kݧ��Gf��s�Vf8N^c�5�����{,R�0׳��,f�߫ݵ'�}���8Ž��x#;by�߫�m#�A�;a�ܙ+�D�+s��-��_J��ˌ^����ߨ`����k�{��N�����99`�K���|=���7_�yRÅ��;ݶM'��^����w�Ls�q����F��({��̨j+�eeuǚu�0���a�g�Gџm�=�-��{��y0܆��}��gG��Ca|[�t�cmZ3I���i��,�ѫG'�8r�t��/^�i�kgN�Nԛ��X�q#:��$߇�TC�4[��k}��z�-��5�����㢇'NR9ڦ-p.k�Ne����^�������m�3$��d���mtޢ�U�4����:\ܐ�En)�g�y����zC��ڊ�U���(�y��N�-�=��|H|L��=TQl��*���4��{Kٵ�\3�V��;�0�l�����
�9�����j%{j���g����T�������ٜ���Kr��A��NU𔽻k=��N��Ng�u�4�����e(saݣ� �N��K��S�{�������\�V�_R�K�|�y��R�^�B���ۺ��-�fxZ~�=�y��'M�{Q�×��O������?U��~��^�~^�ѻ����{����(B~R�*ܤf�/���f[�"�No�9z}:zN�'>�W���yFר�����{�]zk����Ƴ�*�y�����1���3"���H��DJ���Jz�+ݳޝw;��;h��>�P���WVr�!fG�ÁzFNV����X߫�'�;��	M�(�fݏz����Ҽ5*�C�^:�oEFﲅ�<	��r�.����O�t)oU���%L٘�l�{t.�Bc�� ^�p�;���A�O������:�ܼ�eΩ�V^�3-˝���of��]�+�7�ô�3��ǬS+H���K�_1,fY����j?V/Ojq�<�r�^�Q�W���)F�y���K�@��C����7�M���:�t�����ۅ5q#�����Ez�YU����Fp<��<�޾2���-X���㷣(����N��K��^�<Χ��]��)�\_N�ʤϽ����u�٩:�T�,�~��T�����z�Wb��B��w���f����^S��o���C�-*zE��*���3/M>d_2;X����n�7~��o��W�������d���-�uzM�xO��zύ�W)�WM�8Y/�P�~��¨��熈I�t�wdgw�����+2�ǟ�WÆ�nWG��J��}��H�oz�0//G��Lfm�c~#��t��y,X)��S9yG���i���R�^������3S��?/�Պ�{��E�ֆ�p�Z�n'O��xm(UŚ�;�m�Q˗�_yN�=˞'�r<A�k�[��6��ffA	{;^�T��e�u�?d����/���F6F�S����Xu3`1�úEL!�ν���	�x��hK���{Ғwt�rA�.�O��9["b��w6�^�ѳ���M���(r���eE[;�ׅG*�_��a�ͧ(�2�`���jk�ٽ��Fe�47{�%hN�>n�;��8Xu��j��C�z�ڎ<���U���JI�{�*���>^�/|�
��gMjk�uV��o��׼|��[��W�j��?JK=��6�,��f�)�֜��ʗ{{���Vj=�\tCU�������Y�Y�-��V���9<���mG��^^���y<���-�{��,B[C�[���<��+=Xt*�'tW�8H�[_F�������Z�����@�xǽ��#m��{ �����0�^���68��K@�_�6��e�����q׿W!6nD���f/Ut��&0Z8[p����O������7g�[+�I�^p0��S/u�wz�{<�G̼�o�뇫�>�?2}6��2�-�oGJǕh�C�W7���܈vi��9:�٭Ӹ��Q�[���͵z��� ����)���-��eͧ.��y6�`*�3�xv^�x�tYٙ������j+�׭�T&�\����R��L��2����aM��WC���yE�#{^>ywv.���	]&f���ܭ�}*��O.��eA ��@���O��ٲ:'��n��#~��zw$�J{�잛�����N��Z��|�������/U����|B������������wޕ��V�.�)v��6��u��ČQY>���)���mN��T�.$&8���Wj8��>�e{����'��ح����W�<�{����T1�V��Ȭ���^�����:H%&���:JY)z��~�ɠ��m{���y���X/���x�z:��=�J�j���{�'r��W׾B�Aw��f�x_�:e��K���	�8�5x�#�t����7�.U�.�"�l�[1c@��gyt�����|�rv�V�#)�u������yz5����y�2�P���_(�6�����l��y�xŷ�v{���<=�;��*V��u��NF�t�
�����t�Ɂ��T`�y�)H^��W��k�}ަ퇀 �g^���}O:�!�%x���o}u+W�]������ M!e���x���'����\U��qc����4��:e(��sq����2t��b�������*L�Kgj(�*Q#�v�u-Ͻ�*
}�X�m�W�rN3�B�S6�#F�˝]�����R�[�r��F��TUg��e��#o	�A��{����y�~�[>5=<~�e����J��*Wey�eDn+6�N�z`9z�ь�g���{��||�fC�H]^�WP5v�=�������+;��Wg�_tu�}^��1�=��|<�C�傰��a�g\�}���������PUD���q��=U�oٴ|��ݯ!��^�Х;���}��w�0�W�y@� G�fI�y�=ޑ����uq@ގ��?wv�fsIE6��ci\)���yH9���~��D��E����o�zj�n{�x�Oc��Sj�T�u,R�L����^y���������	IR��$����v9����w�ȹ[�ь<+,� ����'{���U�U��/���a���2d����3A��Wֳv����`'��[u[��6��H��c�]�MТVc�*4�����L��{�W��s(�|�y��;�\ݝh]=���f"J���6��s��n���"$*�{Sa���.	��`s���_.�!5s���WD�в�N�K��aˬ�r�\I��e����Nu�3��i.6NVƷ]�vm�&u��U&<Y4A� ��;n�.�p����o&'(�w&ǗRh���ň/Hu�L
�]��	��9���N�nl�\/\�7��Ë��7oc}@�}#ŮQdnU)�JV�g���`������^S{
k��e8w6�kU�j��ZM6lD&)Ea���;P��Y7�u[�a�j����ͣU���^f���
-[���3z�ܼ�{a�gp��Ќ�#��.��3ovu���0I;��k:F��Y�9��X�5j�AUĢ/)�Efow	 ቃ�M/x����^�*i�>���+F����M��՝{Z�b�����oK�x������n4Uk�sg��X_`��`F�PVt�͜)L�kY�c���lT��Z���W�H���Ydnћ���m�NќՑu�{�z��jdQ�\<QF�c#����B0���o�)Nȅv�SxU�����m`�7'Q��Vİ����.�mR���w���V�%{O,e�?�Q�_�+��J�n�|��rDI���d�xSM�0Y�GQST��x��{W�n�Y]0s1ouA��FݗԲ��S'M��=�c�q�b|Am38o��R}a;��蝁8��C��V2_����[c�u(�-�t�CiQM�)	Go���-J�x�&ᷱei�����5[�W�;��o\gtcI��5s�h�a5���%���.��gm�:v��0k��P�+2v�Ż����_^�s��Է7��jÍ;�BU��S��*��H�
���fZn[����
/ MΫ�Y�%�U�[��}��Y�ð��YϖuME汊�����*�j�9�7m]1��e�⌫9k��kj�9���)��eGz�q�۬P�={���� k���t"�;��d��S2L�(���}��e3j������͇be3���(sy�]v���DS��r�K�%_v�c�S0�Q[p������JYImۭ����wp�Ϝ�W���o�.Ծ���ܚ�ki'�Ϡ���u�Ȉ�0�d�j�u�-��DN��9ö�醺-h����H],��(d�r1�l$[�5�(2.^��ػ����ȥR�L�Oj��$ou]�!vk7Cu�PR����;�j>}����q�N��튻/��lh�S��hI�ۤ�MbUۙ�J�y�s-uaw�a��<V�X�q�p�ZMAx8�ևie���Bu��r�~]���wC�[���H�i}�+��#�ˈ�e��[TG����������}�_q��a�M�˅9(��;�B��'=��;	��g�<�@�Q(�BD�������ڑ(H6���%�rF���Q�E�Π�X������l~/;h���?�d}�r�y��`�f�;�7�������uԭ�ت$k�n\�U;<G��>>?Դ����"��նƢ�4�J�T�/"�!Nt#k��bUy��I��I9�I	H3��W(�z2��RR�A�g��/<[V�%�K�T�ٺ]H)��'���� �(�<�+�Ј��E#1�c3�{`�bT���Y�{H�h��:T�\奙�9����}��z�{x|��$D�H-\��JV���ʃ���SG�x�L���>��2�S�'d�4/���f�$�}{D܉\�=����Hz-AB���U=�!�e����:�zJY!Ջ��L������
ٞd@�Q��y��{A&��>I�ǽ��D25���vp��-,���z}^n�v�d{�I�d��i�#^�0�6�ʢ��/a�i�D�_R�d����e�ַ8��:��U����;��oc��GyT��u֬d%�8Lcv�t����.��0�i�a�UuW]���y��y#�~��Dw�YI�����Pi\�#��MQ<D���^�l�5�eO/�!�|��;'#��7�k�N67|�"X��V�Xa�RA��g;0#)�#z�Ӌ*2����|��J�}����L�a^������VE�n�7 �!�M�Q&T��GK�{�\&�p�,�`ڜ��o䜁,��
Rh6�>�A��hwl[ɀ$w1n,�x��}XL��z;)��]�~v#!��[8���<o�o���x����o���{�G��.*��>�9�g���P���ZSP��Up��	���X��Af��2()q�χ�k3�b���5G���J7$=�t��V���Y�[(�e���ð���WE�NI|~�`�j��dl�;�󽮼���Θ�a�p�kh�t�NH��n�>Lۑ)�������J|�z7P���ə��p���?{����؁>�(p��8B���\#�g"�ծ�(/K��|�����"���ɹ�̺��鍙(kΉA��6y�y�!�F0����Փ�wһ>�+�����TG�$���q�r���0�ܢ�~j跚��4�B���W�\=�]z9 ���˔ԃ=2�S<c�U3��*��8�n?^�e��\�i�t���F䩇�eJ��}y�%Kb}�:�;J��T^�����r���^ٙ�\���q�=����`��=9^��['���L�����F��;��1��sb90'�l����c��щ����&��O�Zk^�Q�|��3�XR1Q>�A\��-�:�Ov�8���٣�D�����N0��vv5�d�=����1o��ke0rC���A���y�M�����#���K{f��T9;�ù�v�U���d,eU�x����ڋg���H��OD�𝾨� ��4o栻�a�.2jW���Ca��Ǿ[�n*[�f &L(`5*H݊��66�����[\"�\��b}�����^���*{���SZ�k��	{���0��>y�����o��_�4��љ��W)i���),A���Ѥb���)��};K���?�����ju	}���)�,7��&�� �nzl�Af��'#����vN�������9�䕜��c�y���,3�~�P�&�`ڞ��=s�V��#��G�\���=�y{��������.oL_���тvZ6
�#�R?S-=V-�p.�Ӓ\	�mqW�a���K��ܸ�����Yd���E��w�h��&ѫð�j��v9K佇w���wh��T5��������+eM�K��9sU��d���)g'B�	��6K͢��3�Â�o3��2d%�p�U�g@���5դk0v��P�~?���m�r�j�ľ��p���g�#,EO37�c��(�.<�i���-�v�����a8z��q�fMk�C���1nr'�<?d��k�����0�G�n�?d	�Pފ�����E��Z\	c�X�n��U�l�a�F��a�ة>���� ���P�y�ǔW5|s���x��5V��.������Y���#��{Ɔ��4Op2O��?0C�a�>�eTV|���㲳6!�gkQ�\�L+P-�_��Sf���Bkj`8$��NB�W��M�U�D���g���	�v�e1��f�q��w�1g�ii0������[��_#�Ŏ8A���;ε^$�	&�s�����-� �tǣ��C�o��ǎi���>8��D��`��+�Ri?fF�'i{�_�ނm܈�$p��"<���a��PB��$=W��&+s�J�}뜋�^�1�۞�dP�t:�C��G���N.�T(����3�{>��l�����TCVNu;�\��)Ne��o	+p��l�=7ʪb��D�+�h�)CD��L�����j7!g�M���<5�تMq���Z���(S�J��}U�O*�$�k�,S��Q�s���v�q}X��ગm��E�2�!�A������x�rm��{�2Ġ�Z�][���
�u��n��_`Aa��=+xڼ;������ ;��s�v�ρ� ��lgn��r�~H|5/�V��@�nC�
&q����[" ��U'��	u�Ue����a��j��oei��-�1x��o��ҿ��O�����$�5�/|6��+�}��6��uć�h;�Wν��U��[[wQ�}΃�yK��,[n��}���ߓ�7֦6��]�R��~���Q�χ�K��H�1z�a�ژ���S�`J��o�ųk�%�w�'�ޘ������N��y״�*��g ĩ�"�"�?z�T��z�B7���<�8IR=��B��q��	����͟c�?�i@qKN�`�W�oN��7�B��-���*B_z$ ���yt��;u1�~�R�����cު�����l�GMðV�X=7�Y̩gDlH�&��G�O.>�p�4,�o��f�N�}�W!�c�s�l��\�/��p�=��J����H7o������f�3����N#!�:%H>�P�V��--���\����8�BeBC�Ԥ�["�0�{��6��
}Ro��0i��LP���a�][-T���-|��F�9�?:�C��W�r�l��V��B���C'+a^n�z6��ݹ[?��8�~��+�J�4Э>��i����&��S�Cb�C��1uoo K��;�7vUޚ�Y���۹��Qm5��!S��k[�|�6���˽)���N�T>=�Z���,�m��0�y�T�c,�yȏ_��O��) ��w�½7[�7��,��`lA`��,EH/OX˫�x:�FC���o`_�u>9�o�o�_t��^��op����B�����"R�P�p�C��cK�}&7���ud0�8O���ufqYU�كYֽ%�nu�B�U<~,o��q���	�;�<�<0y�P?�Q��Ȝ�}.eW:�p7r��7ݽ�n0��B#iz�=���<����7�-p��`�
��d0T ���n҃=��4�{k���bkԸ����SJ�%�~���R�)�5�T�G���MI�m��fF=^B���O���t��u9	��z~��j���"{8
��5*H.4�fef��(�ȗ]��!e�/a����20OD(85�K��-�C�];����)]lpNŸ'�#�H������{����������S���?��e
�~�?x*ŋ���!���o����LGt�;�uoL^����HC��[9�^�k�<o�7�Q��,23�늠�6�4-�S���'�~��7%�����"�#G)�l�	��r�8���E�� �q��-�Æ�Lg�o�Y���M�"�=T�����6��l���+rw+��sY�I��:듅8jh��v ������r(�]M�yB5=yv��<��R�w{p�G�=&a�v������r�"�O�n+���W�ۭ]��ѝׂ��C���AD H�A��͊����%
��.Oy@�g�q�3�w1�g��}B��M[����迏�$�7���c�ӗ����JT�B]"��][��uz���N�=�S6�c�R���Fxnou^elt�y��/�F��	�$�m�����2��u����Q�~Y#�<�o��]ng���mf���*��h=�(>�����9�@vІ![SP����\v}��hR�=yzy��u���վ�/r��ɴ��>'#��cN��?1�@=Ƥ���b���'J�<b��������_�^��[��I��a���WU���b6�`A�'�#��P�4���Ge��޷2{NQ�8Ǜ���p9A�?�W��Jg�l�� 3,�r��t:V[M@�E)���wD:���B�Ty�na���[M��*�N$=�ڏ��xap�.�{�X�uWv�wx[�Htf�����5/�f����Go������8�Å��߶���	��1�E��)~-��0�$�2�����l�}�^�����̞wy�7�?l��}o��0�)f�kx��Ǚ��Q�&����+v���|"�����5Y�/	+)��tS�tʓu��n��AG��//��9{�mqo:��i�jӫ�Ƞ���\۴�
��i�	L�={��Y��^-1�ob���Y��hL�Sk�q�{���8?��D�{�x��G��{��	K���/|c�����b����o���_l���$�����X*�}]T�u@��z����n��\�l��!ŧ��Zj��k!ߘ��5�ɜ
G��������׌����}�t��=]۱�+f�/�Xgc>��� T;M^��=��c�9%_�$Dnxo�5��d�Tr��뷰�<�i��h�\�ɰ���ѳ��?�2��`[�ہqa�*��������p罁���Vf��}*UDe�Kf,o��
�S�����f�xV1��%�G�Q��]U���J�#��� �n%t��N�}%�E�b:��a�)���nF�\�=0f-�L�o��M[n6��r�agҫ�}�`
=!����}�Aml�����!�Nw'7u�U�����1j�t�r�����
���#C��_'��� ������wu��v���Xf��k�m��u��b�ځv���rٮN�+����~M"X�kAaՂ��>O=3"�����B��266)͢�^Xş)��f$�@1�t:�n�|�X;�/��2���m#���R]����;�\���
2�XTﬡ�WDQXXi9fΠD���{P�3�u��l�mn�)a����DCs.ڬVS]m����:b�.d��N�E������
�*����x/)S��8���[��Rs8��+f�&-�Z�SK>�]��X����|`Nx�xx�9{����{ޅЩ���?@�*�ҡ��ѷڬcϜ��;=O���b�G��*�W�B��M/�����1�;_whRA��&ᏨÆ�m�����:-kvz�KB)�����3�Ӫ�HoD[1I�]GE��2���B��
A�\����LG͖�sS�������n�ڧju��(�	�B��fc�h��}# �_i�e�0"�D�Ϡe㉟���q���ʯNU��Ŕ2��.���`���A m�E4�b���;5�|
�2"�R* 5��˅S�sY��������||.�4�v���v[b�K�yA��}r��꜒���ȼܫ癕�C�����=�>�!�K'�$h=�z}�U��Z_m�FE��A��)b;�OCv����ES����}���!�L<�zy�6�����Y�8�e,BM��n����)ǳ��=�+Y��D ��=�Cz%{�B���6�����o��L��&N4kҀ9�hoIP�I�I�;κ:�'�u�㰞x�]{�Z�7��-���'"�-;vs�����60����Ƥ����0�W��q3U۫n���J9r�W&�nd5BEB��ge7�I���u����yl�ldq���[��o(��Rel܏6���ވB%�<�K1.�}�l*M��w8�V��SK����U�%�����B�W܇Ggv���
��-iz���I�/�Y��T�E�����	�  � ����$���M����X�'.L|�Re�#5��t�4�8zo��s*Y�bE18���#V���������ܗ�����"V�[�]�\u-4�%���VTX���ȥ�e�����̛�L7ˏ��,P_��09l��E�[nH��]]1�q���9P��)=
���d����4�-SƐgH)���Уb��'c��^+�@Q-���Iңu�]y�2]�\�fllYڡ7Z��ԟ��q�qX�9��9�p�·�6
�H/OX۫�x:�FCϝ;�إ�f������k�z�W"�l�r�[t�߲�:����Bä���jLip|Lo��[�yz%���3����r�<ǫm��������M�ʫ�u�B�8  �D
A�ѡ�R/#��J5�����<]��k�x��s��Ј��M���c�H[r�����Q}�L*4J�g�1k�3p[��U�@~�"��Vq϶��R�V!nנ9:����C*��:0�_x��o�+�r�nm���g�n�=0���������8�5[����"o8
�O,0���za6@�ȼ����ǁ���7<Zڢ}�D����ٹ��v�v�7\��`���x�����DR*Tcc�c,��7�v�
�KzV2P�̧�|�gQ�6�s�T���䙜2�.�D���:��YO	�
u왗>o9�����|��| ��  A(r�w)܈���ȫ����>�o�S��ដ�rygV�7�>�Pts�1�Sl�1��w����)[^o�[z���f��W�n��z#�V@q|����S��L�\��r�K?J�,_>)��m�ɧ1֭a��d�OSռj��0�?y
��N�C�ʭ��ڭ�k�<��O�>������2?Y�A��Q�<e�ɺ�^�{Ռn���t�����ȾSP��������N�����8I튞�����b�w��{%\k4�C��T�
�{��b�����L��i���\;M[��{+����z"=�=,Q�m�ˬ���pN s��>�%ss����.H�޷m�3l��uO�^~��i1t�טwՓ��鍒@�t����-e���އ�����[v�tµ�q�cw����j��QJ����y��[�9����ds٨B�u���	�P�W�P�(mMCワ�q�4�����l�/c���޵����j��I�9Oq���9`)�c������&!�X��c��b~j�n\kb���+�f�Ҽ��_�3��*0y�Xj���uQ��&#t�Rt6 � $ �<*�u�!����8�5p�ý5�5�S��YZM��2����Yܑ}f;�3��UW�t�l��Y㢙S����<X�%v@���N};7��u7��/�'X�n�������7v�=��jS:L�KoUGl�pX��j�mMy;ݶ���2�{x婘u�ouBK}�Uإ��Vp�;ӕ�u9	�-���Ƣ�Ld���j�>���w�7C�E׷������b ��kx'g6��z�7�+�m�ƺ�-�����#As���y�P T쬔���Y;z��P�଼�O���]��>�5v�N�;Mdͧ�b
M�����]��l���[u�d�1�;v̏ӹ2
C���D�]���z�� ��Bk�{���jՅ�pB�}��e��\%���~��D��&�8�(e�Yg3��;l��.^L�i�`���_]8�m��z�a<�54��6������+�d�$���ܓ�W���k�&�}��c�35��E�>VҬ
�z����K�dbմ3/%�v$���9q���zv��u�S��(�`�Z�e�(�0kAC�#i[�����,⡭��3zF��aY��/��Z*F+-��b��nu����:��4�ś�'^��\�Ck���JL��Ty�=��(B��U�����s;"6
ip�fop3)��f`�t���Cje�;�^�Ѳ+`\��������嚟>����Dsn��|O+�E��q����\���VZǵ�.�Q���9{��<o2�Ŕz�T�|��G��Pz�r���ō��]�>��u�ton?��Ԩ�;����r8.�-N1�:Z65���7��������C��'��fź�a����4U�TGG2�������Q�R.�ÆLY[Sz�+�]䷝�E�&��
��]m�Y{P�t�=uwɖ����vC=��n�j-��i5 �ʹ����^��\�q�����`��Su�u>A{�N��f�{��Bam�������ʒ�1i�5�P��%���b�]��d��s�3VX��ę!�2�pݦv���62���sD�������	G�O���no]��w��w\P"lm��ڇXpjGc�2���B�婄��}.�هU�`n����1VֆYr�����t�1����3{��ޗpdH�ޤ>�H��_v��4���-��r	Be���tfJ;�v�v�����,\��Q=Y�I/�b�ZlU�[�*�l��,��ת��8�Z�����m�F1�h�����z�v���OG\�=�ςC���5'caZ�#�^�ή?m7o8��X�J<Z5w��S�1�Q�����[ܑ�-�R�v��*�+��l��u�9�Ƌ��Sh�l�nCF����ǚo�<�NRB��>�:u��X�/����ٽ�����P7M֌u2�U��oed�ǰE���uF������2��L 7o.�#MYm���i��{E~�#SWHH���Ԫ���Qx1-�C2|�Q�^�P�?�����D�$7�s��D��&�鄊u��t$C܏9�3��<�ْ����kυ�<�T���������u���ךX^��y�=��q��(��چd�v��r�"�ן>�PXѐ6.��ϱ�u$ʏ�TQJ�$WW�:$y�J���טto�ޑ.d���1H�
��Fљ�_�g�_w�s%N�R:%���y�Jg�Qji��Z�"�nG��+F�ח�Q���A=�L�(LDB�Ū�{zȏyUQD�âz���*5/*�P�I(XTL8ĽD�ԫI�˒B�hF��ob_طW^]�2�����go�f_����^v�D����y��TG�K�6����&�^6]�w�ԩ5WK�&��_iW^�&p�V�iW��ra�޳�^��=-ֺUY$���;ڮ�`��D/�ۧ��$��y"�LAq�"/�
$��g����|�#����=�#�~�̨�~dt%-�SyΨU�v��$�V"��,x1��^w<���}h��O/yv�BEcl�F�k���9��_vM����8G��=�s4����_��O���mfU=&����a��W+n�EX�S��@R��@ �)� $=��
 ��'�p�| �Xqֵ���?Ęґta�r���p:�3���]__e)����~��{�$O��t�>�v�C���Bw���G�p�G{ʁ��d'
j���9�E{�"F�ӟE\͙w���r�xp$f��\���2_������q�����ͳ&�r�F)8<��w�Q�%�}��z'�5�U��(���&&�vK�9����iW8zL�.Lr���䏛꩷�����%��Z�_��Ca�S-a�ʾ|է�$�<ă�xCܲ�Ù�=4�7��^]�k�������X���X��yZ8u�loVG_�dh6L��H�� �Q���;W���ϰ+�����.��<��o"�t���yK�~�P�5{��\��9�5[]OB�3׾H��xl�@xMx�nEͳ;հ������b���y��b�;��О��n�Wa��[<�Ay3�mo
b���Л�����G�쟏E��᳟)�e��;(��z&����"K���#0Nנw�Į�����6`��B��F4GyL��O����ޱ��YӨ����f��.9W��[.�:�b�h���5(އ�/���'��:R�ٯ���]G�ב��-�i�t�[��î_$�/7H�j��u@޻&����׵�c:9E�ad��5��$��`p�5:۱BmGDQ8�ݾ��"(lU����8�e��|#�H P@�@G���^�{�^��8�D�R"@H� � 	��Ȍ����Uk�c�l%�GP�l'���%V#`�a���Ha������렂0����y�>�ɧ�Ԛ�=Ǘ\�����!��#��L� U�z�~`��L�<�(D��I�9盯���v\�=��b�-��z��Sf�:P�ژ��.�� ���-�õ�8��a�A�bdl.3Ƹ�WB�SKH�	;P/�l+Q5�[��A�v"т����ċ.��{o��8�AtF��T] ��!î�F����=#�t�<��r+/WE�'�N��J��Y���F���N����\ ���p�� �osl��eח
G-n��`�^KS��N�e���u�>`wQ��yp���͎8 �T"O�a1�� ���#'����3��ʢ�gi2d����q��m��摋J���U1Ah��t���i�g����O��޼;5sFnj��=ƼT���_�� H��3c��@�r�iT�/	�w�Xf��D)m�;��o��y���r<�c���@]{����w9�#l�9�-�1c����Pb�i_�C�Yq����|���K75��W~��iM����+3N ��y�%�I�crqy���[gDc3L��o�<��뎽΃��ga����V��cu���9d���gB�<n���m�͛�hv����VV������ʾ�ç*p��V���:���������"��)����r�/w�wr���<)��� �
܁�yw	I���\���j���2=>�Z/�ew��St"�5�,[i�>���x��bU{�Õ�(��:�㦶��E>�#����4�ꋘX��p�^Uh�c��[3��_�{6	�C����;��(���Ǉ<���}b*B���p�yܚ�S%�g�;"u�0xO�l#4��ʜ-;�}^�'ѤЁXtIl0�!t]�mL�����h�{k��_��-���4P�P�j�=7�F\�>�v<{.�K�qe]M^� ����4����Nځ+���zm�9�4_����oz�:�R����7=Q��ÎcsWzۃf~�6b='D�u��P�o�ZŶ�^u�mga��B�Y0bc{�+Uk��n��U�7��XB ����C����+c���}��z���-']F�[��::��\ʭ���E�Ô��6�#8�8A� �@C��!���y�U�nn��(\lm̫���z�Z���I�_���(~���
rT�@�8t�?1<���ƆR�3�3�]]��� �{A�%���q0�7,޽����	v"�I�����c�/�b���� _��ԡ�WY��:�����bi��J�ͼU1�t��zB}���%�{�8����jN��9N�.�;(R��"�Hh����I��( @)D�� ��  ��D�R �P@���w��_�ٌ�z��:v�`fz��U�i�ޓ��p�P�Q������z2�f��м�}�頲��L�8�#�7hDmw���ҁ�w��|��7
,v	0�	�u1ǯת6r����:��D��@b9��iV#�sKi+�*@ݿ@rl%-�a8��4�bv���͏+������$���{�܄~w3rz���������u9�s�q{U����Qة�^ȫ�|�{���{Ǧ'X����C=Yʾ��t��X|a�����/h��NUؔ����`�ÿ��1I���z�w��˄7��pM��{�8�*̿u&G���k���}|+��O�q�]�Ll�{�z�R���[7�����1-�U��ڭ�at��0�F�P�Ia�y���?��\��7�ۊ�;��}iW���?m��G�zXd_)�l��5W)�q�3�>�����V����X���n��^��O�	�1�T�މj[s���[>
f�y���j�dMnE�{�S,�T���(�<�s�z�s���R�Dm��\!����$ 7��g�)�e9���tY���$�GB�yM�T���dn�̼�^����.�60e�h�'��N$�rI���ae�݂L�^�ˬڶ�5��(���h��g{��e����k4'�lN4UR�{�8�mv,�
78��J���6&���vr��N;�q�W'c�e>;3����%IHP@�� "IE 	@�htz��pf���j��'���-�-pPzA�\���nbG��mz-�f'�]��J�_f��'�]�t�6���-�3A(�|�`�ϟV@�^�{��>�碤��W�f�.NK���s���Q�j�Wј�F�c������q�ω��Sd����HU��p�8�����5��Z�-��2�Z=���aR�Fg���Q�Y����B�	��]�N�d!��ڞ���o֗��^备0�s�}&8�sw��[��Pv���W��>�7�a�~4$.d����������s8C�A	P����#{s����-��Xʫ�Ӊz�R��=5�ף���2��\i�SY���A�ɔ�>+��?�z����k�V�k�}p��/|���0��a�R��D�68�W�(���F��P�����~�k/���I��<#\�qG�/��v�%)h�7YE��b�F3|k��O�"m���֦])�&,�ǽ9^^�wV���w��Ϟ��/�[b,C��<�"�j��md;�zFAf��;/z}J�5A�]�	؞�M|n�/-)��0��z7s�(�nL6�ua?.ô�2'Vu��5��=�ڇ0ZȎ��͉:�s�+�t&k�2��X��]�/W��Ǜ��Ic�Y���xz��,;WB��fk��2�`}w/Y[�P].���FoU�ɼ\?�����N�S�8^��{���RAgc��w�0����=�R뽰�V��_t���)a�~�P�5zU>�����i��=ω=�ջ�7z?�g���R2��4ˍȹ"�Ŏ�l8���l���#L����s�8$�Z5B*rc�^Ǽ`�c��:7%Y����}��T?s)�e�<��[c��h����;v'0zUo�=��>��ڬc�v���� 瞓�?�q��[�pa��,��F��b�#�f`�G*c�{7��+�b��^�a"���XY*������%�'�BJ���Y�G��]G���w>�4igH����\�}޺l�)�h�!H�~��4���	b��[��̟K�U���氆/������_�ZŶ�]��|j/Sf�:P������TE��wJ+/z3�R_wv�#G�z9�*:��P��5�j�XŊ`R�1'J�������{}�g(��i����(?�Z��i�B��1����Tv�U�~T��; G��i�D�ىj�
�.n�{�!�C��/���`���`�D��A\�T��U�[F�m�8��GU��Կ
«��C��Pǹݡ,�Iʐ�7�R�}�ޥ���?_,��^�Q���Y4)ݝі�A�jלp�����*�l[=]ևI�%Φ��D�Xi#4j�w�`�/%<���U����'Gٺ���d�rDF<-t3�3^\ǳ� � D�@��$�  �  � ��   ��v�D�l��i������mɊ�����H�TX���Q28)Ap ���[3����Y���sZ��{*�F#�=����Ji��������)h��t���4L��VD{5�뺔F`&�~Kݽ���ɉ����G.�=���HH�BJ�����N�>R�&YV����g��i�",Y�}�;�z���9�x�ݖ����Xf�yA�iX�7{;����GMv�4-�9��>�7���S"��ޚ��5Q����¥��:� �{z�:k�s�C�&�o�w�5�=��`oV�M~�tS��`��dbr5���9ژ�'�ne�w�l�e�ʷ�/C�nt���Ƭ[8�X���o��1B�A�aNEE }qR�K����Q�]}�r��_m8�R�(2���@pZt�A��êu!:�@�_��d������˷��h�Ƌi��`��Ɂ��~�Ce�:nj��Vq�R�ɳp���W�V����F1�vf��V�
v�ɡޛe��R�n:nީ��^�G�B���DeBӆ0�n���l1��X��|��j�
�t[�vD���(��MH��t/l�������m̬��:K��ji�E��'K�$gu��nV�8:�R����Q`m��4�e�_[J�x�0���$��֨�I��ta�����uu=��H%A) "H$$I$
�����䧟ZAc|S��yA|�����`-��Y�[nH����#l�t�/���\ʽ|q���3{�Qo=�v[n���j�{Y"�%�r�V�ʌ�uugOVZ~����樾��Ue������@�D�ӌP]m�����|Y�kfu�u=��u����cշ�/�S��G(�J,?eDu��)"��g�'�����뼦���2�y�z�>**nLw��W*v�`�Y�	Wէ��F�ʈV�T�DՇ�U�I�x���dK�	�4%	�|�}�0�^����F�D�H�B���ZB�s��K3�Hު��y���;�&~�\	�A�8����KiP��o�
��)lq!�����e*�ّZX����\�X��&����%�E1�QWS���7��j�;�k1^�>��t=-��Y�����u��悫u��w��P�(S�3�ß�>��-/]��Ź�'7MH�:d��.f�s�c��u�o����
-5��mc>��/�Bɑ�FD�-n��.��긃��;���ET�:�;�;�+;��	��|k��zë���1�R��8��r�Xq�����7����)u�X{���:�R�u��G8ۨ6��muʓ
���`:�F(�|��0����ϯt��������l�[;7VϬ��RN��	A@$ �$�WD?��݃�O��X�c'�ͨ��3�r�n����g�[�Nx��(�x���p�ڋ��sll����H�%�M@�&Gp=���}>w�g��E�SP���\<���N���a��cy�Tpv3}Iu5��iA��q��NQ��������{��L�|�i���\1�]�
u�O�2��َ�ϰ�p~�Ԭ[�6٧-p6���#�����L�z���N�1�����U�ff�}��&�^�z�;��:-)�e�-~= �+Cr�1�d���j�~E�!&��������S󥗬J��j$$P|�����˨��� 9�(q=Q���}��Lж�oK��,e�\n�}�Z4�:Jg��g��r4LgN�������2ĝ�[K��됳�U(wb�j�T-
��3;���<�,5���
�=cg	�ӽ���_������^/yz\t@���hI�)��X�gٲ+���!�u��[��3�#^qyfl�������Wtt����[��]�1�`A�\B\(1��}�=�w�[M��t�VE�U�V'3;ʫN(ި�����_?^p1p�y2�[����[ӷ"o�@�9��G�N�ّ�
����`b9YM{6^��K��ѾF����AM��ĝ)N�w���HsB���Axg���.d�'F�¤1��
��5�٦ LB��� ��$������$ �{[)���7��b���7�l����G"x����9Q_MK�Y�@�-�ú�@��Ʃ:�4���vf�yqٝ��O�X�0�ÍjT�_-��M�^B����'�楲�ل�U�/-�:s�Y����`��Г��BF��<R�����o�a�n&�=�T���[��_����8���S�x;���u����+�x;f��-�/��b����������E�{��ͭE�=.I~!�=��S�r���o>��Ⱦ�a��R�/�L=�5{�;�z*���8.�]��(�1�\�a�H�&�q��#��p|_����Sl��?�[�l��ى�?Dw��D��&y	S�Q�9/N�"�ɠ6�ͮ��f�p�Q�;�㡉�}[��0�^@[}3��[}�q�z�3\^Ռx�df=�!<�����"���n����]�XΏ)�;��;��w��?�p�����6�+��	��̈́�XEM���3�zD���"U:���x�]n�{�r_�<�q��*���b��M��7�)x���u_'��߾(c�OG\�>��j��g'���wX�[&u;w���sA�@B���SrΗfY2|�N��y.���%us�g[�
^!�:3��m�J]���T�
�ǒ��M+J�U2j�[�{+�9��Y��chko����P�6Ĝ�303:�i/r���Üj��Uc��4�?t=Z^0�d���"P���w\dCǹ3gvJ�CJ�*�*-��՚,���%i���:�^c.d��!�+m͈6ﶛzhh�91eu�S�l�q6�̲�
;�k0����ёc'm6�8�o�jB��W�9���9���-�Qp�w81yf������@�I�~����de�qU�7n�;�k.��r]ݞΆdܶ��|����;m�q0������ǉ�q͘��X��n�U���â�ʋ�\9T������iES!�F2��Y5rSo�{՛� ȰIɣ��Yz{$f�'�J�A�×[�܆<U$冶�NŻ��a��G�J�l�Ā-�έ�U�ޣ'\�c3)��u�ыmK�1u�`��/S]��&�o.��W�������ծ�M^Lr��1ݒB"�qLT�	��Z[Y�����v�[,c�5�ۗ��خ���j��:��WE�������(^]aﻺm83\Η�0Q�0�N͋��3)��<~Z�٘#�y���:�J����|SolJ��9�Y�����L����'��Ë}̝t-�즦5u��0�-tmC��>u�m��������V��	5�dE�U���x��I����zc�mHr���Ax���ct>�@�.��ʞ���r ī\���1�m�x���΋�����\�Oh{e�`��q\�t|`�Y9&D=-�k�J��^�vY㼐�z����y�5��~OO0��I.U�_f�On��#�V����
�_#��-KU��Nx7�@뽙��;t��u�ydN�εyq���kKj��v�1(-z˕u���ܥ�{��a��W��!N�VN�au�;M�U�:�6�����α���F�|���2k�s�Iݾu�iԺx�h4��mf8i�o]I�F�����iú�S;�h]j�2㛚�ue�[�w��֝��7�+�oc�,_u����9���ʸ�	���h��{N�]�]6Vlk�m���i��&h�%L>Wm�ԧ1������#��5��h�g�F1>��Ƀ�����o5ބ�TD)��&\�t����w�O)>w�4��7$�=tp>�@����#\��Ȫ���y�#e�wxJ�1��̽ӹ=VUۑ����o�=AM��w�ġ���a������tӬ�9�+�f���ow��f]�	Qӳd���$7WcĻA6������Z��Zt���i�zF*y�qr��_�Lb���<ܗ��Ė���SV�r�o�4�K��kx��t+��s&1.��S�׺V�V�6���6l�RsJO%:)�=�D�rȱ��wc?o޻���nؼ�´�4n<�D��6���mJ�L8�ſ�x�
���~??�=^֞�0:�����E=�~�؆�ۤuג@�T��<�,Ҽ=�}�[턘}*������R~?�ݝG��z�G�m��e����|��b����O����]�O������(�(�ՕE���ߨ~���gr_[$�����U�?cv����|��v��MB_���'�	��h�bL?�`���?*xעy�����~ף�~��3��$��j=7ɑ�G�*5*�c��U5<��N��oj���{�N�(��c����?c��n~��j�ޏ|x���_8+ژ��K;NF!b�TYr����{��B��aK��̱u�)�k�W^��'�O�y��ٹO���������_�`�{}����"�Ǭ�~�W{B;Q��f$W���%�g�{�{V�y�V��+��O�}y��m�|}H�y3�Dt>�cơ����UՇ���ϾLc���{�{�{�xI�{y1.�9P�������P�ɶ��r������I>l�����(4P �~k��^�^��/nN�m�>�%f��	�-�z+�7���x|���E���4�օ��B�7Mָ�`;���L�{�o����� � � ���޴ü���cP��6:��J��-m�����^,��`N�+kn`���9��F���=�z�)���]%�����;&C��$u��y�XČ�zN�WC��;�����<{�%\�`�Xg24�@V"v:���C.��tok�o���:�xRf�������/�1r�}S��c�R9)�DX}��X%x"�?D6z(H>g�b��=ZB?F��be�{x_��W#a��vz�K�tb��N�[����*��D� ��.���œ�&���
��G���\r�1��M��v�:��>���Km����P6�����nJ躐��݂J{�ζD���_�M#����k��a���	�C]3�9ӵW�U&�7��7Y����.x�zȈ���	�EϽM��]�p��z�^�ݖ����K�O(1���T2��ѡ7w����.]�E��rO_M���*���E���ws�i}�u��>+"o��8�_EѪ��z�*ވ���Ra+ZA���
�*nJ���!�q�
���ZE������1�y�;M
s������_'/�&�+�o��vWPMY�X#�0sc
]��y�F�x��ӹ��V��
ƙ�ep0uE��)\�;��/eIۇ�)������j]c��w�n�f�>�v�uYW��a����]#Oj�4ǽ��&�>B�ʺ��$�>I �$�GM�;gM��K?j�����C��O���׬f��7�xf(�>���{�E0|eE��v|{�F�%�X��c:���z4��g��2�:P�99�tx|M�}�w<�Y17�:������!�b�$�w ��+����/��Ce�:n�����!�^�����a��=�{��Q|D�ALG�L����B���/p�F��f���/�:n63М`�X��ƶ�w}�cf\�P�O���$�a�G���%G_]
�}b��rE,u�v�H��k�ǧ4��j��n��>�P�>�'��l!�8�p�9�(7+P_�ɹ���ُ@Q*aDf���k���o�{�k��To�s�]`�c����h�@�D�'�*��������:y+�?U��{���T�=_��ds�^��u>8�����ۥz�,�zX숀�a�6�[/s�rs�f�����U�X�TP�&;�}�p�N�,�Y�J��<�z4.ʈV�Z���������+U���N�k�A��/�m6j혏�	�xg��7�B���L:��h-��OgUQ���OuI_�d:I�oo��������x�M)�8�CO</n�w����7.ʹ���3++��ٯx�^,zr'���[i��l<��wM,�|n�mc�n|��N���u��%�ع//�\��a�2439�v��m�O�����'�D B�@ 5�>���oqr����&:��&~�\	�A�ӬG�W���j�
�ݿ@rm)l�@PZ�eh͍�O�Q��(1��aƋ?f�ܞ�8����=**�r8:�4���n:.��=_d)�/D�b!��ܯ�rOՑht��jT�o&��5�b�����L[\P^�a]�1�+q������vmU)9�ҕ�����5Y�ې޷�k>i�/�Q>.��O����U�k#����۪8�&:أ6�u��3�r�T�8���[.������G&�q��TN����k��'�H�h����T9���p�;迏K�Jj8����Sv�+�f~��Tj��-J=�9MY�hq��e�ةp���z�.z��ϔ�2�g{F�{<���\2�|wD�=���d`���}9%q�1��Du��\!�[F��NH����\]��rj�kzz���|X��߄uW��U���^b����8pr�7+�.cȪ�ёe�-5q�1����j����L?E�	׬���H��hu���4��d�(l9�Q=u���f]SW�HB��k.�]���x���,x��w�I����s�M�^J�f�i-9;*3C�r���ϳO���U�&Ǣ,Y85@�Ds��R,cEK�{�;�DZ�[�n��5:�q�U��ʷ�;.�qr��+�7����w�����x�+��@@ {٬�r��*;�|7SP����W���3�hՌu1���N{��ω��
l�������J���y-$-� F��Һ��_��\+Q��U�ͪ���(�s���3��ߔ圢s��~���q��NY��@B9�Z6\��*�9��#;N}ېr���m�e�X�}l���;Cu-����4t�xh\V@�x�оPb�F�����½R��X�=&V�!����j������9��.,#��#����bG��5/�`ۡ��כ��'��7���!]�]�Ssl��ÊJ�(-��k��L���=y�Z��;���ם����T�u���=	\�F�)�\�݇���\�F4a�ch_	�}���;�}B2�����G�L�|A�=E,�b��zN��)o�I��LC�O��X֫`߶�,�"J5^+�OWf�	]�o�U1�x���:4�xg���.��s��=�,3��yK�0���VH��l{�{׸�rZ���x}5�>�	C���,9����iב��4����6zX���i��F}ح����Y�U�����8p��-Z�$s�S�K;�u�v��A�9ӏ���6�c��Ԋ
���.6ӷ=:,;=Wf��l�fWMU��s��\�ĺ��A�NJ�n�ʾ;��^�']*�<xX��\�B�rb�%�&�x�Q���Œ�c��)&+����$�� k�c���wZ�vSz���K|=3�J��Q�$d�;t�&s�}!ʨ���l���}=���5�,�����zD���zz7�&Y|���>wk�U����~�2<��C�2�.v��k}����>}׏Dk�c�P~U1]����FC����ͧ��*m���F1B��:���~y�v����c�i���ۺ��*�;����f�d4_�H觼hm��|k:̬�Jޘ��޿���dD�#�Ԟ�o�m�(Rն�]��|j,b�l�Y�t�TQ�}8ջ���k��~����d~�D�=���>����鐣��5ƃՕc2�E�N���h�_���ׯ�s��<����@���di �v:���B.�]��T-ƞ͟�'9{�>��g_�_"�x�w�F�Y\C}��X%yH�xO�1��R�W>�z�r�y�U��c�՗l�k�;��|�a8��:1}a;�P��g~GAP�dpR�x��׵���'�w��umX~��ϑ��!"��#�-��	F7�!i�ʪb���V:E���#�0?��$.Oߪ��eɸ��.����?:��E��!�x/pT 3�a�+_�Ѿ��ʩlc=rRDa�ե�Υ�-9����n��WI�Evjvͩ��Ic&h���Rﾋ_'y�Y�a�W�u���B�N�0ff }L���^�.�<�}y��U��RW� ��Jz�75{c��{Y���bA���)?,"�˘{uc���$7!��ҩ���|v�r��>��;o{���y5�c�Ȉ#�H��	�E�z�>��ӑ����۲�3�������K�=�F�C���O��X�a|]��}te߅,Y�x~�\��b�d{�E�!�Db{�7�]Wµ��yOw�,[��i��zeM�W�pX_�#�ƃ�}�y~����v[6�g���)LvO�aC!N=�Pp��l�c�.��4J�i�b�����_��[��5������}L^N*B�a���;ʺ,��`Fi����ӱ�����zw�Y��;X�֮ċ>��;�	zK��BOp>G{ �8w��]�M����6_�t�|�&��O��K��SexO��/�DQj��<l0v(q��L��QB��B���Ή���\�h������B�;�#u�/�_��w0��*ʋ��d�p�1��㯮��k}c�#���z���^���b�_Qc}9��'*�Rz	 ��Aځ?t���	�;�4�N�:��Ӕ����.�WI}�7n��n8Ϙ�t���Y2���^U�����v�/O�z5��'�.ڞ�ِ��1?1儆�]�P��j������f�ke�&]�t�;�msO�Pa�Ⱥ[tg%��Z(��]1�_q9��Y F�z�<=����]@}��@� 6�ּ���r*{P�Yޡz�u�c������ґ���Hbz���"�};[$����Y�W�����:���n|��d��۽�����NR9G��(��������vSX�#�F�O�C��Y��pK?b�m�YK�	3=gp����g�@]����^U��x䪵��B��1n�D;�JF��\|�m�3�>ݡ�;ԑ��@���_(#G?D�"�&w���/�.��`<aP�P��"*i�#�n}���BCv�ɼ��}��<8O��Z[�	���D�9*�Q�g�3ds�
�Q��_~�>�ї����<�;���!{� ��r��;����w��x��W�ya��) ����lq�3��#�T0˄I̺_����u��­]�զߪ�57Q�*b���-5��5O��p��T��(��B����Ϯ4HBa�;��u���K����ҁ�S�`J������j���s����sېj1�u�������d �{��Wh�����jXd$f=�j�]4A6��n@�zv��(͌�`��:HX�b���5�����GRi��g#�\N=��Ҋ��������A&lw[���7�6�f��DK]S��5kj�����-�Q^��K87R�pԠ��ܺv�V�Ejm!{wad�P�����%���)`DSB"�0�_�	� �DA>��Z�u�̨TS��V������g	�AK�&Q�ދ��lPB�Ը�e�:�4��H{nR���'��NO݂M4���^���=[��n�4\k�J��"�0.���2��f�3f��]鉻x�VE=�ݗ��|Ͳ����j���	G@>���r��}@�.2�*=�T�{��V��˺��y��8���
�����H�ϑ�b��+���K�ʶ�����ژ��;��E<���u5�VMGoݮ�3>[M�t6�N{���r;�M�۟ejX&*�Ey{^��0(i��LG~����xиV�_�0wSeG��f���}x���z��uȹ�����+st&�b�����zfK �`lAƆ�hI�-�w{U�lˁ܌�=0k�C�\(�����:��g��N�7�#�Ө4zd�qO���:s��?��������(R��d�u9�EN�M@L7_�ͨ�xaqh�$O�f��%��_��~ß�����G.y%�����c!y�u��_y�[����N�8��I�^eD��3�(��z����!�~�/�O�;�W�+{�,�̆�D�؛��k
�8�&�'��7�[��^i����5v@�ms��r	i�\�Qk��S�)�Z:Ӱ�t%C�|��P�Yˎ*ׯ�mF8..|�P,AH��"���,p�*�:w{��̕L���s����'�@�PD�I��q�������Ë���*�I�D��w�]ԑ��Cm*���[>k�f=ۛT��u��}��&ő,^����z7����ٿG�lإ��� ��XMV��<n"`���j�}d�����Ƒ�gH��L�mN���{a��y;��v<���Z��9� �S^��O1z)��{�ǮrK��"FP�4���6�w�c�>��ӂ�j�y-��z���I��=���t���;����z,��.���jĨ��1�*u�W��-\��G�f�����f8;��q�Ce,�MXǎ�23>��Gb��`�����k|�1�2��/���w�C��#m��p��*���v��ϣ�[6�+%V#`�a��6���Z�u6w��׺�cpdVԎ_۲*�;����f�M�E�Z(t[�hwg{.�K�
=W��ns�^ѧ3�Y�A�Jw�IB;��Ͳ�e
[��p.פS�qJ�Dk1����u����qlg��
fI���� �7�Q���qȾe��>��Sҫ�{EJ^��ؒ��,�Z��V뻕��)�˲����Gp�$�ޚ��Oq��ML�W�����g�]���^'����ջ��-��)[�o&���u%.y�7������C[��j��v���1_k2�oE�	��'��,D�4�b�Z�s+�}�2���� �� 5���g��ޙ{�C�ut:�[Q�b��~� A@����!�t:5��u��f�[�{77��7�(f�Mn��t�<��r0S����`���%PR �~�cOFb":v{s87[��?X8��c��ځ�akvz�K�tb�Ӻ���w�pAT�Q6��J�^��5�/�^/cU�K��>� ���]Dr+�b;���	M#����*����,��<!������}UV�o�c���4L�r*��jM3����k���=3���	m�b!�=���On��T���z���{" �9LN".}�l����.���`�:����a*3�~�z����Ł˂Ϣ�;�rw�7G������{�]��r�7��To��3��x�KQ��z�q�,C�t)6�i��zeM�W����՟��eQ�]����)q��Y8���~�u8啷Q�ĸ�����|\��Z�f�
�L�VQ���g��k��W��w�bD���:
F����]��,l����f���:P\��fO��, G{��c�V,x����R<���C�]4K�<|悧TAG����ŦV(�-;��Y�2Ҏ4���jN�
�B�=�?�t+��tL����P�Cq��f��u���[�>D�V�vP����f��p�Z�Eb�(�vݿ��έ�Ȍ���:�w|���[�f�D+$�wp��3y5�\뭝Ou�c���;�$*�V�����G`ĝ��s�*X�|�X������{w:L�3�/M�������l¢�xr�7�����x]�jZ�(�=*;y}}ƹ�Y�B����Y7aQ7��\`N����{��vYVA�%=	�4�%�+�#���H������r�u>�{��P\�y��ڙS��"���jn�q��L�Ь���tsL��v8��`�,T��3�ʼNcm�f��u��O7��XX.���P�"�X��5�m�G@ɗ$7*�X��.�V�4�ۤ��x%Wo7ͬZ�É��$óD�3�]1�#5����v�6�fI\�2	@Wo=9���1�,�^�L@q坥so9n[��I��cY��]s�6��Ɯ(�He�Vz�n!�Q���U����:Ɲ⥅&�C��lm�Bs���뤴9��d�:k��Y�}�B�e����Ck�����o`��6�`
�
w�(M\��ǲ�R�N
��a�/rf
ӑ�B��i�ٵ������{�u
��������6>Ƌ��Ԩ�5�ּ�u"�J�H*l��)ʷ0�m��z�+v� ��[*�%Y�7���^�K��.��&����Kt��ckwv�Zo�V��dVͰ;r��Cc�O*u�+�fC��gE�������dkKM�[Mlm�{>�d=�Ja��=7(+��+�3���X;�Z��ՖD��4�#�U�����-5|j��X����M�8�}V��r�����S%�	�<�r�Ůk�'��3�פ�N�|��ڲCk�m�m:��\����+(���_\ev�����*d�=�T�XLB�{�.�bZݞ����;�t�D{Ww{$.�Uz��}�{*,�v����[�1��O&J�Y��X��vFKp�&s�B�:��.�)pZ�r*JJ��Q�nT��DzѵSzw�x��	땛[]xT�M]��kd����Tܧ;�&�T4�Y�ը�f��������3��=[ۏ�1ln�&��9*k��x�P�B���{`K�׷�(�6y�@���6��i�6��m!i�],�����8��w[E��͢J]�aj.�]̓;g-a;�z�!����֫�:xk�q=��"*�����/�U�3�t;�y|���#eD֌{zZR��]�݃w\��Ɩ�v_g.&�.mkfKű����9�cS���V�ɖ(�*�S��Q%�8��t���K
[Rm��7����C���VS;��i�EGl�]��@=<{���{x�f�J���j��0a/����Qu�6bp��oj��3�Z��0�#��3N��&DL�Yb8�8�dD��%�	Hg��uQ��VE��y�n�=>q��Wo�xO^��й���r�! �S�����AC�_��d�}�=��I=�i�9-A��|�o<�u��ش{ǷK��)�*[c=�m�#�ZӾ1��x��g�\�����uyf��~�
��%ڣR�q��h)�a�(G��=�S)��Lތy�h��i�6Ӣ���m��ԎF�}�|缇��eQa�v����Y;Y&Z^��/��"B�R����:�<��%]�m��WU�61u��*K�����dW=m<�\�O{��󙚡g��װH�&ѐ�o^0���bԭ�.�������d7�{�O9�F��c>���"�3mneC��ְ�6�^�$�[�u�n���x���h��l��#עϕ�J��҆�me<�W�;Ifu+�h�C�x���ӷ��9�'���}FͩA���{�\��2)����{�g��-n�{�'}��>���yZ=o>5���)�|m����+��S�rkn��z���p��n���,�Sl�U<����c���׳B��D����EwQ�[ݣ֨2��.��L˝�t}��-��d��0�r׎����+@$�x"@ $�x%ԟSH�>�&D����>��� ��+��;U��2�j�E8�s7ށ뛓%����L�P����̩�`h;(t�z�ʀ��Z��hS��r{ƙp��Q>�t�S���U����v�8�v��c�TToĈ� �p�1�O	q��A°��-x�4�[��*����w���}$y���7�q��NT+��q��D�����:i�zy��`˦7��Z�_�����ѿ�ˮ��V��	;To�X-��6�g� ��A���K6&;�:�f;9I�w�E��G���9g�v�!�u��S�H�jz��*#�N@)f��8�N�i�LhUԳ;�x5���F�/��g�oj���ҷ>fz��J��<�z=�#Ѩ{z,P/�Լ�]�R��zZBe�<�&8:��hԚ��9�0�^����4{3� J����X����upޏ^�5(�����C�|;�\d����N��EM:�pmϴ����J<�{��Ƿy
f�|�W�}�_�Ӭ��44�aF�cV�.�'�IM(�Jp��a�w3��zO��ͯM���l�Լ�G7I�ϕ�g�n���U��\橘�[U�l���@�~��}�^�\�o��L��mw!�:NR=�v��t��E�q+��`p������"���ܛ��j�aƘu�f͸Vq�ѻ�J�q�d��UScs�,z�Fe��f������� ����6FNf�7���cn|���k����S����>j��k��c68�&f�S{M�3�x��Œ���su���v��}L��n<��#s�*b��[`߶���2��R5r}��띔$�<q>�׫� E���`7�E��9�#��n��Gy��ӱ�'F������D�޸�e�7fp���΅#�������E�l�u.|���a�a)�l����j"��ʀ�'���p4���V(�>��Z9��&C.=�L�112�?w���w�q�1���pYg�S����\w��������Q�Cy�ۤr�Y*R_���������=�}��S��1R�c:�H�V���m��BՇ��:8��}?��1?c�����L�FU����������=u<#X{^�G Z�b�^�F�N3��C�a#�o:
�n������<}챳G�Ю|}�iy-$?@��#iE�A�]SP��:�W��b�m4j�:M�=���9�%��i���h����S�Y|���?�WcS���ȁ�gf��U�����*3�5Ks�uu{U��Ӟ�YS��$ϗ���Vum�m�]S�����_�y��C��z+D
׫p>�����^������f��]Z;J��eY�\�*!������W(��U�f��sA��*�ʭop�jË*GӐ0ʵ�;0��G��i��y�M�u�D�"@"IׯYl_g���~�:��1��!���G��ѱ�1�o�Xǎi������fB�5;
{��}�������Z�9��������2
B����kNyW�L�Z߳u��efn��V���q^�\�4���(�xaqh�$O�:'�ď*2��r����oB�igo�s�����Q�;�G�����b�N�8��I{C�..��}�D�͝��:��cۭ�X9c7�ڭ����'�\�NG�������b��77C*���F2{Tn��U{*�ɥx�U[幼)��(Y:4��}§+!�뼯���ٿE��`��,F�pPO��yRU{ͬ�9�L����E��mMƿ�# �8�20)����kjwN@u[A��ȱ�,3�D����ݭ��kb��<X�H�|���(휎��IXDF|Ñ��i(�1��l8I��nT�s.�����F̾�ϧ�o�#L���ݸ�+�u�Iv2}@�*>�*�2������Q	̡�n��c�1{&4,�����p��3L�	��W�!\�dA�����CN��\6T���}{�䚪�WD%�WE�Üy�A���fs����y����	mp�F���D�����-��*������|�7˷�~e]E����,�6�a���Wc4qś��&.�SZ�)Y�����e��!�C�m��̻������$ � �G��d>^�Y��haS����]�ȅ�/�ۇ�<��l�|�,�X�:Ʉ��v�t/D��ʈ���m#00x��诤��X렂6�EC��s޺l�r����)�v�o{�c/g�u���<6���έ�����z,0C�RP���i���`Zς�p.�^�ƣʈ�3y�vo�NNջވb��}���vܺ���8�;y�^WE�]�.F����_�b�#=����9ٝ�k�+�o�ǟZ�c��u����H僱�h+�>O|t��ǟ��Io��Q��=�㕾��{T�z6Fr��̿��=O�|��r3�NZ"�`��G)��"E�}Y�ٚ&%��u�wzh[�bA�=S�o����kv3�z_��֝�(��F2���SauT�L�B��ۋw8��.��,������/uDu-���SH������ULt��C
��Y1S�{�!��2FA�_3D�"A��O��O�w��Hc1߂t;�H*�t�k��0$P$.����<bP�v:���9�l�/�����'�"�׽m���9;e��ʾ�6e��蘘~�r
��-[�4��)w����~��z���(i��׏K��a�$�/��J���[��uL�W*�����7��wr5����a���0����צ��=Μ �zb�����;�J��*;�� ��==:�.����J�5q7ܯ�(��g_<��6�Pb�i_�C'�\_�S�]��pd}�*�-�_z���]q$ߙJ�f�׹��	�ǷuT�X�x��ۏ�����&�f�A�ĸ؜
�JÜ'��/���V�}]H��ձ�m�tX<�8� ��L���u{M����+��O��L���Q尡�å,A�7�T8�s�t(9�R8G-������@q`KN�0{먡z.���8b��7�a8L��3'�9b*Gla's���I�f�B�[>���T�_��/я|���zo����|4��x���(Gw�D��Rj��k�{P����V��}�]>���k�sԫ*"i�A�a��FO	q�R!{�m��]�{�q�oE}U�%�]$R�[E�g�j�=��A�Q�X3�8l,nHA�\Xؘ����4b�g���X˫�*C���Z��$�Q�wJ�n�q~"��ߑ����s9���>>���J��e�t'���k�s�2#�����|�SӀs��Qϭ�Qo�Q�7J�?~��nS�5��PF���=��[��u��#��:'a:OmT��'�׀�r��eY:9PE�E]���)���ru�$֐9�	�˜�޹B�%j���u�Ah��܏j7��Wxݑh�2��ND'X�r�d�۩����k�� p@��$�}q��:�{<�փO�0 C��H�Liq_O�������X���J~��cʐ�^%'t�U�n�Ed?��Dk6 ��R"�� h𦍌�����]����v�~�=��n�MMu�h����C��ÕgָMǣ����F��E	�X�}�>��W)��t�ջ�i����ɰ����ҹ��~���=c�PX*&/�ǥD�7��������Տ#���s�q{������D��NN�0���AY��lq�34��!���p�fe���^Z�>(�StC���E)7�ҕ׶8C��YŦ����fҸ�	����[z���>u@�g���}�8*:m�"�o��b�{�!�8��x��V��k�Л��z�7-@c��3����>w�G�����$��q�Øg���xT�^�>�~]��R�(�3���++�(<����'(���W�+ӹ2R�}�/���\w��S4�Q�+�{g�*|��-�n�4C�t�79��=�ʡ�|bn7�f����4��y����K2��"F�#�Rw��"��xϯ}zB�����>�CLT��:�eq��y�b=N[=zj��*�b�fk�%�N��j�iͻJ��|f1w&l=ei*�w��Λ�m�7�ɐt��$���.��O �Sum�|?�@ �A"���F��fUu�d2�}v���πS6�~�:������	O�����r؏k���a��wd	��*2�ֈ��E��]L/G~�8�0�$W�·_�U���<��J���1�����u�ph�����=�.�1�p��}�v��Ųѥ��Óa9�'fٚ����z�Ole�op�RJ�y6LO�\8t��w����WB�Z�~�ϻ���P�yΜ��C���R�x.�\���g�mHNW�����Y��<!HS�F4�o�cN��V1�zx�h��7wocW�W@���n��~��Jo��=���$z�`�4.)���(���4��b�<;U����{w�m�c9�$u�獐�`��qA�M��xaqh�$H�0�l>&Q
�ʠ����Ҹ���WM������ʜ_���ÍJ�+�qk��b�l�	��m{Y�RX�Dġ����/�r6���_H��\D�u$b۬�"�U0��	���tTƛ���ژXX�Xg�вdx)_!>�G'!���+����_���X�dy�4���;�5����}k�������#\�z�V[�M�tc&V���^J`��U]ȝ��v+;�cj�)M9b��ժ��7&E6�H��Qru$�[s�d=՘�}��.�:&�K�v�6��}CLh��=8�}&666e����A H�Ű�z�Κ�B�=�[Ƕ�:�# �C�6L�
G��[7����7:j��z&%�:Ɯy��]����;j��􊆚�AЧ���z^���%G�8�����y�^��vpA�C��?51��:��X*P��M�ު��
�{���9%�O���%I���`r�^�mn[��UZ��"�i���p��z�tY�p�D�->�i������+���Kq�v��F�����{>�c��S����]�S�n�?#!�c�S:|�*�exF�¢F��Om�DQj��3�b6������}tF�Ȩv��P�]6o>�YWH��VVvԟc�3�W�/ځ,\1~f�����X��<h}�>4�#��\�)VP��m���+�^:�ތʱ��R����r��C�}���r� ����̓=�>4>��q!�#���-�zm�Lũ.���r��=��Mv�������(O@�BN��5����hkXmܸ����c�{O��K_���KwR:<޻��x8#�#�����G#9h��WE���_)=qވ��U�v^]iۍf�&��M��ٹN�����d�7^Q��79%0]��bfԒ�3����U�(��x���:�OM�1�
AC5p	湷.�v��V���DP��S�l/��l"P�ks��
��JC��d��l�>K/��c��Uu���� ��2��a�*ؾ8l�ً����nB��$�U�~:1}i�B�}#�O�_g �|�b�j����uȃl]`����p!*�W�b/��徵#(�S�:k�8x�(��ٵ�\��\�؜�XFAGbI���Z�1,�!���o�\@��N0g#��ތP�F��Jw��e��X�ErU1K�r�0��"<A��Eu�[g�s�r6��Í��8:���]R����0��,#i�-�Feˉ꜒���p(xdW���vw��fnpuV�z���Xu�S�Y�u�C���X���S�ݭ ��zeM�ZjY��F-ūחܲwh��Pu"�ōU��
ۨ�b\f��8x�
e�e��ވ��XJ0z�<�uֻF����bPS�A�L\T��z�B4w�t!������-9�
,����ˉʮr�̿f�1s2�1.��ld����B�%�|$����W�wU6^{�ǋ��V�Ύ���kfr�G�dc�:n�ո@OT�s*Y���Q`L���\�	lH�q~��z(i������T��~\�^۶j�j��دR�IYw���sH�Vo2���'<�F2�^��Y�V�w�86�Z���˖�Qa�e��0[Uu�i����z�l�E�>�]�q�[�ۀkyzK������;�#Ӎ=kn5|u�2��Q��{/s��D  �vp�y�]�?I�joN�J�����p�=��R�����H7�b=<$�zF��Z����н�]�llm�P�^��)�;�2,b�v��'*�Ԥ�XdQB�j��M9"��K}�vB��s�T'SH�S�%�lf$�Q���quN�qgA�Z2W4.�����UG{��q����?X ��cn�5�v�!�{.�����Q��E�g�ꓧr^r�yDk9 �/�H2��&#K��I���t�5.�sfz��z\[��g��w�8���,/Ut>��z�U�G ��-���g^��Ю}OP�>w��\�g��Gj_Y�<g�&Cq!m����7
/�xTµ4L��#��"��b)UNiU��F����4�����V��U�U�~��T�[��q���u��1�n����x>�\���V<'{�՞�}ق�ú���s�q.��]�M��O,1mR�C�oྀ��Y��.��y���~?;?��Ҍ�n����kV��m|�݋�⣛�)]���(r���!��6�y�L�����l�n)�tI�б���,���k^�κ!�)j��F�ݤJ2�	�����Q���
�Wp��`6����J���p���G�z �T��d�ZaoF�h�y7f�c�l�2�X��L�܂�
�In���X���E�tn�M#��˦1w7:�-�K��h����-�Nl{�{}5��:������F}ifٲtF��Mٜ�u/U��j�ҍL����Ҳƞ�kI;�,X��-n۹��{�l��.����*�$�J�i�6ܖ�.tn0z��	1��n�������[����n�q7cn[ �����|Ga��r��K�w�j(NV�����<�Z��(R��K�i���VC�ozn�Z�|�2C�x���]d�)w0��ف��yP`�\�!1�X�4P/�|��7����1F��t�@h�;W�mZ=/LF��.�QY��oۇ�3S	�����;�dԛ�P4;��� �֌ˎ���f� �ojV]t��֤ջ��!�\C�.�]��\�Jm��:g<��P�Z�	5׵�YQ�I�m(:]
�y�p�[���e�!�5�v�'p'���jz��0Hv�:��U���˵�CH��j�Mu���;R����������ޢN�U��Kŧ�V��"|[�l�nҳh.g�|�w'����U�>Ӻ1+�V�L��0���Jc)�J��B�9rCݛ�l�L�/""#�.ܸN�o,v��z����֙�w��<��W@*�
BN���'B�ON[�b=�+Dݬ�<�/�߽cպo}%�He���e,��:����ƕ����eq5{1��1�a�=������%˚MT����ڂ�Tw��<¸�@�c�f��7�Ums�,����ӎ��Ru1e��N�>WKN�̱G�!��|F�`ur%$����f����3�.�l���Q��q�,�u��>a��ȨZ/��qP:�U��.�\�	�W�c�N�Z�;��=���'��@ᔞ1E>����޴�U�O��3qP���!(3:Ύ?���u����i�}w��n�����Z�\;'H��Q9�iۙtV�n��	�Ġŵ��X���H�:e芣���SQ�����yتk|�3[�:�ՀS�\c�9n�m���|uNh�iL��kr���m�۾�t���0�R���F�h�Rݨ�%�!d�J���*�W�"�c�u�Q|�:6�Lν:��1�x�e��a��C��N�]�J�r銝2�_@Ft�o��������܆��*ֹ'T�ԝ!�kM4�:���B2��6�ʵۏ.����f6�b��6�-9�B������.�R}�R@�qP��	�N�r�����Nb5�p�[�����T�n�U �S8���*X�Nt�/�=�u^��[7Iv2��ׄu#'9�A�fq�漎T��L�r���>u�<���T\\(!���R@�F;;��1&H'7�d��2��㸏UG��nӴLPa���ñ�ׇ\_K���1�KQ�.�5NrnE]J�(�j=!方���~?�����{��&u����e>}��F���zRDT��G�{
Z�wd�dQx�Ҟ�2��s�Jϫ�������&�h�c5�j*0�D��¦L��]�ޙ��m�,fr�P�j�ONV-X�y2!gR��}������|<���lj.�*����FE%&�e��o�&dU<�y�@�I�Z�w�Dg�sa�J�Gv�(�	�"��EDB���ȉQ�%D�5���7j��m����oe��篶�-�3����9+&jS��:(Ra'3�E;�?D"���ē�=����m�����)���k�uom�F�h�I�1���F����rY�G(&�nE�
�6�F��{9�rd&��uĨ=��#ˢ��l���hE�f�]�ə�=��I2I3P�#k�{��x�D�F.�eBC=W5�G��ns�%I�r������Gr���?YNU�τ#;m�"�L�������X�"枢�w-�>w�J���<�5v��	���Q���P��Y|/г�I[�3rK �����Z�0^��ܛL��2c���;;�lK�x�IN������['H�m�q��C�	���oOr����Xo�¡dρ��hz�__�{��_w1.3�P�Ȥ�d��x �&��Fo��/�[�}9�xo�c��Ñ�P�*�`���{�DM!�[��^{m��|<F��\s8<�\9n�_}3�>��q�,՜&h)q�&i�\T�F��}�)=�_d����h�cC��f�[(�e?�P�vV�#'�]������^7r�E,�T+��O��vk�#^]!�L�z��Czݶ|�m��#�Z���@�J��:j~;EnӁ<��F���^z׸��xO��P��B:�k�l��S5��8�?t�8�C����[��<4��LQ{X��_��m!����a��v5�D���ӊ�n�5c�t6�j���ǩP���ǐ�we���r:Û&'�`��:B� ��":��.~
�\+
��2��C����ٝ�c�^˗�To�z�;u������6p����B�J��&4�z�q٫6��67�y�Z����-��������3���龞uƇ�X_t	�̃��P�TC�u+��c���"w=�Cg��atMvrqۻ����gk��2��.���7:�v�`k\�oO��D������}���c�z��^=���h�
T4c�2���J���]��)�(�"��i�i�-�Vq��Ω/f8ɗ�
u-o֮��#��"-Ḷ�yy��Ga��1�l=VySd$ʫ����P]a9��.,#��?q�>��ʭz1���%^��?O���������q�/+qx�f,'FPjT�Ah�G�8_�.'չ��y﵋s�|��N��p����� �vװwO�̿Q.�u$b۬�#g�b�Kݻ��lO�ލ��rT�\f����={B��dM�'�$T�d4}��W��lߣ̶cG�W`:}���k�!�y�����Mq�W�\�l�Y���h9�8M�G��[46�t�뽰�ݵ��P�U�zƏd�g�zh�?C�6xxt��,2��a5{�S�}>�w�W���#(`�Eƅ��CKd�1��UM痗V=�gS�z/���6zX�ど�[�B�ݸܘk��_�[w���"���ՙ�;K��KyC�2���Z �r�%��wL��&�c�v��N�@:�`�w5�>Q�W-�j%1���E'�BJ`�R�;�0�P�*���v���d8Lt�gל�o&j�=��̭oÿ�_�%���(!>���=u�AdT5�Sz�kak���w�QBfG����;h�fs��h	f�szL�sDʧRј�9���f�+i�{Sr��w�k@�1O��%^Qͬ
�V���ϙ�#n9�/l�HOf�Ρ'�AFU�skasm�Y��j�On��z��#2�l�fc�ӂ�pH Gl�W���6�2����2=�.��D�>D�|jJ�luͲ�+��I�2VEK.�g/�}��m�?�V�YM�Qލ[ vܺy��'�;y�^WE�6?�}�]]����I��TGớo��i����3p9��bN�����[��<���C��	cP ����z��+��u���\��p����[�
6���<:��;�|p')���E��]�SAsݶ��Lx_�n�ݖ�	��CҢ����m[�JG-n��z�K�tb�Ӻ������nf�aʴ��Yaaa�\�&�9F�p$���=u�}�ܷ֠$e�<�-��n���FT�v�2\E"�^����NC�.
>�i�d0��hy���[.a���AuL��牏Ui���7���Wxy�5��F�݇Q�K�c�3��p�qx=k7^��P���K9Z|�2�^{��)-*;ǼXݔ���R�6�Xi_ч�\{��.�M���%@���F�7w��C�5]�����t��Oḫ�y�us��由�ǖ-���kH7�^�YSrWP�0~@��#�������;X�U��2�z������v&�;x#��`Ԩs)������v�_\v���`�S36�d�c��\�+�\�.so�ќ�)�K���xα�Z%��VZÝ�����Z�������-��L�J킋|p�e��PD������~�����!�G��s)��]�b�)l��IPp��l��͍��K���Uw�^������r�j�3>��`����^�!�}����u�g��	A�_����֭
���7�P.���O��64��>&G�~&�HA��!;���t�ʘV~K�I۪��흜��|��G2��t�;5n�zo���R��Ǩ)��L����(B��֥�N�lFI����=�b��<���h/M��`�t�~���oz�:�R�����b=i�z�ȟ%��GT�s�nV��2�(�{���䋿����8�F'*�Ԥ�["�2�A�y�͸q�o�����ZH[���:%F��_�+�~����3�j���������\�)��\5qY"��jޘ����D�.���/O^�\k�ֆDd<���.��>NR9F�{"w���1Ui��(��x�9��_��p���}�����;��:Y����/@��O���&��Yz��2��c�_V�N���쨅jpA�AH���5�Z5$��9�_������E/�~��<_����9�7�d���ʙԮ�
d�d�{oLɷ%wfGG!��Ls�5y���Sm,����z!�b� ���LJ2�ݗ�����^.���@Э[�+�{� ��TAo��LJ7�f��~IdK_���F��Ȭ�> �릷�����3�	{�O��7���cCf���y;a�j�Xh�s�?�/ƅ�AmM��Y*�Kdu��y�=�Ƽ_�|�?�B���&Җ�NcZW1_#�ճ7'��P}����=t���_�5�߯�Ҧ;:s��ι�8�X����3�@V�Xb�T��C=X�,'ve����+ٯsP�<��J��������������C�K65�q�ʘ�oՐW�pc�����ڵ��dx��j�m�xe�Bɟ�Ȝ�^�W��)���l��;����:�:}�Q�j�߯�c�k��;U_�Z��at�EY�}�Ĵ!��h���!�{=!^��$�\NGy�fd�{yˎ�Qtx��j8Up��n�����/�Af�	�
G��b<4:T�ճ�L��仫�ם8P~����[(�e��P�vڷ�������)��5���ήPr�<�2��X��^�:c�ۣ��9"���g�f�Lt�]����S�M�O���c��޻�:c=�޾��������v���z�f�o�̲�~f�N3���$c���a��b!���<�nAz��X�d��f<ٕcy�ں-"h��d�ܯ�{�rͽ>7��!C7�ݎW}(�
1Y�Eu�x�@0��+Z�v\��(�)���ܕv���.=Pw>�3�di"�|��~�c�y�#8�w��W9�I�	O������u���l�c���tT	�B��P��z����:ش��4���5���;7X�F��E�w�2���i��xQ�X���".�H'ޯ5N�e�	ޜ�1o	�fg��/}��׼l]���h�=��B^�zfJ�[��A����&4�s%r����9�{�z��c9X��4�u���=8�W��`�y�'[(1���F:
��¶�U�n��p��ݻ�A�.���m��;v��+l��2��<	�ɚQ�����8b^EvX��U��_�Uݼ�Z`?�'>�����N������a��v�	����u��
�<c2c���Pl������,��D��0�)��9�����{�Ot�a/,}Kw���L��7����%�X��u1X}���W�в|19tQ�_�����hR�,���*�cg���z�N�/��)�-��"�j���,��b���'c̃���M�uYmz����WU�������*��c��ȶ�v0yKK$8v���)�>��8ת�%~���0������a�$&E��q��C��aP7Flʰw4�4N��L��#
��ș�1���/�賱�b�'�o��5�*��;pqQû/�ݳn�����թ���Jf:��f���,ġ�/��;�J�ݙ�����e��v��;9��?��$��=�=;�~0:q�|P��R;$M�L��t�!��
m��U�n���~����9%�ǦT��	ӈ?Obݮ/���OA��J�({�R/��y�b���������5c|��#-o�ʩ=�虌3���ŕ��9�z>�'�a0F�B�B�*���u�p��<�a�>����z�%�ac|݇�������="Xb}%z�� ���P��s���&'���SU��uݾ�lwVG2�
D�/x���u_���ƈ9�=5��#��\�+`y�	��K�W�s<�E�s	?��@����^,��'*�T�3$�w��ςρ���X^��pߓ�f��������{�XČ�zv�_���e���X;�24�@����x�Ȳ�痹�ԇ�k�!Y���uA�k��ǟ9��v#���R7���Ц;�Å�~����]�o��"O��OE} ��b��=�@��Zݏc=W�9I�.�����6����)�f�ǜ��_���A`p�B�E���ʄ�_t�w��������=;q]�k3�h�M�6�;v�/�a�=X�57ζ
GB�՜�!�rт��o�]�d��v]_�۶���,b���d�4�0po;��L�������&�����վ��P��nY�`�7�To���=[O��]�*er�'���u|�N�;�ؘ��6��S3Z'!_�# ��$�aH���M3�",��C^�s�#_�����Y���'���]������f�c���+�dDx!XVw�����]�e��gai>���N.�s�G�^=�����XF��[J��P���d~�.��L0Z�ALe�3�7�q!��wH�^��>���x=wQ�z��ȱ�,[��izrMEINşꟽ��'���n�~���>���k]l7���:,b�{���Ջe�!���-�s/عA7:�?:��7�b� � �"���������9�b\w���*=ً�"����޾�}��#u׎��W@q`KN�d��㱸e���f���`�I3�!;̏u���boj�ȟ/��V��f���#���d+p$�ǜa-F���[Z05��~C����=��]X+}n��L���{��荽����R{ƙp7��E��7�{�1֥YQ���A{�-��[�З^w�d
qtJ�X���-��X�ܑv���8�F'*�����H<c��=Oƭ?o���s;5�lL�Ű��r6ҧ�u�_S�i����W[�E�T��UV�{	7}~[^��"�Ş9~�6-n��_�C��YU�^�����zz�mC[ڒ%v�$:�;�n�N]n�n�5��u���J:�вTY�H8���|�p�騿�A=���;��G�tה���M�O7Pُ!�N�܌IҢ��=��[��d�����[&�u�o1XX^ �A8O@_q����ף��d<��	u>4��2GS�-='?mo��`�~xv�tj�_�e�Ӡ ��s	�>�4`���Ǝ�ά�J;*��L<�wW�z�VG?�;�w��U}ޓ��O���G���0��h��>F��7#؞�뫑y�;O��Փn0�Ρ���${��`r�o�����Q}�L*4L�T]
g�j�ך'����k��g'���}�?|��U����iK`�v/�p�b���3rV�f�Y�Y�M��s�wE5���ѥCS����9�����qgR���o�ƫd��ElllLK�9~\�Yj��R�3�0,>��Z����T�ַ�Ɯ�E)���z炧�cc�!QY����vw<R�/�\?y�`{k8ߍ�}Bɟ2'h��z�@��`7>5�(�R�c�zzfV�s�S��=>T�8���[8�V��Ӟ7���7����9����d6{p�@�����^m_�J�O!�O^p�Zz�D��0�[����ǯ��=�uq���G�1��!�]m����)X�2�_���[4q��B��;�s���q頹8B��-�ʬK4VY!�bQ빪ͮ���-�������=�.��@�@�:�Y}��U�uu�-����6��8�(�T�Ȱ��6q5W)�q�3�>��Y��r���y�7P&gB�6�_�ݧxb)�J���8w�q��L�|�2�>�p�n20Oz�4,�����b�GR���lԞ�V*��=1zbT��`5�rG��m�)�e?GW�c}W�s�Fm���)M_�/������AA�x(09r��uJ�vע�Z�c���o��<�˅�����T�f�	b���4�E�WWH=���B?>3�Ð�69a~J���G�v������:��[����sw�nWq����Óa9�6�#�)�bGO������{�I�yuP�,OYԡ�Lj����{�^��[�=��=ǘ_����+�u��'`�A^�c�w�����g6���n^k�z�a�/.a���<��8h��[P��3���\�9��c �|ذ�Tw��c7^4�Hu��>�%G����v��v�
��Xʫ�Ӊy9��<0�]LgEI��1�W���o�,D
3~�. ��%�P7nF�x;�G��
'v'YI��VnxN��uE	�N���pO��2�����e�&�����-��:��cf��yé�H��GX�GP��]����N�쩆q�/��|�9�5Җ+x�Z��LKK��&�X�����J>�HN�T���3�k=Iuwit�;��q;��#�܎.�|:L�}6M�Qk"갽)u}�T�Vң����µP��p��7���>t\yM�7�0���1��xQ|�����;����:��̨A|:�mvǨJo�l�M]�����rK�����Ӹ���Mu��C3b%;��*�f��[O���JW�OwL/S�'���9	�hY}i�g%]|�K���횕���6U�҂v��(:I�����h���徃)`>��P&�i輻����N�e9�W�G����=З�{nV�uS�I�u[d����BM�w7gZt���Y�zY1x����0r������ݺv:N��/A�7���|�������&���uB�\�9j����|n��Eĳي�%ۓNFҁ+��3�h1!{x����I�]oC��~ t$]t����n��������	��V�g$��L�]���t�a�Y��u+������7���d��V)���x~С�(�}��[@��<h^v�`�#/{xT%�4�*����J�(�En�|FA�N�O�Fxv��у0p�Ǿ�N�����e��%�[�Vk\����8�F��Yyu����7L������Sl�	wJ�e��)n\����T&6��QY��
���2⭟iɓټcْ�ͩ|f�K�SgX�&�������v탺�QqoN��t5��Z�#7�	���	P��
�xi˓w*U�y\�xx�
K�盗�U�MuC��N��UNM���.�1��SF�,�h�R��b<L��hE���jc4�5�ћ�����k�pʒ�H���(����Dh'l)�놷Ǣ;%e<��־¸l�Q`����0��	��1����b���:v(���2�Y�Ÿ��]Y�1�ו���|VO�7с2a��o;cW�"�3h�Z͑gmZ�2���cp���Z��u6�C2��!��;0��P�ײ=yi�7�W^��+�CR<���IQ�V����,�Y��_�q�mr捧��܉f��
����t�:��̺rm���.劝ډZ2mѼ�vܺ�bԝc�j�+	R��hy���j����pxމ���\���ܡ��%��w�[}�<']�M���I-�J�T�y@1�����z�8���u��6��Q����$���2M5��tS���W=��69�9֨���'r�:�E(�u��onw'S����-nL�0��X�ɗR��G]�N�υ��on�{0��U�պ+{v�G+r�J\�C�wa��MHToÈq����nU��w���z�81�a��M��G ��W�VfM����>π��l0P�F�ؓ�����py�k�fq5\V������$�sv��74�6���������]���z�2m���G���㢻�K�v�;�G*$WPf�#ͷd���IKލ���R�b��ڽ�ox�Y5��Ǐ��HQ?�2m'��&F�Ջ�9�Cq=+=*�Q[^߱&in�Kd���H����I��܉54�(��K��%���]HӉjd��	&P��J��ەu2�7��������=!q���z�dB����_<NOl��!摐�W���r�>q�{J"
3�z1�����i��i��HHRj"HVE�"��*�J��D\�b���g֛���A�,��ؑB�TI�3�$��SE�T�ڟ��Ȃ��,��L��gs�d��-/),$��(�<�I׶S25ĥs��E���H�"Z���b�R�f�ǽ���4\y�^�77\���k�4j3=�hVQ`d-��?4A"��ў�U�kQ��az!v�Ǵw��Y��&N�g��',9m2�]ז(d�]b��2��c�V�N��7��-μ����d7Fm`�
y݇О^i#�)�XB���ч�>��n]uףp�����W7V�1qcyCʰ�qR�w�{�=�p�>J�2=ϸ�W�,�
EW�O�MNVCG��+��K��v�������7�C�J@��qa<�"�j��k!���χ&F#��-�p=G��1=��tU_�ouc�*�v�r�[7�c�Xgc>����T;	��(���\䕄D<�O6f�/���^��HK&�C�����ꭅ>��8����x��S��/Jf����*)J��K6.�u����3�����J�Zc��]�,��X��;��)�e��[��4��R�4���ĸ��#��Y��"U��G�(!>�[Vԡ�&��S��ç��o�ץTl�f5�V�E��E�\�,�X���3���0}%z�� ��&ݣ}F%\�^M_��R��x�f`�7�0�]w�ʲ/�B��Ox������5�"C=&�#��A���v��{��mf�c��������񨱋)�X�
�kY�_����
z�=�^��Y������L� �����
7�O[�X��q��q�AYN�v�|��,��� ��A��x�ޭ��w�i�u
4[�N�x�ubq��.t����)�ؽ�M��u��j�~�g<��]���ܝ.sِ=��[���r�=��`�ݓ'����A �ެ����K��_A�Z�i�y���~��>SKH�IځcWC����
��v:,�^��?)$EY��q��l�ťZՎj�&+���+�s�[��Wώ')��/�N"+m�~�>+�u��S`�]MA���	�)9�o���+¶�=��{���g���O1�uL>ʫ���E��T���t�f�8 �
�<�:%�����T�6Z�xwEʦ��Z��z�����:i���DX[89ULP\'#o�dk�4K���|�	4Ϡt��,�~��w��k3�fV����ޜ`͎�	m�bS1�'!��3
�Ȉ>
E+��7�j+�J/֜w���~dR>����4K�����-�0��:N�1�4�術�.,uNIw��8˵~�E����z\��n��������EvUL\wڝ�<��w�<�o n֐E�cD_v��Ӱ6�����]Q�hv���������|eW�-wQ��X���r����g�2*.zlj�Ȝ͆��c�^�����u�ME[:�jL��ץ�>�����=B�����k+�_�dI2�W��䳆{H��j���.S9�r���,l��s5e�iJ��q'�U���u՞�tB�2<���o'F���,V`�>��x��.���^X\C���h2�ni�{k�Hu�ᨅ�lo_�?u8vʶ۱S4�C�c�JTQ����y�J-�R1�t��>�H;�}����;M��L�ۚ�A\�_�����zw�Y�����IlX���>��b�Y"҂�|�ML1����U&_����j}Ji����9�,�lz���D.)m��f+��;{rV@��(G[ءIz���L���E�:n��s���������=I�۞1�N�o{`����#a�<%C��Aµ��kے.�^w�qg���EH}JOFw��a�)4\&�x������kO�J����ؠ%	��۫e�W^��j�Г�F�縺L0�oH�ք��sN�D�vX�#,t�> �B�-�O�/OmMF����d<��xv���~��3/�����|����9nz(,���7 ��P �ØO���'W�o;�����}���&n�sC.��y���p���J��69UtZ쨄��0��D�)Ah����X_K��`�w��~Q��!�?-��M��dw����3� o�H[c�����Q}�Lzs�J�e`D�xIkES�_o�~�?��A������R�V!nנ9;�R�6�Hb�W1H����7>P��z&���b��¥���x��^�	��jpe��<_5��x ��{��ӸS������w�k����E]Jr=����2�`&l�FЌ3M3}.��lX��>�]d�u�NF%v�ʈW�x�Hz�v��F����O�9ڱ�]�(�u:���� ��w�O����v�v�Ч��a�B��Ϫ]�w5���j�nH���)M��P���W7�0�oI:'U��B-̐]�����1_i�3�TTPAˊ^+��:�߶��O[���I�����ɰN]�רP��G��p0���6���}"��2>�����~��`7Kz��w��N2]<K�����~�[�,C������V��Nx��xe��Ñ�����a������K���Kz���X�t>UѠ��ȴ����&���7n3���:.>����~I�M,�����ؑ(w��N*Tމh�R��L�|�i��EC�V� �OG�N�B�x�G��Ӽ�9�+O�#pħQcn�C[&��rE�v��S�uoѳ�)����:}~�kܦ6]@�c����= �49�m�<vc�d�Ʃ�����5g��r�*���%(�R��o����d:�g=��2{bPx�!�y�S�CZg�.������ޙ���������7ʗ����<둬r6�	�q���C��JH�u�2 �#�4?�x�vA�ݖn͸7�Y8�И�;�,x]��/,J��T�y7L��sq���U���q��c��ە�zĘ��~𺤽�#�d��[�;�o��C�[��4��Լa�R�}'je�y8ƁJ orn�(��k$�7|U��w�am�&Zh��ԁ�� D r�WOr��b�c�o�����_�0�l�ϼ�,5N~�WU�6LF���mR��`��
3�"�u�۪�<���cJEфw��[FT�>���]__`�7�a�~��&:�3�~38��ᮖ�w]�"2BvP���66����X=q�m��ʫ�����(�>��փ((˺��.�[��CÀ�!X����K����*j_��6�l7��Ƈ�����с����&v�����]bY���.H��q���a�m
&X"btd�-���U�R�߶�.�˯�8]c�G$�-�N㈖3�Y�n����\d[;fR�L�)_1>�59Y�[��������x�����k!�J`��b�!ń�=lF��md?pY�w�
G�zߵܕ8=
�׳�ϳ�,}u/�@�]�x+f�/�Xgc ����M^��=��c�\�x��U���&{{ύ������׈��M35VË�K�g��~8�e�U�n������[;��
�����!g�C˜��}�}�LFdT�b���p�K�z4��l��f��y������T~��FJs��f_��` _r�^��-��K�С��[Ϊ�-s]Z�h`4��ʬ?���43Үd[�j���A4Ny�ԃ�Z�E,����7�{���}���ʒK�K�RgF�|�.&w	&�mfз���v3���ܜp\ɱ�򪿁� `�OW�w��ۅ��=�*���@�� dyɗpaw�t��2�f�/�����s���Vi?��Y��|dt7�:��a>V	U����	"��Ha���%{�B����c،xO�&�6�Ա����0�R��Sp��
GE=�Cmu_�0#"�!��trt㐼M��k����ͣβ�-[n�^�Ƣ�Ŕ٬�:P����Eh���8y��	X�j�����ZHs��r#aq�s|V~����3>Iځx��g��`PG, ����&*;���'�s�����9�qC�~[#&+���1�sOH����r����ܙG���K^1�پ��oC�!��R���"�Cz8H>eX��{i@���ULʅ3+3��j}�/w��:��&+S����t�EE�+ʅ pR��_�gp�z�!��Ǟht5�k�s�[:bswEqb���[sH�S�yL�%�r���eN�A�"�h�"^��B��S��Q�X��n5�?���k�ޜ`��P�=�8.�w^���1��ɷ	x�U��g��/��>��r��.1���&{;o�BT~�hg!����ct�{ϲ�f�l�8��,�/#&�ӓ<B���G]��D������AڝIn��m���=]j��1�Gv�$鵼��$�k]w�������S}c&�=>ME�|?A ({U��o�&�o����ޮg���ӑ�/Ƿe�f,b���Pb�k�g�cӸ\a�g���x}Y�������&�c�α�gP���K{�}���g޻��"���yK��
y~��1)Or��D�H�KsøYr�/�u�2���MXW�xC��q���whs�����=2v6�_�o� _���=�b�S�o�f��V����_߇��?!<��2Cb��������+����d�foCȝu��ރ(����N�d���zw�Y��>~4$����H�d��{诫��k�{��Ѧ���򿻦[/�3P�p#�C�ոzo���eK;��=PN-��5Yy�P%�y	�@�
�N�ǧ\�S�yx��}Sܽ��Vl>,^ٕx��/�R^�2�^g�B��5)��'D�u��P�|��-`[nH�����g� NT#��v�b�7�y]�m����C3��e�������ji���Zն3>	;Tuǒ똯U��������r�(r+�,#��$1=P:~�Az{jj5����B�����~�@L��x�^�݁{t7V���r(��\�}�u:O{����-窲-�N���� ��C�v�D<�fc�u�z��vI�k$v�#�����.bᏕ[�C��.��?�Z60��m�/�p<�U0׻��@y�~�����R�kӺ����V:���]Bw��:
��'��� ���N��P&����M���o�_�ь��s��r��L�Y�	Wզ�*��]���8 ¯����H2)���=Y�ůf��>�ZWw0�Xݡ�ަ�(?J�jq�9�&�yZ�ee��*G���}^�V���m�@�2(M*�sn}�� ��T7o��	K`�q!��Loy��¢�s|�=>��Pm�G��ܞf`�	QQ_!�Q@]NCg:�4��]cb��z�u���d���'�~_�+u�K����,1��$��68���Pg����c��m�Ӟ��r�H��7u]K�����	���-5��m�7�]�&|ȟ��z�__��C_C��o)^����g/:Z���1o$rB\bR�(oɋ�qڭ�at�����3�İ��Nڞdzd�e��[վ��S����C��>w���do�MCgj�Sv�	�z}����BV4+�V���1�z ���j�K��+!
�\l�e���[�	.��^��zuz���D^�*�1�RK_U��1M�_LO�H�[/T��8���1�3�P7{h�����fF���V�w�0�E�s�f��ڐZ�N��v,<�^5�3��:��/�V�8�u:�fΑ�v&����,_��y+y��wGb3�|-���X�ߦ#�B_�#v��=[F��rE}�n�(�e8u�.��*�
Ⱥ�/���=��P9wk�ZKy�\��8pr�7+v�����h�]LN[��A�Fl�1K�`��5[��]o�h�����F��hsSP'ˠ]xG��~|Q��,lp������vDNR\�2뚄ǒ��ǴѬr6�N{��|H��)�c������Pq�͐[B���ݼ���Q��n�q�иV+�f	]m��,5����]TG��&#t�����o��q֬�]=���$9�b/I�Ӻv����n�r�_���K��)OP]cu����B��ɮ{���b����JAC�f�����Mu���'��qs1u�Ű�Y�-�a�Lh诼�/��Z�wŊDz�6��*�G�
����{|���`B�䏾Z-P鲫��24gAm��z���^�T�mL����$�����Z��
]�E�c�"rU�A�c>j"$�ܖ�_��x��:!v������B��+��}�E�,��G����Qc[vTO�ymZv�S۔]aq��s��������N��z�[�����>���%k��M��w������9���=���g�V���E�p�[V�^��<�
�0�;a>��z�9>�z���i���}ʪ.��y�sٰ�x��AO�o�w��5�����9_,t�&�+�חV.
ӭED�c�C6wk�T��1���	y@D�
��>ߣ�yiX��-�J<b��T%�j���b�0r^ڼn����!��H�lV�p�{��۵�;���0��ce�����Z�bW+��}�/ý�����f���B��LU�*��V�s����y-��GS��u�z�e�<Xc�H���D�v���i;=�9�F*S�I^���'�2����T�(������ᱹ�v�k�[*w(���{�w��z�u\�Y]�n�y�իnS�!n�dI{됥�yT�=��Ȕ wL�>�ﺫ���V����@c�sS݃|�<��Ml{/�����v�C��DP5����ڭ�y�=����+�հ������k>�x�1�j��RWNŌ=t̹��2�rÊ�����q٭Ӑ��5��O2�I�����t;F���ݙE`�c58l�2�?����
ᔷz���go��m�*gn ��.��ބ�I�]�ύth���X/�o�N��bP�}��v�K�u:h��w<r���MQ�R�
��^�e��n^������LǾ�����*�j��ʭoq���Kì�;��gΔ����L;D�Yt�\�*:��@Q�Lh�N�vŭpd㚖�D�&�n�U�G]_f�t��.��N
c&Ǣ�.əT
�\�0�>�#���a�SMs���}��wi�b.p�bvQ��/����%m��_R]lT:w��7��v�_r��u�'ߙ��"��w�t�	���vg�"wk���f�X��@Ӻ�H���cs�s(m�4���!��fd���л�&�߰��n��%��K>�;�B�$���"{6��p%�v�\��� '��r>�+�s�g��9Y��̻x�V#x!��P�j��e`G*��7q�᫺v�6,�Ȼ�P8����/LǙ3�ɵ-aűҫ�re�IK�N=��c�����t<�aA�4�2E�E��R���s.w�nc�Rmڝ�P�����In�k-S�cI�jYԂͼ]��״��hkt� j<tD�����Eî��Gq��\�M��4<ivq�eZq���%�񖇯_wO:��^�h�nL��m�rjII��i�e��朙.!�_v�wL���ٟl}�У�v�{JJOZ7�� ���:J�x{�o�]s�V��ԭ�}�������/q��V⌙B���ھD�Y�@�y
Fyeb��vu�56`�If��}��l�+;xՁjI]�����YQ��2���/"�u��`�ͥo���͒�ȣ�6�}vI`�ݙ�*k,���u[��o�MI�u'gOܮPƢ����cS.��]}��Vh4oqs�z�V>i��z]�T(q�^�I�yn�z�*�����^�fZ�FF-y��N��7@j	�!�"2m�(54���}�t^Q-�d�-�Ker�����̈�N���*ڮ թ�-�	wa뎚9�͠s���kY�7Nf)�Ͱn��|避[��ͻ΋Z��-�>F������f��ۦC�e��f�rOu��M�xk�wM��[V�̆�,]l��5��xzT�`�%1f1{�b����Yy��gX�X^�YP��7�p�Oh��5������J��5�E��4�X�y,�*dֺ[xa;
ӳ.1M��c�{_d��m�T�l�'�iٮ��I�DD�S{�hDy�o���c��ԡQݾgg+�C�=�Q�g��_5Vq��a]��	����"�"1��-L�/5}�p�`ܗB��Ji���"��M�^n�fT��cg��'�V�h;�f����;���	xt�ݜ�IԁK3�]
��[���G��RБ0&=�x4��.�$@ ��&�� �R��n��� �b��U�EFJ��T{\]���=�#�lC�������9�y���QD�QQ{��F�ɶ�7�j�e��a%�J�n~zG��������$��	�!&TDY���ҤK�NXE5�¼��p�WE=u�Q`������d���%_�q�E2ṩy��RTI�V!��Y�Yf�U��Uu)UrJl\�.Gթ(�d�cۮyt&.#3��V�A�ˆ�E�fJ��UyzzT�H*DAn��AѴ�]�+�:��2�$Ty������VEea�X�5��B#�[U8�T�������*'�.���#�M>Љ�J���P���r�<�vҊ

"(��6��jRe�bT�.U4d��J+E�M"�<":%QA�j�(��B�ܳgiQH�F�	F���Z��쨍E�e2#	X�۪5���j�͟+=��wM5���}�A���v%��؜Д���/�E���4KB":B����;�`L��[�;��>�Q�g+��$"�v�^}Au��b��B�7��4}��%��q��u�5�`^;����e��+d�N��޵��0@ࠏ���p/�]c�+��N|���v�w��Ϣ��}��3�<��?E[��>����5�v���+KQ)��T�����ϻ�H� hw$l5��o�����[�jkM��7��!N2dh�"�3�
���{���`д�WܭQ��~����vl�VM����ҷ&�F��Ppk���u3�Z�U���T�6�g�d�X����$��&bz_h���C<��~�*ˠ6���0J�����>���^V".�ފ����zb�g��i�Ʃ�Ζ]��=C*ʫ�,,���X���Q��N��3����)ݾ��7/��_Hj�j���ܴ�ϳ(o��C��m��.�g�T`������f�H,p��ñot���o#ir����e���B`��ճ����V;i�򵋒�9���t�/2e9� ��G���l(��.e�0u��i[��:�s�[Gdhd�2�{�6YU��\
-�s�AXi��s���>N�hs p�ĉ���\3te`�.�o9$�"�8���7���ݨ���X��۾�b�ON.��@��>i��AP^�t��ܤ�:i�N���U�y�L]/gd����J"�J�),����6��}Iy�V�*�ָ��G
��9g�Wxc�<��3��|�?-�����z�ڤ�m/�����1�8�;g�o_���we��S`Rݥ�:���� ��@��@!�l����CK���x�u���4_���O�t��ϭ4�n��]V�=C���9_�Vff�<��".c+����^�Q�ߕ�K]i�='3��5�䍃�8�Z�[���P�&1<�.�"a`΃��=C���C��X�!c����yh��/�^9�~�ܪ����z"�}0G�r󟌼V6�����bs�$�N�&���B��Y�4��5�W�Nl��z`�g�1O�+ά�KsG����.���+�Zx+h�o����c��}yn�͕Cj�:hW����޵�����+YTE�o=xs �qM���ǛxHb[I�Uz��d�Nԛ�%u+~AhE��^���i��Aib�������%
�c���Mm��[B˾��[�+�ΉF��s�m1���W}���(`���Az��}ͺ;�EL=d�zWR��\�]��	<�X}����3�T�۴��{m��y��04��q����+����˪��b]X^�V�W��w����b��[S���ݞɢ��1���r����g�W��(	|���|��j5�Җ���2ҭمwN�V�͈���^��Mb��;C2%�ބ7����6[X8�V����w���Y�7��'|=9U�8����[[\w�5�}�u6�����,e�N���o�&&gA^�������+�k�+�߇��̳*���g�,荧���b!�����}�~*��k�>h}�����s@.��S��
�ޅo�ɏU������w� 2��׻n��.���O�����z<��լ�/^�����s�3�R���9�T�^67��>�O��z��j-�l�����n��r��{�l��k�� zG&�-��h)O�#�R��S�R����S����@P��v:;.�Q�1؝�t��+��	���t��dNV���3�V��5�؎uu�gL�\�ܣJR�.�\�5����q�S����M��[���h��վ(�l޸�wW�K���/�Юۖ	Y��,�ɗ$̈́��osr�D������F�����#��GyF���_��66&އ�8s���k�45q<�N�Z-uy�蓣��� e�R���/�,��W��S9{��L�K��J9�Ih�]6UL0���e�5�'�:7��,�y[��k��'wpJ�m#"ױ�����ξP��p�U�{
���v`��_=��S��>�l.�i�O��z�c��[���TO�3Ry��W`����)�G��ަ��[��f뵇��9K4ע���`�a.�i�g���9B��,�pK�3������<���(��SW��k�o����ϑ�G����%�DR�"^
܎7��᭭����=�;^į�N>��3��V�	\��{����M=%�������8k�Ƚ�/���%Lh�ºuv�����:�|��=}Q�V�bb�ͷi��]���TEn�I�F�]��&��뼧m�m)Z��y��Z����
=�t5�źm����Hعý�聚���8]^5�M/�ԁ;�P�g����� ,K�$�産J�)�Ǔ��.�uۣC�\*��S��jXE,o��v�5�����vYAy�^g{)��O�ׯ�u0�mˌ6�� �Wvv�IX��^ֵ�خ�y���TՅY]w��Ϧ��nl'�@.�|1���F��ۺ�+  'a|��dC��~����U�����>v�T։�Ǭ���j�攢&��Վ���@�7���[+�ݪ�/4�̪�9�u�ے�vɕۙ�^�}47yW���k�X�B}�4(,oIh��U�B�:�*L�v{�\Կ?���<����'܎�v�V�B���ࠏ��c��/he�OV��;;����=��a*C�,�ܤ��vj´��ʗ�2-��;�w��m���<�=�=�>��5�ç��b��HP�FO��癒h��>�����'N!n��1H9�િ_g������h�z[j�Fz*;�t��"֫үG�������Pp%����ZʯW^UWy��������~�;�4G1��t�q��EB�׽o�;�^���+;3�#p�UB�|�(��;r�E����X�U�FreB�����l�A�[!�n_r�����u)*͜�&[7X�g�o8Q-΁�ݢ�xmM��xs�����Vqfh��-a\�mtNLO"�֝f'�	�>�����]O�.N(:�����׭�<S�5�
/�����l�J��챼۱�S��anz�ʲ�^C���֏{n%{�|ꍥ�{���C9�_���5�q���7KN�����.�"�O�����W�n�ćzϐt"PTd1#s��m�2��J�rv_2]��U�O�&\#�չ�yn�$p�<�_]�\
��f~���:i��u/������SJ��&[���+����C�x=<օ��k��|���j��]�Su��k��Dp��lv��jH_-��:`=��{fS�V%��br򚽩�ɗy���� 1oK1�9���Px��d
�1�~��Hz�k���'+��q�׳�쮽����is�	�sS�t=Cm�Q��n����n���˼�U� ��ٽIڑ���u��yu�������޼���\�p�i�[��ˈ�>ǐ�.pX��^h�[�˲t���E4��Ӯ=B�2�%A�u��:������d7މ�ּ+��;(��A��K�{z߅5�1�Vp�
�֥ӻ��ܻ��7JD:L��$Oj�50f-V����k�G(�w��<j�3�Me�Đ�B���O�w�Y�A���X��V+�����oy��z���B����rⷥԫ�_�g�j@�T�F+�	Ώ)^+��7��t�؜��6;��1o=+�v���7�j�Yc�kɏ`���=^�?��T�oVm��o�����24½��f�wD���7�4�U�ݛ*�������S�jj϶v�o�ｫ������cל¥�ݦ�+�m��/�+���p��+;=�>����wn`�u)ތ����N�0�Ra�:��]�k��U��{�п\�z��O�������u���z5��*m5/����Ժ�z�+�U�Ag�߫Dg���� ��҆TKN��B�ߣ���2��(;c<7�5�;7� 4�������u�.���2~-����>�&��5��1\q�-�ʪY��=Y[�a������t�rX�a���1���L ���.�ԩ�UAk��� l,(q�H�Ǡ����8t�a���^���₽<yv�k�����=5�l�7�1o��-�����S�-�h��R�.�O"+.c�%ۜ�o��}2��WMf& ���%hUƩ�Fb�8tL��p͇^���� �痠��~����_-�������<�@|��k2Fm��O\̀t��zv���i2mW��tw�Mi�	�>�	�S ��۾��&�/�Kߘ��e
Q�e�����ҽv7�1�\ؤ�+��`ML��3��^���!���k�w�4�>��׷�]�ػ�/.M�Q5���7aQ�!s�+4$�Gk�߶K�냞�p15ѻ�w���F��k=��I�x�a�'*��u�!�Lx5&^/J�º�E�����2uo5k�A��ݙJ�P��:IE�4VLΌ�>�y:dP �6���^�p���y�Z�7G%�;�/G�Z`������c�?#�(K��t��H�!�]�s5��vϫͰ�ba�v�W�vZ�c�u���۹�R{Ҷq�;yz�S���Y0#r�s��>�����[�'f뵇��9K;ܕ~�c'喌����l�{�U�:I>� 7s��<�V��������	������V!ݻrwAu��	����'�Z�s3vlSC+:�p���XgS�Y�'`�"P�.M�}��R�֦gj�B��>�Se`�|�:)�S�;� ���"/���G[�6��k��c��쑂VW�3������<��f���g����E�ާ�������^���á�����\��ح��r�VVt��rd�X�D쯣Ϸ����i�exr��>�-��H�Ǥ�2�4F�1�����������y�5��ag�Io��M>]ǯ���*�y�8��^�p�+�Y����f�E�#���U�w�����MՍV�g�ϫ�v���j���3=�A�R�]1y�y�f�۟�2�����7\��mSs��%�Q�T�0��ݷQ�;���MW��v�d8�9C͈2�6nl�W;U��Oz��8�o�#�Ffg�gk-h]����6������ހ����o�[B;��ωٜ�yǗ�w�>�"�wc�M�:�PV!O��hPXށ殧�QTP.�n�V�z� _��}a�J�b�?^#Nc1�����X��^Wf)�m��MC�̾��T6|*�ZC9��y��h�;�皱W�v��@f��n�^��x��D��%�Mok�f��]�U!]��.Mk%<��t��mA���ДY��ٵlN��.��5���#@BS �z�Z��aK�J+<��xvd�bӻ�Tɷ���2�t��emw4���k��ή�A'{�g���X�����4�b�9�b�.�Ʋ)A1�jyq��(d��L� ��n,��b�pA��Ip��m~w�Wl|�G�������vv�N�S !�jsϪ����{_n��Z7�=�P�����%0wE������U��P~�[ `o�ޥ�W^Tڨ�N燁�L����B��\}n��}��ǓEl���
�u�>U*��N+�kީ��1���j���ϰB�R3�w�S��e���U�@^AagE݈�9.}����}�����1�<�����st��7bZw�����L��gU��*	ϼʕ�����BJF�W�S�Տ������Q-����'7��]��4�EZ�]׭DY�P���Hѓ�����T�],f~���s��'���>#(Un��`��~G�.���8�,���sk����:�~k�H��f�W�nռ����3pz8V�Z>�{�z861t�p�R�pnvU��*��]�VN�KE̝e#�!Vz��ɠ����33Y�b o��W�ѾF���>�B��ݔ-oeL����H�5����"�yғMQ��u�m!�(-Ad��;S!�tu{�;�ڗ���mŕ�����$�V��7����MfLc_שܶs���aT�U��i�����O�#��	���^w�>xD�ʗgC�8�q�ִT��ˍJZn�B"�'7l@�����%�g
�C3Jd��{����M3Qj#n:�J+++��cd�ۜ.��2���;�rR�*�6���M��v��"�^�x�R����,���b.8P�����&�4����e�J��
څܳ{�Z��ɔ�he��E���C3���OG�^��j���d /R�f]����}� �K͚�޾�E��9f��h�hd�:�����G0tڙO����<��/.r��	$�,+���]�(�ѡ��+��>���=�����(�j��U�s�->C�B�.�3o$���:)mZ����t���U���uV��xXf��BҪwa����I���9w�Z��M��D8s/�|����p�UnP�k�x8�1GW��<�;��`�i��_Uڒn�wjnV�����4����Uҽ�'������S��`�t9�h�w�ׄ-��F�i�'o�'��yR�Hf�x��NN��6��W3��Ϊ&S�-"v�|�u����_Z����s�1T@���	m��7��*�v,L*l���Uʙ���o ��ަfXG2DD�v�t;��Jnڅ�'5�ʹ3:�B��Ս�����Y�s���w[E�#��Lή6$��r�yuµd!�P�,]Lr�ꃏl�p�ۓt�C��,nb�:Q�⡬�Y\{H������S^M#��GZ��q��ʓ��%@��[ި�M�x��A��B�OTB�'Λqb�]�,M�2��]�]�|/�Y&��F+Ŋ�r����T��)7.l��79!��L�y&��#�=�c��hH�1�ȯq�}Um;��t�*Z��-[��R�����ݧ�Eؼ.Tԧm-[�{�U7��r�y+>�­��L�;/w��0�_�tP{lj��)��)��ex����b�N��usf;]-N��Y�(���8�07��m
�f��V�A�e������-V����r�Ro���T+�:7R�t���h�U\��l�]�z@n������>=`�I([�#z�k�p�^��Z]*�M�@ʑ]��>��N��t��|��:�}��+-���5�:w�{lȄg���b�.���q Fh��+�l��'Nu��v���ʢ7{o���K��aU��:cBSoa�7��l���~%��{{6��֏�AԮ���R�q�n11���v��wӆ�ǧi��2��@	5v	�{ާ>5yR�������1KOQ(�D�"�=u7DM(�2�s��^�^G���o�H*(��iι�x��?��!�=�T��%D�ҋ���V�QM�,�Q<�,�j�E6<~?��OՆ^W��E[��^y���Y�H�gWL�,�HQE<�g"�EW��
/"ʌ@�<�]=p��Az�F��(W����u�I��D�W��DZ�j��C!%(�Hy�0϶9�*T�{	
+�,�JM��=�g\N{eh�l�җP��	s�0��f*夡������Q�&UF����ʐҶ{bU����IY����
�BL���(��2�PB$��Ե����(��J�$��}�̯+#r*�
�	+D�C�E2�ŭ�W���:e.���UxZ[$"h��Z��g#�-_���݃ߔ"u�T�O;&��yzY�F.m�4��+E�I`X�|���}�G{��kt�ѝ���e3j�̤r�����5�_��-yҩ��>�ޮ��|�5$-�}}���[T�[�	�#W\0ߢ��]��׻�a6�EouM����)�����m5��fw`�s&7o������Uް�Z��y�\��J��=���g�wټ�D�?e=�i���-$�b�I��O�}Y�ݩk��X\�lr�]All�vJ�,Z�}�5M�^n�V��N� ���V=AＣw��_��!r��\mí�=}1��c�F,���~�'�-|u�}$���?V��{�����o?�e̃������z�שu���x[��VJ�s:1O¥cy՛hLO8=�5"N�>��qFuV{�нM[x�|�1"��l�T6��2�q�צ�T�q�ѕW�X���\˟?��+�M�g0�e�i��m?eY{1�ٗ;�2"�A��}���_��>�h�؟N�0�Ra�Τ���]���{�n#,���0����o����y�&�Y���$;M��,��}��ؗ<�F,���N��z�2@Mm��N÷�u�3�&Ż�<��mǼ1ե��5n�;Ba�9� �{�`�4��c*��	v�8h8`�g^�gr^�\�C�[y�f��r���1��<5;���{�ߩt�(���'%M���lH���&3kٻ�L�|U���^^D����̉i��������F�p��p����\�v���v�wgs�2ˡ�Be�����z��.~�p�6�|����d�(~,��秩Ovy�Kʣ�;�_�1�
d֙��%Fa%�>ywu_���V��dv7�ʟ5��{�k���GL*~��ӷ���~����ht�t��c�p�>����}��z�S���,l-��Kb�W��������ӵ��R�թ^���cI��Q^����^��F���_@ѿ��9O�kU�wb{��������i~���u���$��:^	>v�zz�]c`d��0�cp�[~����V�ly��0��\����ը魭@a�7��]A9T�u�X�#��:<�e��O@�qU����"{V;��m9*�@�F�'��WR�d:�����k��PtS��4�K���i�l��B ��J�٨����$�>��.��[tԷ���`��)�3�Ѧ��K���Yv䜞:/=�VW֝:�F�O1�Q��R�+�r��=����yv�nwk��� c�+����rI��t�T=0~aK��g.���^�;���g�Rs�aVz�7\��؄��HSv�.�o��q鷽�m�n�`(��O]�KD������W�����l+���ݑ�f��Ǘ��v��sօ�>�P@��8������w���}����,���q�3z��R>��c���~vM��G�0�~�������=e�Y�??{��5w3�o�j���\��W*N�=�t�yy��9C*%�y�#tTz���PncB���j|��r�]�c����A��m�U>�H��~��ջ5��.����J<�4����:^�ˬ���,��5׾����v����x0\���g�v9}���MՍV�ds�x�vq�b-{5勔E�J������h��]TՅY]}���^}5jۚۯ���}����4 �%:�e�A�d�o���geC����NՒ1q�3ӣ��2�ڂq�(�-a��z�ˑ�5�F�HfN���^V`[�ڮ�C}���W��K�lΒ��KGV��ˬ�0t�,'>l(j����78-V����P	�a��yl��RU�}[��߲�}ޏH��d|�uW;�VZ�=뎍��T��g��{�s�����6=�Ya����~c���?ڭ�ڴQ5�oM'�����}��ܼճ�+����o6���T!g��hD��팏
c�7X�{�b��G�/s�Zڶz�c�Q>�;�ڱX)
c*�T��~��6t�{۾}VD��8=����^������O_��{TU����w��+��bjd�]��=8���GR�[7����� }��H6�C� �����tN;�5��U!yJl����Rn��U~��s��ld���2�=gsLӾ��@χ�-�!@w����@t�u��	N�}�S9�+0�z���8e�0c�@NE�O������`7��loy�ޫ>و��*�ͺ>�ݺ�����V=�!�>GOx}�����x�;t��-�d�X/#���H�o�p��ܘ{r��ڹ���|����`�r�h��ݹX�%���D��k�k�x���;��p�g��6M͆��	��.驰�Ky	4��[)J��9I��2t�8�9���Y�`S��ut)�l�����v\��8��t�Q��W�&�Hn��iH�6���&��N'�vy���V8�V.n����>́�\D���,���ǗV�V��=�D���x�;�'s��m����ߺ���>�.V9�����ԙaf6]�FY��Hᐓ�h%�/���I��·Bg���S]��F����Ϣa����6`Ya�I��g�ߖ���~�C&z��fO�s��y7���پ���I�<Ԑ��������*�UwT|�XgGywoM߼�����m&��F�[���!��X��ϣ�U���$zFϮ7)/v��n��u\��[�)DF�m{�J��=�2�����U(l�C�ȱ7L�r���lp�Y·�o�f��
Z���Z�[c��\.E��õƞ����ż"������q��w�=�Q��ڂ=HO��;��T*��z*�\;�*'��oE�b��S��~2�^�y�ý�W`B,>�����t�Y�3q��g��:���Qψ�Y�q����:�X�&�J1��}@uw.M����^�'���RXr��A�����޺bIce�i+2������!v�j�	���pN�#�ok'�)q^����Xq��;{&f���v~������=�OM��?0�X�"�q�ng�~�`kf���z{&�ٓ�=��m��1"���*��`���ѷ��1�O7Ϻ�V��V߲���������,��&�+�n�ʹ��F4�������Ʉ09÷��޷+[B};]�?XI��r�3��O���%^=<,��ѵ���B%�lV!C�]�h�����WYz��)+��]�_��#�~��4�aUyHD2�Љi��8H��̇{'}�b�z�z����"sW�`�_ܝ�Ӯ;��e�Z��2����x�����b=�O��.S0�s��6�7��(�T��������Xc	�7x�s���7V���W\6���،���_ܭ��_���vӚ�fx���ϱC�;]��������[T�����yU��j��)�p}�z����4�T*R����c}�]�AE��K�N˫=]�1+k��eq鵵��ت᫧��E�vI��(��í�[�7-)�/wE>����|�s�5d������VZ$�y�#�u���]�r�)�3H�U���m]FXAM�������r������t;�T'k]�+V�]�.��>�]�wW7q������%(ķN�S��@C�?!�$6���_�jS��9�C�Z��Y�7���Y��Y���X��,��F������{�͊ݓW�}��<&Z��fqfy%-����NU=�]b��DR����w�幻�^-����� =O���pŉq����\����T,����̏A����z�d5��][7�f��b��h{��g�����u����o�{76oQ'���a������'�o��Ͱ�:bX̼����pMZ��,�*�v{�P@��������.��Su�k{��O�͢VY���^����r��V}sEP�`+�&xP~ib�Rx��9����;+����PYԭW;[yﺬ�\K�3̨�f����+�uu��C��W�1pG�#�.��ي�|mة�=�/�P��##��^W*��k�:f�$�ep�5 0��-'uz��X�Lw1��:۹��_��0�'���Y���k�����@�o3 ��]b7�y�*�0����4��^�N�_�{x�{�}��+;F��#-�M8\���@o���FQ�p�>�Kާ�}�;��`O�7�Ӯ
�z�Y�-.��vz݄��F��K+���8�E��nE�wS|8���
}[Huw�`x�f򛱪�!���C��]��]\��ޘٓ�ӯ�����Y_8>���^���׫���5�m��ٓYlF	���~��i��%�^��@�G���G^�̧��Sx�����5�g)�����zo{�����9�{����\��oL�>����I޸*%LO��rŵO={խ�����w[�)���xp�s�OW��O{�.�C�Z�TкD{��TnW��j�Zڿ�����ޝ���a`��uu�rv�}��]�aH�<<�
�M�U�,�?v4Ҕ9Gb�YDxU^�I[1�w���ԭ��s8=�e��ߚ�;�O��#]�
���8���^�Ab.��Y@2]�9|�]�+4�V����V[�MgK�U[�0N�2���y/e=W@��է�,LJٵ׵��N�Fb��e&^Rrl�K��n���{�L�v��͵4��o.�D�̩��:�/Ix�Y3WI�;��!�F�n�Z7�����񧨷�r4�U�,bυM�cj�}���.m�g�I��<O�ە���C+ޓ�W��|h�r�t��O�iқ�~�7���.}��KV�ɺ�w7�����m���ʲ�mA���\}g�*��ڤ+�UW��չb�T���rgO���9�k�)�~�B�ʆ����p}={�띝�����K��Wg���}C����7a5�����e�hsꨯNk���4���=�Q�W��0�d!;�(��e��G�����qU�;;������_P���l B ����5�~X�K�nǲ'��5�%{�j�˻c��|�u�ybպۃ�Yj�K�<80X:`�/��{����?�x��}:<5�l��8z�J���6`g}�Y�O{�a^���X5
��X���]ϧE�3\�V;��j��o�����78�6�ݔJ�����4-���r�t!���ӏi�S�f.�߼	��A�l��[����V>���]0������߱���Չ��.��!�e�|�� ��l���8���r�a��M��Ԇ�����!_uX7Pzd��9ť#��u���R��۽��Cg��qx��K�T���B�L{ݒz�P��=˰�3l_�D��T��WٽnԽ�>^��:�{��~	ȕ���Y�����I�kذ)��
I�U����F��5�\]�1�<��½���%��=�S�E-� ��a)�eb��}��x�r��w�7�r�4<���ٴ�	�}���t6l�L�!��q�7�.W^T��v��y�ǫ:��fZw���1M#"���*�Q؊��}t����~����s{�2n���Ӿ��klP�aWܭ�Ml{i�1�?��k����v�M�U������޷�S�Ϙ�Е��	0���z#�l��d���{�3R��cz�U��b8.X*���=ٮ�Ǵ#XN±���Lt�ߕ>ؿm��u+T���+^B���e�ӽ�p@}����=��u�f)���H� 7��Gk��:|��ʜȱ[tk��ݬeӍ��| +a]W96��ˠ-�����ggN����ó:Ц٬P���m�E���Ke��w�0���v�����F��N����:%��.�<R^�ȿwׇN�0��5c���a�`.�*�[��lu�"�r�5�)���ɝǞ�/C��҅�_,ݮ5�b�N.�P��5����B�Ŭ��.^8���б���n5լ�'VfcP]8y�5}0��T2�W�V
��n�.}/Zѭl�!R`�C��hD2˛�*/g`�%i�P�w��}��Gt-b�[|��~n�^1�g|�2j��C]�:�ѽ��u|Eeb.�K�V��aH;V���#wou��Ϡ9�>l)K*�Bȸp^#>pT�p�
H^�P�Rs�֥@�]�IZ76���.-,�޽�������{�u���Q�F�a��V��o3�z6aЋ �z���>����@��z��m�������>�7�z�c�1����C�B}���[ܼ���	��Y]�z���Ga�
4�����0�rs�NV��A0�㋔�Ec��*]���m����m�����4޻�����iA�m��P�Ki�7�˫RY5����Z6΂�-�
��@����0k�q�r�Q�m�
�ޮ玝�mX����n�ŝ��if���Aee+s-WM�5�+]t���edܫ��
w���b�V'��))�oͪʒfu��ɾk{L53��� �����>+�t\�i3�-���Uk7������Sm>�ʱ�=M��`��r�r�%�.*��Vs}w���]Iˏ)�F�=B��P�*˵ʱ�[��[��r����Y�bո��"n4��WM�����
�z�7;k�CX��v]�6����t{SZ-����nR2TFs���ʣW8�}�A�sz�d�&����R�1��5��t��24��!R�W(�47�2����s��֮�
N�v9���h�
ڀ�ÝD�<�	Qop˾�(垶N/6o3vT���;÷!a�W����=۶� ^H�(��æ�%C�����[�V:��J���z��l�nM����˪��	e����o%�D���ۏU��)���j��I�NY]��>P��m��u�6��� �v���ū"��oؐ�����⎨k3�6�J4.-�qt+w]��;�S�
WPEf.1Jfqv2��K�o�ޑ�Y ^7�N#���X�d�.�ݞ<�}�N	���O���G\�/���I�4��Y�v�:�=�˹�Jp��Mj��y�pMã�����޽�fDP�뾓1���2%c]�n�̧�I�Օ�x��iɳ�-���;j䷒ 2�L��Z�5Ұ��7c�흼}@�uP3�����s|uۿ�#��p�������;����cF��Wl9�$��8P�����k�1)8=X�.uuwWwh���kr��JS������R�E���a2Ī�1Rv<'��PC��	#t�)-�Er4(2L��K<�u��ɜU=8���|~?�3��Q���p�����Ө�ؓ{gsǷ�ޚ�.�R�/V��V�ug�j*e�3称�Ry�vu�=U������]�Ҫ*.q���\�������gy<l�{Xw�]�8i=a\�M���D����X�_m�� �I�1;Ѳoz^�g�I�P���i�	�S�D���J����^Ǔ�{�:BI�U.)*��F	"��Feh��gP�>�=W��	�E�l�'���mm��X��L��J+P�S��R�Z<���U(��L���7�����O+7U��lT�1�b��ؚ!�HzEaml�\���V�3�y)�Z)G�v��ץm�&�[�=��}2�q:����8z7�h�T �KƯ��@EM�7��:�������A\>6\�}!��_Gs�-��y���Xm;��#�˭DHC$ųi/d�d{�zg�ok�����P~F{���_+��-}a/*=�#F48Blz/:�<΅��GWzU}���7uc��y�=�����i�s�A�y�z#�91��m�J0��IѯfWxueu���f��nS��?�fjv*)E�g%ᮋ`Z��������S���RХz��͈�������Q�G��.�n�=�&�L�h��=��7��Bn����;D_v�װ�Xs���^��S����n��R�{hyu�9�e������𺉪��iߝ�=�w�w��[C��~��.���6��z`���v�18�O�G�D��[��c�M'��v
�%��~CU|9#-��+�k��s��+��v�NB�$o�C,!�-5���n��BH��6�����H�J��hFl�f)g��Mҧ��m^���C�IX6�d0��[�Ge�Aq2��Q��V]�K��T� =['P���-gA�}�qn��|����[�h2�Eݱ��"e�Ӥ��uf���ݹ����8p)5��mڬ��z�����v��a-���o{��r�CXz���7mL�V���y��L1�m�1h����T���`���y[_k«���7y9�b{���+Su�lӫ:�ҙ�Y���V߳|9,t���إ�"抯( 0�VL��mR���9^���:؝�P�yi4��j�v������?U�B��+��.�[����S�?�����1Q�r�}����b2݄ӯ��vc����,�w�9q�����0�f>�p�7���6x>��v,ݖ�Cm��i�77%��쭝���]���=#���?!��
}Ci�)k_vSw��|�8�V���3 ���W�/u]��)�����PO�x>���{+�}���	��s��Ɯ�5�L�����y�zxr]9�{��4���׽{T�9��s������7+����ܗ;���^�]lDn>���]�9�Y�i:�9��=���r�V�x'IC�����
;[�D��>�JG2V�R*�U��D���b�!�j�iT~�f�`�CX�9n,������5f
��;%��=���]�|5Y��H��J�Kθ��[_F[�F��ǣt<�MQ19&4^߽��"��S]a�=���>�j�����p���9z��;ҷ{<c���]����Gt�����ֶ��x�~�\�j/w�A~|��>'g/��,EHC��9�ϳ�!����ZT�(Y�|$��G��t���8o�<&����L�F)2�X��Y�p�����xN{&	��&0{%:�K�&}acb�#+��$���#_1�j~��j�}��p��z��¹?�N&y*������}'�9�tM����c�XnF�<����U�����]h
��Su�M�}�ëv�Ȭ�:VV�,�P�1���kw��VA��̕.�^�N����X�m���;���Ï���i�h���Wk����ݣſ�z��+��>�lW�7Gy��0�T�˛��ڋ�]�T��1s3�
̯��M\Hk�hz�J�/�H��]��4!�%q�Y0G�S�E�:��)b�ڕ�-�m�IW���6�H��6u�g{a�}ҭ^�5+.�fԷ6v��:O�,�����bS�u(B�1ͷ���g�>>k}��ϲJf��>��o���ht����K� {T:�-7n��)�v�e�&��	jI��v��t�ٟf屛J�r��>�P�Yt:b���oo���n%�AU�׶n��ofbyv{�\W��4׼�+i������wg�,��8?N,U�Y+M�����ou�z�ߑX�}�kZi=㭪+���[���� :��~JM��*����{���^�MO}o��-����ֲ����K�z��T��*��]���遮A�fu���t�+���J��=��\�Q�<w}j����op�<<�1�`��RG���4y�?������s��:+����	��X3�F�5��9]ⱋÇk���>���Q�ǆ?J�W��;S��atۅ��2:�U� ������"ʦ7����^~ʾ���e�S���b�p���f�xņ<-�����Ⱥ�^������z�f�ŧ2�;��7�Pi���l��g��8xu��7U�Y��N��m9#"O!�;z�899�ܛ�R�ě��0o)�n�t n.�n �a��5���iJtj����[�EW,�.���`���r��v�t�:a��U��7ke^:p�ӯzn/�ڳ�;T��Vxn���L~�&��o�?����9Z��-��Mlt�k.���)��b��'o�.=uQk���p'>�z�S������R�$Â.��=�=���FR���=C*ˡbw?X�~�Сٮ�8���#�j�f��mwI�<��T�:UAz�]������!v>�i�@��.`z�����B�<+��#y+�)rt�6���rGe���1S�[}�q"��)��=ٯ*xz��}�G�[O��q���������=�{"�����Wc������Bu���/����ί���C��>&���t^�����zbϜ��s� ���j�}`uewyΎǳB��1�0uMZLP�HO��G���-���^p�m�ʄ��5.�9r�����=>y�vt�V�ܽw;�~�L�`+����lr�C�P��_�_�7�%G��7�W#�,��r����]Wtz:=��{AO��#��`���L�><V�l��a�9��f�O1γc��Z��s� ��0�Vd��Vf�w��AkM$z�v��vB��=���r�d�ޯ�M)��*��� [S�vl;6u�k5))-�Z��18���ͬ�/��v�\d������=�n4�]L��S�b�~�G�yE��p��0���5��o>N&W�m�X��!s�ʰFzf��V��ך�4H�C��_X�k��Ӌ���rF~Z-~�p�႟���I�Ɯ�w�9b�~���)S��x�n�{|��I���뻄=�{������d�W��OD`s,Z�*s�U~��/Q�l.Ku�~���ٟm����1{-
��y+5�t:����3��u��깪�+�?נ''{Sn�r
��N�[��%_�P~a���6��;����۪�~�.����]ϗa�O�:���v���fE\l(��D^Χ)!WJ�w�ĉo���Ot���$o�P�M��i����-�t�[��ة�&Pw��]}ǲ���2��uބ;n�K�o#����}�^�GkxoF�����Llѷ6�9R+�oi]�����骹�jZ�ӎk�to���	 T�2�]�y6�dY`�v���æ���5a���o��C��a�mM��eo_#�,s]���-2K�g8��#ղ���,�B�r��:Vq'A����W:�3����ʅ[Qv_���=%�i�)kۖ�Fz���-n��t�~�7wv�[��v���<c�,'����j�����o�O��:��>�f�_g�z�}�j۴���]0�G�����.��l��r�d�GO��<yeg�{�}˝��,Sl����WJ�N?t���n�k���y��r/��J�+�ݹ~�k���u���>�Ԯd���=:�j��*
S��!g��r�Նz�j�W�ӱ��Wyʽ1ә�!Z���W��ԃ>�����H�|����n	VS�j
�Է�8�D�ܙ�
�ׅW�0XG��˵}��5�È�w���ɺ��.;B���n �cZFB�h�tc
g��#�l)��{�;�X��qڻIb9[�l-�S����!������:(z��U��βP��Y���m���+sL�HqA��(��Q7.�������nlGf�ꓶ�n��F�IJ7v�RsK��Y��Wvu�hRб�UҤ����;��B��W�\Q��AhcdL�P���c��GggCݷ��Y��Ҁ�N�c�xJC���,V-�����^
���+o�U*��joX�a��-7��c��U������j*g�z(ｚѽ����}9.�խ�>������K��a��ub�E�����t!g���w�_hY#�K��=��+���rE�Z���|�S,��U�z������H��}"��~���,����r嵬U����"9#g8���c���������e�[��ŧ����f�vI�J�Mt�x����*c���zy=�GR��hwgP�0,�{�~��Y��D��睫s�#�!�ڱ��V��ǳ�kZi=㭪3���S����Ng�n�3�~]��l�t)�<�o�{V���So��-����}�mڣT*��wzc2�PV	����k�:���^�����ʽG�̭��E��JB���~�[/�@�C�k���ާ�^�����5�Sы|�
����c_H��_7�[[�K�U؅'h���û1�.�#���]�6h�=�^kl��{[�S.םh���Ř`"�݇�v�}s��f��Aֆ6�&�n]u����SD4��kE�#�g&obt�d�d���
0��t���$�nr8��W?���.�#�F����/H~�tI�m���-�=�{��/|����v@�y�Z-Pbt_�]��x����:��w<����Wj�ѽ�nu&�'_q����l����4# T�˸Yϼ�hr�� T�Ϧ���fZ�y+�b�F�/�Wn���}Q�[�no
:[�<<P�v��!K��ޯ���
�[}}<��l���9���xw���^�\l�E���O�k)�v'ӽ�<�u{��^����/��?:�L��*ŁL<�y������ϣۓ�]U��Ϳ-F�����*n�MS��U|�yC^W�D�B~r�,��^�ޓT�jjf�n�oVy����p��`�!�۰�w`�Oe��ט��ɄWn��}u�n�#�� ):8�C���dwSo��iRZ�,L|8N�f��7�]ׅzxH��O�`eaZ�k��׽w��'��LD����͍��-�� �Pk�8�2w�Ĩʕ��ո;��r�Ept�DР�'K*P����; \U�J��Ӯe
]9�GF^��i�=2���+��9�c��ZG��ea[��մ��z��0x� �[�ýޕ]���n��V��g��D����L��K��cfO���	�H��	��2
�mS���+�w�v=�튭��ͣ3uj҈�nn_y:�e��{~{��Gg_������5������jg��l�����kuM�s��� ��!�7��4#�W8�y&i,�oz����{)O�k�-�BR�7�b:G},@SxOK�x=肣ηV�H��/�[C��l/5�6[���'*��u��C�����AK��:V�,�@�����o �8�PGD���V9"��x��/	���T�˿=Pl����SC�#�i:7�f��!4;��`���x����x����~��exh����2~��'��{=_U�.� �b����YY�O�M�T��Z*�_�BhX갔��1[�B�?���_�DK0#�	 A%���	O���� A �I_��ˇ�I  @< ��pwp(� ��	��!���� � �~;xD{�9� �x��wwwB�� "�w �  � < � �����N �$��D�I@"A$�$�PI(A$� �JI% �$�A  ����Gwwr	��܃�ww ����< 	��܂www �ww ����!���໻�����A  A㻻�{������@�I@ I$�$�PI0� rA$�$�PI(I$���A����������A��0��=�h��N�A �x������^�8�;�(�wp�� ����?��7�}���������.?�����(g���c����c���������H$H$�������?���$H$�A  � A$���� ?D��<?���?A@�A�I���~�_�!���5�G�g��?� pW��������L �'q���� �� �w /q��rq�	�p ��wws�"I$�	% I% B�J$�	$�w<wws��  !�������JDI(�Q �II   � �I����O�����H R  W�q�?_��)��c���!�G��@A'���`7��"I������P�}�	 A'���~���>���D A$~�	 �	?�?h?�@~�����$�	 ��� p@ �	6
����c��G��r���y ��!�s��`@$�O���}��?�@$�L�(�x;����?#�~����� �@~G�� ��$x���	 A'��� >�����)��G�� G������	 A&@�H �� "Oظ:��t������I �	?p0D���qO�7�I �	,������x�? ���
�2��xˍ0�B�����9�>�<���  >�B� (���QJH��
� �
��U(� 
(J�*D@
  � (��@@ �Z��6�
ض�A��jA�Q$�hUQRM�i[bT��(�RT
���E)UU
� ��"��)EU$�_sTH
�>��$�V�E&�֑V�b$��T���!I QUM2"P�����B�H�T!E)*$"�0'�D��!^�   1��+��w\���k[YJ���n���{��u�+�Ά�)֚�A��T��]�ջ*CwT�4��ݐ{=/cA�/�
[��k���"IEW��-�!{�   ���D}�lm�"�P�C}�����#lhP�4'
�lhQ�7�wcZw�^�Of6��Q�$��ۺ+���jٸݙ�k�5l�#+��wX�
؛�C�N���հ5�[sQ�*�V�ٕ_Z��	UEISlH٤�|   n��;ijR.P�*����tv�[(�=R�#Y-�Kc�G�{��

�W��L�t#h�7ai������h=i[��w
Uv�q�ZD �E���$��G�   X�[��ڶpkT�V�9N�*�ө��{{w\�m�w\�i[wm*u�+m���;�[
e�6���jI)B�` * �Ʋ�*i�R��Ǿ  UP����)�Sh�U�@E@�%T�T��7�
(;hR�T+��aTU:.��4A;�([uӪ��U!J�v�R���=�  s�)j�\k�T٭�ԯMv�1�Bv�M�UJ�:6�JST¨��
�J�� (�YMT*�IT*UD��d�/�  �*��� 
�o#�*sQ��m���y�5�<�2(�!�R�`��h
� �cӀ  �JQ	{P�*��;�  =�>��@� ��  F�  {� �0�V��P�r,� �M�( m/q� ���^۳A�iB�6��=�  ���N�P  � P	B  Ж� ��  w�@  8�pP ��� �1�@�S�RJIHGN8l�   1�� 5,��>� n؀  �Z  Ѐ ,ݘ  j0 �w!� V�� ^ �~@e)J� ���JJT ����)���OOP���S�A)J�  �	�R� 0 �)P�U(���W���������������Y��,�԰�2C�ϼ��x�W�w
� D"=�<|���`�1����m����`���ፃo��6m��>���~�O��A� ��E�t2۷�4�R�1�0�c ɸ�i�P���R��A^= m`^(O��|�D����C&�e!��Ɨ�r֛�xJ�W�"�S{X��NT��"e<�0آ@�O.T���֛6P6.��õ��pi��Ո@�ˡV!��I���cܢ��/ႆ�EKR��U�CBOVcmX ��T��;���#W�$�Jj!�w��*b�6�~"Yw�佹�̶���+M<��׆I��!p�J�m�jDw�2mCG-M�tF�[��bUZ���`|of����`���PjOm�JW��㐍�p�oӺiU�Ӏ4�,�]%&��ڗWw���%ǧ2�7OM�n1[�+);���L�?����u��5�E�Iq�u17����B��4%{w�������R�wn�ɗ����-:qy�D�c�BI�O`7Z�aWG-��9�4H6�:�-f��`y��N�Ff*b���t���i�_fƉ�u{�]%*�l`�(��ݽ����Ҧq���u6��Be=�5Rͫ:EA�v�����[T��^h��yvb�����A��:��伀�+u5�K��ؙ�m�3�gI�i4�5|����)l�;Y��.�v6��9!ba�w��r�𬠪��u�.+ei�vec.��D�.���ʘA�un�9C9�Z���ց�d���<[�ն�k��#�nBf�XA�l/)K�5+n���+j�Lځ�����ZÈ�`���[��pd�E12�q2�,eGحQ�)�L�+f�b�m���XmY��(��ÏC�Iƪ^IeK�R��.���%�kv�,���W>j�F&♛O7����t�2��2�2^�SFe�tFY��3XiցLi�j�~Օj�wO���ڴTmܳ-��������Z�Q�{ 4էk3l\Of��Yn��-�����&�K�L8����h�m�Vk:�H��{c3X���p��;�wh�8�m���sS���3]���Y�>m�J&_��v�g�e�*�bq� C2���Y�Æ�&����@H>ēú�%jTP{���;�J%J6��*m�yv6���i	�$��y�\���zV�׵�"T�`��=�c���4�Á��^��a�B��6��-����Z5�Kiku��'f�:��(����4t�\ń�U�B��L7G+8�7Mm��*��W�|�V]KF�z�i�T*]`��ڦ��̚I�	ԖJ���j;@�͎��̶2��WLY%���4��84f��x�<�ŧcuA��4�é4.f$�T�`����fV��*����(��v����9���ڌИӪ�i�%cCd����/���ךm�����N�CUn'g�H����񊲰�L�����Zp�*�e7RL��oAPءkk-��^Y�T.�qXu��5-E�sN�0�n-��H{A�a��Ϛd��ʼ�n鶴&ë�G7m<bͥE�\w��;R�� �Xl[Ś�X��y��o(�b�%d_�Dټ��Nm
b�
�lɘ�,w@WZ©���ʻ�Y��X�m���J����㴄�FW�蕑��i�W^ѐQD�u�a
�.h'N��{$p
!+�sC�N�)�A@�yu���\�%In1k�&�q� �75F
�yY����Lӄn�˨+mYGjP��-��P�E ��F,0Y�
��5�Y�\�p�`�r�Z&]��t.�-؅��6l�HfC5�&����
T���B��e�Z��Eő�s	����
fi���=�Ǻ%+]��8vkl�X3N+��
än�9�f3 ������f������Ӿ͡���{�˻m�3��n�Q4#s&��$էu�l���Xr��6�k[�7.ҬlcX1D�t]k�c ��fMb��4�% �A�[M��[+-�:�(.X����S�=������ą�^������I�v*��YM}4�kk2�ݼѫr�zl�	@sm8kUI��Pf���Cfh�N�=t�ތ�j�4�Ni1��lF�e�B�N��mIv���(Dud!,�r1�P�����4$a���P�i�\7���?���j��C�
*����8��z��3��A���އ��b���7VhEC��t�(^���u$�4, .4偔E�u�6qE��^��0�ӻX��$���z�i�X�V*�o61�����;�2�$嗝�n�����G�(ϲDځ]l⣗��sXN�EU��G[6K�P����)��c�Pc6�K��Vn�ɠ[�zi�x�b�� #�}x�v�~��j�`h��>�-S�PϏ�З5�ɴ�j:2�,XZ)�F�?�`�
�L�n���,^:a ��Z��2ݍݢ��w��	�a�g3����t�����a�V�d�6P��F�]!�#�͐�餎�0&�뻎�_�bm ,���ǖ\�3e�&un�m^�=s$��c3J��`y��!]f4���(^b%�_��vݒ�j]�����K�����ȩV3S�o4:j���u�����A��A�w������/C1����֯vY�>'T�:M��(j��h�V	�i��|5�H'�B���c�z��I���R�z)27�2�6�LX�p��8�5q�:�^ieX��7(�T�*$6�p���(ޙJ�cv�	�5J@eZ��ܳ*D�p�z�ݣ�����#!A<rҧ)�E��Ŷ�"�uc3-�kKi�ռ���E��*Monے�j�z��;R�j�VS��(+ #�OS�n�2԰t��J�dS�E:[UkJ�7mܼj��0����K��+���n��SJ���I5�a8M���V�-SH��NX
\Md����j�4�9!�%e������i�5zi�y �b�=])��.��plV�:Z6��{��4"F���EG�!-��[*4����@875�Cj6���т�Ň(\��V���wi�uy�9��Y�n���=G-��+�2�]�u��n4rѼչ��f�ѦT��� ���R��3z�E�YA���w���)[�.��5��K��ě�&7XV�CN�2�14��,�)��[M�9N7�N��t�[�tS�*�u����[�[�jWWa�e,�J���i�Z{Y����mbb|��nY�J���ï4��*U�Ϊ��ѭ�h,�R��M�j茣m�V�(˽/FK�v�ӻL��9A��B��u�V�7,�,[�(9�En[�I��f&�^jɗjkA��wkӦ�7cT:�ŵ
ׂ�&�� b��Sõ!3q�E�����l���tMц�vF#K�ڔ�5�=�gU�Ѹ�X�,�K���&��T^�!�W&d�ZU]C38*v��uu�QZ�`�d;��z�����ay
jlZ&n#�m�)�-�j��MgXE�Z�u�2�r��-�p�WJ	 ]e���2�e�ڗT��dm~�C+v�n^�.�H���Ztwt�w�c��i�x����;ˡW��Nf޴M[Gn�&�-:?�&��!��*y�/^���oL�;6 @�E��;���Z��׽�nƩ]7"�Z�x��#K;�x+f�"��7X��7n��y�6�Ul���mGN������V�pV�����voM�ӗ��VV�!�s���@��t�`�� ��n��K���B�U�0Fk-�t�U��0Ő;�9�v�ә
J��3j��;aL�N�t��kn6($�ٰnˤm˼�0�TY{�&��Bݼi��	����
��raF����:��ksH!`�Å�"];Ax*Z2�l.8E�P�K�� $��"���*�������n��>
���z#n��˰���3�>�rnl����vn�=��i���P�6o W$J�U֝�`���Y��n�)^�Ъ�)�X�WGs�N�v<Y�����2T+b��9B#�?�d�&f����7AO�e�0��[���2�-Xv�y6�ƨ��"����f�K\	��p�G�*���P}�5��δ�d53��B��[j��,�����1�%k(}b�+��Dm��E�H���B�@�"R9d������ٹ�)����+nL�ٚ3p���o	�{L0�=�Ք�YԖ5N����
����/��曥�ܩHO��G ��
�qӦ�Q�ChܺF4N�� ��@֨(7PBP�yM���g�ܥ��y��C�X/	�Wtҕ�zl7��)�X[����c4�I�r�!��RF�ʛ�u����+�q�B�҉l���m�h��@3u崵���ja2��V�y)�s��3~I��mV��H5�Mc��N^+�*a�%4�`�R͖��3&E1C�j�Z5���0̫@�>��P��0b[���Z"�t�Pv@�Ij��XN�mc���Ҏ�W�(\�SiV�^�i�J��`)����{Sr��cp�� �T��Ū;�ZӑV� \1,.�*: k�gk^����6��y4��NU��7�j��+��� ,�Е&�6l�F�sHK]��-�W��$z�V��<�2 �n�uի���� �iͬ"�II=J�X8�"�����3z7]@ɲ���2�4:�Բ�%}ɧ���ɂ؈[q�7��ϞHwr��Ci�oi8wu��*��$.�U��M84���Jק0�HT7n͍�z-L�kM��$j��c�5Z4����6�R�MZ�.��h��٥z���*��!�*�5{�ʶkd2����@j��yM-��4�R��7)��������� A9��m�̓]c����ǋK]`�Ar����B/s.�gRz�:������q��i���5�,��x	�&�6�e^(�k�����E��{a#���20��V��n[YMD̳Df�V^^�_4k��9tkYƵ=n��%m��/�RZ��	��+e��+^m��T��u
��b�3_�7l�ŗy��8k)��XRM�,Ƙ�&R��D��mM��`�BdB
�]��{W�-EY��9�ħ�$Qn���"�b%Q��]���Ֆ��҃z���J[i�؆��(�{�]̺Uki*=X��%0�"R�ecf�o�r��E"�P�!u�Iטl�5�*b���!��R�!O�PB���,y��x~lb���������b��r�%�42]�t�6�Er(���<{�սd=�8��u�_�n�f|�5E� F︧�����Eѭa6{�ki�a�]�u�A\Y`d�(@~�D�fT�iT��ܼX�Px3X'��MYy,$ٵ��,���F8���]�M��tf+�f��P�b�ђ�vŚ�  ���n��Ywwx��*md��n�yR²���^�"�K���?������圚����S�B��.Z/5��oJZ�u"�����-�?Hm)7s��n�`�a(���Q�%@h\s6U�@[��)��0Q�F�H��� */����鵡Pv��n^��nR���ț	�KI.9[d�Ѥv�����9Wd��M?�UŐĶ�$�j"������{�S"B��Q�&I�~��1K�;�D�3I"�$ǆP���m�u,���;(�Y�o%M��obҮkQ���-��W(�@H0J��DXr����de��R�2�*L���l��}1U�`��/B�Z��w�'e@��0��^�r�X��f��蝚�ͬ�YPP{c*K�l��fЅ*܍�)ۺܼi5��Bӓ�h�ژ�cdXc�5��n������Ø���Ma�h;���鶍a�v4
u�P}vr�0^.�O(Pv��^�x �X�a6�+@����a^P�deҀT��w^��*�Ѽb��6�2�[ӕ��ց�:u&��;O��s��*�n�m.���s�(���܂�I٘�в��V�ڙ@'O0X4�z������I��l0造q�y-��#X��� ѻ)�74�a[D�VAu�LR���r�ͱ�/,b�jL���+�K.���6�\�8����F*nе&���F(m]���
���CJj-A����̀\���~e֗/%��	3 ݷh�"�b�T/�,�������<��S�6�+�x�/P���.�Y���q�x�`	xI-dmdZ���6��7H���3@WJ�b���ڔ�F#�7�3a��L���Q��j�s&��9�κ�1� ��r�)R�M�X&�ww_i�r�4	=�@mf�*VwD��u{qT����'�8��q*��L
!էic6*hԌg	y��Qm�f��j���U�p�f����dLן<����$��m`�5���6��F`��4�ʺ�kU<���cm��魇X�<��ۺ�KhR(heՃȆ�l<�����66�hʺ���Jn6��a����Q�&�r�1�ք*��,hM�Ơ�"���[6���PB���=)<'p�%,u�ga��XY�6Y��H��c��zPè3�;�FZ"��o#ó�򮥙KI�e���B�^�1��J
��*���0�Q�9y���M­��f�x"'U���[D�^n�RR�h����>�8����z&^�*����aw��=GU�H֥��%6V���r�2�R��zܹ�J�m%M�Mj{�h�f�� ��G-4v�b!q��Oa�掚T��b�{LQ˭Ps%�ѕ�b�f�D�V�*[�ңa��ih�M��4.�j��[U� )��0���vl�4D�5m� ^-�6���9h��B�Q�.<;G'�:�G3�e��t��Z�:��zjnT��0<��/�%Go\���jG�R�V�95���T肭� .��i����"�Ǫ�� �@���1�T�!^̖ Hf�����n��X�S3]�DX�7k�b�J�6a����m��o�Z���� �e7�&�kww��n�;�%0����L��OM@�ė�H��-� s�CV��x�tS8 ���ٶ���"����#]���U��='�Թt�d�J�ón�}n�T	��u)̭t�`�H��b�o��U��������5�U5Z�֍�*�ݼͲ+u��.b`�!ݽ1kݏ0�;dW^�]��c�o.5E�Dv̊o+��ޛ�����Q!�U�c@bX�-V�e[KB X@ ��؝A��ԏ*|�s�ma������z�'4��]����F0v�1TQ:݅p�)=���V��}m�+hd!Rѽ��(&kBbF�Z3��Znn���ڋ���oegp?��6��뱠�c��Z��x����fT<��q�N̙�5�8�e{�37��\ݽ^-v�E4�z.���@��{��hq�u[���t3y���ެ@P�]�����׫[��C�kd(VK�GNd{%3w��gu�Yc❛ųGPT�q��ν������\
[�
�W%'0�.�CDx��ڜ��m:ډT�X�Gp��Y�9��&�js���ç�A�^�U�=m�C:3��<�A����d�ޚ��s����/3=[�t<�5�G.��2����Lt���9Մ�j�Y��l3�am8p��.٧/6�ژ�蕡{�ojR��E��oi��:�o:�ц�7��]�o1ӓB���uv����1�v�+�a�\M�b���`�b	���n�Z���u����E|7f�JS�a|	�6������gv�� պ��v���d(J1����U�df���qkr�m��8S��.�4�v��Ƒ92�5�y�]s�A�P��Q9��fV�%�Uu՚�v:EH�0	����D�a��Nr��e�����-�(��S�ݲ�&_x!�k��¬'��^W�;ͨᕚ�7�ն�+&�V����`�d��H�/E)يJЅV�K�jQ�|�A7]���@���L7CF�é;CY8��Ho�g��C(L*���(h�kǝ��=��,݄�a���0 ��V9�����z�hj��!����d��b �W�ʤ�,_l��]<n�Q�%V�����ۜ����j �:��9yt����e�xo�+��VIaQ����S��0G�����l�m��ò�F.׹w��h�؍���KZ�2�X�6m�cC�D�E
��
RYż.��;���5��F�)L	㛨)�������p
��6��=���_�Ǳ=�=[eR�f���n�V�'!�*+�/5�ݾt{j\��޻�k��8J�4�E$��j�(_ms|p2U,į5��{l�:���1��5��{2�!��:���<#��n�rI��@�o]���,�N��dٶ�)N\�-�W�D����W��NBId�S���n��1�\��ng+X%�f4]b4�R��'�9Z�оh��KY��6�h=�u��2���$	��i׻�U';��/3宑����\�c�.�onH�휨c�� 6e�*|�e>���ST��0u[�X'<hݽQ;P�&�R��͌7�.�K ٯpa�ƺ{H.b�6'%����X���Sͭ�K_M�+��h^��Z�wZ�J�@+Ecΐ�hW�O�s2lM�S݉�ܒ���i�����r��*+�&A�N�v��$ֶ{��`��S����Ş	�L�cP�
-;��أ�Ŕ���V�ioV��0�a�ݮ�D�������p�������v��N���x�˵w"bQ@��J �Y�zCa��ߗ:\��rNo*KT%��:�V�j��i*Y%�m�s�Ǫcth�w�F���ݍu�����}�܍"��ɒ��{j�W�Q�Y��+_u�8��֭Qo;H�����L�G:C��?�4݄��.��)٣kxk[;�Ǉ��H.�zZ����%˪ �^Ku�sa)SCr쳽��	������yr����hk�r5�xΥXȬh-�M������j���=�vSQQG/��A���m��7��.ޗM�w��У���Z�+�Ẽ�]�A�ڵE�vN�/>{�/g:q�ΐ�ݷ|L�:��ط�*5l� �E�T����Ba�})�ҝw��l�N�FSDӆw�8v���(!�Цr�_G���j�BL��4�Ľ#���m�K�w�=�ks:D,`���n�4�����������BeR7#Mj�^)��m�>�Hرn,��(�T��!Ko�q�͔�7z�ΘVZ�J�[�B�4"Le�PV�٪�cmEp�9R`*�a�Pܬr���K%g�)W*�M>{3j�Ѧ�܎�p��!�A�d�C��i����e`f�����������E�
n�����')��F��?N�q;R�3�z8uYz��n�(�PW�v:˭��|f�i)y��b8b�c��U��|���9"g;E<]�B`f˝���6��mu�Gz�62j�x����\1M�]�U]��l�:Ġ�_hS�*�)��Nyɽ���]��)ݲ���쫸�^�aٰ�˘�eN�
۩�Ҵ�����ھKhN���Ұn��v�<�J�+�Pr.�]+��%Ip�c�9D���6Ĩ�Г3C�4UMyF��2^��_q�ex��R��U��{;����]v�+��w�F.p����F��c9�:�g^y+��J6+7X�7�o.�wO�]�+�0l�.�d�*\KP��k4�ˮ�Y��ܼ�m�\	i�:I}4e�,V�F��f��[��%���+(��8�,�'9�9bǨ.�t���6TJ�����XH��%�Z�ܕ�
�M���O���]+F)B>!^�[o�G�]�sOX�VӮ%S>�3I[��&3&���}'�k)���ʄZ�༕��S1e�K�Ҧv�V�S'F�)}u'S#N�x�EV�d]p�s6�8�Mv��P��ee3�)�i27�;H���Ę�1��X�fl%E�����,���_�Ƞ���c�ˮ��V�]6:�TS�;{�`�|�x*L���Ԭ�(�xǽ�4��
����pLk;`+��`i��֛�c:�(9�$g�s=��U��@c2����m�[N�U��3Q��F�f�r�x�:�X2`�gmpܴ�� �9�V/��Q�hT�bTZ	�ˏW|pt��b�IK/�"�^����m�rY^�XL��u^�e:-��,՜�{�B	)�u"��������:�]径���+g"s�ە���aU6�uc��@5�GTtj�6mg�n�^
�Z�m-���^�T�u�bV���+E0�@��)^V����BH����vWL���N���`�keYU�����)J�c��S.�ֽ�]������Ѯ�˕�C�U�B>4��s,]c��Km&
�v�n���	A �gd2�e�.�V���s���G�a"A	�b�����u��Q��;��m� ȩ3YÄ�"]s�h%T��^A]0��ժrw����h�e�Q�B.9�fFII�9��c��-%Yj�ւv5a�[�BR�{ݶ����
���s ��eH��[��ig��8�8^���#��$��_,\{��6"�XY��.�.<���C�I��-�J�����l���6B�����5�����c^^l�XSrw)��=�j��*��wN:�������)s�+�mlR�-��2z7s)_^���t�s��Gy����y'f��WO�䙛T�v��Ӻ�-���+noC.���`욟|�!`y���+@��齘O`�vh�,|�:3fJ@c��K0��qP��y�3�D�4��[%�mm�.-ý[ǆ�+B����SM�� �m�Tc���0�.�*�9(R�pd%��S}bq���"�g(��p�j���6�h5�R�4�>8Fb�k�kק�)t�bU��:�{;��6��6N\bJ����|�m�ێ5 �;K�t�k%t��k��]��-:.��n���t�o8-�"�$Ni�6����
bh��;���0n��t�ֲ!����Vs�q����B�;�2�R��\��+��c7I���ܽN�Emh,��"���`�e����{_<}޴ױ����]oP��Z�N��L��n�nLX�=��q|Q�`�w����R�f���;i�+������E�^�s�/�C�"�P��Tҩ�1�w��%�G.�������j�\��fj������P���M�f����퉇��bHԮIōg$/Ew.���"ޥm,o`��;���(ou'�ӰB�ٕu�n��[
�}ʃq������R��I��Cۼr�Ym=4RxU>�W`��Ox��Y��A�/te����5��bo 툱��i��a�Z,l �=�gq$p�kOcj���|�ǳn�����������Ld.�
f���!Z��	�����!�6���F�W��t1u��@�9wE��z�E���� �vC�N��ĦK�$�;t�WV\;5���;��|/J��J��8ث*�;������(gd.��l��D�|1����.ƮH���7�p����A�f�b[C�M9.V+̈�z��IJ9�P!���K���Pݾi2�#O8��I���2�t��{,�DƳF��
�;c�ܮ�X:��H�}1�sy����i���c�3m�:���Z��vn3Aس��w�6��������u���A���U�ޮЅ�������3���E5�_L�p�;�a$,��F��^އ���-{t����J��C��|��+�5q����n�3�����1�<�{52��3�|��G<�Am�\���S��#>	�r�n%�����5'X{I�0�n��u���a��l'4��R�*q��Ⱦ�R�G�v�-�f�r�n:Zm򸣼�t���  ��)M�w;~b��P�:���M�c�:e
2��e��{r��S�n�D^�_1�.��9�Q��{E.�[��Y/�V뢸�ϧ�1�0e�skN��?��Сԑ�.w`�zq@���n�>M<ÁvB��ZgXxq�^u*��0��meX��IyÅ��&	勢�v�� J��Xv_;��v�'p���G")�ϞA�gWXeJ{�;��M��Xj	�H�}1P�B�MM�sVwf�=ӛN��k ��F�j��c��I��؇{���i�m�V��0;ݱ�J��ɩ�Tȑ]��{2�"�: {P�VNS����c^c�֖\��Ȯ��\Hk��;M\�,�畹����V޷WXJ�Dk��Х��4��:���!���X��Il��m��V6ȫI��GqvH9_�c����QW�P�C�W�x�:I��wv�833:9.��DR���U`���ԏw`�-�5��oPEf��'���)n�mYgn�n�p�'_o*�5��]}�E�1ʩ<rɰ��/h�u�#�ͽ�Vv0�XNv<ZTS�xn�iR�:���ѣK�8�.�G�X��l�.:��f�6���Ue�� ���U�T����E��WV�#����W+���S{�2K&1b#[�X{˰��>���eQ�S��k.�Y�x�p�!��`Ufm��c�~ı|�fPƺ�-��ڮC�@�1�K�i��}J5@,�嚓�x��FٚNJz�/o��X].]�3&d1�(\��•�����}�^�ޤ����ClWaP����������J��&�y�s2��/��+5�Be�	%1��u�f!HX[��37([�Q}͒o��:��e0�B���t�0����$vN	�aN,lbz8��
�Ր�����u��{�Ayz�#�3�iL����6�hIׯ���{dfNd�A�g��{�CL7��\g�K���g(ӡ͙ZzcZ,�����娏a^���U؋+/g�U�͸F�zv��g,�@Z�4� ���^|v7(ѭI�r�p�Z��t��Cb1QIa�ʷV�\#��O3t��"��N[`�h���{	AV��vЩmV:����-��\P�r�gS�d��Ѯ���0̦���؞���m�۬��{o���}�m!����aR��#����8��a�彐7z0���WM�8����kM%�����O���f�w;EJH7�^�uY��C��o������Cp��qSD�<f��hR4�7V�K$���:���O�!k��he��۫�9�}ѫ�3�0�U��+�\��M��7߃�ܤx=�3t�z�<�����GӾ��}f���|�1����3���YG�dz6�!�(.�D��z��yt�==�Y}�D$�;
uy�y[��×��*��{8l��k5�syV��+�M*Cy�Z�r!yoOsv������+�k�c�Ԧ��x���4���>7�k6���s2��C*�5�J2���w����X�ŵ��K���t����1u�0�9�woW$��ێ�6N�v!���Uz�";:�2(��Ren=����s�!�ⶍ�%Îf��������:�F�6�����%�Z�^�L.������R��E�٣��z"�:�����'�P�s��d�M�gk*4��os!��ڈ�����ս�0z[7|�`&^,de��24lv�7F9E�;�N��.Wη�S�t]0�z���+Ҷ�g!�������M�.�m�I�y�KL��z�P��:����X*������f��$��Ō�,��B�hO��ٻ;*�b%I�cC�K���8�v-�i�x�9p��-s�!)뮰�қY�λ�ܲ��!�1�Ҕ�W;Gn��E �^�����T�a�Im�,����23kyM�A�z��!i�˼�t ,	���CN8r>z���m��(�t��M�nN�cX�\�a�HAe�ne�ᵨ�����^�65;�� �ݟ(X�	F��ȍEB:]9�6ܫ)D��{Ⱦ�
��ӠzמS�H�����J:��)tC��l�yNy�(d��`�cc������o_=���w��&~��:ׄU��Hm�nX��F�'���ac)��� .EA�����
C!(r�>�媜����Ƕg=ǆU:�xjc���]ڭZ�� ݭ�Y�ɣN�5���yV�JԹ��U|�[XPD=�5����ʭۨxÓ�{�(�w�6�*%���U��ZA3s��a�>�:�o�����WA�wM�G8j��Sn� �4�P��[s�X������5���J_�2�,4H��ԅ�n� JU��@=�[2��N��NQ���ӕ��.޲�|g"�kvf�k�r�ղ��&��zβk�/��Yu�Ix�p��e�]O/i�"لN�sis�A�I۬qR;�.^��)������k��85���U��z�\2UqA):����osJ{��G��V˭4W�CrWt�-�����a���*�,��Fe��F$T��j���5o Y��|I�]ٜ��4eⱴ)vN/9Q�� �=d3��\��,u�2����IAl���EZ��b���G} Yk��-}�=�nJ�����Me;�*���D��й��l)����1#-��Vb�N��=E@�Qu�0���w��n��:^�����r�jQ"���ͮM=�7ᙨ����1�v�ȍ�H	�u�uh�cfb{i�)Tn�Y�gu۴E�'	���[3�<2��s��j���iL4#����9�����>B|��hd�xM�u"K:SB+j����5���'LU̍�q�z~z�=I؋P?vŮT�v@�u��څ�7W��V�S+�h`Gzj�TF�䶅�f�J�͹SY�����T6���/]�-����v2ܬ�{)�Z�C�L]���<�ф $���4v��L�.[�^u�E����`n�.9W��t2�]NS�ԧ
,tj����{��t�����ѧ6����j5��!�r!j2��\�&E�fn3�L�+�gD�W��NaM\�2�ѫW��I�Z��kJA��"�i�N�6��u3�
Κ� J˜�M�9˾�r�3-���h^�����<0�{i}u�WSN��-�P�{��'�{��C���2�ڱ�c���\��TKHpuDhǼ�0�C�<R�wO'r�j�}CNZl�^Mr�v��t��iTNۺ6i��Q���-9�ol��M�l���9ipC)>�v^���s�hFY��pi����5 �|q��d�3�T�y�J�/v|�VҶ����[˫��}N�ER�򗘛�ME�;o8_�:i�n�6�T�y�zS��=/.����� �Y=XZ�u���,�@U�.��7�g���mͮp�h㔩ٙ��׆�Fa�)��;��X�.���l(��+.P���͘�>�q�Mj?<
7jw��+\u�X�q5�
�;��Z'r��3�`�]u4�]�hO��kS[��6�	��v��l�ky 7GQ�t>ݰ�n	��q����[��{.�}1�^��RθXf�<�i֩�$�-|^R�#��V�K�ۃ3N_�.]��Jª�on*oϸ(\��	*�=�Pe����'R����\�kêp�Dd���{����sn�o-YR��6,7XϞ�{u�\��YL᭣7bcǅ�Ō���/Sw��%��oJm�IP���0i݊�f�Ɏ�c6U4&鼱{��#ɭ%�s��D��l�̦e-1��o���J��@b�/z��I�|qǒ���������h<�����\���m�5ò����4�����������Ԯi�Y庌�g2���j�lї��Gp�b��SӘ��F�wv[{P���]��\��X�շh��;��Z����u���h�}�c߄㚸NuLN��xm�Ȍ	!`j�qލ�����4
��{'o>��^D�wm��Ew���=�kb�"���^�~��m����xmVeW���r�vSdo>��t7��>�\�c� "�<�c�`��s���d�!��K\H6�F�t/Za�v��m4�!�Zz'��dP橪Y�w���3�p+�R�eа�a�V���%ehSr��Z�{�tt�r�T]����;vG�Z��L��O+c�z�wRt��՛�i�+n�(M^����+2]�,�M���c�@���^ʍO���,[+���l�p:֛�uڭ�Dxst��`�L|0Ծw���E��w�S�l:���KV��+ub[��T�]V�n�&��`��\���+n������l�����O�Kn��YC&�����l�gW{]��Kq#�k%gb�w�%Ƣ\h�.򁻻]�`�GR%�U���.�<�����;�\��ݗ�4#1���f�|fv,�5����m��E���0�5�AR��)��[�GG���Z����gZc�
�z��9^�dM�GV�����������Tk�v�Evc{�k��Qs��g]���>;�;H}v®��c%���eM��pM������gr���uae����t9�S���?�޻ci��L���mR����@mkV�u���Z�����׫kWIs_�>����� ��!�5s�r�ޡ���2��w�ھ��蝓#��᭄�H�Ε-M�<�����oO �Vn�X7���Ҏ�[Q)(�����1���#|K{(�*��f�AW/Iyu67�w�������l�n�0�y���̺I�E��.:r|���(���nV �D\Ws�^��f��+�+�%��įk��Qnˡv�ZT��7��
fE6�Z���sÝ��m]���erZ���M0t�!�s�\��T㑚�%X��_M9���{8ֹ�p��XT��\��]�;�qna6�  f��� s?;���X��%]y��ܭQ-��]Vi�#����Gw� �Ohm���1)j��Z�{o_IV��LscK-0�W���Ի�i�,i��ޣ�6��qF���X�����S��R��54�n�^���Ji�`26*S��M��w��RS[�C��8�N�]f�ɴ��(w���jS��g�Q�j�i�R��]ڬFn��#��ѐ��L��>�-��rn����(����yJk�ډy;��B�犕=b�
�Af�{�ݮ����c���������$�[B��N�<z�\*�"��C�0Q��Ս�3��9c���,`�k�V�	xN\9�����i�.��[�Ms@.=fm#�z�eLU�ir��5�@�*û��\���<��*U�gB�֮k��,��{���1	M�-_Z����e�i�C�WK��''<il����q���4ھ�a2�h"��{\��쭡N'x4�'pF��b�4NH�v:�l�;�Z�=a�X��WR��.��R��KA���}�U����6���7yc�dK���E��:�å4rN+rb�i+Ոfa�n*ׁa���f�w�U)��ܴ^��Dmv����b[���݋�X7��OQ�д��.@�R���t���AZhn�A�B:�B���\��r���X���8f�f�)���W@�8 .[�,ÛX:�\Ɩpg	g��a���/P��m�z�Ӧe�]j�'Y��)ݐ����&m���ں��:�έ
1�*y��7�s��ћN�v5���wa޺F�.#6ލ����vM��R['sW|�VP���F��l�)񡻕�u*���I�DmE�!1r�g�\�Nq�:�f��G��f�k)��ذ���`�Ε�����f_X3mV��$�l<�4�M����e�a��hmA�6�Z۔��a��IDs�i��Vf�ö��yդs�]��+pe��CC��Mw0W;�)L��o��_e�vh:���U�!d�K9f#M���Z+Q�+y�Yts����V�6f���.����ѫf3�4����3�M�ln]̋hK�l�]s�{&d	�uӢ�*4Eh!�N�m+泹|�T�6>�/v��	��7�I�����c�؎��L�Ի�J2�(P�C|^wр�A �ת����MU���2u�{�^���3�em"/�C*��I�E������!o9��M�`}a1h�Y}�K�z"�S����tr�*SH���R�x�q����6K���a�85e��1�+���Cn��8�MB�]�*�J9R5�h�vQcR{�I�yF+ɚ�����Wغ]�v]CW�n��*�OS[z���
�L˔�(-��L��ΊGV��ؔ�>�	�wWageu:�nCZL䯭��tqx%�i��G;(����7��L`�zom�'���{�v�7�+��:ھ��j��uV�nrgo���5]ʙ����-��|��8�\��S �'���]0r3��&�NF���h2hg:<4C�2�i����;Gby���-�Wi���f�Qh7�6Q �[Z	w&lfo.7��< J��ů��D@��|��Ռ��Q �+I�jWr�ά�Ӕ;b����v=oq�v�.Kp�b��ՊyMѣ2�KOi=�5�UP+�H�q
�ž�KM����鷥���A�ä��A��c�3sl&�;7���:l��C�T0˂ͫ��%�B[�T�T�9�)k��{x��a�^��B�ͧ�'s2����1��cV�ڥ�7f��|[�a�
��+%n3��#�c�٘�p*��/��Ou4I8�:}G��kEio>�Ŗ
��1�`��Y���Z�,'[V���_S���Љ��{�m����[�j�j�m�5W�����.d�W}q�"���↕�J���O�j�q��ow�B�d��`��la�Ρ��Ŧ����LMRu�d��q��1:��N�����-U�=�ɸ�X�ᦰ`��ζ��FM�DD��:�*Yͨq�8�R��Uݑ�eI9n���g>��n��B�wjO��A,b��\�����ǘ2T�����X�V��i��J3�+$7h�*��e_zX�}��*����Oo��*�R�6v�Ky9���q��Xe@1��A�ݡrP����a<\��a-I��{2V���.�7N�.� �Ƞ`U[\ti��;��Tu�
���)]���H�o
	E�9��rV��f�����1�'��VJӔ��0)�h�x�\1O��nh��<!:)���5K����Eq�o[��>��'[o��\J̲��*M�W�G��/�K��x6]]���6� �v\���iCX�|�����2��;~Ε��<�u�&tɁ�иvKc���o#�i���T��b�ˁ��Q�e�۲�R�ٱ��(30Ag��ۻ=��Ŋ<L��B�bu��iR�* M*]�M&�FÕa"+J5#[	B�N��.Jꐭ�KN��>��yga��t@IX����{�K0����ls
�k��k���H'��kb.���,T��qff�s�ۅh�K�����o �� 0��1��ONCIfS����;+�*�5��������x�+ܩ(o7����v^��y�Ή����'x��eḊ:�4a�v�DW.k2�[�5� ��gc�3���bc�g�ܺ�L���ih�d��Q4�K�m��_|/�S1��9�8�b�l�^�kE���	�{�Y5�)�K*4�$	�7v�"�K$R�)h�E	B�D�^����:ћ���X�ݳB�cQ�� �K��-[1m(Z�=[�u*�}a��ɝ� }]�*l�7deD��z:�����	�hP뽑&�x"�����b�ttD�S�v����o�Y�����g�K�`Le�"D�۴���]������M�E��z�Ń�OJ}{�ݤ�[�̤����a�ݡ�ۙz.^�9��ܧz�	���5�q�\��O�:�M�<r�V�[��d�[�e���X�2�`��&��n
]t���̛\81ǧx�S;�{F�q��{��y,X:�d]P;3.YH�2� �o�c|tl����/Q�a.#mm��֚�{� ��mr�0�s&��q�V[s�*��43�	Ʊ�G\�]�3��j5֙@��v��ҽ�������jU�j�����sP���[h>�\^��]Gg���V���˜�ҶG�p[��3A%y��Y�r����bta��)�W�OU[
���kuYWcY"�>���2��9e޴Nݨ6�1�J+N��F��=����F01�ru
���8'v��'ApH���;�T��lm�/V��DY3�@>f���֑{R4��o�V�}ڏn�V(��F�{�7gm3u�\��B���R��-�s(�r��t��P���>kј�T�����cZ��&﶐9�MP����5mENɕ2���4�Vӣ\�Vq<�.Rѻ�F� )�Sz�����ͳ�{y��eNg9�ֲ�u�� !k�m0WwaҼ��i��u���nPu��ĭ]��gE�*�5^X֎��@�u�w�G;)g�laX��W����a��&a�:4V��-�y[n�e���>q���� ���h٦�nU��WE=yʗa��Ŋp�-d�6��]A��sǼʉ*س0��0�Y� �]Zvh.�y���ƻ��f�h�:j��݄h�i��^͔��Gln0C���yD�5f,���������q�5�eabPGuD;�r����(ia$@�uǪ����`.�w��V{"s�5����^U���Kz��*��OA�p�/ApT�dkE.Z�h۬6�'��d�֌��w�64A�Gڗs����%Uz����Z)���s��oY���d5z�w.X�T]���}z���94��ʝOƺ�۰����<��̍w�|�&ө��p[O�.�i-���v�ޑpd�#��71e(����-�+�;u�Uʲ�{�NC�c��Q&�s��S*�r�t����k8IpFT󃭾3/Rڲ���ז
�I�'���2��W9ٹ��F:��1��Uu
���G���왂�mhG8�'�ѽy ��g1J�g:ͼwd=�M��ޮ�o�U}�W�����^���sDP�6�����Ԙ�����J�Kȴ�X�,����'��o)�;jgPR^7�&�x�����iY�Uޠ�&�x!n�w+Ua;	
��|u_:OU��'���IK�n���G}����{�+#�(���89�������Ż#�9@e��.��d� -��
R��j�o!���������"����lK�lD���[�I�ڄ�Iqk��pvRk�z
x�E�i�*��qyqp͕5�r.p�|�*�i���dړ�ncz�'1�������I�Y=/�h�C8E ��+��Ź�R�Q��e,N#&=�b ���כw��y�s2���/n����VX�,T��e���9
�J�l�6Ô��v	�����LL:ic�q��{�	C!�])Y�4�M�έ�7����/,/�e	�U��a8�Z���]r�K{)wBf��۠���<;zVG�c}�f:!.*�bʕ��Is��a�H���n ���u�<x&��F�i"��Bj���1)-�q)��P�@��F�S�>�:��w�c`Q��M�{��S6����ܺ������{�jn��!s�ҕ�/(�ݵ�>J<,�#Wm+��|3{��[��S�ӷ,D*�"�R�Cյ�M��`*�y��\�=�iL���4�A3 �t�h�;�|�A�r.��3\�D�+�8�r��/�QW��n_��:	D�( B��@� S���J���
�P���O]u�$�$S0�p��1c���KD�
��[�9n�wH�"I%1�r�rw���3SYah\�3�� �TcU�QZ	�^�9D�*��E��B����\,�OP��*�''"�.��g�c�x��dRI±���r��Ewt�$�NY'N
�v�A,wr=LL�(5�l�S�RBL�Ee�EȊ4# 3��YAXdfEZJ����FU�Q��*�eX�eӖ�Du��*�
%���BDB�u,+�4�H駞:ң���ڴ��*�/\��
�BgJ8f8��Dhfp�C$�-fl��=C�]�ٜL��mB��*	���j�s�\(�Tt� ��34�RQ��C���PM(�UQ5!B�K����BIE�L30�ZE�!!K.Z��'Q):fLN�;?���^=��0��N��ܽ�uA�':�ǖfaV�$����G�*�;�.
��y/���[δ�o����1���E����s�Uo�Ʈ��r�]�{���K�M�G��˨���#ŰeKb��G~"��;��f�[nCa�i�;C�!cu�鷫���8ՅqAX.��P'zv�k9�."�쯵:˛�搘zҸk�x*1p�T-}���c��M�į�8u�����q`'#������{�'ro4,�T&LeA�����r���;1��3��SؾX~	���r��k!����u6Χ�i?���|{VK�� F���)�c��e
�YW�*���ߖ;�ddE$��p�=����7
�B�.�aU�/WJY�Xݫ������?X�����5&�mP	gÝ���7$R���S�����v�n�s���(�U��Ib�+Z���,C�y�$���A�ޮX�쮵�.\GxL.T���c��)�(WS�;�.p�A^HLL���Y3�����!��[0Y��rc#y���ں�-�\ő�[ݾ�Ԗ_1�o�Q[ �Z�hD�&N��|�s�%�`H{���:�\�@�wY��r���LpH�Qy�>�ҙtx֧wr�ͫ�)	%w!�K&um��n��eK��^Q/x��e�C4�e����G��fG��������pI�Ά������HD�|9j�s��[ٮ���J*!�k��Ҫ�9�_M9c�����ү%����!
�IF�:��R��͖�sKk��5���"��8���芅��h�t��l�7��n1���ĳ�彇6#��FT�JN���QLW�Q12�u��c�܀�1j�"���V�9t����Oa ������V�N�yq"���"4�q+iѸ���^%x?oY>�u�YB�?�Jlֳ���:���\ �������� �~�]����|�ǒ��.�����`��Ϝ>�+�)�&�M���د��$�:�����o�����īu3G��3�j2}]i�Ǳ�YԼ�k�='��N����y�.���f}���.0��Lb�$A�yxRq��S�"��;��ct���8J^�t.u�C���n��jλ~.�j)w���OqXJL�� �WU�4��@
�u\@R��N��h��$9:{plj����ޭ�Г��
�Yt{��m����X&c�<���$Ң8h�Oَ[�S�vܝY���n�y�#0㱕%�o��h�b���P���cԵ
��+��N���Vk-�ZJ���?o��իڼ�cN��<�F2��%H��98�Î�2^���n���m�X)ɓ��77Re=,:���1���r�"�0�pM��>����[	�#V��d�6V:���H�ۘ��� '���R���m'|`P�[�h�ח�
����u&�nN
D�O�Y�mS����s[W��ƹ0�2�D7�_+�j�����q	�ed;whV)����9Ee,���+���:��ӷ
��T�N�2��s%s�>�|!��;I����g�#��Q�Y���&����׫(�w���N��A�E��H�F+�.�v�u,`���1��a��fgbUD�W���lm��6j�rY���A� 	N���2���R��p��pf���LZ�IˌV�3�6?n� �d�<�W��O�<�i%�0x�7XP��w��G�S�5
ow<�y��)6��u�x�Z�<NH��ex��u�j�
@ٔ������@�g��v�����A^�
�,>���6��qj����5��c�0���K��`q\��(�[�C]��q��Q����t����*$Hl�zb�^�\�=�e��Jm��Փ d��J�jk������2��gE��U�����V�q��Fj{t�nl|�E2��Ý*{�,+nX��z]�u��*��N�^X��{�D�Sh�2-��r,`� 1�3)�Spf˂(�u�v9��Y��_I%���M@M��4���/nAL���Jj�n�p�-��5��_Q��T`8�a�0�=w!��H��閼�z`��%F�	v�R����-��2a���?TL��9҄5��lh�4Xje�bt�u[������Vk<+��G���	23n���&���:Մ�T�G���WJ�[=�����>X�F�CjӧR���,U\ˈ�_$o��ҹ_�`u��j�6i�B��c��ܽ9S=�QkQ��S�ICUn=�o{$�ݺ�S�i��ѾYa�ۍ��@�CVo��r��o������ĸ�2fJ\��
\Pt9�A�a��b<�C�L��\cv�Vq�����!��=˼#Uf.�Ok�޷lw�^<%2�
����φ��� k������L�u��~���� �o����Os�_N�q�4yU��QZ�G���!��*�G7zZ�@=U4$�F�"�6Py9�Y܅����J9Q%Q����;)ˮ�Y��~eK�r@�{�eo^];v��1��������U�*�ځ�I횉L��pp���:������kb?/qU����mn��z�f a�i���$��݁�V�(�>���mR���]x�]`���Z�u����$��G�Y]���ǖ�B��×v���4b�:�'c�j�S�Nސ�F�dй�r-a(4����i����:JK����Ϩ�׃əR��}=�tﺑ�馥�QB:���#"[�*������-z�Ӝ����m9�^/Kޞʝ�c͖�As"�7Pr�S2%)�S��tӨܓ�x�rܹq��T��O_M�J��e�e��j�aZ�����Js�b�R��_F����Z�2�'��J���u�#�n.�Nn��*��g��I*d������ԯ-e�u�/?Xp�`��,������YQQ[%��[^�.����Sӆ�N�uE:����g�(���Nt/����j�:����j���t���[;�4|���q&�uwvk�Z�m�]�ϵ�˘�?fú�ZVL��!�7(1���v�Y$����
YX�T�yQk�dg^���3y֯��;,w��k+Z����xxS��&����4὾��&�I1��̎\�w��^<��w�Pֲ�n���u6Χ47{���*t�H�����Κ�db̘ b��N�]�zr:���|̌���.Rg�]}�z�ܼts��� ���pF���M'�l���p��޽��/y�3�B#f�/�z����L�k�0��K� 8�Y�؇2�g]k���*�T-:�ی�9�8���OBoG�*e����H��rN�V}�I}����gu#����GN<q�-S�%riպ�N�7�h��2fIym,!��U*�[�[���vbϻ���s�N��f����tA�"�ʫB(�[��r/p��6W?�,U�zj�
5�-Wp����������w-B��p8G���3�S�7Z:��l���Kd���m28���ڧ���Rks�m��7��l�/�=<Ԗ_�?q��΄��eYZ�hD�I�olȫ�����t��֠�NQ��#���]9�z��X�q_s��^KeC�B@�(��&z��Q�i���pgX�b4�QBD��%8�)��������';��U	�r��q��������Gr��D�$,N��Vl�/r��z��Q	5hd9t�����*su��M�����}�ڰ��N�xW�PڨY(��Լl����q�;Y���ݟ��ɧ*J�iJFE���Lx��CVL�T�MF�H_+lĄ�8�o�2�od�u;�ɏ���t���v�\_s��E�|��}�N�]Q�B�S���mp�< ��F�;�B�c�s$���AR�sA��
�Fkc�'t\���E^�\n拣�>W)��L�wA:������gR�l�y�U���v��ݷ=�n�f,eImr�O]�u�S=|�G��L��՘�phڳ��tȍ�L��"��-�������sюV/l�J*"v}�����X��9xP��h�F����!�P��u�t+3g>� :�3�aGP�^�p1ӞV�}{N�f�8E���b�egh�a){q�.u�C�����;���^}cX�ZƓ'�{kݞ6���3��,K2�Lh>�ª�b��¶�m +�uB.m��뙂�)�Sأ7U�6�+fvԁ��y?[��\Q9�f����Q���+�� O�y"9��J���S��%m)L V���of��話`LV�6x��u�Ec��O]ܛ���h�N�kyc6��N�]�z�P���I�2�^_�&xFf�����6'ӑ&�:<�	`��a����,�����L¥2!��_+��]��N{Ǯ�=>�i�ZpQ��":P�k��[�z�^d��c|��X�i�۶�ڹ�K�����E���&�d�~tT_*�Bi9��fĴ�ժ�3d����& �d\A鄎*�/���-Ա����/�\�=4h+7�$Ө���f���ER�2��X7+P��2N�bW)�!7;�}Qy�����ul����zX�g=7�h�S=����$#�ª��-ε���P7�(�����̳֦�ʣ��� v�-!�i��N�4���H�M�5�&͉�y�ڮX��'��f20��(.éf�<�6fI���B���=Y˺�`Ǻ��[�����!.�ؗ	�8:T�]���[�>��RP�J� !��J�Ҹ�RDg�+xAv��ws/�:t��T\�����q���y6�5X|����'������:)I}�jm���k�:�h*��:5�-���mC]nM�s!�Ͳ_B�S2���m�q�M!hjʽ}S�ˎR�\u�Su{��G�.�R�@m��W�uë'R�WmP�v��}N�����������uƌ��OM��1���C����2�',H|;!�ƪ�C�]H��;#��6t��U�(,���/;�t�p�u�f�ˇ�ܗ��Kr�O6��v��2��GP��V�&`g]I<�^���+��P�ꬶ�ELƈ�q�)�iɰ5��W�}���K,F�L����6��Nz�F�z`����٘>�
��O��{(�Y�H�j/0M�:\���S ��Q4��~����j�X�CVo��r��j��,pJ%�l?,�;%���\�qo��l�IO2��wI����o�n3#�?8�7x���c*�.PB��|O�vڙz�8�̹��K#p;7�Η�v�M�)p�<�8�Cf��Cz��t���R!�-2ؕ���i,/pSr-X�v��zjc�q��f����.���j�����d���1tذ��GM�W��x�"3Ǆ�8Fm*��4��*LE�)�u<��ƈWXf2p�k���ԥ��<�KV-FHQ�L)�f����s�.��J����	�1�`8���p���G��r���h���ZT�;���Z�$ʁG�2g%��=��(?b�N׳}�(�0NY�6d�Z˲�t�cq���1*��	'�:@���0T�CBE �v~̝$lvS���ܷz�$v«z��g��9�c�x>�Fо�G�����2Q4#�jz��D���J#��k�eO��:���<���b�m��se���`����uL�D�����N ���n�k��p.H����uΡ��e���k��j�.	�d�?A�y�G�/3^{g�� =�d㠕w@������.�N㺐w�\�/�z����K�hE���[�)y�Τ�&�b���<�x�/w1���L�2�3n�\��H*��O6�V�lt��.���N� A"��*��cg�ڂ�⠽6vs�qml������ܳO������6z�]:
�����S�ݡt��	[D��4/Ń۞�M/�He�F��au�3�G��/n�����c�1t��c��54i�^�.�PbϺ����uε�PJ뽬p�Rp55���d���Ү_j�:�Z�;�!Ыecqo�J�4A1�ۛ��w�5:˜��~�S"���p�
�UF.V~�u��ᒷ��nj��c[��;���[/:��pT���s8�(j�'�oJ@��҉����v\�?m6���knTń�O������E�����Z�c%��"���;�Վ쎬��c�V�\lkf��ˮv'&�f �eVT+t�7����,xU����Ȥ���gE�xľ�nf������d���Q���ʝ7eՙ�ē��h�����b�{Ȁzf.��;8��۰�2T�q=^��u���~�k���WR}I��#���P�I�Ȓ�7�XҜ�2�Veo+�B�N�'����;Q,>B�S�;�7XtH^�RX�&��Fo6�ӑs��ʪ�	1�S��0t�X�5��8Ԗ_��Q����EU���T�.�|�A~qj��qQ@1s�f�)h�q�������j���Z�#�s��\d��S�B,��+��K��tw��U����A:E�#p�y��
tB�<0t:j��sK��q#��|WE�>n�koz�ΰ68�|LR�FL��2�^��4h_u4\.�2o�J�ܐ��tGl�αV��Q+&1�1�9Uǖ@�4�����%l�n�[����"��}���{4���ZĭpӃ��B��c�ųxv����
0�ًJ@s�r��m���h�[�&�/�D�j��6�$n��ǼP�:���حf�$l<�J�(�=7�{K`�r`�f\kL�6W �	�Z�֪�d���}���q*DG-Q"ξ8vV��^Fk��B��%s�F��%6��
��iY�mn�ᄀG��q6RN8t`A�Ahʻ�{���/#�h�s��:�p���h��f�X#6xL����»�v:9�5�d�ʤe7���7$��u��f��4�̭v��4���s��n�-���YX)�<���u�7"��4���X�[��FՁ��@�`A�y��_Ɇ.\p�g*;l. �ꝛ��<n\�����0�5hFf�@�O�[�Z�19�0X�C���|{9��K�x��m��-̢&qN�o,�s�k��&���J�dх�;��K�*��ar���Y��z��j�e��2�x[6&�5�з)�rAi�Z�8��et�n�H�4���Q�#�l�u%�3M,��u^�dn�7\�O_I� 蔀��v���8]�:���˴��a,k���i�օi�p�j卧2^�AF�2`��VV�ӥVR�����GkI̪I᭜u����V��KQ�6��LnS0l�=}y]�܅�\�\&�c�ᖖR�r��U�нG��<mTc-���w6�TM��i�#��Y��@�z�Q��Z]��+��ӭZ۳�^��L�K�M�2��J�W�A�����#�d�.�T�0��@��7� �X�ɕ�U<�%`#�:UyD�at015ی1s�L]�/i�� rvt��4�[��ז�6V�,2�+�Fn�o�vQS��Gm�5��.�A�s�BRG�����P�nje�BҚl �O�1 �8x�����.J��;uJ̦�r��kw{k��;�muZ�<
i���d����{�#v'bQϋx�晤>�``\��.���9�������`�ζ�[79ݺ;�"����-0��T��/'"��+pլ���՝�����1�4*w�k;tcrf�f,��]h�9������2�:ڙ�8@C�r�k#=	P[�"�	����L�.��uwN��s���:�[Dg	[P��i����˥�nb�F{wJ f��zY��`��Np�V&�i�BF&���a���*�a�<�]u1@��M|'/���|��H2Vf݀)�V�J�d��q�F�9������D(�`U����S���z�� ���FM�r���҉�1rm	*�z�Xx�Y�z�V��;nS�*D�Y;���g32��os���*%�[��,O�Ń�\	���;�r'w5P�N�jȢ�! PA��C)*�i�R���¢4�_:��G�����S	"�3�ȫji$]3:sZWS	YehXW#�)$(�֜*--F�Us�d�PF���%�dFK�	�tI9uLӡ�&dhu�Y�V�S�b�E�ʵ��@Rʂ%G$'2#3�PE+���Q�J!��E\�������8�r�!df
iE���ΰH�P�KR֪+N�U:� ���j̐%.=7K�P�gQ�*����NU��B� ��Y�\�R��]wU���T�cT����Vl�e�BvS*���\�s<�J�J*9rSXU�6UY�V��n�p�#KSMQ�D�)HU$iZr��H�i3�E�qp:��Z���.Td�(�
�Մ��TID4(�Ե.E�r䔕��D!(��B(=��VZ۩�QU�B֘KH�LC�!�Ss�revnv����)��).�]L:��a�zY:�;�Ƴ^*�K��·ҐE���=
�ɶZ�y��~Y�V~�@&$��$p�&O�{�ȡ'�9���Q�ߟ�y(��v�����?[y����܈�Hf!|�h� �1{�LI�D�"/����b��r(R���Wv���~@�f"H�H��}0�� "ݹ;��1���V������0��y����]�Ǌ9\
o�`������F'x�>��ǔ���ro �}O�8G�(npG� xG�_���̹٢}�Hߟݛ[[Om��" ���A?�������<��������S~Bt�|���M�	'x>����7�9����>����;I����y:>I�	�Q+��,��B� ���3��9�q���+���D`�DF��#�yv���s�~������®=}�Sr����x����v���ݷ���q'�������7�'o;�}[rrnw�j��yI�dQ�1@B?��J�{�L��×��)C��">����{m�ܮ��߃}w��o�^����iߒ4Ɂc~�F� `c�x�������<l����9����x����O{��1D��I��4�aH���al��䮝|�է¶�Z����B�#�L>cӏڏ
��i�y���w󴞶���_�ܜ�z=��xM�	�����w�bw�k��6��OI��TE�����,� "u��g�"eEcٱ�Ǵ��X���}z<cS�ǔ��9A�7;�s�Oh{�w�®��Ʈ�!ɇ�z�|��2�On܃A�9�ݮ����ޓ}Bt�y^�y��S~BOW�6�����~�u'ѓ�u���=]���������;ô��?��{�8��=[�zO(xMz����~C��{C��]�N�����0���>q����Гz����ߐ���g��N'A�<;��RoٗW�}�ʺ`Sb>��}�	���7��m�97?��a�~v�O���7�o(��cӼ;۴��z�����ù]���M���o�_ףŃþ��y�z<;�yL.��^~q�=8��C���j��2���u���^����g�]�P���|���1;���?��9��}��þ~��Ѿ;�����U?;_c������G�<��;Nޟi������v��q����nNT����@Q+l{zV���b����|V^�A����n��0"��Y��\L��8A.U�sb�C�4��k�"�8���g�Q��½Җ.V�:�+	���1���'7\��"�M�(�Y� �-\��xڭaX/Ve���p���X�������y���e���R��m�{�"���G�>�f*��!B(_�z�뷔�˾���xL)��}��]������I��'���ϣ�����S�O��~���=&=���/��������/'�nGcz��������/�:���~�b�#��A"	�  �rE�2Dq����Ya�������m� ��bO������`�8�a�C1�#���\��_˘����|~��N��&P��������7!���<�oRq8����7��oI�������������o[����|v�<������N�v���?p���c��W��F�����k��U|7B�
"�2DYO���7�ϟ�yw��]���='��C�y(?'�O?\�����o/�nNC�ww����7��}��0���o�!�<Dh/��'�$'��R����ջ��7�I�1���c�>1w�G���nܝ����HO�y�c�y����P���x@���i7�r���L(}���.��toZ��>b�$G�}�u,٭��+!�z6�^�9��.�D@&4�0$��� Y	������q�v����$��?;u���O��t}~;xM�	�~>���1&��|�	�۞����������z�LH� ���">��yN����m��E>������N�?w���r�^﵃����?��NL.����~xޝ�����&����}��x���N'�=$�Om�<�Sx|&��9��A}�$}9��+jL�We���>���|�P�[�<���@�ox�;|t�������ϟ;o	���ɾ�����&�{�q����}����ӎ|!�z߸�P���_m���I�"�ԍ.�;gf\��	��<��?�s�ۓ����ﭻ��C����(��x�$@6+>��G�1�!����򟝽��I����)�!>ݼ�����0�����>����1;־��V�_P�����[;k=�2�kU#�>c�2~�;Ӵ�_n=��ü;]��ÿ'8����'����ǭx����|x��o/��9����c��$��>����H�w�k���˷&���ycA�uj77��3�6�#8�>,��eR��ϖ�)�f��ݹ,�5]����wrm�x���u@�^�ܤ��u�{�+ܡm'�ӆ�����@5 HҍL{��Na�K�;W.<��r0Z>����|�,�RJm�H��٥[k�����
"�}�Y#�#������'o�x��?��<.�� s����9�����yO<8�ǯ�97���?�y�w���~w$������<[Ӽ��!��|���\{BM�'�y�X�Y���Ŵ�v�\}F>�'��߯�� }I���xğ��ߟ	�'����)�[}N���zC�a�'���yw�Ǹ��nt�N<�q�7�.��w/����<����x��N�ｇQٞ���{u������/�(}>b$`�y�������C������$
���<~0J#+�,�?~1D�>x��_���}��<�Oi�>X��7�9G�yv�w�������H�g����T�V�u[�e{�D���D� �1b�l���@G&�s�����<!������M�}�eߝ�@���xM�����G�����S�O��;�o�Ʌ���}w���90��n�6�n�ks.�����#�$}"$}�����I��>���x@���8R�{v��P�����~��;ߞ�P�׾�����]��@�����.�i�}��I�<���Wz����7�����gf��W���;���}}�#DzozC�raO?o�;˼;��׫�$$��e0�����x~;y@���y�ǗS��7�Ç��L+��dE�]?�#�<cLB1�j��FTLvfj�y]h�z�����|G�>�?pyM!~����~�J�S~w��G�P��1;������9���s�����w��	�]�S�?'�9��$�]���x���#?P�	��DJ��= zu;�Qy������W�U1_PT����������&���������q�I?;{y�~�㷔܄�w��yO*�S}�9����,~^;U���xN@���C����r��Ҧ�����Ǫ|P~e�SKB�:+�u��1�����!�FG���q"1dzkꃓ������~8�C�c��<PI��z�����;ӽ��Ǜ}v�������S�|�
��Ǿ@�@'7D��ֺ�;=>�"4}#�Q���p�]&��7�����_� ��!�$��B-�d�����~NL?�ݿ�����rn��xW�N<�w�<������x;ri��.��Y��yS��$A����!�ح�!y6�j�n4]�� �:�Kt�X�W��}K�e�9H8}���h�mA�+l;�C�p�y��W��-�#���""��o��X�ș�K)�BZgH��R��i0z�1ٝ*���DC{�q��P�%SûR��?}��Wfd���^�����$`����蓼��0��J>��܄���w�����.�����;~t�����xM��������p)����<zM��bO���~M����9�X]�����}{�������z�c��ᆻ���� ��b(F���pU����;�ɹ���[�xL.��Ǫ<|���&����~��w�TD��I&,Ɔ� !��ߺ�b��xD��_}b$�@�g�׀���J��_�Ur���h��c�D��ރ�����V����L.��'o�~|9w;J���97ރ��5��bw������xL.��Ǆ�C�q����X��GL#ٲ<D�D�|�2�ʾ��z��s�C�G��u�ׇ�nM���x	ӵ��<���~BI��߯�}����zv��A�������ߓ��|C��W��{NO;��"��a��{#� 2"LF|��>T�Gt�N�{2���z����>���h�������ǅq�	�w��ސ�~F��������ې?������q'��oυ�c��W����='��P�y=��o�o	��ɥ@�����{:���7�/�w���l�`��ec7�1V��c� � �Ǫ�1�~B��z?z��|M������;���?|����
�z�<
��8/￼�1���ɹ����{��aw���j����I1
P�$�{�F�?�-^�z�|���hď���z$�@��{C�o�ÿ�����Ϟ��;zNW�����;rw�==��[y^�x��Ʌߝ������r��Ҍ��DP���"G�#_��1������S�p��Ѻ>��ɸ]�T.�^�b>��;{O�S�P�z>�r�M?�?�����	�>;rԟ>~Lh�������s}dx`��&z׌���}d[u�t�-w����fɁ��J�w8h{=S�Ŧ�2�����UF[`w_�} �� �D��`�l�l���`T�������pcMO��R2�失TJ�U
]ENH����������]�A����7���fҏgW�#�.�J<>f������#��$Ā#��4]�lɛ���� �ԣ�D�QΙ�����0�-#h��%��k�e���ۨBkD����k�F�C	+X�]:�	/A�̽���ܰ����ܶ/�諭�yi�޸k��7?y *`�ON@�<�{p���J�쉺���	�U��'%�e0��h[�3׋Wo����lk�HBLz!�(M|�[��\�Q�*�l3iSL+S�`�	;���1NZ3R?,UX˧?K,h���i��#J���>��-�v2�y�h�CM�:�!8�T�v ��"~�0��4�S���k��_/�Ş�7��+J�s��� i�v�,�?1K�-D�@��Q-�q ��ixV���>
���,>K��P�@�U��r�H��:U2b�4���\MA�!�?w�����Wq�2g��Ok|�Ȫ���᪆MCn��L�
'�ꜩ���H(�GT%y���][�"�t=��
u1����|Ry_'�C�ԾJU��D�z;�f�j����+]g}����į���_��X��'���?O���/ �zj5�\.N��c?"y����P;�UT��jk�扶�,ܙ������Y�
Oyx�m�ԅ��g�.�~�Rw��J{�Խb(��f����νdV��s.Ip�fi{�%���+A�ӻ-IQ��r6%*�z���]������n���!c�Sx:�:������Vu�����Y�����K��N��-Yr�8�S���u�
�ҙ'*-�4���U_}�N,�7ȑ��*3���D�ٟ��a�uUM�(�;�H׮��s���	љF*;cދU�{^�#N���{�rc0�?g�ѡ4�7xUu�}����j�n��d���R#��ձ��G�go(X�>�Na�m���n>櫄\uΊ��F�3��\K����Z{ V��1��ŝ��d�%�;��fΪX,2k䧙���t��:���ɹ^6-�Hh���Ǽ7�yX#�\��w�{�����R"�k���t����e��2�ۿ��V�f.\����]�ˤn�%t�\E\���&��3@NV��۹��܊2����!�t�d;(D�wO�l���E�o^}
o�xޮIm,���zd�OjL`��}cݾ�a����h���{N� 7)i���*U
�\�j��~2�)�s�c�Y�W���؃C����;Et���`ذ���[��@[�|�'��������v�,Qxo2��-rkn��$Fq��+��'I����A{X�U�R�g�'��-w�)=İm8u^Cp�wZ���g�IN7�P�p�Dt�}��i �Н��:r����Z#G���P Zh��7�<��=��;��&�^f��L�Oh���RE�V9������6��<�)�o�+���λ�N3{�K���VG~�����r%��a��O��i.wV��{��-HeG=��m�p`3l�Ы �4�dfm�X��[*��7Ϲ̡C��U�>�5�� ���Cu?-{ԏX]��
��Z�c�@�'�]m���~Y漶���x;jR�������k�U�8���/�1ƻ���s�m�:�z����thK'{��V�HԽ]���>UWѠl�>�j�gשgݻ�'=�^�1�W,`��0�׏D�AlΈq��fVC��t��ĉ�u"*0�r�dfL.��h�]�Y9ٺyM�8����=��ڶ2$�x�o���^��\�¬�#��٧D� v�2yT�u[ϯ���*��Yv�EL�J#LF���`<�%��l���5!ٌ����qFCڕ�:5��(�P�&~ڝ���>4�58vXw�ن"�)�X9�;���\ct���gP��XmP�{�w9�F#`�Q���.��(\Q��Tm*����(�?��#V��R&.ֳ�Z�1S�Q�R6��h��SMvĸ�@^|~����xޯ+g�_*Wb�:��nY�ɦG�Yȡ%˕�z.��0�m�P���]�5$56����eYtnlԖ��T�c.��\%�P�e���
��֍��)Nu.�kc�/��k��6��)W��	�0���\�h �NyW�qӔ+�A�˥�:��I���%j��g�ﾏ�e����0���|&ˌtۅ�����ۃr�ii'�)��jdЬ��).S����X�\\Q6_³g�r��Ϛ��m�:�}Dm�*��|�U��M%�J-x ��e�G���ڭ��TH��G�1Ս㐭������a�Ӑ��m�̣*�"6;��Y4�E�!9$?�*�T����5z�v*vٌ6Z!�������3ڀ��>ҝ��$������>~�RA�hg�\�܄e���k��1�VY��D���Tv��3M�U"���RMl�Y@��`��p��@���*���A����`bg6��K2N\7�Z#(��yS%�,y�W�
sD�Zx�`��a��t�^aXk�݋��ɫ�S�19¥�F��H�f���p|s�	��,���O�,��~Zk�c�bS�������G'�1Ua�y���VYq�ϻ�&���0<��d?c�l:�֕��^���}Z�.ɓ�s�����f�����<r7�3�J�ò�N�x�}�w�45��&�7ch���<��M��z�;g3~#��*O�:G1<�V��:�e���w"f�0՜�}��߂�TJήΦ�zG��Q�w~�e�����B-˧�4@�d�<ͣ�1�6i.��տn#v�L��zp����㤮��ͮ��i�n¶c��}GѲ��9IЉ�L_�����"���A��͎�@^�p�����;����$Z�S�-L��|�b��b�T�`�3|��t��� <4X���|P�ۘXw|!>���t�@*߃�UZ�d+��M�E��%�!�}Ҋ�qW�H�N`wW�ފ2�x� �#�r�����'�}��y��yLB�U��5?gmԌ��:v"$�5U}���Tʫ�ĥ�AȢS�1 鯡껅�@�ON@�<{P���1�7Z:�&&8�I��9��n��ۻyI��yQ��*b�����9��o�5%��4������&�[s&���y�Ysg���� @�ZsJ���~��U��_MD9c�����Ҳ��E�i:�:Ѧ<uOaW��=��ﯷ"�Љݠ�"�x���w��8E<�Ӄ!�W�
��1����u˄IC\'[�{����g�K@����X��ޭ�u�N��UΣh��|%{��'ˤ���Ռ!����]"b�1��P��
����^��q�	v?3u����Ѩ�:7w��!a������ݨE["�w���B��Zm4_c�\�n�՞{
�"y���Ur��f[k:j�M�0q,"�tk�J���v�=i}��;���͐��a�gB�A;I�ܼm:�B���h���g6;�T?�諭�:�j�RqN�͝�5!O��ێU���p/ :`��?*�&j:Q?H!2׏=�:�h\��ݽ�<&����uu0�����{_К�*ԦL��7@sϡ�خ1d��I��;����wNy���*_�'T����'_[4<8��9G'v�k?2y}j����R�:�']1�7�g�d9�ʻ{cj1{D*�2j����A�������K�Y���V��1,O^9R�X��ﱝ듽s6�K0��n�s2;�Jk
��d���Ћ�)��E]��,��,��]tN��{��Ƨ���a��_/��BJ���H�0��j������h�-˪�ٝ��`̲vh��'�2��d۟���S�5��F��|'�.����O�6��L̋1[����ܛ���$l�:��>���>��^Z+3ʴ;-��T�\շ��:a��v�Tf[9�^��g�u[ջ�1�j�E-u򱮘7��6��V;c��(��7�">f����*�R�ut�,Q��z�8��
�=���۶�ι�_.v���:C���f��П������x�vH���ŋYVxh�ҵ�?�8�,��L|+����mv��К�֣n�|
�j)<���Gi"�i���܍�l�M%�O����`Bl�r�iu �z�wP;n���n	GN�<�fP��f�)��6a�jj�z��v�����5켸�:��}E�F���4������.������=�fyf���M�v�g�����e��%�:���w�i��O��%X�E���H{,�Έ@Mu��]c\Aӻ]���I����)����J��҅ѧ��O47f��5��U1Q��-K��H+��
&9��Qdܖ����9���VPͫW)�n�[9IY̻�v/3k^�;-�B�7@άOG�@��jk�E�/z^f�yr(�]ˆ4�.L�Z�Q��O��FҼv�."ٗ5b�g��4L��QM�nƆ餳�Ӝ[�&]�W����q�12������V�f�P�e��)�q���6����)���D�OY*»2��÷׼tEKq�\��;���5��4�q%0(�.ȫ���A����q�Gѽ�S嵖�]���U���N�W��;�c��l����c&�>;���%�����yNr�g��dF�[�r�+�Rv��u0�i��`8�S���ݐs��3Q�1�=�j��j�*��B<�Hݞ�5T��[6�V����<t�x��H�V�=�{�J��)��)oA4.��A��9#��u4�;�6�7�,@�r�qt���2\Y�Yy�NYO6ū��P�Z�XF�f����Pu';ޚ�VvVV!B��z*�;j����wDŚ���s,���.�,�v�F�oF=#I� ��y�����c���c�u��C˯Z�n��s@{tl��sc:�q��1e fk����t3h�`۽a�����QY��Ve��my��q�Om�um��m�B�QY��۱�i� �����'rW)�O68�K@ά?G�E�]qX��8�r_^_`��lǬ��#��w��Xx�:Wm�ޢ{ފ����E+`��ug�.[F�F�a�w��^�K�AF��"^�E]*J��ҰyՊp�8��iKvc���YD��γ�b��-s���]y���^���i2�z���,U}�'��R���[p�j�#uۙ�u�Vpee+�f]k��T�;�������T�<��Τ�c��k���2��ii\���L��s�f_^h����Y�(^1s����l�x��w5��U�����5���w���f�]�n�}0�ua�/1�S�����Y.���q�2g�{7E�����5ծ�R�,�FYw������	*oE]��,�����̠��{���VR�6�É�n��H��uǻ��,��f�r	+��̕1,J��ڗ����1!i�K��@�+=��K�I�Ԧ��䨲���A�Y���.;�.�Gk��4J�T-!q���5������z��$#$�D�`�1E����[�
(���Ω:�D�"�Z���5-,R�R�"�K9���""*�E�9RBi����`��I�G1$,HB
,2(�Δa���3H�5B�Դ�SYQ(k,���TW*�5(�2JI(ЪH�D���r2TR��\L�NQ�Yha,YUDVK(���#ERS
�
Ќ��Y�j�����ց]�Ge45eQ� Τ��q(�T)t�3S<��U������*�Ȉ3
�,�9B�V�Qf���%4���ru$%K:˜I5e*�9B�j�Hh�&E�S�8�eeY�1M��K(��J�',R�g
�a	Qt�:Z��VZ$ZBfD��Օ��J��+J.�5�e:aM1���gL�������ЭH�(�Mn�"����u�np���"z֬Տ��n�,��)-�]���Qy��>��!�u�ױ�J�����}_}_WܹG=���e���^B�5�mE#L��ҖL���$��u!wC��(Ek�U�6ģKs/�Z�P��mw!���и�^UӠ����@R�R�$�U�+�af¹���Z���(�����Thnr�Nxi+����N�#��Z@�K�����~� ���Y{��n�q��W���"Q�_B��BN�9gD6p��ڬ�؅�%��hg-��ޞa:.���k�H��!j�^>��_+ũ�ҷ�F����K�XD�l��o]�����-$�
�k3�5�.U����/�V��Ha�0�I;2a@!���ي���+w�ܐ꥖�հ�^���Z�P>����X.�s�x��3���XU�@�#�{o�'A�2�C�4C��ׂL+��.��]�a��+�i�^�^ۣ���a����s�)85T�^'A�X�,5�1"u�H��(��c�ӻP�"D�i�|�Z1��Yh����#E���m*a9���捵u��eo�DGZ��������mC,���:-�9���7��M-�,<j�v*������eb��z_u7t;��3��{D,���o1����&՝2\��	$H��C3~�[9v�cs
��v��8Vg��Ҿ�����+33�+@}.�I&���G���{���UUU�ɂ{�=��2���݆I�'���[>�\�'go����7��0�+;0��d��̤�4ǽ�ٹIh���叡�e��0�56a�H�,�2���hQ��ޗ�F6��Y�0P8~�z�t��)�<+!Ǵg�c<�:.�&�=YS��,N�?�O3���������*���QZ�G�����OY�9a�~�y�������*�RO�-�RƝ������x�IUf>|P�ݛʃʝYF������u��N�%�~�r���jK1���zn#23���N�@jˇ�G�9青�=�A�zc�Tq���T�E#,�s0�i���n��eu4._�ҡOvm�o�L�"�D�?KU�)�>B��-��ة�g�{-�X��r�u�vl�c�f�g*�2+�JR$���DĞ}4'���#,0���m1��"��5ٕ�W)�x�&3Iw󯫏$�\N?�U��m�#�ȿ�]��|�K�����z��+��%_&\�J�e^#HwE"�u����3��aY޿?MA���ں�w�Z*Pc�����R|�a�Eˠ�n-	�ۼg�aV_\y���f������5��Br��[~�H����ͳ��Џv4`���䑊.�ļ���6��>���ٍӧO�ت�a���T�y�9����	�"�q9t
�U[�K����du\x
���S��1C�.��!�c�5W&� 1I�Kŕb������姾�F�L��]5a�V�xJ�K-������t���>.u�٦����$��:�hs�O�4��=�Sum��82,��f���\O�q�>�k�=sۧ��zZ�-P���LL��d'��͝@�zt��0�NqUYg�<Y;}����k!����[)׷�S:��ob-��6����l���ӫ��(�⫂�<�xs�����[Q�NDw$��m5]0+U�+����L�B��tڹ�Y�S���%�~�tN
�Tsţ'f}z0ț#�@���ڲ0��Wc���K'���yLB�u\�S�v�H���t���Go)T��[V�ڪY?��"t@���s��D�ˇ�	��J�숛�d����3!c�ר!�`tl'��q3�Bs"+�ai��H��[�Ԗt_�~B�N�Z=I�����U��ל=����N���2cʲ��+�Y\)"��ǖs�۽��w�g=`�t�-�32Q���Rm_T��
��enÂ>Rr�7����u�7�X�{6�Zk,f�z�:嫌���F^�/�������Z���"���?ݢM~�r���꯫�%�(GN�=rWQ� p�P:y��)�V3��}4�-�v��'1[��&���(q���쯜���RQ��څԌĠ�#K'y�as�Sέ8o&kl��8'�t���+�6��Ϝ3���}[�X���(���Bb'�u�.�<�"3��շm�[qvn-��K��r���h��q52:APڨY(�,SWX�u4�M7���EӔ�^50�	��U���p/� �h�
�I���O���6�C��ݕ����|P|C?x�;|X�8��K������UU�L�7�n����G��P�#�(��w\|�*,��svh��4AΞ=������]Q��/=.Woy�5~?q:r��`1ך�[�jM>/;;��?y�/N�Vea�9P��eVG����Z���,����x��60Xe$�b�xz����n��[�k��p0�T�҉ݳ?90�ztt�v�Y�"�z�^μ]��̘��\�3u�{�R�Ɍ�e���A����B����c@�[�Ϝ�����X�.3�A%�c�hY>>{S0�n�Ӫ&���{�&iHi���Y7��ԧ��b2�p?u3e��Ye
�I���Y̛CwF��Ef��QAl���2��X������){i�@�]Y��+yٴ�K�8�7
N:������?UUU}��7���[z&gY/ L �i䋧ʽ�ey}=�V����lX�h���'��}��9����Ʋ��}m.>+ή4���u�CDk��%#̽P��a_��t�������=Sa�!�@.��	&�������%Z�!]~_oP�S��<��WHƺ2�	�6,��WwU�W���T)�+
d��3Q9]r�GfT��ĉϗ;c�׵�[���4����Kp��c����Cރ6���4�j䖔ɸ+w�M��V<��z�>��r�yY�K~ž�B�c��`o%�
5�������T+%�}�� �I�3�mV���jEF�\�*��=}qW�:w-�S�	�N3 [�����Mww.��TPC�v�]x�#�T����Wp�+v$��5���|���C���/kjlhAF:�KJ��Z��������RڸHZE��z�o����?��rn��Ys��f7b�[{�[���c�r�
kfdVf�7p:�WҦ�a��a�rBq�h�mj���JS�=Pӿ'[��&q)�T�w�r�
���4CK�K��uol���*�Ev�� ��ɮ����!Osؒ��l��)��cob�҅��c9�CR�!�^�-kUc�ʗR��ua:�����FM�W�縁)�@���ޭ�^���>�����r���٣'��}VL���)TjimLeA]hT��64��������M����S
0f[�"{���w"�d)���(}q���q>�5۟�~t��ـ+��xѳ&�v����E��V���VX�����M���P.�Ɛ_g�B�q2��z�G�]���1V��ź���}S1�4_l�o6ձ ;s<�|Ѷ��r��^���0E�����[��#4_��踂��V]�ȩ��G ��L,j�*��N@�l�j�ص:���L��ѕ�ĸ}�V<?��k����s�[����c� ����6a��Jy��WU���鴊�{J��q#ni��7�7�6�C�P�t�qFCQJ�+���ogM0k�f���y�nс3���B/��3��>�Ʈʔh@���3&z��xޯ-r�ąԛ���o��g_�p���.�(���ac��_<=S�� Dt��Ğ�@����=�M�>�`J���j�Qb���U<8Ԗcq�U�Y*����'l}�-�x�ru{�\���po�ATP�o��Ag?9u�>w�7��ul:�ޏD�t����C=F�;�r��+�Ԝ���}	A���O�[��+�[�5۰�?Q��U�^rN^� v5M���VJU�(TSm����j�joa=�����U}�Nee/W�1`���tO�L!4$U�*��r�qWY�,�c��ruE�dd52����KԳ�q[�[�S�t�DNqrr��J���L��5z�vB�m�ρ͖�a�"�;����5\��Ș����F�⃮H�(Z���B����߸�C�?a
���l���圧r����N�8Lc%[��2t�v��s�=�*N�&l�1QSGn����ܥi�����!:Oڒ�K�X�}`���D�ie��V��*�W���{��JճY#5�[eat�ڸ͸b*<�15W&� 1P��4��eX���&:Y<k�s����6XE��kl����}(�7"Юp7����bsi_#�鏤�
��r���i�P�̨F:U�p�D�}s�%��V+ �F�?v%�϶>�t�gJf�:��eL<,buZ�/���{9V�S�uL���E�Mt�/�X6kK&0B"NqUYg�œ����k!�H��F�B9�1OL뮆�U!��gRLfmk�5~�a�4ۢ���<�s��m�\:ǋ�JƫW�evi�����C#��`4��zf��љ�bm���NF�VT�c���)0I��Ep$N�]�ч"��7�����9�N$�[�Ӓ�I3]ط39��h%� ��Z9��td2Kh�1�z���0�/V�U��=��pB�e�e�L�_W�UU}Oq�X��A���G��uI��u�a��`��aϡ�}Ҋ��8+��t$�嵛�΍�G��n�א9]��crB��Χ��+�U��ɺ�{n�e��$�؂$�y�N��V�K:�ںE����'��U�,���!����3��w��j��N�#��m��ld$;���T�'���[L�6H\�r�Bk����e�z~cb��{h���8�˜��x��54�X6=  @l�fn�G��U��;u�Ӗ8`��{���q�׮��](@l���9U����Ԧ�B'v��Fe�Y;�R�櫦�b�=��z%��l����B�(��:��q�\}�V�W\���(���$&w�i\�6�{;v�������Tg>�Ƥա�9�i��ǒ�9ω��ؚA��P�o��2v�*�WѝnR!��ӣ,�v����|�F�ܪ4ۮÖ Ѕ �U)3�s�]cS�t�ڕ{��}��r�j�唷Sš�ˇ�B�2d�&�mlcf5eLu��5�1�8�g����W�`ͼ���;/�rݨj���,�Y��S�W�L�QTi��'�ٷ�U`��ۂ��S�X�~�[�1]`�[s˨%[^��,]	��O��u�t�=�Y��
@�Zv;��F���KRPw���磌���z�2ߑ����N�g�K1Aj�s�1���gR�"���2����0�d]��'[7|R��Q���p�PY+]����fVʨE]�*��⇯�'<�%�����W;HŭN]��`��A���NtG/�WǲhH��8ea�s!_yvk�n��9����r���$��`�	_ */UC�R���Y��SCt�ۓ�ۺ�w҉��Z�\�EUخs��Y�s9�H�[�rԦ&����y���:*/g$�F���:4�D���5c4<C$��g��K����V� sVu�ǒ�jy����a\9������#{����U��آ>��M���,7���U"*��X�L�0xk��no���.y�ki]ˎ�8��������<tA�ߑ� >��{�ȗ詅��dTl�M�ap���:��"����é�z�(>v;|�(�Di�5rKh)f���튬{Rd��=��ۭ��"n��/`����
K6�h�k�����J�\������ ��
arg3_��іiН�����&՛����Ǡ���/�[Fob�R������2�K2!}^�X�E�&x����ݻ#��T}��a�;D�8Wc����>&�+�Ző@�d[�"�,b7*�i7�0"��f�H�����@ @>�n��\Jn�${V_�z�MB��p��p���S�	�M�+�T��B�*W_	[�c�A�g�����ll�/H|{�+�I�GΈl���`6�`w����o>Y�ܾ�s�:Ր�I<\�[V�ܴ�����
eƞ&6��r[1�ͪY6�47�o����f�ԪF�'vl�̊� qH�27��xЗ#���mn!�����D3ԑ��y�{c5QH�5&jN̛�3�:�qu)JƦ��(�օD����=6�lM��[n���0F;wp�{�"w�������0|��4��p�p�QPD�1�^�m�O8g`ǵ��NX��z��q���mU1�edW�@p��AVz4)��o"�j���sT�\���Fq�:��n�q��U�4_l�n3m[ ��f�:��m]D����̡Y�.�z.��>yS��	�9�2v���.��T�2Qb5cV�ȕ\�&$S9Q�0:XNℸ"q���>�j���e��a/����pY�G��\y�rG &�Tsw�*7q`�ߕ�����I�i鿹�Z�Ł�SY�]zԥ��\ɰ�m��>���Kf�rM���bfwTw#x�r�V��N�9�>��(m�r����[��ȥZ9���C;����j���`[2��p��ơ`��+���7%up374R��-�Yv��\[���m�^��!�� ��{�ڶrԱ�%pᷜ�oj���i���H�t���ӥ$7��oV���YF���#N
Um1fFr����N��[ò]���r�t��4j��C�fS�ْ>u��f�
.o�ҧG��=C)���ҝ)��n���IV�wk��s���Ԡ���ayx]g�9�<
���\5㖥�V.M\�tv�kn�d$Z�F]>z��j�f>��u�WI�r�gD��Р&�9E�bY�i曰_�Q۠�^d��6�s�O�\�ro��'�{1c�ECt�5,R�N�r3l��g�.����D�h�!�Ըa�z��\�;�N3z]^-T�']�+m4R̭X�9���*]�W�o.Oa����~\�j/7�2����9}$Z��K1�+� �am%An<4��Օ6�wS�}q4H!
�o
}�8��v�-GC�>�b�`��e��;%�8���;���<�m�#�\uqV*_�bY�8�,Bv�j��2EY�7r��V���$u���%�a�fŚ�KTEK��]YҎƝj�;E ��܇A���sGv`m���s&��Q�>��[�l�LN63
l
g�J�jf��+�ѻ��	n�<�d�ת
"�/�I��N�����������3�bN.ͽ�W�K�vZ���z�ݔ����;p����Kb��wk(��-��\�s*:�B�Nw.r=c���[��J�.�]&3!HELÚ���>]!W;a��M����a�ʻ3ZU��p{i
$]0b�cQ�ܦx���i���,C�w��BP��b�!@�vT��+~`��]�=���Yy���u
ܾ/[+�Ϧ�5����ۆ�9@2����1W.���ծ�q�a�U�mԵ���zXgw������2�Ŝ�Jw6�bf�X��ׇ,d��8Ί�"�����޻�o1���:P��%�j��0k=�w�&�X�1�u�	�l�=q��GO�mow�e��Mj�|�sܢ�q����F�A�--�����9}b���$�CAŻ��5�+�S/�`xu$�u�n�4l��pz��UE|��}�P��$���t��w37���ʹ���סF��^���.��GX�0��}��#��GK�$�F.�:�M����fN��Mhn��r����2 ��}���'�j�n"�Y�'N�z�X����BU�@�1�<�r<��SW^أ�a��f�<z���]��'B��.�$�&�J�'Z�F07�w[�Juf������o9j��p���C�#�q�9b�fRN��S�����@�{����L��bܘ�(RnPVwg��ou�6B�$Y��HIZhF�(�a�UW(�$�wtp��@���B���G))MUI"�m4�a��HjDS*5�b�j���cL�DI�TŘ]R ��NI.D�W.��EE&r�P�����U�
.q�й$�$��Ar#�h�p�9V�L�bQQk�y�(��*�+�����DS�39�rC�ag3�K<�U�h�V�P\:�E�Ȉ�2��E�Td�Qh��Q�dQg��Yd��s�Y�Eb�I���G*�eR���JН)�r]�.Q&�ΰ���$��J�&�2C*
"#:rT��̊ԣ��J.U DDuuuaU;����ܮR��*"�����L�d�HF�9r��ZӉ�PHH���(��	&	�$�T"iL�l���ou�[���]�& ���%�[��R�t��ŒC�ۨ�bI9>B�ūtsf�t�Z)�j*��g�W���W��n��S
Vt�+�ea�1�����p�BTB�(eFʐ��-�I��;ZӦ���ڊ7�F����H�:�p�*����j��$d���;L��	k=�bx̒�iCf��>]^��6۽��0�c�rw��q5::�'�s$������<�="�_p�w�b��%��~�*��jK1���zoQp���yV��W箺���	� ��x"����"��Ucx��ڸ��,�s0�X~�ۺy��o!�S=��Xi"u?`�GݳMKH�4�v]#2�A�&F��q[��{�N�0�)v#�i��u�׊���{���0ED6�[�fE|�JStZ��	��%=�^|W���Q�*�T3�/��WU�?c���2!�VY-���]I5��ʃ27��A=(�O��^��%ttew���p/A��c�����K�X�}`�0DpD�@2���t�CA1^����kը�Xk��W�p�R��&��� a2���eY�z��\��V;��p�XC��Sg_��ڼ�vr��:w�3��Sm(Y���;��<�un=woo�r.�c�o�Vxn���R(�\�}�i���g3]8�;C�׎ٽ�fnq�.�����V�])>��b<�ⴡ�E�4Q{W.�Q�}��_}_s ǣ=��K	�;?��:<ٺm��x��ʰ<�u����@9s�|6��9��N�ʊQ��.���s6�p�厌?-�f�qt��;�3{]_2�&�'S鍶�z��8�5E@9|q�w���iB(:1bjNuU�~�<Y;}��g��W���OW�7ǛEw���t/ռ��&������1_cʝ7�0`0���<�s>ҞP_]cf�^��#����\̎���.!�&yT��s��KO������o�0�{3O�ֶ�Z�b4+3%þ�ȁ��}c�+���;�#������}�S#)1��]�W]��1��kR^]S�AOTP����0AGaj���9�ӃD0��Bf�Ls(��'"��Vlܪ��D����$ɲ���+i����ʣ�3���椲��J�fJ��V�jw6�t��ge�n�����Z	<|d���2�.���������姠����#��)�k�t��"��T���#J��>���@Ԧ�B'v�R3�ĉż���ѐ����[��pv�ߘ�N<,o��r7�O]!����2Q2M�o,�,J��.Z�]�Gm�~�"�tAЗ��mvP�ӡ/U�nr@o*v؍�j�:?���Ca�n'�X*.j5ز�b�.���p����O@ ]	�75o5b�5�g/��U}��cz.���tN��ݮ25[9���N�����:lK?L#���1.Ol>k)�w�GRQ�J����0�nDQ�u@5&��ˤL\02j�����0�<l9흑���6{��q񈄷^�*��q�ϒ��|��o*�M6�x0( ��l+�%轺#�z�{�q�W������ƏO������v��t�7�Oo�MTQ�2d��B��vj�5�:��R����$�:����sx��WS�����\,�o�G@b��AخiPH�۳\��V��N۬��Y�9`*�v���:(z͉���[�l����}�;���T�pr��>��N�W_����V�aﭫ3�
���n�qպ(�F����K��b��V.+.!�D^��!6̧:�?���7'�}�|�ĐZe��::�d�|
sG�DZ.�����.f[%d	� ���<��Ja�m���o�j�E�\�ї����8���t��S:M��m�V:�{�#*�LCFκ@a���V���눊��J1�n��n��Nh.γXë
�7N<�]��k���_���kk>�Y�Z1
�0�*�F�m�wE�YR��&Zw�ߴ�m���?^�V������x.�T9V����G~�c:qC���gcջ=��LFz�9Ob�̟	����\g��꯾���i��+�Vˬ�hSFĞD�D��A,7�1;n�/wҗ�ׄUf!\p�;��o�#� ��Y��}q��uaUS�:+�_�\,{���mq�m�o�%W*Z�ي1�[ݾ[����gi����(��cW$���L���&��D�W�r=�N,��*^�ב�ՈA/Cc�ݯ���@c�����[*�ܽ��-v|\Z����j����"z.P ����a��W�*����t�8\9�|wb�8��0TC�BF��; U�s.�:{��EZ���K"`�.u�K��^����I�E��+���q��X%J���m*f��3O�S�u�Ke-�p�~j�@��iS���)��R���ܘ�Z뷮�;s3��ܭ�rHV�Y=��U��H:�C
)V�|:�WҦ�P-��+H�Pm`৬�9��N�j�H�gtԘ��N̖�v��g'�Z�[Prc(���z�w��e�����2�7��)Y��Ks͡�;�rN���Z`�_F�uk���Z�������aT;��Dwm���om VJ@R�ׅ��.�`�S'l6�Ǒ�W�ۅ��Ʀ찟5�a��9DJ��:�I�vi�O,jrY�dM��d���q�N��5�5o&tn����m��n=�j��c�/BȟP���UNj6(&'��=��}_UW�s���#�5*̣�;��ƌE����"��̧1@�؆bF���ڗ�}��QW-aY��ZY�.�+���}F4F���L�Fm���I����'_5��V��9�2��@�[^�ח����݊��Wf�?�t|�t�n���;1��`<�'�h!�`Ylrj��!�D=/��l�0�^��=�6l��_kX��/��+����t�-��l:3.zV����D�oe��u)�]�s�4��l�\+�����<6��upxj�\�^+&������FO
)��a��_K�"۔�d;�<���
}R�ŠH�P���u��і;;[�9�y���r�M��V�+|5�ѐ�L1���{p����D���'�����x�xg{z�t3��u%��P(
��H�]w͊{?2���jK1���zq����F�w�j4��;��\�ɃD�l�5MIB~*a��*�U�x~��W�cx=�^��)-�
��й�W���G�`/�ni�D�#�=�K�
S�)�#"Ɩ�p%�>�-i��D8�|�Y�A3�;���X�N�-R�S�&�F�rc�i�ڼ�"F��0�����%�g����%�ׁ�/��W3L��T�e_hq��1�a��xv�wmv�U��QI1����1�BV��{�aZ�v��#������gbsh����q�G��N��to�x����(��1����S�T1�lR�u��	�V�֦..�[/O�_C]l!�Z��A1��n��
UH(��1���â_Hl�$�;.Ef�[	���3p��w��ų�~�IS%�r��W����N�W*�yc'�����)������w<�uOp�#6�\���\���T',/U�w!�cU�!��J��[����	��?{�ڃ��:n������+yVYj
�V���.o��䢰[B9L�{�г�Ɛ���|k�pUF.���-�!��1��{��	Qy����mb�S��"��|��TN���(E̬<M[�\<��w�->'
���1�iU������Ʋ��W��g�j���Sl�'V;�o�tF<�҄w�UpB����:Gb4�{�x���C��f����w���I��̦w�W_f]ymac�� �'}w7ΤLȺ�⫴�� �S���5��QΨD[rGYԧ[�b�:�nM�׈�ےT�Z��8.��'���䰝)e��1Іu�7tM�]Yo�T[�r�!\ޚyA���Nh������]r|kw0�hW�8ڙ��V̗���Pn|��Me\��(���)!h�/N�x�٣oE�������N�ix
�x����}�U}���N�r�ӣB3	:#�T)u9#�w"Jj���w��x�ˇ�	�x�y��cc�S���Q�6�|pHp��Kd�=���dq�[0Y��b���o�n�P՘�w��-��ܔ�Ɗ���2�j88&�V�ƺ ���t�3p6R?b��f�S��z��ޔ�����-�.�i�r4�\b�2�����K��ď*F�-o*07�f����+�^�k-�Ö
���h�M_�^�3�:�&񻃦��Ҍz�Bdĳs��j���F,SH�;S�\E)�s�1.�Ƥա�]"~b�'a��+�V�&�`| �M^�M�j��3�+�ݤq",Ǭǫ��{�cܪ-��Z���1-N�����X�U�g'�G#Q��+kY�����Oo��5P@����r�v�6��
8
�&K������Tq�$��\u3k�1�?�=������]Q��¤C	����p�"�||�/���i]��~d��"sa�Q�+�� 8�z L`Td<8#Tڃ�	��?Uf�)�:�٥��7_��f�-H���6F�*���Wt�+�kׯH_t��������1�=��`3�z��5�GI���ͩ.>Wԝ��D���am�xMu=�~(.;��Ðobz���-ᚲ�-���������0�)+\Vq�`�Wv�����������0�1z��Wa1��<��8�J�ddju�C���p0�}mY�a�s!_xN� {}y���g3N:�F)�UCf�:�v� T^��/��38�s1mMӑ�?M��3F
�;�%(�F���[DRfc0���}_OeF����Y�`	X���%����sU����=}0N*Ɇ�pz;�T�����1TQ(e���Pghm�޻�{r5agQ.�\y*����wµp�����]os�j��+�)����օSFĪ�D�UD�����
�'m�E��WՕ�%s���^�v����p��2�����'NDq�GK�ȃ����p����x�>s�y�ǧ@�H�)��n�N��؟K�y�Yq��&��ƚ�;��AP���s��ڵ�UoC��\�^:�t�YN��k�5�u[��*�PN����FУ�3M�$�j�>�A�!$#RW�u-}5_u���!>�m���L�����Nbm�%��s��~�_�W<�G:��ԚJ�n�ٽ$�.*wE��&0Gt~ںb��=���iɰrgPݚ�[4wr�;5��@0�l�M�5*�I8uvH�h�S��G_f�݌b>t���qt{[�iD�U����y��e�i���C��w j��d���5���[��͆<��]'8'꯾�����=�zn�;�M#]�FQ�JT4�MD��܎)�>:-�
��VԜLoM5#(��
��+�򙙮Zڼ~�6�/oV�� �O\<LΫ���m��=Щ��P�`�Cn5��rGr0-m}2�bާ����6�E[4dP����N9���2{�W�i��e� Z�={"|A�b����N�S�}�+2�ysY������^v'��q�����`:��m�8�e�u�<�A3VL���>حuSS�k�ɾ>�Q�B�v��:E�3.;��E�~�L}���9������Q3u�{ð(�Xӌ1�������5��ҽ2�+�NRD�S~�vr��̯���x��*�m��(�ֹ�mf�P4���_7͋�I��U��nPz૘Ujѭ�-�y�����t�]�5R��X�m>��s���c?t�^�g#�Fh/N�O"�w�N�@=_�0Ҙ�������r�C+^�\,���j��¦�4��x#�}�KӰ�yfK���{PC8��j��{G�t�9�e_	EY�i��%۬W� �ҧ]�>D�ת$�C3�着��@���S{R�^zT��벫�J��9��zˌp��M=��o
�:$ET���۾wc��6~*\��RV���Of�r�[A��2U��U�7�:������%����wϤ�b���M�B����X1���;r]:V�ӄ�֜gT[c*�(�=�pb��������Zn]�I�ڮy]Qu8�o!x���*c*�0�]P%*���})�2Vjq;R��`���5��J�k�ahP�p�F+�����邧w�[�}nV3��������� �>�I&7�YN��ۻ�,����*nm�<�`����'�0�y]�isƚ�֜3P��y��LL�9�o����Y�JgZVD�0-lg3��b�̯#����3Xǈ�s���ջ��+���@�N���3��� ����:�tx���	OO����=ٗB���"Bt6�N�\z��1#Yf��)C�J2f�x��qbr>k���n�ӲV�6V�z W��w`�
���|{_u-a8�0��r��V�����uYT�� (0����������C2X;��>�Z����c)���F��t�7�J�WVl:Ի\�Mm�%2�$�gC�b����ED���^�K��QJ٧L��D|A��_m��9�2�eֻ�l�!����7��:��
Ҭ�|���H��p�$ѳX���I����Q>&(�+CwOj^m5�[{]/2t�P�;va#k6|L���DTxu��Oh���V*^�U(
��MI��G�ķ���7v~�����up\�M��V�3�>A좡��O��S��_mԺ��]Ȳq��M�ʑ��,}`�Q��\Zi���^�������d��:I7w��0����Y����˔���]x�T�%�,��	i�N�_Z68�k�)	ߧ}���vm�cB�#V���0�!y����6�g�f��^]5y3XO#5�q�e�2�\��F&)O�],f����p�=7Em�֭P�{H�ŵɣ���<n���&�'�56i��Fր�E\��ʶY���R[B�C������p:����#.�]�]����N^�����,k*MA+q��H;�6���`�KN@y�]�\��ш�v���=�)�mnEo2#��:ɾ�w(��� V
�S��\zƙ|N�r�=��a�nP�9�"��Vؙ�)4jrl���肤��]Y+ ҵ�\�r�u�j
L�vj�o%��fk9P�媆�K��V�w9���d��=K2@��H� ��*�����^��i]����˴M�[���<�	���Y�M۳8��0t�����.R�wy�w�G#���V�4����SC�/��kU�^	z�
V�������W��vLT�:�>���T3��T9�Ǣ$��q�iǢ�1�#���T{{Y��\��mN��c�,�Ս�[D�X�_�jNt�rM��w[(��@5VH^��G�ە��s0s8�^Q���X�P����(F��\�����u���ڂ�N��_c��]�7�_u%;�5�C;�2��-0P��V�(j�z�+(���V��ܭ��v4�<����u9L�g����a���ug��]6[E�L�;	=}y�*�d�uh����n�V��k�c7�i�Ћ�3��<Tf��n�l	�W</e�3kR1qɝk�#|�Qǅ|q{腄G�WY���/Y���|���&M��a��ս���}2��;���6����b�B�ϱ�iPe�޽��Z4�[.�EE{*䪞KM\s%�5h�S
���=3k�=�d[�lrܨ�cU4카�V�2�]�h��V;��RuE%*yĮ��r�V��-���-�K�&��m�4fr{yҧ!k{�ص.Ѐa�T)�)=
`�0qMi���[�=sD�6�A	 F���P�9<$�8D�G�G"
��bj�&���'D�JU�L�GB��.�L�E&��*j�����+�$�dr�.wP�
����D�����I���ˊ��ɥ��绹T�'(�=��9PEV��.\�ADQ�
(�)΄QS�d�!\U�DK����dp.�W
�0*tIΐ��J�WNb��GvP�$�-IS���P���N9)���I�!	'q
��K��jA����-Z�:z���u�@r��R��s��Yt�*9Q�#�
��
�!EԮUA]#<3����g�j.��3*�<�0�Ȯ���Tps�ʲE�՝0��G#2]i��9\�EW<�;�ēw���t�Ӽs;����N�-h��6�8�� ��e N>���c�1�����CC*�;w�cJa�ߢ>���;�s�bt�LU���ؓ8�7ظ����X
�{j��ۣ���S6{�l���R���	��D�b�pW6-սNp��[C�U9d�d/ڨ�%m�y���c�+5ļ�p'�+��&!c�J����<�搁o�&Ԟᨚ���NZ�Xʸ��F��P���J�cb�s{��5n����kSaT�����L�l����<�GK+z䥪Wo-�o}�R���а���f�'w*;�][;����
<����!�ԝ���өP^��0Np��s�o:�z�@USh'��c���m�J�P���|T��RI�OA��p���/Q�z���9}�k]��:�-���(�����!��v�'o�3�
v9IR˳"Ψ���ܴ��y�'�*�NY@.X���3t����wpr�X��Wt�|�,UxeBM+�_p0�F���/�j<��
��^�<ܮ�}��r�[�Yz��qUTw�!)�`�
��P��6�����3 � j�q�s�fMզ��#��C�v��m̂�8��u�U�^�띤�jܶ��JT]�B��فA�w�"����ouL�5��
ُG��F�<���]ܕC=u
�5˶�;�|�oܹ�m�u[�p��K�b`�%�T���≮cd��߲#�_����}��y��{gk��-QH����}��p����E,A��M!Z��D�<^����;~������uj�u؜3��v������ш{j�}��:�7���F�M���O��t����^{�����){x�����Te��;7Q�fn�oB��N�on\ډ�s7�qV���TLV4�x�x���?��\B�̉r�ڲ�e5bO6�e}nGs�쭸��W��,i��W6-ս�E��g+恬��"z��齳�H<��Aީ�F��5p5¡���P�Q�fcf�����˸��?A^��z��.�s���g��Za�h�Oc��n�V�8�S����7��i�ä����m��@l��T=�*5W���ٶu�Wbn/`�'o��0JW-F��5�ǫ��b����οj�
~|6��*P�����ٛ�w�!9�ۇ:�Y�*��TK�7283�A0�k#�.�2vs�;4�+a�sS�WM|��ܱ���E�'I�����;5��_UUU1����~�蜢���ӥS_.om�k.1��M=�^�A�U[�6/^y�K���^�;2[紡���	�!�t�j��ֵٮ3�-��R��������e%�bW�l��h��|r���9}�[���GP�]|�|G�N�|lE���M�^Ud��G��aq;2y���Z�˨�=��9�m5�� *{X{��y�D.��hҞ���3Gy�jb+hD�^�t��f�U��5��<aڸ*Q<��@<�\��;è��yٝ^p'o�������k5	&|ۍw�:艎Cg�kmޖ�]�\ԭGA�2+Ǵ��QQu)�\G'F�8F�6v��~�dm��+��s��A7��̵s�Z�ə������oj���5/o�NV���l�WU�F�f�Lң�Ti�h��[u1o���5<�\�	����EW^��X\�_��vs�T�9�6� �W1�)�+���=3 ��d�;�܈�@��vH�q��/-�k��'�_��I�iCW�"i܄�6GI����#��u�L p��|�l=�[D��6�����s��Ω32p��B�A�)>��݈��t��G�Dt�=�Tܢ�WV�7��y=�n��2���`{79�'�;�-I��vS�z�R�%|u*�j��m��V��]��<�d���^'�j�.�j+�WQ��!]�F�c�P��%͋�I����W��r��V�n�=0�z�+�Wn\��(�=�kyp�}:��kg��<�%8�G�&ز>�8pVL�N�q�eWʕ+��[��\c��	����R�*�
ۀ�W*��=�0����J��u��Ӕ�����2/����㡒���n����Y�%m����b���g\*}.�I��-H�z��f�WH�3��Bq�Qm��(�"��pb�)h��ɧ+�0g��T��⌑��;�ZV�kY�
�62�r��!u@��hN3�Dբc�+���_t����2V���Q����0�(V�8wY�ٕ�Z?}5��]�s�+�ӷ)JZ����B��n�:��~Ѿ�e{|���r�>}��	�+_�՘\��u�Q˝H���b
�4���G�Ƥ2$Qk�I-�$f��L��3U5M�t����M.Fئ�1p��j��8�Tѫ��(��@��&�}_}_h�Ug��L̯�=�5o�������4�N�I�a��jĹ<��LH,w'�=yVC��[y����#K��EE�T~>ONΡ3w�s�Д������u�u��Y�؋��ڼ��T~�����r�ӡL�B�K��z\4FU=}���v���j;�/�#?Y3��#��������3%v�{��*�d������kz�$޳�J7ϔ��[*f�^�}����k����W6.[ۄ�v�mm=NY4���9C�O&��a���++o�*��'叙�\طI��UP$���0Y�j�����8�0{��PU���:��\��Q���g7��C#�n:�I��0eq��b��5�;.����:�o��ܝU&γ�^>��ٯ*�º�R�݄'���c�5�P(t�܀о|�$�-��Z����,����f[��j���:�ngCK]�u��;v��5���- ��b ��j�X���d%�|�
��q��Cl%B7.��R�H��w��;�3N+�tnT�"����憁6GI��������zI�U��e�:i��.�./�e���P��FNO�U��o_�7/Y�;>������5���}o��KA��6;d&;���f�����y^#�&�1�:/i?���/����kZ�q�o�{d���mxΣ���C���K�@�@O�d�K_m�9i1z�=���P���Q]O�rӫ�I�!t�	kf�W=�|��RM+�_p1�.;JB��/c�f��Ns!�a�c��c"��k�p���Z�q�7$��df.�Us������p�B�L�!�����E�=���R���cL���w]��E�bݒ��`�ɸ�j�c]�<�툺��uji^�|�9�̞F�/1E<3�M�mk�W�u�pʿ��ڇs8��F �Z�s]m����M�w^��1V0�9�x�ncn���R���OZ��z��yٺE���N9
sm�	8;�3D����^���TLV4���9	�V�n��_,N��,I0�-_W��^�-��/n[X���ǻK��\��l���Z)�weC7QI�g��I�	X�>��]H�N�VqF/ň��M������^S�3��h�A��S�L �ֺ�Ę��ƴ]���A�&5
�-����������ޠW�ۯ5��������\�{+nJaX�f��͊����x�Tn:������І�����'ڽ��.��-z�b�tV���2��ͤ�
���Or���f���9���[�V:����G9C��ի}ʱ��2���JƦ*��4��yƶc���t�[U����L�ŝ�BG�A��B}.Q�weT*U4���|�p�4���^�}m�V���ݫSe�ԫ8e�����4o��[%��w�ֵ���Ϋ|2pTNȔz_�=�6�͔���>+�F�V�Υ�����gkzp����]���% NX-Ög�B����*+����_D�9Q{:���<���ξS���|q�,jo!�9�!t����jt��2_��Ӱ�&XJ��5���x��D5��o�����E��L�Gn�֎����t�+��w���]]A�c���e����19�m�p�P6+i[G������.I��Ը��a��/4�i
���V����F�R4$���"Tvu�o�2�iwEMړ��a.�d�ػz�L�4:�+#pi�kG5��u�A� ��^�>���j�I��
��Kǵ}�j!s�O���=�n5ڸ?k�9�2���Ǯ����X��z�U2�aĲ�5mj�W�Ѵ�M���9UYЗf>w(�lp27/�hy&un�Ek�Ч���CR��8ewT�VdLS��;�r�0Ϡ�L`2��u�;ty����S҂���KU{�'�o���*"ꬽz�Roc���y�c2���M�g�'�9T���!d��Y�}���p�y��4�P�ޏ�z6)��=T�d�dW��s��V�ں���]<�����]�J1��?zǺy���=�!��_�xNՠfWg^m]��)�/�:r6��r�ca`n�O�������B���[�̾��q�׽:L��w���M��J�sx�7k=}�'m�!�+bq�f�ͯ���+��."u%p���t�YN��utr%��U�B\#�笥�N�8j�۝)�TOet���J9�{GT�m����M��ˤ2*�����so[4��h�t��ݛ6��[ /}jo�Սt�6��_KR\+���Ņ��t��/���w�vF��!�@I��ݢ�m~�� �ok�[� Vj�������P(t��>��I���\]����n���|��ӟP���T�}�	�u[c*!�3�!O}�%�R�X����r��uw��ET�c���v��P�kY�
M��r��!t�&�s�&:w{2�9A����R��u���\ղ�;���2�Rn��Q���yf�os��8(Ugw��쭎�� �>��a��q�0^�o���������{ꏲ���U�.ȉ��qP��|*Tf���Bؒ�mi�8\'����^o��_Y�y!�?CI�&�����"���yz�KW���^�+�b���P`2�]�gn��o	���=�eq�՟'P�=�w�s��&���>sϱ&��R����G��q�%G/g;m��f��	�qڢb�󲹱:���u�q��n�3�3M.Dn�Ӕ�C2���H@�;��]D���\o�f�����,�h���9��d�&���\�B7^�P��/�D+�R�7]��EI�w����'y����'0jNf�������8zj9t�,a��`?4*j��L�/62x��:�wn�)�}}7o#HH[d��.v}=��\5�J��ܮl\:O�!Wn�v^��s�m_)]�r��jv�42ut�� ګ�:uѭ�	F�]1�K9�������¬�Ν���]9����Gm�������ʧe��Jߖ�Bp.	�3ۋ2�+t�SNX�=P�>�[�(w 7
�����Gu�F�{�����u�>O_�}���i(���|�`���FO��,M6#	�I�����d����X�>��/��kW��:���W�R�>��b[F��J��������I\+�_m�9i1z�>�Qm��*M&���ףM�Uv\2|�@�O-���j*'g�����w���--1�ޤb�٪oZ���ˉu�c�s���_�����7=>�˧�V�x�B��=Δ�jFQ{ɇ�>�p~R��6q�ǲӏ}��E�S���\7�gT��G���*)uu�����k1R�8�f�(����Y�{ƒ�h��4˒�ht��ur�V.�[|B)eδ9l�;�cB�W(^��&)��:�����av^��4���g�mN�QFD�%�gr����� ��jm�
dXu"w:��fnc����&=`�17��ciuˣ��IR��ۈg�����M�O����|uR<��E��4�_7��v��\��u�[�u���)�j�- R�!7F�[V't��v*�6�o^=���"+	=Ɗ��jc[���o{� Y���ѓm�� ����}�Iv��� ���UeS�7��--��f��v8%�K���jˮ�B�+fA��ΊW_8'���8Ŏɛ���x��B��P4d���b��+�ݳ&���9���6���Ӣ96پ�`7�&_�մ_���D�����
ud,w���kH�!���%ͺ������\�j��*��av�n����˕3��qn�
�ņ%WC����Ӕ�[����gl�F��<nv��R����9�*ZU�Gn����c��!�3���e���Vm�gʒ̃uL]��J^ռC;v����s�1�0�%5�|�)�༬5Z�"���Wk(�=��{�:�\7�R����v���[��B��l�v�����q�4����\���pSy�+�(n�3��^�h6�����\͓�Z���+��z�d8UoU��Q�L����%�:�+�N��w��b�)1�92��BK�)t�4;qr��\_,H��ݘx��6�;p7z�#��s�F�$-e���p��ɼ�غ���C��'4�E�������z���Z�ݾZ1��� ��K(��7[0Z�z�-T�bʵ��hݯ-k��:{�uv�[��%�t^�T[b�_���o*6��&���Ҹ8�mso"�j��.�ګ|�sK0)����[j=�.W��f�Z2�鼨h�e����E�a���hcs��t���m���g�%َ:	H�^�,-ٸ����ȹ3r�pB]��n�z��:�rl	9D�e1�DE�Z�����c���Q���T�>'ԣ���B��W�+Fp��5oS|8�GU-�I�*����^�0ٺ�>fB����2A�dr�ZC�� ��X�x�>�\E�#����)����R����t	�`Ρ9�A��Y���ݙ(}�I�%-Rs�a&��И���ޏV����s��2�p��
�A"��C�/��}VM<�R�z�_Xy�����r�������z�4��+glət���G�WN��r�qC��+�<�`�K�V>�٪��p.�Wc�Y�5A)��;��7�K8����AyucOK>Yzq<��D�s�y�!���k�K@f�z����n�Q�Ԓ�륻Ƭ��..ޚ���Db�+�{^!��
;rHE�#��_�h�;��gΞFiG��Rbj��]m���ט�$� ��H0A �r�����B=J��+*$�AIj�QABq.�Z�*%W�:eաV�L9��E�*�Qh��'wj�4YG"���Ws��)�jЋ����^�Q�!S0�],+��Y�S(��Eh��)R�y�"-@��!E9��S�r*��,�R��;��䩥A�*<���*
�vh����<��B+�ˎ`�^e�GS���ª"��]��B)��.Y��:��V��9Ȫ(wA�$�仮��Q
,�t���e�B�'
�NPNβTe$Y[UG�(���9S�	1Q:�eI��f���D�A�#� ��z����L��3s"��VE�b�Q�B��K�mK�2���KC��r<P��'#�nN&�9E�W=�@"/<��'
�*+u���N^g(������L�*	��I
	D�%	��l������M}�����A�`�3�^���R>^77����!٢�X�K��qݺ7z�V���z���}�|{|�>�C"�?|�q[j�DZL��k�u1�ȞC�Zڀ�Wu�m��-��q�nGs�[�KM����\����8g�=���qY�A��<7Cr���7&����Oer^��H�_��TT����M�yz��}DnzE3�R�>�{P��L��1,l�H�U6��qڢb��pT�g>OZY[�����TVR���.��;vn��̯����T�V�D�±�&>X�; Fζ���Oet�Zʭ�Ku���z�_�dx�V�vr�^��V}}�md�՛{ֻ�	�Lfh����!�j�v���9(����5M[ �Z��2�T��Ƥd��g^�]���<妟[��N�ݶz��iN�ZTڲ:z�h�t���lՌ02t�����yߡ���Ol�X��ٌ����ϣ��X�@c*\�@ԕ�h�/ga�dW��ez�uƮƁW�_���*��L��<�d�mu�:��0Q�¥r�Y��V�Uj^��½%o�
�����.�W�����F�!�]SDg`���k�Ņ+.8�}���Z?L�YC��l�dT���Wz�Q]Ë򲛞�hxD3�1����^��|3GZ8��"�����C�#�]0W�h���K_M9}�f�(�JK�U��ӄ��	��l[(���(b�V��~2��u>��7��w8�$.��ꋑ��ɋ���*y����.�T0���Vw&6�7�K��Ó//�s����k���;W�R���V���׉�jo�	������5ù�.a�B}F�$�m�>W]yJ��Uey���x����U�m�kO��Qյ��_'F�8E6s9\.��;��r�u7�~R��b.��}[�$}�?CI�w�p���%ض;.��g�0�o}\�/y��ī=_T&�����h����-�@N��Ժ�:[��pz{���j�W���#u�fTq�Y���V�?i�k�ȹ���s���D^�x�a��&�����k��iѾ��̢���$�$�8����mk5��D�}�W��'5�`lV>���+�w�ĭJ��P����a�Ϝ`���S�NQ�,o-��䣐�r��2���JR��B;>��9Y��m����w�b"�yR�_b�=��R�#/�pR�ۺ��W9�jVk�^S�=	\j1��5́�c��!P0�.�t�ƼnÕw�c,L���_F҄�k�c�7��|瞅�����r�����[~ݞ�d��v���pjמ02uT�J9��z�=6�f�;o)���+�Q�d�v��Y�N��'d&=�TN6�<�ܽ�Xލ��c��&@ʭ�WֱU?��������)T@�����
!&*ԓo��Ľ�B�}�C����&��_s�;�N3��NQ���;���Yʮޛ�s(Ҷ\ʐ����f�%-+g5��=�_&�T9e ��A0[1=.�C�%EwMO>{�"�c�sI�����
��PvFj��Q2j�7V�^#r��go�7"��V��
�Ө|��O��I��;��02:7/���P�����Y��wY���c����Ί��?oN�z"T��>�a �o�(f.���s4�e����>�wZO0%ޡ�Y�M=�}�?�f�"��h���Ug�P�Q��[����+n�
�et��zۂ���a�Z$a�TԲn��҉$�7k06��ᥱ8;pǇ)`Uk�vL�����J�m*����De���n5���c]��vD[P2��u�\��W9!�|Z]��_i�V��u�'�y:�J������vػ�k������0���n���j�p�1���u{\�����Z}'.�]�{;�V#Ɍ�3ڥ=m�'������U^�h5+x��d��Y��|��$�i��V�󹾶���݉4���W;�Oem�	P�c�X���W6��)�6wژ)ls�d�W�ڛ�9T��*��uWӮ�F҄�ᮔca�
��ڷ3�;9�έ\�sW��C}].���[��[��7%��M���c��0__j����xJ���>�>˅Y�h�d��L#��we,��up[q5e*�Hr�i���T:u4�=�|یp��,�@����*�s��ʮ}���iC�y��'���X�>�_^�Z�dF�ζ�딺2ݫǳ�,Q�"r�%�~�=e�Z4��\���ڝ��n�o�y�qx��QZe�P�b<�	굘��9�=i�x�Ѧ/C]��W�QB��.����|ڲ�a�_o��*��{�ة4�#ݽ=�8������L=~t��x�r/��ʵ-�\�L������w�语?BnQ_mÖ������D�E��ܗ�-`ݿ,֫��)��A���jT~F��;=RzM�����	}�!�5��)+��H���@�P4���\k���Νm��*r�`����=�4���7�FB�L� �A��":����P���{]>��be�x�5F��`�ɸ�p���vD�!����8y�BUq*Pd{"�o����W�/p��=�U��A^[���t��t6X��c�9%5�a�*�GBco*/�Y8��������>r����=<�.s8SÚiQ���n����03L�ے�m����al��9C^)�:��nQ������ӣZ���A����$��p�D�(�7t�ʷzu:�j���ظuoy�ݬ��9T�ʂ�A�:䘍���Z�����������ce�������u���%츔�s��]QB؎m[[�]����`�{9>�A�������������(sm��4��:�o9(�����]�,B��+Ej�3�u�c͜&R�q����ʺ�d�M��[15X�(�Yb���U�\��;M\y�d�MUS!�T�_�Gq�T�sYw���_;�vQ��tK](�ðմ��I�َ�<�ɢ�s_l45�p������.�ʨT�is{o�Yx��i����0(_;�����u�Z����Q葯t%A�w3CRV���t�i����˾��|׆X�Ȼ�O8Jn�2\E�NR�AO���*KE@�k2ΨZ�LB�� �5���V���8��Do~�,��^m[_6*�^cj��p�Ŗ:�?)���ٻn2/m��F�6ҿ�����	���t̢P�������
���r+:9�J�+VcE��1�چ�����}
�O!���j���%��Y���7g�����#\������tk����\S�.k*�.�TI�p�����ǗU��g�"��.E�p�������{�i�T�f�_R�dW@9S'���@�}]494�����N�#G{��qGλ�#끺{)�\�xgN��?��\�yKV[�z�Z�0�0�m�.�V��qЭ��r�؍�ơ�O�&��îP=��5u�Z陦�h�t�	�e���{�^����8yo�Rvܬ��S�e�>��"�Z��}�s˚Ϸ��׵nK�+E��yUӌ8H��q�Wl�D;��vn��Άb���}bV�ZХ�ʙ�O,}�j�h�	�V��^w���3(���;��"1���z4{ʶ����*&>qe&�ë{i���vr���۝�5�\!>��J���9
��^�\(��k��>�U۷
� ��u���ͷO2��f�p�E\���geB�]+�X�m>3����u�<��D.�)]��l�m�QL�)�<�"vx��+aR���ˢ.ђ����u��r� �n9���΃[�(t��
�(:��Y�8��#�w������-���R��n\6یp����)WL}�>
*L\N*�;5Y��j�$�Em&�g9}<��\3��!8Ψ��2�n��w3���Y���xH��o}m�бŊ;�2;�;�t��n���|�p���f�aX�hl毣�ח��Wiـ+�����\r
�I8�rv NeܣweI�[�X���5ҵ�'pm�)̻�Q9�j�>��u�6%l�'"�i���`�pYql�U�\�>:�ov�)i1z��=�P�P�:���IT��������,RbWP@��j'�=A����C\��/���Tc9��r�ꨞ�ᆟ9�qӆ&-����\����� ��0P�Ш%h�6眄H�ƻ�pS�6����u�\D���QQ
��§��ЧI��v�E�[}�jۆk��kU9�e�[6"������F�K������ޙ�^�5��W�zw�8e_�l�D;�Tj�0-p���6fjs9�aţj	S��"���	{�?�o�5=���p��3�͞�=�p�b�!���HR��t$���n�"�޴����1z\��Nd>��1�:\��Z<�e6�i�̌���܇ʾ��ہ*��V>f�sa�7�uv���y�>��\u�w�$�$��H>�*��S��ʄ�>�b�o6s&�$i���4b��鎕^2�V%[ʳ,V�=�z���<��N`���y�b��w!�H�5��JJ�T���j�Ӽ��/jT9[�0Dg6�;��Y�(��֫�B�W����P�I��u��j2f�n��l�!3�ƴ} yW�~�?O#�=����g*�'��<�'e��6վ?1fK�ۤ�Ȫ2��(��z��}p�=�[��܀܂�]�Y3ؕ�Uu����r�ȇt]|���>On������-�ID��[���d��q9�w89�4n��#c�O��׭k]��3�-���b��z��V��1��:��@��~�0P?�W�y�����·-+g5��-ڦ�q,�v���8��9�!uJ4T{5:��|*��2݁S��zQ<���ڗ�Eθ�w�\J�g�⋫�:�^d^��\k�Y�������<�]Sh\U[�{�j>k�m�h7�B(��CfN:�_EUc��ܜ�M��*e�ǳq���s�i�5��7�Nk�6��Q�^�=��X�Mbz�=�%�������_']q��*�{'i��v�,��(��Y�mnb���B	��m�bU`U����nr=�0#�\LeġFw�j�
����a���O!�죙6cP+%����l�N����uN'�]g�����:e�M�,�X���.�8h.���-��)��z�MT��m��N�����[UcϬ�v��;b���xW��
3Խ+�}C7X��4�0�QͣW���yL�S6�܊Ц�o�}<�p��0+�桾=ϽuV^�jڭ��ٷf��C2����#Y�7'�����䥩�1�goz!�>7��n���]�׳�rPw�U���5�`�|)����\���ç��l%��v���v���9T�ݥǤ�6C5��|�/�T�O.6�Z�p��C��_К|�<�Z��\O3 �<_����r��?V�y�L�S�M.om�k/=�H({.�E)N+1Fi�}P(9�L�s7RKd�/%Vb��\�6;ecgN�S�J� 6V��:�-p�R؁AO�����1-�&�g����{��{�ӟP�r��p�h�Ų��
{䡊���l�;/��z�]KƆ��B�\�s����7,5`��Y��a&<�ҩw_n>���S\�c�w�yp=���<�u�м�H����^��P��z5�I�}W��N�]�"��-�F�J�ҡ)fXx�Z�	�.�#��Μ��%�35�Wf��e�+���K�d�L'}�1��b7�gJ����`"G�n^v�#cdZ��i;��dUwٴ�`��9p����L�-��=�/[<��۱��+O?_i����+�<��L(#k�8j<�*R�:-�:
ȷ�Y�������|� �3ihK�k�e�u	���kzf"�k�1��u.�"���8�bA�1�o�e��d�H����X�M̏fϭG|��	QLw��d��<�gv��2�,!���u��V
'E�_\V�V35�s�V�4��+ug34�w7�Uh �����Q:�'F;9���{/��ܷ�ɵ�"�[eios��j��6N{Nn>�+_&[��y�G���x�o;#:
��Fs\�h���W����ѶP�Vr�n����f�ӹ�ͻ�1��T�ni������j�t*�"�+�6�62�y�$��
'^Ӵ�"a͔rndb�N��x�eÀRY}�@von�\kNM��j�^@ogr�Df��ܬre`��(6��J4��[�m#Pں٘��	0S�%��LQ�8�΁'�9na4rT�(��6�қ����0bP�Zh��\��JA
�rc��9p�бr�:-<k�@/iY�Y(q�5�Xo�b��K٫,׻C&��,�#����
b�!��΁�����v�%��a����^˫�+l�����R�>rM��k_;��\:f��W.��M�b����G��)��uD�!�S,��Y�ý�]P᫗*�n�f�/DC�2�ҾG�A�ja
�Ws-WdD�V;Sm�ou�-�	Ԃ�ޕ|�ᕰr�^=�|v�]b�Ћ��u�KtՍ�,&�,�lZ�Vf�LZ 0U��y��;�-r�3c��l�鮯΢�
��(�<�w�J/���t�c�=�;����]Z��Ǝ���6�X�6ν��\��>�$���.�z{#�O:kc7{�pQ`�U���K�(����ӫ�}~��d�?u$R����{í-F�����ά��8vZl��W��hy�D�N$.9n��\�}%���8_'R�}�-�{����;G�eY�mAʄe�����L����x��WX�֜Df�m��x�B�h��;�%�fv��F�*��5.u�G��Z�-�8vѫ!�uü��4ՖV�J�[9v���qR�*�B��l�#���T���]�cZ��h�E�2�[�@D^F�ti�D��w����\��c��	aa[�l:uy7;��%6C&�YOm�F�6��xp)�Y
O�և�v�Ǩ+]�G9��"�r�G��U
�M +J�S�2�Ă�p�Z�A�$�Q�A	R<�eTur)<�D´u,��]q�z�;��QȈ�M�N�$�#@��R*������c���9e,��s3�k-I��r0�#��K��<��eP��ۈh�Q�
�]w'"�����v���⚜����b�3L*"3
��Đ����I�k��9�<2c��#���U�z�,�R�M��*I��f��T�G*'\���U�V���2���<�L3ڒ����\����L�@ڜ�$����f��(�9:�^m(�l-J��Qe+S8a�,%�{r��և��:UqȒ�C�3NU$�F��j��z��{�I�y�eY��"��Yz.Ay9�s39�ͦNVt���疴�\�ݪ�%)Î"�73��*��㻮�0�bH�����e�"�$,���.�P�:��"���6�p�gpܡ�w���N��oэh��M˔�ڃ� �������3% z��$�a�|u�r���[٪ۈ�%G1�wB�(U��W淁�
M�WΙ@.�) �F��Z�ؗQ����MJ���ݽ8��k���j��G�ZM)˩�̞�\�� N �P����m��r΅�:�>�I&n1������oj1��z���q�$8�6~��+����8�WFj�SK��vw�R'Cu��R/�� c��yV.cL�/��]�����+\~�����x�խ�(��+�����ZQnW��;N�uٺ�C&󡘉��WPVu��`7+�#�՘�yQ�s�#����pT�g֚�{��#Y�fTAv=�F���;o)Ӟō-	�?n��cv���z��Rl_έ��:����]]3�v�72��! ��=��[q��F8Qm�sa�{ʻuU�]v�J���[����!��\}Y��Z�ƶ�%�p��B��@�̠%�J��,�7�V)-[��Ֆyg�]�����3{"oe��J;��L�R΢71�V4C\��/�B��mY%��\�`oz;��\�L� z���gFA"���N���u��K��9��;)�L)]�+�[9��ށ�;�T�f�+T;�J�ʵp����06`�?ʧg���*�R��Ã�I���No{���떂����/=���5�_
<����0(��IN�j�P��S��ǯ���O�Y�P�<��[�S�iJU(t�|�(��fe���4�r�ips*D,�c���S鯜��gnBq�Q��r���[��m�-��V�\!��t)!_if|r��E�?��k =�P�*����{H�Xjf�7������
YA<�j'�=�����+湫e�cm�t�wr�=ɚoR��?��b����t6�s_M�ڸ�N� �;�b���mv�ɭ�H�R2��L;ƵP���9ko"�pȉi~\�笟sP�Y�Zc�N%{K�TdM�{��Rz"ӆSp|����,?[ڱY��V�~�&֎#T��5�b�q�ky�ܫ�I�\bpʟ{!��gC�|='�As0{��7x!]�s[s��(˘�F�����=�N�[�����c����Wp�8u���0�>k,��h㓌�w�'e����VVx���Q�8�;���k6x쵞��b��;0�w<�oG�d4�f��ލe݊so%̙Q%�8뫚S��w7��cg3=V$��ȧ�v�S�k��&��Sڽ�}��%�Q�X�%m(����r�'\=�w�f:�����m�ڢ��lc�}�:�:5�=�*'2��t����9d���|�d�����03���y�{|��\�w9_�r�9� Av���삭AZ��˥INh�fL|%��+�y�7xS�or!�j�sۃ[=�r����8G�2�4>{�U�g�w�yM�|���O���sxP�@m�W�U�']���҇�jT�J��.e�>On���{_[��ׅ���aK���n_[���.F�jJ�c�O���쿽�+�Z�R�r`^A���5?aV\t��Aw���@%���Y�uB��nZR����L��S�r�����h����Y@+�J4TA�Q:��+F��3���f�q�Κ�5�/��	4�Q�V�%mR�g_g��㞯J
�p�s�@�k�ֹ����l�-�N��뼓J5p��ڇ�{��F%�+9Ej����cj7wa��-rj;Q]��V�A$�zn�ay��*W4�$�o>��f�R�54IE'>�GL\�W�͗��x�U
��⋠R��/l���Z�_"x��S�8�M��_G.f�|7�\R��Cg�{k�۵4��|��аǶ/V7�F���.x�Tm&
j1?���Y=7G���@�o�<�*�����M,^~�����u׉�/�OcqЋ쉬�؂9�� ��Rv��G�dΪ��#\v��Ow�p�M�J����C9�r������3��[�c��]����uIOa�;j�]����7}���J���E<|ޓ�[C�W�Y=�o��:��TM]�s��w�)��/By��k���&J�įp�~�:ao�;/��A������<��s:Ԭ�򋞄�kU1�P�7�^��{����m��7�z����:�n���5�������lW�yq	��Sɭb�<pK���3����>���6���:���ܷx�S��{+�h�;k���B��jfv�p~'�V��/ǭ�V���B-S�&�����mM��^��+��7�.&h���0&�f�� �P×a8��j����S�� ��\��U9�]�[��Ծ-:��������N�*�\��σYo�|�N��W6��d�z���T(t�������+�mN���(��d<6]�w����4�G��E(��稣-7�͗d���s��m����FH�=ޖ_w3��=��m���(�"�|�0�\�!�;��Ѥ��"v���ڄ�W�9����
��EC�e�k>�˜+�pr�[fJq�=�5Ϸs�x����6�;j�=Jc����u۝-��o^d�݌�
ݠܧ�4&��^�ʇ�z��@6�:������9�K Χ�L��FS}��ֶ�]W�dd��<�U)�m��ZeU�r⥠���E�p�6�}Li��>2��"�_n��q��9~��Za�Y�-��^b����M��e\=���g]��C&�bRD�ͰW�T���H�܅���P�Bs�ʠ�Y�Λ4����f϶
��ӻ����5���1�w�g�.�#wʂ���(c��3)ms��T31�Jʭ{j9��mD/L���ul����������فI�RT 2�atڗ�6fWo]9�[�[��A����us�Vjj�K.lj���o[���vT�e<|��9Q��������ff�G�H�\g%b��Jm8�Q7Y!݅D�|�M����Bk����v�ˑ/+��Žr��E�	?��Um�P���
�6+湱p�>���>�puN���m�\*��^�׶r��>��������t� c`Wet�5a7�G��v�H�ǹ������WK�sª��կ<+�j�a�ēebu��
�N�e��7��8{P�{pkz�:c�0T� r篾R��i���Z��*=�{;S�h5��շg��'}}oi����g����{=䁮[J��A>W���>�r���ې�gU�1�x�VwR���'ۆ�7���x֊������ovږ����<���U�;�O�N�G��s9YXs�K-��j��y���簛X��5���x�]�,nW��鹽G���Tf�ݾO�F�X�e	�<�w�K��^s��.�T=�Y�[w������=[B�n�%+�#�x6h^��5=��U��;��1�&<x�XLlEk<u�YA�qz�^%�fE�c�>��S:�q�n�q%�!��0�P|ؓ�F&�$k�󃿝��(�!��<�ܕ�jDk�s���Íc�]��>�o��c��h�I�a��p�BtD�!�
ڈ�"$��[~��r�i�;eD�zO{�.PNq�+��K �^z�oj�F�S�V�[Y1����[N%�ۈ�NCT��R<����{���T��.�R�6��	�W=i.�_V�d}O��������/9�|���tƃ}37�l{4� ��5=��c��v�����w�ZJ��똽-}P��׼y�7{�<��u���������`R�5�m�;Y�*����A�|}0O<Ow���=T3�l\C���Wnڽ���� ������]g^3� ��b�<�1<�u+�&)g7��5n�����@l�m���r�ΠN�귖�R�q.Q�\U-T�[�z�Ɵ_Γ�5�B�fRt���w]�B�S*�@5{���^�l���W��*m�y���^��xM<�T�n�*�:���b��20ؾ�F�p�,�e�:�|_gnEb;��6�׻g�Sdܣ�T��oSt�Paҕ��)����n�_
Z��x�#��-�
�8��M)>�]P���ϓۇ���zվ[w�f��eɔ[�t�)��
9���+��ljJ�V;t�k�/��ָ� �5��k/�5nA����2��B����b█�j�,寱ͺ�Zy�o��XsD�e���jǼ-�R!OBS��O=����D���܁��n3=��N.��}�+��L>D�W�\)F�����&DZ -��WIH�Оĩ��e5���6�s4���q����(����=<v�zu�b�L)�f�U�t���-�����֓�Mƻ�u���[��ô-n�7˲�_��C��[E}Z����^މ�wbp�
��(�u"���떵R����ޣ�V#�&w۾$}Z�>��������{����Re��8�H|�|F�?FY=�?o�d����ȭi������M�h���!ⵆ�1� R���-�:%���G�v��*fވŎ��]����H;6�jPD'�L��质�X�VW�c�bu�=��ӃHC;�����&��e��ve�_v��t��`��{�V�ӊ�C-�����U���D7�3 �8���2��s��ݸ�ٷf�̨*���0�V�[p��)=/v�F �@�f��͇4�y���ٽ��H<��1q���V�8�{.��X�p�����m(j5�ؤ��t�']�n�z7���֢*� �m�̻��Y��9��0����PUB�Jƶ*��4���aؗ��`��(�3Y?n�UHs�9�z02M��?y-u��c�8P�YN�'� ��ͧ�_�C�%GĔ8R�I[->���>t��^Y��ں�5�G�o��{�^elw�F�3ʈۇTø˚����X��p;����!ϫ�����)Un�؟k-x:�F��Wq���|Nx�)�Wg�dmǦ��s �Q
n|��eU]{���gb��=*�a�E��gQ�|�G\7�lǎu{�����p���.=7�"�%�B�L�w[e�:�o�W��+����S\DDZ42):\{Q�=q�W#��_����V|G���V}��Y*w�K]v�/%�wy�3�3�q9)C8-���¦l�����4�XwEaR����Z0��M�������q%.�̐���Yʕ���o�춮�x����1[^��A�gX�&��Uwlp5�C���%*�p�]�����)-�d��jV�o7ܥ�@򭩓������zĬ1Q/��n���iK��YʪD��.�x.#�wOs!��3���;���z�A�R������t�[�+e������ta��ɽ�����{	�`��J�M�@9�����,��*A������;�
�*�{����u��ջ�a�i�Z+O�o/�<꼎}����G�*'�#�t+��䜿�X:jJp�o��Us3��ឭ�^b�Y~��5+�������މs^��/�|S�ۏ�f�G�3�����hߔI�B�d����Ό��UVYѐi׊���`S�,���~#�Y����![12��g}v'7c/�bv=߿W���^ʟ�|N�c+�g�]���EK�<�mxp7��E��_��zB.�֜�nשP]͛�C���s犢���MŖO���xh�S�WUzOS�C�v!ť{*��Z�ת�+�^�h�����q�A���hx,���e��$�!���WM)><�����܀Sٷ|�ȫq4}�۸p��
�t�no�q���xq���l�JX%M}%���K����������y�me��Cp��X��J<�X;�8G�ЙX.Ё��@ת�I�yvTq�p�K���fR���rK�7q,���o0
���,!M��z����UƖT|�٧�(�v�����򅺆�MT�2���3�ǻE�fe�?#6��Z�{9�^d���/�K�I��s�'��=�c�j��j��X�v��^�7������+JP�F�&�ք��fv�r:�����n��v1]����e�b8��[n��i�R�	v�ݵ�Xr����l �T���ԑ���a�EУ�m�Ǽ�R�e�Eau���{(F�&��oy����C\^̶�&WɅY� {�^�B.�]���yiz�lP��Yhk$4YĀ���Y��ec��!�������<�u��t�{K-S�r�R]����؊�TM.�*6��K)��d|c=!�1?�$�d��Ϝ�2�ۥۮZ
�[b�f�-0ja��;��t%�O�[a��'�vJr��2��U�OՓt��o7)��nsu��Ss���\�׋x��Vv�r ����)Q�m)Pb�j���,vxMCw{��zj�V��t�$��T�\kza�R�R&��2R܉�g����93h�����x^�jQ�N�����:E5�|��Y;�E�\�����E���4
��(į*�;sE�8f�E-MX9�J֋�'T�4<�z���6��C֒K���3Az�����9����;4D�o]$��ؤ[4.���ͮ��x,�r���;�Uo϶��r K'-����W}�[g2�l{-j�BAWf��3L�fj�a�10[앛^j%��A��%��1����L�fa;���2Q�r�+x*8a�b�J�Z�1��!MYr^(]I��b]l=��y�Q��e����q ��Ol��t�&��JY��D�l�t����`檏.�� Sԋq��*Q_�v,���-3��'�+�+zQ�ͨ�[�}�cʅ���N���
�4=o�%M����6u���2.Y�|F1�^ZyXd�p��%�d9yy֎�Z�C9������s7:�Am�@s+yHiRWXv��I��7�T��n�ĩ������ ��r��)]XI��N��wZ<q^��!��3N$��bޡM����f����e�ԍ�K��6���Ih�[���r����\�C�dΜQ�v���8�T9*P��N�C���pa6���ي���g�ݷ7�-d��x��^�7$ްVh}nG��:M�':ALV�t=nL��vv������	�|������s��k \���@����-nE��V��ս����Q�:Z�(�4n�Of�E�A2�f�׶RjsVK�֣�Z)��������U���s������1�}�%+�� ��8#�Wv�Wpr���Z`�����pNl��^M�7�yB�V寇^�/FyN�ˠFP;��r�""���*�U���<f"F��@��@�*�$)Λ�x�{��&Dt�P��,���-l�����dPJ�H���9g�j樒Q�S+ΩFFaI(��O]�M�a�0E.�C��+����h^��(�3:烗G�SD�&2���*�V���J��(�V�3"��Ēʥ�V([�(� �Zf\���9$�OR�2������gN*/S�n�OrH�
"��a��9�ٞ��;��͐�Fa�LV��YqR"օ����]آ��H-,���
4E�TJ9��Xt�EsM�ENC�������4)�2�Ģ*",�
�d�Ur���3H0�#�0̭M��MdDV,M0wn[��.N��zH��\�P�0�n{�Ft�Eҥ6ig9V�s��eS��wI PP)PDW�V��ϵ�Tӗ��X��DٴlQq#E��rv51��'��wY�i\�nՅr��RA��o������1E��^�T�ݑ��}�>�Re���]O���Q^�^��,�>�H���+#n�.�B/r�#�&�����#�%���n�7��ƺ�EC�Rq�ZF3�N��~��^{�{��>�����o�S�2=��Q�@�TDL��H��:�;�΅o���>�^v�zw����H�yJ'a���rɪ]��G�%�ݰ�}="s��N�5#���Be�N��JZ>��:������r�O�l/}^�5�Y[��iH��D)u�}�ӣ��x������v����M{_�e;^��O�VP�������!�^���D��yUɸ��xG���u�?UH7�O K�<lL�ʓD5��9�<�G�
�a�W�x�����k�q��U%c��6����.�Gd�G�����T�.y���xͳ-�{��t���W5~g����yp���1���^��ݗ���=������wEb�m���I�,a;聒��:�UVx�ȅn�+;��^u���u���^�w��.{x]�ߪ�P�� G�Mz_�O}mY���9��ߟ�f�<9�|�.� W�W��C�k�iv�Õ0c<v��--��:�Qx���8���Zzce�n��O�����e.�K#O�*����y�׫�ؤ� ��ҜW��6P@
�B:�7x��Am�(����q��q�y�|��e�tZ�V�Z��4� V	���sV�|�L�W�T�=�z�w���Q�ʝ7�wA�dyL5Kn��EK�<��ob�\:e�{�7=�}`{w�$dEzW�'"=tǑȇj�vD<��t䝢��=�����T;�~�w��s����tr
��\�x��w��KҼ}�=�����W����p�ӒpJ�D��+QYH˻�������c���	ڎ��U�1ԦY�|���ޯi�t�iϷ��VG��{��k�7�X��	õ�S�]�߬}���	���,]u7���|}^��N�8dyS��>=�3j	��Lu���8�]�G�W�7�
�\� -2����F��������B�^W��%���53�ʷJ��� 7��y���y�\7�P�\�j�>&&[�$q^/Q��U�z*VS����ڊ�+�o+�.��=��ldzv�Ƿ��C��zHΈ�z�j�sP��ċ���*W�}����u��*w�j;S��]���j5�܅G\7�l��P>,�k���u�S�fQ.g�L�f��=�{/��ɍ��x�x�N]1W�#�r�x����G_ɫ����ȟ>��ϝ`i�ȵ�LFX���6c>�� ֊�5�;��F�:��j�]��^�m�9�޾�6�i���[{?s�;�s|��=�Yo�Zh��O[�m���vwn�躔-�뚠\Ѡu�<��w{\�gM���'�g;�.�3���e��L�ZrD܋,��V��ʕhLw�p֠s�cĹ��
�)�Q��h^_��k>J������w&/��/��7���e�{#����ی�zFu�}|}�2��5�Ī1�>������W:^7�����g���@0'}�]z��S�r�\p�L�!�xO)�#5�N����j��^�ӑI�do[��d�z��U�}�5R�0g�a��i��k��hOF��^��y��ݸ�0�k�P�"�/�l��9�ޘ����sw���%�Cj�����%�{}2�1�R���gep��NI˅,;L�5����A{����9�h��w�+�w�$�K*Ϡ=�IQ{œq��=���,�U�s���]W�&����(�؁�e�&|2�L��]J�b��C�p��;��7�����/��\wu*�7B4H�yz;��f=�����$�2��g�]U�7��K�ޚ7��G���W��[�&-����Ws���7�����R���'�� )c"��O�"eD��o,PҼ�md�	��Wz��W�>��F���[���9~�v.J4��*��8R�I��Ke�SWw�!�dgN�F�U�����~"�����7}�&�U�W^�G[ײ�t+��,9	ѼǍ+��Yϯlt�4f�Z%c�Ay<�H�Q�a����4f��yii��)p�C�w%�l�|�.c���CR�V]�J��=�Q.� ��{��9�ا�ub�����X�T\�M�z��*�^�i���<���g����p�5�<��$��I���*�^aL�P>���V��F��ʢ�>�������/�:
�z����3_9�Y�8F���e����Ǳ`���R��>G�X8�|�G\7�l�Gޝ�������p���3;O�Ѥ�nmh�}~�2=�>S�n�Q>�#B���q�e�^�\��5~����ƥ�93��e-����5�R��N��2��L�G��|&az��1Q/��n���iK��C�cXmP���p���T|���su�3~���|�0w�d�,��0��\�jsDV���켎�[��G����\�\dO�h�z�����\��~����	�Y4+^T�[,�@���ݨW��*�mA���j5lb�i���~>gyO��m��g�W������=�Q=���9l�t�ϣh������ڹ�w�?|2Xs9I�S�'�.��y֮=�潧�_����w��4���Ъ�7ӹ�3w&r��3FQ�rt�����G�g(��4��NF̰)�G�o��\G��ǌ����MG��L��W�˅��k������gB�k �5�70ٗ/�n���Y�5C�v�tP ؼ�{��������LP���.�}gJ�0���������=|�m<6/Y�~�ӵ(����.�s�pi�s8k�%���j�-֘���K�#]�=X�W���h���X����Wz��� y����7��AY����m��ϲ�-�p>�u�+��*��ӿYd�Y�xk�=LOL�N�[��6�3޺�v߻kTP��q��G��}��SY����Yu¾]�(ݖI�Q_�A�P�0���uN�xY�W���tNz�|�.'���C���{���s}`{����ó蛮
��U)`�;�
=�U��^=�����@ͨ�^E���S���TW�װ�<���9�=g����e��:���(Q��6���ܦ򽀢���,	�x���c]N"�����W�#���/�a��˧f��f�x�m�N��AޙFG��f�A*.����Iyי݀�B�������ت��H̰W��=Sڥ�VT .|�����ab����49J����`Τ$K��+������ڇ�����|򶚺�^����VǏ��=:<\�x���J,�߁��G\�D��Q̖:=��0%�eZ��E*>�;~�+��Ǔ�p����6���>� ;�� ~��n�xT�ƒ�4=f���V�r
�d!f��1��=�]��9���/<9��MY�=VB*�_^r���yT��b�Ryb@:Q���ҫ,q�\���'�s58>�fG�rN�J�����8=�����k;���v��V
�#��@1�g�l�������r�bl���j=��[&1��O��^ۏc�q����C���<�}�%�5�++;\��l�,��ώΎ����WR��{ʼ����v�\,��v�f�EzK��e���3��1�qԲz=/��x��^�q��d�+�l�wU�:9D���Fu����qs4=�����Q��ԣ�	����	�}��b����d�B�ߨ����7�|�����D���T�2����׊'`�lG���g��c����¾E��;#�a�eV�̩����ޜ�24n�%hk0�� )�~���������WǕ³�$�ܲ|��x|k��r�1�w�uF�v��ff�V+R��ޯmܛ�ʀ��=�y}^&�{+�ݿ{.��Z�Ϧ��rt2��z`��Q�S�ddw�d���P'�⺩L��_�Y|�C�^Ӟ�>>ӑ����[��m�TT�TO�o�@��ʝ��P(��Q���b멼�חS���Я'^=�=O�o�\��Ô+V��U�r���3���B��aع(�( yQ����E��m�F���_�
P�!<�����[��V�Q�8:�K0cx����b�����]5UM�f�rc:B�V�<��Z��-Z��=
c�Fs����[�hl���G�s*L:�=����[��Z�ݶ����/'A(ZQ����
�7D±Ͱ�S�k�X�$�Q��i]�V)��D9��g�K^��e���PҮ3޸:}.a�,�"t���V�`-��쐒6�ۺ��Kv���E��m�{�_O�0�ӵ�=�ԇq�������C�.k�@l��##�K������5���T}����Q��>B���[g=3��8}��oΰ
�ͳ4�R�ݞ�<�H�o�=3�Q�ߔ�Y��"e*B��y���܅Gy����O�>#��|�u�-����m�����(O^{*fCr|fc���;�B��{�bT���'�w&-��2L��t��o�Bpy$D�ڕHnw�V&�OT@ɇ�'�b����}�y����w��;���t��`�~RzX|�CDez=�t=3q��O_ެ5���,�E�}�'t�nGG���[�z������yl�-}�H��m塑�U�9��P�y����dЮ�m��NP��D��j��}iGF8�w�������T�x�9�b�|����g�_�5��y�F��h����E��#]�AΖ=<読�W�Oq��b�]V%"x�*��߆I�Mù��d?;��Vq���<�gz����(]?���pq���Wك:
[�Q��]����HC�xЏu�g/L]�.����Щ}2ͳ0[D�ֈR���ۣ��B�p�{�^�!Zl���&�ѝ�4%ZAm���!Et��L|����s����Ωg&+8��l�C��f��鸎��Bg������r<�A��v7��m�^>��_��:���f==��(Jz�~�wƝ�}��\<���S�^�u��>�Xx7��Ez��`���S���� ��N�����{o�5�+�ܩ�Y@u|f<'��L_��J}9�̨�]Ӗ��_ �W��%��������������H}�Ǹ�0�I���{~3
�*�W|��O*��M���Y|��x���;��3�u�#q�TF���p(�� �M/[���EO�������my��<��"�]F�q��z}I��\u�t+�������2w$}�$��u��;ެ�x�z�%I>U���^>���7�G[~��x�W�p}<�� rl+�-�����3~��7�Et��Pfc�6HȒ�;լ�G>��+b&99]3*�^[��w��>���'�ꌁ-�����t���4�{_�U���_:�ʫ�']U	[����]f.�=���:�7�O��g���?]H4���>#�m
�>K5�i��>X2��3�>Gnqe�<;9'�Y�v�Th�e�I཭��;�7���5�`u�%����:��<�������X�2�N�ǂ�#��`}�?�Ϛ�ob��m����}inl�Gne�����ܒ���@��kg�5C[�i�ɕZr�T`����'�8� 9_?_��}���/W��BǴ��ւ��h��9�_�^����i��E�r�qΫ�k��>����=�Q=q�l�������(���>�Y����6t)��6!T�'�B�~7֮<Y�a�O��/<��vt��zʱ��=�[,��_�V��Σ8m�*g��@��s3�t	S����O|�<2[��^��u~��<�^t�r����1��\�W�%�+O�s!U?���9��@y��� VR�~��_�T�����]0)�#��������ٍ���p�d���0��ꃾ�I��=��m���4������]�y���"�ϼw=�c��Hxr�n�R�Y'M}%x����:�bYW{h�Y��Ezi�Y�{*5��w�{N{���r7��oμ;"&낰l��l�+b�������^�<�'�����G��L���1>�w�>d��.7�<z���s�����wk�\WB:uz}r\
�@_��`)�5e"�j��^�)G�ք\y�q}ѝ�,L��}d�O��ʛ������7)����,��PYa��>�6�N�hX=ׄ�ʇ��&6����2�;�	kA��5	�1SubD�[VDՓ����^j�����q���9�Ň�������	�����jg�N'��y�c�W�Zk��G��b�ܖiA*�������E��#���]�C���^�d)��>��Y���"��<�}~��K���W�&�)\���u:��VҺ��ٹV���cx��5�����o��`�7�c=>�O�ztx�����T�&���/�-�;{ۙ{Z�Ef�-��Q�y��5q�&&9>�I��x`�x�s`lC� �J'FU�遐ۗ
�ҵ��B��������Z."r[;gK�m{n<�ꤨ�s��6����<�~����*��tk�A�o�ٓ'�z`i�s�:p;��|xdEsWᑽ>�o�.~��_��%�(�Xb�(��/ۘ��֪G�ϕ]fl��Y*�Lu@�������V��;��_��q�:�K�X�TS3"��9�(�H���zU̽�����멳���/A�0�f��D��:�`3s5v��t�g�H/@�n��ϧ���8�[⟦���:;=�!M�|f>��_�������2�e�g�}���^�}S>�i�*!FE9^��TǴ��ʸv<�Ӓv�|O��*fz��1��W����H�+/><�"��^�h�;�y��U��5G�-鿊i��7a��aq-r�E$���w�p�YՄƺ�ܳfv�G�)ۛ�&�0 � �>rƢ�\�9z�jå�r��f�ر�����܄k�9����˨"x�p��*J77j&]j�a�ކ^�{����ws*�w���3�2�Ms�W��jf
U�m<�a1��?�_�f)*괭��S����;M����I��5�&2�l��
���xH�K^e�G7Ú��9U.�rS�e�qT�C�S<qqg0�B1��-�v*�Ep�I�m79�qY���]�l�z��Â���銉�>42�v��vwz��
�*yq-�v���� ��BQ�T�!�ndK0�;/T�漮���{X� ��B�l�Y��Vq�X1����4M���%������`��"��V��t�1�qD���c0��"y,��N�&��0�G�ø�؞ar7��;�)�p�k�uR��X���CCۧ�d�O��[�;�e�32�D�>Ԛ�y���S��A���'-����]���5xg>4��U�[�[hgm��b�T.+�7�.�§k7p�IB@��vLILk.Rů{ow[�`�sF1�>�W�E�Z�;�?Y�Pnk���u0���ČZW�#b �R��)�GG�傇M���U�dfSX��
�7�؍1���J�7e��Z��������I��q�Di8�;zs��S�Mt�!�hόu1�\��rHζ��v�g��oB|,u��w|K�z��������gܥ�?Ya:���dgv�Vv�<�q��P<ô9Gt��n[sMS�T��ӫ&Wb&ˬ�;h��/�wn���9r�BG�����5��jt��Rp�@���*w5q:{����P�oy��4�m����6�ћ��_��/5G�<W�ڔ�>��ř�&6�or������	o��F�W�J�v�*�8C�%��˝z��S_��i�
�T�by���E���E/�'wz�/�&��b��M}��d��ټ�@���X�m��'J��Q�庺�.���F+��HV���6�W\J�а������+�ނ��p�u�;���e.QW�UŤ�7�Rİ�=E�/c�Ǔ��R�m�Y)�on�R����6���"�v�Y@@������%n���ӣ��Ѣ��c/��z�^�����=�,��2[+�Z6�F�?
������ۨ��{��5mQ3h�T
tʣN:uG��b����cV]k8��8!G��U�ul�%��:a�G%�' �(j�V����찳�WM޿��/&�ݒ���v�C];��p�j��k�ڠ��6�Z{�8/s��	e�U�9���˲\��N�h���\i\+w�b�Q<�J0JJY�x"�5�(�V����2�%GJQ�&C�E��ë�B���!��&�*��獳JE Q�A)+L��G��L"LP�e�%s6!NxE�d���Ii	纅W �5h{��ft�Ŗ� ��*�%
5�gRYmܯ3��8�"
�Q�[����Dh���g�Hs9D�u-l��B�Q�/*H���d�S,�+�ӡ�+��ER�rHԑI�s5KL�2��p�L��J-�;��X��P��%$<�+Đ�H�0�Y�rv{��I�Nh�Uhݢqʪ�����2������Uhj��l�bE�Z�U��e$�$2)=�s��%^��\��%	J檑��C���,�h-��-��e��
YXi��"a![(Uۑ�X�Q�2T����P�\�gN$���t�(*dh�e���H�[BL24�j$�d��c��ҶH�4S��$�,�v}�]�]�fm��dr��46|aoL&U��|u���;%A6wa�Z��	-%��.�]�̵�N�3�cs��rhƔ"��6��bN��������DW��ܞ��y��P�}>'��^>��\?��q����2�]�k׷�˼�쓃גIu(8&ٟL��Wzh5�^�|}e��z'��7�em����(�.��>�`�I���,	ȱuԯ�UL���X���~3�w������׭�>c��'�n<���3lÊ% ����2�㩏L����7��gS�Kj�,�=����l��}�U�.�!�7)��A�ҟ��]թ`c�ڥT��t�Vz5�QO����5�w��ǧ�����{ǵ���o�����UA�S%O '��?{���N1c��T�(�+=�F�o����M������qu�S�f};~�s(`�޹ܔ�^Ǭ�=fZ6\�1�1W�����q�B���_�߽>D������'��'��S���OA��S��^cTr�%\���%/J�k��~Wrc�ő�ӵُӹ�r!�̟?O@�g���?q��&�d�a��}f:w��dEj�x�F�xv�=��۵a�W��y��̤}*\j'Zy�����*���W��;�����R
�׋3*�g�VT����wP2�^�k]���V��z4�r:�S�/���9(�F���q�
8�^0���JmG�� �aɅ�v���oV���&��۽�x��'�`}�Q�ޠ�o����`�_kʑQY>���>��*
���G�rO����a�Z�]����ݠ��u��dy�{�}�C�纬O�M
^ʑ�����OT9�~�X)���c:���ꬿx�L�'�.�/|��K���g_�;�s�;���n�w�ɷ�|����sW��{E�} ��3�h�c�{.���J6r\
{�~.W������Qݾѳ.�-b���aZ��}��Z|���d��2�A<}��1}N���>�x��^>���&�~�x���A�f���b1�s:v�����g��>���2��AA����~iʞ=}�����>(g�����]G��֘�;Q'�Ǆ�*bzeO�LK�<n��S���"�*�^��X�i��g�O�w7���������B����=Qa@��}�q�]N�[7T�z�{�ȯG�븟���+���{�|�do�#q�TF�:��d�?l�j�E�cSx�wb %>���`�L���y�5����\z�i�+J��Ю3޲6��1�v�qY�u�啝���n(���%�es����͖z�6_k�WA�K��)
�w�WM�җ��*��U�,�;�H�����,q�s�7��*N�-Y�=���˗<6���_l�;�{b8�pe�18��gf�dux�r�N�|c�neI�n��~;���v��:�x~�����A���g�v�E�ކ�m��N���2�w�bǕ�)Z�SUݩL�(�B����lȧ2Z�&��:O�Ȩ�U�=�����2T	4���sI�aޚjF;���g�"�|K��F@r�E�,��3�{��;�d���u�z��A��	���{�!�>��v�C�����\6���{��;΢���ԃP���!��>�����kވ	��}�^�>�J��ϣz�F�t�~��i�
|�~�¹�Z���O�{�	�Z���5ڪTЦ|rc�S�ӑJZ>gyO��g^\\5���_����O�z���u��3GK�
f�������:jOp6t;����R��8�_��Z��D��i�~;�#.8��}�U���/�5�՟�q��F��X�|?N�qU�t	S���,
��Y~������NNVӄ����u�=��w\u^��\Ν���*�qB{�\z*]�lz���ONv+^Žr�{v�{���r=t�V;�;�<��۩�vY>�3ꅯ�ҿ�t�;��O]�(�U����eCQ�E�{��S����e&���	�d:B�q3T6���(��#zs��%�2�ܻ+K��-Aʉ����R��3[Y.X����iu�x\��Ɔ]���k�5*�fg�V�k��V�Z��y�9��X��G(̝��M��~�;�ΨC����C������1��<DM��22�$鲷}���$!�r�ٻy]�S>���u�9���!eAf����@^�i����T=>~u��u�Uf�2t�lM�u&�E�_z���zpd�>�Y��c!����޿TO��a������ܸ�����"`]g�'3������}�����*�,	
|@�H��j���w�B�>�"w�Ѥzfʡ�_�/�ӄϟ?Hү=냾�f6>w%� �������E��#�N-�.��=��j��ꋯP��W+c>��_�C���p�냦�^���d��Cpx��^���>V꼧�����3^�=��W��/��c"=>�O����:z�t�>p��Pyh<��Vjۍ���Z����tn)�G�!+�x����ED'��7�n��z� ������*_����=s\Ɲ���^ǉ,z�#pT௥uh���x���M{n<�ꤨ�>�p���~�Q�c"�'3T�m�e�A\���08ɹcl9����tN���>�{�˅�7�bz�:~q��������	������S�H�Wo`-�R��!n���L�� ΘZ��h�e9��cua��I1&��5�����s*���6m"!����]�PC�A�hFF�ՏJm��U���ʖ1W%s�Y]6�;r�g$�ΤXn�����S��=�&'��w��n��Uѯ��3��K'�&:�N3>����"V}�Lyz�Z8`k3دuW�L�P{;���+�yU�����u6t2n���,�M(�a�x����sѩ<mjs�����@
����ϥׯ��?V��~�Ǭ���T��Y9�a�f���}�ttm�]�v��vzVz;���ȩ����=��H�r��>��i�^UÝ��:rN��WJ���
<��؇��<K�_ꍺ޻�}r�6p����x������\?��q����2j�9���L��C��>���(:�3�Ϧc6�J7�V@�W���Y�7�;�&�����wAm�B�p� ��lj���X�>E���~
NhT��H������]~�P�=��U�~�>;o����a���_B yT`L��@�ۛ�RE���R�e��"��V�
�z�y���w�iWꁆ�*�J9D*3��*��e�5Tk�ԕ�'�O2�=1��}�qq�+C#ӵ�ߟ�&�=�#n=UaL�/��]�W���A���m��*���WWf{u��l���d�������A2�f\qp
�q�ƢF��`&���{ON�<��W$�R��Z�Z�����LT�r@0�l
kQk��.:�����P�]:�Zg^3�G,|]<����x��G������>�f�Q���Ts~����x�mx�<� ���p�<2^�s�^��]�j�W�,�t{�����T��%/���Tu�����ޟ"|B�t�� �`��ԪG���u`
���H:�?��R�ե�K�~,[��ԩ�k����#(C���9���Z#ɍIѓ�z}���>�$�"��0���TN���b�׸����T����[۪2�o��]�c��R-�B�L�;�`�Q��d��d��;���4����i�f\���G?է�~�~?�*���:��2<��#_�x��U���{&�G{*Fid�?5�~�2���z�SCY�u�-#$���˥��u��ȗU������9�u�u�C^[���<��RVI^�=,;s=�����˽ /���8��w�3�t�|Nz�<{�J��O6����[ПN�.���j0�&t_��t���Bg�����xa�C�F����	�b�.��2�g��WQi���C���Tn�F3�gMO�Dc(���UzOS�˂=��'���� nj�����!c�Y����Q�&���xJ�Yk��sR�D��[�_7���mE_N���h��s���G�	.�㜆�m{�x��F+��9�J�:Gd�(�oY�Ğ�J�|�r�08��1ѩj�Q���rݥ*}��u E���~��ީ���f��.ʔo�,��f�A�LU����n��'���e_x$:'=r���*'�#���<�/z�d{���s����qɹ��rQA�W��M^��2�#v[ŷ��Ӈ ^N��u�^C븟�_��=N��<���o�iQ�TF۪a�a~��b2sƇ�(y\����G��5%�>�x�t�^k��C�+���z�9���_�iW�� �j9��WM����F��o��3Q25
E$\�\��~,n�:��T�9�6c�V~0�U��N��ϮT *|������z��z��E9���Ʀ��D�^SB�:^<����F�%����:�:����k����g)�\:u T)d��z�lD��Q�<���>��Vg]���U�M�߼��~N���w!�>'������	~��Qd��2�nQ��j�nz-e���{�ܧ�"+e#׽Q�*9�o�!��ɸ�����~���b�;�R`?Rj����ܛ-_�=ĸ/O���w���}]>G��)���˅�߮��P�9{��z�b�J��x�>�"���������vrf�-pǛ�3�m/$@:2h��r�ؼ}~���QC{�½N�M���7�ĝ�Ap#��ŀ�rpxk�o��h3)X�َoR[���k��
�*:ړ�Y$��|���+x\�PYJ����m��n���G:$��C�2�g/��A��V6t;����WM�F���3�\x�>���<���~�vZ��}h矮�{�ޖ?36_�����χ��l�wU�ta�_��;�n����՞=��^S~ԊEl��
N,z{޿�z�<{��vug��T�Y;�fA�,m-��1qB�������\�
Q����
����S^��z����t�qvxw��S��|����G����
|�w�+�W��W��M�� �@�]�y}�"�{+ޞؿSy�<M��26������B��kh���%鯌���WM)>W2%�����z��"=�|}�����ׂ�r�WU�*d^;������^az�])@�İ,5P祳��]O���V*��w�9R|_^.�_TR5��;����kѾ��f�w �(҂�,��x������#��B���W��/=���oٶ���B��t��#[u=�aع,��	Q�1%��,��9����#��j�K�^(��~����O�0�ӽ~�Ը���޸8���C��N�{�Τ< {�u�-a�?�Q��Պ%'�AZ8���r�F��3E%B����ȫ\��RY�>��*6��@6s��f��I��iL���,>�Z�C1�-V����id���r�[l�'E�|)��ӌY�J�UƟg,G�?�SȚ�C��깽�z����+��+��cQ�d�ߝ��z}H�`���>f��n�j�}�/w��
5]pz����L��1�*2��V�\?�&7�W�7���������;�?����ފ���4����Ͻ8N�3>D#c"}բ�+)x����񶽷�j�����2k<=}3Ӎz��ӹZD�纤w��~˰����2�Yc\N=+���j�/>ޯq���ù�s
܅w��Q�H�wf=�Q^��=�Bz�=YF�����pɆ�mhwU�:9D�}�zE��,�z�I.F��w��}�^�����^ǕX�ٱ#���cv���|'4�9��0&�S����/[>5��{#�lQ�W�K�^������/�hn����'33�
���ZU�Œ���F�S۾9S>�/>^ S�?d��)�����/�=?{��;�}] u��M�˞�;Ca��o�b�Z�y����u	Y���%)�ȇu	�W��f[T:��q�c�	^��vZӒt\E�$�D���q]U阸�u,�ϽVD�x��3���>��3��S�J���ǵ)�"��\ن�ٚ�ɒs��:�hA5룋�󜍻�KǴ��d��
��H�ҥ��l���o�aF�{h�345tu˘�TIĵmg���2\L���
;y��/m=�q�#�ޥX�V"�29��d�w�<>�NW��:�j�7ƾG��7�� �,ȱq]J��]̳1oc�m�z��v�5^�X��Q�
�{���yS�������x���F��%W�X
^��ݞ�Y�+�J7��E���U0{���p�z��F}���V��iW���t��糪e���}b�CΏ%�;�FA�y�<VR&��/t:�F����z|����=�ԇy�Qz��5n~�d��M���_G���<@h�rD�>u���h�w�j5�|�G[~�ω�>�q�Z
����xfB��ey��
�����ޙ��%"$�g`��?D�Rq��Ð/��{�����_����o����)�E�O]��R�'���x�dG� ��4�d �H&�U���xи�-��Y�T��r�1(���k36���\�3����fMǽ>��ȇX�O��5�,��0���J�e�;�+7G2tQ�O������:����1?]ȼ~��n��z��X(W���d��d��i�����_�[�T��8Ǜ1s7O�+��oy_������:�q���2��bt��ɡ]���ux�;�~�/���H���u,�E󦝈^��5z^��yᜱ�'s��\���L;%��1�2�W�K��	�neS��گ�-��]���`kt]�6a�)k��(Ι����������f���S8T[�Ld�u�vDĩ�i+r�ϔ�0q��9Ñ�mKd۫7�rԗ����0���h�yu����Yنi��7��6���Om�!��׼����툕���z��Q�X��$��)�pn����}�#����_��$k�y���ׁ�2�t��+
��*�[IK����VY� <WwP%<�LL]#ۥV$�c6_Ɓ�˭ے���$F�[R��kBm��N,��b�޴�YO��x�>J�XN���(����K����O#V�买'wk��G�^jxE� :��c�뱮D�&�\�����0-MV)wSv�Yyʖ���{kfʈ�_Y�������o��x;y�sU�3N��VdC��!vN�z������(���O)bɘ�P���A���S3��=ͷzXS!8sf���7,�9Ϩ4:���>�w@Vy]�0oPl�\�6�ذ�z&���bVZЯ-�@ݵ]tEG��¹e��)�$Rٷ�n]iYD�P�h�-B?��rn�}
:��Eժ��۬q��H��X����%a�Y�NKOn��v�Cpb��.꽦2��|��B,�i��Ҍ�΀
Z��*�P
S��	6f_5���p���8�J�Wl��jZ*m־(�\ٷ�fk�F�+w,m�X3��[ϓ��O�:�{�Ӄ�7٪�,��[��鲱�႖!�����x�<�^
Uy���OS]���O��*�+��9f��\lӗ��!� ��.]��/s2���F�s�s����	�w�)t1j��3���U�W�,�C�*'������y�C�T���u���R�@��cJ/�d����VX�@З&��].�v[*�a�2U���"��t$�u�Zo���vW8f��oiӵ5qu��}�a=.�|��:v����̸t��M�ό�u��i��r�;b�ٰ;/g���HiU�h5�LH9�V�'kiuu����<Ѯ�<䁀��F�[9��b�B��*k\�&e�Xgv�;L�̅QOr�/�[����n��Y��#�˯�O+Y;E���a�v-����jj�T�n�3\�kL^וV9�mp3%���ׁ���؆ݩY]�;\�67p�#��+nYP
�>3$��h�B��o{��oN�ك%gvY�Te��F��ó�-<m)*���ZM�׵�����\�d��݃�բ�F,���(ڬs36�Ts�v`]�ro\�͢��f�h|i7/�pylZ���櫠[ܧ���l���-a�L��Awӟ'IՍ�3s,��� �qJ%_V l�lt�v�;��V>�oXxx�&qy�&�o	z��ԣ{�[�o�����������K��D�EB����:�RWJ�tu�㬔�'5*S6�qC*���*=J����H�,�[�vQ^��MCNNn������y��F��H�X�5L��T��tK�܌#D�[42�8��NZ��aE�{�������窅��$�d{��DK���5Gq��XQ�Q�wD�QK���u!�"�,�SH-�s4B�9��bz�I+�Wp�%*�J�ʕuۈDQ&��U	���B�H�d�I�e�VR�K�%��� ���
GMh�WOs��k��p��z%u<У.��NnR����v�{�p�q�
�����랑IG)
��2���QWS1:DN��faEF�JmB3+���0�E=[�b�����e�r:�`���&D����D�c�w2,�˫�I�)�E���gg*|��,ݺ⠺Doh=v�o`�e��e�XZ�l�����|;�Âq����Z t.Rk��8WM�}Ŀ��7fUe�r�_�K��w�.���~��9��ۡ �:�9�=����]O�{峒s�i�·�Yw�I^%��Y�LK���j���$��b�N�)��Fo����֖	]�9�A->z�g�t<�>;>v_�h�u�|�fuV�W+�N���U�|z����ڸ��u��geN����2�W��'�}&��1��,�;�k�	dd�E�����"ޏW���?��=��ߡvT�A�{L��>zm+��&1��YU��꼡Rǃ��*sٕ��o,Cς��F{���s���~�=�D��QD������RȲ:g��%{�1�'��L��l���q>7���qW�w�9r|����7�DmU��e?e��+�V��5���*�� s��,In�ql�sC8�~Wq���s�;���w�S�Ç�sYڻ�
���7��u����H,�(!S� �<q~,d#�\C�Hvo�cz ӵ�����V��"�Zc�w��>��_�Ps�U�"�̖��50���"bJ�I���~-�X���Do�.�/{�?�^M�*�y�|=�*�3�9%8���|eZ��{��>ltGma;�)��.��.]�"��3.�o����Cq��;�wZ�B����@���L��Ⱥ�����no6hnV}�cԥ�uk5��
G�%���z���d9��C�Y�����j�Ͻ>V|p�wļ�Td	�N�
R��0�b{kw�o��*r��+���+�G�W�{���\w��𿟕܋m׉�@���|�0O��R)d�Dޠ��;���o�}c��2����9[-�����㟶�2�\�~����}�*��{��z���Fn�oԻ.� �=8N��������W;�9]-3��K�:��7�+�������V�s��=��}ޥR3�4�CD��^ś^,�7s������}�/��\zq��� ǚ��v���gǣȋ���U̽���Y������|vv�|?T�fr��4��<}�t���N��yn_c�$� ����B>~����~��7�;=�:mN홇��"���x��s}���s /&}�P�L
����#"���T�P��9'�FvT����2VoF;�р�ʻ�<�E3�3ꌸ����Z�<�w��<�YJ��k҃^��"n�O�K�`�o<����'j�#(�%ILѕP��K�U	e󪆾����t�nD{����~B�����ո���f��5%q�.�n6��=2s��R~�}�9�3��G��g��u+'Z�Dr�W��kvn#x�K u;{�{�TK��[�sF�GJ��*ҧcq���u����}������s��rEeI�._Lj�rXf���Lr�?u�գ�u���K�%�p<��Sg�!�����4+�״�w��꽧o'� �����=�T=Qm�p��|����7���k���ݾ�m/L�=ԶS�ꋯP�}���"=���{�a���ˏ���7+�-������Q��>��8����B�j+�N{�΅~�Z3��y��޿ߡ��g�pt�G���,� 7����v��\�on�3�KdǾ�t��-�:�w���4[~vǏ��ӣ�ߜ���I^��yst�����z_*��_��Ѳ��*�R��^%p�n<���M_��ޔ��x޵�v��MǷ17��
g$�N��͕8*_V���)x���ҡ�mǟ�T��z9]�q�x�R>���d���G��W�}�%eH���@��sҸ��j�/7��}܇du⊪������=Wz3�J�Ϸފ��������ٛ:>_�j6t9���˦�a����)���#)�/����xg�׻#z���X����f�Did�Ѝ�W�����΍��I&_mGP�;�9wVn��n���u�:1m����
�ޘt\Pu^��#�R^��݆6�246ٿ�\�&���'�4�b]
��Ԥ�S\K횗�.�`ׄ�]M ���Y3��P2&�r���[��9ըy�����DU���`�W��׾2�;��uc��vO
�eHǝ�P�ˋ�9Q�{��>�[��#�am-��$��'�|��3�r��9��t�9�Ҝm{��Ǯ=�:��u>��Ӓ]KK���u޻��\2�z�v7��[+�ڔ۞�pa׎X"gV����}����;���9'Eߤ��(z�L�w�^���2�>�X~��p����	KU�m�(@S�}TQzs��~+>�[��a��_#�e�$�,E����ύ�>{��;�/z��NDۛ>��X��w��#�z���=�|zߝǻߌ;�\�j�%T`Y�*�Ѻ^��MUwx�{� 3˧�o����~�/��z3ϫ̭�Pҳҁ����;�rYڿ[j�L�۪����'c�xx@K�g@[�M��l���Q��Wq�,C#ӵ�y�xi+������"W�'����=�4��W��L�Mq�E��p6:Z>݆j5��Ts~�ω�-�������x�&��R��}��TG�њS$�lԶl��2�HUҦ�@���
��F5G����o8}��*TX�f�D�l�5|��{�fIkS���X�p.�Y�Ze�߇ea+1��{ǖ٘-fE
IL��U_�:euě�a�z��Wuu�ܭ0���{���tݳF���Tu9՘f�zx㼣nT.��2��9����� �J����i)��R�O�A���<��C�����]�P�a�-�X�<�KVϷ�ɬɭw��ZC"}�}�Ǽ�������7�O�w����2M"�����b���˳7#�Ւ�5�e*��DW�{���xu���1�'��!̧��X(V���e��#�村�߯g��j��ފ~�8�+�w�r)KG�y_�μ��<��_�x�~��<n=�ChM�R�sQ\���,�>����;#�wj�e�%�:zK��w�.���~��9��ޘ��0������ց��C��s�r�X:t;9ӡ�V]�ʙ^%���=�y���ϩ�[*#���s�=����Vq�>ɝ���;s,e	�
��xdt<���ۯ	�w�Zk7�����\�Լ|�_�(v�;��#�3��'� �BiV?R��C<f�-�s��W�O����`�Vo���G��s��~+#�H{��]s(�Yd��#1� t���m�r��S>�;\.�WJ�w1-Ӻ��^��p�x�o�u����&��/Xm��#VkE��m�K˱뱩�h#1K=�)fZ�ɞ��/�B+�z�&8)ߴJ9d�W��7����v�NZ��u��!5�͝B:v|"\��S4�V]ǣ�(��5t�T���R�I�2��xz���N[a@e�,���,ȣ��fb�P7�{@L�ݪW�R�LVv���_e��G�x�'�Á0Z��Se�븟W���.���r|�7���BԪ�����e�c�0���mW�_��>� )�,LAn��:[/5ՍG!ߕ�_�֑�1A�WE#^5�� =�_?Hү�������3QdiA��Q-�p:_��:��=>��>͇w� ]{���NuEϨo�]i����_��>��m��o�^2+�2Z��S��^SB�R��5z�v���6��+XSG��}�,;�+�����<|�������[�@q�;�*��hmeCHqY;��E�W�s�=�N��Kf�*������~UR9�^'���;��0?T�3�.7ޥR=3��uӽZy�ǉ.��VTTJ��9[>��������������ʇ��|xi�Q1�&�7��<k|�}���H<Y*�����W޾�WKG��)�μ�Y�~��3�
�Q��c�-��p�>Mϟ��z�eЮ/&r��`��,(Á�V_��h�r7�����G��1�Iff���+�g��<�U�/c��'��f�g�*������X=w�"��,j�~�ʚE�TH��oMHjS
�K��Z��������ul�/E��h��}BG�s�n �Uʸ�b�w�q��XQ�Rd{|1��NP��V��	N�	Qɉ�]�:���Х���l8�MU�V�5�k��Z�H��.�tԺ���eN���Ŕ�)����� *����[�����x�C�X�Ϻ��W��҃'3L�̋>��%��{u���{����m_�|iP��k�=�/
���T�N���xVvT�5�53�A��Y��C؇���3Uq\���[���P���Y�W�=^�<����Gr6�F��j�r�?t�s��nd?E�$�!3�UC������dK=����ޯi���iƖ�ʸɼ���w>��=\��adM�d�S�I�`H�wWSg��L�����W��u�gf+�.*����2��]�G��}�#}#ǯ<�d�]�6
5
UX��-�;�
T5�\����r�z�$_��=}HUǫֆ���[G~�Hҳި9�z��v.K5�C�@�N暙���6�+G��u$yt�3���hpϽ^v�zw�÷��\M�pt߫�P̖T���;�-�%l������/�p����Tn+������5޵�47�L8���>�'�� �,�h�Mxm{�w@��ys�}�'`���Dľ�Q��-��+��q��G\&��n=�R��?+
�
k�>�q�z���̵����&���w�X�tPp9���W]�C��R�fk�
�r��k;¦jQ�H�č��'Ը�a��m��ۉ�]����(Yd�S}@�������i�p��;Tk����X��G��w��\�����0C��y�E'm����Z.�����>'�A�~7�S������z�%/�^ʏe��=1��9ђ�9z�Dg�N��2[r�|��Tq�L�a�:rX�����\xesW�qC/�W�Q]���L֬�v���O�=yp�<�v�dk�W���U	��e���,�PɆ�և�z6.���}����Py#�c|��u���G��ǯ:�G�|�{�2z���yU����Az�l�id���y�O�ÝYҺ|��O���0�*���A�\g˭�/|��}.�{�:�]��άw����ng��y�:��W������wA���*�\R۾9S/ļ�mx ���"Y�9>��Q��ױ��zFH��s�sA����'�b�{)
�:rN�d�f���Pg��w���uˁ�rz�v7��j��1S5.�ɗ�� <��z\/�z��vG�Ь��:)�OlJ����z|���T��s9�r;5�zo�P�|n��mi�~��N�ڠ��gmKY}(�����W�qZ{ଭ�io*���:'+�ϞeOS�׫�G���7=�|y��{T�v.J5�>$��C��{� x��:+dlt��p%ӟ]/���3+C���Ud�zv�*l�A<
C���ɮ��8l\��cU��;��:�ճ�䎑Y)9N:�K�FP���ػ"�9�9�p�H��H�^.A�@�����\�EtKp��"H�|�� zE��7�E�\�9�S�=~�=/Ճ�����H����p�N��л�y��96�e���Ə��@ݨ2��x��Ҽ^�u���+���Z�Nב�~�8���8}�����G���w����S]2\�"���"e��c�Gء��E����;>�b��=ܭ�b���r�)uh7�u�W�9�f�L��lԶl��1/ԅ_ԩ�Ð/�GG�Q3��v�}�{�T�[�1v=�k��_Ϡ�w��>u�O�i�ȨE���3�`,��{� ���:ڶ�e_�;��^��yS���#��]Ɇߨ�^��ý���2MB,���L>Ο"��1w0{_e���O�}�'��6��î;�xO�Rc�3p�>֫
ו �=r]����{�Euvx>%�t�m�'tº�{�Q�>N9_�����ϼ��#_�x��U�����}Bp��Z�TZy�#/��ڀp{���C���=S/�⸿�u��.g��~^!�c�:M���B�?�Hr�O���ρÛ�xg����*��J*>;.��пr=����[��ȷ],[x��j�gw�QUN���ʚ5�HMН{nR�$P������Ja�g�նv�[�0#��N�&�4[W�{�)P�E^S՘��xP\��K�N��Z��5�NV�駯���"Ȝ�F�5vd�j�^b���D6�wA�Y֔����s����`�.������%��8����^'Ÿ�3�]uz��S*��f�sע�j�F�x(�,Ct�|G����v�;��#��:n�'����7��4�=�ו�����.eI��Pe�zh47��E���~��=t�� ��]�(�ws�U	TK����!G,��$��>5g���]T�Ӑ�*%�;yb�^���'�;���o�Ǹ�5�̟(�m�`��ܪ���%"�>�1��X]L+���|n=~늿S�i�9>s�ߦ&���V��B���h�3�Dm���6J�� )!�����O]X�qߕ�e��E���Ȋ��}��+�/էޙ�q��U�do��;�Ae@��#�[�8�3bWVY��ǧ��7k��8��/�P�}���c#ӽ~gO����T��^2*�jl��q�F�S>����{="��{�SC��^G�>q�W#��x0���Y������Td	�ө:~�U���?�˙F�{�Ի�R-׬�kݳy	T:֮C�Q�J�.`oB���`�1�����cm��`�1�����cml6��l����cm���`���v�o�l6���6m��`�1��M�`�����cml6ލ�`�����o��6m��`�1��M�`���v�o��6�������PVI��|#gM�ⷷ��@���{�d/���]�� >M���T�41 ��J��$()Zh�P����&�hրj�hh�Yl�S��1R����[kbV��fѴ�����4e�hm5��J�,��m�P�i���+�&��2�k6�m�ڛM����F���l�k�F��-�3m�H�VL�M��=���԰�� w�`_L.���hd1�ՁBɊ�Ɓ��lL�����j��Z�m�� }J�ΠRk ����=�   �p@ �{�  �w   �U�p�4�o�ى,ђ�  ���$�w7m&����A��x:��Op4;zӮ��� v��l�w��t����]�)�m,�V�� ��o�=���������7����롽a��z�zk������zS�`a=Z����ecWk� ��EU8��E|��v�q��֒�w����{{��4s��.�ws�
�s�:hv�d=zu6�ʬ�ɪ3u�  �6Eol��aM�>���C�e
h��9�h׸b�k��{��MK��� ���{=P$Uzz�V��䭦�f�ȵ�  3�P�(W��ܣ��V�T��i���e%@w}�yOwuJ
[R�Yn�9�h֩$\m�Քƨ}� �&�+��۠�!��t��Ӯ�����GU���ʫEi�:�uґ .�۳��;��5�U6c6V�� �ζ���"9�k���)�Xt��+�9��3��	��]ES��v�L< 9�n��Y�\�4WYӸ�U�`%�; �r�C7;F�۩�A��t>�       D�¤��@dh  1�B)�)JT@M0L�0� ���LE=�R�T�@	�  4�~%%R�       T����)��       @&���@&��AG�e7��m�OR~/ɯ�������9����~)g��;J.�C���ǠQe�v��D>!���K�� /�(*�YB��0�����
(�Ae�߿��p�`��ҏ���������2ϸO����$� ��Bab���ظ *!�"a��db��(���!������狟A�_��?����<�[��I$$�I!$�Bx��@PJ��*(TD��PDB��T P���QR�Aj(�QU�(�P��PB�
EU
�
Q*"
T@Q��$� TD����{މUEUTUUEUUEUUEUTUUU�����>=���Fe��]/���S�{U����+~�f�K�2{\�ڽӦ'������nm�Oq�kx�v3���,������#o+%l�oR$,�jl��i�*E�w%, �1H�EÚ������K���"��A*�ջ��V�����F�f�S��V���N�V�"ӷ5�#�NUąѕGE���yGQw�N`s1Z-�jU�.�]�Cst��:phM]�hn�<�D���+,��f�56�,�Wb��Rq��b���������M�0۪ۢB�b.���`�sC��.;�6�*��	��ۻ�7Z��T�ޑX ]WOJ����ܬ�ݎ
+t�4�}B�q�\奖|I۽T���yW��N�XQ"�**�?SX;�D[���`�#n
xo$�.��FV�����c�a���T��O#Y�Q_�k����1�6� ���0�nU�E�	����V�#Gw�;3e6fd2���x�$��/�mޖ��Q�Z��`�V�.M�1��lhц�]h����J�e���3�#Y�]��A�:F���5*ݻ��i^M95�4C�+��˕͊�e][k5Fk"�k��j�7yesi.�|Z�n�wy���*W��c��Z]��Z-�qN�D-8����y�m<I��B8P�^��5/��`�OƒխMZ6-jV\���d4Z9��H+Z~#]#�uH�e��1�0��s5�9*��9&|����Nd��a�"�j���b�Z����ϙͻT�$A���A�V��1�P(V�/oqĎ�7uj��R���s6iʱ���2Z{��dw���Za[O2�+���Q�����y�����rS��/F�j�8�\̌]B�ʲ/#N���H{�U�Z�ԬR��Z��|@����yM�+Gyf��� R�+���vcF�S�����S�U�{t�4��(ъ��n��U��e޹Y
w���n�Ȅi	N4Ki��K����&S4�1�{��	�D���ǮP�P�E��ZU$�ǕN�,�/2-#�.�FEQo!��'UF���9�#�s�5'p(*fJ�(��ea��\D�aU^�^�"X�f�����J'6rΣ7nU�U7V�Fe\d��8ؽ�+],neh۴.b��)�b���}n��l"��T�b�[
��4�F����B��5�XRM׬"�J��v^f,�U���X�0����V���i��{���B�׏�խ�g�O)L�������-Y��;���TmQ��9-�Z��{�sSqH�^^]���y�$k�iUw��<ړY��5��M�����O�ٷvط���CJ�i9f΢V��͛&��rc:֦,^ܒӠ1��#,��.�sj�qL��F���w�������m��;4�Z逸٦���ٲ4���B�˪iP��:Kj\9�L9Yy�D�vT�%7J��ok\t��b����L����F2]Q���p#Xj���d��^	[��&K�l[��e.Zާo���w�3fe�0�]I*�9���5��K�^F��{�N`BJ�R��:���sl=7��ZMᱭ�@�(�icr�e�h՛�K�s����g,���a��)�M�'S�,_0�)�,��Ag���y���x�iۣVP��
;�M��ͣ�n	�7��^h�.ֆ�эb�4f�x0c��ګ96�]f��ۓi��k^�6��;w#2�^9�\�;��{L�^��!.�G���ĩFQ�%h�3��ܫ����5���/��i����c��ES,v��tp���ܼDm�l�gM�>��o�[E8��pr���P��3�RJe���rH�����e�nh����,K0�r�X�b�5n;pf�W/Pt2�՘wt����oE���ZH�;H�4t����+��ҡ���D��������t.�vD7Q�*��r��7rcu6R0�eUAF�i��`�Ue�en�R�����5@-�o7#�sf���*2�LF)-��WUz�U[��n��J����{s�=fˠ(љV��)271�L��v+�Yw����̰]_Ɓ&l��ƉĬ���L<�N0�0Oɽ��@��}�� �1V^��+8����oS�
ը%p�C�.����h�Q@%���U㵄�o$���ނ�H󼐉�ŕ#��ާt��oa��ݳPm��&��[��Z1�Yڕ�(.� ��Z�erͶ�_``���T� �B@�ISucmˊ�)Y��-ݖs[�^/U3����X��f��T��c��L��bU�fn#�k/���Gq��:Ҧ�ċ����N�'k����jӀ��0u�O6�e)�t2wej�v��ֶ��m�o5 �kզ˴K�T�+�w�<��-�hܫ�2��;wr��6�ؒ8+(�W�-�pa�_vY�ٔ��хL�&�0�4���D�'T5b�#�"7y�Yz5��srPӶ��*b��捪�XqPu{���9���G���U��t��ݗp����B�(r/��Ԏ�t^����֭�n^݂K�ʳ��R��*�����Ջ�P�h��)�v�pěCo;Y�.u���,�A�u`f�4��Zt�2oK��C�(ԥ>,J`Ğk��1R�XR[X�����3u�D�7�oFS�a��n�'o.�cb)^n[�4�*����Yy#i$o-;�oD�JT��*�m�ˑ˷f�=�|[!�Ծon��g4�n���K{N�[<�/Rz���{�Z�VQ٠�ͷ���*�A��{u���VI�hч�D��6(�
S^�5Y�{7ADZ���N��Z/hX�.uJ5����YWc70lܘ�^]�Vhg�YoN�����pro��{D6Y(��M^�f�������b�♗ �9�
,L˕����S��ѓ1�]��4)�a�ۡwx�Es�A����V�*��Kpج�lѲ�\fV�z�z�c�UI�h��)�e詗uX�N��b��,�o�<��o6�R�ż���>�z�MՀ�*��-�X3�����[K�e[������<u2�H�#�s+a���*�j�թ�L�n�,��OTAi�(1k�E���ʣgN��v'��C�ݕlTV!W)+�E�hի�xoEQ�7�wl��w��л����1$�tܕ�Ƀ2����;�����Ƣ���&)�n4U.��q)��㵔XmY�Z���1��e�y����8�V��4��u�йc��V��X��$)�/��{H�Vۧ��*��w*k�[[X�/�C!&���7�� ��K���p(�5ѱ����^��[Z�b��J��{�ōm�����|I��Y�-Pt��$�	f�eڽ��\�{����o�I��jê�;{���0����Lr�"��95��W���	����uY�v�f�n��+XF}��0���R��5R>�d��OQg9�t���=`%\��|�V����S*֙&.��
��P6�v/�T$twqe��ч<�cB4Ͳ2�h[Zwe�WC0c��J�@��iA�׻�4m�N��/hd���E���o,U6m	�ǩ�ƕM�V�/r�YALQޣR��������x[�2�A�d�[V5�f�͘1��e�+pۓ�����U����`;O`�/%����P=���W�ʮ��E>=��Ō*��Ry�ʘ�V��BH^`oE�ś&�a�6�J�wy�˸����cڷ�%�UKQ\��H�Y�F�W�u7l9o$H͹v�"Ԗ0ud+�R��X�%g�:��t*H�cY���_��kKT�o	ոe�����N1�Z��#L�m��lS;b��8�&&�R&R++XF Udݥ,�ONL�����0��zP�n�aR�͠-WkC�h�[���E,뼽��J�^��6��*ǚ�^e��j����͊���b/��w1�Ct�ʼ;ZKĜ��y!��1�LV�N�l&�-�Zu�F�CƐ���M��y�$�<�)/���7�L۵�΍ǻ�)GT�0�S.���̤HP�e؃3%�z�m)i#���j�AV㈢�kܣI����[x��ȱ�X�hS��?��3j�؆J���G#رY�)jB,�T7h��v�p�h�J��m*ž�f�Xέ"�Ӵ��^����.�R���/w����k�� ]�G�oE�\�_7qiï^�u�3B��FJ�������<�e4l<�u�A�EZAL�n���,�i�Q}�f�YCh���R#��(�i}��4���Vm�֛/n;�d�]���{���r�];D.�^;�R�!�,���J�]��UH㬥wr�g�(�R4�bo��5�Y�-kQ �;��J�a$���<5H"�1�,s�1S-Qp�EKT�r'�~���?���ŧ���_.Qā?\}���؜�
KB���|_��'�&��,eM��.��%΍�P9s��.���=|ۆQVq"⹁��fۣl^�|�qA�\�`��6(�ANe�SpQ�xc�5�y	�B��z̃N��Lk%c�MX��i���10!��{�WM�\�h�*����#��x�㧡���\MV�޹�nb�
��ؖ��ZJ��ۗ��j{�pWS0��,��h�s�mL�r��Ѷ��񢻝�Tёfei++v2�nv-R�g�!X�]-ȫL[,i�u&��}*�ҵ�Q �R�89ؖ��긳1��uLۨXEnC��=�{L��.9&�Ҵ8/�q��LY��=���z��Z䕨��xz�T�$�)����;��n��U@�7eБ@���kA*�nv��nuM,���U�����N&���m:���nsW�̵܆us��rq��f�Y�:����2�)Ňn�]�b�F,�Wrqk���Q,��Di��6MBo:��Ghre���i��SF�v�-a^��x�:$���t
������5G{�,��jG�z��է�������):M�\���-��Əb5���5-�	]+Y�'1�r)���rƳ�3H�\5�ۏ9@��vٔ2��^5R�\,�h�#>B��߁�^f*f����d+v2��
�M�]9��`�֫O>�j���>�|H=��b�w&��+2.�U��i�례uv��`>%�һr���V�$}ݻ�K(���,�;�����UrE��sr�-�N�V�=��8e��݆�I�48U�J�V�1�4�uF�B��	Wl那�>�hP�Þ����?a9�d)і�$�i�m^���;ۼ��:eg'ݗ�rcC x2b�Qa��dz�GN����y�/���F��%�X�\4�A�9����w�4��ѷ/�CF�\��kݱ�����q���wҪdمbr]K{n��{ɉ�8^��x[Z�L�R�ǣ��p\���ǧ�B�R�GV�qx��>��q���o7U�Ոgf���Y��q3�˲y�B��G��ڤ]I�u�컹�.ī��vp�������{9ͽ�X��˧��C���A��9G�61��k=�
���,v��f��o$V��)v���f*<���ux"����,�IXrf�sj<'7�U�}����['��Az�|�?��G;���ǓS<,M8���X:���ɮ��B�c�X�8F<��k.��Ȳ��Z��;+�If�`�+h�8�"�b�ܔ1Y� ��s��
b�*61n�:ݪ�]r�W�ֽ���ݜW3�7]4+7��!pV�4Ş��6�R2�泷y��U��lO�[Z�PV.�Ҕ)B��\y	[�sy�Ll���P2��Ӷ�n*YL��K(M����bA}���U[�F���1��<[��e��m.��m���I�1��ν�ޑ�5�R`�:���i�{.j�|�{�g�+v)�jt�a�[b&7N�g3,'�	޸Dļ�N�:V3��+Jz;imt}m˙��1�����?;����4ɐV�6����������o�9��*�I�M��(�ܜ�+��<�Z��1�5���x�&�����b��]-;) �R3C2�}�oz��2B�D��]�x A�Ƶ�Е�f挅�����^a�1`�b|t�y7_T�X�U�V�&���F>9H7;u�m�*񴺆%��#ܚj\RMf^r8��ggVŝ�Cc��[�k��e�zuf����mX�:�i!�ͭ+,�R��sVw�C5&d̮U��xo��e&�]j�4�W�l*�0�ޢ�:�s�0f�S��f4�#ו�V��(�x�u������ybхE�ɔG7�w��ּf�V�:�s-fP!a�/maW��5�-a�G�����)}��3����3�vR��*.,�R�I�{��()^��X׃�F���ܪ;���+L=��lCk1���loM�#��hRq,��9ͪ��+�v;e�[�A��oc����Yu;sM��*��$7�"�]Y��[DV��[	j���=޾D��U>�ΰ�!U/������:��<C����Ԝr���u�AA�{{7a۲���{!���V��hȨ��
�N����յ\{}���00���Drގ惙dq��|�!��8r
D�Q١�ڇ�@e�y@I��i�U��sBJ��	%�@���r_�ʸVn'�
�Zbs:�I@��9u4��Odݾ��Vq>�e
�y�F�s�-ŽB�0
,�s���TK�8SY[���o�B]����fp%[��'��JT6��:gɶ��s(���7�HZZ!5r=]X�qgIv-ʾ��#]�H�[ٖ�J�S*-)欗b.��)pԭ"�m�����+6��,�vˊ����lǘ�u�*���x�n�r����6�1�m�&��j�63��].�Ճ��\�Qz�M�wZ��"�v����u@��GH̴2��h)��ujuк��B�NwG�#��6���>�Gb��;��$ݴ2P��t���(�VL�uv3�_;[U��LsC.�%["eN�gHsݪ��������V��vY�֩j��\���'�ww��i�օ���-��8d��tMp,��e�� �����u{*��a�9��'j�Bf��lի�j�eՙ�W����;W3��Pt"J��h���ݣl�vn�6�V���rыO�I�bT�j"��U���&k&�')���U�w&u<�yH+�bʀ���������t�ś4���H�SR�3�gw��m��T�I|����ի-ӄ]X�{Vu�t{�2/i}��EMI�F�q,��d}4�Y b�bRV��30�r�Ct�n\=&�Z���m���|�]>��ǐ��겅уn螑F����4�F�]o<ںI
���4�c�g�sG*Z������t�]����.�<w�ӏC��n��$��V[I�����`��	91�r�iV#�x�f�I��))]���3�aQP2U��I�Sc�ֺs��i�%�'*s�'�
�eD]ؼ�6k�����YI��޽��fs�&��*�K):��)Cdar}�e�Z�w{X�]m��)zo^�o��BO>c�#�9H�����}�f.��PmT�6�
 �<���c�������q[�K��;�������+�Wa�od]���4�uZj�%Rs�`:��6���Ӕ����wF��e���[�+d,Nˣ��A,�މS�,��|�\-���oQ����\�Y�K|�-2��i��"��l���viLf\\�hpl4�U�2�V�Tw�ҒD���0�9EY�����v���y��ſ
��1)ȹYs��x�#����<d�xHW)�[Z��֒ޠ`+�6�sj;fR�&�5�oe��!���QͲE10n�b�:�r����1q���ɚ��ܕ)��G�v'��ӭ)[׷�:+z\�T�p}�\��RZ�*emEx㒴�oAt�]����	*�Ƹ��:vh�ٻC�i�q_:4�
�2\�'�K����T�0�4~�y;g���A*--篭oW�Y�[ռ~�)���
��܂ݜ�v
N�Zb{q^8Z�d�ѽfvg%߀Vc�(˾��vq��9Y2��ڗS��*�	{6�n@97�Z}��uu�y�θx��Ҹ-��vB�N��1�f�)`��f��@�/�Gx�q���|�:ηY�[x�^G�J�3RX�
s�_QqH�խ�T/#��إ�SY�fe�ab�>2�F��òs� ��Ne��&E���n9�i�xc�F�6^ܐ��͖L9�6e��P��H���	 �ƛ{�9(�j9��y�fԕ�
�pc6�,.˔�����)7b��ճn6nУ����l��6�pJ�6!�i�Ҍ��vJ�2V���1qNA��#�L�6*%N�s�7�L��d��vT:f��t�n����.�n��'"�c�$��jk\te�Ie�a���ġR��E{gb�����nw��Y���5#y�M<�ܾV�0��we�����f�6wA�	ˮV�u����YW�����f��n�QfƘ�X��t�֜�A�fA%`+]�X�Ol�L�	4���[�BK3 ��93��hd*���r�=�2F(B�y'#���Il��������!�"���f�{���S�	��5%�擕z���S�I$�I$�9%��-����{8�'���H��/�oH��ʒ�]��e٭�C����PI�z�_�E���Ӫ�m��_����������{��?ϭ��~3��oo�P��_�k_^y����Ͽ�����؇��QR���.Pq��g�#�^������ow�T�gr����1�g*e`��Z$Wd����$��\H�s2d<�Mbک�h=�6(��_M�56��Q'�K���m�rG{��+�@�&+��G$F�[���H�vVd�3��\�oN��t��(M�HM�#gz'� �국g:b��[RĊ���X~
eCG�y%�J�}��S��u^a!4���D�f[��q��Udɢd��a�Zb�[�e����W�Oh�)�N�g#M�6��m��*��1�2��`�Ž(B����3�%�=���d���f���,��uH�0������N���86�譻jh���GBԥ�F�����M�xε��YYO.Ы�Gs���v7
�a
&���m�G��*/�_WU
���TW�����wSV�&��0���'s��;�[�S� �Q�v䫖��v��	�燁p�ܒ)RI$�˒L��$�$���I�I$���HR��l�6qd]�m�i��)��D��r,)�K$u��ʦ8���δP;�o0�t�r��i��k.;9���U�ٳs����X������_Wd$9:t�ogʌ�Tv��f\J9����wC9�g.�iU�u�P�j]�+*q��l02�L�dOr;�	{�Q`�5y�M��P��L�B 깚{8�wGeG�n�Ѷ/*=d���X�ˉ9ޥ����su�/1eK�Z�Y��8�~嘁"��4�zsbfY&�ZrU��<�,��1أnhDj�M����	��"�U��^�����{�Ŕ+n]�.й���%�B�<v��-��:V^]��9�x�<v�u�r`3��w��VʷF��k�5��W%�}]go3��csU:t��GNk����^�+*���k�V�b:7,J嘪��]hk^o
n�.��;x,��E$�$�$�����I�I$��$�I.�Y��P�s룠��EcJ̖�VܬI-�mɥ#�%n���,�TP-D�b�"�Sn��G[��92*Г�10��YW�$�Js��ƙ��
yГ[8��n��#dj�o��6�D��wV�0a���+y7dݘ�v��Nf%���MmT�U���wt%fm12��f�D��ru�ђL�F��l��t��˭��Bf7�{���sJ����n�۹4�rgUA3�j�Ѯ��S�uPZW��E
+,��Dr��{Z89̈́]��7�w��5�Ax�@[V�Ƕ��8ȑ7y�<Vl�̃j��y�H���8�
T1e̼�`��|��˗rÝ�N*����b�S�(¤$[C�����9�q�Nٺ!����B-�S8��@�xι��*Xł5v��܄��i����4�}�)o��0ְį���3Q�7��P�[�9ۆ�gVCI����[l^�<sJ0b�5e�s�siʹ�U@0,�j��3M�v�QZъK&L�+/��M��XMi�:�ڨV�,�Y�7Cy+Kx⫴��*��c���ah鸪>�����:����"^�3��d�g+e�zG:ۗ���;n�`�3M�ťn&n�>a���;�����/�:���W���]�_*��N�3C8�tD��A���Vnp1�1X�h���Ň��!Z2��0�������R����Σ*2��*�eo qj��L�p`v�8%ʻ5��O-�*���=ŁW)�U7��Y�9�.6��U�!]��ȴ����n�i�F�?`�D�����)�1��v���+�����f�޺J��dj�#�|��ʶ;4��3�踓����p�Z�
��$�&)�dJ�Ҹ�]w���NP�����P�;vȆ�q��{
��-ep���u�]�t���@E@�*��a��p-*fs_f�����K��L��,�z��icEu0��:�����@��1���z�KQ���ä�%n�6뫅������wg�Y3�[|vE6����׷���ln����!S7Ŕk9g�X�r��9�����&Q��k[{-�}�ݨ� �g�;��l�|����xF���싘����Hi���������m�TU&Ҹ��\��%�q���݇p������C�)�kS��QTa$-���՗ϴ��� bSf��1>���W�,�YF�7%,Ő���=�hT6�}���k�G'Lը4+�ht�^��%�t.`�6�00��Kn�dJ���+�.�Ǵ��l�E�]\��1Vt`��YM��7��Z
A�[���mY�+	��2r�\�[���_pܠY<��Pr���ɑ��JPX�u&}����d���䕖B�P[z�����q9�����x�a�XC�Bě�̱;Yb�S���Lɔ����N�b=����UZ	Z�j]N��
�Y�7o7��]o�|��,����9Dy�E�d�ظ�Z�.�*]�CCG+��ʲ���Ca�IP�z#�.n�HV�1vF5��ٷ|�u{�U�:hҀ�ݘ����|x�������F�zWU�5�<|#�J��ɓ��`b �o�f�ʚo/�̧��m�>���WL�v2�;��C��w�a���3�J/��(�v�|��w��1Y��c8���Ƚ<�ٵ����U���GTa#B�f��VфJˤ�7lfaղKͻ��
xh����gVM�`���]�,]y6P�uCy�
%4����>����|�SL�R��vڗ��w�`�f0�jlH��j#DZ �����ۣ����{b/U�ͼ�v�#m�����37�D��8(�z��ޥKG���h�ӓ�=n���4�d�pJ�M\���[!�Vv�dX����NY��x��v�Sp,M��@���ܔ�C����(.��.��5�yJ�'���8��qT��-�Z{�s�_m�DQ����h�w�����Q(��|�]��)����ڡǴ�u��[F���T��n�D��;�Uȣ����Tἶ�̔���EC	��R���T��>O�Y��*�%����������;A�r#�o:=�n˜�&�n�iX9�N��Fʦ�&q��0\To�k�#���5�;
����SD�9Z �F`�z�ΑN��mMk���O\��"�P�b�|��)�x3.ƺ������Aq�j^}�[�z��Uj�)��;���⪩!P�wFc՚��h�X� �wv�x�*�Noq����I����v���,��ӫ; �z��S�C����w^mh姷I���B*�v�nh�2[r��P�I�����ufX�������Zgۖ�fZ���n��<����=�v�U��q�x��ժ����l���5Q�%�{q������3^�C�f,5�A�����{/�mXW���)�9U��tm�&�n@�X��[oQ�0f�yWn�_ ��fkJ��K�p�è��E2Y洧���y*�p��g�M�l�n��7��F��Q�ݲ��,%�ں�.fO��bs'f��nWK�:���^�T�Ծ���'R���e�ΈsL�b���^���I�+���m��b�M:�h�2:ʖV�J�#\&����U!��dʚ��)�uc���De-�c��֚��L��_	�.�ͻ�[��]MM�Ε)�t���)2&������.�uZ%��KR�"����\��p����DU1��Y��4I�Ɨ۽����F�&;���S,�N�MYG�x�Vw(0�G	�f噐�3��)�}�kѬ��h��T��
��u����D���Ӈs :p��u��Y����s�{t�s�&�(�3k�;gd=�{r�n�����x��F���#���K��M..6�H��^j����f�E�Gs� ��]��J��X=$�6��л�F�Ø�\��kޒ��,	M�K*S�*��'Z�F�z�:6�s��}F�gC��C�+&c醥;y8=�c^wM�ɢ��M��L�LŤ�:�8�6�S��Z�е	X�j4n	wʺ�N�p��!�ݞ����ՌY�y��)��(�����Ǚ��"���H��n����2��A���n�0���ʬ0LB�+FU�hg�b�ܡI�ƫ!.�cl�#����'�G�����c������1�^N�1��?V�f������Z0G��ڶ�:n�2�5bs+�	�' X���N����G9Ttn��.=`I�ֵ�ɻR>j �#9by/w�V�ǘK�y]&���+�Uhe��f��N5�i�r���d$4w7H��2փ ���$�6k- ��֡���%�J�Fuv��ΰɲ����`������@�EG��̰���b������]��igu��7��dѮ6����[��gP�3U|��z�Q��FI��J�I�fYO7'���J*���� ��ﬀ����u�S��}5�E��x�3r�[���<�M��4��/Ε��Z`�h=A�5�vB#Bւ�S�`�]j�22�����\6ܗd��fln�G6+��y�Wa��b���o	�6.��_ov�"�ɑ+�Mۘ�W���M�W�橤S\noG����]�v�`\�����*�$w����ť�va�-iuׇuV���4�sB�c�R��V�N9r@�)k�Fs��3v�C�״Z\={��)C4�g7��a)H���wdx���GMW��Br9�R-�9��h�d۫���ݹ�d��~��0c*�VV]���Mi��Y��p�E�+� m�2����e��T��Z����	͗p;[:�m �����4�!�r��D� IYf�&�Ցy��gjVst��J�[�72<�:��p&�s���kʫ��N6�B�$������O�GW��3U�K�2D�'.�S%����=���c8�aaR�kZ���ސ�ɑ��iy�2����~������i$B�3�PWԊ�������Js핤���F%��[ҙc8��c9�י���
dj/P�TrlD�l�;1�G%����l�)|�p�M�rc-"��ka3��;�귵��E�F�V��#�Zן)������h�˪�N3�fp�cjT�sY�x��;+���A�JI�1E���f"��m!i���PK�����>�>Ej�-V�T*HKX(��Mb��<+]�w��/e��W����7Q* �%u���jXMD�o��p=J��_S�;���U~�|ȏ�96�&����������5JƦt��&uh�k:ȅ��P.� �#�7J��A8�J,Vj7��j���[���|��OB�n�F���k�ڞ�m��W��n���L��UM�����ocy�E�P�#x7Y���A�MpjҦ:��x�Xz�V���j��+c�� ��<Zo�WciWY7�I)W��"ӋboM�A.g�޹ڴr���ތP9^��.�)q��K�3��1���9+��踲C�}=�Y��V�� F�Bx���ԧ��W->u[؅Jz�m���9��˭�6��U���gg}�,�C#Sz��o(8���]�$�d��Q���)�(=��uX#�)��R���_8{n�T�GH�M��.��pkeβ6�D�d����u�W�tћ�Ĺ5��;��������ȐvBtc�ܣ��k�q������33�uhv�y��l���;��"1���e)E�v}�10��N(�L
��yƓp���<g(Z�$M�iȋ����19���
h6�V�}O�f����J�/ �})�+�4k4<lZ�8կ���<���`�]��]�߷���˪q�3F3�`��d3s��7�`�W���Ԍ���������3���~\�>��4^�вn��Slښ�������O��ݑ3�[x�Gs�.\[��%�(VMnA�o;W#o˼|�=����1X:͕��B����;-��_��{���9&��E$p;=S�Nv�7��5�5�oʥ�f�uw�[g���f�Ɇ��y2\�^�L3yG���z� ��qg@�˸��D_.Sr�ɪ�oJK�f�m�`ZO:~�k�l��ܨ��~~%��P*�����ng �f)[2$wBo24�:]7���i�!��z4b��N�uiȴNĥ\�q!��p���|T:�q��	��c������uQ�L������T|喊ֲ�^�9�z3m�@�ȁʹ]z�M\�z�������4�{�܋{Zx`9	칗��:�N��	D��o$�Ad�W7�(C���QW�yU4�n6�';���X�Pzz
�f�Y�@�d4jm����lOR���E�:����G;��Rr���{L�R�c�[2�����g����ѧ�'�����U��/c;���9��k����TqMkOFeߚ�C����L�Y��Ň7e�ȼ��%";N5Ĭ�.��)���%=����2IX�2K�o��o+�a�B��A����X�e$�3&e�a��vɰ޾��e���U�� x34��z��������^�͸A\A�ݾ|y�/�Z�6g��\�ACt#��mN�����tiq��Q��u�2�9�����"�l㪋�3m_��ΰ�#:%�\r�����Î�r���Jz�O4�O[��9J�2�r��~q�.��W����C�SV(pS���x�]�����a�@W����&��	��z��3̛�S��|@;�sj�� ���r]�uk}:�}w ׃C�^=��Ʒ9��t���'���)VՅp�\�CJʙx�|��2�mKt2"�;�X�m�U��Kx�
�ɧ���u�VW�]7n�p}>����#m�u͎Pj¦)�[)\��3j���4Mhw}��X��+!��P��ՠN����Y)��)B�(%݉@I�Y�&���A�j��7d����hW��e'}j�)Ê�(��295�<\�羮ӎv�־{�i�}��������~�޻��3>�y�IH����':��f�E�aŨ����}���Pa��W}��bF�qyСmk8�V�Q�ʘ"9��7$�q�ֲz�<:
{q���Z�E���eK�]�<�INq"�1�;8� v��Þb�m��x3�j�����^wE��$<�7}�y�6�V�e`���Q� ���'�pw���c�y~n����R�H���GV���S��D���kX{�Y�m�iۣ�ＲJ*�Ǻ�u��w����$U��+�����9��h:��1���I�{+�܊5�*8���e�J�4�>�Z\bgCw�o��&)nLCu���}xx��aj~(c,��'t�i:����f����U�^���-�s��6!;�5�(;!ɗ�V������B�� �Gd��>�gs����R�s�	,��}�U;*r�Z���=�a���7��V�+Ρcud0D�Ga0#3����:���G�Ϋ�r�ե-�Q���iVh��9�ޑ�p�ը5�v5ݎ<�OM��0���
���H���h86c+��HqșԈ>�W\[�����h�YKc�4-�)T�~�:�|�`ok������Q�W�b�������[qC�Y��-�&*��J�Yg�f^S�e� �Bi�KHr���z��=�@�I���O���N2V#�܋\s� ���':�{"�\�4�:_�q�\3c���/�9�1����$��Ӡf`R�OY����gn�L։|�;���ș��+i�����T�[A��ᆵ���r@0��aʼ�P�Rb�B��O�d��۱���]=�R�әh�9��fJ���"�>����{���	�i�ٌKx��0\��_��ж�ځf�O���ݖy��';`Sb��Wfyt�B�� �i
�%�SW�x�E�!����?�g��7!ŝN����gXɆf�Nu�[y!����*�/g.d�A�Mm��+S�mN���HCr>�މ�8���a;6:��z刐4A��[��&�5f��f�/5���o�_Nʥ�K�st-���ny���,����P�1K�|60)�|ɰ��>�53�V���1���U<���|��oN���`4�j�sѓ�����,t�OsM�P����3��e�vhHF1}��ıKYv]��|���Ά�cF̈�4ú��T�Y����N�2�b�B�X��*X4��f�=W��d��l�͚F��11I�`ۮ"�5j]'�v{S�5�'e��
�o3/JWLb m�,�Z"�sU�D뛓*�����-���ko˃�Gkb�m��q�Z^H�h��n�%w����@&�U�.k�i�n����XZO���juzZ�S|��-'Xg���]���p`Q��c;d8w�Y\*�pO)� �8��&򫌹I�Ȱ�?[��_�Շ��\�CM���ycc�
�o�b_gT �9���f��j�)R�7����D��y*�7��;�#��ơl���!9�b�����lʵB���Ύ�����E���Jsq�$���yq�Q����&1M�ń�X�3X��:'c'	�k[�l��d��@�A��!\�,y��W�ο��t�.Ų�ti�T��]'�5�k��A���s�.��UX��m��\���9]��=U��q�i�+a'4\cuW؜O�iq����q�o\��۵Z�h90e��=�+V�!���=I��k�4��N�=�6��n7�5�|Q�u<s��.N���s1(�����-Ϗ�Iu�3�5�Gm��hR�<��U��M.�iܹu�bm�8��'g(��
�"v�sNPX�!�w����.�oWr���;�e�;�G1a�$��o(���ڛͮ���A��(�w�VMj�n��G�]{�[7)�%�$�3Br�˗ǜ�]a�VRo6����Z��B7����K���3�k�iŌ�F[!�=,�R(�M��<މ}��hM���S��t�R�i�at�62��ͪ8�ɷ]�
m�,GN�7��Q���N+oZnԨ�ݝ����_���5!b���o`+ 6�$Hf�l^~���}Β���'3w�������;�Jk���k��fIZ'h'�WQr��:v�pcR����+�����S�r��ھshH� �2���2g��X�����*ے�AؕYO*�G��&"��SH�ƪ����ys�WCV��"�3�ܸ�m_B�0������l�NnIgu�=hd>���h�,�k4�WU��i�]�&ma9��������r3�I�<�s�tΚ�]�ur��T��y���muňvhA�d:��vJ�t�Ho�����5�B��
���n�n�q}o�m����ԭd'���Tq��c7d`�R�"C$���}}AW|�f^KGW:��N�Pv4�Ra����B�fw,��Ҽ�)�42��Nz�p�ܗ���r]�`Z�Dl�9{[�+fe�ʶ�T���pM�e�m��u{Y��|?�T�@�A�JM��[J��
M��_�	�)|��\w���߿���4+��8#m	X�Fũ0�N�d������[>�-߿�߿2~u�Ue�g9|�8\8w�yAs�1�A�*�HN�B��M��ME����t;z|���X�O�5�
���i(���[��DDa��2��o�.Y��'��uRM%�FI�V�YוB�d[�XP��O/��J����u�@�u�z!UU[�a��w��1+z�X#Lĥg�<���4�)�6�鷶$\�=���v�25���,�W�6���?��g�����*ǧ�4��'%��t
b�cT
��ۦI��R;�\C��&�\��/1q��խ�>@Զm�x{$id9X�����fR����͜�(>MA��/j*/r��e�N�^�m�������k����dp�Փ��n�����k*
���{�/��t��`���#�;�%%c �;H\Q�8>����Y������9�r��1�2���.��>:O��r���/�n��0덡��۞0��1חS�������2b�+(�6U�؛�K�v��	qj&�u|>>{w�:���t��Ǵ�2��[�<�՟ (彏�9��Tv$��W�U�~��q�߱��#��N��k" ������ߪM��/]^�Vx�q�?
��-��wyE�70�/���ȅ�Sʍ���\ad�]��I�"b���=�%��[�f�����|�u����k8�C�63Z���9\�5;km�v'Yۛ��H�N���T��u�}�����^]Ğ6#~Ψ�H�d`ń��L��yg�	�����/���6�p�]�þ�)�B���S�79��{�~��*�_4��B߲8�U����Sm@u�\1��l]�y�]��Ƀ= �Nv�YV{?a����/1�+�T��Η� P���Y�������0�9Pa�E2�ϰ����W����X�El2����ɊYQZyM�@N�O3��W��-�"�uxl�/��C�-m'��H%�jK�Y.�o
�L��q+S�ILi���b1��0����ٷ8{
R�'q�K�5�X�?\ڈƖ�Ђ~B�	���N��2e�,�Z)V�f]�7�S�$�ܷ<>ߩ�`���p�z�e��o�Q�e�;K����>��t�7G�no#�j$_�mk�ٝE�-Z,�Q��[���g�ꚍ3����¾��q\��ԫ�FD�#9]�6�դ1�8�$>?I2����U����Ҷl������ W
LFw�>H��w�;Ղ�����s���umK�Uŭ�|���El ;�%*T��$�C3ѓ��p^�X��<�Z�cxxpٵ4����ٺ�ջ���S5B��Vf��pT��:�9�x;w�q|���gљ�Z���	��b�x���_8�sX۔�e�3&R�9P��)8���i����?O\A�aBb"x���%b���A-P�ͷ44e��Dt���Y�>?.(��;��;��t���p������ۻ������.ŹFě}�p"+��[Ϳ ��.�f�h��،X���$��7�1����$d�]��$g>?)�oi�S&;d*�9�	�����n�����S���+#=�/����#�W7�E��
tV= ����J����!|@թjZ+�P��j�9��{�Lg����y<�K@ozD1�zf�����^�C��� �5pȴc���������7�;�yè�b!�Rn+�����1��S�NN�q�;/�q|�@n��/�o�W{��òb��_g7�_���NN�4���%un�Dp�����
�n�E]�I�����|���q�dÚ��n_z�Wr8�N�1Sbc��C�`�K�ޏDR�CﾌL{���;��.yB�!j�C��hM�5-�\��P<��4!��y�o�Ȼ��fjw:��nU��뜞����"�����\�%CȎ 9�b
��BB�iR٠�)ȹ;@�!!g��\����0ǝ���k��1:r����G�P_"�]�y3k�R٥�D�)�Z!�����/�ȭ�A��w��癶��;�tj��5�7��95�M�<��+��]E�VU#�&��nR<�X�7 7��s�[�8V/�w�vtS���"��qyF)N@u��D<����"ܷ,	�nԎ��*�E7|��[8�{��Z�P�D:U"b<����`�"�|�r/`�uJ��`���'���u"��$�_x��n��ݱ�g�ដj7�QND�P��Z�0w"nf��و�
���/�ȍ�W�Q� <�^׷��v�λ�WE�1��@���J��T� S�PwqŊ�oI�P^F��;�)�P4ڔ�F������+Wּ�y^���<��/"��_ wx��ḕ����.�QD-����$�R����n��s��t� ���NZQȏ��HZ)��)�E��T�լ�
��7��!���^E����E>���X���Wٟ{�����$���q;}�QJ\���R;����H�2��!�k?�r#���#<z�uf� ��.4�����mN�՛%YS�o�K�E��"$+:�w�;�rx�Ғn)lP��X�/�\Ƣ&�H�r:��Z��]A��e�nPȾ����{���g�.����hE/LA
�Ȧ�^EjqK�A7�i ��n ��_����W�������T�s��|�X���.r��R��<��'b���qBD��Ej�@N��NE���7o	7�y~y����R���Y-�G�����*U��;�j��Sw1avb�3����wA��};x�p������TS�/Qs /qzg��R���]��iN�/T!�v�	�����iqȧ13�-�η�y���P���[�������RE��V�]yB� �(|� /�CN�!P�iR���F�^wU���;n�r��b��������d�E��Gkp^ŸAO'1B����mz�C|�|�\�{���כ�r>8�1������M��*9����+���v^#�)_&���.���T�~g��3�V���B�#�[D,���#h)�ԛ��TC�;�ؼ���"�����M�5��^O �|޳�s}�Q*�Ȥ� �hM@�B�Qȭ@�/z[Au/jO"�)~ҞE���9�;�Y�;��U7��Hc�CZkEEcmC�q�>�.�f\�ӽ��p�Uɴ������ع4�:BŭU�4��l�����wf��G�k��*ìB(�?Lzf=�o;����t&`�ǔ��;I"���J��<�PM��T�"+�;�(7�	Ƚ��H��'1����mY�����Ssɨ/"��!��e��už�SUJT�3gp* v����j�"y^�;�y廫O/���|�����uKK�$��ڐ��h��)u�y1*-���7zT��Y������E�<��i�_^k���/!�L�y�S1L��_'`TT��y�iA��\:��P��d$GU�[�g8��>w���Qq�R>E̴/zG�b��^��L�s��v��+�7@��� �\쾫���y�c{�l�`��5��,��x���S��y2ڂ�^@�)��^Aj5��T�<�r	���jn�ǜ�'� b �%���l^"\�,���a{1�j��/�)���I�!؅��1^D	]�<��<�{�y���P�(�D�iE��ȝ�m��E�1e�P�R9�X*�q[���J��`;�~�����ڼޯ^g�ߛ򺍢���"t� �N�)c���yWȵ�[^E��d����������+�_��[Y�y�5����LѨ^_�05��f�;�R����P��<����\k�T�J����,v�j�V��ةp5�Z=�s_e7]Ց�98�4�����KQԤ{L�cԯw�5�*�>wm��\�7ŨY{$�7lLW�?k�tj6�Zl+��R��~�L�DD3���}�$�w�"���5�[��QK��uq/�<����S�^E*����A�;5�I*�}���1�ke�GqE���e1A$|���V�Ճ�B��7�T1�O"k�r r&�ؽ�#}�]���*����t�{�^�y.Z�T�L >�z��CU@���y�ND$B�3Ⱥ��4!�Nk��^s�c~w��q^D"61]��j.9J�n�PI��Л��B�\��/a�Ц�I�;�D3�'-�[��g�����R�u7E9�7;�ɘ��⼋�P�.ccw���C"��F���Ȅ��.��g���֭�y�O�� �Rb/�K��/& a�
Z���.[���t�aȷ7C"j�R�6sF�T ����mէ&�3�s�����_"j=�`a����R�b&�Hr#g4ry/j]C�!����(n5z�;�Lc��g�T��dBA��;��f�	�mz%Ey@{�ug�/&�d�
S�|�� �iu�yc���|�<P3���쩹�5q���#ؾKKޑ��(;7�KGq_"k��]K��-3~�ߝ�����f)��t�r-�H�n^�P���TNr��K���T���*`��ف�7U!t�pz5��n���\�l�3A��w鲫5Wy�:�o&��O-M�q���,n7�wg9TEt�2BRs��R�G�>�zg��3���Q�RNʨYAi�YN��Үd��=��u�AP/����1�@?�͝��9�
��rn���Zw7'F��^�}7�8���-3�¤������p����:u�#��Ӡ���+7�I[8�T�z�r�g���iVk(��sW�=�G��r�M�RD�=I,��h��(+���YY:m�	;7*��ʡ�	f	?*�q���[{�n\�59�	�/{_�U�������C��ө&��/l4�Tp��D^��� �*�)�;:㧍G��T9y�By�[�]���6vA��̾����5sפ�ƟOE�*���z�~����~����D8y��J���J}�E`nu��֔�E�f��o��،�r��y�z�o���F��*�̒�5r����)�즍@���eA�E�8�F�傗.mf�ݝ���x�P��6(��nP�Q��}���Q�Ԧ�1�n�j+4���>�9T��Q�e��L%�3��rj���	�`��p?W!�U��o�frN*��Z	�����f�
��i���_�]�V���[���p�vCsl�����;غZNY6s�F:<M8|��>L`���oy��	����ެ��^��y�7䷗��۳�
�Go��}��٧�D�X\�em~!��כ]�C�t��C!0��y���-�{

��V�ǀ�t7�-��k�b b̸�뙴zE�8gMڝ{�~iL��0�ۼ,�Wgf[\Eq�2�cwnjj�va��3��t�nt�/t����Ë�Y���xȚM�%h���/�K��:�[��]�N������8�\)�v������ǒ���8pTY�ݟ��.���M��M w)����Mq��l�	�yM�-��f>�̈�U�V^ѳs��T�ɺ���8�5�.���nen��)�]�v�u^:��j�{�զ$�ܕ(=Ρ�'1t�+);�	'N�Z�m���Y!̣�J��	5�v4�'�%��,=��l��Ә��'ʼh�nQ��njv�4̹�E������Yu`�"�.듪�)K4A�ۭ��p��.�d�K���
��l*�5t���m�5ܦt���¢�۸_f���bG�c�����Z�V�{j������"�Z�0��$��y���(�^�О6q����m���D(0�-��uJ�D�Bi�M%u-�;�a¶#���6c��.j9�&C2���l�}YoU�h�g/GS&b3w�Nʸ��,��9н�� �8&�\���sl�dlIֲ��K��ZS��YR��D��U��qb��H���n.{�9>4k��YXU�V.Rl�Ҍ����c�t[;��lՅ��bN���0Kw!ě.�JB��(b!`Zs��3`PV��M�-\��neY��7ǖ���$��E���7;��G��+	7���<ˤ�wv�Ζ�Vi�ZJU	v-拤��ɝ����FWaq�����]�y&T��-Ӹ��y��
m1J�VL�6w���)Nf�h�K:��)\D�+�7��Ca�إIiJ�^Xݾ�Ǧ�«,�O��9�E!�LsI=����?�������Z���֡s��^L�յ�U��VI����}��ѓ&r��2�X�s���f�y�51S7����[�R��~������d���>AQL�i(����yA|�+,�d��F���QFP�˝�'��'afRF`jA��� �(��Z�j҃���*9��n3���4���l�j���3m��j3٩u"e�ٕmE�7��dM��ض���GNg%T��18���2I��FХ���$��>|cV�}Ʉ�b��i��hʪ����M�+�f�l��Q���v�j���z����ًЋn����S,����c6vTmM�-�BK��k����yv�?R��TqE^�ؑÐ�s���^��q�Y7�5�V5\���k<���U��1��{�W��uc9߷��w�^�P~�0��"k뫯����con3��G)�t��zW �M�&�o�o9��P�۠�N�e�b=7t�E��$�Iv1����T|���̍-ܾ�y�Fn7�Znr��(��`�cG��_����W&vN��|>Uz�bז����dT�����3_K�d&�߭����zc۲��^�M[5=0�?z�T�������Q�L��I���ä�ca�%ܗWn��m�3B	� ���ʲ[���頪���w�[�����/��s~�6�h��R�ܻ�6���#2uY!XQu^ǆ�+l��E����NK�Og*=5ݪ��O���F�O���wk�X��:�{X�Ú����{���=D��ֵ�;��s젷�~���\E^[T;wI��>�F��W��$?�ʠQ����:�΋�ڇR���,��׊�"�/^�T�F}�Dj�鉷�l`�+�T|&�؊�2x�H*�p|�4��D���"���)A�c��I�i@�jF6U��B���x�r�J2�\����S���);W�<�4��,�_ ;޹��x�7�9�٪��@�^؊e[������F?'��K���u�T�;ӻ�g޳ۢ��3Ƈk9�tn��x
^g�$&/m���·)S���]� �(���JϺ�ߴr5���[��i�������o��Ą���d��EFf���jGf�S��n,�;\9�Bɨ��W��(H��/���J���Z�r������O��.�g_rc'�8��Q�v\��$ӓm^�����5%�d�ai��7j�c`�V��{�O����k��_zi����
�����"�8H�z�(Y� ��\!\<���[G�e:���ζ{���l�����<��a2,)۴L8�sH�&-Ƚ�5���ޣ^��[l���!����]�;{q�^bw�O<"搜^0[��me�n�q�h�U������*r�D�+_t@�pTׯȅ:�<:刑*	ۍ�#77l�VfQsJ�;d�QE�q�F�-�#B���or��stY��ya�w\n(,f6
��|�N�ۉ8��|�/�s<�9� �d@�w���;ڣ��\%\^>b�yyQ�*\j�P�c�m$ڑ���	�m����ꉭ���U�/�*��iF.���L��˰�c�ݖ�.;� �V2�Ҟ��������M��0�V�w#���O2O��3�y�X��d{�s֏���8Ū��dT�Ro~\�)y�Y�+[�H��s0��kj���*N�������"~W��P:fX���HρM�Q�Y��UׅH8�7�� uz[c�-D�o�je��Ov���J��;�u�*n�L�Afu[�0�*VQq�X9_Qt�9�j*Rkm���˓�6�ʎSʴ��)��J�h���Z�r����o��o9�7[�,�@=Db<�x"����˸y9��U5d�]�b�q�b`P����M�
ܑ�^���>ۉ�nkΡb�(�mlM^�a�D8hM�g1Ti݀��=�
D��-�]=��^���V)�ycke�3�AEg�|�>hY��wsk���o���JUx/
���t�S��1����ҫ�Gq]*�6�:X/�%�j$������,\Ĳ���\ӹ�V�:P�N���g��]i���^�c b��WN�c�[����y���q����3�&��vf��A5���x��}�O��D�MQ���k�z���U��s��'un�B�mczv'c�	�i-�@q�4�+L����}_}����D�{��D>��/郗���[##R�z��=v��@�e�-��0͝�m��[R���U��SI���.��J��3f6�5�4��B��h���c�}Q�2!���"��vw�J�6V�{�\�Y�)�H��Y�[�]m���^���ί9b���^S�8���!�^mA�t��Nso�����S�qLF"=�8�\nE�]^��:�{^���-�8����&�R��<�����	�2���<�����b&)c�1Xj�^g/���\���TL���h�*���x��Y�MNϔ�-篫fp��m��@�u=�i�=0gL����x_>!k����Y���^��fs��<p����>� ����3����ߣ��8�7�2���
��ά�m�^���U5��`pF�j��B�ri���̍>:��*�K`�c��������-��s���ڍ�X�@����",��b*w[}�Cq��%rڀpo#+k�2�B�	*������1+mɼz�tTL�����:;Cj�ahu��2]Q8�`Su[��Z��u���OJ \�B��H.���w'f��$q� ��L"xP�#��C�5E����tz�b��� �Ue
�I���qn$��r�-����c:�^if�Ls�w1?�V����|�Ζ!�u�(�;re_p�s����6��H�bPF%�p�}f�;��H!��_���>�zf"=�yvi�'G5�!��w�oߏ,�h��.�� �)k�!�솹���f+x�A��8�RԳ�j�e��q�1Hn-�T�z��7X���A����"A)����w"���Y�{B\��t+y�eOo��2�Jh�HB�o��NZ�w�	�c��������b:XgK����5���,w�m_���k�	*2�}�N�_�L���{o����Ҟ���U/�_+Z�q��)]�>�'fK�+2ZӸ�5����h�9`����t���}���u��眚׵�&�/��6e����&(��ҨH���*\��X�C��2j�����,Ed&���q�wЪ��sT�7�3����o��z�����ֱ����u�N�4+L�"��")v�I��g�D'y������c�s]ZVvTL�a-��q<��h�����ߊ��9��PrW���L]�Qff�La ��"���4��[O/�m�8��jؿ<��+�<�,��ܶM���Ec݀��c#�qȽ�vy�/\	�n3��x�qx���^���ߴ
�V�K���a,̟rX�z����=(8��oʷ�w���Ko�?[�������у9Q�����d�7�ڮiU��e6�����+j$h��B�e��B�o**�,�8�!{�Or*�T#1M*��c��I9Άhx���8����b^r�W>cV��~k��ky�5ɾsС�
�
�s{����݅�ے-�DH
���a�����/�;Z���~iNԊŋ��eB3=�K��w�tE�����T����#U(�68Vog_q?Ͼ���8��գl�=c�pK��(��L��Tu���.F߂�ch����0�>�ɗ�>5,|<�Sw�j/+y[R�à�FU�@����ڭ��EĵTm�1���'/{1pj��q��u�ה��EU�OL��z������@����1ءP�+�x��E���"5"�`���q�����u4|r�����uod���ଈ�d��sZ�N�OM�6)����{|oh�����gR� 0��K����N[Vn���#h��+����°�x,h�ȟ�p)�ԭ��R�R�.�-Lr����i�>���4��zO]�Eu�ѻ�"4���ɸ_)���OXʹ�uS��͇{K��0==�ڨ#�V��&�#���ڭd|��B�J��Ż�y��f��m�A�Hkն�]��M:n`G{����aoB�("4��CՔ�IG;��|gf��Xa<�<���UZ�/�UQ���mbł5�VY��`p�k�)��\�NՂ�pH*���>�w�h��&�iJ
�I��';jη݁���)^m*��[4�Xj�1b��`G(���'s;������+1nG�M�綯����&�c@�ڹ��*Q�)(&^���y��Wۼ��I޵!��nZ.gs��β^h�f�e��bu&L���{�;U���e�k��;��q�Mv�;E������JL��c�
U&�E�}��X%5�X!S�rG�-n���\�v:&�4�z0Џv�m���aQ7ա��tNΙ�Y��NfJ�6P�h�)tM�n[|��3�\��i���1��k��|i�5��v�f���g�!��������J�w �S�G�d�6t���=�.���O�γ>`�w݋#��C2q��GWA���+�,�aY)C��[�~�ӨV�3G)͋��ӪZ�9n=��\��F\��{̤Ni�h��wo �KTL�RkZ���z����"�R��5��mKk����{;��ܽ ܍'+'����4���t:ڽ왕�iof�ܻykF�+�Nxm�j���!��5�$��WVz��.B]�EP���υ�t�CeTQ[��I�{����:@Հ.��bIl&4O����sN�Mom�Rۿ����_�G�&צ��Z�]^s�ѽ
,^߸��\b�Y����~�����Y�f-�}:�m�ڽM���])�!��|�鐧��4�s9�dd��k��>Q���b��ݎ��fZK"D"RJ^E��˜2RO�����I��#��4u�����M�<��JL�l����(��ce̔�F��t�D�Yi��jfڗZ2���tZə��lB�8��|<�uw؟'EvÜOn�Z$�K���Sanx�����Y�;��R2TK������g�;�sk�ᾍAgM�}\v7��ՠ�5��g^�δ��G ����{���b#���i��gO�f��t������5$�ǹ�Mნ�.֡���ip�ٓ�8�M��]�
��Nt�#oN�
���fp6Ҭ�v��mZ�֯���_v���1��\�Jhc������)��	!C��d"�C�Ԗ��������[c#�����5�x<zm�-� lƊЭ���tG"_�r݃w�C	y���5va��������Nk��p�orwDiY�6�FQ��S�nꑮ���K�2��;�Q�~�F�\:�[������pʲ��i��%Y;si�t�N�j�����'�or+X�9jN�ݫT�
}(�:����q�f�͸��H�/%���˜w�s�)�2(�W�ߛ�|�5�s5�~Q�*��.���U��s�<sm��-�����:樤V�P.f�tV�³�,�g&�������0��p���!cGD�Û�?_*�*��c�N$�8+�j�Z,�כ�p�^�֎9/d�ܚ����e,͑�2�A9[�����}�^�5{w�e���
��:�R�"n!W�/��q�h���"dUOe��ڣ��
N���΍ALm���w�D=Hˌ���w+���z����lG$�ֽ��c���������!�-Sy0�`�&��>�_qov��с�i���x��R��E�����0�*��Rm�,efdT�9;D��wq8�:�÷���,V��ۛ޵�ou�zU�I8g<ֻޛ����,,����7k���ɺ�}YϘ.f�5��"B�	ؖ0������YG��G�a�Ҿv�����d����Vڽe?9��YBw�j�At���Y�\�����:��s���u�dMv�A�f0OQ�c+�R����ֻ�����2�TpW�x.�Bhuu�=\��z!m7���յJ��u�N5V��-�������Z�H�e�*U�T������s�8���얌W��+p�6x6#ǝq��4.�9>�ӢṴ�WN�.�K'*%x�ۻ��]fh��Oa��V�%�!HQ�t&����:՘���{$'��UF�,�U�Q����(�����DDϣ���D|K_W�(e�3�M�F��]�W�7 &A~�s}��h�Uz�J�=����U���
_8y9�1ZA}�n8]�%�<�Vf��8�b��Qy~�+U^�q�����q�I/�g�X��X`9�� �._x�,&�u��TX/ �1(��fy���=Wx>f��3Uzɰ�ʣ]z$lٵ�Ż']�٦��M�Ȏ�͗Ose���Ùu����A�W��Hſ
�|w�L��o�Q�`Y�:�*I+9d�Q�A�n���מ�H�u%����y�uN�]FxF��H����/���>�j�,9��Hk��o%˨u�a�f�P���ޕv��*#��N�0a����q
��k8�o���� �(-sZֹ��_��_�1�Y�wɽSۢ�w�&��o{}�X	��K���y�I�Wu�/3=�%�Lg3A��k�x�F\���BiK=��΍�:�RR�Q������7b@�r/qLV�T�<!�?���T}�W����ъ�4������;�Foi���%�f��V$�$���\o����wA�+`���@�d)DM(Ѝ��y�V4Z.���g��O_F*�g�Tq�:ګ%��w�koSz�V��|�W������ֽ�$��#�;����>�P?U�
m�vj�u�
 eef��M���0l�G-�W��2J�ی7z�)�=x���m^pի6�m�s\���s�� Ȣ/���'�2~�c�|�=��Qn�m����_W3�w�f9@�d�J��.�mg1�wԩļ⸥���9�S�ø�
���yfИ9Z�f�0AN{] ����}\�o}F�nlq���t��p�h]"n(��E`y}�%�
����,IF��]�H�s(Yc٤��4�Gy1u�����0��*�l��UN~�{�}!�,����vU�06Di6�l���X9���n��.�y����e�fi�e>���u���g�-"5�Al����J۞������PZdjv*��gl��g3���j�ҍ���V�^��7����kSp�з��e�"���e�
R�7���+�KDG�LDDL�ޏDE<_}h��Л��\qˌ2/Мc|L����&�f3�5����y̘e��M[��Ô��K��iI�D��
�15&���̪gt5cc%rg{ K�M#R�	�\�U���e�0> uj�ryB_XS���<������|�o4�kK����7BXw"EZI�񶅮w$UF�7#�s�-�F!ca*�w�����'k�T��|��Nʫ+N`��yڶGj6���E�Zx{�=h��'%E	b3��H�����p�!ڧզe�n��ӂN����or5�}YYU�)f$#��R��y���Ou�Nf����f>���+�]Ý�>n1q�����֢�F��cs|�A}@Ek�ͳ������bo�_��ꮎ�����[_vd�웰���c����aԗ�]b����Sx0wm�%0�����7q�89t�ޣ�Ϧ�u������*sJ��|�4b��QԷ�����ʢ��s����흓{[�B�(N�a�܁���yc9��]ơp̌Pt�\}[O���+ZW+
���3+��p��hJ��������Ѕ��S ��Fz��|@⚑D����1��y'G>{u�P���^�6��n���E�"��3[�b�G�P�E�]�v����l߅�;9�#��c�U�f�4�aJ��0e���7`J��,^�K���#�j�7z�1Z��~�e���
W:�3�_�c�u�(�v�&���U��.J*���w2ًI���n�5�ƹ��~�>�F@ qmk�ߝ������'���|C��ֽ�{�4q�b���ךW��ns�^xh�G���A���PKO��{ON��׬\Pb
�YOy�m�E�j$t��$���9�E�氻���\Y�������=�z�c<����R�B����z��=�J�^��U��5���!.2C��Ļ��	<s��r�l�:Ƃ�򞃨��ub�\}Ռa�J����k���Ӟ���}�,ܣg�	�$�����Ӡ�w��:f`lu���rj3bAt2��*q�g/��9O Oo�N���V�75��6�t�u�~��Do�+L�C�N�Ԉe�~�,b&���X�GW�Ӳ��o�:����<��I��1O��yY㶪xVV���,v�~`��M������-�����P�6�,����+�7-8 ����_)/���a2WegQ��0͝����:�˔\ ��ʛ��"z�2
^cY�<�j��G�z��E�}��<�@iF�k��|sފ��VcO�y�C'2q��B�חxvA�����ZB�^v���o����vwV�>�(�!x���>b챜�� h 49�&�e{�e�p���m��t��s��������K����ѣ���c���=¡>�)jNy�=��X�Y��^g��B-��.�Z�wfڞ��C_�W����w}��|V��������0H� ��)x+��c���2���Oz�4i����OE�.�8��z�e��+`�@���z���z��tI��n�������hn~L!kOe�pc�,���Mi�8z��V{��fD=�iH?��� -�<��Z{P�[F��#c^�/׾��M���wq�ħg��)�*<s�]�茣��lD�7�-{3gK���p����q�.��dV;fw:�A��Dn�j�ƶ�.󹀳"���90[�s*Z��[z4ڦ�1s��"�v�oB�%)-���N�:�_E2�زr�TLf�]*�����c��A�&�MtÕ �g��K��U����I���(�Zs�m��W&Cbl	+�eZ
��faK`��p� -r���ÂZ]ru51�MQ����RZ9Ʒnùy�o��2�VY�E���38��5[CcRS�d�K��3Y ���C��D��kvm��!>F͝��*���ﺶ�z�AQ۵�Q����ʷ����pYA��f�ĩ�	T�T�Ŵ7�<���iP.zD�{�����'8[�$ֆ��Ju���T�VqB�	��&�1��+�ݼ��b�U ]Q�Q�-����o!��[o!������Q���� �ׯ�8�ߘ����u���l��X��d����h�J$���ִ#��9��.�n�kɶ�[���	IY]��WE�sltk�d�7�,+X�b<��5�U�`��m�Ҩ�	�x�k6,7Q���-uB�T5���D���l^���{U\2�W-�:}����o��r1�ƍ�:a�����Sg%
sVE�'���t��H(;f0��fWwE�X��K����٢�uXoooz�O��&��J�.�J�axQ�ˬ�0M��[S��5"��#�^^��(�҃�X9�F�wEvY��^[��\�ν�Z�3�2�۬�;ʰ�)��e��J6f\5=�O1WB$� ��d�g[��T`�Vpݔ��$[�h�(N7��̛���K���I��qsYB��=b�t�A���Ǌ�~����"nf}>��W��,Vب1�ěY�RO��m���}�W���h��OlK��>k�Im�E}w߾�̿8�.�-��j�>N\�4�gԻgD6��$Eg5�������l*4K�{��2rn.��C�9�l[�[F�y;ﻅ>���B"���2n����e��K�ݻ��b�+�)�6a흺;��k�y���L��ϧ����[}��|��a;��Y�6��kΆ����
�d�m폾>���[�{�5n�*o"tN��t���7�����^���w"�r`E��wݑG��-�֮�"������*����S}ߩN�k<��:�v:��f59o)(�ղ���%f�+���s7�k|�G� �_1�����?�Ul�Ҙ��܀�􍨗M�uR���dqf�+���z�����GG�m����?Eo��O7^B��N�`�4�z�R���k۾*|v���dj/b'�sC�74)Q�W��=+ם�T6l��8��b����Y!ye(?���u�����u�.��>���n6n�#!ŀY_^��V�0��$O{Çok}��㨈��"�Q�桯,;�~"��⇦�2�o͹^��	<G�wp$�S"+��5��l!p���90stײ�{�Z&�:0Ĭ�����L��9���S����4�����C�~	$Ą����<>���T�0d�lA�*�� ������o�͒I�Q���BC?/�x������h��*$S��aK��v�$t�4K=�#3S��JKon<75.�`���x�Y��R�7FG@e�W�ly&l�cI����A٩C������7�g[�ů�C^�b�ɝ�cH�OQ(c0t�-,/��7_z�~�@�-LfR�qN�u9�dd]9J�o�Ɲi$��|�+�j�=�0�(�ӋK��6���#O�4�ӷ�L4������~�lU%�sq���\t�WkM��:)sR�gi1��7Gpm�v�p�+ͤ��:O������3��yx�>�e�U��^v�T�Yҭ�p]DC�(�:k�┄#ǵO<���;��|�hTK�jD�s�eYW�2�*�I	����G��o-h���^(�����%k�cN����ֳ�.��#���xo>�'����.;��j��KK��:d�����`�Aށ[]9La�_�P^:X���X�K�b�{+83�Y��ݣX
onv�*Zh̕��g��~7���e�j���ޠ�馺mse���j�z6N��m��c�I�ʾxU�1�o��o9�7[�=
z�� �뻾��ۿ#4�#I�
���;���6{�k�M��U3�{�3.����F��<` aMH�C��&>"V=�ū��[�G7��%�7ظV���a��{t,��3�Ke���`
l�}�Q�e��yV��dH"r�(߼p/"�-ML��*/�N@�/z���v�1Ja�+�ٿ�<�%E�+o�f*�t�
x�B���U�Z|l��zv 5�U�U�z���p���$hZ��T���G���J����	����quJQ�nF,��y��Ը�0JFMę���9ӥ���q"�]T�Lh�ˌ��axbZy�'><r����.uy��K^��f�&F�h!�Ì�4����A�T{{��lfV/r�)�Z赎*ԡ���[��V؇v$���M@N��,xL�9�v�<�/�q� ����u�d��G?}Tz�"��3�w~vSz��7v��k�?Â��:Q�#%%�(kr{��S�BR��_��ޠ���#O&̩DpW,Db�z���r�rc&�TlOM��y��l�?��0�k&�U���J{S���s�YgG�ډ��H��O����*�U�F4�/j0���G�����0⤸�/��)1P3�Ò�ȹ����F�\m9	�Ș3��9�:�N�-���a�G��w��a[PQ��>���\x�W�����ݖ3��M���\��L/%~3�\�o\9���9�P�����*X�m0Lmt�wR�I'�{Cc"�+�>�ii�B�u�0'�Y̝W�q,g6=h�2��%g`�HbC�����:����C3�4�kF���z-���8ϯ�Lk鹥�@eJV��uy� u�<��{�.f�4�v�iëY� ��[���<��L����Jz�H�7�X�u���8�E�[���Ђ�FΤ+��F�R��O�Q��켨
�Z��T[?D�^�w��@�,�	4<�VSc_b�s]��ok��K�ְߐ�(e�0,�;X�!f<h߶Y�����xe~5�W#Jr�aR�웸r�uW���Gn��ƴLa�t�!���V-0��G�T���|���S*�?~�����q��h�C5��Z���}�^B
�N�O'���o�}�	#�g�φF���<Z�%S�3�	���^빖\�绹�9�����G�T|Uu�&���R����I�=��Oם�^���#ðkX���8�Y��8gn V�EL*.F���_`�����LRk������~"�}������mƊ���bu�J5f�iE;�w�Њ�]���%�s%�uD�>���Eu�f�i��l9]�
9�(�T�f�nE���X_8���Q�d��e|���Ȣ_:�{Ν�=�yWj��[��
�0u���4�VR�>y^��*�ҷI���C�968����ta&��|a���]Nn_T�Wc����K��ړg܆�A"(�~Z_�heǾHχ�ҋ>��ݛ{�MG.�HxL~:E�L�i������i�۬=fd��<|�m���u�P��j��T`4��
M�Α��,m����WW�n����YV�as��3��>;���cN��X9�-ܿn�'�v��X�)��Cl�"����dZA=&��To=y��φ�v��@��Y_���PXx����k���ޝ����n{gf�u.��%qC`C����G�҄�8�ܭ��>�~D�,��m���8/D�^�.)HW���%�y�ބ�鯍>n>��!۫�]�o���V�)cm)�m����8|�>��mL���A�Pҡ���^����~�yǢs��C�FG9�=A� 3��zߝ�=7ŪU�bb�<�>8t��pdJ!��u �+\=GM=��q8G}hQ|�@z׊9^a�G��/�!�C'�²=e��^�h�K�Xs��k��L���(~�\���qQ�j��r����"w��$W��-!����c�.8Nx��Ȧ�{۾��n(G����x����|f&v�Ǎ<�<�R÷]���{�׶��<Xrڜ~V)����S^���u��W�77�Ӵ����cj�R5v�:J_T+K͉{Oy�gv��wF�%fWR�}
�. WN
*��2�Lo6����J>p�"�m��%�>>�s��\t���ɗ}z���ʬ/k")��ET}��ՊO⅝8�>^���dW���}���{��S46ǂg�Y�w"SO(Ⴘ�����I�N6�����Zoy�x����cF߫w�|�v��h��$bh�+(�7�M֜=��%�i�:�L���s�k�|�W�B@��3�y�����������o�U��u��)p�_��ki�ʆ)
SsS���;�&e�Q�&�K{q3QQ��X5>��s��U?�F�߼����^��2C��'O�|v͍�x|光�2f��H���;us��#k�c�KB�.!�ek^���
����nO���%>�����ƅŜ:֖G��E�-s��wH�[}���Z�\��r�)v�9�*�#O)Qڻ��L����s6z->��!v�?��5q
����ȅ����r�t���or�O��1Y��W�q�5�}��C�S��8g�J�׆S�%���Ȭ�������*�*	Qy�1%�}��:E'PU�^�k�j��Ρ,���0fS�s
�\f���W�Ջ����ır氲�t�5͸��y�����$��i���	ֺ�T��P�.�.��]�@��ur�k%`�X �'0�B�R��g^���'�������LϽ���=�I`�������*����O�b�������%j��]0�L��ͷ�F�*fj��r�S��ޫ���]in���h��7ns���Q�2�T�&�����21�_9;&���	��V��V�@d��9Ea�M���;�Cs_��w�n8�k �������u�b�$�� ǖ�F�Jz{�������Y2�w��	"��㺾n���b�&��w�\�v��#�߯k����7����S
׏l�0�c���_v���x<�es\q� �u�=F���.tD�Õ+�J�6�������n��}��>^j�EL^�9H^�m�)Ni��7=�o4��!E~oMyѷ�I� ��V�b|��w����Y�E�}N�-}j�;�;��^S�k�d��go}�����c���gS��K.�E����'��ٔj3���&/#���9�Vw�s�=�H ט�{�w��wc�d�|��a�j-��qas��R�>���Plq|�J�����͊Sӎ�Z�ؗ:��񹘥Ck"���=r����t�{�-��+>�����oDg!�#{�J��U�2��_�\<Cjt�oL"���2�,�׆{_G�W�F�fVm^{�{O�K*�^$���vƙ����>PbyYT�B(^n{�9�E��b�	c<�I��+>�y�qxÇt�>8�UO5�1��l+�
�m���� rB�ik^���#�$V��6M��rBϭqv�HsA�zt��N$�������Y	5�ƒ��R��c�{jcw�)�8e�A�OQ8��#J8��}�Ι
+%TV��nb��T���
a�2*\��Wӂ�����F|�=3݋�:��;? A=:;����wiS�I�u<.���9�j��7�F�ӛ�KU���
��U{�:�D2f��랝��\[�i˴��9�Y�]��f[�`#<���X쓱��m	��g:���%���7WԮ��+)�.�9���d
��}#�bzP�v����6�ܘ&��Yd˨���s���,�����,��y�2tٍ�J�C�1t�L��z�4��/8�u¬������ؠ�53PՋ�5t�l�'�5�u��.�̶�*�v�V2��vRYKU�v��o��&�v�YI������f좧2�z��ƴ�z�ᨻ���]V��2�B�=��n�=\f�|2�LO�k�zq��%b6S/�@n��C�Sإv�&3��a�-mM�Xԫ,� 1�����&����vxA{[�@���y*?��4b��{[���r�Q��x��\\1�*T���YVi"���t&Z�3����>"��$|�1v���7��J�Aę��o]Ud�����mͺ��sy��ɸr���J���:��%*�[�Os�M����4I��`,��=mQ�ܸ�$��B[�IG|n���@�1���i��ru��3�d��@�-FA�7Iz;r�Xe��y�s4�F�J!�3!��w�*�+��z�-��vd'��[�Y�ۜeMY����"��nHTR�<zfv�$����N尖���y���jR>'v��t��۬D��g�i�r����=>�9�=D�uEɺz�(���d���2;x��I[�R�nŷ�-�Y�Y�0�tO2^1q`uf� cLJ�o0;6���D�����I��Tz���!���\[+��[%�������.0�#�nl_�*ZvLg9�gΣ�@Vڴ��B�n>}�}�2��e�������G�F5��R �֫���>��@�}qdze�)g�}&��w�߿}����̩�xIM^z�ͽ���~����s�~�~�~��2}�w�*	��)B��:�ì����>�97D��y�x��6!۸�Uwzz�n�_�c���/%\��U�}.��z��[w�~��d���v;<�+wm�s��Þ�Ts���?Q����sr!�_��t,�0�'B��z��FIG�k��l��l�������>��*�bm�w���<=#�%?mʴs_n�%�����*z<�|��Ϲ2y���z����^z/%�/��_
{�Ng�5�	��>$��!�1G��l�����?��{<5fY�/sB��֫�Aw��l�6�)���m e/����b"gޏyG��q���3���\)�5������OHv��k�6�-�w'~�w`��C4W��� �_�ǬRB�epW/�F�&�e�����wu�X�:)0�q�f�!�l"!�G�9n���{=w��N,6}͆5<Y�i�Q����{W��G��������/R*cS�r�q����e���5^�_(T�E��C/T�|~��(�\��{�P���Pd*��0�;��T>��*��^�ײ�}�(�U&.���n�E^x�-{ϸq��H�"u�(��S�����;#�A�������:�߂u���	���7.��Ȭ�����P�!}q�p��yi�մ�������jDH�Z_�P/H��c��wN_���+�߹n�z4�*�R��Tn73c��I���|�����*gL��a;5�Ҙ�؝u�!OL-�	-Q��E$w�(��~�G�}U_5��~��YWE���|s�S#�(��V�o�t^�Y��wP��;��3��P�7���s��z}<ő��ż�P�6A��/��k�[���Gb�C���bֻ7���W8�<��^�9m�7�G c�Юs
D�F�_��OhՊ�tm�X�^~�Ii񖂽��0.��U*�|g���E�P�ѼH�;˃��z&�ͮ1qQX��|Z޹dZ��f�b��m@�"I^���R��,a�;���a�fm�E��sd0t�xø�n�����˭fa�2�|q�z��ֽH[q�Q�#s��BX�-��˕����x5����ܜ|~�5���t���ţ90-[�d����
����ͬT'Fìu��g�+��~M��Uxw�*�x2p,�c�`�M�qd`[�� ܙw��6�b�L�������[#���QcO\
�\n�S0�<'6������Mb�+�s-"b��9�Q$PC<֭�s��/$5-=yna�hP8_�r�����qB<|���RS4(�9��S/ưR��5��D��)RCΞI���M�{uپ�,�{�cy-��&��І�sE�y~?Y�-�/�d��~4!gҳF�{}$��1�Ž�.�d�����5����ޤi~+�C�y�U-&+?�y�ӾB�8P�s(���Tf�7�b����a������C��ON���×ua.�����{���7��G�O����DMtL){[&\؞U�Y��2�ᇪ�w��آM�XtĬ��$an������'+YPz���X�6u!C�KAa��F�̕~��7��1!N=#y|��ݍ�2�$@I�2����q���gm_p�Y�ɶ˵�R�� E�n�����'v��a>���;���r��6�h���z�C(�8.J�oJ���e)�\���Ɉ�Ͻ�����>���������P���{��e�zB�Lt��/���ȪKJ���lq���i9����\-�<��n�9��(2�A�sU1.�ʺ�B*b��?� y?y��W�w�|������4���M��� ���:	ʼ��A�m,�[77�w�h��
�^�_�9f�Y�hcŧ�*�����`����kdzP��ͭ�)ȗ0q.w���H񸙬<��o�I߼"��$(��S}1E�ވ��qe�/j|��OLe�+׵�K�}�z�@�5t|1�����x`��"��y���}�Cð�r����+CM�夵��9�kO���g��s�e�,�3����'<��g�:R�2��&kh�<�
�q.�U0��Y)�2;��7�t�٪p0*��,�zPU[Iq|;���6o3�@l�M�g1+JDn�i�i�+\׆�T؉A,�Y�hK�K��ߦ=1興vx3��;�;��fojTt��F�bCN�o&��3�)M�i�f���U�#�Cq��,��ǦjQ�I8n��z���ʚ�K|%֑^�N{�@E�z�C�w��k{4"(�	qa;�Ʉ9�ԫ��z׈�[��}��\Uك]nnpB���"Q{"isō��`Z�=��0�1��p��Y�����^"�ώ�(n��a�4�c����ݡ*CT4u;M6ڀ�={,�ևym�C#%�SG_�`C��ޞwB_�no��&��>�ƒF���r�"��O���^��G��U��o�i�)HB,�$T�
�თ���ST��^���}��$��t�!5�D�iG+�=Oy#�_U���u>Kp���f�F�1�k�uږF��3-�t)���؅ɻ��BC,�H��ҹ���qʈ��`�nj�`�ֳ\���cs|�}DdPf����@�������������O-?�H+�:���}��f���v��)�W�H�,ť��TF�c���n{]}�+6t��)�����8���EyQÒ݊����غ{�ue���k����t��}or_ԭVѴ1�fj���~w�3�@���b��N�
Ջ����c��ž����d����&m�2��Q@ڷ��w;�E%�~���_�Fe���OG����S�)Pi����{=��M�z1|���<��4.����.DGTr��r͜�T�ܗ��ʙGF�De}L+p
���5B��2�&�~��(���np���K:2�� ځ�$���� �jt��n�l��c�Ӯ#��q�T��H�(�E���=�ذ��3o���Qefk姵K8��ڎ�ˇIp���[�ޮ%�-���/P����q�*��u�H������yٲOW�R�&wUa�X�"��x��H���~�{s;�����GO��vӤ<��O�Ӥmc}<�K����0.�Vzk�7&�?=A,��:Xиث�~��J�{{Y�#đuo�"*Նy��	�H��ߋ���s�]z�]��.Z���m]lH�t!T_;��n��=O"����.��L���j�X0���_̂z��������C�%/�[��^{��.�Н�
��)U)�^�9̤��ft�]p3�M��Zó���zע�aP�$m�5�N�R%4׿\?u'R�&F����XL_�{#Ӧo1F}�q��B��{t#�����ԉ#�s$�j�u������t�f�b����6�HeKO�6��86컽#7�97J��J9L���J����؛�˦�il�N�B�N���s~�Q�P
�ι��[��cz圛��/Xh�->1sHeG�S�q�����ݍa�5-�+�������}S"$4����!�X�ܩW�ݻ偑�T��SB>!�SBE�ԃ�>�Θ��~�����T}��B�zX;���B6@�ly�O���wϷ7�a6kU$7�Ը�^,_�쯓
׏e���u�����G�#�+*�\y��+�?�O��"�B�u�B/g��ƨ׾^7�4�)�),<������DU�t.W
�����v��_q���H��DC����I��{�X���{w��ք�O�Hx��M���Xc#Qmcg�|�URz���I�t�
.R����|�ȗ1�-��s�n��`���-�ow(��ȸ�N�}8��W�2��>�n��L�����WH9ɏ����h���}�;u�ڕ�����.9��'��ne@�p�E0�6�9�OQd<�s���+�U�<���R�9)���sy��q�0�K�.��'O���O��sH�i�+��2�,����t͕x:�{XEH͘+��܃5�U�N�k�'u�' _g)�w;�뚳{�i�(h���.Q�]�3#]����\lE�|�&i�=y�刼*��7GR�d$�Q �ik�x��֮�w<X�S�>CL:j�p�$ǧ�L�i��#����I����\��H駯�~"�j�{�@E�z���}�k��ܫ����ťe��R:��c��*��9�}�3��-}w��_ �t�w]�N
����3��8��ET񁡶V�=xm9W~�����}���wi��ג��������Ɠkj`���Ol��p��LWTB��7�����J��������ӗl�'�I�W�-��u�R��3cn�;�Q<�7�%Ud P'rJ*� ��G蘈g��L���1i��Ϣ���6K֎�!�^�v�*�bsº��-��"�Ϙ���$�6t�l\����������B�{^�lm+>�R0���Zp������pe��O@���f��hR��wcl��;�"���-�F��z=�G�bsA��{���l8ہ WU)8�׮��9q��|�^��$k��a�6�r՛�D]���������o�h1f������7��w�Fzlҟj��\���^��
NN+s���e鞶0�÷�k���TFG-�ӑ1nr�.,04�
лIk.D�����X��Z$X�����ַV�k�u�i^f�C3O��3hI��O�#�V�R�뎟	���eUǾ�L	vEY6i]��bD��/]'�� �ȻA��*3��;2��K(�/w���n�c8���ܽ�r-��JFc<�N������P��vХP�ܙ�	ά�h��h��q
{�Ϫ�XV*�l=��n�5.�!����U]�Ǯ�[��2m^=��|���I���N'J˧��6�d;W�lz�ٜ�%۸�$�R�i4+UF�����j"�9��4�wP[��v�=�)%����ѱ��	��OI.����nɱ���%#��1�Zܾ@S�z��:����B�]��*�=���,��0\����`u�,�4kY4:�xLr�����!��gq*Ѧ��jv�\�c�6�A55�����t��_k�t9���Op�jVR�@�;B�4�4*F˺�5�hdl������l�tgf.	��2(����;��>�ι�sf(gY�w�-ఆP�wF�7����첗�Q_$b�����p[ۄ[.�j�yM��ok8q�	�k��]&n!ٷ�s���P��#%%.�J�����k��ڳ�/z�0=2�n�˶��j���Ŵ\�����5�H�?���=�"����r�y�l%�۹��T��ze�F=?`��l��S���$�����:����.At��a�t�X�!dmvd�Z�i����5��ӓ� ��dl	���(���\Q'%�[Eޒ^q��$o3��+9(m�g[��7b3�n��=�9��r���+�H�3΀3*wL�3T/�1���p(�5�[���ڸ=6��[�u6�X�;6i)�܇2���>���[3�y:dؙ�ݹ\��m7۳��`��w�Hr
�,�]p��f��u�#H���ԩ��&�ٺ�
��vs�!�"�J�.V���>Ș�c�{Q0�M͜Mu������I�~�(gȇ����'�Ϩ$��{���~E?�s'2/��/�o<�̟>�>���#�ϑ�?w�}�����ї�|���G�Y\�1�z_dbG�D~�u�<��(U���c�|}��9����\���dQ~n�Q_"!?V���}��G@�u��K�w��*�R���*�\^9��xG�_ ��>~M���㛺n�ﴻ��B/�^�%�^~wz������pL���__mum��L/����6׮�jO�_U}���e����gھ������|��|o�s��ܜV�W}c���O���7�FdW��~�y��_h��wD'!ί4���Q�c��?�E��o��gK���6S����Ԝ�S��#+Vc�a�����Gc[���'������� �A���4�Q�k:s�){֦�ڕx�]��OGv��Z�!ly�G����Y�i\�J�Z|y��#t��o=����^�B<7�8��}�9�����ƋXw���znU<|��e�U���t�����Jw*�*�r�
��f��D\`kv��<;�Gz�%�<{�T|����gHB�q�#GB������]7�O�*���{
v�j�I�ި#����{�Q�J�]$|}��Ӽ�SXI�|�<t���b%��������6�<Q�H󷔑�9<ǋ�@�T��=~���ݰ&->7�M�D6EP+��Xw���o�V���^�(��(C�a�x�j���<UuN:I���H��ź�LUar���2ۻ�*m��`���7+],�{#d�:.b�K5�:��ή���\̦Np���g�&P�Ea�!ŽWr(B�jr##���w�x�>/�?���T�;Q��[��f��{Q�܆��q"�(��3�{<�Z�4l�m��kϷ�0C�����X��:���ݛ����� �jZ��-!;��㳰x=:g��Q��:\8%ս����6�������C��l�C�0��K7�mB�K\܄��INu�2%�]����7��F��鋘��q����}�T�����Vt��a�[�Ѕ<�1h�ea�M��ɬ�`�P^����u3�!�19�*0��2��+��6���UvMq(iS��u�ۗ��2d�q���w�mF�yW��K.W�Ԫv*1�**܀K7�K�Qآ��l���k�vg_{��Έd2kXR><�A���Q�5}Cˈ�t����^pVi�*�:A@6>���z��l#!�J��/���10�0k*�i)Hv¹\��ީ���++]�
jԝ�ZY�������&;��PJ?���;}Z`ON��*����h�f%���*:��x�̻�%��f�r`���a�xt�_q�����gk̑�fK���ϑT	��Tj��1#�q���h��1���"��;I8��U^i(V��Zp�L�*==/����W\)���/��H�V�.Q��@�D����Q�}4^�R����>i�e$�[ձ�7	S���y��1�F}���h˱&��t��A������s�g�E^Q-$� �vƙ夏��ud8ۼ\YK<:�7՝�B��٘uwI��Ό$�����*R��1��=����ҨZ�:����Du�D!��CN�%R��|.�{z�<T��z=�G��Νў��*�s�5&l��ӵ�4��lЎE(j�Ej�/j���m�V�-6��J��ߣ�9ޮ���w�L���JۜH���L���D�qfY��w��M9?�˫����_������K�ȑؑÏ���EZ�7����_���Ey�S� }�]��EF���1��WDR�}Nc�1��ɋ�ʛ����/U�i�Ǝ`"�ar�(t_�Zy$�&~I����Q��B��Ⱦ�קb�rI}g~#M��;u��woyqj6}�-�~0y3��Ll��h�:����յY��ǈf��m�|�x�CI#H�I
���Ѻ���w��*B�9�b)HZ)���.T�Oʜs��W0g�^�}�f(9U��w������#}�"��`�8R^��0ʕ[�N+ӎ��@�܇9��T%��c�#®N�c�4/B�'>�D�c��j�t�Ǯ�Β�5a{�I�]+5�u+c��}��
R�U�E���K�u�xws�J��f������Ӎ��I��v�>��X�蘭��f��戾n�����^����R��Ͻ:C��_�U)��p&���dV�8|z(E�<a�!�qz���/��Z��C�{%T�%�y�������� �
�u4Q��������֠���yON?�z�a�W��)����[��vb@���P���&�}�ǩq�~b��g}�t�3j��w��-"���� ����$.|�Y���8�n��r_���)�W�jȚ8а/Z;C�v�4��L�]�Uޯn�d6}� �nx�_kڂ�V ��s4<��܋^~J�{��^�b�![N$%$t��s���3��Ip̬�/2wox����)�Yç9F�C]T�I���p��On��n5�À&܍>v$�b��&��#��Q��G�;`�R
�qaC5��]\���z�ޘ�ef��AYƍ�-��F�[>Jom͚�H�G)e���p�������ӶˌL=*��sBd�������g�]��?����Sp�f��Sکr���7&��k	y�����?T}=~�Th�B�8��DQ$fgʌhJPr�<���ܽ������}�2�:��S2$�bӦ�2��\C6��ڏҳo;��xkd8�<���/���tc����⋥J��\��g6�zvD��j�u#5]�����Wd	���=����>"�?�:t��ƍ��6}���mv��9�G.6TL?]c��CHw�*���ӄ��ݑ��g��P��Vs�O��,g�$�"��`�%�凮���ߪ���Ͼ���^\]s�����Hז���@��6삫���S!_Y����5�=ku�B��-��:X����y{M�U=��r�VG��ё#]�n3��ӊt�8b�t^�Yi)�z2l�5i��/�bq�P\��̀r�4�%�ImƌRz=BEC������f�g7��U��Z��i?Ĵ�9�oC����zF�����tsHY�A��קҟ����5C�}��m>�̺�>y�ڜ2���*��I�o,��ؼ���~C����x�{�
�h���q.uӘٹ��.��]wwq�q�ڼ7�3���5n]�T��[l����X�Z,�e�ߣ��������3�}�l���c[~3���#�RәM�d�@�>��v�o�a����UhW"l�F8I�x�!i#���n�+��D<��k�Jό�p��|����1o-��s��i�զxJ1�H��GW���HJ\r}N�yhf�EU��3��FK���k������{�f2�ϱVLN�ͬ����P���H�6��sz�A�؂f�T'b�U�A�8I�V&�����u�����e�Vݧ�{E��PV8L�=TrҠh+���{��c�3���}&�J+���"�/��|`�,8��%����O���Y�������m4�/���b���=a�,���F���p���{y��}j�:sJ�^,��ُ��hY]VUz����_s<�JK�v�n\,���������*й�L�,�!��Q֜��
6I'O��D��͜1����EP������5LD�^w��T^�J�3�x����y�����z׏�o�ܻ�y�����Y�V]�X���L"�	��6����50ֹ��x"�9�W^N���|�(
<]��6�cu�%a�M���i	{�x'u~�iӃ��x����Ǔ>��jcd�֎f��=���̈́D>�y
�|�ܸ�li$in�2�jy]�hByK����s�<�:�h�M�J:j�wn��.�"�N�B;�*�.�p9�5�}pe�4�vu��c��%Z�U/.;��D!��_���&c�1ȟ���R:����4?��R��x�H�1���2%ʞ:�8�<�b�NU�{u�`[�B�t�!hyH����O�^R��vo����A}<���j�Z'���z�N��3�yg���j��>j�me���v��H�z��|��,:F�l�;���[B��}�1�R.8^.=JG�z�c*��F��&JSO�qn��WohJ�o#�ճ\��;jsO�����������Y.�x|�~yO~�/�੐gA���u&j�D�ʙ����-D����h[����!�R�}ٝ�*�b�ZE�c�Cǈ�#Kn�_K�/%F'�_�����UL8=f\��W���X)��ةWF���S|^呹��R�3�q�K�q]�R�An���biD��;1��SQ��u[�(v�(U�ӷ�ι��y�ҫ�[��3,��I����m���$����Rk28�W<�*{�=��j�,�Z>lQ�ԅ�+ş
��}�͂5.d0|�.z�����ˡ7��HT��p�\_C8<��32�mOU9x)�Yç9"*�1��!"�n�.��~�}��axGw'>*zOU�j٫�z���D��s�y
�0̄���*��>�_ɹ4ח�Ma//T�y�����ଳ��id;D�[=N|Д���my����kt_��x����L�fU;�A[�����!�(/�y�������/�qB=�*�ǔ妏������og�MV��~ۯwQpHNV\L���!���Fj��.�m��:���eB��)TB"+���_z�8w7�8F��~8����G׾X����Y(h>��H�r����ZNu�EUm�l��`1!M�����m���b Dے�H|��G��÷Z�3�\wd8*p��̬S���̝}�/u�,�l�O�!�t���Ni��T� $ؽ��r�sd��0=ɴ �z�r�����;h�`4�'A�T�=J�A����q�Z^R�0r��=�u�+�<���4*GeȦ�·t�IGkvn�Q������@,�a�=��y:��]GL���6�m��G���Op�Q�9M�z`wOa����7���9s;^ॲ9�;�f=��N�ۦM��yb
u��ɲP�Q ̇��0t;}������4���8�+	8Af�2��[	��6����G<�d��Y�b���n�/j�e��Ut��k��Z�9 '��2n%u/+F�9׸2e��!O6�h�H�fY!����T���Wm���F��n�^oNꤧlwG���>��K�=,�3�
}�NR�j�Kvj�%t#V�=�q�u�+w ��n�U5t��g��ff
�Uݫ�C@�|�0G��⹳��g#�YR�����S.YcZ̚h�#r�}�3WM�j+��jܵ�'ѻ@�
V��ۛ)���6�j��v˽����3�r��\����׶�s'f`Oe\�y��mvKT��l�3;��ɷ&�6κ�o�#w����3V���n�֭��V$���]���Va���TO>�p�դ'��Y�ۺ��F�l�D��!��Fw�y���� q	:yQn�2����(w�/���챬�|��r�V�uՔl�1�M�b���Y�1�H�78�c*:�(�jl��1f�7$��aon4�i'�1�����4�b��9�f�1_u����L�&��.2���r8/��d8��M�y���~��"���3xY�u��NvX�ʡ_4��uwb�.�$�D_"k�(��5̈���O��|��>~�[}�~��_i߻�ʿ�N�V����;��d0��Bjc�:�m	l)9d�d꟱3�v.���w|$�#�ޞ͗Ϲ��9o0�;4��
����g��t�K+$̲Ӭ�7�7���~�h�c��ʤ�i9�4�:����pC�㭹�3o56�þ���>s|�ZY�}��$ �E]Ц��u�v�_t�{���wb�slb|wv���n��	�H��gu��a���g�9;��"D��pe�Cw�u�gɋ����5�7�Ѽ�T�[�j`]z�/�b�b`�d��*��ؤ��1Kr?T⒟�~�%�?�S� ����	Dw�Q�n;;�C�]]�u����!�*՜��vX�H�0��i&��\�1����WA��3p�b�.Dj�c|��n���N:2�UC����;�"��5��v����0�u���&���p<̧Gާ��Ш��/�􄑄Tמ��*R��u�5Т�7�,7�뙤�G�ĩ �ah,;d��o�Q�l]/>���g��H��4����L���ۮkb?%�
^.��e&%���W��_o�٣�Ŗp����!�5�#�ͱ�+�i������{��5{�X~�[x���C�6�?Yia�Gq	W�I_z�T�k��p>�9����T���^RE�0]4rs$C�zW���'E��jأ�W��{�^˫������t�Nञ�~�_��/_w�����l+�-�ch��
ގ3�
jK�yyӴ��*Dr	|��������y�#:��J�K�!���M���P~�ۮL���լ�c�\Ī��N)Q�祌\C�~�AO!��^v�z��y�Ք�^1��HJ\rS��C�Yw�C�)���H�AJ���)�~��+�{����Q� �]t�a:�/���^�[0�s�k�K����D�'��4�*����;=3>�[�9[�b���<�-�TY7���&���o�x[��ZaúV^,Z����:�6B�!G�#^�o��!�m�ޞh[[��.-;����%�.�z�4P\���H�$�*	Ԏ|��s�h#Hz��]\�)J�&;��Lл�24�XZP�xC��.cϴm�//7� 9�Y�u��C����E�^�ۣE����z�̬��X̐�X���]�\u��Ô�XS�ض�ՍZ����J�I6�m(����$���KzS#�}�F��vdƖ64^"P"�d1���ƶI��=���7yY^	����J���q�Zv!{�~I/��+&ٗ����w��08�*<G��g֧!��ʄ��`���n�u�I@�,�ZC�������i�H�Ν�R�M�}{����q��=�����oZ)�`�zp�
{=]9��g����g����{�!=�Cj�H�?u�_c�~��q�Q��k<���FN\9ͮ��/��ڙ)>Ը�	Ae�,��V�yw��%���7D���DH�-��_�����E�;�TE�<Q�BZ��	s����� ��9�tkI�
�9�ü��6z�1���TFG���OK	������<౺�˝b��
{�G5ѝ$j������V��mۗ �^,MޏE��yT�XgW�`̭}�&��ʻ�ā��a��}B�����[��d�]�%a�B�h����1��Bʪ�u���=E��#q'�e��̕'1xr�)|��/L"�1��'�>��v�ʘ���@�� L3Bo��:3 �3 �<��x�4�O�w��j�*���MO1La�<i�o]G��vn\<�
Yҹ��/�f��q�@��y/6E�=:"�uj�m��&�*��&*���{�l�H�1��d�J�X_�^V}ࠗ�2�õ�'b^�+�wg�����Z�vִ(r^l�:V~�k=���G��H���x�u�~�f��׈�f�f���ڊ~��ǆ����Cd%��PkO�}A�4���5����ɴ�U89�=6"����K"�#-���gP��馡pqn�:�Vl��'�iM\pӝ�®Wu9�@�,��d��Cڴ��J6�dd@	��tE�F�B�5*jN�g�Rw/�f��6J԰�!R8뻡j��S��y��di'�/��"-
��z��x�7���Z�E}�1x�~S���t|_�ZBO2�%��$:�ڹF�,8v���[�(M���e���u�N�=%�O��I�P3��q�gs�;o��ݩW�y܄G���"e�㠋NGP4�����3�4#`L��4�o$O3f:��뎙�z��|��졗��,$0���^ueom%S����w~"0��T��C����=���oT�����{�NLܽ�)HoG|Ti�)KL���@7Xh^�w���ˋ��4��z��*�f`L	�=n��*���_�����8z��o��1�X��ť�����ԼD$�q�������Wd5*{O{��
�[�vEX��x�}=hnV�`E��^�@=|zs�sbE��"�U�����ދ��r#�ŗ1�Z+�p1Ϣ��R�;��h�#���`�����X�ܖ����wOE��:kT5BvrD�߁��ZEFbXU5��cL���t�A���U��V?�,"�l=\x��Ɨ��X?YIa�G�����W�M�3(Ɏ���{),������[�<sY�m�m�H����rd�Z���)\�:����ĺv]�X���HƓY�Y��%P#�]8`�Gg���]H���.u��qc�o�r�u�:�g��������n@��I@c���q#��nDW��Ygw�}we���HW�sHq�6��Ӽ�����C��-�f+���~ȸ�?u;���K#�����쟗%3�3>�[.9���xǣzG�r$����^ں��[8�3�v�+A=�R��K�F��^r�R�Ba�E��~�����ˡҝe��IV�q��$R�N'>Nm��y}��Ȧd�6��)[/���~...,;�Y���Cf?#�Y�<�1<l��@-��K�uP�b��[p/,��sz2�����LoT;�vs�n�N��{�OC＆�lĉ�ig#�jJD�Z�-S�ͥ)v����I�7.�^�i�3�ia-/���tȁ��@��c�!�6�u}��Ţ1��9x<��C����0���#!>��Ϲ�n�rwH����;���ޙ���y/y�^�r��Y��"7W�Ӳ���RӜ�4,r�⏈�,�����ߓ}7٢�����X����f�g��<`�wu/ܬ)�K�eG7m�7ި�B�%�=���)q�<g$V�[��n'ts�S���ĉ�\����`����@Е?N!���yH�U���3���m��)ǪR���_M���Ι
�i9B�����bÃdi����� ���������*�<����L�CB���V�aJ9o*�ᵎ�q�p�#=��0�Yb�畏ry#�X�c��5��Z'����֫����l������ٲ����P����ָ�nZ��Z��s��p�ܾ*3=,S��kK� �b�=)�/�-8��ǭK�r��tu�We5�z)(�B��Ǔ	�����������}�}��+�y��ў�,�,��V���k�K C��zeNt�f������Q���%����e�"���Rqk%����:t�%c%�w�s�\t��:zm
���4�e�ˈg���b�<;ò�ו�wJI��{��r]c`����	��	��`�=j�[�o�}�
;��<�N�E��{sME���)$F��uL��_�=.R���\�EB���BR�iw����Q*>�luҼ^��Ī���zn�%HQ����!8�	�S**��wx��6�I�Y�odA�f���J�m�؛�rA��֤�Dќ�ȷsS��Q�N�׉$�^;����	��i"&�nwd���T�����&~d�ҵ+k��$��~<`�mW!�=��ɤJ����P���8wˏ���}	c��T�sg�:�w��c9	�g�|��L$�Y���a�ZY�17�h�Ф*z��ٷ��I�Lxr�R��,o�N�<~�ii㚸لC�m���o����'��-q� �k���������R^mJv��?ow	�����L-cִ�Yf�7-��s·�d�(���0b�?E%�(z���,�G/�U.�#��Ż�GP�T*�l�k@NsrSWvQ���"m����,1yE�8��N-�?RQ�]�6�ت}nN;g
��b��pf|��n�-@S�&3�A]��Sd��ѶY񷊓w\vvT(GC��<� Yd鋊�b2�}ú����S��[��4y�G�W��"�ʬ�"v��j�##�/L�嬯^�����u×��4�UC
٨U�fz�[�ָbD���qJԝ��YH�ל��Z\����ek�B�v ����V�x_a�H�0W0%g��!䆑9o���������^�I���
�����\XAi�?=>��D�b�m]�u0Do�޴Gެ�jŢ�1Wt��a�����C�kz�2Ω��"�}�ZpU��&oԅ]�AA�憰ԙ����EJҀ3�Ȁ��Ek{$�C�/=�Sk���I����w'����r��+��|�}<撰M�=��P��{OBmָYn��yB�Ī-�u�u��q�^CG�l�݁i�G�vP�E�q��(���B�d?�U�a�g�����w7��M�v�v/���+)Ӕ���x��Z���њ�r�o���
{�9�'
�qh:�fv��Y��ȱA�+����w�M��.{�-ո�I�Mԥ�$*T�y�;����%�d���b�,���k=�õԜ�.�ʔ;��iѹG�2�3�6��VI�TÇ�Ǔ�]��dP�E��vB6S;O-��z��4����75�HV�Qv��Ke�J�����0�vS������M��{���j�9��"t5G�+i��vb�wΦ�s#"�K�7V��\"������z��#,���mS�uϴ�:�{��ޝ+y\�5��uSΡח�r�1��T��"V�M۪��F�]
�YF���ͦ7�ۀ�	˨�eaܖ��\ZL�\6�\{~�S���ro1��Ùnk��f@�#�������Yp���ێ�����oS==쇵	��f�qa��ӱ4_۔��ɫ3N�|A������J\��qA;n5��h�ˣS�ntڸi7U�Z�wlwZ)��f�c:)-�m=:�!�uŉ��w4Pg���Vi0���K5��5���x{)X�<%G�J�y�'Ҭ���@�.#;�`@��˂��b�&,��܆�Ц��o*��D�b��`�E�k�6��XK��1���~��Y��__u���n�+��G�����LZM�֜�]:`��W5Bڜ��o}c��VҚ����V�!ٯ1d�{�x�������o���=�(���8�&�W�l�"��:Gٖ�w���S�o5�����|mV�g$�19	KL�z�u���X��)�hV��u��vpl�y�Jh��/'Az\�!��''7$1ҿ�g�EEtO�UgVwn�ݤ�s���L��1>�[[�G���~���J�W�+7�<�}o��$���4������_��߿~�m��d%��[xL�D��K�Y8�T~�)��*�mx���}}{}vb��dMH��Fe>)Gg����rƚ��Aԏ���[89ی�#@��]^��u#0����&��љ��6d*�|�D���D�c2�iQG�*P���ˮ��W����h�~IQxa���2�j�R�����v37c��ݱ�㍊e��<uz|*�D�bhg�.#[��W�n��ɬ�`
V.�^��G�b7�L^#&^Vu㶝'v4�CS
�w(u[ �hN=NG�����o�p�Ӣ1����휎�gz_�8�@)�,�4'p�[�Zn�G�yv�47ry��E��Rwr3%������diz�b�](j��R�?`sC��w��%��Wi6�g���Eec964�D��S�f�"YY�a���5+����j5��*V�y�42T�W�(��z�2�OnU���y,�k�s1�����5-���9q\��x�z���im!�c*��7j��\��ۯw��z]3��Wmǰ����iN�UA�.귉J��<[�fܦ�OsJNԲqH�۸��T���r�	�j����Us{�*#5$8��[+3]��v��Z�66�y�zIJ���t:<��eh֥�F�Ԋܜ׵���)Ũ7�{r�v-�]pZȒK؞g�?Lf}}C�g}��Qw�ئTLp�q� d��أ_�����,��v�;�iI��7�j���*t��f�����nQ���T}��̽�)�B�1ߛ0�6��� (�2�x��㓶�^ݭg!�g#%�Q��_-�R0>��M�[;:���t�8����5s�=�y�"�/X��yp#��W��ȪY%���14Cs���}�	VYGX�Gs�>OGo��g1x^�V�9�Bq[l�5T��v����	YI�}��y�6j>�rOcc//E2/z�8�u���1�d��s)r?]�ki���aG�K���5
���q�5(c�����,�C5��E,Y}b9� ���tκ�C�N+�t�'�u��Fо2tD���KX�eF뗷���%��QіM��4)H�y�t�ɯ&�VQ��=7�t��H���$��IV8���{�>>�+��GLV�}2fr�`@m�[�i�P��$M���6ɌULVuh}�O�ya��S��B�%���Io�������N�8+�u?8�q쫁e������jt滳p0�b�gRj
{��]�y��:8��~SZ���֘.ќ
�[�4g6�E�}nL�uyY%%F}�$Z�kn������(�1��׌ެ��6ZB�v��ێp�1�3:�PA�P�}��	����kK�>�'�/�5�]�i1�����X�:;qD�����
&_d7gOEи:��)�f�AX�׹	E=�\�j���Ɋj�ʨ����]ɷ�+8�p�`\PW����%	r0��N7j�_=��!��+��D�]���Z1s�8�+,U�7	�����vB�Z���~�֮"cjxF����3��՚2N�Z7^�\�n�F�P2&9[�=�\�io[Β|�,�
&8�m�?]D�Ǯ	��'�WZ���,�|��*�%g(�3qI��,��Q^^~�X�ڔ��k,���> �4�W2�(��!�V��'�S��3�ŷ��k*�OML�D���J
���&��3�3L�<w"⦞dҌ����9��@d�'�]�3��с7v�����^�ml�	%����S�ł[qz.A��yªͫ=0��g�Ź�pr���y�M�BVȺ�@Wl��-������|��"/_m�w^�o��x�*�\nu���`�V7N��!�<����x�B�����o29��yg�L���J&�cC��-�p)Gg��g0�($hP�B�3u���yQ�����0:��״	��/14��3���V��
JbZĚی������_����-D(�a[�(�V�Ѵ�nJ 2�`���Q�X'D���Kq�]��2�+j��t�w�öOY���w�]gA��v�7�S�����ع���L�����7*�M���ή�8
���}~fgθ,.�[���y0	���佛�WC9��9�&Ywx��3�^���q�s&�}��~A�-�3I��l�Ƨ��ݓ+���a��E��հ����3�8��U����M�Z�;6����}ǅ�ch�ލ�㫯�f�A�w�1-{Y���Nv�N�N�M1�oV�Fu�b1t��w�����u}���eIXQ99~�����əӎ+H��َ�Y�k�r���D��[�S�<��|��Q��f��kq}u��Y��/����v�ݰv����{Rb����O�F5�r�.�tPZ��$C
���G�����H�I"�H�0�'��3>�3)4��v��T+�ٗ=��+��vꗳ�T����C_+�l�s�OP$�%:��PӧX�Wf��5^�y����7'EV�/2U���SGݲ-T�-s�f��\��X������|��+�%���⡱r-�Xp	��O۬y���PL>��j�b�T�q-�7q(fD���GEǭ�j3w���G�Jvd�Nf���o;�d��ݳ�.Iݺ�K5ޖ�*����G�C7�*�ru��(�'���.��p�����gh�C�zy9f��'�y�ٻ��4�IL���l%�Ĵ���=D펻7sliN�w���L�t���8 ňv��,��p(��pѫc;LNj��e9����P�rw��#V�GH]�9o���b��x_���%�`z+��|�0�u�w7�<{��𮞡�����W �䙂�����M�e?�8�.��υ���nb�lq�qyC�7̹[����X݉O������6b��-I9Np���;�Jf%lފ����}ǛTmƱ~N�9S��\�@{Ց9)�������� T��V{DTg>�5�AM\n�j�wz�^��<q'���1~��k|C1WdN�2Q�b�3�q���CA̗�bȖ�5��/17Y����t�ej�$y�β��w�*��`�ߢ�#Y�}�hzb���j����-%�:�a���î�s�q�CKW�Cw�[�&)nE���Iw�����~�	��gQx;�b6h.ß1�S�u�4�韴ɸ��On��19 h��>ۈ�1�ϓ-}lWl��&x�w�οh�b��sLV�ӄɝs0�w�����q�h�aZ�D���w�ə����2�d���]���!c��R���s�X�����p�[�����;w��ᙡs��!$�ypL��pD(X�vN}'�v���-y0��Q3|�3�-��]��9��9����oڻ�e �=T���b׻���*�l���Z�7M�x+iR>vWd�;��C7�A����������6xQz��IL����n�W9CM��I�NkQ�#9� �.i�3NIMƌR=9����Yois������cO-�b��:���_'gL�r8�g�w�k�0WQ:y�^ۇW�s���09���;����*
��2��9��;!ȒF_Xs��;}�}�,���� [��\hdL��Ҍ�+D(�����t/3�+�u��cEto*�����z��u��KKi��t$5bb�Z,w,�\��}��
b��f��&����:��.��ڱ8�������(�|��=q����ږC���:�I�9��y�P�����Ӱck!DGќd��.��i���ī��^h����N�N�,�#f�1���\�bRh	%�wkY1ѽ���ؿ���)̗s���{��nBj��8dYN��2��l�z+;y�n��7[u�ƒ�t�rrT�&���H�P�<X���X����n^�8� �䰍R��r�)����v	7&a�B���t�Vi*�]�j�-$��Ĳ�S�q�v���)�{&���=����r=�j �v;T�n��R �_T�z^\F��{s8d� )�f֒��Iıٳ3�.]6��tJ�}3m��GPT�`�ʯ4���6�t���ʍ�; �X�D�yϓ�����y����p��lѕ���F�i�;�2��w����]��B�h�zx����c�^��n�1򭱧v�ݾ��U���N�bMrpoy`�WtZ��/��� m')A����_\Ud9���,L�@�dͳ�鍼��}VSQQ������u�g�	�Ӈ*��ʂs�,[<�����ul��|F�d	���1p�s�S;��z�.1wW+0�Tp��Y��'k/�(�^gd��N_w:�WDdR��Ri:W N���f�V�ۧR��������f��j���ʈ�j��d���ӫ6\6��fH]K�u�B��V���r�n�u��_aމ�uhF^qޢ����%j}�6��u3����4	)Ѽ�.Ұ���gR�/�ʛ�wJ����a{}-��
b��Ix�;�z+��x��΢l�m���F��Ζ4ݨ�]���}Bn;���*���Ēq�Q��guw����p�6n�N���4�ɼ��L���5����Y/W��M̶�����R÷*��9�՞���Ld�e_J��+����{��"�cn�����S����,��k>a�+9s�Ï�Nt��V��D̬]x_�3Oog+���=sD(�I��������^W�"��3#�ϩKɴg�U�g������R����ϥ�=(̢�/&}g;���'&T����K7���RXԪ���o�*���c03xU=#;F�$Z�&"b�|�lB'D`�zUQ$iNv�������E����ӒUB��e�9TK����Z|�'k=�3���zEi���>I_D3��]���$G2�{l�j��U*Uᑯ;2�Ki�w�U;#�f��h|�6�t)n��T�7�5BhoJ�������a��:�z\�3<��\��W�D6�Z��P���)�ޑ����<+�޳l\%p�k=����֘Wn���y/	D�K�=�3[�f_���s�I����]��5���%aG�';2��8��cqH��Z�v�`�A�s�X�.䯺�-F;b
���t�Wl��U�v%�v��e��%�xec��4_#��^����i�
1������+��z��ك�}��?Mto7u9��^RM�>>ĘsF�l�UITʢ�F`,����w���[f7x�6�[}xz�{9�=[���,�No�)�!)FeYň�B3vL�%���Յ��n�P�ugM�{�.�I1��\M�t/f�|�S���n��'ne��w�*MU��(
Xz� #�R7t���v]�Q������쟳#f���n礩=���vn�
��ο��9���
����]�)''&���Ad]W7c'�l!�U����Zwlx����6�neC��vحn��0Oս�l�#5��ga���j�I)�32x[%�Ƨ��移���t-O_\s)fѸ0�h���l��d��sW�ݛX�آ��ԭ�5���ɘ�L��k�Xm��ү2�k6�δ�4RC���d87�'c��ۉN��n!�m�ʱ*�y�6�m�7���;�Jq���me�<�C�ʪ׌Xz$ڶ{�"6�S���2[�u�!S�vO'�n;)ѓS���C��*�\���ӱ�������MK�{7S���.��H���]����j��������}��SW�뾥:�n�C�2b�Y4�r��[���
�##��A�\\��ञJ�����^��C�䴙�Z�Z���+�5�B+�bȖ�`6��YA=�x"�i:�h���D�n�e�ȼq8�;�J��Ht.vbEN�;#�X.�n��<����K��rÙI�yk�&��*g+P�����e�5~b��PH�{Q��rY5m]��a��Ԙ~�T�&v�]sE�*�R�����]=;7s�{�ƽ�b�W/,�4)z���{iU��[à�������W+,��cՖ�\�p��r�r�[!kj��n�"��4�>N��Wx�kq-EIN�$�p��Q��/�1��8K�]I�|�&Q�h���c5�����]��z
�\�ɀ*fGc}�7q�829TD�ĺ٭��e'F��|U#:������Ha��C� fsk����8)6��+8z���D���]��E���z¯P�- [��'��;���\J���UzP�/
�2p G\x&�7�Z�y���>5ne_{ϱL���H�Al��� �9Čz����Sƴ�s�TL%�zA`�^��8�����NT~��t��Z/%�7��+wܯ�Z"#��������D5{o/� ��d2�hMaV-�&2�����-�Z;-n�<��)q�����I=�ҭԧg����IZ��X��gG|��L�ݙs�l�!�o�J1����
�%ު�\i.�������ċQӷ*alX��6$l��%�]Y[���ü��%N�g)�5�9��Mb�0|S��b��,T3#��yj�M�ݥj�ڪN%�Qݡ�P��GWu�ᇗA��6l̂�a�h\j0̘��l�㷨�N8���]���ӾzBK:�_��=�^��Fs��vώ�'�o�vSŰ��F�zE�`�盏XEz�<��Ss>�S��/r�(���ڬ�pGm�r�'a�������_�1-�>���<�q������&����$�?��82n��9z]����lM� �2�ơ�Y�5Q�e�""C���%K)\
�
��ۤ���K,<�#M���P!	�e�顚Hi܇�Nq�$�O_p%eeGt�1�np ����JOv�b/��tޜ��q��w��.9+�������ot�[� �-��o;�%�}/�F�����/26h�Yl�#�-͹���t�h�a_��{ܝ�ъjg6����^�,`Kۀ�9}�Bև�����XxJ��ag��HGRa4�v�2��b���X3Wja��m�MTCJ� T�s�G�̌3� �2諬�FCkd�_���f��ݡU���U�e�;%+p�TAZÆ>]�K��]�Vi�s8,$���$q���]�!�e���$��֖el�`��>�%Ɠ];{	�-�_�3��gKQ������ᱨ����hX��B������r������Z�˲�0�6�K������2����[0���ڃ������Wu��*�^�\�K]|r̎N��m�Mͳ}�ә��ƾuy�2�v%.�K���ܺT�U�3]ի�5&>r�I�eBˍ(ӭ��8���쇘Va��)�m�K0��l�G^���|Ҝ�7�&v�����r$7Ci������X����uw��kb��o�I���@������ڟ�j�s�������;��^��ތz��>�kz���Խ��s.�E̴����Ț��ٜ��4��I�Gf���V�ݸ�ʄo�DZ5�OA��N	�QjV, F���b��eû�-����v�VK�\�����E���	>iv��d������aSq<M��μ<K��h�����Ӆ[YUW��
8�U���.�g��<<kno�U�������1>�}�V�}c��3p)�UA_'�hz�u^���*m�^y�����8���;���#t�V��zUU�6�������5NM�=�t���N�w_�6%��y���_���/��uN��Mpk�o3w-�]d# WIEߔj�Ư����{"�}H�z���A.�4'�vºI���إ�k�,c�gksuI���(W1��������hINn��w�/+"MB7��)��bp�J�p�"�� T����pJ�F�d`����9���G������W(��e�纙�**��r�^i�[!qD�W]u���D�TT�U)P^+~��o�cx�8e3���>��1b���}
�Ǘ#di�H��BMN�I`���5Ȣ���VϪ$�%��M���}�UB���$lJuvb�>6 ��ì�[Ux�lH�x�uL�W!��M�Lk�[GH&rk�Tc���j�0A���?��]_�m9�x:�X�R����-wlt�v�[.��;�ʂ��B��ȐФ��h����n�6S�5�%G�_C[�TWx�P�!����J,:��*�B�x���eJ)� ���JN-��B�>�vm�����<0��fN�X��ACv%��˸z����է�N/z�Fٛ�,c��<*N��!(En��t^QCj��bӻ�F�y���M����g��zɾ��`s�,�������`�j���=%�Mhm��a*"�_1ѭ�!ޅ�*_C\Lo9sMo}]�-<�i�u����T��R��s6`*}�+�НC]���W�����=�[a�F���wʠ./�ؿ<��}g�~'�|�#��q����AR��H��B"�KQG�DC���P�(��x���HG!���6,h�X�.%ɚ���m�mC���<!brb�	EQ@�` �E�*��*QH��PUU�QG��x��!�[8?��?Q"�
(���(���
(����PQ<�
/�DDEQES�(���)�!@T��ϣ!x��{��>
�@c�h:��Z$�j�hr��i)?�E�+ �*¥H$��5���{�=��κ�(*�.\B��b�+����I��`��t63�͆�D6�,[��UD��O*HV�D������x���`k��(��Hy�������`T��Z`!TC�] ��C� �!H�~�>����>������D>O�,����\8�,?��������60��e?ܠ"�l>�jI���q�z>Y$����WE4}��`�m�4O�s��#r�>������\�xFZ��4�?��|�����,����Y?�2�i'�~v��B��8{�S�&<,Qc����B�TDD.�	�^�Ix@�%V@�U�^�FF(V��E�U��?��n'����.z/�
 "�P�$�䂔AJ��R�H`B����?=� ��O@k��`z��mv���)��'�ܦ:��O�W������р�� )����գ���z>c�Qr��d>#_�c'�����Ō�
?��=ï}�z����O���~?��CO��c'r?����>�~��ǹ�r~��~����`��!������Xs��c�0 ~���� p�`6!������Р�P�{�Q��� "������B'Fh�1O�)���Kp��?�X>���>�i �c �� �"��-$H��X(�а?����e��������|�b����r>���������6+s>���5v��H��D�|t�.\�l	8��2"�@��{C�,��:�G?H��!X��������;�~��_�ɰ>������|���|O�>"�1�����a��h\D���_b��a�K�>'`P?I`�������������`�\��>�p%��ȡC�~O�~�|P>�#Da)
�������ď� "�R?�@���8��a�P�p8��p~?��}{? [�?7�k�5�7�4!$��}����'��?K�A ��h�~����b�������������'�ޘ��I�}��Ȁ�!c�؏Ҏ2�Ic��=�
��G�4����O����cҟA�}}T6 X���d��p���b?��4�?c��'�#P��?�c��~��P�O��$!����}O�׽���P�3��� �p��[��l9�
 ��C;��a?B���=�#�}i0�������:�rE8P�{�Q