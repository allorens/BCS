BZh91AY&SY�s [�c_�`q����� ����bH{C�         7�R)B�UD�R����IR�BU%D���HR*"�"R�T*� �HI"�H�$��*��W��RI��i��)%*�(�(�UU"I)A��IP��H� �*�T�H�B��$�H�$TQ(Q% ��a�T(� F�Q@�*%%)�&���*R�E)D�U���
U*(�T���UE%JQT�@HJ��w ��*    m���m��Z�CY�RI`ͭE"�U$�mE���&���P�a[i4�Zm��2M�[j��J�P֌��J�*��)Q��   �t�@c��
t(��p�jC8� ݞ�{��:�@(�� A\�@
hw�֔,�p�IE	�w�CwRHP)%J$�
��!�  ��i���87���e��v �j�u�*����5R�9�C�U+�j{���҅=���킛�e� hZ���*��J�E$�P�(�<  J*���9� (u'.i��@=��:��հY@ j;�� 4�R��Pt6�����^�S�҇A�p�t�R��U@���UUA�  �p iٕ�wt� ]Gu^�iMhڞ���.怐)K��=��G�� ��㗻��ڞ����2 	Uݠ(�T���V0J����  ��
R�,�$T�ʮq�
�	ùҀ�����@S;�a�l��N� (�]���Sjfڕ#ZU�aA� Z����T�T!T��   ͽ�JJ�� ��;��m"�  �L  �w��MV�
i���`�إU*��(�
��   p ���i4� c@h&� 5� �0 mL 6Q�ֵ�F1� ��P�
�T�C�  ׼ �6  l� ��5SA�  ܦ 6U��i� 3"` +� j��I��(	)`  �� ��0 FF��ej &0 F0 �m ���@�`)@a� )��      L�)U� 	��& )�IJJ���L#!���`4�%#F�	����e<I�M4S4�B)� ��j�      Sz�U&���     B��J*� �  [wl�ʙ_[�n�JB��Q�(�I�6�¶��j�>�3�w:���UҜ{U��� �f��%��J��@U�� ���D]�(�Ap'����O�" �Ȥ�I� U���DEó�5��2`�%�.a0����k&�k&��k&3�:��:ìɬ��3��&�k�k�k�3����:ɬ�ɬ:�3�8ì�ɬ������k�k&�k&���k:Ɍɬ:ɬɬɭ�������ɬ�ìɬ�Ììì�ˬ��k��&����ì�ì�ìˬ�0�&�k&�k.�k3ɬ:ì��k����8ì:ɬ:ɬ:ã&�k&��&�k&�k6�����k&�k�ɬ������ì�L�α0�:ì���ɬ���k3�k&�k&�k�k�k&��&�k&�k��:�c&�k&�k&�k���ˣ�k�k��������&���k��&����&�k&�k&3��ɬ:��:ì:ɣ�����k :¦0��
�®�(k�*¦0�� ���.���k":�2	�(�*:ʦ�� �":�.�+���2�� ��Ȏ����k :Ȏ�#��
c:������:�.����0��)� �
:�����
��2:�0�� �(����� �":�Lk������k :���	��k��ɬ(�����)���(������"k
̡������)�k*��&�)��k :ˌ�k"�Ȧ�������*k :�2��#�"k�¦�	��� :ʆ�L
k"�¦�+��� :¦�#��k k*�Ȏ����k :������2���c
��.��k�����(k
̀� ����#���:ʦ��1��k:�������	� �(�2#���	�
���":���"� :��+��k*L*�:����� ����,�.��(�"�ʎ��k :���k":�������*:ʮ� L�+�*k�:�)�:�!���:���+�.2����(:ʦ������0���
:�.��� �!� c k*8�������!��ì�ì���k):�ìì�ì:ɬk3����ɬ�ì:Í��ɬ:ɬ:��:ɬ���:ì�ˬ�ˬ�ɭ3��:ì�ì�ì�ˬkì�ì:ˬ�����k�&��.�k.�k:�0�&�k.��k�:ì:í��ˌ�ì:ɬ:ì�ˬ&��L&��ì���k�k����Lk��.����ɬc&��2k	�:�k��:�k���k	�2����ˬì2��)�:�	�:�;���2~'���
������]E����ҁU�`���Bl6i�4/���l�T�߃8e�,^廛wW�qA�0D�R"oc��]n�#v��B	fmF"]��=E�a��iѺH�"�i��e2(��Ɇ��IlɦP�T��FY�G]*|a����y��
��a��3��kڬUu`�I�.��H��ҭY�H����h�����M��H�n�����4T{R�!:�-3E�E	��m�[��5��0h+5k2@������e=��2�'Z�Si��t�����ʕ88�E�a���5U� �:ҡ�ۦ�A��5D�fQUt�S6L�E� i)!�QԪ캣R��M;k��&ܹe�6�h�{p%HH�x`TԺ�!i����P[v9J�7{[�N#�컎�ix&Cz�j�A=�t�B�\��rӼ
I4�.� m���.{�)i���U��8X��Z�Q��o.��[D�2���b�z���{ws
��mc���`̦-��TCor��h9m̼U���j��"��ج��(S�
cT�Y&,U��f���j �k����{��q�r�����fat��Z2*fh�Y�X�����$Z��ci1Xo�ݭ���ũ��Ry�D0�;=٤	+$U�4��j�%4�Z��ob4��l��B#�6�괩��x2;cq������1JJ6��1C�WH���^�廥Gb*����l��C( Uz��`Է���R�0�nD��6.]��ɼ�n��}Zd���^��e�!���K�������)<t���'�V��ɿ��q�P8��Q��M�t,v&�T ��e]96Z����
�L^Sl�l����+N^���O��ޕ�Z@h˶!�%���^Њ����.�\�J7�1�bMXB��ַٖ(�xHf��6d��4%��A�c�߯#cf�B+ɸ�Ǯ���8�h��E�M�r���®�R��ת�Ţ^&ݺFʰf
�J<փq�!ąnk2<B�YJJ T�KfK�-n'�4��)Nb�y��(�a�W.1@TR$��]	���n w0+�h]aҪm���7hem��2ʼ�D(D�8L8i��Zn�t�����W��R���܈:�(�ȋ5h����KV��ya���M�r���iL�n��nA�À���Y[��r�Ad��0 +C_[�l혅j���e6sl`�L=�J�͠�����1�F�x������ Y�YJK�
�rmG��L���X�u��H���)%�\��sv�����:a0�Z�h1{�F����)�V*8�[W6�nƫ�(!(��yһ�N:Gt�D�[n�\��S_m�e���j�f��8�QGs)�2
�p]%WvX��жfo͝d'P��u�4좦�ㅫJ��R�wDnRj5e:l"5��-����V���X���LU{V���Kl(��:4y4.��j�A��V��c���[ٕ�l+*[�l|7`4h%2�Ի�h�W��1˵D���AEf��uk�~�!��-!�b�����B����Wm�WX�;-���7(P����CR�hQ��ݧ��F�'y[@}1�mc6�J�ti�QቶV�k���9%A5��c�Y�����QۼՀDfRF�g�b�^,+�-���D�ڴ��p�*�c^1"5x�!_6D�E�0+:�f�a[��e��.|K�Zb�|���VZV	U�1�)7zݠ�U�2}�����֢���vlZɳ~��ayz���4j(㙦�1�&�%�U�4�-e�+e�XV@�k%�u b�е%�����n��1Ӻ�"�{����Mص��J��m�x��
Ò��k��F�*�I�iG�b�d�$ͺc-��ҐT$3V*տU�Vշ�����Լ�4!�7j;�h:RMyXAW�n/QA�W������IY,�p?�W��vZ�̡�)�Ӈb�z�j�H�H��޺��wy54��U%֑xC�jQR:�gk	�6��9�a�Հ7���ʒ��&S��]��Z�ܫPb'*�8%�CfV�� ��Gr�֫�%�$���ZE�̈́��ެְ����P19�Xk&L#h�vDν�R��֬�����z��0���$���;�i��@+a�Sv�X+w�먋��nĉ�u��L�%�MY��:Ueۺ���j�)����Z�e��mk;�Jl��ͩ��-Մe�J��ʇ쩱�h<�f�����w�^��@��L�B��������*�G%1t.�m�"�f�e�wr0�U2�X"��M����,L�E����a8e�����޷�ٵN����7q�*&��TݵM�`�"~�qʼj�^R#*�ǆ�Z(�Q�5kE��V���� �h/En�w.6>oq�l�h���I���UP�ș�n��ydkj�)�ۣ�BM�ut4�Tc"��>s+k^[;[M�y����{v����Z����K��VܚJ�*m��56������3Kȕ1r������U��^P���*� i�hC6�K���8�=�^T��Z�!И��)c�ŀ�g^Y����7���]�cc�'tܻ���g[t@T�wka�Ld��)���x*9d�N3.��f��a�Z2��wwN�R��ס���v�f�GUgt��y���u��J�ñV��Fn�FՀ�Z�ܘl��/l,X��Z�Mva�j�
I^���5):�l6�1�w��Ԣ�S�S���Rj�A�����m�A����Yʅ�ǔ 2�@uޣ�HY���S[��t� J[(m
ݣwVAcPM�(i`AF`�ot�0��a�n��c��h,�[R�ܬr۠U`n��e���KbSÊ���0⎮����8�F�g6�z�l��PҧW ������JH̊��@m���������jt%�*�M���+�x���pՖ�,�N(#JC�Ђ�'�jɳM,^��!+�q[K5�zpX�U0��%�:q�ӕ&3gef��zu�%nv�xv<�*�f��u"� k(�J tPn�%,������[����tV��[㭭i� ��tn��N�۔p+����F��ժ�im0�{��c2��-,$�&�G�R�k0
���lVB�F���qS�F�����qh��y�,a�,��`m��-	D�	��w)�r��.S�M@1�j�ܓn,U��vd'h^}�	�f�	m�)C���'j��v/a��u��X���j�-AB���&%z�h��6ƣV�%p@D]�%��]��n�N��kA�oZ͌\"@�F<4ن���4�a�y{a��Q�Kً(V�hҦlH��B��I���x67v����m���)�]��a�PM����*�b�Gġ��*B,Y�TPm�Qj2i�Y`�w(S�n6*�ƻ�Db7Y�V�t�*�����{��3�"	Xʲ-*�XՔ��F�X�6�n�W�"�����怈�ۧbS0Z�.В��ws6�2)�N'0T�z�!Z�̣+f:����h=S뎪�iWOk#�e�,�f��H�w��(�+�U���i?��J���!U��V�j Q�T�� ��4
ͬ-
Ѕ:U{ZQw��/� ���N[,�Z��ݍ���E�6�an'P�6�?�����M`���/M<�H�`[Z)�t���杊R.:�B��l�*w��&wb��yn��a7�<f����KR�(�RB<8Iǟd��0�4�d+Ss�n����,Yi�ԃ�W��B�Ҭw�|$�,+�p����R��v�ź(�P��6�>;Kjs٫ �$E s"�ww� �{*6�@WS(+�vX�G+�J�u1Rݫ���H����d��Pע'S�2� i-73f�[ �T��q�f#���/�V�,��r�!�aZ�w�Օ,��I�A�	L6�Uc�C�k5b� ����,Yk�a�XfF`ԅK�������cF��oSq,!�4�k1�f�)wb�T��ХD��H�ѦR�h�0š�0�hR^i�j�t���G�nV]�C�wx�uzb%�aN��2��r���=QK��5���.�͌�صqe��'mV�bE�B-R��Z��
�8Bt
8�wfʖL&Zѹ�1V��GubM�eQ��@j��M���.�֊�9���a��� ��m�x�!�]b���B�u
v7D�,c���X�S:.Y:�B��"[AX�Y��F�,g��𬴣�'K��7sT7��i�$�ڋ�ve����5E���o,�I�o��T�Y��Sp���[��z�R"3-�T���h��1l�4��	�Fe��C��*�mȭ�&�T���+r^�b�c����m:��m^�11�JMÂޭ�*��(Әr���	�n��p&⸠�E�3~fM��GWm�YIk&��n�t�9L]�x7fhƆ���ݺqk@dwE��a��#(c����*���N���պO@l��j�d� �XDX�b��E7wv"�T,����R��ܴ��է5l��Zn���B�,%��- �V^F��e����b��U����K����ԭw�NR�i#]��ݨsp`ԫhT�����|��)�+\��d��0���ys �5L�[I�ɛ��P���7��t��tw3�h;�v�
�/ )��d�t��A%E��%f̧#�b��4��`��`����B]D��4��yy���1�R�Ƴ���k3��Sʚ�M�%Z����B�x�J`���כW������(�є��e�\y���C"�ʖ�r�ݒ5Q��C��⻁2�j�
�,Y��m��ɛR�'�:v��ɖ�����
˭�7p��`�b�F��u�r:V�2��y ܷi*�5�q����uXQ'����̖*�I�I��مڶ�˂��1���7���@�T5HԻ�&i�����D-56�le�Zw�G�m���a�5��l]��i�<M���`&Іƌ@U��C8�Ӽ�	B�3@`��e:F�rQ�H��,����	��z�[��R�!�{@��7���a���fݦ�;��R"O�Z��e= cVa�.�>��}�@s�Z5�6��w0�T�iZ0�4f�)}����y+(�d��+�:�*��Nu�!,,<��a��֛uG��ދ�Wf�v\"��2Im�ڸ�Jږhj��v#nG�l����\�$[5(^?�R�Վ˼���c/@� �.ݡ�P��>u}󬮑R�EK6��ֻ�u�D
̧��7���Ea��FV�J�i�3���r�^�z����ZQ��%�P�j�M�j�eZ��DW4���Z����w���5�1�]��Pؐ��t���Um1Wl8��0ևf�!n��v�]�A� R�6Rנ-(v5c�q��s�Zz�=�f��e�4LŢY9'-L���sp(�|�ҩ�7Q*b����^7�4�f�AW� ]<�z�FJ�
1�џAw�&����:��|h��*�	ĩ'A0�H�a*�"t/�m��w-J5bb�S��JZӓq��uM`��X��D9AZb��pS��7``��7-y�Ff	IP7qbӸ�ZH�$T�X�h�^�6ٌ�8pI]nДoC�f^��Z�#t��ɛyy3)�����A�X&JQ��1ڧR�T��c3�c�Ze���i�9�
�k����Q)�q14�u�X �ѵr[)�R���5��nG1�M���bedI���6b(*�;�Z�7����WD�u��U���v���}��	�74��YVd � n�6]�]���R=�s)��R�^E=��@+�[X�l|�V�V5o�c�:��b�L��V�ͬ('�.Z�t�:7l}j��V��2�HZ�w.΋�Ƴ��T�x���i�J��������6�c�cv�4:���[�@Q;HLQSY�}u4o`ϯ6 ��+
��#�����E�HP܇�"�0�8��M��!�b��1ut��浔��ߥ0�T��sU�.��&�Ы�sSWW	X��bc�Da�㠵72�F�>��	jar��[Oe�ph4�AP�Ȣ���4j^��H2�Qӷhn�0[!Y����Zt��Y������d���"4=]�y�(ε ���J�Y�m��*���k�D�k	��z���$u)�Y�T��G�ǅ;��۽��|}��g�I໨��h-B�U��+���j����O7d����`G�޼})�Ð'�NXŗ'����D%�q���d١�چ��V��ziZ���4%^sP�P�������GQD�5î����>��G��:'�Z��j�D6��Ӭ;��I	<&�L��Y�_�׶�	���\����o�uHlv�"�4K�����ʹR�ۧ�U�uz�ߞ��RU���.��_���S5��JRW��59)����U���QVlW�U>�sO\��]���F��䌃��x�!����.񹆃��C�2����� ӃZu��)��ÿ{�=��r�,f0D�D���-}�ۇX�yf �r�������E��^�oN�j��C��
<��͉�PV� bd-)�:#�枳�-�D��)���y*��[�����hZ/ю�����ʓ)	�r�<v��xe�����;��tV�sȏD~�1ְ|�`J��=���g޹M�W.���h�D��W�V��6��W�y �5��E�+��"K�C����,}�����Ε���ɠp��Y&�Qp7"�f�,�!e�0�PDp�S�>�}�tt�L�8S���꓿�Ҟ3�o��n���1�7Xl-��KS����
�����!Rи�T֠��^�z"��]A������Ob�0��If�w�h�E�.�b���0�*R?ow^�l#�v���7�{�2O7�=8]�`�޲.`��ya�K���2�x��Oy��P��iRnFi��w���a%�H~tw��=��(s�:g`36
��#͈8PF�|�l��WkF�`WLO�z&�r /E��dх+�sm��qz�/r{�G�/ꡗ_���/-�:u�-�;�&�L^��¶ի�&w@�m]�hfmu1�Q�t������g�oW%;�8��ed��.7�]���ۚi�~�����W�Ҋg�B�٫�A[)�j�n���u݀;ŵo�t� O=����i�&.�Θ�J�i�
݈�9��k���S�W-�C���OJ�l��*��X����ݒ�3�jf�t����78Z�LveD�㬘�V�y,;:f�̗Ҷ�E�*��N�h:�n�T��ǌ0�DD8�N������z�u499�/le�������^��b����d`^����E�hkK�t�H�ose�D������&�^}��v����Xw2q����MZ���v�R�=��	mmi�s���ž�S-��1|��ev�缄�q�����ۮ�l�X��5']m� �	��<����J?:�GxJZ�]�[�4RT6"�@"rz�p�J�_ǻbݕ.�O�T�Ռ�|�3OA��ҥ@�Z5�ҥ���R�D��҇3S�<bN?pc�ൢs�W�7?�K�t�� ����"�.]�I�E�Vfn�����fsݶ)��-�q�6��B�5�sW|�[Ջ�W���u�"�dJ���D:�|VfoҺd�
�YB(6�Im�޳�S���0�&=�;e�	h�ژ�k�>��JTK�rwJ+���o�	�p�=�jg�o��������kau����[��TZ�yn¤Y��ރ�����(Jz�f�-�ٲ8g,�Pf�f	�N�e3{�)`C�մ��&a�\��d��]^+t0���;�B\�S�і�KWt�6ݠ�]�7���Ȓ��2���	��Sn��檽T^��sL�7I��l 6�\5��:�
S���H�wڴ(6��.ٗV�DQ�:�R��KWP��2S}��}��,P�E����#��rI��P�\R@C'j�1���P�aE٣ӗ�)�/fzk�=�Ͻˏ@4�J(���G�t�!�)mj봞l]����(�2o,����(Y��u�-n���|�
�p�i�^�%���^w|w�EF�]l���Yr��^�]`�$C]fC���ɔ6�5yي����P�Vo�i8z�=����+۸,�#݆�F��L��CD.�q�i�f�Kz;uh��ܾ79�jj̕jP�����O��v�˱ʺ�ΛS�V6��H��l��_j����nң��Xza^���Zƛ���n�J
��Q��=����3d�%]�I�H�:��p�� �(ri�q��ZN�;�kjf�@�x3ڒ����o�����O���������,�)М귷N$#�2�v�l%�A&Wq\��A[K�u�Vz�PUdD�<t\L�`���r��M��uLfeJ�UjW{;)�y�Ϊ�t����;���$5��e�}}�h�::��0G���X֑��a�M��$�|��዆C+e�u���󑁕ݲ�	� �u'.U:K�u�>�����7��!�s�˦���`fv�S��rPB]oQ�Uxgi-=ݺ���AC��jp;�h�4U<*t�Q��//�e��w^�=��53�R��{��f�HmA��)��!t�f�k�i�B���}�步O�d�;?-S˦���J�>����t�0c��k/�4P�Xj]�}P�J渫#�z!j����(R9����N^O��u�w:���WƐ����&�u�(�k��M��^|8�:�Ӡ�h�Y%:`ҔzW5�t�WYY�C)�jr"�`���]��Q��MD�]��=(��M=]�Lv.1vR�՜�9�����sO,*r䝡u���d�w��Ë`��0rڲ�$��vk�G��s�=C�,�z��o��2���v�Y�{�A���WYIX��X��)ɲM�JU���z��:5��s��x7�RR������� �Է�9{�)xvﷻ;+2��c�
���Y��4��ueup��e�i����u'���^mR��窲��˃[���[��[�g�ԛi�'�K(GhT��S�a:/jKUnvw-JIV���x\U�����{�ig5�3�Ω��IR���m���pf����}�t��X7��Y�NƔ�gn�p�nvM�iXU�q��:zм���WfS�Χ&��s��ʺ���JF�b޻}S��xܺv��R�2,���������ں��AJrЭb�˶�P�!Hq������9w�����e��jk���Գݛٙc��H�ә7iOr���,��ΦrH�Nek�{ʺݻ��Z�ë[��@��N��^Ʒx�����������YW�,&�ܫLT�+xM=׫�-iU|l����R޳����S5�5IA�����.������HL�U���Vi2��݇�4�a�3+&<u4x^��Ф���7��uU��|,,�6��w+��c��1iF��/��n]�y+8�B��ab;m�^�!��ZԎw1��+��u��`ǹt��v3��b�䧇��c�T7����#y��S6k�Ť�^�EJ�Վ��tްq�xV�������v�2�f��6�fПF�1�bV�vIk�-ʅ���A�h#Du����{����4�R����VU�B}��9x�{��)�y����@��.�=�F�ɺh��h���W�Z�.A�� ]�9����ċ�Ve�$�b��9Q\*�����E���[��lkN��N�V��;��YV)I��b򺮹X��9m]C?#���g1��9�V��j�j��es��XU�t�t���U��3A��C���ɤ�|S޼�N���}*��:_j�ff�N�s�(T�/[�jG� V�-l"ҶkYP�rvv�k^4���������X�}�����M �����W�/	�����d,d�7A�[}�g8���x���rҸ��һHwj=,�E(�v�����W]Kv���ζq�T۴i�� ��V+��R��Uۆ#λ���h����ݫ�u�������7ڈsy�;{v�l�L�4�.�1��R��re)!�Ҧ�����ê
Ժ��/����*s�@hlԊ����Y�r}z�3yeN��{k�*Wѹ�W[�����*Ȇ�cu�u%G&m��&PK�;RܥOk9A¬�c���XF����u�]�ƒ�-�z�1[(f�����{\�v�u ߻2iV��8�tV�&�{�%��"d�Vӫz��pчiZY�kzT��;	��u{�sSBj����yV���N��fnt��O�N�Ǧ�us���M�R��������{]X,4��ڣ�@�_\�G�2��ù#� �&�ʱp̻Rs�T9T�&�#�a4k�8��cႻz�k&�ƇS�i'	���#�O��Y6�u;sg��B���Vu!�^/�4���,й�(�D�:��t*�uh�M�@�8�k�!��Tt����H�=A�67KgM���WQ>f�X�L�-{�i�:w�֫nl3q�c�����'Β(j��l7����ޝ�U�N�r������ko>ed���/yh���45j�8X�=yV�e�a��隟�8gZ�uګt��+{6�?�ɉP�ܵR����l���3������=X��Z��T�+U�$c�Jљ]��ڗ١��8�nn�o)���γ�;&/�3�rF�k����wh�O�3%CH7��\�6���S	�w�`��^Md�]�4���e�R A�� �c�f�.Oo�B;�"[=�6�#�c{e3�%���	�*�v�����u性K��tvwm\� θ����C���:�J����y��6f��;1"&q�h�:��X�5�	ܧ&p��w��됁�JT5S�x;Wf�
��Ѹ���JY*�k5u{za�૾X�(��tӻ<������+�@���h0��d�T��}|G]���B�#�fj�Κ�Ձ�:۝�0�m�����Pq�/K��.��U�7.n���>�3��&,o#.푻z�&fwb���Ws��<VJ#ǔ�wR�C:iT�|o9�D���cG��Q�]�d������� �={�X�]���.�k$�j.�K]�Kl;����Ls�yI7�6��m�3H��1h�36����*SX�Wi��=F�BR��:�wd�W.�Fiө�� �O�����5���W��(���=��2�����&�/|S�]���t1�eo9lu�4����|���.��l����R�\T�mu�ъ��b���u�]6rK���k�^������Lƴ"bܵhV���WVqՑ��w�fi$�Ez��*u�S	=H�w�2����m[�:����&76,W.��ް]ǸPx72�q�����hҺ�
|J3��Q-���w&�b��<��Z�
,��iv�4Z�U��0U���Md�\[�j���K������VR<J޻\��p�`\��S���Wx��
c�����������t��L�yjD��DW�&7[��o*��͗��+`lW1�#�C]�]�T	�l޶8L����ڋk"��HǊ��������[�M��`�w,���Z�y��jJB�{�,��w�,TL}�-��-��'��M��z�^��Xq�S��7m�{�/����o"I��vi���;�01N�Ke�ZruEvi�
l�I6��s�!�6_u$���^έ�؍o^�|*�9W�������r붓{��NZ���	�d.�k������.:5��s�����,/:�����Gk�����7���q{�2�qf���]n � �A�!2��1�$CE�D.�/��F��^Q��B�����MN�M;2"JFw��!N��*zY���wtٷ�ݕ��n�c�*ɮ�z��ξ�Re�Mˎ]g�|�]NG�4�7b��掘o��4uǅ=�=����`s&�9��A�9����.��R���'YϚAlko{#l�3l�3��dU�9�/��n�ՙWW�5aPa���(��.���z����V5N=Z6	�n��ٔ{Eh���������e��nmm��t��V��\�<����Mǰk�JU�C��SS������J���V��C�{�d��Zw}��X�P尫�ˬpe�19QS��v�U�o`����a�rVM]ǃ�Z���o��GTq��\�S�s��}���WIW�N�r%H
�a�6�vm:�F�fҳ��fe3B����f0ۓ��&4�p2C�d\N���T�r�f�3z�gEc�:�ݡ{\B�wK��:ʌ��=/��r]���j�7{�J�(G�u/gn�i�t2��M�^S���س�JV2)����ʳȼxZ��k�n���4q��nή7��-W�3M]���y�LBq���6n,Ͷf��d����W=�2�S���iE����Xopw.�9��*�֙������]�FѽO�L\U�=�i}�(ͭ����u;�|�4�����*:���Y�G|;0K�9�#���Sl�t�Ƴä�*W��J�|�1n�/��!�a4R!`��PWك^5=k5Z����dƒ`�s}C���ޮ΃rq];6o'o �[�����ok�7��5�oSܜ��\�=������kH�n���p�n[Ml��-�ţn���Y.�j@��s���(
'a���W{1�X�S*���A��y�D�e�RBw^�� ��{\F�iˊ�*�`�q�+�0^���,�Ɠ/8��>*�UQ��I�\Ȼ�Z�z�ؖvi�=*�W_��D���u�̦�"Q���4�ވ��rn鷹£�KǗÍ^'��-#�b�F������+9�w�-9���%�zq�	���%�8>���2��[o�n�*��g<ͺn�t�+n>CnJ�W]��xmv�1��J�K������E���ۮ���Lo/{Ս����R���E�N�}]���]6ݤ�W���9�ڏ���p�"�}3&X���2�;wu��br�sܫ�.2��� ��ik�}ǉǪ`�ť	��8����j>�rK�f�]��Rn^%�`��Ҕ�npw ����;��:�5-8�={[ȭ驷����m;�Va��Ǌvk���U���\��#X�=9���u�-�WY��C:��z5|8ԋ�uv�x�s�&Ƃ�G���t���U�����.H�m��bȻ��%N�\ɛ�9s�E�M3�\1A��w�"��ޕ:�U(����BHJmv�%*���$�{��8#[n4M!�G�?$�n���B�'E�D�4�B�Zk��[��j���J!FfK�	�@�! |o�UKB�h�Ce��c& �Zm�4�MѦ�%��(��¨Y�}�V�\�g"4I7�˻�q�`f�?�)P"�7��%�M�IQ�lR��Q���E�$?7N��i֢�R�G��U xu����I�
I���`�TS|�h7*Y���I�@�eYg%�*��hR��8�1J�a�H��V���"]�XZ�.�����L���t{K��j@��H�T#X�?~�>6\p"*P/�%7�˂�k��L_LnQ�˘lp��s����z�ʼ���ڲ�ʈ��p�_��Z����K��P\0`DBu�v�B���3>�*�u��i,�@dTf��&�k�� �A�B�Ti��*(��N i�u�A�g����(2#򽩎�������l�t.�h*m�H�r�4]:N�4	�L D�i��	��6C���CJ�R-L�����5��J�Z��� Qݬ��x "�`a��iUOpfD}�@��yl>.���B�����~ �j�����]���G�U�ڰ�6��J�r*�Os{F[&��KG�d:N8~PS�-	��.V=h����Ͼ��)�ؓ[��2r�ڭZƹ�7&�#U��_�	c7}Yv�mȆ���T��
�ۍn:�y&AB�l�h�&ݳ�ǯ�\b�v�Ш�h`����i��-uM��H�������#�`I�Ũ�����F�U=Kh�r���k��i�S�wdЏ��"�*ٝ����ݑ w����,}�.]F�̨b��ީ{�*�.�q�+qe}C�J�[;eN�û5�nJh`N���lWȠ��̒'i����J����wC�z�v�ꪬ�K��o��'�T�Ï%�%�i�![�������)up��	իZ5��\ye+ɖ{s}Č�6!W#jJPWk�Om��L�)��L�u�E�`��2��z>Ty���ݔ��9�6��$eT�cS7ӫ\f�Ɲ�j\����-
�nN>���"�Ǖ��h9�cW��t:>M��0q��ӷ�ڎ�3�Dy��^ҽ�Χ��7G�T�z%s4�)�1V�`��؅��ۻ�ش>ڴ8P��������2S�ݸ��ݲ�V�d�Xso��g�C�����������ǯ^�z������ׯ^�z�z�ǯ^�z���ׯ^=z�ǯ^�z���G�^�z��ׯ^�^�z��ׯǯ\z=z�����z��ׯ^��z�ׯ^�z��ׯ^�=z��^�z���׬��ׯ^�z��=z��^�z����z��ׯ^��z�ׯ^�u�ׯ^�^�g�^�~�_��������ׯ^�z���z��ǯ^�|��yq�}vG`����l"X�u�eV�f)��H��N/rw*5�U���(��dY|���@�r�g�=g>�e����v9�`��.���c��52��fA�*-��.�rm��-�:	�n�4/7_<#�=I��Q���j�mmh6�e��6�@ġ�t*ޭ�]XVd�Y�W�}R�����z��:x_}��E����[��+�2뜥��Pi;����T�x//��B���|�j��5�v����A�[궍,����i㷸�'6$i�� �g�Ɍ�p[��md7.t�g_]X���c^�S)��i�7�WNf�����z��BJѲ$u��%�����ؕN��ى�a������,��K�'+&��7�6��]�	r)WĆ�_Q޽����@�0H�B��6X�1S�&,�i�;��qȷ��]��f�|��өɷyh��{����]��-}X�Ւ���1�&I��c�;'��w�s�|s��WX��ABq�.N�)]���f���v���ۻ��	'h��}��6].L�o�/�VY-;*Jߟ��m��RWjk{��"�F�έ<�V�|)`ud�xΓgm�hN�v��H�}B;�lF�c�(ꢙ�y��f:;����ϛǎ>>>�>��z��׏^�z���׮=z��ׯ_�G�^�z����׮=z��ׯ�^�z��ׯ]z��ׯ_^�z�ׯ^�z���u�ׯ^�}z=z��ׯ^�~�g�^�z����׮=z��ׯ�^�z��ׯ]z��ׯ_^�^�z���ׯ^�=z�ǯ^�z����=z��ׯ_^�z�ׯ^�x���~�~�_���ǯ^�z��z���ׯ�z��w��XDs�¸�E��i9��󵴳/kF�O��;�Q�9�]�Lu��ͻ�=����GOI�f�CO��e!�^D�{�ՙ�/��ss�.�z�-.��Ӓ.o*�Y8[:�d�ԫ�@���Pb�ɮ���Q��e-ǯwBhw&��i�p�g��}�hG9�ƞWu:��}�Y㦈f�(��ZAILU|dd{��Y��I���+F���X��X#p��ys@����x��M��	�ܙ&��`�"�.�5�6�M��Vt���|y��|��3ja���}z���-fw��xy��s���b`ۂ���:(��[Ÿ�F�U˸�� 2�Ռ.J1N�f�&��om��o�[Vf�1�J<�ʹ[bB�Gf�[����ό��ZT�]NqB�+'�����RW�T	1�_�v��.���|�u���$��Æ��V�ԌY�n�\�y�uMS:���j��^��Wv�1<HQC�&�#�2� �U�d"/q
숒:",�P�y�n�n�cԻ2�u�0�ƦWvɜ������Z.��$M8��n��;�k�n������Z*I��**�2�/z^i텔=n�ʻ��Z�7�ڂK�j�f�V
��|��|��<��ׯ^?�G�ׯ^�z�����ǯ]z���ׯ^�z��^�z������ׯ^�z����^�z���ׯ^���ׯ^�=z��ǣׯ�^�z��ׯ]z��ׯ_^�g�^�z������ׯ^�z����=z��ׯ_^�z�׬��ׯ^�z�z���z��ׯ^�|z=z��ׯ^�~�g�^�z����~��~�_�ׯ_^�z�ׯ\z��׫���_�iqX7o9�;fu�=u.�u�;(�S'�B�VLߕgx�8����g�U���Ш�+8oigAX���]�VCʴpZ��c[LIՁV�WQ`#�kbͧ��aԪ�5�[Lq5���.�3�vթw'��})����K��� �^�u�F�\�c�C�^�F,�u�|���@y:���*!���W+6��V��I�@��@�G۽.[�F��z�
�>�-�o�����\����BBi�FE�e�÷�fMY�]uv�ǜ��i�B#H�ҹ\�a/��A������֧����i'O�/[���É��#����wrU����k�V6�2��P���픇mko���i>��Zn�4#��^�[�ˁ"���(=7\2�����k��i�1��wGn@�>��� FtY$�Y[C����e�**�]F��.�f�t+����H�&\S����z/����kX�[eWm�v�]�׼���R�%����sr�.E���e��)����g;y��E"tSd��^Z��\Uܲ�awf�Cu�M:w7�c���g���V����]��	ɽ{�=uǆ]4Ļ¯qņ:=�.���&�~�4����Z3��p��PZ���V����0?�E���>��	���D1�9�- �^�!�,�x|y�|��7t�s���ߞ��|"H��t.��ƞժ8�=�bh3�>�ԺI}_�n1&�\���3#U�Z\Eہr�9)��k?W����&�G9Ǻڦh��r��Sk�����o�a����Xn��Fo2��q�Z�$���t��\�˨N�B�Õp�l�,
�UR�4�.����u�R�;�]��,���ܘ��y�w��þ��)
��c15G��k�Y��.��>���}�*�6�f��J�JX���7wko���b�{��Tr�.�`��p�_�*җ���h9w��1I�����Wu�v�JTs�f��>ѕ��/ot�-�)�4N��d�&,F���q@��)�6�ȟ�O>��r�ġ���}Y��ܩl��	�#N 5���Wˑ�Ż����&��m)�w����+��gŅ�K�u묶�j*��ղ�G't50|��ծ�\4���;)��뎂w��>�&����%�;�7����u���r�d���G�H�#U�@ܻn�]<,ǝ�gm:��x�X-�|���4>��}�����m0�-_#{��4#]zU�Ʋ�}��4�R�_V�Y��j=C���o��\N1��s{3i̚8-��U-��Ȯ�c�i�ĭm� m�	�B�.�K'��h���>���貮��44"b*�������-��2��ch�+�g�S)����*�� �F�:9he���*��"2��C�������2
J୉}I��7f�������}���!�jy��V:��X��ww�݈��\�7��Ay*|P����4$%NDͮ��^���$�{���D]�ԊT���T�Z�V��n�U��wJY�.hU�N���S2$�u\ONɴ�J�U�V�[Pa��NIM�U��;�U9�"`�/���!����]3��ݑ�ij5�uĹ`���%�L��ãf��llu œ���k���Nmd��s��{y�o����*�e���t���]���v\Cy��m!�+��S���n�U��gj�f�v:�TKB�����|���b��\�Vf[�Mwm���u��Koa�J��|]8R�����eKC��Ի�z�>��T��ᛀ+��1-\�ݴ�n�����Uz�;Kmcw��4-��Y�B��79���f��8�dx�f��3�QqulԐ�z�_N�w���@3E&�q��o|fJ���m�gm��Y)�hm:{ˍ �Hh����#�v쾮�se3�n�m	}}p�ۡSRx�n�Yy-N��%�j������&�p��i�8I�n�U��kv�_|�W.Ƿ���Q>S��W��4�˴�C�m(T���\MZ�m�5��\~�S�����&�s��Ra�خ��-)ۊ�Ü��Eu2�p`���,��sP�;W�S2��P�eT��d����Gu�qAd��weq��W=�Vsx�9�xok��&m^�}M un򶨔Wn�B	g��Y��$�.V��A�ikMg_[׷��v_d���K:r�XՂ6S��{��M
��u����d��ΡY!�.C)�m���Ҋl�0��mj��"K�`T�wm��pgd8tL��3t��*s{�kh�UU�Nn�C�J4���{�pQ���I}��}2+�����'fb)�h6�+8�M�m<�tƈX�I�T4���GKH�u()�e����㾽\�ֺ�P˼�������5�"��/����8r��c����G]]��x0y���M�:a]s;�\8�D��y�m�{.����*�|�{J����8�̧�|�X'�m�j������]�� }_��WX�2�1�S&Tv�jwk�����xz�b�q����g�X%��Q���J�����˝v���6�U;s��*.]q���\թ��[�v`ͳrY���e��4�oU�f���U���QZ��k�	j���m�N�g
f�Sx��Ԩ����w����#z�Ӵ-�u�P�,�/�&F�b�����Bł�EVO��z�0���PRW�d����@k�9AGG���5�Jh�{c@�{a|�f���{�1�;�J�*�ېg;]j.����<`n
��1�������j��.Js �tK�0�&1��0m-�OP�	0��{��fN�ڷ�0<e�J�s��iZy��(��1ڡ�i�6ͯ��,4��b�:�V��� ����kͮ��[��îcy�f.U}0�;FoP/J��5�U�fp�L��^��g]���8D�o.�WK�^��w��&��z>�v<P�������EM��Mٛcd���1��E��q;FV\qn��];\V��58;�ٜr-�Z�~ٿz��p*	]/ �N�w�4�t郴��7�c�b��i���Vol՛\�f4�V�t���5ۗN%�8�=���j�K���v��vP���;(�z���p���3ض�|�]`
�o,4T�:wwSY��%s���Jwyy�ʝh�M��g��ɽ3��k,nVvʘ.��Dk�a���T\��v�R�.k-N��8n���4:���i�c���y����2�&�Ʃׇ;
�xlH����+9�|�f��l�*��H�%ˀ�C��:�w0��_���2szIr�S�İ�ULᓸ,�jEӹb5�F�V��l�u�^0�9�\E��)F�8�3y+�*����N�5������e�v�7�nZ�̵�[Xb�&�˩ ��1�a��_Ў���?*ٓ!m3�ev8{c}r�eRj�	��G��غe����L����|�i �e%7i�o�o�ġ�VW�58(�����R"������P�^嶻J9tf���\H�5��CT�m�;]��٭�Y*����mu����"�5g�l�9��@9D���xDRvoNcork���J��D �7}����IF7�pN��c��0Ɂ����t�S
������{	�W���ƺ�^ͥ�^�s�x�{ٛ��X��Pg	��:���l��eN����X3�l��DYw��Y�+sz�-h5}��d�B�aQ�0���K�����ԫ���A��x�!�+�rc��Cm�t��p6�o�eWf�����X�h��,����)�qSnԣ���LhTʛksr.�x�˧��x��%'�i���R�Y��JoJ�S���|��V�7ُ.��Ӏm:�+��/	Y"n�!�����r��eCb�ۨƭ�y}{��;��ڙuڳ�,ѱ-��Q�V=3��p=����j���^+7FN��"�%	Y�.\���8�e������*ڀ�����r�Ev��s��wl7���� �a�f����
猉�U�9X���ka�Xw��^4����M�`�$g��3�7Q��cYN��x��7�)������/{y^��y�0�kݩQf�og[Cn��[0Ht�c���T@��M=HY�a�ǯ##O>Ƕt����m��=S�D�ꋵ�JST;w%ժZ��rbF�]����s%F����&,�Lڱ'Z���;������t!'A�����ޖ5̗����l�x{2��M95B��7sP·�T�3N=�J��8T�;��YC��vV�\;M˫K��Q���D�^�x��n��v`1>�+��s�Q��d�����u
��gt-Mű	W�Hu����SD�TL�P�A�v�q�t�������<ת���M��Ԯ�Yzʬ�0S�@ft�5�m�o5;QV���];r�=)������+��a�[5�x�Gus��B�ݱ��I8+�bfpG���P�F<�hB7��6�����nZv��͕�`#h�N��O�WA��w��4���Ofwmv���;���4�Na2:�{�`���:��*��ͮj�����q�n���}�F�b�zr1�R�M�)qŬ9�u�W}t�,��Kt�%"���Ŵ���]�2���:e)Amu_q��'�U�E^�6E��O�b��J�WN�f��3`�hZ�I��h^G��Y�&�������n�J���]�����Oisb���3'�Qzn��t�:mj����Z���DW)�|��˯7j�ՠhk�v<�P��ɴ�C4�wht�x>���@��* �F�B�U�t�� �mI��ʞW��X��]�!4��|���A��C�@�ofX�46-r�Z����=�I��q��e_t��k׫)�Br9D�ӠM�e:D9n�o-$f�%�;��Ü�0��bX&�e����44h���5��)�=��Pg��PX^	�[K����wKM�)��phE���ʚ{l���v�\s:�q��t����H��	�:��s���uM�Ƌ�fm�*`�J
�y	b�ޝY�4WR��m7��}�%Ђ���nrb�����o��������ٮрWZ�2Y�a�l��,	]��&'�V�\�����8�8t��:��
_v�U���S��zj���랍i����Q>[1���N���6�*���.�V���z-�K�7j�w2l;LD��m�fw%yM�Z�[�X:�vT�8{w8t��}Kf�]�x:X��aĘ�5`;�Br����J���fU�v�`T������#�+wV��\<���SƉZ��V�nO�J�e��k�r�]W;&9�z�Q��Y�U1_c|��N����cu�1a��çq+v�Q�[&��;:�>"_G*�s���]�r�돵4v����_Xsuu&��QT�����-��4肮%�$�$����е�je ��AEM��B%�٨� F45���>y��y�U{ys��̯9�Xp�܃9�7|��{���eCU��dda���)�eM&F[�[�LQ��FEa��x��x��Ǐ����3�������AI��w0*��L���E�XM�nv�
��AXA��x�����Ǐ<z?�fq�k�g���y���r*,��}���E���-�-�P��1e���Y������Ǐ��~����=��i�dt��,K0˛��`c���1�(�����a��[&ɹ�IX�y��d�Fc��dr�ز�C��l�DQ���]�H�p�@�0���stv�36�7�h�nr��lB#l��j"32 ��v�wq1��*�0!J�J"*�"���u���0��3,>@e%T&�cf	a���J�0"�̌�s
�l,�K3F��
���*���p�9�����3\�2u�̣3,�(�ڲ��L#sˏ
r�y�l�1����fE�s4�5e��t�,64�Uڹ����h!�r�	����#m��M"��r��1�rM�u6b��w�XQ���h9�ۮaXfۘ��[�E{��� ��!������!�s*�'�gm��kp<����I����$��#��ƍ'nf4r���˘F��f��i!���I�\���`�\�c##���sv�?���Ns2Ji7}�B��le}��8CG�f�cdI�I�k����`��c��3On���ۻ���9�-L*���Z}Ԕ��y�v+I�С��	���ǣ�"U�2V�,z��R�]k��,��"��ɮ�X�t�$�p��Q������8r=��߅�m�wU�o���{%�=I�����k�g��9��V0���ޝ���;���l�ל U�^k��-Vv�lӽ�ڞǹ�<:o�9����\FǴ����J���C�2�w��y�j��]zv�7'X���M1�wa���Q�s՝��7`��L��E����{��v���uQݷ�}�i��ޯN���'d_�����t��f��+����8���=�'�ݾ��j߼�4��w�Z��ߧϝ/>��'�ү�����ds�7��������v[}�.u�i�n�ӽ/�C�9Ⱈ1Zb�y��_��z�^Ǭ��0��4tB �>�}�罼E'�AQ(m�6/0����^��S�mw��_vY�`0��vw9�۪�PE����t��>ߘdVsS޿vi���M!���:�ɾ0��>y4��k^�+#�6S���[�\XMJJ���hh�Mc�����̴�@�yL)���i���u��:s0��gvЄVftW&Mv5��K�Mq���y�T}M�=;���VK�ja�4�ť��k�{2�v�y_}Gs[�q�9V��V}o�����\�
+��e��<�U���'��B�7�+t	��7wK���u�sz����L>_H�@����$n��_g9��f��xHO�/{���'�t������_*�E{�^ο!�I�}�޴����ϯݴ�߃�7W3������ʿ=z=CP6=X
�ie�Z�x�j-��}������:����:OS�vϏ�y]��n��-���Q�
�ψ��QZ�у�y��t�/��w�)W�>�������?
�>#����u�_u���0 ���{�v�����?l���"->��w��\��o�Y�8����5�ٯ��Y�w�H��FC�#���@_U�>R>�x.^]���<�.վ�D��o�����hw����z��ji"h�ޣ9��޷�5D�ҟ��>OjNv�[B����K��� "��tcz�R�Wc�Þ��Lv���x���ݥN�$�}��ø��]錭a��6����o�������w@��^=�5>���>����Lm+�]�ŷn�2;�n�aa����ww-bX:Ʀ/�Xb��wB�,�{�_P���8��U����|_^|���:W��L������Z�/�[�E�#l�ޞ ��<�ê"=����;�����:2؈�3N�����<�VE��s:�3��>"�������3]S�a����/�`�c�n�1M��8\<eb��;v1ޟX:z�n8	�9Gs�
 ��t}'{Ӌ�f`��Wuj�����}�;��v�	����=�a��y�F��i����'bC���z���1�r<ݤ������k�]�.�k~b�r�/��Ӟ����q�{�K�[yK�[���,q��q��cA�40k��ƅ�˩/W�Iۺ!�a�gO��&@����oş�G�~�5��+���#:V����w�!�.+�U����Ux���)+^[��H�R]��^o[N��	:�_��z�k<���=+�R��V���zG��^a��n7�*�z�$x�}��E��>�Eֽ�3��Dゅ:�:��Ow&�;9�<�b���WL�=�]k{XwECr�[�Ũ��4r���om��*y���<�Ve��#��=u�Zǁc�!^֦���_W��bl�d;��2OEH�l���z�v���o��7F\��=���A�aN����i^��ڠ3�I�I��ӓ>9l�@�L�>k�������aɩ���UF��h�z�*�*l�����'�C^飇 �vfz��|���y^f? Fn�D��%{���L����bM4 ��zw��K�y])E�)�۝,�kK��Q ���V�Y	������1�{��|v�lOu�y;�r�^��v=^3�j?gw�yl8�,ONQ�gO��v�ߖx�?��>���㛃����DU�4x]�
�����M�x���f숯W���^hdd�fH&e��Gk�q���D��{��1����c�!z�m��������S�~�R�����1ɓ�u�k��N_{5�tf��/2�k�ލ�}��p�ML��38��گ�,�k��7 ^B%4��_�h�RN7hma\D�w7������fu�0_V�7���W}�yu��
)#O��P��A��1��U�S4T�v+N��a�uǈJGCl�ޭ�_��{"h����5��h�-i�ƃ���"��^�7W��o�V���%*�+u�F�D*�F����7�VnIƧ$ �X��C|�UF��k�>潋�����;9_SYۯ�n���o��N�U	�}�'� ����W��پ����ȉ�������zh�<e0�H܆��c��ᕞ=���ΞI9Ι�����8�����cڽb�߾�}F�w�|��P�U:+����*��&��47Xh����o.�"�{$��/�ZD-�y]�o�
ўon�܎�������h�>�����"��y�q� ��ܮ��v�@+�����8|4O{�U=��������<��^���o��=U���j�޻���$��/=Q��%c��m��[8�N4�M6���t�~��Nk�rW�u�
��ww�P �6�=�Vwϫ.��)���^��'�:�K4��hO��y��������v�E\����=O��Û�����T���ÜVo���g�w3��¬��[��*S���n��hc�S��%��ωh�  W��d�=���=[��)V���f���*����u��W{�PA��3���Egګ���eq	gY������P����]�Õ�cg3(J1�u|'b�I��-b�M���P̝6��yJ��k i�^;��������'N��$�Ђ��v|��������j�&Fg���8g|(��ǫ��y��>�e���lna�7����h�y�5��n�qb^#��k����+��z$���»����s��2�Z����oNP�(�����[��Di��K�
n��y���V`�f�[��#�g���
#�ԯ����٢�gY��ݹQs�~Tr���X-�	mo�h��rw�{��;dL���nk��z{�6��_C��14��T�cL�޿{��A��t����W�W��ۉ���G[ٽ�|j����-���H���Yy��n���Sw�j���m�7W9�N�Y�~={C��O�K#�W��YV�w����VX���_�9�E�dXa��Y��GFf�.�u��&�/{+}ڼތw>B���Q��I��:�W�]�O��oz��`��4��p&�*w��mz�ҸG *�^��ac��ïHε�o�"��1���H��%��w���d����(�%d� ���X���U�h��q��>��v����ب�v����΃o��Hc����8.4�������
�N�Z��~�B}��H=!�����;�J�cWFmP�ye����Y55{��{���ڮAvJ�ߪ�ْ{pR��H�t�u�^�n��k�S��I�፾��O������, /޻����^Fg9�^.g˯��(�I�=�&n!����r=�v|�r|=~��?{���{G����վ��ye;�Ro��>�U ߜ~ř��>ˬ�1�W]����T�ԋ��ҧ9��|���o������,�ۙ�rҺ�/&tz�KʴvȎL^n��'4���Ķ\D�~���]=~�!w��8�~ʂ�ʾ}�$Խ�)�Q{~�4[���z��}�k�nv8�׳'���L01S��f�>�0���~����Fλn����^�5Y�_O��q�tOY]�ƿ
�gf>�m��΋�N��i�~��_ ��Y��	��w��]��j�.���euǰ{ޯ�9�d��T�z��}�Mvk��>�I�ja<3o.R���q���cІ�J1-X����4�AA����9a�����og*���ec�;�$��[���.^S�ŝZ�;U����h�J�� �9�c�
S�j�{�m=ʡ�W�EA�'k)���|��ڧ:=���5r��w�p��2߆��b��)�]������ ��n.����cܗ�����f�X���¥f��,�}�z��,E��Wf}�3�ꎉ��R��Ce�1p8�a3�V.'�X��f�7R��c�.�#X��5n�Mwu��:�gs�Ӆ�����)���I�ſ/+�v�\�4vݫ���xK�6��^X��	���<�7�4�;^E_��_׀�ߌY�^i|3a�-���d����w��a�w��g|�*sP�}���C^{�W�f�w�*���.�u�"^�fN�&��>Eu�߽�Z��
=B�Ϫ��6�/g�nUw�t���Ta�+�������c��0��Ƙ�S���"�}|�=�}�3����3���ɛ�U�v{��rm�����D��{�qr�AX���!�oKo�&33����.�g�?o��uz{ؖ��e�M����)^�������Ǻ�{ƕ	s���͜	ˆ�N�&�c�j����X�>Q(R#u*Ȁ�hĊ�d����HLjV�Y�݉� �A�x���bKMwm�lW���3;`�إ�$�8�%�U�P
��TY�D*�,5d���|�z�vm�պ��&{;���n	7 ?l�{����N�z�j)x�}o�wL��<}w����&[~���s�W�*ڛ���[6'}���}�xw���l�24��z�Xȣ�{�����˶��k�+����oW��.���ܜ�n�(>�i����i�~�Q<�,�6
'~��nOw���|>r��bZNzD��Rz`�6u���[��}g�=1�wz/d:����2P��k8V1��Y^xh�K�럻m�vT�<�s��y�����|k��a�a�v���q��5w��q��NP=gϙ��`ͩWU��W�u���B�Ƅ���#a��ྐྵ(�וh��������z���z�cG佔��*p>�<�Y�O��+�o"�0	�q�O]��g�3ٝ]�#�q����1R*����U���{��&����B��놮4˯^����;q8w�,״y����זe&
�ģGwo���Xs;^�N�-�!�2*��61�t�F���V>�q�s��D��^���7�X7�Wn�S�9-�w�VFcn.�[�h,���9q��ٲ�X]gX$��R�����6�pᳰs;�w���>s5 ��{&��|=oޱmk~��É+��]�ta��Vf���B�PqQ�Ou]9��T8}��sʽ�Y(��nnBPs���q^����|G�Tj��г�,�{ru��w7��=WNڭ+�gl1߼�U_g?��q2{ڥys�8���e���z�k=�__"����L��L��ޛ@]g>Po��R��p�7�c�w3�omx����/9�t�5�9ozz<��� tL0Ϯ��z{|$�U��&��s�Y�cӛ;v���~wf�MY��{���#>�w�eo�w;�Wy���l�ί=v�������)��>��\b�ʰ��s��}�������g�����p�B�;��)�G{5�o0���}ps�\憾���]=�G���C�x�=�Y��['{���}{��,�~�{ߢ�� ��{��+�>�	�������D�'O*Cۓ.Mn�H��)#�����ג �E���x:ֽ�r��w3��T�e�D,k}��;BR%�Z�]݊�^������KE椠	�aJm�`��\�v��:{[��B�>|����ۮW��ɷAY@�����A���;
�k�<Ʒ���fszxĶ1ݧPpmfټ,�Ah�c���]
2`����Y[�M��U��<��]q�*G�	\�?����¶A@#�Z�֮i�6I�;t��Z����Θ�k���T+�>��0���\I�s@X�����8�&�3�g�j����%)���,Y��70�<�]���z32��ĵ�hb�=�����''��FM��K���M8s�����\��+�	�ӻ����O�[Pԫ �#��/�"�<ut��Ns�zW��f�s�d'��q�_!i#���t��dڽ�u֦e[��.�(֛�v=�J�.W��	���}�|�'�7i���˫���h�Z�mP|X�<� ��2B��%�1�	Y�up��ܹ.}f��(�/��U]�˳ �Kig ��b����ͥ��K��u������CVF�^��*��/��+hA<�ѽM���K�e������ʠ{K�G;���v˔|JO�8y]�I�kA�x�f�X����縺��;1��p<��0�׎��/�
�"
 P��yoJ�&/�����F��0yWa���P��S<�m�ׇ�X���er�/0������Vd���-������Vp��0y�8�[��NlҬ�1��ƽ�]"g9f��뢢t+��L���]����ͣzx�
�sq�e��ݩP����U]�3V��N���w�}g�h�j�=���F���9Q�iSU2̾/��S1Cl˦j����w�y�����G�owKc���	oӸ�,��f�i]�09�{�<�Q���v`Fo��K��V4�ױ��U�v�l�]�����r�Ҷ��[GrT�'�����⣉��V����v��sK|+Q6oV��t�^�Q�j�a�;��8��U��<��Su��l����i��m��y+V(eF$�I �f�H\���o��:�B&�Boqu��4�ˤ�]�{r��5���G"�@Ԯ�$�y�,)v�4r�+p-�W���p
�Ly������`��<��y'���jh�	�g:��eJ�x"HKL]w��=D�+P}JȽ=�5U����	�%ᴥ�Mn�E�)=��7\<�k#��]ƃ`!áѡ�)��	���hv���4��dk���q���3w݀����4k�`P>�m]��/eZ;�vN@i��~{�3�;�8mￌ���d�fe�	�1�"��|����2"2w0�p̎f5�F���>:�<}}z���Ǐ�����q�^��aQYzi����FeEY9PdPP�g���2l����t�33���sl"h6z���뮳�������Ǐ���3?�{��єT��JJ6��0ܰ)����̲L����/�&�A�1(���p���}g]x�������Ǐ�����8�N�l��MlfefdTR�v̲���'�nP��L����wm�3�f�dQe��*4322+l�+,ɣ'7�LBy/$¢���c��p���i�N�Em�d�f�Y�n� ���ʪɳ7t�.ni��e_c�r,�4��'�f������f6NYd��Ȫ��B���ϸp��A��e�6m��+!�2�0�9.�A���\���NJd�Y����ff�<��U��6yD@FIFYa8A�69e��`�#�o\y$�!�U���e�a�e�TXfFYa>a��f�DPY��;fY�C�VLE94eFK�QY�~��䞪�{T�7vImC�% ֵ.j	'r�N��m���\:��^�{R�C��;�{�l�{��s=�O��!�Sg �	�����1� ]���3���"�GU~_-��:ڕ�'�:��T:!�C���ղ02b����#�_Xe5�ֆz-�e���fPs������g	Se��3t'��	㣝��w��ˍ�$iwY;�\�x|x`'��yL'�8����G������.����`6�f�	�L����k%f׀��4w�=r���S���@�v���\��=m��X�ϑ���[�#.�I�p��?4�dƳ�q]�����{v�����_�bĘ�3���*�L����>c�.T�oP��o����]G�Y��j*c��o;G	�=�4�/� ��^9�L��l�-�
�-m��]�=�fe��~zp�W�}M�ٜE/j��8M'k���Rq}���s[ ����,GE's�]���P)��S��]��>�k� �|���Pd<LOc�/x�/x4멼@c�b�!/��{��5z�`;�q�&�"��*�Z�TZrsUx^��kP㓐�'����V�p��h���o���Y �͞i��=/P���c$	f�_O3��S-�9�x1^1�wT?:�O�]+~�K����zI��� ���<1o3sp��M\��v��%����	xF�/���{<��'Fs��P��uL���:��=۴B���t!��&Y��v6L�ܭm��x�X�=|!cۣ�9��J���Tcl微��k��ыh���{8�[J�תA/pn�6��m�q�-.ص�dX�WkXl��9�>�x\�a�e�����~�7�'/]� ���Ƥ���x��cfo-pv^3���@O��Ny���CP��ff)gH^	Jy��7�� ��c�;��^<�~�����~f�y��A�ݤ�����\熍r�����a��5�u�����}���"ԊoW��a�,γ�����Ms8a����ٽ����@k�`��U7O1���T��k3x�� 
c,����F4��i��}��k{G���'�B�@��I1b�k�54��=׺�*�/`�j�vA�=��<y��9�Ļhk6��͹�o�	r��3EƸ������
�>�f�{nF�y���9�߾֮&w9��e�{�?$	�����O�a�og���8���`��9������94�0�78��n����+!_S���&�=QF�~9Yt��jW�9\�Xc���_O(�^�z���|�f�^U [4����A2��6��Cθ�d\d�d�c�f\ٚܜ�]��˞)xx�G�����47C�N+��x�A�7��j��(J����R�d1R*%�fV������������1ou�y���V�a5б��7���f)>�Y^��Kh]���Nl\:�	P��)Ȯݟ��n�SVe��c�d�	��~
Y��2�u��6a��s�/˽U�%���J��>w�*ϝ�7ΗT�{}Q�v�'Y�:����ğq�-�r��������8�:�w����Gy�P�w:�dA`d�K__�0���>{������}?)��Uo�<�8��<bUx_>��ƇdH	���9�.z[ R}Ò+4����gн��ʜ�AonQ���ðW�����/7+�n�Ӌb̲�bӹ=\�Xx�^Q��"��6�\����L`�ت�۪�N|o?��^֍vm��o�F3���l`6�<�~��X@�һn9O�����'_���X��IW��<q�Г7�9���vlk�����i�px�Jum��]EK4������ȳ���L�F䷄�5%��x�J`�����R��*���
��]�(�A`��B��՘����
z�rp;�������y�	��s�y�2*� ��ڮ`Q��.Ng�H��� k_�뻷��
���c���xLv�\�t7��T�c��as�s{wf�|Ʉq�(� �����-(��X�ί<�V�ь�8�ޜ3l-�͢f��3�[��}��+��������>d����C�7R���EEZ��h�.\�I�wz�������߹�[�(?y�Y�?��A��sK�nw����>��p4Ϸ�����yS(6)M�`��%T���A��̤Yx{ƶ�� ���,�S�!y�TnNñx|2"gd/���2��"��J���m���	�]>4���`^�y汝�b�.�Yb�hl�wQ/8Az������d���� �[,�S�o��HK�)p�r�T�u� �k�W�KT�q��l�&��g9��]c 8�m���t�	wڛ%s���c>ͣ����w�W��a�e7���ߟ�g��~6�l���|ڜ�[2ɒ�[��wT,��G����xa>e8_��wf8y�yƓ7���� jb��vo&죬�����n�Z�[~>�J�`�8Ͱ��ݽ��wa2� (��s����E�S�,=�G�z����_�E܇m�L��a���S���r����s�&��d�@l;����ͳ�|j`�'�j��n�)UM�Cy�4H�5��i$h�Uǋ�s���I�kӑ�{�ٗ�X�oؒ5_��	�ɱUa�����F#M���f�x�
i���Y��k)۟��}<�x{)�_�Usq��-�Y��B�����R�I���8�p���j���w�7Areg)}-��|���:�٥�i�-X��yb9�*��e ��P*3&</�F�j[�u�d˜��\�����TU�p��fC���f�-���5?D�L,��w`J���0r�����=�Gd����Xl�&6|�]�vM���@���23�?]�����w�2}9�ʗ_��p&���y(�}^JO�Al����&#�x1E������P�+��Z����9h.s��6҂��|��Urz�]`čocl����޹��nH}�~y�����/��}�ʒ6<�V2��m��ϵM� |�}�ص�k0m��"�	j+[���fۖ�
<Ȕ�l���f�?��}��ٝ�-�̮�nmtp���:����v1����������ߟ?�?��`㓃��٭�˛X�C�^<5���Dt�u��j^9�������hb�	iLQk΀�D�{;4�WCl�-{��P����P`E�S���e��CC��>� qp
G�C*��cAΟ8n���X��y�Ywvn���y�sN�#�� ��kQ���̃��������3�����皁Sͅ�\�g���^}�/o]t����p��ߣK��M����#���@�g<%q�� 1�ˇ��n��gG!�//%���{�����7U�R63���[�w��i3�m�]e�O�׸�\�jo3;��˟<��)���gLF�n#�����,Pi��;@��c&�� �vl�C2Ǡ�(u�0-��C��bJ�.2y���n�1(����%�Ǘr��;my��z�J�y�^ێ���h����0�'A�]���)�TF��_��d���ӳe�=nh���R�����?��*�-�𰕢�
j=RE/8ڃ>8#m�l�M)υF�c�����(����'�q^�x >z�<�H�,#�B�3�����9vYy�g�ݠk�K: �K�:���q�M�d�-���T�q��s��2���H̲^y��l�kH=�2��@K*p��P��PybZ�SL^wp�kT�}S���^�GN�ޢ�:/
���h0L��hV;�^����ӺWN�8�9D��	[�HGt�K�p�.�o%u6�hsGlb�e�"���ۃ��Y� S�of
o��R�Π'ߩ����)#������;�}y�y�?�������x8�+��׾u/����M�
�ǻJu����F����u���n�&�:'�����
���a�i���4z�c�
;�o�%R��	��W��X�X���Dc��q�v0C~˻.v�T繢�v��*��6�l3���b���l���щN���_�����A����"n�p�~�L��ۂ�2�Ð���vC�U�aasЗ!��[�&��i�C�0��F�if^FFvs��|^g���s/N��J�ð�{�|�Z�l�B\E����܉�=���0�aF1f�~�!�1/�צ�wf�aE����%���>�/����@u�aF���ޑ�iPk��m�_������"���B�u�=Y����m�?>�0�8�S������q��vuЀ�O�<ۖ^��+�ȍ2'۰S�d�%��zC��}&1�ީf���kNS,X{S�`�C�\3�wi�D�y����21P�z[���-�-�ƶ�S�&�X�+�!����-� �w�Ce-B�{�T4���p����?[�[vZ�F�mL��꘸���I�����fi�P���JF���W�ޒTIvخe�"p��͟k畏WQ�z��i�W|�<+{f�)xR"�������������7g)�%pKQ�OWW]lyy.�-jn'r��S[��D��Yh�K@�jg@��:U]kN�H��A!����W����J�/7�
�hf`��N��.�}d`o���y�>Y���=�^@׆�*�炝&�q{�:�ۑZX�EV�!�� ��&L	�p��fמ";�ڄ+��	�wU���H��.���N����u<N��9�r9�4��T����WӞm~��v��N�â�6oת.=�۸���k�ǲ�%����Y�����s�\\r�3.z_i饁u
�F9��&4�Ь����5�/��f�8�"���e�n�Y�wmL�� 3���?D�P'���v�����Ly�碓�{׆�����@.n�ƫֻs'�c*�` lAa�&���]��{m�2����|f�J�d���&�kznI��d�z�l�e�����qb��v�
Փ�瞒��b��_n��|��1ר+0�k1��_Lf_RU������A�^�˟�%>٤r��g2`
�O!��=�	�=�{��;��C�o2��l�T��.�{͌7�,�T��|h���	����JO~]~�m��s��l/A�������d�5�,݃}�}���OCK��><_��mV��uE��<s�����C�Z������ɧG�poT��ރ�z�Ż�{�;y���-wT1�JGW�X����X�nڼKv���/��L"��:�9��`m)[hL���Vg:�Υ˯{��kgr��Et1��9\�VkKN7�簧]a���\�:*n�Jݪ�a�d<���=���n����������]	��fw�F;q�U��w�\O��z���l��������ܬ��0Z��D�]���&�Ɨ�}O��+��R.����y��FkT~��Y��3���6�Ɔ�z��q�;������8�xЀa"�_U�2i����Gܧ6g�M�N,��g�q�.Z��q�gמ����~����H�(��<r�d������^��im^�1ASG��i-�k�O���F�]�r�ƧL7�5��?�7�=/�<�`�K7]�����ճ�>Iw���X�v�4�^Sy?�� �D�DSc��Bz��ȼ�y�AçE[��7����~�k�%��n8������X��Fm��Ky�B�wW�m:�B��z���p]���8����#\�u_�9a5�$��lٽ��*������{��Ս�똇�zw��{ki�m���Z�{�qѓ��<�
m�$&�=[8�v>��CM��k[�^+2��ݧ��f\��7e�����_�~uZ��p-4�s� e��&���L�b�{���Њ۠@<efl�3�2�ɽ�-Ώ�]:��� P}��UΣ(���B\b6f:�r�Eo57:X8�����7&uۼj:Nmo.�wW}ٳ��cK�q��{��x]�>s�3��D��$0d<�;x3{��{հ���D�Z���'L�e�⪙����l,�`S�L�����4��t7q��/�
����m�I�h�ٯ6��7?=��œ<�������A������JR�$n�>�xT��Y��$A��.4���J�����6���d��c�lM2��5�򍙾�h�-�C_8�MQ1�>y�m|e>�:���nr��%W'N�رV�O;���I�����,�� EH�&�}��ei����0φ~�3^���$�z�L�ځ~���R��K�r�Nm���L��td�}br�V�O�P�>|�5�.���E�w�e��#,hǘ���3e�f�h��C�Z�ղ��m�ki�>f�c�v<�f c@}��]V�_�dsۣ�y�4ˠ^�ȍ6TAO}��*�w:9O�����Q g��,��t�:�i���@C��vE���|lc���6��ơ�F,q� ˁ5��s�)�;�׆�Z�N�L�;����5�p�"�5z\Y`T��f�;�=�����mU{���d/�׸ �t��pb/�8�n��j�����0��RP��@�q�H<��»%s�=�o�i�z���:,.o��)���@P&���UD
��� 
�7��:��Q�f��d.7-�[��q�=u�IN�C��c�LBC]3W3:�8��vTۏ�߀�a��hZ���~_x�Y��K��-�1��>�;�\�/-BG�Bi��nW��a�#2�vn�v�D�3�t:���.�l7!�Y�im�<�����������U>5Lڨ���2�_7ݟ���F�'�J�霳�L�Y� gw�G��o�z��/�Y�>��M6߻��+ߌIx2g��Z������:�ܿb�配J��i��C�Ҩ�4��]���74�p�eimSm�)�ػU8�<�D�{���	�X\����;�\��ˊ\l����ռ��$��ͧ:���M�y�¥Z�����Ş����z�cAM���κ�����Jq��Κ��>�I�+��oب^	���ev�w^ŕXgG�L9�\]L%�����ϥ�2~��l}A�7ق`U�N�(ƥtD�����a����[d���F7W\�Cg��	U���V>��/���=A��6w2ԃ`�=�B;b.�#��6{dVm�	L-sb��yvŊ�����[��8�x��]_��K:��M�Crd�$�g�haƸB%�8�K��g��&��{��x��!���>~���\�u�zgȄ5Q_�.��Y���L�q�dާLʇ�צ���H��u�<+��<��پ0n{�/����7�5qLu�x{����5:N���S�]ՠӴ�7`WA��ڴö�wcA-�Xs��ŵR�4+E`z�IuZ���@S���[�P�x��'�]�(W'��)��Rk'K�P����n��\-ԃ:)u�nl �
�� (&�.���f�U���ǌ����7��1_Z��}4M��](���������kyٜ&e�z'%�ȼIZ�#7i����+R�3*��Z�CZ�y���\+ Y]�*[��9��T���m��bh9YB��+uS*��n��-w.�,I�7����ǉ�!V�*Xg3�N���3�@$��I��.1jä�E��'>1B�XV��ܶm�B�r3�����{��]���v����V�Dr��|l%���}\�bY�a9XE.䶖_׸�d���o_i5%s�z�Z�j���gr�7"���r�SWmv�]�ղ�Jx�(ˬ���(+.Q�˒�����}�Xٔ��Z�s�Ĉ�۝э)Q/�L9]:3������7w� w:�1]
XG0�&�uJƻ
=Y���qZŲp��G]^��:�s&�'C���I��c�B^�۩�;�]gZ�k����p��`h�Y�**YYM�xh���y����H����0�*�`��X�+�ӛ2�o(��q�eu��6}�o�L��2,VRL�2^d����2��d�޻ʼ�M"��������I��|&��WX�%) J�<�����U|��D'!��5n"����C��}���Ju��}Or����QN�h��U��_G��:~k�郾���]�2�#��B�%��6R뻗���+~��<��۬S0��D5җGȆ��o���Z�wn�6d���Y�9�M�k��
�"ʝ��Xo�텝r��O��}d��=�>�W�-:�_\s����jd���M<���c�88G!�V� �VoaU�|��P����
.�wi$�_�9z�J[��1i����L��X*	 ��1e�t"�Q�>�6�Y�`9��feQ��6�1	Q���n�%^�r8�&�j�G:/\h]>�c��vO
��Ms�k���\��!=���+qt���jGW���5m*7��u
Cg+�r]��	g�S�g`H��֜\��^��u+z;����*�H5Q�&j09I�8��ѵ6���6�i$:�y�.�$���ꈓ	h̭W�f���+�kC��%�`S��6�Ȕ�e��X�M���g�ra9��9Fś�ؕ����f����e)�c�U�(�r�k�����Wݡ2��9���*'��.c4�$�>c%:���J�"��5H�������˺xEe�۹�reM�Q4�K�)�;�:��B�M[�K�U�oLu�+��j���.\�K<��bt�P���m�����J��j�� >TC�t�
BS%����*t��$4c)���tҲ@��(�@`�-T�Ձ��BP�J�HҦC�ڧZJ��7sp��w�Ku���n���+&3&��UN�[��m�w�3#3���v���"�$�_�:��������Ǐ�ׯ�����Cڃs4��l����0�)2j�(�3(�3N�4��e~}q׎>��������������8��~+��(�I������622,1���nQ;�AFC��8m���^<x������������_�3������I(��l�l�ir���22k#$˱�U���r����p����>a�F��S�aG0�K;��V�Xfr=�̾)���f�Q�XY�EI�n`��f��i�j��lǛ�ifs2�d2"�͍����E�D�NT^n���ae�A�g�i���r�<�)-��r"�6i�aA�Q�|�6,��G"��� �2,³3%�<�;�2��
���(�!�,�bnfY5��&X�ld�DY��FMf�Yfd�U���FfTBXbewp����{��2L��p���q���$�yn�e�?=�����_=�np�OUn.���x=W����U���u�>��=�0�Ǘ��T��KK1�������OT�v3 ��^Ս.o�O�����ʸ0-!J4%�O}����y���>}�s79�L�2�~��_�����J�π�d���?����g�E�kpf���ۙ~6��:k�0�����LPǤ� i�#W0��0��m�e��i�֨h��0��)n_�7ֶ�����"�V�X�����9�y�`D:de\ySM���h_<����T�i���iVf����\Ð�5�(g�8�}�*���i}����{�������[u������k�2hܮő+X��9�ёa��L]�?s˾���֏d1��
��U����9bV
Sצ-~RV4���^<��m�z6�"-��5�8�Ǜ�;F>�Y�f.�<I���E�Vn&��;o~U�cV\7��@{1����m�CN-�(�E�2���6O=]�Ĳm�W�ف*"�`7�aKȧ��	D�������r�y���1�"{��r�5�{7�}צ�)?m�:���>k���M;Ϯk:im�Lu��b��ʌ���&w��*Qp�%���qy�Ui�E;�C���c�[�U�����J�`
���j�K@�3�x�>9O����ׅ�W�V5i���<參Y�qx�RsP�ym�rNaG���ܷ��LKS3.�sm��;�{��|Uu1�9�$d�\Z�Z�V5����)C	�`*n�8�;�b'Y0�F���L�6<�u4W@��3��:2��{�y� 0dH`�#�ҿ�������U������3�M�V/�fP��'%�[����X�S�P럪2A�n.{m�R�9Sܚ�A��v�����2���:�eL�LW8�yw��/>N�͍8�.�����8{��t����{�)����_���e-֡c��Nӭ-QQ\�-6�4�Wa+d��0�BT<c���y/"ё6c��4��p(�ds�g����Q�M0���N�ŬXצoM;�!�;�|10�<k>尥D�]W������j����tG��/���ԛ9�}]��kc���0A`��'�ͥ�h�����w01~��O^��Ɍ�a��Nb*�����$?�~Yߐ4�.�����(RT�}����5O��֒b���.����k7���L'�Z��Y'ۛ�Q�Ge�V�Þa^u\Vt&��3���T�ؗn>�d3t��v׀��o>���䮾kT��vx��D�l�R����w��}��g�k/��C�w�+�U������'A�G��R�b��ƫ2�wa������H'�s��q�f�ߎ��o��[��M�n1M	��<bۣq�͎�p�v�ѻQ:u�1C�S��#Pw�{��ZX�S�L7�<��3����t��e�e_�k��,��b�\�����O�9L�ovnH^���k���cy�5sR��R���W3)w�N�8�Mg��<���X��o&���'{�k���L���!�2B���S�o�[y	��w��k�o	�I@�{7���Z�Ic|�B�	���r�2Gd�U�@ځ� ���OJ#42���~;L�O��je�lT�t��ӽ�-�������{+vw^%	m�����j�UJu�/ҩ�VbŅ�� [T8��0:��͝�v������w��"n2�S �1y��Vyz���]Т�(� ~�ɻ,�,�0�L[���A���ь���$��c?~����eM^�j�nYa*���E�l��V0�*r2�F)��j�qc$����4
�����?��4��nx.�h��W��wh���n���u]卞��֛���T!L[���N˰���Ih�	���<�R���<^�E'>����|��C��	�X���J����g������Ý���QdR�oM�'�&�\�zvW�=������¶�^%{Z��-�P/��#`n��:eb��ҝ����~t����}����I?gL9�KYx%?Eܶ0B�hL�׺UmG��k_�����R[䧋�~͓]f(:�1M�@䭻�`��St�a�=ǱI�i]^պ`�B�E�?;��\��F���(ne��BO����ަ��XY�k�D%�f�X�+��<�+�����p���d=Sm���(��ϟ|��w���}���0IO�a�!�D�P�h���������yg����)Hդ�Ñ��/��z���H�C����k��G��yn��m����kYՒ¢[i�]���`���D�Y��[�=�W�U�fX�u/s����ێ�`���<6�v*�j�J�W�ꡉ0���=^���K`ny�<)��vg��=LD�9��{����q�t�0ga�D�W��1ʈK��B�{�������������m�m�SΩƭ��lj�%~�_��9�׌|��Yd�tJ�a_<4�T&x{nVޏsm� ���g13^�]�z��슎��0��U��F����@�Ψ�s�R�U�k�UN/���㍚��е���x�,)�O���z7:&%����a#�\DO������Ɨ*|-U�6�پ}�����=�u�K?�<O"��6�/!-G"Y6����dW���nP�ӳ�qh�z��Uf�<D����,[��5�݌P�����)�=��(�P%�J�ǵ�����BU�X;V�熨wc�Ǐ��ͷ{^1C���E�0���(tJ���Bn,ћ�$Q����صm͛n��U��-P��z�	���v!�3P�'��Rs[,k'|_D�r���Luk.� ���J�]���N���('{ܥ�]�R��[֝tI=7T����kV�o�B���Ҹv�{[�$њ�5�O�㥨)�{'WN�VG�uB8�'���P�.nyᇾs��o��
C	�0aLI(J
w�^�k�װ���S��wB/�*��j����oG�Y�*}.�������
ĪZ�V8n��댶����!�p]�_�x�Ү<q�ͷ�5B@�}M��\��7�'���E��vOn�>��b�G�q����s�/H��ƶ$n�����0J?��FW�6����kR��~�g��)��Z������%�-0Yr1?+�IώqD���	�C�泭e�����A_�E��e�=�p�U{�Ro�²_==Y��0�K�-���k�[��+��z�k�uH��dЛF3p��5����ҟ�i�7�)8�="�}Gf��F�@�]�*�܊��O73�ζ���-��f�������ؠ8eO�.<�ƀ�X������͉�#��7m������:#Xm~��J��x���w��tu:A�>[��vj�3Ż�����}�\��ly�`��yz�e��\�Xi�W%��hN|^]�u�k6R�2XX֛8`k��TE�)j�� ��MD5xc�~�^��k��o1��6�qt��uC:|��~V���`���?�F��AN�';XB�'t<c�Z7l�h��������vM��e/����6����7s,�*����Q�^ZwR�ƒ1�%H��#E���@�I�b]�0�a�B*P���K��*�u8�,�63y��t�]ft�}�^N��vMⷻ_ʯ���A��dW B� ��B�i@�?�����=��~������o�Ox�ڮ�}7���(zF�?\�Z���pt��3�f+�jil�ĸ�[9
B�.�A�"Id�οh�y2��0�h%t+�k|�"EN��9bj�Cdd�>*�h��g�Н��T�� �����lu�����uf�:�b�u��}������ANТ)�"7�V>U�X#���U?<4h~��Լ*	i�&Ok=��S�@����gț�^=Y�+�NKվ;�i��>d����L�߻����$F��O�!
�J4_@�O�)=�e�ؔ�g�bL�zZ�@�vkmW1a����*u�yW�\p�
H�x>?��P��^$���!�S��\��mAt�my)Z�/˂^Rd�~�K0�>�71�K�x|>�vw����>��<הV*�"�8��6��YFK#�g�F)��4#�o�W�O�`��#X*��~X:SKM8����H�E�B�ڤ.,�:{z]7�������G=g}�)N�u��
�e��.�ةK����Qx������<���J�6��<>���@4���<�>GiB�����R���)
�tȂ�E]i��C�%��0uۣv�ju{r�!J[���վ��[���Z�9�����a4����	�b��&ǘ^�>v6�)B4wE�Or��J�7����J�V�U��VB��$2���o}���+�3�Я�r�W��j�hk��_�m�x���0�����tݒ��\�����|4`�R��r��?l�;��w�GkѺ~��#�r����*����O��U6\��F'�[�.�兆�Y��ƐK��Ͷ�az`[1YL(���0K��GO������屻H,�ͮ�[p�SMȈ����W��3c�}�f}͒��t��@#Sl;�+��p��{��,軕Fd�s{@õ��'wQ�Z�0�rT
��Yȼq�.�;G� ����m���z��n��� ��K��p��3�ɣ�z����h�5�9�~fl�Or�S�S�L2zozb���`gJ�a�*h\�k�7E�_<9sKy�n�H����ZUZ6��:/����1@��L�38ۑ�m�B���Q=V_�y�Scܨ�Z��/0�S�b�-�xy��2�{��;�[62Z�3���;X�{^P@����tBd/T���QLPK&
v���`�U�ER����ߦ~����'�uD�tr	mH��@-�������_y�<�נ��0�_�U<�9�^�L����{s���~g��t����w*���c3c��$�Zg8�md<)z&+3,�@\���4U[U�N�k��h%*�Ud�"i�J��׸���R�!�k�U���O^��"�Ǖ�$� !I����=���{Zt�k��>_7���/y��>|?�z$��(�	"9
	JJ"ߎ�j�J�6��gy�5���{e�H��j����O�ȽT��1���"��D��k�aѲ���]K��Ok��0��]^h�LB}h�mzgc�)W7�܌��zb���[,UhΛ�l���������)�ǁ��=6�{�;��C?��g�.�H9O���*b�O����iWj������r�
0��9G7-���R1��3v��@~�G���0V��$k:�)ս]P�^�2�V�^���l�-\��	�Z*���[!����nl��ϝχ��SS�pC"݇2�s昽z��ߟ�T������x%ݿ+ߏM��oM����'���.�{���Z��Bmu�vǇ�,&o@� ����dU�ß���3�Ĕ�kdnC�M!�Kbi���4復.���Q�v��ɖx���.QX��s'�����\��U���ݫZ)
mCP�c�(��b��p *����������c�k��MA�gEGk�W�%D�fA,���f��a����
X��˧�vf�
Du
w�ն�����������/�jYaB��t:2��[�Yj�6Y'9u F�P��@�h��}M�E;�Uj%�F�ܧb?^.þ����@KBkX�
oz��vE#�ι�z���W���3x���lA���k'<��W�=N���-p��/��8�SfM3���t�r3yo9��g7�0��2A�a�`�$A��8��U��.�?��ٷԼ�T^y��@�/q�;���������
 �%i'�M��K�`:`���UJ�����:w��ԄL�יq\�[�:X��&Ė�\_{�5���[����b��l����a��SW4����0E-��n�uo�К��0*�O�1*۝�֪{b�
z��{\���l�%��;/^C��q�)��
�`'�� ���8��*���G��Q�Bժ獥M��H���a����:�p3��>�1�uVs5�h�WKtF���ՓY�����X=3i��)�����z����	�������8F�w���y����6���;�&��`�%�i��T`�.'��ҎP�pڽ!�������W?mOo5�������錞Q��>-��4��s���\���R��ϧD����]I��g��k�o�_qs���;�iSSC �	���/:���@�2*�O0�ڞ����&9�Ϭ��f�v4�au[I���;s���`�4����T��b�='��"F��,���
���4��WV�{(v���R!si�WCUևÆ��؊���JlA�5����%�{�&�?�z�W�[�t��ގ�L>��� ���wԹۡA��͔�t�z�m�1<׃�V��%���,ij�(S��˒NF�]=����G�:�{���������)�*�0�(��<�{��5koZ)���V���t�76�ݛ 3�wi|3�0g�:�<��T|��u<:�]��h7�ٸ��-��ߗ
�K�x�>�� o��Qô* ��<L��Lw�3ẛ
�Iʩ��m$�y��v*l`�z�2,4�WI��[B~���2hJ�>+Ε���?q����۸��ܥ��L_��o�|�����5�yO�&L���A`����]�LۺoW?�T,e&5H�SL���,.�1yB��Kո�����g�d0�B�H�����ނ�|��货gxZ�p�*`���[X�'%��$�]:����݇�F��aӮ]�y�)p��?�����L~��(���t�`���<���
y�eH���ޛ�9�z���T��xF$d.l�AoMόR6J�..��vݪa��N"���V'�~��~*{��4�}����>L�����&<�犟#��@�w?n��֭�,�g㔭ePg�<�A��\�^�[1J�t���3X���ߓ��S ��%>٤r���ڋ�O��O���<feh�K^��n��~�����^�˖�63rj!S�œ��V��TB�H���*ұ�A�*�5u�jЁ cxZ6�)��wr��5�T�-S���-���,�\k�mIW4��v2�>�$n��1�ڝ�������)+A��*ҭ�Keނ![�J^��	b�u�}�$i�J�ת�����}�1���.`X���F��DN�l�/�I��_V���Μk���$єO�7�r�#�J���Ĵ���U���Q�s��8���yh4���`�Y��.�U�� *���j��r���|�y�t�V��H���d���*��l y���b�����#w˝n��A뮼��{&�ʤ�k�[كY+9̣�����%�eڶ��?�-�����o=���Y�M�k�We�!�rƯs�|��$�u����J��y����aEe�{nd�HZ�ջ3���"Ce�ʫ	����z��v�jM�G�T�N���TFNf�۴�E�gvA�$M��aYk\��U�.�`�z�z���mes�u
J[����x�M^v�k1YЙ�
�_T��w���G85eЏxA�!�Jj��VYt|f��q��,fm��;i�=8"���֫s$R�"�聺ڂW]XMA+�H7���(���N�X��R���iN���Aj�1��L9��*�bZ��o)��Dx%<�lu5a�{zn��(�kt��8��R�V�}pC���t��ʾϲ wyCN��*!U�N\��W|7ݨ]�`�����f�\���~S{�*G�e�<,�;�����������Mzv#D#��x�M�/k�e4�d:��>�X�u4E�
V�bpг+�$�7*F�],�8�7�mf%[�M<M_r��9���]BP���j�X6��:d�Hᔒyv�]��"&��:^Ɍ�Om�%�ܮ	F��'N��>�L��]���\O���ɜ��G��(,@7R�C%�'�o�����$K�#4���3�U*�c��]Odօ����v�v*�ӡ8n��Zo����F�wN�]�m���[�6Gcη)b6��3����y��6eɁ�<���`��X����ʭM���R���γN씵"x:����{�y�W!�o�ncY����r�Jx��<4[�`S�Cori<�x[R�o�:�ぼ�	�)M�n�H*�ӽ�Q��6Uh�Kv�u�$��,�[�Į�ݵp�%-$�d䶮��X���S�2o��n�4l͸˶�ʚ�mZ���kb�i���c�]t�����Ԡ�Ҥ�!H�j�[e�]�F�M]ZUkQQ�9�����ʂ���6�<<��EY�t��۝��@ɕk��N�Y3�M�;�������7���C�4�<畖�=����2j�l�f�0p�&���\*j72���V�֘ѐg��q׏���~>���>=���8����,��,�ɳ"0����ʖ���lv��(��s2�2�Nm��^:������������?���q����3�N5d��m������13
�̒����x���__Ϗ���������q��{��#gi���&�����7p�*�0�&#0�,�' �eQE�f�fcNdPV�m���&ɅKY�$�SFF�l�S�f�}��bY�P�d�-�1�3tط2���afdETQa�4�>����nf��[�i�Tu#+s���X�·0���3�ط2
i�ƪ���2r�>fk�Q��Q�"����+�<�*����̳���D�c��fdUG���aDRy9�q��cp�b�1��$*���##3wJ���1�3p�h�#l�Ȫ�2Ȣ���2�\��0+qp���s{���(X��=ùA����J�u�G�G����;�_)�k�ӎ����/�n���M*�ʓyu#�f�[_����W��Q{�P�!���}��n�n7�OM}A��ż���r�g�=i��q��Sq{1R�Ϸ����\݅Nc�Zֻe�s��e�Y�T��A�נ�LG����m�yO w� C3Eʎ.;�қ�8��y�Q����\���i�Ŭ�V?	�~@�U��xPz��4�%������db4*�I.islI��ճ�V;槷K������1�,�����q�<w�)��@#ˬ���2�c�o���c�+^���-�e��=�1MF=Y���Mi�1l��ޝ�����x��L%��s3�Zzs+�iu��(i�f���8��ܳ�;���������G~gg/���{���s�Z��f�:�A��S�1�����pG���V2U|f�f�UE��)����*�l�:F`���|��d�?i_4�~Y�Mڟ{�m��K�y��8\�:_t'�Oe��?u��ޫ��낎�B����,3�,�ly{�a>�E@����~����a�P���,a�)���͸Yro�5�q�9�uN��Cu��]�ɢ���V�F{
c��S=�;��o�����1�Fnb�]�O:�|Ai�VUM�#~u��H��ԯ2�������Z��Lc�n���v��u�Q�{G��p�-��C!�L��l���p�[����l��'�E4�N��f�Lǝ)�G S�jet���M�����6�s�T��\Qpe %R�w����~����n!k�h�o	�¹��0�G�^�?cH�M�Dذ��v"4��b���ͳ�М��z�;������jqK'�1,�ہ+���+2���=32���v�q��z`Z��AgOk白�X���{�lj���XO��S-�
�d|O-z�V0)��M�>�/.�z�����\�/;��E�\��O�C\��ݑќ�̩����.�P�S�݉U��b�L�1��?)�M�"���
i��h�%.� ��ڸ	��ꅮ�n��-�����0�iji��_��Ws�!��7]f:hhwv�����D/r��W�d�ߗ�D4��(R�o4u�5�>5v��j�U�W�G�.Q˯�$n=�ۚ��F���]��`�Aa�-���J�MO�*���E��I)�[��@�q!�E������p�͞��*D�tT��ٺ��[#���8���]���[�K�C{Zz1M6�k�0,)7k�rB�y��iG6�#��cm����S���#T��m.�d�O�)������Q���c_�#������B�d>GH��H�Y9�}��R�{��y5q���	^
��10���u-�#��X<j)v_yV<���l'���9�t��m��6����tA�*7wB���W;�7��ٷRQ}�gk��(H+���?�~WC�[2�LA�Z=��;�:�r�$:�[���/�۬Wy���I���B�h&X"s�?�P�F@H`�QG�U�RJ)U(Dw�}�~��~{O��v�O��QdW'D����xS�L
���>1�q��5���2�����K���g�e>�(�W5y�,3��?���z�����s�L�����9��.ȯ	�fÐ�`�+�'Gr��ݶ�lsdN��u�(8���(��1������C��������W��{�X��3+�������Z��	���Q�f^[�e�0#���
���Ժ|�ڙ��.�n%�3]7�OF�9����U�o��Ȧ��׭;��T��蘜z�,�e
�vp	"�Rφ,��#	��2����׸�`L7����%J��A�x�Z ����	u
� �~S"ܽt|��Y<n+�4uH����A��N�gf���&���ݏ g�G2eη"�z4t�ޤ\�l��E��浪s�`�H�ذ�l��zkg*�߃@���8�B�AYf�@r/��s����k��V�i���¬f�[dj:���Vz�B2~��fUMЪ�zKfyis�2�2K'Z��&,�R}�J���g(m�MІ��8cCa;���[�&�A����ۊ�s~'-��=s2�!5`2��S�uu+�����PK6�����y<��(|
  I��x�d=z�^-��rZ,j�9.	�b.�[pԏP9���r�<�o�x�Ż�6Ũ�@�	�"��,2*׽� ���۫ݦ��A�aN���ɫL;W(���R���(�3��kf�.�!ƻ�����|4*��bs,NvWy�B��χ�V:|]_�L:��������X,�x��-�%ɦ�p1��ռ^D�d�R��v~2���C>K	��/*�O4y���:П�0��ǀ��Nf�2�����C7���t;c�w�h�귕g���tW�W�|*7�]�Mt�hi�y乕j~�1���gɋw�Y��4�C��"9����M�z���[(�Ⱦ=]ɉ�t ��
L�r8Vm/9�P��t��Ҿ��Q����_��w�=-�m�`�=��ڬ��A�p�<�Z��2l�}>��8�}��/ �AV}L�ޚ�C�.Y�$�令�Q3����&�XLL[.�F8=;6S�?���If׿?8�Ee��m�jw,��c��Y��K�f��y良���I��S]��rj���� ƸȖ��ƹ�`fR�����[j�|�%���G���~w��K����)���+z�C(�}�U�Ŧcz���E��p������_j�R��@�a&K��v���q�̝x�m���0z{g"��:�Kwڮ��+�s��z��0�t-ʜ����洵�Ǘ|`���t^r��ůu�=mL��]ƕ�0�]��A5us~z\�}���ޟy��+���H`�� `Ȋd��ϝ������!������˭�3��Z����玑U������z����&���۫��|�M�J�^�P�����Z��do#9�-W��L�����Ғ�g���o­{�kc�\Rm��~��K�f���������;'p��L���w�Y�+�Lcз�q->{�iS_@�F�X[7�ݹs/C�J�A Y��-I��~O�b�s�P��M��.��}��Q����Zo2!��}�o�������C�����|�!�=c��`=��S
�uIn/���7.�l����1E�ll�����٫3}*5��*+��Z��ķW���v�~���Ű3�fx��Y�\�\�����N0��W�bu)��1m�^/��!�3��s�&"
~���ƅY'e���/��m�����)r�7���*'��b6����4C?7� �E�*���T-�5��C��]�,ꩂƜ^�Vޑx�X�;n*�
y&�����r�6��9��fC�
�C����{8:�y��5J�!R���u9a���l�2����uĎ�z ��}s/�L�{��gH ��x��|^��"�y�6*�mU���^���i������].Ϊ��C��{\��=8�t�t`I;�W��#����;����nk��Zhf��u+'��e����f/�]>س�Ռ
I�]i��OM�y-�����.����0 C"���
�!HH{����m�vg�G�+$>:/��'1�FH�{v��s�l�6���Ew@�i�*��	�1�+j�Ms\����Y��%�!��ߞx����k�J���][+u��R9=]�ʆhp�P���TK�k:2���V�RG��*��b��8r��s�!��ˋ�ɛu����\:	G��#T۸yF��N�;a�aہ�5��=K���4�Ow)��z=����%>����|mt+V47�}��!�WE��H��v�"��f����Ȕ�Kxv�j�Ӷj�jA@�=M������)�^)b�f%P�k��1��
̱v�i����ڜ)�5��8����v��=5�Ò�\�kd�Aa#�e2�U2/}���m����ۯ��`����Bk[x���O��n��F;�%�\��<��C�]#S�y��酂�Sw0����f�9s��jK�W�M��P��<~��XfEϷ���q��w�v������:c��CMwZA��ԑ�M��Ÿ�DQ^�d��[H�+�Z�l���2���P�tN#h�G���u�w�շp�T���[��Y�V6�[0��VQfjQH-b���9�<��a�U��H��d�Y��7��f\�w8v��ώy���'�RhHM#@+x���d�H06	2���Vת��*��p�u��M���-�JorA��eoGΡ�O�	1�^���Wn�{����tS��T���pܳ���-����d82� 	J+�/>��zz}��<�y�3����ހ\�7�"?9*���9�مC��b��E��@��Gy�8[/�}-˻'쫗C����B�YY�k�g���Q@ܶ8�Z#(tl�x�6��f�=	�\�q>l��Tbz���檦X��g8&~_�Nǡ~���W��χ�TV%Odi�=��5�X5�����ga�ѱ�z̦xg��3�kU`x��A]�.&��Hf�QQOs��s�=��� ��/D[X���͓��,|�/�`T�^���1Z�7`[cv�4d�WcW�Ms�m��F:��z�]� �34���3��H��T'�ʈ?�>	��ߖ 1��/~��.�%S�U�N����{cs�� &���X�o&�ެN,1�X����`k��*=#ɸBs�z�j���J-�Ү�=�
}�p��M��Q����Y���Ƙ�D�j�=�;��:��f�^
/R��Z��f�X̩�wV=�k<>�Bj�x5O��M04"Ul�38�p�h*u�^�1-���a#�\D<!Kk�U^���ڝ��ЇƇ�"��/"��ƭ�o��	B����Ũ�dږL��Ь��C��g2e
������z���Z�B�叔Qq33���W�%3t�������]���H2�')2� ��:.F�J�޷}B�gn�o�ʡ
ó�p;�_L�M	��i벩t�U�B�8.���=YkB�]Op���H���2B���ࡼ  3{��̎�F�*�u�f�d�4�ỡ�k�2��&��4�mkvz�.�k��xh���x1������H��b��%��>���T"<�b��ҁ��)F0l��<�9�[t��"�3�]��5��g��bqLC���Wl']���v=A���	�T|��!���!�{���w^#.nU3j�̅aږ��b)>�%CZ@Vr�����+x4c}�s��z�I�u�w�f���r������JoGj�(�_���F��R�P`3�0	�l^ڪ���^u��|�%S+���ٙ�����SQ}/]P�7�>�*�O�q��q��tϧ~�����=��dX���?��s7'��|���{��'�&ymj��|�9���:w�Yf��a���{��*�~���>�!���� :�
?��kyL3�t��2�r��B�h�:��nB�qK܍j:Dm�B~����?Q}������e|������ˉ޼�vY��ʉ��^��"�Ћ2#�|��c+1�܄���1��(]Bq�޿Ҽ�Y�L(��7-
;a���;����m�N�,�G-<�O���Җx"�a�U��{ͳc��$:`�#��
xDo�PZzA��Z��g��dr�����o�q�v���]��p���#��z�*Ƌ硕�(^O��7��a�a` �!e������U��*��H|^u@d3~Ǻ����m��\�
�-�E���� 	�M|K�Hf�8�cw�:�&)S��y��c��2�yzs�l~!�������HR�Um�(�s6��;��11"6)�	b����[W��|�"̻Ed0�0�m�6.�k�y;h�g;z�U�~VI�U7�S�:D��CߝIIW"����%=�y��?���YB�
1�Y��Ԉn�^�m��(V^��*	�q�]tDk�ź��y�q�b')򬫄�-]���Pt�5���5����)?a[CS�8�w.�^C�����zz�!k��p����mtͷ��z�ل� ����`1R���:�uO���ꆊ����ߞ��`��jΎ�s��޶�B�Z�0Y��웺��f6+�i�穚Oc8̀�|`��f���E�@Ӗ-�4;�fP��f�fB��B1�w�;�K&�|�2��M��d<�	�p%��+��on�83�>�jX�un��4Ω�Q5ɕ�l����;���ы$H�\W�����!�]N���~���B�����J��Ǌ����aңBܬ�̊학�㌁�g&�:�n8�;ڏ�����͉�V�v�b�Җs=w#}��f��9}8��s���c'��[�~��(���L�� S�m�S��LfJd5`_S�����S$0d�� |��ߟ���n�}Z��#ҙg�bzmk����k4y�j�^1�^��/��e���2y+�]��t)bU#Ô���Tw9m��K	�!s�F=�����4��i'c��W�/J�YE��7���t���
&�ί^��-�)H��3ёe�N^�L[=x��;�����[R[���.a��%�L7B����k_e� ��
1���]Ɵ���|���v4;�g~��M����n"��?�9�]�ɱ��69���U��U_[ʬ/��	�L��1\�kҋ �%���}t���"T�k8�r�q�E�;F^O�Zj+�)��Cڊ���iTԀ�$t�n�LL�z���6�r��>����\֝���/w��n�|<�p�]m��Ѕ�gn/Ͱ�86׸��)�=��a����UP]���V����G��rϤ\��÷x�nǖ��hzF	�IoL2n�n�aO����幃x�
Ճ�m�WK�̇ڶ��|#m�k(q-S끻6�g�5:�i�R���z��_�N��VlZ��yuUR��$������T���)=�,�;Z�>j��]ҬA��Ք�T��h�sqW*���qB�Ϙ2���^e�0��<�����֥I;�Ҏ�%���&>�"�����١��qt�����έ���WpT�X�__��&ݽ��jֲ��a�+J�c1��N�u+N��>�^S�Ζ�Z���?��dkշV$y���oS��9MOr$��N�Ƅ㴴����XTe�b�h5�b�����t!��q޽#��qLK.�i�R�𔮲�R]�bu�t,˰�\񍗽	�Xs���d����پQ�0M�s/^G�������p��5r>�X��W(o�)���L�\k��>��ݲ�eb��=\S�)t[���)�n*\�+13���E��������J\��!apj �s��W��b��r���
���+�J��Ver� 
�"���Y�d���.����w�1�(5�GlKp�����
���"�0����^�ؖ!���2r�R���V�+(���3ke�Y{��[z�̈��J��M�y.P:U�����-
䌍���#�Q�҂�dbܷ��]Jl߷t�u�u�2�X��ZY�m=QR;���ڋ���/zŻ����wp�E�(�Wua܈}D��N͎�j����h &8�[�v&zf��L.G��w2�f��E�ҙ��� E1� -V�^(�\���ر� CE P�L�tA�B �
���n�J���*��ڭ�R���%��Jo6�:udG�T������S��9(�ڭ���s'tȸz���T�L�U̪�]�4���e
9R	�-�u*��z+��xJ�ʋ��-�}24\�]J��wԴm��xۖ����l��hP
�C�GJ��|s���]J�f�*�A�] c$[�kȈ�gZ�:��Sl���)��Q6S�����쏋�]�ax ��&\I.j�=����v���:�� ��\�����bHv��Q��؊g�S�B���󏷷�E���$���GT�ЭT/n����f��3�����v����.����!���`Y�]Mf������k��1
ozr�3e+�3���@K��1��V��u
��l�p>���lX� ��\C���K�k4�w��a�(���N7MtYu����&�(�.l;��4[�;y�.�:țA��C_���Ρ��:�:��kn��GU֪�
��!DI����`����Pڸ����\MW1}�:q���Xr=#jY����*��P���g��[�;e�u����-�fΦS�eFe��}Y�0�
|w�JS\�jor�b��He7V�Xr����7kX��v����3+5V]�L]
w�K�����pQ�g].^E��^�ċ��G#�����󼌣VJt�@���)j�H�D�D�jK�IL�l���F�p��*vj[��e|���	���F	.�
]"���e���su���s7��wm�.~y��Ou�͋��{E�ӖY�71���Ԋ�̈pݛ���UY�8U�wv����_^=|~>���?G����3�O�3��p��2�����p�7
d��v�nfٷ�ǎ�|<>?___�������j�����W�KE�3,)���U��3LYeQ�5�r�3��}~<~>>?__��������a�bTM��a���c�0�q̓��XsL9�A�0�&���f�QG#7��&.�9e��[�g0��2h��*�',�����晙�ea�ϙ��c��6f$_M�f'0��4ȉ��aQVFE�`fY��c��|�-��/�a�VU�T�7��|ܶ���
h�(��
�
��fE�³2�ZF��UXy�2���QIU���I �XI�FfPPDe�f`d�QfX�NXUTԱ�MfaFFU��SPVYE�7��c�EW3�1��9FU��jA�+�E;�/4�)d�m�_o{i�w�6�|3��U�G��ֈ�Շo+2V�F��*�����Ю�u����haW��vŖ�^�����-�e/�ʊ�N��A�a�eT�2�K@	�>?�3��O9�,~U�~^y���חzki��{O�[_�@�9a�)�ª)�|O-���GI�ܙ�Z��9���k�Q�&�x{na�<iy����NÁ��CH̭�j=;�t�D�B`��ٕ'�6mS^�ʭ��[n��X��p��3�Sa1�md����U��iE�^��]ش�n|�BL����Lsm+_�k��ǜOXh�O�S���YЁN�5ɩ����fʖ��I෪��*5:wZ�y�n�c|Tc��g����dD�mpQp�Zb������7��u�ɽ0�7X��- Q}�h���+�G7-���R0��o�:�w{х��coUt!����)~>�|����r
ϛ��'�	�P�(�����O��3��:n�?7�-ڻ��A{]�s��'�4a�J_���/�ǎ��<���/���f�#ߍq�f�.~�Y~s3Gg�q*�h�d��~��\�w�>�F� b��4r�E�
4�c��	��s>�al�ǅl^�հs�ab�D.z�.�~�5W�(�])�%�#�m
��C�!Q��\���)aǮ�ųF�f��Ыf��*b���n�e7�?vj��]�;�C}-��!��OZ�cW$+��!��c�1�\�v��7Oj�� �Me�+ّ�ٹϚ�=�hB��3;��߅q'�����צ����S~9���o/�}���0ʂs�����߿���}�
���T�������1�-��"�QI���m~<:0�1�|P�[��Y���8��S�HS�u����l8Ϸ��3!�+:<�f�҃u���
���Mӧ�p7��ƝF��\�z�����Vx�6��	y���=z��wP3������GU_~���ۮ#�,٘�~��a��ZH����En���o���:?�/ؓ34����mQ-��s	mܿ�=��0��+[W�m
��8�#���LS�c�|��&���-���QX�s-�Hn�O70�z0�:������"�8��{m��v�p��h��03mX��
�Վ��������2�����S��`���
�./����(LN)t��<�ҎJ�L.N�z1���8���7"6�e.����)>���k���9N�>���.]�>f�%�/���:��E�k����#"��(��#q���P�sN<1i���CVJ�>�\��.�/�;y樎�	������}+��C��C���`��/�Z���g�����4���ʘ�]�W�=�>���8�_0*5��[#;g��-��u�����^�YGo��c:� n#󢈃^S�Lc>�&��n�Mīir�embx�eX�R����0���=Lf\L彳��'�5�e��+al�����p�\ހj&���������p���,&�y߇�������s>i�.��
C
C�x0����²���#���}�ϴD��Ac�fg��s�i�w���9�o�3Ù��?����u�U��B�-W0ٛ�"vJj��6��X��	�su�ݎ�A)->�n<Dy�]�<�`43���%ƣ�I͛M��xs�l�e�jv�P�y�y�_��^��#r�e�f�̛l�ע���*hs���ԚJ�V���������>�ܽfw�
�K�x�>��\@�:;�Ѐ˸� �����`�J����w��c܄21��r�]��p7L�e���{��UIj1�yo&�J9�x��Ŋ�'���k��炟ɫⲏ�)岮;�hNY��qҙ�׹yTŵ�w���=Z���c� �.�w�1�މ�ѿ:k�D������V�,�d��㸻M.��]��p���f������R%�t[�牛w�KÚc�R,�b>�:;F�n��@m��%�ȿ���_Wi�L\u.�,u���\&�J�Vj�jcn2��{!t�F�}����LE�n����0����K��,9��k��L���R}����8�S�n�[)�����v̹]˯�m�=X���m7�2'U�y��Q{�̮�����to)V�80��f�=�"2u�>�~E�{ǽ�)�k���-oN]��@f�ٽݖ�G�vĝe�m`��B�QR�����X.8��3�Qa�s�79����C���	�0��J���ӚN�OW�E��\H��i��-��wL�Q�T��X��Gʙf�z]a.`C��B��(<� `F� cT?'�pCe��1Aקٞ�P����~㿿/��f�~G"�v0w�]�QF���
���D�@�y�W��|]�����<�}�M8jC����R[�C�'���Q�f��\ֵ*f�*V��P��}}��qӌ��4C�����^E�#f��6�;S��:V���ͥ��t�FK%�s<�@���}w�q�ə���^i��4ݙ9u5�]S�ȑ��M䒑W�:x�y�^˧�Tw>5�(,'�֢��Ί��@�O:<oM���r~ռξ1/������Ao^�ac7���y�|�}�eh{�S<�_�hϽ����|��c��Mu��M�w{�0=k��ƾ�nߌ���+�c�������t�EY]�i�>�iSYN�c�m�vlt�"fXl�u,����>h�41Lk���m��Ӿ�Ϻ��]�y���n��� T! ~��h�m�^�'�yR����.��O@k���Uo5�x�u�T�y;�^*���kV�if�{:�Em�o�
�?D|{޶���n������g6�xd����2wz#���@^R
�Ub��;���I�y�����7�u|kXM���[�ʌmn�V)uқw��p���)�7����EPT����o�̬�˛����a�C���<0������[�
��|�9����4�f���L>��=z_%�9�$C��O��~��ǃ�+��)����}�������%�c���s�	�p����ٲ�tñ���Y��.A�N3ܕ�� �U�<�ck��R�M�lh������nl)]
oc.ݑ#�̼�z��j�jY��R ������TŶ������=.h�O��GyU�mC�Y�e��c{t��"��w
�Q3���1�ÑNǃ&2ɨ;�[K�Ө��.����ꛦ����{$�yg�㙏���߹�r������yj��@i�^�	��c�h�e��I���U!�C�Է.4s���_X ����`���'P�.+e�Ʃg��*|�9m�	���������%\Pzɫ���&�-IN�@o93���	��ZQʹ��4ǝ�Ӽ��&��]^�o��)=5�&S��Y�M����e"�y�6I��W'�̴�7c��������6lф���[h���ȯ�CO�+:I~���W������G�����4�*/�#��c-
��Z� �qW�h�E��7�\d�v흁����6I�t\�oۺb�$dЫ�t��o�.�����l��!��SY�u3+��Xr]�a3^_K��'.sxQ�(��%0c#�9U�"�X,�M}�"�uk
k�����De�����aa��Qr��7�=���y�{ҿO��y�4��f<�?A/@K�:j����Mx����=��z��a�
7�kbD޶>vlP�-"A,!�k�@�n0�l*x�����z��&�1���Rmڐ�YN��|V���&������C�3Z�F��T0q�]�`t�Z錡��:�<���/�l�+�zTDS��dot�!��mlw��#�4�I|s�O�� 텝�l�2���y�	�ɜ�Vvep�"�N�������udߛe��2m�4O���jW�m~39BPa,�#�v��)Ak�k/i#':�z�/L���q�ME�܏�]Àѹʅ{� ����{G^��ܺxjQ���5#�h�.K����~U ���_��>�TU>,���q��b��n5(�V�x�R����Ķ��I�$4��;k����B�O��W͵S��W, ~�_U���ߠ���W:�ߝ� ��#�X��E���][u|M��Z�׆�[;�D���;�s����rD��g�kR�c����.凁�0�+���\�룱I�	k�9�v��:��l;OG���F��N�����2l�%���E��o��l��W�*�#Xm�C�����3��� U����B�!��?��ۮ��;�����q�_W3��F5.t�K����8;�g_ Û٤�/@�DJ<�g7��H�����]��\)�:���ݶ2��c
;Tx�ʱ�_�`!��|��~}��������(��;�P���V��(M$��Tט�[#p���L���f1&�j�b�Y���������_���z�C4{
�j��F,�Ry��x����n��m«(�G+Y��5e��E�ey����u�����1h�ɨ�v��"GuJ�8ǒ0��6:���ODR-OX<f�L ��w��F��?b��W�&?��>/����9o������0��fk�����(V���6Px��=|&�(tc��|c%�Qz���{�X��զ��3���֞ս��������՝�]x��0�����bF3SlC8.��0������;������.�^��Ntrq�OP��Y��UK�>>�4/���tWx��c��3߯��9EUHӛ�*%�P@ȋ.n������Es�-�m�>���4\PsBntX�;4�q.�JO�U�p�,m�b�����>��f���՘f����pa���8��&�\�4��ŦK�c�����+O���3��xJE���K�h�qy�{r8燠^tn}B�x�uT������K'�]���:�V*y���Ă��e��[DVL���1+�m����i,�yc��(n�&�qsv�O����@�bc�>�?7�G�mݼǞudq6�n�u�n���]�y����o�)#�&��Wgbj�y>�t�e�sm+͒��}����χ=�;߿N���y�<?��VFa�4{� ���!+��)f�j��]��r"��D-2����b���jĻ��rb�����FZ�/T�\�%|�{|�.������T��3a�O<����-��Ԕ���Fz{��fT�g������dG7�y�4,a$��
���_�vW�hy=�M��X%t+,j�aMKr^GT<>���g��{3z�Ү�s"ꑜGj��J����-�F������0XFؤ��;��jv���/��(�z�'��/i�<s|��ث���~�_��?<W:}�R}§ț�l׏B�e��ƪ�J��޴�[�O����}�*C���"�� ���v,����70���&�c���˟�������9\�k҆,��sK�<p[������Ž�GY�Vd�q�0��R��]��zN�R쾁+��C�e�Jn�v�!)8�%=�y���y>���xM��!4��A~Y;i��f���uP�
�Tb��@%jkX?��,���h(E�;<8��~���ii��6i��F���YW-ڪ����&��\u��C�l����=X�U5;.Nt*�d���>��*��M�R�2�+��|��,�S�6{3�@��F�=N���`�]�˹��-���.&��{mu�g)"چ�T�)4HWԹ<�;pjΡ,;��]��+Nn��f�t�3����h˜]�#�hD��9R�1��:�p�:��Y��}u���R��@L"�sw.fZs����?��!�&����Il�{i���vE�O�����^�K�S��M��u�g�ӳq��h�45��x.kֲ�C;�Us۝;���?U5 �TP��Q���-��:_�G??
�ܼ$����gu�q��a��^�M�v6��P�c@Y����^]�k�1���	���E�Ƒ��P�qǹ�T�(�n$�n�S�ql�1���Y,�ޠ�]P��@n2�ǘQ��c��c�=7+�L���)��7�M�:f%�_ lw,���H�'�c�b���L<d;�K<�lw��y+�іq���ӻ�u5䩬��l���sz��8�>�6�B6=N�F�z��x�����&�_[ݬ�ۖKk(��xa�7�n����H��)���M�ԉ�Ս�+���� ^�Sb�:���y��[�)������E]{�|�ǂ�h�[��ĲԦ�km{�~�`6P,���g�0R(�5s��n�;�v_��`��e��_����<�Xwt�e�ڋ��<�Ȋ��m�n��g���<��&�QQ�0(^4RwaZ��v	����k[�c��
��'�o7	|�0^4t��=9x(:J��������٦�#��z`�ݹ���.?��M�rgUP}VW'3�{�hgZj����=�xp��boCr�gHb��K9ϝG`[��p���'w���ߜ����{��y����0�����<��2��J+]�XR����L�,#;����{ߓs��Ů�@��1����(y��DsT0"E����[�rwE!Lg�:>ny�qO�x��a��JQ͵�k�X��@����F���{���t�1lL>3z�]�Ź���fKz}e*�M{�'yc����
�nj��8��~x�S��v�ƮZ��i�,DG6��zo��C�w���λ�k�QQ��c!@c~{�N�	���X���9�2��W���P��ݕ� )���4jΚj&��hVyƊ��{��ʦ��O�HG�=Ì�H�.D���nf�z���C�(I�K�azǤ�L�\��MZ�N�.��슠�B��e(��}a�;]�C_t`�@a�$aG����>#|/��C�l��Qb7�ѣ�1r�e@��l1����=#LD��1a���b�<3`N�V�'b�Em�͔xf~UO��\g}̼��d�nh�(i���$H�%M��!>s˾��I͹)uh�r�cܘXܙ�^s��7+��\v��;�ߗ�ߐ��PU�󰨟�����v��Tfҥ�ti/u��v�G+Fs�\����_�ݷ�=�*ޏ�n�wM��Z���V�JFʋk�UZ���*���=o%����bh�s��L���"X��ց�]���5�E*�A���F�[�u��ꑥ��R��]��6S��f�j�l���e��Iʽ	�����s��Z,��}ǘ�I�Û6p��Nl»O4e%���z�5>������S��)[Y���׌��潺m��ja2.k�e�:k
��'�&�|�9k�"��0o���-���-.�[xF�i�ʂ��]֯6i��D̻�h#ҝ��=ɫ��;78�e�"!O�Wi�bm�uM�6ܻP�\2��+t�Yu5�ؕ-�Ͷb�|��u�1u�9����u�v�Uӝݍ��ӫ�lU�5�ʾ��C�ɸ%v�m#<|�!���t���[a�u�C��b{Z����/�z�ER��ŔN9ݶR��w�O��	r��g3)n��B�&����f�k��g�p���cjy��k3#�4�aD����s$�y�Ծ���r�R�̕x�盇Q���g��ৄ������^�����d�Q�4�N�����I+�P�޲hL��ݵ��+=E}]�9�yx���9y;�Ү�g[/����Ys3��FӆI\�b��P��PO�i����V�V��mCUq�ݳ`h8��������j��[�UבK]�%N�|�}�O�0��Q�g�g{���E�����N�Tf�R��t���S�7������˗���|�jae�}�'����6!V}���:G��1{z��!�]�9+
:�$���dJU�R�;�Nd!�[ �����:0�ijã_�z����b�3��h0a���=��#����M���)�r�^N�*���5��V)lG!�gQ�@�d���j�u�׋��:��I��ܜ6��A� ����:h����ہQ��b����u<�N���/h�}�Jn��lYT|M�%a��0���*%��W]��������d��xʣ7��ə����r�N��݇�!}�ݓ���n6�n��Y9�MD�G(�R�xvl��ڸ%^���F��p��S��sެ®���F���ن��B�ş�W�X��iz��Jwuʳƥ�PgK���w~��/[��UL}��ƔR��z�y�*f��)N��t��]�ZN@um��⒥-�(hM*a�W�5Ry���;����Уvm�F�$<��0�t�O�g�ib��Kl���A�YOw37�����%��%�ȹ��2��L���e�9n���v_db�oh��7�1l �#�r�C0��g�'�\��D��n��4�F5uZ�;ouʙOH�1���s���7/(�K�^�a�:cA�;u�*7���YŸlH`��e�>�[��z�KӚJ��c}�ƻ8��b�^L'*�P�&h*;f�g4�b�l#3&�,���0q�

��h����̢����^>>�~�>?__�_��q����h���j��aA�&PTD՘fc8eF5نg��I2��3��>���������f=���f�DT�˛�7��;lÆ鑘X�{�F�fVQQ�帔����^?_Ϗ�����������~��De��YY�t�c**�����(3(ʌ�-��,�����.fEE�y�e��%���k1#cu3321(2�2�2������e�TfX�LDE��Tn���F9eS���n�y������NFUQ�QY�%YQ�4�e�0�B��2r�G��e�r��`a[�l�m�dTAL�F�A��s*&'`�����"��n�dD�UYeLS�}p(ၓ�aEF!�L�	��2�̪��1�f7�ӄa<�b2�,b�b�pƛ0���9��9�W��e�y��a�f�L�Ue�J�����y_eL8󺻜�%������s�5�KH��>�G�tf����&�:��s�.�{�_����e�O~�_~K��?��s*��mT����q}#�tg�<���o��)���v�Ǘ��
y��gv/���5%��2���<\�sw�#��lP&�"��Ɨ�P5:���L�� B�qSAe%p�tc�l�l�sv�-�VP��@����0�����n��2y�UBʿ|��Zf~��;g�wUy��?cȣ�u�)��H���u��gh��`ך=�魟�rڟ+��rk^#yi�٘٦���h!�ʞ�P��S^ʄܱH��6��?Gk!�6<�.CE[�f�Mu⋙����K�l}�^O3Ft�h�J����	0ZS��%8��B���$9[B6r`����}J��^��a{A�J~�A��[�&�+�]���
=�E��ǖ��d�湺��`�sv���_���Tz��(�Ն��*��,K��Y:��6�K-�0xxAT1�twa4�oI�����ӎ���=)���"EV9�	������-����E'i�.� �{�ࣅӑi)�Wӫ�	�O����j��������v�����3�4
�� ��K�������L����>�������E�77�7�jc����v�T�c�s����=�(���dr9/y�{��f��������K��!y貾�[-�ZX٤5B�e���K��u�1v��*M+j��wF�=c��;7Ѯ �/�_
�_
�<��� ���UH=z�=<�^#6|>��$�/�z�5=/�m3:Ľ3� ���HV���yՌ^����]�g�̐�p������:��!���4�8�0����З�A5��V���'�w��7��QT,��AQ�񪿤���-�mcY}��ݕCls��``f|�"︡L�?Wve���I4�hס�)DW�Uh�J?�:K��w�(}�"!e��K�a��J����߽�[}��iW\[6�Hkͻ�6��yח�"c!'�Kտ�5����+X��{���âf<��QͰ���
!�����!����&�JK�~T�W�T]�Z�8�<�����s���tm��A�=Y��@%u�g<��Q�HΠl]m��l��~9n�g����^5��0��5�ZW��t�_����$f��n��v]��	�ɸ�ō7�]���F��uE���@�2���3Xʞb�8ɡ^脟,��GT���Ɨ2��^Y�N~�~��~���g	��Y�X-��Ldz�����UY�{L�:�~?�u?{k����S�+~L?����H�ﹽuy��"�h��W.�*^(_X�)u�(v����k3E΍/�wOb9B�,�)�J�@[�����c�Wv���u�n	�8i�i|T��܅Q��-�5�$f[�Vi�*�g$9 C����C�
��a�YsM�6��Ἄ���k3�?�!����9��?�����>Va�~�}��3��_��1}͸��C�D�g���}��c��b|ѭ����j�U^�,��XÌ�6s��Ժy����qBsCH�@hzg��Ze~)���_����?[����K[zTˢ��50i�j�����2�c=�qN��Z���;�f�p����a��5�Gz�6�Å��Bpm���R'n��g���*;�e������^l~lٸ��x�b�Q�[���o$p,���<��&cK�C'�����_v�[��ć�J�6�nn��yn�=qMx�b��<�f��1�Ґ�]0����[p���@�8��ܪ�/��)k�	zcWTvS���p ^Зe���ܰGK���K���?�l+<�'�r��D#<܌�vf���CX�x�XS2�TZQ�`���Z}uI}�~�I��<�O�����F��ya�;,��[��i:����|d@�ƫ������ܶχ �*m�O��gOC�^���e���;���[O|�7M���i�ۤ{ )��ȼ��5t-��Θ��6�(�wRq��+w��W�`�����z=K"�2��cuڋ�����69��+]�u�Sm�@�	/�U�Y51vr�D���i���ccEԝ�J���-�䊔*۫}�,0�F�(��K�^D����x����&:�⹴]]����m����3��;���g�����1C< ��梯˪bZX���T�M3QLM����	�zʡ-�8&B��ڱ�Y�<�ECr�Ӳ�$C	��?(Ӡ��7>�U
W�����K,��n[4����K�Z��-Y�X�;�Y?J�c���UK>0U${񹊿?k��A�w���ֈ�{����v �S"�rm��M�^���"���*�\Pw4ԋ�-z�?���$�F$'�m�t�Z�NbK�L&���w�q����w.5��zk�M/t�aX�b]8�GDY�'��-E�d/zCϷ�s��\��|b_Z��*\�8v��:��gGE{1|M��/��z�u~z����D'a^^tb%�I��^�c^��k�
~�U4�W�Q�DS-�7���X�F�Z��oWV��*w^`l�����0~a�6�T�dۦ���5}:����ESanK���BU�"/i�t�b	`��f��03w{dB~/r�Κ�嵤z3���Bl*�*����qb/4gW=�ӈ�4�]8�H��66���zCϥȔ��s{Kȷ���P'��N���ѵ��ۤ��5u�j�w�.X�E�'Pc��%�죽�i3����W�6�xd��(�P�j���.�Kb�q%ڲ�sBݺ�R��{��]��ƥq)L����rt�y���n(���V�]��ww������VH��I�P-�t�u��LO�����^��t���Q�L�N"�Ȧ�����)K�Ny���-h��_�&��5Ŷ'�w�Vro����"�jDg�W�yV)K�'U�Rc|1�VgE5>䗞Zk�[�(�36��a��7@-��C�Se�����c�����d��m�Mn�Nġ(wU�ᴚ�߮����V�3�z��"AQ��{��i�|�X�}A�3�}�����A����p��w̥�za�V+]��G��o�*�*g1��+��2�w)�v���+fǲ�n��a�������X�R6_���=��Vg�\q����]�,ڸ�C��,;�5�A��T0r�-e�e���Y"t-�w��ᑉ��,�E��A��v��I��"��s��C_oY�z�5�d�<u�s�Z��)?^)�4��Q���)�qx�ǃ�r8�$�[6�lmOEm[.�5����@V�'�^�q��J��BbqH�������"g��b>B��W��:�I������.��
��OUq��FL�h�ɵ��#^�� ��{�Gňo;�zA�5�v������ �[1���@�*��l�ii�zG��釴dڻA)��S�BQk4��3�T���^`_�e�Te����Z)��r�~���������m�ހ=u��%���q˩R������mI��Crͬ��$y�q��U^.�8#um��g�����y���v�ʗX�꣧���YB|�/�����.C��M>��w�R;�9�kܠ�zqww]M�4�闹^��B�>��oǡ�J�tV�k�FW�ɏ���~��Cr�V�y��(x�O��5�"h4C4@���a -�&�ۙ��'{,b}"Љl΍w��:��8�*7�����_�P�Gi��V��}��S`J��a�����Y٦`�~&y�ס�����Qu� T5P9��I���/���އ�L�2�LPǢ�s���N+I�P�!��5Z�L[�^}N����4���Ti��[�*o���Z����6[��>L����_�;C}��ͽ��d�H�厷��X��s���դ�EP��Q�|�!�)��v�Ϭ_>�����ב��V�xv�8ԄZ�q�l@�^���h�][�3Ɠ��(���7i|�����Ⱥ9D0+�lgv�A�p�9�\���UHnͻ�mQ0�/fda=	z��s9 ���r��F���j���|�<`�Qn�S�y�:���l�|����IL�̦˦�j"0��A(��j�9�ca�v�f槖�%;����}�,��Õ�����5�!ޏP�Ј��sz/����h����DR}�Q��H�9;4s=9ݐM���]U�u�G��W!���떩<���6���v��/�˽۫�UɈ�-�b���nY�����7����?��!�����yΒV�̜�Π��e�����3a�za �I]7��ƪ���(���W��� l�~ڃ?_�3}eʶ(3���<)Z�,�u��	��rs�)��H�
��ua����w3���vUò5�8ޠ�[[$�1fV*u�����S愧Ȕ�{�7p�����#?V����2T�ư�8M0ͤgy�vL���e������Ĵ�겋ԉ��]������2���S�n�6]�p�O.��%C2נ|�2/�M�A�I��#9o��r��IM���7�����Q�ڜۇ/����:�/	��󾖔�دseӓHC^�O)�_*����� �%�g�Z�lj�.�1�#X�,�g�v_��>�iBb1�=0a��=��F�V����z*;�e�����\����}1��ދ�9�n��jg�J��b�T.�[�ϙc�X�>>�E5�d���KTmO�ծa�@�b�٦�!�ضr�]�ig�����6�a>�,F�u��d��
1�>A. i�-/�#�����X�j���d�fj5ί�ǎGAm�'�^R6����
F�,�CFw�M�֧GW�֨�<>�|\��oxfM��Z��S��\�y���m�l����z�u����7����ػ�=�q��E��7w������41�'|��~��xS[�k�t�>�� ����no�]ٵ�(��gؗd��E��E*k��WS^�wD�,�������w����d������;�>�|uQ��ȉT�pf>M.���OJ���0��p��6���we�_Z�!6�,`*m�I3l����S��xjF��J�)�n�_+6�Z���/j�����3o��y�/1�71�Qn���i��f�I5��g-���5Hg�p@կߎ1F�L�m�@�6p���0f�n�c��]\w3M��f1dz�z$���l:&Ǿ�
�%�L7氡J���ږ.j���Px;�%��?1v_�������{�:K�l(����_�ݐ o�}��~U�+���3D�芻0��-8����2�w��*�C����V0��2`��6dS�r��5��=��M�iL��s���yr$C��t�4'L9*��ؕ[m����-͏Ux�aа1���~|7�w;pn���r^ς�a!�_u.����ci������)J�ֵJC��J�et5Tɾ��:�{�w����fC��]���R7֭,��y�,Y7,���;��Λ�*x\%�o]�񬼔b䖄f�Q}�^�t���ɏ���������:��Kpr�#V�W�Nw
�黙��f��0<�<�.��3o*�
�����Ѯ��xe1F�����*_��K���{6��=����x��}������<k%�Mz2�SI~�!�o�
ju��C�'Qn:�6fK��;3�e��;�|� ��Si����9���A�����K��-^���|薬���w	v䭻�t�^o,j^0Y����l��]��N�0k��;΋_�L�����$U�k�3�ʺu����Xfk`�	4(���O��Rz������=��J�>U�'���	�A���~��Oy��2s3i�����X��	�t��\[cP؎/C�H� ��z�Xga#b����<���Nc`��(n-r��i�,_ŏ־�S����|��'�����p�q,f���wy�?�=ѭx����B>?��'��LT������c���|+�b�'��.��s��N�e�Z���DU7f��=�E�C?�+j�y6��ֻ6�xK6��ߌq}TPV����g�����vř޴����4Ƴc�_�-�eC	���$��o�sX�����Am���O�w��<m���wu�oN �ǡi}�;;B��7� �����q@	�6[_J܁��oy��\;�ר���۝I1���S����������W�u����D�V�-]Ox�����X�a��6��>�����,ź�Ȯ��+몱�<���0n�X�\!��%n����^6h@���gU4,�w���̇{k���a�?kΕ�.�36�\Z
h��@s�ǯwBe�~�ń�s��Y��w�(����V?�������/w�n���{l�q�/_�E4��oH�ph�cO���tQ��l	���_���h�M
�wY���:�u���K>{�GDz��>��3G��3F%:ͮ9����߻INa߯�n��%�-��
���_Q�V���>E�P���9����~�z�˔��K!f�ۙ�?�tts��?~�ۨ�i$a�B�� ��@�҇��rD��/�Ai��+.���.E1�]{*&�WO2X�}�Seo0��!�4j�vg�O7�zw4��Rw�J�;/�{%�
t�L	���cӑgg�Lso��[�Gl}��� ���hcnp�ѣ�i�٨_����-lhǢ���12��V���2�q66ݽ��Lζ��3������NU<ġE���ؘ71ݚ�3�wi�dy���WG��ll� vA�����j��s;Ӫw���T�2�|M>*to�������r�w�Q[�Gf��\�)�u'L֞N| #��&�3&����F��[�C�3a�*��#yu�$��At�C{{:��y���Ü݇��[�$s��d�Ok�-�}a�"��=;k��b�6�b-��WeJtde� X����VEy1ꔠ���XUb�dL�쐊�X�iL˳OC��;5n�n9����4)Ke�֪��{�*�-jF��O���΢m�� � Ǻ��ʂiEs�hj-�3������-1�M�Cl��,�w$�֐�����15]���v���ۢ3�_w\9�-,_}��fP]�W.\C&c�yT�٨�%
u��u��FnX0w�C���>�h�ͬ��
� �}��1v��C��#��B�B5a�������+�;\ k_t]�i�]��K�����C(��-��yr�Jݰ���@'jRlk�xWv���onn>�j�;v��}�r4wO:e��8�i���k��A����{.��85�����Oz��uf֚��{oK�����k�"���f;
�Fs�<�#z��AC��9���d1ӻӬ�O�+}��x�XhK������tT���̕�%����<$�h�����zV�G#Ҭ��t���-�lNa�/�NpX���]w(���l��mv�%�e��*&�J���3[(�*]�8���8��)�ڔ�͌�����ubwxO�Ԧ>�3���-��GX&GC�,�Oƨ��[n��j���x0P��K�+�n쵫E��ea�fL� ����|oYt$W�������,^�1�c�0�p��\���ŉ\�TGG�i����o�3:S�r��|�*17�U��V`�R�5��g��5�W�Q�Y٭���[ݦ5j�ֶ�;�;����]�^���u��}�8��*�Z����Je��fm�Xn�v "ͻ���i�F�7}[�.��R�"�N�)��Z2>�-�g32�=��,��G�y[���
��ի;�o&�MT���ݗ���� ���ݗ"�Ҩf+mED�z��XWυk�� �6�v�l��"�ky��#�0�_���څ�b�ܴ�x�/i�5�H ���u�q0d��.�q�Y�\��{����-h{j�[���Uf���ʔ2_7Ԡ��T�6�:Ɲ���}��]�#�-*3�[������$�� ���>�]wVtO��G}���Lk��jb �p+%��t�4�5gWN4G� �Uأj9���V�V���y�-s�)M���r�v��_<_n-��$r�<�yh�W�=����4���}�o4�U3^�I�F��ӑ�"{If9|�L�+A�`�Q<�v7�!N��˺Og��Nv�cmu;Z�q�:�u|⼽���4J��E*W��7Nb��B)��{s�C�w�:�ܼ9���\5�e] +�8��䡥V L����m�Į�hHj!MA�S��i�sw�0�ۖf�iͷ婶I�P�"���"�-%�6^�����A�w�m���b���LەT��IE^df�y�iSG"���6���_�����������}}_������e~�)(���M�*�3>���'M�)��C0�b���Mm�0���]||}x�������?���߈�����w�E,����3*&��&�"���3r� ��,k���_�<x���~���3��������XnYa�G9���##, ��f3�Ȳ�XQ�[�EFɓeF��8�Yg,���4m�|�Y�����s
����1��y���y�F��&τl�U,�̌�f�wm33��&�h�d�ɚ�#	"*���wO$9�.XRQY����DEs�����$�
���;iE�2*�r����-�Ķ2�L��	���ane96ay���VS5VF5D����1�"l��d�s2�"��z�ld�S^K�m�1&NNA�:�, ��(xYU9�9�c�$|K*���j�Ɯ��0Ȣh���噹�_w�x���M��WRZ7(�F�ڊK�;�gfm�=]\�W��;���$C��F���U�N^^ uSm�I�`��s��?�4�y���ٟ{��?[�cr��d
�Jfn^Ə�6c3s���|����ۢ?
?�ր���}w��4�@�S�3�f8ܾ�q�]:�(^j�d��%~J��<Y;�QU���)��Ebj�������He$"o3H�2əy(�q[����"-�J�[�f�=�ÿ.E�f��X����<�E����Ae��6��5���q�6׸^��;E�kk}�5�O��/ܧ]�|1N��L/F±����{�v�#=�s�Y�yQ����B���xP.�\U���z�Jn��4�0�X���"�b�����ʽ���Ō��{���>g�H~�j�"o�E��'�驧ry��O�1m���M�r�m����|�\b[��$^C�uPV��h��LH���:�p	?<7:t)L�u���#|�j����4J��gP�u}�B����{��'����?��2鎽AU_�����
A���;�������,	�D'�E訦Z��(��kЎXۓ9���t��m,�k��s�mC��GJ~\u�����f���FCȭ5�(t�n/`�J׳�͵$'pԵ���P�!�P]�NbW�ӕ�7m�b&;u��4 �*�ۆ�Ղ�k�̏������x�o���[_Ɠ���K�тn�����v9y�+=}����,ا;���|��e�)��hֲ~r�(qu>Z�#;�ԣ�u��Z�g|��3���|�<9������t�O��9�R�aH�Z�g'l��_�c�<�,�ҔX8>Pd�X��`��=�[]�Z~�,�E�!�&�	B�\A�eH���?K�iF���ge��Q��,%%���z11Z�t��kk��5�7r�B�`�����!�<�ye".y�>�U�L�d^4cf�=K���~�t�L�7W)Ǻ���Ḵ6%;,���+ ux��hU�C��sw{���-i4�Ǜ$����[���vQ��cШ��}�O*�`�m��^���Ξ��P�7�򆽙��0Hh�W��1�e��P�^�W�����K���+�7��]���V*�+k��v�X9Jk&�OCoS6C.�M��6݇��g�O�s�6j���O@��`��&����7Y��,�=�,o��.�Op���p�T�t�d1�>�4#��UZU6By�+{.Y��ۺ]���; \�M�8����e��ư�Sō�����6(���o����N��Թ�ӛS�o���S-�mĬ��V-��w�m��$k��2;켘ϩ�E�+��ܧ���=�V�q봉ҙ��ʖWJum>d�H)�93ŗ�3tpG1e̜�Gs69u �.n_q��<7��p� �2ntew�>f`��=�J:5)Q����/���h+v����P[j��u\��w�U6)і�w�j�/ݝ\�}F5P0V1N�Z�U�+ۯ^+2&�K>�ҹ��-ۊ�N����5��xWm	�r����aU�Ȫ+/6u���n��.�Q|�3X�fd��U�i0!�:v����vy��sB��v�Ig)lzx���,��s\3*���p����]>kR���(u5Е�"��r��lɮ�w����k���;��#�6�9�0�e��7鎉i9�7-����e ���巵���u�y,�M��!#Sf���l\f#U�]V��=2K)���.Gt��������ͮ��\��@���޼�������)�3hE�{X}�I8�/���fW������l��u���w��VK�Һ{i�,;����BQY� vt�Ϭ���j�|��/�n�ƶ���eu�lVJ�ܧdG��q�W1!�+���|�㟷;��C|O��M�37vs���af�wq��a�/7�bgs�N��eAɴ�W|�sR]ys�Rw.SS�2����0[�=��g���ￍk�C���]�ߟ?\�s�}��﹙������H���R��n��1��鄑�0�xme��H#���z(v��fm�c�q��&��_�-�ܦy+.O���T��'�v�[O���#^|�V޿	4B��8�'���!�G;R��^�������*��oZ�Or�13�:2V����۩�n�
��J��t�á^5�2i����[�n�e��.��UVMGc%�B��։�bFxzl4*x�m��ݗjڌ��Q���K3ջ��usۮ�.��{|U텖�!+a-�N�ƍ��z6�[�3��Uۮ���G�:Ú���+}��yB�X���q.C����F;��r�"Tn��rk!n��V�J�6w"�	�D_)�
c���'�����VTu�����@B[0F���_V��0��.'���[�߷�3��$[��#������;.���c�暈��ҹ9���GJ'����2߾ab�����e�e�&Z7�AOE�����#�ǩ��3���/��z�ߩ��y��pt*�@E|��GS)4�C
���������dE�w��>ѧo�����V�D��t -��� ��0�K��0U�F����&L���Q#P�A�E��q�2������3{he��x�}p���ڻ�z,ɑ]IW���9R`h��31e��v�1��{��16gL�7� \�l_�����dE���H�!Z}������`SJe����v]a��A��3�i3��H�Su�r�y��zyU	�Rm晽b�;E�q���a®�Ww��Z4�{9���WM�d�k�����(A�>^�6;�T�ƻv�F_H��M0f�����qs�iJ�εӑXK9��h@�]>�W
���ɺ�)�������&9�V���2x��X^/f�#x�l�	XFY_s��x��Å"|���y�l����$��m^�8��ُ^���p�P\��QY��#M�k7ә+�w��̫*��ٮ�"�����q��}9w(���@�U����K5����kMl����D����ZV��WH���u�*�n,=g{ԋ*�t���lHxk!����@�|�D�ڗar5�ԃ:��r�Q�ee>*�h}>�us@g2��p�'&�sxk��ƗP����/�]�Fyg����}9q�J��1[Ř蠔�6�fu�2ȑ4Tx��1ϖ��ggS��E�3B
TU�Je����}w_]0�y��ג��>����3�7p��V��c�0��Dn?O��+p׹�b�U�du�nuy�r�:�.b�^�Ba�<��j�Ե�,�:[>�2��^l9��2f�2	f��ʴ��%g
G6��d�\��.�\�L��<�ueYXk+�E�� ��j�q]�x��jݽ�U�<���,��t���-��6Ǟ�}鬃 R1�:g���(���{�b��4V�F/X+Y��z�X�X 5t޸���eOlZ3#qq���2�.�����U^i�͏|,���Qa�Ѷ���͏>{SHe�b5LB��}��Vs0m��Y:�B�f�ø����z}z �4�܎�nz}cO���`q��t���JY��%�s�W��(~��zi#͆(��>��g�4%>}�w-P�[`xgk̮��!/ �3�0y�6y�O�<��cA�ձ>x5�����_w�b~OIS����Ư��������#�ҡt�8�ZŜ�a[9������V�Bꕆ�$E�־Ы#�ٸ��]��ފ�0������K�Nww���&bgTl�e!�L������v��>w����{�y��?�0��b��R_7x➾x��/�E�����fr���9��,r��M��z�0����µ�Z����Ebt�z&�ׅ�.�r�,#<� q��ѣ��e`i.;r�6��Z#��΃,���g�,�S�(;�z�����|�gL�/��{2�f�^��)�-\�u�T�-F|�pr�g���-��W�`�����]���)������0��^�9���x�W�j������3
~W���t`�H�Ϫ��xB;IƩ�'�_WЖhJWP�70K�e@�|�e0i�6���Os
��z��e]�8o�Ӛ�oF��s��&3n����M3X�.0v��z��]�,�&��ǽe��
���h䌶��h6�%�mL���Gk�H{��rg_��c���`K��G�S��ޛL��~+�؞�����ǧ�ݙ�9�\�ܯx� ��<��f_��I~ޔ��ŋH��IR~\~��F��5�����[ީ �Gή��m$�+�O͜�:���D�6����#>��RF�ݒ\g�]tY[(�\'X|�b���2�;�yb8Cŷ�����.��l@Bw���l��&��Ds�_e�m������}� ���;Q��+��՟x���(����'p�7R��B�wf�捇T]�*�懻����a��{«�&dVn�
�s\����x+<��H�mq��O��N��t����}c1ϣ���ս���{o�.�a�ok������炪���*��m���v�'�x5j��z�v��˷�{a�@'Ix�z��U(�����������������r��3�����m�7�M
�M�����C�=Vcaᚧ���K�h���a�16U�U�#c��t�6ULj7N���3��aT�d�u~��{�t1F�?4�k�`��ܞ:�M*�~�.��$�[��x���-�Z������z1Rf�����{-�xNnˮUJqTw+�c�q�d-J��[2��ק��z��EEse�xl��.͝�/3\Cm�?N#���ur;R�9'jʬ*�zy�
���z 0��i���>f�N[��<L�R!���K���3�t�6�-�B��;��P�+ޡ/H�a ڤ�Q�)��R��7���	�U�<�������QԦ�m�[էQOx�붜5q�B�\#Z����]�W3C[���:�0��4�E|��
t�MP��9��O�C���0����;��~��ߙe�p�KC�<�zn��N�*낁7�/D�%���g"�k6�u�c��H�iW��� �2��U�!v�!�[����ܯ�޺��;���B�Ŋ(�a�d	]yB	�5�����[�Y"��Y*�eu)oo��"������t:6=^���7BK�~�nRGe�]����:D:�uW9��S�*��S�֪������eu��ށhFM�y�z1�����y�"+/c�s�'�9�ol�GV(�ū,v��Xu�I&2�f�kn�4a���G���܇��j�oP�l��iN���3�Ʉ��7~���1b: \»�]�M��~�m"����W�|	����qk��yD0:�*u�/Y����=�W�-��?�f$NK�5a3��B���Cg��,4,{�e�g�Z7Mq\�3�V8�y��>p^��)O����T�
���mZ�B��Vm��N�Q�l=����c]&p�+;�)l�CM/�F=�a�Y�|��P�k�����᾿xo)s՗B���Ey; ��=$���X��WY�^9[r�k繌�yt�c�iб1NF����"�/�_Vc�T�'�^LM OT�d��6@�,'�o��|56�}Y���5�uYVM�M�4M�WB��<���9�o)�����3��)�c�����9���K���^�M�Lzg`$��W��Yp��%���a�/�{ZM��,^7l��� .�#A�ݐ
��S-��ؑP�.Z$�vuTC�n��ӻ7�!� �h�f2�ao�@|Ϋ����"U�1�1��^�F�*���W�Έ��U�0cۖ��`ٸUl�Wq>lj|��9d�KL�ƞ������]�zu��� �?�����>��a�+v�*5����os����4�ϼ�5OjHUyg��嬌B4#f�ќ���G��ȇpҶֽ�'B��b�ԓ��x�<"��f�����!��!��.ު��J�h��=�:V�w$Ǻ��K�"V�}T}�g�+ǝ`P��v�3���EdG�=f�R�+c6��g�*�W ���$6�(�@������yCu���f%�
J$�9�����w\�כ��u����Պ�cjCN��mt�/+3
��������Ï��gR���V:�w�g&��;��T{��;�Rs��4��R�׫�ڛu�D��k'�ٝ@���lW��,R��1��J|��*��M+e�{]�7v�!�.d��s�!��s�%�lwu'��������nE�p�n�l�U��mu:9:�Җ��u3!F2���M-�UeJU{Ր4pZ���R�[�c���ϚW:���9�+[�P'̨��Ky ��F�]��\J��1�G��!�/v��yWU���ʽu8#ovpZ����<�R;fU��a���3Wk�GB�	��aw�e����|�dحqc85=��G���8=$"c�lL�0��ޮr;k7/n����jaH���D��ˆ�Gδ�����3G/F�ʏo�6�Ev�a�I����W\��xJ륕�邚��u/��m���'h7/s�w'6�LT;����ݴ+Z�5K; /.��fVzy�x���/A��q�`1�WW0,���Y�(�*
<;&S�b�'~��x��[1���/����#m�Q�Ʌf�m3[�n�g-K#�4�N���)A������Sz�A�o1p��й�mJ�M��b� pWet�@P�$^d״�#�j����V�,"�Z5P��n��n�y��[T�R��ƛ��k*�t�����Џ�dN�b��k����g0N���%�tΪ�e!w��]�i&<8�l�B̚��= �X�\�bzIyv�[�P)P7b�x+b�r�tK�Wcr��?[��o�dvRt�vwE�P�>�,�2�eU�Noo�@q"��}֕�������![oZ��9ŧ�Z�/�����S-�,��sh�9q�+z��y��Ns��n�iI����CG^���:[ɚi�����:��ܽ�s�D4���(fݸ��m�掼���W3��)�
��2m��E��L�wv7{z���h���s�@�]mV����*FD0�v��:�зUn#m4Ӈw4�ŝGs����w}LWfo������
9^�YX1*�gu>m��\�EAm!]�qT�h�V"�_^_n��aͶ����<],���Wd��Ɣ���#7Ys.SB��.�i
 AX�Y����A�s
�nhʚ����w-g�l^c&�A���R.�������
�aǿC�"U�ku�7w��f��7E&:��Z�:ĭNm��	����v�S4u��NZ��-�6�?�<���c9���Gh���	~�3 ������`J��!����!+��!>�W�M[����s��&=�RKp컩�J���i0��CÛ��6M���9�1���d��J�u�5��[ި�J�u1sB�n=�&�( +��AB���
)h9��D��UIFa�`�^FUm�S�?�����׏<x��~�_��ބDv����v�s���Q9�EdQ���A�9��FG��1%%�0����q����Ǐ<}?���g�j.�̀��,�'s�H"��m�fD�s2��	�b3�*,�
��h�2x��:�����Ǐ_����fz��Q�"f(��&������I(�̊����~����0��AT}�j�j��=���*���(��G'&*l� ��"�c(�f7~��< �c�9L�EQESLTddQ0���IG0��"��L��*�m�TUU1QT�1A�dDm�1TG3"b�Q�t�a%���8�fErr��)���#�����(��Q3d߹��m�3)���0�&
��3�0���n`�[�4�9&�f�I���.�Be�UMfX���E��,�ͷc<���vv�����ɢ������b�Ә������h@D1Qfdr���R��9���մ1��Ɓݦ�I���p%'F]�"r�3]�8D٥�p8��8��;2�\Bn��횷�D�K7^����<�q�@������0��#6�3���]s�:�t��/�"Ŷc�4�%1u9���wb*V��E�b�b��>ހ��ņ$�k�@����M�]L�ʷ���m�5�9w�=� ˃�O�s�q��
;��i;�۝�=4D�T.<Ҥ_\�w'j=���#z0H�FC�f�F���ĻTV�:{p;3��W���5X�="��H��3�׹�H���(�]��3Z]5e�����[	s���|�"
3�7W�2�I��  {Jl��v˽�VF���b�r���i�m����e�ӡM=ٟGW��uk�ɪ;��E(�ѷ���]ӑ��#�����~���5[U������� �R�5!G����WK!�u��f�K?r#f��sg��+2��q�(-�vê̬��mlؾ�ޙ�꘴��W��-ѯWJF�S�Vk�h�ϖ�����n���C^�oD�B��Ļ�wF�Q�q��'�'{ɭ�X��������B�mS�8�jƑq�U�4G� n�LR��^Q3N�;��s���E����9B�Vhg��7�����v'��B`��f���w���;z��XF�?�����f����M#R��
[�Gi����ֹgߑg�c��~�^��1�Χ �y��Z]8kp#!d��_sD�]^c�}F)e�.�{j�E�%m�=��a�do���ۭ�O#z�р� G�S�Wt�"�І���c#�'�������~�%_H<	�C�y��)w��=���j�K���S�����S��8f�T���w*�OZ������`��C�Kꉻ:"i�����u�j ��6df��������	�a�ݴ��R2+_)m.M����!������= >,���I;�z掶a�<��q����V�
Kc�����yv�(o@�f}vme�����k���#�ݻq;���[�2�lXc�3*�EV*�����zo�ܛ�;����p��m�ԁ�ؙ�_<BQ��^����S�R��4��zj�әs� L_t|��>� o�V9���p�+{y]AA]쫵u���h�.]r�*^�yؠ��:C'��l�Oa.����C\yA����C���V�<	Y�QB�kл�����G�x��5�o�n�a2t��:xە�~�a6�,��L�U� T���MdY������,7΁��ĉ��XU3Y4ˆ,x��j4���SL*;�t��B��=�3Hf�
��!x	��\�!Q�w�t��e��P��Ϻ���99�ϨW[����wK��SV���[I\�qZ�w����E'7ۼ2�`�i�=�!;�cw�E��'�W�-���`������{�N��vn������h��B���Hr��<+���-г�{���z�k��^��8��Ш�8o+�kyQ�,�����W.�m�\)%�mx6�g��Y;U�{�˷�y[�S�U'J'�}}M�!.�#�U�4Cj{6��֣�ѹQ��V���R��-�Q�wbF���rC,��V5J�]��=��c�C;�峆^{������W��rT��}�b�:���S�R�z��0)sf�ښ�Z�}���:���i��-��eGwO���M����S#��L�h��}��U�V�)��W(S�+mV�`�fM툶䙘gA�h�5�])֕�[��^���I��w�Ѿ_P��������YG�[���ݸ��d{��u^�O!��;&�
�!ˡ�Z�6�`ǂ�`�oU�qs�r}��k/ !�{��-�kh9^����L���S��J�>��aWC�Nm�[p�RѹY�tB���ӱ���}��;6kff0!_�ˊ����{������u��f�����.s��Ւѐ�A�|Fq��<l�������Dݓ�1�.H*�mn�"_�/��eP��j����莑|.v�>���k뻮��o(��z0dMT���Ϭe�
���P/S:�b'Mpl��-F���&�j�J����-����p�iQ{���SO2".���wI��DM+4�z����o�7��e�U�����af���7x�*�4uu�d�Qu�jV�c=z�ռ
�����"������xg�ۨ��2ku�FOP��h+�7L��K]ǽ�p�nQ�;Zd*f�=ou'��^('���*r�(�qM�w#��4����xe����>fC�*�8���eu���-���e����[�b��H���\�^ڂ���8a&uŠ q�r[um��miP�t���}W4��V�����퇆��1(�:�"���v7F� z�[��C+��L:��x1�;��P��U�3S�E���?|Eg�Y�e�8酙���H��x..�����v�=�m��{H+�pGv�.(���wM0�Ĵ.��rx�QmN�5��Lc�ɻd:�YǗ/Ӂ��1�`ɷ��@�
�2;�j��(�qU�#j��n��h�r�A�y�'���FnZ3>��*�kk�z\��غ�'(;�;__b���B�I�oH}��吅/��3)M�s���7�A2�N��=��z.������?�y�y��������(�g>qJ���3y��[��L04A&�z��q�K^�G��3������i�e�+��Ķ^���Gyz��q�:���5�{6����	�,h5+�@�b��o��x̖�k:�lׁ
��ح�b���Oޝ~��ֳ���A�ory`�� ���T6�=�]���aXr�7�w{*�
��~H`��5�υG�o�]�N}|�B�֭M��-]���y��k�m]x��pmz*�x���8��Ó�;`.�T�g�Q�hY��,eO7\w{�A.3���6�PhX�ګj�K�Z�$�K�ɽ�VJ�e��t%.,�՛�&��]p�
�,����Fk�Ú���g�1�T���.7.�6ī'�{�^�=Ꮍ�vxܚՍj]�N��7*���oVL��*�m���f�\]3��Dv��l���挬�M��w~�Q���h��I��)�.ﶻM�D��3�]�����K)��x`�Id���۵Ef@i��^��y͝U��Y�M]:��Fz��H�:5�-R^'!VEK����[b��#����o�Y٣�/Coz<%ky�r���	hˆ��y=��;�[}���m�9-�
Y΋��{1.�}6)�0%o3�=�O[��m��Y�x�ۜC�����U��m��,��3��4
��r��P��m��	��y��x���_�8����2Rs��'�i��윊��K�5M�?G>�t0��r����ڢ�j�`�=���g~��ۨ_�ǳ�gaM�p�C"�����N���}�[)���u���.�ւ��E���e��ΰg	5g"7yb�c�fDȐ�
�=5
Z=�u!lX|^ʶ�!ɹ�����s���H���O3w;��ʒ�Y+&h��%�|����ݧ�IR
��E4� ��R���ifs�6d���vp��A�Ϟ[N�v��#9�yd���v��N')�!�0���5:�<�׶�����'�����pګv�M�^�Ü˵t����vkޑ�O�GD����g�C׍z#���&�X0�]�z�j�����ٸ���vӢᏰS�%�ֻZ���ܦy�W�����xx.{h�<G)H�涙�N�Y%[4{�z�j���wDb�>���5�8��ӿz��DF����X�|��&/=I�ԣl�qRp3�ӫu�G� �J����7W�F���z�q�X���+%�sE�hܛܮ����B�|�i2B��O4z�.J��uSږ׎I�&��ƖU�]Y��,� K�o8f�p�Q[���=���m.8�ϟ�pu]�{�V�6�Ѭg���Y7ۻ}����][��"N�M;ě0��,�<;,�yV�}{O���5=l5���tT�g����]Pn�]x�v���D�\���0ҳ]��H�ە�����8��'�t�6 ���
;������5$��Z0�S����-���\i�X;�ES�T�X����ܤ�i眚�L㧂�;���ܚ�y 6�&��ݴrtM�m���[��D���A�-��nǧ���ii�Q�(�������nR������P,�<�/Y�T�̝�0���"�h��]�5ԕ+��>Qp&�Ɇ������S���f�t0�j��!q���3�V_k.wn��sc�'p�ŋ�f��nO
S�΀�]�~`Q� Mj7��3
�X�j���6KGS�i{[�kl���t���M���}W���Z������ t��{��7�`�.�w��<n3m��� �n�`8��Ȍ��!�1J��-���&~��	t%G�?��7����P_���U�<]}6Ǵ@;�\;��������V��5��Y�}�bq<Y����/VN�B�U=L�\�l�<Lޞɻ9�n�5��N�k�|HLMm׮�,�͒�!�=���y  ��d�2�y>b�ivR��K�P��ٺ��,���4����+i���Q��Y~֦���Hq7O�{����|�����Q+�s���>jd�;os��wEv�@ӝl��b��`�J�We��
}������&��e̮�o��I���>*��^&ش��@b�|�jDt��ԕ
����;��Ceme���W��������*���B�!˥�@EG��ݟ�lCk�+�ú$�����#ׅ�tV� ��9l�^2�wB��ym]o��bn��w�S8�q���5z�Ѕ�vm��+61VM+��or+}�d����?<����R����˥�|�eVψ���2��riGF�+�K� K3y?g��N���M:��e��_s����,:�m�D��]�t�Bµ{��Iʢ�d��Ẻc���Y�qG��Ϛ���q�����[]��V?mI�Fj.^�˙�U�_�r��wq��a�Y�1�֌�t��^*�Z󕇵^�wU��-�g1f���Vψ͇�o_��A�7��#���jMi�jQ��Ze�h�*s�e�SFZv@�6���=wj��C=3��E\���Ftk.bV�Z�^{� �kƚ{B���� v���6Vqkk�:Ek>.��XQ�絃����9�[�:�\d�T����!�φ�����v�3��ҧ  yo^Hy!X����S׮�>9p�f���}U1�ӫ�f�P'�}s��p�w��f��y��x�>�v÷q�=�B��z݁�s�li�#��6�"�}�y�F������׳ݶ7���m�ڱaO�������h 6i���D���.��4��qh��c��5��h�n����f��m��p��rb"�xEҳ��Sym��KzI����Ƣ����"�3G�S)-�C�G����[鞊���z�c�|[V��1��'�Ng���y-�R������x�k�{�nUXRz�ɦ���ެ=�fŨ��@���S���=+mY�U�ݦf��,R��b��S�Fn����Tq�+�s�<\
Xg_���R�(��E�&�lӫ�}78�k.��c*mذ�+��V��
�7�!���%I��r.{1�a�f�1�k���+���#�z�C[�*���]��ڗ!��|t~a����oi,[(z���b�>
�h)��:9�J�b]sw��Nჩ�ut��ޝ�y~��*>�`�-&70�!�1�Nv���O	�ٴ��˕^��ٔ�1Ox�Т�҆TT�����u�Z9�aܪ,��7C|[S�h��X*���%oz*��Ρ�(9�Ӭ���)ds��� S;C{�!�L9U���+SW[1�v|�0OEAfM�J�ҫ�< w$oك�Mmu��x�U�"��k��xF��Bm�7/�"S�*wB�^d��7�NR�ۥ%m�J��.�[a��֍(��$��V� \�[X�>@*��՘oK�
��40Ԯg`��c��d�Һr��zF%ር�+�����i�Z%
ǜ�ֵK*	E�e��SؗZ\����:�p\����{��{dAY�iw��Q���^lZ�}¹�Aq��]�x�ʝDW,K��/���Cj�ed�1����ث�Uvv�>�K+2[��"N�v�����
ISF�ğѡtg^�;H��Ӂ屏6��{��'Gg��(o&�k_�Ûݲ�E�ݩ�+���cn�-�}'O�:Ҡ�]��ZOH�^S���'�9쭜�j��<$i���S+.�S��P]����|�hf�[C;�VWS�YՍ��+������ԴՆwo'����(U��	9e:�١���Q"�#V�ٹv�cO����ۦ>�7�u�R�z�d)�~���a��.�R�i��qX|�mK�F���7n��2<����!��m���"�a�)n�͠ ���d�H+�i��b��{����i�ᓳ�}��7�/��z��k��~x���n`���=l.t�;*<��K���P*���9Q�֞ɻV{�J����s�:�pݾ�ɼi����Mկ4��{|��_�'\���oe5&�^�\c����Ge���C��q_rY\� ��1�A��k�X[L������F����3Vm��R��;Y���*v�D�m*�V������{���1Tm]b{����vjT� �l��ɧi,���{ 㭋7��0*K9٧�Z��c��K7��9�u�S��3k�e �=���L)�4+d�
Wcˢ��Ϟ�nf>�tn[VLn<� ��mw�[�V������{'y�v�A�����Q�P`6��{��
��p�Z���U�|-l�a�)v��1���K�4�A!���֚?���9fr��,�a����AFM>�	WFA4_v�"2����t���M�mGx��I1k��Vz֚|x+�� �ڗ]4d�x���h����.�5LϷ�F��L��8Y����&����,3"��u�K�>��3�j��YI
��Ê^��;�Pw�-3J-����11+%ږ�ì�h;�9�)�@[���,ǝq
5��E0CE��U  ����A�E�AQ� �nP.��d%�L��ʓ4qR
n�m��r8�f0�@�(H]���ܷ����G7r�|��[�n5�����9�a�?�ޛߦ�_����C�Ę�c��I�t�h*�+�͓kp��#����&�ӄ�u����Ǐ>��G��f{��~�?n��7q��K�A���f�T�da[��FITTTS�cAr�M��㯏��<x�~?�����a���EM~�70�ʫ��Q�˖�����AldTI�a���^>?�<x�������g��.�c�V_�2�(70�ܳ#��~�7&9��cG��a�J��2M��'���dd�NF0DP�LBLT����APL�f1Rm�D�eIf8LE5y��QTLRL��C��$��eY\�J����L�(6�(��7C(&�)9S�ѐ��TMd�Yr��c13� *J�l2|�e�����(
j��̥ȭ�������rȒF0�n9Qrq���`S����d��eDiPD!E1da%Q\�/gl��)(XYi���c���I��-�y�:��Swv�;���)�K�;9�0�,*\��Y����Ry9Z��nĐCYje,�qFelܝ�Vm�[�ɵm:Ȯ� �P6�4 "�& 3!FiiD����[..�D&@�5|��<�+'�RY�!�r���w1.�}6>��!��ON[%�oF�YP���.���O�tte�%_V��x��Ǚa����5�E���!�+��3lD�l��`aYW�,:�W�	^�v��>�ɺyELN���x���<A�{�!��hw��3���3��v��qi'8)V�CPʛ�Z�o�F�Wo�u��Z./�r�6�w��
�
��]�Ems�����m=x�t��j9!���&᷺Db2 ,3v`ZȷÚ��Y�=;WgS���H螖����8fmŸd��c�U�$�����#+�o�z���̯6%�8�⨿��f�H���2��'�"d��Z�vOt��׮����GڽۭmrC�o�� �����?/��f��vd=//ES*���_a˾Z����ʟZȹX�7����/Oˠh�׋�ԥl���R2�_�[�ϱA��ht�7��,�u���3�6�h�j��"��}�X>=�H}������Ț�����7�]j��cs�R� n�W%3��m�뒁tW)�ҋlOwYʽ�x�M6��1���y�eTd�@xN�q�i�ը>8nɐ���t"Xj�
�y5y���f%Pa����i�U�צ���<jn�w�sĮQv��[��Pt���ǃ��ua�9�NF��(��N��ٔ�}@�Y\(J�sl
�mK�KS�(�fw�����������3X(�b�v݃�"����-)�*�:r�����ȟLy�\n/m�t�a��ॐ%ue��[����^�貹��Ucn�)����H���k�P7eo_9Hڃ�A�����kXr��CsW<���:��L2.6����i����:zgd��UVD�,��Me��,��\2�G�ɀ8o2F��ՙ�Zr���C3�g�h�[A��u3�"�N�=dN_{5�Hf���3��G!iff�1Z[=����ՙ7ۜنb�;U�<ޖ�5�M6�x�Z�p5ش	�W,f���D���[a/̶;r�K��e�i���DR2x⚠�˃��V��$S��yn���7+�G��,����T$
)�X9R�3%ئ;�]¦�����Lc�4��.�N�J��U>�Rvv��e�ͥ:e���uK���ͦX���s{�h�7(���oݦg{N�����X^2O�]l�Ŀj��[u�F�P�Z�U�7n����s�oBNڬ���Am�}^�����ۙ��o{��5���m���V�j��{P}lx��-13o5��K�>�������)����ش��^B�1�fة��\�[75����ݘ;��"�X��[��g��y��f�GL��J�Y��Ϋ�h�� �{jhlqmv�5�qonH�n�wW�>3��n��]�G�HK�3�=yg���6x����N���rF-�jR�W�]�����s>�j��7u	7�ރm~��%�ze�A�Xnn��t��J��1|��n���h�w�N�?[��x)���&��� �k�¹6#��en��5#zj����\��ۦ�kC�/!�A�r��k�K0F�h��䧺��'觉n35�ùCiP�}�kx.�L]>��YI�`��͸��c��&DuÀG1k�$7�w>�]7��=�zϖn���
��7��Y�9��׍:��U��<��ċK7
���K0�[�ړKf$�Ŷ�B���Z�ūn�i��y0@x>Np�����7=ye�����u�#V�d�#gK��\/<5Es�s�9i=Ŏ��+ӭo� 2��R�w��'��:�!GNu�t����r��˜�Y�>�~�����Y���]>f��p���6��sͭ�:�g.�5S�n�C��A<�DG	w�q���w{�Y�-���d���Z\�X�C�>7Yy�bm7��a�ta��k:k��Q�� �צձs;�[``�M=�w�>�9���!��
̋����o�����og�)*|@�M�������[�ټ�sa�3{�d7�Zp�S�l��2F񮦵mtF�7Vsh�]Uv5�֚����`�:hN�~�>*�/�]�G��̴��փQ1�~ ���C4qR7S�v�m�x|�{
�9�߶ᙉz�r�G·�̎�4����\���=�T�QdjƋ�pbg�R��{��E������md�B���Y׻Ҁ�/W%,-���q���4=��^}��~d*D8(	aij��g�Ff��<'��I<ݘ� ��iT�`�
;l*Kow�o&2��o:-cn�z�ͺ�oU^Mc��x�0ڱ.]yE�閖,�GI���Vr�q��'_f���k���0>d�������ݲ.s8a���c���3��߾wF��oG:�3��WŔ��@ȣ@o,�YL��趸̸�����]���Y����ib�ˤ���f5�4��H�iEu
|vӯv/h�I9s�k2'�x�PZ���P�tKlrT�^6���'o��S��\�Z���Ә��n�7�W�Y��p���t��W���]�c�us��iv���'���͆`np^9+�wo*v�,���f ��}}��q\�:�b���uqͺak�{8�T/�9"����d�"3�	��]sr�������}�''�o<�񊆒���+����X����c6|������T1,��
�i��s�cZ�2E6��w��ۈ�@���u���˔�Y�M��͜��r�F���)^�v��+�M	f�e w��[�'�F#"�6}��v�t��t���a^_,��Ľ�����me�`3��EZoI�3}�g]�6��C��m��t
�4��|x�n���=媱��E�=���I���������=���yw\.ԻIؑW+#�}c��Z�;)����}Av�0��׿=<{����Z��pɝ�t�9͸�shkg1��;j{�cEB6c(�ԻI �E���6)}��������Y3�o7[{n�K�WU�v���O��H�'+���
#�����gMu��S
E�����=�O�CJ��g&�]?��O�w��{�XT2=�:F+e��"2gh��O�d3�!T����mS!�j�@�i����ϯ0VelЖ�n�(�q��1{ə����r��Sv�7D�������g-���1ZN��K3k�nt�򬢳*�X��[ 1ƚ��\"b���Ktf*錻Y�Ƿ�\��)wY��6�������Uڽ��Z��e��r�ͮ���+|$^��أ���o�d	]YQ֢{�9�"�ܩ��:�Ȏ�ٮ!��L��\�݅���)�~q#s�|�%��0���O?C^����׶����v�6�\1��~�mn���lMJ����V7��L�6r��ȭ��ׁX��}�ˋ����6os�s�8�>�fq�Q��v��ZF��i �qs�oC}рɱ>�R�k��Up�� �]m��p�\1�5x6�C�;�и�����j�z�0���@���{�ܳ}������a��}�@�H�k�{">ޘ��1�5����c��>H9g&jv�j��V�h�+$`�p;����{Q�QnZ�E�`�|���
�G�=u��[d�o�Nǉ��w�G0=�7�CCq?ǿc�\9�s}=�3� �p�'�a���`ӑ��5�M��%��wc1����T���e�N�5��������+�
F��G<M�V���l�u0�2��+s۸�G�Nns^��D�TU3��� �$l�"�mLs��:n��/�������\��	ߧ�,��z�"f���y�_M��U�u����3f��d�X�0����hF�=��X����{�-/��*��)���dӛ}��)�#��+�I57@�*��<xt����[�s����^�y��~��}�p�(���5��m%�Z[�ȣ�ɖ�@�? )�7s��k<�!�G�ꅥW�D������m���KTicv<�K�r�`�-�δK���{5L+lu�Q�J�{ωˮF�1�n�\�5�6c��L� <*�]�7U��?>L夺�Svz��6AWk׻�2��= 5�a��m�֝����#s��Y�:חs��k/�y'�8!VR�����ɘ���Ȇ�y��f嚙����&���l��=�(
�v]�c���,� �]3d7:m����A{���W�
��H�w��B��-���<c�KNɦ�
I΍�ks;����AO�j_��W�V��H��&�qӷ{y75sV��媻
�JLL�V�;ne�D?@w��5!�Y�d���k\2�$���x\w��e�+���1�V���vff`8���5]W��ĺ��:_g���V����F��<�>�%���۝����=q���&؆�SmM�S��q�����dɌz<�[Ծ����4��d�dW��`�Vf�v��8tvx.�����A�Ԃ�^����*G`����׸�-�Հ������0pm���"���d5mY�c��̹)�)��+I���f:���*���OPJ_���vIm��l�q�9��d=�{ϘH�b��ś��˻E�G ���a<��4}[�jՀt��JM�H���1E4�U�	�Y��ټ�z�Z����W�d�t��v�!�!�x�ȋ��'�8�uӳn���=[����g��3��@i0��;f�{����"�&��5QO
�1�Z��-pQ4f+1@�6x����q�4P-����x���!�s*�߲���_r����@��<�o���|j:F+k2�AKQXgJ���g"^�V�14�5�6�K���b��'U;��	��
̥ݰ(�S='=q�{�g H=T[%ZQXo_����R���x�Ɇ��V�l�;^�Mگwc�z���f�b[���T������h�S[Z��}�S��G0)���f�c��Y����+/�Ճ���-:�7
UWX��`�-L��j����֊Y�w$s��<��_��d�]��S�Uy�[�N�jIs9ʯ�u~��υWF\�o�ǃw�Ӯ�����8c>�nu�P��+i�;�J}���0j������X�9��}D�;��%n�3��,�,(;�֫�(%�5)�^�:���z�:�h4�tvn��W^gNX��t�(d��
��6�,)Ӧ>���\su�YjX�~�����g�A��@CҟDa�b���CJΡ���V���A���/=V��9��;3���/^�^u�}�Й���Hī7O%�=��wae�����ScǺ�Vy��.|�Fٛ�0��W�Q1s}�k:�� �$�wHn���-�#�#��ZU�[L�%H�y���؆;ͫ6��L��������|��m��w�]9�2"��a����K�#n7��[D�U����lR�%�<�ǺuQ�lñ�v�x[s���<WeZ0�8��<����Y%[o�I��>���{M0��o�1X'��vU6�z@���U�e�p/#�K��C;B{!���2�dT�u��UȌ�I+g�k7�dfC�Tz��JJ���V_(�cUCNm�SL�ol��$�ܵ`)�H{�cP��!r�-o}���W�J�O�:VB�ח)����j��c���ڏr��k(h�a�t�N�/kc���b�^��WfWd���	�'ϳ�
@۹b��m	�x㩶1�������ȴ*�[>FS휡+�U��fk�b')�=/0)t��1�	T��傮w��ͫ�ߣ�w�8(]�RS��7�4��[Y�]���/�h�L��m'�(��ج�so����R��즓�8U���ض֬ҕ�W��̤�rbS�o7�"��7Wv�r長M���u���f\������b��ٶ3&e-�fJ?^�t�1h�RΥ�V4��*G*��-�V�`tbs4�1�Y'7d��q����cI��	VW_Ps��J���i��p�m�XηqMަ�n��x�[��1QQ�*�?b�9���v!��HkG�g�n��
Å����P�����]G�������!Rw�G���S�V���{�3����	���#4[=�$Mv�j|�^���O��wX</b�/@�v.]ќ�}a�z�\���mخS�m�!�u��g���.�+�L�c�jejm�ۉڛ��jQ;�Ly�[�\P�f�C*Q�%_|��MCC�}�Q�M��s�C�B���mG��0�;�"Y������W����&{���}���[��w�����闑�E�Һ�vꮹ��qU��{�_����}��yg
��6?F��w�������s�p�~���W����06���b����Dv�s���HG�7��LK"VfnH����fn8W]�%NG�U%����G����\���aH���wabe
��+���E����3�2EZ�ծ��0�0�&LĨ([Vs�@�o5[)�]����K�d�BV���wz&f>��FDxkw�+:襘6��uL�m�������u�L��I�Wv_;r$F������o��oF,E.�Qg,��D���g�1�p��F��:5tT�B�����h��}3����gC������6h�H�R.�r#�w��x��㊲GJ/���w*��� Y�_oZ�4T��G+����|��P�Cͻ�nZ�C�0�ٗ�͡���asb�^쏪�[�l��O��<{'$��W\WM#rk����c�+FQ|��A�eg�Cr!ot�kLS�%��Z7��+��X��x��=�����έ�K��"�lf-A�}qH�@ov�X�w��tҵ�僓]c�؍څo`H�J��N���؅�U�6tH1�Ԫ��f#����2e�4yW�U�f�S,�Ƨ��&�a�h.����{���9��a�<�U�q�<�%�w�;1�I���Lǟ�&N�z.h�o7Sf�yV�B�N��ӏ>m���@o/;��yϟ}�rr�m�@STDLEI�E{�6�HFca����a-9��<z���Ǐ=~=q����vj$?gw*J60���QI���*H��ncAAC׃��>?�<x�����q������I�0�h�8V`�~�������8nl��1Q� ���}|<x�������=�{��AQP�G�,9`QT�IER�n9�'��ʂ���g|�7�͏$�Pnfnd��n�YM�ULU%,��\�6
4�Y������Fß���c�6����D:��L���T����-������]�a���
i<���71l�1.�@Qfa%!f&In!�UKe�JV��@PӐ�&JdQF@aSCFdCUMg0v��"��)��NI�d13��9�0ܲ�	��C���{<ᔱ���62�-���EFI�d��VXHV�!�{��R
S��I���=��Xܬz�=�i�s���ۋ��z:�i�Ѿ?.�١��\�rZl�ô���{h��z��q���h��g�����w�0�IW�IcaW�m�x�=�Y��Z����{����X��&9��5¿&�%>]�f��� �{9������]49��Ogks�mɬ�����޸^�b#x�l��QՕ��Qe�ND3M��6�z���z�p�7
w4z���QM��7P�sV��.��7o�� �s�?�޲$�s�����zD.3q��JexY�Vkȝ�y�z0�x\��V^��DP�9���0;z�8�oTAF�8`^�����x�ݤ��Qӹ�iJH�Mۢz�X����Z�����=$�EncK�e�n�j�AɆ�gf�9�j��� �{d���Oe���o�|�iP�.�˷��o[��!����ǃf��3����^�����*�BH�����_�sS�r8���X���޲����9����JUߧY�q��Y[���&��F����cK�����W׵+52�$�丧�t�ᙷ��c�7X~g:�(B-VjYS�����c�]��ݶ{������QtY�W}�wD�&gY�O�e��+�(�[�/DQ֋�w�S�W���r�{�Mܘs~�%���ފr�D�*0��x��Qv1��#�P����%cPpp��>��3i�K��Y���*��ث���\�e^,0M�ǘ�k?u���Qs�ّ��f\�1U!�Ԉ�u+V�,��OF*;5�y��ޔ�����ts�X5<v��֨�a>�m�zq���;k|�.|�}S�o37o������ʯ1�N$w���5x��Ps�ʆ�:f�}�*�^�4�M���/MR���d0'#��Xdm�N�Y�-Db��>�;A��+�/��y�'&����j��yk�P�e�,b���z��R;Wp�yX�+H�}ƪ�ھ�a=d1��~w�+ڷ{g��K4���vZz�����tDt*��uئ2�/=�Ov�6�У��]>nxu��{FAh��/9>�����r�����"�E�u��u����\� ��܄IZP�y��.��
*
Z��\L�m���ެ�+�(���}=+W���T��L�\��v7�u��T� ��TL4@_�dغ�V���L��v�뾑\g8�ݵB������M�[+c�N�N�r���'X��=.�g-��b]���7�Oz�s{.ր�m#E� H��1H�U}E���B����� ]3���ai�q�gY�ֳ̫݄T�3���.��?�.%�������نng`]؊����3���;�;�������tw�dJ�ۋv��6�Eɀ���gA-��ss����\7V�f{���F�	��u�9��{3Y�}�������5�5霳a(7��^��q}ʂ�GH�9f��Y 2/��R�͋�=L��4UL�����;^��S]��W��l �b��:0+�����3��&&���S_�f.1Ih�E@�������>z��@q��WZc�7z�˾Ɗ�jj�Sd'�+ V��;��bȡ�F�����_V���@��������ͺ�YW�-B���I�k���I�S�R��ؽ��v9����3��� 5T2����i�6Җ�L����fg7c9GW�g@�Ѧ��6T����O-�nc�80�J���Qp}�)���c�~����O���n��T�k�]��Ⱦ뱉t�g	�x��ë%�|J�R��i$��v�ө����u]|3�)
�F+������U�kzW�����,Υ�7RUlp�iR�?%�3��[�WmQ�}��ȿ�:E�`v����?g�R�U���پ��s��1O��dvUJ�-o�j�;��Nʔ��Ovy��\�$�;�,�E�����dq.���F��7<�D`1�z��P����_��!>q·�+"٣�U��%�5������K�Sy
o�H���.|�A�'��Eo'U⻖'�\8�M��l�wt�o]&<���>�fDF���ӉVz�����,˧8<Ig�|����d�w�`������p�������Z@e����eOf�65�g���<enn����#L+����t;�6�{�`!���1DF+js��uq���ެ���7�Ix6�A��63<ɻv�**갶:��N{M��$�?�^�l�g�ۍ��[8�x_��i�E쳨y�fm훙���U��-8�˛Y�q��)�t��h�9��-QW��G�<��q�]�P�p�]`����<֖tJ����\[�㦈郯T遺���yu�a��0����1�m��<(
�e����&��{��%�Fo���4�����^�=7loHU���ᙃ��X�)h���0�"����V�#t�p�pZ���>���U��e�5�Exe�PȻ��{���d���q� a�W��}t��,r�����*i%Bi�q�,4��}�.k4RCT��K+U��g�L���`��x�� |�~۬�����7�]{aH;@��Ox�K�	;@읫�Y@��J�2�H�%��I�uiͻ՜]�������m�S��s��ė�5&�,Ȑwj���'Iʣ��baV�RA�ݾ�-,����y[�
ȕՅ�y�t<�{v���A�ʛ��)��EL��P�u
����ݕ�~�+��Q��mMK������՞�^'�C��l�f�\���7l����s��c;��Lxe<S�wgv�Ѐ�Bs���^S�oK�E�=
�g��5��uhfm���2F��H�Ѷ�xW�ۡ�P�i,���.�P�7�uz\���}d���X�&�A�Śgd�b�e�T��]Ci�ٚ7���߳����Į�����)�z�Vq�U�x��l�W|e*���T=GF�Z��f��;���������sPv(��<<��d.f��nm�'���EJ ʀzcy+�ݧ(Y-�gc��t��Ì0�z#��@� j����s�����fEO�WTw@j9#4�����3�5�6'���;Ig���sv�?���� K�'us�c�+�@����ߣO�4�&��tm�]7��fi~�e���ŵ[�x�j��k/�7�=a�8�l��Q��U>�V8�=��7S�h�'�υ��u��=���<��|��ZV"k��qJ�u��n�Pp���+̍.׭C i2hjƯ<�m�!�g؇~������|��l�c���a����K�ۓ���W����U�V�-���o��6�^o���v��@>�H�آ�1�*�YG��]j�e VeQ�em�z�z���]c�5��}��y��C�Xg��~݄�N�N)���
]Ĺg���P6�����>����yrǧ�u�A��x�B�k˰��Q�܋5�I96�{ْ�Ìm�u��H����$[Uw�P���!�*�1E�?���=�t8=�r�1�YD��.��{BoN��]�&�nU�\�k����:m�U��v����V�:(P)�>��2��{�]���4كӬ��Ê߆ȑVʥ���gυ<��\Z����'����ۈ���)��Yӝ�\m����Ҷ��sU�1�[,M0+:��d^��%�C"*�Wi�7��&�m U%�f���8�s������A�oiv�)�쭻w��8�f������8�����?t�U��a�[�M�eZ+wX<E��͎}�r�zjWE_*��ɶY��Ֆ8��!����3������<Ra|n#6b<�q*���dN��r��^\��koq/��X��k� �4�r��r����2;��4uM�٨��-g��ˊ�}h=./$1�Z���3�c��3Y����k���u6��;3}��`��B�/;Օ�|�ո'o��Cg���/�<=�Z�E���`���Bz�n�Dp^�^I�nj�i��#֩4�E� ?�a�ڣL����9��8�ݽ�K�y P����)eH-��-wu~ў�A �Ud̲�c@�k<��L����-��bB8N=C�����]f���G�_x/)c)^�\��t�%��;���7�6f-�j�+�j�X'V��#�w�I��
�	��Z�MA}�R](�{�C�xT��擛}��{s32����R+�w��\T�F�ge���P�U5�0���+uuṈ���6gm	HT��i�!F�[ʢ�[t@�-w��\8F�6;�6�d�@��<j�Ӫ�nM�^�6]��<�"����^������5#����joT7U����W�X�k��f`���'
q�۽{��}����7$ݪ+2$^2�g��\��p�t�;D�:�͵==�;�-�G?YER�Њ�6��zy�к��q����L�z�ޭ�6�E;�wv�\�z���<��q~`O=*<�U�y�.�!�ht
W:��fΈ��:1P�:CJӗĸ�<�	����� �z���أ�{{��^C놭.ڮ �P�D���o'U⻭@��u�+�:�ݯ��lA�96�M�u�E�V���1.�=�p�����
�6���
*�X1gaB;�Gw�}����тE�2Vt!�Y���W�ٗ璎�Bx���RC=Le�ߩ�+�#c�2�6y�gI��$�}��^��v���wל�r�L��V7�gW"�k��b���:��-�W�z$W�������h�v�:�~@Mh�$*z��y�Ja�1�T��Ml4u��֎�P�G��v�Oct��wPn��8,���Z���}�=��O�a�����}y�1��������l,�lɧ}���T���`��ùӼ��-���^�>�n3�H��O��)��;n�[s���>�޲i�HzG=����v�"��1��1�YA�!���g�]��7����&���J�����d#�o��|r��Fx��Wߎ
 <�o�[�����<�r��Aj�ȣ�"�Us���|���KY��SĈ��N��\��lx���ďiq9�H�Y��o�_����
�-C��D�v66��Q�`�goT����:�jZn	���Y�]�sP�a���/\�7ۚ)�p�I�1�����|'�p�K�\���pQqko�n�����ѱ4�_k=�|�w�w��)�WU���vP���n��A�������Z>��*��s�\R�r0�j����+<p͆
��9t�QG�_HF���+v��]Ϛ��/�y��3@%^�t2��u�������g�2�y�l�(1�]��|k���ܻ=���~+2�9�{&rLV�����A�����d� ���ީ���γWT���5[m����\Glj�mF�_^�Z��/)�uí���lRS���y��ph˦��z���H2vx�ߏgB�N!S>8���ݛ0�'�b�dF흅�7��wA�l�Yc��I̾��"�}|<���_A�eI�x�t����wVW�e���J����y�L�R�:���:���j�y�6�Q�7c���W�^Xq-[4�T;_ͦ�v��a��;�w������'*;���$46\�����0��B�.��ͦ�4ٔ]B�yff =a��]�_��z}�i�&Y�nB&}|�F=S{�{�SלS�̥ۛ$v=�#�{FI�b8Ѝ�g��<�<�L���b���wv��ٽq��(�*�Ԫ(����PC�  9�&��z8��j�Xh��}�ta��BU!T�%R�B!�!R�IA�)�d!`Bf�a�� @�BA� bE�B�P!	dpBE � P�u�BQ �%`pB � B �$B � B @�h!� � �B � �J ��B k*�(!"�B��!����J���J��J��(B�������B�!(�B�
J ��@ ��J ��"JH�4�B	B$!��0�B$!��h�J�!
���@�0	H�2�!
H&b!�$! �42	J�!��CC!���B����"B)H�
B��$!"�0	J�3�}+G�q�C	��@QY D�U��1�3���1���:g�������=a����I󦃊R�>�/Ն~=@��Xu��Ӛ*����D@c ���@�N~��N�;�_�����7�M!˽,/�}ĵ�S�Hp�BJn0T�% RX� �I%� !R%�HYD� `!�I�I��IID��I FD$%BF"!eB�I�T�$R@�H!RV$ed�	 �HB I$�ID% �	XD�A�!X�d$ZA��!	��hFT(�FY���HL�@(@�D�@"BeZ)���  $B R	��B$Q�aB$B��D&D!��H�
D!�	�H�`H@�P�$�D�w �(>���� ��2��
"����3P���;u�	7Vм�i��MB���ʁ���_�)~"vU>	Gx�w~Iy�s� U�!�8�nޘ�W`" ����� ��Hd7`E U���@�^%F���
�)�T�75�v��� U�����b" ��1I �~f�;M�}�0k�4�M_}��
 
�-�:�� 
�����v(T$L���!��d��9�x���-`��ʢ 
�sF�~|�z"u ]�����K�kL�Wh����o`P55�QE�׋�U_~\B�(���
�2�� ��X�� ���9�>�
��/�
����U)	URQ"�R�IT �H*��E�$*�R�UJJ�TI"�!I
)EIU�T�IE^��
PI)) �TQ)	$*U%J)PAEJ*��ER�IUU"�)HTEDH]���T�
� �(��
�D
*(���Q%Q�U$�($�*)@�T� BT*@IEAD�T)	"(*�u����%+  	��he�i�����5m��Z�6ūi�մ4l[L���[�e�յ[Y5Y�����[jR���J�E��B�J"	TEE*�  ��@(P�
��B�
P�w�(P�CB�	�8�wcV�,���1�3mE,�0� (5)�iPP�SK6�A�mF5B�P�QJ��J�)B�I� ˔�Q��mcB���+*
���+T�5�L�ղ�	�1�"��*l
m�Q3V�f�B�e��[a���[����B��(�U*p  c�kJ2�ڕ�ʪJ-�(�0�i����Fڪ����[a�
 ��b��5�E6���F����
UJJ���!)8  :�(P�R� �ke�����U(�+0�BSJ�	UYM�ƀcF�XY �Um�Pc5)����J)P@��  � ��k5��-U$�SU���D�`�2Ҫ`�BUVT�`40��kB�Pb�mI(�*QD����p  ��QU
  �  �L� 
Y  �4 �`
h6K  �څ  ,�  ��J��U
�KLUJ�  k�  C`  6T�5@Ԭ  d`  ��P ʰ  -Q�h
4�L  �L  EJ$�*�	J*��  &�  6*�
�jV� nm  1V  ��@
6  ��@ɀ���  `ҪU*�T%H��  �� 4b�  c  ��  Kk  j�  �0  U� d @�5�@ �>"��JR� 4 �{FRT��d d��	�&i��~%*I�� "�FS   I���5  1+f��H!'�f.z �̖1 50D'(ć�����v��-JڱC�}U_W��$�3���B�u I$���@!I?t���B�$�@�@ Byߜ����?�z:޷s���Z�ѳ�1�Ɏ�z�-=0:I\@��r+"\����N��Vv����M���Ж�-]�W�t�"4e��4�K)j{m$^��j%���u�Y�'�BIF☂b�wSVü�� лaK�r���6'w[�Ua�ML�������  8ZVJ�A�������a&xX�;�F]�Ǯ̩sƢ����h�7�]��,&��6oiQe�lË\a$M�♢�i`"��jc��3�����ϕ��V�,�-K�7
8�-y����>nQ1 H�	7`eI�m6��W�q�bii��ך*�ʊ��ҸC��ad �$��5Y��ћ�@`O1ИCtC'�[
�Ɗ:ԃǲӢ���p�e�pLZ�ϋ:%It���o]G|�Wj�N���V�P�VH��]f�ۼSM3v�dp�:	,�&J���ʐ�j�$�9����!�c`�r��קe^��3j^c̺�Tec�P5i�vL�^�I�Ȯ����0�(�
B!�[`X�8^V�Z����ƴe�0dq�[zF�b�,��+th�p�\����3H�MZ��D8ɏC�t��X��H-���6���Hdx��j
1�4���x|ÙW9�4�H�Ne�+Eb[�B��kw��4���+v���6��Ȕɲ�L�j'��z��T���0)�[kKׇW�]�+f�ĵ��g`�1�	6PGuݷ���=*j���r]�s 57�㝩� �<�۵�ѭ����V�&�P�gi^0f$�1�g��EY5�QH�3pQ2JP�3 �u�c���u�۫��b[L�t��EE[��:;ZST UjiY�4���mh�&	t� ͋.�� y�+7Q�3Kw�m�7�1��a0b�����xv�%7j���`Z�[��<;�f�"�20��WM��PLU��X�HݭG,f�Z�Ō�#�F�K˧�U޲��I�aW�!����s5��kĊ��Q]j�I!f��F�����˂�ё�,e`��߭f<�7�ʐ�d�mdh�ܡ��3G
�eMVB��j�5J�aR!��ݤ4D��D��j�ێ)Q��Wm��L���ô&�)����,8C��N�r�Z��ئ����3 )���&�3KK6�af��.D-!�v`ȱ�(����n��ds2�ʹQ7p�Y��I���@`y�qC�9#�~��a��F��i!Z`B��[u�v-:�J!��j�ú�^t��t&�A��.�ڶ[�%nC�L+�J�k���{mb�����Bzk*D��'L�c��蜗q���§F�ɒ�-��K:��\9m���?�fC��b�wb4qX�Y��b��aV�ߵ��e��p�$܉��ڹq9/f��mw�6�3Y���0�6����-j�����:�CI�VJ�f,�@��o)?�f+@h�֫K~6ʨ�[ܥ��oC���Ի�@�JZ�ˀ�wOvޅ�+I�v� �sD��.J��4���F0]�шf�&hLK:l!s�v��LaZ%��$e�V!���sj���Xvd��ǀ�$T����72n֪d��NЌQnG�� 7@k;���M5+q6��i��)���8V�E����7��S�ӧ/�(�u��v�˫r%�r��9�0bFh����4��Uք�"Z���ո�C�l�U�ob��v1��{��q�:��@j�m����2��X̣�Ģc�L��l ^m���Z9�6�\�jm�tGZ���7�e�znó{���مѲimB�0k޻�cf�{g6��!F�&��LXjګ�53F�MO6U�q���V��5�$
�4�[�*�'%	��d�$�Vs�eZ����*��m*w��ǒ�c6bc��A�P�2��a�Z�+�!�'/B"��+L��up����d$c��5��y+v�ǂ��Y�k7a�;i:����	,m���]C��M������`ku	�.�j��J���$���M]dg�t��(��\ܵv�͘��m�֟��nۑS�z�RbȾ{�3��F�#O+',J3,�gqZ0-$��@�Țg4��#kE5����%��0֘m+eܻ ��,|�l�.oh
�z�Փf�H�Fŕy�e�ɦ:(M^�N1�$��z;Y	��.db��8@��Lv��8�e9F]�T�q���	���k1�t��ó[N�}l�f�m�t�k0�<���Iv�1�z�k��J܆�Y�@Ä��z1��k��bJ��2���� =a�IܦX�X�I�ӋN�!��6S����7 f�H�mܸT�{-�9PS[j������7/6�RѠ��ԫHT��{�kid+�\���ݍ�-�*P\m�I��l��l��$�ܽ����݅��ܔ0fbZI�P�E�S���Ӡ�A7vSm�4V���l��"jW2Ap�C���͑hF�@f��g��.���.8���cI'n��sU�w4un�#�S��p��.��JC�6�V�4V����U`nއ)K-��&�0-��6��0�6��7v��c�\� J�)a�3)���S9��V��v0��v��n�:i"񟓵#�h�.��uzv4]�Mj��ܢ�%Rn-�v�2]��I�9�lTE�ʄ�	[���rH��v+�@V&�B2�M_)VoV(B�_:���zƓt3^�ɳ!�@�@�n���or���QVV&>�N�J�7�GHǘR�*�Ve�u(Nh�$
����nXV��i�u��Q+u����z,�Q$U�Ʈ�1
��WAԢ�9��i�7�6(Ѡ/kk�x2�c��m�[�� .�5�4��U����{nE���զ��NlX���ݷik���SA]�T�R*�CMƔ�q鱘p!:�X���
�V�iZ�Z��%���R�щB`+q�j؀7-m��o�����0C0�Gb�P�\V]\B=��Q�J�u�����B��0������S��
�T��*A; #e����8t�x)@��\n�ueL�{i��mvK,�eӘ������y�[$eֻJeZ�p �K���&ޝ)G�&�HC�0izv�
Pe�P��R����p��*]%�v]XͲ�y�+d�I)����F�]jM;�ru�`;�h\�XRJ�[oA�� �-Q�v���kB��#�!��J߂6D�C�%��p�ݽ�IZ�\��6����(NLi���s/J��`I�����$mk�J
�g%�-����Z1�����3��i8.l�j˓0v�MҠ�Ҩ
<�6��áf��ŵ�P� $p���fǔ�r��К�1���5yF�j��t�S ̻�@�1 @�H,�I#�ūi�ͫ����ـ�2jɲ��YZ!�i���l-	�Q��$�u�J�j+MK6�)9��%�3�e�E�����e�|eu��l�,]帥=��|�٭��X���ю����Xh:�\cC/r�R*�giE%�fk�8e�OX#2*��Oj%��I�o���{a^�2J(�b�@.T�B^�F�q-�B�E��֡�(}��DM��kIY/.�������*�t��[��F.���V�/H���#�K\J���m+����ˏ�V��6+ ����Ͷ�Pl(�bCi�P��V	���J7��9�A#��`a:�ag�Q&���R�m㌫ts	_k�'w+N�F�3NQq�KuY��v򝊌�B�רH�+Yl�˦1���h�)r�%�uCs �2\Jk�;���)������῝[��c#���,�J��y.�x��G.�`��!�ʁV��=�e*˼��gXnc�XH=yN��h�
��GV��⊒�{�f��u�	���N���$�(�����H�f�+1Z�vҫrlՙ���+{/w)*�F�,�lC�-v�lo[нMO���R��̹P�y�!��ڃ7��q�.�◙A͢��)��:�qch��R�1�E�h�KF���A�^�u�Ed�	2]�yXmV4(^�q�� M�Te&v ��w�2�Xj�bM�w&�޶헕�K`��ۨ.ILk�w�V�ա�͈⠨l���a���jbr�	�6�lJ����Jʕ*ߦ-�P��i���T�bɩfKЎ�&�Fm�䦶�h���Ѝ�ŜwXm���za��	��ǁ5��"��ժ��8:n�KF
J�G2�9��@n�*mCWt�wW�%5��s%V��ea��lj�ɵ�5�ia��թ��T�b�V	�ůI��W%f�[2Ӣ���hh��}�t�)�3Nf�\;��dǑ�6��v�˱�ړq\t�T�<�#d}y��x估�,D-i�*�n�o3Fk[�NkY0U�JS�הE�x�X�V�.��O$�V\��D���ӵ@i�@�[[X�Tf���5m,2�\̒�U�4;4V�a��j��+ISJx�Rg	��`�)SIn=�C(i*������V2��OXW3]˫n��6Ԕ����6��*L�.�J�Uɵ�p]���B+.+n���ܴU�����NԽ.:R�h��(�"�h�����MxJ�&F�.�Z�6�ɲ�x���>A��V�5�p�xsm�k^�BZ�F���c,�'Jt)o�xt��n�µ)�+2e-7n�����ݶ{t�4�ځ��@�ީ3"4���̀=�F�	2��+5�e3�axve%'.)�[�7	{XİjZ��է��.�U�$�܃f�z�Ԯ�m����'���:�
5��&,�t�pm=8�5e�W��0mP�A*o0��4/6�c����l�n�J9��q��J"d�pm%����2��$�v1���`�'l�OmV�V��
�5����$35f)+2i��5�`L�{�� 	�t3V�~4�0�5��jVӴ0< \ֲd��y��G��ڐ�-��;�I��i�e٭�
�����e=�����K�ܴ$
�Z�^ւ�S��l4��8��T����6�Mcn}l~��W]oj�*p��#-������E�MԦ�-XSqY��*�`��ݥ������T� ��f�	"v/��5�2��bm�9��m��彠���Ȣ��cm�hzܩ�a�
�:p��y��*Ӵ���Yn�N��)���R�Ә��^�:u��5��+Z��Kz�b��t�5�(�`��M�2�`R倘à���m�S% ��j�&����[dB��7�fb���N
#i�e�ɻPyMh*Ӓ9�yp��,��[7]hۛ��!�
�PVl��f�晑�+X�F�19�*�f�D͝���"(/.���g�p�p��A�U�O+/R� �7N,iJ[n����n���iÙQ�YlՃ�M�Vqv��-����Ң��䫼�hiS
f@�լ�;�2�]�R2�N��2����ѵ�쫉[����d�tIfnkuc+ 4�ŝkjL���ޙ�+E���Ԭ���ז���[��QWM`wri����YI&��A��� fX���/ie-���Vn)a�ڣH+�lYU{I&,�u�4�(��lf=ĕc�ZSp��Ch�x��٬:l J$䡗����x7Q�w�e�B��=1YhVnj��yR�%X/�ط5�%%�-�q	F�;ymP�ֳvYW)�Y>�Kj���������zD���N[�K6�k���{�D�lr-f��S
����gaU#�HL�e�D�s+^ӐR����J�HTr����f��$f3.�ygLe8�C�-�g3����@��� +�Q`��`5x�+Mc#��[�;���qL�`�b��E�$ف�jĤ:Q.%m�Ҟ��o-+��4<Փ1L/D3`�t�֫t�a��k�n��k6�Kj�,l��/�W���(E�%�teSԮ��լx��I��hbɍ�{����� �t)�n�J�Ad���jAc�x�hM�[�v�8F*�ř	��fTcU�)�t��˫2��O&�,MA��ؔ��[���QX����	5cZF�̢t�A���&�4v�l��͉ �˨��W�JԙNU�!�7[+3�,B��D��/�wt��͡�5�:��"8�n^^��(���25�4������敔�y��lV���h0�b9x%'�k7R���33Zô~�D�o䤹�`�lǅ�	f�tėVج����+{xH^ɲ9P��h��n���W�'�0O�����h[�QKۚD��j�8�MU �`�;�p�6�6�iPь�[��6��)I�2�V���w6]�e�i�j���=l{ xe*���n�Q�tݝe�5ke��{�CLL@9�"	z#�#E�ĩŖ�V.I/)�t҄��,Z-kD(�Y��B��O�]��*#�ꡐ�3q^f 驒����)̵�P��!�k67�꡴1Qx�f��&���ꭤ�Q�B RWk*�`�a�Z!D���*��MJ��#yf�lҳ�L��1h�g"���i�-�r�٫M0V��^<�9��Mf���b]�S�޾�t�tr�
��~�k���L�R�)�d8�$��*�YE!M;p��5�c�)C�dӺ���^�Q4cjV���ʊҐ	7���-��֦��6ŗ43�bwB+���P.��]���V���е�ëg^k[vVVKNk*���Z�6���7�%��d����@�L������׮�aia�k��"еU��.GyCE���Ǵ�-q�BZ/5�D6����ՎX��ܩ��6�n)wb�%��
$6C�w^6�[{L�U�E�z�ɮ������Cn�m��]�)�D�m�n"܆]@�.�V��Ԡ�v3L�ko@CE^�i����`�
!��ĄHdGX���Xw�-m��=� йeX�ެg��=MC��Mh�C�)Y��Z��m��⋩s�*p�lp�[��E B#��ۏ�$�uuJ���%pH��}/�|���&�ܒ�0��/{����_`�3l=Ħ*9p�Jح�T;����vޛ�N��D9�WQ�Ąod{U��H���
�v�m�<F�fԷ�P���|��FZt|CmuDtˋ�'�Ӹ�vշN�4����B�:���;��v�D�{�^�5��ꁳ+���pEv"\�]����w����y���,[��pq��%�˜��+���Pw+um�ù6P؍�Gl�N��()�6��P�`� s����������ڍ ��fH�f��g��̴�^7��ڶ�R��K#�}Slp�d햹gn�V.�yβ�z���G�t�!�R�kAW1�P�u�8*\��ŧ���Md��r�r���T��3��U�ˤ��F_u6��P���9�oXsQ=ڰ K�,�,�;$.Gi��pͭ����3��23{�D1clH���kU��B8��(ή{MW5�s��op_
u�����Z�e��C�fP���$#�>b�����2��N7�.��9[��^(.�M¡W��O�b���Y=��%�κ����x��(BUµ��:���m|����u���A 1ه2WW��A��e���i��)^ 6�/\d���sw�D7�J��i��u�����\m�˕Ѯ��lM�yf<�VJUؤ�E�p=�N��	};�9��\7��f�-r+y�^n�1-���Nj%��jl�qL�|�4�u2��iN�ڿ��K���ή՗0��j���6��pd��:�e+��@鉴���d��{��B%�Rގv��/�[4ftX�Z]�3\0�msw3���-]�Wy�E<�CZT����z�ed��K����^�����-�p-0�s`崦�!�9�:�Z���֕^E5��yd�V�Ȫ�Cɱ�ѫ{��v�U��y�7N�n��|��m
��I�6ds���
��&�}�v��%K�R�k_|5�:j�{�b����|�Y��|�n���m��]��8ZD7|�k]G���l,�+<T�(��@9���.uI����r��\��hfV�<�l����z��<���a�^:�yJI��rhcD�]}w���Z��s4[��a�]�9��h�)�v��3��F�h�ߔ]��#������oH������P=�����n�D+*ь"w����X��q�������5oJ��}F�/;+f�-:�r�G�pI ��KX����p�EI���	h�e�|N�}�9�>P5t;�\>Z�f�Q��ڧ,BM�
iԸ�Y+�U�� ����wWQu�`8�Z�2�U��$G�ؖڮ��B�\ݔvS�q(�:� e�_l�esk�j���*f�u�o�U��#��$׵�P��=x����ƽ�ɖ���.�-�Y�R��˃;���ϖН�Lޜ��+�WW��&��i��D�ւ[��7�H����w�e��T�29<b�}�8��sAg���ua�t�|:��!f�/P��zJ={2�J�p��M��*a����S���q3�Mv,��U&#�8�R���Ev��v����v�b^�J�TR�,5�!�{�T��AG��E��ql�=����和�&�s*�����h�@Y�B9X/�"���(�ݨю�ڼS�f��ѩ���f)+�42W�P�˽41,��A��<3*�K��Ͷyu-�b���t�y�6�5�4	)���gw6�D�r��r��M7�u�(����
|WjR�M���R�h��z��ڑ����o#	�3�43y3v�>�f����3r�SV�!Ƭ�f�.���:��68t˧�30��6ʙ�!p��ֻV�Ԧ�ۮC;9�=�U`�] ,���ߐ�a	K��V��c9�ވ��>�����j�ި�)�5��ܼ}��+�k@�`��|k�{�u��E���>M�z=��>ɝ��Ħ��A/�p_��_(��1c+��A�% ziӂ�kP&8���J.h��zotU�uc %�;����*P˦�-"J<�KevLYCgb�U퐨!�����F���	�ٹb`$�WuEzu��u����l��N�Jf���fY'l��pK��=]��顁>��W,3������2�U��-ST��8}�+
���YBq�޺C��"�����5u�]��<�}:��ARN\ۖ	jъ*���V��N�N����F�n��Ы[�C��Ӌ��SE�p�g0h��G2Wbt�	�f�oE��.ߘ1��v�é�J�YI|�[m���n<�F���U�c�r̾9����r�����]�\Wj��[ɒ�w:�z��Ӿ��;��:�%X��������.ne���J�K��Y]���w6�h��XT�MWV��
�s��<�ڮ�P���Ǖ0��-'�duB�Xt��;��&���{�l�"�� ��o ������tl�u�A�abQ[}ݦ�b��ۆU�5��e�Ŵ�	�y��BYf�l�[�v��k����,��RƁ��	�R��zT�C3��IMz����e%{P�;^��X�7���m-}��tpV�-<��%�\�+��kn���t�a8��:)qR�{�� �z�/���Iw�XV�s�6$�z�%�/%��Y�{F��5�+N\�o�r�j�'+���˷���#x��Vl��T=�V^�B��dkFw�uu�A,ב�5l�u���]sT�z\9�H�T��Ս���M�@mV���\"S�[7ȼ�ۊ�ۊ莬��mZ���0}�������fU�j\��������r�N.?-��h:&�w,�4!C�ֻZ����[��g�@a�Z��AM�6����d�-�fZ�â���b�R�=�e1#v���lR��e�2mkwʆ��G�u#��S[r��C+S�=;!�t� j�D��9�w{�̤q��U��.�Ά���s)Q�p�@��K$�,Kr��ҩW(�0���������c��������
_��%"�Ø9��©���./�^-yLg]oNU���w��yL42w��#a�9F���S�y�Iє�u�(E.��f��mq��yJ������c�K0�H�+�\��b�
c��5:���R�<��.W[�ҷln�O4H����.�v���h���p���fs�0�8(A8ELVվ������5����۴�W5-�F�5Dg�r4sH�vi�%ì�R\U:���&t�T�Q �����LS��'f
�3���C���ٻZ�4��FP�n�e���v1L�f��H2�Ár�$պ��;&���`9�,�椼�߆�mx֌1_WR�x����j��1O����t��n�.�e�u��'8�[��g+��7�Ξ]��YN��̽O����ڛ��V( ]Xw}txuy�2�4{\�SUu*5�c�!s��]$9ЛG�y���	�f�%�un�w�޶�;U��C)��6�U���kz���JQpWc�Z�k���8�ܰ(��4���C�����J����;M�jf��b-H5���f��1{)Dৼ�z���q{2��u���EX�|��O��`��U�,$Wl7jQغ�]��8�����]��x=�6Tu����7Y�]l���w2�2�vR(܆^��@է(tA���-Z޻%���ִ����7����r�;K
�������b@O��?L��,�S~��g�C[�rٳ*"8�N�O4:�݅����i.�MnΠ�:�%��m�ʾnU���C�|��sB�a��X�wf��y,�,n�m0޷t�e����{��5l>��0�j����j]*�:�[Ϲ+�b��Ni����z&cr��]�;'&E�W\���n��7��ut�>�;>pk8Y��Ë\d�f^�����G|���$t�Ya]LO7SvAy��J4k|U�63��
�d/��,|ޒw��a:�Y��e>��9����^R�xWSk55����M�έU�8uur�X�&���AhU��۬�������M��0������*|���EM�]<��ƽ=%w��D��K�<t�7���pY�8����ij�Z��K������[���5�(Kuu&�S3R�֊����V��o�Tw�;�Y��w0;-�Z��}���VS��-���v�헹Yw��u'�*�TJэ"�X����%�J�]��P�*wA�uM�r�Z0=�y �c&Y"\k�13�T�Ⲁ�ty�+n�r�1Rܴm��T|�J#�j|��o���+P?<w&��G�v���J��&Sfaߌ�-K`t�Q�Ȁ�����!R@Que�M,ϖ<�����咂�^Rů:T�r$+���Z��慅�'<"�X����xѭ�Wen��yK���=����dAf��N�[��W(�Z~���n��(&�����<8"�usNo{v�^>=�B�t��������x�gd��Zzw	��Hڝ�E���Vc.��N�g�@���')s:�Qu��wd�{.m`�#rk"�-]���l��a�Z���q��u�W[�I�n��`��8�嫍X�T���4�`Ғ��ǶV��,6��غP�j�n�S昨�ʺ���G6um�j�L��ڹ��b*/H��S�[��;�w������謒��"�R9����<V�jj�yܨ1�^�ȷ� [1��
�Q����B����y�me�cЌ�c�]B�e���bRi���Keu�n����݈���-:ʋ�֐�m ��1^V먂��e���k�c��r�n�[��rn� ���aM=V���u�s���-Se��SUd�����p�kl�q��"���4�=m���Z��p�.08mݣ�a���oG�� �N�찄�x�5Ì�[�I).u���R[]Y�2���`ˬw�4n���eVJ8.K(=%&z��eV���j!��.Q�%��9W�F�n�˳;&����Gy��u>wX�AS�������)D�ɂ@m��y߼����,�Y<|��M�@c����N�.)>vH/�o]��v��r���.�>���媜s��h��n�<��ciS;��Nvp��٦5�>㥰��NM���C|��#o�д�jWs:�Q$��>-��!��*���r�'H�o9�xC��(\i��1N�e�e,٬�|3���T��16ʉ*��f]��[/�f�.�"+z�]t���q��n�������;��K|�{��|ʘ��)V���Vt͘�ȆPWзqݺ�T���>Se���t"Y��F���>�kk�[\���ĭ���P�`�i���4h��0>[��E�y�7�����	f��w���:C�&��-�q;�f�q� D�72��u��K��ȼ�k�u������\
�=.Kne�y�@}x.���5V���SC�KM	,�|�NKR�������i��R�]e�M�;��c��X��Z��|WPe�<o0��V�D&Ef�+.�bB �V���N�dY����g-�I���r��,p�w�74�~d���8��&>��7�]0��Y'����D�#��@��ƞH�c�}�a):"b������,n�<��ҧ�E],(s7�g�
��wD�����;X,:S�XzA��m�:�9����=^:�ک��~B�]��ӷ�f�4z�yܩ�"��VQ|1B��sqH�YkA�+��o	�Yz���]b�K=ɚ{�Hگ�>�P$ٰ�Ik:�R�jf�zTJ!/4��k%��W�هPL,��k��c�s#�eY̏cY��`�;p49O;�`+	;Φ#�r���TmE0�WhK���NT���h�'������#�Y��]e\�C
�Mr͹N5�Չ�R�m;�k 7�Є��c�Χ�i�؍�iZ�83�V3o4���W>�u��p2�qg.�9C�����n���{�f̺�h�[��*۴9��1�6���S^�jV�Ԑrɒ�Ea��(.�|�䚼�}	���t��3<��h)�����n�!N�Rn�7�j�'Y�_����k�@��ն��j�ݥԛLдz�e��Q��@�#R�Co��vp瘑,��*��3��Q蔔kkIJʑ�י�[��q"�Uܥq� �4�,'*)o+�jڦ�݉�\ԍ\G*<�S충�g	�lS�)�ꈬ����M�Ej�q1B���]Z��κ�����(�t7��]B뀃z��i���).�ʱ��IN�T�:�Ӯ�c���]v-�h�3�xy9��:��`A+mnJP�]Gz��]�Չ����:<U�I-4�4S�㮶�7ܩ�%��4��][�@и拡�Aq��j��qob7vss�٢� �70���B�/�1��-3�uܧO-�����&���ہd
�_Fk��*9*n�c.�ĨӸf)�:�v��)��puv��Q*��ڗ]�_9k0�I�����zC���3�e3m�EQY�{OV��CO���Ξ�%w ��!0�Dvc��Lb�^�z�j�r�#]�1c��A\��/z���}�қ�g5�֩�C�7��Ď���8���޺yK+_,4�^� �V��t��F�Zi���U��U�۹J�B��L�@f^�'-cx��9��Ѹ��+���+4�_`	@ΗǊ�]�=�l2��+6����\0��/aH�{Z���gD]q���4T���l�j���גe�P��X�Jr�a�[���4'bp�z��H�+��V�B\�Poz���3�	N��Jbz>���}���â���ydC�����v������s�z;����Vb�Mp��Qs�#�뒝d��6�gB��yx��*56wJ{s����֌B�I��%����W�ou��8���S�ף�>�V��%�R�ru���}�h�*����_s~�߾��� I$�����'�~Z�^����	���k3i���z%��x�+J�	�x�t�����K����/�J���; %��L}��ƴ4V:T�D�8����@�#!7s��Z�ހk�q@�paM�yg��(�W̊���Y��V�5��kkIs�i �ł<��4�v4�jmN���贾��;5�u�p��.��W�*+"p�7��^i`�~�}M�j�k�ft����W�x:�v�.�������i����[��-r�ո���Ve��}0�]���e�q�|�ֵ��Y]E�	�-�vZ`3�����Dt��l'(&���֗{&�����h\�6��v�B��wB�A+�J$���ӗL��G�Z���!�k�������[F��	�}YQ�Y�-�Isqia\��
�*��w�|5��˭��τji���FEQ�x/xE�Օ@+�+nh�8)քV�]�tE&���;�mk��}kW �Cd���:;����N��ЋGDV�	f}�����x{i�����5 �O�n��-�:�s�[�6������-y]pw�^�b�X�p�]�fQPdw�v9�C;�ީ\�V�cD����F�Vsn17'm1��[t����N�2�QA(���:�M{B�+@C�Y�z%)��gὥ�z�k��$����*��{.j�\BT�&�u\8whn��iĵ���V'׷]ۦTĤݖ��8S�Դ�k�bʕ���u_N�st�{3R��E$p�R��./xg+��褵TFV'��Xl�֦wVneu�%��H��6D7��p��Ӥ�z�� Wv����Y|�_BsQ�J�d˙	GE[z��y9���N�����eB���Z�Uh����g_]�5�gr]�xbk�hi��k��V��z��P��)9yϹ�T��_!Ge�GNE����߀�b�]��yR�)�k+�v*�7��m���n���M��r�Kr�k��Ǜ�3�����]�����d��+ig,� �L�6@�T���n���Všk!Mu��s�)P9G�<���.Lɹ(����{��$0�Gr�Oe�L��5��*�ĚI2�Ӊ� A�AI�tT�KeV��u��:4tW�އΘ�v��C)c�n�ϑ9ۏ��������}��P�5�ր�;)`g�]\����x�����6��nQӫt)��!�]�|�.uڹ�u��π��C�]�y���]Kd�b�Kc!�ӇJ�J�Ѿ�B�l�n��H�l�΅�E����8�14��6+/���N�	�ڒXl[�-�/Q�uv�C*���C�Ԩ��|�m�Ѥu���n�k.�n�3���uT�������p=!D���E>��Q5�P;mǝR�I	���Y�tGU��P��0�$���EAX^Y��U�m�:|SV���噔PL�����F��	��m�GB7g:C��v��u�����6j�wE�e�|���.�h�#qK
=�j�S@��u�x�T��*|��t0��&���Fgy:�/b9{z\���_,�6(�df��7���ʱ/���ct<����b��NZ�5r�ͧ-J�P"��c�'�T���KCyr�5IXj�m�r�-���gQ��ͫ_y>֚sp;Vk�fi�b\��TmX���u|F74�g[�\�o`֚
��ѝe�qV�\��X��)V7qƞ�f�W���u��̱�H1�<�r��� ��Wl[��2e?�}�u��s�YZj��s�>EMIY�*�%Pܸ3�`��n�G+V
]�?0tfj5u��ji-#��c����ҦB�LZfb���9S&�J���{JF|RvcW�>�Z��b�>���q*{Υڒ�or�c�)��+������qdN�����EW0۸�]g;��frܢB�o�����#z�����U�Ԉ[=�1\���=�]p��%h&p�xq�HJVuY����0����_>W�8]�V6M�i�p�Z�&)�D�|��Op�b�-,���[�r�a����V�r�5F���N�g�t����G%q�u�U寘-{��G.G�LC��E[��c�&6��f�\�xZ�eh�؜F�YӍZ�X)ͮ��rq�O�(c��c0���/�#�mĺE��=>��b�5����r��u�F�yL�|��ݙ����d�����oi�0�[��v��'\�.v�J����"��M��.
й�M��01֛����_���^>�����Z�mt�0�0��t�"����n��ǹ�:��TR�v�]b�b�8bW�Yω�#�*;��fClW 5{�s�z�q���<Ն�7�I�O5��6ѷ�aYC�_Mj�=��h�W	,I���K�>�6�5]�û-��r���3.k��@x����.;�T=,b��R�L!��e���ȭܠ�ڮ�vq�s]u���i�R�H���^>p[x��!CTv�̀�7�M�[��bH��R#�e��J�8�����ԻǤ����.y�E���V�G��}D$��l��(�`Xm�Ɩ��j���<�Gh`�ʆ�E�:�к��ʦ���t�lϲ�u���ܸ���[�t��R��b��Ф�:�;�َP����ƷF�\�U�8ӊ���5]:��.=���r�oMڿ�sXli=t��.[�V�\l��@��,�ŵ.�(C������"�M�}��L� ���i
����O�#"�v��j�π�i���ۡT38k��P�8F]]]�W4X�,vX��8��<���,R����[�s8P;������ۑ�L�>8� �,�X�>rqmL��W+�X�s��ʛ���N�_��t^R��a��{�G�%!X�V�%���5���_��aU����uV���\�*�V%m���5n�I���7M�SewMѶ-�8,dk��61�����"J�r>Uu����1u!��Y��[ê����|];���]���Me���@�!4�j��AT7�2�C�r<֭�<H��3{K�X������3�<n���ŏE�Aװt=��!�ں��n��}g��XX	�O�o�� ,����a�0�@J��;ZWKXo)�8v�P��2��*��o�s�
*fpWh�t;:m]����L.[gC)7%��Y���v���b�e^��A�5A��BWs�rg�a
�:�%{0wl����NQ�CE�m�|��/do�*%<կD�N� ��Z�w�W{4Qfd��`m���G.�b����B��®��EC\�5��=zcX�۳$MX�΃흢�fV�Km�)����1>��n���ɓ�![Y�B��̷�u��ߴ��Ʈ��"���A]�rXaP	���{83'2K�7��]��*;�V�v]G���e8kZ%5d&�e��;]q��V��J�F�^��Cs�H�j�o�9�
F�&����=������6R�ʻ�>��9ܳt[�k�iG��v[ɽ��}�-$]��e���^����h%�	2�FK2_]��:�ރ�UY�kEf����K
ݼ��>l��r�'�n�
���W��ZT����~"�j���\�VC�vb��1�[4�1P�7zg +-���Y��t�,�W�2�����v�;K� ��P+Pmb	[1���j�����)�ԧ kh��h�c�ڸZyf���E�Mk� �#4�6)��`ٹ�r
$�KBv����<2]n�k
XzUp���y').YvX�=F�_�	�Ccz�E!J�x����q/��Պl��M�����F��^ {�{���ƋT�A�&Q�8���PL<!gA�E+��Ζ*��U��x�0�3[��QD���]0���Pn�� O5r�ay��4���1�����#lZ$���f����X;;�}�u̽=DX�SI�{���\2�|�.>�aإ$.�pQ�%Zu�S���oR"�}�S��>����L�	��ĞY��ؠ��kXژ��R�$R�k��zky�ި�^o_f�)rWd,�}�wQ%=V�-��-'η6���H:U| �ƺA�m�	����ߛ�si� �f
��s�j��57{^���ɕAt��2op��JT��$�]���ݮ�K�͵}�����J5�k�}�F �)$�'����6�xt]dB�P}�:�RP׽�LY@=KU�V�;���xڵ&]m�K:���c���f���fA����@����Κ���zFBmх<2Y��0'`o@�j���t�����I�.���8��X��w����=��/{�;�
�jw��A��a��֫r��C�����N���cu���F��{!Sb����������^$.��j��栰�v��v%��H��C���������.�����ra���͟>��*�֧��elU�s�ۗ�9C���w^]oWo
��=2�k��w��<6R�l�����K�<���]3��cU����l�/��8������H�>���d�e���a�
�lMh��Z�+v�l�M���KXv[�ѻ�Z�Z��il��ݪ�-̉�� H(P���=������b�8��rTZ���S䆓�!<��COS�Ӓ�v�5��:C�����){��֘�U��(ٶ��w>o�ǚH��y�������}��L��k:Pت�:��ܰ>�T���{�Y�@5�t�۵u���}jY����;"j�;u-���z)%���y �v�W�(���w2�r�j���;����[J����8@��Fr�p)fY¯��䳾�+*,9�*(;k* ��W�Ǻ���X���[ERf��Ԑw���g'Co^�%��UR 5M��G7�}�
b�r���iC�B����7{b�8$�s��կn!���
��(\��Ux�9Ԡi�O���[VF������#�B�8h��]p�Oz��&�7�(o܉2sB��]s�f���݀vˁ�ͤ�	q�%N9��BTDSu�χ�g���{j2>�.A[ǝpTA����)���a���P�ـ>2��sM����6��gP��g5]�Ҧt���+]�h�����4�}k�/�R�-����k,�.���^�֧e-Ckz���cI�VL�j�0��(. ��H��F|;f��	�K�VգeU�5���ˊ��uk�=m�0$O]�q�)DJW']p��3�y��
0)ݺ��S�<��*�WB��sb�­s�ɋn�|��W��tb�-� ��v���8i���aC	����@j�#�jFd>ͷ��8��tFVv݌�8�6k.��r���'E�֥Q�[c;����mt9�;�P�n1���l"lKl����n�����wZR�Q
�h�\��Pqq0�(6r�T[J�_;��j�́K������� w��fdp(%9��ZTMdOa]�O�����1;7q
�u|����h��/�s-$���	ٚ�>����6w������][�c��7A��%d��V�V�p�
n?��d�ˮJ����h{B\�k=GE6�s�h������V/6���^�Z)e��tm�u��27۹2��wI.�s@`	פ�
����j�^@��&���AJ��|Ӹ��!Z�9%�$�8'_L����Ε{��Sh���:PJ�D���3�2Vh�.�yN�L=�/{�
���ιoz�� z���gg;���5�2�Ѥ/g]铅M2�b�n�n�X\�6��K�W�Ը�C��z�)Jq�;4!Yt�n��͡I���j��S_R�Vx`��n�ѻ�mƝ�)��v-CEѤ]�Y��u���RrUЭ,��n��vq��oXU��]A��e��*݃iǢ����p_j�\����ȱ�$��Z�+��c�+�J��id�-D��ZQ³P�l����W3�x���1��|�l�`�{���9���vI� �1��Ve��"�������OXp�E�6��1�m͵��;QXK�x�v�k)ۂ��aL�f��#�^��&7&�,&�#��v:��du�*K������.L����x�l��tk�ъ��\�-Nd�X�rf���/����3J`u �V�����Z'bu�34����)�s,^j�j�����<�m�e5D���nc�vޖZĥ�Ӈ}�����:�PV̓@�n/�o�ջ_v�i��]�RyNf��w�u(/Y;i�ܫF�ޮ��[�C
\���M�������So{����0�Yz��C�p���PQ=y��m=[���Mr`WV�-_Y�ؕo�����X7��:n ���j*�C�Ӯ���F]=����(���ݤ�q��C�LRoXI�k(]uC
�I�	;cvlSẫ9�1\�l�O/ u�5�FW��Ȓc��C��]\�9{%�Pl�"A6_T�c<�
�����=�ZW�{�����G,Ρǒ�⒱�-�;�A%v�hso ڙ�5K� )jTb�mWY]rU�����"5�d���Nf��n�{����}���N�(v�)�A��ڱ}�,aG��s���]���ۓ"�=G�E�Ѽ�FD�]<�B�N��&dXڀ���(�P�{~���%\=J��U��uSmp�X�y�%"�5�gĵ�,g.J���:l����a�\w�c9�P�kF=k$�ffR��ff��4À�y�(@�l�2���hS2 
W�ξֆ�T��j�����ct�Vc�}�7��@�0Y�pUE���Xt� Ę��5�.��{��h��@nt���p�d����*oG��I���龮\*U�[L4��-4"5��,��v�Y,Z�/����I˥�C�U�B�EV+-�x��.���NL�ER��i���rr6kZv�@]K6��2�&���Por�׿Y1�]��[u�խ�y+����糛��ٝ,>�]�T�,D���^����9��/��u��sB�P�~>�:�g��)�t[�z���B�}�v��ͩ0oE�:nwXfq�p\6<넪����[��@R�Ҵl�J;�0��U�3{����ɐʴ�Sk�WL��!w}\܆�
�ma���m7��,���̬�@���
p.vs�*b�Xs5�r����vx�C�kF��rKٕ/��@f�k6��a�X>��=*�u)`m�7��R��T>Ν���;�T�C�/&�6��[0v�=O�e�Cz�r�n�&a�Ǉ*N�Un����pMߔ��մ��IgP�X���cV����fV�V���Lt4����� ]aY�/����j��]�Bgi�m�5�����`�n�I�:j�o:��o�W�N�
�jeF(-
�圇mȻSU%��c��+S�4��Ķ0�չ��M\r��$�����=
��/�u2�hmKt�9u �M��h��q5y��0���8�X�5GK�Y�v��;�m�c�jV�6U뛸�w�e�]��	�u�������:㕗�"��|9��MV����6c�R�ض��MF�Ԅ��0�w�� �f�)�]er�I�X�ݵټ�k�hIո�{#(��������O�)Ҥf��Y»&7�0C
{7�+�a�]�����<��{(�d�W�g�>Ǒ��E�,eY33�i]%�ϓ�g��%)���}YkKUw\z�Vt|��䛦�\8	�(w y{H�Yq��-d|�����,9eb�(�����dY*VCLBz�2,Y�*ܥ�,�"�Ae@��`(V�V�V�SJ�i�������-Vi%DB�֩�D�AeJ�\Bf���*�� ,�!�H(e�
)FTLaY��eE� �Q�Y��U�d��
*���b,���P��%k��4��"�B�B:l��Mh�L�b.%aYR*�"LL�¢��IQq[l�j"�.XCY�"(��DU1���%`VE�jh(,U
����&8*`:���+ *�E���*e-Yu�4�J�BڍJ¥��AaE&$�.a�m��h"���=I|��=}����+�Yڲu�	sv���A"�%�(s����ղ���y��ӏ�����;*I�4
����F*���br �Ee-�lʳ\3ֶ���)׵���~�.���A�_�k�>y{{�-�{L`=�h�C�����[�l�s�u����Zj­ WQ6�7�[�������z����ׂ��`{��<�~�P����������
]4)�G��xۅ)����/;2�50Y��62N�NC�6c���U��*��ˢG�}h�){��'P}/0sP ����6���j!�zn!�Պo(ፎp'���}/�ܩ�\WV]'�V(��҅�����P1H�_us�`ku�^��}��ގ��WS�^�S���o+�]D�8��Y�]S@��^u<����Ƈ�:��
�r6��'| E[sW=Jm<��fwC����~����#���h<���oˉ���vˁe}��6����ݺK�����m+���R����`���,٪&e7�/�zWO�.?:���U:���(U·	��"�yu[��GY5)���j����g:v{���
�I@SY�r#=�yJ�˱a[�x`��黻2t&�$�U�$�d��3���z�Pʿ%~�����+����=Y�)�c�#gxv[,�;�x:�I� <�wx�ޔ������N��LlN�"�xr���9̷����̝z�\+�NKkPq�79�ͮ���}2��U���+�
�6ܾ6�[��]B�
��9��&�q�E�	�+��� T�o�;��?+�W��=�: ct���������w[´�,��%�p]T�<�a8:�ʅ�u�\�#��+�rTq�x�ͧ��U��ج�eߩ6qc/�W�#VMWM
+i�#��'�;va)�l��g*-`�J�͍yݕ�*�۽ E_���FB�*;�YB�2����*wd@)������ƃ�vkm��x�s�C�|�C*�'~��:�v<���`�MJ�[�A���	yx�x�Q�*�veVQ�-�U�*f�N���b�t=*���[�<�f�^(�'��F�J�P�����o����s�_Ic����(o�Hs��LTs���}V�ؽ��ȇB��@[5������6�N��u�T\�W�MF��f�B g��dYa���	n'p����ަ��}�����If�]:va��}_^��S;7����D
���0#����-ӵ��*ͩÚ�4-]��ʞDw�]�[o:�f�|��yƝr!�Hؗm7���R5�xl�R�r��t�h��ޮR>���Q���T�G��9����7��v�i���������q=���w/6rA9�/����Vur��	���{�4^�`�[kt-ţ�dT>�0T%�tŹ�e �Yt���g��b�xo�z�o�Ȗ�Ѽem������\*��eg�������2S��k�"2�|����4��f?e,B!a��,��v����k�����r�Z����,f���_��(�B,BG�e`=�U`c���[2�qeZQ�`p�w���2�l��5�����OuF_О�g�{Gl6���ڬ��{�wFi�UXS�@��0�\��U��c��%�N^������rrVT�m�ü�f�*�U�����?:��Tվ<���=���֍3��f>�^(�,[�F{w�`P}�Q�i,�$�Ne��\I��x9�y�{]�L���u���9���3�����Z�n@�f��௭ڹ	�D�*���Gx䦐G����l����+fe��u��N��s�u�6�h���³�t@�V���b~0t.��S��`B�}�xu��A��3Ӹb�B=��<�T��d�9��S��AVe�u��w�8W�6��{8C�1�ә-�#)l�2�7"�Nz�Wݝځ��{Nq����u��L�Y�q�͟\HI|3U
Vl!��qi�����];�faJm��uv�]�'W*aw);�/ws�Y���_S�+�����|:7R�+�G��ޘ����P������eH��! �����Y�7�y&:���C96�������ʇ�[��;'�%��)&MHb��0�[���M)x�7uˇ)=��l���Ղ
���W�Y])=���t0�g#�-���m�jb�+��֥�IUZ:E���۪�6����{¡�Ϧ`�$W����:���x~ԅ,+1��2�]RP5������ŵ=��|.�7E۹�!<��|�*��+��C.2hGcl@�"cj��$i
����'�5TD�t���#n�,�Ϝ��0��C�ۂ�DߏZ���G|�ޯc���֜8,�ѕz�����J�� N��5�ӯyq}�dp��3U��*>g�N��*,Ub�|�t,k<!7�>�Kº}�!��.ޝ�nc�:��<KS*��Z����r��L���xK�앀��9�Q��u
����\��r�����$�Wm�=yz�ץ^������gZ
q�Y+�`>�|j�`�Tg�ˮ�4��s6��ė>�tb3;[���uIj5W�P� ���]�n����K�id9��Vk����r�0e�*�ܩQ�Z�b;7MT��}�a���5!b���r=@_�i&p�����l��xp�+�}�O3��e�\J�_'ZC]đ�..�qKWk�]G:�Y��o.Y�c\@]I�(C�iB%�;c �Ǯ�
�:��bDK�s� v���9���ދ�a䲬m�qaTD$�#�&s�?`��(B�R衆
�#�f��}�/�l	m����D�ixp��.�%�����)�g����N�wk��&�8�`��2j��WYJ�*�ө�����n"����J�p
�/��0�ȍ���@O��v�VxX�;����vf�� <�"$��3��`�E.��i�7n�;�S�U�m(r���������K{X��#�AC 	��2ջ�. �c����WהB��[&�J����q�[~��u}SkVo+�`G$�h��H���U��i��^G�Q�°A��_vE~+���{���Ga,���?G�Y�ͯr�Ϯ5Lb��:[����r�͎Y,�`ab�fj���y��f�{�jz�ѐ��r���`�e &7{��j*}��
���w�T�X�l�ԫ����'T���qWUC�tAaYw�u��b:b�������n���\\��Y�öE����\�CE��w�:�Q\�+]�m7���Թΐu�D���y*��*��p�5{$(n�U��w�ys�]d�����+�g0�4v��A�Y�v�)�t���E�����Y�uso����ӛ��=nY�ua�o/�w9��x=���6�9�|��6+�O<� _:�hxT�@T�S���h��7y����1�">�a���]8>k�WL�W�}_�����B�T
��^H�ޚ���uڒ����L!ێ��<�5�Q�غ��EM�g�V�[2�׀��U2jec��ؠ��U����7�)��#^�pbQ���/H�]@B�� Wa���"�\�m�8ʹCr�c	����Ffƅ�^����?�f�UϽ�������̭������*�&�b��*�P������ܖ}�l�;�Fn�����ۭHe��)ݏ�:/�����xz���M���o�	f�zJ�]��:���u�s�nPBk��r�Yl��"�%u��ix�y��W^}�ԧ��G|���pR�}�����*y���v�I�ڌ�72�<��o���DdB��p��}=8�`)��q��&�-Sn���;�-%_T'�Ys��8�(��ۃ_Cʂq���B*-���w�mO[ �!\r
�����wkMr�<y�.���;[�p{t��:�%[}{�tܹJ��u4Q���;�+j/*�V'�;�⡵�j������`Q�Q�&��j����VZ�����k&lm��ɜ�X��N�8R�� d���P#��w�zԑ�d�|)m�{�6uu��/6C��(:����B�ޮ�|p�}"awK���K�W[�9@T.�%��g]Mi�+���}o;����J��}�EШ8+<<�5�xA�yW{���0;�(�2��%L�Q�'e�^7�4��,^�ۤ����ק֫�^r�S��=]L1�
d�(��P��|�Prx��o�o��!;�8F���78 	��]f�~�@��S�z U�U�IO�(���M�9�.�Q�^@k�!�����a�U��2��-䭖���HU b�����]]��ӥ^z��`^�-��?p���ۊ����#p�`���=b`e��!��s7�� ��dÅ�La�������I��E��_{�~߼ΆAJ�@s�U�훯n�K�o"i6���{�+��r��fHtȘ[-��R���������T7�G�P��n�]�7���څ�܉�h�|����g�9ʸ8���t��^/�0�ch��;M7s��`���#c�0��R�ۋ�@���[�׳�y0�r��[}n2��1�d��z�P�l�����ZW�u6K���go�(�6��M�Y����>�x��՝aK��� ];qR������0v�8��7��K�1�����N�eh��6���!笾(S�]}"4�I��J���leڑT��w@�#{�a�>2�i��f>�X�?Wvӽ�����2��$��̠����^=�H�����F���X�s����6q�!��z�����^�T�mY@wF���H���cn�*�U3w�[���&0\��R5�P� Ζ*��.��\c�"��R���
�m��P�+%̞ԙ㲉;�c�K�!���>s
��Ü�K[���_ն�� �ls���;�����=I}l�5>~�H?���2�
���>B�Iճ�U�>0
����n�w|N���<L��B��>��ݐ0r���p|�~V�+�+��پU�'U��o��ؔ��1� jT6M�4 [��+���l<;��6X�1���gr, ��H�t[�w��;�UE��`�n��r���{�0�L+;a�����qk��PA��O�O9�����b%eu��Fu�.#Kd��_SwY���482�*.Z�����0�{z�8��Y��<qX�kr�a��#zo�mTD�K�:�uȵj���"9�0��ѭ�2v1n��R��:��v��7vѤrΤ�:+\��(�֏�h��u�}���o��B��R6������T��0g�S��-�[�ul��W]�q�d�5-�`�B��;k���Ҡ���(��k��	�P�tH��O(�=Z��[�Z"���O*�ꯐ؈��^��	��luG7���U�
;Vcv`������6�e���Ҽ!4�c�����3¢�q��,B��d!��</Tƌ$Vҷ<�lW}=<:Y>=��I��^��\U�M�"��e}F����Fiu���ޟ�ў�Y����j�e����F�c�[�����]y ��y���T�����va���ȷt�oRK��0��q	uG\T������B�HSꠍg +���bDK���dB�X�y^�~��s�X�	BN�1��Q��_7,C���q���6�.�˶�t�ry�k�&*z�B�}}G�xIj�|����ok���#MDY��Z(��jd���Gv�Oq��2���
T�@�)���sdlz��	~�)֮Q6�T��ά)h��ofA}4"*6��䤀�.x*T�^�&|p���1/+�i��L�yle�>ޗ*Wqq�xV����FΞ�P��E}�O";'�"��O�=Ov㧸�Vy+ɘt*;��կ��:W>ի����	N�x|&q\�pJ�7�k���Mt,r���w:HpR�箑��`ħ]���u�}[w9����,�ʜ���=�jt=�M���@���\/�7؆R��W���s7}�Ը�ẞq�'�yټ�N�#��8���tP��U��R��)&��膤��\��4 3S'����X����5����t(�G�$Z�(��3��U�q��4�Q�m�hy�3�"�p�:�e�=Y=oLk�q��4�K�7���k�!e�EF9`�FR~޷��s����H��2'~mY���jp`�����RWA��E`�GV���XV]��(��)+���Ȇ�8��:���AU<���N�\3���fl6�Wq�R0��+�3k�y���/�xR��J�ߓ�{��3��x��5�}\"�*�ez[��[<rמ:��2�����p��n8QsL��MGc�qs��tS�>�0C���T7(h�}��\B�
*l {*�	��p�g��z�1�蘽�:{V���C�c5��t��Xxm9L��ō�Zc.����)�T�(�W]��5��t*��J@#�C����ZU�g�-�]<�Y��TF�T}���5�t��w�omn�	��gر����U���|y�>���}���}��|X}�rE-���ƶؿ��o���h����+YP`3P�5�#v��}�%�N��ƜA�J�$@O+r�@��]��]	�u��fbN��-��3�ț������o�;ráOi�қ��7-lM�Ǖ��-d�9�>_(ܟPno4(�%(�I�k���V�t#�d���	�E���-��b��}���k��Ɔ(�ƅ �+嫹x�	n�*��	��s��D���ΦhÀ�˨���˲�w.���n�u�voI�6�w�"���9���B��s]�u�ys���t�f�"�ѝ�;i��R�y��+r�I���I�2�U�'p��Ǯ����>�&�R>�p�+7[�`35�ww-�O�Yp�����X��k�61�釹R��SN�hU9�x��9�+�w:�ʒj��:۩ko+�1e,N�y�i�ά�n� C-pt�m��]_Q��Z�)��Z�,��he�Y�X8�e.-W0+�Z�7�Vu��Lp��v�ᏸ��}�J�X��QWsfdy�IʳX�r�1PH�Y�E"�gJk:�:dg�S�$U3�/jŐ��n�p+�x��Z�Uս6�\���T5Lj��%�&�E������B�fT�`
XM��as�JJww/[0��q,8�f�L���c�u���T��9�f�^CgW*ُGP)t�p/�
AĈkz�U��_Y:�tU�8��_��Y�������&G)���5�V:wc�^��h�,�KU���Ĉ�mk�j��ыj(�>��r,O-�N��I�b�U<[���G\Vi�JNa�µwU��i��:��[fe�H�(pe�7�Vɩ���ۖ�
�dZ�}#y�V��u�]2�;� &������2w]�-��*��TT,��V}f�7�.�_(nΈ�U���Uhhs�֣na�Y�K{�@�c��|�
AΑ:3q��ʥݖU=��
��X�NLi��J A2`5��II3(���
�ź4��;1�S��t`�NGg��^�Z��w���W��`}�f�w���ŐO#E��h�"i&�t=�R���F���r���,�5u��<�FYӢ&����fn�9�ͮ��r�[{�|�0�����Et�q3�]�)ڥݢ�L�bAq�.��fѽ{�t�"�7�ι|�,�&�9�����l,�m��u�pG�:��3�Enκ ����X�EX����ޯn�1!�nfy��at���
x��C)���&��kvv6F֬�����y]�>3 ��VNWYc���+V��y2�pyo�.mv�7�J��M��@����y��U]3W	Ѕ��3�o4���.}4�ඞsx�]�wb��ͭ]A Q����8����F�q�����S��;�CWw3�=�/����L���p☁]R�۹����RÚ�pI'�t�~�n��u��}BI�[���]�r�����)�Btz��*G�Yb,��d}+V�&��;�ߗ�o����B���I+
5�LbeZ�ĩ+-�F9AH�ZR�a2�
-�c+"���6�R�Emm�5B�@�ʬ
�`�8�.[eE�rմ�cn5�2�\b�F,���""SI����"�s D��j&�I2%cn�0h,�(#V%���e�YڬXb��LEq�G�-�
�B�*
Ĭm1�+iq�ʂ���Ԡ�Q4ܺa�2bb�mZ�*([E*�f�2�̶�b�U��j[�J֊�Y+ELeµ�KJ�D�����E
�b����k�\P��*J��Fйh��mhʂ��
cV�WN!��
�Q�FUAuh�&[QF����J���Yb�[Tmے�P�X-��%��cXi4�r�-JʋERP1wm��Ϲ�����v�ճ���B�h���Ŵq:�cF;����57zh1����\�m#����}»ϖ�߇���޽��3Ԃ��m3<�+1 �~]fH�8��I��1�j�i��%`|�f��8���
�A�&*���:���=CgWj�V"�"�v�<#�C}"#{��w}��y���}}�����P�1Rs��I���]��z��4�Y��ޡ�OI�'~fCIY*�jZ*�_z�&���x�N���}C��gi�;�����xãˤ��8����^gz�5�}��lϺ���7���&�� �C�����1��zM$�
�����H,풫îu�6��7�kP�ڰ1
͞�&��8����fE�Vk)�
�}��?}��}��O;��<��{ԹW���\I�z���d3Ԟ8Χ���6�U��OI8�`l�_k}�8��N�c�,���++>yz�i �p�4�ĕ%f���
��'���:5zg�"!�" �VF�K��>�5��8��_�?3+'-�v���u:�x��0�|N��J���ܛ�ĂϘn}�哦bAz���I��c>Փ�����w��J��>�[g�"D1F��]c]�n-���pw��!�
��5N��A{C���ͫ;IP<M�k�+�i�ah
$��v��+�M�{�W��/_}���� ����&��UI����l�@>�>����*|:4Nwk;U�ǝu�8c1������&!��3��1%g�z�C���$I�kwHt�!���Ag<�b�P�4��*c�6j� ����u��'�ןd����s5��|��t<�[��~}��~���P�L|d���6ͲT��7�1�VϽ���CĘ퇦���+\I�g��Ag�:q�Ă��LI�*Oz���8�!�28؈� ��#�"�K;T*{=���w��4��
���g�*J�}̛I�+��&t���L@�*n{�orV��Jã�J��ɩ�a���|d�1�]�!�J��wa�)�Ag��wb+��}#���in�zNݿtm߱e�L�~|�X�3�jp�>C�
��}f5�3�bx���3iP��N{��Av��s�C�$���>��hbJ��2gz�i�_-N�Y1'�Vt����[�O����j���łF�\�-mƻqV)�)��,J�4�ʗ-��.����grm]�:2��f@�Է7'��jp�k��ؑ�� ���&<:�齕�leaVmI�q���:a��\�!ܴ�X�N��n�殶��>�NL=1�h{��8W^C�%kΨ9w=p>�z2x��!~�01��֨��H/��LJ�U�2T���������+�w�m��b|����z�P1�!�1��扴�ɹߙ4�'�ca�5���Ag��1��|�WO�s��pˮhI^��T��a�I��ĝ{Bl��C�<g�tP1�a�x|��I�}�C�>d�������zɰʘ���`��f����;��x�S�~c�d���ܑM$�
���J���c=M'F��IY+57��<I�6ua�i�V�WHi'�W�������L@�^��8�v�Y��d�N2!">�&�9������}��#�퓇�u����*I^���&�M$z��
i�L�=��D�>�f��^��j���m�C�q���g�O��i �����C�6�_�y�܄{�(�tϣ���G}���@!��LC��;a�>ä���.�s���N!Y׺�Ro>����fea����g̕+%Ws,H.٬���cWt�3�La�v����.��&g�{Zݮv1�#��C�bs�p$5�}���!�|�2y�1�Ag��3��h4��*o�u��:H,�}�& T�'��a��~��ƱIP�����4�2T�L�{Eߪ=�p�_D�����H�  #����1����8�I�z�H,���ĜB�>�3H%I�:����v���G|�P��l���m�:I���ԋ4��+<�v������w37�ڨޤ�"�}� ��=~�t1& k~�Y8�v�Z���&�gr���^0׾�����YĜ���&�M$�u�2_���C�����������""�`+Vm��8�t�׭��Hv�C*T���J�3�bz��a��ô�3�LC[ϐ�՚IY���Hq%|O��i ��eR'�W��Ì����_�}C�>�(G�*=�]�S�#�p�Iެ�}�ߞ����풥d��ҐR�7��4�a�
�<��C�=La�vj��H,�ިx���݇�;M!�6ua��*�i�Sh%I؈7ʣ}b>�>��5Mș�Y���+�p�ݐ�̼�����i����;E����ӝi����~�!���9��Z�\�U<�}�3r�����q��,��q,���W�R�z���hiw�,	�mq���'�2�O���y��76�$6�7�m�(} �GލN�6°�=�g���J�hq1�3���VJ���̲z�V��$��'��e����8���v�H,��n�q
��嘬��I�]��;�����W��o3�Ͻ�.�v�'��Ƕ z��SL�<x�:�f'U�$��4M����^'g�ޡ��:IRu�)��z�t�f���
z�ێ[I��;�q6���|�]]e7�tf�w�@�C��f��G>C�1��<�b���6�$�;'�a�hx�C*^��q�1�!�Ծw�1 ���jM!��ל�V��C��o0*��i�w��5�1^z��˚���}��#�!��1ď�OY���>d���1�>d�@��==��|�R��:��*AT�{�xô�i��+�1��1�<�'���͡ɞw��bJ�}�[�_#˾���u����g�G�|DE�b"G�G�LJ�Ο�`�|�&ӝSI��LH.���+�
�û>CL+
����iIP����?0++%vu�@�,�3�}�&�v����<�9�k~����^2�5��>�D�Ж͈�D1(�zI\I�����iRv�1 �@�g;a��gI�1��I�<;��N2�>C�Ę�I�NO�|����/�*�08q������������2��rs���a﹵`):B�>�z���~�	��k�i��fE�2_���ˤ��L��3i����C��@�)��>C��^�PV{�t����O��=@� �p�0�OP�I��p4��b��;�0���J�����'I��w���`)<��4ed�� _���%ea���f�*T���@� >5����3..�_�zT?��S��p��P�LMyg��6�Y�{->f��%@�_kB�8ʇ���0�5�Ag��nN�8�'a�`i1��7�0�+%W�
�,��AAO�� �yLg����\FG��ώ�N��%C���4����8N��,=a��$���e{`T>g�S��|�&$���R|�'�T��d�+s��H/̝Kδm���H�� ��|7�	��e�;{s"�O�m>�P���P)�i�㺪-p]f��\;~�)�qz��߷0� �Z�/
��M�����G
N8��Td;{p�m��*���B[:�⒲���6�M�����+B2�)YYvԂ��b�Z��wb���,�ۣ*ȭ���}7�^H��i�Lg2Ɍ���;M�P�M!Rz�5M>�̙��c�Y>M"�Ƴ���M1�Sμ����/���g7��V6�ؖ�m����ǙwB�����X �5�+���"b��f�\c.A�t�.%u1��0�7j�:ޕ�ÁN#]���e���5<H�|&&"�V��&̱0�eb�I��ں(��C-��Z���\kW�������u��O����������o�c��:�:��^�B��tgG�c�ŉ�Q0�vl���D��"� 5R��i�b4E,�@w1;2Lm>��|[ϵ��6xa���Q���Z�0����k�oB��d��#���'{Q������6U9�YF,u��*����N��6z����0��i�=�p1��@�Ɗ�]=�4AJU�#�^]KC&����R���Q��{l
Ɍ���7���n�Wh�7me�A��x:��;K�Y���j��<�C���vܹ�ٶ/Uv㌽�m!�`0��;Y�w�+殸P{�~ߒ�:w"]hӪ��x]�\5~;V��]��	I�f��2�����L1|���,Y¶�I�VdO�����me�yX��om\���\:�w�Y��lp����pc����2�"(3E�纂��6�
H�vӤw�����[R�!��\�\����;z��W9֜���l�a*�byc�tfjf�@��R]ѱW��-����>|�1�n��4ܡ��e+�h�A8,��)]���h�9WE��ڣJ��N���|��T�PvS<�io&4R5�2ۨ���)����I70�S=G�N���n`�/��!��<%��ҳ��X{�Ƈ����ҥ*��kg�;�f�[n_����]��{�\��J5\ zu�Y(B�s��˯�Q/����0�;*qG�c^����w�h�N�����>� m��͡�{��kG�U��q�ܽ妦fV<N:_-<����J%�/���%��~R�k�躩�a��=���w_���n�Y�7=(�\�5����T;��l�wXd7`h��t@F#��x#�<>ޙ����`��r�%Y�ZTӘ_Ĭ)5_s��. ��\�7 syD7�Q WL ��Y2�VVԌ�]ơ���I�#�����n�n�TAޱ0�!*w3�?6T����m���^����y����Rv�6O�U�G]r�X�1C��X|-�O	\Q���<h���A��{p3�����	2�.�aC_����=�6�W|����4�D�6�Yu}z�s�W�o����\]>+�9�G'g�vSCٻRP��.>�w%N]��Yvz��A����D�և�<���֎NF�q�������t������Uqb��b��"�[�!ra��:�D�J�X��ہ��/�.������̋�J'x���Se���2R�rR�]fU_���Z���x<�����o)`�f��I���U�t��U��!<X�21�@�1�p\@�,�Ek5�%sJg���S���ܶb1��ݒ�3�]��*!<뉸:#D���ё.'�����[x��`��3b�#��*�gTƢ0�Ɵ�Uˬ��m����U�A��Ǖ�S�jo'�5;��"��ܬeR_d�*.g�ɗ�d%T:�;����gKg��-�o����&� �I�����<~�G�p�<���*k<xKJ�:�p�b�xw�W��]�KToܭ;�<��kqq���β� 1��t)M©�Y>_J�sx�ﱿ�Z�W]�نΧ��o/�5����,nt:CE[��C"I���Hcd���H�;K����+�+\��F�ȕ�rM'������:H� F#n�U���yQ!` $z(P��-y�=����{^�t:�����y��-ܔ7XJ�Q���]�u�,.R�n/U֢��l|+T��J�����-VdEu�{.��]]yC��ٖ��ԐĲ��kwΟQ����g���靵��y\�Cm�؁C�f����ЮW�*?�>��0�i�Z=����x_��WgK�ӘA�3�V;�&��tX�_A�6y������� ���u\M3X�*{Bg~K���T��a���!(�n�݈u�[k��˃/i��	H���K&&��H�����i��1K{V�WRyU�a7VvS��3twK�C@P��Ŭ�f^�70�FV���9�8�;H`W�4���׽�U�<�EPH0��Ԁ��MP�s�p�<�J1�;p���^���+3)I�:t���7[c�2/D^��CT�f� !
n��r�Ͷ&��&XXH�8*�ͣh��8���[�:��Z1Mq�UZn4�fgDGt����SZ���F�nT�Q�yS��5�&0=Ս��uTf�o2�	����p�u�V�W�g��>�%Sկ���F�5qZ����Py���V�z���d�T���戫�\���_�0���h{'׳��G�4������]�njutfE?�e���5�Q�,�ayU��WBƳ�~9��\�!���ɺ�����9$����VvO���^��"��d��.֮ᣒ]���;�Y�����Db|m�+{�s_&��)��s�:���DG;ps�G)�s6�:��c�����L�.��;�,���+�-��R��7,����ig[ũ��k����Z��z��l��Q�<��f���?����Ar8�O�y�]tH�3%������{=����H-.��B�g��t�
o�o*:��ҏ=� ����:�G�Yҷ�.塔�R�bl���W�Rӑ~ct�7,E%V�Y�w�PA����OPI��^�t<�@f̑eJ���\F:�X�ԺH�q����6�S;l�Fo&���j�����<LJfʐ*�Hk�K|v���^Z�c��״��ok��;I��39��ڛQK��+�q�I��G���eI��	���Į1�
���J�u�J�5w*��:���8�`�(N�Vg�E7#ܶ��_�B��^a�$�o3���Sr��r!��w)�فh����� u7���; TvY��ʷD3zqYj�22Z����v�l�/�A1bcz&}	'��!�8'1� O��9��~�?j�p��O���Y�!]_m��l�&OiA�_j0�	���ܕ�o��M_����WD'1���H��4W�oH�[�F�,��Y�����\��`"�S�'Rʻ���#�0���}솓=�^��Wt�u�W�Sw*ޥi����5B����-�j)�7��ZU�6(�aS�o ՃlC����1�H#x廪����{��0���CsfrD(�rZ1qg�Y���\�b�y`)�y8�~���n��矎����yF%� ������M]�w��C�z�@�0��e�B09�X�Q������t��j���n6������:�{��O`��Wq�r0��;_X�Ɏ��u�l >�^:��M6��!�[ W��c=Z�D&��P��?sn����hL?h��Z��{�r(�s)OU��'vDq�*aF��p5���������-�0oϲ�[�Q�*p`=\6�"���c�pn��-��p�\;����DYC���4�
jC=�Y��b�kw�&�2b�D�%���z�X}��z(�J ��iᶖ�g/�F.�V��^��g�YJ'ۄ(��䟜����
���eW-`v� ���	��:�<˷�پN���~�Z^���j<΢�<���
���?6l�����w>&Y��U����ObՎ��,�Ѓ��H�7��6�2+�ߔ��b�z�҄��{e�Mc�{Ȏٍ7�����r�~f��(v냶��)`u�l�Z��a�W<��٪������h�{�7�l�|%[H�d�kid4�v��HZ�,���ab�J�d��۱Ӊu��[_�O{;{�^n���MR�����E�71FV��D�p��������9Md��cg�o�y['\,�f!��=�݁�*-�Q�.��!�(�A$hm��}:��T���C��qρ�wN���53��|\�.N:�����y3;��t6&�2�T����;����������CX0�j��c~'�ƕJ�ڞR�<�M����eb`/K~'ĔkD�z庱��l�B��٢x8FK�}�T�g�Y�|�+����vY4�;��9_e\�Xa��p0��s�@����c]Qdia���Z_ν�2|�Ɯ�,u�e��Z�0�}��P��{'^$�p�oU���'��T0.R���2)�}ΰ1[��q�:�.Fo:$����-q��)oG%3���5�@ʌ�`U�-�8�� >������#p��t&a�biۉ'�=�%Pۿ`�t������������^�;Kw����0hzY��|,�͓i�kw��xx��1�7�����3HC>��G	|R��F��l�q�SGT}"^��[��z5wZ���oDmZ�o��v�)�P�3�֊F���T��n�S�n3o2,�j1�)��1�r�is&���Їr�o�c9�ڵb8gwh�v���/f��Y�j��Ƭ8(���#qm���
޺u�S7�T{0��m06�T����[[B�5�\���<YqH���A#�mh7k�s����m+�:�b�_S�#Uv�F/w �33��ԎX�L���A�t-�j�2����������Բvp�n��V���0��Ļ�F!:m��}Xѣ�o0�]�Ϗ3�p�;	��ٝ�-�Gp�[*Rƶ�v<̰��í����M{��X>/m-69�t{�tr����#*��y����ugwEZKmL�倠����Pg+,ʣ)�H3݊��o1���Yfn�ި�u�\�����,Ǎ`�Pmf�]����u�"6`�ˑ��[��o�)��̡�����ʧ�� �5`os������[� \���!^���z�������,զD]x��l>�]�,ϠɎ�Ge@��*�e-�3n۬�ͭ��h ӳ}��]A+S	VuIx���K�+d���e'�4��;@vr`wO<.�A�;�*oa�]����T#����L�������M-�W5]�IM�2�⯲Rl���G�GV�u,�*����ԧ^ �2a:˹�R�lT��H`[+�I���r�GY,�q˲h���7ɓѣ�[v��X:_\6�n���ð-l���\��Y�;E��� y�7U����1���J���f:ٕz0���n��{�c��U��Y#�=�i&S��4�-�ݥ]\�m��Ě��b�A�.����]a��Z���k(q��lEW
b���J����<=��0��� ��mq�W�ԭI��Wu�#on�	�`^�e���u�w�n�f��n��D#�J����pn
s]��Wп�xk�K~��p.�B�d+
�>�͈ۢ/�e�-�U�3�+b�n(c-r�)��k�5�#�F��C,�#�JzwiBjbN�;����6�4���j�#/yك�u_R�X̨�\�o~�V������](�V�<�k�G�5o���\[p���!�Ʒ�P#�S���{S(�c4/G6�{v�Ю ���$�����y��Y�2e3/x���*;ϳ]%���+\t�*���+X���jP���)y]�@t��.���?.�`t)���\��G&iMWtQ��ѽc8Gϟy�q9�;z�.J=,������;���;`:�����;T�t����,=Yd�6����E�WB���z�}ֶ�����j�0��h=Y�� ��8�s2�����4;�yN�U�{p�5�_Ma��	��U�ʱZ[�lY�k�ңmt��+�|�#Ok9s�s��������@i-.]��n�-��.{;a�����t��i�1�!�x6��WT.��C������رd�N��Щe���*�ar�̦*V�nS2�"�*b�*KZ*�0�2�e��Cp�I�+P�mֈ���ۊ���eb��偉��,ֳ �kl��9fe ��Y��ڂ�l��Tkj
J¡Q���l�QJ�mhV�MD�Jʖ�-��nXcPĘ��Z����[E��dY�
�PʈTQ��EX��RU�X)*J���ɦ�&"�3--���QJ5*Tm�kaP�X�币T��[Qj���R�UDr���PK���I�������X�W�md�*�[dP��CL�)B�QeLb�(.��DQd@�|���IV��z�B]���[l��>��C�.�!m��]v�fD2�[N۸�,��3���Ѿ�:d��Ó����!~�������W�2��l��~�\P�8����ᖕp��eyK
�t\oA9��H����*����dEB��3�lt����檻%/�K��<w�X��ml�r��S��w�ܺ����8^(�;s]���uuOL�WSP�x`���	Q�Ѭk	&�oR�ޅ�Ö�܈ڄ�G��_Wܩ�G~N@�f����멋/*$,F�3��)'���x������AQ��5p�*״��n��Ea�����Ep�~B�_�!��x��xߦj����`�F�
:,dy���5>�\<�!�^Z��W%cǕ\Yoc%��	�7-��(t��Ȏq��/A�@�0�ǭR��^&�>�H:�^Öz�¼#��8���T�\��y-~�K0��;W�!`k��>��I�4M�N�+u�ei?LS��XP�)�P���z�\�`q��[3+���.�l� -�k�B|7!P{M��)��ɹ�_��y�-�.�f2a�Q��ldG*���0KuL<�����a��x=;2|/3��9��dP�)�+xعn��{s��R��t�Vmy�O8=jns��3NPu�����E,�v�7)\Oh��s�2�{��w�M��Oq��D��l��q]��s����b���tdI��Cx�����Wi0+R0-}������&y>����ó����d舸�p�U� hl�/���u��G�F�����M�Xǉo�u���JMh�B���ݵ�f_!�o��TGqv�AMW#O5��I�vg�S#��!){Ӻ���|
��˶��4E^�U�*���/ʘw��Dz�b�ZQW��p���ɾt�ɜ�z�eh�Om�ʊ1P-�/�B8�ZzQB��v1�����.�\���\�݄h�	u�9��p܇u�o�_�XZ3j�X|�#PqҾ���:�7��>-˹���UBe�Ύg*���R��')��Lh��Vp���B͐%T\)�)�e�V��ۧ=�pe������J�1!3Q�j�T��i����b:Ӷ/�V�Z��k/	S�g���	��HY�c��FT�0*"�F.0��X��O0�OiZ~���1����uvq��.�h�G�� T�$�����t;+�Jθ^}�+�;<����] ��I��nS�����fQ�L�1�KF����*�C���1�
c��u���N�7\ĕl��T	*C(rԒ�� �Q� $��y�=�f���Ch�)gZ�;ؐ���}��k���e�s�/�
�R�ǝ]`�+��c5�$���� Z�(sˠ�쬗ڷg�t���hՃ|�#�(��_.��pn��R3n�}�̺5�[��C�)Sp����u�+j���2�E5!�순��X�[�U��[�yg��'ݫ)^k"u!L[}V�C�� �C �����P�
���}Swm���G�f�1��b�[�����ȿ��Y��T���m}��r�qS�o!t�wB��Gș�}{�+��F励��r����zgfk
eG+��c"9���ڪ��Q�_X�:g-��R;��3$� f��q�;(`���.p1΃;H	޷��Ds�Q�"^�U���5���űu�'VM
mm�1����pʅn�A�<7�aYu|�(�\j*­��9.*�7�)+�) �B��H��Yv'��'�Cy�������§h�'k;[=k"���E� .� 1mP9gi���tPQ���BYGN�*Й+GZ�W��n�'Ow6g�!?{µ r0���'�crễ��e[���h`�7����=�A����qe���nջ2]��8׊�c�+Ӱ�
�g���w1��֘΋�j����Pnn�V����L>�����fĥ�{j�
�Z#;�xu��|!�@x�vԬ�4�9�c�i]�f]e�FV�șR����ԣ<[ڔk�Q��11�LJ���ְ��7g
+��Rt�ܒ��os7����1�j>J@��[�_U}�ո�L���T�Ux;�v�~3�;|(Ġ
��"i�ZZ=t��Lؿ�A�q��}�(�z�-���ђ,�כq!���8�f���*�	��@	��jk6P�g����n�*\_k��g|�j%�܂�?7o!�=�_�~HәP�T�)R&�px9M��Mց5�^w6��^�W1q��I��TY`�����P1�*�Sz���̩�Ns��6�]��S=�T�-�@\r�~A��BS0��/+A���
�h��"7����������v��UF8(|~��g >9�e$���U/�γRm����
)�vA�p�5ep� ���8��;RD!�~�R��@(`�%N��C������ ص$�����A^@O�P\�<N���Z��V��8�1C���ޚ%	1]�PJ�3�����t���ü�a�Ȃ��5��&d�ӑ%���mHW!^ApV3��W�����nLT%E7�X|�Ƌ�TY�N�6��r����2R�rR�]fU_���k�4������X}�V����[si��z:����(���B6���@�h$^ef�z���Ѓ�����*=�{]�Z؟���b�Dj^�^�/�gi��s�Rܴ~���Ҷ�J^�md��t�ku�:��\"[2u�m��2.���}�3g���-�����Jӳpv�P%�����'�G0�~�;v~�8��f�n֩�%\a�/�Ƭ�11��^J�k�)���_�z�Vr�*�Ζ�������Ǝ����f�5W����b� �W�zΙ�*�&u�j#`��}gV QL�,b&��ᔧ�����:�~����-��{���ܦ�5ժc���_V���鑵��l���}O��8�\^cQ�mv��甑�5�p�����0�@B�St�	���-*��%�}k)�Rī��e5ϧ�˔0\n�g���P���U���)\�Wd�_J��e��Ov�g��;��B[����?��B�����c�]!�:��/�ω)�2�Fk��Yk�.7��cC\f���(�L��ڄ�_m}\�$r5���bp\��/�$,ַ1�J� s�rB�N4Y��v�@��C���%���0���#��#
�r{�]��.�v�B��v@�՘�ʕpuF��ޒ�*�-�PWwk���}<�
5�Ф��3/��=�/]d���,[(����O��kt�Y��I�PKt�����2w*��f3Z��s�|�/��}��-�ZM��0VG-���k;��-Π�h���/"���8�h��8I����I���nRØprw��IO�����L0�!����!��W�_}�َzu�ti��O���V��2聱�%#�בRɉ�[Q#c3D����.�TwW=j������X�urn���d'D��SA�M�Nڷ]���?'�h��]=�J�v,��ݹN1I{�v,:΁�A��
MP��ST5�@i��Աۆp=;`Wcy)��3��)5�0A��a3Y���j��o�X4S�a���M���c8g�?Y��=Д�7�7K�eD^Vó����fkLGt����kY���|7*~�R�z��TKr�7Y؏WR�*QXA1a�p8eNSd�
�+̫�3�G�N����g�lo��R6�����b��_����#���m4��0��DU�\"���~4�U��V4=�c��/���;}�{s���v7::ᬾ�QF�0��%�`���Vk��P����jw�Ѣ_B�bM�et�ю+zr5L1��-ȉwb2���u���ѧg��Oo.J5��N̠6a�G���J-�5s,r9���(<6��c��9Vu���Du��)G,�Z�!f��λ6������N�vѝFf�f��A.�_�C���qFC�܋�ε���gN<p)�K[�M�D1�Y�c��Uu!cb��;��mǩ#ʷR�vb8��;݇s�j'1q�j�?��\8�a���i�PQ�xz?G�}�DLӹ���^����8�mDM�VA�	��յ
��Nj�c��2�J���\.��y�Ml�fqoW#�^�{ݝ �'�y�)�1������`C����4�#�R��0"�xn�x����s?1�\+'�c�x]b��e@U���Io��k��Z�c���O�ӿK^���b{%j�oxv0,c�(�"�х� �h�Дʓ htz	\c7������dҍz�з��t����c��ܡ1Hjw&@zj�L(!��rce��.21�m@xq^�ɍ�&�`��oj�ȅ;LA���������*�;�C�T�oTC)]M���߫�E����ka��b��oH�th�ɪ������l �&�PGK�;��UNZY')��#D�r��u��Uk��p�m���Up���V���V��P��#�ã�Bq�-<���I5��`���1G%���U�"�\�3Q������1�\�7�E���}�×*�Jg���ޚ�2�=Am�A
�f�p���xAaYu|�(��7��߹g+�Rͬ '���Ȯ�]�x������2M�;+��{L�Wy��PR+^f�}�# l�VN��p�E�4E�-�<�����s9QI�w���!�\���^�۫gB-���R�.��1�i��;(:R4��=qM��yw��#��I���L�x�Uj�Y��ވ����x� �O^��(V�*2��`l9�*�F7��5�{OD�,�X���6+G��!��{!S�kz�v�0���� D޺�r6��Cw�)�z�{0?�wXx0�X�����#�������l����j?mJ�%F�ejvɸ{0��#t�(h��F ��;*�ЏwX�E"���x�YS4}z����ީ��a��xt������SV�գ�JI���Q���4��0��
$�#Y�?��������h��6#�6N�����s�ŕ��=�ᚵ?_\���S�q˘�@.���z�ǝ�>���Z*��{���yѣ���t�81��>�E�����ݫ�0�_ч�9��}U#D�H�{ZEC�q-\���\��uCUQ�
T��7��@�Q�t�C�?)]u�4�UoZ��a��s�[ܙ��yK�_Dm|��h�W����yZ
�@!FGI���m�+n����4F��`@�n���Q̀_ӐJ�Q	5\9�.�E��ul��t%���	�BRÆ�)�EB{��#]"��g�+ʊ��C�&^��,|��2tC��4p�FT��oM*�E�:��h�a�5f9D^�j�<Ķ��Y�T���E�ڝt���웛���[��х���*~���>���򦫳N��ݨ K���R�e�"`!�~���;���z��P�>Y���u��N�<��hi"Wwۏ����J	�cWz?#��j�dQ�\����卓_01Q��-��ycX��:�Ջ,��.c���w�f0;���"�h	�%����}�r�-ɇ����-n��2��уEj�\t�2.#��O_��Ǆ�)s閏>^cNE��Ϸ��嘞.7bp
�S��M���+ϜCٌu���� ��L�iUC��!<n>g0Ȩ��s�:a��l]d�b�s�=�%����g�������ʥ3��t�ξBS���q��v�LN����6v]�Z=7v!�8�X�>G�D���T�}��kymˬ]���2�D���{�_*Ğ��G���o��F0BF�^V�Le}����G	|R鑵���D���9gl�ZQ�?7���,>5�Q���G��`��T�8k<xJ�������K�\ٞ���Z�{��zX�c�h�E9co�Y|7AW��0�J檻%R�P}�{�^{ks���Q�p�ȵ]��#�s0��*�`7�����+yV"�i�sW�Q��͸�Z�cGgs�p�v�k{V���$5��Z.�}z��Y�Q_[c��ʔs(*��)���'+^"�M ��������	�����5��`����}}
������xT����<���/~~{\j��Բ���4爹gT1gd���2S�3ՂY�Wm֔w:݁f��JE�Qr�[�	�_Trt��rj7�'�T�3\�i���Z�u����8#ƺ��Ymػ|=B��������
�2Z��Bn���L��c6��|��g;ܸ�E8}�E}|��4��	L�;���1�!)u�m$��WJUQ�9|�:WY����nbE��5&�/�JG�"b~Ɋ�LLRډ�)cu+!�rv{39"]�뺖��dgp&��!�T	���!t�zM�N]R�]���?L�'ON���ƽ�B9%���5��
�z�!|X���d)��D���c`Աڶ8Ǻ����}(���e?R{�6��t��N$z�N��()̰���č�3�����&ỳ?�*(3����eE�`w���q�����.��3�����s&Cɽ�[)�ʔ�k��v~{�S���&0PP8eN>*ׅs�+���xU:J���Պ�w,��V7���7tۤ���A
�;/n.�jՂ')�5unj_9�C]��hta��+%�ѣZA�]+�UqF�`�9�� 
ܣ#���kǊ�$;�^3,9��b�J]�Xs/څ��T�w����6��c���[;Ӗ��m[,e�J��-��TL�x�Թ�*��-�g$�r�)d�E,?>{V^�0�f����U̠W۔��t�c%������j�^c���HtR��<�Q�Y��-�	�C:.�r�P�m��Ȓ��\���o+s^f�v�:�U���W.��ws�W-� T�^b��Qò�u#g�N�f�44v���@�Y���3�ʕ�*G�$�U�<R��Bqe�D������\:�O��е��guls� +8!t���qu"��ou��۷��(HaE�ٮ��VӠ/Rt�� ��L��=�zN �\�-�t��:�߷wԩyv�K���Q�%e*�	we񩯮P�@q�s�Mm�;¶rjҽˊ���]J����Ī�}��}���Ʋ�vη׍Ⳕr����*���zMC�ê^����3�Ī�"���4-*�o����u��(�
�Irj�Cӱ.��c��i6�<��.�o���PZ�i����>�R��w/���۸�(���#X�:ί����m�Uz��B�m��Z��)hM�Jb�u��ʟ`�5N �:�$�3�^]1���/]I���QV�{	��ɷ�=[�o��&���g�ypTdeˆ�>���O�q��SƢ%�T�d`�]��3pA0�b�����'-pEl*j��F���i]�<�Q��V{'`��%%r ݮ]��m���:�;G8�b�B��)O&ӕ�v����)�7��ں c�R�Ŵk3T�����o��nF�]�nNͷn��m�]S�;�w�G�`��!x)5�t����W+/ �붠�r,yS&�ȷoa��ù��<�D���8TU��f.�n_=t�z;t^R�,8,!]�Rӆuvj�V��F�˚�XZS���J;9n��7?:��m\m��Y�߹we�]���l'POmN�T:��\�ʮ�D�C����-�8��G[��ZA�̾�mD���!A�P�н��ңս��!�{ɽ3��qs����{])��nT��s�n���И���V�%��̚��t�6���2x���5HmC�3�EH�&M�N�r�LS��h�ٶ������y��ubI��6ˤ�s��"��bP՝`�y7�b�SZa�|6��Y�Y�����R��N��Y�G'Y�*Һ�t�U�R]޳\6�v��Ԏ{ҳ� ;�y�1�'ua.������ �T[զ)z{1���P����T]�Զ-]Ý�Y��)@��A[GfL��$�����{�^{�v��f6(��--H�j�+��j���k`�P�J�Tr�b�"��1*j�Z��b�jB�.R�cLl
Ų�J�-
��,Y*���+�YjZʕ��E��i*TQ�J���V`%a�̕�P�*�[�D��՗,�S.�LD(�-��VX%�e����B�Xb�F(c[F������YR�-h�յ��m�[֥FUmkeH��TV5����p����,Q�Q���2�+DT-(��ж�TZ2��eY�V�ѴB�T��TmnZ�DrХ�%j�jQ-
nZŸar#��JZ�FR,+�֔V2�b���X���Z�%k-�m-ki[J���Z�����m�X��eE+*�Y�]w���C#�''���p�n-��fp���i֬�Y�ӳ�Sz��JyˍleE �۲��-�ss�a.���������� ��}a��f��	W#n�,�ύ��N�� 3�"��D���L;�$�vC�i����]}�6��� T]�f/��j놾�<a�V��s#�3+�������ʞU�EIܙ\�l��6d!��<)���m��/��������t��Oa�
��/n�	E���omB���}s(s<�~��A��})��a�5��ym�X+y�y�{ku��s�z�}���t̀�UF{���Ą�F��W�Rӑ��7Ke��ܠ(���z3���
p��=�@���/ ��s�x��=���"Wn轴�	F�D��������3��\>�(T��W�&	�M_O�^�{jز%b�3ؕw8������q��N\��1��qUY3*���t.�i�$��q��wM�)k}�ȼв�un�q�nG�^Z$�Z��$�p_�i�~ N�{O"5�XW���o��3��+#�!���L�#���/�F��X�Bd5)t�mt*v����q󂤮��J	ǦMk���y�[�p����κj���
]�Z���탁�Q��J��+*�u�d��|[���@��W���--�ݸIv����h�8�g�8��\����j]�IZ:Q�]_���>��5%np!�c�`��_�Ñ��s����>����,�ٜ�!��ս�:�%���=C�gX]�������X�'1�AWڤ4FrW+���JW,����Xj��z/����d?-)q^O��auZ��@�"K�WS��{�݀�?�]	���S����6���9�~>}�V,��y�AJL��I~}'�L��b�tWr����9�x1���Z{:M~���>��Q��En�ɽQ5���7���x�f��I��j�P�R�՝ӻ��<��"n{�p��D(��F<��{׾]�׋{�t�(iT��+)�'z�vd���	8/0u��V��qW�_+�U:��ɦ����M�*�|ui�]<�}����C��;�4*�ʧ�b�窔0vQ���%��}��V[}��{P��_ì��nWȨZj.R����� 7[Xsp���u��v+���5ZPM邦�{S���׍��q���^�K$�Yg��5�ďf�z�<��46�Bm��顖{]n�����F�����kŝ&�tIgy1���ʂ����U���'Xs�Õ���Oc��vܤ����M�0oP��h�z>�舏��i¡��b��ݴ$���x���~<���7c��Y�����`��3�b��c��|}T�eV��
_u�qܱ�˔Rr�`���#��uo	Z��C1Snzg���e�؜��G[�y���8�aTʉk;.&��z9֭򼥿mU����c9���#��ʓ�۞�p&`̜чq���n��s��]��rel��do#�Y�f��6o�>��QЮ�jn'V�c�t�u�P���>�Pc���pe���me^b�zqc�����a^)e�<���'G��Q�>�3�� ���-��A�����o)D��XgA�=/=�
�����bWn�T�����hQ���u�Aq�!�6n5�.�AU�q��W���Z�����8��V��s�7�:�c��뽵	+�ںK�8��z�\[AqӋ��-�Խ�O�Զx�߼���}$���-/���mlO-=$�D��q:��A�ٍ��c~�?:�G�7�yc�51}wQI"�oܢ�qs������"��`��mv�['z-;]1�|o7����L�-�i�uН�:u��$���ķ��\SP<)Z�=��>�茹}�T�ݫE����7�Y�z���\my���Ǒo���X�qѷ[�kt�Fa�q��}	v��pj�	q���K�T�Ρ�C���/M�Y²��|��K�\�ަ���S]���[��H���h}��?fl��mnr5}�6#ENPͫs��wE�Bn�jշ�ՓjgW6�]W�����w~t\+7�Xz������2WW��F��P�5�i������3�/��i�8����ܸF�t㋯1z~�g��.�|G�ޥ�𳍰Qmf�"�*7����쫒j�8����`���O�+[��~����^r�+�z���E`�CQ��BQG{�����}���U�H���2������)��}���IC�G?��Ř�!wW�L�nI�-SI�}r�;����cR���l�|��l'�0���/�ͬ�C���2!*]݊�#�������/��h��aa�ǥ-#h��U�wm��A��3����
��2{k.�l�75V�5��[�yoh���b�FNO���Vp+�_C��m��^(�S��5f:w��IZ���sf����Z�PV�']�ܯV-�F�]9�ż:L�ܩ��k�#��ʸ;��k�}�U}Q���ή��j���vt�j�ޠ�SV�����_.�;L��N3b�O�uo���O��)�T�򱋽�8O^��Ơkf�fN��Ovw��r���\��q�����T^c�7�b�3�'��|�9�)p��ы�n3Κ��<��rl�mh�Ek�Q��K�{i�I�UcIէ���T�G����sk��������K���s�����Mj�V��4��|ֈ2��W�碹[ٴ�SW�q^��������Ι»��Am�u�i����U��_iY���z�n;ݨ�����|�L��	X�w3�ۊ.f�MA����*����F�U�<�MC�U�>���n%\<|藧�C�<�bU��ʅ�p~�މ�|��Q�UDh���{瞬�bT�bE���a��n�qB���n$ܔ�k���]4��#}ر.�X���)ɎY�{,�_�{tP;�����b�&G��kA6�e�gO��A�@�3�Y.�څ�s u���m�Z��x���V[/8t(�3u�:h\�#EVƚ�L�����	��-��[ؓ�Ȼ�)������iS'S��V/CP�oN[��Uᄣ�^}'��Ϯ�.v6+ܤ�!e^�7Z�n.r�
��S�ceTa��F����{t��7�e�<����L.̸�n�S���:��U��JQ�j��b�3c�OnS�iN,k��k2��]��ML���f���u�J9�":9�Z�����;�ɶ��hc���e[k��bǶ�����}�� �MP��=��}�㢯k���0�7� ��)v�|�R�aw�p���),�tw1�9��k&s[NT"�C��ו��/��UĴ���W���sS����p���>M�MCX2���du�U��^�̦�Gf�k[=�ӛ����Ry��ΐ��g��t����50�^&���د)�\>9����]U�1�k��Q<�䯛ިj�j��e��(�{2,Z6!j�,&��+\�gR�^��FuY:��ʼ���Lnv����ygL!�7�=2�4;D�hm�â�u���rn�1�upC��KT��ް)��^_5E���:��ާ{�-��;&V�ѭE�R�{ݩmn�Ch�.��b�p'�������ԕ�jw]�)zf]Q�B�b�U��㹱i���p�b[�g:*�Vu��P���k�Y�,$X�5�e�Ue�R�kyF2�_S�Fqc�[�֛�7ثq�m�}p�%WЦ�77'z&�*�,�qU:8�;�Z�^��p?I����Nj�6��WW�$v;p�j"vҔ,���MwLSn���nF��n\Bn�-�˺�>��-�q�R��	S*���=qW�x�R�����L�!_Zk1wDV�E�kqܞ��r����ϤV��bꉠkG>b�@. EoW��?��u��s���� <���#+�_�b&���H�N^�0���J�F�����>��Ҳ��΢�<��6����mh�ޑ���窸�����/�cyo�}c:,ߗy�|p]C�]l3q,�=�5;;o_5MQ�m��t�/s����U�x����X�+^�R1qx��ꛋ1:�	R'&�09��$Z��֤G`�*�o����]ɡ�r��-�}���dl�@��Ի�`s�@����m��>,��FV��c[ƍ��ҹ�J�l�_J�丬���U}�iO��a��y73���YEj!�Bj�S8�,Zd��/��>p�gP���C2����ih�\����7)]��!�43[�hQ���q��,k&��c���x�P�&�o�)Q����T����R�q���'�g�L,�`b�k�u;��C�,��H죊��:��9X�j����LW;zl!1�c*V���jkJ���\^uʻ8��:�Q����L֒	{�w׵�y��h���_.�K5����f�����o�TYŵu%�	��mV�QU��Q[ó7�����;{P��%1��bPU����o3���\�/�eߤl��EuE�r�K�jyx��Ȧ��*�7�+n�PŬ��K��6ʫӵޒ��Mz�Ь��S�#%ws��:��>�}��L:�	P��զD瞱ۧ��S�*��qP��ܔ�U���Mn*�M+��5k�U\ƨWJB����w)dP��۵:��X��f�y� ��<W,P�G<��O3#_$}kV��h��G�[�
����[8�Wy!t��2�
엖c�.�p�[�t��hT�{�,�N �����8����	.���R�#{�~����k���T����浳p�r��WS���Bz��/DX���	�~}]��?f�t�j�v&+�������y��� .� _ý�Tب����s��V�\�C�����9Ż4���л.,�`*^]���Z�b���̎��:m�7�5e�*}S�Z��:j�E��Ƒ�u�̮�6b�ǎkVN�����>�3����PԢ�Ba�O�Y°Ը��{f�U�:��g1��D8�����������v�P�Xׯ��[�������f�����T����P~ަ� ��Y�l��q��4*�b�Ys-<9Q�nW��`�Y�U��b�i��L��@���᜵vC��{�c����ކkf�}��	T9ą�k�B@���6q��&��Zi�����'�_5}��R�o��iʨ���.�B @y�^?l��������~V�^��C<ߖ)/p�{��Z���j#KH#x;N�[��G^2�s������x����pO�f,����u-��V*�\�+�ze�B��ݩ���7:�8ڒ^5��5,���U2ˣ��D}	gtw�(fV)�}g���VTjo.��_n�Kk�G,�aI�=WP� ��z"h��ͭ}Ȉ�>x�`�nO�[�f�*��L�s7w���z?S�+̙ꎤ������9[��*�w��϶����k���3;eڶuQ�[ݱ��m�в�8w의)D�sSx�<;1����㪙}�Z�I�|���q��7NW}a*�+���Bz�yZtx�0�2y���N\��Lu�+���|�1N����t�k�\wu�JK���f��x�N V+��e��U)��<���*�biJ0mD��~s<�����5�x��z
�fXo2���a�>j�@��AJ;-��N	�|Rt��h�2ىre�yQl:�9�����P�5���WX��
N��4T�v�y��:�7ճ�ho�?�J]��g˕����|&Mؽ��}�n��1�1�.e��� �sA��Pj�y$�eh����Y9|-���n�{9<mZ���+��b��S�M9Y��;x��EX�#��Iܣ�|JD�u�]4�`�Y5hsC2 9Ѵ�X1'�N��M �dS�5t�/y���.49�Ϥ31̩��X��4���hݚ�)�:��L^U�����X�=c��a�3��5��x�ھ����F�;���k�i��v��+�cf�b�����*,pU���V�*���l��`�U��aY�|�|X�cvX��
$DM��[mq���J���P��"ˮ����Ї X1�1�c�P}7�f�]^}��]i�Y��z�;�2�]O;�9<�.����
��g��5���YZ�l�u�U�C��C��z�����mMt��⹾��%\Y%,&�t��oR�P�ޅ�[󖒣�lw����˃��N.��5�˸v��;��+

5s_ۍSy|�����E[�X`JWy�RY�(_�9���ǆ�iM���@�]���Q� wp|Zu�,\�N�s��s��k����3��l��Ƅ2u-��+�7�VZ4��:�x�.�)N�ej��]�>��|�+��K��(�y�G9�PF�^a*�gB���ss�5c�ź-M�A�3��&�Ζ/��-�R�ɵ.��59�5�.YwX/o��tP m�٢�.���(�w3���Guv�S/u�syA6�v��i5������/��x��x�9×֯��\���-��o:ǜ�1Q��^弱qC*���C��֭q�:��wa��6 Z--���]Ӕ�׻Ro��m��jejZ4�è9s.�����=��G��r��tT��y����1�Ve��5���$.�{o�� D�on�l�)o=�ĆV.탑�]�HP��ٟw\>Ǒ-٧��1��v����U�bΫ��0K8ђu�}oT��ݥF�҄bU'?�k���tJ {�U�z9��&�cW.h�H�}j��)�b�P��'|���l��l9m�gvr�[l��&�2<���*��Usr(u	�JVA}��=IZ�-|��QJ��V9uF���M���G0`�u�l�ݘ�4쥴�W���]r�
�<��FZ���BfI�lQԨ�λ�yVP7t�h�ǛC��z��c6��HSw�kOB�.�i�m��;jQYFhS�NtQ��6	'u�����qv8̪ܘ"���u�����	4��~X�اm��{P��7�k���G�cm�p�YLaՌ뭚��N��\�6���v����j��$ÉZ�!�t�/�pV�8�f�S��2Ÿs$B����O[��B�77o��5Nt7�,Nʉ����]W�sg�7�ҲL`VN�ۭ�������,�����Krh�����������y�%8�����,�!!5J��i�w&.�%�k��m�������Uv������r���0����x�����x��\�w��߻a�ِ��]��e^�/`���ѯ+��|��dI�;�*�gu��]v�8�x��Ȣ*�$I4���F6����KB����`�5��-
W(��cSL2��"���1�����-B��YZ����(Um�+D�+c1ƥ�E"�*���YW)F,q,�.\�fR�b�	Vت���EL�EUQ�[�c���E�)�Ċ����iZ��C,�Ę"��UAW)TB��b�U��[J(�\ʢ
�)�bVV�UT�L�EF#��e�����E����\
#�UV(�b��"��\qb,��X�\lKeƢ(��*�mR���(�5��F)U����Dm��1L��X�����
"���\���e̹TAm�Z�Q�-��DQQ�$�`���X��U�F�W*��¶1jQUE+Q�(�4���V[(,c�Z��]��pS�edU�>z:��y�F��0��0�atv��ᡐ�3N�m��W��wN��]w@ެod������g\�I�sB��_5��H�����{���e.+�`���7���4�{���!t��RV>���X1����\[�\F�+yy:��z1h��b%*��]���i?1��V���<�^���S��`��}o!晪�䔨F&�뫜ڋ}U�����b��6�����3jtc��Q�sZ�m��睁��V`��%\�s���8�1G*�KʍM��������G��K���<��Fc?z!ԳA]�3�U�Ue�R�w��"^,b�(͝ջ/���i��[���v�ؔ�$v"n�E>R���Y�[#�f=At"l,R�ulg+�q�oiM����}��������.`�]5�M#n�.zT%���.�x������=�r�����Or�LEf�� ��R79���<���rnb
LU�yq���U)}��r��1N��u-�c:J1}ܮ7��f��k=E������T���G+���B�䨙���.l]e ��هWe�)�i���j�DR���٥��<���Wc��)��*8���$擘:�⹉��ӧ�:l�u���3kz�m'ϱ����h���������'W�G��=��U�2���C����B�Z�|�
��;U��t�z+����KA��T����9�I����󯚞7��Ol+���SqԞ�˘�f���l��5��:)���A�9U�����VNO|�7P�d�w �pxT�F��^b���.�pꊌ�9Ü�V[�S_kɍ�q/~MC�3���4]�J�j7ON��ö�=�=ͯ��j�f#��ު��45�)�niEQ��`ڤ�Z�����Ԝ����Y�^���j�]M�S�/Z`������ܾ���3�N ���u�qh\t�Gص(�Q�2b�B,,�5+�]WY�}���L�~�\5�\6���{��%���9Gi�1F-�Z{{X(��ǭ���
�i��;ͯ���}��`J����~�����a9�>��-�q͢��������ĥ6(�U� �������|��^t�]L�r�p�޲�����AK�DÝEm[jn�Zo2w:�"��3o'7�G7��ڈ��,�,[Y��/p_s:�ϰ�G]۫Uy:��Ϣu�􋢥GP�}�}�Fq��=t&^�պ{}���o,iU�Ȏy�dl%$���FP��ו��k���	�W�yX\��V�S��|�dS{_B��|l-��\Y�"��m�AV_;F��u��=���N.)�F�gM~}�nwr�}�^��;JM�4�+����`���1��a'��YRv`�¢�Yq���$�J�;��k�Ӥ��:�F5'�d�]IXv�^K�VG{H.w��M:LL�♼���u>}Z��si�n�[�1JQ�f����X�9�o/<Y���<|��&x�x�W$��h��,c��V�J,��[�:�Z����.U3�nH�j
�@r!�t�f��
���7��P�T�rwV��I#�-[ݵ���w�Z�>�-*���,sQz��ޠ�9�W7�L�;c�������tDx�yC_o�l��<�<�q`9��o]��!��tqћ1:	�Q�O~�y��⑴�\��p#���n=73%` ����妙�ȥ\�$oT��.֙�+�F�	��À�۔����+kiثI��y�\���m����Hj�"ݝ�PEH�J�Nx�&��;uwۉ,m.�kOGN��}��G�k
:�Ed����U��Yg�z7ױy��'1x��i,�sBoJ���rU�w\5:��{UCܩ���F���z�߂�ϊ=~��!^$7�엸%� ���Ew,|2ި}}8��5�u�W�*�0pM��S�&v^槫-��V8����^ꊾX�[}�����Y�4M���n�N��:
؉��.���C6�՜V�iY_jo.�۟;ݨ�kV.��T�� ����y�N��q놦��kUg�Y|��S��>�������k�٧-��jb�Z��;��y7����a�r��w���ϫɬ��{�7u-����зn{_)���6�b�U�[rn`��w5/N��UMU=�sVqOC��/Ww+rҸq�*Ӎ�r��K|z|+y|.�]#�kzm�q�#���r�R��J��.wx��V�p��W�2~�H�'.Uᆮ>�q�uP���~-�0]�8��y� R�Q1,�Q[�wI2�����9������SH�U>�� ���
4nj�j�pVi�Z����P|�cx�n�`	���N���u�����t��ы�e&�ާ���=��J�[��ߺ������^\:7P�P�Tߢ%L�N�.̿�'1��Osy�;�5����cg�L	ؚ�r�ֆn�w��&�[�p̅Y�æ����&Fe��o�ݻ��K󾛄�6R��S�=�)�����ʫ��JVks�����تx�4����.z�{��P�A{WA����p_m]W����\�J��Je_�������{S��t�Z�����:9�]���#��m[�U[h�(�����Z��OSu�C��O^�\7��Ck\��5Ϯ��a�4�j�Z��S]�������ڠ�u(��x��#�s&��P�V5T��ȷ�ϑI^w�*+B�qq釨�z����ڜ|���>@D��x	�M��99���h&��9c���8�c�Qʢ4���7gU3I^ͩ`e��
G~9����-���7'%}���u�Z�ʈ]�zs��7^dK���[5�EL���A��ed�8�efZ��(̹��Z�$�ouLǊ���=�Y�$wGVJ�:PY��X�8̓+X&m�lp(����.�B�G�n��#]%� [��p`��1%Ý�e:t��3��}�����ڌk�p��~����{[`�|�g=oe�J܆�aOv[x\=�H�Gb&���B���w#{Q[�ZHM��l�+�j�jy��&��M�u��êEB�-�apk�9lY�m��:�l�"�8W�1K���]4�P��q�m���k�-�iH��<��Շ��������<����t���.�H���=�Jyz����r�p��sg_lVxW�6:��_j��zd'��w��Vꨅ:�P�g�V"ڬͅ{ݓ�J��Cq���bUʘ���rʉ�ek��!U�z��d�<i�N<�g�2%9.K�^�nt���O��1_t��YQ��]��ֱ��"59��h�k���s�:��6=�NC�n'���pe��W������'�}��;�yEٴ���9ɋ��M��E8T@ul�2�t����;�Y���)�T{_?;���q>4ԇ�46��ǿ\jn�,#WۺrD���2�7�w&���[�N��ք�X�#���	2�/`���)QjI`�i�!�l,GH�Eb�7�M�h8��V�b8��Z-g6�OF��Sw0's�����>��-��.�u4@�[t���>L��U���4����DGսm��rzD��}���Z����+� ��
پ�N���^*�ucq-���WzY�OT�Y�Y�V���qӊmbߗR�����j
��F�����u>��b�{�o���C~�m����EQ_:��P=M�4�����NGi��i�/�әoy
����<\��y�0%_�u˾�P�!�_]oQ���U󍕍���i[Z����}�󷴦�-<=ֶ����yg��3E������^ƓC�f��w�}g�}es��j��{��7��70��Wg]J��o��B����)�:
��˅�;�_�O�����W�Wu�b�ەe8�43�e%�{��f���[����B]�[rn`�­5�����h�d����A��[<�V'�COF[+�t���S��H�����T!�ѭ�Y�^.�Wz��e��_\7��c�V�FE$9��^�+:��B��؍���	�e�zw�/�k�5� �����$��.�	��천�f�͵W-������i���K�c�|���ݒ7!����b[5k۰(c[���]۹*��(5�
=��Vl_d|��1 q���fu�49Z���'RP��Stq�_}B�v���ŋ��e��;u�)�W�8�6��wP�1'�wW��3���=c�u(�Z�byd�Y��W1�:����*\B���O!���&�Ont)gvn�M�e=�k*�9��c9�Փ}a\&&~MCmf�t��ՕknZY�Վ]��D��6_m}_^b��f1`3����A�=7�{��y}���܍q��mD58У?��A����T^c���Z����9B��մD��׻�3Y=Z�>���S8����ܯ��ʃ��-�e��'2�e�C�L)��dc����uӊ�z�c[���j1�ʆ�nۑy�]'e񽰪�05N[]{��U;����-/�+g<_w���=��3��[�U������
�]��*�8�-�-
�7n�۟;ݼ�J*T����go����k����Ī�*�q���j�����ѪUF��hpն��ݓRW[��[���fJ�nr�ٵao�kl�����݀����ZW���q����2�]z�:Tz��J�wu�rɥvm�^�ϩF�"��U<����Iǭb�B�i��R��v楷�.s|	���q��G�Umq����ܿ���^�E�l=�V�Իj�[�׋��\�Bۉ�3��S���O$.��v]힦vU��g�=O'#R���y�����5��+ë��r�u` ���:�v���qg3\��t��N�:i�z�o��-�v:ܫ�%
�f�0κ��b-�M4�S7��������^�P��a�8F%�5�K���sq�������&:���Ň��u�����Ju�6���vl>x�V����$����]Ä�[fO�\J��	�_�\�0�h����^4I�g�-{ř퉡�5��t:�1�%�U�	�vX�B��MMZe�������4*����_#p�32��O��.�>bB�:GVx�xr�Mod���B�q���B�M}��\m��ⷷڇ�ʺ��!�AM�������b�m�����;���RTcCjƝo����K�H���*'|+e�^��hJ�TL�-�]�{aԿ�q}�%�f���L��w�.oS��kU���b��5�wC�C_�$H'[af�5ț;��(a��^�0i֫��I�YT��tç@�CQxqw=�Lɔ%�����a��q!���.#iõ������.Ã1v5W�o^����1YǨ�痨�>}���v	s��V��2�${�=���}��誁*�j��}7WR���,���g/<9�V<�/WXă2��XM��j^��K��y��U�\⯈^�]S��#�vp�o��ޞ�Bݎ�7�Q-������*�����ֲ�$#k����R�p�|�QZҞ����	��!���MvM�p��ĪS|���>K
����J���T8iu�ˣU��c��ɸ՗ˠh[P�ð��[¬�:�U��9в���A��i�Sx�b�*�˺�>��d�M�X��Iߤ�N�=�qG�d}�k��#��O"�eC'�=�~�/,��E�N��s�����Pw�J����H���m���TA���^��r��]uf��¿��U�+*c>������Z��>�q�Wz�&����P���u5(����I��������[�7��mj� �p�mR�����J��:�t��`��Y9Lx�6�Z<�q
D���cs��]�Gm7� ���`�s����|Em�Ѹ`�)Ȣ�N}�8Gy�g��]�pxw���eߍ-]=p+��Dǆ���(�wh����N8�t��}v�ϡ�T�l����t����F��^���l7�=d��'"�8�8��O	��*��5^���6&\T-�颸ѬY�tiwGv���ե��;�C��9��M��f+ŴJG����w�q�'R�;�s��9�J����YMY�y�sLS�K��zG����y�c9�B�^wu�{ŧv�8((�$�Ւ���#�Y*�e�r�#(�,pAWI��VF�S��9�P�t.��P�;*8�)��7���vl�����I��utU�	IeN������tm4���i���	��A��ft����kM>Ee�}��t3�3M�R��hS�vK�W�\��婹}
Sк�h+��I*wa�/�f|��Ewgu�N5��7)�{Z�A�8ёA�nh�Ó�\sR�t�A�
Sr묀\v�5ۃ�q;����U�"�Ҏ�ٯ2�j;����Ү���Q4P�ӹEu���i�h��T�T'�X����߷�-ǻ���݌|o)�8e��z�C�D{��h�4GQ��%Ese�"qtU�����,�S�Vvᐬ����xF�А�Ʌ�Wvs�s��Jʜ1�e�\���,�brJ�<�@dLh|:p��Ƹ ���.������s�]B;�[�}[�����<phl��=8��ͤ��C�qb*�R��I���8���
\k{)h���6tV.�����Y��CnS%�u�b�F��B
FVtԧ^o��0|�y-wI���;�W��a9����Z1�ݕ���!u*MΫws���SB��E���`t����w�������v.�8���:����/z�ω.c��1�4Q&۸���ڥ�I������-ej�Ary\����%BaB�͚�ި�mG����Sۤ�n�k��Ҝ���w���鬽8:�ܚ8r��&�л25&���g&��v�tɒ-�8m��k��_�ESx��on�� ��v��(Bҕ��f�������o�f�|�z���n���]�}�td�{s�#u֦��z�t�|(�\[��䷱
��x�r�u�aG�\gw��%�"(�1��#r�$E_E����l"�A�w]yz+���)��i�tg(�,3m#��J�R\�LsC�����Ú���j�3�����S�U��'f���M�j�q1��N{�.=�.u���ǝМ�:��Zyt�wU�q[:����BZxč\��X��gc���a�ŉ5���c��Xq�=c���+.6��"Yt�1�u̫'i��E���=V$�f��v$F�a��u=k/7Z�M�_*�z��d��� !qP��^n��y�g�����F"*ň)�*��c1��V-�TDq�%�UQTAJ�Z㍥Rۖʖ\J���*���k�D*X"*"�F"���Kj	Z�(�%�b�s+�U(�Ŋ��Rő����.\p��`�V""��r�Re�ȵq(����"�)e[\�,Pi@��"(�D[eDq������["*�*���h��V%h�Q����T+X�4���U`���Q+`��eb�0DQs-�0TX-�A��(���Q�����1EE[[R��QX�B�`�*T���"��mDQ���`��)H�-E+%�*�˘�,�J�J%`�L��(��U���b�h1�dQP�Ղ�mDR�,b�TUQPU��X�5*c,TPkAa�L��F*,ڥ��bł8��\YDX(
\sIEUEL�b��B�-�Z����UJ�,�k]g�,<�uu^B���f'ۙr���X��n�uN8�W�wF9mw63�����/8��3�s�X���E�r����}�e��Ұ��M�K��)[����=���l���f�U�"�dS��w��bb�-c��ke��ݰ�w�*�'N�P��NC�n&9۞e��.Qx�Ƴ�cL�\�er�x�ޙ�x�^N����i�k �t f��{�o	�i�w �-,쨼�W�j#V�1��T�#T��̩��:ę��jo�s����67}.ᾨP\O�?�Ŵ��oϨV���홶6e�y����97��J�)�7��_x���mx\*�.:qC�U.��[�s��;&�a��R՝�/���?S�����v��~�/՜r�.o �Cs]�����wr�.�֑Fad������Qzд��|�5���}��������]\�<��[�Ț��X�&�4�OP��ڰv=R�^��k}���w��w{£;��Z�9]{�� ��/��m��H��GO�V� jyq��숦��ma�i��X8hH��1X��I�F�i^�$�.��(�;lr�B�f+�A�/��SY�G��*���D�ο��U� �`�AZ:��g�Z��S�5��{�������H����Vt�KPQ�,6�؋mRxf�-Κ{����#���A�=kJ��Q�s�3=�Q)�������w��K�\6���GS�a�}#�n?�'Q��Wc�C*��;���#T�!Uw=%{[�'$繦��j��%p�W�����OI��}�5��e'�&}��zw"�:Z���8�Q�����1l@��fx�ޟ�������AM�a<��v�S��!c���[�1JY�y�s�h�
��l;c��A�Ɉ��'"1�ۏ����jK�i�y
�R��uW5�ξ���*���:�Kܼ
i�ŎwVO��jb�%�fW�Ns�V��o�
���m8�-[*n>ۃo/-l^31�����0欿$��������ւ^�����7�Ob�7��v=��ʼ�xn<s��=�UFv��W����呪u��[�9��y��mh�E�q��NE	�e�4fdi�F��L+S�b0��:�V�Pu3/A�du�� ;	Z��Euǜ���S��{%��h#��js\t�г�X�GH�Υ�Y�G�o�#,�Y�(��;��]*ú���*�+#��ŝ����t�r�WQ'���1�Ŏ�������롮����y��yz�7��_�}B�ک<�-W���¯}=f�����{��܇Y�*z���z|�WR���-����u���������b��zi��ۼ�of�^�X���Ut�ո�]Ҷ���y���3"T+�<&ڜ��k5r�t;N�sk_�Q��O�ڰ\�����'���n���yܽ�b?>W���%T)P�����S�s3-�kZU[�;���p�u}��ݧ����SM����^5+��d��O^��^��^J�:7���t�<m4���یq��7c�ʼ0�P�2ط�+�eaqr���N��݅���][�aK�� ��t�^L��0��ŃZ��ɷ�5��9a����ƺ���c���ܼa<�=�p�(bc�5��?V�1Q�5�a��pg4�����=~�tVVִ��*�qjt1���z�ʳ����ͺ�����PϻαnV6�0J�c��<s�-��v�t�%��7�>��
�Ǌ��=�'�m�v��1��u(^X���T�<�)�T��PB�O����;k�<}.���v&o�B��paV9�!vlYVÚ�8�泬doK��9U��u�wwf��CyI�z��h���:�>�����\$�����[��Bs�Q�z.�g��Q~M@�fޣ�L>�7�.s:��ȅ
��OoS}�x�u�3���[x��ث���ɍ�28�q�HO:ح�gjGsn�Ei�<�h�K���lޭ�<�^�����a'ʣ�o3_/�Ldϟ`����~�yPq]Z�s��}W瞫Yy����W�쑁c��>�g�3�T��jt[T���6ӡ�����D/j���0v 5�IN�G���q�x<Os�w��,��:�`H+�ۛB�_��\��fA0��9��k����T��kx�&�ñ�����CȞ�I�'sI����Řs�	d:�v>�j����m�oiM�Y[C&���]�0B�G�>���n�wD���Պ��5�@��>[����WX�pah`�#U��V��`.���\���3�~����퐹Y8��7�
g^/9E�w*���u�w������ͫ�ɋt��N�H�.��ں�z��i���#;�+����aF��{��/(b�\�}��z�l��+�T>y�'Hz��{��T��u2�9W��<PUK���q�v��rR�V���.�ԋݥ7<o�X��M�w��Y�It[��F��*�%P#�T����@]�x��[Vl*V��%Z�Nrx�V�)�.�#�&T@���'����o	u��M�T]�u;8�ޥϾ�=N�z�uBxU�1�!v�Xl������['�7/���b��׻a��oPT��q�T5�r���7bx9|�i@�Y�qÙpn��j���6�-�Ŏq�}�AT.��P��L�Όҝg:�+��i�X�n�H��j�^=�Z�f��^F�ڎ�Q+`��ˊ���i����/�LW�=S(⺋x��'��W�`ju9-��L�X�	g�;���F���\kC��f��[=V���E�8��}�W�(r�aoxU�cԖ�*�!@���g��:���l�S&�x�|.����C\��Z��x	۬gt;O�.vH��U�P�o+���Wܬ�Z�'2��Hj#�.�,9�-�4�#^M�P,�_j��r�������~IK�꾆�>C�U7���<��)޿ﾪ����Os���ܨ�V�[z�_Mcõ�OOvA�P�>&΃�z�Ԓ��u6J3�y���b��GWs���a��}��`K�e{iA�f�Ց��o]L�s�	���,��w�V֦��z���z�u����S
�����x��)gAN �H���u��ʬ�z�p���5��8����A�<� �{����}�͇��J�R�m�ĥO���WV�F>�{<o-ׂ��M���/��]���{YݖА�:T*�j��*{��t�{���=03��P=V�c���ү���^(���%7�l����YQ'�������pe��.�#r����x��uTB�}7�8���M)G��a��"�r��x8O��f*mĠb'S��,'1���OT��:��U~7�#p>���S�{�j�T�=���^
1��;)�[�_b{��0��n!�z���1�ՃT�h�{��W���f\fN�v�� ���b�1��Й�����W��E4�&�6����w?)\V>8O���ե�CU`)O>�7ܲ�'��E��_˺n�u����e�h�����=.�Q��2���Y�J�N��`te(J�1h5}J9N�P��W���j��+!zȘW}��L���-����%�ٯ�9�SO�%��q��X�r{[N���7���F�2���h�\�YhGh���{�������Q�4(�G�BYg�{g}��^c�^� u�<kg�nu�����7qʹ�GJ�o&^���z�D����5]��aq_�}�ĺ���C�['���z'�g٫�"!Z_|���䚘���J�������>�{U�A�yF�T��$���v�s�mX�%+��w��P���j�ya��}��U�JϬ�q�B���$[�0cmZ�[Ĵ=�ō^�CV���녱(*C�&�ֵVyTY|�F=�c{��(��o_.�Ʋw�'ݑ��+��ȅas�fS�z�T��R��h��N�Z�����o9.�+��C�m�B�n�����׏Wf�
2�s00�mI��Vq��H�b��c���}��Th�ӟݓ��.��2n��7;	�8�wiչ�tv.��5�5
�����Q��')xm����ʼ�ǟA�h��C��}e-^���6G@I�N�:8��:t��]�3{����]\lYڥ�m`����G.z\�ѩ�j�sbisSq��=i�q��]�k�e��'g�@�:9�OU��4���TB���ہ��	��x��+[��Hk�r��Va����A\��ƚ�}�ч��W�a*�������2��T�[=���;A�\�*���-�\��a�a��Q��a��_τ�˄��+��^�I���s/V��J�>j�����7M�+�1�!v�ƖT[b�](r��TJ��r��]kt8��ەs�e���1)�m�¡׻���/�����?[玴5��hY�p�|�m���~�9ޠ��5y�hY��:�T˙�滗�C��Ã��৕y���k�qE�u6uHq����qQ��Ɋ5��kjN����#��Eb]�>���'��&F���v╮��������V����}�V��~8���ݥԽ��Ks$��~|鵃ju6��yv�7Mf�%ǽ�NA(
z�,\����r��qgm^m�b�r��[�{ѭ��f�Nȓp	�O�.�H̆�gv]#]oG'6�f?�)��ג�$֩3S��%ty��e-BO��m�ö�4�\{�}�g>o7����k䕶G��k8�]�D/a�O1��r���31[(��N4�kLu��q�mD7km�����\MC�bS��2\;w9�z��:��/���ӸM5�󷨪Y�1���]ζ�'MnΦ�Ͷ�vm�7'6)��+��rɣ�����Rkx�6�I�(�"�.����.Y�a]�k[�m����k�����]���녊���`nMOܮN⫝̸+�V���5�߻%̨{rnJ\+�\�v^�M
��!���ԫ���+{���;:��y�r��a��rʓ	���,'��T�X��ոX�t�p�Gt7�-؉�h�0���YS�b����wm�����g'�2�+����W:�2��U��ו:�;�*L$6{n�*�X���R+W<�kݰ�cz���'N�P��NC�n:X�>��yr�Įʅ�Q�5`��Z5�f�{�@��8с刹:amZl����g[�G(���jxq� ���ŷ�yY�ϡ���B��3e��&��k�(u6������ig��:��J���K��X3���[��[�f:	Zj���h��ӎ��<�@������4���w��ZR���/f�_�Ԛ;`>�=���x���V����k�x*ʛ~�;�ٷ�y��֭q4��[�z�끇�����iu���Wr6��kFޣf��a�^A�u�TE��'����%>/^��,��5^�����z�>}��F��z������~�
��82���5�^�#�rJ������9K(�Vl��y9^�f���m�C�TU�f{'&�l����2�F����赁�gC�!����ڈk�u��Fvܰ3hV;��R��x|Wõ��B�~�)�{O��|��t󠇴	q���ǽ5��`3��8.���J
����X�AkQ��@��M��ks�O��]��4��ս)��ݭ��8�
l���i�W+��p�g@�0j�@��9��Z��1C�kj�w��q��T-�70R��!�]B��r��G=�4�f��z�wj��oa�������i�W�]a�/c���[��%���Nᝰ��swG6�Ձ;��p }䲕Z�=���H]��Zl�Y�ց�em�N�Rnq�b�@����|�] B�h�qЍ�!�.˄V>��u�a�C�rε�2<��#uu���]�Ob{H���u�/r�'WP;)ɍ7W �*���feZ4�t��t�Xwy�'�[�C7��Gl@��;V����or����X�r�s;�`�͘&je���+��^`��%���jF��љ����3{�IgU����V�㮞�Pm$� ���ŝ��ϑ�hҫ��Lx9c{����y��X�/����kD�c�o�г�0֫RP�d��)�d]�k��с��p���q5�����Iu�v�=���n�
x'E��ulL��Xi%��
Z���]�-Ƕ(u=d�j�V)m�����l��Kw��|*��*_A�],���	�l��u�s-]�c�L�����u>���T�V*qtL�Lvw
��:��һh?��	�Nn�
,<�j�\�h6Oy �qv1x}j���N�{�"w�-�k4�Fm�{4�c�1�V��Q�z�7�*0�x���xns� ̝��D	}����r�2`
9��s�ä=������wW�I���[���V�R�״�f�Ԝ�H��}ۭ��h=ǚ2Ĩb�/i�A�N�˰��J�������j���;h��.jω"��t��c�0X�x��^����	�S9]�|�M�� �N�6�C��=��R�2� vu��T֬�o�s�#y�>z�4���˼���]n�{.YDvҫ���M������2�Y�sm�'eO�I�yf�a��N����vl��νd���GP�n�V���;�m�����bo�NH�}��[��.����0���gO��8��������]I�;)媍�[zx�3���(��-ܳ���zFj��4���-쭘�6�v0P.	Y:�J&Q���er�@)�D�h�n�UY�k�BE�򻿙���ː	�V��nC���ui9�4_;+Y�9�L������q,���^�՗�����-ҧBLu�A��gv3��n�M_9��l�c2���==r�#R`ꕻeh�@nJ�*�9�D�v�I��xT{��/*�X���̊����6�Db���-�-6�ڒ"B��3"�-H���A��KNy�1�7�GU�A���m�|8�����H���+�:��^���5���nٶ�]w����Z��'��W����[\8u��;��3)d�;�q�r��F�6�N�'�������u)/�f1$R]��K��'��R*�w.�k1��M	T�pX�����I� kؐ5�6:ЗS�Z��Ȼ`�I�CwE�܅n�:ke����o��إ�{�}�E�Y��ځ䣘d��^v�Z��DAX�{�f.�)���
�%=؎��*8�RN�Ѭ8��Q�Okza���G�:��P�������X�U�*
*V�QA`���"(��-�ڒ���Y�0X�l�9@��q�,X��Vt�uh,���
�"-�DEQb"�12"��B���KZ
�%B�9eAb�#1)B�TPX�UE�X(,�QTb�Kj5�R���V�Ab�d���ӈ&P���[�R��֢*)mT�EfeX[Q�H��U+KJ�����b������PQTTX+XV,��eJ�X�Q1AFڑV6�����JȲ*�cYAJ�"*b� ���4�m�(��J����UE�V*�"��Ud�mդ1����U"��U%dS1X�bB�ڣmE[B�2ڌ++Z"�i���"2*�T���im�*�j(T��Z�PGMT�M8��*��� ���qy��[O\�g"������wc�� �q0,�Ջ��[���k���^���WX�����JYPz����}�K��<��[��ݐ�ƻ�Tc�k^Ӥ��nVJDjG��ag��H��ζD���^�W��&����n�u�|��W�8�n����#Y��Ua(�ݚ����t�ܖ>�>F�%]藔B��Y��:�p�CvUԭ�is��v�8.e����0enMb{��#y�M����T������YQ��$q�Ө�Ad*�q?+�1��i��x�S�1��F��nL�Q=��l�Uܻ7�T9�B��ơ�-�#�-[*D�͈6�1^3W�2s,�Y�tw�b?GF����|OjC��j�78У9��Ж\y���a�ul��)�j�����1���|�A�������ەJ�Tk��#S{�FN��I��J�o��V-]K�A�eE�[���o�{\ϳ�FT7�^���G����F+�5]�T9�.�纺�m1�՟l��w�\螤�p�Z�~k�{
WbWj;lJ�غO���\���^TepZ�Ҭ���u����jU�(�;�`�p���$��L��u�U�c�ч�c�o�r��D�ٝ��v�!n�-��2�k�œ� �2��8�����u|r���O)������6;�G`�=Q��NׁT�/���!�o�q� ����ܕ^J��J��Fo^T�c����y&���"��`*�*M�N�v�&�܊�1��_��u�ؕEZq5+Z�<�	i�������mOW�S�M>�O:�d�j���%#гbn.������5����he(]��,��Ux;�����hz��}��q)�{��,��qNȡ d-���dPV�e�}����~7�U#+��~���6�U���x\y��މH��F����<|�}/�ܣ9����O����pJ��!�^�� ���6��ܾ�ſJF�>���j~���3����]̟C���F}��C�2<���ٸ�SB�������@�~+�a��b1��ҋ��|t��;%���^��Ȩ�T��>,/����g���/�t�X�
��}W�ټ���R]�p�1�.?;�7�����׶�y���3�bH� 6v���I5�+�������td%�9E>2=�g��V.s�S��yNK���n��<�ITs��=�`�:�d�.uvȻdQ��1)�e���*3�oJ�1��e5v[�SW��[��e�$�җ�kZ{��{��:u�uZ����l��+2f.j�^8`�s�<�Ʊi�/��:Cseq�F��d���K�m�q�9�6��}_t�aoh�LY��}����I�p[Lz�U���V}����M�,��9RĊO`J�u�+�ބ���}�����ꅷ��cכ^�}��f��R�_�9����<�'�5�+O�Sac�ߝ���޳^BO��t��v���T;�ڭ7����u0�Z�`L�5p_��Ӿ�f�Ԉ�B�)��n��66#����83M�;,e�V�+��+��,���TB�Q�B��=�Q�������������|z�=�F��\U���|/����9>��VU1��d֗p��B�{óX��R&<�&<�B��)��z�
�S���N�^Ǒ����%�[�Nh����� ��R�jl�08�(Y8���_�鐣O��~S�w���uj�s��>0�g>O˥Z������F�r=V}�9��3`eOx�Q�3q�,/g;�Ŕ������{!��9�}�~k�hS*�8��+;����p9�z�;�8�c`{�n���J�u�Pѫ��8NR4�c.P�!Js��ڔ���{�������r�/A���,t�Rݠo%��ͨh�U��5�ǖn$P���v��C.'*'2�=`�k��W��F*�3�In�K���u�jiUѝ��A-�g���Q/2ܧ�K#����@���P����e����%�u}Eobi��j�w{���7��zz��F�b�����	딂�Wݪ!�ZF+�w��>�2���R��w���J�8������W�w!�g�Z�2d@L��g�?�:Wx5i�T������'�2��B��E�T7=^�GӼJ>�Z�e�O*�<���`����~Odg�H���a��d�\�:0����Xʄ�h{#�J�1��O�>�8_{n2��ר��8��R^�ԸyƏ+9麍ی�LLW�m�O�vi�6�U����׍ßP�N*��w�{$\�_p�ŋ*�FFˁ'۞5�n"j�;����+tü�t��K�꿺�4W+��US�g�Y�S1"�NW����xȟg�^�`�o~��x.�3��n#7j�׸���F�?UA��T��
=#|�S�eN{G���\F����Uh�3�6o�IG��~��2�3ա�N���8>���"}��kS<4[�������^�ۊ��҇��=>�Co��c3|v�	�	=�ݾ�آ�����Zo}#T�`f��/������W��j�w�Y~�lYl@w��}���L�%�CW��ʈɭ>�L�7�@��G���ZU�>�eh����C�Ƕ1���������Myw.��U�4:G��J�튁v�S����YKEU��NڷQ�<}��dR0�l S��Py2^�7�t���y��U�K��iv�y��A�cNTݏ;�i��/%�Na��#��r����
)�S�,�ҕ+Ń^ts�o&�Q�j�^�>9������L�73��GT�:㟯�|��#އ��;���v�a��\����;��ވ{H�ҧrf(��\;�2��ɖ�sʇ�;:��Hط��u�W���2�z�4(�X��nK;�{�;��`>��`M7p+��rܭ�(ⶡ�۾YW��1��Wy�E}���謹���Ы�Vʀg���yU#��gKדY
x��#�z|��zX�iaV���#��
�9�k�����=��,f�Ke%��pd�x-� |�^(f=b��U!������x�Fς�����+^,o��H���/�pA�(��O�ĨyV{Vl����\_��N��{6*�1O��t���|%�#�|:!�U��v�
�N��3i_���Y��)K���辤n�*+��L��߁��}[F���0��G/
𼶗�{���������ʟwGک�cӀ�΀w�@b��f�q�D;���K��5<��q�,@ݾ�T�yws�>N�C���f��=�:���2@��:�/2ׂ㓓ṳ��`�^Y\?b�E�T"�'������VƬֳ�龘1nnWoP<ۛ���>�ն�jC9^���@V�5�Ǻ�����u.w>���p�γVo�<�~�=�N�z�ܓl	�e��)�����d����%�<���wAE�;X��iJ�������'�zX�3�|,��_:����N��w��{|r�G��/I�xｽ^2�쪻�A�O���J��'Ei�=L	�~���;끾�z_�j�\{�gLu�i�$���%ޫ���_7�&�����#M�U��iCћ5��\����`Oڶ�2!{k�{��o�:��S�Xء�ZkE��'�<	ʷk�mR׵�K��S�]�L�/� �x�����z�Q��n3u�����4�tw����Z)�{�Y�V�*d1{�����n0�e��<�W�ҽ]�x���wp�C}kNG���c�ƾ^n�g��Ac���]``��>���(ޚAq4��L�r���LyL���9��9�~����O��:�q��<��Pͺt�O�S=��p::�L�^�_�dQ||?Dd��U��8�GFk�Wq�?Q����z�1ͫrF�dbM�|���>���UHʉ���x���anz�x(��1���w�����H��{��ۏf�ٵ���h���5��#�n	�o�T�RÐKGّ�U�qaϥ"~���F ��ôx�����;V6�
�B5p���������P��I��o)�&osA�%��
>�qTY�6�beѝ<G���;«z������).�<y��me.6%�m��	�۽�rf<ȝ,u�oGV�$�U�C�uzM�SN�n�a�9�Ft����{\��b�%۪�����`h��~��^���dy�� '�qJhT��9�-�ǰy��Y-�}�F�˾G�l�g;]+�C���w�-�/z� ���e�_[�rE��Gŋ�0|2�j��s�u�uA�&��$��5����6*=o�����3�8�(~�����B�!��t��j�95�o}]w��+kΗ^!z==�"�N��</�X�o�{�c!��'��=��^y^���X�`������P_��)#��g�6��v1�󪝤�C�����顾��s��w�g� ��8�e�.�2} ����JG�L<ﲷL;ͯq���3_m0U���n�|A�"�R�G�sU��ٜ��BuBE}�������b����k���i�6��@!51�-ǩH����ɥ9�1��#��LJ7�ۡq�h�������d^K��y+��毬׿0����V�f�䵐&�������
��狯?\y.���/m�.����t2��8{�=%^mY�r�8�>=���)��HNo�2=�׳��z�����~�;��-��ӄ�}�%ʌ�*�SC*��z�j��9�T�ߡLk�O��l�B��U�ݝζ;!>�zQ�X�+K3�L��&�{�SV����N�9`t�q\�J�7	�xs�{6�3��0G���A�=�*�vW d�����	�acf�ZG;:��;J'�-�Ĵm��W������υ�γdϑy2|7���ly:��mϼi��d7��A��}�|���ɇ�����"$�.n�����@���n#&X^�vX�X=�#ۢϹ���A�����o�g�����}q����7�`>3>��Ex�Q�����G�.}����4�.�_r;OQ��hW�]�ѡz�^M�e�	���ޜ�22�[��KG�����^u~Ux1��po�O�4�z��]$W��S;�8:/��@����]ƙ�f3�2!!�N�{q�`Ǯ*�����<����l�ƾ����#�4�.#��8�#M�K��#*�P*��9���n4&=�w�L���W����Zwc�!��W�����
߶�a��F���Vg{a�Y�w�� z6��g�un2�11MVѽs�ݐ%���xK�5�~�Cޗ��EEA�W�9��q��N��@�qˀ9�H��=M�>���0�=]'C��������c�8��߷�\����������R�9���^bJ9q��]�g��n�;�6����fJy_��\��	��t�d�o:�)8�-s���ԓV�� Y3�Rȶ�9[��׌Ǩ�>���3����h��#pU��k�Oe�����R6�%#r��Z�k)'q��V^�q��sP�w��5vٕw��B� R[�2+��)��������t�;�V�Ec�ξ��9�}�U�h�/e�����x׽TǱ�5c�����Zn'e���hv�~���ژ�����fO���3����ϛ��3��G�v���M��Ӡ�
�U�\��r͋���g.��489�/�b�+Mƹ�,���Z�g�������*���\��0�`Uuo�7��J��z��8u��^Y5��ɝ�r��=��lV�{���Z:,@��l���{&����%W����������M��};����=��]1dγ��'�C㟯�f��s�=o�u�foٯ+�����e!�w���f�	�r�%��&�����\<3d��=7��xy3�~����Q\���/Ez|��q��>�[.!V+�ϔ�{>�z��e���~��xzuË�$��xr���vo�C��}P㜤V�+�o���_��+�e��2f����ޚ��&�F��z�|�+���<��e�Q����7���dA���w�F��n�`�S��ab�V)'۞0����<c�G�8̐�e2��r�s"6|}���C��2=�\��@�;Pg9�IV��n�K]B�v���PZ�S�ems҇�0�cl�ir�����+S��*ˢ���ծ\��K�߶����Ɔgij���/��9��R���,C4$�s��Z�5��]�ݵ#|7�������.eA��`�4l�/��CU(U�3�`z7tT+�lك���"b~���8KGw K�S�|-�W�^���H��8��og�m
�p/�@u�;J���W��=!��@xW��11O�hޗ�ݟ	��F�S9��쎾��k�t�y/:��.��ϋ� '�6g���U� �76H}~���
{�,�/۸Y^�^��Oq�j�G�!z���^��(�:��~���.�O�#���4���ɡ�f�s���bx����CL�i��}�3!�:���:{�z�G�ʛ7��!���P��FevG��YPm����o't���Zw���m0&�g�<6��@ϺV��yu�wӖK�Y������h>(Ǣ0k�r$��N�{2}Ņ�Zn5�뎦�,�d���#��a��{%O�8�_���w������i����FYUFV�;�WY��r��᪞k�O�Nz��^������n�.S�G��C7$���CJ���Tb��q�;����jÙ���R)j�񀴢xc�O���Wo���/c��!_C��sa��}�5��<�=�Ll�#��;�\��UfC�L�]��ۦ��x�EX8��\aT��'1j�����Bibp����]3;7��U�x�ҷ�eꥁ�*��-�
�+���h���K�)HgVǗ���FS�s����>�$;28���)�Q�.�yۥ����U�t=R�CN�=�d"�z��}�7����Ih�q�x�-�0Q���%��J��L��g+*�%u��AҖg=���sWrȖ�[��,�L��iC�˓Nǅ壺��3Ub�oC�>W�@	��nVG����pt8�Dr�O�o<�)Ʈ ���R�u�]��$�2v�@�`���
'�v��C��:�5/>t��^,&�9[f)+��RP���[�o�ʵ:��e�%q���J�=��>�Q�jw�-�v9p1�����	E�r�慺��i����crX�#�Gth$�x�e��)���4�:�ք����b�~;p1I���3�c���]��̬m�rgt���`<��u�
c.�+h�Y�{-ѡNX��D5]�޹������MN�r܎j��d��x9̶��U��A��4ew-�#׷�u3}Q��^�/tT]h����=���n�8��;m�Θ�'O�v #z����6�@�_m�'�@س�/����E�b�'����yWw��}��Y݆�k`s1k���AV���z�{�]8���ɮG������
�n�ܻa.r��u�.W�'��ʍ���y[Q7	���0NG)�I�Z�x�AyYv��*���t��f��y0,]ݔ���q��wL�ƌ���ܸ���x��<m,�kn�F�Y�X7��'�����\� ��Y�7nQU���h!T�l�)䡔h�u�b
��īmW�k2�ò���t;�B���i�؉��ô=�Dۉ)K��g��p����=�rb� �VG�-�d��#c-��m�u��u�uʒ�9u]���S��r��q����v i��'��U۩�����i^a���0�4EyטE�� 3��w#H��.����;���BR_h,SF>d�a��y�R��|L"�u�_&v��O`R�bz�!c��tb��jǁ�u4v�*�㔝��V�ʝ�( �]��81�������6��NbmIƗm��T��*��H$�j %�g.Vpe��-��/5-ם���%��9X708sCq��-`��0oIh��©�1Ԛ�l6 cxʮ�R4����T�3��Wn���h=�қ�-�C��ʛ�m�7k w�Je�^� X֙Ќ�"�K�Wjg � �߳��
�ƻ�ݾ��J�9>Շ��;��7}c1-��q��m�2�*��P}"�ׯw�<�d�XM+��[V����c\�{\�3�(n���z62I{���M�����D(��Y�LaLm�%��1u;�ТȖ",ɳ�C(w7��u�>���*%e��F)R�VQ!FV��%TFb�DTU�E��E����eA��U
�U�QP^���T�T��((�֢�(1���Jj�����++R���AE�VV
��i�b6
A�q���� �X�
�"�4∦�����()1*Q*
����+!m��\q��H����1&6�5"�Z*���CPR)1�dX6�
E"��%ZB�dեci1��
E*��Z�5��E��l�PX*�S-�,dU�؊����(���,c��f�4�4�"ȣ��1��T�T�
��%a��U!1%`��UA@U.R�
�&[j��)+Bڲ"�XJKY+�Ld��-����B��AB(�H�X(�L
1[f��1����ʂ���H(�WT�r��\eL�Ŋ�P�٤>�	��f��f�̙�v�VNÜ������	V���K���XX�k_`�z��řhr��$����_v0uh�1l��A㪍����ҿ���L�1dϓ��4�^ӏ��R;���8��Q��W��
E������V���e��/���/}T���DY�,vL��U��8�GFk�Wq�z}��_�=� xH����gw�{ie9��4a��R�q] �*�eL�@�W���;�ա�?:c}�w��?x�9I����Աx
�m�GU�n��@nd�:W�a��[P�]w+��8�u5�~3q���<���)l�^:��[���y�G��{7��|_W�������$�����d�F�]�>��G��Ig�v���`�=�@��t��Gŋ���7��#,�,ُp���y�U�sϋ�������K£��+���K��9��`W�.�DZ�!��w.Z����2Ny{a������h���zdo�|7�2����p�x����;rF@�|ʠ���*����)�Od�Dܿȉʅ��m���O�I�tݦ=Qʬ�.9����vo�����OH�n^�x����~GnA��%�#�����0��ͯq�����m0U����Yk ���(W�#���^�?tt�8�!�!���E�p3ҍ�q���;Z+R{�m�����W��s�������j���Zl�}Z,j�����%3�|���	3�tޱy-ud���.9���mқ;e��t|i$�`�ڪ���T���;�C�r��	<r��ӳ���w�U��K����Rx�34nV�]��:T����G�|'O�2�'�������Q��e���ۅ[��^��to!�l���>[s�G@�7�@��P��[���To+��eN�7�x�ȟmh*:;t��M*>خ�]�¯&uL\F�	�����r;��_��׽����G�c]-��)�f�qj��P��Vg������\��<�3��L��t�Ug��g�������q�Ҷ�i�a��3��;R�gЫ���{���&�s�X�� U�S8K˩�b��?f��5I��U5������1�g[��T���X]���z�9���&� M7@TZ���6���&�=bm]I�h�<���}M��5��.�P:#޿_�B����Cr�2��NDQ���@����s¶s�����zϷM>�h�s�C~�����8�;�	�^����2���� 4n���5�]�U����Mn����S��c�s6}�}���_�p�w�G>��iw�+�N�h�O�z�^�}��^��ٙw�Y;f9���s�sQ~
o��Ww�2�=��֏:�[�b�{����Y��>o�ѭ��W��l�2��b�sF󃬧5�p���V�;�����N`CYalvye��V�\�fB�]�dE���@w����5Ψy��B&q��a�_�Ǝ�������>��r ��\�l{}T�/�)~���W�@~��*�0�8Q��z�/;U�3�c�fzĐ+�A^;M�{�+���U�u�ށ,er�%�o�~34ks��^���;���Vv���T���z�4���=�9P�'p���t��K�����S�"�]S��N�_�:*���Y������Y�?z���R���V��J:}>A��*3v��R{�z�s=$��į�#�����i1\�-��uG�_��`���p{�����	@���w�Ǟ��u_��H�#ؿXe=�Mh��g�ʫMƞ����#��o�*}�{ݷ~Tp�����2k���u%]�r���P�}�}���kO^O�i�r7�|XQ�@��^�O��W#~X�*<<�y�b�ˀ�� ���;}=~�1��^�DC�8udU1��Mic	��r��#ٱLK���m�w;�X�z���v�"�ݘ�o��f7l��K�VET{b�b�gY���O#�C
���l{��"�o��j��Y�G���o��:�]��=���}B��l7&b���Cxe2�5V�/��!<�v��I�H����s�Es�љ�5]��VK{)K.r�/��,1:Kсd(���M��qA��m�It����.�*���5;�����O���s	�K�ݱ$���u�qp��A��Nxf�{c���]L%��R������A��<�\�i\W����~mSЪ�={�`[�(�txн�����{�LvgNM����N����#f�F���:H�k����_�_��
ʖ^�d�"�z��Y#'��7���鋯�芩R�Qr�G�,+����$c�z�����lnэ��g7w��\��:<�%xق���"W������>	}}\���C=�\���U�l]>�d>�Z%�+�����T_S7	�>e(=���14��� ��w <�q�=�0PZ.�|�w7Z���}��=�b��*�x��A�쉐���	��մoK��_o�����s𴫫w�H�=�
b��^7���«@
��������L�,ߌ�cn3h�D���XbW�=�ܓ�%�¨����0���ٸ~t��UZ=��Qy^�5�u��p4��D����w�I>���FN�5/I���l_-݆���a��oު��.f�z���𪙱z}ka*�?��������=����ٵ��:+N��荦*�ǆ��@ϻ�ʔ���Bz`���#r2Ǫ #��D�G��0�l9���4��w{w@�<�E���|�~kBsp޾5�n������[�V��8�֖ff:����kB�N��-���j=Oy�n�t�*��,s���Bm叶������S�]z��D�.��r��M�3���V�K��+�~�����_kב[�Y�<��]��o���L��c��H|��/�~j�w���� 9��U�}�po���9>��VET<5[P�=]f�����\Ƿnkï�B��wx��h}~�g�V���W疇�<�R�h�����iS�E��U�p�N�ѧ|&��f�T&���L�����9�OŮ���q���߆r��_�h
W�X+\^%z�6M�ʩ����a`y{���)�^K��惾.�����w�>�p�����,�ay�c�u�,K��s�u�3o�W���"� �����E��&P��w+𫞦������=�h����[���輼�Fr�"S��W]�'�j==@7�U#*&[ U�^.�XJ/գ��Θ�6�&�t�*�~��u}]��]�3�H��dxaY�znT�=�!��X@h��a�Ƴ�s/ލ&�OJ���Y��ǡV�l���H�G�&�=�1�5��#�l�ٸ�4+����i��~�x���9�m[y>�5��	}���_�G�x�޽ <��n���|X_>�V%;*���������g^p�+D���v�'�׼�rP��=E����_Xg�}K���s˲���򳸲�YVY��Cny�*yGw��z\]C�],찅�Z��q�ڰo8q���N䩒����zs�r�;��h�F-�bN�K&�j1ԡRW'%o�W���u���wN|K�IxTz��W~9���}'b'�@;�΀���,��2��p.L]Ƕ:� �ߢn�;���i�_F����V*�u�s�G�W��`z@����OOz��q�G|Q�������,9�b����[.�|:Mk�k��c��,o:������;���������X�lx��"�	Xn}>G�"z�ۓ�a�O������� ��7&{��_f/rQ�=��ު,��S'�ު){!~BO��v�v���uC��6�Oo�Ԉ�WJ}Y���)w{}Tj}� ^�V�9�/�LK>�ʡ����y��Q[3�4�N�~D��F�f�u5{�5Y��E�q~n����]����N�ǫ~�z㑿<W�ʞ<���)x=����"�X�{]�7�	�^�{�UᕓZ}dΩ�d':�8��~��Ǌ��}��7*�S���A���5{����Ӥ�ļ�tUX=����:��ϑ|H\6|φG��������( ^��|�k��z}�j�s�l��Ͻ�T��.q�9U`O�<���a{��c+�=ƪ�%�@����em��$�>	G��8wt��N�dV�}�%�?mG�2�P{Yf�ռm-k&��i!��U�#������rNYX���ʱt��&����kk��5��?��������l�%jt��b���m�V�)��%K�T�_Xt��uӘ@nJ*�C�R.�â�ߺ��{>~���).
��;>��z��̰���M���u.����7�} �����ې����y�p�9H�8���]���~�_�b���2����Eu\�C�ʛ{�طyiO�z|��6��}��u�H�!�o�tU��ȿ���E���^����{�Z�	KE�G�z�碦D����,7�l��bW+��ģ~�/=tF{y/H�
��^�|oZ{��D������║1N{�FJӸ_%�C��W�>�~�u]�)
u���Ηʊv�ˉ�,�T@�T'��M�=���LLSU�o�s�=����������_�9V��/;��O�O��҂�U@����5^G�'*�V釞���^�Wxș��m�9�2�w;9P��:�񿟝�9���*!z$��>�����ڇ�s�M�X`n`�x}��ϣ��3_mG���/Û���(o��U�Z�G�����Z}��j*�\6�w���Z��lޟx���,	�W�6g<@\����*+_��J��C��؄��AF��u��r�+G�cʒ^A�D��&P��^��r�a8j��M7*�o|:��*�玐]Z�_jrT6�vл��Wr��; :ܲ�^����e��#&끨k�%E7;EIu���lY�G3z��YE�]�%�-nD9T���Ɠ����k�ٕ8[�HI�v#���>�ؔ6�v��ɭ.�X�7�o�祁���
��zX8���4wqĵ럣G���;=��w�^���Ͻ�{MǪN�*��ɭ,a;㌁��T�m�[ b����H�e�j���r����h���-�-��=�-�>�\uG��F+�/&u��ɟ��N,��gj�.K�+�5=kN������χ��1=`���X�V��yJN����'{��������O�
�^�(�ϣ�T;����s}+�-���p��u���9E��z��e���{1�J�{�!b��q^`<ځG���l�h�w�������w�}įO�L��exo�Pb}nT�Q7�R�]� d�����"�FTD��X�>Q�¨���Sfz&w���7����7�obK���Y����Տǟ#�>�K�4pu�m��f�G����TF΅_*�g���c����s�x�����?���~����9f�\~1>F��U"bb)�{NA-���}��?j��ٓ���'w��.d�gЧk�����w�̂*�x��A�쉐��	���V�՞}u�� �L�%L�fW��_n��ڹ�2�f�ב���;��j���zЂ5�	f��4p3����f��-ӧl:��}��M����u�ڷ%N���U�9���;�Nv�i�{���;����#��a���/�����m󒭣ˊ�cg���5o6/�#�k��*���� .~���]p��u���{_����T]7}u������I�+J�qzyP�{�?Y�o΀�.fpy��y�zK��3�J��z��ع]eFO�^e��mhXu��eDi~5�2��:���x׽Tǧ=�r&A�ZO��N����}<}��iȟ��ǲz���wO�'Ei�s��������λ�@�%�/���#Cʱe��{F��O�ڱW�t��8�O�GL;�qb�6kN�{e�C�{���J�}���x�C��o.�y]���W���=ƴ\G���9�udUCÓ�c=]eUvmi�����b}�H��H���<�
��<z���+���C�G��A�Igz'գJ��,g�; T�;��vs�R�?}�<�@L��e��~�i��K�]�ˎ�p����'QX�����leMV?luczw=��^��-:�Y)�(ɟ/NBN�V�i^/������U�����
9�7'��~V�uN��x�	gާ@>Ȫ�&"��s�X�ɔ=z���h����q�_E>�jGq��=�'��Z):��#A}.���}L��}�n�1�C���-}�e�l�pjS#��T;7۷�FG��_	�;�-,ABNWk�^f�Β��1�}��R�I^!�
J��^{��IR"��9��Է�TpE�U��8���Y�s���E�491v��"����~�a�����*'��Y�rފ�Q-�*"ԯ9��6XU����{΃�������f��Ǡ�)��RL?_�����٦Cr��b*�!R�K\u���`���0y�.���ԫѻ�[~
�$s�{��7����n������#�{�@�t��V�8�v����>�.�{Y�����B�w	��Y�>��� ;�'�uNH�����{k,�^�Ú�ѹ�L65�"x�9�|���%�K£����>�g�re ��{l�s���6���Z�������mQ��t��=�+L��s�=��X�T*C�m�Z^��R#�w8v�3`��8 ���J��`g��*;g�������<��/�'ä�F��f���}ʬ�(��Q��̯Vob���=��k�C}���"��	XO��ޞ����}�^�q�zx˾��=�K�^Y�.�`�jy؆ǝT����Z]��z�P����+�Ƨ���3�f���T=��1��78M�ֱܠƺ������Ҁ���Kվ#<��F�ݻt=��c�h��L�xf>��j�����:�=�d�y۱��u����IB%6���W����&�m��(�ᑫ�r���ԋ���WG��'��F[��Z=w��]qN^u-�x�N��1ىLRgJ��`Lf�2�zGaOz����B�ss�`s��[���r��i
�>��c���+�f@�g�� �
鹓Q�v��͏i�������2���P��Si#Z���/�4�nP�r=�w�������z٤�qpp3��ͨ�E-wQ���->p���uA�k��	��^�Ӭ��S�s<E�����Zͪ�=��T� *�v	۳	��U�7ɧ��N�n�/� ���3����N�l�=+�/5�U��R�:D 3�*�ư����|��`<���oX�X̮)��8��ۜ�g0�Ms�r�|��,r��ǧM��� �X��*DϹ^`T(&�:��W��vE�5�T�"j	���]z�d��]�О-����lYJ�M��- �N�`�b��+R��YO�qW{��f��'k��u u����k�z��e�4p�[8L#�Iuę�+�9�b���׆ޭ�ȇS��Z���8f[ǃ]գ���h�|;��	S����h5���V�ru�3����#���#��&*e-�O����H�<R��d���}�Ţ��<i�&�۰�$ɽ\���^Wa��w��pN�w��M4ۂ�3�1���EQ#��wD�:�M4]��#e<	}О���F��,N:�9܀��b�6z�䑝i7��[�M�D�%چp����@��ԹX]v�ޘ;���7�cCב�=�鎧��..V�N�N�AM�ƪ���x���9ڠxؼ�}9�֋n���L�9Z��9�^`r�e��F�r*�A��S�ۈ�@u�]us}��֛s��׆�'f^��Ы��҂�j8��RXl��WJ��Zm���Q�ގ�x�3M�ݹ��YO>h���x��y���j����t8Hڗ+����4Gu&X��˽���"�,xjZWW�Cu�a	�;t��C�.�:�L�1ޥ�om�*�
I�t�?�,�AA�2�އ�+G� �����,!�����ېL�6c��t����pn��:4��8)C:��H��e�� Z���7�`Z�P�_%�f�pv�-��栴Ue�n�Q�$֔		�Ө>w����w�v�Q��eoG/�����-�ľ�rk�Zn���Ɯ��W%�ji������]/qRr��`Tzn<�8�\Ƕ�O�p�ﰡ�l���50;a�=X3���������@��s*Z��z�C�l*���v�����޶�Ŗ��lU}C3U5�|]��ؘ��z÷�!�d۹��Ƴkk�v�v����*$}o!���V�7��ъX!,zm�κ�윴}cG� C�T���b"Ԫ��AdP���PU�J�K�r�j#�D�c2�MaVI����a��k�Y����"�)j�ȭ�+%aX��VœP� ֓�,H�X�T�(\ִE�1@PXb�VE��,�Y"�
�+B�,UEbe*IPQA@Y5B��,AE�

@U��E&�q1f1`�E&j�0X�E�N�,�Q�Y*(V[W2�Ċ�AE$Xł�+1&9h#n�@�
ŀ��B)m�+Bb(���c cq
�4���T&���R()�%)jJ�
Ƞ
��(��P�*�kQR�FT(Ȱ#�V
�+$Y�J�c&!V ���" �IZ�X)EY"ʐ�����Zb!�T�)�ńX�(�T5�;�wp�sz#�6֑+�e��wA$�-����yu�V����{,Xu\���$�[�:�K���]�(j�G}%8���!f����W����p7�����oS��U���3p����۔}�X���>�g��/n�׈�}���^Q�Z]�L�.#\��͆���3��W�N�x2)LL*S>��ȥ�j/��*�^��ܶϏ��-����eU�1=���γq�>E�t�T6|σ���zq\?d�z��ױ���m�o��q�T|a\G��������2���ҙ��a{y�|y�(D�S���f�'Ͻ�����ތ�Q>G���ne ���w�#�*��MF@��n��^�>�q�F��{��)�ϡg�ⓔ���#}`h�z�~�,��ω@{��VxE�×�bd�����Ͷ�����w�ix�y���'E}~�r.��E���7o���*'u!�1�4|`�;$�>�q���~5}��W�3I�����kdq�uX�/�{�-���H�Kf�n�4�t�:c)/Z�ʯL5>Խ�0���5зv�לw�����,�Rl��rCɯQ�	h�M�=��1�MVѽs�ݐ%�2����.�q�Z��ܣ�t��Xr�N��:�mͧ�U�V�۩�4'>��I���u�pu�.�T�~�;m�j��}���t=�T��|�b������f���΃���,޾KG�%�1*(*��>SRw��ݨK�����nᆻxf����=l�������}�</9J;�W�(y�W㑮��9�8��\P���@��5^G��<ܭ�==&�9M7�\3���{��T���=��1qUO���<���9���J;s��]�g���r�T_�>U��{��7��3_mG�k��/�"9�o����޻��9f���s��o��'��0�,P��XPm��J,_�օq;[7|=�$8���g|@��z��v��O�>�TL��ͺ�;�NQ�=�O���%���OO�~���M>vz�E>�N�{w�4��pŁ�9[�������O�ƴ���}�{ _��=e���wǣ\����{r�u9ɶcI��/��$U{ 	��/�8G�����F-�l�D�wIYQ�5���ɝf��QЖ��Uw\�h�U=}��{�R����}�}�\{+î]��r=��羗8�����5�o��t����/�{�~2ٿ�g�L�sʆx�����t��Xྔ����^{�6V�? =�x��򫃝�C���2(Sw������٠Ѹ�uC�Β9�x�;���k���E���1�	��Ղٚ$�j�3�W]���S��x�9."��:�W�zN��B�*>ݡ�y0�J�׮��/�;�{����k�}s��f����Kk�$�\n
VQ�X�a/��Q��0&�ζ�mu�l��G���:�j�xP��/X��o7��K���=*���j4�t��Η�4O�i�;�ܺ�}U#*"]0,��}��{�|��a��G_#������8�f�&�w��䯮; t�,_�1-0X{uRL�� �^9��(��Ϡǡ]ߕ.�=���yޔ<�W��>�H���dQn��Y��n�R&)����݅�6��V�U�ի����a}-U�h��y���t�ʸk�]���~�;�f/�]E�L{'.ފ�����i�x�=�&���x\{ʯ����ր��X�=t�����#�ѷ��=��bu��HA{�莫u�t{O��qzj9X�w��p�z@�*!̱�~��/؜V��;ʱpv�F5�˪�^�7^�u����Co6�z�'|f�6X�3Q��r��{ꏦ/|���6{�@g{a��w���=��ʛ7�H�zr'������gFN������*�Ǆ����X�> ��s�ݛ���g�Ѫ�ʟ{f�{�ٍ�����8���C���/6kM�7�^T��s;a�v{�s�=��������Z:��~/}��_�z+����uLó����=:����kr�݆MT4�^c�M,�Dn���b���B����fD�xf�ۢ�bi����%�t�*�23��7p�����U*�I*�5M��n��M;���{��Tf�V8�tM5	B�U�ԇ(�^�>���t�C7��4�g��a��/K�CB�m �pK}(aS)�\�n�̒e�j����3���Q�,m���N{�����\w�u��<��)k��6�GG����>�V=	k�9�+|v�p.f��uFL�1q�>^���4��|�i��}�Wt��k�}�;y�W�����*��V��*@}qU�LT�"���,^L��S��h�1�w�r�<'�B��A{W�=cU��4R=�ޫ�ǡ\�1��]�@>�"�&[ W֥x�ͦw���z7ޮȳ�z�S����z�9�%��:wM{���
�M��2�����gҽK{)�dtǱz���s�R^I��Q�Qu�X�u�H�ԁy����~�R6��p�L�9 �Lhn����Z���K����xs�_��	�x��κ���\
���p���`��uNH�թV�MD���cc+Z4F��`@�~�DLW���x�闦�xT{�3���x�J��=��P�a[�ݕ��U���۵�#�$y5>��#�r���w�x2����m׍�V�κ���o�~��E(e����C�=[��v&���{R��oj�&Sj$f̏�W��ft�+�Ƹ�n��)b�}�>h_K��P����/qk��ݫ<g ]=]D_Q��Y�C�h���N���56dnG�e����:U�=#��G
�MG�̊=�zL���G	#� G������x3�Bd�(��?�����F�
����G>��#�9P����.����5�t���<���Ӌ`1S��}y���/}���G�\[r5��>c&A� %a����{'�=�[��׸���������lf���=@ϡV�9Ҧ6#�Q�o����U	�e�x�Ϩ#�;P��ݳ��-����^n��oE��kS8pk;>�`	����^����Q��eh����<�����J�=Y�ޥU�����J�2�����,��@��@m�[�տ{��Ǟ+����Y���`�=�V��>C;$������T�a�/rg}1q�Bs��f���7����)Aeڻŧ��<�zl�<��<�9QF�K%�^N��~��/&u����/:d/��%�*/s�>�i^�6=�M��ey�V�7#��>0��2�f�R�	��D
��)���K1���#���&�ݪ��5���E�~����{�c�z�ت7�~��G�z��� �D�d��w���΃=���=�axG��}Y����;��$s\O���}@h�z�~�(��~�8o��h���-ɻ�N2�HM��'�4�Ys��}e%hYis��,��λ+:��� �QD��{�i�4�T&�|'zo3���w[Yj�ݜ��bL�ݱ�zr��L\Ԡ3d��wb@���i���ƺ�[r��[����Γ�5kGP��\����}FFT�~�Z>ݘh�����^����L���8&�=�)u(���_�s_���Q��ވ� w��/�n�D�s�>�XZs#e���T;u�����%Ʒ�5�ڧ���F�u��+ڲȯ�*�.��7�۪D���t� 1j���ا[����n�﷚^��F��~����;�.�Vh�q�[<ja��c�M*~���/�w4�^��+P��Fo���R��c<�Y,\?z�����Ju:��.�^��W�܉ʇ���a���t'ޛ���1����R!{d�Ǵ�����*�P�T���ޠ<��ݎ����rx��W��c�4�k.&�F��:�*��#�{Qכ^�|_5P�j̿�uG�^��<n=��g*l��	!ט'2��;=�{֦fǍ�h��g�^:��2v�o�,{�a������fs��:,ݯmW��ߦ�~C;�^׷:n;ޣ%q�V�d�c�+o�k�xg��3�i�ּ��\jT%o��F�����㞪R��U�ߖ+�����<�z#�'���2�kK3�:��dM}�\:���]��JS{_�;���{�rǴKͅ<���7�6m�u#�����ӥ�wT�h�$�vv@�j�ӳ����Dd{6g'$*_^ιgX�� s��53�v��eN��F��&R�J��"#�X���j�����_@:�a��J��ef�p�Ix�^}| ��(������������(����>9����a�WLVRB��_L�I6{:�.�3	�|�x/gT�:㟯�s��:�=����uv��{��ES7.p7:���՚���]��*��(�0=��\a����Q��s�9��=�/��8\<T���dOgLGJY���^SεY��+�Up��6�?\
��'/"6h4g��D)�r<{�k�q�g^����at	�����9j�+�+�*�.��f�*�}�R2�]0*.X�>͖_V�m��0���B=�K�-����F7͟}�#ME�w��E�ىl�(=��
�W�Ð\�͟|��j�RV�{�]~���~>����=#J�ypE}~�nG�O�y�T�����*��2�d�I�b˵Wi]>�]�y�q�u�l�9��+#޾�g� ��^7�TSG�&@zs@���s�>=['����P�:�T}��{���ڼ+�y��������R *�{,
�y���"G��ez�1.9�.�F��ѷ�DuE��5����/M}��C�~�f���G%�h�^��H�=���bi�HO uN
7�vb���\ �#���kk��t�_u3Ot�����{��v5e�}ܠ�ö�_m���M;���Yy|�����Z2�ծ���2�����+���V�9�җrX�cg�O�/k��0� ��NKy���d��l��gC߹fd>n�}0���S�n�H���k!l=g�C�W	JM����O����=_��d�a�8v5��f�i���R�����^�{��h�z���S*oݵb�=�/��	�7>���N�<���/6kNL��E�y����"�r��&���*=���p�׀���["'��4d{���>z'���F��Fq��^^��*�j�u^e�E��g��Y��H�G���������]��pW�y��<�R�$�?u����M����ש�����E�wq�ɝs��+�X������~�K�}�]F3Pߵ��Y�74,7�ko�}z�]�G�?jVE� ��x
�T52���ϗ�9�u�9��Z<���̯HGwѧWz}*�����>+"=�3p���� ��DY�,vL���^��Sх\ʫ~�Iz��}�Wq�w��nW�<B��a�tk�J��"�l�H����܋�U��Nt��
�����R\/y�މH�o��z���9�j��6ɒ8d}�Ɛ'z������G��a��o���v���b��b5j�����a�7�10o�V�o��Z:,�%q͞��ƺƁ^����|w�<cD��bge;��|�����X礠�������n��.v9,"�i<f�H6F/��]�G��W�S��e�+�2����5Q]ŋ�ש#��R�dhQ�^����;�2<��d�S���֯S�./>+g��J}gIc2����T;u���/z� �=�E�z|����oU�{"���������<X��*�&����_���ߵ/�g�U^7����k���B���u����?G���e�"�HG�n���=Dz��#~�;��_r�p��a������N����D�d��G�7����;���y^G�,��*��v}�_���<���Y�{6��t��k����&����g�rJ����܂+�	XO��o˪=�;����\'��Z���+az��=��f�i �W��>"��������^�H_�BO��v6��Y����=����ϣ˪l������`	�V�Kվ#>�b��nT���B�8�1{�|��IwC�zO1�a�|�K/�k���t=�X�ߴ�Q����U��}�o���n؏3]����{V��Ez5m�7�{�Dw�mh+*���&��'}1��'7�G��k��xy�ة����H¯
˛C�Hh	V1�΃,�΃Nq����L:޵d;}�ce^*ڏ�	��^��&���6�Z{�>fx��A��D��"Z,j<(`��ڷ,������*V�̇��!g!�%�����<�u�=ӧ*�m��|������x�;c�Z���%�^N��n{Ō'Y�ɟ"�*F�Э����ʻ�'����6|�8�W�ګW��g�G�*���8˜��b��h���\��ݑ�;�p�����<���b�?^���O������-3�+�����e��{����W��(m���)Á���_[���6��_n{�@N�9r�;��@`~�S�NQG�G��C�imf�;|}�.t�5>ٝt�"�%;@�KGۛPѫ�n}I�HE3����鎣�����f�>��]��ۆ��R��ޮ��L��Dg6�D�>��XZs6_�_uC��g���Ol����f��:���>%��a^��tD���D��Q�����L����Zw 2�ֽ��� �7;����[a��Nc�^���z� +�=�5&�D�	h�D�C��2�LLSU�J��:�نks`n_����]��\6�Փ��gǾn�bzr<�����|i�sU�+'*�\Nx��fUftz��m�n�Mp�<0�u�5��u}^+�V)�j�|_���P]P�s�/D�wb �=&`j�߼2=���p�Nh
�͵�2.�0PZ��/pۃ�?��8�v�^�4fV���ZT�v�MC�s��KeF� �ր������/�۹�0�jLwYFf�X���c�j�\�x]+�4�s/�wRh���ٔ�.}��uH��2hGs0uހ�&��]�]è^�KB������H�ÄR�HR�V��/�LԝmG�m٣��F2��t>�9.�m�i)��Ŀj� c�V��r�{���;�@_	��_��q� ݖ�)����q�V�T��v�9'�4h�t�p�����F^�o�K��^.�ww%s�=m�\�pi=Q�g|���|�F�/Wp{sl��ދ`Qv��׳Eg<Vþ"�p�(G��������|(Sh��9E)�Y���X+h>˸�*r=��卝juf�s-��Bg}�C�1�g��^*�.2��Y]�L�k�	�y�z#0M�̶]�,Mp��j�쩮9�m�WKSO ��N������ս��9��nV}��޹f�cK��� 5�TYݗl>���V#B��y��/]��66%�Vd&�9�Kj���f�ݧ)�����+u�YP��/Jŷ�\�u�60�w����j7�@�Ƶ�v7��4�t���������>:�+��U��lS�.$��p3}[�g{�%�
C8�g]o��I����E�a��8f�$:�I.�����2�]�ׅ�)v�2��u�j�Y��ʇ��qX�P�o\���d�]Qu��3�4��";�8���پGAQ#�h:{06��h��t�Mv9�^gS�g@��5X�jA�+':�
��>E)1N�Ϻ�1vI�S�Z�a;�ɂʛ���������Uϭ����i�x��y�
o�:��(YD�Ю��c��.9�9e˫��u��9��
X�n"�t���]%d�-S����AƲ��ٲWh�M�}�&É��5��c��i�YZ[��")
�S�W�	S{{��;F7I�@bA�x6�Q����"�!��dT"��b�-�Z*��2��{(�#/Ӯ�FQx�ې�Nd��&y՛,�QO�f����s�%
d��$C�-գ9�9��%N�)[w��vvv]�p�n��3q�m�T7����'bn�`��J���o�Zh-��9�v��㰴�X�YFiN;t�Yٝ�7�u-=&R@Z�{!E�\
󹜉f��[���X��n�P�P]���'Ҕ��_,�)��Ң ��]Ǩ�I�GC.����U�3�6��(d��=���u,�ȸ��́�jXr�_a{u���2���r���59Vfe
���}������h��{o�r�d�W5����=�'������v�R�ή�����=�s��1.mW<�oW(�%d2wf��d;�ŢH�B�B���q�,J����ʌ��8�H�*+SaN4т������2�0*f*ъA��F�ʦh���ɗ#}B��.��`���9z������+�'�s�q<
mv����v>o}����ɦc�"�YES(J��X�AT����,�5"bV)
��L��A`�,F"��T��PQE]
�!���R,�QjVD�J����DJ�E���
(E��"2)&2T��ֲT��YAaZ��X��p-�F,Qf$��U��*Qb������)U!�%@Y1�Q���,QH���h���1Eb���Et���X�(i$��"h���b��j�HT����1�1BQ�""�Q�Ŋ(* �
AĩQ`(�
�Q\��X,J�f$�Y0ej
�E ��U`,X��ȢŘ��LdP���#1��6,dPU%d3)Kq
����8["�̲j��I�.��i�� 5��7�d�W{��ʱ������e�R��=[c �4�T�]�$y}Y��p�0Ќ@�t*Ǆ�^�มj$�Y#��?h����q��
�6���&kj�[{��7U>"�P�n=�]�ǭ�ּ�wTu��`#�z1S㖕��b��\��ǜV�J���R�i�
+�G����tV��OV8�3Ǯ&�7���ۊ���p� ��>��o�;Le�֕y>��\�������,swfjl����>K=�n��9@��s7�sU��r�;p�T�)dU1��ZX�ɝ��vV�1.�u��r����*��q�� ��*�o�����e�����F-�l�D�wIYQ�#*υ8��F��v��K�=�F�g�>��~�a��ב�_�O�lp�!(+��bԫuy��ksq���u���*�~W~�6��6q���%3y2���yP�9��J�K~�_�6������s����rb�,5��l�+�]0NQ�)���>N^F���	y\U�Β7�G�����&=q����J��ϣv��@���p h���9�/%��G�e�Qա��]T7���df��Fz���W���q�^9��F�������^�Ƙ-�`���*��^++��ӣu��3��5�B������x�J�Q��sV�՛4����薲��L�߯U,�Y;c�y�rm�ܐ;�l^��3��Yғ僪�șض����Z�<��-�j�A^�����]6���ໞov:�U���j���r��شO-X�w�ͯ_ʕ�X��\߈	z3ِ`T[b�\G�O�8<ߪ�1|�L��"�6�fT�P����b�#�'�;�|<�q�s�L���ׁ^�hg� ��^7�Pj{��i��@˘�/=�>�h�E'[GG���0���{��^ʠ��t ��v��
�����l2�ٻ���cݐgq�Dz�;'��*#��Q��C���6o��@y��;̡f�ε{wR�+�o����)�t*|��r|6�kC�ͯ	��4��c��3!���k�N��{/z�ߨ�ǣS�<o���{E�Y���,�'���z�����댝����fα�6��u�@�g��w����g=P:7���q�ڱV��t��ށ=���HGn'j\e{�	�W8]�sd����]N���&�����@L,���/u�)��ۯ
}��_���9�uNO�������^�Z���^�g�YQ׊���7��T���s�59��N�Ї��E!W^�G�/fS��Y��~6_���ѥ�Q���w�g}7��7�,m��~ӟG�_��e�q�[6{����m]z��*��YΔ�oK�R��ǽ�5��N���u�׮ƒU֋���(��r��p���+[�Ǝ�pJJr%�G�K��z�}�!�r��o8�Wb�NR�9z;L�1bB
*������/�4�P�jY�)��tDX��8�teic��w��J��r�>��]�|VG���X+*�	��\<%9�ɟ/O3!����M�a����S�n��.�{b|,�>��R7��Q���,��uL�:t슬�"2�ȱq�(z�o�oeܫ��E�ϗg��G���{O�ޟqs^��@YR�vDk�vn=.�}�R2�e���i�2m�fH�.:Q^�9^�^��=|<3�y�}�{ސ1_��a�j=xbZ 8<26<�	+�6'y�Qo��si�Ȃ_�͘j�t��z�9�u ^}��4U��ȷ���:�q�/.�����gy�>
����f��4+� ���@�~5�I\7*�EyO�=X {q~./��߻;ÚvX�=���.=!
0|:��'�s�w �r	xj!/
�\{���
O6�O�nx]�,"{�z5q��RT܀�{`S˯Q�*�=�7Lm���#�V��|6k,o���q�f���]�v��Gz1z�Ɍ��P��t?NX'�]�n}�gӕn3oC���f/s��ڜƒ[3�^��zlg�9Ւ��:���@��/M�3� ��V��O�잨��3�}vO���.��;�$�7a��K��S�ݷ�xk)&[Ys7��mH��8Kf.�z���~�o�O$b��:(eξ�/���r�v[K7�-Z�o9b��)��8�\�+p��'L��3�:0'l���]�q&���k�rU�K:V�u���V�n�&�i�:���_�}Ψ����[%g�T$TCBP�/�:���vt�12j=�#��^�K�����
�6�M���M�0�Z�`%���ʘ�n=۷B��x��M��;g�0'�o��(����d^K��y+����>?)���� lRu�.�������}�T�6ҳ�']��y{o�ǒx��dU1�5��d��b��!9�G��U{q�����x1I������L�E_�}ޤ����q�;��-�����[%��*f���b�ɝg��es��bn��ϗ���Cz�����>gs�e{��*���zǌ+�%l�I�\��Ԝ�YʿUe����7"������ςy�S��������:���:��Ze�o{�=r�/�8}��1O�h������5~��
���[0�Q�w:H�kb�ߺ�h����>�l2��
W���:����L��ۙ`{�(�ʉn�7�����4j��~�����#��	\����@�N^����Y�X�Gm�ȸ�T��L�ٿ���TȘ.}��Ni~*���`�	�W ������=ck���l<N�zp�uduj�e�n�7�{��|����X	Z� �7k�y��P�a�&6+s5������wes�j�'�jby��UΡy1o_]3x,tq?zh�q����TYC��q�rНs�b�m�v�����Q����|T�g#��8�>۬����|͘(=���3�tg�Ҵ��S���9[c��yޟG��G���鋂����8�{rTC�����͛�{y^&+�y���F�bc#�4/��}Sû O�Wܪ�a�Mx�����=q� T/g��95^G�yb��E�T;�g]v��J(���t��^:�:=�ճ�}�p��Ϗ����g�B��2��Ye�+�!"c�Z�tjr<h����lvFn�{6}����f�j�wu��d���o���/�\c�(R�~�ٷ�����s4}蒎\K����c/Ӂ�L��,{�o�,	����u�WT����S�Ԧe� {�?Q�z��o�۝7�/H'��D�%��c.2kJ��8v#\����#�ތ�Z}j�π�|�d
�W����\����������]�=Rp�Ȫc0Ζ6��wW�<T��8�^�>�l���ꐷ:� �]^��S�S���������%G�{Ò��wY���WB.)�u(z2gY���a{#�C|�~ӑ�u�{~�W�9�C��xv�ʯ�g/����~��טd�8%��}��w�y�%�;X]3mĎY��gE��믘���=x4�w��qV�YqL��R�v2������~$��8�
3���o�Y9#F�[��r�t�agf����/��eZ��yY�>�}{��;���J㫾лd��/�������{�W�0�f�e��=���w�9�_dn{A�r;�̢�o��7�s��H��
{5���]\s"��n�U��/6h4n#��9�G��ӛ�U}�n=��qQcK��nW�_��
ʖ^i�>.@{2E�,rǑ�F�	�c�
o,]���{��??r�x��V+L�x�3�g���'��&%�fn�B��Ⰶ����w�z��پ�g=�_�����;u]�G�ԋ��H�=�TE�f�g�O�����ɾ��������~dǣ׵�8K���>�=����[9V߁{��pʠ��zɸ[����?*��ބ�D�-M\�s���1��&&�մoO�{�ó��+���U~9�@y8 S�5��Q5۞�zښQ�~ ��������[�p1��C��l������l�7
�ï��͑�˯1Jfco�՗{�B��o}���=���*�K����G"r|6�ͭ�'|f�e�2j4��F�f��jwP/��G��9��w���/��<n=�������Ĳ��?�x�������
�޼��y����W<s�1���EA��ʹ~��u�{R��/D4��\U�W���f�4�'�o��Ы��s�	��㗣.�����>¤�p�Y��3bط+��c����,� �G�*%r'�����I�{�'c�#A^�(\���q�d�����a7�f��	�CqQ]�F�P3�]�[k�����"���V*���Θ�xZH�8ra����L�)���7Ƹz6r�ͦD�����Zo\�����+*�/mx��h�uׅ�}��_���;���^�ʩo�o��0��UB�Q���������T���vE��|UtG���'hp�ql�^P}CykU��C�z5m�u�J��,eb���梨0�f�e���~�i��K�]4��8f=uw��y����=�գ�[E���\�`���b���&S���^*9�7�m-ZY����=���g�R�h�{=C��1��Yeg���mӠdEVG�|��v�YT܂.�Z(�]��A{���c����}�>�p��q�¨�z❟ =誑���G��5;�j+����\+��g���C������L8��JG�}@m}�_�<0���<�L���q���Wy}��x�\
ɒ4z[�a��QP�B�H��K�6r#ޔ��X*/֮F�0��Ѫ�C��9GwTe�ϣ������̣#��%���D.�C��x����k�4���<���+��E���
ܛI��_�ժ�)����ˮe�z�����x�Ǘ����>��`Z�PA�BVa���+������K{+ک3a[s-�׸_U�5�oP�`��]k�k��۷�X�SE�C�7w��w&eY�܂��=�eɅ�c6$}@�K,��tBr|XP`�e5DM9�;��� ;;W�ǭ.5��?]�~��T��}U>�>s:�I���t<��p�h�}7LnzH�E��"�5���bM��vMte���S�u-�w���߫��/��C�K9����>%Y蛟#��n#+t���cT<�݋��>��Dy���9�f�k��r�'�㛳쌍��}�#'�j�#����|��>~Ϋ�;W �N(��P�=���i�q�^�qޞj6�R�_�G:��.7���z�H�^�Hu���.~mh
�'3�ŷ��e��}�j izT<ٜ;�i~=6z�m:~^����%b**|�K�����S�Ԍ�!�=��<��o�TF"t�{�V�,��=������]������v���od�{6�\����H�}Q�|��+�o���{Dw��ւ�"����kK���L_��'7./D��y�~���m4�|t֎��}Ο��q�^���+��̔JD�y�Up=��Xd`�.h,wB�u��	����S:���
4���yי�\���ի�����w�&Qr�r7NV}��(��=2>�lc�֤F�.<�ľ.�U�������ZΓ���{���]Y��1X�0�I�~8��tP�T�<�Њ07��
�5�����K�T�0�M��*�J�`��hg���#<�Ky�����o%9roT̨!twU�۹���/HǙ�d��Oy��wz'���W�\�A���>��1��\�+a��oې�7�'����t<���?E?P��t�j5~ڇ�#��j�}`h�V����^�wc��}K�+�Tz����9deD�h����>چ�D_uC/ԑ��kt�eH��u/9>Z/�N�T��3�.��ٳ���L��.}��Xo�e��_���π���.�	�*���*�B�o���Q�zF�y�*U: \G�O������=㣭#s������Jw�6}�r��sxǷ�^���O�9�z� W�nAy�D��7P��UR�2=�É�[��dǣה��}��q�|2�U�ŷ���S��@������
��]l��U�w���c}�w�b�mcB���f�<��3[���o}e�w>9����5A���0�ond�܏r�>����Ȓ����Av���n�;�������~5�y��ꏈ.�H=rY�wGbا�����Z=��M��q%>��'e��NQs�ӡ�잎,��^L�L��Qܶ�̚��b�X���*�@��zls��.��wS�Μ!����"�7͸�*T�A��kTr��dC,��&Y��Y�g&Fm������`�`�깋gP�pA�|v��CV�f�n�6 �ef�1�r�e�0�V���l����ȳ:�29)������T�|s�����W���J����JvX�ʭ
�'´�����r������eH��-S�G@��<�}j�zx����Q]��nx�Ǟ��9꓇VES^���@���T�Wg��Ӌ��ޙ�o} k����`
�J��޹��>�b��F.�ϳ�3�~~�y?q�5�����۵�o��Y���)��+��Ľ~Ө��{+Ô�!�+��r)m������[�4=��9ЯMϧs�D�X]뇀��nX^<�a�.��7ҼR�t6�~ʺ���=�W�p�oh�C�CG�b������P�`>��6�7p*.|��٠Ѻ�ußc�}7�����5O8��Gt�xyջ���R���2f����R0�`e�G���n</f&����;��=�}%H;�^��c#�
�9��F�����X}^���ĶnfHOå��������H[�g����̍�W���Cwkō�yS>������1^�n�DG`�Y�7���c�oнBng�����%#��a�}ӺX*�۬������u��������@!I?� �!$��BK �!$���$������!I?h!	'��B��!	'��B�~�BO��$�BI� �!$� �$�����B�~�BO�BI��B�w �!&�1AY&SY��{ d�߀RY��=�ݐ?���`�� ުBI$E*JJ�D�U ��͕R�TR��T@D�K��P�)*�*�H�QUJ��Y5UX;T�I[i$���M����A�3��6hZ� � ��f�Vl�Xj`� s����f�֐-�V�%KV�5��p�ۖcB�A7sAl���#]� �f�m*�S : ݲR�n�ӻ �a���n�:+ur�!��8ݵ,��m���-ai����d�*p6�fX�[1���
�V[&�Q*@8.�SV�6ki��mf�ճ�\wfm�if4i��e���Y#(M2�v]�J6iZ��m��f��ۀ     ���T����4  h2b)�IJT���4���&M#&�0# #	��14��~%J��S�	�`�M4���0# #	��14�JzH)h�	��A��=F&�m2�jO����A�Ͽ9���g?�.��~�
���J!� UP��J�UX(��(
��

 ���#�J�����>�����u�ԯ�`���<�BR��� �?� @��@�E
Ua����!�~z������R�����&��EP%Q�ĺ������?c�/��檹eB����=�~�N#��K��8��؜�8�5������=�P9�E,�-��1^�Y�k��w.��j�$��ɭЀo@��N�F��sj�^�/(^�Q��i���@n �e;�4u��(�W���)��Dӆ�hi�^�W�F�i��!��y׸����V���HU��އ($Rŋ�K�OB;S*l�
��{n4�]�w�i�)]\n��q��M5o
qn�nͰ`�ۏdݥ W3,�i�����ҋ�nH�$Fa�����쏉���6ba�*�m�
��<ͱ��%VQm���<��h�.XZcbEve1X�7�2`_��nv�Ɗ)ꡋvڭJ��̀���112�ٌ�U�`�NY�W6�p��9ǕKo��n�b�M])�Tq2��(�r�̱�]H��b�Wkk��f��F����6^$�m]��)�^�5$�(ޕ�Y��J[me#�]f��^��^� ���q,,
���me�Vo,���[4�Y�ad ���dZ����1L���v�0�͋ 7zݑ\C6���K�P:�b&���T.E���"�V8M��R^�c������vp�ֿ��T��Y�a�j�u�ުr���H�p0:�Ԣ�ۚ�*�e[��#VI����O��	W�yY��Z���xN%GJR��,�1,�̚Qf������&�ֵ��@#�;A����nR�t��J.޸���j�l
�]���ލ � ��d�B�6�-7[gPȳ
�R��9p��5�oaq�Z18.Y�ɔ��y�6��ޫ���3j�Ӣ���q��2�=fև4%LQ`�N��#�����rQV�H9t��܋Q�u[̸(�,9m�m�1��[�b#�������6��+
WX�^iB;ޣ(6V�SZ����^|i�q^ж�[,3�@A�OU�wz��[�(( ̺ug�W}gJhmE���je�8+j��ծݥ�V�r��`A^a�#/e�F�KX�CR�V5�*����4v;B��An⚝��`�hC��ЍԳn�>-9-�V���#��,ZZT����ԇ�E�j˚
p�6�ڣ17r�ؼ��ɉ	D���+ks%S�Z(���`%��8�B��vvĲ�wD���i�6%���!����.��$;̦�w��c0|�U	�bTr�
������{��V����Īơ���O]�t�J�oQسcݙVj�U�wdS,һ/N�Q`�h�W�f!��C6m2sU� ���[L��:\��xh�֣d�SL��M6-����twn����j^�q�jV�٬n���H��Iz�mQ��q�~Y���V�`m"F+IM��~��IGnn]
g��H�ӛ4�������:3ڋC�v������m�W�h��0*��m�Ʋ�ì��Z�7����J`�N��B%`��˳!��0�.��n�ŇwB�ZX��ʦ� �����a�RM��lA�/F�&�Zv5��E�3k�W��om�Stتkm5�h��@ս]fh\L�y*��L��2e(��[��9Q�K��8c�m"崬^���ײ��F��F���Q�M�2����7+�Kt^яsIV.�%[�x2�n��cET��s����H�w��f�YB&�A�-`,��3�@��t�JX�1��@�n���R�ӳA�X���Xմ�WybQ�0	u�mbTV��.4�v#HU��
uEy��p["n������&U��]4MH��35�I�\K^�fb�����fIKE�(�J���y��XD��X����U+V�)�1�D�'b��4��5=���u��޹/7��c�a��_��BUr�Ɓ�iy�(�&$<�������?a��Y��w|���ogo����o[�]|)X�$P������ty�ucN� k�syp�npk��w�~����p���B=���1$��y���"����@�5}��H��=��m������99�_h�(�"��+18��(nR��]*p�	 �3�2��, ����	�%�\��K.�޺�|9�흔��fv�(������v[�c�74�œ N���Bͪ�;+h�u^s�	�Jq!?��N��
���������G�÷Fօ���J��l�����x`g,�(� �N�#�Ԣ���];-��Qՠ�z;4�Nv�,���Mu9���=7�Ł�Ӏ6�ش�G��y��
�"cu�$�e���_moԹ�L�HU�⹔��7��qmJ)V������
�>w �˓�ϋt�������.1����R�ڍ�P�%vm��SO]m-���v�)�n��tT�зI�L�B���;d��)�E7�v��u���}bLTVn�t������v�X��t%����)�l^-]����=D�E�S�өg���2ӷ��O�f�g�f,Kn:O��k�^1}�p�q�%f�+�iˋ�� �JM�E�L�]H�șZkx����hv�����R"�M�Xk���:<N+=;�Wx��Q#`�O�C�tU�8t���*в��.y2��vb`����\f@k#��9��ȃc*S�wV�bu�nn�Y�蔕첊9�7���<�W�t��f� ��U�V�J|��_E�WX�ot��;BY-p���B1�:n-Ϧ�r�#B�8V�Hsa�J���5e]+1���*�� GNsJQ�F�#{��nn�ܾea��q\�Vq�O����s_��-���It���.#�����ż��d0г���{W�
�l�r�����[��x�U\*b�W�C`V�K}��O.���6�P%�sU��7&������{ֶ�%�����k.�DU܍$w,J���GOM(tm��)���
�ޫ�H�����|�Z�
�T }{���"WYO&���G�X�����#Ⱥ�
���©L�P̽O�ae<�`�0�S&�w���I����-(/��\�V������p�k+q޵|xFټOT]WY% w�w56����g�\��b]V����Bph��u�d�:*�L��fe�h#�&��݇D�/Z��=���hN��d�:H�l�T���;���ͬ��x��e��g�^���]&y�+:�N`�G�ӷ��X5[50�/P�7��˄M�,��X4�4{6�|	;fT�I�]Ev=׎<&���Fu㤝�ZJ솕u�`�J7]{�+�(!Rn��&q9c9�B��_<d�R�J��΄385m�eK����n�3�YN[��u6%�U�)��Q�k�h��7D�c���:bs��ؕӖ�-A;�8���r�*�Vp�
42�
��	5q)1�8wk&��Y1�����e�#W0wiGx�m�@��S��،:�5����Wb�Y�}�m5>M-����tR�*��wHڭO��vV�㧤���$ ���`�t��P��8e��_X)�__kj�y�+tDC�lɒE��5y���u� >R��:�����CG;3ࠔҢsֵU����x�
�R�Ln�/|�7Ʒ1M��[�c��{�vk�����Ӈ��U��j��U���Y��l9�gt�cv�/�\C�o�u_î��\��}��[ѐ�w};D�Z�����m�p�nDa�qp���6:Q4"������֊4K�7��9�$S����b��rkrl[.Y������:��E��s��,�RM�[�Q��
۬x����+"WVWs�̫N�,w�2;�T�>qb2΀^�Ί�_������ߪ�	�}>��g�@
� 1��fh(����P�l��Q܅QT ~���tӺ�?����?O��XA�7�ox���	�����O۳�5��
�h�������v�_3MmFi�v弮�U�mܔ�:�@u�$�G0.B!e�;�W���V�L�z��4;N�eZ�����񗣈�a����c$we��`�Jc�i�Ȣ���������+�s��[{�s�v�\$B�N�2�\/{7Wboc��W�kO3��qr���jy;Ay`���b;�@�@��]@�Diu��<��g�ŶK���!T�ڰ�K��d�4�d�7����8�P�'ZI�+9���'�hU�gcrL�kU�ɪ��a��̡�|P<���7�Y�N�V%:]�1T�J��	�8�޸9����*�\�SF���w�5z�����K.��\0���I�g��u .ԬJhu�r�e�c�VԹь�o+��B<�ºV�Z
�qz��]YƆq�mu��*��9EK�b��[��<D�W�j��Aښ��2;.Պ���:8[٣c�t�VI#�vsa�ua������Yףp�S~��'Lq��.��w_!;����OOF//T%�'Ws�gܧ82ͲT<�
幂�֟!yZ�M����O���Tl )���NI�!�4_�ܽ�I����x['�:j�e��C��. �r��T�Cn���j���;��f�;]%�۬�N��;�Cq�
���$ɮB��t�ʆ姢}!NI��ֈ�����p���b�Ĳ`�tl�����Ì��3R��-N2����B஘�������%-�����&5���c7��C��:�>bpu��b�塘PR�*�(�uӤ�k�ac_V�-s\���C�Y=ƞoP��4��8!Mf�=
����[3թ�M�Q��כW�mL]aIg+��{�.͘I����]{M�<�l4HNWw�*�n��ڗ���m�6�_r���PY��i�2s�u�Ƹ��ܱ"����:�"�^Q� ��齬�/�o�j��!u�[W6ij��ׯ����C9����vb4*�;{��|����o�Պ�'5���U��<@�0K3A3�Ɉ��9:�fr��ex��5ɸU���H�Z�ln	�l[�������)dMd#�KJ����</�3�_`�XS��	ҧh�BʻB�Wf��Z��%q�\:������F��2c����7,�:1q����򯣎�Ӻ��+H�7�=���J'��n��j#{*+m�r��uh��<o7km�	��f�0�&�a&���u7y���V��E�)!��ًI����rJ�̼D0��c}�9�p�E���mB�%Ijޑ�;���:�
nZ�ќ<��wcΗ�7*PɣQ�
��\+&�����V��e�v^fIE��ᄀ�5�Q�*$��˅7y1��R�/�]KT*ţ-�gt��4��^�yڈ��]su�S��X �ٝ���s��89�w��ob�;� �A�5nUʺ��an�Eٺo*�5�`q��O����`;�w�b�b�7�i�Ɇ��[����1a��諮��6c�sp�d�]�c2(����S�����1uc`G˞|c�.���7�!YWܐ���Ufo*K�*�RSU�7�\�j����w� ����.#�kJ�vfe�\S5���k�rr��/6Wi�-I[�������M� ��٫����2�ToZp��i��D�;SC1���"v#�kMn�35`�o��b<ꂜ���+�1��{c_i�8�ʛ5�)�>�w�-%z�s'��m���Xw��C��JՉ D��9���#�zk����q��>�-�ڽ:!���2&�"ؼ�������*#� R�k�\�9st�E&��N�ގ���Gb�.:��ye��W�UAT  �P��A¬��("��*�~��k�1x��{ɼߴ9�:\�^��K�R\^��0� ��7�g��(�ǩ�>�Q�s� ���4��t��d�w��'&���ʘ�#�uF!�v�Pn�s�(��jG�	Y@:+��NXՑ����i�s��uy�q��1�K�8\��P�l8�^�[*G*ȳ9)`��;|��U����b����i�2�Ҭ��k��r��Fw{�c�o��Rӝ=2��(E�]~���w��# 2,I�-��n�dp�.�2]�%Ji�1%�!$���1�)��Ԑ�L�qv�&[	d��EQ�.-7j��B4�R��Y)�"$b�V
�u.S!)�q�H#.B�\��h��=�����[)�����������?����MT���W�r[DX.�WĥWC�UN��	�"�
s��(�O1� ��%�)f����^͈wc���+����rŷ�k���;��̤�se��5>S�d�p���~���e@��sH+O�C-��Y'6>�3�TH��s-B�\{�H������Q[k�Zu�^�xK~�V�`�ዼ����V���MS��腚��ۑ0���ԯb�sCCг~^�^�>@�8������=X��1�9�fZ¾�}�����. �/��v�wJ�l��R��O�l��}o�a������Q�:�Oz��@��+�����u�z��_K���Kw�6��cyI�^ٛ۵��!�9馶�c0���&V�󩣨��(d>�L�kju���y8(S�+KX�\l`���iyQ��&nnU�����ͺ�,�m\��z���fU�(�I�訷"�OZy�hu�Ӫ6�L9����!����P��њ�,n��,��=l�k*��ǹ�t-ߥ��A���껷���[�:���]S��jj��=�����+_s�-]��ԡS���ͼ�3�����Ya�T˵�{�k}��u�n��dg�Nz��g?K}3b/63W�Y�}��<O.ټ=Y�JH]�,Jِ��:����(�ڬ�R����ݥN�;�gY��ykmc�uI#����"ڥt�s6o��SiY��Zq@U<$�!^�j�]]cJm)t *}��՛�ww75��!Z{q�5}��|�m%�A�]5]�ݧ���z B��rl���F竽���1�;v�3��ˮC�)5X�fn�+43�_OW��n�%�!6�S�5mC����H����F\a���Wv�V�V�d3�� ��l��}5ة�[�`<���xAޏ�X���^��$��/���\�
��t���ԣc��17����	K$�"�aypa����{��n<�6�8'��fY���l�j�z�w]��%�u`giGgۗ�	�U ��[�]C���T��_i�`'�����2W�=v�>�z��5o=�)[S*ڻ�܉���W+��6ɞ��U�;����k�L�F��{<��
`mz��;w��U	|G	ݛ��s�a�=�)�m�yd� ���;�B*� ��F����!z��f�'zĳ����m�^�lO���]�y���<�e.���R|Z+	�[} ;}k&ҺWy���*�_J#(ފ6.�z���w��ͯ9xb�s�1=�ޅOg���D*X!!�-[q|)��%���ۡ�*��n3ns�Ɋ�꾿o\�Z	J�z��g7�Y̏Vs�������I�
�k�5������v�7Z.��&�cV���}N�J�W�bs����z��=�W����Kl��}�OuL�Ju��LЭ��ݓ�Ԃ&>���!wc���M,�d�z�con�Gs�`���²n	^]�=���0a�B������5j����ш��n�L]\o�1W��1�_��~��GR*� �qc���7)n��]L��Q-3Uq��u���VL2W��F�����!fg(+N^g�J$|�v�P�����폱�����.�q�
�Ό�w�s@&�yXsu��;Ap;]Kjц�[G�tvf
{mSy�+�mJ�Vn���%\��[Z��vj��F���!�
���N˺�+]kc颦�'�;�sG"(�^��0�{������R�꺩B�n��0�pW��0�y�c!"-��b�VS�˻��4D�i�
��ن�H���u�ې�*T��* 3&]�Z�E��f�2Jߒ���R�����(�cd�hqc���*���tť�
�]ՓXnб�j��c��2���ƢiUɒg�%�UhђܗHB�2�Fѥ`��RǊee�<�$�H
%
�F�I$�"�\�c�[K�B��	%ܵ��EH�4�B)�p�G$�u��L�a�M�Z"��˻. �j��%��PKcP�+F�%H�F�b
�Y�1��ӋdXő�KD�ʍA$���e����H*ńX�����t.�л?Wg�!%�����=�,��p����Ɩы��#J���g�w�E�z��~?���b�p��1��'�sq�D�t#�5>��9�����~�,�v���fń���"��hܑ���C[|$r���p�Ķ_�]�Ԏ�A��f���+������/s��N�"����Ы��/�ϊ���I���w�L�㪾��%��X~��2�b���v���y�I7�ҙ��7]�K��T��Xym.�N��U1��8{<M���o�s�|��:t�٘�o+�t����W����trrc8��L,��ʹ�Ç8�T0�|>�������u��V�c�vwL譫�{"����)\���.v��̉	a��"��z��IѼ2�������Ɣ��Wn���$�\��qU{+�8S������+�j[�ʃ1|+(ۺu�E"ߌ�ﲖ��E��Ny�R蓗q��
T��:��Ud!��������8���O܃��n�t�;�f��?�7:�Q�/�*��e
�Q�k�/O�uGƪ�	]@���[UXJ��e�,̪�vP�h�_3*�@�¨�W��MVR��!mu����Z@�E�R93��th��U�*��q���dJ�%�+U��z�P̜�=�UP��`Z�*�%Uy�h��E�Ua�<f��5UF���C�AXh����(���|ә�h4Pi
6���=(�_�q��(QģIZj��Pg����J�hJ���V��
��J�|H��+hQƃIU��S����5Dj�UAhPF�->HJ��T���W�<�h�UW���;��a*�4a���U�T"UZ�J4�ib#gނ�=�=�i~����1+�^Q�0a��2�S�aͳBv�ʸq�NWLV��yn<�+��Ȉ��	�zeP@A(����(�%Q����i(/��sݼn��!E�CMU����Pe�%P[T��5�|ּ���8�5(�P^a��HWR��J���Pj�5T-U	�W��|�>oeWZ�*��tJ��+mWƊ�T|B���VR�4��Z�J�n������Q��-u�A�(�Q�5AJ4�j� c0�4�Q(�J�1w&罝\h�	Tq�EW�)F�UU�U�-|�ٓ��b�¨�PF�-���R�j��A䪮��_��ky*��i��q*Ҫ��zB���U|h�Uj��h�����UTL�(�w��:���(��*�%i��|ϱ�*`���,��s�Q{/�~M��;rFO�7)^�=@�b�G��;����g��୷I.��G�_G�]���w DњϦr�}'���n�ޡ����\bpe�=�-h�0�R�&ی��(��v�)��:�=[[B�<��mx�]K.��2�J������F3�	���)��oוr���/7_��Ԕ=:�s�싳�<�9���|
 ʝP�}����D�|�}�\|f�!��ڌp��D������X�Ֆ5eĨ���r��ճ���y�����³��͚�i�Xtڬk�׳g,[Dr�K&<���'�%p{�;V\3����Z��Eh�"��8�ᢼ%0Cx�6�t�r��k�y��޷$��24Έ�rϾ�I����
���f�sȍ�]V��!R�����E�t0u�&xV�7���%���o�e�`KC�r���i�k����TH�U��.��:e���tA�}�0j��q��B�(ߌ�:�|���<�GO��;-8m��՜�/�}�V酇_�Md��voG�q'
�,r�r
����R���ڐD��u�R��Z�9怉����f:.�������ʴ�g���}��0{+���3��b��9"la�ʴ]%;�g	i��u!�=�9֖"C!\�@lg9�[�2��\�:y�o~DG����f.>���sՔ����v!�ޛ�R����WY�CɌ�nL���p�͜��R}���vVF�J����u�0�zg�Q�ˡu~��\��eA'dG��g��93T'.�����Y���No��d��`յ�����>� ����fʵt)�ۭͮ�u�v޴��S�;�*_�f0���p����%ׂ&��k����l�l\� :�{y���W�x�D��^�`V��������S8���)���T�T!�eÜ�|�����N�f�\�*��N���������f���8+�����+ʻ�Pw�<�q����ShOJ[y�4��;��K�bH�k�yŗ�a�"��]�0\(Y��Ǒ`/f�4�&�hD�.�$]�e�t��wB;�v�U�,�c��Z��X�5��)� Ù,���d�MJDN�]����Sr+Tݖ�!yPm5�)V2�U���:�f��آ�&~�[�@�Q
�b���g0�����W:bE�Ҭy�ӆ�F�*ʍb�.�Ue��$H�b��*��)UPiZbAA$�\��V$�$��Va�����$�K�)��J�1���KDqE1�5kL5�0Ҁ�KE��bA��2JQ��Pĉi)���2�b]��܅ĉ-e����ŶDEqql�-�H��K�"���>������VwZ��ԸN.��V"h�{����f
�f������'���Y�&��ff9�ne۠��_��q��dԯ�X^@�@�r�*"uM�8U���3�E����l�����Ձ�'/���k�P�7:$b̖��_�P�7�ۏ��B������o��}|-Ub��54G[VV���HQs�"��K�+H��D{а��-7A�eɎ�_fi��btx_no�ϭR�or�\��&�]w��Ex��k'��\ƽ�s}�s%�X�+tWqZ7:Y�ٕ�ι�3�f���vEv�@�+�:�j�Mހ�g�r���_]�x�qfثW�������� a�'����[Y���{������6"�6�h�;����Ư���w�aAm�J�>�,�˒������}�����HSq�ѳ|����I�څnS���P�C@t�P!����5>XV\!�/2&�C̞\�����Z�D���쩥W�kzU�ս&�����[Ρ;��r$�9����=꯫�+�u��~�K�<���۴�ꈲ��*K�xm�!4��,Vu�=t��E�SU7�����w��81ya� ��UG��צw�o�e�����ި�N�o0!�NT����D	�X��^}]=���k�5G�S�=?g���$��_o^�į�~G��Yϴ��C���=z�VA��M��p+zk��N��K.��כ�\�Z����)��\��1�&�)%_�.-B�m$F��33ٕ*��}�9�}��Ѫ3+!~�� ��\�: mD����9�p�F oǑ\oj"�'R:O|��x��s�c�X�/WT��t=��}�T}���}U�7�g�F���o�\bV>�=���u-Լ�0�r�q}�Qs>�ou/j�]{j(�i�-.�y������T'�BiWt.��k�Ihv�^S 0����[}����7 <ۭ
��tiVG�v�@h��"�ݻ����f�X�b�%�&p(��Wd���R�����z#������b_���JQ�3��.>e�+�څjU�0<9�c��t������g��~�q�s��a�FW�&L.�,rV��*q~�S��ܒ�U��\GZ�����D��m$^LĬ����Ok�b�5��j��d���5�G<��ʕG���o_r�{9�b	n��q��L���"#�9��d����c�C:���㺨f�����`]�*h�]�Z��X���1+�����������X��)�h�\Fd��'��l*>�&�O�܎�^6|�W�k/�켙��PP��X�i�͉[^*s��uV�C��#ޏ<��U��+�Û]�S+��Ps��N�>����g�>�7�/31�"��4$cc:��� �
�H�u��5��׋ ���%v�d�,�ބ��E�"�>M�%;�Z�e3cr�w�-�pw_,�n�A#��NX$�f�Ka����{�����p���.���7�G��o;Q���s�-���+9���y� 9L�Q���m�nM���-Hڬ7�_~�p�u���������Q���E�l�F9�[�ˀW�Qg�CVA�����=�gs{f���mfب�(�z���e���w��U�b� ���<�:.��\��T9X�8�5f#x��:6�(�rU���n�7�}k�Wwɣ$��Oq���x��`͍6�T��뙭ej�вK��|�L� t��W"F6�i�[H���ѽ¬1���iC����!��b�ƁX,�t�|�X����U�juu��� ��=��r��$�X�jڬ��s�nC�uL=��� Y��9Z��1z(���H�h:T��+*BjF�	p�^F�m)yldqG��L�y��"����"���j��]�yo-X^wia��T���X@L7�u���L���ߕ�!Q,4^dU�oV��B���t4e&�xn�Z�Ɣ�+&2����YR�|����R67��v� �na�K�	�U� �]�\nI���˵e�w� �EȶH�DV�nZ��n�M ��*[�P�Z��-��jԱ$��D�\%(��d��d"�ܩ���rȷV*��V�r�]����dE-c&%�ʄ���-$�"��R)!wvF�5%�c.�H�%�.�F]�2\����y~}��+�_b�ܖmtZ�A~ޏDD'�o��{�*V��T/�f:���`��N=�G������>Ц��������O�@e�ק�F�2���J�^u]���#�b��
�Y�&��=�a�b���h�fS��	�s:�ѳZ����Z�eä��x�w�m�C!L^ŏ�X/�5��C\z�P����κҍIw}]�c�%]җ|ܼ�s�CZ� �>�@�T�U9������k������O�\�]�r5��'wc��O�掴Gn7:h�řk	��w��iCi��ɜ{�:�r�!�^�B�4||G��X7�rw��pԆ��+(ZT������ޡ���[�x��0��}�$���g���}�����cQ�C��I��{�����v琝ŕ��Y����T�1���Wuƙ;3����}ª�Z9}��#{BP�yXwǾ���_W��w>~>jQ�K1*'s��z�k��0��)�8}N8jp������ي�4G�īܶ�^"��6�̽w~m��ٚlvѦ5��y=�Y���{��J�6�Ʈ��޵lϯ�s��O4c������[k��ze��C��׮ZR�bːÍ�\�˚��{P�b��|�Z�p��?��������3��̰�ª��k���b�?�t�Q'�K,?4���A_|�-�*�=f��G���E�2j�䮔�tr���G��A�ʦ=�}0"r{�><x�����篜�������\�}�Z�hx��\C�Q�W�Ofb�:���9��]]Tn����_D`@�i:�*&�ݦ��>��<�n�ɪܨ� �jv֤mM��5�gVu6�p�Zg9�˘�h<'�c���s4�7�[�6״s��x�مK�������c)�Ͷ�6�&�2�Ҟ�|��e��靨rRt��vN��u��-w%�H�xm�,�8� ����G��ݻL'o�|t�V���������.}umnBve�%hM6׵+���5��M�\���ᧈ^eayz�L���;���Yv���C~�w���R�:��O\ni^�y���o�0��z��h���>��{�;~��&w�=J�"hNY���9�WT��³���UX���w,NxV�wj�SO7k~������c]k	��4�u�h}|P�Xk�hy�V.�Ϳ�V{�9�	P|Y�.WW(��f�g|��itM�RY�sWg���9[��㉴<�^�^�����e5ۑ�5����u"'�b�̬$bz��e��͙M�H��r��je�����P��놭�HM�-��g���6�Z�8�L��29�^���]��q���y2�p�Ow�h����Ĭ4���C<��y��bڴ�/��[��{�^_=�wߛ�����R!�& A.����G�V՝�cÅx_��Z*��5{�Y�]��^.0wi8 7yE����s;nl��Y����.�jR�����+Eh�+D�^0ct��
��z�
�����OM<��%
� tx�����*V�"Ņ`�k�̏e��Z�G�J5�s�8�c.�)z��y2�2��3��V�W!�J3�^cQ-SP���s3-��OS.��i���7��<��*��K..c2��e�&VY�q��*�ZX�<��;�����X��\`���쎁�g�o>���S��y���\���ވ��w�2��ϲc'�^����Z��|�h��7�Y�Z�M>t"�X(yc��L|�`��[Zp},�ႰS��K8j�\<.*�޼_A�s^�霡ִ��&[�:�'p�&{��o�nܮN�3��3�ǽ�_��X�8��6��۞�r9���'�<ַ�(�Z& q��X�Mrg���д0�a�O'����L�&�z�+(h���T{zs����o����YW�G..p����-�Ҵ�3�;��?

���4|��N�ݵ���Y�۴�����j`ў1��|kY�N�i�i�\I�<�x��+�.�2��r0��F���h�����ALEi�7��&^&br��S���N���� qZ7ه�ݚT�؞ԯ�h�9N5�S]�^�y��o�݋Jh�i�ɗLNIw�o%�|����D�ޡ��(��n��8�
�LR��X��\K�y<��ę���S��й",��"ur�w(���}_}Ny�*�~{���e6����ws$��ZcX���78��ˮ��/�7�>�4��i�SM]�a���_JX���g��c�+ ��/-q��ۭk�Ώ4�fay��Vw���[��y����!��G1*��xco��]�=Cb�����q2�U�S��L��`�4l��@I��޾�i:�[j��.J2߳u��q���ekWe��G��] �Y+���<`����e�L�nB5�,�eKrYZ1��!�0��k��E��᣶�� o2&8�
�![�"�x��_'z�`bZ��=�9��O�% &X����Vmn�ըǰ� ݮe�tE�Eo�j�w�bP��vˡ"'"P�fe#�;'6{F �p�l	ͬ� ��1u�\�gVi�WrV\}[�E*,\��Yi۬�YnM�1[��-��.�u�T���V�腦�i5�5�Br0��Ү��5���>��n�Su�ţ�=�����oX��v�,`V�5���wc�\�c��#��u��=��Ru���[c@�}u=��f�j_b9YV1��E����}�Qk�hn������;K���"깅@�� U0�sU�ϕX�u2�s�q{�w�}F27B���/���TKnK�"$cH(�*[�����&!is�I2���e�d��ȵw%ݭ8���1u��I)d�����[xK�����.!%�D��w)��7��f�5�,q1q�Ť�$�	wR����F�d���h�	""�剖Dł�k8���ݤU�.���X��\!p��B9�a�_�k����}��S[�
�V�8/ע#�X�_�S����Ɠ����3,��u���6�&f[4F�Ӆ�ד\tMw���q܇��J˶��5��	�ƶ;Os�y�ea�i&[��P֡������wwKV��z���{yN�nCP���z��-�����Z%�n;:�j<kW*c0�q{z�&s��S���`kWZ�<���ӎu���|�䘔ds��c	�I����or�fL�I\�O{��/��J��;�u3� P(����vco�Vf��Q���%�����_}�}��uxz�;�|���a��{KM3��H��A��PX|~4>������,������X�)�Uc��ȯ��,A��?0����0k���=��a��ͺk��)]���|δ)����k7je6�+�����l|G�^ա�W���UR�Ⴛ�|��!j�v��rJΥ[5�M_�o�8�Zq,|��~�u��o��yJWn��J
�X�\�$vl�����W���j���t��{�
�ݒ>�����sn�u�)�m��7�Y���3��-�|���W��!����chG��{4�"V�զ����x�N�e�e뷆���I��b��LE:ۗ�]zVu&ݦ�~]mu�C�k^k��1�r�ԯ߷���9�XDÄ7�h�Ѭٗ3V�]1b��hb����i�K��̭'�\<�0��Ξ�����ƍ4[n;r5oyƱ<l㣔kNW�n$�U���R�}'T�]O��q��Gw�P��3�Dz#�4�������aP�!�_%sz���{Υu���L7�ִ����x4sVq�JTL��6��5�o�ޜT˔�ɫ-!��m�w�f�btL9v���m�h�a=Q��û�C�w8�箭�3)�ōK5h��F��)㨍�e
�>���6ۖc����.��^��8�e�Z�ֹ�Y=8�Ξ�U����L�Q܏�|WR�_�@����{(	jK����+v�maPMjF)A����������ٔ�m#����[�>�~�9�k����C㖭ÕI���G�z�Ẓrpպ}��g�;��Ǯ��"�Н�hiƻ�{::ц�JV��������^���(�ky��}���k��8�۲��8�2�:Cw^ק���q�ð���{w�×�_s�36D"�,�G�ˮ�c�ߟi���W�Mh�7O �4��O�d�̴��2h]ܳi'\,��rfCu�s'D�l�}UU�zb�����¥�6^qz~n�w��M�J�'��ZMt���>�����똳ɤZˆ�L4�=��9��=��2�L;�&���	��`�ٔ�Yī�C�g�םր+Y�>������T[5�;>�d?z��,Szj��r�����h��[KK��}����qu����)��v�.��=���j�
i�!���qI�8|���״������xUe������ک6#'pSwD�-�u�zc��;���*�2t��T~vi���^�,۴�5+�ƻ�<J����&'�:E��v_��;�7m9��cCp�i<N.�>��vlm||E!H}����9�'�#ou��@�Dm�X����q�l)�J�"���P����7��]�H']�t�"WhvY��w��sP�湘i桍Ku�V�x��]䩈m[v�xךơ�Cnuٛ��g]L5�5�2��+�+7B������+j�覶��\\s�H̱�/a(5{�\��z!n=�C�~Y��r�~fV#����Lcw{�bk���L&^5�2�<���9ل�Lù���<�}���kcXB���~�q45�vw3���-s3M[XI�XE7�i���W�f�=ܭ4��6���7�{�^���_5|�\��ѫB\=3����|��5��<��	���w��lK��g!ם�ӎ�æ��s��u���>|����M|9u>b�p�ߏ=�g�e@s�0o��[��es|.wDzs3������?B��߻���>O&�c�F&�$������ζe8�5�C�r�n�5}��e:��n��ܬ�B����ؾWa�}W����*�*
��2��nȑ���sfS�%�M�8����y4��!.�o���Q�9w������1�bQʐ�}͛����y����TƠb�X&�ҩ�X>�!�3�B����s���COu8�j��m#@����^񩼩/m�r`��j��1x,�ΕF%���`Y�冭+������m\"�Ծ���At�'ue�%� ob��QìAƹ�X�KZ<��]��jΑ�_9�Er '�v�nz�g��|����cO����c~�vz�A�b*u�UqM�7Luˠ����z�p� Y�즪/]�p�l�C|���.m�]�9T�
tќX�:�ͽ�(7���H��OQ���t�t�5��Lc$K�1��r���Kn�x���C�+P��K]��2�[�u[�V�px:���D�/�ě$W�Y|��ٺ��n�r�o��r��J<6�0��ڭ�b�m�NK�E�M,����j�.�S�(��(;M<�:Sn�4����Tĺ���h�B�0E� |�{{u9�yB��^�����1w�[ޕ��� �	\K��FK��ToF��>��ʱm������}i�;{:,�N��ڵ�4,����턕��a��--�z�K(�b:O���F�x�z�5문����A�	`���4�i���}R�j<9�cO_]�0�a���L=ڻ�����D3`�
�:�y���zH�U9HWJ����C���(PY�g�Y%�H��0�n�wq��d.�6�r�Za.�3�S�QU�RT��d���cqm-��"�4�̎ �Y�F�.[a���bA[�����Ӌ�"��*Ԑ�[K�wQI"7wuD�˕dL1/R��q%(�Eiq+-�a�!�ʲ�Y	���nTQ�2%Ȉ��5��w�OLV����]���	H���G-}�!~��2> �<oB�Z��w����Y|#M��Qh��<�$�TS�Ε0F����g��Kǭ��#4{�//gPE]I���#H��x��I��<q��u�&�^.�h�9蒥�9�6����q��Wy��2�t�VV����Bi�r�t�.��z"�e�C��;�a�Ϩ����k셓|w`ظ��ܠ��e(����%/+k�,�iX]��v����o8���M؋���vR�
 {�4K}c�i�y��qh��)�o�{m�]���l��n=����M&��~���*�r^��!Xp�25�̱����WJX�7����|�H�s����5k��9��US�˿-^	��(���ha������s���U�_h~�9S� s�/.Z"{wG�%T��/��0reip�=��W/o�[���y=|n��M*�#�ôg����cϙ�ȀBZ��MA>�G2��/Eg����7yO=�yҿB��>1�_j�u=>��0c�����Ug��ӽ�"[bb�T:L]��"T�5\�)m?��a��ܓ�E4r:�5͑�:J��6���!�n�Q���^8��v���v�LQ��bb6�v/	W�Vv|��sy�|�ŉz��"k�7��oc=ّ]d�����g.ɤ�_��mk}�f&,��ئ�������f��>j7x_p����{��j��j�u-T��m�� �^��M΅����:�,�6,t���Z�,��uA�_U�)��M��,=�˵�`�w��fl��(Q��L���fQ6A�U����y��࠸�u\�E��wވ�@τ�U2����$�WYk�2��J2��λ�4��\��#Z\���i}�O\��5���sg�v��1�2�j�z&*h��RhCCo|*r�7���;]3��s
���e =O}*�;�cI�;��O�i�<��r�oZ�Z���eo}��\6��3
5jf�c�F��Y*��N�����Q"��Vl/�f�ph��1��	�l�p�@�m�*��&f�c�V��t�l:�2
j�Z�%��r�k���Ns2�s�+�y�{���E��`�6C.�����Z���k:��zT��~۷��Z�鎖���%���=�k.��8AJ���}�)��{6o��3�	�b�]驪΋�]�R��{�q������8[Zop��]{��Mu�4"f7�M���9�Y�M��0'��LJ��ٛ^x,���Gۊ�{�P��c��[�ջbP���(�k�+���9A&��h��gr==�}肓w_ۂ#>q���%�vD�;�{�
��Ӣ�S�: �ʙ���E��ܸ�	�ǛU�N��R��.�A���9��b�'vfT��b�Ѩ����K#��W�1@_�:�'M��V<�;xΞ�Ցۇ��j�P�oW�o�+��db�T�f�\��r�����������&W�?ex�~A"��r�ߊ����+.���|&X�X=<4w�&��k��l�qV�G�;=�����k�sԶ��\���F�40s���^�]c�>s���K9ڸr�1I�Aj�1έ���o����Ş��|��Z���H�T��pesӭ�e�YTè��L� *N,--�����M1�`��k��@�����чqȃ���ӯQc"�k���6�d��-�=��f�|�s���8v�[9l;�����{WӨ��t:�YLF�S�ko��\�gui+.bEM�����l4�GWJ��v�+{v�R�h��|��K�ێ�q]�٭o	��cA��̫r�V���[N[Snu#�o�P  ���x.�Yc7��n��s8%�io�V)��
��+B����ۥq�ML�a*]1qn����\��,cB��F�YX�Î*�!��d"$PѬ�/˹)��x0;W�<ĐV(@�i$�����Xi#A�fL +�͠�	�*f�ݕ�]�`�Z�
�����kC�	�G���WF�KeIR�$J���DiPMb�RH��ڸ��M�H-�"���I�hV���cZ[DDAY*(ґ���24�*�!�
"���p�T�LH(#YKKZQ*��VvV��nq��!�lnڝxL3�����F'�Z:-��}=���	��q�I��+�"�35%O���8�{D�{
��Kæ1��!HۊUqI��\ůZ\6��a�����g��k�PF?_"#�9(%�c�ʶ�v�W*]����ĵ��#��Dcж�i�: �q�������=��%������L}�!��{�q�9�WZ�z󣔺�Ft�HJ��b���"�\iD��W�v�j$��V_�[�̢��{hx�Z��>�@j�Lx�,-u*3^��������\��3��T]2��}m�x�W
��G�q�F�Ыs,g����\�C�;նQ �ǂ�������� �ƠLI�6��YM�C�շ�h�gz���b؞\`�T�T)��~{���N���k�޳�^�0],V�xGENt��g��1���0�4�VT^vh���b�:#KctuV�Ł6�[�Z�D��VC֞����z$��N��:�7�u23��<Sg����ހj������g��������6��9s(D�=�\㲐4��т�e�!kݜGq޹�tĵª=V�v�k�K+r7o���Ⱥ��Cf��(Pn-�5N_n�f�4���gY�����;�yL]w{�oRS75��Q�J{�z,��0���ٹ�w�������u�& �G1�i#�l.�����Irk�P�t5G9�ЫBb/4��U���k&�{��>ʐ���[�i�N�Mv͇7����w�2ȧM��Q��Y�l�ӹ; �(�zy�	�5�T�ё�};�_��G�q���-E�z�}~ŗhtE�ջP�j9f��`@��*��ޱ�:'r*��J"��4;rr�Cϻj{�S�{*ʙ��af5��c'o�{�/���9��8s�/=��i��rɉޥ���s��G��g3+����:�
�M�*�p��O&d����t<��ݩ��zn�\��b��:��&��8RU@�a�2�{}��!�.�ר�쮓��8 U	E�7� :�ʴ*-=׏W�d����w��Xbz����l�>>$�a�\����^�W�д�Q�|7��z^d����S�o�����=Eg6�3����#�s��mJ��ۘϔWw�ka� g㪢�e{M��3x+�� O�d��*ƈ�b�N��8_3W!�^F�D���+M�a^)��c����U��:}���!X`�V"�Z�ҩ+�֭xza�,R/}O
�7Qv�6���ϻ���`�U��{7���զ��l)a;3�R̛�9�6�L\��p��Gofj|�sFuJ�ΗZ�;]�Dc-������N��=����Be_>*A*�Pd�|���AWn���ȼ��I꺬��W ��� y"�0�#iL0.�{��ih[O���,�\�Ľs�]���X�|�2��G���B?;�ѽ����z��`��w6�$�ƞ��B���]y"�s�W�z�tLŊ��ev��o��zl�ߔ8v���y��6<�u�H��Ɨq�B�%[W�ш?k����>}���^����y^�y[+�m�J�w��ŽI�R�e�U�8����RtE�l�DE�vN�wE�pVr�����a��{�Gr��\�և���C67f�APV_ڝݔ�r�}˝Lt	��v��:$�i��@��ȏ���˫Yf�,홆�tX�0m��s��e�;b�t�V	O5vڶ�����v6�bI���x[�ʎugb�yA�T���)�$�(�N!Gf
��r|�" �x)��7g2����$R!�*$Q��I*�$�#B�9.�*�N\��qQ�6)���H�	g ��vM�g&1T*�Q�1�Xܫ�լ�JO��,���gͦ�N�
�[@Rx"B�72���j	ȎU�J��B���(�w0ُ5f͙#NX
*��)��В�iZjIE'�[E\4��TF�RImZYr()lE�U�F���a�.8������R�ҋ%JZPA��b*��\��T0ƚU�0�e�#p����Q��$��+�ov��ו�L�9��8��S��b��2�X���ίhTk�%�d��&:z��4��o}�̓���ح�s�o�DH�"��G���TO5l�o��'i�x2=�=�C�zw1�I�^+u���0�(�ۥe1��Y�ㇺ��9_��X���v>�>����ǝ��n�oC �(~����c3��;�>���v�姆���鼺�$�͈M�1�t���F:�Oz���8�;U1�zy�B�}L��/��CU���DvS��]J�n��������{#Ff��VT�p�E5AԷ;\�����}�ł}�noZ�)ou�Q�K�8#ܹ)����k�hel�*��u���������� }��K�g�'q��������K5d�05���e�Ȼ������v*�fUҭ�u�I�-e�i��k�Sy#�+?+����Z�,g����g2r���r��bU:�Rƅ:�yn)$Wb��뭷o3��Ӎ�L��N�\Eʾ�j�n��.���Č�ⷵ�8wK2�)��<75j�Y:k���>6<ŉ�Q3j0���5<�qۥ�a��.�uZ;��'Ks��{�����Q���H�v�;�SΖdݪ��������C�l�}�)Ij�8���gG�B��g���Z���)���q��B	{]D��=�/��`c��������@G��i���/0�*P�`��TY�Z��3t6��\O�;��s
Z��+���/p�,��V��t���1U��ظ=��\7�>=W��d�ƽ��+�+bٝS_p/���:���2Xj�#�_�S�,�j�u�lM޵}�e������xQq�FE�N߹��u���=�)��8�oy$�Ԇإ�']�:�%ڰ�Xፊ��w�^�@6oJy��,Q:�9w�hQ[����NW U�y�]y炶�G�ts%on+X����rK퍮���#�ː���J�pz��{0�Tq�w�L34�����c�>�hm�r�z��1r�n��Ü�����VuK����,�	������h]���c�⮦�[�GG"�D�u�[X]�R��6�U��K99��r�r`�3ӥ%8I��ӝ���u��)�z��7z�St/-h4�%���(��AoL������3������\��7ѕ;���i�#|�``��Lf�e4u�Y�{�U���-�J\������
v�ti.�����4�H�#LY�Ay���[��m�-
�U��d�=ÈZ)Z�FR�.6�v�u<�Y���Sc��ȏ�����z���;��w1P�h\3r�]�nǇr{�-dnl���泜�eTdó�����8y� э�
y�Un����EYUڕ42/��.�:�c�u�֥�9w251sÜ�B��d#J:J���LpuRgR��J�����q��=Kv�
�-�)�~h��>zw��\�	�+����⒨�\�W����[>�Ub�y�=��Q6y�/;X�0�=�c)�x��N���؁����ϊU�M�~�3|�q�b��w�I���_V7��kۑ�j���c��3�	�͵��Q�xڇ7#Ջy��b����_s3��=�W��؅���FB,�3/��Y�D�ܳ(z��8C,k�r��@e�w �7YRh7��!Օ�+�n4p��E��U����=�7$��n��8�G�n]���v^�{���7\PT��������J�J��s�ű�Wt@�Ɋţ�Qc7����.���H�PƘ���O����2�ڈQ��ń�yB8���3YX�W+*�f���V�u�]�$!xl��0v��#V�) ����f�d:Mʹ2�&)Q�he�¯=�.r�HŴ�H@�Yt�$WF�������r�r7s%��#w-%����$aT�En����A������F֚c�"F�	\ ር8jjf?.�����z�eIPR�q,�	`]�\teD�~P�Vf��-���`Z�{2�L8K�3�c1vj��.�[ǻ^�h���=�6$[�hQmfW��N�{*X��<��Sa�R)ָaU�Ow�Z���.�C�Z=x�!q{;�"��@ǆ�{SLS`�s2��R$��ػf��x�txN]J��N�{v�grt��2E�9(����e������Ʈ����B�$�����qx�=�2��q)�-�U<t߹=����<���4�Ԃ�˺�g
�>�RnCp���1ve�q��ήv	��0m�F��rֽs��Iuma��*�y���wvFX��8kvG�g��m�S���
9�5NK��|����
��2:��R\xw�FB痤ۥ�~���_f\\�یfȡ�������*:�ЊlKY�*�&-?FG��,R�-�E��"3�|��a�6+,]%ƽr� �-\��TNTt �b�k�C�.�w���˫�E}�hP��k�-����B��Vka��[�&�3�s��2��r�n��8�N���t	�������%�����Uܠ�2�K�3|��7�=�ؒ���F;*q@)t/����41���+/:�T�����N ��V��� Cr�἞OwҧSꓢ]j��k�j|�z���vf�Vz=��Gu�N�$�&���_Gv ����OfL�h>rL�EF\�+�{K{���؝�o)O!�u�8��I��!��;�e�f�=]/��ޮřPD�������+=����g�)=,z\�BV�1�^#e	�k)�(��f;�šs�p�a-��tt(�,��+s��_E�0pLpu'pI'��
��`K����Ɍ�X	Ù�6�uı��Y9����M�GP7
�a��ө�x���7�l��5��f�8��2e;t��;���{�S�6�O;^�R�y�y�uJ]�^Iׯ����C�UV��d4X��EuĎ͐���`ڨ�MRK��u�F�%�����0���]{��أix^?8��YK�ӛ���\7v�y�%�"��/����c	��ty���w#���s���ׇ�����&'�Ǉ��*N��u�Sw�|��O=�2zQ�۬�aw�z�b��5�it���Np��ת;��d��v]v�sPIPhܜx�����H�@�|�|���8ܿ`�����ܸ=�;�]�Ʈri��Z�J^D�lXq���V�<8Vu��蒅�Luf��Z�Ni�k�9��	@��-I�1e2��Qȏ�ҫ��W�	ڛ�~9�z�U5t�K=Oݚ��S�ݾ�~�9{�*%Mu�:�s<ȭ�)��r_{���7
�><���,�E����u�{���+���l���ӕ{���������!uv��򩴷�|Zf���rKr�)vΠ�b�V������/��{��:�(��n����]8�^Ulh�r<�nxk����պ�;�t��,�jȧ���W��7�ng;u�l��.�S�Zl��@��2Gr_gC�����w�T�����/h�����k6V�w�Z���Lpֺ��u�@��>�̻���m+8E�4���R�и���|�%���,uY���:AfU���f�e!�d����g
z���vB�R�8ҍ2:e8u\����%�`�`I�� �k�S�R�IHȈ�Cv���{�V\L�f�O@�bk^���˯^*�iآ�ep��	/(�.�$��<Y�W5��K]�L�E��u2{��{}��ɵz���S��u�[�Wg��a\�`����o/]������#{�䣺�s���Ssl�``�m�r�N�NQ��s. -u�Ev����n�d���p�וy� ��O��;3Eb֛W�Q��i�Y���l
5�J�z+�7ys��+�K�Q���j�˦/�И2K������F�8�V��l�V�b�bLL&$���a#jB��^#B�r%�A�$#�kG��Q�d�č��A�FclE���ӊ��۶�L5vJ���Xф�-�E��|p�z�uQ�.�pr��W*�g�l�|"��u���<x������H��Y��a�k�q��ʳz���$Os�>Pf���nv�W+F�E�c��,�M���ǋ;�Q.�.�~�2�n(����AQ~)�n]�mp�ﻨ��븂I��Xi��� |{�z�>��0'r�9F����T�e��`�1�\Ϯa�ح����"V����R�9v����>���P��p	���u�D��#13��v�<q�K�c�ۂa���§�U����<�t�i�4�Yk����yo22y^ID�::䂸��ts_O)�^}r�P4wK�2h�=�������S��2����{�ǢsaW���GZY��밧DDD�o'��zN� �v�k²E�jJ�a&�C]�<�3s3�\T��3wүVWW)f���m�)��h�4r[�\�or���^����je�w�FjNf��\��e�&�	y�-,��.D��ڠ!ul�wxT�{gP�����Y��J�X��*��۲�|<:x��ǫH�k+��
!��/��z��Z��^��^�*`�&zLbh��/�	��J��Ή.���̾�Ӈ�wu
�ewK=�V���
���v���#*Y{a�ԯjx�[�rő���K�v��q��/'��У��51�i܊�n��7W��o"9qxs0Q����R`3��/D��ɓդ�a����Dm���ao=�VN7�{5G��ac�.���9B!u�(L��A��c�G�>�y�$5�*x
�����
ٝo9��mu�o�d)Ywhu��	s��5f���f�	��v̘�3k��X#�w��c�.Ů�Jܭ�B��^P��5-52�s��Jޡ�.-ĂH��4��d��*\�����(��y"' �s�ȱm1D�E�$�	��S/={2�r8�M�y�qA��o�{JV��95�X���k��T)m�z���+����9�I���4ܮ��H>��ܗg_
�i7s6���yݠ�\�E,��B]�1l7-`�0��n���7h����L��&�k�+�|���A[Q�{q���S��Df���{![��q��)w5w�]r�wK��gT��YX!�PM�����D�`�S�W.��|��?!*<*b�Sƭx��Tq����fN۞�,���upN�|���9+��~|{����#�׭��͹&��&�O.�i���|�����I&�½�����S0�bV��J�JvnXX�βs͹��j�L�u;�K�U��rY���7�m�6*1���H�BeԸ	�J��7���.��&MSu����jw�ʎ�����
�P�P��
;��rM�N˼cx����j{v����!J�;�����v���F��bz���E9��_��-�6w�M�g]#��_!�<6^�n�u�y�E˕m����ϼ����O�"����(�
*�a��
*���
 t
*��b�AtW��%LJ��A���>����z�� � �T "��0���vVcvҩ�G�*��WѬg� d�U9(�u}�[UAT ~�)~���g�ϻ������ ����Ε�e��ɟ��}�RU��p�F��h�pCz�8U�����@�K+�Ѽ�QT �G���G~�?O��J�h�Gꢨ� ?Ȧ�TU ��(�UY��?������W��W����?�H���������βW���C�(� 9��9����?)+�@��`�@�Ub��R��oJ>ƫ%J?�C%�A?�UI���V~Ϻ�4�����(q���e~����	_������� N��!�>��TȎ*�*����0�B��9U���VM}D6�R����&���}_
�C���QT }Eh!����>���}�>����(��߲W �}_��|��v��������W����?�~����+_���)�@]@�����G�h�E��~��W���Z1�	���ת�+t�?~��k�~��U.@�J2�~%}|��}W����_������ʪ�� ���Jy���R������
�\��C߻e��*�� 
 �Ie~�(� ?����� �L�h�~P"J����t~]Ю2
����Q��aUU@�G�Z��W�
���%�P}N��(��$��lj�4
���~���jP���U�]�+�ՈUwfr`��@���E@j��g�~��������� q����
j����}`}�����W�~�O�G�׏��>������~�����~���TW�������*?�U��(������1��%UP�ξ������UK�J$!E~_����?���� �_��k���������~߁�ҿ/��YGҾڪ�����Q�4lJ�]/��J����?#������|�gG�D���ܿ��q�7]<W�g��e}Y��� ?���(��@����7��`��n�'�Ҿ��+�����7�j}�2��W�Pf�?_�>Ɗh�*��ST�)>ª���u�O�}u���>�*�������B���U_��´VsN��r����;���&���Z��J����U������H�
�#��