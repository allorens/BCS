BZh91AY&SY�.��(_�@q����� ����bC��     7��j�5�L��	R3*�-i
1�h��P4�[V+k(jmT*�+ �P��d��[eH��d�5�%hV��>��66�[H٢3AkhUi�=�uf��f��V�F�`D$���d֛M�lֵ��lb�
[[j��6�E���Jf�����kZ����ɰ�U���Ֆ�fcfkM�*���3e�%�Kͭ�L�j�i�f֬ى�����̵R[Uiei�٩����۬���j5���|z�J�   ���kiV�6����6s]�uks�,�Q�C\�vm�TZ�[n��6͎�gV���9Q�mZ7s�iclۋ��ֶ�l�l�)4X͵�ֲ�&�Q�  n�Pt�n�f���;�����(  n\�(����F���S[  Psq�@ �n�Ҕ)��ۅ �z�z��RS6IE�QE-�V��  w;w��� �=� =Pq��iC�wU�� NwQM��=�  �Ʈ��(t������b�� � ﮞo �{y�X���H�����&� ��A� 9����Cx��� (W�x�d+�b{�7�)A���k� 3x��: h�x� P�x��� ���WU�]�6�m��a��i���o  Y۷��� 6  �L�F��B���p��Bn��*���ҕM۲���ht�ʸ  ;���  �^��6�[TƆ�V��Q�  �x: R�8
(H賭�	�0�m��:��l��`J �q� :, *�\��GN���%��ȩV�����R3�  ��� 
R��  �2��厀����]
PP;��4 V`����b� �u�Zu��#Z[dh5T��Y���    ^��  �q� ���Ϋ��� W5S (Ӯ *4` ( 7;Z[m,F2h���  �x �,  ۶�� �� "� # Lj�(�R�;�' �n��3���
�i��vu�ke��   }��N���  ��p n� 4��t��p t#@��4� �  FY@��   @AAL�%TF�4 � �#COi��Dh@  h241�L��T�� �� �?��	�  4 &��%�Rhiꞩ�@��20i������!44L)�1���@4ڍ�mѿ��V%�xm��#���Q��񪸧�һ�=z�x��y��/�ׯ�aPW��
�����p����?bE 9�$y?����#���c�� U����\���p U��=���p��UA_?c�?��~�9��졙C���L�S�2��`l��������l	� ;e�G�A�{e|0=��l�� �ʽ�/��{lʝ��l)�"vȝ�'l��*vS��;eN��T�;eN���{d���aN���{eN����
vȝ�l��;`N��G���l��v���l!� {d��@�;a:e�{a�C�@�;dOL��"v����;a� v��l�(v�XG�@�;e7l	� v��l�� v��C�P�;d�C��� v���l��"ye��P�;aN�C� ��+�(v���L��"v��l��vʝ��l{`�U�x½��
�Ȝd�{a�;d��E�{a>2e{e{`N�0�<e� �� ��
��S�@�W�PS�S��A�(l�l�l��l�� G� S� S�E��"��v�
v�
vȪv�
ye;a;a;e;`;d�'l��l l�l"l��T�xdE<0
v��T��
q�T�U����A�S�*l��l �l��l���D�@��D�{eN���=�l��"v�>S�T�;g��l��(v�=��l�� v���C�&A�;e���;d�C� �;g�Vd�C�@�;d�C�@�;X���_����������&Ƕ�W	�_��A0lcM[�k�
�Q�M���o��P{d�_?��D�����c�)�g3Ļ�c^��7UhdҘ��Qq��Ԝy%�X�����������@ ��1(�K����c� ���p�Ŗ�yuy���m9��Qdڎ�B46�d�A Ós	͖p� ;�\���D�U;� L�cT���lL�ܭ�v��w,�G��=Y6ِ����a�W��"�L%J���1Jŷ���{����i��ЏbC��/����+�i�	�H���)��df��V��RR���F׷��
rP%�Iy�7�\�S�+�sC2�Uv㎦]�R�02�,�z��X6�`y�ƌɶ�&���U�2�J]ۻq�hӑH,��X�JCm��#k�;L=t�aa���U�*f�߬�L���x��ݚ��nn�c\֜$k+iV�1�����3��1��O�m�n���\M<77hZ)`ZЉP�x��ݱC��B�4�R�Aֻ�xx=�y�K��V��IL�j�f\��Κ6�8�2�Lxe���;̓w�¶-ߌ
 ��
9`��@�E�[�m�ڲ�э�f��,�}d�����Ҽ�
��o�CY%f��e�ǳs.�#2MJ1�;
츅�:fkv�H0f����B��	�&��UsDz�
�O*�`������ǕJ�L��7Qܬb��n�S"�4j�i �ю�a��;6qZ�Ǵ��onbSUC�e �jV�Cə�7�V� ǖj��r���:��꣉��m:����{�ɺ1)���b� s*˕x��6�0�zձy��é��f�ڄ�b���n��b����S&i�w-��*�O6�r
�a� kim*�"y��
J���[�7e�o4��6�/1��٥Q�캷E�� ��r5�wP��1�٥S��d4nݳH���`n�5�$K�՚u�Yy���UlE���(+.F�H���ˁ��&��|�ݠ��E��tQv��Y��*��xz�(P�Jȳ��� �����7K�5�bB��l&��XT��"���fkK O1SШ9m���k�x-L��庆��*8��4��"�^�6��k[{RF�ͪ�r�;�]3Pk��n݌ja�7z�h�;d*�rK�`�X������A�R�G&������Q�{F���t[z"���ïL�f�곆
kJǘH7OPjᅗ�շ@֗�j�
H��7&ǖ�m�g
[�>ݮ9���L�N�5|sH,����Y\�۲
'�l����� dj��>g,p�k�	�[��w����Q����fT��iV�����>Z8m��42��E�y��gE�L]ܣ*�Ƶ�c��1�b��B];	�ڶ���֐)U��o��V�-�L!�@7��wL<���b%+za�-�ܩnV��q�V�������w�A�iըZ2��2�H���1�\,]�ݒ�^��`�b���@��U��So^���1eM�07�"[��.��q�n��bj�����*����h���Ym����e�[��v8޶y=l�[�˨�̥����oQ�?j�4dkZA8�ag�1m����ŸTܭ��x�Lb��n��/b5"u�R�����֦���n�SO��+I0U�R���v�m��nh�6b�Jh�zo*�#ui��SԔt)\t�а��r�e����;�E��ܨ"3r�:�[���f��7��� N=��,��`�Fti*�f��$5{e��0R��"��Sj�b�n�iR-DY��Eҭ���%D�n֗q���n��$����o\7]E�5s�q2f)j��������#����7��Xc��XJxZ���ܮ��)S��ۖ����]����AQM��P�ӬΧ�n�7��Ϯ�5�@H
I�(��[���A4��b7�L�f���c2�vH�2ʦ)����w��Ly{+vXx>ǐ��ư��ᬫ�o(��z�>@�wt7fk���dC4��`M�9�e�5�[Q��a�V����k:�2�j��{%�vݐ��V�^�1ȡC_4����n����b�����n�\�rZ��ٳX�©�sH����*�O��l5=řF�n���$���*��%�KAvN,9Ls,��:5Ym w~�D&/��.����Hc-�8��$HY��VZ��\YKsC�r�:*Qq���yYn-o�5"�Sˤwp���Xj"q6A����Mڬ]�JS6M�:�v�8��ַMM����wF/ݙM��I�顸5Cl��a3�Mw{5f�T����si�HTAJi�^��fѷR�ʔP�Z.��r���A)n��2�?���*7���زʑV1WQ��a��dZ�3鷷6�X���I7ZN���tj�N�p��Q=�cU�v���96�\�Л3���J_!���p7i�&�i8cBV�W�Er�I�]���6��v�
����dm�����n]nۢm�5�:�����#n��2P���'	���L�SKwS@�R�{Z�7[�*�A;5��Ԅ��3
�J:0�B��g�sN����n�6at�:���{��z^�c��4���j���h�ur@��&�#��ڰ�6��	�׹�+���s��ܖ�i�ʹ�8F�#�y���XR�^5��oqG��]x�0�R�+	��m��(-�.���yPܚ��Zc�之\�<��˕���H5Y�K�q�fl�ǒV����c�"�ge�0V�ІA�j������.��f�t�C)�H����W�骴��4ۖ��y�y���u-���L��r��0H��
ɹa�f=���.��/,�"��76��96J�	f��V��t�1����3v��4H�3�J���x�*�YR�7o,�1\U��R�%� �ۢ˼@�e�(aM��Ux�ۡ��)0�qԉH��Y*���^:w!.���X�(^���+u8��3e��a��4�/CY�(+%ip9o#�.�2��t0��kN��j�mf���٬�GbL�AsԋƉ�̅�eH�l�ԼQ�dk��iƎr�RK�;=z��GH��7P�C��x+��w�t��1 [5ʄ�5�i��2͟��h��QCZ�kV�����w����(�^�(��*iL[hTشA ��T���D��V5���;��:�w)���������n�c�m4Nixط���v�`:��t����%4�@�l�+t=P�`T�N��=���Y�Ϭ8��ed8�(ݘ�Ś���j�Dvw�N^A���KKe�4�3c�E=��i��ա�)�R˗L�nέ�C����Y`SO���v�i�Z�՜�)2���5k�WU>�ˌB�I�maO�X^AE����E����`晈K�*�Yߡd��{X\M�4Qv�2� �#ѩ�;%�`S���u �5��ryZ>����aa�l[f��ٕͦ�ͣ��#&��;t���DݙM��5�E4�[lݺ�Gmm]�
�e�8JD�V�8�#a�:���$��gE�޲z���e���w�3$�6^�E��"D̼�Z�͝�l=c^���Z��(PR�"�B�m-�2��-��":S1�e�qiI��L��3>����	�)��V5�!C+N�>:������[kV>��-�Mn[c�� ��Kө�A����h=i8���$)�������:�Ū��P����X2���� ����_e����[�!c�L�V����6�lo++:"	�nA�Z��;�M<yq'������n�*��蠉"�R��Y� U�"C��PM��a�r팵i�K�4�VR�cd@S/$�Oc)�7>1����D���Le�Zބd�ۛ�4�n������{GM�[�gpK����G(�KY��Z�æ�TvZou����S6�Ŷ�6���!Ќ*�Y#e��� �oaguT�q��S�����jp*Z��F*R�yi�փ�S�/r��]�yT�h"ȴ�qŎfHZ2�H,��I��J��W;�����Y�@[]��j����%f�-�+��<V̲����e���Ϟ26�ȉ�X�;yX-�i���v�snF�#�/INIwn^u���I���.��N"\���Ű��L�2�-�cK�8�;��Z}NưK���l�˦h��T9�5�ڏop0��6K�s�N�n3W��i���Rܘ��ƄZ5�B)H:�F�v�.�Wo�GoZr����ʸ�?����C0TU�ڄ�����ɢ���|4b��(n����E1�9�5�}��w(�-�7]�q7�T$z��PX'&k5Vج��Yz3�iVbS�)!w�.��r��)P;ؗ��@�d�k��z��o�O-�n��1�{�,&i<��-�T�p��j؀aV�Х8#�����bn峲�Sc�i�ΜQx4c�u��ͩM64���N��q�^�m�4TOPz�F���^U���q�0^�Y�������j� �EH)�V�"]�.f��wkQ�c8Q�B�D�+/#���K˚���T��ի�6H^n�)��jJ+��DV����#u��Y:��
�^Pe{VfZ���U�Ւؑ����V[�Q:!��ޗ��*�D�B'�Y����X�fo�'i`��l��ͱ��Uf��i��.�R(a"5��K9*,o\�J�L�в=�cs!��)��Sݗ�ٓ���5j�y�j�����ƥ�`\�/C�b]��yJ��B�Р�dn�^g4�'��Um�Lc3K�{P阢6����8$����`No5� ;�E�%��&�/b�	ѭ��w���13�D�U%	p��T/M�]nar6�ܢ˲�^Ԛc��<DX6~�E0�,t�ǫ`U�*[+��4��gU;r���op�kEk�YGN�$���7>R�J�:F�n�⛷7��L�b�BA��hL��n��"��*���cV�z^�k�N�`G+V�I$P�l������̔��*�ƚ!X����#6��^5t��emEq2$2���w[x
���)fC�V��a-MwVr��V��Zˣ���o[Gr��-�@�$��$^V2�wcU�N�ͣm�h�-U��;�QC[�l���1�=&,[��	skH���r�Ov��V���y�
�6l�qd�A(nõ������J��0�p�4)3En����/k!T��#�W��Ʒ(d� ��9{(c	M?l��M^�1����K�k�h���Ӗ�\o3W5n�=���*M��[2[a9��Ge+�֬;�6(+j��Z�愌���aT�t�3cE���90�7s0�)2n=�Swip	&�l o��"�h���Yj��
�e�
�6���P1:Nj�U�V�i3��۳2��6�3%Ԭݹt��y.�d�)��
y�"Uq�:���RaR�ئ3�^�%ԚI2+�e�"�^�(,l)*<�9��ln�ʹ3FA���29���ʑ$�]1j�ʕ�I�\�P�J*Q�����W���9��щ�8�R��w��̈Ĭ�T�V3vG� �#^$]���ϑܤ�9��f�A{7&S�;X���E��f�O>[�M �k���i��i�)�t�mk�E6���7[ lO����B.�K��P�m���y��V��ʉS������#���Z���z���n�#LYR�"�ѥB�j֗�U%��E���<��\�����&n��F��Ӕ���,Y.R���4��^d�n2�7Y�P��X����ְS�����b��=�hz��Ap]dp3F��5�HAH�6��jP�%��n;�V���̘)j״r�9D덄�X��*EM`��*���ѻ3;b�5�]�5u^U�X���L֛���-��.M��h�Fa�]��#���Hni����M,�J��/�"��d�4��O��Q�	���Kc��r�;��|�����ǵ�;2A{E��Fݬ�%�"��
����cz����n�#T��2eVZܻ�d���P)�
�����4�B�����Q�h���v`�! d��|���h�ޗ�,��P�v��S�y��7Y��uj����HOI�SwR2��&���KL5���Y9�Q�����ё�5�m+�/i�
�O�^Z�e�ة�G��nM�^�[����u��`��G]��d��j�ݭ8��w~;*��r4�Z�Z~�7�4�A�B麐�.!�(��'Wt�/NQͻ�L9��د�l$4�I� u��ָ�ee��.`��S��$��=f����n��s\7�u�G�')	m��ɦ(�ht���l�5�^�K����l�E�X�Q��Tr+���ݽ��Q�)����nK�	t��M��"È9��HQM�o�Q<V|�k���cK0�4�=������R�X8��m@���� Vɽ�Y3e�Βb��nc��Lî�l�����R��SV����"b�iɘ�gv2љ��xV�kj�sT۬+jij��y�z>va��fQ�n��F�* �W�Ѭ��&��0ia�b��y-m�P���zA̛[H&f���Z�S#��m"r�ʷ����Mn������lL?1� �Ӗ��7,ޡ������R�0��Ԇ��Ø%��rѲθ��e�Ҹ]Z�7u��P���  $6ѝ�X��9� $��H�Jt�K�*s5��1zW�t�I<(�� X8樢V�[D�p%+�yf.Ib�q��PZf��3Y|c/Od��_r-[Mi��MD豔R�N����)���=$8�]����R9�l�H���&}�;n�"e��̩7(���S'.�;��ڨ��R,�c�Nk�3�e���	��+�k,�-�DU�B�l�{ǐz&� �q� �ѕw�� "�E��b���W�VP.
�dhV�Df�a$>:�ih�:����p���LI4���&e"\x0��8C}Fp�* pY�`$ɶ���6ӿL�M�FH���W�}�x� ������`����?/��՜����Ɇ2���
I�VI�I�N`�*�Y�$��G_V���d�u������.�N����7f>�d���N)�[&�]��̔.6nT;S]��I�8z,���.�Z5H.��MfMv	��[�0+Z�a��*�.�,��W ���궊;T�Lv++�j$u�\��RR$�.d`t�\�܄Ө��Y�L��$��+�خ��.��Cy�{��P��aP
�M� �Rݗ�C�@��0�,�]�C4�3F�s��̡%��R/��n:2�d<���o+!��u;����y첯�:�6��a�;���!�J}�[,g�m�E��174����+J���u*��f���&��F���H�M��bN������8��7�䣹����Ջ��V¥�1|:f4�+b�M��֙x��\��T�V�4V�w���8Ju4��+jp9 ��;ٝ�r����|�i��$�z�s��R�u�m��F�����-��.^S�0�rU���6Sk^@�f�`;lH�k!t��UL(۾U�˚9���Ǧ������"���;/��*�wXռ�`ܼ�k2���ۧ�	�o���v6�1�L�3���Մ�\��=ƴ9b�@��Z%
82��"�.fT�y��A;'�����ӭ<��ݠn�7U�Of���䎴C��t�;�r���h��x^��n�Y���f�hĜ�Iá��4�����+�6�!\Sӑ��m��xF���b�gS�_Q�`a�|����_
�L�U��G�֋G_�lv6��+u�靍t��6����ݣ�\����2�Y����VM��/qΣ�#w36(��ׇ�����M	��V�9iKN�;��LL� S#Xy���>HG+��R�Ai�oSjc�uV�XNjp��+�,W'���/�w7r��)�0�r�:c/(��oEO`X®=w8�_z����d(�;�%U�")5g}�{�3C8�"�57��7rW+3g_vf�O���3!����¢yn� �z���Ҳ��]�R+7��#9� 8l3{δ�f$k3����Qz�����Y[֝�������Y��4��i�;BNN����Q䮮�M�c��I�ۏ]YF��mC��i��]&0w��WR<���Fnc��YV�"e;f�e╝�ip�Y֛m�(��"�O\���;4���z {�-�q�/3��e�N�j>RX7|M�{u�Zk��j-�Y"��r]�
,�`���**�Z�Ou7n.U󊻰_O�NmZ.ͱHSr4�����sa�ɻ�['�ۗt1�Mޮ.j!*m��.�׶�L�n��Ar��� �L�"�)���j9(��]r�����m��2X'�,f��n$	��yn%#�؈ҳ������ɶ�j�^0��$W|���q[�����a#��R�a(�\ܛ�8�zr�H�������+wvV�/�=���,k�Q�%�ua��3R��rN�ۃ���\�ɪ39X�jp10�C/2��r�s��)�|�*���BWvjՖ'wV�7�܁ȝ�k����l�z$��=�C�-s�w{����6u�Uj���v~B����I�u,HC��:�XhodE�^P�q%.ga��V_7D-��G5��$��K�����I1N���q��u�RR��Y@��N�J��r5��v�af�P�e4�j6��݉)u<��+�K�MI4Ɛ-��uئH��B��g��5���غ�{��-e@�)WK�4��I�)��-J�i]
��E:u]�1.�	���6H�7d�����>魊�L&u�٥K���l0�v���� �e��y\XkY���ԥ6R�F��!	+8wG5;��)g����i��w�����趸��:9��O�avo�v_>��(�&��rY̎���`)������CZ�7o9|{8�v<���*R�v�4b�p��'�;��{����w9wәc%����4رD/p�_3�0��u�fF�R�ڷ	]���+y{��;;3��PnS�pet��[���|�Q�
�3wX"�$FX'�3;���ܢ E�oD��ĻF��h�[�R���$�j����nB���hj:��E�t⭷g5<|�R�ZD#��Y�*vų��yr��T+r�E���6QH:�`��l�D��&�=��A�\rH"����*@�QJ{��\��5��+�I4K�B����� ɯ�<�B��K/3�};�r����݅�n�L��(�j3��#՗�[��%�y�#�N>�����[�ڛ��l�Q=�6��BS�EU�Ei����t�6���ɹ1Vl�3�޻G�OТ��pי6�=qu����}��ڸ�׭�W<��p�{I���A��^���]Yz�\7�<Q���sH�9{p�J�_V�f���֎�F�8Gz%�yg�8�c�7}��k�I�\&ܭ�JN7	.".���ң���X��q�v�D ��K��V�S�ɍ֩W��_P�CE.fJz}�1�
�{G����l���e"RG�+�5.r<R��n(�y����/��
���2&uB�!���T:�Y�+�T7iQk���Hfl���v�rR�L՜�fU��;˅��<�<7��*a$4	W%e�/]:s�p_C+���gBVT��B�+��G�����q�y��%�b�T�cщ�����$���]�� OcF���w:}G�Y��,�P�� ���t4�VU�,� 7W��i�^a쵱�}Ƶ�u)�T�Ǣ͹��V������π�޾�h�ù����G,�N��ƛ`�ϓ�k�7���=�<��m��N�`��y��]un�SOe�o�b�k�G�oF7�%v3�υg��d��3f�Ux���{<�[�Ϩ��]]qŕ�oK��ʹ�"⻼����zA0�RfK� zr:t�Y����g���ҭ�+yP={�@4�gQ�j	5��zB][���E�zt�b<�n�T��'L���׸bѽ�$�Uy>�ީ�������0^�D\H����׸-�V�%m�8nu�h&�u��X�%�麢���o]�×��بӴ-}��-���c�����R����^CtCأZ�D-�0�9$��Z)�6y%���϶���v��;���,42���/�L>Hef0��fH�q-B�Bb�9v��[b���Y#�m����jw�G+,�qK�OF�̶��XV=f[4�p�a��� K���!�E{�8Y�F��
�6_nf|~�y��ju;)^�l���x��$�'H/gK��F��]�զo�WDi�Q���jדT ���I�O(��m\�Ֆ~ݨL)��R�L��Eƾ�U��t9_T�K�rֱ��4i�j�엊̎Q�/^��V��V����6c*���[����z8��C&�#�C���5,ZFtj�]f������F:X�8b����uŉiY�ᶸM��HM�������y"�v1����p�]�U��b"r5�^�8nU�T����rw6�X����9ѕ���!k.��	�Q�$䚇_e,:�=�ˬX5^\���ف8/B�Ylj{�y���`�\T��Sv��s{��f�F�M���2#%�Ƒ[Kk��Z-�x�@�������w1�S!u�CvU�2�iv5N�LwKI��h�T7X�yfD���8��ld��޷�7��2]ֶ��^��9���e3�I05�yu��>Ҭ`���ӡ�Aq�Wh%Ō�l����l-T�޺�xl=�f�n�_G%
��������&����&BeS�rڏv����B>0�3MLձ�\0&�ѕ��N��:V#�:�n�:ڶ�۹}�L�@9S���yƥoP�,���\v���O�Z�Kǽ\���}м�Do��T�˱ʀHeoW�Tz��\�+���'�r�k��ha��u��8������sc�9'L���5p��ZÙn_$�%�,i��׳*��ݍ����9�\��G
�&^U�#�7Io]����ء����-ϝ�Eݵ�w���Mso�{��ˊ�
ˤi�&>;Ko\�Np�|��K�p��	w��Ԫ{}S�]S��	�����v��_ �ovN����kʘ;Gy����͈S�Z$u20`(��0��Y3��6�Dd�9�϶�U��M,���X��r$�ֳ���	���;���x����±D�9�,oQ��5c���j>_I�Z�N�[����C|�S��,�Er.�:7~��t�k2��^�zj̸[r駝'n8e&tnӍ����q`i��.;u���XBltѓ(��MWs,�9+��ݽ��i��W�)����&�X�6𓨆ހ�q'9�sy]i���Z7;��9Lˀ KJ�k%��9vX�ͣ3����ü���3:,C:R���ca�࣎@x�;��1���T'm����U�����6h)o&��9ܶ��*!71�6+��Rq�V�nnӒj��S�2a+M�����:;��-�骮Ф��+m.,����%�z��8Z�r�sX[��l��-�8K<��]��us�;!�
SP��SP��hUk*B�OZnni��%�mV���pq�嗑Ȑ�(�5%w�� �ݛ�Q1T����7W@�_Z�yI��ֵ�C3</�̅i5՚����o�];�;N�+VԬz�\�8�)�;3D�~�������u������+<�x�<	�4�W���f*��w`��컘gb���tB�D��y�djk��!����쭒��y�|}6��u�$�����9*��NF�;A5���i:/�-oՄo�nS��P�d�+wvdw�V	��Ew��斪�8��K&��w��æ
մ�1� :'=�����^3�ָ�3S�ǫ�t���c}�m�ċ���+*jU5���Y&S�O��g!v�����a�x�G�}��;��p�.�{;�9^��̈`U���o���o�LZ�A�t蛥�`�U,S��>�P�r}ͧ��&���:gw��θԙ�|�d��X�h�`v�R���P\b�}[��u�͟ueAқC���ݔ�Ӛ�֯c�$u}6���h-7�q��p�X�gq˾��ǙR���y�H���ڍ�/�%�Q�͛��Z��;V��ml��e`O��\����h���M+��W_,�$�t �h�R�I�8�D��s�ȹ#�EwI���l0�Q��{@����)8�Z�:��ɑ[����h"+%[����qpY9ӘJ?fffg'*R�:�0��V���l���.n��-^�]c��!��e侲0-Pݙ�ߘ�E�[�\�%�W]��z�wsFV�6Z	k*���������9��8#B9�Թ��uB*\�
=���^�S�����@����h����C�6�W2�w%xQ�Ҥ���6���l�D�pՄsnl]x�h��� NԘ$'ܐ�X���flҫ:.��BT��Ye�`�ȑ'��j�(��w��i�`39V; ��O��^�k�.}K;���2��r첷�)WT䪺IJ>����ъNen01��}ϸ+�u,�*��;�f,��t�Q��-�S��31�*h������P���=�f�\�mub/MA��s8��:��)���ׯZ���9�fV^$�VW*=��Oh�m��c�T���Vu;{|��,YW�����j=;.��}|l��E.�O�J���g+���=���~6"%$�%�&�IԘ�2u�#�f�pf�NX�i�zw }tr�����0���g��x@�Uӏ�Y�^=��}h�;}qA�Z��fAJm딛�]]��rU���+b��X^O�H�����B�tU�m#�𼛼(a1��ŤƗe[�$����d @K�	���V�@�};]�3�s�����]�Ẕ�]P�߹`���DX�e�%r��������z8mŵ6�7��JT�V[�Y�m���|�`�H������GV�B��۠V��v�I{e���1����x@K���"j��j�C���{i�����]xϷ6���4�Y����[�Nڬ	H���go���[��&w��z�����[�')��&,����!�U19���=��<�\�T�xm^�}��FU�X�*���N������o+&��Q\�V�<\�"ɂ�Q̱�_+�Hv3�b�ܡ�2=��\�I��sL}�Sa���������H�[Tv��v�^<dj��ˋOd�\�}�y7C�P�|Z�E��l���(�W޾��b���oj��틍h��@t�J�=z/fǎn۳V��Y�<ݬ9����� %�T3(�i�3j����'5�SX����ܩ�R��ė;Eʸ>�i��ho\V��dtv�����WLU������FX�J���&7�@7�{��7���3M��$�C�uh<G���i�c�V�=˩%r{C�ܼ�)�QH�n�¡jjVMo�}AwR�@�k^3���O����4�b�"�]��w/\yE�]ԋ�N9 ���d�7��ؔY�a=�9�<o2���n�w`������w;{J�m�85)�̺��20d���QH�5�*��G���RL��&��RFq�ue��Χ�jK��-�l�%�%���}�M]���/���kz@�᥮�f���\�S.�F>
���zm��瞍�=H�#II�}d�x�x�z�C��>��#���y����3�|O�sl|��$�:���|��q�k��z�>1�F��u��4������7X���z���}�{��>����_r�z�x���>��%'��&�Iy�|�ܼ�	�آ"����?��Ј��x�z�����	���}"�߫���=&��v�n��1�ƖHY�J��x�m7v�.�ƝU�YBY֪�&K�1�U�ɫ��LT�i($���U��wUۜ�okt���"�;�|/rDCqX{r����NS@?�<�����FgT�q�J5l
�zA�(���@��iDUiy�Zjм��{���X����̢I�r���i���b��̪�	�J���n���]��QN�@����$#^Qd��^8m#�YQP�����L�5&��w���p��x�T��V�uS�)E�5���u��L�:�}�nIG;�4:ѧ,�1�J�T��⌙�G$դ�L��u�W"5D���sd�Hs���6TU6;8l�!̊��_[��*6
d��)]���)�?"x�a��IK�9�3;~Z麃<e�4�h��:裛
�u7���`ɂ�=u`��RAu69j僊aO{6{��N��ZYv%�N�2����ǼԢ�����P-m��lv@u���N��l3�<5��[x�"�)d�d��*6���<j�7K\�b���$�[*���$�,ށ��3��J�e��u|c��wo]�*�\l8�m=��w~s`�ϵָ�&~W��.�`!��1��UsLS�Y�2F���Gp�f����Ҡ烞�.çAr���A�u=K�9f�XzD=��Ԭ��#$h�ĝĨXAf��wlV�}��i�D���2��-�>o���8M�$[����_��d��]�����S5�Vr`���Knr���)��gh�����s��ٙ����ǙL��Z-����\ݷE�\S�SLnwJ��z�	�l�Vj��*6VkC���T�f6&��rQ�̃A�b��E܃.��힩y���n���|�*�x����ޙ���{ۊ��dx�O��=��5Y����-���M\���]zs~@9Wc�;h�wd��}�Q\�*��ce�ݷr;} �*^Ҁ�;%!�F)�,"�����i*kY�1@'�BFo^���m�pD]&u�0B]��������Ǝ�"��%��zyc�a��[���gs��O,�X�cy�CP-G���&��H�@Î��k��ou,=��`�a�ɧ�ly̙m)b�Pm���PN[h���g	!Z��ln�j�+1��kGsc�gW8�!z�{L�kZ5�aÍ�K��0�o	;�S��gY}��,74Z�^P���+�[��������3�8�8��t��`y���kE�̴�jص(��׋^#�8�wJ��"E�32㢳Pt�iu֙yI��f�>ɡ��XiU�����ӭ1��y��A�4^ۡٔ��b姢��q�F^���J̣O5�&���+>�˥{2�Vty�g+J;���r�b0֜3���g#�VL%T
��w����໕l>�̝&g�iW�Yt��J��^`ܬ %\�Åi{Z֛���=V ���b��ԙ}5���SoNۢ+�i��WYx��*��7����KЫ���h�o������T�F,��E�.U�R�3l^��\n�戧8�ݥwс0^<�)�SFt��iff�o+,Uw1�j1�m�@���K��2�u���u+��8u����'T�Tڜ3:�-��<m�X�/rjP�Ko�n�ɀ�W��EG�R������ p0.��c��w�bh�Y��&�̛�[��<��N7>�):�@�L]���Wd�*2�8SN�2h>#��X��[(Z2KV��VS1{,a ���U��wW:P]:�N�U���\�ڶy�4d���식��N�4e��� ��'N�<��}M�d�����-HԧB��s˰GJ�������+���!�( �t7���fŢ�gd��ľ�[}B+]��S�T��w	 �t8l|�\�1���,���PB�ΗAtμM�x�J�֚˃x���`X�5S8x!���歈��}q�n��5yt���l�Ɩ�n�ݘ�����Pŧ�w��D���T�c)j�.٧wYxь��8����g�y.sz����<z
�Rp�ŧ�6����΢w������s5�cU1�X��2���9�UB��.��E�
Ǥ�&�4c�;����,v���L���Wz5h���$p̕�2Ixa�a����� T��*�AT.�X���멥2�J����;!���As��B�l��ζ�x�Ws��w�=!�:X�ĞLqvq�Q N�54���N�Jed�Me˜ʫ�Z���yn�+��*:i��9=�h�1��eꧡ��CO!�;���G�z�q��xh�s����a�b��³����w�*b��>��@�b�s!u]LP{�AםI�>�=QX�q�.���F_qڋ]���oB&e!��9��������w��g�8�e<dU�f�m�R�1S�	j�_qB|�Pn��p�{fd˵4(����2(v�k�Hc{�n��Y	���I�s^M����\�)�:�$��f�N����*K��L3{i��	�����Ym(C�c�Y�p�լ%�PW$��a���i�ծ=�u�A=u+��G�r�/�d�wpwi$�Zb��R6��/6�&�{Rv�9(	�ԩ�G��W�1ͤ.j�	�]7HV� �g��Z"`�56Q}����@fEW��.wۃ�p��WK0�e>_8�۳�(h,K��е�U�]��͙���jO���:��$�Ӛb뉭C0o�U��>k5L��W�����i��V��(�.�h���ƕl����7��ٍO�Sz��5�ы�M�{F���I�E��<{�v^��M�]�v	;"wNr����2to��]!ٕOz�7R�����+5�%	�{����}o��OI��������Mi"�|���2���m ��ʕp��B��j��z�-��æ=2�Q�W�u.Ȳ�[�� �tANN�噚C�Y@�od[m�m�؍=r.��{xm�/OD���2bX�!aV��%�t�Eߌ�d�:/v�Z�{V�jp�:�usl���h3�u��+����zu/�
�bUΉ��4�؝ھ�u�C�6���ͫ6�\�{�J'��� du��}M��{%�	l�
�;�f%�%܍���m����[]O��L嫰�/����4�tR�AtWn�I��1p2Cڱ�f�ݚ�U��ݽ�r�^Fq�k�Һ�(�SoY�z��p�헦�Xy�k�p�򁌠�*��Vb�A�f$�l��tbV�ҳ��,���G�9X�����E�4�깙��W��Ӕ�wf�M��E-�8�K����(��[�����2��;��H:��]k��	�[I� ��q�jU�ṍ��[/OYb�
�
� �۬nt�-��[���.+��b=)k{�AK쇍\��Y�lڬd�W�Bv��.��C���BZ"�Pw�z�Kk�U7�!��-#N�Z��n�񿙃\k��$������oS��R}�N��G�+�X��}�&��qV�f�繢��f:���F��m�i���oᩭX�W%�3�eh����sF:��N��!�w��J���T��i��ii�ڪ]j�j�2��d�*�OGةM?ZVԆ�і��K[Im�bv�v{�3�����e�]�t�ZCz�4������t)}
���x6��l��n�W��z��&R�sg�t6¾���W���n%�0N:u�ѵhKO��t�wF0�79�[�7�MN�����k�\,Nߜ{:���K[xt�`#��{R��`����,�'m��/[$� iU����Q5d?�r�^R���Q�"�����B�����Z��M١�:���{è��f��w&;gd`P˵Gar��`ԋL-?K��t{�7�B7/{A=���ˣ�⠐����LUKݒ�>}���,�w�}{J��Y����8ڵ��:p��y��m.�5 Μ��khp6��tL���r��4�2���:g&(�zfY��_^k��ܕ����%�4�����ح��9Q��ot9�LK��&�Ř	�l�jɲC�Ѯ����UA`�4��T/$α��ҌV��V|)a�ԇ��Db�ni�5h����]���԰�g~��W�K��lrq�V�C���ɝ.�����	W"�g<�-|���*G1��}aa���S�ۤ�AuwDM���U�q�v;�m����%v,.-�)w3����r�I:�cL��o�<b���cXƋ��:� Q,N�lܾ].ۧM͕�\��Z-�����̧zٕӕ��Zs�Cq��&�S����	]B
6��|^��t�I^t+���f��R=����zP*�E��Φ���a���5z7i�d�G�ܙ�kN�4���"�Z#9�E���Wl0d���r:�P<k�������1�U>_˙G�q�d��'M1wp!�S{�S�l�t�n�u�e���F���q�Y��x��'Y���1��I���J}�m3Fb5�;�dܗ۶���anV^��ͫ���r;���V��_)��F,���;�z61Υu��&�t�wdԊv*��-Rt�����9(s��nn�j�]AP�y�`���ϋ���6����j��J�����2�Q��̊�]*V�gu��
�%m��v����V���,q�Q�K"Qe��yP�HJ��bܒ��0�O%\���qn�9�p�Hҩ�Y��9�#��o��}��X�.b�B��~W#+�*�����s��ea�ƭ'l�U��P�*l��b#C��BS)�����q�6@y�(�����D�O|8<��c)�Y��;q܂�d����.gs|f�:��F�`�²v�q���.�D�xPsf9u�E�b���Kk�%�~�V���\�ܼĪ@VR�]k�]J7)���u
��]bw FX�8q��:f���Ֆp�oK-���5�Ɔ���l;��l�Z�#�F�O��ěy�p���]feX���XEZ���]ԕ*[W�����t�rf^�Ga8ns=�2#��Y�T?ܴpܷ�4��[����9��v�w���\�~�,���9eD����u�T�4 B��v�[ݩ�+7kq���^c+s`�q���y�Y#bw�Vcvm�z��^��W�Z[��6�>�ou�H�|=ؖa1�X���0��n�uA$ʥSk���й��dx9s�X�e�B^l���Q��ˡF�*q�������$�����`輰���0B����f;�;�b�x�F5;�w��nҘ6֙�Iζ�K3�	�hS�ּ��F�NW�^��̱��Bz�L��dǎ�IW+6С3U�njoZ��w#ݫ�;���r���Lf�q"�T�zrԗ��N��ⶌ<:�9��i�'��u��gFs��{�3)Z|���"�1�I.<�ϧq�΢R6n�I;j�;�6-��X{H>-��q���p
��Ӕo_gq.\E[�*# ܛ����ͣ(�M5��r�_F��X����LpA,EN�����۾ۛ[m�T�tK\���%�Y}����S�V��)�Rܶ/"��]J�	l �:1�P֝�t%�VS�����ۨ0��m�
���H��l-�q��(c��J �u3�q��l�NMӳ��UJ14u��{�&��2�]"��e������+0C�v�*�V�@� ޽�k��葜�� �pzG���h̗Yv��ǁ��N�a��}���,$�׬�ܹp_r�Zwe2MË��[��2����+�j���ӻK#a�֫8s������v��q�1|�B�_ʝ-��x1��Y�V�k�-wl�+Q�g1�&ijP}�Ò�"�Zr_ǝ��-8L��c׸jm� ���5Z枝��f��X��q
����6�g0�F�:�sr�`�O����)|��]����R��z��qr�ī[׵;�Y��v-^FJ�,��*>�S�mK�m�Adծ��D�Ī�4��9��qzj�eN¥�Z �h2�E&�\P�mr���oH����:���I�L&�[��GJD�i��W+��֩��S૩hYKK-��>����7�mC�W�%��}9�huv�����J��l$�-V�{0�u$Y������sn��2Ղ4-�K�j����!���i���]
&��beLLF��.8��65C*ehf����-G("���P	�*�ͮ��=Q}��h��+U�qCw3�l�y����s����_�oSZ���q�l=x�Ki'���_7zQ�tK�T���h)W�tF�McY�O/�ɬ57	3�1����l�\�a�B����.�V�-���.�10/����E7����&�+2'S'��!�Rۢp��;ʙt��7�l޸&aY�Egtɻ��U�D�B�g�U�0R�6n��S��gf8��yӯs�Z�1�ܠ�%V����}1�Wj��ogP�8f��l$s�J�6Aq�5
o�	t�Νu�E��n N�V�-��#�r�cT︁N�{�5�ƅjm�j�8'� d�XX�a��͏r�>�Y�&c<�~�; xk]pܕ&cҵ�A+%�m��ӆ'd�e�.�o�5	���q�wR'M��ALe8�)�]�+�h;y�R����� R"ըN���y�<�&`wӸ�ხh����BT�$�J�Frm̦x���v���5�k�k-v���[�r�r�}��{�)D��Pv>"�N���� ڶ�,���q�fG��#;t�=KY�oN�(E�&�ȪB�5qtiՎ�3�91�5e�\�-�UUϋ��y*^����n؝k������B��#�����dy��OPw�)^�p���Jt�s��AU|�f�y�ٖ����h��hZ�o���kU�yT�<M�� ffٝ����ɷg��f�����/�����?��?������}�ޟ���W������o���~t(y4��	)"��A���:�2���i�j(�fd0�v���;h]$�Є��e��p��!��B?�D���Y	��j��Q��������^'����G���p����^D�4��Ĺ�\����Z��i�ۖ� �K)�Ʀh���#m[ݰ>���O��hm����T�99��VM��7_uᤷm�+���D_q)�',��Xr��&
�u�3_<LQf<yC�Ihލל�ڙ��54iLC�`X�-��\��@��h�%����9]q�a<ƳYw��j=�kp�i�WPqb7}�yDݫk�L�jg5�;Ȍ�R�_��tT�_L���7%�է��Ŧ��dMt�ˉ���T�L������Pb�Gם��U�����3e)NRV���l-L"�GaӸu_U���i,H����C�ћ��$��a吆i���F��ud8�U�>�;��6�p�>�+�H2�]�;�yj���V�to9V@SY٪�\�Ö쮖���2�Pĺ��}�W=¹�Fʺ�@��\���xD�xT����hy��#�>&V#�njfɿ��JY�⚲#�n���0�����=VZ�������1�n:��Zmԭ��T�b�徽=䆬ʳecui�[�z D簝��r�%-Z��c��8f��H&�m�JE�/V��{��3]���G:�[�����
	v��yH�V��q%vm��BG�U�xG״t�V�V��"bb75�qٲ/^�X<�˾��|_�P��%7�2'H	)Á�D��qB�8�P��4Sa��%�(����D��5
���i7H����1��q$!.')��%%0)2"�Te�R`�Ŧ�e����a2�(F�!�`����ˈ�ą��`ƂF|�Ѵ�F`��M4�!6[��nas� i���B�A�QIQ4PMH�U-F�5����Ӏ��Ѧ��"��v�P�4�%4�CE�T�)KT:M1D�IUJR�ɦ�-�F�4R�J4��Q�: *�E;cAFڂ`�q�h���hi�i�����
�Z
�(j�6]HP�B�QQUA3l�(���"
"hH�(i(�J������h�J4$��`���Z� 
H����Zj�kNjD�"���@��hf" �D�8����h*%j�!�b�*�����"

*���e*!bԦ�"�*�)���IT�QEE1&�I^@�?�� ��0�H�$�.R*����E�[f%{q\�]om��m���)�w�t��ky9�o��2�����|)P[q�&�Zd��9ԭ�:��	1$ �� 
q�	A/��\���h�c0��pb�Hz�=f\]^Vu�U ��)IƩ����܊H���f��#s^�Ό����O�{�ft`�>w"7l�FF��k4�>��k��۱�x��4*t�4���[��ιOr��bF�ls�mϸHs���Gm�O�����AJ���{k)'�ۻ��l�=��Yo�*��
3�C����#o�\�T��y��0�M xz^�y�zǓ��A�ｙ��@�.�1�}���5�ƃ��;Q��sM�Z$�q��|zI#_���ճ�tb"/�<-�F�j���j�]�Wfm=춡�߀�$���T�8�l�m��/��(n6@a���{3K��b�D����V�U2_��}覕���}����?sP�.�҇W���L��8t�\����q�3�Cg�у�T���k�n����&@�mvH��O��3���^�s��7��NPve�}��cs�XO���v���PL6W#���"4[��snh�ֲ���t�
�}.ؖ*4�ղh�ƪ���v�'��,PK��g%���'l�u�6��=)��˗srJ��wǆ�v��]]�e��X��ړ��{��6�Ju�N�g~�D��e62s����n%Q���㦢5sҭԵ^��HיJ��G]��,�{��f]J��R}˞}~�����@
�liy9�`'��d�zpd��r W������¨���yRIN\�㸨�3�vX�L��tӋx�Ue��5��<�s��/s3Ջ^���.��{��/��>��0F��Z��-�jo{&<��ѳ��|��}F�{[����;4h��n����b[Onzr9�<��>�_��V)
�*z ��yb���� ύ����L��e����nM���@
=N9t흷WG)5G���Նy��x(;x�"k9B�]���?r̓��u?w��]϶���WB)�>>~�lA�w��ϓ���y����m�Xd�$�>^ש����8S�j6^�$E��soǠɪ ܊9�c�e�vI6=��{����ɳRt���Z~�y����>{{�Va7�3���Ԫ8�A:3��G��l'����1�,����;K��X��l�$���|j��,��Íy*[UY�mN��9|f�}9�m�� �像K�i{φh�=+�'�:�UK��U����/��������r�DO�ŵ1���r��V'�M��=^ϗC^���������!��g���xw���li~�I�����������27������7�	ݘ}�և/��۳÷�����)����Rg¼��Y���S'k~�K�h��U��2d���������Q�"��7��0�C���n\�O�%�9�\r���ȅ@��ó���x�ym�Plw�J=�,��j��[�7/lE��O�]���[}#���9q1�����5{��$! �6�;ܯ7|8I�ݴ��n���h�2S��9.*3�g���Q��27=����E�{�Q4��(d��j1'�v�G���Ow��K��.����9��ZE�:[>�U�lxZ5G�D��c�z�"GYMth��m�7�&pi%�os򺥻}�w��"�-v�%狀,R�>��r�+��tYX�j׮UH�E�U)d痴D��4֠�@�l:ܚw0�N��ٚfr�k�@֗o.C@�Z���wƻfR��簛�/ei`P&�U9R�;]�]DU��.G6~�v:S�7�Ǜ�K�yV�lE�=�5��o0��� :Nfh{�f��S/7������$`�'��;n��](��b��7�5PH6�3zksM�-�tۯ�-�szp��\��P�e/J��c�����~Y;-�g=ֻ�5�1$G�؈��I�x&��4 �ڽ�s��Ţ*;�3�H�������#/^7dM��Ƶ���]�Y�)��My����U���.�eשeW����y�rx������g2�V�8��7tMw#nz����fݼ��Ez��Jl�y�a�]<Z�0����X��q٠�x�=���=����Ǒ,���_yߜ2_�WI)�o�;���C�C�;\���yI��U7i��K�I�]'yS5���<���������y��߫�����ڞ�w��i3V�?�2^��^�ʭ�1��$d�'o� 䁹� v��em9y�Lf>���:�1�vXb�|�`�Oʻi�LV�o�P����d�)c݋+8���,x��/%wu0Me�oU&)Uhg�e��K�U//�R'��P���Asw ���)�
獧���<�U��Z��=�괱S��)d�ԡ�kp*"��ޮGX�L\����c�jmr���us�G�7 �U��^�V�+��+�e�1��g���h�e9}�w=��������)�pʑ�㵾+nb�*f*�3�VoC[�#� ��<����{�7�:uoX����O^�K�c��+�y9sD�����d�,�����->��z��w��6D�i�tu���P���z����mvf��e�c8_�����DԚqy��w��=�Eg��+p�US����,��4H�������7��V{I3�&wa�]�ݪ�S�շ���󾧻�E� m����H=Czw��1<ӒXQ۬�����/wr;-̊�q�"�8�h�o�v	4��s]M��RC��iI�>�V4I�1��ukY��^̶8[^���kg~�ݞ8ͣ�Y��d�N�h�y��mOOS�{�RC>_'��A��_���J���^e�����Qwk�i��v*ޤ�)��<8���a�(�_�(x`�ѩ��u3���u`6aI���}׎������Q.f���>ZxJ#�޺��v9y��Y�t���/4��K��W9p�\�Vd�Lӯ�+������}����w|Ot���8�l�0�s����IX4'�O�>�Z�g�T��O���b�T;�D�{�kƷd�Ǻ�O��$<������ۭ8�>��ޣ�t��L�W����/e������i�����`q�oM�A��2�@�7goC��rF�Q��OS�`MC�������FD�{c�ƒ�bڇ�s%[�j�4b鴍y�Ju>H�m�0����ÕW�~��L�_�)���j�WeN��*C0'ڤ��;%^�7��WG 3-�7�H�iX㼨�r�'�{���ʙ�S�}��N�=��R_8���Ļ���=W[�S����a;��oZ��2o.ƻL|GDc��&=3����2,�f���bL��1��:��!��̩�*i���{��KS�t׬��������������d���W�T}�Jh@;&v�ڇ+gN9���B��M�Jm�GXԹ�>Į6j�*w,�ދ[ܷ���=G��V򚞘�+c�	��V�ąo:���F�F���\��x�p�|9ѿ�hRX�}e�{.8m�͜����,Jx;;���@�����ճ�n=b*�G��-���`�)?|)a�&X�����]��Qsfu��}��=4��8[����=�r%��ڜXj	Zlש9\�{�W0��tMc���s:��
�c,���7ǲc��B�h��U����e6g������ɳC}h����4�r~�Oj������T���e��vy?w�H|�*�!�?QI�M����	��q{�<>�m�\� �ˆ�o�_l�����<��{=�ǽy�)T��ӊ�Rt���Y�9����n�G��l��o�vNӽ�=��>�x:�ߚX>qC�������,�����υ/C�4�5�����P��Uz+��uSY[Y1��A��������x�_'^.������^W��>e����MKf���ׄ.\�!��룛W.����1�w�P�̖��sh��xp�4sض�}�h�V	��U���͵��t�d:檀�}~�f��slOLx8��u�3�+9�ƷGEfD!��(�NK�(��^l��)��;�L�"�YU#{a[���N܆I�z%�1�{F�ԏz��6W&��J��>�H��n�]��.8���ˇ�Ps�}�����Ps��T3��߅vzbI4:oh߷^�y�����&�<�7b���)h�Q�~�;�>�#%�sψ�Tz�jv�dd��"��0h]laC|dW��QT��^����[쪌���I^�2]���ZF\f��FMYf5��z'x�$���f�;d��J�^�;t�������n�;ơ"���UF�����A�ޒj�IoW��5��Y�����^�6��
�����������"6ۄu��I5�x&��5�<j��o���wq"�N�csC�%�. }��ߤe����7d�a��7��~�T�{�B���wb~�'_��?���<<1��{�~��A�ɍ�ޑ�˛:��"ڳ$��#�\y��
<k�v�}���)���~f�[�̻ǝ��˳�K�.\���̐��9q��r9�Ե��s@f��]�.i���~��V_d��������b��U����>�b��|p���7]�<P
�Z�^V�(K�6o��H.��{��MiJ�wM��Sj����G]�)%V�v��t���twp��N�ңW�L������'�A=����]��e���{Uoh&ǈ�
�5�Ūn����;�~�>�= ���e�y����`�|Ɣ��j��w��qo�S�wK}B��>�9 N��s}�t�{�uQ��r�H��m�]V�q�CI1s{}Zs��|O�q��YQ&�1{�j��rƩ1�~1`M��i�Kp6�ܬ�̠�B�ߖX�W�R�^�{�ӝ�S�+�~)%a�g��|f~�i��+v^2��7��S�s�^�7Ke�N�v���35����'��Ăuɱ];� `�� �0�l�n��n��ol�Sg; ]�!��q4F���
�3�s;,�X�x/�����7뼭���|�A;~
d�\������}���#��}��y{׾�K��f�F�`��Dx���P����i&|(����og��W_^x��[�
s������#wh�l����ML���S]�ƥ�cNa�F�*�%�흌(�+k˥��{��(m�N�W�/.�Xc#��X�Z���؝l:�_,�����*�ts%'���E2�A�=��=u9�gc��T��}��ͩ�SOL�:��Dm��;>m ��+�0�S2Uں|�ݾ	�x��g$�̷궱�q"߁�+G��2�Neh��#I�#N�zc=ZCD7�&`�i��[tx�>ʕ�C�g%3����/U�g�LF�yH2�{i��{��||�f�}B1 D^,]�����(��&���f�b��0���/2Yخ��	����#�>ӹ��J�Q�������"���B���'CQN�=2{������u~(���L�<���N7��g$C�Q,t��i�NφL�l�0rF���q��5<��%�����,�t����+oc��5����"�e���4:	�8����5�dJ�;sy���Ï���T[P�&Ju/*�zX]:��4�j3+�3`͜��LvC�m���{y��wDv
�ݮ؇>����=�>�W������>>>>>>�w���������7��1{�sQ�"2�\Na���������c8�����ue�l�Ե�ٛ�}�E���1��z#�˵��]i��v��V�g2H,�� �'���NȾԀ;�Q���/b�,f�ep���-�,�C4���z��)n�g\Ɍ�������� �ir�J�+(�Zĥ]b�q�G3
�9�J4{�÷t��%�F&���%�E�s�^ p ��oo���ն8:���kF��t"����6�V�29Jnb��mC_l��_a�G�l6��r�p�x��zdz+�#rs)-V3�U�W2�S�0��3E<}&�����Ņ��*\���(�w����{�M9Z
���If�N�Y�g;��Wʌ����}������''�x�;w!�Eo	�����Y��x �H�+���H������V֌P�Ǳ�G��ھz�V�q�dJsR�ԩ�/xQ���H_ʥ��SL����G��5Ƒ�w���[[BJ8�²�E�$(�5F�k�8�1� ���+m^�AU����А5(���4m�&��X ��f��$xġ��_m�y\e�rp��e�n=#���f]î�,�=ӏEIГ����ZT�=�����q�=qo)p�m���:Ywr�I�{C�n���kX��r���p�ɏ��n�]��,w�ea3�
: ͌V��O�`�w.��9s�{F�ȣGT�
r�l�6�.��j�ڳ�
��s���؝Mb�ͅ��Y��V���s㙲վ~����]��wC�ㄧ�>�w|6^]�3�,��[���O����G��~�������wU:����heє����������+b��dt��j���eA2�b���Cx+X�_-�.-ɌT�j���;�o:r��q�;1">��j鵈VԸFk�S�$;���	�r��Zi�XHQKz6��ދ ��#x�&�<ӶK�a]ù��'S�+i�dg,��QU��YC�}�`d�����M':�=�=V��X;�./���]jvs�u��[�+��3wl��	h��vƍ�Q�(>���+
�l+ivvs��kp�-b��E�A\W�L���Gu�lX����7��T��r���̀κlԝī�m��$�6w��S��|�j('.�WZ,¥��A�*�2�Z�E��w���&̒�#U��vr�2�/I�`��U���<Ԭp��{�=;��0jt��,s�N�hQ�ʴ$��h��L;M���XfkF����_V:�0�[Fy��Ƈ�}����Y����yzE^�M�Y��4�=W�f�<8s�J��{�b>2�����TS�g��s{����EG���&pݏ,p��|�ڍ��`丛#u�	|�9N8��6��7nM����k�s�&V�K�ɤ
�h�O����6r�V;����5�s'���j}n�&�7�*>DCZ$;2�%@�v2���s'����]\�N~�����ȄI ��i�����b(M�
Z
�e�&J���J��h��(hh������
J
OR�)(������bt�C�P�4�--�%5M+V�)��
�Z��b��@Ru �^JQK�!E1<�CMU4SM-r-�$�BbK�4����1�6�T][d8W%�3N�ՙ����15�N'B�[�t<�41kF�u�UOQ�#D����\�*�m���A�J1:�֍6]:���jm�TA@m�nZZ Ƨm���I��`��%:
[�&]r�3�PX3���Z�1A��3���1�e��fjNUQhִ���e�tr���T�rW8�l=\���0RbE60R;E��i-�
5�֢X���رIl��PU�͇��>$��}ӽ�?f�\�Y�l��bOC��S�`�۹.=��`�f])dl�+� L��r%y��bt�}x�[D��|}"���{<71dQnMkl�����g:XM27k��F��8#}ǩ�|_E��b*�᝽�Lv�ʩ���΃�,���r�l�О�ǵ�=C�F�f����s~d7�ӿ���i��������� ��w��u��G��2��l�����FFS���s�ܙ�RR͇!(S�@�{c$�xL&_2�i䑹�h:���@�}[E�%�E��𠪱�V'b�=�Jlomn
��S�5��쬏�]Fh��R�aK�1YR~Ykc���O�8E�Ǽ�`!��H�T��<cc�l�V���ֲ�B
*%�{�Fi�#)��6���`s�:y�0���'��>�bO��.���: �[CSHBNJ�?D�Iؼ'Et�eI*L���j|��U���]5�1C;*���E���L�a��L �Gd�>�ކ��)? b)9\�%p[\Ø��p+yy����yG.lT�.���P#[�=`��?-��pnO5'��a�:l�&-8�����N�2�����+�.��B���	�?K�����r9��� �\�ՓM�;UsYt^�7�y�<�������u1��g1���Y��J��֧l0qc����L@G�5_w����RU��δ���s1�6DgL���=���h]��Vπb��ku�R�$�l�d�-���.�#��R_58��P���'EC��E���n5�yQӼ����=}��P�x��݈k��M�G�EڷW���H�xQ��X�˹�C�~92'�7��L}��4ݏ��l��vŝ�~٧�{��<%{�3n�/����Dc�A\��ුh��	����t7'&�J~�TxL��C�pc���,���LcYc��Vؓ�^/��:�;wA���TG�'�f~C�z<�B/V�sgn���������A������X!Š��[��m ��p�i�0�2}�+���Y���>���8���k%c��s��"4���C���0w�I��u:�]`��
��E<ƅ;��Uؼ-Z�>��s����R?0;.���܍�	sձiB2�3K@�m�v�gְߕR��[$�?��~f(?x����n��`����Z��y��O��r�Jb�VJI�|ض[�,��T��!��˚�T@�ډl/>�g.�Ƚ�v��i/V��L �Z��OB�	eA#X�_��^��8fA8��B�K#�,�f�Ӷ$�a}����y.��g�5����s1���4)X�E�5+�m�tޟ7�=ض�m�E�эd���xGw��+2�7��e�ןGJ!P+�׫2��DJΛ����5����7�y�#d����|��=6�A�Bn�n�8��D�1�T%m�e�r��Gǅ[:�7W9��m���Z���؋Z���ȋ�u��sdc�On�w=�4� ���+*ߨ�:�?v�d�C�P�M�w_(P>�?�?��25���i����%�1t�]�N�%�61g�R�ޚ�qa�yS����v���۲i���h4N7�HB �vH8v!��˷�Θiԩ2�0����F������C<ͻ�\.P�t�PV#������5�T�B9��ꀘs�8�]fa�����f�w��X�W?J�zA)�_��>c�������+�\@\���fy]؆�|�����]�O>��i��""s_L�ٔ*�5�*�rW<��E�Ґ	�~��"ɤL�k|����?V�Ύ�p�b��1B3�Ӷ�5Ӡ:��Վ��j�H\]���Y�̨��a ��}j�=�x��`�>�P�+!��ٺ�/��(0|l`'�&U�#�k�д�8�cҹ������'X���ًB����CC�(��l��!�� (;�4?��'Mb�sCjY���Ú�Ԩe�k�wh����b̵E��2� �δ9��-le�S�PgY�"]�p-�D&�޶�R̓���������ܟ���9E��fqz��[��.ݏ^Jf�z {����j�~Aև���3�/�0���7�ś�X)�MD6^U)�4�m5.x��kl;s�6��Y�`�J����������nJ|���|�Q�Ef�9U b�n��J+%��3�[y�&5���񎝭�楽��FA�+�ξ�/�8P;m}|9�pJ��NEn�vn�ڋ�y�q�W|9�}�{�}���h�.��>&
�C��ЏL4�l���3��(=��3=�e���dT��EpwN/��U�k��dfA!���\��O�2�5t�ê�vڽ3��|՗�(��s� s��q>���{��cV�L5�jR���Z��Q�Czq�L�k�kֺp�w�di!��L>%�!66~g`�s�����ږ���D���&UhФ�S�7���)b��5ם��u��/�� b�|�I���!#��CO��W��������s+�i��y�B�א��[Ҙ��b6s��ո�!��y:A�0O _7���f�D�O;�<����ח���u��K"�<S �%I�ؾqA��׵��	�b�M�ީxnv�U����T���%W�R�{"����t��7E2������-N��50
&N���}G��"prf� ����Oa�F��P�⮗�f-?5���]��	p�j/�Wے�l�Eh�v�'�[>RPa���M0Dk���d�0-@��d�2�Gr�g��Ԁ?���y�Q�yv|?k�Ul<��H[ ,_P�7�~OvR��io+c��.�akܬ��~�`R��#�o>O+�����~�;ǁ�V��'d�rK��@:�ܠ�N�5�mf���\˙�[�K7�!�o%���O��s]x��:��:+���{�ݑ�\B���w�M*As?�~��j혖��TZ�aJ�a\zW8VDPKV�������=����/-�e3Et[�(����X�C\����[�6ɽ9Kbs͆�5F�e,�y�1L�i��)����3��;p�tņv26<���h�^z�f����Fs�Wae_�����M/{���_�1�IC�@8Kϰ� �-���D��A�xO3mFp�g�1oj.�1�f�	.�vN�K޺=���cx;N��Šǥ� �u��O3pK���������~֜��Ȯ4�9�����j��I���twH摻�����,��R]÷���Z���Q���u�V͹�ה�z�m��x��֖�ɓLde9������͵{RTͶ� �7���m�'����IhŌ5��p/�6�U��?WAH��|,�a~�.=<(*�`���'bϖ�f�5��x��5e��M�Y�d�J~��
<��I�e�I���08E����ā����Uw���F��e򖪴�k�<�9���K$���+�&���|njgJ),��a�|~�f�zUw��յ3~�nH:�r���9��E�Ԓz�
yeH&���HRd8�na��B�a׋1�-�Yc��o���ʃ�Z+�o٭�g�{v��N�\�X/��Y'�>��u1˧�;e��3��n*�iE����8ї7�S�bn��/=�o1�{������< �{U��ڭb}9nͿLs'��vQv/�;�� �E2��&��GG�����y$���`�`n�0eN��n��//!�ͭ"�n���C�Y�&OuI��b)9\�%p[\Ø[�����}��\�;�R�t�<�!�[C�zM����;��EΨ����/^ŧ���n3Xm�I
��4�!V��ۯ!@#4�|_���XE�2�F����bYs��ɦ��:���C`�p�����hf\;���=��>�C�ćO��E���B�a����}����
�M�Q�h�B��w��TvP-+�ɬk��Rrִ���U��B��`2�-ݛga�����G��`�}N_�Y:'޸;C"��馅�����,s����ۓ�E����;�s���ܪ�
�Ռ�kv�1(е�B`��mP鯞��2}�2�J.9���¸��LW5�X��Wl�?F~������6�.�@���L�,;(����|"ac�ڑ����� �D�j��"�uE�˂L�-½ۺ������|?U��R��}�D��A����I�z���8;��3,�47���,��n��P�������;㌅�]�7x]$�3O(�QS90�4����{�VE�s_�`#*��u7�S�
{��r����ٺ{*|x�����zC�AY˻.5,�N�I�(Ӱ��g�s)ws0�����E���%5�K��vL�fֵ��՘�W���>���=_W�U8�)�d��`�̓;ei�m��˰�TC�Q�7&]���6����;]�`0&P�`��d_=Us��������r���Tٙ��Ӫd�
�X�Pd�k%���>l[ 7���Ϲ��[21�C��p�����ͩÁ�/�Y{`�NHJ��V5i��at�-@�T���3ю�Ơ2������N�:�ૉghn����Z%xbB'�e	�3^� kp5�x�s2�:�F�+�E���AvN0Z;6����+{���l�a���\s<���R�t&v��v�=����~~��=���W�o&�-sCt�����V'%p��r����9Шt�z����C&�v�۝��J�&�^aZ���52������5Ǘ��V���_�ˀ�t��-Ơ�cH�!?W���Y7���J���շQK���d9T�z���]`c�V����@r���D5�!�R>����eᄬ��zf��a"�7��'$IGi0�����"�JKva��<;�͸�n[�Ұ=�s3�*5����p:�>S#�����|k(Y���.�%Qo
gO2�
�XI{���9�Á�oQSh(f]Oi�zAՒ;�)G�'>����?�`��(�S!��[�C�90��i�z����ml�=r�!�f�]��2t���ӂ� ��ݮ�V塤�*���avj�� bY���x�!��e.&����<@��.�t#x�h7����[�/c���*���<<���p���K��-s���	��X�R9��i�V�V����y\�⠗���9�ia<8�����Z:�� 9����;=!��it[L�涥�m{��j:�x�k\������~�jm�.\�|��c-���\�s�2%߁p��x@x���R̓��noI�{޻Xr��D�=�:y�0@%��9K�ǡ�f	��|�@tg/��:�B{o��t6C;u�أw�n��^���a9��<PސHz	@A����H[ ��m�Ϡ;^[�D�5d�Uj�GV.����Q{%=�/Nk�g�ts>̅��vA�,��r5��t�P�V݇_$�O�%����V΂���w�%���t�^�veB�P���p��Iݩk�����B9_S�b��ʽ�S<!	��	����v�βW;Rū��J`2��!2ok�U�-�PE�'�4�h�CK�'�(_�y�qU�eO��`����?!<�'*0����>�S�Nn�ٚI������5����
[�<JsiI`��^q���j��xOV��C�d��0L!@�����^�H�+`w�/��]��Q�JN�s�-T��Sܓ�tfc�&c������E���՛Y�D"��3�[�p[V%k޵|�]޹X��mj��x�Q�֛�K�jJ�*-v;.E�ʬ�r�*�}���܏,��WɓG�ۍm=� ���z���q�N�M�b,}�W����e�bY'Y�ʀIRaA�/�P{���ᯭ3��=gZz�s�;��|�3�]:��˱�B��FGdQt��*�]g��
eAoT7P A�-N�<� 1�Z��)��1�~�~{<z���P�!p͌�9n�1����:҇@⮗�f-?5����ћ�����9d0�f�o���+{� �})�p��!~:c�zz����L�x�C[8S�t$iKׇdw:����rVx5�،J�������kg�T��0������/��^ښm]2Z�pR�[�u�?A��/�f~Rv���Q��^��4�w,�]����P9��y �����;����t<�R��G�m����O��\��������y����Y�z�p�8��p2&�K5ViZݲ�}�_��О��P��-��ұ����-��󯧴;3�u�>�s���C���X����W���<hZ�y%Ĉ� Y{Q��`&�����>ނC�ghy�u�}�T�z�W�T���?_o�;֪�q,�K(d&�{d������H���f����K( ��o0��6�+=�+2��A�Ø8'�]�h+����,G�xK�
�л&0�vJݐn�~�㙧�8���2�ln`������qC<�����<���up\�W�g룣��DUzIr=t���V��֘19�$���Y�۩���߄ompn~۾خ�������\z;�R��p�U����xi��a�CR
H�a���*�zy�ݓ6�9%L��b͹��_=lKحيX:f�R3�5���ͼ�_�\+󮿩��(�
Q��a�uJUX�'�뺢�:s6�6?-�#��м�4%6ZR� ���4���gX{��oV�^��;�
H"X[xϡ���8�S���Y������f����I�f�_�Mw����{`<�{w*�E,��e�ü��7>��Z%/٭Ls"�H"Gf�`�a۞��^ɹyt�d����vO0Ssʣ�E�����
= �5�=�=2Ͱ��$`��L8��4��E'+9�����Ͷ�ʫ�DJ\�9���p��2z7�#ϲ@��C��d����������sۼ%]�t�B�y�-z��or`�'�Ԍ�	���E�2���D����������c����^t[L����|��yԶ.�O�cr_u~6�����ՅC��:�����w��K�b,�ؒ6:-M���ok�R)��6�V{�Rr��&ޭ\�T�f�m^�{�����_/O���|>�ߏ�����w�����{}>>>�_��5UO:�6Ol=�d�+IBe��mL��ǽV��} ٕE�B9�|��],5:�an����_d-���NK
��R���2K��KY��0��6�'�WzA�%q����2�>�D�]���g�a���Z����t��.����53���9�G ��<%r=����Mb옒�VF� ��9���> �+mX��	7FGˮ]�tʥ��
�8�[%>�e֭�eM��_&��0B͝Cv��'{%K�O
�p�x��B�٩b��6�iN�Woe�'Q�_]�<�]����8A0��h@�[�V�i����}��F�-�m�4�]�P��;�Ӈx2����׺ì,Rͮujnv9n��w�Z<ɩ����y�7��ߏ�!7���q�2zʙ��3M��ɺL#�U�0iȵn��{��W�h(mS�߳A��v�\�ק4tǚk�3�5N��K�A�L�I���t\H�NES*�}��.��� q-���RށEp��
���\����T�Ԗ��e��mH����`�ۙ+��;�p
sr�(͒���O���$,p�T0\��W��oPY}9����g�S��AS��Ѻ/'<������V��a\+Mʙ���2��ut����j(l���C{GQQ����[�S��xg�HEJ�9�n`�C���l�|r�ȶ�F�o�j��(ݲ�nVgIh �t�os:�t��u��I
���V�Ūh��Ӕ_�Ys�k)��;��;&�YS�c�͈�/zB3)��F��1&��8HU�f��8r�u���E���o漆q� +��u�^�>�����z_��V��!sr�4��W	��duҏ7�}x��f*�8Ѝ�*;yi��m=ΓF��v;�{��q��$�|2}6�]qn���T��P)� ��v'Se#Q��V�f���cw�����ݱ�����H�Z8�Z��f��Y7�"C�]�S�S�j��EL'xe�N�5%g5v{�M�e^c�Fp�{�9�!YL�΁\2�B��Y�aK4ܶ�@5n�V�f\W�	חn)0qZ���{��	�%c����Sq��2]���6�u�u�ɲ��ɴ�ܝ.+"��V�N��\Qz>�-�x<kә�����Z1��c�o*�k�����eyŭ8%���׽x+��Mkܫ���m�u����/s�u*#J2�x������|�ΣQvoF
�W,�p���BZ����x-��y#%vJ�;)�4�[�Ra�3kL{c''L^k�g��7�Y��+�#g��]/�E�
��GIm��gt㭥�H���YϦ�)Lޔ�nS<���.^9���.���׉<�y�5�W�9�J��2p�٦�}°�E=�C�^n�{\ ���.5���)3*�i�7�9xȉ�L��2Ku���b\�{�l�ĸ�EEX�l�*d��g�˱�����\0 �R�^�}�ȶ�ư���Z�r�G�-.��7�r�ZPE�g��v�@���9��>�@����th
R�l�1��l�4�M���i�2W1�A���`�"�	�M͹��$�n��R4!4rxV��m�@ru6��:-�{�Q�[m�\�����SW2���u�U6����"��l�S��ꭓE�S�r�ƓE�q+kEr1AHD�AUE�T�Q��AALI���(
J�x�GX��%�W
�j�:��6zڢ&Jyk��(�(/x��UW0bj*(j��"�����Zi���F �����E1<��QE��D�T�MRE��sj":�94E�N��lƪ��$�RDA<��-�v�:�OS�Z(<O �QEUGW ��J���E=cu����H�����)����9� ((5�
(h�
&����;׮��nU@�B0�Q���{_�qK���ۻ5�7FsZ$�g���*�v+w])#��\9��ڱcz\C�ة��.Ƭ�vK�zL��{�E�AT
5m��I�(��D��pJ�S�|��Ԁ!@��
���sz��~:+���o?Tn@�������j}ǯuC'��j�jéL8�V�ǧհ^y���`|f���~q�}����������9�Bd��-��\N���V�JN	9�a\Z�^y�ۆq.�>��I���X�-MA�"��<x���0(-&jV��ͫvCk��hEx���ޥI�4'�ne��9j����3w�Ŧӷ7����"��..���l���~2�\sH���_T�m����莁	��(���[���q�X���Hi\���PJq�4;��0Z��r��������H�����:��ƼN2B�ͺ�U�&׳W�j$Q�A�QY(5 ��g͋dދqL���߆�Y�mlC�A�9��vs�]���^�P��nr+S����	�Z�	eI�z1��� ʋ�-�"�5uw����ܫ��ב��2C�^��0LN�H�:ɨF@�
Ѓ,~/)ծ�%*�
`7�Ν�^�����u�vN�p�����\9��g�[Р�5��N�7%ۄ�Jnj~��=��N��7�qUI��8t�Gv�ErT�iqw�la#�-��0��� �M(��ƿ�E�x�lύ}���X��ᔤY1�3���^V�Ӷ_u���:S9���Pa�jQpO����1^խu�dA[3��wul�5�u6a��0{�>�,���ݡ��T/%���\���X������61�%�԰eG��R��
��z=|�ׯ^����u�� ���@)���#�/T�V�n���"��D�6"=ͅ��-ᄍ�B1�����nZ�Q��3n\Z�xtd�(a5ra'�1L����o<���������[P8Z�e�v�d�����9�MƻgV�t%�]P�U-J<v�
�rW<��I��RX��5<;�������?F]�L��q��t��Z���$����Vh�,dY�:��RX���U��a>/vYF�'���aZֵ��ˇB_��Xnn���p�1��#�hv���D�������$���ts�vL�U���C�U�Uv'Z�XFs^��`��ft69�@|NkjY���Ú��@��&&�Ncy;��j��s��r�`'+�KsQ���*���^��$�0������]����QKNµ�����Z�cҙ�r5�(��4@����#>Ш�9�+�KJ���&F�����x9�&v6#c�{����d��#���3�xހx:.d�N�U�5��;�j).��0ݣP��Ĉ̔^�5�m{��1�(������B�F��댷M��yǧ���\�u�K7�Lq:(z�~�����V	�\�u��Y/�e����$�u�g� �{��a�4ǧN ��8���0+�@'��٬m���A�j[�#S���7 �c���bVE6�2]Z.rPVе���R�8���4볇;���}� }������f o������s���}�0Um/
UR���Ԗ�ck�W���HZ�veAfP���A�5�5}-��s�^ �ɄAq�]_k��^8pO�-�����2W�ږ�n"X�ku��W�My�#1]��w�N�����p%�(������fy	�eǞ������.���T���ηw>�s3�-����2�&�!^~��ǡ���O�N�Sbt��	��M�1O�����m�-���S��I�1,��tղĖ���C΂��q�n�~�f������Q|���� "1�/B]S��%Wey�E��Qu�� �U�P��0i�:O��m9��b��?E��3�]y��7�`2̚a�C&�p[��vl�(qG��1i��I��W0���KM�ת�3���ں�z�K�<���G�0t������z��a��2�r+B*��%v�94݈-{l�	�T_)t7����Ӈ��#�F�70e�ѭڸL��G5f+�%k_AG�T�vW=����{
����9��@A\9�����ψ�ˉ��k^��,]�K���J�Zx�4qL}0>熍4�)ʟ0��Zg������#�]�i��ml9��;\��Z�Y�L�T]�]�D��n�n��]kT �-Q�w�;���H8f��Q�߹rX���xB��-BH���Ԝk��c�������2[���I�i�vm��T�|m<�������3�^;r��F,3��`3?�6Ld*��uk�m��<��-|𞇷��A�k��K���=$?qנ��I�ū�b���jS�ƒ��`��R��ָ�f���f�D�c�6�؍�$;��Ť<z���^�x/n?��\�O�ꈨsF%��->C �!�z��ǳ��9�p�4u�aۼ�i\�������m
��-Shh��R�_�r���O�QN����k<�vI_Ԙ?�~����p{�*w��ѽ\�Y�%(_�_�N�L������cռ*���h����/�������)7��{<+-��&az��zIBSe�A���/)�~��:��z�]W��l<� �B�j�x�"�ss�A�� �=ƽ���\���A8��%�r�1,�t������t������f=�|u���u��bS�e	�`g��A�y۞��9�N�@�\J�[:���TukZ��ٕ,����8����|!'��mQ����v
{$É�I>Iʯ@���'^��0�j�m�e����\(�dԻ�G�G��v��V�V��@�`m���	e���{�����el�z|�Veuz�Ʒ�.U��l�����tk����9���"����ʫ�w����E6�9�i��ѧ�b��el�gU�}�� <<��x 7�>��}���1�L��7���	�*(���B��f�0M^���������!�m�c�l�O5:��ۈ��۰�+��t4=��n0�.��NVR	u��w ��=�.�G���ׇ!�r/�=
g ꉕ��S�2i�F���vQy��5��%Λ�h1.� lc;l�	������N����_z����7j��L	e�ɬk��I�-0i諟A��l�l[�6�i:h�Xj��v��ýqQ�c1Їb�=���>��T-Xu%�PcYc��������j�c=���\ʫs/�q��z�뵌�g�
����L�D>���d��d?�\r	��
�@;x����L��PHξ���ůÕ��)��/��q���Pk%}��N�x؛�|.�z��p�q�Owz7����*]��(0�A�^��x4ȗxy�6�~k0���m�3����h���7��o�[��.�%S4PJt�P*q�j�&a�[�Z~h���dS�`0%�[FE�-~̪T�1�x5�����W>�c�+�(H88�2nd�ԗx�4�,oV���Ϝ��|��OU�L!��䳹r�����_<�f�9�/����z7a'"�D�n?(��\���\�*ݬ1�B�:D�poz��t�'�������f8��Ã���~w3%v��Z.���w:������^gY�IĀ!��U�9�Y��7�;��ꪯ���%"-*4-B�߯=�{��(�}��G'�|Ǧr4؜�ƭPA�mOA9�K*(�g� v������dp��# ��*a�(�0(6"y�P���mQ���!��A�=�N�b4)T��VNj/^y����)��VÚ���x�\:�q�����f�t���v�#�SsW��2O�Y��G=Pu�Q�k �s�dS���QN.�t�Ǧ�����F4äL9��r�����)�VXמ)�r�MQ6ݾ�P�gd�@2���h�.�}8^���n8��i�'�+���v��hVD�u��8�{*Rz�Ⱥ�Y��6�Ms�w�~�E@|l�V��J�D�uY��"� e�>�%�9�uo�i0�%s�Q˔��),hv�������t�ͺ*/n]H��7���w�`��<�ր���xuEs����1'\Y�<��<ʬu��Q9�T��>y�*�������[ۇ�H}e,[�} �c��w�еaB�6��[��}��x6Z"�Z��u3�v�/�b�?�bi���]0B��%}ᯌ�R̶�h��>a�;.�61���-{�q��9RS�W�ebX�D�S���A/�%��4/:L���RR��Ҷuƈa�Y����5�� ���W�K���5+��̈H+8�1M����뗆����N'g`n)/E��侦�����{�Vp���?�� �!B�*SJ��-(������s�)�F A؝�C��x����0���d���z��Y�"cq�oVs>��A���m��w�)3M�EK2[yE��$�q�co���4�w��)V���+�j�!��=?pIcʙ��,�oshG�zu�
���29��f3"�xހH~J(��I>�8ȼ[�"i�����z�#3ecN���A�=㌌�I�j/���kNd� ��VHB��~f�,Z��l�b]��f+��B�D?Ƀ�xS�~6���m`|��cS�Ak�A�[�Xq�
3,7�9��8�{�I���w8zӌu���΋�g�!64��L�������Է3U��0����lb�����-��ƂeX�
O내{���*���R���<���	಄�H\��'�;�#\\���Z�K�o,�Lx�N�*�	�T.�1�q�=�;���.`�5�*8_VX}B`pO"˴ v�锝g�ĲN��)� ���_8���O�9�Q����t�J5}3��6�DB`��n�Ƒ*��F��a�as�9�P[�����8��U��w�n�����bF�ݹ�ׇN�Z���-t��wfH�?�8��i<��3ӣ]u�3v��e�}�����>��u1���$�y@{�,��+�3����dDo�U��3zM��bݚBډyi�;�����uNř�.�2�J*Y�߿W�W���R�T�
T))Q�@��
R!�;��ǟ_�����>+���;�3�ˇ�Bݛ��-�&n�2$�;JU��^�ŧ���w��Y]j��O[�.ַ!�;�0�}�d0�t�Y�>�f��urg�9B���1]����ӡ�����S�%�U�����T�n0���:�����mJ:�8���ڞ�[�����Tԝ��Z�R�XP�]+��PKܺ���w,�]��GO�p8t�#��MY�n��T֎���i��L3rz�m��T�ߓ�S�3���;;r�k�,3���:�k�R�nե�F �?S�yO��;��`3n�J/�Ǥ���:���:"صnqLX��\�=���Nup}�a����;�h|a����"T�}��t��c;���.%�zZy��&�m`��a��v�����
V-}7Mn&U�~0����=�OS�x�s��4��4��+rt�ow}��O(����T�p��y6�=9<(0�u)p�~���X��F���̆���zլѯ']�3QӘAqu
Y*��l �ڜ`�������i�wH�x��,:/~a��B��V)�YJq�y��m��k�+9��*2�ef�WZ��*u��Y���æ�Q�a�}����Πv��g/z�$+gi}�lnl9������u̞��۷�z�e�c96�;�,+ՃTot�*J ���"�ai�V�bmofm�3�R!@�R�2P ���pj5�?e����p�4�!{l|6�X%��<���=�eMV��{��8Fc�M<�o����WA�t�q;��<xV�CxaK���Er�>ǵ���N+��i�|�f�\�I��F��A���§�kSc�yt�H�#�K�e	�I`�(H#�>���> �%:��E2�����
�Y;bc�-�����;k���~D����'(G����"��0�{��O�
ޛ#��$>�ƻn���6\��WR���s�e�>G�d0�`��!�n�pm�nO5ùI��2JR��[��n�;y�6��r^��A��]rx��z���k��C�.8�;�t��Q�S]O��1�{��nC�W5�yW˯%�I��t���^�ha~l�n�"MOw���8-�^�ltvdJs�Ԋc@5�w�)9ki�oJ��j��5�ݛQ��P��,սF���}L��
��y�d��n}�2)s�L:��5�=���l�g�n�h�)����w+���b ����֜�-�2�J.9'3L�<��ٮ���j�I����5�;a\)�t�p��c5H�m�۷��t�:Ҍ�L���yZQ��h���p$�»3�û�uF��(S���c��Fn�#5�v���W�Z�[����*?[z�S����CW�&7��G���]8�e%z������_:�ϹC�
B�@���*B�=�������<}}_=߆��7�q�.�h+	ɔ�>(�����X���k%�!��'.�4Z��y�������
��j���Lq �/\�o`C��C@�q�"&uW}.�]�5Ϻ�N��R�S�`5c��}�����%ځS��R&a��Z���o`K��0'e�31Õ1YM�*V�U�����q���z��ն7b��P92jb�0d�c>��2��l����ܚy���ĺ;#4۹�ֈ)����L*&�#s�X��PB}ka�-@�d�#V�5���ڹ�����Ϗ�b�~j��r��fpB�s�)�C�;X]:ɨFB��X�(���[mZ�B)��f��W���SP]��^ꋇUq��$AoB�,��87"<'d�x�uy��A�63^���Vᆞu���F����1��GM0�ȶ�C���`D�;$d9����5I2��ה͙���|������{��`$���,c1\�%>�"h��/@;�0������k|z�13xs�)�X-�	���E�%��CvL���6Ⱥ�1��>y�m��f�~}�O��������x��>�w�����{�ޏ_���v�f���k� �Z1V�R�%��õ1U.�B榘�>&v-���ɮ}7C/u���P�Y-_q�;���4�]ZP[Xf(:ȁ5�ǉ}9ʋ��lH/ʹJ�.t�\.�D�:�e��E,�x�JHӈ0�Wy��#�tX8]����d��h*�<%�`�@��G������W�A	���5ϱ�h�r�jnN�q�w��἞�r�zt���nHM�(�R0۔�1�+�nJ\�&��V��F0mف����0��úH�ʝ=���+#�Z�X�YL��4����U1,���)��ss!��U�y�3��Dܼ����P��|ia�59��FT��E%�g5q�F�D.�4'��u��K��x\Y�B�r҅�\�:��b�;��`�+fG����;H�W$�\ %��:����_]t��p��}jub��%�d/��Z-�"D�Λ���:�g���X�v���±���]��#C�A�j�z��y<��xbˮ;��U���l�ٲ�r�lmޛ7@�H�^kRCq:L+p��*=�l��eG�0)�֢�=�w2u�#]Cη�$0f�����E"*mX�6�t1����N\�teIYȞb�3�;�ɕ� ���Y�Z*��H~����8��/��S_��F�^��������T��X'e<0�(��$��c�v�W)q��M16
��F��M�%�v�Y�&��6�8�K �W��yy�FG�Ń����#��2a=�������S�e������{b��_PS��a�פ��^U= �2�1ں����-Q�"�0���_&��\�n��M�K7��gC��kޘ��
�����ϗ�o(���҅֭h�^�nw6�q��c�vm����,Y���ܰ��e�aӽ娀N�0�a���Thp�h�T�'\��yw8KKEj��F��:ۇQ'j�(U[�.�o^��t�DrN_�U�>�x�n�m�2W]g]�'Y�>�2��]�~9]DRE�X��եY8eM�y�ΨM����62Mtj�h���] 5�(/i�5p�2��߳*q5��"��HN�	L���J�*�:�zh�m/�YX]�Lu�/�c1�*���Xs�8�ڱ�xv!d���)KM�	Y���%���{�2����=H�iُFI�:�� *!�\n��{���.�v���5iҕ^���Yݙ��Э��i�E�]��҃$ -�����	Q��p\Q��s�N�C�G
�����G�T���a��]Fq��0�5����O;�M$ί��2Sx�j����3Ms%7�c;ҵ�X:%���^�w�%0��bj�wG�S-h�h�3��ە��>!n�n��)�
��\�m��PO�I� 1N��L���7ha��fK���#���S&�ն%ڭ. 'o7�SzZ8;m���Wn�]M�Z�¶P-�ԁ�@~��Q̺[�3PrG6h��
H�Վ�z���T5EG2h*�
���ZsDTN���4S�1PDMU�͘�4Ѩ�e�������!�8X�����l&�h(,Z�"�n�M�lP�TA:j����<�Z��JN@򹈃��m�4[�E�E�:,ƃG\�'m��"t�\��kjJZ71���-����)��)����>.�'�9r�P�5LAAH�rA0�liI�vڭ>.9�u�Z��4c�i9g�n\,':�u&کu�r�=F�5�3ɤ� �C ?��]����o<e�[V�N�
�\	��&t�6�{���G@�CJ��=lO�>R-���hz���Gd4�E�gw>�<���������<�R�M(�H'��]��}|�������qx��r�З��C�ТvS�/�����OI?��]S%EP���1b���w��)wfBj݃6��s�M��uEs��f�bN��T�,��T��r��,�^+2�؋�{������P ��w!2|B��/��:���.�wʆaQ7�M�~{!m{m���z���)����Y�����\�%�s!��J���`>'46��l;Z�g�&BMuu��g`�Ӆ�)�H�V�k^��Ӕ5-�G�az�{���z��`<{D&Ü���T���Vz�u?!�,ܝ_t�t��-�]�<���>�_w�f{C��ŕ奥+;�5��Օ�X��-1�o=Ρ�?0ب�����=�8�|!�}�A!�p�j=0����ۻ)<��>v�]�d�u��,��*�3?�(��-8���Ľc�n ��nHxm��΋\^]��Ra���90���^d*.ߚ�L\9��g�`���$��K�TcW_���Ƥ�,u������ٸ�p.r�pc��Nq����H���:��`!	��`�,���-�d�q敫��-�����>�ߺy����(d@>^i��ƶ�)��f�1RnS��� Ꝙ��.�Μ���'V	�u�+�5���p��C/��;2����|{$�a�6]j���Ƨqܾy����9����s��RLE��h���nV̲�$?��>��)��$B��`<y��� r�au�e֡�6���*BeV�
ObWe=�m4��Ol�{d���Цf�w���I|�Z��E�CUy��?��s���xNR�`YEP��R�k���,�������k��/x\k^�'�!���� ��5��):�1,���eI*L)�/�,;����b���ѕ�Kk�B�t�@�̜���ρ��	��ey��=���J.�s�2Hpy��=Yv�+P=݊�yKƾHL����>����#�УgiC��U���K�ȶ�We�eo6��嗉�ƗI���\?k���{�0t�����Cjh��$�0-C���N6�a9������gvɗ���4���s�@di�����k�`�_���0U,�Ǽ��ѕ�єxE"�huVߝ�߁�ZÏB�⠗�{W q���'k����WaBe���{��g���]ݑD��v�M90̱��qM��eRb��_7��>�z�;���,�F,3��=P0&�OG;&�躮�ӇZud���y�ߧa���m��J�ڃ�����G�{ٿ?��m��T���(Q�����lf�����Әِ��;��D�tyI�wE�!�ִR�b���~��Uf7�o��]�b� ��XW�ŏt��޹ۼ�p:���V�=.�@�ݦmb���b ����:�JAZ�mN�;�Kjp��_>|�?<���eG�HL% ��(�
�)I�D�G�׏al�q
��1l���Q.�L46����f�D�b}�ciނi�p�57٣�j\"��Zi����;O����EC��D��Aiid�{d��;�~��^��AɴC{�2/��߫�ܧ:ƹ�3A1�9������ɴ��6��5��ꉡ�9��N�##)��mW�=�Cfmun���>�u�36ĥ,��eT��	�$r��͜OC��WH�x[s�[#���i�yсv:��B��.�y�q��2�&�h�'�Fq��|��x/rˠTLD���2+M��:H������5l��h~����I�4��(�kq��m��-�;�|���Ʀ�~t=���`d����WR�,� ����v��?9�N�Z�f��2������ښ-	nAn�kk�<�"��?���8P����ӠNȈ�b��3�Y&C�[L��m|�L +] b)9Y�"�-�a�@�az���=�A�"l?ڞ�S�m'0Ww2��M4�a3q�t��LZ~Y�R	z���Fi���@]�������C�v�n[ԝ�Kkݫ��9yW N��lv��$[��f�0��tB�p{��y��O��1Tp�WOc7T���F�J�� ���f�_V��1)�nط2��k����q
��z$W�O��3g8�]���N�݌p�-N�%�.���|��Z?���BR� �	�A3 ��7�7�y�GJ6�uh�\��[���z%����;)<זH�R��w=y>;���v��g`w��sdl��MV�V�;<-���D;J��W:�X�V��	?1L�z��}5R͑�5B����s�N�ܥݛ��2�t�@�mt_�۟tv��Ba��1����{+��~f��%�4<����oV��Ň�Z��:H3�J�^<o�оPc���A���\ء��m���9��-R�cɠn�y���1דߖ�4C��|3h{�����`��OM;��&O����6��m���҃C�r;B+��j�v&}�>h{B�,���K�!���������&<�Z�?kā�M{#���{�}�2͵�$�PN2H���o�}��<]l�wj�Z�xQ���+�6�BPB9�[�.|W>���M�z�$R�A�p� �F3�E��\��[z�N�>��/|V�~T���2�$s"×!��ƭPB}l.�sj��X7Dʙ����9�Afਈ�Z;���=^5A\e	��i]:ɪ2=?B���=��}f����s��1�'����˔�L�;T��_<G�0D��+կ�}�t�W��|�rA��;q�~��q�ta�6�Q1[�b�pq8�ЏJ�ǘ��Oe����M���i�yл����k�ɛ1��rړ�Qi/�Wv���_>�}��
Z�I$`�f�f�3R���F3�3E�¹P�r��[XS�������-�A�k����!ۅ�T(�3��|�X���������tD�V4-_�QN.�H����қ�oH!� �hcL��[������n�a�j�dN)��)�0c�E'H��N�:�n<����N�EŐb��K��h��S(|	�z` �{ K*�5#����=�P�0�W���g`>sez۫A��#=:�MHĿ/� ��{�G��L�.��'vJa+��yj�˔����B��6����=ݛ�G�M"_��D ~��_�H�[�׺�����e7�bN���,�l}�<K�jW��xvt��H�k	���P�h'��ߋ�C�B�� c_��ꃛh$Ԍ����!��,�`�!{V/����c���%����a>[bu��ÿA��H�%�k�?/@_��j
}���VG]�p�*��jjT��Mk�a�r��nj�=�{�����p�V���b�*��w��Ǽ������,�fI��K7�,7�bK��{}��CQ�ƅ�g/�a�)UkU^<���Pf))�YQ,J��ϕ.���s�M���(1�u5;ĚuwW��kX�-�:�[	�c�d9��� ^.��Ā'����r�Sl^���3q`ivk�p�?�}R��w��
����A,W��^����� y<�σ��m1�|����{ǯ���/�bP� �����u)\��2��g-y���½�s��wS0��C�oH$:NmG��V��h����̂:�B��x���`3?��2�.'љ)=�_���_Fd�d_c��A3&k��%S������-š��^i��ۖ���sC���R�R��ƌ��q�����bۨ½:�5A��x�;�����Te
_�Oj���%�Mz��)���0G��ެ}̉Z�o.R�[Ϸ�D�ƽ^�RŘ�	�yHL�֍
Or�(]���ƚxk���1ld�t�;+o/=f�9�����}B`r�5��������ħV��	�T.�g1�}Ǆ�E��B�M�]�<i܆�_�|���y���^�锝g�ĲN�s�2��&gm�\	z�Uy�[-۲�\/?\�z�֐��/�	��!�;/�B�7�h�Ϸ"���t���4J��Ad f���T��چT��,�^���N͍~���L�#�УgiC�ΔED��/[�2(`}���ˠ�Zr֔4�0�Ʉ8{����SM�"8F�lėS��]GbI������ק���I�������������;"|��ۈt'1vN4������V�:����w�-Wqut��]{k��	z�p��-�X�7|�u�1���V�$�V�«Z!��}5���t�h2�ښ��S'Q��Y���#��� Hd��V��	|A~�q{�-�2�~{S��yh�R��T�����c��.���Q
�y�{���H&7A������3f�j$�ڭ�zޗ�T���X���Ԫ�ǥsߊ�^��+�eu۞��:C��z����]{��~��٘ew���Їb�&�����6�Lm<u>�)��׸�߹��nY��1ls�͙�����ݦC;j�@f!���D<��{��O�7d3l�Ny>���!�@�k䁧��[Y�*��;[���V"�5m�v3�.�C�4>
,���t�94�ΰvȻ�MBbY��gg(�ףw�tS@�%u;�O�w�~��t�2��{d���^=��h��[�x�hK��e��1�2�	d��YAP]����~h���;�3�����Ͻ�J�wO��2��iʪ�Jz�6և'Tͧ6PeB��y�k	VPz͜O^ǫx]]������tj߶esK�Sٮ���I���7;��q�-A�U�4���z3R�֭�,�_{'��8�<c���v����.�	�`�1W5{�Ђq@q�d��3L��=�F��ݩ�	��z�É� TЦ���p��n�=�-ٶ�b��D�7}1f���n�u�G�T�+uyc�Uj(H��@�נ��s@�9j�׶8���-�������D�x㜴r���u��z�7]�ZyZ�eo=<��;]sϾ�����~ ��i�)d�!��:���*�J[���^/l������(����,���<��Jt�hoʍR�=�0���R\��"��R���ޞX��9��$zf��Л��vD�Wu�f4�I�۪��d��8\��'�tE+9�R�-�a�@�az���a�<��!�w���ִNg!XcKA�ZԆ�4ε'�uL1�M���b��
.W'���a ��h���Kv�x�������O
��Y����˞�VM7_i����E�H�R�䣹����qxwn���=�Q3��u�'�s���v!P2C��!ؿT+�A�,t5mvt��i�oVϴ�Y�E���;��KA̾w)3j�@�ͺ��C���ͮ������4-_�Ja�ƲǼ7�۶�M�Sd���;�@���A�܈44.)��$O�ƾk�ڭ����^�6�>�v�TϮ��fu ��+T낂~�a^%�%�@/���� s�>��v����&94���!��:;z��%��A�ϖ�8�j�.ŧ�|О��ʹKO��K�!���\��m����������E.���]��M��xj]6&,JV�����j8���e�(�[%j�S5�!�� �����Sy�z2e$΍<66T���3z��K��-����p���fͤ���#h��ȳ=�o�|�̺�/�@QIE1 D�}x��~��a\��o���.��m���@̵Lѽ�p*q�j�&a��29�=�x�&��,����8ըS���, D0��I�k'�ۯ8��0�q@� ɨ��#���%��[����a�J�P����RN�1���@�b�)˃޹���r�vA>B��o>p7-��6/Qx�9����X�J;�������("�Iq�1<�!u���X��o�@��љƥ�2wM��Hg�\b���hR�%���.���z�Y�g��AA�k�5�I�3�=��-�&eq��*���%�Ps	�{"S�	�J��]�:q���-�P���xH"1����t4?hi��f��}Ya����z���Θn�2�pc1V9�RzH��ם��OW^c\�ѕS*;Y��A4F��t�	��<�@�]�a�vT��|f�Y�s ���:���6մir��~��N��!�LH�!�ב�w=K�~�:�
'e0�9+�Z�r�'��}��.0���}i�N���j���F�5���T,;]���6�^K���lĝqy�n2bY�y�ť�Y T�+�`���f�� }d��G���e+�f�S	�j��]K�J��.ABbum`Q�r[�۸�Rzﶒ��Q�)���^�@�s[���M�V,�#4��o��0���٫לL#/u,��{�>�� ���o�`�T܃.d��L	�,k���H�NV��0x-=Oǡ1�o=`�@�meXǠ�1T
ٹ�@��ҵ��t�{*	{kU�|��鯹XK�0B��%}ᯋ���.��^��Mnn��Tsl.��jY��v�a�@J��q��;NP&���8��3��"]�۳ri�E��B���Zb4b����B�;0ͅ��n�w(��8ėn0�m��ClvXƁY0�9n��U������i~��I��|��P�s�`�a̋!��C�J�J���ԕ���Kp~�ݿ��*ó�5�L�`��`L�\H�$����nƴ��>��Q���^��&6;������8��VH�E�H��t������`��(~�~�JK~3�����d��i{{t2���:�C[ x�Z���,��*<��vE5��tS���?���6ph)��+8?e�Bi�����ږ�������ʅ�B�ܮ�o5���z�o 4�{gl��قێv�T�;�.��2	ħ� �=���G6��%1��N�),T"�]��c�o��������{�}��W�����|}��?�������:\����#H�$ԁK�XO���X#���+{�M�Xգf��qgH]A-��R[]�N����U�I�I7b6�L+p�@��tN@�i�^'��@\tm�	>642���2��{\��8��.���H��1Oe'��3C6`�|rMMҍ^���O5��Ի�����,�	�Mu͉�Ouq�C�k��9h�I�-p\��u��{r���N �U�+�o�7����u�ZE����2m���(�٬a���{1�#d	w�I��tz��>٦��u
�8j
H"���T�P�y�4	��D�f3�p�Z��D�Y%�u&���"!�Ek�])r�DG1�KykwQ��źe\����9�wNM%��4�b�j���Y��4�՝+[: ��l�̼s�$��VF�5>��_���4�ǻ�|vFy�d��f���x5'[j��?�� �Qm��p67e�)Q��6�(�n��)��V.�5����ݕp���n��Τ�&�8�'q86]����ݯ�wu�ə���A�8���eu�]�n�捔��7'@�6���i�:l�s�$c���չO�b���̽�]���#/��(��A¬\��I��rV�YGOMbpU���W�֥g	���5%���w9�8���n�N�0}p=wa��J��j�Yv�l0=�u@у��q���E9+B�Ei�������M+�N�i�L�Ŏ�t�d,d"����\����C��7��32�3�E�{��ֆ����\ld��q��O5z��ă�ӎ�.�V١�GRVX�ps�w^qPq�{��;P�zP�K��em�3��0��H'���F��e`|��9�o�%eA/S��=B��H���rѬV��Y����443�g2.#���8=���w�wS�P�Y[�Y��n�ͣ���������sZk^`�ze���5g��.=t�'��c+[�	B������pu�ӅǼ��t�d���{�pS����4w��q��w6��ڽ�!F�Ӥz-�7���C����l1Dң�'��[��zY�M�����}.7���ۖ/];�XS�PA�b�㻕�:�q��IW�f�[�m�o����2&��Ci�4��Ŧr=74e�]����ӌ)wU`}�WL�$wD�C��
б���ѯu`�7L�w���풪ܥ�I�'V�#�c���#��r��w���*���C��y'ty�q�D�b��9�{gM�2E�lt�1[b8�j��в�C&���wws�����eRf��P��>u�'u���Ϻ,f��Oq��D�n����ذLJg3y�s�����[�����ęX�e���S�b�oouҽ?k��M�X��u[�
��tB�1e;&�bӸ��x+�S�qaЯfK/��L#t�K�X��g���c��Mn�9Fb���%���lִ�Ug���ս���(���$Oޢ�|��h �O&�9	���[�5l���^��r&��CѰrI�!�Nl4��(�����9<����[:JH�5A�#O �xMk�Ǚ�)����[a��͔�H��kK��������#Iːs�mTs,l<�Ns<�F�.���)�����#mF���4�s� �5F�A�M���������X�"�l[k�'��F��kA��ڭ����(71�71��͞ʉ�e�ڂ��r��m�͉�y��\ۖ�/ �U9'FŹ�1�6֭���C�,A���x=��QhC�ʌ��.tU¨z����p:��ѷ�x�$�͈��а;�:��h	Ek0�-)8�OT������0���5l���J�į�J��@1��NIa(��	�D-�#q�h�sp�uˣ�o��)���]��'RG=�pG.+#Z��ͺҷ�Ɉ��=���C�ndC�z`>QC���g�L���Iֳ���@�t��Os�m��X��[��K�\W��a=k�HN͗�~�Qx��	��+�v)�������0����C_"�4�~@�Srޘn��_��69�P͍1�uL��dI��Ք�������f
_����h��b���I�y���}b��;�XG���5�����w< ���	�|�����)�����ZJ�/Adw:�WC��,c��0���zGA<�Y,�u�䡜1y��{*i����B�`���{)���ڸ�w,�^��*rk���^�͢��F���B`<�ݙ:kɆm���\eRca<u>�F?�j���6�Q�mr8l� �d�b�,3�I�����:/p��v?V��ׯ��c��X�:L�p�;7�n++�h�p�uw<�.lZ�X�c>���� 円���T�{��f�X	����$�3M@�]/0��9�P��x#��&�D�=N�����?_�%�����2H��IϘy�^���\�������K�]�-.�H:�bl��{��Q��2:�Fɣ�y��aJ��|iV<�6�!��8��[T|7�"�/O��if3v;WX;�S������/sE�xӟ#7@����7ݱ�i�Ծ�Dd+��6���o	�bl�\��O=��� �7���T���t�~�^ӻ�������K(!C��p��I�m�k�<�-����kz�U��5c(��sb�}:��3mZ��m;2���H������O	o`wہ�K��:�vN���vF{X.��
e��y��OPUX�+��W���M�2�&�Z3I�Ҍ���S�է��r�s�z���o����~�`�耈yղ��\����%�s��w�빈B0L�V��I��T��k�Dn>753��l#!�@�
$�6P	��|$>��/f��x�q7�M��R����_���$�-L���O�p�<��ki�%,�Bc�'��C:Z����h�}ۨ��Fe8P���q�&IuFfӕ�^E*����z0� �}��a!�[��.','Gg�dm���b�)�R{T�t�.K�})��^�J��v)�a>ހ�sh�[�-�V���ࡁ^aq�"�q;1,��:ri��j�k�vQyYYK����|w�6�sUҘ��#��ݡ흇��d0��C��ƺ�W?��2)��4ՀwJNZ֙6�^q���p�S�eCj��b��72>��q5�N��-����+��)�ٷX)�a�}���Eͽ�n�����oz�^�z���宠��>r��;mn���:_x�|�s4]>�ܛj�>5��}oer5��S����RG�j��g��ީ���Q�7m�'��X �>v����ϵ�hZ�:�Ã�++ �-�w8U-���z=8��1m�}}A��k ��.+�~>(�-�g��k˼�8C,Oy�s��kPyER�
���- ��[��m�;���Ds;F���=yT
~�/�z�u?.��_u瓸hG��eش����xFc��x46D���r�Z
��}�:Є2��	9�m�\;����4��$�7���A�ș��o�i�3Fun��N!LȻ�&���S���4(!��ļMG��v��ءj`�,��&�b�A�`�b�v�'�yε��ד���b��%c�x��� TE.z�EcW�A	���u�PŻ2�k��֎����t�	m�WV3�;%��΂�r,D�S����M|T\��Y�*?0�;�@��A�����uS�I��4)_�QaL���,���<69�$Bos�f��̌
�P�]3^��mtl*׾�v솩vBGd���P~��=�)Մ�P��S�����Ш�7��<��� SG�I?i�u���W$o��,��D(���C���,u�˦�X��fPyV�
���(��>�=��񋋎�ŧ[�U̬��&�t�\��� 0������m\�+{Kk��F�+�")]c�K+��܍.�&��z���H�s?Y����o�������n�l��0�ҥ2�0~�I�"hӅ��F�:�n�#�w���d{��Y��k��TcÔ�C��g�}�ROW�m�u�`se1r�I�)��"�QC��
^��/\���!��B����П��Q�gi0����Ei�a��ﰛ�y��l�'^�2X��m2'ߓH�ıZψ_�$?���Ό܊1X5��vF�]S'��z�9D����ygO2�
�XH/v���n5�pC�t�f�Z�L)r�(�~B.Z�ӷ[;[�)
j@i�K���zW9NK�)}`r�c/s�w�pÃ��0Y�7&*f�,�������/G��|�mK2��Ø�R	�.�����{�5-�y����T�i4�*&�J��i�!� `>L(<A�6'%ا]����<��.Ն]�=q��ܽ�/2�ke�=5��a
���(\gO �}A@���>���ٹ�Gu3�eⷤ�7v�7\����CC ��&N�5�6�ʆ�f`0&P�.'љ)=�E��^�kP������z�~�+�cr���47��(ђU� �.����:��82�Bkw�"Es<�b7,U)�%��.�[3��/��};2�!(�v@�ݗb���
[N���ч�g,����TDg	�:4�ly�M���"�#l�"졝 K9>;�N����~�s��Fs=��"tޗ��Hw#��(��� ���W��H��t�u]� ���zzs&��B]=S�\�ۊ���$e!�k��5-lJ���� �eȕ�*<����s�^�M�U�ß���qj�Zu^t`Ռ��.��]bv�����Jl�R+FD��+����u��V��%��v�e��^D��9b5헹ħʘ���b�j�	Ll�N�%&\&q����"3B��.�`���w
L�P���F#]^9u-��}{U&�p�����~)[Kl�C�{Ɂ�!r��-�,+��/�P{�����3d���sЗ!�{D��0�wJ��ƌP:���9T�0�,�xn�Ɇ(�rk���T_����|�?ǨF?�����F55W5�֬\�2D���8�*�z����PX�]&+��i�;���,#��~�z{߹O�v��)W NF�Y�w��,���'�d����(]�Uz#��_���zY�Azp���2S������͵�Q|0>��O�����l�:�����XO��|���uO͡]�6ǜ{FP��������6���i�ڹ]W��Vm�	]�X4Jrf��������>TX_<�q
�{ �Q
�n_�P*��炴e�Ku�L}#�M��,J�^��61KS�����6������T�!1:ޭ⶞�̮�q�̛�ąWc�P���V���LP>���ra�q�nt�#
S����|gӯP�{D��7
�:�����X�˖eC��;)�����y��]��dl�}(�����u�;6���y�`}�要�Sώ�-�ؑ�.�����Se�^��fig|h��%�\�լzRg�h�v�L�f�Š<z���c�?��a��D�ǐ����e���p�*l�|s%��/|?Qy�w���#w3E�,%��r��o&���Yb� P{��������+�����:O�#)���ϹM�RTͶw}H2���R9A�f�'�5�]���$�cCkR�H�x����{��OP
�%bv+���%6_��5Z3I�-�k�l˦z�����F�R�^Fcս[�=|w ����� F��C�f�A8w��{�\O��#3a��� ��w)�0�����|j�t��{w� ��Q%ٲ�>�+`�Y�T��j��h��2���;�5�s]'�D�K�K.IRkk�<���������Δ3k�Ǎ��y�I����$Xf�{Il_nE�ܹ�kh��U�3f<�Agv]h��D*M��pxϴ&y��[�(���(Zg_
����aB2����8��z��2O񦡾�T���!>���6��b�uca���j|o:j��m4�>�<�cԛ��F����e�#���wR��<@���)-�a�u���{a;�OsL&���ch�h���!0�)��E��i9	�^��O�(�r��i��QS�Ӫ�}�l�@ �x0�a�	�q��ǟ:�=Vݝ��E��e�Y#Xˤ���$�r���u���������s�xk��.�b�k��s�dSi�;�'-��z��&�y�*�c��}ވj}3��B���e�k9�D��AC�\C��)�Fu�z��7>׻MS=��^���C�hm�j��8��aÞ������5\������(h\W��|m�9�s��b����&��"�4��d���%��,�=��typ��^VQP�>��F��.cf�1g�/D�'�ڑ��������f��q�b�1��Aѝ�硎����!����<�J^2�,V�!r� �<4(��c�q���t�3,�4V���^*q�jD�5NdfO[\@UL۠�j�C��o^4����r���S"��_Ү}]n֙� �B[���麦r���բ���ܕ�,4s�̏Od�,��[U�q�֫dy�a��� h���6��yӵ�mN#P�î{�t���N�W]��l��ݳ�c �W�(�*���IխЃ��2]Z�V�w%a�	�k�c��8g6U8y�@gv�Y���u@�KU�ǿ:���2�je_��WX�0h]FNI�C�=0���Lcͱ�!ﺑ�h3/7��)�_Y � ����.�g��ذ��vר`������ÞC|����MwX�v6m�!8�����ۜ�6�r�W�X!�U�d�WT\:�q����s*X��9�.3s�Qf�1��}fY��vInjЙ'�D�W�W�*��WvB��y���-�����[���ob��M�ƴ�r���A��n]�4�Θi��&@�LV�SQt���2\���S�S�-�uj�7eT�6����$!��}��G<�Gy���ܸj�%=Y3l���&�Q��<�Tچ=h��6G2�ǐ�D��\W(��!��X=ɗ�wOA=㴘S����C;�-S���d[�S�$�Qz��zKGjO�xwf�z������t��^��ζi&ۻ)�Z���ث5�f�f4�I�J����<ʕN�߼d:q���M
���
:8G�s��݋�C'��li���#�W�MVJ�B�⠗��*�a!m������y��Q��ڮiS#�-���-+^�݅"!H�/��+���b��1b��n���:���WN��&H��-��j�oL�7P�w��v�v�!<��E�Q!�"�衽3%�\ʼ�Nı������n�����{�
�H�V�R���;1�.��nǶk{��Ȏ�G]���7Ko�&j�W,�̥ĢÑ�C�ꇶPk��if��I�5J��q���Y�R��@�����������C+p~�#������:a^x����v)��q�T1�ܢË�v��]�<&�Cz��*�*}@�Y۪U��U�l��^]��t8_!�>0���d{��]���ُ%��x�z�0��'8����!�*����I�ʇD����fq��5W��.&7e'�zǦ����Y�'N��5�l�Xu�R�:�C�r9׊�P�k�>��t�u�,���a�qw�}{S:�f*�C)�wʋ�UԮr���iR���,������@���46)����Uy,�=��FZy<+B��A	�g`��l[�v���?)��)	�hФ�+�����xH�I^�m��L�f��i�}gh���i.%>T�HOex��ا�����6^%:Jֱ�4����}��(T�z�FNc�}Ǆ��|w��ڂt��	�B~�pFv/+�x��N��[�{�l6�zcL�/��-�%J���lg8l����-.2r|��_ܯD"�u�`���}�_A��@�~U9L�k3�(7�ܜ��o6']@�S�歩j�w���m%Z�|���Ju6�m�[Bb�U�3��mmt������qi[�oe��a�7�k6�Ί��t�τ���9�S\�;�\�g:�G����;΍G]�ҫMs�:T��{{��d����{�W:o�U(���ʼ����:��|�<��*/��N����k��T�2�q�TcKB�"Ж��hR����S��^��$���.��IĻ�l�?��α��s\���J�ےE`��
[A��S�������v	Te�dw:�R;��@��c��.1���*�.�}�����@p��յ4�o��[+R�XW���{*	{���9�J�Ǚ���)�k�,���f�{`��7p��G�C��i�L3n>�E2�f<�1����Su�c^�Y��]�ݏ�b�ӭٞj�ۖc^1a������x���k�x�t��n�fٵ�1;�}13��s��|������)�vQ1^�tE�j�X�c��hl..%M�y�s�<w���m|6~�{U����X;w9!�qhO�i/��ӻ雗�xg���,���`F�W>U���ȰC��/G��CZwqS4vA`{�,��R]�ȳ�O~/8��2�o'K]�A�:N5�t�sKh.�##)��O����͵)S6�;(2��2]r���|?O�۟�������|��������o����Q��C�o)�uzp)�K}N
��H�7�%�cd�d�Q-��)�SǤ���Q*��L\
�o��0�i!����֣��X�m�JE�ZZ^Ǖx:�����z.�N���]���u���wY���I+,�æ؍`�N�����5t����c�j��M<�5w)nX��;���w�.���d��Q�T��s��R!i8A�op_y�r�)�%��٠���_@�Q���F����.��,*^]i�VE�7hN����A�7tچ�Ww�-���,,���w�u[գ4(s2�̚*�7��};|�Un蓨�pKjGP�ue\���J�YU�ջ'�[��ھxՂ�-r�y\�����r�3�����p$��S��M�ЯNt;e-��hm. �Oz�1U�{S9�m�B4!�_m��kFWM���!�a�.��g�E�}����r�t-f�[2�7Z~����Q�������ol�d͙�,��-�dݧ�+���Po`��X����>pǎQ��ٕ5��4��'aE�q�kC��n���=��/���������=�(*#� x��P�F��*�ZhU��Ѡ�Y�#G�;���:m<]�РCL:���D���o�4�<���|��Y��:��B{o-�˙���ѣ��]D�љz.�
KW9B�˺Ĥ�������"���(i��L���_I�6!����]yJ�3rCƊ��B�zܧ�`���}�J��C�,X���W:�u����rlY���!�p����(.���������i�� !�n�o)�v��~=���!�.���X�ul�'�Z��GKZzQ�շ�~�ќKg����p�gfǡ�C{Y�ȚY�6{��e�ǫ�1��Y���'=�J����ܩjꕙ�D��G�E��G۹
q�!�K���|�,�Ba�340h��?.ڇ�zg)��&�A����{�����'EmR�o���5����5�''Q�� JZXɗ�ȗ�%���R�ޙ�u�AF֙����F�>]N��H�|�.c�wB:���$���q�&�1^�+uʱc|Y��F�*�ڛf�I3溺�NbB<ʔ�Iܮ�ux�u ����>��r�V@�0������:\�v-�JdΧ�1n�N�k���U\�����Y��qL�$8���_	z*�ݨu��U��<�s�7M �&���3�]� >�׀c�Ǩ�X�.������\=z	��nKx�A�źu�(�C�-�+��� ��Y�ŵf�p�\3���p�,V�{ը�\���o5�ﶯ���i<�˰��h"�����+[V������oH����-wE� �����]��k�[T�M&��n�u��P`���fȐÕ˫���	�.x,��:�Q�$����̝l����9�������1��L�Rr9�G �6����r�\�3�ngP�9[&��"��0nOy&*Ks� �9Q�֎�:щ�X�A��M�T������1���V�PQ;jۗ �bk���Z-k�ŭG
�ˑUFڊ�*�3U�ms5˗.#\�\؍��U5��s��ش���\6�TQ%VΊ��:4�����b։劢���S1RRm�Ţ*Ő��p���&����r�9Ay��1�&"*.mE�Y�����ېj�s�"8IQlj"�14�����Kb�"��e�Z���
��Z�-���1h���T�T����Ӄ�����MS2F�*6�r�O6"*�������L�r�@��؝���D�n�����s++�)�x���e��r�Н��P[��K�
l�zr>��1�+���Ҋ�d�V6N��D����3��Z*qmä������V'b�#��M��6+v�E�c��y�������ќx�����ј��z�����A@��fL�ƭ�E���w�H�L�g�N�yH@\bYc�(�2�e5>z��VW�ԭ'�c?'�N`������O(�s��s�Ŀ
�B��K�s�'b��)�$�5���j|��\�� �5��=��ܴ���}%3�I�}�e�kBc�_d;��FP&��r�)�\�)P[\Ú�����ٻwɦ\�eV�+���7}�K�#��Bm��gs}\�_j�i��mO@����2�K���:�B8�<�v��1�v�&<ѽJ��i����@`�Z}G8���\�ՓM�;UsY�E䅒5��{ʝ���6�o��:읒H�լHt�yċ�^C��:|B�P4.�uP�urdSM[^&-e��2�_b_YKg3v�p��
]*ޭ\�O�ܳm[��٬��ǂ�(���ʺ��!/ʲWf��ص�s�ZA��L2�e�`w�}[c�\`���Ph��(h\J�Կ�W���]�LN&��/#8f� p��&�@����SO����4��������;�2�O�0.u�r�o��YS���'u��`�PWټ�>��j��YLE��+en�*��aN���ѝ�E���0k�C�+����Vn��+�	�0�u)��'`�cvv���CU�i`�������a��@8K�6��1�Q{�9�5��r�i���gt�hZ���D��7�#X���N��3Eی;�c�ĝe�Nդ�g+,�Eb�#+v�}�`��
�K�!��-b&u}S���;��e�f�����EN2�e�.N�׿���r�_Wwg�����p�m�;ǰ!��Ƚ�\����kH�	�)�*�Z��_6�fty.�-�R�g��e� [:y�������'q!�E5^��r���݈l��{�?W]:�At�Z��	�8�Z��z1���/P�3b
ȱ\eB���K-��nXޜ�a��M�Wn��̙��}�C,p/�Ru`b4)\�,)�vK��L\:�q��l�J%��G�a���wH��0`�K5��'i���{$�5y�$�b%:Hȥ
x��*z���c�\�[DTr-���Z%)M�:1���@��`�Fܻpi��L7t�L�1����E'�3�M�L蟯�+_j�)�r,�w�����7Z;`F#؄�� �y�ȦTuT4��I�|��|�<��3�FȆ�q5DM���\BR�?*n`�bہ�)o��h��752���{��W"�BoK�Kf�H\�.�d���S����価t���4mi�6��(����ց˄l��'eG��Z��PU�'e˖�η����YP�Q��bS.Av~�n֔ťe�i�߾�]��h�K�c~�+�%�r� ���ڠk��*O��:�
 ���R��V�v�K�_9�P�g��,�I뒒Ƃ;P�Bxwf��8o�G�?&��k��_z��Ū-�ԍ���f��X��E��<ʕN��T��}�P�Z{�CS�^��ײ/���a�#x-jg�mHM���BՅ��_���{�PK�XU�V؝nj�n����ݑ*-��^Q9�Ѩ0A�3�O�9N�jY���XsP:�`2��:{��Oi��^��:����?�w���Z][�g��.�Z!0g}���쓫���rKbK�V��s�{̧����u;t����1��ݞ�Ξ@חx'C�whO�0l��#�,�G^�fZ�:�"�T:�Qo�HD9Nm��e�N�U�6�ƽ��`0&|�Yq>��I��k�ε8�B��5\1»|eF5��c�C���B�F��q�����S>,;'�Tz��D^(�����h�Z_�p�6h���kWt�Kcv�=�eT�(R�#G�={zq���C���^!xߖ�Us{�n_0��eC:�Dj-͜�oQ���=r.�J��M��Yxߚ}�u��:+]�����'V�w<���]7�Hm�M{�2Q��.���Go�]�h%y\�z�/T ��P�L�}�}�����}��Fs�&r�i͈ts�'�lz����L&v��b�.��nj��sؤ&UhФ�x]r.z�w(��뼐-��.ͧ��;6�s�[ռ0)흣�[Jq%�B{*|���v)��%1��)��k9jx��s�-�MXa��FwsE��ϝ;��X�����x/���x[At��8#|�c/�zȷ/��QɳLF��S@?&1,���e^IRa@>��w0�[[��"!0\�.Cu��ʧ��c��H�d"P�F|E'L,{�J.��O�ٱ���R�$A�p����A�	��4!ݥ�
ڹ�j;��;a[Z��Gexص��C��*�{/I��%�yt�~j8�x�l��r!��V\�ݾ���0{li�p�ƶ���g:nEh%Q�������w=ydg��c�7��R3��}�.zj�#�t�Q������j�uQkejUoyŹ�\�PKܽD<��״���Q&.,�#�v�eyr�����H ��a?���h��q�wΖX��+L���q8!��mԳxUui�z^�>�z ��j;r�K�gb\3o�!�:�^�a��<�p����B��u�-���"﷩>����گ�0��:#��9��*��R)����X�#\�	��f❋���t_%���G�: �`3�g�x�vf��w��:�}�2	�ɣ)��
L�s EWw��H��oHk�v% ���
�\`}�6�cO�L�m���?������JzZeY3~<���b���,#���Aڻ���'O�7u���s���t���c#v�����ᅠ q�v-����l
k�2����S�?Հ۽���{B�A���Ƚ��{]�1�w3EvI`J�r�w!����yΛ|�*m��̚��p�C�,��T�� ���||�9�����͵IS6�eV��&�Z\�^^����9�`2S�����C�EA�U��.��-�Ò�"���g%ޝ���%6Lٶ�,�"R��^�U��/,��{�g{��z���o��'`p���x)���<+�\R ��*��9��:˱ֲ���QG�L��$f�_�O��$�����&]yV~+���_���C*W�q�;�fհ���!��_�S��ħVH�T����#�y�ȸu]�c�������,9��.1�rf�QJY�z`�R;%�)�d�q=�i'.��"�[|�X��~��������<l���C_�y��X@�s�>�� �F�03�ܞjOgT�[&��LZ~X�A.�	�N���#�־��vމ�h@�}�}�Fb&�p��� ���gX��bɴ�q����	�ucu����]�0�>NcpD�L��_
o�t[:���Md3�@7s�|�n�\�^U��k���8��j�uj�(~���Ku}� wos�6V$]�Vh���B����w����XF0^�ֱCw�\�VM7_j�k�����:}/e�y����z������H2m�<��Z���$^�(��t.�G��P��_:�MH�6h�~��N�gMOx2��k�l@�����6�~W>��f�طvm�63��A�����b��j�X�T�z��4����f�Ja������O�_��\`���#�?q����A7�Dd��Ĥ�+�������2>��T���df�P��Q1\�
�ԏ����0��ʟ�g���W�|<�lya�b�Pi�n�uN΁s~ۂ��r��<k�aq���r��ǡ^s
ˡ�8� Ax�A�4�"`�]1m��v=ٖi�(oI.�U�&ZЋ����G3ϡ��=.�1��^�<� ����
ȱ������WXݭn"r-�w�O�Uq�	~́Y(2F1�sgV@�t�9���q���%'���׶Ӻ�c�dѭ�B���BLV5a��vi�2�%Ռ����C*.�����g�=��&f�6,��bw"R=y�TU��lP#i�GWj�Pwo��.��Y�}t��&�8��zm{[òP���K��)��aO���k�nس��P<-���iY���������>��L�v▮|wCx ����KV�һ%�a���I�����%nr��I�����x}���;}�ӭ�B2=?B��r�N�b4)X�E�2�lꋇB3��&œב:@�u�#��:�]zas���f�>����&I��N�#B�ʢ�]ݬ�<�˜���j�2U0B�[A��oD���!�e;r���s�@�K��Z &*�Fr�fgsS=�p�"��[�A\t�zw�xa��PB!���'�pG>�ʻCR��&��Ɇ�8.���n�ɶI�08����9�B\W(���?j�5�{�	yO�Ӧ��X�u���Ӯ�e��B�E�R�\���)=ZRX�Gj%�y&�/�ƱO�Xv���B�W���.:���9��e�\�=�-X$�%I`Vt�*U:�A{�֯sۇ�-�-���\��,�W�c��@0�WT���������\�_��U�B����E�*�-�T�\���|�ؗ�?�G��q�Bg���3,�;h��u*.���q�i��u&�� OmU0tq��>Z��f����a�O��w�p0��[0x��뜗d�X�n��E��wT�b��.J���	��-���=�~;�gܴ&�mI3
��\Cˏ�ge,xp^m�'j�]F�]a�l�^�k��ߴ�y*�
F�n�C�pdL�|﷔�D)s���0��c����kT�S� R�{��u���-�?J���\ŕi�-+�j�T�s�yv���>��p_��T�v=%ު��xF6P���:��p�hy����e�?��,)3:�,������P9�0D�O
��zJ>#�*v�-m���yc}�Aq=�JX�Fg��n|��L���ڰ�Q���kNd$� ��VHB��[�:l1p�)�D����=N�������s�\� ��H���{��j�Ɇ��5)^���,���Q�[ӌ�.()�ҟ�[yx>@�S�E3ǰBli&9���9�B��J��KsS��/ܤ&V��O�.��R�8��\7:��͝ס�V������[HN�4��p���^!�s7!	����,0)-�q�u��Nx�C�?ƞ������@j�O�bN,���pB|�f�DA(�dhe1z^�m�s�.3%:��%�u��˒T�S�_8��s	����$Ia.��.t���&�S{/6c'*�+T״��G%C���0�0yγ�����S���^=2�˟��ff��8�xN�L��0Ac^�	��l�(qU㊺^����~d��>]&��Ƭ��W�~�h�&)��)J�;�6��v$&WM�� J��CH��c�99�:�����w�K��M��]��H�m=�uk�^�u���"��9���X���gX�Ri��/�b7p]�Ҝe�� �ё㰰EN�p�2�ٷ��c��D:�1�^)9�@���k��4��k�SE�ɜ`Z���v	Te���Ю|��vx0��QC�_pۼ෵eON;�8!����u����U�QkejUk
�J�}mm+�jh�r���/��u�iWrʹ9���<9<yF�������:)��t��Y溆���{գ���\�y<m>�«��b��1چb�����|`8w~�Eݣ_�붋�\��PD��[�w�m<��2��̢�lc�_�8��LW�lZ��!��ýy,/2Z����o1�7xp$�B'ec��3]&���c451F|�Ŝ�M;O>�H؊��Φ�ћ�-�]N���t�sKH��ZD=�O^�ǳ��5�w3EvI`J�o).�Λ�d���)��{F�թi�<�V�k�����/H�|�nIf�%L�~eWyc�P���4���k��wߡ���AWٳ<�ክ?s���h���ǧ��0G�b��s�I�6&��[".�a`����[R�&�Fi=�ޘE{�b�)?,�'�~c&��������w�m��c�܆���>�
T.o��Kv__X;���T�n3Is5PH����u���<�q-�Ui�U�]R}�m@.ؼ�������9�.&������f�p���]�5�w��Ԙ���{�p�Ӂ�q��n�e��\�1�|��*��#���S���H��k=f�����E�9����I�1,��I��Gc�P綈Q��4*F�p5��6Y�V�ܽ�}9nͨ	�`�iH��^~�N��xN�]"�PIRkk𬮟�h��\:�4��ҵ`�zyٻ}۵2��x�vle	K1�0�)�`dvI�;��O�9�NVy��h���n �89��2M��{�}���?���B�t!6И�۹�_A�0�-�jz&-?+I�[�V�m����¬���ǀPFi����l�Q�>�#�l<2�}5����|6�źy����2[�O��)��&R��w:lw�Ļ�{c�G��!��;�'�T+�-��ϢH��iE��>�sF� �/A5�v	�_�����_���vid���P�d��:�?��/�(c��tm�m��u�Ψv���a�Ʋ����9ƫ�K��@���)vk���W�ő��]�����涘t��C�P����h?Q�I����0����@/���N��ٍ{��k���C�R�,E��pQ�>���o�R5���A�����N�C�n�������g�����~?������{�/����Vgi�l��)o�29^Έjv��e�
�]50���iןn͘C�	�5�6��+�R&FP����9��Z�RΣ��i�]0��UuL��P��Q�Dd��|ﺙ��������]lQ싶 ���]Np��_���u�7:�;xh�����2�N4����1�8_wQ �W6ä���t@���^�������	�0K������6O��h(�#n!���@ҹ[]{{G��Nu���f��J2r�v94-:�i�6;vp�W�;n�f��W�h����mfty�oVݝ��u��֥z��0�Z3�v�y�p!:��Y]���j���w�wr� ��Cx���>���+kN����Op�4�c�,�3"e�t��v`v����/�PǸX��nZ��w��5����EBA0==��
�7�0Vowt�ڱt�.9}�!�b���a�Տx�H#�g/+31���y;��H3a��f�gt8��3��U��c�Y�����	Q�%��y8���T[ά3,Qק�|�B.�q��{3*ն�a�RcEdX���5܇f��{�vm�B]]l#C�W���e<�xChiYӘ�Z��U�*�	C �I�A��N��ej�z��[)���ŏiat�u�v�r�H�f�;&�n8vIoEk�>�r��d}��mu��+��kr�GB�nv�tbW�V�V7����'�6�f�ëu���ۑ�qV�ReێZ���ʁCz'��ms�3 !��o.Y\����TBs;1Z+��9�����F��1�^��8j��G�D�B�d$*�Z�l�Y�:U�v��B�Nm�V���Hc�[��״rX�^:�c(у�W�1f��bkIΑjA��;[F![��0m��q���F��b;���⠒��I7aA�s��5֣\��tvL]���f���ח���-[f�{D�\�V
ᗼ �Ky�
X��qkCM�ַ�iX��I�w$����1�V%^��U�)�)�LT#�q����LVh�y��I���Yvjf�HR�f��j>6�g�b����)OJvot���A����*;�q\M��n����0��Ə\z�������TT��:Y/{B"��\.hX�B�K���V��V��qȐ$��hd���4�PH��Y�:�r�Y�Q7u�B�+e�5�Z��#�ـC��n�����V�� ��k�}�{vG�����Z�X&��t�턑Wb�;��y�T"��A�]J2VDYw.���s�f7d�� w�R�Z������d�Dǩ/��s�L��fjar��;e�F�]����K״_K,�UӂVԦ�`�
�dg;��Qn�����\�Lv�ii8םd�]�-��*.�X_cꂞ��e[�_-��U,sE㘌/-��ܮ���K��"�hd��Vi�k�(��~�(��O\��>x����D�ڊ��vo
yA��
ܺ0�:���#[ob�S�rW�����)�����9b
ւ+c%15��1����b�A�+����m���4�$EUSUf)���M�Q�b��j��Q͎[�,g��EES��Q�;�W788&( �j�+�7	��T]`�ŬM��\�"�&
�"�����.gW-%T��Z�$��Q1')*��%QZ��M�j*"�C�h����c�*��IS�1$W1���s���(��Y�j(�*i����" �Z��"��PS�9��+m-MZ�Qƚֈ")��i婦v�EDkQQ�b"B���d��
��h�����'QZ�%TDDM1LAV��*j�*'F��t`�C���j"!�Y(�b
����EQCD�LC1p�*��M�5�E���i堈���"�
�"9�Dgh���i��E���[bi���('F��4U5���^���u�uTn�Q�cM)�,��É���[��ި�f�� ��EII�E�����56��(4�-�\��:�q�{O�>�z�[<t��m�k�e��
24��6�!��Hd a��h�E&�)��E0�#�!Y{�SMU���,��kA7T�!��?���Wڥ������h�� ������o�a�^���̿Q/tX;N����
�w��1m��F]�[�_�C���C`���!#�U����Y*���{!V������86������(8��b�\ ���>l[+qL��sӼNI�/�kE�c�;�e�V^�(���cͶ0�}ka��P%�%Ռ��{#F�d:���7�j-���[���{�f�j=���N:���v�;�X�ˢ����v/a����)͞�%J���'�f�m��_sK�o3gi�y^Q��"9�]C5ߦv��n��M�A�$�b"T)�F��琇q��z\v����;{<��j��a'"��@3���t���!��˷���;�RdbBL�B��Ʊ����j�k@�t�4�Yvk���CG��<05��uǇ)��?��Eg�Cr�|���'j+:�So<
YJ��`E�*m�u�c�|���Cl��=yߘ�V~$ uXk��+ݺz�O�Uzv��DZ�{[[B�����89+�@j9r��PX���0��٣r|��ojm���4��VO���I�V�A�¨�7���d�R���YxĦ�ʊ4X�
�=������_�Z'���l�(}�>u���^�݇}|ww��߲�5Ř2����B�'H����� j��/{�V޷S� i�D�����#L��;�Ep�Zz c���RsbNP�`Ĝqw�U:9�+�a ��Gh�:l�����ߝ������e���Xv`�ɬ�uH���4-'��;���{�PK�Z���Mݷ!�:����I������t�����g��f�.�@}Oյ,�kݴXsP;~J����s�͘��-�hN�l䭨u$�jv�Cv����e�Pg8�i��\={D&��s�쓫��Ɵ++�V�&{sa�y�0%���.��L˴�lk�[9y��gGzt�zO�![��Ÿd�:����2���9S0��^(wH$=x%��˴�l�tW��X����qm��2r�R^{�_k	�`ȗF?N'�5�m���|�(8�ns�`��cOO���MC�.<��7p;)U�̳6;#(j�t�S��8�sI�_{D�K[V�!k�t�(R�%G�<`!(x�%����r�R�T�C��m�Bllva���s������Է5y��M�9HL|�;��#�r�{�k�Fr]=�B�Fc�M<6��; ^�0���!>��ا���gͽ�Ou���M(ޢw����ZU�Vż�i��G̚7��c��N�F;��[r���u�nyki��{f���6M��3��`�Pl6�[~җ=�tt�33Dvi�����kݧ���W���W;:��x����XơX.���F �$�wk7~��h��پqm�?;w�����c�EP�ػ|_q�=z��Hqm	�i��~��$}�0��������ĭ6��k��$��\�s�2��&����}�K�̜z����G��a_��:uc�R�H�"UvQ��Ȣ��E�s�2��P�_��hw�u,��;��Gw*&�"x(b)٭��!7W�n��B���*��]/e�?7%�.�̺m��'z�Î��g��3��������kH�#[��SI՚�`X����2��;�VQ�*e��nIf��]3v�ևy~��H&7C<Ah��G?��/��[SM������*��m]ޤ�u5���|���+�>E৹{�iWr͵�l�t��:ǈ�.���&��lG����Q���;kQj0g[�u�6��O���T�2چc����A��぀�y�a�cm�豗f3���Y��
�OC�ݐͳ}(����ZeW�Ń���{�]�c,�z�A������k���bT�{��f�X	��F�ci����$q�v��n=�o<	mz*��oN�XD���F�]��x�xcZ1c�G38��-��BL��mVF�Yݭ*��
�1��{�I� �b�ɗ�RqF��Q��Vee�꣏3L����S��;�^��mX�N	[t�U�H
\�5�����\���u����j��'$�� &�m���g޿��?�̳�t���2L=�O��ydwP֝�/�vz���r��̄Fl�ٮ�m�����:r�Wܥ�`�
X~0��㏾ٶ���zK�dͯ=��Tͮ�[y����������Xs.7!�6q>4�����=����/B*==J�%�����F��|۲�x��u��)��RC&�bS�g��ݾzޭྲྀ;��_g�K��-"!�9�5�V��/l�A׵l�*1W5�A8�'�L��$f�\�I��;��<�{w����qw���DV�B�Q)ٲ�9��ƐD��<����'�ħV�E2IJjn�<�Ĳ����Y��X��5<��d�[̝��ƈ���L8�wQ����r�<�X�n�}ܶ��M�w-aL�y@z|�>�h�B<����|��8ו���?T?�Q����%t_^�s��N<:s�.O#��#=>�|���ҏ���?}(�]-�ީ���VF�7Ys��[��'��k(U��Ϲ~8��qO��s�J!��@B�y鸿���ri����+[X��K>>?cE�,Q� ��G���r�y���LE�D����uC��[y��>ߙ'��^8	a�����8�et��*��z%l܍7�&Ý��ˑ�Wc�����/�3�X�%\Ы��1i���MG���p�qr2�p����{�͖�7ln�W�r��E�t^i�E%xe7����C���=4��=)8����z)D{��l��H���dชr�7�_��7�u~#��wf�<��\Y�Rb�H��(�é�k-{z}Tfu��a���Ue[�����jO�i����Bb�Y'�v/��h7���I��]4½Š�b��m^<m;���O&xu�����1`Hz&\�����^R�d�wPny;��{�Iv�'�C��ݲ�Sb{�ii��̷�{C�U���6��g�62T����>�ǲ�vY|�iyc[�����f����T}˥�@/�i�y��[!�����E��=Ų.Fi���R�`���W�\#){3�ڵ��b�^�p�䌆�y6ʺ���;�#^�p�'y��X����/k��v$o!:c���S���vOV�K$�m�A��sop<=&]}�	U�Q�����޼�q�3$:XxN,CƻJ��MB2=?A��r�ʅ�B�)�9�����Նc/i�6�s+��y����A�k�0����)���"!2N]�:og���7�'jeo�gد s��Ld���n'V��VVb7����{���'X	���V�J�����]
�0���4�N5t����5�bWyו�:ʮ+jm�y��
�LSeb{h�*_IvL=��Z�1%���6se�:��|p���.�c���>���F�%+�Ţ��~��N.�l�	�8�o��������L9�n]�4�s�d]�v��R,dĮ�C��aSr`&*�=�����P���W�+�ȟf0��<��uF<9�4�7��Q��P1��4�&���JO`q�d]ct�����<����ÁM8X�<d8��`����Oz�(�X���SS���P�c��
9�[�9r���\�HO��7!�ɹ�㔔�]�Ӫ�7��&N=�H�����]�P4��`�E�,��T�u�����(��>*v�U=��A��K�B\0g��t�t�<�An��ʁ<�-XQ+\P�ҹ�r^��v�.��H�dJ�c:�wj�U؝j׷s�p3_���p؞�a�f�����UQ���鐭cyݭR��e:��p��Ks`=ֽ�r`3P����~�9.�<�p��4FF�����ݲY�r5�(���^�.�{�=���b���ҡ�y���M���ɺ�}������&�Y�H�VU���~���}����3�����>�bU8����oMV�9��?(�$�rغS*���#X�r�$�Iw�����Fo�cZ뫫��ͬ�o��s4�>�m\�756�Trf#0;pq�9ΧR9�q��^M��k4δ%9�D$�z�E���+/�F���g{6�C;����t�塨/��U���#��5	ؔ�&/���kNd�� �VHC��ϛn74T�&*����<�u�ï�� `�sE��w"���K[jP? veAfP](sڗuhD��a�����áy8��宿��)�1e�,y���|��a����a#H��Y������k��K2�,Q�A�_�]{L��p�l�G��~5b]%^�U���w�Q�c���˹�f��~��x�B*���F�(��8�֑��Z:v.J�5�p�+��;�<P�8��%P}�gW�-Ԏ�Qa��<cI�.k�E���A�C��1��M4x�}���`ї����U�z�n(�!Ɋ6���q��o����ؑ�GU�J���".�[�o��y��l0�7��*������[T	F%���DP�57��;�KRvz�l����n���NC����3��L���T��4���*���_ef5�����!�&ࡀz��e��9�����-+}X	�^��	����g�ea+{�Βcb�����d��ٵ%���+C�Y/�wi�D_l��*�Q�킯1�W�Ft^T��U�-�W�	�����eC�9[�W\U�\ow�?�uMwQs�~�:�"f�fE��O��#��N1Z�rلe=�V�
���WP�;͆�o)���/�3�r�Υ�_��̉l���ؓ�W���M~��ޞ�m_�.[����G]!�a+��9	���ި���ގ|Fϔ�a��t�^D�Ѵ:��q#�vv5>�h;Om�c6S�p:�)+�s&��+��X:o(��tC�o����Y3|�t������]�{�C �rt�����Z��0P�*&MvE�A�;�61Md�;�#�s� �$�T8ӛj啍��n��`=��X�ΰS��/�tY�+.��
�D����'8OZ�{2@��2( �^쎤��o"��FN���1k��{U>��q��$e:������UJ���m�̇����L��k�R ������6�G9:	T�Jo���ف���ŕ�VF}'�B7l9g] �bt��-�5׎�vg����tՎ�6�g�o��-���T�O!_�7[��vQ��v����l�q]��-D���p� �cy���X���<��2�P��
�ڊ�1���#��4d�0Mc��#*�W
��m���uHP��#�rV�>wJJ�r��"Ze�MK����H�\Ef%@����!lBێ�����,m�3NV���o�!�ot�5+
�*�l���=��������>ٔ��|b�k��6t��soT��̑�fz����%	w-����Qf���-�o�i_f�fI����Ȍ�#U*M�ܔ���i@5C6XVz�e�\?]�P�
�a޸�����=��Qr�y����<��0�턴��,��l�s��@m3���&�0�!l�ó��;x��M��o&�kDF�wP���β;z=�Q\v�(�G0���uz�W����r���t��ә��h��u���3A�إ.xEL`d2�����h��2�K�����y��җ�(<��"BDF�nYK:-Ί ��*�;���?���=��xV����S���czl	���,G���s��+qM<��v�q����fY�b�-��?eª$��ww�!��:�.���]@��.��Jn��1��0uK�n�����kk�5�;�["�-���L�8;�[�®��Y��B�f��+=�G^��{5�P���#���hO���H��>�n��Gj��K5���ದ�VEwK��Z��&�FEϵ%~��	jU�A��n�5������\f����͔�� {d;��,�_!V�ʏI��θ��h��-Fd��<;:�W����� y9���[�<6�Ƞ�R^f�k������\sOK�5^|��N�vdH���B�h�{��-�j^o$�]�R6�yΘ�o�RJ��)"u��Z�̋� F~�	u���M�ók�2#��U��DG)T'넴��-�RZ_wɺsb"j���	��W~�ʷ�+�O�A.����ħ���4i*K�A�t�������$P+Tݴ�,nu��>�]i�46d�4p�]w.D,�SJ�{nt�a��3.����>�`�Sb��] d���4��Ӌ#�|ޏo��������w����{���o�����^�`��.'kے������q9��Ѱl�'j;��>lV�n������a�Lpp��t�Hgu�BIF�F��_t�r���~��3�lzn-��F�K��Z�Р�憻�[��*�u����fAv����Z��K^�{	��^�}d�v�R��E�`��tdk9*�K�䚟r���@R��.u�P(�"�_yu:��F�#�u��:�R;2�.�|��ZqT�Uq���$Q����V�ԇNwCS�׫A��z��I�K٧�Pu�Ṁj�c�hV7�Y�	�������A�����̇�z⵹�ޚހ�U�w�Q��c����U�x�i�Ge�2��}Q��i�G`�0;�'w���Ҁ�z�5��[x�T�k���T�1}ΠH�Kl�#�{"���L�o�7���#�C/
�a�ʏse�&d�>q�̩(�5R��ɔc.L���2���(�1�_0���І�����N��u�f�u+�E��9��:�2nȡ9n�;��L�h�|p�}��ji�E�̚w�gK���WQy$�aM������p.��u�{lZ�)�qy$�G;��O���}�����+-��g+�>��#�l�u!��ʓrF�K�sc49S����x�Y��f�ongR�|���Z�l��휔��^�Uª���n���qu�5���[��>��8�4��0]h$��J�u��s.wX�1�a�
Џ���@2�h�{ovPe[�i��n�*֕�Pn����c���aO�2�k�.��{_7����A��n�⋊�������c�!���<7'2/P:��N�f�]�дՅ$�^9�(�);[ޥֻ���L��7ep��ɹ�>��e�*�P�Zt�/�It�
�e�b[}0�m�N�'je��ZR|y����1-ߊ��Ov�4�hV��
)'WR�Wx�J�L�����뻕7U�<y!����4���#T��D{�ՙ��qb$غgP����!ŷ�K�Fr���ۄ!��q3���H&(�U�v��:�x�\Fz75�um�蝯� �fJ/%%%�Nܲ�̟����&�
4j�"�ׅԷ�s�裥Ղ7�=ۍ�Z,=Or�tYe��6*��9"������'sz
ʳ�U��e�ņ�ٗr��v qe�C0����A[[Ql�Y���$�o>��܋�#��Zp`��s(J��b�S7�+YI��$pec=j�\�3�E��lX�i��{AM��,:���o
�ll��� �X+w�+kT��T[�5�\;�n@��ې`�tF�<�yFxS](=�������qfg3H;��1Ri����\�����7p`բTW����5�hkk1��5�it��{��F*r�:Z�SY��_Ms�ʁՑ����g�,K��4�|/��w4�Ӑ��+��pcf]�fwS[�q&u݀�8���ժդ���~�O��R@�m�&��-j"ֶ�5T|�D4E͍�EQDm��`�IY��h�C9�I�(�����kAF�UU3�N�#m%1m���h�����͌�"*��j�L�U���((�խhѶ)т(��`�q6)&�������0M�Z���ITP�0m��Y�j,lSEi41��6q�*��(vp�QEATKTm�h�f���8�bF�N�*"�"��"�@b"����i`�F���
������b�F�f�������*#F �%��(创l�:tAZ�TFƊ*)��l�AMPR�m�����AT�(��
��")m��ZU6ɤ����f��.�'Y�����JMb-���Ѥ1��U%QIA����z��r�M�MXB��J� ԕ `������XE�#���9�w9��CS�����]X2��h`̅��-}��SÇk��?u�l��txo�G1�1e�W9}��v\���!|9�u]�����bg�8����{L���ج�p��[5猾|����11ų�����ã��2D�,nI��`��6�}�΁ �+k��jqۖ�5�y�w3ެ��ۣP̶�n�	�$�KA�Q�y~�E��ͷ����}��5�����d=%"6�k�v�a!��h�dN�Ml�q��[j��6v�[��KՊ�ܻO�n �UA�3 t����[`B��vPe�[N�>M��܌{�WsO�6Yȧ���!n$���nl|�z种�сwc����ZR�B듷r*i̊�@�ȬrD��ֻ�ia�Uj�T�!�$��
��F��N��}�>��ʭ�3�;�z|k��I���nۡ��z؈�o)Ғ��Rd�U��r�<ވ���8k�c;v�ȍ���ҷ���l�-7λb������򜂡s�~�[�G��%EB�H��b�|�U'fog'�gd53Z9�̈���\��h|&�mG��k��s���-��b��R��;;70&�h��[���/�TYeQIkV�����}3�� 9K�P0:�GYz���\U��T�,���=���7l�uz�����S5�0� �1&5l�Βq9��F�T��߮��]�
�]���׎7�n����»�)�l�lWv�յ�L5km���`�I1$�ɵ�XV�8T�7��7�8\dtΩ����2��o?�oSv�U�5��؎���(�n,O�/��J}��b9���..5�;K�^^t�`����It�[�V�[#�V�1�v�t����=�l=�rkm��,�gt�nS��gvb���c��&���<Fo6��FϻE�ı#�n��so�t���;1�J8.�<:��Ӱ�n���ǁX����.+7�K�L����hR��p6r����t?$�+$����˼�/g���f���b),� ��YK^\�6*T�3����7blp�X�~�Zᆮ�j���L��6�#�@�p�?d��xU����&���]�8����C��Ǎ4����������;��(G�F��wi�����:I�4��A���sNR�8��p�X�*R��DQ��R�6���:h���Ҡ��0b�N�9{��8Yi*��p6�~�D����/.j�ˑt��W��:����㺜h��[��_]*Jq*�\d�Ab(.�@'�Q��4�hl4#o���E�<2��ǜ�+EY"�~ե�ny����IU�N��X��ّo��Kc��g�����ñW�R���$ʕ�/���F0��w�����*l��#�t�}��!p���Q�ڧs�t��,V�a�@v��j����{��y�����f>��rרO�V�Y:o���c2�:�o;�+T�+��g>g�k��n�����k^����`�K�w��C&���3#��MrJ(%ܻ�|���������﮵n�|2��dA�ʍ97Uܒ�ޞ���6�p2��*7���������Gf{pңu{�uh�=�cg�����uWJ�lZ�d]�-'�s���m�'q�gIgh���IC,f�8j#�{J���Jf)[�oW��-��7�ZD"�4D�n�b4��q�+�����W��mԼn�c��w����ٴo֫��gwws;2p����PgE2t}�h�N�Dk�5{��������Kz\����c����lP[�ͯړΌj{��h*a�ݳ��~���7Xs�S慊��������w�fg���r�/Y��3X�GO>�cF�壏<��K��g@����.�h>i��nN���3|t�̲}�HI�Fi֎�-�`�?J��<���{d�՛�A9s����
�'��Q5u@fdZ(u��k�D��\+6��{t	x̀��x�;�ݝ6���df�5�����Q6�����)e�7ƅ�5@%�ѳ���-mut���fT���3��p,B�;�������+�r�t�Z���[�u���z��ۿ�Dt�����	��.D$+x_���P����6J�pc8{qD���'�x�>Z��u=�E�I�%p��q�F>���e�!��t"l7?�)�)2tL�����_�皱<��]��>�,�CxQ��ˇe��\�/[�wEB����<�\mK��VT�5�N�8�x:jtjR⾁JƬ�Si�{:W#���հӘui�4�$(]�1�qޑ:G�<)� ,��T�tI�nIYu�;�|#�ĕԚpWU�'e�szw����*��BÜ��%P�+�Թo>ϏOK��n���N���zÛfbx9���my�E����W��8�$Q��%� �:Y�iU�9�[Z�ws>�0B%�k�9�ޭ�I�9�]�D,�Rf��N1��V���J��t��@�a���s�S����J]DNѠ�3Xlp�u��d�ۈ�>�ƕ���-��-�7ͣ����V�\d�ܚ�Y;2�������J�K�2���>ލ��lѰ������ފ˒��h~�$�zµ=�T�����3w�5>& v
��ng���lՔ8ܺ�YY��w4h�Gt�K"��w�f[n�D� q-8)���I��u��l����y��q�?�(�,��S"6�����3	!D�%�.��6fVuɉ�7z�!W}<S��8����X}�F ;�����%����X�q�su��і^�:�+��g�u��"��H,�j�ᢝ���cH�uR���S:�l��;���͌���_/C���b�+׊�@����lSܣ���I9��z���͒�hm(��BdD���2�j��\��n�̬����Aj���OƟ^Z�k�p��,��8���+q'����޹S�;yú܌$�RUiJtk۹4�@�dזLZ*�u[�����:�o��Sc���wa�����J|�B����P�UW�n��L�k���-͗V]m�:��z���#�[;ǽ�) ]��h�Sup��˭��ݶƌ����懄Y�
lGp	�c��e�^�g��T��E<�l���/o'8wwd�
i���5�
t�,}[�s��8�� �حiٸǭ;3'�{�n��� I2'�F`v���w�7̈*��}�+D���n�t2���}����gûLH7^�4Ot�k�S�gCzo0[��jY��3(ok���<����OA�@o%�Q5
{����z��۞����9�*JT��
���w�χ(o)�c��]t7�w�'�AK#���?C��ɉ��Zh�ͦ���l��^���d1���\��Y��>=�`����;�}���w6�9���T%i�8�P�P@�����M�{6��n�n��X��w�W:M�]�]��1ռ�6�p���:�nX R�ܓR�ͱ�\�j�vՓZ�Is���v\��;wu��S/p\�j�|���m�؏W����n�v�u[���k�7fJ �P�"�3��Cפ	�#�xW:6q*�����#x�S��]�-�"&��M6��m�%k˭�g:��]�w�lF�<1c9�ӏ�ǅ3�r	�i,�nE������l:T�H��O�j&%�v�D���ͪ#�W�Ld�R����^	i��Y_��8�n��U.�'����+Όg�jv,��.2u�z�z�ۺ�=��\�N/K��~�u�79g3����++s��jk[�������ޅӝ�.��Bz�&��c]f�ͩ�)[�l�
b*�#q�Gb�mH��f�c6�L����(^�P�%�M*�⋂���t�y@B�:B<����ڤns����z�S�L�Q�q�n�WLN�ƀד>'��.�v��.���4�o��ݼ��F��2lk��Mky7�i�ܦ�u�r��E2���yAh;���}ӮAW��Z�.�݇��5��X� w��d6I�՚
�^P��Ok[�dE�pv��A�^c�(YցIov��"��P�{(��U0�czo
�5olr�ͻ���v�Y�i�ڳ5�3��E�<���2�ט���[+���>����T�ĕwU�l���۶%.��Cf�Wb�j6=0+�Q^J�z��x�.��ot��i���Fd�"N�MO;�|�o@{;�_�����I^�I���9�9��5&f��pvB����CWO�'=��;��+�՛�=�tO��3Sֵ�h��5AH�wӾd@~�hl��;kd���}%œ�B��밵I�{Z[/{}�\�Pc<)�sX�u[W<��=̩����<�穅���m��n�`��v4Nkr�π�#����/��x5iM:�Dm_5B����箜2i�����@�+=�YJS�u<�2�-��s�#�uћ��H��k�D��{3#֑]��x`J}�^�C�W67(�ծ�"��g���/���U��ET���H�NFjJ��4T��z ������8q/|?q�'VŐ�_��c�>��lF�K��\t��-n�+S��T���$��p��9�9��0X��G�G�S���?Q��X��u3x�H^[���glp;�gY�t�jxWsg-�ra[Ȗ�*���fd�y���Y.
�tcc�[Ko$��]o_���������X���VZ/�=��Y4�Ǔ�f�V���:�E������UG�:%�M3�B�-�+x\����ә�T�ѝ�����Ϩ�~O�"��l��N��"E�Ij���st�]K��ٕ��t)ab u��$�v�%�y\�����T�w/ķq��U�B�;9���pv�� �jU�>�����W�)���잞�*0xm��ד3�s�3����*C��`�Y��ؕQ��FRKu��"Ii�y���Z+8��J���l��N�dӽCfJ�6d�]W��&�{���vPi3�v��=rGR���y힦7?�ހ�\�.��]�TP�޻4ݔ7/;�*�|;���V���J���m�n��h�#z��L���X��GSG,�w���m�'{�H��x4��>��$`������t�m�L&&h+Y[�:r9��w]�т�ȵ�&_XPi�W'ŕջYy�0냫�7u�l�뢻|�e�%��[Ӆ��E���h�u��9�e6��tD�zw;H���驖29�&m��;H9����H�Vb��:��OM�t�a6���g;"k��;8p�5]F2S���6��$H���{��M9�d5m�m��*x�N��H�q��^M�6;�Fe�{7�HD� q�h����өQ�����_�u�	>����9�ԕ�ں�����P?N�����;4!��/9yܪ.�z�k˭�z�BMw�3 t�.+���-�fꫭ�x:�<�u�R���.ƛ�Q�[�],�V�<,$��F;]��LbhO]����X@���H��UB9'n榜ȥ�w2�z�/=���fލ���|�g��yB<Vh�;Kr
t�4O$��n�Y3\������5�3���7�Ʉc���[�Gt��t{����;��΃3Kt�l�n��m��X8"���'���u�ݎIʑW��~�|�o6��u;�|Gm���ly�8A�,�ղn��O=���z��������{���w��������^�W��NWM��e���<�^{F�e��m��+�����`��!m7��3�D-4v�twM=I��Ms��,ùDe+��a�ǭq��f;�6l8E�;VV�0�Қ4�u����'v}o�!���u�����j��̑�q�4�vIY-����Z�b謨D�;��Ld��T�Ηw�36c/�y�	�T��r�����ss��ᢊ�eX(��a=�P^���M������f�N�a�Ў�)T��,i�k��A����;�P윯�4�(&�F�}�6WwL(��&�y��.�6p��z��ɋ�&���ł�-ݮ}�"��vX������D=�.F��Kl�G�M�,4�KGA|�l��h˰���7s�l�o�1��Օɨ��k0Q��w�qRP��E����y��f�<��K���������t����u�d�X��o��B"���s!U�Ǻ�[Đa�����_t�ʖ�Da8�Jm�)��/ON���l�8Vv�%�Q*��i2��Β/L�^V�qs�؞^Τ�ͥ2�f�5����Ƹ�?h��pھo�l]Ί{�7x�֔�Hl͈3�SӸA�y�G�K� %;{�]�)o�r�Z۬tC��PJ������6S�H;��Ј�k�|�o��e����0��e��Jo}pÖJEu>��#{��.�aH�<��f�X������")�F�t�5�pj�l x���Μ�etYg��GK��ݼ�vM���m;�E�6��0Dg�%[��v���N�).�Hc�V�fڎW*R��;��2T�$E�/:�}wЉ|[]z��4��ټJ�,�/��:���d`,��U�9���;a軒8n�v���\��l`�dr+N� ��'�y���m�F�~t�D֏�xxP�s��o�t��Kҭ0L��`�[Ss�B
55����&�yt3�Bk2dط)R%���<Q�"]��٪��c4�����y�|n%Ikvi���d[׮�+<�\��.O~�M���V�����1�i�0�9f>厞N(�;�����-XṶY6-R��+�wrN��
�����R�Ξm=�K#��3�3��2��tXs5N��$ѧk�\�4ܖMcy�V��42s��j�ԛj`�qv��L�ҸC���{�ژ�qL����ԟWs�f�)K{k�0��0Х��v�D_m�4/&r��k9�9ו���h{�{���t*-{��'��/gg.t�hP�6�ʴ4��j�V�m�JD�6�Mٳ�8eL��^.���*T��m2�WU��S�m���\mŇ-�CF��엀�+5'��Cnvt�4��wG6����9�o�MP���T9jQS/�J�����8s��T���߲�,|\�ޢ��5n#KV5�UJ�Ӯq�4���ܔkl��B�XƦyH/&��"�v쉮�٬ukb:8.e%o�n���y<Ǹ�4TA5Al �I4�(֊N�����pA�PM$PKV�
h-�E�[`��-�E4QF�11���V�P�D��QLRPm��*��Ѣ�b��h*���klU1�������
"5�H֠�)�����(�4�LAE1h������*���&f*-�SLE-STUU&�KIAKMF��饪4b�)JR�j*
)�������J ���vuM��U��V���"�ib�!b*����⪦jH���&�`��&$�J
bӡ�"���)
�"*�b�����TPS�E4b��6�KMR�h�4�Mht��M-$T�"�$Z6�j$�����"(�`J����1EEUD[�4�}�}���.#q3A�*L�6�2#-�?��u����_a�����h��@��&�9V�bw��>�)�FDk��q�l�v����Ko��*���(GRL!JD�iBʀ�HR�C*���)��So��[��X�����Ww{�u��;����˓��kl0j�7��(�w��ћ����F.r��Olʕ��P%W�	�&�a[���0��C*Y4mN��;��V�ړ�:hl�R�3�cy#KI�S`̋�O�7�+8��m��Ԭ�və�|.�+`n`��4al�|9��8���-�V>�L[!�����Jg�g!(}��m�͵�;`�y���J���zMEE�Ͳ;{b��h6�@����:6q*���se��}�5���C1�Ü����8�@u��JF�?NC8A��
��E\����,\!z�3�:��N�IG�X���h�e)�rY�p
7��/m�)����}w��

숶Ԑ�}��M%�H�f��t�a��oXR]��]����=.�B�3W��T_���j!gy 4)�X֫ǳ+���Fx>�@2�zR���fU�����SMK}�ȜX4���Oz�zx`8��b7o3�3���v�-��_b��%4U���&�'Xb,�W�\�X^�ѯk�Q���8�5u���4���m�C�q�u^����(�Evl��إFbM�b�^�7x6t��c� �
� ��g���jP�)PHʋ�^nUޞ�Q�vui���V�j���r*a;��b��j>Kwb���TP��Ց�n��H����N��^�ࢩ�u��*S��f�34��V�7{y܍3��Oד �\zΆ�x�t���j/+^y�2�u��3���5���ׇ*\�Z�_3�T�w7G�_.�`�Ψ��޽�B�t��}�+�*;a���<��令.�,���P��|��-��4ݕz��G��^CQ��g�kjuTq����WrR�w��4�wj��p�}�}����-U0}��޷���J����luw��C(=�u�����W�����m��o�g����W�F�����T�w^�~�1;d7��>c��1�_O��x�Xc��=zg��3�w{=4�Y��XrVV�5�ƅJ�i��)	G%۱��6WX�����c2�i��AO#�
+�q6�v{�	��J[�}�<'}�b�ɳ�فe�.ޢm�I��'R�"����.K�ɺB\-'�sz�|�{�-qv�7�s�6�	w��p�������u�q���;'YfG��	��y��=L`d3�W��dLr�=��[��\��R~���f��S�.�@��$$F{N�r�T:. �P̝�Tn���O�ͧOcV��6"�(�ݤ�7632=|H���V��.BV^ɧS2�{__tveM��(�Q�,�1��ꧫ�6@ꌋ�jK;;����\�sd�ǝ��.��ݬ�X��3�����!@vr݀Z5��Bjn���J�pӸ�.=��}g$��;�ْM>zj��5A�y��ֽ�ȉ������	���7$������S�ܷSّ"Ϩ�Զ9c��ĩ��'��J4(l�m��G$N���#'o�T�e�ҁ��8�/*�V����
�4L7�l��W��rV�\F"���2��)E��`�np�-��0X[�����<뻬=]�U qtM.�z�2X�]Q�}�ݽ39m����̵5ŵ�Z�����qO:Yp��YX��ZL�y�.���w�p��
@��Uy$�jwcʌ�k\sr�Ǖ�ut]�28�W��g`�u�`��k�9��D)W+�q�p��p#*<�/������lǙ�R��H��4wT�6�w'���.��Y��p��j�͙-�Ɖ��*^���klɮ��j!��甒Ԧ�U�&����-���5�����ڢl[��+r"7Po;õMI�ޞ~��:uz�Q7j{V���n��m��ɮ/Y,�l�Zxt��6����ޥC�R4t�i�����a�F�"YLtJf�յ���Dm3r��Y���F`��\k��ō�;o�݄[D��Sv¸�����\�Pσ��<*5�x�p�n7�H���"�EkC���CV���8ךm�-3���O��kW~�m�//�7cل����н�u����V�x�q}�I�y6�ڑ�Oa��;�J��rb���k�g��f��ܰ�j��o.���)
�%��/-H4�F�?���,�".7f0)�����,ښ0�##9X$�b�^�%��ɩ���?/��dyv�V�!\=p��%%�\���{i�wYG4<	�5k�x�o��|H�I���S�W������x�*�,�8�یZ��P�Z#�1=�}ڗZF�'�s˱&c��|eZb��aWn�˾:e�NI�\�!L]v���o`]gka|�G�d�p�h
�y��|.�������!E/?V Gb��)��<�EUx>��8���g�oAj/���A�q\{��� ��b"��t$�u�ؤ�6g�9��a9}�`��MU�5ө�T�+hO��{���=�J�cR�w��,��P؏6�wh��n��u�M����,}[��A�S�B~÷ѝ�qۄ���׾��w;�b}Ǝ�H����f;[}]A���y-ir�om�7�Q{�5�Qɴh�ڡ�Q�W�$��6�M0q���7��5j�1e������p���FFL�C�L���ky.�Q5�Nȼ����l��J��i_g�!�a��#ss�i��=χ+��v��m���wu��
��]�"���g����nHܝ��؍���NE2�X��u{M=�춓Z[��݅ ��c􆡮��;��gVll�U�4���K)�n��\���c(nJ�;N�ܼ����2c�����]hȯOGHj�5�n�{Q1t�蹽����9�5n�AH_9�k=՜�]��}s�n�Wʃ-ݍt�&=��ъf
�.�A�Y�v�Mܧ�A����g��?y�F�1�Z=�(��?H�;�]�,O̷��'qȞ��U7�K�w\sy+�[ ��#b�ϲY�tY�n����ո���1�ij��S��ȹ�P�@�J�:ٴ��S�U����.�4wN6Y�9�C�
�`)�ₛF�\d�D,�AO�A�z��s�f"���)�rr�f%��UL��.�g��ѳ�
�8��R��*�d�M��ѝ�crg�n�ڭ�ճ�@.�O^El�p�]���X32�һ�Ttf�ۏu��U*H����]X����t�����k+n��~�~,�{nr��e$9q kɐO.��e���H!��w;�u�M!����v�S��F�<m���Y�X/���|�2\�?o�Y�1l�vt[fbx9"��)ٕ�:nz�b��[\��K�Wc�y�RǦ#d#%��lMg\�CT�y�5��v
g���V:gbd98Wf]R[�=��9��-��T%��'
]��:���]�����H�Z������j�չ����3yӜ���ˡL��=L���I9]OpI��/eǔ#w���Z|�:8������Tr���o�`F}���������{C�u^�J�ޘ0�shh&�z�����#�L���N��3P޷�1F�{gp�.Wg+��L4]�֪[ort��(d����p\ݔ�셽��{x|���M{�O�[��1>�VS-���-�>�c��h��n�Z%[�]oW��g�
lgo4q�S�M�Gp�sLp�n;ǟ�'�ɛ~Ŗ�>�0�k�;�yW4�c��������t�̲}�H���:�,��r8mP��n�#�p�3�/eAV�B�vK����Z$uve+B��������ۛ��Lwα9��q�
�XT�=T�z&�>=^��r9���pw=yD7�5�7���t�lv���Y�Wa�;�Yh��=M#Lؗ6�yt�M���}-��$�zMA�TfOM<	� z<���-fz�hj�ò�����������}; I�J���pf�GRݮ��-^9��բ~OM�n�C�5�c���)�',��8�ti�J;��W:�[�k��f�[Ab���7�ʓ�A����+�r�gJz���f{0#66��mI"Η$T�<i���n�̪��m���Ԕng'�A�����^2;�Q���JK���_�v&Z��Ú�6I�`T ~����������݆�O�-0��ԍ n+re�����Y�T� }�g�n��RY>~
���]�ɣ�Q��*���z��gD��m����@�;yJ���k�Y ?�k'߇��y~��'�n�ћ#��bg<Y�Җw)*�d���a��H͏0�`WS45�-t�m��<�(���#Ԫ�ӴhY#N��Ǻ���6���O�8�X�d:ޝA�+�]��{&��p�>q��7>�(�H�ˢq����oF�:�4E���x	�J����]�V�.��8��S9��'Ô�����"x���1��Dc��j�u0��A7Q���ԭԃ�'�f xTk&���ћ�{}�~��T���~��(o���3O���bvʗ[�����ld%a��~P���;FՋ{����ܵ�[q��Ⰾ�rv�9��ҙ�9����T���	�ulT�I�t����h������]ȍ�v8�&=�[�	�˸���=���٣V۵�r�N�⠳�����ю�G`�hu|؁��`=%"6���\cQ�-sX��s��i�c\��{���#O&�����"�p_��q�������0Vdm�e#��f�▝A+�]m���"���:s�b�N֮vk�Ý67:�O^t`�!�! wb�2 g��FM�5�mU�SNpф��ۻ]��C��dV�6�܀�XGb��rK�����R�wP�Bs�TRƽ��͚��MZD^�Q����'ׯ��eZ����Ͷh�͙9��\Ɠ�ʟo�5ӝ�8"�y�[Bx(�ee�hk"c���wGLJD�(t%y����-�-�5�� ���c�h�ަ8ύ4�Wm6�lT���{�/�'�Ո��:_����WG�X�}ޡ5V���=\f�l�
#b4�ٴ�L�.�x�����Lq����vb	�u3o"�$-si��P{� �6#�j@�*P�tF����O/ ��5ȸ��bidEDprno$N��&&�L��p.޿�㫠���%N���_&����nՇu���ħ��|��m9^yz���?Dvatb5ٙ��������i؅�����>]~(��
�2/�j�w�E���'A�;���?/W�8!(q�φ�ܑ�ԫ�V�>�7���k�I��j+on�y�Y��E]��CSh�󠎇�̀�7���b9n�}�hZC���[��il��1���}��^�g#��,��g�H�=eL�ך'F�CC�����Fz�����g����g;�+�����R�����k��V�vW�]��Ox�B}ȴVR��(�8vw�?��S t̥�w�j��=[�s�I	h�J�:���T�b��e<f�bg��	֑=^�~��ҿp���%��D+A+���)�:�vv�6�ȧ�7:�+��4�"�j����kgͨ�=;p�VڲD]e@�����c��_�����n�­�'"�G�����|��z=�#����{���w�����|�}^W�������^j8�U���q�W��;�+�+�8�}�ୌ��r������������w6Y t!�0��*R�8RѸ��M�3X4vd�z�A��+��xPU,���X�rP�br�D$E[�/)�]w])hx�N��>jT�]eu�7�Ӯ��nl�tp<q�D�_sM��tRz�v�rR�iJ{b�	i����^�	�a�u� �ڊ
��J� s�67�k2�"�&m���c�>�8�F^��`�����N���#�(zu���]��tu�xAu��ά̠�[��S��c��Mʒ��v��f�p|�AA�|���Fc��@6����h���G�ڽ�����s�5k{���v��k��a��$�z�ӫ��b만ܤ���i��Ggf���mXr��.���i��,��yX4�kT�F�� �$^�8_<L�tu�]�7}��)[tpI�a�9^��IdN��'����L��� �lR���쾊�vR�B����a�&]�F���z^�m�N6�!����g*dۄe�&��8�a�L���i�j._N�r�J�ܨM�g���,	I�0�=�����:��Q�qWZu]7S3/�ީc.A����I.���/�:�ưzs{��sv	�Y'M�m���wQ�o� \���Λ����,ܙ�L%�E�ٚr��qiN&��E��Z.`[q�nz
�O����Ka�Sr��gU6z6Ve�{��1�������M��Nmf����=��3��=�3]�I�x�Y���n�Da�PP�������%,��!�k���I�0��2�y�^����<��7�������3]3�G@
�f�3Fz�>���-[��K䛡Z�U6!e��yk(���UE�q0�<P�۪Я��{�1q2�RTo�����>Q��w���qT�N�Xr鉶��B#�0IFX�)@��ې�O;R�1а�ww%]��˱kl��J��E&@7z�lqc�7h^���ym�X'��3;=����(z��h�������YŢ''V!��&Lyk&K2 Lu(n�ۉ�VMmfXR�@�o#�����y�����$�D{+����X��]/D��{
L����z��0���e��m0b̀���P����.4$�j��78:0X������\Z��w�p��A�����y#*���j��f�PU��gZdn�R�A�� W����Zl	}N��%T�WS5�z,�ַpw���O���s3	k(_
6�n�r�|��S�Qˡ��궄B��<C�����*�ƻ����M;�^A�tr&�{�ۚ���|E�3�岰��])������p�)k����6�����V]����b��s���2c�8KO�����,ˢj��L��Er�/�M|��T'!�ԓ}pfcU�T�gsq��@[�S��uM��	{uS�����V�����H�C�)���
"H�[+MQ!KEPQJ]��Q�%EF�1U��(*�)
Z)
I����PTQPUD4��14�SAMD:AC����1%0�#I\Ơ�� �
��$"Z"�H�h��Zhh"��!�P�CDl%$(�����i���"6�4)ATD�a)���J�i�bhb(��Y�%�����LZh�kZ
"&���T�[i�
(��"�
����KY�!���
��h�&$6u3���3�QJ�D%!k:	���T�ӧLEAT�%:4�TUm�֛m-����l�&�@PA-R�!�^Hi�+HbZhR`����6��CT�)�����v3{����7���h}L���n@�J0Y�:fz���t�d�u3�.�C���L��蕣SvR���=j�k[HgJ�ɻÑM\6�ʺ����mxC���J�H�y�㮝O��.�6�
�Kf�!]�W=]m�"���R'��)+ˎ������� �}w���9�bgT�=��
|ס��i>�l�<er���0b�����>�}����ϴ��88Ñ�btTw�3�[5�(Ku����Qy�\�{�:��ֺ���C�3�;�W�&h� T�rS/��y�w�Pҝ�T��Ov����^`�l���}=��U5�����$��6�=<�k�����\���K��i�e�4c|�}��s�t��SUA�V�����
����a=LvW7��q=@�(1�g���_WK�^>�����3p�C>�\��$� R9G	�nSǞ����9�\3��w����Wc˕�U3���U�{�=�d<�x�!" �^����T2��N=l��Z�;?t�n��P�gXw�����+z6�k�Wx�gGN`���j����6�[�3���Ԭ&v��ʧd{�'A|ޣ�\�d�Q�&H{5m�`��!��P�a퐭��Cf�Y�"�>�^w@�G���	�,�3&��A�����Ԁ��3��D!F {�^7Օ���u�����};�/�a�8!��+��:��'pE]t����zZ�j���M��ȷk�ݏbD�����\8r�x��E*�]� ��Z
�� ��p�d7V���S��j8N]$ �

�.4zM:��{2zi�i� yp,�����n�������0Ƒ���ѩ.@�%Iǌ�|�#r�cy��5y#j뫸�oYɞ����P���,m��V��rT�������R컹�e�wk	j�n��2|�n��!��s���eP�/�J�2���1������ni�ݜ	�4�vc�==,1��_���O�tu���*�fE���~�a�K�X������&�/XH�\^5��0}��a����o_�d��e�54^;����+%E��4cb��U��ʖw)�[��t�|�Fl~����{��O��R4�{&b��L�5\+]$���9Z�v}�n"k�Z�<�b��i���u�.M&�m�S�U��+(.�ͩ�7�!��V����W�������;NoC(] ��K�t��v�z4��G2WR���Z\�]��ج<&�	�ZJ��J��V�KA'I�}[qª@i�i�`�6GJ=]�)8P��^�.9u��Ԭ*���=M��6��;�毝����gvz'Be�2�8J=p���'R$]9CL\�������F�k���8���p~���m��^�~�n`�����G4:�ݤS�Mé�ky{�n����}4(��nyڈ/���F�o�;�@̶�j��L3�{��O&﯁�͞8*5��}|΁�Y�-��ھ��N͗5-�Nn�ʞ������6D�O&�yjz)���w �+�6%B͘�����}w��f��/V�+lAR�Iu��W��[��k[EUU��ȵ#��y
�\/�"B�*�"=�B��� �J�G$�`����?f�Y��l�IO�};p�܇�#Vػ[�S��<�^�g͵JWn�hvD�N"����^�穌M3���Dd�Q�"oҒ�?�n,}�����w�p�읁��GWEٶ&֗���#�^��A�b�9����ו��u�H�f��q$�}�Zދo��(6)n���W�Yt�Tߐ`PҔ�tEx]^VGmN�
fs��}����{=#'[���G[.־���)��oS���Œ~�����{���)�u�i�@�U�M���*�ǥڬ�Q�n�w>gJ��mҖn����)���e��ڪZS��av]��sF�"��vUxOޓ���]�䉐�?HF{[}<��.-�4D�����E`�B�@���ͮ�9;�Q�xcIݓk��jɜ�C���\i�-�������3��L�~���]E_���*�k��y��%���V���"ȪO�����q����J���|6�s�mi��澕�����~��5��C>�@�7���!�7^��F��՝8t?)��,T�&����h��u�hwF`<+$����^\X�|Q�c}�Hي8G r�yĉX���X�g"��E���z�!f��m37t�u�YVos��!֕]7�{t]�9�IV��E�%^�9=���Є�|�����^���W����H���b�6�#&��zXۣ�u�����Y�<O[�)�.������v��I(�d��r��,J�z�^N��k~����}tnnd�28��&����h9Z2��z�ћ���\���r�ѓ��8󔾦e��1_E,U�~51�m��vnE�Hh�@��iPH�l��6���fT��Stj
��P�r��ظ�D+�PJ��f�gjӣ����k<�2}sNhPATP��</V�`�����|m��gyn������K�e�FUB铷r�u"��p���Ehjaw�Å�q'���f�	��b@��xM��{y?z�U*H��뎺u#K��6N�om	��ɔ��Og>��6ӇJ�9�ݲR��Ƶ�ρ<���3��r���73ѽ��뾙�@�
>ڔ6��M��d��4�X�<�_#k.��&�q�\I�c��F�JB���$-�#{b��s݈�Y��zu�CKCf(/|ls��w���Z׏[�p2��p͆�θ��zuT����`h�^9|�Bh|7����5�j|�݌�a[�3d��w���_���C7������$�n��,+,$E��i�X�O�}ݵt1�L��O���xt�a1��R{֦^�51�� � �翍�2:��pā��=tx��U� �.�N�h�Kd�n^�d���o�ʞ��w�T��_M�f�;-P�ڡw/m�wk�2��7k�<d��?��V��g`��!������.}ƨ��S{��;�n6՝��AS�v|q��eW9>&:A�3���k��mhv�E�Q�B�����pc[W)`w��#Lp���<w������dU�S2��u���@�g���/����Z7�s,��<�ѳ3�T��z�d���>�wձoӡ����h�j�fG�:���[e�e��-n�W���t7�Uё��OKX3A&��x��get�W�\��cD����Dv��8A�EJ����>=pD���*�X�OVi�hȓMy�;�_\H'0����W�;`� �d�[*������/��KL��&�}SPIyB1�@�"�ѥ$SĤ��9�7~}��ٷU�wT	^
&��csC�:�
�5�w� �� m�n�F�rI_<��*i��,�)�L<d�[`����T}���+*�1/�q�
c%�Eo���4��p�1��
��a����H	�o�z��<:�K�t����ʺ�u���=�LR�l�a��ĺ>��a_
�;><�H�=��iwz�J{��s~������+�\y��+0�l��+���=[��VzҤ@��L�6��S��������t�#�m���/��G�{��95%Bܷ�#�U�ҷ�}=�1�K�VK�]"@�3�2����AƝmv�~�v����X��IR]���B�7<}��l����h���i��j�k��}T�@n�T���gr��vM�C�^嚩Лw2�onO~`أ�,�d���W(Y�Vo�Wૡ=�jm��OӽN銹夦7=�/+��Bk0+.\���@�F�.��i��}��F��Z\��-t�TP��Z��|����f��ƀ�$JΘ�	����uf��n��l��r;l�W�0�@Ǩ{�d<w�>�b�ѲґiJ�ܓ����~�TqW��z����w�t���0lR�-ٓϔ�W�w^�ڵ��\#*m/;��|�Y�Fȑ��M�y}v��`���K`U�\��bvO�B��T�\������]**����ݥ�Hz*��M1\'�]�@��p4$�f�̧ʺ߻�Q����-�$����$Ev��+ͻ�'������[��W>�%$��mvr�X,�%�ϵvD0��X�/�9�Y;/'7�ޡ��'����Kl�
�,K���jE�9�3��g1sDe���9�Ċ{a�p���;HW@�J��*�.�S5V��sN��M6�h;�:ji�[X�nɶDj�6֖��G����t>S��D^��<Rx�Q�ɹ�c M3�YDfBP:؈�e�o"��v{)�rݘ�!�}'��㤪}���N�k8"�:+hO
���%�?D�c�b��E�B���$��H��t�������|�aN��S�4�Ԩ������*���{����ؑ�GU�*�4�9����ܜ�v��	�k����W�^G�����خ��[TJ0�h'vA��s��1�C6A�ۼz"Y�n�`T8[ӳ:��T���׷��P.ae�T��7���to#�����~�p�0!�+S�j�7Q�z݆��Z�#�U�l��+�W�p��Uϓ��û;@X�9c�H��O4�o��0����s�<ߩ��+�a�^]Z�)$�=��U���E����OU':�K�4m�/g-��-����g�&3�c$]�x�y��"����f�#M�S1���g6�ۢ���K�B��V�
�l��8�qS�����t���m���>ٜ���t�c,u�̭�Mg�;_4|9��y��w@�+��3볏�p������١[J�ﶛ'NN�^�`vZy�q#=Ŏ��h�dnzn:��t�F��>]Y���,�:�7`:H�M�+�m����K�	�"Ւ�N��v���_vX�=Ɲ��]*��\�a�Q/����ց��Қ���tNLͧW}��:��U��aM��L����6�f�Qq�5�����2_��������d�=j��˰5�
�:0 �E��P�B Ӫ�c���m���|���]��8r@�J���P�d��N�U��@.r*�=l���p��"y5�cY��!غCjF���*���~���Gd�����&���1vEf֌�"�p��!��ddns�t���q�������+ޡ��C&�v;���������u�=g�T^�T��Fb��sI��,S�Z;Zv�i[H�i埱o>Y���f�u~�F�:��)EZ7cU��,���i�v�E;w�;4�%]�jm#;
�v���F8:�N�d��
��į2��%1/�����vP��66�N�x�%Mq����^Cu������p��ݸ�}W*A��ao��r7������3~���ߞw��&��Ґ"Nn�r�w���2���@u�voժ�q�O��S,�g%8�$�Usm���� �3@҃T2v�?�x��#y�E�6a��iO�p��>���S9�:z
�c�x�O:rFX����J�-*��-["/c9��f����xn�N��[طN#��-��$��;fGPc=�-q����.�n6�;��i�c�{�ѯ\�J�p���3��#5���煙}3�{R^%4��}Bze���r@�}�ثF���!�����U�i�5��E�}�j��,��+�`S�����DZ������z�S�EC�S�Ӱ'�O"N�jL���[���j�ݺ���7��4�u$�&�]���/�{�� W�� ���?w�#��>No �!Y�fE�`Y�f�V`dYV`Y�fE�e�	�fQ�B�`Y�fQ�V`Y�fE�BE�V``Y�f�e�	�d%Y�f�`Y�fQ� �Veb`Y�f�e`Y�	�f�VdY�fE�VaY�fE�aY�d aY�fE�V`Y�fU�eYVdY�f�eY�f & &��fE�eY�fQ�Va`Y�|���"f &Q�dY�f�``�a��fQV:��^�T\222�2(0(0�:Ϝ8DAQAE�=C� d@` a n� 2��ʀȪ�*� %� ª�*�����0�2��ʪ�*�\�� e eUa�U�UV d�dY�a�eY�fE�`Y�fE� �V`^a��eY�f�@�`Y�f�V8`eY�f�eY�f��W�^c������
�H* ���;;�sz��׃�:��G��=X�w����9�������u���Aϝ�}�f ��γ�����xU|{eA�EA_��H��� dޟ�_G�'�C�>�C��@_��X�~A~�?��2K�����������D�����?`~��lW�����*,�"�*R �H! D���I K BH��ʪ�H 2 �*�!( B �  J���$*�� J0 �*�" A*�0�H ��%�a������'�Eh� ��A�?�~c��n�>���ߜ:����~ʠ�����)#�s��؊�<a���q��b�
 *�3�~t?b}����Or ����
����C����������p~��a  
� ��������_�y���`�����	�}�D�O��t@�����P�_�?PW��c�F0s� ��lCU���`v?�A�C�@_?�~C�g�� PW��������_G�N������?��={�=�	=~>@_	�gף�L��à?7�8����I���UA_�zO�Y��>�׳�
�+�?��~���}�!ŏ��d�Mf;�X��f�A@��̟\�n��BEJ�����U"�a+cJ������
Q%�UT��U����U0���@%��5[l�4ְ��JD�J�̶5i�����dm�5�l�6İ��LYV��)�l�5�+j��a-*M��nͣ����ٶ��(Ҧ�6�n������-L�+l��susl�&Ͷ�ikiMiSYl�ƪm��.�ukU�K3Se�kJ̶ U�k[T��m�V��jf�*ZhRٶ�m�U�l+%�X�Ҕ������ܳf���   �kۖ
6�mն��G^� z2��M�gv���iѮ��pꃛ�e�\�� ���ڲm��{+]�꡷H��-V )�ggQy�Q�r<Ƴj�kYIT�V[+cF۾   ��>ؑCB�
Ƈ�W����#lhhhP��n�hhP�B��С}�o�B���/��_v��� ��OgnU���z�W[-�m���%�z��Tn�;���F���'��©Km�lڻwZ�3;qӾ  ���Y2r�m��wil�Ճs�;j{���i���;�:6�{ww7��ڷU�Lsk*�Z/W{��.��o;u�ʴʖQ���J���ٳF�[[P�m�ؙ�I�� s����Ǯ����s�V��v�^�����K"��vj���sq�mOF��l���^�����=�8�{�.
�����{uQ��{�6��"���-�S%�Z��w� ޡ���{ڽ�#y�����4+����=T�M�f�K�]&L�T��uHWm:�j�wb��ҥ��wP�v������Mkbj�Ka5�w�  ���DGUn���W��{-�Q^�z���X��v޷��%���*��5�4H㺎�cͲ�X�Wz�m�"�WsZ�mcm�;�I�2��Zk|   �ǻ��ջ�U*��{c��*�.����G�;����k��AE�w�]�т�׳�  �]�@ w\ێ��(s��fj	(���ԙ��j�F�   7^  ]��  ��8�V�to]� P v�n  wgMX{�  .��� �;6� 5X ���84����-�cmlҵ���   �� ��=oA��n@4�w�w� ���h� ��� ݮ  �  �{� i�c���  �����6��Y�$��V��em�   �|�@ ܦ@�'{N = 8:��� ����  ��.@
!�  �� e5e���t^� P E?!1�J�A� �{FRR��  5OOL�T�Pi� "��	JT   5OȘʤ�!�4�R$̪�  M������������xx��sO��Ճ�a�AV�W�f�Ȳ����kp�鯾�諭���>�����Km�Ym�,��m���Km�Ym�|��%�����d�ږ[e��g߇���5�_�Utww��<%V��^�ժ��c��E	2S�n�ƞ�v4m��]葷gm�rbNJ�V)n� (Sh�bB��Kd,ǂ;0a�1����0w̑�X�a@^��!a��
�LwbI����!�1����'L�I�QMu.��ޚ�ð��r�WP�b,�l�����u6�ڙ)�ݙ�cF���Ęˡ��mb
�d��Z�B�+mi��}�
��b�ЛB�Ǵ/.��ѓn�,8c��u"��p��h�T�yk@�*bf�J�F�t��e6+Ưj&�вo�@�`}�6�,b(�$��3vZWvZ����h�j=���:k+"���@��T2C,�Qx�w+y+����
���p�P�d�Uݫ܄#1#�h��^�W�F"��G��d�@���Ĥ8�
�d��%�L���̉\z��Ѣ�54k6�B��C�s�P:��`���l�y��]kǄ��i��G^����S�W)<�[��W��XVj;�7�L{*�S�V�����"���50�,R���8����B<�ݔMm*R�F�j���˅�SrP�z]�:W� 5�m8��cd�^=X��#l	V~��S�+b�v3�K ��[$WJ��&Bp-�2����SY����]�����hF@&��&�GzN
�1^D�[(I�j�5����S�L�Z�������d�{%�5����ڴ>���R@M��uӵt�{*c��&��e(������H�k�Ni/]�E�����ܙ�{V�
�~�[zbr;�ډX���K�EM5�ؐ�u�iP���Y��)�-P[�fܗ����0�u�u��b3,�MJ�{)�%J�,�[ZIn�����i\kwmb6�I[y���t��(����������{t`&��Pm".�j֠�)�Y��cU�Wq�Z&��r�l°��A���&O�ۧ��T�%������X��ʊ�,��Yy=�j�[3t�P8i��dmq��)��#3
@�JZ�F(a�3�:h�l�MR��[�w#(X,��:r�x�e]+M�Kf���v�H���K�	�6ޯ��F�N�Į�rK��;{���S$W���A[� �M9��,P���r��)ږ��y 1N�ma���E��ۺ��@6�l�&![l���Kh�;"J�"f}I5��7[�Z�,�7^T�G0���T>���n�f[�{�R�/��06[���#h��i<��&��E*�,8JzU�$��aՋ���Kh8��L(�4�^K��E�`
m��bG�t�_�=8��3o�R��p�TYH�֖��Vm�4��6�iR�Ȭa��K�-J'@�E;��а��T�	�������Ҭ�Uh�O1XK*;4sNe �ʶ75L��ųgۡ�́�.��ȥ� f�0��C^���
��*�Nm7>�m ���F�c��K	>J�0�bmڠ+v�T�=z��+R$=Z�I*΍��U K!ɍYt�j�=U�kp�O
'Yi*Y�䨴�6`����ThZ��Y���F�E�L��G�ܰ�{�1��,bfh��v��`�8��2p3nB6ܗ��l��AR6);�%&��K�Y���6���P�	� Wc b�H��ܤu� `e-ڻ���"`�L	I+x6^=U��Gp���r�l��*8t^3�>hګXm�V�ndhY���J� ��������Өz�68� Ǥ��'.��5��r��$�o�*���AzUi�6VhsZ����l�؝Z!��h?�ze�r���n|�H��	�r���������S2�qS�XUm^���P����5L]��RݰkC�u���&(�7k%,� �ze�E;[�k^�!�4�W��*�
�DK*;g���?eVD�i��rXy2�=�FҬ�cA�j��0�{2�*ƷF�$���y�*���G�E�e`���V�р��GqGU���%��4�i��:�[��f�8��Ec�4�Mͫ����Yo&�t�L`��ۻ��N��Zʎ���-}x	�b����:���Ԧ�4� ʄ��hE�-���<�-�_��x�0-kBL���G$劵����G9�'���!LN�����CkH��"��WD^ȫ6��+���BU���Ʋx(�2b��1�7`U�s#X�$E�V�$֢�f6�*ZD����б�,�x��&���P�Gi�1��ө�Z�xց"%9���ط�9�ėm<W�d�z-�I
�������;�׷���RI�p�',3RJ{I,Y�<��Q�.7u4��;ƣ�W*�b��2�R��n�Z5��WZ-,�Jo����h��$�sN��G�~3�ĳEE{�ʔ�JE԰�כFܹ���H�����n��DS6¸9
�|&la��o)иil��D�bdoEj1�cXt b���إF��^eȣ()R&��B�v$�hLfe4ǖPբ��&���J"*��1�8��1V0�L�Dԑ���I�9����!���hI��-B�;�܅)[e�ʀ�v)E��.�MU�f��w*LS���QM{����.����^'9,�Ƕ��P�)V�^#�RaQ�%��D�M��7H�V��y�.H�ׇ&�WE�T2�^m�Z5�ۚ�7xq �kXw��كR�5�b�m8��kj�vf�9C"���9�`��)�e�p�%��=�ۆl+\,M/-��LIU�/p����Tj3����Z�:���ɢ�0��!GQ�V�r�9�e�B嚑=��X�m���Ͳ�ҳl���G4nm�j�͘н�*6��ދ�f��q��ѧj �V�@K]=̠nh�t���������)Z�j��P�/�bE�l��5xU��̥Mܲ�a74&�i-�Q0���A	�3j�X�ɩT`T�o�Ac��Z{���E��=GN�C7��$דj9V�ʙi��f�n�z�� ��v�je �ӋK��A1��4�cI��&�  �s�EeB#R�F�����$DV��X&�H���q킔�.�izi-;��6Pe��n�:]��m�w������k��i1%�d:D�&.�hl~v��Ld�������d{n�/��Y�+`N�/U�1�f��P��f�q�
�a'�xQ���iʻ�ϱ���m�dʂ��.��{F��2�'��i�Q��Gd7.l�f�%�V��uh˴�%-K^)FA��3v�#-�,��+ݹ�iz�«���{�Z��`+Wb�鵱R7J]KL��fi�$a�V0+�_E�N�4!Iӧ�H2��,�LĒ�䣅@�F&7"����cK���8��f�n�� ڻr��9R9�hWfe�땂R�����X%$��r��X��d�)X�I8�Wp��ז`f��+`��I�\tp��РܙVk^���Q쪛��TDI�bsUfH��21Mػ&��;t���SI���"����n����e	���Mk�pf�a���V�l!�Ӳ� �+/g�E��3�iT��f�O�l�M���:>������A
�	\[R�n'���x�33X��/v�m7����L�L�i������w($�<4#/�Li���Y406v��]��Z*}*�,)E� a��&VQ�1=UC*4%�y��ա7S�r�D�9�Z�8���dI�t�j����å<,������	�x,��P��=9�8�aBth�^M���a3��â@0e%O6+.l����������9� ��^�����{�*����Tr�5cV�v�K�tdDݺXe���U���ɷ���*�x��[n$[��D%��d���.�	��N��.��̓���7w�Uq��V^�V�n�տ6`���*��7vΰB��K�P��ꀥ�7~�G�t��A�m]X,%/]^<�>)�L$j���@p�ʷn�/h
�WX���&Tu�������ҒUrd���l!C�±���
I�i�B;�"��R̴J����V�e^���S��+TѤ�Y�2�3����b8f�6�T�fB��(L:U^^܁���i�b�Li]�y5�+)K
�F�4��K���T��yi�fŋT��d�����q"� ���mkX�P��/Q��������fk�-�ͳu�mֽ�n��ɴZY���܎���9X�v[u�t͙��ꊎa���9 Z�>٘
�h��+�YN�h,��*&�f^m�T7���EE���U���#vxlaL8�:!10(iea�lݠ	�uw�+V<{L\Q��^ަ�Q����ah�]���iU�ĕ��$�R�*���`õ{�� LO�cJ���Z �gei�4Tۻb�Y.Z$�� Ֆ���\�V��h��Vc�e�̭��RI��b�n57Fe�19�ha�M�ၿ���0<�vll�K1K���巬v*��{N:MS
Azx���
�2��V�WWfJ1?���O���e�^"���9��vq���P�.'WS��f��bb´3bu�z��7pVI+���t�.�W���֐H�뛮���b�Z�����=�f�����o��y)[>�ő�-B��!�5`[Z����f1 b���+1�6�r�����K^#cP�ij��Ƙ��C"��l W�eª�kY"��Y��+�.;����)�8*��$ԓ2t�4{I����.� ����
�Q'c+5��W���Jj�ϦeӭJ`16rý���P�T�`<.�����m��1�˩[����dxo`�}��j�k��C��[a���iP��V����p
Q�NnVSע�fF�A'7Y��������W�&��F�J�c%=X�Y�Fn��w� �X"ڔ�f+J�ܕc�N�M�e*w���[��pJ)�K���2c.<CdA��;�͹����l�X!�`2�<���Qep�l�C��Y��7R��z��YY���ʰ4�)�c�db,3eU���� a�-�Y5:YoJ� r� ��P�C6���Z�y�V���cj��!Ǻuձ«(Y9[Wgd8��i< �,��ahf����P���U�[QJd�.��,4@���e�ܹ�a��O�+qF�a��1�s��x�pnwvre���,���ee�kQ)IyQ�5�ڷ�ү1�B�I��˦��i�nY��v�T����m�f=�ہ&�V]!V�>Y9Kt��i��b�f���3VG ��f�Z��m��ckRmI���5U���K�X�i�V��MT�����u�]D_�Yl+OwjL�m�=�6�n濖��7�lfp��c���n춠��T��P�a걔s)ooi�v���d�Ӊ"X�0@`�W%�1A�FR�9�7�9X�,j,�vk���ޘ*�zp~O`���	W��X�UĠN}�ٻ�����Q��ɹy�����lX�e^�mA`ѡI�*��[�Mbxx�F=�{yg�=	3���t;Ʒi�����2Ճh(D�Z�@z���-6C�z]�s&�;R���� YA^�X6��[ �;�E�r�Z�YN��H�e�H�S5%L7r�ĄA��ȭ�(Q���,`�Q�`��K%�����ͳziժڇ@.�÷Q54E5S�J�uz�����6��,j�x9/�u]4n��k2�Z�Ajǀ���{sF��/e�G�ZM%4�L��݋2j�ڦ���{jU\S��Á�0�3ϣ��.�-��1F1^@d��&f�j7G]��B,������VрQif���eH��+�@�e͐�m��U�FS��Y{繏��ol^GX���ޚ��,VH��;T�ȣُ��vaŸO����^�JEA;;w���̺F�55�����\�0MZX���b4'�kUZPZ�pyyd�)�bJEm0q�jе(�6������+�"D+T,^R�Y2,��L1d��rX���<p�9JTy3Q�kA����nIYF��yt�N�:��F\L�(��e㹔�	k�v�a�m�n�b(ԂeeAxpËYV�eͩ��E�E�ثZ+Kן'B��x1����m-%��̕�},)��CxͰ&���̟d�Ԕ�ո���m)�F��6��6�'���wjMF$��Z&29#o6LݖN �(�H���r:�jC�w)�ݧj��U���)hJYg!���k�;j���/9n��f뻏4�J��-�L,��k/�[�M�����lK��p���e�K����ecԨ֌[N�V7�Њ�*�n�[�+�hR�md����"�"����Ǒ!��M�Q�2��AXu����C�7�ZP��B��%`Ħ;�(��#^m��B�0�����[�m�Ŗ�"�M��$wyN�R������U�"��t ,�k4�9��5��u�,����ُ]��f�%��Ѥ3fe�uCݥ8�Y�!�����n�n��E[wR�0�BQo6KF�]��(AG[Zw/1�М�����u	�1Z�z>0b��hN��K0G���JQw��M�su�� F�W���)�4˷X�X,V�<�=���$ur#�/u�f��ek�f�*܆��v��]e��B�c�G,LQ�ֆ��z&�m��c)/*�8�v���@"�+d���� 2n�F��#A��Ԕ&�,O/>Uѵt���8Kfb(��̳ZzH0K�w{.K���d7�M#FԠLؐ���YܘM��yJ�Uę�[��ܵ���N��7�)5hU�2ҭ�1�e�
���H-׳@���v��
̼1��h@V��R֦�X��YKM؛n��Y��"��3v!T�eA�C���jZ���}83�qos����{]�*�u�7�S*K�}K��2�Js��{�~�񚢽v(T�2�:���m3ӂ�y���F��/N+��eښ�kW;�&2�X�mY�[��=���=�Ӗ�_B�[��R�|z���Vhu�t�0�b����{�u���|B��C��Jol&�7��3�(3oC��u��,���#F�3��!������'gpUf�!��ng<Ո��UnMn��a@����Mk�=�����:��B�A�O�n:�Ȁ��%�;�z�n���S������[�� ��Obu>��K�	��.p�k�bJ�`�K�����������4�n�A3��^�Y���v)�EoU���4l���ũ��+�] !L��1��%h�_�\���"�\�(��mӾ�éѼ[{°���:�
���7�K9v�g-�i6��h�^��<x���u�R��l�y�mƔ�_��`��;|�o:nͽ�j�����\�
h���$�~-�����8G��Ζ���"�9�a]AmO�v���7 �7V�k��#8m��I�l>S+赍܊�ݘd�*�H�������Ï��zᰭ�K�V�Y��{�3��08��!�8c���MZ�OOB�8�ȭ�uc[�yx��r���<~�VۚdâM9���X��������z�۷j��|�nk�hCX'ɮSs��c���ޮqR����L�t5�\�Y� !й7J�,��o7&	\BﺉU {�9We��{��7G#Wz�z���	�8q�N�Q�7�9E��n0��N@1s�ҕm3���[�N	s,���t�73��ƶ���,��}7��:L[_z2G�x���\�U�`�7z���/���ٵ�z�;����\eC� �`������|z-w�U�?��ؚ/�a��C�����y�3�[�~�3px�5�\�J�}��oq#��4��;�qS�%�3��V�I�A�"�S"���Hq��R��l��m�G�<�6�\�m��N�u�R�>}st�7)�pT�p���u�I���V�ٵ�z�H��%���OR�u�2(�]u�;t��@�2���s�H�/FX=y�b��9���m�.����n���ÏW���2�g]W9�IRDŔ9��2�� T�����Q����?@��X�x���c�VDF��߮�;��@n�˱Ʌ�i��Y;(�KX��Ŵ����sɮ������;Y�_����E3sc'�(ug4>��ξ���w]��0����V;MP`V�;�H_�/�7���l�]��$���(c�8e�:��n�?whRef�
��i�W�_l����f����E��$����և��Q� 0�n���f(Xz����E��ܒ�OhA��u��������/m���q��i�\X�̌ޱ��u;Vq���[/8l\]�b���!�Ի�b�)�v�u��9Y����X_�����������A�ا�,`�I�y��N�/�Y��]�pk�[��u	P�h���	�lyQ����\^3�J:T{X��d�O����� ��v����b�����tA�:��/7�]��K�YL�{�t@��]��� �4�R���j�o�/�7A���(zx�;��X�]s��r��'ec�D�F9��ԏT(�W��A�2ە�ٮK���*�+��Z[��=s@E�]L�YyY�Fř��>P��Q'� �/I9&��*[�rh<YLV���u�����;���u�����������C�qC��0Ӝ�m$�&�2Z)�;x�����t;�b;�t�Vv�݂+��-�{�\�D�EN[��:��E��co���krZ}lm,�)���X�h�;}	�Mz�knv��;S�\�L8�-��+�׀b���;�+{�κյ�%ay����]�A�vjP�?v+��YQ���	|�fFȲ�M�u(�MI��Y"�2��le�R܏j�8�3-�3��)���..��{r���>0��R��6�e�M����J�u�-�.����p��C��T�]sڜx��9�Q�9C@����:��AeCSz���v5%�2�nA_C_;M���n��+ֽ�s�1YI�ҙy�U0f�+�f��j'/_�Ǜ��g<|�������,-���e��q	����%���hЩ�ϸJnă��0��{�q��1n<�{��#Bp��3�z�p������}��b5�j!]s7�e]jΒv���}I��c�o�.�����qa���-������x��a���)PaZ��ӯ)��`�5����7�v��A�Ҕ3{��kN�@	��C�4]�0����.�s��}�HvÂ:�в���-�x�Yv�r��bb�8XK�%�)�];�We��	�s;v�Gt�"��
i��b��r9����#�mi��;��"��[�����w��b�7�U�Ǟ�i鐃[~���4}c��I�V�w�FToi'6m��D�g{�w�ʫ=|��շU����7>��h�GWʱf��6���8۱HݨTV~鱰� �=���2µE�s�ר��Ļ/���h�:�N�9N�Ga}h�@�+��df��9or�h�}�RV�NkKO>GV3�z�GE\c�w3w{4�%K+ʎ�.�<8�����K����oM��N`��G���5`�pn�E�h�|+{N��91eѭ�A�
Y/�Wp�n�]��:�`���X2VV�[��ڟ�싖�`�$�YY��f�/�5��i�����tv�cX�8���77ڞ���L껨��Z��,�$[�3M��kFs߫cr���:�y�UϿ��ª��\PZ�ѳ��e(1G���U�I��g�ȗx9��s�#:=p�C��p�cV��V���t<.��D����m�9��$�E�o�Χ���8����hSl��������)���b��5�uӓ��q�(b_g|ɽ̬��n/L��~��^���ͧ�p���ǈ���r��-�K˺p�c�g�q��Y�.�1�y���[�og\����Rwk�˫s4��kffK]�`�Ny�EtwaI����y�ҧ�C�XP}O��[Y| ȹ�G�n��ff�ή1��;{�V]h��	O6\��Ņ��#�ִ�'��>;�f�o��pN(M��c(K=�����P���A2e���#��a��	����TJ��Ӏ%�=ywOR4�;���w2�
W��ZZHX��<���H�l��]�vLV�8F:�u��+��#�`9�����e>ۏ�!Zz1��k��֞�;��XN�^割
��^}�y�CJ��W5u��mT�2�X�ʻ�k�鬭����q`�*.N������"����Y%����w�����W��nz%^���v.*%ٹ��#�f�l�g����Y���w���:�F���l6r>L���܇�*&������EMņk��kP���g���h����j�m���uyґ�}�Â�̢X2�� [�ӱ�x�S�u˳��N^2�{�G����~ԟ���l�o/����^�����qhY��y���z`E�h��-w
��'l�O�˷y�&E���Ҿ��I����"��ݙh��{y,�>|�uQ�i�52vT���q������"����[��sj�Wk+L#�u"�ľ�4��9=���$J�6�>��V��7	�J�D�UԙJ�7��y��b�aT�ZԈ�.aSh=��� �ښ{v���_�|�1�R&9��Xr�w�Θ�k�]Y����E=G#�zQ�T}�mlc���y�2��z�o�)�$�NE���'C�:U��-)�&[X2p�GI�۽�z��4�m�V�t���2������j�kT�Y��9�ЯR���)鲙���圾�F*��0���ս�����%|��ĥMC��ҏM�ݳ`��|�>)��Z��wTдM���o������N��E�xv�N0"�=B��z*.���#w�T�'s=�b��%��絸c^+�H{�MK�<o��y7�s.򊩗�% ��WV�g,�qr�>�Ͻ���A�C3��օ�ݣ��$� N)�!��c�:����ŷ�^]�x{&�|�x�UQg
�Vṝ�2�W9��<�e�!Xn���-�-�z\�~�CT{_E>�^2��L�����u��'N)��òdi�~��M�Xh^�/�Vqv�'4�!������6�K��X���q�6Z�t37dq�cmXTUě���Ê�y{�=Y�}K��7 )�T�%g��<ʫ��1��e5��h��L��Kt:�d���D.M�ٴ�C�+�v9�+�ܼ<�#��f�Ω��r��)�k�������S���{���w��r�b�K8���*r��ZzSxv���mL�u�m�^�����V]�d��������תּL;��_�������Cۛ��ܰ��g���x�^��=���=���j�D�T����9=u���i��\`�dĆ�JYٹ��u�"<��&�RS�n�[�-h�FNW���7�1���}��S�3K}�y:�
ָ:��t8���ٰ��u��A��
λ6�����q�mT�:���:DơN��g:󁅴L����v73 d�h\7��g5sW m��O:�����r��rb9�Ut3���ݾ�&Os��s$��/@7�p������JGW]X����,����	Ԟ=��0�d�|P�B�y�F$�хV��7�L-4�p2s�Y���;[��4̽I�W���n�t�~z�/j��f��F-�}���d��DpƲ"�z��wVYuz��0E�:LC�aq�pω̸��`�-=�	���:�����4��C{���t�.#lg��鄁���{pc[8ѬB�"��C4���������d<qꡋo=�E�ݸ������I��WX�څp�fgR��|\��U��e҅�b��K�.�P� `1�|�]ۋ5�Y��:V:�m��b��ՄV�a��ٌ�yDuYPhԤ��OA��#��Re@���S�A |]��;K�k�S��}P�R��Lv^;!�u��s�B:Y�z�`r}���m�y�U��ټ��+�m�<:ZX�ϟm�Qk�{��
����6-�Dd0�j�z��딍 CdCI�|�����[S>+kc��ة��� s��昮��` 7)�����,6��X;iޕ3���TAuw�.k�m4v�E W��9��=��a�����5+�A�y�O�n59Q3�[������x�^�me= �/4X�Qr�o��ʳC�=Oq�ፆ��h4��D��Ѿ쾇9nЃys�aԷ��v��V��6�I}����ۗ\�s��M%�۽��Ԅh�8`�#u�3��&��t����i6��٪K�7�.u<�ʊ���q��!B��T�9:EG�z_I�F�~p��yŮ�' Q��P"�q��c��׳�=�]WZo�؞u�]0�Iܢ�w��r�U>�U�6��:�n��t�*E���t��W>�uk�{M�z�
'�&m�7N���[���o�soq�;�"���;�ʛ��Z�0P���j�IS�k���㍋�Z�����j�w�M!S�1-��J���Ѯ���ך�F��^��0]s�d:MD��h{��H"��4�fPF�&����a��$:	}��������$�X�3�m��,�os���d�SpeY6�(�p�5"�)�GI�ʫ��<��M�e�Lg�2�҉~G6Z��wt;�M�j|�T�@��Z��D.1�lL�`#[5�]�KnL�{��S��o��qY�.'"�P�b��FU�s�|o^�D�t�P֐3�Ž��}GF��t�U�̇���>9Lӻ1��r�uz�M��Q�t~wC�eh��%i��+=�Z;��`�ד��&�e�}.P�:L�;}{��g��6�����ӽ��r���^^6��3��d-�.Cf�>�n��!�rS{��6��S�u��'�U�b(�B�Q3�>���������8{Ɗ�ީl��VM<ɚ�3���&�C�����Nּ��[3ȓ�k��]D׺MC2����^KNi�uQ̛��ۙt"CYbXn?t>�g*��%�!MRa4���P�hJd�cX�`룂���{�З��>��F.��+*��m�/$nkUӯߞ]������ͫ9Y u	��Y���w��y'ɻ4�沬��u�Æ����o4������5,�Yz�K�L˲U�+����G��x����w˸��� L��Y\ȭb��]������xL-��YS��n:*�;ي��n�z�@�N��VwȾ��||�i�)�� xO����w�M�Kv�G�;xe�|k�X��â����K����f+�I�e-�K�}FbsKt�D�ίc�
���z&�YS�����<G�{�\�[^�(N�Qxy^+V˭Ә�^��� ��Fh��#�T��垒�ay����Ma��f2�]�����8ʅ��n2s��DI�5�[�pw��`�}^@A�}�M[��E�,��k�-H�-]��e2R�0�0̴��S���h�Y026h�x�ٴ�ͧdX
��k�X@�����5�hs��<��Ez��<�[����Z딄��]�^zz��:�('�9妇�ۥ2*�y�j��G��~�ͧ��BZι�U�H�!h�桾���n�J������:]uvN�g��l����ܪ:Z�Q��:�i���Sn�J�I@A���خ�It��Wt���GV�t� \���]��/�����U<^J��x�v�o���'ҩ�-�-
�W<�G_a�o��2�	z��].�X73O�x�oޓ�%�Z�~�.�-��;J�t�|����?����|>����}�����xV��]K#G���`��n]~_3h�:<�����ܛdm�R��p���֑������l+�����\�sza��Z�+1�=�>ҟT<�<<C*6��k�Ւs0��������'�s���a)���a���M�����.����a�ii�ԎB0�[��1���o�捫�\#U�
����֚٘�j�"�������;��GA��TC���z0nķ;zK^>� �V񆃺�(�%^_�MB���$��\��� J�I��sK۞h`��3|tp�;�4:Av�ړˮVs�o��=���6g�h��͂���WN�h�)�b��aVd�N6����զA*�+�ܬ�]
����l.�.���u�`וׂۍa�Jܽ�r�b���P�X/�O��T;�@L�V
j��Y��_1�	OE��xD�vdk�7q���Uoh1��Y���fr�*gA��I�kC��V'�'[�wy���{����KO��b�
=B��H�]V��_`�,�I=L+�+�XD{2�}|0� ��t�����U�A�^���`^t������oE o7��a;��er�]�ܬ+쓻���w���Q%��9��C�ѧ���K��c6��
��V�1���ur�mb��h���ddR�Rea�C�ۅk�Y���)-���v�>=�����������>�ԫ�V�5���%@r��N�s��f�ky��J��u}��;)���St�X�>=�J:#�R��m�����
�����ή<�j����Ttq�u���^emFrA�ֵB.v?�H[v�i���Z���һ[/�C*�uj�xL�PVв>F�̗�dYΥ������I��[��jH���,7��!��ˣ�C)jK�fd��^�Ȱ#=Jb�(��y�]��qϜ�X��{УC��@J&�o9`W*
���͢��~���S7slKS��<2
�6v�-�;O�7X	�5�ۜ�`@�9��D*V�B��B�_#��;|�V:�r��M���y
�^����D��:�Dֆt>��l�t�R'�o��2��dỾ�]B+�c����S,i�ݧ4%իl(Ue�G�J�eѦ�ƍ| �x�={r�{Đǡ�No�����xs�Q�oۦ�:z�
x��G���<:�7�{�TY}3ڮp���<}=k��A�%Kӣ�O]���=}rدc���J��.��mV�ά���
����y��0>{�H���|�ueR�=Q�]�/c��yX�r�s	�Qe��+x�B���;�X7�U��M(o�6����zmy���m�{�� ����v�N�Own "�G�3[E��T�n���|)�@q����*G|3��h�eké[:��ӣoD�]��nS#LW�qoo�]��9��gM�����c>�r=��4[:e�uԴ��pr9ǄK�����𰎏���ۘ�b(�*�P��|N�m�w�]�{�Vt���$�����<Uj�k���)��a�p���܋;���tz�T�o�%����wl:wL����L�XP����M���2���Tm���V�ٖJ]���6�mP���=gU�v�!�v�X]Y��5Ƒv���j���<�\ӥ�W��F�0q��+�e
_:z�ٌ��C�3�p����!���׆�tX���
��b^,�]�ӛYk��o��N��h�'��U<�;��f���w�:�.)��3A�F��f%�.%Ft��N���-X�ܺ�
�ʄE��<�n%���O\���;�|��\��h��:N�yQ�hC�e>=�-��zl���� $���v����ԺX�;��0��DfXU1�9a�����g��@��9��#]�hY&q[`ԝ2P��7��:��;���Q�I�Զ��Z��ܾ� �r��	*j�}��'}�eD���k�h�\o��|Ev��j�̒��Ōf1J��ϲ�V.�$,/r��
������Ҥyz6�t7n{�J���!�����J$˲Mg;�b�Y۸�W�J�+��� CK���sk(�v����<�0��$1^egZ/Ow��!�Ég�o��^���ٹqԦ���d��*��wK+3)�	S����i�ƚKF;"�3(f�8a�z�:���%���	���	��(3,����c�+ی"��l�CiA��2R;���e�_[���ـ3�So����q�:7��#r���?c�7�s]�e���:����l��s�W��d�Υrx1�uh�r�ы�ڍ ��P�^�+0J��;��5�S5���K0S�|!�W�E��ܜ&-s����B��r%��]�-�z��<75'#6��*
^��g~�|��GX��;_.�ȱv�7�l���W�U��|�P�zZ��0�E�;)�o����3�7Eπ�_pS�\�X	,R���9��nwl���s2���H�2gl
UMniU�*�X���]�ږ�Th�F=������Da�g�[�5��8�TQ��p�_#5�WW��n�v�I}���;p�$h�쭀:96Tѓ���a�v��O�.<֎�t��cM.�c�U����5���5̭�J�)�=е�}��q��nO& M����v	b�=���-���o?����z�Lj��U���}]X�EۅϮs�0�Du�k���g���W�c�a-�H��x�9����)�_o1�w�����p���(8[��S�w�:�s�n!�(AӉZ��w-LݥT���M�0qϛcP���6�� -]Vyt/#�Ρ���3���微��$��XZxuQ
=�ŜF�ԝe�0�<�Qh'u8�x��D�ǚ%ʁPF/(<Nd�ý�i��R�����N6�&6�)�[a�6�z6,�p�5,��Ыs7�Pw�st�L�Un�^�=2�6�+�#�Qahn��|�ݖq�vd%C�nZ�Ӗ-j(��^��i����̽ۻ}��i��	���$8�f��X��ugQ,���i ��yc�͹���흒G��L�eƕc�bZK�쩇��o�6Ւ�^��pu*�G��P����M�u��: � o}���[�L�� Š_P��T�a�z�f��L�'�c��|Vm��[5��Mc�u(�h��<�u���X~>��+�rc�ƚ�4�M�{b�6-Y}r�
��@��˖�hcm���[��N��u<��4&9l��烋)}�6ɮr2�6�[����"1["�2��:�-$D72��t��mrd^���qv���{Z���X:�@س)��7�r�[}��w`=�+x4xt=o�K���,���*L�t�*4t)g��+�Y�y[��v!U#�c����n��;�c���X����X��pڎ�91弒\i��M���e��Ttn���FFu�u��l�1��k4n#\�K*��1[�z�5�C�9yL��lb݀S ����LkH��\x�P�T���6/��;�{q�������ں���FfP9�C��䧛�,��d:J��ju������|�m5�^O3��u��]�A�}��&���V^�Κ���:?r˶Dʃ]K쎊&?vkٝ��e��u�9i�����W`J��&{���&��r�'�})�4HeP���n�Ф���Cg5��'I�$�Q=�h��C��c8���bwrc�YC{�g���2Os�pb��ܣ��㛜�
ಳ �nY�u�!in��Y��u�"Z\�4;����!]ebi�����/F�.prc���J�m��=�ˢ���R-��m�
��,�\͸4�S�cC�rV��3[�h�L�c�u���{Jvs�qɂ���=���`Z��=Z�U���Dݨy
h��٨��0<9��i{2<B�G̅5�����/)Z�+p�d-�����bV`r�l�27�N���|�z�Y�AJ
�ܹ]Ʋ����@�@5b��T�9Zǳ9K]B�s����H�qU�/d]�àJ�R�R�mVr��v�i�x@�]MS��&Y��S��'J��g]r�!sGh������̬���N	�oi�g*]W�`pt�6
 �"�ݝ�{���.�����l���\$��Ў�M!�8;}o59ΗI��� HJS7	����͎�׹x�Y���AT�����-�Qjp:ugfD-(9�B�PF���|�^�

����6�`�p���?mݜ]�p���6ntDVME��k�P�"�ƪn	����h���w7vڏ����#*!e��R#����^������H��l����z���!spn,^�'kNt%�Ӗ�"#a���;���v38��`�T��ty�x2�.�Z��0v�{�f��h�����Ћ.{�
�=�8K��i�[[[is�%�1�7V�
�X��^m�J�9%gs��Lv�Iw|xc!���y���ϓ\���\�2�v�t���ۣ;k콈��h�u�"1O�.�G���k��7\1�Wb��'OY�l�Ul�^�W����3��K�q5�V���(�8���b�oV���� s���R�jB�eB뛴�7�y�]��+v)�A�?dL^�<#�E�::֧���c��JAf0l�;���ٌ�V{Yֈ��1H�%����3�۷��흛�G׍���T��%�
�is��ub�u+Ǒ��SyP��}Ԇ���	���pes�e�2��7Ѻ,�<�5���,���^���N�N�n�҇h����C*q��K�����lx8@n�
#x���޺���N�}��3U�ˠ������ySWB�/9��m���\I]ĸV�x�p�(Ι�(�bP�����~9�ɓu����QFҵ�r��;cK
	�+2:�Nft*���tdݢ���19-ew\���[l�j�E���n���mnW`e��Œ��¢1V@��O2��<���n��׮s^:���2�v�]��:��6q�v69���f��n��<^�M�7��Bi2)ga�N���.�a�ovo:�v��T�5��a
v�խ��z]���F)-� ԕ�mLú�1��&�N�ǹ0Y�1�/��X2TB��x��Ԫ�_#Us�^����\��rl��j�o���od0��;>��&�򾕻e�7�Ld��X7��M���B܎�CΔ��#s���f5$�����[�݂�tuݲqӛ�x����m�9�t�|aۯ����:-e�f����{��I�NMk�������o��|���12�4�	�K�pGs�g���z���GzG�/]��{ωK�W��i�G^j�V��F�R8+,�\,�7~�5�k��	��Nc�r�r̎w[[l�-�0�.����4�|S�+��6�g�ݍ�Ӆ��Y����(q�>�jl)�н�z���H�Bdɥ�sD��U�$��H�6�a��6��7�^\&0��29E���MOX�cΣ{x�}�H8SI�[��l$�d]�
�7)�Ok��A�G��4D���/`��C�;语�#�o껔Y��xVl�>_-�.�U���w��<�p.4(��Wݒ�Ƨ�78���;���ޜX�a�2�.���x�]�3���ٙ�=�Qzx�.�M��,��^n��!q��h�,�o+�Dq�.*)q��j9��i�b|�o�]J�vio0���oS����g�k�(N95�3$*�)1�d\75+��fu��γ��W�)���SC�뎹ݻ���w\o̶+��j�K`�sQI޹6�NMݐ����T:�cx��j�[c0����*�s��s�ľ85�Nx&1T�܃�G���^��X����V�|w�iށ����!��Pؕt�h�F��"YY����m^U���m�sw�X�jB:q�^�;��r{��A�.IV�U���h�X�ÐiƩ]���s��9�9-����֓��y�{��w=;�-v�t�l�ҲԶ8���d�ǲP�-��@��|xh��{3�2���m�+���K��`�q�^A��vz�s�R�����ءk�5 ޓuj��ZJU���P,����n&p0R�yY�ݣh��8��{_#Y��[�.q�68g���9��VA��}��|
�s���.��.������7�Xd�u��[��E�B^֜��
��єN'�F�F���o��l^`ٻ��n����}���u^�K:Ģr�D�dX��=ۥl.y�Ņ��@�ob�"G�&��b̫�h`*&��@־�ٹR��Yc��P�ee�94@�a�x��칚ݾʲ3p�\�*� �iK��D��(�B!	�9�X.:YG��BK�-A�Y�`��C���V�9�5%�
����f^��]&iϝ��;�xغ�1Ƃ��1G����w-��|����(T��s�]��t�Xw�N������p�n<h��7�"�.ԽyE4�K\7�級|��]��7 �`ζ�Vh1M�\�������E�䮶ԮZ 2��ʏ^e�Q�4w%�{e�6P��C+3���������整��a(N]���u�{Yv�Ym8��l�sVB|���u�\�j��C�{P�WC�6��"���6���@��J��I!�z�߹w	^�h��o�nJǅ${	�;��('��ܢ;���H�et�@����I����j��7�l���E�|ĩE`��^�cb(޺� ��v���ݹ�A�2;tڡvnt"��7��:�[>>�ub��J��A�W�HD�@��Zp���t��_;A㶠�j��>�Ѕ�ǉy=.��m0xv޼䗫;q�" i��.�4� 5�rmZ�i�,��6<:mS���sL@�$�Q<.Ұr+|I�|P�}�Do���ks[P�]Wv��y����(��5�k�>xOYB�rɆ�	X�8�ws�[��.����+:!ގݥA_���}��|>����cuϫ�D�;��J��������yƝ%A�-�͹O������=UA��[�{q��<5�un� �lv��GN�n�:��U�s���!�Ȏ��pN�U���x�kc����2����n����>+�ΡB���}w���~�z�[Y$��5�aA�{\1�=}�T���Xn�,�=��:��(;r|_e����P��]�a���T�jMj#�km.'s��;����d����N\6��h����m(��s�ƅ[ޟ\n�6�Yc+K��pEK�z����c�p����T�͸�N�m��7W����Tۣ��j���.3LɜKE3R�B�ʑ��� ݑ;��Wtv�s�nv^��;�Ada���!�2h7��W����~�cb�nN�e(Rۚ��T���\����۶%� ����pܩ�������юh�.��I�z{f���d�9��Q�����@�֯lf��U��9C���˭dC'e��n�[t�Tu��i��g�݊����s��;r�-<���g�r�D�7A;B� �!Ӌ�乼��]:�VqI���o�=/�uf��7�Kb�7:R�S�l��uؠ�nd�����(Tшs/M���N1����ʟ ��A�o�=9��&�tp��DXE����#U��"]�{^�~Ζ�SU0{��]�k����=��Ã�m�y�`�B �$|L$*m���i�D�C2�"!��X���I�$R EER�!$X��
T�\���23�"���!�"m4�Z��"��D""R+i��l��̻h���#k��M�B�D���"��-���D!h��T,�M�ń*$U��H�%�!JUY�*����ɠ�����H�H�ڙ�"n��K͈����9��$U��8��H��vҨ�)b���N9H\�H��R@�P��H��BEU"�6�R#��i�d�Q2b%f�!3G4��1��RE"M���8����@@X�mB"D�i	@��X��"�d�!K$���2T�DFh������DYQBx�DYH#�T(�����yAn�&�����v�N��v�ɹ6ML6'I��1�8��.�{S٧���%��(��ɓ-��vWXQv��R�����Y_߇I@�~߽�^������M	�zV����L���jb���6,�&Z�����q�(z��}���T݅�mA�����z�J��p�<�c�7óׯ���6���nP���Hm��yf��Y�W
єbᲅ����-j�'5(�oT��Y0�X߼�����_�	T&���=�k�	����c�M!�fQ���d̩���U��]�z�ғ8�gT'���������l]�_��G�h{�̺���'0��E��E�=��roJ7*
�N'f5��Vk�/��w�n_�Է����&W��Ov���'q�����s�W�$��C\��d�������F�y\�v�K�>��������xB�=��$r�V-�>��"�N����W��@�7zWh�y�^�6����h�v��>Lw�n����������V$(}ɔ��S&��k��p�^AW����+��N���y���57��9ъr�_3�3��D�=(�[DTO ���^�r��)]0��E�B<9'n��&��U��go�.��7-�w:R5gu�w�yB�ˊ�f��X"��%�0��K�ݘ\�@�h����1�#���P���S�E��k��+��Tݎ	}��:� T�U ӦrK7�/�(�LX�Q�U.l.e
���|�UW��)�BG���]'x����C!�I�pD�l�~D��tlexId�\�����yx�9���Y�֑c�:pT��xE�L�%�%�6xW/ j/�ג��L�ӂ|o��|��
��ׅ�3p����p����1JiF<8�ީ�;��,д���>���DC���Յ��Sۖ��6��9��v5C�݉J��ΖMg]�b�<�i-��)�e�OD<M|��*����Qph��z�MV�O���w��5�^�ˮ���U/����أ~��*^�Y=0���$��U��kE:skl���w�.����n���8W@v��O�3U�~�ܻ���%`zSo���q��m��4ƿpU
K����~�]Z�;���JԆ��3�V|a�S|;�r�A��e�z��������[�xA��'=q�^ݤ���+1�&�b�^ﳼ�7�,C��E�VI}�J���K�rq�B��8F�/lm=�T�}�8Кt��*��=��T��%�'H ����Z���$b/=�j���AZ-!q�����%)�=ؽ��ȉ�w�f�I�ܵ��g�lļ]M�Jz��a�Sl����i<��������]�(��a�OU����_h����կ�K��3���Y}LGg^��PK4v2�c}�}�av����\�t���:��y�,�P��Ѽ��N����=>�c�>�V�?��:s�U<Vm��˶�/�֥~�NC����]Z�*A��{�ґ�4���0}��<�FT��'"M"ty�KF���[��HuU�{��j=YE!9�����p����pr�N�����\���ź�λ��,��"=l�tg�vY*�W]�{��^�B��.�N2���BZۑ�Nϕd_Y�8�?�p�*e�m_h='V�%��\M�#am	��G�
xOL�eE�~��A:�.���b��cޕ^�t����A�4p�����ʄ�Z�$:'���xc��^'���,���;�8f�U[�h�f�0�RJ��.�O�H�u�Ɛ����φ.�����8�Wը���Mw�7�s�N�ڒ��V�爛�|%a
�RO���m	�qq+��Ӳ����wD���7�"�o;�O�4�X��-zJD&/D�5�Xjq!�[�1�^��]˝db�׳z��_4g�ź���z�ʣ�����*^�g������IX���9xi�{Cm��`��P�����jfr��I��%il'�,9w��	������],%7��{�^����G�z�����wKE��y�֗�(���k}�⥙��;���k���V�V��z��1p�������W&��B8v�ђ�<m���]���R_?X�i��ubR�~�.������A�UbJ��c�a���G���网����� @?Zʐ�x��~�b@�κ�O��|r�P���s�f+�7���!��%����]����@Y��ʘ��>���>=�����^]#��Ż}p��[^7ϴ��5��t�@0������ds�h�0Ei@��Q�ٹ�S:��[�kM�wh����;�7�������Kmk�#�������_��})`@u��yy~0���I)*ϫ^�Ϯ���ԡ-�v�"�S��-����3d�hp��Y��;�ν�V��%'=wg(x�g�T�ǽ�U��R�&�l�|$�T�3�U�����3��v��;<׸t��g.�P H���*���)��c,}��삶�������J%�w�^�U]�#����7�ĭi��E�$�_r�Si�������_Z��#xj�DہV�Dm{�>x�n1�*���6�e��_u@4N� -��ɠ]E����՜�$�f��=��'��)!�O�)<�Dz��h%aËq�p�{[��qm�vׂ��7bSzc�,T��sq�hti��S�E��&Nmu���V��QXź�R���Lq���粛�.d�N'����M������ԯ�]ފ^'yy�ځ�{VIH����r*j��Gyv
��n�' 1�O��cCuv��p�����!�"����'.D!^�m`�C�$�[*����&��|��o�P�T�L��m����E��j�ߋ�g���_N�,���GO�+�S��vEYC��&\]�1u8dG}�J�g�n ��K/�����6;��U��Ja�	����%�V
����:�=�,�XDSZ���j����O�u`��߾���z;��lܮ�<����u�{�0�,����q8"���3ǔB*��1���}��Z��S���}"�ѥt�ڰ[X�sޥ�9t�S�f����FU�>����L�5´/�7"�~�G�#�dn�IT�wq��`���]r^S�u"�o���uBj�[>��Mi��E�k�4�Z��f߉�o�vv̈́����nt�}b�<�x��c���.�#*V��U�ޏ���z�W�b��+%`k�Cw��۽�;���V+t�:q;1�0<%}f���N�C�y�X�n-�w�j(E=�oӐ/��Vm����<���	*hP�2�@OPnZ�.�}�b N�w/=��V�Z�8��z"�b�/�
��:�Gv42B�'Y}o�6��':�ĭV��6i��RWܤ�p�������E�$�D�/q�S�#o��W��kH�YzGS��vĸ���=Я�_��x6�ץ�󇸐���-|���w�;�%9�{�dz
�Ş�Yv�Q�Q%���N��Br��
j�7�{|7/ՈTos�=ޛ������D/2X�Q�:�ZxHw&R[b��Fu�ﮩ�
؞P�oz�=����E�=Z)ˍ�}-a��!��~ᔽ�/�o�X6��`�$��j�vJ6-�ɬ�g�W���+�}�wy�_Q�i���j4�s�*��C���k��[�Q�߆l5^OdTJ䍭���Au�^9|t�H��7���%�%�6xW+��J48���S�.T���|�4A�R���Z��ht<�������Hb�Y!�T��������0煞J��>�c�(�Y_6�-�Sږ���mw������ՌuSr��Q$������b�k�`��*@�,��3q���0�h��?�aʦ�|q���>ʑ���+��������Gb��:�/I,��ٿ�V*㉛Z)�����O,`ž�׀Ik��'wC�P/k3|�=z�$�D�F���pz��%��yvC����x�줏+��J��N�y�J_2�9�v�#k��&�e卒�L>{��j;<uc�y��cO+^�]|��G�m�B��:^S���3 �rV���7���υ�=8���gy����1��5�����+蕁�L�^Z߾�5V. ����W��}������Z��!�m35Q����5�<�d��ɾ��tޚ�I��}��	�:^��ԋ��+�f!=t&�������d�ܖ!���b�{g�_�{E��.it���=��Q[C�ϽKN�<V+��L��� �]�v��[}ЃPٳ5�s���-��^�rE�{����G��9z��|N���Y��y.9��U�>�W��+͹����s��;�^e��K�J�t��t|~��T=&}�/ÁY=�
�%�o1��-ճcn9=0����W,�o;)��~�.����H�Ig!�U�H\�[�V�Ү�o�a7O��=:���?�׾/b<W@�����vK7�p.���1x}���2!��,�A^$#i-���&��H�C�k�*կh�QB�B�R�I��㖌��J�{�ó�Ӱ��V����_t_
�jX��aw���
�I���:��SJ�OU�K����
e@[c��fa�;�_��Yr�����7� ~����v<�%�Ys۫8x�v�48u!��珉7�8�}�k��[�D���u�'�
��|��s��-�1qӒ��0gend����_u˕���ǉ��J��mfj�w����횰ꓫ�Ik�~-֔1=^]���>簑��������o;V����i"��	S��o��؃�'�٪mx�!��d�oj�{ʺr�Ny���И�˭����e8��C��N��"D&/4��0:�H�hTP�V7_C����#~�y�f}R�6}���b�ˣ=+��#sʗ��6x5c��I=�]��O��ۓC|Tf��'����ӥ����_������t�p��vxuR(JXY��N�mε���'1�\Hr�:Ū�ʠ��y]��p�ٽ�t�����K�A�G��$�T/"�X���>\����u�*a��4)��m�0o�9��;~�Ub�K��4�`�Q�Q{�
���݂���ك�#�L����2������^�֨��W��LzG���7���z*������f�tznp�+���t~��J�Ʒ�~��K�^��W�S�@u�`5�ayP�ak����_TN�]m�՛T�zhB4��`�r.�.���	=�^+Wu�*�D�W�u�!M[s�����Z5��w����glwtm,�{��>05�v�xY		+..\���WӋ�@������D����Y�<3�j�#��N��1��,=��M�T�����=%�ʸ�]���"�x\��6W��,�n�Wf�"ܭ��E`���W]S!k���R�^j��6&l��_�/�~9�1y��u8<h���U�m��T4b?wV���c,}�u���=��z^WZ��޶1>�;ou��ޟvI�GK��O�:�\�����4<׾y��9�����'T�O>�H�n�4������f�2}���W_Q&u_ԙ4t!t����U��<I��$-++��S��~�=˝P��H��'��T�4�#�yuԴH�LUƈ�����jp[�ow�|eML�0�+��Ǔ�"��J��\��o�����T�
���tb}b�k�!�9_����{z����;��3�N_gN�Yr��
8�~_�@�˯e�q߂�ǥ�>�)��S�A�5؅�Ze*�|����6;�3����J?_�v�򏚥s����W�'�>�G���EP�t
�|}n�˵�x����³�;��x��+� ݽ��U��O֧�(I����Y��]Q.�W�{���k΃��-i<8I&�z �+ǹ8=Ҫ�^m�%�����ʩp�Э{�k��+]�'�b��;���I��WxWeo���~�[��`�2L��0�;�3[�����A�wIOXG��m�i�7�fBF�p�o�ݙb�E��B���I����[���w�ew*�Zi+�:љn�4��ÿ����M7����Yc�u���L�\+B1p��_w�u�w�1�����n�h���Z�u8�n_��P�
ع���~��5���j��c��J�����u��rXz�R�>��%�����9.�#*V��%��`���p㝇!�"QW9+��Kܲ���}�3D>L�8���\��k�[};��ޟ	Kϼs&��.�9�V_��\�ڜ����,�/7�:o�,��~��(N��+:���Wg��3پ���l)���\2dt�6�MW��º|��xm�-�й�\I�t�+S�����,��lKxxǽ�}[����w��i�՟"�,H�������y!C�)-�T��>1u�Z^k�]mM�U�Y�=Oʇ\��V5�N]�j��glL�|��`�\��&���r��d��N����f�ω�+Z��E�c�Ȳz_�jE���}�I��(}y���ܱM�љ����7�&	/�ʉB!5#kk����H����*G�"��w$����DU⾠i55RX,	�F����;h+��W��L�6 ZAE��ff���H��ħ����8P,�3B�dH~"l����{/N+�e�i���qu9�Ir��?��c�\�t�y8 ��s�e��-ܧ��X�:}�Bۏ�Z�܃�l˶� �y�i�V�ѕn��3�n�{�i�j��֒�<Z���%qQ���j��{;W�f�}CPṼ�=;yN���љ�&^�Q�X��	[��/�bS��:�w���[Bͽ^�����x4c�����v�}˭+NeX|�Z(%pY���+�β��aN��b͆�gjt&ھ7K�qJ�q�/��OMX1J�U���/�u�s��+U�j�-sCE�]����h���,͋`��	���o�6��x��ʼj��FP=f��V����'�չ�V�W*yV�	pfhʳy��!�j��f�չٰ���lh��Ku�aY���|�wLc.�[�!��:m��B_2/;�I��v�(b�slX���_�\��(����`��{�ŗ��_l��~��W�nH�]5�U�u�)\�lV[���&k�Tk��ݙ�&��C}ZGf4�MFo@��ٙswFl7X�#R�e�l���ʝᐱ&{.�������z�δ`U8�2�J�ꥡAp�)b�R��Μ1vu���{�7d��'�#BW�x[�n��:�q�9"O-�v�v:fӽ��ݭcs�foN聡�Pd��ϴ$q�͟�xd�5ne���G��DL��]C���ru �M�]K�U��h��Ua�F���R�YW�]�-��"��kR���Wn�	�G&w��
��rnֱ9��*�h�!�Ӻv
M��R�U�[���o�<���8�hf�Q�e�WMEj��ŭ3cF�}�wXx̊WvP�^�%�"�\��*A�)�2{�YLl2�~�]PH�.���jk+cX���S��&J���k#`�e0}R�7�`=�]�5���"�kj�%�fk��_RX��O�+ueqObۗlk���
�:Nә��:�E�-3���)��I}��.���(�aH�!��\����W���Z36p����y�!Y�W�vޞS�c����n��l���ݳM�˒|6�"��ޥ��������豥�����#p�Ȯ����ocȄ��V�A���3��2�@ox�)d���lySJ�Ftb��q:s�q*,j���x�-kp�d��Ji�- �mc՝Սu��Sq�-�ȱ�pe�ۡv)w�M\z�v�֩Q���ݭ���#a���$��`Oe6�ɹ�6e@r�r�h��`�������1��/b寛�u�H�;`<+*�.�1��V�=xݣ�!�t��L/�����=����v��[|��?{�dv���&�@CX�9���^]EW�h��+B�ڂ��xM���os=^S�9�W}�X��gE�����e�MB�3�c�ݮ�>��o�׆� �� ��k2脅){����P9�TXT��T]��L�$(�d��BB��
�!V�A�Q!1��bD*�D,DA���*�$@R�A
�tq!�
Q"� H����,N5		��2h �$�A��I$A"J*�	ƴ�"#�L�%TT"�Q��DP$H&@��D
���&c�h��J���D���.Q*D��"�I2d �LDE��R�JZXEQФ"(��P$��"����	AH�m1PX�*@��*�"(��rk2�*���X��'6R�HѬ��bd�H��
^,ԉ�����wϿ����mXƘ����Wێ�>T�ͥ[�6�
w� Y�Od}�����u�w��5���٦��oX��	�\������r��y��>�g�W��a��:�k8��<IĽ~�skK�׉;�t���İ�~�[��/i8���^	�n�K���I�X��ſ'��t\�$��".#���C��>���e����g���ʦw�g�Ks��:~���H���U�#� #�o�{�RΗ�n������,/I���/�),&B_<�q�9�սsK2�z����Խ���I��<Y���r���$����Z`+X�~�����ة���Q�@~��>'�~�����;_�w5�/��󴾤˖��<�HK�L���v��/I8�$���$�8���U��'���~YР�B8�4������	��	ص�~���|簿�<^$�'iǿ�哥�'�����_�;K���|�N���,�Ϟs��_Rq8�o���:Y�d����������{����'�~��<�[�E�8>��Dp��ͻk�[.�y�C�s��r��%�{;ׯ5���dwz��_���/�7�w�n_�8���>u��X_y�O�><Iİ���]ZBOS�8����[ך����{��Ӌ'�ۏ����1����=S�s\������^rO�e��'�O�:Ki�ϒm:�nI>�s�O��_�;��$�'o�x�|��ygI|I���~��S|�̾��?{�v����a���[������D1n'�1������v:*�H����,��|Y�t��q'�ix��q>���s�t��gSn?�$�X�O��:Jz�V�'{�����-���'�����_e�ws�������'����Ꮠ���U���	8��Ę������>���~�ē���rt�����s�}��?,�Y��״����.���?i:_qx��O�9��X_/�OWĝ��{�i�'I�d�擞i}Iđ�>ڙ""�>�>�#u��~/�׾S�����ﰏ�����C�&/�dQQ��˒���ߩ��<������h�'�rϫ��[�?$��oK�o�;Ӊ}^8��M��N����/��4�~�ia/��b,}���Bʍ��`��<����y;���t��q�r���ir�|����x�o�{����|�[�t����y�,	���O���~Iı����-�z���I�oN/���Ϝ�ĝ8���M�B��TG�T~���p��d�C�mm޽�Y�[��5m��� �=�o��>���c���$9�,���.�G����
"��Ycß��Of����'�A�g�됆],��8�WN"���a�J��L���8���P����^=�˔�](��K�JR�]c�Ae���κK�=�s��!��7ş�:�[��:K����o{K���y�V�������;_V�k'��\.OVq<K��|��Y:_S՜O�w�'�>%��W�5>,���'_�>�2S��o}�}��]W}4),�v
�q����#���~ZJ_�$���iž>��o_{�?%���I:Yr~���O?��<K�>����$?}�I(3��B�������ƿ$�F~�� QG�� ">�I��K�4�I��ԝ�^�OS,�:������/d�t���'}��|I�X��o�~{��_�rI�o��yվ�_�}�D[?|��#�I�wk�7��q�����8������)�|����4����X_��q�N%��HII�~^�7Ic�iru'7�����ěiK��o<��~��^���_����}�#�>�F3�O)�B+���Q����|[�~潧I�߮/��d��N���?-�s߼�q/g����,���擮��x�$���qrݴ�8�Si�ܖs�y擵��sK�３��!������&�<?�:^���>%��:Y�����q'Ia'���R��g�8��kϚL��=[�=�'����i�ս���.OVs�d�O<Ӥ�o�K�':[ēǎ.L��nO�؏{z���ͬ�辫�"Gѣ�#�z�%�>�}K���Y:_z�I�}���q,/�N�{���}^�qd�=��%��%�&O���N�����q�O9�;I?�,���^��żKě��%�e�S���c�\xZ�scw^�M[����y!|N��ܒs�NE��/Ks۾r�s����~I��-�/��Ŀ|��u֖e�/�޿u�v�'ÿ|��g��g$�O��y/I!	>��6�%�������z��ù:<+۬i�8�}�B>�C�D�s��q|淞k;�$�,/ԝݯ?i~$�X�z���/�ܿ:��'i�߮/�����2_gս��ϝO�a/�3���z��|�K2���z��[��.�?�ξ&l8��׿�؏���CQ�U���� W�q=��t��rXw<�{���z[����8���gso��,/��c�}I�'�}�OR��Y���:���L��>��~����z�~��$w�������5եA�ٱ�%�.����ǫl� \��1�F,�u��a��:����Q�D�|�^��J�PJ��Z���/%�Y�QJ�E�!�b ��n�2�YS/�;��Z�aZ�48��8�c��Dө��%t\FI|��cB���d��9�Ǜ���k��}��f�䪮��}�>�>�=�ޤ�2��K�?���/Ź$�����I����$����v���Y���q/���O����$�x�y�ԟS���>N��^���'��g�L���	[���W<������d|H+�}\Ľ��{�ߝx��I�e��u�Vq=}[ļO����X<��N|�|�_�;K�S��Y���ܗ��O��[���gs�%�&��xwy�'��I�4�'_�Y�!���p�T�e��Y�M?�h�8}�qd뛋�����>��sI8-!'���z�$��=���9z_��ռN{;ܖ��~����I�O�`O�������_�8�֝���w�$�8�[�#�C�/L#=��U~���K��������g�N��d%�{�n�-�9����4�o[[��:I��/ջi?�\��nO{Β����?���N���g��w�/��a��|��y~'Ԟ$���{�]T��g�>N|^F��3������_v��I��'��5�$�&_�;�s�~��_Rg���o^��������|s�/���z����$�?��޻XX\�;���d�;Y��/�=�����b$Dp��;;�4�vs>��g*}��іe���{��O�S�a;�����������afI��e%�4����rt���������K:O��x��|�i2X?ky��'i{I����{�z����V���lbf�z��o�TW����N����~�^��4�%�7�o�{=���������Y�N��f_ϗk>:Y���[���ŜN,���-!9v���Kk;��'K���/-�>y��-��~�;����H�޾O���q���'I`Og<�ս���IĿ���:�z���Y��$�2x������O�{K�L��$�:B_>Ɠ���9�Y?8�n��_���֒q|[�����җ���]S�Z�l����yŨq�Z�q{[����r̿SŜO�ߞ�/��,/I�N���2~I�'O9��.~Y�����g9��O���9oi'I���=�u޾-�^��4�z[���~XI�>���J�V�Ս�e�1�=���͸�I�x�%��;x�aar^��:K�?'z��I��O�ğ����{���$���z�z���X��r�I�z_WĜO��\�t,�I�w��'ic�/���"�}""(A���i��D�u>��S]a�ϴ�K�U"�>3��-x���!����L��M�����o������u6.Vn��y��A����}�n�0�"�Z����f��^"p�Q9����u��2vjz<�]M��eX��� >՝�c`�|(�)8�o�I�,k;�~N��&I8��������?��o��[�����r^���{��9�����{����&�K2y}랥��g�����Y��g�#萁�Lum�o�\�{�}��9�P��=�rN��N��Z�<�qz_Β��'ͯI�X_|�|�u�K���a�뜟V�t�$��;��z�O�x/k����������s��nK�Ly���� �ю�z&�8��`�0}���d����-�[����s%���m:�I�/�'_��K�4�_����|O�9�9��_��,/ru�'坧ԟRqg���,�_R�՝���;Ki2|Oᛵ�ڻU�,���/'>��k�?}�'����9o]���%��sޤ˖�6I;��Β��&[��w��s�}I��[�|�O_�,,.I�x���qg��pY	|O���sO�|�̿���zI��$}�(��^l������?��Jp=��/�OW���s�O��R΅�Re���i:K��d��I�>?-�I�>��S��fO]-��k:I���_���I���I������oI��%�9�'���˓���}����!?w�m�bUF���
��o��,��\O%��|��e��}_R�qg�q?��ܒt�,�8�����N���UT�lǡ�̭uPt�_�}� 0�C\���Fk��*�{7Êyȡ�2�V�u���J�{:�7�8%���`�[d���ۢ�Q>�m�s�pb�w�$̺��s-Pf�"rf���ʦ���*�p|����ޟ���
��cݦ������._٪L�=�m��T>'���s�>Ky�������V����n*ލ�B];�;���q��ᚭ��܍�Qq'���ưW�{�R�κ���{����!�@:A.�ɯc�u�rm��l���>����(������Y/���h��������t��h>~8�
4�Ϸ�/n�V�Ȅptl}���fQ1�d33��H;��N�9��Ӷ@t5}|�۞�
s0�ͤN1N��__����|9���Tz��~���`�.jäB��<$C£�w>��<�<92��L�����=S�o)����%̠���5��4͚�oӖ�b��W����|�O��HPEc���U�9��0�X�:bL�>�ʆ����w�d����
E���g�Q���ʇ�QQWg<���/���Մt�y[�,*%z���G[�ZE��J���轩��u�px��9g=~䠒xW ���Z�A|$���rfqv1���8R�a�ʪA�����N����C�-)%a;���D�a_6��|)��^��]�;:wy�I�gޑ�+ٿY�[V3�X����G�	<|��4ۥW����E�y}L��]���Y�]7ݺ����q�К�׆�|�Ϳ�H�]��%��>�����U�����ꗛ��'�_�Rv,���'şb����d�C�Z^����x�����%cҘ+}�7ڶ����v��ܙâ ���vV9ѯY����jU����& ��S|;�r�A���j���-יB��%MY�ə�>��	��n��m��8�6�==r��9�`�[����n�u����<��3�V~�)R��s������ �]by�����өN�kf̜4�e�����t�ёed���J;Y�����U�l������}���ַT��ެ���Q�Vl�Kq����_����Bj��³��d�rX��Z�3]�j�}�2��w�p��Py�:�}��̕EWYt}�械�]�ww��W�0N�RXy{8��I�؁�[� =p+�n��׶c�G����%�U��hǵ=NH+�T��r7�9�S�(��j�/�(�WҜS�z{�{�r��j�Xpy�H\�s">�f�I�{;���GM�~���㹝2���������j�
�ҁ���"x'��f�V�7�͓�_i�����������|�>tWC�xD��Ͷxʧʘ/�?N2��
��w������9y�Ԓ�Vf��+ؾ��<ZK�d�w$l-��7��*կh�q*P�a��G+�<7N�:��[��j�)b�}(qX�n���&��~��A�A7z�#�~�]��Qѩ!]c�r\�Ͱy۾�W��Q�[�[<���G.]�W�N��D���&�J�o|6����c��3�b���ƾȬ|��嶲Ua(��V�$��XB�T���t��`�B���V�90n1+�����gcpWQz�!��U�^�?;'a�abDł7�*
vu��7W�"$q���7�We�V��ᱚ�r����6�832F��|`�;0���/�Z~��hJz���/�tT�vjPك�[��`]\h-��}U�����y^�s?�2,"멵�t�H���HgN�k��8��dJg�^a׸p�2����W���z��\g@v��uh���.�7���\�3Ҹ�
߽��0�����6���^ӥ���%�1�{��[����.����)��Ո���������}�Ww�a{\o[��yPk�@�-����R�+�=TRy�&�k+��l|<]y�8}n�cY���yru.�K��{<dJ�W��y��� 8_ySdhS��۠`������K7����UcB%G�JS{{޻	6`�E�}p��Ġ��|�5����6*":��٧TOCz�A���_P�y�A��f몹K��&�mP��?	��[�%��ֻ�	������C%�r�6wQ�'���K����Z-���K���fuf�2^���t�*�H��q�^�s}�J��G"����̻B�T_2;����Ujg�]T"�k���*�cT����l��]�62V߽������y�|���y��-�]5� N����'��3"X"DzM?~��d<Vu�3F� �U�]JT1hiW�����U~��ܶ�Ϥ�w)��a����am_s��n�2�	)�q����/Z^oǊi�G�K{f{��+������ل���9�$���Vt<_jͫ�ݺ\�c(7iv�q�{Ͼ��un�V�w��]G�����ﾁK7R��G��C�#A���d�r���,;�R�c�I;T>���׵m��m��]d�=m��)�=y�Z��__�t��>�F!�,���z���W�I�� -�8zd�����}Y�l���8q���=����UCܚB��IH����s��V�4�!������<N衁vdl����R2�o�gi����r��|{)�H�7�bU�{Ζ[u�ތ���$�Փ|9uE����a�5�������#�u�9xzQ����N�,����w2��"�w����}�|�ȯ�_;�|��А�y�yN.�Nf���臄�Zͧ�*X�/f��+�U_N�q)�ʄ��E�������*���XO�qh����B����>֫�5Ҭr#Y�4�����k�b��nJ���ߏ�3ƺ�\�V���ON��v�<�e�3qO����t4�]�s���)xb��_��J�֕��Z9�����x2�_�f�� D��߯��n���z�;��e_�L/��+Q�UPw����i�y4����O}���K~�J�=�'q�(.�9����O/��"�ۨ���fv���ѷʹ�C��:���j۵�_S����]��sajǵ�^��:��} ��<(jQ��y\?g^�O7[���N�ш9-��L=	������_w=�A�瓬xGb���꯾���$��SǥpE5�֤0�`��{u����r�g�u�o�pK��ʕ�tUO���۝�gBj�}��y����WiiU�|+�x7�*����5�-����I�p�Y�n[����|eKmmJ�ط�ǢVm��C�{��
�*�T|�O�����VԺ�������ič���ܷ*y�WJ^z<4���HL��8Z]N�~~�-z׹��4�:���q�+�Ξ�y�)sV"�<$C�ëէ���L��>�yK��^w+��Մ���x�hC���i�5zߧ,�F)� ��;s;�� ��f������q�s���p�U�ER�L4�G��������"�=/�"�<��?������ɛ,Wo�=���Oj�Z�\	=��R7����CXGr���R?}~Ϻ���+��ȳqܣ�V�������\�E�|�-W"w�HUt���}C��.�2.�
e�zw��;پ�5/,#g;]�ӮHA�ұ$�&zX���+�խ�hSۖ�'Ύ�{��a�yHwg	"G��ޜ�Z�Fg���
6Z�}c]�C�S�5��4g��9��Z*�	޾��6H�d>�{��'�:Gn�`ʝ5웮����t�J�pya�r�jP�F�U㬢VV�(���b�-H_V&d�+�a����?0��AV�l>��1���>��^��xA!9w���w�?�Ƭg��(��A\ ��1`t�I���~����v�_�͢��F���iY���:��y�������K�E_N�d��\�P�C�+^��=t\�7l߰Z�eB,ϏX��_,�p����X���x��C�+藢`���|�'y�oW��h�,{�mH�Ub����N�C��������!�L�Tlÿt��R�����%_S:�
>���zomr[�c�̔W�@ݚ��U�/�x�7/g 7�tg�o�S!]��	�V�@��W{g��ʹ���oڴ�Y53�l��CG�~�ÊǺ����Z��RŌ	)I����A����ǵ�w�G��oU�N��:,��{����ہk�Ң5ex\���^����{��%J�S�v�{�{�r���t�hb���m�Www"��I�cXK�{U-�	��*��0�@ژ��"��V�윸��3AgMB{(ʦ���F	)�XԊ�U��L�o�U��g�-5M
+��~�{G��U/5��J4/��Gz��L����u�ru�l��R��v��᎖t�N��/Y��x���,ў�4���vթ�uӇd�k�׹p[����QP�h���.�HbiO�}>�N4Fk���t��1�/��U�+�ߖ�({SFj���OK�d���*�ꆕu��+)>=H�H���k�|�j�+A���u,�̴�1�/ta����ե`r�hv�Յ���s�G(�����I����mp-��*�KyLf���8Җaŗ;��ĵ�%���u�%*�f�`yu�o��9b����E��>�G�)SI謬+�1�f����#����i�yf�aA��=;��;�B]�hN�Y.SA�(5�cJ�f\��xl&:�&�z������8�u����tX�hӀ�6�<�Njd9u
��&��7<��NB2����^q��(ĸY�ʱRwn����(a-���R�w	�(b֞�W�d=z�R;T6���'[�8�7��� ���-呴{%*�M�T�$���5��N�6(�P���<�<(̔T��U��Ҭ&r���_�1ݖ�<e���Y۸}�Iw�P�T��#�'�m�y%��|e�W�eaAHԜ�u� -7�:�a�E���94� �^��X.�]��}�f����zy]�� �B7w����rd��׏xL���?zwY��v��з�v`�n��U3���qt���)�y[b�����7�>�T<R��r#8�O�.gL�a�4t�.	�㴪^x���q��{�r&]~�w���I���}�ۗ�ײ� �iX��m+�v1�n8	�ﻹ�ܸv[�\p�Bp:���3XD,�o�<c���5��j�B�C+1M�7)���i�(��j�SQ���(�1&.��=o3���놊����4^1��liSz�u�DM��l��50�U��n���\c�c;���h]4}㣴
�)?���d)��ܾӕ��0�=C֮�Uՙ�wnOz���'cǯ>p�rj��dv�u�����C�2,_13F�vi缲����2�s�_#ne;�OkJ� ����}-༣�U�w���n� $��0]�$��Za�!���M��O�������(�LZ�Llo'q�[�:��ꏘUé���4��Y�Õt�ǖfF7]C���ᬡ�jD;U�(�ǐP3���9���=�ڻNQ����R\>�Jt��6����É�ۍX���!F��6^����,�������M�C�LAswv�YdL[q:j�������K��}g�
��P�6�;��͏#j^�l�c���0X�[�z2�.T�%o�t�4DR��N�c�������n*�8�!ڱnMMXjfw>��#`��ȸP8ZllT���w}�t[�C�"�V-��N6_�][q�&0[�R x�0rs�Ui�� z�;*��.V�3rR �W��^v^�_�5c]�췭�x��I$I6�4�FX�P2�b��&�,P���8��4B""AU�� �@UUCk��eEdȱ)$
"b6�"e�椚
�&\�M��n9"8�PJ�D"���j������E���3�M*��@�H�iM�����B�sj�0��H@-�iDB�D�&ڜj�TB� DDDYX()�U��^iu��&^Hm2BE�ʫ
�B)b2d��"!@�Ni�k�� �Dmv�\�1��!R6�f��#4$
lI�&��HA�M6��(�	���;��h}F�f���Y&�q���2�1�w��0�4�oZL��̾L�\�n����m-#��N��Nu��������c��V�:��&�>�����8�(��
�4WrF�[C�{��aO	�l��9�9�T|��7����G�\hNK�xJV'N��}I�?	�	n�-�!�<<;]y�<�d����Ǯ��3y�Rr��s��r��&�G.]�M$�>�Ik�~��+���bJx�Kb�{{8���n�k��x�_��[j%�$NV�$�'���&�O�^���mۡ���(:��[P$	W�]S��ߏS�ڹ!���ޖ�$��C�+"Q��<Q�U9��d�H[�Uح#@�J�s�;xTB8�]�xoS��]�q�B7-R2}ۺ$� ����d�ڧ�:�}��Q;�R5c�V�t�V~�����R����f��"w��N!���F%�������[@��^'_�-Wl���y]�U�:��/샵�Qz���B%^�u]q�]�<�f+�|V�P�}�]`bie���yn�}�]@�n�<��W���<7)]+4�w�l��V/��ݿt���5,��(Yٞ��x1�>��~R�iY��f�n��'������ �v�R�x-K��՘ї�U�̒��/.(�Sm*��U�ớr�Ar�A�u˚�H��Xg�%f��g��Ɏ���W�<5�aU�f}���x�O=/��yl3�1B���B�w͓&���"�����5���}_W������q�di������4���*������KE��t��ݕ�����eF���}��U,��>}Kz����U;X}�ӳ:�mS%�U�E��+ �s�v������q!t�Ը�(��·A�����/
t����X|�x���,�Ov��OԲ��>r�]R��*�A����	~q5]l�[�c����.�Oٝsͧ�m���Ӟӓ�s�,��_�
�i�ir�ɤ��NA͌J�v�)=Z���S��8��Y~GԪ��b�O�t�:�F<���=���K�ρd��� =������M~�'�z�� �wX)�z���i���{�{��P��d�����G<%[T/�����Z_�;��GpsP"��ӇR2�����#g9X{�ǳ�s�!�{j5�	T0�����e,Q]�g�%OW7��G��_s�b!#����U�R�=~#�|�z_YN!��b��A��5Ks=ɩ�G9)��N݊�-�T:�C-2�ߩ���f`� 宔ƴ�b�j�<	n�W:w!p�P������w�X�M�N�le>�Q]�U���E�XZ�Z��׏���a�;��֯;�X�R��"z����
3��H�5����������3���7{�g-�3}���$jwzW�S��������\�nN�R���w_X��%0ʄ�ϭ�\���&���Qz��XO��6)��>���<>|v
������g��#�Z��	,��J�����3ƾ�u��z�(gj������}}Ρ�N���1!�TBO����!��Y� ����`C賛5����us�Dγo�{=��wPW ��k�t�C��mv��ѻ<���j�����-r��{7�Q�-W_��	'��|���mtN�4<W��i�8���.���k�K=�u�o�r]�G�#��1�a��jWT9�}�i���ZZ��
�'B��^�����Ms�U��(R�I��y���wK���*3���Kqn}|��>���,,x��+� �](�-8��E>Y�;����z�ɾ�]���D�����R���e�_v��妒բ�Ea���u�㫣C�Z�ٛ��������W��~�y�\�4�_���"������+��秨ou���)4�y�IT�d��a��� Z��6j��@�����Yuɚ��o�cUt��Z�rh���=�=�hU�_Asg�?�=�~�53a=]�X��N��cvW/��w�E>�~'��5J��E�Tp���D��B��q�,EY�X�lb3��jq�s��Px�yo�]qv������^ٶ�r�.nDΞ]ˢ�`戽V���q�<��y�b��/*6�?|>�|`�����Aε?��^+U�0�P�ˢ�����E�����H���v+�9��b녪]=�-F��Ǐ��>�	B�$�OwD��R6�G[���]�｜�]!��h�M��O���5��/�/	�¹��-q �����4d/�Q��Q�����rQ�aѿ`����~g�m!���%�>�d�AD:���am#V�2��S���*�U��QU��v����X��J]$�*	P���C�ӻt���_]ǆ���`X]�˓�e��j�'_R�v�j���Vj�3��l�W�ΐu9o���%��Wd��[TuPW������\Z�<J}�uaei����v/�V=�>:^.�� n{��_D�t���=�{ͽp�擎�o��A��1]̸��PUc����<&����q�<W��]�[}�����su~��{�%�����o���H�9�'2Q_yvk�5^��6���<p�x�wr�:�WgH}�D���3
��_D<:U�ճk���hM<M�|Uu�}���5��C�U䥆�ֱ?P�A�rẚ�$��mǲfz$�Y<9z�H�gL^&{yoR�\�F����̜�νŀ�x��Д$t.s)"[Ǽ޳\�tA-,O#]lҦc��p~�z�S}s�6����&p]}�����[�q�2YE�� >��]� 2�fpg𪧉nR0�]������Ǵۭ#��o�r�!F$��N�w�z�%-y&��e�I�P�h~.��� ���@_�QD�'ۗ�;>S�����+�3	�B"S�p��*�0z�yh*�X=^�Kyb�O��U n�G�o��z�J��J�Ff��9�ߧ�4��8(���A�xf��,�e���Ef��~�[�4Q��	{��LK����'���?	�d_X6G�]aS$䏾[C�z?XQe�0 '��QM���V�ZU���;<p��q��u,]�(qX�۰��5`��T4w�/��[��~�w�ct[ej�:���튕'�	^��\�OW�Q���#�� q��iA#�9�K佄X�lz�c�·��g�9�md��$X%m�^�{�����nY�8l�1�|�~�I��4H$6�����N�=N-<����K^�JD>R�%�ݖ.�n��6�\����d�^� �)���Mh��]�xoSծUx;���(��q��~��=�R݇�Ҙ���&���q�x�s�ř�}q���-)o����Inx�<�qbi~�e��h�U�ye��4������{N*��Q�ifocI��j*=�QA=<^�Q�j�<+�eq����xs�r��9����� �����V�{ʗ�%��Ec���*J�4�b�p<�}C�)v���;�{�P�xB�^�ߍ��6~�Z���JP�ڧ����A��Y](6>y�Hx��h|��F��B��9O�A���r�P��p�=�a{t� 8_ySdhS���۪���c2K�h���y �^w���^
�as��2���X��|�5�����ì��Juzb�rz�7ٛ�fk3A����V=��4���J�o�׹�<J��g����ei�f����ΩS+)�8�\���N��7�-�K�iy��N��ԙ,eD�N(Q�W����wt�#�w~���p��}[��3��_
,Z��YU��J���i�~=�ˎ�LsNazߪzn#�]��K�F�T����>U����tׇ�$m/�U�|%4�J[��ޢG��~{w���T\~��>���I�9�h3�(��_��V��>���&�e|����U�n����3^�U�]����(�
Y?T�1gJ1�K%��޺;���v
����iީ)���乨�f}r�� �{�z{s�2�+񘚧[i*7�h�Z��D������b��(^zԅRs&=v��s�a�/thZ�w��X&A��(8^�f���^Y9�����N���B���®�M|�T��d�;����҉���������:�2��'��
L����Y��<ug9p��z���*�=����Ih��|�5���3=�r���b��"��.��T��l�#g9X{�Ǔ�"�mF����V���b�Øvs�8�#�+}.ڣa�&��|��"�N�8/��t53W�ܵ<�L�s�V���Gi�����k���_���u�r9U��Am�h��/�9�V�� �9]��u�p� RvO�LW����=E��_X��A'c�G��,"+�M-�U��e��̊��^١c�:��}��*[ҙ����Gֽ�׆(If�N��U�3ƇTK���;�۩wL�CQ_&=C�ߎ��կ'(�40�����{��D�S��������l?w8�"����t��U]`�
��ᲅ���G�s篴�7[��`����uBj���T��W�c��۩�O��PV��."ʵ54�Z�9XzSV�΂��n^�g�W��Sd����+!M�s f�׳������U�3�J˶��4�*�}�<.�N�<��R�À߄Ս 2fW�C;E��B��~��hӳ�*s#�f�q-.���3�p)`�J#{W( G��xmt�fD����?B�wy�JY��i!?=G��2�Ur5�N��%Ze�B��v�^��v�KI�}v:�y���>�O��5���㣽���}���y̞3މ�+�d5|��T�>����n�ћs:v�(��t��9f*�Id����Va~R��/������m#o+����~�y����[�V�h\����6=;'g�R���ǿn
�o���c���$>2�&�̖$A���������2���.�ʍfqҬI!e%,U2h��<.�����Ze�5���J1H�֑�u��à0Z�8�����5P/�����F�� p����͌����wyOK��H��YB���,�jrs�%�W��>r���~��!�I���Q+�ԉ���qu�QJmө�}�w2��_L)�^��7=���{S;�K�K�M��(�Ɓj�"ajC�����������Qi�["��'�9Z���u�|`���R�B���$�'�'�_�(�_�|ژ2�U�+jok�#��Y��eI{k��"�g?}�j�7BR�֔��\$��hx�T�P��n�Ү�/�J�ټv���%����|���������;�zGb���]��$�zj�������ܮ���[7X��۶���M����y�=N4���ݛ����D^<��6xz�0���!�Y�Y�W�����_14��EH�U�rڷ|#ɜ?���<᷸	��T�6u�*�f0+q�׽�r7��O:`k(]�[�kMk��39Ïr�� >�o�n�<0{���C�&���e2,�?��?:W�<%�pv�ww��W��oi/5x�+���̿�)���r�C��b
��g+�
W�^ �����Ki�2�7�o�Q���嗱�=uj�u���e��l��M�8�.�xjin���Vb�]	��{77�s���Q�nոNRZU�_f�*,j�K臻ɋ�u���j�s%QU�|go��r��y�o���ޥ��4�i;t���o��u�m/�Ǵۭ#��o���)	�5��+��v䱾������%�]Q[bT�kE��U~	E�ҜS��p�AI���`�ȫ���HP���3|�@�\5Z_��u�e!�WϵK�xJ'�:0�=݉�&J鐾�����^�>��xt`��x�o(�P>������O�0k�V��W��:�i�|~�Fe��%��#𝊳���O�:�+�@��[����{�?^���=x¹�~y��>;�yq��N���%+�n���&���	WP���K�=�����EN٢��4q͝}�ܹ�h�������렭�t�ɒ���A�6�]G�/����V���i�Z��7�@ku�QYWMk����@r4�T���]�Ԫeޠ1mԔ�v�`��lP�V��h޽�x�rA%��G�
Y����������z܆��9��$7Wfq�1��
�Ï�z�-�%��MA�v�XuI�f��=rwr����l5^�K_3��V�1=O!����|��r�O�U�H�J�¤���9�sU��+y����E��>�H��Qk4ā"E�.O��P\�ΝrԈi����fb�ד捾��Nl����vմ� �ߕP�㷆�:�k�ާ�\�2/[*z_d&^����TѪBt�B���UY��ԧ��Q/�<N�����3�_���
�sW�j#d��UG�y�����7�{�1˻!�z�%BR���s,Jy�&�����+�+�M6�!���OM��[�.T!��Å��T>���!����>r���z���F�1�$s��p��顓������E�Ƽ����gS�۾�B	�������:�_~�h��s��@�_�#�"�\��+���k�yw��U�&�j��Gbw���Q*#���1�{�09ñ��?{x���[�l�K������KX}��N��ͪd�����h�P��5u��Ȓ��i[`o|��w���ֈ�?e��"]u_^�\�/�j�nj��vLF�W��{P�ϭ�,ң��j3��+(���]u̹9��ē�ɽȐ�贬�b�R�w)��}�s����]��O��oT���^w������72�An�vnJ�UL���=�\o�Vr��l��:F�F�X�8�Z��R�7L5�(dQ	ZW�f!O;�rOJ�ɼ놖�4䉹��[u������J	0H�-����u�<�c��%�U��T2���e���Õ���ʙ���3;3�ͬ��c�]�1 �4�k�Y�NmL=2�+w��:��҃��]$�l��k8j����ukv����S)V
���bƛ}r8*_S$�uҶ�[��U��V^��}C�o`���Q����؃!"���rk踦�Vl\���^w*#������x�~�Z�(��P��Q]����W�[����O"P�m��ј�#�(9��d�T�
�U"`�,��9����N��̰X�h��4X��I���@�4��w��a�6wѣ�;�1�Bo�9l�;ƪ�b����Z�7���P�#.b�)5�Gsc;Yaz���ؼ�Bkz�\�5"��Ƨ-�U�4��(�r���Ю�I2jN��U}�fP�"T|�{6̗ݯ#w$�|�w�����}ܻG��+�����Fu^	�}Q3��r���fLn����&~!�S��n:�J�{�B�O}p�7	��pW^4E�];s���j��ө��Ok �8�y��Q��D��w�Y�?B	�<7��nV�f��P���̂���M��v��7\80\���D݆u>R�nq�c��\#R�&���1
�{�;��$���C�E�ĝ��V�!�^�	nA�������,.���,��Jfʻv/��˷ 
�V#οB�j�d�,>3�mzϽ���{3w=��:o	�)�r�<g%,+	i��� ��b9҆u,��4�=�������x�D�ȘFb|x�A}�q''�c6�+j�|xd�g$�_Z=/��fȝ�B���3Ǭ3wN>��� �)ƻ��3������d�ޱ�R���H<Q�B��e�-�Y��{]��l�R����e���urUv��;�#�&����sM��q�=91�[���L\TĽ�։�b()��a�XE��^���Ȍ�^��}�>���joV-Ƚ	GOy�5x�a�e蝬�|��.ל%p�Ljc�;5����>�^�%;�#�o���{j�����*�욶e�9E��&S� ��w]����ُO�,ޮb������m��,��6�D.�r�'���P��g�S.{�M�J?���gg0f�ov�Y�i�CG���m�7M��J:��$��U+pQ�9�-J���p�&�b�'{p�,��Ƴ;޴��N���С�N#N2�\��V=����4�Y�t�|�h�EH-4���
H�R�6�Ci�	&�BfEUDE�͜�h�Ɠ6���L�6ȋ��T�6�M��rrD"DR)Q#���i��2�rḺۛe�l�"�]��MsH�S�����fH���6��f�g5�����m4B&�M���&��^',�Ѵ&�Em��J�����وm�D$L�A�QH���Ms6M�J(B�@��5]�m�� WDL���6�"44�i��D]5ۜ܇8�,riHB�h&��b�0M�m�m����� �A���X����ؙ6٘D�m��XBe�m0\mU+���"! ri�Ti����8#��"mG�B$%|ADc���ΪW޵ݰ��ּ�&�|��2���������z�=<c���*dg�*�g�(B�묮z�&#	�q}���}�}_Ty�$�o��I�,o��}[��3^�|(�l�t+·Y\#������Mg1Ǎ�����uN��{ ������)��dp��]���r�}�MxyF��S����»�����z����>�KU؍��xt-=~Te�W��ss�nGK�ĞP������L�כ]J���z�X�m����
!Sk�
;��#�2Y/W�޺;���v��֫�yv��YT�O�^��K��]E�-���w�|-��^����P��g�R#P�'�ȊT��q��Ȟ��:��(����|t�8��g9=��)�H�����,�Zk1V���tw*��U"�rX����*7�M[����F�t���b�]C_oȈ�5eۼ���;�_\��Ò��
8�~��\��zW#��U��m�t�"k��*w��J*:�019kZ����,κ��w�(N��G���E}ɥ�T^���>��W��Ϙ���̯	�I{�/h3���E��g��#�Z�	,��T'TϚ���3�7�7p�'yw?��\N*Y�)����^�NJY�YV,b:�*�L/cL����`�I o6�����x������:Pʌ�v���3���ac��;u4kk+��<�\��rܻb������g����zlg�PWU��8���3�/�홳��P�����}��uo���R��/$�|
��gf�1�A�:vS���G���,�K����;�m{Xn�d�Pv/��pȔ�
�!�݊?Z�Iõ[�������!1�gz���s`�ޱ����b��⼴��� ̯�U��ճ�������;���GM�t�u�޻�����zT�;��׼jV]��W�������v&,����s��g=���l�N��5F ��*S�)���V���ˮ^�$ߕ} �5���+��3V���Х��m ��j�����Ew�{�r�!J�h9��Zc���f�"����O{�7I@
H�T�*���Br���������13�B��<$C�÷W&��g�R�c��uYHo�M-:	8���uѥ�C�}@�m3f�[��t���<�בX��<�ߗ�A��ߴ�I��m=+�r��Id�=]M���wy	�V��w�ͮ�J$��z���<���j~�*� �z�MX���D��ԍ���:�N��C�=��&��NZ��Zw!�U�0'X��c�sf�Vu!���k�([8E����p8�r�{��X���� Q����P�n���HV4�*)���;5e湺���S�0��$Z��� ��t�{�" dͲ���$_v~����}�@`���7�9N?}��3�V�]6xW/��Ak��5�|X�q���dߕG���[�ooZ��/p���Gǜ��>�-�=�CJĒ��}2xQ!��puR�s�g���G���m@�#T��ׅ�F��9��ocV1��]8(
�E�2�{6WB�]�jW:����h���.'�@���:�T}��]�m{��|�Ϳ�H�Q���T�`@�*},\�3�2�^@�q:6�S��?����W�<%���s���M���c����N_P�����)��K�Z9MU�܁=@���C���W������'�e�3����q!w�.��Ϥ��3\��y�����7�||�.�{�M-�|}(��!���p˾c��x��y���fj���;ГnK����*������&/��{_��q�$��8};i�M�jǁg����i&��}�Xi,�;t��m�B%kU�L���Pݘ�lɻQ,�w�߅��oF�����m��X�W%���q��P��Q+�N)�������%�1�*�n.A�cydȯ�+�ޛƗ��ޥC�
��:�t*}����w ������� �p��ཝB�1����{��j��-棘J�`�o�<�C\>��f؝��3Q�-훬L���;D�O��߭������Y��Kxg�����Į���Wdտ��B��6%T�I�4t���/j���`�u}���T�Rۏf�|�E���\��z�X6�Ԓ�O'���/UZB�v��2A�3�ꮾ�>�e��c���=m7�:񋗖4��7�~��-���-m��'b��� �k�Q%��ʙ4WrD���xuV��J���7�"_���*�1>F��]���i"�V׮������S\@�>C�w=���Ύ�Wf�d�d�� �I�q�s�+�T�|%z�-�-�K�M����X�z��ע�c;��V_�Ff���A'�~��CS�1��9[�mD�Cj	[xU،�� ��mc��A����_L��lԾ6L `r:"�g���<�&/5m�R�9�]o�)�[mR���i{Rl��r�HuƆTR���5ʼt'�S5ve=�$��-�绷
篨�3t��sʗ��6x5c����O�_`2��}c�y�m�g��N����%v���|�r���.�ċ��|�}��x�N������/�6�/�u$�#ɂ���&�ub)�^ō��7,hčY{iQTU�z�i�T�z"Z�L�Y�t�+3�0�x�,��Tuu.�:۽n�2��}�]fjO+
�6�̅����zv{RR�N���u�o��Ɇ��|���U��UK�#������M�]N�g���^����2'f���2��ޗp��C��/]�L:���Ӝĳ��k��vEGޞ����V��ojW���a�����}އ*3R�w���,͗�x�6hοS�/_����Va�-Q�̏;���SK�	����#�N(�J�*6�uG=�rPt�e�������0S��?�|����a/������tgW�L���%mdXzw���A�����5���O�[���͒�a��t+·]�?�Xx"|+I���
/6{��r=Y�k�iߋ�+�xL2���]���g ��Mo�$m�"nG�%�۹�ՂB���l��~���c^��.���;R{NN4̔O)����Î�8 >�^�����U|�����j�O|���76��w1gJ1�K%��G1��f��U��A���p4��tIr��&�t!t����~;ʜv)(wSH3����~��8{{�I2�ò+��"=��\�~)�@�[Diּ�T������<*���^����>RPy+�h�K�"���}G���f��ݷX�n3�#?L�+P��~2w��Q]�#��+�,y�k�^����{ʰ� ���[x:c����Q&��a������s'����I�/	n��˰��J�f�Յ��6J�thZ�Y�v����cypmy;�4?�]J��\��l��������cR>�Ӫπ�v!ڌ�͎��{+z��/��Wx)|{�ޯ��B�J��,���'|1۱V9S��!=BR�i-7�1l3ޏ��e�����/�]�=���0��_G�pP��h�NXDqims�Cz�T�Qs��1�,��}����[׺�^Їo6�#ܮ�$�����*��9V4�C�|�mӜb }l�|ش6����j|�'Ά��dv��{ܵ�&R�vov�Z��8�0{��v��O"l�嘍 ��>|3�^�b����ۖ�K�>����Qvvtr��MW�A���g�鹎�Cp�g���:Q[������'��3*l�/bN�~��s�:J�l��=�9���?	� S��e�x��g��sGò�
�'NB�<��f��7��7[듩='�k�Ȟ��|�v[D��amON�Qݿa���2;�ݒ�ҳ���y�һ��q{6�˦�t4ګkRo ��f���Kͽ}���ve�O�G���z�KVpp_	�n��B[���o����u(Ʃ�I�2eǌݏ=�=�;	�@�go��^ۆ{�M��g9d���jﭰ�#�h�?}����P�B:�����,��s��#;k�7o�T��<��&��d���*����.}��F��B��,��&羾��ۺ�nj�y�����y�o)�~y9������9�{���wө0��ko��y3��5��p�6_�++��ה{_���N9��X�݀l��u#zE�^���z+�p>���w��v1��)����$�72-�%A�|j}����$%����
�P�Yu��p�v1���~N3�,f�,I�����Q{--͂�Ջ���z���R�b��߆󗱬o�t���l��Lu�.�����׶W�禎��`O��M�ǽI�U��M��5͞��F̙���k'yg�v�J����?o���{y}�-����S�����w�����5�l�W���e����(�V�ny#�y��nX�ҽ}a��W���rċ��z1�i�@Sk����I�л3�X7��`��G����Ȩ��M�ʻaܴ?ug�J>�!�S�n��%~R=��
���;�v�����J��q��L��<�5c=�w�xX��=<�k/3#�M��}��w����P='�v�;ʿ��+�Sܟ���ă������e,(o�VיM?U��ɟg��e)�ϑ�{���+ޞ�U=���5iZ��43G�Ύ�x�~�>�V"����v6{�܆��[z-o���f�S�5��/�om9�{,)�o(�k���!��ɴ�v,�
P�ݽ]N�y��T���^�,�p��Ҿ+Z3�V�]��v��8Dۆ5kks��u��>���N���|�{mvd�|�@�v)n���s����!�������ǫ���ꚅ���~Q�Ir�6��P��P'����S��Z���8���{����	Jʊ9��#��qι���7`�z��|��*�.�a:�j��d	�{8��z<�μs��'w��ӷ$�72-��wXK�~��v=۝˫ҏ,P����:��g_Lϯ���-���^�ݳ�rϑ@�.���,Ǹ��|�7�eY��}QQ�p4:�`��)�3j{���u}L���_h�N;�tܫd��k��N��q^��GH����_7�I��e:����\�d�!G�\�����s��8Q���,ˈ�t�{.����
���p�s��ﾯ��f7S�������[��T/�li�	ΫϷp�2r͞T;�����z[{������V�e�C�t�s;Et���OeX�>�\���sϦ�p�\�PW�nmu��W�_�A��xW�<�gk����&xxma3W�����S�[^��zS�}�λ��}�R@s~�cf#_���]����ѡ�n3����j)?_/mg%�d��UNy�Z}<<�z�����-��y�'4}^��`,	���'��A��S��n_O|�M>��u���c�g�2_Ew��߾�����c�W����w��[==/ n�/l�d=��'2e�M����M�Y�e��������;�,���e�9ۧo�aW�9|7P�ܐ+���?yt�B�M�q��J�6��W���v�X����;gڥ�Ra�<=�z���qh�z��sIcx�Ģw� ����N7�������
��K�o;w�2���+`�xk�6 e�Vl���o���L[ul\�1��W�zf=B�ۡ����^�fV�5�k�62T��h��4�_��F��-�S���7�K��|,w9���`Y��{1�[���諭����gȂ�Y�w_¶�X���|"�<&������{e��Z ��9{�%���ua��W>��Ro������jng�A�dgc'_u�@�û���L�A&z�o�S�I�[���߆;��9�ԝ���y}��٪91-ʼ�g�m�IMSE�}�_(P	�6uǘή�0��G�N���m�X+�^���½ھG<)$r���u��W�I�Քw�ϫzV��&Br��O�s'/h���E8����Mxrkl�_��=\����4�`����,�ꂼ����K�N���2��-7�7Q�����_��*K�I�g�d{~�o�s$�����l��<j��]�[J�Sм]�%�"y����3s�n.~���i��w�Yx���U����<�ag�bn�dm����P{]�t����*�;�_>d���j��L֚	������8{Z����B5��3 W�R�o���m~X�'�[�v��Gv���S5���Qu�jawb��ӊ��K�y��;���#��n��FgZA������5�
Y�=F$����w�XVq�rAQ��>���N7'����΢��iyh��c��I#�C�>Q�p
x�E$����vܬS�a9b9�Y��F�g:]dQ��i���]� -k��>�#f�;TÎ����<�������A0��u�5:����� ��)>۫� S�����E2�����ih8r?{ܟ=�V{5tm�+b�59�ۭ�����`�z��9u#7�a�Y��E�5�ZxI';�º�mc��x&x�֔���(e�l�F�+u���8�i4�}Vb�7D��Ժ��հiΦ>u�ga����t�Z�u����=g��S����Gy��f*���,��K����Ns-�9�G+�z�-�C�D;���".�m8/)����VNZy�@�ݪ�Y��w�Ң%R�䋠 ��w�^�
�c�t�w����m�*�n��S�~ph* �`��z̪AkVi=��8��%�Ev掜�㱒��
}�b��h�Cw�1���P��[��Ĺ��e�̚���L����=yp���%��|m��V�a�)ӭ},i���S!<�"���t�u�4�l�m#aրw5cvݔh�M�f�q>�U�������j��p���u�ހ��V�f�jP֞l�HWj�xB�9+��ʍ���'۽\ێٵ3�����צ�=��J/W����#pzDm�
�ߣ����\E]g0N�f���!��Q��	2Nކ�����*�=�7i)��9p%�WS���ǖ���(`���f��P�7�c��dX����|�bK�v�AĻ�FJ���Ջ+��;4�5��qJ�� V8�R;ݹg(�/���'���N�Ń�%k��ˆ���dP���y�#mK�~�{}��r���bW8�g��ڹvp!��5A���8��	�����M6/&� ��u����Õ,VC�muJtèFZ��g�dv�}��Y�J�ǚ����1Ov�N���8�ኋ����{�tu#����Z	�"�4o�jО�1P��pt�s�y���tN���n\ȩ1C+Q�D�B�Q B�%v��MZخ�Y�ýN��S�A��1_!��.@���MxA�;9� ߝ��s��M��û<�
f�z7q��'wq�gs�&Y�����q��2���*� WIsa�{��uW�&���/"�b���{Dz�6�a�u���ot%w&/e�˼�S�:�o�
�w(9NrY1iFm(6	v�ru�/���H�5�2���eVL�F�|�C�I>s}�=Ϻ�Am	��(
�������,B\:�j4\S#����hPV��H𡙑_'\�,~U��[���gu�`����f���L�GI��.UUCi�Cm�9��1y)Dڱ�i��ʹ2䭑r��Y�6ņ�66�]�8�)2h��Dm2�m��h�h�	�^n'4�2lF���f�Ɉsj�"6�ڈ�1Bm�h����M	�M�sD^��i�!J\��la�6�afH��6q/%q����3�նN9\���6E�i[\fT�i�6��ɶ-�Ƌh�ؚ�d����TD�"ɴ�4d�ML�Úd�F�#kBf�ؙ8��rm$d�L�H�b��]�Dd9�r�9��4a2I���&Fi�q�ٶ�UI�q�M�E����¹�K61�rl�M6�f\'��_
D�����t�����N��"U�'f^�U􃦦(�ڕH�����=y7��v��,�7�Q�oz�v%�l8�H��:�������S��mO�����{���s̷Ă�ɾ���p��`g��#�A�)���A����ի�ӳ;޵�~����z9�"B�֖�8�6&��C��/��:"��S�u�KGE}N.������y�Ή��O�!��J�Vz�ڕ��;�������:�a��]x�*rY�Iu�+V��P�����Y�y��%�)v��RP+��Juְ]�nޙ=�M1���λ��m��;7z��J�˃y�#n5���ީ=��huuuQ�R3k�[|�	�i���=�@����M�(��4�g�!��ol��N>�����={[�s��<��N9�=!�Sv�C��"A�>x�Q���#� ��gq�n�`/:���#~{^ɸzd[	QSE�OW�|v��I��C�5~����.Ϋ�VΛ�|^;�e��7���`f��|�j�5|�%D�����?�P�ڴ��Eɑ����x�

�#�j`Xuk���뢺�c,ʏp1�;H�*��Y���x#|w"��=/����Z�v踸qb_'�m��e��Ś�n,x�:�=F_O�6zZ7O��y�l�>�����Ң�A/����w�`%b������{��WI8�W}�Oy5R��gnOr���3�2�i2��*��ǲћ�w�}���5�:����f�����Q.-z�l*�r����f#��=�g����V=��Z+/7��e���V�2����+{���Fܙw��l=@���sK��у/�h��:�8��y�n_`��{��z|g��w��s���8��WY1�S�F���@ޜ���N�{�y���S�g��uSZϤ����}�z�U�|kf���s���Iϣ9�_��`W�/�N��������>���^W�m��n��G�� ��.~�{U�����Û��k����C��a���������0�}�z&k�ad-�뷔'�ƴg`�`��!�/�Xi���{����Ɯ6�y�:S�k8v�u�d�|�@Ρ=��=a� �Q��W�0r��Z��G��^�����h]K犲�����7���X�����ɽ�6mׇzu4_��zzaĄwF�$�j�ǖ칛��@/��1��t+3B�a׸�w4�[=�F�F�q��4�k{��#�ۛ�;yQ�+���=�ֳ�c�����]X�&�N1�@�Ďo��{�	���Z�)�\�>�}8�{����Ü�ϭٗ.m_�9��#��qο�r����:���qٝ�&�b=�u&2i���y���r�zv]{ہj�#8�͊~۱�
,��V�*���7@oH����X��,s��g���mE�{N��^9�[�ܚ.z&K�4��t��꿫�n�<�W��.�9Im�xj^ڸ6t�rq��!��g��+�|q�;�Cb=�\����O
�F��Ő���9x���g4��uՈ�*Đlw��������9 �s�H�k�'R�K�ټ�R�vVu__�ʦ��q���s�b.V���mN��ǳbt�狇�Y�ۨ��O?D瞵��{=9���������Pzw�������zCxZ�7��3۟#�.^��e����҃r �2z�F�}7�:��r���Z,`�U��ސ觌n��RV����DR�J��4�����x����א�Z�[�&o\�Y(/.StPܑ<�|t�Ì��ǲq{V]���,�C�uf	Ӌ;IvjN���&�F<��GD'�oAQ�W�k�m/�ʅ|n�X�߾9��\K�q_P���P%��Cs'E����nN8O/L��k<�{ܜ�y�ZB��U9aͬ�)�c��ɓ��nK��g��բ���l���}Q��پ��m(C�\��[�W��n_�x^N�<�A�N|)y�o�5K~�70ǒI������2%Q<�/bƼ������߰�k`)�ҝu����j�=4Ǟ {	��E�Շ��w���5.���۠)=�޸�ݷ[At�H�V�B켡\�k��u���W�}$Ֆ7`���h����wt�w�w��̛�佗��>~�ރ�i�8קk��ސ�)�h�ﻨ(RoM�q��i�������
�����..�o!��8�>�#�P��bȤ�����y��8�>s�Q睐%����F�S��Xˇ�>ڮ����`��H�-��l4/.a�aW+����(�T^T�ӛ��.ʘ�{�!�&��[j�h�8�l�ʵ�i�uPF7ajCr�=z�fu�0mJM�l�L�n`8ξ�ҳg
� �q���RoC!7�k���A�x�k�?���BWW���7M��~9C��ge�9��oj��`�d��.��My�n����#!��u�[u54�)��5�s'������ٕ�hӒ���)�Z��{>�.Ø�7����u�S2�s�T�6�f����X+���w�M5j9(�_Z�9rʯ�Y�Cr����ק����/vqU����z��^�0�\�5t�}��=�A}d������n����ߧd�J��	N��+D�(^N���9
�;�Iy��v�缲��+@��j�[y7w�M�����)Yb�������܅G3��پoz�����U�[���T�R�/K��:��u��ң�R\��\���n��'�	N�������^}j�����s�Jr���;�ɤ�&�YB<��s��,�{m���Ts|��f�s'p� �v)7</��'z�{���ޘ�4�k������짮mG�׼Fr�"�W��{kNn׮�mV��̗�Y�98�o7�9����=8�x	��+2+�O� ��=B��l�������2��Vn\�f�L�Sv�9�%�eܠ�f�)�m��o9�� }//�����������X�}�@�g<��v������uV��������]�p�*��t�;�V���<��N9ސ�~���l�ﻯ�{̿fUf=����ǧ��4.���`/;�2wH��rN�2,�Qw_7Ƭ߶^�N�
p�#����	]�S��#����}����\#�+ڴR&������5H5�f6������@�Ob���ʸ��Q����O[�U�V�\_�p����_��Ѹ��#*u���~�n��9���Z���t^��f-*��TF����IF+�)��U:�u���"^�J�ƍ��Nܚ'E�)�v��ϣ�`k�?|ܾ�8"��޶��Y���,�S��7����V,ǰT�]4��/�����*v86s���k�e�]!��Tj��d��.�қ�ЧW�^Ų�f�zm�Sxg1��s��ԛ9���vsz�|��ۈW�u(q
b��l{�$��Pâ���ٸ�A3^�d�@ߜg�_����t�v��xؾ�xR�uraR-f�8I�]{�ك�:&�nT&M�l�:2��x~ܒX����3��feGSr��}��؉n��l>���Q����}_���W���v�v���C�};j�Y`Rp����v6luG!�F�z�W�M���{.[��z�}qm5{�.��#�ڠ{����V{�ɵ�;��I��E����虯)����z��	��k�<��`�<���ٕ�8��{�`�70Ǟ��;���{]�]v��La�h쓕�6��G7Ύ1��/7�~1Ӫ�5ɾq�<2�9���v�����e��G��%W��������vd���(�G���8�X��%�vm����j����Pr�n?�0YoM���y׎r2wt^���]v`��M�Ös���m�**]�t(�{o�����ڥ�+�6���R�9��}I�9�^�!��h�=�� �u;4;�6�tn][aS�ޡ��JmJ7�Yܽ�*��q���`��C���wU���M����]�����_�$�,ݹP��-������~*�����`�^�9c��չ�(^w�j�I�թ��`������n��>�Hkk(�zlV_�/)�(�_����ln�	Z���J�Â����ܕ����4�I@q3s;���L=-��?���gbYҨm]nK�Y�yݕ������p� ��5�[<�s;�9L���f+��=�ʧ� �$�|r����z�(���7.���� ;c�Xݙ�l��������$�Es>���Sk<����9�7/Ӣ��c�.#R����7��+�/�;�����z޶\���1w��S��G��s���WǛ�nN�_k͓���U�K;����י
��k�s�~ꛟT�cMN��i�U)�Ȧ�+���׳:C�������z��ye�:�O�
����;kR�&�m���)`{�Pp�N��*9��f�Mw�w����׻x�ox����e�Io�X��V?Wq�%�Ry�$��S��^��~�{ܼ���<�tt�9*��2��@��K��m����o�T��4Ǟd_��Jb�=�|��K��mbN�=���*z�Ra9��WQ��ڰ��Nw������A7o��A�U��aKc�'7Ml�KHL�^��rR�&��QK/obz�.W�w����1�����h^P���h��nBp��D�sq��%��$,��N��Ej�.��f2�:�_'���%Y��1��7�qN�����v�]��#LNf��^&�+1�Qؽ��:{��g��ؘ@��m��p�y��N�j�nI�u�u`+�^�{R�6����<x��t!G����sdg� /����Z�C��v���~�/lyῤ�*�?G�Gp���7vgp�p��WhofS��0*~���d�ӣ��q��,e�,�y���k��[;P_��@��U��SQ7ە�˱qT����AXJ��tֳއP�Ɩ��HۯR�'j���|Whw���z��߆k��ITʹD�7�a;���]A-�=ޔ��8������y�֌��%���*s��Y��z.���,��G}�E~���9�`t�������sצ3������u��5û�zO
��W���W�r�]�F/_�����s-9��Ģ��ݛ����j
��Fs�:
��NB�=�^o����/��n�$��;o��5֕�sm����*pt�R׬�Á��P�!��}���Y�^�;�x(�_X�������뤾��T��^"�s��[,�A����^�w3/��d�d�yWP����nĝ�|�w�+\�a�c.�8�3o����R��A�=�yfR�w���v7�!u���~c�f���nb�xܮ�Y��#��#9���*v�����Wo�B�rYgLaA�*ī������{{eQ��܆����P3��/��_oԻ��F���O?Wv螽���$��������G�9���Fs�G�Ѭ�����a��!����V�i��|6� y=��/7`���wө1Y���P����#�\/�y���َ�{�s�����>�}�=!ț�e��f�Rz�k}���l5^�� ����w��/:���#~���M��d[��*z�ˁH�ha��g�0K��w�e[�'<�������7������%e{���篋�O5@5YM��^��s����L��/MX~}�ܛ&];����=�2��M/�����Or�W����k;�{w΍j�M�<����E:'d¶�d���&;��n\B��Ed����<�^��Zanf^<����_q�Rc�)��_U��;FJ�w�l�WM|��Z-8�f�-���x�^>��5���l���%Y+n�(
��+x�
���`�X��s�>�v^�ȣ�o.�(�1����A 	��#�ʉn �BO
�����3Yܝc�S�Z�68�I�h�Uթ;u��(':��u�1�&��j�3l����[�̶k^\k��.����N�$�~7nS��aݱdkVp��M��`�Ј���3�ܞ������H��ά�}\Y׆�ؤ�e�|��"���XԲ���& *%a;łћx�Y�����&-�f�Xo�v%I�u�Q����m��w�f�r���������ܔ��q�F��3//�k�+�� +�1��w�-��k�T�6����oo^�6���`۽.��z��Iҟ3�2��魾�Qr�5��t���j3��~�<I�LO�Ǻ���X�޾K쭷	�5M0�6���xEqw�⽙�d:G.�*��� �g����7"��5���;\Z���K�|� OGpR�o��Y��TU�[Xi��Cφo[�ُ^<ؒj�6e+u|i	|X�7+��$`Nt�9Z�XWlv`a�\�����mg]p��th'��i�>A��-c���묜���A����Mm*�˨�[SL!���u�c���<���G6����4H64<�w��wX}�^$j�9Y����)���:}��c{G.P���q���Y��ƙ�z&�zI�s싊]� �\t��bk���A��(n;÷zW=㌴Cs��u��^ڸ��@®3z>{C�7��|~��P�E;�Z������czP{$1X�ŕxx�J㻚��|�
�*��T�E�|�M�G{�UN�8��*������}wq[j��f������sM��C�X�<��k,o!F4E�pۗ֕K!�e�q���n�h�=E.n�=�\��y���h)���hu*���Օ�>ʓ����5f&�����pۛ�.pV����
̛͕�|�����"�����L�+7t��wx�ɤ[�2e�d�,�������{{ET��v�c��]Z�
�.��j��+R}���A˔C;B������w ��{�����ڵj��,&��}��I��O_`�][�p�4gO>V8�廕4��P����b�.pfdS;n�o4:�SźI�Uy�9k�b�}:fw�{�C6�u�Տo\�Q乒��s]����7[�pǆ��r�I>�����y�.6�xN����
�V^�F/U��P�kgU��JtGڳN,��7{u%u�+|�3b�d}�)���F(����yej$.?;�n��� ��%|BH$$��o�r��4%,�8�#$m1�١j�����i]�F9����a'4E��8���sNrs�k�Ӝ��ĎF�ږe�qsni�"p�m��i�E ɦYļDq.���.�"d2�6�ͮٓk��F��798�ƙ�6�L�$�Ba#jI�HW+6��#I��.]���aQ[Fi���#h�FƂ��h��&��61��r9�$8��r\Ќ�4\�H�	���M��324l��5�2f��@Y�ʻE�I�h	�1��k���&��3Cl�"�]��h�m��M�s����M�i�m[eC& �\�Ѧ�6�a1Q������n@˖F�teA��m5&\�,̔�ɦ�j&�Sf�3&Df�!fD�"sht�1xӌl��m4"bM�M#&A��ƓMy�4M"   �/b\T�Ĭ!����ds$Pk4_ooKA�ֽ�����H���>�k��N��E�b�#��̰��o�.ȭ��})N��K���]������N��bH6x5Ycf#_s=_=������^�LAy���3��>�M���]�V��W�������a�m����Yⷻݝ�R~����K~���O�{���M�pt{(�7/T�G�y���l~��:^Ի���)(�K�M�Og1�#���	:>��t��]�X�K�V"�5�4k�'�8�_�nB��Yuبju�Y�>ѱ���2�&������Bz��a��>�uZw��;}��Owf��w����.�7&Tog�;7�gP��e�d��n搜�9���αY���z��-�j���y$�+���U��|9�s�5��i���I��>�l��=���t�ɒq�2�#����gI4�ɣma�#ϛ�^���R���r.�@m��f\��c���>�������9� �4�F�]E<[�0��o�=�Z��݃��SF�G����*k�0�6����㋖������v�!�˳��l�\�+��[�g<�ַ�5k2*�;�һ�xw�fI��ϳ=����K�ի�|$����V>��r�p��.�m����B�ں���j��w�6]��b�zl�G�U|���Cޑz�˶K��t��0?Ax��^lv���Қd������}<��|��ZY�U�NP\��'��=�N���kpE�"�6$�/�=��4ݝ)9չYى���3����}>1���/�J�$�=C�t��������n�s����O̸�ʰ+����p��']\nI�5�[<�v�o���j�N}[���C|'����mܪY&�k��~~n]_�p5bH�}V��˳�㵢a�ާ&�5��m�ο�fnN~���k7���+$���eY����4w�1\O�&]�����`>�3�9X9Z?)�hf��`nl�_����������q�b�}���x��tF��QQ�������w�wC:���=Jts��9
��G�;5�3�Y}aw��Q�<�����.ua�q�� �Sa�ĥ-
}�,���z�P��9��������:�p\R�ř�����q�d�#Su��y�� b�V�ݩ[������e�ҝXo���e��o:�N�:�AC�k8^�^ؓr�5ǚ��r7l�������ʨ)֣����p�G!���S�ϼ�iBDZ�{�M����Jo�p������[Ⱦ����-�����Iީө���Զ�iK2��#%>��|N�n�\�u�[q?m���G�;�-�������8�N�:�Ǆ�]mٻѷ$צ��=О����w�&���̰��N-�U�u�{;���Y��ؙ�,:n�6z�}8���A��f�׼^H�b�N�P_�j;鳲��t^��$9�=!˔������P����o]b[�TV���A,�B���ܿ�<��^����"��TU�E�&��>�׋}�ѐ�9_�n|YK���gMG��_�:?���_�X�R�WyA^������(��co�l����oy�65.N���Yp����Z�����qW���x�h�S���:���#�)�����_�z�m���A�.\�K�Z��,C����C��z����]���R_��O�p��f
� &hލWr�s�l���U��\	��֐2y��,үȃt�:�	��ּ������I>^��.'^G�_t�I��{�v��<=Z}Z�L?"����}}���rr�Yv6b5��=�s�ṮK��Z���k�ڡ���w�,�?i�\�oܡ�U�/�YU��7X��@��<��6���{�c~���JV{���{NW.%Z�ڱP�Y��u�=ុ�cQ���8��߮�|^u��e�[xg1_^N�'!b������z�[P�,��~�h����J�ώaw�_5刱7�1;��zy!�+�Z�� F���!R��_!7R������ɣ�}a��{ }]ѕ�V}��d�7O|����Dm���~m�T����k0['OO��)�+X-tb�aG�v-�����(�V���;˰.�]إr�7�B���:*ގ(�[��/����b�;�\���uc[����� {L���g����.Qon�=�6���'���G^��s���<��qα�X��J��W��h����[����n_4+q�ܖ���y�|a��F�cV9�/�>�Äw��7�gxgn4M�.�e�+�y
6�zP�xs`�8.��3
��BR�����u��\��;���/z���`�K|٩h�ĝ�����^ă�`��s�껴�fkI�z�~��h&����������d�;%EO�P���1���&���:w��0�&�;Vz{�t~���0��^(�:v`ix�q��%Ł���|t���\�o��6(׻I�n��N��϶t�rq�2�k�\��NX;��*��z�Q���-���wpt{z��}#���Ы��VX1�=���g��SS�r\�.�+ �����c����ܾ�O�-�2�y\����Oۃs��uxo�g�I7Y�������mQz|g��w��w��s���4r��oէ;�/��v��!w�Oc�\�ޥ��o�rSI�J8��Y\vna�;חw���m"A�֖�8�U�p!*�޸��۵()qͱ��)��8�=l7%�\�^�8}�)���Ŵ8�7��A��x���-	���1���)��:��c���3+(�PҎ�ז��9�$A�/��u�Pqd�Ň��WE��W4�0��jl_)�c&�X�m��y�u��qD���3�ɒ� �5�b���E�)����2�s�C�}�Lf0ǫtk�^)�rn\���f�Еo]��O3��+���%h��Ѧ3)ϩyح�e��[�!�0ǞI�
�m���;מ���o'��7��L߁S������[g�����&����G4����g~�36�������1@�=ƾ9t���K�F9�=RUߘ���[Y4�f�<{�MY:n����4�����~s�侸d2ς�G��Y�n��Ѯ/8�[�\�uׁ�t�q����p��b��9�=%V����b8߾���9�$�'���u���t�MArn�}q�l�<�ݪSy����>��I�C�=>�|�ml̶��
�O��1�]W~/�������X��)�uՈ�7$<^	�^:�ܷ�<I6�q���N��o.m���O=?&����.�y�՞��R�S����gk��5ێu����һ����ud���� �d���ߴm=��&'�l���x����h�qY�VI�d^"�C˅K�_��6>�7��@�wu�ם��d
kH��O�a�w.�W��{0���l�vMfg9բ4P�B���v�V3V({��]g�r��!yS�Q澵2����s�Y�
�z��u�:�oӻ��\�{ޮ3�K�[c^�Bo:|g�P���ry�����{��� �O�sQR��,]��Ci?eB�7[s����-�[�r����V���Y��Ԟ�+��r5��Ϳ�f��ye봎ז��*�{�w{ZJ��v�gb�)A���N��Q��پ�M�>�2��[967�UY�\��	��+iI�k��U���x���=�V�<g�=�:^�q!7�����v���`���wo=䇞���#"���/	�-�{rN��y�l�2|�7�R������6�8�N�����5��F#܁�3���vl��u���wE�3-^cl�<1U�����w:�):;����_ސ�O�]�p�r�5<�M�C�S��[X��O�g+
��̪ynօ��8D^��E�Y�H�˗�WE���|;�9�H�km�#,|ލؐ���k�A��KWݵ��'��㖏_I����r�9jb+ٴ�x�
5����+�--5f<���I�qAP�u��ɑeK�~�g�Tj�����ۗywZ7��,�ە�vR��~bv��j���~G��/�E�5��=�~��u��Z+B�2�h�8Oe����u�!�Ef��v�5�A��^ʿ��m�8�5_7������w��T��������6{�*�nܴlOW��kj��Zj>hd���D����b�}u�twW������t��[~3s�;�da���3��ҿo�>�*q���W�ʶ����ܮ{��d�\v\�y���	0���}^��ꙗ]4�\�m��S=�;�r�wj�pZ��e��!ꡏde��E�[(�PW2�Fs��Wד��TfL��Iy���N���-V�a?zu�S�uH����ܪ;����R>��=Ko�=[�#���r�+	�m�;��Y�{�����w��Օ�b�j������R�dy�Q�.J�\�K�v�c�(}����+�,F.P���Z�Kq�x
9w��]ɽr���g}�d�b��6�i8~/���ջ^�8v��ۧF���%]���2�l�}�C�c�{I�'V�!݈p����c����7�(!�нҝ6�n�޳|��#��;e�e�h�N����%5w��4�73��z�����8L1��I���os��d�|����O��]=�ػ/R�`3q��f��;��~��D������g�Ot����v���Uc2'����;�܊mj�g�y`�s��A፛ۢ���Y!��PrΆϫ��򈷤oG�����_�N��ۮϩ$�j�`c�����"������}`O=��yW)t/;F�<������'t�jt��c7$�bz*��X�}�����7y���+��ٷ��"�������5�KB�	b�Q��w�P����#���L��r]Z��K�e�olk�����>�INf�G�W�g�L��np��]?z �I��	�X�9/u�k�m���V�lI�����^�쓼����o�1���t�eo A�:&��F���AA&w���D����Q�>�ީ eDg��9D�x���(=������}'k�ڭg�h4�nt�������Zs+[ڲ��n��煉��;�Y)�E�x85wYoc7�Ţ���#��g��2�c���H�W2�[�Jny-���>�|^�Ҧ�c�v�+�'r�����Z�?�F��|�~�H;JZϮ{*��|�Cf|���O`MO?<�+m�mΜt�A���y�i����$�ih���X'���+�x{���F�L�5�B	ݬ�!`T���G�w��a��
�g:�7�S�o.�>�����b��G'�I�9��2�[[^{ܓ���{�I�[�|)>[߱�~��a��$������dپ�#���<�Ҭ�}l�I��u����u��'�i�=�=}���*]oo�8}�����2��t�ϱdm�f\��j9�oQ�y����]&%޽��}bg,i� �ߦ�.�C`�G�FpFx>���j����V;V��=�\�;rL�d[`Ji����)wa��s�^���z��e�\�c���$.<#���˦gU�Pk��=�1M�ٴ#o�t��Eu]����2v)On�C̄[K�8�Q�UC���i�4P`�2Ͷf|�v�p���^���E�� �6��kE^�Pԗ{ܩK ����NA)�y���_f�Zِm�n�rG&��Mo����}k�¶�"�`�k,�ٸ��ӀYյ�|�u��13퇪Q�:1wd�+n
��e��yӂuCl�0��8_{wDnE7�PE}H!�l��=��y��h}�vz�a�3���dxa�ݒ(�T&p�q�r�e�2pT^���u�YG��V�_���9����ǆC�T�n�6�Ζ{�w�Bdׇ�f��w��^K�o����(]9յ��s"g��-���Х���W|�Yx3�Ç��������sj��1�x�m-��pّ�g[�=�=6�44:<bf���hl��Έ @�ZV$���\5��������M���4E�'�ZɔZ'g�	���SbCt�+W��o��i��5.,ݥ�B��v���C*�!0�r����ǳ����ކjq.�8we��MLwP+j7v��b�����P���fS��v��θ�чd)��4�
�6���} ����;B.ms�����GO�X�{�w��da�2�R��c���,�R��L����H��"SX�.V��祥MG�>�[T3�Zk��J�Nzi`Żr��.�����*.��B��9	�h�Y�,�W3�k�*�̤�m��9���:��׽�����;Fl(���6�#�L/W�!=a�8o��8ڦ�9�:��H�}��{T�g��]�|�]˶ͽ��]�W�nQk�U�>�.��V.Q]Y�
�T���pz��wS��Ѹ/�Rzӛl+8v��X�z�	D���r��6+�!G�K�ڟRj�E�:�rʵ����ԂS�jnA����x:��\*M4Ѐ�����ঠ��ޒ���M���y.]����1���
w���	-���o1g��]�.��w0_J�h#��[�&�.p�4]����1�MdFR����+5I�=1m�O63a�r��M�C"X_oQ��yLt��on�Z��0"2ʗ˒��m�g']<��l��r����b��������5�q�5������gDCyR+e	Cv�`q�'O!��91�^N�m�q�.j��n�N��	���Rk/_}4�KeVN��Tr��}�PP�!�r�≢�Ƽ�9�5����\z5Ծ����2J��o锝���B +"�	ق��#��XB�����7άs�c�8Ү�7R{�A�q>�F�){�-���*-��v�$ł����u6�.p�l��;p!:�a㷘3���}g��{�P�v�\�v�������]@�}e1ͼ�r!	�9���,�v�8v̝w�-�qa����r��f��?~믿�߾s�M8�Au�!mL�V��i�$Lē4$6m[]3&� �i4��)!U�l��"�2254�i�h�s��l���HY��6�Z��,3cL&]��fFͩ����f�m���ٴ]�Fڳ]�4M�3F�m�]͡#��&�dM��&�m3mf��54�U2k2l�u�f���BC6M.�s�9��%i�Y��DBf�d�6i�)3M�k	r5�I��m���Y�f�3M�6B��'&��ճm�D6��	���4H�v�fa�m4m6B�5ړk����s5hF�6�3f4+.���m�6�d�4Mr��LMuѓmuQ�B!26�cH���r�5�Y��5�l��lmi��3ff�4CPhč�漜Cd�s��\*��Z&M�!�b]�F�L�З)6�4��Hɀ�Zd�a2@L�	���2���͈�k�&fF�c$�!4�&F��/'��߾r�#s���Կ���z�-/ݜ0=�y�5�td*]Og*�";E
�->ȑZ�m�H�e���L'9u�gn�}�k�2������_8ߢ���n�l����ܯg���~&���+��a�?*��:G�NYc�K�I�{�2�"�A���v����W�C�U��Hv��+]>+����l����VoK�uV��7$.�x{�ח&����c�1�X�Z0^�98��H������ ��?*���-ͤ�+2����]A-�=ޔ�����2�=��ʡ�v���_9�G����%��N���(|	�ON�{��m����F*z���>�33c~��t��2�[d�.79ɹNpN��9���='�|n�.�;�2p�ۃ�8F@3��m��PS���)���AC�i9�����mf���K{&.�J>��rΒ����p+G�X�Yb������c������}���zr�W/:�Ȍ��Rų�jz���9�Z�~�Uu�&͵�ۧ�nv��q�@�֪,�+ۃW`�{hڶ���lb_����2��V�}l��'W{���n'65���(IqIϕlч���}/pŅ>���Cw��yţ������x�a��u[���'�3�B�WЂsT�s������z�B9���dP�NR�Eo_ԧ]l/�7k��9F�f����Y�;myvR\���lH��0u
�9�`���p\h͌b���Y��:�'_*}&{�=��ۙ�`?7`=_w�`��父�t�t�޽��_���4����uXRu��;d>���N��U�;��㠮��9Ɲ>���*��:�^wݳ��8ߢ��3�d�j�X�w�ma�o���<k�(��|����k~���_v|y����>��R�!������6&z��\��&��+���U�N�O�w���	x�ǲ����7��+�UZ��l��xW��Cx�=<�=���[��ԧOi�	^�q
����#������g����tg��X3���^��Ƚ�C��}OJg՝��?-\���=�ޯS�1����1熋YmQ HJ�E�ײe^T�'�����̼ܚ�ó"-,O�B^�[�� �����|nR8��I���\��w�9�xw�y��V,�����җ�"��(؈S*��т�Kx�jQ���"cIL�W�&���������t� K���4��G&S�ǚ�{�9ݱa'6��X�zwu�ʐt������=bn��Cs�+{���GKܓ���2ḁo,�s��Wד�����I����w����;u�&t!������d���P��7!~�!Ցw]�M���ǧ�2?o����E�����P��o���+:�J���u���S�ܝ�k}��^S�����N��{k��,�N��
a�&{ݲ��N�fMJǋ�A�-�RX�a��I���opu��:��~d���Q�u�����������j��݂7�_�s�m��3��va*�k��W�Lv�tρ��n�J�4{����-F���oQU���nx�����{ 6z���A4zl��)��ҽ�S&V�A���A�;���^k{����Q\�V��_R���0�,.}���M&o��m7�7�pt��g��q���G81+������F���W�YYв�72�);@�k�u_<8�[�'�D����;�+��<x�&%�T�����łq���d��j��]��.:�y�³0��t�U���q����ڦ�Ƕ�h����[$>gd�,OEM�Wp�zJ��R��mf���N^������N�$�x�k¾v�}���j���Q�iװ>�y��ʁI�W���oM��KuՈ�bH6y���F��>씴L�ƾ%p���Z��0r\���쨌��Xn]��ՇZf-���4�o)�.�wZ��X��Ϧ���76�gX��b�&���U�j��+7��P޾��T��G�տ{�c�����|-P�!'5=��nѥ<)
��xt>�5���	����{;fs��v^=����tz*��TZ��!�z5�u�� ��,�^���r6t�7�6�gլ̿���+�V���^���Ay��g�=������;�=��V{�g9�yL,�]q�����[�26�U�eE��+z�'��k��~�!�0ǞI��vݺ��}�PD�du"{w��5Rʿ��Wv{��hm-�����o+���}̿}}��5�I����w�{l�0���^�b��0Vi��-L�����1[�����>ma����W�15l��ĭ���{��{��:��	�&IǾF���':�guG�`�����/��M�s�]�[g�u��2{���<0��x��_���s]3�y�?�=О��@�v+i�N��2�Vn��V��!n�q�%t�qz���g����zl��u&n��ۨ�Zy��rUޞ����:&��i_[��[��^�"k>h����S+V� �׳O1n���7��ΰ1�o�q�}���-�rE�%EM	�!�w<�_�o�W�����]�K�L�����:t~N2Y������=`5���S�g%��A���_���MM��\f���%�=�æȧZ\@�cJOv��,��@a���ju�>�v�{fx��`����ƹ����^};:�Qj��r�e��!yS�(�Uh��V.~��0P^{S�m�{�r���S���r�?K9c�7��O�E�w4��vz�4(O�YTfq��G�wU� ���vԭi�X�����W�K��5�I.�=�t����\��������v1���,��'��2W4H-挅�[y�Z�B�!�-z�pcq��C����b�Gv�»)����;N����n*/-����u���fw����뗹ny:���P��?e|��֡�u�����ಣ��8㵗뼀��V#����g��'!S;`��|'otϧ^Q�&�V�}*��+��e��@��z��&'{�LWcqyې��t�6�~�����1���1eϱ�ε�p�XO���J�7ګ�ɲDɮ=�o�18�1���\�V^ڊ]�V��{]�Y['it�3���3ܴ�6:����'\���yz�9�zc�d��s���9���d�s�])U������Fg�J���S_gs�P��Q�|�;��W�2�ޚPծ;�"����W�@^r���u���U�'g��#��qΫHz��l�㳼/���J\Gp�#{����ޏ0��go���E훂N��%�8���kj�S޹���L��|j}|t��^�}4?>�e��6~ �1��,�~��ٯ7����5n�jZ�v�,�_f�\�"�`�꺳2S1L���b�h����]9�Nw;<-IZ�}3H�Yy��.�*;�a���T��{ݺt�O
�c��6�d���e����#�u���U�y{B]Zya�~�����.E�mɢ��T�k�{�ئ�{r�ya���� ��M�fu�7˝�:U���<�g�k�J����:ǲ�n�x�Xx���+��F���;o���t�X��j�g���������^T>Pp>nn��W12�ed��`Vv��k�]��7/������������I�ϙ�
�-^���OMy���za;�X6�{��V����^ۼz9��G�:�f��z�n�M?V,��w��
:�A���|Pd��f9P��
�OMԪ�s�ր�S
e׸��6���z�����~U����ո�zx��k�����Jv�O����ן`�?{�v\n���d8�]&\ǖN���膶�\gO����'�����t��>�Y�xzM�?<JT{�/ W��g�`r��jS/i�6yE>������h�82-I'I�Ȼ��#�V���{m��/΂qS>S�oP.q9��4�`��������C�3�<6��<.���Pg.��5t��iq�d-�}%��*�MX)��7��;tZR9¹a.�M�:�u�>�WS�c��
����f3��@e�u�r����}�%��oI��)�Ҏ
�zn�۬�糬I����rֹ̀�i��uܚ?u&q�ݼp�e�v�
�� ˈ3�H>G��R�����)M	ϵ;cG������A�m\=���>O�У��au�Ѯt�?���H�K�`�*OwO���.�v���Ĵ��k)��7����^UK��T����'ZT����qW�a@��i7���V`U��>����H�qs��mFM��h?�O����:᤼s#��L�5@	M|\�1�h7eqyuӻ����G}ýǜZ]
E[����1�;H��3�-�s���6�@��>fj�+��jR#I{d�P-.�3qʱ�u�EOOa����>3��������Y�s��P��"�8����~�^�n}�7���Xp��^���4'�{��ԴާR�}wF-��ɿ��Z�1^u��u9;��9����2K�T=1���}��جT�ߣv�ۍWx�$��_���A�:6c��^e7���[�&��{���(���[0�lS��uҴ�Ϸ����a�q���}w��j�qU��7A�c���<���H��r�f�9�
����ƥa8rx!���CF�%�ˑ�*����v�c}]�Ii���Eй8*	w~���u��A��l�V��v�v{�q�ha9��B���J�B.\����`�r�b��xӣ&P��̚,9�RJ��Q�Wm���ɦ}���g;|�v�Wl����uǺ{:�ߟ��wև�U~�~�S�Ξ;Bz#.}�~��3�g�k��0���@�E�}c.��JMy�2Ox�/&\
�Ʈ�T�e��S�g�ڸ��Vi����g2|}������GK�rjFz�ލbe���U�K��>��`u�l�I��l�R��B�����p��}��|L��40�N ��t�u2��j����V��`��x!����?z��mD��4w����r���u�7�*;}R�I�3	��=H]L�ښ�#uʿߋ���"K!�^�s��w��
�ۈn�������D�︢OQ�P'���_ճI���+�k���险�'��]�W�Q����%��=��y�#�A�z�� �j$�!)`��g4_���SQ�����f�걈�"�뉸����3�{NCrp���r1�FqL��@z.�ʐ�#�}������!�ҭ�N�c2��b���%;Hǡ϶�9��&�w�Ꙑc%�N6��CZ��*�(��SQ�G���B�W3��c둗ϭ�<���|�q���iں������1��Z˥�;3Od*X�y.�cR��Ku{i���fC��(�_��o�|��N�J�e,3�J�	_�R�A��/��2t��#��T ����?d��o!����47���,D��.��޺v����X�^����n�x���J��9�x���&a��N��D��F�+�o�ԃ�j�1p�]ГUz��"�F\bZ�9�?�<�3q���}(��d-7����[�~�����d�㢽�*������xG5WG��
z���r�^���'��|���g�N�po �ΰ_��*+TK�7��zo����{����:���~�W�}{(4}(������g�vY_����Jß��zN�ҙQ�j�eፆ�V��5����曆|������+*=���q��%O?�gC�8EO�ษt��gR��1�T��9�:�{�Ռڂ���kQ�����<��{�xû�g�C(��a_�O�(]zkԪ�����ZfB��8�Y�����'r6��o�Hf�7���;.�Y��|�1XU�'���mx_K&L�T#�z����gin�\j꛺d6���ȷL5�w��7:3��T���D�5'��=P���&���� <��{@q�r���+��F�O��eg��}>�j��O�G@a<뗁'Z^���c�'s�M��X&��w����h�d�t�(J#��u���`qB��w
V��#�{;e9���]�=x���Me��CщI���d��qU$|f����	k6n'�nd� �#���hI�\cz��_�)X-��Q�z):@&��J�+a����ĝ��S����/�����ȗK�,j?>���U�X��u �кI�)���O����;��x[b���b�\p/M�A+|�׼����qN�ԭM�l�z�-��=On���&��i�O]8�����xgX�Lb�a\�e�b�P�V
�C�%��.�:67S	R��z���q^�-�8�b5O�H�R��M�Rjp�˶X�E��ظn:�RV��Q.-�1uds�ѝ����BXe+x7B�<7
��Y
z�.�;�-�Ce��,���gWL��i����x�/8!2k�6qv �椱�^�������&������6���{.�U�X��R7�&�㝜�6�L��c�"y�o(莣�޻�fao�Q�d'p��@�E�n@�;Id�yD\&Yg6L�����Y��w�	/S?�7i67����t�' y��q$x�J��"�S�^�!{szPEm1ܧL�`D������ͬ;o��89���y�D�%vѶv�4ݔ{xT�)W��a���X��kr�<gg9��[�Pf۰�	�Ǳ����>|L���I�m�LV�Q�&ㄌ����v��Л�[W{������=:���°)�M��k�����#8\��+O��Ӏ�ˉc�7˳��GpZY��*^�*�$�Ĭ�sq�C9n��G��5�3����2���w�bȨH�Aۅ�c��
�SJm5F�>]ZL�rvlIS�v�J�� *٭1̥I�J��u�=���������l��R5z �݋����n�Mu��V!�]��y8᪏c}F��%`���rXM� :� �o�=�d������?�
�n��

���=�T�IOm�����\�	�˖�eű|���PT�p�{b>�L%�{�'�7v*c�ݏw�WE,v�-GVK(k�5��Y���8 ��1[��������m�i����ޞ�>^�ВM3O�(p�ެfI9���/B����� �թp,c�,Ӻ��e)��t�Xv��6t~ۣɱ~<_$��ޟo�i��'6r�����r�x�"kM���j�VZ̡:$��� t�9v��=/l˛�_iT�IJ:�L�!w�f47.�O���V+���x4�|���q�B�3���&ӣ�J����Nn�ȗ$3=%����b��k��P���O�4�N�zM�.����[�sz�*p/UA�h��|��Y��8��k��\�d�u��X��bwm:�{w���a*�Z6�����2{xJ�U������]�k�Z�@Zc�g/e2�N�%͝l�Wۘ��޽1�s�;����|8���TO�2M#f�FL�eMqck"�!Y��K�$D���ƩL�Sh�	��E9��R��X�#dX$,a	Y��bm���m�m������m�HXLTf�q,�)y�je�+��& M�ZD��`�Y4.�4�D�*M��*D@ ����m���l�TE�)5�����Ƌ�B�6�"m�4iQ*)j̚Er&C�9ɑP^i�R�����"�q��ͬ"�*L�D*2J����Df6�6�J$PɬH�
�5�.H��]EAQ*���2�2h��$Ѥ(]�L��v�B��TL�m���TDR���R
�!H��f̀�"*&jT���*���"�!`��]!S&T �QX�D��~����sAM{�/u��&���^��,	��e*GC������jf��z
\qA��U5�F��y�*����Ӟ�Μ�˙�{�/�S=���}tYT��f�oO�\�V�}�B;p�� ϑW �<n��蘜��f���3P��qP�φ�2�*�3�;uu��~k�8�N��7pr:�գ�
�i�����1N�l�P@N��Kd����pS��k�=ڴ=��lk�3\��fN�!�:��%�۸�7�D�#%� %P'I��v��eq{�Tb��w�`���X���Yy��=rz� ��2_�fp"o��h��K��d$l�Vˣ��\v��U�z"�f]�=}�TM���q�����tm�\��0�#^�ғ5҉�	L���ᐸ�y��/��w֞�L�ʺǢ�*zvϾ�+MƧ�ͫ�7�<ɓ6�~F�W�_�MF�#��\`#&��{���uh���x5�>��xp]c�b��KM�\/BN�z>�✛��T�ר���ثQʙb]�t=�m�L�����]KÂ�V��ͤ��w�ǣ�>�br5�h}}!AO���E�;�{w�~����3�fc�	�0�+���T��s�ր�o랗���8	�7�O�̝2ʙgo}b�t@w������*����%��u	���_���/~�T���`L���.v��u�6�1w���3,�;ɩ�6>P��s/�����XR���d:T��>˄p���̼��|vs��a���T� ������%Z���2ӮE{�X�>�{\//�#��J'2���/��^��EL�Og����m1�b������
�� �r�j����Tb�IN}��gO��ܲxe����G9#�����ǎO^Ny�q^�^.)��\}2�+��pԦ^Өl�����½��8.ԒuϠO���e�Z��=soF�2����WL]k�T�sA`r�q(���!9l��)����>�/vz�
'����w���3��f��RA`�,ŉ=<��z�2�НN���Hg��G]gx�F��K����}�q���+��f�8�O��{�r{�|���ފӼ3=^�p߱}Xv�^�JK��˼:�����9�|uR�W�Q�@}_�`�ZH�̯pU�էVS�9"&|�U���W��$��AS㸝p�m�n�	D�>� �2EĥZP��{��M�4�z^�|è�o��N�>s>��g'��n�s�f�S$�7�ƥ"k��N�>����Wq��6�{̇-�
�������ټ|j2����_�gȔ�&���͏h�a�D~#r��+��-�U����P�.l&%X��Yk�=��Ŝ4�%�5_:�mJ����ׅ�;���Jun�ޚi�WNB��f������ea��S����q�<��i]\����+�ՠu��P�o�W;iP�h��_�����6��y�^vz\���
���hO����Zn#S�Ά�'FJe@�6�-�zJ�9hm�o;2��Ǻ.�\8S�2JN����C*=����_�^�뇺]ᇀs�܁u�q��Uu����p}�c&R:�O�,\kʐke���pNa��9�WJ��z���V��E�P�W�7�u����~�R����3=��~J~�w2/c%%�
��/|�lO���df	�O�{B�5��:M���n_[�US�Z��L��!�jY��,
XA<� �\����rmꍏS��B�*�7S/���p*;�~�L�(�DR��y�q��7�ޙ��oz��ϯʧ&�G�T�M_"�L��	��UR�>�d��0�`�s���鳾��\f�9����8W�8�0�}�n��̱�J��|gT�W}�Յ�.�"�Hf_�����f���{��W��>U:;Y�����u�U�ŕ��SK�Ǳ��}�o��u[\b�C͋:�۱�Tz�hpЖ�{ �۴�}>�O}�z��(�B�٤��=��e��'W51�<�U���.�����@�՞C��{�:Z��l�^�.�fw{�f�No��6135�1e֬Wk�˃=�Z��}L�1wm\8%� �ӳ�wy;�:z3�X膣rh�8���҄%����l�ǐJKuv�Y��2ս[�}y�������y��椵:�HXy�T��T��D��� >����ɡ��=�h��C9
ٯk�\;����gO�'����L����>;��܌���3_)�Q�[��k`h�S8�q��G�c�9TD�ep7��L���S�n1upҝ$a9��G��7����xW�U8���=:̙L�U1�ch�9t���\����)a�c둗�>��9}e��SG�މ���ax]��u��F@zs���#��Uߨ�5t���3�kݪ{z�z�H`=/=�������wS<ePs�d�e����I����N�2���PV�x�d�;~W�/���yӽ:}KQ�q�\kY|=��7��7�KC�C"5�H5�K'��|������>��s�'�P�yiGtU�R��9�/M�n_�;ܝ�bt�q�u.9�_�W�}l�x�w�z=F�_��[[�ӧ�w���
t;��1�]KI���L�nZ�jL�1�ӊ�Vk����^i�w�����:�[��}&Qq�:rp�D�
��p]OS'=Ԁ�j�3��.�k=T����%���hOM��m�dU(i�P�W�Ƒm�8��to��^v�a�{�z�p���P;����k�M��f���['T��M��I�^��R�C(���6�޸އ����u�r�E��Jq�\0�݀�YG��z�jx:$횒_M	~V�꟦�5>˶�ʮ?�̅W�������xQ����:;�d]�ʝ�)E�T)��WF}���#��u�4���ީ�vY=�³�3�
��U��P	h9�b�Њ��DS��W����W��\9Q�y��r�����h��(����5z�eu��U��������y/JrF��/it���eg��7��j��}>�p���J�Ǚ&˿Mإ���ڱo amGI)K}tQ�j�U�jV��!��c���ꅝ|�魮ȘC�t�|��6�* ��<�:y��)<�|�v�_�����k�8�N렧[�ޡ�cw���)�[.�g�6(�.:�d��E���2������I5q���T�f��JFzi���i6��N���:��d�Q�@J��11<�h�l�/p*�CRR��e꒺���*�NE�����.������󸚅2�z	��?J�tz�Vk��S7��Ơ=OQ��Q���1�	u�6ۮ�� �P�����Q:)�"Ȧ�B;���띪 �Xs5��;�������~v����3夻4�2��g.�tއ;yN<T}h��>9t�{ǩtuޫ�`�}̙����o;h��Ò�ȝ��ܡ�z*׮�pM���̶���Pݫ:3��Ao ˔�NW����V~���OD�ޗ��Sۇ�m]ѿ���2[r>F�Ti~�9o�+�V�T/%ݴ�s��5n(����Xp��ʞÂ�+���ZoU��z!'w�=�S��T�U�Z�z���{�=��V����"���za���+�����r�'}�m �*�1������Z�NdߥE9{�n�Q�L{g�!��k�.͚�[�<g�]�j�^5����U�糭 &�9����� �ܮ~j3U�xU+�3��2���i�k��>�m�r�9����s�O����CĿm�c<oc�ҧI�� WcVE�O%'�R�Ų���m������d�ˉ���+P�x�]��D�g��:uH�l���f\��'Z��ܷp�^���y|+�l�N5cݕO�J�/��E矆�ȷ/�%~K:	h���*���)�Յ�.�6�+���{�j��^�/k�9B�����y̖�x�����'�qBOO3]rQQIU���S�4y�t�'��K�я�6zM��otT�!�ͽ���VD ��Ϛ��vBh��7��m�U0_C��%����ʷAW���8��\i敥s"�ѓ0�#��7,��)�hι\�֑}�A%��s(r���DGP\�.IK[c�_��y��������Y/�eӥ�R�5��3+:�a��:�ԍ�37�?����-�_m��x���/��\�}v�2�3�M�7?w�󷣶�����SG�!�=y���*�b�\D��P&
U���ee%�N�F��G������t�����q7)��3r��Bu�I�x�F[�Bk�2T�q %!�&�ݲo\��nbJy��(���|^��Fq��ƣ/����ϴ�r�`7��.�����+����$r�f��f���D�+k�\WS�s�ҙ��c�ϭ�l�%�\�%��k�_�����"=�oF�ٝf�EMA��Wk����Ȋ��~ޥ��:���0�:2wE�ޟZ�����:�������3Q���$��'c���%��J���OM�7i��w�nyo��U�Vn^����JC�7C�n�����2l�z<an	�1�N��]+K�%,�h���w����>���*��ầ�؝g����O*�]̋�J'+�|9���P�A~�u��z��_f�)��y�,Ԭ'��3q�}l{�UOI�5Q��Ѫ����yb�����l������1˦��j�������xe4��<o���W�g�D��R��|ڸ�j�����ɯqC�ʇ}������tz�wJJcT�F�
�P3o�n���6jfǗ�q8!��uS�=VY�8�Nl~��\źi�J\��a�m�WVѫ�[0�S���x����^-�R�E�^q��-I���g�A&Y�Q�Mљ���6)>+{��f�7�IA�����_%��KGJk���ט���/ׅ[��t�`�)�go�rD{�̬�qϑʟx��p�8�{}S����\
�t�u2��V��iuaz0�`���"�yõ�=r}B�p�$y��{�f��}�mq�T>]QU�ŕ��U4��{
���C���돲��K�ODs�S�Al�c��v���}::�'�}�z�L%�g3.'ܭ������>�U�V��%�xZ%����Zm�T�S(-�ꎐ�R�b�`u���FſY��8�����~�[V3���}��)�3�r���;���Fr0���}�/o��x{:p�R
.���D�A�@�L���S�n1up�D�i�m�q������:�T�͏�ޮ�$e�>�u�TZH�C�H�.���\���*��ۑ���Bc���ޞ6�fh����d�l����3Q��Q5eI�1������zWlߣz�w"��������O�v�YNG�5wB㚦K���Z|��A�܀d-7�~���mfJ=�<�7�3�֬E������S5��n���}�j�׻��a��Ct�
�wu�+ù�.$���v�i��2����z!v	�����$Z��چ�z��V2�Ydl%�X'w��I�}��1�s�&�|hT��:'=��������z'zK�n��\-:���mUѸ�'@)�큥��� s��y�c�|\K��w��l�x�j���^�yؐ�Z��S���5����|}� �����s�X���L��C{u.��n�z���ם��>��d����Ld��'��or��Re��q\���w�ʭ�݇8sA�̰�l(�߫��6|�99s(:8�O�࿪z��ΤD^5�cʩ?0jc\��d����d"�m^Jh{��1q�T�(�˃0�B_'�p�R�	@�m��+���)Fꫫk����e�g;�U�4����g\Ν��'���/�;P��W�.��}hg�LR��]�Ë�0+�#T#oŻ"�Y<��E�a�}�ntgo�F]�$�#�K}<�����Q��\�/�w����>F�@,�UP�9~+	G���}>���7:;~���ۏW�ɫ�Q��|��X&m�$ˉ�G�G]L�+�J;�U�ԩ��rZq��sθ[��}P�xsDn����Ѯp�l* 	�`L|:y��);�2��
�n�`�X�q�l��vb�l�(ʎ]^��O*�xa��-�i���J����Jo!4�b���Ň@	'�^��t�����2��Y�n��2�_uk ໏8��W����:XHr�T4�>e�]&��i�1��m��������7��e�ݴq�z6q�۽��,���Ƨ��8����2�-�rQ�����F@,��E��js>
pr�\0{׌���I����s{q�ɳ�M�)���u�M��q:mӨ��d��@K�0y���ղ�����Ģ�^�>��äU��b�H�p�V�.x����[n����M)�3����G�G8Q�o�Ƣs�vb�Cj�^�t�i��j�L��Ѩĺ�m��0�#^�ғ5҉�)�ieݵ�l�W������O�:�s;g�Ҵާ��UG��y�&�t�#T�ى����f*�i#��U���6�l�r�늞Â�m�~ͥ��U��$��bqNI�..箺�k�=�j�dO��E�ύƔOP���������q\�I��A�ܻ�`�A��әma�ɧ��7txͨ&�r��������kީ������s�8�x֭�����k�iyF�?8�?���~r k�<��2��<��V3O��p���R=}(��3Ƌ��W�3k��ݢ�w@��>E�L�'}�`
��jȸ���ʘ��ԕh�5����v���P���DD;|�G�`-ʛ�ūhܳp����(Į[կPx`��b\j�Y��U���%0�EH�r��R��<2���w�G����V_�$Q��:����d��`@g1\�*�������2Sj�)<ܡ�v_h�o��_/��ݱ{/�Z5.�k]{W|�l-u����[��&��J]sw��#���LO�5Z�t��F�C$�rV�W�e����[w[��t��S3�\~��B��X����T\��yo����\����̽V�w���;���e`㹃%iH����Mf�
�R!͉�mP���Җ�͛{�j�UƼV�Q�*���z��j����ו��sKf����w��L3I���]�[��ˋU�"�l���{�YB��ᲂ}w{r�r���7rd֪�q�a�y�N�6r�D��ͱ��z��%v��jk9�F.F�/��D�,󍫲�y߹�P���K�l;�7��Pa���P賺���m�ֺM|� ;�yp�K/2P)�m�&��rc�Q6J�\�����$ɷ�����s7|(A�����Ŋ�NiATDYłA77��~�Y��S��KU��l��t��d����%��<����`[��DkmI�������ȴs����#f�;;Wl[�f�����+�S���3KS�m�u컛�u[K+$�� �c�t�vV�;y\;ub�T�e�WC�d|����0v�U���zMot�OeLp뷨�m� ��!+2�$4`�>ݰ�ּj�VՆ2���YeM��kQyv\��y
	�5r�։V�+��&F�����iü���Y�4��u�ә	>�x��fNA��:�8t�ڕ�X��r,.{�����S�,�9�͢�=]v��Hnج����TͦhRJ�y�؝$�k��݉�v~���ہ<�N���k�r���R���y��ŰCnqlY��H��G�,WЯ�+aݦ�b��Wm>lV�����Z�ui�V����I0�@������f��%q�)ǝ)��u��Ӝ��WݣU��m�maiq8�	ק�46m���V�-r`y,΢�␍�ED9�;y,�3F�0
Z���w|�\�V�to�l��T��e���Ϲ6O��O&8�;���"d�E��ٚ�#�-�j��`W1^�u�EA�-6i��gS���ɧ��8-i��L,ʛ�|pu���e��1�c�1��w�)O�<,��z�`&�^�h����&f"W7j�_2��9��զ!�S	6IZ��4:o+}�2��{���ԣ�S0��$�� V��6�Tc&#zfx"~O �M�qN7� OY�L�(0�b���o�f�ŝ��;�ꏴ^MI�0�Sg����}�vp�n�2�N6fo���8�t��ԳIg5��V�DL�s_Y*��y�
���p���+��/��2��^l%*O��>>�̙��]�m��18�vﲵ�H�-�rY��_�����&��T@�M�Y� � *�M�L�AQ�|hE
Nm	���mf�b)rd!i�"H�h ,&؈�"��	UP�,�0�*dʑ�em&ERB�R&�X��2�b�ˉ�mf�4&T�`R"e����P$�]6D$Pb�	f#s�����h��#I� �m��d�B2b�i	
"�Dbf�4a�\��BR�B!��M�
�@��*!���T���M��1T�jD�TDS.��
A ��(�Ĝ�	""sI��m�E�h\�i�	3M�Eb��Ƣ"�¶6��ЅI2'9��TP &L�&H�J��	6�*.c.nQXU* �"�$�aR$.I�J��.�H�Lm��`�D�@PUd�.d�@���L�m*""�")*����4�j�r*$J�$!�o�}���]�l�acm0��5C����A{ܑ�q����q�4|��w����F˼+̊_Ḟ��=�A�}9%�cy���������AS�)Uq��p>ٗ\FL��e�w���������VMn��`I�\��;�>�2l;RIu3�T	��e��֪M�'V�,��V�g\ƭ"���1�����y��q�G|e��$�2��_.*z��E���t�X����h��9"=p��이FХ����㩪��g�±rx�I�2��{�wN�WP]��A�Ǵ�,}��>�l�S�AĮw��s�h�>���θ7
�B���F�����?�I7Q���z�Nǲ)�G��7��=��}q7-��yϩ��N�i/��êBiL�5�S�<ݪ~��۽ѷ��7��~d9�X����>
�8�ظ�e���E�z[*!��6�@�>f^��::��*ϖ���qE[�R"M�pzH)O
���wå3q��F_���n_Ͼ.q���lW��E�}~���e۰8֒<vk�3\�
�%N�B|����Rө̇����k�@�$��dˌk����'��vCC�ة+���_�(N��b�G�ڭ~��&��%ߗ�s�;z�~5ylT|�3����;��T��l>U�a9�>��:�Ia��>[��g����A_���Hx��dk6�`�!�aj�~�$�sv'̻�Z�r/\�V�o~
�ZН♢�WC��R�ޕp1�>7�6�6��k��GʧFW��횓���<v�Wr<܅3�	�w��P�ו �l�z�zam���S��t;tH>�,=9�K�7�[7*鍏��>>�k��w��7	�X��ީ��D�@>�E.c����ٜz���q��8�/	�ϣ:S;���B���/�{j{�T���s�,
?؀�ve&�WMUb�QO��ENq^���<o�*G���)�J�:�zW��]�z��sʽcc��U��7�-)8r��c�&tt�'EJ��p�tFl�I�m�1]0؎�b�����=#m�m�>�ͺ��4�m�3�|O�W��i��/�n"�PEhsAs�<�c�>�lkڜ�`����y�p}�7�+��<h"N���A��.�{�FF1��=��[T���W~�_�v�b7���x=�=��Dc��7h=>�N��rx�qD��3
Njf��w��9��8����'�9�����]=���Z���Ijw���Z^t����A@�z}��d��3���`�q%07+����2���gE'�q-�q��g�����އ��g�����@�G�A(h~�2�q��)�[wr��}r��<$s�uػc��¸�.5��G)57�.�r���ץv�!�[%��[�xk�.���fJ��qX�*b�R��������y���:7��g�����E��;.g#w�>7�s=���טvo�o��?��>* E�$l�Z������Ό_Jv��9��G����}j|���[�%��'m�#"��F�����'�M�U��"��ڑ���R�0����ޏ\��A
u�g��"W�?WA�^�t��v��@��?���f;��73w8n�"�������KOD�=��#Co��\CJ�/��ZwRDt�vHw03�\M�3�t���͙q�u�p��-��-:���mU��r���`ihzhf���:Y<��M��};W��V�׭��.
�t�0�VK�����;�u���N@rW����y�c,z;�zo��9��6�3:��(����X����Sq]KI���L�F嫇�U4�Ǣq\�߫2}�Ub��Ï�۟z���p��_�5��x�f~��aߞ�����~'=�H
�k�����Fuiw7�����Q�����gN[�_��x�sCٰ���d�a���s!U�a~��)�xc^`~�Q�ۑWw��Ḳ�߸���U�@?�u�2=��.S9�J�f�|���ӶY-�'�]BV����27a3�[��{(枻r��J5��; 9+7I� v�A0� )��ќ�K��]�b�LW�h��HC�Άh7�op�3�5~��&�X��
�Ysz�Wܥ�bX��M
�8f�x��,Jۇ��|������Ob���P�7�u�h�Y:�������e�b�?�/�d�ƨ���FjrVS�8�w����>��o�F_�(��f��f�;޹��\ʎ�3�n�\��Wp���O�{%���p�O��c}>������V�N]��3�{�ϙ&_�P$��e?@]P�*e)c�}tQ�V��^�oO��ei�c�����^[O+��;g����;\�`�,���e1���f�)=���;u®%�������OG���>Ix����.������T�+%� wW�@1��E��js )�׏|~<}������v�/�O�����m���v���N�N�i(�*���;E�N�4�VM`| =/Q��1��ox���<����M��@�~wJe���!#9����]m�Q��뢽�C�n�F�e#��޸l�kF�.�tnu��@t��׀�WJL��V )\��qNO�*˅����D�pf[6z|*V�
���4v��Xz5=�~��wF���2n!�@k��z�^�oו[_�JΩ�����g}2k�1�dx���+��8.+���ZoU��y'w�: /�X�?�a���M4d��~�;wN A��O|�����,Ռ�"#��衜n8�fu	�dù,P\k���u�p�AE�<Gl4��7����#%^�-Q["��T)0峲�>]�%�c4dȬç.�*��B�\�����+U����3q�n�A��Ip��������,����2�)/�Er�'}��䝬[�1Y?���e)��ڹ��i{�5O?�Ճ���X���S�xQ9�f9�	�0����z���B���ip��|� 3�S
�ޣ9�s+�άf�o:���h�g�l��!ể�m~���韉~�h
���8��*�7�L�'�J obVGI��*�[>�%Z;����rw5�KSb%K�;�;5��h�����C�3�+e�h�6e�X�Z<��nᲽO�3@ޗќ;�'wK��C�#���p�}%�D��2ï�΅u2�b�+U�����p�+w<[�hU�l�=X��\}+*;���3��ܐt���u=\Ϣ��Q���Į�D�Un�p�h��A���G[U: ϙ�p.O��$�@L�H�9=�3;�}'���w�m�l���84���P��n�y���c�8{�x�J�E������F�UK�ݗKێ���^�Ĳ�t�`U��뉿���|����'\4���n�	�2T�^q�ߩz�����3/�b!h�݂����wu�����V�yJ�p{"���{*;����ׅEOט��M�>���@ʝ�n�%�`F���p3t�-M�Ƴ���zXI{�����$�Hˌ�rA݅�ԝ�ϓ'�/����2��up���J\$L�W_3���Q���|�}����k���a��^ж=�4F��cg��Y�-L��nN�Dķ\*�qѸ:S8��{b9��6ܾ%�}�O��;</U�U>����Y�w��f�^S����R��(k��yo�ħ~}���a�:��tG��*�O=��ng��1�-9p5����e��5���r���v^	�/�w��s!���:�x��x-�k������ȿ��3i�v���/^T�_l�z�zam��1��w�|K�w
�^o�r�?w��������7/��9�����{�6�U����G��|���/@Ayȟ/{m����\���S�pjV��gJf�/��*�zO�j�WO�U����a�o͠L�n�������^����P8r�e��S�]z��̞7�P+�����'"��=! <]�c�r���|;(���Z��^���'\��tt�'�"�P}8J�0�`�ᕽcIq�|Kk������I�>������N��}fP�@3���|n�PE]��>�/<EQ���`7��%�~%]O[h���h���ަ3<�xn��e�>s4�>+�H/���^՛6��;C�mh+,�����G���%7�}����W�z�6c���Դ�Z�!ܱAo$m�=%&�I��M8��
���E�';�{Ӯ��f�u{���OB�ҁে�t��S���1���7��I���&h�R���G�[W����t{�x��u_�o�#��x=�Kg1�:��gGl�ǂ$�v=��1�����tO�Ÿ�
ڎ���H���w�v���j�d58�H�/�R2�U ���pcB�3��k{���2܀��J�66R+�-���I��ܷ}��B��=�!�8{=C���G��3��nv����52��8�D�"e*�cJet9��up�Jv��W���S����I���"�g��"���)�����3"��F��a+�m2y�ОS��|��T�e+�P��w;[��BUz��z��a��Y_9�D�D3Q�*���2�퉘�	������=�[6����=W6��Z�s}wB�L��X��x
�?\�](��d-#ּ���\���KQ�z\S�����3n�O��Cj���:M�l/��X��i��PM����gi��^^%8��g'�g�<r+%�|w�·/������r�����~ל͠p�x֜�&)P��[��p�F8��7�]XM�t���X<�k���b��� %�+V�H
�ﱆi�Bvw�.�ӿ۱E[�^�C�g.�,˶xF/.X�R��B9����0��.�G3���ƃT{��k��v��;(L�
=�7r���:�_�˙�Х�Ə��8�^�2�+�i:}��n#r���*�zb���");�9��F�B�6�����^i�|���qg'	c��
�*}G��~'3� eɼ1�Tz���+��o�`qU����k=�n�f�^��z��D�
�%�B�+�Xg_ݻkЇ��y���`W8F�
�v���i���3��U�4��ó�S��'�VLo�L�c���H�����S<_ս@5�dGXJ�Q'���t�^�w���O�EGo�F:�N�U�S��k��j��&I��u
⌾7��o�������ef:��TST��aJ���H�=vm8��ar9�6O���'I�,.�W2��辺(ڵV*�ԭ��k�����P�lL�M{�cQSXƟ6��o��`�<j:��(	�<���e"���2��
R�x��q����tz��x�q��p����9�ah�(� ;�� 0�����S�<�J����g���w`8�T)��[=)�C�}�Ʒ;��:���:��d�Q�@J���]��M5t�<���ر�Kh��Нox��>��]j���]B\���<��t)－o���}]�����'ΐ�u�,�OV�k)���:��xXf�$�Y��2�%��aJ�X�%h0����^����<޲���*�G&N�̌��&�k}�����}ߺ��r��������5hyˮ%�������k�2�x�Y+"�=R�m9��fk��V�\B$?�mu�ǫ#6�2�3Ki�m��_�:`~F�Gz�B��e�z6���ft:�-J%
�3���
�^�
��W3�}Ҵ�}�����o�y�'�8�E6I�}�{8w�o�}X��L�̟l�;5��a�*{	Ŵ��m-7������IӺ�缳zj�qw�!7�ߜ�o��,��_����Y=C��e`W�KÂ��U�����g���T�~�Yoԕ�����w~z�ޏF'C���V[��b׽S�{ �s��0���z�����KB4}�Ⱥ��=�l�J��UN�nu�_G:��}�k��+rѮ� �hn�>���$�=�vpZO����u�7�L�'�K w�Q'{���Q�gВ�膶�?��H���]ȏ��vqF_��DuIhGk��zV&=���R�^:qn�$M{۳�`/3q�qʟx���V��r|+I'L�U�Ю*e���T�9���.�.ja�n(;{/�}>Y1rJ�Îm��Pi�,�j�S��mexj�k���4툳wl�M剀�`ef��UշYN�8)�Եwh�)$�`w �ܚ{��cP��I]���LYvo�m	���`�F� �/�kŲ��n��o�����߿g�;�M\=���fx�֤��P$��5�%Y���Q�{��ý^ا^��\DrVƏD.��c���j��ϙ�b��,��e?�Hϓ^�l�C��q�V�\s���[���������c�8y���J�\@�(�VOk�7}�s5�{��Wf�l�U���H�ς��7����K}�ܾ8���\<u#.R��b(�{��Z�Tn_I����pW
�%K�d�#�-V�p6W��=Ǳq�ˎN�>s>���;Xo�_G�b����] ���@q�3��2J�f��7d���\Eu.:7>)��ƣ.9��3�ޛ��;�ng1'<�Ģ˜�_��_)�H�����ck����ȯ*�7��Z}� <2�Fݱ�w�ݸe�ӑϚ���;2S.4&=
6_��\Q;0�����x4���d����蔠d��6�1����N�E�y:
e��9��((�yRl�z�zah��aR�	�z����B>>x�k��Y��i}��lh�����e�X�#Z��6�U��z�{>�0g��)���?;��T`m��
�ݮT�$7����*1׃OQ��Ɵ+�Z��%�S��9%��4.VM�p� �	�!մ�����*o$�df�墶.;6��;R]�w�E��r�p���hXAP�lr�t��a�����]t�^��!�Z
 P�oӺ"�j�V�N`�-鵸���:�Dg�4v�2]p�Dⷩ]@�uv�<�9�rMV�v"+��\f�E��,��,APf^/�6��a�ҋ��5ն�Uͪ�31����9iX�֖�.OQ0<�w0^��S�	!�z�"V,�no 5�]N��;G-W=XQ��m^�m*�GA����4;G>6%JU�XC���	˾@�)Czt(�����DX�2Vs~/�c���b�s�0�g����77���N�X2ל�{\�́��5v�:Ņ���sZ#�8�>�Wέ��\��t����S�zq�;wU�{�u%m�Coe�8Ar�`����*�/�+WaV��Z��$G��k�%[~�G#�hS�s�ᇑ�y,55p@.wU������ioU�����ӳ�{ޕ$p,^���a��|*[ԯ+y�=�z;�I[�wD7k��H�2��b���-�>]|s N���}Alڔ�lt�>��W-\�'�/%��i˲��`}��v$Ja�tݹ�.��3M�pi��@<;:vk�A���=ˤ���0<c˕7�{�6j�݇N�c��,A�]�JC��Q�s�(�%��Y�1��8%^qfj�,wa0|YB&΅}`�K�.WQ�͖Վ`��qovV�aw�H�D�m5t��}j\��o;zB�5{cvl��s�&���>���i��ľ�7������b�������\�kn8P��'{1:�P�r��|���a�&�hۇ�5���%J&b�xd#1��pteuY�:��Z��P4�㺰�q�!j3i�gv>���M\�Ԟ�^m�W;�o�: ��ih�O֍���{*K�ںk��0>�A�/	�d�m�wA]����,��jh���]�xv�;��rJ��}����|�8Ž8�٧m��g�k }y�&}���7-m�2̢��NG�����'����P��V�̀f��8t�����X$>0چ����d��I�.��r �HpXx;��s9z��C��G_S�<�����t���ga2 �r�7�LWK9oMè���O��:�9�p����D�͡��Ջ,�̢qu`T�;L[�Y��!k�tђX��N|��ƪT�iլ��+c=KP笍fh��"�K7\j�{�+a�;�Y�n=6��3�g���n$�Y���ڠ����c��Yz���fF��1Ӯ�3�Z��Dl����g˟>FR��q�:������)hB���D}�܉�& 	�]q�/um%�W����(i��[��W��w8�u��|oI�=��|�[1����Y�n�9�m����~z@$
K�~!6��6�B"ă4�6�m���JLʈ6�5�����	b),(D��3.�m�k4@f�p2V.���2�D�6Ѝ�"�@�bQK��D���!@�L��D�l�2k��)M��#&���D�	h�"D!B�ٮ��v�,m�"rh)Ds$�`��L�m������h
��")fm�B�Q*DVh� �"ň�!m��TL���HT�M6�6��$\�4H�Bd*���&�EL�M1P��AR��� �!�D��dRBS&�U(��e�"!��("E@�2� B&j�!Y���3f*,*!�"�a[]bͰ��ԛLMQa���&��$	�"�j��jH��(��E�D�Q�֦�m&RB(�&4�P�l�I
DDL� " P!!j(�I�)Z�3.�K��ǡ�����D�)�eޏ�Rr�.fJЗy����g����6iD<ɍM#��]vɼ���]�q�t�9�;5�=�Ua[�����S�$�'�>Δ��_[�US�|�F��Dj���E8������>����q�U����V��\����+KNSK���&T
�sWЪi2�E��w�e��{��`��m��iuFn��.#�g�/�C����R�ຕA��(b
7�>�5°_���F�Tݿ��"��S�����{>��;.�{�%��T8
�}uO������~��tmf����Ë�1G�Ȫ�ތ.�!�r���n�=���ޘϻ}S��N�	�W\�ȣJq�G]Vwe��y!$�ژ)���G0�xs�-��c����O�ӣ����K|��E�tפ�<$�1���8��L�UPY������CS�$���uH˥�S��X��;'�K���l������,		S��EzՌ�)�D��}��g����'v{�w�F�Z:q�n�eÚfk�2
5q�DL�ZiL��
s�.����p�Uu�ˊ>���a���p����s;��6�'\�22�F��J6H��}4.+�s:w^;������]������EB�C�nT�/p�ֹWA۷�2<!����n;�5���v����Ttc/+��m�%|�_=R۳NV6T�l�)Y]l�
��{Y3�S�dݑ7��ɨ�������Ȉ�tyܨZ
��._k\���>�wOV�p����+�E8ԮF[}l ��,�3���j2B�Q5eI�1�ك��<��Xn�f�.�=Cj�^�qJV�߾�H;֮C�UiS%�,|�ǀ��rDt�uW���s �52\˾�>���#�\ꃛ9�><�_f�-7�[mU��r���4r�x۴@��m����&nʐ\t�=@�n�9*������y�?pN�@j2�r�����N�rC����k�A���չ�^��Ʈ���	�_�^��J�
���\Eu-'N�L��W��G��1E;"g��:Ux�%�y�k����^i���3�|Y���e�������N������9�Q�JOF��^7� 7ݾ�=�O��{?U���qW�3�in0xx��+�o(�O�ǯ�ׄ����NX���d�@�a�c�̎�i���3��U�4���q��7��Ov�/RFsDľ�Ž#=wn7K�˨�S<g\��i��)Y'���t�R��O�G/Gm%�]Oo=��۞=я�L�K�tx����ў�we�e@(�UP�K���d����������, ��!C��R�(Z�q7��tfݎ��ڼv�=T�SÃ��W�Ê�#A�`�f�Hy���N^a�wǦȑ]E�3LJf���r��q��u�N��`�F�ͭ�b7l��k��芈d��$A��o�lOn�Ed�-��d˓w�V�t�ȷ�����l�],v��@H}P��R�+�J;
�X�J���-��Ds��Gun9�DN�gt�����ꅀ�<���� |
`t�3ce"���u��U�պ��A�W�9��t�Q�<���㏤��7pr�R0��G���[$I�i���ϖU�f���͉�q�v�r��]���mZ�>�c[��z;����N|��j8�	{��;u=��N���[�a�үQ����� *�Kz����ա�.����D�n�n�a]�˽^{^ѻ�S�Q-��(_�D*]��2�/q�{�	��h�e�]n���~��5�Fbl8����dr�.݀�]t��S��2���O�D��>�g,���:�T>���o�\����~*e�5�P���<L��P��P�/�&�f٣��ς���8'�ћKH�%����V�U�Os|6Qڗ㚻��✛�9P�^��_��ޖOW���'ةxpp �(�tN�}�ޱ�QM@����S�.��s�ޏF'C����V\=�-{�>7� ݊�߿e�_�[�$�� b0Z]����%��ڠ�cL��3*���_Zv�]�G��?�b.&�hY�N_�X~���=\=7�w�̥8��S��C�'k	�X���lؔ�]�IN�
�qZX:���7�90Ф��y������ޔq��U����
Y�Zd��>y���y�cЪ��2��<��ہO�z�2�-v�_�J�����]��]=S^|JL�w�A�w�2Jd��I{%����K�:��%�x���ne�*��o��]��'�\��3�t��l�F̸�KG�Y57�V`�v��c�l��[n8���Y|�pI�u�\?Q:=m/ܪ}O|���悭O�����>Żѻ���Gm�/��Q�>��ަ�� ϴ�G�7�Z�������S���@�3M�U��X�Q�s��u�V&�s�4{����tۆ����0�\�<'���r�}#��^>~���y����%�%u۷�."Zw���SG�!�=C��8mR�QD��g:�Ѭ���G� v83
���l��+0*��b}q7�{����Ȅ놓oH�۽��w�9yo��^	)�鯑 r�����R�������8��{c����s>�٘�ˁ�3J�M,�O�;�xz��.w�[�#4�I\nJF����\*zW�:S7��g���_�칚
���y��H|?gJЖ��o�I�҆b,vS�`J�R��%�i�rn��(�,��7�`�h�{Z~S=��d��)Sh���؎a�����n.'�T�΋Sׂ�:�<p-y�����b28T,>ח;�ޜuꫯ�uNq�a��2]����+Ŧ��uD��%4k�R�D�����p6�*T�4.+ʻM��q}X\ķUS��D�=��*���]ы���&��_����W�T���9Bw�~�.Om�<C+mo��K���ǁ�u�o۴��ڮ� ����y:
f�`�~�b�^T�[,����I��yXef������k�+;�U�o��z_oS����2��r��O*���������#X�xT�����ٳ�P�����jV�8�V����UOI��Tj��5��h3�ևumϽj��瘸^�I��p�VC>b�U�I�O�w��j��9�S����6^���L����_�Nw�zWގw�n0ߦp_98r�P���R�ษTO���(��β�F����m�^t@��I��)�g}��5O����TῬ�_\A�=_:PFr7R�{���O&����y��-��{K��]0E����Ct��s��7�;��T�(��6��멺y�^�n7K�3���g������X��-�C�-� ,n�,.}:9Vf%k��x�癑;3F&��dg�eY��U`-���ɽ�~����|�H��2۹��W��F�Ǖ�*�^>�,�����d�a��t�&_Pʋ��+����r���]��'���f��[�N��7��f��*�d�l8з|��&s+wS��oR��G��$���?�u�I�j�7��U�V��!����ZF�y�B�l*Ki��l����
���%�Ht���	S�l�W�Ռ����o�n��z=����W��z��-q���Y�-98z��q�FiL��}�G.H���A�)�Z�mr���ê~=���[���+��s�C��&�w�ꙑ_)��uL%ch�9��'cќ��
�s�-�)��.ӍY�G�q��g>�em[��Jbc�1Z���*N�1�y���hK�ufk�Z�^yfKu�o����~��a޵ro��kJ�/��_���	�H+*R��� �l=`ꊷD�d4nz��%mfEd�v��N��c��WF��t��큥�v21s>S Ｊr7â�R�H5
Y=@�=#��ؐ�k�A�����Te�]���Z��"F�V]d�:8�]02JU0|���s7������8ש���ZN�F�O{9�i{���n��Ƿ���*�ZcЛ��VF��=o��g�Ϗ}>ɖ?��,�[8:��!c���~Wo#����ˇuݗD�	�ZĨ�K�K�N+�����A ˤ��F����.D�U��$Y��u��s/�����$i�&O;�+��OH87��0ܖ���˖VQ|��b���	 �83�yxP�T��z��y��=۳^��7���&�*@W׍z�*���ϩֳ������׼b����p�Ne���F�{}�VP�Ǽ�5ѯ(�t���N��J{�dz�lr�Έ�\3O�ok��w�t�P�f9P7�i�ף1�ꚷ��31�5g*Ҫ�:��MP�������N�[��\�^���3k�^�8W�8�r>�Hwr�:j$�j �T+�2��VʀQ��+�^�.�|�K+24�}g�<�_z�'3�P��ޗOi7:;b�z���N��`>�WS)K���(�B�V+a��tnF-����=j���!���CθZ���GA�A���fll�PJ�
�I�̺�C��?Yq�ԅ\�|0z�k��|w����uH¸%� wQ�2�ť;�K�����k;����Nd@S��:ტ%�h3{HgCu�K�Q8v:�@�f�g���x{p�k�5l@I�D���WQ�����Q�oY��=]q/���D�ͺ�;[�B�7�hm(��\K�L�ʀG#�d��{N��J㷽P�Q�������p/�%�'��r}3d�_�w��H5�gR��V�,�"WV��C�-�z�RN��ë�d��k����p蘩�U�&�� ��	\�ۺ@K��/������_�ڜ��G#m �%�O��}6^)�����w�����#np|��wpotys�6��3^�]t���N�3)��Ǣ%m`���9g8�+Sۇ��'�&غ�7�^r黓�]	βd�ɺ_�������#�P}<6����࿫�k�L���ފ4<Ю�l�Q�WQ��V�q�S��T��w�oK��,���]q+WRy�����ٙ�}�&n���)��wћH=ʫls�ތNF�宬�{x,Z��|o�(�ς��8���r{G.���+9��;=Xz#:���[�T�Q���e{�X�>�{\=��di�q��r�7J�z\��r�̸3Ƣ�q^��u2�=�P���Q�<��[�际��O�H�2����������|�l�	���	ᒒ��V�������=�.���d��+&:O:�)W'��Ǽ��$W������½��8)N��΂Z=_�T��>FS�=����u�z�U0meVBr��j���������RA���&|Pwչ�͖�'n����ȏ�-{���=���j�Hf9�|ڸ{�3�aX�<x2OHe}��qz��y�Y���M����c`���ث��E�LK��!�w��1=M����@����Ԇ7W$���
 �⃥�k5���װvRX��,oBو�/���{!~���%��J�z��}=x�k��t�V���<�����/��J_E�/7@]��h;	�j���nߴP-:�ֲ�=������p�S/�w�~Sތ����,�@@Zt ��,��+0*���D�K}�s�|w�N��z���㥤�Bnv�����K��=5� ����)V�W�
�8�.5|��e�LO��-�T^ks'<��"��`7	��-ϙ�I+�A�H��"e:�W]K���)���� /�,��ٹ��(����ѿ��Ĳ�%�6�6����3���Q*u���âa\Ӛх�p�5f�s���5:���1��vd�'.�|�FEl��I3�(Nӣ�w�e1mv߭��>yF��/�:��ݔ3�U�<���~N��l�o?`��� ���%k��S�f���^^%8�n�������[�ƍʺc����k��w��+�P����L���;*�߽R=p��� �r#2amz�5+	��Δ������UT��y����B�X�=~vFۏe�j�?�R�����z���?c�ջ߀���Z��K7k[�vҴ��+�`G�*�K�V�*�+�>o�"R���f�<�U�L����vEZ}dPN�<��¬͜�!��r���}@�=Wn�\՜ȯ�K�ͨR���j����++^,-��=�/��r',΀�k���8����}1��U�VIQ���k�#�S�G�ڸ��s��xo�8;�6o��Қ�����^.~�����E�1]-L�q�n#�&X>�t��R��Cw�����7Y=�e__����^ś�]u}��J�<����#;�]]XX�G<��峫�u����LWo�x��Cv��m�o<7����xI�b�����e�n���wz�w����Z>Q��[7h=7�I�H�"���'�!_х��.O�G$�a@�/��[4�z+��fݽ���?d~�m�\���^3)/�j_���ӿ�)d���U ��z�@�������0ll�W�Ռ����oY�U2b��k5�]u9E��3�q98z��̣8�AF���.�)N��)�2�h"�c.=5�>e;Tn���7��)�F9��E��'[w�Ꙑ�(��a+Dw^�;�k�B����ٳ�}V��)Nq���1��ˎ}l!�ϡ��%z������_�T=�x9��n�[U����ڸ~���Oo�x^T}^�v%�6?Q�J�;�n�S>2�=�>}������Y%�[��m�K-����l�[�-��e�Km�Ym�2�l�[�[m��o����,���m�K-����d����m�K-����d�����l�[|��d�ۥ��,����l�[��m��o���d�����l�[�[m��o���d����m�K-���l�[�1AY&SY�h! ԮY�`P��3'� bDY��JQUAP	R�P�E**��$QB�!T���*��UH���@)
�JH��@H*���P��֊H�" �
II
�ԅ�"��i�
BP��P��e�HD�"FƅP�UUI$�6jU�JC`a6��*$*��Q��i���0��)*��QR�"�THTREQREEUUCFQ
J(�4P�*��D�EIT"�H��J�ER�  �����i�EÎ����4�d5wj�UV�wM��6��m����U�[p��u!n#����;7uZ��멗f�Z a�΀�:�a�J�TUUDD�  W�(i������-[ֶ�����nu������V���E��� h �=�x
:�= ����(�Q@ 7���@tP  wx�@  �9�J)"�E
EAT	� 7����T.�k��zĚm�q����c�{�!Js�j��-v:�m���U���J��^�i*U�Q��+Z���9k]iָ�
�PI*EREB	� 7�^���.��k5�s�� }�4�{�"�N��
 ��z�Bt�v�u��:�N묷m�u�v��佞��w�[ 7RF��Z��$�	T��T�J�E'� ���wnԳI���kԶ{s�ݡ�K�v�v�gWcm���r+j�u�nݨ�S;�s�t�⣺kW[j�7m����[m���SN�sn�49�i�s\��$��UEUZ�U�  m]��ї%�c��浑����m�IWgM�۵�eGm��\�l��]�6�Sk�gp��;��M6�l굩n�����QVө�-�����3��v�E̛5HUR�4�  c�٭[�ݮ���R����5�q:ݖ�uE��ݧwnu�9v�UuZB8��ڷn���8��Z����w[�;�۩Qm�nE��wm�
��m]Y9W:�[N�JEP.؊T��EV���  ǽ�m��P[�̷Z�#���7mj7n�]���V�s��n�9uݪ�ۭ�{�Vm�ݻv�l���%�t��En]�,ڙ��r�˫��֡]��ۦ +��#
�m�Q!*��  .��zꝷ[d�N.��n�Nu\�ƫM݈֮�maL:�n���k���ړ��*�uۤsv�Vڻ��(ݭK�v43���t�i�᭷N��t�8ꢊ%T�TH�K����  �^zݝ�T��[��H�n�e`huZѵ�*�u�wcknI�I-�vhÝ�L��Q]�.�L-h��v��l�n9�m�2e�o��y^�f��vw| �=��2�J� h��$�%  !��1�J�Q�P  E?�SM�ɐ�S�Lb�� �M%OF�U5!2A��?_���#�b�B�~]��G�۽�P��Z<����{�&���E�[ko�IO_� A	&HB!!��IO�$ I?���$ I(H@$$?���{�������ߋ�+��Y�W���F�M��Q\G&��Z3-,���i����#2C��k$[��u��[��i�J��:���1z+\��.��J��!��c(`J�i��G4�,f��5��$��%���MGj�4ݍ�b��\xF� =�[޼f1�t�a�˛{/)"�Y�5hf��	5+�@�����g+.�����*��q"C��j&}7-��R ��vd!աՋ2V�D �*{N���G����.��oX�E��a\I�i)�j�R�t�zq"�U�*+Cn���U좶Q&���aVL����J�����%M�*MU�2���J�1K�����1�0e{�ck6�Tq��m�ւqգ�4��I�2�[�ݺTn�N�A��kF�,���o�[��)Ĩ	B}�P;�[�/u�z�S��j]̸�f�,�ʺ3+lP��U�sI�C�+6��E��tY+&�-,l�h��MN�Q��j0Z��h��&�;�j-ac����z���J�j�9A�����,�n�tNY�x��ǎ7���j隷��՚�z,%�.�͹z�JR�8��򺅌Kҙ���R�r'{y&X�w�(l�u��4�4�v��2AN��a[V!�j�F�w(��5�L+��m�=̫s3P-�Wxu�CZ��JW7b�P�O)�O6��z���H;�{��g4���SR�K4b+I����c����ZbI�Kr����̼����!�A�V���@��&.�ud�z�!ʂ�f�U��)�F��!�t�Y����`x�;��1��^
DMYQ�n�(�$5KB�ԡi�v`P��ioR7�c9�\�^i�[n�d+f2�<��xΛ�CD�>l�	Q��h�A�1�B	m�C0�h��{vˑE-�nbJ�ԣ2(���e�7AX��J��O�IɅn#-�i�"`j�U�ʘ�f�m$Jj
;��7h
+m�������d���[Y{ �t<���
	U��8�c��f�[P�u����	3v�V�;��l#\�%Z0��2d�N�R��@���ɛ�%+ȷ:�Z(l9���EЅ8���%�����#1S�u�W���HQ�q6ҥ��[�Q�D:�0m�[2^`�u)� e�TCH�j���h2�n[��TMR��8�;`�`�dZ��%f�o���Xn���)<�X)Z�TF���j&�P�3rf��j�$��W-�q���2�n��~S3�Zǡ�B'kA��LTն��a˦6�5Р�*ńtZ9����������!}p�jV^�D �O����ԭ"jE��k"X-F��ã������~'v�	+y��kڎ�T0.��4�̧ՂQ��92d1D��tά��ҍct�%m�S+E^��( )�nS8��ik6(���/2��^O�lW�X�?�1����i#����Ш���>�5y�� S���Ip�r�5g�3Vi���1��x�v���-T�QR,�#��%�U�eb���n�lWKf�%���r�m�1f�nEV��N�mER�H�M]�2��h`��jܓ�#�=Kl�sv�j�*,�y�PS1���y��ڴ����R��f ��2`�"�f�������sB��kd��x�%<2�u�[�R�[�V�/E����M;4V�t�q��Y7�d�0jr��3��&Kz�d��qkݫl����aB�Sq��&[f�P�и���qE�U�Wam1�ݔ�|r�50�Օ�$B%�K�:բ�r�Ek���fhaB��z^=��ޱ�kk�ʒ���f�[eu�IA+��5����x+o!��)��L-�	 Vnk�a^j\����W�[� ��zC2e��WF�^8w,�(-wm]]n@��3��㈭iQZ�7��^��V[th��+��lm=R�te ��Yj]���%C񭩬Iu���!Bͫ�m&ͬ�y�70ֶ�
�f;:�J�v.E/��	���e!liYM��6�Ю��p�^�QSXμh��-�U-��4ֱP�k�F�n��r�1ڊ��́d&n<Ou��U	�S�W�m90�
Y*S��arм&�Kі7n\H����!f2��1Nm'b��ktJd����>{��v��J�&Y�JAdWy[6�܎�l��4^�7N� �70�m�զ��`���
��j�+0�u���W��5[�a6�L�)D�J��
�)n��`�]F�Ǘ��]Ч�VQ��Al��s�1A��:t��r;wH�*�)�Y�U#*�u2Y�twb໢Ȧ\nM�*�\�)=vټ!���=4H��@/�E*�j��'����*�y����Ee"UBL�o1]��w-�7ݺԜA�� PfҐ'�5-�wQ��$�҃���
����WrÄ��*�dyh7W�u����x����u޴YOe���"S{�%)ֵlޔÖ,4Y4T����iE�Wz����(�w�c�f��G$Ԁ�v3�kR�К��J��Vj+~c�K­7cmN��$��T�Vfm�YN��Y[N�8�4��@i�]D�- �v�.��MY�)�P�K�N�
ge�P��;jP�6�[٦�T��U�,0%J�J�hy2�]�Wyaǡf%k�^;�����'���v��;��e��,ͫE��2vMw��U�n� ��Ti� ��oji��,ctj�����FkC)jk2�cyQnh�f������LG(���� J�Z5Mn�ȭ�[J^'��n۱_v��Ub��~< `7D��A�-��vE<����:�m����B
��J�"1m�ŵ���gl��3��fź\q�r�*�8���z�r��:[aMq;�^��ѻ��L ekL#����z~�$�ڱl7����7wP!��[�
�4.JaWr�p�Z����ʖ��&պ�m��{�R�%�w^�W�Z�,�������ձ//&���Q��;�Su ��N���
kK��A�~ل�x��U��G�ij��r�*X�ԷpѬh���r��l���ˎ͚�ۤi^#+��BK��NE���쭼��	��6K��VР���%�6�Y:�Xaђ��-���E�oq��<c�_LX�N���\Z�贡g19{lK�s�uzSJ� ��n�H,=�2���,ı�ml%5t�����)Q�C�$��N�R�c2� ���[�(o5����e8� F�Z{m�s2�����CU2�2��#��F͌z�bݢ� �ي�a���3�St�{����$�'��C�2�g�ڴ�Cq�
jb��k�W��`��� �
��0u��s$�/eI+#7�&�w���6�ECb�d���3V45�3W��Թ�\r��5����l��6�w��R<v�ԍ�L8��=Ҝ�{���$͍˺����;F�sCdv���K܎ؗ�\Ą;��F�D�w@	ݶ [�m�r�a�U�3a�ά!WŜ=�XI� ��jD��K����d�*V5�j�@e�*��&�w�ZC%-���ncMl�{RV��@�-x�$��c��9t�5�-G�ڴS��$�Z���։��6y@A�:�!4�e�ՑN��Re,Ɛ���{kcl�K+s0Sa��W���e[X�)a�j��	a��.^�C�ƍ7�n2(YB�����Tس�*I&�H���0�lJ�N�;�Y�^����Zbr$v7v�6��c�B
8��[z5�kM�
ē��v�x��	���+�jP��#Lwd�N�� W�����Z���e�D=�&��ح�.(@vJ���J���]Ez�CfXe�t�iX�ţ*3Y\��P�v��Q��3+��8[3q�i�fȗ5nj���3
�S4N--�a�J��h����)��mj�z��4�tu�-��h�ź��x�0	L��&V�U��MU��y���F��ަʹhCa��H&�H���U�X�֚�VdT~�,��T���j�`2�d�� ���w+&�L�T�4ҏ@�ji3��ь]m�s3ou�[7Z-���6�
g�݀3)�7�kpV�c2�c����Y+;j�Sѵ�Gv.�!�*G�Y�C�QeX:6��%E: Ѷ��2 n�;�"S�o#���E�=i��n@�V�5��V1�-�.k��fl
���V����,a�bU�af�JRQ�>d�S&d/i��U���b<��^����Z�F�����҅����̕n41�A��b�����4��ʓL`$�m��aZc�L�أ�u��kl��P.�ĤBp�n��!VY�xjJ�@��� )m��Ť�6Me�X����������#`�˖T9FY[J0��f��(,�̫$&�R��b�� �.��2�&�[o�N<ӶM�E<�-%�l��Z۔��"�@f��M.i̠h:��4�n�B��sh�W�*B���U�[�OL�)�m*�2�$u�n�i� TMYE�S�1��p;ۙAe��������Ӻ��T���<u7&5�R��$�A^a���\��"Y��H���B���x�����(twJ�����pKߖj�72�+ƆkX!L�M)ӇMkn���jf�f�xB���U����j�YD��������Jޑ���n���6˰�d�ssEr�`l��Ժ5s80��ŗ���P�^�Ðn��U�H�Õ������S�$E�d�ov*���u� �BP4su��-�2�;�]`^�)ǎRX�iJ���Rq�W��*L��+2��W-27ƷuEvY=4�k/qc�wZ�����)\�Qm1Xm��d��x�Dm��mFM`[A�?h���V���LK�,�l�%�~]l�&����R�@Q3P�h����e� ��^,R,f��7��&(<�4-ԛXQm��#���2� ��z�.JzlщU5����K�P4��\CyN��2��n�	�n,�tbO,9��������ͨ��C@�ܺ�A ���H��ux&�Wj)�A۱#
��D�i��(9����B3�:_=O-K����Nj˺SD(�t*��VB�:{��q��*uxI�F�����i*�`i�R
#n�U�Z�j�T̈�gB*�^�m-�X(+��0&;w�q����F��R�]c���U��`��[�
Қ�c^_�m�#X��s�����$3i�K5��=�xN02,1Sի ����fӅu�@� �{�ݕWn�Y�۷`�B�eDU�t�}���j�q� 5�
Ϝ*K!㽨ص-L;V)`Mzc��[d����qCl;`]:�G"v�t�p`�n�Ь��Սƀפ�.��J:UMd%c̺֕ѱ��:g3u��k4�L��5$6�҂7�.��5��U!e��V��E!Iʂ�

A�@��[���,("�z�����o4����Fo�c�-n��@]jR�z�!��dsrf��YJ�Ƙ�z��ؤ{R�pS�LD��V�t�J�A��c-4�V����Rˠ�:&��5��9��;'L�&�y�-j�\���gL��ª
����P��)୽L��a�J�N��!6�jS`�!�2�ы�j�Vҗ�Uǅ"���FS��ֶ1˦\c�}��9�Z(�5�uՈ4]�6�L�@K�d���Չ2aэ9 ��3Y��aQlǫܺ10B[d1��d�YHPYwuK�����2�f9P�+N���Q�*�;@+5"�慘�������X��s0�٭���$�u5"0� U��ѻ[��@v��w�x,�,�%0L����Z�Aݥyq�CԞԣ�n�
�uZ�B ���;t�M�G�D9Ԇ�r;�h�)���AL�Haz5|���ˢ��	0;P�,0&p7/���������.��}ԡ@S�^m�
�L�i$�b��54�i21}��d�juS/^���"�%	u�]�V�r0�hv�BF�Yr�)F=F�k�V@�V�cN�O.mZ�
��҇)d�ͻ��
¨b�����ݚ%��1�3���u�1i�vҽclS�o#�ᔛ��m���9��Z/mO�%{`8�q]j��}h#U�M�6ʱ���8!��{B^X9D�EF�6f������*��O��̐�Q�c�j�K�O
32��2�[af�S��a/]/��*����5�I"�B��\���4��r��N�:�2�k/]ȶ��N) ��F��`!�ѩ�٩��l�&4mX������Q���mDvw������W,��ȅ \n��4�nSɊ�%Mʘ�f��5]�wV]J.���[I���Jڽ�;���n���t���g�S��/F�rL�&�5J�>�0������e+�������e��KC�SÛ�R�e��TZi��Aۥc.��ަn��4&Nii[H��(���q"0�j�2�`5���Hf�0�Q�v�|��[�6���Pi��[����e(Nւ$ɤ漽��R�(0GaTVk$�n�b�������ݣ{�V�Snհowim����1�oC&Y���xaf����Қ���U8�v.SqY��hmޔtMY̘�aA����d1!��Zb��B���X�:�rU�o� �:r���!JR�t��@ى�����T)�E/����{ �5�Ih��^����`�f��TrRۡIDͽ��
L�<o)��@h�[�����C��J�a��� i�'4���Q�KwQBT��/0�ک[t��@�x>3pXQ�i ��p[U���Ƿ��n��'�Z�V��45��&vl�#2n�y��O�hVjk��DɘL�Cs�� 8�LC%̏o��_1Y��WWNi�ޝ�ܓ%bw^���U�����
⵼�~�j�Rj��[2�Αը�̽�ԝ{�2�kТ~��h�n�rI���\�׾���A��0&�u9C[�ʊ��X�U����
M���*[&�����w|ك`I���'�V���>̗ÁjJv@jcV,ڛ]J\֊�*�e�}`��.l���X��Kzi�}#Z�,�����9AoM�!���ǧ�ib��r�ُo2DY��#�3�vGx��^�OK�:�����m��ݚ��N���v��Y��}u�Re�Iu��-а��F��h4�:wZ���m�8�:�:U�Pv�`7���팼vg+�jk4�^��n�oZDf�V@�������\��%�-9d��j��3΍��̔�Қ���Pe5%�܏FTp�'���u�"��7:�L!�$�s�\���t�$��=�N�n�V�YLj��E�{����E���QD�^�빻lq1�f&�r�άR��ț�z�}}���׎���3���=9>�?�$�����t��q��/��lV��]��i����/.D��I3b��¹#����sZ�����Д�'ίt�p-�Onl�Έ>��#g����Z�m*���3�Ft�
9`i䥜��y4^+���ggD/cN�}���EV���ݛ0���jv>�EN�o�GT�2�m'���Jm�ˤ�ufkڛ�҃.b�Q;�F��&u��!v�d�LN�˂���w��u�pb���'Kԥ�1Ǭq�.��ks�|T���	oi#vh�|�]��Ó)�����\���������d�<�Ռ������<w�������]Ǔ,�]�aW?�%�b�t�a�Qte��Ӗ2��G�V��R�^h�(��V'�H�+� �o�R��wD+��xj��i�F��*��d \�$r,��5�T�0
����)���Ұ0G���RG��ݻ}x�n�8�͛�!鲕J�]�I[�2���S��H���H1���U�#�Z��:���O6tX�#wg�z�=��ԋ�TG܂(f_U�=%eU�-@A���#}���ޗϖ>������'_grVFtr�9�̴�y���V��s��(�s��S����`��a'�,+ݫ��ٮ����l��j1q�{�f[�1s�H����7�������-���c�.���g�k�N��jne9��#dH���!Q��ڶ���7Vwh���k\�K��X�+�a�W/��}9y�k^�a�q�m
�{�\���[��p`G9eWXn��\P'-R�x:�wp�:�T�ڟ1�[���:�ʘx�:�-=��g�b��6�U�;��eEW3�SjV��yw�p��R�7u�1]�=v��3�Ղ�c���b��ܩ%�]B`.��˄�w>���	���1J��B��6�mb�ՃO��C4[X���:����x���fӏ�����]i�ྖ�7K@���:��ȗ�P�ݽ�h%cf� zj�f7��.Xros�Y{*�A����Hs��ʇ<�������e#�մ�b|���h�uw�JR�p�h��\�:���\�Z�".[��)��V��x��W�m쭃vz^n�ֵƳ���MI�u��J�+o��d�g!j���+�Cqݔ�I�%W_R�SɜP+,p8kՏR�����Tj�J9A�E�fegM���:��0�������J�Y�h�b}c���U⻮�g��ʒ���FK��"�@�b�T�M�%��j�����
��6뺺���o�.�
KI"��g�'mE2-5�s1ԣ����6qGG@0ʶ�q�i��.�5���Cm��,���G�:��(9�mw��0ӂ��Uk�}r����P�
*��q�r�!Ӧ��eY��%��V�@t[�ݸ9f81�7��{�+�'�d�)GZ��Zhv+{e��=|��4N ��_t��H�,V+��}H��Q�tvr��ܻz��̖�cwM���O�9�����MA�NΫ����+���q�[�&���eVs�����]ƅ�2�#7��7mF��WIZ���$���� oÝ��x�Mh���ۃj�TԡX��7��C�����%��l塛a�nH���CV��ض6����
�x�\���
�j�����kc2�2\9��zmY�s�a4�I�>`d�A��Z�*�Y��t�hi���ArW[�@si��3k(&0���x����SX�t+��WR��]f�+;��q(XF��P�2��)Xv5wP��#��֬�hXT�����&�5C��4v�[��y��D��&ف����n��rA-��=��Ni��kt�,^����]�T{}r��vxց�y����,�hu9H����Z��ə��KG8�v�������i�1Kڀ���va֮�J�"���}mn:|�hu�a��)��p	��Mto6e���8�P�G��[۴�4��a��`9ܶ�y��4�m
ΦXV���[��3��vqǑ�d�ml�S�I��^����� G`�.�<90{�BaV�Q!��]wb�o7�u'r�˔�y���eգ�V�^��ŝS�� e�V*��0�]��׌a��\�5�5ˍqG��v=s]��qE�n]��͡u�=�L�Fuap�Ƌ4��9>�ޣ�����~��<�X��ҟ-�o�e��B�IvC�У@���J�\��C-�9ׅt�Kw0WM똵��+�ѫR�T2�U��ӹvwT�s��<k��2�w"5}x�]�u�!b��C�gAH���Z��� %oX�t#z��W`����:C.챂09k�uY��n�)��.���]�Oqz,b����K��Ң���`��W�̬/0p�:!�oo�,T�y���X8:��m���A���}�m��T���K�k
*^�}��6�N�z�IK3��dZ)�fe
�᫭�VT�G�.�Z��p::�B3Eu<sB��v�L�ܳ��"���K�J.����v��K[T2�|��W�v>u`��K�h>c+1�r�v�ʵMr
��Ӣ�g��${(^*����D,f�9wck�Y��!>QJ�-v�dyn�K+4��4��إ��.mZ��g���$ڳm0W4�СK9�NI^m&r��|��Wk)����v�&�^�)�@��[�;tcq����v�c��Nٹ�^��a׈�`��Pk�i�c�t�f�ݤ���ӌ�dj볦��+�.��Z/9F
�yP�=���܅�p�Hn��a���f����)9w�N�7W��ޞ��D�ή�"��Pep�bR�8�����	2��:�_ˀ'+�`jM0�%�\�6]�y����)�v���1�0u� ���wdG�a���Z��:łZ��{o|���{7z:H;�~M3�S\w��n�ôl�Lע&�n���-Z\G)��wok5fv�[k�޶�
\�Hx�Ɍ��k��jS,�k8!�Qsm�����X��8�Y� ��+E��S4G���+��E���{�Dp�`�v�+��a��!Q�Lb/��D3vQ����C�QE��;W�퀻#鋣��Ooc5t�OI��# μ��L����*J����v�u�S��{;;�:�2���ףeM�]�u�r3��5;�����`�Gx��S����mN���ܕ����q�G�;��xA�a�5X�ܺ��obKzn��i`Z���L	���`��E��=�kט����zsB�iH��kk{�b{Fov�
e�b��RU�����ԇl�y����s�Н*�(ko�vG��rwX���1�u=��h�v�R�\4P�&�����\3^�L��B�4l���T��|~�.�195��*�=]W���TPuH-;�|�]@���=؞ݜ|���/����΃ȷj��Y�����*)����F���rqkl;e_N�`�����m L�)���A��1@fu�s9i��۽�˂��n�Ⓑ�tjņ^�"�T��ӹ���g_Rd[#�/ڹ�[|����P��Z�H��_ �oJ��
&f�*�T�j�JΦ�h�-`���GS��NB<�x�*�:�]Y��T�Z�au�����*�j|���<�(��f󊽫����yR.�.J7S�`��x�×ɢ�u�{F�N�s�ޡX1����-2�����	���:Ƣ�>}O�I۾��e�q��V0u^+�'�+o��N����݆2��Nr�}EQbcT]�z�,<=X�I[��̹]�2��h�h�D���e�@ň�����1l�����ɝWQj��*c;��8���}&�ku�K��pCPs&Q �p*T�N�/c��o/���g i���
�]]��v��b�JXQa� v���r�n�1��r�(�jb��
k*�Y��M��i���/un��a��S2�+��s20f���/�^��:�����ܜFڠTtn,������[��a�ؔ����0�a凚�.bɄ�Sz��`񙬇���m,	�>�md��[Ź��O�wP�[��#[�̷�x;n���>�m�㼶��w�E�3k@�9�,��r��؛ov�r��T87,�}���7:���M�{3�gwT��;{9Worq+:8A��[�s5�J�	t3���z�K���6�l&�OV_|���A-[��T��2jSD���������S��n�Ւn^ ��l�\�1��Nr��������s��ݿ���U�7(W��uٹ����l[e�� ���DT{�n��ʛ�bӖ�3��u\h�4me���KK��ςIʝ�y��J�4c������@g8�[�ű���V
/#5�ekY�|����5��;��g9�7mٹ�oPz6�'�(U�
��P��Ԛ�`���l�>Rf�"��PY,A"h�t�'mq�I�IA���yg�Nq�@C��ܧ�[Z��q_w�k�Բ��j�eK�6�t�nc���go=h]b9B��Ogj��hnb *vk�R�-N�����r!.2Yό�{B]MtH�f��e�l�\헝En�&Kݏ��;/��qK��,j�Χ�\�Ԇ�%�e5fR�}N�.�U���;�L�K�b\�o��Y3.��1����zs3ڻ�έ�gk��"� q�B��Ub�+LO��]��o--U��V��\��Bb�M�Wm�ٔ��Ks�B�_e"�[����;کp4�� W ��mH�'d��۾�Yx{}�d��M3���n�,V����B��|�ì`ݚ�:��cO���%�G�'�B�g>K��%�tDK,.Y�4��0�,mޜq��x �鮄,]p�8� 1���i���c6�Z3XT;.��1!��2�p�Uڭ��2��Z�@�ÚsH��-0J�ه�Tޫ�T���͗�w�	��b�h�|����\;���.�.�חc5K�|�>j���
��j�2;���]�*���QiarL:oI~���ךZ������zRI�o�����(����P��
ؗCQB$nG��7���fRB:l�Y��Ŭ��7FM����/;l1u�D��a��\�4]��0�[����,Uի'4���y�|Eˆb`�y�>�i)����[�����CMt ���� @WR��ݚJ���}��J�BHr��g%zW+p��i@��gq0��AyO1p��]Xz�u���(m�Ui�ʘ���]��L�O�`��T���l��e1��ȅ�bf�:��8�X�����֍H/�9��.�U��}���g�4=ް�gXQ�%C5f�܁��t���(���|�j���\�X�ib��ԋk�5܏ӂ����)�|������l�|3sY�yx-���K�7�oZ��6\�9Y�=A+�.[�V��[繗D���=M,eE6+�c���Δ�����e�fؤ]�ݳ6q�;��z"��|��c�8�x��&�MVKP��f�mլ�.�+����QѽKy޵��}c	���[��n��j-���<��嗀Q�x���q�CЖ���A�ø彗`�ΨN$��m�q��:�ΌiN��[��/e�4�)�����:���_=��������uԏ�s���Q�Ļ�A뵜�RR[D�`��9l��O�ǫ�I8K�a�����c���0�T5�Gj8h��m���J�IK�P�ub��~.�n�s9t��]�ջٸ����@�Z�b�9�����ë0�][������vK��ۖ��*�&�2���^��D�3*g��R���V�Յö�ok�Z���^:[
ϓ�yA�v���I�:f��t6tʹ�zquu�&��ʲS�Cr�a�z!XsWw,�\�N`AV�SUZ�8�N�����	ak�'Jn��s�X7�V�\�pF���Z+As@n�r]�V{jꉛ:U1l�fwW<pXHކ��*sé���3�C?>�p�ӈf��aq��y�q�q��L�-����
�jA`���eǽ1Է���ѧ2���o4���-
���1s|���F��7���gS��A�Bx]J�0����ֽ�}�ٲ���&��34�w�-��A����Ã{��u�>z¯5��x=��ȓoo`3����X��'j�:8���Ksj���/�;�e�GGo��u!.�&���v����ou�7���>�N@P[�.W]��R�M��K��x��Wsy�����SoJ�g7ۢjvT�U�J.]�0��>=}��+�j�l<^J=g�����7�NQh*��\)����ˑ��ZdfX��YLb��/�S�]dL{1)����Y8Z���ui	��m�ss�����yۦ��K���y�lv>lY��		�	!I�ޟ{������_��S�7�����{�bDh�ƹ�.h����ޛn�������W��;��Ő������[��wC��|�S"�����a�F;,ܭ#�;��t���=�
�h�D�v�@��X%:�{"��h�t����ӭ9X�K���\��#��s"�
�����4F�������݌>i�����Z�u���	���Π�.ã}�5t�v����_jķ��<�aC�i�:qe��i�z���;��:�'+n��7�1���JpC�)8m,}��Yݩ��n�\�+yGjeG/Ha�J�9�MX���1wR�����Pߕ`��ۚ5��GuS���,�8�xc�ge�ϒ���3mqȥ��
愩� �;'N�V+F�F���;65t̝!��@pv'�;F9S#y� ���i�M�a<>F�87c[�Y���@�X���4��)�!>����42��"�8�Q�!±�ڽ{���%b�˽&ٸ��+s%��+Tw1�[��\�)չk�ĸ��u���&��߯$HC�u���h$g>֦�քA���I�I��l�����;t|0���l��4�&��óQ��9����Yn��,i�On��4���S5�];� �^4jY�9�6�xef���d�-�*�2��K�Ų�h��Z�I�|{NA]��U�c�l�w2��i����v��ݧ�Ռ��{��UjydwWש��;�_�m��_�pf�.��s��u�J*c%m����i
�X��o9���vuf<�3�܆�(�\���evS*7�q�2�!�p�N;r��;��.���$��L\�W�-�s������R}�{ÃA*4���V��3�\��~��M �xpgc�-��Ά��5x�$&�|K=r\�]� Ո���մ��Ņ�y}��� �Zc�fM�����|u���;��d�N�bZ{���iv�
!-�w+�}4-�}��\�]¤0�E��+��m�si̝�"�"��`z�>t�: 
[{��D4Ŧ�]!�VgJ�2������~o��0��-�(u�X�ެ�Y�9F�Ҹlhi�O�k{�]e�<�l����;O�*���7�*���j�6�X�1 ���"��C��@b��s��1}��^Ǐ����o`\��7�MU��"�b���_sU.��X�u�(sU�G�E��k;i�����o�7-Rmϑ��f�I�.C�]#8��a.��6��G8_�ۇ9�̯gDoC���PôR Vs�4+|2(� ���Z�˙PBf�Dx[6|:(6�-(��q�׺�%B��J�K_q�յ�5c���=�<���湁Xj�t�gC�$�u��p6�*���hE@�1cc�uX�+^^e��+hE�YE�	�Ki����b�N�t�n�0}��:��=Q����E@о����7��yoM�a�y ���t�c�o�1.�a�|dc�y<����R,�O���3�4�D&�r]ur��Kg]���b4�\�V��`T�J���"v�c*b���u#Z_�*Gr����h9��xi�^��C��{�Xh�����x��ˤ*n�u���4��jp�+]�FA\:�x�ʗX���Cע���լKy�#�Ź�M�^����6N�,9h�9��Z8V�Wd�׸���6��7�(��Bv���k9�Ҋ��t��1��9��Sv��ûS��� �+��v�=��(��,�K]�8K�D�c�ox6�n�.�N�+?d���]�]YW�S](2	�)�����ɖ>�%�f���\���>;�x��_�[b��I
�*Eܦ�Cc,@��J<Ayх{��zx��k"�:���Z�\j[���]�g��LWe��b�Xdr���T#��Yj���sx1>��Õ�k�+7�͞��)֚Uݻ����A�+S���^خ�D�}eZO�,��#V����h=W���)�l�R�)@�*]h�*[:@�:�:��̵��-t�A�uu��W�v
G���uK<��ݬ�0}wr���mh�� ���
���ޗ*=�R�tݎ�(����g-0��/���S�v����+�%]h��en��tC�'��.��:�SPmX� �Y\�B
Ea=N�Ά�w݈ʳ]�g�E,���T[ܛɊY�1�B��:��O�B��2�p�g��+@i�q�L]�̘o4$WY12����Z�9^Z}�D��;nes���;���9{M4�e^9J!.�7mDi�+��<�L�3t;�>ݡT�f�4ƌ�¾���Yb��F�wLg�Gzi�Y+��22y���n��򜡤�����ϵ�5��r�8�J3�M=W�-�V��Y��*I۷i+d���w��f�ފ��j51�hY�:���w��Qw6�%�@��!2pĈ�l���GeLfv.��i�Բ��]p�X�Y"�j#�U�R��菙]���|��f�+%Ь��>Y�ҩ�Wu�V=:&�xu֝B�GA�����CE���E���-����u��v=�Be�v0eA.���1ҰU��6�U����Km��tm��
�P����*�(mjͰo��4�)�Bl8 v]LM]�i��s&PY���
�q�q啣�0*��Z�%<��������P��0�Ul�"�����N�ck�K�5���(u���&Nv��9
L[4`��ǵ�nG��F��]��Nn�o%f���i�`��3�펀
7	&�v�j��K�͖+��*�+�J�8eh}���#fӪPn�&�-���i��y��60��Z��l�ϩ鰝oX�T�Zu�O̏��əQ[���8"V���6���A�[Y�#�L���	���M	oK��ה���4觙�E3��u�KQP���^ȫ��%��%X����9�yb�<��L����-CL�1=�)��D�q�P��՝(���r�PJ�>�AV*�'W��h,e�{�^�`�v�]�-%��3X�s�fl�4�@�Σ�ǲ��k�2��B�]Ӯ�B�ͤ���٦�З��짤u]ۧ�hn0��!|{(�tm^�{����b���O�n�ou�	�j��=J�]�O�<�Z�)[��\u�+/�H��8qsT�םy���n�+�`�y�GC�N�u��ޡ�uA|�>.�^d:�e�Q�&����]���W���҅�f�r8]"���ǫl^fV`LI�.XʘAx�-�5�)=]�JTř���D*��
�qp}��νj�^|��9��L�ŵj�fk�p��)/�/[�3�Q�؇!;v�e"+twɪ�4�&�t�M�W)h�I�t_pY;(��M=ʥ�bj�kD/)ۙ@I��M��-6�X�7a��\��qa�҈]�v��LϮ)7GnP�ӕ0��dP(�4[-�èJ���ܽ���] �x�O����]�,hr2�4��!�Q����� L����X�Of[fS���:͈c����I�Ӭ�K+"�W�6��ֳ�9A�_$�S1"��}װ�:q;���z���z����e�4���˛hѓ�Ur9Lw�krp�d���  ���4�s}�j�a��6�����ו�N���<��"޷��M\+u��6I�]FуL�=H��Z�O���Yƃm�ck�-�����t.r�NR�z�F�k;��H��"��GҰ'Da�N쥠JT�W��������V�T���PT�u��ҁA�>�;�ؖNø�T3f��ڶ�Y��)G�l3�,�g��a�녧���H{��ݏ.�IՁG�6��B�k���ȩG)���԰�U��lw}�R��O#��H�^t�57}#T���k4 ���G(��J�����2\z�<����C�ш�t�����
�z�W=�Դ���b��l鱶8�ai"�y�k�QjYO�j�b��K9�Z�yQP���I�e���l�4�Nk�*�w�8:�6QK{@��oR�FE�G���M��`�Q��b+�.�+����^�8P�L�7/����U0(���ʹ�w
�bB�c���U�J#Sٴ����S䔼�%G�j����Y\4_/��p�+
\vs��]]�H:n�
���:=F��˻���(�U�0�M����t�g�gfUq(�v޹�rx�mn�&COWP���4Z1��a�b�,�%�z+	��V�,G�YkiA�MG��p!���L�}2N�sU��Kr���7�����>��\�i�eE�Vڛ#w�7m[ŀ���5O��_^:���;���B�zz��'0�i+�m];���J�٫wh�����M��b#�Uĸ�OhT!��x5�ju��V���1k�]��}��a�)�b�=X�闱VR����:�Sa6�-����2��n\H%MOf�O�M�J����Qn���i����ޙpS;��5�o�΍]�}���%��g�;��ڌ�]�n3���1�vc1�d	�Q��.���y]���oox|�;�#C�<&�p57���V�"�8>.�
�޹t���s��k{93�P��Z����{#����P`��b�K���|�D���Z*��D^�"�N�H*�?*p�s�q��M4���	H1���*jX^��30eqL��i��}�!c����Ȧܢ��'0�>J������ɧ{neB8�z��x�q�eCw���Gu[�s�`�����|������1�������է�'5ip=��;\ZM���x�;��b_h�zh��̨vu�+	��5{�3X����rJ?5n'�r:�q(�v�>�8�G�b�U+�U˯�u�1�Z9�)�򍚅�XG.!��.�U&r1;��u�ei�#ʅ����D���_�*�ۜoy��(ؙB6�l��1]K�H�-A���!q���r3ORY�[�|a/&.��tnc�\��'vG�+��Ĳ�R��.^��:����,K4�:?���L�f�&"� ��rR�w&³���{5ͭ�\F���o+)�rg��9��i{�y8:��3���@�p��r�E����<��b���k7r�?r��ʭֲ��cua�uwfQ�m]s�7+-���:z+�u��g{���.G��č�2��������n��n�he]���ZHK��
E�.N�z�l�;#6Zƈ���&AX�xOv����%���'���UBM��"S��`��l��ef�"�y	Yi-�p�O�F�,k��~*��xiZ�� �kn�����-m^�5���B7p�5�&�m$�QG���*�r� �oM�տ�,�]19����w�.-�����ʺ��}yCi��7��F3.�ܐ�uM�U��%t�$9ʕ�O����vm:{խ8Z�
0��s6���y;�e���wdU/��c�-�)U�J�$��*.��_�wD�S�y�PW������2�%�cZP5ӫm]�`�ԗ�(NO�f���B�u�.un�(i	��c�����w}eQ��
�����tdyH���:\�t�ت������5��}I��WA�
M{r.���ŧ�nRأ3-ӵ[�p�]�J�w���â�����o�}����;���|�ݘ4-#�^�
Ư�E��'O�E����̘&i9��Avm �r��؁�N��w����� �/���t�ܕ���g��[tŦukY�1�i9
���ڔVeh�qM�y*��u��&@%P����BuM�3 Jrt��mU����M�A��Ȫƣ��$�������v&�IJ.��B+n�w�/e�@,�i|�
읫�~I_��mO�����=�k૓�E,WՋR�Z��f�L�C$�rb�dr�}4=��ۘX}x��5F̔b�cP_m\�ѩ��I��!ڟkHuEwY���f��m��52��f��\sf��)����U)����<�M���`P{���J�fbJ�oq0���K�bs d�jSt��t�p<����k�X�.nf����4��(�T�j涏�m�Ǜ5�3x�A� �� t&��K��<y����az8���l�@������ǣ�Vp�����+��B��L����=�Es�i΍�eKi�Ĥ�̈�utT!X0�\���>˹\,ZA�A�s�7A�z�ҧ)O e2���ӊ*�E��A�*9.7�+r�4�j*Ƌ��5G	��K+�V������E��.�x���V+�pW���;ث��i#�����]�sd�5��ӥu��/y+!B�r؛'���p ��'3S��(`�M�spL]���u�(�#y@�$7�M�;�P��R*��Vѹ�Ī|w���!F���;M�S�Vs�Ӝ�e �[�Kz�,Al|�Zb��orm�l�i�������ѫe^���"����U�@ݦa��ͳ(Ι�����ҷK��VӃ�Ti�zP��&�6黝��aU���9*s,kp^n�	|"��{�f[㯖���5>Ǜ��:0L `�3ٌQpW!᝽E��^"H����.�Kuu�scCV�MX�7Ehr��:�7^��hV�mIIgq��g�E9�Kt��%vF�
����4��f�֣��h��J�΢��x惊BZ���s�۝�Y�J�������#Z�.7x8Hf�|GAϣ;�;yZ�X���x9��D�kQ�f6�Q'.��p�f� ^5.��$a��QZ!ʇy$s�:X�V�rZ;H��+�R�<�O��j�⺉�c015��AYQ�%���4��^�Ɋ��f�އ�D��2�!���3e�*��۸
>6݃Gs쌹��T�s-�:�Z�PT���a�|#z�|�kX��+
���[9�b���=ɮ��Fa˕�����q�^�� A �D�z3�k�R���#a�����m�oO@wB��/�/
ݾ�s�My}.��ާ;`}�:��R=�S��2���0���ª�gPf��
�/T�%�k�	�(��:�G����<!*�[)�m�G��m�=+r�<�B����mf��8(M���kx�P�x�������k��ܲ�G�)љ�bZ[��D�s)��];�y�i7�K����8c���1���B|x��=%�[��W	�z֮C6��y��h�c�]w�n�v59���U�j���R�H�;�B���I���y����Q�{Vq��.������^,��إ���5\��'���9dL(L�ؖl=���6:�u}��˛����k��1:�x�V�'���hw�;Ü�u�r�w|�$媑�.��7m;��2��9�y\%�2_O+ˡ��o�<�~�~��4�m�r|���Â뜉9�����U����vc���p���Y]ozazX	*V;O
껔�l�ݑ4/�hfw��u�}fʌ�q��Q�������Ղ�f ��#�k{LMJ�f%8FY���-냒��0��;�����v��gR\ȅ7D�N���Z��z��d&wٚ���_(;���ܟsS�^%݂�����2K�r�9w�JT�	�g}��G;#֩�����O2����vq�`�@�����l�j�ӵk���љ����y�G���E�"�eB��+%F�J�U"��"Ŋ-HQ-���āSX�	�QFJ���2ڰ
ŐYQ����f$r��mP%H[BQ�Q�R`VVC�b�YXAAHE����XR��5
�E�X
5�ISj����V��,
��Ԭl�I�%b�(*�[%J֤�#!�0�%H�1$�̤�*)��\F�E��iPSd�Z6$*(J�0��J�"Ȧ0YQej�l�RVLVe��
�jŐ�T��T����� ��,
�d�LpE%j���RV�-�+XTd���PU�
V%q+��TX�
��*V�`V�V%��X([d*���dR8�e@QRUj[�&5�X��8�51"��d11�����b�?|��-���4Z�|��M*��N��;Z��B�L�\$�%���į�=��M��V�ǉ��y�KL9�G�ZW|�f��+��n+c;��N]!+�a�t�[�5�.�]�݄nj�n�ny��.�N���g�qƱJ~�����X&\���b/��I5��9����f�}�v��]N�on��.��y�J�������>�x pd��F|`��R�T��|oqﲥ�K=�_�X�|k$8{�rz�fB��)�O�^Fl`�S����;ĠO���z�~�{�dw����ZD5�u�G�a�<I=/�@n����s\�r/Jַx�����qc�j�h�l�[���{�B
���/��L1�/$��M{�,6 ��P�ػ����]{��m#�)����� U���מ��<�|V�������մ�w��bZ���h�F�'��tٯ��2D�{>�Q��.��;�Tk��+��r��^dZ�� ����{Q�젋I�XŪb����	ũ�.%Y�4��Z��O\�`_��{U.�����\����חMa�|�_�V�o�zP�\-�r��1��ˬ��p����� hE��t�YEv�d�^^_n���:O0���]u��Z3�u�=���F�9������E8[ա�[I躳ET�ro)b�{��k��� �j���!��12uP�f�n�)үt<#������,E�w�x5ԥ��T�5���pnw��_���͎����3	_=�8&�J��=e��j3~c�`�|��q�^��֬y�!���K#~		%	��Kּ�9L�C8��7��
f����)��x�{��*W3�6	tF��t�z�0��}`��T�-��p�ؚ���dM�+����%��MO�1<��a���	b$E^�&
@��{�7��{x�ޒ%�x�0��H@�1JX��޸��3��R%��y<9R�r��
�1�9���ޗ��y�Wj�D�fqyb��g'fV	�Drǜ)z� ��=^!\j+�l��,��t�ǳ�̻�< ����
�{���ڸ��]3�s����*��<7���Xj�����$��ޤ�����@v6<'�a�p���<3�G���0�׺�χt�I���F�a�0[�u���ve3ِSd���qUm/�%)�8f��T817��*]��K,�简���
���:~=Por$���"R^2�U�������,x̻LU�^��"��0Y�8�M�M�Mo
�Mr�w���6!�,n�Q�U����Y2��G!�i�nV�Vε�eC��Q��gƳ9�����}�x&I��:��S3T�\�%�!�7ê�����N\r2����j�k"����5S�Ź�:�����͔1.S�n�mY/!�QM>�յ5�Tw�5*�)1=��:��c}�	�b���}y+��q����`�Vr�¸���d>������\*�^q���u�Z<8�!��k���{���^!�ف1�+�ʰ�u�o�J�Y����-���/���OHwW|1���ޭ�d汊�j��XV/AC���}ܭ%d-p��!޲�9�_8_#��r3�;'�%9���
^�v ��*����=>��>2�Z=�	�/ �?kݢ˿������7�kr����b5)�z{�]j5h�&���:L�-&:"�q>�6
����wo�k���V�$4L3IM�X�i3���ZG*`U�E`TN��j��v�s���3f'�������2�o���*^�
ݩ��]-�/�t�.���z"2�^�j6w�V�P"��՚>WP��y��,tX�X-�4�K�BM�̩���.�!�kX�B��T�=撵��ħ���N���^5t��r>��GY�2\C͉k4�ry��˼��j$�:�*%��u��O��g��/�-oBnj�f���{ZM1m�2Sco(}æ�s�����\5*�*�=(��z�oh���x	8��ǽ\�:�}��Y��8��D���L���9��^r�	^�@v��06�μ�R��q�`�vߖ�V�������A�&���ȵ,�W�n�YB��ͅu>�3��U���4��BŞ��'G�X��3>�ǃ��Ck$���q	�`2�$�,��0�߳:쟬f���r{��fΖ�^�6��I�p�y��&+����r��<H<[�K���`�G�~�7~���s���!=����R(L9�%<A�<��=��2Fm<�T�ΆuD�v���VT�X7K�/*ȇ��E�Z|+J{E�-����<5�(�q��=%!^�y�;�Ry[����p��ܥ~��k�UY��Y�Z|+Jd�Z���#�k��8!��T�^A�WK1*�[i�=�r{fE46��G�u˗�@�ש`c����˶8�VK���d���B�@�m�+�q�]�^����y!��L�<Ԯ�}��F���X_Y��D�z�|��.;t�ke�s|�Ƕ��Y{�0U������4�B/O��47>�F(ue�6Ϯ1Ǥ��f�ט�x�_w��5F}�XP[d��r�j�.v	�w'[�g&\��?�+v,��4����p(G+vpU�u�ʗi����}]�[�l��h`[#pc'
�@T�>P�u���4񞕤+�מK �w��1� �2��mc+�u�ik���̸	�뻖f�ma�z��}���&��w7�v�3�A[	_{�άuc�Y�,ؒ�
�х�%=��v�XD�u�E��-�{�&W���\�ŷaJ�Z:��)�L�����{�o��&oE�h�Q���j|�w�������r�s���'u^V�T{�3�ox��Q>����$��>ŀ<�]zSf�ީVy�#��E�d�����Z�ڕKwz+z��~��[�EןL�Lڠ@�]Uӯoz���c����\8�wO�>Jiy�G:����."�_Lڪؔ��G�������5�~��f���e�.��ܿt�����97|���$w��y�=���󩦇5���0�ʜ�&��^�̖�G��~{�f.�c�^�`�\�r�<4L�o=��32c�v���m\�d��������֯�T=���޿O�ƻ=g�؝���:����ҟ�m�-l1H��F���W����6B��Π`�Zt���q�h-aw����U���k%��.�]���\�s/+H}C��]�#�r�|�e�U�#������viYeV�s�����U�r��P�R�W�J�Ye�vb��g!;YZ�J�gvq�J��(��O{���{X�@nl^�y��$_��,�>h�y�C��?O��/b}�}�i����q{<㥑��y�y����S��;@ܹ������|d�
;\.�{\�� \X�?15Ǿ�OM�Psݮ����mǝ�ys��/:6����Qh�.�7H=q \邜�cxYb��*���d\��o>ܝ���m�֮v�X�'b�X���%p����f��M�+iz�y��:O5��u���F�:й|���;���!��<���m�I��;�b��̮�ק�_��]PAՎs�F��͈4]����s���d8װ3�{ӣS��E�.4�T�tި=^c6`W���=Y6d��hc�WX]�]%��5���u��9 �97�n�w����e���"�ڳ��ml/���3��8o3=�K�s��̕�BŹ������Ck��%�i.X�)�5��(�f��%�o�����w�~�LE<R��*���G�ƻe_K��Gg����� =J��`�s���weƬ�RŬ���K��E�D��i�2+{H��b!��!�'3����i��E���l{�ײ�݊��/zb��3tǏG%��Q&F�*9��w0ZiV�/{�.���v�Bnj�eƪ�z���ٸ�(��)+۝�������t�s�,n�|��W4��:_�[]��,����2����t�t�?,����s^i@�Bꛎ����eF6꭯?�	�*_��ڥ1Ρ�ճ�<��o���[�1u���=�����pV㎗�L{Y��V�	�D��p����z_&|s�۟�z�).�'���D#���\c�rwP����їy+�羙��"�ԯ=fb��y��:�OޣX�/����1�x�-T㧖�u����7�镗�V�>��~��^���S��������&�Ǖ��>�ܮ��?^�9���p.f�2s�u&�~��7C��O;��x��jx$<�K�)�z��j��͋�4I⭞\��7��U�v�u�<���Ӡ�p���//,�2:˘����ı�<Btr��uz�f��n��<f�3�s�l;��9t�le���3Y�B�����}|L��px;ضn��/�4��H�빖�*ޗ�`�VT�[�l�å�i��ͫ�/��ۤړ�6�̚�I8��.M�m��&7��F-��ZZ/�݄�(�*=�q�؁�������3�z�8��-zv����߽|���T�GX_'7�I�y[�Jn3�V��/H�y�7�wٴyN���Mw~K��D���J�ϐ!�x����盤c]t.W����͚�㽯 �ո�]x&Oz�S��9�2�����S��A�o{%�����[ͼ���/di������z��c�٥���^�M-�y��}= kvUhnG���оr��~��6��L~�{�aSr�O3pWC�-�Y��ݱ>�U~pU��	��R���b[�[�O%'/?i��2�-�W3��Mg�|ꏧ���_����ݎ�ߵ��t9ݫ��7k*��/�+6R����N�Y��[Ɍ�%f�����EVOP7.>� �>�*�u,m�wPQT|�V�0
�	�w.a:��j��S[���{�����Z���<� �5�j���k�,��,���8�;�N^�i��.š�	/m�|�=8�l�S���\�[�R��lbO�oRȨ��54��I���CKR��v8��Y�tt_��z/��u�~�t�:g��N۷��T�����S�zk�����M�a{tr��Po�}���>��3��O!8'�r�����t~q����u3䅺�r�ͩ�
7��z����W}>�4y�}WԘZ��095D3���]�,����7�.:%羳s�M�z�/&�>nN��:e�@}�.U�Bm�͓��}h'7�_��X���F{W-{�)����lB\�zKp.й���?:.7ɯ%����*�wCz��Z�!;��*="�R���b����g�ؒnm��x�d��g%��v�ީVy�S��0WU�CV��a�z8u��Ey��k�73��]y�Ȑ��]u=��^�H�ݞ����p^̐���`v��n>{�IOD%�v�rUېmܶ���X*h�k��tT�2l�õ�O�Mi=[ b^�h���o�[젥1Ĩlk���0�{,]�9�a��e�h�43"�JA����=SuҁMC��Q�,ͧN�d�K[�]sGО�U��s�}��5iT���:��{� 佫}y���ST���BI��Cn�hf	��v��>�|s�V�|��{>/��W�,�{�L�Jk��eGN�ٵzFZ�I�yG�|�ۣ�5Š�]��X:�Ut���[Dn�qJ��Y�<̚�cjr���J���Rc��zǗ�����Dfy���BM=Ւ~���9[gݳ�ڸc�D�Զ�w����;�$�zR(> �+K�ܱ%W�`�����ߦ'`)��_�A��"�/g�q���m����|m�;
�-a�K��o����չ��${�as��[���Yz�Ř�=ɮ=�'�F�7H&��M�Ox��R��W���3��^��n�\�:AꭩV�k��v2�m�{�e�����W�4��	؀�:Ǔ���H/��t���jR���������ob���ìhut:?U��r׫�op]&�|�߲;�^�
�3�J�w��PI�Q�ځ!�,����'kl7)@�x�T.=��]}�-7��S�~k�Ғ�	\�mw"B:ܺ��I��ڗ�9���l��ئ��tɡ��༒k=�.�ѭb�y8�gFP��Y�6vc�_^��G1n�_�C%�����c�m����F��G���n��m���|�W5Db}hgNt�߰ٸ)���B��L٬-i�4*@��Nt:�-dZ�mI9��KM 3��;�9�6����d����m>��XkQQ^�1�i��0�8���weH���ϧ�W.�%v�r��V
���eF9���P� k#f����^�"�D�϶�|�����
쮻�(v�(�� �����,�h]s���vҶ�9�9�����������X]�٫�¨����f�n�#:�C���s
R��a�����u��g&�n�O�YG_�}����-���y�����B��\+"<ZT.j��l���귆S�E�-������u�R�ջ�8�����NM�f��,���w�eډ:�R�E]Ntڸ0'�
�wv��Y�T�ŵۖ��p�w��[n��oj4�e�a��L⤛[Gt�g��ʺ	�Ro!ڍ�5�IiK�����чVt1�����e�./��w�yeޜ.�ki@�U���O��s:,Pc�͹QX]���7��[֫a������:ˣx�7���L��ۡ�6�uNeY��9�A�X�Ke�eΝz+�56 ���Ӗ�V�¯'�C�VL����w��.��A����[�����4u�ދM]_9�κbӝO���"�fq��6�Pf�H�������=[�Gt�+�MiReC��4�
5YS�%u:���5xh�v5)լ /B�0�c�+d4��֩�v�4x4�c�d����G�N�o���D�DWv���*L��еR΄��tX�'�Q��H:5p�9P6U���ե�������B�{T2�d�7)򣝶��L�m�;�.`��Ӡz�M�+�@�Xf]�L�\��}F�G+Kp�<k�]�'���˫���L�vk�����|
��ax�Lآ�a^��+�s��(�0m�|*��1���wZp�k�hOT�&4��Wn;2dprN�QX��f�- *����d��q����}�¨�榫M�|�nť�{3[�*���3@_1Ւ�{d�˟u���Zv������wVr�7�c��Wa�ޔ�� �}�c�U+���e�tz���k���C's�{�C��L��\�CT��w�l9a����bX�Ò�#���w�.5�&p
�Х{�$̎�A��rs�,�w���%��w�^��2�s/2�`�v[��	MJŜX�`��mV�'�1s����|r�왓�Γ\I%Y�W+�����RTET�J�#J����H(�`[d��,��CHT�0E*Jʒ���*0�PF�`��ejܰ0YUDX�U��̈���[-�J��mV�Vc���R�«aX������ʃs.Ć8-�R���%h���rʋ��-,Z�TY�PX*�r�1T#m�1�	D�-TW)Q����"�J��[j�Uq�R�9l�q�U2�d�Kjխڂ�*��l���U��2��bƖ�B�%TfSPZ��,`�
��1T�#" �(�,BUˉ��±TŴX,X
�"(���,"�)3
���R,X
A`�Lb2��a+\j��B(1-�
*��!���e�1�X���&&&%J���!�QHU.��1��Sr�F�i]r3�遑\V%V5(Z=K�[a�v��e�B���\�����_=j�M��t�Įz��c�����<�p���;;��|�b��<ϺSR�k��AV9��3�hg��5ֵ���~�w��2O`g�����{<�S*X�FE��w�PN���ܨ�7G-U�*sDk����鮒�3����u���3��gJƱ+Z5,go:l,�r�¶2����ah?:��x%�v3����ٴ+ڒ�5��{�O-� ��Q�]V\�B��n�����S��a�۝�W=g�ِ����AɨL��U��{,q�^���LU�\(�qjF[�ށ�E�۵W�r�%=t����+�2�Y��eQ�Xe���޴��-��(�k�-���c�ۭ��R��k/6�23B���x�:�u��r�
.|w"����~��ϟl_k��c��O���QN�ΖL�5��y2^�T9�N�oj���/r(��8�޽s��U��z�2�&�X��������є{�ؓ�o��E�����*%�G��ׅ����] �Gqf�]XE���i<�ӴEk��*���	�6�8�G:�Aݰ�W��d��j�c���ۅ���~�6�����7���ٚ�����Gk���>��]]�[����'��6�kkޫ��T�^Q��l.��2���� pzkE�C%z���H���Ѯ���W�\��2�8�����s�m�{D�ދ��L����~X�>�cK�'dE��8��[��gc����>��N�uGσ�WJ�T�رբJ���T�cܣ�����u���n��ή�G���vM�#�ǵ7����r�KI���~��e�CjP��Sjկ���y*��ڟi����0H��]c���+I炊��AՄ��w�o�)��=���@"��,Z9w���H{fwrO���R�|�-��?>ٹʽ�r�%�o�yFH~��ods��}i��ŭ�"��2$&�k���Y{f���,ay��"�O���f!�*��s�0KQ�6�$�М���%�U��_^�vz�'E�TU�G���b.��A`u^b��n��̒|x��h��6��Z]�����ݹR���|���-y^]��Nh�/}pBoJuR���"�H�8���]�qj�f��V��.�i�_U�)��-��孩�����4ޠ}u�>�k�����ˌ�ݷ��������kvUo����m�Bpz�V�鋳մi����{�wgƙχx��I{3q�$�e% ����u z�yE�^/>�'�^�W�T��O�g�������S鵮
Z���ۛ׷�9��I����c3ݢRco}�xy�,�E�C��Q�-�Ǹ��"����\g�t�Ou�ymw��_�+~�n�_��Q���v�RJww�r/O����y���|�bk���ϻ����X�y����5��ywT��^�QAp6=��+��ӱ�{�U;q<T��vfa��As���ń�����8�u�?8�s�
r{�������.����(�S���ۯV�q��WZ�� ���}6���a��꼗�-��X��$����`kx|�-�k�Z�Y��ݠNܖ�ls�s���L�[�	Ź��	:C�	�6�\�M����}��(�X�:;Đ�v��wѕc.��g�F.=�Z���{���Z�y_@S�g���ͺ�j���^�)�4�7	K<�@�|0#�Mb�yۜ�ryy�і�`MRӧ�[�;�;G�?�U}��H�r-+k��ذ<�̐>QV�w@�S�\����ٜ�z@�՞����j2׾`ȕ{�@Os��p�ɪ~��R�Ͻ�S��v�˜ҙ;����n�ު�'d/;����3��]y2$&5_h���5tf}&�G[��Ī-;+�9�嵱>q��x!���.�U�󃐹7]7+�*dɫ�̪ٞ �Y},���Ώi�~�B*�#�m�i�ܧ��1��^[Q::�em�:��4m����l�����q����;I�'zo��t}����_��|E�{�\�l�6�8o?h�����$����~d��XT>d�+}HT�2w���$�O��+�$��'|�?I�8�4��0���C�<�=_�}�J5���G�'����_Ooo
�7����8��|�f�ϘM��k|è,����Y8�����x��6ʇyHT�2o�{�I�M�d��sG�	��'SS,:�x���'�7�����o��}�z0���a�i��8��o m4���}����5�a��5�0�'�;�IĞ���w m�l���6�uS�3�u��_}(U��~LڰC�{�6�����q���X|�q:�yCI>Bk�m��:���6�Y:���xI�CGy���I�<=�d�T'��@�&����2��d~7������O��{�ƾG�������)���:���;Vsu�X��zsC�gڠ�^�'5�F��f��_&V���.��ur1R�h�m����t"�Z�!������vڠ�v�V��b8��� ��o���\��^鶌�\�o9>Uzy��W���T����<�w�z�=`^�zԟ�6���:��=�:�=J�!ԝB~��c'Y7��8�Ԭ��x�:���N��'����q�	����<���[��y��?2}�N�y'Y'���IY4��}I�R~I�T'���Or�0�0��T8��2~ف�N��k�p�'q��ϧXJ~���������o�{x�z�w}�3���<`�OY8��v{�>a=~d��O�N;3Y%a�C��=ed�!����N&���6�SG�Aa>������_���ܤ��]_�����w���*Oq�:{����a��0��I��:�猜d��9$���]�I��њ�*M�=ed��[hu���ԍ!��h��|��W?=r�g�9�~׽���$��`q����d��{߲B�u�|���u�I>;܁�Ğ2o���6����z����T�H'�@��@U|W�_��m���3�U���?2|�d�$�tՇ�$����}d<�`x��N�C�XI>癷�O4���^$�&�9�$�i�S�d���>���ؗ��N�㧯��W�U(N�ΡY6���hIĜeO�u=5a��N3�>d�C������}�'Y6�k�μd��f���4���o~�{��<�;���y����I6�d����u~��(M�IY:���|��>g�XN2m?Mo!�N3��q�~d��N2O_����d������~�*�25����-�l����P���u��i��,���xɹ�0I�?�IR���q�d�+'��Y>�La8ɴ�y���I�N!�7��M0���9�������X�_�}+��ۇ�8�9�ˇ�N$�{aP�OPY�w$:��5�0��:���T�'��VO�4e���d��k�����;�-佗~J��:�GI�}�;��^�%{%�PG�"���赵�����W���`�k	8�*��h�W�lD��F�+igP�ˬG`��
�>�mC�$Vrwʿ�5��s��|�J�T�WY��S��#q"� sBz�$��.�1�lT����_� ��[ϒy�ￓn�>d�wd䟘�:�*V����	���&�q!��!P�&�Y�i'�=��O�'k�2K��X8�����z��O'u>�������~�d����t�ì�d?k̞>�xé=��d��N�����IR��{�:��+�9̝I������N2m+��'�?�'�����#�s���_�~o��?�k}���x�a��N'rÌ���זd�!�^a�u�Ĝa�ߙl�'�s�$�a��a�IS��ì�J�k���6��7��;�g�~;�k�����׺΁�2t�^��m�A�%|I�N'�XORi�2�M����8�z���:��=��O��'P|?o�'�u�����'�o���o��~��wZ��9���7��O�Y����2m�ONs |��&����OX������'��z��=���ԩ�Va���2�q�l�C��Aý���{����޷[ιF��A��'$d�J�nGȓ����d�'��]�a=t�$�� ~��~a�5�C�~d�k,�$�*~ՇROs��9���w����}�u���P�'�(�¤�&ҳ����I�/)�~a:�w�:������:�o=��$�$��k$��`~>�����q��!�?2q9�s�9��ϻ}�����v�O�xΟ�u$��1C��J����%a�N%f���C�w�;��u���d��O�=��O_�jsY'N3Fk$�6�{����~��5}�������������q+'䞳�Hm̛Me1$�f��O̓�F}��'�5��+�u�;����C��2wv�&��o̞2sm�u�G'w�߲�;����������9�O��~�+Y֜aR|���i��N�����MO�>g��Y�C����y��񓌝}C���U|��`���}}ڤȍ�_�Ds��HG�zd�ʹf��&���{o�)�7C��QY}4f0@��I:Ct/5����k����y}�͗�WZ�6�=��yK0u`����ϝ<A�pf�Ƨ�Ț��Md�&Ƙ����q�)�S�טN>|��W�W��V�u����{�g��<tɶO=��g�O�<�VI��s�IPP�nϐ�8���l�$�'SS$�'��|��'~��'_��8����z����k�?yߵ�}�w���'N��q���M$�d�N�x�Oua>g�M�̋$��k$�(L7g�VN�d���q�����q�F��}�޿�V���zJ�#��N�\�W������>d�?!̧�OM�Zq��P:�I��'�?>|��CL�;��q��IR��x��|���|?W�:U=�/�������s����$�'��}�}��4�.�4�����Iרy��i'Y'<��~d��<�p+�6����d�,'R{�a++	�z�7�;���y����~�]�%d�X2�l�d��5��q����i����C����&�k{��%eC�w�:ì���~d�
C��P�OPY�w¨}��������#�����֯���ROw�0������'?I������Y8�~�>2i��ovӬ�a�ޤ����'X�J���:��
���Of�3~���r��4��t|�$�~9�?0� }�%ՒsvE��I:��2OS^P�'yOY�M0�O����N��w�'�T���+Q���&�_���t[��@W�_���'R�4w�<I�M�a�w�B������I�O~�$�XN3�&�Y?'�,8�<z�!�'Ou���:É7��Z�����~�y������?0�'�/o	<Cl4s�u���=�N��+!���Ĝd���w ���O�v�:ɿi=k&�:�	��'��2�2OYS{�߿w��{��=�}����}�a�0�߸q4��O?{�m$���x�:�S9�SL��}�:����'}Ì�d۴��@����%d�����ֲ~d�o��_���t�� ]b�?��"���U�i��6����_��_R� G��6�إ�+�+E0oq!���o,l����-���	\�gtX����}��ծ��;+�ӗJ������qP� ����q�@�}!�;,Z�VXw�A��}�?wg���� �����;n��$���>O�P�I�T�jìY&O�08��M{�m2u*y�y	�a��é��<�d�'=���d�'�̼��_�|�~�ɻ�U��Vi,����ŉ���l��6����P��!�~d��2�0�!S�����P�'R�=>�!Rq��S\�!8ì/)��I�We~������������M���Λ�s�o8�IǬ���N2M��a*M��d���`|�q�q�m�5�è,'��}��N2�5��*N�w�T�L���߯�.u�ߕ�oVg�N�3�|��4÷x�Y>I�w�$��'XVI�{9�$�6��[R�q��i�Ԝf��	�N&��O̓�F}��>��z�u�������>�Qi��̟2q���d*�vw���'Y4���0�2x�ýń�|ɩ�a*I�~'?d��	���VN �RC��O~�~��_	_~����N��~_g���~z�k�Z��i��:g��s�!�w0<d�'Ϩ{ϰ�'Mw�>x��M2x�	�u��O;�B|�d�<�V�~9�$�@}|C�}����m����ٞ~-{�f�o�{���ƠN�d���?k�q�q4s!�N��x�8�<~a�?a�OXMs�:�'�>@��'S�&�~O���a����q����o�9�No�Ϝ�߳���	���J�l�?I���'?SN2m��o�2N'���'P���8�u�;�0�$������6���:��6�������s�k��}���}���	�8��PXO�o���I:�IR|���)8ɶN��O��O�o'��:����/4���'�%N�����N��}���y�O3=��^�~����7��O�R=�!P�&�Y��`N��MN���I�9�IR��YO��*N2m������q����;I�'{����O}9]e�������^�o��<��T��$р�3���*(�.״��ՍI����j��t����|�[�@���XZ���o�{��u�@u�M]����
�Y8]��{d���	�[a���K�� ��M����N�Xk����W�z�o�_� � 9�q����U���O��?yOq����������B��M�a���'���5��I���+�$淒,����2�&�S�2q��Z�n�3��g
��t؟�/��:���$�'N}�6�d�}�a>aP�)�ISg�ì�A`jw�$�M���y�*OY?���N�k�2J��9��Bx����~��s�w����߽�ｇ�'��P����^a�4��I�v����/��	=C�h�0�	���u��P�;�Oq&�P�9܁�M�hߙ����uTz�׮���,�O��o��˓L�N�a<~d�h2Ì'��x��Bzk�6�2q���ܓhu��/����!�4w�:�d���y�Y8�	�?g���_�t��+O���?7t�m/�;���盿�L�d�WĘ��Ğ5&2q:d6ϙ4��:�=J�!ԝBzk�P���MO��6�:��~��N���N��'��{��L�>�m�4o�?|f���5�ϸsY��M�~x�{�>d�'��t�rN�O]���i���������e	�~d�h2�0�0��T8��3���u�G��*N$�*=�G�~��������{�y�B~I��{�$���y�Y:��y�p�����?Y>I8�5�Vd?��+'Xq
�z����)��hu5��XO�<�u��W����~��������Y>J���T�$��5�rB�u��ï�'Xyy��>x��O{�O_�5�d�a>ML�IRm!������R,��N'��y�_9��^~��{�|��}�k5���~C�����$��s��J����x��N~�
�������u�I<;܁�Ğ2xo�Bq�2k��VI��Y*M�>�6}o5�i��϶t��g�VO�,:[�6ɴ���6������$�џ`u������8��hzw��I�s���'��d�`x�����_}�P}�[�w������5n�Qv<H�vڗ���OsM]^f�Vʦ#犛���_W''��}�&��[@���h�w�]1��Ng�i��n�M�UU�ذ������E�ࣹ�ov�G��Xw�չMM;B�ȃ�q���ip��>����0�hC��@p�5��/�@ z����.���� �#�T���3�>B�|���h$�O��
I�N��X}l���k��:���	�>�:��	��μd����=]�߁���/|;8��_A�}��c�^u4ɠ�$��IPP�x��u+&̠|��>f�,'6����\I8�s܇W�N��ì�o������<޻�~.�����'O;��l�I�9�'Y�O��ú��C�M|�Y'��IR��n�aY>J��I��}���a8ɴ�y���I�N!��������1��uw�f~��W_K��9�����0�{��:�9�n�8�hw�
��M��S����M�̓�4s̒�I0��
�����q�l��K������f��y�s�u���d=Bw��4��N��{�Ԛa��:�*V�s��	�����N �;�
�=Agݤ�$�5��IĚ��d��$���><�{�����?oz������t�&? w,���z��:�k�4�ɦI����i��x}�d�+����J��2u'R�I�OR���a
�ԛ�x2��n�������ھ�c	�N��I_N�7dXx���ja�I��x��'ڧ��M$�u`z�̜b��	6�Xh�0�$���u��YǾ{����ny��}������Cl?2|��f��ml�7���|��M�u7��Ԛf�P�	�u4Xi�M}M��N��O����4��'��$��ߜ�\�3]>��y�����6�6�w�2u+!�����m�O{́�'̚�������i=k'�N&��m�M3A�q�z�?jì8�>_c�T>�P�WT�\lή�o>����>A�����O���Y�$���d��'��d�'��]�a=tw̒�x���O������!�?2u52�2OR�B����m�u���˯G��X��ec)ʖ�^n��0�A� �v�$�g��:\[FU������n81��:D�^sB�XYXlZ�gkL��us�d��ލ�=Ͳ�>P�xb�D���r�MN�[,��yo�p�3���(�mց|ۣy;a�8�F'/`�]�U�l�<���'���:2N�ܯ܊�}��Uuv�'�u����D�a�t�ɄRk�V�[�{�n�>đ�AHn�q��r�pLŜގ�8�λދ�Q�w��,z��Šp�VԔCLjkE|��GK�E1�;��֗l�w�j�y��a�D+���9fkZ��cB�R�kWǡ�&�����a5���5(WA����[��m�U�ݘ �r_<��(u�!;�l�S�](���CT��9���M��;b�+���ձ�e?�@EV$��_Ի>��ٗ$�6Y�Uo���]$�Sn�m�ɑMr�=�2ļFu���FȾ�E]��AWYU;m{C��g,v1�7#��P���[��Lw�-C!�&v�/�óL�R�\��y�fԫ@Ǐa��S��W=����N��l|��t���Q�VG.��K�c,��t������<
ɛ`Fc!�H�׳I�|�Z�7e9LvS5���T���M�K�a��ݒbɳ��V���M�b��U���n}�ht :��RX�]m�%�0��g�����я{X���v9`̝�w���,��6�o��/��u�$<O����
�LVt����1/N�/	�O@2hT��[PSʛ̫T_sy}d͎>v��K��M��	�SJ(u��+����0��x�y������	�b����!�O31��:����I���;��eggf>u�f��F�Q�q�T�(�X;^R6xÃ�^Ɖ�j4�r�z�rǫ/w���Hx�@�6KEh첦M�{���-�(c�0,�+!�w����:^xM5�Wʸ{m�!�<�5�;X̠N[�l�u(�|f�BRa����Q�#9�`v�ƹ��꽧x��t�`B��,������wu�-��r3�%q1����Int ���GY�I�fK7D!ܬ[������ _2Y���qH
�r��yG��Z��"w��.\��*Փܧcew+W �ͅ��֖b�*tI`a�F�u̔���ݻ�ę���\�1£���W�ӳ�5���+_]D��4z'b�~Χ�y�8�Q@ά^5��ڕ5�]ظ����]�M�)qGm3��4
[O���������cu}`H:m-��շV�/0��n|�*u�(��ۑ��{�/�igg�y��n��]gj�v$]\��J7q�.�M�\yҰ�-������F���mkZm��.շ���p|�tyS\Y���e������9fQb��q�=����Dn^�ٷ�X{x�Nt�n�;Y+��:5V۾����v�B@�p�:M۵.��C�T�8j�{IY\��T��z׃��g��`���|��J!m�-amҋ+��A���lĕ�V��kRT1�V��TPƲ�*\�U��0%IY���m���H�*�Em �kQ��82
Z+aP�G3!�H��R�PQS.2� ��T�Lk�b�Ƃ����P��(b(��2�EIZ�e�	m	��[V`³-�(bC-����@�)��K��LB.3�T-
bK��r��(6��QeLqШ9am�H�T�%�Q�2\�E�*��r��D�Q�aXT
 �5�UDB��b�(B�mR�[H�cZ�9E"��`��R)�a�C2�`�e����F���X��L�QE˘\�e&26�\�PQ�G3T��S)�����"����&��Φv$�f���o.}hv%��\����K���;2����_���x#����}�4u�fװ4��[� D{�s;�wm��'�)'���m��r':��9�	ĝB�g����O�Nw�����OMy�q�z�f�J���R�_�m�޿�9A��;��3ӽ=o}���̛N̸�<C���C�)&��2q+_{��8�Ĭ�=��w�w�$����q�'̞��O_�}�/�|>�����9v����f��_u{�~�앇�C���VO�u��Ch~d�5�ēhq�?P�~d�:ϲd�V���Vd��w���~��'wa?2h�0�2x�ϳ����{~��{����y��O�$��VI���쒰�!���'X~-!�:���SO�q5?P���O�g��s�!�CL�d��ݐ�O3C�����y�{�|�����vɕ��_����'��f��?���s\_��4�y���W��:n1z�Ȟw�%�u�'9�ɒb����T�J��>_�r�@iL�o�w�5�<�K�gG�~�<�K^�f-Ϥ��&D��������<ѓV�j�x�_)V��ܾ�U������r�������BMB`��fש���X�RF0ɔ}�P-��r^�mm�N����Ub9m��znOw�;��{M��ڥ��՞��R����{�ˎ�ٛ�~ILJ ����< �G�)է�ت����J�κ�f�E��im�n��vF)a�c��2-ڌ�m��� ��t�Y���(����r�nn�-�Z̇��[��˾�Y/�7��E�;����tA�/.�[��ha��[踫����T�����	 �JKg����z�fW�_�������X֏d�[��y��͘��A<�r)07������ڙ�*����G^�/D;+����/�>�&�s��{=�(Zy�l��E��ع�0^���!=�w�w/�~Jߧ�"��i�X~�@���z<Ǝ�Q��jc/� �z�9kÜt��sv߷^�&�o�:�D�r�^�[��z��yQ���o8_8��{�8���a^�V���k�]�ϑw��wp+N�Fu_ɋ��xw��_?8�s�^�~;4ǐ���z;=��{�\VدTh�`t߮R��l>`���ؗ��4�n����](>K)��X������t`.Wvn�zԛ����u��e���&d�I����9f|�jX��أ\�����ҫ]��lN^��OeV��$�<�Q��x��.��<�;��a<�@�ɧ;�ϥy��K1��'�ٿb��\8-^E�a���#����7�j�uX��U�S��@]�>�v����Y�E��&�lL-Ȏ}��6�w%5�<@��ou7�Bj���Y�T�G�7���� >� ��O$�U�������x��77/;� �L�|�]x&E��ٞǱ�}'*�^I��t�xQ�� ����΅���F�f�6V窄�AI�s��xn�K)�j�լZ�+���^vr]J���ߤ��R3<�����̞7�оrj�q�R���e������(��B!s�J�ֳDt��?t�Uc�2���%=�zڶ�ecZ&X-`O�P�\��{#����={v�\}өpU�q�$ǵ�֯l6{�w6��#~+ɧ�Y5��;�b�<���L>�����:B{�w���8�NӾ�$�5v�z�BC@� _����`�{��y��:�M��"�I���e�OG����o��߼XZ�W;/�jK\-���N���k�-&�����&������}9��^�E��Qz� _U����H)�㧡/xz�*uоJm���2j���S�}.=����#"I���2��z��2�\�}.���ݷ�z��0�@W+����Э�npz+p��lܛ���bp����� ��������P��1����.S�5��:��eG��՘L�j5�Z���HҞc�}:�E��qJrb��V}W�Ŏ��1������$6����ko3������/�Ӕ��\s�S�ߧW�}�
���1�z<�������u��r -�G���$�������K��%���˴����r�\��U���F��+J�X�V�{*�G���q���/�́nLJ�r���خA�Х7�;�S����s��ծ�GvOmM��v���.�k]xrA�n�!��Y�ȇ�az��-Y	˾����zG�X�8�{pqkpI)�0;Uu�`�־������nR������z{%oR�LE&G��쒯Brj.'�Z둩�"����>�1��r�פ<^���[��[��IO�Jͯ��܀c+�����I6��� ��e��j��?wr��t���7�&=���A|����3yQ��=훗����#o���7�u|���kj6�څl��ن�:�m^���٣�=��y�5תՒ�T�l2��s��l�ы+xKS�Ĭ�P�/7�Z�)�ic�/�*p�垷����w�v܊�yK�慩�諭���4�/���5�ۀ�fϵ�^߇�9ʾҼ_��0>ص�Ut��n�Tើ���ɒe�#�I���l� ����{fܜ���݅`�^�$�����gjǜ���=׵�|گt�P����m������R�n���9暷��/wp�^��.,��ܚ��)�S+,gU��vEa�zT��k��Kت(���IH=p9s�
=��N��}G�S�&�n" FA��ѩ4�������~����p~�G:`��x��w�Z�B3��	��&�S������G�"u����t�{RzmN&���y&oZ�w���Zݝ�,к|�:�v:��IO֭z��r��5�[�/{̕�>6�_k25�� ��E���8�V�w@��b��q�p�f_@�,e��~l�RW��W�r��,�d���h7�T��*���\�ieg�E)�:BI�݈�� '.��{-�ƥ��Fn?7��U++5̯P%�������Awλ�SZ�,��!�7ӻ;o�4���V����riT��樲�B�,q��o!ܽ�Fli�V�R�����x�N�;���>���w�~��^�,�{����g��<�Z�c1n	"�\A��oAxn^������*�|{��}���_w��;y̖��m�	*�''8�Kݔ(P�zy�[3�����^�!j���7eU�#�m��w��p��
m�V�-�yժ����qx	�uL�̣U���IG���Ԟ���!O]oMg]��g�BJ{K����I����y����%[ŵ�V�����}�p�s�/c�Rc�ݽ����Գ}�C��N^;�4����jt��I�g��}�-�}{���qҞǻ��w-��fW����gQ�iKRy^�*U�:�]��;�.,ϛ����v�=�*��u��+����R\X�|M��ۡ�J7�yo83��=E�<
=OD��3:Z��>�Md̏ի���/;h,�3��	�/C�ަ��E�ଌtgf������8le�jt�����J��*��5X��[�!u�Fy�ѩ�h�S�x%q��i*�d��^]�`�e8P
���uu+�k��':�k�9���czP��z��L',.G���J��u���e�l�ي$�e���> }���䚮H�����+v{�j䟏�V��⭁��Kɱ�ݴ�ё�cՊ>�z�C_J���U�gτ^�xs#��htzJ۷������\�����e.ځ�9��uKf�Y3{2@��<:�أ�:���&-�zl�r�^Z��'}\�k8��}���1d�I�sյ�;�xI��2����B���t:yo�77!y��y�x)^��ևT�y�m�Z�y�ܩk��EEe�l-w��8��j0�����	�O�sl+j�}���)�o��T��9�0��_o����5O��������B��n��Ds�NŎ���7��
Jz�Tˈ�S�,/}j�Es]��Rz]�!=��=�~O�lI<Ġ�3��} {K����ʓ�&T�e��ڄR�5�SE�7�������]�RQr�c����G^�/H�V;ݧKn?#���P�%�]�W�$�J�+Q�ݹ�rW0o�[c�6`?�U����%�Q.Aݺ>�z`�np?�i�@�v#I%k���.�q�Ȑ��J����-�".�\e�obO&�?��Y�m��*l{/������ۭ�?Q$�oqR�銛���'�;T.�j�s�[���<����>�ǵXs�Û?\��u��x�w��z���G/o�{+{S�d{����^n�����JN��2,�QS�[���Ņ�^v�����'�Z��׻_e��s�.~�;R����?15Ǿ
O U+�m\����JUk��@yw:j��{Z�Uo��8Q&�Ũ�b���D~���^���׻���Ee_K��m�{RR��qΘ)�nuf�O���ӎU4��} ��
_��;���a[E6=O�Nߢ���}'<��gK�g���,�.Ŷ�aJ�tUc��Ɠ�+^*=ϙ�7bWO9g��iTZ��n,���MT����Tؐ*CA��":Z�vt�s9�hH;ӳGMO���z�.s5��'^L����u*�<������S��)z����`��e��nWP:j^���<t V�R�d�`ԗ2q"�SǓl��v���ܨ���Fj8�J��/^���������;/{���f��a�]X�-��!����G+w�����ae�&m�{1�)�������^����9��K^����$��E<�������ξ3}�x��b��w-q->�`��΢�#��Ϥ�М���q��ʸ�(��4�|�k�=�{cS�����Ǻ�KvU_��P&����A���B/�F��&�ӐfVE�����b�z;�L��UX󂭸�̲�uһ�3�xn3$��*k�iY�Rܛ�6{~tW���o�G{+J���ޣ���ގL5��ނy��
������G��ձ��h�9�h�ly��#�.�(��3�+�G}����uSrwmTi/vf�̕C��Y��Rn�v2K�],�o����9��_�p1z�����pMqo�6L���m��ݩKy�'���>��]�J������_w��A눸�
��~�{��7��u,V͍���n�C��:f�����D�2����塰�H�9�8�ݗ����[�C/۱��X�z��=�oJX7��9z��u����Ѣ�e3#��*b�oa���v�������M��6Zn.N�n�LۡW�%��!���I(c����Ȟ.zC]qK�b���QN�MƓ]�$��p�0�i�Bs+a��`W��|> l�6Gճ��ytEV�S� ��	֮_/�7H=�=�jA>ĞQ~�[�
���땜�N��ï�c��H�����AG��Dz��[K���se����}5ы��S��_L��t6_Q��߅N��8"Y�9�su�N/�����9�{?~�;��Nx�d��g$�7t5z⬏��Ҵm�����_
�>
B��϶z\��k��_�H��dJ`|oi$�G,���o������v�ٰ������d�Cos�*����r���8쇺y�Nꗀ<���^�l��zN����9���Z*��y�x�n���,���[V��N�L�^��ZJ<��>�q�#�#���??E������Xތ/����Xj�*O�=�[��g��7����(=��͑cՖ����{M�5�V8�	1�`�:��ӕ'�/}��s���qT9ݽz
�`i���+���e�_
�4�W!�O���2��3VV��Yk�N�­�|���	E�������M5�-���N��dݲ�U��I"���Xm
�%�K.��L[����#ʝ�`l�p��%��R��dU{L�v���5� �X�M�u�u�p�J Mbջ����:,d�Ϋ�9z�(*Te�vr��4%���@�^v�YE��^��y�r����/jpkP+A��tn��P�ٴ�/k�����ܔ�7�Gr��n�ֺ.=�����(3t0�����rvV�5��X4��Z.�����c�E��VX�ں�5%�����8ރ�¤v�Ll���ٖ�WF��`Ψ7Cӷ%�jƲk�&6����ݾV(�GX��������9;�~�X���m��8��ȳ��t�%�k���eS���8f=��&�+M�[K{�'/�n�Ix�af$�ÎDe-��6�"�5ZI�����T5vU�vdu�n��B�:�>�|�:L�׫��Q�m:)�q�q�텼��8ʂ�㡑�4»�'B]5�5�;2���tn�о�Vc��\���ʧY�A�.1���x�;d��N��;Z1�v�2�ݤ�7U��:���N(-��0ӭ���s�y��sz&�K2���V��\�΀�{��U��>�u����g5Hzm�O�0�]s*`ڵs��I9%+Er�L���v�v�U�\C�E��O��,.�\D˖�w�j�������
Af�-��SV.�U��y�ɩ��_u�7�����Q4��+ulS�3������*-$.��mnf!�6�s��"��>�����:yW��B�[��x+��qg>;8�DWo$������Q��_G��׵���W�5�Q���/�A��dE�b\B�eeo5:��o��l�����A�X������t�:��]EZX����UgY�X#�\�rz�p�5�>H�t�.Y��,��,�d#y:��\f󖴣=*E_\*wKΏ x�,�����UWm] `���J���A���H���6ˢ�_ �P,H�]l�9�����=���-�"��md3Lķ:�0h�izk@艕*@�f�*��v��5T�n����_K�톅w8�L�5�r�?�e�l�yb����նE`eM���G%��Z�K<(7�vWS�W:N���c5�>�EV+Q�����L���!�|V���.ɽ쇉��4��d��$J��Y�!,�N����"�1���t������m�j�U�^[�bX��3���9�asX�F���t�Xy��gU�f�@ؕ��.��t]/S
��N��4�']u�jv�K\�4F4oB�WfPP=6s��/�w���À̊q��!f̹������\��U`G�Ip,K�*uC7� v
=z��\5�m�2BS��7O����������C�	�U�
&��dYKLLq	X
��1�"�n2��1��11*f%Rc�c�
)2�V�#�X[�J�dm��!���T�W���-hcm��m��J+�VB���c�[2�e�%-Z[QF�Ō�e����ZɖȲ�Z�[�&eU%��J�U�J�7+!��E1+P*()X
#�P�\��QjQ�)�q���m���,Pĥj��Ȋ�ʙ�2�2�J�&Z��(�)KjD�
�h,.R�V�J�ы(��)�+e��bT�lPP����0���S��(�ʋ�"�"��K���R��V�(TɍJ�F��TW1�eTb"�q2ܧԁG�B� /E�u�[MS���	�V��u,u��hĹ����{n�5�x����3m}�٥!�m���R}�n�W~l�{?�}���ޛnG��y���g���p1{�G��q���|�r����A�|I��^�E73G����UMG�V��ژϯ� υ눸�q��G��+���6<��W���A���ZĮ�>j��Ƀ��.��X/\E���}5����	��u��o8�}�||%�B�>�����r�ަ��mp�N������^�d��w��>L鵚��� Um��F�[@����~��uF�=�#��������[��I����䲟�Sí�����b3�oz?Gy�V�����c��D$�S�霳K�;qI�2]�P�k�}j�@+7W���]m��8���B{�,$œ9U��{�|X�Яf4�>�ae�+,Q��ϑ-o���!y�>v��}&v�b���F��ҹ�Gvg�{��ev��\����oo�@w��8� �[���L�b�U�mv���ľ�#5�<'<�V��AX/M�d�~D�u��=����S�̆�n�"yma���x<O1L����8c�B���e�Y��i�\�eN+)Ve5ى����fg������!���CL��V)���>����kd��w��������dS�	檵�V|�j���͌�gn���xgמT��N�����/���aIOB�'O� �J�_��ڰ��1C��}�{���O��=�y6lO�U_�e	
��c6���`�.T�K-rԽ{�E�׭Ȧbjhڦ�ծ
�q�+{�d^��58��i?#g�W1���g�~u0�'}� <㣧��WV#勓��=�%���ߙsQA���=��y�u�9�S��_��Ó�ٜ�B߾rzϻ�J�Ok�i+����C�W��a����Fm��/wxy�{o]�T���ŘG����)<�R�;�ߨ���S��޿,�ī֦�=���@�NRz�.t��9=�ӽ�k�*��ǻ��@�s�8�(��k~���[�Ժ��j�ד���H&���)�ӈj�O�;/z!_]��
F�3�&��Ά׹ JwU��Lqm��3{un���D��ʏDձ氨+
�+P��I�u�m�w9��vXnD3@w���{��M�Q�3�ʜ�@K���m{֍Z�]��$�f$���_S&b<�&��FfIW�r�<��t~�����tn���0�����l@sڹk�6<�$�K��zD������3{5so^�s|��u�A��i�z��r��7D��=�}Mu`[�w{:;��rkR���,q��ʗ.�z����t�����4�ݾ�>�����M՝�����<�)^L�a�]J�}���G�{���}���u���)�9�>����s�"�O/����VnN��Q�/�'	����{2i��z9 ��Rdx!��$�Ѓ�W�e�rS��-�̙�ᇧ���O���.K37��k-�Um�T��$���$$�x���C�S�8�*]����ܟ:���5v����;�%9C�q��;��h���}���n�pLf�+�vV=�K�,N�Y�ۚ��XZY��76���/H�2���uxg������{�x��/�+ts��w��wCK��L��Y+��y^]#�5G��a��z�si>ڻ��R<��P*��g���1�õ���V�*�d�\�}f�Ժ��uҧ�sVU���w��N�\�i�*B\�OtwF�TK+��fo.�G�꯾/4�'�r-�v�sL`����<�=�vsr��������d�[���t���U>S������ř�q�	�=��o�`�;�91�q�7���^ؿ
�~U}Q���88�((�*G9���4���u �;E�=ŉ���7y7ೀ��w[�d���9og>�1��Ԭ-2�V�C �Gg�7>��h����R z�'Y��7I�3�_���63x)0w�S��v�/'�/T��v:�t�sZ�����]�K��~U�O9������؂~�~~��q[��ENAՄ��tV�<_6KK��=�Oek�@�=���x;����(�J-�C�Pm�&��m��o�j�t�������c��G.y���bܒ.�"�h���:��^s��e���6.�jս��Yթ}��d�m�Eo���Y�Җ�Nc+z�=����U�����Jx�6X	 9�g���K�c�������4�WlP=IB�g;�c8{�c��c^>4 �S˚��kk�I �E�=�@���hxQ�������f̡%+%�s���L}W\u^o;���H��vI6�pc'�����o�:w���U��{w��Uu؀/e�d-^�iJ~�w@%�=�$�7S���gVfA�p.a�NXj�*��*~X��,�c��:-�	>=��NH�(7h�������q|;+�셯n]��Q������^'��3���-��m-pU㎔���G^���ec���3���=|�o4���\;�}�Vzۿm���Ⱦ�y��}��8�'2���VnNG1�
��]��Fz�(�v�3�~��.,ϛ��b�}�Ŭ��n�(��݀-�����ޫ��$�X	�z#��V^��y���t<3=�&��m���q�^<"�!o�Gnz�B����;��pk��Ιz��i��'ڢ�qL��ܩ�;������CDa�ONY\6o���[yɽ���W*�S����.d��YOjrV�[��c0E�4\��٭8��E��ةҫr���m<��Q�l�����6̣Q���:MB�'Q�3u�����wV�c��2JD��21���ny�9\>�[�aP����|y���C3xt��S��^c�#5�ЫJ��dqz��O��*�+V�܃�������N�d�^���V?����==N{����f�c��EZ}t��O-�?3��7��/�O1�t61Jmy[�����t��&I�]J�_���s�ߔԭ'+pKv(� ��S^�Ҟ�_V7;/;>ׯ��S'������.�k]y�y�`v�F��zu�-�l/{k� �I���)���F�����@�m�T�����!����k���r4p�v��kY��-ޥr����&8.���U����k�dO��)����'ˠ���+�Kt�sNS��ˡ�qK�e�	3�Yg�	0�Ҙ���}�	4!�׭f�����n)�}]J�1:��,�ìj2�踜���!\|K�f9K_�f�l^w��,�rމ[h���Uxi�*��[�<����'�����Q�k,rI%��&@���Gc���$��^-k�<�}�2�K
dum�+W�J��E���m�,�r�c��ɒ���É�����7�<�2�B)K[���(J�Q���z�-�:3��$j���w�&���Y ����K�����s&f1��v,2�r�:S>�ɕ�i������+�*�PpU�uK�]ӱtn�ڹ����-fE�Ej��jk��W�|yQ������ҫՃ���2���X�]{�+0&:%�2U/:�z�M"�"��-�L�I�����A�,��u3�ja�x
�^�kR�ܹY]x/@�}W}�<�g��N�ˣ����){ޤL�,Z���&x5�s�W�qM>z�� Hu��Kh��Ż��{��F��w�GN�E�~��.�T�tc� >$H
��a�#QPsɗ�Q�5�������g���N�S�:�Zl�tRo�=O~Q*x-�	��bx����l�h�,�|D;�a�u';�G��s��c����x�) N�=OF[E�n)����
ZS^��e��~��o������{�YU�ѿxᨢDP���AV	�x�:h�ĺ�ڶ}B��7ܾ�l"�b�]�+�V����^���C�$�3��3>�� ��`Z�@ ��4mD�X�S�d��}��4��P�>d����Z�!��l-9%�*��(��	��ʘ����6���Y�d�w��(unn����3�z�W�z`~�!��YGF8��]�8�5ގ��"�T��ٮ�wX�:�@�\%��s]k:1שS�q�<qXκ�ٲ�)k���z.�nW`k�;��\o���u��
�Tߋn�P�v���qߴ	�sP�:�0mY8_@���H�f[g;'�Q4�<�-��YNn��A7�u(G��ꪍ�Q�/o�����IY�GY>:)b\.��c�R�4�b�I��ua���/���w�c�f��=u�ć��|V}��.��K�s��k��ǫŵ�{�ea8��n��g��e�G�2yh*<��skƪ-W�V&<s�I��
tWz��O�o��1Gi疕R��CZ��/���X!�zN��@j�%g�[��I^>K��V#K�P�s
{;�嘟{̈k���a���C*Y���&N�@�}l ���xh�&��3G��q{�Z'���kk�؍��r�9������ �z��>�3��S�5ܮѾyKryE�����/���K��߾&�>J��)j�g���^��� 6�m�.Z�8��R�{�2�nxgl��5����;��/]d���
<mg�"��+b�.�5�=����hj�*�w,ӭ��Qj��VO��:��r�\�<B;V%!C��,�׉Dz�:d���/�;��㽮9^V�\���龮=Q������r�Y
]���.P�(W��s�s�I��;/W]b���E3��ZT*��!1y"�s��7��YO얥d�ݔ��{N/asu�_�/�h��[Fܳ�g^,�F��k��[[�F�)��w1�"�oGv��&�_Q��0Lе�ܣ�,�7W*��o<��=k�S��}X�*��N�yP0�����E/�f�bUt^�R�τ��F��
���b�7��mv��)�y�/ϲ�@A���9}}���;�3�����H�n�m�Y���e,9�ڶ:�7��]����Aɉ�����O*�}`��A����.�y�"Ŵ����x��y�.��ؘ/X�_y��x�L��؉<ɦO�ܦ�)\��hg#[� ��ᖮS�����'Uϣ.�%^�m����;���ՒF��\�y�o�MSx]V��nٱm�����n(���ee��7�@Ϝ�h�����;�L/ i�U�$4s��4%f�wYG�-��y>�\y+Ғ�D���G3���'�,Ui�a�6->��5�vۻ}�����<�Kԟ��fc"�t�� ��մ5t�NT��N|#�[KsT�+}����{IG:^�r6��#��8�\^^Iꋭ�^��#�`s3NC�]IY��J���C��<��4�s�`;}gJ�bɭ���>6���������������͊�9oI�k�X*Ǟ܉��DXng����¯e�RZzk�EǗ�[
ֈ���Ʒ4��ɕ����r ��Y!a�_�z�m*�F?Z�eK/���"�����˧�:�^X{�Y����:I\7�4�e]de۬����Sqr�׽�X�=M�҄�Ew]��}_}_Q��ޜ��9�Jv�?d�/���:J�,��t<m&)h2���\'-����fɶ�;��^o�����v���Q���+]�� �P��wƄ4��ӡ��u<n�KfL�3��:��~���=Z'�K<����_��3붌���<���+oѵ���.@�Y(=��N�R�dە�]�5���Y3��~�w5��JxԥM�X��||D�]�*�v)zכ�fqڊ�>�jy0����S���Z�Yٰ#���v=����S�tU�vk�z�9���c�����`w��޳��h��a�)�j9�ͫYK[�9���w���f�GvE-<L%}n����5�>�_��`����z�`�ڼ/�{;�zMG�y�U����3���	B�r�B���e#�:�7�]��>�	��Z���.jV��7�/2��z����	�V��UR�U��(�{'��X��[���tװ��y���ϻ�JK�C��&*J2�w�ĭS�X�Vjp��3� ^�����t��pB���>k�`[��c�E6�W���.�<L޺w[yB��݄N�?,T9;��������7k67̈4pf�>�J�[�Yρ�-}ݼ��ؕc�)HeK�+�U��.G����H���']�;���&�)P�8�-λ�U���� V=�Y4*��p�RS��5�\�v�\��Z��s�+J2��K��{S��Xx�Lc(��w��yy���X����I{��jf�l��nK�э�L�HQ���'Q9m�V.�_uɏ��6�AYA�*[j�I`s�[��P����$�#�lGy��;W��钵����U�����ޛb���R���8WK�Z���ܘ��]��6��ͮ.�@�cYݮ��e����3�� Ρ��V��j�]� �m�k_7\���b��������S ,0��o962ي�.��d.;�s "��j�Z��<F�`���lG+���Cc9C���>��S�-��gj�]Ι���{m�gj+�j�SMҨ$	�c�qY*��a-bWINn�L�ם��ϭ)�03�1�L���;x�Q�(n�Z�K0eC�y8V�yh���4q$���L2��Ķ����4�<Z0 ���F0)Wn����X���v�:�Ѻ��!������y
�}�Y��r��؍,��S�D�4����̭̎U��!��EI���L���gk$�h$�];���Bs�VeU<��[��U�^n�f�}m�u�Y����}B<�����
N��\k����m'dޗ�}J'�T �Z)�9�6�����<���ym����0�ޥ�Ab�^T�� �GU%Wl��k�6��-m궊�vP����R�K��k�˕w�qj�,�]�Ŕqps`��yTgs�Ev�s�t1�r���#1K�-^A�2Ro� ��:V�z�����i����ᙓ*&x����ݸe+{Mv斦�}����a�*:�e���1��A�oP�q�1��{�\' y���*�3��C,�b���+�z���0u�2�9Y����+����Z�I�:u9.{�B����DM*̐K���b������Ք��bZ�v[�5�V8���y��l5�Тou&�=qXB����w�u���
Qݗ�N
�ڱ;�ٝ��.<��A���-�7w�CiM���ʣ=V�=]:Ha拃��w-���5#K�ͧ�5�p!R��L�A�Գ�Ȇ1��RB�_@o����3lN���Z��4��p��'m��'f-�h���E�x
��lT^�oT�|,eiO�1�ٺ�M+��Wk������0op*�F�Z�_[سr�q��	���vj��S��ud�k���kOK�1�%{��4�:��r>��ֳF��gWS=k�٧���E��l�qe-�"���H��.�	�P�v��Hy�Z��o�k�wU�UŨ�V�׀#�Jy S��]� ���I��`@�*����G�>�"J"%����*�I\�Z�"�
��`�D�P���5Q�̬��[J��VTYP(������1���K4��*`�p�E���b��YJ�D��)U�(�F��ԪԶ�am�(��Ks*1�K`����Z��R�[V#��Kj�E�h�4A`�����\Aڊ���X�(ʊT�ZȲT����6R"��leQ��c�%�����er��k0a*"[dU[[
�e¡R���ZV.eDC*+kZ�*P�*,���e�"*4�f%F��ʍ��Z��E++��-�-+-�F��mYm��R-Coη�������=)P��iѥ3R��_nZ�v�s�B$r�μX;~V�����k
�Fs3(J�H�u!?Ͼ����.z/w�"���Y�۟Ϸ�ר��͞	}��@�WKb���t2K,��a5�����G�������{P�x1��{"�}�5X;��y�`��A����S�Ź���Ǟi�,��u�+��N��>�ʯ:>U.&8/��<xd�s��(h��=[��:O�G�k
j� W���;��d������
�`����S(WV��>����<;��U��;n�+�
�W��,.�<#>�=K���c'^�0f��/�^u��z�Q���y�����B�K�:�-n:��?Cb�o�a��~���,O�
[�*s+*􊮳'=�ok���H��V���,.1^��e�q��*����v�Tīt��j?S*���Wn�}!�P�.]��9wh<���<w �Ȑ�¡����,���뫯w�7��鏯��3)q�Zl��V�Ol�Sϔ^*ߤ$d[�b$K��������ƘW;yۣ4�3ᮊ�*���J%�@�fe�S���qM3�_�o�����K��6�;ϳ7N̓S�av�i�[5V�b�3��%�m���s���*�;�sk+�X���D�L�+�=�L	2�Y�[R�����t�5�}��l�Tz4ZmӲ�>��\IsE���}����לa��=Y_	$�
լ}]9Ku���BGZ�~�_?I����F"k>wdW�A�Ͼ'x���*z�P�Π��X8��<��V+�G�#�!��v��A���2�[�2ꠕ0XH����e��;�o��Qj�^�,l+쐠�3�29�\6�C���>���n@���Wn�[O��c����<T`a�1YD���M�)�͇ ~|��ϏS�H	2`~�!�!6|��NGHz^�_��{ R�SY�߸�&�R�zL(U�X�/U�|%RSğ|0u�}6�7vyz&�Z[������CuѺ�����>��*���c����_�3�	��'�(�\�2����mQ��Fj���2i4lM�8C`p����3�名X&Ьwu�_;��������>���S5�*��@�V����p>$��쥋k��w�10i֙R���~l�~7���Z�2jBW-���Z��Ϫ4{\�'>��a.���W�0�̈�;;s:>Zm�y/a�-K��KPV=����C#�N��jWi�~c��c3�V��t�#����A]_r��*w���ظ�6�k4T\+��5uذTPY�Iu�բ��U|�c��%�Ϳ^d�fx[��5�R�B�+o��yz��Kd���'�Mq�\YF��h�y�`Y��[X��@�F�#@"�uq��-r����}�R�*�{g����PU��0�@���ôtcUW��rϞ�*���g�����hnV��y�sawۉ��m8]`X��Va��|U�#2�jab���nX��BA%|�G{'�Vn�s
�����)�2m�ԫ�re�,�44c�u���t���FM��(���mO�h�eoAvńOO!��Wq}Fqbe��5�B���������7�z5�=��A���C�rd��&/��*�y�+��Ŗ��a̲��
�vw�����]ɔ'N��"�p��hC����'N2ê
+��a_O\��$9kJ�3�*��3���/�A�*��d��Q�����;X�<JV��ŵ�S�i���S��;�4�N�����H��#��QVWw����V��}��E����A���1�u�n�n<�q%k���p�^�˔�,D"H�G����R���u���OM����uO@�V�xo]W)r�<�5I�oMa�=a��t� ��R���i�{�J+ʍq�u0���{a̼�>FnVdkS({�Q�{	��k;�7�xRs׆+���������y��q<��������hG��RNᱦ��+7�-V��Ƚ����K0L��
���e���7���ַ����ru({�[�F^�I�ew�|>����w�'�#��瞆3��	^y(�fS%�w���U]�H�LW�	^Z`Sӛ�v�zܯZe�^�Y���D8��@��2V	��9�l����o�<�9ݝ�|��|< �4!4�n.^I���T��������9�������WF�ɵ�.G�i��Cs˫kI�?w����E�D�;I�ϗ�Ԇ��N�&u�ȸA<��\��{��Et����s����g޴l�6K�
l�+���R��+������4��3�e��sI�-L,�3f�q[]s"�o|F�}N��".Ɯg��Z��Ot�7y��<�]X���9��:��jq���ؠɶ�t���<�dJ��_�<�=���uƈT�Y���a�5��pyzN�2�6���:x�:���vȴkdz���3�y��b�]�pq��:�*y��R��2$*&�v�7�&�u�Nգ��Do��,oY��	�o�Ҫ�9�׋�ގ>%U
Ǟ�y;���p� ){B��.~ k�U��El��nD�Z�e#A��.��r4G�.6=ا��������ie\�J�W��T/pjS���Z�l��]O�K(_`j���u(�e]�<k�9Y�p�{S�f.�
I���~����.�N�t��\�e�������4a�|�t�ź�9;3=��(�>Ѳ���{�ܞkLF���~�����j��L�_yj�HP�#��,�<K�ig+��o�bE$o_�/.�������]:�7/2�3r7�!�#&z�`|@�,��a��zz��x�R��^��ge9��$��9Wn���DX��i	UF�	J���������� Eu>%�J�]�n��%��n�R���@Ə�u�W(������sE���|'ն��M@T
� �˅�ߥ��U�0bS�{��Q3��ǥ�X����[Kq�ʿ|�
�`c~g={���|B�t8Z�!u�ܱ�v���'���{;sX��w`�p^�=�떑X����do�FY���`uP�7]g���
on�����n��G���;t�����U�}�_�\9�V2}ױ0&:R^y'�Z�T�:l�\
���;Fױ�3�
�+�z֧S-���/Ł5�C|�K�yLݔ<x]B��y�
��7��b|Λ�v��0��O�.kpb�xK&�͏T`yv,,���䶼7��wwj���ɓ`O��R�q�)�:�K0;�즞)��T�qδ^dN��<�j�y7*V��<���樵_AϹ�C�W��K��}�˼�F{�5Z�&#����T�yH1Ho������o����=pr7���7�ŋ���!`o���v���&}��<� m-�>}fC��=���q#-M�ZP�ߟ���7ߜ����ִ�aTM��a�8�����?x�����~]-�ϟ��I�ѾZB��~���9���!X�n����xR'a��SYmP�z�{��y=bO)��<l�q��x�]%^�\V>�ܽ������"��[A��N�5/��s�ų;/����i�M0���������FW��u��򪔾�WT��R��	Z�{}��/Y���%kDX�P�e	^g�?�s�	k4���0�W+��J��O_bWu����gz&�c�z�D/�<���	T+E�~3ï��8���Rd��!Hmk�c��k���㷫��ڇq��r��d�,�ӕrЫ���c!{���SĔ��u� g��j���_>
oNgU��ӡ�"��t�dp�f�yT�U�2�U��4�Uֽ�j�'�'1Pb����V���u�1Y[MP�B�]���c���J2��y�:�Y���(�t�{��_���V�^X���]�/�ɖ�[���' �0����X����-w^�'�Zũ���S�[�RĮ49J�`�ĵ��}:a{����n;��0�����#Ek�TQu�@In��٬h؋,ᦕ_e״ɒ��ǣ}�t7�%'+����O�ZϷ/p�|�mD5�(לh�C����}c��%`���a�a̘%�SB��J]������2_��)���ac�P�8!��@y��ɾN���A�Zys�tԗ7=���h��g�`{`�����K��4���=��^�p幙Z��u|�y�j�����7�U~0T
-?���b��@[ڹ}u 
�[jޞ;�9����Q��{�+�M>�NX����^#
��о$Z>����QuOiw���L�k�2�p]���Nm�#�*hw'[T�_q��ţ���l*��V#��#��cW���av>�n/<���K������H'��
=]��>����5�$k�`�r�S^KO�����6CЯ�HL���nSӑ��7�*h���-��M�M��!�z��}�r&r�C@�,�(�V#j#�G!{2i�w~e׾Ӭ!'<�=r�+n�k�����x{!�h �ǔ�b����y֤(���.�6c�o.35m�Fw�*"����h���<�E��ؚ�陶�����:��[6<�>,�GG� ��J׼�����ջ>��9{Jg��+R��s��D4�@l9��t{1��8��{�s�o��ki3�X���4-;0�U���?��u�Uo�z��~���<�pH��{;��~ZѴgu�5c)��3(��yĺ\�9�o�]��E��ȽË�o���,wI���x2�����֊A˔�,F��3]_R���R����/�2|�k��]��H։�����'��d�ʷ�a���݊c԰�ﺮiQ�<#������,u�[�z}w3VB���&<�i3)�BJ���â��
��^9���ֈx���ZM��d\]ꦸ^Ww�<o9d4Ժ�W��z����X�"�',��Yx9�r�9y�7��yi���r� �iU����u��̕4g%PT�4G���8�xHQ7!Ǽ�n���z�X��Y-�L8Ms?m�D���Á�
�jCY��b�mmˊ/9;�q��g����0i�s=_d��M��F�p�Y�^��
�{�g<��aτ�i��}GC�+Yl�ju0[���;�c�Gף')]��ש0n��C��@���7���}��bvnZ�m�~�RO{4�Z�^gl��Z���0F7+�eAF��,dU�q���&�**���� f�Y��s�5��fЬ��U�,h����<c;N�6�n��?~g��l'e�k�����q:���.�z���U�&ſY���7���'YK�E��.�2�����1=o�6���:�r�A�Y4���ڛd���%w��\��C�4�8�HT��uÑ��>���")͹Xw�F�bt�ۗlM��O�_Z�w}HJ�����G�A�I�I����q���aBy���;�6�S�ses�w��v{i	A|�X��H�����G�����Z�_ڣ�bf�|^�eřu
�}<���gj����G>�\��������ʮ.�طSh����V��㞧S�2t��-V�S6�HUmp�3:���T,P�"�,x	�	�&{(������ܶk<o�n�g�>�u� 4#������z�*x�"W���DX@
�A+��l��&fwN����l5�\ej^��V̨�Q��p]��Ap*��Ћ�V�����E5<gU�T�Y�����~j?.��0u�	>���K��
;��|��{��z��A���v��$����J�Fϧڀ�P�yp����ѭ����6��[/|���QG^w,8@���k �3�a[f�xuP!�NEӉZ��bd�4�M8���0h�8�Ughn�P�h�c<4�XY]*�]��3�p��H�s4_�D�m��>��na��c��I�9yն��(�7��+@��ΕL�G�x��F��R��7�~Q.ֽ�"Qi9��a�C�[^�BK�t�}�:���Fw�c�B.�x���B�#ۻ���t�o�v�{�B������ +�&y�;NZG�T�kE���N{iނf�{Z�}�q��{���'���h���������0�Uz���u�i��;���e���ez�yU�۫.^�sfv{޺�qr�P�Д�qϖ�S�0��N�k�C����f��SY����9�|��������o�n����h�� 7�x���	r�C�?+�r9��ټ����t9ă��N�����\r�Z=�	���m�)��[�3Z�k4�Q궑�JށD.��F�48���0z����(=
%O�!4�Љ�S^��y�7[��]O��d/=�`��]&pet��暈ӱt����{T������B�GD�.o�����\�W����{��/M���-g+��L�g���Be�d�AV�b�k�ͥ�ǧ9^Y��72��#�X��R�/��4�	~C��hm���H�+���d� 	4{=�^w�p��^�)���I3[Y/qo&2=쎻e��P�҈e��,�h�=�ૐ7���g0`�;�ЩVK��V�EqRۘ(����h��vf��Q���Q�B�<���������9���p��e;��tm�[*k�w
�q������2�QESt�V;:�5�(�7��Y���X:�}�1L��1ܲ���t�钻�E��a�$� Ѯǩ�g�MF7x��c ���Z�,���U��+n��Ҧ�2�=��Y��w�@o&΁��=�e^�I�e�6k��ե���٤p�5�ʜ�l�ԁ2b�Qξ���&�V�zT�NދW�u�L�{>Zy�}h�� ��t5��^\�u+p^Yo䱇��eAD�5���>�� �U�6�(:��������k+9Q^W�qz�<Y�:�IP(/N�F$���SNA'TW��嶗Z��KA�� ��h7���p��n����Dc&��W[�$ɼnҳ�sD���v7V^����ihv>�7�YU԰��P#�J�v����-b�Np���ۆ�YI�R��ڶ�uM\�AR���\��ğE]Q��Փ��<$���ht�y��9�w8i�Q�q9�u�9g��/���������BV@;�2���N��9	�k`���Yo�;|�y����s�i1n-*9S,�+w4����״(�ŃP���ݚ�"�]ֳsXv�AϩD��X�u�[��x�Ζ�`�(ؤ��a��3�̶>n����LᏚWy�u&F������e�IdB����pD�ۮ���x_<+1�H6�`+���ާ�[r�Vʃ�Z� �@+VV��E\T3&��,�8dɎ�4�}��9���SJ�R��#��\��˴�s��C1���|��On5{𶊴kl9�4�})+l�����!�\q ��=g	�Y)�(�&Ӗ+n�ʼ�C��]�{<'k'�r	mm)cu�������o)g��Ir�VR3x��yc�N�EU.�ab�m�#�=O�{����T�o��W3_u����:v��a��=�ZJx�ˍ9V�w8w�����^��RZ艴+޶�֬��p*Gm�2�a�JҭP:��G]<aTͬ��M�Z����f�I�<��Ե��9�t�J���k�[�7F�$�{�M�O_`Ƙ��0��yژ�ؽT)S!|w�cޫ���[��jy�3��e��y*�woP�5+2F��j�٥EeoT	m�`t֭��������Dؼɨdgk��Z�5`L1Ψ��IG�˽݇%vv�<D���ȏ6u'�ټ]{�����z섷
�<�jBH䑇{J�;�I+t�\�
<;M�Z�WRhY�a��^I��}��1,9K�[U����E�h�b��N�3;��-nӐ�V�nXհ��ղ�_C;,lRi��19��pP\y���lLa�ײ�uv#�n�����m�b�XǉѺ8�4�ˡ����R�єT���fR���X�����ڥJ��m[,Ɗ.[-iU�K�QA��(��B�+Z�iYH�*Q��Zʢ�J)mm�Um*��(�D�U[JU�"[kc�S("VV)kX��mX"؍�Vh�b�R�
T�k�)hکbQ�UjQ2�EDEDUťm�Pm,b���DU+*ZQ���Z3-�m�b(��UDZ���"Lbܰ�D�V�-�`�`��J�+լZ��-ZR�ՉR�Z��YTR��űTJ��R��ZV���Qqp(֭�h�4��j�F1���hT����,n\\
���idm��Ҳ���[EkK[+R���m�*�UF�TT�#mDE�Zն֖ږ�U�Ԭ�����J�j���*��U�*XѫJԶ��QV˭�,cs�A],��Y]w ��(���/�r9:��.�"ѕ�X����p�k$Ȼ��bJ���y�l�����Y� ��V3Y�[�g���3�3��~�i�N	.a��>�^�i{dzf�{�1+��<E���O���n�!������g0���&S�?j̼ӝ�C\l�J�F�6v�]>/�Y&Բ����_��A����wo`h+�����.�&��ݒ`�\�حY����^)�A��#N��fr�{>�l�-�����n���{<߻�֍	�S�s�,F@�In����byhL�#�p��y��e�$�g�s�O�t�R�¶�)�L��=�v6��Z��/8�ԥO��ѯ�z���ڏ�S��)<����ώu�˿q̻t�Z�gjA�|��j�T1�D��C��zRu�M�c�h�-:It�LG�0T�2Ι�|�e�NC+F4�����0�9���<2�fz_!%hEvv��I�l!����9;]`b�cJVL�9=��ث�	Y�0՟z�ۗ���\�+��>���
qM>�NX�����(m��N��"���t"�7�����b���v����Y�V����+I��J¥`���++�
�ce笛�E�n���x]+�w�v�}[Ɣj�aʝ�L���lZE^�[��9�Թ�Ŕ%G�ǋ�Q�^i7W}��m�r6�;r����^*�s{����A�&�ޫl���sPr�ɶ�>��˔���/��ä(m�r�r^�F�jk;M�^z�/D�m,,2_�Qam�
��$Z"�X����r�k2����|�mL߽iQ���Z �Gk�ޥ�jc;v,"�WL�LN��j�ˇ�$��rK<�zZ����YdP�2��G���~>a}ً�Z���[^��
7���-ˉ�/y��W������Á��'�E_���Iu߅���M���6�Ps>�o6מ��+��L��.�'�x�N�aY2��xXmY����d�e4�w�5M�g�m!3ׇY^�WsMtϴ�l����
N���֊N\���u<�Ě�
]�=w�b���{5�(�f-��+r�j��/+����\<���5X��C���:]�VqZb�L������\~ns�n,�>f�	�C�z�c�`'�J5��LR���9�Ev��C�s�V�u�/G7���բ�W�e��ks֘(�^��>
�c"�{)�@�^s%o&�y4���W�+7]E���eЭ�X��1W�n?�����I���8��{Yu�S5���\ĩ��^�mnt�m:�bN-���j�s7|E`o�}Zy�3g{��X��&|��9k�t ��[�XE�^d}8�K����fj�D�ͩD����E�{�w;�>��F��b����U��e��Լ���S[�=��,�e{=pOf�HH�7�k+��jY	ʝ{
X�n/Ä�:���M<��Y��bo+b�E�O[���~Ȟ^�%دm7�����cG�ZG*��ӣI�z��K��<w^�.�}b0�=���x�j}�W�[��om	-�����X��j��/@�Y5Ѹ}��%[�J�^7�9ŏ�ܻ�4�&�
;]hE��g/����h��ѕ��v|��<kr_'7Gem~���o�;d0 8;Ԓ�EV
upX�w�%|��3&�R���ە�{�)l��X�ށ���N�&�{��z�hWT�n�D�����FC4���a�kI�=���m�{�xϨhp�9H:EV5���i�]N���!�*_��BRxu��χ��ȵgv&�"��jy�6o����`
z��B���&|U��꺶''7w2f���rwL{��מ��j�6�	v�pry���p!�&bڛ�P�+�B�	d��~�:*��O�/�`@��^V�~E%�y�z�kD�!�G�3���D�:=����QK��;��!��>^yk��5���Q��`�D���

/���nX�w�rwK�ҩ�wke���n��{�S+�p^r��C��������ε��ר��S��E,�Ϧ�q��ܼ��7!��\&(:e�[=^ܽ[�u�^�{V�P����Bˆ,	�{�H}�t�d��^B��'X�r�;k�*�t<�����d�S���6�!P�T���W����W/A���$���(�@����W�h�L�;w��Sv����1�	֍�O�P/�R}�|��X��Y��O&��8@�.��.�m�3��E�V�%�:O�vt�˔�yg�3H�;(��f�/b0r�s�#->^P�p|��2"�0k� �I�|�j��kE���y���A[��������G�{��U0�W�+Qu�{T�/�_������LgF�Ֆ8�	Y��|��"c�^����h[�KkX�Ct,-	p�F�/m�.�9R�/NMjP�T�]�x��3�M�=��J�(�����XϢ^ *~�O(�P�˳�k�
�����^yYsD�f�a�<w�cG֫EO&*�GǥRXI-���T�x ����zi�3�i��?�ɽEY\�:'�k{�M�yu��%���y=���y��؊�*aK%W9i�kH��i�W��6��9.�>�y˫,E���n��;���h����֫�1U�)�<�{Yq:��X` H�s�����Y/C���}Y�F,͊qר�}�l|����'�x�4�4�9���j9C��&�4�;�� ������ʽ`%��#j`��o%r�Zg"��l�.�82��_�c��V �v����/�o��o�/s��E��m��\��v^�
خ��y���zX��\˯DB�HЫ�馐;O��>ǁ��%j����c/,Xח�+q�4��~R�����s�%�*7�c�&�^V�?w��A簲�'ۂ�� ��F��9��5GYBg���%���������2�W��*�t��w��dz0O��x?@�_o��]%���Y�����A���>>ˮ����j-��c�]�T7e��	딄�$�&���-�|n��U���HHjIi��δ%��� ھ񔄉1Y%�).�W�;�Ӥ8���i���J�
�T�w���ƕ��v���.�� �����=%�)}���B`�#���g9�{tq�m�W5�̾�c�>5KO
Ҟ�ઙ�Gy�ڈkPQ�8Ѯ�)�8#_ �8�[SwU�j3��`�4AHY�N���"�J:o�ҕ�3��G�wv_:tmF�*�����J���@C�G��e�.�2r���3(��,�{� {��!/^�.D*!$�.ŕu�p�u�*0���i�b���3��k�7e�s���"���V�\Y��~����H�Mu���#�k�^�֭y��V-w��	ޑ�&�4Ү�}Z4h�W"6}�ᄹ���/Puإר����h�id��z��>�&�<�]��V�{���}ko��XUf�@A!�n������\��9Zu�ql^jFU��6���ۮ�q`~����u�g:��>,V
ZH�}k�A�/(��m�r��y�2nƳ��
�i5ոNMR�.v	�ܛn����.W`�\Bk+��W��7ա��7��d��7w�	�EW4��%�[�p�]��u�~��kaUJh�}g.��&[��Z��-2<'�v��)oĊL���H<���'+p����jT�4p�{޸�GuÓ�Ow&�*\Y��%�}�gE�;N�#���F�aOj���]޲��Q��M�x��<,��n���d>�\*9�V�:����Cx�$�2E:�l>#����h�z���wʓ}'M�Ǌ��5b���/8�%�"�˘rxXi�"�s�L�̦�)]m+�u�9R�vg��Y�ʊ(�z�33��5ݬ-��Oh��V���r��`���Q�3kN�q�gQWtܢ옣z�*/&���=�d�P�̓�y.	\X�o;B#P�<���^ۘv_H>%I1o@��8p��'q�ʰ��ӡ8��][�n�sz�,�����X��Og�9Wn�,見��b5d��]_������ui��ܻ|7�|��F�a?[���&T�<�� g�U�FQ�_K����؆g�#��)�{�~W�# �{�ië~JB<�C��t3;�P���U1JJ��߳i�۝��A��w��\� ;�XCF��z����F���K�x9��R{j _z���n�
�b�Q"����(�õ~�D�'h�i���AεA~�x^Uqpu/$��M�G���u\��%^�lr�y�H�2�+�J���Sǀ>x� �j�2��ZǄ<?g��n�S>�'U)smq��lU��9�|��^f�S��x.^��D�{<�tF}5�|w%���zs�:J�����O�y��A��Z��w9���PF��VAj�����Bqju0[���F��E{��1�M��X�Z�E5���<�߶=���k��B=a�a��z"��h�e�{N���T匮�ӗ���t���r�������7�243�h�Ic>������c������0Ân��ιV:f,>�0�U�:r^��<-X����N^��k��O��锈4U����d���z�h��M����-�]<��ЍfK��.�+Wu��v� �b|e3(�gg3��Do�!	晆�T������ƣ��;Z=Z�U��9��Z���1�1���`s���9��p�X:�m���Ih�i
ӫ�f��0X8��=a6����*���â�D.��`ַ�>��!ׁA�E:��*km��i
�ej�鯹�O[��jW^y.��&���o�;�~�(CT$�"����H��k��]�����!�k���f-��1�����pV�.82���>��0h��I�߭�3�(W.T(P&m��Լ��z:ݽɕVb/,_W!���X&�Y#�k��ͮ�f�6��Ȍ�g�ல��7f���Q�k�L��:UBK=E}fC�A��q��t�G5!L�����e�=�fN����-�-�U+n�w�{������Z<3�Jx�;3y����:$���<������a7C��^���$F�����~��0u����0tPn�{U)����P;�"]�9N�yOǫ۶I��@�a��/�|#��}��T�Ι���5��h��2hO���H��y�4g��%b^�F�CD�s��p]�I�|
���Z�S;|t�[{d�y ���Uy�pPh1����tHm�hg�JXzJx��T��U��_�U{��å#������V�\��K->�+��R:�דY���0@2�TT5����L���B���x�5�^k����p$��n4'h��C"+��o�`�O\&��q͝�%�tĬ>F��2���V�{D���њ��2v����h+Hu�d�榌Jn���C�(g��|�Tu�i��>�60-N�ja�xS���}���Hv�~��o�'5�U���bW�+�&:Uޣ	����,X\,1]�Y��_8r���,�$�w��Ͷ��wh�/N;�<<3�:�V�0�7	G��>1%�ҟ�ו\ y[�^�����i�#]�g���N���Տq`Rd4.�i�O��ྵO��j���ޯkoح�o�d��D���u4��"M��R�3�:U�g�����K�9�ws����/57$Έ��=��LVѕ��S���A[�E�.�o��#����2���IuOZ�A=��毬��`�e��,tC"�-�4�K�BM�̨'��9�&w�4�P��oI���ֽ����z�Ӳ �H4(Ӈj��Aי���`�塞����`��7���/7kZ�FWu�+�OrSj��L��G�%µ�c�����8�s{{��\dd�R_=�~���wY㎛����;���L�3��yF�|�]g@�f[��
)�{�m��|V��3�-�{,wإ�u�L�;K;M��+m��&N��^UpR�,U�s���R�KF��֙�b=qх�Ӱd��z`|Qg�鸙��m��O^^���ƣ��ꐛ>8��x\�2�7��?
}v��Q�R�b�٭��~O�#���L�g��P�����`Y����^)�A�y] 8�W��ǵ6,��t�c˵�>� ����z�umDX�(s��Qb2��d�t��S�G�E�������Kʲ!��Qmi�)��u#8;��P֠�K�<5�C���m+�Bm�ov`�k���M5V.�o���2%��*��/$��l=KO	^�V�I{�tO�y��D�S{�פּ�< �۶x�Wu�NC���*���&M_<�:����ǁa7m��ڼ8���?ӓ���A)p��Vv;G���ZT��	�mpEI�b�{W��[�a�2����粞�=8��zV;�/�}C�[+�>Fmߒ�ɽ1Ey~ܿ��Z��!h-�'z
�qeM��aJ:��c�U�4���vo��S�;���V=PP��B͉0�=��O�|.	�=7��/���h\f���	9+�iim�n�i���]�8vF'S�w�h�韞��������k��!e�6�w��m��pp���"J��J�:�t��F[�K.暲���Xc�1��z��y݁X���������-�D��U�%Z���sd���^\#�7�&Wh�U��[9���w*ʉ�溱��.ǔ��7�bQ�n��ܰ��&q� ��m�X���N�ޮ��F���:��洪�c\Ӱoǫ��i�P�EO�6c$��ΰ�&��;�Op��]b�L����j@ղ��rDͼ�vg"]�쀍�;6�wj��I\��Va+���<;f����U�)�vM�G��t�d��V:mq\�c�n��]��zd���ktWd��.�n��`{��n$1KiiF����F^Lk�%5��WN����BQ�ǫ��]��VR�Tn��n�{:���w
&�:/-8��t�kө�p>m=Vrέ�
v� ö�v�q�O�%�Q-孚2�;8�5ƦP�8>���˩�B�}��)�I|-��{��A|�qn�v>���-v8�6�G��ib��9 �H��c"vH3����̺Q�k7{j4��36�]o��n%'�IWK��eZ�1ֶ���\y����9`k�+�FBEp$)��;�v�>eR-�Is�W���.��c�]+��7�P&CܢKb�b+���R�:N)���j&�ah]�R$�u2��z:�df��\S:����/{�[�$�.�p�[σ	�� ����!��&{�����0�ga|���	��G.��V���·�]NȜZ��U�Y^�S#��U[-�1WZ��":2�]n$6�b7���-�P2�9w͋��˚*�����t��V�I,%��h2ғ��B�m>ݡ�����$��ڵ2�_W`�;M������̥��:����PB;���1�q�mD��ma9��6�6*r��RevM�tѨ��j]h�lS�MD_ܝ��u����ղ.)e�߻u���U��%��D�](õ�!��VX�����u�Ay����Wa�.��Ov�Q:�>yS-��Ͼt�5��������vv�
���\��˵;&w%*j���<}0~[��z�*�E�b�n��Oi�oݵ���+ۨ�e.��cqr�0��{9�{�䰮_�����"�4��M.�/,��Ϗ;Į�͗k.�L9&�&Z֯.c���7),�"ю;�"�rI�q�O_|�55����])���v.��b�vEenr����^�ڋ�J-�W�kX���������]��[��%�m������z߬�k*V-����QX�q������l��{�W o���]>���8��2���yl��c���K]6���p�Yݍv �[�cM�u�$��+��7Tx�g�j��O�v�ޙ����^l�:�q�C�q��q����sJ�ڮ�Ԭ�XƔ�]�zt댰Wa�6�����/��D�KT�����Q�	�f(�m���Q�[���Die+UZ�ij�Qc+--V���U�E��m��k[m�jejض��!��[J
���V+m--��iaZ[X�F�
�V�KZ6کYJZ1`%j,hҭ��jTUV�,Q*PV��*�mQ��Ye�[F�J��*QF��V-�m�V%����J��!KZ�l��Q��-+���ڭ�
�)JƢ�QKkRŴ�ѭ�����%���m�ŭ-Q
��KQj6��ԭm-m�������R��R���X��+#h�B�*#K�*-��Kkmb����TD�±E�-�jҪ-A��[*��TmfZ�0m�KTiJ��VKT����U�-J֔UJ[*�ʊ���%Z���J$h�+q*(&#R��cKF֖�[[e��6�Hv��V���j+#wN�Dl���7���E�̉�P��9�ۮ�;���#�5�� �c��\\OF�������oY����n�w�䫪����
$8�L��]M𝆥/����ǭ/;n�+�}Ҧ��w�q\�.=d!����N�"�mQ�H=p��C�<"��<z�珷�@�vv���P���U�MY̘O��FH�B���6a�B����o ��9��v����eT�{���;Y.a�S.a��a��W��2U����6v�Č�Jzr�afש��l�~�_�{6�>�']�b#²e�'��IU�V��z�Ɲw#��ݚɵ�y�|�:�}�ڍ1�Xy}�Ȑ�0�7�@r��8ʕ��9x���߻x5�ך�3��T2��Z-��/��)@y����=An�	�y�ϡT�-+�v[4r=���c���?�����"�Cֲ5�x�屻��3�4�)�D����b�8>l=j��Ɋ�0��5��ɏ�*z��B�/����^I��`�,n�yOV��x�iT7���s��K��y���/n��^��X�W_ڳ<�S���
�%�2���Wʵ<��Zu�R�Mse+?�qI���}ǘ@Ľ�I�V�������DN�q�E^���	�i�|�1j��Nȹl��_$jf�X9$�s�7i	��CQn2����/�=�%����̪w1��Pw.[��I���WOn\vI���ӆ���]���Q���1�P�zsN��{ʙ�;�5���\�{tؤ�n�2�U�J��.}lEnf���U��5}�E���-����-�L����ef:�_�Ĉ(e_T��������V��9u�svp~}+l�z���Q/�ا����c�����n�`��fY���,r���&{�Dw%��Cp���u�AjG��W�w�5���=�>��Y�P��]ک�+���n��L^>��W�i]��*H�g;,�kY0���g�S�
��͜#IW�:;�U*<=������x$��q|�J^��B�v�<u��c�S��|��: ~0Sj{ƅ�D�S=�}}c-jr�c#�K�ȥ���P��/V��άf3���fh~���B���;v@Lw=��y����P��/�#�}ul,W,��Oj9u�Լ�i��P��B�tMW�=����3���w�����Z=�St�ԍ�]Ea���Q��tܭ���ܺy��fV���5��� ߊ�FN�:��}��֍�A��u�v��x���I�������"�HY��`K��,�Y��sjuINf
i�����e�_RT���A��3�B��ڕ�A�Fc��_h��W٩Ji�g`�J��e��V�w�&���	��ʼ1�6<'XD*+a#�<�ּ���S�<�*��38���j>�占I��
��c�Yg�8��:�o�u�g�P�����u����)��纺�;���V�*D���'�;:WۉJϟ������x��n�sn�k��\��o��#O�������M0ub^�F�4Os��p]Rg��)i��t�n�W���{�̏��j�6S3�>�-�԰�GVِ�m����«՞qᬛ�7MW�S���4v���'�{8���y�rݚ��6�j����iX��apI�ϸ��Z�L�ߦ
����̭6�Jԕ�T�V��>���Yo��@`��Bc�Xϧԗ��Wx�aK۵A�������ۙ]o��s�@z'�S�^�1C�0�ۈ�Ғ���tyy��Z�Ļո�y�~��	����/��C�N[�݂Ǹ�)2���>&C���7��շw�s3s�M�^m5^�ҭ2�$(��ӟN�$ر�r�3�*�U�r�Z�X�_���9yO�t��=���Z�CL�21��7������f�Z
����7t��8���x���4Gm�2����h*��Khq;���j��U*���d�s2���{CT�w4k����-ɖF�J�2�^8��pⷝ�;&5_0���C�W�������S�(�ڿ ���d���:����3���V�d*y��pm=�4f˧�`n�s��K�=nK�Ů�~!�١P1J��fG>�"�sǄ�)Z�ZA|$�����b���VZ$Y^�~��φ-8�J���O|���L�U
A�F�;����ei�߫T�]S�n/t�F=G�����L���W���2����,�[�x��
�~�S<f���EW@P�^/[���u��i�g"Ɂ��		�������I�,��]��V�����`�[�wG��=j�*�%�*�tD����Rb�K44S���<J��Z �}�pN���gX����]�:}K���x/�R�p�ӣ���29�Qb2��[ z��4�,Vs����8�r��j*~KB�+w�^���B�=�c>��g��]E�AF��q�;�������Ӳ�^kj�����n�h�m�x<L���~��k*^I\<�ac�-CЦ��Ї��8��݅�YZ�K8G%�:ݻ��{I`cƳ#�u���y���4��oY�fV+��u}�Ͻ�
�Y�Us��lS5=�^3�Ȼ�ާ��ns6�}A�����}�S7Y�T(v8���=�����"�R�1��%],������-��P��Uњ�a��줛Ҹs�x��d�*���U��`����+F�{+���~x�p��>9���<̦K�g��n����h����e��%c��\�l��`�z����cǨ	]�q����Y{n�r�}�8��
��zV;��a�
,�t/2I��Z�œ�ܗ�T���P˂�.�5�j�&m�s�O}N��c�R��ʙp)��9����!�[�^�G��+(�PP�<��ׁ(+�aa���v�XD��W0��FR���<yr���{-N�p_����r�1r�S�$Rf��-�񓃰�;j,#�*T��_("���59c��oj��:'e�p[z�BX *���=@��A��Y_Lzx儅f*�{흯5g�f�WO9{0ɷg��e,9��l;&�|��I,Fz�W��v�y�׿q&�d��[~8���%+Y�X��
n^q�K�E�	�0����"��L���+����4�$�j�Q.���@�C9�s�˨��J~�B���K:+�\�u6\���u<�u�[���5+8_�;�z���F��j�����$>5Pߙ*Am~��"ݞzhG�.�j5� !���s�T�u�ޏR.%�&�m�k�����/q�z`!�͕��s�̭��4r� 3�u0hを���)
(�[QYw�I�e��e����R�F������gnGaaf�1��\	��s{������N8���rs�oq)���c�;֐��5�����_X��<���ts�C0wL�瑛�.��=�WCo��M�׮�T���&}]�e�8:�"�#�fS\/ܶ7r{!I��Aty}Y֟[urr��|8���`0�ӑ᭥��V|0V�x6e�x����FPm�gtֹ[g��.�G�H�h!�=�s8&���o�L~쵈���~��=���1��Ҟ�C��gs��C��g�Z��ח/T���j:#�1�P�|t�3�
�գjc��c���3,�	�<m.g8�+~�ip��ju0[����k�����߶�6��"��M�
o+���/�j�9gQc����(+m[�r��EmN2�����we�~���B��7U�����L��x�P���;�b� y�Jl����~�f��|�̣��c:ε���|'��&k~�]jʩ��x-Ĳ(!!wkG�HV��*gl��Ӧb�:�/t�}Ʊ�b�ֽ0�g"LR�\��*�u����9���#�fM����h���B.�#i��:J���)�VS�ھn_cT�][�j-��W@bG�^�;N�7�s^5u���Lu�b2gfwS������X���������dU��A�f���g2<Z2����� �B�.�D���q��W&rR�~}�l{+�i�[�l0��j�g�=��OT 	.ȥ�o�qgof���������h�*|e��b�2�z
�,������}�=�4;���3�㺌>k�/���Ե�.�9�]
�NUYP���+�ew�b,��!���6�ш�.��@��/�Ff�9-r�����"V�v|��0.����e��A�C�w!�t�g����S�k�.Z���og./^��k4]�3��*ʗPt�؃i�/�¶8g��x�:�A��3��m)w��x9Ǳ!�NK(��.
2{·}%�v�w��~	����*C�����+��:�<�8FdEWa���R��@�h���ݎ�w�t�k��v�vY퇴���5VM�z���6jQ۬���N[�<�|G<��� ��~�}��/��A�P��}���:#�!�5{LR��H=X綥��6�d+z�@�/T��V�ǆ��W$���no��?;���V�ū,p�6"���2�V �X�LV#a���M
UQ+�*����ǝol�6�������a����Kt�vQ�^���ǔj�DE?Ssu{���������}n�N� w*1�7��п.0c�8�6�{X�r{X�
wD)����r*-����vwd�wsU�	S���<�����-p��'�s#w�Qs׶��xO�Fq���Wmz{�����j��3�ܭ%���Cn�\BݷI��ۍ7)_>G�L�Wӊ�3%WK~,x��κ��YAxO�g�XT��㳆��7�;K�<L<ZWkhK��+4�l¡�D�N'���d[!�CO��G��W?��N����mĦ�o�������|�U3�jBk�<pN�'�ŬfԺL�ϺU�r�`�W�ļ'��~<�kH�/�X�K'�z��Y�hV�u��SO��)C��r5`<��pm=�4d�K3�i#��j��ۘ��L�e�k�H�u*�'��,X�.E�|-�4��~R�������<," G^�#�ƹ<��jx��t�yUJ��`]'db�kƮ�>��}Lk+L	�Yԯ3ѫ1G���:<�j=\2��GWOd���x\�&U����%]�g�:�j��~�,�R.i,�)޺�=N�j �B��Ϥ���,M3���b�C�v���s��8ⵧ\)׷����U�_�*g+;�$�p�x)1RC5��H>oK����ޮ���=E�tk��f���f7P��4Da�̾i�wr�K�֜e�NW:T��e`�����uX���wH��l�K����d��K�[�[��*�ɚ���6�]l�l��i�v{3b%����ʾW������6c�|�]�I�룶O	�W��⛶�"�ÉO}\� |X���� -bƜ��]g܏c8��'6���!^5+5��Mf�S���x&q��]��c~֠�ES#���[����t�z���f�w�U�Ec��J���\/��Y�jA���X�궻��o����~�FV����V��L�;���G���1�&�:�}��<�})a��8����=�r/O��@��2�nfV�%�~�#Տ��+���yw�C�b�Ui]���۾�[��/�~�l�}� >��&}n{)ӗ4�8_g���YJWp��`3��������xg�q�Ԣ�˂�.�5�=���T��s�O
w&ۭ�/Y�U�,��b�آ�M*�x��[DuxP�1Y������]2P{W*o�a���ڕ几��guMn���w�h�9ݑ� 	���3�Hq�<+p������e�p����1;�|/��_C[f�/�ۀ����xXIلx �ƍ!��5�ˠb����{�J4-�\���G���!7�}��}�n�;Z�um<K��k��^�_JE)��;�W�"������Z]M�;6�Ȧ�8U��q�>��a]q��ۤ;�]N�H�l:��<�ۧ��b�f�L�#Z`�9s�y7Ym�9Y��c�L�ô�tv���0�	p������CVEN���z�r��?~SϜ����J�X��2��$��JV��-����d�!=���\�3C�[fR�\}��f����Ԅ2}K��s��k��Dzj#<u�Q����Ruޖ"<+&\�����JhY3}L�#�Y$A�Wĺ�w+�j��LkV_r�#����ߙ����ۉ�5���[Y+y�{��D:8j���JO*�E��e�Ձ)^~��=�v�fRS(�W����A����<�a���T�w���U]:\khm��3[�i�H�^�I/���/���y����urzd����j �Ք"�U��xa��`d��LSu��>���`��4�D�����K�%���<���hk��c��bm�'��mjۃ��O��m��J�����w�U�}n��]K҆���!���0H���q�N�9��ixM%����F�~ؒ�B.�<�`.�P�7=ᲆS��.�S���ez;�p����1�,g��<Y��ͽ�B�r*���Uލs�P�ǰ�S���[��^�6_w�Y���)eb�2� �wK��X:�y����Oy�3yV�c©��Hi�S����ᗯY��k�p;A3�&m*�Ոa�p�s�����zeZ%���/N�PA��T��b��Ǻ�J�����5�YQ,��U͍���e�{�W}7X^S!�x���;P�Ň����KVI�	�.\�seEDK�n�C x���F<5zH�h���r�n޸�^���E��!����Χ�G�Fh{]Yj:��}��Jp:�k	-ݛ�]���M�8�tQ�ĵjQ���.�J�g��W�'Gm��,�͜�ɔ��*��F�(�b�k�V�y�r�n�]m�4��b\!0�nF-�E�W>�kW�
�P�FqY7��*ifuYm�|�f}q_[��Z��5e� gG���N������FR֢�+�]&�uo.N�U󗢭���:�t���z�A-sI�j�r���X/�eu��w�eـ�cm+Hp�����-�6�S]�&�Յw�k{h�-��9�\�a�r\�E#�Y;����,�t��權	����3�4��=
��ͮ�yib�C�W�:N-ɦf���s�m��WQN��E͘O&������Ծ�F��֐��
!`���R�?�sDy�r�ԫ�"�J���@���v�U��ø�-Ұ�8b�ҍ�z�9�x½߂X�I.�Ư��E�Bb�u��Δff���
22�e�!be��meXI��̈Č�+v6�n�8����N�-ݺ���Y���2��mǽ4t�mi�)��e�������ٷar5|�ךS�@d�R���4s��TF��aԘ��u�;�{B)�gys�Rݣ1���3��|�fY��������׫�l��Y+�+㢍
�9<��F��o�b�b����b��鸉F�8z���)5ӁT��e.�r�q0�,ގ l��Ma�@��z�ȶ�]sJX���_w5��D��P��m���ɣ�6	���N��'F;0Q�bad\.M�bx����t&�n�C+3�u�i�ZS)�'F%*�holuq��7��WI���;�\�Zha㼮��w�ɝ�x��lX�FfB�8��su��F��5���ފo9�4ږ�`�QU�2���e폸�]t))H���cnٽ�j�%"��;رn�^mml@*}*v�M��Zo.�]��]�w*]-���T���ƶ6�d�z�d�ZzPyw 佼�ި��U��w��]���Ɔ��l	dЮ��֊�n��.���ʗ'Q��ջ+%�Wv���jԾ�/+�:}���ᒡ
	�6Q���֎�j
�.G[�4�Y]�3/gL�k�2tD�]h�vNp��gs��aT��)�n#�����<��]�.��:V���x�8;�n��dt;�ճk*%+��r|��ic`EI;�������ͬY��<����o�4]�?9��>�V�
*�)ek"[lQ+R�U�e��m-h�*��J����ڲ�9��m��������ib+�*+j��Q`ҕ�
 T�E��U��YZ���D�P������J��ThȰ����mZ(��*�B�b�TR�*�EX[`�IRTPT�(��-(Z���d�qPF�ij(6���cr�-�jQ�Q��PF,˘PV-��Ymm��mAdm)6�V
6�+m�VJ�@�)X)�*�j��IiJ�T��D�U���FTiZTm��[`�
�[@\AT�V��AT�mXZѴR�"���"Aq�L�eZ4jQ��Z�dZ!�3,PEaY+R��Y%k�������fb�E�d�X��")m�YYZʩ
�c�\dY+%EX�V��V�-�QQP�
EP��2��j~S��鵴��Ml��*5��h�#�|�eq�Pͻ�f&�ub�ugep"�MB4�[�t|kC�������L{&~2o�*Ţ��}��|m���qB��AY�V����L;}��ɷ��km�ΈR�h�k�����FF���{),gҩZ(����0�%R���~�w������i����������.y3[�B�V}S1�E�G���2�%��W��܇�t�}x��k5��e��>��&g��a�Mk&�g3臩��v�x��VC�^���x�Q�L�V�YK��X;Q}�*�-��Fx���!��	�y��}<��a����@�W�o�۵�9A���h�;B|z�yWV��b�6\�_���e��{��j��L�;^�>iZ���$ӭr�|�B���
�'>��Yun�g)fVM��0}C_�������ZYz�X��Z�-~^(A���=eT�
t.��]������$��3�2����Q�z�>Ŏ�4��#�e'��J�\0K�	�T�~�5t�v,�دۣ�e����5�����OW��T�gú`$���@���b��,��U[Jg�=��b�+8je-X%���CQZ*��q���a�����u+C���Q�.��WZ�	�/���>�T�Sf�a�os�{ۣ�B�'�1X�r��u�p
�i��J�/��w|�1Gv=�73��U^j��͇5�Tm�4�U��=��>˭�=��u�sek{�1�[��ّ:^��=SGX�egtD�5��BD�
g����ҷ�0هr�[Ю���<��rM������R�-�~��>��qGE�:�� ����(/�����s=�f�e�j����X�q���g�V�ʖ��-���<��Vח�@᱁��W�����g+[�_����Uݒ��(rݚn�o�^=�ǱB������.�ɴm�]g�<�_M�p�۞Ǭ�j�0|�}t�V�]��E����}�2�'�*�r4$������57N���BV��Qw�[������.�kV�T�!�eNճ~��u�����Oú�s�:��ԕdQUXL[��޳Q�Ϟم}�&S���ȶC�v+N�M>Žm�I`�Bg����7�鱲���.]��o�2�SNN�'����.�83�ZGs�ԫ(Ǐ#��m��ҔlV���J��'������k��y��[���:Z�0c��}5�īc�<�1.ϞW�v�m��Pb��fe��.E�n�K��#A�����}�����_��4ǅ5M!WAXT+��v��`�dIjI\S�!�W\7s�u��I "��n�]����ӵ{í��Aҳoz�M��)�-�JJW�:�G��Xλ�*�}t��;a%l��Z�r����Ž�a�Cb���Wdܐ�P��.�*f���i��ӛS|�eM�z�s�UV(u>@���jk����Y�:�wh. �~��i�f�+�b�R\½�M�0dڸ=0YJYd��إa��~����e����kl������_�]E��)�	��!8��K� owɯd�ѭD�sܧ��L��B�۫ҫ��tT�VwDIO�I��,��I˯��*�/�f����3�L����"L��<U����$X/7m��&��W�� |X���J�ձ�YM�{���5�$$OWD�v#{���\���yd!g�gQ�3��]D�{�a��T]v佋κ9\��j�^�̏}�a2�̊V�ׄ��u�W�J�gZ�Z|+h�Muޏ"6z������*}���s�e�<�ʝ�a.�A:K5� u�+��sG%�&���x�{ܗ
�-���8��<�����}����:+E֝>����"����Y�k�꺾0\�EdUW��n��uJ�ϯm��n,9sŁR�/MԾu�*� \�9��Ju!lF�h��J	�@��4������xh��Vq�ON��6"�ńސ�m�S&U�����4�U���$c9*P��Ն���n,�m9!�ӣpnV)�����20�`R��9���%]����m�Hɻ+9>U��9��'9s�G�(�"#�\��^����!3m��T�d�@fj�{)>�LծwV�{�.g��l���Xu��������]2SڹS|�5�y.���[�5+j����ʈ\g&Y�Q#]H�\��|Me���$+}0�^fꅽ����PjW<!��ޔĪ�Y����ç�#C�0�U��#���A��sX#�7/h���6_~%&+߫��? xrW?vV��8�zׅG=%l3�.��+y�NOչozo�����s�.3�h_�HPx�9�����W��n^q��s���fQ���]t�Zvx)����:���kI�_\��)\��M�kaϙu�=���v�*�]OA��O\ޗw�_��k��P��܉"��Wīw�|�իڍ1�5a��r�%�������gݞ���u�ʵ��	�-"oT��)�V"/�U��V|��/?vz��F������q��J|�-=΀�ggCa��H-�9T���`�2���������l�Ω��������\���k���MÒ�����2@j���,�&S��̡�(�S�[3���^�m�X�qzg-��0��e� ��؆.�2=u,h�շ$���2��v���=��H�ݣ^�k�).�h<�u8�w�D��9dq��Æ�)f�Oݗ�w;��a;�Nk����(D]x�xkkVܠ�*}ו�"�������S�{��lK�<�z�������P��s�u��.u�(�6տ�{�EKͮ�����q���17�
&�w��Zk������#���"���L%C�棢2k���'2��W�,2)����'��{���k����*�>����+�\'>Z�L�3+��b�0���2���ɑ�p�'����+�~F�K�j[dS#�Pb�E ϩp��Nk��kK6�i��VŅ.���g�������ۏG��0rX�4GP�,s�UC�wu�������k��O1�8�\�f����aY���<.�_�%.�rC>=~�ҟZS3����"�[�`�5��1��L>��s9��AEV54���s��S�D��\<]���������T;�A�st�'��a�Z�E�ʵ�XU~�нѕ��7�� �x7ܸA�u=�V<x���t�ź�����K�=]��pe־�%q�4`�ˎX�<��������n;��97����ʧ�����o~�$�e���e�*��{OP����o�\U�1{Փ�h��]� 7�'�΅����^��^y�R	�5�6����;j
�KC�Vv�n�m[�9]��'�u��j���c����N?>d�w�s4vq���w3��(W�r�B�p^$�3�b�r�9K2�lE��8��jo���ޛ��O�����k
A��FL�+���� Q��t�x��i^�~��=h�X{��b�wӭt�=;�k��x)/!Ф��J�\2X��bU+�"���Yc��`�ϽQ(1���k�g�nN3�Eb?��D�z��1��,�� qUm!1)Y�~��]��|yN���{���+Ԫ(Ԥ���T߇X�egtD�5��R �!%��v)l�f�Y�٥��8}�@X��6}>���N�2���<3������� *�q����&����oe�9�QM�-hBx/�&	�mKх2���FB��T.^����W�E��'�ċy����9)�d��w�;A,օ��0&:RW�%/:�p�{M����v�,d��Q�r�[�/�]�Ԇ��;ǰ�g?
�~x,J��a��LtI���3��4C���
�-kޝ�<��ۂ�
A��0���\I�k�񐺕�ث�[L?��<�%��S��<V�,dw:6���DJ�&���B�#�,��iM�Ƕ9��Z��̾yԠ�xtM#�������a�_7ˁ�	b(�ű�~����و�:�"f�VXܧׯ��!ȹ������ve:4M��%�[����k)��[u�a4�s���kqm��3��mծ�w��tp=�
�q>���@����1�9ړ�Y��ᮼ��
�	�v��]�o��Q*ymHMd�<s��D�Tص�ڗI�%U�M�Ӧ%�u�iz������خ "] :���<[E�}n)��C8NF��.�R��,�<۳��&��r���VA,4T�5��,WPb����9���[�����i!�w����{��5gr��u��^q=�U6zi͛�3&�=U0X���)�j����τ�1'��ōr���a�v�ˈy�k4��l-8$��]׮xA=t�ށ��#��Ӟ&+*�O��Y܈�ԫh謳��>�!5�s>=N�j ���	,���N9=Y�仫Y�4߽팵�#��M�5�l�n�B�Ս*��tʧ�tD����Rb�If��7�=yG;sF�5;Ӟ}q���[$�=��.�������qK�c�&Jx��xW�VS�9��s�,�� ĉ}�O�ٳ]>�Yfg�!���B�XL���@�ً=�܋V��lfm�݀;�.������3�S�w[���3b�r�����2�x3Qَ��]��v#\*H�qk���u��g�B:ܺ4������� V .j�-��w�C�Z{��]�U�MK�݅���U�z��gQJ-0>l�fu\l�(��:2��X�������5^0v=̊�j�6�q2�'��O�vgq�rX�oa�,飸)N����:�V��a�P��k�d��c�}p ����vΙ�]�����:�M���Z{y�^�VKt�vd�� �/Pp��;������o�?���={�t�Y�;o�bn��x�]�d1r�g .��/x�=]R���u3�v�`�i��p�>��b����4w$����v��g�
B����#3단��*�p��2=n�.v	���f�j"���t����v�6/Yɗ+�^#�#�a��K��0%!�����4b"����23��X�`�D�>��0�Q}��B�92�^���|��H�&�2�� 	���Y�=yu��G�����}����u�^���sZG�����(��o8��n����Z��6Q"����'~.�;��y�>��CHr/a���5���r�'��W��>$�7�P����6ߢR��}-�ܵ��K�E�F"���[S��
�4�``;��vy\��G��V��YP+�Z�}�ol򔓩�6��·���z{����]�qp=78q�A-U/��E�r8�/�a�'��p�AƐ�W.Mk�;1��MJ�`�6�5D���j�ZO&�[�ss]F�����6��Ƈ=�����2K2�����@�C9�q�Q�b��!I�\��nǰ#�hIn�W�G���*_��$X�Wġn�����_r��Ϯ�^�F�ZA\����e�;�YY�� FŴ@��v*�M�V����{�rǝ솱��:�\�Q���/n�Nr|n��S��zN}�Uj���t�k�!�X�	�\�I/�w�Q=�ݒv^'����L�::_a��s\�2
^:#�[Hnj�M_��V��+����<����>6�þ(vofA;�^XeΊ\�z�+\�L��3�n��U9�����᫴��_�X�h��V�X���:��'��x���ǧ�ث�_?p4=PK�5�;���t�����2@|���`o��u�u�U�B���b����s�:��[�LU{.n��x��.Y���
��o�c�鲻��kԾ{V��:�@c�P��0{w��,m���N�F.�B�q�| �K���_Ǽ�Ŀk��N=)FF�p/D��DUh�RAiyƽR�ȯR���MS��	03��"���q�!��]{����8��u�Қ����{��� ^���2>0���)�!=춷�k-� ��.o\k.V����X]v%���#�J��?tA�NR��B�V�sw��+]w5����K�����`_�3Ľ%�g��R�땅�̏	�aOn��aܠ�p��:]͸}xam�5{�=KL��Tϕ���|��f�}:�(O>ɇ�+���a�o'��F	����=�;S���Q�٭
��g>����A���9���t��<�d˜	�#I�.G�gJ{:#�L�8z���DV��WM�b�E����r���^{j���ח�"���y'�u�祍��hw]o��P�\�P�Y�x�g���X�\���+&�Y��\B�g!R%�c�X�^g���(m	�3�vT� ǨxG��	�|e���V����O����)������r��`�`4����]�=%Z�,Jخ����8V��S�9�N��Ly�]�W�p)n���9OùT9�$��(&c!,����BbR�E�IK��g�}�֛w�Q�Z�_Oyz���=O@�����*D�������v��v�#��1��m�gҵxi��s���Y�7^2"�0*��j�������~��y�����\M�X�6ѽ]�񲕨�-aś�`ît��֎�,&���!h^�����=C��Ih42i��\7n5�u�N�GGJ{y��p��o�J��snI�gc@�8fw
뼠6�ݗI|:�f�9Wt�J����*�K�Et��h���6�}*��L<�+�\��E��S�;j|�V�>f[(�P���x�E��A�Ej4wOVI}X�[C"K�E��*�'D]`���/��=���^s�zJ�r�U]ugb��M�yf�/�����On�n)+5�BU�ڴs$�uy�}�"V�*J�O���ΐU�- ��f��+O V��}ZI��<ʶ��z({-�Ԇ"�����:�!��Π��ź���@����7X���{$�)�Ec�mƵTڱ�h�v�xv�4.���t�6�o��G:��"-or�%YǌqW�>6�3��3;��2��L��Nh9FE*�ƞ )Q8�G3EE�_k�Л1WT�V%r[��6�_����������LoTB�m�����Y�z=�ׯ�B��L���ZΑ�nk�ȷ57v�:��Zlp�k��Y�<�ICv��5��1\Yh�;��H�����WB��:�
�Y�ֻH��:���G/�"�n:�r9'|1=�*bɰ�ЩH��t�P�ѫ��$�W��߲���ĪXm
�egaB$��:���y�����3�XرVQ��st��B��ι�C�m���v�t�,��)����v�5ڵw7��6n.����9��gK�/Wڮ���>�D�e�ޤ�RxKe�w����
��%u�F6Жܙ��ێ
�lb%�N��mC�� ��s�w%�󕌨��u�a�	��Y���{�*

��[(��E��Z����U��d�x+���:��퉆�qc{<��2���`b��Z�]��ҵ�a�M�-��w�M��;��x���|��;y�۸tқ��GsO>i�*"�&�v����oB���_��k˯�|ػG�w1N��Y�ݵ��d|Fl��P,R���n��J9i��|	*:b�ć�+K�n�;���!e=���a�Cf�Q�{��ΐ͂UM���CU�i� 즻j=g;��fsL_[�QW,����F�z8COx�jt��lW���:��ؗ����ˈ�&��:�Oi�(�,J�^m�k�2��8�������9đ�Rj�/�<�Ӝ�A8M�S&]�-�f��L��R�wW�w�bq���MY]�KVpp�NTcF�<;G�f�}����s��PY�rs�qƻV?��JÞB��S�ڿe5]u���X�2�V��vof.y���5��J�L�R�=G�7��IY���yo^�Ӓ���T�ď��(p_ZL���#�B�����\�z&�3��G��o��C�+��:$ի������!��V� 
V[b�(��R,VT�Y
�A`o
b-d�J["�iDD���k,-)��V*����
1m���mB�l%`[IP�²�XT�IU`��X"ե���T�ҭ(V�+R)R����QP���
�
�+V$U*,YQd��aYE�a�b��[B��"�U
�-�d�*%IX,��QIZ�ej��k XT�T"���)+%H�@X"�"b���Q���@m�"ֲ�V�,��IQeB�@XXV)�"��XT�

�ȱHVE�YYZŕ*E��U DR�R�6�d-��Z�%��Jŕ�H�J��J����
�,-�	X
��`�+X(�iEm�Vʐ�Y*�+ "B��
J�A�(�@����T��B�:%>��e�S�t5ڒ4"���ӞZ�:�mk�-���A��e`�X�����z��ew[:�2(�S�d�Iw]�{�6v�\d�%����aWvHSk��"xL	�=�-��6��C7�Ty��q�rb�M����wJ������c<9-Yc�p69��~�`�uҤ���faE��ӹx��:G���l��S��ژ}^�zrkR�ܿT^��^��bXϥY(��F���^�|�^��	�d/��+�L0�_8P�3 ҧ�� �Vz������[����}��(��}�����8NU��ʘ��� ��l}fC�N[�ʔ�dF�C[�L>��.u;#����'��֪=O~Q*y��!5:��b�Ǚ�_R��u��0`��.�
��	�V�~�"�wĢ]Q=�6��mY����	~R���;8�t�G�׻l���|`�����e���HЬ����,sX�@�"�'�TM����w9hj��HW��=�6zi�^��O�l^��H��Zܦw�5o$��pp���^g�c)�_�������0�*�������y@�MR�j�Ax�y�����مӫ�s�YmuL�k_��W��TW�`L�.U��K���t��)u�ZX�c]�ui��U�N�{�I^��nR}�P]م4��`����+�(�y90��Rk�XmD��ඟ$	�8\p�P���׫J��u�P:�5����qL�:�r,��HmeIgǫ�DF7�>9�����VvD�:�"I�e�~8._P�]m]d3�*g+ ������:�)�`��E{����u��"���C��u�Um�O���>�ז�����	�.�<�}��A�E�����<�q�A�`��p:O�vk�疄��G�<�������!�S�< ǽ�����+�_{�'�O����֠�Hyǆ�C������<&ط��+�	�<J��;��I���%�4��
jnԿk�G�Q��W�s̜��a#4@�ݳ�pΝh��\m�x���u����T%d�KfAW��@�Pp幘=��d�w+t��{.v�����ǖ��?ti.LK�~���RV=	Ӏ��=��+������`���4˄��701s�Êg����m���ϳ܆�g���l�>Fe��P�b�.�5�j�&m�����̸����bW|��o������)W���r�/�ڰ��%�Y���
�х�%��H�6�yU��h<{~�ڿ[��y�YK��>�'ƭ\���W[	���n�-`t-�Ỵ5���G,�ޭ\INn�ӢЧ��ya1����B�Cԅ��|��]WJ���x-�Npr��޽��f�����G[͉��rc����ɓ�^��q�����}\ �����q��d/Ox�(m�?)3��
��{$�{y�bђ��'+p���;J@Os���͵}�t�dhu^a ����m+o�X۵7�\�ִxCF�OUf�O�O|���ƔWS9{0ʛpV{&e,9��lK�`��n[���ǖ��+%�O��p��������sm˹^e�-�ܵ�VK�j�'�����z�f��ֱZ>g0��DU�L�̦�)]�i��F�e��T�z���~�����m��B�G(k<+��h�W��>�r���aq�^7M��fX�ȑ[#Mg�߈r��0��f���� A��)�V"/�P���Ĥ"D�W�/�)�Cˏ�����c���FOm3u*��%[�ptUZ���Hq�!��&�
�	Ŕ��dOE�[���Cw�u�D?��N}�
s �0�ӟG�p�u���%)��-�����s����h�'��=>+��qx:��x{>����h-p!����6�0$�����@ծ��o��d���]"mq�xJ�����a�8?��*�ފ��l��3.��H��P3�k�u�cc�V�V��x�i�zGv��0;m֢_+��D�����ݼ��8%Y���=�r��j�M� ^��
�y���wkWω����ȭvZǂ���[N�+�q���3�o�E��cҽ��Գ/|4�	�zB_����#����d���w���>�*���i���ͤ�P���$ �����m���y�=������N�̯xsA�5���d��" ��	������ZZ��D��K�� r.�2`ו��O�a��OU�D`�.z�eN^з�o�yy����ی^,k㚚���振
�r��6Y<��0��"Pq\E�&k~�]n�I�D��E\'�����W;*o���� ($r��	d�[��6�f�QY��Mk&&s*!�b����s'���iox��Dtď�ٮ
�S�,Q}�*x-��F;�����S��VV�o��������#�w��[Q�]�KO#���u�N�Ͻ���^,��f��)��ɳ�����ܵE�Υ����(?|�P�@�W	5���b��ћ������66��� �L2'��p���f��!�5�	�V����0�tH����}�WB�W	�����!Z���K[X�w=ZhP�z��)�t9�"-_Vs�2���>������s1��5x��h��h�4�[t����5��ݼ��W2�e\N�N���}��x�.�R�AY��� ��[6G��۔wn�.���Bk�6�I}�f�Γ���
�	�z]3��i|$��?R|d�u�+�]�@,-��=*��g}&����E�,�8����<sNS��U`�%}%�D���K,��V���I�0"P���j��<{Fa8\�V`��ǆ)pv{۞��m�LwDI��� �unCf)���n�ħ��͊��4�Ln'�u�g��@^tyT�T���~��)j�26�'��d��~t�J���1c����j���)��׍5�	�F�ȼ�C���u�ь���*��Z�M�m��}�U���\>3\xFN�W1�ܨ��vi�;5��	�����<>VR���}R����1R�k�Tf�:�-����N�&�(o�[^���ߵ�i��G���|k;�ͷ�_��G���	Y��p�/��Y�_8U[��iSόA��z��Ԫ7\�A7'k};�.�%�~�+��� 	|�*�p�UK�f���=�
�"`��ح���*g���V�{�X�e���J��6Oxũ��������$H��ӟN�'*�N�]�y!�,�n�we�M�x�l����3'@�l�=hU��Z���w���j���P�/�nH���5�N�^�\���$���Wt���wN���`����u���gP��Ȕ:��{am�I�v�X�^�����zR�ڟV`m«�$�S$}6r�;��riY�ʞߨv�*�#t6�ıK�v�Y���[E�n)���<*[����3#=/o���pkF�z�����=���S,֦��)�ʢS3*��4���`��<׹�^��_�z|�)Z�	hu	9�euM��re��7�A����4+���Cޅ�����l�*� E��������qL��Cai�.a�1JU0]�7Fkˊ�'Q~���0�������}v�;>�Lu�C�=��s(�'�`~�!��YGG��R���Y�/���L��GUc3��<�M�d=9W-h]���W��3���"J�����X�'kŻ�Z�m��b"���B���u�'�}�}e���yt�pp���V������E���]���Xߍ��@�# t�����y~��|t��W�|~���k7°�饞 ��zq�wQ�G��w+���AF��xk>�)�95Jݺ��"���W�	t��k������[�����{��<�u�a���C*��L�v����=H��R6	�/nї��l#N���R" �;Zn�m�[ߚ��܌��8���3ge�^R��9��]w�I�-.��{�T�5Ҋ���G=�8�et�P{£b��8��($%�#�&M4�����E�f�����_;ܴ��;�l��nn�@���0@��t{={�>̂��P��	q!��r�(O5+����o�lp97ܧ���l>���e�JJ�B|p�����%v= J��be��V��L�V<�:,�LL�k�34������aB�P�W�|�Ϯy��t/ʭ�F>!*+�Z+E��hon޾�s��*Q�yO~��c�J�g˕��<BjåC��,��wuJ��[o�.�m��h�sA���'��ڕ��]��>���Mvču/���H�)����5ϛm�^lK������˓!#Qu=5��<
�闽��\:z24:�eVS��'��݉͡@r���JB�p[�f���Lz|���Ӣ�;Os�a���(b�F�4�Vo�+�E���bo�п��d���b3�X.���A�.��~�%+Y�X���f�U*�f���/�K]�^|����"��J��4%o"8��xs�߆ު#�g#[2�3;aޱg����k�	ox�{ޯAWr�>v"0V	�(!0X��$�0Q;nО���^�^�i�k��$:��Z�>Z�J�ֲr�q��ݮ������3L�y�킲JN|k�{���X���]}Ƒ6/~�L��i�&.Jc�A*�:H�
X9�wo����WO�\�>������8�qXk�b�ڹ�X�]�ڝ�/%r��Q�ŭ��6ܽ�ay!M��b���w�yU/>��� ��A����yUbp=�����}j��f"�s�ә��
�ͮ+��=�tL�4���dB��@IV��誵WN���wp�kf�4�� ��^�6�˃ջ�6n��膓�k���0��5ꢵ��N�l��[؛���+|����OU+��3�}[�ǳ{2	�}�(DtV�,d���~��*��ӳ�sɵ�.G���p`dǢ}Yk�C����cҮ>p�GW��$#k�� ��R�'@�v�28��Y��r���<���ZFb����IP垠����9��1G7�&�^y��ksz���`b�o՝�m/��O�e}9�5}��߯|F���$m���3��1K5���X��Щ���C>|-�s����[�F.z�NW��/�>�:��j�Iu��W�Y~E�[�o��[��*UY��EQ�0���0��"|W r�4�!u�&cg���a�!��6rTvf���x�#=Wv���ؤU�|�d3��Ef}5��v�	���Q�e�]~A�ف��E4�,��s�b$�ټ���]ƨK�4�����;����nP�������}op
�wj�i�Z0,c������������T8��o0(8>y>Z����{���DMkK���#��af�9e��C沽|�/4��[ƭLT�|.��<B$?�	���
U�S�L���@C)�y��M�}�����&��Y�8}��T����=�H������=n��ќ����JU�����6��py>r)��]��^A�φ�����M�Ã(6E
��tY�{�u�u��ꗁ�ޮsu�v�.���S�d`�5�^g������� Ǉ�~�e0o��?�)%�yx{GNb����!���8���s>�`4�����R||�j�`�%j��J��7�f�o��;{9��&�"+[$h�k�<^��0u���ϻ�J\�T��V	,��K9��%	ޗ�4mǩޜUN��'X;�|f}�
��!'�����K�F��+w̒��2K�p�Uʻ׾�=�v�EF��UЕIaa��`cY���X�i���ED���g�V�|F�V{k�
�CÈ��y����[7ciM�ϻ�b���� �et��!,�ChvS�#W�Zb��{���� t��{�W�"��Ѯ=�涛
��.���v[��㘼
�X�t:��WTOX���p0�Χ�u���M�b��mÃ�%���q�Tjm.�����P�܇;��|��(�#%�̢����Q�0j��f�J¥��f�T���])G5V�8|�>�-A�h����L
�!�Kj8N�e�1U�Rq�	_u�vc��w����p¬m	1]Ca��}P��r���zO�o�����
��#]�]8�@��w���5Z�&#�K��R�OiWP�%�]���[��m<��б=��easlSY�יo޽=HV�E��%��Ė�O��	�/ m�;��؏���i7mg��5��ٜg��K/�!��Ǵ��[��aD�>�-Lt���S�c�[RY:�O��Dj�ݨ�W�i
os�3j]&pg�H��t�lW�Q.���ae�b�����\O�)�n��e��U<[.��M�\V��W/vz���F"k|DP�+�1VO3(z��|����C/\�kfv_
�y4v�\�i��+\66��ٙPOE<s�y:̞`x?���ۼײ"����{{ԭ;5U��E�e}��	^g�cL�%������!�꘥*�pu{7,VKE<�^�˭bn"�Yd��+:)��������P��N�ќ-L�.Z��y�#���iG��ڇq��.TD��YI�
��b��l3T�g%<I�@�*.���H\�ο<��*����c�v�Am�m���H&T趺d��Z�2����`�ۭ�&��Tx]ErXګ�fwa� ���#Z�����)᮫��q��x�s&Ʈa�����ŹĒ���78M#/&&݃|���`6�`̝��y����2Vf���Ӑ��;�е��z=*P=r�a�';� ɳ�V���C]���57�;˹�V�Z�Z$h��
���flց��.yf��W"�]h����e��­y0�B��M���9�}N��y]��O%��A�GH�3'iI�z2��hGŸ]���:�r�J�0�#�/Cޓ����JWV�hQ��]��4�֊�Kt�u$i���l��r�U0n'J�ۛۃ��L��s�-�Qc`�a˨D�AQ�L3L���W�#�9N�˽}(-�r윺�2��
�j�/b�:M�N��3B��oM�JlT��[w)�Y8�uZ��jϪ�� [閟d� m�)"쩜���eRʗI����e��t���mn�=̥f��ݭfKh��ܥ�'wZ������ܬa5#&�-{���$1��cu2���Vki8��@��}�;V����D)<��V������'۵p�f�.=��VH�(�f����}zZue60�'iKޜ&W`��z��
�e�v|r�F.�¹Y�k]�#z@�.}ɝC)Իyd�u:���f���їIbNm.�:�˰3u�fzهh_/y�����4:ƖY���Va����z�A!��1�p,��˷eټ���rc���F�]����]۱��N�����J��h[��9����J8��99t����m��+MV��h�k2��]�y�I�L�����.���k�j�QG�����/l���}"Z\�����u-B�ծ���{k��Xt������i��]��x�e�}�P՚�9��Uc��u�^nX�L�.|q'*G�鲓ϟ&-�UϹ�����&��\�o�����|*$*�e�<E�l�w�v�v
\��9�i�YR�#v���-�Yq�R��O����B>�t�ʵr��Z�%}z�u�R x�.�B��xF]>����YU�a��]1����F����|޼Ϋ����eZa��b&)rc,[�/3�y2�]�p�����*F�X�(sCF�;�����f�v�=��
�jԏ�ԑ�������\sh�Z�j�_:�mԩ'#w��<
Q�tYc��J˾��A�V�N�k�=Y��^��<W��]��u�㱙-8��4�y�je@Z�W.l��,��������s����6�;��;kkl��+(��AW@.��V�N��R�j�"X�x�`�k������)��q4Wqզ��N�3wA]���X�:��ud�ũ�V�'3R�N������mi��}vЭ��\�*:�s/�|2�S\ra
Z�����0��wl������ʓv.���>�*� ���ԅAa-���$�
��AeE TP��*�@�Um�	XB��E��++%eHT�)YKd�YR���i
�b�
ʄ�%JŨ%b�m*(*��*JŒ-�� ��JŢ�"T��TD
����V�IZ�k$�[Z��Y*��-�[J!YQHQXJŨVV@���i`VJʀ��!Y�6��*(J�eB�V*H,��"�I
��dX(V!YP�i*,+�j��IXPEP�Щ�TX) V�V���aU��R��Z�[b0+"��PRT
�ŕ�R,����*��d.\dR,̪@�iB�mJ�@ƪE
ER�����u����6������ٮeS)Ŕ�� ̦�\ȕČ��T}fX�B�K��8F���֩]ڒ�W6(�6���6�Hn���݂�տ��Y}��m�O�}e�-��pp��c��e)���٠8�����K�s�F@������S��E�p�@��c<��������^'��"֫�����r���x-2�~"�[�^X95j2�u��{��[�wg{2Z�Z`�)�]k^B:����k��z=�y�;-�����;��DA�*��̞´1+v�(�������p{̂����l8K���2Y\6��z3}5�9-w#۝�����WJ�����W0�v��UV�r���UGK�\�ͱ�(��w�����j��A/N;PӅ��y��x�*�P�W�|�Ϯ.���`_�[��k;s��Xٸ�WE�hD��R�9�N��ɶ�c��b2��:G�鏑/j��Lj���I�9���б�&>��b=#��o��E��:й�W�#]y�4:8�j�y"���q���gp����T�S8;�谈=5<����oj��ʙ��`�v4ZZ� ��t��D�1�K�� %��.kU�L�[����^]N՗�_s����,w	�����%�뷝(=�iާLiz.��G��47p):���%.YV5�;+�f]&��QfIW�e��|�7��]rpV_d����4��Vi��Sw�^���S���fA.�&1мtչx}o�um���X^�y�K�3�X.�����ͷ蔭g�,[L!dڡ��l�گv �-~W�g���Ռys}<,5��EX�f�*��k>JW/�ޢ�,�����/��I����fybu�e']�b#²e�
`��&���Ie	�z��g� ��wi���k1�$kF��;���/!�2�^��eJ�.�JO*�N���	mr�̭�6�<��c˽�uD�!z{����n�`�	^y��
�*J/��ѣZ��8j�R������޴���d\]�cx���6n�ħ���*�s%�0��n��7nNY�H�佯ݷ��+�A�Z���0�xmK�<=�_a���w����o����5�G��2%�z���Z�L������4>�+@[�T�Z0�&k�Ԇ�rD*�C�n{�n�}{��tԨ{=�:#����K�9��+Ӏi�T8,��t<m)��J<��㔳ϒ����mQ��P >���p����Ns��ʸ>ʹ��w�ٓ���D
7q��IY������:��M.��+��t�i�uŴ]���9.5��Χݚ�fVj�w�78ӌ����u�ĉ�Hw��;6QI���9�W�~���d������x���s&�]��5�@=�P�DNYվ����J������2��LV�W)���Qjq��\C�7�+yyu2��S=mn����:w��W��~G�Y�(!pX�y�Jl�M�R�9�+ ..dxN��h��N2�4p���ձ���h�htq4�����w}S Wt9��dd3O��0���0��vO
Zloj=[����X��m!(&�ƻ����L (�8pX.�ƕ<�~#>w�ͼ��A�樎	�	�q�8�cػ�2=�gp�|%4P��IvE-<L��t�ź��dɔ_���ܔ��֩Rx1vh����7�L��c9]JD��	���°Pl�p^%�;�I��4%�����M�>y���N�VM��28��K���na��L��7�1V ����x�Yy�^w��m���0Y�1`H>(w!�t�g�������I���j�`�%l�������O}x�����gUՏ]�Ep�f#�<ԧ�����^�1)�$�.
>�3 ��׿r�ݘpe#a���S]�
�W'e��H֔�V,�I�Qqp��颃��W[���N�IV�1^��uЁkge�Ɨ+��Qg(3�����J?��uoK�t�w�n���ɖ��{zu��wi��`���s����wֶ���NJ$NMJ$�}�<��u�}�v��W�=�w����r����LX��o���y,vQѬ�M�2Lp�QP�*�����4h{ⶽW�W���&���Ɨ�Ba�%�i��1�9o�X��[[�Ҥ�n����9� �_��&y�;�r�/Tϻ|t�v���q��߱Wwt��o�/b|��^��eoZ�����3��U���ɾCt�v����-�n�o�:�	���Ð�lԑ���eX��튜F�-N�[S�ü{�g?
�~x,MVoM�;�iz�g�9�%ɉmY62��f=�u�7�>�Wx�aw�By���=9�jGo�K"��Q��~i�ń�g�
�ah���=),�'G���紼 u��7G�0�
5�J��h�8m���}�)[�i���pRd5�ح5^&C�}j�}f��(�<��&�B��Y���=��u�:��j���Ŭd4��u���@�]+�t���'<}>Eh�ls�n�V��Os�f�â^�>0��3��j�y��y�<�g����f����]C����Y�OZ�j�c@�Ji��b����`�h��\ٳ�)8�{0�B�_y����"�瞲�A�1$�+7*���z��	�YS�����p��8Βwv�h�lL������=s�C��r�IIP%v��bT5��n�(b�ǃ�v��'rb�����cf\��sŜ�^�-��D�po�g��پc&Xw���ކ5��zЗ�h`�@pX�]8s��}O�=�z)�_����6�\��J�����{{rt�{���`b}�W�$b�Y>�b��|)�·�5Mx3��A��`hkח��;�wReqX9�`��v�ǫ�&τМpO���$��f���hU��Jx3���{���e�S�]Mg��$��`xϼ�g�Y�H.�Px�x;Ȓ�L&����G��oOx��Q�t�����n����g�� }E���[ FH������8C��3^g�e��>)�ƛ��k���}�׳{Ր�e���@�@���r����B����!�&�j�,7��˼����;�^��}-�r�J�t�,.����rCF�l��hwt ����1Ӧ�b8<��GV�/.�ʻ�����,}�x-���8-���P@���1p�sؠu7�NgZ�c^Ai�Z4i�d��=V��`Z�!�y sۓ.nu�����i`��s��� ��)q���2�R�Hb�1_ �E�6��$]g;����޻긔��$[w�`�}�GF�V����̕z:�Yo�Z�9D05!ɀ,�X�U)�y�ޢ�f���(��v�qEǳ����=Xޚ���4�B/O���x�?uυ�#0����(�m�oԖ�����ה��PoU�N	�P�9	ɶ�Duz�}"��J3�����j=�~$.�N�4���������աz�����%=��7�N�QO!�+��|U�pL�\�F�B��Gz����ߩ�x�]N��&m��UV�2s��X��az����#���ʷO�^�)鮏Z]v�\����l�&�X	dm�� �&��奻�e�ࣺ�MO756z�	_W8$�w�T9O��Ï�r�jȫ��W���g��Xx����ͷ蔭�J&�c�8���?=��ǝ~����s�ɗ0����E_;4�@[���������925�S|uX�+ktȱJ~��Ί�( &��d��
%}nО�t�rͫ<����}�[��eWo���b���x��}��2��7��v*�E��՗a �D�{��?f��|�Xp�<�d*��+1)�N�Fl/��t$�=Q�2�y��Ċ$��L�7F�E�_Y�]�ՊJ|�L���о�Awi.�^�eI]J�~.�9עsuIh���-,n�]�ǵ��p��5I��ڴV�嘖k��NP�[�
�>�qG)�Q�F�*Z-"l�UΏ�ܭ��+b�ilV[�s9tńs\�9��-N�}��BT"��f5�xe\\]��C���#>�i9��>qAO|{eTI�į''�<��6��G�ZC`h�l���sr��ofA<��e𧤵�mc���|���m�����d''^ä�x���c��q�?Ki�V=*����2�㹷�]p��\�zݷo��D���I�
�w4���4z�_#�y^�t�Y�	|]�&xY㾝�^�<{���LVW��N �:�ī7��zD�s��ɪW�YO�n^fR�g��A��ޒM�}{��L�2�/B�CWa��������h��ѕ�{BMh���M�"�6��>ͫ�C~�����!=e�i
_Uʺ^��a>}frn���\��̇W[d+���o4:c�@�ss�*�Z=e��P��ݡ,�H�lT�d3���M�Z���=�)��N���{٘kBgυ���i+��i����Xҧ��ƶ׼�l��;���{���A	U5<ѓ-3�je�)ʞ�u�(x�a�,AKt>�~Ж�]V��>V<��	��x�fp��@;����5B9j���V�7{v���:�iY��/p�����u,�^��NY�o�L�Q�����E�<wt�*޸�Y�꽾��n�Mo\Yq�ZB�쮵V�(s�I�J�WGR�NLN봫sI��y��%�[�K�`�s���p�=&�z�C(J�hP���;����rvw��F��},^��r̮�d`�z��K�඙���!�#>��:e����v���pFHh���@���V\1bA�C��Hge0#�HT!���h��y֣��b����;Lw��c��H�+at��Q����8�^�S�I��Fi��v�smGy�;w�Щ�g��EU�����~��1X�����)�=����⻫�|�ѐ{����<�$��h1JE8�7��8���L>�@^tyT����'�z�;����R<z��=ȡ�c !�*�0���L��v���,^��`��0&<ْ��˛7��w!��[s
eT�E·�Tr�L«Ճ�<4|��a}��p�P�+4�{2|T�ӢV�٩�x��ʜs�cN���v�{�#a�>Z�B�#��S��ɭJr����uq����jo�6����V�c.�3��i+ �ap��!޲�9�_8U���ju�lKo��W����W�<"/N�|���:�Тs^<<L�Ο�	���^��X��aY�Η��ɻcD�Zb��g>���$�:�]�N��S�*�pn��]k}����[υ�����Uq�%8IV�Ew]z���p�2�jL���{��+T�:�E��`|bKG�?0������D�
�D�z����<� �Ԃ�]]��w�5�l���V���!�/�S4z��C�E����5O{�wA-��G�E��8��b�3e�gD-#< Eh�Q.���z\�،�tS2t�i.湜{��o�߅]��d.���z����5��E�[J�gnvKS�d���B�Bc/,Xֱr2�w<z^�}R�HW�Ow͞�sj����]lJy,h�1�=˱*Ӓl,���ۂ귉�����,8Voy��E0k�H~�M{7��}�o�G�}:C��e�N�^�"7��7�\+QuB�d�����c��GG�v]��|YCjܼ���w��z}�!���GFDr���<I*
�P||6�,���cb�1Sh�&4�+��'�09WlV�f��A˯$w�%�
�}Y얟�Y���bW�{,y&�ދwyW>��Ƿ'�Jx���0��d	q��� �hu�U���!ö�e��k�׏M�Y�9m����ڊ�ڳ�C*sW��|D�BF�>Jȋneu��M���a Wvu*-��nh`'%�Z�t��ӝ���� ���1��բZi�]���VV�mAT�gS�݌�o(:�H�u,p���'NU�|.���OZ�,����ù[EkPQ��xk!�zLvh.9�����^���DY]~J�ˀ�|�|)�n`uzy�=`�R�&O�s�W��mz^ftkT�����r�A81�]���-�'�p�]O/	�ߨmSŢ�S去��u�`�%�Ч0#���}�֢F��3:�;~�����!����	g��~�ʮB��@#�,�=$�����@J-�e=����`�
��/�d��t+E.$Z>�^z���&�g�=��^v,�%V�\D���K�];)�m���F/������҈��2��>|��ַ)`~��|Rb�,2�(=��7�	�j/��R��I���g��g�yu>xwU�*i�H��`@n�����[����l�oN&[#��W��߼��5�,<Oo�t>�q�n4P�}d!*xX�va�j�A�M=�S���/�֏�e�qt2�k�ov�廘f��V�!����DЕ��'Gi����*�GF�����$���$ I?�@�$���$ I,	!I�xB����$��H@��B���$�	'� IO��$����$�	!I`IO$	!I�P$�	'��$ I?���$��$�	'��$ I?�	!I�	!I���e5������!�?���}������   P@
Q@P*��
 (�)$�DDU)Q($BQP*B]�����9�*��TI%���@U�RB*�)R@ݜ$prP���[d���WcSj�nݠnt:��*�r��wT��J��Aܱ]ks��.��m桻;���\�ԅ�����48��:T�H%V h  l    2   ���mէwf���M�W05R
Rͫ��5 �"� ��t�fJ���m����V�2�j+X0*�U �;Y�P�viWbٰaIm�[ej��*H�%�uT�25Z)UZ[*�հ�+1
IZ�,T�J\ !�����X��A[j%���� L�"�)#p1P�ɦ�̤QU��٤�h�V�6��R%
�. ��-�VcFkY��Y�Kk`i�Y��(ъ��Z����Hm���e�dkmZ��M8    &2R���h�M�h��"�0IJRP�4`� �b �0�挘� ���F	� �"��!�R�i40�hh�	��d@挘� ���F	� ���IA�Hъ���LLM����_������y�r�[m~��ƶ�x����QEUP����g��PUG�?��EP�EUUEx4UUT]U3����?��kiT�!U��
��"�*�*����UJ��P�4QAUTi����?���?/��~���PUP���S��l3\bO��vO�A�A���_�����d����f^ede�X�:�b͢�[(+�ֻy^JF��GM�W��V��dRj�H�Zc�n���PKG``�d��j����\d�W�ڬ#cU��+���r�b����Hl�v�W��j�aZL��V'�P��	��H�����DwZ��4�	YK)IN�44;[�e+-Xt�*\�,S
��n��a�bE�����)�y�P4�D����l�0(�f�[z//*^̥�ڭ��R��?�����y�ï���ʊD\o�LS�R��ܚ���Kt	�:���#V܌n͡V��L)�Jd;xv���h��)��2���9��l���D,�\���m��3�#Kg7u��sH�H:z����n��z��-nS��\U��@�k��� 7�K9��-�Q.���]r��'t�qP��X�BAr�̆풅���V9gM��r���-]n#h%n�YP�(�//m!@\�(�sv�ne,��jmM��7뭲-M{g+m@p��	�@"����*����e9V�赪� e�j����1V��X��м��F��U�ۊ��Zǩ��O6^����P�Y��n�IV�"�ܖ�a�lLFRodg�go�B�%ʗ���ܻ��V�s^i�J���*!6��fe����gj���w"ٸ���x������\Ţ�m�tf��Y:�N �0\T*֦�e��0��z1���fl�Qdy�X���u��U��Wi"�[��J6kP6p,g�Mɂ��&*�+j˗%� z�0���O%$�y����F�k3R��{��DkL��/2�I�(^��Lre^�nn`��q�������,�ަ3���Fk�f١�l��xÎ�j�I��D�����\`1AX��H�^��ɛ�7��B�]���8�&�xJ�YfK�b�Y7@f��,��M`j����9��`cC\7DX�4!5
��;�lЗ�b��rU`�0�bI4lj\ʎ�ې^G�n*�wܾ��8 G>Y���l�J����̈V�	�W��c,5bYX�ea��6^�
�HZZ�C�[zdn��[ـ�E[��Me����e+���F]*yfF�lY.j�q�jԬ�1�GffFs���Yj���h35b�L""r6h:u0*ښ����i�yksrJh����m���'�򡭫ـ!y�'7c��ܼ0�x�ci���t"�����&�����? j���Ȉ��8�I�)���0�7���*�f���0���>�*�kn�D3�{�۾��4��-�Mflv^�ϲ՗0	I�M6�۲�j�v���+77������tmW�@�-�>���%��"�)q�Z#h�y��f�5�&Җ0�8�Nc�ug3��,�h��FlqF���2�Y�"�j;�wSۍ6hQ�
z���ؗ�3hKr�1c�sK5Q	V�Պ��ܱ�eJ��,��:�]�ZS.��hn<�=�zΜ�*^*�,Ů�W��j���#e��٢jm�<���:���b�f��+XU�I
�sR�YlfK�z1J6�+�m�a��he�{`Ѻ����Y��#s1'N�hU�k�$�
�Q���< io�V����}ץQN�]3i��-�by[��2Q�P�{���g)�A-i�3E�G(Va���6��34�VJ
1k�"ĚZ�ە0YQ�i�am۩�iCBFNm�,੉D�[��ǖ/2�)��&Sb7D0���3	{q3��72f�4*^��I�c�;����<N��;����wO���w���d��rTE-�"��h�CDss2$z4|�X]���W戰���P�bS��K�u���_K˽yH"��$�����*��T�`�jè��
��ܥ����I��G���X�����m�ݬ�,�1bX���(f����G��)���yWR�ڹ��T�^T�Yu*Fk8իӊ�_=���*��� �q.���4��vۀ���Tn�v� �Ҵ��^;ɮ;-�ܳ�KV�L���7c�i�2Q+r�^-I��wi��#�b���cX���(H3����ěЍ	 ���؁�{7@~f?���b�߱C��Jd�)Օ������A� 
^�ݔ.����ohi�E�F�S*��죊��C4AJR�1j�5;�VF����,�H�Eۀ;�IϞ�����[U�+�6��at�k_h�L��	/��E%�[E�(�͸��f�dH %�BP����O��Pgэt+r� �i�Z�;#-ʛ���+t&��^�S᝸4�Ƶ�����Y[Rl�zcʻ�z]^�%-������$ݺ@Y��ۢ`�MDH-8m�ydM���Q�#M�f�c�Yj���9x��5h�έj�٥��e�F��rQ�)VMb���n7@%�T�9����N�Y������H���O�F��@Vf����f��]��6-��ެmXD�;�W�aآ�w���ú�ݼ�!�A���M��6�c��ee�m����)�L׸��3��ܛxE婛�F�n��B�gWi:Y�e2�⻏<[W�:�4l�j��C��T�][�� Ő�N�e*izn4�0���n)so�[��
V��wܝvQ�8�(��ł�U�A��3v!�1�)ej�S��0��7a��Xf#ZrV�m㵆�r���L@���nn�[34*Z��7��ߋ_�?`co�q4%'�>�]ć��ϳ�Z�~��9��;w� z��r.� T-c�%.2C�$�G�����2���$P���xw�����z�C:��oha3:�3w�Zhw��u��t�on��Ɲq�]͎d��
}�CUM��+s8�t�y�6��b�PQ���GXk��v�*��_1sM3�/
��[�Ɂ�f��tI�}W�4SP�{���6ʮZn�T-<��-JE�J>����u}#w,p=��N\�3/u���3֕���WK�_f(�1�/��q�}�3�n�2i}enAw*HF��x�7r��5Cv�m��Y�$7]�bڼ�«q<�FMO�V���@^�Y�n�^M�u�U�SP�|���t�Tx�]&M��=5�p�kp���H�A��ӱX�`�̚���i-7�0���&L�8�l�v�x�I�8ve7�ë:,�N9o�=k�`f�:���>l�m	gs�'ΖV�Z�jҪe��r�1W)xX�y]��]�ݽ_[�8�R����79�b�B����Tէ��zk;�G3���_	˷%��S.f� ��t濾7pS�r=RE�;��5�[%M�dӹ�tN7zN��2k�N��.�{n��RՓ�n#Z#�m̙�!����gK�Z�>��\���!�
Ē�d+�T���g&�C�ʂ:�C-ݹ)��m	g���V3���R��Ƶ����`�e�u}{�������#y��s4��\R�(���d��7kc"��BlJ��q9ۗ����`UF�
����π�M�s+I����Ye'�%��������<�ȷ7Y:�:k��vR�^�Ȫa�nE۰�@�;\��6�L��۝3�!�]w$x��a.�mK�WG	�o��{�wu��؀	�&��J���t��u��Y��>��R�MK �`�������d�����s�J,ݮN�F7Y��xohGUʋ��Zܵ����m�{B���1�jY9nk��[iwshc]��J���r�R�ӓd��^��2����S�OY(�f�z��Պ
����u�<GoG�V��c^��]܂��)&�c�(v��cu�,ͭM��[�wga2*�$^+���=%�3t�i�	��C�M�o��{�)��K�J�����㽴�ڴ�lੇX*r�ବ�l�K.�c�Jd��fX�45��(-�c4оS�s�m�{o8f��Az������e�ޔ�'pԆt[������.g�U�fo����}��� m)�vVv0,x$�����\�ڟc�[F�Uf[�����e�@����EQ>����F�I�v�G�XDWH<5��'����9|��C�3�0���:<iv�����_76G��R��plʲ$��i���k8�V��j�M�^m�-_U��������x2n�cj��¸���b'��O�
�Yj�4I���l(�;�:��Z�j�4�v!�Z66����i�+�f	2�Z��P����.�3q���[m���z6�*�nʳ���|-��[�Gl2_)dU�i��uJ۳ҽOV�g~b�<I���"�ǘBcw��#5��vH��k%�o�q��Qs�
�p�r��J��Ѯ���r:�2˰����{�)E�0az�"�̭ ��^��:�(�[�K֝fM�Ďn� dǑ�n5Z�κ�+p��OR�Qb�gٶ[*��J�ص.��v����tN�3hG���Q�1I�k��&�=�z���ЕdU��d�k�����Q���(�f-<HS�'[{�F���Y))��mwXcEJ�j9����d�n]���})Dv�"e��Sa��iخ�%<�w���^_UݷVtf&�@C֎�8�{ō�I�g\���
P�U��b�p�7Yn����=��`O�H�m���
4d)��ud��K�Y���c�������[:��5i��7��:��)������o�81�S�ߧ7�݊}�ծkùΊ����:����v�Vf.�P�S�*� �֫.f�]��Í�Z�G�pcU���a�؍oơ�]�l����7���y�E����A�m�[-o$�B"�J�2����nm3��۹u���l��b\�VޜY/���^�uI]ǫ�N��0N�%�3�S�"&~عÃ7�c�����vm�����S�Q�uN��k�[���:�����̉��l�M�:C`H�8��p;�\YbN{B}|��2�W������۝@N]/�=�%r����k.��Q[�9��JⱭsض9iD�KR��+����ӌ7�T�3�Ώ.GݼD�KF�驨��Ýxy�[ͬ��y�|ƳQ/L�;�Vv�9:f�(��L��	fgfx�����G�/EB/0L��2c[�.
p�9�sU�������<3/k%�W��!��pW-�.�FX��i���X�NEn�	C:��)�sG*��&�:��;BrX�g+��>���a>RA�$��9�&l���Y��M�GR�'��I&�I$�I$�I$�I$�I$�$�I.I$��z@�S/���ݔw����Ҡ �f�aGj�25�w+���p]=m�I�Nˏ�wJY�5.�*c��t�d:�{�����,��m�y��)P��ý��RE���s6��lG�z��ۘ�$j��.1o8w��Ij�ovn��u��{u����a����2�WI�Tb�nv,����o�°n�w9]���?���g�Ө��T{�肪��}B{7̕AUUT}k�A�j�~a���*���?G>�����κ>�p�p6����.��]�
��ea�s)uXQjۮ�������#q^�{ՙPp�}-�.2�38B�_e��'[J�A����x[lu5蕵��,��u�<�h��3~��9d=B�Wm�X���+۳ƻ��v9��sm��!�t�]�Sj��9�t*ڔ(F���!S�)�>�3�HwU�vd��0t#`T�lֺ� }���˄!h��V�{\Ai��Q5q���/�u,8ũ��݌�	h����Jc�ru3 ���r��z/fNуfS����G4��k-�]L��FS��=��9Z�I����.
W:=�4E�cks�$�%*�C:�� �n��R�0(��*��W|�nl�W�{yCc1���n�÷d�wYT��_��՛�*uX�E�=W��0s���@���v�r�6r9�Vns-80�lF�մ.j����C 	�2��v6K�2S�,\!c�ńɽ=}��� �0�ݣ6钶̎�z�c���B�̤�{s��<��9�]�}@:0��ZoTU]*�'gS4V��$�+n�(-'F*�6�.���Y�MӺyu d����df�	G�ט�B��_}cz�����p4���\;�F*�ˡ}nG��m�&�A2.�]�n�.l��!�$zE��rX�Ϲv��N�/�]���7[�ĸJ��+6�x��.b���m�˽r���hK�X33mGt`B��v����j�:4&'[�pd�5] `��a�Z�A�5D�`�3�pX���	�;���S�:䨂�`��y�ʫ�0V��#�2V�t�P&��;�g]=�ѧלG%�~�X��te�����-�W>�N���f] �$��CX��=��݃f���7�FSY��nG%�`^1s�ٵ�\Vn�ξ�����nY�A����Kn��f�N�W[�|v�"�s�����4�C�E�V�!�����}Ţb�]a!H7�N4­��J}un#��b����om�t6x�	��XN��ne^L��&[����$a��/s���Ok6�hYs]����m�D�N����y9�����Na��{Q9c+�Ѻ�[ege��N�H@n��j�JqУ�Jb�0��uf�r��3�W[��I��Kհ�1�z1�S�K5V+�]��}�;�����K	Q���R�,�ؓ��Y�����}��k�I�WK#�E�H��a����T�WdW,�G�U�`ӵ&��y;�ej)����F_�w�s�$��L�(wF�qn)�.�dx��/lZ��g:*��Ր�P���ZH�[jmF��au����GKY
���nY���1	O>Yw*�9ER���Jgu�+��bv�x�;df7(��hҳь��L�*�]G��Oa%�E��k��+��Y�p^I�����q_r�d�c��`j����}i*E�ݢ'NVCڶ+Q{h�������A��Pf'M�Y�F�ً�cc��3)�9x"�C����h�@�����Ѝ�&�|��*B�3� ���׆�f�6gbd�������x՜6eOL�Ĉ��g�/�efn�LټS��ڵC4T�l��oz��9w�Ն+(+M���V5��si���6�[���e�˙��^"����]��;|2����Vܰ:��b��P���	�Ʀ}��`Uw>G���V@74��M���p�m�.n
�oĎ��vd6���z�ԙx:õ���8α���ɝإ�!��%�f�ʀ��9&E�d]��Vk����{��l�������[�s��b��;�>�uEg�5&S2
�0V�+0�J��jfJ˵��2�����o���O4d���u1X�_�2�ڸeu\��Q�B1��U�� ��f,WXW��Nd;YV��gV���w�Yki�x��v:�#d��痺�]W�Jf��Js����t�6��\r�gk7hT�frT.��[2��$��Ԍm[��⭗��P_����7&�d�Z�Wa�#ɝ�j��t�����f��b:�`b�)]�/���N����,'�d����_ǩt�-���$� �-V%���T���}8M��B=�k2�ԝ�f����Tqŷ0��h�m'/>�52,ǻݫ]���[>W2�5�Ji3w��c.������*�g���xrMc��o ����
��t��xX��+��ϧL�e���L�(޾��SJg���iɔ��z9-��b���T�ܺ�棛��Q��
�Wt+�S�y�%�ɝم�Ig�ɼ�M� ������w]A��j_4�Bu�Gf������x���\��+�J��n>��F�"h=d�$�[��dr�pꫠ}yc��7��EX*�t����C�0+iA�96uݭ����qMsg.K�v3�Dޜ3jTHF���+4�͛Ⱥ�p�!��ڟ,T�Y�c����3.����Wsܾ���,RLy�\"�sua�ve�হ7P������	�7��t�k������Um���h����E�*�K�u؃)*�[�Ь;�]$����-0��)f��JG�;L�h�A)�� ���:5e�鵕*xvVf����6N����o:et[f_Y�dp��5a�Ew�
���a4~mEgj� ��3�ٍpڻ2�y��=N�YDmx��)��������k刻
��j��Pg�~�s��o�������}�[�t/���d����@�ѕ��u�\�No����������9���_���Ҷ��&w6�wyfgJuz��ܛ�ŉGF������B���;�g-��9X��t��3�� T��_l�cT{��;2��7;���-;R�>�zQ7iK��#�Z�9dS~e��Q�8;r�.��+�+DbtV���I��ˍ���,�������f��"����/"UԇΝ�N��aJ4PMB�:�r�Nh۲��*D3�E|�ӎ��﷜k��|�1�A= �(جEZ�׮�J������[�X9n��JȵR0V� �UX�V�IBg�`�V���BT#��8���e-����R6��H�Y �((�5w.����F��$"QQj*$KAcKDh�*5RH҂��h܈���
-(�T�\"�#Q#G��{�>k��y=��sF�n���t�w�EA,W���$�f���_�����?��)~�1�7;ψ���Q�Yr�S�\�>��p:�KHXہ,X���O��]o���gF��^���_=�pٺ�2=<�y�W�>CvwN
��<]�T0�_^E�]�Eԣ[��<��Ĉ��eh<�����V'ۚY5�bC��Z���8��A?z��#��^�������Q��PS)��;�uqs��+�kV��}X�mݪ)9�*s�K|h�����ܟ(�w���R��Hv���u{�nLpEM���� �R�H�������;-g	n�.q �3e���+N�z�n�gy7�^e�7g0�l�\�q2�lo�,!Q/,K{_�u$v�;\p�9p����:�q���w93�a�CP~&F(��5��&���kG��Ѭ����]]�;N���HZb�p���G�̻7ݝ�Ԍ �����]��J��UV0�k�N�y�B��5�g���5�=+:���Ϡ��*��Jm{��y�N����t�ާ�����l�ZN�W���{��������A�����f�3�Z��:�SG6�I�+�:��nT\�aj�.�e�ʉ5�ݯxjICň�[>Z�`��!��]0d�o�xAZ@�n�T'`��LM��=f���{x��n�*/N�W,�{�u��D�S���:�wW}�������-1���c�+q9��f�w	r�B���-�F�t�/�@y�|t����M���Q�,'4���(W��6b���Vsʝ�	+,�f&�Z}ܴ�$"v�#`3�ॱ��J�r;3�6�䎵�7��{V�j�[�.���<鯱���g�@xùK*����B����8�n�Y�P�QQޟm�g7]ݰ1Wl��,��Uү�j�k��'X4����{gZ����~�����pՊ�Amңb�z�z�ݧ���V���h��U���by슼/���G����=�V
C�`A	7���o1�^V	�k2�C����8wr[ۛ�}+�[�� NC_Z�x3x�>&�������ϱ^�|���b��m�}��޻���.��Q���]X�D�7=4�ľcs\ϯ��m=�u`gC�_:.�R�
#OZ[�~�F��8��洃���nS|7����,�#Qf���.��dǶ}�[{����і�G�!����55T/c1{Q�5�O*G�B�;|��:�n�V,o5]��h��(����Pp�W[E�n�m�}�M��^��'��Z����}�V��U�/�տw�������S)�g�Zm���x�����\7ÖCp��i�V�ڙ��Nc�繛N��ӄ+�2�#f:|r�v�b�C���za�]X+A�a���1���� Ե�{z��T\��z�]���V��@�q��*q��DT}@R�,R�*����/�{���W�:�50�h�=Y��N3)��]{�fW�&����N�CY���ד>~�+㙝2�8�QQ���S�|���Ϸ�C�M�Tw���zW}X���@�K5Io"@�X�V���=>.#�d����S�L��u]u��s��˦�jjڬ�V]�l<Ng����u���a��3*�:=�b�e��9�{�3Nb�i_���D􉎞u�UoZ�����4�ۜ���e�mϳ����U7�a��kY��2��O5gK$��c���8kmr�z��[v���{��ǻ�t���#Z�,˶>k-fBe��1��z���!�@�!�L����>�P�%u��Mm�zy�C~���g��zS'������8�[���I��2o=Y�胗n�>�fȗ`�\J=��!���6�_pC�b���[^�Foi˟>�ᒲ�^�Tl�Y�z>#�
����Ƶ9�`ļ���j�}�xA�1_`@���5����ފC��ME��>�V�}�J��P+yb�����b��]B�ū��O�Z*m5d��f�S�ǚ�;�y���Νp�+�>a�m�\(��U���'v���6���,Kj>k����r�k�﷜��ۧ
���1+�y^�s����q��Vs�㧉�����5����g�Im]����t<��)k�QF�d䈔S����t��a�]:�'���p�!�,�Q�Hr�hk�CJo����O�C�S���6����]TH.��_Ӯ��U���e��w.��Z1/0-��!��Z�y��ws��!��e<�Ic����������C���>c�,V�6��>��4T�e5�q6�6�r���3r��wڣ�.�8>N��\�����R?.ޛ���C�+�>����5�Uy�ꧯ��L�I������X����N�{8k_7e�rײ}�vf,W�6�M.�&�[.2o��f�Kr޿nM��]���:۱r�m��v�௚���e�e���8��J�����얨����^s�F�A2��}�sR,t�]�}���P�t.K�yf9�`h�4���ο��%���׬�g��)��M��!o��MB��ƴ���4��O5�ŋ}�]���%���m���mjJÖݡm����;�;�gA��se�w��嬴e4��P�7���}�l��B���N;��NW��T�����ؖ��u1���aI��҄X+F
˺΋�\�L[�N����Y��{��ob�}��+��&�W����A�w�z�M��)V�U{p$J��Eor��~�h��8���=����ea���['\ɕ��B�4Mm���r�wn�J�c�Z�qfezo���l��Vؙ���E��z��RJ�6�A{�&�F��f[է_�p�5!@�.���"�4�p8iZ)}�17!twV�m%����v`�]Ɛpʎ���v�@�5�iTEj��&�YBTf�F��^��	��nnk/8�;�;�W˖����G����Y��q�T�{�s�+��î�Z�ѱ�r�/��P�գ��:��|�O��s�آN��3�*�14V�138<�r�tok����<�8���w6�ө�.#}�ro�q��u)d)w�L_R���5��Ly��aX�A�Q9�)	�IS�&P���w��	�݇fc�4N��ɱ��������G��h�r���R͑7�feu�n�����=�ot�9��#d�5#�묉�ʈ��-�9�(�R��Ftᔝ���۲�c��P����_���tQ�}Bi��g>|��7���8 2�W7�z]䏻D�n�0�c���1�c;{��9������Ɏ��6��R$ij��)��H�K@�$�"Q&b�A����$Q���0�Q"A�ظ`�%E{�`��X�V6�"[L�RB�ոL�])Y��R"���KQZ�4��p ��*�(�[e���-��UH����h[T�*+K��(��+)V\����[�Q�Ab0�k2�"���ăNd�׾����k[�s�����v�f�v��m�O�}$R�v��[�}ĭ����Y�,��Գ��WFyǜ�{��q�����̧�zΧ��>y����i�֮���m�m��Rze=5eܽυ{g�+j2��N����3�-�xx>7vvD�s�j#f;½�����S��ڼH�2��:bV�gVݲӽצMr���$O!in�����''\�Me���{-�k�U�m+ӗR�e�p�Z��/��r궘x������\ ˳�����szέ�kp�W馵�Xk#ԃ��쫁A��� 2�e.v��_���sS�Ib���_s��ȇ��ei���� jtT�U_P�
k�����8RWL U�����n���L+~!o�B�*�^]�ǹ�6Og�ᷩ92�gң]t�u�{�hɊ�y�j9bk���a�ʇ%NνM�g<�ļig_��?�V�"�� �����'f���}�����ە~����t�8i$����&�t��Q>f��K����
�II��q�M��g��ݝܬ�Tx�ZZO����h�t֟���4:��)T��<a��5s��a�O^����U���=CQ��i�y��9g(_�e�e�6~�gMϳ}�y^W�ݨ�cZ1��}(�/s�'�\�/zYL����X�瞿�ut*�����U*+D���o�s�a�9uԴ�R�G�u���}Ƹo����z��6�§󆱈a�Y���{��д��4y�d�4&��a�ƭ��z��������S����/F>���䬕�y�Ýʞ�䉞�q���wZx�����U�+.A
R����{vn^x��7��e4�2�hi�]��:��o;�Lnvֺr�rg%e�ә[t���{�{or�f�'�fV���lv�'n�#H���$����<RG2s��a�Q���p�lmV���|�N�C�Y�D�p�W9J�7��f;�[���Un�J����x��u�����M^��S���q���誅>��)���\�,�^똋G7go�2�QJ_Ԯ�u�ӆ��{y0���9��o�*|f#���3W�\ab%,ӎ��ny�5f4`Kk�i�:��ӓ^y�i��Q�1UɚF��P��z�]���\���8k���5�޽k��䛆q�=�{Y�s[v��IĞ����;�2��W�w��oP�Z�6�msY�y�o���}�+z�^<kMaˇ�[�Ž��M�tlZ6p�r���:��g�G�Wn�͋��u����&*a�ʡ�A�XN�(������
b?Q��\_��L	�5��fCM���s]�u��a�R�ww
c��Ϥ�L	�G%�7K���z9Ir�!���w��~���Z����u���8��a)2�z���W�-���x�ސ�V��Cr�׹��/��n����3a��mZaN�ٔ�r�93���{�[��x�������n��R���&��G����+�����������l��|��S��ǎ<k�Y�1{�=�o=��\$or$Ԭjy/�~�쨄�?�Ԛ�-Rt��/视E}l�+~� ����~ݳ���!�YފN[K�A���q�qh�
RМ�(uD"G�	�ƴ�H�L7�Y�X�n���n�()}O$�ؚ����M_��}C��4]^��؝�u����
����+�f�ևI���]�q��[T��1*vi�֥e'��m���5����L�%�1p��[t�1�3;�sW�ky��i�aW����ukf�ϭ>�\���\�9�Q�:r�g�;��^��;���7 ZG�m��7+�^��w{���ߧ�֯�����V�W@���;�1�{�,ۦ�!�mm�Xt��y~��ĞpM�\�ِ��.��sF�vYk�-/q=H��Gã� �Ԏ>�W{Y�o4���%q6�~z""(!�7��? ���.��G^�Ǎe�3�5�sy�.W��w�]���l}��y�;�I��

����ԫ|�*fi&��묅�E6�б���h�p�H�
B$L�j���_!V<���^�z����H�z �[���L��ּ������ٻ5�pk�8s!;(�X�c�y��״0��-<��G��КC=�����6����W%8���OJ�&�%si�Ha����&���>
�)	/�t��H�f�z{+��'Ə8�_=xɇ �#&l���e)��������0SZ�� ���8��SH_@UKֵ���v֟�/�)��	���6b�}��;��x��l8�Z0����es|��3�,�l���\+���ھ�Ӗ��<��Ǳ�ؖ��M>O<̭j��m�m�1�t��s�<<j"5�r�>1�NÀ��|�O�e*c�ۢ>���ה�q����\ݝ}�g�0eĹ��F�=a�n��v�_=��2�O����\y�U�ɖ�C���غ�y����B�&����s��.u�X��/��u:��ec6b�u����xe��w=�2��I�vމV��Jb���z�>��f|�2>��ʑ�Ly�]��{���Db��ȏz=7d�#Q��5�꾸���q8��Wn�m�s�s|7�K���f��"������pȶ�Hx���=S�)8Ѷ��,�3]�G�y{���gJ�a�he�p�v5l�9~���s8��6b�'�e�s���ị8S1�j��ҥ�鏑&�i���G��
�e����X��K�ZM��=�o��m���7/�������Ą7)��}+ڕ�{����iֲ��դM�滿Xk���^q޹=�����y�X���Nv�9�Ӯ��i�����X)-��N�o�����?]]��2��]$2����3n�*NM�|�X����W�W�,�߇�[jje=�Yv�[h�|s�^/~�q�`��}t�q+ϓ�%n���0�rsw�}���˦���~��~?��Xq0��~Ӿo��K[�˅�V58��Z�9�wsچs���"���a�C���V���S�瑸Ɂ�\���k�n�w��c���ʆa�meL�r�qvoI�{׵��!�3n0zj�4�kR�03�����
��8~����b�`�����ܹ]�O!�_]z>�vW�w������^�]�YǸ�d~�
�w�U��*���
K���w��^�%��)f��u��Ւ���!�4r�x�:u����Q�u<*+6,�+�L�k1 \����S<�`���]��}�Bm�4��4m���3f`�ڛ���"FQƹ
	�I�(����ܾ/ W�*\3��|׽�7$�ML^�ɴn�l�lFc9�72�@��粓�]TY|�Ķfu�A�8�Ʀ��N��Ȳ�r������P��Z#uT���7,Z	����A�Hgo�\:�Y�,h�V� P]���LD��c�u2�t��d�n���̫���.�)�/՚��ukjW)�V<t���r��U��sp>��jT�F6Ń�+Ը���Qa����ws;�8�؎n�n�()v�6�)����;����C�c�4JZlk]B��892囸���4(+�T��&B3q!�հΰos����aŸ;on69���4��B��9���6�pˇ9ޞ4ا|e�2NH�H��1|���]�l:Um ������0�L#2,q��4��v�
�m��{�7%9�d��a�OOs�:f,5)^�E���z{��{�'��]U���w�V�h�C/�.��m��wPZr�2���7����)L�%+M2QZL��$Ĩ�M-\�4�Q��Qj�	Uis�]e��5M(�����QZV�
[E�m(�*�娩mq�KJ �(
-H��\&b-�T0ԶBF-D"7**�)����(`��X���z���O�K��D��.����+Y�c좪���w3G��m2��vr���X>M�5���q�rX|�9��\4���R��*nT��c<�q燡���ks�����M��������_{�q���%{�ۦ�!�M�c��&��^���o���{Ҫ�J/���-V��q��Cz�J�N D�[h��j��U��"Q���G�J�v��k���w�����)B�)B�-h�w2�҅+�h
-��%��4y�!��E�
kܕ��@_�CIQ(Sчs��=��m��Q(Z>4D�J�� ��-F�4cG"P�e���e(R��U���F��D����S�^�����{�E�D�~4qJ��(R���ġh�DK#Ƃ%
�񪈥
Q3vP�Y�0��+�k7w����4���J��v�D�Ch|Kh�DJ�h>@QJ�e*҅(Z��F��Z��J'.��=�vG;��%G��-<�2��m�A.D�|�ܣ�
U��iB�)BѦ��h"P�a���-h�}~:|�j~k����;�iĎ�����v����4��3�\�i�2��R�]؏�奛w�|�ƹ��
(��k�҅�4D��+�J1��V���"�J�F$(Z�j�q4e�4F��(IR�(Z1��Q(Z2�~c��y�o�)B�(�E(Z��D4����.�h�Dh8į!�4HR�GZ#G�"P�X̫J��b��B�=�I�経��V��頉B�fB�(Z#G˅^��m�\H�P��o	B�/����u�!�B�(Z��E����GO��6�u*%
{�kMTh���)B�(
)��-a����m�-�U��0�)B㒪�J�zUZP�g�;����}���G�iB�/��HD6�8��(Z4�6��6�J��@QC	Q(R���]�P�a�5���X���wU��J�����ĉB�i���(|~5��P�((H���-V��B�(u��Ѧ��[Q+�D���������|�<�E�D�viB�x�ZP�a�����e���1�U��J��n(H�m�P��m�Z�J�?���]��Zz�)B�i:��"P������{2�%D��-u����iBѦ��(��b�@�C�Q��{�ۛ���q��Dx�D�@�$z�DR�(R�)J��B҅��%�u�����>4F��(Z>&ڶ�4D�&3��z��\�̺�|J�B�~J-4�04D�kmTJ�4GJ�UR��J��B�.9M|L�
J�H�%���oZ���o���#�U����l�ҍ���b�����!��|�����BG����/9��Q(Z���҅(S-��-��h�]B5V�J�4D�J�j�P�f�E�֪�%
P����-cx�MM��S0�J��ц��(2rZP�c�JJ/Ҏ�J�D�h�m(R�"J�C�Q���P���7�1�2�J�ٔm(-*��C�*��ִ�Fk�%�U�G1��������䯈D�J��D�J�Ԣ�6�8�%D��(�e*4�JP�Ʋ��F���)B�)B�tZ��=��k��VR�+�_J�h�YKJ�@�D/�*҅�ǥZP���R��ƈ�@�]B4|h�B��)B�;�;z�m�E�F"P�h�!iB��Z�)Fd(P�Th���
�(Z촡J�U�҅%D�h�f������Ꮧ�coʴ�J>HP�KT��*%
P���4u�%�h"P�
|@�B�)�-�Dh��PZP�����9�Y�]p�F��ZP��iB�)y��	B��%q�i��-h�B�-h�h�h�|J�B�(a*>��/osy��r��B�}���P�[���P��iB�/Ƃ%
h�iB�|j4u���bP�q"P�E����j���{=/�;^j���4D�J���UZP�cr�J���
P��h�P�N5V�)^B=h#A�F�(R����a���a�7&~zr���b;�+z�:�"�ٽ�ܗ3r�M��hC1Ub��f*	�
0�sG�G�苲}�P�_I�����- e#C�Q��%
���C�P����������ӌ�9�"}�U1`:Sj��ښ���#iMτ��-:ךߠ��1y�w�zo����V�fڴ�� ��Re���3��fӍ�A��{ܺӶ���s<��g�ȼ9�ۤ����[��\C}޶^]��F��SP�w�����V+�N�d�����G��݊F�����]wSW��F�{M��"E�W����F�X<�s�8�:}|�ǖ׃.���x�y쐂���@Kx%W�+�䭚`��)�e��43�VL����s&J����u@w���x�9�8�>�r&�� �}; S>C�H��lM��ʱ����+SI��٦��O}�o����DǬ�mm�J�݀�>�����R�'������U�!}�h���en�&w5�qx��ƴ�71P+f�2�����&���ӟ=���e�<�mm���\}/&���g��s+n�&�ܕ�mKO	��9���9r��>�����l���R�t�����#Psf��1��}冯�À�V"��g�s��ᵳ���y���<ND���s����69����]�z`BwM�C`a6�)!����gm��Mλ�}@�p��ֿ*���	���>���L_.�X�uf'�鿛�~�6��3�h�uzS1a�b��~߻����8�r����DJ�ӭ�_=�s��wDKp����Ԯ�����Og�ݾν�>=ܢ��:�fU<�h�ўT�߅����W�/ꖽ��)c�}�]�|���\��N�o57+��p��s=����/]'Zi�GɇX���W�y��Y��]݇Z�)�4�B5����u��y�MJ�������N$M1c�<0d�`[n;����߭Z W�:�]Ԇj3uL6�2���
5� �eI#��P������Lx�#�]]�uI��*�u��_T	�w:^�\gܫ��J_�x*�=�X+¸S��3g�Aº�T��K��pu��x���sө}�[MB�Z�\j��`�n}�y�C�+��L���>���Cy<}[���oжrb�7�Sܺ��<1������P��o��q-�N�=������R��ۂ��`���%�=���q�DT]�>�]A��Wíwy����7��a3����%>�I��Т|}~������-�[ll��8�dBR�]��⻌]�ҷ�Gp�/7rݼĘ�'Y���W���3A�]��H|N2�R��N���s8�q�OR�Ms��6���)�Mc�/]���L�8�5	��眕�b����}짚ć��W�e�!��ɷΓ�{�c���8֧��5����y�a���Ԟ��o���[YN8ki�%����R�sȑ�7�uC���>C�WDV�����g7�fp9��Cz��r�ܬ\2��!�����d�u��i^
���N������pj9��yBė2�-��OvV�:�8��K�H���z�d��[*�7]��j��8��%� x��+�{�X�|-M�������Z�s��?*������'�0Ka�R�e�qۗΏ��f���gw�r���e84.R7�w	|����%i�s�=���.�֬�]�p�<��,�����_�����i�ƹgSjJna���sy���GW�
�r��u�)��zٹ��q���v_�[1���M5�G�w�N޵��[m�ݕ�vq�)��[�%�]��`�����UA;����9�s~��:{��l�#Yj����*5����u�7��;Z�bk��Ƌ>�- L���MҍMZs;���\����3�������;�Ԛ�W,�K5)\��\�3�X\����m�;ϫ�|�����ۭ�r�n������h��^ }�z�����kF
@��56��;�s����9���ܲ�<�2��w^%���Y�}���r�R� �P�q��Z̺��L9S>��)�P/×�C򋵊w�9�$��p��X+���x�ܘϱx����8�N�M{�ƪ��r�n��Ϋ�p|���x�|��uu����o�7��P"�h����+G� TX��]R���`�6���P�Zi��Ķ��9_W��>{��o٣2nCb�A�ō�ޱ��=q����c������nd�%x���Ũ.\-2t��Ƈhv�ĸܖIS{8KC$w�oe9v�o&;�JV�,5nޅ�û�_cw���^��p����ӎE:����f��6�@ٖ+���ܔk-�H�aM^S��!�t^t�ӭ��U���y�76�f�%��!ד9�;s�(L�]F�9v�����w�02h�3��`��f�
��'D��JeK�dzݩ؆�X�3�Kd�k6~G!�tĮV�4�/��ϑ=F	( .�?�׺l�MA�d�pL��kϚ�j4�����%d6��Mʔl�Ӝ�gN�K�t�}7bČ�9x)E�"G~�,�8��2�ˡ]�zLc9'��j�W�������#�������<�io��C�r��"���|��]����h����}YVo��fZy�e�����ڹ��+�����s��}��7���l����*�W��,�|�Щ�u]=����4�ے�V�.�nl��q^Yv�,�Щ���Ȫ�2Sބ�V��r{g�T�T��{$��y�"s��ᠮu\Y��.s�'�U�̰��/i)�$���[,D�F�%�(f��iJQ��"0�
&n�DLB ����F��H�R��2ż�w2�[E�i�ث@���-��R��@����FS)��܀���W ���AV0Pp�Q�s��*��� ����"�
�
#QS9���,�̀�A��n^$R�XG1�pՍ	��.�Pbf�	�v�=뙗���M����Vɳ�R��^s����>���7Ay��[�jAħr�?�{��'�1=��s=b���ɸu�	��5"r��Zᓺ�s�W&3+��붲�0��{����y�gd�2�a��l�'y�N!�Ѽ���"D8�D�͚v׳�=�cr�o����z��(h�#�m�4��k�}���]oY�ħ�p�AÇ� ��2���T+����7��\�\8��x^�������ޣp�C�[�_��sC��괯�Q�����deq`B�n��Ű2�⽺�����g˟>ٻJ���H��{�m�������K3��ו�}qM�97�a����֥�������u#j{*�C;7t��!���IF����x���ѥ���Q�^��S�Ϥ	e���u���Vv��O��9Qw[7�̦(?>c:�x�2�O5�X)��;F9E�ʦ���ƫtV����͑{{4���nͧ��[�t��&�\v��.�vS�C�m�p�EEʞ���ۛg�)��@>���E��#��w�q��
�$� ��ؕ�ك:�@5s
����1�)�&�p(����\-*�����O^oV��4So4:\Zmƶ�hf�)�ʿ]���B����2�Sܡ���n��̎�y�V(U_s�Ki��[�R^�=s�����yu����R��r���tU�8��fm�ٔA�7���r������6sOw/{�f��* ����9սU ��F���������?A5�[�価>0a~=�]��	��b�n"x���`-&p�~���>B�%���x���䓊NT�l︳�<�V�D��X���W��ONL�К��g@%b��.���^�v�c��z��:��A%������zr=z/��t�v{q�3:F
�TA��yz�퓔����۔�9v�!�_;|0[����ֻ�.]5�5�W8�عw*��?�U�}_a#3��kn%�4n��B��Q��u�Y5%-[�}Ǜ�C�]���9zYP�b��N5�
��Ѧ��گC�:�[s׾F�=�	��d	�2�d�I"�5������ǲ@���u�u�5�ϖ����,�Gޡzۜy���'�ħ��+���{�:w.�yl�A��b;O7]Y�NpU3XO���C�*K#Ճ:N���5��h"�%��Ճ�ʀ��W��}Vt����I��X���v� ��#���?8R��w�|�/N�5���Ƒ�Y݄vz�d����=���ELE~����􇞹��l}����%~C�9<��׬Z.*o:�U�Px�H<�w-�e�j�mw��S�=#m4D��g#b�v'dk��)�ONeF54%�W.\=Q��
��F�^��k�2s�K��8[�ε�κ� �t�#%TZ*�s��Dz=�Ö��;7[;D?����KK.�vp�MWZ5�Z{)�j^i�j���14 �� mr�e���/M��i����Q��s���^%���IG�o\m��eb%��_���q��p��p��D�<F�xS�lm��	^7�����Pk�7��uv��B�=��z^N6;Xy�諤l�2��sh��� �wa'��h֋���:	�5�y��rsTNK򾪨�
\�>��V�bNd�㨳�lm��}�,GX�j*�r�QkP2�5���ú�[�bn�j��^[�L�����+�o4.�a��x�m�S�c\\Ǯ�_�ԖND,�}��*ϩ^��6�5�)�f�����ƽ+��8&�ع�Y���% P�3�[�9�ld�ֻ�����,�0�b!��o�K#��=o�Qu];���Y�n��F�����ޚ�9&��~h��_o8�2S���o0L<5�n�j�C�����9�Z�
�Ŭ�sݣ��³��)���⌬��fz�U<�c�������.[}�\�_���}C�Һ�+{)P�| a�{<n�Fu��,�ejJ�T�8+�9Z:���A4B���zcr($����%��Xvd���s=�T�����ߍcͷ�5��O��l����mJ�/w��P���U_}~Җ�_3��.��]�)�<���ۤ\�ޕ�,���]��*Sx�S��f�}C�@�M��D���4s^�@ʐ�*��4�7]�C[��T]��ĺ��p{a���5	n+ENګ?�.���wˇ�=1t����E�\Y������H��}��l�Z��<l���hu����������H��O<:��y�r��)��Vcup�̫�R�fjݐ�2�f�}�j&��.��$7Y��]�`�(���A�,� ����Ԑ+GV,���'�b5��r��)yMt�
��<�uHwYn���(���-��TLU�Wـn�S��؂	=S�F�����&�u�_m����e���,E��uʬf$��b�=�\wF�$�3��Vܬx0jقP[�Q��\�5Ǯ�ATo(� �T�ί3wPK�0i��CF��w`}'\�t�JN_w�h���0�Qu���-.�����0ҎA�ۄV��h-���N�m[A;O��i]C/2�m`B�UЄ��y��M��a����+Q?�B+�`�W�:���r��_v/�r��,�W�2u�8�)�3��u_qgMscI�=� ô���*|!
t��X䬜aF�RŮ���%KZ��B%y&�4�wM*Z
l�ԑVփ�RLJ��e����� ;ҩ.�:���` �|��׳��R���^�;��5��8�������G��'�%�Za���!��%E��ؗ'��3dUJ.JV�"RA�5�1p�b��4��EA�w3 �(���J4"�F��"�S�ULB�HDYB#CJ�JfZc)�2�T����U���Z�(���#JF	m��2�6�T������E1 7"��l���a�D���K���p��KE��b�0�0B�0�"������!2�̊fX�F�Q��XcV�[�B�ً-�3��u�x3�=䰭=84���u�8ꀏ��UUf�2��F���[��i{��!ËFJs��e!�W ���v��gcl;ð��EJ"�N{���y�5b�)E����t�OQ-nԈ�׊�5i���2�{T.�o)�v�9^�򲨇��x_O����en�1�Uaն��+��+V�]�Qq=��B`������U�7�!kܺ'bu���U�B��������_�]HD�n����<f�;���;�c]���KS$�>���,�߸T��������C���E�X]�je��\�OY�����B6C�d��[��X���hk�ռTN	�����$�H�����T��/�B�9@� �m#ݷUua���!��z����-�;錊�}q����Sޖ���z��}����W�uā�V�dc�j�"��:۵vo0���^e�{�r52mcf⫑f�勃�6.�Ɔ�j��]ÛWJ�f��G��a:T����� �	T�?�v��,���P�+�C�����9�n���e��#���{�3?LOex��c���w��A�~��z�� d���X����0����fO �'Hb.�ޓ)�	�`l�3��Wv>�1�c9�1�D0�WZ�E�5-�\BIu�i7��2�^)yOm��]l�� Ԭ����*�y�C7����z�R�{�֨�S;�:�;��-B���Y<�ͻ��(��q�yגr��q�\:k<�q��9���O�-�[����:`u��#%l��&`�sC"���gJ5���kMd�Lm�����-p�A��hU�,��k��OQ�ٲ�NA����Jv���;M��u��(̪��C�4q��챊�{[�
�\��K��ׯ�=+��o��+@�:����<�ޥi��[��w������ޥo��q[����Z_n�o)]Í�+h�p���F
��b8�I��Du����=諴r>_����w�,��7ҸgϹ���<�m�ߟ0�����޻{�6����\8zA�n����=��n�w{���0���hQ���Z��G�ևud�E�8 &OA��}M�+}�gc`�a��X�4o�U�m�c��%[kY�^��jiMჱ�[1��^��y
;��wTЗ�<4Y�y�0O�hmT�%��pA�:[j��UԺ�ը���t�/0��ѝ�7{'Z��UUfh3�k?TyV�V��6��:�z����<B��WIb���G�&�c�}.��3y��gݠ�x.�䐅��'f����*��Z4K8��q�k�ˍ�&LJ�G`�K7���e�<5����m�k�υVB�g6���, д竰�M\�����j]���[��du�]鯞r�1}����x��K<���u�W;9��$�r�f���c�+�����*���k�,��W�Y�ܐ�L+wJ_��>۱�<�q����ư�gͭ����Vj��L�&�2�B��qr�f\T]��
����/�z�@g�y�\�ge��9bp.��Fu�}n���S�+۝�i�Mr�ud���??L}ۏ\Ĥ�X� ���?-�J������#~�:"I�\�)\Yiy�ϱB�\�F�Q�՗y�;h��>��b��Q�*@V����}�U�Xp��b g���P�t]pc~�iL��lܢ3�ƻ��Onl�ބ�^��aվ�����y�4�<����W;�J�:p���42j{#L�z�D�[1@hkil^������q�U�
�-�f6Bք'p��N֚�0��	$}�y�E�u���ue=�Y;M�Ƀl���us��1J��`۴�G��ec�u~c�h�x�+:Bi���P�������9h2�Y�FX��p��%J9%��zV%۟�o1��VP[�,���������B�̿�[�j��2��l�l���������}�)���V�����Qv�X�x��x�����R�mlG����`�����'�z�Ӕ�M���u^^��:�|���W�~�X[>�{���N]�t:��j_Y&�,Z��k�`0�ٸr���907���
A⣐�s�v���M�<X*M�v�������������q}7Qs~����ȼ�@��eL�ޞ��x���F��_.�/C�.�r�m��x�r�(*�{X}�+�!_�ko7��T*�v�g�����R! ���mP�;��[Y�.M�,�Y����=�U����h^����,}����HG+;Ύ�ж��9�;�i�e$�X�.5�	��H�V���n�i��&�)������n�)�l:Tμ�
��ίm�B�/h�a��Ƹqm��r��zb��ފ
B�j�'psR�wn���(!�L�����1{�Ju�.����4�N��D(e��s~F� ��J�x֦ru���ugk��f�E��WLug�7y���,��%Y��S���.�rL˰���� ��K�>�|�ui�}�c�n�9�:�!��=3���Zm-����{�Sr�EHނU+���IK�߭;�i�Avu�*���;�:�,���VU__��des���fٴ��$e��b��O.�<��e7��U�����M�y:S�+T��D4t����ȮФ�eJa-U�ph6�f�=q��8���:9ݼ��}��|J4f�wF>�>��l�t`cdw��)���J�T Lb�]tʱd*.Q�aN+��a�1on�P�1&���7`Y�+k_1bM%�ftwPb��`OJ�فoE4CEM��E�Y�i��a�NV؜��,)��+%<�7An��0%�#$ќ'cON]:�4�ԝ���yL��Ȍ��3rwDVv��7��"�l�'Wl�;�Z*�YFu"�Ŗ��h\4�l�(��K�CA��%��V�Y�*--81Z�F��r�\��DebU�$�2FC.48e��]�W0���(�1*�лa��V��Y*$d̵E�R�$S2-�-HDZj*I*"��E�Fڅ�\!ŌT��E���"�"�%�#U*H҈L��#J�!+���܈܊(���3	�H��"����,n�S*"b�V�����Q���O|�7��4xך�}�~!��3aW��\�ݰ��] x֧����vf�*ĭ�X/[c�x��Q�\֘�}<�'�ҩ����$![a��Җ�vs���p���*�{�ȳyP����+Vܯ9�E^έ=g��Wb	* ���b1�q��4�t�Q圮U݆�4��㘻=Z���*o���T�c'�;�=In8�o����Ȥ�7ʍ	r����n�dW�N�V�wq����I1�'F��0#��`�lʼ�Z:�!3�� ���l��~����ej�u�&�H浵�[C�~�o������Pp�Kʲzة���8��sP��ƃb���	�WacQΦr��:Y{�o��U�ʳ�բ0C���޴��1=G'�c�[��o5�m��Y�^TA�O��6�x+���h��^{�9�2�a����6��o�\�����0=L�f�^��i�2�kR�it�v��]��6s-���S�]�P\��k�{S��H�ׅ���O:7��N�ΐ��W�Jn�d�4�}��XY��<��غt�� �X7�}��oqʊ���X(-�f�Ư�_t��w��y�`���y����R�z�w��I�Yzqis�ˮBy=}�"�D-��be`[�BT7{)��h�!�=z��S��������u���乊��dK���u$�+գwc}e���h4I=JgVծ�����tM<���Ș��vvV�|F�Ű�D8xh���d�����c����Ӊ�㑹Nx�!�G����������q5Sd�Qyn�WWf�O$I؉kLM�b&Om��\��x�[�{/����,��	�����g
5�ц����RXS�g�t2�[�޽IO\�f�QA�0��^߼�3��f�l͠�ܦ�+�i��/�-P��ccP���F�'V�����,������f��ɵ��_l���_'H�ǻ��n�Ĝ�̤���]��z�,? s�ʳ�ݑ��%���w��i$��MKf���c��1�g��3��Sd�8�%�S�քǍr�k5�a}��e�����fV���|���C9�`o����x�;.e�	3{��ѻAq�	y�"��\ű`^t�ʍ�3�X�	��f6��<�=#���� ��+k(wvQ�H��"�K��m>w+��ߩ#��/wo��_teV��G�o�!j��O�Jm���s��a��c�sf6�K@YPS��v(������ĝm���w?y�m�3�e-��Ue��;�Z�9��6-�p�KϬ����e#����vR��x7�{��|Ac�>S��[G
]�ҙ=��iZ5�t�w�ᩂ���tK\�n�#Ke�U�^�^6�9#X;|�k2`�p���63{�������,f ����=&����=\�k�2v1ݮ��h]G`�Tj��O��5�f :]�U�� �V�[��Ή��}>����lf�#�:�<|[0_���%�����
���6���vձ���0��H59/G�+���SR��0t�Ҏ;����j����G���8������n\�ߊ]�rV��t��tÞ�n�ظK�{svRQV��jf��(���*�ܹ�����<?YK��j�)�0�.�9�q�8�~d�	=�I����f�)���L{��˾���z�f�?4�wՓ�A7?>Ou�d.��'(k��n֢ro��ȘB��*
�L�h�}Xi�p[�w�c� UЊ*`�\]5��יkhz����-y���b�����w�w�>��D�K��7Fh�r��[+)�H2��8h���j�0Rz� �Q�r��٫����K��s�8�2���������st���7Zq+x�}�HJ����1��Z�Z6�z)��nyQ��o��[W�w/�kyIn��&5lkTql�|�J��E�X���`���j����̻*��~u��O��m.=JG�٩}ʷ(U�F��2k~�<`;fk����cU�Wu��������p�7U�����jg5t5g>�w���M+:��9�99c�����]؃�2�N��?W׺�����V~�>�t��/�v�9P�����P��,�{N���q�<��h��Ʋ+z��m�,�}q3ϑ
O
�u�m��r]�a`�-nu�Pc�GX�"c�r��M�C;,�<����u|�.
�wz4������L�F���Ww��@5��%�'=�;:ՎO�֔�*o/fp���*&�58f��m�ugط/��P�IN��T��c Z1�:��g;��9;'l1��dZ�8':��(�q�6���	�����wy�}s2����x6o-�Ƴ��X�.J�3�d���]�
GF���u�f�uw��W<�kvuFM�J[��(��c����!�����1ѹ�Z���_R%]n����f�H����+��+�|����0�e�u8S��y[L�7kv�c�D��́��TP7�o<S=.��Y��ŕ
9�6"��	Rm\��!6dnb�<��ˤ˼�:�m���1�t{u=r�K���s5
*.��[@f�1�Rt�S0�^`��b�q]`�y�(K��c��;� ����\:V)�sOs�qL��\���^��Y�I��k��CFِգ��f̕{��g7U�^��:�y�	q[���r
	���;�RG���b�F4�լ;�.-�ܖ[([���Vd��PSw��0U��fMCjqP�cr+��n�H����$�s�N&�^���;��e��^\�H�$�����1��[-��Że7Z[kM��!p#lK%�Q�,�%ܶѡb,XIL�[q�Q�J�aq!��\�F��m�d.���X�V�T[ctʒZF����"H\�.I"��rIM�4I.
Z�E����V�0�J�D�e��D�.�0�H�[Q��e�7cpăK%�R���]աb��D���X�v�7*D�]�H]�%��,m�pUb�e�9ؑ+��c+M��y�6���ە��%���>�i���țY�[��l�0vJ�-�p#�ܡHm��7l]��//Pj���/�J���'���iC=�3���,�^��*���yKa� &�Pճ0�֗��ft��<��>p@V��ތ�v"&^�i6J��D�oEo<!��;�iɄ���H�5��v�۬v�3I�P�#�����K7+F�w#�mN�z[9%��L��Č � �
�v���+_-_�|-��~��P|h*ݡ�d��)6�v�%���Oۅ����͍�;���^ӌR��Y¦׆ze<�F��@��}�*��-{f�q�0C�y���~;Ev׼��&hA^(��F3��ˍ{��v?-����^[�����{y����Գ/!�+`��Z�IR�7/�ل��6ӆ���W�ВN���.�.�wR�K˵FM`�z<Ec��ƘYٕ�L.�iw#��.�������W]�xMac#ߍҾ-��Z���jM{x��SEz�n�y��ߌ�Ҙ��}���Hb��î���B����������i@
<���[�ިo�2-���w�������\��KA�kr��ÎZ�ۭP����[�I��ӗ�-��/���;���^�t3L�� ��#�*{�����cUt�R�ꖞu��hX�D�G���o&_�����t�	}�;{�DG����&\�:2unGg�>�</���N,���@�`�C��a�r�p�����:�b������)�TDεNw/.���E-�����f�kF]?9	��\��s]�F��q�e�
�1b���F�s��ڎ�~z	#�Y�Z�c�S|�|*��R4�P#�
>ޠ�ߺ�?Ix�<���+H�W����Z�sE[�2�c�'C v���sw�ʾ��Yj�R�9v�Q���>�{�vA����R�ԘߎɌ�k��+,e�.��-��brm�5i��5;7���4���O{4��Is���zծ��?y����[	��'ۙh�ͨp�mu�hFq���dB���q�a�՜Y�Y:�|���6����q	��<E�>'����Ӕ�U���a�ޚ�x`wY)���p	�{�EW;�-��43�r��n�e]�@��ކY�����K73-冦\�ܰ�u@}��z(t��~:3�ɡAM��s�1��#�v���}�8��xu�ױF^M��Q�*^D���&���UǴ��W���-�ľ�TU`/N��y�ܗ����*Bmt)����^e�l��z�����wkt��e.Sݎv��)��O&���{t��̪�ea����`r.�P���-<^޻�x�z���ٶV<�~���3��ЁT���a�ϹW�� k�K�n��_p������wkz*�WZ�â�"=�zG�� k�n�v|up}�Q��w�i�r_�eo,{z�Z��t����م�y��-�i$��[��@��gP.Qy���s1182��|3�ѼÅ���Œ��=�+"a<�}��d�Lמ�z�	��t}��p�b�^�'z��[!��q��(��Q/3Q�l�Z��dM�*�M��w�
�Kzv>��3�+gz�5U��U�������G.�@*�,�����B��Mp8�� U�ɺ�z��Á����[�\M�WkN��u���ۗ2��7,������_fܭ�vb��F��3 ݓ{����F�`ZFU�Nղ��1Fa�Cܔ�B��Ƭhu;<�B�j����qw��̽6�s�sG9�o�o�C�ieش��s*vM��tC�vxu
��T+m�7�ݑ�ߧ��|�Jn�[�Y�
,�ʊ�w���������	��hr]��{�gEo4��� �]�Wg��W�en���[!lu_.&^�M��,q"��͔��kօZJ����}}���&�c�ћ�WA�>]�.�Ш�:,��2z[�~�+F�1���VN�L�r��0ַ�4.9���&�Lygu���ς�O�-��8u�lSo�7CQ�ȩ~!��9��Jo��7&�9�79��V3,�\ڲ����ݤ\J��fn�C&`�:��"u&�L����%߾מ1A��~�-���\�þ�C�4������m��y����T��=Gd��	)$�Dz�h��`Gv�e/M���W[�
��ņ���AC�R�J\u�U��Վ�\�:��ϭd�]���2^�!0���~
��=�*�.�Q�iX;�w���sHO���K�2���L���V��z�0�~�r��s�_:�Xlt3�ol����'*8�x�Yٸo`�w]�f��a.	2R{��j�4��J�p[�g����n���56��`�������9��:L�/7��bА��@Z�8�e�A\�^��c��p�Q�L�)�4�p�O ��Q�s;�平oN�<M��(>��xۂ�vg"LL\N��R�.�=���fIr�H�����L��N�R��9��0�q����j��7�pv�tkJ�pk��
�h��V	ݫ�,�%6�kNň�ݷ�w`rq������$�/3#����I|p����H6��*���޴��ҏJC����Ë�{�m*��Xv�q4u�IV����#�4;o��0�&���=	�j��R��sx�Zw��fg_%�RNJ�B��ʗv�쮃@��rK1��hV+w����)}Hs�)���f�Օv��0�պ�mWM���D[Q�E��y�Hr�:7mgv��4	b�!�&�+�����8��G������ƍ;{�5Ӧ;�����i����TD�eݖ� �Yc�L�-V6�KJ�%�B����J$�Ĵl��e[)�$n�)!����mF�$���(���D�a�����0D$��"�FS"�j�@K�����0�.,R�6�.�$��H���F���1HHb�wwu"I#vKXfป���D9�5W�Kt��NWH���P\��RʗF<��9��4�d>k��ػl�a�mv�D,+� <��C9xﮛ����G^t����(s�1l'b�Km�#z����>�D�Yf����`O{��);�ȩq�K]�n~m������˟�����'֌�O��N�^�_�`��A�2����0׶X<���a�k+Ã�/�s|�ni�4/�Rx���e������8:Ɗ�n��G�ΉV+q=&�=Je�{�<�X6V6#�4���9]~k�MÐ��:�����!��k��3Bg�l�\|~�^�C:�F�>�w9gwv�f:5D7?m~��y��${�ϑ��ڸWt���=5+����t�\�e1Zͥ[$"�sov�po���}���}�%��ք%���~�!=k����]���vr=帳�<�J�������At�0%��n�f��S��>�ю�̭[Gx��H���W�������r�#�Fx�-ӓw�&��}���~��;x_9үk��P+"C�̚$��݉��¼�g��f�pu7�js�4���˃����� `Z��	5f��cȉ�M�,�˜�F�i��Φ���[���F@�W�R/:���k���Y�û��������ᆶ0Tt�j��-P�U\E^t�3��QƷ.̔%":�.�ӆD�(#�J�+^����m�}�k<�3=5B�1^��kA�x/?o�0�?o'�lp4P�<N�D���:XKV��Z� �,l���(k1v2����Z��)�HY��*��#�σ���>���{���l�����.�ô:&�ZQ��S��q�����TS	\��U�p�x����fؕӠ�����s��\�3�/Lޏ��t�W걞�y��-�dE>o{�b8.�.�A?��g��D������[����jG��ʯ��}[�y��y5�����Ӳʭ�J!vٹc�x�"g�r���&ͭWei���KC7��5vr���v���u0W����N�3_���M`Y=�9�
��jGYQ\�������[W�
p�tc9��{�X�xNe�9�gH��1���Y�˴*:���#�j.�j���|�8 ���9AwX������mk��4���=�֭��w�B��}�:JǵiE㗴�[�G2/7��D=W��ֽ�Ť�g���a��e���t��I���L�i�C�^�wwL�+�=*�A�(�wu�F�������eL�O"Ċn���y]z�o?H������g.��n�Yq׬��=�E8e�ַ֜r���Ab�#�]k����~wv�F�.�/�y�؆���}���T��%�9��ob����D
*�ݗY��k�.�M)�ӽ�2��S�\+�����͗Ŵ�����6��P�v�]7�Se��ܔ�ˎ�g��v�&�������Z9ᵽ0�g��ސ��`�n�xN���C�`!lt�d�6�&d��_C,�fS�����E�02�7'��[ld{�=/@&�lmO@T+�U�UK
����LU��Bb63�J{\`ɏ�XV�'v
y��kYg{�]��^�Uy�_�v4��נ�ɓ�g��s5�jiw�V��/�N-�D��u�v�Ŝָ��SYe w)\b��LC�r���-�wZ��=�sNq���3^��	����^罿G�-�������x�� �Dt/���
F��E�^��{�Ê��ƝW'�v+��3@��T�s��r��Ct�	뛴h/�Mg�Z�{y9v ��Ĩ��]���md��d~��9�5��>�?Nn���������Lw`f뎖ne\	x8��1�l{`h��jz�>��$G�/Q�#�'�+�<i�2j�3�{��ȾOw ���Wry�ev�e���:�,o[2E�;[ϖ��V(�G�-/k`:�@�oj/3\�w*���9]]ک���9�!u�]2|�7��V�R����3P�w�ز�G�j祉���^�yj��E�g���zZ�}���hSoXU,�"��ލ��|��tIk�՞,���e�!�nªg�p+�N�.��]PB���N<�l��u^ǌ��:��G2!���ͨa�҅��Wס�	��νq�9+χ��-����у�{������O��M #���U��u�#�JN2L�U���u�2�?�("��nR���F(v��w{��B�%����.N�*&��U����Y;j����jJ�.��X/@�\9�ї��z��S�c��j����%�փ�Ci5p{�3�ۍҺ�K�o�B�8]� n�lT:��0��#E��k(+���]�@m�8��J�W���h�`���q�4���tⷐ�<��v����!,ߢ��Ҫ�pI�u��b��a`%�#/9��#�����OB�Z>��N������mѩ���{�M�Ŕ�^u��t� ,U�.A�ڰӢz�B�(J`
��	h�-w\�e�/z������6I�Ӱɉus����ѩ׸�jy�=����\r_YS���u.�oX�2��sf�
�sZ]����̻����o�m��e����slEW}Q��x/[$�4V���EM�}xҩ[,�.�2�i�Z6*�&��*C�7��ɖ��ZW�k$�U�FS3Mu��vu`͹�����QG���:��5%%�=w��#[H:�/1t�
5á�ú��oO�_.�#��O)Q����F��*�uL)�fN�Mn9�Vn������32p�Ym�.�i�$���"5$)�$ZR��4�T���]�+JHHƕDFIN�%7��%�pQ��hZ�d2��)�p�H�R�.�VԺ��-*�e�SlŰ���e[�iv�.VJVB��4Ֆܦ�Ƣ��x�qd��F�,�\�۴��lFJaB쀒��|�wَ����gt�.]�w������ъ9����S����m����1mQ6��	�OVz�r�ε�KT)��V�*x�q���j߲
]Z��a�r� �J��'}=�N,x�ke��6�f���1�ݓ��v�m�~V<�HM�N����[l˒Hz��4��{�F���É�n�ܹO��:�@ѹӴ(,�Ž��`3��Ͳ�쮵���=xΞ�wͶ������6`K�Ov�-�*q��&��Z/d��c⮼�ذq��	�A\�ؽ���Y��'kz�v+�뀝��|r,ox[!�k���j�\�tf�����J��Ï���ଡg=�P�;���y-��w�۩�X� �%�ͦ����VI�y��d�^>�mu�*(����l��P�Q3��NN�7��)D8�d��}�Q��Ly7�[�~���bl�u�B�t��p���`�vz�7Z�֍��e���_A�Fd�"\��܅ i����څ�L@�,����=kb�ZzglnY���%W
�<�շC�tw�^��3X�C¯��j1p=�Z}���d.�;1�-�b��1�x�^J!}ӄ凳�]hW�ry=�Ξ��k�2ϭ��3p��MD�'��خ=�Z�>6���U�H������x�5�TOnc9�5�ר��V�UҬ5p�{E���#�6��z�~K�x ͘�G�or�PM͹S�"Y������4[�7�5Y�<G�˴����0+��Zw�zD��"��`�0�!��T֬In��7��]�q;�0t�y=�eb��x1��鑋W��Oa«{R��EZ�+&��o&�nU�NQ%��E����0,�W�i�h��+��5$�����ĥ��5���t 3~}�S=�f��i�s�,J���"�yq�7�����y��h\��7Q�t ��w}���;-Ȭ���@��"~���H�r���|v�#r������f���n�z- ��P�K�s^�X$�ON�V�8�Ƴvy�ͤ�`���^A�S>��-�ɸ|���ι�6�iJ{�R�c46�7�W�'*�˹��s��=M|�⤳Z�$]�Ίc:��5wʸqw��ȸ�.:ؤc+72S���vw�v��Յ���@p��;�?���cܤǩ����Eܹ,Bm2u?o��|*{�?0Y����}����ŕdd���(Z⋩F���K�����7�]q�J	��es=q�A���:�+#'.�=MP�全���%W]{��A��S=��$��n�����o�_<I�żL�<��آ���|u�����@3�o/e�w�3����� u��ְ	z,iv��	�f�[k�]y0�ҥ�܁�E�K2��Y�V��}Y�M��[7�U���;�xvV@��o���i�F���'k��9ӎ=�ޘ����Og���HM�]o��A������ls�^}d�T�Ґ�سB6�%y�]
�y�=�[ٶv4�����۪#�e^h���Z7���L�=�Kv���y�r{ұ �����]ޘ��\o	����J)�G�钡Y��>�z&�#�%��^��Jc,i73�ݕ��n
,�B�{���]VO!���tЎ��	�\� X5�F`�˽�N��l!���8LʨiF�S�r�ܼ�����|h��`3��;�H�|�	O-�"����o�`b�Fg�[{[0-�q+�f#�پJ�Z1z��)���^��R	��L`[�����xW����(|𧊇^��OP��5ƣ�VJ�`���9�dItP'��0��R��s��FL\���؝���9�"��,������eP�02�~m
w��Zu}�ֵ�l�OE���[���%������#!�{��x��f֎ֲR�!��5�=sЯ��8x��
K���*����;BK�������V��-mFG^�{��	���������|�^yʴ���-��>�vDѓs�9z�5]�۳�\�[-
�pi6�K$��i1�� V�����U�)Z�'E�b-; t�Ѡ�<ռF��O������#�/v9�M���J%��;���H!���έP���A�4�8��E����l�*��Q=X+B3/S=�����fI��6&Q��p�0sw�	�a�7��]��� %*+��7����M�f6/M+��Zq�-}���n�~b�Œ������ݎ��eg[�M���n,�м((���6Y�1T���f����Xơ6�{�b�/	έ�B�sO]3�X�%sy���J�	��U澂���^dףlb`'@u�c�%f�����8��|l3y:�ˉ�ޒM����dz�o���16�ކ�AپW��}e�W9��ӈ�c0��;H fb�h,U�K�V;���$w6�2e:jV���� ��s�%9�i�'���#u�*����G2�ˌ�͜��\E�~��T=S�� ��c~�ؙ�m��;���]�^�qn����]���#-��1N���`n�|��/����c��'���ǹ39�YK�n��e#"@k5�{xV���D�����H���݈Jv���1�.YO�t�z�N�������Fn�AE�H�Һ<�����D�V7��b^���de��#�V*�R7+���������ə�[���n�� S4���6�sE���ٴݣCf��>� ͢,�C%����录0m\ݒ70�\�_@;G,�8����s�	�<��C�n�5���rF���KAB$a%�˨�ZAF��t��Q���E���B�$�"���"U�.U��hZ�a.�yı\Be-��%܍K�	)I$KF�ꔹ�]��"����.U���S.PQ1$�)P���%�X���;h�8+=6dވru�[SxZ��U�Y�#��]�__�mw t����������~t��`C�e���5��Uy�}i��q����nW`U<7����ᆛ�A5Ƕ�fö���{٣;&�vjT����k����Du�Gzj6_s��s�������j;[�0ty�v+����xވ��!���e��S���ݜ�Ou�[u�NhT�/g\Ww��t2p����$J��
"\j�_*�.�l�	��q<S���e��vF_��Ꝏ6Ƌ�E�����"EL�Yp�=�����ak���7��>�(�����#����8s��|H!z��s;��=[vZ�OxKO�2d�r�F�"9��\21��"Vf�R�k8�_��~��6���D��{[ٺod��礼6ӕ뎌`���d�o#J�§km���]B�p�9��d�c���^�&�b�!�[��SD<;Yg0�;Z��i�R�G3N�	u�U�n���<��r�����iG���3�By�n2��jq�X9&��Z�'ZXJ�FM��}d��F�S�2�`�1��@�H�����Zꀲ����(�������ݤ��.�����J�cf�jb����C�ڜ]ݸ��k�]�x�x�l+ܗh��5���� {�ς��צ���\�2-!.Ȓ�]Vo_��0��ϰX���0æq�T����ۉ�,�h��)#&&��tC��Z�Oz��p_e�}.��+��yN�х_��7ZV�f�Wy]�K�*=Z��9�ά	�{7�[���{��x�+�'�|߻v�d
4���I�ڮ�eg�>/��hG��=O��aeY����Z9�T�y���>
�e�H�jP�/^��n���Bh���)�'�Ft�����o�h��ɫ7��(��5=���G��p��;��M���.|eN�]��bߟ �s7�C�`�R�o�Ms�j�f���vj��h��t�=S��\E5jrl?NA�.�@��l����vx�3��U∺牶k��I���n�;��b����OH�<�9ʜ\aY��>W��v�g�R"M��e��xgrܜs]+����`��Y�~����X}bCY1tY��|��!���W�f�fH���hwg��/�bh�t{;Y��?Fܖ���浹�=��M޵�����Z�í����[Zk��I}zq�,���R�1����8�]��p�6�:�rŤo1��܊���`�>Bz��OK��h7y]M{ ���pV���	��B�-��
W��G��߳st�/6�>-�''��+y��:kNs�F���7�*�p�3TNJ�+][��^�u��Vz3�]�>p�(X�O�E�I{�D$,j����4]:|�9NK�����C����~N�䳗F^!�\4��}����y��S9vk��ePLy0ÎV�G:���ۗ�Q]��3�o*}
^ɲ�cSs�������d�N�b�p��זM���	�/:,�qQ�{c_c�"�{C|L�Vbx�Pz�}��Ӣʽ/�g54���y:�b��Gs�е�2����Y��M��wV���������{��c&4Dm-˨�ۘ�xv�cr�%��U�C�`w�z�L�&��)�kn税����s�-�ZOs_��&�l��];m߽~�))Z���5{�͊ԛ�^�y��˨{W�L�멶�k�$��ٲ����9�3U��WU���î�s7g��KC^`盹���r c,���mӨ�xB�2)�C��s;ա�#W���������.�QS��L�e#�6o�/6ng��_u���`ɦus�΋�d�oo	�Qe���U�Yg;�����}���쒒I�L2Q���&�"���ݸ=^G��2�e)��u3��C��N�,�o� �����Nl��-r��>�g�C�w�jY�7P��ͯC�k_�ߩ�)���\o��p����Wa�	G繦����,*k:Z���!2��M�� �M�r�C�T]�����9G˂�����צ�wAY��Wc]R���6d�*�Q�|xfߎy����8�e�.���ʍ��y��5-:{���hY�ټ�{^fl�0�;�f3$�>�^gl��&����{�<�^׉�N{ų�1��b��ԚW��9�<���wj����}�ݜ�u�L��3ݷ�s������w�?L#Un� UU��}UT�U+�PUQ���t̛��vJ�����݂�d�p�������UTDw��P�l�l5ϒ��	U;�e}�PUQ��e��+���Ng�?���5_(������R�Q�����C�U���͵�c�f��t}	N����f7Ҩ���}W���������5A� UQG��U Px5^��*�����-�J�?a��W�Q�@��������޽������̇��?mPC���(������g���� �2U���~_�-P����Y�yU�ɫ@?�ń���T����W���梻�X?m�C,��W���(�
����c�>���V
 ��?�X~X����Z+�*M}M����M��2W׃�>�� ��>�Ei(�y��W�_y���_Ъ�?ދ_
���H}�*��a�������?�?o�h!�?�����O���PUQ�)�J~�W��_����~a�C%��~̲�T����~��U�W�G��t������������3_��o��q�B�*����ɤg�R��i���C�?҄��U" }PUUQ`�A��@UG�?�B�?C����%W�1��������
+�3A��}�EUF�G�j�O���C���}�ʪ���j�*�l@?A�kA�1çJL�1%'�uT�5WU�C���$��l��rQ�6�2U UU,?o�~�����(������?�S�W����%����?������O�G�~�?EU�W���}|ħ��p�����>~���?Ə�a�Q��G(������*�����}�mQK�
+��֏�UT~5_��g�����"������Ep���`U�ݺ��4�j��?��T04�YV���~h���~��C���:���o�����j�����c� UU���X�h�������㬍O�u��}���C�?�g���UT� ������:J���?�����}��O��PPUG�U�ȯ�h�c���aZ�t��Vwr�d�J�J��?�@����h��]��BC�t�T