BZh91AY&SYꩿ:�g߀`q����� ����bD��                mʠ�E�%IJ�)@�A)(
Z¥T��$��I"��BT�H�(�� ��Њ��R��@�A)�*�R��$�4B��P
�Xt�BE
*"�)RU*RR�E$� P�Iݺ�H��z���֔�*� [�R*�B�mk���6ݠ�
�
��J���`���L�J!��I)J�$HJUT��q��UUCz��D�X h@� �@$�� a�ty�U���,Sn�5j�F�0�w ���ޯ<����Z��Y4}uuZi��뻻�������j��oN��J��b�l����IJRJ n�υN�C�y����㤤�^t���5%{h����R�2���׷X��]�^�ox�J�ձ�������T���4���Z��=�N��O���U>�]��*�J��6�U ���>JJ����C�P�
������u)K�b�qy��CT����{�}g�BJ��y>��2ٶ�*��ϟ}*���W��<���r�h���zʄ�#Ͻ�|>��J��7>�|�R�R��oeTB�i@Ka�+}��*��羥*��i�O=�S�U_py���zȝ�����<�JR�5����T �����(�����U
��{���J'�f����UU{�Q
�Sm%J��O�JR��;��S�wܪ�ۺ�t���u�R�!x�}�`�ǯ;ҕ+ъ�p�ڤzN��glH����s�]3A�h�q�UC������hz��4�]]έ��H)�J��ؕi��"�>�*R��Ϫ�S�U�Jh�wѻZi�]��� �M.� �/���������v��.7A!Fra��UBT��$�����JT�S��@>��=X�sO���u�� Ÿ0 ���ִ*�r�@0�����x< \`�(kwP��B�ђ�	@����J�π�_.�9 Wk���Fj�t��M������x r�]� h��E wS�w��� �	�����7�*T�@�: R���@��c��4��Z�����O=��E(;�å w}=���� �����UU �ZK��
�}�)@w�}��t u.8A�, �-(�6>�� {�p� �m�⃠w���:G�   (      50��J4��d�0�F����1%*J	�  4� OLAIU5   b  ��&��J 4     L�$©H      CSiRHM���I��  PdK�5F��?�w�� `�/��SmUS�$�/�fP�_	�67���ePAWvM����E^�����_� �*��O�����j����
�?��$��B��XT�� ������~���������F6���8Ķ����6������6��%�-��-�al`[`��[#�Ķ�-�[������텱�&�Ķ�4���[0-������c��-����cl8����[��[4��[�[alm�e�����cl-���m��i�l-�����6��Lm���ǌm���6��q��alm�����6��L�6���0���:e��%��i����[al)�����6�����[cl-������m�[Lm���6��[-������[�[aM���[0���Ͱ�6�L-��-������)�����񅱶�M��a�����[�[e0�6��[1���[g�cl�`Salm��0�6���alde��6����[�[2�[�m�����[8��Salm���6���)�����q�l-�����[���alm�l-���i���6�l-�l-��l-���clm���m����[alm���6��[clm���Ͳ��1���[cl-�al-��-�����[f�[c����cl8�M0���[alm���i��-��lm�����[`[M��[a�6���alm�����-�����6��i���[��6��[`[[clm���6��[4����m�����m��al����6���cl�al-���cl-���[#cl-���6��[)����a�6��[f�lm�����cl-��-���6���cl)��alm��cl-�����Salm�l8��[�[6���Lm���6��q�li��-��M:hF؃l-�<b-�M��+lT� ��-�P�m���l��m�`�F؃lP-�6�K`-�ةl]1ةl� �6�b��؃lG�F؃L��m���Kb��،b6�`�R�l@-�6�����`���m��b-�B�l��b��F1� �m��ةlD��m���[b%�l��m���b�)�6�[b-� � � m�6��-�6�`��F�lE��m���bb����lF���ثl�"�lD�Q�"[-�6�[b��؉lA� �l�"�4�`��B�	l��m����b��RةlT�*[m�6�t�m�6�b��lQ�� m���K`�؍0[`��B؉l�-�6�`��lؤbl�
[-���K`l�
[-��[m�:b%�RةlT�*[-�����*[-���[b�l� ��F�#lT�� m�6�6�Kb��GlM�F�)l� m���`�Rا����lE� �-�6�K`lQ�
[��"[m��`��ةl� �m�l�A�
[-�6�[b��ةl� �l��t�Kb�R�#lT�"�l)���`���)lA� �-�6�L���B؉��m�6�`�b�b�)lE� � m���[`�R�lSLP� �b��lE�*�-���8�`0R�)lE� �b���+li����V� [m�lQ�+LD�*�؀[1D� ����E���[`�lE�-�1 � �[b����Bء!l -���[b-�@�*�m��؂[bl8�B� [`�� �*[c���4�b[�ǌalm�����6����[`[�m�l-��l`[�lcl1-��[�:b[clf�[c��-�lt����퍱���-��-��%�-�����6���F�K`[ؖĶ6�0m�lm��-���F�-�lKc��`i��-�lM6�[`m��l`[ٶ6Ķ����6�L-���;`[clm�l8�`Sclm��-���6�٦6����`[a�[��l`[ؖ�6��clcl�clM0�6��6�ؖ����%�-���-��#��ؖ��'l
clm�l-���%���6���-���F%�-�lclm��K`�cl`[`F�m�l`[ؖ����-�lK`[��b[ض��1�<e�)��-��-�li�Ķ6��q�lm��h-��-��6Ķ��[�ǌ`[
e�-�lbq�l�-�lm�����6ƙlm��-����-�lm�lx����%�-�lc�%��m�lm��-��������1�2�[���a��4���-���)��蚞6\
i`3��`��~�{,*�*�F>�$XTx�
Fۺ�p�e�fV굸�|]Y5��(�̈́�o�X����ؗ�+��XEn˷j�! 2������V,!
J
Ő���{�w2�,ڼm��n��,c�k�i��ij{>aqh."�A4!.F�wei�c�oCwFAz6l�M�
��\�Q7��C%�&�}�)Ď㊶e(�nI�tG��[kN�˗�ˆmq���p�aգ{y2'<�%"V�6�#��z�˛�h��НˢӺC/ 3f��D%�2�.�"�!�p�c��y��9��;��\�$����kѤ5��wFAߊ���"�D�����	ZOl֩�܅�xM��]�2L�.ޛ���wVh/���kc�h+9�pl)T̗uxS�e�zزE��6�Ie�:h�*�	N�mi�2��<)�h�R5�+�V���5v�9���R9�Z�"m`zȒ�,���3��[ F�ئ-^)�\n�f��];�+z�4Q�-k2Z5�wS]V������X;r��eYg`7n��*��I,�%,]M��9�+#��~���ol�TR��\���Da�	�E�h,���N@v���L�"�b5dd����q.��ܺ�t��AM���£)kE��\P���1��� �XoYՃt�J�ՇzA����w��:.��k�n^Zhik*Z+EP:���u4:7ݫ �"vm���ci�
��ґ,A�+ڼR�/	v�s6�P�3�+nL*��V���F�!X	J�&�M\�s�0�7���Ղm�(��׸oe�N���NH*��n�	㼕Bl���	���D����x�ƜWA���.(��-���J�x���ECa�4�FcX�Ed�6�J�%D,k�1%����^#6�{1�����ݗ�@��*�ye����Sw&�W��kW��ZM
)�O��,�߶��6ͱ/�q�,�kq{��0ݫ͋�^���hݽ&�͖�Dh'[U��`���V�WLm�ȍ�!��4��O+-�Ek��,�Q�C���Q��^�v�Oa��7v7Z�&Qm���)ʷsdJb2:[m�-4T�M4(��ܶsRӏF�Mݭ�v��4U�\�L��$�zm뉹�&�͖��h�tA1RY���٤�*V�3(M�c�zO�U=�j<w-�`1���͍��n武�&f]bx�\��uK�%
;���{�k�MIM��PPj���Ӄ1���(���I���N2�h�:�B[x�w5�c� гaP�4@ݥ��^�5ۄ�P��zj��${H�Õ��jʌ�G��<����w�
]���
�����5��[�ռA(U�9�($�s/oCII(Sj�	��U(����)� �E��x�J�c)�	b���T%Zݻ{R���@fDm�$���Ƽo7i:�m��Zq��U�4����q�t0���*�
�%�J�,<�m�	��-��a3��R�'M�G٥2���cA�gVG�X�V���r@(�����k��Ɇ�M@�E�Ĝ���b�m�$���:�F+2��W�A�b���YBE�2cE��"�9we�0I����E��ɭ�[��Ue���&�[���ՙ<n"Z!��f��HA���y��J�m3e����~�R�T��&�dK�sb�<Q��!{��L[�u�6��*�4Vv�#6���N�g�����J�U�nP mK� ��gE���I4����qLy�m�S��ܱ��6�B�;C.cyM'�^���4!�D���j	�/���ˬv���	%�%`	H�G*VDũo ��C��յ�����jt΍0��ON�׃R�ҕ�e�I#����toAQR�ZELT�&�ݸ�V�+�]eV��=�TŘ�`�Md����bVd^�Y�ËJ.���d!��0�� ���B��<�5��R˫���T�����D#��c����B��3p3Q�Z��y2�'`� P��F]���٠�����b7�.DuЍD�1���0��"�t3\�i"И;y3���K�`1���
T`��z�Z�W�s)e���J���wy�8������n��`Ŷ�n=a-:/v%�e)��V�U%\�>�<{�nX��6�n�َ4Ѵ!ӈ,���g]tn�p�i��w�U�Q��.�G(�%�7j@Ҫ���ӫ.�n�#n�j����|L�0�8���"�o2���Y� ��c��6�I��!�ӧ2ݫ�	V�]ӛ"-Q��4�ݸ�Xk\�G^���Қ4:A�y���g�+�U��P�I͐�sVn��i��y�n�Y.�"�"6��y1K��&��ez:��n�ZD�cYB��X��q�úw���YZ��7���q���
U�41�dޱ��2�1I�6oj�ZWQ��2L`3�<h�T�y4��L¶a(�`7zbi�PJE�=6�<O��ܚ���B�2����W�rLĥ�H[��*��^ s/n��;.���Y�����mU�clC�P�=b'���f	u���:[k�����U4�"��fPB�檁:�J��]B��,��(�a�@ZZhk�n�&��Dq9�q躺5��a֕��V��[��۳V��"Z� C	�@�n㊱�.��yY��ё�Wm���H�W2n��w��lTQ����{ �%���M:�����)���2�S�سV�
�A�ƥ�
;�X�Cf�ǅ�v��!w�7�G�fa��&�kW#K��C��ն���x�i$��x�XdVE`��ұ�6�d&��(mfcs3�[t�iF�׆iٵ&�ѽ�J��]���ɘ�Y����<%+�g�3���KI�n�l�Gt���M�bl[�ݠ.�ڑm1��+(Ũ�����-�����Y�$��N�M���-�Ź��%�۔�#��P-�4�6���aQ����j7��`K�snN4�H��1�q��T��A{#�v�jI&��*K�RɱV]4\y�:(V�ۃvI��ú�sh��N3�^�ٺ����y����L�c#��%m�,:�7��ɺӬ��P)��d"̗r�fP�w�L�R�蹪�h��U�ӊ���i��r8����n��^���]I�6	�+4U�mYB�TA�{DAE��ZJ5eǂ�2�ٗm��)!c1���Q�Fc�oe��v5��/aZ����%�����=O6�k46Ɂ8�y#(�8��%dV��V�Ec���cV��%���;QL��ǎh{�jcȉ�֑���w�e����ض�f��D����A�UV���t�!yA���F��+�FXS�a�ש����$VAe}����IvK'j��'�M�X�з����V��/w0-d�3���kt��h�N��-�է�+J�r�*��l�1�փ�eMGe8�yhU"k[����5�h|�\9m�/,��S�����c4U��o����9e��	���b�U��{�����ݓ>׫"��;��e@��d�ml�̐��F;�/j�
�ͽ��Ĵ<~������)$�(j_e�F�՘�*f��A�l�֝��{yچ�8X򪋭Rk�t�7`��-k�Ӡ�k�6��q�b�պ�,��&Õ/�VU$][UW��nM��3+k��]�ZۡǴ����X�P�9R"J[��/̫�V�m\����rE�:�
�X�D�J:ٸl�
r��
GE2Ɩ��w���Q��p�,�b��b�����=�IR�%�HFBA���Y����Ӱ]��:v���ш�V6fV�N
��u��(����-���ѕ�_��d��m]@4Z
�Tcy�H�F��S���=��#�P��j�,╤���A��4��kT6)�I�ʘUG�)�7�Yi�
f��74���6'�Zhb���Rm���#bH�̕�l.�ԥ�.�jSï����V-�*=Nc1է*�U;�i
z-)x�ª�&�K�f^:I=�Vf�V�QYM��h��R񟍀Fa[K�+p��r�5 ���f%�X�U,M����[���7
N���&�L�JM�n��.�l�����ʳ,�Kp\-�:۶�Y-C�l��N��e��T��C͛JZ�x&�U4j�Q8�K�j,m�0��Ee��b^��7�Ŗ����^̹h�l6s�*&�u�bÌh�VƠ�KVL8���CR�4u�h"k6-Fn!��nǸ��+�j�:vu��-ȁ�67cu>k�ׁ���O��W�&0�2v��J]��j�)��^���yJdy�ꚦ�f��r�U&4�2N�t+�V��֋�ez��܎�C/B����[��l�������
��:X��#$B�v���ղ���0�J�5	���٣��0^؇L��1+�{H�ZP�\�L�śF��-�][�[F�P�v��cL�.��-�2�U���b9�^ǵ��v�{I����*J�M�-"�Q����Y�B˗���v)��l��y�$����D�0�m��$��Z�;�	��ca74没Ո=����
�w�*���$�<�ڵj�B��r��\c$�f�{���7��j�`�rA�lX�,9&B4��%{��U�%��J��ܵt-�1a�SFRxש��dڳ�6�;sC�@*��<F͢�F#i�͚kK�F��m)�v�QFҋa�fm�����n��LR��M&ܡ�qm��u��`q�hlҴ��ù��
�����\�y�&�6^^]m���]�f�or�D5n�D�GJ84�s�5�����e�Ƞݨ�S"���sl�b�lٺ�-�H����a��7RXw)��1*�Eoj���EzJ�فa[�:�@��j�k�չ[�1�vܫp[v�c����'2��l�e��Ca_K��܀=�%��͖�y+х�7��Rݩ���+�#�$��{+e��`�K��+j�K��pt!ԲH��f�i���֋�������Ev/6��d�b�c�W͹�KG��v�@mJ�#�uUPÂ	N�`b���&�[��-[n���U��1 �Y��n�k���n�C�I����&6ov��2I7��ID4�<S75�Ҥ�6��:V6A��6je ͥ�~x6XJ!���e�h�
�>��f�iG{eA��������z�])�ִ�Y񔩛%�=�j��Y�hBn跗R���"���&�VY4Z��@h$�T����fѪ�`�2��X�9�M�z����[����Ֆ�اPD�[�$�:]����W�d�ᘸ�M��.-J�Z ��4ڌ��ZΧ%du_m�yD�vK.�(s;�Y�oH���#Nr*��^�<���{Oi�d:K°�;�+�ƈf���s�V^ω$�m�2��.ϑ�m����s�Ea�̡xe�e_t�Ǚ<a%�I�{N���!��7{�	
����;�2��#�$P�y�ͫ鼌����,�ʙ��L=���{o��!ei�!��yb�1cZ���ibN-�A�;k>_|��e�z������ٖ6��8O�p�g�Ѻ]݊e#�[".[g]�2ϣ�'�c�Q���E��dR�����VV��V�v��5�h��q�v��&e�ɇ	���vA�ȳ�3���/�k�^�{�<�m[N�v��%�*�&C�6���2��D�/q(�V�D��%dPu��(�z��7A�T��iD��$ڍX=ՠ�T�d���B'J�0�����I��U���\�f"x���vmC�c<�i�Fa��Zz03��nfb#ei0����/�R��^�[��PP*��j'��0�]ԭu���b�S\J��P�>DWx�Gh\���y�ťC!��qٚs��t9�k�����Ѕ���4�J>?��b�=�0�;��%��ĭ;��ʕ���yji�8���f��:�BQ��!t�R����g!����v�C	�vˇt�s1M8z��q�a�K�۶�P�`Ei�wOa�F�Pl�.&���Kg4�:�	��7�X[1��Y��"̲�8H���W���K�.��8��h�ƶ'���l�g�l�=�4�"�q��z<{p���U�PZxŨ�°�b":fȠ0�)E��od�xV����	�q�g,�+G	�uէ_�Q��N�6l�'	���!��4��]ƶV-�-sWZ��b��֜I&��☪&�ĩov����$����Z9R�齚^��CI+NfE���Զ�uD��e<UI�T�D��$�0���ZyI%�q�a�v��+1��к̡,⓵�t!fal�:O�D9�a�7eBѽ(����b*�^d9�l��rVe�z#ťq�t�x;��L*ӄ��iF��"�a42����c<�E���k�J]�5V�����Iű$�"im���\N���[j��f�gr`7I�@�U�2�E�kpmH�KmN�j$�P.\p��=Dh�@�Q����qW�w*���QH�D����bt���m��<�g0ݕg�0�(�\��B��8�\c9����=�f
����"��`�YI�T�V�d��O�iWSiZ|t�@P���,G�w��D�b6I������7�BY<q�EՅ���^ԓ���/Q�gu2���>�8g����;3�_j��*]N8\KT �x�UګS�hoeb�H�����hK�v�x�sM�h��˲��qf24�Z<IE��q�K���p��֘)��ҰKWI�Z4����Pޣ�UѺOC��fat1��Y����idT
�ڤ�&ӊ�(�U$ژ��%��4�%�{u�8�=��,����%�P:U�p�n�gt�<K%��=�P�YӼv�ɖ�x����Z6P�2������L�0�$�V�F�T'�Da�/����z�¡l垇����w\z�d�q�l�qy�7�g(6b*�ҙ��]�mxW&��h㬫9��$��7E��V�,5�]��]J&�$���&ҥ@�p�f��T'N�(f���a3´�y�E3�����<�Q�a7�:��J��Z��Z�*��?��$v{�����_���>�
�q��_������"*��w�;�T�����o�����}ˁ�&���*$>���}v�s�D�Ͷ��XQ?f!��-�Z�f�����hK��w3G7.�"fn�O���vC@��m�t2���{Hb��1H�Vt�I��ɻ���;]4<�W�T�*��݂o_S�v���l�U�tk��[��2��i���X��̈� ��Ŭ���I\5s���[҉�6K怨ij��<챛܍�q�5v��6^�����Z}cylM��OQv��k(�ҍ ã�꺼+���dO�ل�shs�vDr��zl��Un�;kP��5�h��-d�;L����일�Ĕ�.Ɲ�7�|0i4�z��msu}�3��֯2�_f@f�������U��u̮����;Pe՝�:�9.�Y��Vh`޳|�ȅ�E����Xvf�O�s���Rm�Yw���q�o4;5<-��x��ŪV�{r�,N��=gL[ÔtfF��&�t�\:��`q���gx�&����%Ub��u�%�#n�к�$5��/Vt"��>��#91�{�b��i<͹�ⓏI��cb(Fi�C7f���$n�a�=O�nݫ=�1�Џ#G�s|�F�i���:8���.�ٸd씉N���X6�=5]�����Af1�tSec1�ڪ�S�(v�h<��K��{c�:k4wU"+�%�V�t��ӱ>ض���Wϫ!��@p�:�ؘ�M���W;u��1�.9/O
��m�ה�9������8sK�0��]�ueLتKK:���R��Vl����&,���ne
�3F��e���^f=��2�wc���;�H;_�Д�_�z{�w��A	�)��qJf9�&�9+_N�v����o)M�J�es���3f%��ĸ�-}��Hn�8���[��$8�&�w��/�P�v���;l5;����Ɵ<�|q�5�
2�ҷ�3��}�u^���q�t��:/�god7�˰Wt��n�cHԋ�y|ճ�E-z��yS~�Y)O��N�\�[�]p���ĺ�gvj�j�j23�9N��{z���K�pn�LaҍjM��x'|Ђ���]�v�=�1�����I������hj�Vr�[Ǐ[�hӹb�?�i8V�Y��sjG��f�^B�l��O�"'V)�m+^���Bћk6�+GL�4l��tF�9�d«H�3Tv�mi�+jv>tiצ���� ��	/9������W����=ʗIy���<������X;�9���p�v��z՝yB=�ιW�8��d;x˙�)��1�;����)镍R��:&G_AhZf�Yf�tF�ӧ
�����kK7/WV�eM�Ϣܓ��;km<ۀ�ਸ਼qtU�[�z�4���Y<Ż�]�q�^i��߄t��@��Sf�X�j|6�2"������M`Xm҆e(���j#�q�`�x����;�NNo5��=���J�2���2�wv�[��`�w�=��] pD�Ҕ��z0��I�S$�XI�;��d�9)2��{����Sbb����q*��X���#����wX���rK:ҭK]���6i*�o7w0j[��ZT�F��f�;�cӜ�1͇8W��Pc��*3�ͤ�������_v�:K�p���7(t�����nI�v>*�z^	��Ӧ�D�^ӊC��oL�
{N�\aS�r���V�'��t�}w��
����5-V0F��Rq�;Weo���T��O��Euw���o�V��i��rM����D�jqv�-Y�+�&)ݧd��]�%x��j%<����zWx����	�V�`�̻�w]g�q¸mU��"Q�����r�>i3��Φ��6�_t��xm�y�כ����W=?Dc2�oiZ�FG�J��� ������j2S�쫱Д.�<R-���y�+���,�d���7�b��V�kYU9�B��WY����9�y:���=r��\C��r-���:��x��Ӽ*�d�g�u̽���goy�v����4R��Gj[���V��D��r<����^�(���v�ou\Fi����҂���7#COY��E��.k!���Cmi���g�D�}�˵�k4���[�fgaW|�Y��D$��jׇ
��0I4�:�/Ď����Q��uA����aR=\�dJܼ�;r˒���j�T�r������)���ޤ��a2�:y���MVý��wD=]�`�l<����^Z�Q���n����k�=�Q��&�z�z�b��u\���mL����h_W=v��D�}ֵ�BR6�|8ꩽ�k�̬2� ��^ջ:���
�K;+B� �f�B��ׄo�z�Xy|%��Å��5�q�.���aH턺�=|Hp�N�����:M�}(�lK����1�7��קP�H�jL��8^�wPς�/�t0��Y�LM��g��8y��D���A� ]������3�hX��!�-���malj\���[/_'{:9;�.vs(i�oetC7�����ot`�-���P��]:�P��]�X��xeyY7\���q
g8�Պ��q����`�JM��{��mGqdwӼ��]Y5�@���v�b��]!"��k�w{HJ��t;�}N���K�ب#[��,ޱ��\컹�f��ǉ1z���d��٦v[U�8��-yNR��6KZ-�g��]oW+n�3Zz���v��v#z�tE4.��4X�}�{1���Vn�h�y4u��G,��W�.�tVf���)wA��nބ�f�	u�9�sseCF;�v[�W�WI[���)6+sne�li�E���ˋ4]+*��j��.�I�6W��Cc����H}Oi����jY0;�{�O�C���vt��)lnUw��z�;�������7��ǽ��]�+:�4�t�}[˗��T86	g�.!�0+�D�1�d���������]
��R͚�@����bQ�,�l4A��2�.dn �Z7rwm�fR��v.S�=wuv��D��e`�1&&�Z58��Zv�f��@��9CF�>��\��%���Z�ݴ�-E�E�I�,M�����o���:���%��hQV�|��|�R�a���9f��<�qÏh�]�G��]Jqm쒻m�����񘃛����8;:��3�b|�W5�v��MC���&V5����-��r�[j���C�+3�$<���
�b��R4��ڷ� �m��طj@�\���;4v�H�k'62XqP�ܻA�7#3�Sٷ���7�,�����mT�]�3C�y�/�� ��oNDv��"�i�	���Pfq�g_-6�K�*eކ݋ߙ"�n���ү+q.(�a���|k%�<�w���N�W����س8�x��o/W����6{D�M�*�I$�_)X�8N�'�\O�!KF�{����2��-
L�Zili������]���Ỳ^G��gݛo��H<y���^Z������]�ȶ�C���"�;�oNb�+��͹�cq��7K'��\��v�Ju�n���]���S��;˶0t�Xh	3�v�������c�����.�2(��&�u%7�Y�j#V��XxG	�.��V�@��M��0wu%�.���v���Cb�%h�ȣy��ܛqX4x������WU;�ڠ{31fS�Ň:�5�ԙ��S[�hq�y�S�n��]��hڮ�t��F��dsҦ�5u�4�=�"s8PG�U3��V�l�]r�n
�n��.��o*=�uU��0�h�F�ߎS)#\��(F��=]���jJ�"mw([r�d��
��&�$�&�R�-gV9{�d}�\L�Ii�������N��K��o�ld��v4_o03�8�x��9td���tX��x���V�^��tٍD�b�z�
ŤS:��]4$���.�s[�U��W[ �V ��}�R=�ø#��W�B��"�n�D�'�p�=�b�]�6(|�)[��f+��B[��ضu�"�vW��;֧WM��5��9�:v3�t��{F��B�m�,R���C��-�]ӈMfs�g���{%CgQb�dE�&��몑X3�j�-Ky���B�Zde������l[��_9x�p����V&$t�����M��7'V�=.M�;tR���d�_n �:Gf����ӛ���Е-� @��fY��f��/~�j�5�w���%ˮ^턷(���-G0&8����9�Wi��-]�J�R���D�O��$���2l2�]-F^eN�Aśr�c<��O!跊��o-��(>s/���t��2��an��&���}hP$]��ݻ�ӡy
$U1ī�]@z��;���j�Kִt�B<Jd��գ�/��L�k��a�z�V!Ff5Y����������ݙή�Z'p�(�#��4Y��(�|�(�Pmud��՗��]T�9Y �/m`�n�u�܋��ܳ6#B��\��:�=��{fkg���4�Yˇ4CuT{R����.#��\�^�mE֧U�Ozn���C�����)(����(^h'��[r��kam3�zg{�*���ʺ�ZE�W}�^�X���-걘ck��Iṃz���F�L�c��_V�����'�sJ�}��DH�ħ���N�hӰ�����4v��ռ�[s9�SN�z�4
����[���=O����[�%��Tɛu����z��[l��e
�xFd���
�����9Z��]W�d[(*[V����[���o��0s�c(h@W��jL����bL���Ӓ���w��?vo�Kj��$������r�(���u����^d:�(��ɭ[]q!H�򉭹s�^d}K0-�:�n�{�ՙj��(�y�m�V[�_&�׻϶����ώ��wj�{q��zV�ghWpz�eX�tB�����g*鸖G���ʻ{9����{/{��0M+�^��t�ձ��ͼXz�84
��F�c8��&�0Vgk�u�
їvV���x��@Ȯu�y�q�ܫ���h����.�`���L�}��2�Y\�E:��V�:�� N1<�y/7�(�$��F��töD#)��|���ud{��9�慝�
��p̫���^�U(�)|����e�?+�j|����!��[�}6�.jXj�6�M����7�{��U��N�B(A��6x�G�ػa�\�[��ƺ˫�MF�in%�2���®N������������;a���}h�}�Y��+�TV�b�ԍ���k�
�bK���\zs/�N�ثy����g/s]9���0���8N����D�;�����>����<�˞��pS�ޛ�د�ԭg�+��{�S!!��� ��UР=���� #���އ�S�sS��(@�=�U���q��~~{�~��}!;l��ȣ�$I!s�7�dܸ�e}t	�����&Q�����'"rn#yB�j Q������<�n)|�Hj"�A>�	�C�^@*{�	�7�t���?j�20�/"��zb�(��"TF�\�QC��	�:����*zdj�)��u��$q�*	���ȣq�I9=U��n����B�����Tv(h���[W������ժִ�p������3rl� �@�/�zmI+��7��;9u���9YMMI�kF]O��[�Э�p��p����j}<E^���z�.��%���#�.�z�$���
(�����'��(�
��~�V)�EO�O��������������U���ߦ���᪾�4�YV�{�]������i�g�����Z��U�4�_-GBnK�����:��k���ͮ��I��;AY�KbU���{Gi�d��C0ն��Mwh��w���E�L�M��+8��Ws%�L��,?�$s����z�k���6�]��4v\�-�^��d�ը{�k�:%t&C�T;��9*�}���=���D�L��Cx��Y\���<�.P[�\�%�=;�����ͫoBֵ3~�*xf��v�����'��cv�-�.�U�qgv����e�Y�{:�A�&�Na����WI�N��p��{J��\�i����!��ʻ�*��84�
c]ܢ�gk��P�eX��q)�-+u��5�Q�Yٱjx���1t9D�ڶf_Ȫt����-YV�m�ҭ�L��4�R�ξV]57��h�n70�p��Z��n�d+���)�e�����a�qvz+J]�22������F��6N�Z6�d�0������*W��Z�U��T�L�{���	��b�O���޻�eq����q�Ǐ<v��8�8��8ӎ8�8ێ8��q�n8�<q�q�q��qƜq�q��c�8�8��N8�8ێ1�q�q냎8�8�88�\c�8��8�8㍸㎜q�8�8�n1�8㎜q�q�q�q�qӎ8��z����׮8��c�?R�
0�Sq[pmT摎I����{������S	rPC�悶AUUK���VC���B�T�]�*�;�Kc���;��Z9��vs͡�:�\��Q]�T3k���l��a��ӂ&��R��Ô��zE]�u�2H36�x"3��s.
b�
���kQdѱm}U��s��C�`Q5��[Z�υ�WB���F�EKC$ZA����7y�:��t�[�w�F���<0����f�֩L�����ފ5�0�A-!J�^^`ga4z97��RNJ�ѡdާֺ���w�a�����Q��t�ѡ�"� I!�X*ˡγglHI�uV��˲fTU�i�CtE�&`�ƻ�)���c�-ى�<2�wu�!)�v�y��˦���	�J��ܙY#Ϻ�U8w&^�4:��R�����C���+���Eog;Y�Ƕ)�9˄�<q1�끭�U�Y�����V����G3�텺{Etb{9�'Νn!3�O���J��u�z��0��2��wU���>"5uy���=�@ͯ�/�r����n�ν��wt�N2��4����7@�P���p�*[�(V=����G�8]
�;92VU��1�w����"=�7&�z�x���q�Ǐ<q��1�q�q냎8�8��4�8�6�:q�qێ8�q�v�8��q�q�q���n8�<q�t�8㍸�q�q���q�q��8�8�8��q�n8��qǃ��8��q�x�q�q���N8�;z���o^���q��e��os[��s��鬔.>��U�(��ZG�I,��YY4�a�:NJ���[&�,wn�#ǽծ`|@w�q�3��׉I6����uf�Dyy�/�WK����u���^���0*Ko�E�*��bz�h�X����}X��0�ƉE�c�K6h�m��B`��=O�����$����a���$e�·yׇ�uܤ8{xHb��	� ��'H�*��A�hᮽJ-&b��Ҧ�i1bE�<=�0�l�h�Ȫ5�H��ŔwV,�]l`�84�ZT�(�o�9Z���t�ҝ��+fKR� �
��y��Ģ�P;�Ĺ׃�j�H���A�s��5[��s�*��V�F|7u�隣������r!�S��3P��oN�f0���ц{�^.+CC�ȇt��0ʦ(v�7h�f��y�da�U�#Btcq��Pǯ�qA��4 �i�Ɋ��+pS�garf�q{��hb
�SU�kti��G,�u��F�h�� A�b�e�,W*h��^Y�]9����=٨q�9�����
�t���Ww��s;�dq�k���=^�	����qc�h��i���1i\zHʏ���T�s����^j΁���0���v���	��U�#X1�Ó�k	}_:�Wr�B:�ǃ$�B%�8 �Y�[�Rc��a>i�b�@`0�SȀ���A�";�����{B�K���y�U��V� "��]ς����]p�t��@dFD���C�L�s�w��.V+����^��_���v��Ǐzێ8Ӄ�8�?88�8�8ノ8�8��4�8�q���8��q�n8㎜q�q�x�8��q�n8�<q�t�8㍸�8�8��8�8�8��8�q��q�q�8�q�q�q���qǯ�z��׭=q�q뎜;��������^��]��u5*(����ª��s���os,Y}��Q(<%S����f*��`}���}�x��w.N��a��Ja�3-��{���1�]-=��hWS�k]k���[��� ��Ix���̨Kv���5��.��5Q�pܬ���f/ iL�v`,aP�ޒ;�YP�yQ�Z��ܡH���,4^&�.#0�B1���q��&p1�NE�on����:�����,�YT�V�������u#��PU8e-<L�ۘ�a�]]Ӛ�/Ez�ǉ*Б@a��ݵU��Л���*YlI$���m�m.����1��NB!;6��P�����c�i}$69sF��Aj6���s����25�	�^TD��f<�$�g,g5��V]�ܠz�(H�$"��+	y���c�:z��[\�͋�w�4�F�C�I7Z�\g>����
��<��Gk,tb��9�+��n�Gp䲆=~3N�3�=�5u$D�W[Y��{��јQ��W�Jׁ�ގ�J��mh�ٝ�;� �(����F2>	�Z3�s�է$�U��+H���n[�P�)�U��� \�� �Q�Ȭ[�_n�ȯ9��37�xg3]~x����׮8�n޼x��q�N8�8ێ8ӎ8㍸��n8�8�\c�8�8��4�8�6�:q�qǎ8��q�~qƜq�q�8�q���8��qӎ8�6�4�8�?88�8㍸㎇c�8�?8�i�qӎ8�6��8�׭�z�ׯ^�q�q��.��}�jMv�W&��ɫ*�K�瑪�tr,ܩӺ�THo�,Ҩ���X�C�csU{�\�׫��'��M���N��bJޮ:E�H�Ӱ���uV\���8v�[�l�ؔ.���t��~�,��_m�S��*КoqV��>�5U<-�>�&'��{��{mr��\��O1ںgE�w��Z�f�LY@�X_+i�t����-��5s�kyy��WF��C�)��{�������2�t�xn�'�r Vn��[r;s(GK� ��㎴j��\��q6SBnY�qkF6uuc�����R4�R�b�h���ف�DS�\:zc<D�l׹u;2�S���Ӑz�Ɨ;/��._�#��8�)�4}���R6`G�>�d�WSL'�>:ح���9���Y��Z�h�J���F��Y]��Uj�b��!�Y�Ss�Y�c\����:�d^T��iE�"*�wMu�nbz&��B^r6��@f»f�a�l ���.9�����9r����q��݉m^L�1�V�YϮ�N�ȣ���wAY˧S��@t�uU|�Oa9���3ֲ�8�#�j^C�k4n��˩Ð����v}���N=q��<x�۷�z��q�8�;q�t�8㍸�q�q���8�8�8��8�8���8�8��8ێ8�Ǯ1�q�q��q�q�q�8�8��qǎ8㎜q�q�q�q��hq�q�qǮ=i�q�n8�����qǯ^�=cׯ^���q�8c8H��0*@� $�>���f[�ٓG|w�2��I��-R���i\��Dl�)��wf��ძ+�3b���<����*SwB;��X��ݑ+��n#���mm�gv�fwN�a���m�D�1�&֍�Ty�� Z��MV��U )�\�$���v�v��B�[�Y.�ݣ�*��g����H���X��O ��3���<�ʽdg��Iml�����ow5������#�z�*{�ذ��5�v�z����q�[�f��qn}2�ބ�s��,��j��ud,#m}�n��8���u�eIWx�ft�T�������m�2�W  կw��houXxVJ��K�4<4�	�[ˢ����r��=��X���7*t�L��**�`\ĠۘÜ,��������Jv�J{��v�=�lb�u=�WwSv��SJb���h�C������o�e7q�.��1w����R]P����Zm1L�&���[�U�螦8�t���������H��p{���Yc��wCJ�Xу�MV�;)��b�u���u9��l�Tf�̱'$^YN�N�W[�Lp�k�9���}��ۃn�x�׏\x��n8��8�8㍸㎜q�q�8�q�N8�8ێ1�q�q냎8�8��8��8�8���8�88�8�8��m8�8ێ?8�N8�8�n8�q�x�8��i�q�q�q�N8�8��q�q�8�q�q����z���x��w�&�n��J�]ˋ�뭜���n�S���dko{���5��Wj,�\�,�\wd��������:���o�����C:�eͰ4��g$ŏM'��\��2@�������򰃂����7�ٺ7�1��]��
�+��.��Sb�7La4�5.�HQJ���{�9gXAgc�ƶ�.�KOw\H���ٶ6�Ls�� �	�HG��끪|/P�$3c�٦
ѫ٤Ws�3d�|m�7��;Yu_7�hlJ�VN<̇z� s{b��We�w��2�x�}ۉ1�ڝev;���p�W`^8���-�s���b���K�
�{:>���f��T��&�2�`����d9��;4�1_c����fΘZT�m�o��ަ��?�.���r�x�;�f��#S\ŋ4k�sGK����|oM�R�ʽL�o�+�g��sLj��ә��+dUq0
)S#��a�}��9ںFv�ږ˻���ڛ&��ө'k{չ�]t�2UI�a������zKU���# �wU×v,u;Q�X݄��'2ɫy3'I�{Y��"Y���d��-U��.�F��]p��xഋ�y���h;����k����cւB�8x�D<��]vҾ��ǉ%dWr���xIi\��r���k�b1,�A��k.�RX�Z���K��f��&��}jk�T{�&Z�!3Nr�#f�k���n�I�z��ɸ����^��\uMvb��U�Qm�F���4l���A3�Z����9��d�2��{��+>����9H�tƢK�J�����V���\YN�9��p�n�#|�^�![Wut��֧K�g mᩰ}�P��Q���7s 'f��̻�9���;O��h����-μ���p��,[�8P��8�*M�N(���v<Ĺ6��W�����AǤM;���{�$K��Mö۝Ҍu�R6�����R�ʶ��vE^Ų��_vm�����C�f`�i��MYe�B������eK��D^i:���n�YÖ1u�P�Y��콃i�)a�I�x�<��oh�Q[Vn��5y�K��z�$�(Y�՛���w6��sBIgp���8��R��}�.=�\����񮧕�'a�E�7nc�3�,!kj�G<M�c*��vY��2;]ʷY�ܒ�d�����X�jݰ���s�������~uʻ�xNMb�& �Uv��� ���n�)�#s+��j�|n�WKuyӥٛ��&�<��,�����	o�;�j�A�k�z�n-U��#,��.]�B�艺����6�-\�'_JL�nUTC�'5EOl�85�)���Q���ӫ�źv�c�Z#�ݐ��C,����7z�E3�ԍ(���z�-ewA'�R�:w��b<r҄�6n�iqW%oR�K���P*�&�!d[|7�sl"{1��p��+7��,��2N�2��M�jȱ�̥��V�ΘС�p�.x�}��WK�ݍG��䫆�'�k�6\���@����8��7b�X�]p��<q'���X��ݽ}Q�ia��շ^k�ûr����}*�e��Mmk��`���ܨ'`ya�<�f��srJ�r�1FK�7ՌΌE�we��֎	�]�uq
��	�儎�ЩQ�˻R��݅Y�uhW+���x¥�16ؽAF��E�պ�\��u��"�ܬ0�>�IIۻ��p��ak'-�1�<B��1��ШK�vV9J�T�0���07�U��1����}��횬|	����i�g���	����9�\{��-*��2.�_+�]�k2�܍g	��A|�v[z�sU�]��r���Q�+���6
��S�{N��E9�}�K���f�]��z�6''_V����=��[�zԒ��̳��-�^,srRHu�uv��P�uP�|��-�2�ƃu4`��w�.o4�'6���Mf.lG.�*^<�_ 5R�@:�H[J����X��o.��m��Ix��������ni�PE�<4�ReM�׋9#2��E)���b��k��̹���H���2�����Z��7�^��i����2E�EK珥e���Dc�@գ8I�V�.+yA��=KX���*��k�.���wg6�W��J�:!�n31�Zc�ItR�w�������:�'�-\�����EOe`s�IZ�	tѣ�E3E���]���(Q|�d>t�܊��V
���V�k���� te�7%�d�U}�)B��9�P����&�+�f�[�������}]�_*��������Ƞ���3���������y���a����Uo��ӌ��M�@�D���eT���hDT��3��p�iE��i�qH������)�	�dj��i)
+�qǮ���q����G��*������K̐4���^�T�6Y��%3��X�q/�tL���p2HRI
�ϩ�B�m&���B�@4хȸ�f@ �	"�*8��`�Tj���I��h�¾W<S�'yܾp�yw��T������I�Q�%��eQ�O>���<>�9�N��%i_.�M�CP��D. ˉ"�M�#2<ܮR�4��������;ʷ/���#!K�8�R$�h1!�]�(�HK�1���ss��6�x�"� �r
d����"4E�O�����5爉g/���;y0E��p4|p"	��*# m�yH�T��ZR4�l#ے�P&���CD��P�p0�P��p0�L4PJ6�A��p-5�-���]�E��= �,�	R�N`։(�f�(uf�+�yl�#N�"L��-n��S�ы9댴�l�ޤC�wb�Ӽ�C���`��B̻�}���-��YZ�sV�ng~l���h�Xb����ێ.sy�nǜj��9�$/s\��P��hT]��/;w=Q�\��sa��pr�,t���t$1S�ҿY�w�1��/��^��x����5���0�53�N4%�yN�����\k"���4�Է�������&S�y��=Y��*�"�ސHw5T'W�+�Ux�n�1f3y�h;P���t��W��;DI���u���7�p�1��ypN�XLʆ��V��ge?%�'b�]Wl��+�����!r7�rJ�ю��ėE͸���ɨ�����z�g(��i�}��*��ٱ;;�X���O�z����K+��0�dٗ�oWJ���V�q�8��"�+d�UՑ�%wwO޾��]�r<BUz$k�9sN�Tb�]�H+IS�;�wq�gz���`���pH�HHK$�H�
28�A��1!�āM�t�����FD q	5�(F)Kd8Y�)m�	���EA8b���d0xTJ4�Q�Qe�L4����ja�(�
(�i ��U��,Cl"Ae�%�B		"�pB�&Bki���P���qܐ��j����SN1��D�(�P�%�IF$m�M�m�'� �	�@[A��Z�2"EL�-� <���B�ԣ(�2Q	���Ar��O��ሒĈ�#J"�b6���1d�.[a4"!H�a�K0D24�b �DB�Ir�����&2dʀ$A� �@��)�GLp�m��,F�M���Iq9"q@�Q3��	m���%�Ȋ	��0@R.��
,"ф6�r@�!�n9����+���	���M1Z��.ỻ�*y�/#�ɇ���c�8�A�i�8��M�Q0�b�����%��h�:S<(��N�KHJ%Ғ(
�E�2�m4�a�f
�@�
@�1�Z@����b����ӈ�DI&ӕ�Ȝ.6�D��+�xPR3W�u��7C�<wx L4�\b>8���1��b�Ј�&6�$�	u1���di�(�����!�>1"�!-��j�=�(��@y㈵�dD�UD
�0�<ASE�`)��d��IF$m�	����SN1��EjP���cN"�rB�]b)�E�pB�&Bh��ED��1J;@QtEL
(�i ��. �EB�0�i�#s�2��8�A ܐ�C�D�L�֪"��LE��	�iHl�Lm�%"�8R\hȄ �06�H�����X�L�!	J��I y(��Gm����L��e��0G"AȤy�A,�	h"� ���B�kL�.U$�:���h�h�uUQ�A��6��nݻz�Ǯ1�rd%4T$(���$Q�z�y��AE���QNe�;]q]޸�{˷~y��6w=�s������ذv4��;v�۷��q���r���S��m5�q�B�' 2X0��Ugc�s��*�;)�PV��*. ���Q��cj-��9���Zӡ]�\L�A@�96�˂ěN6r
���Kɤ�C8�U�;ox�/���,r(�!9U��y���R*��WA�CQ������]�v������1��3�	D�J)
B �M�����Ʌy.q��17��o\�;T�b���f\���u�[θ]�@AkupO<�:��/=��K��ν��o7��~v�۷o��ϘǦO�BS+�-�q�ݝh#&�W��;6y��l�J�S������M :�=ז����<�պ;���Q���)�D#���Θ�t�����<x�z�����ЩkN��$�"�$�C�k��=�='E�I(�����?jS�)�{�O�nq�B���۳���΍���o�ͷ�=�|�=��Щ#�MJXU
�c\ᘦEEW$�;��������6Q�g�̊	�f���Ub����D.S�Ϫ��$Y���QE�z�c�.�M*�+_bQ������=,���
-RL��_�ϦJ-�&T�"R��ur�as2�!8_ip�L9E����Ser"�S��~f�/C���h�)�M(�KB�(��-F0HE�	0��K��&#%��lC�`N�d�6�(�#M��!��%�1��l����<�V�jyq��R�Ą��`��K/]f���&G-e>�H"L�%*�dX1�Xr$�@�@ƃ-�b�E�LPI"�E�
R���[���!p$#Y0 �ds� �PM�����o���T@N4��K���JA	q�l�T�I�*�)�
 �PA$��������)9��ʓ΁��)8Ir&㏅@�,0P&���:�\��h��QU����*��Q�e��g�6�i��,��D+A�PF����_,j��{�8��ҫ +��ᥒ��W�/�su�����@����z�u!��J��z�U��z�t߄��ޤ�������͉�t�@��ʊ7uD�ʐN�ً����*w�s�$	^i���ṙz*<j�jYL��E��X�I���cz���8�g8��S5�t�%*`}�B��vd��aZ���B�؅W��#�
��Ow��.�Gd��}��u˾���_n�<����,t��	A�w��ܠ�8;3)���ӂ�����͞~�C�p�;��U�b��rA¤:[���^�ɜ�����ޕ�0�0���6(�k��v�f�2����R*@9��9o=wQv�ي�Z�]	�����ʻ�ʻ�u�{s_�Ľ�DT��l���\�ݼ�.K���[��,|VL^�[�@�w�R��駗�R�v�C%*߁3�-Y���{U�i���5�׈^�.��u*�B�������@��Y\
�c�c7P+�U��gD�Vi��� j�{Y���|3�Yu�wһ��R��x5����1�v�}�Ӎ�S5z�ٲ7��^a~k[���Ϯ�k�Ś^&�6v�$��>+��Rؠ�x��Ѱ$\/=�07���kdD�dl�ͼPn�a=뤷�pl��ӣ���Lv�)�y6���j<�y��c���ĳ��J�7���dC��l�^��y�J��y��T��O��a���7�׾��:�R�	�'��D�>/r���`��G��6���_;��$]k��}vy>[>m��ƲV�ϷX�0��/Z�$�,�V���!3�p�[ez^����X��C¥�V�[
�cx�Bc@3[;!+����[-�33G�!��f�ܴxy=i����諹M�Oㆽ�Υ]�Qx�"�s_-���})�yd�M����g�u�Xt���0�NR����MA{v�
��Xr�C4t�l���}pd)s�,Y��ҵ��v^_3�1���k��o;8*����1�̗9����*�!Dܒ��\V�A]�Z�\�v��Ƀ'����z����Fi/�|}Y7��&���Ӫ��u��I���m��^�����
�b��j*A�p�t^�G��*&�w��t����v�}  }.�;�ml_f��s�W-�E�GoR��Ϣ���ˊ�3��f�M���Q���&-T\�uBȒ����T�ݟ� �]�� {��V�q��V�S����8�x@>��+�9O9O�
����4�F�[�^�E	��KzkƏ�;f�G]ɻ�mF2��/��t�[5�-l��+s:1^�@V�Ǣ�n��z��{�C��7]X�t�f�7}TŚ�յ��z̖���ʘ��NY������i�JZ�Cㆴ�Z��&ZG��9�J�٬��=LU|}7;�:��Kͼ1J~�+����ϒ�� ���*_8M]<_f5����9�-����HD3u���}>콗�Y��u��L��Vw��d�EQn=>�0� T>d+�j�x���Y/Gv*���%���O���/<�>r]-�5������p�^�G6mp�� �@{կ�I�9A�ޣR}�酗ܠ(�2����O�]u]!�P���u���j�ٍc���e�^~Z�{�p�������g�V}!���$̊�	�ْf��c�	5z[�%����WmV�iU�y=�i�x�Jh�toӨUյ��a9h曔�h�Դ±�o]E�nk�ˤZEo�	������?�R9���,�u`��I��7	!��n�ƶ����Tla��p "�5VR�ͣ��	Nl\��g��6j�F�'c ey���:�Zk1�I�15x���I%;+73Se����6o�y��ݧz��Kޞ�"WޭS��bZa����E"}y{:��� ��jr���UJ͒�hz�}*#c�{��e�;wF	�kkA'&.ݕ�,43�R�˩:��AU�r�s�o ��e�����#l�ۄP E�2���rD��X�V�V�ѳr�U;ޘ�惚M���Ѧ��wI�#ft��0ɡ�5֮�q1�[�t�ֻG'2�E��@˷�o����q�y><��	�Ų�;{�FvZN&�I�"&^�:N�V��Z�<�:㸦����$(��KR@�+��~�g�#&؏����v�J�l��c�U�z�9��,'�y���׃|���;a�!���k4��LdV�ƍ$q����f���Y�ܰȼF�{)�B��\��|Ϳ �:>���Y���{�;��f.�R�i�S���!�X�&�N6���u$�]�%�4��V��6AT$��Xl�YTb�����2?aϭq��y�Iii�B2`L�Km��s���p��\���<�n��AM[كW��M}���) 
��ӄ�L��`�M�IK�(oJ&��<5�Z�S�*��^�5i5��6��(�F֣;�p�g���M���w֜�O�3�V%����s�W��'���z�n>盳�����u�L�Uhi�y'��s~�>ڕ��q��ex��0����7piٹ%�������X~^��q�(CS�p?VUl��K���s�2��eX`��٣�q��v'�CΝ����)�w�1����WoU���Q����;-��2mR;9}�8�w��WP6.Ľ�@Z;>դ��	n�!%�AHs��G�W�W��K�9��/UDk� �]ХP+k��j�8S����N��e>b3TsT�b.,�l��lS������"� J͑H����;���UӉ�'#.��j�q4�A8��`Q�1��c-+ڥ=i��>�<�t���t����~'��{<Y�gR�aH��}��{Pmh ���si."��l�����_�9��և���
��s���A�t�T��H$���%�2�9guw�?E`\f�xm{�ϐ<�0�!�a�N>�ޒk�~��g��>�n�|7��9�u���oj(��3Ӷ*�+Aq�1x�:{��`��=T���J�/��W��U�'�[���=����ԅp�a,Cl��﷯�J�4'@�}�^�;{�~�	\�5��JHR�����&���j��J�U�G�P�!+T�Ȼo�>�]Y�d��!�{��v����z��ʩvfr.��X��Kg7{y��+]jjEd�n���]���nД�����b���GV�W�:����gv�,/ut��ѯAYYid�YGԘ�� @�GS|�.��Yxr}���-�,��r��Q����*l�`�כ��z����@��=�]�^߳�m�w����*� �y�6����W� �[�l�gwnXQC'T���݈3|��^eY-�Ġ�sR��FL��+U}�L�-�mmM��7�-���Kf���>�AΨ��j��bڟ6�I�'F����5�r��h��Aީ �d��v+5�S�Ϊez��߰����ݧ�E�=��F��*I2�
BnF�5��-�Ԕm3f�2�`&�5�ugm�d��{� *���~��4L�A�(���k��ݾY�iu;3W�9chP��S�;7>�Rj9�K�?+�q,���S��Ogv2\��&˩oq��40-d�q�N�����6
V���v*��g�A:B!�x��Q�[�}<ќ���1�-<+Bt�+6��o<ܼX�>�q�xw��#�GM���T�8'H��0 9:��Zӕ��[�?������f��fuƺ̋�3+3��C������ �qNê/��B�ؤ���<{���AZ��p��z�^&���$7w��g�r���cC"�Y[*������!�7fɚk3c����4>��K�:ч�@e��i|�^`���"꘩6����1�Y�;�3�,.��?�l����ZM'әe��x��
�8�(�/�A06�8�v |��NK=�e�U4�8s��Ӊ�e"
��AxW���3��'2��,�ʏFx��Tsi�y&/���dT�zue�t���u�M�*��ͱ"�n�M*5oV�m���#���0zgT�3�ٞ����7V�`�٣��5�ܬݍ�[5oT�=��T�]{�H!�y����[��4ocW��,ԥ��ݲ�-�rh<�L�;W|��A ��vB��zY
x����'��]�Sg`�E�eWc�Ɛ��޽�>��	�Y���e*En�����M�;�P�P��#ȏQf�v�Z%��� �m���N^�ީQ��	 �X�����A��i$�L�$��q0ȇ��D��HC ��+��'sR�����mV������ǟl��̏q�̬ŷ�s�!2^D��;0no�=6��<�cE
�8.��]�R�v�}���M�U e�3�L����'`�Vh�ˌ�[��u=⺼,���a�<���v��Q�����ox�3?��m�e^��e���i/-�lM�@2�EI�W��~�;���7%f݈ȝ)*U[r�\^@��@��>^�qB�=J�tJ�����1;�J��+���a)h���Kg�i�*y�e졲h0�y����D�Az�r��BP��烙�V6g��J��ǳ�v`�$�\I�j!�&�����wd�z������bv��{�P���?*c�$L�OIH�&t��I�û��S�Z���d���Q��A����7�t�si�y�Rs.�Bw[
�t�a��bj�(��U)�</j��1�?cV��	�,Pe{��S$�j�*��S�s��;��[B�q�R ouor�ʇz��(��L�� | #��96�o;I��|�F�v�f����O�5���:e�%�&�̉�t��ܙ���ō� [輛���I����ʙ��[2t̫��Hʿ,��Q�F�\��#9��~ɯ�������ş���&6�kۨ�)�/4�w�f��L58���0z9���'K�m�c�
���V�%���L�ed�;�R��P�h�5mjh�rJ��+�a(<eJݛ�'}霻�%+��Uƫ�	#&����"4�كOh�I{g���c�Y���mO���;�OOU�rV_}���5]8��'x�����!�t�7NFU�
��C�'KV�0�1#sɮ6�ܬwƔ��\�I>��u�ݝ1�S5��n��k.��x�ƻ�-Q����߷�{V,�~X��ra�	j���P���U��N�h]	�4Lp8���/�����L����������L�*k��s�*u�9���͖�n���#�s(�O�*�[k�>���[�ŰL+�xJ��HZ���Nn�n��N��Rg���$�nE�7����Q�јm-C����NG*X�� �e�i���C�re3E��}vBob�޵�Z=�P��,��S��oy�ŋw7'K�u%�!/�h�VXt��-K���.��'1�)��̾�΋���р�W��ڀ�ٹ}C�k����~���v߻H��C�_f��ָ�A]�u�SPt�}�z��vLvE���̨�6�����(g_UVg�[��f�n�͝ИOud�{��V��(��q�Jj��w�cf��o�P�A˾+h�!��9Zb#Np��<�*U����m�q�0�@��I��� �ƶ��u���ݱե��;3�,���ƒ��ڊ`�cS!q�-T
â��E�U�+d��s�%����
�Ys����Jv[�dI���ڸ*R�ʮ�N
v�gư��쫻�}7��[�����2��1ҳtA֬J�%����T�:X�^���0�p;�vI��񶦬bU�6At����E�*I�s9D��{��Q�a�;f
�-��.FYqة�B�~�pVx{��X���x��\�^�aV�7��&�1-7�'���-v���Z��Ջ$�Yk�����#wԡ�݇o\ȁ�}o��z	]zEM��w�v�_B�U��Őۗ��a�gHJ��7Z���P*�E/t#q����t׀0��.�р#F���B���N��J9�1,�+�b5��L��Z�GC�RZf�{�,Is��yJ_n��u�*��Ӻ��j�%<4V������9J��K'^��1]8��[7*��/,���m$��ɽ}֦=G{��L+���AbYt�v��o&ְ�ǁ*�5�n��T\�6�:k���h�m�LֹO��]�"ju]�bѺ�{+:�W8�n�2aU�&Y=�5�A�ԕme�0-�4DvԻPj��U��w�|+%>���7�We�wV4���1.�w��ΛL��DfVʺ���	���s��܂k/�����(D#�����4nq¦��f�4�X�*wB�Q�{f��\K'���J��Sɏ������W!�i������'Ճ�N�Tբ0���V�;�r߳�>��I$�顑�S�/9e?�U�V���Y
�T��O����x��nݿ<x����c����*$�$���$����_l��˅Y��օVe�'((��s�v���;v�۷��Ϙ�ǎ�d'�@ReG"RS2.XI)l�%eET�B�{���m�x��nݻv���|�8zHB�A"O�#жt��Ik-PR��!,1CH.�O�cN������nݻ|?=q�磑_�T������@�IQ�k"�BP����dT��HT�rQ�7:��;c��?<v�۷���4�=E���j2BJ�j�s��AK
��"9z���#���gL[�Q��gv��7���v������4�$c	*wTy�P�R��,ʪ��,����kx����I�r�G.jr��ʐ}�����U\��"#�"r��N�qP.L�������8TG�54$˖��#�G�TftȣZW.$��Q
�I("1o}�=���TQs8b	,(��
�zy]���X�3**�B{��K1w���4iy���q���L�jH�q��r�m��翻�l��}Y}�9�Z���0j����ߓ��>�-�V������������h�m�N�}v<�G���0��Z�͞��[ۑ֯���~���\��xx+�;t�<ߞs�.�����ֆW
@�F��}'Wۀ-M�H~e}Ϫ�*�w�}��0��?��ȱ�L����\���s���.퀍��X_�f	�z���v��z�դ2�E?��wu��W=�S��Q[U�7�%1ʔ��� m�qZa��v�1k:�#��g&t{��B%�@w���	���a���(��< �k����y->�j���~+tEЏ��+���&�_�Q���� �z`8s�o�\&,��������اx8=� �X'��PK3����Д~��6լ��@�=�X�10(�k��ǿs�uV�W4]���wo�gn=�y�2��6I�3�6������x�-L��
|�0O7����j���c���ɶ ki뜗μ�Z~��߀��{~�~wc>}�����C[��ͭ�{��WL�����]#�w[͛��;�o��"�O�SR������2!�L�Ǡ�?g�*�r��=� (:�պ'v��m5����}�R�)<zx[I&��u��1t2��N�t^wF5�D���]b˫ض�E�bA���ȥm���O�5���l��,���<t��-0��(�8�2�3��~�;�������/��-��`��7�z�j���]OD�̊����R<`7g��+|�@t�@|{��Ҡ�0�Γm���׏����w(]l#Ẁÿ]!���,h�Ku���s��g�骽�w�7���s�����d*E$ǁs�}3���3��|:h=��y^Gӹ�ʜ��J�zvu�D�g>�>=���3����g��!�9`8K�� P�>������ k���0#"�	^�	?�T��2jO��8o���W�و{��M�@'�a�|�x�@vר_zw����k��9ۯ`���
`���x��c��Ҿ�sx�� W�� K��A*���ˁ�@V)�� ���A��vp�ߐ�}^T�P+�n�Y��m���C[/�LX
קY�:m.f����`N8���Y�<�'�L��{��������c���_������ⱇ���y�ڞaש�Z��O��p0f\�?�0km1/A�/F8��^������@m/�� #�g��P�@Gʦ!�R��/���=��|)��x#�y�z2cLv�b��LǄ0.���	�+�I�@���^�g�߃�?m&�D�C���m�g���M��g�y}��y����ȅ�#��^��d�4pU�cx��k�2��Jv���e��[��{ ]�BC��5s��bm���wn��:}�9v��G�\�[&��[:3�f����N.uI��o=�r1{/����f�jH�)���41�p�G��j�A ��A� j�}�-߄d1�Zf�"�h�,q�b	Y-��g�6�q4�*o>�
�SW�%�
�;�O��8�����P����+9O� ׻����<���'g��AS}3P�����Tt�7]�#�����O��#���c�3�:鼘���*�����v�r��0*���޾��
Jn�����1��So��=�s��%N��Q���); ���eOl�*�b�z�Bl}o[t��%󅥞��W]�_\�DC���D����eN�r�t�3��{u�>���W��y碮 �4% �k�������ظ����
��l�g�.\�ƒ�_%�b�}��� ,���p��M�)�(�H�끬y� �[{��}w>���b$;s�:YZ�<���|��@sތ�5����c�b��<@w���S��s�}��fff����=�B6#�ا]B�j������*�^���> ��[�;򸀇сsO�gwH��zK����-�%n[�B�#W���h�U����A*N\)��]?<<� u�� ��<D :@��  |q���,{��;Ǜ՞�W���{vq��q.X��60�2c� FC�����Ch� �~����
�پ[(��G�����w�_�z��е�ɹ����t��k"�Z�3��ݙ!"�`	u�� ˖��`�8�Ҥw��|��w���U�N�oşi��w;9q�ܝam;YB�G�]E�R��u]-�+TM��&]IK��\���`���MPP�`�wW�d�ޯx��,�:�;�
i(w� E�	=!�J���|��=�W�i
��E���z�$m��7{�=��i��}��#>�z���+�@�X``��8�sߛA�|����]O��!�S}�]��p ��1�as'M����<*j-���<�P���ZxK��x6�|�@�Qp,�YN�	P��k`\��sr��f�'{����>v���r.5J6ǽϟ	�x�ׂj���0�ѳ��3vW7��_�7n&��'�,�F��i��O��:{Ƅ Q���2���p�+�`i� �Z�U[��p�+�Ⱦy�Y
q�7�eУ��dM-�� j�,��d�U�����;�w�}�ŭӳD���vJr� ����hs~�uP��=@��q2j���x	�����>򫏃�^�%�ߩ�<�4<q�՝�o�����s64�B�C m�8^F�����L����� ����eE��R;������<�Y/���K��̻�����zǹ��$]L F�4��� ap[Ɋr�\�Ժ �sc��\�/��V�m�6.c�1�c�B�s�����f�MK���D�<wO+Ǌ΋�}\�Ӻ�M���R5���]�ExU�9��}d]�ljT��ޛg�Z�ܕ����)'�a��O�S�������B4�����.4@���ݾ˸f���|�]z%\Bq�j�9�Qȵ�/��uܗAĕ�r��wg��ξ׷J��5M`�SCJ7���������+��??+�,�'i��L��ht��@ހx��ݐ6	��2Ľ��"h_2\sz�㪮���y��������
<0%z	�P$@j��I��ߐ�"��|hD=3�6D�kŚ�m��1����iop~�e���W����ǵ��ga$������!��&��W��A���\l׼lf�F�E��kɣ����#��>����ϧ�|F��!|�r��\�5���:t�@���1�秃}�KO����ngN���e��vH>���R:'ݰ{�� �oI����-���,�U��ݯ�wH�u@G�Z�hh-˭4���"��P�Tx;w����Ћ�:y����zG+(�|�����͈?�F@��1��.�դJ���ߐ���+>Hp��o�������H�h���J�`d�7s��'���]�84��������t��N@��~��i��zY+�f�u*�nY�׽K���Ш����)��^)��Nvv�c���]��	�f�� �W�N7��(%��`'ʒ1"��N
V� S\�>��ό�R��5�pw�ފ`-��?�t��ZW K.��7���6��i��t@p��Db�������F;j鞛P~�8�)L�EMT��o�}��ϯ$���A��T��Y�&��
o����y<ag���4A>&5R�*ޭ����k�n����+De�j���d̓��f�Ţ�A`�"Gw�^���c�/�v���ܟjf��T���41�!��J�*��*¾@�7�k��ׯK0,�34��-p2�K��z�
`wN/l-޺Y�Fl ��@ض����ȁiF�?��֠\���r�m�����! k�����Lt�U�|����,̊���U�|:��;�-���A�'�_;�u��O|�;��8!��HŰ-�����u���@<�	i�rTk����2���xT����=��Y���3��ZqpO�z�x<@Ü��ڀ#g���K���{n�
.Pɽm=��-J[�����~o�*�ڥ�X|0�*׆�;kx&��>�]�0����wt�=mu}�}/�1��k_�c�6��C�󿃣��άK��0�|��c��a�C5���Y�����S���҉<����pexk��s�!\G�u����n���$d���4��2���'s�����;�9j�0�s�=s��`z�c����v�q>)R�iJ �MCB����9ev�PxS7�7��٦�O���٣�a���UR�{k�j���N5���k�O�
�*gQ���9���=^�ZG�����@�=GPF<w�P,��"@�U���3�7��z�}��Ul�Ʋ��l�en~�+A5����W�G:ˮƝ�"λ7�u!B�ko�2.Ahk�����8��AK���S.�|����l>|��U�,wKEt���{v��uv/i�\F�[��D���ٵ���~�ghi �.0 ����L����N5!0�䜁�!}u�����T��$aDcK�0�P��_hGƑ���DN$�l���
�����}�P+7���<H=���>4�f��,҇I�a������X���Ws�`*�t���Ō��[�c�`Ś��-1P�z|���XE'�ސ��^�׋R,����I�ƈq�î<�˴c�v�A�c��l(wĦ�ę��U��t����=Hf��z9_ 	�[y	䴭Y������㳵�l��ܼ>����3�N�¬��`y�V�w�����^`}�-}LC>�Mm>��`�����F[���57Ci�eF��oT��ζ2]�f÷*h��j�0ro�X_��$+u�n��<���1w�]ש��=Ru�6�7�˖�����$��a�nc�^q��CE�S�ؘ�ˌ���;B7���m�tƧ�P E7k턧�>V���T�Y�|�N��a�:���g�4((����W��TH"� �(�d�_?z.9y<Gz�L��������X�q����h���TMq}�]�-��H��z����������n2
=85�l0mS����C�a�ScR0��c�W8�r����zaػ]��Y����:=K���|�
����G����q�+������e+��I�oJ#��ٜ�j�f4������]��L虮��k!�}�� ���N��7�)+����gp�ڐ��Or��f�Kf� �p��>"�cj0JV�9������~O�|��gM�ɤFF�ܿ���>�l�T�m���_u��),.b�#H�͊绢�|�w΍:>D��I�� ����R3�R��ޫ����;�!F�Gym��KE�H���Q��M �	����ZA1m�{�3�4��5�� u~>
�{.z�k�v��C�7ݺ��n���i�lco'�D=��A��OŎ��}�+��52|�÷[�^�rSAټ̆��=M�kj����H��p��L�z%P�m�Q��\WD��:-��c�^<��}���{Hs����Ϲϊ�6SߕG|��F`��5�F�F��I3l���okU�k�zzm�uh_}����������H���*3�܊��(J�����.Ӏ�-z���Z��I�U�~�S��m��z���R*#���ܤʿ�0�-}�i�):;^����Xs_�]�y3]�ŽY�������qy��jT���f-���f~C~��>W�z��4"N^.��QH�����3p�aܫˏ�[��Ve��;r� {fn/�J�EL�0�|��p��7�K?/�U�e��~�{#7%�[�P�De��P�����وon奷�/1���T�R4�����T@F�1]��p����ca�8���ܤ�:�m�7�J*�z�`�6���������m�S;��-X��,O��A������
�A�� z*Q����{pS?�>1��o��qE7uE0<���!��V��t)n��6s��x`���;Wp r�ׯ^�{�a0�ƧX�SM�qM��m��q6�CLXYi�������Pq���*}�6����NS�z����X�G[�V�᤭׫Y9�G. <�fE��4y@��Ƒ�fe�r�>��%�(k{Wv����`s�wz�7X3{ܕrť����c�i|%��K�z�ON�����>O�W9|�[_�}Z��|f��۠Qt�RǕ����x`���~nY�R1��@HiЅ (=���|wx�]�>G�:Z7i�r��w�Y�v��M�.1�UϓV��@���Qw�a:���_t���q����sr"�o��~5��--8����%�AU@�wR�VN^���;�t�cd�и�������/z�sά[�v��6yӦ�y���=�� �:F��-��YDP�G���]��O8�w��.�H7/���Fv��T�\;����5�l��:�40K�fe�s+є�dz�h�����|���*D�����q�u��'P�)�v��Hۛ�E���;ӭ�o�tO*#j>�G;=���3��(���+�����]
 ��r�����>j�QE5 y{&��`�������'t�Fo.iB�.Ԇ=�P�+���W��d�&IFpa2`�	 7 Z��������W�Y�_���K�L���e���s���Qm�`l�4z��Y�@�V0��ɫL�̓��H҆hCX޸��'Q;��#�����*׾X��)����O+�^nK9�~Ѿ�=��C 	4� �=�S��c��,�3�w�O��^��On��c�����K��k���]�ǩw-}w�����T��i����kK��ʦV=��$J�=���������%v��>=���f��<��e&���w�6|.�= ��	�{܊.�d�]�e��;�
Om����4�ߣ~������dPyXAz����h� l�o�|p�}�:bieG�_J(^�Z�w���Z��8%�G�~�p�I~�_$ �#7��_2r�@&����
���O�#�|�ݦ�+��b�e@ͨ�%���ۏ����\�K��7����	�_��AWx����L � �������Ί�$w�kxt:.[��h��l�Wm�5ݼ�c;��x֘t�m�bp|�)ӣH^�o��y�`U�v�>>3q��Zγ��B�\��?T%z��J�%�%��2��ٖp�\e���8�Ql��2�{��'s�9�c��Xx'4���텦�K���H6��)u[�����VB��^��P���r��A]����;�����[ZeN�
�3h^=���AW�4C\;oF�\u�����T'���e�G,��,��Z�����k*2Q�`#eN���q" X��r�L���")�˧+�p���׉m��k<�ǾUʥ�q1��V��k-��90z"ջ�f�h����Z��I�Jaý;��%����mb�=��F�:�����2�
H�& �ww��z7^ڹ�b��P%�b�NJ�ů+ٴ)�OǗ�ZU�0�������n�7���=uGf-����ֻs�C��&��p����IV4k�f�O��t�X�z�<��;�a��fY9R���_�,=�����༬\DP�A24����͝��T���P,u�H��M�AY�o��]���ft���Vl�����s�9f��ѵ\.�-L{�[w;���U�_x�"9��D���ҍY��9\��Pc����%[.#�q:��qփ2�f���T��c^6r��E6�����U+ε�ȩ�����+A7��q��K���]��>���1�s�.�w	��Wܑo���oL��F�[��qM���V͠�[���޺PW$��uG֍�1r�i�A��J^!�*2B��t�r�����Ij"z�(И���$����l�!��yk�][��b�����&#��~���	`OX��H)l<�.�J�&-�JD��D~wVp��:�C���יUyN�t��|��[�/�n��w�f1���2S�|4�=��y��s�)�ff�O2[�����ڕ�Ԩ�풮͎u�uL5l��T��)fR��
�Z)@ś�E�͖Ԏ1O:��j\��Ŗ��wrJ�x�J|:����Ax�U���L������ia;A�ٗ�cY��u`�ƛ���I��EQ7hB��'����Ɵj�����Gip7kt�*�'�B&H*�S&͡FL�V�n�z����+�A*c�>8�K9��Ӹ�WC���W�(��0Y�zy}���,����7%�9"������Ļ^�˿:G�Up�r���\�u���n����p��as�ץ�<�pfu+��qO]GR��ݩ��l��X�v�9����ZŇ�%=��C[Lq�2�ܝF�b%a��4���G���ͼ��X�]���:Rח�N��
��!t7RO�|��wr���hZ�Ӆ�f�T���+Ӆ�8�aY����㽃e�Q��m\q.�׍5��vc���f�jg!0�E
Mbk��~<�U">c'�s�`�W"����[�۔T\�+D�#.��BD��1�Lx����v�����1��Є��PBBaU+}�]�\*��P�q*����$�R�dh�d�����~~x�۷o��_4�0�C��w��W�#�G�vU�}���l|��t�L2�Z&�tpi�$�P����t��z��nݾq�Lz�4BG!���[�!32��D�z���NU�1���Ϙ�M;x��ݻv�|��g|�!���\�ZD��vE2���!:W%VHQUj�QR�1ӧn�<|��ݻv�|��z�nO���J���9S�r4�3"��*&j*BR��M�c�N�x�����;v�߷��Y�7�~�����*=>R�Q�a�:Ľ(Zy컆b�>�>P좾6EZ9Ĝ�T��S)P��#R�r�;5���
��G����kq(�%JQQv2�sH�T�G'�U}2;���*�>�����!�C,�#���j �A�	|h�H���Q�
eJ&M�a+���8\�(�|E�e�҅��Z���|e��!��*��Xt�)�wv�pʙ�&�<-��Kb�]ʖ-��+=%����Z����V�]}ph���7���V�a�3����R �FB�q9#�FA&p�L(I�&�O��$b !��D��)6�l�D�Ɗd(q8��M�#�d�!dIH$h��M��\wxË�]��iKμ���\q�C!Ƥ��Sj�!`�H(�r&� �(��)
j&�8%
j>Ah(�r2���m)E��r&0d8�� �A���A�,+H�'aLl�`��{9�WߌxQQ�_�F�f�u�ְ NRk];�y�x�t�dV�g���;�(O-"��J�M��_=����@��:`����g����C-�b�+�[�]�Bə�V�]��j���a��w~~ a��E�U兑�|��M�g��z^!��s�{�]��xXP4�M��:�f�Z��<�g�����s�B1��G��׭m[�鞥ƻ�{2�u}K>r݇=��t��z{�{�<��0s�g�B#�N{�����$;���[7��Gsω��"4�g��_i���T�3�o?1�Ma�S&o7�ĳz��`,�*y�($�2<;�4�G<��9(�ln�}C�7�o7���츞w�f�Ś}�0�'����l)^���.e��9'dȔ3����^ "�]J�(l��>��`b^L���'�`�.�>I������|ux�N�����n�
<��bx6���z)J��(g��;t��a��|D37���^_�}q����Bh�[�v� �[L�%\]�+�Uj����w�~PZ�	�^�)���ĹN�S[B��0��v�ɿ�؞���vqv������;jk~\�}�J�k	v���b*��,g{�u,,5a�GU1��h:�V�z�/;�_Ol�c3�F�-R�C��C��>�����k@��?q�����@��Q4�Sھ��qNnQ�Ε���T�;�e�Ƕ'��;aş(5��@�o��~�
0b	"j(P� �[��Tuw�w�g=����e���|��{,_�s�yC�S� 9��ĸ!�+c7��J>9рqd�x<��g�1]��i�-��w��
��i���'�g�s�C�Ϫ^7CJ3�Ǎ@�¢��r���iw&:'{n�J���5��[���Y�󅂮`a崹�����L������z4�	�XѰ������|��}����@c
�O�{��"5{�'ѝ�'֠�z4v5�����-��C�i.��V�{}��1��~^�6Q���gՓ 9�|����U����i�����9�%��>��g�<꼍TȎ�M�W<vq#��@$�0/=�R'�(Y�<}~�.$~6N�������5,�~?�=�XT��`$L�	�1B9�;��T_y��u��Ƶ]!�	���`.Kz�s�7�y�	��3�:C�=��6�W�����%@��H&(10o"����Z�Q �N/vp*Y��>�������~��F���d�x�ߣ8�sQ^z_-��b�Y�m����R�k���;�i�y�"��O ���Ȗ!��ٸH;��I}9��C/�@ޯ)ܛgO���J�r�mL&�xk��'18uv@�sH��o�����/PK,�p!]x�ل1��:O�!�8|+�^��
 �e�9W҆Y�up��˩�SxM���i�Js��x߷��͆���V�
}%Ӯ�-�N�X�g��}\�>���1�H1�5@� C��L�������0I����#^��T�eÔ��b-|Q�h ���!��x�gR�Om-��϶����i��]" ��QΚ�9�2��)���y�)�7~t~����8�1�=UNoc�)���q���h|�$���_�-o��(�e�b�5�cN˖Էo�S��{ۉ�M�vgd��|a���~����Rj�5�mg�[�4[�>���Ge#�:����M��'�'N�Ƥ�m� ��	g��7j߾:zWL���b�nι��L��s�U]�=�n9q��P����kW	���Qi�C;��7':��آ�Wf�X�=׍�86q�ڛe4���b���� 0�~�XY���41��(V;��z{�P[='����:�L��ŭ�^w�wo�y�𔶗�ަ	yܰA��*���Q=h.����s�ނ��{ʄQ����.�E
Ȫ]��z9���P�(�-A8���;@�/� us��8DG_�mJ<� ݔ��R����x�i�8p� ���$�0+�y��d\(hT�f�f�ؿ6��|ԛ��?4��UU�K��f3�FT�j�շ8�E�/��~�#gx
ۧkEz�Cی{��N��g�,�	S�Tѿ"���	��G�O���� �4(�r=���Ŵݑ�[���+��լS�[:1�L���F�'��}�|}��9�r��>0+Z'�\���	��L�a2�83�6$�"-A@'��������ߵ���%z�-�#*��z�OSD����l>��\�h/�A>D�u��(��{w��������y��馽��>VX� X���zW&#�C��su�{\]Ѐ1?{�B�i�ާm��^����=���4��T�9�{�_����=�5��;���|9�G���cj�R��Cu./z�����wڷ�=�s�ѣyA��%� �z�ӎ����ٮ�'�1\��ۉ��=m�� 5X׫gzNrM{CxW=�V��v��v?b�B�ʣ���8yy���]�F�G��S��G���^*ގ�1�n�v`�<q��mz�T5g������ ��1�yk4�^�����ѣ�9�Y�l��βS��H�Z~�w����sU\���nO��R��dӝs�q_���ߞ����A�n)r���E4��`!��\�eAwm�wdoy�=6� p�zfBHg �5�f�<�t!� o��( I�q����O���#S����1P*j��b��v����M({�U��|=�������G��^���~�p H����,#;���;�$V�\eޫ��(<os�l6���ֺT�m�����7�4P�K��T�.;jd���f���.�[
�"�MT��p@����M���O��z�~�Ω�M�5�L�J�I:v��k&'Y�����2#�Q!q;8�=
�\��À ���9BtB� AR� ��`�s'tG%&���S[�$B����6�Ш�E(L*6�M�N)	l"�m�Yq�	H�4>w]������a����	H��K�=u�|~����}���|�\�^|������4�M�/N���z��՘f�&\�[s	=t�`%S�-��cw�pQo��+�|��g亩U���xhaͯ6:�g��r����C�ws��N� ���#܀�r�۽�lP�� @����g�5��ҮO�w��]��9
>�ps�A<���Nk��O��������w�-�b��άH#�a߇�G;�!����׆���=X�3My=�\���-�8��mo觯���,b$t�6���g�z��߾�^�%|�>g������z���q�`�W������+ %��ܣ1�b��鷞v�3��5U@�$�H6n%�RA^�>��,�8�� �����g~�&j�>�t�~�
��38:m���xO��d��x+��zڜs�U�0�,�W�����k�R.�f�6o{'On�t��%Z�ԨPA�$"%��'9��7
����p�|��G�\�If�h���ȉ�8�ԾS��R�{۵�I��ᮗ���TD~��:��ʄ�L�8ȭ����:��߸olwC��*�:�WNg.���stvO܂��:��Ռ�����P�事��ɕx�-�=�=�e|P�a�A$����+�
"~�*�zt2��NF��§���On�:�.ﰵ�����37��C���t�S���d�����O�����	 ��`t�1 ��>�{_�3�Ѯk�W7\�,лo���~<��E8�C�|
�5�+��۸�ѧ5���3rd̽»[��TF#�`���q��z�5|w>��6k��ij�}�>�jp����wW��A,�m�[�!��W.�"����tѿ7~Y�;�D<5|@Z^7�UOe@7��0��1.������ZS�\��" �̒.�	�!	�xc_b�����{��v詖�u.���넞����F�X��Exv*�0fn`��zkw�dW��� ֖���PNBę��Gx[
�8�y^�`׺,��߱�!'�8����{�o
�.�ո9s>�����pW�-C��QҐJ���Mx�Z�e��|� %<��
�b�K�glkj�����wit��=��B&p�?���=\�1؉Һ���o(g�pq-�h/�xԤ�����A߃�(�+��ol��߻���r5��6�ʳ�j�L0�-�sb��=|hU?���S���]��������c�ώ'��M,�x������~cE�|i|�|�bG�*(��c�䚮5��\�
�t.����aR��.h��6��ZJe��r��Jp�R�I�Us*e����n�U.���t�:<;^�˻WM{Ύ����5m8cxN�8�#�w�ס�&IG�ܩ}7��~�y��w���r�� �H0P�(`A����bC<=����AZ��N�a����dU�U>J�ͭ ���'L��X���5�ٜ����Gh�ce�_��cٷ�����z�6�z:5��ǽ�,5�A�:ʞ�<�@4x3&����q��AnQ|�g1o��uw��p������
ϯ�qc ��ho/g��J����{)���v�����9ׇ\�>ጘ.f��2&���j����L�tb !�.�*�|.Q#�t'�ҩ?NM�q�9�d�����mMQP@�PE�2A�7���k�bJ�W���O�o%d¸v��F�ƹ�4��-�k3*�c���v;�S�'���P��r���:�g�4�����{%����H��$wO�_R��n:�� xN��!#�����#�K�
e;^��Ȝ��Mi��ɰ��'|�y�,�p����u٦�R��okp�jok3s�e�o��e��w)0F"W��V�%L{�fѽ�}r3�]G{����9�����-G2��2Ǟ�E7R��v�:$Q�N_̆'�e -ԗ����s~f��
pǪF�@�c�?�Wt}h.�t:l�,%x�u���0ëdD����q(hgn��mW7�=4C:����0�c��=�t���-�X�/r���G��o��U�U�A��(���y��A۳y��aY2K;��g�a�u��5Ɗ�:�����Xs=}�rv�s����}���� ��y��-E5CB�*���������{҇�qQ��!}��+��!F��DL��� q�}J�i����z�z��hC8�z���w��e=�g)�t���՞3���~����V�C�=]E����q\v�����D>w�Z�]S���((��E`$�j/���s��|	��O�����%��:�4x�9�kS��n,=�m�t�W$+��؇��~3�Cgޏ9Z�����
�+۾�P���f/�g}��;�'�t-��3�am������41t��lz����e�j�>�n?�6���laq��a�_5���&�~��Zz1�,y]󯕜U���K�Aݐ���k��Y�/~�y��	>�15oH�o��ڇ:�3���S:7�����!a�e�hs.+�,&g�'����1!y�i�y�<��Q����J�ADx>���ˣ1z�'2���b遤E3�𳹿f%�s��ЇG�7e�!���~%��K��`5���_�;;�}�X���� M�������@�l�3�f�@�[w���L!;6�0Q"��0�[��SϨ�^F������yA�`����X�L��[���`4"�˺]����_yCX�-\���DUP }�".rUT>�DC.������7s���uyf^ή;���l��m-��NVŧ{�5SJ]W*��z����!Ƞ~� �
��`�U
��`�&n�5SI�¢(�� H����}���9��J	���H�aND�I3��2C"n
j"e����8�)��J����Ɵ�E>�Svq�ҟ�ė�o�O�媢o�|w�'�|OB���Yݾ��pOq�L�	~W�b���e�I%3���l���3(}��L���̺��zim��ަ����[G�y�\W����<KH�ۏ^��N�z}���k#j�̧�f����xSDtk �dCU�p(��}�g�:�Pяv	�p�)ab�E╀;���
����C��}l��σ�7T���g%�����ˮ����)����hcc�?\�Dڹ����,!�=�c����S�r���ֲ�ګ���:p -	��};+��T7O�"�5U������?P�5Oy��j'\����<c{��7�
�3����W�#XkHw��//D�w��Z�M�sr��ޙ~��;�A~a�����}k��qa�_=���p�py3�ܗ�o�����IY��ԢR����6��T�=���%�R����s�.�ښD�+;�{����f|J�޳�tv&����.��Ls��c43��s>�Mb�o<�^��}0Ȏqk�g��שg⧷V�R��&!����Mf�;[�9�T�-��KeYLky}��6nïi=�݃��j��u,�>YG�x����t\�:D'2�I���Q W7�QC�������!e�y���zU���蹔zlY�����5K`;Sp)��[}Zh��� xr
҆"� `��CBP
V*"�_?>��s9�������Z`�3���� H!�ew��.1p���/�/����A�7�%寞|�Vt?X����y >0�f12'Z��'6q\+��p�}L��2�瘟9�Nmn��v֞�m8�����>�ޔ���-�̼^���{�is2"�=��%�n<��;�=�!��xU0J���5�>�f��
t�ê��\���H�t3X��t�\���{��[�5}|R�6~(���7ºy�lės*~�ub�+�T��"\C;��q�"9���u��T[J�<�G��G�hق�΢n^WF^�ޕ<6.�ó��Sk��QK0nxz�Ǔݨ����@U����	]��'~caW�G�~ߢs�ǃ7� }�͍������_n��zہ�7��B�ӹh�W8a��r��W.\��"Ӊ��4���n��1�w����>���t= VP�z�+ÕE����b�$����*�����2���g:��{�xаH���f��E�u0�N41�<�ܪ�_U�b0��O���<-`[ɪ=3�*�5^Mm{}��mX�TV2w6���,TB��}�}y�յ4�v��VD��]�cf���[:��do�!�t�-�ꐒag���b�Vc�m�W�j���`ڪx������^�V�r]J�R�r�rhk1��W��+������7bH‌�E�:s%�ET�viw��Ě�>=�V۬��}z$=Y�Y��9���τ	d:���M�݈Pۡ�@���6�iإD�@�\8Ѭ�/z�f�5u��7��
���V+oVN� �7l��T�hG�J��Y��I[f��uɹ�8{agX�NU���;�,���c�\�iW����rP��4��%�"��V�@�����u+5��7�̜��W�E�����ֽ�ը������e�E��J�����Ξ5�>�OTA�����T��$fl�T)�@���oYp�wK��5[��FZ'ϻm���f
��3�r㋘]��']���s���Ãf������Ѕb��+z'�&�%`�j�^wi�]'G�\���R k���T�����!ՊB�B��zoe��6�&��&-��g��BӦ�l��](�k/P�x��r �����ՙ�#��<%�@əj��}k�����ъ��^�nG�v���hj�,��#튍B����)�	Bc�9ONb	f����{M*8D!+$�n�U��'�$�C粰��:���,�%�*d���q��h�;Dm���(�]�:{�x
�U�U�Z�O�UJ�x��z7/��R�|��	�f�f>[��"�r�j�M�6Nfw_h�G��z��Q�Ŧ�:���>�7R���3!�ya�4�
���]q�3iHj�p��U��$3���jwk��kT|�
�U#��V��)i..�n��[n
�hLy��b�u��a�rr�y�����&��M�#�VA[�G���[7wR����7۫q<�����6�@�Vnl�X��̭
u!77( #��F��m��]Nu��� �s�����p	�q�SO%�[U}%ՊFos��C7X��+i�bW�t�z�]��G����(�w;_LVF���R���u)���eD��C(�GS�dT}L���[�˼�y�x`�7�u��ϸ��I������n���W�pn�|j2���j��v�h96�-�,%�M�7���e*|�SV[c���hr�����Y�ˑΜ�(�)f�!\�U��@귕��n��`��e묥t��]��KJ�I5E�1G�;�b��8O]�̼�d7��rz�L8��$xPH�"��i�&S�aU�o[�t��O�?6�Ǐ�|�w�=�qТ{d}�"��XA�Tr�U���"����ݻi�ߟ�m�Ǐ��>i�N�B���R�j4_XQ:�I=�����*�.E���sm?>|��o<p|����@��}g}�y]'�8�JiTU�T�!��DO��wn޵�����m�x�����1�|PI!%B�T=$���ǔE9�D�E5	N�Ϙ��ƞ>|��o<pq������H�Dr�UVC��\H��H�#��"�+���iӶ�6���m�x�|��M>�Z^t*|eDW(/�%�?b_ �p�HQU�D_"r�D^q
��k���> ��Q�yYr�r��)P����<��r̎]�� �'PK_>yú%Ȣ���(.P��}׌dDUQOv��J)P��� �T>�
.�sA��l� ֽ)���j�*����<t��)
ޓS▞���J�<
�ʄ-ٯ���?���Q��P (b?�T541A ��@5C倠@�綧�to9�G���/�j]U޿������9N�黹IcK��ĺ�g���L��CW�G���qէćЮ�6<�6��q�"��'=���"�d�K �X�N�^�|f�wt[sP̀P`�5�¹���$A��[b���ߠ����G�届s5!ZA���y�I�8���X����L8	>��L���TSJ�������m�����.�!�R\(��vg�k`��y����gy�4�#w�dME�ہ�C��P_��֫����>�U��4Ĳn�tdy�ё��+^��3�}b��s�JT$Qp�3��f�0��\�-݆�}��o7EGkץ۟�@�ge�0�(݂�ua���O���虳V��U��f>��hgO�|�5�g�z��z����`3N��C�X�S�GQݽ�мs\��7��T���v�� ��v5�g ��yZE��~a�_k�C]���JHh�Ź���/+*b;����Y��@>��}ݚ�_mDE��Qcx�W��ȸ�p��AKuv#>�_7r����3%��&��3�N,#�H�W�^T��M��lB���c�	��h�j��k�ݒ{��9N�Q���7��}�>�����F��z�����o�;f�����uc]JG|���ˮ�#sܽ8�Rܼ�٭}/\?aV��@0 ���� �1  � �*�f��Lf�X(t���� <-.+�7�����}�D��%f�dN����Q��{�җaS�tGP����^@���<3@�,�y*���w\��ۧ��f��>zw���m��/��</��K؈w��j&�@��p�k�p
Y�
��>i���[sЦw���1L��+P]�n�f�=�{��{K'���/��l|C��\���(�Uu��|�"��ݠ�[q�L�]59ڍ��	d�;8׺��`�9_>
�LC��^���������6��}�x� E�������B�
�Z�@i�po<��ni�&���K����E�P���1�>c���}�����c�/̺��F��8��]73��@@��=4W%p���y��k����|�Y��m�;_wH��VǓ&�p��ϸ�����Üd���`��`,+m�dS!=�|�Qћ({ϯ�K�<���M�͔r||BE\M+;�`?�{�L P��!�;aU�����8�|SOĽp,H���]'��G��~M�P�`o�_�l�.b��皰u}U&��b9���&��������k[͋)�1]_M}(�c�5	ElE��wj�$��i�FlF�'�d�����_&}��oױ��E�Q���D��W3�������=���k�&�2�\��{��͆v���3y;�;���rUk�a�!
0a؂��C�(��*Ry�-}�����1�-�ِ'�S>�=N�8l�ƒ�� ��b"�)�"D�	�3���"!LC��p�!�G$��B��N����&:����g5}���{�8	�s�l���1�|�������O�����Ɉ���s�x� \���i�����p�֯�>sU�2���pB#����][؄�����<y��zA��ޮ��I�Ή��2 ��<���eU�.ݗ��Z3�
�65�;�>�a�&V�	*�/�͉�:���X��.����i����~���n�Y</���3�+�$��K~]�$E�I�f_5��=@�m{�{~X($|�Pj���3�Q�s�\cA�sws~�����%G�\�?4w9��g 3�M*4y~��i U{�"��@g�bv&��1�y�V�v_�nCfw92��	�11T�Ϙq�w��5�v=`�E��0����X�d_˖��[O���g�ˢ�A����L0[\-��;�ؼ{�����#}Sb�\�����3}9���b�����͞���	�Bۻ�KkϾ/<����*s3?7j�	��؆��	�p6E{�7�~[�z�n|��و��ef��1\�}ߣ<j����D�8�-�ge�gtw�c�zo{ڲg���*w��!Q#8u�䙶�UT�O�$R�K�"����1�E��u���~�_��j*1���CH1A������{󟕪�>� �yې�P3f;\��s��6.���ďR�A#��z��G���y���p?�<1��D��=��~\���]��ͧcX������6W�9�Ft^����O1O�|�E��|�\;��t=D>�̛/�ﾚD���f��]c���z�˵�g�N��sQ�Ϻ����&NU�QO���k�4xz��)�ط��Y�^'�y�O�����b!'l�����ݫσ�Y���и����d��=���cp,%�;��60Qk��p��0����r�}@M��z���������n#[���!%�W��aˢ~���}
��6�u	��G�E1c�:LaSr�u�B���f��G��l?rTȀ4�k>V(.!D ���*'���l�Ǡ
��a,g%����/�b�;����)�(<��əhQ�C����__����a�ܟV�]��ez$�=���;�6Yd0C,]j�|��.�I]���iJTG��*ֆ�;����;ɏ�gA�k�%}v突Ql�r��"/�������vZ��k��q�J�P����t�G̱��%����>U�Iu�>F�F�P��R�\��n��qCIHj}]�{���dq�8t|�Wċ�پ�WS���_j��L�[�`�J�OЁ"����A�hb��CH1E�3��x����d⟳��;c&�1�TMA�g�Y6l���W��!$
W~��	�{�N����y�� f��[?�����
�YA{��
�=ܤx-q#��]8X��ߐA��5�7����c���k~"��iⵝÿx���`�e
O���B��,Vq �$%���x}}�����穸~l���E8��C&6O��_4%2è7C(7����/:��:�:����@��&AIQH"��.#���|a���9���t	!)�CƊ����s�%�,L�?WP�r�n��5�J=����>aӮ�Hk��j`�L��������k�Y��/�M5G��"�n���1���s�& ��-����=�͐�_�[+�����LVd��lʐ���b3�X$;�_����(� d�����1�¯%Ը]T}��2���mh{����Y��{<_�7�o)C�c��^IP�)� ��h���3G�L��ݤlS����>t0P��Ы�:h<�#:��t�X��OQ�2 d3<w��Sݴ�e��<�����yy9iXV�E�}*��^_9y!E���*��EnW9^-�|$�w�5V��<5Z >�f3%��=���w���u��!i�C����q�g1�Z��
��{��a�S��y�?�����41P�`�@�P�+�O�5ޅ�W�fͮߵ2ua8���2y�C�!d5�\=����Q�:�5_i�j�k9�_<�3&�z{��2��ˎ����C]��z��K-�C3O�29@��y�|�	EA��X�;M�G�ǅ�q�]��F��S�dG�O�,�]��T5�� sWR��"�3���Ÿ6��Ӯ�ɩo;��c�ρ���4H
���}�.S���E���a�@��m��>�i�f�	�Ϙ?/��c�\MJ��<"4hZ|4���g%�,;��u��	G`'�@��\z �1W�nvlb���)����]�t��������O�-[��7Z0���<�ת��/ n������-�췞k����`�}	Il�y����n�0�k�����M���8�[�h���ξ�'L�g+��`<����

'�7��ucu%6� �qW�ۑ`����5�{$w��"�[S�S���WYM�x;�5#w���� �/���|�P6Gt�����f��d�B�|A��Q`"W��W�����"|�6��3�K�3�$uc3�	|��������h�#�J<ua�#���Q�AX�A����e���ͩ�s�\��:X��/���o�o�����TW�}���[�9�NQP�c0d=s;��9���� A��)���`�hb,��Dy�@��5u �	a�I1����~�}��5�H�iģH�HĈ�L�\0DD�b)�~�%*��H��bL�O?���@����
�|~�}�7��@y��|�� c���#'���XCv�Y�����|�[�Y��S`#�G��l�|����E��`�Ρ���>>ƽ��tOh>J��"�|�X�t�k�����o�������|�x��P�M㰹�w��D��Mz��A�);ǔ����'����fO|��=-6��Qӆթ�m��R�'}�J"[�hD���g�H�g���0/U���终��	'�[E^mL;@p{%�G�w>�V��l��� �M�L�A���� �H3�kx�z.�?�ѱB�]�s���}LP#N�џW&{�Av��Z�]3��3���K���Z��ti��G�(�Έ����
��íچ���	#Mw�}9�9g�2�W����R�f���=*��z�E��(�[	di'�}�Kbqrz��8����\s<(34{������A(�r$��i΋jǹ�S!=n仵3o@�࢈���$��-�H���ۑ�f5J�*�V�[�mGNO*�L-1qw{+T�yA�M�s�p�}8�k��7}x��F�1V@N�N2��e��hX�'cY��Н0H�
h�Q6�I9E�;xْ<[�rX�&�+77�Lp��o1v��q�����ݝ��/� �@?C`�@��@ ����<��-EJ��ߟ��x��?pX햓= �����
��<X�:�'R���3�����׋V�b�O]�>IO���wd��׳a��|�~�V�xg��d>���=_a�}�Y{�Z�]��%��!��KCv��/��Y��:���|�PC͖�	./_-/�͸�EB����<9���.}�y�0��u����ன��EÇ�u�ev�&�b)gcr�"��]r�v�8eB�n8�F�,�.{��p���M���I%c79y��Y{�~�4�*D���C�Jy�_O�i}�����S.� FG�Ǻ{m@f�ه�^�j�Yʊ�6�E�҇�����A��XK�2;�~/-��|�]�Ao	jc�M3��%�OV�3�����{o�v�rI�������kɜ�VsΆ�g�� Ԇ�i�!�GZ��z�E����"�i�RUkJQL���`�\�ف���r�6}��־�DU��j_-�^˼}f��{���6�����SC�B@�B��[;/���<k�gެ�����X��%��8R�il�X��*y�>���b���ީ���Κ:�IE�;so�mM��ȋ��^��N��*���w\ɱ>zo/m=��*�+ گ�b��$y�v�e�٪pZZ>?���C&2gL�vѝ��F�dh`�E	I�b�竿���;��
Ϡ�M�_�0��Z1;����ջ�JE_H����w�>�̆�}�:_ä���O8G�՟��;�fqO����+�·,ӝ!%i��Qב?v��z�}u�|��1�U���H>��D����_v�  �!����`�Wfc���ا]��\MC��*7�~����*�3�;0���`�K����{���P,\`� {A������}����#���MA��`a*͏:w��p�=�S���Q��}'ON���p��"E5[�[�n�Xv��n����X�����M(~��%�����3�����!�#�bFcb���ݜ�W.	���k»�r��<���q��w� �*����m�;d8h��tz=�����_H��ޑ;i�9��n�c��݅}#Q{��[�H'A�OǢ���T��O9����U��y�}�וb4o�x��s��(�q�;;^�נ�^c>���9�r����0��~���X�������[�(��d>��ǳ.썏g_��#��xl��Ya�2�gb�� x�����C֚ v��/��ԡ3u���9�{�����z��*?��sJ�\��ʖ�s���I�d�Y�:�?��0aP�(~@����2%B��2��b���x��w�*�����?1\��������%��?��TC}��� �ǵ34r���(�9y�fP�䤐_:�M�≏i�lflC`o�G�x7��M稛x�ǙNPf>�����}j�f��J-��A$�2�&;-ᡏ�l�z�l���� E%;�i��*1�`5���W9���9�y�a�2'
�����5/O0�yk�b����ls�3{�*v1�Ɣ�(H�P�%$kn��J���h������r���D�yaJ� �gU3��3w����Ks�V�������<{��@f�7Hfi�:���h�@Z{;����;���L�1�|��Z���B�
xYݯ��tg_,}�EyWcX�Fa�H�����xW{+r�=�%+�sN���wW���+���G�-�g�Rv�#��ާ l���M>��:��|=������^1-��^a8D�	��'X�5>��E���ǢD?�3ɚ�\a�p�sy�t-����ʌQp[��Qs����v���B�o.��S�]<�xx���F�^(�b\�~�m��ޯ��}���*�(���&t؛ۙ�dd�����k)h7^:�8�S2�Y)��r��y�|B���6�P��峇U����	�U�d�LGyH;��r��a�qT�knCKE�]���y�aab=F��o�Ԃ=�\�˗!L��`��zhز:k��9�&�̙m�Oe��&�h�ɪ�l�.ȵ�O0K���xP�-�ZL�"q;s��h�ٚѰ&N��%��ʍ����KĨ�J%Z-f��Whm6.���=���3(�1�%����VVZȬ@{�S�u��l8�;VP��GX�j�f_S�{�v����r�HB�k��t�G5�aF�m �fΥ7�gE���î��p��9I�bG++)`�.5kb��Y4Ŕ��=s�ܐ����zzl�K)^��w���^I�46��.�p]�hM�䟭vS���1����j�=.��d��q\�Z�����)5�]��I��s���.▍tN��5��N�� �oi�uu&��}}oX�Ne����%^�s��Fu;~�d����5��('^��\�cm�][�b�5�6mEP;��QO�ˢK��_n���e또����m�Xη�x$!����e7;3�T󔲮���W�e�کB��1rj��:rЇy�E>�X�]T8��>�q%j�-�S�R�R"~y��Џ�曗t��B����=�&o��)�L�̼�K{Y(��r��*>�ve��+{�ه#\�������Y�-�\���^�4X�Ĝ]�"���Z���̧�����՚�lE����Sz	�Ya�qɴ�&]R�r��%��U��&n��6E�U
�aa��tI#�h�$ΗS�L��V3���姆P�,�Nh6�}N�Ғb׽LP��e�ۮ�q�UF��>���|�Q�+ܯ��ܠ욓�\D�f2(�ۃ�c��_U
��]��¶�����|^cZr�)��.��a��]A]���j�!pv��%����5ƍ��[˾�|W^�N���X�z��G5;���u��y^��T�Q���,-�;�)�f�
U�w��7���m��#��;O��j��}��j���{�mh�w�}�n�b��*R��ϻ9�;��u�f�P�mw=|�����+mD:��.*�,��:R��_y��i�~��Y+�/�8��x�]/(����GY{�h�Xn��sA�P�[:�۽6MÊc}ӛ�̂\������/]�H6�M ��6怉�$��|yXE���?b]��I̪����t�ج����~7��c�M�t�����x�����|v�bȹ=�!�(TL�G":���(��U�ARu�t���o�?6�ǎ�>i���e˳��w@u��
"�t&��d�(.Tr"9t��o��Ӷ�>|����<z>|���> HH.�(�YU���r���t��*��r"��*�Qa$�Ϙ�Ӷ�>~x��o>>|�o���~���ʂ
"�-lYE�c��r*�$�$>|�N���?>x��o>|���~p�*
+���r�"T"�����B
9Dd��22[�4��n�>x��o>|���>�$"��Hd�FBQ���TTQG+�)�oQ8U��\�Q˕Qw�C�r���(�E�S�'D8r!�|�x�Ҩ�YW(�ED>�����*�#�W#�PG��Ϧ~�|:�9m�8�4��m����F�2H�A�`��n��đ������P3N%
b&mq��2p�"�)8���I(�A��@�&����	��;i.��Y�}��m�\�՜�<a��w��Do`�GBy׽�������;��r��ԏ�J�b����r���h4[HPB�4�q�KA4�8ʊEl dz(|�f�;���<{�)����0al�[)7%���qFT���rH[@�ƚB@�$�JD��c	7!<�҅G$q������(��p>"K($�I0	���W����D|����O2W�>1�ABF�N1$
>B���e"	1(�	�7��� C���Q(`�@(`�Nr����QDQ0��-4�L��H4]��l�K����#�R2J�I
%@��=w3�xܣ�Λ���������*%Ä諢z�k��>Na�n��G�]�@mOVb�k��q���b[�_jA��GuS\�kz�!�i�Hx���$�\S� ���U����+����iם�\�ֹ�Ul����RJ��^����]s�P\4����q�c]����LYh����٭��o�!�D,2���-�Oև~���M�Np�7[7��&�p��N��z���O�z-!�EO��ȹoUi���u='��v��zoK�N(gx��H�y`oq��[�-��n����-��D���k���n;��6oA�-�PP'�:�K~�9���8p?U{Hb���B)��?7�i<��UF��~9T����2�s�Ɂ��8{�z�Sb��v�	�0]���i�!�=֏r��_�[��=��?`_�ڲ�%~]-��?!�{Y��c�l���p���>���s��5�D�'"�|Dk<�c���[�S�/��l
�e�,UYU{{�/9�����h}��O����3N�4z<G�o�D>���U������.�y	��=1nG�N5�§�h����ܱ��^'mm��ע�V�`�:E��"�1T.��b����-�8WrCpR�b���S��+�9���:��5�v�ޔw�̝t�v3���e�bi�s��	�ɽ�#8��l��s�d�� =ݓ�Tp��f����kde3�m�5=��
���P�
�	`
z
��hnoG'�te�:�ڴ����Cp��e�� �SGy�A�-ŀF�;�>ݩC�π�6��`��C��Tjh�E���Dc��K|�S��,�����O�^�썎���mǯ�å$�4F���7�[�����(�⦰��Ġ�
�*���� 8�kdk��fxT���&UĿc\�Ъ;6�0�k��`н�O@O����)�N�����/"y�0L��Ţ��<���y {���b����|��DV��yh7�N����0}����c��0�HJ7�-%�}�ú�w�_c���[��t/������̈��¬�3��;�`�.�~|M�O����ϟ�^~%��!P)�9��q�Ex�s�^��<��;f��5�E����ͱ�l�U�mk�L�l8�k=y�a|�	��i��'f;\��{�����l%-ܶf� �|�f��r|���r�'
>9��
j�`V���~>=�����¿#@*������lμԂ�d�0|��"��[u�x�<���x� �˾fp��l�m�w�6,��|�W��Zzb�Sq��9���B++Cfzm�C��>���t�Kg�; �b@�5e�gs<<�\G��$%B���(���g~����>��g����]���w������?�C�o�H���i<)Uu�r����}��EҞ�ӗ>�i��ͮN�@���A�3�tV�]	�����#�M�~��'5sV��AH�����"� Su8*J��I�yٓ0a�,6'p�gTy�0��;�� r7�����Lb�q��Ukv���vhʦ֑��7����*5Ɓ���֊�}a[by����D��h�A(8BA8gSL4��yS�O����U�/qU/(�!$��T`��X�(��-tB{��P�o��v�V�]�LYk���?g!;���|�!CV���^�,�����	�.�s�g�BxwKk:�w��%:��ϾUZj�����4�i��v2e��cVsqU�a�}���}��$�Q'�KHK�D֞e�1P7^��t��;�Y�^��b>���H�X�ӹ{v���}ډ���
�p5z?�!�L��m����7hi�Z��22�E_����r�"��L]����D{����g����S���T
��{�^N"J�]�J���6�kT��'<��x���)����E�N�;��ъ���u�����G����C>����(4ƽ�f�M�С����Hb[���Ht�j�
ռ�^Ώ��6s�m\œ3��Ϸ�ݓ��Z���C��41H5D����T'HT*)z������K�Q�׺�����v|`ϴv�-=��"��F��������fK�4�W&����_x�ٮp��{��bC�� ��@,�_}�������x�����4<���|�ԣ݌��5l�V�_r.�d�*E�n٦�%j���H�%$Id@x/Ӈ�����R�Y�$W)t_>_ΰ�;��k&���պ�ͭR�7��Ս��o�^������w���45��pv�����M�'��L�4���G����_/��n�3L(�Ǩ>�0ĜE����I��L�ôQ!w���߾�D�۲ڽ���SA�w�`�C�w�=�{�#�^���]����n1��/�l�@υT�m�:Z��5���Io?zb/���FAob�������luN0���U��x5�B�99����>0?0�X|g�p��"�����gX����I�<b�(���ꏾ�����-��<�!G}�<j���9j��~�Q3�!G�`pS��6�3\OZI�{�OSm!�b�Z�.`�w��;�4O��T1A�2�r��﫠*vl��K���%�ճ�Ğ۴+Ou�×�t]�����S���⧞��I3 �z�!�s�>�b���/�Ýùq�\/����a�&(��LdO����Ufc�㦫n�����¦���D���bA�@M�.q�b��[�q($@���h�".z���wԨ�S!���	�d���L� r@�d)�"E̂0B���q��32y��Y:��apx?zq�����,	3��W:Dk|�q�y������>Öo����,��t0!�wgRw;�I0�Dh=p�4C�s�tn�<�^c���f){���`ڟFp��ۏA�}Y氕�Ö�{g�ڲ��:��t�Llq�A��Λ�"�	S�7%3j�U'���!{h>���ȕ*<]+*���K��I�Z-�od�/��8��e�T�<!%�H3ol|Xu=tXK���`�������t�u�����TD��0��M]݋׬/�S��qB�k+����H.��.��0���n��J��F�ї۝E�;��� �����\�{�gʹ�n��?b���ʢ����Y�|2nc��t�(.�7��,����ú{\V����������*�O�su��/���!������H�L�X;�,�;�
�E$�C�H��pٿ
���_� �z����l��B�2J4����%��k�𛧒�Z�D?O��/}�{[!ﰏNs�]�h(I,{ʵa���C�*��z_���� d{��z5�1_Qr��z�&pW�q�ϐj��9υ������i�/V��q��{����g��^���n��RO$�c�/s���˛�
�6ַ)Z��w>�����.#�p�J��M��	f�N���Q���L�|�<����U ¡3=����I?OꍓU��i����	��B!�Y��������9��SO�����Q=-ܚ�v����_�����(���}d��~׾y��g�O��F���+7z�s�������ǳ��w�D�g���p��\/7N'���](v�<託�D�����(�=o���1�9��8��{<��k��}�a�!�B�M�8�٪6˾��MW=�O�y�\#9�b@{�E�|luzi-��P�0+9|T�6�Y�̛{qZ�V�l���$��"jm��-�2@�wj�����;0-3�*6�@C��o(S'�x wo:�Y�hc;�Ht�M�����叆�j�)�ʹl6R�kk=t&f-�!&j��X�)j��w��W����OD�\�(��SȪ�疡�40|�O�ދښ�ܯ�W�c뜢v���
���gH8�P����fr�k�s[{rFd��*c���Wj�;u��;8�i�_>v��.�߽0��x��n�S3SP@���W<��;-����&I$ף�͌8h����6��М�t�Z�'�|��z�X|8_R�{|>T!��"��
W��x,g�y4_5��+���:��=��a��0.�����6�e�:�p�^3�J�4�\��u�?��)w���ù=�e~g�+D�z��A����ǎڙ���[� �������>=S^��czd3�У������%�oG�T�CO��M5�7�j�Y��su����E�����0V�%�@��r�P��vg�x�XF����W���l?k��\��Ǥ�����w�̟w��S��,�H���0ć_��D�{+=������+����r��1���7�ߗ����DʔhBSh$�i�d����ɂUk�ŗ����dy?� �����4xf�=�'Z�rn=Y���}�V�Myłm������o�Z�!��>�	A�\j�T�]pq/e�.�7u�%���#=CL�q�`Km8JAU��J%�bv��%�K�v��������f�M������9� 3 ������
�T�cW�a���:�X;��ބ���wwLWMS�~]��y�����!i���F�<~��.�n���܃�h.�l�}���Ž,9�FzXw<��PxX_z�BWo�dW�~V��4_)wP�	q+�=!���9I)�j�w�5̫����$�����˨}�iܼ[�l݌��8�]����V��ѯ��s�����/mH*w3�Az�*]3t֙�&�U�S��fnŰ7}N����N�8U8�fM�
*����?�8�<#�8� |D.����{K��o��͟Lc��]����i��H�F�s�M������ �gi~G��lD=aKi�T/�;p���l�N�>&ZU�]��m�=S�]�w�(E��s��mٹ��}�#��&آP"�iC" ��$�YH�F��.�?Bȉ��������vUY��m��A<���iF>��ɉS�Ҕ_=����%������X�{(.��q[۔�$�Nl��JC:2��!\[�_z��O���x��N>,����ϟz
�(���������}��ƺ>^HQ9�D���H���-����ƻ�����|m�Nh�K�����Y��`����x��(|E%�њ�>�Vt|[P;�[l�����&�__�����Y0o�d^�����H=��W���o��uZM�1/�D�9�?)Wr�U�Eoa�V�'Iă\�Z����`i��-��=0��gƹQr���Պ�92vދ|�QB�2�.+�s�7��qu�B�u�<0n*;���e�X�G���.4.�n�$]Q>�)Δ�y��Y�ؼv�ݎv�v�Z��rV�;��Ƞ�Mq�v\\5�����q���^ɇ!l��V���Y]5L�����ܐ�d�j��]/6�)���a��v]�._|f�M���?��5R�A�`A��B���)1n�
F�R'�(Ib=���݇tS��P�фR�E��D(`�Á##"6�@@��M0�)��
�y��]����>�`�B�i?>>���=�?{�����*�=0\[Z���������#�6���}�
�|�"5�k�WP��<|���k��{�0L�-�|9�ft^r���ZJ�{��@P Ԇa��o̤C?���R>VE�����9�lY�pR�~��qT�Z��������OW3*�`,k�<�#�Kؼua�D�M� ����:9P��}0]-��<p����<zݙ5�}��Ϊ\GWZ<X�cp�p�Ji�y��v�v늞��<���&�o�7z�C�����H�A�0o,R���7N�uٰ�x���ۄ�u��2��4��Θ<�	�WP���xeAszG��]6�}�
y�O"R�6e_z�N�X�Եz��o�'�
�6��%��g[\���;����a��IM���d�������)Ud�W�` |j��R��/{���Q>�&�����4<�4VG�μz�ca�]�\�孮�E_&6�^YHJ�ϜP]$^4g;�W�D�w��o���5��ɚ/����I���K
׭�r'o��,GY��#��f�QJ��sf٠ ��� �������x�@��#�xL�It��3b�^�����9�X����Hֺ�<|L@�Uwk�o2��c/^��к�щ ������ ��3��y����:�x�sji�G\��樂j���j��y���1�nC��JUH�����M\%�s��n��5"�F'�k�>�.��Щ��oj��L
!��1�S[5�]�i���ctl7�����t���|.�f����?1ޯy]q8����b�]M;��/gf�!��;�<y�6w�"뿠�
�W&�����ӝ�?�������_kmó&�ϔn/ᡢ���S�ᤃ���t�� ?B6&|�s/nF�봤��X����]V�����zbH#wW�s�g���R:}V_�Y�󷏇�\~���;ğpG�P-�LD>{~[����F��~�����Z(o]qu�V���5�B1�x����.����e����ja����.C(����w�[�wa ���1�|�<��ygM@�z����zۥ���4��:�R�zx[5�z�~��5�b�ǅ��궽Gf燡�ߎ���W���u,�Lzǃ���^NCD���o`���X�$i{��'������Vrؾm�"��a�f�ų���RT̍��'@wrm�G�������̬�c"#S+��{��Ѥw�^\�� ��V6X��ce����%Σ�T� �1]wVB��q�Ʀ5Pb�Y}�˳����u�>�J����Ŝ��ku�͇x�+(�VK��:�
��#�����Jƴ-��*Dͫ��[����{o5��/e�]�C.�ڷk!r���\!�����;��ϻ�e�ٽꀌ7�Q�Ǖ��S�w
I��̥|&�L���+Lк�s���%�F���Gx֓WXF���{w0�j���脝��[��W��x�v�D���|�^�a���c�)�Mmv�PA�q�jm�](�L�hHm�0e	sM��3�����kξy7v�Ҝ���q���(���:�ww&�����\�;.[,R�.�)��Kg�S�B�@����k_mғ,!|p�����v#9���bp���inW7^��Fa̷x�.F�1��wu�]r�&	���Y�B7�*v!�����G�7[w\Kܸ9�V�DY��u8�-�\w�q[sK؅��{�W���`��X�s�Y�j�Ϭ�i��:f�5#Y�;�5��[V��cK���@3d7V�&0Cf���~��j�_�-7,���~o�C?v_���&�Ɗ"ݤբ�*�aH��".�b�}���j����� ���h2z�ڪ�5X��-Y���z��J"{ucV�|��5��Ix�C���?#N�K��Y�o{}�zv���B()Z�5�� ڵB��=F�������D�"��:$���y��b��Ö1���;��T�O��c�l��*�%���\S^v@!e-�/0�&��RYfW5�,"q��F�w,�q[�l,���P�.�xu�H�B�2��8E�iN�=Ej0Ǧ#�"k��qO~��� �uܶ�U�9�{����8Z�x��g>��04�F����S�s:�y��B�qL=z��ڮ���h�Lq["�\�c���j�*u:�1�<JwVb�1�(Í��VT�>�+B&�uH��I��l�c�z���KHXx#6A��@�V�ŷa����	=��^&�R/3n5N��b�����P���dΌ`Ȣ�W��w�j�VX�Γ�v����*⨆��_m�R�I���6'V�,��[��Wz0�}��Х��[���ji�)�Mx��]����W6�jpc��p��Pѫm'�D�u.cw��:��P��|Yȍ��]�;KhIC;�l���9ň���'e���}�t�ƫ/@g[\ˬBs� 
�B�DW�
����W*dG8\">���(�����7�η���{�~x��m�p|���}�I5*@�2
���{���)!*���U\<�9@\������m�m����m���|�=!U��9��p.r}v;�c�0��O�|�N�??;|���m�|>|�σ��5�c�RI! ���QE9$DDG9�Y�Y�Fj��>c���?;|���m�[�o�߷��Q_q"��UșE��o��"� |��ӷ��;|���m�|>|�ϓ�u!��
fo�Ҋ���!�,�����e�YO�����=~|��ǏͶ����>|x��#�N�c ���i\�/����&s�%\��9�3�.vPDD�۫"�
eT���N2�L��-g*�\�PS(/��Jui��A�P}wc�|��U@�n��U�Uv�B9�YEUEȈ�L���غ�ڹ[��ꊴ1m�Ef�Fe�>�Huui��>}�-G��K��?�����j7Dd�k��g�c��~�'4���o�X���>U'Ȩ��q�t�g�P��$��{�}�is��ƞ���;��z�v�?y��)qN;���"*92{��y*&U=T�&�63�a��m�Qp%�*��oj$�@_iY�3�uĬ�?zľhMll~�ϤøjS{���<�b��ݏ\�@f���=j|�Ǻ�3��ڭ����/�a���s���v��G�IRˤ���̕�A�W}�+�� �
��c��܈YB��i��7YO��x��V��Sf�^q��`jc���j4TK�5˫�f�H]a=cҲ�sH��.|����As�N)�y�B����逽��r���&�'e�A��(C��>�4{��.WVG'�U��zR"o�Ϸ�C?v�)��O?~cD?6i�	��='L�w��VT��ŉo�{�G��=�x߳�N;����ă`h����}O����M[��i��s���U<'��0�Oly���gX�t��G`~�����~�Ps�����^pZ�N\�ǧp��W9'FY��Q���u.�v�y7+���Ɩf�mj�Յ'���F��#��߯���w)lK�Cr�*2����e�k�w�[��ڬ��+W.�͖�	rʕ)ӫr��t�i�߀��#�������w=u�zxrП�i�F'\��H��bU���y���4��-�p{yv�n�$���D�~���D0[��������>�0Xfq�Н=~������϶�XFې �L��=G�(^��&�������B��}�~�N��r�uƆج�M������Y�Z��O���꤯9�pa5��<2�ҏ}��0��Ulfr��	�N�����{����z&K�<+}�Y�{��WQ�b�\���GT��F��Zv���E�g.d�Z���$w�{N$�7e���c���`�7G�Q��n������K���y��OC��ˤ?P"=���3���Xl�v�$�1��M�/�.�s��N^d�Y����O���7�}ns����t��g��
�un��ۗa�M-����S�� ���\�G�J͆����8��ݝ0u��Y>��?�������6���eaS�Ê�Ȁ�X�y�����f�8׎Kc��K�yAǬ��󸫺�S������Ǽ��vÕ�R�s*Pޚ���v(�}	��,]��ɼ�vb۠�!ZP⦗�]]�r��J^���C�m]r���Υfoʥ��)κz���Oq�9������[���:���4���As��ʗն����?B8�A��G	,w��)�A
Ui�m!
�AQw���{��7n*%"̉(��Fi���T����|5�ݗR�Iģp�
a��I2���qv��Ͽˡ�)��������&PC���.������63߆g9�z���fh��q<�tt���;)�Hl(b\�R�t�9��hs�\���H�{	8��������o�{ք�CtO��Bl�&�����=Fٺ�#'�hy�Vz�^��%���8�q��'�qu�Іc�z�k�Oug5���'t��H�� �%?yF�'�y�z��|�Wh'���U)V�5m�L�&�m��^�R�'`�@���C�e>5`�Ζh�?������k=�Q~\�f��UŻn#�H�i�5�0���s�g��p<~�Q,"r㳴<�����K�VV�'����X��
zo'�����EI3��S��.f�	���F���U��;#��rI��}��2���4`f�h��?�ӆ_d���B�X��m�oO��a��@���������L�OU���]wPZ'ּ� �+�t��h���C�0N~��ք�Ե�樴-f�!��l~�ɼ,Y0�X�`vjX�-GW�B�|�W펳z�SX� ��	qN>���K�����VK��O.���y՘�΢eۗS��FsV��T���&){�����#���A8�5������S�?ʾ���b�������X�'�T���<Ͱ�͛e*T�Җ�:C����,z�"Vvտ��!XR74ӷs��ݛy�*�UGQ�>�U�4qR�L�CMP�1a��}iKE�M�Y9�ٳ)@	H6��<���u�U���h�۲�$�n��i˪�P��% l^yu���J�]�3�.n�'�m�� �}��RL�o:m�V�be��+�}��S׵���{��t�x0J�s�������gd�M�`�@-5��ړ�ᯯ���{��w0=.s$%�}76�%SQv�f��O�}ʖ��H5���"�(�Wx����mi��׻���:�ŦX��^R%O��2��������uI�{3���y���fcv_�ofǌ�?���%KL/G�3rG�6<�vϫ�
��4h�o�/�M�����!*G�z6�T�K�7���#Y@�B�mߒ ������|��a�Aߪ.>&�KJ/Ww��Em;l�b<���u�^��6*=i�+%[�Z6N��c��->'F�X:,�ۍ�����8a�w� ��y��6j�+���}��=^�ʗ�{/��7o`��~��I�p�����]�?����Q}���}|CH���k��ϭ�8zҀca�A����oo�eICvm��{���)߇����qS߰��4����w�+j��yJ���0i�*�gǢ��~'��؛��U����D�V����X����|�����30jP�d,'���A!-8r�G�x`F y�z��p���5SU��c9�`��
9��w�Y�]��}FI/��V��"���q�>L���a�Pp�����[��2���� Rhrɑ!e�Φ�}wm���{6n��f�=h�&*7ݽr�qy	�;3���t��S�v�w�m>���4:�lE�MVf*����^(G����X���`jUc�l��t�M`_W�Uz�_j��L]��Y�o�y��7�O�lUx��q˶}�zLve^� l;�hQZ+b�ǌk�Y�[���m���Fe���]��Ѩ��u��,�}V���'p���l��/��G�`�tx:�WwM�oUv���wb��G��qn��w�[��76���y����m���X��u��gs����� �2�h���~~o��ޜ��9�[Ĉp�:�}?�N�G�FGfݻ�<�r#o����kS/�oQ�Ht��l�|�ހf�B^�{2놆Uݹ�w4�A<�D�
M�?�����UދU^��aڲ�}\fpIZ6;3S"������W��,��J[~>��B�$�r�+�  wE�E�������׽�j]�`f�L��;`+�X��Kֱz\�C7��#3�:����.l�\��0�e�)���W��i��e���W�^�@��/d�p�{0;�P�U�0�3f�b�lű91S���Nqԋ>@Vk�/�K�{l�8x��Z�]b�Y�]�zy�R/3����{��9`� o(;>^���z��6CZ�H�\�F���DWM�u�ʻ�JZ�(h�"=W�N�Y4�+e��kj��e���V��/�׵X���i�7W؍�C������[���r�T�����Kn\[y�M�>�*`�B>�0��@�y�[���u�p�T��r�n7;	�W��eT\��2�m����.fI��(*��^ �<H�ɉ�B�GŖS�f��}��i�0:@�cb(�D��K����]��x���n���;��7�g*jx��50g�
C{���Mҹ�r�c8��S<w����z��O�o�2�)Z��5���q57M3���xn@�xcǮ����'r1�V�u�[����t�.םsf�m��m�U\��0 ,m�#�e	�3�4���g�&��骽fvn�vV����6\���%U|U[ɩ��?Jx�f��clI�(��7ssN���^t�{�Ni�=�ˏy_vԈ�q�$��l�}��s�b���:��$�����fX�못ڵ�8wVHW���ت�ד¹��d�.�wilv篣;Nz�t�δ�Z�[i��'`x vs���h��Ke;m�Q�
e(��y{���:�.����8`�FwX����*����)�aT*zY��oEyz��86
ie~�BZl��M����7��@i��W�'��ȍ��⸮���X%)����J�5Ո��ΞIc~�z~��G83m[�U��Ҋ:5�@��j�v�p)n��3:�2u�o^�w�@��d��+�-d�q��R����x�<C �y��h�H�^�M_F�&�[H�8�"Z���;V`L�r ���"�������1��e�{t�E��f6�3���]=���P�M=��Ynn�cAꮳ�,�������\�}Rm��
�}}%���4yJ*w|/ʨ�]�Ю�B��d������d3<Zϋ�(HL0�������%�R�x�u��f��~����̍h都.���#����q�1Hg���3�i�yÕ�zB�2�! 
,�I�C{���_urɑ�Y�ѽT.�25=�W��z���f��),�ʮ�7�չ��=�-��k��ֽ�ʃ?�=P�-�M˷:�*7��zG,X���IW-�I[����k��1�����Oݒe��%��->�S>�=��oaqM��xǇA����������m��w�3$dP���/W��T5`o�?\�v/R�����g�d�"}{������	�U��c}��r[{�t�Z���ç�bo+sdi����u�2�T�U��[�y�Ř��N�d�!��y��`<�Y�N.��r�3!Nh�}j{r��(w9�S��ԙ`���W��F[6���T�.�m��$��3ԛ�쯚�s�:͑ѭ]�N���S�B���ޛ�;���rګ܊�h<�˴��-C�����Q��օ@���rN�.sL�z�ON�X%�}�3rk��1�r��PH�����G�h��P6I���A$��G�4��Mh$W����y�;%����)��O�����-�m7t�gx]�8��!m?�g�T6u�Y��R�q��x�7����f�LQ/�Xf53��_*�={�Ĭ�M�V6H�^󦖪̈�y�[G��3�|�{d��FǓ��Wy{���O�q&hE�p��fz��j�#��pݦ$g3ų2׳�U>��g(�Ԏ���=9�EѽdW{dv󊐕�kS����J�����ow����'��wr�T�l�H<��3�)h��Q7Τ_=���BXU"�����~�ʵ>
d�YDb(xQ��C��ꠍ)bn��ѼZ\NFT��.�v��E�n�1�z7�9+7�s��}W�!;�+{0]Ɏs��͇��<=�L8�ڴ����V8�+���WL��ߚ����:K�c���1/'�z�3ǧ��,�|��
u�����`#=b����m7[gPjy>޽����HH2Jh�j�m����oP�5�|�� ���{G`W�Ƈc�9&g���D������C[���C����Sz;#�1�c��$ՙ�y�:e)`n���4�ﭠ5��}�7[�W����;�O^#�N�<�hf���e�v����k�Y�Ѕ��j�`c����'P�}�֧�+��h�vYj�q��Ƀ3XP���x��M�r47f�('mz�*�F-�Y�9� ��Ɇ��e�D��1Q�^�h$�|��/�8`���>���\�pƳ�w��3Ϳ���	Q���J�=��D�R�3��C�E�Pwa�F�U�oH�ݗ�Q�g�����(a������{�Fb�cx����4��Ք��n���(��@g� [V'
m�Lg)7"����3�eV�#Hkx�>�Q�l��f�O���n�\[u\ٹZ�Xۼ�r�E�1��'�ҕ4��C3F�ƦC�*��޴����c�o6�Q#2���6�����ze.]b�x�]�:<�9n�$���mw�o�����x�|�ݲ��i�pت�9>��Y,���h���a6O5��=%B��q��Y�➒S�����)SnT�n��T�m�%O2�Fٵ]ji!˴W���[��9�.����ԝo"įe��1�i�A�Yy���D/,�w�� fȺ���✶q��wZuf�{��z%�I ;&u����LOvL5����yOd�&�Vvٝ�
��x%�_8�A�G;rRN��uV���,Q�6\HA(P�fB�J*�����J�be�ꛋ�R���n�Y��԰$�H;�lwR������DVi�$8K�.�[K����Э�r��z�E�u�sԳ��s�J�>���c���pl����۩��^u��f��N*G�yp����F4t�+�M�
=ޞ��Y�y�N�s��AX�f��X�R��r��b�D�9���آ�_X�d"��)G?,�,5 �܌ZTx�oT��q��dΧxأ�� �XIP�%R˲���ɭ�eѾ�0C�{md
�±��뺖�f(��B���%�ڕY���8*��(9
�T�\�YJ�e��\�#�����<ҏ+�]u�"@���#82���E&&�#�Ҭ��w��t;�z�2<$���7獺�Sv)���9�h����ƅ��jS��u1��M�ԏ�q���5���Sq]K�_��;H��SNr.�+�(.����k�ZK�:9�n�w^ڴ�P�ǂ�K�J�+���aחR��ڊ$��
9ʴ`�X%��[��U�WT��խR�����clN7�2e���Pc���fκ�[���u�Gru�'yl�CMmX�ھA ���y�e��Ѩ���V�(wwr38�sO�q�s�K��V��_rɝ�۰�Q]��l��mfr���ԇ:��l���7A�3�K� M�I�y8�=�왥�ùq�D'D��9�����L�C���GK!"r+��}��f��/Y[ذ6��Ǽ΂7��F	���-Q���Ɉ,o霜�^^v)xZ�y�A5����_[:�@�.;0g,��w5+{3rm�l�HK)��  R"�|dP�.�˔��\*"������k��v�~����<x��o�1�	*�d�5�EAQ���g
(#�UXr��B$K|�ӷ��>x�����p|���>��U$a'��ʌ��:L��#��E"�.ADQ_\Y�N��Dv�}�۶ߟ=|��ǏͶ���9�A��Ҝ��ˁA��Q�޶���.�O��U"��w�������nݻm�����|��$�T(��(�Mi\".T+�y#���51����Rrw{z�O���nݻm��1̒2�BO@*	�9�P�QT\�N
������ӌt����nݻm��1́HB@�H1�(
9I"(*�U\}dW*�t���ّr�t>�aA���r�U�"�EPr(��,�Ѭ����L�#���|}3�E��r��UE��X�(�G.s�b<'�t|���t�
�7U#|%"DG����޽q�g�x�[�q<>=/t�!$o�	"�eq		�,�1��!�R4�,�2Q:X��X�Z���y+��u{s���\�5�(Ҁ[J��y��[���m��j�:t��^gqH�)���B�a�̀�C(�@�8�j���lLR)3{N�)�S�)�L�Jf0�A3��`��O��R�\I��a����z�)w�z�d�W��������	th��J �F"�|0���,(bH&�.3��2K4Pn�E�!E$� ��)"A(B�[�Cv��Ä� H����T����l��� i��{So_�F��0�"��"A(�@dM��|J2�fc��D!\�xQa�H���b3� {��c���Ь����l�g�Hn�5d��X�t�8�oT�%��SF�f�sD�T�,�ع{g����du�֥2�Gy���O��0}�vY_�6�p��KQd�
VĜ���3U��]��w����_���X���4M��X�=�:H6R��A����P�]!W�Y���'�&�����!b��ɴy�6*��[��z���ft�O5�쾰�J�)JW^�+�~�c#��J��Z�"+v���0�c
���}�Uj��Jӛc����nc�W�4�Wh{�ݴ���Z�zHf+7�
�
�#YaM���'�{�	N����g���:x�*bd&
���=x���W=C��3O����jf7�͝�T$�����/4ș�[����c�g/��{�?<���i�63��s-��0q�3�ņX��-z5��̳&l�z�k>�ⱽ��t�jn�:�u*��:3[�W_u����*�ᓆ󃔺퓭L�SG9@Sͬ�W4��|���7��0ߡ��o]w�m�H���rϖ����W�q����[;��:Z�s�L���wR�@��æ�v�3:�$�γe�K���]�s��)�fK�����Glf�3��sXF��\3
ӳb�+l+�L!��d��>��`)�4�}�~�����Y�r��W9��[������0\�H�-c&e���@<j=���[O�n���u���:��2#!����ƾ_}U���~տG:�
�F�&�KW���Sb����Jm9@������d2�3��B{6:�r1��y� ��g��L �/@Q؄yӝ.ϣ:ojk4��1�Vpx���+�������3��s�|��7�0��
������a���=�c�L��5#��V�<�\&��߬j+;;Q�0�f(���v[�6�V*y>����Dp��(<�o���`0N_7qB3�ܓ)�x��[\FJP��w��N,�}ת,ع���:<�h�Fe$�9�Wx��Am�7��̛�׽s�����ۣ�z�w���=M���x����!u�v�CQ��8n�?S"��A�߽o1=�c��z5М^O��μQJhʞW|��6�c�j^��(��*rM��q�y�C�����@��d��K%\�u*�͍rT���z+�a�}"�}�˸�/�Ȩ4k˻p����]��vХw�r���dB��|�S�0ܞ�	3��~Ƽ����+y������-���q;~��܊��UX�gF浔Ɯ�ב�^��ۖ�\\�d��{ҙ�Yɽ)"Yp�&�ag��KK����':�-z�����j5/�A#���1����-Q��W�6/�@�}T:-�f��-ve�F����$�=�79d{>�y�c���<�n�ҴZ�����ل�K34�
X���+ꄺ��T�����w.��Ϲ�ۯ����(���@��7UOǱ3���fD��D��Fw�	��Z*:��9%�y�����.vB
TOusy�-���o4m�#������=��͛۝s�a/'CJ���$�e�惐m��ï1a�>v y0�N��FyĻ[?�Q�5�vl6#��5�jQ���VT\�Z6&yƔ�]���<=�ǫ�F&�4�^�v�������������-�M�<i�Cĳ<N�A{�GJޖV(��R$�]�o|�D��Q-������v�,v��\V���:��������CR�f�_[TNfv�m5'9K�_z�p���26jv�,��ݶ�T�~�[��&�r/���epO�w���fݜY�ƻ�jMr��@L��ٯE����GV3��sP���Z��J�X,f:
��2��w7"�P�h�ޥoQ�
���lȜ�%����	�v��w�cӹ��,�;��h�Q�瓷�'��h�O;�&��0�B/��8�6f�Y����;����=�E��×�8�m�=6�].r}�1M	�^�p��z�9�[֐�����]��۷䄋Ȧ<�9i��`��v��&K��w�ۄ����Pnjj�f��*W �K꬇]�>� �Y��O	Ռ^�t*ދ�ڒ;���M�S��ß�8s�[�!A���H�"b�)��������a-C,�i���c�$��L�RH9!���p��e�8��\�4�%8�$N~a]6�����s8�T��m�����y�vT�F��3�5�Y)F�[�VzA�n�q+b(>�l�j4��Og��TX��m�?��_�d�:��b=Y��褲���4g"�y3]�3H/s�K	�Ϙ�l:s(���=��Tܹwc��a�S��T����_�6FH�}0$�k�dGG�淏Wד�G���b�qJ[iA��#7{��!M��V*�����n��{�L���)��̐�ȴҏWwh�wvg_��#M����;���[��^Zlv}R�&s2L!]t-=s=s8D?��%��4�6���#��Y�?	g�ĉ�R�|0��e�@ē���@�r���~��s�U]o�����C�Ƀؕvt��M�ژ���-p�Pغ^ �%@���z�����ġ��L-W�����ʊ��z��M�h�2�KX�oz����X�qaso��i�P�u�2�y��D"�m����'�T:̊��.��z2�^N�n`w��'D��ш�of�����3�j����_��#ď��@���Y#��#�3,߾�;��e���`�0myG���]�֗����GrR���]������7u��q���C6���_c��OJa�M� �p9%�����	\��^p]g�;�eKd���ͻ���5���ڊ�v�@C �ʀ��һ�2g�Gv��gTs�j��Og7�3��*B�ІCh�x؞��&���&��a�缢)��{co�,�r��
��?TՌq�'b� gi�����6�������K{��?��� 	�A�t���`�X�v��j���<�5�U���	~�~�����N~���g�g�Pb陙�36��G�ίp\�/V�8<ݬ�I��k3I��+�L� ��썝,�1۔>q�QL��@����V�b6 <w.�5��Ӿ��0Ƕ��,dG���Ƚe�үӴ�;kNz�RdP����e�h�~%���"TW-L�:��JߎS�{�B=t��^ہ�uk�6� 	��:&Ag̊n\:��r�u;xL���T�k=o&�-���<�E{ռ�ѺZ
룊gv�&��(�߀�Z$y�?����{)����v�τ,3b�.��`t��@q� f�1mi�v�u������wS���g��i���UPL5_��/��\Ʉ��{��o3Pm��z�1�����}o�ɏ�+�*y�w]Z�ʾ�
�])g��緗�\y��+�=�U����}�U�������\!���	6s�XU����9�c�B�;6^�KV����i��z�{��#��3��Gg*��.�6���,���nr�FM�$�!��"*Q��IUJ���vJ��w���ƬS��d
��`��7 ���=����=�K�:h��'ώ{�n�h��ƁD�5)��Ș���_�g�����vn��y;��9aZ3��֮�F	뒙�&��0���r����I�����&�w���4���("\f�d��zAI��vb@�SU��n�ַ�Ｆ�W7�Ot�.]����ٵHxz��r�^�� �v�j�{[M�8_=�'N*���Sݹ{�nvr
b�qA��Z�DgG��(�%�s χ ���횳|B���^M��3W��Q.����޲�2"Z�N�u�gsb����:�sL1"�S>���^Sc5\�I9cKV�m���Co��{*|�JL���.Ş@�j�`�B4�������׿������lk6s�}�o��D6�Hz��ni��#��k=��q'Q`r��Vctl2�4��m 3-��h��U���ʶ�ot�`W=��mSMUնr�8���z\��k�b�8��\��}W����g��A[K�כ}:����i���n�Jj�z&e0�Xgj�I�Ө �)m��X
	*���JV�5�nt�o,d�ki-r�OC��2�f.mw;	J�TVUym��6��C�_$�vхz�ep�s gu�c�LW:DQJGu���s����b�?�D�`��*���.�,�Fj���J^���#ݱsښ���]�56�TW���O�I$2NQDW'�߿=>�9��;{|<�ɾ{"��n�ێS-��y͞�����I�nY׺����7��V��*���hX��W�:'?8H��!�����瑍�UA�)��f2)��o���Ї��\p�M�Q4*�Q������/��%Qn50�.�	T/�K��︽�lxղ�� �F,ޥW�v���ՋM�@ғ(%]�^���&Z���Qwp��v��\{�e�%�L�������u\��l��oI���������G\�`���͝��\Z�en���7��|zL��F���8��\�]k�FSk�FwWm@�L(P�37����{������wm��}V�/�z��P���`�U���[�ڇq��m�1�+�����<j��|wN4�aҰʪ'w��kv[�"��wp����cc���u�SI[)z��lb�"���36X��h�Q�^����3�8�٫W�0�l."fXI1��,N��	2�׆���qIa��pQMHhWA7m��<D 삾RK��>�f�2M��tUy���s�� ��c�Uf8��^y�ǈ!�9����;34zg�pN��S%�c|$�K��i����o�t&Xǝu�]�)��4����Zr��{��������plн73���G�1˽2��a�ʵ��'vv��8�"�+�|��=fd�"���p3M�ö� �{�0����wE�=T��9�wx�a��uh"w����B�S(�9Q�5D	*��V��o9��>�����E&�i��Œ�L��]yoG�NSM�)��6	�]�b#@�����K�C�W�+ȟ��h�����<Y�縕3���ߘ��-䂟�(���p��7sK����V�}@$�^Kv���y��U���V���!��1�dl]w��b��{wWP��kgǫ��W��'ڶ��k��}%vxFݛ�Y�QI�	r�e9���[=8J���S\�Q�=�8L�j�z��ܙ#���(J�����դ�wwn�W�#��~�s-�D��[<�λ�=ǐ{���⣶���0n���F7�h4Ub�wږ������4NA���69�6���
;�'ӝ�}|����%M|)�:���b�R=[AP�׆�ڻ�.#��R�ݽˢ��mYѡx�o˕B�Tw�W_M��}��'u�v��p�����EI�q0��
�!˰���l�/vbW2�V,�7q-�ZV�f��{����{�j��=�*�v`����\����iPWI�;�>Ň,N��ä�un�KsNu��l�a	�֖�*[%�U[/܎�.��r��H<}�k��:�	���/ܥ��rV�y��M�I=u�I�d�nI,f�7#���]S�n��@�&�ҝ�J+j@Q�d�W���y�h�%���7��#__�B��Eev��nR};���f�d<�QȜ*C��'4F��@��X��l����w�ké�����٘7n<�y�2��-��Y8?.��6�rх]����c7�ea�P��¬���Zu澚��۝-ͤ�S���
�i�5wff�Y\�D^U�3j��VU�j�m[7�`����U&G�+3�7�L��h�*F�2�vڧ4eeI$P��́|H7�a��_M1���kr�cr�!�Ӌ��U����$Wλ����p���"�=�gɹc9ܵ�VGB�W���&wmM+�Mp�*]%����L�1ΙC�f�X��1�Y)&ͥtح��^h�&�@�UiI�&{�c�&@Y�{�v
��I
���l���rBqB�4:e��샹@�5�dĬ��)Ӧ8�����%�t�S�g��,27P�C�meCb��^����N'mR�r.&����.��@��>\l��m�FtG����?e��H��$�Չ��,�w1�.�N�#�s1�Y@��fù�bM��
͍�d���5�\�Iu�*�4&����]۬ߑyg4j=+c��v",��b���ĥ�J�:��cÈ[������9�w�z��lNj��vJu�{ӥ���X�B��	Σ,IQi�Z���u��-�V��`���8J��-'�`����$�-f�Uus��mܽ��A�Ր�L�F�PĨU���6�)n�G�-΍�KC�9k8h�E��8�[&)��0�V&�.�Hk>���k-uS��б�˛Dh+�Cf�TS�J�!�]�ԍ�-��3�0ۥ�����CS�Lպ�wX�O��E]w'1;�)�z��Q������*Pɼ�0N�;-n%�i�k-�``+�oqۗ�(��;JP�7])�\�AH�"T�gt��f�ֳ}r�tKKZ�kj�ƹ��)%�o6#�s�^�e��ƃ��̒�)�����c�8�`���k��aE�Ro2�4��ٽ�kCһk��\ �c=���ϯ�-����ڽ|;VL�h-W�-���^�vf���C�b��wk;�օ��\�QD�	B���PU�'���#�v��nߟ���v�\>c�!�Ҡ}��
,���c�D<���!$HBJ�[��v��;v����o��o��~�����J����$�R��>�)̊�]Dj�#{�UU�q���~|�۷n�|��~�����(���NUNg�ʠ�HBI!"��t��x��۷nݶ����3�$!!$!�"�UQ�£�~VE�Ӽ�,t��ݼ|�۷nݶ����o�Y�F�2��g|t��&�dԢMB�$������ݻv��Ϙ�zT�,���B2��s�#���qdy��*�UEP�#��)�E*?�|}����*'�O��2�*�_�z�H�L��L�J��$\�;�/K����ۼ�(�&q�99'�z0�9<���Y��RI��d�uU0���9�����a���
�֧Lm��¢u��:Τ#��v_X���st��2���Y}�;��;.�ߌ���Cw<������Dexh�����H2%��33O4&ܻ9��=����.���K�yN%���Լ\�L7j}�n�.���R8�&�����G�7�a�=�Љpv����1����W��T����I�E�^P�K��_d6U�7���l�����1����v��M���C\�"E�-�	)$q���^s�?g��se��d ��C����p������c+c�y5Cb
 7�E&C~���N���W~~Ѹ�h�3��c�zf��G���?�>���=����zcf==FU���6�ml��H<�C%���`�eW?.���M<`zp����]t�ge�5�8�-��NU�dwXw)J��dvS>�К��;��G�O�98�U���v:b^RO5{4��[#����.wҽ�}�S2׏�z���!�����:'�����.���Z��G�:Z���)�a��o�07�UB����0�:�`����ƹ�x��a���
��Ü�C\1�W!����j�����p�wg�=�9��37�=�.͈���;�F�,�����=���@��<�a��غΨ�C�b;�B#��E)[�̒���U��[͚�QԯF�w����ޟO��j�@�u��v��z�7��a��3|��W���J��C�M@I��L����e{��\]��=�}g�;�9������5��������n�]������[P���}l�v�̶nۼSe���V��R4䝞5��*i�␋���3�)j���D���Ou'���k���@�X_��]����f`�%���<���&�F��}���6��#C���FnL ��a�ʉ�i2tv�wfq��E!�b���4w)i�		�FC_Op�F�`�a� 4Q³q+|��ۻӋ��F�������N��O��/����Y.�ks�V=9����������T�~�!s,�Pر]��r��̒Ⱦϰ���I���1(]	w<�s#w���H��=�1��1Ҕ�c��1oik��1��T���iW>߾��}#���]��{T�����n��Fn��&��n�M��>�7n�S��34n��O$���hއ+md��z�pG�4A� ��|���!��Jd��_��}�v���L�TZ0�B8�%Hp���`�(�.K�9A�"-RA��l����B:QD�Q"(�#�/�����|^1��#L��bg�I���J�&��x�U���{��"gr&q�=�=��R�.֯��n��/������O]M�1R����n���z�̭��kw���Z6�4�ly��A�{t;裂t�����I۞�����H�-~��xTD�J�6�*ۼ�4>�1���s�,q�e\۞�S�PN;ʘJ��h��f$-�X���)�U��e<>�n��nE�6��v����+�u7�a��t`7�$G\�cF�a���t�m��m<*�))�<�~ӧ����+��d�{zn]��g⧗s�_Wo��R2�@��$�.�>�6��KT�����}��9��7p\ǡ�-��m��Y�wV;r�S�IK�FL�m�2�T�T��Yh��ƈN��\��	�؉�M��ҵ]�s��AsY�.���_G;z����zݽ3̋=+������,��8ɹAoioN�Mi�hT��t�U+o��j�ٓ��۽�V9ꒆof>u9��=�a ��w�,�t�Ѐ��!���r{�C���[�曓D�9�%eW�J��37����p�������Q�Y}�._j�f����0�)�P��U>��2��M����;rn'�<wBmعw~ӻ�A��8ɏP�y�Q��k!���n7�Y���z���왺7���O~���?*T��b��_�!@�Y^4�s���᭭�!�t�$��4T=%ީ��*���u�>3d�E>k7F��7��NT��3��9L�"�
��9Gݰ}U�-t$�l���MxK�x��n�&�i���÷��{!���7v��M�����H0Z\ߑ>�:"j}蘲����<;:���v�]H=vvc��VU���7�{�ttѥqW���кu'qDWAqotҡ�]��-g�y��g;���b��o��Ǵ5)���EM����	Ϡ�է�*n��}�T6�m�3)���3�r�>�p���!G�x]�λ�p����	�]#��#yK{j��j��\e�� �[�/��)&�P��3!�����	K���	�d�9=03��'�K������ۉ_w��$��/0�{ỉ���Ԅ
����q��;�癰���{�d�t���J�YJC�TQܼ�����f�W/W����d
�9lvu{|_�g9͚讘���F
h������{F�A��l2�{���}9�����>�L�w���C>)>bR6Lbg��yy���ޥ�|&��4C��h�3�mz�G?SVpDU-��H[��Pk�d�rjl�Va���?��8�ˮ�{Z2��sɅD����+vz�-�M��d>f�4��,��ǂ�2�l����5nD�I(��s3�/�`��X���{�g`{���sH����w��H���l(Z~�O�)U\o�����C���PB��C�b����0���5ϗ4R�,�So����Uz,��:^~q��k�Z�%l����؅�-2�؍�OdĨ%�6v�|�n��~Ŋ���u�+���Aw�`�D�}�$t�6Ӈ��>�Wػ)�+�7\8�6/טh��W��3�_ow��W�[���Z��%�a ��Pq��N�M7n��hx�������A�e!�_(w{�ƭМW{��5���c�<��6Z���c���Y(��i{S�to�T!&l���`� m�Ͼ��]~h�ܕj�^�x�f�Uz���V���n<^�H!����2/������>�U�2��﫺ݩ��<�3a���o�.��k�h)�E*�~P+C�r��Iq���z���WK��!���۳V�򉈐���Y�>���៪�[��.�6k�]��<zo �mbo7��}Ȩ	*���!�9�����)_O�?5���(��̟/X��q��}�xd�^��w݆���Y�<�Ku-���M���4/#{���q� �r
�	�Mc08k��J���ƶoI-��"�T����3��g�� `3��܈�j�M;c��b��w4��ɜ��ժ)�����-2�U���	�+;�QqU��;�޽
��r�=�֎�ٝɼո�<�w6��*�ۍ�V���Ǡ�s�{��Աѷ�r�G��519�c[ ^ q3����H��$Ji�hS���*�~SN���EDʪ`�����N|��/<|{���S�.�u�x��D�Uܱ0�;�
u�uM�d��{}�sm,/K���	�f�����h�>�b��OLb�f��g��4z���-�>����<1�	$���y]3�d��l���׎z�WV4f��Z�����-b�J`:�k��#z��f_�]�Px�;bu�]\ؾ�Z�B{����7�V �ޯ)*ϡV�j���w����e��I.���Yc{��7�g�_o=�k]O!u��a�F��UXt���L����*@J'�F�Lx��\�WM3�5A����s7h���:s\�:-�yV�<D��t�/i��Ak�Xv1O�9D�(���D����\%�����ɻg�����ëc�G ��%c���6��S�G`��K�-W+�H=V��b���?|m��h�C�hj�"��Gw������ݚsf^�X1�uڝ6�mF�=��[��y ZtW�X�F�>(��d����L�]��v��ݜ�Ζsm���z��NhcBE+��n�D��\�O�Q��3��G���� �Ν���j�ϳ�H1ٕ���[Y�.+�+�u��v�z���[l1<���݇p��D����|k�Nql�w۱��r��' ����v��G'֦:P0b�E2�t��f���`��D�g.��0 3<d�䘼[��>xt�	�7:��s���m�Ԫ!���.V�~q5$jj��������L�LR�-���u�h��2�dD4>�M�U�=��Q��(�2�z�u)��(��نa�6j��Ǜ�вmIu�&�a���zE�V�q��Y��6^�<�ə��ݠ��,/�F�03����-�gV���M��ʻm��"����YL�6�QW�"��j�SV����q���G������<a����:"����=5�uf��5��{'�_`q!�$<���KE�Y�'%I�s���f��"Ǐ�ݎk[�5�̇�����Y4��pM�����ډz{{�:�3���wޛ��6�'/S���٘�V�]+2�44�)1wۺO�� x�U����Q=��5�^�v{��v�G�����]^��i�L��m���7��������)l�5T5�����/��ɮ�^��C�*���K�z��&�L���)��ct�a��e\>�ͭ�9����{�b+��nF;�)u��ҿWR����5l�\,�=���/���b&� �"
T�d�Ce��W����N@��ݏ��Ou@꫟iW�#^k����np
�S�P�.;�Q,�3�Oi1���w���]�CbRIEM<l���hp"}>|�����y?_W0D�` ԧ+y�4]JWi��`5f���uA����57L�����$ic�uaQ�w�D��������j��Æ�v��}��g��х��߻�́����	�0h�iVq����-�M��)T'�)�[ًN+K\�9|�-��{;�=tr�"�w�CP�y��]`�hix���ro]GG�~���l[�g><����.i�o`�����[�:�{����-�,�ͱ/�����M�f��w����o�����u�F�uc+ُ2"a��S�u�ﴳ�羐�M�qb߷s�vL4��vW<���m��eP�quӟ���ދ����۠��&X(��vr}�~O�	��M�1wQ�ճ�çp[se���+{��w�
h� �ג��Ce��<պ�z=���]�I�;T|�ݖ=,�v/�a�{PH9���7O��w�<d2G�`���oGm���B��s�7
�t��+g��^�j����ݱxWcfQdcT=3WM�oG�ɊA��RF֮��ͯK��qX��F[e��NɌ��#��Y�έ�� F%s��ޫ��Tx��ǀ�Ҷ\����聱�<&�s/J���e�?��O%C����>�j'�k+��>	^��Og��[�z�����l	�F�ǵx���b�v~�#J*kV,T��ӆ�Ϲ�d^�J�O� ����5��!vJ�Ew87 ;v���z�Lr�+�uU������ݨ�T��ɢ��꫼��l��y؁fz�n²���9&��ov�W
�א�8����F�X��4����x�]$��ָ��O9�upn�M*^�RʽgB/��xB�����}���>�y��,��ʑTtdЊ���Mު����-7Btʭ���ٕچ#�.f���Y�ʬ��wW6Ɏ#Π�]�f��l ��µ�k�*2\(Ǳ�w�WY��v��y���h$�7��/��E�=�<.\�^[�.����NVaT#����uWu�o.Ϋ���v��R�Ƚ}��9?P�՜�+5d���܎�C��.=�n�{�:�� �n��CO�%�q�,=y�ȍ�ڌl��K�ԩ�ε*r�����}�%�zW]5�U����KT��ӭ罙����xg��FM��3�K�,9�+k�33�SçW �ӎ�]n�K�i�ԯ�l�+_�b��NP�@a�W1�G&�oHy�+��V�E�j�hv�&��<*��<�����W�(Ʌ:q*X�v�ŕl�!�L����-"V1QȈ�I�B��jvk�R�!"W|��B�0�w*���{/ P�^��AL�z�s��&��&�R:�_9ҧ�!?��?D�_�q�a�j��d)������;�3��C}wCV&V>�Krn��gw5E�ktrT(�����ڼ�¡�g�*���N$.��f��f�Ѽ:S}��U�m���.��m(d�E����Y�i��9BŔ��9�����4/�/����L-L�M�&���8�aͫ}tx6ʾ��0�cv.�CQt�����m��t�ηw+�N{<�C��eqݩxWΙl�ib�W�9sS6�[��aE��6�rZ*8���F�;�cYL��sI�Ё���Ѥ�$�9���<w��JO�.�4�qG2�r�G�0سp��}ʹ41ڤG}��5L�Xv�ǁ+aR��1�׻h��N�;�Ŏ�Jgd}IoJ���g9�!N�Y��5�6�9�����5k�evvPA�ed(�l��͏7�.���9���]����V��a;)H1/S�G�d�V.d�VO7��W.|���X��W���C/��ڍʈ�=��V澺��-�+]ܰ�3wE,ٔ.��������Y�J�����t���݀��g1u������ݝik۳��Gh�-�j�s�T���{���VUsK(���fv��P�"8�(�D��N����
$dd�R�$����t�����۷n�q��>c�N�yD�zS$	 ��7�h!4ɔ*��\�r"�WBo(7lq��m��nݻm���~��2�<Bvﶗ��(�
���C�����ѿ�.��<|�N�6�۷nݶ����g�I	'yq���Q�$�+R@�(�)�D%Q�Y�N1���|�۷n�?>>c�����MziM�C�*�AeQs�U��f���_��3��o{��nݻ|��|���zv'��T�Z���8$纄��2�A!P�RjJ�EB�z�N�|��۷n�>��~߳��O�!V�h'o�/����PG1i7�ۑB�Jꆉ;��V����pԊ�j	!�Q*����W�z	Pi˜�8�$'�u�u��-�QeKκW,���+2�6cwnwv�g�����r�*�©$����"������WιX*��X�<�.�'��>�wyED�8&q�X|a0�p���	D��D�Q�@@�O�ܧ	�Q$6���$'"�	AH���#�IBH��Ɠ!#�-��Y$8�"9A�R��w��N�ܽ�����Io.w&{�4����7��ن�d�Pi[Fx�g�8yV*����u��\�l�H0�
H�"f\MN3,�(.D�("�<L��Ӓ���*�D$Ȧ�j�)�*A
0"�� �0ALӑ$È��r3"DD�H�JKe\M-Di#�����"�@�1N�A!H�n8���.6�Fq'eȜ|L�	"8RnR���0��aA	%	BD-F$�U
�͓?�!�se�Y5a��� �4)A!
~NgМ�8l�R�Ą��Б"���<%��I�(0L���䁢䈸�)�̐�$'������������_E=�����%��9��5|�n��h��]���x�y�E���L���K�Z��s�hT[�BNl�����w|{��J�P�g���xxz�����3��G���Q�j��v�湫ޥ��j���E,����H�x��a7!��ܓ�ꅡ�Fg+��O�����p!'�-�����d�|�F;3�΀�}�k֔_`͸N��^k��ؖ��H��� o l��f�I%�B�>(/�'~��~��6z�H5y�ص:�v���g�n�E���ϛh�6fy��^�z\<����<b�^��L.�(��u{�U���u���i�Dbg������{Q7uE����\��5�ݝ�y��!��u>J���GL;��.�p�˳_��_�����99Y��T��&�����e	j�,Mq����=6*� 
��^��MR���/��9��,��q2�t�"������d�FDГ���6}����� ?��)��'��L���zzF�f��h��l����\����Y�Y�%x�3��F��:�̀ך�MW{�7^��(E@򽬾���WV�����i��'b����Vgt?F���;��oh*N�
�b'M�J�?����7�C[�=r���r�-\�e���OQ�OS{���~��`�ot횺;V�um��XO.Z�YZ�%ǅ���&�����f�Pu�q������q��W�Yֹ5�E�u����|�.�pIe�d�K0w����u%*U�+:(�v{�a����ڴX�~z0�4��C�%^��O�|�} ���q�H��dgoMYA�SޜTs� �5�z��i��;�)�ۻ&��ny��g��F�Ю��sٱ�9�f��ZT����]�@���o�\�v`gl
���%���(�j�3��}n��`�r��j�R���U���o����kJ��Z�1�A�/N|��]�������|[���s�h�J�3$s���U��b�q��<	�N�����q�t_C�j�A�s���h����wQ2�F�X��w�i����Ɂ�����'�47Cې�6D�8��>�8��
�)��V'N��ƃ��N����&��%i�Pi��E.{=�3�X�,����r��v���E������=m1�u��v��j�]�F�^�i�xB�x���y{�����D|��x�$�ɍ���!$7��y�;�,}�_�ߎ��C[����w1P|����a�v����77�]|��fQ��@�P�G�Ҝ�s��l��f���|����'�w%�Ou�R�n��C]��vC�C�\���x-�F^^=�p��fjvY�~�ݝ���U�������ϟ_z��n�s�� �y�H$I �AA$�}��;{�sx��B��������̢͎E�3���s.�e��C\Mj>�,�fS�E׊����Y�8�#ޞ�A�ά����d�d�8�άK�Y�J*Ht�zfo��{&�U/��V~��>]���pO��OFWs�ԥ�o$W��OP�-������:(F��>R��k�j�V�*�i���c;��V�ۻ���� ��W����u��ukӵne�^�j�5�<_�e�,�&^:� �r"�9̞W�u�>dy�SW�W&�MS�GA]<��Uaԅ{�^�Q:����@�&�UT�\�w�gZY�BrF�|�l�_����u3WTU��
d>�(��z�u��="�Ɩf`۠P��w�b��ܰ=�u�����q��\��+��zb����g�����3+��1�E�[��߽�3���A�}�!�����ީ>�9gK'�{�֤���4�jh�u�#��M<����f�vy���z����n�,#\�%4,�����>�r$��w��u��{몣@�&�i���θ~��WA�Ml�̬>�ތҬ|��|3�d&ϛ��̼�>�L;{�D��%�*��Z���N��j@��AC�f��{�_�*����ݩi������}���@3�6��[�&�R�Ͷ7�[�.�X���  x	�JuIL�ϲ����� c��%�s�ݫ]�`n�}z�m���+��	6��nw���j���G� z��D*G�����*�l��M��^��`@���4����*$�\*_B�T&}n��x9|�Z,5/�w��ƺL�c�nT�P�K;��qt΋�V/�����ܣ�����7U���o�+&2���@��9�8hʂ8���*b;�V�+1�N7���Z"�Uާ�M�����<�t���\�����>m+���S 1��.do`����[��^^Lo7nC�+l��Vu�ܧp),ހM��;�w����<���ei*��O`%SBD���x�d�s�C40��솳y��A1��m��.����ۀ9�J&��3Ćx�%u�fi��=V�5=ִ�F��S)5Oy�o�M���tθfs��
{ޟPRN+���X����*,�;�ը�)��dk����E�D�̮�]��*���%@|��=u�ʞ���<�ShCe�n�/=r�.�f�H�.#1m`K���M�M��2���	"_�4V����~sҼPv�U�Fg����͊2�h�R�
ki���$zn'��5���vM�a�KBu3l���h�ڗ�}�t3䬩ܕ���z�D��G�cu��G�v���U�}&nN��_��� 3g���Y��Y��ZH��	�m�G�>nguZ��~�U6���y�B���!I{�5��黣Hpx��C%�b��Fuי�_dR/{����=E{�����S��G�A}K`���x�N�s�R&=�U;����ԗD��U������;��]"1g�I�%IW]O�о���|��y@,\��@�I��}�96�ګ#B}[�n��ܢrgr��y�������x���z�*�홨� n#w3��w�z�޲�V{e�C26�ϊ�C���aU,�z D�x �z�{4�������9�-n0���k'X�R�3�;�r��fux�������3�f����C،��n��h��uN����c�7��k�n=�[��A���ÛO�cs_�uB5FZe>��ѱPa�L�m����i1<�^�)��=����c=��Ǚ>�C��h���痯^H�f�C�Ůl+)�λi#��-�A�=��p�m�]�ݱ�9���ug��=� {O���/��K'"Syـ1=�N1��1�
� �裧g��s;+O1�ENMn�=}���3�`|��q�߻L���]��]YyHe�xHa71���1,Y�'=2�d��A{\��@�U���k��3��#��H�1�N���5�j��
�G�����>�UQ�/P�V���q��4�\ �����)���W����/���f2�s&���m�X��UU?]��b�;�]���(��_U�L3�e�ǍT�.^�8����➥�{8E���x]��"�O�]m�z�7>�`�� �T�P�0�̐O3�K\�t�g�3H6�H�����M"�J�}�l�y���hF�%�4�h�F�Y]DF��Ԉ�O5F�d�Fƪ���{�d5e>�ؔ��x[%��k��a�ٹu�"8]�^�oo��.�=�N/�ڙf�3s�$fU��T�0p�\�t��]Gr.su7�v���ҸT�p7�Z�uMÑx=�棁��u&�'Yb��5�w���l:��n���Y����E�f�C����
��gwb`�  8��������y�U�0���k��m�e�_��;�{��9�ȸn������D�N��y��c��%�깞]U~=W3�����]�"�B�ZD�XNM)
M�c�m%����'Wn^F�s��į�7����z���=��R��2�<�����W���V�(��ޟf�"��smo�����d�&����ڐ��=�@`������9��E3'����!���K{{j/Y�3��y^�����̆�M-��OQ:��Ԣ&�H�oW{�G�	�\zA̮����B�}�w�0b,2��w�
(�Mҟb�䨍k���|���S�Q[�uH>�q�\4;�����u:���5.��}�v0�F8l<�/oS�X����라-������ d���֦����m��5ox������̏ʺ��A'ۗL*��<����'+�Y��~��S% �`67W��\�k�Z�q[��V>��}aM�5z"�N,S�w}*�>�[Չ݈�`�i-�4��N&�q��x55��+$G��}����{�!���!6A�XQC	��\�3���7�Y�TL�> Ke����Ғ%".�fbRB�0�L�$L�� �;�n��MCq�*��=�j^�w���s���!�̈K�Ř�}P����^q2�9�l`8�vZ<o�-�Ѿ2��;"����*��6�77mtZ:
^����g�>�X�u�E�"�-���6�^�z��an�?�aGLM ���3�hH�K�5>xR��װ���;�N�S-�5k�*������\���WvIzUˢM;��C�W+۽RU؈�t9 5V�_������^s�cVHϨ4��5�kj�p��ti%w���V�d3�f�=����X�7~���<֣�!�quW�Z�/k��q���/x��)���6���"�Eb�\�sO��U�l�Fu3\��{��~�}6����j�BT����|��p���h���������,� u�{yt��}�&�3�ə�xݴiI<�3x��3��ɰW8J�2���<*�%�����j�Z��XO�3����=L�w&Vu��[���仧pnh4��t�iڶ���k�ȅS�`��oZ띃y�zk�����n�R���Lo�J�{ȏu���F�z<�˟�d5�N��Oqw�^r}�fA���OV�!3�H�2�����'\M0�TҺ��tzT��k�&���ٴu�2���*��/��0]^Q��|��z�׈fs��Z�˳fT���㓥����ّ��gdNI���L��Y�K����l�ls�[����1�oO���@�Prz�]ÆVp(���[~5͵|�Z`ML�XԒ~x��F�]�ږp���׾�z�"�/���t�/ߊ/�eҡvlD���9z�R7�M4L"`Ӽ�M:��ʉ��G�{����:�\USzj�	8vf�0�;���3*�nK���C�m7������{��F�.;���eˡ���f��]��WvAX�\�MI6{p5�1��~����es����\����ϗW�����=a:�r���)�lB3o��u�fq撮m����Le���1$�&븸+��'�p�=�;	��Ej�pʽ��N�Wg��Q�����.J�[JQ��j�݁f�X4�$d�du-�����5�r�d�zY�H�mu�Zn΅n�S�}-^�=�g�ʐlK����ݍ�NeA�6�������ݬA����y�LlS ����5j�]_J����Y��ީ�f�C���3u��jc�<���CWEI�*ƧAXCK��u74�#�\H$�S��U]��]�����zZ��L�k�{!0������ՙ8��F�.ۜ�t*iPn���Ik*�}B�r;W]�r�U���,����R�D.$�2�'y��/p��uб�y�i+c!w�fEj�N�<�=���[u-X�T�wzë\�	�E�1Ǝ>�Թ��ԮjTr����}zY��ԝP����YF�������SP)��.�sv��:m�e^d�`�,�L���J�z��6Q�n��ӣqv�kު�JӮ��	U��Z#39n�$�7��Z!a�DTDN��w�a���zq�rۤՕ������'IҀ��H4�Oj�EbΞ>D����B�*��A҇����[k�s-�Nڈ�l���N�'b�IB��t���(�12�a-e6�I�'7i�)xN&�/���Uд�eiE��В�JMN�&KŗL�	�)\5F�j�b�d�X�X��JGT鼶�av�n�Yw�������#�4Z�쑵;n���V�@`F���ܥ�
0�	�l��Z�3�/n*I�t��.�����5U����Q_֯C�7.�m�S1�o�4�Wk�8��ܫ�Z�2i�:i ��^3Sz�u��8yleP��6(��3������O<^��j��L��Rv��s5C{yg�S��z�yL�]JgSY�}'WHP���w�Cy|F+/osPw���8�ԴE#b��O���V��1��g�f\A�Y�Zr��os����XFɭ��.�"7���9���7R��q��������r�DUco�LF�\�+�KE�s���ڨp���lL�]�]L֎�9�Hգ �̃�ܛ�����S�ֲ�t��� �WuZw�U�P:x�[P�V��n.�*ݔR����x_: �J�,��
߂�\H�ݗ5o�I$�]��(]6��wN����;��ɹ�.�7����#O�I�����T�q�ֆ���Y�e�#�ޱ}D�	�{v��;&.�"cc�a����ܽ��h��\���)�B�������\��y��;�X�U¬D���&Ff2N�BR��Q����i�;~m�۷���~���g~7ߟ_��3��e�Y���»QHд���LI��e����|�ͷ��;v�۷�Ϛc���!�U룄��'��.�d�%��ɕ�3�G(�rp�~�7�ӷ��;v�۷�4����d	5(�j����$��}:y2��4�]�ҭW�������nݻ|���>�J��D���ar��zU�,��HETo�0��r�Ԣ�=hv����ݻv�����z��T�I�ߩ;�B��֕P��T�?�	��K*�a���P�*�Q$�\x;x���nݻv�{�u�������Z_�[�M!�#���̌�k�֒t�Ap
��p19d���gEj!r�������t���I��ܓ+����y�ܜR��eI%Uf�N��4u=��W5����L$�UȭJL�
É�_�L��.!HH��R�,�5U����۲�9�afCn��V6��Ok:m>���u98(Kl�'�ݹ�M����4����9�VJC��z��	�^n͈��3��%{�l/t��]��Vݲ�F�5[+�W�����#&�-QBd/����������u�ʚ��D�^[?'��;W���"�~�=�E{-	���+̀C��(�����`k��/s�⺸:���UOkk��q**�>���;�Ƿ#�hj�wW��OR,e����U�ߧ�kYta���d�׀_@.�����WwR)x��jn�6�j���]�z/k'q�Ջ�S��S�\��y���I�{{����q��Ѷ7��U{X��A�0NM,����:�J�T�`Sר�ݻKql��{��h�V�R�{:�����+f��`���ި��N� 7A��˗l���.���ݓ`�����P�`z���/�*�ک�_�񐊘?�3%��S_�:lr�]]K($�N4.�>+/5Єe�f�O�� ��ӊ����s��D�nv)�����}��ɳ@���KV{oHݻ���佼tE��h89wb��2�(����y�y���iS�g������,G�&��w����]���&��Td���ooa)��,ȼ���`6 g�F�LM���l�q���Y�ڎV��x���;�5{a*�����	SG�5��<�`=�B�"�Y5uT�9��/%og<�)���<H2�����e�M�Ӝ�]�G ���%Vlz^`w84s��m�����5	F���/�N��[��u�l�/[�2�����=6����1@->��w}Vu"����2�۷]3�.C� ��q;Ҏcꎎo^�l��a�*�*J�ܮ���l֦w����rq;�9/s#O� vǼXJ���~����#R&�Y>^��`{�����݋�ݗx��#���kF��}Y���1*� �O�\��
�����ؖ܎�+iG�w]���ثyWpH+Q��v�����l��m>��1���X�J�ph{��;�X�7�O]�0mξ�,i���C^�5�sE�k����L@��E��r)7I�vG����PZ��=��
 z�^�Ů�	&!q�Aȶ���w3Q�!�cM���IBF��R(K*F0�
%�D����!�f��/)S�F��7T�ԗO�g_����5�`����L�ޖI��V�]����gu�mfp留T��UXΏT�tR���#ǁ��.���lǪz�<��u�o��)��њ �ƣx(��#��>��1��d@�M�f/�������$8���$2e��|7L6Ȁa���L�՗62~�'��� śx�u9�.cXgw��9M���3�^N�K��@k&cTWJh��K����ҝ�N}�P�+�#ޏn�@���U���F}z0��{��zW�y�)��iDi�B:ezX��x3���V�3�[;�F������H*�g�vwo3��2��[��6Oy�/�`RR�m �v�P��������Mo�'��dd5�5������i
ו�N�f�!+,U�{��o�^ l;�\橖=���v�}����Ǜ�r�`�K`W[���sM�I��)�<�(��o���Y׺�aN�VO�O��7չ�ۏ��ھ.k��(��k�=z�*uN���aCr�Dn7�������.�� ��=���1�&��U]�M~�c����W!뢴<S�dz4��v9J	b� �w�ܣ/��]��۠��.������"���F& y˽��殞�{ò3�ɞΥ�ʵAcL1�!��l��UV��3dm��´e_Q�;��=.s��b�k�Z����?�tѼ�/XPn�3�x���=�@�͑G��9�u���qO�3Vo��G����X�w>N���+njK�:�S)�����3�zjh)38=�}1����A$�C;�1�1� ܪcyH��Ψ׼{=�t�r)��u'z��-��/TA� �2�d�`�a#�|�í;A��צ�74��V�rkZx'0�rcͰ������v�螌��ת8_L>�/G_[��wfvn�_W�U������=�N�OM2�9"M���]��o�ep�N�`1�w��(uޞ���o�n���Y�>T)��v�7�$.��Q�x�1�#�{G:f��Ի��ۇb��I9{M���8�׌%�7�r����x0�U>EbmV�y���ϟ|�����J�{Ff4�I�O2�v9��U)�G��Ү�j�,�,sZWU"� O,^����w;�w����®�������A�e�½~ZJ	<�[v�`�L�����a`{�V�_opK �ǣ���@�aΟ��p��Oof�gKO�@��ݫ<�N;-h�d:�(�E�)��}+x�e�s��~WveU���n����������0e��P������WC�^�K���6q9�f��ew=A�5��l����b�N��و����)�oY�|جg�5`��PIK<s�W���#oт�,��k�n��v{Ƀ�7{����F�	t<����_�^�H?���jEp&^��W>s�>�D���j�5���Dhp�줂�y.�=d�T^�SUUm���W���f+�_u�ސ�ge!��|q��#�l^o��P�����t���f����o��ك���عv�����Y���x����p]���}�"� �Ӝ����۪���z;V~�4,A��w#M�!�3�D}Z����G&Ig�����j^�#]��]�Z�x�B��e����H�Z]u��}EG�ز�ϟ�Ƕ�=�����p"/)ׯ�e}t��A�Å&�޼�ɳ�N:� ��Ym�b��*`�05�m�%��N�@�!K��nł���0S�}>�hQ�4��w����$L3��=9�k��6���R0{�V�u��5#@Y��;ѱ��V����o4��v�H`���659��M�Z2��C�����l����Z�q�%�<M6���ۜ��������톆ꈾ�̮N/Bot^7��i�q�;\^�R������������K����U��t<��Q�N:nY�Q��uVϒ�>��]��i\T��C���,��F��<�1޵+�=*:v6<gֲ��h���v���cz����SZT�aқH���߱��.Nf�%�eܷ���ɹ2��R���p�C
 Q���|4��g�w�Y�fN����'/m��Mk���0�lM���ܗ|��r#���j	��{{�u��Ew7��� r�� ��Ia���Q��/�{��k��
@N(d|eӌ�J2�1܄��8�TZM�����n
��*3��B��9ff9y�U�T=�Y���.oc�yf\����]VЄF�h~�ӻ��*N�t���X�SH��Yg��w/{�r�C�����|TY0.ͥc�� t�h;���^}�:|s�9�V�6C`�N�Z���U'6p�h���k�{L����]jp-Ofv�7��>z쑒btfi|!�o��u�-��5��fz���j˳�yU��q,w���>[��335yrx�>�t�������ev�M��U���§�=��T{vDϫy�%��8��Yg��캤[������ o�w��t��L0�T���;���Z���7�/��Y�K��j�5dY�B��[B��'������U��������k@=^]z'�7�y>W_.�H�v�w��P�[�sn�F�H^�+�ݩ��[<:�
���[.ߛ�႘��+�>���A���9@������i>�n�ՇW0�הc�N!���!}o�(X�:����oen>|��X�XI̒:5�MDg��=,=�F,��,��^��:z�Wt	��$hE�.�Y���7,+�Z}����4���\L#~VCGUק����Oj�]2c)��I��`��O΋Nz�����#
Z�pC���NQ���*]�2r��4-��UK��T���oq���k��T��lی-�缣���������z�o�c�M���β���"�,A�༫`ej��>ԯ�Ϯ}�{O��*k'�L�}~w�^�ZX	K� _��a��<�K���������w*�3�cWj�m�f���E�)�l�	̊�4G4n�gp���,��2]y�R�A�+�7QjY�=!��p~͑Ѱ+�{6Or3��Uz���_[�+R�)������t�ff�y��]L��6�y�������5��_�QA�30קY��9}�ˊ�t*�5�ʸ�i���
�|��q�ox�J5�G��^f�!zj�����矫�s��=m'�2�M���q��c��4���2a�]St8������ҩst~ {�Cv�ʱ�Z�szI�D�{7#ͮ�}ʤ�>���8��V�)wwr�ܨ���,dρ�`�f���d�[�p�ÿf6i���ﳴm�3���53Vfnڑ<��%ם.f�B��D�}�_������Ȏ�>�j<)Z����a���,��4�l�Y�3S߼N��gͦ�]�x��(�;q�3A�h0 e�?l�V]�G<Wzxw[�^S�c�"�Lo�.�+�ٚ�{�G<� �b=��]��cw_�+gBU6L�z�2ꗹ��Z��E�.�N�ffo�����P��ui�s���`�)�r��Sl5T<����0x�������z��cԫ�X(�=�uN;��n��1�i�s7VV�-̧�v���EVU���=��WqQ�>�y�t�|ȶ�^Ny*4�n(�ێU��	*?�v��%/�Q��4�Ar���Ks���/��]��{�i��4�ruGHD"F� �G� �UD�ۈ�|�i�c�����T��j�t��])�z�q���* {C��޸��0��ogv<�9���x�K�a�|w°�ex�{�l��\
2��C���Ok�^�tю��1�ڋ���*�2����O��l��o��wYV�?^c��WpӻA���[[����H�II�E��^o���g��A��/)�w��m�>��U9���ՏK�"Ⱦ��uF(Cq�6�)����$5�	NWy��J��4o�*m�{l�,	�w_��~�Ѱ3��Э��fr$�a���P�oj~��L�қVy�_P����mKw�R�8oe���2���]�,��^jQ�J��|36��@�͋�.��\c�c`i�I�u+y�F,�P��2�;*�>��z�9^d�ݮ���a����д�\R����}�~�b/:l[�1���aM���A.�<�_'̆#ce��]�����\�*��s�?��G��ڿ�G�Uk��@QS��_���
���� ��� �X�`´9P��p"�@`� �B
����B(�� ���d`T(�+ �����,�, �@B����"��*#La
 �$"
$"�$ *&���m�P�B �B*@B
�B"*@B*�@B(��B �n�B�A ! !  !D ! !P ! !P !P !� 4E BATQ �@��P@��A��D`!DT�� !�@!���@`!HDT�� !�J"��B�@FA��@`!DR
�@R@TִU !HDT�� !H+ �T��`!J��T��`!E��`!HDFA����9�
.g�*�(H�"F($��
��w������|���C���?�������� ����� ���?O���~���������C�?����@ ����TU��w������O�E���~��C�b�����?����I���b|�������?�@�2�+�4���RARDT�T�UI��� YYF@E�E�E�E�dTd@YX��AaX��Ac XDVE�XE�XQ�X�U`��Tb@E�T`DF!`�X�@1X�E�E�cdE�A`�FU�d�D+d�DX@X��DXE�E� �F+X����F	dQb1E�EdE�@Yb� !`�E�@X`DX)ad��XAX�@XDV+dA��1V @X$E�011V@XbDXQ��1��VQ�0V0E���Q�`DX�E�0 �@X�c X�XDX@X�X�X�c �F "�E�Q��E�$ ! ccab	�X�00 �@*�XFE�F EX@Yd���@X�Y(@X@XDYdAb�D�D�A�ADdT@ARAD�Ԃ�*�PT$h��
%��������(� "(H �2
�����p
����/������A�p�}�k��*�?�������Չ����O���a���M���
�
���'����O�� ��A_���?��@A��~���*�
������A>�PP�+�\O���|�4�ب �?d?��?��EA_�$�_��0�7�?�o����������`|4�*�����TU���p?����?�����	A�u����}�ބO��A^%�H����J@���?��4�|�<�� ���l
�̀ �?��������R��b��L���� Qq� � ���fO� Ă���JHB��  (�P�)B�P(P�  
 (�AT ITR���P 
�P
��سl��Ll�Ѵc`��FjƵ5�F�e�X-mm�$�U��V�&�jZ���)���hSLZD���R��MM,�VL��(�A�b�kZ�6����%S͖�V���[-���Ye�I��Y���3kf���,�TU[e������3mi�Z��Z�af�md՚Z4m�[m"٫j�-Kmj�iRԗ� qvz��TjMKj՚�fղJ��n\e5������Z�n�:�k%�Jλl䴬����]�SVTZi�4Қ�R��jJ��֪�[k%��h�����Y��  sa�P�B�
U	�%â��(P�B�U�C�t�IU�5K��JZ�B�ҍ�b�l�45*�v΀�[
N�i�Ume��XKe�l�e�R�ml�%�Q�VI�RKKj����  ��h����ܱM��M��V����EjZu˥Sm�G\v����N���+ew�V&�U�,je)��ͱ��M�[%)�[h��b�6�K^   �T���U���T�U�9�R���U�I��N��CX˳\�Z�aճ�kmkjf骊�rt��d�lu\Ჭ���5mmY���f�cf��m�   ww�0�Ue-C@�H�6V���2�J�̱#DRֶ��u��&�Kkw.���u��Dڭ�)�VʶsST��l6հkL�ͳZ��  x�6�&�b��j����U�;�  ؖC�h� ��k�p  5�����&0 k@@��  j��2նfUU�Yi5Z�K^   ۼ ����(P �8 ۊ� �ۅ� k��:P Wn ��I� ����:u� 3v�65�ڊ�%��m2֌�� ��
 jX  �4��t�h ;��  �m��
�7  �+ v�`  6]p( j�[+m"��[j�-E���  ǀ  {/n  �ڶ� )�@6�`
 l  �6�g  t��@CX (P�]\  �\m%�m�H������f�k^  e� M�p�V  n7:  ��  #&�  ���@،  �V�  �n 
��@4�) @��a%%* d ��D�)4��20�~jR��  "���F���  �J�2���C5!8H�P���P����Y !9���M���C%?t1����P2�=��>�Ͼ�>ͷ�ϛ��`��m�lcm�i����lcm m�m���1�p�����1�����������	����np��nW���(M�p�ԥ�I�̽8yܥÌ/�۝�:�;R��+�oie\O\-(SUm�tE���s=a��'�.���v��<��׈����F��{�"+ǑӶ�������U/i����ɨ��Za�ֺ��,�Ɍ)�r]���W%��t������+oG}����wJ�;�[�p�[�r�]ub�Di�Z,�X�o�
X�h��w�LmpœA�׉o��r�]ӹ�Dz��H������ɰ$����Y4؎��H5�M*���S7�-�P���4��u�M���.ɰ8,b	�z �{s�]�:(k�:�-�SS��B�� �L6�5߅�J�^��pN�d@P��#u�"j�4I;�N����ɮ�h�����=[e�jf7·�.i�K��+hX�A{���.8�@��A�H2�1�7H�>��(\�'�äT�q��
ېf��ε���lɜ�!�C@Z�T�
ŷkZ��*R�҈N�2�`�VjŘ�dD:	Ƀ$�W}n��f��9
�K��f��>;���ќ7S���{Wk`��� tzst';uwË-�|���/l�vp����D��t�����(�,���n(X�����븷��BW�c��`t��J����ƯwV�Os�'s���C�;B\�P��/k➽�8QHot�Ӝ
�Q�</:DUw8&���I�v��*���
����5�	���h�X�'̀��v��p\��5A�8ްi���Оp�Ĕ�t�R\���1+�o��Ci��w�7X�䦂��.��-I'MҖɊ����.���Y�+����up��S�4�a�y���?�77
�tor�����!�8���W�ϓ��á�]'���,�f^�o����9�^���a(�@|)H��.�'/
�����b����ހ1
���\��!F$���-7�'���4��!kM5en��o\�yu�����LyDm���d�F�j����T�G$�Og7-g}(t�^�c@��7���kJ�k�^h�a�B_�gT&�O:��L�&1�n�_8�I7{,l��PLk_H�{j�b��z��x*a�Zw{/���Z9����mWw��	�;u�q&Ľ�i�h��cK��3�n�`Ct��ǝD�z�e�rE�@�ˍ�9N���g��/t�7�4��c�*ě�l��-@d¶�Y7��x&�#�v�ZZ0v)��rf�EB��y2dK�1�p\E�η�%Y�'��R�b�p2���[�Ⱥ+c�e`�~�^���)�5�L:&r)nj��:��o�Z^m�vsz>�m��u�)Ai��:�eޮv��-�j��i�����ܖc���-g2"��ބ�a�)nnv�h.�]v�q�ɼ*=V�ٯc�y�0j��V6]�vnRv�8�S,7�l���ߢ8@' �\���̷4زsr��D{��}�wq���]���d.wbap��X��w�t!�eQ+ �1���q@�-;�+�!q��\T��'7�N[�훻[��t�}o|녁������D��7��n#w^P���X��I,���J0�^2�f�f��\��J�*� �cq��I��NA$�<�v�d���;��I�����d��ڃnK0s9��,��(!ػy1��ؤ+	\���9���UX�a�籣۸�n���Y��5�ut�$�QKc[�+��%��w����P[�~I�\�MtXsTz%�{��т�.��;���R�dԓ�1�4�u#ulx8m�bs�6��i�NBі���	ƪa*�k8iE��ot��������;�r&L�YAol�iУ]RxFE�rf��L�pӷ#��	`V�Z����p2W\4n�c�>{���u�P�!f�8u�.A�F��)K���jGV����^�v~$:D��WF�	cB�܆	p-CF*�bX���G'ΌUȓ�&n�;n��ِ>�Z�cd��Wd��Wu���/$�&x�1j��=�f1�S��EMnb1���P��Jn[�$7a�c@�U�7Q�e���>�)�سs����Qٱ�5�Sr��-��yv���l�0�[�"�$�n�6�!&��\�T�ê��+ˆ�+�"��nq�N�`YM�s���މ�#,7P#�3��AW�w��!��;�G�L�X_!��76�C�܋K�6�C����� EmӈKE���U���oǍ�h�\˖-]�2!�����էVp�(���˓�Ň4���"���>��Uŷ&F1㹰aA��1t�D�с�ǇZ�������1	/]�7e1�G�pzcɞ-:���\����T#��Т������&E����M0�.�����)�F'�r�3�Ѥ�Vi�sh�q0�vX�LOqꃸ�a��_��@(�7�8�NK���S�Ƿ� X���
xl�j!0�3�P���45٣��9kVX�{݋B���h�n��v���v�J3�}}n��f��ͼ�{p�x�չyi��W.ca������V e#t�-7�5f�zW1�on�O�P���qbkʱ������Qm�s��P���c/u�n��]ZS��Y̦��(�o�TLM�C�>]����;�� ����㺟��~9P��.�^����듛	{T�y���޷5Y��-ǥ+��r�*�tC��TN�E��!��𹲱�B��V�5��b���3��F����@�Ԍ����\si��R���L4����v �wwA�H͆��p)�K���F�8b@@� ��Ϯݽ��A ���&�˦P��nӇ��[}B�,�\���5��ۯX��g&q�w
����$�iJ�;�h�¾����0�U9�h�o�[�޹���6����8f�D8������w/h[pj�{;`ˡg]�� 3�T�#�X���;7 x��9��2��J�f��>�P���&��u�l��]��Z�0"��h{E6s�VqD:;,�/D~W�30M#h�u�vn�w'�}�K/��6w8�Ϡʌxt��7�^�g�h�o.t������d����%L�ۆ�5$p��rw)}n��i{���<}�^rO�÷���A��4�37L9`��A���四I�]�vcl���وG�T������&�zE�,��P�i3&���	�µu�D��V�7�"nA!����YrE��[=:��`C�'���72F�����C��6f�ɶ���p:�X����$5|�^�2A�5wc�g�=�H�I%kgj�6��j���fk���p�.��;$J���#��3�젗�c�0��V���ڄ��۵f�1��n')J�'<NZ����;[اj�P�n-��5�q�˨�\t�����
�B��.�6��z/�U:3��Dֶ橂9�]L̐J�f	d)��w�L����V��Ӣ%#�&��78>shln���فD�ǣ��4G�{jb��j ��@�c��r��6�" ��se쮃��b<,�h�Ѝ@�Wt�2��X㕵p�7e�L��������L�I�O�-kV �P'C؆>%^I���hOhE{;D�:�B��7�1�5��M���;�m�����Ma U��VVw
c_Z^���,��=6�^�-�������Zm�.�H�� R	��C��w7Uy�9!��М�(��#Z��U)v��{'C���p��Q\�q��2�_#�ʽ�LY�(p�ؕ��F*c<���66�׍�{&��x(�u�0G��M��)粌x5��8�M��b�u�]�� ߑ=�1��.�{�r׺F=�湚۩��.嗞Z�B�Kq����2V0��>�X28LR=;��#sH��'B�ù�Y&�-����4kj�ut�-�!�j����y8l�!����.ԕǲc5�(��V.b�<���pLTs���%��z�v�5�oiZ,�׶b��%�0���V��F'��r������j���@�.���TѰ�nԡL�p���6���!�I�,�t[3���J��
Ӱm�:�5njT�N��w���mJPn=G{v��ǳ�a㳚3i��.��v�;K�!�gc�J���G���u�u� �{�������DL�X7�+F�E�sk�V��Y�ܚ��pO�i�a\: $k�RN�X+�>���ш�>t�xnr�p�}�2�s�
\*�(AI�Ȋ�Ũ��Z�> 
w9���jW�p�lKWC���@�$l^U�7��m#�Sp�������n��f�u�}-v���O���Mc�:%K�@]J&�F �p���~E�9r;�8�;��//Y����`Wkݪ��ؤ���T�:?�i�Y��d�#�<�w���I� 9��d��o�v,�%�t��t=�t�Y�������1�����F�M��m	�2��Z�k�Q�i�\.��V#:�7���y��c�3{0�N��Ù^Q��#
�x9�;���A�lK�\u� �+]�g�Y��Иv勦��.%Ӌ7sE���@�0�O}��=��!���B8��\ ���e#H�V���1cbOD��aE��%�QlX1>�Z2��������3A�22���@���K6T�KI���r�&bb�l��Y��e�N�� �D�gnL�;V�2���8��@עa*�	�J�ۗw �P�h/�0���:��.,����������9>Q�p:wwY����tt>�ay2�/r
�#>�z��ƧTC
ۂ�\;:�w<�P����kR�*�gP�R��qUZ։�ݸ�UV��"&f�-)��g*9�^�N�/&���<������a�ť�7�c՚,��^,��9̩M��H�����t�W���u�y1�1���ϫ��0d�2�	Ǳ���B�n��̀%�t���L)�V���A5�tU�R���Z/$��ا��)��c�xR��N���n���^�[ͬu��`=�H�޷ZL���`,[ڂW�d�x:r"�ʝ��^mP��I�N�!w6h�P3�
�)j2߹�a�90&*�n�]8D�JUi'�E(�a�s�>�n�����"'c�ꋫ��r��l�b�Lgm
��^�7-hޭ� 2i�y��\2p՝��4A��Be�����y�C����/k�J���������}��y*\aY�2�,�]��|z�pi-n��QӸ.U�T�W ��rVqW�L��f�X�Z�Y"�{AW;x�����t%�1Z�f��D�+3!��F@��MS�47m�^��J�*��rJ�_T�>�v�v�	��Y]����]6���i��^��i{���1��x��	Fjb�^,6�pX��D�4:,Q��<�dr�qŚ9q:��v`\d%`Rn*^�a|�,-ۻOVFs�n��d�
������8���g
{�_�O5}ED��o���V�Y��n�H�_��>�7.���2�E ���P��ז��v)z����[���ga�B{H���#�%�D�Y�=0�7H�;*�t�%������&�3k�+����ۡ��F�74��Pm�u�.FH�k)3Rʹ��vm6��e�َ�aH�u�$��a˸�Ysy�.�*�UL=��P76��OWa�m&piћ�7ݒ,� 3CF�� ��V��6͸�WKv�F�,���{�s��جA�����`�x���6	Zr��t�U��1�k"4�rln�u�"��v�C�v��gc��tve���F#�B	`S��wF��3�(}�r�$>7��Dnw ��x�5e"ʏ<�O<�{D�r�Z�U��, �=�@�[�r�/|Rb|�D����mlnY�%��[ec:VjR�{ԔN��F����0��c �[JLS0Ki��5����f��u1ΣÞhu�4Ȿ�}���/����o�jg���ۚd{]3�=�����<0,���{���>2"c�ŹAQM-�kX�r�t�ń+���k/|Kn����뢈��s��I^�50�Mq���l����C4� �n>�{ԛ�۰��{8&��}:-�	,p]wC�y{]NTV� ��bΉ
藂U~�"������k�n�M��� ='��̅R�ſKu[� 5n�I�s��m
���[��5�ʦ����;9���:��P[5qU�kpfq{�6�`V	�-)9VݹG��1��X[�n�"�t�c{��Y2!��ˑ"泐��7ʰC6�v!|�����-���W�y��a�{�R�Iy��`��hv���$�v�[n2����i���Q�����[f��{�	�3j5J�g	�>A����Q��K�8`op��\%3�u�2����8�����ǥ���EĂ�t�b������95�s_�F�d3Tʷ��m�Kpn}��&�:�:��$��^�q�PJ`�H#1����vp�iG31�V�Vo��&�6�C��h��{y�����{O9�˗r�Q��#�POtn���m� �A��1e`���ur�n��\��5A��9g>��֟GW-1��s	ǝ���3p����&A��;˦\i�3;�W'X ֘�&�-�ۖ\����䛪������6GnM�/o/]I5�7D�@��&=t4s�k�&��
9M�Đl�uj^`������u��Z}ä����2���k-��έB��G��pa�L��y>��潘���S����i���kyދ���K+�/vm�=ѩh%�+gx�����.4�.a�	�@�;@J=LS�R�R�؄�1�eh���n,8�C6���+��"���^�h��#��D`k38c�Ź�y\4�rP3��QC~j!v�=��!/�8;���:�\t��Q���(r#�@L3+'l��u��M�Qʍoel�F���-��D�oN����P�C܀�ᬊ��m�͙M��^|�-�ZsFq�hr����-WuGB�9����:��7A�ja}ۿ[6�y��@�P�r�5^$���N�oQw}���32�6�� ��]V���=޵���څ!S0nW_o_ߌNCM�R�H�4D����O�^��ǯ�v�.+�wU:r���2L6z�r�v��0����A��q�ɔ�S9Mo[�qà-f���d Sw������:v�цQ�M#V_P���#�ʚ��pͼ࠼R����e���;�r�D�����[�5τ�u��W����V��OA_�)�|s�ݳ6A����1]�N��6YU��O"���t0f�Oa�[`ъ�
��ی;�����Da؆��y�� 
4�{N{�l}�b�t����Un�U��7�6�=M����Z��9�H�0�g�7+&�$����&����k�y������k<�r1c���o ����;.��y_G�W���/��4׶��]�5�G��So`�ޯ�Nd[�S��'.��
*S��Lu̷�m��v���ƶI��8f��&>Hsȟ��tl����,`��N�s����(Qa�� ܔ���Yׄ�+յ|�2�}:�2�K=���	lb3�(Yi�p��!��x���S�^��kZ�yG�/{���h��f�:�Oi�C&�����E��� ��͓���;���Д2��������l��Ք�����ܱX}��eY������ �b-��Dm=}���:|��p���J��m^rЪ����Y�r^Hwc:��ui��Έ,�zEҁV�޺أw@�1u�C�ܜ�ۑR3P��p��hԘ��ֲ��NF�s�1B����.�9�:pE���=��;������t #U�%%i�6�iIϓ�ٓ�@�߶�޼�;vQ�[��6d�P�z��e&F���Vr��L)�.�\���t�R��C���jm�BV�u�릩�����7��)��Ω��*�V�c.���ݚ�:��Z\闦U��Z�4��,)]��PƏ)�M7R�:e���$M��4�U�ik͏,�r�b5���6�ӌmJiԮ��=��d%6����H�^�=���[�x��N��-��b��R'��ny͸�2��p� <�zWh�n����J9�|���98e�WA h�7��ߡ��E�U���r�f��Wh�aǖW��`pMwz��U1Sǧ3 ډ�$���ƺo/ZKG��伷gd����.0�V���eqa�XV南:b���+������1sS_\�⮥���� �.K��Z6|��&I���Øu�H
9���.m	5���Zd�H�Y�O��D��>��C(���C� sV
w�v�����i���fo`�]@�=]۷���� i�շ���z:.ل�;�1k�飇	O �a�'���������k�Ӆ�ni���븋���`2��[�$�m��xP�����V1��ӆزr
�g������>�E.�b�I3tD��哨
!�&X�]��71ue#a	������;g�঄i��|Ƀ6��!ܫi�x����:�xo73.����8�y��J�ݟ�L�b����bԫ�[^Y�B��U��p�[�C/*]�S��.���d��/#�oz]-P����֬���M�:n����>fw��h��AXN�Ȥ��*ؕ���yc��Qj��V�҅ZE���\cWy��ʸp7;����EX.r�9�Q�\�#��6k�blG�Z�al7��Xu��>�Q�hgf�l\�6#���ѧ����j�t�h$)]���+��
����F�oA��	����In�IМx��חr���x�whl�׽q����*�h��lǱ-�t	p�jt����k|)�f{T���[���p��]d8p3ǫX���I>O�����#���!�&��u,'q� �y8$"��K����:��g0��+r0.��L1J�:`�ˏ��|���G&ڦE���H�펮Y'Qw,=27Ŧmf>ϫN�\�����Z=~Ϯ��-e�O�1\�F0nJ��'�4�?e�{>X�.�Y�iǇ巑K'z}t�5$�M���rva�5���7����I���p��@�\X
�~=�~i{DU�1����Q�j��f�k@���˺��gb���=�1c�ʞ�:�֞��;{2t{Ԅ��_�L��f��ݾR�;O&G��wh}�-*�*�Ov���3��w�&&=r<��j����|��WC�:F���9�d��Mg�Vnbቭmv���H�_m�+VzI.�\���@}2qe�����r�ra��8�92�{����>����бW���i�#XT^���[yW�eu4�Ǳ��DͷI[1F�kJ��+J�\^�J�
��}��V�yR8jx���/�y]�a�z�(
�|������䝈�<�gD�)��]��L�)�#��\{�]�Xǔ��c�Y&��{�'����s=o�����/�xΞ�
�Q���/%�crta��]���V�����jm1�^x�jZb�3��'	WT۩�X�ς���C�A<�Z4>:��S��w��fT�c���T�Բ�3�v��DY�2��G�ś�����]��Aw���D�o9}}����L1vұ�9�+���\��R�5զV�)3�2���$nPk���sz����+��E��X�ۺ~�c�O�#�q1�.�v�c�.f�&gVs\��a�ѷ�䴮�a��S������$Céj�w�@���T��(ʐ[�8ԝ��s�kl�PQlO�	���;V��OI�n�tЪ;��/qi7j߳��֧Q��Q�ׄ}�]C���d#���.0o.�-[�"9,���vT�[u <�I�{`}�����T���VkxjΪINq�|�޹F���˩��fv�X��K2;��)QCʎJ���&�w/~ɦak"v�'�ǚ��O�Z��E=`��A�Jt9��_�@�I\���ҁ�
�e3pV�\G�[:�C`U�+x����
�5#ٱ垫:Ǝ����ͅ���o\/%�9�)-*귶��i-;����\�1��&�L���h*����6є�c�z�=ݝC-�w+�Ѻ�<���s�{{)�}c���r��[��]k�oxGP����e'�v�w��v���dj�����y����M�Šਞ�*��
����S�ĕ*u�H^�JU�E������ݥ{�YӆR�]�R3�ϥj�^^m񋲝\g.���3�"�Kxz�"�mAh�J���f�X�ެ��Hx��s�R��4_@�E�����aܭV�e���7�(���A��"[����gUӨ2�y�:�Ӗ
���� ��0]%��y:WJ겹�}�����݇%|!BjY+���؞�td�&�p��G�tM��3F�2,�ܘ��`��Y��#��zܚ�|n��9	`w'�k�� C5��<���,7�{y�s�k��6N��6��t]��Y�`�*��t��N���/V����v�]��;[�d\��9ltog0�t�*�oZ��7�iȄ���/8��h��L'���F���� ��:����$k��`��̙ϥ��a��\�s`Ŝ$�T��V�K��c�,SaŽn5YR�Փ�S�!�h�n��Vp&��^�J��:A�n	{��u�~é7��c]Z_��`Src�M���Bʙ,4+ۘ}a�j���Wb����3Yd��Re��u��=��3kZ�P�ہ�hU���`�A���u2H�uv]Rd�-���ɾέF�;䘫�0�Ƌ���1�b�5��ٗ��-��7��ו�j>�|����.�Zk)����MɨwP�yP���EKI;�;zejJ���dɸ�i8������p�Օ5چ��%�3@B�V������t��ݎM:�M���]H-��)eӱ¶��Fk)C��E�F|1����tΣ�u��5WJ:����(g`�q���4���*M�* V��m�B�j"�wW�`�q�Œ�̾���7O;w�B�k2��jЙ�l�<�({�-��K�:h��7*+�~�o���1M{u���Ssj�E��;1Ib�\�d^:Y�҃*!��f��d��Sb.B1��V�R�w�0�!�n��'BbI/1U�c�[�WX-��R�6�uŦ��,��mjv8'��
�8�E���Y�WJ�3���h�<�����}7�Iܠ�< Q/x���e[�|�&xN����d�nw�Tj�@�����<`�ee���:5w��NѴ�Mu��]Zͧ�m�qm��QZf�$�F��YY㏈O�S�U �7�K��u���T�@i��NQx�d�V�̺�ڗ��9x��ˬ�}�rk͕�,w7��k�uJy#�ͤ�ګ��N��3�l@�$饋�!�.�e-���u��y@�"�R�$�J�[�m2�,ͭ6$�WZt��z!^^��;a�[S�L$R��4s��87nK"r@�#G�	�մP n�N�����;�����Ժ̵y��A#nb������l0���튛]gCS�zu���r�"@��a{����s0�ז��Q3��.?Z���{8�O�c���{�
-S���aqh��o���p��w��v�m�9��z�i�I�����V b�i���+2��ku�eG����]&0ķ*�wr�g..B=���4^����Xh�L�-i[1�;ח��������N�
Y�f)�P��_op�D[����F�V����4CmP�c��>hN��ŝƷe�������jh��8i��D��t���Hc���{,�f[��C�t��J�VE2F�<=�z���,m��h�hR��R�iQ�m�1eHww��e��?Yڄ�h3�]��y�p�Wm$pt+��~�:��r���}�vM�����t�n��l�kͭu� N%�r����׋��i�^�C{��
�.m�k���7��2�}����!,fm��;�n~aZ�n��|,[Ȯu�}t6����J�!l��|�*�j��݁T��:rå��Cn��M�,Y�A�����f�GC�	t�&9�s���6u���V3&��+m�l��̄�;ڥf�M4�QBK;j���z�� (p���[��C2�>֍��֗�Y��p���>]=���Hmr�J7�M>�Vk��G#��'9�۝�f�c�c�(o).K�w��VA'D�z��sZo\�u������]rT��nG��ἳ�n�v�55JI���������[ݺM�~����z�'N�!�.�na��A�&�D�7M�"�b�F��ӯE��8z����n����gLyS�L��4i.���.�Fݺ�i�s�։# V�nh�VU��tz�ŝ�'=����DZ�;]��3!���0���[PӒ=Ux)�/Ob�t>�|`�o5n(����uvG;��q��K1ç[;N�N�ըt�o�}5�{��̇�z�0p�΄���=��s�;�>��������U�Q�7��h�ë�aI��.Y��Lo��S�z��$� �jeS�A���g�ӫ�N�mfȣ�C�Q�"�n�9Bop����1��u�
�Ӯ7�,�:�8)'����i]x�S H!u%}��&쳸3�f'���w֣3y�ox��1�&�;�-�p��L^x��G�^6.�?�d{4t]Q��6c� T���\	��)��Σ�T�6�|)b��X�U�C}��%p�$~�C��;�!6����uvd��9S_ �um��9�Y>5.n�*�)ֲ-R���#&m�{S-Fh�hyy�Wn�O��Y������A��t�m�nU�Շz|/��x=�����ޏF���z���5[��ւ��Nz;rϛz;�+�_�v-������ba�w80�1��y�3��q��C�&�ʖ.&+�8׺)���@�'����m����Vu@t�b�<{C,y����q����j�|�z�Tj�p�r붰�'��=�6��7R�G�m�ݪc�Y�a{�ipi�3z��ՒA��
���Gy.���L\�F���Jqgs��Y�ev��u������Xԙ]Z���+�I�t���Sk{�+��X�zΠ:f]�(��MQ2<�+��S/��<����::�Sy��w��I�aN�����e�l��5e�|�t9$������r|���q�rxJF�[�(���1������{/�p�xp(gr���l�cz�|ǔ+�������*$���X.ّ�x�%�\���o{�O��F�so45��0�2�8��:u�>s�H��v�5��7��hG�M�F��>���Jl:R������!x�7q�R:�nj�mNBs�uy�۾VyxsH�����{56˹�Y
�ֺ��M[���C]�f��>�;�:.v���P��V�{*�p��.�X2:���}R�րr-����T�^�<G������Åug�:����d�9�jD���>V�q�gt��Ҧ��-���=���Ђ�v�䴥�MW�W��Fr�G��&o�U�ܳ{.OXPn��?g�O� v[�j�w)������������Z�ì�t�����G�DnŚ��R�o2Jq�}�
)�7�ƾ��������}U^����{�M�B�@��[�1�{"���>1���l����"�� }��"��Km�ޅqnq��R�bs�і�_L;��r��L^*�r��UŅ�^�q��k
�)�R�����+"� ��c�i�5U:R�Ӎe=m���d�<����E8���<�RӶ���Ѳ��2*�|e���R}	��f���z��ym�#�� 'p�Z�襎=��̼�E�u�kE9��t���\$ͮ�*�Cu`]�]�rn[̷B9�O9xnj�r1��\Z��2������I��fJ�~�j,�ҬL!�dqd�Ń3sv��_7�w:wI�reB��ӯ�$깥v'�}�X
Y?9$�#�s�
���z��$��s�l�-5�oz�_�����Bcz�ye{��Ϊ[�ڇ_3��P;.v�n��6�c=X����xoQ�E�je�EsK7�E�u�R�d����Ɩ�X�}A������@�fP��)��षR��^P⚏���7���b���c��r�����]f����]1�(�������yH�t ����бL"8!��߃G~�j�^�fp�e�o*n��)Fև�����=��-V��ͨϙ���/`R�!e�Y%=�GA�D,i���t��r`k�7p��E���и��Kz���d�!x��n�RCm��#=�򭪕�N�@m�	�ܡ�n�Y�l��3z�:�j�7Z�͚��'���J��f=b�3�jd]0���R#o>�k��*�9���6�=BJ��Pvv�n˹���朩��_W��l�a�Ʒ0��f8V��fTQd���X���]�K^kw�Ж����&.�h�=Ϫ��x�N�]X�k�`e��Օ��=�G�i5���{D �KmI,��W�Y��Y�ۓ�c$��{؞A�ޠ�n�nz>}i��B;�of�F#Ʊ�چ�R�٭����^9Gj�7o�/���1���Y@>ɒc��f������CźN���4q�x�fe��� ����Y�h�}�k7<�ONxΚ��+�ׇ�5Wp>�{���Op-h�^hj�%1e�Ψ�e>p�B�R����A�d:Lu9i��x������ѯ���}���\U�U����Ky[܊�m�r9rmɺz��M����C��6�J*;�#U��
w*���h���:k�fh| �#`��\2�5�~̗��ԭ��Ð���c�e�*Vb�;v�v�n�9 �|X��S��_�*��r�NYtQ�Ch]8K��� ��Z��nV�Ǣ%�"3]�GL�V��6M�N�. �m�a�r5������@^fރ�w�6�C��m�������Et�׮]�,�|wԐ*��3ק5m�^�.R��%c�%b�K��C��y]W�ᛮX[Ɖ���R�k����f��Z�K���"��f]�ٹ `��K�Đ9]h�W��ε�Bs�'��|�P)�f���l9�X��̈́����7�cӂ� j���S�q�mi.�f������؏q_ֱRᴇ�`��Bҷǫ
2@7�䷦�U6��b��IXT�qE\���YO�G2�+�Ёy��<�|Q���"GA�+E�qo(J/X�,:P��综��^pj�Z[Zh�tCxm,�L!����y�#���u;�AVtn���6t�[�mM�s�Eu���*ﬗ��-*�55��w��l�آ�H3E��:)sį�P�C(��q�鶄����V�}Eq7��<罜�յ�[F^�wK������q}�k_\��������U��Ĺ� �<�:&�,WR�C&u��eK���IX�x�I�0v��j��UZ�bؠUzQ/��@���4n�3�C#\�j�F<�Ŭ�!���e-�n�o��7%s���7o������A�ލ޸��x���{ܳ7cV��Ԍ�ʵB�)ъ]�
��y)��D�V���Uh�_2�b=�Q��]rk�X�k7
���I����(z���7��e�Wce�8q��L���⸋���z�R˝rνVY�u���k�ʒ
��WK�="�'6ds����}�I��BtfLc�h�Ulu�L3��}�*���_s1�i^�drZ�p;NF�sFS�g�u�u�t��Y��U���aͻ}��B��R6�*�{��{N2F,g-]#*���
]ք)L�PR��ᜪ�Һ�Zd����Ҕv�>=|UL=E�Zw:r���!��k����֦X��TWkt�sn�liˆ�N��_'\idf���&���fm�y��MAzN���)�ke����Ijα��6�n��E�ya�~{�{���i���5�S���v4s�i����u�x�74�.ы}c�<�cC���
�Z;�>���w��k$�w�9�^ŀ�W��mg^���z.������t�T
�K�yٹ��o$A�t/^�#t�"�sŗ|�5��3f�ˢ�8/OZ&Ћ���=�ߑ��%��%v7NT/	�v>Z��D;�"b�ϙ���q�kO}� ޭ�N[�C�b�N\��<��*&W5:Q�*T��c���\j�:�{��������̏Sn���`rý�N�U���3������[C�93V����<�w�!Z��vȦ���u�fJ.Wn��Z��a@>b��\��!,ä�\~Y��ʇ���=S[�vd9\cBU�rj��]l���Ϣ�x��xwk�o�k�4h^cbE�9�F�Ò����B�� ':ڋ5u�������>�8Y`�H�������gJr �^�
�{�v; k��Ϻ���-�d9��F׳E�o���v/�������2��Y!u�]�	��Qݠh��XX�����#�BR-`0ծ�f<��vX��� ��2V"s�<�*�]�9Z�c栬{-ui�֣lw�S��A�2 ǲ�jB^-���(sDka�����7��aO���Y�Y�+.��6�����S�k��d�O%^vv&�u���êx�)DR��ౖU"U�c�9^wN���SKx�Ů;���!P%�p�6�u�F���83υ^"
���ŗ!|"��	8ҫ�mv*Uo#f��9o��2��J���W��l7��:�2�ؗ��w]�r�$�	��pvY�V#�f��r�	z8���Ke�!3��1] jm�t+(�w�e^�8�
@oU%-]*ɢ�$ޝU�6�E0�sO9v�H`U;#P����7p�8^\2�НZI�^��v$&�|:�J��/�a�m��<���t7�v�l��h�'�mR���k8�
9�tn]pˑ͝h�*�Qi��K_,�[{V�|��2�=��S��|R,#�3Ba�#[Q�F�0/�w�5F�J�it�D�$�����P����O���)�]N�Wֺp�ʷ�A�k��Vy>ӌ�����,ޘA�YfƾU�(�I�\U!�m���WO������:ԣ�R�Ч4!k-���֐�*��l1:۾z��*eV;8�3謖5|eX	��Oh��b�3Fv7���ݩ]@�\ܡS��q�^5ЎZ�֌5b沗�{U�b$U��C=>Vrb�ԋT��T{�)�1�ۖao�޺i(�]��y�Lbw7�怑����|Pt��h_R`�#&ő[7]�BXK�F����Cz�\}:��[�W�^��F�s����%�4L��v��j����*�����+��M6m�^,=��L~i� S��{�ɨ�	ӌ?�AhJ�E�s����p�h��td#'F�QY
Wk!,�zd��@jm樾VQW,I�n,���Q<� Q�׼	�V;Ym�)�)���c�k�&�,��G9Do$���ی�q����2,>>��oz�:k#z&�k���r�7%)�4dFe�S�)ݑ��T��toO�4��8�3>>+ ��·���5{Dӂ
uXt��� M��hXp�R�E��7�q
���.�V�
�%[�z@�[a�����wS�.(p�ᝃ��C7�9e�
�q���g�V�V�N60�>}�r�i=�]�Ƿ	�K0���%�hRK���m*T4�Z����� �����Ŋ��5o�ٚ���T�9�+�+�X�v�fAF����� ;��#���1�w_�v"���6\�E)��T(��D�W��Nzq>�rd�T��S�6�æ�la=��=
S�7�d;Z�dT��k7DJ�)�l�_e����+�a�.W�o���N��u��|rT��ĄRw����C�N��r1��4�u�bY�/I~�F[|O@�Xp�g����+�]����.��f�
�a)��٠> �|r12��2�2���t�M@��vgH!�HFaW�G�yX��Lt%�+;TQ���da%%E�>neM��ǳ2\��N�ׂf�)^t���3�:BJ���Q�׳��̠�,,s�Ԙ;�Aڲ�6���f�����S��6u���a�86�hgkC�fS�"�8��ZSe8-�
�1W!<�y�k����YN]���x޸Cy^ L��? �?o�h�t�Z魘̦;/ȎS��I�Cl]���]��W�r�ٺ��H1����IԝDa[��D���c��&Ը�
��E��B�3Dlc.�T�r0�'�ґ�F�@����� ��'Z$e��_�1p%��s���k&X���P���=�o6��˩�th@�BەwX�۩�W.>ά���э[�|�L��t���ُg��M�;f0J�&v�Zo^�pѼyr�2��^tͮ�d�\�On:��ƕ���QJ�v�'5.�7̎�mL��|Rd�{�hU�}�ШbzVa��F�@��^� ����kb�ş���>m)Co��]�:F��+.ڣ�-���L��[�Y�P��D��T��9Y���3��it�]�7�z�h�=����=�ww��r�2�}.�,�#25Ɋ�_�G�)<��d��a�Ǐv(�B�*�%��eo%*y��\x&^];�N�+��>Xj�n�:�(��>��XV��
�������H�
���e5[*%qh�z���!���y�抨9Ξ����J�'�/l*S�р��sgd��.�[�gm��=,cVJ�0�Ge���ђ��}�L�Շ�EK�Օu�/���^�p\�"s:)��I�:or�3��䨞������aȅwV���u]Lֱ�{ �z{g`���z�Cٰ����=ygm2���$��mX�z�S��Y3 ��@��y���>윖L�tVd�rQB���4f�)/;�r�k%XޏНnZKp{��լ��
�A�K�e�o@N��Ђ�G�r�HJ\�:0͢�okSpT�x's�M�%Iah�V��M��oohF7���-n�(�@'+�>�J_ Z�{�J���t��Y�:[)ҥ�{�dxI(Y�4n����('o�C]_j�ݚ�=�����螬�:�Y��in�!ۡ��rRp��%����}�B�f�;mIc*�1PN��cV��,$:t�<N��=�.�'ڼ܃K8^#��|��id�5Ӷ���\R����/20�������1R��
¾�;^a.,��Z���G8�Q�YթY����S�)�@��n;ل�m����^嶬w�0�nœ�l��wDù��h���L��d�
��{�	���nM�b%�w������ׯj���P���x�p�����A��.x�Ͱ�P�[[�.
�[D�V�P�ہ����E;�)Y`�Ν��7��fK��3.�=;e[ԉ����ؾ}V�ZD�P��'�3$&�5�jE�F��7�Jt�}7щ默N�\E��%rPM��%e
Xk��̩�!Z�`�� �W1����0�н�w,a�}1M.��-��j<�aq���R	���@����f�c�@���L�!�Lu�8h�9nt�5��s��4�#Wh�$��Δ���Ń1;��et
37��Z�[���\ބo��YYY�*�5��d�G����طr�(n�p�y,|Y�iǸ�L*��lN��w��7�uޝ����H3cnZ�����I]���}�1�V�.�3��׾�7['.���*��CI+7M�a��'RhLJ7v@I	���[�����3EjG�;�=7�T�=�wb~���l�wl�@¼�l��X�3��Ilw�%	�Q���gS���H�gHh�풗ʷ7c���>z0h���K Юz���S%���W5�X!q��΄{͙uw�*+�k�v�����A3��a�I�/s�5����'9A�NE�n8�΋۝��l)�i�:�MOr�@�L��� -�ޠ�:�t|[,���7���LhH�7��B𤰥��s����/��jV���Z0��8�������>��J��������5BX���*����ؐX_k�v_1��G��D:E]�&#���<Y��]�3�3Q$�72��N/!��]�A�-�WK�
E�K��]fWlN.����`�u8Q#~h��[��D��'+��?_%�9���̚����y����Ȟ��O+G-�[-�:!���Bh�2�J�fR�c9�l
���2!-�#��<nM�Ni��=�vջ3�|%�����Y�Z`3���"�)�"y��Ps���7�I�fZQ���X9�8f����0��&����N�3�禓����2���ц��=�!|�Ȇ�9�k>�a�g�Vf�9'Jx��*a�.,�{˅YG���/�v$C�/ClMs�Z��.�ۤ�q�j=��3��� bɣ�.�L19��T�.pt��ӹW�H�)cn��$܍�ɉ<���ouE�ujvR��"�����}�������9.{ݺ�b|����ϣ�ce����q��c�P��r2�w�X�E�.�i�`��m��L��2��%5�r��:�
��`����J!`��;h@���ofr$!p�NE%�q�X��t������33�ϳﾹ�G�vN�7}�}��.uʗ@�5���8���3n��QsV��#�bxg��R�p�}�1N�-�7�{Z��@�#�H�n�s5���H�9��IF�/�m��u摢��\d��c�u��-mY�s��oM�U���o0j�qX��f�A/9�=��u���Z�A�� f��Y�o.�a'�6�j!�Ef�<�*�Q���F�|�t�	(S}?�w�eJ|�l�*���e��v�C7/ H�^�E��Z��5f�e�������+�}WE�"KݭQ��>��o'���%���N�b�X�oZ�WJ��u-xK������5��.�S+��E�X��֔����J�z�7&�b]	3�d��z���7d��%��2��͐�v��'2�e����bb޾���6d����k+���:p,YJ��(W`����q�E�MZ���X�T:�vAB��q��[��T:-S�V��*�*n�m���m>.�=������Dqb�O'9�Ùn�V�J���M�2�y���z��'���R��9��S�`�Vq��-{3����9<��ɴm���,��h%��}j�A��˅��K����Q�_*w;��9��C�q��A�p�}�v��7Eќ7'�f����Y�4�,�tj܉�����'tImol�:�u7n}Fcg ���>$�%F��+"8�Ɛ$���\��ʨ(�tH+��Mܖ��D�)���E��A�:��]�r%X]<��QNL-B���$�'Rs���J����ivjL��	�(HN���p�I��������)̎u�.�AL�ֲ��4!��U	�"s:gueS����c�R�.�Y��Gwv���=K�:r���'*��EP�RE�r�s�s��E�!�'QΑ�w%�����.PTNT�(�J�$�@r"J��L�x�E9S�:*"� �r���8�E�3dCHJ#�d$�i����a�:��
aB�r��G
L����1PJ�/!�\<�# ��0���n�F�t��y&�VH��uݺ���e�˂WN�~�6m��t���:
[a�,���4��׹͉NWJnU��ݘ>�N��K��U�Q�_��;L�+�"��Nx[�7�)Q���зk���`yã\��u��E 7�����������OY�ܲ����r���9������ �%co�@&JI�ZN��l1C����Ϗ���Ë���V+ҝb�JD{vV�)�z�ĵ�_Je��V�Qhd�C��)Bi�@k���ah�z�2��JZHq�ݛپ�1W�r��PQׇj�����1��
�����~ᚖ��G&lU�6��3b�����%z`��rp��[�f� ����a%sb&NE���;�*�Zp�h�Y^g�aG��W�=�SS&�����
U� ���r?q�~�^�mZ���J��v�A^���mUf�΢ŜzhNQ{>��Ԍz���Bi��|0�l�dM�ګ��N�
b��zi'B�؏�.J&Ń�πܓ2���^���-q���mT����鸷Ë�`ax�ys2�xt/�d��^���SO&}~s��<ߚ�^���k*�I�f74E��l���w�{_�ͫ�TN���⦏�Q�.���>%�f�v��٥c�:�E�aw��pL�H��^��ӇkO�Mf���s���D��ӝ��8V��9��i;S� @�ս��B�}o=�6�"+$p��OVm+���B^"ǵ*�������`�|�Z�a�b��8��L���:Sw�u���]��t��9�{鮰 �����i�f�z��5�����R���1�;>CV�s�kf�K�U�T�S�����`c5��Z�c�5�N�~�0,޽,\^��W<�fv�יw��5���>Y�q|��+@.�z��޼����fW�7\�`b5�x�����Ob��fJ@��*`���\���m$zm���L%c��;FQ"dʺ�pC��G&ɤ�k����1�H�4���d�H�Q�G���TL�-l�:��=w��խW{fI6��&,�k�e�>�o��#ώ�)
`]�~dR�puD��d��yn��p5���B�f�Ϫa��R�
tǭA���rt理�ǵ��`�@*�h-	���y��t�b>�w5c/�/Vi?#K(��E�F�|�Տ!	bgH�6�"RN��y�t>b;lda	��*s|\�B�H��s�a幷��*���WUq���쀽�J"[X�׌2��wh�x��4o�YJd�^�n.�&º���3$ۺTt)ut�2�a>"7N�VJ��i�k
�P�(I�,��)�s��Aқ�Ӌ�U���T鋫�l8�O��:#��<	�΃-Mט����+_<;��qsKr��Ww�-]V�H[�澧�l�#�61Sʬ:�a�5g��f�/k=}��X�h����T�5���ί9��
̢'C!W1B%���5K�tm�b�g=�gh��1 ����oՙʴ�c�8��2>��[,����8e:��6~5^�Dtn����-V"��T��?kc=�}����R�5`�}�Ļ���][�����X�|��֕C��+gm�m�h��st����S�a�ه^�4U_>Po֔��bCʿk�k>qO���wv�6o9Oe����\-V�c/��EU6�p�����`c=UbPW�{o�eTU�}�?�F��g�������M�A(� ���������$N������/�lj�Z����REy�ז�}��V�SfF��z3VR(2�*��_�\֩	VH�`4:^HV����6��tnZx%fīu�d��^�P�>g̕���`s�P��	�AU�X'e7@c��fz�9��*M�nV����b�Qj`�+�������룎���W�.b~d�����sa�h���$oE0�娻��/?=�ڊD �'3�̀`bi�A�Ov���&{1�*�_HcUk��2k�vV>䲆Ư����PpX{}ץ*��j��|���)�;m�%�僓�o-~䊱*�V���5N�>r]�ȁ6Ө"�I�,�t�T�D�A�|��2�����T��_
�h\�S�B����U�l7���S���J���]a���k���D\��ۮ�O#-^��&p�z��o�;����
�(��]|c}�+�S����tV
2[Q����ӵK��u�����"h�b�B7��X�N8�2��4���ŏU�i��K���;���u��ؗ��e�pҁ� e�tS0�4<�D�YP�Z��L0T:�B��(2�հ�jRwu�u\���A
en/}� ���eJv���|�f��J�RZ����2*E�b�g��/g�1'�gI�P�[�>�����Z���8 U!��^�vUw�5�i�~��q�7b���yV
��t,ףHe��7Y�G�� ˭����ky�
R��dˍ���w�*o�=�a�niz��W%�+�GB�/��`��bc��:�^P�թZ�ٻ4m�Ζ�ױ�(���zkB����r�p	��|�.��}�"O.f&A�X��ޣ�:��۬Oe����꾲�t~Tz���#ά��L�S�n�4����.��r��&1���@����9��O/e<D��rU=�Cf,�:ΦDZ�|�.�4�fT7l8��u�u�sG=��4oMs2붰��6�q�h�� ó6��<:B{&N=������s+��/]C�~{��c�g�,	��hc�(4����[ٗu�w���i+�C=TZQ�9��7!ak"ْtK�PtWکHoT`V�߲̉�o���*14��{&�����6�{�)��u����&s,B�Ll�Cjt�6ʲ ��/W&���P��T�we=�4_��b�ڜk2�
n�Ɖ��8BA�m�@n�,�)�����wi�:-Q m��tFEQ�F��=
��MŇ*��˪
��U���v-��է�'�IȗJuо�ws��F�Y�eK�O�e�O�F�.�>��.b��\@�W�y5i�1����o���2�@�a�T �2���(�<���o���k�_��WL����ۗ�09wH��P#�"ө��܈APX�uŊ �J>�ZV��R�����ɛ�.�@h��¶o��6�����׮�yE��ڙm����4���#�o2I��w�j?`���G�įL,,/����TW'����t����=�Aɸ>�PH�W)6ވ�g\����Y�5�b�\K���o�Z<��[�i�{	,��ege�.a"-������^lB�;��s�����4a;���껔�+�+��~&z]�@�O]��͢t����ݮ�f��*(�żx���a[�rDb�p� ���BvH�Ϋ�[����vZN����W�`���s1�H�iOa���I� ��@^����+�ߧ��^�:.�ԳS���a��h?o�/F���F�X��ǉ���Y��xe���X�k�n��(>�#��f]�^�v�a���H�O���8e�]� ������fR��-5N7���'"~�]3�^}u�Nɡr����p��[�����PQ<�6�+x2%��PPh�ˬkUn��y!k�%����[�v�D
	'�5�N��(��lf����y��\b��^w)��p<�x��� ����]b�Մ=�ӟ�gB�t�QJ�K �k�Ʋ��D�LV���tx�^�R���K�����~F��g윍�G*XӞ��m;��S�3\K�V6�W#��6FF#�&)�u�8��P�a������Le��f .E������U
�l4�x��w��ȼ҈�{�F�^P�?�<N8E5F׋5(S��JǪ:�փYƼ���ŵk{�K��)q��U��3�#l����H
���vp�S�SۑAb4ʮ����U�E!��z�o��(KW<�hus�ϋ%xV�ŝ���՗;��v �b��ڑ�
�úp��i*����[���-o	�������"�E�R?��
�n�h&M�#:�{A�#$��.а.>=�mUƭ۬2|E�6�w)�k[iTW@MUf�NN�q�[˴��*����U�x����`����@aJ5������h�x�uz)Vi�s��4)k
i�[��B��e
����
58�� �l� �pk5�M��ž�����!�qM�y��z�W���-?�A���"D�A��@,E����W���m�p6߄;��򳷆�-Lg=y�OS?��B(�6�� 1ELgPM�������Z@�|�#"��$�#{-e8@s�d�Y� qg1T�3Δ��陼���M[x��k
L� 
Ft�(6�W1�����1��r����6-�qޕ�*F&9[��g=^�^ڮ�a�i���԰|}��%���t��ֲ��ij�f�{�jl!	�[�y�l���Vuid7�%�>�HV�^/�s�N����s�k��o�ZW2(�1�Ӛ�T銁����~s
X�Ad����bCuƘ�j�k����^�}�m���p�V�ų5��a�j*���U�~��3-t7�A\/Z�������ٚ��я��
7%k�鹖|zƭ�<���p��}�թZ�/qP��_fD�RAR�EX��)nM/K+{Y�kf�Auڌ������f��'�Rg:�Պ����,�3e�W֧	�q���)wRST��=B+w�j~Ɵp�y�rm�y�mv>ނ���.)��[Q�;�)�� �l�M��,�\�엍: ��8�\��vZ��\�W�������+	6�!�^Y�l݁��>LVB�L42���__�c�%��D���C��
�Qءu{�lU��Od��>�Z��o/gs�k_���֊��#�3��ژ�f>
�u��	����=�7n�Ô�QW�',�խ�H�2�QfТ�-c����/
�^n��'�@���'S|�ޜ�M;�R�X˚����L,mQ*�8�P���PP��Oe�q��� ;������{�z:9T�*��Q��tSu��^�G�y���
���\�;Ƙ�/|}GS�Q�����l��*�u'�
� n�i�>�G'���[�y�S>�~E֚�EV*�<�3;�ZE�1�� 3h���Fh�I��/;�G�'Ug�n]�*���˝���?N��Of�z���3�C�3a�+!��.����ҕD��cӖ�Ɇ	�L�ߦxe�[nXW~nB����u�XVn�h�z�7T�O�ʅ�9�^��_}Kp�4��D�<_��~�t,ݐ��1ܭP�YV��T�.��;��z���]���i`raIk�M���5���ᐕ�v�VM�wN���rW0��s����q��T���/v��A�=�^��Ҳ&@-o)rMg@��/ -U�>��VDMD*��Q��&Ҭ��-��
���A�e+i]�˸l���^��HՊ棡Ƥi�K<o<���Re�?�����W�^	w="����I��k�?zu����`|;+�M�E1o���\���GB�/�Ϲ(+�fߚ��!�mI�v��k*�8Z��hB_2(JՓ�5�
?�u �`e?K�v_E�݋j�kMi��ĳ=8LN��93�9]Ƨ@�1^��O/
q_���.f�����0&�>�1�gt�6Y��}ҡ`�*��CI�p3��b���,4�7X�eN�z�/#�t�/=X:���z�ze��W@+<���J?a���mz��Fk�;ڞ�&x<4��U�"iV�����q�ۜ��(x)֪\=���cE��,ڜk0<�պ`����tK��)z�v�yՍ�V=�~�iP��9�l��Y���E��jw;&�3,*��o��c����Ai�����Bp7�
8��1Ѐ�����'�/X'�#t������(��}�V�L�5���$�c�5sc�~�09��M��$����m'A�5=j*P����4�QVHm�!�^-�"�jAD� 9Zc����l���1>`ɒ�
�cm������� a����Rؚ�����X�^\n����m��D��#���vr�7��f�[}�Fuq��c�ѕ���L��{�p[2�9K:u�xmIo�&�Ws*��`�Z �DQ�@�|���F@/���-�.}^��W>[9�Q�gT������R2��E�N���Q�����ģ[�*�U Ca���Y��hx�i%3r���j�Fl�����
u�Z
x�_��. ������q�v��ԫ��~rW�?u���0�Lg����v���įL,,9�� |x��t�� �(�h8҅����S�֟�W5��w&�p���>���W]��{뻧��RC<�!M�<���o�zoAGݺm����US��g��3�쿖kmK�P���)cH�g��{!��{�b��ɬ+�Lt!ze�}H|���,u�P9L�xIwI�L�����;��\�:%z|�V�l�[,�@��_ �A6���:��9,���>}���H�J�&_k����~�<�6�=R?a���^%\=t��%ҁ�C}�>��O���P�5·5�^R��tݣ�ؓ3�ɐ�����ݎ^ �X���X�4��n�s�����'`(3{ʄCŶ6�cg��9�ѳa��`}!z�{a�ҳ�܈�ǹP˥ZPM���	qh��ح�K��-ˤ�	m'4GFW-���m���w|�1q7հ���8^N��ՌkƇ�栧w7� ����0^NAt�0f�ZVq�L���36��J*���K�<w�^�p�v�D��p$S ��ꂵL}{&��R֖J�y���Ŗ��P���h�8�y��p�}ܯ���£��,�wMUӟ1�����ƍau����8�N�.�wn��l����Gl���Od�|�`�,&IOw���9|DY�-�r����͏�������{fx��$�N�_&���չpq���6�k\k�fӶ|+��N�{��V��w`1/'����]f��8�٫�X��\{�z��qQ���f٫׼s(�z�]3�f��/��]G�g�2�48J����T�B�*���+`�/)M���� {�Q�Z{Ǆy\񂕅��#�^��/��n�ж���.�n�0����n�L����Zm����U�߭�}��j>���of�Cr�]�7Y5E��fn	3���.���� n��oF�qY��:t������O;n՚U�3>*
p��n�Z:�Ϋ�WY�ʫ�!u8�G^���AV�c%{�ӕ2��j�ū���t�&�uN�n^Qz���&�]S;� Y4q̮���R��K��';k3gn=�s%�]�w9�Be��V�V��1��p?w���{^�D9t��w���8ֵ+�>��NWSQ��S��zSՕ؜B)� 4�@��d쏒���!�8��� �Dl�):[�3�?o���7[�;a�ڃ�o�*�}��ܔW̎�+d��	 �+E k��{�jۀ�ƌ�I����x�O\X�,'���I/��>���5J�7����A�#��S��u�nY�������}F��ߦ���*Ps�8��8�F(V�Eg�s���Ƕ���ҵ���������\J�����Z\Ł�Sk��T�B�,��,���Iwp�]p
�M���T�5�������rSw�׹��*0\�]�g��j���ڻ�r%�,^s:�JIGǦ�/I#���x"˧�������5��v�V�X%+���e'G���?h�����[��eu���I�K���ru=���}��V	:���j��h��]gq(��E���^8J�$��Us��a�Z}}��#c�X*U���l���{*���\:|ӽ���mL��u����[�Zg�l�K��lԳZ�yb��]&�,��,��;jrC�u�m��nN��C�v�oc{�^౴���ƥ���M���i�Y�Ú35��͑[�W����3�(�M���\�9��xB����u!���ա��E8Z�-oWכx}B�j]%*������0+ۋ��)�ɣ��G��^7��[�y�{��1��Q��*�\IkD;���}W���u
sP�R�	���WV��Z��ahj��9勨ӹ�Y媖�pz͌ю1����|��_q��I*��-�=f`A�Mu�
�k"����J��aFs��R��4���6iQ&QNn�̪y������aL���K�l+�\HC)�r�=мI �$"�@9ˊ�3u�L�.DN(�94��eU=H��ˎ�Y,	YI.\�����9�B�rJ$�=�\֐\͗
�P�s���n�*8^Bp�`���L:b;��cB��uS�f���O$��e��	2�TR��wg��*E*jFgw\�Uk�+:e��,͜�m9B��J%%Uwwn)&d�T(�� ��hiU��ùӅ
OWQ�2%�^o�lV������o8�]b\8�{&\�zyvU�9r�S�y�s1��������{9�}cO�N���_�n��x���O)�SϾ�7��7�����@Y��=��������x��뽡�I^���n� ~K��?��U�HRO>>q�7��?��f�nj��q�q���{yv��/��5�mC�r�~�M�	ޝ�߼��pyw�i�~����������ɾ����p���}O���y��<>\�=|�ߐ���=���A�������<��^S
{��ș��ʯ�l9���_z �A�ϸ?#����s��NM�	9�������;J���𛐜]؟�Bw�����9���|�;r
R�kմ�ޓ���}F'ӷ���ɪ�1���N-9v�G�X�X����3�{;�oo;Ͽ��''�®<��97����;����x|8�������]�N�������{I����+�4�wޔ$��?��/חo	����]�����ێ�z1��%�y
���6�8���hnn��������|��7�<?\|C���V܇����x��aw��߭�?S�a~�݁?���?�o��������I�����Ǘ~w�9Ih��m���l��²U��9<����H~;�����'������һ�i�={���4�O܊o�!�5���|�ɿ!>ݼ�G�789��;������}&z�m�&���}���yW8y�4>�E	Ϯ.���:oC�&��Y��vP�����}�վ�������<zOI�S'�ߎP������}��.��ې�o�}O	�!'>�(Rq������&����@�@t|�ᘎμ����e��eQoƳ�}~�99�����.�� ��+��<+�w���Cψ��q����8q��������y�����Xl�®����ސ�{�?\~C�� 3Sa���1�!���ē9���J��M��C��뷗yW}M&�G���S}B|'�n�0yM;�Ǵ��~�����N=}���yO�WoG~�yM!?]�'>������O���ǟ���]���Y�Ͻ#@�23B�>M�Y7E��u�e`/���Ԟ 3�<㛏��hfe������<�I;x��;˿!�����P?$�}q'������'�����w�ӷ���{O(ri�������
xC�k�'���m�4��I޻s	t��TH�J*��FŶ��m�h/6`�k���l�Wڊ�ꙑ���щ�l�J)%vn��*q�u�d~�Ӌu���N+�ו0���}70�c� �������4�_I��D���ݐC;e�O&�r�Ls�_4�y	�Q�+�]G�;�3)������.���Ͳ�|�p�=��e�r/s�B?}^��HUxC�������_��ےM��wϖܘ_�=������Y��x~�����O�?<x����>���|���S������9?������ߟɹozz��ɉ�T�����3�ٍ��O�}<v�����Si͎M��ϫ�P���> N�׿|}q������c�����>��>�z���m�=V���غ�)uєn�gX�6p�`�?|���o�i���9�S�z<����NӼ�_|��_i��I��cü!�4���ro�O�~q�|�(zM&��S��@]��w���i�>�|y28�N<��K'`mG6�Vƶ��k��P��f�Ky�f��#�����Ho0�m�<;x~�&��<&7��?��_H'o����$��v=>��s����}Bq������EM��Tp�J��f����`�X��c뾧!�4�On?����$?�^��>�����n���o>>�C�{;�'N>�_w~�þ�I&��݃�a};��8����ag}A���\~O���T;�����U�خjPo0s�}w������<�<�����O�9�׻s�Ă��������xM�	<��z����ԝ�;��	�o��^���O߶}e7!�����y��yw�x�`�v�s��l1!(ܳs��9�7ϑ����ӏ�w����z���������O��]��#��7��Npz�rē!'���;~NC��{���= rN�}����_)��W��w!���,���z��V�bvc�%\�� ̃y ���<x��&�zO������ޝ�C˾���v��V�o�O��x~8'~M�>ݼG�����[s�<!���S}|y���zL/ |������>u�U)�}Gr���q]A�CHft	$��y�þ����;���Ԝ|O~-�4���/�����+�&��z��<!�4�O��x@�������I�!>�=�x�89ރ��z��h���EO�Ζ�me�^�k�g��G}��$���מS
a}���>����Yޱ����P���s����S�a���>;�x���|C�raO'�}�n�'�9ǟv9��A;�O���I��[]��@fd�glW^\�HQ�Ϋ��n6E���� ��p��Bí¤�1M����k�r�]ȭϓ��;}Ѿ�ʻ�{�f�N�}�*i��>�F�����7r��j�f�r�J��ۚ�e�|x jw%:�;���٭�30�kV�J!w;On�S��P}D�	7��9��~�[~�|SH~C�s�v��<�����Į<�>�xt��w���^;���;�����|�|�{O��0���>X��M�<';y>[���t.�˪��R��Z����/ܗ;���a|8��'�߸��q��N=�;���M�o�Nӥw�׃���ߐ�������P��w�~E9����yq;�r}v�����ǌ
o�O�S\�5�c��3 ��<��v%w(�¦��m����k=��<���Ǵ{�<D�f�t�"�;��L�[/2ʄ�`��0{ww�}��ؤ�Pg�x*aaY��]���n_��;��r��ƀ"�Nͽ��U4��g'��b����d�� -_�����Tì���m�P��N�^�*ڇ޽[���D�O�	8*-Z~��xQ���s=��^t,�%�֖x�:�!_۾���V���|��F��6�3�{TV�M�h~�Dϫ�Êѫ��_Ԫ以d���t1̚$M#P��h,m���*%��|E����b�m��J�˪1�',f�O��H��ٻ�3{�xQ�W{��2�9g!���<�gٕ('�(�C���M�Ή�rߧHٚE�%��uV�G
Y���a(͜��ٹxXj̒�R2aA�o^Y���nֵQ�e�D�	��F�e��F�m����7��`�)K�gq�EL�\��7z<��;��3:��"�;�l�<��BWz���&f&���=O��e��%'�Nz�3�^��kNq;ŪΒ����q�%ېazC�][�6�H>���6X�-I%*oz�����4�ϼ��[k�-s7�ϡ�O~�w�%�&pY���y'%����W�>�Or���6�V;�_k;n��g���Y�@��t�kW�oUJ�����#��1mu{Zd��e��ɭ����UO��#�;ں��Z�&�ÔK!U,�0�**j��3{*�C|��L��C�: d$� NʇG�������բߊm���E.���>����]���MXR�y}��_y�&y[�����o̫�������Þˠ-��n�K9�^Ӯ�承U��~�B˽�
�`Gʸ��~��w��;�F�V(��w��z���#�pY���k�W>�Ò��kF�{������h�Ol�ɍyu�v������Ӟs�S���6��0�uᵉ^�0XX]VE�E�*��Ժ�wa��k^df�ڡV�RO��ܰ������C�V=�������Ld���(�@�{�i��'eKV7?h3 ��p�����]z+��{K�Ɍ0���v�ž˵�,�>7K���mGtaK�S�}�m��vvԕt��wr����C̹�kzu9��T���%+:<�<�#}�KfR�z�Zǘ��ױb k�����ᝋw�<t������[#ul��u�k�w-�J�ʴ��4"X��7� <�$��/31������s47��1����9!Ze�}%�T3k2H�LL�%�N�WOtw��+��ޙ��H��^KO��wEzP�׃
����s銼/�e�����{X���\�U���%��֊>��`;��E�0a5��~�+\ RJ7

�}��9hI��̕�z�[G}��o�S�l͖�� �|�@��OC�T#o��k��Dt�h��+�f����~�
��w�\0�>�����=�T���.�`c5��	��6���ul�=4�*� �/f��$� ��ACa�?+�ZL5b�f)T��˭~����[0�CPu5^���<�S����KL2�ۤ# �� �B� /k��w��΅Pm���4Uy^{&x+��+ݹ�kF��o��;D���?��L��)�]{�d:�ct�|�	�W, �^���w����x���`��ө�S��!��ô�{vg�L(@ͷ��-�[2xe�N�&1F@��M�<K�TХ�)��nc�(!e
����rt꧐��p��w��,��4|Z���TdK�\�G��]:��q資{/�󒷝��m� ;N����5���-!����|3�&V)��QZ���>�;F&y�]$���0D]���^�3�0�iT��_hy�E9ܺ�m&���2�=8���]E���:j;�Uϲz�]�z�h:�C�qM�vi٩�X��^Š�J��U��xg���9pF\�-�hL��l'*Y��d!��z��p���c?g��0��~5H⽪C�o��P#{�B�W���;W�K9�(��	�q@���G��*��a-5���)��^�kӻ�Rޠa<�$������W�5a��&� ��єA�A�c%1B%��Ъz3�FR�, �"�C�z��Ow/L  ���XN��!��i���]\�y!t�{"���o�v3�~:7��_�!�	�҇�Һ${���U�`fEL�ZY�%�3+���_�Χ(�����:M�>��޷.s2��u��%���B�������0�x�Ad�����+�1Wug}���m3�U[����ɔ�*&p!L�v��P#^YEU6�p�����e���=X��V>�j4��t�,h�ɫ����`�[�C->���Y
�8T�w'�PZ�;-PwO�Z�o���ѽ�Be�V���U��b|�-GC-2��ЉS���}���1!�ht:kOF��rw�֙V-�N�֜eR,:���)3�� �r��	�]0�=ܢx,���r�.ʩ_
	� J��Za,�:;K�;"�r�C���q��\�G�3��3���s{W���A7.z0�2T�[|���w �v�m������Ma��[u��_R.�J�����b�b�U���Z��]gs�uK_���*���~3=0C���Rtcm��60'-�+W����.�I���7*�K��`8��h��V�_�k�Vb�������A�xS������R��"�/B<
�h�VfA�W��|+¼3�>6^_�����+��ݻ�7N" �t���<]���E�鸽d|��(�����\7���{|���ۜ�N�pw0���\Rr $h� -(���䄘�jJ�����NO[=n�C��}3}Y����fF3�������$�a �Q*a�%�P�!�\��j&r/7�tO����bgb{�����if6�N� N�F|-��d�$,�|m_1������b�����x*՟gK�T�੆³��.��>~T3��/u��\ؓ��/"�=�zV��.0W��a�ё[2�X��z|7qS"&�=�� ,xV���}u4;Úr�d�{�%�'	���泇���{)\?g�������� *i"6�kt�+>�G<����ӻ�C�c8yW[׎VS�LGxs��S��VŮ�@��3b5&Qqk�W/7RUw�z9O��f*^��fS�S.��-'������(�1��m��<(0sH�t9BN���S/�'H �bw.j�ը�N۾\����f�J��T��q͙q�y�4�js�����vW���=�/_ԯve��M�$���ÇV�IfMI�qzS2wA����������cB�+&�W�dW:��pW3VP��Zp��7��}��n�Ѯ�DI�m���]��v�(*E~�7�8{b�;����-ؖ�u�-&���RoB�,��p�fC�F���u��5�9{M`�k��Q�Z=Saׅ�+�%���P�}�0+my����83�q�]Z�=y�颼ý��b`�;ʬӤ�,}I>����T�Q�T0/C��	�<�|t���iz�u��T)Q��3G�X�.`�	��\�uW��"����}0���*�yOh�iZ�
�����}��/yxə\�֊�	ei���[%R��R@�w���	�h�E��;v.�]E�.�BA����/�
7��k�]�y3I��d: 3�[��d���g��J=b�z���7����d��=�T���+Ҟ)������<k~��|cۑ&R�5*`� ���lҰǏVU�yҎ����r�\�mᶕt�s�k�w絲�r�X]'
�$�w[�2��!2�T{v�z�q����Y���_��Ѽ��)t�i�G8w ��_;'ܷ��{�?9�k��Lwpfy�3�v垮���)��/�UU��ɪݰ��b�c6X}���R�����V�8���W�UJ�k���Qe�~d��J�'����G��J���Cr����/mׅ�W�
`��ȼ(�� \�H8��^y�c<�Გ������2b�K!��o�r����F.��ӊ9.�="U�,f���� ��BkaOp�ƥ��h �[����6��бE�Mv�Oz��KV���V��#@kjo��ˤ����ܶe�Tf����D�����Bt�$�0,�8US�,0Ȑl���{`�+�y.�=Zv��ī
�c����V�$�������E^n���It�}L��7�ؓ��u��^2���f] 6�V��ia��R�)��a�4H��|���5v4b'�&H��I���{�*�Z��O�D��r��L�mw���Hj��zs�[T�%�3�#�yZ�	�� �{j��#�^�����fT�H��*���'��� KT�`.ׄ�Z�����G�J�^�}PX��8ߢ��~�F<�A���5i��T熷ٶ�x�v�ل��a��p�ιcV=7�u�E�J?�W�B���kQ7�IrG���}KIn=X��v�ޝ-��C�m�\I��yn-�	3c�6t�jq�d΅����k�Tn�8�MR@6��J�����砬te�%O�@�,5{t�L��MV�c�����˛��Mp���O��U��쑆)��6쀃D��#S�PF��}Gu�Y05��;�5��W�^ʠnE�w�&a{�3���g�F�O0:���!ױ�@8��ݑ���g�ެ�j������Z��Ȩc(ӟC4�Vw(��0�:��Y?w�\�C��~6ycWM��;y=]�GX�|� :
Q���ُ�Z=u�Ƣ�<�|1�&N��8P�ZSKe�1���䪢�#K?oz���U��hz����ӳSqW���AN�TU& �')�ީR�	���!���*Y;�@n?�֤C��`�C^a=L�~G�f;EZ���w�j�\+G2���fQ��F�
�\@�|�}�Lwz�Zjϐ���Fk����ݘ������ye��yn�X�^�	�Fl �DCf��|�I�ʡ�-�н(��ɉ���l��{�~�T���/ -��zU�[�W�4�׆n�Ch�'q���%P�d��,I���j�9�)�9����e��E�Ф
��i:��'�d�HV�������V�Q�ÐZ����zK�Em[�}s���WpCi6��I&e����Y�hZ��ŊZ���f����1��x�%ͳ׏N;�h�P�3<��2�
��W(�gF3�����g�ѱ���})��p"�sM\�3Of���� �*�W)9°�W��M�� �>��˙�(we��j9\՝S�I�gP�[9�g;��в�7ۑ�%�Ux���Y/T���۩� ��'o"�t �/,�7�i��كn-�f*�7{�5��*�[�<���Mf̈́�g���\;x���Nu��S���r�NɟqX�\(w��G��0RE���ͩ�z����e�}�%����($�tx'<�oa�Wt:��F��/n^RÇ��|�bj�&+�����䙭.��] �!����R�.����p.�&��9i����ak���X�Yw�M��0�U��;�N�D������E[��h����4����Y��� ��x5l+6��u�z���ɵ��"�Q��������828��fGV_V%4�:��rj�sL �*r,���w0�{\}��^��Q�PᾺt����%j�n?�8;$����ym��|�e�^כ���P����io�w.�epT����*����� ,X��3�#�]�q�^���K'+���l2C�zC ��v*z-�V�8�~��}=��+�*�1?MEOD�9{�S� �2��5��q��W�\^�d}˙�MD�z��آzf�`G{78�.��4��u�bn��1$���Ē)�YY}�_9�lxؒ��Z5���W ;��=���x(譔�b��v�:-"Wl� �T�0�mi���xN�3�ۋc�6�L��l��1��G���kN�33)n[�6#���T���qdڵ��M4֊|+fx���]�ٹ:�����<��x�<Xp��bo�P������$��6� �K�����&�Yiv�d�I�^ah�}��Oo5�l,�V��y�y�9�sY���L4��}� +F�X�jh��*9D���S4k]p��=��;(̩F!`�~����ٯ���n6�k���rR�a6��r�ˍj�����w0.՗q:�}q�6{���p�"�k�7�ҝ3gRTmT�ȕo��5sѼY��-%�ى�]�ل�>n�K�!����V(�����&f�7p�s��<�lL�BO;ǅ��ղK�u�R�M�wP��S7Z�?�9]�w<c�EJ���Ö-���D��ڵ'ctOr�Uצi��_u	f�؅�q�Q��ݻwV�pw�4�[I�9ޖ�R�l��U�RQM�f���[d@��R�Ρ�kJ��ê�<�{0`�;��nsmh
A��ώW�P
�A��x.w`9ek�����wu�
U͔5h��V�Hn�l�Nk�\���ӵ�۬uC�-:m�"/�E�=�9n=�����\�'��ќz+��6�6&W+u��	�雔�qUḑ�o�<a�tT3ɟ'́�L��5vo�^=w�_l���q�sԼ!U�����
�r"�Nr�Αs��W&\�HLCJ���Ȫ��
�X�fE)P9E#�Z�-#+��8�nNU���TI�*��h���E�R.�bg;5�N�˔QʝB�Qm7t/9IYȠ��D�%Ad,�r�͘�$��T@UgEE��S����Q���i!£̃�)�*,�Z�QEJӕ����
��B�M�p՚Щ+�����9��R�-@����WQ(�+�tȥ����V"��#eR���	$��֜����
��s2�2	2�AY�t��R�\������r͑T�N�Eȸ���q��ZЮI�����!��0�d'Y�r����Q9�R\��a�*!6PDEY�����㿼dU�������1cRTJ�Թ��[]���X����mǯ�36�㇥.����-�S�]��P:���jO������)-d�T&�3f��8�r�����m*��.����\s
MA�iA�ϵؐ��x��,rx�#0,�=^�m�k~f?;��U�<È�U3~\*���;v���|P��%y�i�*�Ε����ą1�����l>�^냅��k��]����!�����^����-͝&.�\.�Ks�^*�+��_�6�K�x��=�}f���\6�\�o}�S]��O��.���De��8�B�Fyث�x'k��y��_�_��5��L'â�"�7֝*��(h�,v�T�����0��Nρ[�5�*}"L�e��׺����ʇE���5����aŭ���	S�u=U�/Cg�xV�,d`ufa���;��xW�@͙�]]�D����QY��"�k�s�޿�U8�n��.cܬ�����Gʝ�(�0W��v*D��o���<������;΢�c�pX�OE8G�0��Z�mԜ���A#%de=쮙~��qV��j
*�WB�߅�GƼ d+̔B	�^��1�P8�&^�?y�����7[�o���$�CAtV��?/Q�xS��=�!��L2�p�p��!�1;��[.#9�@S��C�;�fY"\����lU/��G.��Q��p������<�2�:W^',nLw��ξ�)��A����?����ꛇ���̬��t�F^���%͆i�P� ��ٴ�Q�S��I\м7b�����p!n�&��� �pS�r�Z�=�A=��b�@���?C U�Z}~T.���(� ��;rU�D��S�����0ا�T��a��� Z�;��n*a�d@d�h{o� M~U^���;y�6��n��K�[�{����?{ ^��Պ��q�C>�����
�B�ζl`<�;���X�F�J�Dy-�}�EW�d����d�hՈzׯ����k�]����1�pL�<3��()��0뼺ܧ�^��Ok�S+P
��Ƚ���*��������o�C��:Y��ŧ�x�걪�޻*���AP�|v���^�0/��w:��|X�sۏ��ˡ Il5��Ӂ�+Ǫ-�����%����s�b��9��ƛ������O��ǐ��:����.ס��G�0�a=�qߖ/N�|O>�yf5���i�U<|�N4tvo��Ƌ�V,Y�8��<��-|(�>�w���^��q��}�����
�9��{��CPT�ִ�b)���{�����������i����5ʵK5{����x>uw�7KE�XfI�mڴ�cmƢuf�����>��������X�2�ȽpO[�F�6'r�g{�����ꐶ����d�i�l�n�������b/���}�}Đ�:��/��v`ߗ��|�U8�Y~�ѮއY5���^S�ʮ�B=��Y��F� �d��6h�܆}���\﮷c^�:����l�'��
}|�J�P쭃eIAV�Lh�O=@w����l_?U�~J�'�w�U.�r򯧫ʧ/zj�SC>}�Ґ���ڙ�[*�[�yҤO᜶�i�Kh�mҌ#X©�unZ�ZE�`VXޯL[]㯶�S��C�Ȭ=�Q�'��r�F�Z�o_�h矫}H_z��z�/O2�}�v���?T{C���~��@Y�T��
�J�u7���ZųaCn��Y4��Tml���SY,�
�֬���z>�r9X3O����>�U�)V��_t�z�1{,c��wt���1kr{�����w/�6���#Ӌ���Φk[�מ��`a��w��@z��ݬ*9�剻p�r<��Cs7�ՇR/���0M���,���0�?F.��.M�C���kY�a�[�^җS�$��2�@V+�tHo��"�����n�c�v�6�ZŪ�l_{��7�ᓏ)@�1Yo��xG�v��_?Kuo��3�t�予���v�>*���rOxYW,{�b^�`_kΪK�3��d�=�;B�h��)��u�X���s$��t)�s��{�e������k)I��Qm�Z�,����Lb3�JI*��NY%V�s6��*��'I᫩�E.���bT+��u� (+7��ս��Y��Z�c��)�{���v��;'�њ�-����e�'��V�OB��r�XE��ץhQ�az�jlt�E��^H[j�N�}Ƃjq
�4�����cS��:�����E��s��m����K��;ς�]^;I��T%Nt
ه����3�e��	%���I]SV�8.�d�K����FOYW�*�z�Ƒ�R�b�݃�r�ܓL^�0������EG�zR6`�Z`��M?2��U��bB��so��Zi�ݣ]j�p[`T�"f'"W�l�����.���9��#pdĕ@A�����63뤹��*��.ٟ�M�;X����b�F0��G6���d���r5���1�"=A;�ʳ�j��u��3(Qw�\�I��������o�B�2u���W�٫X����:�͖����{�Td4k�ޮlzU�a�vK�Փl�wL�����|QūԽ���N�����ʹ�)�Ԩ�iiT� +p�/�LL��6Ҳ�C�W�s��zuyulym>�S�7T�3�0�I�R�p先�L��m�Km_V�Ը�F���};X��<&�[��A^���yWv�'��������y	����Οs9Vw��}ޠ�C<����ci2�uH,�mԎe�Z�>�����ѝ���]���l�<�s�)ޭ��{r禿����f:�R?��M��{�B�g޹'�3H���Ӫ��9���|�n�l�4�)w�����7��®��|�R�X�^��#91m���2��h�%o��F�M/l�O�豒��&�gm��kA����)��l�I_{)��g�����m���[�*Tn��S�+���r�;,Pͥ����w����g�J��Fm���q�ݍ��qP��:��!�ьy�z^,湌���.1�g'e�6�J/z�e�����2��j��i��i�\i��9�m�WrV����y����s7en])��̖��J��.+������k*��{�Wnlj�!���)iֹ�{��3Q��	K<l"�㍨yl�������KW.�X���/�c�ay�ی#kX�Ĭl3��L3�zmX�r��:�$-�Y�NM{�W�^�9 �ROY��S�&��}�0ˍ�'ߏ�z��}���W5a��XV��R@�V���Q�:�H�I���U����DG��{iN��*��Ȅ_�j����U3�*���p��b�~Ԟ[�j�h�Sۏ�w���F=����Ji�f2���o��Y�ϰX	DR��z����M2�mŘf����[R�q�Cl)��Κ]�v	SЧ�4&ibpГ#x�)Ъ�=��욽�A7�:�Qs�XӼ���W�B��YxǼ}��BM~ܞ�gw�������C^u����V襴-1��}�7��.�WT\�z��&�{XBL=���=&�&�9�u��zPkc�@ݭo�}"�{���4�M�2��AκnV,B��r<�FW<��U�#��u�j�U�./P9�Vǵ�.NR���1Q�V���U��T����V�"�0,���[�&��W��U}Uy]���(��3Z�������Ւo�n:>�;	�a�S��s���b��ut�z�`���t�&��nI�����C��ڥ=�OV�w�jP�[Ó�����vC|D�*M��\�՞�o��7��E���b�vj�5���8�/Sk�Kwg©#����e0m-ݧ4��L���hè�w��W&�ݷ4Θ��N����=�\����)}.]���`�����;��O���z���8�~8�쨲G��0wjL�H��Z�Sjgh�蹅X%X�r3������BݢdԪ�l�8���|M�&L���v���*FL����]�Yua3��~4�H�e.�W�/��-��2�q{�w�O�v�i>]1���%�תA0ͬ�����x��U[@�#n��e? =Li���<��ꚬ�('@}^����&�
�ɍɇ��G�5��F+"��푻h���k:�,Ɛ�vIʁ��[��l:��ʵ�u|j����åav�����z_Tv�Ocj��S��`����`����CW�������l�&06�N`�!�s��%m��w�\YB�
�c�w/u^�%���m�mʊ�^����f{[OH+JL�w�Ӕ�[Nʧ^*�e�.��V��cs1���g���a�,�[�O�1��M;խOz؝n��Y4�J��-�vN2���ѝ�u�a�W�9za���x]�牵�ELV�f��cb��yU��Im3��c��	���d����k!=��~#Ӌ��������d��(�x��<�h�ug�^��r��!p�U��rs�:x����aw,����i��������b6,P�Ek��I��ceK=�?�l��Gg��t/�f�s����\���==.��W�z\���2^��=+��s����%�;L�7�K���>����ױw�zo��_�~q���K$xk��,���['�}=�/��n�^���ga(Eʽ<�������W��6�m���Ӣ���b���.�|�*����a�ڕ����<7d�Mz��f��W@���,�����ys���.�����<W&�}BRg�"+~�H;J���K��ʴ�� H�wŜLw�[Rcv�>��ý@M]n���6�ykp��(u۩ۥ2U�zt���o �I�Ok���6�{�oy��c�����1��ѐҨ���7�pZr�۞ݺ�-Wx{{s+m輍�rc�z��]����}]<'Wm}�]��%{����{IAr�:|�5Ε����m���&p^��/F�),��	��Y~��c�lԢXd�[*�㘑r�bO�ڛ���u�r�:�X��*���u�e�] !�i8�^}�]:����w��ߓ������m(�[0�H7I�+A�kP��g*6n׷�R6�5w�G����S^>��>~گ?'�� �=2�$'�OO.�M�et�b_{���������E��<�c��)��V�Egl���׍�}�V�6����G��~Σ��7����;���kgK5J��vC�^ɱ�wibݸjJ߽�[F	��9]��]��{�Q�OP�r��ӏТ }��~���J�=��lX_���c�s?d5�{�U�~��#�Rθ�#�ɓ��ME��&�V�oNa�Vf����K]�nR�f�mj�Ǵ�~Y�:�N�"r�|��9Ѡn�u?�s:�7�Pu~x��XS��h�$eʁ���x��m���*%w���!�6R�k�ld2��W�UUUx�zؕS�pi��~���7�{��Yrۨ_#�J�w�j��^%�:ߞ��}�r��Oӳ��IG{*�o~Q�<�g���8�/a�}At�+�������f�+��mĚ��6��ož�6�y�eyh&�>�?�ŽY{� ?Kx]Es(W��(l�H���]����Byn�=�l ;�͚7} �w<7��=Q߬/��eO_�U��g����}�������j)l���be��S�Zc�bP£Pg+YkU~zá*�b4�RۅC\�>��6�KU�E[��z���ޯ:Ҫ�o��3�޵)��hi�|�is�q̷ʴΪ��٭�gVc�|!>�b�JP7C;�D���U2��,/�=�ƽ��{�jy����V�k�J0�m�U�\!����tR߻�w\��1L�Ʞu:2�_���)b��ci�A�>��u�4�����;�sZ9`��m]
%f;��N�=���v7Q�T�1��7��&wݽ�S�9W,)km�J�����Q�]�r��h�3�2�|���i��v�{ز���o��1�X��o�8[����֥��'Wmުg��bgv:˃7/��-O���J& ��|��Y�{�=�0�`	r{ds�BnذoH���3�e�(l!14��ӛzS[�5V8��`��(����,��Te֪�!����FeD4�{��}����L��}p�������ɠ��=�X<��7�
�$���n!���� ������e��5WT�ӷ7e�+�a܈�o)��Ϫ�)��+���8Er,��D���m`�."��Z�0����[�@,����e	�m�K��w�ё;������陼���t��8,���=ڝ�o}9Lx^o����V�b�ٷ<�+���$�j[6��)uZ�j�W(��z���~����Ȳ��ֱ9��+p�+�Vw�sCP�Bwz��"\f����w���W8;���۸�Ӓ乀*k5Qɱ���]�/M<��ɇ.L�E������N�����jX��qH�5���0���G��/ie�T�y|o>�"n2mvu��;bKs�զ��n\��V`�El�V�^db�^������g^U����|����h�K�M�|4��ڧvl򤁼*���|�V�py`�V�"�;6m��[��������o��r�Vw`f�+,�z���2N6�Hi�u�3�����,3@h��]*�'���кs��+��:�&'���Bsa��ȣ��U��U�~�k����g_ T���
o1`G.��~I��^��}.N�~����x*��k�)J����YE�"0X���R�)���.Q�0\�����J��=le��_^��^-,��lt�����څG���zy	iJjc������ej�ܭ����f�����K�{X3��K���j��ʇ{ri��3���9
�m�M9t_�C\��&N� D���,��ݻ���D�x�m:�]�Ǉ4�}�If�ȶ~�v_a���鋅�jRkWVj�ku�^�yv�knp�6H3a��-�[���B)	�8�Qҹ{e��������^���+7��ܝ5�(Sη��f<�\�g�ױ2���7�q���逸bA��J��|��a�m�2��u\E���b�:�r��S���O��j�g��g>8X5ۀ� ���̄fNi��z�V�R�(�P|T�a�;v�kk���X��L�����X�f�d��cӠ�ͅ��W���r�)� �A���^��ۈ�]ٴ�<��{����q
���/D)3�2��U\�J��s�KK��8PG(.J��ÕUT�(�Ȥ����Qr��EEEr�\�1N DQGE#��L�R�AeDN�fE�Ȫ�
Ց�U=�� ��'@��N�W*�dy%Q	й�!0�T�TY�r*��AE�p3b�����$*���Ȼ�G*���TPEU��/wn��Er��#0��9Ȫ�B�*���s��p��D�sR�wp"(s�x�3:t�h�d\�e˔r�<���0�TT�	�[
��EUPTr�"g/0�G�S(�2�wbr�8r���,�*�V���T!AFHE��4�Q�+����RwU��s�Q9!d��*�Gt �H��9Q9ȫ�ܱ
���h�r��.�ʠ��i�"�V���R�p�DAjr.!�9Qʫ��]�tBa�(�ZL겊���$�Eݹ3�w}AƽJ�/G����oP��8 Apg:�\'�`z:*�9�̔�l�#��Z8�A��)񌆁��]^������R�T��OV=�o�{����=5��UQ[T#�}����Z�go��.oT�<������N�/b��g����qy��=�V�����s�s�����ys|�>iJ��}��u.�[O�j�t.��O{&�{�s�`���髣L��$�
���o+���߈]�G���cZ��R�רե�)�QYS:z�S�P����~���O:ϟ�ӷ�ٝ�{ݿ>����w7�Nܽ��t�gy�~��6�`��W��m�K���t�����G}�:Es������̹~bI�n��Z�E+'r�f�Z����^�C����	>�P�yw:���]�t�$�uim��b�УN��q�P݆�ٷ.���x�n���ŀo��^�w�ϩ:��*m��Hx�8Y�P[7lV�%rW�h��.ټK���5�_q'����Ad��;�6��7���N:�8��P�绯KW����J��n�ۼu{u)ε��-���wM�o�G��36���D����TEnVg;Õ���]�\�w��n@�Q�}u�!�}�KX���82�,���Ҏ�Z`���n�'{�!3$T�Չ��w��d���Ց"�Ҳ�����T��7���dZd������;4N�x���	j��"��>���E=K`�0�b�V^�X�,���tl�tvml��/JʚSsޭ��j��ƻa��..��3%�&��S-^8�����J�YW���V�7�ê]���<�%��yn{-��6S(s��$5[0�S72K��h?�H�����Wپ�O>fC+b�v��ұ��<y*���&�Jh��;&�n�������W+�/�^9Q�MJ�5>k�	��Ħ��[�HI��S�������� ��z�Wǵ���u.ߘ��}Bt�߻|���3���،2a�N�'�0�I��j�*�d�:c�{����|��ӧ�&�-�����?T_�G}�U&l�U�b�3��8�gs��GO{��籞���g+(̽�������6�x(��Smu���ƶ��ӑȶ�|���u,��*����Hs�᫹i�Ztj�Fsb���.�OrLq<��	��I��%��k�"Y�W����,�4q�����mM��@u��C�3s��CG^��P^�ل����c3^���k��"����:N�ά�Ÿ��i��H��"�bVgk����������qw�<�j�Q�׹�z����yI��݆V��cmC>>;
͢sv�N��T��8̯G�7'<rw��M��h�����C����˞y��sձ']����/\ȕ�<Ӷ����5���[�*����~��̎v2�u�*�f���������N�Ey�nUSN�v�ƟP������eV`����~��R�r7�reA~��s�++O!�{͛�=~�n�ɷ��x�l����-���*�j�V�^�c!�=(�/g5M_�2�j��(����	{^���]���A�JF�lH��Y~������iɨ�y��e\N��NV�����[O���d�x����O_��3�eo��!S��ݦO5�j���c�t����֭E'��K�}�����8ѹT�B� ����q������-]KϩUL��~>�S���=��E�oަ��&6��9M����Ɗ0��E��S��z����6Ng�ɓ�$�%��N����Q��d����/r�u�	-%���}�3��J���<wdӼ�#�:�K.=�$�'e�sO磌���s3}J�x�4s�ː;�r���*�:�Q��E�����O����]{�g�؄ܴ>���SNyQ���c�vMD/i�NĠ��>�Q�m��"j<��k�w���
�)ۥ&�U���і�Y�;�G�� Zt��&�eA鮰�u[�}�:N�(�n�k��ʄbus�*Y��]��C�\n��u4�^��[�'��r?�u���5�������ϗ^����g?)o7S״���W1���;<t�{>-k�צ���:>D_J��yo����R�1�K�V��������9���s�ݍ���pwBY'[_�ڳ����������VN�5�mb���s��y=`оlw�º���+o���]0o�z���Yp�g:����Q�n�;F^4 T�-2-��H�:-d��U��w_��ɿ_{����y�8�huN�}�NJv�#� n?i�.��=׏�^��gV�l��W(�s�}��/*�9ٺ}���8(��Z\�����ݝj�cP���ק�t�f��N�O^�h��"se'�Yݰe����dU���y�[s��Z�[�X�$���ѻ%��Iq�'[Z��fn�苘jk;E� ��G��4�Q���7�����������[s���5٭6JlR���jP�O���K��^�'����d�U�<���J��Մl�a	�0O��H��Z1�Tc�AVR(�c�TG�[v��RbT�VڰkZY�Ҍ#Z5U����t��qF�������܎�!7����~6[�UT�Z��^�([�J�%�f
�ԅ�h��%s�Դ(jSF*�[B�|SMC�1�Q{>�����j�Ӑ�)�.)�=�V��X�6��{+f��Ԩe���6{�yjP�08}��ܗkԆi�C�u��E�Q�M��N��fJ�%e�*��S�B;�Z.^$�$'��x]�g�eQ�#H^7�Ҙ��~��}3��l���d���:�c��o���\�C�9.��{�e[����ֹƮM��d����c�<��R�|^o�϶���*a�]��t���%�4<��f��Y{Gm��N����xF��N�Vp��;=�(��m�i�p�kx�C�S^}��U��v��d﷕��ћR��Bu��W���f���M�V��h�S@�YS��ScKY\�[����s�B���/e���v��DK���{��7�y9��(OFr���J�nE&�;��[v�W/�0�;�r�ׅzn�^��eh�ޤ��+�l�Z�M�ihԎ�
�E�n_؂��U�n�3����y�^��.z���i'h��4����[*6��bin�ԼC�o����yi�Ш[1LL��Z�r�ǵiM���6��駻O�t��$��\+�{��l��k4�sٚ%�B*�.c�ޏD�]OmcQ＼������n�(���@�Kپ��*�/f�,�M�f��^����C~�K�Je���J��?�@%k,�b�Z�kf�[�c��Ӭ�ɂ�#
�.�����ҀM��Ԟ�l=��bl�b�T��l�;�`��c9O��^�.qm�0֛��zM,��juM�e��I�	�gj�n���甓&�r�z-�%4o���}ykJ�z՚��P�7U쬚xjTo�mlB#'D&(Y��i9�d�^�,v`�����Jglp����}�����B�uέ�z������{׻�`ۧ�Q��gWlt��*�r�����x�dW�������E��%���g}5T�󝵖�������t�Ml�BpZ9q׻"]ޡoi�g{:�������3y�f+6R�F�M�h��|iz>��:]K��<���Ξ���,�Q���}�!����;��׀�^����BF}0q�<��˪��՟t��5�[�^r�͡$�_��\�2W�v�kS��T�Q�r^�NK6:o�g{^ޔ�J�=mf���a��^[k�ƧSi�e3�^�C��䕕���s������3�o	��V�s׹�z��̯n<�R��d�RW��'w�\S�E˭ɯ'zf��f��i�M��l��UOy}m��wG�R�$�J��au	V2�̴�46�^�LY�΄՞�h��Jm�}�sOW�s�C�z�����صý+������u��V�Ț��w�ͿZ������8��Ieҙj�	$�KQ��iE�ؠ�_§���j�w0��\��k��tZ�դzgnuL��:-2�P5�G�&���Җ���z�΁[3>��>����_.��c�,{�{�:FI��&h	��w]��ڋy�j�d���]MT5կ���黜���O�a�ݡAt�G����9��5՘V����p`j�6���~X%�{�6_b~���5�V_Iq�{�uĽw��7��#U(Z����1��S�4M�[�)a�Ϻ���6��Z��,y]I�==���&�����ᔹXϒN���!?��	=&�{P	����(fLdb����6�K
�-^����c�t�!�Zu(�ʌm��ך��D�u=��x���hwW;~�G�qj�^��&u?o��kf�˛^�3'�8�������+n�Zc��'��ua�<��I�T�g�0��H&:�>�ʌ1�[i<?'oj�+��%p�u=�o�/mjk��Q���5L\�T��eK��L��C2Q�:p��/�]0�T�^u��C��~��c:�����>��^�+�/g���:1ݿ>��~�����y:�t5�Y�Q)[��ua��|��X}�g�f�h��GO]k���v_�ݎzk�sνpS� V��;�u.��Q��%M�\���N�x��w�mҏ�ރ����Q�9��g`~��`5�.� uƇ)�v�T�ˌ�:��Z ��l�~��ϤvH+�o,O�.O���L$f89�!��o ���/+Wooc��L��x1Vm)��Wo��t��`L��zy8S�w!�q𮂎�ȥ�sJ�UUUTI�vz���@?�R�uЗ��	��K��rϸnV�U�{���Ib���C)���7�屑ua�S릠�(�m�==G�:�5g�\Ω�wύ_��)�ɇ �tF���w���Ҥ3��g� �P�r��3��{��e��:�ܡ�̨��˻YuW=��T~�*?u��Gsl�t��%�\l��e�������2��+�/�q�փ�lC$6�M�Y��/d]�����)V*�����ɀ��{9	K���Q��Ӧq��׌[b��IWs��[Z���8�$ݷ,^�嚞iKT�ڰn��[�v4����E�4g*�i
d���O[S֤x>��y��5Ib��c	������Nec�%y�gY2zeJq�֩G�mU�S�KF]x���1�Q{�&/.5�XJC���׾���%\�վ��U�t~.Ol���Vm/ ���m�J��y*w�t�V0g�1}��(��\��0F!^0�[5m��M��5*J�34�����^���k���=�C��B�9�M-��>%n#�v�7��2:��m�m٩�z6���7{&�߳W²oZ����.�=)�i,f����o{!�:Z��� �̔Q��YI�a���Zc��Nj��[�V��N������}Y�ޠ�'%��Q�n�.��&����=��j��9[���!��G5KY<�g�q�o�ùͥ���.�T�.���'{�ɱ?_)^&]�����6uL{��K�.{�w�O�^&�\���++_��F'w��P�(E������R6o-2շ�+X��+a�we���x-erϘt>5�6`�z{���o����H�ݪ�w��U�v�t�Q���(bOryh"�ީ��{�Dc��r'�>�»ٯc�����k�+��~��Z��bQՋ�S��
�N'.S.�К�BU2L��f�j>CZF�ˆQUR�Y\X5j-��TX�W\��(�VN��y��U2�)�$�]��
�+Ϛ|�V�W4V��Pϊ�c����3��-Se�i;���Y�x�ZW(�C��Oe�;I�X�L��kn;�
3x!Q�-"�i�F.�S�e1f��[ڪ�j��]�rr��&J��˕yF���j���ZP�4v��Sw�KAO�]��wQT��2[׿s��Z�W 'dX�������5+�'m�}��*3��P>H�ذ;�;{f��{����*W��Nv�"o�n���G��3�ݎ!�2��g��qk�u�D��y�"b�uSY��JqR�`Ӻ�v��Y�Q�u��n�3��Y\�S����Eͳr$�Y�9�a���Ө	����ofQ�4>n*����e3���q�E�W�ѳ"x��O����ʓ������:ؘ�p��[��[�"y�TQh���
55N6z���ن���:ES�����<TUMZ�q�k���!��3W-�z>��AF_T'F�1!*�s�4{=fg����Opv��K���,1c2>	9P9V1�L�v�lƝ���1Z�`#-7�f�������r�`G*�쭡euNل��}NDV�b�tq񴤂�rT�zN9y.U� �{W��#��FR&3�oY/�[�'[�+4&�=\>ҽ�|���b�
�kU��c���v�er�Q��A��Ƀ�Q����3�N?;�$M�{sQN;
��,P��>w]� /�3rsY&����͖>�'7��R�j�VH��F���5�a���Yz-�`�S��J;��ځ�X���Sؘ�:�|�� t����8��z�KF��I��O���#��O�x`;����;��<}T*L1-�p�K�G:]1�ڽ�:��ܧ�k�LT�ڎ�GFv��1����Gl:%�![$���շ��g�%��:�x�,�Z^�r�/9����i�I8򫫻�XJ���
J�J�ݛ���<��f�w(�h��kV���ig���ƬFr��ٹܝv���ź��������q�����
6���_�ϊ���pJ���s�m2�3D]���K�tM�%�9���0�u�-��¹qe�<� �2M��$�ڴM3�T�'���/c�y��o�+4�E@�O|m��2���ձ��i\c���r��:��e&��/f������r"��oJ�R:���u��p]�)��յ�ja���=U�h�/���N��)���
���W�=+��\8,�#��8�8��|�X��OZNgF����枅���:y��21C�ii����|�j��#�6[$�����1�}-�N���,-�O�M#^�S��7r�鑞��_��O9��j��}�mc��Dx���7z�_h���+v5�Fg8���ު�Kx�<Nҙ2ɽm��)���uo����|gJ�o�b�d�2Q�Z5��tIr�� `��^�g�v��m�)(Ԝ��5��]��{ww6!�wT���b>��/-�j�J�t��`��I���4��)�q�No���K�m=�MV�����U��>��`s�od������p���N�6-�#E�������޿�w�Ƿ��D�U�DUI%�J(�$*�C�0�.QҡE%$�.�GH֜��0�e�X9\�s���$�T��D+��	T'"��\U�E´�-�������%R�8Ur(���9.��w2��r8�Ep��¹UG5i�e
�,��)��ÑT�p�$���Tr����Qs���p�U$r� �^� �zܜ�Q*Qe���슋ZY�3�UD\�8UET�G+��AY���E�DA�.ETQ�sR�\�˘�U�4�(H���U�ą�seW9p��֗I�BHgBT��G*j�˦AE�z�@��(*�Q*��uK���j�E©�A
��ʹUL�����R�����8�(�ɕr8��$뛎�¨��)	.�D��UM��
�`UP�*֓*�LB9QUʪ�p����?�;���yD��� ���
��&�!�N�j��(����=�_n���c<eloFמE�&n�12��(+]-��G{��������&�H����S��|JQ�l�.�W�l��W���׾�4�g��%���YyAK1���&��EC2OJXl�Z�K�&�
��̡*�_r[*�/pZ:\S�R���0�z���`�՗�C+ڸR��t��^a���Od.>�I{��ɘ��2�R���YQ�e{}Y�w������4�פ�JN����P���QP�Q�=�iں�;�T��N��L�I��>桋��_���}����W9�P�W՞��������7iP�0��;��&]qC@�z>'��f�jr]M�r�^�r2�Oz>�B�Z
���zq�!��W���U�gn9=���yT�<tgT�]t�Os���W�f�p�M��#��v�>�w�uy��up���*w�5/-�z��;�o���������.V::ʷ<]\�����w<��~ъ���}����.�|/0B��,@�(���`wˏ)�.{f�����e���Ӷ�
�̺X����hT���p`J�Z2���2|0֚�gVi���M�ԧjZ�2o�����Ǝl�wM��ln�IGg�[��x�D�λr�:����_����q��w����r�+��<�yĚ��mxJis������P�=&���saK=P�C1�`�7�?{.�oD�������D�q�n^��Lq��3�z��XRו>Bs�8/�)��vD9hTF�I]�7�9���bX-�֮bs��g̡�mRc-`gh�(�ӘQ�fX���s\��dOfq���Sb�8�H�g�	�>���TR�-ZN��I,�wm2y�5(��3�2#q�Y;�|��y�'��o���[3���A[W�/G~K �/!q�����%��qm.�+��F�{����>�F[��R>�l����0��4v��l4GTW���a~(��Խ��}3�n�+<��p�I2C��
�槪��1K�]�uȨ"�Σ�k�E���]��n5mx*[KU���6D����'Ӻ�ul�+�q�C.J��k:����V���~���Oɒ��%R�;��.�$�[}Fʆ./6W\i���Ɍ񓏯{Q�K7|��e_��J(�R���;T���j�D��x��x�sn�6ɫ{��=A��G�_P��`�.�"�B�hd[�:E��f��x�}����'j�U)�ٯ[<�Z�YUi�ٹ�6)�U�IU���Z�����l-ܝx�j�T,�p��y�mQ�4�v���ztk�{�!O�'B�^�����\��߼=P:lL�A�{}ƶ���;��S�w�ތ���<��%�j���o�R?^a��ݕ�j>�]����˙�t���������h	���#ɓr���/��޿�_���	��K��wA�/�N��[Y���[g6S܅��JxQ�QO�֢si����:4rn);�m/>-��#)^���4磡���G�_�)j*}�����&�����W��8N� o��7,3j�b�[���Ǎ�m�Pϴ�-�ޑ���8�Gs��>���5X�f�c)��5|r�����2��{hOW�@�)��(��������.�[2�EM)H����]�/�ߦn?O�e�!b�b�]o�7���n��@�i5H���Y���"|��Y����M�tzi>ߛq\Ѩ����H�j��i̫gx�Z����mF�c{��\j�݆:�y5�p���H>D�xvA|�A��F�5���pb�͖w37��V�u%I�[�X����ƚ�ݷ>/}r�O4���-X5���H�7	�C�����n��� �mNG�iC$��f���������E� �����3l����E홑&
V��G�e43VhQJh���;��[Dz���=E)�d��s�谈�[;Zԭ4��cV�0͚�NF�R���[|_�m�>��R�T􁔽ӭ�_z�:�|{X�!{iuNw���N�Z��~����F��zX�
��[�U�=\���J����h�.7�Ҙ�~�Q{�^�;HZ'�[ө��Z�:�u����~�\�\��u�~�N��vgz��x)��=��6�˿8����e�����W33}��uBJ�t��=�O�}�:�2G�����WUM�w�fj��V.>���p�����)ۈdԳ-@��U��1�^�������c>�u�}=����.���ƭ_q��q&x �@5�Ix5��8���4&�ҘՋ�ƝOK�Q[!����SY�fRٝL��n�;�PG˭�	�%�-�9�ԩÌ�!|�ۼ]kagt'V����6�l�#v�7�jBu��#�WU�r���y���W[7+��W��#�_�D]H�Ug�o�l�Xiw������p�{�?+;E���䫎e��4�Ǩ�|3lUy	LPY3#fա'1�j��絧ʇ���{�kf�#[�X_KQS=^���y�e}��ͣ�l����z-�?bkr�m��5����)2���b쭋f�.�����gUjjl��i>���-z�]%�-��Ϣ�핱��%����ꛎ�q՗}/�Y��a�����S'^��nh/��dB��5�i�=*��Z};����L��7��I�;��o�3Ԏ-]�5�A�K�S��{�N/ygf[�7p��M�@l��Q�&=*-MK�z��E�S�5�6(M���'m@M�Y����暁RSV�X����g���6Ϛ�]�ymWV��A������Gý��i�=U�K��&}������7z���tG�e��X&���h�+���;B�`�'2�\��dj�+�њ���<n��v踼�T���{}�SC_t��-��-�9�Bb�i8����K��5�C��u�)��'Q�v+���he$����.�P�n)�/`�r�~����I�}�=��_���{|!u:/�n�K=�6�c������0��(�}�{0'����\���.�ɱe�gnS������o�
	*f/�D���.����%Lb�J��sh����I���z���m�7s�l��l��r^VYx��CZ�x,eg�ƴ�xoǺm$���yzv�αF9}����[6��^��;���+f<�-yĚ��oR�5W�Cw�ܫ]7�b�G2M��!�__%�Z�mZ��޷��̩����]\�%��i��ՙGq1[!kSb���N�F�C����47T[2���;�_��n�\-П)�&�16ZR��0���,��0�//Z���QEM���[���'���`���6YٱBs�`��D���%�z�oR���E�-���U/+.�Z��g�B4�`��'���*Z�=���J��{�hҫ��Ts�3��`�7��?e�p�	zޗ	O�UI�&��sP�'�?��E�5/��X�����܆U�:s+��*l�!�v�4ཨ�6��}�p=�^��ݵ#�2�;�@�X�zA��oV6�lt7F���B�o7�"�j�TN�����v�?3K
�H��ޱ����{i�]K�L8����0��~�,.��}��̳�Ϸ�x�}��}��ΫeD���n���z�Wy���^�^����~�+l�=EC�gQϏ������^-�F��.>���3�F��?�v�ժ���)��6�e\5�D�X�b���	�G:��ཿQ�;~c������s��<���o�γ��3F)f�c{�<g;��{<k(��g�c���lk���I�zz���Lc�u&���<;���s�%��usܒ���];}Y��Z�{:�Ov���;*k�c�X߽�^���}P���J��us90�����{������ku��g*�+Ibʬd�C��=�[-"}Gf݇8�֣dB��Uǻ�d�x�3�qx���c!��v�(�ڑ����u��v*�Y-��Hw�ug�Q��6��ƓSu��ϟU�^��y����X�au�����W7]{�uk���A��'ؚ3�
��y�Q�� ������
pͶh��;V���|ʊ����N��|p��,�����3Qu��l��{�!T�-�0�C��0�UU�`���襶�P�m�L��Li���-�{s*[K\�]̺[U�6���yЧ��3,5UHٴ{)�<5i���(jGD!�#4�� [���ڵJZ+K#l�>��G��Ul�m�%��������WO�/{N<�6�fQU<-�ޖ�uN@��}y��Ҳ`+'���]a�����]�]�[��B�$�����?�Lrn�hc�������ڙ~�O<Vz������ѝe�z�eq�͈'d�^�ũ��/TѾzov5gD�IgT%ﷵ�/`Ǉt�Y�j��{R�+4(�)�	T�-�h��L��j�����
����g�y���3W��z���;<��ϗ�>a��_��	�L�����g�<�𕪏��!{WT�c�~~�S��;˵ԟ�ʹ�)۽q��1N��:���j�O�K*�,�9�t����|�eu&�n�j*�u�yd�R�.̰���w��먭,�ފg)@vS��=��9�� ��=�]'Z�u�����]c�Й��M��'����9�)D��:sAv_��ݝ7���终(���˧y�B�g0�Q�3���I1U��KY�Ͼ��ݾ���(<'�;_~�i�W���8��CY���mQ���<��W��	:/Y����k�W���w=�a�~�G3�W��T��u��캻�E�����z���tf��l�+ۉCL-���՗,�S�(^�fK�H�zW�O�����T���Y����vA��5&;|ܾ^���糅�(�]�Y>����0ŏ��4�羆�b��x�އ{���h/uy[�M:���4"���u׫K���jվg��y~��k���\y��]:�;�a�����z��8ו3�#}�ţ���{vİ�J�e�cvOd���y:)Q���6�e6'N���c{'�z|��`��.�2}���?>��nc�2ʤ�+��
����ۓ,��\�3|��0�޼��ǝ�^>`���x������D(�5�iI�6�թ�h�"��e����z\��y�4����:�f)�mmJ��6�����g��m׫�)`�\��2}�$�C�K�˓������ �hx�rL���%Ǝ@2��`nȳ��ݻ��]��e�8�0P}�cy�L��5�o�n���O�}�}>O=���H�������qj����*g��>�O�����X(��9�d������.�3�s�њ.���A=G�Q����7Ơ7%��fM�z{��������V��z����N���Zwl�ʀӱ-�S�L��0"Ћd͓C���-��[�2j�����<��F��U�Wo8����#�9��������ӊ�]]s�J3/�����p/]�I� ��H���mt�^��}�{h��/{��n>�Vοy�V��W<Y�
�딅k�L��t9%���:��P���n�z�l^�^��W��$�C��;�*�g�G	e�;���
��}���ÿƴ�xm饞��7�\��4�1[��[�wɕ��8�1JAS���uݟ�缰,��	��i�jP��>�����ukV�e� �<���:�a�T��Qu�GCM�X1?{.�vb�����,�ў���b��f�L	�cr��4�8�J�i0kf�m0��f��Mmk���gI���[A�睞�������:�ݝy�aaC�]�7�t��]�U��D5�15b�w�qv+�ޮ�GLFrt����/n!,��ܔ�Ƞ�w"��݁�oZ�*m�U�"D���c�a��K+�;p9-�a'��$�g+7~::Wkr.}An�*���׻�9�ҕ`?z�۽�u���i�#�g,=)�DX"=��Ryb���ꇝͥ�m�
�ͭ��y�)C/8Swv������F>�b��N
�����"����xV)s�����Ѹ�Z���tҞ�yvX/g%���$ܑԙ���2��"�s��t��{����L�]��٠�87�c��� h�S�ܮNհ���Ǭ�n�s"�j�9�.�WZ6g&�Z9�M��F�e����;oT儆)�o�}|u�n��x����{]���H�����j�J܋���U���V6`�A�yn{������5����9�cك����[�99�ζ4��yoE����q���v�!S��X��ʶa��X*�AX��ڠ�b,(�ϵ��y��oSy�e�[o�ب^��
u<u��ř<ߕ�]��$��Ve���Bç\��S��km�e�k�'����ny�/��9.�����=,�Ϣ�Buckd��ԁ������A)pTgw,fgV��|��w[�Gudj�ג���2M<����λ�;�R89"y.=c&�)���r�:e��9I%l�d������u�ھM�ݾE��0��������ԺbKpU�uc�����Ǻ�-`\j.ɯ�tGn��@I�V��bWf�D�Ѻ���{D�u��O��6�n4Li�Ӆ����Η�mo){��\���a�ӄd�4aם|(ӳ&���RwSr�{k�d��hn������1��I8��"���5�[�ӊ!�--���oZ��SI�er\nf�����l�/I����[�׏@��̰��K��V����m�)
��I>�j#�¤{m�y��.���Yt��*u�Y
��A*|cr%��0E"À�n��{�滄	C]�"�\-��$^p��7����C([��k�8rOi~��h<��i:��nq����"�1r�WT�W�8){/�,%E�X��/",�8���fm={Wv�zw�6*����� �s��W!n�61P��{���j��xhWvT�Tu�j�ZFF��䳰��ʡ�bm=�gmn��*��0����?�VAk�~�-О��h ���q]Vԩh��:�uT�1v\L�Y�k&L�o}�%h�}ܚ�:����P�9��#���t��d��+"qM�����R:��b��Cb�d�Q������xP�Ӷw�(9�>X~P�
�UD��N�\L*NQdDDz'
�ɉ2����*��fQE"��
�U��@#��U2��F�I�����L�\������r�W��DQˑkY��E*'�QBAgC��DQg�]P��\�"�]�"(¶�5.�Rn����T��.�dA� ��Q(,�B�*��.DP����rIR�aȺ�r�r �r �
.�9DT\.\I#�\*�QENI2��r�\�
i�Bqɷu��F�L��\��"9r��%H*�TUy$S**(��Q�� ��"#��2�����A֜�UA91�;�E��.ˑ#�29We�r"�E�9�)���߿1����Ϫu���[��]�t��}�[�4t��X�u�ŝ��(��3q,�
�Q��M�q�g�_}_Oi�]�OT�Y��A����6�m�R�Qg�l�kU"����jj�[ṴȄەj�P�3���.؂v�|�	�G�&�e�-�S��{��x,s�����%˰��ԝ���J���c�|A�Sb�bR�l����Z�U!L����)��ٺ�y.��VLd���#ʮz�����S�2��1t����y��%k^��J�~�hc�CO��Xʥ�Ǽ}4�ɪ�C&�K..�i�+ӰԶ-�Cږ4=QmP��4���V-�Խ]��|�'zI����wn,�Ok��l�==*���*2�EձM5�Z)�E�a[Z�jw9��Hr�Q��zR�����N����������%q��!�O	�t2��
��#HOO�v���UEӁ����S�q�W#9�['��Iv�X�N�X��.����|{��'i�,w>�Sӣ\{Ֆo ���RI�'G�]��/���ͤ��Q^˷�؋��uE+D��_����8Do��Ց�6��V��@V���}�F�i{݋�m�8%��zTz+��Ni���^qgE<��P�\�����H-wX�6�薭pٍ^؉���y��j�X(��~�n�s�J:3�m��O�����̞�'|�D���S�-�~�s�a��ivo�^�O{Ϋ��/��zTۥ���O�}��N�u�0eD��odx��Jɳf��y��C��V	;T�^X66�C��m���S�=@YxF\[�L�(����w�P�Д(U(�P$-�7oo�=�Yuq�t�wT��6ױ�e�)����-��[�����j*���{0u�(������\<�-\�Ч�Tf|�����*�pχw��'�;:���xEKg;FP��EJ�Qg���'v
�ٞ��!�⪤�s�DbY0���\6��;�������J�ڱ����~(��X_.�nm�F�k�<�ֿ��=[ހK���"�t���
P5SG�c��۟�K�)j�����ލ��5���zgg> ���j�܆�>�)#.�cԃoSeCj��yz���x����+xR��6�]�[�Ӡ���w֙ū�O�a�f[��T�D�Ege��5���z�a��vk	���[�Sr֡hPm�t�V�9�)��baWgx�W�y��󏵌V����Ǟlt��ף�iۉ}zx��`M�r7��$v�dc��1��N���Y-7��>��ũ<��*z�V�0�i��G�JaY�cj�1��Դe���r���'s����v��Ƒ�����,��'o��y���V%�x��&s�S�=6��J��+�����6�^��;i����ٹ������Y�lW)J��6w������e�`���{�&R�4����lzJ͛;�T�ƶ%yoi �W��c��uD�.{����2�6��U?K�o��S&�L��vz)�V�vI(�4j�Mu�WG����ϨuL=���L֯)��K�,��VZU���ڣ���vΑ��vߴb���\̝XjN��^EuY�$�֏�-��w:�7ükN����������J�m�F�ӛ+;�E�P�-�Ϲ��fu+ю����Oe9�����~ّd�׸��\g1�~E{-�:0��ׯqׇE^��!�D(#S�(
��pE�Otت�=����Ǜ;!�M����j�
��u��'/7�M�v�eü���j5|1�@o��h�=קp����@��F!a����bg:9�7��Ȏ	�]��3�_@��5�`{[�&<è�멑dޝݲ��#��|yu�9bt��#\=�f|��m��K���G�bq�]oH
��(B���'ϰ�'�7�_� ���Sn`KR~Æ�Gtv^T8���x��I�rv��A�.����#y�>?0Ræ 1����~���W7��7b" Զ
�Ɏ��m�!�m���B���^�����>��S�H0�98�|�T�l�妯��ű	^��n�/4Ys5�,9�zt8&٘�9�6�g�� _�UY%n�os>�=�Se���5aNls��P�g̖Vm桖5�E����[! c���]눖܄���UƘ\�8c.�a��0��lT�;بCᲜ�����WNSu]DY���|�aL.7��e�N�rnf ەQlsv�ŧ�;ˣF��t2o�_�#0��=ڎ�*���S��Zqi�E�7l�vRV<]o\qGSvCn~��%�K���ʃ�Y[�)~��v� T5(T\,���&�����*Fk�*=������vNG	��Pz��cUd���:[g��#L���)�p�J���X��b�y�6\�;�:���|F}N�7��3��CWd-9m*�n��!��[�/@�)~�OB}{Ϟz�������[�S�s�Ô���[�_s����FL��!�au�?=���E�Y/�O�1:�
X����or���8k��z�RY��kf�Y�.�nm`n-���h�GJ+��Z� �*�0����>��;�J}�C{w���{1T�1:�YA�2�?> ��4����*����L�/�O��8mo�e!�ox��6U-���k���A|�ӽ�G'�π$�ѯ��S	�����-z�vY���+��.4�U`Y��̺���MY�\�zzT�G�:
k$$vݟQ���ݶjo��������,�X鮣�(]@lɗ��4p�m��k�|��[��	�H�*y�\K'}r����i��A�BE�����H+��N�d\�ua]�t(̌>w��`�|I�]2��<s \az?���@'g�^j;���;��,#2�r�if�*5���2ƺ��:~Kv� 몋���1���8���~նe�>�
��kX^�l�ȷ0�U��l�,k���.W3�;���m	�J	9������ �l8��s��F�b�YU�s�k*�{v\ofa	�s�7w[���4Nm���T@<ݽ3���+�͹P����.J�L��2Y�.l*f����+�sP~�7��;i�HM�7���� Ob��>������4%����L�Ϣ��'��[��S؋/�d�{�6.���j_����oT���|��k��MP�F��N�*q���@'�$�wm����x��U�E�����x�:(�4-q$�h�,��P� G�q:	�^WP�3��0���邒��4M���:Cy�1d>*������"��N����ͱsK�7���q����c��a-{9�j⺥�����;����hRFsk��AP�f'�i����gxP�u>I���ruϲ�LpyJ;
��+/�_K+��jL���%��/�2�wq�U����a�*�M�Ʈp5K6C�.[:$F���'�=;�P�ϴ�6l�XRہX����{���@<���-E�jw�k����-��Q�i��~�n.�Y0~���b�Sk�#�VM��px�{� ���F�<�X[SΧ�.��Y.ڼ͍+[r���>\��sQ]A"���Pp�Jt#��Ȁ��m����^u�ǁ�o.���7��5j[���.$�s<������Vsq͘n��n�;�	�gH�[� ��WM�`�y�\��W�:,��c*0<ӤvZ�0)g~Ãx���2�#�zU3�������m��캂�+�-�vDm��Q��2{����F�Ц4������	g܎s<lJ8��LGFj�0C�_i���6<�.fz����C�}��S�U/��������m��~b��t��N�!J�i~�÷��T��S�&7ZUeoV4�������Ϊ��W�˥[�ʘ�upuxԕ͍d���{���=s�q6�I�C8$���$��rۼ�![��`|�󭮕5B�3i��/�B(�1��c���.��Uv��\6wq�ɥBU�m:6�4
�3����$�t��?�ݯ����ҥL,���y�-� ����.p+=g	Ta�dC+��y
y߹eS��81��kn��zQg��� e�8����8�X�F#v��8:��|�B˼���9��4��RN��n�����]�1<mlG�� ?�8F�}��#�����k��<�����~{�&�7{.�d����t������Nl,&�;9�<ye�!�͝@��<B50f��T��r��W�.��>�#�_���i�����-�Q�^�'��"��������Ml���~����Xy��9��M�NK*���-i����V(Y��ؔ�<|��11�Z�4хB���^O
�S�7,�,�&�NS<�{�6SF}��.[: ���c�}�G�������-nX�E7m��>f�! �����@E%T�>�{N�OjsH�wy�:w�>h�n�g�7ݱ#���*J���[L�\�λ�#
�Ӡ��4��D1��%�t��ή�:��drwXU{BS�$E%f�S�2̢�Y6˺-}���� ,`���:��Bŷ��]���a�\Ŏ~��x��M�8J�$L�b�-�FI�A�3te��c�9���bI9�%��nE�����1�m�{��+)2ʘ�j���Y7�A����PF�tvz>#�����<��9�7:ڕD���g;��**�T+�۱�Y�W�y�W�9D�? ��� KT�iy�H�S��gڶ4O�Tr;��/���%�[9y��1^^����1�x�xe8R��1܉���u�柂�����>a�pr]�E�6w7��Tn*iތ��b�����-�'��p1c�s���GUP�&��Ż.1v엞�3t^���=Yj�=��{ܺ���fb��;�"zO+ŊF墠����Ti�4J���ٹ=s��^�؉'7��jm�؎ ws�� ��-TGA����n~=�����x����'�Ss�y̸��+��7Cc��i<�y�ϯ�:GL��/a�q��`Y��7v�V���wUu�LT�A���A9��{
%�>�J�㡣˜o<����e��~�Z}g�K�u��D�ӗGrs�5c��c��MF�jb�k@~��Xͦ�C�l�p�وtD�?���q/sxq���*fr�⡷9�g!�6���n�Ou��"����-�����}���%�p��ޘ�����B���쨸+��_�P��t��ٟ:�"��%�m�-��a|g�Sp�d��w=�r��ݚu�t��#�+�皵��-��V|�S�gi/��R.���a��oU�R��x�nn��7�����Ff���GL���F�+��FB��T�e%�t��.Z�o	e�����շ�һ���~�V�g�3��K�z�Ü��4��B�� T5(�/,��|�ϵ���u5ә�����Be�����/]o;���O]�r��Pt귲R'��~�&�.�
z�W��b��֬�}:��w�3N�J�w'͑�D6��YLj2ͻ5��l�/Kj�wD��߮ڡ���+�iOF��H9E�Ӿ�jwCz�$$g%E	�c�7^������i�����J
2�]q�Z���g3b����)�Z�D�T�>�}Fi����/�b}Ӭ؟��%����z�μ@��:��Ƅ�����~*�˄�q@+|�k����aF;�d���f��a=Cs�V�5��;�~t0��D�+2cA�:T�G��anBFY�R�<�$3j���fP9�L�"?��$s:�p�i^nΆR�p���N�jN8�����D��ɰ�=�5F��L�����j��\�`�"�h�x��;c%ݦ��ן���b��A��r��芹i���!U���ة�^tt�bk.^�'�AШm~'�m�i��7�Y���n� �y%�S��q�b�;^��.�T���TSs�l�&�G�g˘P������{{B=����p���0���|��{�|x��t�~Ǧ��e�Cy&u��ܼ=��3!A�q��qpj��/�3A�M�۹��L<��$e�2�`[[%;vK۰���nԼjE?,��ܳnUwh��l���egK���).�"%d���	{662/�?R�6+�������5��1�:��t(k^Ȅ'�j2΀l���l�]dNfDTvQ+E"�����;,�u�P��9ͅd�;.;�0�Ĵ��xw���Uc)����O5�@n��^t�p����L��*�¦����k(qwŖ�5�KN�	�%��Rg�zv�k��g>q��3��^���0�(Q��ް�:�A��W7u�۷�4�C�Dn��������a7�����j"��䵷+�O&�N3�rӽ�:�QJ�m8	�.���]>I� R��q�>l� }�S��Gi�0&�/��W?k����x����c�C����ވi�\�];�j�V9U�tH�j�A�Lu�O�g����ĵ6�f]p���;-2�\�c?�p��20��iz��g�/��S�ㄠ��D�]AW��p���m��أoJԽset��-�{8)���;>��t����"yU0��A	sڝOE�:Ogd�I0�cl���X�����i�?a�Q]<+���5�I�Pʍ�/�hfi�q����"m�1=V���ҳ�g!��(aƩ���;KͶ{�fG���hY��ܮ��e�9��Tb����b��x�C0�&l�R:pZQt��g��#,f�]ԟQ�1���q.���Ӷ�c��U��N������ x	- ���_;r {��ީm8�.фɶ��.!9^T��-[�K�.k�;��z�;��4�5�d͠�֥��p��Y��zA}�͇/��ȅ����U���fy�[��f��E�V���v�Lޠ��b� P|�uf�S�A�r�f�k�\.e�ֵ���7��ۭ�)*x+H�91�w�Y��p%\��	�R7��D^�6n�C���I��r���ݹ�#����i�v�����vz�z��;�[�8�]��R'gh���7�\�l�=�t�%�΀�sf�F�>"������蓮��h��\��3~��ݠ.�V��Տw��������������g<��\�"�Mͭ	��ծ���{�</�%�O-������!�9�����Fܬ�Y�� �PJOiꃆ�5&��Ooen)pwn��:l�����4Ⱥ̃��9�(Aر��ؒ�N�i.��U(��ϋ`/i}�$so��9�sG�d�)��h[% ���	2lxp��{v�9'%e�ć�.M��9�:7`�P�Y�7f�����74S�J���C�/!��3�%�f�թijG|����)���Kh˧bd�����,͏��[i��@��&�75����ҋ�2�ڱ���y1]L�����N�\mwZ�G+_�d�b4���� F)ǻ[���<9b���r�i�ald���;mX�K&l�vF姉�<�yJ�Pf�='5���Wh�q|��;��6h���f�A��ys, �7�9�I��|X���^��Au<_�Ϊ��<��Y�x�u�[Ҁ�d�]�4�\(�vt���� �V�R�jW'.����id�B�� ��_Zۂ�7�rF{v/�&��"�&��;%7�Y��vhdT|�X+����5ٰ���N5��5�7{{g'�T��5X�W2.��*a0^N����m5&����5L��܊2ح���̶�bΫx�Hi�l�ݒr]g'ƭ�gp���51�.��^�w�ɐE�[X����3u�\oI�	��kÊ���y�Bם8����x�s�� +�|��{{w��($�V��eER-i�J˘r�'JΩG,��B�W=B[�NzXF\���a�m��q�M���q�v�|�Sf>�V3�q�#�����>7�h�T�e�QO>B-�.oU��[��F�䒡�]���ʼֿFz�X�3U��P�$�o#���ئ�.���
�U�;��F;���v�pB͕�ɺ�Ŵ��9�u�T�v�i9-���)DAWb�76��>��{�ۉ�6n���ݸ�s�����<���|�Ǉ���R�8_Q܄��K&ʘZ���{0���|�>�(�O_h�6\B�#�t"7�'r�JVN`o�HtT��6�d�|��Ϗ,PPW�A(�*.�W.EU�#�TM2��&]3��S(�'I�"*�ֲ��e$�Aa�$Ȫ��M�<8�PQp��
�J�(eE���¢�DATʉ����A<'"�;/����r���e5�W)��U QL.TAC.$Ċ�\�Ȉ�I��Ls��90��t�Ar�kN'._�����9��X�(�U�(�*;(�9�
����r.tȦ��)�W*��- ��G*eT��I�&ANM*"*�$�wnQ�T*��s�9糗
��C�EU�D��Uӥr�'�J��[/�.hx�]*
���(��\�q+*i"��$AE��5*�ŕED�3����H�Tl�$��QȸUdSπ�/�M����Hn���@�Y ��8����ˢ��<	�����i\�����/2��N�,7󙰾�\z}O!Flf��Vuc�=��݁����~,R1O� wE��Mhd�7��m�l�ϱ�hS�A��;�j�����	m�î����ҩ�J��Wu�l�nxYi��B��E���hQ�Zn�:ّ�g�hԧ�U��VE�kL/4U�v�� sNٖ��%'�@η���4���1+��Rs���m�L�C��ev��wx���̪閮A?1�@+�@U��vXs��8��v�T�0�U��D�:���D˭õC�@ܚ��4����`��N���t�oLt�4l:w�j�:�W��ۮ�%��R,���t����g�z3?W��c�Cl6��v\��:�*�?O��.~����&�[+�PZ��Ӊ���uꏮVI�d�3i�_.쎖�,��CW����.q��d4y���3>�y�3��+�q	�&y������a�L�oe���<�Bm�)������Ov<���{.���ʇ9:���)9��>|�:�7{��Y�h3����_�5�����},� �lP�S�9}[���J 3��UW�lAs�*8W���(K�ue��k�W�D�$%; �����۲�j���ϕJ�2��7@��?*��nM�*}��g�_c��e���N�RiH�!�Z�����Q���Lbϊ�B�@�� �j9˲�ZD݋�n��+�Ce�gU�=k-@/`(����9�^��lP�2֬�	�b0e?E�:�����NS=|�e0�e��n��ω�+e#��^�-�8~1�����Q�^��=ײ�{��鞻��*,X;M45%T�-N����)ô��鍜����2���n.7�͝24v��:ʝq�(���]�od�/�>z6h��O���l�۽�5J#������z�+�BB��l�*γ��)P貮掓t�}��4�V��+����N�Qj_x���#�`r:��&���;���6¹���1�1�Xݹc��EƧ�o��F�*�*
�������'�s��9t�1Es_%�w.*�9��[�"G2S�b��e>�'��pǯG<�����z�k�\a�2kλ�E���-m����x��9,���O��H�Q
�s����S4\q=�b���TJ�w�����,�=�UQ~�+�s6�L���s��M�n�r!�\�1��_kQ[DQ�O�ݷ{Q�5����ۮ��x+\;*l~�v�<�y�ϯ�:GL�	m�����Y��4�{�.F.)�^��c6�J]E�a�A����O �>�R}�n���6��5�-WY/n���ˀ�+=��)�ܦ�m�5��.t�-ډ�2�J;j䰍�w��})b���F���c��nkn'wovK���掛���z���tO�8\6��y��C,��K��f�X �KE,���KM�����4O8�˂u���-Oe���;��/p������9�J��^�Ov�f��Gh�FK��.�S�5o�-�j�YS]DY�+�<� �?	��M����n�\�~��z�;�eF�˪1̷kȄ�ľ�{
̺�"���)���-� +���y��-�x�]W��a\� v\�J8b5�ڋ7�g*r2��2+6:@����Ocd	�S-C�7�T���Sp�k��v��/�V͝,]o;��>{�n鳕ţB��)���pka�'g���8�U��yѻ08��wB��i�і�~���w.��T�~
���������j�[��|o$���|�8�n�<�����44�*.&��jwC{Fр�]���'C���9`CЦ�17�j�]H�=�P�&ғ)��trϲ��'��	�}F�Ai�d�8�t��Y�^�u�#g�Q�7�L��C�Et��tUYp���@,zhׁRϊ��\��얺:w�15���
�2Ou�G/��ߎw n��folǸo� �3�(��\��k9;��V��r�=�e*�YA��j8�<�JU�=�8�p]�>�v,��or$��n�vj� -k E�s_ш����)�
�_%W]�n�N7��[Y����F3��9T����G�{!i���=����3OJ�+Ǫ:
k$$v�~ߌD��~�0��V2?(h�Pc����h�q�&��x{�w��q�g�a:gԜqS]RD*�PtQ������Z��.��`gd��r����p��U�b���6��{���5�#����:�e�S�Ae^[f��S	��w6�ڋ�z(�|��rE��W/����V��,���o9��d_oL8}�E��n�s�C�,k���w�@�p]����m�t�=E֟i��x`ڨ��s�,�tF�N#���	w��@�4Ǫ ����
�����\��~s�eY/pˍ(�5*{_V���x��D5���!��"q�w���TH�Ρ7��Xi�28e\T�Ve���^Z��"Tӱ݁9��.��ll���f������_DXy�u�	�~s�O1�Y���#L�K��ΐϕ��6�Î�)G��_<���eSz9�^l%�L�.�'��OE��X���zp�S�s��UVuU��������G�bp�9-8��u�B >��>J;
�r��hj�}��<D�7c�ӏ�i�3�	�ܬ���9�}�i和��7xIan����o�/8j�E-�s�|������q�W��a)н��|g��$��]�G.l�_Qa��*v&��������d�0s����䶰�[�R��¹Tx[�tY��f�a�'X�i���a�'�?].�ʥ�ӽ�p5Kd8B峢D{ml����v�r�[r�c[Y�Ӝ��<�b�g��4�>�v����y�*�y����S��M��,[}!D�ѽ�Vs�I�7cޝ��C�譛�pQ��!IP�X���amO:�5 2y��+b�+:栭	��.۳�l��l�.�����\D�lJ*�����*hفZ��]�c.��M�8�`s'�x<��;-O!C6lf��Vu�9����L6���e�F�E��xm٬��̾��c8���S��9�<�Ӊ�#�~ÃO>tf���h�;ohq�5mh垉��mU��y��	b�G\�*``���i֛�f�F>a@��sǞ�������k?<���=��~�/��1�P�XN���r7��õ�4Һz4J�wL�l��"��'<���+����R=�y'	� ��T� N�E7;��;�;4M�s¬��Yb�2<e&�S�+�7@v��7��w��0S ��1~���D�M�����~��J�wYX?U��i]�b	�(�M��S8ژV���Gម}��h��޹��k��<�N�ƈī�y��?Q���(�܊���b�����Vn������N�^#�摅�e��B�i0/�"�߽���NI�����o�B-�>�2�(��[�0���y>�Z	�u�N��5Jq~�+�E�O�:ln��s�����+ٞ�.{�yEĳ}�(�	(��:��̋����/�3�"��3[��3���^=p���n�0�+�~~��bٹ\�jI%
)���]t�^�&ߘV?-��A��/�<����[Z~�����#:����D�sRP��Fn�.���;�gP�<����;��g��45K񆼚� �e��f������:�\�Q��;��e���0�f�2�����Õ��g^�9���9L��w�{	�������%�	Y'1�-H��O7d ���Qyd�-�rS���b4Ku��ӃW��,�~I��4�Ѿ���E�u�ԋm~�N��������)l��{S�T댨�����7� �e�T ���Z`��s1ӏW���u+H�@��>�&�p�%��i�ǐ��!	Ԕe��P�T����eDu�pzt����hCvQ�=���l�9D	j��/>jt�Ϯ�#L��G�?a�o,�-J}k�	۱����]��CLj�Z]��i���2�k.9<�ǟXvSF�
�i}��j3
����70�(;�_��̟�}&N��Ov�9G&�(�y}L����KX�k�֕؅$�ջө]�.��d�M�uzsUn�t�+��\�y���6��E{%��ܓ�9e�4�k}&t��Y�-��\�Α���6�*��Oޯ��e��qBJoz�=/����[����}��,��[��}n�jǯG<����D�׸�z���n���eر/��dD�o�j��{�
v�����R5�$B��O�z$�}G)��������%�&��N'˫QQ�&��vCt��iqNq�@-�RD*��#]�ZGC�l�@VL䵦�3
�/2z�����sZ��9L
�j��X��1΀y�� �鎂@����Yu��e	[V��9a��;u��3*�`�w�G���u'��D?:�\�y����;�-�>�2������E�9�=)���Z�u�&Y][�YeMu�Y�>��p؇᭛Q�����q?���5┴��)ٖ�{�6�Pg��C�k�G������[�y�w��\O7ս}���q�Z�ޡ����A��vT\f>ޡ��� �%c�7]9M�oQo�U��6{�r�f�#qo���8.;����O��f(e{��4ҷ#,Ϲ���y�kQh%@��1�w�&9�+������Z���ϰ��R����/֞��島���od�obv��jh��@���%iď� v����y�A�T���Y�)y���*+�r�ә+�}ϴ.��e�xɺ�Smm�a�[G@Yj.a�phJ�V,�s{��Y��2f+��@��43:m�\��%uK6^
T�Pi�@��vVn4�f�]��ݙܽ�e`:� ��(T\M;��~ҩ��,��!���P��{T�SmF��;��V����*9��g6�i�$B)�:tiP���w�f��ެ�	��#�]��䅗�wa�iCd�n�R����yEN)=��\"�N�Y^}���0Ծ�4�Ӑx&����k0҃>=w�Ofo�
��,��%�z8I}��v�������.(��a&;��O�Ȑ�7]t4�n�*��ۚ��]?,�m���3ea�i�؉�R�S�s��HH�����oZi��e��{�Zk*wC<���k�~���m��Xxv�i(<z��P�N�Ή1�9�/�w������׆X6�����ء B}�[�P�����q���?yfI�����b��h�MS�1�{��`���2�t>���rE��W/i?��F��=��X������v��du�|چ�p3����J�0�gZA���g�%�r-ͅg��
��3W�(�Ô�2��Ə7�8���Ƙ��!�zz`<�X�&�b�YS3[��03:��R/~KV��p�o%,����݅]��uĠu��hmC��Y���;1���_���Q�4��N�x�d��k���`��(���(;�rAԪ�u�g��om�[an�4;�WF^�.6�7���+���JƑGkj)Ge���������p]�a4#����Θ�p�tG�
�C�sAˤ�����ɨ���>M�U�ٞ��c��!���E�,�1�7h2��:���"��w\Ж�~|{���-�f ���wvW��,���t��n��=^��fӋ�����,#��\�-���t�Lߗ�X�
���^g"r����&{��(�>�m]��z��L�p-Kd8��@P�'�)Eg.}�2��*��@}���._ph���u��*��g�=�:�I��kS���T�8B峢Gv1���A���H~����t+�4_���F�dNQ���?KPIU3��g���x�ݹv�j���y���M9Z/ĎӼv�B5�V͊l낎�8���@,zf����	D�)^wy�!<�o�bkq�n�)�3eq�4˟�ϔWO
�ڇG-8
��oSa�]�*ޮ�{a���y�&����:�Gu��Ә[���a�"���z[�eB��N7+��<�35�|�%G�� ܦ��,ϐ�Ц2�C�5?#���k�a�-��uՒ;S_e�{���n��8�sT֝[r;˸p���)�ֆ�k�E���Q-�m���h��Z"��;S`��{x��,�ݶ����ﱍ{�>��o��铅� Ľ��>M� �H�m־���f��e�Q��K7Si����J��lfv���ʿԺ�"äe�ݟ�h��b[��hQ�Zn�:��	��G9���gi1=�=׷[1W�s��!C����{�M����a�ᦕ�ѢW�`쨽=�~����WUu.:��\�XG�y�s����L~eS� K�vXs��8��tL�sy2Z������Nl��w��'Q��b��n�'�;��9{�H�#�ߜ�B��D��F�}Q4��ض�M[��W]�6�O@�m�A�eއ�le�s�˘�7�:��?>�(�-A��ś���r�d���:2�"��f��/�p���nٰ��~�}�x�յQ]p m�9VP͋ăU*6	���d�]z�+
�Om��mxDl���Qn�U�����}�v~�o��"���_\P�d�FY�g�n|�%���e����-i���� [ރ�b�TLuS[d+P�W��:��Y��:+�����JSߠ�Z�b�4�����	�'��+��­�I8�4�B��u��ݰ4�]A	�(Ǝ�{���ۮGD5e>I�[p�Zm��M��(ң����V=��d��ރ7��)R�����t�R v�eN���aɰ5H䣀S<_w���b��R�#�}��ن�$���ѹ��;��o�1�%R�ͧvU���Z=!V-i�9N%3]4���u1�EӱCkS�Y�
�s��$�{
{�YsDձ����ڢ�ř�Z�I�޻jT�w�=��K�BGhJ�=Hаt,��f�뢎Ac+t�w���Vn��<鄽ݎ0:'a����Tѝ��1���{t'0�3���.���*� �r�2��M�@��qD�֭����,�ݖ�=�'7�k���
ǹ�Gy�/dN̖
nR�����QG����7�U��]"̓��;V�G4t��{�y[�Q���(�Є�A���A v���g��u���d�����I�J꾾��'�vh�[��j,�ÏR�����������SMֽ���)���w3�MwvE�*?��kvG@��+in�:���Ns��g,��0]fw=�ONk;;��0����m�����ޔI���.�K�w\]�m��R����r�n����n��X�D:�E�w��憇t�uŽ �����P�J���0����(��vNV+ã3+v|��}X�ʝA#k����m�˷��0�1���[�G��k�&��8���+�`�5Dȏ)�+<�gw���y�;[�GZ9ø&��[��¥���g��a��}�<�o'5oU�ad�E�B�w�uXرK�qfO�`k���ٽ>��@�5^���D�7	����컇\�!�R;��K���-�qYu%�8b	��R�&�;��^����:��')\�* kd�.q:�8���ru��f���w�&���y�ci�~h��;x\ٛ )��,���WV�S��0��i�C�������dŹؘ��AL%�����|�l\�\4�7Cxح�.LuҚъnj���u{8�s�Ӣ5=��ީ��`c%�nN�{x`@�a΍�,�7ǹj�4X�e��P�4��	��}t��O����.�:,#6��q�{g�(�W��1�F� ��)�K7�$
�!_�+)�F�*n��:p�(L�Q]�̠Z��;Dxp�m�[�ɓj-q��f%j�)-��jl<-�E�ih�`^����ڇ����R��z�=�b���鎓5��T�06���s;n�Y���4�����z�Ow�z�K�=�W�W����X��z��2�Rg1�̰X��&Y�n��Uꗎsf�����ý�5��ߧ���ķP����2�s�y�����;�tp2����܏�:u�MCj4�`����o#Wnण�d}[�<O]�޺/C�ܺp��7�9ȸn=D(˕vnm�)�rZ:t�w(>yj\��I�]�\/uQ�Z��kױ߾�# � 0b|d\.h�9r�������\�*�Y۞8�P˲�7��ʹ@S.\
*�(�
(���(����ʢ�]*HN4 ���We�Q��˰���Ȉ��ӗ"����:2�l�U9��P�i3D�Y4"9L(��AvUPʠ���.G(��Q.PD]�e�"���9��J��
���s���v�Q� ����5�
x�".9�
��
(�m2.��tiTG
`Q�9S((��D.�

�v�&PaDQ����Os��.S�I�W�*xtx�ęC�0.����dS�Hs�xNAr�L��t��W���P'��
���	��-��+D"6��AC�+w(v�X�i��	�̸zl�M�o�jH��nȗ��l[��\ۛ`^E��U,k���>�Z�u�{�A�g�;�;M;.Έ;��w�v��`���#OL^��\éU쪌��!�:p��m4�	�u���K|�H�RQ�kS�2̢�Y,a7������)z~l�y��`�iہ��[9�hRg�(c�H9
�R����;4�9Z�-�p���R����[yѵoen�"y�T�6
�uO���#�z�Xw[D8���ݔs�0��~�A�}��;�uB|���Ӽ(�ua��~��H�ҥ��ts�&�R}�p5c���25���q�6H	���j�F�i��jӸ��=�FO=�����WL-�T'"���B�F墠��5ӌ��գ��5ݭ����F�)�M�z�v;v=�i�W�p7�`�ʢ:�r�;
8F�?<E��N�pyXi�ɍ�����������ٷ0'Ժ0e�G�2�Ϯ�y��s�:<ò ���"v�"J=��Fr�d�2^#��M�ַ��a������W�x%�����f�żz �WE^S��Y�کa�Z�,3.�a�7'���-�e�,k��2؟xk�8F��
��Yq3�:h1k(U�`V�
Y3m���+���
��ڸ���5x}�o<�P�ޑ�Tt�cr[��xv���5�	5���ӌ8Ʈh�^�G�f�}�P��+V9�l�ͫ��t���	��ά�f�\�n	q�q�!*��������f�sȉΰ��c٣��9��9ʞΙ���������i�g��6�PʥގY\q�\����6��,���4y 9�NM�bg��~�;*.�����3��e�dR�Ӕܰ��y1�@�@�Ί{H�>?2<���m� }�"Y(��mE����|2ܮ�ȭ���u��]���,u�@�'S��S�봳_8���\��y�8�O�]�LLVf֘{ޭy3ۀ�d�g�i�d
��
��jw�g���Uc�Y>��"5l �Q���׈L3:�rKL�5�((�sv4B2��Jz��%B��Z���t7��3���c�ӏ�:<Eh���z��	I�m���_G��,�9t����)�Z�G���	j��e������u����NE�͓�|�-u���ܮ�C�WO
;P課�'�΀X�ĜS,29���5��|3p��ߛ��s��C-n}�������OOO
8��H�!#6����w2��_U��M��@�#����M
�����u�&�M��ì�*��*}]RD2��C��;k���t�Y=ykM��dF�_\���^&2�wb'�)LV�Z�{R��Z�\Q���؊��LL��җ�{ė�[w~,�g��j��3�$܀����]E��E�Ww=.m>��5wwgO�*�W�ĝD��Ν/^I�e�J�H�;����O���Y�l8�oWFP���b�.H���B���7`�1��:_c%ݥ��~SN�w�U�9�o���c��yR�r2b��A�v�E�#�J���R~�P��k�<#m�L<�T_r�����Wy{U��3�6WU0
��_�`vᡛ�<�V~/~4��ǘ�����̋E��s{�h:;v��ڠӰ�ϊ�%OC��4.�N�0:��Eܲ���4�J�⪜��y��}���_��t�2��I�k��=�è*����(V��.m�9jU����3��.�dma":�UfƄ]�����K� ��+��?vĈf\�]�a����M
y���}���7)�X�u����+
�[Ћ3i���a@?������a7�����Z�G|�;��-��q��;�ƿ5݈�4���B�*�����kN��q�-���c������3 d=�ET��Ғ9�4.��Tޖ���fY�B�U�!��7�*�M�Ʈp5O�!w��U�ڦ�zDW8�ˍ>S
�S6��+��h��	���GOCHIU3��zH��G�`����&3��j�����^>�Ԓ�c����J�Zc2��R�7�+f��Pۗ�yT��g�?	[ۢh�n�jWj���*Rm�o�>�\�b�6GnܼZ͛�;\]�����Ӱٻ�,�@>�3���'+��>�%��ۍ��yI�C��<<�y��Do>��r���b+:;>����Tܭ� ;�?���@u��ԭ��|	�7�;�0��	s�K�Rاh�\v�����Lv��ʵ )7՛O�]+����9�72�t����r��S�ರ��xig�8�,7��v�(�9�}����GCu&@���s.�J�k: �E���t��h�����C��q5d`ST��<.�~\bo������{t�Tym��!;1R�9(O,�X~Fm��,���c��$[u��l
���b�� �<�񮜩�ڽs�ǘ�rV��:�e�C2�O,'z'�nF�=4Xv��Һz4J�w�`i��Zf��_�V^��˔ϧ��G	���?��#�,������>�G[��yt�'�2ۯC����'��g8��;F6�CgA���o��s(p3���8G_%���\O^�l��g::�U�ax�VK�k(tle۱���Ƹ�؎AT �/�&��]U,�����o���x��e\T��̏������k��?<����a6�߶��L�.����=qz0��Q�0�狹3ߖ���0xin�B�����(�v�b�̀s
�ժ�ɽy��0gKb#;^7]!�:!�o8ؘ���,@MB��N�����"�G��l[��nt��`9m��;8��R|I�l���NE�������WEu�4տd�]��(T���i�c�Bm�3�(���S}3=����;ˣ��f���gˮ(O+�i���:�cF�2k5�l�D
���l�\����P'�U��i~mQ�W'�pq���	J���g�g^�9���9L��;[�L�o.��w��/̏0�2����: vm���dp�k��Nt�ul�1Qb���httm���l�� �f�UL�N�����7��Ιͧ�>�RW�ԗ\���ˡ����y�qpzn���&IR���f����DKSΔ&�֞�c�Jre
	�����̩�����V�<sDm�al�)�1[ %M4zr%�_x��S�vi�r3�cA�׼{ E����o���EƩ�nv��VI����ѳ��*�*
��O�mㇻRتB;[g)��[g�ώ��:��� PxΌ78�)>x����x-��T.&���r�7��h˞ȧ��t6�9��Y�9c�`�% pR�]RD*�PD�Aℛ��R��}�6�aV�?��������:�C+%?=�J�{:ͱR������a����z�iܼ����c̓�J��z�5GHuI̺��_B&��B��sA����`Xl������XtFm���u�tPͩ;�kN��!�5����Y��ʚ����8�Y�By�H�%Q���n�{��,m��pc��b"{�w����tk�S��e�x��z&s��8����0&��P*�{`;(l~�v�q����Öcb��(8�l瞝�����э�����e�L�x�w7����=�Z?>_�mD��u��K�F�t�[�[�VftAK��D����`!d�qˠ�|�y���E�]Ga�O��3\!�;�m����ѭ��7�w�ܢ:�9�f�Ƙ����!��o@�g�����UN�v�_���w���X�{U����s/�рP�	�z�'ې��ʋ�>)u�}9~w��J�"bK[�b<<JȽ��� Vs_7TE�f��_<��� vm�!'�h�KЅ}r�yS��v���x�ӥM����n�M�(נ�(����_�-��٭8���_��(`��#֞[�\�^�-�!ǕVIU�#8�]od�%uł��$Tz�*.%��Ѣ{J�B���D{V�Y��smo
�`�V�Dіsd5��G�NK]2W/���cD"Q�S�4t��Iq$�;N�oS6D������&���:���=���8���v��o����jY���qѶ��b==�i�.�Kk�)N�v���o���@���r�ѹ�o�Z�a�ww�Wz�s oq�zu��&[G�m��$�ԅ��3N2W<-`�.���u�rSƩ�y���Sm�y�v\n��N����8O��)l�]�P
�e��3OuH�}G'c�qK��^�|����%�����Q�Q�4��p��n����6\$�ǟ@X�ѯ�r�y0֊ep��#'�d="�N���Օ��tשּׁ<�v�ҥ
f=Q�SY!#u0t�m-�\eT-����M�GD�n��@�Ea��m=q�y�v�=)���!lX8��7;l�s�4�l�Έ2��y�����TwE	�*6ͰC�ّ�����%?}M��)�]-��zͼӅ�����WT�<l'��L������r�i�l��lq<\���¸Ƴ��=N^0��c� �Ξa�uS
��XK:���������n[��-�zʳ�\n�j*ۓ۾�ME�J���0w@{��`��>;;�1U �p�q�%�I���eZ�Ι������y*�dk�C���\6�٘�-��g9��3��%�Ĉl���8⬔�2�bZ�lL����1����;��«z�yk+�se���M��&�����"��u����Q����{���'�em�r)S��o�Ub��2jw˚��Mݫ��r�4\ʝɧ��-�ݼ�5o
�}��k�b���#�w1�yWFs96���g
�G]�_T�5}��n�)���k�~��u�;�%x��G�p~��d���_Rlq�-.����`P1�\�����+S[Ћ3i���a@;z�U0�c���2�R��4��:&%Ğ��|���S̕�Yjea��DI��RCWD��Mt�&}i���GU�! 3+_,]4>&��O��ˉ=����0�O"���/����F��6}�XQ���\KS��p5^]�9Tڲ��־Y&x�'��#��Pzh~��ڻ)�A�l��H�r #��-�E%T�2!��D��u���^�tI��#Xb��Ϩ�B�8&譛���v@�t����d��f�l�X�r:��Ϊa-O8����Z���u�i�=d�:��R�u����&��� 2����I����t�yjt��S�Q����!a�,r/��B�V�~m��լۖ���_甠u�Xq������lxm�C�U�Fú�c��F��yB�_��˭����a�q�/���5�n~0�Z�i�Ϣ�	n���F�i�b���u}�i��3tѽ}k���6u<�O)��U1ʡ<���<�Y������i]=���0{j~;�Sft�j�i"�iA����	uA���ͭ�w�u��X6)՘���|9p�LS��X���}�Zڢ�� ��l���M惼����F$w0sb�Y�yy�y����b�ֶ��w����;@�ʻ�'A��k<��1r�N&-ry����4�1O�<��pg���y�%��;�$o|�C�2�r���vŎ��T�0��Xk��m�쳜���xϟz �
`m鎂��Щ�˰$l6�F�h�Q�O8;��7��F���3���Yw����}�睗1<V���	_�咼�������}̉d���S�pɨ����za�l��^.��FZ��3Ǉ^d�`m�zOc���^Į��ؤ�8��Mϟ�[���+
t�fm?|t��g�j�e�n��@M�P���穹�[��ء-��e���6VC3�p�}u&媍�v�1ˠ��ya�Vۼ��EwF .=� ?�<�y��W(��o��d���g^��
k:^� <sM�y	�����/�l&���K�����^aGG��N�XW��K��Z�zz�;��l�%2�����t���=ӽ�ڞ�GW�:hK0�O�eS�3�؝����A`��)��27b�3��m��:�A;�H=
��y҅���Sd!"���.�F�m���+	�\���.��S5e�B����"��W�T8i���N��K锏p'D��]A�z�3�(�o�C]��]3T�r_,����xO�8�mG&��v��Q.���o���yG�z^V��.���f��9p�@�s^�<r��n���6+_[XtI�(���
���W��:L�J YM4� L��V�WqC���C랂�f���׳s�9��9~N?�OSp��v[���I�í�H��RAZ_d�K�w���5�b��(�\�x!>~|�>��9vA2zT�̻���r��j@w�e?ɍ�{ظ���K3����r�<R��z��n����=}���QC���LB�3���F#��nn���!�:W�Y1��M��:��Sb���5D&����4�1+�rW8�� >�#�u�k/eU���\��w#t���r� ��M)�0'ԟ���G�dK)<��:�E�2���ׇ�/rK�0\�L
�9`:�%�4+�GM����s��D�G�ׂP�P��;Y/��n�B+`�nn��Y��X��Srq��O-�V�VYW����8�1-E�5U�k�1w]UVo6�t9L���H�k~����22M*y��E�'�g�����YeT�V욨.�V��bN�tABѷ� v�Q�Y�޸�܄��eE�����!��?@eٛa�����1'Ax�AW長\w�Y/hm�~�}�"��r�6�)v��&�Ҿ{�e�]��q,:ؾ�=��/�
��f�ѥş�mk��MI����cr�<�⩑�(�q}�t�T���Ve<�: �Ӕ�뫮�u�7ó��Ӹ`�-U��˓�H�Pº�K��k��6r;�t������l-�O�DrJ���B��9a��F(�3i-ْ�L���CB���y�����������lh�\�;{D�n����K��Ҟ�"���L��Q�)ŕt폊܏{kr�|�䧉�0�a��5��dU��+��E5�]䄞�wR��I�(��e�_x��Ko23�W�	ق�'\Ӷ�0��1�MP.��joj[�#8�D+����,�9�1�:L>7�F;B.��~�!���#��q�ioz]s���f�����U�b�S��Ԙ���z��DQ!�=1v�S�v'f	�y��QEmb܂W^_q����g3�t���]�X�r��}Dۨ���i0�긓y��9`���ޣ���jiYפ�U ���
i�G����7
4�����<S@*ЪUf�6�n�s��2�+�:`�s��,;V^ܘ��G��XSő�d`���I��
ӉO���1|oct�Y&٩�v3A.�gk��dξa�Z���[��H��wb�˛�yo&q7V,��������������M�9Ϟ���ٷDЎ���Ҥ�MU6k�G��o�:�L�)�E���hA�w+*�d����-9R��ɝVì������B��C��[M��d���N�;$\����,YR4i��ʼ��D��
�kGG_P��o��Ǯ� Ɂ�=K��¥�h$�DS�	�v-\���]Ձ�[z�_$�.v.�t���{`8��sQ��F��Ьs��9�6[���B�����e�|[;���F�*���{Rw$�ɦ)�0�^��g�ʜ�<��wg�wr��L��E���|s	}B�A(�*�M��sL����[�@�M�3�V.7|�|���2��|if=�
t{�*�1)��<�a:��g�]["���C`>�r�;�a�Z�J�Ŏ� ���`�OP�=:a��8(�e�FrRjb��xF�`#P|�Vּ�k"��M����tZ�t��֏P�S��8p멣AԹ�� BvU�YIفE����S����;|�Z/�
�-qgr���&�z���3��yb�ܭ{l��є6���W ��X�{��N���-)`�4:Q��ˮ��"�;�n]�U;`O [S9.��v��oC0m���Ϥ�d%!���-7�>�'��y�K���WWeѼ���Z�^ب�A�	P�����S�[|��0f$�ل}�}���	1�yӹL���\.ϊTa�.܁
���L(]lN:�$P^q.q�q������v$G.e�)̀�@�k�i�\�(�S.�L��\"��B��<Ȋ�U
dWu�"��S
dz����E&%v�T\P)�)�\��]�ʢ"� �EPv�HnqH�4�@�s�쉴�;e�'1Βy9�����l�&v�P˗aT\�&$˲��r���!<�pL�DT]�9��ʍS�"u�v%vQn�9W��78�t��8S
I��8��N�u�����J'
e��'D�T9�^�{�Dw#��-Ck���`�R����r52��$eoDo^���1+*�|�`�b�}4�;K�U¦�0z�;#SA�vd�����~"�]9L����g�_f\6���+���7�d�>��Ӷ��gZ�4����2��*�"��A�^�E
��/,��|�6�Zyl.:�إ��]o;�f��i��V�C�{y�ѯ��^�i��e�'��[�)���GH�Qq>�{Fiߴ�f�p�[#��[W�����d4��������ݕ8�黭Km{���k�i�4�e�:J�E�Ӿ�-N�o+0'v��gT���c�,=���+��M�}��8V�-���a<�ӠS�0��$SFl��&�:��ܙ׾�<���4�/�O�F�b~��(`����E��W�$�Ǫ4O�yYoz"F'���_b��_>]�
1����k�eC)fލ�6VG�УB=Q�TH�:�ګ
��jVԚ�-�%�X�g�����-���0�t<��uY��Y�;��'L�s�[j�*ܥ��r����OE��,cL$h�����i�(ʍ�w�P�����{�v:݌:"�U����T�Y4�E�e���
k���*x� N�u�O��^��,Dҹx2ԟ�eB�q��7�g�w�n�>�;�X��Y}�s�b$�$�?g���W��u�cr=[딌��z�d�Rz��.�{�u����h���5�2D��_we�$��)T��|)=@m��7^ъ]����<³�����^~q�����wXvu�Bh�=������w��k��M�nǄd����p��L2��\v�1~�m�/D�E�9/�O�+�WO������x�3��%�d�s{��P�o9���c���.�t@tРq�.~Y!W#�#��T�9��J��KՕ�=g�����0ͳ0���e��ݓ<9������mMF�Q�YU��כ�@�G,��ƌ���
�oQo6xqw��o:�D|���"�چ����w��#t��m�jću�;�d���x]5�V���e�8�|�������8��e�Wd�tUQ��~�P�}t�ZY+�i�����)��0�ƺ|�-i��9:ꃊ�e�UL�61Ͱ����(>�g�Ej�u��iWbg�'i����%R≾4���cF-~U[��*�p���E�tH�հ��(�=M�����v����dO,Ξ����jn��=�3@�ѵ5qL�m��_3��/��~��PZيhN|�k�5�C����	l낊�pA�~O�.��e9�Ҟ�hG`N��;�L'����\%ϐY-�)�3eq�4̹������sJ��G��-eq䔽{Z��;���n�df3�mN���[�z0Wd�S��6(=^�rݍ����W)Hg��֍:��ѧ!Z-3RJp�IDO��t�6�4o�3��t�#5�=;2-a'g%��P\0܌�ʊh��|1ustG����p�e�g7�)wu�&Ӎ�3Dm���]f�y!Ӳj�q��^�Y��� ,}�l����x>5:Ge��r}�Hyo�%�����7U����J�<�NK&���gHͺ�?C���ThQ�i�����*TR�&��tf�
����ݮ����#��K8�]�ʘX~F}nϡeE��SB�i֛�;Y	
��:--��=c9��Ϲ	�(�7��,@v]\��[\w<1�"�^������0�ˉ��3�����׃�Q����ƙ)�'�; ���OL u�;��I����qwֶf��s���꺒�����D�1��3gA��� ���ú�˫6D`s��)��b�9~h˒N�c�n��pu5�axkt,�Ŕ;\;*f�s����玑g�qL@�=LY�j�4��]3ⰻ�6�o��?�~F��'��4z����g>��
l���m�.��Z����-I��O0WQ�����܈���<摹g��O5A�db�?\��gK?�,;E��淠� z swTh{Ov<��m�qC�ь��~qG%�K2�Ӓܩ16���J�x���&чBzkGr��[xE�F���w<�S��i.l�I�vԙ:V�7�۹#%�u�Vq�s7,F�R��2��Q�4�2��rel����"[��]K��o���EE:��c�ޛ�$ㆴ��)�nI�<SO�Y�_� /�#�� j1��Tv]
hd��y:+�����JS�Ts�)����^�fl�ہ�W3vM�<ӽ��Y����΀S�.��R8�اE7m��&����K�Ot93�W���U�TX�U4l�IU3�S��ijw�O^��)Ι��>��N��vb�ɭ�p���ǌ�k�k�:vY�l�(מ_By�l���TD�<�Bi�i��<��Ё[�E�睆=]��Hi;cE\��4ys�3�[-��j��h�!'^F�i�T@���/4��z ��I���1�ٓ�"��Q�7�����f�z[�����}��ö�!�|Y >�s�ј�`+U�=p�	��T������O���f%��0�j|�ݒE����q,ˣ�YP�)<������v�U=��U�����by�:��K^�ݻ��d26���@��j�8u3\�U���7yBD��n:�a�w���r�\4�M��g���
Nz��7O��L��2�u��ͺ~x��ov=�����N�r!D��1�q�Ȭ�Sn`O�?a��(V�z�������~��xIw(�#���x3����ѭ�}��;)�8�tS�F�]u�wnX.$�Qr;Y�Mj%*\���+�_;�V�����!Y���fu���W���	�FTG��
�p��µG�o'<��Q���*Yy�a�]��}��U�9Z�\�HfS�*�᮶
�gnՎ�����l��
��C����|d�*����߂����0R:`�~���~�,��0+�����dc���:'#��������(��;4���ˠt��!s����a�7t�!�8�|�<L�][�Yer�g���f��k�d��^Fs��ѣD)��:�x�eq�z{��Q"}�B<oA:�/�-�z�9�S�GC��]�_4�2�˼�"���q��:8[C�����9GYu�	ޡ����t�T���O)?E���`t�d�f�	z~������@ͼ��K%1��:A�����׮qx�j��6���=��z�
@�jQ8^Z��iŧ�.:��vۅ��V��oWi�ؚ֎S����rZ�]Co{6�GIH���q4t�PԡQq,��h�=�o��,� z�ܙ�I�9��w�.4<��\���[)u��m�gtu��)���@D�T\KS�� >g<M��{sRq8��2�=;
�U*4ry���=-�����3����jaF1�t�'1۞1�e��8��6�$����_����[����C�Et��tU5�	<_uRQ%�DF*�LZe�]���W��跕ޣ�Vf�K�{c��kmzTξ:�M�xN�ʈ6qMO;1��c�-�k�}���9��Թ��RM�R^��r��/!��Ʒ�t�JiK]�P;[e�.\(��}@��ڷ��ї�)���S,.�W;�S�Z�Օ���t�[����	���]���(<vΛ�39U͛y�ˍr/O1c�n}7D�����Oݯ5���a���N��Pڭ�#K/�N��T�,#���u$B��E��x�rE�OtءLeFٻ�̌�N��{E�:6�;S<��n�n�I�U��~�O�)n�b��@�b��1�1��� ��+%��<.�ku���nE�Ҧ�Zڣ=c{��N�[ƙf<�y�ϯ�l�U0&W`u�k�x��g���T�z�-�^z�Z�p�k�C�fӈ��l�,k��6�0��ޓ{2;��p1�����B�$����ɍg�����tU�͝��
u�"�[��9�zʲ^�f٘Bu��\@<o��:���T��q'r�
��q69��]���K�輸������e.��:[�De��*���dz�~���=������`���E���Yq���ބY�Zq|��P�j�Y�/��Z��f��k�����U�)n0���vtf'�v�6E�K�k�+�i��څ Tz�'
f�|�-i���1g8�j������J���nAto���u��7�*�L�,uڰAr���Ӽ:r�9f3u�����k­k�y���	���4���Tv��W3���h���~��,�K<Iپ^Yp��p]3��� ���Ӹ�*ػq�8�Q��tLU��rn�ݴ��1o��˂�Zג�}�t`ﺥG��Ǒ�����KJ��ן�3	V�4b��qՔ���\ř���ۙ�n5r���k�!y�V:�u���4S7m�Ѵݍ��z�c��{$	궲q�g�;j���I�V;��H���w-��8�=[';`���/�W@4�%��Vk��L�1��;�-��S	jy��K�Zr���Q�a��9������6!Kb���E���G:��Zp:�p�C�O�h	jy����;Fv��-����\s]����S;�-Y�'��͘m��n�a�
kvt��p�t��|�F�1�Z���ƍDZs��6�-5���B���x�M��2�<bzvYĳwG<�k����0,O�:���g>@Pg�����s}qp}
1�
�����{%)��U1
�<0�o�E�7��tf���X�Ma��q`l�Z���x���eF=Y�8KY}#�w�dpauH����U����ݷǪ������#8�d{5wE�g�����vQ�o8�_z ��\�^�ʊ�j�	�����Z5���Ǳ�ޞ[�3�#:k�i�\�\�]���љ�w�r�$w9Kd�]�ZPt+�*<��j�Ժ7����<���D�2��1�$G��WI��<��j삫\͓0Ɔl��o�â���?�?#wM@ӢK�g���������в�k(~uu�R6�*̀�p��̡h����Z�6�y����l ���
.>�?#z���w�=��>�9π�\ %�gkmCnb���Bmq���9����sŘ�Q!�:���x�5o�-�L��XP���=�-Aq�[aT��zr1�K��0�D	eO�F^�'��b��,�l�Y�~qGe�K7�8�ƣ��ry�5
�F�qW̔���_8�͑��P�y��vM�(\��%�\>|��T�C8֋�6��fV�Q=C�G8�)�i����a��c��΀6��/��-n]��lc'�S9)��L���v��س$��Ȑw#�@�J��}N�����ڞ��������=�Ar&2�����Z�ĩQsZ'Z�SG^.�+��� B%K��#f���TE҆S�����W8}����=a�uZ�Zq����3����1ź����R�y٣!a��yh9�s����p��m�U�A��s2y�Y��4N'�9M�_tt�A:��.y<�ò�ffd�hk�҅Y�Hq�w�ן�8���*�BSH67�H��2O�]��p,#Wv���G��{Ks|<};.�E�S�|zH�tĮ�`��M�9�<z�X�+,��'���r4x�t)S
vU�=n�ᘘ:�"2>�qm����m�k��7�%k[�X�j=��{��S�U|̥��:i�
��Z�*��q�Z�zlSs�N)�O<����ڶS�7]y[Qo��~�k��n���D�4��Pˌ�;,{�Dq�q(��WT���!m3z���.�.qA�w� �@X;�������L#��
N�d7K�F�`��/�M�Ii�ޭ�M�Q�z��W2�F�;N1��:�
xQn`kR~Ô
d6�7=) �#���׽ kS�W���99G�v�zc��>��d�Fw7����c�f��:ÿ����ג�B�xC78�hf��y�^uR����7.�M�l�u���دVg�3�
kG�QbK_��]mJ ���!�1�[]�"\s���Ɗ��>Ρ7��{��gV'c]	`�1�Ɂ�TNMC_]�Y���q��c���<E�re��i���b�fkU��U�kȩ��	_���� �dzD��e��^������aY�byDJPצ�s�A�N؞Xx�;�i���Z�~2��f��=ڈ�Q�Q8^|��|�-iŧ�.:�إ�Lv)O,n��-�ީ�=1�`��{K %���׈��&�t����-���Ի��^�A�%sZ�5� ��Fn;��8\�ݳ����L�Ӱ0��4yQ�ȸ�l;Λ�j�����>s�YW@#@X|�N}�n���^y�̎]���~�k��R,1�ݗ�o�fe�}��?g�kE����+{%#O��GH�Qq-�w�g���S�JL��x*�9E��j��c����[-���r�[{�gOH���"T*.6��g��37:g�jNN-��Z��'����Y8���Zr�B�1��k�R�L�D#.� �f6[@D��p�9<��9��6�T�-R��i���*8*�}�e?�Q��{�zxS�}=�p�1��]��w�&���BO�S��^K>uS	�<�w�vK^k*K6�n����4݁�c�=��	C�e=�T^\�h1JDs>F9��r2����SGD�l�4*��t<���^k2��#���{�H�)^�%��I��;��`��LB���x?q��ez.H��-���7`��۹�L��Z�"h��)�s��fw��aǎ>7'�
Y��X�*x� N�u�O���P�M+����+�~ٝ��y;95�z�Sq=#�Q���_L��}���a�U��g�4v�/ڬ�]AS��t&��)=���#��O6�'1�;eD�p��f�ss��>;;�x��#������B����=cE>2m��<ّ�W�q�7د�J����C7'~��`CVhLm���^��
��iL�:ct�m�$Pz��x.�񥽺�����9,��^I)VDj;5NN떤ǆ����.�(z�Vƻ��v�!����G|�EnĽ�;�X�2UL\�|uZͷ6�X��s�ɒ�:4�;.�󜰘��S�<\�f�D�v�(�u�}�8��1��|Cي�4]u\��vG�fgp{P�.$@��lYؓ$ .ţ���x\5�gw���4��T ��������n���	��<�����3_n�U�uŝ�2���]*��Y���-Skb�[�;�.�b`�iJf�I�S6)'��-���c���բ3��e�q��5p�����OK[BA�<��Y���C�I�)�]؆�K�%F� ��6kΗKG7wn\B@<w�H�.�3��è��Ѻx����'�M�U�k���u�������6�ֹu���{��Ђ+<��(�ߒz
�ɰ��g3b�U�:޽[��y؝�/�VW�����K�^�<��ڙ0
ɂ�-E< ]˦�����4�7�����ٽ2�@_R]´�����_.z�*���Z68=N�!_#�������5!�g���Y�g:�l�9�%f����5Vͷ!43��u���3|�{D�59�1,�nj8�"�hp7�{u�Z���ג��{�xS=f�mc�Z�1�a��կX4��/&�Ss}�Ի����ںm+���f��U37@1ÍV���}�KyyhTZVW_Q��;���,W:��({�����5i"�WarK��6�5w�]Z6B���Y������*�ٻ��&����Jض��׌Ez�9�k x�2�T6�e�@���+�?��ط6�֞++��3�(z�������{�s�Φ�&\q/}5�uwH�z��n�J坎B�'|%���Ӽu*[���n�� �`����.m��v���!�x(]yv�"��&��6�y5
Z��7�N�� �H[�7�r�� ��yi����{���y���AIb�]�[��>"r��Y���]k���Z��t��3�Ԧ��̱h
�j��v�r�ܳ�Ǌ\�];��tqޮ��0&��UeL�v��i�8^�+\F"�$�qu�*9u9Z��`y�V�e�wBnt"��V��2�bbe����s�;d%�ӘhYWB��Ҋ#u�Ҏ{	����:/�� S�x�V���&̑����dӚ�%��3p\�5�Y�e]�n�e�J�9���\*�=YF����n]�tJ\�>�ҝv�xԂ��\�Ƚ�S��7�q��\�e��f��W �j9A��9��܋� ��C��4-7bP��h?��D]}S!63Z�Uh[�������"�����l���Z؎�Y��/n�d�e��:�i�gjR�)C�+o��r���;Vyv����85�G������ηO<cs�^�ˑ/N�[O�����pZr6,�Aޡl����'l�mef��� X-B�lrp�t{���]�����v���n��n�T��"�w`�9����\��"�]̬%�UXY	�]!ɹ�wb�I$� ]R������$9ؑ@J�UUT�hTAWf��r#�(umÎy��
�)!��k�8dRAy�
r�H9]�S

�yӹ�r)! �W() w@���(u8Y�Q����eP^w;�NBA@eȇ$�r(���
�u�PD\
��˲��G���#�'HЦ$R!�N�!V�`�EhJ�*JQD.�� �'9l��(�	%��))Ĕ�!&z��
)ȺE$�T�'Kw,���8;����EXE��� ����$��1��\��oJ l�F�ތ�Q���~N�>�r����N��Xx�d�K��Z�q9Y���lj:��D3��F�lq�W�]�r�����I�ڷ��n�+q�E֟�Ju����vПn�? O���<�1�~��f�؛���������fY���<�,����(qw���|�������v ��,E�<#og
��$�=N�UD�[P�`��~��uq��ބY�Zq|��(�{M�i���v<O��w�wD]'aL�з��]�M�eŖ�+�O'4Rֈ�P��8xS]>Iն���s��vO=JU�)�q�F'"뛡 5C�t���בwj��+�?=�;Q�&q�a�o�]�7QS7�/���q����V��!�>Ή�a�h[=��dpбѳ�����q�����fMV�f��i\�[@������N�7�c�����w.T��|��cM��(��Tu���ծ�P�e�t��@,z�zyU0�y���\%ϐY-lS�g�W��7tB��+�����ڷk1�>��ځL�x�A�ղ�h��� ���<Z�#��Xo��8�~8�}��4�Uǋ���DC�ū��k�=���tt7g��t*ݝ#g\x�0._!Q�FThy��q�.ֺs���u*u�Y�	��^p9L�f�)m%�C��-j��7[�%z�X���[=�;u�2E��*������.}i4��m����YqA(����*��I{�!�c�Ʌ��7��tT]6��M�U���x���JÃ7���[��Х����0�Z��i�
��S���Y%�%nݰ={������I�5\�F>aB|����`�2S�)��b!T'���<�+�,I��=��z�uzesN�������=bu�,��p~�odҎ	��a��@%"v���+��z�U=W�����n�f#Q�f��k$�����bUm����`��gmlwUjxiv�u�V�k%���T��aAy����/���:�S5����)h���u�{~�P̘��6�n�2����jg�[	p�� ��[�g��g���[���f����s�.��[D�a�TLS+ޣ<����nƶC6�s��7s���WTs��2��4ܿd�]5�V:�kmX�J�:�dc=��1�! ���Q�^�'��"��mʬ�a�?8��C��=%��8��ٚ�9�D	�2y�NK+��8����G .��x��~»^EA��6"1E��h��i)ʿ�/b=����.��_�U�;�<�L5�;��Q�]B�����^W��-��l�[�ݑ�����=�|ftUN]E�?z�~ti�Iśl��)o�{{I���2���s#�63z�\���M���6��{K�����6bNX5y���p�3��c+�		�L���I��N�#�T��ັ�&��8���캊�u�_&7���z�e�_�mӔUS���E�k��@G�*�y�{N���ڟ	m�U��i��=)yڱ�)���)�#���v���������:�A=z6hi�TD�Δ%��i�k���;='r�cs�k��<v��$Er��6���El�PڇE�����J YM4� VP��-�ט�f�ܙ׾�/������-}��;.r+[�z����p����"/*tÓP����9
�� MK�/4���5�����ʼݒE���.%ts�+�c�[����	�ABV���m��3-�ѯ�:��14��)�q���e>���<,d��;)�!A����/6��R��4�P�A��E�]6*��{��]nܙ�#N�f������U�ʥ�U���zS�f~P�]RD*��"[bZGC���"ᦔۘK�P(ST�<Kk[�ܾM���;�#����G0�a�R��� G��C�t*��fF9A((�N��*��ǫǞ���.�	��:8�s��v0U,6�#����Y����g�W`=��ג��EG-ҡM�t�u3���ɽn��]l�[n��q�����H�����E������Z��/D��N��ٲP2)���=��&k�ܓ7�@3wn��z6LtO��O�%�ѡ]Sj��{���\��R�K���L�t�!�1�y{Zj܅0Z��jlO��\p��I(�W��ys��9�"1u����ec��[o�<��O�ߤ��-Y���SM3=��*f���-g���B >�G	mw�"w!��/Pc�i��ʘ=���j�أC>rJ�:6u��9�YT�t�7S[�[͔��aL.=� o<��K�����e�U�׎��VDŉ�qxy���`����P��(�/4�|�>����#�csG"�j�r��>�m�ņ�\Û_/��:�zn�l�ۓ�U����?\X;M Tz�*.(�DG)�+=&g���z�H���H�j�A�?.}��l�]'Kl�kL�DiO����@��ڍWbɖ�M:���@������Z��oW�$$gȊ셧.T!��S���
�tN�gE��'��\V��B�*S��0�ͩ}R���ӭ���n��Q�m�!ѽ<��@v�\��V�����s"�S�p�Z��G�S	�<�w��d�没��F�+#M������ޝ��^���2���Lz�AMd����>���� ^:�`�:Z��^Z�!�Su=K�pQag�T4�M�}Wn��έ�
v���N�9g`.$�P�ړS��Ԋ�j�</�N�Ha����T�]]�Uޘ5�TF��Ǘܜ�\�2Ex�Y�v�O��$��W�Z������NG�%�~\��f���k,�b�o�?�Xt0�ve�$\�T݀N
����a�o���s!TB����~FM�б����M��*6�����A��r�2��~�=��l�}v��q�'�t��*�r��Џ����T����R- d���ΨT5��<�t3+��T6��=��|y���>���T�*�xalϰ;]ݦ��1<W\���;;{}��/9��m�t�T[���z'͐��pP�n�<�n oA؁�h�@���0����K�p�Jс[�� Y��w��o~�����9eY/nˎ�:��2� ���e��<�s�N-��|����H��!ä㊳���G0�˾��x��VOSvTɄ\�UT��z�!������۾�]Q"�j�Y�g�}>~��v�8{m�E�����[VD�c��^��V^��z��ծ���������;*L��A�ο8�{P�
�������R�O\<	޼���C^;$�s�}9:�#���x=)�«��C:�d�hU���ݓ���n�}�3�c���v�a-�q�N���s��9��tH�m[<��GY���CE{��hӹb����Y�+S��W`s����u�V�8L0�F��(�u3w1��ml�إᒀIѦ�뢺��U�ޮ����0����d��]�rz\͔����9���$�R��vi���ò�W7'=n�dY{��N��QҼ�-��U��՛�e�/g5�.�����IL��5�e�߆��tb���<"G�_��vr����`������±^���OM�zyU0�Tƣ@����%�)�;E�U��=5"�s,�+Z\�Z3'�>�Q]<)��:9V�&O(e3F�
�>)�%��t�z)�)���cMV-m��s��y�u��m�����U��l9����b�s�遲ϐ���}X!˼iI��Dec�	��6M��Ptu�Y��a�,�χ^|�܎�i�T�?<2j��5�>��R�S��[����Y��NY�}��$�OL4.oc�%��c��Q�)�!�uOE0ֺ̼~��n.;l^�������q��~�-n�=��@�5LYI�g�oe����N� 7ս�̹i�W1*�/:·��<�$gP�Fq���/��蹆���%Q��쳜�2�o�Ge�]���:� *f03+~r���a��h�V����Y.l!�;u����⫘�j�� ��פ�v�L�v�p�R�_�L\O���9O?������_��x/�1(|lW��v\SN�[+�(�R�sa�(�oJ�.�;��������~��K)��Bb u9s3/��֢˄�H�Xjv�>�Ů��+[���y�ٵMr�e׏o��p��>�\�ZV�O���df���#��>��[c"���V$�<��
������%��㟞{���ҷ���	�~��6���:�x9�z^9���Ogׯ�[#�vׄ@Η�+]�o"��O!lы��.c�2��Wsq�)	2���XѬ�����l����r8q�P�y�����b��*����izY7)����j��'i�M�3�S��)�Z��}e0�e�߅�g@������Cո)ޟT=�Vt��Ω�ÐZy�b��ۃ�z�
*��,X:����g�m;cS�j8JT��Db�8I7W��m���;�^���W��v����� B3�U'�F�Ш���(F� nd��w�ެ뚃��Wzz(%O���t�m��<���v
-���&J�ݔ���M�}�m\{�v����H�]qy��vZ�G#�_F����r+;���S���5�	9cw<�b#B�[zpTf�%6�aߵ�ۨq#��T�P{K��Tf%�tב��z��Ӳ��@˶��F�n�:�c�4�Nq<�����M�.r:����2���e,�qȎ6oQ͹ˮ��~��p��Ӫ!����Q)���f_-_gZ��E#n7����N���
�0�~!��qz���yP>��t��!ݘ�|�d�umt�L1e�<��q��փ��{�mAW.�r��)@N��\J'�H8;�r��ս�<g�uj}(~��|���eQ
������9M\utت`k���
L�n=�w�,p�ұ/n��ӆU#�_Qw3��l2�;�j ��|zcx��A4����O�q���˪�b��Zsg�WN�n��q�Ѯ���7�__�t�� �?9ٟY�L��E�o�4���AQ�r�^V�+&��0E�s�tls6B���f��i�s��N\t_�rX��O'��n����z�Uk�6<۝�e�����'�^=p��l�p�w(�W秺 _*�Dǡ��b{n5���ʪ�XThs����ѻ�Ty���ӽ���|� ����"w%�u��Dz7��`~��R��rz�����[P�l�h㬂*k�)��ufZ���&��{��Y�󴧯n�YصWr9�f���v�`�k��<��'�ȭ~�'iD�yf�{�i���v����<)Wf�X�8�
��7\v�=i�fSv˝:���Mr:@إ
����d6cc[4��U7��zFk�*=�����מl�#V�,�9s�(���]r�[k���t�x��uА>��7uT�x��U����U&�Ab��XUy�u�?j�t���jz��T�&e#Z��]2� �;L��s^k����/.Ś;Y������au��Sŕ��<z�I��S����֭���g��|73�I��k�L�W�=��'V����Zȸ��͍͗�n��.&��f�~Ց!#-��U�u��ء����}�:�����]�_r����-�������0��L��$	�}Fi���%�,O�u�?��B�̶�;�Y��UM��v�I�i�/=";Π������ǟ@X��(�au0�����ךʆS��Z$Aiˉ�c^�n��з��M��`����q�ʟA�!#LX�n}6[!M
����Oݯ�0r�j<�.-B�P�h��V��6s>�i�=��VO=0BU����`�W�rE��M��V�2�qc�>u�<b�+��fF�;�k���q�<��b��& �,��i�=4v���-�UEƞ}�ו3qO�`�e9r�f��9L
���_N���/��l�uSU<��n�`������oH����Cb�gɷ-�Wr\�Y�=�,ClB��������@�4�;M�}���֢�Nk�� �N�q3d�����oMw,���9ͅd���.0ͳ0����53Z.�ڀ�rY7Z�/�2V;��Q#�p��P8�4��)�()��ǟY\K�k(�0+xl�S*�qbX=�XׂT��J��(��wg�"�]ݵgAU��s��y�eB�*�#V�2�jׇIWzN�_PXL<�)�[�F���Q�'�
oێ���<OK���+qZxC�o3P���<k$�Tn�{�ۧ7p�1l)6�!ч�Gw����5�Ʀ�E�p��Si����wlОڇs�O1�X�����8:��E��e��|n-�����Х�c��a>����ݵ�-�th������(��B�+���.��C�����y[#d8W��S�k��[!�\�B ;j���v^~SC2��4�������л��w��3ۙd�a:�I�ه��|g���r�lΚJ����od��W"��J9Y�1�a�X�Y9���#���j=IU3��(��:��#y�����!\!���qJu��@��+&�{U��� B���d�UL(Ƨ�.��^��o{Q��:T����}ӵJ����`��Fy��1�*xW�T>���I�� YLѳ��MF4�v�S��Ʀ7�b>-��<\�0/;��;��ز;a4{���w��9B��p�GLj����P�3�x�*7�:9��pz)�{	>Gi�[ϥ<�zϰ�/�9嶅���fuUװ�Y��1u|�הq�`�}��eM't�1e��gD�ZB4��!�L�x�����6�6��0co� m�m������m�m���1�������`6�6���m�m���1���lcm����������1��`6�6���������pco��m�m��lcm�X���������(+$�k(%@�a��B �������'�����B��)T�J��@��UR���(�*J�	J@F�鰱����haM��J��[0���R�UM�����P���*"�T�E%*�**	$/f��T�	IR�!*�-
IEۀ ]�T%�`P*�ib�bjb��T��"D(��B��� 8�WJcL� �gB� V   ��  ��������
B@�\ �V�	���dheJ�jm����m�@(�Ֆٚ�ͪ��4$�a��,�� �� �IAța����M�6V�m�V�ն�����5�[b�,*�n�mjBنi�2P!%[�� m�45���ک����D�Yl�+6�ɦ͕��vs����P3��JQ$UI-�w6��elZ��S%�-ݥR�����F4�4M�@��(ԬF4Z ����Tj�VօZ�̔lă6�hY�AMbJ� �dJ�� и ۉJ��h&�([eR�)�1)D�V�L�$mmRʩU��� m�Dф��$�؉l� @*�̅[[ADT�P-U�)�� ������D�k(M4�4�6b��
���  L�b�$T �4i� )�IJT�L@�� �2a<M��b44L�L�  j��	R��2d���4 4�)M1	�#�=L�?T�F�6j�jA&�*R�6�h10`F ��q�f�ԟF�o���:ʗ�}�`N+u0�_8��-h >�K�`  �����Pp �5>d* �%���|�����@�>�� �5UT  ��?�� @� ��0�CH �W]�K*ԣN�S]�  ��q�1�;k?7�ٰ�R����߫�s=e������0�E�I7�xUY;��Kee�sL�*f�-$�Xe摗t��G(<
26�;���h��bY��N�0f�-���J�2̢N&��#�.�&�FZ�Ө�Z:����4�{uv".=��e�-�q��+L�X�o+�a���d́�*�����|˛Q,��>)�$��i��P�f��I��j����P9vP�nV-p��5T��om���I�ƃ��S׵ZQ��1�7��^�L�f��3�-�@7�[�6�!+ZR�S�L�t������b���&�"��813y�hH�+4�
o�{2���Q�.��ɍN� ��z�ءv�x�y(T��E�kJjKR���	Ѱ&�,�� �t(���Z�O�����]"� �0Q��R��1Q��*{r0�f��`a���rە�`۪�FHi^^)�X���"�v�<_bZꫳY@�SU�B�#Çsjn��vn#��o�2����v��Y����ZKKWY����-[�ԫ�Z�m(t
��i7gj��*�yu[������f��򑉷!&���RSI�SL$r�bYf3/䥊[6;bG!OoFӎ=�q��ʵ76�ڮ9�;�n���;B�0�B:f�t�̂�-/	��G�Ŝ�7b1���ܬWn���Υ)���ړ�Vpъ�hq�Û�(���ڛ+r�el�
�MV**��̺��@�Ҳ��z�嬧��5�&�b1���26�
���%uN��Sm`5���kr�{�[��鵔5�+6�����-�+q`��.����f�T�;SuV愘�UA,S*��[{�f%��䶱�^���曍��x�)R��T*�仰fG�-ڛ���ZҤ��Ef�yc��geV3kv��0$�T�3r�y�a����J��\x)J��U-�0-bl/j��1^�K�� ���eZ��U�mJR�Q�K	(iU-m�o�w��0�"�e���ȼ�+V�r��^c#iEWCN��f�U� H��y�Q�*����U�*F���
��T�5{+dsp���b��B�^w �ͨaut��+�FMp$��^e��SoD+e`����1%�3Mܴ�7oj�X���t�n:�GU���ˢN���J�n˻qBƼ�7��0ڈU,E�rDBeV�!��z�hn�V��xr�W>0�WA�ΙUsF+�Z�@�:�n�٦K�x#x�;ml�ٖ_I��;f��!2��/[�HĚA�EL��E��v�ӚC��de��gm<�nKێ-[5[�Jm⭙�^*�ͻMl����l���U����e�xu9Y�����J�ûe1	�P����űh&v�X���Ww:m��g:��֊=��1%7q���`Ǥ���[�ʪ5Q���]�YG �q�mQ�a�c�heYx�~�j��ު��;z���ի����]*�jk�i��wP�5ukQl�i�j[
�A���Ѱち*I������Ե��"Y�r<(щERzm�I,�X��kqL47d�,S�D�@NX�Z�!�I��W�ٵ�I�#5���2͝6�\���iK��t�����˒��H��cI����d�ň��'�J����:��Co�ÕU��X��wal�($֘�Z��ݣ�
�B�@��.hjJ��0�v�x�؅U{�,���ɦ�%E�EQ`k�[������$��IZ��&	�(���N
x`�&a�dV/>�CgT�����E�.�&e�����<��iX�R��k.�k��ǔ���2��3f��!��UЙ��0���q��6�3`��(�Z)g�"�,U�)�����Ǖ�H�S�7�C ����]�el�v1M��4�m[v^dN[��h�EssKOE]c��wM#rPG/d�`:��Ʒe�YJf�l7L{Dc��ۼ�]w���	V�>�*�v�B�u8�a��xX�*���˳q&0P�6ՄcSjT��u�ٰ�hu�+`����F��2L�wVv�X���y`�bP�*T�q,�b˽FX��FT�#��+6�&m�b��Ȭҳ����αF�N��9j:AkM��/\f�4=0f�6Q��id�!�����f�n����ì�nѸ3X�%���hjnM�w��.�\���6�YՎ,�(Ofd�b�ٙ�1�Z��٫�T��w%Ġ����s�����d �4-5,,I<���v%��d�v���&e*Ƽ�Fɺ5��I�T�5��h�i]��2�d5n�h(����)J�^�sM���)a���i���m��>GA�bE� };BSˎ�Ѭ��Q�b���ֈ9y5��V J�s4�zsj�5:(cV�b�F܈:U������n�	I�!o%�V������d�82eG�ْiDlв�E���F^=$�J"ZL�8��R�m�Ph��j;�mM��#/2����̵2�)�ywEmw  ڼ���aBZ6���2.G��Є�$*`�Z��є�/nļ�Á��SA:�dw'�-N��� ���;�^��#�����=Q��.�e�*��m�7Z��EZ�\�����U=�������ݻ7/@��ӓ0:1��Y��+r�H�4���QrU���:�Q!Kj҈2���)��`�/2�ې���*��k.1�S�'0�S��el����Cc
�M�]���["�Fkjb����
��M�HS؊V�gp��ndI4R�F���k48�#��죿miXKf�ъ��V���dq��n�n6X�a�p6�C�ɠ^�ێ��9�sS[�pnՊ@�L%Ve�&``
g[�����G��u�Rm]���nL9�3(�"��V7h�7jT��jvK:�^�uB�d2�S�JI�QKR��vڳ�su�X�[E)g�r�wR�7[HT��U��]+QX�f�Z��en��!.MeR	ŷB��`[��:��jQ�¤hd�7v\I&��u����b����:�*щ;��m�*��MG��
�t���dn5��Ј�*�H�q��;Ճ]��E��)�u	��4�mЩ���x �df[�W��3Snh�cP�j=̧�LO-���1���\���nj�wu�԰p�{K7��@��ڠ�+�3B� �!!�\��M�q�8�l6��d3[�Ӛ�����p�q"�1��;t������r�B��lb+I����*E��VQ���Y"�ϑ�uzY���Y�zP�LG5���U4+IL��wr2P�DAh�QF�!9�b,�x�Ȧ͠���[�UN5-6�S�(8��&P��(��̠c�q�����n�F6-+3.���1�O��%\ׅ]M��Ա�,j���J�3$����m(՗�����6l�tb��FP���+	�_fZ�p�VNn%F�����6��R��(r��1.��mQ.��gv��1�rk�ٸ#Cv��F���i9W�2�,K��OE0d�c2�����ڸ�)*vo&�;gl	��}Cm�i�j�r5�D��+	�)��ٻB��:N�r� i�y�#.�^�=���Ѯ��* �I4�]՝���V�:nä�E�1��T5�dF;�B�ZZ�Z9��4e[�z��:�юٛ��;HUZ�:�<��M֪��(h6�b/&�#��ɗ���H�p'kgM�1`���1��YC�`+-n�.k�T�T�)�V���U�he�j�w�s��w���?X?/o�?1�q;N	�L�31麨�~@��?"p?�t�O#��n��.W��z�����r��bfp!�Wo��Yd�ˊc��#�ݕct��ͦ����6������u�v�qp���"�Mg-���r��|tC�!T�3�m�Ih����&� {�->�ܩ^]vNo�;�Q�e��:޶�ce���)��ѻ�_R@S������p�$N�Ϊ�,�ޥy�V���u�ѵVkJ�9h��b�8��`{$˽� �rj�-� F㏙�q����q5yq�c|���ݠt�=]%M�E7�\�Mp�[{v-`v���֨o����GD!}�!}���:��ۄ�E�C�Ҩ����K�J"?����9t�mEz��s�ϟjW��(���rG��Z*�����
�v��g(C��+{%J�#�g�,��I,�VȠ�t�V9���ޗ�m���v��1�I�����]M�t#�ǻ�N�N�ʐ�ƕ�U��=�@�*{�mn;��7y��MNw��P����X0�|�t��j�˫e>y|%v�rq��T�<�;8S�'U��EfF� ���������`(��ǫt2�bc���h� ����u�F�����檽U�:,PFge���G$'s&�6�=���[�i��+�\nL���vJU��G+-��˶#���zGoN�}bV�[ۨxWwr��ͮ�Vi��!�����˻&Wؐ��C�����X�I�}t^2���9�Ub����1�� r�b�`�R���]��#��&h�Y���>� r��f���hĖZSE�"m�1&����()�����.��].��������-WB�ա+��w�u*��u̪�����Q�Nx�2��̥+R��t;A�]ž���a�N͕B����F��2e��sI��C�m����EQI&"�O"�,����M���>X�+x_�j��YʂZ��l�c�ẵO�=N%��;]	����<�ͧ���e��n��8�*��Bz6�w,��f{W��̘N�i�(�^��`7V� !g����Y���]�S���,�N�(s���|s��MA�q�XI���\}.u= �G���x�eޅ[(dG2�r0�E�{�9�TخE����ڻ-aڼ��r-V$�q��j�L/�*`�
�)8�N��	YÅ$�����a���%Ǳ�g+u������T�؞�N҆��c����G���]����I�}��\���	�Y(E�R�D��!��-��wuҬ�F���R� \�����(=5�;/�x����*�0�$kh ַU��\�]+�^�;[`\�=���\y��d��\X`JW��hZ�Ӭ�S�X�֮bl�b���
m¥�7J8R���J�F��`�՛t9�E�7�af��ᝈT��N vV��N4�V�S���<�.)�&�1j�λz�Y��	ua�ٙ��G�Q���K���W�"���+ =l�+^\+���8P�1:ru�uy��K���p�Q����yM��-b�vf�N����Ǽ�	�B��+,&����j�M�[�T�͖�N�i����;_a�������D���]�J�g*�UF�-��u��p��⳹`U��cm�m:u��S�����\�j��pk���ܮ�U�>�*M��,niz���������:��������*�m�&��ݝ�y�҆���s�a�Gѣ�hN	�[=J��L6]�Y[�_.�#�374�W�r�9�草���Rj�e����GÐ�tteE��� VX�V�ѩj��ܝ�SvPf=D��܅վ�U)av�J_9��u���e�X���A�Yo�De��PR���<��S�^�W7E��3��so;�c�Aԗ8�lwE�&��:�'t���O�X�wm2�9�*eZ��L���I�uI��BuR�Y���q\�ہU��`��mE&�U�VO3W}��j}Ԯt�x�C�[tY2�;�͊�km�vh��.�C�^��U�Δؑu\�wWS�k��.��L�J�tj��S�r��#��	��NZÏ��׌����9w G2�0�n���+����Q��$�@�j�@�!|B̦{����8y��*ɮ�6l.����g&��{�A�&����t!��Ŋ��9Ų�@]O�ǽ�7)�y����h�]����r��oq��:Ò��#cmm�ԫ��e_P�[Oq�)S�2��!T�:�TRxI����<�$�بW�"�?�:W��b�G�/ ��bǯ�9%Ƶ�J���"��b��X7�5'�Y4�!�Q>����������U磮��m����Ŷ!�u�`v�j�5"��yT^�-�>�m��;��*�W�N�cG-�v��
pɹtz�T��q�t�wn���fi�J0�Y:�=R��Z�������U!O6��!J����r�n�A}�jt)�|�N��5ʛ��%�\�*�:�t鷰�df���h�(�z{�hU^;�$����Bڮ����H"0E�^��I[�ffǖ�cd��QCj�K��l�k,��ָ������m^J��p�Q�#�yU�7TH�uJmImv;�ekG��<�R��͕`��Ʊ+�,��Sw�9EӢ�uη�2����B\�O-�s#�V�`�8�a�R�0���f��FbH���5�9)�A�j��yZj�8Y(�N�yԴ�Pn�3y\�W��V�t��;K�'![}�J=۹W!�L�m�ݫ�gm�̴&ĕ��o�xaib�*}��]t�N�^b��6�P��-{-�z�6��9�0�f
�B��Q­ܐ�S����C�]Vr��ϟvF⬜�j�<%��#���l<���̈�^��q�_��sݲ��MJ`�Cw!/�{���)���U��C�6��@s�G��Z��S�E���8*Q>����sm8�윳:�CD�������"�,�ܾ�;ST+u�7�����޽��y�d�;Xd(��O{��ɰ�V\cP���ŋv
{��f�
f����{�/8���	.��+��S6L�p�e�ڙ:���#.궣O�*\7MqF��*�H�ޣ�/�"/��&&�度%����Ĳ�lr���dY�'�v�)}���z�hiݙ�bJG,����[`���pd��ͥvu��K��Fݾ�Jk�U��nKw�d�v�ZVƳ��I.u�8�Aq��V1cܒq��&ㆲ�M�Mw�������RŒOWC�(7؞�J��tj�d�2�n94K
۽�ؐ�ÍEs\��e�sv��ǶVGv��@w_B��C9�g6�PҮ1,[�F�����3/�*�S��q��L �Y�ٻw�{A��c{�c�Ț�U+#�Z,W+n�T�I�U(e	mY}��^��r�⡢f�~~َԤ؞3����k�	CHk�ڤ�}�,�-K0oaw���;:JH��SܴΉ7�#vi2\�
�a����� }�S�r�f��Y%N��|n���4M���yW��s���8�!sOV^��dN�ͤ����jX{�m�䶭Ѭ�4��Y4��.�G�&`�:�-����^�v�wT�Jm���I$��IM��ޒy��gu6��I$��IM����$��RI)�қ}���I%7Ҭ[��T�y.���t�ô�*fw�_nvMM�F��'���j +i%UY<R��Z�IuG�<�i�}��d�r�W5���2�Q���qCW�l����,�Qs(R	Qr!8�eV9���ݚaj�2���d��� #��N����Z�D���_1 q�Cy�իtKv�ZU���lyV`�y���Pb�1b��q>�ՠUc]WZ�Z�U�$W�	n�����P(�&��2fIJ�;��1��}
C;t+| �WxyIO��3v���n�d�X\��q�o\��oN�q�Cq��1���=��Q�s��:0`�4����8�yv��J�tұ?L������j��$����x8�`&��-P���λ�����u@��p}�<%�������Һ��l�v�iq�;��;N�05�mG�E"dO��ܺ�����m]�`��K;F
� �Ǡ���
�A�_P�"-V�bT��en�
�K�����R�Vb���R�H��8r�ڛɑ�ƚ�v�6�r+�v�=��_�V��(	5]ں*ɹ�{!�bi|���uV.��ef�bh������ȍ-��g�ɸ��7[+��U�j��K-u��sT���M��jtT����S�F�wqO�ql��ۂ�ѠZ9�s��慝U]��F'��4���p[Bh��#WW$ڒ�DYz)d};y]S��Ek���g�G�����yj����&q��uwF��'�E�sk�9Uy���D_P�<�_f>-���=Ic�8�t��˫[e�חײWb�Z�F��koʾҟ���V+�rj9���P|�+{���Lж�w,���]TZw�vf��Ќh�5�uɼ��Ŝ�"�d�ow9wt���]F����\~F�F�f�7f��uq��,���H:ލ�`u��8�3�ɒ`ox�s��8�Ť�%R69X��*��r��v��ʬ��dD,�*!\Qa��@�0�'qDS�u�;���-��N	��_V0�8�v�n�_I���t9�U�L��~(�ܷ�ښ3�B�����j�{�����,����j�d��Q,��t&��V��jۈ�R�w�^�����.s�.���㪖���$h���;,����r�)�#�/��O�t�M�a퓛GlGh$`/��S-�_=��wh"�w]+���{�w+5�8�	�u@J��v�`���u
�q�Ӑwk0I��t�Iyn)U�nӮ�ɯs��Y�ѷʕe6�����\���2�a+�՘5ʎ���pf�;�����ؙw��n�9in�sVh�,S]t�Ӆ��2�8�'�&�V�,���1n��²a����^�=�*O6�d�ara��u�A�u��D57�)ZH�Of��\��SW���鮾;�;O�G�� K���3Ntw�,͏�u�e�GkjV73U!Uմ꺨�%=4&B0<UA��Ux�է�ky���x�� k�wn-�b��Z/�vV.�+{d��Q�u�'�7��c*Xȥ�W������:tv��J�n�5��w܃���WN��j��yӡW��^�Me=<�CD�:?evtB-�w���p\V8c��$��ʺ
�4��RP4�f6o�����x�ь��µ�FB�M4���3�r����v@��MO�\�!��1L¯ncn���6YoM��o]���z�:�Q��
q��� �[C�7/�.+�%��So;'iU�z�ȥ\(���&��2��c�Hbe�2`,c޲�N���;|��u˙Ӳf�WY�}{|��:�R��c�}��@ ���&�P�A��.�R�;5d��X�ҭ���Jʉ��U�]�N��8r��觽�ɥ�)��u-�4�Q�k5��t[*��ݒ{L	%�r-�9\�+�m�}Qf�9?�ZXUz���$���x��O~�A�=���eB%n6P���Z����vVu�wS����Kי%�(�y/�r�����+2n���T͕��5���o��3��
���Ŧ��Y�Lz�7V��3y�5e�b�l][��{�N-ޢH��y�Nl�
w�UˣT*��n-�`��q�Xy�
�j�n�Uj���q��ܑ����J��Κ���k���UT�f-��;�\�3�ᵅ�J�w'�R��9��jj#)vb�,�ۺ�/X�$��&�q�4�X:��E�*�Ww?��c+�M>�غW��h*pT��ّ+���u�|�bet��8�,��}��]�Y{JMf������<gЬ��3��v�*��3X�:�#�6�.A��(v�}B.�����WO�G��tAB��W+:��e�r��8�.9\F�K�:l�ǑJ�e�"��謍��^����E(U���Bޱz�]�p��w�&�>"G�:	ҋݴ��Ըoq�0v�{ϓ��Z'n�Ps#���ǆ�\Mս�����Q���+��Ő��3'T�p8��o�ыMv�H�'BY���c��:�b �l�@��|8��|y��|+(#��d�Ca�篭]�H��/T����ᓙ�m��=Ο\2u[�{F�������i��T��5�uf�IB0)(��8�S�}��t���=N�V��2n˥kYto�%$A��n�%U�z�r�ϵ�U\��\N
����h�u��������:�_'��:��@�T�<�����;�	D�gZ�93�@�7��<��-S�Y����5�l=N=��d�r�v�kκ�RA�������]�º&(� ����TK+��L�O��mm�wO������s��b��9��m�M[�Yyo#��%�ZE��ʈ�{q��IWBEf����]7P��Wu^��V![è�{l�N�=���WU��&��L��_9"H.l���4�����昽*��y��"A�Ky��e�ޒ��r�Yy���&MeCc���'i��6T�(<zE�J�Zq��2]�+�j�ivs��@Y���`T޻����w(D�gqvH/Wi
�	�����ҟ5�M��c�PY�B�v:�M���b��E�\̮�A���S"�.�Q�UK+��
Z6x�8���T꫋Q�HMRT.���l�r��f�Bl�
�
������xTd��B��o��Wo6e@�Sq�J��1�Ql<���]P;7ϲ�Yj�㗔����m�Ħ[��T��N|����BT�����w+�M����SӦ��_V�O+t�������Ճ6�8Ǔ6���J&�p��D�q��
}��IU#�Qpe
�h�_�C�b�-[VN�nG,r�9nh|vэku��s�HWs�5n]��N��\Ddr�X&7��hJއSs&���&[�y�49s��e���G��|v���;p�|5j��������B*Et�9u�d�����h�_:���yJ��m��+)��%��:+�jD�z�oR�\�S{Z�*tY����U�ǣN�H%��sjp���.ә����}�x]%H���Qt��_���^a�n�Au��S�!�V̫��uz�A��fG:W4n�ҏ���j����(f.��S/�Fh=b ��Zm8��o��%�SCSά]��.��{*e�g��Ou/��#c��J�GL��O�ępZ�N.w<ѷw^�	eh���]n(ԇ��̮�j�V(gM\(*�?x��>���zjzn�vY����-<���u��C��L0ڴ;��Z�S�h�R��.��]8��:�+�=8]������%q���Ff9c��m)�N����F���gv����l�<�V�/Rn<Pi�ƕ�č��w�WP�ʊWwIU�o�
���;�m���뷸c���-�HU� �Ǝ����{��c�F^3gvgs��CKNg";������y����y��۽=�	�I$ `���2A��ߕ3�����3e_�)��RMU�ǝ���u���V�e��YW�2T��6�+�����Մ��j�!�i��)��t����=�m2���^,��r��[�(c�_O�Ǖ|$�F�e�{;�k,�"��:_H�4�Eu�Y@�]�H=T�M��u���Ye�t� ����K-.ZY7U��.t��ư��4s�A9n����eQ���9�� ٦��\�.P̱B��ِ��C���Gnl�A�������7Ժ�VȊ�M�m7�]Z��"����k��]*�UCm��m�KYt7n���ʘJ=%�*���h<��b;�Cx.�"/���Z�N��ïrl����K�f(���U�b���v�/���z)����׷`�O*�w�7�P%�p��%�f9�+���6���;�����`޽[��Հf��@bRAjH�$�oK�z�WSξ��$���7�?�%$I�mb��6���UTekhfX�E�[j�E;J�Gv���Tul�z�5�qň�6�(��,�Җ��E,c�dR(��.uI\T�b���f2��`��U�1��lJhcr����\m-*����dU�)��
�Z�MeV��*��YQB��a�f\2���B��[+t%�噔�f��8�Lj��-E1̠娛y�I��r�1��DF�ԫ%j*���!X�s)��V��[UUS�&i�X�o�q2.�aU�j���kKr܈��X�(�	��������Ok��Ww�𜨇��c�f�َ�7�3����eG�Z���~;�S��w�����:~�P,|��vY#��ȉ�/��.0cN2�b�"��g2G�P�ޥa�e�w�q�]!��׬�VNI�[��n	�z �UV��dz�q�\K)�ԍ-5��D��v�f	Ks6i���J{�._(�J��� �A��xR�3G|v��L�}�:���q��R(:U3C�PL1�Q�B���x�(+��9x$����tJ��g�k��U�9q
�-����Nɮg��NMr�5�4mb�.���Z�9#�Cǡ����|v�Mn���֊8��$,�G%K�藬[���ӏc#љ�����P{oF{7�5n�dI�`���R{{-o6�
�da�v�s[�o�p��\wN���Y)����L%N�^��+�v=X�iu}:�-MOhR�G���q�|�1W\�_"��y�!EՌ�n�����g��}l�W�:jTIN�Jd����!nC�;N�g-Vݎae�痖�T"vq|�WQ��TO>�}&��Z��ղǘ��q���-�-9�.:e�з��Ő���1�x�o+��:��5W�qMUD��خb����� ���)'c�eR�����q��z��+!���-��P��g\�^���Kk���W(����#u2��π�a�RL���i���e.\��.u;Uom��bogu�nrR�%C�c]uw����-�h���g8��;M$O�f��>��*�X�)�4X�t��:��h�x�)����A<Śl>� oJ���񀢉s�j0T�Ȑ��ك�0�D�c|�h%1>Ut#Q���w�Us+V�/��#7�Z�.�;f�gy_{w���:�s����z(b�Lp��~zJ��zy�#ږ����{��k�*7�g+�)ŢI({]5}s�þ�]\����ڎ�v1��ߪ[�{s�a~�G���Ԧv����=�u���"^���ۚ
���;y�;`��y��e�����̷lV@�k{6�+�SkRݭ <�z�"�b{���ѩ����c��pbm%yO(�4�x�.!�ɻ�w^l��in�̥���b_X9���c3��p�[���n�f��2��+3��.�>�����N���rv�����`q�� ^*�ݨ�%ZVol��T�\I��=KC���<
N����R�缺f���6�#����s��z�h���b\s���i>��׌~�@xyLLGNg�]��Ǟ�8
�n��5�*�Q}v_=8Ŕϵ�<"'"`v�w���oڜ��r�y��Czw�]aY����":�H9e2;	��և�[ۜ�
d�_Am27�e�:.�l�s+�B��ҺC �~x�{�zo\��8�T�8�s�N4`�M���EP��ǎ�gW5ܭc���#�Emrn��\77�T#|SLx���3w++/�����U]Gw���F�	��V�,ꨚbC���B���aEM���M�6$��>쿠�G�N��Wx뽮�*4��of����=�N���^؀T�	�gz&14��8�����{z$㷛�z�;9\Q�ޔy
V��>6ov;��uU>4R��|\�[,Q���c@m�nϝ�f'G��syx�ǽ׎��������|�1�Q�1ۏ�"�<��{*^d��AnH��v���S�����n�u��D�����n�ξسCH�er4&��Xiɕn�d��p�7|�yWW�<t���74Y��cnV�כivs����;{"��G����Yt�i�d�oe��-��7u�s����`�7݂�.�u`n��˥9�	3ˇ��&�����
�a���Q����s��s�l�{
���;�����f�%����}P�;�[�^Y��Z玔���Y6�y�:�gp�2�1�S��͉U��=KpFÃ���wj+�`g�fג�x:�,bb�?��w'V21����܆�9�ޙvi^�]�AS�}�]�a��Ƒ��rh��\��l�6e��{@^B�V=0���n�H�c�QC)��~�,��ۄ+w~=��k�ܗ]o���y�p\��t�!�/�K���ҷ9��X�7'�H�\�0xQzcP'�;p\b�������m�E]FD�UwIgeMZ�W�[d���)��ڗ^���Vxc�����T/�^n%�'l���w&�����c�g�F��Of���6���=5y{��T��&cZ�w��A��6|��]F�tH<D!��tw=q�UrW�^J�{vm�I��݇�j���r�w"Zi� n�^��}T;�2	��_)BȊ���� YYi�+z���E�|')�d�:���zT��n��tQ=��W�f����#����f��[��y6t�Y�y"�xi�}|��k59�GeV�����6ˋbPx�s�q���/���v�u��������I���ӳY���33n�<�~�A����]U���K�����^@Ǵ�F�P�f7G����������� �G�����h�v�~�Ȓk���>z{ʝ �V��~��!�x�2�կ�[�w`#��m�3hfW���T���=�s(Gu�\�eHɜw0Uڲ����wAۙyhR㨣����C��H$��b����w�aE�&�m�^w�#�y���r�U�ҷޛ{É��J�����K�䜽\V�ا��B��L
�V�Fn���Q]vB�3����a���[���/�q�U|���f�U��7�ׂ����BM������ ΋w�X�.Km��U��AV�:�-������ q웄.����{�r8	�ݘ��}����	����ݻB���b�:���nv����7�Ͳ����W��b5ZϱQc��{�>���qg���,i��?\~�LP��}��h����h������Uh��Ws����1"�UVh��8s�l1��CM��M��Nj��1nX�e��k���Ҳ�$��.���C8�����
�"����յ�r�T�T;�ӑ��5�5W�/�v!U�J����\xR�V��b.���!Y4����-ޣV[e8�fN�����n�;,���t���ٷӪҷ}.#��K۲ّ�b��*�U`1Ra�{�=�ӷ1�h��Iʂ��w]��/����绫���w��_[uj������,�t�RuP)Rknr�/kKMM�k�9m��z��SuP����ɜRe�x��J�HvGA����ѝk� �3����pp��B�6�m�Bc#2�rS�'fT|cpL�y�GE��5%��N��5�����?:�[���*{�,\F�����o"be���i��Q�L�u�,⪺C0'��p�J3b�ۡR��0(�5q˦b̡+�HZ-�VA�y�N������vRP#ww�;��H����+��)9%� �b��X�?cO>T�UH��f;��,��ud9u���pTX��%GP�_Pk,�E��N,����DӖLq:Wm���p*,Pi���.Cs&1dˎô�q�uN�n�W�yr]�w�|k��R�0�5�Y��T)҆��q��F^E�uC*w/�<d#a���iSJ61*�"�2�C+$Į�e�d�r�Ev���a��R����w����"��uP����% %m��Lkou�N ˧�_��3�}WdJ��Mf�ʋ*��Tc?&4բ�3y��ET7J���YDX�r�G[����Zf	Fֵ+E�����e��
4�\�9�d�Wy�Tuk0�Z��XʍRܰ�A�sXj�-V��*�1L*��2�\p��pͷ4�q.aifV6�����V�U\m��e���j)j[bZ��.�n��[��1+r�`�-U�Z���j�#m7�f�U�f�`�[be�e�D����lhܵ���%���8�\Z�e�j*�(T�S9�e��+�ư����q���t5Q���(�A�V�(���E�%��o�0�s����>'k3�-�=�Q��S᫩v�*��ڶ�	RKX���xC�Օx�bă]ͽy�U�Ǽju�U)��V��q��@��݄n�ҕ�s��.6��_4�Δ7{�c�0�|���������+��Z�Tfژ�W_%Q�gpzV�⽈�.�����,�����=�o7��<h���p�N�|X�8{Jd�h&oR7��V�E�צ�c�َ����+�Tb�wdf,[#6��μ��7���A��=6 u��K���9�,A΍�{��z��﯑)�"j��W�6��}!8�AT�g�e�h�~nk:��xTl鬣;zu#b�F������E�#`m�'�9|k6���=oޟՏ����;��1����.�]�m��T�h&�0Z��F�Q��/������/7�y�7V���vU��W}�wG���uc��Q��&ܥF�V�O7�ճ�S�yn�#^��l�.Y�oS6!vw��i�]y�Vι�3#|�k�~^�Q��20�cދ�zvx���B�4Я�g��<j�x���6I��LolWEH����]���kVEP�7k
�9�!p��r4]\��yi��X>�oG�Z�[�9; >W�Nms�
���UF�7�J8���g�9Q��f���؀8^c��B��;�B �;�OTm,ٮu�׼�^{���|���ci:@���@�!�hi�0��d����@R�I�s������>��x��n�v��!�+$3�t�ԓ�w܁�	��c$<`a�,�0/~����}���}��Rm �,=H �zȰ� v�G��L�d�큶bCXx�q�C$>���~o_}�<1<H��09�o�)<`Mya�"�aݐ�	��d
��>$��� x��w���~��y��zI����P��3(C�C��9Ն$��݇��CĞ$�� v�<��f���w֭��f��߾:C��Ձ�'5�� [d��<@�L'�{a4��k��Hbx��<���޴;����v��v�+;d<a���Il�C�m���s��:H�^sY���z���x�=9Bx��;d��N}IY���NN�'�4�t�I�"�S_��{y-F����y5�Ky-�T�ۋ��+aɛ~^�D�+܉]�e@����(v���=��"r�4t��¸��b��$�b�ɞ��s�i�<���;B}�� q����T��x�<�i2�́�I�m��誯zf=��Y�1��8:�Ϙ��z+$�����l�=9C�8�4wd8��$�s�cg�t��a��M�{��� o)!Y8��5C�N!5��3�m�>a� ����G��'��)�>�و��~`w����}��{��dY!��1�h;�x��m��!�f���6��=Bs�@�{��֜s�}��}�4�b����:dY0�i�<���0��OMY�!��!��t=Hx���3��|��v}�_=}�%d4��O}ް���2,%<��q$��h<d�� t�v�!�<O;����{{�I�H�N�v��1 tÇ������t�ϩ<Hq&�!���;���>����>H��N�T���t�����C�Y<aR����!��'y@8��ߞ��}��������d��&�Hm!�Ї��Rv�;Mu�$��EP�<@<d�񇌓������׽���N0���	+<C�Rq$��I�'!���C�P;d>H0�oܷ�;�z}��,rD]��V�I�y,3u�TV�z�0��EW�dw��W�H¾���?O�W�w)��:�jw�!c8��4��Zj��Ƴ1"�����c���n�z#�#&!�l�Ht���P4���C��wB)�������{�y!�;I1!���!g������	��RN�V|��z�>d0��i��>�λ�[�s[�|����$�!>H���E���;a���x�6}d���$�R|�<�������{�w��3�u��i�NuBaC�x��	�ݐ�	��M2��SL��C~PI�XI/�����z�>�$��&�,I���P���2�;Hwx���t�i';������ē����w�w߿y�f�wM��e$:@� ֬'�;ġiӣ}�����<d=I�I�<�{|;�����>8�>�6����2N�:�"�=d
�L�7�<L��tɯhx�5y���^����}���t��$;O����t�x�i�s��C2�&d��i!�!��:d<N�=1}�{�|����;Ht��VM2��;B�!�E'H i���Rqi ��z��߹�{���HbI��zj�ԇh2	��L����x�o������I:y�	�C�������6}����XR�z���P^�Ռ�G�),7q��>��nD�3��w�KDF_.�j����l��7�9=hoJP�,��늮�SAG.�O�=��n�Q�G���1	���l�&��āіC�L�@��l=O�Z�:a;���f�������v���$�I>CG,� I6�!�*Htr���}a�OP��H��嘄>��N��K��}����|��<�� z���d��CĐ��i�C���HAL��T��^�N�7�^�����@���q'����OXz��HN�d�!�Mua1��H��7�N��&������w�x�:A@�!�T�L���|ɫghC'��C_P��C�%N�b���0:�޻�]�߼�<OC��zȲ!=d=`,�k�HY�|ԜI4�q$�� �v�2A�^�{��>o^|]��aY�z2|���!�l��uC�@Ω��<I��@�"��<B���=C������y �Cě@1�� �ΨM v�9d�>��OMy�Hx�hd�!�tyd������qֺ�޻��L�$1�}� iq&�@�$�N��'=a"�و3�O���>�U�٢3��&�,�O��#�����:��_t}w�7]m�阕�寮��v	ʂ�&j|s�w��+��w���u9�]\%�-f_p�r�T:����t�wPw'iZ���~p�0(�q�ƿ3�9f����1.kN��T3Or ��)Z�o/��Z=����?{ڠL��[~�=,����������`ӓgp������R�2�]q]1���R�9[�3����Ox�o�1��enmn֙[�	N�����}���c6,Ș|���q��Mxx� ��ܜD��$����.���V�R�s!X	�p��U�]zPrR�9�ޢ6�����,����}�}�cbB��B^���:-	'�{k��X���ų�K�;�E�O3W�5�2�>�s	��]6���ﾪ�B��u]\}V��F�N���鍼��e+�m�o��ŕOsI��`��;\{���>�6m�K����p'�?�-��������@���Q���x�}w�Cgh$۝��#�V��.֬��-�ʷ��6�qg�9�Ľ�[���x��ɾkD M����E����-W)���א�؅g*Hk6g؟��Ge�u�s��1|���*�l�"i
y]�yN����w�԰9���8 ������&�5�u�쵴ss�ݢ�����
��K=w�e� ���;��9�\J����=In.j�����vQ��ߵG�~����q��a}呰A=mQ&dC�w��]ۧ��vJeS�j��'��;���>�� =�ҮgLk���\�����HelU��B�Ok]������H���\�"t�yd�P:��)
�f0���{��6q�O����q�'�����8�n��u�L���W�~�of�4ތ�Q�nz��h;�瑷�f�;�Vm!*��i5�w����J�vZ�=�ɶ_S��D�E��w���3+�9�Vٮ�ar�I�Af����O�+3�ohkp;����D{ނC���n�{�_]g�g�e���ֱȠ[�ˍv�E�q��)!
�-/W�O����d���ӱ�����h�:?����� ��p�l�$�;�l3v�<�ʅQ��H�W#�X�;^�+�<�:���"�Ne�J�Y����~X��͘6%���㡢�V��SY���@t]�������b(��h'��2r2��5u<&hMf�����˯z��������?߾�n�ڍ���A��})�m����zj��V�2��E�v쿝�3��r��2�q��������9L2�r���o�q%���ٵ�q��ߵ5L��"�R-�2�m�-�������+)\�Ź�>�{�>bt�C�r�_Q�I��۝�0�{m�-�v��Z�G)���>;�Ӫ1�d����k�Y;{sm�%�K<9��2h�7�uU�3a�KiM��y�����r��n��"�Z��� ��ƌ��vu<���2):r���}��t�E�W���اG�ٵ�[���)qi3�$ޭ72�p��1����+�wX�0����C��Y�i��m��{�,�(woM≝7)��'Iv�prX��7���6�WIS�k(����뒻�e��mHl�J�6����ڬ(m;57t�[�(�Q�oAPlA��0U-�O~S�_�Lc��'���?S��<��[�ܗJ�����f��K6-�Wp���Ԃ��U"�p�N�5W��*k-�o+Z�,�0��i#Mԩ��n����^P`�E| (�����:�n�]0v�#���j���Q�"�8�]��*�=/-�Y�u�(]%��X�M�α��&�**��-*e�*��l�.�fq�ʤF#2�r��18,F	��7P�9�8�&ڻ��QbѺ��D����N�4U��n�A"bT�b��WN�@�ܣH<ͧl�["�I�)]J�`���6���E5pZL�@5C꼬�\�B�nj��J�
�M��+�M��m'1ec���֚�wX]4��{��k�/껪���*��4X�ёb0EZR�eb"�c��ƶ�A""�1�A�Q��[H���2�,X�E�VvPQV)�V,����"Ԩ5�*EWv\�UB�T�-&�25
�EUa����`�$ZŒ"�Tcir��U�������J��QW��J��n�F(�h����)"�d�.R�e�����UZU+*"
�"EY�Tuji
��b*�E�`al*��+4Պ�"�"(�U"���ދ����/��t���Y��:r�*��K'F�Nwb
̑ǭ.��=�{P{���;?�Tw߭����S
>P�Nq���;p1���"N�c��nl�Ӏap�os{�C����ԯ8���y_[��ȧou�1~`a��n�a!��]}�v�� �7��<Y�F��Z������qT���x��͇���z�L�`4]j�m�)q��ͭ]{\�MFr���(���2������:�&��p�)D!R����[T&EM�_�s�*���ӕZ����E�'JŖ�5�˾�ބ���4��s��Л���K���֋��v�V�;$����z#ρ���y���;џ.N���o�:{(�B�e�}����#��y`[4�Wه��f�/O>u+����[���c�q>a~U��V8%�;3���K�sΝ����v���c��]y��4�ᓙ�� ��z�j���Ԝx^�l�8� ٵ�Վ�62�^�6����8�C���=kC59�kw��Iy���v��89���Fk�S{��ך����S�X�mSb�0�\���$�/��J�2�U�2�9s����Be�Y"&��AY�6��P���<Z�P)�7s�Cyr��_(9:��������ޮ,
x��lvw/���=�A�%9���j�$�ٙ����S�/��S�E ζ��\���xG�j���r~�l��{�r�-a�=�1����4���;c(�-��8�b�gmLL��&*��f��6��y���X��䧇��*7��lSY����igI(5�=�̱����vm�9S[ E]A�		�7$� @| ��La	VZ�zayY^_\+ƀ�`��N¼F����F�O��y��Ex�� �e�"D �<��!���D��~��C�y��n�G]h�N�h}퐥�W��٤£&Μ�2t���aV^�t��"Ϯ�����i��Ĉl����h���Z���z��vdr����İ�8�k���{5T}�&@����^B��������^�kD��ͨ������ 4&I��UiY�A���]U6���0/MG֬��+�F
�h�(Q�U���{:�h6���T���y@�p�kb�%@�S�W��{�M�|�!��O���6k�f�&H���j��gg�$�@��:d�<C<p��1"C�U�`,Yy�[7ozv��N_�<����B]
�n����e*��~�S>����EE�7O!����(\!^WLw�A��
��ڃ�8w��Q����S������)�������$:f^tߑ�c�kx��ۭ�*���c�-5��~Æ��2�ٻ��h|�N�ff��OLEON���"�:}��_!WhfS���+ �ƅ�y�t˫��t�p�DaK׻���o�Q������̏R�ŮS7`�����IH�{��#���������5�xF�Ցai
uAFy]����]¯E�\�����s�=Nbg�	+��C�EƩ}S��Z��U{�����uxm0�L8�2�:J�3�	1�P�'d�w.������ӟ��m�ɰp���C����ًCIt[�zoy6lӺs:+g��I�C&z������9�����0R�!�B��P#�,ۻ�f�:�W%A��d����v�<���^��%Jᡉi�KXM[���RXw�F��۝�=Kb�U�b�5��͋2!O�fn\��u�I;|S&x��4�9�������+(|�
[����A�Ͻ��:_R�|A����l�MTqo�U7��m?��&J+z�p=w�yx4����7O0\D�)�>�ys��[Æ��mu�������A��Kt�vf�D�ZK�z=�G����ٹ���j?�Eg�.J���<���ӌo�:?z�/�|��
P� ��4E�[�u�.�U�5���
(_8`_{��1ݰ�0�--�!��ǧ�K7t���r�§+R��(��H�t��W��g�&�lW{y�Y��Z"�||r�jGy|�Z���:WF3����1����^���Aq��ƵqdiҼؖ��-,���:~�m<��mM�<Џ�%�����ƱD����
ޑ�s�f��<��A���؂;�>�%��"E��'T�kڋ�}}�����Q;TvG�C�s�m�l����׾��%g2򺟶�P"&Y�wY�Q� c�0�����!��-����Xϸ&��bL�Ɯ�ٻA�3�l�:�ÑU���������T�lIZ�J����d�%�*��uǇ:uX5;���<��Dz#ϤB���q���}��-�90�0N�����N�x�g�
�b*՟b�z��L�A��f����+���{����x�x�S^4`#Og1�i����X��t'�`��@&Ijjnv�z�]���U��+��MEpۻ�g�}T(ժ<h�><x�Vn��v��\�z�e+|�z}Ӑ�ЯT,alޭ�6CK�����2XPS\���F0g��W[;$�9ؓFqT)��d�n��}D��3�5��mڜ��5a؆��2^��Љj#Ԉ��s����z� @��+���/�:,R�#�ff�\���s��[l�O�h����O[F�8x�[�6�^�S�Ŵ�s��G��T�sH�<���$��;��w[zO��cZL�΀H$�S����|����o(Jf��Y��)ll&Wi�v��.�{˄Z�&���az�ڮYcdG���r��B;jJ<�p_������4�-��R'�T�k�r�ӵz%̫���tnlh�I�+���	元�$BE�X~&}t��Cϭ��w���Z�1�q�U��"XE�bu�f
��u[�Y��2fe�:R��L��Pn�D䙙B`��� �T	[N^�(�|)|��Yߘ���Wȸy�o��M~~0�&͞�%����*i�^\�e{������
��	2��F]�<��gZ�����7Ag2���v��E���M.���z�>�Ǭ-;��+mS���v/��F��m��h|�˺�Y�gs�4|�IU��W��+(��.�X�i�j
>�ZY�^1��2L!t��<�ť��&s!BM-xi6�'s�2�ꏽ�����5�,�!�fadh�Xն1�X�x`Շ�&S��wJ�M�
���\:B��R��T`�j\�Z�
�U���č2O�ՁOh#�����/t�0��N�HW癞�/��G�~j���e��T��2��/C罐B��(�#=i���=��oF*��@�$�ˌڅ+�+_���(��'O���h��$���_Y�󵜇||B���9�/����9\^>4r]��sE���_���W|�_�]���u�[]�R�,��W������W�b�Vxא�	�Ɔ({�����dz�ۛ��'��ȟz����R�|�t�AO��l�g̋��eJ���,��*�Y���W��/^�m<�yF�,�y�,����{)��e��->��[��c�@�h�QV��V����ʬ��8�0�^?JL�jا��ޑ�'�[�m�C˙ʬ�]�a�<5z+0琄ML�/��YV�x<�z�볮4h��!�Z|1	�f�>!K<tx����RFhҕ�n��=uw)<����ec̤³��!M�߹V��ׄ
�_xѨ��-��|����e�������%�wK��
6m���s;��Aƪ��G.� �jǌ�8�fC{	���Z[T@E�x`�0�9����R�3Ң�J4�t1&&-!�n����"%]Iz�d>�(IM�sU;*MňҀ�1U�NL�理��m���u:i�H�US�()�JD��" ���OL~��XR7s�[��G?�z��v�4���l�i*8��X�He�����ꉈh�k�|8�	+�P}%n<Q��]�w�&�}���.o{�]t�_FO)z'���ΐ�Ժ���-��b:�ۃ�)��E�Un�ۨT汦���U,���w�:�fkě�1bSn]�6�K/��<��tSI����/ǥ �n���'�W|�!�,�KV�.��\�+�ٜ��݃p�[�_ �n��/q޳JXE�����s��s7Ev������GyEV�-�.d�R���r��.�@RV�1v�B��a�U��p��)����;k4��ا�Fc�m�e��a����!c� ��T����b��m��=!wz���k0�Wܮ�Ĵ:���,��Ν�v,�ڹH��3{yk��9 5�<��Pr�lHN46��~x{*�$\­K�y(���D��Z.����\,���Sb\2��)��ʚ���M�C���R��h��jȌ*�g�J82��i 2�C���Z��3���r���Y��˻"S���:�J�ZU1E���P伟aG+1IВ���@�e^��\�<���82b���.�*��\.����h��H���4��ˌT4L����a�����D���&e,����(�M��k)X��*��Zʪy�Ju���&(ةi٦%$.��!2�UpL�l�H�:�V�4ݒ�j���w���m6�m:�E4���~ ]V�ق� .�1Q-++U�mEZ���m����eT�n2�*2*�M6�8�r����J��F�6���B�j"$P2ذ�F�j�VSU�eJ�b
P�Y�Q�"MZ
:���Ԫ�髺J������X�Ck[X9h�m�QV,ƻJ�
1UT�U�*:j���"��i�Q�XV�t�(��an�T�V
1"��E+\ZТ�J�Q7er���~�y�>���k6ͨ-i�|	���v��ԧ�b��5�ve��^�DG�j�x�ѻ_�ɨ�cF�}K��2������8F��]|�r�n�n˟	�\:}]FN�T�&X�T�Y�S�[v�GF���{M���	�p�MO�Qְ���.x�7R+�]e�`c]�Cځ=�'�ڑa����6�����u�ݧ�d����]-�&y��;�,��f^��aܫ����Z��4�{�����p��2s�5sy��Y|u[�ֈ��/�{P�Fc6�Klu*���X�^���ex��I�9k�a�_a؆U�����I<�/?[~a^��\�X.����l�f�;N�hLK��.���L��0�x��[jl6��KK��=~d�����ғ��}�Ω)z���%3z��ܗ��G���)�T��(g.�:o�\ƥ�V�
oq��x�4K!� m���xY2aJމ)�V$7����W��֢��I3Ԩ��ޏ{�:
��'�������~ �xl���ærV!��lЄG�!���hD�ՇH�*c%�����u��o��|ЦDH��<�kb��]]Pq��GI-�Tm��_8�/zr{+'������hU�/��}��������qjֽ=ܰ^�^Y���_*��-;`�B��rC��wn{P>��@�k<�#�,��<���D��{�ݽ���4��Z��!������\^"SxGU@�$�r{9��]���D�lL��Z�ɐ�)��+f�Lٮ{��c�l4\c�Y�O��@�Y�3��`G��p�#Y�'�	�WW}~�%��Vi�HJCu=CO��o|y��:�7�֭<��!�n�6�m	������{�˕��["���z"3�o�b>���t'<a�Jr�ЍB����zj�wT��X��Ey0���	�mz!M8I��2m�&_I>��o�5�}pv�����<�/��2�$!��y\_R^2q��&�e|C��vQ��[���O�}b��`�Q@���+}�>�~#�.Z�.�a�J�j�dY;��`c}Y;=�h��@�.F�E�%�z�G���T�����-*��E[�;3.cf�=(�y�qi��Mf��Mi�x�<���w�*c$8��� #�V����LJ��7�C���)��]v����(�+���N��Lo4y��3�2hʏ/�PK���6�<..5T�C�3w��z󫄪69vC5���5bv�b{��ا���Oޮ��bš%&�.i�2��D�I%��G+�=f,���*2����d�l��UVc��Oޏz=�A��)~J`��(!}�i=�q�\Z�ܲ$��9�ҡO;{n�~���0Z��D��h�DL�L�1[<j1��:��K�W���T\YGv|g�������p��G�׹^�rI�~բ�]��wU�/��fj�LN�<���(�C�� ��x 9W��.#-�!� �����^���Vַ��>}�oֻ��0�oe��.v|��f�1o�7�X�s�][.n5�r(��|p��5Q�&h�2�lY�x���}+���=n
�K(r��~�\(F��W��W���;ซ,%���;����p���u����ɀ�H�ϼ�x����/5ўl0�6D:��wcq��s����A�F�W4���1��ʷ���'�n�=���.:a��ސ=��6�y�fI.W:M[ə���1r��DD{�G4�\r�~��z�w&cZ73v��XQ�'�2ma���{�I�[�F��<dL����w(||k�d��0����g��ߨ	qX���o)3/^`U�6k�,�)+k7�n?�)�US����>2d� 4��ؑi&����x��g�R�n1��1��&`p�mJ��*.]f���M¬�5�z�3kn��+��t|�3�������g����:ZU�<,Bt�q�Dd�����8��Mc��D�3P
���+�{���y˕��g׎��H�r�C����U!�ANuʈ�=��V����J�#֍�ƅ�}�M��rgMA��f�[Sx��vu7YY�N{�%�Z��;�K1XR���la�W�j��{λ��G��`�ZI��*o^LW�Q����$���-�.`⋏"ٷr�8�;�� t�Pp���B� ���A�Ԩ�ވ�G�]����^?�l՟Fc��O���:+0��N�۾s0�|9q��
h�h�b���_e��<\������b�V�sc�r�Vk�Ν4�(%ǌ�e�;ړ�lp�B�sw��E�#hx
N�Չ��r�x������ڂ��<�'�^��ӳd��$m�P���|��\����Q~�.�gϺqe8p��W���5�#�%f.)������٢;�bi	�{Xy��.hi��V�E��6a��8A����+Uj{rF��Jvi�U�C�*6zE׬+<~�W����k
K�}[��Q�}kڣC��B�Yg��"�,4B&P�:s�`Jd�Wp��>x��0ʔO	PQ]�6�/�jtMRzܕ�&��χ�>�МÊ���;Y1����^�Q�RkXz����+-��T�7�1���}ց>�Mb�܉��{#��%�-�v{}��^E�XD�	��z<=uA̻oKWl��:{]{�<��w/>���c���B�-:_چ���#2�x`ւj��K�������ʃ���l��hdo�<���]u��7�)k�<|С�-OS4,�����U�7��^�����1=���n8G�f�冧��6�"Z�}��ٯ�r�|�Q	�];8�W.�=�3��s�7���U�+.,#ݹZ�.�l3F��~��w��d����AF8ѪVv�FV���
���M�Ǒ�^Ԫ��Fg��Vn���;*�9O{fQ�[���)�F��wXYp��E���I��sW���:�V����""'yn����Q��XI�XQԃ��陮ύ�]��u/����1�u��)
�G( A�B���{��w�3R>��y����ɍ��;<�DJZB�Ɗ��܉���S��*6j�3�fw����V�.5As��v}�3�j�<��x���fUGNɨ6��D�[D�t��_&h�~�	��Q6�Ш�{5�^������x�!⚙�	ˎόCA� �.�m�k*-v��0��U����O9|��N�K.�׷c��s��} 9B�r8vX`��dj^"��S­���Ռ���锲gY�AJ��÷�Q`�(f/��b˼��ƦL�M�-���U,W�`�#3ب��'T0�TzU�A�&���t�w�L�Uj�ۏ�\��g;�ʓ�	�sv$~��G��o�Q�S?G�6nT�B�N��h�<׆&j�nO.�T�a;�k�՜.�ׇ״)�V4;����K�9-6{���ݝ��u^���w��	�����$�VP�<��q�����	
L;vn���(^�A]&����̾�+���.����1��^���l'0鶨���N�3��j/Q���C�hF�0wV���hח�v?�e�fq�D�J�'�66|vF3R8k��e琖�Ow[���-�� �ӥ=0eD�2 N���%g�tџ
^ǈ��RTh��X�N"{q�xNͭ��8xe+|`��yCD��qq�!J׼���|�{�����Z��|:QE�X������uy/	Zg^�[��U�C�:g�;+yݐ�wm%ۍ��[��bZYz����Wnv�r.����x��Җ����t��R�1&ftS��1c�&b���:�ģ���A~��DS���'5`���ERx���������i�ur�Ju`3n�]��R �XCdZQ������ن�Ș=R#@㸡�Zt��8x���s%߷ͽ2�Gޏ?`(�ӄa�3`c���L�[�uޗ�y��ʍV�>�p�0� �$
�m�[�9]���/�����y]�`c�qY�Fƭ-�Q���v~����5�ʋ�J�]-��^�N�0�{����Pg�/!��\�d�#�u�n�g�R�V��{�?-�kMI�UU^{��g���֡�>=/V�i+�^����N�?��3͌�F�S���bT��"H�E+6������ԋ�Z��g��6��q�^gwm�!���]��Xk`=��l]n���ov^)�c�g2�T�c���\�bVx�k�ya�Od�xy�SR�E�r����/	�4����}��P_\�.�k�hP�_m��Hz���5}o�L�˕�@��#��̪��g%m����"���Ud��j�ݩ$x�f�@���aG�kw�q�uSI��^���]D�DΏ"e>�7-�M�4U�*�}���i�Ko��S�)ͧs�V�����+b��i|�J�����芤�,��1���e��!��9�s� u�yJd`��P�d�r��{i��l�ZVJ˃�bt�$�����s�(�]uu}�,��nVS���;���SC/����ѷΦW%�����L֚����{����	�f�-�56�g��~�n��Kp-�"�aD'&��d*m��e`���r�]�nt�=V�Ƨ(*�g-ۘp��^I,-kx��9���M	F�@�F*��0@�nD�V�A�]Hޮ���x��O�0Ƌ����7�Ξ���wV{ �(� �r��q�\���#.�^r̓���S�sw�<D�n�ޞ�51B9��1�b�(����t�۲s �G\�5��ܪ��y-��	
{aU���G4!�}���p�Ws�=1��f�YJ�jv��I�]����_Ws�Aq7�OT"��Y�j���	X��,��nU�
X,�ͱ�aδ:�j�(�uԢU�3.�{�rI$JI$���RH�)������f`Kh���N�X�\k-���[lDAx�qQt��e��,��XU���ZU���IM�0MڻJLl�E����ƶ�Օ(��)TDE�2֫"�%J��)�\�v�UV�.�I�����TQZʢ#+P��QQU6�k+���ƺ�����lUEJ&Z)�Lk.UPwn��PQE��Zc+��1�ݢ�M�me\��j#��¢���������������mj����f�)C�)GqI�m#w�ܿ^�D{Pפ���]Bj���k�i	�{`��G<���5��J��z�$�5���c`��4֚Q�ڃ0-�A̅��a�Ie��Y�W�$&c"�~v5��~5��t#�g��g����ls����l��dA��Ôv:Õ��{3^�'A�y{�q��m�(r�n�o�C�\����&CBdw*D��P�Z��Vy�Y����z��jDY��Bbϊ!�Gghy�0^$�'�����KK����:>"��^\����������T5ɟ4ĺ�w��>7Q�Y0�_�?s�@�z��b�d����Vڞ�f"X�y�b��"G�͍�����{Υ��Ѹ����y�:vK[+��QJUnd>Tm�W���Z���T�M��z��z��I�=�*8㵇e��>����G��i���뿃<p����f�<B���U:g�� �d���0���j�B��y�*_�T��H���y���s������DTGw�׻�4��q'��B�tE�k��'N3��X.b����TU�p�a�y�'�n�<(��D�rf��roC�SSq�������^r#󟼨�l$LCܡ�6kP�3wy�3p��QQFTԩf���*�G�֚9Q����Y�0)�e����R��B&}�*�������^�Pz�b�)�����j��3�%*�&o|�����OM��R�e"�̌��t��I��.n6��DL��,���3��fiS���V��i�hdx����'3yF�u���Rq�U�f�6
�g����uh�Q��k��۪���f�m_���&�g�HdCօh�ϵML�E�e�uGP��������V��ٗ�;�0��ǗR��-!���'_�J%$��l��mC����d����J�:��������eT*�dʂ�E�A�78S�g�ޱ��4e_�>e{e�>�k�L:`��c��[o��'1_]YL��w��u/x}�
X%����B���2l��5��#�5�:}�� ��F�cYG?���F�Vw-����>�+e�X���Fc\%fL��tg6Trd!Kb��=��x��ߕ�C9|��po�;Y/�:Q��y�{&����!�:|A9��{�b��D�Hl�s�����t&�pWd1b�sƼ��u^X�����,���5�&n��o�Lǋ�T��k:9]��p�L��}� ozlɓ� 1KI}�� �ss类jUT	Ŵ>�꨹�<t�Ԏ?W<Y����j�x٢0�����}zƤ��>|t�4���VV�����V��H�:P�<t�3��c�W��������s)����A[�5}����A����A���H!�Ǖ��j,����C����q�IT^0�XA#�x��Xc~�o_���k�t��&.�9y�؀q`"����_��~2��5Cؑ3ϏDe� �L�DTθ�[Ȓ���0�}�S�
rD���E��5�|,ޝ��6�ƭP�xdA,d�<~ù{��O�{]p]��$�y����0߬[�{~�r�ݫ���V����|�^�N;�&]���Rx3��oU)q��R���5����O�d�1qV�r���mh��u����s����~��λ55�T6����Fat�sƲu��~�73#ҥO��'o�|�}�}��O��?D��A�W��aZ���̬2��W�;��!�^.��/]?�Z�w�M�p֠��c�m�˛�ڹ��4@�������\�MI���1~���88�v&z���Bp�B�؉�A}x�	_-���yW��[U��XgԼYZ�f,n�0�:A���k�M!����M�>��GJ>Ԓ�Ƒg���aCW�
�pJ��yۼ�D�2LJ�r�ʒ��'��پBH��gp[�o*U�����B(;K��D��21oA�+cA����v�8IO"�
`�E�gS��ꉐ����:_!%gRw���Z�m�������]%���U&�t�y�K1�ӵ�Cj�v�9KI�Z�8�㗚�h�P��IY�\N����=�����d�
����S�"�4}^V"i�R{��M���)�O�\��{�o�t�	j�g�)ի��YFli�N*����T��j�4���U�e�j��>6Q���%}-�{ua�7�����A^HF���%}��drB�n)�a�в:��G�Vbh��ɛ�Rz��5eŝ
}��^L9�6��.qif���O��3HC�7�
���5�|��(��oy{х��N�z��>Eɍ,��ڝ!n7u���9�e�'��wL\��]+([��ZJ�Zô�k�S*������J!ܽ�&�=ω0�ŅR�R�bE��Y5%�y6+�.zN����̯p�wT-ښ���E���So�(��+]G)��K)nR�/�v�Mڑ�Ϊ�ɶ�K�K���k�N�F�WDkz7b�����U��H_"~�DAaE-�f�7"!�O�5&D2��bb�I�]o5Q۝A�G�
�k�`����Lų.��Ϟ!��Üx���i�exm3��TA�_^0ů����ٱz�vv��,���Cm<^8a�U�
?b�	��^�M�Y(g\�����.5�P�zD��VhI������o��W��T+T}�Cܨ��~[HN̝��E;S@��yץoNP���!�܅e<>0����L�1��ZެZO���li6�b����v�=�B������ݦd��Rڨ��D�ʛ���I�Ԅ,n>0bS���]��M�e���o>�,졡܀��� &u{��i�J�e��h�
o���']���fP�I�˯w���9�%Vkw�Vi��܎���v�]o�e'�m>;��s.M3����*�X����8�s]R�a������|<ä^�F#�w�n��K,�{�l����}�xSϽ헵�pm�̡f٠����Ld��,#�����|�������=�Dц7jU��y��r�ց+U�#��0bgN��U҉���1��^W��MY��L�q&&�=I����l����z�����kW4||z!-W�f�������V����gf�H�Zs�zX�H���:�U\���F��V��TyL�
}h�%���M�:~f�����1�u��"�'�=��!On��!�@Ȫ˫u�Et��n�#^��9s
#Xs��9�e>`,]ˉ9z�+�P@ER��
���_�y���6�����=�S��=v�&vu�m�̱�;_�ؒ>�[$���qmwÉ�Y��r�Ϣ�8��;�h���^>No�z~cf:L���V�I�0�3�s_	jN�4���a�:���~p�:~�F��m��j�}�;�uHի|(R=�� �5e��@�g�a�͂��\%�=��n�V��燺i�F�^�,��M�2�6]���NN��E�����n+5���:h4N��Reg�״ek&�զ��c<EҭR�t0�x���Vi����l��q��_V��:~7;�[f�ܺ������qT������Utv��(�Xw�{7��N�n��Y̜?xbj�ha֠HNVȁ���5�K{ŁX�B��dzL�ׅ\��#f�a
���7H�@�&*Cb3J���Rc@^��,��^M�oܕ��������վپ^ 悞��,� �s��|^�ё��W'��-���Щ"��q���薯551��d��2�bQ�����vL�T��;�J������^�Mg�&��I�r�!D��VY�$Cn�]o�`��P�L$�VG��dA��B"��W=���RE�%��H�n��5�o�!=̜<{�:J��iG�z���	��G؉��@YF�W�b�@Qg�פ��&K�y�;H�����r�|Iiv�h�&��}�7j:�]w�HE�4��ck�e.�xyaG��I�j*�w+�"f�;�fɺ�<.^Һ�v���Hcv6�g�>t�`��.;��Tk�#�p��k���x��������9�HX�|�߅R�qڂ�`��_SS(׻� С*f��w�+9�Vδs�u��L�3'o&�j�t=�� ���MW>��9�0M��H�B��M�	C��MP�v*���p�p�S�j]�){4�^�\�U5�VU|z��aa䋬;��OWJ��V.�T�O>�A�s�M rp�Q ;��bɰ]n���/���j��O�/%Jݮ�-3G(�c���B�=x�
x��e&ط]�n�v_q�N����&d�*Τ  )�4�V�c����o,Z5��������il�x}�k}}D�O��#+X�I5�d�63.��
0`��_S�WC���"��`��˸Г�g��K��}A�mIS��yŝ�l�R�P�W��d?r���ER��Љt���3��qY�ׇ��'	P�J�K;x0���dr����b����J��{��n�Q��N[��bjVSW��yz�dA�m�e��\��[��c�f�rXf��V��z�uI�U���Q���:��U�Z����۬�OT��tf��%tAʓ�S�D�V��ջ�=&92�/�S�R�#S	죋kw:�Di�5�.U.�pa���;l��TEwL���@��I5j㵲����.ۦ��l�%�d�i`��$�+c��R�е�����I��.��Oj���	Ŭ.���e�� A�.�"�R]q�DR4��߹5��W>ҷj@�6�HM�^�2VՌ�}�-��IE��Y��LmT�;�����M�=�`��V�rL �a������w&Z:�;��[��v�1�#������ɝ�X�*\���Z�gc�yU��YEÖY��N
B��L�=�!t���jq��˼��wvr�Ao*ErU��7Xz���bQ���@��ʢ�ʊ*�����E���Dn�ưQݖe	��ԨȪ-eA�h�E#���YH�D�X��)�b����DQQ��A�"��Q��Ddբ��J��)7lD�*��ZET�"m
�*�(�cR���s&(�ѻr-�ƃ�fQX�R�T�K�sZsNڋ���f2�fb�eȵ*ň1UT�(��j�?�U�{�<���Bv��q�r�Q�|]�Y��!��Z��ݎ5���Ѵ�)���A�j3}5E�Jr�F�L.�):]J6^�]���2\��f�?a5o�DQ�4a��g!R`��}��,KW��<�_���]wµ��������@�B���,�2���k�����[߽�R�(���"�W\9�Ï��C���v@"6���!͊��������c�qʒ����!��u�V���ʧ�H�|��	|��;&ub�&�%���Zv��9a�j�>W�a��vR�g�J�ƱQ>C�5���f�͚6��QrǴD��V���'fQ�d#��Bǐ����51KKq���u�穮��2�g�o�*��v=0�r���%n{�z��۶���d��hl̹r�û$���c.MdNgF�ɼ@�M�Iv�
}�SaН·�K�Օ�v�G3��ȅ�.�S&�<ʛ?�ش��(�A�Pج��(�S�*�0jؾT���iX����Ǆ�ln-0׵��������5����skM8`FȘͩ��ѓ&zYBLd��>���4s/w���wk���7N�!B�P3W]$Ә&�o:�R�m)�O(�u�[�پB�'7W�h�ⷋR�{�U��cR�X|y��/���+#L<�����+9�o����20�{��O�1��k�=���m�.yy��G�a�PŇp,>:dL�駨 Z�F�˝Vv����F�}�\G5�B���p�REA�ѓ(��ȓ=>p+9L^6F�h_֫��ICˈ��7��S0$���n���::�)^HP���zǇ�������c��p�	�l��f>9e�]2�V���ÅU�O�ה�{���Hĸ�I#u��t!��N7t�Y7CL���U욼���D:W�bZ����$C��le/�䪥W�̾~���j<�~ZX#I��O�׹ф<^;�wY�X�n����9���=�2F�ǉ9�oA�iF���h����]f�zt(�;��s�ʿ0(�AT���k.
�[���9L�G굆�q�gq"3��z|G>}���ٽ�A>�/!V����y��D����|�<�%V�zU�=/�)�ek���Ⱦ�[W�!v�C����J�ĳ��!��m��X���g�:eퟡ���v��[��Ke��]K�SBF�M���aٯy��su�BIS��'A��ݙHsPa#"��sFx��Jr��=����
TzP�ͲE+���	z�ßW���	�r�PW��{����޾Ky�]mT|*:FW�(��B�\��\c�Z����Xw���G�W��5�q�vô&!��&�qe�����!�N���:W�,,41-J9?k�>��>{�����8��I�GG��~���ņn �nE�`�+�<���H �yRcg�b��=.7������9��/�-���y��~{���w|{��
x=yO�чS��!��D#D�AO~�K��8�
h��%����tQ����ڨv�VP_y{`%�D�\{٨鷗پ$��0�S�j&j� ������+�:dJ�ھ\��]c�s�E�&i�W+<'N^4F��x��'T�����9�6���m��w*	G�pص�WN�s����2Z�ұ��x��W;e1߅��g�p�VS�H�9�N��J�;���D��sWsߐDg������W@�nN�F�+��<{����ug�<-|����J����b�ܔ`��	�!\�;��2{]�}\.�ݸ%�>=��"]+Ƴo�{�
�["n>��J������C�K:@��̭b�b��)�� �:S>��J�vbߝ2&�]��n;�ֶ���4Fa����{��j���)���A(��F�������ٗџ�%˘;�*3+>��ww�Z4qغ ݟ<@3����x,����~&����ü��-��H!�vsAN����� �6X�!��kqæ��t�ld��n��ٹ��Y�Б.Uh�/=0b�_��>�����*�gΜ����N����^�����"UHaJRJ�[v�(����`���mྨm=d����\�ꛓ������z>�{č�m:��q����G��M�	����[�.aGIm��d��3+Hsq\��qA�������R��z�n��u����	dq��<D;�Y�j�-,���vS��ڇ���b��i�J/�\�!*��.<7=5V�۽�w�"ȳ�C6�ʎ�0ʸ��E����k���̥ځ<F%;&[��5�.�uuT����<I��A�~��P��`�[ɇ�8s5�F/V�o�����KP{]����V?�[��զ����T��xz�ު�r��1*��j�-�VU�/82��یu��k>�\%�;G���l�n����V6����s��;�N�լ�r��?R�b���$Bv�NAW��]!Ȍd�^ ��mI�N��������/9�UI��ȻfKk6UI���p�ck6�]u�K0�ͪ��n�6��$��Wa�����Fz{4R��4o�,!7 �q�~wʎ����H�k&�:��,�TC2��,!X|t��ּ;<�7}x�E�D��7���튣#ʮfnyط0��g�򷯩ߪz�OVH|@���զ�8z!-W���"�m=yt��đ^џ93� ���� dE�]��*�2��Q��ʷٌ���0\��F�X􀏹Y��j�{��_��n��߭��[��4<I��8�:ZF��)�q�:ym�nu��.��~���;*�y�+m�W|��$�����u� L*�Y���9��$p�N�ONèA(����>���܂���"���=y��BЯYCn��Oj�6�¹��Z��s3*-Q��<i�,m��j�X�a��)wބWbi���:�g�r�����ENñ�w^�+e�.I����;P�"ǵ�R�w:=��զ��m0�6�j���$�}T�hw�<>agR��Wl�5�\a^�;j?y'�y}��_]<�����#"�y�a�<i�'���^5K�l0���it����/d<6��z�M�D�}��\��P�ltH���l�!�z
/龜|s˱�ݺ�j�����"b'�}c�KR���H�����%Q��b��W��gH j���X�i&5�j�c�9����W�uS8FW�D��C��ij$h�1�8\_K�ꕏ��2{/��ݐ�5�[ܫ���gø�6
S+��ف��/o��Շ��I�u��7e]��t�mJ��6cB�^IS2�$���Æ!�I�}�V�Fe�]"��3��n͞_G�w�w�
`�\��9�U"u��"D��k�ڹ�kÔ�CEp�����6��)��1��"�,?z��	^�Lں�&n�O#��|U����DBȯ*���eWGU��=�pF��`MD�oA�Vx_%��sǆ�6Sn.'dM�)J�j�Pg1yo�C\�~XR���q�C���>0��ëX�+?JY�w&<�+��'�"dWԆ�$��s_�����N�>k�f�>䮍�_��Yb�t�Vj������z�rc,�׳z/+�˗X�¹u�ndݤ.��s�!��Qr�ԏ�4��ύ4�%j�$���g1w~s]ܺ�b>g&�dP{�;��'t�V�w��A���ڶTz�u�����Ȕ�)���a�f�*F.%}�zլ\��}�����|r�<����s���u�ʩ6�jH�(�1B�ZxP��ͣ��C�5竪6�>�=�{�,��NM�i);Y:����.�b^C7� -R�>O�����]7�=�<�����\�ӝɕѱ^�Cu=GCW�:�>�{��J�{�ꝏ��k�
s���xA]�]�x�I���k���t�l�!67y�q-��E�nב7����$K���5�N!��23co[�5��+;pM����R{�Dݔ�J�������8�<\v*���BvU<�T��^�KM!x���o�����}�+k6f÷�n�FX��Q��^��aT��E�Ц.9�1��y�I�t�aMp]8E�Z�O4�|�v�xMhv: �u���E�<;���]�W�
�Ւ�6����ڐJ�3�J�,ټ��`/-�ʴ��kWJ�G��g�ǳ�w�QVG��ۤj��1Q7؎��t+<[���}��em�%̩����4{�:�Z��Y6�cI�L9`����;����`��<�k���dV�F~?Vڴڵ���]�h�m.�8�s���i�4@Z�,���q��IWQ��8�3�T�Ğ}/�-���-��'L�}t�u\(�qk��:�vǷ�;�Q[������O@�ڲZ<'A ���s�<�^�'�R�x``�X�Å!&U',�Xe&i�ĩԖ�F��_L�QJLStd�V.�P�k>,H�>$fS���d��d.�e�Q��X�i	�)(0hHQ���,e1��Q[_$-�c35UO7(�rӼ�M%��*���٨�����6s��%�CIJ5S}F)��*�4],/.VP%ɇ2�Y�$��rdßRl�˼i��4��aj�,�D�b���G@��*U�e]B�U�J��
��w��Q�X,��e+�M�8�SϨ��ᡗ*��f)/�0c6��9��̱v/�R��V�4HƮGUN�ҧ-�/�f)D;��QEuB�Ɏ���p�U;�C�����5�[�����Z߈"�Z�Ya�gm^��U[KTY��֔EW$�)U�",F(��b�*�-S-�.&5iSv�Df"�c+��D˙��P`�b/,̱E���9h��m�iQNZ1Ub�-,AYAT��F��[r�e�\��CJ�A�GL��,�1��pEUA(���eƚ�*e���08�EF��+�DCu�߻)�p����:��4qf�lb5�,5w�����ǖ�}ݝ٤O��J����[}��a��q���%�x��ʪ�&��"���2hķ��_�.���v6����A4�כ�uWHW�s���:\��q���(S�ɽS�'�i�>�W,{U^F�ɽ:��v��yT���w{A���\8���=f�b�&��A4j�F�"�W����e��7L�2�}���\�un>�/m_C�������\BV-��h�c��9f�h�p�v���ˢ��a�M�kU�ƈ�֒���+BH�@������<=*�>&0��R�K]Ҍ��pG��5}3��Ʌ�u�z��bf�UU��E���[�4��q-���r����n�[Ns37��)=�<Nצj�Ot�C|�yGe���H�i������T���t�b������U���7ng�����x��/j���{�Oa��?m=�L~j�km���������$!c���c�8o��z�͚]��{�ex�3ϓ�5�\�%{��L<a�[���Y�h%^��ZU�U�zj��h��&�Sm�,��Ob��y��07��!� �1*βb[��^�D�W����C��V��=U�4�q�!,C׊w%Q�CJ��IN�#nj��WU�qmo�wem�����嗜Z��?|R�0:	*�w_n�N\��w8�@��N.�t�1B�3���Ъ���n���omT�s��I�`F��C�@gwr�0K�1��o�H�[}6�/�j��>����u�^f+�����N݁�v�
WU��[��������"��{Pҳ�]�a�r��]���W��RZ�Q}Z���,[y��_���^�c����u�横g�X3&,��Yms��������|2��������4�F�������+j��{��v�8�E1yJ�hV�ɡ{������9���'{�a�CU����4�]���}I�%:8o��g<����nt�3\���b]�r���4����Q�[{x���Q����z��+��b��@q���=��4�;;����T�EZ�#�~��SfRiR<F������-f�P���������O�zml��i5�p�y]C�)��W]�Ϝ�{YXq"��ޱ�5�?^,�l�Js������G}!��5�]�z6*��xz���L���؇��8���b�ϨStD�����b���^�����Ex��]�=������a!_�����ծ��⥢�p�{��5��4�dY:�#ft�[���~�5��4;b����F3��1�ű���&z�s���uMs��1�ͻ5��_l������S�^YRn1��eh��w��L����C��/K��΁����� ��x��)�6)���F˴��2�k9��V���.��g�jݼi��x���(��N��y[ዽJt��x:�8�Ǐ��g�,%�ې�j��{&؇Ƞ�=Vw+)œV�A�6q6�FB�E]!Q;ʳ�"��b8�^�?U'����������)6�&�\gkq2C	�R]i�[Wo;닷�2sg��ujS�oU]n�R����Z������}�>0�!-���"�j��q6�A�e;%F�:֪�|��2���-�ǆ�=�t�[��Hh^]:ض���(5^�5SΥ7%7����9t����<��_JpLo�݋�ZK�'�H&M��\$S|��̵=l��Y�-�[;GC��:j�N����b���V;;��(��W�)e�W�ڟ/i�u��-�;w��o����q���l��≴0�py!�/��k¯�НF{#�pVҺ4����B/�s��p�s�OM��֋��Tٻ�+�v���0&�����Ri!I�k������tr=�i/��Kțf�V�Ú��&�K�.�Ygkz~��
瘎V���d�þ�jk��s��ez��$�K���Ī�U���i�u�Ѹ�_����'GGT����'�z�t�Dkڋ!���77�,�;��nA���fϠ�s��:�tپ��]Pt��[�N�AE�㩾8�8%���=�i�d��)];N�2]�%�d���G\;��ی����H��.8֏e������ux����Ii���]Jʙ�ZiWw���vK��uuWXo�kW,�Uǭ�o�ǝ]6=����9�
r�22	En����Vs[U�����1�^{7�yh�Nc.��A�TuS[[�͘�iZ�)U� �ʼ��� �J�dF���!UVDN7��$l��01�-�]~�7}n2eꎣ�ww{Qc����Ug��6��i��9�$��=�y�U-�b��ݪ�J)���E�֊>�<c(���~W���9ԶT������@i�*O"0 $��fW�$��l�q��((��c|�sΪ���o�F��D,�s�:,����I�F�wkֺ�0Q�Hb�틎uܫ��+xqsts��Yٝ�n�����o�nE�V8�C|z��)Rs�NoW7?W�s�s�����}��t�:v��=�g!,n,�@:]�X�b�]�k�Y*b�¢�r!j+t+���bi��r.�2��8"�O)1Č�wKg��R���QT�i�I�[(��W����O��.�W�Wy�`��$Y���u��bfލ���i$tV5y�d]��t���l�D9��)7�?��:.��*n3�+��k�e4�ؐ�Nlm�z�9>.����i�N�X@"��ʵ�]�'C�qcSp�'T�fkJ��=�Q^j‷q'�%��<~1���$��]��՝i�ѩ�ֶ�3|�'���9���U/a�?y8Q������vV��J&��{�og �ِq�ר�W �u�6������nn�`5����b�ۭ�1/��ث��En_]Y��u|����Ի�{�H���p5�{3�EzF�(]��y�w){U�_L�X��ʣ:��o�K��]�t4�� .�\�\�aN�Ϲ��4��.�R$�n��y�y2��<K��m�!�A�f��ܛǼ�8��*��V���T�j#��s��yR��r�Y/#��M������"�1��)����Yw(Ȏ.�����׍S뚞�ޑ'eX�Gv��C�!�~�f�\���vK��ĮP��o�i�י6�ȣ��l�̌.���q�z|q�H-9N,V�w�p���LW{������3j:�&�8��_�CD�����[}�=�)t̨r��Uռ�=�A*�u��x��[? �b�x���8Ӌ�����r��ڻܡ[D�m_���B.��ddnu^&*�dcJ�2닶�Um��Z�}��Z6� ����Kv'.�4AXΰ9=5��Tr�qvڦ�:�+�1 �<���ٟ�le�m�śH�gcsw0���HIh��LR���V�� �uZ嵟*����:�(�\�����
Ąo����ODݮ�D��d�ŌaB��7;���Lf}	F�##V�F��-d�h��1UJ36�1���U��������`���"��!A5A���S�/���L��U��I��UU)���	�^�)NJ���7b���ܫ��*%()��<���T�X������R�*��,�]�0�4�i*�C��:��࿩Z�0�����D�&����4j[�6X)�w���Fs-�l<��i%M�:ӷ�jm]SѺ5��Aydd����%Y�J��ٗ�2��	J����F]Z˖�h`�rU�@�J��)$�Y$Tn�Q����RS�b�<i$��vZ�j��>e�H�ҫ�� 0�S�!m�o�c,��y�9����*�F�R��("ۈ��3Ck��؎���q�������R&Y��㊑E�N��*�i��QT�Q`�0�)��X�툃D�*F�Z���m%UE �*,�Q��e����(�3YTA��-��n餘 ,MXXѨ��5��
��2bԵ�s3�V�U��&�V�\�+L��`��J0�6���? GĢ>�<�z]d:et��^d³�hjV�G��`dɹ ��^�W��Ofv�����Mu�Ύ����q/�`p�"ƿb8�� ��I���F:�{�*�f�>��4�q�d.�]j���N�5��@��-�\�o��^���ۤ���y�ʆ��� b��Ogf�jGa�h���St�7��s���=]�'�e5!�z���Pc�=�e���k��d\�b��R��Z��dhM�+�r":&E�zùj��<�ގ�>K������r�4�{�3
㸮{U�.-㎀k���#H�ay1�g�rL�"��,�7E�K4�js��K���vUS�F�+��}+�R���Q$�,=0�חM}rm h�s���r����t��׶��F�(�)��f����������{񋱼�Fd�[n4�Kۻ���mT{zlt\�i)�byE4�qz	�Ί��'�p��7٨��?=�s˫�9L��F𝴛ҋjN�u{�ˮD�`ݭ��K�gw� ��P�{��Y�>9}=��yLU�y��z^_Uwh�s�`w\>��!��k/�v�q�<���u�Xs�\fc<ɦ��΅b����iY��7d�95��m��j��P����u�+Q�*c��`��z�,囻ſ�V$�[ɞ��qw���{��B~�3��#�������_.�u�a���h1�T��nmj|���NݓfGݐ99��ѧ���t�?v˗9�����I�4��J�٠�T1��Yġ�U2󼗾Z��g��yR[֤>ua�{"ʭޞ*{8!��OQŵ]�@z�H����n��f�j��O��C�N�aܝ h����:Ȝ} ��j��M���m�FQ�7��n�)�,��N�V$R�c�-f��/�iWh'U�����$-�\B����/8d�\M��P7s�f]w`TmXE.�zT7��3�܌�7߾�ꔞ�4��X�p�M��Y�)��@(�Y8�gP』K�X�x�u�¨�	{��Ty�\��Ƿi��B��W ������?gF�{c�L�|=5M;cN���iga3|�>�̝0>(�P5��?Y]�jK���`�V��pz��Gqv�z�q��=�����(�~͹�WH+
-4�p�<����x�KOkٍ�>�M8y
�`tt��i�&9��]�g[�3�ʞ�\gJ43C8 �c���k�'��Q}M#��e���=��_V`��g6M�m��u���c��ن���V�G��z29�� �|�>���W��A淫��������$D�=F�UGhҾm<���nE���+����w`���w�i�{�O�ȭ�^��N��Q�A�.���:�~@�}5\�=~��������12�彎p�a������ӷ�b~د�~�b��*ۗ�yU��� �㦹ƣ�9u�prna�]t��;���4t����
�ˊ$Z��+0��ܜ秫��sh���B���a�g#�{�W�Y�y����yie��c;
��$�W9M�f��7k�c²G��`cJ���o �ի!Z&�t��g�M;�M1��ض�R�^-&�󷄚���+_z"'�	���]��o^�8����XT�mzz��t�/:�3���{�(3={���ǁ�E{��+"�T��;�p���Ru�K�{QJ��{H[�y���z�jzey�ɗ�Bl� �h.}:%_C�yJ;[7��܅P��'1�����>�e�&�J^s�۔F�@A#o�/����ۺ�Kq\�FK�1��:)�i.���z���v�UG:�ٰa��#2N8zL�ݺ��Gv+�ܻ�č�0��*m>2�N�jŗP�{�>�DA�v�����u(hzD��xBz^�HN��z;��W(�����ױQ�XNA5월�sN�5�(GY��by�n=t-p�9��S��f6s�>�cb��5³w`�_v�Z����?-oCwC��-�6��18;G8j�%�;�E��[�1��m���o7Q�OZ+r`��}�l��\M:�w�/�c!� ��Qw��j�k��r�=U�F��\��̱}QkC|�5x���W��WPq�.���5���-�q�G��p\E�X�t�r�9肼*�ZJ�yE����ET��%	u-f�v�~�զ��]�s<[��А�Iˌ�\F���:r�y��Z��M��cu�����rU�+��e��svS����g��a���	C��]r�J�/���\я�*��q���w%c���W2u��>}����	:��(�80Hҟ��K�z����Y	�#�s��0�g�g�)gc��ݨ�
��t�G<��-�����)��k�k��SM�E�͞�����^��Yu��lm������VK��0Q4��A�X��!�&!t�KS�.u9�FK"3x�A��z{��j�׌;�fe �����t�{�e�����	�22=]����gEF�؝P��<��*WP\����2��,�{�z �w]��zT��Ջ򋻽x�i��p ���G�V�F�#wg8��Oy���^�\Ba�`��V���ĕ�����R�j.�3f4�}�s�5��1�P��;�����ɺ��|�7��f�%�ƙ3#�Q��<�V-T���]E }�����c�R�y�ê�NG=�T�H5^*�(]�p��+�Ĩ��X��UV���ct��=��d��������O�꛳v�l-:�DvC ��6m�#������[4f԰m����G������GҺ�տ]��Z�m��Ϯ�R<���V�{Ht:3N��a�u�΅�ݸ�uԮ�=iw��1�a��B�ص;��>����L��\��No�-�@��\Q6�"���'S��_���cyŽv��[�y���Z�&[&�e�o�1G�(��ݚ3ۖxoh'���1V�b��n��hyQo��5)�4�9] hS�6��w}����<��]	��	�W��s^.��>i�
�k���QM§7������m��,*��m���x^t[��� v�{����	w}���M�Vr؍
�C	�kI�7+*��9���z3+r���iJ� Wc�ϻ�������Qæ�Yx�Ζ{9X�iw�q���,�n��]-o��FX�f0��m��H��,�����ʖ�4���973�׵Eh�DGVN�����k��ٻ9� ��>=I���0֖�-�ɣۆ��t���H��<�r�ۖ��
��Mq�����OJ/4��	F�-ۼN�N�ϑ�V��q��F>6(�Knus��x�]z[���lZ���y�8��*䄺�ee>���d͂*m���nӬRs��3�\_yh����j�ќ�Ƣ��n`�dM*��&Xד���Ty�W	-�؎��p���uW-氍��n�,���nwM�I:�Pm�me_Y}MS�z�A"�΋EU]���Pٰ��٭�aѡJ���"�uw��˻t��B�+�a��ae��L�*�-�j�M3�Z�cwY]Y�eӸ*�L*\.�8*��e �]P�wD�\�j�]"Z�+$M[lbx�,�)եyd�Q+2e��J�`�ҫ��PMU�9�Ԕ�<w�m��輣Tc�D�v�q��۠S���m�n�a��.�S.㣉S�#K.7tr��6R��IWy�˻�X�7x��͇+%�D�H�s�X�r�����"��$���2�P�]��]����*�Keb�e�˻�ěm��m��ֶ�cʙL���
�hT�u�f"�Kjʶˬ�V�0q�2�\�P��W(�fR�R���0����UZ+X�
ٔ�k8�&�$���7Z�"��Re�k�!�Ԩ��iVf\DX�+�\X֡bj�f&*�c�9�b5�((�*(+u�53*ֶ�h.Q�Y�aJ�b�[eEq�
#�c��7LsY�ȍ��"���%m�U����-��F,yh�u�b-�7���8�m,H�1�*9jeP��TEI$����J`��yN�S��ۛ����y��z^��*��9S��NخN_��x���������3��@w�>��.X%y���aA'���BpA�{n'pĸ.g�K5]�W$!G}d}f�mn�@�g��:=S�%_oVtQ19=�-�|�=TG�I%���?OB?r�)}��>TYy+����nE@��@p�4��v�u�}겶u���#6�i��Q-Y����^.�̇P�� /�W�u.��V���L*��!��*篳ܟ���zv�r3g8��Jaᣌm6����,w�V�P��|����dp�Ȝ��J�eD�j�F�9E�Q�:�pN�z�}G�"���t�}�<����=��o^v�T��o��4Y���Z���S���	�%9�f6+�ң��DAS/���p#,~9�C&/MܛG!�w�a���V�_Ϊ�U���g���l��4�ڶ��1P.���P8�/��� s���:۞
�)<N	z{���s�ͦ}W�����r۫+D�[�� �|P�>���vU���)��U�8yQ�P�}��6�jR�����)?y���&#�Ho������;�y^,�EvaBY��6LM���tѶKIl�V�&����}�Dֽ�/^�9��K���W %�3r�91�ָ�\��������}�K57qɔ�3^�{��9��8f2}�o>Gg�5\GwM'����#ٍ��W�i.��L��h+�twTf��%����<}^J#������e<׻ʠӻ�9��$�4�Os������=<�����sݱ�PM4�hu�*�,�b�xhK�6n W�!���q��"��n��p��a�C�!Hr�c�K�~[2ė]�}��EƟ�� �p[e.��W&� ����o��0��n�=�yH��2�l�}��9xr�|�/^�ٲ^��*�ǵz���6�[p)ԭK9�/M�C��k*�]�����{��(��:��{N��c| g"z�e��|�k�Ѯ����|c*ݐ:�����0�ʂ�Gƺ��~z�8؃n�#�sc��np�k�Mr)�Ϧ���p��"~�^�GG�us{g�SA-8J���>�'8�d����@���b�n������|Y��
.1�vq���l���ps��'����8���-n�ȗZw7���ݝ��.M��j��P�3��J�L�n�NLdI�gq����P&ÅE�O ��}Z�s[����GGr�Q�b^�f��^�!׫��6waa/{�`��Jg$�֊�յ��l6�x�\�I�wIP��oZ�t���}K��>���pxx$���L'����;r�]ח��<��4_��jҵ���U�B�̘�o����d���mc��]P�q�D=<�8����\���t�
Tζ�:�IF�}f6z����7��z*�ͬX�s��|
�,�篚�I�`ؙ5�F��<����x��� or.
s�����F��ZCr�Yׯ�2������:)�8d�$p��x��v�����G]s޲P��F,b�5���Kx��.|��ٳ��̉���ҽ[�Kڽ�/�>�F����'��	KS�.��{��L�e���hmi
����r󜽽�K��Z�ٴ��9�úZ�Vgn=v=+/v�w�۲*��*�d�<D�P�8}�4�ld�+�E� *��ii΄�@�w�w�1�L[�ZsT|s�o�Ɨ����)�pv67 ��mq'�y�Л��f����I��n^��[p?8��S�˧v�a-�d}˺�wҽ��.�%���[{�)��-2�1��Ȫ��i]7Ϸ�,��"����39�۲�6B�*�,{��P��V��L/9v^���mnV�
a���X�W�a窸zT�,��$��cTAS�>�NT"� \�z��Tp���pͫY�bbm���n��hWv����lF=����䙞 5̦�l��Or=R'�0�bןM{^����r��
�����q�fq3�B�D��B"�0v���߸�|D��y��&��P+p�}r�ۍ�=`�#��MGX0ma<S��f{�~o�i�զ���>���6YK�j�A)tf��<ӛ����x`��-�(a���\�3mH�vۦJ�6����.��oHuN���o/v��<Tv�g]�X����u��,�)�N��Q�N5}�j����^�e�|�]1���J�Y�>�/��}�6a���27Ι,�v��OJ.�K�k@�Z�a���h��n&8�Q��ξ{\#a�ɼ��QyP��j|a�����S�
l��"�>��7^�Lq���r�8Ax�,�5R�Y�u��K9Z�s_9�|�����ڌ�͍�O;x0I�7,gՒCuն'bk�ơ��v(9�Aٹل)�
��%��zd�::�w-R\U@3�$!8�ʛS��V�wI]�3��m�2�gF��M�Hk�	�'V3��o;ݍta{㽏ܫ[/6�^�������ܝ�]};��<�XE�}�)�Y9�u^�qݙ�K}��R��a��sFrt��>��t�b.^�gbGe��(�oF���E����1�xs7*����Kt�	Ԯ~Z�b={�9m�"w�rHw�_*ų�+�0��� ��b�Eue�R!��.������;�8��{�/�Dn����%����Rw���Ns�ձ���][����YB�n���]wc\��]_�Pɸ+5ՊZc޽���!V�s��G4#p��Ñ�tH��:o�R�@���2w�H��⃃>i�D��&7���znw	]����xr�^a��Y%d�rB<�˸�a�(���K��9ҙ��o*H�a�z�C�4oX�]a��4z�Z�{�3� ����h$ۡW�esG2A�7�ɇ�����%��ݦ&ζ-���ܸ�Q�X�:�|�Is/�7�s��>�Y��p���s:�3�y9vٽ�ۅ�:���Ĺ�wjz����>�#��_I�;���L��� ֝��w�џl�n=5�bXI�Ĵ�>����I�֍��#�X��E|{��>���\�v�MY@�G;�D#�d��]J���ht+'UAY\�[��ݎ�6ֲ���)����ᬶ���r��y����%��BwIϱ΍iw��}:+���6���Cy���Ӳ��m5H�*E]��Ԕ:۝�m�θ�w���S/��k�����k;r�ҕs'�O�me���<�.�7e٠��еu՟#�We ��)Mc�\��H�s�Qޫ��.��N�#�g��jJp��Mܴ2fuJE�ʝ)�����I��tSf���h��] W�����s�L����qt1Q�o��4�)1N�����3+(�Gp7Ǭ��������'��+\���al��WJ��U�8��.Uk�C�4�u�,�u
�6����hH���4=��/u�g���l"G��K�]$͏l�J��\=2�E����r���F�!i�ҹ�[����h�ӔbΗ�@��sZ[�;۾ot�.�mՖ�`�pP��wu��}�c�$Y�]�Wz��!
S����ԭ�ۂT�Y�Q ��}���;����A��c�+e5{�+����,e.�7�S�Z�+Y����R��c�։Y�r5&mt�1���GX�Z쩋f�d�s]�ѶI��k+��p�yY���d����� ����lP��ca���}�� ^<�.܊Q]X�jW��S�v8�۬˃���*k(�p��Ew
��Y�.'�4V�i+���rɈJ�%Q�D�����ܻ l����.K�H�ad�:�Z���
*jb|1�*ư��TP\E
��V�eB��E������e+�b��,e."����CN)mb ��Z��c�W�,Q-MG(fU0J �U���4a�q�k�ڔQV
��
�QҲ���GHX�.R��ʕ-�����,K��ݱֳn�IV���\mmM��-+�G7r�%j�cq*�1i���Tt���^2�5�řJ�e��T-�R.�)5j��-U�UT�F�ʕkj(�8�AiD��H��*��RĢ��C,mT�R�����Umh�nٽS"�-E��+S�(�מ���UP��`�g锥j<z�8��ܬ¥Fu�����:���Q?�p0��C�k�K�)�<�t�K˽!���^!�½��wW�f��od���z�ʖGRq�.���h�N+C��A�k3d�u7Ϥ^�E[���ּ}��f��zz�I*P�Q�Q�� lM��k�.WFE�=�uc)�z����<uY�*�4��| g��j���=�՞�U�ȬU�����(,Vڴ��[��66��Ȕ!����CA��&���U<���/r�Op�v�vg��̿p�;x�eS�|Sα6�רmƃ7O��^j�\ʦ�i��ۧY��1F�sr���Ԗ<2�Y�C�O�cIZϞ�r{�Y�`e�j�L�ْ^�}x)�sӛ���ֱ��Y���̺�=�l5pz��y���i�$�-�Pb�6*�x!�;�r�p,��mĽ����v� u�F���;��xS^��Ԭ����^ݫM���� SLC� jȜ�>ܬ��,g6�����D�Kt��}}T��3w���Q�)�[�i���Z�b��1�1�اNr#��e��I�)�����\+�d����#���4r�t��`�&/W(²��7��z�M�c��Be֪��Ԫ��#��үwRĭ�BC�FN���Q"��+��q�)XQ�F�{Mp��E�*ܾ);��nb{��{�d�����L����w�
Է�
���މ6��gzax��=�%��(�����CКc"������k�����e�(Pu֎ޝ��>s�NT�'�)52����7H�t���mC�zl�f�Q��V�2y	��{�n��j���pJ;�e��]��k:�tu�t�!�mc���Qx㠠#�P�3:���(Y#��t�V�"��^oV�f�+^�7�n
��Y�lw�������Aܫ�3&`�yԕ����Fm٭dx��U�6<�F�A�>���8�U����*�=��/M4/=�W���ګ��!wkFp�ʮ���aL�A����4���%{I.O3�z�A���W�8�#�m7�0��}2�T+�OkEu[��_gW3&oX��ĺB�<���g/�鈷C"�kuf�8c|]��u����y<��U�'Zl�>:!�k��j�[�Y���K�U����cc������ښ͑�%��Y�Vi��R%{�+�!�G����wt�w��,�X�GD3S�ފ�rk��mX׹{���Z�-�u-�BvN0c��󺺲'/pI�I�-?�NU��_����bqYu�m����w���	��!�{�z���O]Ҟ�_-�a써=E���A��a�0��f�������F���Z�U���oۡ"��]��xT';���O�.�bʔG�H��4��'�{SI^��� �fD��}wTU�kK6�b�|��u[��zq�ebJ1�����"qѸS5n��-��G��])8w3��<[��r'�x�ey��hfB�޷�zA���y<;1=�A��{v��-�B�wR��c�s)�Fy(�[��s]#��ӽ�*R�u�j>��>z}��˱.��-��y5. �o�F��>����]��:�G��m���t���j��(���c(�G/��zx��� �����A�]�b�G;�x߰�s���ȃ������R{�������X5ͥ���s-�]�݋�i���Cbr��ә�[�J;e�����FmV��4N�-��j	���R]c���l/r7�D�>��Krd�+$�9�͛7��,�ܸtB��i�r7�,�|���k)ji.`�2�ujݓB��Y�t|ر�]L������ה%dg=n��]B���7QUڱ�@ F�T��x�;Z�I=�G(|�a�ՏW>�r��Z�t�t`n6:ޓo��fWv(JN���b��������맪:/Pn�E����
�Ѻ���{N^\yڂ���;��1�d2Uim���u�`�;Z.Sک�ثt�L#�����۳X����\���x��+g1��_zmz=v.����S��LJ��1�p'�b�y0>�Y��
��ˡ����n73_m4���q�=,bZP+w���lpѽ"�L���'�d8�aڴ�Z±�g&�;/��v�h�n�n�+��	�(�ҏ���CV:.�f�#T �'�~���{�U	b���_E�o��Zي�tͅZ0�ՅۢB$�Ze��:�3��}y��Q�Q�!���S���s��($�6�c��[��k�훈�y�wҵAJ`�/H�岹��`oH���V����ˊ�E�8Dp�+�0����}~4�)��	���=#��-ѩ�o��n��E���]E�W.�H*wn1�$t�V���C��e�3����C�6��xJ�b�ʵy�n�E-}x;�s�=�c��ӞTC��-!|��q"g�������3��aF�*s��c�I�S^�]�)Gv���]�kӎz��{�fk�:Qw�@F�9^
�����.��ޡ�4�%�`�>繽b^�����D鞑���+S{"�g��<u�<�ui�¥�<�c�3{z��W�KqmH��{k�N��.�RR�u������}[��v��<�:R�0��w�-s^��U�K��ea�s��׉V�Я�c�(3U�u�3�l{;��-�4����������Vf��7�u��Jۧ:-"�?�p <�"@O[庠x�	��LW,q�)��S��|&�z�ŭ��r�i֨Dd�G�F�C��ռ�*�̮�j����K�s:&�=�;��ь�.θTGl�T-�Ry��>|y�Uo�f���Q�;]�5 1�m�V�ml\R�W���"4+t�=B�]�V����`v�~�9��/x�-K��[�Z�,+I�L-BQu��i��$D$J*����-  ����  ��څ�I$� >����y?�[tP�_�e)h��CʅlS�a�$Q�Q@D�! 7�٭�̎�	M&������Һf����YH<�\䪨 v�1`.�#\g}t�헪d���)�+]�"fՆt�}ﭭy ���{2�ex]�Ib��,J�V�`  ~I�����c� ��w ��@� ��j1	%����E9����k�lb{T��h�����̫�K�$t�  �����n��@�Q��x��,�<Y�F k��F	�%Y���i@���d!���8�{ ��4Ӕ�6`��ȁ���&�� F�`7�K:���*�� ��@�:U��d����g>�j�©� ����  hl�e��4ͮ�aM��� ��ɽ(~	L9���)��?����;'w6�HѼ!� ^�N2bk�y&�t��t�_i�)#�V�SqY&�}�%�"ۺ��"�����u^�3Ї2�;�&�Y�UP �� !���tC��h�_{V���$cd�!�!� � U���%U@��A�����D�dƘ��ɼ��HAQ�,~s ,5�" ��3fF�|��L\(� ARCR��nF��	�E�(�H;��
��@�)� �al<���w�C��@ �Îӑۀ�j���8����������s4�bl�sI�r�4RLz@L�Ε�˃�(��N��ZO�f�����UT 7���3A��IH���|��U@K�P�S�>���a�G����5&�0fi��R�K�l,�G: &���r�^��ٖ[r��dG��/�s�!�]=N��� 7�J��R'�]4,��v\ Ճ�01wA��D���[/*A��� �@ ��/���dx�~&��� ��aҚ��M���Ջ2[�B�O��S�K&��zBB��B9f���w$S�	��q�