BZh91AY&SY��(��_�py����߰����  a5�}}������UJ f� W��h *�F��  ht��*TT�� )J�� ���@��I���V��R�E
)%*��� ���w��ɀ��TU|y�+�u��z����{�i{��;��ݓӽ����x�=ѯG$�(��/G��^��i�]ۭ����+ϯ���[tmz���Y����G;V���s���ͺ,�m�{��h}�#��!
�|E�����=�T�>�w�q�˧vq�����9΍����{�n��˽�{m�F�X��Wzh�/\wJEm����/>�h�vl�.�<Wz(��{��=�]�٪{�m����^�{<"vkݝZ����9�)([� }��
Q�n��:wss��y���o{ҽ��稵���l�k�Uٻ���z���;n�u=�� }��'������[��n�T������n��x<��om]m�������< �@�U�� ��N�{�^�l�n뻵gyx���uk�WV텥ev�y[�v�8 |���}}v��vK��m�l�f�wn[�Ǫ=����N�ٞ�͹ �  yT��g@�Wf"���������������wOwq&�ǣ�pz��{�{¬ >(�罱�}5w���.�/z�M{e�{b�ޒw{/]�-����{�\�� @
�R  ��-��   (0 P�  �~�z�J�A�hɈ� � 2�OЈ���4a 2�hd )�R�*� 10� �0� 	4�h�UH�    "j�ML��&�Sڧ�)�ieyOSeQHJT�0 &L��!���?)����,�]���RV0K�/�g�I���+����c�?�
��eED@��B˃��� ?����������������9n��F8VB@���9O�V�U_��HŒ6�!�(�ݣT�H�Y��~����?��'��|�_��	�۾u��S�O�2_O�G�`��s弇�M��;���M��oy�)�.�[���������f.W�yw��b�f�򥺻_
Z�Y��v�����ٽ�pٲ|g�]7�}%�z-�N�
JN��}	��*\���>��V��������P��]*��5�|G���ѻ_p�]��t���%��o�������q뎖d�_y�,[cr���VZ~Y��w��J=��o<<u��w�^8���f-�Y0�k��:w�J����õÇ'�8=)үJyl�?//c������K�����?//m��wCr�R%��k�B�!ڔ*lB%�@��І���s+Z؄Cv�XЅ��EC!�,ކ&�*�.!�F�1���~E�V�Z�V�
���b$<R��""�s#�B���wkb�۔-��hFd12�DT?�\C��bT��|�F���ԡSb9B$��~�7���b�R���D�Z�!�!6�,��!��"ȁb����;��؁���(2"��N��\�"Ԣ�b!��׹��^�O{m����G|p��-���v}�;�nfDz����~^��C�Jg�!o֩>T��͝���;��������zr�=��F.(\=U�~�o	��\b�>��^��{{n�f��sH��ON�m��v��1����">5�k�>y
�L6�b5໘��cv�g6{"%j�^�p/*��_1�-o���ޝ�[�����_|o&b�j��ҋ~��tG������7���>��.5yz^����ŭߓ^���mw��RcO��c�m�9ަ�ym<ƞcLȈV�DA�gD
t��"#H�݈�u1�5D�6#��",Ȏ2"�1C�G�#�q�Di�ˉ��LF���z�#�����TD-T�Sn�ղ٬�s�v�Bp專�l݈9�=�Um�j>�8��ȏ/v��gC��J�q��z6�ds��FDE�DjٯNps7�l3!�ÚB�N�b�B3�թ�n|�F7��.�����vۿ��������<^\Bb*�%�n��g/-��c}�nE�ެ���)�o59P�5ۥ��F�ʚ\��uJ�6yA�v�U�S��sG�/z�'N�x��C��;���}��gC�w�����ݮ�yݯ��s��>w��<7���C�B�N<�
V���S�T��5
��	�Bq+�'�����M���r�Oap�W*��oҮ����^^Y��k�7�oǛ�6]'咩`�ז�yw��.O�}����Qj�����og��$y&�;q��ƚ�ozq�on>�lڲz߫U��x��=����g-㋎L���hzw�飸p��Z�)Wɓ�NP��Z!j/���!rM[p������yD�-�Լ�,G[z�Mc~B����2���&�D�!i���cp��n�X$!-�>-�
Ep��M�!�

lB�-lB|7����B�nЬ�ŋD+G+Q�p�m�B���X�b�B�Z��M�
�J���*�b�ɐةAM�\��rPy�b��yo��/'�ݩB���y������z�m�!r9j�}Z�$#��G֨��л9�.QCp��p�X�!�B߹	��lB���b���F�!7�V!�Zp��\��"�]�)�1V	���b����N���Z"�gڙ	�Y	��+�=Z,B�+��)�'�\��R�S���Zp���J�yly=�O��r��*�O�<���^X��֬on|�)����p�yZ�~^���_���>����%�^B����(�k�D/[�6ኑ�K�����=9��|_���Nb�����ނ�%{Ζ�ϖS������Ё�w�ڟJqzjǧt�Nq�����oU���0���k�~�/���>�DL#X�ȍG��ɺGҚ{���Ü�1?-�DD	��M���z�N9[����{�j���1����68�<�{u��_��;����;3����M�N���������2�p�v��oz��;��|rA�����tɣ��0Պ�~���kZ��8��T�������ʔ}#�;;����;�z|k�p��������8�|��B��r�h�m��L���B#)��4!0qS��Y�!R�BÜr�Cj���hB��'#�B�Z[�]M��m�)��e8�����N-4,hB`�X������GjP�Be�����8�#a��P��NG�Q--��H�q	�6�	��B��ZC�j6�Z���4!3\��sn9
�p!V�-5(k!3
՜�\���l8�е�	����hB���Bmj%���q(�Cb�=O�w��'����/[�����S�zw���|�v'���[�����yg���|�~���)Y�xt=]w�\z^=9�E�s���_��jq��v�")B�y�}��*���㦝�ݮw����ӝ��Ν�ه}��1(CMJbmk�Qx���sbb�ϟp�����4�R��ykz~�p���</���fk��v�^������B�>[������T����!KBԽ~qji��b<�j�~Z������y���=.5g1R�\8�v�B��|E��Ѽ�Vr�7�F��7��FFa�D)Y��ԗDA�k�pDD�[��!��1��1e��;�{�~��/s�ӧ;�o{m�b#�G�\F?FD_TDv����o���i�DGd8�s�����9��Ȃf ��'�e�E�6-.#a���Ӣ;�9�,�qv�Kާ>}��y��~϶�b�t���u���+Kq|�fk���nLAn�q��g1R�pݶ��"F3]�T���l3��Î���qZ�5c�9ک��)�7/���"3����;�;����X���WNqK9�<9Ə��8�u�Sl5�k�=�=�=��;�g�X�����a���{���>��ߛ�ѽ>�8��ŭy��5��|>�j�k��d=W���	���b���O8��G�R)�Z6���&���c�b���YOv���
{�.D1�q���)�p!�#y���)@�)���8��b��&k�BH�T�>b���B�	�1
�p!�
����|C�
Jp!a��\r�N8���츴*1��@�X�GG�8��p�T���ϔ�m����ԩ>b��B�r�O������B��!��h�q��)�qhTc�m1A.��q�|S�
Mp!g5J�����5�s��S�>�ݨb)�+:#�����D8�y�Z=SV7*�T��#��-pqkQy-St�t���N1�j�b���ږ&�>��I�§'�o
<�ɜm(��حQ���b�|�w8�W:��z���LF<s��n�аȍ��1r/\j� ��l��#[z�m>gڲ�D<V؈x���
t��"!j�hm�|���}�F��G9�*>ͣ�}�w��m��w����yGq�����ǵ�kT}�bdB�p(."K���3]�E�3��y��XV�շ�������o9N��7
�lDFDD�I�vlFFH㾖�7L�[k��K��w$�ᚶ���^_��U(|�~:��\��	�h������O�C��~��SI���W�g��m4I%����u�Ϊ����_�?5�r.ݶ#�ӻ1��>qx�D�M���g���]�����^�;�3U!�>�6�{k��E��߅��f�����b���\�2�3'(#s���_������0�ٹ�g��~���gd�&7���M��LS���\YN�i����8=u�d�ˮ�7g*�l�*�wג�˒gqF�ѡ?{>�߲YЭ�:��g�XϢ�f����[���¸�eP��mf�������r~�{=r��=���O;7ə�$��������U���9����<gM�}<���k
F��Nw~�?7�~��4�~����\ƽ�۞X�!�}4˝��O�g�^���;��F�m��W�}�!9��k;�!�&��Q���~��~E��������$�&zV��w~�w�cM��v.���M�r�Wx�������36=�&Kmv[z���ɘ\��׽�}��|��5���~��S�{�~��q��j
��[Oiq��u��i�:�y��!:cvgr}���ɻ.d��`��<��{߽�����z{�.�lX��E����߾��'b�|mgK'�nS'��<���y���<EwUC�fZ�ڷt�S���V��U���l7�ϲ;�$�����w-���[�ɧz�:�o���m�h��z�ufչݵ�-�5�8ܷ��ｻ���L��/��'��k:N�;B�d���z��UYw�l�s�DfEw(���(���_��}qw{r=�K{�tû���r�iDj�!]����Q9���;a���5��y��Ku~�:�lKp�3�~���Y�^b��|re�\�R�N�<���Ō��y��V˖�w70�c�뜙tN�ݜ�ܬVl���ku[91��ۮ�f.�n9�_��2�>����v�5�>���U�+b��B�QX�K7$���rLa%�x���pے���z-i�6��� L�5���س�������6��sğ�,�5��l��;f-�?w�7����;���/�ٳ�/��5e���p���CXJ*7�����k=�?7G�������<\�YOo\�=A�^���E)����lr�Xf϶��>��Z�ߩ���2�����~kΨ�D�����r[�nI��+���݄"��I��F��l��+ʘ�&��l��+em�C�����[������q��E�c��gٓ~���L�G���{?eʌ�w��͎�Wsj!x�ܧ��Զ[^��_����vb��;�s�l�t1{~�k����
@�/C0��|.s�Ļ 3��6�m}=�oz=]2}�=�:L�س�72u}����]��kzg�	���t܍�^s��"2}�N9�]1��,6�y�����5\s��}jS0��*#ǃ�l���؝s��$S��_�E6e������Wq1��q�?�\�먝U��+�X��#y���ո�[�^c�lE�vw5�����2�<n�
$�\�Ҷ�&���m��2&.cS�b�b�o�ĳ�/��r��<�fI'�a|Mޣ�}�E�08���iӛ�pB�͕��|ly�t_]+�L���]Q>Y����$������<�7q_Ss%���usS;�X���ʬ.(e�^��>3y[�7]�6NN�K����;�J�{b���^id���a�����ͪ���P����m(/�\Y.��ѣ��$��]����#��ff<-�}�ǟ�Q���wu�׶��_ѩ�n5���٠}2,ې��Y{0L[����uuu�o6U\��xv�ΊJ��>ūUӷ�msr4�֯m��k��J=w���+��o���xO%�}��&)��;_�nQ;uC.C��Ŏo㺵os�˅_z5-��~x���~͖-��U\�_׻B#Of*��R�ٓq��B[�j�F�)8.��ސ�Vu��� �Ν������~�XZ�W{�����Ŋ,�f_ڟ���0�.����K�ݒ��e�8���uc$d�ܙ��A��/��G��݆��l#>���7��4���i���v�L5���?f>��Nۙ�<fd���vw�d�Xi��-s������gg{���>�{Y&{}�~�6��Qs�n��~�$gK�뻝�}�.z���y�<�㛚6�����zK�����I隬���Λ>y�������oX��>�^�Wx۲��ȇ�E��K:�5&T;��%֥�ǯ�^���;|����{�ǌ?�w�v�%2�ѵ&�Frh�ܘ3��/���t<�*{ճ���ҶӞ���y9n����y�:IQZ��0�J��o���fm:�\�`q̘ipS.��KQn�YC�c#�O�>��8r��+���̒�1Z��Wl�zwU(��}�2��oe����wyE���.o�~�3/}��L����h�v��:U�f���3h�о�&-{�73f`��;{�jYq�����Y�,�}C�{�"�5#9^g���Sl��d0d���Og�O��N2����r��_h��̵w�C���|����B�<j�=Fꬳ2b�W?nI���tkD��{����1z8/?z�P5����dֵ��)rf]�N�r=92f���sq�Ei41e�(�2����[�g�P�3''�+���4=!_ݞX�9�92f��ui��w0F{߽��څ��T�T)��D˾�U�bYYz���9�X��Ol�
�Y�>��c���_��o>�^G��z#k�g&b���>��7��g>ޘ����ʽ���3�fN:��'��k:}~~����˗��[�R���o�!��ޫW�O�~��e?v8�L2�G/L��~��������U]7�mz��~	vw���}
��~�d�'���_�E�Nv��q+7��ݽ�u���e] '7zn���ʒ�6v{o��>��f���d2���4ɓ7L�Q�����B��wd�5c�,���{"�}�0YW{��od	��U����=�[\��j{��l��;�uj��n�����y{Y+�fe	�t�u���7Epl���#�#����q�S7���0�>�l�3��1�����޳u[��e��^�|��}��SN���z�foxnw���˭i�]�o|שf�D(�z�ƽv�L�ٍ_�u�����2C�{	d����W�����~k�M����bj��:o\��~�\�{f@�٣̛����lֶV)�l��{]�#R���i�f��l�����U�V����Nj����3�r����e��1��Ld?N��Z��l}��0/��t��[�������/�/Y��m��(�j�����+i��Ӷɿw����?:��{;�C��g�aD�S+ٱ]��b���찫0�W�v�1A���f�M���vm�]{~��V��e�����>͐�%�yy�λ�����D)ͺm�&��y�Z��ڦ����7��sUH��\S+N��4���Yٻp�i�Nʉ��t��eN��6�P�c'3�|l)����2��m��vOL6�O]��f�⁆�U}���{���s�od݇���>����'c����0��UP�nQ��"r��s3d?vw�ܞ��?K>���~���܏ӛ�܇G��C	��3߷�O|��,̇�ogN�빛ej㗱-{�מu�m�OM�_��w�����HϬ�%���*��Z��޻pʽqy������";���<����0nɏ������׳1X���ɓ�g��ocr�c�����k{b��{9�fOu�w.�(ح�,3�[�w3�ݴ�SY3�i��rWwf'���`7��v��ڜ�*����s�#�n���R�.p�Qu�M�ɛ��}kO�wƏ.�X�:^��N���IHy�T(n�Δ�3�~>�{���_�y�S:�:Jެ���t���nr�uGن�"�\��O�������뇶c���Ԓd�ҟ�~�_�����?�W�-8O��������~���X?�I^A����R�o����Wt��xB.:����*�NU\�#R)�F&T:e�!�to�>w�~%���lgi,m6��^'j(��pc���f&��f;Y���p��YdF�:b�qI%�{�}��vۙb�vBm��H�1h5��7ckX�a�g9ҷi�ѥ��\ۭ_���{C
a6��锣=�s[�!�G�C}��[{ðI��^����-�76��U+�Z��J>���
�yٳ�i`☳T�tkٺ�s��n�==���a����b�_,�S(��eǅ�Ė6�mh�m�Bfݒ~�d��.4�hY�5M��hb��khQV#���P��Fg#��{laHc����z�L���$�*�"�Ws�L���l���$���Ḗ�ֱwT�W�f�O��2I�ݯ[u�
�a��9�_Ӕ��>7��!=����:�[%�-�.lf�κH'K[DTm���0+T�V�����km&ҋ�֪KS1�ct��[4�F��s��9�e/M�dֳHŘ�,�QK&WQP��9�q��A5k������1I��f��)�ˡ��&أ��W��ϋ���X3%�y�����i:��Us6��E �1i�zw�=^���!zмrZʴ�3��j(Y���57�6�t�%f��LM1H$sw�+��JKa���lt�4s��;h9�2��Ԑ��u�XWK[#P��,� �2�m[T�њ�[I���.��x�,���7Q?1��B��
��*�C)[���k�kr�G�^�x�� �b
�q�b�;ޤo!�IeIXbu�����!�uͥ��I%�!�5ӗi��\��,#��4ae����P�`&���Y[�Z;|Y�Ć��H��HYW���|C�h�ќC�m��9GTfq ������ܲ���UU[#�G:5io<Xd��*�b�5��m�ɖJ�`����Rzޓ輘��ٻ.Q�w���,|ʌxbcr!B�b��/.�qX�eVX��v0 ��h.�}�`�r���X�Ibڕ�j�"��,���9*2�G�G��u��M����R�
H��"�[�+ĄEh)"|�Q�ċ�{ú��]���2�N+}l1f1Z'Pؚ�o �4	�2�$o�,uf85����2!vI\�������'[ّ�2/gǴY��nY�X����ީkl4��X߻�{Ɖ���C�"�<����a+��2�N���NS��Z�3$O»dMiC6n��� N�eqY���uѐ��5�7Yջf߽�"a��n�ƒ�-���bI��J(�b�b����w;}�(~��l���"(���_H}�ˊ�?!�_���������o�?����������A%(���/����~��n� H `@�H ` � \� `       � 0 � �  ` ��8` B 
 , ��$ 0@ ` P`` � ڪ���  Ѐ 0	 ( ��T���$��+*�#���E$����%BIQB#(�hET��$iVU�-��HQ��Ȥ�6�# D�h��6hl�h `     p� 4 @� p$  �     �  @  ,�� 4@  C� `   �  h@@��v�@     � h@ O�K����KP�ɴ,X��"��� � ��l��"�"զ�M"�[	U"�
����ȍY�ĕP["�$�-�ff`���       �  @  ,�$ 0 ,�
 ,@�4�� �   �  Ѐ�  �   �  �HX�    0 0	�d�   �  h�3331���Ў��*��R�؂�E��R# I1	RDd<e@����H������i)}�j}�x����      �  �  Ѐ 0	  8` ` @ ` @HX�0  ��P�  �  0 �
  �	p@  UUP  �� ( �   ��|���!YFE�J  �,�P� Q+	Xx�q�5�U-D���ZE���%�I�HuC����I�j��ȡDE�G�AM0��*B�
��a*Ld+�S,+ P���1�_���A�j��'������������t??���?i�K?i���~��f�6p��4p�t��c��z�1��i�1X�4�Lc�1�1����6�1��co�v����m�lcm���|��1���>c��|��cn��c�m0�1�c�c;clS�X�1���ھc�ϟ1�������6�0�+���>|�1��0�+b��v�lcܷ��ͷݿ6Ǐ[|��x���^6��o����6�>c��=cLc6����_�1�1�x�>ccc�x�c�a�08��:C|ف���O�ͺ�:��%�[t�mv�Ŷ�9��b-(����a���;�B�_����d �Dے�B4������T��c�TKc�T
N�+'6QX�	!�h��{����'GJ�Y����*c�̜�I o���6������D��yC`����U#Y�&���j_��hY�f��$`Vm��K��޾����%��39�݇ftade�����}=g�W[�2�
J���d�¦ضh�Z8,��H���V���)ͮW4�m&�Ƞ�w��L�B�D�֙�O�!��_���ᘛk]X�M+vIf����d�Wr��fl��3!\0Ʋ������R��e�⮴�U�%�Z��`�B\�m�Z�v�A��SV0��#�ȚZ��4Ib���i��n��FxY/�gU�턢m5�k�oc5�1���mlHC^�o7Z��k+5n4��ےhM}[���r[�e]7�-�{WIp�3%�=4�MOzW�u}=6��cD�m��M�5F�����ID�M5�F��]��L#!]����%��mu�%�OZ��;��k��}���^Y3o$6�I
ÌDu�m�K��vI!7���[�,����D�ka�8�_Z�Ġ�D�y:��׏8�!��m��)iKh�VjD�H�#�>K�w>���{�   *������� p0 UUG���� �`  ���/�K�� �`fo���}��pI �>q�8��N4�J�cӦ;c���O?��0>�Q��ZEba$(�I��AI�h6ͮ���BׯHV���R�_#D��	�s��숑�խRݢ3-V�f���_Ѧ��Mu�U���&��^��d[p�l��ME�pY[
N�L��V���]ȍ� �OQSgќ�z�lE���Ѳ�I�x���R��4�$��Ͼd?#��5EBJ���}��G�s����[e%�~Z%������:��Ta�+��j^���!�۽2?�*J�gS�Q�*�n�)��M��k�C������6�3jX�G���jX%��-���{<�I>�g'>��a��	'�2H�QTS�G��0p��n��cJ��ct�4��xS�&�� 跊K[�%�>mUP��59�:��<9��pJ:��!��U<ٳ鷵�cQ���g�� �d؏�<���n����(�*�������s&�pj���/��6�(�`�3$�NG����3"�˖�S0�<7t{�eHD��#�l�b�|���x!�����S�Nۗ0���=z��ƞ;v�O�|Ҹp�+�ݱ���BS�!~�>A}V;��"� ��Ѧ�Y�$0prB9��N����(��L��\̧2<7�}��}I��h2�[N��9.-$�\�)b�԰��3l����l�2l�ޝ33�B}�`�!��}(d��GT�\�\N��L����j�pb����,�9��e�FF�%ko�n:m�4�1�cc�liۥx�����?���)k�� I���s�zl�o���syW�i�a��K��� �KuiڰZ��d\8،��ȎI&9�ۏw���s��6��4x	��C�:m
Ԭ3��|M�cb�[G!�c��n�E�E&�U�:�����~Oa��l��u��nk�X��h<��V������_omH�˪�Zs�8M�1&�R�x�o�6��Æ1X�G�~	�� �)8�կ��.ǗV���͵���('�̍�Ν���py��J��B�'��)���>}���	��Mw����ѵ�k��V�m7��)s"v��P9�����$��f%�)SC⹎��MJ"�YV���n�}�� 	\,��jƝh ��)C��Gb�*�W�����pm�&c�f�0T�GLM������'6��j���چ�u�ix��Κ����m`��z�rČ<:>�-��k����5�h��|)CS�Xz{����'C���ѭij�F1)B�`|x���A�Ǣ8�ۮ�m}=��R�l���!��ߟ]���d&o̓'p`�L�4Y�V�+�خ�+ǎ�m����ms�Z���JS�UT=,~%�ӥ�m8�o�*�O�rC�7���%&N���j]�m q�&������l���{)h�>͜���'���S	u�&e��e�����Ƅ��棉��%�/��ѣ}a��!�����V�m���{(zh�a0K�)B��it�r3�o_=v��֜i[8c�?
~��1�Im	Q]�Ua���?��0�t�e����OE�b��xS��2C|��-�M�A<�t�=��C�����Ʈe����Kmh�l�ъ��������<x��8%��gW�yw�j�2a�p���͚g�Fڳg�f�D5��٣���s�T��r�,�,>��г�j��>�v��Ǯ�i����1�"�bUD,X�������q��`�Hz���� k�J���	�^>���}�1u�F�`U���!,!,�����w�,=�;��J�T��9:�����d�se���h4x�#1-���S�������eip�,��;�Ni1��>Ð�Hn#������o�Q맯^��֘Ҹp�+鎘���i�[��TAEc_{hYk��A�[R�NB�4M2��Q9�H�D���&��8�)XJ*9Ib�����-��JHf��VS�=2_x���m��?<yB�z������ ೘�Xՠܬ���J,6M���HZIЅ��b��� eB�cn�Q�D4G�c�u�J�3,Q>7?�a�7<�<=�Xf��(��0�w��'���PN�3��I���Rd2d�_C�T�dԳq0�355���z�j4��9�|�"�<�rta�p`�5':z���J��!����
`v�W�sp�ffW7#2�[q�4��aD�L�+e�^=)C�8�z���!�V��ҝ6h�Ҿq\8�+�xt�^<t�u?��EިV9WīP�1UP��Ҝ9C�}9fD��=84�4It�CG�ߡm�QE�||z��^��&Sm%&SN�vw:��*���	�6������s�%<�,^���G�7�ɣ�a��ٶMc�u-�<tv��i�9N����H�(������>j�urj�,n�������:-��/��Z�9O&FF�m���V4�궳��V�k�qv�����5q�4�N5W��ǥ���|WӦtzt��^�����t�M�;W���:=U����|ӵ��[��\\_�v�/��Uv�+j�v��_���j�^+���)᲎��_�<��~i��6�������W�Z�z^�5����\Wk���v�.:zfA:'J_��pz'G��z?�8at!��F+�����\cUƸ�^/�ǍqƸ��N���=������GõO���ѽ��Õ�^�_�������~��=�8;	�:��h�N�螎Ζtpz?*lh�X��\]���n��.8׭j��z'L/Nץ���~;W�����N�U6t����S����Q��Q�z�W�bx'��1����;����ng�ζ���g�^e����݂y^��ؼ�{��i������]��;l�A�㸬Ý��෦w)�ܾ��NC�y��z�{ʑ��vZ���x���qP>,��Od��K$�m�d��du���14sO�U�Q-����ou_���ş{�d̮f~���I�߾�'b���Zԧs؟#M�^�;������wZ8����N�%��>W��O��ŋ���9�l֛�{���oݯ����{�}>�� p�&fO6��仺;��ǻ��{���D32y/�]����i�z}�{���fd���wt�w{����{�����=�����t�M��1��:c�����|<B��btS�EEED��S�Ѩܦ,*���sW^�G��`�R�ȧq�H�)� ��"��`���tZ��Y�Ԋ��aғ�ڝ�y�Z���@e���5���_�7R���	��j;M|���iEV���]b4R噋C�;�����p�t�޹����,�W
��jjI��k��jrYҽU*M�1Cޤ� l���6@�A0�,�bg.e5!�YeC��bX� s��,4D�L�b`ISrU{I��@��ȶ@�y��)�A��e�ƍ�)gM<m㶜~~W6�e>0��t�Л0��EF)�x[Kim-�'"�̀�t^�u�2� ��$(]Z�a��R�:ϡΫ�N�~�쩕iouut�Ma��m���M|�d�a�w^ v�n5��������ܭ���5��ɇ����� ~>TN֕C���u��̄P��R� Z@��462}?~V�C$3ؾ5eJ�U��;4��S�Dl��җ�/��R�L�ےX�Bć>�� �0�@� �E�-�a�I���E0�AP�Eh�y q"���J-J[<Ri�o^;i��+�0Ѕ(R�iZ��j�X�z!#zj���& *82�7,Y-�k�@��ʹ�<B�K=�{W>\QWmON%����0�̌����X���LxjJGᷤ{ƞa��yƳ�z�q�	��.�%�̵��%Kn7,&'h���3u�e�m��r�:j�����$|�k{pz��}��!OR�DSl��;H����)fN*#�z`�aN��HI���k���тF0
"� o�II<G	�N;h�$�ɣŏJk�4���kD�H`�`B'�.P�����@��z�4�2E��3����2n�$�%�H"�~�R��e?�jC�+Ց�Q�'a���C��N�44�Nfd�M--.�u�c6خ[�`2�ID����-��
4P9,:x�nSز=���M=U4�v!i&e m }� �۲P�U��OX����cƘ�<Ǐ�(���#��e<o���UEH�R)��`�2��=<F��H~�X��f�ٱti"8�d `�Y�"5�HP� ��)�d�x�(�.��R��)Ām6�I���m!a0N0rD,���0m�{z��b��/�D8T�N�K"T:^�/%/�m"�`f.�9%a�P	���'��T�d#��"��]j�xeA�����2C�6X
=�(7��g&�XC�	�I'C���"�嚇9M�\��?5MBy��s��2��c� �"�X�D���NMP�W�Wiy�%
6`ɃE�i�+���c�1�۷�4��?$�פּ��[h�,�V,<k)�R�[KiA	�`nD9I���`t����`,~��89)E��J5�63��x�:E���/��UU%���I��L���e�.��2hO�<1ɩP����M��a��I�>�}:0(!�>n�gڷ�:k:un�]ѓ	L@ژ���dENDP����W�E�1~HH�Hl���шٔ(�H���ū[sUE���!�.B Be �-�v��J;)�r֤YO�������������C$=�>b���l��*�5v~�ԏ��,F#�4�"�Ca (�Hm),`�ae��6E�=1_?��~?�1�cLxv�ۍ:z�N�WB�ĔEj�k�L�c��(���E>����[JQ����,0��$;�b��D�`�FR'�:�ɦ�����凷��N�$tT`HFK+.�;�KՓ�Ō�]�O�f�Y��^/JH�v�v)ċ��&�+���I(n'�.���K�.�˹krGeB�
g�[�qZ�eg(ܪ�;W��%:�jM��L��Nڍ4������)�B�SeF�(!푂J;)�CC�!(n'$`��`���܄�H������Ԕs��Y�F$C�i2}�в�)2qZzXr|��J�dw�,H|�|D��o���ÞU���N)��|Ǐ�������V1�1���j㧮�t����n{`�>�^�H�m1���@�(C�w���\V>�u��k���u�u��-l���h��V��|#m�%���ŕ>�e>�V��Ԯ��,�K�<�a�d��sj2�ĐCi�t!v�H����u��m��i	=�vvIRt�ݙ��5��%d5�&��/!��/AP�X�6�����@�d z�Y
C��l�m�z'�%9aa�=L�*P@=,��wTI�Λ��O����ۮх�@Ϧ>����2oM�e����2V;JT�����Ux��S���Z7�	�'g�*@��h�t�"�b�>8����==�Tb���`�؇e(|$>�KL:�I�F}�*8�t|KP�{]�qUm�U	Pw���lX�*�^��ja� p�:��y�zBC�۳%��
`�5`)F��40�߬m�A��L�"z폕�6����1�1��WM�:Tn�e�j�ְ��J߽��}��-����碴5��
�Å�	�30OD9�[!��|nf,~��V2)��5YڝڞL��s%Ux�D�ލ�r�$$�D�"�٤ᇄ!ԧnM�dF�y
BL�i��G���"l����xq:������~����cDH�7��4m���Zx.LJ�)��VY%�t�/��/U���B!���d<�ҕ��y'�~����
5,`ɨ�ז�\0�����jBB]�@��[��.J�{L��� im>^�,�t[Kv���iƜi_�1��:c�<*�/�U^\�&x���Ӻ��4�-���	�`�?~��pO=��a(~�I�d�N�K4���x�1f�m�i3$f���"R������8iF��խ��lpB���}�Ta`0#m�,i�ZT�KXF�u�͔��|�:i�H��p��擥�ݤ�r�ݓ�nª]�S!�$JO�va�C�	���l�<�\5�p���|H�a��Rx��M�9&�D�:ᣡ�CIF��}��.�~�ҡwM� t 4��/�����=!�f͙8Q�!��A4!
�Rj�&�yb�߼ǻSJ����B�g��'�χ���1�`�&w%'�3'��p���8��rC� ���m�CJ{i�%e8>����P�����sZ�$sk�������u؛�������=#����eti8�h����lLd�Iy��*J��F\�)r
���:R�CA�{����G�w
���W\���覙����~��7��O��Ծ�;��r��B�	����	�Ή-!�����:�i��5*�.�6<)4�x�0M�4���E��� ~��i��Ƨ��������t�����}/�b`�4w��/G����i��t��/k��<�:S��t�z'��:l�����z�V[���r�jb��/���g���qv�v����q\^.����ZW�n�1�h��x��k��͸�n4��v���[i�������������:^�����~�J�A��z3�G���z'�Jtz;^����uũ����z;�>8_�~:_�;1�z=0�^6���qq�\^8ۯU��^)�:3GD�_
tv=��:p��\t��j�8֛ռ\^+j��x�+��z>����=Bm^����N���x�W��W��:8?���zj�/G��~>/G�æi��S���ø��gK��ʽG�
l�M�.�hpz(��^���D�?E/J��0J~)x}����0��c��U�|Fn�5�����E��߱;O��D]����u�;�}��;,|�z���ݸ�1a6)��6��6س-��Y����n��U�2f�b�]��խlY٥�=��Ǟ~C֚u�5l��s;UPO�5LV���s\RH�F}�u+�����k'UPU|�z�\Ɩ�k���5dZEVZ�0�\���6=ض��F�퀾�����m��Ẫ��!6����˞���0��[:|��R1k�#����"��I�ˢ�ݍ�k�1Ծs��U��a6�Q��I�� Vp�1DS��b�j,z�M٣2���r���vc�G{t}�L;x��L�l5:�u���ɒ_V�[l�+4MaXr(n��7MuAB��눋C{\�gآ�d1�eoS�פL>ŹN8��*t�S_r�f���s<����QЬ2�c^���qP~���/Io��\V��MvKv�2Lmy�No�����|���&2z�,��-�ߩ�}Av�w=ܶ�����ɭ4�V�we�3�D�-���a��[��L�Z��q|3Θñk��VGَ��bv��v-�qKʆi;UE�ƭ��6݆��]�Z�'��C[��[t�PbtYE�*<깃�hIM�:kf�����y��[d']�PّWU|���.�0M���4aNT��LZ\[H����W��-V�n+����$����$3�,U�Y�a^~���=l���ե��{z}}*S[j�b�T��R0����T*�1�@����P�䊪�FMe&ƙuH�Mj�/|���*���P�̅��/�h�;�ߘ�{��/{ޙ�<�wt�w{� ��^��33�K������ � �ޏ{�3>ϻ����ް	 {޺������.\�Z��m�q�1X�4�n��t��^Hk\P8��[�+�5ܙ�G�9h�K,��G!`�����E^���:\H�I���uԮ��o��osk,���ݣ��m���r�>�֛h(�26��k��愅�k��n�%�V��-u���5;̜�ӄv�#�)��1��$f�\>,�I5���f��S9���+5$*%����N&�'h�E+�ɹ2�H��s	i��I������"L�%q2Za.��6�[}�5P�UCHa<N\'vS�9�c��椵���[k;�}xt捐�E:�-���I:�Ô�֘�
0�8�9j&��z�2�/Ȃ�Oc%<!�ғ������Ҫ����^U�l��-��u�њ��IHJ�a�*�ӂ�;����l���$4F�/�i(��C�UTl���Yұ�X��|�c�V1�R�j�V�5+��^qL��W_U�kZֵ(0�����<�� �d�p>Ee�*�\���F$p������x�7e��L�GœX�\$d�L��E�R��6e2:8�}�O��A �&\'�]�[�������Oc��:Q��ت�=�&���,�p�v%��g�ʒ541�RN�lbt�1
3��ӽ�^���e�gĚ�>���w�ݴ��s?iU7$������-l cv���Kf����d�@J������*e�@���7V�G�%؝6h�F���N\~8ⱎ��+�j�ǭv���$ 3��v�i�OL1���޶��}kZֵ(�"���K#?H�D�����L���\eW���:D�Զ�|���a��d�p��!�B��U,�FL�9N>i/e$��l�
�$cPM!/?�~q'��/�핬�<ɤ��t��-�feAQ3#Q7x�r�y&�$3UuwY^�!�i�?����x4gg��]-�1&�h�0��o���R��t�;I����4��I-1�N��!Ё�nXQ�6������q�ʬ;g�e<�f�N������>���������cI�C�&hѓE�<t���p�q��1�ۥx��LW���N��z��kZԠ�K�K0a���2u�ؘ�������"�4���u0�9���v�^���+-���}l&E̖1]��;�����d�m�x���q��Q�9>X���-�N�,��XY��n���c^��?(�mL����L����Jp�#"��{�S!&p�[O!Ӹ2i�p td�aN����=7E���C`�u9ia�%��,��n��@�s�0E&@�$��Dƈ�͔�iF)wrK8�;O�:��i�%�˨��|�۷l~q�W�W0�����<:l�/7pЉ�����ґ�H��8fp� m�u��)	,3U�y���>�G�K\)1n8%�1�s��}���-���M�b��Y�Ƈ�EE%9jpNE�C3�	j�5X��,.�QR�7b78k�m[��H�QT�3.B��1F�m(��0B}I�5�����!\4��+����		=�����[`�G�L�����
H�!2I�׉E�m��H���q"K��\KHz2<1��i�N�@���V���>�O�@�;�a6㍟�
"D��-)l�&�zfH`��Չ�=�Y��@�MX�!G�N�Q!����E��8M%���+&�<�8����A�"hpR�L:0jE9��{���!��^&	�Z�3�L��0cG�O�DT]y�[�٩vaiF�Sl/)���IA�2<f�XZ@�'�JHz,�Tj^d+�����v�Ε��~?q\b����!b��wqф< JY4|kZֵ(0�8a�a�f�
�=,����K'�����}��-n\��|0�jvɲm�v9�Ju���8��T�cnIK"h�Fݝ�U��A=��i���*M��iޢ�	)��"�!��U@�B�ں�M��!l��Ű,�A7;���QKE���Xz����iD�o���%�FXY+/&￲�%4|�<�i0�SX���J��?UjY,�N��}�0e�I�?_y�h�/��/V��~�����ƺ�7��(�$<��R+�>q��?4�Ҹ�q�q�K��!b�QSF�AZ���:ֵ�jQ Q�������^�kiM@Ѕj3�	�Ƀ�!;~p�!ǀ�����u!y�aGݢ�17��*����K�hP>�C�CϾ�����֫t�e��������
�����}��>�JIl2�2BL6` YDͯX�>�)w<�����kmk�Xp�ӡ�\��ܥ1�J:���SG;�G�B��y<[*�Z�'�ř[�p�h u�F�u�%'�b��;MJ��C��9�A�<��k�E�ՙ�M#
2Y��(�D><:'N�pÇ����5��ZMm�a̔cԣʿC1�cć�L�a�ҢՖ���Fb��� x��L������c�42��O�Cs���ޔnex��nI�1Xpyld��K0�k�����CF}i����%O�C���BX��1rx�I�(�L%�Pu����"�n�
���><R�CI�I�ueܢ�Ve9�Rq�!��ς)VPc	I`�L%���ҪW�.�Pd y��X�||�#�|��Md"�A#��R1�P���!������?A
�0���a�m*�'
5@5*�<t�?:~i�+����/����e�[���e��H�H�i2.[��䞧�(���o:0�rev���9 '�#��+v-��V�}o_��ؕp����ͱT�뵺[6ƚ�L3Wi���,g=66��f��&�I!L�ĚY;t��R
!Bn+����1�bhKUڴ����X��$��c+g3��l�d/3K��yrm�Rh��!K�����F�N�ŭK��$��I<v4�r���!�bHF���M6�` t�!�қߝQ� Μc�P�Мy�N��
F6iM��I��tq	I�izM����I�D���h�/j�g��#6�YG���=8���5�DK�����!AA�B�~5<��*�)A����������d�D�願Q�T����eְ֣���l�C!�3��y<8y(�t�b#7�0���b����{���;�>~
.?+����1��W�{��wֺ�:%*��'�1�eJ��v����E��I):�)f�Ĥ��E%�
6İ��	�Ӊ��S�n�&�FBɻpq:!��S���/4���!I��
�P`"��N�_'�.�+	�I�����P@��e)6G/�#!u�;	S�*�]�esbdx�2�Yd������R%m�䤧�����B�.�lCd���,�å���j��+û�)z[-:)e��F�����O$5A4~�Q=?~.�`�����γ�gg�;gKÒjkQT�,�W����j�q_/���W�q|�Nץ:l��O��}:^�N��e��=z=�t��M)�f�W�뚷���mX�[�1X��.�qg�=_��|�]��8��z����cN+ݮ���mg����=���'O��<��4Ӆ��x�^;q���qx�Lx������Ǌ�K'��`�G��:'G��~W��<���|a��x�V./կ���qƜx������zp�poG�΍�h��-�މ���Wgj����:p�Z��Lq�ץ��\��L_ˊ��+�}��6>�x��MT�Ή�e��
|R�gG��u��x_���z=9^�G��/N����;:^�NW�NG�
wզΗbx&b��:UFtQ:	�G��UG���.|w����������עo�7LQ�8ĳwo5��U��������_��j�޵�˓��ݼ�ϽWk�����s�_JK���!��=��G�1z��=s:�t����v�{���/zh�~O�Z��#M7�W֘�j5WE'=:��ؽj2��~&n��Z�>�d�������� � �`z�ֻ����ް	 ���}�����P��U^������ޠ��u^�=W��nݾx�n�i\p��8a��тx��v��a��Zֵ�AG�P�d�� ������m�g��bx�%��0���!���r����t|,8S��ާO�Α'ϒ׬0^��x�I�<r|���%8���a��O����,jY%��1�XY���9>b�(gΘJ��ِkd��Tŝ)���S��W�5�<A7�
�^�Y�
��L��Osea�=Nx�� �"�T���%����O@�ɀ��`y0\2t��i<�@�Ui�u��ɡ�i$�C�ɨ�Y�8�O_1�:i�+�Î8�N<<���1���
��
X��i!��~TTTW���Ӄ�ؚa|-�.���(�dO���B`���Ul���&�'�	�Ϣ1��!�r��\~�-�65-܄'��q'��!�1!dD�=)|`�Y����-��'�UUg���`��M������d��1]
홙�[3�Xn���Dvd�4|u��$BS%�p�=	#��hك�i�)��IQ�1 �x�Ĳ���B��(�<;m�Q�����R���W�`z�A����Diih���%��-��q�4��8�8��<:x��{�������E^��)ꔯ&H
1�F*�Vemb���0,�E&*�'�&�>:;V�DC���nYn�SٓX��2�\e���-t� H�n���`!��4%��R��P�M�9,Yc�nt�RjM�޵�(�J�\�r�6����g�Yv�%]?��"����HJ�u0Њ=*����R��N�3df�m�\BH1�c�4�6RB%Ü)p4��J0<w`��5��'>�Mţ�a7���a0��>Jr�ҋ}�����e�H�x"}�L%�iYHq֍�g���apt9i�v���!��A2M��,�Β���	%.B#��K�Iʪ�̽3��:<�6R}�ב	ey2�)��:�Rg�|�Ӟ��H?'�������Ƶ��V�R��I)-r�w������dO�~$e��yA���!fB�Qi���䁶&�H��K��앧�<v���~z�O��+�:_��E�Yʰ[n�p��t�	���-�����:���(��)��`����xc��W�&@��'�C��c�6i�	$-��E�}g˃7�o�Y��ؐ4�C�=a�	N`t��8C0�,"��p���a�t�Wf��>��7��>�Ƞ��BHИ���!�T�E��X�B�	�\�r�[�`�\�Q�{�$�)�fI0�!�>>�ߊJ��d!��Ig��M܅ݙ�,�G�v%��8C��;v�����cO�~~8��/��!b����(��"1��I�ʵ-޳��Kim-����Y?t��jUD!]B�0�2AIeDc�5��D*�	j�%�����v�����~f����u��esv�>6�k�`���eq㧛�[�L7z'i���c�i�8X�fV[�!4�l�(�	R^>��|���f�k��D�q�J!�8r{{�Sr[�I��a���m��ܪ�=��G�-B�����Ԟ%@	�2�g=*˲&i�ٴ�� ɨtC��s�{LU%עH�K�:��� �\S:�$L�e��Z}e$�`ѣ�)���8~8��xt�^8=U��+>#х��QQQ^��	I�M�~	w.��ٔк!ac)�fOL�)�h�@�|!�\�����:��a;Su��Q��m�RʳM�Mvb88M�-4a(�Y������<ұ:�9RpC04��&��P���2Hm8�O:8�`�ؚI�&��RD�N�t����ɳ�!�OŞ;�W��!��/dL11���h����e���NI��*��%M�HC:�Jp0�MRq��J�h��ۧO��[~x����㎜q�Qb':�>���E33c�C�Q_=	��#�i:Å�\�+�%']x6	c��j��r���9�+pu:ƈ8�19KJ�mu��筗F`��ҍ5�4]�>�.O������̓}!�\�����4&��Ct*���.6���|#���=���P���C�,d>�$2��N�w{�*�*�^�'C�MO��0e��P�������<�،�����jx��u���6^��S�M<p��J�}��Ct��8��N��Mh���N��ɢ�1��;|B��h!��]��.�d=�o���)�._�d��V���)&uWS1�&���(q�)e��=_��o:�s�SF��5���߰O�84�O�L4`�e�2h�G�!���:tN�0�����<;�_XV�i���ɌȱF`ʍ��b*�J�p���[Kim��K;hf�(���TU�2h�a���m5�������D��o�h2R|�Y�څY�`���9��$<�i鲒�%&���Mjs!C|�������f���DK�zt� ��g$���(#�RҒ��ϐ��z��!sD������,�Zr�tD��P`���jFl4�<=R��j��F�������{��hC�0�22��%����*����|�NbI��Fh��/�\b�~p�㎜t�÷J�Q?"D��8���	�������jT�F̦R)3�YUˢA��o���ƒғ'��	N�6C討����Ғ!����f'���3�i23�֡�<
	�m���mƪҲ��Z~[e�b���ZBg6�ar�tX4�0,�	��72N��	��3B�O�7;>���yin~G�>����Ch ���fL�? �4d�L}�oj������e="ʃڤ�Kr��������;����s�/�1U�N͈$OvIm��4�������2|Y����+���q�q�N8���w�M�H÷�y#9��٣6d�;ϩm-���V%01>Y$�a�J_��%�C�K�&KZ4R{������J�A�D�Z�;:)0K��.Hc)�䁮?&^!��
&�	8̇��&C�*�v��2�}-ɔ��`Ӑ�@i�<��|�`�l��k����Nt���[Op���4�,��<w7��sx���]�7foD��!ӥ+����4�K4�����k�H��ONՓ�/��nIߓ�4�]��ژ�.,�,��]���qq\���:p�GgK�kн�:Sӧq��<��Kӵ��68=�j�N�W��:&Η��z3���ҝ���W����G�K�(�N��N[X���z���⸸�.+j��|Ƨˋ��N/kś^.׋����[Y��q�OZk�:���\^+��5Ǎqqx�\^8ۧ�ҸN�tJt���,���N�D��^��li�z�W-��N+���q�����ix^+��pvl��N3��ӦlO��~/��ax��?��&��z|^�ӥ�8S��c�m\w�r�4��v�V�G��f�x"}_*Ή�Å�g����_���8��N��=�������3������M*=��=/O�����/G�Jt�S��辭������xY¸W%�ū8W�	|O�B������_��4�^���M�R�!�F�>�>��ջ��v�O_x���/.��?c�}��w�F�_�]��v��fW����~��d�Z�}�Wͨ��v��=�>Z�d�Jriw~��Y��;�}��[w�t�:�a&��MeCu��n�ߪ�o~l�r�3�1-M�W"rǄ���*��"����z7A���fd��r�A��|�y��f{���k���,(��n�����b�n��!�(Ne��<
J&�u��!3�ؽ�1�c�m)3*�$�6�����;u���-B��!�f�O^Jk��u��J���<�˻�g��X���LW��h\�V\���<�A{���>So~�65�s����/웫-�/\7�:u5��m�I�rFv�(tj��Ƶ�R^�S�)�n�{�A\�|%�q���j��g�������"qA;�7S��ݰ�}ۣ��Uj�+���,�v�e^�\�ݕ�O�f��kp��I��g�F��}����b޼�Յ
�vOk;�2g8�K"_�^�D�����31x�̟_^M�L�.6ِ���6F�̽����q�� u�"j'�{3C�{+����'�o�i�ud�}�9i{�W~�/�~�ܴlG{W����Le!Z��wN�]']��*$�1WM�
a4��hII���%]a�/h�Q�9U���9]Q9~�24�"��T\&Q�Jƈ��� N>ə	�0#�L�KF�S��1ah��T���9vei�**ݒ�q�X�ٺ�tÇva�-�Q` 䊢����Q�4��uҨ���"cN��@�E�=�	�I]hAd��{��Lb�%S)d�[�Nj��勹uV�j4z�x�P�r�"�����䶪���/�g�������� P`@W������}��  X��www_w�@ W��=��ݝ�H@�IU�Oܹr���.��j�ÇWt��+���V�ϋZ�rEv�KGQ��Nl�۳L�B�8��E&�e���t�mX��L�YKY.Wu���dɦ6˫U��a��mGN���lؐ��Y�ˤ3��Ϻ�����=���h�H]m"�����BQ�q���8p���D<�sD�01$2���������z|W���98�>�	�O���6�k����y=?|6ֵ��&Cu���Ggr�t���>�!�n��a���CaA�t����)�6^�L(��<���!���D��E^�����n�f�c-m����FQ%�j-���a����ȧ���!�ߣ���Q>$��h��w�18ij��i��l��t���Jp�h�t��:tçO��}�;�]/�ც��.��Ya4�7ώ��h���!�Nͽ���{!�|d;����F���b�<�P��p�ae4vd#��L�31?+���f�O���l�|h�o����d�sG.ʒ��Y�d~�za_X-�Zԅ�u���}�(@�߿�z|��)�u�Um�#�F�y�{Ǹ�>��#ǌ��0���w�~-�����$*0��|�����͟V-��GJ��s�Lr�Ѵ\nz}=9�p�7:�m�j�t�۷�mҸ��x�q�:tæ<'�����d~�7�g��z&����**+��ǽ$獣p����͈'K�pٹ�4,~����x��ª�曎�q�d���q��̧�=�C:�J"/Z���������,�n1ɍe�bR�UR9BDrI#^]��Y=����ӧj��JY~Z�jԒx���&͛o�d���:�6S�$�`�M���ZQIL�q�~�DN'��ñ��-L���R|��Ra��I��Ꮯ8���O�cJ�x�q�q�N8�)�>b���#��;Y�슊���'��,ôE��
'=4�w�f�<W�z��c����]w.~J6�FbкY4�ʑ���9,�����G��x�^]Z��`�<�C��͸6��rʪ8t�O���<��:6"��(���ߣj�����]�!f���6�Co�a {&C�II����Zh4C���S����5��J[rܶ��N�!����CnҶs$	� �m㷮�=t�m_�8��bQb&�|'Z��RZ�������
Ǣ�F��ڬw��uT�87��38�	�6�rZ��G%�U����^ب�ad��kr�vVfcX��R�D	�`�lH��niJ��4imav�e�$��f٪[���XQd.&�FB5���1L�co������Bo��#�Z�
����+&S1̠�Z���Xy�S�`�G���N�
rUl�Ϗ����xo㓷Wu�2C�M�2�!a���}�c��Sg��[�CpCAD;I���dی&r���Y'���FJa��>x�0�G�{%ܶΧ�28�L-��e��賈a�o�O�h֗��D��;�2�\���1ڱ�0�N΁*E�������S�rM	�!Ϭ����TRb��]�2U��8l>(��2l�ei\x���8�ç��umU��&�&�J&������QQ^-x���G�'�8!�>�3*�7�>#�Ӓ%������>�I�9)�3j�>2�ϡ��[�g�����Q7:vzC��*ێ�ҹ��6u�Qe�GL�1�����&���!v�2B
,��d2�d�dY��K4�ۖ5F�C������t��;KO�<Iׅ4h!�Ƶz�tC���x��sI㉨L�z�ܗO\x���릟1X����0��h�<4}�AE�E�N{�[Kim�f|hݏ�fp�[��׏.*��S	���4h��a��m׏���9ܽyi�d!�~2z��k�R�V�!D��^�q�SKy�l�����SjCLR�a.γ&n7X]������������/�>��]Y�)�T��\K3�Ѹ~a��~W���f���W
jHUUUG2' Ç����},�>�]�(в���!"�0� j2+�p�m����1���N:cJ�x�+�t��a��Q�-�­���q�2>ܥ����Q07�"k�$�`m2&�,�!�2Re?�>�o�|5����:�;(�q�dd�Z�{�n��qS���|�BW�0j�1r���![��a|a<�M!��Fq=��6l��{r�>���q��!}�Qx��;�����^0a������>L�p� B
����|�~�Ǉ�ߐ�L�!�u��:�6q�o�i�O�Wߎ8�8��O��!b��>�(�d^�nj�Օ��8�"o,��n]��>���}���b��)믽<6ik���P��9�������DT�51�2�b��-��oX�ĕ,���᝺푟��**+�A��eY�5���4�Bۮ�����%�3��$cD�SJ�1uސ��S�Λ�Xd<NH������4��Jkc�ٲ���#��#�mŶ��C��}��V�b5ɣ/А�g�S�^����6jy�~Ҽ�)U\G�B$J9�ހe(�L���Q�[�M\�����!�Ε6��JqO�q<@�?l�?�^��c�i�CYv�95EZ�R��S��jzh:n�2B�J3�bJ�d+~�O��f�qƞ��j���Wt�+Ə��4���}����L�w�7�N�L�~EEExHC���x�m�O���ha�Ȟ�ֻ�s��\0�D�f͒Pd�jEe�5��wa�/������mr� �I����Hy6p�I�ϒ��I��� ��F^��֥̑Է�ӌ�iѐ�_,^�\�/��RH�p�rA�W����Xf%�h�i���{��I�4��J�`�EFV{?�<4z��_==S�����;�)ڿN;��J/�4|�Ē0�y�4`ٓ�2���1�a�cLc0�6�=c�a�V1�1�������ͱ��|��l|����_1�_=|�������|����1�1��<v�J��1�1���c�a�1X�+�1�1�=z�1�>m��:c�1�c���c�;x�cx�x�o��c�͟6��1�>c�6�����8�ۧ�8��n4|㍶���|�m��n�8����z�6�1��z���0�0�%��T��x�{2Tc������b*Ǚ�6d�L1.�n5��\Qv�{�������ߵ�L��W�e^_�j/�m�/��������z�Ö����nn��>E��3�V�߾�J�F}�n�>6�뫔�ⱎ������ܕ�f��]r�қK���7�Yj�/*!E��� sUӷ�OD�,v������"��T�>����VWY�=�  �	*�u������z@�(J��z;���;ސ �
 ���^������� ,�$��W�J�˕.T�B��W(MyyZgN�Ӧ0��0���{9�)m-��(�HQ�,����@�6�����Xd��tGw!):i2!�h��4�z��i�q��x�M���Q=׃���a�g"NI����y�r��2�	�2��"�]l��)m̕�Ja��i>)=�F	����2y:��&�=O�S^M6!�ɰ�����OD�tB��.��&�p�Qݦ2���L�)�ɟk���UWm�0!�٧�2�H��]�B�����;q��?1X~x�㎜q�x��풉*q-�����9Kim-�D8�Y��&�$��6Y��%�;ا������{�̷��֝:~��Yl��X^��Q�Ǹ�o6hJ��4��Υ=m����$6��N	g>)���?W�%2��O����ǆ4Xd���ē)[�~��Wԅ#�Ad5���6e��tD�6�!>���������Q�є8d<%�����O�vƛ|�J���ât�L:xhL)��:>��ښt��A\o"y�4�Ӛ�ߣn���,�A8��w,�+���"X25������S:�պ�>�.1��&Ȳ���U@��D�01��aa�Mz�(�%��,RdwQ��@d/2Z�X.����M��M�&��e�/���n����e������0ETe�*-�m��X�� ���s���2&��sguQ����HMQO�,�̐�t|��&������&_��h�6�@�f%&a�ݪ�9���ZR����p��6i2d0_a!�n$��D��n5�Ǵ�J�wV|�O^���~�6I�n^�fG���m~��y�4W�R����Te��2�|��ߛ�=�?���`�6z�U=[N�:�z��O�W�ϛV�+�/�:h�<)���؁�q9����Ҫ�4��uޒ� �I�tI��n�SG�mV&��?
���f�Yi��`}�up���K/f�3�h�h��P�ݔs�f����n�#�����p��a��L����2����m��SÇK6�9��������\;:Hl�Ζk�r9�s
88�NC�l��/���nh�ߌ��^a;�h���a���(e4��Y��6lΗ��䬈�۷��v�M�t�J���:S�4t�ИS����gɊ��i5�iXc%��R��HQ�Z�����>�EEExO��2�%ͻ���4����6�z�6���ÎK1��*Q�K6�N4e0i Y�gr�쫺�����A���墦�--$��-���[V��i<C��ᠼNe�Ce&�n��D}@ɣ0�1,�u��~��r54x0��r�~s��f����/����;�Y��N��	��I��ӎ޼t����ϝ?:Wx�8�N::tтxSç�-j�K=��<Ӡ̿��**+����a$$���u�֮����a��`h�`�I�Y��I�<NF�T�.T/7uR�-�ˆj��,�VP���l����J�
0��V>��ǽ�B|�t����d��%�eJ!a�g��L�όM�ɻ4&��ΛL�8!�	���d��F�!O�y2r�>c��=��<z�����������/�,B��+�")μ���̕�4q����#ǉ�2�w@.m�Ln4� M��G ���� ���F��G2X����b�#�nC+!�����%��i���Mַ.'B�q���Q�+4���)��!q6Rb���^��X�wJ�%��2+B�c�!V5>�|EEExO��>m�ݴ�ͶȎi�ڛW+J���V���e���Ub�y:x#93������{�2�PD�ܝ ��i�<�X��Iֈiчͅ�}�I6�{m:J!E;[6�J0h�,��0h�]���~���� Y��&���zC�䤳���6�A;���,�ab~�W�̴���(氹i��MÁ�|��&�Fl����S;-ɳ&������OD���fv�^������qƜt��+ƞ=�u�D$i�0E����[KkG7 A4�0e��"�0QF�f}x����=;�ay̅(���y�̘KL"|�E/���h�]�=�ѧ�$|<b�k�=�zBt
&]��t`�AF����ɒ_=!UA['{dS1&Mc�7@�Y�Y7kE�z8��I�VA'~���ӎ�o�6|��Ǆ(�[��UQE�h=����)�$!��}~����ms���|ssf͞pѣf�����\8v�4�:x�x�ŲYel����TTW�������\y6���p�.�d��>:�6�L�B><}��ID������&�$��M)�Nܑ8+ć<�#:B0-z�EY |>�'q_��Sy=2nw�ы�|}0�`0Rh2��I�����g'�ܒ͗�2�OW	Af)�UD�Ǔ�>*UQ4i�u1�SUO'��i���X�z���n8�N:q�n��L__|���o���#p�j
!e	>ה����
�;TF�vxn&�,�C��#�R�9���fk3V�ec=c��B�է���]�U<�G	}L�>k�����ٔ��`��ҟ'�Hd$^sg�'���M�g�*V�Ȕ�<6:�$+�B��� �f�ݘ�Z���dN�p��yɾ�%U�%����{���O��o�r��q���<vp��e��':p��1�;x�;V�4�1���Ǭv�1�Ƙ�Lt�<cx�>m�lm��6�X��[m�o[c��=x�oX��a�����c�>z�lc�a�|�>x�X񍱷����c�;c��z�1�1�cg�6ͮ�=z�v�1�i�c�1��c1���i�1���1��6���6ǭ�m��1����Um�������cv|��t��cl|�b��<q���n1�|�Vxǎ�a�a�a�<��;�e�uC�e�E�d6����󼹺��.����b�y��ٺ���N�1�?�;ט���b�ϱ��*�o��w0G����m�	��unG6��Z׍Y�=a[M�:�Ut�L��Î�*���f�Q��y`{^��d�!�n�������ط��wV^<P[N�5�r����J90)+���a7�!e��Y�*�ԩ�ġ|[H�2@hz(bnͬ�0���x�}@��@Tu��>ɋQ |)ɾI�%v���p��˵q
��0�&+T,��Û�	�c���>k%F�D+��V^���սv��'�[��J�oӅ��dWl5Mp���Rw K���ړV5� ����g1^XM��4,0������v��(��W׶��߬����>�uٍ�,w�l��&����ݞV	u��ٶ'װm`I��m�jd�ɾ��u
�[����.7꯰d�iV����#.H�[�%�Y��XӪ����嵣����W�Ę�7�o{��i{r�FY��㺪���*���Y[��Q&�Z�Y�PB9\h���ELXiI1&�%�K�dfSM*�B] X�u�IV��y�M�i�f���m�>�ǥ��MZᵤb0���z[I61TER�[vě5��+cWk#	3�m�5�⑭���!2ͧJ �EJ���%q[�3{MK�Z�	�J�.}�{�V+��\����� �(F��4��c�R�t��jb�*���s;<z@�(J��z;����ހ 0	 *��~������� @
����wwwv��  UU{ءb�ʗ*Mko�t�;q�q�<W�<k�����a����ؑ��FJ���l�Q���0�-��K�Պ]j��5H�P���م�m��\�\�b��U����v�2Y%wF�c^��B-�tcfl��k�b�f��`C:5�۰�[�˵��s���{����Sږ۫c���F�a-���FIvt�I�RI
�FL���8l6q�
��zBW��+�����^��}����ݼM�=��0��� �d� s������Vx��.����ӆ2W��		�ɰL:�Sߌ�<7>4�Y�K�M�Ʒ�L�yƝ�2OXQ��BQ���'j�r���'CAf�`���m~���F�tJ\�h]r�,��o(5Yd��*~>,���80-4gN9�Q'�칧	��??<|�_���q�8�q���}���Ő��-�����4�{����bq��Cn\�q%Qnt>l�`4�^:�lK~}g�J�l�{]n٦��!t�d���*˫.���WE�:�2���f�:}L��t�e�B�g�>OM�)Z;P���[k���C-��4�i�'�F�ǳ�0ټ�x��UeK,Xh��Ia��D�Y	��7���7�L�3�ⓡ�	rA�͚t�s�U���f��0p�m��M0�qӎ�qۥx��s��]�tFʂJ<�)m-�������m*IeTx:�Ll��Nr�KY�ٝ(����ψ8�%��>��$ќ]�mv�Z�q[]#cn`�p�ij�Z�[=�v�8�tz�^2z�b�W.:�����F���>L9����v#�ٗF�B%9yp�ٴ���ic�Y�y�tk��e7pSsG��<V1�m0�q�:qӎ;t�x/�I�$�����I��TTW�8ގ$��D��D6��`�ѦOt�/D�bbj��3R]�;�7v�e`P��0�^ϛ�Ehc��u�Ӷ�rz������6��U^!w�$�g��ag���>2�!�����SծkVcT�gM�l!��KCgS��D6~N�m���T���Գ�wc|�x�E�����n�9��dd�=x���n�;W�?4�L?v㎜t~��)	��}��^�ط��E�����I��֪�"��׬z��4T�E$r)y�)�g0ʬT���u���W�I}�-z�zݭ���j?5��X�[r��t��x�K}m�]l���f1�Y"h��Ș����nH�fW��QQ^��~2B_��30ڮ]d�N`���������g�2d,��L��k�Q���A�/�2��aꪪ����2,�2k����:��ΚKAfM�oȼI��U��m�u��G���n�m�,���ß�� �����5��������y-��Lm2o�SEE&?��zҔ��vd'$qF}<<��M�CGY���?x�����O_:t��q�6ӎ8��8��n�
xy�Tb�V.�$���Ҫ��J)�ioƽ��Y�'>�'F̅�;iZ>�Nh���v4N�Kp��$��@:Tjz��yᾘtVz��'j�j'���Ϗ'u_a'�m~:px��`��S�w}�F*i���5�4��֌Y�0�m�%�hMJMm�$�������|�]6Þ�a��aiĿBQfǤx��L~{>6��������[W�Z�'ƍ�q7��4|l���q�6��x���ǎ��Oi�{�s2Wɬ�e-����|v��''#���m�+r�~&��uv�,�O��y.2��U�{�浣vM�O=,�>�`)����4{���&11ncn�$����\�%V隹��|�����ϩ��lO��=�؞٢j��J-ɰ�N�n�$=ʪ��i�Tl�z��BBM��HII��3�J�ayİ0<#e��4p��L�ɇ.lɒ6x�GO�N�:aӦ��3����$��>|EEExO�qN�EAI�.�F{>�Z�'Xp�Ó�aO'����<�Z.�n��Hj٫]n5-ηU�N���c5�L0�fj"��|y�)�rnwKg�_D�$%�>8��#�Q)�<��6&fKO2V�Q�H�Z!n��aA0;���h�5�E���4��.[4y2�C��r����ْ��S�>c�����:W�i[~?�4t�L:lИSø��gr��j�B�ڝ#Fꛟ��N�"�bd�ʮ<!!�Gj�'T���Ɗ�̓�9��{^�3$ڢ��j��5���fVZ�����j6��%[L�
�ۨj�����#sI�z;X:�n��add���;�x#����!��K�ig����m������GR6���D�v�Y�����n*h���	�oǧ�:��=��<��WZ�Ñ�=Y��T��52vl=?{�a��Ҷ�i�^̄��C�gN��$8���"e��ӡ�xy�d>÷�i��M�>KM�J�l�\�]7�᷀d�06�����'��>?~����f.f��mu��ckVRI���8�N��?�ަ�{�����o�6���8�<0飧M&�y4�=H���QI�۟K7��EEExD�q�����<�p�y�PUP�jy~~M��oĚ*J1�9�e�y)΍��	�M���!��^�4_�	O�9z�8�Q�m�Q�&����;[���%5�Ė��ic5����w)��$3Ys���������|��6���*[�79��p��h��3�4��|�����:i��c׌~m�m��1�1�c����Ն1�cLv�z�1��>v�����o�|Ǯ�=i�1��m�o���׏X�X���6��|��Ұ�1�1�lV1�=i�0�1���lc��^1�Ǐ6��1���1�v�1����i�Lc�N��z��m�cli�6��m�[z񷍼m��n��x�q��n�|��c�c�c�1�X��q�m�i���0�#�Wn�yء��J7�jݪ���=R������*��q��;��[��5���Y��;�o��{{�o���)V8T��ɫCY[;iBܭ��#��f�����m���*�]gM����ת��R�3���f<�">̹3�����:r��傝Q:�oJ���狩Aث]���U�#{.q�֜��N�@��B�����FM�yVfg��!5ڦ�"�e��C����������T���yS}�Ӝ�����  UU{�wwww{�� �$ ���y�www{�� 4  ���y�www{�� 4  ���ؚ嫕(Z�r��\����:xa�GO���₊��-����^�m�a��a��ԟ{ͪ�WYtXp=���3[<(��͏�V�a4x��l�6Q��\}�/�j�a�ٺ*�6���ʺ���.�/KN�8B>�o�n���m�n���=�E�n?M4l�I���A�@z��IA��\�!�!�G�{;��q[��-��Ϡ��[���r=i맏��q[~8�<qӎ=`�/��ǩ��-��R�@��糒�F)o2���������F��wBm+�0�Q=A°��J����}������qb.��s7nk�c��Z��T�1�0o9�*�]�S�<{QO���&�nv�p;�#!��i�L;���)��i���%FC.�%�v�s�S�7o�·�b�jd�C&�O!����a��vNϾ��h�vn{�IN��F�ΰiþH�)�I=v����1�m�qƞ8�ǎ=T(�:�Im����r��q��%��G2�/J�&Ʒ�&$�뭹�͉R�J�Ʒ%��0��%V�)Y2I�cY�E��+KL��DX��3��ԺB����m^�����N���QQQ^2h����$!��d��IfIn�s*35Ė+��&O��m��dN�,3���l�Gs��]�]�ʇa�����0��y�sR2�?q,��.��g=!��Ԑ�xٗ���K&C�!����+pܿ,r&��I�:f;<7!��A����pW9�Uq5��g2���]eK�n��wK߽��Iߓi�fJu�B&0ģ�Y��ߟ���q��;qǎ��^[�zJ��B�ք`G�7�Ҋ��Ra�	g!��̩Q<�bHir��O<vv�!��M��GS�v��m��Ca���W-r���~*ϘP
���|��䇌�"a�Fy5|�c`�mvŹ$�%x�&d1]��\mօ�k���z}
q����#�,^����>N+a�S�zn�ro�V���y�p�_8�|Jw���=æ�0Q�Ǌ<Q��O�t��f�����j��˅M�|Ȩ��<a?����G�����&�.�Mx!p�C^#�ɲ�)>M� J����k�.�M�<9������V��~9}���o�8�+vu��_�Z�����Ŷ��q4����2e���*�	e�I�����-�q�)	$&�-��&�#!��:G���XJ2�Q�y�:4�M��S>L8t�G���#�~8�;qێ<t�Z���n�e��e�{Kim-�w_���{(@��ݝ4�l������̮~��'��l��9ș�GIm�Shb�V���n�����ߺ{�{�fߟ�N%�:��aڪ�>2a<���l06������p�TD�Y�����ܱ[��m�ś���3�9�S@=<� S���She�~7�m�����Y�G4�t��N8�N4��W�q㎜v��j�-�F�L���=m��]吝b��+���}���B��]X���CB��$�g�Zf�����rGfף�k��`E30�M���r��0"��;&���V�`�kMH�����[#��t��,�Y��KӚ�u�K�E�~�EEEx�<�Կ3V$!�-�.��!z�P^*�\�$f�&�>�]�����>j�E�d��?lD"j֎�na����=6Iv�]�bi�xD��J�z�P�zw���'Ɠ�O=0�VßI�֧�"Ȑ�������Ҍ��C��{�N���b�Y�˃�c�ƙb��M���,o����v�l�V.H�Kt@#E�������|k�
�,�Zp���:|h�G�8'��N�:aӦ�e�s�
%)}�Ȓwܨ�����D�L�"��˩UP>#��Ua}�gi���PCG��x&+�ږ���=K�2k�ɀ�H��p����z�q�)
�4��%�0�$����gK�;�8�dm�~��R��f�����.�.�4��5ށ���W�OT!
���C	��i!��Q����y�>z���~c��J��q�gM:x`�/�yŔJʕ�{�
˚���	�}Kim-���Hd��)����.�����2|��[��ę7��<P}��5��m2_�1g��UֹF,�V�H�֗�3"y;/L]ˍ2͆��>�yV��mKn����M�
d!�0e�H� 5m8aܦ��p������9�v�����k���nծ8�����+�q�v�N�&����6,R���Z����T��z_�tU;r�M�{��5VH8>����ğM�Җ-�u���H��ٺ0Vi�(���������G�Ι���3�������ǟ�8>Ϫ�F��p�|u�zg��mK�]�pÄ��c����%F��k�[�A�}RD�c��z��t���Zd�:nI©��Ҋbm,ǒ~�Hx���oϝ�~i��m��m���ϛc�Yl�+���<c�z�j��c�:c1���>c��|��4�co��z��1�lcm�m����lcl|�O���6��|����b��c����lz�=c�1���oj��1��6�1�1�m��1�o�N�;i�L\c�\c�\cx�xΖm��1�t�lx�=|��1�lx��1��޶����X��om�������o���8�1�m��n=i�1X�;c��m�c��Ǯ=tҸp�Æa��g��W�[��;M̋�YV�v�6�m��oY����^}Ź>=3��k�Y�ݭ�3J����b�ؤ���dμ�����,���VX?sﾷ����s {�آ����F�Ͼ���N�u�j;�z�tDD��nN暌f�Vw�X��+�[��[-ت��w��t���4�n/��I���L��.��'��W.W"	rYZ2��Ne��Y'�w�7?M�OFb����ɃOJ�K�c��I�r5E���Ѭ^}f>�J�e�\���ٳ3v���ty����$�N�Kj�n��g�غ��Ϊ��k��г���-�ّٓ��w�����5y�X{ə��"�b�?H�~������y˹�U�K�/���0�9H��o$�=���X��Z/�m���ZkӮK4����]K�6�\�����pgW����z�1�c����|v�1�X����s�I>��E6qU*�&��*e�'�je��)�mL����jA��ti䤦X���b
�%vh�ւrV�5d]�m�E�jr:��
s�ު�*w�1YI�#��)�.�CE�f�l�.�X�]�2�RiX��ZUe�����*e�3��;i[Y�,v A|���u?5���il^�u2��ǖ��P��E>�� ,�a#�ޝW|����#4Yt$���Yh������/zT�Fh"4X&5k���>�+�!4�֭tyٓ��%Ii�v��ͶMKv����$�,�*4w߼���{N�4c�i�0��o��g��
Z�V�ˋm�����^�7���q)׮]�Ժ������G���   *���������� 4  ���˻���� � UT{�����x@  ����\�r���\Ҹc�8�t�ת����<��3�6��CcKd��n�״��5��� �gq��}���+n8IHV�q�Y�&!�*e�p��o\I%&�T��Ů��H2�nt��%�Q%֎�R�B2͉Zb�CY(փkK,���c�0���**+��I��-�l�K]l��kDn������J�N`���\r��#�pŘ6�h���lm1�L�:��8ka͚<p<�a��k�Ojܴ�֒fFOuᯣС���2�t��Zo�����Nl8��!��Qd����S�RV�bL�0�7��=(��/�����K�{^ب����p���Β���'��������j�Rm�lvӏϚcJ���qۊ~��>�<S�a�U=$�W��6�i�0ҿ&�$$�}���`�G�=�Q�UW.�G:�#�GCz��'�RԐ����񽾒�I��&��'�O�RP�oC	��D�|�?9�����sg)�^��x� 5�,+���䐵c�%"�l�$������&�~�{�;6Y��}� m�QXM<xxN�w����P��'���"����j����ݻq��O�+l1Î8�GM<:lИxa��'%�D���QE�>2Ǻ�̩m�1j���,>	���:������2�9\�*����zT��~�C���P����'���^�5�7��t�S�C+�f�U���ZԳ�w���>w���Mɴ�'������m5YC>*��ģq�Fæ	�Fdd�7���O�˪n]���w����i�`
Zm�n�:cO�~i_�q�iӎ���b�Z�D<�Bc@�1�7D�C�a�U<��}���[���JSD!�?-�o^����(a��c����ϫ�����>|(z���'�����,��e���'Y�i�L/P� |��]�A���潆���çQ��M���=}�������w���S��f7$����-��hEW�9�1���ޑ8{���I���ɂ�4p�Ƀe�(�J�~q�q��q�]�������W鄖,9,2:��I��<���$������|]D�d��Ĳf�Zq�Sb���f�\ŷr�b��2ň,�yi��1�S���+.%�� ��e%�%�ϛY�-�D�1��u�cթ�	���-��� @���s�ݬ��%Z���!x�߇�?)�p=���T�J8h�����?D�������j�=�7�iS�ө���e�j�����df�jށ��<�Ca�9LM1�f[��i��w2��}�g�U��L`�0��ʣ4�:t�۪m+��`�e]T�a��Rx�}�O�Cn��)���kJ�m�����4~>4|a��i[??8�4�n8�ҽz�z��D5��Dq^uc�&�nx��ʩ��|L�H~M3.���Q�06ny�6u�Q�r���Y$z?4�O��7�'�a7x��.�	�0���	
�_w�ٟ�z@�ƅ��u%���FBvCWcIPXI$����8�$�sTM��
UW����a�U�a��&��B!>���d��9M�Oi���ś���ꤞ�8��I�5����i�%Y��>(�D>����ӥ:xh���f��f��+?R�d�Ct�1Qa�{D_(���l��I�|I�o�x�î�А���N�p�u=s���G�<���vf@2V�+��HQ�r������IFu<g���S�g���e5�zT-�.��H�z+��ɲ���ވ�a�lF�6[narS6z'f}��8�
N���?��mK^)�i�����?������?=i�Jُ�8�8�ێ�&͘wǶ�"�#�c�i_�EXvo{�¸������(�と}�K�"����U���Y�u� ozՁPӶDȨA�RE����k�r�Զ�����p-4gE6�	�}>$3ʕE�/^�����`|�M_ڗWc��o�ܧD�{�"u*�i��E�L��a�Ȓ�$�OO��p�q�~|x�m�˹6x�Qҍ2`�g�:Q?8�8�N<v���WO]1��>��k/Yz��X�<�\D��̈��
l�0yQ3Yfpj��#�,S�
�ډ� �(�0�}늧�n4ᶎXX��T�X�s�(�+6��n��!�%Ȝ�hQ	�I)���[
}�=��_K�֡J��r9�� A�sXc�ˮ5��Kvv3i�vq)���v��ۉ���kq�W�l]h�?G5Ϟ���a�ύ�Xh:�ϋ^*:1�m����Fxx&K3r֍E�M�@��$6�8�3�$f���'���?qg�Q-���b��_��HK8�k-�a&���1I��E?ŝ/�����?'��<䵣�i�v���OZcJ�q�i�n�q�6lÁ�j��s9�(�̛�r�7�,4���A�Ԫ���t��m˟IJ�G�&ݤ,2�vgR4�_�Ç�OUQ(�h��	��͆Mq������~�j����	*Lf
������ʃiɐ�?I��ύ������
&��\}�r�McUCć�H3S'���>l�=�
&��o��u6u�ҽq_=z���m��lc�1�c�1��Ǭv�1��1�1����޾|���lm��z��Ǭc�z��c��_>clc�<m�co_<c�m0�1�c�V=c�1ٌm�c�x����������c�c�1�m�L1��cLc�<c�1�xƟ6ߖ�۶1�c��X��ox�v���c�+i�m����q�L1�i�c�1���<c�<qۧ8p�Ç>U�����yמi���_}'5
��=�j����Y��Ҧ��fJ̮�]M��]ݬyһU2�7WM2|6>6gk=&j�?�)���bӫ�]s�k~�J�2Ґ����~�_�\�^*���.��z.� �Z�K��4k���;ד���Q��]�^�{��>���O)�t��˥x�-����:��w9ޒ�o}�Ŋ0�'37��q�C�^��h�N�nD���"��jZ��-&�=��  8`UUK����� � *���������  p�
��=ϻ����   UUG���-\�r��(M��:q۷8�ںz��uiE�5��F��j�B�f����q��T��|
��8u1Oi�Bꛡi��y�ུ���@�i��Ӄ�^�#^A9aY��A��Ϋg�4'C�qPy]�|�t�܄��r5�##߉6��N']�-u�I��H��ƠM%h)�u��J,�G�>,�F�!���:q۷x�^�t���t�V��aϕUMtu1b���ӝ-:~p�Hm�kM&�İ��J%n[$�����j��Y?uf�֒'	�<�0p0��I�����V��t4����ͧCǋHm�qӶ���r+}^N2P�=��a���4�EeV!��SI�Cqc���AD�f2�y�u%���>0��G:Sm+����qӎ���ǯ��O9l���O��oz�6�7�,4s"S[[V7!*�
r�sf��5U���YR��C����Z�F�13a�A[+L��ev��n��Θ�XBHi+R]5ƾ��9��h�H[�.'�΋.am�CI~� "��ȱ��5�^׆\�i�\9ed��ofy��.GS�P��9�K�,����8���6s�O��q�X{���<�m�ߎ6Xl��Z��n�J#׏��/p��ut��ᔴ����622�0S�����$I���֢���ÿDS��K{<��C���|/���g����iv>V��nZ�ZT)��++�R��yR��y�����A�=\�~_�m��V��;���v��n�i�+l~c�8��N�q�z����b����Q�N�R,���-B��Mc\�UTg��f�~<;5Au�k��a[O���=�J|h78�z�*1c/�c5a��'���[G��ɴ�#S��?\�W���r?mj�I$�����{!��y2��h7�O��g�t��km�mݸ��B(J��W�������!v��JO�(�=Ul,������6y����
ͤ�����3�����x��:m��V�8cqӎ�xxt���l�D�����m�YZ���着��&��7����s3�gsK��lÒ���]]�sG���������ߒ���}���73����㑄�(rEq�HT����{ěKiM�ӏM����1U��T�W,�-�\��Fxx����*�6���D�9f�g��d�1�*��3�/^��&͙(���=t��m+?�t�8�ڛ6a�=s
!�2>�UN�O7Ԑ�!{$4H+2p1�'�6�q٭�yz�묚٥��?q�'��BQ��f��İKF��w/��0�{Gc����kǊ-<֡!�)4N;"ypu[1�	!*��UXq�?p�Gn7�˻.Uտ`��nHd�U��g���ga�花FwP���A�h�-��L�xكE�(٥l�~1�8��n<x�ڴ�ӌt�\	��;��J�BpƠ��Vbs�1n&��f33�$�[6���I���U�"���E#C���A�df�.�S��V=�Ŵi��+M$�m
���^�7��b���+"1�I����໬����� 	l(�e���m�"�U���K9�݊�\�D��%�Ř�0k�А��
m�	�~:��ɑ��}V���s�_.I��n7��O�^�M�÷�r���ɛ>��Н#&��N�9�h�-�Ʉ�M9t[�~}UR���6��d7��ٵ�wRrnl5����2�U�*�.%զ��5��ut�FRGA���Ď��p�͞FC�NO��j��������������8��?�����ct�?JS�<x���d�Ef��O<UT�`a�Ɵ�\0�|��	��t(�4q0���C�ܨ����Щ��a��K�h��C�~t�]B�4���&��v��츉\��Ye���ȩ��5�Il7c2K���E�����gɓ�D�*h��	�����_2�!C��##&�y=VS�u���S��:aÆ��zS�J���Ɯqێ�<v�<t��NB�egSd�Zڧ�*����r�R��_g��{��Xm>�����>�Ī*5_z�EW5^#��jF>�?<ʓɗ&aK�\.h�*Y�N���r�R��kC��l6#�pj+Gp��xL7��RL��2�:||�4t��M�]Ɯ`�f���'h�t�2�O�I��=y9ƞ���1�4�a�1���Ҙ�<x����������*�1^)�0��5��SS��c��ߤ���L/�[�/�Z�ro���2�CPٖr>�pԟ�s��Wn�����>�����ߏ`��urc)i�S��{>!P�t�i��?q��t��>M��r��@�����<q��p����Oڒ$$�ʨ*��H� �?�?�?�Z�v���z-���;��KJb����]�2������-�"�*d
�"�I*n��E�T�(���Szh�)TR�),�RYIeB�R��e*�KQeBʋ(���%R�,���R�)eE�*��U��*-�YQeK)eB�,�T���*,�R�K*T���J,�RYIeD���YIeB�*RYK)QeUQeIe%�YQ(��KYJ��ER�)T��P�E)b�V*�YR�,QT��X��UB�U)e%�U,�*�R�,QiT�P�YJ��,���T����%��X��eIT�J���R����e*�)JX�R�*�T*�)JX��!eE�eR�,��*J��UX�(�DA�H�1" �,�ieU*�RR�)UJ�URʩR�IUT�UKUd���(�U�UT�R��)V*J���Y*�b�K
��e*����QUJ�*J����X�����G�����U�UY)Ud�UT�*�,R�T�R��R�d�R�R�U)b�K%UU���UU��"0B2"#""2"#""1T��UVJ�X���%U!`�����Ȋ��R�UUU����UDdDDFDDdDF�0B �`�����Ȉ��""2""A�"�"1��DF	"#*��UX��*��*�b��F�#��� �D����A" �D#B�V*��R�J�*�eUYUVT�VURʪX�RT�U��*�b����F�X���J�J���V*�YT������b�VUR��K)ib���YDA�(�#��1�V)*�U��X�R�R��T����R�*K��X�i)VRʪ��*j�H�H��Y�"�H�1Qd��J�$TX*t�h���EH��TT��!Qd����Qa֓��D������i
�"��TT*(A$	�OJ`Q&F"U"��#Q*,EE���*(TY
�J��E4�T:B��QP����!QH���H��Y5H�EEB��QH��Qb**B��QI*iP�*)����TT*,���TT���Tҡ�**%E�TX*,"������B�����Y!QAQaEE�$���AQd���Q,���TTJ��Q`��*)J��TY
%�*)%E"��H��J�Qa*,E�d��,�R�T�%JEJ�K"���P�H�A��b�*$@� ����b(*�H��a,B�$T�
�R�
�K �R���JB�$T��XEJ�DT�*PR*
PT��T�)R)R(�X1V $T��!P�I)PT�%,�J%*IP�E,�R�KJ��K
Y%JE,%"�K!R�)R*T*Q)P�IR�K$�X�Y*�T�K
�%,�K"�IH�RĩH�
�%,�,�K"��*Y%"�R�R�Rĩ`�b*X�,EKK$�AH1BT� �`E`Ā��!H�$̠bD���V��R�JQd�J��*�R�JR�JR�*�R,R�X�*X���K��H�R�d�U,�R�b�R�R���UJ��)Qb�H��*X���R�Y*UK�ET�R�d�J�*R��J�X�*X�T�T��R�J�R,�d�b�*X�U*�*UJ�X�JF	H�"	$D������a,A��ab�dB��"$`��"$`��,�*�b�T�X�T�X�R�)B�)KJX�*�R�*��U,��Y)b�JU,�
���K%*�JU,R�eB�e*�R�b���T,UU����[�iJ�UBʱK�(��YER�*�R���}��%)b�K)T����R�*VU��YUVUQeB�e*�R��J�ʅT�ER�R�(�P�JR�*�)J,R�U�,UR�e)V*�������V*ʪ��e�R�%�Qe*�R�E�Z,R�UR������Qe)K�,T�B�T�����,R*��UJ�K)U,�UYR�eJ�e"�eR���*R�T*��J,UT�T�YJ�*U,��eB�ʕK*�K)U"�U%�K*%�eu�ꪢYK(Z��K�*%�K�*%X��Ib�X��b��%��b�E��X�YE�K�*%�K�Qb�uZ�,QT�R,Qe,R!uIK@,��b�X����QE�,�YQe%��T,���ʪ��T��T,�,���eE���P��(���)V*�YR�*9BCHr��A��5�b��H�:
�����~�*��
!$���2B	���k�I���_���s����G�O���d����3������������d�'��#��21����N�肆?���/ڜ4~_�����3?1��c���d�K�����a��S��op���G� T �����������������0~_�b�(��
�������;�h��ІA�"P�/��?�7�����!���?����֪� s�Q?��������~�Ա�:�����W �PL$�!l_ޛC������������ݭo������Hj�?]����c ���3��o�cz)" ?������ ���H�� 
�"�P*(�?JF���`(��e�*$mi��W �t��]�
����_������U������A�FA�UP�T��DZ�AԪ�$YU��ƿ����`�M��3�؁��#���߀z� �"���P���������G���g�X T ���ʖ���b�^�����C?�����������Z`+`��?���h�?�������~o� ��ο'�����O�6�?A�t��u��,��>?��w�?�}�p>?�Ӥ ����ET �O��U �w�ց������򠫰?}��>?���p��X+�S�P��TAG.V�I!�l-�X�}U@
@������ڦQ�41��`i%%��)�zTМC�G��n�k��r'�h�Q @��?����?o迷����� ���h_��R~���� ���9��a��_��H��������~��A��C���?��?�ܐ���G�����a���.@̧���T DO���uTP@����G��_���<�0�����Q�?M���`iF�!���x� ���n���H���� �n����,?��_��s �k�~�ʪ(��
�+�C�C�&�~���Q���"��0�t?�������<�8���+z0Q�z|������_Ѐ�D��_��g��+�����?Y�1���Wp����t�J
�
O���������C�Ҩ� ~�&��g���H�
Te@