BZh91AY&SY��8�l_�@q���"� ����bI��         �ƶ��H���*��Z�I��0Ф�mQUD���L�l�E��%"��R�%CF�Ze���(dR�+U��5��Z���!JR�+VҕR��2�6�R�XcUU�&I���Vk%��S2���lj֔��,ՙM�m�d�@m�fڍjBMm����OZ�-�d� ;GI4��J�p�]���6Գl�6���Z�klք���iQ�kYmZյa�3Y5���[kj�ɳc+T-���ew�z��U�Kd     ����j�] �֫�������v�M+�4sw9��� V��n�, s`v�:�&�u��{�r��.g[,l��Z�M5��*�  ��@�PP�͸JSup  5�^�*�;� uB�V���
��  7}�<=JV�>� 7e4�.ѱR��[a[m��jI�  d=킀 -���J�pԚ S8�:@��t@�#��:�(+��Ox:�zS�z
���W� {m����u@ ��5)�2�2U��"�^  �w���ֽh����(wG�� ����K�a�B�jӞ���� ��]��q�� �G��{Ǫ ����,@X���6�ͩ�4�5��&��  	����ޗ�G@I��W@7�{��� Vz���н��7]=�� �����i{���@W.׮� �w �^PQ�&U��m��8Fl�  Ϻ

V����ҀYOn 
z���t �g��Cs��M 0�(�hl��(�M��x����j�����
z� ]��J���b���x   3�y�Jovn]�CB�miɅ ��� c Q� .�` @R�6 �nsl�kcZ[1-�5Vb�J�   �� a� [��]+ P�� 
�9s�(�;����N([ �� i�����Z��l�ֲ�!��<   q�}��T(��8 �up �� *��=�:�� YݮP(ۥƁ@�,P��ܧl #GL�[k�k5�ՖU����  �(/f�� �w  ;����}�\ ��
hg�w hwg  Ns� 1��T�      }    j`�J��  � L ���(�@�C@i��)*�� ш  4� ��R��2220�M2b)�HRQ�m�0&� ���%$'�Q(d&M)�CCjP�O_�����w_>��8���T�������7��J��c�GAjה9�A���������_�@dT?�PW�QUQ_�G�O���p����������?J��?����?몪�z<EUE�����xB�� "�����������a��̎as#�̤���as#���0��`3#���G09��ds)��f̤�f2���`s)�L�f6e&S2��̎a3�L��S0�9��e3#���̦e3fBe3)���09��e3)��0�es��0fS09��`se�L�fS2��̎ds�\�L�W09�̎`s�\��G1�I��.ds#�\��G2s����0���.as����0es+���I�3+�09�̎es��2���.as#�0����ds#���G29�̎d3$��09��`s#���S2���fa3��fS09�̦e�)�L��S09��`s)�L�fS0��̦i�̮`L��G2��̦`3$��09��`s���a̎e3)�L�fS2��̎`3	�L�f2��̎d3)�L�ff2��̦a3)�L�f09�̦l�L&a3)�L��29�̦e&�&e3)�\��3#���0Les#�\��W0���9�es#�\�� ��C2L�0���3+�\��Y�2��3�0���.d�����\�� ��d��@��\��2�+�\��0��3�f2��3�\���L�`��@�.as+���� �.as�\�L��́�2as�	���0��̮es0�W0eș�3#�f@̡�G0&a�f� ��0+2��D£�Ds �@��fDC0��T\�d@�s .eQ� aE�"��2
�D\£�A� f@� � fE£�s"�`�*9�W2��ȣ��3.e̪9�W0��@£�s
�aT�9�G2�L��@s �`̈9�2�� 0��G2(���d �s(�`3*�dE���W2��A���0��3#���09�̎dsfFes+���0���.es+�2&d��̎as+�I��� ̮es f0��3+�23fW0es�2`��@�&`���0��̎ds#��Lf29��t�&�~���c�?������=^X��3�>�;�"�Vˀ��/I{�6�֧gm[}��*In�x�c�uk��x�=݁Ĉ�v�C3�xm�,�,ה���ܻo,��U��7�48�ɚ���8���`�(��"���[������¤�-��n��pKu�1�F�2���HV7z���R&?[��`ZJ%�\��9��iK*���Ȑ��C���b���^*�4%�eD�Q��'H%�F�y�X<��t����p�������m�,m��պ�\����u�}5\��4��R�y�E�Cs;���]�E9�^i��|N�yot�Eo�$Zw�|-�2�0��K��l+S���yrdDD<P�БHyJiEV�HQۤ�ùV2^S{	���M���Lc*]��5ᣱ���&�8�7��ii{�3F6�њ�If���٫V=*#�E��EL3+jSCw[���;�.�J��b�v��i:�d{i���fl�rfޅ��Oz3tJm�ff��*M^պEEzZ,$R�R�&�UckJ��Dɲ�������(;�Y�B#CaUg 0�5��V���f)X��,�yYj��R'����A�hC�[mDj�"�A왴�7�\�~�5wm"�סrś��M��GaGu��@1X)zU�֖iu&��ڪgsJ�à�b�|0]���/���t;�>��p�M�iYYYǁT��^f��P���(,�RiJ;r�3vk�1��su�2�9��/��=��n�z.c�LM���-���s6Ý�B�**!˲�`��-L)��&�Y��Ht�����?j�*�v�0hTTj�7+�2�3^jc�V��^=����Шp��U=�K~ͳDəi�a����ɩ�b�^,LcGp���1&��5����B��F����ٕ�
�v�m�&š
F,�C��"������]��س1���P�ekѱ��l�X���S�W>��Ul�D��Pt.��+ma��Wp�O�{��@�<�GiV���U��u�^�+H/*�v��Y�1	����)�T0ڄ7"�-�o�a�F�ذ������S��k���bui�wi��]��,�k"oiI�h���I������݁X:R�W�9&�z��!עm���kBĪ�꣕���֊�F �b��]C4�7�6&�R�k1�P$�j���M(&e�(8�1h�[).��Url�{ٛR�m��hr��mS�OP�O ����k3#4`n�ѓa&�b��36���&��tS�"�"�d�%I����k�1=��k�z�᎛�3r�/�P麡�[�.�S̭#p<QlI�Ǣ���eS&XQ�ᚵ��VeZ��}x��TL(���m���w�k�L��gV	�u��)��!ڰt6N�]u��o ���Q��
G����WMxdË)!Vc�x����V��V:�f�,m5��J�[z��V�ض �-R��i�o���dh;1���3	�t��MV��z,�T���w�h@�&�4���É���8�a2�"+Y �]�s61FK���t��Dn2�9yN�8BJ7��1��jm���D�W�����df+K]�'p*"��CM�o7}ʒ��{i�Y��U	kV�{,:��ι5�- Ɓ6��a�e�ա�m;F���]�ݩZ�Z{Bnѭ$���M�ǎR*�oj;.f��+u:V�tMܙ��F�u�lх�����Լ�t�1��3]�{�ވڈ�J6هc�6�!Q�����!���b���͔ �7d��l^n������Л�rIO4�԰?s3A=C@�X��{I.��V�ٶZ�J&�N��I��+6�ضf�KBׄ�fO7���  �<�-�۬��G����\Lћ�n��0�U��M��b|��o˫_��J��9D����v�9z��V-�f*70Q���a�K7���n={A�����S��k�p٬�ӫ34X��m˚��$6Q�kS0V����eju)���.D�ꦱ&�*��5V/�1�|	����hj!�U�
ł��N�Z��ΆӸ�.�[�t��2�K���*T�V�5�˘koVc"γe��wvK�Z��B�Ҙ����;י���opD�RMK�x],��'eiz��x oq�ctŨ�kO��&h^�A�ڑ���I��Z�b���= �Y.P݃$�D�T��cko1x���ܢ30e9��7c�H��!��Zl�r�l*߱��X*lيA�C�UXux��i]�:���|�k��،{E���b��U�ţ-2(�%hR���c���hn��ѝFvU0�+3*m����ͭ���=-�Q���T&�h/�ܧ*ܽi-�ND�^I�����e�ye��ja���3"�^�I��Q��3�dä����ڪ+E���U�$����,Df��<��4qަ��Ȭ�Vp���"l�r*(�j���݋��0��9-�ԙ�5�Km��q��ǎ���:���o�.�7J���fi��,�)�m��c��u�Zs�v��c��(K��X=2�h����C�m�u��%��R`�S-�;w��`��U����Xѡ*zZ���&�C�G���͆���t�� R�.��wL#���y���ov��5@��f�M(�$6��eeCr����>����ډ�Z�6�y�6D�5h$��H`�4�v(K2�1R�L���\b�ך�ʹ༒b%=yZ�M�<܅wD-�V/EǄ�v9ι>�QYΑ-�оyI�X"��	�҄��R�&��Mj�&��s�S;�K#o,e5�{k-f`N�Ӳ��Y�B�m!;sGtGK��1ǅ�qћdm1p��;{!�	��i&f�p��Q���O�M�j�W�!)�d�[c����LXKK�;Cv��������6^+��G:ٽz�F����lN�dв���h���i��.��8m=�u{�${@���t��z־�����Tt�A�1��u��Ӗ�d�����sH�6�
��-u�L�n��\d&�j�z���w*�)�H3%�8٘��M�3t_�S�	��w��:���'XV9��rzooAET*�,���Ylj�t�z��/*��d9.���E[�Cp�Fjm�G][��H���%:5�c+D���/)���挠�L���.ؕ��A�l^L5�������"�(�����[
&w<��Y��p�������䄣*�kT���n]�O]�]��dQިl���z�x^+��4" b��˺SH�����
4�n�#V,7P���Fj��e6��\�3+Zz�A�vb��+%R5�̷��m���r���Y�Pt�C4�0C�ewu�x��uKvc�1INɬ(�	��q-�l��2��v��n�����e06l&�H%LT0�B�h�ж��iZ%a�ܨl��+IT2윌Z�$G�t2l8�⩃IǴ1���|��	P e���d�_�˼oޗZ�H�ctZ[xN
�aA��:�!Sz�e�Q�Ѥ],KPo#IGA�1��M���عU�b�$�fZ��Sz��{��T��j�ĭ驵�w���ۢ�#��1�S61nVF�N�d,��ymRG6��+�;�%�`��ݻ��f�j���`�Yz��k�Niͭ�M�լ7���B�r��鳪��HU
�Ű�/P������Q��&�������2(+L�⥒��Z��]���k�l,��f�{.��ĴX�B9��d�t<��6L��`�.��
y f��[�т-2K��
���n���ձ��nC��R�ifn���w%�gR�6��1��w�t�{Խʆܖ����)H�m���/�E�!�$iF�&�˱6Q�ڼ�wmEz"dR�lP ���	���<*�S̈K1֠q5f��Ҏ޺�)����˒K��h6^��M�2�e�J�gU]�#*�+3Ψ4GU��v,���M�H��弁��C���w5۵q=��D<�q��Rr�@nC��Tc�V���kC+\ܺڸ��X�Ӱ�!��i˕m�(�=٥����QV�B�6����d�4���;V��1m�̔J�قd��z|�Z�U�2� 3BlnVÊ�k�IhL"l]:�E�X;F����-&�ZI�t�l�LM��̔�r����z,�*;�ZD�c:�VH�b7t��ʹ��d�"��^���(mZpaũ�h4�^�+�hٰ�4�Գ�/c�wm\Y�Ci�kF��� ���b�����;B��{0k�aJ6|�y�[��뻅+w(
њXŎ�77K#�nK� f�"ynY�`I�q:��ߣ5*����6n饹�ƙ��vM��˲㠝t��W2�l��F4�̬��/$�rՁ���V���v�����9�3U�W�b���zI,��W-g��t^����B��(�ʻ���5��"п�.lY�#�R�敵#�
]���6�oJz#Ͷ���r�Ÿ�6�ۡ�&0u��J����V��#����u��+001�%�c���n�lh�r�Щ͵���.]�q�	<��������kT���N�U�Z
�]�x�I h���[��|��u���� �9���w0^&F��V�ȷ2�U�sBØ���:Gtm�aK36'R����̏k
kh!�n�9qZ���T"�9�v�K
�یV]e��u�6��7���~;���][�)M�t�����V��D�lx�:�*:�jR7A������O-d�	�&�ɥ�&�ku�F�.��n���]{T�c
rİU�6bZ��kec͊i�MiɊT������^$47�k�$
�-�ak.���e9y�ޛ%M�eL��^;���I�=�iu2R�j��2��)��{����m�f�]�@m8�6�����A��xH�[�0����M�V2#�^ef،ŻR{b�c׏$�i3��vj͜�D���wK��H��!���ں5V�%رY^ct��n[��X������ù���\�+F.�Ӯ��66��6�n�J�怣��ڦ*1�l���"p��f�f�"L�6��4kf��]^m<��Z�!�2P�2˖�Xˑ&r�e�r8Iͽ�fCy6�%ց!+��y���
Ygx�l�w�v��(�'�RB��х�(�ѩm[iS�����+
��f�M���1 �Uk�g5$�q�@��p�P��w��/9�X�,��4!�3K�Ӭ��V�4�V���U\��)$��Fd�.����*��4����&�K�"�t�U��i�)UlN��yc)��7g��Ǧ޴��0��U���/L]}��ճe�/�Wp�J�49���-� ޘFiZٻW/^kK��������c�0�ӪeC��s$Ԏ�h�ӻcAN�X���aܣWe��������
�]�Z�A0b���u��ճM�Ї��b��Q\�!d�a]bk71�b4���앃"Y�-9.�z�$�`�C6�Ԧ�3�≩p���nm��Z+`�ϫR�!�kR��cm��-b6Ի�Y�b:q\�� cv�[��=�"��( n��<�Z5�����r���;�e�AWpf-�ե����j�jmʏ-�f���Y�����M�҇w̡ŤwM�.���Y���}��� �v�x��T�f�n�6p�pWE�'�AVHq���6nEk[�f��AH����.�m�M��pV������~dm�z�{��`�������1���BXݘq�u&-b�l�OL7��J�H�L�b��6�Y��Gh�{�`��E{R�sm9�i��1LKP!2���+V�h�q�s���L�x�ߦDw���ƽ�X/Y�{z"t��2�0U�oU]O;�]���m������a��܆��.Q�JaB�+Oc.�ˠ.4�z5XVQ�Zn�T��7$��a�0�4kj-��h+)�̞x���-`��K�Yh&�z����L�����ǖS���]]�;�{��M���ʳ$�NG&�e�2ͳMA�0¯n�γ%�PXٳǻJ����}�e*)pk���D6�\��T[\70j��YAS�{����Nl8U�cѥA��CxM���D��ͻ��MXu�G%���(Hz�G���i�%壎��7�YP�)Y��Xjݝ�`��N�R:I[K87׫\�`�ܤ)=����<'frtԍ��J��P�]	�x�6!��a���>`��r�����8�My���,� �ˣ�13�+Q� �z�dz0%C��=
�HH0�"́a���=Lb�l�F`Ch�Ȱ�q��g� @�3�w�@AA2`_V4=�"�(�7Bg�w�����aPU]�+�L&�xQf�h��l��3�Vnz�/J�`Aah�2G��m]C��A��,"����fO+�R�i�#���"���GlONA\UGufI[8��0�j͢k#x��*���5�0�K�`����09��� Tt�w��ɲ��RS<� ���,[	��Ux)��*�c��2�^.ypon)�U��! `0H ��l���٫u�_A�zvNhL02A�9�U�A�A�E��,"D�`]�p�����<�\2�j�CBh L��7K�8(/�ۛ��(�"B�`�'Dϴ�q�]�X�R�d�d!FQvUfH���"�.��A��.�����c9�*γ,�H�!<(�y��¬�S�faB�1�YxD�6:�/���Hv/�������+�2�VV�k5���{�`i��X�PyP�3K%���7g8�5��$�3A���¥8�C@*E`�(�zOP3�S;�6l���E3ݙ�ψ��!Ea��L�eX�,\v��tZ�B���GX���EɰN�����e=��z}�o�ݔ?�￟�Ъ*��~��I$�I$�I$����dǗ�]��\lA��������ӹI&�n�R�4��3'd��X��*�man��ԧ\&l�i�%�g�
�c��VstP�Kx.���}���;0�I��ʉI����'q�q�0�C���mhm�RΊ����Q��&j$��*�0ّq���r�����6B��#5���x���7���N���y���mB�6�:���	�8�Z��x���C���Y�L�b�b��H��<���bg+vp2��p�ˇ���]��7t�f���SS��M�-[z�08�)�F�@�[*bz�Zt�Vx2�Q:˲���SxS�:���MvAR�+�^���k!PT�������͌�Ԣ�6�Ew�#:�u���A����2���b��jk�}؊�Cw�ɘG�{�M��JP{��ˍ�C���>.�:�+V^1o��={�d���nnZʚk�B.�q�fp9��AXJ,�#�f�JVSU(Wu��徜�	d�t�}�[�:����v��VtWٍo�z����
�ͻ�n�e��qtn�'���.ˎ�m��~��k��+/
��t���\�>��n͑�I#�G./kf��%�Gnm�t������N�`I�w]-6��&O;�K�[{��b����%rD�}�-�h�{:���-e^8^�ɬ�������K,��h-��L�hڕ�]�0P%�B�v���|�d4�E�r'�,wR�)qOe񥨰v�lH���R�}k@z�*���4<rK��b���ævL#_U�Z�ܫF�[o�fEo3��s]	�����l.�AXn��,�'���K�+���D�
�ո�,��	��t}y�ܫ�m�dr�o�وt�b��坌g�����'
�����tɺj���@a-����]�I�)�L�MvWdޚzY×J�"�8�fX��}��-Fr
r�I� ��ַse0X�����ĕ�|��p��A���Oc�9�C%E�l�{Im���-�eu�+�;��fWr� ����Uą�jvevF�E9��t���y{[�,ī�X��B�&qQ=*eK/�N��IĻZ �;�m��̛��ܦ�87Q�9J�8�@��=-�6�N��|ek@�o��t%w�ľ�%�)�[�W�x��ܢr�Zhi���[R5��Gl:m(U2���e������ïm�8;$#T`�M�T������G>4r|A��xB���T�Ĵ�$��9�`˜Fc41?�+X�����mVO2�=n�ƦE�-WܥaOX�LK�6vr��j6X�'[v���f.�@,�x����V�tC�=��^u�g0A`�,w,�a0�`���+���}�F��jP�˛����&$��RB���%�5��S>�y�V�Ý�	��мq�rU\;X�)9Z�������d3Zz��ʦ���J�wO�*��Mđ�����7�c�VpR�pFyl�pWܚB�˻�U����LTǷ�[Ѳ����W:M�!�͵��qܩ!y+�M���V�H�����B�2�X�kyZ�+7x�H��q�Z���[�������Պ���f��ԪC0�4�}�p��BgמtwĻ�ݕ�`����C�[�<*��.�ʇ���j��h��Yswh�\�#�ޝF��\��6���i��.d���r�xy���F�Q��j��[\}E�|
/��#\ڑ/��{���j3x��5M��k�x�� �f��(ǁge�~��3�:eH��)uu�t���겇�����+9�uv�Ϻ�O�jpn�B����\��rRuU��esx"�Å��̪���f�Ѻ)�]��E@�/V�����;s�;sf%=���߳��V�8�]��XC������7���f��D�A*�(�X���>��tC"�\�f���<�X.����Q��E���y�����᢯;��=9����i�.f;�eQ��h2L�!��|Ҷ�Q���XB	A��t���Cuwi=l_ϭ�X���bq�/�cf1�n���;	k��:�	������E��a%9�7&��Yb���z/�Q�-샢kb���^
�p�����zDe�w��y��V�$V���l��h��	��,tu���ɽ[��7N�P�7�7f�A�\;|iVtp�t� �~鲚N����h7��H�i6aW�������$/C�}zZ&bE��N<سog�[,�������Z�ru|�	r�wO�uY�7��H�j]�p�;#����iȒ{X:��vk�X�È���=d�g8Y�\��j2�hu��`�/z��`�v�B{K����[�	&uЖeX޳}۰]�O	''vk�RofeV���ʡ�]3�wt�S�i񛮱*��8�7����9����y���J"ݵ�;�V^k���P��"�Sj%�S��s�K}��"\T��*��ƥ^C7@Gպ݈Ov���ٯve�]��-��e�L٨�#:���j��C�9��3ztv+6��l�*�����3�Yo+�({s�:��[�9��Υ�����}(�Ll���j7ޛs��QU�}��=��#c���Җ6�ݐ���"���N�oc��/Rʇ^�e�]Z�Wp�R�$�<\I�����k��%}��e�+Sn�:�x$�g��"Y�w
Ba��ɱ��4wZJ�bC��8'��J	��>��i�k#�RӻK$u��)���7nb���m��`H�3�0Q�-j�KOIӊ�)�j�g�E�7�t�l=����b���=�9!t�� XWA�t&KkC睐ӽD^�N�@���lw$/�Vɫ�(�	>�l"��dY�]2��9+��\�A}�����Yr�n�dԕ[�3	=�3w�E����r�hY���s��έ:7EKx�qiL�v*����Ӧ��X����`6t�p�x�.��p̩�C��nqd����"��d3^�/�﹯;}���ۧ�7�J�E�a��C��iN�S#\
�� ή��R����}g�<8�ҫ3I���:uwy��o5�SF��e�2��m^R�A��:�p���"mh��'8z�����7yB+��lG�E����s\�GT�V�h�}��Nv�XR�����S��|PT��Y�y��1��тM�ƪ�vi�j��P��	�-�&cw�KX���Ǌ�Y	�K��VОxW���;6��K��f�,o+�rwr4�p0^�E���R+sQ���Y���ފt��%�m�hU��A�ǻ��J�9i&�K�7�Z��
��7��F���*�ޑ4A̝�����-���u+�jC�,�[y��e
�'-D&����;J�͛�p�E͐҆+���y���T�ZE���ܤ�tǖ{�]��e�ۤ3%����݆Hב4�庲��p��ѐo8s�r�B:�'�*���ej����avԡ¡��l�m�w�px�ua�
#H�vN�v�y.Cr$�h��-5�Vl����(�\��NQ��jKA}�I��Kp���(���ʐ�s�_}W���3v��Z�ql�[�smЋ$�B*�.����Y:k�6��!ݑd���p�<�Ѽ;xờ�%U9���ʶ5��|!�u�"�[�Z19�ȇZ:�v�\�wE�ek����N�'S����.1i�1;��0{��炱���U]���B�){O��(���XҖ)*ǰ�C5*��莢heP��-��أ�s(┹�BK�M
���w�����c���5������e'��e�u��m�T���*l<��6������s&�D7x:[C85J�+x��,^Z+qr���U�-짏]ּ�+-�(�/K����s���y�)��Id'��^�)��5{�7X0ٽ���s�$�����=����g)K뒮nӅwv��I]J�%{;-W^��#�Q�J���F!����l$z�^c��']�7X&P����8�c<������8(ܻ56R#�4,�Na��t���v'&v���˛���yx��,$���y���+)�8��;�ķ{D�jʽ|e>w���ŭ)��f��rK���t�M�Z�y8ݮnZ'��+63EM�B�^�x�,@���TB��Q�ېG�j<*}iQ�-\������:���J�ō�N����!Ԯm���[����U$�["#��NQSX�n���Z��}J��ø���S3��p���)�tܐ��}!1u M܃��5�)��\�`��NJ��i7�>���=�b�g*hm^�"3��6]Cڔ���[�8D��<��4н��Y#E�}q�V[y//�J�()���г�2i�W�[�������q�Q�ȫެ�|'�wor�f=į�<��x�`�;�[��3����ؕ8�'1���G�=�5Ѐ��ٌ��O�2��%��Ne�w�>�I���6c�j�~�85�]��m>,��c;2�gk��6�f]�� ]	�!��r�@ΝV۠h��wqɽo'TnV񙙐�:���:7r��ԣ8xfIJ.�+����E1-���j�e���b\%��Q�D�ħt������k� �%i9�E��{c���.Ԓ]L�}:��ܨ;�����	wyL����"�/ϨR���_5��=�G���l���)בzZ����;���ն)nq=�=���t}���_e�:-��Z����A����2��Õ�W �Wmp<�2־���������\,���r�b4��T+Y$�����PSa�r���ے�\��&�2ism��]�O�%��d<Ⱦ��Kut3`oo����#61��xa3��Y�lT��1�ɽSTj��i�1��6켤�
%�@<Rp�̄g=��s:�^���tt7*�J�kr��Z��bm�Bml�"f�H�k���樇qD{�4n9|����=R��Q���Vfv�̮L�!���[�hRw��˶x�r�x��6��fD_*��mr��LU�7����˾�lT�xfT;�4m`<�-��Q�Nֵw�%�l�(V͵����&ŪEݗU��Nz"�k��t��x싰�t�v�-����V�=�Wm��J�N�.�s��~��56z���MP��+%����/'r�卲��:醡X'-�[fC�GؼȈM�Kջ����+J�ź
�"�N�ov�s�ڢ�nhK�J�ۂ�6���;x;���լ�V�+d[��Ĵ&!ej0n�o��{�l����ܥ
ĝ��DX9�3M������p�c_d��+j��e���]��&�)><�y,�]ˬ�t�]m��������$�ܭ�\�8Z�Ip�˗��v#K�st͉�	p�-B�K�����a�*T��I�`���4 \3��oQ�
�L5Ғ	<Yf���৳WuJ��/
�vr��I֌��RUu���e���.��VP�gF�SNa�R�#�Q���f�[ծ��w�eˑse�u�2�@��6@��Z��8t��rJu�sL1�i����-tF����#�:�G�
�~�9��wM[bNM}b��1��#�G�(Y6AK�b&K�l&�����;�����[6��Q�}v�I��vw���W:�;�b����H����� �YZ7#b�	u击��®���7�GL�l����	O:�F$��6���%%��b����_s=�p�GlK�X���䐲���'1����x�B�\t�gd��.fɋy�V���%�i���_p�&B�	n��&ƃ�!�ː��'����aּ�o%fA3�sjSSky��<]un�mB���[��{�^�����F����U��@�r��ˤ��2��ت`��br��۶�S�ɻ�8:����D�:Ș�)ں���=n_v���Mu۬��F7bȧ^	�.��!dp�W��w-���}�;�v2�]�d�]�D���i�!@�v����β���N�)��KxVS�u���] ԋ`;�^
��sP}�c&tF�a�Ύ�P�D�Ҳ'��G5�%g
*�����k�d6�W���{N�&�f^�����춎#��ά��bU:�[7i9x� ]U���]�3�v�B�n⧓P���[R�١a����� �ݜ�t�.��W��o�<�څ��%䵏����s	�r�%�m���J�R{x�.n����Cjq�o����5���	ym;Db5�7ao�(�u��U]xcZ��l�;�v$�E��G0���fĮ<��^�zҹIA�UR�<e�R����y��M��;˜n�"�ͨ%ެ3\�jv��7N,�Z���s����k�$lB&)yu��]���y��I$�Ih-�6���?=�N�~K�a(��^phS���y�!�����������r�I�p>^B?�a~y�h!~B�n@�<��� }��y)�W���%>�_R��|���O��?!^���͐��y��>�����G���+���P�?.��!�z;��<��y��/y��w���<�!���UEG�������}��]��{����AEG�������߽�����{/U))��d�+��>��<��wN�^��{y����8qr�a��5����7\�{N�����YhnQ�.d�jv�� $VKX�v��)���Ӈ"�o��]��S{�骼�r�ޱ�RnYv��C��;dN�X7�@��O0n�VA6�1����p6�@կv魝iGt�ig��#�5-H�[y�B����KSɨe�c�m\�+`��u�e�tɆ����hgV�	�^�a�(�	�c^���q9���"^���l��.#�kĢh�
o	��X�{\��W$ѹi��OѢ#�\L]�ïM�,tk�q��q�a��2jEJ;N��s"��x�e�_tS�U:QuV�,�SRY�e��s�9(�U� ���R�V5�K6vZ���r�}|����.���J�/�(�]f�}�'�:]�z�]n�ftio;i��f�J�٥�Z�t �iJ����]����Tipա�wj��ja�m%Nѧ��n�sx��ꢻ]�ѭ��dN@h�h���iޕ���R5��v;1�я����ub���ie�;H�F�*�B�R�A5�����ڊ��	�\�z��I���XW��G)�˫����;��fv��p�F�+-��x[�zP��I�&m��Ek�a��}P��6�\b�>d�k�h�|���A�e⪵�^�LhB��Ñ�����߉��=|oǯ^��^�ׯ^�z�����=z��ׯ^��G�^�=z����ףׯ^�z�����=z��ׯ��^�|z��׏^�z����ׯ^�=z����ׯ^�|z��ׯ��^�x��ׯ^�޽z�^�z����ׯ^=z��ׯ��Y�ׯ^�}�z��=z���ǯ^�z�z=z��ׯ^��sׯ^�z��ׯ^���g�^�g�^�z�����ׯ^=z��ׯ��^�z���ׯ_O^�z���ׯ^���z��ׯ^�z�z�랽{��{�ޞƈ��c�K$]��O��+�d�z��L�}Q}a��M'N֬;2#���1�|	��r����֖u�FL���ܡ6��+Օ��׻R�H+2[1�j��h��>����k!�t�I`����j�O-�R�n�X[̱���J�U"Uη&��x]2K�ϒ҅G-�|og����8�kv�c�֦L�z��N�k��:R��i���oF��c�h��
�nF��`�o�b�*���;��fb�#�\�s�Dv��˒�[s�WհM\}ɚׄa�j蛶PL����{W:��+Y��m�`�K��*#j(&L���]������fb�;�<�z(�G�;��n�d��i���[�t� ē(J�~��e\뷙|�c#K��'}�,8s�g^�jli-1E�O>�8�tL�n@�u��x2���Dq[�b�Y����hm��s��s�%YƎ��#/��k޼Vn��{�fN��[�6��L$�ى�F�v�2U;L`�O1L7%X@�Ŕi��i���Sޣ3^q�L�<��a:EAfR���I���ciՎ�����jt
��ooz�.�`U^�Iܗ¥���h��^a��]5�k��\+uJ�x�B\i-}���" �t!�q��r�W֫���gE����uv�N;�(�|Ŧ�iӣE��u2�W�։7�C��S s��[]����}�?����z��ׯ^�z����׏^�z����ׯ_�z����ׯ^�=z���ǯ^�z�z�랽z��ׯǣׯ^�z�����=z��ׯ^�z������ׯ^��ׯ^�z�����=z��ׯ^��ׯ^�z�����=z��ׯ��^�|z���z��ׯ�׮z��׏^�z������ׯ^�}�z��׬��x��z��ׯ_�^��ׯ^�z��ףׯ^�z��ׯG�^�z��ׯ^�^�z��ׯ_Ǭ��ׯ^�z��{��}^m�5��%Þ��MsuK'�o��f�7���:W;�M���5]6+����-Z�#�OM��+&h������V�'$�k��5iU�k���g���|��ě�j�(�n���j���"�-n_Uy�g�P�'��J|Q����/;3�0N�]�Ҳh�Q�K18+.�uK��˛B��Z�U�S0l�b�����˭=r��I�uYY2�9�T�'"��'C��p���d�|i�/y���(�lm��Ty2�U���ʲ]�������Wy��N<�M�5��v�W�C���3��׵�5@<6I��;���Y�im���j����o>�Z��
����ف^]�O'�����7D�hn�۠n)vxaY%m���ͱ��̃b��]]p�[�gGN��[�^���1�D����r���31Kw��M��u�P�|go{$�;�˅�Z�������3Y��;�}n4;�tMˇ3� +����Sil��p�)	���uTj��MӶ7O\�Xsf��-@��b�)�� ��FK"�ݔA�i�c�{����
�xu:ȒM�*�U�мc��Xz�_9,}�&�7�H�����]v¡�7����P,�|1&f�.[���÷{��{C��+�y�~�H�L�V%���妌2c��U�W�eA�[�c�a�ǳ�C�����sx4�. �ruU�r̚�G��J�}M˽��0���áN�;/�tړ���{��]�:?=V��BPYz��k�E��8�G��!F���s�:]�M��7ZL����ߤ)���q�59dM�΋���)N�g�t����P=+2:��4��	IE�|2d��]!Q���qY�k���Vs�b��d܋�#� @k,�xz]i���㉍�b�YV"}���A�pb+����wG,}#�Mh�5+P����q�ms�6���(�#@;��*,Sy"�Yw8RoT3��]���|�Su�� �c�kMS����x�_n�[b�)TZ�T|�R|8PrU	��$�![I%X�R�2��tY��ܚ���.�o���^c��SjN�@�yW�g.�7��ݕ����e�أ�x걢��v����vZ���L��klvVN���^E������GH�4�8s.�1��Z�.J.�crJ�-v� {�w��i��B[�d�r�^
;r��B��4�f�6��Sg���L�?8�tiÝ"S�JK�c#�҃�c�G�:�*�Esqd�n�2�y��R�/�	t�^Z2_e��y��ns�V�ML�� ��x.&+�r��tF�'���[V�f�:�Cu�'���*���ȨQy��Q5KS���4E8�sU�wO���-4�V�T�,��g(���1`K�T������s���7Dס�V�8+h:��Q�3�O50z�êg��e�)�s1{]7��I��x333o
#���h�0��<�yP��AeEp��5׸:�C��h��s5*������ٮ��)�e.r��ʦs)�4�2�(&�����gV;���H3��:��V鍊ZAU�:0'��6�WImk�$L5]��w-�Zzv|)7��u�+FoȂe�9��Ҏ(û���&�,Ÿz��+!���"�P�Mws�hQ��Cz���Ʈ�r,ށ��(�ïwD���U6\������cJ�V���s��)�r|�Uu=Y�I��C3c�=��]f����F
�2m�P�4�����j���oL琳�N�ӣఠ�u�fԯ!Y �f�8���(JƟtk���rr�m�G��9��V\ӑ�e�D>2�=5��9�"Y/(��V��%;�
�*�S\.�r�b��2�9�ˀ;���Tb�^�I��R�(h��	��jV��wA�v#]�V+�ܱM,���̸�[��V���J����@x�n机����,==G r�J�tq���Ҝ��QlcX4�B����J.���eshPSi�yG���4�@�g.鷭$>I��,fY�:�Եȼ�gA'�Y��D��D��]]�;g�mՈ"(��4�8�����(Z�tڇ8��sQΩ$���tT�����D'���.��G�]����]��!�*�}[�׊�Ia��C����9Ƒ�m�֔��[S$�\ub/;�59J=�`4n[[�2h7�
Y�9usVm�W�m���ˍ���(�c�k�}�I�����VV��V�OA�M7lh��P���d�Cb>�Z���Ir���&��Xʮ��������*.�"�z�^��Qw#ٶ��&�F֣N��6�`%͝�Sn��&����j�9��c'k\������y���>Oo&��s��s�7�k�*!�!��G���fWT냆��;��'MMf��u�m5�����(�.���k�x�
>��O�G�_f�/ǵj�$��֌
���e-܇��L���Ӫԙ�%�=�fqX�9n�6b��5|��B����f��UF����vd�Xվ4^E+el*�����i�ʔ0RK]V^��Ƴ>��Fգ5u.R��h� EC���A�Is�2l�7,���`r�����D�GU�q�+mYȫ;�Y �TWf�x�^�<�w!��.ᎂ��V�Q�7��v<��Ul��B
�EvR!#1<I�j�ˇ�+��Vdlf��x5�ĉd*	f+W|���u��:çם����C8�.�F�-<��5.ܡ���1�Yi3·[��E�q;}��9�jf�5v!fg���$�{��xmݺt�i�=9����qr�8�݌�q�����V:V��[Xdet��n����V��*\;�)�*�K��s[�#k����'�G5_U=����836�q8�eiK�cp����K�M�̓E�Q۹n�ӆ��q�����Ζ��c38G�uQN�k;���VX�a�"��!��6sjv[{\&��t���wk�2V��!��]<���4�\9��u!��td�[u��-,Z����hv���p��cU*2Żc9͗E��v�m�o�\��ӤӺ-ҥ�kK}�c�>�l.��Xb����� �g*��QE2 {��*��L�t����u���:�:k2L�%V��q�k�9��{��/� �Y�#{GEt'g=�i"yv�V��=$�)�qXQѵ�7��zh+Xs,�t(֍Q�4֘��뻍��r7f�E�{z>��x�M�����=�<�:�Ҫ]x]蜎ƃV�ƸIWc���N���Xv��3-�s�9�����cݛ��ކ�2+so�Es�f�L�o
�QI�C��ڱ+=�N�q������iw*�-T���Iie+f��{N���bWKT&�ül��n��[��&.�R���j�%Gvえ�"��Nr�#]<��������]�OW�K'>Q<3d�Ah	��z��Q@n�������vovvI� С�|�:{�<��N���U��L��5�����妲�X����;��<mi�ͻhS�̥��Ȧn\.�V�lM;�%��7�N%D�;�P��g	lY�WP��7��%!�U]h�������7����9:��#�^��3C����#�����k�̳�+}��U�{�9>"�_oG��,;���i=�� Խ+k�8��H�ϴ�,���U6��s7��'`�/:ރL��u|��ŗe�O�ع�{���Ԛڦj�X��5\�޾畎�7��O���n�i	��O���ڄZ`��9)��v���/F�5���wvK�o1�b����f�9�ېQX�[�ri���v��i+�[����ݽR`{k�j����u�
�;b�)���'U��YE�f��%Ǽ�]�	�cLV����Y+�C&�KY7��"�������iSF+m��Cd).���άˇ�<�N�ʪ�uE�hu����aD�*���E����Hч:�`��h��n+شj�n����5|��'E�}Š�Q˅�uB�c+kv�e�����h���( ����-F��R�گ=��qm�}"�;�Ӥ�]R����r��+��kS{vK)�p�Z1K3vRM����!�\�E2�w�����s��ޕN6��D�.тv�ܰ�웅�z��Ⱥ��:L��6:�VN7Bu���-ͺ�{i�B�r騎��X\j���Z7t��dX@��:��@�+9.��rKX%�Q-�՛��D��Ɋ\�X�o��	����}�N�rUgQL�a�uCyd��� ��T^!�m�1��ll�6��ō�&R���ݥ�^�|8�����-��(̼���ݼ*m�L�t�d'r�ӷ{	��u�LV��ەA˺�(V^���p�z��Q1p����A��\�Rv��U��9�j�t�<߬�&�A���OJ�OuU:��nX��ؖ>r�W|��u/�����};q���t�k3���8F���9mp<��v4���oL�UT�/�ݭd��3k�&�j�0�%]^���gٍ��FB#�p!��ո9�m��3*P&��[�+z��9�r&��Dӯ[e��P���Nv������r��ّ!�t��;^lM�lv��HJ���zVp��襼���h��
]
üq���A���2�z��l�c�}����w��V�t�䥙U��=���yV)�oa���ő�{�{z��$�n���ͩ��;�h��ʰ���,L!�}�J���Ko�<��N���3�q{*8K�Ҝ��Ҁ�S�̎�zŘb�T�9��V�k�c\�y��S{����ݨ����r���>��Zo%�٢�!�mk����m�T-)��NX�J�3�gr����=+Bݺ��h�l]�-Yz�j�
$�M��uѥ�Ƚjj2��:��-J|�Ho�kUEXw�6��>e��;�Qח�����ʟ5*չ��2�*5��Y��Q��i\�.ż�A)�y�")�x��Z%G��(4o�4Q���-�-䓫����DY�uW����EQS��)B�wd�}�2���}WAXngIR_W h\:�m(Fs���Q��G9CZ,$�(޼� ̬����/������|�pc}g�y��ٝih8�'�D�@WA*��bY� �0�:<�x# ���K�i�t>��{o���[w���u�1�w6����>F�f��k�6�cu�js�x���5��R���N*(f��Rj;�1��2⻱�a�aP0���S��Dn�xҀ�=�{�\2���L��U�1�hڛ�e��fW�����y���~��G�����ʃ�����������W����z�7��O�b�{K�J�q��;� �r��)6�!?(S)BD�Qm��?�J�S9!��Rt8�)��	(eI��tف!#H�J��`jH�N�("S���_B�"J%��aѠ��H�cl��`��h8�h��&�B�.F�18��	
����P�V��T2F���?�"�4�2Ci�)�
&D�l	
�0�I�~D�`�$Y(���@�e��g�N��[��8�<*��kok�υ��hV&��:�3n-�t���;�MvG���C1��,����8k�^�[�)5ՙ�Ԩ��٬e�Y�&=�&��Ժ�V��"pU\�v�S^
�`=�M��������Bf�=��#!���F:n�Xt6�'���S�od�5aك��0������v*m}���ʸkWt��scN�Ӻ���ʦ2X���DKMaq��,HOV�T
9��N���|�ݡ�z�iO���Gr�C�6d&˽$ U���\�覎f�Lg�v���v��\�Au:`+˷���f���W}ݳ.H@�
��ꂶ,G�.��^9&����(P2�K(]%�j�� ����W��ii#�u�ǐ��x��A�2�g[i)���(IhjS,�]���9�9\g2��W��X���|��-�5�v$�WXٴw�����.�f�������$��k�~�r=��'jU�+oG�c�6a�^ncs*�&��Z���zzuH�Ƥk�̸^�^�t��1�y��]՘I���z�M�̹T$/��P�#�뵛�p�����8J���:
��,N�f���>�z��ړ��z��=��ǽr�v�o#,B��t*i�A��e�����95��p7���PH��&BqHc�)	e4�dF\[I�����0� �`�����8�B �n�i'
���l�K)�х��	�4Z*7P�%�i��2�,�B50�SF'!!$���&DI�e6\�����	��e�M�Z��%���&\R$�	��ܒ0�(Ě���
��ӊ?���!Ɠ�$b2�FRD���H�a("q��0'�S0��a�a Y�1iH!l3,��!D�!�P7$��~���-��
B�_Gk�a8��A�2�-�dq��D2�0�E��I0�)IiB��&b6������,&�QD@��ȢYl��$L�f2&)
C$%|���	���T|D�aN/��&SP �d�DP�ځ���F�2��<ݣY����ꪗ�Phڼ���1sf�1���"���}��O���ׯ^�^�z�����}>�O_o�=l�gkAMEF�&��kl?,Tm��l��7^�������ׯ^��z�������}>����t-<��܏+��M&�T�IDG6<�f���-U!W0h����O-��I��W�6�����u�+$���)9�O�.l�(6�<�'��
<��j���6j"�&��TD4�LP[�Thѧ���s��b�Ѩ��h�Zf� ��K�/,��^[��6�h�����HnQ�F()�h*�;�2hNMo6�yy�A�Lsj (J6)`��j#F9�xR}�y�\"_Q�r�G��:btѶ)<�C�7//Wњ��r�d��<U���fw�\ц5�����`��J�ss2nn*�����`o1���Q26JD�ڈ��$��j�-��7�� ���eDc��&	~��T�(1*R����a���CT�M���\"�W���K)
��'d1J��RݙQh�I+Umq���y��R0�&�-6H00�AHHF�4L2%�h��D�0��f(ې��I��@��Q�E��!	Tk<�~�W��L�{3�+$�᭄�L*m��a&H�s19E�m����J�=�ɖ�EX���1UU��s���<zm�V�z\�q@��'׻�x��blO{7�=��ۿF�^��g}Z7�������=����B��������$��H�&�FNz�0�w7S����)�&��H�M�����rN����hT��k����k2�>�6�f�J�������0���3�+t��_��7
�ܓ�S�g�/$ɕ�R�+����vt�l��3-30K��d���~"�^gl�O�[z��'�|w�K���5�����Z�*U^�^�ް��~�=9��[�z^o��ﵿu�ЛD%@�s��h~�K���h�@��|�4<�7}>k��;$~~�����<���k�9[ݻ��w(��5�K4�*=u�^7�M�ؽ�3n��/S���>��x���׿~R��/��}�{y�B��f���a�Y���&�%���F��H��}p̭}y--�e�T�sj��N�������c��R�>�� ���1�ë�Ʀ�N;ZK�B�ơ�w�}R,���o���h�>���%<z���c��p�]��	Y�.^���6y��>���H�.�0=-���V������Z��+�8VU�)���^�(@�$��@���Q_+������<%߂�Zf���o{tO.�ɞ����6�D��P�rh��~]T*]hMW�w�U��{T,�}�Yrx��P�$_5�e�~���G��2����s�m�f���G,Q�/P֧�Μ��/���Gm���e��Poީ<=>�L�f.v�ދ;�33;c�􌡓�_�w��Qdw�u[�%R�J��/^�5����X29�L��&�>݁:��i��:��\�5�'���Q���7]�j���*OR��d�&<K���s�هT�$f�9��p˱#���>��'K�m����T�w��h�vϻ��6q���	8UJ�n�"�"_1W�%l��
_C��B��]��K�t�	����=Y�ؗK)�앚��)s�Wta��iQ5R�uIx��x�>t�^��.�;hJkx��n����K��{=Wc��yL�ךEP��e]u�$�<�vWMC:�R@�;Ӷe��N��ҫ}~�_��9����o)5�@�����c�V����� ��$��w���b�W�{;m�s�{���4�QX����U�X������r�����ۙ�S�z�8���}�f��e����Pn�p��e���1�y��������M�}���&��y�/�m���>P^�,�.��LWok'�CbE�Z���y�:H���^=��/�=k�Aу����FM׬��T�Q��'�1J�S�^���3��Gb1��E? �	�W�;U�vu�:��z�}��}3����.)rW��p����չ�{�� ���a*E���)o�f!w��o[��{|3��W:e��35��=����G7�<P75�W�ϩ<߰��5�_�o��=C�����y�8���x=1�軠}�tN��햦O������zT�V}rr.�|}6��f�W�_�[���lT�ޕ�>{k���.����&pr�GZ(�ʹwv��:a�_�I��/�}}g�~jlË\dqB�+���fV�k���� ^����Y8�����U[��R��ɼ�o>��8��V*������'�8ښ7����� ���)t�G����7��%s��E�i���I�~n>~=-�u׻�����Q�$̃��3Lޮ���nի�k���>�X!x`��D�^�l��G9$��M6�>��
�>5"K��<��Gc�!�RmP0K�Ůf�y�{�OOm<�}��RD����v��z��=+���g����O�k �˱�6M���|���Yh�vi��h��3{��c�^���Q�+���7�~�-��^[Nz�Z1������=p���'�g��3�X4Fٶ�d�/oF��୛v��o�]D��b�l)��<���~�bSu`{@��wA>�u>������=/�g�����~羆sb})��d�;�x)����.UI������m9c~���w "zoۃ�a�X׽=N�9V�j=���mw˖���<k����	%q��鵆�Ȕ��ߪe�[��3j�F�i8�����|��׎�8v��I��}��4AA$p����.�f殫���u�z+����b�z�S/k9��$�0��\7<k<�y�k�y��N��'QF��?w��}V�>�j��1��;�x���Bm>�����.:��)�Ս3^��D���
�}3�@�PD�o�Z��{}ѽ�V��
�{�n�;��y��T���NW������ {����+�_'y���Ŀs�D-�n!��zf!C����gҨSg�|�_ ��@�O?>���9�	�Oo��<#Քg��vY�s���ۇ8�;lLo:���2,�z6�Qᇍ��T_����vZ�e�9{Պ��p���|�I�]�=�?}�Ѝ�s�V��C�=}=�7�=��8�]���'kw�=�7qNEuy��v\E��V
[唠�EL�	�O����3���SF�i��܌ ?]�ܷ3V���M�p5�,m�n�%Q��^Z3ow�������*��:7��f��z}���c��l������W1/F��	;}�F��x���dq9ϲ;���X~���,yη��l�=�:m��.�1�|�d�z� 1�=�:�]��֎�`���R���j}���J�E����r��ZB=�*��Ȳ-05G]^L��`��Ge�}�-�Ұrfp�)��T�b�Zb�o���rE��rnK�[iT~W��`�֛����}�g��g���E���/�a�ۍ�(w�i#S^5pR��y\�$|���w#�IӦ��u������{�̡�����Ev���z�7r����)��ؽ���	s�H���3 ��If�sf������&� 7w~)}�A�G��^�B��{��;�����Um����x�������rm�M/��$J!K���~�,��t�)��rO�{Z�M��#������>�����R�~��N�����5{��z�HT��N'mf4@���3��������&��]�����Ʀg���#�Zs�I���=O�����d�5;C3 f_E��h���_j�`w�c��=Ygr����o�|�ֻ��YĊ��:@�P[����ݳ�;��<��ξ�K��۾��c'=-O���576�� �ؗ�ɊI-c�]�z�	���9�t�Œ}�p:iًٰx�ΫA�w�d�Ϩ�L��pY�]t-KB�a�5>y�uB�Ы���;�x��1=[Ƣ�}Y	|�PO���6s���F���o!�׻�y�;l��2��W�̾�Ī��`�W��}+S�]����b�����>ޮ��c��/���D��]���34 $νh=ۻ�7t@`�%0��'�~�Rۨ���\ߟ\MK��Ǳ�3n�wX�p"�n�M��$�$��>ދ�7��ћ���È��}�c=�{��	��9��$�͜o��{�*g����jHz��2��j�H�䗻���@����c���o���&y��fn=�K�'�rOu�����>�p-Y��'�-���}齋����K��t��[����ԗ�ާbJZ_>�%{�㯰2��ީ�ׇ��:��[��qMMLɞ3�P]��~� r�Ї�f���HT�S��E��"C�=~�<W����ݎ���S�� ���fx+gt��ݯ\����7��RƧ�}+�f9Qd�1�`����ZN�f�����^A%�;p�v�=��h4X���|�	�m<���o�Jm:4���Մ*2�/tK���ޭG�����Ԏ�{�!����Iŝ�����p����Jܢe�Iw���j�VGo5�޶�2�H9l�a�M���@?����>�ci8į1��`����bF�k�ϤɟH%��C�!���	�o��C��yLQ<��b��}����Ȓ��p7 ����P�z�#/��Ɣ}^Ǿϕ防��=�g�߂=ޜ.�ܞ��-���/'�'��.��r�k���ܯ7�tN��p=�[&Pс��ޓMl}Z���>�;b}��Ogڳ��}����Q1ʟz��ӣ�a��5�$�i�n�ن�[n��r[4��$��< �����X&i��Cy������T`�k�>xVh��v|�I�~�I3�{��ޯ��ôq��H�o<�Ӿ�"��;=�={��+\{�cs��n<y�^�S~+���ztط��s��6��N��x.�������������^UyU�:{ޏ����|�{���N�i�x{�o�=��[�M�9�)If�7�b�'�W���a��<�`�du�:����Ec�[oWf.��ޖ,��Rm�W�v����AW#�(�y�n|ԂV�ZJl��7nJg\�������4f��5��cq��ҧo��]���ut�"�������m����N����$�Ǯ;�N���틮��_�u�]j�pw�I���=x���ޒ�����s��>'�k��c,�>'����~��L�ųC�<�d���_?g{��@���`4BϏ�n��l��e/j'��.Yy�@��tY�ε�fˈ)�?zM�=��ՏE??"�?{/ԕ��~������+������5�����~r�Ά�zz�b͖�4d����(W՚j�ll3�'��`!���d����$��"�j� 3�:G�-�k�$6`G����9����z��W��`د�{��M���~�GB�2|�s��_�!��zf(p�~,���,LL�痽�i^�__w��pI��O�Xվ��3���G:���u=��vӥ�n�C��3�q^�!�dЋ�>U	7B������z�ƕ�s����t��ķ������`�/o�f�t;��Q�(�х�~GX`.[�����,�iN�K�p�����l�y%o��>w>���O�C�C5�����!&|���7�Xὰו� k�	��γn�]dʕ�C�n���Q�O��Sr1�ڝp-�u�W#�0�뺫�#��=Ή�ٶ��d�7��ꇯ��p�MQM�#�����o�;/�6��,��A'R���Rnʪ�/{ޫ�����ܖ��z��R�9B�l7��/���"������I��mM��MPx�ޒ��nIpI#go�T|��޿3���o��'%m����m�\�u�����d�9ϳ��Ќ�����K��qB=�z�	���D�[}��26�bz���t�Ǯ�����׳���{��!?P��x.�1��Ql���J_����>^ܺn���﹧�˚��4(>���L�ǼT�O������_{��nzU7�gH%�^~�����4����a�ë��/_��>]0e�һ�o֗^w���G��zGb-#��!g>��zX6����K1�z��k߻�~G�|nH'!%��
�A��8C�_h�~���5� Kv~�a�	��ͽ�pj�Ӣ�i��ڂL��[x�V��j R���P1P��I������,�ۧ'(ʷ��"c�N��t��̫HBR����f���U`h%<ط�Xn�"�=Ҭ��FZ��"�n셴�b2d�w+���c*��FAo�н�
�S˷6���I��Ȭ�F*�s�x&򽣄<���	�s��{{�l��!v���Z�4��U˱��&��v�䞬���t��0�t�U.�(J��&�c�u�]�������=ϕ��5�(z�*��tS�հi�q��]�ݺa�����D�!&=�B��/f̬�$4�Fu#�-<�r��z%$�Z�kHI�q����<�9�;�J�^d5�*��!-E�n*5��ܔP9cMr$��E����0��0�mk%bk�w^J;6Uǃz␇n��e��:ջ77��,*�Y�"΅���pt)DmX���Y�$C5[���v���N-Ŏi�ф��9HmkٝR��Aɗ�"�B��	��kSnU鋻s)Ko��]�&�[�����.�3���^��_u�O�7gf�p�i�;����2ճ��}�Tc�֢ʯ�v�ycCO�b:�^�r��T�%�#�wZY���qr��p>�3%J[�F:1&󒊘��5�4Wut�8�GYZh�wFg)��z$�Ʃ���g_.1F��+s.6$l%T�fS�j�LpSVѹ�CΞ�o[u�v�$,Z�r��ޡ���M

~�{��ǹy&�4���4j*sf���;Lu�(�L��%�dm��{�^���\����uL�C������F���@�cP*u�e��]�V�W8�C�{��2�؟;��u-�z\[�y�Ӏs�&z��l[5���ނG;�ى�W8�<C��/����g�^�$m��e"^��8b�����w���2�s.�[TA:��2#h$2s)�Vգ�N��Ј>���w�e�<䪋N¾�����j��.�T�5q�G�^i�yC�99.�t�I�Ҷ."�n�w��ݣ�X�6�Qʷ_.;�k6?$�sj��=�ξ�UQ�����A��I��z{g<Ν&��gKˡ�uq\[p���Q�^ұv�0�D���oXpR��%�D&�7����;4��*4B�B8�J�Qܒp�tB�+�Z��� ��y2vL���֤�9wSs�廆��ܣ�����9�I�ϮX�8]���G�R6q�ov]t��1,�Ԯ)\�u��/I�NS4#�D˽p��vD�C���r�<�O���Z��Z]�n^�DɕOu�N�X ŕ���PŎ7.m w2md/Λ;��{_��DSǏD�ך���bc5�kk�7���7;���|�Zm�~=U��]�q���q�@��Q�������Aj��c����/2s���W�lpH�n��մs�[I8�������>s�kX�2θG9k@w�G�c����O������z��^�z�������>���ߗ�r|j&�d3l���r�4�l�m�^O���'�F���(�ʎ!:��q78b�O��<}�߯ׯ_�ׯ���~�_������ׯ�~Q��C��-��Dld��ch#��������\O8U�s^��[y��G�Ç�2�Ŀ'�B_��C�
�6�778�ŭ�Ʊ`!���Ae�X�4s��P^b��.>qc����7+�E^o8M�'4<����<'�6��d�9�����y�'#^1�ɤ�#o1�SZ���j9r4p�E��*��r�Q�S���.Qs�s��/1���nI�2>l����AO�����X޹�lAkz��Ά��Xl2I��A�j����$��6+��i���m����`�S�"�Ek���Z�lkl��g���I[�=xf���)5�^�Q��G�P@s�71��#����Ŋ[�������%�__�qz�]�æ\���e�C�#�Z"�	���N)R�ӄS��,��l��s���溓��^��g2G�}�����[n��k�P�T�l��:����݌`탺	rC�7��b�i��g뭳5^Q���?T%���M'���f�'ϭ��m�z�U�+�5�n�P����׏�A
�).�7�i�!�{��<��f�aj��ۛ�=Ձ�g��<��eO�>0��~��)z�>S�m#Q�jf�e����8�	��aI��5s��!^b=�>[^Ϟ�瑑N���m'��W�5���^��%6B�<�s����ޭ��{�P�m���E�*3�=[෫o<��p3�b��i�L@E�m=X�+�*;�߷��a�����PĲOa"}V��&��,5�+�R��c'�<�f_�3��HY�3)C��Ð;>I�\����>5��H�U�ʓ[q�<�"��t{�x��h0b�FGj�3�|�@��џK7P�Sq��I�;���ؼ�)7N���k��sQ1�㖊[����w%a��c�SAaA=�ژ�l�sIz�a�vAn���O�<�A/{v��[pǷ�K\�R�ǁ���	`??�����
5���s�ge�s^�ln�-|��Xە�]ߦ�x�5���q�O�T�2Y�ŀ�#v+��	F�;����<�I��&2$킦���u��:�K�H�*먧_K��yv���j-�b��z�6z���n�ͫ���]e�Ləǳ���y���x���t�}5�#W�������n}ݴ{8�}Jm��T}���e�3�t�b]��XQ��r���q����N��!�!'�9f�r�n���b3#K�_������1�Pe*#�A�t� ෝٵ�52��+���3ڇ��.�)���������^5�׿q��u���<�_l?ӗ�
= �AZ����g�*����{����C�&��K�|���>�m/�Nf�W��5� ���j/A�J\��z�݊��[Z��5���k;F�Ìd�v�7���&$���f-#�p���M����k ���b������5?�_ñ�8�����A���a��"��K��d��F�e���&v�~Cͪ-�7��e�m���sͼ|���;�."�����q��ܬh�M��˦��vC�Q�8�(�2j|}��\��lg�3gP�Ξx�xxd����S/L��nHxڴo{_)q~C�yL��V���G=?����|ŧ�tR�g࠷���*.Uפ;B
cwDw=gJ�g���ʃؽ�y��}N ߦ'瑯��=����1���Wαl�*U&ʞ��;?3��~и�6A��k2�Q���^��I]���yj�L]�OY�\QĈ�wuvd��-"��׻ ��ˢ����T��Jֺ�;i<݃�t,��|M�'
Vv�',�S��j���[׃��^F��e���9�sB5W������o{.W����BΨ�q�eɳ�����$���;づ*d����|�:s���Q��j0?���2.�9;7���`����	�{bS�Hׅ��H�@�:*&�f⏺�0��޴=���WE�*���HP ��q>�!���n��6wR���LV;<��w��%.փZG�q��O	�pc�e<?� M�C|��4kO��!?P�s͸�[}0���/ښX��flƜ�=�#����Jq�:�7-/#h�\��ޟ4s㼴 �7���n熄���
����]�V�O!�,��Jh������"�����߶�~M ��X��CҠ!~ v77g���vm��u�{P�a���_L��(�bN������]<�UW�X�G�]���� ��y=fӋ��O�U_���P����������KuL`2wE��`t�+�҂^�ū�a@�γ�3N����J��]؇������=��O��!q	�@}N�a���#rKj��jT
n�Ǐh�.ե��Q���/��7���p�Q��̽s��^�:��.���3��m�_��u� 3n��Q`�\�T�҉��˾gU܇���@�'�P��F{_���b��N�AU���L<��"��43Bǚ�a�����ٻv�2I�W%�1�����=�\璊}���őg�s�6�^S���u�u�GN$36��G��pD�,�4qs>�zS�qi�n��M��c�����7ђ�����w�C��_5�uv+*�51�+��sq�cd9U³��O?����}��������u����$=x�A�G��h����ok��0!��|����쳫�.3���؜u/e�� ��n���}*�!����0Yn���>�E<K,��b��J�����Cך�ෂA��L]�kܾ4����� �еt)YTu��E0�i��*kS�,;�dx���� ��M��6C�Ay	�P��ֿ<��`��L�֍xR~�ѭ<�����J�����x�\�Xgu�cռ4�{gd�_��/�1���3��6��W�H��]�X2n�^�#�_��L���IW�ߣg1����	�[�Hqm8	>T�!<�} ���.�t2h�Bܓhy��q�g5�;3��X��.���8�e�%I�)�Y
w0����H02bϽ6�/OZ�ӹQ^�wt���8�;"MvR���E�fpn�d��0����-A�6�z`�7��vTNB(�f�#�@ ���,fԉ����»�� r-?5����.�|\N)�jd)B��z���ܞ#�_���0~mi��jbK��T��;B��.���QWC��������4-�"��.���;�9��B��2�љrP>رBY�����n�П:ҽ���4R&E��|.�fU�h�}2%�h^h�����&��j�hlⷤJ��}��s�Q%�q�p�Y;�ks�`����>^?�����s}Dy���������Z`8A����0e��0�(�-L�����Ԓ�Pu7�g7܇���y�SV��#����]�hp���}�:�#D����g�h�i���՝3���`�s9��L�N���,Ƽc�k��]>�O���}�MrOGH�cɾ}/C���[)�3S)=�{9s3����3r����^=%�o�����ųìC���%�Xlp;��Yi�N5j#�3�Q�"�59�d���@^.�t��7k_��	|!��Ӵ���N����3�V�AK�F�Q���(x�3��KLzcV{�j�cv��7s�|]}}@���.���p�n�������/���ky~�-31B���Ŀ?���#~��s��X#RT͖0�[�;GEDɉ�K%nk�#�^�[gm�u�9ύ3�9�)��hh���E�9���X#S�^1|͖�f�(��*C4��/��,hB�Pd֌J~Tgz��z� /V��$`�as	y��^V�%.bx��t<]�B��P}��&%�{	�V%*Mm��񹩝>
{w�#��
u�b���ʴ'g��g��,�8��	�jB�k)��7Kr���gM{����7W��YNC.�o��v࠙��Rѯ9}㓠{�OY�������e)�E����{{yK**��2�m	|\�1[���u��p��Y��^�[�\���������m�bp��qj`�M��;dӷ7���9�K��H� �IRkg�m�p�:X�oE;�e�196�f�ǮC܀���`�fP�1����0f_v�$�p5�V����mי��e�2%W�uZmaa����<�- [!d6����^�ئ	�In��b���<)���}��k8��^��\D�u�*�3M�><���=>#����G���������Mi&©�ޅ�������\��q���8�jc��:����ޱR'\��v�ݬ��[�m��<qƱFM[]񔜵���=����q��n����@A��.�;;c-*��5ڇ��vg�צ���d���R�Xu'����?��@4��l/�Y� Q��Wty]��B"��w�9���P��󖄄[[" r�^��>n)����A?`�V�����M?��
rְ0���ݹ*�61Z����0F0�'Mq0q͉�����ۆ| ��ӿs����f�'����B������=��hw����ճ>4���X-�?ߝX���s{��̾��g]/7�ATo{�q�x�x�'���ib�i��,*�S񇇏Q�Q^�Zs	��j������Z�xۺX(����Jfw ���eE�H����m=�{��9�b�f�&UfʡҌj����V�Yч�`�������P������l[��MO(' �>��w?m3�cf�X7�d�����/��Ju�1F���?sͼ�υ;ǰ!�ok�����EZ�nJ-z�zua{e������r�W�3���Z�Y���.�,8!'���S[s.�@c��˵���sN��Q�9T�[N�!��	� ���1E�z:���D*��]�t��u�?ߏ��br_ngx}��8'�w�田�O��|c��mrہ�����(ʤ�d���ԌP��ʥfvl�C�X0k��K��!�z��Ⱥ	<y��o��{e73s�I��Jui�o"J8���QSy�zz�!�_��(R08����o@�c�@qp�2��`84�t�O��Re���+���3�Vjθ�=%�k��2(�&|Xg
��ZdM���~��?~<��喃(ծ������ը{	�d;*y=#ɼYu�72��6�Ms�w�~yw�vA�okH�!���k�����CU�j�ڇ����4��7"UvV�]��Sx��f\��J�i��Bxw� >;�ы�oR�1�7��d���@�X�%��R(�1'_��E�Z�s��X
+XH�����������w��;�ݚ�'�=N��i�,�7xl�B	�� ���q�ٗ�D���9����{ �tM6���&Zk՗OD�c9���a��{N��ǭ�z+�b�r�feU��Q`96X�XYw�Q�k9r�s�/U�D�pv�+fF���ߏ���Fk��7~��`�����1ng�j��>ܟ�����J簖zI|e.Z�׺���q��gc7�gJ7�2�����k�Cc�D����d��,5�v�@��w�<�Ž��f6�3��s��j�ͯ�3z=��^_���� �"O�ah_���ہ�0̓��f�m��H7�ݫm�&�:���v��`��p��θ�0^�3.�HD[��m��}�A8����H���ӋdH+�v�*'�����y�>5S0��^(wO�!�&��O#.���TD����#�������@�U*�k�j�����ݔ�Ľ��P��c����� ��\9�q��d����s���NvV����Y�3N� DS��8{�K�4�zn���JB�ð��t)�����Ya/Ş�fb��7:���}꘨��g�| לl�G:�=�yt��Sk�xJloX&d������v2s���=��t%vP��=:�֬z���p-��`���R}�/͈W�|Cu��sd[�nA�2�n0f��=���ħV���2k�J�.�g1�k�<'�kѰ�A�5�Nd�!>��E�k��3��B�=Y�c��R}7rF�b�V����A�|"���	��V�4�����c ��S�GfV�ѐ�Bce5��ҳb�1��A  N�5u��v�p�V�Z�f��#�H���t$8�
�o�c�eX���J����E�$�<��#MtԒ���	�������U�b���pGֺ�(̤�<�%�y2��T����� �s	�_X	�<=2��������<[XE:�A��2%vIoCo�"�����7(��1L���⽞��]S�*�RN��8��Z���9ܼ߫��p�f�r�`	���P�v��9��' �!t�~g��v�쩹��%vOV���a��jܰ���M�^����.��KO�b�?��=c0aTe��#��k��̫zrŷݝ]�d{8��h�5[�X��
I�0�	H�}h/ֺ�-�6KL�ɬa���P�'���7����=�{�r{��P4�u#htY��+�0�����|�����;iDX���c�f+����b��z����i������ܳ-���dtg�`<h�_a�/�o;����d��x�s�8
]���ٷ_H/��Ly�%���}�����8~EKۅg�]0��'o^o!�����\��J�׆�~o-���X��{�^�"=���_E��F�z�T���r����b�|��bJc���F���V~L�Sٺ H�Ρ}%��U�B�ܤ����[g��Ւ���-������ڔ��3Ee<v�D�F�B�5�W���,��dw�I����vU,�~w$�t�0tyy�è�h�+�V��D��M�ٸ���T<b��VK����s�c�1,tQ*ϧ(�mu����m��od�`���F����x�<x�QET�E�?^�Y
����p��sͼ4�^Y����j�	��Na���OM�Tx�4C�U�,F�<j���z���5gE0ok� ���8�n�[�}�)�08��a�yp ����!�!Ov���u�ob�/��f�-hyA�P�f�ߕG�c
���ޭ����K�e�,-�a'��M�]���G����`!>��֠� pN(�=�f�X��5؈�p1�����\c���Q����
����&t���࿁Ba0S} ��y��%:N�讑�Q�I���9�j�vf��%.;�q�@/hx���6�����0Y��}M$wQ��Q��]�C�J!eWmmdu��nN�s��}�]|l:��尻=�������w�3˳�Ch��/Y� W�r��A̽�}Z����Ld$����0�z<����OJ>�4��T'0!��߸��/y�6��=��ڐ���!\�c/^&;��c?��z����,��p?G�����\K���΄�? �״<�����7���MϢ�,�A�]�B1�ݘ����n`��@�����&�cW�o	�<�J��6�\yf"�v�<"js'��a������N���SMd�5@��ݚ���RW&�jի[F�L*��4���l#��P�R�RP�èN֧�vWv�~%3}�4P �]����k9l�8�&�������х6e�C�5�H�m�!��
{�u��|�������W��	���ZM4Y9�*��7��7���^�o�XŦ�vpD�U�9��ay�#�9f���?u6�T����AJ:��{�B�^�V���Uz�]�;6!+�R� �$Niޤ���]O�m��R]��0б�!������u j�K2�j��]an�����}o5���.�&�.����,7��}B<;��\�.�*��ٰ�.l[É��9�{����
�&��mλ�[:�an�t^cu~/Sy���Lw-�ӵ�W��}�(�\�0�PZZ]�n�c<I�#A�}A	5t�]�}ۃ���$])Vzu�U����?���(�����|ݮV�v�n
Qʘu1z2���ֲ[)��-KW��Y��!Yc����yVoOY���K�#���i����)Jb�ˆ�L�3�I�!V�j��E��X�����#J�m1O�*�2�����헱���]x`�N�8ok7Y�>amJ�x��ѓ3L.��푢���U��Ե�|N���UM`����\���æ���B��KYЩrn4xm��>�e�õB�7�^���>��p��ݺ?S�u*��y���|릫0�+sਜ��z��A��1T,hM�h�l{���x��~���W+��w8nVA�l.U����2A�oI�S�C�uyty_g9Nۭ��7�S��{�n��N�'D���.)WI�5*=G�nh;]J�U�.���j����MIG��k��{3[Z�Q�NKx���BTY���tc��ݛ��>�:��턭k�J��{�'��㸂�=�UW{�%�5E5U���q�J���R���qÉl�g՘f,�c�Hf�ᖭdhbȖ���w��U��0�;����˕��&�y�f�R�k�-p�Z^��$jK�ʖl�R�'HW���M���v��;��˧V$*��]_pX�a�8p��Lg��;7��6�Lj}Zl$�X�ؽ�slU� F�򋮦<�5~���FVVM�����TUE���D�qʼ]9� ����r.�����t҆�Ñ�;2v�&�L7���1Ќ�2G�('��=��C�������z�U:;���777' ɼ�[���jwQ�9{��q��h�)le򻛷���eH�g5��]Z��8�M˧�ԁ�	bd�:����MZ�dΓ�*�ץ��.�,J�,c"�q|vR+mc��.G�oS�����:t�G�Y�I;�^���j�,��y]'�+/h3wD�Z���oyFVĶH0�^z�瞏����^�k`�VՍ�t�s���/1���|�7�O/��ǎ|}�߯_�_�^����~�_o��������{�G�Ƶ<b ���^�8�&���Q�*�����|x���ׯ�ׯǯY�ׯ_������~�_~�/�V�t���sgDC��3G��Z[_#���6�/5�LA�gO4��X�9'���y�*�u��N���P���D�A��f��-G0��<2SI��*�,b�Edڃ��͓��@Rj(��m�B+f���h�"��j�<�D@E\����bƳ�2QZt&��Z"/X8\�X�A���b"çX��4[$m��E�D�[a�(
Ӥ֘-�q��jb�H�b�Nf��<�O6���4TEͶ��$ֱ�ƸN�N�-���[�"֝�+:��t�fٶ#glfh4�cd��m��^�����q�	)��5�H����YN0�-�1�
�A٬���O�ܺ�����$
CC;N|�ň,h�q�1�Rj�_n��ܕb��p�;pu]+�w��	_H�*""1�*B�01��pKi��
\m��9$Dp9$Q4
H��B�	��� 	L�`f�G�fY�e�_�7���G�����J`������ƌR|���b��&aF˖^Hn���O��� Q(9�~?A��z+���mv*K�a�Ʋײz}]~5\����ݙ}p�9�ג���݂���2����!1`&4a���/��h?Wm$�ݨpha|Z�x�朗n�'x\�յ4���Y���gO<������,	|ܙO��>(�~08�b����n�m}� 4"��/�<F��4�������z˳k ���q#�E��y��["]�om����1m���w8W���"�{�M�Q0�ocp����ޯ	X 9��]�E�ǌ�H�ִ��6�v<%�� )f�%� �Eږ2���q�2�%�Z��oO!�o���{6*� Ũr�W�3���l�ێ-�?4�Ճ��Gu3��e�Ui`��m.���S�b��uA	� �-V�K*�F������h�aSr����-6m��絻���x3w�Ф-���>���^�`�5�K�u��M�r�0�ē�8D�$����z�s�B��pٕm2����+Y�D[{|�P`fL,v{�nP�[�� �'b�[mP׌z$6^Y�i��<M�܎�������>�h=�� �3�	�G��� <^�j�X{~�!�[��Bdy+�6�_���ޘ~���F�T&X1֫{(1f�S��0Y�^coS|�Dt��o��������ל�*�e슈��s!���s2ڲ�T63��J�Bj����u�ڍ�]}|�� �}����z<<��xƂVj�%���<$:�ԉ��k�8^��m7Z
1���S ��5v�Ot��(����	�Zچ�E�|L�"����q��Ln�t��:	q\�@Qc�AkڊRN��W�{�=��P���4S�/)�:'�[��5w�d��W�\���:�]�xw7 ����1�| N4ҭ����{Ck?�ύ��`X�K�9��B͘��,����y���a���[�
�r���w6�e��`5á.5��T2g�Lr`kd��BՃu�c����-}	=��������8�}|WٽY�G��0��~u�{�)�@a���F�g��L ̳rKm�P:Mu&_��K0�W�`�w!�.�N?s�����y�����lg��O�I��	��&��X�fM���L�9D�`���Z���;&y�J%=x��;�a�2�t=1��+�?#߇��yn�=ݮf\]n�N��#ų^�!	�;{�� fE���	E@A�F@v�m�F&���3S��4̀�ű��7�!���@\H���){��zj܌î\j�ʨo#^k}�M�ç+Kt��sͼ��<�K�EZYXۅ�ZFW�;�UϹZ?yO��;B��]���m��x_uwg����K3ɘ<4�6JE|	��or��hg>���Y9f�n�65d���*�r�|�;K�p^+����\�5D��Oe�t�6T���oW5�������{���z ���	$�������C���g���G0�a�q1q�j/r���&�[HԤ,{ ��t)\��/���7�y�{K�z�F|]0-��tS�~8`�����m���l;�M~�(v2WF�u�Z�C�{r|''�o�+>�1KTQyD;,�x@�O_�/諭��o�Og�Ɓ0N��u�d{G2~�7�?D�6L�	�IP���ǭ}ocBz�	-�:O��?<g��<�������~aD�X��c��3�؂\��%����J}��5�c-Y)�~���B|�� ��tn�e�بxN������fC�5�(�`��!�z�D���0��%��5(����PZj.e�DaE�Ld>ì9ݹ+P�8r��"p�f�BuLx���ݒ�����\��)?7�3�p�0y�m�U��~��<u�en%��&���G��!�ƑG1�=�tf)�mNׅ�*���C�5�3M�ޕ��{^�ج�1=��}�^�$����`�"�� �ֿTĶ7�L�,3[2��چ���9;Zuq�w�s�PK�<��5�8s�N�����)�N��9�?���- ݲ_^hP����C#�1k6�^��&N�C~9�TPO���r��x����ƥ^������i�V�nIp�f�c��e�G���블��{L��_t��'"0��
�S��]���L��hr-w��jb]q1-WW��|�~�}��z=�x{���[�{���=����z�M��ҩ1��S�z��O����4��,Īu��:8y�3�\Ğ��?���Z3R!�C�:Ǳ.��>��w'��ş�\�㰂b�y���-�b��<4�<S]N�U;�G��8����\LJ��x�X��ݬa>�t�H�G.СR�YN�p�����F�wu��5��[����卉g!���!�Y��'�^�dZ��^�ۆ�U������Z�t�*o:�Z����-ꁁ{��y��osP�L�e���>��R�������mZ����|�a�!ۇP��f�L�ƅ��	��#���8��vޱ��xt�w�-��b���8�K�XU�ފ��=��	SQ^:��&{�:k�2'�Fq��x�-��$���	�3���;�0k:�}�C�60�pK�gK0m����\�����f�7��#4��)O�3�Gc�W=�����yx�@�K��̴��x�;���f��̘,��A�'��p�)�v/	���ʒT�i�ۙ�}QEf�N�C��%��\:oP��
��Rʹ�V��gd�q�1��;��Z���S��YD�&Y�]���*�l��:�*e�M�%e�l�V��g�T�������#�'Y���#�ٺ�Οe�uϧM�Q̋U[�Z-LwJ�I���:�ulA[*]`ղL��s4AaiL3jR�'V�u�v�s	���+��z<=�#���{���(�k�I�<L�-^߹elCz�n�d��~�-�͵��	�#^�|�>�h�B�Ȅ��� ��%�/G��Ows�y�W���2ozzVo���2�Zp�R	z\�GW��a>=�-��}`,C��%����u�"'�0�Qn��<]�v�5#���,�������̱�t��x���q�����w'�{f�tgT:�ըx�cġ2%?W�H�U�Սw��%9`�4�~�s�����]�N� �78n�����:�Nn�j�vg�oC�<òt^��_'�q��Z�Xu�׿x	�u�U� x�@7ox�-2�\��z��a��C��B1�p�X� �;��6'ɿC���4h�I���@��D��lG
t�KwM��:嗩�[�Pװ� k��������?ؽq�?�W۴���4"z���3Yn��L�zP� �a�X���:"���x5�%�&`��~�D�'V&-���mn��x��b����zlp���F�7�Ǡ�6�7.vfh�ikmjNKͼ-�.��A��[�j-w�ԕk�ݍ2yt����?���i���@�Y��r���k>�c^��e~S�T��f�����^�9��߽�e=O$o��ʈ��v����ɛ�Z��}����Fm��f���ԷS����e�r���g�n��khC�)��e[q_������&Y�"�j�XE��
ʙv�:�l��K�/r=�,�b�U�i����N𹡁�(�?��D�ǏV��eof��x��C00(�yݮ�X~z.�	����PB|l.�zO�W��vr�Ol�y�v�Z�݃dx��9^0��/�y|6�s�X�'�W���}�ܥ:��$��r:�XJrr���C�G��G�xz�����O������]FN���p��ͮ��F�K�N�*F���=%���	�Vy�`�I?��E�Ñm�q��cG���i�g�U�5�Fn�GK�+ n���!�&!�mu&X�b�@���x�xS�_=;ݼ0��<��֨uO�u�����W[۰�P�0q��_��Z�i��J/d�2.���J��6��W 1 u`	Y�������L����ٵyIa��Ө|X�%��O?������/,@̹I�(,u)v����d�����<e�~t�����ͳ耛KЗ���''�qş�[­t�)����F�s���%���������l���)R
�_ ����BҾ(s���pȥ�$��W��\�m4V*�w5}�ߞE'�����~}��|!D������_��$��L,��D��2��m���_�k�<� �Y������&�'���oq8`���_N�"�rb8��U��X�yA���٣���1�WA״eUHG��U՟N�j�H9�����K[���$�U�����;/��,��i�^��ش���mr96,uwy�|��_��z���<x �����i�4�P�qq%�-Q8��"���Һ�����}�����0�W�����n�m�E؅�a����{���睛��T��/D�1נ	��/�Lptg.��]�."1k�W�UMSwm�"��m�����;?��ݠ	�en������n&��f±����ƀ�䒗�V���k2���<X3!���� ㉋�OR�oM^̀1�ِ����%�r�g�B%�.�L7qe���l�ݳ��h{�B�^6~f���߬4G�ߐ��W�!v��JB���1�n���<ܵf�.��>^���" �O:��c ,�f�2�Y��@��aBi�8�y.�U9R�<��e%/͘�Ӻ��؎j@!2�F�'�G(Q��y��7���S�;B-�*�Mt""K�S���B��6����� sS�y
v�	�N�),:JE>E��h��?� �
���F�����S��{������0)<ځ�Ga���HbY'��L��*L���UD7�m�������1vM$=��p-ܰ��.C�d�p$wW����J.��)�-4;z��mU��"��g�z��xhk��Iܻ=��Z:��}���,�vh�m����T��z�>�[.F�����N9ƹɺx��j�r��k�\��]4���v*�{ЇF�m`Z����#IGpʍ�1g(������W�䛷�:���8����_������U���n�lS|��������C0���Jn�0)�o�I�ކd�r	�O�����Ê�Z��=&�P�/HZ��ME�ϔ�����������	������0��,qXYt�h�ud�E6u�>l��<D�o>���!�`��F�:�n��L2G5�p7\=#Xw��C�B�7�mX��Bz�t,�e�%��C��X�&��*W=����(����#+_�����+Ø�=���gA����2����m-Cś^z�s�Vde~�4:����=��KU�>3�p� �@���a�L4�h�Gz�wsJ�\9T���ᆿV*�g�g}�b����Ab-�^��"ۘ
��3�zNT�]��muC����јy4��1�-��y���/����7{��0v>&z�"tnKH�zY�b�D�n�=p�>�NDT?V@�@�"ߚ��$�%�ލ�v��f_P�]kfh+��������z˖�&�h��K��ش�9��lhg�U�榐Q�qi�}����1�L3�隢�p�kR��=���ޖd�Ĩ�	�.�����1�dt�S���,:/p�X��U�B�"���v���)uF��i����ĝ2�q�)�N���K;�� �MWG6������|)�c�q�%-us�r�*Dt�"��eLI赔9�y<�\��d겭�D�
SNǨ��$d��t�}�nm��]ܷ_>����T^<x��~����;�ϻ�_&�o�۔_����w�Eu&!Vo���=�,	�7��D&�	OM^����OE�ս[�p-���Pw��c��;U�w,�p���b�X���kS� AqD��K����+�
�(�|főw�.��Y=�wk���������Aq^O��WI�Vt�B.�Ad��ħVR)�y�K۲ם��7�ي[YzH�����8i�z��	~�U��]�[�Çu*I��h��q[k�Nu���vvp˵��-E�0,��v^���Ű�G�9��Lpm�]�4�3a�av��Zv��2�̥����ԓLq������#;�]�E�~wX,�B;Y�d���f����$�6G���Sq-يD�Y+�h��^�Q����I�>���k�5���sފ��l�� �Y5�;�`�o�s�4L���J\,srz!\�����n���t�qƗv����@d A����W��\����8g|ֻ�&�u����븙�|��V�����S{y�������7���K�Ы��h8gAki��E�]��ᑺ 픜	�i�;3k4Ű�����*.��ܲ��]��-&]u�gp^�kCvr$IXktD��!���QE������V���^�mT���*�����t��:����T��=����)��	h��]��h���<ߝ
G���-�r=���V�ʔ�D�^��]=׾�z��������x�����<���aZ��/�z�����Q{	���>(�����\�������n�նm���gv����A1<���Oy�!�
���;(��A�_��Z�10��P�v��<�/�������	�1��>��5�� �^)�!��˱ljO��m��oh3>�v�l�:�wE�-T{��o2��c$�7�˛ozE�(8��!�W��B<�䌆��6ʆ��t�SO�m���*���կ=�]�x(p�T����.��k��	>5� ^��ʼ
5��LpL�\lv�M�m\�9�LT9����a�8�x琞�4��נ�c��i�&n���Ӽr$�A��}h^�E�5a��2�-L�D�y?�����N��� ۔��]޿6ڂ
���lyӘ�����F���ѳ�$ȶ�р7�C�&H8�s�I3�`"����v�wɐo��!T|���[wz��RL�~��f�xac2 c|a�5n��ӵY!v��o-��&��.}Yl��`ܩ��LS"�v�`�XF�GW�����6�x�������3_�&ofYˏ�ܠ^���&΁��|�x��&��Q�a]97r��F������l��S:��y^I|Gp/��oo(���;.B�n���ږ5�Nąl90Ú������kg���hݧ��gv�Z&`���D&f�iVdj��j����.���*0�(����9�m�*�V���o��h����xU[k<�:��y6�_4=Z���Tд�3W�(��n�5�W{)#���O9�v����y���G+hT帓xSͰ7��ꉋ]�}�����دD�;�F�2�!O
v,��UjڃU��6�u��Fe�tk�ڞ'eT� �Z�WW:�=X������qSר[��㙩����1�hO���έ�@���s"չd�w���jr���b}�o�`��+�X �2���ʏk��k܈G�WU;�ܧrZ��̚:�G�o8��JQ�Q��YS�y]���-Vu���9M%��K(ka��ثtK�ʈ,-7��=̳	?22��gDoQ%f�^�h���X�Θ�4��7�3���dٕ����^��"ZCiUld� ��E�%�Y�a��"�YC �_C�0���Io��]=\B�DK�͸j��nu7Cڏ��%����y�/ݾ�)Y43��I�@˯�O�G�E���5�o̉�
�0���}\���ic�[���}�̴p��0�+9������NEV�Ǒve�G9h�7�嶙��'9�IF�b�Y�z�^J&��9#�u�a�ߗ��\���dt�.������bw_�=���.0.�Y�:��$��_'�/��
z�`�O|�-g$Oh�n����)%�������6�$��fݒ2�UMDs�qވ�m�MJ�V=5t�7O1��:S�>�/�{_�*�c& ��r���`��T�=�n���iY�������%v��M{ui���XX�.��lz��oIr�>Δ/w�.*J�*q/����RpΧ���\�T���<�+F�Y�_G4Mr��H.͜UV�sс`�<�Sd��3�imS�K��mP�㙙G�}ZPoO7:n�w��s$9:����5#嘌��3'u�6r8���-z�<[R��E< ��2'�Y�o]�{ը*��Zܲ�bї'u#{t���tz��b����,P��L\5Y�+����θK�ՆwL'tE���<@]פ��)2�f�@&5V<E���Y�m]�ǋi��\��q�[�����"f	0��v�{np�j��V�T��5�-�WW��#��e]�������=Z��0⼟I����*iCi��&d���gU��re�T+]�j{���Ϊ�ΐ�"�@�G:�T�Q(Ӆ���+�t�mu��|�f�`y�db��:Ș�i�^$-:����N�������;wu�a�V9��}s�T���M�jj�km1Vء���tUP�>�><}>�ǯׯ��Y�ׯ_O�����~�_����Fƚ��61Q�G˞�]͠�����cN����������ׯ_o^�sׯ_O�����~�_������ȯ�˖�FKc`�77ᵣTSI�6�y&'F�-�ʚ��h��F�kU�[��\+j��Uys���-�9��4SKEEAE[Ƥ�N�9�h��ŋ�m��A�#�H�Vlj��MDlS��S��ӯ9���1QTQj�ūmE\�#i��&٧�W�cK�F�Z�����o9�M���j���#f�66�6�q�E5lb�G8�(�b��4M]���z�8j���ڨ�b,`���"9r�k[`�mh��^��TSyZ֩�����&(6�fY%6�?g�{*�;��Y�m�������o��-�p˶;�����_w�#J�)�ǫ�<�7�x�#^\=����|�
	����ǏNz����������^���nO��E�
��L'���]B.�U�,u)vQ���R�sV���p�5o!Å�M�9���/)�T:�@�qvJ�­t�)���{����-��Nrj>���ںu�� �DP��7����#�&��>uY��C2�I�*�s��w53&�����F�y��?��U��\E�L�hr��s.�W��3����wY=�x�4Kvξ�;p�y^���w!S�
Y���~.#7ޡ�څyx�+���2G�ph����M�e�U��{�l�!0̓ϳ!�$nu���e�^JdJ�Ƈ@�>8!�|�Z�����;G�_e���S�����rm7�00�n�C�~o
*/������vT݃�*��;ވ�hvv3��2���g,�xm@�:��_���~��;y�-f�s���U�A��1ήح�9[�mݻ�� AK|�+5�GmMP�,~����D]��q>ۡm:����{���Ch�~[۶�ױĆ��7C���p�L2�*���%�x��#�S�$����~�J7�g�:�a�������_W�5����ǔ	V*�M���5*ԯ�7Ҳa*~��vT6�#�0B�"��:�1���Cw-I���g=7���B��i��/��h&3��*tп��zL���%��>Gy�[���S���<(�x��������}����w˘~�%6Z2&�Z2)=�9S��8�-��i흡��k�V]K��՛]�C�@���S�	MDħIA�8LeR�o�v�4��>�ģ�?�wB]o�1?���r��g�1�Q��S�I�!��פ��>P��%�{]ʒT�7=s���}���樢�YE������'�\�!0�z�������]0HԢ�tS*�dI�i"��ioNލ����j��j�0T_q#А|���b�|��vw��\Q۞�c�Ϊ�Oًn����8�|e�*�C�PN%�v�}���a	�|���gg.��KhF�
;F�(�#.z����6��z���>�UiP�z q�W�v�L���G?�����5z����L����Uۋ�:.D�!���P�R��(%��P��a��z���6C�%N�����E�#1(�[�����C�yfm��M��O��}:�LsH;r�#�
��l`��3'
��Ө3.�X�^a�az�b��<���E��/���V۪Yx��ވ0$M ��㏏[��0.6����l�{m0ݞ��i?g��(�0��ݍ��a�XN�*`�f����YN��]�ͽ�4�����=�bS�PWEٱruhrS-`�3�du�0��L����.�E\�[�ml<�mo~]�j���� '<x
"y�����������������VB���J��й���D�+�2�G{���D<�q>�Se�)�3%[�{g;`�_��SAF�a�N�����F�]N������P�~Ȗx �Ѕ�4æI���oF�ݯ FfB$>s�!݋o��r���@���(.�ob��(p9��q�����N0>F'=��SJ6�t39g(�^�u�1m �T�e�c���	�7!�H`�6����T�w�-������ȹ[WW_`�.�c�9��M�z}��M�	�5Z�OE����oV�^��Z�
5i���M~v���������Ū���\��?$k�̮R�Q7}S	.�,�	���vrs�Vc�!ol���Ď�	ฺn`���L�H"NI��L��xN�l�Yu;�{ɧ�{P֬�j?��v;k���ǘ��~d�k��=!N��8O��Hb�=M����|'�9��[t�IIa�������a!���K����86̺�kL��b��:��9	 ���`���2�'�|�G4�/#OD������Q�~&�(�Û��s9��-��m_��T3P�C;!=ͧ+s.6����Z��B �u�mv���;�㜺[�aL�áN����(�	�@ۚ���9�t��G�ķS�[��V�޹�L��{:#�#�Р�dV�ea닌�����s;9A�F���}����УǏ�(���?;y��?_��}��M���eb��UvI�9!2���z;�c8���j_[�6V�U ��ښ����c�?s�B;dN���"�����RqK:y=_�ύL�j�T�z̰I��_�9O}�$Q��.̻= ?0�'�L�'E�_[d�B՘�Ë>��������ݍ��a_�$��^g�|�Y��
���S�CЏV��hZ�x�\ѸX4�����o�ݽ��@���5�%�ܵ�3�}������i�ֺ���Ӭ���ԍՂ�7Y���OP�bK��ŉ\��^#D�+��M�$�c�;���r��K#�WI3�W3�i�=�����26��Q.�
�� Ǧ�����y��[!��PG�D�d����������p���#��^�SH�C��C�
�A�0�)��eʞ��w��y�&��g.��.����ݮ�XXp ��մ�T$�c�� ^���`��2O\ɞ������ �g��[:�ůN}.�h�	Z<�Ϭ9�@|��g�V�j@���#��~ʾ�o(A�eLY������C#�m����+5FK[;�;̜�o��s������-���侩�%�'��1�Pt8���&1Ku��E�CR�[���Y)��^,wұ�b7��v�����	bvΐ��M���O9�[}�<ߞ��ߝ����� ?<Ax����P)P"UO>��{��������E�᝴(��a-��N7/T\�|g�`��РȺ��N������ә��i��������E���̓ۘ���4�I�ll�	܋hUӍ�􇶏'H8|�e������ѳ5�իn<�7 cX��P;�Jb9�bP�E'�ZPh7=s���������]�_���Z����o�� ����!��L5�ʞOd�2.��i���6�Ms�Jx���!Nv'yv���np�];�����:y�{��.k.D��L*�d�yj.s�F�2�%��41��gtk�3���Ƈ��
�|A�����o=z^K��4x�qv	TXw�u�=�Gyg~�$Re��)��z��z�`�H7�s����� ��4<����~�=0��u��]L-�S���w�S���I�^������|D�\�C���s.�W��i�~�N�t*�� �j[&z���]ڙ�Pk��ڕi�k^��Mi��0���s>2�����s40�CN'Cg���	�-=�z��ӳ^_J`I�.JL�����ȕ�-�8�t��GLSL�ȇ���E��ޙ�O+����
��Eq�r�٥Z0�otp���y��Wa4t�2�U��tjQ��ǍS�(>x7��������E%��w۪�꭬����֎�������Q[ ǲ�ʲ��-��i�-�9�+��We�S�<;}]��>�#���x���ǈP�糧�nwWg�C���C���C�{aP}s�~��dRW�[� 3�W������fm�*��U����zxl������2?~Č��Z�C1ᙏܙ�|��݂��j��+i-]g�9�+�ho c^�P�<Z�R�]����K��t-���&�3*0�b�����GS�1�Z��2��뿙�zq���C��w�e�=�C_��A�
!y{��8�:q9{gr$����J�R�|�%�ɐ�P�hR{�P<�oM4��N������Md�{��Z�m�eA�� $'�>A�m��S�X���(��$�]���z�Ξ.9�J��=)�=�Z*�޽�X�8��>�/��%�_@"{{�!'@�2.�E2IJa����
�Zv귯��m>��u�p���[�`��2�>4x�y �����]L���.#�Uz`�oj֤0�J9j���ޙ����S6��=���<*�P)ޢ6�-,�=���ˡ���(,it�~j	Ė;X['ł�pZo����~�t��BJ�u��0��ފf�^e��	)ݹ�D9���$T����FFU�d�d��]��&�hcr�6`W�[ԋ�n]���,�;쩍���k�[�p�;ܵ�F�n�F�fӁSQkO�v*em�S��,���2-�z�/)�T����_�����Q�Ǐ@��x{��zd�x\�<���q�����9�&�����4�a�Kt��7�_�X�w.�w�ʌ��nJ�s�q+ՄϚ�l~�L%�˸oW���dqt=�ӼC��Ĳ�R%�����=����)�&Fk���!�P}�u�k�j�nn�[̽�C�vN�D;6[ϲ�M���C��O��k��@�G4��f��]��{e�j�o�ѷ�3��b#��By�Գ�|�nHf�ܔ_��+$���߲'��������Oc|�j@��~?��vl�����Q!�`r\H�Sx��|d�>���`�٫B�4��Z��Tu��{9~��9�p�~����}�2%�<�h\sLg�2Or��Y�ؕ�W�������I�G��4U�B��K��ش��Ox��#�ZPP09�;�.�U��e�	�By�"�tk`̊�lO��6�5$r��w�KH��k-��0�m�=E�չٜ��M ~����<_�.���?yO>�%62jO�(�0<�n��'�g�1��U���g<Eٜ��7�[�<�""�kP}��J%�=���d���qO���+�>�3�Z�&��v�6�6�fY}��DP��U�ba�'�jw���~�-����;�
��QR��]!�Q��~��%ܭ<;����lK�5��q�9��Q�ً����r��z-TM�ܱ��%Uu�sVL�G��\��s�����~����Ǐ� <�=�U�l�W��^�7�d���ΞEFC��P '���L&
E����.{~��<Zݒ��f�
]׼בˋ��0�ȩ!���ݭ�;dvX�\���\[W�)fv���5�41��L̛�~��[wc��|�=y��5��:���))���|����ŰA��؛n��k(a�����.W�/��=�	��@ŧ�nZ^F�=4�{�?O�[u�]ꑩ[����eA8���%�J�l��B�!s��)z	Gs�eǆ��輻�<�6�q��`}S�z�g�S;E@�`��>�MƄȝuC�Ċn���l�gu$�y���¹��V�`_=�*2��������{�_��D����-"��!غ/���hZ�Xqg�X����8�l66�3j��4�l�/jٝi����I��A�A��a���'ͳ#��/�ٵ������y�/SDP��=���˭xו����'���4e�!��?coT�u%N2�=��;q�!���
&$�ŧ��.�d��l�vD��!���Qhh]U�Y6nWQ8�
݇l�f���;�y��љ�^_9�H�h��\t�88������܈MO�oB�ߩJ:f�{��V*�Zʊ�֮}�nݪ�9p0��KLU>�i��ȫ�\�k�nt�U� �"��t��;շ:�=�T��?�C�����<x�J R�M��!o&���Z��1����֟�nϠfY�;�j*B�ö����c�kI{:��Ѯ}��3X.!z�v@�"�Z�-�&\�/��*��\�ԑ��:wb.�,9rz��1B�Y_��IX�6�-V��h{�+>}�-�kit)�5-�WR�eb;z�ڼ�V3�1����_��ft�%ó��{d�]�sp�kf�ƉX*�r��|�e���	�_�Vz�k5��]Qp���hAo'0.'n������4�ǆ��XnN��)R�b���.��:�B���b�m�4-��?����;O�C��Ydl�.�Gyd�SPo΃n�
�2���d�@��wHmz�!���Scƶ|Îe���d,S�L�9�U0�q�o�w*y=�b�M3xʏ~��v���ș=ٕ��j�|�r�M��]y�6<;� �c�9y�v2'�vRaU�}M�-G.S�A������5Ǒs��[��zhd6H�Քp�7�[@���y�^K��4��/�mq]޽?��p{T�Mu͓���c)T�[��r��V������@�����z��l�vV���x���cSC#��_Yg	�d�qf�;P��\+�f����!Q���x���ӮwU�w��f�V�\JR����g_r3���F�د1�_��Ǐ�Ⱦ���������X|	�L������K�kNT�x�}������Wь?�][�f��`���3}]�q/q�t�u�PK�_�G0=Q��N������; ǆ�5���M{=��8��{i!̲B�U���UM�8�\FMi;��3��k�!��-���|��V�ܼ�I{��ޱ�:�l�ۛ��yy���2�w��a���3"N�������k�Uy�٤c>��yw�~8,�P8z�y���G��x$~��xW�p���r������M)4�����v�1h`�X��:3�P%����~�j�}������8N�ĖUOW���V~[|�>)~���O���_�;kK(�B���~Bw+ɐ���YOJ;@��jK���e��=������*���)8��f�0�su���
e�b��Wy�ەL��O7����T�;H��L��4)=�%�G�1�ޭ�S�;o2�	��5�ߘ�fV���C�e�%��D�|��4�:����LJu~]%�j��w�9���]��<�P%;y�EV�jX�y�W�F��l	�����#�y��7�è'g�����1����1<������5�1Aj�4�*"EE���W/��2��G-u>9�!�ٮIr��4�������f�kB��� ��ڰ+�L��7&�Z�v�����-<��M�"��ب7�]J��۩���7�u:�j�*�WЭZ���P�����w&�Z�F^�\sAހRQpN�H1������xr{yW�x�{z�cf�ZP��8[��0jW�'ufWCϪSw�g�G֖�ݦ�C4�l��iGJ�s�;O��K�u�.�%_!�;u��rj�ң��A�����IU�wv>Z+y�c��U���ݞR��R�ó��0�U��a�,�*���NٰS��jZБU�٨��Y�����MNK]V��c���Jn���u��{�+����*��G��G<���N�D�e�
�N]�:�:N�M���r�z��(�q&�_����	��J&Uqxۇ�h��v�7����j[2l�b��{y�
:�#U �&�Ժ�e���Yԙ���f&)F1./։=���iJn��s*���VX��-�m'�&��f=�3 ���&v��8����/u4�
��F��6��z��:�4b�&�#�)���W���K̆�ܴ��rS��j�`�Cܼ�d�Al������v86.¹���9����5R��%m#3�U�h؄.��3l#�	�y�t"�N�`�������v�.���f��6��Q��ޭ��-)ۃk�2ەu������u��m�3�}B�����s�y:��Y��3�>X�KY�vlQ��wl��a�_A��VY��(�-��PMٕZ�ٗ:�w��j{�g@Ȕ��H_KΫ6:rs��C�s�9:��Ԫ��O�tud�\��dG�^N�eu��jf��}��(gғ�A�5���a�.ΰ�90wU^��ݎ��oDg[�8���˛s��gCY��Ś�n�=a:�B	�Ƽ��T�:њ��O�f%;�'vx��:r��tKܗ��b�:�;oD���/j�wkdfM�+����B��@�p����m`���	��G�f��Mp�cUP�V5��Μ0��l��8N���ʾ̎*]9o.PL����í�{�WN�V�[�5D�r�����h��eE�2��
��2�n�	2E��W���Y�sn��PuP��x8��ڇ�!�#(��&M��ʏX!����򲆮:E#� ���y��i��+x��ukɪ�x��e���w$z��ѺK{�v�,ffԎ*��Ƕ�C4f˭`Ǒ����ۋ
�5�M����wC(��훜�u���.��˪�Z�b���
�˫�[-�ww�]�Qk�	�!v�Ęqh�Eb�l%��b�i"��U�-�M���T�o����Ǐ��ǯ^�޽z�^��O���}?_���U%��4DS�j�"��Y�V�S��R�QT�j�h�ĕ1��>=|z��ׯ��^��ׯ�����}?_���5�*��"Zm�Rh��Mk|�EMʫӦƪ��ѣѤ�F�ڵQ��ch���E��M��5MEF�ө��S�V������R̜�m[j�j�1��xF�g͍ka�F؈
Ũ��#f�+3d��F5lM
���msU�j��6q��sh�p��h�f�nִTTrK�j�"�3MF�ն�i�ţKU˷7 墇Nؤ�(������Q��0l�(ô6��3�Pb�UQ�#sb����QEM��kW*�E�AE�s:���M���Fؼ��كU��(��cTS4�k�@/��,(M3�"���UDKbE�
�'LG�O�L��Fʯ�쨯W���.��h����]��>��}J��ӥ��� ��+쪤�Iջ[.�v��"�wb��:TI��>@�L�"p��%D�Qļ�"Y��)��1
���2!D�q�!�$aRҢ��QD$6s��y�<��o1�W4A�?������8���JUJ@�O;����Ԝ/��y=�7v�7�٪&�y�e\EJ`g߸�_�b���!g�X�������a�`�I�/���Lu��6��_ql��&��1K�/\S��'�j1�\n}�?j�_>�eA��<��E��H��7p�%v�]lu#���S:hu�;�ׇzhAC0��!6��M�/�Im������u3��|L8]�*^��O̓�$.��A>y���0|��2ll�p�n\�Y�M�
f�uwkV3�]N�-���7VвT�r�5�ג���?cg�T��1���uH�g=���sW>N��zbX���M���mj�q�Γ���>� �dnz��>��3�g:��52����r���a�y�PYٛq�o&���T:�x��޿q�N�/���0"�H� Rƃ=������X���3�/ld��!v����vO��!�7!�/�k�\�I��J@v��V��ݮpʼۋݑ^�LH�dجC�{�� ��0/BNf,�	|d���Qɉ�jc�U���X;/oD.�-�pc���۴��-}�F��߃����������N�يM>idv���[��U&��Ķ���0���6���0�{�1�>��gU��
�����0�#�LV3W������Git	e���P|ؼD�뮮9� ө�<3S��#�ҲBr���͛.[Սn̨�WG!���
�}�d����N<x�(D$�Y�ȑ׻ؕtxlc0e��~��fX"3�KE]+��qz��=�6�ӏ,�,G4������_3U�^�^�T{����\�z=�mŴ�*���a�X&ԎPz�l�zǶ�h�������Uq��㽷���e:���:�!���!E��%{{6=�D&�	J��j%=���I>@���Q���t��A��8.�W£�,-�.{ )-V�y�.(�?Rn��������'���+�U��\��^i��= �����L&
E��+���]j�V��sYc��n~U�j��0%�IRkg끃�.W?����҆�>K�eyo�6=M�9q������X�É�T��LU���*,9�����������	A�
ʋm~�J�n4�`P�Cr��F�L4�G1��LZ~X�G4��<�ð*�j�Q0���y���)�U�;w�]�.1���!Ꮍ	���4*�%s��	�����3�|9�x(����ثo���wR�3��9���y C�q�&D��]R)��z����'�9<���
��"�,uuW�q�|�B|a�Z��2Z����/G�|;s.�����^�䯳!�!��P?\U�z� ~����\W>�� {�(zv8$�Mv��Xw����^��}/=��uО��S��Ԡ ��W@ޓ�lfﯝ�����o��<x�����7��`��� �ګ�rJ�r�/|u�U��H�$��Ҿ/�y"/�Y�\rF�j�Iaï2{�Ȕץ��gA�=������Ux�i��������|7M�P�Ƚ{�O���ߏ)�~\;;+���8䟦�P$@;@��_����7|������
v��Q�]fn#3����C��Pݠ��;pРLIr]���y�!=�߻�%ezl+�Ts���c��wo7�|����"`�v���wg�3/�EwI.�
��H�e�A}kN���E��E��p-U���1�uW<rC�����g�W���.Y�_��*�b�U�(3-�-2��4V�+��z�K��Ա�p`J�jU��% wL��W���cH���J`�sfiW.{��E=�`5x�X�F:�M�T9����(aุx琞�Κ�M��dj��E�W^�醐�ɝ��pe�iAehȕ�J��유��眇�|gA�z��ȼI88��� �g3���O���r�Rnf�,��{����R��}�a��m
�q�� �w*��Kc��j�>��^����O�B�L�5�T���s�*�������(G�mUa#Uw���O>�3�2ٱj�
��G�͞v�Ղ�r=��Z��6�Vl=��;�
	��A-�%�FD�칡+��>���W�}�?;���N>?��x���"��f����0f޼5ܢ0�)��H�!���[�nt��I�y�zBe�J}	7;��s(�x���N�ԝ9ۻ��$�(��#8Ƙt_�`�6��v���nT�(�1L���4,ɛf�\s����>y��א���P�mACȦ�ܪ/Ǡ�A:�e~"�vO�� -�*�W�����:Q���-(J�����#r\8�`�D@M���]gQ�B.K�S۲�s��s�[�Cw�0�]<�o��ZDW�-49ZH �=�-9��К�)�p�ɺ��u��t���]��k����$d��J	{e/�4�֮{w�p�3V�k�9*j�g/�y���U�<r�`ڀ�Pmݙ��]��Ui�k^��H�Jw��.qi���54@ׁ�5�r��٬Z�2�=a�	���V�bc]�=n�6�b�����7c�fGW'x��c�WLպ�z��,P�Ϗ�};������)�EE�63i�@;���� ��mw	�C��Y+0�����42����ٟjt��X�+�1 ���OB^��ّ�^��i�If�m��*\>��Μ=V�nI��4�P��}�����a+����W7j��=Cr�ѽ��q���n&�+b�V:�D��E����}O�I++���2Im1���k�L���,^���R}���෪����x�b��X>��	�O��8'<x�A�5T>C�9�6ɪ>����:�M~q�<(Prw_H5���"n�a$~�yo���W!FG�n6�7C�zc �x���t�=�Iu��<�X�
����^��B�N���ں
���5�q��p��1����<+/�y��P����"�E�X�ʣ&^�	-��d&V��O�Gkݹ��xe��Ws���M�<j�,�t&�q-n��Q��݊���Z��N���1�$�Z��.�tCss
&��箦m�3��IY�����p�_�F��(>��Kݟ?/w)��bX�To�H��]v�o4���ZP��X7=s�w0_XX�k�.0T�/����
@��>���=B�^)�ӛ��\�DԦ6�K9��;���TX����w��;_F?��Ѯ-���.zp^�,y��:V*0�ps���zO�K�q�0��'���XG�M�NY�l��B��e�$�n`ް������`ZF�*~$�|�[��k)����XZ�3ʒ�����G��@% �YS�{��-aɇA����%��NУ�V	�a ���~F	{��Jx��ϯ��3�~�lܰ]���2��ПT�Xec���bꜻbf�7w��jtX��04���g�L�Ө�UJz��2d1n�ܺ3�X놻s]��5�7�������6nf�q�3�3;�9wB0�u�܁.{˯iu��tұ3ߝ���v����O(q�ǀ�����f 0�J�ن�f�`��H`�,t'�v�M0��o9}6��U����z1�{t^��1rM&�1Z{M��b�C��,���^��ƃ�t^�o���2|�7$3d�J/���l�,͊���������C_���Fԩ��TI��G�E���*��%��q0�*]�\���`�w_�E����I/rD#�M;�O�P�Y K<!~/�odhN�kk=��w�kN:��Y{���̳B+�KE](r��/^��E<6������m�f8�W2VWnޚ�Z؋p��|Bc�^F�[N����zc���	���3g�ʲ����-˂ý�����xȧx8��Xt^b�� ŵy��ȯj"^�(2kO	�E�Wv4�:2�*�b���֭�sպ��E��>32	�u��" .y9=���� ��Zsl�=CVD���ǘۡ���X��UyG_�����)ZLA���5�7#�F_1���t�&`xjq�߷���t��=��Ju~JE2�$�5����ȸuC�� �ɲ�.��\�\�{e�:�,܃E�)�b�g���{E�f���f�w�wK��5�#ya4�d)hu�
�ŊV��&N+�5V�-؃s
�S|[Z�'l��x����9�o��;c�y�]h+�Rt�{rnK�Ĕe�c�>��>�<x�U�%�={?=~|������0P��X)'a�t�I��&(t	Z���c�0���cX\��53�9'v�op�|��)�9�p#�F٘i܎e.K�~AE����R:��4�߯4��l�������Q�n���:�&^���Kmn*��{���3��	Gs�V�>`]�W'u��#l�	xw�}ga# /7s�x��lL��T:�Su��kT�bm����G�g�;{i%�uϣ����"X�A�:�
汢��*����w�1C�r6H��l�Z��˘b͉,��#>�S:�9���d;�����у��T��5���͗�7|^��]'�-,��ڙ�P��l$�ؖ��b=:����-�02l�Ƹ�����٧�c���޾��<1x3��05�V�בۊ��Dė�L3%˸â,�53���L����t���ۍ�}�p�d�e�����ʃTo���Ϟe�C�@%ڊ��O#.�J�4�<�<�P�a+;���yз�x�d38��&�|Y�;�i��W-�'�r�������|W漧�؇+?[�����~U����ލ���@�F�Y/�9�ե�Xc5w�o�E9�x7���(�Z,��d����		���[bkw�ꦰt�ں��GqK�w�ͻsj7�$�j�yN,/v�);C+8V�I�MΪ�=����ޟ�ǄP��ǉBI  ���e,\(���������ٶ�zv>��k�NP��/ wN�5=�,q�6�bn���l$j���|�ȘA=Z���c=�q"-�u���<A�)�=����8���Zx����Э��Ѓv9.�F�+��8���֣Qp�Kэ�zD�TCI�������Z�I�����<���%�1)դh*�)I��l�Ǧ��䚇fG K�;����cyh{lbC�b�F���;�Re�`&J�t�Z{H���r0�]�ʵ�u�}G%ٶ�-ȯ4��Za�~��G<ۈe;}P��ʞO`��E��U�g��k.�ttV������p���tWĊf�����?2k+���ȥ0�&�H4����|�Y��K�oT�(,W)�ø�Ȉȏ8q���l� &�z���X�W�H.�O���9��0�:�n���8�,-ts)>
�X���zp��@������������{ogN��T�MҲ��Y�:��\�9/LG�|G���4�p�����k֨��%�U��7QwR~��(�ܴť���T�*�o�%����/��[a�!Q��UǧIF�7xa��q�Z���f��@�'�ʏ*�rū�n��F�q\�>+��8�=dւ5���nY/�s%��L� �|?@?�<x�x��@���H��^��N�?n��Z[��M��]FT�<�`����U,��nэ�
�G[��z���޻˓�p��R�l'�{`N�49����!��=�T���Y��8�)���3č�ϿD4�Z���na�;d�*,+�ė�LW�ο�٩�U�6T����ݾ�!V�������ޒf
D�Q�jȠ������y���#����N�_�{���044�e�A��5�� 38E�эT���2u/X��mir��݂�;v��� 3���R\IO-~˄^�o\�+����N�=���b ��'a���D��;y��c�.!I���j�HX��cC֬
o2���͋a����46)�!�K��h**�{3�Y��)�8��ۍNT����,!2�F�'�@�^=�;�����iWTz��\�?m��7�9�>���Ʉ5`��!�mN�y�,K�u�),0�Y;1�3z���w݈���3���l���ć���_*`$����^�wL��ea5��ev�e��q�˘㡫=6ȥ6���\5TBs�p��`\���7���,5��2�2Z�=w�^�H�u�>��r��T�<ߏ���8���G�U:�'�����
� �ջ��m�J�C�8O�z����O��?Y�Ѓ���9_��[��OE��k9�56�9�bvd��|���e,��X��N5�y�û�L��홪�y������ǏS@�g��â���"��F�C�Yp��C���,������f�!6����n6����]ۈ;j��H�^܆���ا�"�Le�Al�ן-t�{j�q-�d0�w�f�M3-K���g!�`�cC!!3��6&i�вT�rF��	P�z���zw�K;�B:����t�舦,:=ísBb�O��5B�WOU��ܥs�	A/Wq��fgi��-s}=Z�S��6Cr:��"��;3e����+��+@�j};w��0/n�ݭ~���^͍i[r�#��a��v+G0����ӞT"?�M�'�c�A�!ĳ�v������S�.������ZC|���_A��5�:RS�\C"T�y��./���՛�����?-�`�#�	z$@3�Ӵ��`?��P�^Ȗt;n	U��V��oR޶�4�ǅ�d!�z��z��=�fDgt����(�qX��y���X�v�g)^�[;��E~�<�
���b?�)Z��iJ��Y��6�2F�;��gh0q�F��>�6�V�0�p����|+gb��'QJ勮s݅`��
I�������m�H޾�ۄ��i9F���N��e�薫�Q;h[�O�RER�QU�x8�k:Ŗsܫ]��:�i�P�v�*NT��C�\�M$c9�D|�A#2�;���ЧM��u�:�J����>�c%.��<� �4+��n9�_oj�rr��[�.���sڍ]]�m�ଷl����b.��c!֘7/����^+Vpd��58ʖz�Z0��^���f��P�T�5�Ԇ�^�V�J����>p��J�/y��U՚���-�{wCC��~�t3�p(�4i�'r�C��:R�ݲkh�+�8I�P��Z�Z��F�nr5Z�g�������gM�C�JvIX���e� ��᪖�w:��g�gY��_�k��T�T��Z�z���m�5g{dJrv�{���-�9�a��%���圯Ow��3Qݷ���v�}���q^45J�z�jJ�C���V���}m��(�j�s�ܘ©o���!&T��N7k�8x-�8��H��y�w7\�-��I2w��f<����9Y ���9���6�{�эTȭ��	l�O��s*��2={�$$ͪ�6���gC��|t��)U[G`�)�Œz�r	U��5E�ujQ�f�.�v[�U���r���c��e�9(�`�]Ԯ�.���6��H�<�ةH3�
Z3D�x��2���;\r���p	��=��X�~g3��M=�<��T*/_ߢO���~����H����f@��G����yd�3ZD�u�^ެ�)Mq�Xj�q/y�Bn�k	\��U�r4 �hv���7],k�Ż+���vIɟ\͆�/��d�\Ϩ�u!Ò!�h��������>�bl��:�+��n��Zm���j'MIWCg^��ټ�������֙����$��(�U{��VØ�w1R��2�	��`�h):v!��P.�z�r\�]�C���kp;��ņ�#]�@��S@���1E�y�{��0��]l)�`�{������Ψ�Yۄ��f�j��ˢ�\��5l�2�������k(\��Guv6�j�I�k~S0��'qʤ�-3����n�<��)��	������,1y�h�+�6?NG7x�U��6�4wjhnޞ'k{OL�8+�(Ƿ%����,�ݵ��eE��f�񋌥��:�Ҝb�K��Tk��e��	�B�<��WНf��G��t��dzsZǦ����"�N�ҾR�2�#�{;q�|;�)��Ln0�T��Ŵ:�<�d�2�Ŋ�Pn�)����z�u�{-d4VԢЊo`ا�bw2�Rw&G]�����p㎉���!YO����s����܎Ki�Y.W�İ�_Q�	4kRm�uF �.s�����܂�m��rZs�L�#z����������z�~�}=z��ǯ_O�����~�_χ㢪֫Zq��%���lI�Uh�h��Ei�Z3ZL;jJ#g��Ϗ��ǯ^�z�z��׏^��O�����~����iX�LA�m���[i�:��Y�͊����8>y�(�����h�gm�F���"����F(�jj`��Ͷ�Q�ṌEm���TPQIMSE-�D1A\�Q���r�s�X(�F��ճF�U��si ���sjJH�֨��E$j����HD%<����;����Z��[��"�"Z��G��55F��eƊ����)���y���<M��h���i�m�Elb�g#\���D�b1h�6��lgj�Uh�խ����ѣEjJ����c:h65�F�5��lFb�-�6æ؋lN�t�&�ѭ%j�X��J�"5��b�`��kA�����ؓ��-f����|�>ء2%�|����f\.��7��н��pb�x�T��6�m�S�*krθ�g�r�g7C��v�7�G���h�y���	? G��J�~��&��k�M0y��e����[E�E�.=2[jn+ڈ�פ��6�C��l��V���!vr:�:=X��ׯ���n̂qub%��@<��
b�kf�_8��vDVK�]��V9��4�=�zi���%b�.��>�U��JV��}�~/�~B������y̓ڮV�v B�'��L�ߜħV��e@$�5��;$O�d\:��@.-��၎>�ɶ�mݼ��;�d!�e"��]���L���&(t/5:S�5��l9OU�=�A�^��U;]�&Χ`�0X0��#�;-��m�l��$�?�}�	�A��������>�0�l�x�uV��`����-�Q�0�s�ge�~��K0CqP���4HL���	0��	^U򣗽�)�k�q����G�ȯ6�!{�?����~��;çV�]��O����u�}����.:r<�s�򪑚��61P�ZC�[�4|�yTZrͯ��9�9`����C�Q)�L����O�&�;A}�����
п|W�g���N`6|?M�ʵ��?���\�]U���6 b�U!_p�ȏ��z�D{N{�ޫ����3u�;�ǟ��[ަ	�°I}L�·1i�N
?|����S���wn�>�n��m��9�͋T2������i���e�ГL�v;fήRd�3]t�m��gS@���� ������G�����a���{�����4���k�1~��x7�ε�UwIN��Y��&��u99�����^��F�^�Q.}��o�Yѧ���E4��c�Okz)��{F�^��bĹ�D��on�AwSC�Mɪ����h��w�!��M~��/^�������e���-L����x�1M.��0?U�-Yۊw2�m�>u᎛}�/�9R�_
/��"|"�b��ƛPx8~YQ�/3X����[�kn��!��m��l��_E��.02N��q����'qp۲G����d�������=>6�"�	eE�z:�H������ft�%�)�9��lvl���~��Sd��D����e��gK�)c�0�U�B�),%��[pꋇ�{k�5>�-��DM�zx���+��Ф* L"�>�#nSkS�&%��Jui
�)I�؍�`�z�Z�%@����ӻ'9մZS���<��D9��[�N�H��T��1��+�)>!�T$z����� M�vd ���]<0���F4�r��L9�[�e>�ꆟnT�}񁜛:�DFj�W���D?�;:;�^�CDt�u��P��/2N�#��3��t������e��P��[Oxn>���I�;7$�,M���7N�R�m�[rK�P��ͬ�=7����X�7`a�3�3�D��y���y��H<}���I|3��5���<x����}�o������5������3v}(e����"�_S]�|�i:^A�_�������;�B���e�^�7M�ح���3��gm�,%vO'����'I�*���nC�ˇ��و	��au�D���ƙ�j���p�?\�܃^��f� -t�'��Wz�K�c���}���A��e*7�F�:�'���8�-��X����1'\W��\�9/L���mF6�;��s[H�p�ђ�o{��c��!�G��'-P��v묺��ݩP)��k_�j�hsv,�zd�Y����������9�Ԇ��Pg݀̂
ǴBa��`L3$��#ۊ�
ė`�ki��+٣i�o�y=T��]�͋�|ke�����	����ݡ=����˰��56����ցq;���-g͏�������k�9JL����<ğ~����?lW��`�*���_0,w�B�1�fB/|�U �=>d.6�5{�.u�=b9�k��+fVU��ip��٤�%�l��Ө�X��0���J�}͘D5뜆+.��K�_��G�0��[�j�{�.ԧ�!UB��i�CE��d�%ώ�8˒JAa��mx�����y���V�z��~:B�&г�=C	\�����s���&��o��������\1�3�f��vV��}���^F����q,�zdB�����?��0������K��.G���7�29���אl�	ʖ��M��s*�hR{�Pܭ|k[��8��d�]e��ji��B��m�>6�Z�D�B�W�i�S�O�Ij&%:���ӹz��	���g������ڼ���k�]���}\�S�ߞ0����X���=} ��5�2�s:vhMYX�1vn�/���2O~Ίd��ü��)���
(k��'�	�ש~�}�+���ل���~�@�S��	�N�Z5(���T���0q�3װ�M��o"�P!��U�ݽ��R7Mǹ���;t������+�C�pN%�_<ѭ�lr���Ÿ��n�;y�1�</r����B�"���ӸM�J�/Adk)�%C��,��c!\��Vnmj��w�*��4O�
C�8u�hLKa�'hS.��a���K�}�L��;,��L��WfNnf����-�*�T6-�ϕ���: |/0�aٲ�}��l�t�qofE>�tWv���k�F:�4��	?O�:��:9xN��T\w�坵����В�3���J�*��V�hk�J%�T���/JY��N��_U�S�*v+b�;5�;%�4�[C�)h�`y��Z+Ԝ��p�f�{xTJV�Z��Uj9�K�8����̭�*�ֺ=�fc�O�܊��'J�t+��|_���s�JADG�w�w�Ο~~��B���=���ߍ���l��Fԩ��m��=���`d\62H��2r%D��ي�����+v}A��mki�^���ӱm��y��xg���.*��J7��!,���a�.z�oF��^��}B(wI`h���r�Q��3���m�"�)�%��sn_o��P�������n���˖z�-�IS50�qQLV�k���?۫�j�5s����w�?�=F`�5����N�*r=R��7C<��DJlv�h�plTz纑�y�jd�z�����z����n��(aᅻ�ϡd���M�*�M�㾕wڹ�}�	�bY'HĲ"R��Z~��яl�����A�	࿅�/fPn�=�+V�v��I��nz~��;�뒑L�R��\X0E}g��]��&+�1��򟯶��pgw�����R��.C������M�:�]1H���Û��.bp�Ѕ�n�/{r{9ϝ(, l3>��G6��ɸ^v�ʥ����F���2���	՟�j~?�;I�Q9�׀��K+h�u�"����̷V)���:-C�A�N�6����y���Vs}����a���zm{_��>��K�g������gm-{�^�¤�^uE�6�K<�ke�2��E⢑M���v$/�MU�S���3��I�о��������7��+x�U՘޶C>f�O�-�,�G6C�|�D<5���Kmn*C�W<�ې�,�vc��y���*gfmwgG+�N�)�O�1�q>.;�K;�d0u�"7"u�L	n�e����r.��\���km�2�����Ɨ�O��z����D��W��yF������\�W��g�'n�����b4-Y�,:��k-{'��FgZG>��v�;l�t(�E:U��>��7pܐyӯ�YU�xf/�fFw�d�7D����#h���nZ�{�f�ё�6��v�7',�9<(�c�����F<n�)��A�瞻���}����v����F��~ަ�wa���n\��v^�q�10�ס�9�4l��6&ɜ.�9�7�F�Z�"��L��|��Ӱ�Z���o
����  ����Ƚ�n=3�6���0.]me�����_8^&b��PjH�i��e]���=;��D���y�oL:b_�Х:&I9�R[���t�yI�i;�5�@�2�Q�g�c����C�p�h({���H5���'�ͦ�-�v�����wk�$r-t.�҄«*�n���y�>Un!s-.�9w\��%�7����I��+ؐ/;:���^�йV:k.VS�N���*a�h���R#��b�0p��#��bu��y��zں�}�yy��z���
�RX�6D
�K<�m~�a�\дU�U.��!j�.�QI#���N�����O��,{�0�Z2%B�a�� �N7K�=O(	ws;�-��Ǟ��h�?=~��?r3�c�s�M�����ט�_�F�u	8��{]f�D̬���ͬ�Y�֣3����BN(C��j9�i�a��J��0%�O��d_Tf�_��u�\����?Oh�v	�7A �cO��~��G=�vW��ꆇYN�St�d�s5g�f����s������i�7�'��6>�E��]؆E�\�Y/A�n��8�ڹ�{�+s
��\���):NX�ʡ���|�H݇ן8B� ~:��������E�v����R��WAW���~%����]<�UN������zw��=	���%�S�gs�-nL�C�	���|^�ڤ]�:�-��iA/l�����։Mt�/�v1ǥ�{�����Xyl=#���38l��ves�>�`��RT��5���d�t��A����ͪ~��;�K��O@J���и��7���d���9����+�o�&�wc�=�Ս-r9�)�{�J�p����D'Kں�$�iWL=��vp�+F)ntmr"��1^o���Fh�����7���6n�o�|�-�k�X��`�
��Uz�ݾ"tY7�s_jњ�M͐�;���5y+��7Ǻ5��\�0��&`����������y�`7e+<Y�.�'_������&O����sW��I���=<�S��ӡ��joz��Ő{n'`�ts<����E�CM�pӱ���/D��u���=����o���<ʷR��B�����p�j+�,�����׭����f4�U�k�"�m�WL\<��8��3�;vp��[zp"���p�]�c�;R)�Q���a�ի��)8��b�nM�Ϟ�\���9��C���"�z��1i��	���P�˦�D��-�	��
Oy��ebV��gfs���A1��-������1m ������{jk���D�`�]���ү���/&�!�7-����q�S�����b��.�@��x���<�ʘ	=���6���j�u3�����3���̲O`.�eI*L)�/�Xha�R���4	
�F�Z�p�4-��,,��C��;�[i�r7 ��~���"�t��y�)���o����)���?��G7x��jG0��F�p��Ђ�^���R|���JH�3��	�O�a(,k˥C�PN%�Z���2~'��rv���P���%K�K1��\�.i���!ywg[�Rެ�t��ZGa��{w��W ��V��r��w!�mͭdI���q��p�Bu1�A�U��O��>Y���l!�ae�F,"��r�2����]�v�Ξz�|��;�����O�9��H@3 �|�1����J�4{a���B�"�S��4�٦�߉Te�֫Ӭ�)έ��y�v7�Wm��{��WR��T��/�~���^��3����{)�w)\�m���Rh�D�nb�=}�+���:�� e�b�>ΟVy�4������_������[X��þ�^������5x;���zu�}%�j����f�J�G0����>kNyf�F��fѰ
l�ҏ_�ve���!�Od��Ǖ�Q������E�[�DY�@�*B!���OJ{/Jsch�-��NJǆ�=۴dv�0v�t_A"�&�����w{f=�uXS�[�,�k��-I�Q�40˱����EV�۳����x���{��qf[6U%<�g�ks����*.�?��:.@��?0·���~|�_F4�H�5Y����*��l������+���:�k>y�eVџ��I�[Xd���	�<�O�^��;�������o�#������D��g7�,�ǡoV�^�ٝ���L2b�pyRVVW���@2<k�5����¾����1{���0�U��X�n��#/6�uB�X �"�d;1n�|K4���s=�U���l�B���5��+/
��f�k&L�UY��^dVS��%B���;a�]g=�gM��;�޿/W�>����ǁ�BJB� ���y%s� ~Umt�ĲN��d})P���ơ�l��Sۼ �{��s�+Wi��r�Y-L&
ӆ�@��<�a2OnbS�JE2��&�������b�b���xm���xP��է���\^z��;��G0S�&O���O�a1C�J�%E�6su���ڻ�|Y�}�U���K��}{aA��F�?7��6Ӈ/�i�0�ő����j�,�"��f�\*�[�f�!-]� �İ�/����X��ƽ��#L��Bs�hn*�/�A�x0~9V��f�-/+���^��w=X�;���;1��`�D:n5�:�a�q���n�C��1�s��ݝ�t5�2k����G'��}�FV�H�����H|D�����Ů�b�R݋������.��n�����Xw�����3��j��HB�GCP�9}M�0�-��2")���/B]���*]�����x��	�i/��K�,�s�����1�zp;�2O,�Yڽa@���~�eHL�t��ӸhQ1%�vb�y��5[�}Fu
�:%�rq�F
ޒ��ڢ�k`�J^(�I����Τ�3�� ꝲ�J�e��p4�c7�!���˗��)~ޓr�����y]�o[U������6��"�̂eu>�"Oi�@��*���l����V���U�Y��8���:�R(u�	�1f���n)%�5��[�Z)��+�J��nr'���7F.�魦� �6�"����z؋4�k�i��c-9�m:����'7���[kR�o�.P�vX4��u�B���٪֒�Jsz�v�)�j����đhɂ����ݱ�ˋin^][\�J��ٔҎ-xզ������
T�`�IUyάq"8 8�\o�Ӆ��n����+��_�so1̺G�t�K�&)�m�f��ڠ�.��Θ��t�9[�u�Z�I�-H�#Z˒fk[�]+��$5L�JQT&h��u���h�;U-��zh�q:���M��wwu��윜����7����;��qr�V[{��Pj���{.���̷�n�3A
fU�f�9;^\N�1�׊"�tM1����a�JSN��Agh�uYb�a���)�OY+N<|���yǓ��5�W�V�O��46@�]بRI���ֲ�âɌ�l�L1��qSkLT8Q��^���c�z���{��P�����5oR�����V���"�YU�+����"�EMl��<�m��q�l��2�	J٥�i���"��#���`}&,�N�N\^�}'J��@,e���z�h��5�x.�y'}�$�����_V:9''q��5���X*ei�՗;�I�X�uY���%��g�pWo%s��Q�V����9V�³D؁7�'0f�ٝu�7.�L4l��
oe�4K�չĦ_B&�R�F�$*�x�%Nz�:W7�obL6��a{����+�{�I9n�J�b��eY�l�l�9���ù^rd���&�/ZI�^fv��l_iA�fwZKoj�Շ*ݤw�6dȝ���$PK��9�n%S���_ϝ��0}�y�{w�~�Yw���N�gM��b�e$�v���Wqt�N�ŷ�Xֳ���ɘ��-�v&��\܋3y}P��u�zM�.�ق\�J(���cV��E	%0��6��٢Wq�Gz���+�],{uܦmG+�$��]W���_K�Lo�ܝ�s���� �ʀ	��$j��'D�=t��A���=PAF�o����pcO�T�x^ κ=Z�;.6�*�T�u]]�!�����tr���*��17�
�ZV){4R�������AR���%U�r������Y/��:si����G����;0�5�.�=l2��ʝ��{ ꓸ�fd��x�+6,�uU���떒"�l�Zխ%剡�͊.1�ѣg%N�j��t�W��Ǐ�����z���ׯ^�z���}>?������~7��q���Q�lV1�X�����D[i�l�DT�16���ڱ��O��>>����^�|z��ׯ�_O�����~�_��K��!� ���61��(�*X��h�:J��F-���ACf��Ir��N��U51PET��E r9
��h�(�(���)������9���Ӊ�,r4ϫs-�M1%ht�ÑK4r���+jY�b�����,�T��\�Uk�<��b���S�q6�Sj�Y�m��Nƻb�f�"�����9����������T��MPF���\�E���l�USE̱-RTb�U[d��ڒ٢�����b���{�>mMU7����ח.D��QEiѬl
6�b-��tPU4�ͩ�kh�՝EE�m�5METUD �T71��@E�#~�u��l�!��E��4��-@�eD-��]�����-�Ù���Js�Λp��6j��z�k�Y5�:�r��N��k�7�<�-c�5�Α�u��)3��)O�Q!@p�Y_1'��E� ���Bd_�I@��[eC� �0�$&��B��\P��`��2&ى��%�L�
��H@��N� �_~�}���R������Ͽn�~��Oҷ7��۳��xl���0�8h������������h���Yg�k�6	;���;�>���
�1����V���#��##CO�����֟�)ߵ�t`�}�; ڳ��%�������ĥ=�S��X���}�V�����C�PjH�i��e]���=;��`@��;�?A���pGBYxc�T��#�Õ	����=����	�C-���=�q"�*��ݷw�lt���Y����B�"'�H����{u�����=�a2�F�+�E�1�jը�B�8�2o'VZ���l:��xL�I����#h	�N�.6�6��,KߜħV�����y[c�Ȇ��z���r�V��q��ld[B��o@��Œp�C)|n��8wJ���h�E5hm�[eg\dr�טȢ�8�B�;�A+�ȃ1��yၯߗ�M���-�2�ލ��g5��?Lgv�W�K.ڛ>Y, �2.���J��`��=^��O�������r�]�H'��� �eݣ]ۅ�P9"MnRaT;%s��I�~nK�C��(nC�ˇ�r�����h�ɐ&Y�\�nƓ_Y����kyd�it�ΆA$���{�p�6��Kk��LM6�Jf����=RG�O�o��	��/ϱ�N����Fj�7_t$f��^�b�J���%m��������W�6��%uk�_���������#l��S0,��"�ǩy.hu*��E�g�u-t�)����kml�=;�;ͯN���mQ]{�܃H<��,!c1����j�bM��zW=�(%�*�`ĉ�|^ڪ��8����}��Rܡ��]\K��� ����b9�\��H�f둗\�5{�*���Y;�3�����{䑝#�;�k��D)������^�	���&3(�oq���y�͛:��l]�a���]]��Ȱ�x�\a��0���6:3��Q/���t�֧�dz�;����)AW��U�҆[N�d[<���~Nn�4|=�ٚ�.�%C%~bL�)�Ǆ��-xZ��w���˒��N}N�cZwO���_B/@���#>m�Ʒ��WL\9:�Y� �p־�q�z�����B�#2k^�.#$mжҠ+}�o��,��W������r�J��(�0kO�fv2z��T�_��b��-�]3)����|d�	ʖ7H��d�L�4]�B׼�̖�g���ޤ���ǯ[ռ4��;G�1l�C]�Tx��m��xс)}�z�l���q��)r0��6���ӷǩ���-cwZݔ�4�ډ��c��Â�Z�IE�����银���^�<��mP��pr��z�nu�hl,][F����E��r�dtw2�j7�5<��j�"=qՊ�+������~? )s�8[�[����⸛uiI`��R+D(�u�Y����0����B`$�i�\YaǦ�F-n�>+]^���N�\�2N��	*L(?E�{������}�k��v���n[.���۩tفY�JGcz(�ahԢ�tSZhu `㖯;�ש���[i)��5EQ�5gS�
v`��5���t�U�H�`W�ڞ��	�O�iAc^�C�E�Y%M����3j���O����@��}#ZD<'P��[mITe��k(=�q�v�Kn�nw!4��4�Ӿ㇢#zXtï3G���dl��3�p٫e�Ks-��=�ѱgw���i��/�#ԣw��#�=����ap�P��VB���� ����{yN���;=!۔�T|?x��+.�����㺧���/�"�`�Ğy�Pz�����ӸN@H���̟��uCs��W��?e��J;/;�r�\�h�EϹW�H����wo�?:|3��+�u�ya�`���~�*S�N���Py���䇞�QҪ���E;[�幤4j�<�u<9��ޞ�G�Fҋ����˗ia��{�c��fMF/cyU���:o�xf�-�Tي9!��1/��s^9����?��@�F:�������}�����z�XU�3�6m�]��F��E\��{���$�V�u[�0�ɫ]��y�lgiylS͌�{
 ��{�5"��jH\3���]��7o��w��P�EЫ�M~nNk�*�{e�P9�oc�opw�̙W�b~Rͷ�.�d 6�]�i��|�f�tf��֏U๧3A����s�3c&�Z���]�^}#��=W��V�d�$eW�&A۹�n�U�|~
(�ˆO={&w�9��hAJ@��$��&�T�$���ֶ�'rDMh���yĝ��g����Z�n�!����~�[�Pb�E_��t�5�Bݡ�&����+9�1�mu�!k�ۧ1��=�ܧ���c�7��i7ճ��e��vs��T�\�e���1dGF�2"�*w[k�[�Wv�te���J+�wN�n.n�_4:��^u�"�[/k0t葃�8�E�­u�l��^��q�ue�U�>�v��؁:{�^	�Gh }�"��'�e���k7w8б�5�(Y8ɜ��
*'o�L���'o;�Ps3�d��k/�_Gӻ g�H��mҷ�welUOSOM��h�ƿ7������+������M.�lxv����$ʻ͊Dls�3z��3{;>�U�:Ux�R)n��W�#Sw����W�sT���-Nژ�<2ˋ�p#'��tr��}ZOt���Y�]�0��S��*�un���j�:D��6�H�Ix���;$��/|*;�E�#1e�u�:z�H��l3�����%�toe�=1م� �s�{k[�ـ}K��tI�enځ�/���)�F��7z�^�Z���1�v�5�q�#��x嶫���|�0DF�e�b�;7WQU,�7Ww�����#��q*����e)�n����u�-�.��#��h�ފ�xg5�'T��W���;�������*6��v����>�-�<k��w�T�ŭ���]x�dQ�5�)ӍF��+Zk':��L��EK8#Rsw�H@����,��D�c	��ܣ���*O�o-hNf�q&���j�#8�D�.���+�A4�y��v�Rjv�[C!Z#����D���t� u��R챨d��'���}�Nª�IB�ol�hT��;�l�9�,3�Uv=��K����:��J\3�ޏ?���������)�V�U}��ڧ�[����E�)[��V���ܥ���λwfF����{�-�$:�.�ke���X@�K��F��	�ʠ�8�w\��O��ʊ�� r�.���R���ϏOH1�P+&a���8=��<�;��T6s#V��������O������r�W��z�J��l\�ݬq�fV��V��`�UH�D#�N��C�r�j}ܦ«���*o[�ڬ�'��Zr��L�9C�8��,��@���m{�6r��ݴ�^W�8����'��J��6��x��5S�Q�Ɓ<�1��-�+u��OR�����=�������%͆��Ý����_P��%���j�*p\6l�I��}'�I��,	 ��z�!�>�ndt3��E��V-�_����mou䧓طoͲ#-�w��9'�KA�Q�/�̇�E���)������V�Y�be�+�Z��v(���Y��c��K��q�����W&MV��Eh����f�_k�
�fױ_z�7Ѿ�V���w5n,�g��]Z�ntغ��J�&��l�BE���9������������?�nut.Y���6��/����&�f7�a�\w���y4��P�-<���fܮ�oxM͝�|vC(������2�1"���JT�����{x�#�3Gv[}jG�h��n>�I�2ef). _My���bګ9Q�7�/#���o�`��z�_���f$FM�����B�es+y�o3H��N��sϏ�t��3{׉�%:n�Y_����\����V��j�f٭�:�u��ҷ�|�4�TI�Ğ� �)Ԏ���}7�T���:��n����g���{j}�>��I��}O�hf��lƉ���4����I�LG`��d�w�}��>{��wJԗt��Fݱ��&�n/��oM����K}R�`5(����b�;�q$�kȻ�S�<��8����{@��3�9t�G�3�������L7��!Y'%u��+I%諫� ��s�NǒDw/T���v]Jx}�Heջ�G�k��ꌾ�̿i<�|+�V���{��r&'a+�eR�99�\����H���md7kp��b����S���p�w�k��O���	�:�����{�=�"��LT��l���˨���c�.r������<����!Pn�-�6a;�{�6]����9����]~H��(A����G7��m�N�s6B�x�xvx�j�0:�-6nq��g�W�+��D���^�(vt�rϼ)�Mw&�V���h��ue�-%�3�|�q;�������jm�nyӏ�����bU�>�g;�
���I�������;���4�~P�zW�7�}6ӭ����!�ޱ�!T��GGMmˇ�����f5�p';Y�V��A�J�8ӗ��Yl�������]�nQj�Lofߩotsw�>:������֫�ͬ�{�A�
�<�y֛��5NM>�p�nM�@=vw�H3�I�����tc����1�2!���y]mC3��O'W�xG�Hm�$G9���$���*R*���iuM�7MR�<a�G�ܴ��kqVo���:˥�;yΛ�<���yhҊ�Vܡ۷�Q��^�#�ޞ�=�X�&^��=I�O6���7 �waə[�5�N�ۇi�A�0�륧�Eo]�k��]����Tҥ���76�#������|��9ks����+_9.i��9�r�;ja|���w���;dN��͗߼9<p��sT�s���&p��z�F�Y���k{rH�ԪS��n�z��
؅�#���9����jy��֪1��z{7yq�ƒVl,���T�7C[���޿D-�uw˃8{�����)�n��h㝳�v#�:�R�9�q����h�3`���U2�FF'�W���8��^Q�������	qn�'4�ۦhҀj�v�a���#S#���[Zw7z�{vC���6�e�<�z��;=&��;=O3
^�gN�����l����/�!�#^��6�Ob]E�?o�տyə�^�J�wq�K���O��m{_�H�g��0he]^�In��R�_fE���3��c{��5HH��&���מ�1 H����T���l�]�8xW8Hw"�jC�=����9�7��B��w��4�T�<LDU���ܳ��Pj�ad�[�ݽ|]����ܬ�V	0{;����ݒ���Tä�1��8$����*������v��1ŵ���vؕ�<��V�Y�S\��2��8�ܧM�f��8Dނ�I/�S�l�n�|M�udS�}����1]��L��ȿ�W�=w�Ǫ��%R�Y*ƫu=-�_�^�U��fm���]U*���5�E]��>��QGOV��Ǧ�,���N�_^�L��qbyߠ�3赲x+�J3�=$d�m�7����\�gm���9R9z�$U��]Pn}	�2�PA����d��-;;W\�q�B�7z���!�5^|��N�݀dzE�S�}���
�l�98s^}޺�;���rIXn�)ސ�[-T�ku�:�9�sP�a�g�2=�$U�������b\�G�Ը�RKK����SWR�>d�͛9�z�;{��O@�M�Q�6Ѫ��I�J��t�.�CU0h��ڸ�9��v{����7-9WA8�ʡܹP���QAV�;v^���Q|��WT�zL�b��aǤE{�VQ�\��Y>�De<���Xt�Dp1�͇{���nu�Ԫv��:�;Wݥ�-y��C˺�_7c^��+��}�;����F��[E�|ʗ-WmI�_�1�[m䡻�݂��k'K��m-4�d��S�y�k=�!�ï��[��b�}����ytQ<�̕',�w���z���&�ti4�2��&��ׇ.I�P<n�RL����Ӵ�^��&�[�)�W��&#��Z����w��� �.S���٩�J�H,\��v+&�s��rS��+6 X��W���0]}u��z��0e��ci��]��������ۺ[��NInؚ��n'���^Jx�\륮nu�͙%[bK&��Jt�O^꼕g08Q�X�M��"�J�F��Ц�2�F#ǩ�iF�W��[:��c�*o�w�٫7X�_��o�c�}oL��f�L%W_f�lἾ�!o8_1ΣJ�Q�׊=��g�O}`�b^�fӃx��`��"k:�#)��}de$���|j
XFC�v{��W(�muj��j�w���異8�<�0n�c���Ph�w-䭎�]`�Lt��!�պ�<��[Qx�4�S�Ư�0W�sX��@��k�f��\��9�#_nPp]�ܲ�־�6����sm9ڨ��{Ku����%to��h���K;9'�؈�B_��!0��RHL70ˆ�Y��eE��_Lm�U}�}�
j^[K�u
w����׶��X˲MVvl�`�4��0ùmV�7��(��t��D���.�I[W�1�3W�����ZPI�]��Fa++���@����㝦clZ���J�N����Y���׏�)4��N9����
޲w;t��Y),��_�C�j��pT��Rf��u �s)�;���N�|�*����L�Q����Ru�d�dn�ԫ�-kņ��3t�����_2I���z������
�]�9��F��k���5₸s��R��!X�|z�u���D��Vz��W��&�Nwe�ۈ��-[;,PD>&�Y��
ʋ.K�9iD�9BwP�V]��(�yًO5��oU��M��έ�#��n���%d�MN��y���T��,��!:Q7���7�]�0�a�����5�u��TT��v�n��J=l���i�=V�#lZ��vk*�9ՋhG7������ruL�����_A�UDx��G���y��e�Ǒ�5WMi_U�Aə�QR���@��]�u���S.�.�ZuA�(�441V��Sn�z5j��pv�v�0�G��YC�-���54��U�zF��|p^�t�K�Ҧ+�7&��z�O6n��f<�VY��7Q�N��e�u��>Y�����j�������s�ф)&����:v	I�s�b%�1Q����ut��)��t��Μ�?_��*��������U%#r���

���&`���Oo�>>>��o��׏^�z������}>?_�����cF*�6�Z��h��Z5~cL�E#Q4�G,�`�lm�j`��?_�||}�߯_�^��ׯ^�=}>�O�������M4�A�����s�Ƣ����"�"ZF�"*��$���4ET�T�TQ-,PU$T<�A���Q�AI�A�V�C�KW�9�*�F�6�h��!�F�n��<浛mMEV�Pբ��",gAS��奠��l�QLV�UF�
��M�1-�)咂�klQIT["
)ih���ʦ���)
*���(,Y�1MS�$��mlɬT��UգEh&)��"����
"
���lbs4PV�+l�kS4�8� ��b�s���!�����1kTTITQs�*��d�btj�td>Y��i��������[߯_=�q���X�5:H���Pn���R�b��f�&��>aͭ\��5٪�v�uWG�m�_W���~?	�sm��I���Rd���ۗ���M���į���lb��Tev���5���ڭ�û�ڹ���L�0j��5Xa�pa����O/��&����Y�sso���{�;Ci�����DɐH8K߻t��i�g���t�N5[��Uu'����eP���7F�[n��q$O��Q�/��Mظze�s�&���/|�B�dp�^��3Rk3#0��q���y3�i��á1;Rqi��O�)�چ,{�5����R�}�Lc�F���N��:vξGu���m"������T�?GJ����3�m{֕{/̫F��Ρ�GrJ��(F�U���5map�n\�{���9n�3i�ύW��!���쥂�=��T!%M�w�L�_��:�YE��+�;u�j؝�z"=O�"F�)�R@�]�gĒ|���-��RǕN�gf=��d�ٛ��ԺcE��Ժp����eGĭ��B�:�����޿����%����
�@&P��� �[��P�,�ȹ�7�"Ʉ�=�sk�`BrhU�3�C��yv��Z�+����<]K0��
:�]��TZ�������=|�ɥ�X��
�u�ݎKQ�P�������3���4Ï=ѭ�ʭ7�pa�d����S{p_A���gcu-U�z1�+8WI��q���k�<��jko�uy��~ܧ�wv�����4��	i��o�����bA;��k��>�8o7�-�ı��jt#�Tcf^7M������k�I��,鋑��do��#���ynv���xŷsk�G��Z�+��s���v�ot<�N�&��Q_�4�Z�%ڒU����ڇ���l���7>��Ò���ݹ�+��d@�+��VfM^��+�G:�ǰdǐJ�����`��nYrJD�񻬍�||������n�m1��dS��2 ]~IP��;�w\�������,c��Gn��-���VRח7���L�̈	ک�tqf�S��.l��̭��Ա���-����]tY�.��h���5j��N栽C4�Λ!��wmX�`���v
���Cz�xU_8��D��З�K�x@:sv%�hZnq*QÆ��K��s]�|���j�h�vh���O}����r��D�g<�u=�ΧHꝂ>��R�\PH"%�WF%�vS�ڳ��A~�ݾ|7x�N�����L��6Y��7#���ne�l"�vn�^���B�P2��z�דsNh~/r�u:jZ�W^����#0z�)�����O��	���BQ�u�|K�b팜8N�����V������Y{�;H�n�h�X�8n�;�qQ��ّ�?\�s jq �y��N/7��ۜ�;�%��#�g�OH�[�7}S����5줋�c��c���+3^��a�]ްG>d���.��|��PF�+e�s�l,��͔ -b7���f��Y�B(�n�v�/����9���$u�e.�Ռ��q�[~	���C��.�s'�OT�Y~;��q�#eWs��⦖�����`�F;Jq9��x���"ÄT�6�,ҡ����������]��(�K(�eU�N���[��KuL)��n�\��Z�Hf�2�e�5ЊG\�Mh����k����bAV�)���e���]��W¨|�&����7��;��;��E'U��Sst�rƼ�i��`����dC!UF�o����qE�r�f�lT�������1+ ��:z����o��/8��gM �R�#|�����ؗP/���V���no����k��Cv��Q���l�`��
���T7F�烵�TV�en�v���;���Id�WL��}#�<%Z�/����DV��m=��c���H)�=���yY�z�h�]�������,w�N��2��U��.��]|A�HO �{W>�n���T:��g�� 8[����I��o�h��w?]�uR��C��Eu�-���B5Q}}�s�w�����#$bg+�K0�"��l{�~��g=L���=={}�ݽ]��uU̞�xLA�S�7B\6�?(�8�:�m�;cGwn�+<�J�EK�j�-O�'�� RJ��KÑ�"���?*5k�ąKO9'|��	+ҥ"F��ES���G�6
�y=��;��Wo]���:��(V��)᧻��R�v^R4I���A�۾��g��3<�)%�B����%�`i������i=;���P����_��R�9�bo�E��^�ל���.�N�F;f�#�ü�}���������~���X�6�l�;�ǯ��_B���q��-�ڔ�Z�ƕ�7�a�����x��5���5�W��B�� �S��l���Wa��P-*�t�.��Y��J������o�5�{��1-^>7n�z�
�$�\��\��r�v�[&z��4cC�Ogi��}���Vww��񃑼0���y��J�`�1���=��M�ݸ���:���J{|����ptW��l�b`�f%�]��[���ڊ)q�'��c'�{6�y����S.�}�|����v#sh�nF�yf��=@�$��1����m�ퟱ�%z��.��O��O1��zM��^r��6e����H�9��x[@���Cy�ܶ�W�˒����t.����#9Z9�U�h����k�ŧܨ��^m�ñg�x���܃[���v����g�UA�C�������9��U����0��h^X���,Kp,���˨M⯛�1�ț�U����ce�������O+wl���$�)>vf[.fw��b�]p7Q�{ʳ7׮q��K�H��.�å�B[웼S���g)O���-��M�W�}�����g�#�S��A�����'W-YsNge�)�"��AZO3�s53�EU�9�w�{4�y%B��R�oFm܊�sVց�&�4�ޠ�)�Vv=m��/[-���^V4�%:�w���HgX�P�2��xٻ2gN�[D�Jq|s�RM�s	-�I�mP~�b�Ä���{۹=���AgLWn	૕����<��ia�V]!�nc��x0`7�6b�0�����>�{�66mM��4KpY���/�'~6'y�Y���Ђ�;I�t�=[��z����+��������y��~>�T�;�Ț�ϗT��7��R;}�'3LO��wt�����!�=�	t?9�*�ڭ��4�^�_�tRI6nkꋞ�d]�����zWK���;�#�i=ĕ/O�����fI�µ! �e��s�ϋ+yN�'��v����QYC�)�>��w_G#�Wq��3%��93�Y�M����:�Z�c��}>�;�D�l��2�P�46�*T�(����wuv=�:V	4�O3enU%3`Kq`�XXo6�,�-w.�ѫ��i�$�pv��:�B��>����~�;��EL+I K��f�l�X����d"�9e"��*]3�����l��Ê7O_��=o,�O�7���=������sQً6���������h63@ ��K:�~�I �t^�/������1�Ū\N�������c�*|�f�H�b����E\����#����[�h;�o�\��x���h�eO��s7 3�N����`9HVw��fof���2VR%u���By�4��4��S�]2���mJu&Q��;�UEKoT{�q�g�k�E\j!]��Px�-�.%����D��|�Yx�]�;`,P����`q&���31���3}C3���:rs�n������|4�9���\�xt.�6�i�zR��a;xC�S��i���p�֛5A��uә\@7�f����j�|ꍟ|�K���&�Q�T�����<��;��x��B��j `G{2]3}���]:���r�ջn:�4�-�]�7�w���e��ʰ,�$���fP���]77���67,3"Y;�O�ڰe9"���ַ�b��.��Y�cѩ�]o7��ؔxA�}�H:X��D��o�%�3U8�������>?���ƽ��\�o�i��4��� -�=������m���]�7�ٴ!vc`϶�흎���}ܺq��ڷ/ϔ�����b�c���P���z`�S~ٲ���M-��JV4?.�2�ɩ�d^��ެ�����8�b�/�K�S�f�{�OP/�h�E��$U���ӝy�ٻ��(u]�a\Y�;�aΥ^�sl�r��`�R��)�ܺ+3dq��S_������:���H��BG��c� ���G$��~�/�#�:�f�m�����������~/>2(��ǟ:�H�^�=��$Sl�c�'��Q��q�;n}v��2��l{�O����q�(�ط�К0j�^ǌ{뼝��4�è����Њ��eݢ@��8����&⼴���̗g��Da�7&�r�(T���C�OW�Y�u����4P�Φ�	;Y�C�i�1��[��gV���D�2(+�^��a1�4�xI��z����	Lk�aw�R��Z0f�׉mb��dhʧ�ܮ��Jٕb�ˉ�:��W�t�I�'�tm��]>1N�"�ܺ�Kt����Sf��v�^��
��{������R���$��P��ӭ�qn�7���������zߛ�~&ܧ��� �җ~��} �rg��O?r�=��/SL��
�$"�2y�-q|;�T���i��~�wݧ͋��0�y"�9&�(���0H�	+]���d�*��w;m��:�m���m�$��T�H��j�3�|�zr�2j��{5�흝3�,�����-A��͹��=(��H[1�zzK�������b��{rN�y����t;�E���>�Gf�ߖ��%a"tET��0�`�Iʓ�~���t�9���;K0�>��r��$��u�����v��s�f�)�����#(�^��g�����@`�'�ؤ^�R�kr�;�q
��;���h�i� ��J{A���n���hY��M~/o�ui�{{t�v����v�[�Oӕ�ɑ|�G���W�=^���-Z�9/,�n��#�G�FA\KXN�U��azU�+�I��}6�{wB�^%
�|<�_�a�ڟ#T�̗T����_lػfS-��a�ED��L�:���el���D�!��ś֫�	�dv:���e���G\�����~�/?���cu�җL�k�@�� e�5�d� ���Q���mԦ����#ٷ;�iy�q�k:��EZ47F�v>{����
M�\%Y���M�*�qB������>�����pGD!e�+�W���33'ǣ �8�q�t{*�⎷���8y����R������F=�G�����쩎s��W~��m����Z�#��Iu��yjni�쳡OA��_;)��D����YU�[���ܠ��:���#hʨ]rv�EM9����><���P����B��e7�W��#P�e��,�/���A�z�x�3��_n��6�;�-�ꛈ-�o�����¸�g�Mq\xwJJ��U�dJ�w��٤`��\���z���/�Y��)n	�
��1{��_��U�g[�m��|Y2���A��ܓ}��v2m���p�VLjپ�֝pgb[����ND�v�{��0�(����V�RJ��+���9@Ү����Gо�U��8����#+�o]�Ky�ˎ�ԦL�B��b�bGkC]�G�X4݊z���qy��!�c7J���(?vB��*�һ\���;�ˡZ��������~w�a5(��y|f�Ǖat���{��y�}� �J�y�3'-���L�J[��a|�6GvDG	������D�"/u7v7�v�M��/[5�'���W�n����*Jɠ��qL�=Y�di���o�PIoys��	�uК5aj�{��v7��k���&���e�uMI,�m7XU�7Q��)��u,㶴ì�*�/|�bXf�Wk�����][i
2���F��We�ԟ�|����4q���[;NmI5\:d��>�����4»�x�����o3�/:�j�`���uT�*��u���3Dv/^bt11�� �6��6�[��(�����5]�m�x�<���C�u��!pڮ�'H�_l/d�<&�hÖ�=s{(�-/�Q8^I���8�O:�WOwϞ��)��e�X�i�W��ut�>���K�bI�v�^,�g7�|�$���<Q�\��{v ��ثNb�^���V�H����D+neV��͚���V��5����q6�3���=+ j�g����'/�>�}ɚf��L�ѫ$�{�Sy/�h8����G���_�I�s��<�ߙo��v�~�n�����-�)�T��|������oއ�ټ�<��sw��~ݹ��7-V�����lw�UQ��4�˛�TR�vN\n�xt���j�\�Ev��V��"�԰�W��]�+����Ov��VO=�iM]��cv[���9��oo�z��0�N3��}4�ዪ\���ƒ9�e�1���n���":�}Oy�s�P�r^M�N\L�=�7j�EV!��H��ԗ����p�\n�k9]ג�n�:M*��5���S
�.��>[�.yϑ3n^ٹƑN[F�C��{I�u0�٢Y�J�(��B��|b��u˹v�o"Zf��+i��1�W-<�����+�6S�̪�r���#��d�pTͬ�L�X�a��\��.���I�%����^��UٗN$��y�DAyܨj]�E�n�:�Z#T]��7�+i�_����Li
���6��&�ٽ��9�!C����uh�Ș"�m,l.��I'6a�C�
�dAt��^�j*���t�JXvy\b���.
�Q۴�����1V���v6���e�>t�Mb� �4�+9Z!?��bK.J��й_9r�K��sU�u�Y},\;��e�1��s��)�S�Q[���T��A���Ɖ����7���M���,�q�C%.5x��9�/��q�w���oj7����#��<٪R��M���UF�2b�gY?��*��<ƎF����R����������~��sׯ^�|z�}>�O�_�������h1��it��)֖!(j����ikZo��������~�_�^��ׯ^�}>�O������?"�����6%P�#EDQ�ii����)�54&�5�!TV6N�.��;�bM& 4ձ�
4�\��h��0�A^K�$�3F��b+Y�����MS���3r54��rt�ұ��E4탑��DQ[6�����()&�(th&��AUDQ6���"�CT�>�PU4W�lTU^cW�Qo9�hy'9��`��<�QTh���Y5C�m��^`�c˖'QTAM\Cj���cm�"(9��"�J���NG"�<�j�*�mE,S$�z�.z���y�/nm�y��Py!y��G���#��E�Ԝ�sj���Y, �҄�hIj%"Bc�	AF$�ěđ1�D�u��Z{Κ��Tɖ�u��ڎL5n*����T賂��ue�'b6������oyVJE��R�)��$��A Rq�f8/�҄�����%Q-4FHJ)p��$�d�DDP�̉�`Kh��	@�BH�2&"�������!����t^��g��GG^d0�r*������}q��͑�,Ք�%r~�g���WG���5���7���[+5�gs#��((ąx����W���q� �^g
0,Xj�U{�wn�m�?�H�[��A�W�WGXC���&��t�ײ��ߛژ���N���zsuP��L	V e��4��l�ϱe�yOV��!��o�ㄙ�~�����'���H�/�CQ����?fLq�['ۈ��=ïg:�J"�A����9��cV-��~ M���V#-N`���%T�d��Y.qꦏ4u�gvn�]��;-y~���4+���O5E���ݝ�=ō�{������<U�<�VJ��N@���,t@$����9����=��쏤H'k����uǵ�>�C��Z��ͥ��u= 6[w/��s�;B���w2�z@��Q
�@�~��]�y}���t����U�=c�ߦvh�_β=v�:�k�C�������^�91kJ��[��NBl�W�kG�?,�N�������<��j8[��s��n2(t
�>��zG%�E}�ɹ1K�31�e`b[��oM�sew߾����R����3ˇSB������ah�I#	k�vs�ǜim&�asy�����U:ʶ@N�����ػ<ڑ�Q__���漱��38gm�#uR).�����S��t��Nj'�u49|�j́up(���+���;�n�#��D��	�-����
��!oK�M!��F��a���{�H�{֊ƭ���'ݲ�w7CY�c��n���ۼ��\.=DSL�Уgl̍���R�	wN�b�5��^��7]�q^왎wf��ú �zP�#jvMu��Uܕ&p��Mp4�+_�
e36�����������^�S�0�p��A�ł3ѷ�4���գ�I/3<�����Wz����I�~�;�x)�P��<���G�_`�t5o��ș7��a�����$X����oa�sH���WL�YeGY�M�3�5�L_�o����ɔ�i+�V)�>}��G�����B�U]�\�Ո�kI�]nEN��v1aV].{�,6�cĠ�#���W�r��T��ì���LU�_�������\VLq��iQ�V-��d]o�&Tĺ�Z������Z0�]�3����AG���]#�q��Ko��1�/P3g�u�]�-j�2���g�h�Ø�2���DH(�=��isӞ�s
c�D���/��(s�ԃ��s>˸��=B�� �B|����4��i�ge�����"���j����P*�OTY�uRW|�=�Wh�c{�ݱ�v7vz���3���i�Q.g;��!7�nR|��V�qCmLӬ�w�U�\ws��d���.w�*���駉�p��
����'��oen��������q���R�EO��M�Y���ܑs�5Κ��f�C�2���v��P���7`�9$��������j�*�1����P2�ÓGX�P��c��m:�َ�r�Ҹ�k��./�;�����FLi�OeV�����%��u�F7m�v��g���v��2��	w�u(ZԫCsPiۥK��b^+iMT3iI�ۉ��>��2@��{)�eLA�ӭu�W�d۷os�ʜp��kL�Q䝭��6<`�}'��N}C)	��7N�ΐ�N�2u#��.�맚���}�QM�,�W��z/$zM��<�GH�m��o���ޯDм�Ó���/[w�%��x�.L�n�rD�Q^T`�����z�`�o@a�����O�G i\%j��t�u�� ��t�{���X���[��n��~r7���lL%���r�d�;��a5��Xi?NV�����٠l1��J�p�]T�_*�w���4�3s�)@x6j�b�,�^&I �c�L��a�k�؜�Mf��V���:_�ʋ�#��c2��w�	��(�̏߷���br+i@�i��m����g^
6Ba�\׀�y��� d����M���/�׶No8&�R��=��P��=�_�	~�YmK�Pq{��������]w�܅+R��^R�sNg�,�PE���t<�ٽ���5������*b�=��_qH���R�n�k=W���T�m������٩����,ʮk�t�`u4�L4U;��;X����;�ު<Flb;�C�R�Ac.��En�BJ�:�uFG2
Nn���Dբ���N��*pӽ"���=��G��֗`2Q�[+P\8�K8]�a��ކ����������8�?y�ǹ�^v#`(X��[�B����)���A�Y���{�u�m�ˇ@$�#D�T!%M�]�כ&#z!�+�{v� u3��x
�ԗk��tF�{�t$��a[& ��n�'͕�{����I���y��g���:��Q�\��e����b�oaZ�r�zi�s�#���>n���7{���l[��g��.z[���B��dᐊ����ݲX��+��W�A�:�"erw�HF�[,���e�;E��@h�v�nk��Z3��/�%��;�mt�L����<��ڞ�jW�{�$��LA/��66���WRD�h��	���.�
�Dj���sz~�ݞ�x�@�8<�e�_Q�жG>,��;D�wayQ����:D�8m�h��l>��x�	���lȀ�=�[$nO��/�<���iS{�6�l�#9@���63A���³^�Js[��Splg�"�fcq�K%�����/N��u�a�_9짙�q6XϹ��+CLQ�Zi9����<��W�#�COͬ��6V���s;��寺�v��Y7q�髮��kH&x��[�r�N�^	����y:�k�1�/��X�����}��<rj�q�Ze(�Ai��(�;�9��A�
��#�ƫn#�ޫ����}����m���D�CG"�+)N�9��qc��9B��*��f��s�����ah�U�z�2=�p�\�q��$q�ie�)��a�̪j��OWm����t1��=�ty��U�1W��,2��J�g������t�^��9�s�~ۺ57뎰GN��D"q4���2$�ֻ��(!츋W����~�>��#��mݍZ�j���N_�>�Vo�\����gɢki�wY�z ���׷U$��~�����O[� �:A���0)��\�C��o]Ɲs؊�{ֹф��ƃl���'����l5$3z�g9/���_[����`��`�+_*���K.9���'�T�7G:���Y5��ɻG�.s�:C7���v�tnٌkc��<�jƱؚ
��?8��C�UĠ>b�$7`b�^���n/�N��֍Y�#ܿ�q/�澧(��yk䫕1]3m|8��$	�V����d���n]���ŷ)�Y;��z��E��<���gV��Cŏ6�Xc,,�kp�R�{wW�_dqܥ����n�Ӹko��i����;��|+��=�}a��� gӲk�tvU{�*[�(T�~�^��Ļ������y��Z��m���7�8H�lz�,گti��1�r��-�{{z����cN6{o6Ce��0}�p\׈�,l�"M[þ��{�Woq=�_eW���'��=A��N�g��ٗ5������G`ۓ�F��6�Rz:{�K`:(��c��F���sh�m��98����J>�W��)a.� ��%{�yu���?F���ɭ�͜�����F�1��]�B*�r��=�����]Sm��Oy۝��;l��V��p���U=^�=1u�#����4��1sic{=��<t���D�p�΂���1�:T���J���6��s_>&9�����������Y��Q~m`�(7x���nV��~�����O�{�`�)3�Q�.�{my��W.�k�v�Z�Z��XݧO4�:�O��81�2U �C�uI�|�d��
�U��Ր�aeuny�
��`Ù{,��J�c�m'�j�j_p���>eqQ�gP<v׿z�~�e���T��F����ϹO�? �R<䚧�nU�~�#��.��ɹi�X�������ʘ �g��7`�m��_��O�>�O[��_���z�G�6�˝8n�+iUp6��H�6(��sʏJ�5%+�R�j�L#�z��1�v1�C�d4���G��϶Ѫ��ܤ2�k<Q ��ׄ�����#8�:]O�3����Ü0]ƄP��@t���cӳE�a���=u3H
�w(�nɽ�2���;���_R�p�O���ʯ��F������ڴ��EW�__��F��sH��	��0�t�#2�dOw��8ꋮ]C��I��e���� v�n5�a�l�ni���n���}���xW��]���M&@$%�Nc�/�;]R7l���ƕ�H��,��5�����A�]V���w��F-AY��T���w��:�����y1�&ɨ���\�T��k:�s��\�l��T�!�[��$wY��s~`ڬ�5���n����&j�Fr�a-��b=�͎���]w7;U�9��Q�A���K����9���V7߽~�(��<�Qe��碊�mB�T+M�oVu��!g�Z��@�g��B� ���S���#:ҵ̥Ƿr�(��;}Z������<k�X:)�D;��ty�ǻ=��/�0OӲ�K�-��%%�~ٱ�^#�Z!u��G�W����e���/�y�!��k�p�s�v� fg=��
���zMA���M8���ز�UԠs�{";��8���yY��A<�>�T$��+�A7VVfvT�^�Ѫc4�\"w�R�Qg{o���I_�I�"j�A��9�Zz��$�o&�Nu�lG���_(�Yu�.�"2ne���㛼��xI+�t�Y�=��Ŷ� ��eպ=���6�9k����k��[� m�{f=]Y�e@��:_��0;N��s �y��)���0��d�ް����5������pQ$�]��q��D'�B�jlV����l������J�=��vg}qCwb����o|�iϢ
�����f�^%�Sm��t]D��#�+R�"���T�uʹb�)�J��;s���O�:�Z{�vs��}�C)��W����R�ʍ�U�4;�y�ށ9��v��qr�پ���JDF)��4"6��Ζ�D�וtű0e��f�ٙܒI����P+�B
��"�/+�p�[ s����R�a�����������FHk�L������_�>�5���͟��{���([7����#���X$w�0V�G�c����ZQ��E��/X�}�����S�KI4�v	7�O�2�wB�N�D5[]�nN��峈E�8�`ӻ���PJПr-��z�6m���G�Z;��s���)�s���B�;w�!��uz��Ҥ�4��'�ƜB�����}�rM���}
�X]��T%>���+W�� �i��ƻn0�6�y���c#�����κU�h\����X��#:�԰ah���ݫ����ֈ��^�kOJt� [w:��[<3�9�E`� �!TNHP��ޘ����l���^�(-7J��2��q�]�Y&KC�,�&/�P�CD�7١�\u��<���8]�N��λ�N8H#TWF���DX;٥����2�[J����wn���;�)��]0YEG��J�,sV�R�ia�y(8v��;��z�̚�
�r���R7[�[�ݨ�I;����n��]��s!N��8J�ѻ�4�#�9�����-Nu�bS߫.��O�e��r�����t������U�}ȔqJ'#7��w��ii�)��FH�o0q��wQ�o]�q_w�(w�e��mq���"��&,��P��d7wۍmd�+�A�8K}�H.�`�o���������M��z�i��"�;Y���0�ݻ�N9��p�YՑ��e�w�N��ѐ�h�v�E]s���Z.�b5vs=��8U�@GXb���n�T�l�&�����8V*R#��=W�[�n޺��du]��ң��pQoQ��3I���j$��=2��[و!]��uCy��PON󣧌ct�|wo'=Z+���Vء[-�ټ˦s���ɱboU�",�	t��̀�J5D��=�UE]^��ZZ8:o{���9����:�;"�e�0e�L�_iD��WYd�б(�m���4%wL\�*#J����D���#(����-�*��jU�+X)N-�*�yj�(��6j��iG��+nD�v�ķiz��n���33UBK�w%՘��%��hx6�d�:�ލ�w�+9�Wۉ�F=��h���~��}�uIi+ս��)�ʈ����-��S��I�]]�v�`��}3�V2���ְm�zC��|� Z��;��ĉ	O$Ӣ��\�&�F�%n�M54,�E�I4p_F)�g<���,~��t-O>N��6v�ϨCB<M�a�nR��4]^@Ht��:S��ы�7�����G_Nz�n����`5yYm�ު�D�0����Ӳ���}%�+l]��Wn�Kcm^�+�Su��Vuܶ$nR3�;.���n��&j���V��p^n�i��j�G��>��Ԕw
W��P��$9��5T����z�}4;�H��!G��[���Q����zH�'��L�L�j�vJk��� 9�q��Ż��2S*pfU����e9]F�u�ݭ�:)S�.j޻p�[؎=����u��2�IUq�2�e�'|��2��
�z{s+��뾨�j!���f��+��F�%AB�[�؇�*�kY�����i�����7�Y��JZ$E��^�a%u����l^�D겻�`.e"�G[���B�kJ���䮦y� 5�pJV���
Q�W��{�e[/d{�u��,hgS�'u��Y�:�űa��98%]����f�&�6��ʐ�F���ua�V(e���-h�j�9��
���꺹	@)i���$�i�I!��CG�Ú��"
BƼ�"���
*��kX�v���O������z�����z��ׯ_O�����z��z��ys�֓X��1UDQG.\���<b��h�&�'*
Z�s����j�&�5s������|}�ߏ�����=g�^�z���}>�O��������*����(����h��h�=��>Td6��=Z)լPjb"�(*�c�v�yÞy�V΃�y:)(�|�^m\.gF��1��BQIIy��MSG�QZqRAQ��'DLCME0�A%x��c1Ts�p�堈��sr"(�
�����i

*c��(��H �ZJ���׆&���q��DM1�ns�Y�^c�9U勜��Hj�����(��f���A�jH�y�<��Njk�K�ӧ�8��<�ÑF�(/pjJ�ռ�.A�V�E��UQM�bb4��<���<��[Fj"�^s%�q���h(6t���ع�1QEU-Q~�C%t�.׃T����nb�~���3==�M;/ut>4b�*�qb�ə�u��f5$������*^�'R�t��y�ޛѵ���n�7�o͚M7A�T�I*��^���>��ǝ b�s48��v��a���OҒ�ܸ�m� �\M�����d浳ɮ��δ��Tv,�Al�)�+<c�Z�&� �B��F׻�*l������;W�;��4���j����;j%��[�]��RP�`�9�B"vvN���Z.1�z�o6���k0M�ǍDb�3��s��K��o,u9���Io�I�������X�����6�aާ)�k=f���·tm�7�����Ոk�k�{����l卿X}�k��z8.�������퓙�Wv���ոK��UŎ����Z�h2��p8n�/Ә� N�m����m�6I��;�߯�sCa�]�=�4L�=�=��Q��	[�2V�'j�w��W;����0(��Yq�^i�љ|��H�����;W�cEM�3���3l>^L�u��2����ݾ	
n_s+K^�%Mq���4[�KI�2iD���kTzv�����pO&V��P��%��WTb��E�gLf�P�t�K����_.]*��i��z{#b�%J�/7�ߛ���Kz�^���:�g:!
0����Eg��|A8��(�ˆ��u_h����F�������0�aP*��[�A�<z.�
Bm�7�m�c7�Y�5_MP����kxb�Uq�M��s��U���D`y�MQ�&r��'�������d��zM<�����M<
�g�����E�����m������\3��~D��	$W9&=T?�Unc�}�`�UC��U�Z����|&�5�,m��	�)�A��XV�a`���f��޽������
�!d+�أo�������"���ؚgm�=13�LtV��VuԞ����
�d��!tQ�OWb����*U�d5�@������<�d��΃�Gh��K�_��l�{e��ս����ʭ����Q�jm���0�>���U�yZ�w)!U����.�|����'��%&>?>\t�Z{E�Y���8�M
�;��rv�3j�Y!�TF�Y�6ɭ��䴾���D����qL��m�CWl\[JfU9���۱A��ۜwbr�.=P��N�J�Gi��E�T�z�R�L�j�q^����W&�� w6�
�;�=���h�׻�izw�=�}O�}J��r��k���J{|z�z��o�ꕶ�2ݜ�g7kNn�Ȍ�p�{�@�<�v�k��r���p;�y�����1�0+�1�v�6�gXg�t.����ǀ��^R$� ���e�S������ӻ}�DଜQ뎡����\a�Q��F�F�e�fin��m9�����^�����Źh'���h~��� !e�+��볭a�OXwx�HX�t�t�f������yo��-H��C�J��3�w�0����Q۱�dC�T}#��e�@ȥP��j��%��e�T�2����E���Vw0�8VG�A�������
�<R�at#gj�YƎr���;w`�ns�}�H$�;��&}oS�`)#��A �#^'���^��̵7s�;��m��^f��'뽖74�\rD%�m��������v1�.��x2������Sl=ۧ:?�-���B,D�a��H'��^=��3�p��d�[Ő$�
��y�1iu�n�o6��3�r��yWN{�����g	�F��N�.;S�8�,�΄���bI��+o���Gnu8g��o7����-y�_a�Ĕ?_K)f�0��hĳ���<
�X]�H�����2���e�9s�Z4���R���u��m��f�3�O!^f��v�01���O��lwJԗr���(��Ll�Ď�zn<��s�E������a����V{p�%�x`���A��^��S0�7:}K8����c�nP-3��N�ae��Wr]IR�=�wpųH=#��޻u���l����#�=�k$k!�N��ן����ˇf�O�a��e����`g3�h�A}�>�q�[1��ѻJ�]nu�v��7�f	 ��j1��Ͼ�! ~^a�Yn����ooN|�{0��[9
 ������A�<݁z�=>���Z4?^a�}�({�<e�=i�x��B*�ǻ�󺉠R�0�E�����3,U�;�X^zNdܕ��a�PhX}bn�p���c� �������ɜLdZ$�d)/d/n��ʣ�\���'{]:�s�I�}�0�q��<���3��T;閼*[��@A�ǿ.Y];a2[SDh^;oR��\�_MJ�X��V�s�݃~�|~?E^��W-�46�!T������Uq�
;n�ڒ\�O@*H�
aYl�1��$Mܞ�������g��MU�D�^j!V]Z�L�2�ګN�؃�݇Ƕ��4�EG����*�&��j��oy�6�b9��5 L�ET!;U��pl��\'4�����nI��S|/�e��=|'����4�׉T�$����	uz^���`by����-��޷�1��ns��R�ܫ�m������Þ�|}7�N�˽�|��Y4����\@r�ɈڧYI�e�)�ir��Vs��i.x��LU��U���M5���`�=0F��r#�g�mL���=e)p��3v@�o��wMv^��sĆ}��VZ=��:��3�Ӥ��[{G-R�uծ�I���[���Ѹ�}�L���j�e�z�͂7�fkBg.�̱9;�\'`�����׍�<|�J��}٘�G�40�<P���fR�Z6����B���9�{��P䓣���\��Y�bQ�r�̆j��1�6�3m�jw3�!�:�J�l�cq�]y��N�oV7Ӈ��SH�}��y�����6��{�`�^O>���g���͐�{����":�]�}�k���V�W�s�]��5@F�������;$��7���L)X��(��x������8`�ُ���?WP���Ѱe�����l���¬�M�e��Y4�wgf�y�]��f
Pŏe摡�љ|�;�.�W9{��לt��fu9������ ��Q��#qc.�r�s���\������{�����YFu[����J�OP���E�z�a�[-J�#·�6��9��(�T
8��7o�P�]	�&'���1YhV���'q�wR-h�
�T�|}����~�u�}ғ�{2�$.�1�z��6��+;C�Д�DG�pe,��D߃J�*C�j�-b�Xk�
�K�n��s���DxH�oTq�W��@�>��(�I$�)��M����ݺ�׶��ν�҅Ke�{g�ɫ/0M��}�TȘB�B�-Ԧ$��!Y���ُnbf�F�O%j��H�د��`J����ou�Y*M��0p��$���۔����fK��ኺ6�^]��2��g9q��-�
����޿_�����BwW��ko;�f)�7����Lm�M[����Nb`�����/����Yaʩ��]X�� ۞M)�M�b���뭎��-�ώ��,:{�!���]"/ǧ�c��^[��߶���;}�Wg(�����t�.���!��`��7�օ�E=n5��.7ۚ�ns�ۙ�=lQ�V��)��={=L�1��3X�3�WN�[EMf�J�����;j�ޚ5��x���Ou+Uǧlu7)���zj�����݃�#�g`������HO1_��)&�f����(b�7�����c �>`�F���9� ��J���R�T՗u
1vF�dh��u�7E�����C8@��0��U�[�_1<�7I��ŝY�y-��P�&|u!>�Z�P5����Ϲ� b�v��L�T��h���Y�ƻ��+��E���'O){�U�O�wB�r�4ԑ�$UX��,v���YG7~�����Cs�Ƕ�M� !����9�]��g�����9
�s���`�mA�ۭ�U����F�g6�Z�S/�
w�V�T�\<8�緸n��\X�Y��]�ƭ��q��u����z�~�E.wS}՝wq�C�eTa�
ҥ!.��gۊ�N�!�<]�.���w^;���e��G+���r=�>��ѕB�*u�Hͻ�;{�W8n]ٮ��㪷��p�n]dXj5�H2z-]Fv�ge@/:���xy�Oo]y2��T�w��sL�\rD%�@��w:����ik��Y���n����x�������O���Q�Et���9��Lǫ_o���������J�imҤ,���[a��A�E�kd�l��Lh�ێ;��$BZk�}Ԯ�^<��^Gu-V�3�'���؎J9��XŎ��k���{V���j�Gp>�&��bB�0N��6^��!v��������<K ,i�C��"#�zz�_g��.H��n��y����h�޼�� T�N����z�@����z}�0.�/���q��u�tƵLr?��e�ً ��o��ڒ�86e=wn��r+�;ۼ�{��$��͐�'uQo ���Y f���������&��f��y�}�r�]!Nd�ͅ^�7O"r����t�	)o������D�W7�b�|����>ގ�=t�� 3u��;^'�����@h��Fl���k���������Q���������*)��&�?%���6�k�TO-O�u��#�̝֞"	����i��< ��c#�hEl�b��d3A��u}����*�d��o`�0?�e�]QW&��u�;����Z�Th/}�#Lnṳb5ó3l$e��D9O��-`ρ��)
�;x�Wnc`FWB8�fvA��ۦ5�n[o�3�PS	���VL�=��B��M��q�[ލ�7����w	>����[�דsNhPATP�����+
:v��f��wD������T,�T��N!�.̞�u5o��Nh�[���W\��}۝g��襨@Y�-�n�h�J�J�?_\�����|�ˆ���dE�tt��� Eȇ��'H���)\Kl�yw��2��񛽬�^�D
���C����|�I�[�WX���S(_a|S�5�@s�q�\��ks��
���{i+6�T��5Jd���X0�����UtX���mGP�;�B��w���䊉U�T����سf�u�z<�oWu�<w'����4��aن�N`e'�e�J�ǩr�2�u&G;]�zD�����ǲt���.@Ak�~�!l�:6Fڙ���a^�U�]=��z���#����4�Av�F[Dy�.�\]�_�Mu�K7H��xW���_';�;*H9�E�ig��슦�#6ހz��\�P5����؜��|W�=��������������7�k�,�\X�ʸǃ�8f�89�g$v�_eql:OQ�29��1)�v˨���W{99��Ċ ��0* ��_ӧ_���l;w�Ŷ��J�몑#k���؇����C�����(���*C��3���|�$���N�a��ʣԖd��Cތ����t[���^� =�/7�|=Es�#/r��ޞ�Mɜ6���9��޽y�������?���d���+��((�������@?���?�E��� ��>�{�E̢3�
�*� ʰʰʰʰʰ�0��C*�*� �2 C °Ȅ� C*��2+(C*��0�0�C�*�(�0 @ʰʰʰ�0��++��@ʰ�2�0� C� ʰ�2��+ C*�(� �2�2 @Ȱ°ʰ�2�2�2�2�2��
� ʰʰ�2�0�2��C
��2�����C ʰʰ��^��{��VV �!�a�a�aXe!�a�a�dBV@��@!�}l2��C
�"ʰ���2�0�*�"�
� �2�2�2,2�0���C*�*� °��ʰ�2,1�+ C �0ʰȰ�2�2,+ C ��ʰ�0,0��(�2�2�2� C(�*� °00�2��dQ,�J*�&T �@ �a ``a@d@a@a@s�r``ed	��Q@�@�& �eDd�4Ȩ��!0�� C�C( L3 �C
�C
 C s�M2�2�2��Ȥ0	C"�2!��;�W� C��0` �Q�U�p(��ʰʰ���0����8 �U�U�U� !�a�a�d�׸���A�q�_��*�B ��
�D����?��|�w���?���������%���a�fo�ߧ�3Kc}�3|�0y�}~�����TW��������U� ��c�����O��2����R��?���肪�����}�ȿ��8����O������~x�����_�� ��J ���3*(J �@�ʀ@ B * A D�$� $ !" @���  B�/�$. ! BT �  	YU�  P �`@RD � @ � $@E� !HD� !@Q�  	@VEBU�U��eZU�P(�_8hE������I�qAEF�B� �@(P�����w�/����������>��U��?��}���c��?I�?���������������C���?O?�>B����U�?�����>Q}��΄�����������/��Oǁ��!�~��������z8A�����+~��?����������TW�����G0����Q���������C�� �O���?�2UEz~G�����UQ_��A���ψ{
L�Zc��`����������|��~~�?�Њ�+�=�L���@� ���������'~���
��1����*�����=������Z�1AY&SYIԗ� Y�pP��3'� bF�|��@    >�    �:         T�@  (�  @  m��K��݋f�+)���3���wl;�k5Yl��YZLKiYn���Ml�f�U�5TUw1T�L�������U�j+-��5�O��"bZ�Z�V�Vm�Z�0����h�[��kD٣ZT-�M��K�liۗR�li4�ѵ�,�6խc�l��e��m���Ӳ�������i4��  ;�W��j���gI��-Z����:]kks����s��]v�w�y^�.Z�ݞ��k�N�ʧ���ۦ���Nꛕm�Z����vө�*�Z��[[-[�st��eRZL���֖��R�   �c�H�Yl(V�9�ڸ}O��B�
(��ٯ
B�
(H�s�p����wO��X��Wk�Y�ݷ)S���5�֭��gj���)V�[zSW���݅�qr����jw=�T�*eӻZ�Sm�����   ����ڥWg4s]t�t����n��;[��G����t�tnk�R�T�n�mж��j��'U����sy=�b�]�um���W���Vۻn��{�J�N�m�{M��e�.湦ʦf6���    a�SO]	]��;�ö��;�Z5N�#��ֻ못Ej�M��Z�j� W����W���/98�Ko^��w[�UT���;n5(�+Z���͚����|   {�4�z�:��h�z� ���{�Hm]:;Y��w{���)/2��Z7���i�U��k�M[R�f Q��m�a��m6�m����57�  =��=��־`
]���{ѕP5����6�N)շEZ����{PwQ�b�h޷���6۞�(UkU���҂��Z�d����]gv��k&԰>   �z�հT��QTv�{m�ڭ( �]p 4�v�  ,�  t� ���  :N��@ l��P(P��])]e�V�R)UQ�m�  ��� hRj�  !�pP(��  ��  ��  ��p  n��  ��0  ��  g:�Cf�mV�TLmC+m�|  ��  ��  ��  <��      ;��  ��  T`  9�\  m��  q��{���ƥ�i�͍��>   �|  7G  r��  �Ө  A�  :`  gqp  t�  
� t�U�  �S�)J�4 2��i�RU#@24Ѧ�S�25)J�  ��2JRP�S��Ry ��R$̪�� ��������1?�-G��
'����2�8�j�FT���Z�)�iaRUE	�=�<<=�~��}����6cm�lm����l�����1�����m��m�������2��J%�w@J���"+�ɲ'�FBt���� тp�n�;��bQ#l�э���R����7h�N�f�����c���9���Wo}sX&gn�#`ޝh���|z�1����/
�tM(-=�>]��V��^h�$EDL�5�!�w�G[�6�Gc�{Y��%ٍ��nj_�fu!�.Ǣ�x]�˷f={��$�\�*���\�c�Eܺ�{�^kgL˷\嬲�v	�c\��lc#nnl��x�*{�4�ww#G ��7v���RY��teԍ����v���+�tkf�ӕ�9��E�r��8�k�h�7w#xrnR��Oqo,��Xr}�<��/[l?nt�l�᷸5ą����}���&w$e�I���A�\w�;;��M���M.aI�7���Q(�G^��ogN�����b�\����9N��3-�����.�%���R3�X\���p ��˛��ٮp�x��L�˳Fn�lُ,��h3t'���*I�+�����{9�{��d�j��ͭ���7����y�q;����e�c�4����<-�__+ʳ1>�E��rC27�?XVpV�i	����d��ڀ2wY;��˪"#p(�np]�l׊����m�K8��S���oM��G]|gNH��;>〓؊���t�guO�vt�5��u���ۣ:,��ۈ��D��84j�b�(l�պż�B��Y4ыF���˽F�V6���ʣ믘� I��ދea�:k#(l�֡��/���l7�S�Nt�:�S�nC���at�n���q��n�μ:Ո�xޒ�D*'˙��fd�`+ܢ�Z��sVk�ޙ:,�jn�x}Z2��f�ǩ �t���(sy�4����y돰��[gfp���wk���Hwl��g�*4�Ο��t�S���Yע%�:R�ܽAL);W�ڵ>Z�V����;����gZ�]#����Tqs�&+�{V�����=����g#S���%F+5��:%Vf�É)�\}M�g}M��m'l���YK�;=�@�c"�,��!�4m獍�S�0�tc���^�n�\��7u8��e
8N	�S��F�q]j��tق	w ;ocXq���V����;O>�Ot'VL��a��(2�oq�'P�ˣ�������s���t^L�zm��Lz���8wU�p�o�F�|q�hQۊ��Xa�D�;�v�;!���;��B|7[1Z��.�v��Mnɷ9���'6:�}��kpٵ��4y�%��v�8kq\�e�~E#����M���Ei�o���!a��R�u}�3V�B�{{Kj�˴`7t����x��@D�հ��2ġ�+�[{4������-���#B��)��ڙ=�c��b��n��;��-�7�22e�1>��f���&��877ND��LJK�W��|����s�'m��q㗔MLӹ^��r�Z�ł���7p���p<s �ŭe��C���ɸ�=+��q��@������ȫ����=�qh�'� WɕmuR|i��VqB�(gf�Z���5]�J/cL[0k��]{��lgn�!r���C��ou���ЃAz�]��CP����4γ�(%��$��r����ro-,Gw��y�m�d��Hܕ��BѹN9����� �ƻgi\7�5W�w#�f�M��@��r�dx��	3k���q�t���`H�>ѹڞY�	�di�CgA� _���6�Y*S�JV�*lw.���r�.r�.�9�-�w"�۷�0]�t����ܲv�Kzh���N�oqէ.�b��>�hsx�WLÜ@�������Ʃ���5�.b�3��۸����5&�}��qNX��	c�M;b�al0���DbɅ�����j�mMgN黀^{+��C���a��n��㳺u�E�r�P�l�&�ۅl�ܰ+k��� �`3O2Vk�x���:�r�gL٧�;�|q��=&�k���1W�,`9A�� wn��Θ.�OA��Tg �$��}����owS������=�]j�U�a�a+��	�'MȎ��=^uk\�h�K������5�������sZ/c[��
\���u�0
�坵v�TT�����4�ǎg
��6!����;���ǚeRV�xs��h=��[��4��$�Պ�mX���n��z�
�(��=�۠��hQ����N6esA��pvran������хQ�1��%Z��6>g%��i���:�P�pw7�A���w�kp�B��F ��7w v����YX:v��������-����c��&#��3��D����#���;�1�`�	˄�Vl���iñRa}��ٹ���,�vG����<`-�V�3iطvt��V>�����Ψ͘�6��\�b�s�.��FƲ����v��c�C��}� V��޽=w�X�Z^�y�ў4V0�;8FQD!35�[�ĝ�rh�,p�N��4f�&LVq��^8{^��i��
����Of��r⚞��{tR���{/�<��sė���Ǳu���t�9�qǍN�^��&�d^�i;�V���7f�퓻-�ԩֳ�U��o������6�\�dՂ��3�Wl�����ɭF���a�i2@$C��mkWhӧ�5�ܪ͠5�`[`���O52�yUn�5t�F!D��I��3z�V�I����Ӯd����+���:�c��{%�{�s�3N�Wv�
j
ju����k�ZC|ɧX���&W����8�(���#;e�z�tW�����	����r��H�;����`X3����:�WIx	��@�gS������Qe�����0�i*�I����.ش���c�p('c�S�s��m犹��-�+zIqۭߞ�$�^l��z�7r�1)iאlB-u8xnG���Y���n	!��eH�1&�\-֣ҭ�S� (.<n�*�*�yRҀ��v��6�ԑ^s�Fۜ����_v�yl�F��Ȝ�W��F�V
��-�B:�o�� F�hP����C:��#�e�r���FЛ���İι���S�J�;~��gzN�k���T��S�ޗ�WӞ�\D��`�>4�z��+�$���R��
�q���M� S�0��N����9 gs���8��rhV�jdq`�������ږ��vM����͑���thl�q��P�����d�jK7.���Z�#�-yҌ��3��Z�%��ؘ�0�G�Tx'��φ'͈!.*������y&rc�ۀ٢����.�)b�YM
�כ�uL���cD%`�1*ʼ1�����[�����8�T�ot�Fq�"7k��n���F3�9����r�2R���^�=���}��*��K
w9��=p8��=sJ�CE��\z��[�˛�t��G{~P��gc�@s	�i���
c..�D�8c;��"�|+U��:�	�)�58�8U�]�>2J%��sSR��9?�t��G�6�۴���,f�	vMԬYxL%�[�%���J����m�>n�)��p����FWvr9qi�� R0�%�ܦ��S:��\��pcAOM���֕%��&�%���3�T7��d;F��&�niOBA��x��nk�N�̜]Ę����r��h�,��u�7sx�ŎE��� �Y��X��|5U��]<��|E�j���L.���ؚ���^��2��7�p/rvS�zf��Z;�)`~yF傳�<;#/�����Ǹ��~Gg[b��}N]oG�`����$o�wg�Ls��6�t�-'��݂�a�˅�s���F�Z�Z@��ln8��GU{5I�b���g*�m��<�@Ê=Z���Zf����\<uژ/_�$�O�o<��j' �"@��D���v	z���H�9���|(qK�v��ԮT�Ls�|�zk�r/���@#�(�g)�6���һyw��6t��jEه4\��q����
a�7�cr�N|	S,�V�JΚ�����Q��;{&Xq.�|�W6#��n�kA�t�wu_��&���6<�ݑ���!�8����n=�H8$#~e��{^O��,HEEq6L2��&Q�;����U�t�]z��<n��:7��o2{�1<�a��%ڷYWy)��"&�s�5�r�����sg[�6�����5�+��ͱ!�]�1,є�zFr0���/
����w:�-�NfL{ڱ�Î�)7�����K�-=����c=�q��T�9x���=�3w��D�@�q>�#97�%���k���ů���up�{x����P�1��EY��T+��)@�أS�����7&C�Y3��:p�k�����9��M]+�/cvAԞ:퉡T��^ƚv,+��+���`$�V��΍��ǫ������f��6TGN>`�] �#4kָ�Ϫ�P�ؚʡ������B:NdHA^�ݳ��"k���`�\D�:��YN�zr��7��.�K偖6̠�19Ӵ5,�fō=�״c�:7�l1e|�������9&շzj��=瓛;͗�.�k���{No�ݙ����'YX���`�m�۵W��(�-��U�Z���s)x����Iۯ_MA��ͦ�q|�ѳ���z�l����5��[;�2%��]z�F�خ�}ϰ�(�m8�çf��0��»9�i�}D^%f��:J������;��)��hr��.�<���8sA/;	�;o�j�Bv\:-��E���4t�����{v�ء��.��+i6����$�sBf����q�g�LǙC�פ�SA�4TZ���Op1Vr�h��ª�Mv"{�^�n��@秒nymʦ��C/l�#�q�۞��`�~{�������ݨ����I�U݊5q��Ԅ���j���Ǜ�f� �y��44��,�j�'V;-N�\۹��juޙ
���@�"#4먝�"D���i>$Z2j�#y����oUM�&A�ݻҧ[�d��WH���b�c�'kS0��C[ڹ��|x�=k	��_�p�t"a�K�� ���&&К�7%��^��b�W`�m�P�W&��y��sp��r`��Й�la��jV��m�1���νDxN]� �t%�Bu%a�S-��J�-�x=�i3%�ѩ2{��<��״6-�N�Иi��b��JƝ1ˏ���o�m;��_\����u�Ô]���2~[����K��L=�9��M�{�Xۗ��#��m⌜�[L|�e�]�s��6=G��pY��v�:,�4�ǲ���3tμ��BVp�V�a��S��D��S����o ��`:��s������~��y�Ms8�u��0���oK��$��sjL2�[�n��>�i��-ˠ-ܳx��*��aX�o`�m�khv���m 2��=�<�<�b�a|���t�~��l��d�V^�7���T͈���#�hO�����	�Bt��@�!5�xŚ����׍�D�-�X{�<~���gU�#$�P�$��90�p�Hw����R4�4�*YCw�I�搒�殣���T|�]�fؠ��6����Huڭށ�D��ш!ʎu4�w9�^���b�.�y�t>�M8M���Ы�_l:���zg7��1�T���E�ڻ;�f��*�ogC��.\H]8��!�m�k�� ��Xط;o�-Z�6��t.5��}�7K�M��Mhm�h�<����Z�)4N�y�ֱ��jXr�m�9n��,,���.���d"��f��r��A>�@w]Kt�B���t�xib���K}��}���ck�\�	N��/x���f��0y��7#�)�oL����t����]��/o`rdE�Ÿb�ݖ�\ݝ�v����q�V�Ƌ�Q��"��E��c�E�/r�Y�@%;�\޻��=�.�7��&��\8�i��e�n��z�á�c�ɑbZ�D�fZ5f��������&���M��<g��U��;�^��<�ޛά�bb�]��[���0\{�5Wy���-�:�n�ܗ{�Z�ͫFN��R͞o\��7ɩ&�{sK�`�8���{pM�D�`�5wC��x��'[X'���Bծp�M�{ǳ����ۿ ����V�$�WdLk� �X��-oKf��w�㜖��.���A��ip\V�mgWN5������B�a4�������l'���E�ݦ���Z�(A��U��]#�y�͙-
�+v�v��쪮�w�gkP�Cl	�Y��:r&�����TB{��2�.+��t�f�Y��83!$�V�[���9�G�K8�q�]���k�f�p,�W5�hu�pB�aYP��pi�\�{8��ۉ���t�wi�i�V���F�;�p��I��A��[A��3M��/ `P;@�5�&�`w-�ԈG��ւ�u�v�n*�qH�h�g�v�{���q�!��7E�]lxX�`��sz{�CXʥ��H�hnp�+�(>Gw#�\|;�f�7��6"�tֵ�l��H.��(�f#Ge�ٓӝpj�K��PM��^ ]!�t�
Tn�dol���<y�`����Ӊ�n<yr��`f�S ��M�0_nD��\�x͑\	c)b��+�9��9�O*H�m��1&�j���]�{�Q��Nm��G+��� ��Ν'����rܐ�cwp�vV:�B�J�]���Y�]��ȱK,�WWM���z�C��*���d��7�8�C���[���ڛ'}�����5T�n u)�%jX�_�y�{S�f�{��3�aZ�Y���ޘ7�%��Q�"�؎������g�Fâɗ��Z��/!�۔���އ����9i;�U���o��.����m�>���W�;-=��d�Q[�)������qJ7}��)�T`Z*N��/���l'6'����;�rN��R/g�MyXI�2;"�ؓTN❖3m'Q@"�+3R]�땁���֚�A��7�[�װz�^0�u[*�H���:�7�y��4���MB�x`��jӻ����coR����o��۟#o0I����,��I���8N�::���d6�=��80^�9�,x�rulJ�&�L�����'�V��7Kح�$��֓Hq��t�*�.��/t�f���p�vhG2�xD9�1��[)n�͙q��b[��Gq�G�g���ľo5��"���*��n=�6���4ث3]ݧ��Xfʜ#;���y��V��To�w���/kn��Q����.�ɱcj�I�]��M��L:Ӂ�N�4q���o#%��c�7w/��=��K+7s�/_.+%)Q��|�
���/��βR�}�&E�c��+h�+Ɨc��KB��iqv�fLe��;�՘�u��P�3]��9d�C����仛�9�gP�$
7Y��"Vfٻ՛��2ƷN�S���s��ʃ�@�Ž2���w<{V��C��[�6�g+�^���h|=�5*sӁw���vnzL8qb��৔�݊�4'�v��y���8D��MM�}�̇}�9e|��
��j�0uB_U�'�h��S�4����|�y,���9E�X({�A��R�q��Z�bD{�G��QW�Ӳ��,�z�Sj�B�(2ve�夈᬴ruok���7�6Ukd�篡�E��I-
W�$tk�f�Wn�EBP|�Nec��z�v7V����S���sL8f+��Nw-����=M�T�̮���%%=Bu\��w�.V�o��'��6-�ω�VOC�M�zON�oZ��Y����NU���XK.5���{-e�ܱС�f��n��`g��f�|( ��A�ڥn��"s�{7\o�V:�r��p4*��PT�e���ܝ�Jj�I��L�	e�9��Hn��<��	_��{@�e��P�K,#9k{�+���̲Kϡ��
���9��RoL��4z&�|#�E�U㢮��u��ۼ�nr�QI9��w�A4��\N�`���"�k��P� ��V��R�u0f��IB�`ѯ]Y��|�օΚ��k9c���
Pe"�����t٨�$ͻ9�k~Ps��KQ� �ùG[a��:n�'~�{yP�F�AdY���.A$]g-,nC���J���b��^Cc��U�:�[J[��|'>��B�����(R�L4&����Dj�e'e���w���9�˭�۸%
�2��k���#� ;zoaZ�v;�8cE�j`U�>�s�y`k4�C��'G��7���W��׆�#
Lwh�CV=���:���q������a��ńZ�(v���<<'].��*:P'1���0Y����٦w7����*PHEz�Ks*���g`V;��I�SD��VA�hKGC4��aПO�'ⶫ@rU��7����'n����/�pN���J��Ti�pS�r��P��VEmVJ�va��x6�)Sx`��¨�k����̜ ���kYC���)�Ì��Xc��w`�%�n+�qՖU:� �P�)Y����8n�Y�:6���6C^�	��CT�.n{O�X���K�.���g]�����)�SW�T���S��Ll�r�b��B(ƹ	��i�AA]kJ�j-����".��Z��͗���r_r��Y��$�8��U�3�pi޷��K��f�
�\�e���2�Mn�lF(�i�k�j�5���u��/|�=�: ���=��7<t������&��Y{��ǻg�wPl�R'�Ot W4��j�Uη���}��y�E�Eg�}/fzl �\i����%-��U�ݔ��t��Fٳ%*h쭀R��Mx��!����}�Zc��e?���OUۏ����� �ޫ��ˠl0Ԓ�c�/u��`�q֍��1�"��Y@�g�`���pwg=sjk�2�-��gE嬩�Q�뻣\�7"Q`}qk�S�
e��K.-,�'7]����k0ł�G{�V��������Xb�N�%�S��T�.��'2���l�X�����.V�珝_<H"�?+�$���~y�w�����qc �����X= "jO.���:z�yÐ�5�LXlW\֞Be�ִ2@r�E2�m��.�f�Ϋ���b��m��kq�ͤIK�>3ȱ������k�hw��N���,I�Ÿ��ݩD�R�˥TR��p��\jvӺQs�i��2�nb��Yx젏1�(}iY�/^ih��jӓ ,�,��
��r�!�&��xt uc��䪲���X�n��<=�иVu-sE�Q3�+o
7*��F���.=��e���fܿ��˨����	��ja;�2�������^�˱T宂�Ȑ	��e=��JYY"��<(�x���Z֌���n�L�KX��sve���7V�[�s�kS�b]���M�݂�x������l��P[�)��T+]ږE>��@嗑h� 8�����p{W� M\y�</��E*���2��[6-ϗR�r�}۔���F�_es$�[�4��9	��l��0���%nc�c&qTӱ�y|z)�s��3��-葠��,�:�yw�N�D���B��A���N�S]��1���8�����_[����2��<�sM>S]������779c��>�~~C�I\B�F���w��Z�K(s�b�c�f��������n�'7��B�������s�V��������nv��|��k%�'9��)������D�����ܷN��vuGXWA�G< ��]��xV̐�Y���oh� (�M���]��Ϻ�҂��2������"�!�q�bdΖ�p�"#�R���$��<�Φ蛡�T-%qZ\=�dP�*x���k<�'�	�74��0p�fӨt����[Y*�,���q�V�=�B�������8�n,�g̵]��g��f�2w�9�eu���O�v�ޤ����[��=��R!���N�[��K���D��Pk���VX�۹���u<"�f�����)�T�&���"�E�IB�F���v��SF.7�ߚ"�x�o_eI��fV�x�X�;��D�"#hS��Ѕ5��{��Ԛ�Æ��,I���t�÷/��}��6���h'z�O>=ؙ7,��������6�u�g���*�7hɲ�i@n�G�j��MG��S���}��_b���-�nGJ!W�|ǻ�N�U����9�����I&�$�Vu��n����%o�{��>����}x���k���b�#�e^tU'� ���=��X.���e�r'+�[N��s�Jg�N$��v8!Α���7�[��ѷ�MBh`�CW���eޙ�H���{4f�X�n=��g�zH�a��\U��l���d��r��I�{�k�X-��noT��j���y���c�HH��i�'�yn�)����a��M�=ll>�T��U�!PV���Y1>6�
l�nn��	i�b���X�)�Tͼ�g^�/�_z���ni��,x��@y2%�wϣ~19��=[Ǥ�k:�5�aX׳vepB7�[L�����l�r�4lٰ�Õyc���q�)zrGxt� �,ay'��ָ�A�}��p�M(�t��5\5gGl�3HGgD�P"Bs �f�ۆ_I�PŊ��ei;Cl��xq�(Zc��U�����3	�֝�zfgk�q��YfP�FPY��V�K!�{ B^��9��X�����	�B�V(z�q��8��V�����L�3qc�jmm�z2�s{�R!��7�q�ޫζU�����Ѫ���2��N��RE�\/	JP���m؅S�J��n��LXd�̗��:�B��[�~d ��gL�<�����'�X��x�>6{�(v�yrg5u�y��ҟA\�b�w���"�(Ew-�������=J�w�0RR��ן���ZJ�����{<����T㻛 ���^w"7�5��́$�EX1wu��jw����/I b���P�c�ߣ�^���X�뢖�C�=��-v3��]�3E�8�Ϻ�b�V�:��tw�c�$��%=��T�ٝ)���Kz��Z��ԅ��ޡx��q"�p�K]��}Y�ɷ��VI�N*�R��Da�s�:����*o���l����wj�j<!�l�ޅ���V���ۭJ�� %��"�tt���]���F��{�|nњc�Q˙�>�y��	%'�P`�R�P�ŷ)��f�[��c8�`�}��l�^����wx�K�c���껚���U�+v7 ,��4�8T"¸��\�V���R`��άÛm��C"l�Wu��[�s���.͛��L��E�Mr�R}>�P[����^e�s��XּkY7��z�jfMڛ�D�`6J-6ն*�Y~=:��Ź)5������n;.c��Q���p�p��ea��ˠ֛�̀����Sd����vW9T��8�ʞ@��ܫz����<��h��]a	��x�P7�H�gN�H�
 Z}�:�y7T�S�X5�1�7�7n�β��5�nu-�hec�"��������qus޲����7���j#:@3Qy{r<����M[�|-�7�R�rqV���Z����l;0n�ͭ�>�Re�,K��6ګ \���үx�^�<�n�"ke�|�hի��=1��H2���7�V�=�0y�����p鼝 -�m�G,K�J�ŏC}$Nn���+��(�+��QL�� �t����sp<�n�K��7�wz#1s��#c�������0�`���}jh7c�TӁIxK�[���e2>{Nq�6�>�5��bo����0G���.�"o_�7ןN����K�
K����r^�[&�=����(�З��-��ٯ�[���j�4͖OI�X�5Q�ۢ��?��t�Ö��-K��X�@0z{Su��\�������񇴰����ʀK$D�����T\�{P�D�a��R�l�G$��47�Ej����}��t�ƴ5:L����W�kqV�Wh����˳)��)� 
up�T�e&�L��ދ�}򝖢�b�G"�w��k^�!t&t���ʾ���oj��y�Y�C/����1kν���`��Z����*ek�5'����;���x�T
����h��Le	͵wk��e�eMk���OA�6Qs;q1���.����7�o!{���m�ǘ h�_]be)����"ژ:�c|[���{���5���,>�:�h,�R�Q��{��:��3ݧ���7A�e��K͏�z��u�U�x���mĉ������Ysh	�e�X����Q�s�yw�en�ވ�z�n#���"կ�XpZ�%�M7Y���OWh돧�"2Ud/|�Q�~X�����{F�68���C+//n��i����zQ��l����D�v%�,�eI٨�|r�w��Ez��LOu��	w�V��Ic���o�D㼪���,q+EKp佧S[{-�/���cwf�U*V[��odR�FC�\�������+,T�[���c'NK�I�[{���)p��g�d��O���2܋��@\&@���ſ�ݸ�mU��r�Ө��V�R.�M%��2^77N)*���U�`86-�ZE�w|V����˷Q]��R�����N�yy����н��kc�1��x&��5i%׳:v�W{��t��k��*�[�E�F��}yy���F��AL�}2�����oo��$�͸M;4��˩V���V�cw�48��|^%�����^�K8�9S�ڻ=�>ۤF򆯦J7w[R�Qu��gW"��b8[���d��T�y`ټ�q��
���9;�v�z�:���DR�۰[��]n�oy4�n�J&�Z��ʳ�wC�����̑Y�y�_>�[��Z�D�o����2��QY�U�(�f��u[op7*�1�� ��un�%����7VZ��]k���.\v�Y���;�ՙ,E3(�h�,��pt6�00�ܾB��c����^=�q�pN�ǉ�7�k�=%�[�L1bWQ䇂X���+]�cko��$~]l��Ԟ��tTs�%�H�z*�P�����0�[G�j�&jk\�U��8eր;����� vZj�h�|��I� �LjO5�{}W1�2uVq�p�v���b�MV��v�Asr-�0��羽����wW�����څ��2NK\_)�j�n�kf1u#܏��=�89`������nܫ�Ϯ�á���,��۩E���&�f�����E[��ܕ�?�ώ:yVOS��1��3�V"b�f�Yr��묇vݺ�gw,1[�}n�;�����d�&mӭ��Sٰnt���,r���{�i���O�fu��۫�R�펦��(HB*IA�QȻ�r��c=�A��ʽ�{ۣ�r�a9G�.���/N��[bm�)6.��N�t��6lSa��r�āJ�'�v��'gE����96�Iw"�*T���F6%�fWt�.�~Ji����n1&�Mc*�I���3_`������[��Nl|��꯾������0��`�6���O��������Z+�{��3�&c��:�sm��ޘ$�Q
�-��t�Ҥ���U��J�k�+���]6rV�X7��&�4�Zq��S=��G\GВ5�=�<.��\��giÝ��B��t�h0�4�q�4���:c�ރٷii1��b�`�t[�Fҫ\�k�t"\���l��j�'8���������a4N�Y�ۭc01[)�}4]j�K�3��,��|�Kn`;bN�˜����1v�m��^�)ns^}�ŧ8Z�)wy��u��(կv���xɁwN�#���V3)��¸�;nxcB�-��}VHބ�Ws�5�m,���Z�`��ж��9A�Qp{(Ӈu:Y�!��V�Mq���X�ED��8Ns�<x��j���i�������(��
��{���lC�+ډ]8�_l�Z�@2U�����*�U�9S�Y��j���q�䮃cQ��Һ���O5.�.Q�����7��:il�idm {,ld�2�t�	��	hdV�;Z=�$��a;�� +��F�mS��=�;VV�����"�j+�-��۞8tcp������������@�2���x�U9b@�I��i��K�Y�xj����=�(�ś��֞�V2S�o�}�79��W8�#�V���&|�كD5�凷f�H��b2֞v�w�S��w����D3���/E�q�z���7�]����Xܭ�K���oF��8#��2=�.i���=�.,}���xnol�71���#�O�k���R�~���ժ�X��t�� ��E��dQ�:�V����Q�*����ӥ兮�Ok��x#-�Rtw�D���C7z<
Ź��$_ϔp�u���1=}G)sBճ�����c��x{��� �x�/��1�Ds�/O��������[��u��b�hQ�����+\�j7F�u�$-�N�ԧd�ŏ����g��5X�	ެ�B_Fz���Η��z�7@-�>�R�5�)X�-8��,��<:�GUzz�UhW�R�HwAT����-�Q��.=��J�Dܦ��,�u�`#Ŝxq���o1�i��G��f�"^���4�޲�pZ��.*悙-�7j�c�Uؾ��y5S�*a�����3����Kv��n�<�*\�O�Əs�#�鳽��Ki��돳�W�+~"�}yh�M�ȧV�6&���)�ֶ�OzQ����;�Aؼg��o�[uq�r?C�6ׅ{75�g�]�z[��_I0C�tz[[/x�
o�2�1�d�o�����#E�^��wu#A;���4�X�+��2�}B$F����`����~=�9�tG�4t��T�㪅 �9�d8ml�� (<�y�;e�۵���}Z{��@Vn;Fm_�v�={hd���.q���3�-S`m�ئA�z[� ���Yl���vz��4S�H�#]*����e�n��a��$dی�*PV�B�\��)���5�2������,��	�L��D�vTB��� ��w���&Jk1j43%d=�Yة���� x�V+q����cz�g�w!�t�*W:Dz�k!�ȬW�:c�s �%u�j�Hܩvꋨ�T�388Os�q-���
�K���8[� R��� ��wpqkr���f��W^��g���ܙ��������V�r��)�O[�d�J���J<E	�_�p�A��׊�L�׻^1O�5G�ڂ����(�KT��oZ﯐�:^�.[h]1����]{-�=J9u�x��]�}bcw���F���F�׵(h����U3�>7�َm���S���Ⳙ���Bj]������]鷛Q�K�J$�e	܆.8ʓ���wܾ>�p?T�]������|��P͊�E�\=������"k�k^ءB�l���/z9�����s�ɋ�*%-J�V�WPX.�N���v����y\�T�It��c�ܲ��;��}�}�"W�5Lwub����*��vV�|4�^y��]����޶�8.��qt�"�U�/�R�>TZl^���<�u I|J�c��r��9���~L�/���������R)�7�����0��:Y��r�32�=�K�w0���D�(�5]욛����;V�F�<��Ӻ6��^����O�p�r����M˲�]���n}������HG=��b۫���g�[��m6znqPɥ�j�U��vcn�[�]���j���L: =]�K�	0�,Ju��htqaºe���^��}��"g\��w}�YH��D��3�ܘ��fԋq�SWw\B�*�-yվ���|�WG��<�:���!,"*��<T0��7uZ�Ŷ�.ĻGN���o�&�	�D5�6�LUt�#jgP�J�����J��M�ɑKP	��(���+!_i�����ܥK���Z1�gq���0\Uݔ��i:�9R"��P�J��������[�@�Ď�Kֹ������Mu/�B�S���(�� ��[�t׏Hg@B�]�zjG2������֙X@�۬ٚ(��M)��ꯃ�E�҇�i�},/9���I�u�x=�#NK�=n�H>�ضw/ H(��Ǧ�P�$\
q��L3x�w8�75'�In�Mr<�J��휼��W�K�/���V5w*��̙�iBò&�㹊��VQ�R ��x�J�y1����z�*U���Vt�AJ���:�.�З�cŐ2r��&�n�W��኱��0��
���w�����[����,#��2��N�oM���T˼�<L�U!d �E�
81���1\#���"�3�����.�ùu�^��v�y?�'
�$p<��ٺ���Vn.�Ʋ�+yR������X�K�OC��[̫Rܳ�_*��DI��m�0�eSF��1K����Cz�ּ��^.*��ٮDr�2S7����+ VΦ��;h=늀�z37b3тq��F�hh˖n��f��%4�a��5B��=�����3��]r���C*�3��D��<7ϴMVM7@ĳWCـ	e`���دs]6�@���8Gq�w�N�-�I_C��h��Iz;����A8�Ʀ1i�x��҆��W[�[(�����Bު�3��n�_+�6�	�7�L�;�V`WLf��[�+��V��v�Wa��;/��� P�V��i�&ɴf^f0�5��*M�Ȗ��ϰjΤ�gs�q�ʍ�ܦX>�.�k��K}�#{���efF�)⻽½�jop�{uu�(	0�A��޺9� 6Z��h��yk��+�������_&��'3B�:�~�G6|3�2k��Y����8fp+f�ܷ]�P��^��;;�ZގJf����6{~�j���0��sZ9E�RM҃!ܰ�wtH5`Bh.�ޜGP������D9}��;|`�)��Y�sg-�b���|D��x����`��F&n��@�E��'�36F
����zA	��gY� sAr�����"�d��-Ds�j���p���oV��4{t�+�^t�a<��e��T��9�Qu[�.i�Y��Mm�4crB^�Ϊ�r�/�cV�1i1D(b<%YD!�{ޟ>��@���!��s�G��x��A��ة{��E�n�\]܃ �_-%]��e38o�k���!�9����HĚ܅K@��>b>��N�p�sD����	|9�ਪY�����-�)2����v��AJew$�	�S�;��AF�
��1�w8�b�����P��0���`4lb�oT����B��#�؇��5�&!��9��e�R�׮!�kT�ʑ����ʲG�7�*�% ^�[X�U��0�Χ9�6���m�;���w�bEhˮg��!�5��~�c��ĴYis�
�aP�u���8�ӹ���:��Ň8vY���๕4ԚA�����W�imA�n�Ν!H��� �x �ޣT7�
6q(|���u�gؐ���$7ڧ�]��,݁sz��v�Y ����mf([1����r��W@���+�79��cx`�w���Ǫ�����.NZ[t�2�*5B��U��۷۰����2P9���뽋�ɉ��=�í82�L[f���\4QMǍV9���ge=IAVE	�wN��Y��b��|}|̫�	{y�����#j���W���4��.7�"{�\��:��$�GT�%��nF��������g��m�&�6�g;�
��w�Z���u�]���9WO��Gy���۬k[�ܴ�O!�^z�fyxsI��E(��O��:��v��v�gI��4�1�1S%B�q=�˦���q��)>.�vX��59�R�}�pPiɴ��wjn�sQa�c_n���p��L����d�s�`�:X�pR=Wn�Sd�#wBeZ��\+N�f��'�n�]�[���[��~���N�>�7���7ہn�*:^���8�3B�>�a'�cu�:���i� ��t��3-����Z���x�N�	��iYz�D��Go{d�{q�u���G��X���B�{����{�s���Z�W�a)�7J{����i_w��P��wC�5��F>/�6�,qQ��fڰb%��vY�����5�����Ox^.�u����Oʱ�~��eMθ�^�lM�'%]��<�ѵ��$�Y�X��Tm�Pr���qނU��&�|���Ѱ=x����Vu�[y�H���:�=:QuxYy�%;ȯ1�:��Th���𒱥+�n��jU��6��^�ױ���%Ҧ�\�(���0���L}�Y��Mɗ*��Ѿf��:�J�י� d���w��}�#n��LsA�O�Qŷ%<�L�1��[�uw�oFx�ժS3=�}$�W����E����ِp�h  �G:������tń[��/6�'D�CmH���}g�Ps���������GRju�Z�vA]A�ή���6��5ǣ$��nY��#���#��%�sl3Ky���r�q`u��ӥ�ȶX&)b��w%��hH�"��@f�%� ۏ���
'D�r��Z�ZJ*y},eՈ��T5&��خ�5<�	��G%��':��x�luOm6n�\p��]
8��B�����������wB�R�(#�q^�O��x3=�$�+GQ��ߨ�##yL�4#�P����g����>�®��vU�O`����h�'�w�g(� ��d���3x�����+�;#x��=ge4mĠS�p<F��n��a�{:,�D�]�5\meJ�Y�J�M�4�P�Vn�͂��0���#����i5���u�ZeN�W�i�|��#��.�.�AHS��r���F<�v��7,G��[�I�r�u�U� �K��b�FkA��n���Z�K��i�Fk�{���zv�r��aTud�kR��.s��]��!��s�1�>�������ڲ�}�90&��]R����3���eA(	r8�erb��R�����kk��b�+qK����D3rT2 �e�e�6�-|�.�sF��t�ښ� �\(S�������'��-sĪ!t�i ޳JͰe����+��W���Ӵ����׻�p	,�}�+ �h����=�~m�3h��0ץ<mI|������������������vk��,|ŵH�=|�zh
\�Xe+�W}��Ƭl4�,�V���l�Ve6{�y4�J����沅�^�λWP�o�^$��FAKܯx�}�f,�%��H> �kr��Ro-�ӫF��'��� G1ʤ2gp��Y{i�����=�̶�#y�J�t6h^5�����;�ʲǷr�CAkD�j���C��+&M��Z�n��[��FHVu���nȫ��H21S7�7V����(ݢ�N[��'q�5��!�ܽ0��^��ڳԗ_�,� _3�cA�ٸ;Jt^��Rv�$F��q�n�Vo�-����3�}���[�S�@�yz�θXGZ���)����1Lc�w<�@(贕i�7҆�U����o���Zo��I2��w�yᷪ��[�&�z�W����h�û�0S�b�,r�+��3������(�:���k�Q�?��;�v9U��E)��;��A伬T�S�2�C�1�x9W�Xw�GZ�n�x�b�:*u��(]ǖiMsS4�U�Y��οk���LWa��a,��qEF��X�r�� ���:F���"Ԧ��A��](��,��n;,^�����7���q�|��Z|w����Q<�B�Ko��ϥ*�wX�� ��F������Q��T�d��(�}�_f��k�����<X�c;���q���0Y÷F >��02���ND
=��Nۡ��S�.@��U/�sf��J��}������tk�b��NH�Vw�-ML��U��$��vo��9���O1]-��8�/�����fjD�~1a���⤖b���QF{M�v-5�8�|r��D�sJ�cq23�V��������ׯi�GWTxU<w�{��Er���M�z&�>���7��xy7�k���7�{f\"S6[��cfnEQP�yXt.�M]��]b�FmV�W����yԩ�\J_,9w�J4zh�,�����nB�-:AA��kYH^�����1&&#2�V����RcV\�cf�r{ �glf�%l%=�VWdf�7@��i�,�M�
w%Y!�J�h�M[��|�uX�y@�b�f9�Ceڣu�%�k|�9�=�2�V���)�l�a�l*�=����j�fT��Ad��8�k�|9Ә3�����q�xs�7X���
5���!Ą�sJe�gٱ�]�޼�Y������YV��GK�I4�7��q�jn]�N�q!7���-9ɺR�>����L�`޾,uܛ�W.�E�w�=>�N��t���F�$mX�M��:�Sw�U�Ci��|��ٽ�v��@��4%T�|����>�R�ۭ���P���;�s�e�-���������RVժ)o6���J|Vv���ُ�}ݸIKc�P��nX�b�uM^�K=�TX�v�L��G���&�B�s{ M���#�L?��5)��B�}����̧)W<��]v���X�����@�*�&���ꨓʺ,�۾|�̺��Rf���&��yQ�g�*�m�#O{G`;��m+������$�z`������[]n�R��b�e����{�>LT�w%c̗;�+kQ#��pS��q�S%背�M��٘��<=��ts�;��6�:1�3��꾜�(�,.�ulθc¯n�
2�]%���3{�ُl<�ӟr�]��{�΋�si�i��gf�w�f�͍fۆ�J���۵��ٙ� ����=tJח�I�栥�݈��»��4oN��;ƎH:In���C�$fg=Kn����`�lv�,*
"�G��n��Z=<�b(
���E�y�QWQ;��=Ty44S.u.,����v{4�ͻ���/�qb�f�]��k�����Ľ��|i�5&F1r�G`���gf�ٍ�N>1rF��^�x>Hʾ9; ��1hU�ˮ�ujp����۩�� CC�,���!\%�<y�x�8�("̪Hؕr8Y����[��
��Pb�QE:���3 ��ȮgK�U^s�y�����CS���U E�un�nQR��T+�D�!I�np�^)(���-6�U�p��9��I�r���`���"QW�'�r�fȂ�HArN���RH�9��^���j�OT�eR�(�UhE9�r&��@���J�D��(�9��8Q�
��9���:�uq�tͦ`dk�91),U�K*ISPī4ڒW2�gLD�3E	n�Y^R�R��*�!��$SP�D�I#�f��s4Ȥ�3'�3�\�T��XHNW6�Ik<��˅�K$CEKeI&Fċ�RRek�8��s99TS$P�i�p�	��%���☞�ψ�-�4��e�b�ٴ�;��U�*�>a�!;����Ɏܹ����u��v�j_)�Ze��%s��M�ڪ��Է�9���Vf�e��ɪ�Y���de˻wz�I9vD���2�qkK���S��r	^,cԲ
�څNN�v���i��b��)�Cݸ�wL�X�M����'�\�&��A���:�MI��#�|r|i�a�q������@(؛y]���F��>�aل�N�����5�s��&2�1ч������c=��y�NbRH���꽶K����ֲϥҸ�)�3�ՎY_#HkwzUC@7�v����f�/���ս��1�W5�─�|00&;�"�y���]&VS��M�7���Q���/fr������P:���Q���������N�q��Z�`e;�oc�t�){����]�Տ�����ݿfKf�]��CY�{��b���~ʙuC��f���E���"��Kb�*Bۄ�\KT�,�
	����Ȇ�z k�jt��Ldޙ���.F	���.���D1��θB��^��J @P��z9�"S0��k����%�no?c�*�]��/Q͙+t(�ڦÙz�t(eXo1a���6�~�WP�����2{�Ly��7)ؽ�d���]x"�ݎ�����l�oi�_Q��u��rZ�p[��(�s ;�v�j��Z\�Т�J�Uqr9�,�޺��;u����--v��jN�q,z�t@�4BZ�&�+KM�`�-�U�o"�r�k(	`� I:��q�"�k�8htvϧ�Z�u��H��o��ꘉk�5q�Vқ��V\%wcœe�j���Q�.8�%k� ГT��r�E�Nv}\�Y�lϷ|��z}դPb�����m���}��-4�����T�׀JR<[�H�y�5m�S]��f��ьa��
4�~�<G��m��y\)�qp�¨��B�s����@�_>�"�L�=�n������K�5c�OO����<��zy��rS۫�fHo}C��6�<js�%����Jyp*����Z��X�	�������\�.���w�~s�U�2��d�Y�Ѱ���>����q��s��U�>�#�Wf
Vߋ��٫8A���+y?cU!��cm4T�s����@���u*|�3�sCx�+o\Y���f��7��6�7R���n���ɟi�Vg��5 ��B��ex:�="���	s�<������y����D����Wbݦ�|���a����F��1H��B�(��S��<hD�'0��05�鑻�1�=R�]'�s<���$�q-�RXQ6���{��Y\�8�,s.��3U��2N��\�z�z�Xj��ͦ+P�&�|�����Ec�ó#ͧ�:�1��%�i��U���D ; ��9�Y�^Hot�ܺ˻��䦈���Um���e��j�
z�Z�Bq��KN@�;0�c9�B�[�ŵpgv��Z.س��}T��<���2�����Ƒ�����P�{�����G�n3���`nK�
L,��5��l}p�:C��t6�d[�#L7���c"á�ۚ)���'��H��TmUD����(_ЪX�mm4c��+`;x��x�������jp_xkTx�_0��_��V��{V��b�5���4����
Z�W�tk�V���7�%���]4���S\@�����3AT���ȩ�&�ϸ��4r��^F�_N��T��S��;�*w�p�$8�Zc�!��H&@L���+N�]{[�(�\˜֢��#Z����1�	��-��2m��ցI�2E��"c�au���.�$�W'�Z�P�9&c�y~�}·�����5��Қ������(@��(��z�=�YNn�%�n:�K$�Åt
4�{�f7�4��Z��M�� �˛�<�E�����u��-;����W�`��R"_d���t��E����W&8ӳ[+"�ooH�9;�� 0bkAZj�R
�԰e/���q�ۥP�:<rw(7+�v�ES-q�[�E5���+��Ě_R�ƛ�fL�NoD27����ωJ;_���D�i�+�"���X>�l���NB�O���l���^��=PhT�#�L�
_9�6�\�O<yg���l���{~~����6�R��V��A-����论�hOȲ��<]B�WܥN�{�Ѣ'	q�\!��Uo�s���#�l�fO���*�����m�})+��y�����qř�@Q%�g������<�f�k$��%���>c�w���~�c���N���+�҄��a@sQ��`�S���xE\�zoP���^�3;1(vzLkqw2�e��֐� �a�L���g�MѪ�`r�8nS=�N�5�c8�)��f�z�^��x��<]���3�̈o1LC�6F�A �l�����E�[��4k�.�z�^�+�\_��\@�\�ڱ%���=�k+uW��9ʁ���.g���s-�nvm[��v�O�_3�9��!i���R6ӻ��6JD�;%���㺲r�N��Q�`u�z�1l��b�n*�2Ù�2j�^��R'<�#����;���}=��(��|���]��37�5j������7��fx�SSd�-<�h�ų��S�}�PPn�J�����So�yhY-S�nuf�4Evd��i��z�\�E@�n�4�E��ڤsc�Z���=Ѝ뺴j��": �Ā�U�����:+s>\���B1�i�W��S��(V�UlQ�@W>��F����RDv�N�oxue�⸬z�Z���GxٷP5\n���퓳�	U��E�c%[5�Jv�*���c���O[SsMu����P���D-���Ӽ���?l$���`s`%u�����Ou[}w۠���� =�m\��Z��܋�B�N=5#H���<w��]�U���|�Fe��\79�� ����V|&m�=D}yO<�D4v�}��!�;���"+�g�d�R����������ӑ��M�F�2&�yb0��9&�����o�Q�y�/7ܢp�J[7�j�����V��e��J;���H��
�!��nȠ�8�[ru��٨S��G��T�r㶘�d1�K�q9�w����F/ṓ:o�+m�e�x�z�ϤΫ�=C)��	y�ʯ�O񣤱���y���^�yk��|�����s��ߣUOC5�b��{��.�;�7W�G�*���!�n��[x��*2���g`����ۅ����C�d��O���:����|<���Z;���:Lo{9vݍ�@��e��v��q�7r��Ldm�Gc�O�םb�٥��un9$�qG�f�T%R[����6�#Y����g}/��ن݋���ӑ�e�09ugZ���#��nZ'
�5����zC�Aj���;���L�J�x�־\��!��j�_��y�1q-S�+o��	�4t���
�Q����MSڅ��bJk�i�Bk�[�5%��>!���p��s���P�& n֮�Ikt7���6?r���=�?\+�l�_M9c��-v�h�=e���:�B��(��f�n�����Шf�����L�~(Q%�-�k>�2�T-uÃ����5��'����j��܁ZR�� �|���ƘeC�>�=3��5��W��@hʑ�C>r��w
�B�;��:篯����C�ٽL�lNЉ�1���[Em��B�̏q��0.H�} ��z����@��_�p/!�`E��W�]s~�Q�G�-��o*�h�[�ƣ���w�=�9��Ҳ�wm���#���I��wA9Û5x�$���Z}�59p�g�zU�ή�ǩ��tI��?y\���5;.����Ε�qZ$D��H	"4nv�X�B�lc�w����Z_[e%�����D��V�5*2nt�`���;K[�&��'uϭK��5�v�ys���Ż��>�0ljI��>��[�dh}�����g�{��,WR�}�y�*�����
��#'"�P��3��Yϝ�9GcA�Â���1xx1�h!�/njt8��`��;�ca�Վ�����\���ޒ���=H0ς~�UR>�1֣�MQ�:I��8�R��J�9�Y꽩�ev���J7z}[�ϲ���Kzn�#��v��ʒ�=>���A�;���L*�����+[�(�P �����_=�:�1�0�,5-�(�N�d��aغ���&N/���z��Gv`s ڮk�����ς�B�{di��Ma�ƒ%-�
�.���tO��.[Ύ��f��6B0�� ��`�9���7)������a�F�6�;��R��3���Nu��n����IJݚs]m1��1�>��s�����*�����6�U����5Z�!�8<<ITg@���eL!_mUD����(\*�0\5�ь}'_,�W/	�;��=K���x���\<�\�cהcA;��V��j�a���=#�a92��K�k�O[�n��j[WM�Z�l3좉5)��J�O֥u��	?��~{�7팶%��w�+5<!� �{�[��Oq���±œP��N�ҹ��(�Nͮ�>,����qT`�-*��H�i*u��*Æ���]y&sLȭ�n��~�vƜJ|+�&�3��K^{؉:���R��Z^dD��2����+ro-�w���fd�(��9��nw�[��kii���㐐%�-�ReML�r�����_ٖ���ci.�*{��8�7\�P�L�H��a��t������w�ԡM��Х�W^
��e鿻���Rb�I;2o���v�a�-C��T�e	o3so��~
��Q��t�����f�{ܗ�/f��#yos�Rp���Zy�[ػZ�o�I�Y�0ʁϒ�4�d�]��_����^�OT8�
L�
�H6�"�Y.G}��U4��52P�/ゆ��F�z%�*i�/C�Q�ʋ�y�lS�p��y�Գ�r���yy�dذ��Sƹ�9�y�x_��T���ٟ���ʭ4�D�fj:��l�[��K+`<��O\g"h5ƹe�k�U��5�c��_]���vzX��jvP-$�Ԭ|���q2��V�]7e �f#;�s,�t�yS�3S�F:!�u�<���V{����U��|�9�q[vcs��]�_�S�P��������=�no�q[[��s����>�
5�a�^s�mKo �]ǔ��	5�ʰo9�|V����B#�b/Q����Ӏ��R��-41�yX.!x�bu{�k.|�b�1]~�l,���3����I���|N���w,�{}��նf����k.p�tS�J"�	�n�xJ�a{50�F������l�l��v��ac�b�5��X��[�w��2BN_�M���d�kV$� O�؆��UCxs��~≺[Q��b������sSU�u�K1���!�{�#m;������7���&Ue_�@���k�t�=���ND�.��͑�,�:�㖫��2'�Q�1:�|5��c6�d�AX���"�i��J���қ���xB��ޮ�*v��^�E9��	�������{�����:�h�k�d�� ��w���9�2��,+�<>�K��1�VY�c%_��ѵQ�@v��KOz��-r�24Gjx�sh�ϋ�B��@�������r���z�Ԓ�K�(R��1�"�u7k��\�(ĀZ�}�KB�:K��S;j@]P�V!ƜMH�#ٝS�1]�jllk��)M$	����ω��u��������^�F�|����'#�)ޡu�8�s��h/!��K}��k<ZÆ����^�������;nB��������{��r��\�$�`��!��R��˄G/��t�<Aݍ�sq=���J5ǰ����M�g%N�ژ1�6h�hl�d͏7��Le4����
�{;��ٱp��Ӛ� ��a��m��0;Z��BF�8){Ku���=SS�˖�ڭM*�М}S�N�͔��d��B�:��n���B�#��b�_���8<u���]X���X��鑧�� 0�qS�~�R����W/��5F���{�m�MPV�%oJs�dxib{�۠շ*H&g�X#1q�����	�W���;�(�I�WD���؛3~9��/^O�F���!o�\��Y��d'�-+#`./F�w$�<}Z��Ùn�/���۴O{�	�ޢ�]BF9A�ϠnT3s.�V���	�z<�y���n=ą�<+{��&{�~	B���!���ۄ�_��1���,�����ƂMix��=Qs/%��~��=��?Aip�&��|r���D1��θ@3l�F�A���0fp��˻�x�rKd�5%?_]Seӟ����X�q|Nq���N����V��v�^^,s5M>CQ���'I����{؞� m�a�C��}<���wFbG��y��v����S�ԟ�B�8>���1�:
U�+4!�"^R�G;���;���/j%g�8'nh-?sxX�oǽֵz~#��������S�7��o���8�[b&Fb�;����T�z�ڈ�w3+]+�w�C���Wzq������nyn����^��(ׇ�繴֊K��YǨ�P�Ӏ9sUpwYt�ל:%�pM�-�u���={c&�z):�������cf�+��v��Gw�z'�,�|�K�\hF�g\����� �o0[���R��&tH-:eK��ˏ"G���!`@�]���nsi1��6��g�ԍ^��jPتY!y��cv�q�i���^�V�yLL�L�{��sY�Ci�;��w��.�X�7�l��k!{|AKv7�+2���_V�1��;��oeI�b�[Z�/@opݙ�NBS�<�����['�w�XK�]w^*�I��$��#�>��KA$����6}hr�t�W�4��תө�^k��	����������:h*�Oh��[�t���jj��~I�5%D�1'Y�ƃ`���z��gB4�pw�ܝdr���Y����#��Ή�m�bv�Ήuz{z�c��
�h�oK�[�6����5ƨ��k�d`8�oG]��g�;�%���5<AC=��ǎ���Q��S���$��_�D��X;h��@йoG���GSG{rrD^_}4dV�ӊmö��4�,[Ի)Ի���;��������ʇ��6��a�*��Ǳt����S��ӓ�7���;�[�u=]�%X|���unW<��vs���|e�=)���V�	��X8K�"�WZ�B�%_e�a�n�w�{�]����`�K�Q�ǖ5̽,�}��inK��AZ�7�L��V^��i�����uoT�#BuEHѼ��+�Ӝ�A�6�
���	���K�,��jq��V���P	�$��r\��,�����xo��+rVMgf���]�x��4��yj�WNv�mf���x�D�r��T�sXqJ\\zp����.>�J��u�8�6�#}TD��|ތsW6��t��r��m�ߒ��ރ5$��N�nI��J�a.)�a\x۱�ؔ�^~G��J��ױ;t��nL��,k�'�n?���R�80�t3B��z���I�����������a�s[q!����
�k�� S�֣��(+��t�[��}��2�e������ W}��a���8d�7y/�M2�=�GcзXG�U��I���;�A��t]`ǈe�[�ͩ���VZ'�OT����AJ�;h9�za��º���]�!g�4�h>=�G����C-��w�>�'$r��ױ��D�2��U�OZqԀWZ�n�y����11���M�f��;s�H�\Z��Ρ�ܟ����dF�Զ�GV�qW>�&�qRq���HG"�-q�J�r���II�a�,�M�Y�)� Q��s�&t��<Nr$�EEUIY&Qp�J��<nLD�QJ��7sH$��s��	�r
�2L��@�%�ҤP���jFD^0𩄝
�)C
U+gB�A���I�2Q
���)ag-:��\.\���D�%�[MΥ*��LH�S�(��P���$�d�����N�Q�U�x��F��sE�� ��+U*�%V�*��uDTɧL�H����A��U�R"t�K��1�IXh��T�CʋV�
族qa�a^	iT[JYbbsX���!R,&��djVaGJ�����jXF��e�C�����35$.�r6�f���dZZi�X��3hH"$Z�Uer-�۽F V�u�[a�m�J�:2]Eu,9�� �-=���dQ�gn=U�X�{om��#i#u��9�l�8���o'5�۽�c�q�����e����
�~��(I�M�
�];���GHN�]=���w�7hq�J�]�c|���a�?;xy��@|G� ���_|����";�imY�!Wm｣���p��c�D�#�O�G������=��n��V��;}O��ݤ�z�����@�7���ٹ]��bwG^p���7i��;���?�Dp���%8#� �#�=�:��t�#��樥���k�A#��{��>�%ێݞ��S�~v�oS{�v��'N��~y� ��BI�y������!㸟z���p�m�i7��8���t��	����"HG���� �͡�k&,����ԧ�G�"�DE��#�{Ӄ�z��q�=�޷�>&q�p:M�'�s�#z��N�~o}�ާn'~}_ct��$?���\���I�u���>��KV}� !�jr�d����uˆ�r�E����1��L��������2G���z��yq�τ��[�>&x�����㏏�8�_����(z�C���ۯm�N��>{���$#�a9A��8C�@d|�k�};R�����^�t/R�~�� �>���0�&����GJ��i��x������vw�t�;q8�|���ߐ�]���G>F'x�y�]m��>&y�6�����{��P=d����������'*����%�C�|Y���F�����t��q��n;��'�>���t�UߜtW��q0����}v��$��k��C��y�&�	ӵ��t�Sz���:�o^����~����/�����Չ^�u�����#�(}ޞ��ӻv�}O��?s\t�ߏ~��E�D#������ Y�6 �]����#�x�i�]��>!�o�$��<��N?�<�q8�w�<�E��s��^^��Ϙ���"<}�ѻ_li���L?/��_�:޻v��!>~�������q�߼��[t�+��㉾;�~B��X:w���;����S�����w�n;|C��P���jafw
�d]W�(/��S� }��I��w>�_m�N��sލ I;u���n���n{�}��>&O]�#���q0�G�|=��]��߿y�v�]�x������<v�qRv�x��uC���*�������d�of#8k�����}����a���o� ݵ���$���u�\�.��0`�{�M�
���v~f+���|I��)��}�n�{[%m8���9G
γ+ݍ�i�k�����I=}�w����(i��0�{0�8�b��YS��w��ǧq�V�ϩ�a~����׎]���6���&���ރ�z�r��{�I�'������8��O������0���9�4�8����5 ��,�>� �{͟�u,���٫�����8��v��,;)�|@>��4������8�a�=[L�̈������?G�#�}�xz�����p�-t�V�w =C�w�8�S�A�	7����7�q��[�q8����n&�w�����8�{�hv�z�v��|�������z���}��o�w���}">�ל{�f��y�wR��z�9�q�<M�{�\#�����v�S���_����P�n�>��uˤ���'��� I!�徻�~�۞F���ݦ~v��｛��c{�}�CK$�]z{�RO��UݻN=<��;O��<w�{&���v�s���F:M!?S�޹���1;�vy][q�:@���j���/�`\��y�����(8��1�h��e+Z���g{sƵo:�� ��v���z	�
��=�ݾ8�;c޹���}O]����>�n�v�{z��o�N���|�#n��#��ۏ<�O��n���=;�#�N�G������g;do���3��>�>'�W~O��ɯ�����ӿ!㸃��N&!����o���!��}�I�!&�	>oz�F�'S��s�}Iĝ��7i�����B�{��M�#�>��t�����#ɗ�+���Q�w�=��v��i������t�+��[|w���6�7���7�~��A�#�M{��qӺN&�p�ǩ����=�@QC�z�/9�L?����.��\�.�6�$���#�@�OX����nyc毈t�]��s���a�?;t���;��'I���v�?���!?]�߾t|L)�B~����'Σ�^{�ܭ�zN�~=��a�o��c�]��G8�>C�1����:L.�{a��ӵ�>��N8�}q����0�������}C��;�=M����8���� �/����x����ʅ��Q���>��������j�Հ�x��	��R��G����g�_�DE�X�B�������&���K�?�+��V�|���,:��xL��U��2��sMC�r�ad��[ك�
�7ۛ�GR�4f�k#�*�b�F\DG]���D����]�9�k̮��k�6䗃��"�Uw_~��t���Π/bwN�z�������.��C�#�|N�t�W��&�8�C��es�bw�~w��}C�v�]��;�z��ûq\!&���J��<���Lnz)M&����-�hq=���׎�=I��\�I�����O<���4��/>�ѻC����|���|w��o}�����N����t�������	7���9���bw����؟|����+�t9ʳz���ג�}�����pzwqߜ}N8��O���:We?{���m��9�w���@��uso];��n~�}���
�����c~C������W}v����N;`��z<#6=P߲˺�����;i����'���t�7�w�����s�1='�ܭ�'H_Ѹ�]�7���}e0����߽�����xw� ��'�8���[�I���>��7����q>���m\�_���fߴk�Xҁ�`4��hq˳�e�O�8�ԝۅ.[�ۉ�!>��n���έ�$���Ѿ_��۴����_|�����{>�z���Į���t��G�H�C���ꫨ�ͯ/:���_���������}N&��C�wN�8�,q\HI��nYL>F�Q��H$��N:O��n8���!�i|��y�i�BL?����m�>���>^�m��1G�gg��o;��ĝ��:wn�����B�m�>c�y�\
o]�����c��F'x�j��ӎ;��g��8�q��.�
�(�
=O�q0�c��q�;���@Ϯ�(}������܏Y�C�9C��;�þzn��0�{�:��n����o}�u��ۊ�>o~���'��^?7�x~v�7HO�y��j�S{�`��ۉ�,�]:v�o���8�;�j�桊@ G��y��뻝��|oG�j��K�E#��#�}ｷ�Ap�>���=��'������^��'�?!�9Wz�8�C����e����޶��ĝ����w��;q7i�q�v�Nj?@ ���(�{�y�1j}q[�����t�'S��Ӆ��2ɾ'���%~�
o�qO>�����N���������z�L?��7�]ӽw�q?��t�?��vy�=C����S�b�X���b�E^�q3ޮ�B���QZFz�6�����eoa��:��F=����ވ��UY�i��U��3�1�w�����:��N�iZ��5z�ͣ�wk	/wz	Z��2t<`w0�"{�ۮ��#���3n��ݝ!��wJ�0Ii�1*趛�N���<�F��E��.�v���Ϥ��W�
���w�����i|�ޠ�i	�^�;~N�۴�wm�t;z������7I�B���~�J�S}w�~�i�B�1'��s��?qާ\�'8�8㏍H�(�Ǜ}�=��?�G� ||��v���0�o���t��I���v�{叴u�7�8�^Q���7Hq��v��?;q]ӻ߾�;v��矼�}}����~�]k�Wb�^�ItQZi���ܞ�F=D�� <��\���RT����Ez�4�u,(�Թ��#ѽ�iD��!%W&������������妎M�qN�J꾐Ubs�T���|�w�)�3z}�Lh����%�9��M��m�uB�jM̫0�p}n����Í=)�|��&}�gչV�������u!���*����p.�|���Lf�-��͵M�|�N�0�a�*M��P� <|�O�\i1��i�m����n�r;�Z�(��nT��L=���?m��/�`�a�:�k
�%��A��8������N�����Nl-�Q�&��տr�Z��^q���R[����������N�n �r'������;�Ԕ� 8w:���L��ч�W���=�P�̻IZ��r��ǡ�؆�����4[�}7L��K�y2�����9uJL��PLVa����3g�$/3�	���u�Ј.��J��9��KgN��}�'��J����9��Z�P��>m�gR�}�%��t���s��N���.o|�U�a:���O�6qj�P�_��#��M9$�걅��h�Ξ�h�=�L�}(k����g��1(�$�L�(�q��!���g:�V�g\�8����D�	�:�[�Ie�ȁ��y�_��2�X(�\V�K[!�mD�v%��C%X7�:��}uI�N~��,p�p��H�Rt�,}yp%9�D�n̬��D���G�7]Z7����
I~	g[���xl����9��ʬh֍��y�-�i.y۽!b��{P:��w(ɲs�B�CG��9RN��t^J��r�/T�q$�8�8r��M&�@�uo"��!���[E��	��QDhx\nr��}oy_P��1��d��k�i�p��(��*��7�(�(�X�w&�t�~x��eFK~�1�{�p��<�����V�2d�6�y�����Ǖ�Լ\�l,�o:��^�-j��_�	�z��;�͢�ӟw&�>�K�:�_�&�ܸm;���9����P}���-�OT�Nw��;$(�!Ԩǣ]$+����ɠ��T�#5:c� 9n���S���E]�|{c]�<�\n�c7!�V���m^,������Ý��X��v�7�u$�Bm���6�����6��t���4��:���ӧ*V��X A��3w�JS[�/����0�p_J;E��.9�nݰ�᧠y2gwg)���\郾��/��z�O�|o�م�SM@C��@�u�}`�evk�{}{�tW{.39���vdz=�ڰܽ'uQ�����>�V�}fx�4�p�ر������ p�;"媆��F,2{]ѧ��yMx(ւ�9���Ŵ��4���헞i�����h������`��ܫ�u�n�aYlW#^���yMX��
����oc�^�X�� �{@K>��2�o�ୋ)�p5���e�l�zZ���C8�ۋ���3������d�<\V���_��1Q3�����d�	�Z폭�t�cʿ�u�ATڋ�:OH�/I����x� ���ZK ��VbD�j�"�ƙ}/l��_Z1p��Rb~^|��Y��&����,�c
���k� |/�[�I���0{T{&�L����3�\u��j*�El�GnV�m�M�9�6��BQ%Nq #>`�J�c7wn��o�1ݫ�̈́[|�Yƴ���D��'Is:!���k�����Dҙ[�#���Q��	4pQ�,���lԤk��K�,Y]���z���IX�>�F ��h�g.T,�>$�aM�^�ٸ��ٻFZ���wQ��봆[�u<�W�u����h��"���	]��2�/�U�J��u'� �@I�s��ʕ8X���N�	����עѽ̟��3��#{��$V(#�u�e#�cj�r[1����Kϑ���d�@�׭^��}R��P��t�]ɮ�P�`�PXcÙ��W�Έw�|jLW�'fM�1�tt7��5cIfNQ˽�^��E�Ï6s�<EC܁FC�Ԣi�7��7��,�h��9S�Y�\���I2�N�MBS��a��%�1� ����R�ZGY�e�ᘜ���;�%ɩw9%�#o�Dq��'�q��܁���D�\�mX7�Kjgg��G��p�F/G�I���W��Aę	�J��/]T�U<c��#R:*����r��9�.��3<n�\��yvR��3qE2Qb3��GW���D�q�Y�Q��uk}�U!fq��1�p�"�w#i�{���-��������s=�U�'d� �gFr�S��ȩ��Z�tZ�
;/�@wi���^�3/��;Zf� =gVO�:���
Z1�^���57�ˍ�%�0t�z��,Qb�Gې*�o)<�-,�~�|F�و#�"{	&�v�њ��VPpw'6T�I �)̩��h�,����+˦��#:��E��H�r����70�Yl��`Z�jua�RT*�]�0�;Ak��<���֕gF��ɴz���tA(����V����	��+�#��(�y#��R���;�;꯷ZMo�w��5�y�c.�n������`�)G��[?�CY[�e�+!��P�N5��sW�0��?qR��5%��{D����f��=��-���x�5��o�ղ����c�8K����#S�ߘꇶDH	��R5��-P��=ҍH��5�����g��ePT;/�}%���Q�?��8B��-���*v��^�E9��Pۨ��\�Y�-L�*� �|������kH��J����5�5>��W���Iu��9j�#f��Y�7ǉ飊��Z��5��u�O��\U�2ځ���^J�5����D�17�w;z�������\K`�5��z�~�1-j�GiX]P!�E�Gg\�^�)L�Z�*����R��F��ꞛ-M!ǌw>&�P:���p�㈛�(�AUU�%Nz�jT���%���rJwu���7���N�NF�@97��ڞݽ��s�W���TC8x��H��л��TS~Ꝥ2�^��4�7�>Ѻ�R��/��|^m��wWhFd�+Z�D W����V �]��D�˞#� +�gmo�_-��i �D���Ac���L�9�&!����U��l���'W����[��j�m�Ƶ>�_�Rp��^�VW�xW�Aj�K�I/����vXu���ܾSh���}_}@�%<�w�%_T��WTy8�:0�^�>J�.4���Ɵ�j��=���̕���8�<T��_/U��!&�:A14�Xc�%�)�x`b�g -(�����&�!Ћ��X�۞Ϗ^��g�3�m�"���������Q���M-�O�o%� �)�������6C��/�����F��T�I�φQ?
�ĝ�&��+��.\����R s�#D0�~U<i_�xs����p�$�i����y��ODvgk�H�b{���	i�R0�5����jK,X�c}P�8ˆ'�H�=��K��5I�C4.4��@S�����6*�j���-v�h�=FX���ڭ���\�|�L�k��dh��P�����
I~	g[�Œ�/c�~�3�$���?^�;=�"i_�7�o�z���A�W�>�b��H9td�~YцCB�L⁸��5�02�����D����2�3�<��&GD� �"�'-H���S��bt躰��tv��η5��]Zv��K)���Y�wʹ:E��i��ڋ��C$�����c��-9w��IK���B��3�jw8n���U-�ة��8��6��i��/�N+hGu����6sǰ�17R�(Z�D�{��q����視-����p#����T=�Q��C&�u���f��E�����㙈E�}Ҍ����5[�{��{�eɢ}|������~o<Ď~�����2d�6�xF�O� �� ��s�+��]2��e��h@����Kt��^\,���\c��5ˀwZVZh��f�˽\�����"����a
;a�F)�"i��mA�&y�;�=~H��a�\_���ce*�ٳ'�j,<�o��2��;��}c���^����׫�f��D����H�QB,��_ܩ�Ϲ�v��o1Xp�[�=T}Y�CtW�a�C�s��s�\9K;ŋ$�2�$O�΁�ςۣ�Ok�/�]���[P�̜=9����ݻե�G��j8�mo�n��zh���x?w:�^�:��e�����+窶O
�/:zk��;^�.z�(�0��[Ó��1"5�SrA��*aL^�g�S����Mi�m�6�Wwf�&�u-!Z����Lk �#L7���ٯewo�����q��)ŋ7Nb�`�� /)v��5����{G1��;t�ʆ^�����m�wM�h��ٌ�kÙ���a-�B�q#�!�Ɛw���D��bM�W���z�%���1*{��v\1�CF�_L�T����mt���VȆh�U��W����g�d�/�7�cKUnE:�+y�j�$6��&�♜j�������^1{���oo�p��C�Sm^�P��qB^���+����Becc�Gq����!�����l^EQ;�<�1��C\��a|/�����M7#��\��w���Au�����IE*�Wɳ��Z��]e�}��Kk��A��kT�^Ѽ��T[����^r9!��E8�z�# 	�V*l7f�Q�4Q�c�qb��-
��iH&���\|J&��\��9U��CB�;��b�M+�N4��OC��w�_:��i麛��qw}�vW7 jM����+����F����O#�A���L[��L�YԴIz) �����m����h�J��O�p쎫�����'�g7�*/�z��Z1��
�$��/uz�2�f����XrNm����ե�0Ɠ��qv�G�$��}�C�oܔ�q��Grm��DQ7�/9�K*^���1�06�r]�Z:����55�.�1�C�.��Ў��%�y�<B���Ҁ�:�ǚ4C.�:�Rj�fd����{�[��N��z�k�b˛�s��B;D��9�"���o��674��f�S,�3J����6�z􊷉����Z�gPW����R�-1� tv�*�ܖ�^�p��lNg.���p*�fP���UZ4��v�vR�_y<�p���XsFI����AM1���:nhW�,���Mc	1�$���G�rlPq�tȫ.Q�[���s.��<���JrUo<��{���һS]iJP����ò�K��VՋ	�581���;���-K��Pu27�na����&
+,��3�T,�q��"6��YY:�5ˉ��+y+˾P��J��X�qx��&�:r��9�ζ��wV�َ��n��Q���"��ޮ\�Y�x�ܒ��,Z�»Y:��h]F:���3t�ʗ���C\��������Y�7&�T�i}�q��0Rc���{�0��Wsxe��ϯ>����暛7�� Og*�sM,���쬄N��f���.h����ZZ&�q�00��~[zh�Z%�m��)���56c�+�7KbtbR=��B�1r�s���n7LXW�[5c�K�:wK3q֞ݶ��[�E�[����*�ג�;�z(�a^s��AU�Йs�%b%^�cR�F��R`e��CC;|���b�Gd�y��-��e������k�����A�̒M�ڼ�`���4@����}�����K���n�C�`�dT�]�'��Ÿ��^^Ԟ�܊7}�ޚ�k��(�v�����h�\Jƃ��S�t��;q�ӊL�a��������@�|�$P�j��jt���ΨuJ��Q��b�r	h���.TFE��
��QV����q�J)D1#2�T�TZK�-�M*6U�:
���-��RȰ�ĉ9F�H��.��Hf$b��eP��(�0�P�Ki��Q�h����	k@��uES	JL� ��T�K@���*E"4P�	M5��-U5-!J���r%S�FHX��:YU���̉�NY.'86�ԄD �SL"�s��p���*C,�DE%�"�b*�УP������ZuL�JBBE!S1+�-1����"��h�B(��ĵ� �:I&�$�%s�YJ$+KD���-��L�K�#K�EN&IqD�<���ʌ�Z�*�a�T�JmZk��DIE)X��-�Ӧ�G9Ha�CkL	I���8�[2DI���IR�gNf�1(֙K-
,Ȱ�
%SD�,�:��2�0ˢ&Z8��4B5�")�A�R�Y�H��T��Q5Y&T�Ƞ�P����}?=�m��*��&��z�c�oE-�)죻0U�F̩pj�̣�uTW:}���K�����m�Ǭ|U��I������x��ӝԄ�E~�.�]�ֈ���$�xH=�.CM�D�:`��md\`g)+{���8og�����c���zGH�Mߓ	�d�眷,v��끗O���=�k����QMS��jr�+���O��&�.5�� �I!p��z#�u���Ii���1�!��[��$�#��tCG�`6���uV*��d����-^�/�z�{���[�(GG�q���R�B�n��l�a�h�p�hXU��8ɗy�<��p��C�S�lfrW!Ŝ\��<��s�|fLo�'d&tJ��r�sn7:sE�\@�΃(���e�����QZ�TX��w}>�<]��F	PKU�v�%]-r@��q
e2������,�i��.Ϗ)�>��u���6�s^����n�P#Vb�t��[�y9�v�� �l�"=k��(ߘ4ڏ��V�s����KuzI�t91b,T<����Z����\F:�;�燽s^c6p՝5Y3E�?��v�6*�ˬ���@��:�]���ݥM��1w�]���o`O��9�U����ޫ�w���N+y��uj��j������ʲs7*e��Q��[Ҝ	틲:�MdΠg`E8�5w��3� v�T�}Z��8ڼ-�	���� ���>���p���ѷMڰ!n�`m���$r��:���׀y�!��_� �VT~cjIW\��ST�!�o���FDk=���on `w:�X;�2��pv9[�r��|����d@�rU�"H�����*�Z���C����Cb��ǳ��tZ���v���e,Ŝ#�m&+�nT2�$T�g&���b�B�5V����_t�ї��y��v�C	�1��Ά���}q��;0�Cě�#�k�ܣ�I7�޵s�l�g}S8<�g酪����p��zn�F�{;�l�Q
@Ӌ8�U�tN]O|����7�~�T/m1/�ʰ��m\U��xW�L1�s���n��wV��ظ5����S5)�@�"* �|�6�lx��ȡhe�}r��Orl�m�`�.��R0!.{;�����T�{��6�F�F?�B�u�2"ez��O~x��o�뗣�[k���I�.�\\j��(ե��+z:DH�5 chg��m��=^7.��0��'$�\�J���<��x���?J�2�9ñ;��z7V��K��˫?��[��w�4\F�ےA7kzGU�2������6b��}����-��:}�o����\�^l��Wi�{�xB �s6�QJѣ�̬�[�e���r)�V7���ꪪ��������($G�8��	*d�fX�W�sq�j���v��b��
X�M��rњ�|�+�JL!RỆ"�<�15W&�<{�K�pnB�+��6��xZ��;���N����b��<������`�ӂ�;�AS�K*�AN�`��7��P�I��N��L��s76A4o�e=���M��/�nD�����vc~I�k9ꘕ��S��U��f���4z1�*T�X��a�i�Fuz�>J�ޓ�}�8��-gGv�$:���x��L��1��t4�kwPPj��!��UsXo�,1_��$��Q������Jl��W�*P��u�i���[��(�Y�U@?P���E��d�w�y�_"+�E����+\��1�1�Rg�o���;�U�ќ�H� !�X��-x棝@5�a��F����Dl�GmS:bƈa�u	�Q-S�����MY�{ia�Z׃oո9�v�%%<zK5�2a����)ņ���]�r��cv�a�)��7�Ac�Q���nN���<�nW�y9�ͺn�A:L�#ƻ#޼�4^���VA���R�j�m�O�bt*s+]�nn'X��LCváv	"0��t/{^����6�\hg�珶Lr?�v��(=��_l	���7׏GK�+�����G�}���
17܀]�?|��dJ8�7 ��������R�����Qx������1�9g��*�S�Ա�e�P0"o
>�CI/�g[���{]֍��,�<b����\}��@oޭUkM��f%5�!b�b��'�D� �x��d���n`���'p���4b��m�+�V�9�f-��ɤ�Y<�E� �V�9j4n��w���;���I�������ϥ���#&׉�m�ؘcG#�wlS�g��}�<N��3�f�`��?5�b}5\+���'_T'�$S&Kj@�èڰz��Pf�0X}�ۤ�	�LZ� *zD��Σ�_L���bi��MT}<��O�ܕ���+�΍����s}������)� ��cl!Gm�F!O!O/Ƃ�n_Vb�N۫��9��9�d��qW=�fL��v�b�^�#Q}�^�\(�x)��)���Ί��1.p�����48[ݯ��mXo�zN�5t}z\�' ~�V�|�Yb66uΛu��;]5,wV�̊����8��o.��vU����OO�c��T<��v�9�f窢�7����l��}��Ǘ��˕:�8�9u�r��R���Y�;u�p@ՌT���wbq��M�r۔��v�f��j������UU}M�>�Ι�
T�������,�`"�N�$�_=��t�B��f�e�,�!jlt�Z5QLs. �Z�/A�a%��ќ���v|�Ы��#N�p%�`�������+wAYmI�Gia�-�ن���)�c mL^��2��Qt�i<�{���Lo�ъ\1YTE�U�c�+���a��5��b��>�j�F�p�9�L��S�Ĕ��m�;P��}�V�G��$��xK�]�@|Ƙ���/2��te��in>�.f�R��F[\�@�0�Q���@�E�
���U[���X�l�=���o�9�����D=}qV��p�S����u���s��ǵ�� �I#TCH��٨8���ӫ�X@��f��'IJ��Z9�QS��2@�!�B��=.[\�efBYU۬�L��[�B@���r{
��S67����ظnc�19�d��V)>�)��_n�@/@����^l"���d��1���,ǈ�A���)��!�Ƥ�c$� ���U���T���n
��7j�*��oj^����E�η�f��cc�GgP�]M�N�)>Z���z,-e�PtZo�`r5��_j�b0E*�i��5����X�:ԩJ%ž�;�Ћ�#��t���U�02kf�����}UY���LnsU=6G���j�1q�� u'����=�e��Q"��vG@��ۮm�1Y�9.�wC����fL�7����&k��������
Ϩ.s*��5ښ���V��y�B*�5lh�4c>�t�br�X��f�9�]����({��^��lv~J�ߓ�M��cxGE�	"L���U�N��u��.#T���</�ʂ0����M琞7����ߔ�V�z�Lm�l�n�j�2t�鈘�}p�3̀C��n��[��R����(<ź9��^Lwq���1�~�8p����L��R��o㲀����<�`��Y�^u��B�9����ё���u��!LQ�ΰ���t���f������zά�쵈��b���]97���RSF��޴"YL���pk�� nT;S(,�9H	�i��$r/+����B��l4�Ha%�n��ݱ��L1���}�N�|o�Y\D����F}\�ִ�y��#����Egz�S���Tga���Z�ƹ�h�.�xo_\���Kr�@����U��^��]t��}8D�N98-�+t^W�����Ʈ����Oo7��m�Ϡ$6u��r�xO&ј��p�O����>^-�.`��l�5�\S]��<{���ݵ �P ^�j�#��{��=�(z���%�o۬>�o"��� <����w_f�IV�y�%����\vU��;j��=�#-/I��j݋jf�[��as{w�.���%��[͓�������!��o�P���B�Uo�|��D:�OMy[��(�p}PV�����8�0���J����#X�R'�dk��b���޲�CƖ篽$��T��	�J������:DN��@��ݑ��:��+LH:���;qE,�fyp����?T6�x̰9�
� nX�K���2=�\���s3��%qy1�ۭ��.�q��#�fmO�pʌ(0ECr���)��\Y�Lt�{�U"FAeʅ�/k��D\oڵ kDC�o�͘�_wM�\�V��&�m'T8E��'�0����y�(��f0B/�
^���L=��H�yʲ&=cuא��ի�����V��i�RS���Zi��b��"�$*<�`ӣ��u��*p���^������m���[-�\�o����7����S��s��.
6���:�5Q�Ɩ�Lz%�)�|Q���5��_�^�K{^A���%��cO4�ڎuc.U�W��Q���R
��mغY�ü�ߘ��zQ�27��?LǗ�z�;y^x�u��ς
S닊���2�{엂��h?Lln�2D��:�eЂr/���T�Te�!;�K|���š?}_}�}�S�qO4t;��#��y�ϥ�3��٧��pU����]��L�`��f
̍ۻ{Խ�{�cp��XV� +j���3���=F���F�ݹ>�YP�ȗ��,Ҽ���k�yl��4GIO�Lw�gamS>�cD0�Ễ�\KT�gҶ�K=f�ur����R� r�!YIt ݒ�;�:}�"㚧�E
K]�9Ie��!�"�m��7�;*��i#]���ӚV@85��%䴖q�@����&!����c^�4t=9W��5���GRc�z`B�v�@�:A��G�"o '��4�,�{C��Ff>�칗�-�|�b-�%fm�8��-��븛��J~B41w O�b\�����3su\h�l�o.�O����s1��h�j!7Z���E\A�� ..�g���kM��4��E��=��C�.�c~�KxTm��C&�m���f�0E�1�Jd��o�<N̬~��,�N��E"�ٔ	�\���LH�خ�Ǹ�w�z�TIJdɸM���"^Fe��we�k9�CO���;Z���5N�	�3m�e�E��<rӻD'����P6�s�\�ůf���W�=��h0�,UzO Y�l�)�W����L�O��nm�SFu�wZ�ޜE��J��q�D�Oo��[�Y��|��ֵ�V_nF.��}�G�-�I�� pЧ�Tūp��x�`=yK����HTv�{2jagܝܘ���6�[�6��ꚬ����5�K����v�֥4�@���鉟�,fK~4����ѳ�<=h][ٍ$(�v�쌈��*��_E7�W.�b�?d��ن;>U1�k3�]9䔑��m!��]C��+u����b��q�j�;J�Bp��Υ�3%��u:N��{˱O�%�1R['�� v>�:%UC !�Rs�ދ]�%�����2T�� Hq+����jaأʞ��V�_�:9�w�w�>1x_(�&������C�o�tz�b��SMb�����}�])��c��yL^���z�O���{>��	�l���X_@��W=<
#JX�ߢf���c^��*�"zV��'�^�僥n`3��U��ʂä� ��՗u/ZV\�{�;�I�~�����(),Xք�a�,�1��M۸qD������vZ��^��� j~�ٵ�y�
�f$��{]Sq�{uк�Ѭ��W����Iߠ ��MgG<
�x�|NWpF�<�!����N���w˨��2��%\Z�rL���+���ʈ�KMPu��H��I���f����vR$.N!�$�����>��һUz�s����.>��q�0�ثt#z�W0MrgK�kk[
*��)�����˔ ���w+���ْD.5������.�,��Nv�M��jf��t��*�9��>\��~��í,�~H�sVm�5�v��ڄ��9���Ч,
!f޼U���Z���h��9�"b:fI��z�`��B=����yӈ�O!ѓ&w�+z�HrL5�Yg!��k��P��Q1����[��+�nz�渙�N�Ƨ�U󅗼�B�v��.!5w"�&C�l�����A����Nڡz�Vd�Y�3�$bz�y%Zq�ۛH`�4X_$��br�X��fӘ�M�Q�����;����FW��D\a;�[P�o�:+�����7�m�� ;;	:�uPw���xC~�{�W����:;|��(9Dw��,�|V�*tzG��-3��+�`?EvH���1��Cv��Kw�/Z�����a^4٭
���Uwχ��J�ì�=�@V��q��b����5Cr��eݞ���B�!T��ԥ܋V�wOr��95v����Z5v�L�E�i0��=&K�}�R[^K�.L��}��3j����r�Ү�K����ai�����==�.��|�wZ>c�i�ˡs#*e����7f��xv$-\�uc3w5�{<�|R���S�Hn�Vf<bf�U���o0�u�J�S3v��78-g��+�����MFl���m{\̾�̉����&w��}q�iw�^���i��,ɛ}B'.�:#b��m
"�Ulw!�JP�Q޺��g�2p���<��q?����.�L} �M�Z��AC�S){�����ce�:m�;����TX��;�����ƪH>xE��P_oR�G~=��'t�y;5�^�e�`h��7��ʆ��z����T��ҹ̷Mp�7�������.+������L��61s��U�f[����l^l�����5Y�/27U����e��FP}�P��w0�����ִ�nL_f���O���$��+.*�o WD�N�e��)qN&����R�W�@u��|��m3�Y�d%���� Q�����J��Y-]��_������+*�~Xq>����gy�*�����WW^��~��, ��\�k�/��X��aD�b:M�W]D��#G#Ub���;�q�vq)�Y��s�OE ӁFĸ�87!���m{LQM>$5���ۭ/�ًC��3�^�HH��xg#��F�k垽��Eu\�-2��\��ga��]I)���q�byc1�9W)T�n�2��Oi�Ą}���*���GF��0�����Zwk0P���2���ێ��F���-j�|͉]~q��A�n�=\>�\�~��1ir������P0��x�����X���5����|���yù���E<y�ť{jY��bg��&�ɻ)�/����6ՏTW6b�G�H糽ʁ�܃�8p�:G=]�ls�c�32��{�P9���N6_7�m(x�su��s}7/�Ac��%瑰�8�8^�����/,gB���ה�o�V�+i<�|�b�_��]�����.�6�V���{=�L�����y8��ǲ��Yn=<��9|oI���%ZW.���sC�B]eZ���cDr��z1+�9x'u2��OzN���(�'L�:r8�u��{�̒޽����rU���n������f.��,ڴ��%r����ȷ7���c� �^׵��E�Ec�]�.6������so��1���u��tՂc5��Iu�T���y>���"�vnh��Mj�9g��9���n�� a�x7ڠ�z�\|��d�W��3���خ����)��;�+Z�ܨ�+���	�t�M��t��u퍹�e�ٝ�(_י��qT�s��̩,�Ɠ3h(N��{
��1.�"��օ����5����s�*/���j#����uv�9� �b�hP�L�1�U/u����A�DB$��djbfETR�D�ӐE�iI�&t��r�9�"D�j"EJ'B���rYhAFYa�'5���D�fb.\8P�)s�e֚�b�d��BVV�fYf"�$TGjJT���SVY��$�	D����9ȅ�uh�QZ���TFrD�$��ӖI\��L��IL���!�̄�IT5T�C5H̻T�E���BZ$*�',�T*L�-�H�,��ڔjȩs�W�Ԭ�
��l�J�r9�r�,�V�J ����Ι��R*%��U)V�E���ʐQE�Ej�KĎerR�+E"i Uf��*��\X��Qjs�]#h�Xh��l�3e��I̬,	D��R�jb�V�h�"�s���mMicY�V&Zl�S�Q��Ts2�D��M�sD��4�P�H����jR��HK��̴�QKV�ZY%�"��b���Q	,��!�E(Y�I�,�t�ǜ"�$(�4��L.���ͷn��^:sj�ܛ��4Z�`pc�IzU=��PV�����}(J��A�:;�2��X=[#7�E�Ҹ�w��ﾪ����q�]�L��	c�^��T<"�F��!#��X�$���zdkM�C�udժk�v�o\Ȋ����V���=�lD���s�s�1�F�jĠH����O#M�I���=�������i�Jˬ�#j!�P���[��-C�A�}N�|o蕕�d��#Ğ����ǯf�wɔ�������(���e�G����z_�b��C���_K���3�V��oI�i���K�<e$<��!<_���ToǙIL0���":ahMT.�e�ƙ��'�f�Pѽ���*�#6���<�ݏ������v|��f:y��Y���yY��ټ��N�>��D�û�h\)���v��f��)�3�A���1�nS��j�mD��\n�7�+�k��ot�@�"$j|����%�A�g�D�7�.uT彻���W)5�%�T¿�+#���?Sn����':�z�}���65�S=��0�^���<��ْn3^�ՠ���}�ѯ]m>ylgɪ�7�l�0�
hm�~8�Ol(�R�y��:Z�< Uӵ��!�R
�W��-��חS��R
����b�us��W;��ra��Lyφ�*J�D�L��^gK睮TV��5��kYI3W��,%Ж�����NT��xB��`=i��L-l=�����_}��WգO9@�S��r��s.G���B��u%9�Q���&������o^4�yKR���9�5(ox!�aaK�i�`>�50� �������A^�@��i�2�Ʌ�w9
Ey���Պ֍������$*�Ɲ�!�/@]%S�K��D -�ʝ�[���e(��������k+c�X��j0��L�F ̨�0��|P���97��s��Y2]^�%�iI�FmV���<�g�������s���9\-L�~��˙G��������y����g
�ދd�zIj'1_)j�1
�]p��u�Q�R7j0�������Kb�xϜ��V�Fu}Qc��P9[T��Ι7D0�ߍO
5���k^���u_ ���E	U�37wA�g�k��z���oI~;�6tc�/���Q{�ם�w'�s��5��q���ԅ�\��/�	`�}�(4��躅Kd���bXM�V�{��8�=�}��gU�P�7p,5��A_)X;���Lg��
��bmsY�[v�q0�w�#r��2�!۳W9"����9@75D�iҞ�z�b��}[�U�q:����#�LQ?x���u�yh��P��f��{�b �ё�z�(0|acw3	Ae�LM��ݛfܫ��G��zf�cѪ$Ơ����s:�{?W�}UU�b~b�?{�%3fy�Pw����o��Z����p�51T�w.�m��қ�ζr�I4������ا4�	,�[w��tmdr\�`�p%j����S�[�R�z|��;�r%�-D��V//U�P�.H�����{�u�z�_d�j��a�}F�L3%��Ms�ߝ���kc�9I�ꆽ�?V�?Z���pG�j�{�~=y�/j�ۭ�3����w��$	��gB5	�C���(��;q�j��{]y��i����U��ǝ�ٗjݷ/n18f��;p��5xr���}��gVd��Y/q��-4�w��z�d�EK�d���~�~E/{�q��_r�^zJ�*9��k+�\{Ss�)����⧽F�1<���LX�fT�>&t�{���Zҁ�m�`̨;r��gҡ�|1GP�ϛ
%���dT��]	��2k#�E�������~/����]H��:ܷ%˅�c{���DJj�X/��
U�pJe#EKiEp���-b���j�$@�-�F�R��r�iӆ����P�y*δ;bTBuJ�
�r؟V���a��ldaI��꯲E9{��'Z4������(�:m��C�߰y��*=��3����^+�bK�]h�H�<��{5�k���D��UM�-��Vl5�o�A�|�<�;䜴�����ՏCv��{P�{eg+��}���_�|kR�5jw�:(��oz��[6<߃ٱ�h�}�B��$w�2�|�#J���-<h�?F>�^�*C�]>�T�i��Gkb����TC�S��Ѽ'��9����n�i������m����K�il�6jRux.����
8�Yꭼ����i@#[�sL�1�=�A�Ϥ�w��[�k乤��"/d��2s3�wV���5�)�9����Jv�G����m��)�^��ˁYEn;:���=�.P,'�F�L;�\k�#'�k���E��"��׳�����6�^�RUK������Tj"ӆi��K{��xu�׾�T�b�SCX]Z���=0,���/ɧ�j�ɿ|��b�9�8�%���Jc��}1�Y:���2w��|���qHh}%wn71ǟL2� un���vE��Ŝb��eZ���\Ndc;S�m�6�k���1�pJť9<��˭q����꯫�17%.�N�d�_~�٥�����ᚋtΧ��4,�>S����5�r��:`�&�U�Z�*�g:�Ծ*^ZN5�987�j��2�������~lfQ}03D��}=ᝪ&ޱ�_ܑ
u���*��Y/z�VM^�}[�����lꯣ��{�U�y���`r��3U��M�����jl���kC"%��y�5<��!�6�І�A��AS�峠�݅	���᳽cy�Ȧ�>~O�9�G�b�\��L�3��2�+z���I�zճ�1��7j����񏢠�4�J���ڹQ��Rx�"���R���V�T�-O_�=^r�'�<0Fs,g�v*t�{z��� ���]�)����r�ƶ��4���9jy/��p$�1�e-�XS�w^ۑ^տ2i����u��\��#Q�F	<�:ҁ���Cur '�NP�ei<����	��č�
~�z�
��ͣs��c[�a�,�w�~�������W�h����F�ȟvm��;o�O��/2������U���a��2=1�H���}��}׽�n[Ir�^vz!>�OڇT�]Χ�b~X"�'��,�&�W����[����ѵ�W�2�6-����9�5�,���hR\a�Cz�1���J�$�{��OfM=�K��\�kB2�\+��銅L����NV�<�������A{�S�'�f�s�i�6���8l�#��<�-�H�hQkr*ف�����7�9�G���]k��[���I6�?-��P��^�g�_��]�V{�~���y�~����>�W#�S�=���8㷣U�z��7vo5���_t�W�:�^Պ�f4�s�-�p�È}��r�ZOZ�u�o���a˅�0*��Ku���J�
���{��N�t1Gc᧟63�x��[���=uc�sB��3���9�;�)ָt�_TNOT�}_qъ3�Zy�W�6�ԣ"�F��6<����`�]e̚^*�Xq��Ҕu�K�	�e�f��Ir5��=����Ty>�1����y������KSl��&_Q҆�oj�O��\��Tl���MY����Q��;zm�����nX�Sp6j�J�}7Fn�G�h����U�W�-�=����8W�@c��UD��*9T-��ᭊz�m>���ڌ���ۏ�ש
��oZ�.�+@Т�>U{�|���Z޹ړ��Gl�2�7�)�;M��4����Xt��$4��Kui�u�:��U�ۛ���NV�k���:���黁a��zJ�(�cr�\'�͵�E�r9�n�z�y��B�gC}����eJw|��r8K#6�R�T9�n�pX�b1*߸�[�}��o"�	����91p��#�j�o��xڽ��	F�<�k�[�zS[��\6�6-��1I�A�GL��{q��.�z�>��a�X�ڶd�sQ/�{Vos��5*ݰ��p�˞��7Y��\:�^��B�@~�٭���������]4w7�E��C}�(�����Zp�6�kF�"b5��sr�s*��F��-�`��ν���A�=���3)3ᥡ�U�G�u���!=ȱl����]ƕ/�k9ފx��W�/��t��Xq�w�J��W~IO�z�no���Ԕ3xۃTޚ��(���k����y,>���z�믬�(8�F���3�;7��$$D�q��������&��~s2i�����V���'�tη��^�c'�o����ʙ�tV������\�㯥����:���eK�i=k9����mD7�s�Va������S=/�gZ���{�8?[�)���#�8�[i=��QS�;�mciu��Q���ʼ�Π=��`�s�Úk%�ժ�7y4y�Z�Er�%��?)��gM��!�
m`���Q�~�U`������c��xp{�tj�4���௵vQ�l�N+����s��bf7yc�7�6�dףoiX�{.!�o/��Ci한�XK@�*�ڎ����$/=���X�}7ڧ�f̏-���C���؆�8'{3jǨur��X����}�򑺦v3S}�P��Z8�r�m���Ѥpu��q��	\�pr�H�_k���?�B}���bm����=ez/�ó�y���ˍ\��w��8���N���ox9��FN��*�� �8k������ue�i�V���-�oT�������聜
o��⶷X���P��X�f�}�?:�bp޷�ٺ��>}�7pB��	��{���>�3����&�Q�C�ɍ��R�ΐ�4}=��y����7�3�;;;� ��b���@���?����D�nk�Y�+��{7쏰ZՇކ����rpd���O���jq���N&:Q̀V��*����o5�
��Q�3Qo�f%=ۓW���r�i�5���͸�p��k�"y�5ZC�ɗn�>��KUr��;U;�Q+欬�I'[q��5��gS�OO)U���)7�eci@UX���1̵�q��'�Ź�~jOV���Q��٘���Ϋ�֣�o��7~9q�2��Fb���+����Q1X���KL�}Z��I�Ӡ��_9������"�Q��W~skv�1�2^��
|\�)���B�%�Qk�-5r�6�Oy��c�*�zz���p�N-���N����ڛ���b�=�1 ����W/�YYˬ�)yz���y-��:$�AJ�2�H�7j\�w�q7��ٝ7&*�A)Ymq�6TڼP8���T�t�!벲�=r��';�L���!�ʫ�毵rIʚ��7��̾XC�݅�ހ��[�>�O��wz[I��UUU�U�E�x��?X7_IݩQʢ�W�v�7��>���\�G���y�a��'������=tv�\�JD>[�SKS�����{�l(�a�kG>��0�pk�����'��Ё�#�r�LoH�9�V!��Y�o�����Gy����z����̧�x+�"�V�˸�'�ǁ��Ԕ�/5Uxqs��{���xι�9�1�.ʺ�O�3=T�85�-�t��rY��]P���$Ҹe�v�1I��sNj!g�.5�b���c�p�#]&���sbud�n�P���̶�5��adKt��X�Ogg-RWqH���{�Z6�NKy5ڶ��;��I�͸ֱج�O9����x���P֋��ۣU��~�ݹ;٧�o6*sڕ��h�}�éoOR�톅���u�� z�����`�PѨ���y��k����-���fs:n>��q��>�6F��;�;tW}���Ձ��$h�N��P����w�A�5�M��7O�����"��6ni�)��R����Zc�Ћ�;�S�{Hb1������ds]�T��u��+�`}X4-��m��*�ˣ4�>k�>kS:	4�ܵ3�8e�{���wL�M:U��3o멻�ʛ�=����Q��_P�$k�6#M)
���R�rѴ�Kܵժ=�5�G�s�6
� Z{��)茷�V����
���R���� t��ݵ�6!\k��fe����lG��[4|��^N�a�.�Ʒ[����f흜ŜE~���Ubd$kwq��&�,�j4�\=略���׽�c<I�-`f��ðb^�Bϲ��` 䫭�6.a�S6�+�8�V����.;���͓6�F�-��ղ�2�_U�:�T��S7�,��n�i�,��j����m�����\x`�]���ȃ*�J��XLݒ�����g*0�v��JrV�V�V2��m�!N)WJ��lj����Ge������u�Vv��%�WJ��3Uſ.b��ƻ�4��.��:U�&�Na\{�$Ѵ��\�o3��]s{�U�����V�o5�ṟ�V.�&�v��%�������^1%a��4!� ���=�y�YO��`�%�|tE4�K�*-���g}���=��j��LÕ�{��iX��,��Ώ�KQ���+�Z��}q��&���|�kbdwt��ƚte]<WS_Sy���MuST\�~��=V[3"�xE,�@��%�a��}Z�Z�w⋖� 0�W�u��Q���Ά�c��T�b4rG�\㑳o�Xy���Ą-iQ����u�}�*�}�P�2+1�<�q�����NP��Ӵ|C����jf��eeBu�'�&��w�Fۃ-&	�����`���'(�-+V��뻰�[M�|�����N��Y���W}�U�*Ǵ�n�A�t��ޖ�;i�ֺ�,G_i�Ra�#Xr��jm�J�ֱ)��b�RC�����h�����۲�3�J:�V��ii���:$b�t���4����n�nzg2G��6�b��_vjS#����v�{g���A�@�oEE� �{�Rva��vF5ɪf`ٽym��W�
e��M&앪W��fI� ��okbPݔ_Ti޵cS}���� �6^sP5@4M��ӱ7�XK�ɽmN԰��x�̝�5��t�[����M�MiE�O�nA��[F�To!�9+qV���1̊oa������B�"��ܑX��LU��z����ܷ���@�C�4n"q�v|���Ƣ�Na7��<���,-,q��ٱ�ůN���*Ӛ�q[�F����}��X���v7e�&�u6���u�f��_1�ȇ5�D9�}�Y^�8��J`>P�^����'�����.>uU��2���$��4�"	E
6&U��\%V�"Zi5��%(���:q:UUDD&EGS��]iIr�fu��*��b�GSB����i���$,��aE�Eb��ED�Ur(2i�a@VU�"Eh�DgB42��aUx��g,�	#�YUUD�m@Z�9��3���0,R��1R1��J��YbTR)Q�	LEH�����UIҰ�W:VQQC��\���Q����L�r�/������5�Qh�0����&��8D&.p�r�re
�eR���I�g<�i���h�IRS�(���E����T:�*�R5�9��(�DQQ�<u�W8���*�!:s�R�%3:&Е�,R��$QI���"q�B
"r��йAӑ��*�.Q\�YΑd�DU��3�P괗9!�L(��H$�
H��@$�F���E\��q�f6�I�Ñ0fJ�:�C���aNb:��=Zj,���6�*�cFή��gE�pr��a�Y� ����}�f^��Z�HQ���/n18�q�Y뇻U�7�r��������"m���o�����>�\ғ��vc�pT��OZ�u�o����q�����4h��}|�Ӷ�ҥT���h�ϛ/\6����Cէ���mi�D��ΰ���������OT�}P1�TQݭ9|����˾U�I��8�oR����X\��9�uT��*9--w�[Cv�[�[��l��� ��)���|&֫��BP�9�߳<��wvk�)�M�y=�ݼ���?Dʓ+=i��������h0W� 4�-�6'9�,�׌(��y�N2�f�������|/{�|2����1�那d s�-��g9���ҫ�b��=���\#��!��Qm���R��B�v��vJl��Ud�b�4�������[�xf�M&/[P����4�C�l���e�Q��o�+�T�����wK}r> 0F���r��T%�y�;+4�a��1ihIQ�/.�{�>X�}gn�w`�7~'0��,G�r\�7{F���K���4ӐNWB�m�"c�\E>'�]�q��M��?������uz�-��:���t��wP�K}5J�ˏ��Kxj\�6�>/$]Ъ�+��޴��KT^��ȝv�+g�]Ao<�}��/n=�ǲ�`���ȭ�ۮ�i M�Mƻ�,����skت����;c:�O˙�rR����Mc����p�6�m58�Q�LJ���؏M���{5?I���4yE��i"�8f��3���5xsX�Ә�v!Y�Jx���1�������ڮ��g�|T��ֳ��{�Rx���0k+Vk~D;��J�z���s�U������ҟy����j�1]2E�b��ޘ"�n�뼧�4�,�p����a�1]���yr���r����VO%�]��`u��M�N��_f�z����C�J��$�*�̵n���x(֫�m�o3�\�-�P�7�6�\K��_j�[ E�l-�Vj��|nv�tTm�:���2`m�ַdr����tu-���	׆��%m�6'���]��������.���{o�s[���Vs�Y]K/\�/:��,�w;v���,�eb����u--���/EL_>�E97'h��1�3>�t(�#�_W�_U^�^��S]D��J{�[�zǡ�6��Y�ń����N��1d76����K8�ٵ'��sP�<h5��8�7M��c/*�©F�zMSO���7�Rv���]��K�>�r���ۍ��࿲��S����Czg%B#���zL8KE���8����jZE���rC}۳YZ���o#U[he�����!q�h0y��Jח��ȸ7�
�tS��hs��j�|��g"b�(3�WW�l-r�fl�k.u��/��<�ڹMuKm�|����)&�\k��&���u��MҲ�G��2H_(��_�?��M^=��5'�8e7���q�b�ݪ.;��f�kVl,ꁖ�%fW���j΋ڵ$�n18f��;25�8;P�畯K�|��,�Cc��d�S}PѨ��tzn3ek���}O��η�5��Gvz�y�V0$�D��L��~p��k[�EBs��76���l���-4����)m���8�E���a��t�ג�u�����˲PG;���vܮgo�Rs/Z���5�%�܊9X�����E��.���}_T}z�-�����1V����������̣�nr�{�*;TrkOW�a�9�q꧗�Ѳ���qe<}����ާ��m`̨*��Ss����a�{׷�{�4��q�݉���A�͌�����}�i�=Vm��1]���y�_	��H����.���N��+�y��i��_6~��|T�8����^9=�V��(� �Ԃ���TK�T�z�4ކ��-r�⑽���}�|��tW$��n���l�.U%*�/��3��=���Kۗ�4��ȧm�]�{���p�-߫nJ�'�B|��_�e��5����G�
1�k��I����;�QY^>��׷R����a�	h�ϯ���s
,^K��S�y����+�Ŏ��uNj�]� �:=��uFl����9�7�N����xjM%���a7��i�9��%��I׷Z�����
˺WKՇ�2�3����-���i��-&�ݸ��p.gc��\6��]�6�Yg�$0(�8��ӹ�`���Yʜ��|{�t�,�WNͩ��	s�0�p�oQ�j����r�*��5!!��u �R�_��U��N�u�S�rW^�K�Aꚉ{�Q��.Cj9s4����q���Y��݅�*t���V���	�Ub:{~G�=ٿ5����=0:2z��O�������������D^z<����y�|�}q������ء�e���p�[�i�֐�6�[Ѝ[p53�>z��������;�9��Tެ�k�m�-y&4b9�T��\���@��-��Mt��|KE���殙8R>���>���pe=Q1X��/O(�[�������WV7���k�7]۝8���uM�W�����b�9�aD�}6����(yH��^�|�Mv�/t��!��6�B�YG�%C��(��֞DSME�u�D帬*���x��,�7�Եi������_I}Q*9TB-T@ƅ�YF�>�F��z�yHǧ��N{�|&֫��	B���o~�󝚝�o�:�ǐ�����<�4.�}t\@G�:~�l��ŗ�)9y:����.�e�J�rއS�v� *x{�e<ݮ{j�\�,��V�ob�ݬ:��LTS� C�9h܍�۾+9����ۨ⠫w錩��M�����wuZ��菢 �g縻�����Z�5k��6��X݋	h�APGp��]��%���(�3#-��ͧ��:{4�<�kZ������N��}�eJSe�����{�9�0����u��_OD9}�[��o�U�6�R�˘�{�����$�z��./�F�֊����4b�&���ky�;�������ӻ�Jm��u% �zӚd)��{���O��ne��:[�i.f�N�'�sMj�ۼ���6sC��*���6yd� ���}��/lE�ue��j�]ה3w�!N9Vn{䖍�0jq��ȝqQ<��ŵܕٕ��]4�T�Ke־S*�.���\rtj-8e�7�
#>�:-j�nU_)��\U���'��wmd�(�͊L���n��oj��Ð	��c=ۡ�.R8�C1T��X2�S��|T��<��԰�q��4��:��3�x�;�>��tȳ0��r`٭Q����̮��eON���<���R����-V%y�#�������{���W���p>�Ho�%�w�0�Э��b;�>��ͽA=�դH���V��m��*ƶ�_�UU}��P1�^���m�I�Uuj�U��S�럻���T�e���4�}���4iQ.I����s�j��e�y�@z; њŖ*)����\��۬֔ц�5���W�6�S|��i��C�aM�{�_����&�o4��l�\lT-嶟\K��s���w��=7#��42Ba{�����)8���Z�c[ǡ�_=i����v�bcl�M�f��;[��}�{Q%��ڒ�yJ)ۆ�[p�=�y�2�Q��j��|�(y-��\�PBQ!���K�S�e�r8�q��/�FJ�u�v'ݨ�I��R�SP�S�}�&��W�s̖#؛c1xvx���2 �U���9N!����_:�5�?t��4�>���k��_'C_U��k�v�KV=�iS��6�>i���q�q�*oO8�Ɍ[�㙹�p�i�yfx�k�V4�/��^�����z��&><�q�EN���!ٝ�jVv�@��w����|�_S[����TyVj�*�2
]�CK�M��K��3�v�8{$Y�S�� PU�#��
ռ� ���-�ќ''t�?}U�U�~T�1�LƳ�Տ�7�ͨ��jy�ڒz�k�Լj�VOV���ĥ�b*�\WsK��9n�/s/��x�{�;��N�q��Fng���`:�φ��/��\G�ꂛO9�o.?k���mZ�I��p��怮�6��,��z�va����f��؁o�b���+T^s���빆�����ىyz���J\c����=�g/��P}�3M�T��:���^>u�������0���<�'iI����wju�mr��;Y�����Wr�Um���n5�����|��k��y�3���S�Ͷ����1�=��)�u�!���9=Q.F�����o���?3T'>��I��(�m �&�t�Qފ'�Y��f�k�ћ�������7��>�xw��r�N��ƓU:�!\��{9E�����ʤ�R_+W��m�^���Y��7p��� '�]me�JE���zHeo�ʌ�-��g���]<�r�E��:]8�x9X�t�:��ы/��� B�e�t����6f�<!�fmLM�ӕ��ގ�)����O�V%H�Qus�6An4jT�Ŗ���h�	˺���}˜�L;Ɣ��C඾y�o��������*�#4�����Ɵ��)7�ݩ{8��k��le:���?w��}-p��ᮄ�-v
;˒9�nޯ���rҶs^�}��9�:�5�!O|�P�9"І���Z�Z�q4�j"q,�--ᚓJ�|��Rob�ӚbvӀ�?C&���w�+���rR�"�"9Ԕ�B�6��3M��q�����1M*6�iI����j���������G���j%<�՛�����Y� .X��Z�9*��[͍뀧+\Y�g���v�'�ˏ֜rx��FgL��g:d\��q8����jr/�Tk"�T�U��y�6����P�/I��q3�ǴV�jL�?t�/�x3]�U�S����{�c�`㙻�6[{�mk�^:�x2�\V>}K�i=k9���>�{vmO0����fg�La�������R�ø|V�xg@dX_a��o�*���a)0��{��/���W�K�~5��s}O�����K6��>�d�d�KL�:؄�Oxk}j[�F�������� �����)��b@zc��)�����(��+#�L�S�Pg*ܛ�:�SQOb�Py�c%����\T7�u�,���Չ%q�-.hu�Z�k)���,ֆ3/���NT���y'�y��0I=�%��O�yN�t#ʰ��>���Cҷ�!ם�EhT�O�f�J��p�r˄����+:�]�TV��T�T��u��Ӵ�5��xҚɧ����j{p�5�����OB���aJ�:`�K�*�"�ܫv��׏�����͸WET*[(�{k]�>�8�Bt�P}t..�8k�h����.k�u��dW�-W�u-}4��Z8�r�m�7��g���|�ϗ�.4��_wO�%���w�u-ᴓJ��l�n.�Q�w���f<��mbQ����بSJj
c�.�}7�2��KxjS[����f���JI Nl���N��l��n�[|�>�|˭ ����
�z�ׯh�28t���EV٢��d���#d��m��*N27hɆ����j���݊́�82�×mvr��g*�����H�Ïf�]5N��R�͗��Y�$�Š�K�*�8��c{2���h9uPt�v����ŷ�<ޫ١w�L��U�ّ�VVS�΅�E򻣲�0�t�Z�[�+�nv��Y<>�AMd�u>�4�����p�c;�����ݽ��M֋��/4T=WԚrჹ�N"^v�����.pη��~��H��h�-�bw]!5W%��<ۢ���6�˕c���6���Ħg^��S7��C��k��������H��x������ �ETmp~�E���:�v�+���Md	���;�ozU��U��RVd�%YA�z����=t[C�2�C��oH�^W7���/V���]s'$y*7v�c*�,֝%'��i@K<V�n��`��U>�9�e)��ܮ��d]V���G�����a�Qql����zC:m���@K/�Ja�rŗ�����H�F�.j�N�$��\]u�wZ�VĨ6i�2��x��'N�_,KfM����r"�<�.��*F$;Z�^gc�Y1ow��t���A��-��򧽾�N=Jc3�k����\)#�A���G�&UZ���������㡶��F����b��V����N���mhB���
]���;^2�+�f�%yA�ٓU�9��$��\�y%Pa�[���;�ö-;ַ�_Ze-&�wvl1d��(�EߎAO9�(3��Su��)g8Z��[��I�]��׳�?6;�dFw*2�e�.�Eb��r�)�WGy��k��D@�f���ھ��n��sm\-9\˶�D}��Y�å�P�n�̡���Sj�Pg�^i6��C���YrQS8�GU�xY�nok�˝�>�t6��<\��H=�l��R2��{:L�q����x��vf���Z[s>銓a�93��� Sl�(��c�]��SIe�K� �x��2��z,n�����R��Ki�YD�rYq����Չ�8�����]��Ç��r���V�bn����$Jd:esƹ��N)���B���q�Y�oe �L]�b�k�0�i�b.0���-�i�);O�q��l�%��{�w(��a�V9��̨�X5�A���y�tK.�+N[�Е��G+�� �X��y�0���!J�j<��)K�>r�'���1g�K�H�_����:/g���H��J���Ђ\�=��l�\��˝�3�-��h?H���܊u^mei�`�ͱud�ƒ�i��Ws)�JZr+� ��̏!o�ys^���%�;��ǳu����<�� ��x^A'`f�r�^�-v��]po3;;�`��͘%�1{��c����>#6b!��o�J�#�$���%b�:],4"4C�Zh��Fg"+��9T˲��.QE�R"UU����5
�dI��t���+BΆ��
#�үW*�(�I
�YVK"#Vq2���Er�fs:��՗J��Q�'j�G"̂�QD]2��U���+0е(�@�#��@QH���J���+��*<�8���ҊN%�b�.f@,�'"�dAI��G*�9�UEF���E2�r���(*�I�Is�(�*쬒,�hh�"
5L�9UGr��*&\�����N��T' �D��!a&���.Ur��iF�K*�8kU"β֕UQΨjȹPQ2��ˑ&	9� ����!��r6�m�㿮�t�T	�O1w�rG�,K�n�i�\�;�_2�S�YX�uF���{�����
��e�2��{?����8�	��d��[ڏ��BI���|DƸ��Cf-���W��lJ��_����[�f%=�c]��ou[����Zp�6�kF��&5�ёڶg:�Dʹ��*��W!�l=G��V=��[{4�����5靸oj��}]��6Z�~}�(>10����מ���j{h�~"g��I���}��]ӷ���+P܋��6Z�9�V��U��`r�����[m�S6{���T8�j���~O�HJu�\����=��*C���nj��J���1�,���62Zj�_f�7�����c�*�P#�ҋ�	Py�ҵ�nz�S�A�r�bB�������Ϭ��]�TV���*?X���V#��c-ɏ=`�iu}�9\+T� kyoCyp�=��ۂ��� 2²�耎f��y���(��hND$F���5
S�������	U�טt��|��ǃ�*�|=��ڶ-չ(���:|L�K'<�h��c�nN\p�U�	�p�BAÕ?��ɈZ#� {�I��Q#��vZL���Jo�M�U�WQc=A�Q��. ���f\���k2b0Ҿ�:�sitc��UM�;�ˋ���>���A���
�����].R�z��9�Bչy�=�����܎�g7�:�����!w���%��'��w�ٍ���QL�v���mD�[�֮>g5��w|�N��|�S�T��|Y�2+Ѕ9�s�'�n��|�#]8�e�{�i.j�|�8�b�>N��"�ԇF�/�f[�W�>�j�pud��ɨ�n� ����I��q��ȟ�8���/�\Xy���'O�z�t�����qQ趩�w�&��֜3_6�Y#��q{.6J���)޾P3�Ő�0-�@�E��{f�Vl_I�I��V�N��}����ϼ�N���������^��n��1�y�2��wՒUk�x�B�S���v�����f��eA�L�Q78;�nf�F�J]��):1��+0��e<|�������kgUF.�ث?.�Du'��18:�Xq�KY��ov�!��&��I3�O�YQ}�Zs�"�[�k�b~����2�8��0Bo �k*��w������}����¶b���]];��j�<+k�~�/,P��1���okL��o��.��� �f��V͝�'$����m�{��8�g�+��]P1D�.y�c"Zh������=�ķ��h�:��n!غB�_�T7n'��T.�/����(���|���p�zk58�5��k��v�ʜ��C��Tr���wCy���Y���h����?o),)Mz�{�6ng����8pH/�*�f���U��EOz.<�%xq7�=������[p^7b��_7u�ͅ\��Hnw�ϭRm'�ϖ�MB�ؖ5��lc�K`X]��A��������S�9&w��MA�>�ZI�׹��x�ӪsP�M�I��SqS
��n���iDbvf�Kח�*[�k�W���!�b�M�����'z�\��|t�#�4Yz䭹�M.Cj9s4���E��%��qu5˝jJҌQ��ȘjЯ�3� ���X[���MGl��/|ނH��M��;��k/��2�&kp��=�+]>����u����r����.�Uŗ�(4�{�e����A�G/�Աr��F��Z���_f�p��ٶ�d���J��b�w������n��+�Z������R��*�H�l��ڶ&��n�����r�-��4}�ā��k�o5�徳ߏ���ݹ;�K�O�Cv{�5�[ם�w3f\-���'[F'�[p53�>z�X��3y`�F����$�55��[�勫�w�jҗ��k�r�\cڦ�kg�\q}�uۛqx�uoc��w�7�R�ev���|�x.z�}η���d�����T#�eoZP3O?�`Uas��ʔ�TQظi�͂����]e?Ɲy{����a���U�=ZrDI�;
������W�ѸS��~�si�-5�d����zl��z�Zt#�P��ܔ���oVe�
g�:�~缎�s���=��i�i�|Vu.ª)]��J~pcw��`#�����&oS��{p���B����k.���z���t1Yp�m�2�*�S�K�ʃ�o���T�lҔ��k���y�Ӗ�R�4�*�����sz�4F5eԎv���Ҧ��A�ú�O�'#a<��
bt�#�R�/��s�|��*�ݧ{���W�u��r����I��o���[��񙢜��*+Z[�n�\�[�GZ՗+e+n���I�ܬ<�Q��f��������ü�MRO��5�h���j$s��wB��N_u�8�q��gf�Qٍ+��K[�@��f�:{��:�������Է��$��R|9��=���~���^�yS2��]�@O��neƔ����:e.�%��K6���j&�?�5�m�v�1�5Pczx���V�x���w�k[ݬǈWn�'�\6��|�O��$�5���|�w��=�k���u�aF�.V��8qx'�q��OE��{�=^5�MNS�d$��cC��fη� U�}�n���꧳r�⊤�j�=^5��gF��$�F�y��ʽi@�]Vm��ȵ�1T��X2�;S���wK�/�����a�	���k�W&��Ks}�s��+��2�[���|]����yY:�^Z捕NN���x�>o7�ϼ�#����ʿ[5WK�b���B�o�H��J�W���{纐t�� �8<t�G]�������6x�m�s3��is�89 b��v�W�vt�4ݭhM���z�l֩�l�z�n�~��h��t�w��㾜�/Q�Ţ%�{���FT��%Ƨﾃ�Ϡ�\қ��}v@������C����W�A��m�r�������Yڹv�8�6�vW���1!P�7�����g.���$_m[w�k[��z���k�]R{�&_%JTcvކ��yͧ�Ň��;3-u}w]s/^��>]�ۊ�hb�*��I�v�dҔ���o�	
b��u{�:�k���$9P�7B�zJ�/�]�t��S�1٩ig���{ڇ8ށ����(��`�،p+�[j2�ܞq�xg*�9�ɮ5�y���֥���J�	��_:������*����˨��+2:BK9%7�\�v0���.i����q�p�D�v�E�O#�m�fs�{m�<�H��!gK��=���'�RL5��adc7�(� ���䀎�ZT��K�ˉO&��sƚ���2��{�����=�6pK��٘@�hÜ8ca�fң�S0i�&�h��ō
Vs�j���s��t���fs�5�K��t�J�mR�*���ȷFr�u�%l��(R������*Q*^�4��Q:�GMR��9�63f���k�o����Ku{oZ����<y�{8J/٧�����}Uk��v�lú u�$�)fOC5v�$��oB5n�ۄ���f��߅����m�X,q��&��;޽E=��h�[I�r��q���,���۞�3{�/����1\��[��G���Г=!I��u��JϷ��j��qpS���oC�ꇹ�U����Z>Q���Z\;i. ��9���|1��ظT|��i���ٷ�������k�7�]�
�"Nl,��U�>yz7 o�$)o7�M4�
��Kn��]X�1{�ܶ��U�Ͼ�n��Y)Ȅ�[�Y��4a�ܚ�Ԧ���Ժ��_.�aJ�6J��|�JD>WR�r�TK�fN��Ÿ����kuk��/���9hv�
a}�T�(V�|P��t���E���Fsmú޸t�i��K���_[c)�%
c��О���7�c2�%����޹���R57�n,��F�B�TXGZ��,؛�k/�·���R��-�1�����>L��0��x1�1�"٘��&�:����0s��	]��O6�=B�@�O]n$��(�����%7�^/;W�&Cc���T��cu��>��)��#��k �Z�CR��k��!�׸�hx�9�%>P�]Z�����6�R:&��b4�kd�w�r[�Ri0�'��\ �\���}2�RP�sNX��7J��/f�]�T���r�ӏ����7�+Ww-��k�SgcZ�v�B�z/Ξ��Eٿd�f�Q;x�f�B��*�׫R�z�vK��-���NWѮ,��:`Zڀ���e�`�]�u��7��u��Ku>�������շ��5m�ڄ�)�Uk?]Tk�3�"�}�s�X���މI�7�x�L�[�*����q���=�%��y�����[}����+�)#S;�3M����+�Ec��T�Ryzu|���c�Z������Ƶ�.��˛-}o><�tv����U�9>lU���V���xs\�#�����sm�\O|������3U�ǿd�:�Se�mވ�b�bC8���%t��r���N��Pwv%:l�/&��]�c��x�U~�_0:̑.k���yt���I�t�+��������2�l�{�-�Q�ǐ&w@�8BN�:���^��f̡]z�:7N�2�Π�#��ͬή����U��w����хW���M5q/�n�P�i����:J��K��;�6D���t��I�/vw�kb��oOT����]�n���Tͭ�W=�S�R�;q2�X�g��V�ik{o�YoC�����n��ሐyl;��.5��*@�#[펺.�-�S����ϟ�y�"�&vE2�d^����X��}�`�!(��?<,G��o�͚����ƽ7Mv��R�'������\3�q	1�T� ���*�®E{W�b=�'j��k�˭n`�me9k��?��O��ا4��bvP�L�^U�o�%I �܃ž��o3J�-ѵ	�-�3�;G"S>��|�b=��x��Oc髳�I�Jg�N]����w �>��`�n5���/V�S����2g"֥<��k�*e�aN�~�[]�j�:6�3�6�kF�g��{qڈ��yX}~���t���.{� 9�Q�:
�%u�@`�+8uylId.���&#@LY�9��Aw��hK65@jj�u�"��c)ԇ�v�]�/Wol�Ѩ��gur��@�s&%r�tL[�%B�P�%u�[��Z��m��UU@��=�����S]�>��\~ױ㼒��n'��I���e[����^��ufK��\k0-�@�Uo�%`���ֿz�

�vk��ػ<��hο|�^���{�_7�r�eAW!⩹��w2��Ъ�M(w���:a���<�x�!�L�'�G�3��D5i��m^�K�t*���V�+�O��Cuq1����KM\�Ͷ�W�V�������Y�__Z�/�]�D���\>�/�bB�hoOKլ�몓vw\���.z�rN �k�yԞ�|�Z�p5�������h�[�m���^r���/G��A��r��*ʾ��D��j�M|�<�_#"�o� }�u�����[P�7-�

a}�%|�Piu�].�r �D��h��j*�^�4ž�lgT<g+�U/*;��^�hUK1+��;8s�ݍu�6�<�}�
�_����w�k�+lo$�5�:%u���!%��cŊ�1��_���6*�gyj;�y��+����C; ��� ���#y	g+s#�!�׵�A��c�	G�Nζ v*ݩ��u�f��d����O^��jG[�09V��Ʌ��!OEt����c�V�i��P)�Y��3��D�Sz��JT.v��Ά�n���'G�)_)�����G�,�Yk��x ��t�(Ь��U�*VE����X��u�@e	`<M��nͼ���=9���x9����q	���q��7��k��|s�F�.1�]/��A�\���`h ��8�b�[��`ku.��o"�����Է2����ҩ]��d͊�q��@�*�C��z��`��wn]�մ�]���f���,��g���<�#+�8���o.��$�e�#��ج&����xZmXhL�/C����\����0=�XSF����8����_UG��Y$�mѾva�p�*�Z/hps]����AN�i��Yc��=z7ޛ7J�j�Q켝�'*�k�)Y�,��\��8	3�F&��7���m۵�Ю��i�Q�/�=V�5[�P�5�dw��t\@��D�Z˅�C��w�Y�5���U��Z�)M#��װ=Xb��=+]�p��_�@�]�~>�r�у(a��e#x��'eo)[ZT�6m"�V��]�K��cX���^R�T��Yl�xJ��O��$%l!�."�,[;�c���w.���{ׂ[�!H�+���a)8_n�+���gǮ���E���+��7]��C�{�y��[�@[M��vC:-�lE���V:S43��q��R��;Ѥ�p����������b���e8������@��4qDF�S�EG��*žn��נ�ܒMxޅ^w��m�� �]�:�32뷹^�����u��&SRLC�Ӭ��PX\�� �y �7��^�u���cC��;l����B.��6m�u�%�9�:��kEY��̫��t
�*�\E�ޛ��G0�|�Q�{����MڙLyXVm,��íQ&�1wr�x*�֥j�1����]whL�:�+�O�֐��i\]�9YubI����wb������ �2kͪ}�h-{�k|����V<�#����U�].�W�s�Bs��L����R.'_^���Lӎ��6�щ�N���F����m�D��u8oV�k��FDj�L���Ӭ-y}�r��o����5���W8Dh��;�H�
��q��A\�i(r;�Y��Wd�b����Uz��L�Gr���0����ttMl�[Mk��m�[e�V8��5�Ïn�np��s393�i�8v�d-e��R�F�Q�|W�͚�Lʽ6��h݆����+������0,�4l�����Y`d�ٻy&��O��W�8�5��SK��+/D��N S\?<���~����"dDA�"��s#��QQ�M�s�
+�Qh��8h�"�WQ�J�2��
�Ar(8Qʪ�T\��B9Tf3R#��*�S(�0�q
���82�eD��\ ��.T�9vAeC�L����TPQs0�����E����ܡ�UTQUUUʈ(���P��T�R�҉��
�"(�*"���ys���VW+[I��TR��UvD�(#�*r�*��R��UUB�*�$��Fk�((�(�S���(:q�4"�QU�u��(�E2�Ȩ�r�r� ^M'M�u�^�(�n�r���+�Dh�É��ܩW��9��	ʢ�.�TQy�QD�Sk�sR;(��e��9�EJ��+S$��������� ��D�r㸧�yip��7S=u��:�dgGs���vD��c��C�K�h���o���6��h���]����k��0�!t�Gϊ��v�{�P�`�,x���
��-�V����
�����ZJ!�֘��N��qf@TU/������ݑ꣑^U��$��sV��ض3�0��gb�02������ӗUR%,4"�#9���p>�>��a��q���]��4�s�ݧ77��_n�c 1�bՃ�G��m�Hz��gk��TD���d�
���j�jᵛ�е�B���P/���q��;q�S���'{�r�hsI�1k�;���ﻺ���j"�3��{U7Q�t�-�f-�ys�{1}!Ŗ�Zw<�IB�MU�s����]��Y������^c���Dz�u�\����R�˩Le}��k;�����7[��z��[������Os�o�3�Or�܀����])����ldKMט3Vj���Y�ì���s��V�oD5j�=�Q��y���/~��ʮ��O�O�%=楜{���cx`��AʃB����mݱ}��+b�u\��␆��kGK;e�B���1�c:f�,G���"��]w-�]�(���u�q�Ӝq�v�Ƴ����*��F�R23v�Xr�K��m)S�A�3����ba&C[LU�W����"�$�ě����]��V��TrZR��*a7U���y���4�|�'��>�i�����+@ق��|�$�Z�̑����z�|��x�R+si��C�ֽ;眴;n($�ޒ�d*�����'��Z������m�5t�ç�P��ZZ�d>���2��%p,!IWAac���r�/
���W�W#%���͚rҶs^�7�)�;�sUr����v�/��v�<���7�t�[�7��X�'}�4�|���Q�1gݫOZĢ��7�JiM"�����Z�nN�|�+�GR�Dq̾J��Ip�X�6xWf�wO��,��K�ۧ{��)����L�l��⩜�7Ѯfzhғ�q��)��G!�-mn7rw76'�q�7G����Տ�m�i�>.z���j"ہ��s����c�ӑ�z3�l�]6�ng/9�5N�y�&��=� ��;V�G�Cg����C�.��
��v��wCE��&�P߻s<G)I��ey�٠E�L�:w���*����]�ԏno�!{H�H_R��:2%`n=Up>�	��n�ʛ\�g$���%\�ǲKkjs�g��~��{4�){bq���=x��O.��k$z䒃�=���|gXngֽ�0�l����ʗ�'����H�
�4�ܗ��*5�+R�|��+��k��be{�U�yW<:�b���P�ފ׶��U�t��Q�v8�꞉�s~Qt��}a=��=��EHα1�]`��T]mj֎���%���E4���ۆ�W��i��;`����͢��N)s�;�yë}��{)\lS�����{��VEy�ydZ����5ă�uNpQ������U�5>�=�/���%�<�Պ}��м����u��G�Au�1��_z���S>[��&���7�F�I`� �H���]D�����V���+|��K��]�##]v���͓ϗ#>BQ�G���d��C"*�0�In���ҼUb5��W~�,Ce��{wx�߯��gs;^�+��Hq7�{�G\G�튷2\� ����?끰_f|�CFc�	��
��^X_g������.fЭIV����V��9�<İֽg�:���̝0|����3U�}W�6�L)_)�g7����g��Z��j���s68�,�y�t�����77,�K�d���T�����ג��V<�3�%�EX��g�8�t3P�sޖ�.rVm��Io���11��OV����:#�W�W�%��T���=$LK�!Z�nL?S�7�ב��3`�|���C}�>f��Tu���}��O�����c5�S�g�ϥO�k��غ��^���N(�[�j��:V��.�q�K�G��ܘ�߬�~>��PF�zEG^܊�&Ю�uj.e/r���أ��b�-�^�i���c�!+�g���E��L߽> ��q��7.��u��ׯ���l\�>���Q&=�wL;�V���si�:��ng�_�_aB�̵��7���cL��;>�O���y�܍Ο�0y��P��QzN��t�ӭ8�ʡ+�go;���v=;U�'���>��Y����#/�����G�����+��
"F�u���vO�$����O@��W,��}/վ+�ʍ�
��D=�l��{'N�L���{��l�y�>�˻�+�.�����F���z׏�دS�y^W��k0�����vg�`�{/�l�_�C�Uz�ʀe$��Ӑʱ�C�5�(|=^��?�^�<���1��[@�߂V�V,2����̷y�P�\��ü=`7D37-w�48`}�:-'Ie-���θ*�[��X;ٲ���wn�kΟ`!���ձh-��p�[X.[\��H!o���d;`�d�?z:��
ۅ߮�O��W�wݺ��Wo:\gis��%S��r@�q�F���vx��f �c"�R7S���t!����Ͻ�}㾎�Οz�葵��w#�Ԅ����h>9>�A��,�3Ĕ8|��l�L��]���n=�&}���^��<�ϵ���;��Q�q�U#}� l�P��j$�$7P(z[*�ZQ�����c���v�5�����[�ZG"���;�IҮ=��~��j��,����9�"���i=r;{;�M�>�V�3<g���H,�^��gޝ��;��{I�~������иs%��ٕu.Sw���*sJ3�V��
����)�u��@�7�Dk���1��G��g|K�����畝o��������uz+�#=%�BZ'��D���n�[5k��[N�𿟕܋m׉�n;�eg�z��޾{]�ҍh����^��
��z���eEDK��9E��^m�◲�3;{�j:������*r�$	��Y��?_���hm��.A�>%P8;8�W�t�z}��&�çӆzs2{;��M|��㱿]��~�=&��^��t:<���\t�h��+:=���0���#p͞�WN���b�\A�V#U�>˚�)�q�q��u���KJW��b`�v��.ef��|9���͍f�|Q쵠y�\1(���ך]K2�^�I�X&�z�O�t8%�b���fb诮�r���@0oD�4�s��S�j��߷���͖��Z�y.k�c!�Ew�o��%d~�}�����ӟC?���+�����J��=�������N'$��r���S���#�"]/d�_�|VǽV9yV��"}�PY�w+�~Ԕ�NF�'v��ʁ)�ɭ2�]i������e�e������<����%�y+�g�^�G����������; ���U#t���C�F�D+�ޭ��=08�����joݎs���y�C�g���k&GQ�N���hʨwF|��27�"�5���߆���y��XP�U�����B}>��^R���<	=Q2���P�wMP���^��ϱ.���?�:c��9_���hW|�߸�G���#�'Ǯ=����珠X,��9fO��ͽ��d�>t����K� z���R�,���Dz�HU��hhϛ�[G~�\g�pv�wl×bQ�o�Mܵ�5K�!���A�A�:`>� ^S}�2·޴ȏW����޿�����q�E��dMLT�<�+���>�]��<d�H�U@�%z���|}��Cw��poΘ?DLڭ�UT'/»{��ԡݙ��7�Y�Cu��ƃn�1�/�i$��g��'�c;{뽣����)C ���Υw�G������0,زjX[��ݮK&]��S��SB)0�8�XJpřeS�lr6p�]�+�$�i���ә��&�84�y����_�*�s>��d���� ��QȢ��_���������ҳ��lz����n=�R��^ w���+���,צP�3�n ��R��Ub�O{��w3���S�f��ޟq�yP�Wro����� o�T6��2d�)�T��;�_�����wln,|�}��ꗧE�Ki���|n��y	��f�EzNx�~����=^�1��>'ĎЕ_�P�ϕ�����5F·�T�:%�'7��Cםw�����dg��C�9�U}��P����>�Z���1�Ǜs�����a�;���ODS�o���{�~.�z	� i����h�����a�cd~�ؼ�m0j;��Յ%�j"�>쨫f�������2%u��^^���d{�ݮ�^��)Ͻ�\B�Z�]%Q�P��e�=P���R>��x�n{<��$^@�>�����@�KԼ}[~�~/+��{�m�s��H�Q,s���q~��V���;�=�Wo�/EL�/����3���W��ui������;�,��F�Ze���r����V����KkF!�f����ʹ�<:�[�Pe��l= �YaP�]����(�V�:ӏ1嘺.U�mò�Y	��|�n';r�[xٕaGp�����(���mtI��#����=#jy,���RxGfP7z�3���<z�p��5-�����/���$�Cj���C�V)���B��7=�|z��w�6S�i߳��\�Y仐�1���t�3ğW�X$Y���]D�ݼ�B��������*j����/�N������[,�Ct��~�\{I�DTf	��@Wǥx��j/��+��:��e�;���䔓����s=�ԇ������)���S_<fu��@/����i�=~�諚q�O�n�׼�z2ϗp���m��}����h7������xֹ�X��IjnI��ޥk�f������T�:7#�S6�
�����M���O�G�w�����<H�y>�7�mz���=[n�����!>��@�`���4/�r���z{�Dzߕܘm������{"�؝�𘸫�>Z}�Uꎉ}� <�u�Iv.a��Xb�|��dS�i��c{��0���[�2VrIz�'�U��O-�j;�^�dV��R}��U&7�
��ڐ:<��ɟ[�U�����r�q/z�o����B��O�*��ǧ�>���\y�܍Ο�"7f�����c�P�?��-�J��p�6tu9�z;��Pi�Uw]x�W��{�5�K��~��¿9W]B[A�\�L�r��M�-�r�[��;�T��8i*:x`X�t�J� S���l���g�Kġ�q�5����+ݒ��1�l�a�`183��7��?W�]�L�	��ü�az�
��np�{kd�B�N�����~ԕ@j���ۜ�c��ҽ�#�=����p+�Wϥ�/2_�|V��q�o�����N�y�V+��=���1^�3஧h踯H�;>_�]������Ez��ȯ+������\Zq��W��J�q�y��IV;�G﨎��(e|�b�|��\6hyg�]�E��������wdcݐ�^[�S�R�����0�L��g�<?�*��R;U>	�ǖ!��z�s�>Nd���������%:=L��#��?[�K�A��,�ĕ�a���P�"��d�����N�������1�ws5�|�m��zO��G����j��Uxy@6K� RC�C��)3�<����Y�sCx���qW�ZE��+J���W�\��][5p�Af�AT��uK�eTd�mb�kY�'�=X�����3�m�:��c>��_����i7?z���z��h_�;�����i:&���eI�Iy���)�x�|��;��:�W��}��������4\���%�N=r�[ufe��K�Ȅ+�Gf�-���ؐ���{��ځ���5���jZ{J��zS�����'�`E
������.+�'�F՘jW;���S�]�	tα�ԫ�H�j�`�lT����T]ka}�J�<��0�vʺ6y�s�R@z:��z�<eI�2G��'��K����[5.�<Ӣ<򻐜O�3)�ߡy��}�s���Q6��5z��)�.�R�rz�����TTD��Ӕ_��mCӎ+Cwtf}d/��Q5�c����1���߽~���ދ�aO�T���ο���.��B�2_��8�9��o���n#:���~�㑯���|'z�,\y�ɜ����A��R؞b&��m���[����Ѳ^���Wѝj�乯i���Ew�F���V����Ӟ3���B���Yد'���O���}3�T�
�r��G�殦�ǂ�]/d��_�U���rP�V����ο�1��������ceO���Iݳ1�*�E��:v���,��� �/_���1ϊ�krWq�]~J��.vtf�'ԅǹ��9p����Qz��W���rQ�#�Jw+����P�O�h�'&h��_�?{��c�+և�/)�25\�'�I^5UC�|�O�;�:�욚
9�I�&����,��q>>���9�W�x"�p,���OTL��ձYQ9���\ኔ�,��W�w(��=������{z�L�
�K3���9Ha4Slv�.�=P�Bv����ڢ�L-�F;Pi	�]�)�ZV�&�B�JED�v����Tח���+�ۄ�/V�����,n�3�x�����/o;X���${�mĕ�ޏ�mHz!�^v^�7*+�7Uu6�o��~s;!�fR(�f�����-ƃ��-���ѓ�Y�f�Q�D�y��n��K����5��2�8h��ߒ#(��;��)dgq01}X���)�9�'�]�s� ��D�ٸ%Ëyk��|�GZcvR�4Lt$��P�H��oh$���:���vd)f{@���#tz0+���X�ɱ�u1�aMa:�l��
�su)˷��s���Sb��Te[H��Zy��d=ޥ��!P.";=�es538R5��^vc��0�x�6�0v��5�o�%-�;�i2�vg	�E#ɫ��]u�:+#
c�t���ͮ]�ll5���#��� b-�+�Ps_y��:S$������$��K�*�J��6F�ݪ��LV��]9)��`���P����bGlM)K�e>��f�^u�OoR롕�m�6���T�Bd��@]h:C�Q3Ӂ«5S���8`�4��.�f�-��C�JOwOH���.g � ��kw��r���n-wl�g�y/g{����O{^�"o9q�8*�{8�D�ӯ�ŦG����[`p�P�V���?g�m�����u�$��5t�-��}�!K��/	�2�ٲ�e��enM�� yV:��Y���?3R��[�P�;��-.S�p�7�[C�����s���':��:�I�Dn���2��=m=�s�j�E��Mԕ�<���x��6�ɔb@x�ܕ;���E����x��m�+�tp��z{z�����Oډ ���#�_qH}/K�i��J���$3�˚Jo����7�1���a|<��7_���&&z�j�k���vz��9;Z{�Z]��)lc`H���
C��t�w�B����������Y�g;��D��rj�`u,��*��+8y��t��ga�4D�
��	�����c�#�B�ŷ5���,)#ᗶhX3KOY7h�Cp*<�ʡ{�R�I���
*�&��u��i]a�o�)QeBFgS*����3]����ญ�x������3ΐ.u+=#냄�!���d��pt{	�Z��FNE�6�J_q\�xl? �P�V)�X����DĤ��bSr0)^;.�ͥlӖ.��j��仳ȫ� ��[£�]�����JE�9@dY�Y��mQt/���mqNYj�W�/|��6�@�� �h2q�l�̽��rec�T�P{�L�\�67v0�)��X/?d�R^V+C�JN$��z�u6�Z�{�*�y��
��Y��n+�y���5��<@��Fk���s�76�9z�"[���R���������8��*������V�G/Pt�T
�zx"&E��xە�Dp��Ȥ��T9W	է���$:fL���0�E:g
P���Yr"���Uns�\x�r�EED\�	��M�8��9TU3�Q;�����g8Qr"2OJ��BC�B�P\�<x��b��P\q�^77eȹr(9�DC�G�&8��H��B�����	�^�UDd��EEQ�@��r�:ay:�S�H�TY:��AU�.yJ���D���]�J���������='PB��x����Br�M*+r�쌅�&�<a�(�/Q��Z�s[BuYr��B*���+#�NWV#����*�T\9E]ӤTA�$TAx��p�Tt���$@@�ڙ-�	��+�(2�<��7�{�2lq�M�_T�o�uj�4D��u�i͟.|5�dc���W�
�6f�8�jqI-	�p��S���ݘ�����<ub�;��)>/�D{����T=P}[��pk:="�1E�«�n�"v;����O{�,	>����O�"=~�*�^�4c}�h*��z��D��F.�{��N�N��f��va�� z�o���W����z�C��L?N��t�c=Gmvz�6��L�'��p���_��f�� �=G(�>܄j|���|:w���[-$�9�r���Ŀzt4�+�g�(Z#����Q���;C���@B�%u=�v*�yp��p���~�~���	�|�f�
����7���g��S�����`:5�W����uܒ��p�T���{�qI�G�?;�7���7������O�Y�
exL]��1��M3;ګ��p�Nu=�E���ͧ�*���B~����^��>�w���o��ea�(�gi�ؒPFY�%������t_��Iی�C��VvF�H�I+��5�3��=*w�¿J��W�]�5�f���>'v�3UwL9����:�B�`
����ӑ�隣���o��L�Wa�u�qՖ��M�U��:��,���i�k-
�Fi3��Ȳm���i<�[P��-�'Ϩ��_K�j*ͩ�	�T��,���
��7]Cv��Krp� ��2s��|�����b?5��Ӆn�}Ic穩���=�W�z�r9�ԇ�2�f��wl�<5��w�Zn(��'U2U.w|�^v{�;� y���s�Kޓ�W�7�r#�u�d/u�q�u�VE�����Fz�e�~�G�����_.W��>��5����(� jN���b�p�^Ey\og�c���IB�$��>�Ju�{GFg�j��ǫy#�+�	���e)���H^���^/ w���{���N}�K�Y�y�yau���<6�]��=zz}y�CӦQ�_I�x	���ԪB���<ub��}����=,c�Q��g{z���o��u$�w��Ӛaxd��x���AH�G�ڜ�Yu�o8P�Oנ�~�jgs2�����;n���p�����~�Ty@�>,����@+�W|�CDD�T��~��=�����q^��c���=��!��{�G_��d�;��$x��ڵ�FVoc�Y{�$}�kX��>|�G7�l�L�x�G��A��_q��s$�P�KS���{=6��[�QO{�Z��=��qS������ƿ�W�7��㞙��f�
����_�%d>����	���[S{r�qi��y�h��V��}�+'�Lf8����7F�z0�6�s���^�cg�mzʹ[�&�J�8��t�d�{@jN^�
��y��.(��z�ʑ���<^�ŝ��7��|�d�a�_&Wiv�jN�,�3+�5oxTK�f��zV�����%�#����Ŷ�fM��>��������g�W/L�k�������F�a���	g�iFm1֕�2�܎+��K~�۹5�]��J��tϽ���o"��z2�>%h̯3x�����h��U&}n��˜r���k1y!F�cк��u�G���U�OO��C��͹���|#qv��O��|맵NL�k���S�D��S�o:��3�%��֧�L��s����sT�:v�^�7�E�T�g��˓���g��Ez��G�J=���
�[�q�x��)׼V��q˪~._�r�w�	~��Q���3���\�E���&XR\��=Ҏ�X�p)/Z��3�~)�^W�2����>�KaE��(�1�O�|hY)t��x�Tϑ��rV6hydv��z�5�Q>�ꩣY�{��.D���WW���k&Y�Ğ�3ƌ�b�e#2|�x��>�./�nV�sW}�Z�7���ǲC�G�l{�K�A��,�3ĕ_� yL9�=P{���9��nt(��s6�2Sx,���Vқ���]ԮÐ��Q:�$�J��SVM��c-�]��R��;�#��_3��Lf��ʸ^ z1̺G)����s
��5�����9��yC'������{F/���b�rX���m�{�M>Nf�_p������z��"<���g��������w��p�Q@���cN���چά|���=N����X�.��)G�֑�s;��'J���gG������,�+�Hx�p(�wu[���/�$��d#v�7 ��3"���T��^��g�z��Ǧ{I��\�-�#�𹺉n�@����yY���F�u$%q��SBY�P��;|������1��+>/��I�Ϫ�=����֖��s'����TR��)���c"_W��Qkf��]Lz�vG��jG��TF^��z�H�G����>�����4
~��
���d>7��TT��Ӕ_�Үp-�0��5;��9���v|�m��ήM�c�鸏z�`sC{�u ���������TlX�%�m�٭�J��>���9���U�{������n#=u�=�ݖ.<���\t�kq�^��E�Z��5�rG�"�ӡ]e1�}����^9Ԫf}�q:Ϸ�^�?~���G����n�j2g�4�k2�99����tlR����{���{ dK��W퉮پ��w�5V��B"|�]~���复�	�=쒏�dUIyl��q��ك��s�[ 6�Ov{U#�teۗay�0�z�-�Ktx4��ޡ�D�|�쇸��%�KG�J��1�el.c�;R�xD��%J4ݴ�E�#��[L7�y׳���\L�RR��˽�
���q�gIݳ0�O�bpΝ�)�V6�]�G�J�ù�n�y�o��Go�WSe�z��9�u!~��(��g	J�3}z�ϦQ؊rW~)����.�Y���{�,/|+"�ҽ������+և��{h\5�#��<jJ�*���t���O�w����ʫ�g�G {�Ǻ����{��g��>�}^u��{h<	l�$�����#��;=�ֶ�9,��*2I�ڟRg!�o���}�'���t�����Ӟ,�p�>�u����!�� t@r��[r�����_�
�W��}�h���TU�~!�Ԟ�.S5�=����2J4���=`��@�o����Zdz��w／��ت��eW7�;���h^��߷���^����,�"U@�%z����ۈ�62�#u�v��rý�mD׈ѻ��e���:<M�z���~ȫs>��FIh�� ��QJŕ��P]�}��˹Z7MT4}��p��I�{ԁ�G�x��k@�{/��9�L�fg����#~y�rB�� V�i���43E�ژ�\ma�BQ���F�g�a�"���*kwQ]7:b,O��o����t\��	�Q"�[\Q�nϥY�.�MNĝ=�k� ���c�rR%�A����o��,֌�L�[Ǿu�E��zfJk�ov�-����Q���u���x����6��������c��d�{ޠ;����#�;��9O�]zª݃s�j�r}�q����i�>���|n��x����k�W��g��g{��V�$節�}�@y��:8f�Ǐ�Q�<�ևT�N��s������cu����F.���t��}���n_%rX��G�iZ�Ez���>��az++�n)΃���y��'��7I������Ѳ�`��}	׻��z�r9��R�ݹ�t�ۈ3D*�u�Z\���DZn����%.p��\ �[�d_ҽK�g��1��7�����_{�t��\�(m�L�3~�m��fö�ǝ�u+�.��W��W���Ѹ;.�rN{��:�����q��}�_��]%�|���=�G'qG�U�Q�$Ϧp8%�S)L\E9	����;��n=�|}�>����������=F���I��Ȯ^�{��4�3���H=QX �X��T��O��x��[�_���5�S�Kc��9�j�R���6�g�վ1�%��x���,	"EKf��*V������yF�{n����xGQ���-#���\N�������[�[��g_L�^�Q���z���9e΢�"��fc���+�Tۘ�ٍ`��J�\��pOs^o5�1�e���.9�kg0��6wݏ��8�X���Y�S�����]��^�h󗹛{}�I+���G��x�)8yG���6�~��@�>5�" a���G�x�I�s
D[ݸ��&�6�O;y��+>����\:����;�O'�g�Du��ثs%�" jj	*�/)��zF5����0|
ҳ�cȧ�Tu���>'8���gMց�U_�\9�X<��F�����{��w.J1����}LU������/��!Q�����z|�������d3Z��G��������J|�VH�;%�
�T�{ƅץi��u>6���\?+�1m�Y����b2�_����[^�|�|�-��F�|�B��}'� \��>��ތ�s�5y��_�]�ap�\�c��'-�O>H>���)�?O�=~y��ѕ �O�Q�A�0�+պn(�>�9�JIS��v�_Cŝ�ߤP�>���z��u�G���X����b��6�nt���py��C�B��Q3}Tv�GuV��V����t���Vu��.g�Ks��;�Py�_�{�['Q�p�nY����_{;O��A��묪�!�Q�;.-���@)ϙ�G����Q���;8=�t1��&�dNc�1#�oR��'[���f ��*4�b���u&n~�{��J��=�@7��^�]:��3��uAl�*W9�u/'IX?�)%*�*�k�}B>{(͌�mۢ�(�/%�"�jBk_p�XRH5���Q�����M�͛���"�@���n�ӷ���3��.���r<�i`.���T%�^>}/�-����5��x�v.U�=�,�3^��C��(вR�2�P3ŉ'��9��#�1�=��_^��g_�����y���l����s�6������f�*X�R=U>	��:A�%��T������(�U���>�܏u�z�����φIe�$�3�*��h�:hگ_N�*��K�4�a����qV�ߴ���;��{UHۇ�@�[ S{C v�S뼺���k9.r��a�_Bʱ�g�1����Y9⴯zN�~�\��][5q֪+n@�M��^�vdɯ'�{���ET�0<끰_��h��*Ad:��c�:�����}�o_�rji�鑏��b�A�C��h_�d��=�$���Q�v8������J�bc�\�F�Y��r�w;�÷{�[^6}��'��l
~�\U�3�(���c��z���j�]Ly���5X	�$17~���\�[!�}��r.!�^'��>�� ~��
ӓ� �|l�**%�n��������^r����K�6Rx32����yW�j����o7�����-�x��_�Y��ϯ[t��]��[�������}N����\!`�����<����W�?}�6nT�IX�.%�vS�Q3{)Wa]�Qt�6f�t�z�Z��䱐�q�G\�)%>�n��Ǹ��׶�2!�����ҽ��}����F\�P�Ī�p>#�Nw���_�g6�Q��r���[��/�F��7�u����w�#_�I��ׄ�C�Я972���U骟�:�Z�r=��W�8|\�WgC��cn��:o6W��u���K������9�o��%u�ՅL���۪�;5�������3���'	������(����{��.����}�`�l�;������d������&�Q��ݹ��;�fT	�,N�,��Ci��P����Y̙��m��%6[z'w���S�s�C4��ԅ��\�B�K���Fz����U��}[�쉿bDg��x
��o�[<��~�Sy�z��Y/mkjG\E�x�I^4�E���[�Z��V�w_�z���P=��e��z��#�'�ۑ�~S��^>����p����U��b���\��$�(�B�[�ڟRg>x��[�~��'����I�����Ѥ�2՘ܿZ}Wk##9{��Þ�p5�z��&���u/�G�ԅ_�ֆ�����et^���f���߲�$@�6��ؖ��f�"ʊ�,�q�@����x`]\��ȴ�Xg"�ԛp�y3'&��n�Y�ިe���lLT٨_�{�����T�>t)�b�IQ�����Z�_N�ji�K	��;Ź:�#��4�F�h��7y�6�N�[����9zr��sŗ��pv�ݳ d�iA���-� ^�}�
���*Y#}]�H�<wg3��>I"Nzǜ�[�Ը�����q�\U���e�	��]F�c�ƚ{/�^/�aEz;�������Ѽ#�������R'�3���?z��U�"��3��%�g���,��?U���޾�εFGa�{Q���*:�W�7�������h�ׁf�3�=����6&��'������>��%3�vK◲���ܛ�/���� o�uC`���P�:�D��HFҧ�e��
p;���E����|n��y�~����;�ɼ��g'�v��[�ԣ��
�R3��Gٸ�,�a��mhwS�:.)Γ������Y璡{��|.����ϐ�9��.T9��ό��_��N'1A��a�e{�ӝ|����ǁ��z:���q��[����z�n�ޗ��c���A{�nF����*������V=�t�v��r�|���\d��o��W�x�.�K~��{��s���.p�6�#�ۛ5�h!Y��U��6��M�5_��3�ww�~7�������/�^�ؑ��{A��.=�?`9̆kSlD�O��s!�������'l
�=�I	V�[��M�:�0�M'kjqSo(e�V�NnucK/-��=�a��v�Igj��^�JA�ձqH#HU�W�>�����l`������1h9�Ww97{��2V1i�s�nW�@���.�?jNj�}$x6{����o7qe9cv$�YӈK8�=So��P&#s����w+:b�!̩��`��re����5PT�����Y��e�8�wiU���gT΅6�vs��%Ŝ��o/�:s-�,��:U���(��T�FkU�y�%�ˮ�z�xq\�c�jw�><�Ma`����T���)����Zk��o�ѩ��u���y�z�<��c��S9����xWo�H�μn���<���NŽ]��7�V�-(��Ƽ���X*�~~����JP�c0�#M85�~i��]Ӗ��3��B��rC���պ�J������jT��}ݠ=ܹ��*z�<@���os�Jpޜ����jڹ��wy�4��c�ϖtgKսu�I�;"��P�YtD��h�J�,�	*�s@�qH������R�
/:�y�Qٖ=��<��Y��K�a�
3��_\k���N�$ծ;����J�Z��{`�N�\����C>���YοS�C�w>yQ�}&F�q��$l��lU&H{�c�}"B���=�Mb���}��q����qp�2���HL8��ժ��r�g<!�]�R\6��<�.�(ЍW,u���V�A]rZ�{]GK���.W}/��U�#e��wr�X��KK@�r�2�o[����t��q�EN0����\w�K4`5Y[s{6�{�<v���n�}h��A�)=���<���/�F�kY��A��t��D2[T�
�[�:�Z�&��(��g+��.�Ռ�!�\�gK0(�y���\S}˴ir`n���ŀ�mټ�1�Bk���F� Џ,ꈣ�ǿp�[oxܺ��;��t�Z4uMS��b����5�|�~C}���Κ� [�Ы�jA[�B�O��-���>�k��<>���%������;�l
ۗ���N1{�sre�����:��F2:(�VN�jT���Q}�UŊ��b��c��q	���6^MK�.�ǳp���:�
>ay�)=oՏ!<T��w$��t��9U��5�8�S�t����Q:gR�u��JC�**�h7/v�?��"Lű]��an�3o�[���4���5��N>��KR�i���=��R �-��4oz�,��X!����Ӈα+��˙L��N�_�Pp�[3�l���i��o2�d�K������;�J��X����a��x�	�Ҕ�ge�E(���v-���ܽi��pQ�/E�-�.�ui��	��G9���Oo3lIX����W�l���K&�WƇ�j�x��8��TP\�	�eÑGr�E�q7:aDUW*�����W��E��X�D�+����ȦN��
n�7NRA�v�2#��EAUs�aERHDr���vs�z`D�E2��;
)%ƙ�ǜ�Q�h��q9rE9��]p�"���剹�US�Qq]<G�$A�X�.r(�w)ʪ9����˹�8�G"�*���T�Ъ�=UÜEA�8r�<�ˑ��Z�8W���\w9� �E\�L��L�%+P�YTS�T0�'-\IE^���
V�E+q�,�� �g";(22ȏL<I:�'P�˅�.���U�2N�q�r4�P�q G"�s��R��\��z����	˄�$"��*�dEP�{*o;Y�2�T��w�5� m�[a�0�&�F��z ���8۫[�|�<0�X:�c��foW�d��<�[f���r�)�M�3��5Z�`��>��nϠ+�
��/V������+��=�%����|�+�Q���vk�� �d����I�DL��L�w3�1t�'/����O��{���NG�/�U�����6H�,���jB��^��Q�V�񸾒T`H>E���H]T�9ǎ�U���p���Hٴ�a{U-S�7�)�>�od��C��au�1�Y�g�*�� $H��l�u�D���#pE\�^���a��}�\��*�^��{�̭�{e	����`�>4ȁ�p.tR�����GgՋ�b��܌�x�z<j9�y\U���s��{cޤ8�������ݱL��Q 5/8��1��Q�:����+��~���	�qq����m������ǧ�A�~������Ltϒ�}ޫ玉����C�R[�Ă��J��ѹ�_���*:�W�7�O�>9���"=���n��|��g��Rk�3W�U��\����J�V����Dy�UI���o��8��[����%S�̟{g�sȀ�6+�� T+�'�\���1Q-m�}����c�'�䁯ue�����Æ)O��S�guT���w�6-[΂��P_�*n�� ��8V	ժ��F�:%2�㨙�;+_h���2�ҋ2��2���i��{VsqC2������5�ۮh(�+���=:ul�]�d/jl��7�P8�b=X���J������+��#�+ޟ z��+M�ތ���Ī����}^��g����z�^�j�)�3y���u��g��{�}��<f�=V==9�U���6�o� ��=��S�R��M��䵼�ס���o��i8V���:��3�'�����UA�{��~���؞�^�N(�orqD���}��~�ea��ӡ_ՕZl/�A�p)o�ǲ%�/��{�Q����
�*�ƹ�B��P=�}�sf|3�l�;q2�P�஧�t]9Sge������x��o�-Ĺo�8�W[�G�;��N����ϮQȳ��pe��x��3�e�ʌ2=ʵ5��)ד�ꊧՔ��k�5�4}`�D{B�7�����!�]j1mmK7x�����*���e#7�=�j/�ܛ�῟6��E^�H����~�}��u�z���{H<��Y�x���0��mvi���*��\����Q��qS<9�S�^��O���!����R6�~������Pf�Ƽ}5�.9j�=>�K~��t�V,�w�q^�REC����'_�DB�^�w���^<DC�ٳ��g��Z�jF�h����%��a�B��,�Ȍt�c�2�v+�"^]�j��^�;���59&Z+�����`����`!�G����k>ޛ���Z��#c.�gL�6A$��%�f�p�ν�s�{E�^}�G�[}{�S��#��ӆ��2
5�����o�_��h��ʐY�[f3ӽ~gZ�5�P3�����%�<�):��Wv��̖jI\	 ��4.)�x�|��;�������G��5��������E�WQg�zg|K��ƣ`S�z⭙����A�0_O��-l�g�Si�S���y���h��~Wr-�^'��>�� ߟ���r{A����Toy���ә��j��Jg�����f�.)<�����?P����q�|�ێ�e�4�į�����n㺕���W!�;�>�⺷M�z}�x�*3�.7�9�@zM�z��{��)�
E�c����i@�S/�:5�����6�^���ex�u���.k�c!�Ew�ǣ���w��5�e-�W׾Q������oޜ�gN3�����
�·qS�tJ?�ͅ����,�ِ��z��2���ޤ��9^��U�+~~��<����ݻs�!�'v�3(O�b�kL����R['��~3mB���h���#�潞b�O��W���l��[S��g	J��< ��v���]��!B��~�9*�iu�i�xC����S���5�{��*�r�)�Q�c�
��|y���Y-X�y����Uk���DGg\9��a�}�;�2�0�y��������܎��8�کR��c�ឭyoa]4.�(ѧN�!�(��1fm���B7$L��Tqs��?u��Y k��A�]Kg���~�<�hx,�{h\5�#��<nc><�C=�7���Wǯy#�G�r�.����&m�S w��s�'�ۑ����NEyׂ�{h;�~K�7s,�P9��Y��,\��U�����T�s�O�3��Պ����ȟ����֯�l�5Vܣ�\�w��ӜW�ơ��A��R��|ܡ�.��G�ԅ_�ֆ�kJ1�X�ˮw�ش;��v�ڏ���W�\�]�0�d�iA� z�� �/�az�����c�nE�K��{��*�cκC��޿�z�q����]��%��� �=DbEeTQN|�<����ܑ�q���G+���8\7�lg�ԉ�xΏoޮ��~ȫs>��FIh����"�*D�����f_�n5G�zuVQ���;W�u�f�i�����O��@��X_������n58a���Z�Fd��[�:=fu=8*%uh����ѿ�K�%��?;�7�_��q�z��R����Y��V�����`�C�EC�EMA�c�zpz�V���*�6�J���0v_�duB��;�����
�`绚6�s��+C�-b��	�z;A���n����sG�פ��i�k¦��]G���sR��YE4�_��=��a����̱��8����٩�oR��R]���[彂6f1X�m\�"�4v+ӑ1j�´Ո�m"޺���d�ϙޒ�97~x?~Y�[wCoʎ�||J�0�����*}�D����m!�}�xZ]�ǳ'
��y��(��|�����;ӛ�Y��/�{6�NG�fc�釿VW���z8L��<k�J��'�z� ����Հ�7^�K����R�ۑ�t�ۃ0�E���xy�޽�=�yvK��S�f�J�LKZ�.W�x��]F>���\���s�����Wk�����P~��5UB���#qG�<����c]I:^>��C�N��7�^���F��H޸Q{�R����I�I�ȵ$�O��x>��򘸧!9��^/z��O���׷"��ᴻ7Ү�������ᬈ>�F�Ze���Q�"ĕ(w�S��!�U��2��{n��y�<��1��^�{�����;�ps�1�$��V����"��[/�H�sUg��t\y-���M�6�8PS�V=�#��_���7�_�=�.O�-�0�*�}�_��zn��q-�$���{��t�d3Q�o��W~�,A��#�ޤ8�������wlU����U�JȦ�Bf%�8�ߪeN�4�5Y���"��^1l��(L��Ձ��讧d�Qe��
w��з��[��Vj��5+�Jӹ�M���-���$/�pﶃ)�XI]����	n��{Дf�{�57�'u$`|�^[%V:jG+���Ͼ$3'v��}�؄�E�	�m��9��w��w�OV�q޾_�&'$������|�pY�|�IB�Ԕ�q#"'ޤ*��ѹ�~6�
�mW��z|��[z�S'+�|2�/�SԖ��s'��Z}ެd��y>�P�a���D��^���K��z�����~��k��$�>�1臭ٓp�>����b��B�
������tK[z%�a�;�nM��A�.�z-��7��UcG��܋��zf����<�+Oz.d��*�d���a��zV�d����5�iV�Y��v�1�Fu��ϴ��g������htG�m����;N��!�ǹSxⳳ��ˏ��>�>څ9-�p�����W�꽤�7^��z�[��^�ʚ��Oi�>�ҁ�rW���t�.�:=u�Zn /�D��o�ǲ%�/2_�|QW�n�g��tW�-w��F�E���}�͙��9�2�T@�஧�t]9SpvX
�k�+��\��u�*��SGۅ�﫩��7��Y��(�%+2�W��.�|�Ӑ���k����뭉6{��&cBc7Tmq���mwR�t^r'(�t����eZ��/a��$����/Or�D�8]��n������b<������Z��Jb#�#���W���6��G�1B�`Ż��z��o����4UZ�oWQ)(��*-v/�~w���������!��1��Գvx����K���=�Q��ӗ~�[~|���}U8=�ˡ
�kw��>��t��^���%���e�3Ĕ�wM_9�J+k=}��R�D���qF|��L�&q�ۊ�t��|��q�=��ڪF�Ux{t�y�M���D����5I.C�J�t���<�z�P��VBʰ��w�qW��֑�s;��'JA���� ��j��R�J2;���V�AF�AU}2�7\��2�|�P��ـ�½�u���Zף�7���vN�>���pz����з2Y�U$5p$��4.����B3����q���ӷb���k�w������O�������1�6��p��J$��OY��}^��������Su���j�>�s^�μ�;#���]ȿ�u�}�xπ�g��h��]���ӓ����Q�q� {�"��q�_ZJ��u�d/��6��m/m�d?:�7���ޯ���ދ��}9uW;ِnW{V2Nx5��؊u�o�>��;��Yח���~�=&��]xOG��k�&�/�H���K�����,����d���C-A>��F�utj�:��=�ll'}@�w�\�ld�ٳN��\�p���\���:���.�,4eD�I�� ��8t����s�����K�O���LK#�Q}ί_f3U4iFqrh,��.���a����Q�䰮·u���K�t�l�εp�"\״����;ԅﯺ�/��d������	Y���o�ߧ<gN|�㳷?��:����:�X	s=.Y���Z���Ѳ�N������M�W�ǻ2��3��٘yP'ȱqY5��%�4'j�O���Ow$��ѳ�z!�.%y{<�W�����!�s��B�ϮQ�8JWf���)]��[��\�wK��S����TY��@-=�>�Jz+և�ȗ����#�~23J���Z=WM�V˽J=��$Z>�>�We#qG�7�>�a��W����>>�uC�K�:�Q>x芀�vWmv�dWw�P5��D��9�Iꉖ�j���2�����9��V*��q�'�����^�/o����B�e��p�zs���Y��9Q���j�r�}.��Dz�HR�Y��R,-��J}�yu���\�hc��W�v<��W���ۈ�ݳIf�9�6@�W�^�;xy{B^��q�#^B����������R�o�o�'����l�f�� pȈ����s�������J��60�xEm��w��\��=��KV3|�%[2�VP�JW<��c�mҕ��w�;��CƆ�M��7��U���p��&A�x4�D��u��e�WYĖ�W3�b���.�̼W(��.��VӮ�dK���$g?��=%�]���iM��G��V��i��8\7�lg�ԉ����z!���zk����X��㳓�ձ��%I�>>�&_S�#��7n�lLoD&��}�J�Ƽ �18������nB��p�J\����7�,Z:T��V���~;F�K�B^ۏcU^7�9~&J�{-m�&�v(�^d��oF�l9���z��x��;,u�N]JӢ�ׅ^m>6��ù�n�^d�oVh�E����KZBO�-�'���������l��58T�N��s��2dMW!P�ؿ/g�;��H�D>����W�#_�o�������c޼����1�*�a֞ɉ�_v_�c]e�%{�G�WN���`
��+��u��r!��zZ���+˩�v���p����{{�&.=0/�!�̍�\}O���
�*���}�U�� �DwҽK�1og��pX�և�"�۩	y5黫,�nw@{&����3�N�:��U�⊀�ap:1H�y�S�L��S�&&Ϣ��dZ���z��.Bϣ7���-󮒆Z�J��XT&x9'�cb�����z�Mzfw�,�h���;W3>"Y��|,�/YW{��n&V�/�#E��㕥p��f���3e��X�=Xt*դ�H�{Os������<��� %*�OjS��a�'8����A��d��ڶ�;+9ܫ�,����GU��)#6J��4�z�5��v�v��w��ߍ�gϥ��"��<���Q�V�f賈�e�ȱ�R�	����c��[��e`�ǝ܆O�Rݤ4{�!�cs�Gǽ�Q�E��ǰd�j�J���&H��4?u�z<U{і��F}�}���q��1B�����>�2��*:UǶ��7����.O�2 r�3wL+�ث�,�-�LDt|ry�Y�y�U�^X�9��=��RMǷ�#�=wlUJ��}������$�v�_�a 7 7θ��!0�P�
�����r#�;��;��=蘜��^��l�ۭ(���k�G�Ib�I���I�HU�K�r8��|���ͫ��D����:��b��۽��M�Ni/�ցP�Y�C��(�|��.{ƅ�^���u>7�:޹������s��C�w]ɋm�̛~�@�d@u�z��+�r����}�c%��}���`��׏�V�R|�ףަ9��wП��c�L�z|��ȭ7ތ��|J�����|dg�i��=�~�aʜ��+K��c��^[�W��k����c�ӑ�uX��͹�<�[�+>�X�ٻ@ز�#E�c�3��%=�T�em����ߨW�xU�O�u萕ybo檭�����^*$�p��ďѻ#��;�;��񙂷z�ȸ �7bU���N���.�6-�Gϼ�	Ͷ.fp��|vm �^��H�Y�!�(��wz���*��,J�Ι����r�ZF��vS�*	פ��4��Y�7x��ӷ�P�Ź[wp)Yl�^7^n��v���ǁ5$�|^,q����]Vo�W�<�ӮYh�'DLfVnD��m�S����j*��݄�F�i�)�a��]�DVM|� �fλ�����9�$&R��y��M�ZvFH�B�@���Z:�͌Yj��@�ՔO(��{Yq�v;�oc��y��������� P9맹D��sT�}����W`Pc��27~B�*]Ǝ_Cz۝oynJz�+��ÒLk�p1�ξ�J\{|���pю>��@>Ujo�`�'�K�ߺ��;���.{9�|����䆖���X�:�K7l�����#�:x��p4��C�j�Î��u�Y* �����d�pn�C��[������|$��ёC
?�G����b��d��������眽3�i����z���֮h�˽�Y�]f�atxQ
��� e��I�"+!�F^�tr�/#�����(kN⣑bɷ�r'mhÍ��,����G/���؎-��P�y��':�0ҧ�wnenq��g�Wޣ�l����A���������+31�#N]�{�"y�r�Z��v\� �H�E���G��}�/M�p�gm��l�n@z�	z�s�e�2��s�e&��ܝ�ik.�R:E�H��Q�WA�ٳ�.���kZƹP�'a�<��*��ކ$:ނ5W�۫��UN�	+Xq��qT��B�'�!v�E �����Jf��]&�=���~�-a
�G���G�[??�kG��u�􁽔�d��:l���j���h{oL�T� �͏��*r�_6MMhS��s��B���pL�� 
�4T�ƿ�te�C�\��qd��B����I���Ⱦ��.�xVF╨M�>6��y�W'"����G[2P5�����EÅ���͙�z���q���_'ˑ��
W���|78(��9� �S� ���b�@b��N��!��`2v^��e����)�;B��֞9���b\!�Y�iVR9ׂT��vk�����݅����LDn�f�z�|ɬ�!37�Jw�W2!K�]Ԇ4]��ʱ�ՑV�5�B�k2�'4m&>��[�V�ػ��덶U������P�%�sn�"�V����BP��(�6˨�R�b�(�:�47v\-�/#G�<�wh�֣�E,]6�<��j��R ��E��%v�'H<���Eip�'.�Ԑ�KWX:t��`ʶ��y̷k#����ӏJ��wR�K�!]�мl<t��r��&aE�H�"q�W"p�]��\�9J��-YTF.��w2�Z�PN\vꎜ#�uB��XFQȼ�Ƅy\e�3&��N*�.AT�*M�Ǚʢ��"��r�t�m�s�"LM�E��E��
t���A���i��+�q
�dTr�͢Z��T�TG�K�.���n�ʨ���ҥS3��3ViG*�A]:���HRa帮^R.�0猥ˎQDrexQ�`W�(�'9Aq��*-+�6]�e:IE\r��s����K��r��Z.P�
�E���"�QQjˑh�9/+"uSn0��d�%p�*q���sBqE�E*�#��)g��u� ��s��8uO����,�r$�K�p��B��H�R�pP]�UDb����ɚ��x㗈�m.��K�
д :5�,4{-c2��A�Vkz�O���d5�f���xSׂļLO�zL��՜K�t��g���Kp�׳��=@���n#:��3�'�n�;�;�P{A��x��F���^4��������p9�V.t9ɞ;W�F��|�=�.ix�7!�4cɊ�}�'w�Ҳ}x{�ym�,N��t���ǲt�̱�&x+��Q�S��6vX6�8��y���r���jl���e��?��q�������{r�Y�R�2�W��.*g��V^���߲�����c��$��
;�49g�}~>�^�?��C�>.�k&Y�<I�3ǈ���}W���j��Z��m}S9�uR���B�w��>��t��^���%���,��h�d�"}���E�\��I��Nz���3�o�Ax�Ƿ:w�>d�οu�7�U#J��`u��^zw�:3�ڐ��p�����5X���]*�G!ߕ�z}I���s����ܫٟw��>�G<Y~��dk��kâ�|��*�@�7<@/�ϑ����H)��{�o0߲�~�� O��#�I�G�{I��\��]ߍs%��RCW��4.����a�~��'���]-�W�M3�ն�}��̉�["�Ӻ&t56�s�n �T ^|<#��\9��C.v����R�&>vrjjs�;�{$z�<=k�w�H,�7ڴb�%�)�>�����"��]s�zw�]�|�t����{��׋��2�f_Soe�Q�z�po�g�y�#��_��+>9��wļ����z�!����2CW�����3�����iL��Q[�^�A�i���E�ۯ�����@�軁P���گv׆�9��r�K�ur��|}�>��9E3�q�p��^���~urq�@�����q�44���\�ϵﶦ�ucDN�i��8K���l.��[��>㑽/��^\<o�|s_�I���>��1Vu�Q��O{��ЯzM̻��(�>`l�s��^��6W���j��۔vg �,ep���;�|�V���GѾ�𕟿_i���s�t�?����?������9GE�)�N��}֙'&
;[�/ܷ�;�������/d�_�|VǽV9g��1{�nx���;�a�	�,n��Th���N�U|�^>g�Y w�e��}hr���b�O��z��9�u!q�}r�%/P�����w6b�p�M:zjHz\�z+j���HV6�x,�
���s��1�W����^usU/�:�����@�_�x��_IHѕP�(ϑ���&_L��}>���^{�p��j0�Q���}^���n�ʎ�5���/i�/n�UK���i���yvq��N�r v��.&>�Ξ�7p�@��ckc�CN�]X�2@����3uΗ `�1:4�T�u�1���7��mc�p͹Gs7r�ڕ)꧶5n�R�Δ
�6���5���=�|��V�+��=��x'������*�$�1�T��8�Պ��;�EP�C��������&?
0 _�(a�A�o���Y�p@�Pe��l7(g�.���c�)E˟�>����{�������um�h������\g�pv�wl���Y��UdL���n󻌡��E/rG��9����A�W����޿�z���D��]��%��Ttl���o����{�_���~��tu���G������3��D�>�&�~�p�dW@����ju׻�@��j��3��-���Dľ�F����_u��i���M_�߽�@�>� ;���s�&o5u]�T������o�M��.�F��_K��R_�QZ^�������������ށ��xnw�O���ｽ@s��m��a
a�4vX���늕�D��
��|Z���*b�}�
O�r�oT��֢�}�+�1���^�q��@<�R3�M�����_�j�Z�S�:�l�F��U���)-��Kѝw���vFk���F�k�VF��X��*p��|N홏,^=W�"�{��c����w��Xg���}��r�e�G�����Y��D�o��j(���ݫ�(D��u	?�׎RNF{{� ;+(j鸯oE�8V��Jų���9�,Gͻ�ˆ�Z��@�}Yg�;�Y��f��C�BrMwܒ������3����s�.� */|��%ׯA�n�ޗ��c��G����Z����ك��yγ���? �aa��u�*���_�V6���d\�R�.�K~�B��J�
��<��V$�z=��I�E����ឨW^�F���y���
�k�*t�}Sg�yQ�=J�{k��*>���Wu��B�c�;%jI(�|&x;��򘿩�N_�s�e��"n��U�U�{�M�X>��E���~*|�=Ⱥ�m��Y�$�2����,_�*��}��c�.}�F��#^ڹ�gU��޿C��8�Q����Ǹ9��Y�x���}��u��׫{[5����a#�N�uQ.լb��~�{>g�yQҮ=��鿽��ǲ��S�^�z���}�< O
��Pz[*��j/��+���;^G��z��n#���8��J6E<���(���w�W��J�d ����u����>�F��o����m��}�u�v&_WO���Z�;�'���3Z�IaI-N��"~��B���ѹe��>B���S=�^�5>�7K�36����i�3]���1k�[�Y����9ˬ�
A��J����)�o"�˺ȺVGn\�7Y+�w�eו ��)N"�J&l��YȳQ�ySuTY�Ͱ�c1��ǡX˳%^=��"���Ү������;Db5����$�'�'�e�|s�;�}�ցO՞$;>���a�
�TK��q�ZiE�#c޳�r:^׻���F|����D'�U&:~�&ߧ�;��2;�(��\�=b�\	����B-��4��5yp���L���DR��W�m1��Wx<1?]ȼ~�雏z|�;��ދ�GO�^�,�QsN-Z�kݮ��vxO�Õ;�b(�>��c��^[�u^�k��MN�|��`y��JՙJ����b>�i@��I�@87�ݨs��z"��t�.��q�j�2%�{In|7�ׇ��G�*��V�|���{���b�쭓�
t;�x�y�\n(����o�|�=�r=�X��W���\��@�Ӯ�������QQ��sfx<'��:��Q�qNG�襁���w����9Eߖw4w�����k���z��ȯ+��������=�G"���e��x��65+>�]T�y�sz�,�u��0�@٠�@�lo���sާ���!�֣�Գvx���/�W!�;�ݫ���J}
���`����3%��Ԉ�|��>�	��纈�_�l{�D�����/Z�>�����6�2�r�s,��:�'8��ܵ�bz��µ�6^]WÐ�z'��UʹȺ�I����JUw���-w�OA}D�M�a�����=��|��+6�[�m�S�7��oM��V�t�ew7�4Jq�����9�M�I�&���G�Q%T��%*�Q�̒���=��t��r<���d{��q��lFgF]>��zBԹ�HO��?���� SRX���J�EC�+����"7�0�{�Q��W��.��uݝG��'J�����][5ndk�qD���p�C2����U�K"��n��C�{������uu���ί2��=����\z��h\9��B�!�� ⼦�Nz&*�>�Ë���R�$kʎ�X^�+#�W��G��Ϗ��׍F��~�\U�3�5
d���y�����{����q����u�n(�l�����N��_?+���>�,~�@��Tz3^������2�W�o=���dr7����ÿQ���mCһ�^��W&�1���߽~��_��	ȫO�3A^�\���le�5��Ī���g��n��/O������u��o�Z[U�Co�L�t_<��E�52|��{n�OcwB��M̾>9>
�:�Y^qR��7��]Ӈ���ui����bi
=�N�{Lb~���UxJϿ~���NxΜg�ٻ�C�T~�j3B�����濓�,��]��Q�fS����g�����OD}��᷷%
�/�-��(̻JK��	onI�M���ڌ���cKGq�Z5�k:�E��7��5�O�#=+�1^��SG̢Hp�&C���J��okT��v�-��lfʺ��Ӻ�nuu.�_�j��W�t��3�����U�^U�Ƿ2�KgIݳ0���@Y`E�}n�O���u�sL�t����B�hq+���w��?�^�7�}�R�}r��=�ޥ�s���#�%P1�}z���R7����t��s�~�<�+և����]�ϐ3�㞮P���J����ԏ_�<I�Q%�ѕP�#!�L��U0�z���O��"��*��/{OM�e�-HBngT�ވ�m���]C������wS-�\T��8�Պ�p=������U�^yg���3�t�}�=�|z����|}[���� [e�?(�7(UM�:��ym ���f�����B���������Rt��z����f@�,� rߌ�������Χ#�+vJ�䔼� y+�ς��޴��y�����z{IQ�����W�+~fK=�Q�G�K��Ub��o.P�	�@��;��n(���"�n���8\7�lg�ԉ�G���/ޝ_���X�&�� �ˀ��W�L��C2JF���}��2������LTrj�%}�z�>�����f��><�����,q�Z	�����o��J-���f,�犮<�2��@ǒ^���^��xs��4�����s�cH���9�\�>�}�_A�X����T�[eӛ@\r�=�P�4,�%�4��r��@ɮ�]�����h��3&f�}�:G%/� N��ց�t��s~�B������R��U�K��7�񴽷��'C���=��]-��>�>���2m��{�qޡ�#�Ӳ�\N]JӢ�ׅG?-�����~���������ˎ��w�3_��&�����롾Rl���Ta��և�WV���3�3�Z�T�K��'n3i�q�xn}�_�w�#}5�+7����ٷ:xx�Ƿ�=���`޸��K{=��3ٍ�e.2΃���*����V��\�B�X�s�.�%�ˎ�~e��q>z����ѳ���GŪ�]eV�ĮL_-jȸ��^ ��{9@;�E�����UZ��yO�a�c{���9�)E�����_|g���n���l������?k�Ϯ,�<��Jh�p��_\6^W���G�c���IB�$���@���)���!9���y뼏Z���;R��Q����ޗ�"��<��F�ei�n�H<�c'}Vbz�1���F-XҚ�X�6�}��X�ޯ�z��t�^��au�1�%���$��}��9���]�{��8�n���I��B��ₖ���;��p͟o6�\�F/�k��a�Oy�;�>Kk����1g�ħ+�,l�9����p�����@,�U�f������7wʭ��ӛB��I����hQ%ëI�������O��O�R]ۚ�G�o��?� 3�z�bRV��~���W�[�GJ�����޿\{}��+޵u1q�O2MWr�5�>�"*�1�'��@Q�^*��h��y\U���s��{ޞJs�dJ�!�c�ݻ�%,Ԁ�H�UZ+�d��@M<g��p0_B5�Lo|߭��n&E�r1#~����{;��]���OV�{޾�5�[�Ib�T���I�HT��o�e��dVH#io���A�w��Q��iD��/Go_���ȟ��>�f�
���.O�ҙ����h\���Tե��Wo�L�Y����yz����Y�q����:��� b�rz�0�C�<���9�,�p��('���f~CO-��Q]�c�܋����z|��ȭ7ތ����p�U�/��<I�F3�����[�⏴��7��ז�Cu^�k���U�OOV_���vx�֐�=�=ۑ��� �h�AݨwY^FC�p��~7�u��ȗU�&ײK�_�e�j����}"��=�P{[��I�
t;�`�t;�ʮ7W�F�ˁ��<��h�����\>�x4?y�:\�)���ˏ�f��ޞ�Ќ��]�cw�ֈ� ə�EYzMf�"��q�\�\�J}�!z�}�%�n2
�;ke�f1=�&ftHL�gc���	o&zoU�����mnuu���܀��������z��o���rϡz�q����=��Ib��T���~�#@3�/Wy)�+gǧ�w}p+�k��ϥ���q�������{r�DY�R�2�Mh{�#���[��Z�w�=3�7]!�cf�Q��!>��z���J��u����Գs��:3�\�3�Y�y�G��^3��!u2�����<�yt!X�;���q�=���l{�z/��=���$���;���r}�=2N���$��>UAc%��>x��ӿi�'�vžπ� �կEw�;��9��Cn�k�W��Y-� r���؁�l�YV8����A�{��������3�_�~��^{�F߮����24��*�@����B�;t̳VeHɊu�~5�y��Y�.�a9�6a��޿3���n�p{�U�C~s%�$���faAu�Q5�I8v=�9%>�sCԧQ��{�F��W�Ǐ����ƣ`T?g�*���j�i�~��ܮ[��v�G������^ңqE����T:���bӪ"���2|����g�A�co�c`�6����co��`�6�6cm�1�co����1���1����`�6�����m��1��P�1����1�����|��co�����1�����m��6cm�`�6�獃�c`�6��1AY&SYc�L�Y�`P��3'� bF���R*M[��U����42�JT٪B��5�L��6�Dm�T6ҋA���6��%DH�m�X	k+X	�ڵ�eJŵ�+=�R��}tqekkce�&�Am�ĵM5m&��l�J,L*�u�E�6������\�UQ���ZfZ�-e4���f��wuVȭ��b��j�f�$�)��jlMd�զ�jVV��ck+e[6�,��5�i%��6�"�M�Z���Ml٨�V
��f�V�ٺ�U�
+��  ����҅��� ��;� ��{^�z����<��U�q��^�tO�G��5��N���^��J<��^��]=,�mY��m��2U4�kf�|  w{ꄕ[xy���N��5�;ݪozc��F�.�[�@ ��4h��N=� ��m��( ������  ����z(��(�.�8��� �Խfh�ef�k)���Ե�  ��h֫���[��OF�-�=���uם���w{�������z�uU�N���]u�޼y�ո�.���=U٦ٷx������!�b���w9��62��>   ǅ}5F���g��zw��4�ۻ�.t�
�ֱ�޶���׸S�Zd{ug^��h:��ܴ�����y����w���z�7��Z�[Kf�MD�وV�U��  n����m�/v�:���������`�y�[k{hY�y�н[lm�/9��WN���ۓUw���]�%H�ܽ�+�{�lZ�X�C{i&d�EI�����{k�j��  �Z���v��2� 4]���{k�:9�:���J�{�{oN�YMv�m�cݓmt/\r�.�떇7�� ��n���m{��m�oOm��ʓ�ݷ6���wi6��V�j�z��  �� }e[.�=�fa�S���9/e���]���wwcG]g�{�kOw��׵�i�v���n��ۻWN�zh��w/Y֦��:/O]��j�n���*��i+5am��-o�  �>AZo�Z���z݂��y]s�t��n۝�ν�1Kx;��Usn�G�[�f�z�{�P��¯.���(��^mw���v�wl�w�P{m5㼖��V�*�V�h��۵�ݓ|   ��} �l_k�kvԛ��<��Gy�{���9�5�e=�GW�w�A��hU���^�k�{�N��n�ۼ�� =+���={�'A���i�eG]Ս�n'�y�jv�  ����Wn��Wg<s��0��m3ˇ�luЮ۲󺽞-t�v��[��vV���zkO8��/Zփw��W�Ҷ�Z{{Q�٥����m�:)�٭v�f��h���� 5O�Lʤ��!����S�����  M��U$�� ѐS�A*T   E?����F M)4aR* hhx���g���O��o���<��ζ�;�Oj�,�^���u<νϸ�����/���INg�`ILHB!!��$ I?���$�IFB		������?Y�=�������Z����##7b�3rf���_ץ<[aE�(UʹV�4�ҫ@��,�])�tN�P��M{ǁ��`#�^-�� ����3��*M����z-[���X�ё�"v�]�N��F�K١��zj�I�]ک�E� )4�<@\�����&�>��P���Ů�F6�+5�j�q���R��-�G$Zna�Sq僫Q	Xl�$UM�,�w��m��%Pֆ����&�J�8�����lV�h��X��k6�hU�	�kwu�=��O/6I�b�d�]��n�i���h���O 
eJ*��[��GF�2䂠��=Omժ�bRw�.��7�4F îի�T�ih81lW�1�b����ъ�*:Wv�Ƒ9������	W�^�ʚ�B[��dlxK*�N�;���@�vDqiӐ��U�������*;BU�F��T0H�֋A����RkBQi<y������>�F��hT赵IH�$��#��C˲�����^�kRv��G&5lL7E���/Aڅ�5{ @���m��M��aYO��x�U�̞�0�:�b\��#�(��׏!�Z�X!�
BV,s$˫�/ �%7� %������Fο�Ђo.s�X�0�է"T��A�.�)v���9e:����L��vu�C]�Z�F�����v*g��l��ne���C8�^�ɇ2�������[Q:׶[D�t�,0���;
��ϰ"D��J�*�-P�G�yi�
�i�P�"�t��&oF�ra�غ�5[�
�mQ;�8,�v��q���� ^�Pw"��Z35��+�L��N�#
o����;V�f�5��۬Ö�3��xu
f�6����av,�rc��%mSy�Ir
�I\ӫ#�Z�I�	X�֡�`��!��J��"��j�5`M�E�j`R�XSOƭ�OK�Ӊ�F�KOf �X��r����P[�]a���xּ'F|���FMyY��
���ۭb˻.`�����7�Y�Gdu�^��ll�bF�Y���]H.=֡Ņ�[r#�n�Z�T4[�6�����R��b�P0�ٳh��Xé���Z�/ T�h
mc�k��MP/���ЈE{g)�f����ڜL*FL����Z��)�"�ڡM���vaB͢�+�+��v+E�Ph�0�:�`����h�D�%BNe�̛���L'��Җ�b�n36�	��ۧ��t��d n���L��ב܆6�'w MNH��+<W̽E�ǳ.�L�O��#���6J�6� #w�o%[#S����kKt94V'U�r9�[�ؖ`1{�$N�G����J��������Vk՟jIK���䤜چ��T�#��	��[��I,����l@k[G "�4�����4��fl:�z�刭�ӎ�J+9h�Y(��������0\�H�ۣ+BJ�ic��
w3J#�BE�{ �$Ь��.�๬�M3Z�Y3#�R�<��iVi-���Fd�t��	��@W,p&"Ax������S"��̣�ҍ��շ���R������̰�
�O4�
�K�i͠2�1(��5{����>a�X�_b��t4�#�KC'��j���A��
ub�Ǜ���X��;T�k�n����a2��J�nKWq;���R�$��{�F\�ڱtT��3A@A.3l;*�U-^[h�d�4� ܽsCR�ۃm�J8B�z�3f3���VGn���l��3������&ŧn��^n��LL״܏w�커rB7���m27j���R:$(ɘ%#��0��+ǘ�Tk 2�`m��6vn�<�8°], X�KR؁e�A�Ix��/o*i#(X�6��U�Ҭrޠ����A��n��H��Y2�a���5e��I���=�)�@:5�u��c�\3GP�`Y�WaG~I�n���"0��z˫���(��#������<��M�[��kV]9���+��J�M�kA��j�X`�[E�	n���+6�F��EB�V<���.�)�i�\���ұ�ƺ;�Y��ӷV��c&YшǕ$mmXzuQ�����4��įe�5�i�ݒ;��	�n}�|�cyϵ�7pI��	����'���N�v+4�L�V����,]ƁY�Q�J�.&�wB�H�M�K�b%Z�Z�u^�7�T�o��(ٔ�V���C0+n�l�V\�y�Z�q�!S�J��e��`��:U�t�1�6��_]��9��*Е7���Lc
c.Q4st^���� �,�pAiD6�n��VQ�Vǀe��*�`Jt��2�X�%�b�ͧV���
����vs�t�ЫdĶ�feEܸ)㹅Xm�ne���uMP���E��T�����)ae�w,(�&����-4�MSB��p��O����z�WY���T�eֳ�Ҍ���v��ַY@���
�VØ�7 �(���N�˴�)�'�@cgr��Fٓ镙�J�	�ܛ���r���Y�r�����R;Ј`5�$�� J�(\�m;T{J���S��l��,�,qX�d����h	,i��,d�cUuy��*J�)T��;KRрp�GT
ͳ����W�l�gφ�'����0��a�(�G���T��W��ZWy{��x�*����Ha:�fa�2҆j�6�Ȓ��\��-xjR;��Sd�E��%�"���y-���c�@ͺx��R�V\Ď֌�E���]̹f�L��h�O1ݼv�e`Cq��Wr�d�b	2Mn�B�DJ�i�m�7Q3x�7H��+���uk���=�І�å��]
�.�"�-R�՗M��l`�c��d�L�c!(�U1n�ܸ����>j�M%�����[�b�$L;Y�]�d�k�
Ũ��T�.Bh��)J���GL�ʉ:�����tF�d�f��)B�"H:���4�Z�E��,V͍�`F'�����m��d��c�*ı�u(H�kwK�U�<
������1;A���'�n��X�e)���յL�EEG��Mύ�ul��u�˸l�����c#(YEFV���[7P��(ݷ�G��d!��5��̖2���l^FUdѮ%6·Z��� �����ɱ�!!A4O<އOL��>#mI&e0�p�����1OV���:�cRN�pX�d�.��G�Z�)�ѬKSu���VM�)抭�1x6a��&����W-ñ�����@���/���Yt�K9�ke��U��l&��b�0<��� ��fӔvCD���ӹZ2-��e�'W���mP�h�(X��W���Ӗ�ԽW�z�5{��m8�1�e�h6m;n�8�²c-�f��
�{��f*0�jU�`mnV�#oJ�@]�@ܼ��E^�5&���%�iVM �u��D�ӧ�wJ�v��n�q=}��͟?��9ٺ\"#��q�̱ۛ܋跴�����/�m,l��8�CV���LwKL��-����@:nVWWQ7�RA�"�죺��s �6�d͛N���LId�ʙ-�+�gKL$��*āvFm�\��u@lJ�VjݸGv�z�������zK��<s/�zKƗDF66���.�ݼ����w�0��Y�j̼O��,�Y�̓�wE���7h��0c�n�.m�ḅf�ǆ�:4����ފ V��˚Dn�,���,��/mk�)VwM �Y8r��f�FPѵ�0虶�ڥ;���i�ۄ�Q��z��p^`��>Ւh�Nd�6IR�Lg%�Gh�tBm���#%���oj�d9N�՗*�-.��Sj�V��a�Q�\5q�v�e��j� ��a(eJB�v-/�{���0sP�,<�+�������p����Q����`���L�7,�ئ+8�e
���/(ǒ
�p(����Wݵ����X`*�:�PP
:ʟ����R��ǻ4��)�� s�ZYkwa!���h�z6FK�t�3�yq���q=(���<��ہ�Yd �1�+h�%L":f���vV�	RMٛz����ڋ�f�k�QS.�-O�V,�Ҥņ�nɢ�h]"Uf�c�Ol7s�im�'N�v�w)��J�4��jܻ.��Q�H]�#-NV�P9@�Ksw5�4����Xʲ��1�%֗X����7�9Y������J�"�*X��Ux����ޑ��40><�5�$H/;=�V�̓.J9�[���W�R����*�ch���ǂ��t�7 s)���ڥ� �;PJK%G`��-�qXՕ����6B�Y�J�4a�eK����U�=�	�J�o)IVL�r�*�;Y1Iw����+45loa��וE�T.5B������p��`�7%k�J��r�#��j%u�`
�rY���bQ�>q��0�Ԟ�"H6+؆����7K�rP�n�Q[�X)HeѲ��qTPi�N�j�}y[�H��-h�ʌ4�*��wp��O3!r�w���N�vF�J]���)[9p��Ў��ɚY	�SMx7���u<OZ�N�����S�-�%�W���֛�i=�ƪ8TQ`ɥ��O-c�K
�¦ޅ�Id�oKE�镴6�Er[�(��D�Wf !"��xҬ9B�*@F��w��l�d9��O�e*�F!���hL�VNj�"l�r@S�-J�.ձ�;�s�`G,�l�Gn�}�p�GN�h�vbD�Ԣ�);�L����ݼQ�6�^'9W)����F�F��b';������=$VQ0���U����]e�s�l�	ehѠ�sz���Ч�EkY1ӭfrP��Pۺ6�vA��"YyOoN�dT��F]�ۋ,��ت](YwO�q����9*͒�	�YL.ֱN��=92�J�Վ�֞];��vmZ�2�Z���@��a��p��,�tf�Cq�w7wW���!�&f�)��e�CE,kCj@hT��5�s���8P�e;%Aj��Wl��*T��Y��B�6��b���PG��Ɉ],L�r�k̉��gu	��{���ݺ�s5(���f��NkN�`�9�B�(�NV�vq����������ʑRնhS �xѺ��r)(� ��K^:Ie�c"!���R���T����T �ddպY���Z�Kk�lX��u�7&��CV)� ���̷"��<�tQ��yx�'���Emh2�V���Aq1X��P��i�րi;ˍʙ�L��Ѝ�è�J��Ѧ�#��C��cn�+_M��٭7��!��,���u`�(�]�鴨jK�(�&�ۄ��X��m��,��GX��5W�/Iv���]�"�?7tEP�̋ed�!��ТqY.�
ǻtݽ��+s%�V�V�&���% It�E�V*�n��4�aZshja,�&>�����d��/vsi�K-���.�`J/����][�R��YW������Em�!e7W��r��ZT[��ԫ��ҍ/h/�#z�6�2e7!���� 0Y�fV��ҁ��ƕ��$Q�؃�����4;���`^^
g�ŷ
fˍ���y��F��p�E���&�쬛y��,5YD0�,¥3E��kz�������wR�:9,ֈ��Z�`�X�	bPɎv0�̼�vav��(O�b8������.��tmlu�{X/*gt=Y.*
\n�b]���h\c��޻6of�%��υ��a�W*�Qˬ��$L��)m�Si�ڬ�Z��!"��ېh,K�������k�RM	P�4ީP�
�n���Î�M`�۷E�=�3Q8��8,�0����יD�5 sm
t�9M^h3�%冞�Z�d��pD&�]�&2���oAð=پgQ��_n{o/2Q�*W�@�ev#���x4PN�H,�[a��Q�2jE�2����Fh�	[(��e!G/m�[�RQZ������b6Uƨ��7N���̗ �����e��X���R<��K��-��4��Vlۅ���1�oj�7�����:b7jZq���I��[�z�)���=��d|�h%"�0��� ��|�(l$�*�8�:����j���l����"�n�fQ��F�q���X�GY��˃X�mĶ]JsY�԰2��m5��摱7p��V������	U�s5E ��q�7p�È���������o��%�&�[�{�iM:��FJA+�a+��/j//3u&����I��ڰ!�%�SB�f�ݏKV���sb����II��c$�"S���kN�bۧb�Ob�C��
��AQ\#p�U�����ig�Mn];ٻtܫR� �:��.-�\���YZ��~۴
�ՠ�뎵�%�V�l��jK�!Z����k�ɂ�1"r�M��HG��#K,�3���b��7)�X\	8M�t�����QC��D��!�x�`�fk`(G>�o��N]�����#�,틘$MX�Qa���m��)]%b��vn�^M�-c"�t(�(�Ֆ�� -˖���$��pkJ�1YXv�n�gu�薶^#�2�TJ�T��C3�Vq�ȱ}�#�j��ȩ؇k�i�{���<E���g�)Y�D��=�Ū�%v&���Höj�,R���1�Sf�t��6r�S:���Fva�X��5e��e�	r;042��9e`N���b�j�^P��1R#���"V�Sj#�>g@E��+�@�)Vc�����A-)�MK������ת�'B��y�w��!�cC�S2B�=��w=��j�TG&�n�4Ż��#%ҭJ)�f�V29���'e��Vܗ|��.�ǥ�bn�xiޫ
�[qf�G�����m�R�ε����{9�#��`�����qۻ����-z�>�g����|r�9�|��C�Y}� �nq��{��:�*�����~ju< ˼�n4�NW["FwTZ����q�u����g:��ٜ���»+�𻭊�,��;W�����+O7Fdt���S\�g]pS}���Eҳ�Hu.Z}ܪ&��n_��i�udB�jpృ�"ldL�l��Eep!�%����F���ڂ�F��H
��.��mvU���ŷAݾ�\߉�yg2.I �p��Wh�:ɬô�pn-s@��B�R�1!F%^?���%��`���,��ϛ��jVb���9�z�r�`���}��p�I�h�J����"�*�/�U� �ƣ���.7Y���%���*J���Vkew]Er�o9�����)w,u�uY8�W!�k��!4
]����L�/{H�{��P����2]��v_U��kOk��4��rnv�q@b�[��T�
�<�����c��6׎̯�!-��>}9��]��}]��l��E.����:�ϥe�jPU��>�F欩YP
\�\��2+*�wQ{ D[��v��7��=�GՉ��|d鯳�`�j]ec�C�L�4N�� / �[F���ǃu[U���J�S{uR��};�o,<A;2{��wm'�͠�条t�]{P�j�]���i�E�KrZ����2��u�e��j�H��i�8H˂Lƹ`���H3J^H��]A�b��*�CO��ճ�Y��78�;�{�rܽ�T�t�ub��#�J�)���`*M@,P�2���|��(K2��jȻ�4ݑ��z�U34N{S��c6�F�}����D�2CC}���Ht'�|�Y䳆�r�6OhO�Wy�gU,�V�s�!ش�)����I\4t{�SD�cpq�EY#��xܘ�P�5={�x�uiV�A�fD��x��3�ֺȡ� ��Q���:��i�p5ݓ�h��;%��ٳ.͒��N�Y���� m1:���<�6uʷ:�B/�<���y���, &�3^�le�g��Lϖ[��z8>���ھ��F�������C����%*{Ε��Op5n�YG�o�O�B=�fݫ��%��n��a��Zm�{��%y5A��n�ͮ�93����
�������Ǧn��h^�nk�X��R����.�e��Aݞ�%E����ض�f�Ě˝*�!�c	m��q2^o*����k\�CQ`{׳��Q$gI:��c�Ư�c!�}��|�c��*�bb�^"9��S���k�qgh�'d��O��n��x�
V��m��e66�e|{�ʾ��il�;����|���Ov�5�lލ���aN���9 ��UY׎T[���:�n�<$�tP�i�+��V\0"]u���މo^���9ح�6��~��|:۩d��K��SVo+���g�P�[����'�(
׊����R�&z�N� �8:��}�I3m�$�B�FDn����fP�t#�Zڲ�;�!�����{��/oc|;��)�Dǖ�[�Q.#^u�On����6��4��S���YB����`Q(���fR[K"ŰhGT���@�.����*M_L.ܲO�8yIc����u+��d��@(n]�!2��3��Ku /R�`��j�N�p�Qq�c:S�]���!�J0�n�!��a��+.���������1m���2��}�S�L���n;G/{	k~+`óN��	Ű�f��-�[t��� �+Od�
����0�.�����>�k5gr��s�0R2�D-��R4����ثp�AmZ;L`�vojb���oq�f���]A�p�0b\��8�*��6V�/[�q-Sf#�b���,<��S�ml��1�jF��O�k2��P�p�N�b�h	Li��f4*��79��T�R�O���`����%a�6�7�WJӜ�~�^��8�uǊ,䏜�Iᇔ���U�W�^��y�r������u;�໅�ޙ�8zj�el�5Ó~�3��	^�� C�w(�nT��N��qpAA®nˀJ6ޅ_W ��K���6��=ҩ���n��RwLqW��ө;2�-������1�V���c��9�hM����6N��#ݦ`v��Z���^��Q]�ƐE��J��m����C��o�jX`��D�]x|�yC��47��/��v���m�fu޻}�#jqx����Eg�}�j�� �-�Rk	�:$��������#��z��:���8���:G�:�zm�����PqٍԶxv9��۔�j���G]1��:���rT![tL;[�v$7]��d�����j���M��X��&ukz�N��@�Y�Q1��o�
1uǍM���۶���)c#�������h��2�"޹��h�����G�G����[wŷ����`��y�����l΀v�Y�-����U��{�/u�>�ix������@=�Ԟt�^�L�?'�6@���B �]KoH�f�	��0F��a.��Zm�徎��I}�^��l�fP{�+�g�]ؓ,*ߺ�N�i�����b�G�s�yiJ�[a�	,�����epa�ǩ��4b���	��G�� s.���K�Zc�7������e�`cH���v��<�v{7�Ev]�Z�x���3�fʻ��
�Yn�5sJR�N�|�c	���4{�Z����I��xe��;p:��!�*�۵Q�Jc沝� �(iv񋖔�3C�'G��[X����Y�sK,j��o��>���&�(]��|���Xj]!�a.3�(m�@��h�k�=�&���I�*�w$��>�+o�~Ƚ���㲕o��5K:��+�6��!��r8�"츊��<���vQgp�^01۬���8l�m�x(;�Q�z]DͽM�Cw��;s����U?&��Ռ}�9`�:���Iu�)a}��g&^�ۅ �'�YR��U����.��IYk��n��<bqa�匲���U���I�u_g# �)הy0�Tu�{Q.���ۼ�ȝ9�c��<�ﲝ4�V�X�S��+���-���-�0�Ri�ZJ�6ш�]� ��f%]�;���}���Ӕ��	-��җdq��2��r�����/��1�hC��{Q$ۛ�m=�!QD3C���ЫӺ������U�"��j�;¯e<;bh��o�j]�aAKy-J��0-C&�J[���$4�,K��VwG^�'�ө���גe�wz�*u��\1�w(� ��ˮ���q�N+w+pYѰuCI��S�C���FZuo�C_�C�8�E��u+@i�'�`H\�{_�+�ʀTzp�6��*WV��Qh�3�F��'Jy�c����e��;7N;׼t0��sx��&<>��Sے�-��R�<��/6�����5�l�:Ś4����H��ЎB�쨩���Mgtn(H̖N��>w_bя7�U�V�m�/ȍ���kn��Y�ņgu�N����$��lg��=��v�ʴ1R��ٴ��W���v]��L3-���(E��q�y�7��}@t^��1F�5��	��b�wdt��݆���x&��]J�1�i�u/��
u]�V���cu��ű�����,H�����i��}�Gw��������h�|�`��-�.\+\w�>ǁ1������ݙҫ%��o�̈���g73y��1���:���JV���O�=���^�▧ci�`)�P���r�,n��*K�hіܝ5u[:��}�oHm�gܮxL��ym��FxL�U�[. �j�r-�1��2��_�@���5W��z�ۧ��g{����#u.�с��+Zq]izp�u�)���I����Y�cs��R�V͉�Üj2�� .o���mo�D����*�O�g�2Cu�T�ku��{��c($��������ݞ�ϩ��Ή4Mt��gd,��u�2`㋨�q�h�<��ڂN�}�k��/|��-L��8���>׫���m�X�|�V@l��s�	�\�ή����n1B���`�u���Y"=w���<��h#"�xA�f��6��馽���^:���\=B2q׋��d7l�M�����%X��g.ŝ���p�{����Uy!�!_��9�,�����L'EN��5�渧ت��&En�s9�
:s�pI�w9�xA���N�D[�9��"�.M[��N���.����l:12��qeolKnge��ԝ�'ڧ]���H���.�-ꠃÕ�2J`Z���������1;j�^;ur]R�gaS&�Ix�i�֦J+z-u{r�(ӡWKn��cZXvv���X[[IwU�b5���t=���+;�^:7M&�΍x��ϯ�[��X`��������p�}���3mw�q����7��aݙ��[��4c��(�����Iv3%�T�#4�#�'0)e��l��mnԸ\��օ��8#\g`�s����0��R�\y���s�9V�?ns�uP�K��w�k2�Nu�)*꒹��9-`zn�t?:���u+��[�ׇ=����G-x�<���ɛ��'K�`�8��A���8K������B�4$1����^�V��{�YͬT����UȬُhL�"� �}AM
]���o����M:?��|���Ţ�4@o�Rxh����2�G� ����U�X�4 T�dLo����c�j����{�Q�;��uc�J�{1r��2�m���U��J�{�榊��!�v5zw�gI�ho��q�,e�ъvKЕL���er��E���{2�/1C���MP�G�*�u�(e�������Z��-�5�ً�U�yq~�oz(w�y��	˔��H6𮴛�ͥ�Ո4�U�XY�x���R�n�Љ7��W{�Wv֭�5�bp7�.� ڹ~����_R��!Q�Ȯ�hs��\CS�XfU���K���F�g΍ܦM�9�/�)C�0���e�)	n��b���*��b�S�D�c�}�S��8}�L�3fw�*��U�����V��:H�"�˽��Bѕ�>���.�ܺ��j�
{fدҌ��Zk:��W�+�V:@�ǲ���3�Ǘ7�_��F�x]���O�;!�1�K� .���7�J����U2���'��W�W�g (d��u-s"֣�����ӳ���w��&���?%�Z`��qd�����6o�o�c����b�{yQI�1hN1�f�1��PȢ��G�3�gt�K�������mMk!z3뾐�B���Ҝv\����S�����ʯf��~.i����£��k�c��7���[UUn�U�e�n��_}��b�n��T���������,�1�ӌ��CY�X#MiN.�ʰJ9ҙ�(s�K��U��Ԓ#YDP�P�� _RW^ΥqV<x����Wٹa��	�Wc�z�T|v���<�w/�{��': jv�;�J/�� �m�ώ��$���J��K�VAy-<�'NM�۱ג�r�5��K���Z"����],�kK�O`�可�gNx,T�z��ׁ�����J�(N�lu��$��mB����P�0wW^T[Ӣ��&JKRy���/ެ�Д3u��mYw��t �1��@�-���(O9R��f�=_�{r�`�+�L�C%��<��S~ӂ�\��}��=�Sw��,>��X�|�2�5]{�Ր f�c}� ��hA���T��ɽt�8-v�������h�p�7�s�Tᛴ�oK� 傕m}ٰ��*<w�GS�z]�d̾�{/�#�ws+�aҭZ�X5,���aэ#�+���0�s�R�{��KQ��z�zɥΟ;��PCj]Ni�˂��|Ք%>�Z�LqLЫ��I�I
;j��(qÂ�����v��^.�6�K
`� ��K�/�'V'e�ve�t�X+l�FL��PnfJ�5�H���=ԗ�j,�r�ށ�_��P/I�֨��� 3�[a��f�r�}X�������Z��I+��	GԶEQX	�t�Wׯ*�e�^��z����Ub��WB���+��C��:Rx�~˭
��]�=ܱ��oj����v�wqh�@{�ӻ�鸧���0��+�{-ђ�1�ʊVL�ph��[8g��ry��T�~wS3o��*<��r��]���Pg+[Z>��(`]k���t��h��]^)�������j|�J��ݑ!�%a9Xw�����꽯��S�s��)��Es��]�Ȫ�U���=���U��Нcgfw7�S6�)��.����>�78ϴ�2?>�h����?:Ĕ���}u'ٷ庺k��p �X�E�ށ�����i��=!��PvvV�:j}N�mlZIV:F��#g/sG�>Z��D��g�m�W��*�� w�m��ja��j�'j�A�����Do�hJ�����R4�(w!� �Ќ�X쮫��U���m��}VK��&�Su���Rν}�{=�|�a��x�z���kA����M|��>-�Cw.;�]d�'\���+��S�5j@ݫ��Fl<x����du�By�r�G���%����(���jh��w�I��Y���ڂ��w~�n�j�ͽT�����]�^�������lɈ��r�/�Ccz,y�7ՠq�3b| �K\&G��J��y"��4w'�D�ï�`��ޞ�{i8�F�o��U�Ĵ����ۭ��� �B�=�}�|5�q�k�EG吤�Xv8WM��2j�Q�S�����5��٤h:�!M�7��c�5���g��(�6�e��x�����@8�� t�h:2�.��`��\��v컷*�s'�s(��]Ze:ƅq��@SE�Tr˰�\�(��^�?}�+�v��[�Wl���O�+ڮ+~h|��<=�C�i:!Ҭx�T5*�7t�`>��f	|uG��u] �;m��	�(�n
s�/ɻ��?�.>c;(`�(�	s3q͇5�{N�W<�cL�WB5@51mJ�}Z��Ŝ \k�74.<����w	�8V��>5e`�ʈ F�=|r�O���6��J�M=WA𘸷�t����X�xq�O���t���TS�]Č�����g���]ŗ+n.�z2���C�����k�P�w��ɝ��?md�y�W���Yx�^�����7�rL�f9s���.�p��u�;ӀĦ���g�:�٪�y��{]��]��)1y��u ��0�*�B�8H��{��Dww}�V���ƹ�sj6g���Hp�1ݥc�&iS(���	�)�N��W�N��lL�6�.�r.����d�C܄O��l���E��������k�%vNr�,<L�uw���@���,N��F�7�Q�)�a#çg@�7,ץ^�߰Ny�C�w��7�V���j��I��=^��⻷�{��7|�4�{�iķܵ�R��*^��'���k���V%�e�
��NSl��f.��ƙ��;��Em*�ܦ+xAQ���G+����[{�pu��8��w�H�{-�z_uE�ܯeh�?,��$hLV�cZb_nM�E�u�K�p=�zhQ�u� ��)զ��6�'G����i�*|�s\Y�﷓a��#����rNG�5�ᦱhN�֫؄4~�U޽��K�ݎ�z�G��+ȿt����/�#���嫽�tKx��"q���IZ27��^wl����9�V&u�9F$�� ��l��8�`N|����z��tѝϢ��\ KRߟh�R͆�2Q��oX���-��u�??�شwOb�����w9�nX�Z�n9H�z��{Le��j����{y�GD�9��C2>Ӊy�x#x�7'dY�F�69��W(�ȥ���2P�ѱ.T�}Ff����,`�b��b.�7i��kM!��^��cJ�6���1]tg��&�9R=�ǚEҳ�D�ӣ�x�o��c/z��չ����?,����B\���xX�z3�t4��ʴ��� ���Rj!��r�O�]�LR��̷ŌJ�k08�3ǥ����nf��B�ɻ�1�0IG>�ֹm����n�9b< �ݫ�<���9΅K1����+�.�N�n�ڲ[��E���8̱1��Y�Qz
̃�u󴃦��W,�c�\3K|V��lqC,��6ob�r>���k6s)��t�P{�G�y��U��%Y��-t^��9�5ng}�C �Eϟe&VL��;�t�{�O�#�E[n�&�p=�WF�VDyN�T�hj�ٍrQd�#���6Z�[ڷnr3:��Ԧ���U�Uϋ�lI˳�0�'˃���j��q��x�]�{�@���}��gnp�Z`o]t͂`|���/M5m�B�3]P�$6f�oO����9�G�6�����3n�D=�H��=��O`�o�xv7Ux6gZ8��5�dV�A�&���^�"�r��T�&;����s�R�K*��y�	M��ם�Nv�P(>���B6V�Յ�n�e~�X�W�M���>�h��9����k~:��lP�y��z���IV~ �!\��]չk���:q��zc�#�h��'���)�ԮV��l�Ѻ�+/O�ګpS�hHc��=�f�i��J�06+٧2�0���8���ώ$i'i)�A�)ވ1��|�,�ef�k�������^�N�]f�5c�|���@�R�=�.@� �W7 �=���v���C�PZʝ�-slKyus-=�cI��˱R�n�AOB�N)�����5da
�1��E����|���0^�O�<���Iܽr�e^xxn�t����w�����z�C���=7�ltt.s߻:��XNL ҹ\�uzkڰx�F���"�OS��^�=�ecS��հ\� �Sh��ae^H����B7�{QD�W��ϒ�\���-�f��F]=�1=3qi����{||X�K��t��wI��ۦ��Q�h1�ivs���ݲ�Uw��k�{%�* ��r�;��]A��(:Ǟ�fn�e����E8;>���-7Ou��u�mۼ�ޛ�Lr�w��j�S���$���2k����`��Μo�0���xvm���][39ۮ.�7���r%b,�i�X�W)N�}��hb�*�kR���!Kr\��>W�5��A]���1=a�vZ��n^��!���/�l�#��u�}�5�I�Si�(F.�����(i#	v.uu�J��1Z��[��]!#�C���U�Vn�z�=9��r�j���[3N��6�Wuq��eh���0_���f=��W\��%�9��l��g7�i�[��=)��V���@k��ػ)沱�X�峾���T�3�)H�<���а�S���ݼk�_���J!���VU]�JUz���i]lX[r>J�����1���:sp7Ѱv�F��M�>���`�R�MS�=Z:�Ф��.!������\B�Xzsn��:�JŊW5�P�K���4�.+�Y�!o�����L�.t�%^�����L��3%v*�r��5��7�����Va�Y��n��D����-�,�.�dn[�����#���"S�`0�� a��v���p�@���x���둨��X�[����a'�G�9��VK�N��B�e��vst[8���I�l���
E�+h�υR����3c����H5�0�p���E�<z�Zry����W����mk��혝��x��0�j'V����b�X�bbi���/� ��b��彩��{)K�(>ޓ]z�7Br�ͧW�ƞ�M5�Ha�)a��$v����0}ۅ�68���4�_ K��{w��sb�D`{t2�?,����zٞ���G�^�!�6M7�W	��s��F��fPҺ��n��2�2�OzK�i�� rv��Dqb���8s#x��j�%���9ō`�5�x�v\7&N إNGԝfL��cQFA�,���SA���;�p
��7
��*ͫ���'}�O1VmW*�k]�'W�ࠅ�[�&�IcBK��4i��U0R��x)��C$��5��^O}:��a�H�V��iP��FK��6j��|A�[�կn�f�Q!W�~l�5S�����s"�������&v@ea���C:�+��@�x���,ʹ;��Wm$R)�o���d%s��,e`��9�j������o~{%�y��mX�Y��/{6�����Y��~��k���N\�<�ei}%W�����O_N�إ�&�Ae���Ε�U��t8��EjR�4!e'���w�{ג�f��FݱF�
-˅v%��NI�r*�,�}�E*�L�&B=��D"tv��>z�P@e��#��gu�NO���/.���{9��<�.�/t���]A��P\�ɨ� �钃*5�k۱��i�˗�B�c����%ηz|7h�u��|_E���Ks��*��Z ��Z���w�b�3��PT�y���uu*I�;�p���k|�X�[�$�k��{�\/<�\q�E�ѝw��3�
[�u��pbB겳}))�]��3�Y+���>��bգ���N�(�}�k�RM�]�_BQy�����DJ����.jΛ���>P.�pŋ��b�C�gL\��떯��5��}!}�y���s�է�׽\�LI<5p2n�3:ЭB$`q�+�+]�e	Y�C�C�4ڻ=��N��@�iCr�:�������t��h]5�f���i6m0v�5�F�*>�v�=p����O�mDk�z��؝��'���.~77�b�|��}2�@�y���[%�@�z�[e���Z7����m�)n*F���8y&qI�q�� <�	��}�ʄ�/@��BVHX�Y�;��/���kA[�KF�Kx]n�n�j}���n'y�y��*'V6�p���	]F�	C�=�}M�ղ�w|�k�NܛL����W�z��&�d(�(+��#-�4p�I]Bf�>��>�z���DT�P�׵�vۦ�b����Y��`Į=�;<ۚY� (����ʎw�����&�X9��Ǟx����OvS��D��þ�o&.�*�W3�V��Q�a�~��s�>�ܻǖ�����:pq��[u%9���p� �g��}���{�I�.ܰgVY�V-�RN�Ov�:�!�8�0ӾUK}FXk��'����W.>���J�w^+��$�
.�ʷ�oC`*gJ,a�o;W���ӡ>B�9  %�f�ww ��큊@�8����R�����3��X>=��;��zyv��S�m�Z�!ۛ]I*����ʆ���/�v��:P.��O��)�>P��*�#ћ �s��+2�Z�C�aos�ujSqVh_w6T�E��WR�L�-�Da:��'�c��~��<��]�_ga~��d�S4��L����OO,D(�a![^��;��pޝ���nH��l��f�.�N:�/�)��B��L0��}*.w�����w��}4���w�P�6���ή�/k���\��6�]�,�	�w���B�f���8G,�?.k7�w�u��ط:��s½���,]�#�S�vU�����P<�0�l>�6����v�nXj���Wy��P�~�+e����j
v�}F��}���n(s��h����xQ6��aX�m�w�gQ�;�*���g�Q���n汕s��%Ը`��l��UҔ+d��}����}�v�ٞC�C!-��Z|��#�EF��[�qo])�����Nrmľ��\��2}w,�c���v�cn��X�X:�Z���c��u���{UvXF�;�H��M���j��v���!ٽp�:Zs���`|'zSI�<�@Ρ���KVxCq4%֖����'Y3�y@F����V�v��cɔg?,ׇ��=���#o���X,9�N���A�oGX詾������8:�	1�0uV_PK'j_O�]�;h-vs-;u�}��Nz��縒*��2c���u@��[��!L�16�ə.�݇YR�.%X�Ǐ3��G����yN�s�C�}�hAnf��c�jO�c�k��ݡO:��ؖ�������1A=@��Q��}��H�}x�=�ws�J0��.�#+r�ճmJ:r%wjnlS]�i��������f�`��@9��s����d���!���;�A��WJ/�d-e�:!���8�(ec��:�D�N�����:�8sHhs����[i��G�l�t�O�]徙>�D�K�7K/9ۉ�g-)�\�+,.�ُJ����N����َo`�ɀ�Cj����5�P�B���#@s ��L�\�����W_QZy�"��5��Ļg�!j�v0�#?L}K3���l)1����NQ�Lǵ�9�w��H�Ny�8�Z|��-l�A1�Q.|M����x�>e]^�x��=\MI����7%"���N�����n�}s7���E{y�;������F��+ppҊ/�T���ԗ�9��9�bp��1j���bҫ��c�qʙf�u�^,�˓�-9�3�&�.�|0�ܵ�v�uӏ!f%N����[���X-��C
.y�n���Y���ͣ���Gq��Gh2E��c����5�î�ؤ�w�z�3�8�
�}�$:��o*b�bB_ob��4���`�:��h��E��2�f�3��D�q�fj5��V81'��W>��f�o0�	�Fr�J�vB� �WHaŘ�^��Ăm��ZCk:�VpZ]������ziM�,�
�pOC�|6i�u�+��P�/R��+@i<�ĩ��t=���4%���zYd����P�BsV�û��/7�����'�	��hE�Cxe�4M"���_H�2��Ƣ�ռ��(,���7�n�P�@�*�a+���˻�t�B���ԝ�wC�z��îΜ��Uw\w�%� R�naуrL��D����Uwc�<�S�8�>��ȧ::<{���@ݫg��u]F��5uf��=�0.���=�2 �o*c3$F�k����4&<����>A.���8܉���6es�K���}����*5�r�'���r��}���$��Ŵ�9�UǕ�G��ogI�C	D)��C~]�_�q��lc��6���	8Roi�okWl��P�LHs��wDΗ��Zy1���y'��q[�A�������g�$�v��O=<V+��/x�B`��QO��Q=�h�$O=��ru��vJ���(��C����\�n�>�CǱ�b���Hu�w)��b�Z4]�޴;����S	(0�m�k�+sn�P#p���(nwB��(9�V+����L'ip8;_�mqt��U�yf���9����lX�ol�����̸���]%���I6Ab�n���y):���qe�����)N�F��<ag�/DkF:w9q�|Z��u������DC���{��q�j����������c\�v$,ˡ�*G��Һ�ӳ��C�O&ު���Pi���ne.f�N�k���d\����QF���3��N1����5����$����'6x;X^-ﲡ� ���NB��v�E��⫥���,�SМ��wp�=$l�tI;˶1#�-PD��u��5vлZl@H���T����_`�xA�}���K�8�6.<>�j���y��I��Ǡ5�m��lI��G�O��l���*P�D�)=Z��y�2�=�A�%�]���f+o��S��������H�c�q��#��|
�x�Ӧ"�'^�:��I�te@�Y=`l�K��
�æ��ƅ����s���7٣q0�[�+Rf��:h�#�����4t5��t�CQ�sz��4-_>��`
�ed���M��V�0s�m��.�Z�d�L0�m_Y�h$%-.j��R�9\M�b�N��B:#A�ґ��{z��J�{�'S�T�4�;��E}Ǭ^�Y��=��f�i��B��N��s�Ϋ����uQ�o����Ʉ�
c>�7�w�ͱ��k���uvJwU�)��Ȝ�{�f�>�޳�G�I�o=�#���!�)��U�$�(.y��,kH�~��cB��3�+k����1z��SM�'37;+�]YH�-���7�j����mȏe7Y�	7o���#��[��edH,�U�:���Y��OH���U�a�Q�Sw�:����P�}ke���>wF��{���x�Y�l����!F>��ѷ7mη�w�� ��Tm���G�-�E�TR��X�h"��1FTYʊ*��ePDba-�\&1b"*�m"�2����a��V
֊���Ab1���YcX�k*.�b�QQqeB�KA��Xˆ�[h��#�B�ֱb
*���UFVUk*TL6a(��h#V$UF[E[j�(��T���"�����kP�dmkc[Z�aµZ�F�iT,b֍J�Z�b�Ѡ,[kJ!hT�UE�
����[J֥�-�,AaKQ�-j%�ATKq�.����`�6���Q�kR�VYm"���[a�Åb�mjҬ���K�(�յ`�-*b�&�R�%eF�"Z6ʷ�H���Im�h%��X,U%e�j��-�������0 �+..(�@��Z�n��٫Ȭ�}�����%頃�1�O\}���_E�٧c�g9� �7^J	�"���=L�JHt�>��fSj޷4ȷ?�v�v}����BWD��J��f���@
���IpȞ��<4�����;a� g�BX���gX.��%�>�P�(P�yi���=*#�VS;Vo/w�.����>�f_ެ�v�=��vZ3�0�U4��pr�OxT�Z��+����������M��e��RP��=�K�;�5�"��߄���Ԋ����S3}Dd�'ނs���k��qKϥn�t�z�*���}�zm���ܜ�߄���Ϧ�׾�8�p�Qw��b���gS�=�st�!}G��iǾ���[�q�OcӁ���գ���_��?K�y����f��}���n�f��Sv�,71.�l������9��?uI��Թ9k7���/����p�l����~���k�|.M�Y���z�a��!�+�{'#�}�^�qmm��q�p!�l��ų=rӝ1�=���7=u֫)v4$���j���s7*�W[�)����N��"��2�U���3ܡ9�p]c
����R5��E��p.n1`��7jo�)���)ue�tަ��#��ޖ�|�r�%6[��窶�RM���)����:w/E���.g_t��Hp�&�T�����O���d��1�����~.�nt��w��+U���Jw��N��z�v�����c��%��WXO�g94�w�]�?j���l�H�"����9��qn��]J=@tQ��������ǉ��3��o���xN�Os���yXwcg��(�����{A���t=Pkq��N2������Z������o�Ę%�do�4<�����}�w���6N�@�ڸ_g�s����Խ��*O3�>�̫>��U����l�.�W�C���V)��=W�ngs2���O�#(�h͡�󟖸Q�>�j]�	�z�'���P~ǟ{L���ޜ/���:�z�w��2�X�Iu<�ò�}��j�/�Fo�;�ݚ����I���MH�[��#>�uY�qތu��$g�$��|�%M��_���os5����wz8Ew]pR�����5�H�ΧX�)����<��h�����/+Gd��O%�������ֻ'���}�!��<��w\��g���/m�yU���KsH�\
U���ys4��Y��C�Ƕ��|��r�*I�;���헮X�7�����v�gU��8ɗ�7�l�!<}=:��Y��S�ܕ~�2����m����Od���>�2խN;���:��
X��Wس��SƮ:��,w�A��*��{�}θ]�ھ~3���
�_������+=�YR�~6�}[��p��*m��Kc2�oQ^��9�w@"�����d�Ϫ�Wi�`/S��˦�p��~*�����fD}yUIӎ��d2�rt���z����GN���������*���Wn�/�_�~ǥ��[�s��'u�غ��o�w���P���8�Ӧ�o\�)��{c�Ow��=�zf���-�W�b�iR�o<\���[�D���(�vٜ[��l��_\�*u�g��K��No��~mT��
?NY�3�5޺����y����8b����ݩ�^!O0|�s�ݤ*��;S{�����U�����~b�v)��ng�s�dU��YL^��R�u��ܥ���]����>�3њ���z�I2�����=|$��]�t;��i���
zԍ*|���ú�6�̼��{�G�ՙ����w՟<�aLò��4�u].�W�2l�j�#���]�[��\�^|�=�$�Lߔ�,;%}���>/eX���t_�������M�������m���WI)�����q�ͭ�÷(�,*��*�{gN�`K��z��̙����dㇹ�l������WL똷Nĥ�1���/=���~��@\�c;�;����qܘ����ڕ��m�\�!y�� �.Zte9���Q��b�r����{+�Ԕ�ʑ�hОw���9��n���y�މ���7����zdA����;]MK�VG��B�Xˬʑg������ϻ�W�z5�߽��#�	���/D���LlWr���ܝ�˪}�����9w����H�o�M���Xae�1�G ��o���^D�v�fH+�{�c/\.k�5'�M~�sf�uը�z?{(u��-�������F�BE�L�֘���fP �m��d���r����)�V�a��%�I��c����"w�Y�����o�"Z�=�<�L)e��J����"��I��EH��Ģt��R�Z�r�f��J�����W���l>���^X���ڝ�a�6pjs�o����n�Or�{d���z:+�u�^|�m��Mf����L啤��s�Ư�n�fg���=��B��]��裮ιhm�ڻ��V��b�Δ��Nݺ�olN�׻{.nՇ:��7�D 9����|X�oe����t|m�_���~o�w�K��2�Lݐ�����UvR�"��KQ�5Gί��E�3o4��6vI�%�=Z@��ւ���7��1#��ǰ��}��b�2���;Y�#���܅�$�wy��{n_k�:��N�G`J��ϗ��~w��d��N��V��yh�y�j�ɣ��Bnl����-{��t�kb��5�TߟnZ���(6G+�.�~cբټC`����f��;~:#>����<�h�P=x�̩�w8�߻|�����5lk����_�8��@0Ip΋�r���ׇw�LDy���r��(��u�b��s9ķ@�����4�q�u|m��Q�3����Ut͇_sY"ˢ>���r԰7 )��Wd�(����O<޼�O�mËƗ�zd�{f�/p��e�EB6X�}�3%�n؝���]}���'�c����ͷ���]M>������g���7��8���h�ؓݹ�櫙J�n�3���z���ɏ��Phz���lX�l�\����ٮw�fBJ��Z�W��9E�;��H��`OŬ��+����o�Ca����Ɵ{D�=�<A�S����<�=Ա��z�6����k]%��0��z;�a�3����ws�(*�z����>��D����Ņ�N���%��WXO��{�j�X��%0k�s}�zBdڎs����&����<w���d�Ǟ`�s���u-�Fe������t������u�l��x���w�����rIӴ��}�����\��5�o{2�}Yo��`��v�X�Q�/:��w��pe<���_gn��矄��Ϛ����7)����Chp�"�X�_c�/c��vjqB���1���\g*j����ɀ��j�u�Y��3����}�훪�yq�����z�>sf�>ƕ�xT%y9^����=��B�Ӱb�٢���=}�{cg��D��)�$�k��|�.�wC/x��k+ϚYP,���ϵ�5��Z��������I�w�]�M��Jssٙ��W�:�m͵.:'>�w,'��V���<�e�n�%W�z���8�ׯ�2w[tŉ�bC�e���2�=[W;�{�9�~A
�h��N�k��̟ٝ8�n1r=6:��˫�9�Z�m�c�n�zy��oA�/Ԟ���yS��ٮnqrcӀG鵵[�f�^��M�nl�MT��`)�.�}yQ׶�unK�_�f��ǻ,A|T��������ꮉ�,E�����,�]V�{��
�vr��س3�T������ֽ�ܗ7w���h_��Oƾ�lb�y��햺��8N�eo�Z�Yڟ)���&��G:T�ToF鮰�R��ly�>�|L�˷%����t��������ށ���������ϪE[��ntM���)*>]�e�>Ӿ��㜯&'��*$�kz5�]~�ϑ��ݓ�s2�>Y���j�7~�W�����\�Y�#qc�7c�x|���s��Z��u��Rn�����.͵rvu7ao��R�>ʶ��	f���!��k箛pWm�>87�z[ɻ����S=4���]Ɗ@l鸷9*�k�ﲧ�v{�w}�|f�����)y��?ng>�mk%��׽�8�y�X��D)�2R׫��ž��e���=����3<��";o�k�y�H秅o8>��}Zz��ٸ99枠�z�S��3�eJ*��n�r����)��9�����K�ON;�=W���0���_��ǳ �q�IZ.I��Kݒ��v�{)˭s����=&����K��6�����*b�/E��e�	��NJ~��T�]i���������7{F����ɠ<��!zl���UKʯ��v菳�0o;�6�Y%e������_\�c;�3�q��q�O>׃t�׵�[��-{&'[_e9ΏO8���uKo�>�zb=V�յ��f6������
t�
Ou%�é<��]-������HMh��.��B��mI��oO�U�]2q;cg�z����]�J�`v����ϧc��O�sϱj$����׳���i�"n�)�)mvZ��Mn��?Sm�~�������c�����]���;�b��n�l��Q�j���~���^`o�2��ѯ�����ň�v��t����r���un�L��8�xOle��,�޸��G;}�ɻ�;��aeh񵸆��O�����?|z��~�=�Q�=r�s�2gM~�lޅ��W�fm��$�nlvN�������Pm�k8Go��nl���O��֛������vݑjf^�X�0e/�N�<�Ş;�}y�c�"��|Ң���fէu~͒�;��s�n��]r�3�k�kb��;Sˌ��u�����pdv��)�����s���Xu�x˔B�v�>��J��ΛNaL��&v��ʞ���y��Ꞷ�gT���*���d 5�=�b,�;.w�}3\���������ݞ�꽳��I/FT��,GWO)�����ͭ򀸽IU�v�ލ���ڝ��w$�=8`yo�sR^ѻ��k:��*t�+N-��r�̉��+w�ͫk��=R<45^G����:�<K�mN��>� %��AA՗}��q]u76>�v���L+)=�eݜU*���y����@��F>���-�w;Y�G���S��\j{�3�����pw��ʁe�c�tm_˼��t��cφ����T��������S���>vo��u��e�xr_�;�`���o �ۊ6O3��P.�>��٥	�Мع1�扸��۽����AǶ���4��~SVћ��
�J��*�]�pW��2[�ߜݿ�{�ǰ�/.���c7l��Y14���ъ�w��]u�pen;��8���h�vĞ�w�yiM�������[��z�/���*��_��+\��r�q��;¤����a�?KX,�/d>5x�
��¯F/|zz�rp3p<�-GX��w�U��y�V�m��L�������Z��]Ew��y[�oK�=��n��բ����w�<�9�͗�t�����T��p�sr��r��W;�;�o8΀���X3��=�h:���BC^l�`��U��O����������Fo�%Z۞�u��V�P~�N�wݡ�i��j���/CUCтh����ڤrC�,�d��5N�DomS݄�D1�|�o�桼O�)ZF;�&��X`��s]	7%si6-�E��v�VP&	t��P��_I8�AI
o��[�\^¤ڮ��&�dV-b�c��ͩҷ��ټ��<�҄��'��x����e�q�fp�뾢$�5��RP<�[��8<�3-��ό�LwÐ:�!ޏ���>AǄ��S�na�݌��:��AW[GhԴ�v�.�=�(��e�?��n5B�Iϭ�)�UAe��e;�h�S��1b^_s���цq��굁oK��Ww�"܌1��p�E�vx,{�EF��0���ob�c5�!y�RBsx�r���x]龢,s�ݮ׫;Xݤ�i>U���R���WY[�����l3�4��S���G���5vo�Uy��{�G[���_*��s�D=w��r���P)n;H���5M���ْ�\����{��s�ͽУ��d��Ws[/Nhc���
0��$�%6�+�s1C��m*1\`�:�aa[�G,o�Nn��	��j��W���q�rm��JMv�"y��EeM�Ӆ�}~fｫ��6��$�
������6����a{s)�!��譝�͓ǖ.�7��=b��S��Cl�N]ׂ��Nu�u8��tu��x_^8Чo�1+(uZ�B�hu/���Ns�-�B(V��f�V�/;��)�ʊ�Q�)�'�F���-������.��g}�m�۠'�ZQ��0%�:<�w�5p7�ʹ�N�z��x屘��(��!j�Oδ&�G�fJyRO	��=�ʅ�et7��pʮ�B�y|�;��n�1sT��f⹧�c��l�аT���������7���
��v�|r;icV�)����;{����&��ڡ�CU}-<x����:�� �1�<&�5�R�,0t�rw9"W�a��<!��<��LӾ��my����fq,I��>��wL��w[B^s����cA�O�nd�N�� ~�Fei}�]�x�zV�[�h���0�OPCws:�7"�I]�q̉gM���/�:
e�Ś-�B�Z�lmr�]��i��-�#\�]��o��z���F���-�~��[�7����9t30�3�ӹt6
JeE׏i)�������K/\q�!���A�GH��)�t�eh8�t��{AV���f��\0V�B]� ��
M��O�AL�Sb1�@A�{,����W�s�=>��`����w������|/Tv���z`��}A匡Z�s��Z�}yE$ޝT&��Y�8:�]��7X;	�9ڢfG��s3+�A�YE�6)Ԗ�
.��	��yP��S��}�(���*��&-c�c�ZRa�[n�TY-�dE�Ym��0PhЭ
�2#�(��J%KZ��ڶ"���)�����*�Ų����m%V)km�ţ+
��mQ`�X(ơmZ(���V�Q#iQGmX�V�X����QE+E-�R���Vl�[X�����V%�,�؉K-mE��5F���hR��0�T-lE�	���Z�ԩYZ�ƍ����-j�QAb�
�Zŭ���b
X´d���@b�UkX��
��)Z����µ+RTVJ�UP\2��ԬmD���XJ�j�m�,XV�E"�%b��I��F
�H�Zԥ����@DbT-���
��"��X��(��[b�aR�*+,JZF��
���Ş��-ڎQ�����2G�}�������צ�����.�pj��¡O�sQ���jו���)��>z�;���O&�s�?����:�1Pє�%`9���U�3(��m�;���'V�ל[�ӥ	���^�ֺrr�qs�ۿ>�^��k�m�>����?ٗɿw�u���e6���^`�Eott�ʹ��ٓ��.|����:h�]�;lw9����zu'�zi"��<����3�k^@��`;%c3
�kW�����n�δ9�q���\����`�+�,�#ό����3�Y{+�W�Y�;��^jWZN�����9	�:IILX��$>��˘�U��Ԯ��T�z�ok�orZ�<�����cdzlt%�u�b��`ыB��c���^OS��e/w���ߦ�k�����Ǧ<��	`�q-_8/i�o�1z�	o�-��T�*q{�|��Ys�]Ѿ�P~�c�k�mQ/��؏���j2�%{۰.8\ر�MG��XH��6����U&��R���r�e:���A�G)�mn��l��OC������_kзhf�G��%�ub_y���o�S�We�v��E��l�1.�T�=MӼ�rK�%yu=N�>����^�vs��o���/����:�κ�����UiD1��^�v���ē�J�t3xDd�}���:�L��8�I������ǒs����(9�`Z���G�au�����ӽX�[?A��QΘ\��4�v9��.�W�_4P]&js�.�q���X�?|-�#����ێs~����\�o~�Eٽb׫q��Jn�D� �����s�tf��{�MK�^Q字JС!�5����n۵�w��D/���r�޽]����}����RzҨ=oŝl5{�cs<�s�W^��9�g�B��}Zz�6jV��^Yo$<&`�m��o#��r^���d�
`v��1fz^_>v�}Q����ޮ�鳢�~g�>}6d��>�����I3T���0gف�����^uϫb��	z�{�b��#�Z��J��͡�i�y�q��Y��j�&j�S����L��ԭ�iP���agr=:�o�o$��v��q��=��BcJ̏�[�daG8]����e�p��;e�,Z�{�H�N"������r�ҩ�I�PS�^��տ{ë��"�,H^�s�&\��^<:��a?K^��1ppyK����}��;�<�4�_���U��`�޻�Z}�k7y��˰�ۿ���
L�}V���gz�t���%N���l[:�㷝��wL�+�_�⽂/�������;^�Uqu<w��7�Q|<��y�~��t��}�>�\��?����m���;��LN�����߇)�8�1*n�������f�󝾷�r{������g��i���z$�ϻ�=���|�n�c���r�N]��#���do{4/(N��rcݫ'c}=���۵�j�s��ٷ�Zs�5'�M~�J�s&b�Y���<������a'Iz]1�/�����ۛ.}F�@v#��������7���t9�sz�>�i3_�p*�͓4ҽ�Z[��n\"�d;����'���}��]���2�s[�Zwv�3\�SΧ�'>LB�9U��6�x�f�k]��(h;#]��)r�o���M�q����w���t�6��ޣ+|w\G�]�W����+�����+)�q�lE�o$K�/D{oo'������������u�<Ό:��}[��1����ض�d�3|��<{�	�~��s����DG����@L�`yhI�M�Ϝ>�s|ǜ�<�t���{�\����Om�;C�d�O�m��Y��Ci=t�ٿ0q����ޤ�M l�q'S,�a�zw� x���}�I�39�IPP��ӭ��q�y^�w��&}��{�����J��T��d�tń�&��8�I��~�I]2��'O����2�4n�2q��;�I��&�Y��p�|�5��{��0k�����y~�[m�,��y�*T�oT�2�y�N�u���g��O=��I���RWL�CSz��	S�3��:�q�MX����p�޷�yUݦw�_�M�Oc���7��x��:sx	�4ə���,��=��T�&�My`T�d�����(M�:�Ohe�'��a�ֱ!�L����|E�~�gA���-J�\�V_W�5���M0�OwO4�����T8ɦL��T�2xw��e�u�3d�Y'u7�M�`xb�i&_S'�d�!�ha�G�GЏ��>�׿)�/w$��6?/�0�d��� (w���$��9���A`d�p��M2��y�'̞׾I0ɿ,��s�X�I���������Y��n�#������'�Up����Y�O�u'�{�&Y6��ox$�C:���y���J��{��N$�*�� i�L����m$�?{�V��¯�����	�Y��\}�?}���$�:b��I�f��M�<���񓌆O=ğ!�N ��k���9�:�2OY�)�M�Bs�bY5�'�y�g�}�߿�&�a�*]�A�,�Օ5^��k�W5��{��HX�Z�v��y�n�;ة
��*űM�o ���=�ڏ�Ir�Ȋ��ٛXQL�R>�����^��K�ݼ�.[�mq�.�����&�K��a�f�J*�R�����k�	������_�����e�i�I�O�Y�I�Vy�I�&]!�M��}��&��'Xzy��N��s��I�=�0u���Mk�9�xs�qo�v��w���c�lT~���f���: |��<��IY>`d�&��ğ33'��'S8��LyC�,�ϰd�&u�	Rm'YS<�q'X_;�����t��g7��=zz�4çq���}a=7�d�M;d�︓�'�f<ĕ �2�|ÈVC��&�A�a�i�|��I�d�V�<�Sx�7�y�|�L}��O�"��6ʝ����<�pu�I���Iēޖe��S���8�q=Ǹ���C�CL��`yl!�N&qL2M!����;��0|Sz�����;����2�d�{1C��J��{��'>���!Y8���pu�	�N�Τ�Ğ�rwn 6��y�a�i9�%I�CA/���?�<_$�J�<�l~���{���!�N'qd�I��͆��I֡�M�d>�0d�'~���������'Y2��h;I��;�$�x��=�����_kX�Bgv/���u���>DA:��+'PXyhI��ff
I��O3a�I�e2u�!���'|�b����/Ι2�ct�f�4��yڹ�7������������̋?}�羰,�hg��*
�"��VL�i&�i�0XM�u<͇Z�q�o�Ci4��ox8��O�!��i��������V��SkU�����L}�����5�	�&�w�`'P��&;�d�C<�$�XLj�aY4�������0�m�������L��L:I�3﫣��(��H����c��;?� ������I�ypx�Ě@��q
���Ag{d:�̚��|�u&y�IR����aY4���Y8ɦN�L��!�y��{Lo}�s��"˴w�~�@_X{V�eh��P��yI>V�:�Y]�sn���l)[�V�&�B��{jF�f�1�l�s���D5O����(!�/�,ʑ�#g�}͵�˥�_�j���â������/z��2�¶Vj��M��7m�yՅG:��!��qr�.�x��ֱ�IR����d��I��{aP�'�,����I�O��ɔ��9�%d�tn�d۔ ��uu)�+|�P��m��g��#��G����P�d<fY<d3���q��{�㬒�a�)�I_��N��
C��8��V7�Rz����&XO<��}��#���ۿG�}�����$��Y�`,:��OS���u��|�d�&�j{�3,�C{��!��0u�T�{�d�VC=��d�V��x2���},h���8����?���}�x�I�&�d�XM'M���$�31C�S,0Ì'�4�<d�N$��ؓHe�h>�k�OP��:�>A���8��G[��;��w���OR�;��4ɧI>7�@�&�3�}���8'�4���ń��L�3q�|�2ì8�}�$�
��|�Y8�k~���;ͧu�����g~=��O��pi�I=C�\��N0���d�&�Ry��O�|�ׄ�@�M5����>d�dŜd�%O&l8��w�Q�7����{�2y�s��or��8���sd�VfsX	ĝC&9���	���'XN���4���u��O�yd��`{5CIY<I�dŐ��2u=�;{��u�������u������q ��t�̜J�Ωd�Vt�� u����:�w�:������$��Nw�I�as�+��w�����n�L��nD�5�s_��	��gLRC�N&LS	&��0�X�q�iX�x"ì�~CӚąd����7�u&��m��ݸ�|�_�{�J��C��kS��O����|�~�~bJì��Ȥ��-!�d�g�	��L�P�<I6�d�!���d�'_���ąd��t�$�&����x�)7w߲��}Z�DOL\�^����]Mr�m�VZ��E��б��j�ӥ�z�TPq����7mo��u�i��V��{�b��8�X��L"A�r5����I���n�^�qI�I�um*�����e�8�Y�b*�5+�)1�g\ܼ��#��cڒ��_�8�ɖMr�i�2}�q
�4��<ĕ	�q
�H)=��q��FI��O�0�m���u�!���$���Y��`��Dڼ����ӣ>�Y�~�sx��&R{�bN�Y=I��}�&ٖL��x@��s�*
l��IY=P6Ì�LఇSXj�&���u}�iK�����ߝ:�ż�i���C�D��I��;�0zɤ�<��e��9�'S�M$��;�u�d�}���fs8����IY4�����&��z�J�~�m{�s��ӝ~}����a�H�3��J���=7�N2M=C��0e'Y'=���'i���qĚAf{��2gπ��I�)++	�o�Ǽ������|޽���%d���l�|N�XN�i<��_�N��_`��,3�ؒ,�o��a�I�{px���{�B�ĚAg;@=dν�~s�Y���|Ϟ���|�����);��%ea5�q"ɷ�1I�$��1d6��y3C/���qu�@�u����I+*O��ԁSÜ��N �9�s���0{�}��}��8�*2x�븐X|��{�XC~Y/�Iߦ�"ɧ�1a�Rz���P�'�u��I�w�&Y:�ٽ�&Ш{����_��bs~߳��y���{=AI*w\��N$��1=I�M%a��`�a�'����2O3�q%��y�E&_Y:�Ň'�S>��N0�����~�¾
~[�"ﭱ����=Bq'�/f��O�������3���8��l�؟$�&�=w i�L�;���$�?{�|�$�m	��O�R�߅c�E�����������������1�N�O>Ad���:�h/����9�u<d�gӜ��N2���8��M�I�` i'{�	=`|}���}�V;����^x���)�{���q�Wi�Ӎ���,���x2��yn���A�v9h%��M�%��5��$�����9���=�mZ�T<�:�Ekw�2�Uu&2a������T�7|h��.���՘
�T�\a���%F�����_|J٫�u�����|ɤ�LP�I�T�f�i��m��,�7� �d�T�y�Bq�X^S��@�\��'>����:ɷI>;�����T�pl��:Ӵ��}��Wœ��Ȳa��y�!�x��3�8�i
�L�m$��X�u	�b'8�9�	�ayN�d�a�cY;����>���9߽�����/�����$˖Oɭk�:�4��T�H}l4��L?ɊI��g�.'�u3<��	���m'YXOw�):��3ϱ!Y8ý�}j|mǺ����秝�����,�L;�u�	�u��z�ɐ��!�o6J�i�a���Aa�4�q�����bé�$�Xm&�Xh�6��>Ǿo���]k���C�dۦvk���C��i&;�u'Ι=I�w��q�=߾	&ٙ�1%@1�q
ɤZCHq��FI�g��־�F���k�ߋ�{�6t<M�M=���&��9�:���>;�@��g�`�ğ2e��=�x���w�L�d�~����*
���Aaߵ�������o��^�Z����$�'�$���4�I��6d��A�2q'��l�:ɦ=��I�M�|g����M��=︄�2�=���:�ߞ�<���\o�1��x}�=��{%ABi�J�l�:b�Ԛd�d�a8ɦy�k$�xo�Ci+�C;�'O���)�'�&���O|�ýĝL�m�y߻�����>�1�������x�<Is�d�!ӹĕ*I��*M2�zb���d���	�'����&�y�pI]2z������O�?J#��}�5��Y�%'U��I�{=����oL�z��︅C�M �<�u2gφY'X{�q%J�cW�+&��31I�M2u���	�����$���5�Az������t.��u�~����l:�ރ(Yn��a���flSM�<k�t/�e'q���0���TY/�R�sF�Yq̱�̆բWf ���mB��Մ����v���!з�Vt��}��������=��@�����m��5դ6�
�|a'#�=Ν{����=�m������d�+�{�i6�a2s�2��N��q�H,�y�'̞C���,��=�=ĕ��w;ċ&��<���&�z��a�N�������ʺ��.��� ��>�}�}����,�C�{�%eC�S�,�����q����z��4ʇyHT��k���,'��͒�d��X�I���vO߮�^�ƿ͋���������|~�4�t�>f�2É=��@�2�����C�k��$���`�'�3;�ORq&�P�7�@�&�2wy��ƪ�i���~D�hR�*zR��_�������I��L�f,:�i6̞��N!2�3�aԚ�ؓHe��/��I�C'9���$��r�d�T';�'�:ɭR;2}����_:���w���m��x�Ӝ��0�`z�ӄ�d�zb�z�)�Y�I�Ve���ݡ�'Y3��&��'P_O5��I�3�bu0���?$������.���?;?�������2q����g���M$����+&�5I���'��b��<d�gq�|ʙC�,���N �o`�'���"^h��Jwy�W�]�����~[/~=	��0��pi2�i���2q����pq��4���N��9ǘ��e��2�xÈVC��&��S�Hu(�����z��ߤ�T2����wG�:2q+����N��{�$+'Xxw�:�$�g1�Ԝ~a=�� q'Ι9�q'XN�͒��AC�VO�u
~�~��Q��p��?���~���ӌ�hq:ya��i�i��XOw�)8�ϨsVB�q����a<I����M�I�'�v�I�L�߾C�i�y�*M�.�k��c9��o���{���B�m�B�C��L��N$�g����nqC��}d2o2q��P��ąd��t퓬�d�{�4�'�<}'�}�������
Ŀ9�+���kf�FLa��wt�����������ħ� Oh಴ˁ����x�d�k�^T��
n�����2BlQ؞S�������{���>K-����3��9y�{9��Zrtz��'wa�����;�%���͛r>��s=�<]�\��VI�~s���1�:�d�i:����I6���f�i�	�T4��,��x�q��>v���4�x{��C�}�e��������g�E�{\|�4ϙ2�ǡ���I�L���:�{���6�!Y4�����M�3��'S��m�'�7�!��t��i~�x�;������,�w�Z�����{0��	����&Ri�s�2ɶ>v��2^��Y'��q%J�`5N0��J�P6����O,'4E�/����@������&3�-��Rs>�2�i�y�d�z����,:�9֘d�O�5��4����u�51��	ԙ9�IR��5x²i� e/������B��+��l�D�e~\�Mcz���L�m��x��&��sX�]����:�*Vs�:ì��l�N �4w��C��Ag{HT����}�e$�Nf�R��u~�o��9˜���;�};�~׸�_}�:E��1d�'z�0��!�a�'��CZ� i�d�C{�Y%J���0u�W���8����q
�4���H)=I�|}��u�g���vr��~��{=a<d�q%}I8�E'Ϩbì$��0��N2i�u�)8�����N���a6�a�k�:��*y�0u��Yy�����ɾ�X�ݹ�~�k�:a�L�a��*O�<;�u�'��߸����L�vE'��2��'�S�0�	�|�2u'zg�I���]Cﰁ����e��\��׫���ze���6ɴ��y��dӤ�s���M�w���'��>���&�:��XO_�e��d�%O��u�O �4�d}�,{�g~X��=�{Ve��sZq�0�>A�1	�N!�wY���9�u��Y�:ɷI<��'�>u���M i&�ɆN�d2ϙ<Mb�2O��apk�{���a��MgW��o!+W���	k�!=�u<sx�������FX�]��WH�a˽၀y�v�c����Ў�%A��\���F����͋���^)+ΘK�98�Gt���`5DY��<�^u�����iU�/�{42�{�g��sA6m�KҾ�uc���Y��t�/t���>��!��-Yܽ��w���ɗr����O�d�7 ��S�Ov����B��[�k9ڜ2�dD�-�V�;6���&�ӽ�����#Z���v�2:��`��X5F�ۜ�dg\���D��������/�g=�7��ffz�x�7�z�8��:��4b���ʺ|�_%FxV���7h14E;f�rI�p ��e]�Q��?[\%el��R�$� �Y��/�1�G>�ÊYsP���%**�i�טo�>H;�HuK4��=Q���G���Z7�_=y�K�H�> �c[���F��j4����~+�2�#Ќ}i'O�j��e�;9���>��v�IR5u���EXdor�G�M�I5�(����-��:�b�W�M��W]s�ie4"rN��.�����P����ge��4	���8V.�I�_=����J������()˪�:id�k�>�n�BCU}c~���K�������]�1��������v��� ��{����@�D��}�t�.S���*)*pV)�u�x��He��i������nN���2g:�D(~1��\5=�Κ���@�UrW,�,�{$&	����:��.��E`���ݽl�l7�/Y���6�m�ԣ���[Rny>2xO_���.-�Uv�}���B0-Y�hV��ۀՇ)��{{�Z���VA��լ�y�gKsZ�&e
�%��Ԅ�����O��8;��mYk$�;�a�鮰vԾ$O�F�l+wn�f��v���h=�z�[b���ork����wHn�(vr���I�ɾ�挮wr��$�y�y�x*�ֵ�Ō��|#	�HD0݊Rc������������\h_nH�I�p�;��<S���w��K�*�=�!�*3�q�"؝��ǻTɅIY.��W��ėou�U��Ŷ/l�I��7u}9�mh��.M]�K�S�j���P��c���aMz���j����
�Y]��܆��KOv�gV�'@G�B�壴)���6x���kY]ǽ]豝=�Sۺ!P����%ld��#l�r�V)��h���]^�Q�r�b��H<��$k:{ȯL��� }S���fs������Wxu����
��Ҝ�jC9�w2,9��@^[���S��ǞOZ�����eثۭ�1��ʸg]�K�-��YL�6.���44�=�J��A7|c�45g*e�}/DY �[&[��%�f)Y�z���밁�����B;�����e,tiD�|Po���"��2�:G��g9I���P��(VJʂ�l[dUX��[E�ZV�J�Z

V4��-T��REZԬ��T�
��U[E�Z�)R�"���b�2VTlh��҉+QmKDPm�U*(Jԕ
��"��+-��-�����h#B�`�PmȲU��l��e��PF*
"���TRTY�+Z��j"J*m%-[m*�@�E�`�X�ʬU�U��T�ր�����R�E��(#R*��U��[+ZP�+Z�"��"(�Qk�km@��Q��jA�-Dd��R�TiXa+j2��Ԥ���,X("[d��T
2V
(�R���eh�,`,R�����*� �TYPYFJ�X,
��)+%aZ�(��U�B��������@�6QH�IZ�AE�%!m�J��@��A�_�$��脂WK��㨑��J�ci��e��W`۞�h�7wxG��{�M��PL%��6,k1�ՙC��W���Mz�?W��k��AI?]�!�� �g�bM!�}G����S��k�����L��Vr��.x>���鸡�g��l];�O�z
�V�9����'�i~���M�=~���մ]�D�,�_�k�%��A���5�1���l���߅m�͜x>�ھ��T�b�xiр�v�����no���L�|������'�*M���xzâ�Ί:���:����gny�>���:�O��ޔS̓gK����rL�g]�<e�(�gN.}j�OrL=�ý���y��*��˭2>�m�Ω+j\���d-gH�����R���Nqw��}��%�������*��=�%�ϪOZ�'�&�ɰ��;�_o�H�x]�������P7.>���$/DK�q֠��I���k<��"/Q�������j�o�w:VfK���>��!wR����TPc6�f� �X�_�Λ���?*�`���Q�K�K͜��λ��8%��Ĝ]ab�;�7�R�a7���K�;��F��n���z^	�_]L��(0�1)�Ư�뇶�<2{�
���eH�,�t�K�k]nWuf�={�/���S=m�g�If�t;��1�e�WA<��*=��'ɿ>���î���w_M��z_�ݯJ�N��lX���3�sj�;3��S=yo����G�h]'6U;�=pgv�pf�����ӕ����YW,�P���ّF�������'��b���n6�f��ny�k9���qf!��߳ޗ�o[5����z]��rW��Ł��V�a9y���k��/zX~~3�.�ۙ�!�Sug �k��38��B�A}�ٷ�XNt��7z�]~p]����[��'���">ʢ���쪾���Wp���+�auEH�I���i�_�s� Xz�Ӣ��ik��ܳQ�FצuL��J��0}���Ϝ��){�Ӧ�sKw𝋬J=E���:Iԟ[��~����fɮ�tum�y|���ӺX��멮�w{<e�(��^. oڔ�3n���_1.�������3<���z`E�d�<�ǓJ�;[�������L���{�[H�t�/�p�\{
'6�����Ld�ޗ5/RMK�Ǜ��	r�]��h���e�w�\|01&�ǜ���{NW����:��>�M�a���#���u{=g��x:�bN�O�z�zk�F̜�9b����xrn�.d)��s���u�g�{��լ�}�y��~�a�6zSۢ�CS�`@��gKʾwZ�����;�AW��u���.�;��w�Y�sx,�I3�)w1�:�Y{+��W����0���jJ�1��=�9	��Er[��&\�������J��'0����`����%���Wp���|�X����sw�9n��S�t�w/H�X�@rݻt/��g���N����lI;�}����
��Z�Re=N��	��V�-ת[g��u��{ҝ��':����p(-��3���Z|�_VK�Ꞓc��p�N���NU�]^גU�Ό���.�����_n��+��3��y�?6-g�_��Y�~��W�5�c��9�U��rȽԽ���4��5db�قZ��X[���4��q���Y�e��'l%أ�y�I�[�V+�Re.R�����Z��d�X�6��͙��}sN��6�!9vM�L�<���+Ϭ).�ԆE����{i
���}��|u2�$�d�?�t����'^�'L�R���P��y�k@ɥd�=��_�T�s�{���c~�o�3?_G:3w�~�2FGN�YK�4�CW��u�����|�t�>5�#�=.���ޜ�z3�M2��ۦ�3�Z��O�'�u�K���u�ܛ��c����^�<im�Yy�t���u���U���\Ί���@_S��,r�z�厜Ȧ���6���YW��۟\o+���LQ�3���փ�|Z���ۙ-�F�������}|��N.��){�K�+T���+�gM.�W�=�,Wu�Ͳ7+̛���Vw|���̕q�B�.�+�I0EQ��5�2ǚ���w����I��e��vڞTu3�i�|"�/��!�&\��J���WW��Ѐ�U��7�/J=��%��>�t��oZ* �e�uk��� NZo����r���0�V�%�8*�:�W����ޔ��vq4@�2!�|ZY-�����dr�_v�{-N^�6ю��t˺�կln�����C�E����:�˭b�Ǫ�o:����I�Ͼ���J���nȈ^��������Rg�?_�v�Y�=|��5e����e�n�E��y���'p���bu�NV�z�'�)��Q��m����*�5b���׶��A�G�y�lOc�sw��W��g��	�и��<����zH����zrr�q��s����䛻�M�f�Ǿ�nQ�X}�;<�o�Q������ßV�`'-���s|�ɻ�U��Ƚ{�N^�Μ�v��x|��uu��Wk��86m��Nt�ԞϦ��~z�F/����0����_J6"��'���|NCz���o&�������Fr�ѷ�����:m�غ���E��K�Ԯ���ssd�yݲ��{�u��]��>���{�vu�!gEr�C��n�0�{t�1-Ԫc68ͷ����_���x�2�L�'��D.gI��qYy���>ö�crcN
�I�s%e)�o������F�՘D��Jz�2K{�ў�T�^&zעe�����'7f0��xj�F�Z��NoC�{���n�K�=-Kݸ��5�	��8���"�̃�w�t����Mt��D
��WsV�-3OoM���ﾪ���N��O�P���C(�k2cbVk}/x\�՟L�j`w�=}6��j��;��f�B��ꂦ�2���;�lJ���=�$��>�<RN�m,��~�׷�Hd�l��gM6R{�u�ݏ{��2<S���V��J��p�ڹ�5BsL�����km|{;��}fd���+���z�Rz7{�9�;�̿�=Re�󭭋��.R|���ˇg���oop�W#��~�N7�_c�\���sD���6���2�bU�m��^�׻0ܝN�;{>��0{=|0wl�h{�����s_��kQ��i��x�«��鋺nj�/k���/�Ŋ�F0V㿛��������穉g�*{���������z�O���Ŏ��V�\����5�;�1Ӭ����b�M�{��B����`O�}l/�d;ųa�P���8�t�>���T}"�42�X�V ��w��� �5:1G���"ұ���p�`��x�Xv�Kf�E*%�/j�j��S�f)��ec#�nb� �޻�]�t��]��q��v���NAҰY;���F6�VV�-��Wo�s�� � ���o�x���y�?k6i��O���[/�c��n��n��B`��t>6ˎN��S��y��wb��pe*�r�,j��V�O3z��fqɳ�s;j���Ż�u�G�:)�A���i�7f�sm��W�����������멮�q��0�Qo{sҲ���k~$N�b���:U�t/g�Ou�����������	�/c�����~�y�+�كg���t�\��{W��h���^�N��k�@A�a�ٝ-9���� ��}Nz԰��+�gIs��ըG�&%~ˊ]�c�E?R1����ݟ5Op	h���j]���+Y캣��iA\��ƥ�~�n�˙',���:�u�_7"�-����g�]K���{[$���pc���=���ߠ������ngt&���q�cӃe9�J�T��pzS����˳�[��3��-�ɟ6S!������)�Y9����a^}��w���m0[ߵ���^Ύ=�xP>o/�H�S��ԝj�̜����K�Ų�s�l�JK/	���c��Z�vz�d�N�93�!xB�jcIR���K�[NWﾯ���%�����-��d�//�U�[Ͻ��3�e���6����;�����<B�oy��'V\��k��m�}�GʛR'��V_{�y�[�y�O��dJ,��]=魵U:L��(�3~�v`�zr���y%lx��~J��uڛ�Oo�;�=Nw?>�]�g�{<��lZ�*�:ž��`�Uk`Q�%9}~�	19��޹i˙�?g�9�.g*7@w�;�z���Wz��^�[t:V��m� ��o����*9ј�~�s�`X]�J�<��0^��ה�П�>���UJ�	񯳄~ǥ�ɵq�~�szR�s��ze�y��v���\�B/��H��Rբo����MT���ψ^�R�{m�{�Co�Pt뽞=a����pC�}|���z{�V�F��<��~�/ �滟[�*�VɂJ#3��>��r��kU�.�<0���m �}u*�Oj����ow�d_wk�`��<�E��3�ޙs���D���-�v<t�x�� $��߁�ug�{���dBQy2�>Yn�Y���B����yg5E����r�[�͓�m�-���Y�lV��V�N��ZRo��/=WK���^*��������x��4��]ޞ�����侪��|���Κ�We��<�ښ�'9���C�-�����ϥ\p���rM���z�d�[c'e�rd$%(��f��>����d�G�*b���C�����u�s�o�$�J�T��{-�-F��VL��Кp�3>ѻ�-?r�¯�m~�+�A!+%5%�o���)ڪ;-�κ���Z��y� .�}��\^V3�Ȏ>�پx��sf���|/���yn��X_���mԳ!x��[����)�������9��r4�<�Զ���,Z���ʃodi�9^=8uoB�_�n3s�v�{��	7wJ�`�����'��}ܚ~=�V�5�Ak:z�Ov�ײt�r�g�{_�hÛ��R�kh���`/V��q�l*��Ϳ8\��5'�@���jn�WUj��,5ջ��^:U��eK�<�Z�鹚��jnJ�:p\��Oג��Y�˥6�t�a��k�.�]��Δ۹��~���e�q���#k/��Mq7��s��9��T���(r2��CO�v�9i�Sʌ36X)'��s�>���|�tK��r����w�qa�N�]L��U�4;�?g��w!v�>+�==-��N��o�ײ'����b�b_��V�>&v_�a�c��n���Oc��l2�oU�Sۘ3�k�����u�C�Frx�>�V���S�ߡ�Fe���N��t��~��]tλ�O�pbҏ��xk�5�N��gz��������:n5'�����^ԕ���S�X�[����pN�#�y����)�������;075�Ү<S�%o�X�A���n�[�qiO7��>7�؀����d^�ؾ����X�]����b��1�8�y�˿g7f�A�����S.c�e}ò��Y�[�{[~�4C�-x����^8���7��l\���z�˘������lL�(g��vg��]$me��zm�����8�&=1���WÎ��Ͼ�xؿ�V��;%غJ�9�J����N���,����{�<J�;*��N���Ot���<5�6���xv:夵��$��-����}Z;���{�<��efr�I�<����um�'��+��.��_;n�X�
�O���C;2!=^!g�d���K]�K�M�eJ��7t��K���T��3��eq��j2� �aYC�;���֐����85�ƨ�8�{NL�`0�u:���V�;�y�+�`E|0�G�ws{,�|����Y�0x�e2�G���K{ާ)h�I��U^�GG\�Vu��H��B��oc��+�\7/):t��}��s�
�}ջn�;�;+�ɡ����1�G�p�/���y��:�\8fA�3N�I�
|����-���o�b�Mܴ/�a#;�-]AVE#G�3&hm��LVN0�5e��vL�2I�&��|ڠk�-a��ftھx�^B)�)���Jڔrt=\����m�pt��2�<U ߌd��B\����4�A�z�>���W���L�S8b������{��qu�v��r���r�ߧ�Snk���έGt��-�,��7q̛ͪǆJ6���oL�%ej�!y�WI�\F돚� ���`�'<=�����p���5�P&�҅(���6K���a�u��B�'�f֏uZ��$��7Sw^��OC�l٪rz�z����Y��ƕ#�.	pU�4{�<��u���=�|Ӡ1�9b�\�{#Ohhpu��˜#�ٙ�.���s���/ﵭUë�]�#n��$�\�bӭv���6?OG��҂���&�/QW��'e�d�W���	�\wOA���h
9F��T�YXy���ɧ��U�]�S*�KJĈ��c02*L줸�9%٠\`L��:�W_��`wk�Bv3`��k��i��,�P��s7u�������K,[��/M놭Ɖ|�FvRsѱ�́��U�5�ջ���2�a��n%��^[���������ʽ�v�ݏ��5��u��˷z/'q�:��|e���G1�
�xvq&u�n� �>�LM�T&�����N�b!����׸��{���)-��j�f�ud�� 1����\�Tx��w[w)d�G���qI�.7&��2�н�����]��K/C�n:}�u�_v>�&���?���6&W��8���=yǋ����<�r՝;���mP��(�D�T��c!�H��/��nѫ�_)9�'�\���C:���R���6�F!��]HΠ�R���b�&M"��!�7b�Ȋ�[1V�5q�sM>�2�/)j�Ouw�e']J<F��v{��/1��i�oB��D9���&s��v�Qpb;�]-&��N><���WG�P�j�A]:W��^�V���%(`�wA���olX��l�%|L'2�u�k��
5�f���k�ݞ�?_�m*��lZ�,[h¤���B�E#j��-����ch��YY)l�#"�Ņ`("ڠ6�[lRڰi[(5�*("�kTZֈ�mcl�ԋ`�+KDKK��X%��AkijJ�B�PkdZ�J,�b���jVE�T
�-�E%`�b��jUKJ6��J�jŕ��k-�kE��P�Y)lUj��eVV�%V�T+"����"�����mUF�ԋ���Ab���)�j�*T����,��Q����A`�R�Ym"��(���%�lYU#ibVT��ڲ-���)Z�����YQTF�����J!R�j,P���DZ�Kh)b��������
Ʋ�iX�@D�#i%��J�Q�����`)*J%�U�%��j ��bԩX4�kd��,*��-��Z�>�	W�u�;�y[.��ܕ�\�ޤ{Y�/�euY�b.�\��h@s��'7--�a���W�k�����|>T����Ϗ^ ����/*��z����Oy������-W��-�
=g40�v:>U�fy�˕~�.�ь��/�<�6'��7x�bW�Xۢ�Ǻ->�2�]ɽz�M;�i���B�����
��}��	��K��%yfO�wn:�s2��`6ת_��2�Ac�[#K#Ϊ2a�>z�;�����R{�{޹=aY���ʹ�K�}}Pk�iw�Tz���޾�vY���������59�Ӟ���v|��X}��xn��P�%��i~�>��+�o��Βo�3��G9��N-�ӱu�(��}��=�<~�lq�>2q�.��ɹ�N�`Os���yX�9L�oW�^8��ю��dzW!Fpʿ�N�F��U��*�u��sY�ÙX�죾�{[޺��nĞĲ:;Ft�\����7'(3�}�:�Kk��/�o�1o������{a�6%�+��ՙ)#���H�u��4l}�j/R��.^Pn�=˧"�>����8�wO�����O>�&+=>j�B1���������T�4�BƥU��{���}gvtI����v�[Q�yq��������˹[rn˔Uw���^�r�`�=jXv������{C<{t5��^�t�Hv���2���EOpHkE�$�R�`xJ�{/��WJ�]b*�biTŮ����K��|�;��	�܊Ėă�d�ԗ�u���ͻγl������Om�����ǔ�V\��ng�К�AwN�W�_`��䒛p�׽r��Ww�����A9���q�ϕ;��r�T��c\��|�Fu]���8�^=��Y������8��/e��~�3���[�/{ϟ����x���z7F�O����M�G�w�~U8,밟�}q���P�?X��#�=�I?*l���n5�}�k=�6UOL�d�����OS>���Vֽc���<�=J&��8��s2uKz�0�z{!�
�xo����u�>)�{ޭ~|�6w���3>�d��2M�Q-��(��!1�oV������%r��0*uEf}|�����J$wf)Kgl�me��$C٣�����Bm�w)�k��6EF u�g�P84��{ԛ=��-�;{w�~��㾩Jd���oDs�]t��HU�P^���u����=U��x�mb��,I��E�-4��7E�x.���پ�J2�\���4���tE�H}F��v";��k��%	μu��n��U���չh�g�nYuСZ �r���������s,�J~X�\#�����,��x+�ܯ91<�f|.N�hu.��G�ݠEF�O5=�C�����}]S�
�E*����L�ɖ�s�9��+�7�����j��Kg1LD�ba�hs�I�Gօ�ǣ���\�M�j͊��n�R�עU��p�^Z�L]~28*`�e���R���q��]y�vk��Ϭ�K�.f��;��0�'/&Pc$G�*���4ڗ^��U�j���d�8����vK^$��DFmr�K�pЃ��ua��Iw�E��$�F�n������n��y%(����\~$��:�^Z/���pߴ��2�ŵ���@�-����;�1fLR[����p� �@��{�6�bt���������^��W���M�n>� V>���MzQ��|
>���Բ;DU{&JbVط]5�"\/�����I�����e�گ^�z{��C�ZiWu��lu^��O�������[��B-��ఌ�ޅ�B�e.u�J�2�sޙ�����C��<�;foc�!�r��?(��섯�[�Yʏn�涳v�MٟL��u�J�A`8D���z����Y��>|�ss)�:teS\���ly�`8q���[=�P���ܴ!n�ϵ^��U��v���3Ϲ�6�}Zsj�;~�"���`�3�Bҹ�p�+{Zw��:X�;+qq��H�y�ꛗ��a��IX�'N����{|a'>��fS�����^0��Q���'p�BD~��V_����o=cz�f�����ҩ,�v���#|Sip{W=���X��r���N���oA�;� �kڡ���Yk����6�N�*3�4���^s+sޣus�=Y �H�Z5v!���fiYg��m�sdpgB��̑[�y*�.�K=����O)��8f�����1Ͳ �{��Z}ᷱ�.�����q���6�No	ꃣo�1e�H9]s�UF���COs��qB�u�����O4hr�s=�?�F��٭��I���bX�\[X(&E_���}�@���cȯK���Bx��h÷�םI��\4��N�@В��].^�~��ʲ='�</L���-��T�N:Ш���"�#�hW<8F����.�J]*�˕�Lhu�7��^W����A��۫C�[���g�B�P���@��,kj⎯:m��c���5_g�CĞ]��ms�2���N�eI�) �˫��j]����Sg�ͷ��]g7�cO�>���]���X�+�2�C�<����I.Z<�~�L<'ۈlR�9��X%�I�E>���<�='���o!3O�τ�ܪ"xM	c�w��|�7���Յb���>�M����2荀90%zd��}��?%����ף��kЉ�����)��{dz{�ڞz	O���0L��^���ƥ�
��������bw�,��0�C��w�u��&��7�F�B�q�+��ݳ=����n��pP��|���Z���׎g�$}�gtͥ��7�7��j;��k��[\2b|Dv�{�-P{��d{<�2�^�B�Ȟe��3������s�G��X��F�XxS+ސ�uY`�jq&/m��k����a�Ŧ�;��K9�:�� ]���=P�zg���q�Ք��-^!}[.hN�������H�]ӭF��%3�T<e��9C�K3z�����²��kM1�x{l�AV��^��([�&7:�h�g�L�bk {��`��:��zq�O~�K��օ��,�9z�oI�Z��e˳�W��W�����㭋�</�圍�6�cX3}��ۨ�i�X��/A;�K���^�݈��#)iƛ�j����k�-봁#c��F�j�uvI�6K���m�q� �b�����]�o�⤘R���C�M�p�?�����/vO>�N���k�ª�^}uD4��x���N��>�8\\ק���h�|:����Y�S��G�)��F��<�A31��C�N���kG�޽����ь?'�R���*юj�q#ԧ��$u�v��ɥ��]L�3r�R�W�c�����?z�N���oK��G5�B2���n���坧~��� ��y-��r	�ѕ����]^&<�+3����*+��
�t�j=r�ܩ�K9�HC]-*�'f�et+�<֬��Y��8�05�Z���F�"�]�^�՞0��*fa��H�őرO�K���l��x߹ٴs�PZ��ٹ�;��lwL	+��
��`ȓZ;�-"]T>����5RN';G�{��g����F�h���^�P�s�ZK\�%��%�N�t5(<����nq:,��[�6���{~�dx�%W��#�<[x��\t����Q�Me8�����G0�'����n��^ܥ�a{VeKlb���R�`�,m�Oً$�۞�ڇOOm�� ��~�u�U]���0�}]��VT�Z�%�;3�}��{���%�9w-w��}}QA�]vg2nf0-_<���ύux�W+�=���>��i��)����x�ETcuԻ�v�I���<���{�]~��/9+>���dN����AF5B��>Ͼ���srx�/ʎ�m�97�7W��=�������xbX��K�e�F�u=��<�J���_���9Z���r����Ե�Փ]�7�/N��:���5c-'�3���:�h��Z<y�io3�n��Iw ����$�\��r�R��8'�-�l^Ǿ�q�~×�5Bu��/5jpUq��\^ܲh_T$�"[+�Ҋ�Nj[�킙�Lb��z�:���G�g�����IP��s������.�Q{UFǘ����"�?N�����\Mݼ�<�ܓ_b�+`Y�u�]���5�M-�Kb�J���v�Q<ZK�z�R�zh����wx�r��j�bS��a�G~ζF�lХC�e�\�ϨP�y}i�'��<&�{6L��vH��jR��ߥ_'<�<2K�Wr��S0��D�:D�q}�b�Ìӛ%ou����B�r��5��u;�^�W�Ay8����L�T�p�)�ʥ�*�>��n���gK,�!��lK;��x.,�X%���:$G�*ES�{�^�ז^LO��bտm�N�F͹mS�g&,�E�rġ�+9�.�/wu���"%b�7����_v��R�''�ȑx����L��M,7�����X��34\7}_�/�mԹGa�1T�B�*��8<�3U��Jip��{2L�������'���7��M8?+"$��"6��yh��ᮍ�c}gV�w�%fEȮ�=�*�E�`x߿��R"��/+��ك��~�����=e���^_��UL������f���8��wgU��
�}<��B�����|���[��}�͚�[K,�\�//��:���ܞ�˯6{Y�ִo;����**�\�Ϣ��,�"��L���릡x�<'����3�o@̨�����!>��C�_�qp��E�J{���M�����ѣӖ�<��	��ޮ�雍�d��{y��}�<�}UJ��L��6���ZChsI˱�:��`O;��n>�<.�\�ؚ�˻��B�=3�����|���|�`/����#~{|a%jf'*�@Թ�4w*�p���WAGm_��w����^VGQX��S*_c)�B��H�MH�6������V^k���b�v���/�O�S�S��N ˥~:h`5���{�U*3��M }��/�z��,W>�tS=�l�e��a��v3�ƽ�>}����f��\��;H�j�5c�ˎ�H���}��Sb�;�05����j����
r]%���G����@�km1�`��s5����gh"m�N�Iؚ�N��֡w���ȕؙ�~�t�%�-
�k}����Hx	}%�Κr���|T�t�lb*��W/=�a�|��U=��_����|�<P-��w�����V<��o����=���+{��3�2�g��&����%yސYU�dz���e�A�u �N�˒m?'��P؞益�]p���I�P�w^Gd����TΌ3C:LJ���O�u��M(g�1/��}+9\RУٵ�LT��.�K�P��o���ϕ�:�U����ȍ%����S~��@r��I�+O�9��k���R�h�m�Nf���9�u-[�E�b����B���\e��p��Vjgm��	$�׺*�P�<9n�L:ѹ���g�U�N	>G �!ؑ��Ж8Wy_ԟ-��f��4D������e>Seq��W����+,�COR�D�ea�|8���ީ�w�b�7�r�y�I�ݓ��{��q��y�Wb�t��`��c�d �xa��Y&���'���+o�8���ݒ(���,�s�>�sj������u�^�,{ٍ,�ml\�єī�������fN'Bq��^5���G�m:��c��������uO]�J��f�����E!{�o��������o�F��h�ُF�3�G�-v�B�9�C�n�
;F���l?o�)�7�ܯ*0kɻ(JU��UΤҩ{5D��
����I����^��c;�xܩ�ݧB��Ec �����u�m�9��\�u�f>]�?����}��c�w��$��`��;��NF�MOja�t�$t����{�����I�}�C���s9�r���݆��]��r���5��.���$b4��>�U�(J��76HjH�n^1-�����'C\b��̱N�(|�X��7����p�
�G�Ҵͪ�L�ܯ�1�ȴo��w�oS��\�ZbU�E����7���=�f�V�k|8?���V���v8��u^�"U�$�u�![�`�qM^�J+ϲ�5�8�f���q]���干�*����>�2���L�uE�:��nmlC���ɍ��s��.�2N��'8b�w�=kb$M�]�k�M-�S/
f^SJz�h�=���3���r��r��_I�#�f�k�c��o���Ȱ"Я%�R��Z�C��\�ͮ�Ӭ[����q���fi�T��������%��HZ�iH���9z�
eOne�s۔�uᜠ��9W,},#>�� ����$5g�;b�f|� �6���m� O�.½�����:�51�槃�I�hˣ�j�~�J^��	9�C�g.P:T{�<Yd��.cf>nu�<
��'M˵޵(��:�����]%j8FhG��E�.��0L�ӄ��T{��G	�ؔ���'0mևW���b��ܣ��钴f�Cщ>o&[�)��#�Kk8�umN!f�B|J�Q�q�s��I=g��U�ho��^)j�(>��=���@dY{�����>	��޻�����')���=�1[֯w������Mm	BT�h�t����m�F��\{����kZ�*Rc#:5s�u���np�Z,�Ԋ˅�ՙ�U7�K5:f��(����=������;9܊st�]F?{����
������~�s���ܬ̣�m�kwi�n�AЎ$T�q�H˒WƬ=�5���n���g-g�ǝҢ���J̻��xsu�j�l��;��͔�b��ʔ:U�L�%�j���ܛa�:D��M�/V>+��k�U�pŞݮ�B�L�i�O*�Sy;���YL�C�$-�9���|��]˶�Ѧd�ä��}����v/��0��z��*�`0Ǚܥ3��]M�٪�V-���Ư�K�ʄe`������'@.����8ͶM��A����ulZQ[mW\� 3Y��p�#����M(�.����{�~��J���:�x���C��\�q�S1��	'n���l�}�и�]u˹��X��m~#Æ�R�G�=�r��#������[̣�����q!X�����{�f�������0����N��!]]�oU�}�PT�R��;I�,�(�Xy��K�SXs��آ�F�66Qc�"�mZ��O
���[��)�bkB>�;��2<�� �P.���˛s�z z��t.V�w+��V�L*U��L�sa�iu�R������o���a��5K�����t�#�X��;@5��˒[�h���
��W��i��sh�M\�k{�kHP���y� �gb���n�s��s�Q&�}F?u��[�fXF��gX4	�ݻb��<T��1wM�%�x�L���D�j�w,�װz�m$���� �b���]�����w���_es�N���m�`�;9��v��:C�h�|Vž����k�̥j���9��DKWcJ#��s�Ϻ0I�E���uF�uS�p;�w��i
�1�����2�P��c���ak��3ܨ��Os���RjV�6�2�4N��[Lw9�rWb��ᇘ�w�=wr�����Jԩ8�V�w���.�t�矀0ٚ����"ѡ�l�/�ãqXı�e��j�^��l!,���m{��I�h;����t�]�gĆ�:Ƙ�'r��f�/'6�X}ù	}%�O�����>Yd2��cmE
�ZQe�TE�R��-�bF�h�5X��,X
�XUih��X(�0�b �%�YREPm�,DYY#h����U���*(,�m" �KJ����l�-�X1�
(E
�R*��,YZ��T-�Z�lU�������U�(����[E��X����*��[eQ��
���YFV��Q��
�ŁP�+6±* ,++AjJ���
�RT*#"��EV"���Q��6��QV��!R�(,�A��6֫kU�E�(�b1��R1X���PP�U,�QUH��*B�X(�X��b�T����*�b�VT-�Qb�T�`�ְU�QT�,R�)5D� 6�IK)N)$�Z���dM;�����x���>C!Sf[C׵3�����=+�3��O�ܽ��}�Q@����>�*��l���"�R���\z���/�wY�3��%bJ�+�L��5���Z:}A �鯷:�f�)bb�0��
��k6��n�<-�I&5�aX���Ԯo��)�\�,����ŉO�J:�w�,�K�Nyp�K(p�v����t`�3s�mP��3=�a*k�I9�+��r������0��0
�8�+j��"����-t�](�=�9yS:)��ώ|�u�2�6g�N�u��������K����4���nS{і<D�=��9�Cbc�2��^!�����F���6W�� �
�s��"!�,�K����ko��l�g��3�
� =䚋���W�9����^3�˄z�c>'`k��G�y������i�����ꄛ�Kec�Q\S��Է�_��&W`��Ȗ�u�ء�>��JU a9�kS>Eh���c�R^�C��\��"9��mp
�ޖ=���}^����8�����<TG	4�	lS)-*��xO��YX\x�]:&�ۨ�<T�}�[Y`�"<w�[	��9V]:�}3V����*�7�U��4�w
̣�3x��	p�}�����N�gӎ�l�K�6�鴊��j��y)!YZ�V�����P�ŜL�*�r���j��R0$J�߽���@�O������|>�lc!�*l�V27��,�y<��sP�]u0��M��C��`	sS
�T��E��^�f���d;�VS^��p��*���I��������`S0�(��s�I����ҝ_S��{u��ѽx��"��A��[�:�î*�A��^�T��2�§���"���+�܏�q�E#;�4��D�����c}|���v,���WcN	)Z��k�n���c��垓�^��
��)%�#ؼJ�*�.�;-,efk$��NP8(L~�ݩ�Ru�{';7~ґib��lD�u��yh����e�\/Nb�Ɋ�;NtN�/{q�EA��J<[D��$�D�V/r� �
�$�9�.�!��}�]w%�v�:�eH�2�;S��SΙ�����dv��V	�n�},'z�X����o�*K�����9��6�3��[�}{c�cP��[K�[=��CǍ�\h�|�ЛB�^t*J�Լ������ta9W63n�9~�!��9��3���3��ee$ũ�q]��wVc�a�
�[f���.���
�>�y��U��Dbm����:��޾H�M�՜�",��<C�I!����W����W⻤7�C�#eC'���!֤�uUgu�ڬ1�E&����(�W��y�$5��Y���������*�qd���c�>����-tJ�B|p�sS�"/k�$�.2N^ӞQ��լ��i�B�vG�V�F|8wʯ/dVnl�"�GԢ��vS��8���ԉs���ٷ�{�V�ڷ��\A~v65Rm	�Om1�;����i�͑ԝ�T7ѿP�n�')�ܘv\x\F_���eV��Lsl���X ��6�:��u��:�Y�ƸK�y�r�W��^���v�o��d[S�뱹�m��ɖf�N�a��yf�����{:{g%�&8������3<q�w��kQ��a�e��u/��&�����y������zJ�l�1��]lun�^����	�=I$��_�Lư
	�Wƃ���LC����}�o���4�)�gK�j��3�#v�eY�i	�ږn�G^��F��s�y+�P�˸{�����L���#�t�Q�|�u���vVx��V��-�dB��-$+Y�J��\e�p����L�`��FW���W]'����q�2+0���.COQ�B��K�!���gҮ"GB�|n�BIݗ׉���]������C�[�Lkr���2���^g/��M�R��u���csia؁��ɽ*h�軐um	�zn5����&�x��(�&��|:��ЭG$����V,���8xz_K����sF��]ۄ��s�лY����nCҟGV��L�����fwL	y܊�}��!��`�d�XlÁ�f�p}�!8����n<���A�G��T�͌�y���Ct��f�,+s "Zg�c�t�;�_����{·3�J����\F׼
�<�<�sj������u�X��`f4����w���9Y��ݬJ5�L�볣}[I�_Ki��X�������������Jە�\�ޜ��# r�(`��>Sa���X��GE1¬�~�u51����G)?���0����O2W/��9:Xz�	��uLP�:s��<1f��ZWY�恘6;γ�`y�}��'��9��P����`S��R鉚����0���ߗ0��G��ܝ'G�����*���;��^�,�s��9|׾�h{�f2�����`�w�4;ٓ��F�toIq�uDu�>*���:�W<�,�qs^��|�!���	��r�C������v�Zt�qq Y�1ݗ��v!�Ӟ��q� �T��W�^\�K>��Ii�ћ�
YY������6�8 �$�]�g��]f�%ئ�l���%k�R;XҮW��'�>A.�ۀ��;�˥���{��Й���V�F�6���=�#k*|H�֗ �X�y�3�
�;�J���޻锭����|��&S�b}�s�K�zׁ��؉e�����l.�^}B���Sr��Ds*�Xq�U�[7ȁ}��X'�cM�w��c��MB�jWK�쪾���<�cܯ)����xy?a� nX��Y�{�5S"�G>�p�d��$�5��3���)�3�s=���������q_��9Ϋ�w��؎� ��Wo���՞�R��8 ڧ[�z�. �)��bV��m�GP��_��xc�卿���gJ$���]�h>�0���o�.��6�^��u�Nz�"Ǆ�`�&�@Tp�m�v����c0����W��,$]�̄lnz�1�^-��2�N�e�8�ez-�\���`^Ɲ�c�v���8������zzk�xֽ�T�l�.L�5�w,���R�<��X�c������v��K�л�FB��@3�e����x���Gy��ϸ��{�*�Eh�\f��N�[{d�/Y����K�}άR����kP;�fg��b�'���wk=�6UOL�m48�`�D�.���Z�S�s�)�B�\�֫7E?�j��_a�X�]EV�|�4/杞����7�p��s��@�R��ōЃ���ۥ�Yó����.P�z+�ؕݢk6DB���Ӷ�*]sqw�^o�������3�)�u�sS���8�~���6��97�%�����Ը�/� �W�6;Ԛ���s2uKz��LòX\�P�FoQrz����P�6/��,�RX������x ����We���5䖴�U�u���?����x�?����3҄�TU�Z�ŕ�e�ԫ��r켪�#c�P~[�-Q�=�yT���Qd)S�:��r���M4��9��8�&��N�6�qyt�2W[ۿg+-�y���v�=�>�=�������&�#��a�*�]g[#g6hR+(�e��$�#!A�����B�ʞ�.����}
�R��nù=��ve�<2��,�+u�f�v6�k~][�����'+�8�v���Χp늳PlEB�c�1u���[zĥgM��w�̤3�4�%.J�K�w����]Y�qgb�y0?�ƞ��p�8v������[V�X�>�9eL	��U�Dm���Rip�X��hac+3Y%��ݻΈ�:�P9<"n���dĔ��˱5��P�a?++���l�]��K>�.��-RuA��w��p���w�(J�{ٰ+��s�.^fbA[w#��/0�i�0�Ji�}��W�����W���T@�6���P���Ζ蓶���<�&�ƦA�=�/.�*�bx��(��&c7q9Q`��X��}�T���WW������jE����l�J��1�lHi�lt���^u�Ś뭥���r��F�K��Ź�,�M7�m>���	%kֲ�hꇊ���(����g��"m�>�}a�/�Ǘ�%!/�������sդ�{�M^%Pey�������}+�g	�A��U����[��K��ۣ�%{V`��R��T7�wϯդ0��5�S���B�`�����1�=:�;9��֝��鿆�WSW���u�X��"8�I�+i���m�N���=r�M�u�e�yC���z��jh�
�K�F��^z=Ai��{{�E:�U��ϐ�>�{8V ���'�9Ʀ�z/w+-r�{����U��aX\˕��ޥt,O�-%�0G�6ȑ���|&�l�k�uH�x��pg]�t�Η��yߙ�U�Aʗ�x���N�a�����qZ��/���pjf3v���y�^����w�4AӦ �au Ԯ���<��Nx�VZ���2��8-�i|��]n^n�V:�Gm����k��p0��Kv���g�F��й�ܦ�;Y���i=d�Аq��y���	v�"�{�����;�=�y����h2ߔ��1�ʿ-YȔ�}̮�,�N�ēwE��Nu�}ox�?o�� �p1�kdKGZ��M���A�\��T�k>����t�0�C5���� �/�\0�Zٻ��n,fU��i��1eO�@��H�V)�.��z��Pt�!,c�����_;���u�%������֠w�����z!)h<.T",Gt��rWN���w��z}�!{]�ۚ�O�L�Ώen�F?�a��M�z�|%v�K�!����]�χ�ߏZ�{*�l���i���������;����V>���+,xN�ʊǄW~�%	�&#趖�gs!~�=i����+������x�j�j�cR�pXW��ό�ίR���Hty���J{څ�{��˖�����[G�y`�L�ͻ�xo�q@[ZGpX�9ss9���W��W�Jo.K��{oc-b<>v��V=mpɉ����fst�ڧ�je
�_�m�����˲=�v�C�1����Xfui������R:)�<*�o�"���L�0y��s�ͳye�|�%�^�19vs~,=C&���1C����#�'�X)m��tt����Ʋ���[5V ����7g.�%�@c)8��z���4�[Gv�\ҡL죽0�$�cc�g3��m�U|w��8��w�|j�{"h��9o{��F�7s���7�N`ZLW"��wk�ks+��=�{��(��~�����K�|><]�褝�x5�B�n���kifX�s�>���3����]W�D�*�G��������g	�%���U���*���P���-l�T8��kӍq��3����,�̽g.g���0z���Σ�?���U\f]QuO����5NJ&�첅�]ӻ�®�ͣ���s�Ր��"��V:U.E�tp+����T^��ث>���vDB-���ސ���n9�l�|׭x�ce%˴M-�S-�єҊ���Ԝr��]Va���3�{�4K�6��ç��g��o}%���kR�K��z�_�%}�+r����΅Y�*%�K\�7,k���늖t1!�����`p��6����>���^^�I@ϑ�=�iǂ���u��n`F�u�����Y���`�#�⽽�7���H	�D!¶H�g����W2X��<_n�RJ�B�$�`����당�u=��5jĎ��fe�/�7����=��\v�۪>τ��$�y�+�^��w׹��tęd�˃N���V*(���OFI�\���)�;�.�M<*^p^b���yӌ��6�]����)�����M���M8�����}w��zz�1,��o�<��ۉ�ډ]��Ӎ�v 5���X�Ҏ�"|{狎w����2���O���C��N��ɞ!^�wi:}�=u�j�p_y�g���� ��J/���"|��/�	W�p�.L��F�T����Q���;�T�u9NK���0�|d�u�g�'x�S��d�?m�p �݄ym�G��o��Eh���o!���/���o�^/AN�+�E�S�r����ޖX���9ނ�ק��-�z�)Vs�T�Ծ�ǐ.ٮ���!~J���^K��Iꮠ���x�Ϲ��9}��/��ք>T�]gKĪ���w԰1'�۞�0��%e%��$�{.Y7�}�u�Xҋrr�Ç�*T���������z��k��%�<�Z�şWU����\�-(�,^s�Z���g��W`'7{ ��1�D�TsX��':��kyG��਎4�KA��t���mֹ2�kP�^C�c쒂ӂ(���]�)��"G�����c���u��_����"�dh!{*n���A[��6v��Z��C���֙�+�y5*6��,	9��nJ���s��� +��R��.�v�5C����t��p�G���N�P�q�A��x�S��RP�ŃI�XT��dʸ�<�{P�Nu�]pT����E��U�M+�E-�Z�eN\%+ x;�ѕkw^��h�Tg�q�c���}�о|���I�h�e�r�CTNR�Rꘑ*��!�C�zL���Y�[�����`�Kf.E���F�^v��d:8��{�0�<��Y��X�+i?�u��2d�c N�/:�N~�G���;���&so��+YY�ʳ�GvQ����sRJ�\ �sԵ��>�����iV�v*d��&^��	u�PT��qm�r��0�7c���D'å�\�.��� �
39���	�C��E��<���N��@�S\z����F>�7�>��Cc�pܾ�������ݛL���9���{�sQ��%ނ��v��Zg�-�%^U�.�Ṩ8V3��SVe�c]�1��]ۨ����P�5e�`R��.<;L��(�Y��ZD�1wf��4)��n����K�'�Պ�]4�]��];�S3���WsH��+�9h�X��f�ݸѾ�WS�����UO��@NgSU�G7��6��g��+\�G�n�ڵd#��c����
|���gwX����S-=)��=�O _&"fK۾�q,|4qeE�c�__�#)����ڕ�`��0^�_nY�)6�N]�s+��k���X��n���7_}�A�w'�Qr��2]�&�U,�h@85�i�;r�R�W�y�=�7%��9��<���]����,��.͜�媇�;�$�QܦN&{�y����x�#yZ�=�����nL�b��8gk���'��[�Z�T���K�aW���z��n+�a�3������~�o+Z�8��8+�:�'9˜x0N�ZLEgb(Ժ�ûyY< Z������m-�a��Յ�k5����%���f�j��ֶ�A�C�h�J�*{@Xl����L��3+�,Z�����?�O<$=��yI��<P�=^��n�؂~�{��V�bo)fR�um� ���i��&�녞�9'��v(����ˮ-�f�>�o���E)����~�:��;�J��*bb��,u�l����]�v�ij��5t�]��=\%J"�6��ś�IoѢ����uș ��x)���4�����c9������Ò�h����P����ee���e$!�h�U�z�f�ὴy�~�h
�×	�M�ȩ�n�B�EUԫX"w�5X�{L:��
�0y>��ن{�^�b��	ܾ���|f
��w-������d�����Oc��/�L M���/	�w�k�[ۭ�Qq�M� �Y�vpM^�mc��E��4�D':Eݿ���b���
枫;g��*R��9<\�e~rتޭ�g��=\BŠ�����r�B�N�^��ˮ\�b�6�!X�+QDJ�+"�)Z��YDQF5�[T�ZʢEZ°X��j�TE��Q�"V�U�b��T����)J��ʅ���R�ѥe��Ej"%����Z��µ����E%T-�"�,bE��Q��
�DDH�2*�(Tm�Q)m
�Q�k`�Um�e-��T��b�BZQTm����1b�(Ķ�@QTEQ����R�Z�����+�b��X��DAj�E�E,J��h*�EH�c����QD"T�1b��b�UR(�E�Q�QUPTQYQT��(�EPV�b1ֈ"�2*�PQQDD+aiTb��,b"�F���VUX�Q������*��EUQ�b-�R"[c"m�J���PDTX֢*V`�*(�*�Y�{�Ϛ�n4}�����&�
w^�����W���8iGuu��@H �V�ӽ�s�C��%�V�`��sU*����Q�7W����<O��D�"vV3�k9n���:���*�>r�.��!�W�)H��f�^��xO�u�R�!}�$�#�x���l;����şD����u�[���/��V���^�h|M�RPz�����2�Uґ�,+������;>k:�ӌ ���0����)C���`��R#A�)y\���։���<�_��g�}�M�z�o�3>姱gs�V�d���Kd	���yY*,(�oҭ���3�����}���ӂg�����O���_ڼ4+���ǈ��԰Gh�����G�\���]>έ9y��+�H���(5qͻ��V�c���ş5����8I�cko�;��%�N\�j>v�q#B�V<���O��	ʸ��JP�kuO�:�'��M�S�;r�c���`���zL�B�� ���3w�Wh=YN����"8���O��i�Z�����Z���7*u��eO&..�2V�ߺ\8e
�Jˤm�O�������c�2�ٷ�R�W���b�A�|֢����7+�c��g)���K�O"b�6��+ee��.Q�aYӆ��K!m�'�M�lZ<_a	r��eʗ�w\%P�".�9�l�fA��ʗ*��ݮ��}w\�Px�6���^xq��[���� s:�m�����V��	�������hzq��^���a�,]p�R�
oz��'qo9������TI�P�p�=CL-M�0	ƽ�z��v�<���{��6�X�,����h0%�"Wr�v
w�X�e���v#�s�9r��^�L�^��z�~	��Fw=9�V���DԔ�+�6�]���wR��:������q8���z�vKx�3��w3y�]N���n�H�f4���ƃ��:mbu�Y���ew*��}Q�GoU�c��Q�������>�����Z���|߆٠9��Gzl.���|3���m�z{�3\}|�-��j���-p9�ʄZ�,Lyi!Z�rWN��#d0nZ.z�Qt�%�}=%dZp5���n�FEf
�D�Wj-}*]�<&��#ug�l�j�oyןn�ԧԺ)x.�g׵�v�"���J����+,��ԺQ>���g;ZT}�����b���[膵�F�ׯ)��2^E��؆}�,jX5�aX��
x���N�n�^�C��g.�okZ�n;"8�a:��t�[݌UL�Hx�b��76�tq�ɚ]�9|+��G�V���Kc�vF���ݷW�}�<��q�98]��%$Γ���)5��{z)��sr�9\�u���Yw
➋���������ZXg��`~���T���xK92��۸g�׸�>��5�׶���bS�g�R��h�c$s"Y6�.K�i�����&Z�zQ�[G��eU���O������Ay��k%��>�/��r�f9vG�;���\��D�w!/��ؽJ��\E�dyv�W^7qt���[6����N�:j�,��N]�ߺXz�	�麲5�m����&,PZ����ji=���f�z�]Jn_�(��k+K2����u,x�޷�����ϴPyl'k>�20O��Pa8��"��C�1*�Zk>{��eΨp'�&u�ǕxٶE��o��Uܜ4�u#����-+I�~:�i0�7�=��ooμ�,y��]��׽8�dX�X��r��#��\\YA3/�i��+������=����[�z��&5}���aCð�H�%��4�����3�9龾�WX�����U�S�T#���ߗk��5����7�����,`"D#CZ�I{�Ȱ{���5j�B�.���˽����}av��tk�7�u�.�b[VɌ�L��ukͥyh�#�k=טļ�����6��<�W��g���k�)9����^�W�����P�CV�}��8���s�#�/�S��_]̳<|3��tĖmߞsm�wU����C1rL����偹c\W~=�5S�9r��.�g��}�_v��ȏ��x�#u.*R�N�]�����f�t����cW}���Y��[�UA6���w��^o���I ��3��[�xd��L��o���0$�IP��t�s���y�qz����ܡ+�:v�O��F�'�h���@���a���k4E��x|8���H��r��ŵ6x�$��g
�v6$�kR菔ܻ�ߩyND�:�,���GM��Zotee��Om�G�q��\�U��p�.L��{��`����Z�^Ջ�.y�]J���U�YM���1���;�}/�z�t�=�ŉ}�J�[�½��.�c�ng��,��C[�:٭Σ���X��v5eG���`��6(2�٘)�����z���#E����-�A`��3���V�����t&2RV���AB��Ԛ���N]ä����a^�t���=^�(e��	�nU��(�RXI-���x �;�?z�s����˼�=UG�N$مѬ�F��,�y�\17�Rwj�@��>��^����us�.F3��|~�'_.����5eZ*��ڡ� �4�Zt�w`�_r�>����3o���2j�����+���ҫ�7M�޵�|��X<��}׆>����߇zޭ�3�L�J*�j�KRؗ*/E*����t�����,�Y+�k7�d�W&@�����G{��^��o&&��ͳu:���%��%����ȚcWV3�*v��O��ӵ�+�y`u.�5��^����6Xw\�Yy���\١UԽ�mm0��e�Λ�Ƒ�ς\��B�v2��9]S�>u.qV��s���$�gދ���}�9%��$Y�����hGH�Dq}hPq_�ƃ���M֮�����P����28]�ǜ�����lǑ�c��O�W�D/���/�V��p�<vZӪi��<Kƴ>�/�̭V�+�������-�	܋9W'�i����-V�F�a�K).jϋ������%�����%��ȡx"�`䔈�nJ^W����$`��<ϔZVln�G��,�4�kn�σZ^.�H�\�U�cDؐ�$�J'�'��zאy29,�g۽�s�;D��o��i�T�g�q\>�^�����<G>�԰Gh� :�Q8�@@򱨍��v� \~�pa��ղ�{Lx�Փ��.qf�j�� &ɰ'������|ů��u,���4�b����r��a��4�_)I7��Ab���s�퐫�y�ڷgN�!��ze�角EI\V�s�W�6�W:�Gy�	r���b�d����M��Xͻ��V�c�������d�΍n�2�+��4�%��<�W�ܴ �[C�U��a/����/Pj֐���K�\�ޣ�8۲�[G�J�%by�=��֝�%i�z�]D�v�k�w�욾���%]�ͽ���l�g�Q`����:�=0���uQ�h��ե��W
�r�����F��A��S�zou�~6�$ri�ɷ����{�M�8���;�W�Z�A� ^Ί��8�=2^�="���u2�Ѓ+e�r1|�<#��Y�y������1�қ�Oo���t@��Q�({�p�I�]����e��b{�Y�����ʍd+��.�>M�{���=��"�},�5�+�6�]�ԃ���3R�=���e�OD�zx���c�u�+k��뱶��g��A�\��3�	�__��6��EZ�ȳ/5����^F*����^�3�g+�ZzeLY�O yh�H�WN�w�pn'^������{J��T�pc��yB���rg��1�w=�yǧ<wԥr�Y�2��N����������7l,tF�2YcU�R�%+��kZxr4o�LYR�P�,@�:xRѲ�b;�&��%�J�ej.�әZ��1~��j�*f�KNr�ܝ]3��q���-p9r��b;���υ�P'W��3��v��%�:hv{-��z���{+>�ј�0�U4N�iA�S��"����͙�]ִznɈ�
�W�.巀]��6���#0w<	X��h�vCORɜܢ�?d7��$��S��f�H؈��k\\I�<o��[M�:�epXU���=O�@ُ.q�g���}��fşwB0?m�b*u�Cl̯e3c6��^�Lo�T�D ��o��zV��G�Y6�.J��g�g����/*��j��;��Zn�lޖv���e�g�/�Dk����Χ�T���L��w��`�k�_��G��k�Wl��f�)�{Y������)��39�}����3��uh��{���'�U��f����N��݌[��օ���+�Vˀ��4�YZY�N�(Z�0���ua���>=����;Y���<gˍi�*���T8�����P�Zk�E�.uC�b��K�fX� r�9}(���M������{�>�ҪA�ʞo�]{5n��c��V�� U�{y�=� �^7�)���*����X��� �>H��kɦ�3�w/�&��W|6Y�z�<+`L�Ѻq�mf�Q��ҽOk}vޱ��s|������_Z�z%Â�B�N���!�����.�}T4t3����k��{~�[lҥJ�e�"��6�P�k���#�.-��f^;��d<��F���bvr����f�4'T��Z"d�<�˕������^�$K�_rih6��~�S���%�����y�I̦G���o˝V����O�7����;x�E��r�w-�5�!�/}b�ӯۍ�n҂���P���,?;\���~Vf��U1q*�x\�v<T�p�3�}V��Zݐ��pρ�H�-+>�"����4��K�^�n`F�u�S�{-���jt��Z�G�؟.0g����
�
�$p���w��xwY�;����T�Eg�l�Yk�Ni
���I�����̺��+>�j����\7n����]=�B�$�����SZc��[ ���������_OXg>�[�;I��@�a�R�5x|���X����ݚ{�E�u�$���=z@��ڬ�`� +$�v�r�;^��Y�5��x���F����{L�q[��Eݺl�۔-�0�[]��[t�������c�fA�v���q=����٦�h|�!�z�����T�S"����i%����w�i�����cs������Xi�}�[�d�����ٷWV��P���O�WA:]@�y�돺eMFz�T./ G�8�g��]X_|�V|pyǈ�Ք��͓��H�6oz=ur�_�	�\=����I_*��a��U����9�
�fp�s��q=QΡ�y1A��(d�9�af
^���ew�A�T��2}JmT:�@�r�ME���+��P{��/�2���d����Ǘ3!�k�<+%&�qx��$�z?0� ,�w�O�`ŉ�ĝ-��e���Ģ�r�rޯlδ&J��:�ª���n�{��Ӟ:��}ՊO4�M��"ߧ`��ެ/J��بh"���N�1�o�[ny�����=PDy2�\�򞂛��$y����1W�u0��C�馽˽�=1ny�� 5�SS�:X�/�3��<�:��:����në�џ2#�`�*���խ��n���	���t�4Gօ��A�Y�ugS�u�ү܃�,1u���y�����Ws������v����SC�	���җ%b��Ԭ{�uɬ�Z�7�}�Z��á��������ޮ7���ѳ7"�)��l.<�:�మ�ȫ��v�ϲ$N���T�� ���y}�JW��O�bo9D�w�GXX���հr{��}n�j��6uO'�R�*3wsz+/�kU�'óke�.��}�vk���Ɯ�JV�`���T�p��I*�H��T�"��yp������Z�>�kma��]�Xwz�\dP���"Dx����=�'����`�S�TX����Sޝ�65�� ��-��'���\�U�cD�S$��(�X�ׂ�n�we0�wzZ�hdT�Ϸ�]�B�mk=��S�:Wk�
7��x�E��^�
�cڼ)t��X��M��$W��[X%WX�[>�/�x_�U��S�WC�t��xϸ���^���u3�A|�1\�N��O�A#�A��,eRՖ=����J�J��ͻ�ז���YN;tz��s�W� ���=����]c'����\8��A�}ذgTX0{�8|���Y��J���9�:R���ħ�}��cq��hχKe�pV�3>�/�R���޷g��I�1g�9u<.;�s/��{V�)����J���g���uqRb�4)����~:k�Yy<H:|��y3w��\ ��E���4���N�e��a���τ�^�_���}���j+p/-�I��nT;���鷮�,M��������o@}.=�X��
�E�K�r������H�}L�O�s��{����Vs|����
��;Mg����A�ua�) �>�F
z��v��
��J�p2{�LB�Pt5w;��}�(b�c'q�m]1�%f����-�3�H�}��\\����i��˳P�e����B��`�6s��4��ܧo(�#�ɣ�L� )��/�/�2B7��'��>D���"W詖�:Q�H��^�tޯ���E�c�)�c��Ū���ʭ���5��CNr{"�\^-��z-,v�n�/�:��S}�P�H.o�ʖx�۷�.G@z��E�ɳp�h�.�e�|1�c��ʗ���W�V�>c�Իh�gm�U��fkY
K���������P�w�R�,�C`�u}�Ĭ���O@g�WwW[f�[ջ��t=}���[ٖ�Z9��R=�_�y�{,{׾�]3���i;�I�c�yL�9�ò�u��i��.aR�f��W|F`�.J�?*z�K�@���)�.�x)Y2�X����1��f��x��w<������S�M�3�4 �wդФ7�҅�a	+ln��O6k�n��pLwC{ʈ�*�5GO�]���1KK�/�Y�د��FA���G�v�Z˹�g�^�3Ku�-W	$�R��K͕��_�����k������ĵD��� c��E8���`����;6Y�`3�!�z��H&���s�s{�w�yE���잉���L�z (7,R�����_K�\�[��`��|�.�r���;(
�w���5S�}�<ϓ+зR]����5]�@n�y�s����J3.]��X�v�����!��r�bo$d,<���{��f�gn��a��^;�O�߮�@ƞ���aA��Y���XT���-�/�,�p�!���.��+�hG:��c���^��+S���b��a@��W
G9�r9������N�����3/�vD�����]�� �&���|�9'�W �ڋF�x`��֤f�U�b���^�7 J�o�{𢣏4 ���f�F�&���c,*wa�6X}�y�]N��]��H�<���l�[i�<�p��@5���jto.�8-��(�Ӆ��|$�iͣ_G7n��,]����V��pn��e�b�X���nh��ss�b�6=��>)�@�
����/[�Ɖ�)tC9�n��:�]|�]�Z|����g�}-��.㳞�}�`�����h5��vM��F�52��Goa]�(�S���e��Ci����L����8n��n��r��DҴ��cQ�|'Y��n��e~��zmK�����Qk'3s�B�QJ��;p��c�����0�����G;{V���t���Q�v�-��Lr�r�]���
д,K��l�o[�Q8�o���&��DJʪ�*��DE�AmhUX�D`���TX�Q�V,b�AR(��

,��b(���1X+�"�J���UQ��AJ�D�H��*�eE��1U��ETAEUJ�*Eb֡YX�[k��UD"1b(�Kb��������*�+EV,U��1b�F,�TQ-�QP�d�X�Q���BڃQF����1����m%cTEEEm(��ʊ((խ�DTb��Ȃ*�"���+X� �UT��A��(�PA[h�+R�V"�"!R�QF[ee��V*b��*6�T**��E�*6�T
�(,Q,`��E�!Z��yqlػ����;«7�j��_���WYC�B�e<���YI!���7�;��%R[�Ga�>�v�=��"-��}�wy�Ɉ_���ж��'�v��J�����V<�fl�F��d˾���[.��:�rp~�jl��lv�2�'��\����h!ŞH?T���{�Y�ف)�!J�����^A�=}�3��#*]���M7	t�����$�k~���%z���Rjv�����P�� �q핢_�N|�Y��%LB��-o�<,<-\�J��.�M_Ig���ƣ�[���	�)��G&}���j��҄���P�Rŉ�夾�{ض�i.�3��[s.w�n��ǲ]��=Y��z��v���/��h����rP�^[ƶ����r�+��R�,��&���9g�yw���׋�B�c}�O.�Y`����Vfm�^\�;vO�����c������lDp�k\\�y���l57|�	��^VgW��b�М����X#�t�λ;����Z�6���=S���=wU������8�k9�����q ������;~0�U��_z)�7���?Ki��X�^�k�;�(�Η7|��{�1R^Yƛ�s����7q��IS.�a}�R�N-h�Wu��;���[��t��jb���`��愫�$�z.��q�q@���I	5Qޞ���y��S��swH�����C��1\lc��5�ќ}}1�yͧ~3�*��i���'�]����:{p�ktؗ��5��'�Ͷ7Ek�z�f��dr���c:��G�8��ى˳����&���13��x;���	����T�0>5z�R�Bӡ��0B�\i�ZϫK2����K%(��Ǧ�����/�W�<�����ȣ#�8Ȗ3��Uh�K�V����#���G��:�n��T��X��J3�8��S۩����L.��:G���!�Ih��Z�K�ZpM�m��*>���9���j�l����5�ƃ!��c�]�V�xY\\X(&e�n�ri�x�O�\��T7�N����.{���_5�BK�Q"\�@Aĺ<^$���oz�O|פB�
�,erR���<lu;~]���gyY�����o6�RU��6��}od�"�M+�5L�P�z�P�~v�`nX��Y�{��b�$U���wX���ܯf�r�:q*O�g�n��0�KJ�I�ׂ�>W�4�t�����"�	�nÝLu�m��X���W��[�2�e��2/u.�PL�w-�Y��ٗ��sB
lK��
���-ML��{8<��Z��l<���Y�Yf�;Ҩ7����v`��BRR����Rђa �j��B~�y�|��ym/�3�����/k���䙽i������ڔxxa�lx_XD/�
�H�k)��d�׺ǌ��u]1٢leM��W�JzW��`蒓\1�'M�2������H��Y�^�t�l�ߕ9=�'��ô�|���Eڇ��K��aIA��JƵ/�u_�-���>�f���٧~�.����{�1j�ׂE���i���F=�����p�,I���}w,��[f�>��h�ۛ�V���̩c�k��R��GRɈv�����v�沛2�r�$v���/�gB{��T���?����5z*X�ya�B���lPW�����^7*�u���uw��;4�V��!�O1�vb���xa-�RPa>����k�(������F*�k��ރ-?qs=��*nf��oW���w���B7 �7�p�x�Ih� "�M~�<a�x���9^���L�;
�6�P�Bp.[��R�X�*��T8���-j���lߑ��ۇ=ݜ���=ll��ć�u�{H���w���':��kyG��਎���}
�3{.��ʰ�Vj�oP�H[���/ru#Y!�&�V�C眶�5=Ϭ�E��wp�h��Y�G��dg3R�o�ݡ �������ls���Q�0�E��O��\ޜ����	ym;���(��b�e�9��d�n�4�9Cmi�.��C�D�.�)S/Ӵ�
���:����h˞ɡ�O�e�uʵ�{W���z�g�]�S�7�������
t'��2�*޵���Z�<b��E��y���4om�~+n_'�5�Iᓞ���A�G�@񹆉���$����W�q��,庰u;�]�Խ���ʧ{��Qڴ:r�z�R��|'�9�O�>�i�.J���\1T�uڛG�r�����d�-cE�4�'],�Y�����rJV�`��4ڗ^��J���f�Z)89��r8yy[�;��w���3�[�k����탒R#A����`I��<�i(s o�ݿ,w;|*��^ٺ�,�m3�T��j���k�����s	V1�=�p�l@>� ?OB���֗o)e��o�y�A[�b�C���y���e{���k�
7�#�g.X}��C�w`�r��+��O�&���"��B�H����Y��넫�!�x�ĺ�ؼj�3����r��fsv���p��W���ͻ�-3��d���y�p���+7(�/<7�Bwa�̂��Y*6'�*����7� ϽG�X�4�g_==J3[��\/���a,�P�@��6��o!5L��3Rp��4o��^9�p+�c�[9���S��$Z����h�1oN����|��wذ]�D�3�Bҹ�p�+{Zw�Ҵ�Z��
�Ŕ�J��+�A]�L�����jTkp��D r��Z��|g�B���Av�,�¸U�[-�\�l|�\}���g�U�����"����
�=6�:��NhS5:��3�5�t�f��y��Ԣ�7���4<l6�X�Cf]�x�:iXzj��2��0|�v3.c̝�aOPgk�	ٻW%�޵�ʣΩ0.5��	q�DsV.]�z�/�xp�_zi*�|����E�r�9��٦��s+���G��Y�i�\����a8��T�����\�f��bwZޔj��P�{�n+�u�fŒi�s�t�q.K�LƲ�dc�b�_U�=ժ�:|�J�sjQ��[/פ>�z�d��Q�2�%0Pn�Е:Ȅ�x�(m���I�l�'>%qw>�fy^�r^=�r�yl��]���x��g��/1��"�������ߜ'���I5���e�=`z�S9�G��u�3 ���*���>F��7��au>��-���n�$��4ojt�Yy�v�[2:U��m{YQ��_Uڵᢺcō��.M'��76��&������v�r�������`����Bٵj��G9ojV�����."}����i^�D�C;} �ȯv������ޣP"�����\G,�/73���{��+vN�%w�(k�c<�U��{q]���Bl0�������k�P�O�xm�L�ʻ��_j�?z�5z����7YE���zV�J8Ņc�d 3:�<GL���1Lv֡���,�E���[|�μ�X��ʬgW�0cu�X��g�s8�3�,���U��֭�����]�q�W�W�g��oo�cbkV��A~�.#���$�#���P������:<������4�Nċ�=[5��,�PR�.��u"�Ϋ,ڜJ���˳�t��]�����{��o'���ᯤ��.��ze��{Bxb8�:>U���B��9�i�Z��if'S�7bq��᫊��؊��7�k*ws�;�O?��E��i�U��(q�(u���P΢�G�~R�B�xn]���;c�M0��E���3A�ͩ������t��Ih�i
���wi7I\
_{�r��5M^�Esϲ�5�}8�d_ӱX��r���\\W����Է"��r���#4`�Aj�̴�N7���3r�C�ǖ�OJ���+�����O4u�3�yb)�sv{0�M�n"�{�]Ѥ�3����'��D��wDⳲ�B��$�B>]���[����t�����c��e��4eM���h��vwPx��;skbe����r���x�-lD����c.�����]3���Xz��>N��(T.�.'��.���r���i��;���ogi��e_QZ�)���ů�0Ь�P �
԰R�(S=yQ(_�.\ܱ��+�늖t[o�p]m��^�h��>��a0�$��KJ�I�ן]���<3��奺��tEd
����қ��'�P��W}�B��ࡇl}S3>��"+�k1�<5��^�o��ZJ�.I��[�W�V����\�|t�P�K��H��^��ۺ#sQ���ؼ#������w]��k+��p-���4|�=��c������q����C��RD�Ȇ����g��i�t`��@�p^����n�ǻ��ԣ�鷻��^��d'8T~��ڳ*X�c�b�x�x�꺧��C�,X���Ft4�ʲ{/~E��/y�b���AҸ���h��pz���>^u��u�[��4�}[�8x�l�T,����1֩$ё�n�
����׻<���n-�����fm�p�J���ˉ�Y	A��<%ojg�g�T�{޿M�ֲ�6gl��s�YY�׸oy�7��Qm<lZ'��r�Xְ��!�����wU��#]	���%rW�2`����wG�ݞ�g�ʩ�l���U�ST:����_P`��d�b����ӏ�Y�֩��b��2}�-��Lxf߮xVJL8ۈ��,��%��l�}n����J!��i�ٺ��&?T$�D�W=��9���`�u�|g�	�t8�Ĳ_��˂[��XR�5~Ns���s�U�2�ىF����~X��v�;���(Nu��Ʒ���7u9�R4��M[-)�4��0`Ku<�\]'I��OɩP��H�'�8��o{<l'ON��C���n��Jgz�x%��F��sS>(s����]S�K�^�*��������W7�O��w�nfؕr{�����<���&�:D�q}hPqg���P�ի�7}Q<��p���i���WE,���.�u�.XD-�rV*�K�w�}Z�+r�����;�Y����׼v,�����i�%+Z0Ibr�S�-$�:R=����a��}��5Ǽ��)JKD�'��;�I �g���d���nJ^W������)z��9��ebN��U�����V[Vo����~��N!�Ķed���Y y�<�!��ޣ޾�.�Fڦ��Y���~�]2��*M���fn����o���q�/��d��Q�H�͇�o�v9�t�a4b���Z��h�OA� /�^��r�Ǖ���N�:	��}p&�������t�Y�-k�J��h�
d����K���Y��<:�q���Y��
5����Z���:���c>�^�~�E�^e����<�Aj��-�^�c5��0f܈��L����j�O��~�nxө��g���_������$�{�Kk��� �v��7��v�<xƸ!�r���'����"�ϞZ������U0e�� [C�N]���-+�.�	ޙ^��e�������������l�/��w�^հ����Iϫi�����K��.-�s�����ie�yXZo�/a^���;+E.>�̵�]|U���q"�T�A6�����&*sB���z���av�Okang��������Ї�I��λ��tҰ��3gZ1��ax�r�_���˿{�>�3��{"C=͑��ж����$G5R�w��%~L�5�w<��ݵ{���Q�hσm��{��3�:{g%�%Ĺx�� �k����aU�^�j]���M��8�Ci�ˉM�k< ��'�kټܷ��$] �Vke'[�ѝ���fۖ�8X��˕`�9K�5���hˇv���p�[O\�sk�Z9�JP�܁�cu��|�lkUm���:7�y�w�mq��ˮ�宫v���j�S�է�A�z�˸��W.�l�~�F�Bt�T�j����Y���uF�%�?�	n��X�C5�����_J�^�S��eLJ`���n�2��G���N_o��r0�J
�e�T=��	u�|����,��[=g�(K\��9W����Z�S�-n�R2�I
��%E�y(6ϙᵸ����D�A��B��	Or�GX�6>vv�o2��сЇlT��: �ζ��h��r�����;�բ�d�Lz��{P���f*o���3U���i�Y��+�p4q	c���V����j����tP��.'u�,��rXԳ�XW�2�bgVG���{�B
�����xK+:��3�i�gz;Rj�ݥ��<��W����L7\E�pX�}�1��k�r^i�H���jݞ�Kfd�/A��v��t�����F����'�Jv�{�[�c��Df��e	�_jd���b��3�C���=w�-p�F��F�X`�U{�}z��s��N%[L����>��a� �H��G��O[�4�jQ/�cr<Vj�L�r�d�x��8�wi��%+@��������`�$/9��D��Ǯ&l�VΪ�ZP�m�Y�0=���@��]!݁�?>V��ۈk��iQ�<���>6��&5���s�ܢ6��;����>�vۗ�{�Ҷ�~*��@�7h��U�y�W�L3&<TT��x�Cs�:����s�VهJ���[�����n����2���x`�и1�|Y��)��Bz�\a�ފ����dAF�g ��j�5�9|��n��Y�!�� ŽQ��]�+�;h��Fՠx�'�9;8T}p��;0�����9�v{�s�)���n����hr���m�k�7�Ok�.JwKj�1S<}�Z=ӷ���U�{V3�q�<���	�p\�7���q�lz2v�8:�n�ڴ���FP��+��9���z��%qU��YE+�x�Xo3s)�:��+jf�F�˒��O�-�sͮ�ԅ�X�RMP���2�]���ϸo�u5WK2:�K�|7���y:}e�z��ʶ
�Q�ϥ�ׁ�	�s�݆��|'}���nGp� ��G�X��*�<��1�0qOx�w'и��^�b�T��c	o5�o����>P�p�A���[
Ǽ����1��}��@i.u�d`:���ϕ(���*T�Y��VQ��bR�i�������uJZ���b�ډ���>��(r���7��WC,���o�w]G�T3i3��!=/*q׳{Lif�޸8�d+�˾Xӫ	�']�SmG�gI��5[->�J}���i�u��䣻#�ys�mgx_&���J���{<&m�uo(����aI�0^��+	��7�"�2�E@tA��ƞ�އ���]���@Pa�ko�tM��7q'�q�6�ɻ����4�Jà�oq�,��jP۬�m}֬��V��)8������5s&u�D�^��v�T*����a�z��\��j�م��Ƽ����;�iex�R���q�I�=mA��̧��t�/zY�[�~���dq'<�)'(`gF�v���Tlo���O�|�I���������ܜn�j�"8v�Q	�Z��]ԛ�s�1�t/C扺ѽ��j�:r�C���7�nc��t�r,]F�QVL�'�j��ʠY�g2(�^]uSo�ZR�5V���z����Z&"i��,��Sn&ioh�6n�W3�8�Pm�Db�s����c�������)�;1����i��|�1XI/�j�.�ǉ�͌��{nA�s�'syh���]-��Sܮ��D�g�=*2���,���`(�43��Z�V��k����EE��F�w]@��B5��,+v	���V���m�l�����Ǝ��`YN��I=����Pf��N�Z��$�Vǳ�:�+�n�f`��\�1ӱ��N�X�R�Ⱥ��mh��6N"��>�:�����Jű�T�-,DQR҂Ƞ���UX��T��"*�[k���QEe���U��*���Vڌ����imDm��1U
�j�ڨ�VV�Tb��"��j�E��V�TTb�F(�E,b�*QڱZ��U4�PD!f*&-UQUU���ūij���""#\Z�+m0�LFca�Aepʘb�"�b�P�e\R�.-���jQZ�m��b�`�*�����EQ��S����������Ub ��Q+b�2(bʈ�T�Q�DUUQA�QQDY�
��,U�(*�Qb�0Za�����1�����[A�*U1\$��cF,���J�Qf-�qp��E�X�QqK0�E[(�EjTB�U�)E�qe�\R�*��(��iQ�����'�����l����;��jer�R�G���2�GTd>Y�:5p��	4���zG��9��NZ��s�M���Ϋ[���l�	����!R�t9X��
�pҙi֖a�V�=7�y��\�Rt�YkK]C�ϭ��.WH�妴̪�M8���3�ɘ��
o<0:�6M��LrȂ�����/�S۩��������x2,��3�J��f^c�cd��h������P\SW��Q\�쳅��{Ӎ�E�;����\�H���r��ݴ����^�m�,�R��_�:��C��v���8�{���K�k���_�(�9缓�Ö��og�2�w0�	��(x���P�e��җ�W������l:U�۰f2���Ȭ�Ȼ� ���U֧ڰ���A��Ik�P�{J�����+3O7y����������f��������) *��Z=�|�v���\�|֛!��Rt��@j��^�xb�&�zk_{��Y�a��S3/
GK#�]&v]`���gn���������NY�e�,���0$�	*�I���)5��t��/���2�Vp�=F������ؗ��°^K5�k��/1+3�W�\�j��ՔMdO	�z��X7���p,����-S~J��]Ms���V�~ma���r��A�U��{�v�\[&� ����t;S_�4�-�^����Ӂ���vY_l�� �o��Mۃ�G�w|�/;�±%��%cZ���GU��e��F����纷A{�天\�>��/ʌ5�Ze���4|������w	"��_���a����u��g@s|gu�+-�<'Q�2R�.7�G�3��,x__���V|X�~F��9о��[�I��G�SeN�&׹��Exg��^k��r�"���`��UX�;��t]٪�s���lWq�3ڸS\�6el�h���-'�-(0�U�B��^^�����y����8�P`�t�E��qX�d<�?(x����f��ݴ�<Zm��Ǳ�O���n�ž~M�r~e˖M}n��y�Leg�iEb)�L�z�Ϲ	�����T-���{r�w77x�%�<P�\��J�H��A�c�E�N�|%	μ|'�M����^�!LV��Z�v�e�v��D�v(���Ӵʉ���\#ޓ�W��0k{�ƣ��l$��ἻE��u�=h�v�#A���
9���L�S�R��p�C�*ы۷�᭎S|vu2�e��o0Qʝ�������fr:�\��%F#���ݞک���y�Y7�&�}�cn9%�P�U"U����f0e��\Ya��r�v�f��3����k/XCU��L��Y�z�Ay��R��>]��[���zj'��W�=�{Q�ݻ���$�r��z��
y���'H���W�F�|�7)��u�����mH��2d^zk�*���襝��e҃*XD*؎��V�zּ^��irⓝ=��_���W��\YذKɁ�+��>���%��*`�e����ٖL:�9e��B��+i�W�T=jό���Xwz�\�SD���dKk�ѱ�9��8��	�Z��0u	��+������)�>2�}�-�Y+Bf4I8�U�d/k;7��P��a�EQd@?}#�ׯ_�5/ic>�r�����iq�j�����r͆��r��z7Z����`(���E�/�lv��{bϾ�봉���p�J�sƝT�녍z3A��;n���g�s�x։r�Ł�����Y7m��7q�~�]�5ZL�,�D�=N}1���;={ѧ�y�z��X+h⭇~].�Pq1�0���D^�ʦY��y%4{���9���oۭ�_j��2��>��8���NV�2�t��p�3��pˋN���7A��х��ڱZ�#�ŕѳ�+�I�D[�Wi���4_�1��$�f��NX���=㳶�^���o}�p��\(㻾�p����}^Eԡ���g�j�:-�K�ܮ�=JN��8���"�4�ce��ɬ&x��<�e-MB!�b��j��Z`�9��R%�M�As�FT~���C�67��߉�va� #�z����:i�4!��~�Cf��=5�֌�������u'��퓘u�E��9�<3��hl��#�:���[�ߛ�<��f-Ew��麸��3��Gɒȃ���_��i����dp���_tK��>A.��4tY���K��v��D+���,ꮉ��ܡ��y��2T#*]���I���t�q.K��ç�I=��=�c}���Q�>"|/M}C��j梴��^���,���,�(��ɒjE���Y~|��v����f��QK���7ᮭP�#�pO��<����m�W���{#�?j~Cs0�9���R�"�C��H{a�J��y��=Vjg�����V^/R�1����U���̑���N��Q�Їn���� U��=����O�բ���6�\D躼�_���3yQϚ���!��dv�ؕ��8��%��]&{ړ<=k����ۊb���t��O�w�e.w�*�Qn��uw\M󻢲���Z�^�	z�tw��~�u�ֻ��1]7�N�s"��g��Xp��/uX�%fR�������3�IJĺ�o�reo�i�+롚i�P�� �@B���ʔ]ʙ�h�nt���Ι�W�o�^�^km	��jY��,+���xa��`~���T�lA����r�X�]l�L��4���c5�Aɫ�P֑�k�ǳ�cK&ע�Ztɳ0)!�O�w�NN�ҝv�ޱ��z��.�^/~ˆ�j�8��ȏ����IvG�y�e\�˦��Q�KM^��!9�5���G�H�J���>��VX9���ϯm���9״j����R���K�����]��qJ��ݞvC��W��<�H0FVˀ�i�ZcK�)S̳�6�����9�x
)�C��ub_��ʞ~)FGp,�c=*�U���U�:W��baݩ;�1�w�"ґ��>{��ꄹ[��C6N��eaL�]K���A�a~�@����k��\��6���U��E5x	Ԣ�}vx�����"u���r��*/-���A����y��e��ݖ��C�u;sj�L���%�^���yN���1<�ź1��l�^��
��r������K���q>E��=\���s�3��C����l�^]c%���3 ����Ս�w!��>��EФ��w4v�5�3O�F���8����� �
��AųM5:����wQq�w�y+[�d��9��=���wr:f��}כ��fL޺xp\���e��}{=�={Y���O��^�����E.l_{���m�l��!t5�].k�<7*��>���;���ֵ���#�Z2��KY櫜�v�Y���x����Gˇp}S0�EF|5�ҬRqu��G��2�ܙ��¸9�T��Q�6����dA�Ev�zCVxb����a��Ƒ���Rge��0!�|wh�}\��S��G�Ǟ;��Y��JĕW&c>��\1�'H�U��$}����W����y�@Q��i�j�׆y3���pXV�2+f��e#s�IcOϟ]�����ɳ� Q��wT�8/5,�x���0��咷��${d�7s^J/N^n�b�ׅAw(�ؾ�^P�a{Vg�,q�M}�H�=�����~��K��S�l�ͺ���ܣi�1�1}cuxG\{��4�=ԕ���X\u�[�q^\̢�S�SX���ݨ��u��Ҕ��á���;�V(�6r�o�_ۡYܪ���:�@�]>�ٕ=�2��^��e:�j�Hч�/�].�j��/�xxf߮x}���Q�D�\c��&�q[�@:�ڝ�.� :=R��'��4�u�	+�v�|��_scsq�F9�N���x�]���a��nӨ��P�8�{N�]������;ߦ�]�Wh��g�Z�}{�v�=����5��:mș	[֧AΝ��«ھ�2�m������Z=>���p��2�=�3����(6
gZ%	g�gv)ix:hg�7�����n�b��W�.�ʨ�/J��]�N���^4��%��df3v��E����*#�$��Iآ+�wN�8*S�jT#8N�a7�+��x�}�-�yQ���rvx߃�ֵ�#���"�#A#x��[ޫ���Z�-Krz97t{p`p>�ڑ���Z~��~���̦o��&�h�s�I�8�����Wuyw�eaѾ��_Ef�@���:�î*�A���z�9S_���p��p���d]OY��}��e�����jy��6�t���6ﯗW�}�v9���$�kFIbrR�Cڷ����:��6�t�}����_.Z)4�k,X�Ƭ9�֒(_��2$G�>����|SéΣ�}ݨ���O�uG*��^]7.��zpz��Ayހ,ka���t�߻��� ����r���f�t�Ye�^�_7<i��>2���ƪ���� ~X��w�@�r�W� Vh�]ֻ4s�Zܼ�2Med�f`�0�I=�ti+���yvL�{+�y#��N�H�C����a���\G�y]��J�i��&��ٹ=��`Gv�˵�$D֠�p�_9��n�sX��]�yD�0T�@�z7��e�(���ೃ�}a�Q��$��~�i�۝+���OM	�l�]GzkeS`�[���|����idݾ���ѡ����-����>�S4TQy���Z]'A�0����b�+յoռmt���L|��;W���, q��3��u�l�8�)&%�Z�,�Mr��I�[ĻV;��0��V��һ��o�Z=������l���g��I�<�Oh6z��Бzg&�"ӝ�jEpl�^݌V^w�A����=��^0�
�\����6GRwJ�̻�񱎚W��P��U������g��=NA�Z�jGb9��τ�^Ձ���`wh�k�p6����\���pj�[���z�3���i5˧W�I�����A��,�4
���;������Y}�],��"�O��R�{n:=��.�(*����>�MÒ��[>�����o8�����<�%*���,��A��6���YS��,v�z]�,�-K!��Cu��~>��+���В]F)Z6k%�\�r��q�gGm�n�+�9�.�l�J.�Q4�ܸU�s�>�}�v'�w历�f�]�){x@9k6n\J'Q�/���>�z6�^����oN+xo\�I�)"�U��%z��8�@�ᷭu
꼛2d!,��3�������M��xs��k�@r�#�X���>�����u��'>y�;�t��g�'�A^��U�&�pZO�:�/ ����S;�@�Vn�Fj{�C�u��nA� C�W��u[�v�qT;b���xM	|+��|���oٷ��/�E�r4U�[�K�7����"��=J:G�+�q��K����Ӳ���|�_"����ܵQ�g^r���C�P�\5�a_�s "ZbϹ�c�1��A�N�O���Xe�.}=��vM���8ӵ��T�{��P눽pX�����mz.K�-:tM��o6"}}Cc�J/<�}�>���UoɮV=>��?�'�+X=�(=ܐ�5v�ZX@+;�d�0l�Ȥ��V��}qn��G��X����^�ϔ��P��g�N���VA`%((/9���U��<-����0��Squ�뗌��н���kK�]B���Aw{7[�hA~�	L�T<eԹ�Rǎ}����T��ȣ#���`�K�H��@�9.�u��ӡ<m�𩽌R]�i���!I��Z+,ksx�����^� "��J��ّQ8��u����Ur!�Z�U��e]�{�s����?`{�.=L�HxM��l�9�.�<�Z^��Nz$�݇i�� P����n�uk��ט��l`�����x�e���C��/���sB�����pi{o���[-���Isb��{o��U���wT����<�u(�	��g�����a�:��X�epS;=w���iM�(���3�Ǣ�	�c�-!և�����&og�L��z�=��"���i�W9�gBF�l�Y�4�BQ�e����Q�q7�S������-���z|����/�W���8�s��y۷�X�(BjWK��=�eD����r��;hy�soC�~�|�y%fi���.> ȯ��r�ܩ�K8l�5��e'^]��K����.܌����YZwΫVw;�dA�T�HUࡃ/I���Ep�g����kʮA��.t|��x��$�T�-��|a���It�W&c���Ih�2���&S+_[�ލ��j7W��z,� U��ؽ�Pл����C�)$��aX��ĕ�jS/��=��{�ٛg�Xy�	�����/�,����C��������}��h�\t��0� ��g���$���M�4e�CpA�^���%]֝�ʵ_}rb��6A��ʴ�t@���"�wsh�k��X.�-Vf��«W�����f]��t�j�K�h��8w�Σ$8��$�rewW[���mX�l�>�7Ԭ�w�0핂��Y���s(��:_0ik�������:�Ô܆Z&�K�y"�L���0�91y�/*��}94ֵ�̡�������3.�R=*�;��휚�m�W��J-USXz�'=˵2c��L�t��V������1P��:��#�S�lf���z��R;NOg�0�<Ӊ}N���<��{:�!u�U�=[���u��4ی��9�+� ϻ/&���{-h�!���2&n�R�.l����z���-k&�Y���D0 w}��)��^4���Ԟ�[�xA�F~_;ַ��L�P�y�e�;�X��+�յ����č�W�3swT9�!�{G�D����d	�UUT�Vxa����+��c��rf�M�}������Ȧ�c9��l�`Gh�M�$&NQ�7"���-�t]1��4�kjʱk��8��[��w�%V���r-��3��*>;Q�F�����{S��n����u��[ռ쮙f.n�r��tܹO��D��7���E��5�b��8f9������E�	�U�n�]��Y�v����������(��� 6&q�W��6aK˝M�߶7��r��ĊO,��A��Ҳě��.D9�u'Ѫ�,V������sJ�Ǯ�չ����c�o���<t�V9|B��h՛����X9���M,s�F��=�����X"�w�B�yN�TI<n�Aj��I���]ζ��R��I���~�씭����&[��㣢��{�'PF�	WB����?!��4}�[��nҶ��8�p�em�,�M�<#����˛�n�w���d���ρ��=��L�{� w�;�����/x��ģ�f�qfIve&ϳ����Q������4!��R��{y5r�Ogu;r�B =+1��W�s[Bu�2Q�%�;T�>�,�ݛ�P�� ���mݔ��ˡ�Yxwh�-�m[�Km�q�d-Z~y��������y{;�?+�ffo$z��h��8�%l�U����������:SN%�ٷ��6]m��3��{O[��I�����|rt' �}��ۅ�,��Z6������v<m�����^���Md��נ�Q��ws��:�qT�ɫ
���$r�8E�WL���;�uN�)���wI�z�`��<�𥧼��^B�h0dR�Ρ@Z�:Lë3^[r��@�J��p��v�bE+M朧�Q}r�{���ȯ��R�ȋ��3���w�̆�R�;�����*5ΰQ�p;n�g9���'��p!����{�t'�i`Aov�s�
Z���}�S�Fc`%n՗�ݏ�c��x�{�*ZQ��"�K���(�m�(�F#m�"�"5
��b��b�-�6�*1��ᩆ�,X�*[(
�(�Fb�X��,QQ�ȘiT�)R��-�
�"��Ų*��EE"
�V0Q��b�1%�"�AdQE�(�((�
%j�������`�-KZ(��"��mDEEUf��J�ڪ��(1*�����
	����ZD%�LZV�0�X�1U"����EDb�YiE��L0��"���Tcl���hUQ"�TU�(�b+UPQEQ��C�C�U��,p�E�* ��(#���X����Ab*+EUDb�QX�E�T��(�*�J��EV0kEV#Z���#0���*��"X�b�QDX����ƴZV��מѱӰ�v�jY�����f�ά���G�.h�r���<u��c��%#�<�zf�Si�}�����fW�ts	#�y{�6�W��^�,PgQ�2R���*�����リڳ`��!�3������zw�5Y����#7({�5�X�����+�Ư~�cVPdK��;Y�rh��>l�kH�LA{l��b��.'�=�7�/�u{�_Ƭ�Uz��UOn�P�-��өׇ��|�J��I����+�3!�RިY��2��ʍY�8�u>��]�Rǻ:^j��f�Iqu(���I��D�V���r9]�6
gZX�%8+�l�g�'��Z[C�U��-kuYx)WR���4�����Ǵ�~������m�/=��w�m���-�a����*��8��2r��V�G��.f�OAN���]"�蜙���8��{����6X|kQ���ﹳC��!;��R�����e��tު�vF��j:��f�W��9�a�K�W��g�L;0�<�$�#��[�W�Oa��z�H�б������5�o�]�3����8U{�R���w�R��O@����)�&��Z��� W\�unm�.�}w+��,��q����.�Y#1�-c<!GeӼ�0��<��=	�߄<�)��sN��u|��C�qvN��Z�������}�j���GyN���9��ѮV��ۻ��S�����1er]�^�'�]����3bo��Vr��Œ�`~��i�*^P��^�z�k�v�3k�̤ȉ>�F�t��Rip�E�����RHH��"�`�,���,�����7��~�R"��:Q�߽�?<�����N�pMUfp�Ëo���i�=�E�qb���N��K�{{�9d�/�7��$��D��m�f�m,�������nx��K����u�ɘ����ή9*��Ƞ(�x�E��Y�&�س�����G�Y�
�})6G�������:��BIv!χ��^�س�����idݶ{�:t�uƏ��F%�/e���#����ם�:Y�R^K�r��7���\0
��
s0{��-)�P���ǺƏz�K�ٝBTw�#��e&M��>\����":�I�+i�����5=0�̿L�f�K)�y�=)��3\��rݜ7���/�������У���P�gze�û�Cn�>�9|:EQ�	Ʀ�C�p���XZh3dj<�EVz7����rw@���XnYFe{n����p8�Ҝ3_V4O�����uow9^���$����R�N�=��J҅[�C������ö�̨�0~v2y]�N���,3LE�s��ܥBU���C����m��D������x�g��oO1�c]�K�}��=�v��'�i����ҳ� ��G�ݢͮ5��K�v#����s�_~�g%����R�N|��O���	���G���U�Ӯ�pۭ���Y�\K�����=r������7���`Aaԃ�;�,��է�Cb{�n/��Ϧ`�Y��ng�j���/��+�cЕ����M��;��t���C5։~�8�Y��%LB��r31@�P��7���ϩ]Ӭ���[ȍ%�.^�~��ʲ='���]��~k�$LVi[�J>�1���ȊX��H{Y�J�:�/�=c՘xM�Cbt��/�7ޭ9�~�8�e��W"[+�(C�R�]��߸WyXG����j�ߤɗ2�T���h���Ҹ�ϻ��<�QϢ���=Kv�ؕ��,�Bh�=���s���E ���מ�ރ�m�L�o��հԡ�,jY���~s 8f&uGh���vY�2���%s+���r�n|���~^����7+֠<�"��c�<�q718t��p�NԳ<(=n�y���RĲ���z��k �͘)MI���s�h�p������ԗm�X���f��[�I��:��]�\ة�ܤ�HK���h[:z�]�b���\�����{S�r�/��g�t�1���42<��$�f�r��j�#�BJ���[s���Z���v`��v|`��q�W��x�z�z{͊�ީ��M��@o.���2�5'w_iˋt؏VƱ����W�!�(uBG�����X"��z�r�ܜ��x=)M��z�L�7U�몗��4/a��m�Z�A�9���ɑR�<3���gΌ�[}����ZY�;���c�=:ޮ�P��Wh�kMi�*���pn�+�G4y�3{��dJb��ZbT3���=�Y�\�>u/���q���;�e����Yb�PB7��S��ȡá�/>��:�.)��N����d8��s��E}Dghqe�����۹���)*�ݨ��)�\dY�̱�켪�X�v���8˞��9�WǴ� ��F{=�lߞ��=j�Q"X�h�Z���yB��2�R���<o����ĵ���ƵWU��t{��a�n]��oE��r�t+R�\�g�)��	��㬻��O/��̓&G��/�J���*Y�R�(�r���ѲHC]-*����1�n.����,G2�h�Yx�s�7t��Xqu�Ӡ!y�M�,=���������} �Ϫ�5��~c��/�>�ۍ8��y�<�·>���I��8�!-�/���6��4_���o��H�ñzm!p�eY�=G���'гG;Bw�����PHi���{����� ����!�<0(a۩���#�	��s���=|�v���8;��3�]̖:�Y���a%"d($�`���\0}%�����|�S���:���p%/	�v��!�a�Mp_7n���O�|�/��S�%���]�8r������,KZɮ���,� ^<��t�8/�Գ���_41��O{$z�
f�^�:���a*v�"��+��r���^�,Peu��U�*ϸ�ɐ�.O��'g?�������%ѐ�1t�u�u沛>���Si����_]�;��z{�ss}�G{��^��"=��9�Cbc��k�՟z;�o�_������j����65���y�'��4Y0jS��B��z�Q`w��9�)O��	���{�CԽ���-�]4���l�)Z���M�Iq�.Y5}P�y�Ke`{J+NBarޫ>����ʴ�1=��Y�P��}TD�[���/)-)���/q!��u�؈�ݻ5_h���i�?S�5բ췠��Y��s�|���q�c۪һ~�p՗��yk[Λ�ܼȓ}��f?w>:ҍ��^c+9����[���^��yݝ����\֛�,����֨���}���8�-��X�2����-�a�����q�q׏��[�~V$+B�x���'!�T����<2�\�s�L��D�{��G��+6Z2{o�O�e�|�Yy���͚p��	�>�B�?ST'[��L��~�jv�sU�J�&�C�ī���9��nJ���=l�|��0��"L�;�]�ޙϣ|�#�!BE`f���[�:�ïe_��՟9S_��C�L	�׎^E��Yt�����Y����J
����.\���l���O\���3�,�tU�~'B�nh�ś_���XZ���%o�f/-��X�Ϋ-�0g۽i+2(_�/��	v�����mٻ�`�H���G���`�~��,��T���N������j�V\r��^3���l��7�&��D�Ğ���^A��[�t�o��ȃfz���+��U����m*��\�b��ү]�Q����r,/R��*nn8;��K	��ts-�y���y���ݚм۰ϭm�:��Ł����ig�k�:�� �+�pX�ˠϨra�8U��^���Og_�C(�RC�V4]��ɪ�S7jZ�  ��z>�7AeE�m�n��ݭ�r��S�/�#�j��:)繛�$�)�E��x�����,��rlPId:�Ry�أ��]���矬�n���ȅ�cp&�� �+T���C"���gr�~�~0�K����k�Haz���9�=����<��G��<�t��$X���.�.	Zt<5���X�O���	�����G��.�^�C�"Q Mo.=�ԯ\s�����e�ڼ'���|�ص|�X��QJһ�_S��H��WI�/��t�Nѕ9�����'�l��T�C�N57�0��e�B֚�u'b��w��~Do��]�Do7�"���l�Sl�OX�:���N5�Xz��v�6�l��\��Y��2���'=tȶ�j������&Y��b0�s�=��ޯ �\ytY�f��X��]�����Z�Ae���.��ع&�y3ܡ�������P��v:��r�ʌ�gtX���H%.J��f5�"��u��b`��T���v�z|���2Y�N)y�7�����i��J:�N� }Α�P��wX�K����g4�~�'^��7���D��*�2�\�A�(Gt���%b�q�������­;���o�	��I�ZnOgO`�����g�g+���z^��U����N���ڎ��\�BsQѷ&����i��,lp���{�t���|��ˢ���-Nʹ22�ʙQΐ^��<����;��ۯ6V�)�P��;�no/��+�3Yݛ`���\�����>�\�V^EV�8$4��;u.ȅ�(M+��R|����LqK�f��S��uh�L�����fwL	_�H��VX6�����;�0�0הmQ��Ϣ��(�F��ߪ���Z�1�E����;��K\}�2�bgV#������Z�[�3=��^1�A��Cn��g�1�^[�P눽pX�y�iV ��R��V���b�V7ݬJ5�M��e��V���Ӫ\�zU������N�x�z�y�E���ż�(��7��
���r2k��\[�L���/R��."�2򐺽^B��z��/lk���̕Ɏ�).Ü����ޝ�����K�F	�	ᔎ3L�9W�������ʹ�f�z}��<�Aɦ�iifu;��jP�)zg3�x=��#�-�K�]؄�EF�3��S���sp�U`�-�]�<"U�E��縋!ΨZ���}����&vJ�/mjK"��3܀�<yCF�Ė�~HV��:���a�}��;�qU_L
�5�B^�	���^lγ�;�����ý����{�
�,�/G�N��h�,r[E��`W0k/��^���ܦ��¨7�ڗO_ceNK��cX�]q�6c��\�g�e�Bh��W&W+�\��Cv�юd�6�"\����5�[��q��+%��a:G�����,��v^
�؇'Nz�!�|���Y�k>��sx�f��.5�BK��$K�h--˩��)�c)�1q|����:��9ڳ��נ��Mo,>6��M�;x�E�H�gCZ�<� ��SN�?q藮�����{��J��k�r��bVf��U1q*�{��L�Y�d���Ҧ24���M��k����^N�5>��f�s���70#q�D5OW	Yڳ�.�@2�<��w7�m��t��L����LV)3��=����j,�R&B�f0pII����F7�Z7�v�2x���,� ���Th��@�
ᶳ��5w����C����i-r�y�s[H���.\�y�WC��a�n�����r1>�Fϧڀ�,��\�1�|�z�b|D���f%��2��F�(�b��>�Ss[���6@r�Nq�k�3܂����5�v]B�zVR삈̭�	�|B�֯�Yb��x�ώ8��C�[q�����;ܯ��X��Я�pm{�jw�z��@HY _�~�]Xĕ�|�����o��z�s֨)�%r�����>׆V�����_<�76X�*�F���1���弴��n}I��V����n��(�Z�)Wn�Y�q��7{�Ju)`|�R�9���5�N�>o���W�l��^�3)�����z�Mw���u{�_t�8����Q��3�=Z�s���z���TΥd+���ME�;��t�d/T�aC��-{�ˋ�Q�̨������I�a(�>K�>Ih�����^�;���FC4�Om"�M�щ�~~�}{���M�|�6)�hL�#���9���֊��$;�H�`U��c�O��7{ګ���5F���B�;c�`t':���[�<TDi��KA��آ+�ۧi��&�U�V|1��׹�{ ���0�g��0o��j�멇,"`�+���h%�L��m{�#����}@��[I�]S��p늴��I���rT�lO[9�y�0�.d�5/���θ�u���I��-�B��c8�vr�Y��{�~���z�ʘ��w�	J.W�m��m>��c�y��nF���X�du+3��������!���u��}��Z�ܷ��ˑ����zsk�����*�I*)��~�*��sV�ۘIU?��v�7QezOu��6gM�(v��)U���=�V+�H�(�o��W2{�q�e�<'=��j(��W�ܳMB���ԥe�g.���4�u6k��k����a$��%�|�{_u�i8��l���ʾ�v]$��9����0t;�y������9!G/�K&�蚊}��ɛ ��Ik�2��^(��qᷩ�*vZ�sy�ڜ&�U}o	�W��sI]h�ņ1VɵZ��&2�@�0a/aܴE�̵�0�g4 ����uԤGu�:�Dۇ{;�q�]�	*�6�=qA���yt#�o��Ͻ��W{{`~�+s� T"�_	�j�]����S6Ƽ|^s�ՙ�f*4��5�,"ٕ�}'��v
����)#���-�Hj�nN�9\�e�ǧ!�pWԞ֣2���ǕmL�m�0J��>gx���;�	�&�5�Q���eX�۳�'E"1Ǫ^]�9u�<��m�$��wYv�t41�!��6�iu�/�����o*agM��"P29a���*븳C@��ޝ�G|���Y�b�����p;゗mf��U�m�����9�t;�G_�mr��<Q�o^cO ��ٗ����|9�X`{,�Rv�6�(���q+wI<���}�;G{x-</�R�V[�Җ�ͻ9q�����A�0JzVj�H�ut���s�a�-�x�
�#Q�6rt�[���e^�W`��ʍ�+�矫y_3t8/:ղ
�����V�Ҳ[�=��:��YŢ�=��F�.�7����&-�˛җlt���I�-����	��X-�b�E&��Aѱ����z��v�t=��ϲ��4eP����=�����f� d�'��]����R�Y{-�l!0��Yo���IN�Z��,�+v1�����NH[��S{;O
3�9.�QX�8��OU~�6.�����+!vS��0��%��0���vI|�݆:o�\���R|���g�ɧ˚�cG��VnSV�."|�{e*�DJ�Nx[��6����t�Ig�&��A��T�o=�j�3��ц��-�����Ӟ�{���UFg^g�G��}�p� �������b�o7W��.��Y��@�}:<J�xms�[|�]9�[��G�i�"�T��a�<��7c��=X�k탔݄)ڳ�;�:�������]��j�w�Ԍ��xh�;�OO�<:<��Giz��P�����PF����`nn�*��O��D^7��7u�n�	�ӭy��^?g��ƆOA׸O��-
ג���4H�27L�.�r�e1�+�Ž[J)�Ҹ���jws�g����~��pk�}��8q�z�7��\��gw6�� o�����I�-Nxr:��K��=���`����X����x�%�f��v_1�ԷR��4�й\T���1�����  �Pb
*"�����b��Pb��D,��0U��KB��h���ŔQUUQADI���A������DU��AV1dU�U`�TU�Ŋ�p�E���bV*֪�D��DTb�E��"CŨ,X���*���b�$RѦ0���1�bV,�h��Q�1�%E�m�mE���V�j%���Db,Kj�Q-�X��P�AQ@TQc ��8��UX�+Z#EX"1���EDEh��dF��)UD�UUb��Y�(�UUjԢ��`Ă��1AE����
)0ʊ��h�
5+mTDSUA(�U�,m���UA�EV��*1UDb �
8��V8K\8�
��TTY�*���1����������P��,űQX�P� �>���.7\m�b�/���� ���h:j�ܪ�O��ՏL�m�3m,����r���j���3{D�'г��u�"G���������C~�H��r�����<�%��\}��
L���q����Y�=�*��!v���^�n�^n�P&cDؐ�$���~��N}�͚��R��xk�fj��V���z�J�W�ߚvu֨0�po�<GX^��;DT��{P�,<�B��'Y��On��1ma,^ϟ����n�8=���𽱱g�@|o��Y^o8H�� ��]�y��ծ�^k�l!�i"xn҃	���R�y��:�2�zJ���xq?Dq`�N�N���b�ϫ}2�l1��3��A�ڧZV:&�H�������j�m��k��u��)oW���ڽ=/�{�.?p�	b��\]A|�w�^hV�BWn/|޼'ϒ�\DI�'��1S��N ��_�������V�ޤ�lqn�����w�5"�:�[��W�&���G����m�sBx{m!%va0�r�M��3Cv���a�N����̇>H�ۻJ�&Y��;���<��(oz�4����;G[c�6`6����<��	�w��'�m��L@t���|�vV��7��_�k��8�sҜhF˔���6�]̓�����ԧvor˾=ú�pf��@���^�����zj��\���]\6(���d���!��
Ͷ�'v�6I��3"@J����W9�>��W6�Y��K�,���;T.{�n+�u�x���\ԁ(k��=³�9[��}<��Dt�R\',"���:�M�:�k������ �d��Fr�f�:1���qu�B�Hb�Ӯ���y���/ixl4#����*�o��zܮ��,k>��I��BZ�j(A�(FZHV�\�k������{{��;�;�����07A<��ёY���U�N	>G���.ȇBp]�z`��{�y2N��/=Y�p�Z�x�.
ݩ;h�����E�!]���;r�ل�^�c9Y-<�}��d#^��F�T�x��Ac2^E��؇t��\�9�3:Z҅��َ҇t;JzXm���,z4��=B�����1�^[�}B�u�X��E��d;=^�}���݌H�UwZ���g���~jݞ�5[m:\�z\|&�g��x��k4�o;���d�7K�=�M��1��2Wi�=z�J�����tStxU��~��MWE�u�`eo�Z>���vD���2P�����J��b�öToop�X�SA3��t���9�@WGu۫�o,f��Y�[;݉u���?	|g|�[�A�z�]X�^췂�q,��֏%v�a����Y�t���Vw�=[�O��f��� �]��fe9�}�	��m\L�ɛ�t�Ӎ^�v����gQ���Oz�D��[��(@B�ۀ�i�Z�ZY�)����c�>��v����(�N��w阕��جW��Um�E!@�rf%Y�Zk>{���{W��^{��Ծ��y9�,Ʋ>�z{wǝ���0O�
Q�t�$9�KD��#���C��ywөE	��g;mN[)�>��o�=��bz�t6�P��r���xY\\Hf�/P�B�������W�h�E�������Ӗ��;�hB�p�D�*�9ɥ��]L�T�y����V[�I	v�z��3���3�{�4K�6�Xt�cy�o��Y��ĠA+��5�H�k�\�������U���P؞��7+�7���=�����.�S0�ED>�вú]�k���ztɼ	(#8���������/x70#b:ȃ�����xmY�ʹէ'5㞚��M�/;��bǫl"�����5ᮮd���Eo��%"�-�1�z��U`��w�Ȃ|9V"�*	*�Ң���cUoi�c7�S�Boe+$=�9\�<��x*C닫�+�g{$��.&�ު��Q�����	.�\ļ'V������W�-�
�W�$M�]Ǐ�sa��q��5j������x��u�{z����f��i�V$v�� ̺��yL�@T
���\v�ۣ��J��$װWI�}X�u�s'�Bޡ�χ:ư��!��nF:��xY���I�	�,�czq����I�� pc�d�J�;��%��[�uܲ?<��^P��/j����4/w��^��՛S��;��+�kS��d�?oǿo˽�F�����\~�s�P/��4x��S�j?XMI1���Ҍ�gչPVK��/U��S��Ղk�F�\�;�Ұ"��k�Èֻ��&�ᄴw)(0�\�+���Rj'_8��̇���V��?=�Ҕ����K{���DÃp��^4�UW�\�h_T$�΢[+Ҋ{S����3updq�����{�ap�,GK�*U��6�xu�+G_ޗe�TiI(=��#�={Z7��>�4un�"G6��UM���^�ϫ�����|NC-��.:�,�T� ��F<��N	T��n�w������0J�sP�5,�|���f�/�
t �Aj��Iw��yN�/�w��p���<��
��@�G�0��&A��o�npםx,�;1l�0sf"�T%J-�(��;����A~ݕf�<XU*9���هPs���2`�L�n�T�{\�Z�1u��57o�s���n�U�n���-.���o�����](P�c/�3����:��{G��M��zE,��?p�1� U�u�7��ղ&#q�" ����+��8���r�Y��z%_��Ճ��w�{�vKo��FFR]t;������{�"��t��
�_¸b��������v,�`y>��1��33�>�{/'OV`�JV�7Bj�SÕ�*�|��'�E,K��Ŏu������vL=�xU���x�p3��:e���?���0{��>�E���3�]ۮ���k�~OC���F��z�bb��h�\�U��h�
d�(�_�.9�.e��=���wɟɅNt�xyi͟]�!��5��^�9C�k�
>q�=�X^��;DM��f�W*Z�v�x�|�<��ץDWt����f݆s�[��^�ر�����S}L�ʇ#���Yh�S�Ym��X�s�,'i�,�xY=<�Lo���mVq��n���0_�{[Ǒ���=�Ɠ���o�A��1�g/�Wh=;}l�d��H���B�z#7k�f�Ds�����#Kf�����]_]�lv��3SJF�L���ҕ��:b���T(�Q�sJ�Ӎ!�'ٽ�G���2	��`T�dVѺ�g�U��=}��m9�Mh�;�����,�e��M�ݻ�9n�*k؊�:���}Z���6�Ս�K��..���|{�=�Vȯ$}J)\U�
���1�{ڭ�9/�f��Ft5�,natۨ늓9�L��b�W㦽�����ԛ>���sN����5V�����ܻ`��Xzj��s�4Á��c�FWE�&�a3ȱI"��ӱ̌Y�du�Dj�]��N�+�e����G���j�Z}��|]-��f�1��n�e��h��
Dt��!���u/��&��`��s�~@���.��]�rﻃ�)�l�qd�n�HR䮩����|h=5����	��^��w��V�.���Ĭ�s��Ꭶ!FZ������<��F��/s��5ڠ9��Ғ��`ؽ��[lv$���>k������Jփ~�
R��ĚY�i>\�Ok�����u��W�n�7F�IY�+>�v��+/"�h����b�~�vD8�j���#/�ܛ[��h?R��E.�r�Y}�\Fw;	w�y"��+,COR����=~�I�w��+2�Q=��#h	[��5�Z4wH�s$.�������;>8�m��E� ̑��n��������tb]��΅�'�gEz��Vǫ���qy`�\�"��Nz��,�˫�Q�V��l�G\��ͷ���{�.E��ۢ�5n��������H�Vk�!����m�Ry���[M�:�egAa_�s "$�>}w!k-�C��Y�'B0:��� ���B�Y���ġ�������~����.�F�kވ�ur�K��LN%�80z����k�5R�uK��O����b|D��[��5n���������2���r�g��PϦ����s��`�k�H�Hp�9��H�*\[�t�޸�=RuY�G�F���fS����z�}5�}W;�L�#�'�2��n���6�[����wk�5>=A����ި�M2�V�eӹ�:�<%�_a����k0F�x��1_�O�>�20J<t�x�E{�)V���}�E����6\�>��^,q�L�Vz_yv{�>�Y�)R��3��LS6R�l�2,��3��T�� �p�.j0�^�o4��BUZͱ���;�3��{�N6�P�k���#����3�G����D�a���!mŐ37��2KZ���Pre�=��s�/�����l�D�.�5�&��k���f�i4����w����v]��C�	f:��=yf8�o�ˇ����E������3ZI37�~���W�Ӽ2~8��R�K����X�~*���+j�^WX��闼* �R�R�8��]!�o\�v�.52��"��)\��Vۅr��cs��o��)�s<�}�W�ov����ő`"\�A,�ܻ���M�|�ו\��P��䙷�k�r��bVf��+����J~~|�[
ԕ ���J8�W6{H�U%�,�{.���}�.�{����:ȃ��]�^�����|�3�q�|9g������4_XD*��G�y�L��W2X�֢��V$�B���Yf[��S֯=�%��)5����3.�ϟ�Y��@����pMۃn��3���j۫�ۑJo���(���YG+ݕ�=R+��%��k��h�/P������q��H�@{��ɻ8����#��v5�%X�I��oJ�uܲ�˶�~k
>]E3�d�v�qם�-�oztk��#����u<��U��	�g� ��&����uǳ���q�Jo��}"�ז=�י�wEĜ6z������`�!�A��ٙ�;��}�q=S]B<��;5lC�5�/yڮ6����[�1��=�%ᄹ�T����� w����M`n���zgi����d���繨����|)b����k��KӁ �}�F�x��ER��:�!�7x�]ܭ�s��Si����<1z�sr�|N�>V��b��B
�}._crOazf���B��oK���Rm���^Ae�`]|O\�:�5��o�������.�g>�V�>������/�����ؖq����׵BM�3��ʓfS���~ֶ;��("؇)�p�)�k�zP��P-P	j[����>~lu8@X�6o{;�6�,9-g�ME4��(O,�"��w��':���Q��#O$��m-�u�}�s�{���.t�O��t�q�]S��p�{Q�y41f��k.�����l�3n��sK���3�Y�}�4�4������}]S� u.{�����������gΣ��3�_ָ��w��M�&�t�4G����A��[�S�u�� �"�z��o��Gi!̼�����Z�o�~��u�/�a�،'*�K9B�;��jᗰ����H����׻]z�:�������kFIbrR�C-$�$w�T�"�U3��c�Zn{:���K��	por$��=>�+�IH�ܣ�bOf	��IxgQ�r�p'���ƶ�{���	.H�E}��洼Y�-c\�U�cD?�� ��u��nS�lٮ������*(���0>�8�2��?��lK����r�<�5ݠw%y̵�*n��YZN��j�h߅l���22\���7��z�
h�BZ�V���Wj�ۈ5}�j���v>�V�Ql�u��#ͭ���(ʱī�jq�Lʑ��o��ִ�n���>Ӻ%�5�x����ӳ4���R���"E��Y�:�nr��+��'n�y~��%�c�b�d���<'�9�S����^�س�>6�[K1.�s��̝�k𽔠ѣӖ��Bejxn�K���C�6��_�Hcm�ku��A�+��������h�c�J�%<��������:oP�u0Ux�$֕��__T�Ň}�4���ָF�srxZ <X���>3�t;��=�_[���W
L��_��S�-��,\K�~���M��-�NH��MH�P�Nn�ʛ��joW��C���!/�#b��x�y�^�ӹ�~\��Z��V<�A2o���1�W)���	Ώ_�ݘN>F5^���n�E#��L���":+�������^,�=�v#�=�,�C{+����U�-�S�6�/���"h~�ˈ3��NR�o�� �k�u/��K��̱!�_U[�l�{�?b9�{im���;��r�����U�a�Ѡ���Un����`���5�[���B���IJ@�$��H@�XB���$ I?�B���IO���IF��$��B���$��	!I�B���$��B��!$ I?�B��!$ I?�B��!$ I?p$�	'�$�	'�����)���fi �l�8(���1%M��P*���A"T�IE)D�)@)J���J*P���	%JR B�I( �"*���T�)J���B" �D��R{j H���T���"	U�ڪ��TUP�J�RB!$�"B����J�UB�I!)*�M��V�!*�@�J��D�DH*TR���R�J�R*�J��AP��T ��D(T���D�5T�Thʂ�)I.  �\4mZle�EU�Mm*R�MMal��3f���Rƛ-jJ��F6�aR���5�l5��MT�m�����&���EMJ)T����*��.  ��(k)T2��VU5MMm��U6��jʦ�6I6���e��*�յ��+��4�c+)�JL�m�4��i3Ak*���B�R��)R�UJ��  ��

(\:�(P�B�
(Xv�B� ���B�w
 4(�
g\(t(P�@л�P�@
.��(P�B�
7[ij�Ҡ&�km�5m����V�P�*�J���U   �T�-�mZcb�UJ%m[f�h[j��eI��� e�h*�T�m�m��Z�f�����eUJ
��*�����J�PQ*��  N�٭+b�XjZ�cSY5B�+��j�k-�U�m��խkm	T�d�j�J����XP���*�ҫPm��Q��J���	B� \   �ְ*ն�d��Mlkm+R�h��h)�VZ��4�R�U3hKV�%�mYVڦZS`Х[dmF�ն�(ZK6j�[e+J�*�R�U[j��T���  9�mSZ�+V�4meXV[VڔD�F�)��[l&�V�bZ�jM���B��Z�#h�PR�i��e5m��P
$�Q(J��)�  8
�� �h�
�j�@��+ -lEi�d��B�,l26���H)%D%D�$��  8���ՀЛm�QVZ� 6l ��� *�1T &�ҥEmX
j`�b�)EB
�k"��  ��F��
 F�P�#(P(F���A@��1B���f��@,��� 50�*�F@h�0�{FR�   <�4Ѡ���@��@  &�CFM0i"&ʥS��`x�P�ؒ\�)*+VH�	�NABc���fo��������i�*����	!I���	!I�@$$?�H@��	!I�`IF		��C��Zxjf>o?��tS���!�W@�ʅ�v�t�Y�]nm�R��ag h��LG��4�[���^Gzŋx\6]Tn��/�B�#����_��L�A�w6���ыv�R��?1b��Ol�Z��hBRF1�*�B�auߞ�e�U�z4k-<��VY��vT�� �f3��h��xK��ƢsSM�f�r��W��a��Ո'��̌�v��t�T��%Ӳ�K6�M�*��s:N�P�ʂ���\����H�^)I�Ǩ�6m���t�����ګt��e�i:z~���Oi��Xg�)��Ve�M�z�G"�s��Z�	F2l
8&Pw�܀�]d��[5%�[�s6
�Q֕3rҥ�Ƭ�*�Va
ۉ�/����6d�V='-!���Q��YB��.a&�F���H��V��v��[��F�.�}e�wmM���n5Y�m-aZB�����B�B�7�����1�iݩ�:x��G%U�J��Y�)X�#�v.a�-i��m�����&�=/p�,7��Z�w��%K���)ut�IV��1�5��W�fCa{���G	��E�����I7%�E�	��S%9����ԕb��nJX�֨���w�"́�O6X�gX��G0��(|�$ed���4n��8�pM�s^�w��d�/(�RV�����ұdX�͹�W�������v��I�]�R�|�ŭB��(`�i���B*�͵ya�[��ܕ&�Է[f`�^Bm�nf5<i+��kI襈U]�ye���7v��{��0����p����Swp�$�Jk�m�b)l�4����b.��t)]�)�G\f�U�����{��m�B�8uɯ($r���[Ǵ�P�CE��f^K##�n%�5Xv��);���&�����k whIX�[��PG����<8�wD%��i�6u��st�w[A ��26���1a/
�Gvlr�F��$���\uI�eC��6Â£E�ÌB�g5tШ�ɕ����Mh;�E]�h��u��M�v��Dg`5�s-!w��>�H��b��ۤ�̅e�)S�2�����.V��g&=)^ÎU�yU(c .l���nYŶu�n�iڙ��Gؖѽ���r�l��V� �W�lXf��b��ʑKm.M���d۩��nfX`՘��U��Z�Y������P����߫�l�Y��0
�
�i<@��UkYA:�����$ѕoX��Ee�I��[	L(�;�(��m�Dj$�372�.�I���KS�b.�e1��YQT�E���6�ڈd�j+5
�Y�v�dE���WX#g�lې�Mx�&�6aup�V77w쭍!r�U��@`�����nQݺ`�>F ������J�6�(��M�{q&ZN�%ܥdY4� B�x5�9��pl�U�f�J7F�92^J��P�MSP�nTB�ځ�pfۢ��Y���jW�+Q߫k�q�f�GrG�R�y5E��h��n�7k�W�ssX3"�t���f��3��(���ЭK��lX���l鳣�ڶV��Zv��R���r�=���@�)���F��:�'J�Hl<so�pe^c3#ܛr�9z���Nf�k���M�:���@سVj<_]���D�(�� ��`�D5S`؜+rh�Ψc� �B���a���j��y��潫���y0nZ�����[�a@\��^�t�X���I��,��Xe��c͈�enG&Јk��� �l7ciP#ER�
��ɬ�ʳr��r:9A�r�-g,���ݕ��0�mFjE��YW�����A%m<B�@t��Դe�[���Ys�h�0��5Hi�uC�SY�UKC(�{��*A���ک�ʻ�J��ו��.ۭ�o����@=:&�&������������cX���]���1
	�p�M�r�j�"��rR�M�� ��x�Ԓ��-�۬C0'W�y���&<��It��J�׏*S�in�ҽ�F�)��.L��:�W�1lB][uy��5�~8-���L9���ݲ�*��^Xʟiц�K�����i�ݠ�ƍґ�1&R�Y��Lև�@�v�0�ɪJ��V �U�N)nӑ��V��FfeR�J5��]����ѽ��B��je��	^VP�L�;@
t���!+t���+Z�r���V��v�Fj9��^��wM��
Y�fQ�D:H#y�񩚳I�3S6Jɚ�ڡ�SI�Z��Ք���7��Ib*V�WM+73�ŀL퉦�.�mc��}��`�Ux��m���sIWK����������q��B���˺��x�D-!%��jުkY��Z)��6���(����M�Zt��f����M�k�+�\cF6*���f(��TWcr�!�����ѷ�3q�+��7ay%l��8P��9V3.�MJ52a���^i�0�p�Z�����A.cٗcc�BD)�H�H���Q�2��ǧh��;3V�.���m�0�8�0dݎ�܊U�1��\�Ց��Y��v3,�ǎ�05B,Mj�0jM^b@�R(3vi%�;z�,�YyqQ����f��Q̐DF)�����L�m���@ԅ�a��)覦��kIZ6Mti�t��{�!�j�$6�6�p:�$��"-��aK��jZ8N4�(�9������1�N<�6���֝�j<TٲfXrm�wS0k����%���VJY���"�kij'qm踋�!�5,�^V���:d;�@�f��cM�:2^S��l*�[�݉����cr�:��ܖ�,;e�����ص%d�VA5Y���T�b�ˠ�K�7�l=��/Í�M���J�,,��̦٥	eǥ�-�WZ��:̶�1Z��m�5����v��mh�Rfn��<�[_\wiV�S�Z�kZmV��yb����Im��E坫Sb�,1��z��p����M���H�hÎ=�+q�;��pn�2�p�;�Л݋&8u�.�U�R�0�������Y���tkQdc֜��h�P��.�0@�0Kܑ �h���&�.�*�5j*��MHfG0+�ҍ��B�7�A�+1cQKX��JMb�xDrʖB5i2���ɉfsA���*t�E{�&+�@�Y� �%��u^�,EV��h�MB�"XĦ�w�iv�3e����p^8��Q��b�q^,yˢq漥$�V)��	.:�$xt�΄�۽�cTn8��xn��1�r�{�9�Pyf$��S$Z�i��, �5Rd�q�fMgLNG.�����j���͙��@ݑFLEm֓Xj=��A�W6�ǡM��FƧh\!�W�����/; 5u�L���,�p��Su��5���Z4K[t��i�R��bU�7e�N�$U���y�K�JIv+TI�^)�z�%�`ܬ�X�H�XJFj�8JV�wx����n�iiK[v�(�bQc0X�b��	�[w�Ȗ`f��kDq^
�QIN�=����A��;�QfF��zn�Q�H�M�ٱ�yM��1�"m\ j�-X9�6kN�v3�r�F�Ƿ�[�R�G�7p��Տ�]���]քMz����Tַ��hЩ�$�O\K��
�Ki�V�so#%iXm��Hn5�S�>�>%�W��z��(��PZȨ��͒�*1�h�E(����R��(�Rͻ�t����(@ͻxifh%Q�B��&�ku�ʼ����(�e��pR�c	�6�Z�f��ۦ�Ah;ϩ�b9�(22�@��Hiv%��9�����n�6�a'	$��ϙ�C/�u��b�Xb��(䆆\�Eԭ��dWh�z�5 ���QG��f���u0�ُ `7�PZ�[������dI�$�� :(=ys3&�����T�;6=w�=�@���魡gX�&XrY�kRS�E'�r]�v�bC5��+i�*�{���A�Hя1�Dsz%<��T��d�oZ2��n(��V�(X�Zl�n�z�㫒5�;�M��45/V몤�mIv	����cU�����o5�{����w��i���f���/&O��f��[����n�(��}CG�2*��t�Ԡp��j��[�V+�=2�w&\),upI��dǌ �`�FL�sb)�Sb��'��&	�r:ݐ��u�u�É
�6w(�X�r�;EM�#�*�Ov���(��h2�8��j��̸�kL���ֱad5�::��j����,��)�fm��e���b�Q9�rԬ�=����/!J��G3�nTil��U(�M�QQ&D�6��yY-�=�IQ�L[�x.�R�Kd�goL��B��V��1)��n��j*����b�ݻ�/�X�<y��2ju�6�e06��.T�Qf	O%�!��z^1���*X��Ѻ��L�#�7���&�B$�ա��se�r���O#J����,m�[�C�f��|�$�I�pj�qCYx���l��9�f3yeQ���'b�]�G Xm���dd��wn�6���W��P��)��iq˽<ߥ�XM6֭,��W�X�w+��X��kc�Ci�n��$�bǙ-ػ�X���E3Jڼab�A7���.$��cEf"Q���]d�Tv���&" j�Ʀj�Qi�Z?k�e�CD���ȗ-f�H���R����d�Kyi�n���eQ��]Dp�"���YaY�jx��C|i�8���X,����ˊ�3
(k�ʊ�1��5�/�@Pm�F��'fC#M݂�������V�D|��9�1*�][Y(Qݙ�40�����-`"LiZp�u�4�͊��c�渞VQ4ܙ+LJ���`�N�#*E�t�Ո�Q�ǆ�#)��ӦX�d������Au"��Yˉ�M�.�l�Z���%W�7NQܫ�gP��"�B]�����ַpݤ�V¶��0j�ʺVm��m���㴡s��K�o,m�[[z����Iu����h��ܭövid�����+�[h�ۙ����ZXH�?808�f4n���ͭ��YB	���	`�ɰLŁ�f�-+�[OQܣ�m�yI�򮬵f�@�ҤGXT�&T�[y%�VUe������hZ�ai�i�6��I�m��C��d��Lb�j��c�0�B[�����d��R�h��ɬ�xYb��M�6;��bwJśU�cC�+$�fɱ!��c�6�&���8v�Mѕ�0G�V�0�أW>�*f�n�e構U^A5����D%K�7D�ӵ�.�n���ږ�.؟f֗hG���aK0�f��{Q�K6�j�Ԟ�q�c�Y�k�p̼��U�6�Y�f��7�A�c5 ��1�mf/�[D9z.�hO$�n�mm-*�aq�[Q5(%G[�yUxe��uV����{��7�;c���ۧ ���YƱlf-ߍ��I,T8ŕU�/D�@��#���z�=k�uR����E�k\�i5j��3"�^�2A�����+��2T+~:,�64̼l������и�{���]=&kïID��ʻ`��()��w�YOv̭���k� ��F�h%
q�3/c�5ٔrY�+.�tM��^:A��ú�K���7�V$dљr�rSW����d�h�ejʓ@ �ʫ&a[DZ&�U�X���݇�-���R`�[�`�n�t�G-	ux�+�YE]\�R���M��ia��0��ޥj��5�^ъ��Ė(��U)d"C�+*�J]\ޥ�X������Ty**cie��M�n^�K7Kd4�/*����L2(�̵�;���;�6o4���:պ�5��8�s�f��*w�1LC8J���TLX�زV�V�,,R�OazeGhл
Y�Q���G3��9j�JыL����(�0�E㐛yx-K%�7�p����Uf4j�ٱw �����Y�*��!̔��j&��jiM̨`X.�J�#D]�Y%��F�FTr�p����j���Pm:g��,�76^B�hf4����f㚌��mm�kJF��X� ύ�I淖�zsI�Z��H�3A�7J(�D��2L�{��WFڤ�%D^^+Df�Vkt�k1]ӷ�a�+����u�7�2�BY�˥SQu��f��R�ACE�f솝Zwdf����P�.ˣeq�H2,��e�5k��^�!ǁL��Aݜ�����D�up^�	a J��'6\����h�Ǒ�(��N��oOv|�q��P�2j�b���2n��{0
(8vn�-�y�Ӽ����)Ӊe�@K�[u6�5x���T��Ï���%��9��jU"o�.�ηbذ��Jh��v�c��x�Èѱz�)-�Q���I�#n�՛;be��3�T����m-J�m�v���xU,utu�����Vr����	<�e�g*1NۙT�yYb"�[J�TM����.dͺZcA��W�XHj���`�CdTwYtڳ>�1B�ӥ-hu���#8꾷�5�c7Zt	۹gf�D�:X,3��t(L�;��[q���b�9VA���.aٰUDj�6�p;h35Y�*��g.�0Z�EJ�����F��	4k�8��2�mܙ�-��X�kfӎPi�qM��+�bQ�f<�駬qʲ�H�Y���й[)KF�Rx蕥��y�In�-VH�1^������b�,�D�h�������۶Z(ڑX[dPz�&��5yiUv�ykM��T�5�Xp������ϦbܑM���9y`6a(�Yu��&��2��M��&�Ѱ�d���zw6�K"�%a#~� � �8D�&�T��oQ�E��u�m�n9#f���� eB��N��GB�eC��N}}�����	lӋpiI,&���l'�1Cu�p�v�������խY��᎒�8�Ż�q�U�\RGZ.�z����-f�6��]y���݌ܡ,P8>n�v����FeJ���a�.-ޖV�����LKp�Vn���\�ɒ��)KT�[.ܫ<�mP�Ի4ӵ}�Ǯ���)n%�
���'B�hQ����EG�f)wh�ˡ�Y�Q��ld�����K�ə)��i�"8N:��V�I��"=���0�_5�ܣ�cQݭ�R�Ʌ��[��:{�Es�VV�W��MPk�j����i�I��Õ�a�U�(�wyL�g��u�\Z�����,�*��A�v]u�ý�5��l*9�[�;`�icȆ\97����J��s���Q�i��q��c�����]8�Uz��n�nʜv �E"�v�Zƺލۉ�����;� ��i��is�K���_q$5bҚ�'��n\�U+�TmC6ԓ틑����
}Oc�Z8�3����nk����@��������V�zgl �t�`��9��Z��1��Fob���9��7��ޠ�R�@:@r�r��p�hB1p��Xn��J����dz�!wFp5�hY��X�N-͠]������b�c氟�Z��]��؛PWV�96��"�Q�]��ͦ�s �c�����>O1�;�M������������w�Ȥ<���8���M�Ȧ>\g,K.Ɓ��.���
�p�݈E���V��'/�y�4���m:Yx]K���m.���/Uؾ�ϊ�d��a�*�u�o���˾a��X.t:�TYi.۾
�MGX}e��i��bk�OyԨ,b�՝3(�[Й�dh�����\��|8Scل7�s�q4pB����Y���|B8��v۸����E+$����%����
 �<���L5��X�f��j����AFf]FW6˾��^f�:�u]�����smU� ����]���wm���Gqi3�y��;�'y��Ng�:�d
�M�r��.��㔝rԆH�ٵ�:��S�h]��:�)�>(��/�{�$9-T����{�Z��|q��M�p��pI^ch:��Ǹ��*�%yR[Z��b@�����Զ�e��X���%�nBb����˥Ck��B��`�LX��VȬ.��Y�Nd#����/s/{TFu���ϕ�?U�.[]��r�G�ni%q��TYO��ڌ�|�ty��m�2cۧ���΄9pi��K�qU�F����P��|��!��LZM�t���.P���P��I38���)��Z ��	��s�\�E��K�Y�xP&
֭QwEf�F;3�湇��zv��vi�бYPd��n�4��e��V9�i�+x���)1��Zq���3��W�V��gY�5�L��]QT�/��L�n��L��DI	[�#{�)��j�]�yK%N]m���k�m��Zs#ve�8�N�:��m8q:�K���庡R�QE�Z��o*S�dgu�[G{nM58UC�W���r.�����ooN�헆�Ҹ��$�+8��)_K�^���r��J���F��[]+�a�6й��n:
��M1��e5 �ΨA���҈^/����`��]���g�b���u�̻A=qY.9���<i�C�H�~t��җ����P%6�A��Y,+]��62�c���oM��kM��	C�w3_ukqҳӺ5����n�.����M�
��o�\a�m��)2.ƪ�ZE�V��5�(��܍H�ɲ�]�����tt�f7Ri��7�ab�m�c��
����/j�5��s��s��.�qN�|�XI�5�]Ӱ�CK�\u�l>*�Z�:tCЎ��m�/f���n�ʒ���y��g�L�ң��3sS���fP��N����V�1�ٱ�'�ׇg]���U+��kz�U�ł�)��D�w!u�U���W٫�vh��!fœ�9͹n�0]pt2����`��r.5�fgM��@���΂_f�{4�(�*Sw��Q���e�1v�ĭ휁l*V2T:����;���\(�듑����Уc#+gN���w���h]7���+�575�� j"On��]�W����)e�D@���U�Fa��*w��Y�#{Z],�.�aVi�o����@7�b�w����@E�w� I��U��u��ͣ*5�����3���g/<�a7I��S�N��M��,&_�gŖ����^V�W\�1����;,��j{����w�C��2�a���s��ww�E��Pf*.��W���AgnY�+�YlKҘ`�����RW8�3��K�_:��#uT�̇j�������ޫ�(��E�IA���nۨ�\��}]<���暦+d���P<;���oE2{jcS�k�t�:;f�,�Z�%խ�Āwd�z� �A'N��Y���V�r���AM`��j���qU^yfu�7'$-`�F7�q��;c�����|D��ʕ&(���7���ړ����&�Ysk��+�Z��7�.q3kJ9�u��9j[T��+xa�_s-���[׵�L-��Q�P�]�u����+�}:s��}wC2U�f`���m�MZ1ͮ�X�I�R���L�r��K�.�nV��7���ZW�GG���׭�	7;kMl�c�xb�\\���)Tb�r�	pV��bN�v+�;�\$z��ƈ%�8⣜���JVz��AI��b�s���A�;`��/S���gf�9�A��k�T�+x;� /sf���+�X7q~��^��e.n�3ڌһ������8~�[l��v���7���E�k��Q��3�*�u�@�)�<[R�+c����Q�ۻNuGj�\8�2��e�\j�d�[zZ#t�}��~���\��R��Z��_7�JJ�L�7�tٙ;�37"%h�!9ZN62�0�é�ʾ7��9Յ�Ԕ��/UwS�r	X�s�I�:[+ax���G���XyN��ڸ���Rd\�5�9���<�XY`99VH-��c��ܬ�ۥ� r�`���S)a����=���D�)���F�u=�C�ziW�ҙS$gX.*�9Nq1M.���.�An���r=qOM��.��A�p�껗��J7��4i>�Xon��s�11�n��$��wQ�01m�Gn,T{�[[s��\o��WC{��ƥG��#y��.��󝙠&����IؘV��ޥ&_U䵻G.�Q�<<�ꩡS�z�M�w�Ug��۶,�G�7q�#����u��X��h�Iuۖs���G��Iw�2�Jެ�ح*(c���ңR�g2���9�%m.MS�u�-����M���v���CV�hjRu�����\ee5m�m�.�:;��+ݮ'�Ө��;s	�ζ��L��V���⭘�Z�M�ˣ�e��H�+񔤲���U����Ǌ�r���m�E�m�Z:�eN�Z:i;�0T#��Y�d��zu��@e#���@:b����)�w����x����W+�#���j�<y��cB ������t��q{�\�{'s4��k���Ӌ����NGJ��n���!��8\���78Z���k�/����mdoQ�Zx�]G�b9R3f�wjK*��.��m�-���^)�8\s���]��朡��{�u�5��J�h��f*���4s�)]���|NTy�!����a��¾�*����][gD����٥���:���G��g�{sP(�I�U��۲{Y�N����:7)n��vu0�+��fui�O�+v��Q8���y�9�������r&�w�%�B���j�3�߼!����)(B@�#�4�D+�^�Gv�:V�ǈ��l]�ԙ���P�_�\�zg-
��<���~I�z�o'��FnJԨ�)��[ug	Ɖv�G&��'��''�VR�⼶w��6�bt(sC\���vq/�CMN�xo��&V<\(-�����ݢ!d��]I)��Ëx撟=ve��Y���r^�"���,քR��Έ�Z���ϯa�P�S��1�#�$;ٵ֣}h���	R
�-��r�VE�q����՝u+\K���4���n Q���nu��,୛�k�-r �V4P!2U�o9mm!*x�S�+���Ջim����{�������p��u�Kɀ���9	�+p�s,��j��tL��3���ӕ�,\���� ���ۥ��cm��j�Kk�̚�`Ӷ����@+:�KYn�z^��qU��5ۧ$Ӻ� �\c�s9v펜��z+9��	hU�\s�q޸�UZo�ј�Q��%�x�Uq�A���f�ҝ��9zM�Y�l��}v�C��V�Β��3mb�=�}(t�9�c���:j�~�L���S0t�wh`��G�@L�ٍ#��oB���w��Mb�]Rݡ4q33q��&�;;���*��2.��TŮ+U��I�I��,M{\����ٱ�6ȡ^��l˱N�LT�BI{�;{��D��QG&9mi�WZ��Yc�d����k>�C����}:��{��\V�\$�V�5�c��vqE��+rT�R��6+D�U(o2<��M�n�ktTg��!���bċa|�t��������+�1�5�����r`����睨����Qi8!��6uu�L���m�L�����ʘ{n�kR�M���Cr� ����k�O�S_W(�C(J�r��G^<yK3���z��!��?>Lߖ�>�}�ʤ�{��;�0`��M���+��WNz;��&f�TB��̾��&V�7������Vɏ��i��W!q���K����	�=p�-��j��!��mm�X�]�cr�N�#o���^ڗ�%��ɪ��8�%M��p!�����]u\���D�%9����sؗg���7�/0���OQ�7N�rS��hT?]M����u�K^��H�f�*�oU��;+1q�K��խ:8�g���\]+�e]�H�Z����(M�
8�n%�ˡ��Sv����w+��Ŕ���w��y�عط��b�3S5���*TW�{3nd�����qZ�8�y76KF���gP�/����*�]ٌ�сa�Պ;��Zx����fm��YQ-�Gd�g&v�m�6�d�v �+���S�pӭ�>/h��+5,�n��Z�q�2<�t:��p���Vnn��̐ƮD�1�ޭ��kM���a�=����=�W+���C�~GF�Bs+c]�GP�]O�t�1��,�-U.�J����x�,��\q�3t9�	����=|�p�b�9���>�浰�����zG�Y�Q*;�YXz�e��c'�ܾ�����:��Q&������q�g\���CamŽ	�Օ��i�c ��S����ti�(�R�y����N��X�Yj����|ek4;v��k͋��ŝW�n�Huz(�;�ZF�oz�U_N�M��Uwi/��Z�y�rw2��a�]r;�ڢ1t�:�@~�u��ޝ�X�v��7W��{7�O*Y�TzƋ�-��)�컍������o>S[=�$��#1�'���+4ms�����[�3�.D�i�1:�魺��`�R�{ʟ���~ݶEqV�.n��I���SSՍ�K�mI�ڵs.ɪ`鼅���	������*����ٸ�W��c��I�	�˺�)��	��B�>]��M�Ht�����fR����ͣ�ӹl�����ƺ���=y4e[�ۃa���9�()��oB�U���t����Υ87Y�Y�ƞ�q5��;:T��s�}3�͹���'�m��C�Yy�K�Լx(c��Gl�p��)'�[�q.����l�7f���k��D���k�0� �'�R!����߁`���m�uc#����o�7�In�C�&^]�Ѽ�]�튙�R�2T�}�k���e��p� �v*ȷC>�V�Uέ�q�|q	:�Mw6EV]kR��յ��w�q2�m��Oʘ��Y�;�8���t��l�{�)��ū(9�jT~j�S(f�z6�y�O.���3q��4�e�eH-�Y&�����*�|���s�0Ʋ�X���w��wEv"��h���eW��WG�\���q�[3�����v��]m(����-!�͘sv�Epŭκטµ��4�p���}���I��y���1�mԡ��T��32�ȩmF��@�t�
�м���:8�`v��u�xm�"Ɏk=��&[�{{p��n9\����5v t���l�Y"rheKr��Q\I����p}�o:��5h�j��)��tc�I���W>�M�o��Q�U1��Dz�����Թ���09u��>��&�u#u��bጴXTz�;t[Ru�en����x�4YG��j�ITr���4k\�\c�	�할�簖o�m������N1�`���;�{���xn��똎�΋�9�$���Ƚ�y���GI!��D�lM�0)p}�0v��N�;�������y|�u��܏�[x�PDG�]��N����
�~�ۦQ���[Ϟ�q��0b�]��͡����ĕ@�kt��ܱ�&tX2�L	�wSM�^�࢝L������WX8���$�f�ȥ�]�gWt�Fd�Q<����-��n_*�S�/��y%�O���,�9�d:Opo�Js��3E��ם]���h=��]�� ��Ԓ�[&k�!�%S���!
aZ�W��L���(�0vۧ˯%��������C#&(�U����7�� �yJ���'U�)gJ�yi��2>Z��K��(�VQ
ѴyZI�2�$WF�$�%q]}�.H$��E��Zޕ�"�7�ǲ���w�D��`��3�Ir�G��^i+�|=���=��x{�U}��,��9��f��Cm��6+��(�]��u��ںS-e�F��n�}��q��Ʈrȧu3&��up2���(Ӻ:'#rR�M�p�������u�����\6#xnM��U1�ل��OO����0Ђ���:XX�إN�V/V� �[�"���͊)���Ь�xŠ�^K"L��Պ�X3�I̜*MyJP�6��Cw���|�Y�Ӵ���"//� �r�r�;��:gP{Y�&b���F����|s�&������S{0�ކ�kw�!��
'3�XCoj��whG�e�ɢ���GA2h1k�X2��5.e>�G�z��ۏN!�wV�,]b%���}�W�y�"���)[������o����ŀ{��cm���\&��f��/Z�J_[2�W1!Oa�6���bi����[x.��wk�X�et�eIae��0W3eU}7�u19Ix0StV�<6s����M8���jc�2��z�%�R��{R��I���N�q[��Y�l�����L�۝zr}�ZͺL��Y�֘��P݇w��"f�.��[�El¢y}sdb=�i�uL��o���wI�7uƵw"ܝ�q����,u���N�85bjԓ��
��Y,�GhX��S'f��WsZ��=|�9©m��t!��Ѻ�+5�������h݋M3x��l�,i��;������d���M�{(�O�9�gbVo�Vt��\�.Fu����G6c; 
�9m\V)�v�*/�h�b�P��(9�CK3B=ަ�w�I�X!��eZ�{ӛ���:ET�)	I�D%n�e;�$�eG��fB�|�΀��� �-з�*}`���L�m\'M3.]��K�[,5�u>ԕ� �I��5�����D�)]mk�؜JVu�)��������=����q�o`�g'R�C���	s#{�Ν�/qpY�U�8+4���XiZp������f^�]ݮ"�]ST*v���#t�Y�\Z�dVe�&�y�����"���J��M���d�C�zj�f�彤��(@S��%��`O'o�[���I�ݗ
��)�QIi�;�]������blWˆ�x�w����v_)g;8���ַٴW)}�k:Ø9��b�M�&ɃF=����ڗo{\6Kͩu��k�L��ל�$'R������*w�SE�6�D��;�ޕ6��-����Hqhrx |;%j::�s{]֫9�9�B�(����;S��R����v�Ӕ��m4�2�bT���\j+d�Ya��5e ޺�:V`-Nj������}��
��/:,Żb�-������ޣқ�lYm���r��Y��[{�$n˧�h<�#�xyRL7����-m��[��Zw|�s��8�W��i������޿��&��IW�f$�ؗݚ�wG+iU�t�#RrШ�$޹��ƮA:V�
���WݳV�d;�3aZ�|3jf}�#�6%Z��(8ζ�f����7xF�rt�,+���L��Nh�Q	]�*eμ$�(,e�w2�\Ij�E�*��YZ�@ۼ��5�G�n�`9��e�&sL��#Էm��x�/q�h���/�ݫ�ݸ�k�ӝ.jEr��05�r�^.��a؛*��]�VN��ۧ�C����ɷ�9���37:u�
��T�ھ�F�QSI�����K�US/\
��j/��4ro#*��[��`�(�I�V_-��'�B���/��l��㼲h��#[ڒͷ�]���ÐY0�o[�����b��P�}{՝v�p�c]λQ�o6m,цQ�{o���J�.�6ά�`�7�4U#|{��'���8�U�%��*�ѷ�@��]�����X#1��p���j���t�%Z^X�Bl�'�t(麌K��KQI�]��R,Lʰw��o2�o̧�6��������(��Z�S��m���R�C���d=�Z�8�0���z�j�i�������P�B��+t�:ޫf�g|��5妳Z��f��G4�F�#[74�9�g�h 难Xm��X�J���U��LM��I�h�.[<r�Al�L���'P\t��w��XRS�[V��$��<6.�gi��̖��ʑ^`�5����f`Ų4s)�oq���G��/P��\��e�;�֬���M�܄��Ɯ��)�F�"����n��ؠ��4:Yy��=���5�,="J[�s���j�[���2��Х��+���T�$4����zn��7ה�/+U�YS���Ά�ef���m������p8�4!��-��i��l�6L�k��zb�I�\����n�e�+;�Wa쐼��y}��s��l�f5�ݐc+z9Rf�ݱ��W*�b2�p"�n���k;����/^��현��6z��(���0���Fwa�U��E�c�/���$5��Q�#�;d��ʌ��}{�����
�j4�rg:W�^�muv�J����mc�����MEu�~����{.��Q�4J�[A]��\���e,�E�懃�7�������U�T�2+y4��4%�d��̬W2������re֎�9E�`6O)tD�����k*�:C��;=�h��\���<z{x�L�#�;o/9.��d�[8��q���4d٤�Y�:dG/���P�ŕ�ke�EΣ��ݺ��lQ�H�4�p��&�ѱ����s�Vq
_l��,!����e�GG	��gYj21��BJ8d�F�,6����pͦ���5OS)Z˴��<�3j�L�!V��{`Y
�r��u�ɓ�YQn �`3Mu�7����R�}}w� 4cN�-�|�U�8.,`�t�ɋ����X���	j��R�8��35]wu�dN+M���)WR��&1k'wD:���Z��Y=����Hq�%�˅7	�j��'N"����i���FE&.�۱�5��wbq��xJ��n�#�[M��@��Y��(��t�g-z���Nͮ��3�
:Ght���=>4�_-V�C�Q�2�����J4��� ,�ސ]���DMXs���Y��JU���{8v��WFa�ſ	B-���R	�&�0�A����N�%Z*���8�ц"�Z��(!�����d����Gy�3�.Mã9a�%���G�󆲂&b���W֦��!�����=i67�Cvx��F+���M�`�[Ekc2�v���Ѵ;�35��D�uG/N��yL�ǋʳ%l�V^��\��6�T��qdԙtΊN�4��[� ���r8��ܕ̾��]!����$�̻���eďn=sD(*\��n���,Y�R��Ab�4�>�K���]	!豠�goS�˴�$,���r�8b�-��Z�u����돤�:�7���j���Ş�k����i�b�����p\�Zӗ�Y�Lz�$��z��p�b��c/�� �tu���\�.��&�oU�Q�9ܬ�"^ge�a���)�c޼�;	!vK�<8��E�}=SP�ՓQ����6�%V����{2�Fe�,�b�.�+76n���Cg�|t�k{�Hk����n�aꗇ+EYTP��P��b����kYr�u�a�Դ޹G%�eA�u�:�!��̣S�Ua��AO�P��v�4n�N�v�Xh}]4e��U�Ra�r�5{R�1􂢬�v�XL�8��0j��Y�Yk����;mi��ͪ{Ioa"��T�Fm�!՛�7 ���Kj��G��+�r�������1��u\�� oy?s�����yàzr�L��]�V�mԌl�
�;y�����苑,˳�3%.X�S�P�{.�]�m�mZ�LM.�.�]G�mp��nȝYA�� a��ewv����&�f�;|�R&�j\�<�j�S8e�K�!�a������C��.[KKͷ�E˥����ǭ[�ʒ2���l��-�@�u���sR;��9��;N�{uW[������ef>�5xuC	����SwMk��dˎ��`Ԭ�ζ�<��]C��Eݷr$���t��E�hX�bʶ�1���Ƙ �0�x�����o9���R�Sܴ-n ����5m��#*�w�w�C#b�8>�$��4V��&��wz��k���h�����؊8�Jf[���<�c��,�ףu]�`��e��<���_�v�����V�ƥ�:Ιn�;yՉ�T��lW[��J�{�I�O�e�s:�u^��nɮZ*n]�|�#�R���䱉�Z��'n��/C�^SjPe���A�q�X�\��K�r�h��G&��,%%���2����y��t(��XՕ�f���!�2��Y(辒�;le*; ��#�\BΤ�&uK�e�.�M>�����{V�!��6�"�{�Ȧ�����{Y3�eWڻwA6E��Np9����4��e�]�ͨ��ϸ���bUĄ\+.U���E�;��l-(�m���|r�����+3�R�]���koV�0���[d,�lm��%J���aeڰ3��1̲�=���ʂ�s["�����h��᷺�		��� C��8 � ����}�<6r�<���{{:�]���Q%�����nЈ�۷cB�P�	f��bn��+���0�]�>ˊ�sk�CSc�V��ookUۛ��尝=�X)�߬*m�����:���$jۖI͹���W+�8i��ua�%���vR� ̕\x`�s3Ʌ�#jި%`j��������׊�u�����OQ��:��̓{NU��:��㢪g�[h=�
$�ek��A�i��mek���eZ�z�=�����D��[�v�S�o ��o1��T�s5���6�n��zۺ7�����4�^,�:�\���fR��;vT]���t�ȕpR��-Y$�5�v
]�:�ń���<�1]���D.��Ž�J_V;w�.-�NR��2��޾�׹�°�%��K;�W��u Y2pUb�&���Lr����kkj(����pK���֗|Bm��Z�S-S�\/�*��M�9����,��ŏ��t��XK)b�H��l�-�^�:3���(lָg3f-v��n��.*0Y����k��U��.��e���;�;��.��ɏ; �S#7�/iH��|��թ%os��N
�Y�6<j�S2�V!�6�Y��$V�S��a������NIA*��b)�\,����}s�ew&�p�Wa.���Y���ٛ��{V�墨�2�1���9%���:�[�҇<����<M�.�γ�3k�I}������!{gU����J�kF�ʲ��C:t�b)��H�pSn�c���ќ�2[F�Gӌ�.�u@GE`� ��c|�����:�:���#Ꝉ*��W3��.�gIC�m�6ZF�0�O�v���1��P����㺹@n�'t�����"�w���x:���1JN�P� Nʵj�¦���+�2�t�Ӄ�p���*�kA��j���{��g�M��əb���nW�a�#"�0E���y�q�!�X:�L-�k���<�wj���nk�=W����[����7�>� ���l:R	��>�ٶ����D�a5�):�u�kZ5�Qs;�2l�y��V3F����J��P�R���!Wj5bń�;wrr����*˾S�C���[�|V��[X�ӂ�h��nI���p��kP�µ�ǽq�X�h8��Eݢ�c���]by.s��U�CB�e�B�2ak�s����R���jS�{m���hme*R�������Y#`mNr�؍���ð��D�[-��(�Y��\/�']�ى���+t~�Ge��M;c	$�x����b��CPH��X9]����ס��f���]��.��uͱ���碟m��8�p)$FJ�q�TYsǝ��7!<���T[�n�aK\p�ˮ�����ݧ7D�¢����p��3Bi�t�D�6a��w��KS��n>L�xl�B�Q�4ۤ,�_-�y��O(�/��[�N�F����`YP��6�b`�L7�,��Ty�УÝ.�#�ތ]�\�
�^^vθ��b�\��c���c�+�k�gX($�\]"E��I�5�,��C?i1۫�aDͫ��I<D5��Q|{&�`��6vU[l�4n��ž��dz����x�5�q�� ց�jH�{�#ڇ�q�����6w�[����!6��2ধ���e���κ헒��в��+��e*3�g?�@rA��ss�#�{(�;���` �cԎ�#o��#+��.��tJU�Ddu��	O_Jڹ�E�ynK�]���-'p���é`��䡮J� �PR���av���:y�Ex�e�yq�0�:o{V7�+)ӮG����w�����07��5$�#�4b"Y��Ǖw�,�ڭn=任y����y��nHT�n���%j=��{������i9АY������w.���W"�����ÂGx�IFѷ}|%oe��"�j�}����ʆ�1t�9�x�1�ݟ^��[}�*�R�5��-ti;�ͲV��V�:Ό���Ȯp�]Y����컸3�d"�h��x�41
yh���a��7�Ԯ�;��˲V�Y"�e�qݣ��}}v{�ɽ���%fa�ج���bz(B�7oZ��3�y|��B�S㐤�V܆H'��u�ON1uƋ���ۣ�5T��L��)K��j��t���{����w^̴� �w\�)��vѼ��+sB�ѓ��`�����U@S�r]F�X�,a��,f���7!�k�K��`Y@��-�ft:{�{M;݂(7�g"����	�6d^�ӆ��@�@�e�Av��zu���yj
�sYÔ�ݱf s��I����B�xMa��j��A������F�#�������b������J�u	���=��y{#�Ȏ��l<]ή�]%�M��jcn�@Ů��*gwo��:�{�dY�:�o%-�[��
땼�J�zi9�L4�ER@��M��m��.�Z��%Ȣyh��n��WU�c��������WQq�qʫ�-^����ڝ�,�8���c�ҭ�%�)Kz��u�H�Ү��"c��ъ�K�k�Pj
QUۻE]��V��������_��� 
���!��
�������i�ڳ���NytaU�ҡV��>�3������7���I"4���%F��g�V�ٔ�R*��Vf���&E��1ű�6+�K&�6Tv�oj�k�����*Մ��]1�#�뷗R�p�cu����z��Rk�Yݮ�j�w��*q��o���>�����3r�m�o��=���ܕ,�Y6ek�%I��A�͖��@�=���ʊsz�0�U�3׼y	�c�u{]�E|�r��N+w
yM�8i:��=b{��H��ѷ�O\j���8p���58X(�>�4b�����ij��w{���;/e�Ʒ���V��Y�5�x�N��巷��v��p��g[Ѓ�+Ru��B�V�Z�KnT�6q�ޢ��U:��w[���Y�ķ�̌�o��<�-��2s�'6!���ꭝ�����*]�%�@:� ���QR��#���,	:���w3��s��O�)5�{
�Q�����
(A Q_�~�!X*,kb�u��["��Em�֪,b�B�h���B̥+Dc��T��ʹcUX�ب�5j�P���mF��X�1�TDb�[�UA��m0�D*�A�WiE+(
�Pc�U�([Q�U����Ԩ��I�Q�Pb�F!�����q�e��mEj�"��7w(V1YZ˦�cmn�rւ�±m�JԌ��щZ �S�ҩ��Jj�"k#VV�+mVT�"�%B���[Zت��2#Рŋ���R�,X���Z�m���cl�Z�Ji(��AX�"��m�����X�)b�)U��j��R��EX�J�ѷ,ɉ��e���i[-DFض
�d\-&5rʱm
ZX���-j���`"���6T�T��K�.#��~�~�lRa<���ג��oJϺ.3�zuH2�sj�>�����;�ݻ�0�y�ʝ,�*�4�rDr5�s�����y�D?�����.g?�;]N>S�ߟ�����������Xz�����q�~��pKJ�5Y�<��&�.���,�4�+�K��f��n������qW����+��5�htU3SE��MV�jH�Q�NÅb�̓�ޕ�> g
�C���ͯj��b��c]�o�q�/*�K���U0-�s�q�;�C��V
�;Ȩ�3"���=Z�2�+��P��y�iu
y�6=�Pp�Φ�v��L]�����j,]X"�\�iaF^է���K�a���f*30ۊ��z�f���ט�7j*"���d�v]�F��溻gy�e���v~>�BO�1��l�ީ>��3+"�������	*v H��bT�0�ם�zwNƧ-+�ϪM0f���оB¿(�'S|]WO����/�\0�h���m�}��~�/�)��06���:���Ld����4�Ep��V�3��uZ�s�|)�d�����~)*ҲC]b�F��������sL�%X���v��w��p��>�82%�C���unـ�����K���)���!Ɋh��6>�Z��[���]��3�w��S켻�0��O��&�-�ҡf��VPT�	�N��ý6:k4:f�1�E!7���	�"0����WgZ�mD��&`�&zf���;t�n��thiY��^���˵yV-^����@"$��~�V�I�^a!�1�=\{/��< ���x����\��!�^bנ-�Y�U�o�{d�P��AY�
�Q�!Ga���r����65��IbaR�͘&5�\٭���d��� ��`a`>(�����W��4������T-H���;�6}Ap�]�f�?hW��w�g�wrA<�����9n�#�U��s�����VqI*2*�l���}��0�/�̮�L.<p0��.LW�&��P#�Qy��rZ�Ӂzk����@��xae;�cw{	ȑHR��D��j%a$�)s�o*f�>8�4�/g^�3��#9x���,��wh�w�)��Q�u�D�S{�3k��Az�c�Y�nd�%z�`�v�*��8�(&��8b�-��r�̡�Aߣ1�ׂx����QUd�;Hz���+Tǵ#j<ҭZ\���7/Xј{��6Cf�X�:�s��R<��;��Ut�j�s	W��&�E͉I�$7jN]����peC1)�pI�:���o�lĶ�z��9V\3B�p^F�R�
��û����Y��"98�';�&�=\�kpmJ:��k�=U��b�W�:�/<7��{�B"����f��LF5����W�s�x_�N|n}��'@v�cSG��pxC�*>�f-VFƹ�#p\���U�$��\{ZV�O�r�����}��Js���'�y@�b�(5���_u����Ĥ�A�B��i����Yڸ�\�s������k�l��:Y��ʴg���������W�2�ܭ�y:�[��y�Y��^H���9�C�N`���n�0�����'���ᵃf��U���J���9�E�Bí9�;���Q+1M�'cQ�;j&�{`1vf9F�=xF�ׇ ��u����x1J�4�gM1��O�!�C�;ܻ�Qd>w��_7�����da�aחT����n��3i��}���ӷ|��f��{�,J����p��z&N�|�Ҹ/��@��\V��I��7�uJ��K�~�NNs�r11J:S �]��۾�bJ􄇕 �Dp���k��,c~�u�Z/GX:�=��2����5�'3�
yL�-ۧ~c�w2^+�lZ�.��.X.�����&�{��8OU�q��؂}l=��!�*�es�����pr��~���A��ԑW)2��lQ�/q��z�ʕgt��'/��\�FKi�߱�r0l���K���(�]tʌ�ojsڨ\Jȥe`[�o�6և��qN@��t'`;��.]�5У�;NX�	NE9�9˩X	{~����=���Y=�����ጟ������2B�[���*,i��/Bv��$(�{ě�GhL��}�K�����ƈ���ۉ` �.$�� >N�\��*:F��\�]48g��{{�Z70�y��H@v<��������z�NXB&��z�R�w�
R.an�EE��ɷ��j��L=n�t���&b� Xf+�@J.ȭ��|�����ɢʩ�y�{3+UG����x��y��vܲ��1�ψ`{�qP��cu�L!�^ ������t�~3��_��-�oR�N�oc�^{����c<ݳ##���}5�V�lڜ��*�(0����K=zVl��+�W	�6HطU��۶�4��`+�2R����3<��[��r%2�V-3�ؤ��)��/�%k�s"��E�Ö�8|E@��3y�
����Q8u����]�5�gW�����S0����G'CRl|he��h{V�*K��6c�Y��Z��5B�qf�Vp�^���T���j�f��衎�*>"�9�.�\!ˮ��^\r�M�\��R���[�A��"�)%���m�F��	�Κ2�H35b}�!ƈ���S\=_O�{d��[�q}��|J�Z�#D$b�M�{�q���ѥ+5+C6�l`V�t�=;Aj��ݳ�5���(�P_�i��5�\2)��b�,O��c�22'QX�l`�&3(���ȣ��棄���`U Ԙ�0�Aqc��]k����z�̂�r];ا�%�f���>��Z��8�/�V9kL��c��o���\eצ�*���������V��ӓM�P�Y�^yþ��sh#���I��;�0�����4�3��=������N�`��eB��:����L�@A\��;圑>\m��G}HQ�b0s'3���'�Q��R]1N4��;~��P�@|�Y������s
N�[�*�d�o^��+���O�_r�ֈ������@�z��}��5w�X'��1Ң)�m�^���:�;�+�w�����%B�؎l{vg�ҋ��z����l�[���}zLrq��1���7@�%S"-[zI'�۝y�-�kt�f�f�,T���7];�nK��^ag=��s���v�Ѭ���F�V�g#Q�
�0d��h��RU��,/y�9*���&^ZՈ7B�&г��\�x��I�V�nY�M�vWi��@���,�Du�_�ѹ~�,ʽ��4x�3�ݨ��о����9�UW�잾O��i��~��TҸR,�46}���u],կR�p[����5�D<o�u�'��/{/�$|]�ݦ��P�����,;�5dN�,��*�}l���vKe�p��5��7�����.^v�X�A�{X�R��K����Қ)���	�r`�ۜ̈́N_ku�$�7��͝�쫴 ƎT�e��Cý�p﵌Iמ��c3�#��(��Jٝ+�v�z�ݡ��='�I<!)ٚr�w�x�'"í8:5�f)h��ꔪ�޲|e��ɷ���Z`k�J���R`\��(Q*Z�,b��8��:gT�֢�i֘]ʊIN��8ѯe0��-��]4�>�1�
�;�ʠ���z���D�4��F������+6 ���M3hQ~'�8Dx�+}\o��/�r,M�*�W�U�-oyl��JKS0o]�����T�:���7T�%T)ΊU����`.��.�L�%���F��bٚ¾�U�wIs��ɋ�w:���剋�UkwE_(s�Ӷ�ƳW�46��4�͓�l�jv_e�t�5��\=��<�\I��VV.֠2�sw�;��C��c��E�뼥'N�:<�r�iUu���d�5�EE#FۿsN�WW��i3]�0�r��u�|���/VE�B{wPI&�f�K���T�X�Y����ҁ�N�#N�g�����'"E)@�I�>'F�v��o%��^wF�.��9�3h�`�����}n���S;�!�`�ޭ����w�䄷w}���<)�A?�\� q�;A��2qf
�O�Q;9�$_���c��I�4;I]~�UY����=�;��`�A�|W���:�tl��/�c�������6����1f��D$%�ژ�k�z�9I�lF5>��I��0���+�I�b����S�n)����*�Qٵ#��%<��:q1Or�皿tϸ���^3B�$n�"���#�Z��FI��잁�nb2c��x_�^~��Bm�h{.\�O���r�=UUJ������@�N�w�9b��Og���pt�bk�L��c���f��Ft�Q�j�����z��J%��>�8M)���.��j0Si���u��5�`�c�8�_���N�۪��y����n��t�&y�<�]�m3/��c�����1^��nʢ�Xo��2�Q�#*r9v�<�$��I#=p*��>S��fj#�q�o�wb�Ff9/�l�fv��UcY���G]�c�%{]O��D�N�}@�ݭ��דg�_i*%Pf�������Jw�"����GAk��M���O��𕙜��ey#��m3��V��$t}�o���MMB����i)8؈,�Wݬ}�%�H��n�B|^���Iؽi6��ZVpc�}`�쏁~;<AWy�Q��z�j��ފz2�x�P/�jԛ�S�B�b�.t�A�F1N�Ӿ�z"LM�-���Ng�����d�] O�ElשӉ�6܌��&Z��w�'�As�*�ojpj�q*c�+�fT�^��^��^a���\g�/�7�
+=�gx���HJr0[��s���q<�d�����%������O,�s�+�?.�g$N��D�K���q��W9iӇ��I5uM��'hӢ�<>��t�����t�@�a?�< ���E؇42TLP���9�F�C��_f��g�rJ�^��9%�qs$@m�'������1��)�S�������E��N��XH�����Q�C�0�ވ���Z�%G����������N��ZP3f:�3d�9�B���b��v`�*�̗�N̾�K�]�Sd;���[PK[tj�βs��R�ot������c&H�
{�D+�9�[�M��Q�w��ʤoב���g�P��;��[EMV�ӿ�N>�y[΍(qN(c���ƥ��z�K��,�C%ÁO��ۜ�u�U��E�;���[b�r��s;��^����6�ɩ��u�����=}�����1��j��WWB�����g9��ct�ۂ�����g$E��$������@i�0&�V;oc�O���xZ�Ol����g���E���YD�9J�\���$��'�4ж�r���Vq͝�J�nj�to���gF �XOg�^���J�P��E��*��移:�a�K�)�k3`<��r�tش�7Yj�9�rv;�+5+C6�o�fc��P�Q;�q�k���Z�`��0��M%9�r�r�i�NW1B�O��c�^̥a��z�~��)�����q'˅)�P�Cn���
X�t��/Uf����aN��q�F�N72�l��x�9�Eko�J�ʋ�Ф��ÿU�.�`���ю��V����;�Z������aԶj=�.�U}�ODS����{�A6/N4k��{SKy߉O}x��n,,�)�\;G:Sd��G�)��/-B6���2,��/_z�����P-�X`���v�Ջ��T;I
7*��7N,T�\v���T��K����͜�wJ�.�a �;�c_�"�D=��Z!iCM��W.Sl�4h�/��v^!
���X�#|V˄��^�-
�� x;�\>\cA��AB��&?Qa:�{�p��ꁟ
�	ΗAFVz�w�{�[��#a�8.)�vv6q{��g<b/Ee��>{q�Ū��u9�50-Nxr�q�S�\8W.8:�7�Ӽ�����F2�5��p��s\��"���f�w��3�U��l{v`�Sr�w1D'lG@�9
���������j�?L0�:Qk�GF��x�*���Xޕ�+��Dx{ϋ$�W�J���.ͼ���T%��bt����!�}��,ٳ�T�lW��`�y./��	�
tn����]��x��}���,�vtbU}5d7�eA�|�+򶬉�|]WO�n�����Z�g�L��QG���y�6ݼ=�c�X�R���3��.)��`p���s�jlj��Z�e����X����]�
7�!��<;�١��C4:f��
��R.o(��w����g}�V0�<C�Y)>;_$|r�ny4����0i�Ѿ�1K���f1i[b��׻Bx���4��_
Z�+�7�ju˪/!@�����iG�O��ìkw���8e�W��jJ������)��2�lHrs6���h5�^n��\���s��95���>��`ҹd�J�K��/�T�,�/�(�ծ'���5k�u�s9W �ұ��؂Vf��%<_iG�+i�f��nid]ټ���ۼM�#���\�+���q�Ɩ���"嗥;�y��ABFme���7B����fH{%�yB��kׅwk�R�=t,N�u6��+�_tQOCI�NYׯ;�a��"�o���ǆ�	b���ۅ9���o����wod�u�vݞ�S4�
����WU�,��N�I^i��!̭��2]�4��v�uҝz��c��X:��w�?g*���yэ��̔��ŕ�ޟ����zwRݹG��[��O�̾�Բ�:�w:���[�����r-�}����SVT��z���<�:�#��:��	zD����l�b7�>�֭[{��Z㋳JeN���h)hF�qqw^����[g���f�]�-�X��������`�7��V;I`S�ٗ�QR�����:�}��=�Ɂۮ,��A��u@ܬ��m+9-�����ko)RVru�Գܩ�g a:9�����G0Py�
���<�\�,1��Sr����٤|��I��ܗ��E�㧒%<Ǧ͜˩�}{�M�g)�AT7�j�dM����ȗ	8��*�c)��K9��\v�%`)2:e���R��U"Ȯ��Q�/[�؆�m�䎾w}}��-�����s�')���.5�'O�d�c�]����y���z�
��7ɶpҵ��n]��N���b�b9�Y�K|�֭�G���n��"ƞ2Yq���F�/7b὇1T�͈��T�8��6�V�h��[��8/�y�f)u�V�˘�S*�N�;�̮$�܉����Y��ڼ\��9����U�}j���SDf�`ܩ��=��ڝ���$�r���������o��)Y�9��e,���5^I�mT��UCvEk��.���E�]��b�s�!X�d��4�lZj���M�ë��mI{w�o����-�R��CM�r�/�33W�Wgf��sU�#b,��r%v�3�Mz�oE�W<H��X���ג�=|�Gf��j{,]��%f�c��Ps�!
�d[�A�/Vݍb-]�����y����V���bNo4�m'wݼG9�����c��2,Ae*� ��G�HţR%Vv��r���/��xM��	Tup��ʲ��}�s�GAv`����S�R4�&���������3e1H�X��fl�#����3q� ��o3O���aDɽ7�i�6霬ntƷg]�׌������p��of.i�NuV��tP����[���%���"_d�N*t�]�]�iP�8�E�r[y�f��k�J	��L����&��M����Dmf��w�O��{�~ A��A��
QZ5�311��EZ�����TEB�U�3��mZT�*�lZ-[U�YU�՚ʥ`��U�k��ѥ�f�Xe��Q����#m�����j�Ը˖\���P�Ѳ���R�2%Z6�.�[h)Z0m���ՋTW,���e�����
e�nT�V"��I������1Z�l�m�E��J궕)J�յ�m��
*
\��u�:ӌ���Y�T�ʱ*TZ�e�-(�W�S[R�e�-iUD,Zb6Q�k�\U�u�5]�"%�%QDEETQ��)X�iU��cp\�8P��4���,EEX�u�aJ�nE�lL�K�YQf�)�L)mҕ�Z��n9�6�Qj�f�GJPR��% 	�(W���mf]/�]3�_����6x[\{�^ջ�Y6 !���}Q؝����X]��)N�u�u��/A�{9��q�x�,=��ԲNy�_�1Y�#�>	#>�i�9�W$�OX�e�� 7Rێ�''$J�JVJKHY��We4�mF8:�^c��	�16�]����RS)	���׹E-���c5E������M2��(�@hx���h��LƳ����F7	h΅�ߒ��P�Z��~�gj��ӌ��}R�]�rTڵ���\Q��=��jӜ���"�-0������T875�]	AJ�\�5q���$�)����6����6);������*����N�W��ImQ� �����̬�==�kvy�e4H���ܺFu?��[�4Po g*.B�vNL�8�\ywzw��/s}�K(���Y�.q��,��tU�x�ډ��9"����M�[J��Ē���/ �3Z"�%#Pp_��(��Mѳ��bVJ�Y�3��l��m��:�§X���t��?����w��Mă��N���+#��u��5�V��yef��E��'�8xiƻ��˾�r����D��8R�ޖ��Ώ�"���-Q��9ZҞ敦������z����q��_g%� 3����V��:��}�H�d&65�T�ɝ�����[�VM���9�D;��5q�;�a�\S�F�Nt�a�t�b�ܾ�x�t��驁x����ʇ�/��������d�.��H�V�Z�Un�_k[���־Wκ�l�����^z�M=����F��L��Ǖ��Xd��\����LCs�E�y�=m���ٖNq-�kEIȥ��=1s��)�+i��赀l�1yU���J^f�c��۰UyNU��E��̦'j�|5~ϙ1�fhS�}�H�-tө���3�����li/�ݫ�>�̵�x���W��X��dW��z�#H��m�
t��Ѱ�^˃��ܑ��n�Y��Kk��n��b��k8�:��Й�m���S��_X>;MշA��e��y�<��|�M��f���S�C,>=_g�$%��ʇ�Kk��Rm�^�:�䞭hv�s�>�n���*sԩD�nFũ0)M�*��u�*5�ʐ��l�������Q8�b���1b��9/���ׇ���w�RʍO1���*�6�@�]<nV�\�d!5�����G�ܒN�5k{��z�	d�ח4���g���&q��k)Et������n�D͐��K3��1дa��%E r�80�i3opj�j���Չ�k����/���΢�Z{HǗӦ��˻��q�]rS^���+�?!�,��>h�����.2�����먻�p�V����w$n�oU�QN��ؠT�����.��G�H���c�+	���}e����\�]�A���y0�N�;q�*����h	�i�T��d��6�ou�rN����uw��ƣ��]b��[����k��8�7���Z���4D��O����ڄ���n�ɳɥ1N��}cH2�K>��p/��K7�Ɖp�P}DFܷ7�W���8�*�'��,�o�n�;%���=HZ�(9n+ivҲ���ϛ�����������q��ޜn]嵥��#َbr�ޡj?�p��g�3�Ip�nێ�ӈ`:	����ؾ<{���q��#/��X�����5��%�!g����|�ޚTnL�}Y޼�en��`S���B��כ�{ɕ�;�^���!�1����E��$�^avT�[m�Uvy�]�i��BG�ŧZ����ڷd��)Y�Z<ͨ����Ml߁�fĿ��1:�)$&.��F�I�^�9��2{����%#႕f=˙�]u\%�:�O�J���0*�b�-6C�-!q��jek�J�q��_%[n��6_p:�W�h�,��2U��oj�43�ާ�҄,-)�Dc�95���7��>�YPE��"R�Sn\dS��P�S��g��Z�^̥a�M�jI�f�旡��lxPxp��66rҏ�3'OE���AU�Լ`��(��������E��~�^���3��j�-i�_͎>�Yv��]�ϥ[�c\w�!M���sv�S�����(�]�bڥ�Oa���|��^���ק4����z��]�z��JG)�%Æ��тS=�ڃ�'.!Â��|��.04)+Ld��.���}R��K����Ti��nP.���pa�{���ˀ)	V2���`�c2=3��ǌsY�9���G����{ʅ�DNT3��ޯ�ǩx�n�S��EՃ��L�ʺ���,�r���h���g������W�8ð� �Sr�w1E;b:lIՎ�n#���l�kH��رtE��*�=��Y��Tviգ
�ru0�� �Ɏdۚ����ϼ�7�⺵�?w:���江 �!��͟z��˪�f�z������Wcw��D�9ֲ�������݀!:�iu5X곽 ��2�T&&;/n����Y@T���*��g�yy��<<+jē�3:�W&�}�e��1"���}�����	|Z�Y�_^�]��rlDhI��pN/�7�wr�O�Uta�u��њ�ᚶ�d�>lXw��'Pbωۛ+XY�����}��9����v��� ��wo!jv_���+���P���-)��c&�*��q]�*���c�
v,�ÿVU��}ʃ̸�xw�6:o���8+��f���V���{9/L��y�{�fc��-�#���t���-��iש�a9i���\v�]7Fql�,�o+��׻k��f+0h��੭!���0y�Wċ���w�TI.�팭�d�q(��G���\�UF���1}�~Z��u�J0W��Z�yzj�w�:�U|OMZ�Md�:��DY��� �́�A��3(Q�'�8�FZV&�c�x�:�NT�kY�CնU:�2Bb�,��`룕Mˋ�@�|�:����c�q�͍��Szc��N���n��k\��ѳ�x�	�%Լv�5��.2EޡO�Ȼ+�x�fu� M{��+>���ZEj����t�eS��N�g��ړTD�-��笨db�����+����i\��f�r���2�u��~�,�Us΄^��S��[����Խ�G6F_���n"9��7/��J�zO:��S$��u���]z��yY��tU�i<0�6���ӳ��,ekn�nR3�;����v�++�c$i<�q�N��fC��g�(7�3�!o��Y7�����㏕���UVYP��ވ���Ñ+��08Ş z�N,ʿO�Q;9����&TN2:�����鄥�PP,JBQ���^q�5�X�O!�Cd7>8�����N���P�qG��q�oW�`��䍍���P<�']��9��a���)˺N!�Y࣯sз4���i^�F���5��g�8��=���_�e�����\\�v^o�����5�wE�yV�=��n��h���۶�uJ�=~A:{<�;W��`^j��
�M�c[�Y�<�~�Um=>�c8�Ϟ<�l�x+�땰p>;��!��"�<�N�"�vb�w�#s7�
d�XD�Ӳ�3K���O��R��w�~Cj^�ϥ�Ji�٢a��X�(��Kf�l���9�5�Κ.�`ٚ�A�y�#������ye+�+6Q3�RG����כ��k���n0B�w����ȯy�_ia�~[Q���#
��y|���"�<+i�\���pt�M�v�VYٛ�$�ݻ�E� _Ѵ�����K��M��{�{U���ky��Í�ƽ�C�uJR�W\y8��36���]�[m}�Ѫ}N���ݙ�V�74�a�J��l"�i�R�yI���Y���p�W�ĥ/�Mbt�M�P���Ⅾ�t���J�*������j�w��r{c
xN-�0����	��6�X�V���*� �*�3!��|��T�L�koVJ)ԇ�&��Z�%ߨ:�P`K��J&�nFl�<-acڻƺ���`u�ˁx}���Y�����k�v1
���$b�l/�����ʁ�\�qx��"���׬��N1l�;5��wNl��,ͩ�jw�ALG��ykG|��d�k���Ї0{rfo�q<��*K�n��]�g<q�"lWO��O��H⾯��/�x��'�Y��'�s[q0ŚJpA�b�Y0�N���L��b�N� "TMx��¸��2��Y�������2ٱW�61���p*cy1I�/}3��J����q܆�-ݽ�Ĺ� Vl�9�9\W�v�NW�q�j�堳yo�ÁA�sb�J���eY�y�7}ۭ�����=F׊�~^���걱�{z����`�ʋ�U&�T����V�z�$u�����'ANgb��R/�Y�F#���8�v�wC{�@q-�cm�Q��cmTfg|�>������^*6�-ޥT㉆A�x&q_n���83F�%�r��.�7�����:�,������g&�!�ns�+q�NWuK�60,��U[2�l8�q<Rk����z��D~ν�s�iZ�c�3�Ft�_��J}���Nߍs#�u*���|���(��8R�]2���W
�^L;Yщ���Lҝ��f�{0AEV��Y�a\��d�,~U�=��m���uр�$}�bӭ	���q���Ѡ��zgX��S~�&�z�y9���.�U (0�{&�����r���,b��ڍs9Ɣ�8�eoF.4RJw����8�`�
(�Z�(�8�ܗ8�@Y�K{�*�=2��).��Mt�L�au�S�S��j+��UTLhRjj�Q��.�|�ڋ�Q��k��t��W���%O[べ�{bc�lO�/�����M�/N4^Y;Ǹ����y�S�����᠌�	P`�������Ȭ��(!Q���cGˌFg��g����G��vu@�x4lf��1=�.���pa�{���2 ������y��E@�ݔ��;[F�n�
S��\���o3$���jUf������h^��`�;b���桱x0͙hL!����+����������ɝu)��=yS��\5?��ƞ�x��5��:_wg������c�r�-�����#)>��΅v>�{��s�� ��ͬ�B#Ɋ����j`Z��S�;���r�d��U��z*�H����7�l��nڊb|�H3.&�l*�rp�c͏g�ð�{����"��L�YO�#�Y��AY���>,�G����u�_��3�ӫFiW�B����{��`�ZI���-b�<�QQ`�/�q�Κ����r$���g�o�7U����h���n�Qw)�ܨ�]��W@���s����!�3`��V��6*v�,���h�]�p�.;J�c�RL��=�W�;��o����^�fH�S��D�9��I�R3�!u�P��X����1c*�q�C�T
O��`l��1��隍J	�M�W�B��'���\�~���}��1 x琠Ց�R~;I)�r�w�n�r��AO���ʘ��n��QQ(���*�R��z+�Qs�`�~0<s��֐�p�9�������4�q�.J$}�T���_ޮ
À�C�x�c�@�rjBb�1�QRE��Z8���=��s`�Ql�X���3���t�7���D���K�tu��d���J����	'L�k�����{�Q-��Ͷ�������'2��UG��r����Ǐ��՘u�UY;H�6j��pLJ��u^oS;��G��ur���D�0���M���=-��O%�H��+�5�^�\DZ��X9��l�:�W&5)�_��|Q��~ѥ�5�=��*m(�`�0�Q�V�1T����b�,��3]����T���}�t�C�l����5+�uvȃ��_M��z,�)�8�T/Z6aތy�~N�eC�sQؕ�	�O3M��<5vk{4VE��?�>^=B9�{�K��/]b����#��|~�kC���-�=�ˑ��`�7� �?ȑƾ?g�A�����G(5p�Qr�$T��]e�ܪ4�h�E*�Y3�,����Y���Ñ(eq��z��}2qfU�x��`w�t�r���O>֔AYLi��S�n��rм�y;�q�58/�|����A�6r8�g]�f�k��K��e^���^�`����;��<98�،kG ��W@��'����.�.uV�u�<e�dUc�`ު���yg�����]L#O�~`o��Ã�7M��Ք|ac_����Ox
5@�b�)��/pU�yɎ��!�� S�Ӟr,�\{�i���4,��b��Ƹ�d�y`��֐[F����ٜ;k7�n:5��@�g��L��՞���ya }��G-ۿ����4��g;�!�`�:q6�c�k�kx���1U�=�P�n�n�2�i+��7�QC0̵�j`�^�w�d.j�v�~
�Ƞ��s���� 6�J���rmU�h����v�;�e�սU��Nf���[l�G6�4���2f�TA����kv�����ӑ�ǟVL�t[�Ý�� �»�:YB���w���5�ܬFt�<nr(��V�eH����}z��Xo�6e^��O���{3��N��ۓ w����7��m��yY޼0������=;B�+�ڑ�Q�n�8�,i⪴b�#]�XBH��ӽ�m$��m���Gi(��=��f��us��ڎT�C��5zE��icU�L���W���(ǌug��t���Ö#a�lnw�z�T��r݇`�C���#R�2A�U�"�p���3j����Ϡ��P�6�oa���$��	���9�9�e]�A�S��O^�̞�٫<���M��*٫c��3aX{U\�m(.�f��5�����:�;t+#�������D����}xi&m��vi1y����t�F��]X�,�쥈ؙ�f��R�Ӱ*�%������T�1���:���5K&�;{\�%\V	Õ
�=q�>'�s3�.��ā���_g��jy�i�+Y!8)WF潡}�Z�y�����-�n��o�i=���0R�2�ɟRD�BmEÍ.
E��ۚj�Dc�ؔ���і����Z���O	�o�k�t\T�r�+�R�q�""�<;y��f��+�;�V>|Wgr�L��*�Ż�J/tj���-"+u�In��Ϸ;�h�1T��]��{HC�g8힄Ծ&��ɷ���N�06M�cWk	� x���0�.����]�X��hB�\����r�߲�5��!���vwQrڵr��Va�>r�����Xa\`�`�Ж�rm�W��v���6M�[�-����m�g!�[��1v	z���n��=�W��Y1i!��J7V�[P�ݶ{&1����gP'j�N�⡸ﲔG�E*��r�1YBT��z���(2wsgeE�z0��>�,�����.���U��L�c�ȫ��Q��}�����v.�v9��YZn��M�-�ⷧ�8�ЎM�UP��:^�\ľ��b<���m�YM^oF+�T�ql��8picə����<�UCHuen��]���k�}��I��j.m�|���*�:��������&ug���)�^f�%+�n���N7�:q�@�'#�WA���.J��
'p�mj�z˯�r�sA�H�dQ�EB�r��3�����ժ�Sv�utѡ��R���]ǵUÕ0��{b�O����]v���s8$$H[���6�s�ǁ��]q�ַJ=T��-=�o;C���ׯ��}�oS��WN}��"�ʻ��{g��t�wv���H��(/�V��-��Z��Z�k
	�2���ED�YX֋u��
���5���T�5XYm�JR��T�c��J)Q�kkX�R�U��"�ը��Y�U[�⥴��KQ�ť-b��m��,��JU���V�im-m[T��*R��U-�������5�5Zղ,e�[QR�J�������kR�R�T�����X��"�KJ�F�E�h�s�e��iDT�
Գ%�����UKF��jV�)D�KV6ԩVڔ�X��*�Qm�����T(���V1����5MZQIe,U���+V�+[m���(Z,��V�j��Ѵ�--PUKAB��j�[e�ĶJYIh�Akm�3-U�Z"ʈ��t�(��TTE���V�ZU[hڍ�"�R�j� ��F��F1��+Z�L�1-m�+TQڥ�m-����X�m-�*�p��Q+mG"�R�/��'rU�L��.�r0��.��� �,��gP�=����V�kХ��ko�Yo���ʗg�ȝ��{��.ǼX��ԕ������v�Y?9�B��g�2y�i���1��+�O;��� {<�f��eC�/�}��L:�Vu�3�:��Y�u?g��ʝT�곕�w"wwã� xC��sl��?!�~��a��"�;�@��a��d���ǈ�'�c:ɼ�Iɻ4��
Ͱ�y�oD|�Ss�a4���*;�I\qT�WQ���Y�<�����S�>q�����7�B��L5a�u4�Y���>O��E'������i>O{�����u�)�@�*>��3|�bM�Sa�;�'��G�0<!�Vvd?�������Xz��rO]���C��i���qC�d���N���掠T��ܧwa�k��a�纇ڤ�8���sXi�$�ĚJ�{�1>d�����H?�4j��q��O�@F[�>Ik��}��k;=�;���I^��H��yi1���c'�߲k�8��Xu����R��ڲb�q�{���'��'=s������_SL�,����"�����o��{���~�_�)G���:e'�ʇ�۳v�uP��M$c7�gTXy�i6�0������2���E>�Xb��{�4��Ɉ����%|\ *n�Q1�~;w�y�<R�`t �q�Y�AaXq�f!�UR8ɩ�`
�N!S�ydRi�q��̆�HV���a�u1 ��0�b!Qg���i<a���S|��,��?c���;y�;ݺZ��ǶG�@ԯ{�C�6�ud�<=��a�3�Kf�q
����E��>aSf�Ǭ�q1� (��/iS�&��~֤���B���a��I��bz~W-�MP�2�U]t}�����h�G�	�x���Ѥ��d���wO�T��~���ua�<��u6��ViXqƲTR
zp���8�!�Re��N�É�4�R�3~�S�� D���0��{��Γ�_$���H�g�����'����a^�{�km ����|k����S�<;��=VT1�9��HV�W|�é���u9E3�
�J�K1�P: q���~�C��7�t��~�W�ÇG8{��]���KgȂ!�|�c�H��A39��ܐv����:�i>F��{[�D����YP��7K8�#�+����D�9&�7�J�Ե���&nl.3��B�y���P�x��<�]��5���!�(�t�A�g���ʕ{�'�� zh�91˞�P<"g�G�@�o2~aP1*��&�������*(|��x���y�b�d�>���p��
��Z��m ��7��H
�LB�w�:���3N3Ϩ��R�?�
�~�ھ�>]����@1�Q��;�c6É�q
�������N����'�}�E�'b�'�i:�g��b{�%E��T��<��CĘ�d����(�z���f8������[z�_gƄ������l}�8E�;�i>@�6�?QՓ�_�
�5Cl9�O���{7d�z��=���ALd�~w^0^!R�﬛M��l1}��h%gU��rW���Ϯ����Ke����<����������߰yg�Mj�ϱ�T�d����J��֕�����g�i=d띰�va�
�d��a���Y+������QH)����bN+*M��>]N���ϲ����0������qͳ�&$�M3�4�TP�9�	��?0��|;̞$l1TY��T��J��d�ʊ$��0�6��+:ɹ���V�Vk�z��'S}���P���}�#�xD{c�HiUI�t��OP*O�s�7�B��y�3����1'�g�?&!�+���H)�f&�(��i �CybŚN0�M���u
�9g��2�J����~���.�"<xL�}�����<�Yr�'a�=>�@�+�J�d�&�^�ua�m=@�>���d����SL<a�)4�&=��g�1�6�TR
x���޽|P�4���gL��� ���~�a���|�@�V|�{�M<d��l�2)�RW�8���z ��2wT����@�+�!���J��u�
|����}��m>dӜ��s�Z���$d���y�i�������<&*<;<��6�Y�Lk'좐_2���'��a/ԅa��C�L`~?s4��1�aQOC���:���~�(m �a����,�
������7�o2�酛)���L(�·5��(z���g�9��'���Q��B���w�,?#�Ag�5�iUI�P����^�Ì/)
���3���i�zO���=a��G��ޯ���b2T�S}�7^W�th��wQ��[H��y=���;��QT]({/۞ �����;iv���O�m!W�|P�����<kwo2�\bM�(g$�adb|��ua7��m��vw����)3��E�ڣw��q|\+�#�5�
�5��?{�xR��-��my��AO�<O��q1H=����m�<N���:�I���[4�XV氿P1'�ެ��N8��7��ҽd޵��2T����'Si� Lyݺ)���v����~���e�'|��zÙI�m�n�:��?[P�?'}�C���VM��5���5��J��S�*�1��Xk,1:�J�ٴ��>g����/�b̮����l�˻��\x�|�!5��̟�� ~I���������~gܡ��$�>��2x�o�>I*��}E'�&UY=a��|��s�3{{Wq�Ηw��>����@1�}� ���M����6�|�����,�
���1�+��&p��!�8��:s�J��+:Ϧ����
��{��x��9H/���Y+Tu���y���ϴ�]���ߵ��CI�
�:o"釬/��t³��8Φ'���É�jy�	���a��M!����{����Y��Oܤ��:�f�S��r$f�T�I�/�9�|{�_;�y��\R��xnȈ��*=�f���<J釓(��2T>�5��bq�Ն��vOYyCٺM0�;����:�H,�M�ϵ�OP�<?|�v�z�C���k(Laϩ�����s��켕�Q��=}�=�!��ʟ~$����fH����!��eCivi���;��
�������J�CVLN�z�q&�i'�T��g�����4¾{�I�)�Ag��go�ܹMh��ʗoѧ�kK���Q�}ʽp* qS��C�.�
��;�������xw�3�~C�<>�I4�a��¡�1 �͟Qa�Y���g�P�%z�a�m ��J���3y�}?2	P�6��4ws��� `{�	�}��I�sV~��m����f����w�d8��H{M����Y?s�6��|��L���sĂ�Xbbl��LH)�k�,��P�N��^pP��9�(��%c����=�G��(�I��<�i��>ޡ��h���>�
A�N���p=a��ONw!�Y�%I�߰4����'��6��?e�l��y@�fP�<��[��~=^�t��]rTyU�Z�п�R����:���+�Y.����M"x�m2����s�D0'nt�S\�����RM���w{�Cjw]w�;{����Eġ��I��=�F�0R�+Ebd,�WR.·��ܻ�P��Mt��{����ȕ��8�"��Ag�(�I���530��/�*y�{@�c߻�b�P7<��m�T��%OsZ �QI^���d� �γþ`}��ý�F�x�(����ݱ�C�����̍h��q�&8�N��i>B������+�z~�k&�M$٫��N�;�P��&'�I�~fM!ԗ�Cɘ�8�Vq����4ͳ�c:��񺻯������U ���yz�2�9��{��o����ă��\�:��Y��g���q6��+��=�� (�P�馻@Ğ�]�Qd޻�*���i�a�r��P�|�P[�R|�O�6wXg_q��{��k-������{��k��?3��<N���Ag�>O!������;��3�8�0�sY}d�Y��<�p��Rb������fQa��h��&�4�yE��]0��@į{�|�뭟o{{�|JS��sW���"<�ޘ�P"{�'t�2i'�w,�Os�m!Xm�2���%M�|���I�TY>�dS�O\`�C�f�A�������4�Ĭ6j�1��%z�u�������{�3�}��<����6@���x} bA�7<�I�,8¤���4��٤���@QN�|���q
�K���B�����6����i�d����)�h
~@��{s�}�������o��y��ת��1%���՚a�Y��S��,�:�3;a����d6�����a�l:�f�W\�|�C��o�wRx���ɾwo�1'��ϙ<�a
����t��=�Y���;V�~H�Js�xlyǅ���>���%dUU'�*|��ְ��q�^SH�L����w'Si�0��H|�E!�{��x��1�P�o�L咱f�O7�>J���~���_�Z\#+������-�:=�>�@ D|>8a��TC�~èbA�(h勦aP1�d����<��/�N�'{��J��dמ��)
��s	�u1 ���2���O�����{�ݮݍ����|���`\{�*<"�a�����k����x�Ԭ���6�g���a���R
TP�9M5�Pă�G(�{�0�oT6�H{l�*
�u���i�
�HT�k����ж����o�\�ۮ�X*UJ�<��+�y����*Qhu)P�3���@�E���|�N���K��5
sdO�W	,[�,�<�/���<�QJ�9�|mm�b�z(�
̰����
9�+��଼�F��������"�Q(��,��<<=�[��8�|��$���!P���¼d���'��2i��]�w)��u�
q����Cė��s!���a�4�Af��3ә�AJ��,4���1&�����xT�8T��]��2j�p����J���y��L@QC[����Ǩ�����g=��Nk�f�u��{�i��Xk��ҪO��K̚I�x�0�ڸB��!���?x�G�������}��e���w��g���b�!�TP;�����>O����풱f�����R>���1~��f�m�N���ݰ���h��!ְ��A�s�����ͤ��mE�ɉ����5��S�#_ƺQH�*�@��S����HVO�r��|���k2~I�Ğ%E��bx��o��!R���<a��b�_�~�6��*J�<��Ch��)���m��c�E��;��z$��@�wYݥ��>���φG����I�m!��;��M�(�a��'�?e+'�ܐ��?0����SL=���~d��<�R
x��l�8��u%��O��6ê�gY����������sk���2@���v���TR���gx���C�s�a��"�;�@��a�]5<d�״Rc����S�4βy��=7f�~aY�Osz ��J��o�w[T����򗺒?lDD8`dx���M��|���7�B��L�w��:�H,�{��6��TRw�16��bO��� �d�]��a�R��(Vk�LI�Qa�*w�O<���"��w_|��9�}�<�	��#������T<9���2TY�=?fM (�d�y?w�@�=C�O{�C��i
���>�'�����4ϒ|�M%Gý�'̘�6Z/�T����4u�����D��s�'N-b \xR�
���M��gʒ��2M"�S�ߙ���C<=�&����ՇP�s3H%Hr��jɈ
)�|{���'��'=s���!�
�ɮSL�sI�ח1�n���w�����rOY�%q��:��SԚ2���eC���a�B�^s!��Af3g���8¢�ߟf�l�O�����^�u�"�}�Xi�P�<?w&�&2b�����~����*����k���ӺM�����������Hw�q��u�&�^n�ўG]�.���u�;��7d���#Ρon��pVhK�;���Ū�;�T�1��w��9���`N.`�i�[���ʙtH��������&>�NMW��9�OM�s����|>  &�s$�.s�Ltl *�t�G�2k9��������UR8ɮk URq
�5�I��3��B��~�}��u�LH/��a��>B�ύ�$�x��1��}>�k��מy�������y�� �d��=�3��1�_ya�g��b{�"�l*g,<�i'�6�d���T��"�����&�a��&�;�N T��0J���z\�	�U�?
꿲��~3ݥ/�c~��z�������8�O�o�4�S�'|�p4��H<����x�0�V���a���Y�a�.��QH)����a�1�-�2wV��\ &���a%�:ŝ�J�.��d�
)�y�q��a�߲�����;@���l:½d����.Y�J�3�n�AO���Ğ�*��9��HV�Wg(��i �yȈ��<&@������V�|�L����5�����|����=gCwi�~a��������p�~N2c#����J����y�b�d�>��w ����<5��F�:�s���T����h��x�8���������s��^y�o�;}�^�{HV�tSL=g���1�a��?!Q|X����5���6�ud����Y�q� m���N�Y�l����J�0���y��<I�VNv��Oa���޺����w��f�d��G�
�1��L�|�+�H
.!���i>@�6�>��'���+�j��wt�����vLg�?8��i���Ow�u�� ������{a�zw���Y�e����^˹�]�����#G���������������&�a��T%d��c�u��)��²z�q�z��4��u��zn�L=a_̛���G���+������vf���}7{�o��RO�B�Dz`���2!XqY�;��:��Ă�/�6ϐ�=aQC���i6��14��;̞$l1TY��T����N�c��Cԕ��Mٴ��Y�O?�ϫ8<�{�fZ�J����1�1���8��ϙ�}��T�M����'�����08�|�*��:�a�?&$�}�<a�1!]��4�S��N"�C�+,��d�~��_A#�:ه{��BV7�tV�~�;�2@KR�e�TKї;��=sط=��?>P�2�̕{�w�7�����#�X�Z��0�&Y����\�7�ge����;/1���u�\���eK��YFdR�"ۮ�y�Gx�6I<�Mv��ۤ�߇�<=�V�t�|k��p.���Y?���(��
�7ߴ�|�a���N8��{>�@�+�J����:ɴ��Xq6��T��w�<�|��yM0���|��l���g5�^��u�dS�����|�২��b��
���������t�&�6��}�����ɻb�E%x��=�������g;��6��VՇ5gY*s0S�'�@� I��}��{�ޢ����d�T���!�q�Nygg9�m�Wo�<��>a�SMd��R_P0I�eA�%���8���q�ɌO��3�ugXTS����:�����P�<#g���j5�������ť���G� x��{�u%}N2c9��$�>����x��Vc�G_a
��ި�����oY&�T��O�*Lg���a���|������p* 2NΧi�y����-g��1���=gC��E ��|����&!��w�bͧXc���M��
�v��̛@QaXh氿P1'��Փ=���}ἆ�6��&浂�2L "F�#��GԳ~�;��?{`\ 
���<C��q�t�y����r�������I�9��QH)�n�!���+&�ܚ����an�:���URc�%E������Ï�;{�pusG�յ��ƹ��),�����aP<J��}�:�Xl��E:�󉤞g0�>B�̝sw}�4����Nw��� ����kv��Q`ny��q�1YS���G���`ICs�h�/7�Fwq�?DD�>Ld��Vz�3�
�i1�a�����,Xb,�
����!�%z�d�~��(q%|t�k�%I��f�w�=������l��0"�xD43L��{�<��Z�%�󧬕UC��P���Rf�싦��X��
�Ɍ:�&'�tea��4y�H���ܚC��1!��rJŚN0����1'n�vs���f��V�'/��K��,������=�]��CQ��=v{g���]��ٚ}�����U�K�CC�Љ5��g��҃t	�,njG���g�e�����{�����3��i�RR�2���n�`zw�v��9��R��Yf�Ʃ]��TX�J2R=liJ��Mlt U�H8�*���"�LY��ӑE�W��;�o�Y�eV�Qͺ���xݶ���kh��Kz�+�ݱ�S�ph�a�<[Cֺ�tnv�fV4"`8I��J�Q�\1�x�3�ݨ��о���gMg�Ǫy� ��q`ٳ�f�ìU��η�#��|��[ݪ��2%�����������,��Z��=���v���^!���D��X�YJ��*����5�ߎ��$�t��z��ڋ�iV����l9a x���!����_�(}�}NN���a�x8�<;�v�)M��P�Ck'v�|Wo>�cu��G&39��� ���'㤞�n7<��� i?V������ז�m��Z�8:5�f)o���Vk��ǎpT֑ӇF/u�ʷY���s�RG��(��)�1bx��4�)!Us�≌}�'\��ZМ�j���/o)�΢X6�IQ1jB�	��5�Vˈ�S~�b�m�@>r�Y�4̈́(ɘ�g��.�F.8N-
D(~#DZT'F�3Vي�j���b�(jf	�gj��q�#z�}mFL�mUn����j˰�e\�{����`t��C�q����s��k�����xv���k-wd4�pұbܾ�t0��/��GwDdW�ͽ�7�D�\�o�����c���D���[u���)u6־�z1�^��r�WL��p=��.9y�7xh�774Vq�������!Ǟ�z2���S,B]v-��R�EY�S�i�r*2ѳ�x�w�*�'�^�>����bA��9��ۄe��^Ӕ��3T".��[�aI��7�ܼt�e?Dcŏ{p�i{�̲q{�u`5}�c����X?g�O�:�[�T|���9���|�*ӧg��P0�(k�6%�S����]z|Cϐ\-��WƅW��Wl��f޺l�^о�aVc�u��L[��(Z��9v�q�58/���^}��-s��}��5��ͼ��m^��iy�s|��s���c|�����):��#��͵pŎn�u+�¦T�WX�-
�{\ڐGu\7%�t�b��/�[&M�G'y�U�ЉH��̾ج��>��9�5^PR�.U�{�N}�y���
w�Ҙ��n�ӳ�����<�Z��즋����#��x�b��t�~[�]W�[�N�q��Ɩu�IIo�w�[�a�[v�zY�z=s
�s4�v�z/dxgv_�,��=��-��^}��o=�Kө�����]>7]�*�EM���x�e9׻��t�P&yf��Ӗ��0������=維��4���*�Wk-M���7j����٥��7�� R)c�W�#XV��rN{AP=Q�,Wxsb���ʿ��w^�nq�kH��*�ѹ����m�9��:o`p�t��;�b�c�R���1R�.[���Z��k�P�1��p���x9�r���aL\ݙ ˣ^�@f�4#+�ݗ=V���"7�=�tp���JO�s�k��k!Fb���P��]/e\%�Yݰ��)%9
���q(O�g�!�τ|���N"
�9lV3��
�����k�&�)��ov�+cnd5�ъo�~�ׯ⴦;�;�v�~L>|T����.��QQ�kӣٺf�R^�e��y��ĸ��e�W�B��/�����^#�cǌ2gzk���Z;�)^dd?iՉ����e��9�]�T�N�(g�DzW��ة��kr����6�z�gV��O�㚸�����v��!E�3�9��h����H���a~��"�Ι���v��"<6�[��ҋ߼��gVu#�[w��P�#�y0�����a5�ˇ��^��^c�+�h{�59a�V���lb��6�\�a��y1��	ڹ�*����]����	42΅_uEzKK��n_m�ِ��m�a��X���T��F�R���(�}��hVI�p�d[��il6�	�n�T�jX�[�{�2D�����OC5���_�04C�}���ph��.��s]��I�Ԋגn�S�[��c/�˴;��	�b�,3���fe�/vْ�n�r��K��t��rE�b�dk
����N$��r�	Ϩ�\
v<��g�G��
�E-d��V��t��>d�;.J��w�˸�Y���׍*�oQ���̙Z��K_=;;b��/��j�kg	���g�Q���Oo��(��*�|�<��*�O@�9�z�a�7�t��X��)�V���nV�aЗE5��(s����u:�0�+)�}a�h��fX�`�;-���:�x�Q��x�زa(�gmJ��~�*��t���-fh��@i�z�΢�{)�e�AX���D�^+�"�)�F8����&j�7|T��ge!�vC4c�fڔ8�w}hԤ�p�އqXl�����w��U����Y�Y��͛��(�)��b��x�`�� 8���.��]�7y>�Wh����љ�@��f�<�Z޺��v�W����W�$y��x���g�#P�a�\�i�ś�����7�(Ȱ�s�Y�
�ּ0{��ټ���I��;�X����/�.�[���r�6��@��#97ԛZU3���Nʇ�ҷ�ו��]�`pj�J�ݷ�.�3�a�ɭ�v��|߬o5���x�H*���]�oty%�+�k�J���fc��ͭ��V�q��/eoeK��'{l���5s���J̺���Uކvi���{*��<� ���]�uF�#~i�>����6���&#�D��7˙�᪈�tr�Ck����;ʎS��['再�L�'G�KU:�z΂����U���Ы��Qs�ʙ�6[9�B4e
�)1��qݩ�:T��2E��{���c�9��,�m2�ۊ[�w��l��]���_4�,N�Ὰ��+����w����aW�;ޮ�,9�$'"�����|3��)`t����'��K��[��,��;0�F��F��h�Y�W3�b����gk��1)]�;��i�a\O��U�\��ӵ���o�}����(r�����xnQ�":=�s�����W�B�o)�2�- U�u�ԫ���N,�4C�^��^����Ed4j
�z�h�rՕ�iD�1V3�W�`��J �B�&W4GF�.X��/s%�*�M��wSv�ޣS(sӸ;\Y�os6�i�/[y���P���c5�{,��5�Y�k0�:���U���\�{�t&�n�Cz�g�V�+G7��J�ʜyPe�ɶ�c�e�]p.�j�K�&:�)XN���>�[ٲ���<^�qR�#�VB��y�z��q���Oٕ������ݿf��!�,aH�H*�kD�����%��DmYJ5m��QlV�h-Zյ�����P�R��F(�X֨�[Z!Z�r��i���Kmڥ�D�eD�Q�QR��Y��nZd��Z�إ[Ҵ���Q�*�Q*�Q���5��EX�TE��Z���-T��J�V�F��R�ƋEeR���QmE[l��+*%+AiU�j��f*̥m*(�*�Z��*�ĩQ��T֊�i�m��F4����s(�JR�Q��B�[eF�̹-�Qh��k*(�8����*��mYQ(�f�X̡DX%�@DDD�Xj�-j,Z1�`�m�JP�kmP�*#e@��X�ҶV�����6�r�*	m1kee�
#*5�"��R-J�KF���kZ�J�cSM1.!���[jZTE�P��m��T�#--kKJUF#UQU(�V��TƷ-b�l�X�DX�F���DQU�ҥK-�lu�L��h���������>���4b��ㇺv𿹪�x�9�`a��Bv�vu`�t	��t;w���L�����̊³;"�1t�*�����x �wy�����b-� �f��+�cC�'��1�L�������D��U�(�)ɹ�0o4��v��)A�`0���������L!�0/�\c�~^�����C��o��ţ�BE�uV��R�(�/[�bnٟu����=�-G��0,�4,ε��V����3t�)-��+qрj�0�WkZ���v��q�p:��~B�]F��<9h��=/_bV�6X���U^��*�`ڻaI�
��;��k:12�_?v�3��^s��Z��B�J������x�d[^��3�i��)K:lZu�7{<�[�;5rD�A�I�w]L�QH;�f�k6�o�fc����p=Ew,μ�F���P�2�Ћ�;��0����o`P�;��]P؞�7�����Ϙ����{�� ^<x��d�v�����".��h\��f����w�OTߢ�A���F_�� D�����p�S_)�R��VU���k��c��U�`np=:̈́p{�ԟ��XoK'�Ɯ��6�BS�<�F�"!�L�1��*��]*:L��w)[�c��:i���=��Azm�Jveo"Jū�f�ovN<�y%o-Nۥ��^9:�\�2D밐���N��.wp���B�YXdۗ���2u5�LD�����0�2C���8z�� ��=Z0Ҿ'_L�9�ؽ�J.4L�(�4��J���;0sɞ��н��T	[՜��6���6�b�.	��/4|��%|�C�������WYÞ�~��*��2P�Χ��]ν�U'����|�H��&O-���y^�C�8�����J���N'J����<��7z*ZuqF|�!���>se���>LV�v՟���9Ƥa�0Ǎ���IAC!驹E��z;�����W���h�a��G�sWū�q}�U��yƍf��(���`��r0��[v�����9��:jzg���!D�|^Ļ
a�јZ�K��9�O����l�^3s%p[���љ�YXk��Nh��ZCIb�2T�o1U>��'����6*v�6Vc�^��9~=א�'`ųAl�;4(K�J4�ե��-��qlofP��*�T�9
&6�D7&,e]�9Hb4�[�Բ?R3�8P�˟D���~���r�L�Iϫ�����'��;)?$�_p�H���?�����
�߷W��y����M��=#��\��z.���In��#D]n���S%Q�Vj���cs�+%�1Ӣ��k���*ȳozQ��
w�Z���_m�=��z�Yӄ���5I�-��IM �H�ofU����۝�v�5��8���xD��W��x�ڮ�:���3�7�y�a9�v���i}c�_����x�Mi
�Su��;�ͩ��)�纅�>���]3���,b�'�=aΙ�:��	8�=�׫�'\�v��y�b-3T�ku\��mg���M(ϫ��>�c����r��E)>�b��6�`g��vB�4�Y��tF�E�YU���H��`P��~�EZV&��3V�1Yj���LW_���C���i����J��99R���{~Xv|߁� �P>&�S�qȨ6��w���&�aL��I���l~�h�w!��#,��r��ן]WA��*�u}7M�̅F�MgKr�i徽;J�m򅵥.G0���և��t�|{�'�>d�,��]>��umF`��.���	�n�T��K�aU�~�E�[n���)��.�DV��)T9Hm�����׏�+���.y`��af
͞5��vy���]�8��J>�'`�=�����~�u�x���ʽ���������tl�{����S�����B"��n��\-��iz��[�cܞ�`|�AAOV���>��K3bOR{y�#�;��j�`��}U�C��2��2��L�T��D��j��w]�=+\<u�;!���{ɂ��8�t�n��V��@�9�
�Vw(��͋H?W�x <�L7�W�nL*�E|��S5���d�W�5ͩ��p��f��q1َ��:^ƺ㸫�ӷ����k�@����%>�.��`^2hy�Y�����K���ncrc�ܡt�gD��F�]�M��^{C�u���gj�<�lLU���C�8�ꎗ]]��\�]�m{�1�^ �-̉R�ЯI� ��T�,�R�0�}�U��,��T����a=S�o�ʾ K�('&-��]���w��2��9Z��DZt,:ӝ[�飮���IA�-��^�ܫo�z��Z���r����F�ۀ��'��5μSƁW��X��dMf��죗~����(ԩ�l~�Z���1�u�c�4���'O��@Q��+�Ƴ��q��ry�r!:Or�嬙�K���*�@�B+ؕ��J{Z�s��\��{iz�<}ē�_�=ܫ�������Ν�K�bW�,
�PnE9�J�M��(msN޿w'��E��u׷�xM���f��\j��گ���u��9�[B\~^8�J���q���7n��)[�9,ӌ�X6/N�An*��ghJƑ�]:L�*��;��˧{�##j����V�̭/���i�u4Q��*+0Of��{r�v�n�jp��ڔ�#�ڙx�N�z��%���ں�gC���\q/�� �oiw%�-tdW�(q���NnSqNF�i��X9�mN�W8]�>� ����>����d�,<�nDR�� ���1\��N�=u�$(�f���A`�+��r37�r+��|:{�K����B�/��<�� :�.(�oޜ�-`�$�v�0U!�G%<�+*q*SE���Rΰ&Z�*s�J��C�(����i�=����J�6xߒ��u��~�we�%4o,QX������-��f������C�&�g�s�<���φ�mu��2J,��(��r�\�RE-�=W9p�P}DF�盬�b.pFJ���-]lsEm�>9��|٥���v���8�׃�����Cݳ>�5�9�_M^y�6+�:8G9R,���C��{�e��%�	�,]�+ݵm|M��k"̔h�kq�Ft�[�2�#-5u烨��ݕ
�;�n��O����R�5^��Zvc ڻAI��!��yߛ�{	񾂷u�粫y�J̝��S���KA��b}�<E mKs��\,4�^Hb�I�j�=ƕ$p�[aSQ�ۮ�>c���]7��;kͯj^�US͘���N�P��{�yvit�͓q]u�F�`�pӆ��ֹ�0�+�$��^�t}]����|c�m2/T�
P��m^��̀.����9O
l����l^;�C�OzѹU�w7*�>����{��Bַ��ْn>�g�@-Y�[�mD�`ߪ���'h!!��~ɤ�9V9pvPd��c�p�w^)�Z�,��0�x,wj5ϒU�M*�1���6�=*�}�[Yα5.w�,���q�.q�aPlk�2 ݌s�ӽ�zߢ��2��	Ф��2��ܵ�g�茙
=Kka��׊.�gҭ�a)�OG��ba�w4��q0�
�͘�i��-�i7��\�bU~��^�4I�Ƶb|;�'��S=����=�Ge��5�LIh�jkx������g�'ˍ���������+���]X80�������fU߽��C~�X�^ 1�qO�����ܨDy0+�Z��^�D�a�1}��Ui��]n��_,�rㄻ�{��z�!G��=b3��}ݰ�&��˔V.Iv�y�aFu7=�;Ԍ���p�>4
���0�<f�]�.��<���bXuP[<��P�(��<V��ǳN��^9��`�h����/yKO���O��OI�VTP�x"��]̷�l��{5��4w%������d<4��~lv������V9K���S�-��Dl��]��	\z�F!�.���NJ��o��m�V���:Љ��*˅��-Z\�Hl���{]�9���"R}V�V]K�{� xG+G�����`Tlw}w��c��e丼�Bs�W@	*�Y�U�]�`�*ݍ����5-�y�
K�P_6�x��[x���V��.&��sǺ��`�t�r�4"F96�T��S�5O�x���-)��c ��%^C�5qC�-3�NN���>u~AT�
�qc[���Yp?n=��:o��$�zas������������g�0�Y�9]�^�{S��|��Z����+@n�o��Xu�Cj�(��|X��f�ǎpJ�S]eP���M��Nu@~�6ѵ��)|�D�ǜi�R@UF�oL_���	"���+ZNz�'9���)�����j&1HQfBr���+e�E��b�m^@WL����_FI{�N\A��2l�9E/P��XC������о�4����&)B�-L���R������g���s��(�S]N2�g�t	>Xu/݂A<�|�.l�Uz��3BvͿi$��'�ٸ_���Sܗ�N@'�q�L�]Ҙ\x������Ľ�%�d��{,/h����v��䳃۔�������ߚ8�-x�+c�*?�V��Y�iO��Y65�M=-�v�O�}S���s�jr�"�����S�F݃�9g�����\��[�[��{v����gK�P):�����L*���xx6��v_iU[?b�*��G��}�����!9��|��8���t�3�X�*�eǜo��*�-̋b%#��r��*t���uX"�7~�AT9@!����\�:��%_e�}�:5��S���N����g4g�w���8}�N�s�q�5�u�֗)G�5\s���#=
��jjJ6}�����ʯ6z׹W�nf�u�o+� E�N���w_2��t��dF5<<Ĝ��:^����W�5ͩwU�s���ba��9��6[�U'��,���(�UN"V�����S�hy��TE��R�.U�{�I��j: Ŭw���s9��{R]$F?i��Oz{y	��e����>/��G��s����$�t�pќ[��j��{@�1�hC�r)��c�ݬޖD��\§3K�a>S2��>��;�����a�q����/Ng�ѥ4�v�n1Έ��[�9�7��t��~0#r��_�J�+����>��(���ϲ�Y�Wn�:k��<q�u�=��Lyg�J��Ƅ󜱘箚z����4j�y�b�]��̺�A����rÈA� Aup�;1<d��7��Kf�H<����gݼ��Ÿnmҧ�K��8��y�Z�x��ސ����]�GY	�}\em��\����WP��K;i��	�e�n\g��b��
�Zvƒ�� �<�Ʋ����b��zzg� ��þ[B8x������z�����9����*#�:��������˚��}�v.��:m�oJ���}`�쏁��M�Pjԛ��&.Y�ґ�;����z�>=C=9!/�Mr���z�Ҙ^�����Nj�(������Tig93{�f�H~8���U�.�<
,����[�b�qW�21i���8p�Ou�o2�mk�T��w�%C�
L8�8���BS���r�� "9�mN�W�y����j%�V�*;{���,T��<���c��}*/LW9z�]p�
.Y���5]d=��)YΨ-Z���9�����N+ېO�\Qb[��z�ܲa��Ź�=�)���ƦJ�����P���Jj�/����jr�6�{�8+`�R�l�&��'i��s����u��ɑ{���ǐ�n���Lh|d�)���}v�Z�Cx�9R6d�Ʌ��ze]�,�yl�p)�s��uVy�E���QF��ߗ���H��j�)kbxf=�J�E�^���>��힛�=�1).Ն�N+�j�b{�{P�	���7N���#9D��ә���}�\5���Y���'�������'�w4&Y�;+_h���G&����L��6��'N���U��ۍ5E{�����+$�'���zz�2Z:�To�`��ob�^wXbx��c�ddu����j�5�f��[����9��$�3ʀCՂ����\7mGF{N1��@$;oc���c.2㩾�@���ڔU�cL��7z���
c�|�+^3�I�/��M5n�'�W��`<�����{3D��y��8Ypn�=eD��9�zf���f��z��׼�k��Z~"��=ۊ�cv5��;٭䏻�u彽g�k�<kx{gC���_C����Dgp�a��FlF�1� <��IX`9���,b��	�(�.ddN��(=:`c� K����۞�<t�Ң\�p��w$Z����3 盱�qӽ�zߡLP��|te��\p�\6A�棪�(��J?<vb߱��*��������Y�0ܻ�X�Q�ظ��B�Ŗ8��V����e�k.ś�j20L�(�!��Q��m��)���Fz�0u�(�wy�9~��Ro� `���P4|���x���AT��zb���(�� %��F,�"w0b�ǟ� �7�fP����E	N��Ɉ��*�cwz/B�|FA[��L�A<��ko��$��bΚ�WЗ0��7vwK�K��qFn���W8�wv�<V+f�倔�j�y�u�K��*��ކ9>�<�oq�nr��0���-�tU�q�a���*R�Z��I�v^�y�&��k�YP�l8�Il\T�ɲ�oN��u�[R>�c��c��;���*����SP�w�\)�;�ݮ�o�T]m+B�S��s��Q�>�I�:�J7��8䇩�(���p���͉M��$�N����<-�{L;�C&m,6�N���m��'k�@)K�n1˻	�%�6�r��9���O�U'|h�}̌��W�d�k�d8\@��u��1�tܟTD��L7e�3b�7��cW�r��a��|�#�s�kν��,t�U�l[�x';�T�=�+|z�a^�}��Q�X՜wl]l���VfuJ�EC�T�=y*�1��s(I{gQ���q��U_'�.t+��H:Ng˺	��d�9�K}�}�V��6�趣y�˻D.�1vp��{�w�J�����F��W��'<��C2��l=��bJ�LS/��K�U�s�P�r�j��� �o~h����g]��A�u�L�EqVb���h�Β
@g:����)�L+�]��B�WK��Ξ�O/Z9t5s�
��;�;�nQ�x�0�U�\+w01���Е;���6�Uwy�I��iM�w����p��砵�.����8��1�����Q��z�����0w@�ڦ����=T;xK��l�C$��5�Zc���4l���r��X�b���*�X;�����bu���)��]�T��9Y�G��Hlw> �M�SihE��m*�WS�����P^���F��t�A�
���ks���Y�u.�K�(���d�.;yҜ��ŐS�z�-k>��[����;s�����'\���_H����+3ᯩ�T~����<�wɆ<��OzL��ë�£Y��=k3�F�(ޖx���[[�j�ƀ� -������p9� �@g��W@it���g++�Gݗ��{/Ec��J
j����Ʋ�{p3WQ�N�G�����L�w7q��n��
��Uѽ��47v8��=����w|WY�� ;�lCcU�p���|�D\d�b�t�̾�F���U��7�۫�"0��\����*�76��K�3vb1�o�,�G�U�%�e,����k�PN�M��2�Bܗ8F�����u���-��[���������L[��Κ��~��x�U�Jg�*Œ��4�-��pP����o$#�n�X^�h���Î�G0�w{��wMw�_+�Ga;g��ie�Gs��|��k�w��{Ǻ�Mݘ���zt{]SZw}p\�Oq�kw��4��i�4E�ŤJ�ë���~�eKiD6�kX؍E�,��QՕ�j*֪��ڪة�J��iEZ%�KU�Re��e��1��:e��q��8P��MT�A�F�`�k\�̷YE����mKEcir��EJ�J[mkR�"Tl�kTQD��KmiEZҶ�U��J̴m�r�E��TX�E�Q6KkmA�X%ՙ�ij�.[5J�E��n��3���
Q�F��ҥ�Q�KE�V�%X+Tjն*V�*����ز��m�e14�,��Z�ETX���Q�DF�"�)F�FZV�Ҍ��Z��+QQ���ոɃVcieZbB�[l���Vĸ٦�V"UUTWV�%)Z#����PX�"�EXbKB�J��(�� �ږ%���b�Db�k�S���X���mb���4ʊH�D-_JZ�A��tē�y��0�����w�z�\*��TBW8d�wv�X*�W��,h���q۾�w���I.h���~���=�Jں�0�j�b�{Տ,���`Bψ�Qč�j��LV?]��nj"��ܞA_9��/g�摘��c���~�%�:�:Ӽ��>wC��׹�U�ܿ�ŮÂ�8��+���K��c
͏g�°��J���b����8E1�0G4N0ψ�ś�(��N�c�9�����L�y~�*/h�^9]L/�ڊ��h_\盬�Z~k{,�>ܒ����g��
Yl��YUt�Bשx���*�x@���r,�7h_�dy����ɿ	;�XFo��-(8/��þS欉�şU���۞ иa�x�^B�1��K�������jP�����,�Ld�4��q��(}妓|�D�_�FM3j�=�Y��V8F=��o��ٱ�c}�bNW�>�����#�<�5dr�h��Z%��sA�~��}V���Zu�ha9�N��tQA��U�\�YN��,rSz:��ȒNV�F�L��1�`*��zf)K��Xĝ����@�p�9��y-i�<���Y��w���&(��a�����b��b��p���F�-�L�[�M��ѝgk��6������:��[�v�¢%����S��!�l|���.�+����^����;�#�����k��[M�¹�j:�f�j��6pR�Ըe@"g2��U�l�g��ͭ���u#� =�"�[����D�@�������+11x�(�a���k�qJH�b�m�G�[ڌ�x٢㚖IJ�b��)��o�Q"8C��EiX���F��b��~fS�+'OS���4�M�^�0^�fN��R��C~Xv���A<�|�3^r�U��$�w�h��hD�GU�ꍷ��6�1.�㴙��Y�.,��R>\z㘥�)]j�ޕ�cΞb���pάR��:P2�لE;�`n�jpBsqBХ� ( �BP�:�h&r�x4�Y1���]��\�Pj�ʋ����,��㍗w�+�@�C�13����4�M�=�����]����Y���L�';ԋ��y�"/p�}������>��MS��Tx�=K'�<+u@��:��f|}�󕒹U��=k܁+�'���K��n8�L獷�!|�{�):���G����I����d:��g�^��Ϳx��{��SW+��Y�SW���:�LR�ۯl�5�3�y`k1Q�yQ�)��o,Tjy���;�V��M��Ϯ���˾��Ě��%![�����L�
���;f��կ��g>�79�`�.��9��s�n�=��{{6Gc�3����*�4������}�$%�1t��H,PFa��w5T.q�hn�9�J2f2��muJ��� =8�N��Q��;�;�!������ȳ�q�}�&*{���~9>�qx���sׂ�S��#�{S��)�W����LCs�E�^&_��o���X�>�#�C"�n����jQ�u��Ub�G�;�7��@��gU�/�E�b-:i΁�n����A9�yQ�]��o��!Z����]tX�6�h3�Ri���M5nO��'�z���~Z�[���=��4h��ҮD��id�T�d{�R�F��0��j8x���]�E�bt�)����^�CWSE<Zw-����f�P�ݮ�2�)��A
�T�D87�"�%bqҀ���U������}��-ޕr�:�#�s�2�1�\�ֽ��)��s�� ��`��Uy�|��kb^NF��L�Y��S��|�.:�e�|�+��)�#�付��x��q)N��z��*��%B�� �B���!)��t9N�`,癭U��-:����ԟv�ڙ�^{:"~��^���>�!	o��b��y�����z�HQv3�4��ܹ"1�'�H�Ǔ"�)�������>&�z�]����O����O�׳9����Y�g�hy����j�<R�Vc��;�^c� �pV�jļY��൳�<�*��/��%G5l�{���E�3%�o`}�A�Xs�ױ"!y���� n�
d�V�DfR�Y��D������)�ZK�b��s��pxCH⾡ >O�\Qr߼�����G�b3emߖ�wv���<P�m*��uL@6f���4�*p��1��(�����i��@ୂ�K¶X;��t�:��%��P�y1i��IF�{��=�Ь���yX��wE\ʢ1ͽH���՟K���@�Wi��f����ۜn����E���z�*C��kJW�j�/a)p�sq]�UNG1��toZ�Y���.�n�H�[ي��b��i�)5�u�5�nw�;Vԗط��6| [�e��g`s�F8���
�m�a�+Q�c�2�<�ս�RO���c/�y�%D.�ϓߍu�'̱=馅�8r��oi�]��y�����B8�ߢ^g
�ү���Lҝ��f�{���mKs�j�f�8�KsQ
s�*���w��R�}ǩ����ɝ|2�wl���qR�A�6q|�V�<t��$&��F�Y��_3�ʲ�䳹K�X�@0%�^�,bNÄ�b����V�N
0b�����t�.�#�7�NY����������F��x�n�5*�w؃׎���{*�'Ӻr}�k!���OxS��s۔�ۭMS��E^�q�r�1��q2󺭽=�a��-�U������'@T\G�����`���AB��A��u��+��q��";4���{��z�Vvy��r���Ë�s�[
�����$7c�{�_��b�ܽ�X������@�nm�k2����G�^(��{��������x޳�`�����E��s�8a��_��]?��{�H&��8Ѥ��Cڞ����+�Fi��.a�3�;e,��md�X�=Z�B}�qw�9@���A�V�^�C��LOCs 0���w�[�r���T�{n�gM����Q�>�U(K���=�+�o���~>BjN�;�6���ٗʦ����;�9p�\d��{��{���.G�g�ua�Գ�:�1B�ϔv͊������ivoz����l�ƁO�`�h�a��[�����FWj�ڻ�� �i.�]E�8��܄]L,7j*-4/�s��c;�Vv��LN]��|�_�z��!&4�f�z���΍E�3��\oc�����@j��ƛ���צ"�sֻ�xn����KA�XU�Y���'?7m��B�5�vMf�G	����tGf=%�]_��
�f]JH�s�N�wJׁ�r[U�]��\v�
9$Ge(f�F��V!��EX��re�+���Ģ��P7�yWU�X��C��|سGL�*���U���8*�L�O4	OmR�|.̥�̒��m��}���M�ݬ/����VZ4���{�fW��iM�`L�*�k�(}�a�݄)��J���=X!CN��Ӂo<�l���}#fj�lQq�1F��r!�m�g,ot���,�[�9�Ҏ�3BS�uU�iש�a9i�ѡ�4��ώ�b�=POD#��W��z��ZU'�y�!�8ნ�q�H�^������8�3�J�0$�j#_d�Sח�oM�l���([���WW���>�Q�!�	��5�V�qjoY����-Ν����n���#)�&5(8k�X����X��(+}\h_\]N�{R�:�W����p�k��g��_���-���0���������/���0��H�8����x\�wd����d��xw�%���f]ҘT9q:UC�.��%Q�u��<�����]h[���7�ܡ������w�>��%�@��,N��H�]Ӽl����2��g��њU��X:���3��"�Qr�vN
gqƉwz"�7~�@�=���\��K����]yo5����ȁ��*���ԸfԨ��"�oȈ��ǽ�G��	���L�s �q��B�����=M6�{;��<���y�1t�<�2.�V�+ћڻ	ţ')�q�>�ҧV�:J�˔gWt��㝇P��SX���G�h���Ɏ�?�8��}A�L�Y����5��gTŹ��(-�v[�u���(��J��um�/ð����*O!��d7>��8x��z�DSOr��Ma�q��^�u�G�JQ�8�']����'�����d?��Y�9�N��z��q7����]�+PvX�o!��=�����驁xɡ��5���c�-Ю��b��n��rU�1�9�I��r�<������Qʸ��lLU��Ł����qx�Փ͹�������:^�Wu1s�w���h!8�lC��"��c������ΑOk�Q'c&F�Vr)��)w�:����@��-k��N�ctթH3n1΁�u�:	��;E�S�c[1�;eMcߌ;B�P�>�}&�z�t�_[��u���ޯ���x77Ɨ-Y�c2ϻ��>d���Wyߗ%������ #H�����r��y߲i)�i�N�v6�"��y�ʪ���Ġd1�+�Ƴ������'M�u��S����}`�쏁`Wt��X�+��S,)�wQ��.\�f,z$�F2��}��;6���YJgvQ�����`f�9����}b�[�N��.RK����;������v������u�[X�m��Uc2Vq.��ԟS��%�S����+����;����� i��\�sX��jܛ��Z�`,R���L���1�\�ږ�I���APT�2m��*�#.[W�_s�\�FK�q7�v\���&U�.��<
/��L������Q(�(�Ց9�.�斐y���	��Bv��:����Q��/$%9n�)��l��*yM
\��ЪW�D�g�S��(?uDz|}<��`�T#$K\~��\e�y���O_�ReL�ʝ��2!j7ַYyW~���4D����d`H⾯���1K�,	m���^�*c*��s[{��70�y���ɔ >�b�N�<�@�*f)O@�����S�����7Mrj-o$�^M���j��8���N��lL�F@�{��1��hvx�=3���d5�w��;tڞ�X�φif�֗	����oԾ
��ۜ�u�U�b.p���fo8W�9ٓ}I񘧖X��a�[�:���у{z����c�ddu�W^cͻ���[R�&$~�j���>,`Y�4,�P�Ϡ��8k���Cln�:�f�^�N2B`Ż,u��̎2�*�6�[{��M�#��=#P���tT8��#n�9�]W�
��U���qڨ�"����`	�i��/lO�O���f��|7��Ν8�W0�1+��o�x�p��B�����Azfӽ�]	�ϴ7Ӧ��'mh}�t��,X�����_a3�/f��-�IA����nߍu�>e�=馭�Ñ��!�=\�h�}y�j�W���^�6�t`(�0�5zf��H34,O����ڗ��k��O�Z��k-
��評����ԑ!&ش�Cn�j�`uCma���{_�P�5#��hp=ŊiǙ���z�M�q�R�o��r���������T6'��Q60Q��`���u�=�i&�xk���*�A:�%�16�p��w$��-Hq�L�j��`:w�L��V�ÏTݖuF��)_��GK��:���ð*��P��F�^(��~�z��S��2qʻ;��[�a�~�#"��������$b��F�Xx�zǌ�zT.not֎pd��7`�v���O�Y�}y�׬KB
�� g���9F���A��
���㻔�y>��Wz��(���(��S��=̓��p�g�ฮ
Τq{�Dy	e��t�Y��)m��*Jt���$r�q�S�]��ԼO��׻�����qq(Я\;�������5\�^g$�8W5֓1��z�vĮ���D�)M�ӆ�\�&[�-vY0>��uun�'>�lǘ��
��^�ն����n
��
inAN�-�;���GWY7���[
8�Tz��`9y�_DlB7B5�]��+jN3�U�\����Ω�v�}�p`ĬU�9���v`�Sr�w1I��<|h��#t��XMz�g�Gޭ����G2�FFÁ��0��]dn�qQ��:�f���#��ŷj*,&����sk6ye�����ZG+&���TҸR.Ƞȳg��'�X],��^3~̕�V����:�[���'������|]�ҵ9^�KA�U�~H��1g��t���x3�tyj���Q��o��_Q��-�v_���o=�����ٛ#(u�My6W���G՛yT�Y�;�WhA��!<i�����͎:lk���0�����39�;�+��N��2�;\�ml�S��&��B���-�;���r,:Ӄ�[Vb�������͙�2�z�CkO�G�r~
��0+� �E�ռP�f)K�b�,Oyƙ�8.��y=$≠m-%:���Q1c��	�MMB����:
0�NZ�>�z�����������D��o���p_�z���6���ԧ�5�@�>6�b(ZV&�Q�նT�<�v/^vDt�c��ח��`�9o#S8�c˴U��}X�C�aB����~,��b�Ӝ�ݷ#���} Ũ�dM���r�P���j�E��g �RE�݊7��o��kSd�̫F��8��cJړH��|�����2���n�3�4Dl�4��Ø���ܷX7^.��B%���A��B���]Y/
�ֹ�1Yr__R[�n�L����!�\�iW_Y����Y:�8�J�ɶgF�� �g`�����`���n�������:��L�2�s��ׯn�	|u�M��8�׺�v�d[�G*1�΅W�T����s߫��5���LՐ�y�{x^`���>�F�s��ʪ���=c�2"Z�ڦj�E���ޕ��Ő�D�=�U��+]Rs�e*Gx�6r̕y[���>0�B+WuR��5s�ϳ1�%������ͮ�D&�(��s7&q�NU*�]L(�J�&�G��]�aL�7\��#���|��Ly�-8���oBD��4k'�0���|:ɺ�h���yMfaj���9��H]�)'��&n��w٥�|�� ̈�6&��F��b�z[�b�C���Ρˉ���w�oX�s5�AÓa�"�'�����M���W�/��a
5�5t��W�­�jܷb�Mn��橠����4�޻�
�h�Z�+�g4xwP]-Ŭ�Q��.Ulr#lR�݁�g����-��\gEL[��4�ջlL��IC,�����`hسt�"#�ڷ�M+�i��n˟@�)6.�>�utl���f�^r��6�vU�������!7� N7Y��W4�vH�mm�U��.ގ�]ls	\;D}��2%w�+��^<*cx�����s�rUǎK�q#���/�����k/T�n��nF�Z�P�a�xVM��N�)8p<����}|����t�����MW��`˕����|Ӓ��6���n�ӫG��}�܁�kҒ˭tz֕�R�4kO;ֵ�2A�7ۿI]2Qg�V�g��;nͼj�Y�1�;��_^6�0͖�s��۝��:�U�/�L
 Y�U�����YL�j�;����s:�>��%����׍�}/7�G6��ճ#"վ���l1|���3�,�U��<���1ë$���@��ǥ�6�o*�=pV�ڍ���S{o����(U�KD)w>%>�{�v-�f�W�.�pF�aR3JL1R����l��"��zR;S�c�O��{����r�PNѵzկ��Bj$z���[X(fj�=
o��p�Իc{۪��+��c������m�;�4�ˤd��/��n��7sdh��t��6��j�oN1c����d��u�u�Q��4��mej�x�}]�	L�ו�4�ϊ[�5*T�ݴ��]�ʩȾ��ˋ��͂(�U�0BQܶ��ZEn	���5|\�f�稻�-����ܥ�������YDFA���[����Y��*�����P�DX��Qݬr��cr�X��H�Ym��F�����kP���*���[*���T1��ih֋Ub���R�[A��rU��ʪ�d+*&Z�TSMST�DU�,b����Z�,B�"+e�:��(-HTQEPb1��1�hȺeH��6��UH�UAdke���U`�1d*V*#�QU`��iib�"�B�u�1UAH*�ɭP�TT(�Y*��DV�� �UTĪ��F0F,b1Tc� ��T�EA`��DH�U&ZE���TLm��*�kkA���!��AE\�X���#Uk" �VX�2�R*�A����(�-��-[Qm(�UKiiT��U�k*����Y+Q��YX2�Tm����+H���=��7.s��%�k�]�gwgA�o;��r)�/���gV^e��J��U2����p�n=�*�^pApv����;-��Gw[[�[?��(P�����coƚF��g��=� �S���u]9g���q���M�7�i$��ޛ/���W�;���3��)�C�uL9P�
��b3�:��J��f���L��n(f�[�:P2�لi�l�����BsqBХ�EY7���|!g4�{�똈=�.��{6�`r\�9A�����m�Y9�gq�˻����Xy��U���$�[���H����@�d�̫��D��Y��C��ǥ���n���E�X셱8"�*,F����@�C������+%r���=Ãh��7���H���ﺇ����u�G��v�cS�Ĝ�N��hWD�j"����a{Ze�E�J=6�2��/���N&(>�0-��i`�MA�x�4<�f*!�7�r�����|gt�=D;�V�@�U\�귀��N�N9v�e	���Ep�U�����\�g'"y;߰�=��8��+���8�6�<�E�y�=a��xQb�8t��9<Ɲi����lޛTp$0�����lI���UM����Y��~l.����(�Î+�뒬�8v�b�4�72���J]���y���"�ԝ(Lht��4ﳛ���L��!NtW��q��y�Ee�ƝF�$�����֬o���,��}���ʌ�P�4��mz�X����)���}{+�X�������&u�
�N�7[GIq(��.�=��H�vf�9O���&�z�=1f﮹���wX�-i#+��[����]8�*��.Kq24{�R�4�0��j8x����r'��E����˿z�ԑ��I����9��k8�hwk��:m���Ppc_X>;#�Fh��U�^�ӝ���S�*��޺ߌ��4*}��,J����Ƚtc�}R��&%zBZ񜨉s�\#�I���Ċ١F�NnA��&)��i�1�vd���{S��B����U%7^��]��٘W�#ĸ
g��Qw��gx���	NF[�|;��u��6�0Ď\�I8�k�>�X����|s�'|�c$K\~�}�����Н�z�О��X4r�qp�a�O���X*
����dmWh�'K�2׼������~8�-�����Ṏ��ݸ̪Bq L`;�Z�C�Q���Ѵ�Y�t:��Q�^�3'�	7�.iV0kχzz�U����8?,fZ^믮[�/"�$�n�B�=�t�h�oc����Cs��s���wK�G'.���i�L���D@ޚ�=����.�A�6�x�'����޲h�ңrh]�R�Յ.�����E���4,��Q�tp*g�ɉ�|-{R,��V��O�;<f��(�]�;nj��x��hLjY���08�s���ceÀ�H��noj�E�Ԯ���!�=�G6��O����A^��[���^4�|~��{]W��������Q�{1]�δF4�ߞl3��M���I�vP��p��g(gT�}w��mC�j/�ڮֵY��N�<Z�]ڱ��_�7�߾l�pK�C.r� o�G*���V�g_�|��Ozi�-�Öռ�ϫ���Z�V�5sJ�ޯ&�gF���W�iN��fj��+�PQ�~
�f�;�`|�>���2i�q*���Y�bӭ	���8s#�v)Y�[�T:H���)	�����[�Ǜ���T��y4��r� dS�����;�F������D̽	���w���o7s��
aC�(m��%*17*(�j��.��R��An��;*okw�ݵ;���7�V�7�PeD�Ф��Ù
=�]���^(�u�J���$aθ��`�5�f�;��c{�=g��{3��;'c+L�U�w¸��zt��$6�k�_nH�Ecn��sY�zY4Iݬ�21���I�4�v����IOru��x� DH-�B���1�\Vܱ���w�{����LI��#�+٪����?��g��٨��]�$Ϸ����_�/�ZA>�������^��M��A���8M��zK��v�z��m�8��Ȭ���J�������3�F��WM֫tz�>1=O��іE�K,T<�	΂�(��N;�=̓����k�8.)�vv6q{�_����oW\~8+xg��^����|���'*�(�t'����Y.2]ފ�;Ȭ�8�mj\��-��ڏL�߳V��r�hav*��sc�8ð�9�ܣ�<��N؎��`�����������s�%��?X�a�Y҈�]qѹ~�,��u
�U㑀��_���vgv9n�u#�y��T%���X���W��	41ś6}�[�+ω�V~C�z��ޞ�{���e�3�cT��yOv�u^����DYvWv�NP��ZZʀ���5dN�şU����*ڼz�S(��T�
��OmC�ރO��2�/2��KJh�2}���3�B�v�&���]ϗ"[��)Gt�*L_�U��}ʃ�p-�ý�p����:��󃣜�7)t�(��K�$�M��c�;���W���F�v!y�{`��������Q8��UJ��s��6,,⠾to�!Bk�)D�i���iO
�(p]���#��Q�-�d.+㵪��Y�,|YF�Cy���I����+GsY��Ͼ���8��)�,,�F1_���Fu�1	OLӖ|���a9�ZpthmY�S�i+�.a>Q�i��M�hi/iz��>0�pT�CN�z��|�)K�b�,�x�ǻqɎ�*�f��\�SiJ�n�@�ݨ� `5�:���!o��`�1Ƶ��<�m��5���q*W��ۖ�؈�3TXx�́�A�	D�3�J$Gq0���M�/)L�8�	�ܴ��%#:S�~Jp6)B�-L��vv�t�*F@���pU!	eط5*��T]-�)>�C�9�5�EFzѳ�߉N�eC�sQؕ�	�*�:.rM���f��襆����/D*0/MgKs��JV[� �}���w{S�����L�iy	�(�]�[$�1L�}#K?{�A�V��>{�(g���K�i�7,S;�6�,M*	���M8�|Zܞ��_�P5
Dא�Q~��g���>,Ы��5��rE�[*���zc��#j�T'����h��Xm_����5<�StlϏ��J�Js�yQ�w/��h��Aų���3O-��%�)糰����h�I����d^�L���jv	��I��|*/��S�MfӘ+Ϸ�o����V�z<�Y��h�Zy56�O���v��;���nc?K6�t��խ���wB]�aQ�C[�
q�uۅt���QO��������zY��u��N�P��&�n�(��GQ�):�Ƨ�9��4�/y\VE�+)_
�ޑ�.U�-Y�� ��#;��9����1�Ӊ�}�`[u�梲���\]�+�����K�<�{5��Ⱊ�b�^J���e�@�!��!i��C�M����?�݆��6�>ż���b��s��.0<yZ���]>�+`B��zuȷ����k7�wqef�BJ~6���b�݊��2��ᵋK�u�k6l������J�͸�$yW��Ͻ��;������f$Fez��WDg:��}�#��kA��3���6�P�U�rR�ƻ�����f�fm�a��[�:kT�Q3P3�љ��B��Ў|���ը�Jq���1���t���McT�)��^�^61vz��{�1��L������pG>��JvV�Eޭ�Gg�M�~�v'f����Z�`,>=�|����\���qZT�P;���]N]��.�=\�b4�!r�ϟ>�m�ص&�:]�aB�L��f����F����u�N����I����t壻��C�;�ӱ�λ��#B`�8:o���MU������z�)K��������ڻ7�/6��vF1��e������u���'�`Ϯ �h�1��/��̏����r�K��J�uq[�-M^��'ꯃ���G��Z8��^���F-00��K�><^}
3��N{$%9�r�k^*{9�&��[�%���-l�@��ٛS�J���Q_��>�"Z��|}���痆��c/]�혔�m��<Ѻ��L���}��A`�+��a1��$q_Un��g�u��^@�r���o9oNYw���Qo9���)ӋB�ā1�zSU�qLh{�59a��rDy�,��9!wA�j:_���W�c�{���:#�3���/>�N�IFc�_Ɂ��_���8�a�t֗aL(b��S��zo۵�/�q�nt�yl�p+ϪU����,��ǳo�2�=��غʷtn�w�b��ⷩq�f�>?i��C�nّ����rj���̷۽����br��Z_x�<�_X���۶� ӈ`$�s����y�wk��#,N�5n���#:j-���p�,��+^3�O�sޚP�sP���t���^�H��S�;�p0�<v��+.^��;�͈�g����mKse@�z�(�1��;�u���i��j�Y�J�`�w���V�b�LG��W����c��.�F�,O|׽�=����G	=|ԇ&NY5��Mսl�>���^�]��{v�k#��6����T�in�������p��;m+��eWY�R?	�<Yuvu�]�*�$!	gM�N�ɻ��[�2N�x�f�3J%`V	q��tH=2I��GM=13�'h ��q)J�X���dS�������`wj5κ��<vn��7ҵ�ze��ِ�PxpϘ��@�w=*|�
a�n�Z��f���8Lu�:�DU�����Sdm�
��Q���
`ʍ'B����̅�.�~X�E�w�J�?<�
���[Z�;X�������ƭ����~��`���K��P	�K�鞅�rRl��s�oLs����))����p��xc�g�=4/dO�����,�>h�q���S�̩��x���R�aK���B����+��-1�<����+���Y���^�|N���Y�9���V�b���w��*p50-Nr�q�S�]�./�Xj��ҋ,�Sq���+��R�������-09�ϬFu:�@�v�ǳ�a�q��M�:�L]�lG@���Y��Ǐ]=�ر�[.�� l8�Rʩ���n*/4�њ
�r0�������Zi�͸�7��I�~��f����,;xM!3�՛{�N]��
�ۘ,�fq���ɣ�����Hm�&�
]bKHV��w�6J���M�B*�/w���_"j��+������r�w�$^�[
��/�<7|`\6��]&��g�R�X����;b��f�}s�J��:~K�t1ŀl����̜��R��6�L�����-��7�ܺP0+��j�-nvtf�xf� o����g�Y��ş3���)�I���{�nsU���)&EB{v�	T:f��*�/2��ZPh�2~B���sO�ݮc�O;��o��FgU��Ϩ1��<;ўl��1��隼w��ب�4I�ƆVMo׸}���".��*�#N�Y���!	N{���N�Ma9t�؍h8�Te6{�m��y��jqu��_��#�9�Pi!��杨D	��/9���d�[=�Ǒ˪�0e9�:Q�'<�(���BD듂���+11�B�h'.�Y/x۾�b�;5}�R�*u�DE��f,��Cm�ɍJ��X��4<�a,[�E{�9�������
�5m�����&)B�jf�]����8ʐ:��z��;�ځ.���<�����<Bv]:�[�熚�"����Ǟ6w�+%����)�_r��v������onˇ<���z�aAK��7J˔!��+0����Z��������ĺtj�h����1�A}� Y��o��S��9�!�e��̽3m�M]{�Ng��W³D���u}�{�s+���U,;����Ģ�Xy��;���ҥ'�tgP����BK5��ܱ����'a�V��5c0B�������t�eS�Ӿ��7w�3N�W���ӓ.+��݉	y^�Y�=d�,��t�LU�5G�|�q�߳���'��U-l�&�r7W>Φ������VVYP�=w�)*�T9^B��z�_L�Y�U�x��N�w[*�]F�2����)0���A@�JBQ�������p_�|��O!��VFŁ���&��1�u�����o${sg*��ШDS~n�(��B�Uy.�b1������I���3��H��[V�fjG�ҽ����#�j���G���\xD�z}�{��^�P׳�@>�Pg���a��A�X7F�ᐠf��7&8A�B�!~N�N"��5�s��,�eR�������������Ǖ��� �O�V������<��"��c�	.'1n��wvF�����S&��څb��A����a>Q��/\xgP��M�����\��-3���k�΍�|�Vjˋj��ӝ[����H�#�4)�|�gޯ��U��P��_��Jve�*��V���n��F,וqn�xHxC����;�����2���wKx�i�����r�qb˚
�%�ӛ�;�ڦ�40;yS(��R��;UǧG2�D��;�X��u6�3��+5n��R�"�!݋��OI�;������Z�V(S��֝���因�9��+Z�Q
�G����VQ3qA�ƶ�3N�S���J�"�0��5çRݧ�b�����3U�Nm����Z9�H�6+¯0d����B��#>抗�6��n|���r�d̾{��0{<��Y�:���Z�
mU��H���u���]�v*�`�O��YКd�IE����ڥ��v*���k�%�_n{U���P�?;����ӂwj�;;@l1�9��|����T`��ثUmX��=M\&6Wۜ-Ύ��+1s˼:����wkk^��?��\)���	�3	�&�55�]W��Kf�^0��\�w<�Ϋ�}@f��4>B�sI��f�B}�����`�`��`�� �'u.��U�l�ԯ9�O]��|����
�F�KY�h�1 �]���VH��f����`wJ䏺BΑ�Es�j�D�w�i���-ӻ��S��S�b>��|��8�c�Ug5n�����md
�y;)����R�[�-�T�Gl^Gc����6Έ:�[��|���T���̏-��-9�G~�Ѻ̙w�������#�1�u�U<�$!_w13��	��nR�;qh��VT98RȆ���s�v���W�5�hW����8�ʊ�vH�_ugtv���E6��]���'�v1SWY�p�gV�1�mL�X�q�Y�n���p�P<3����N�2f+���oYE�2N�b�uD����j�3�˧o[�2h��
�����L݅�B�[�Y�Q�-�阳c���!ʑ��w�\���e���׵Z���̝���j���$����V�8r{����;��6nܻ��d�t6������XqţS�c�αX#z�w:�}X1�d�/qUB��_���yR��\�pU�ݙ�r��[�1g\�� ݵ-ڬ��,;:�Ó4��p9oU��C;%`u��w�e����ڱ�"�����>�,=�hJ\ ��ǭ>��&ac;��0��7�v���xaY��vgr9W��}�w>�{S��R�
�oS�4[�tu^�g3�z��Ķ%}{���a٥a�ɋgt�@֜�.�}'{ֆ1��;�6�I�oH����=�:N��-��ץd��b�1Ƴ�Y���nf�v>7����0v{T�#��њ((F�%]��A��1+j�MV�����[I���7m� �9eZ��2Ϯ�cEP�d�n]��7I�/]u��q�t��X��Xʫ�n���s@J�l)TSJ����vC��J���cqq�8;U�{��](����{^v��턮�vѢ��U+���ǻ�Q�����,61PjT�0�ZTb!m"�(��kg栌�9E DU���"֢(i!YmX�U-*�#�eAGV��AM4Mfb����FAň*
"�*,P�"Ĵ�U1�����
��[F(�
�*DAAEb,X�IDP�(��!�P"�	YEMYQH�(�UTPST�-U�"���dTT(�V� ���*F0E����Q#-f��d�TmZ��b!X[dYQ��+
��EETUf�S*���b�e�)Z ��UH"$R������Y-�M0�2��dX��H]\U�V�QTPb�P`�D��J��E�H��E%J�(��A՗��j"�"���TPD4�b�5������WSL�"��Ac�T� �["~�H$�I!م�;��/X���*_*�8Ҝ�`[�.�y��=ʫgj��A'���C"9VÛ��t��4�,7�K&�3Q�!mOT��<%�:��z�<��9�7��c��n3�:kT�UD�@~Z���caߖ���[J�7m^o��nJ񸔥�5����@Q�O��(W����֑�o�%�g����	��%�[��aK	ž���%bo�0թ7;ʵ���(\�L���b�t�^��sS�C��nG^H앫bX�Pu�@(0%�R�c�#=��L�Y��|���TG&�F�|2��c[�������+�k�^#�k^��ۘ�ӋǼ��9gpG7-_���;��V�\��;ȡ�TG�w�9F����
[��q���>��p�8�O�l�y%T��P�U�1O��x�1@����<�|�8��@|�s_p��S�{���六��~�INz�rɇ�S�2D��:��J��Y8c��שN~~�rrÁ]{���b��Sy��k����7�i�/D�f���_�F�[g��u�V���!(�cbh֙w;ӻ>��a@��9�΀Y��,���=�V���o�9{M7��\25s}�|�%J�*{����`0�&�u�e��`��o�	P*����r3��n�ܵ@I!��4�EV�D�ޘ��'dj[�������e�.���Zn�V�)�:��8fC5�;��[ي��YD��+b�3x]Ob�ܦ�N)���Ө�=�r�{���-Uu_h�۬��u�Ahz�����\i�L��}������[��3��γ*����]���)}O]���7`���f��^1`��{��c�c���Q����T����ܒ@[�u�c��J�`kq��5�J}�ϓv�k�I�6e�M��b���8]�,-f���v]\8��<v��2����Lҝ �б>�PPݙ��%@y;���D�sЦseګ��4�X�BX:lZu�7{�p�D![�ݳ*�ޱ�me�m���ɉ�*pU}BU"�!A��)OU�\�NVb�,O��c��1�E(��Ɩ褔���㉿`�/�8P7T����2�OyX�;����	��ۛq����s���){���{=������3��+����68���N?ίN3ß[p��U���S�֖����8�S��cY�0ܻ�g�N&)zL
,BX.Ř�8�n����%_��;�t�}Z����0\�c�3��{"�1R�"<o�Y� �����䓋����Vl���Bh6��;6�ڏ^�M�Fr�3i�
�jNKq��i�}�}��ؽ��'u�� QTS^�����5�h�z��:V�@S����I�U,G�G�zW	��q�K���T��Q�D"�f���e���q�C(�'��zU�A5ʹ�	��
F�g��Q~b���(�B�wOs`�n��]WU��/~˿"���ȹ.r6�?/ ��|ٵ��Dy:��߼���'*�:)�O=w�.K��w���\6�{��u<�s��n�k��_���CQ���g�8sC�V3�#׽�Sr��<��A%uםzgL{ė'fq�7^�՚��=0G��f�"���#�p_��3�Zuh�^9im�^8	��M�\^,ԕr#��\����2*�{α:Z~k��W�ca��lo��6KdA���;XR7-�ܨ�UhO������;8���+S�=����;�F�|}�3L�s)�[)�Hdv���ݥ$Ȩa�=א�;/��[7�]�M��^��#(tء�+��cx#:����7
Ѩ�%-5�W�Zr����sկ�OW�o{�7���I�Aߝ�����j�o�_o��.{�b�y
�����4���!	NuU�zw�y�a9'%N�Of�ۭ.Ӯ�\J(l6U���{_��#����"p��=\{E���ǾM&�Ų�*Ⱥŕ�s$T�gQ�%OG�O^�Eb�,z�t>��;���|��j�	�-ZyՎ�WS<%��We�it�i���i�u�'s �pcuN��������kRGH��h��zu�Czj4=��,>�2� �*�&����輔H��F���(��N��:Q�'x�b��_� ��j8xG�J3��g��M��K;��ln�ԲZ䎎R���/D���:�P%��<���4�Tu	�,T�#$U����S��U5�l�(�`�0�Q�նVW�gb�,��3��ڬӌ��GA�$,�;<�N�&��}� ��*},�)�5�EFF�9b�_l�LK�x�&ewJaLFX�{/pf���h��� l*��Y���^£��Y���:P2�����w�>Co�OemQ���\�x�k�p��ڕ���2G���FuU�2Ϟ�
�eC�!r��S�
�uQ��-���d�,�|�K���3����\�>q�=_ <�����n��ວ����҈+*�"�{�c��{����v�W��_�@��A�6xR�o����ʂ�^r�VY�Xy,3��*��h�ke�L(=��}_ܜ�;Z-�9�8<!z훇�e�Fǖ�)�Ł��n�K�t�� �U�s��yk��,����3�ESYӈ��W�~��~<��Y�N�=y��|����[�
�6�=��K-��t#sY5��BS@Om>�N���#�M�z���ݗ�,��}}v �ҏ^�{������M�q�[(�^�����tcC�9輫0��'�]G#���)�e��N�?�@�b�)��)x��u^��5����w��P�m�gW{��M�K������JTV	�[^�%F���q`WWb�����~�apt�bk�OJ���O�皧���Gͭ��QoÂ�A��+9�_?�'�oԼ��X��#;�6����L:]������\�w��6��N���@nof��;�@X�ؿhS��Ͻ@I�^���Tj�+9��)�K6�ڻPD�49�r�S�kjﹽ�ȡ�=J|�1���Y����c�g�5��b�_�gݤd���:j&�(\�yX�qB���K٘1��L���Jfn��N8����z�|��m����N�v�X�V����Z�ab�,�L��F1N����U򨥉�T��7�N�"\Myz�R���NhR�xg����H�9�/K��C�*V�*��fvt��y����+=��~b�qV �F-1��:������<p��w��3EaP���w�������!�{@���`,�6��y�yz5I���e�D��yD�%���~�a^�-�G�"#�u/��1c�c�����4��Y�)�Yd���;2����PݜN��z��@6 ��p���|.D�$ᇉW���:�ltݍB�˰V��]�*�@f��⩙`\s�+��_� N,��ؾie�G�:))z��z��(�}~�ݍ8�ĈAȔ�t
��t�f/8�D���(b_�3�����XQbc�ʎ��u�H������U�h@w�4�N���Q7L�׶s1��[�1jE��<6������J͞7�<B>�z"�;ӆ/ZE�"ͭ�sΦ����aH��l/K�F.�
�14�������zo��q�nto!��4�:õ��<����jޏUs��D���Q��Z�/5F��a���C��C��4��
�r��[�v]���L8=y7W���;��uP��N����J��۪��zՑ�ݐF�Z��F���R(��8c*�W����:R������
,e�Qz�R���=g�yc"w
������m�K������v���^C�yך�ΌL�0���+� �Չ�Π�O��F4�\V�r�(���3Pr%@>�BY�bӤ�dF�0����R�R�+���*���^�����c�*c<8�a[<t���S���dS��ŌX�޻�cf��a�|h�Ҙ��`�ѓ��o��Oֹ�(��]x��<��_v`�U�IVS�����'���{l��h������%�:�i�Pt�;���hb0c�����3(�gN��,��3����7#�:^��僌u�2j ��]D��ͧ0�$K����#!^�ҿPzt��5  �=*|�x�͹ ��.�{̬�#yY��r�ܦց��qL��;�<;ا�oЦ��#�U(v*��Yt��VBw����.7	�ηn�J����s�S��ؘ����e���O�l{��3��%�z��$�G���*X�A����F
}����J�������4s!0�k"e����.���b�VM����
,i��nt�
2�S�^�A�7y�F� s<R�4⬕���mP���������&O+�Hm�ʯZ"r��i�O=w.K�<_��/C�/]-����2����miO���'Z�r�
��i�֢����ee[���ow;F�>���@�.��N0�g�#Ի@�����f}W��+ď';�8s�ѣ�u3S��(�GZU�C�Snqg���Y���:~J�! �͛�x������p��[�rFwdj�Hq\efJ�o< A�ј:�+Xҵ9��ْ#Ӛ+\�.��7ytȱg����pt�(�{ү,.��ζa�.ú�f a�w��u����'{}�����&���;hw�(�ew����Xo�����Å7qc7:��$Y\�^e8��N�S��p�˗��j��zM�Ui;
�悘v�.�y�z��6���$��Q�%�t?P�1Y��xnӓň|<�-���0��kjU�^(e{����j��t\C��]%@:5ુ@L�ѕ;s`ARc&�q�C٧�<;ў�)�ڮ����h��:�����^�_����B�VGO�?���{�nyz�z}=K�j���^��[�w#�,uH~4���1KY�E]EΙ���c�8*kH`D4�s�Ƿ�n��ZT�>��k���8��17n<�9V�����ޮ(�(k���m��b���9�u!��˳�q��B���2�5�V�."-M�Y�y�0 셁M2��#D8F"��eޙ�{���y�;�blcX���b������(Y-L��G*��q� t��EE=3
D����hۼͮ_R5s� �Q��\��pi�r*)0�y�t�2���F�"���&SJ�[s,��)Ê���u�yq�b�?z
��H���{�z������S{�4��[�������T_u�Mx�(X��|�X?o�O�:��`�㲈j��tZ^��݁�9��xB�u�i̱|.c� �v���g;�/͏�*�w�]�-ZҎ���gE䋅9�kz��WGд/��Y��.����|�\m��l��	���r���)�� �F��`Qun��\�v�sV�ʰ�����+uw!�b��P�l��x������#�͇�(�2��E`n��C�4�Qut6z@s}j*!f�E��z�%YH�[䶻���!Y��bܧ!@"Z����.{��8/�|���;o�P�4�=P���Q�X�~��>�����Խ�����/|�����R��ƶ�vV�)��C�K��M5�x�Wa�b�`Vc���s�Gt�7(�yht�b�}�`^��3u�轋���ҺQ-��v+����|���n��G]"�۞��(C`��N�NdPKvx���$¡���ږX�5p����^��N:��^1���`E�O��땰p>;n����^��U���¹����1G��Z�ş���Y����\�;~���.��T7e��h-!>�{Ò��~��٦Kf�c��Zt,:ӝ}��:h��_
r�}넣�f����u\��p�%j:9�1�Wj��^O9�s��"t�Pvx�ي��6��t��*gWNj�ވ*d��D�5�m7�m��-X�R�K^9;*$�F0����h�I��Y 8޾�uxv�8Srf<���']��]���j�{
��9�bْ�m���< K������9����f����W�f�#�Cz�6��we���m���{gX�B�w��0:n��4�\�;.;8V������8��~7`h'E!6�[K��5��5����j��<�b�����nI8w���C����n�ԥe�q�k9���-���M<//�f��v��cQɼJ�`���5!�2rZ���oDM��x��q�g�JJuc��V|��G��߱;�a!{� �`P��ZWP҇g/6�s]?BN��7���SU��w�o؜!��j�#%+\�4�����l�ӛҴ�R������9�-:�s�lp�?e,�Ĝ��l?�ՔM�^YHzښ{���}��������w�q��aJ�-j���2�5@�u4����4/+����_[���ȷg/���=�h����&��t������OV��[uo��:M�]�%)�_�}~}go<��j�Y��z'v�V��Q�;\��K�^gY���M��������K�wp�T:��+vv��a�U�䚿:��i{NT��(�98�T�b]fVk}Wׅ��kV\� 1;|ZI���(�����U�f�_i���,�s���q�k�tZM۹��\�3��w����p�o�gl��V
iI��g+�Xū�{�����/�^�YE��ځ��PK��hc\ת�Q�)�Ȣ�5�T�m��o%>����V�t��{h2zUܬ�SM��Y�S.�����>J�\3� �4��9����濗6�j�ЮoIn����++��<���B�"�M�@r�5Mڱ�z3WÎ�)�kx��[�K�Q������T(��[�aU�Mɜ��e�Ň��\��k��C �b���%�PUᔯ�%H����K:1[�)�4]]�3��y�,!.GKy*UIH���ݑ���\䖍{�Rr��\�LB�CzW^�����!f.���ۧ���Q�zEL�s���K&�v�����i�5%��X��'�ʘe�6{���O`�6�æ����]��m�[l଺"ҭ�#��������0���x1j颓�V��m4�KD�Ɗ|��� ��:���&F�tٹs�C��H���h��=�У�7���z�b�6 �e�*�6��aN��\�i:�0�$Н����B�{|�S�k�m����YI;Oc]t�u˙��nN�P��n�I�
��dأ�׊���F'>������-��%ڼ��Ѥvܘ*,,>�A�1�$�vGV�a����W�`����Qf�!h8yk��y�s�!8R�n�w�O��t=7�o�J}&S��磫�l�ۥU��Z��i3Wj=��BS���+Nk��<�`�@_e�u�%�����o)VH��r�
���dJ���Y��J��O���;�o&_,�WW�������s�q�s�ݪy]Ң�4%���Mbε%X�w�V1w��s��Y��/u�a�bY�l�NTb�kL���}יgQ_1�f\h�S�wj����N��ֶ�q��X(Ȗ@N�4R��W�^���:���y��}$�2q���H-�opw��b���Ug��zIQ�G3����[AӔG���*�"���h/�ʣ�%[�w\�9ֵe�5�Q�F���-8g��5��7 �����=��n��d=���z�ч��*����ONR���M�s���66�t��G�s�8�Ң���n�7:=�	q[�kk�f�[&�` ��.R�A,�-�96J��+����#q����������l΄>�`���M�O:@6�_<�ebp��53R��@ICr 2�l�3!E�V�;+f�u�"�Vٱ��x;Z����:���dy�ʵf_3*!
��mh��z:T��ㄉ�+q��<���֌�T�.�N;S��{$7�<i�Iڢ����~2翾�﬚`,��cE�"�*��U�9j
�Y�UV(� �����E���YDQE X�QE�QAVV��Y(���X�j0P�*$m��(*���AT�#PUZC-PKB����dA"Ƞ)eU�(�)PF$m�(EV ���("��J���
DEQE��R(*����
ȱ��DTR"ER
EDA1F*1UX�ԭ�2#DQ��QV#�(�F
(��,ĔE�j�Ȫ**�E"�F�DQPEU�"�Ĉ�EX��DV"��*�%Um�
 ��AUDX�[Z)����X���FAPPDe��"�Ƣ�չJ���H(�F�2,�X1QVEPTV9lAX�F)���x��up���F��3{g:�w8��!9+����:��{���nҧ�)v�Z��%JI�Mπ��	%���=+?{�Z����9���0��C]�d�ś[�9�U[܊^״R�QJQȺ+6R�5�T�:ګd�M �G+o�m��O��I�fO6�N�C�N��R6��]R�2��,߲XK:i<�oi۝;�sq]���C\�S�������'iʱ���V���Yη�eׄ��(��7'�ч�<���4R��z��BH�ъҼ6�@��
N]�Y����ު����[�+���X���jp@��̼��-η����˝�K1~6�}�gƳɥg�z�M��^C�^�^�ˑ�uSK3�*v����ѮwS�]�i�j�.���a>Ճ��ϫ�!é)�ϑ6�34�fz�|p�\�T�t���9�ZYY�eߥ��m$#�O�����"KU��09��z��݁�:�(u�5}Lp�wv�Tt��!mt�	�hF��#b7�(���L��.x�L�>��/r�����baЙRӘ�X�In���U*��\�KJ���pޥ��$�B��q���E sB�jY
�Z�M\�̹r�+rW�+��@�{:��S�&��>�ْVn�u;�۠�<R�N���7��z��;v���a�+콽�9��#	&7��$5�b45$)��TKբ�k�N�MU�m:��MB[��m;/qL6��M��͆b�����Bw[}���J:�kv�Wcf���oa�����-%5��x��յ�\j�wϱ��u��h�bo��ժ�b��m�&�y��kf�ͭ�󛢬�<r��'�5���~���	���.�^ٿd��ܘvu��;=��Vy���(��zu���б���:�1a��_��O�{`�û
��}����f�u�n�KikmXS�{[FV>1V/hN6P�<h\��̻�)E������ԑ�I����D&��:uhRzN6��`�zF�uKӶd��A�B��f��p�T;M�M�k1j�����ǎN�Pc�"����ɩx�(��Wk�+���1��؎�xșggg72�S��N�Q���۠��sl�s�N|x�;��2mh�»��k/��2����d���w����]�oL�-}`&楩���*b���Weս�Л��Z�i"Y��Js#��*����6�W���ѪV��&树��ߛw,:���Yj�Թ��5rV�1^�R�WT�R�ya�h�%�z�7�����]�0���.�䵮�_��/q���U�-�<�Ns{m,�Q�[��\U��b��ɸ�h�ɲ�AC�zAjA�U�5Z*�<�W��j�{g��_���o���K8Û�8q(j���!�գ%��i������Kn]��q�o�K���ܴ1��-D�p�����W���75����XVQ�3K=����n'ő�D�j1S�*����f�v]��r*A,�5���hf-�f�W����_[���}gnAQu���>7��Sv�m��a=<�D��v.PS��Q�KEc����ͶΓh<��A���-��:����z���������׳\ȮuÝ��b̭��ћ���	�T�����݋�v �����6�����ĝ�;8�����*�i����T�7�V�+��۵�|�Y-=���*��2g��U���� 0xO��J�=]���� �)v��h|����������kɹ}��󡵩�7S�����*�Z�7���M�}ї�s��[��{�N�Xn���y�V�PB�D��L�[K�>)ym΅�u����x��}����c���y�w�:w���9��(X��)-l���TI��|�ﳳ��KKbSc�ǁ�v�N�
OI�ىΫs�v�oR}"K�v꘡$����k��c��cYK<�k��샹�M�wW���S��L(` z��ߩ	��m,4�O�q���ю�#6�c�6�I�bחv,
^���|J�S���d{#W���Љ����6�wJ]�i�y+/�_���ĮVzJ�V*�KW9N	��:��;�ҕ��Y)�K+ ����Y�w�x��Aj�*�Z�P�SwڹN������)W1��ib�[WbYÞn�N'�&�6�gY�S�'U�$o�>�3^�n�6��;8W`KA��<������$�,��;��[}mz-J���]�H�'��4q�;4`M�o���ѡ�2���22�kxu�u�q<�|ΡC��"����"x�1������v`'�c���p��^�:+k��ut9�i���L��1-��ۮ�v��7bt�r�wܜ���}?hQ>#�MX(m�4zՑ��.%��u�훰9�6�6��q�lz��AV���N�֎T4_4�~�V�1+�҆m�����vY6��[���C�R����w�l��pu^#UN�x+71g1"[��1g1%r�(�e��a��>��^ɉ����0g��]ΒZ��ZBN�V���UGWN+��s�������c��;���M?��F�Q���� �
�Is���V�VO}�6t��j������Ky>\u��0 q�{nb�Ht/���79���%O�I�^����+,�K	gM'�7���r"w	U�9s��ь�t����2�6T�q��K*��Jƫm�kvm�Rb��;Ɋ��V��v��������W��:�� 4b�L����#%TUfg'�_$w�?��(����ǎ^��ZX7�;R����\Uzz��˽A]]=�/�7�����v�\�@7'��
�����Q�@�%i�a19�8����� ��YK�����n�f�o�i�u4���'��9S��]���5��f
�+:ɺ놝����U�Z�w7�i7�	;����h�G�>�V>X�g��Ʊ4���u��mܼ�{���"(>�Y��Χ�nGq�'_@8�U��dV4�5H�Hd�}�;ټJ�f�f�uD�q:�\���>�bCJ�*��U�>V4�7�-,�e��ꬪ�8�q:�UR^9�Iy�`��q(i��o��Yޘ�Z��ay����V�����2�j����؝�N����r�:�Pr���YuK�
���ч��}�7�ñ��������z��GE�X&��{o��-a��+�+O<\Sښ46��ٿ348:#Vm����^�3:͌{�˂���axK[EC���h_-B�Jim��%}4�ũ��)�Fmm��.N���8+Nc�m���a�=ְٰ���FJ�۷����-YT������N;XmU�r%�90��]�k�7���4c��Z#U���E�[�ftn�O$Q��g^�1����G҄j����f���㎧�R�"�
��|��r���:���֊]O��t�Ž�R;���+w�:pa0R�u/���ō2N��[ܾ˶��5�V�B�yo"R��Ѱ�#��f-�Κ���/hh�@N�y[J��͌�����Du�iT��M*ů��8��ӷ:w��e>0}b�q��O^�{8�7���_�����^�3�&1<�-XM;t�Ф����{dk0i�/��Σ���ذ�'�U�la�ރ6�1H�0[VϜ���I�f�E�`�sķ՛�uH�`H��tċJ+��W�����L%c��cY��_U���켒i�-Nj�bI��W�T�(�,��a��=������.�u�n�6T�!q�.���E����5�+]B[�����Ӝ�950^�g=��-YN��y����B
�H-]"�X\�zfW@���<���Ie��
�{�x���ܳ�=�M��W�$!���R͓�l5�<�s��B���6�D�L��Ǟs�h54B����l���3����(2����Ƴ��wn�m�swJ.x4��lYSw&M�ag��x�w��<_�a�Nvխ��ůdW�3������=��fm9ۮ�Q�d��|�o2S�� �����&o5ٹ-��F���m@j�ncͩ�֋�"})=�u����9��*i��s����{�K޾��qL[q>,�Y�5�-UَZ.��>F��kaK���i��Non�p�x�u�������S�e�I\��;{��ﶻ��<z�l�����^��X+f-�3m��&�pd&k�s3)W*+�39sW��=g����8>�Ý	ݵ�����7F,k�2rޥ
�+l+e ����7k{G<�{�A�)W�붤���7o�O<{ϱl]ͿQ4J�����|��v��ӽ���8�Ŋ�Z�e���	�<���[��d�&M#����T�'��7I��N�I�=�s��ָ����ו��-< �h^����0s�v}�R�H�-X�'���>Z����c0�2T�6�p)1H�����Qm+4���cB�����}A>�}��[Kc��g9{/=|d����)EYn�k�"_W9n��?n���p=�.���+6��^����b��×��I�v��뤦�f!�X�%c}v)N��l6r�?�p�������ЖJ[f��q��ɓ5��׭:��OW$���t�1ٜ�3ӹ�8C]�u�e໱ʆ�Y�nqT�$�#������9[�zKUS�&�b�ңs�JuS���y���X��ɩ*J�-FF��:�
{S��G��$��-ie`���}�;ٱ�܋#�ܞlCc/#[��agZ�7}���t2m;� �9�-,[m]�YÁ��7�����Srs���>��jFč�����5��0mg�(vp�ܴ���������O��KU͂O��SGVP���5g�^/�JF���x�Gw����l����5Pe8;�OG7�����:�Uɉ^����i����F5r�i�i�C<ۚ|FՆ�fً�P#Uzw[�ܩ'�+gWgs����v1�Ҽփ�_1a�����>����E��t���J�U��J��+�ɇ=X�	�f�6���['s��WS�y�^F�'�������3�������gmP���&�]ʛ`v�;]i��A����3U�o0�4�F��qիlW*���mQY��t����
��LuYmc���f��U�ݒ�lnH_A��2���2J�nk�t4����U����RN_^)D����wL��38��/36��m��y�p�LÍ;aH�.!���8.ᾧ�2��ʗ-�J^,߲XK�S)�i��0zn����N��'�nM3)�ih����X=^��6P�,���j�٨��˧Ɩ�X'��3v��Y��l6��:Z�9;=��`�	:�4bF����r]<}+k�����5�������<r�|k����R��g�G��z�ξ�y��&�X�g��Ƴ�4���s��r�C��)��jfN<��{�9�[���b�Ж����i�k=h�Y�d�}��d����d؇2u�J$�jq);���CJ�5V|�LsxK+-��sbg7������֭��\
����X&��k��-�+9^�n����/zLK$ao04��%,x!�	�w6q(>��q��k�8iHp���gt�����-�~�
�{�S)���C^C�梦������_>3���.�9}%M����٫�{�^���͓�0K�K�9�j��U���<
d���3c�Ί�-��Gi�(��G�}���8��V��
�Sj��Ӛ�`��ˏcx��p��`��
H�R�r�L;�I�xo�]
���OaR�3G8r�]qKW6�!8੧�ڇr�)�G7l#��q�ᩡ\6ȫO.VuG��umJ�9��݊>Y��.�t�Ne�+[n�#�՚��a�;����T��Ul5}����Ҿ{��oC�>E��W��KC��M��f�PwAQB���{Kr�&���ݭ��F�P]��nqn��x"����6�r��Ζp�n�|�v_@����0֩��ɽf���(*%�V�P�ހPU���gU�k��]ׂm�O��B@���pR�s��8��X
�Nuk)�&-�w5"�m1��͙�(�c��y�˨p|`��d�ΔC����֎=���&z����F�|~��S�k�S_a��<�Sh͸�6u��gi��A]���0V3l�\+q'�˧[�k4��sr7���]#L�f�.���XŦ(n���6�OS�(ˮ�C�[y��;s����H�m�Z��΂1��޻��".J8-���H��q!���֚�u`�\�"t��S�#�GNv�C+��Ldo-q��ӭ$=5�=���[a�{�t�8`9p��e�y�:K��G��X��f�aJ0���0�Zc�����T��<p���;�AZM��<v�Ќ�{����C���E�t�y4Hn��Ii���6�<N#df�veaD������A�f8�f�tIҋ��wE��F�U�w*�gV�]�$�9*N؇a�0G9��Ys�����{���ܓ�7�WJ�!g=���B6��}L�;/��5h�w�c���8]�m��_qњS|tR��bH�6.87�ʦ�$e�1�Tm��j��G��zM�u(.U&*�㳹-�[���FV�y�V�6z���;5ƜZ�����wwq�])cxs��K�4��8�rЦ���Q<Nt�؀͸��z�u,n��rĠ��Cs����k�5ɽ����Iכ��z9�Mġ�,�y��d8�N��½*�`ڥ�|���ɞ���F�̄�)V��ţ#����[�u"�oo=[�s�{��ڬ`�|����ib�ۥ��@�எ�-�G9���s�[�"�|&|u�-!�N�}����m�Z����=.nS������6��E�z���WW���<�)�+z`L5��wKU���$�kr.�i;|�jm�xU��K�V�՚����x�E��f�ay)@=�� b�7q�����!hWy����6[�����ztl�{9Y|������ֹ�M�f�sn��EÓS6�9ǡ�+�����U㪒�\иb���O3&>�׶V���|Xé�#���skfh��q�7�E���9-�W��eZ��G��h�,NJ����S_e��3��Z�2�: n*��;(ft���*�<���h)UQcC�q��`��Qb�h")YV5�"1��QeeE��%��Q`�ܸ26ɉ1U�YTb�QQb1b���"��H��QQ4�Յ���V*!R��(�QQ�GMTa�j�EQ�,F"�Qb��Ԫ�*#b���������c1���b*�����D*KmQ�b�UQ`��SEVEUQ5d�(V0GM�����V,b,A��#,��T�i̱dUUU����s*�TAUAf1�b1b:B���"*i(����T�1U��1�PT�����*UEH�QCT��
�($��(��Q�f�����X�0Q[d�PQX1�Q������q*"�Y(��Պc*��Q���+Ri
������s�y�gJ�淲I'V��s�o7�.�"wV�����rĬ9���n��
��h��`���U�u ��LOꃨiF���޼�7�m�.)�mMx&�Ն�fي���,=6e�NWf-ֻkK���8+71��5��/ܵ�3����X��ۺ�2<b�;�3ܶ"�n�kF�fR�Z�ًo�m��&�y��kfY��nwy��Բ�M���TU�
���U8�`��l��iܘv֑���Â"�2��>�����9�й���/tJ��ȭ�c%�y��JX�3�RGBO�i,m��i۝;ͮ����E:���̷��
�)�"��}��;���]��1j�N�s�V�%�k��ͨƣ����K��|�n�AS:�b���a�ރ6�{��cY�m�nJ㘊�!.ͫ����k29Б��$ZQB�W��V�L%�A�����N�m��_t���!�������T�JQB�,6�h�P����ӒַC3�r�']e��qM@�G�;h!W��0n&a�wW��b�p�ط݆�꼩4-���D쐹t˭wW�AX	����,ه^��J�	�����I��E�����m����p�7)u�6��{u��p�<Q�ӆ)D˝�0�dL�N󲻹$�T+Q�ĪG$��JgL�w�<�DS���X7sTwzq���-5��ʇ�{����w"�
'�r�Z�@��Y�j;z$��S�p��LBKLu-\�j�	gC�Ӂ�AĄ5Z��%�H+8�o�����~�֜�z�4�(�SU�m�	j&]1Pv��Nw+�sǜ��(fD�symI���ǅ�1a��Y�(�ì�β���Xq*�J\��ة�B�5���so�^+��o�b�������ON����{N��Rk�zx�����a<��y��s�\��ޮ֑#��Xm��9|gMXdP=�`�5w:����{
�.�T�����w<�A%`뷞vz۵�����蠅�h�GF�yQ.���C��-���\�Os��c'���4�X����;s�{Cy�q�\�@�2xk�� ]��G%boӛ�ե�d����-�µ̊U[�Z's�tt+}���܉X�^��o���ͼ0�Z�s��r�[�4���ibCn!E�Q��ÜҮ7���f��DT1B/��2�#[����Y�����=���طOtR5;aKZ(Ӽ�o&�[�I�v�v��Ν\f�ݽ;4�BD�H��Ug���5HT��%+�i�m��-�Nq�K����˛�ij�);+��H����g���a�k��w�vY����k9k�+����>r�^z:'��AAN�(�X�ʛ��ܚ�;��e����z�s�	�e�+�N%R�(��0[�{g��۾k6�R*Ѯwħv!zq���YX�W��Vw��Ԏ.Zb�ͱӤ�겜gw=s��$f������9�d�v��6[� ^,��.�����=Y��N�J��iĎ�v���תo[�0m`��MV�&kx��[��j��%�ٛ]����0G(��hl�s^�د=������wr�z��攌$^�RHcq7E���P#UM=x+6�b�R�\�e��6��bYC��v��XBϫ��5����"�p�r:k8NPʳK[k)�X�;�sk��U��q�:b�2�J++����;Ϊ���4sЗK9�k̝��ɋ���D|;���f���R�w#F�B���MXWwN����W:��(��i�y�_[s^|F����̀�h�^̩K�����=���m���~^�1kw6���a������;o�f�5�C�出�>����.�Z��´F�M��xV��[xm��;�]�G�F�6���u`��l�� ^M�2rͿV��)VL�ƶ�[f�iܩ�y���vJ�<tՄnz���QZ�g:Nfk���J�i��J�Y�{%��t�}�DDp����˱^��-mv����ӽ���|b���N�,��K+�ҷCl�J�o��ԑ�I��7��-&�rq7'g�����:=ݱhpB�ٛ׳ϸu�����M��x�,޳�k9{-A�9F1Y�m�<��Z�1;p���D�q�R�-p�cU���XJ�~�65��mܶ�yYלT+�3HE���׵W���L5\ ��lѴK��J}�)��n#�l�{�lT��"+3�_#Z����z3�;@]@J�#}�RҔ����gi�+n�J'�q{�������.�+Lp�)����Ȯ���1U�)fV+uM�Rf�ɷȶ	ۺ2��-b7�ᇵ�\v�M<yՋ�M{��fY]ǲ������I�'��9;5��N�Y{�Hi]WT껇���9�-,�o"��f��ۭ��~�x�%z,bp( �BjG5t��kw}���\(N�K^��((�Pl�m\5o�:�-:��A��!ʦ������8��f�Y�UNf��gy�2ū7��{�S9��&���<MEM B�᫴��vl���v{_�f�3�����hņ��M��ٰ�T��j+��R5��-�\ːK7hN��ј��^;�wZ����Z�SE�V%-?�{2?	=����Ѫ�v���ŷ��;�m����=HU��U&���_-[Տv��x�r}���-�|�zr�b{�)>˻����{�Sǹ��D[��x���ˎ�3�4������l����TC�x���{p�78ε��%X:i<	�n�>s�{Ch�|`ؽ�E>�Bef���Õ��Z:�3� ��س�;m�����ռ�$Z�X��R�Ok��H�C�K�6;^�6�`��F��83�[���c��X3''x�G,�5�}I���s��Y0���'s����H=��LZ���ᇱR ���C��Y�vʓ����K[<��o�\��4��t�|�#��v�ժOImF������̬��y���,H'o�LB1�ZJ��oA�k9�W�f������oQ1�To$��1N0��@�ɦ&Ҋ��F��g<�H^�»BQKsN�iֶj5�wd��Y���9�A+N��ypÌ֦���'��jtowK]+)ޓ~O�^��c�	/i"CJg���;=[�0ʜ���,^�����L[K+ �U��8���Ȱ��9`W����>ts%�H��0)u�qw�:�{�x��2�<��N ��& �r��vΓ��ckx�U�O�[�q�k�K⚸h[����ٻ8��l�f�J5Ц�C�1+V�Vm{�ε|8�x�b����h�S�8�9��7<��=Ha�����+��X�Vm{1m�׊�w[j�О�yX���1�ֶ�-��@�n�<��\�n�jnS����ү�c���wh.���M0#��Vm��ټĭ���=SLwxmR�ђ;{���䙜�#� �K���-ݗ��S]�V��t�g;��qrB:�e�`���wiD?o)�Y����������v�
�^�Z�q����!�����5(������@���Y���:j�Y�����κ؇L�x<�yh�2�"�Zޮ8����aX�V�+=a�[��:�~�w�ը��ǯ�x+X�{��R��#X��X+h���,�i��:k��q�5���8w��o������v��4��%�i�O9�x�"�x����(wJ���Xᮢك�`�	��!�����oA�hFeQ9��}�i�;�Z���jO-x���LP��:�Ҋ�U�N)�Y�y|Y�:�;ʘ牖^�޳�����'�Jߪ��8Н}����G_(��,�c#T��&K/�k76�I^�����1���3�;�yp���[^���W�{�iee�V�X9��'R7��ɍ�Dd�η���׶q��Q�D1�����,x�w�`��,y�Q���X���Tz�YE�-ƺ��]Xڔ��f'���M��,�h�U���v⏯b�˾z��U��]�9�̖��/>l�I�K0�� ��ssYd)�d��k	î�,4mX��s�ґ�z����oib�[W�yf�^
����s���*����Q !��v���S��n�6�r�ejZɛ�Pٱ��8jNRU8�&(Ny�rB�w4���������%K�>��rշ�}�t��i�LR�n*�C[��j&H,ʔ�Ǘ�Ɲ�cqe�d+��=�Oq2ŕ��ܭ</�����m[w�l����P͍#pc�N�q�ڏLv��ڃ��𘴭��M�S��뻞�=�Ou�Ն�,��X^��Y�E��v	�հ��<��7�������;��qK��s<u^�G(���r����X��S�M�ɤo+l�6�d�n��	y@bQ�%��fr~���iz�&U*��z�+�g!��֪4�"���[F�k�Nf���iߜ��������z���!s��F�W�:�,�5��=b�[��h��;�Ñ�a�x�3������)��딐z�wA^+r���x#I�V�Վ�8�<��']���;Mos��'.�FV�׽�t�Ȃ�H�vo-�ZM�M�t{\�Um]6�g+pU�t�0G^�1Vw9���KO^R<�jxm��3M`�-Zi�t��9;��`��u:�9on�Uڎ�=��Z'�N�2y��Q�`&��^��&���kM�f�3y�ڤE�#���J*�W�ƫ���&����lk93i ��q�+�x�9�q��>�%�F���\4�5��.��59�9��4!,��#pńx��Ww|�Wꮠ'U�>V4�7omN"�x���Y�Z�9L^�bV����N
15#��(��gv�s�c�\�қE,�`i�o7gW~�q�6'|ӊ�Aġ�'�8l�E����χ?R��iw�
�(���:M|!��EI	�ZɻY,��8�[����տskH��+N�^��D��AD^�'Y*ɍz$F� i��m���k��60^���^Vb��j����������pyTü*�T�t��c�s�w�t�vh�{�ù�4�#ݻ/,)��c����x{�ཿ���{��mp����[K	閜��z�R]�OI�dW[J�<1λ���D�"��*�mNoH-Yr����:��;�v5gy�9��9M�}ڒ-NZ��7�N�N�����瞻W����mEȇ*f�س�a\����T{��X���m�?*]��x�,�l����k+�T��af��`X�l;]��X���f��q�4T����>S*�*���]�k����$2�m��i�s�{|�A{�������5	v���/L�\����r�ilJo��&���)I�.����T��ܫ0��e���H®�
�h[J��oL�Y�Z����զ�o���{���D!�9��!>LPڼ(́��;[46��ÇkZ3��9m���:$��	�RL_5���(1���n�=�RS���f�l���roؕͥ>^�BCJ�U�DgNtq��5�R��k��N�v�iee�I��'��܋�ˆr�-��;ו.���7��J#2�@���bX�����b��mC��(Qe��n������W[l�6�s��ݮ�\�)����e-gm���.��wkOQ�
&TNQ�env
�u����fd(��:�z��\��L�ń�D�;̐�5y�i���xjwj���Tqd�T�ޒ����M��-���)��!k�ݎ9���%]`�h���o���E����إ!f�Y���:\����A�b��M]�6��QU��7�Ǟ��̂N�"�<w9��U_-R�21r� ��ʙ�S!YU��s���a8\��Y��gD*ܛD�4�L;�Y���
h�{-��Y]��f���iAu#��h�xӚ��|����Δ̊u"�]f�R����;�Ekt{��ٚ��r[{�eq�*��X��+�{Bq,����t�GGJ:�Ф��<[�؃�M��k[Y�k�Wk{t�������x�ң��PW���Y��v��R�$��Ն��"q9��G���*5zfR"�-�F��46��jm�@/�YsKrqr�Xz���<2s�;K�rU0f�6�9{����j5�9t����fhl�����:�;2�l�lC4��<�����b�i���}g0�M({��՚�w)�N�+�7;�\�jj=�b���C�c���O2>��z���&������.����oc"u �^7Ms����q��U�WN��ml�Py�pY	k���=EXj�t��ĴJ�f�t�
�}�W%��y�4�J;��Q���%��t���]v8ԭW��;�9�����9V)�:٧������+����↺����Ǳw�,��τ���i
�t�;9�ݳ�Wn���T��<�p
t~m��h^).*��[�����;W׼�Cs3�h��c6�E}�ŵx�\��؃ۼ+�`�C�Sf��2�?��S���S<��m��z4 ���o;}
s1�t�ocd�]��o1�'�`WΦύ�)8Ӝ	Ꜳ�y�����;1���K���kx���ٶv��a.�9P��aZ剱��@���4H�`�̫��eY1I�PvR�\{�`��y�]��Ő5�yG!M�C3��jhF����z��ŝ0ؒ����v$l֕�bʦ��*��!���}�NV۳�q�-��F�Wv��Pμ�ap4}�L!h�9���S�-B�{aq��-�$��[.��u7D�����]E>k3O�4պ�B��+�{O|���B�V�<�����)t��"�U��kzN��Pw]��iHw ]yC�#R
� �I<����-�t��!�Q�b��7O:43�Ő�6/���x�ۗ�ͯ/Z����s'8aB�s4��wJ�j�_*�wK�"2s��-B�K�Y;��{
U[��t�\K�TvУǯ�����3:d�/L���Ӽ�}����>'�AG�U�	�E	���PY�Y%A@YQYEU"�����\B�*�U�QTEX���X",�QX����`�cZAEH��(� �(�H�j��-��UV*1J�*�(��-�ĊA�@UW�Av�)Ձc�1�T*���U�i!ueA�L���[Q�
�d��DU�j�F(�X�A��#"�F*�ز,QbŊ*1ݕET�V1EEUF.�V
�b"!�����Ү�AvʃF���������������"�f0��`��#Q�"*���dQq��E4�J#X"1Te�b��E��ZV*����+�ov�+-Q-��**�F�kR[DEb�(��UҢ���`��b*��]3҂�\f�����cUa���N��;t��8�l��w����	�q(Vbz:�e�
]�w�4�0�i9 r�����8��F�,��:�_֝����Գ�x�����X�	i�����W�;t�Jɵ�oR60��5�k|`��L6s���u{^��/�v�J���/nw�ZڊHᮦ���l�ۚ�د��u�3z�t>*��֝��/n[p�����Ж
֟��un���N�n�'*����b�|{ZH����3͹|r�7{,�O<0]��!��pnn�t�s����'vHO�!i��Y�����h�t�fe�hZ��~��NL?3{��6�g��W�F�<�,��uSѤ�1*)����++{"���¿�6�v؝�\�w4�X;y�j�zw��T,.g�9q�h�Ҧ�&,U��t')���`d�~-,4�&��v�֓���[��O>ܚ`�{���q�l�t&P�|�$�m��d*μy��^���\*r����H(ގ}ۆ��갸��}����y]Fu�T;=}�/*�u�O"�J(@�\����Qت��X[�H1�NB��ӾV��W+�}Ǹ^G����pM�VM�j��������{H��u�{2��'A!ȍ�>�/����D2�W%��h��)c����(� z�h�!��C��&m�ٮ\���%���u>x�k1��ŀ9{/=2PF�e�/{z�G���%ų����FۢJ�衏�m�r�\­��Ef���u\t���8��ns]��Ж�]��O��϶��q��C���ٰ��j�G��G�S���w�@Mmt�^��|��6�K2�wZ�|՚tR�j�u�w�k�׈ι͊E���Lu�޾������s[F�j�);sbi�s`�G�9AH���8���8��|���9;Y�qK�'I��<�&���!U�M=�B{�z����o�]���-)���y�����4dmXn�m��u�Nx�S�y\y�Kiz ��NVmfe���u�|�	*[]��l��,�IM����#�Rrn%��b$!uhU�i
����
�I��1%�l���ʼu���2�����>zwRǹӌ���S!\{����޸E�әND�W=���?�:��Od�0���L��<��c�=�ȁk�ז�8���F�v�;�'[��O��B##�)�	ƞ="ȧb���QRf�;��Q��=܂��<R/V[Uk��Sx_�7]��U�{׵W�)�)C�79m�D�����4�>�&{�o���Ϲo?-|W-�Λ��A���N�y�B��WuQu���;.sd�-I	�X��>s���iX��z��k��2��
���M�[���Y8Q\�˧�RޚO<9�VNܜX��y��V#����J�UǧXN-��=�V0�|�1j��6�ǎrU��N{����[�Ŏt$hF�;J0Yj��ƪ��HM.�A���B�\��cz
�Ua�c�]����	`�N��B�-�P�aޓ�IlDgj�x,���㾖W5��f�cQٱ�\��{�ə��؇�9��/u+�7��+�4�ש���U�{�����R
%4$s�
n1��� ��'�� �ͼ��;:j�<��,����)\	��i9�3�����%�]�x3�"�{Y�ճK������E¶�t3ox�o'.W�f��U�;���z�Ň��D`��2��p�	�D�ހ�B�;��t��ZE9��jU�alH�%o�GW,)m��$��c�g�;8���q�6%�	�e��J��Aq�˻Y�9�ײ��z�a��I߷�QL�N�BۋZ���V�T�xj�I��3̹"��h��ͬjh^vU�6ˉ`��K#6P��KJ���%�f���MP#]zq���Ŷ3^+��o� 2��`IG�j�{��ћ��Mc�-Ӓ�ӻk9�Yc:�!��E�m��m�z7OrKPǧ�oy������5�\6F�U8�g�i�^�EpN��*�5�Y$v��c�]��[k{f�X{�^"��U�T]*��:�x޹�p�-S��[N�z�r���4�ݼ��Ν����y;�α
x�����n��ޡb�J�sμ.O_��K�S\�&��:�NQʽ��������Qi)�S�>��BF.�TE	f��`i�ރ6�{��6Úi�e��E����t���S��÷��V3"�ʵ�n�V��v�uȘ�Y��a�N��mM�agesq4N��o�m�u!Eݵ�1l�ح���K U�37A"�1;1�;��{�E��X��%�)���3�vr��;�h>��.�t�����0>�HH�b�]���-p����5X�JY�X�	sPN����6>2

�2�I1D �4h-��Kr�����\��d�}
���J��R�А�N��0n�E���3��q�e��c;tҺ^���=��f�;�h$TF�=q��ri��Tww=R#��g;��^���:5�E�^��圶�ȇ��9]����Z����T'��U�x^�~`���j�	�I*�qw��fg���}J�Yx8��^����hOy9�]x8�u������f�[|��椌$��I�5�a��Dϸa���Vnb�WS��;���X�G�[	�x}lcni�ڰ��;��4f4K|�&^��u3M!�Q�g]��ʹs��y�|����YZ~�v2����^hez�gT��4_e�C�vl��/	��;X���ymk�s��;͛C�-�e��yՉ�+6h���RƑqt���C���D,�Ʊ�=�%M���ձX3u;�^��[=t�����w,�;[���R�v���ydټ'�e�M�:S�O���5��؜Uem�6�`�+�m�G���ÞuRӣE�@����s���|��%<ju��[U�}pA�4��I�j����V�k��uWѷJ���QZ��t���dB���WQ�2Y���ΚN�^3�o8v{�erFw,kԷ�x(�$z�6b���!��W�N����gK�%�-I䛖��ū	��Ζ�N�F8W�h�Bd���v"�{�l�(�%�YU����^�c�6q8y,��a8��QȠ�RX�k�D��:��*(Yw�z��t��E�v>�iT����B�"L�d�}"����+�<��$
D��|����xL�GZr:rS�T_Ts�$���`�@�p2}�kk��]��zc���ǆ����5gi�1�W6��x��F'�� Fu	̇����mLy�d\D�:�+JIunE��.����N=�q���]�n%��jA�+�T�kw؍8�Ɣ�Z���8�m6M�\2m�)pY��f�:m�n:��*I�ĩ�g	���GY��mh����˭�O�u&����kz�*��:�_��b��I��o;��ǒPQz���6�Ĵ�6&�w6B�#�v	;J]ͪ:D��$���\e�X����%i�qT���M���U\5i[��C�7 �����P~��>�c4�w�q�˖����n�Y��^Y{.&ݝ�=��hf1;�������续��J���52�V-y�2ޮRJ\f�.
F�U9��կ1f�6���4�^VQ~o����潍�����[s��E�Ň�/>T�{�>��{8=������ܼ7ۚy$m�޷��[|��Λ��A�"�;M�J����7Of8�۾�|�p�kwn��M&�h:N��{{CH����>#]՞0�P����f�gm6N�-S��S�riitJhs�&��k���`iFZC�^+�Y�|_H���,$c-%�� s���X�96�Ж �z:DHʡ��+s��q���G��z��NɟA˪�F��/��ɝ��΁
�1�f���
��ಬv�U4��]�̄N��iA��&'��Vب-��c��A��G5�W}i �u���E�B��q���j)i�KQu�bG;��޾�T�.�3.���_�X�`��M)����u��5W������j7�.�}r���@ř�폚���Kú��I<������IYN������ĮE�)��H�ɰ*�����t���N�s2��-e��<���ʹ{����!���bdGri�Uc0F�<�s��8�Lu����M]�,��!�	�ӄbۺu�NH�+S�]g^�&��PS}�����#�S8�з�pM�j��ά�(�]ř�Sc��i���om�7����Sמ����h� ��!�VtM7� ��[�>�-=oE�U�G)�uʿWJ̞��?7q�{����.��PeTZ��b�(ptF�̥�����,q
��qL��b�T�g�_�}~}go��k�Ƽ�B���c�2k(��P�l��/f{���n�����$��J���&V2�G����+�������S�;�x%Y�%�#��x��&Y�f����T���1Hx���hL��s��]�L7�̽A:}Ԥ郫b�vjP����V��`=w�l�%����m�K��Ve��}��vz�[�f�[N�b���r���fik͵(�:�U�|6O{'��,i,m�t�s�{C}��/�/�RO��ux�{&00>a]+�4��
i�����v�&�2�B��(0v�����$���0�t��bhvԌ}uDP�m��M������2*a�P���ӹm���0�׎N��&+�����c-��#�A= �UJ�kg	h�1�X�K��u��6�^GD��PY2����ɥ��xQ;ZO�T��]�l���U<��q��
p�G:Y�];�yh��U��*�Giζ������	�{چ���SQg-?+�{{�D�B]5�+:�VC�΍k=ȼZ-��%�̠b^�Dܵ��(�zJܫ�Z�Q
%U=�C�S׭�`������[�y]b�7n	�"�-Mm:hu6�1]w�ea�8��H/7�K'�*I.D弮��f��̯Sv�X�Aw�W[�{�� jh�ɼa�����z����v)�Hn���p�ېP�i�"����/J.���h)���eu^�u���Ǫ��ۍ�ș�t���NE���5��Ep1�LK�ޭ�[sV{�E��Wճ��zy�I�i�V�,�J&�B1RDp���M��6W=���w=R�.Q����J�U�����������m�ͳ5���t����[��:��Kc�����gf,ћe�Js�-7���v�>�d'��fY�*�L3��u�����Re��[9^C�ڂ����z۵���E�7h����)]T�Ȓ++*�v�V�[�n�K�nfNEσ�aY��O��)��{�^t���,\�*��7=&���'���j��ꂳvo�k5c��Ł�v��	�ك`�y2�K坔&!ʕ�}��u���O��4��W��Y�K^9;%C��;=�/�|��9����l�׾�B�#z^����Sty���o��_���$ I?���$�p���$�HB���$�܄��$��$�	'��$�܄��$���@�$�	!I��$�	'��$ I9H@�RB��H@�XB����$����$��$�	'��$ I?�	!I�	!I���e5�;�^�(���!�?���}�����9(P��P 
)� ����PIE(*-�  �;%J(��m!(�Smk�J @�DT
��R���!"%���R�"$���R���kKZi��`�bP��F�i���jP��
��JUK��(��Fl��EUhԨ�@�� �Bi@ B�0��lңaZ-�l�m���fW;�  @  "  ��R�T� v�jH&F�J�(� Rl�QZU�UT8 8�ѥ���PD�����D�����$�Pi� p�P�fdH�[b��f�i�B���)�Y�A�*T �f֨���I�Q [aUR�P�X0�8 6���
����% "V���1 Fh UH*�UC�� �@D ! 	�  � eULHPT�. 3:� P E��$� �j�+F�6 8�I@��1�ʕ*mA4F���� M1��JR��dM@�@ѣ@��)�Ɉ�zOE6�5 z�� dP�T� J�Q� �FF�41i��101��&$�DD&hLF�I�	4h(�G���_�ӯ�z�s��9y�ۛ�<�7�5�II!6o��D��$�$��O�$�RB�!�HBI!2C���JII	�F�?���gEb� HD�s�!$�儰C�Y�II!8C������osQ�/����$I�ƹ.n�������Z��~���u��Q����3��u����Ϛ�[��z��v��.ΚX�B�h�P��KU���H�ubμ0]۬ȶ�Вi�H����kX�@�emEQ�F$�+��Y�������ԓ�ݪ-.Ki:��֑}݁�WE�oM$h-&��n+�$���yDERm����2�]!����3SZV5E��:��բfE/����OS�K�۾��ص�MMr�I.MCk[�{J��[�m,gLC7�J�[�C(�S�Y��R�t�kZ�܆���[���jU6L��l<AmHu�/n��j��$�R���s��I9�1�E�\ؾ������!-�j�m�9h���5R��2��� �{�L�����#T�m��~G%��-�h+�3&��-�(��+�b����^m-�U{fɵ���FZYUV	۪2(nR�ͳ}��7I���@���խ�Ǘ�H;�>�w�I��]KE�p�x˕-�yl�{�]�X�)=��Ǉ]K�N��<���v�F�㱋-gZDe�ޕ�{[�4�KH�PO!K�:��0ݩ�v����H8�:���Y��;yr��u�r�%#�wv��2h��dKc�4ԡ-V={�+���u�Ͷ�B��k�c+�h���dh�FUh}���q	w�Cc��-��ch�*���Kɹn�;����k��P��I�C6���'���hwl�C R�wY��V�@�h2���׷u7w�T�SU_�J"�u*��^�$��gp�D�������7�A��ܺ��OnA�����v9,`D�F��Z����6��܍]���2�HB��j[wy,���]�2���)��-A.�-��i�F��l؄,��uR�\��^��l^��]P�C��ŷ�,y.[w�������D#u-:��ј�c7sl4�ܛR��v��{eE x�k���+vSK�<3,J��$�>�Il�o��yt���'��7hP�E�/�_#��I�� ��Z��7��֪d�wK1*�d�p�屢y�2\N|kA���
n���)�a������ �7W�$�W�uT���ݱ�n�	7��NGv����O)�n���ie�Q��+3,9v"Z�%��xC��۬m}=��r��F����6M���C0#cv�0�m�e�f�V�kyq'���zP�і&���njL��6���s6�n�#%�\����%�����1�{e�/|;���E��u@^����K�FP�6^���?H.J{tU^�b�NSNeb�)�p\��To/Y�Vb���B�AYg.��i�b�������e�55��'\�a���.Q�P��7^f�V�&��Sv�L���7zl
��n�!�n�X����\��^W2�*ݓFM9G�z�d�|��[c��X��X{ÀL5هu��T;�N]�N�B�rJ�+E�j�հm���2d� ��v���u�Q�e,���&��2���ut@����Ս�C/p�� C����!(O�[���6��)��.ֻJ�8#N��d:�od�N�v4��I�5G{���ݙ�m�6fзW�����^���V�
&�.�ۆ��ۙ�(���iU��1�m�S	�9�.�*�{aj�^�`��6�]/�ج&U�g�<x��z��rл#{u��3���$�^��d�l����xP�hpI�� {oAZz��[x��,��!nTxΜل�X0�H����sUe�p��h����I��]����,�l1U���f}y�v�h�vf���0��-b����Ȝ_+6h^�ݜ�4s�ýzc<����5�7�u��e��f����c6�C	��m;6j�:��H)���g(�m:G�Y&mZ��{xlOZ����<#�{6�c��\8'v3������af-,�8N��9S29i'Y-e���H�9������3v���a�h֧����2U�m�+�*:��H[���7F�MX�f:K�*ꥫ�.��RjW*݌�"�J�anJ�Oe��W�0�*�ıPv�)>I�]�k�Y�<����5����ټ�Le�yB���Z([̚��()	�a7uZi�%cô��e�P�zƛ��8��/�ݵ�5i�EZ�f�"�zt�����s�x��z�nnl�u@䬖ȧ�ᵹAQ���$��,�j�+V,����	��\�7.���)��AJ�H˶�ְ�&�D��A̒�i8a�vi�/���t9�2��s/���ScU^�0V�qY�	*ܡZ��Dfb�@�f�Mރ��z�m>'qp˽i(��S`����qfe�V���U��ۗ#N��m^��0�EZH�Q#F۸�<�Iv2�/h<Zs*kc t2�{��R��a�QZޣ��BHZ3,�E��C(�n�ٺ���g���j�W0.�*���5���G�hsV��@m��[���q^�����1j�_�1C�f��i�KT�;[gF6+��-;E��T��Ռ�!.l�.nL�Ǉ�������3���+Ař�0fZ8$/%�WV���²�C��*�ꗩ� "�k��=-M',
w��;�F֡m�if
�բ�
$v]����/7N�?X��X#q6p�"j�%��o6c1^�x/�[����R�x�̹2�]��SBX[��Q���v���CM��<Hx�b��#����-��,�`��7�U^�PYw"n�����(3�.�+%���m����[��MU+>�or�w��HB��^Ԑƍ�8D���-��-�1$�������RjIdA�n��ܹ�\N$�ʛ�*b:.��m���yJfK�!��5�Y��U�d����j���ޡB�^V�(���mP'7O�3�uN�cp��'�U��]���W�j���Sb�m$��4R��Dڤܗ%Cf&���51���H�w�GUj]�P)��_cw����PWhJY�ʹY��T6F����
:��N�&l�5oE�K7K�%�N���Ihm,v�
D�.�os�k��e�v6qq�<�`|rh</�9���U��`��h���P굢�l*�UN��7��]�a��t�0VȪ�Wj`lS�rUV�'-16�]�X���"�5�7Z7,=�L�������R"[�K��o�ЪuL����Z&\��#w��a5�E�_E�
&f�%�1:����ֶ�����\�v�tA��^�tr�1t���_'��g�~p��oFĉ�3�Dui����PT��B��~����<�.�e��ef>�C�T`�nV�}!9�*Kq�����=���S&V�{����/c3S[דoY��7����H�:H�x������N�-���d�;�B�=b�q}�Blz�K�U$����22*�!CSV.%��0�ک97�G�NY|j3��ܓhaf�"6�3 ���N�4QՊf�89|�V���37�,.!����TS�cgG>�ٹw���&����V�}c:��HiHˑ��ٗX��yAbi9xX��7��c~߻�h�_���j]�#$7\ݍ���*VL�V��/'\��VC�^��#Θ@N�ɼź�!򭚰M�g%��k,ntv�ɳyN���W��K)"���-�^����& ٕ�����X�U�)�϶k�n
�i�麥���� 5 wp���nԾ�;ZlX�U���N�o@�+`�w�S5�Լ�y��1���i��l���m��$�I�E��TC-v��Q�| 
�6���[t�1��J�U�z�Ǖul�Pu��$��J�!�y1+��v��6���ّ^;4��\�*�n�ݝoX�Y6�<.��쬭yl�5����?kH�aUm��.�G�Bq�'Wc#��S�{6q�[8ի!给�Fz�&' �ȕ'F�#%�r�����w)�| �|����<���GΙ,vY�X�Tn�N"�6i���.��*+�]��Ɨ�Ӫ%AcF�f�<��yf}գ�f�X�
�e"H� �b��bK��/I2|*f�4��5]th�@4!+?E��ΐ#����֢��jT5���h���J忩r�5D��/:�kݨ�H;r"����Ϳ�3��*���ʴe-\�X#�óa9g@$���kV��r[�0)�v��)Km��ŁU�[G�a��k�L�Lx& &d�¯��)����;s��]��P�*�^���D':j3�{�G[��-����h�5�t��.4������CO�4w$C�Ѷ)�j� k���rГz{7d	]f&6����\�Xs]�ALkF�+�S�1+����wSF�H<�(ov��[WVR���Hu�� e�\t"G�#.f�w�NS,Jq:�y�u-6���צꉡB�G��=%�4��xk�[�����d����^��t��3�˳�C���B,>�wuxl�ϒ�=�35sy`̃om�w\�bh�JU���@�Z�z��#���Bнu��í��E�p�v�U�a��]��ML�����-]�o���:yY7Y9��yˢS��o.�l�!��&�0���ڊwnV\Uܝ���)�4(�0V�.��u����-�z���u�.т�h��`�����;��[#p���s2�s3��7�����Z��p�ւQ���]��amMf*}�:*���֫�>��_m��fi�Y�ٸ�#;*C7os��t��w�b�h7q�9���*1�O��l;XZ$u�Ϻj���B�C8�N�y唝#a���]�{�˄�k[�+�RѨ�.p>����޸�ʩ����C���i$:[tV���͎�+(��WdU�0�,�����F��5=�&��VcP[�GP�T�V���c7���Pe��Aɢzǁ����0α��Y���I ����#���bhȡν�+�Om�F���)�̧�ct�u���������5ݻ�ֶ�R[ζ+竩p�y�j@�&��]��
�LJO#��匥i�ugN��e�ʩ��b�0=���jk7�ۦ/J�ݮn�vu�����7aA��hj�`��Ř�a�2���_9��6�ҫ[��W���謱E��=�G�ʽ]�33��yLmp�2�=�HZ*��EZ?g=�\��=�Jc���}����b3��du�5�'HE1�5����V��a�³PP�tlpU��U�-���)R�:��S_u�kn�-�
�q����Bl��>Ȳ�L�67�� �j��y��l]���¨�Fq�ٻoֹW���Si�n�K��춳c��=��l37�"6�벋�l�2(Rv�Oa�݇jk$�qV�N.ڵݣ�V�l�\��.,����on��̚P�%�wPkG��w��rm�h��&�Lt��H#�Э�������W
+T��9�����B�pyO��9��f7���2�8�
�s����LӍ���{��F���1�)��j7A}Wh��Gچ��X(�+;P�W�71I/}&����_#����=-t
��ٗ�_]%�2��0�%<m>Z�dԳ��n�^�����&*�VPEl�y�/�M��:���Cbٌib��:��n�`z��©�D=�G��:t�>�vNȝީ�xoSX3V�Cfk��}��>��u�+ca��X r���R�\&���UٳtwU���R����Lꕮ�2n뉻�^�.�����Vt��<ߡ�������+�ˡ������"��dw�o8j>�N��IF��8�^��٢��[�ӓ�p��*vŽ�H��C�e+�3����u�GA1b�M�C|��e���$2���`�"�Ԋʁ�u׹�b�f�X��c��w���vg;����L���#!\���q_4�A�B�NT3���$�+L0�3����l�D�\0�/�hn
q�\�<U̐yυ����fq�"��$ֺ3���&�S��o;�$�2���nI�DQ�ǓEM�d���RHԎf䀱Йټz{������$*�J���M��h�M�,�0�]�qc1>�9S�Yq���7%\���<�p�c�k۰w=��U��,ts��φ"5 E:D��t8Vq���Y��V�Mt�ژ�3j�C�3c��nڒH�RI#�I;�M�n�l���f��G��:�m�m�dlׂ�˓1$:��K��!�@�-�=��jº�h��n�J;�Үh�R�Df��:[u�V��^�NԽ�)vt�O\y����>��$*,�u*+ڔOgqް���jn�s,��K��ֻ�4��Y�bۆ.�����O"l�L9Fl�V�W.�%	�8 =oh�b)nԐS��x�Qٔ.���fM,��J��pի�z����X�_�����I�9۶@���Vu1��DF*k���������>�H�X�O��Y�̼���Gӏ�����w���}�A��?�g���� �$�� �o<� �|8�! �������$����������U�����~c@Ȼ�.m��p���Q������uw��[�g[74���0���[zs8�=Me!��;��i�n���z�R�T�˨�2�E�0�D객fK�|q��T��q�� ��曆gƍ�Pi�#��7��<��_]�^��c�t�˕T1DT����&�Y�Ah�Ҏ޽��Mڮ׸*���⌙:4��c}���C��l�7mS��>�ؾ*��EԲ�����"E���h�כLU8l׼�*�ǀ��9	�Qٳ.��Ȟ�֌���::5�qI݅p>��ABv�2^�b&�#;�����gK��6��e�cg1����R�滾8	�E�U��oh7�`w6݊�<���F��9�5Y�����f�J�Y�yȎ	�%I�#Wlm�3�&�b���gCй�Pis�;�#��̰1]8s�`��t������!'H�v8f˙�k��>��5�;�����;�8'fоpۉ��Ϝ-�D̵�
�jl�f�C*�0���REQ��,�s�2V�fL�[`c��3*J`ݝ��i�M�/.w=oiD1,V��5��&��'W�Y���ڪ�˶�7:��V����x5�K��Lg8��X:+yV�9J�a	J�wcc
�ə:����D�Q���r��B�l7�ct���7����xm}0*sz�.�p���t�v�kJmea�2�Q�>�&������Cl�-���7�m�xA.�B���R���i��ؼ��^[�eI�Z�R��]QC��v�ZfZ��7��L8�N��KF8�^Wgcu4w������T݉�� /v4f���{;ck�<pU�)Y���Mqt�q����9�O�uΔW8�lk_`�=yXc��eu魧�c<3L3���ٱ��+�,/e+���V7,h��ތ�S�6��J]F�Ņcu��˜�$%�uw�On8�d��%�	�ݘr��{Uv���!���w��I]`Gf�N���4Z�n�	���\ �Lw5�q��9mm���.ʇ�X�[�qu��6��ҺʟAG�b�U�Qކ�d�3 7��m�7Ś��.\w��T;K�eCm.O��1֌$S��%�[�u*C�qP�km��aO��Hۼ���Vo���2v�+���3�{��7T�wnC*`t��Xgn���a��֡���V�iR���C�4yB&_�ڗ�ܛ�oB�"�z�����R��Oj�m�u��.�שrF:�'YcO<cv���U�^Լ+�I�	�p.�n�7.���]����ݝ�����Ƃ�jd�|sk;���J�;�2�p�ol����2����f�V��O��ue?�K�Մգ�R��-�Ki�*��m��;�|�}P�p]���r3u�y���s
�J��w�� �-d�WѱHL��6Y��O��LV�Y�����KT�8��.�Ɲ�cB\�e���N�,h��L��\��	������V�+�;��Q[A�ȍ卻ك	�!�c)4�I<-�wI��sݷܦ�K�Y�Wr0��)����8��它�q��a��WV�^��\��sq,[�lv#g�)0�v
��U��Q�����Ӷ:�J��%������#c�5����O��c������r�@��n�*)�¯)�睡���j`��C�����w�! �˯~U�I&<OU��ig�S���5�
T��ڡ҇x�����;D	C��uʈ��3��*�A�Ew>4X�(^�]m���$�J�.���d&u�R42�p%P����v�u+].�W�N�p��l���X�&������oV=���6����������o3��3� �	!$޵Br��nȽ0H�<,Q�K:����StB57up�oU�N�]�����z��K�Z����兵fM�uwi�WJJ2�zh^Q�X�u�W<
�X]��i��o-�ݹx�c(����a��f�\������m�S')y[�;�Y� �i�b)�`h�Y:�B�f��=|���� �pԂ��r���j��4�]CY72�,�Y���Ϡ�ճ�ts:k0���զ����%j�E۪Z7-n���Eĸ�{k���}��/L��_l��pJ��G`�**��t��A�5�:۾�3Od�P�$�uƴ)��l�2���ê���Mݎ�"<��d��Jk�I���c�����pa���+yv��P����:��Z�z�L��"������E�86�/oR�D�n��~YJ�D�v��R�T���Q]���ޫ��$re�}�vr>թX�q����;V��XmUa}����v�xҐ�`Ła��0��W��/*���ǻ��,m���FMk�8pҀ����X�uK�7GA2��1xӋQ�L�YZ�0�d�Ar7F�n�ǡ)Z�N�s���4�7�%YUǵ!؜��eˌ�W����'�<�0��ۤ�U(������6�^��ז9����b��Ś��.��(�Kf��ꔩAĈ:����B̻�@��J��SY�7�]Rp[iS�����S0�#f���O�7����]��Q�u�B��P%Y���:�_mH�:���e�YԳw�]n��3h\�rz{S�z���𬷇��K�Wtޟ�a�s�±�V��8?�� 5B�s��Rc���i�W͝A�twN��{U�:�s34�fB2�e��C(�F�"��9�L@EO��<8�᷹��2�@㸘̴�˚.PJ��p�j��e[�+x�0 �ʽ�3Kt�+�#XxŴ4��d�v��+1��طGH:ܣ*0���V 叮�-gM �d�?=��gJ[��Z��;����r�"�`�Fr�ɩn���V�L���_n-чln�u�w��o�ǧb�)��4�ݜu�͍�H<	[��=��%��e	�<�
ح�92��U�;��2�Tj���e�+QSt���)�p3�^cݶB�_r���H��r�-����4�����X��&�snj����~�
v��\�1#�c]�o-�n,�RxbM�W���V�*�.X�^�yjȏ#+��EL���G4�/(<ʻesUpL#�q7���uW�����B�n�8�Ul���	e+cnл%�kSU�y��^�?1�Q��<�L<��PsL.n�r�ĊB�Wۚl��d����S���]ӛ).b�����H�H��@�q�y�	���~/�U#�򏂝����P�q��h
mkk��[@���na���CJ��N��YJ��v�0�sF�n]�̝q�u�5���n��w��rx|lj��x�7^	�ݏ��F_uh�wiE(��P�$�[U)��֩��,G:v	��o� BY�o,k��}�˅J2ڗPt�f�d.��S��4U�5��(���)�ֳ��V0%�ZX�H�wu�| T�]�W�K��}�ЮB�F+&��ةZ��s�,�y��v kF�p��a]+(��I!}:4s��r��}�'.f���əZG}��e!-k��,�����aZ5�ε�V]'l����aZ�2�&S2�����\-���֊�j����-r--�+M�B��Zڢ�X�Z��̦*e�9q1�Z��1˘dK�b�� �������qV)�f�DE-�J�Z�
ef[r�Pk(����eQB�Z��wLL]fAG%22�5���̢�n�FҬ��X,���b���!���.*K�Z��+�ɄD1m��k��5���TS����U��4X x����}��[�/o	ƶ��퓰ޅA&+&A�J76����]|O�6�F��f����f<bnOղ2���e�H+��#�~|g�y@5x�dfz�rro�'OU��jԿLw\1�5�9�ck��&ul|���I� �$�j�D^wN�˅->���Y���x��p�s�n��8��0�\�=���ʶ�� ����G�o�&;gx�kd��������&����S���X>��l�|i��l�9��Z��q���u�i9��?��*&�*�(;�ݘ7Q�YG�ڑ�HL������]�~�����d�WZ����P}�5(�4��zW�4�u��o��=Ҷ���9����fpg���^[��sf������7tx�9�T����og��wo�W0��9���yx\!�a�5p�fv��p��J{���-�(��ͼo/2�j3)g�Š�'bP���������`o�+4���^c�A�f��Bܸ5y�,�)�o���"L�����Maʪ�M����ҼL���'ʉ7�՚�ɪ{��3�
�C���n�3��3U�/�IT57���2+0�njܝ��&��;�vĹr8	0]9k�FIr[\���gM�n4�UQ��xy��P,x<�T8�ګ�ኮe'YA8|6����񛞤
�"<��n`^����tj�ۜ�p�1���Rg���"t��~�=P��k���8�3�}�t��~�@��� �Lm�n)�:�l`��j�-�1/�|�3��%˵�B;�;V�e�#p�|��N�\��G��[���Gq�O�P�h>�h��lT�i{q+z{g�^؜M��D����~��4�+1�3q���/��Q�����>eQ��0����ę�6ܩo�;?IcU�5����j1���2ѡ��9t��X8 �۰4{������o2�^r��u�e�,���ܼ�ErN:�:�:�U�n���W��;�ɖ���hlݶ����˨7��k�u��Aᩚq�����S�O��b��1���\U��rclZkp<m�d:u��47|�JoOkN�����󬢝��4:��	LJ vP����k����%]I��XfѮ��oAv�9t�
kY=)�,-u(*�������IA��J�S��h�K�;ItlS�Q�֚�UΗ�I���z1CÑ�N/������h:p-!����j����Z�q�dS*J����|w-��ef�ޚڇ C�����T���%�Q�n�����X^?���]��!8�*��D�>^%�F����H��ˀ���UE�k��ąz,��0	�>^���5|�E顗Q�8W>��cՌ����m�ۭ��s�ٖ� .H�Ӗ����wg7O�+ɶ�Ίv.��z�[�_!F8�3�xVLMj#U�ú��:��l4y�	�ĴOEx�5�t*�ci�O��n�/�[gv�&R�2{���6x�#��{"_u^�c�a���ƴ�3ueU�t��1w��	�,��뻘EX��ϲ\�y��Z��^4:���_�|#���g�ߜ�!�,��={�v����O����X�Sx��b�ZY��V�=>`mb��c�uMz<��k���t���h]j� ������A��w�g�d}�$���B �l�in��Tp��CQ8��Q[��-��M�&g��hI��e�!D���~ڽX���>�=1pz�9�z��ʂ3���趱�nwL�dC�5��|�۾ע���k�`;_y�&�i�E	L���ِٝ^�T��೚�4EF*����1����P0��mD�*��R��	�#R��ݢP��Է�TZΩK��i�"��5�S���^[���e��n�9�t��H�@^:���給���R�F�
t\T%�ep��L!w���i˙��z�~����� ��y���J^PY銏mf��:Ύ�����U�k�㤻��,��9�aV'�(x'Д4�n�|yMF��c�@��l���<×|���f���K���S7�o_L����cvV,d�^��=����-y`��\<���XTwYO�9\EϬ�:c�5�𨽚2�Ja��VH�wh����H�=5ij��"�e)�8BB5�w���D�QV��zgv��0VU��� D#�\�M��5Y�*�]X��r��'Pw{��s�Ջ��R2nVFY�S��P�y���F��<�2�S/h]V[��O<���ҩ�H<����wt7&p�'���9}BG\S��A�Z�k>��&-�ذ��0�=W���&�7�ޑ���x�釡s&YEry�I�T$�Vr�)�ɼÜ���e���c ��2ݞ�
/z�7c3
ݥ��_�Y<��Z���m���yu�򻏔��k"�ag�NϋO=�N���4�Vo���$�ʣ�㕔�ܘ��A�=a�ȥ���_M��ȋNL�Ѷ��Z�!��7�,}-�Σ��,�Y�������JV3�ȸ���1D�E�.)����]8(p�u�.��b�p���I$�6�3ؚG���v�.@Be ��|%z-��e�pvU��>~�����μ��򚠷і�`��޹I�+N�^۔#=��wpO�����o�3�3z�WL;.���~q�{*����1��;���Z��;� �Z��Ktؠ���c=`m�[�tP�*v���Ћ:�m�=�*�}#�GWl�in���Xk���ܴS1�KhsR�*�B��u7�B�-|p(�/��ܩbh	$l�����j�̵��丰�[ִw�=w/�ԉf��w��G���s�0\%Ļ�J�WF�4�okj��Z�o��#kS��:������^�x>u��gG&i���
˂�0n`��5���ί���X�F�\U�Y�(��η��9>A^��N�i��ؔ�8��f2�1����0��[	�k�D��� �Y�5�S��]^��2�틢�6
356��,��nt�~��>f2g�e�fuG��RWHYLc�������\��70�5�������z�SCu��6:�93�`z�����suu�9o�Z���,L�������̎w�a|\���Q/W��J��|rD��������(bCO�8Cv�|^����;i�G*I�rFi��"큋ggR�za]��V����Z95se����;b:�}�eL�Pj�����jӔR};vX�F
�gK4/%�$�/L���ˢ�Ø��*o-�}�*�Ae���<��D".Bㅈ%Ea|�w��p�v�%V(��OX9��\�%<X�/|��^w�]�ǧ�����S�n(��\�\�.[Rō.5��جZ�h�)L�6��*(��#�+���֎e��DX�-�1D�� ��b��TQF,�rʪ��b��*Ƞ�TEb��j�"���r�X����QDQA� �TTE�X��][][MX,X��ETAİ[K���8��{��~�/����|�<=ub��Ц�M
ke�,�!
I�P���!l��0._���{Oj Z�.����W�������ۚ?)�Ǐ �����}
-^����߯ �;�b.f��l<�<��	�����M
���|{ 
r1�y2�+j�نu�7y�=ՠai���`�L�q�� ���C5�I�܉���g��u��m���Mvh���'c�]==Qu8���~���T�؅�Օc�ogT�a�gQ�<��S�h���W����a�t�M�37�`
�����Lq�D�.=#dY��Aj11y�ϯ�V^*�x]���R8�Ű'D��nw5�9m�\�jW55����m����v�(�f���,��iq^t5mwc�WRvT���_� �<�i�z�<��.Z�&��r���Z���ګ'���!�O��KcU�PUD�-�M��c���Y��5�{��7�>�&I4'k�����4W�q�9���V�]�z�Qk�����j�-������HmC/�噽 ]�Gb�)Нe�N&bN<%����>ʈN\����Å���d������j0�y~շ�E�GVT�0An��Y�3�æ[9N&��>w���B)�԰Hpq�y8h��/żQ�u�+�������um�W#7�R���rȥ���4�{E�7l�OBA�U�M��c��D�m<�����]K6Si�X+v�
�
^��,>�Y��ߥ�9��m�f����Y����A�7*�P��1M)+	5�������vgf����%;A�Ng)
�#Ҕsؐ9����!��c��h"J�_(@zr��̳�l�iSh[�����ԅFfmm�V�^�릋�u	�Pb	w�����7,^�W4Z���}��`i�ӛ&,4�yŒ�a��u�'zM��scX�b^dו�3 ໍ�m��Y��J��/�S!C�SN�-C�Sp5��AY	{Ď�s+�µ&̋��PG<{�8{v}~w�3C<f��]�b˺y7�5��4xV�S�>��3�siG2��eF�pCD�{x١�5�^�bA��q�Ӓ�l��wK��7Q�y��q�k�x]	�|����_xEV4���uN�(+�t�UQN����OO��O_]AWw1ŌU�ߌ\=�կ�#�6�a��	��'&�2��7�;c���!Z����W����J�� ����'��sf@�B//ζe׏�aۻ�ӧzX��i�=r`���ʚ9!\a��f.��S![L⿪��/�,�W5'�f$���]�s-e�h2Ծ�ڠ�����"2��W��Z�t��^��4����՗1����s3-�ӎRG��̅�i�;��`��V�A�~������)J�����#�u����~ˎ��l�k��f8#WI���l����}Cg�H���b�V���[G�ɸ���w'u���^��k�N�Ed�8�24v�8M^�{T\���xjԝ�-c����Qޛݩ�.�vg@̞k#�n�Ɗ�>�1Q�5ұ�s�*&��X�ˣiAr�v�n_��_j:v$NpktR�j�Xd{�RW�#�Ǩʩv6ɵ�6�_��ꏔ��؝��+2BqM�9嘬�Cf�z��T��*�.5yb��1`�xjr��3٠5��%~�WV��� [�I.��`�(��\��o^R���;�9h+G<�W����b1蹳QƬ�O����.����j���m;lѸ{�]�cۇձu��������<O3��L��Q�$o������3�9���U��m�e�KC^�A}O�҃���j}ʙ���-1��ꊹ[�%f�V��i�1q���|t1|����8�a�#�E@$R�w��N���0����z0G��=Il�
��3�+�;��uu�뛰Iz#'���l�H��5V���6�	�N��q��)U�R�*@牜��O��֚�����!N�e��(d��-�*'+F���������8	6v�n�[X��^y^7un�b�������	+w;�&4���ͬ5]P��C�}GhI^񁑓���&��x*��XV��]�V8���	a��X��)t���]VQ9w�h�:e
�tQ�Hf�*�ڗ�B��ʎM���Ů�>�y�ج��^y��m�����4����z�-�k��Ӭ��q]^��s.���s'��ȑOV���e�������쫄����s���{��.X.�Vj�l:�11l��������w+eN�˺<#/]J��s�D���=��]V�ܺ�Ig
Ǖc�ᇱ�D
4�T��YΜ�`��YU���On�PI��:�m�tƕ�<4�^ɵeW,)��v�{;�0�CP=U��O���*�婓��v����M�֛�"Ӕ#!��>ȍu�b�� W-6dŎ��	[�#�R��8嫣ܾ�l܅n�R���]����]'�[�L���{b+�֯{�֙�g! 9荃SC�ꇪ��.�Ղ����� ���� Mx��y�*���ưV�lB�<*�!s$�g�l�p�(�a��\es���&2��yK4��#������JA���m.U�5�1h��"֝;�1]�V>��N�������ɢ�{Qo�x�4A�)j`
���+��Ga�z<��v�˴����B����3J��ͭ\��<4/l�Z�j[�X1R硼�3wP��2&/�*;��r�VpՔ��t{_%�ѱ����H��͝�Gq���뤵!w|�#s��n^�\�	�č��Ѿ�Et�����-����C�9:��}�u�c���ŻY�>��*�EI�*��(�GP�ac5�����*�~pɛu/JM4�q��XR��uc}]@�s��D�V�Y`M*�	�i�yyK�	Fds��g7
��6o�wVr�0��
�c�?Zu�.9��@�fOI�����5���r��{-���ebu�:ޓ%�|E�ܲ5UԊ} �l�xkfvo�,��e�n�(d=�iN�V3�k�N��_o>����x�9�6�۔M����W	�:�[4�
\u7��cXʽ#�YK�d�橶�hJ�{E5����g,�.�K��;5S]JԖ$5��j��d��.�8a�_5�j���i���Y �j��!�y�k�;:�*@��m�\����ҙ�$&u��F��p�B���e��z@,��HN"������ͩXyP�R��H��}��f����$'D:�ܡN��u<�������p$�V����m���Kl�ҥZ�clR֌�D�jU��U-*��b5*T�7�Z��UQE����Q��9j��2�r�U�((EDV9j3-�(�E�����B�+*˙��(���1��*��*�6�T[i+�"��(+Rε�������Ոg�{���vX�)�,q(��@�${�+�jl��/缞5�}��G���+�Kʎ�Zv�Y�w����54�p�o��<
����6�&_�ý*�O�^�S}�1�1G���a��յY��Y��t�y]C�7���F^
3X0��4�}³�:uw cZP���}��t����,U�a�30m�=~wǀ��T2�k��O���ӣ˨��L��n��G�
�سw���]�⛫�f'����3��)�=c}l#W�.���C
W���tYQB�*��18�#�Z�2t2�L�nT�������j��Η@{ٶ�v���bt���"�OA��o7�u\\��ʦ�y~*�$m	RW�;�g(�'�k5j�[m��[��KZϘ�m��+;�����]�7��c��Q��H��R�(�Y۸�C�ن��sD�5�j���y�O�:&�&���n����D%Ս�i�i���2�Qs<�d�𵕕N��Y����_V	��_C�r����.�UܸS��L@y�;m,��K�ۨ�l#���K�:�r;b�8�M0E�Ir)��y��PVS}����Jū��Z���%�����\�9JePAePK�^gŝ��⣘#�h��O��M�*��u��md���6��<�{a��*��&↮���suv�;iZ՞pެ�P$�(zt�S�Y�~��9X�=��wH� f�7��1�]�״�z$k}=�(��;�܇6���^��7S�=�Cb";�2�eԷ�+-�i����7�9��f�5�}(����n⺷}y��j��j�͛i�b;���ao]K|���Q�9����+c���C���?V������j��G)��p��9�s8V(��*��JJa��r}����:�e�Ӷ8���z�j�I�Vء���6��n�c����W(��������@������p�0���z��4l 1;��>g)]_\F���=�-迫s
�8�xz|b�0P��gk�;���W���Ω����(���tiN1|��b/�]��̻qԟn��܅{f(���C�v��9����\"���U=׳J�E��+��@������=~t=���u^Q�V�GH��j+��L�^��k���8;��Z�2�7mO{����ա:a��q����DĊ�4�!43o���4�,�[�)�<��ʾ�1bSG��Aޝ߯yF:�\�M#U���~
�w���j=zb����Yk�c_���r�x��(C�8%<m!b�s;j|H�# ���r�Q>S�S�M:(FN=]��x/ ���Gz��j;�df����A��]Gs�;�����N�K��^T[��$aI?��}���\B�y��k%����$�U?v�"$�����~��`�FN�~F�CDu��z�����skʡЍ�&��t.i��ڪ-�������B�%n��7Y�c.����V���$E����3X�)G�nL� t���g��5Y]<�r����m[e�-Cv�A��5vn��f5��-n\�0�33�^��Z�}^��GQ�xݓ.�J�˃�M7�b��B��~��i:t��u�F=�Yo2�N���ܭo�[;���R#N~������w�?��S+w)����n�y��^�9R:��%�g�����V��T�5F�㷣����v@���^��2��d��A����d��;}ޓ��̬ۄ��7X�b�yq=��t\�%;�ؕ��ۢ!��=��l�V,�v�
�}#��h����og+q2�����;�L~�{�c�1�
���|�����>�VHy�����!��v�xɣvH{�C�'L��C�El!�پ��>dY����̠�W᫦���9$LY����7��.;����Jۨ,����ȩgD����5��NO��UUa~q�}���i��E;aRr�RN�&2m�2NX^���uI��N��[��}��<vI��	�وv�+$9E �������`i$�凩8d�<���o}�ƞ��$wH���N��!�VXT��L���0Ցd�3�!��釉���:�G<��<�]�T�n�8IݲC�Ox��I�L�	˴�z�y�I�=a�Ho���]��N!��O2,��!{�	�Y;@1 t�d:@=d@垲�w����y�; p��,4�;g������Xx�z��I�~Y*�vHQ�0&{������9��:CL��}��0�M�!�z��M���I��%�u��sB)��w�z���7�a
���	�NXx���ݐ=C7d��+kvi6ɯ(�x��$37���^w��~s�=�a���I�!���p���ć(�C�'��,�����p��	�<ߦ�E�\��wx���H{�'(L�3�І$:d��� ,����t��`���ٿ=0��	Y�@��h���~��(�7���4�4]7n�� TI<�3w�6r暷�� �y�T�PN��L�'$�U} ���y���I&�C�N���vp�L���$���c&0�i2Ä���o^w���H!�p�3�NP��p�2v���!׶N����Ї,��=���x[��ǽ�$	�M0�!�6����I��N��$ឞy�Cl�Hv����k<׽��|vIYX�m (p��!Y!��d��N���j�r�Y5�$)���l&��8�~y�vi��,'���,!�:d72�������NP���z�i�����9�{��s��q�$<����d�"�M�0� T6�
�M����S�&�Y��z�<�k�0�d8a�'~Y�����Oi�p��I�Ә��:H���}����=��w"�;}❰���<g��8@:d��9I9-������p�6�����]�}���Hx��vI�;C[�B�M�+!�=a�I�$񓮨���XC���'��042C���㞽�{�� �!:C�Cӭ䁶B'��m��I���&�!�]� ��7�z��R��u����S���x�=�,���3Ľ_!�X�&tWTpvc93pN��)����<�R+諭��h��_~����I�z�H(r�Ę���	��ov`힡�Β)'Hi/����ӣ�o���rJ����!�}`m�6�����x�5hLHp��@��M�(gvb���o��w�~{�>o���@�L�RC��v�ua:Hc 霦2�*NXx�l�=a�x�>�Ǟ{�L�������M�q���09d� �CHr�ЛHLd�<Hgu�7ϗ�P4͡8H��vHv�2p�p��$�%d��N8�C�N���)'LY&0�9�<������ �$퇩��ċ!�v@�'l���uNЇ,���NY!�d�К����\�ռ���]�p���<f!Y�+!�ć(��Hc&�'<Y'l��r�:�N^w���=��I�C��;�9a�	9fĜ���gH�tÍRB�pɞ�$�������k�םk��CyŇ)�,��凬���$��I�E�Av��!Y�4{@ēz�y��}�~'(Cl�1=@:I�@�y���������!��t�8@� {,k�ѳB�;�u���3�}h=�����ym=�2�R�5�5.�_�]l����!�"o^]�o��"�_on�6'4��b��Gu|�_��yXQ!T�],u2z���\x��s�������T�n����A�J��v*i�X� �g^����Kq�dՉ:�M�'7{��f�7�QL��V��w��i�`��}*(�ƀ��s5���m��jTAlP��o�5��.�.6c¥� �RnL�h�dH��*���J#{�T�+t/S��N��%!f����憉V�ASV���Wn�"%�R�ѩ�C!��17�+ɂ��/h�^�R��L�R��qǎ.�7��v�z"o2���E�	���pJE�L�QZ἗sY�r��
zή��)G6	�s�ў�����yv�����VJ��13�;H�4�q	�Ԫ<-���wwOTy(8��]Nw݇�b��#՝.���lU �����_XL:��UϞ�]�.g��X�YoQ0�x/Y�Hg�^���Z�_/_�q��3Z�N�+�a9���6�@hC�tr�9M�<�!���f�+�b�4��M�]*�S�ꫣڨ��h}�Sw9:��sMg�*rl�b���^���s��aȚ�"�nm�2�1`��R-rֵ��u��uv�N Do2V��'����.����U�W����VeرT��R1`�QE"*�؅b���DPDDATX���1��"1�ƪ����c��5`�mUP�QE��EEX媢1A`.YQ`���b�£h�K�G(յ��1�q�Ȭ\���Z�RѴ�(�V��Uj-���qYelUkJؕ*�ѩV���D������02`YRr��)���r�$q0��NI8a�9�j����il��}UOO��u{ފ��d���VT,VN(��������➺N���q-�8s��	��W�Tav!��:��X6�ZW��z�n����r`I��O��'��|�N����V�F��V�z�-��׹x�ߎ�s�/ٴ���C'���57Ǐ��
vr�s*��|M� �|������7�q��p��e�Ν�k��֖�o�k�<��C��]��=��V7��3�/9�����=d�:X�뙄�$��,���-���IN��}�%H�ʴj]�V��DG��y��/�w3���-D����w�����2���x����\��J�y�dY�l�+X�P������}�;���7#��A�r؇X�n�@��B�G�V�y��8f��b�lE�w��������^�jߟ�{��;I�Y0��=&;�$���&�W��a�m���C�|�x�gw��p2�{�V�N�@������K�4I����a�}����MVH�F��d�}M3;�6�H5��[�J�r�q	lA�	NO�U�W����]�u��cb�:k���7¥���F�{����P��{� �(<����\EeEjȫ}U3ٙ͋�E7�m��np�oúw�ӊ�X��j�Y'���F��E7R��Ӏz�p<I����}���w53<����<P�HV���jx̾��%#x�Wfd"�f	`.0v���!㽤���K#�^�h�0/��h��ڀ���%+���Ok��bjVz�����W�ⱛ�6��Y)���U��ma�݆bF�[�^2�r$㟫ﾯ��6�`�@����PDq�Ij-��γ�1�#�]s�'w)הww1�Ԗ$c-�4�RtnF�]׷��*m��4��b����wc'e n1�X���ެ8B��:'/f��&�󡏳�Hn�ط�Jxi�{.�wNEd����������-�1�Xr���>���)��Y����uzXU��嶌�^y�^�棯ĒB��7{�Ц�wHh��U\N�,R�8�"���mQնP�W�ۆ�_|8oWY�]�a����N�&���	E�DDG�i�)��D��*)Wgp�9׏6k�G��,��2�Go����'x�j��(	 �4����W����i\��ҽIrȬ
'C2w�7�{f�~�2�S���#I>ҭC���uJ ZT��"P����U��y��eZ��䥙V����k��h�U���U���c9|�rq-aԺ:�Y��k;[��W8�zr(�VY||3�3Y^���Ǔ��5pӢɀM�t�<9Wi�G��܌"�N7'�����)����\��̹��~hr��t�>���3h:pM�������\�mEpȠ���w��5	��)\��v�||�Q>CݚcyLC�8Akɼ�>�C�ӓ��8�⻍y�<������#���4�k��a��Il�Hg�T�8�v὚�&�v:�6rd��o[��jM�7s��*F&�����>|�r��V�����������ۺ��a|��8�'/p��X"�P]sq8���V�{6�|�+c����}�W���_���@:.f֪�u���)�N��PEGcrw{��1�o� �+�J���כL�	����X����>�@ܶ�=����Nz��n ���A[//�2������ג�!��9�7Y�䖜U/�����9�����{3�o�^��k������]�W��@\PP�C�<u}�L6�xf�����.y�M���0"JAꉕ�÷N	�I���L��o	'bu,�e�g�3Y�����%��km�m�������y��u��aj�ʈͻ�Z�0/Q��nQ��qL�y�*(����s0=K.F+U�T������t�{{v,{G�f���s�h^(\��Z��#֯[�ӈ54�t���U�&��S�����q�ғ�� ��p}�C5Pv� �����smwGq�_K.PR:AB��T^�=�rr�Kc.A�
��A:���KҖ�̸np�0Ֆ��3��u�͙�*������V�z�2v�z�6s{d.�J���Qr7#������e���f�I�� �}��K���.Jef���D�|�~+��%7��: 	��
�ֽR�e#vI=��W-��Շ|�fa�ܽŉ,=�l����ͧ{L�;�|��/7u&������yj�vlZ�ZV�5m(+�}JoZ ��\���Z��8iU�,�B�'��I�K�9��~Wr���w��s��x�_���.�;d/���*�	�k��S���m��*>�L:/������d9\^����.X������G�[�M���f+��O
�o]Q&��&�.�H�}N��+,g�����ʋ��hz�p�wۇX"�^;�x�]yd"�Sţ�[s�P�7{�\�^z�
:F'����/8{�k&�鵷�)�Dt!啞�Yр����<|�{�^����f�c�(�A���Q�{+6ͳ;��Xm�kBQ9�s��B�#��V4�#��p�O�t�]1�%xI��4�)�;��x�3Mpe��e� :]��3����/�jq�(P;&el��Z�Sk�<�S!Ch�Ej�fo]ExE���ˏ�'���ݾ�6WvvC���%�(��.]*)�Ѧ���7��4���ZZ�EɈ�.Yw��+jYچ4^��Z��7tpcR$J�����Ѷ�K;RN�q����I.�Ƞ���z),Z��K�'+���n�2�Vw�K]Ʉ@3f�\�*���G�7-�	6)�`�ID�b|q>������e��Q��h֘�Y�/�$���75aS�{
����&��Mfn+e��O�V��*7�6sq�&_�G�=�.��Y��.I(;��7�;8m�&Ŏ����*D�����Nu��"I��a;˫�,���%,{ϱ�8��ؾ��/5�/0�º)�E�\(�Tܔ�\�p �+��!�ѫPs�̺4�@"��F�ʉ���uR����b��PT�����Ŧ�O��ǼX���]|{��S��|�K/`���y,q�4�X����K	�=R�;�J�k�$֚�*��2�s��/�v��載pMv��6�}}�i��Ot�(,�R���$�)>t3�}r��xoŒH2��u�9�1��hnqL��Ha��^�rSS�f%e�J%��R|�� +R	ό�N�Y �@t���}��{�W����-�Um�ZR��j���mA��
6�,Qb�Q�-��-
��2��\V��s%0���UXҍZP�F!\	��Z&e1V����UDV�)m �Z[F��0��\�p2��VVUU�R�єUm%j�KhZ+Tk�+���R�ڠ�s0�j�fJ�]Z�u\֦�Y�LMe�A.��Й����::�`1��UW-uF��X��̙\�6�T���Z�aqQ��%�m��Kk5��Xj���X�� �0�u����ߛ9X�f��̮�P����͋�椅�?�W��}XǤs(����d�X�$���y�3_���n�`��;�ؐc���,$�(���*��w!�Q�|1���{8tĎ<ʝ�l�g1e�Ih�裢�`]k�����T�Mz�\��kW��]�ς�����x���az�R���'=�7����ܦPp�7ƪ�9�{M+�vķv6+:s��ǋ�СПR��|�����S~�Ô���n]�� ���_N�eX�+�4��1�p3I6�nw��5��]���-�ӫHtJcnZ�.D�s}_}UUiFP>���S
X��~f��-�x�S=�`�vW-W�ĥu_g!���l�����ї!�O��sS=���]IP ;��|��cL�Ӯ7�"x�g|f�$C�7������-�1&aL��Q-irK��������ř���8���zS���D�囌`�]qf��y�W��}V��2��u�a�������̗j.&F�Tv�diɹ�go��g�?:�:$=�ҝ܍�Y�L/�=J�����5+���m�Ӳt;WywEs*�^�q��U�F+�\������DK�w��5���N	���UZ�{�5�!ovm�Gâ� z\�,
x�p�_,��U8.W��ť����q��@C�"��'8=V2xS�(�6:���������T|��e����^�F;()��q�
}��NT����W������Q�Q9㻉N<}gu��Hɑ;k:�ʝ�~��{�x���
�en����;�9Egv<�㲹k4"A|=t��W�+<< Q�,u���q��ׂ��z��z�-q(� RO����Ude��?OehP>���b�t�3���^�2�g�֫b���v.�9Q�ý/�j0�GF�7V�f6Om�7�����X؂65ӓzlqf�Ӝ��qb��b'�;��OY�s����1�����9�-�6���m7Hd�o�n�n��gw5��O��1��G�`�1����	���ze3Uל�G�;���\�ܶ�=�-U�a�6����EgwagO�c�#��w-�M@��lkybԒ��w��u��=���������v�j����"""[�\0QJ��l�������^U�s�D����ע��wz6oTdw��T�3<�ukF�.��=��=Q�C�g�pݶ�QƎ�e���hR��u���a'^oBRb�ϼ�J����� 7v���%Ls��fy�pl�A1����	uf�1�t�w�E 9��qzp��=t@��<��vC63xJ�+��F�K�Als���~'�s���f����'�rW5v�Iyj�c�)�Lݢ��"��_l��ȚROǣޏDR�[s��	��=���ݼ���E{�1���ru�j�l�,9�^d�
hg6��9����I,��]��וb����:.i���Z�|;w�cU���"�VlmNm[��H��|�;��{7�fZ(��Q�����!�n�C�G�3S
\k7�`�aLwwI���E�;�����+e�W>��/^�;ޒ��(�-UYTXZǸ|}�Z�(:��El��zdHe����#�6薙蕼��9㦪�̷np��t�X�Rf��r��������kO�ޚ�O�?�j�;�h��({gӲ��6�Tzѿ^�>/l�m�eD�؟Ϻ��Em��r�u��zե��To�ܥ���g�^�l���g��1���w�����sw@~�[�Ȟ�96�vˍ��:�.tۥ��^>P��K�c�i��H��ԑ�M���s׻[�elt�Ւ�qM_��h�!��pl�Ʒ����h�5l:�%bǠ��	Q�#�wב�4�m&$09��Ua`L��(����n���p�$��U��Ul��۞�v�xVt@_�q%��^vz_��}��n�;�Л�h�'��]c��A�޽��/�\�ΫkL��D����i�1{��s��+���ȼ�{�$c6I�ʭSr��;n��dؓT����{M�{r[����G׽B�Sa�s+�
[{"|�ڿc/Fe1:�kܺ5oG����쇮�3��bM��2���Ք��'�q�m�ZN�|=Ʌw�a�;�5�-� �W��o��tἴ��W,Pۻ3�NN?�}_}W���!��B>����z��v��jiSqi�U�r%�݄�:�6�Z̉AR��fS�
��^��-�2�_M�۫_�d.vp��Q#��{9��5~�5�.i��\7�_{��irܺW�5��sS����3�Y�o�k�'��W|���G��wuk�{�Aل4Q�)f{
�zs({8�LQ)�z�_R�I�뀗- )�
�y�/�F^*��K;҆� ��.�Ֆ�i �#�P3�Vu�T'��j����T��.O��}�f�(�x��4:�����:Jw��]���DrW@*^�N�OL����!Ѐ�B�ml�^��{NR�����Du�Uc�	5Y1�x�C��A}ȅ�uxRz��N�7We,r���y��M�P��]#[���{w~-4G���ʖ�a���@� ����jK�ڛ�"�!Z���}v���[�7�)�qKVi���tZè?���oH�1s��׳y� ��M�H��e��Vu-oKK`�Ki��m��ӂz�Ѩ�-���q�XF[NM��&G�Qo�0�>˽�Cu��١wy�J�+C��=��-��d�8��%+Zu��L���u5u��$�90�X����,5�&@pl7xw���c�\Z�c6�O�Q=�u����O&�⪯�u��.����������V3)`Ü댈�L���f����|�mfWa/6�;�t�1L��U�ۡ#J���7,��W�'��{+&\&�v,G}��Ch�Zht�;wG��ӝ�6��[q!��.���%_bp\�8�Fws�E<�c�tS���,oL$H72ZFR�\��+��;{�A['�(����}c&uK2<[zw��IN��K7V��i��27i��� *|d;�V�v�I:}�f^_8p��a�V�=���t�hl��(X�h�Nr��D�a*�h�4�pu�^��o��.���XL�o'͑`�ȴj�=�u��ݾ���h�A�N児f&,	^poD�|���N�3�(%T�w�ŗ�W8�c+o�����l
o�5�_c\ma7G��Е�����zv����Kl��`���q4��x��QN�W�j�JJ��{%7�u�p���;����LWff��V�o^��W�3~$��d�l �q�����q�\B���n��尭֛��C)�ҹ5����1�aR�mC����Km+m���5��غ���5�mȣZ�j5�VF%.�W������Q��#ur�ZQ���j�iQ؎�E�T���6T�����,U�[U����ˬ�C)r�e�������%)�D�q4�V�1J�e�LjbX��
��Z�Ҋ�1Ef$�Z Ŋe+�)�)�q��6bl��k�ʲ�G̵ˉ5���e]e�	�Z�t-��؂9m���5h��X�Me�(�TKh�-���J���G�9����^��*�%{.:�ɾ"�SU�
�}3c�!)9?�}U_�2f�Yum��|����ҝգ���~�;L^���R*�C{q	*W�;����x��� �����B��s�����0Dt����.X^^�M[�S�:�z���퉝��9�x��|f�_5^���@�Av�]=~�\2q��U�z(Ƶ�;
l'Q��OeU�7V/O�e���{L��1>�!��K���ll�h f2��קN��V
02V�²%��>E^i�bx�_��X����ݻ���LQ_e���M4��L�Z.B���W�VF�\?����z��ٕ�d���K=�k����l`�K����ۉ	����nj�cK���.�ۊ�����0&!^�����I;�A���{M����{��=t��M��������8I��3ʸ�Q[	L�Sv�Z�u`��8�Ϳf<pW�y�v�_sx�͝5�?e���l�'���kg����|�۽�����=�U6t�f�+��RLn>�@�
]v��ѝ:M�Y'�G'O�Tբ�̔z�Xe�2!�&957���DDK����c>�|��|��z��f����1݆9�fW5OO�;��T���.����PΩɯH)���lm�� �
|!O�$t
v���;
����<	�ܭ���j��"����P�vUy�Cv�TXb�)=��ͣB��f�\e^�\�j��p��Q��9�5��5c�u*�/Nz�>5�'�ժ�/r&/|_���t�qC1c�~�������>�sH��;vE�Tz���;zN��Gb�+�ht�#'��?W�}B��[��s�8�`]P=;�E�yvq��[ː�Ƃ������	ko
u��ܴD��N�l,�F��9{��v?��`*�y
�"憪n�55��u�A�^K�v�/k�j����I�Z��9D��}�Ahܼ|�}����:��w.�H]X�piya�6�H��Ѩ@mm���/��2��:�*p��`ra%h��]��hK���/�/Oj�i@d(�(^͙۫����y�r	"�ﺂ+uܾR�˫7W/���z���3o�Q�]����,m�Ms�y�K"�P�2R༲�ۑN���S�������ݫܾ%����6�-{�ս���o$V-C��3]��#+^a�2�U�o���*�>ϰVSY��� c��S�O�[�+n��y�ٍԧ�4��O�v��b���w��go	0'��z��ܩ�xDo:g�so^���
�6���h�Xd���Kz���®o�GP���]���Yg�:<�ˣ��Ω֣mn��|��]5��E�'������5,��c�������^(D�;�8�k"z.2��#n%��	�r4�q�e��ZY��}=����s�^�"��7x+�o����(v��5����,��rH��n��*��f����y��U^�:�M�C��x��s̩��D���������CKaW](*8 b�Һ9�R)ǯ'�9�_"��Rޮ��[��}�y�ڵ!t�ښ�#�[�7X<@�BT����Õo/;5�b�U}�sq�o@���`⻭��I#N9�ﾯ�m��8��N����o���@��۠�}�z����������f��C�֊5��k_���(S���m�f/q�q5}��~9N.���;�w\D�]���(�F|=�z��=�p]�j����x��y��O���[�2�4�x�G#��gvEJ�)���ޯ��>�4~���ӈ���+�3���l!��c���cw�[ӦO(�Q�7eA��;YW`��,�������y6��
}.�X�^��"�Y�jr�����=�;�?�5����H(ߦ�Uڙ�����aݡ�3�I�pi�÷W�������X����P
��f�V��ڄ������M��6H;Pu1�s�4ry��AuO��^��W�a`��t�	�~�OFW�#�F.M{7�F(���:n��ywGU�ۼD��od�;��0 �}�s�մ�{��[��#ֽ�j�M�a����m�i�Mv�fh��G_td�.w�0��o\��z��U��8�a�#RO�|����?�o�&zEN�9{�Q�%���VVխ�s5�wY��4�s�@��� ]=��E�ؖ��F���9] ��g&�֔���w��b:�>���R�;�Thm;�ݱ�2��N������-D@ώ�S�ԡ����("�{6wJ��qY<��7�>$j4��	v�+>�Q¨�������(�ʼ��l�P�s��5�j�1�J��cF0��ԗy��Gbܙ�E���4rV���$+[����U�x7ٟ��._�Lt�ز�WTq���`v́�I���˳�9�����W|R��OkE��yoD�%G�q�훁G��띻�;v�i�D��ތC���I7r�ޤ�1�e�He�"�'�{��B<K��b�\��VCrj�+ڢϮ����<���Ci;Ĳ�����<C\�p�. H�f��V�w��s�3k��sk.���N��I#��CC�X4����{�,�ݙz*�l��s�s�霒�f�%�V���k\���.x�X��n3՝�
<�X� .�u������h�V����UxҨ���������*C{E�Uݾ��EX>�i�JIi�GyN�r�-�+lQA����TqZV�8N�ִM��v��Ƭ|$�%� ��G�!K�<���t[�����t���z8	m��#�"���J�
��7��.U��2\�&�VK��r��u�p�V�牝y�U#^�+hE�r��O�ͪ/1�R�һ혅s99ԞiR6;1=wR]n�5}���� ��C�$�P�G�D�em�%C�-�<�g5Ś�[}3#�y�9�;;"н����*Z�=�@�Dp��٥�@F���K�\������.kb�J� c�����Yk��CU�Ȼq,���v��)�F��aXL.��ݱ�b�+8�ם![���0)ۗR^.�5ҁ/����a!���Wb��9�1C{�ͼ���mZ�[�w* ��c�\��ܽB���݆��e�S`=��pB��YI�{� ��ce�iu���o�a����ji�$fB\/dx�YXԗw�2�I��d�Z�wV�Y���1�fsW�),W\2]=эvb퇥�$h2�j�5���F�V���iz�rfJ�.�
�l�ũk��UU"��L��EK�#�����\1][�H��,(�UW*��Z�-*���r�aR�[[Tf3Y�u��jf��-B�+Z��F�̕1��ff+UUU.a�U1"��՚C�SVGE�S.��.�p�
jم*&��"��qZ�VVf��qSkr�Ն�2Tr%1�&�kF���
��MTi�������5�LJܥ%�X]Q̭²��al��0���Ma���M.k
�(֎Z�U���e˦h��-����ؓ&Sw��0(v5�Rn�N~���#/߿�ڽ�rf�<�/xΜ�nF,�p��r�ͧ��O���-	����j�j��P@D�����s��;����V6����U#OW8�@� r�rss���[�߰�lN�8s��ş2/�y�˪��e�a���XT�X]��:a�ڡP�	N���[ف6�����{Q������jwrAf��Rj��c30����٭7�ͫ���6�T/n������~�/��3zv�ɰ+���k�9\6���S���\�I'���K�ǩ�#�lw�*�&�co�x>����y�-���ez��g�	�u�3����+}�=���Ԓ��U��U����{Ń�9���v6��!�S٧�.�d���2�R�k���i�w�߆9��8��h�.�x�^����pp�geV-G=k���އ�O[��`pXW��E��B�>"ߓֹ�:z���yB�s�εd.�(Q	�q���@XcQJtm�R�<�$��hi{�M�\I�bm��__�d�cG���ڃ+�+�'���Ei~�ޞY�{�Q�˺a�GW��,�����1Zhh���ݭʞ=�Cjz{85m4��Z��Co/|���\�Ȩz�%-����u�A%3�q)�]��Q�x�o	�ǔ`�J�$3Cxw��<�[���+Ղwq���D�i��{�w�	{/�W��l���Я�����/Ռ����ZEL\�u���g�zr+��Ձz�jT9��bd��m�[��Aj�u�����r4����}�$������W��|,هYq����a"�[��h�o8�q釾��0�a��.��]��q��N�硝�fx.;|*u�ֳR,_v8\<)Г�y��4�ٮ: (ON1�]�y�Ĩz =Q���=�i��enE�'}��7TP��.y�X�EvpVo;������F��x_�\�}������s#]���x-}���͂����6�����eZ���Q��D���ޫ�r�Qy�x-e�n��lTެ��-[lJt�Z�-�o�|\�D������+�ԅ��i�ϕ�}�5���0��=V�F�KRT��PJ�$C�Q��'��S�%�GA;>ݨ�����9�p.;7��i�Ԗ ׺���ѫZe�&}���Ь�Ll
������d�H9������X��u�c�%�b�t��5�Y�7[�5��b�!�no���@sa~I<o��u1�>t5^Bz�%ca
��f
�MT���DT�ϫ�&B�aX��lua�<�0i�<��;�[P�O�{$;3�7[�ə�D.p�gOu�ң��-��_UU��_h�R�Y��][�W��zZ��<:&�&� GmPS�S0�d{��Evw=���=é7u9��`�zp��]f�f��Y7*'Ǉ:P�E��/(����{}F��m�GS����'��	f��ec�:����>۵�q��`��8����e37�wE�]Q��o�a�H�!�3�隮���3v���%N{7S��Z��������p�iQҚO$B����{�}����F%�/(��I1Ͻ�G�;��H��m��&��y�f�J}v���������u������>!��a���n�C�q��&���Eyt����T41q��r��ӯm�E���`i��ۤX��b>�����a��L�*Ee���N}7Kͷ�J�C�i7H�X��KΓm�#1���&��3؍��:!]�M{hߢ�v���C��p6�Xn�e�u��9�G#f�ͧ�O���m�����t�A�W���uw�^�\\w`0�p�u�S�OT^���+�	�s}����z=�DKY�Cμ7��w�������e1�S��{sT�j�d:B浧}Cyˆ�r���.�,��2������Cc:wض/ �˸u)W��0�Ù�N�櫯a̧h�q�:ú���Ȩ�P����nL;Z�����;Y�>d?t��'`\�7�!� ����{pj'�2��/!q<
ŕ�⺺}.?q �:�G�㾙����r��>W;�B�x��4V��fm��XoL&K��V��ȸ�O��<��μ. ���*��+ǳvNr&���舏g�V�=�H����n��3k��j��Sc�;,^N\T�LcZf��a�
Z�eR�9�f�v:�� �a�"�\f敗fd6���q�⬍�MB���,u9�a���a�#Rٖ6����]�2���~��Ѻ�\�N}ܶ&�Ұz�
�Gb�������N��uTѾp�FɅv$ʝvw�1�����$kׅ���VQ�ZGdvEc�����A\k��e�[#&�wppmӠ�A��3��G<��M���\��o�l�򚩾�^K֙.N*I�����̔���S��tݠ+0�ȥ�	��Q�J�W�_�m^]l'�[������w�盺��τ�2w@�ń^�s�W��3��=���^d��!D�(�Y脊��^<E�y%ݾ���j�P�_,!y�����?Q]LI*���*�b��0�B��بت���7lezX�[��b�D7яr�|�_�S�a$.�����^������g�?2�kP����aG�=�mS����'b&���[���R���x`KHz�������ofxqB�b���Pgz�U9ؘS3�̯���Ď7礞�~l:���_�v��sk��7Nt����&-xf�9q`ͫ�kvX�N��V��i����]�@��Vm�WI,��^B0L$�ߊF�c�˔u��3F���z�	���LK�A�ܹ0�>���R.���!�ꕝϬ�\m=�����^ʹ�eodBLQe��»)�|:3���S���o�TX��J�
���+���u�"���H�N;_nc��F�&�6��Rh�$B���A������u�v�:�ucɃ��\&Z�{h�ui�Ƕ9�5;���V��2V�{xU�K=�] ���{{ܳ�4_I��wL�1��դ�0�.����Sk[ך��p}��)��
6�&P�J��M�V��ٜ�]c�y�t�b�f��j�7����u��7�\��[`��;_p�9Q�c-�71}ݳ���\ZRL<���.���9n��?J�}��,j��e���ክ�^"Qb�6E�΁�ڧ��2P���/^�An�Q�tmrܠ�,�F��eP�d:ւk�Y��VpEr$��(mU�k��y��޵ʞ�L]7�=������wqP�������X��N�2��&VAZ�i�L�#[�D��l�V�I|8�7��@�&�X�m��7;\��5%��X��{6�.t)�_:�\�}t���o}+���hv���j�5cW�fc��-*X�z�0n�V�m�ikiF�F�Q
����a�JXQ�]�)J�f-)i��E��ʆ5,k-�c�SV�]e\Z�p�$Rڮf	ZT�Kk�33*�`�p�Tr��p[����
feV`�����1Z5��Fcb�b�T�paR�Z�-�un������R�T��-�+J�J���.L-Y�e�+����cEӗ*j�A�e�1�Zf�I�t�2�[jS+ciq�.Z�-V��Z*�_��(wO{���~�h�3��*dpme�(��J��}�}�z0�??��@�:/���1Ԇ^?]���,wKw��ݓ�y"/�aԾ∾TCi�o�U����բW�c_��܇l����֡~T��z0�3��N����#qY�)Y:��]��e�~^�)�e
�њ��_-��a�����Uut!��l"�@�(a�!��Vct�DPX'����K�u�6�w���B���2������`g��ɟ�}\���yi���w� %�����8ޯ��Ж��b�o�]8����5Jd2=��[ӵ��X(ya�WϏ]:�d�7�a�K�]�c����]��a�w7!.�B��wL���7
��3V�H榮�@�p�
s��U4�y���D~�t�C�}�:Y�MZ��nւ�q����зn��N���i�C-��8Qyݷ藅�߯�D#��	��Wy�c��O�|�^پ�!��N��E��C���]k��EM����
~O�����`�r��!~���	���l`�j�e�6�=��cRW��E�C��b�Gzس�r<-q�	�(酑�Ʃo=�ǃő�ֽK�a�E�*��@���^���}2��ayiI���_2.����n��{+�V�����Y���c�	���Z��fի�i�Yl3�p��w%��}#�oMɂ���LV�#f�'���Q&p�<����-2�)6g3E�T�r��Q���%�3���Q�������%�r��C��^t��
AVE�c�?*__�l�j�mι���=��.��z��F���E��FV@n����ՠ�0���VE��4��3�b�Q��g�l-��b$��V�Q
о\C6G��>=�q��<5a�2���-VM���b	�fgZ�{y3�70��!�?�kO���"R	*/����o0X��u����r�-/�B8E�����<�W���${B��=
ha԰��AӇ�h^�{G��]mz��!�C�T��gT)ؘj�o_���(x7nt`�;����YX^��+hn-ms��'n��
W\���Ҙ���ufէӕ	Ŷi.$6Ɯl�x�q����Y�H��A�:2��kk�����l^�vw�O�z?����Y�Pא�\^�MV�ŭ�q���n��U8�3s�%��c$ʬ�]7'���a���E���M�o����x]N9/zl#լ1�T�V�ݡD;B~�����U�,񔅃�*4l��"]�~Zf!��6gm{en���F�,.c�b�!�� �]��6��vh�ڇ41$h��,�A�"�i�!��tY�uy��gƵ}f��A�쁿�RTκێW��F�)Y{o�b�i�����ҍG�6��^��ϴ����njbM�7W<���*��(�̵6����f���ٻz�d�n^��r6�z�32��"��6�X�><@�l�S_ŘmON�:������'�V����ǴV]��j՜vA��pz%S�V��0��?�À��r��i#�^��W� qDz�yJD�Ss��^8�8���Y�*��#�T|G�&����U1�c�F������y�@�;�ƈ��(���<��d6�
�S���9�+EDJ��ƞ�ȑƏ�~�Q�KGv�o�ʪ��j����./�!�6��de��M�y����/K9@~���L;^4`���+�ژ��)�V��g����a�V����C!Y�w��t���
��[/lV'��>ٹ��k�:W��
��lf�5q*��
"�lyZ`SKK�=Pc�Sbw���ۇ�U�CKH�,d��RHi
�J�)�|�5�w�����)}��8s����tS�?+϶���ˠгӴ��n��CKN,>�p�u�e�>�����0&��]<��c"j`j6Ik���:�A�	��r��aӇK6I��{�%S�p"8�H��^-kt�^L֡���m]U���>"�� z�e���.Dq�/u=�8�~�pV/l!���(�E5\�DL�W����o�k���}�3���iӺ�?e/��E��;}�s~�Z�|�|x��HC������:jD�w���s<���R�S��t��R�q�^�Y7�q���*�Q�.S��i�q����\{��؃e�$���W��dz�d"2}��Ε�q�\x�`�����!흹þ�1����e ��X�֔�0�������,#�e h��NW?�C��`��_k�o����yx�7��֖9a.:�*`�����i���O�B�S���	���/P'��هr�{�K}Hx� �/��AUn�!���Q��|��C��`�b��^�4҇���O�vq��'v�� �<|<����b�8�Q�f����"Ik4n�^�3QBh �҈�ؾ\C8Fy�X�]=�o��;j�	K��!��ɋ�_����u���z�7ZԮ�B�l�g#�1��87ț��ܝ��k�ܻ�4y`2�Au��ԥzo����ꐭ�2��b��5Z���-:t�GH�)*/��;�y_mγ�����. ��4?��J��J��RW/���H�
ȣ�(y�X�xbZF�4~�#դVmn�V�8����_��8�!ٯ�+V?ozmn�Ɗ��A�t��{��(���`�޻���E�F�.�F�6}��9 ����*��G�v?���`�,�|�I��X�)�+�{�c�e]U��E�q�@,����x�at����z�؅�}0y�����
!���:=��ۙ��8w�bˤ;��8|Q�k֯e-�a����/1:�9�"70�_*����Be���%rz�ϖ����ˤ�3��-o�
ɭ7E�(@��{{u^��tn^�����RX��z/E�d�kwV��QB��x�E0�:��V��<~���4;_{�6t�,#�܂_ؐ��)�{�ҵc�pd�re���޸�];1�?qӍQu�����N�j��qU�tCw>0r��^!C'��vVb �u��!�tb]�|~eV�ֱx��CӅ^�`e��&͑x��P����@{�.S���3�۸��?YGyV)H��%,�r����2_od{�!}�gH�@�.!F:���⍧�kw�/��"ֈ�ZB#)��Y�+!�[g�{���?8��0����^�X�7�6"V�s"����:����w�-�u���pY(
r��E�܎ȣ�.�!��\�R{��H�޵���d|Qo��\{��j�+�ᔸ���c�l�e�2О񞭴NObOL]�,񇍝�s�v���ʡG�G;a�V��P�6�޼��:6*0�U��:Gac&��D3�=�\��\�z���+�V~v��/��G}�un��ۓh�
CH�j��Y�C��il�uxp��m=�G�lab�/Vb�RD"s[Ӿ_Y	���[xF�YGu
���\|_��.��L���h���n�5�i��H�����<t��ֺC�}�u���+^z�%�V�Z��úED�D\Ź��/w�*���8�{ �t������)��Uq�	�H�F���E���r�z)@�B��c��gV)��BJ���+����GW�w�H:�ރ6ʧ2��V�;]i�\+W�锫6�����Ϩ���QWʯ1K͖�Xd�lc��N'��6}���Gb�%�a�����Gs^���|�[A��t���i�:oL�bZ��yQ\���)[.�k�m�S.�Obt4k��yG:�4;n�Wc��)�Rk��YS�x�͐��-�6T$9�wM';��n��싴�vi㲋�����+Y�s��q�3r+J��ʇ9Yi�x��.�jr�i�F��4!Wz�ۗc;��T����n�S�;�9�nd0��K�5`�W�k�E��Y����[ӝ,\�e��i���i�����>���&�c�̮\7��3�E�& ��q����1EUVT�9|�[�B����p��o �<dV��uc��@�&tT�=Y���Z�!�e.W�n��7w�i�������yG2���`WZ&Ԣ�V��8@�zQ�ջY	.Y�}�q���(v�i�vY�˳--I��������M��S^���*�z�2ܛ��s�O�m�j����KA�קea@b7��9pm���e1ę�WwY4�Q�̺�SV
6����F�[e�-s"ֈc��#*(Ɉ�K1-�pX�e4�W0
��LaQb��#2�"*�-�ar�\Jfa�TUa��镗.9J�*��1�ڣ1G�Lc�TI��c��i*�t�1*��q�����q+1��D`�m�̥B䢊��2�lUE�X�m*U]P�"̸8bTKe-.S2U���e��Qj�%�-bŢ��RS��]�μ��:N�޴s�^�CsJS7���'	&����>y�E��l��d#��/���¨���;엍Y=���x0͝"�Aj-#��0xq�wk�D�G��D{��ׯL��~9O�˞�>�X���s����q'�����4�6oo6���r���<B!]�X�⼇��ϵc�����%��$
f�P���0�"�iO����p�����$�㜾ȆY_C�ު��Jymo!�	�L#q,�mx��j:6nȮ�-���"�Q��*cK��,�N|�%��Ws+�v���5,Zt�?P�dj!�`�����^���M�;��+˯U�ϔn_h��st5!�<��m#�FL�{��SB�8���0E�I/7���Ԩ��������jЪ���z���Ǝ;���v��Ə�����W�Z
,�>�8��2{��tL�ݞ���/��%�#�\i���s_�qaPQZ�wz{��ã��
:są��Z���~�{=:��B��T6�Ǖ�IiAS���յ~�����.<|{�}�����h�}y�:�ђ-�!R�V�K	:l�©9�no{z�y�TWօ��B�G��cP��=�v��B�w�f}�4Y� �S�!lwAg�#A�=<	�_\�5#�d:y����Fϲ� l����V��J��qfNz�6,*�l=
���Z7&��I���5ѺK�eqz�.^�7@��蹗�ȔNi-*�w�_ws�b6��(� J75�f}�^�E��f�<z���#qa�0�M��*��_��hdVE_0����8r퀭Y�K}��O��!�i�CA�v�4l�D>���i�Y��V�!Gg��h!yis�=�1�f,#���\�CvxR�S�B�����4֖E�q�~������v����5C��x��dgڂZ���}x�����}�q�q{�pg˓�ｎ�ҡ�\�n��y&��x��#�:�X�>3���?3o׽��zs����V?�9џ%�P�ʭa��1x��Sws�紝��Wf�n�5��荵:�ֲ��qT��B�����6ƥ^��q�6��ެ�Tp�M9P>*P�X�u�,�ܿ]#^߰(r3��v��N�CГDQ�<����\��(m0�g!�2nߦ#��H�ǈ�eq}�Cc�1]b=^u���Gi}��A�Di�(����"��4.�1v���!��x�Z��;�1đ�#>�f�]�c ��2������q�b#lc��=����Z���ԯ�TB�K����t������/C"�!��c`C`�ڡ�5�s��y����=�ʵB�ψ8���9�Le����6���(�p����+?YGq}^VQ�g��յ��{�T��-Æ'�~fz�r�q�^�(�kF�U������D+��p�q�r����Ӧ��zw�(�RKh"x+�b�n����Ph�Jby�tl�&��c	1�T��u�,�&X՘����!w0ķ�|��W�9ޫ���!����B�cN��g�?3�r	�r�q��d�"�
>-!e�����Z~�E
�ޝ��E/1�0�g��~4:EV���{_���j����pY�Q�Q=C�vjx�K[=ވ��cq��+����W���u3�R�t�|�,���ƈ�T�u4]-/V���;��5��z�7QX�os>_iB0�)� ��W��g�L�RV�{����dq�P�\Xv��=�����D��?]
}e�[Z�c9�IP)q���v�%��%�ˆ�Za�Q��U��0�Sý&�-$�1��FS=�9����Q��6t���+���]yY�<a�\G�<CN��n/��Mx��}�t�w��o2�C����)�/��0���9���{�3�i�lc�0�Q�q�vD��;p2���2�o=�C�P�����n�i
�V(t�/۩e��Y��ܹ�������N�>7ʈf�Q}�����^�}������D�0���v��qQ���͆���ӧ9p��R_a��c�nW�*}*���d^k����t����jե�\����f���O�q_!�f�w��{k4X4����)��0[�y���^Z��J"Kj�bN˧++��:��O�/�D�k��JI�ۛ�]�r�d�)C������a'M�uN�[~6x�#��C�[H�|����EW�/۬�0z��#���F���C��|Q�x��WP �Au�^.!�2���/��+>���_�/Ҁ�!���o���Ȥ��	F�=�)�];��آǛ���<}�X�ņ��]��kҽ]z��oW��8��*��^Cr�C�"�*q������פּ��ł��7��Xx����c�O��5��cF�������_sE�pp�;��dW,:j׵x��1$h���;q��O1��s.Q*/%N�������)�SG@*`i��D��Y^Q�L����Uqe� ���X�Nf��r����u���r��K�v"�P�8F�u}�[�s����9�3-i���w�i�|�~���c��yL(��>��s1�ܸ� 0��'}3���u�C�l�{�w�f��k�)��~�}�,������h�<FW��a�FyvfiY2���}<��VG��HQ��r��;H^��κW�+Cii�F�EZt�l�E�!�g�|��oB�=(��|9h.�Y��H�2��Q����ϖ�Uo_���w��D�C�=�0��J<iZUKҺ��m 	���VGjf:1q�1�{P#�[���P��E��ޒ՛�*,2�pkV\zrؽ휠�Y���Q�/,I�p��CȬ�}2go\�y��wW6���BDK��D]����_�9�X�߻��}f��d�w�(�:q :+��Fn�����RТ&���:f�!����%���c�nV�gUz!DY9Qt�o�V�?;Ab��6H��V��;i��z."yC:D����ǖj�Y}~�������PIi�Ś(��1AHq��ĵ�}������_ȇ��<�yo���c|���%�v��EG��Nde��x鰭��B�A��<}~�bSqZ%?Yd��(L��og��W	�Q�j�Bמ�x/��XD]'~�b�j��c�;t0�$���#2�f��huj�Ce[�M�VH�q���0��9����jQ�ʸ�$���P8�Z&�Y��������'dO��#uY��B��0����x�;'�>@e4]c���oY#�Cկ�Q�H�n��Z�?i�d2&����>|Ib��jy�mn��]��>��&�}Y�$
�+�0��GJ37mU�u$TZw���/�͕"�dN�~t��s�$)�&Lڦ�uC��RU)3�2nzk��D�%>ͫ�ia��_��,[^[Y �ٌN(�BWKw�&�˘3�[7�̊��x��{��w��1�F��G�ͨsa_KU�q�����2�9;�y�q��:1xѳ��aG��r�PZ�-��t�G�z"�ʹ鍼�n�y���.�h��%���;nQ*B8�]���%N�U<@��+�ڄ���P�g�L��3 �`({�I��c�ݸX��*s��ǳ8}iFi��K�\�A����P�5�Ȳ!��7	z�;�%} 뉈F�;S�gQڶ�KY��ZF�bV���8�#{Ϯ��c����"���mh#�=��J��XI[;vŗ�G+��"��7R�*�tw`|�zV~�J�c���<���eД�����ob0+Y'Hs%��8�4`L�.K����d[i�M�(A����&��S�$Է�wE�!՗��>�4����u��^m��P�0<�p19���PZāi�h�[��<Eԣ2i|��W�ex҆<rwmӨ�F���	�{T��d�i��J�E�Y��̛Qfq���y�R���!���.���q�M*C����=nj�j��Z8��vd�'#�wF/'�Ŵ*"#,��JPف���nl�j�t<�X�赙�:w�BM�k0��.�p8n�y^#����)u9x���I�zSv�}��ހu9F]h������V�.�N�Q�|~��Y*���»]%��5���t1���i�̤otJ��^Y�x0�i��l͂9��Z��p��ӛ3ajp����-˷J�s�R[�%�K�T7�c�U9��@ !:ш��2�FڋZ��������ՌEF*]e��e��1��m�s0���̫&8Ҵ1�1�ܦ+JR֙���,�\T5�4�VF�s3&F\�0�XT��lR��emG(��R6ª��2�Sem)1 ���+�4au��)��Km"�r�j-�d�QV��G�W�UM4��-��̸eW3Eq��E�]k�9��z���u���N{���M��C�R5��2�,��m(`��F�ѻ�u.�c�L��b����ah�D=����C-9���Q{R��y�6X���At'G7na:R�D�ʝ����ݫ��_n�O.<x�����4;"�]H[�����	�X��0��8b|��n�e��"���:�?�+�a.4X"�����ӏ}~�a�M���H�	���C��w��7��[%fҲ�������פ6�p���7Oc�V�U��|a�������HHz��+�0К�uaU`�N����{��L��86 H�Th���>{�%��bX�e���&�u;�[;8�5�e�i�sR�����uf������A�7���i3�v.q����	x�ڰ��vt�l^����e�p�{����2�e�#�[���r��_Ԃ�vo��D����}p�Ȭ�P�:@�`��L�3��P1,��}/&��;UY�5x�t�$��t��V5F�/w]y���v_!�����5}���$k�:Q�)�V��5�+n�~Zh���&t�^\t���sw/ �aE�u��~X}Ӟ��r�W=�[&��@�4��2_��םw�n��vU��d�QC�S&��G���8p��9�$Ë��kZ~>Ǥ�4���$����	'���֝:̝�puq*]��Z��<�:O����c+�7�{��&I�6�_u�ğd�H�k\�e��(�;�O^-q��z�!ZӧN���R����ym3�����6~�Z���h��i�������Tw��zC��BD��1��U�<�=�r'�ɵ�J?q�g��/���L�D����b�������o#@�b�:�0�F�a�����v��}D,�V��3��-#Mŧ CPP�l�!�̳ח��9ho���8���P�\u���M��b�}�������.гF�i�B�Y�f��%��J��m�5���|������!�$H�EU�G[���A��{�tB>���@�;�N(��1O�!�l��Wh+p��vi0̀ڸ���5�{�j�
��]���;Tg% �c����򺛽��V�4vgf=1�œ����fo�Wq�j������
9�"S�R�/�t��!ۚ	��Õ;6����Nb���6�9ij�د۾�~#�Z��c˘�F�8IE"� �]�ҏ��d�{B���/yg���E���8n��]��}���yB-�k���O�ܫ����t1�o$�B��>~y�w:"�d^�O��h�-69q,k$!�1�3�{��W�{�<FD8ED��b���ω"�T����Qߩxم����!�YT��fn�'fW�0����y��_JL�kń�Ü�/I��|/
dx4x�+�'��0��4����z��/.�\�Ѳ,)���z����)�.,f��oHi=]��D;6N��G-�:��:y�����یVec��ְ��е�/�RX�0��ء胾�fKU���p���]1��!f�(�T~^�������2�3Ԩ��w��f���Ӟ��d�'�K�3'��}��8t�|���x��#��������l�c�^x��Κ�@�{��/�B�л�t�-oe[��0y�n91�R�:/�Sz���,� ��'�	HQ���U���8�ɪok�<"�?c���x���,�VU��Y�;��_Ak�1c�\j|CK�3C�z��̪<Ej���c�$a��8^1�뗚k�뇡䬋>�d�a���,@���`|�W��,�M~ٞ�\Q�u��b�m��,�l �75=^�f��cu%B����J�7I��zm���![xR�dg���g����0����7�:�0���k���F�(�`���ZA#kC�ŗ���6������/��#��?f{��j6����Rs$���CRf���[X��㇏�l �����T��!��#g�Y�sTt�B�}7���3��Õv�α�KL�#����-���پZj����9~w��@���P��Z@@��K�c:�����,�d�G�{�s��ZC;�#($l��]CW����o�p:^# �g��BTt��#7����K��nr��.TlS_#�lCx�U����|wˎ���2o��,]�M�5��
��4(:fqc����ts�c6�����m�[N�r\������(U�(��
��JcK��$�U�WO��|g���W= ����>�Rp���β���=����oXG
�L/���Q��S7�ٚP�(~=�	�H���"�	*�=W��7�s���$���ˍ��sH�kN��(�r������w�ç���mϹ�E��r�l3Z#b�W����8F�<wV��g��J��4�w�	濯��$a�_i�k�^*#�L�d�����2{@�~W.����ܯ3-���u�ͪ���o�L�)�H�Λ���v6X5��ą�m?Y�x�����m�$��V�9/6��\p��Uøn���b�*��)���7�j�8�)��I#n8)ۭ+���8����j�G���<wB�
��~�n�f�lc�1�:�b՛8s�VD2�8C����(k���^��Y��K�dC�T�B�=B���C���޼�-v������-8r�0�+��B6}s"��U�·GJvw��@�/�sP��	��5��P-�owӄk�a��8I�/���|t��{�n�{e!�EdC���f>���a��h���
��YX�����^�s�i{kW��x/��,7��mf��dJZ<��̻v�1VJؚ�Lpuy1=]'S8ӴY�\~�^#�23��q#-x��8�2� �L���(m��*�����'�{=z���y:�o��H�j5C�bv�E�+BrklN'*d횃/�x��U�E=�|U����[WQ{�^<A:|lr����,�J��!�aE�=���U:-P#�J�z_s��Q��a,0����r�z�Ї�3��}�|�����Ǐ�lT{�/
�ݹl��a�,&+6x���\~�CZY���ӯ���(EZ񻧄�kP�gZf?W!���������G�k���y3��rл^oc�1��M��i���G��,�[Zl�Y�Z�o�9���2���ֆ�t�"�D�6t�=��I��kp�.� ��3dxu0���9�C�͒Ds>c4��l��q[%�gz%SSe�+H%p�b�u�a\����ٜs& �b%���r�tyF����^��sֺ6�}���eMM�#�+��̉�n��'jDJ�*0T�+�������'�!��yi�����Z�	��봶�vf?�(�!�_0p�#f2F)C���� �;1o��1��p���P�1j�0��Y�x{�߽��þ$=���0�QW��+��!�~��9�YYz�Qdh6FjGlk�Cn<Y<��Iw��<1Q�P��E�Қ�;��I�B���UYG;o0�5�	F��=-�,y�e/������7��s}6���d3f�W�Q�i�T�k�=��&�������tgytn�j��x��O���~���-O������-$I	�?/�$I	���,�	$'�?�/�/9,�,�ÙL��?~�5�:�M���')!HJ�D8B��I9?;<g>�M����C���� HO�M��9�����������������x��hp��f�����q��L8���>�H��=���|�� HO�����{�|��� (q'�!I	��'r$����a2��Q����y�8w.�H����!o"�o���)��I �Bu� �����߱��ݓ9��L�>�����o���Bl�D���'�u��ӜH�>�O�������ݓsm������H��Ohk���N2nB@$��?^X�2qҨN�Jaw�\ϿG��Jr)b��43��k	�J���Dd�XA�"Ӿt	���$��>U����?�m=�,�	$'��I�O���O���ƛ2�o�m��g����}��>�����������]D�Wu�8J��Tjz ��-�",���=�!�Ss���\���0$$����?@$�������'�����,�N]��/�A��gFr~�q��BHN'ъ�	�����I!$�c&�6r2O����k����u�b~ǂ�d�8⟬�[�ɣz��4	$'f��[1��3����iC�!S}C�	��Jp��@�c3�*f�j�cD�a����m�K}ܛ�6�x����q@UMD��F�)�̚�Tt/9�a"y��;��?��x|Bg��rM�8f����т!���_��I���}�����퟇������Ӊ�0��OC!@UF���@We��6��$���>=Ϟp��<��n�A��%��v`$AT{�#�=��[!�ߔ�5��I	��>P��p���}T�M�x�N���,�n���	��?�Y'~Hw��rE8P����J