BZh91AY&SY�KR��_�`qg���#�*����b�                                              �B��� U@�w| h�p A`� p�     0 ��*�
�
 �@         �}R� *E(�E � $ �(P���P��@�*�T))%	UH���QJ
�T��JI  9*�@�@P P���1��mMQF��DVp�j��u����{�FF!>���wJWvq\��
 P ]|��� ���gJ�g���[x�F�xT<���r��<�(�>��{7�I=� ��՟p<�y�}�,G��JQ�  �s�R|>�DJ* R�HB�=�E_6��wcǌ�;�ҽdS�����W7�
���U�;���@Q�n��}�O6�c�@�/�"{�p �x����� P����
��4�^G� 9u�QOg lr���<�� u��� z{�Py�����@�ް:�{A�G weV   +�ޥ�*�UT�$@P��
e� 8� {����͍�A���� ݏ=��pp�M �c� }���:ݎ^���� s40���4���}'�q�
y\�mp���9���{ 9�w�t�y�S�� �� ;�@7g�ЛA�B(  wޥI 3ꠠPH���_l���2����@3���%�%d��k���-���&�Q�����`   �JR�p=��w��^=*����`<��oa���`���*��� w`��C@ ��Ϣ�H |J�T���Q�2�' �r@49 d� �p�����<�r7���-n h��A�b�  Ǥ�� pw�p�� �3� ���A�@2��^z�fxv t�d�"� y�  � @"��Ԡ(� 2&*J!��cI��`���J  �     D�2�R��2L�A��A� hс0��JD%EQ��&M1 ���OT�A����      $"OԒ�0 �"����@��G��������U�ß�?���`=y�<(����vC���� *�����
��("�ꂠ*�S����a�i��������������??�?�Ph?�RI$��� *������I��8�"
��������������&0q��bc���&11��Lbc�����0q��bc���&01���11�lL`����1���%�1��Lbc���c���&0q��L`�8��F01��4��b��11��\`����&0q��)�11�lLbc��&11�l�0q��Lbc���0p`c8�1��`c��Sbcؘ��&0q��`����&11��Lbc��F&11��L`���&0q��`�ؘ��01��$�1��bc���&11��Lalq�Lbc���0iƓ���&11��L`c܄�11��L`�1����3���`c��&01��!`�8��01��Lc$!�L`����.0q��11��L`�8����`�8��0q��LbS��&0q��`�8�bc���&0q��LbGbc���&11��`c�c����01��Lbc8��S���.0q��b��hq�lLbc�&01�lLbc8��&11��L`�8���11��bc���0�bc���&0q��q�bc��11��bc���c01��Lbc8��11��)��\`����&0q��
f11�lL`�8��11��1�Lbc8��01��1�b����01��Lbc#bc��11��bc��L`[��&11��`c��01��bcٌJbc[`S����&01��Lcc��01��bc��B1)�����&11�L�&0-��Lbc��0q�ČLbc���&0q���bc���11��Lb�#8��.11��L`����01��L`�8Ď48��1q��b�8���q��bc�Ƥ#�L`�1q��\bc
bc�6��0q��cc���&1q��`�8�����11��LbF��.11��\bc�c����11��`�8�0�.11��`�8�0`�8��&0q��`���.11��Lb������\bc���&0q���\`����0q��d`����&1q��\r�#��0q��`Ħc6��&1q��\`���Bb����&1q��bc#8��&1q��Lb�1�8��0q��L`��c�8�1��\b� �0a�H��.0q����)��q�[��1�l1�S� c)�$`�0�
��G$ ��q��0T���U1�HDS�H� �U1�0Q���`��q��1)�.0�(���� `��PrB 9!��HAb,b��Tq��1�(8�(�`)�q�11�0A��q�1Q�
8�(� \��1RHDG$ �� q�1�
��S�� ���1�!lT2B5!Lb��q�0�
��S"cL���1R���2B(��S
c b	�@q��1T��d�Q1��1�"��L`�`)� rB(���cLb��U1��1A� 8�S$"&10� 8�S*d� q��HAS*d�q��HA"�`�S`�Pq��1T�"�!Lb��q��H@G�rW��Lb#�@q��0T�(8���\`�`&0�*���cb)��
�� �1S�#8��&11��bc��0q��\`c8�ƚLbc�8��0q��L`����0q��b����F&0q��L`�8��11�L1��bc���1q��a�c8��&0q��`�8����0q��`c���&1q��\`c2B$bc���0q��Ka�J`�8��01��L`�LLbc���&0q��bc�c��01��Lbc8Ƥ&11�l`c���&11��Ld`c8��01��`�4�I�bc8��0q��a�c��t����r�y�|������M�x���!��� ǅ�1
؅)���͙�Ύ��a�ػ�R-Be�Éc.=0p�[�n��]�wj}.��i��7dYuf��V���f���m�c��Yw�Kz>��Ӥ�u%�.n���F�/�,�h7��!3��c�pm�b�I,N)7��+�Y�T�M͵�z��� �۝6�\4\�U�ݡ�ݪ����|�ͨ\���C-$�*U���.��g4 �i
�z�9wavO�ű��v5�=�����A���d������a�⻵�f�9���Ǝ����s����*AÀ;�����>9!���Q&>2���[(m��"��q��$£7�-�*b�9G)ݻ�ѽ݆����[����N��*<h4r(j
n�	��Z���u�;���7��+�;[�¾��Y�� �𶜧"r�ЇLi� ��#���7`לm�"�i�QG���jbL-�6PrZU�^v�!G�|�t-%����̐�7WgA��Nw����N�ς	KWno��3��$�:W��]�dW� 1�m���~6�Y.R�C;E%e�h<mw&�vP�pgcd�a�eH�G r�z�����S�5���O�rt2J�{p �X6#9�avJ�ݏ�v)�NhI��h��QHqC)Qo�W2�7(���c6ʴ�����>o�v8��㷒�l�^��PTN��ݔ���$����SƳ��9���҅kQ����ۃ���GLzB��v���������"���ʈ�����M\����pj,n�Y��}�r씺��Ug+�듄�+m �G5�*:�XP���Y.��\.���n�4�U����%��#��Y�'e�庾���%˷~{{�˃��{wx�	���Z5�3��d:�gN�y�N<�h��V�n�uӚ�⛷��C�F��Lqu�0�Xv������[�qp*;;�2�50-�R
Q�T'u\�ú7݀ IZIr�oj��T����G6wv�Yb�97-�L�)P��Zo%�v����l��=�WuѸ�q��!M@wL�������t�����-��F��9���$��nL��`ls��"�S+q����1
�`,����&��C<�N��g�Ͱsű(�j3z��wZ�o9�Wk�H�޶E}�Gwf�������{I�V[x4{D�ݪ[�M���w���g�M��Z9'b}�W`����KVi`���ވZAܰ�g(�p����q�B�zw���Hbt㓠Ǿ��r[��\�`d\;���,����������_���[ ��No�Ok[0w����9�����{t�z6��.�z�z��bO`#��q%�q�z<ܺ��N6X"���Hg(hvU��U�=��c��р�'�m�h�&L� m^f�|3tًZ�(G,�M��!p�[�B泳�ir��hS��w��Df�g�&�]}���԰F�U*5�ޛ�p�Ox\Ԕz]�p��\8��g5�Kǝ�%j��u�_��gZ�k�i썜�2;�n��ӹi�qKw�n��ɫ����f�y�l%�J*�ڟ�e��y��Lz(��-����&]*��37g�!1>���%Z&t+��`��p�t����)�¦��;&h�
�{ٸ��]�nL�5��:��&�ǒv�Hއ�;:�ݿ ���~X���lq%+�)ù��kx����sRqɹa����2Ц�soV׊A&�4�ƱB�p��<��tax��:q���:�9�5v�`�$�h�Ѓ8�ᲥIۼ�����`��unח��
�Q���-�tkK{���#a���]�.E��$G4E��:YE��嵿�"Q;�C��:�1�F=��}�t���a�,�ӝ�Q�6| 7�f#��u�>|bWq��4 ^3�Er>o�rr�v�0�.b'�$�d��������;wq+�[x%n�������&{#��T�A���k�-}��p�W"tt(�"Fs�����{b�)97�rn0��7�=��7�)�
��j1�SQO�ˊR0\1��V����&\�^����%WnnͲ���Ԅ�����[���Yk�;�h��M���f\���njw�F���h��M���j�2�=Kx��y�Q��q/��dܨ̂�.�����{ӝ7��Ļ�.Ql�7|�k�^�[0�=�~y��l�g�=�6�v�9o=�^֪cs������%�.{ë�i���J��_Љm�!Ћ0��n'���5�)�����H��E0�k<ݚ��%�l]u̗wX�dխY���ud�s�wN��4r�w�I28I�;f����v�BT�)��"��EjÀ0�9�Aկ��CQK%��;��Y��9Ob��3���C�l���;�Pׯ�NNp�r��ۋ7wїV7	�L�s6v�
\��S��W.��>�Wu ���L�ܜD1dd�	\Վ��B��>�:Uc;6�;�ygq�=��E������׿jp�]z7zv���>���73�.ɤ��M��ʴ���q��>������y�;�\�>��1�첁�����~Nr֭� ������V����Q����-� T�ؙռ�C�r�^�P�F̡Ӏ����TN�[�n������Sf�H�|V���W�n�܍�k7�+��g]����l�Zsb�kZֲ.����9?��iOoSy����9�2ʋJѧ����/�&�]ua�#�9ԄEG�lͷ�-���j���zu;R��Pa4�d�fp{E�u\�x(Z󵧇���^��{v=r�vt�4ϩ܏W�wl�7wTpW�&v����@ƣ��Ly���T0��������('53r���9u�����MɃyg_(5,�g�\yóN�.�@��dä��BG�n�����h�v�{;����v�\:"��1�gݼ�U��'M�ul�
%tл_b1])�Ᏽ��u��7�^D�w{������D�Y���҇ͯ����f����Ý��W;+���qG���t!K=���[sz�z0c���t�W�ݷu&[ ��cE�y�J����9�f��3��t��޷��G��$g���]o�+�4�nE S#c|�Ǡ�wcX��s=���0��b�&����'z�v�ӎ��e����S*@�ޥ�i.�z�Z�l�7Q�7mͺ�SV�ʌ��#m�s7�8jsFB��,zt�9r]����M<gӅ�4Ŝ0�[�Ow�~���yn�H�b:�%Kq����=�.&@L���G[�$/L?�������QL�R֎`��/�Cv�NQ7�^��g>2N͕gc',S�Z3W+V���o�pp��&m����v��5<��+�ѳ�΂�	�C6����e�R�R��_)t�>���rwc��p��Vho���!ؗm�0�Of5Vu����+vw-�3�����"o�d��������w���i��ͻ�&T�S
r���ݏP�%�g`z;�����p'f�����N��]kr��Ʉ��\Z���U���4�a�"wi#XA�N�$�8�����{.O5|���͠�b�~�
�!�W�y�Tr��;D6tD����d��:���v+t���Ҽ|Pk���9B�n:A��dbu��eF���t93V�.u(dI��9���0� vB�Y4u|��\̚Rd�v=�L�^���뚡���Z���:��p�95-������*s�]��;�q1K$��V-˒>U�����Y�Uk|���0���*dO%mp��*�����u�x��Ε�7P�#��`�K2��z4
����Q�����^�̔��wS˪�"���s���I���VoD*�WSc�OP�`Q���+4�o�]���nr�[(o=ݥd᩾�S�@|��l
��u�/]�i̽�t<��^�᫇����B)�F��w5l"�m/�>y���Bv�
�˻u΀���8�̪��X\\�p�i��w9<[ݭ�F��B+gJ#��I ��t�ŝ�S�w�>�X�ɻt�,�%`�2��*Rж沍�qH�Fón��aA�)ٷfV��\2�נٻy���a��ۇf>k�؄T�����1d�¹)[%Y1�!��w#��� �xC��9�/-�)!a.m�3z�ˆ�Q��PY+�2�FD v���]�Wl��˸g|��U�C�0 )'C6��3�tBFUܰl� �a^�̠$]åUg^&�9ܗ(����@Vܙ(e�cy���ú,%�Bd��+���3Kx�#��7��h��:[c$\�A�9bCPK��nRn�E�[�E�Tޕ �`Èt����8�@�����,���M[���vI:���G����:��ҹtP��˽3��a��. ��Bμ!���=���w,�GU�5�.7Dw�;s�N3qh�W`�.��k0r�u>�&��OO�;��"��cޗ�[��}�L���Җ(��86,�ש�U䯋
�v�f`hq�)�P
UM9�F ����St\y������U���d(��CKsh�L����Bͫ� 7\

�<4�x['7WpՇ_�?L�u���Q_3�T�`��S+m�u>�ъ�wc#락p�3u)�q 6j��a��wG�AP�+ބ�fo7�����B+�C�"��o.ζ,M57)C���]�� T���X��p�sz-�V2�l���0dҎN��o6���bm���U������9Q!�O�Ό�]�}�c��7A�I�s�����܀��p�[>oh�1���n/�)���>�	�{�⯇gs�*Y�[	E�T:	�����S��ΆP\\u�<&�L�����a0|�׼�պPh}��x`z1�{���g4�,<��8N��C�٫S����4�+�qn����h�������?.���s�n��w�9v9Y��bӈlZ��d���rӭ���Dk��`{��N%>f�Hsf1�.��l�6MՎ`n��Q˨���Ɏ8��V��ֺG�DI݄ݥN��MMe��$zk����`n�{����wA��Q�yl��i�2�����8�K8��O�J1��f�v�X�]6��<={ni��1-1l\8�S���ؚ��¹'+Y~.2�9�`L8�0���3��=���`2b΀9��nB
�|8s��g��k�:>�;iK{c��fL��f�V���n��C�i��l���;�v�b�~˃6v&�-��������QyPA�.?�P�v��x5��IN�g7���{J��u��2Lף��b�����j���qQv�w���z8�d��i�{�.�s4�1�nH;:�	�/��ݮ�į�2=�:Ў`ZgӸ��J�������M-VZ ���x`��={�>�ziC/��M%>�u�K'e�;�t�I�;���Jt�t0�������z� ��0@< <	o���l5��d�t�^ �dR�l]@�^�>z����R;&�I4�.��.�L~{����
���̯�3��H��t�� �At���<��O��.����%/m�x�zN�H�6�i8'I$���5��{���*�H�~p�I�0�QǄ��/l�f���w�t�=��/�.�ٲ�K�·��=߻�0 �C�zY|�w�=:d�⥋��� $�|J%I�a,�^�I�k�;Od�k�\�~M'Id�pN��;q�o����g�!Le�(��T&�t���mp�&�I���OO�,�#�E��w�Y@�y;���|�@�I���C>�l�I&ǰL��&����}?�&�	�I$�J/Œt���I��X�����]K�q$�N�+�U�j���"W�eOp�ĒQ$�:M��Q���a<gK$�4���{��i�(_��M# ���g�D�$�"u��$O�s��=�`�}� | `�٧��������~��/�~w ���N�v9IDR4���
�����<܇�[�	}G�z_��	��Ot����'ĳ<^	$�x�M2J�Y(�N��u�d5����i<^�Q8'�O����Y>$��{:k�t  ��3���w��Rt�K���L'I�4�L'u�g���K���2�`ݷ�E��I�aU�O����/��O�yRT$�e��x�M�t�%��0���x�H⡺n�I��:摥RQ(�'c����QŜ�R��ϋ�L�1��%x�-���Q<J%%S�b>�BI4�/�d5�OEW۩��x�&���,�M$��'k�[�*%���ǯQ$�T<ϑ�w�i�*�t R*���x�?)4�}Jb�x��}��ԊI%��8�V��i&�
����qH��K�Y\^I' 4��Q���c�-@} �/�7��g�Vz^'I��%f�x&���:T�B�KB�<�t�p,I$�x�I;Sp	�1���/�x{��z �c���*�E&��W/�3㴿�|K=K�a������g����w��L� z   �)4�N I��x�`��a�{�"i:K%�He`�M�=ſv�%�?#�/�~��e�+��[,ey�����[� م=�K<N�	�i8��I,�"F�y>$��N����	$���i�I��n!'��i}f7�!�>���T���<�zoCГ	L�w��:�I$��v��x�C }�y�=�t ���C������%Q�B[�,�5�̤�0F�	���,^nڮT�3���SY^��	��������Ż����m��z}���"� 2 jحj��EZ���UkF�bִm�QU�Z�j�[k����Em�-��تѶ�EXڪ-b�b�j��k�F��֍���UV*��U�l[U�Z-%�Fխ�Xմkk%mlj����*�ƣm�kQZ�m�+XմZ*Պ����F��k[EV���Ū�j6�FգmZ����Z֨��Z��[�Q�[ZƵ���Uj�1��b�_�Z�����m/���_�O��y�^Q���m"�y*v��Q/�>BD�2����W� 6�'{w�)؝˿,�j<XY�j�@� �4��KRrQ>�&l;=�J���w[ M����@j�lE�L��v<�����'�������3��l��d���j�Q��/>A/)C9� ϛW�H\<�9v%rP�|�r`D;ǰO'n�{6w�ὤO"%���U*�(ߒp��y �B�o0."�'ʒv�2��y;�˔�I^g���.0�Z�%��; j���v��������
�� � U��8�]��t�ʹ��3��� v|����2|� >F�Q��r#� rU��/��)�� AZ�zf|�V�qE �'b���!r��jzG�M��<���( �������`  "~��B{�~t�?�}<?ye���?�����?������������ӑ�t��noo�Х��y�~�0{�2K4�������]�M��(�u{�b;��y����Q�A��Pgf�9{�8=�E��ӃJ�9�DZW����U>^8Z��`�=��~�ۯ\lٖ11r�g-9�R^���k[SW�xK��X�2��sǫ	��~�z�J��o�NПeO9�Z[�fb��i��l#�w�����5��qC��ڹ��x�d~�y�+�i���i��n�Mf��j�rO"۫4��n�:ƙ6-�(�;�f���AB=Aq�Ӛ�b� ���N�����sv��EhWp�0o�]�|�f��;����=�6�`u�1�y6�s���F��=f�A�ݠ�=�&��6dc����F�i1������w 3M7o�@������l�n;O��5k�*��œT��Ae� M�Q}
������e�Oyv�,��Rٌ�˚���nm� �[4p^:w����GϞ��V�A��_<^�Iqw	���)�t+�3�::啫�ViI"v�p�AQX\�#:�c����
c����_��d�d��ӯ_u�_u���]u�]|tu�]u�]u�G]u�]u�_���]u�]z뮶뮺�u�\u�]u�]|u֝u�]u׮��n�뮺��]u�]u�]x뮺㮺�n�뮺��]i�]u׎�ӣ��뮺��X뮺뮽u�[u�]m�]u�^��u��u�G]u�]u�]tu�]u�]u�]u�]u�]u��]u�]u�]z뮴뮺뮾:�:뮺믎��N�뮺����HN]|6�^]��tK2�y=�{蔄�3�@���]AٲL�ۯ7���`�۵�YӍ��;&n)�78�E�fR��X�O)�|~ɑ��o�Ӿ��5U?o7�\nt�L��׷��p�X���g�ޤ��7v��K�߅ԯ��������,��{"3"|��~ܫf�@ �6cS٧Ѳ��ú���{��vx�`�#]�y��!p���`u�� �/V��,Yyty3��G`λw�>Yuw=]�>�za�w`�ߡ��ÃY��o�ν~��j@�KʏC�"�`��ڎ��Sظ��/o!�TG��{6�iȣ!P�R��/�ʬ#��ng"t�
|�䷩o=y�>�wE���y%i��Y��8vJ���{DB��Z��$���������}#=�{]�y��^�i�z9s.p�LWk	�7�/�p#�<H��0���r��a�opЯ���åƗ�����-��j����qa"Cj8��<q�t��f�>0{'�9f����W�#Þ��N��ٸ�����Z� �F`D�]����xW����%��U����ɉ��.c�F����3ݡ��|���|x���׏�]u�]u�\u�]u㮺�n�뮺��]i�]u�]|i��]u�_u��u�]u�_u�]u�]u�]tu�]u�]u��u�]u�_u�]u�]u��]i�]u�]z뮶뮺뎺뮼u�Zu�]u�_u�]u�_뭺뮺��]u�u֝m��u�]i�]u�]|u�]m�]u�^�뮺��]u�u�]u㮺뎺뮸뮺��]u�]x뮺㮺�ccy����S�,+)��%�Րl+�h/틯���xYY<6�*�'�y{����'ފ��9��w� F>�����07@֕�r��9��y(�>7�\p�c�k��6�I�B	��OU7��!H�>������N^�[��(���E���{��3�%S�6v=��4��Mu�"�-;��Z|���wܳV��K�v�qxG���c�'����'}��כ�8���+w76�i�p�	Ӟ��ޙ/�]��{t�����,<a'�7�1+PM95�܅���F/{/��n�����L:�)[Xq%n�:7��s��!��ӞD�9�S����H���؟t�Zك�FJ�G8�={5g���HԴz=>\I�C�`7q7�gt��x�x|B=z@5ٛ�y����`���ዶ�s.=J$S����:���n���&������(���LwU�����G[�I�t���b˕��G���3��z�3��Vn���!�by����&���g�����N����8�s���>㽢l+ *5�9�<G�9#�g���ga;�u��ڤ�>?���~?|u֝u�]u׮��n�뮺��]u�]u�\u�]u㮺�n�뮺���]u�]u�]u��Zu�]u��]u�]u�]u�]u�]u��]u�]u�]u�]u�_u�]u�]u뮺ۮ��n�뮺��X뮺뮺�tu�]u�]|u֝u�[~8㎸뮺�u�\u�]u�^�뭺뮺뮺�u��뮺믎�Ӯ�뮺�㮴뮺뮺��:뮺뮾:�&wɛ�F�[뛻��p����d>8˅��ӱ�.��q`����1�v�w�`{Q���%���V�.1�\�\�����O���q5��6=z.��L�A��i��}M�\����q�=ގ�q#����.�z�f���`d�q�bXb���O$|ۆ1��t����dh���>���]���:��<2��g��˩.;��V{���l^Ͼ���s6Pv�i�X����l�V߳{۞�f���J�w��5���3z�����K��D�hkD Q�Wj%�f��H�d�T2VO���|	T�����4��o�ǫ��G�|����<<��r~���{݂^��r�g_{�	�����I���ZG���n�;*3��{@ýZ�{��8_��6
PcYA����<��r ��^+��K�٣,zI^��pn��v/}ښ��v�{zv�Hk#9�P�>�gK��H�[�nz�3��-[�=&�$���Gc\�M�z�<
�˫E��^�纆B�� ��e��m��B!<D�x�r��qe����0[82�%��q]팜��y������G��7�Dي�]�B��e,�4���;��W��E�/"g	�\�>�+s=<g�3��of�2�W}��q���_~:뮺:뮺뮺�u��뮺믎�Ӯ�뮺��]m�]u�^:뮸뮺ۮ�뮽u�]m�]u�^�뮶뮺�]u֝u�]u��]ti�]u�]|u�:뮺뮿u�]u�]~:�]u�]u뮺ۮ��n�뮺��X뮺뮺�tu�]m�ߎ:Ӯ�뮺�㮴뮺뮺뮎�뮺뮺�뮺뮺뮎�뮺뮺�뮺뮺뮎�뮺�s�.�^O2N�q�]T.y��}�N��W�/`����U�K��e�s���P�7x#��,��~>|�c��.L���^]���G9��E��e�;pX>J�g>��|���[��
�Ɇ�	�'��'!s���sx��A���/ ג=��@s?r'g�@0�����t��7�
���;}3�Ͼ���ox�vF� Rr����|��N &�4�D����S�O3֭��dY������t��E�+�{�'f�L�|N�Mm,h¼��g��6��S�b��5��}��a@2�g
�����􎞅��{<��þ��D���؟����:3jfB�����3H���T����y����g���'E�~�>���-9�r����g��H����6��g�� �%��!��!����^W<�����{��|[�inE�~��ʬ�`��z�Ywjs��X���k�4�����M���q��5��x�Z��F,�Dr����p�_{���>�>8#(F]9"1�Wxb�؉�S�e�Ԑ3*�q6�R9�Y���6�9���`�7����2"���y�@���W��S]���Dy�`���t?P�r���~�y�{6wG�}�afz�f*s}���I�f���	�|LŲ�\��m�2�R�ñƸ줨yn���]^f}�'�/��0t(�V~Nn�Z��n���T��ԅ�s/�wq $Yà��Z��R��}��0|l�p���_���z2l%��剈c�����z=��<<3��t���5ܗ�}��%˯����{��b~��_o�J?2�LY��Zܴ����|ov��l]3��X��"*�k%z3sUDJ\��9�����e��3uk��z�&�֋s�S�{ϣ_g�/,�XM����w�=��rRT�=�����U�H���y��������{���U�\O�;����+��h"{�D�;�[�h�{pK���=0�3��n�� �,�yu᣻��Ks�x�N?i~�.��d��{z��#�%�30����M� zy�o`������Ԥ�\�(>�=n��x��k�/9��s����~��r�G�Kw�~��:?u��|}t�]~��
�=ƴ$ϒ��n�"�������������L�p]�`�sS��18*�[<2"�oxnU�o�\�g�\�-�ia�'���{��t���bx-{��nO|^y���2�=ˌg���>�������⎛�[14}7�T�Z6p�}����9�[��������;��yޡن�)��X�+�X8@dY�)HQ�b����=9�O��V��ɟe�2��31���s��x$suϓ��tsկ}t{޹�,�Uf��Dt_H=u���#�4#<���E�p�g�+��L�$<+Xn=��n\��=���f�2Y>x(�@���w����~�y�̊n5��|__d�q�J�w�ONhf��а��v� �8&�I�|����ҹ�!ٌx(=((��1�1%L>��</k�|j���=�{gy�ږ7qo��{�������n�q����"����/�m�Cm�Ao�μn!�E�]�(�4�V	ټ�|�c�&�=�ۈ�M%���W�f>R��)�y�����|&�|���>ff˫3"�)i��/�_��h�v�7�8Ǜ��F:�ܙa�2����%�g�r�����Z=ue3�ߵ�������bnW�=^�#�<�m��	���]�	�B�YO�<t��;�fׁ�����&��������`x��%���Eb�5�L��R
j�'�,��)�]��W�����}ݯK��Uv����!ps�=-uq�$ʽ��.W��>���g��_)��c'|�\��>����}������;�m�r{a��G�����)��,�0H6�Uvo����������0VORw=SW��n������O���D��;�qK��������v�Qa�\2z�{V���:P1�Ig��vd�M��MۛMꉛa�܅�5�di龊y�^�p<����	��.�}����2t�*�s�K���;!͗ݤ�E�y&rU����ћ��\�4&�P0�����t�Ǔ��?��6����ɐw�\�`P̃.��Yx��P��x�&Xxi<x�"g���j�;�����V�X����1��cqc�����\��g�z��n�`����˶_D�U+���s����Y�T�[a��g���L��J��͹���W�zWa��%9vX�����C
��0�Ņ'�vJC/е���P��e�-ۗ� �0���I��&濾��O�J�7NlԒ��юaLzL�$�%ݛ��R�M&�߅Y���b��A*�k�:�s�ˊ�Ρ��su
.��4f���5C��s�4���w4�t��^����ݭyxi��������q���C�|��sJ�}1C�yu�_OV�2v茷&$��(�,�6{x���\M*�F�ub���S��q�
�;�%���ߘ�Ǐ'�����v�{$�c/V������p&��=�oe�oӾ��l���[⟲�Dϧ�y痳����}z���C9��A��Շ�\�s��W�������輕�o{�>�����/q��M{����v�BF��]g�&{Ĺ��vW���}ϵ�ʌ���q���_I�yU�;ab�ou�ߚsd';�Qӕq{�����ޝ�=�r��$h�vI��{ݓ�J�=�T2F&������D��8o!ϖ�\���Ob6�6{�t�ΡR=/zl�4ʸ��)������C�$�g:���`s�\;�ߏ��ɾ�gnȵ���G���z����I͆�e*w�`�>V�Nlw48,��U��U���q}���>������۝}�ް�X�7�%�ݞl^@g�_��υ���R�9�d
-��-��^yvj�؏�1�yp�=�q�����Ȝ����X1
��j/%�׀>�A=M���E�Ũ{��n���9���2�����d����W�/�G+ПP�dC�ݳFL|����	
fw��ՠ�}7q��������F=���O�����	��t�+�+s\�L$�EpV3M}y��^�Þ��;�B���2+3�~�GM�h8a��^m#t�C�������C]�g��#�{�l�E��\���:�+�<���tv͒���⦜��ܸQi�/xu[�<3ܻ�x�)��$L�ni�:��f��U�;��H���{���1ۣ�9��oY&ކ�V�nU�q����F0�EGF{�{���c��f���=���d�-�L�ޭ������K���Au��3�����J�%��[��FL}�y�>��<��;��A~�$����s��������>@�J�����8��r�f�{#��z��r�|{$�˾���U��
������XH-*�*�������	���5!��=y2�scD�
��3 �0�7���y�d=��x�gM�kn�h��c���-�-� m�:|�!��DKY���M(�[���D�Ro�=��{`��ZI�@M�Hk<��Q��}/r���J��CBƃ��IkĊ���h~��O���>]�9��=�X��%����f�|}�ێ��#�E\^���&]]�Qk��[����v�G�{�ɧŐhJ�{&����轗^����n�-�q{6]��_�z!�Ոi^^c��ѫ�v�z���$8BC>v��yU�g��~�W����?�~����迈#���RO��yY�rd�\��\�/6����s�?k]v�G��	�YQ��h$���w���X�3n���s��E��Bt��s��6�(�Km����ܝe�8�R�t���[�~���w.�kz�5�F���gs�	���=�xw�����K�\�a��zu��l4�ҕ���w�4L��u6��Hi�5���Ke��׽;�s
\�[g�ܫ�������qk7PХ��X$��ӻ�4N��k�Yf�l2�qo����z�A��������v��)��Ĕ8H��kii������v3[m
��3�x#.�we���gF^d�\hE`ǂ�P�l��ÐKh�X�S�W����ݭ���q�lo��u�d,P�[��|w�7)l:�n�ۉp\P���rP3XG۷�\��Ռ=N�۩��^�8�{����:�e�퓎6�S:C��������nQ4mn[i�a�&��u5���v<���E�7M$�m���]`c<���ۣ]��E�����[��Wo<یl��p)@�ѭ�G�{{-�;1�&�lMbC�JCs���!�O�u��ɇ2���I��Ycp�E��H�X�k*�\P��.IAc�Y�,�N�u�:ʇW�ZM���v��!�-�9V�z脫F�lZ�!�5U.���3f�LJ��sʞ�ۢp�7QŔ9ϢC�݉�ó��� dQ���@�e��K �#Zb̺j/�{;lr[1OX�b��u�rv�����M���r�iÔ�a��z݇SQt��4�m)�,Ĭk]C&腫.�<����k	�g���H��j�5=�{�npY��M�A�9A��4��4[���;ke.��ɶ$4�m[c�)h���kɎ��^Y�Y�7u�L��xTg�:�u!^�����e͈G^�m��F��� 8��4&��,�\T`�k/m��i�:��gr�v��Au�P�X�ueqí�9<3�-�g2l��;Ɗ-�@���9HGE�g��c����9�nqn:뭲��8TF�k�c�uH�uḱ����R7���N�bz0�N�YwZ��Yct��F!�n��)(ĭr)�1tf���1��	ap�'z㽮��R;YZVj	3f�-6�nl��#�e����ntģ�e��1�\{sĸ.$s�D���<esl�����"x����@�5��z�)�7����|�v񫅌����ʪ�N&�wl�4Q��b&����� y�]nzz�瞸V�l����t/�����cy64���[���b�5Ŭ����6�4!�l�VS	�ڎyRL�ý��gn%R]���÷U���[��q�l}����a;[���ns㐌�;�������Лm� ��KJ�b1Ĳ۔ɬ�0��7gpR�����u� ���+j�\�6�g�	k5�j1����b����2�G�e���*���r����#n�/[�"^��v�sA���u����m��u� p�>��Ӗ�c�c.�����;��sv��c�T--C]e8p]t�P^���|�{t�k۰w^/=v.�\�Ϯ�^rWI���;��۞�]�v���h�d����K��q��N�3�q��auѥ=m��,s��S�1s
	�`�]�[T�5[��PŲ�i���4��x��ʥ�G`$]ab�`uM��-qM�b�kvL:�tsOX�S����ݶ�Ov��f-tv�%4L�3n��g����R��8�ۖ;]ю�уn�q������_5��|�iOE����M۰<��q�:�7n]ڳ�=��N홁�u��A�G[���Ct�:�g�eT��6���m������r�qY��-=��2skp,z��5��=`s�1ۭՋpj����9��vY]���L@r��P��1cMuBk�;��s���kf�*������78 9����n������-�9z�`�'ij�Y�v�S����V���v9v��r`���+Y�rȷ��.�˪���\�'m��8bږ���-��τ�uI�L��>���O��v�Ѱ=�(sdoT퓍�.��Y=�F������;lk.��MC��e4�U�ŉf�,2����X"�+��'���)���w[՚|@9t�.�����Y8����n�d�7��<9�rMukO[�0vwT�79#q�f�^������m�z��=���&]��hCGS�T֬%[[�kф�hⶹ8�m�N}2�@�d���ݢ��,�9_=�9������]Z�s���t�I��5�&���a���wt�,����į�ˁ(�{�t��v�ݍ��'��q�M���n��a�m�U�xUQL#k��4A�j��Ů������� �{+�q�e�c'D��z�:����=u6뵧\��ۍ敫�����ݩs;t��՚緉q���x@{�wi�Z�M�A�� �<�u�.w/]q���2�'��<��Pa.����f�{@3��4MLDt�h�����@ʚQ4um4%�cF³5��ztN�ɦ&"��\X�B���񆺜�0�
��%�KZ�k��C�A�q5�;hYIf�Y�KH�����ahtQМ$��rC��պ.m�nn���踅�u{l�F댢�������i��t��6 x�!GY6�k��mr����$�	�h��5ӡ�m��f.�{s��1[V�-���U�۲�݈��6X&Lʕ���Z��u0m����f$n��:��X����Ճ,�Pfd�]��y�i�Mۭ���{��ǋ���z��������n���]oF��f��+h
8�%���ejV��#�0�&1��fd�cRj��һM��cB�`f���h�.��R�;���!�d��뭭�lg@�8fW ������(�-2q��k�<���Ƣq��F뇮�n������Gp��),���άǅ+��2�f�X[��*7SWA��;i���� +���͉J���k6�H�ڙ՜�N�U�g^3���k�%ڃLtCi8퐎�g�܂����Ҳ� {p�T�-^
�&���Q�w�
4�7�0��+q�e)m|3n;�ὄ�����z�Q���8�lۣ��e}�U�f����X��kg�^�;(��	Uք�����y@\��P1,"g�eU�٠����a������Gh�\��*&f�qc,�n���ɞ؞�/<���;'&��I{��L;]U��8�����}s�F���p�M��pƩ�4+4��I���(�J�4s�N���}�����T6˞j����9�]w���{�=�lf��۱�M/l��1��1v^�l��ݮGa�M4��#��i5���e�.2��gg���=�J�c�u(�����8��]�q>'J�̴f�p6���*�uT��u�$���l�$�xhq��=rvWJ�y�瀃ji�j�/��A�k��92'6�a,R[�Y�D�g֗��:�[[rsn���Zx�7[�ݡ4���ۺx��a�d�ê�l�9�V&5��S��=vx�{c�-�.��bSB�:F1���t��m�h30Iv&�q�on8]�Km����f�N,5'5��kl6,^	f�S��9.P�^��4���XK.�Һ!
�Ѧ-e�gx�K�M�3m�z�m�����ו�$�я#��2ڸێ��8��o\`<�[v�;�^:�e�g�7]�(:�VQx��GgFWWnv5f��7N�`�Rjw+��(](�g�ϊ��g �)��'D4[�a���q�8��,d4�j6:Vf����2��.0�ޱ��ZHk)��8��",�|�]'�u�qE��j�J�R85�i�!^���l��<�w_}����i�2]�u��9Y��Φ맨t"n��wQ%v��W݌�v�p$�'F�y; c��d.��vQ�m˅��b��1�C6nT�6�Ga.���G������l����{[���=WYYMςB�J�]��g�S��M���Z�|ϫcb@ ڝ�:iú�;��=�Q�y��d0Rn�i�<� M�!�	��YDynm��f�R�7d�*��e5����n�S���:���y�ι!�����s]��&�W�6�w=rލ�&��m�uq�m�`�����t��x`�{Fn����k�����y�#+����
	0�j�v�lIu㌸[���T=7�\x�-��[��EӶ�֖�$�ug[b,�lq�qeq��S
��s��s]���2H����an���cj᪪����UUcT,s2���z��UST�UUUJ�UUUQ�7e���e�i����DԸ��>�7��C1\c�͍ѩ�c]u�ed�vh6,[/L�a����:�;n���C�U��?Ǒ������.�ڲ�&�LQ��W�1��K�e!]��Aiap>{knZ�q���]��#.$e�e�֨ە�)bLb	�c�ּ���,,�����"M�$9�vl q����>5�Bg��z���)ݥ��R�͐\:�MAn������[H$���2�Y1�_q�v�=0�L�)R�_����Ԗ5ܱ�fP�Q���o����x�:wPvP�������^B"Y���N�#�����Xf `��
2�c\�[n�3s��N�p^PI��	*��;��\���jK�X�3*���!�ӛ7������b�x)��}�:^œ(nH�Cia��V$��1��9Ѳ�;,�cڱ��\g4V4�kn�8����m�m�2��yeK@���y��D�eͼ�u��^���6�t!KcL�j����Gm��pg���4�/{��Av]T ����t.#����e�kӫf8�T<$���?ue���ƫmC�W���_�&�l�8<B�.�̦��`i�Z�v{#l�='$h1=��^���Ќ�؊3-�Q����=��-�z�{�;��<n�܋L�#TQ�$T��$ bz1��_u�G]u�]x��Ǐu� ��$��]�H�!�BF2�Ki�]z뮺�뮺�<x�㮿>R�2I$�#!!��!i��EQ$����-CF4��^�:뮎�뮺��Ǐ:��Đ�a���H&���ղ�j�ô\�N����8���[͚^)A	H�F6������뮎�뮺��Ǐ:��'�T��I�d�"�3��;m#���th5�v蓚��kn��v�n�&�^92��E6��2D�s��Z<��5�$���t�K��ܹ�@��v7�r+X������r�8mh����w����\��uE�N;�;��[!��1�����vr�t775��wK���I
D�+��9���	P��۠S]��D�9�h�ǋ6y�]݇wl�ݮk�N�u��ݨ��x�Σr�7su���p�]��f��N_N'׫����`ѹw����������ywc�cQj4X1���m���x�&����~9Fߍ�+�\�1�������̿z��b�k��{M͊����+�d�Ư���o��w����a�����vG�(S��ݏ���o�� >˕�v6,{ҸG�����{��:����n�ݛ�u���r�m�2=<q�ϳs-�b��i�g��n�{����PY�j�͔˛��z�U���3��'*X���n��6�����S��0.�"�\[��=q��=f噃��1q��Y^���a��M��evv�CkT��6�ط���<�=n�|�7rѴ�ݷ]ܝp1\���z�ی�=�ol��ZmK��������@t#���"��n��x��/h�㊪{��r�Q�G\x�n���M��v�����i�۟S��+<��d^�8v)�y�ۑ�ܼ5Űnإ{n���ۦ���]����Zn(jn���i�&���	J�]�"���[��E"x�c)1۵tq�m���ɶ��%�ˊ1�<%��G�E��u����\����{�{0掗`�`��h�拴E����	{/\�m�{���В�v�ζmЏo9�8�2oU�`�';l����s��2snb��//e�Won1H�6t�Cg�uێ;Wn+�T��(��H�]��n�������u�sڬ&�mR�� �PBl�KCu˶�t]cخ ���ѪJx�-�l4��l�q�� �IF��4����sհ���d;�s/oA�9�i����ڌ�&G[� u��{�s��.���:{*vn�u�7��Bֺ�id�{��)�d��f��]��VT�}j.
6�'2tdB�nkn6�O2t�mջ��8}�G�^�m��pXas�SL�gup�kc2k8s�y���kP�D�@���`�U4�5*�n���m�碷��:�=`t���vf^��Rm�0�v۸��a���ssj �¬��v:��K��ʖj�b����c����)$�`jM���A�w�Lnx�X��vM૮�����0�]ߏ<xb�`2���Єy��ʇ"����a�ߌ�%`��!m�[Z����Ⱡ*�
���jF
<9j[R���D�h5,#+�+e���,i+H���e+Ť@�Umlm�K+-*
Ġ2�֕�e%�E�x�Z�k	J��	FF6H�H%���TEo����������YK� �@Ł���S�w^R۹���G	M&He���Pf�8�.65P�F��6�%��e�O�׭y�ᖏ�O}�:7w�v���22\<������MZ픛�A�&P�<�b�[����&�Y&�f�cfT�e��4�kn�@�^��bJ�VюӉ���_�c�`�w~�����������{s3!�����>w���lj����/���ʂـ;L�^����u�;hm8�ў�	�;E�Ʃ�fګ�UU3��~;���3꛸ݩSYuO�i4�d�RL*��>#*�]7}����MHW����ã�$Q�Z����gp-����*B���qrH7�ww�t/h7��c�ĵ��� ���ֽ�@n�2�9j������{t�ߞ��O{б5�˺��{2��v���~^�v�D_,S{���H��*o`�^�ŋb2j$(v��,X���m�����U`�3�l:ճ�&s��sf�k�tFۍ�p��)�FH��`Vmf��Wn���K�T�^T����q�*�b۾o&��5��N�oS��-��gf��H�[	�L���;�Ygsc!�E�ܦ�>��=뀦�@߹.ӛ�-9������_���,�A���59��j6j�߫,�˝�V�z�3�k�ڢ���I�!�:d��.p�;h��7N����]v`�"g�-@�J�� �j���e6I�\����˯5F���yYB�U�O��	�����o�6���h�3堫q��}�Y��;����F��i>��Wٞ�y��r�2�α�̫��*�f�k'D"�On�S^�O˃Ŕe�^����2�;�@/mIo��?<Kz���
ϙ�>w"x�1�`��	!�*���M��˵��k:թ� Bey����k���m����ٞ�tHr�g_s��C��}�M0����T�(�y{���0ȩ�̽z.*�u�SX�_F��|S3XQRc�	;QL�7���M�틌�L[>�O�,m���V���Z �."��hǎ���F;f�����o���r+e�ڪZ���s�ks�%��R�ŀ���H���ּ�%�L�3�,Ŗ�s'���Y������u~a�km4��֫Ӭ��c�j0=Z�be%����g_H"�pq��~�f���u��)r��i� �K�c7j0��7VNn�ў�����k��+	z���'s�ez�@^��������c4c����x��\��sb�g�u�����﹑��wV�X��Y Ir�
"
KX� �bŀ�}�!�z�o-��z�z���g�9q�F*��n顱*�{�������O��=߾� �r�1tī�fzz�e��mڃt������ƍC��<����!τ��ɺw������7ت/SaצZ7�l�L-��9@{��� 8���ݵ�o	5{�crq�~�ў�CE�iD��*��x�����Ҵ�~2>B�-�z��\>Yb)	(��ן���{u���Ӈ�dq<���v�p���cd=(�𧱑��.�ث��'Ȁ�F�ԯ�߽ŧ̚R11S>V3����ۗ��)�~���
�mض:���啛zv?�1K�z{�C7�a��OǖY=X����.�p���'�%�[��d�P��SI�ڳ�p�÷�C����b��|�1|nH%�� �|��E?O�����<Լ�y6p4Қ��U�כ��P�B�r�� cY���.%�o4�`v�kt/gt�5sRa�1%r� �c���^6�un2�'[�����;c�=�^ͬ�B�����[�s�s�(�meS���ַ�N. ]��ҡ�v�1=g��\<p�K�v5���0�Sl6=��ڍ��ۀ�*lJp�"������M��E��@�tyf�+�7!��(P��m�6P��_7_}���tŲ���o����7je]T2���f��FG�{�]�ykm����P��d�!E�-�S����V�-��؉!D&^_GD�;{�����ޑ��H�}�w{��RV�z����/׃2��XY������ti��9��/�ھ�|��"����~�*ɺ{&։|"=zg�E���K9����+�A�"�UW��S8ع5����z��j�r�[�5j�ر*��}�����K��(m���@lp̫`�*�&؄ٔ�����崡�nfx���ʜx��ўZ�Iܯ�ϐ��!r�_��v�������L�E>$E)D)��P۫7�Ϧ2t�s�=��7��k�[��w�#�eA�YjM��	�*0E�(Ϳ�`��-�F!������2gwߙ{��{��V�^��^L�b/���zf�fI�AB�u�$�?����~���[{�W�!�'�1oJ*|'r��&�5
.Zcw=B�+"�d��U��驻��Lf�	!6˱L�В�<���JUYf��J���VfE��o7N=Z�i���,�O���K��HO�06V���4z�v6룭Un�2J�\�δ�e������
����o���u^��b���T��9Q����9p6�&�l�j�~s|w�,��۸�����V(��ѕZX��Aؐ��h���7w6�~Y����T�𭯿y�'B�-�b�	��J8,`5F�:�k�y�1�ދ��k��op3���{����O=ߜ�(���#�0Rv��,��9�e��r�3n/�췫�V��.�T�2'YU Z7�^=�M��D��>�V�f�ܾ����ཀྵJA�/�2k}#�ڇ��\K̦2��Oj�br��/(�D�ј�z�������fV8��"$K�(9s��l��mۈJ�u��`�!\SV��ug��Ǟ�ڃ�>yֻ�<3�7n7�췫�V݋��p��_�G�X �@E��Z��o[�t���Z��z|��j�#�޾R���`�ݙ��&~�1|~ݮ�J[���^��N2�pR{���E��FI�e
g�����:�� ���L2qNr+n���e�]��S^(mV��6�۹J��<s&w�A��[����t�o�y=�PAq�{<��_nj��t�TF��4�FU(E_���Cq�,X�,`	��	�2�&gG��]���b�d욉ȫe���v��'ʶ�mJC��ϤJߚ��me��w��\�l�d�Ң;YJ3:f���9��;��!��xM=��w��j��cZx��3��y��"};�>�����"���襁��ܫz���g�/�}#�`gPY;�>�}g���$�w��=<��-|>m��1��~y*�ާ�l������q���*6�Ue�ؓ�6 � �B���	���X�їz�6k�j���׼�?������v�A�9b�VN�4�j����Ϯv�]�U�[<��\	����<auPfr/b�����_���{ ^x.y)E�/��T�;QH��j�O~y����y8�ԅ�����ys�Ǐ�����۲�1bŋ :��=��u�LS��E��~����8X�l	��:�1�=�1��g|w�\�th}tx����6�]��a1�hM���"�.�8��y�7]��L�u����`X��P��ͻ=��c㞣�����Ka�>���޽r5�"n:��}��\l�������K�[�nF$�K4r�8˂��k�#����6�Q�����~����?��|n�=�*w�s!/J�:�{N����.�>�q̋k�Pf��"-Cnݼ��)Z��F�ۆ�C����*!�<��yc��}��;�S>4g�g���j�ݷ�h��1}:?�kk_I��g�1�opP��3�(Y�c�6=켺��`6�5�ϴ��L˷��N�k�~��|V~�X>���ozξ�ۻe�R֙���L��L��M�07=w:�5]��񙜶��[sN�|�k��G���N���/��_Hj�z' ��vX�іh�#5p��zi�v��ȗϹ��	^:YR�Z,M�e��=�n5ѳ��
q��F"������S�z� ���l��UڪCA��w��S�d�4ɤSYM��O�����i�R�g�t���.ީ�<�-��wo|���xϐ�X�$z�Hۛ��ÇxO��$O��y��{��=Cy,������,��͑�L�اͻ�;�>�M;>B�%�½��9�oU�W��i��L&�!e]�N\�wp�2���:2�h���	iS0X�N���V����X�|����L=��L�֊����h�d�0?pg2����,��6���l�Ld�
�nVί*�U�6ߐ�%2̐w�~�����_�1 �M�E&�@�qVƐ�淚��f
�g8+����
���y�=%�Km�v�T�1��nUެ�:3^�j��x�4`�{Θ�zJ��sJ�ە�Y>/9[[3s�j�E�2�C�{z�>k�I�+m-�ݣ�Bv��������A�>�k㺼��J�.�ix#�7�f���� �y֫O�#.��B�$�7���pLF�&��Wo� �K'-����P�}��MSl�^��μ�z���+|��g�<�ەe~�b��}�f��)T��{h(ؓy�^�w�u�7�/�2#7`�g�.꼠���-K��O;�y�A���S4{���_�{���Y���w�����"bv..�t�D?zo���[�=���P�D�vd(�}�q��c׬3�޷��i�}�䎜��/��<��1�9}�;l�xq��a��k'=`��%P����m���ZE%�{���=��_y_��uJ��x�~t,��`�7=��Z��K�4`��c�|1qma��ʹCt����8�q���Љ"�wB+'$Z��˂��ܽ�i�x��<�ͣ|=ν��;�gV�x_��{9OF֛JJ�}�$�ݸ"�)������X�M�։�����cԮ�q������ Ώ�?P�4���0���ہa�:�ն�a��w7��3�m�н��n��ݘ���.�d��3Yz�4��e�Ǉ��
��ӕ��x��?s�M�#o��������/����y�Ƿ��7�7�}_6p)F��+߈GGP�{����:j�Z�[�����H�O$�ԑΊQ�£t�A�QjMEK�兔)x1�)U�1��;B�9-�c�7%I�*-���rhkI>�I���_�q�O��;���F�ϱ�{yB˙��B�
�X�+��*0�H���\�$��E�{�{m�]|~>���:뮺�8㮺�����Ͽ���W�X�id�wX�	EA��u4gƜ}||}u��������\q�w��ߚ߂��62j�ۚ��k�d�-�r/��i(D4i��7o��~��z����������8㮺��$I �-#5&�.�5F���F$5�ݹj���F7�ӎ:���_]}}c�����q���|ߖ��4QERm��h��4m?:���,PDh��k��b�=�ܳ�r�!�;���&�S"�Po�j�ͷ�,b��+�b��"*�Q��)76�ҷ���ۛ��\�{�x/k�5���b�����zh-W�������h���-���{U�;��w��$|ªJ��
i��i��JP��N��;�x�s�z�ׯ*�+XQ�#�y3;��I �]��2��/�S�C���f� A����X�8b��zm^J٬�p�ĸ� �',=3^l��<��O`��oߔ�>]��\<���h��%�9�/ָ�҉�{ !s�^���MOY��k��	��)�im�����Co�/j�D��n4k ��$:0��\F�����\mt��b�vZf���欢��y���7Ʌ�ɐ���;v�� ���8����Go)U�9�d:aK�ɫ{f	��KgaDI��q;�.c;�w�}��r��b���E��LCO�a��n{�o�w�|g�1�7m��y;�i@����n�+���"\ݢ�@�<R�EM8좮�1�
f X�jwt��h��l���໻��~n	@.����r&P,@s%���Y�Õl�T)[Z��&5(0�/I��sT�w�ݏ=��=V;psHpvӠ��y$��+��\�=�^;�ަ�UM˂�$��<�j�'eN���ᵳ��ٳ;����:��ܳ&~��HH��4}�AqN�����]��߯� �M4�M4�X���-4��_h#'ʌ�'{vJh�!����z'�d�u<�z��"�0d�>��O�~3̤͇A`N��l����/S��ī��=i{=���֝ې��#���*M�����O9���A�ZɔÚ7�Ð���8~s�y�5<.���1��=9�q��#1�2(�R`��k� L����i���"o����{C�[ ��؀,Y
�,@�N��s�z��UNsO&%>B	��p�� G<�w߹~1�7�.&�!ظ����S��1�3��-L ��.���Ѹjzz������A;�ݓd�fS�52pf�d|F�������q�C�2qg���w
�����O����	Xo�!���a^Lщ�,2�QL��.^Ӗ̬�5�����Ϛ7��jb�c��%�՜�W8���m���c�"HA��S������3)���0�Ow��;Gcr�]�J��cٮ�sܞ��Ox֟g��w���Ի��{�����(ͳ,���b! cXM\i)��i��iW�I[��ޔn��qy�G�/
+@��c#L�[xήwV=�h2U�Z��j:u��i���n�;��F<s��h����\����b	e8sʃ)e�]1��L��������vj4T5����l��-�� �I]6�ҳ5zc�m�=�{��㶫*�l���#���$s��N�)�T�y�����j����C+�N�U��^��y�Cs7I�;�ӒG�� ��Ö�+	i����ۧ����%�[E���nVIJ}3����~��� �wf�t�]��C�t�|�]. �$��'{���033?  ���roS*�b��A��.E׎ش�P�~k 
���(�,#|�
�����O��Y�����d&ۆ���܍~W'36�,=ɜ�i.�L�$�bP�+�oi��U��V�ūݫ��z���G�v�֎��������^��V{��ͪ���1�JX�pKAĸՇ��
��$�-.�\��q��Vo:&7$��ͪ\sb�A�����  8��U&k���QT���U8c��θqW��l��xk��3uY�>��ww͗�����Cm��M���ao���rN����a�hK�AWj�`@ؤ��\��]��"^�2qCqӐZ`�^�eTᩩy�t+8w>uo<����J�?#�;�����;omva������"�P,�����:�K��Q��*#��s̅noi8%��݇���3�=}�3+kw*�����
��>��ʍw�Y�~o�Y����SM%4�SL� �В1����/=&��c6W��uR�,�( �l��pf�YX�j7w<ڀsڸ<�y��	�����y:�c�8g�H�;�`����w6}]�Ww�������n ��$4�g躋�</ң �h ���4�eb�s��՜�,k_ �)�Lr��e������D~]���|�&0�T�n�Twݼ��� �Z���,�FG(X2P:��7rg:X&3)��(<�XK/��.3pkB�\��P4����la���X�5`�^*Z[���N�������2�Y��� ����*���WY}���W|�Eanß��}, m.ŇR,��h��P8��A�Emv��<e� ڜ��a�xw��;�)곚�0,k�9
�,��5���z5N3 �E��pl�����1pX�6L�j��g���}dU�i�>�H5:���G�DRt��)�Iq�;���sU�6D�kG�.�B7��/5s\��'�Æ>ow>Q��������EKm��7����b�Rk^[k��G�ή/�/o�hK�X܀r�s2����Ip�I��\Kɝ�W>��1a��`�2�NW9[��sګ��XA���y��������`�K!�+X���H=��>�Z��}���J����a,@8��]����OU�(�T!�b�^@�h�!T��ʕ������I������M���˪ЪL�E���Y�8 �s�s�AC���K	�.YD8�Ac��S��4�v�NR���\�gU �2o���XPϵdH{��,;t֙ڶ'e��)���55�DB��I{�i�d An��Uv]ﶽ�j���8;�
gL�������v�z��d�̀�PMej�5��!�z�������슸� � 6� � ��A)9bB!�D
��)��OU�4��LrS�!����U8zd*�A4��>ȥ6 �B�,"pG�3�c)�=]��ܝQ�(pk�w��v�C*R�2����T��y8����=���F�ǶsD�nyj��/{�^8����}�哊<�F�h�b�Ϟ6�U�H���Ao����m�7�m�$cm�)q"��|�����N�Q���L.9�A���`��$_#���������0<3~���׹�U�5�;p�-�D�a`JoM��i �h�D��A'5����ڹ�\�Y� ,f�L�:S5���%>N|�����Rr��lg�N&�>l^���;-� =$9�\#�޵ـ0�LGyÂ�J2��a2���L(�n����1�mg�a ��.̈́;�e�{۳�c�s��٩ò
�ia	4��o[y+y����A��{���f���3�� ߈�=c���)�+�݊��9��ּ���Q`Fہ3�L��j�m\sE��޾����XVBc�NX���;��*8\Uf��e�d��<��ݗ���k�0�@]�3U&Ege�T��0�DY㹁<��C�fHA�z�����^������;-2�y��������x���,�x��0�w��v�Py-#�
�]�v���W9;ϗ����r���*"G��ءm�ڭ��h���b��Q�E�!�L�v���^F��<w`׆�A��6I�n����豨�΅�k5��T��MX����ѻN�
,]�X8�WCF��<-FSr8��D�4),��Û�CfT�H:BkT5K���WN�����`�ɻ8�]ߧ����uؖ�ݬ5��Y��Z�����(Bi98]`�İmm���G	��! �m��]�W����<�F�)�^%JQ14n*��3E�3�=�>��e�rˬ���`�KJ#�]0k�gk����$�M_��@_+c� ��B�	���`�ͫ�޹w���ْ�=�ӗ�~�����I��%���L�l�,\�����)ذܜ��6�� MR���9����[�g5�L	� ��`�Yf��������#a�;[!��v�(b�P@B�Æ&�B|O��{[����^��Pw��6�}3�<*zNmRa�A�!���NCI��>V�Lm0��P��v 
(j�����Ɏ��'����(e�,FŁ
/�ǀo|�Ɍ�W�&O����>r��'.�{[�e�����c5)Z�)M�*�X2�[�f��p�L�p�QE��q�qU�%	xo��~tQB��	�'.����j�&KWh����Օ&^V]�;:JN���C�mߤ��0�
cR�����a�ݕ���m�9�(5O
OV6�^0h��z��bc2����e&1�a�������ݹw	�~�7�Q_���HKW�S�A���D����lC�,�+��f>�O�ϼ��H� "j���0~̟��# ��xڷ�BA#m��q��ڀ[m�� R@$[l��kIX�j�Vו��L8P!���l�������WZ�|���N�"1^dێ����`��FZ�,	ݔ����� ��o��R�k��5˴և����[�ŖLوxL$�dʩ0�+���.⫹׽b�0�;�ٶ���$�{ډ���{n���y�Vݠš�%ń`�y��׊���R�Cd��'e�����S۴��!����0"S !��:�o}�|�+�/�� �m��K��D��o��
�Z�>���� ��6�vX1F\��S$�f�1�ijXGb�:K'��^JrY���o!L`�@9j�X��t�ѓ������9�!W_��������I	��Aa2��|��X"'"�U�����ి8v"�m����=�S�snWAv���c���gt���3�6��Ä6YMR\'C���]�o{i���==��ۮ���=᎑�͎[1�٩���<߰Uv����|�O��G�w�m;��X	y|�����uh�mC� '� H�G���đP#m��@#m��I�m��I�PMpkʪ��}������|�.�+[-�@�L�2ᤶ1�^,5�3�_�#pv5ȱa^�.���1��y͓�k����zs�a�,	�&D��4�:�?�i��S	�GY��m$�D<�p T�Twc�S3!��g���s�6���r��[I��`��)�i�=1n�o�yi�k�B�쾮"���E� �!�������m�C٥8�HMvC[�<!�����{��@p��� �,9��`j�ק�ס�Y[ ��q���6��
�X����� ���v4B�AQH4��DM{0B�������؀q�˥��]\�ק sa_Ƀ�,Sn;5��uި}�^�/%ɢ�){���8�g!ܡ����Mc����H�*�AIUz�&��j�^h)�mp-� ���e8�A�Ю�D*�����m��a�`j�8�U�gG��pdz�2�3�ɔY�nM����G�ߛ ���٩	�PҺ����8@�O*O��0������^�lM�C�v]�9�/��� ������m�F��F�lP�
1�۴X�� $��H�,� X?2���L��mv����A�� ̠&��Q	�!ПPf���p:j��>ޛ�^�sÛ90&�"��q%�0A����aU@6fr��"J��v���cN ^�z��a���ˮC\K�0;>�c�l����2�%c
!�37�5&���~ &5�i���u�!��Ő>��4�NCJC�&�ͬؕ�Vm�j0�&�q9;=������) ��vӎv�Ϟ�n��&D��,@�'4�d��`��',	�@G��uwW�ch�`���u�s�K����A��.$t��!p(��m-�N��v��;l3im�vX^ �d�{�{;q/}f�G���M�@�'����ݖҏ�|
ȑ��^�O{Ip��I�{���nK�0$x�/ۓ��͞�^W6Rn ��Wi V���݈L�����^ 0��{w�dO���_�C���p�����^���N�OQ���d�vu#�ӂ�60�&��q,w��ֈ���ŗ&k�L^�@��Sog����,���sh��x��Y9���r`���u�	e˴����.
��K޳��Cw}���#<b������v�G��y�C5yMY7���v{��Q�w8=+�%��n�_Ո6�q�,^�Z��A!?4�.��xU��~�_ӟO��-�B2�OXlU�N�<sQ�iZ�sϷ���;j�{׉���w�=�#5�����'���H����kgy����F�L{u�۾�㛯��*e�jcM�g 3�s��rm{�b}��Q���,����7�^�oO/����Z���ں�����)C}=�Y^����Fk�h{<���n����|�w:z�yM��Z���<��WDȾ��y����X���څ�\>�G҇�<�yFn���Hw��+w\�0+s�e8|f���Y��� s��]{>)M�X�ge�%�n�[������{�	�p���b��Ov�1��v��y���/S/������6�x��Y�Q��ۜt�{��	�Q�|��L�5�/+�W�9��d~��Dg"��}a�R9P6 d�<�lM81d��K,rfEplcX�[�$r�FO�7��y�e��<2��F�9J�E?py��G���u/W�%�X��N�'jr9�	��^FV�f�0�6�P��7����l L�X�BT ��a mR9��5��xƚ|x�������}}}}}z�8��o���M���S6+F���i.F4Ӯ���]|u�:믯�^<x����C�|��H!"$�	"vT�4ӎ���믎��]u�ׯ<x����?!"Hr5		 �-7���X�4���4Ӯ:��]|u�:뮾�x������S؛$$FE$�<����yޕ�Y1b��nV�6mx�TW�v��sX֋�}�j��{[���sX�j�6��F�_�nh��u�Wb@�Z�`6	;r'�b�b�3j,�o�E�+y�"�m�J�d���V]�a'{G';�Է4��
�x��~�N���9���_x�Qw�JY��c�M��W/N��x�c��8���3�KXl)q��Ŗ^jk6����6aˍ��OY�^u��A2����M�UWl�Km3��0�g���kn�\t�@��	;M2�WXj����av̴�`0ܢ��͎�qX(�g�1Ξq��nO��f�/M6���i�뙻fBƨ���Gm�$���jp+YflEXl��
a6�^�ص����7Ma�4R�f�ڏ'`�b��{3�tr;u��wM��'R<�^, �%6�&eũ�
V�ٻK��ɫ���N���*Mɝ��N}g	�r{�<l(A�S�����s�C��q�H2���X�#��sv����[��Y�i�9��������P��bfT�]�����Q6��� :b)i�7y�$�'�Ta�5�n7O$�]�n��E��K���f�=�b����&�$�7<�`��@Qǩ�unM�`ڣۇ��cL�k`{A�z.Xf���ܯ<I���Z�_nA�l!�b��a�Mcv��瓎�6�\Q�:����Shdi�6\km��Si`GB�jm(AM`i������Q�<�e���cuk!3HG7/��il#��t��hrȭ�䮨��Cs�r>7WL� F6hkcG"��4�Ì����I���z9fv�۝]7��hE����.lX�g�v3�4UDԭ�
�C�t�:m%Y�mA�5��K�%�����,3<�qh��[lؤ7 u��@�JrJ�����k��{Q�v�P�#[��/>��=[�c�L�<��=��&��U5Uq%��έ�y89C\���]�os�U��)�[������#��4������K����;�<�գ��͡����m�C���{��;q���#:]`f�.ؖ�RSCKaE�(��U~���P�㭠���j�m��"�M�"D$U	f%� ���nR�	h�~^Uv�O}��}��u~|֗RQ�K�]͝�Y�8*3��v�����\�s>�R�!p�w=����"T�����yl�'5��E�i�H2���n�Ԛ+N6&�si�;-�����a,�;��]l������ݱxUrQ��h�%k4�ޖ[gvv���8����&�i�U�i�m��;7���҄:��d{|l7��"�<J�^�|�ABd��>�a`{Ħ�`� k�3�U&�����Xw+j�ƻ+��oo�4����yy//z��7��B��eD@o_N��nWi1^�t�s!�;it"�6j`��-����1�T�ذ�L�$�`�a�B�T����ga�%�@bQ=��W/�j�Żg:B	��9�qa�������Ɠˣ�#d��p� `D�����Z��:n|�6 �^I��n�׷�s޼��
a��
 [C u݃�%��pRr���xr����o���Hr�v.u�Us<��y=��N[pl�7I�������5���<a�z��n�9Gn���Q#��dI�G�����K&�������Z���� �y�,�ᡎݠ�����<�^��0��o�|'P�s0��V���Y���6�m�͝�����s���&������ې�1�XM�Y��e���z򵲥�aܸ�S��ͧ��ȹwa�"He)�������.����9��6rrx���_��ƦE�IMǨ���r�.�����3�)��=VQ��o�
��_I2Ǧ����㛌����C0$D�D#o�`)q���%��Ucm�"� cm��BED��@[�l? }���=�j��/j�D��o����2�����H"������QV��0�=�@�ǝ��y�q�<������	������W���r�n u� �,�(�RX���hy�c���1 �a�ˇչQ���|�\�\��D�\�iLde�{�����8B	�DUH?p���@g�[�{�ޡa�����+7+��zjj��t��ə��Â�K�=.�ߣ�'<�X~hyY�Ty���mRճe��:*\���s�j%21��`X�((�A�H4Bٜڽ������.�cY=b:�=a�1�W(.u�ND�o�G�+��[�g�Hq,��_Go-�+ ojXx�ErU�Q���|�\�hebH��Hx>���n�f�r	~���ȓZ�%��*Ȃ��  3�=�ޅ��hW���������v��%��2�w��I}�6Xw�Wlzni��j0_���S���
(m��F�m��#m�n
�Ȋ4�~|=�=����ɩ��bT�o�H$2�p������T�r3������v��HC=��ݝ��N+��3m �?%\��~K�ʝ�#�))���[i��ǎS��u, ���]n�L{z���{��
\�)�C	b&2L��&Hz��z�����'>�n����.���f�.��j�v�͏lT�B絛��K�"^�]���i?�ce�1�N �2��<;*wz����QaUo�gg�N=6kep#�3�#���0�aT��L1�
2Γ&c$�:�-"�3�,��{�ݻV�ӊ�@���,z�v,2�FCy���f�Z�3��L�Z10�e�R���T�''��T&,z<�������@��gf�1v+�b1�k�lE���U(�)2��f�J� � �Ań5��!��������o�z�XW+���K�G���%U�郆;�����.l����=��^�Ywڡ���u�֩ݰ:��4Mo's�*W������b#�~����m����h�m��#p$Y	��a�~�ݣy�7ò�$ǽĎgi�u'Uf���f�h�]W9��q1ӊ�\9{�d� x�Ʃ ��!-9Ї�
�p���sԉ	��&�A>𕙼�.��iڤ�)a8�0�,1�n�hD�gg��:�� F�$�� ���1UN������1{'���wO}���k�X.��� ��j� �̪�<��W���L?N0b[д݉�����3��$y�-k�f��D
��u�f3Qc�<��H&�8,&��B2E���Ā�%�(f����y�{洱�t�n��b8�o =i�@���ɬ��y#m
`����A�(��.Ku_<^w?F/d��@y�8@� ";���3�c� it��� @�(��@ ��42Ƶ��ʆ�Jx��ٰ�'� ��3h_w>g��\�GR��-z���2�'�yt�~���{������h(r������j��\s4�²�����D0D����A��?�~F�x�����^�� G��jm�ط���؍�B6�wREdE$X0bC32��������B$L����{��:xN�R�+�2M�f���+�ݹn�:�]��j��5�_[1=��Gm���J&.��9C8�]���,��^��3�YM�kػ��lbon���y^iU�tݒЫt�n�P֭�cO7�3uh�`�7a�R�13��1�r=H8�c�^G�	U�S6`Mr�]R��6�}�����5�~�0�29��39����X�/o���f}V������cc�^��W	�9���a���/2�aYw�K��:���ײ�>�L�w!,#|��s�j}��x�n��nG=z)D���MFK3����k *����v����{����@m����=�%���1{'�'�;@�!�1�@"}���߇�0Y�A��}
�O){�� w����O �x�Vv�g��Z$�rah+�hdǙN&�(���t���{��4��΃���oLU��4�_���<��;)p�&帤��vܾ��̟XE���b��N�����3�`�Q�9���r�d۾=gv�c�'P#g��6X�0�p�L�8i���?vN~����?Ch�V�L�sW��nCCۋ���n-�ْ3 є@>��#��wXS&V�ެ��ow>d_��I�������������,'`��M�&N���|�$;����_��!��{��P�H����wFw�(�b#�	�Z(M��ۍ���i���ӿW���8��`�F���z��{�65>�N1�+�e����Y�s�P�/7<�:>r�*#l��قY�����5�{ߢz�#�a��� ` 7�u`��������d$qш}R��7Q��p��hJe���㊦� �+.��w3��f0���K��m��� ���n"F�m.2 �� �"���(H�����o�����Μ��ϊ��\5NF6���]�����Fow�qC }�g%݃�!�ҁ�~����|�r�������?FG�����zYfy�|ƪ�]�v�F���wEGd���v�� j��2���V��ތ��Up�� �Ʌ��z�����~��<�q,�l�h1��{�v���2�%����C�����[7ϊ�g�h3�d5�HSH�]&6p��蓠�($�:%��	�G�뮺����M�l���X�������l�O�G�����9�㱚�`�+��v�FG�ܴ��:*oo��~ z�G�:�y�8R{t�~�c��@U&�^N�0y~�_���\Q��&�s��iÿ
���笋��
<��7�bޡ �)�/��3�u���p#-������������Ǖ<���gλ_g�z�G�u4���rk*�.���v�U\�g��ȿ���{�\�4V���׼����T���6�pF6�j\#m�%�$@�@��ڣq-��ѵ�jŭ*�WA�	�������^h��A˱��� 5I�`NM �Eg	���9�CH/���k� �/5� L�1�Tc�Vv�FG�� �Hq�-��l�� ż�,h��7��y�p�'�V13���w*��kk�m4� A}N��x�����~��GX�3i����0@��^^L�𶞮|�'<�����,��/��(����b�l�BL��Y�n	XZm2�Y�|�*��KI;�~�a���g� �>�gN
�|W�6�s��n|���Q��?b����ew�^�jwpDՈ�>�ȁ�� ��� �D"+���9��7�=�����D>r��3U;�-��jp( �rS�vA	L��r���K�w$��*r�މ�Hy��z<�W�wq�"�7�Z���s�I@�$K� �a/���v_ݳ�ȳ�7]��|�zn��l�>+κ����C4`����kY�P|"}{�wR�~I��}�<6x������o�(�� �����N����tx{�(�����F�m�B����� ��P�2"	"	 %�zN}��ʞ�[eT��̨� �sr*k x&VD?������P��`5c��3v+5oFz+��<�d�!��wi#������l�&�s�4i�Sp4��MiC:B��tZ��an��b�;4�x�'e;C �2�'2��EfGwr����
<%�T�s� n�D3�ڪ>A�2[���=�-`6���C�3=}T�7ϊ�s���57��Vo�w�&P{�E쭫ֶT��_��{v�4ν�|��������A��/,or���Th�g���@�C�U;��y���X��=J�7�7�Si�A��^�*߷��\\Ms�ƥŻ%��%:3�@7Z�������H
e��W�V��;&�����n�/f��ֻg]+ne���9��1�d�u�3�m�W���'���^���3��Q�\뙻\�M^�r�����s���R����f������%�wY���'�p�?6*G����21��m��m��DK��"�p�ϲ`~ў�������!Qh2R/)N��n�:�'/�r�5�5���i��׶MS���̛L]#��\����>�y����۳Xsx�:�ń�J�rE��4	�r�iB����B�d�c�����4�X*ib+���A����Zom�v
cPtg����;�g#ź4@=[^yn�i[Z�g�ϳ�,�{Q���y.��F)
.�P�v�O���K'AI��@lb+K8�)9N���8�j�;�y15�j��͍����R��O�,��y�f\]Q��;ϯy������ʶh��ư4�:r+�c)��@8 ������~<������!$�;�*�����dTMhv���B!��L�xW�N\O��3���I�3	fةwXE����R��v�oE�\zģ�����}���߭e��n�M��Px���SYNF1�Mg����w�n�.]��!?3��p�Bg{��GD[�6�Y�;y�k��Ӹ�y.�Y7�JNA3)�)����Ynx�e��vS��%W�;����L�p	wA��["!*��|&�d���#�|�<-�($GX��#θ��A�1 ���.�f[�������a����%��@"�ݨ��o�:�mu�ͺ\�r����V&����Z�)�1�$/[U+^R�@�;��B����g��,H|�F.j���yݻ�

�ݚ�lK�G�+�tZq7=`����'�����a�!!��s�ܒ~��!"�$i�l"�m��.��n# Ȥm���"��?a��3��|��������-���;Yb�c�O����=YS8�52L��NZrH	���fTK���z�b��e�R�xX�4o3��-�isb5��0���Bjd$*p�D��N8�uRB#<���wb%2�V�G�yM�Y����w��+��4:�Cu'"Jb	�A�y�R��]� C�{�C@���쓛8��kd����Ebh	wN�S^�[�Y�����/�s]d[5&M2�ySI��#�s�v��7��r���/���X�A� �ܙ2��^w�Z�;�����'��7ꓸ')���A��j��f�°����b�ƭ��đt�Ņ&]��=z�\u�mp-֝�#��!�5I�{S�� �T��Qq�Wˠ�<���T��<��	� �y�ې�g{��_�S�;�`[���|1�=�p��_�m��{����4�/�nw)��-g&�v?vs՘��j������H%=E�N��\�؂�5z���{5�Vޫ����=�����YԳ.�Lg��߷���ye�)�H=@:����;���-T�7����=���n�7ƣ�g�=u�\�R��'���Ӕ�}�,�lG�yTPw{}PS���Z���������S�V9g^���^{.��!�*7��|����%1������߻��S��������{z��u쵹����e0�4�tEyz���CLw���vy��<w��k�{O\�w�q�=��.�����/l��aؖ�p^�n��7Z²�>)�ٳ�|�����1��nU�=OB�Z��/^�Y+_��[b��07�O��ߏw��Qhw���,�E�uX��:n���Vy��wz�������;6k���&�,�^׼�>W���ª� c��b\�,�xY���8�߅;���3x�&o���r{&U�tز<3Z�
ͺ"{No��G�r(��S���]�xn�Ӝ�~}����CxKE6��$��q>�{n���u�ݻ;l�
;:���c��==p�[���|���/�w�9�z���w�G�������ءo�����Y�� ��d�~*�X4�r-�����9_=�f��="���^��y���;;7}�ȃ��0�J�ӌ�X��i��|�*Ɨ��	cW�>~
�X�g��*�`R���Hm mbr��TR�5��p�#m�������뮺Ӯ����Ǐ__]O׵sk-��yڍ}*�A�4�n����]u֝u׏�^<����|ߺ߰��s㗎�i3��&Ũ|���dI�co[u���]z뮴뮼}z������M� �+B�/ʤ=�QcM�뮾:��]u�]u��׏>���4�Do%�k�܍�]6+⾚�����$�V �ҵʊ#W�ub׾�Z5zom\�y���^yŠؤ65����̮$V����	>$j H��[Z�zt�����w�~5������l."H���D�Y��o6��ű�j"�F�0%��	g��'=��u�gm�����&Dϙ�%1b�ǡ{6����8���])`E>I,�s����Q�N�<1� >�x#�A�a��h�q��D A�p����6qS8tɣ�=���R��f�֛��� �Aعʤ�jM���7��^E@�1a |b���C��R�ң�,s�C�ngm`9�=N� ����I��{��4	�5N�uv�/��.�͵������|��1 �t�"�݈���,p�H�����8<��E%��>���c׽<$�X� �*o����#�B��u��
L�T8%�	hd������ئS���&�&��8��{/�=u���-֝2Y��d���O��E��TJ5'ng��4�����@�悸_0��8���)@�#�����$/X�����X��r�)���>���S��=��җF�W9�(��w��W>y�7bb2� � ����dc����	#m�� #m�m�؉pT�$D���I�HI��B��;ER�k/J�� ���*n���'ҝ���7�����'��b��b)�a�@�T�Ҽڗ����c�S��$�ܝ���S�e�ݺ\���#��lQ(��q�:B ޿��G��&�M^�^��Y��s�	X�/zL��:֐q2cx��fS�$�c2�X��O1��A=�!HM���^�A\3[k��!�Ȇ����T����i��Vc��ۘ��A�N����T��U/W�N��BA��c�����^���"V1��v� �!U�2*�^#"J&���N&w��4�B�G��zv��g�֗A�Mc�vҡ&z��NŶӑ%A�A�3.4�N��?�����=�y���{���+�k�6�:b�Qͥٽ%���H��vȎ�tj'ѽd��A���S
��PxL��/,����&�=���W�q矰�O���� (�5�r����^�I�$�[|������q�m�[m�`$� {%�ϴ<��/)���D�S8R�`͒W�MkM�e�ҹ�dЍd��{�B�tTjZ,�6he&���hdm��}nk��Y.��-�`ո�=�uG[��s[�x6�蹇�]��O ���	n �(�6��ukH�m/�ӛ`�]x��n{�=�����n��U�mD��I� ��pO��d"�+�G��$��}���a��}��[��2j9�Iff4-��M���5�BD"^�=)|)�J� ��Ϩ&�R]��|3{�����<�D�:��c� �Z��fP�'��LP"�.>�X���Z�F��H����{ޮ}r�OZr8|��
a\L'4����'e;ڂ�j<�P3�I������B+��4�"ü��g6�3�E[n��������]=����a�ix�2��k���*���7���Wt�{�i�5(;~'��ݞ�^�:0E���p��]!YD�\;3���5y�ǧ1�16Bfk��w�<"��7֭�aj��T3�_���@��h����p�����A�k�px�vv�$ag�ƾ��e_���g�%is#�Y�1QL�|�w���9��ɒN�uB�=���o2��k1ɝ�L� ��ND��uފ��A4u���L�3�<�ڨ������:W�~���%Ovx'��������'ȩCʧԼ��� IS2tҐ$��; �QT���].	m�7�����3y��W��KF1�	`H�D����q��v�?Wt�{��E�@���1��CRʜϸV!����wl'<  A.:)�	L��8��ENA"fcn��D���A �� �d�p&ekƏ�0��:������gPa^�T��w�8|�C@"]2knރ���|� �;�&�x��X�D˻85��]R� �-b(�T�,�fōc�fES�Z�]�q�I� �ShA�'SQ�2���ĝ������t���44f�1j7Pam�v)���ї.ł]�$�l608&HV�2d�R�ic�:�7�(Ȟ{r���Q�!F�L��L�.�O���P30�"��'�P�R�:Xxj;oX��/z5p�i���1��p�Uz$��x�؊L��pA;��_$p`v���&��&5՟���»�����Ec�t8�y�psc��iCL˜M���=��v�bA��ϙ��IG.�xO�1���m���m�m��[�2�ǽ��i�}����+��lG�p�x��eÑ2��}�:UA�7�/S;Rn���_Q�<ݶ�qYt���_�u�ײ�k,����P�Q�-0��0Ԃvz� �����z�����ne�g�^\����C��#-&/�e �Z��������}�_�ϟ6����)���b���6&�Vh���D�j��.}B���u+A幐'8 �dRr%2��w�h��]�8�N8I��#��J�	���	�v���	�!�Qa�F���\'�G��2^Rn����8�^x=��n�8 �&@̩����G�DlPi�m/��pw��� �8yTC�G�T	m��Q-�=�:pS����A����ͫ�8!1��L��JibeA��PV�C��1�*��!���z�`ѷ�����i��1����c����*�pg	Y2��ʝ�˒�Cٕ()����S��<Ƚ�0]�=��v�ˎ����O����'=,H�h!�4���>a�?��m�ձ��--�ۃ#H��[��p�!�-��W��Q�r�C�@�*�&A{�����!6{;��������E����Na`��@L��ᯜ}2yG-p� ��$�Aˢ��������Y���`فGGl#��K ��{�|a{�}��yÑE A.�����������D��s8<Q�������)��2��k�f{�����N�fS� ��wF�=Y�~���kO&�CX�;�Im<�[�0X���k��	�.AM3�M3�"&�ygG�e�
))�xU�����t��/ A�!�R�i�pZP@��遦L�B��B����� w\q�5����5���"Jb�֖���׬ai���c �' �T��D fT��|7e5(�F�7���wG�g�F�s Xܦ�02�8"�&�q�r������b��{?�	�:��#��:O?z�9��x������dbb��Ѫ�i³o�kj����b*��Ă��3�����m���#m�\V�~����n�3�'���,���ڽ�_:_�Ie#�a5�M�a�=ͽ�<К뛌n��m�:�۝��G����;�^Y��k�\=YS�g<�^n�4`ʍю�fl+6�� ��c!CBmt�j��9gnx�����He[1���9�$G�wbv9è�,u��jh�\�d���KWm�l6m3�C�v̫M�^=�e��g�n~�Ehy��"D*�J��ϫ�j~����I%�Qh�p(�v�V`�8$&Qسi��m�a�u,�Β�����Y��c>�Zv�wbd��7<Uhڣ�x�%�zm�T�b����)�#$ o��'-)�vAL��PU�F�1(;^W`����u��X�m�^��
�]��׵ab<��W�� ����K�ĭ�z���Z���W�! R0ײAɯgG�g�H���@8PH9<�$
eLM+�%�O����_����qI�b�l^���8C<���}���pͅ#;ָ�z�1
�d������� �ǘ�@O�ieP���!v��ag�":+�>>=�t1�{/��竹C�w�\����pi�v��UL$K�Ȉ0I~���>�]X��vf�-�S[mM�瓶ں��^��뀛 ����TFX1v2��BZݜ^NU'n̝G{=˼���n["�z�}����G�0p��������Ť ��bq��Z�_ތ��̩S4��ɧ�}VY��f�U��8W׉q9n+�>ȳS3*ҹB�[�;����m��m��! I"�ϟHNy����v"�!ޝ/1�s���ӫ�m��w��� �kraj�S��}I� �&9T�4B���ѼV:�� ���G�{՛�9���2@�PI.�%L�zB�V�c���D��M���Y���L�z�s�{=���1�87+(�AȼV]�h�w��`�b*Ńp`�\8"e�oL-�#�p=�^��Tz(wa^�ckW A99SS��
��{�����~���au��:�Wf&�!�U;o<�
�]u��yޔ>Ϸ�yIO���v�$@ ̸L���"�{����4�&�JqB7�rBcLU���wj,��ڂ��1>����=8��Z_gbuy�{�ި��=��&<"�s����]��Xi���9���;���$
� 2�؉M���g��Ց�.��C�E��=�����j��x���"I9"��$k�-���3���o����J��y��@�>��7am��m�6�m[H�A ���N��
6<2�+��H��`Njr4�2�K Y�y�c%��N�욇A�-m�%x��p���������:��6	%O��Skk.�؉L��N ,5�UI؄�y�ơr��5A]��E�F�//Vh��8��n��P�U�6|�7��Һ�rX��b0�h�!�^�y�ۇ�m�k�5�b𱳎> N� ���������ك�Qzq�l�bO^�a���i���3���g/i�,j���0Ż1�y��m�)P�"�p��ۚ#WOx�l�v��6ÏRO��r���h����'�;E�tW�O��c���C�[�VӉ��A���}��{/���n�#Ã$2��A%�<��n�IA�b�1�KHsaep��7ҕp(�;8@�'`G�V}��?��OP_/�B�t8��4�J��Qm��/�t�r���|�����;7�{��VO�mL�s.���!�a���gr@v�ہm��F�m�H�����q�NyNA%4� �ʩ���ds�B�w��^{v06�8���ŋ͞��\�d"������2-؉lv������[��z۟k�պw6.w6� ��sNhz��jݰ�8`+&�8 �@)�g ̧�9ò��L|x��Վ����8-�<Y��p������F�LE�XK-�Ԙ�.�m2�z�Nk��U�H)�L��8���=]�����v�S8�9�;1Wn�@MT��C��$�ܟ�=��`2G@��n^R�s��}�=��7϶�*vý�l;CGp���d�r�{|����Ȓ���@X���ܭ�w������f��v������^;�v�w�oaL'C��C����g���L�
Чl�?�붗h������}�B_�d����ʡ�i���IE�$�Ž��3�)�(A��'��Xx�6�����=�1qҺ{ڧ�:�l�0M��ȥfs5c�ۚw��b{�����^0kƌKU�G{f���_�"���su�o���M�ny�	s:s>�me�@���{�pL;r�s�KuN]5e��9���:��M����t�v�k����p�c=��FnV�@��CFR�������d��^�x��툖��;�����{M;�`��f���]7;Z}����!~��qk~���(�D�(��N��һ_�n��s?	���Z�b�T�pۺ<��ŋՇ=�0��[;|G��;�pq}q<D�SK����9u{p!���E˳gb�r9͜]�X�.�������m�C޼F������m`����W���'k��SM���zTw�A���ɯ7_��x�w�8x�a7�G�ؐG�sY8)�y��J"w���z�鵢��=�1.,��{�X���KxA�fvi1mF�k`n&����-�H݂�*���f��X>:�b�F;��|���k�]��opʋ���fz���u�{���T7��\޳����������KR4x������I��ǀPo�,נ���J�������O��o�gtx��0��e�.QX�9t�X���D#�X���c���#�՜3��Ϙ���t����^�WOl�{����u��7�bu����o2���)6��׋\�Qm�Wߟ���ou����]u�]u���Ǐw��~�W�\�b�DQ�dd�T`z��u�]u�^:�:�>�x�����d��U7�h��-�;�s����6��]qׯ����]u�]x���Ǐ����=��h���!P!%RT*9�H�J��Tƞ:㮾:��]u��u��ׯ>�����MJ����TV��u�¾6��گJ�E{�+��y���^-m����Q鹤�+��s\�wWMr�ww}�sm��Ҽ[�7-!Q���o�k��nn\܊;��W�ҫ�5���9m���-֞�a�s�n�c _���2;�S��.���,�is�&Hh�,�����득לݥ�&�������G��^����B8�F%�WZ��1anmVnR�|㜭�tc�"��6K�� ���0Ke�;�:��Gn�/ �WtU��yx9�
^`%%�L�X��r-4G�eͫ��\��3c��=Z憟\`B;>s�jӇ��R^�ݤ�m�bSz�d��<v�;�ä8���]/p�ԣ�KM�[3(��ls�Fgέ�Eƺ����<D��ksfc*n<�cf�<��,i3��\�������ki��V�������E��h��S�wl�4�*d���Mt.4�&3�K4!ˣ��uea�@�T$x�� ���ɻ=71��M)6������vm��%�|n�x1��qƗZ��8�On��>�vE���7e�i[�f��X1���&�F]H�r��g;���a�+�����7��qV:�e;Z�7Н:�&
ل�մ���kRhЗko(��l����p��cy��Dm��-ր,ݼ�ǲV�l]��]����{q��n5��]8=!�/��wA�t�������p8���Z} ��l&6�m��8I�fh�dn�zwn76y;e^�8������	@���$�>{cG��b'���r�ޝ�Qd�,�	^3Am0\*b]]����_��䧺���o��q�]M��lY��\��8tʼ:w��y�ݫpUn6��)˥�pm�cgŔcug���mi0���dz�b�=
�p�x���T�ۧ�+�m%�6���=�� tx�R6l�0Kv�^��힩v�b��� �nێz�\�up��9��ޜ�)�1��Om��ɜi��Z�UPj�����<�X�ú9:n�}�������Z���:;tj������:�5#��/h�7�����7OS��;۫�p��:��uq�����;}���po���;.��q�Hn!9�/[۱uqkN�A��������M4�@4ݲ;�×�O���Æ^V:�;��\!Pi����4ScsM��]���u���#0�Ђ�tb���=�3%��g���q�Y�lI7n��H]��4;]<;�ӵ��u��E[n���1�m�ܖ�	WU���۰K���J3Tke,��#m�AY�N�������x���v��'�b�:���S(��9ס��v�>������w��b��w�;��7ѓ4A��{�p���n��ò�ɢiڗS��"�І�(��>�	�c��89�A�#<\
�H"eÌ�1b���<g6Rn"8<��x>���8MMS�$Y	"�̫TY9zk��z���I&��O{�+�c�8�9��}H[c��������������L����g�p���v&H���r���%1+��q�X�����\[1܂8Ze��)����8�Z��|�z�  ɴDӁ��$L��Uُ/�xC���^�/�mj�E�;F�!�ʂI�܂4B�ʪxy05RY��ָG��u��<=�g:X�!���8S!E؃T��ְW���>��?�*�������e���,pp��1���-�̮5x��pH҈;.3�������*�s�����I���\���Y�˳�!B�&eޡ���dԐ�DA�x��v��?�=Yw���D�`�K�F&s��ӝ���r�B�n�����3����':<P������__�m��j�m�n^�6S��ܵ��b��xC��!��Y������Ȼȑ�w�p��j�[|��&K�s2���@ϔQ���~���E;��i����s�s��(�X6��n�ve�,��)�8<��A�UU���ز�>�#13�!W�+�9�����N[�L��5�>�(���I�I̠��撝���0��ҹ�zkY#���lE�ޞ�|�\�������"e�q�P�U�T�;�磚3�wU�^K�q��MiS�Y��p���O���sn���̧X��8���]샢o�g7��+��1�co}��$��w-���S"eÂD�X@�Ә�-L;;Kؒ/���Az�d�?TC�m. �,�\�7�H0�]�*�_�� �s�D���kU;b(�5N�|�\MT���*Ǯ�cς���S��71$�m�U>O�i֚m�=:=>ȗ�L�Y�u��B/�\���v~ŀ�H	8���x�5$,nl,�Hw���ks&L��ggdɓ8p�!��&�5}Q6���}�
��;8 ���AșñHFe;����ֺ�]�:[ڡ�,}+3zu�bƉ����@�Rf�@���;`a�C�ɇ%�����(�<�P B1#�6�|6Lh�"|�{���q>n-�ql��#d�]���S���?އng���;�,4u�s)a�z@5h�g��Dg���uz�(&k�D����Fm ����%&P��Ǌ�<!�����d�5���w�j��3�j��(�����Y*x$�������4ƌ�g9��r}��>��o���r� X���!�� �;#{��}w�t؏�s��Ek�$QA����Q �T���6�ݼ\]�$w��J��/�jk_2!��\ŲӘb���r�+�Z|�n��{G���}(8 ������W��B��D<^���Yc=�L_da�Z�z��xe�̨���B0{(Ld�-��D0|�xi{�O+���{Mz!���1��9�&��E�Z�}i���m���,���	�?��(g�B	@��Re�%Jp��ظ��%�DT��Z�r�kP>�r�/ۛ�ǰl��y�$Sy��`q�Qd�N(@_�uI�����������!�K�����S��Fk���'�`�)��s��\,�W.P2�ؙ!GE;���~ȇ�ۉ�2��r�I�`�x�{_�N�G�����)���[e�����AQ$�-ڃ�^��<!�������#��"f��gc��Y�k�يF�@0�!>x �73Ө�����RH.}�1�7�o>���w��H�c���d��Wl��5.-��'��	�F��b=��CNC���ޜ|��xzޭL�)95J��░�d�W��$ۻk�@���cv��[�)�e�:�O�v���{������u�u�%���6Eۇbh������ ��O��w���].�{�����}ӵ�z����G�������麴@5�7-���v��ɓ&L�L���z����~\�ʢ�ѳ�9�����U��u!���X���^\����]�i�!==��kP��l��ٞ��-N�AZ�s[���gѽ��������7s�j��ѣ<c���z#�
��<ݺ$総x��fWvY5���tOgAXa,֬�;�wR�XK��H�
,#� �x
e���Y�w�[�hk;H��Cnc�M����{t�}���Ϸ���Mt0J8���N�/��d�W�V�?R����XC��G�Lj����n����g��g�1�$cmx:��p<��,!��y;�,���9�C��fH��{ L��l�v'
vK"��7�5�"�)pf`[-ܱl!2��:f�f{��m4���.�`�� �Љ� Ļ�D�AeĆyl���"?J�3��W4�֖@Q	��wG�I�$����P��Ĳ`���T-I�3I�&e?�sw���2��GY���}(A=7�4w�e��	��& ��✐P��*��g�BiBd��_�6u�RkR����
'g.X���q25I�2RUN+&��[����c��|�DL�/6�!ݎ3�Ǝ��:ۭڎZ�])�������/�b3s�NI ����w7_"V{�:��]s[@Sw��R@����je��$L�F�;A�A�yWǘ<2�<�<����(nv��t��� ��Q�����/�O!ZVU��5������]^�~���eRv�|0%��Km���2`�2`� ����A������6���L{E�^dz�n@P��=��������a��8�4��bbş
c�9�W""��/�!D \�I�r����
%�)q� �eA̭b(�3O�f�%$�M9�Hw^��r�w^�k�6Xc:�f�uy�l��X�M�A�J�8!2���EFew���,�P'ڜed��L{GV^c��<�h�A�v�C���u,�.�U)�CG

�� �m��y��f�=�GS�Wai��.VY,��t�Y[�.�E�#�5�\sX��R���ؼ��;����248^t`]�<����igE��g�gi�����H;�+!B��$�6�FI��4z���=�M��2�-�a��pN�A��9ټ��D�&LD�`��ߟ�9>�
�>�������6Z���m��ۇ|�-D�M�|Ǩܫn����rœؤ���;����pf��_~�����!T��9�?P~�s��9	�m����֚i����i���@9��>�������ş���A>d%�w']o����/-Ñ�vv2��.F�3T_zw)p,
e�T)�*�4�I"��0��2��2���H@�h���C��F/�v�c��gOy�,E�-k�� �8g3.��|�m���}����h��]�G�`۔74�Yi�։��E�� �4hw3]�LRr0�2�P�pH7i����z}�]w��ƊbV[�́���h/�*��\��&<�,���C�ƈ@�OuoX�=��S�o�&��ɩ�b����}���}�A ����O��j��x]�����NJr(��B&]1pd�1h����dZ�E��B%�I��>YӁ�o�����pA�-�!� 	�3�n�go2UN��x1��j�B�iMl�Jf�^����D���p�� ���:<��5��zS�	"Pw\*��r�?�^�������\����ӷ[-��yx�£�p�J����صTj���h�?���M4ݶ�M��!=�F��a�,�<���Jg���E4��'}��D���x���W�k�o�{�Ov�pAbZg����Zd�O�W�~��N�Jz��Et�T'��$%֪qs�j�����vx��4����<��<��#�I�A؀N�,]�02Bb.j���rΞ���A�qr���Fq b`�I�w�!JF��%2���ҡ�����;�M�Jr	�U����M������ ��b�P�)��*$��o�6+ř�f��݃�!UI�D@S��f�@Rl��9�n{Ƥv��b�R��~��OV.7i�L����A�wLD����ڽ����M�l���("e��^�Ds�O�_9nd A��|��;��,�D�"]�Ȗ ʀi�5I�0���n�Կ�gϵ�`ϐ� � �ձ������|������\�b��D S�3��\�;�S����4�ƍ�{6<1y����T����B�i{=�PKއg_��
`�\eŬG��b$�[�sM�E{���oB$|���Q��5��%4�[m��M���!C�p�����r��"���j��q�>Q���Q8��n8�Ms�Q[�K^!s-;�f��ڝίD���1�������m��6�i	�S�t]����U��H-�ݡ�-�)�|��y=�;�cm��AF�1�:a�u�4�b�]��J"NMG@�С��cv��'��� �x4�t��v������;{�9�����Gd��{'�)�@�I��+����v)�
ۣQ����	`�o%ǂ�ݪ������u�n�5�1��ؘ�������s��,,j���"��[֑$�=k����q�>���ŇerSb�l�A��bh|�% Ao2������L{͕c�!1�(
��엍~�����I6@]��
�����_fp�~K3t�����ж�!�܂j�W�ح���s�hee��p���	'�1��%��Mn�U&o8�7̝�H�N	�OX�jv�r]{36���鍝\��ZrA�u2-�-���Zr!�,xg�L}I����ʜ9�H^˳H�����I	�#�v�9�g��_6Wk!0m 3 e�`A>ew؁i��xU��g�<"Buj���;��.�D=�
uq�sr�˛C]��߁���}�e���m23)�L�<.����Q��{������׻��&�ر�	�88B ̻�"� p�pE�{#x�{=��x������UUݹ�k{���:�jBg���x�f�uy�s���J� �]�F;;<<�<���^���PM#�$�V�[�m��M4�w�?~v�eH�4����=m�G��ݴ���glL��[:���痊�N�5�v]j�	.1Fq0fĀc�|q԰	��g�9�8I: ��^%���_^���h�	�1As�g(U;��22(��<fz/�[1o�3h2.�a�2D�)�+�{(����p�H����$
yPp`�"��b&^Z(��%�93�����h ���{�_�3o��=/�K�h�ψ"L�p;:2�3�+W�O_��6lOo�	l�Wd	d�Z����&k��-�����z%w�׌�\�gK�8#m�vp��p�[�q{g�x�l�zb���ޔ��Qrf�9a��J� ̠&W����p��І6�q8�7��w^V��Q��{���G��c�vTA��w��T�j"Y�`s�;���k�	3*�--��̑J*�]>t�x^c��E(n��q�-q(���xW�l�\��K������9���Dzf�_t���&s�!��ݙG�_{���֖��#�^W
t���I��wt?G�@У��+��g�g)���}Zb�8,Y�ڣwO�s9#�XEK"L�n{_"��4��J.��t�c�^+�6���"M����������7"���h������(�I۝��WV��^mPF�/s��%����G��E������@�����g�s끱�Ogc�{�K��ad^��|�YZ���b=o-��.2���ܟ�Y�|���0���^M��5���8v��&rw���:�`�yjO��N}�w˼�wZ?V���L\=��%]�3�D�AX�x7��5����D)ҙ&���;�*���8��n���$���7I/:�$zx,��L���Ձ]��}���t�;��N�[�-�M�wݳ��]���|�a��%>*��q�e�z�Q.�����|�tЗuн�5Ֆvx�tj�ɔ�v{{ʞpM�OS��>��F� ���{k�ϼ������5Ó� ������p�>�j�N?e��->m,�Bo^��������N�X�{z�	y�)!�׭{L��z�HY�;NN����e�-����vԍ��yMճ��X��挸��Y+�cNY3�(�ݐ>��)�J)`�-:����|������r�] ����TBv$M���x������΅�P�Xc?t�G)�,��W�d�͐t}i���xQ�R�ī�/�5�Ǒd��͗	c'�˓ �S�d?q9m����o(X���a�ǚ%���/�[�/&�ם��oܥ���������^�-�Н'����F���,��x�kIP���,�.�a��3��1#��\�p�(^D�+J�ۅ�˾�+��,�NK&�"`���{�����>�
�uAH�E�4�����㯯u�[u׏>�x�����a!=�����"l�/9����8=}q���]x뮺ۮ�x�������U�2E�)�2�r%{Is�ȕ.$��q�׎�:뎺뭺�Ǐ^<}}}t�.H���d.\�)q�#��"H]\�*��m��^:��:뮺�<x�������g��oOM�/y�^|�tW6��a/)L(�ɵ%�,��Nv׋�wuy9��\�+�ki������1�dצ�Q�Ư���&J�y2�L�ʆ��;���拚���}��_;�"�l�܃N�hmb{ʑȕ
��MF�I-�֚i��-���pY������=����W]�:����jӱbE�P+��BK�;ѾY5�x��n��jA��*����Ў���O���-��lA�,�Rؐ.���y��-k��jd�\ͧM.�T�Q�c7^����3&)�z��8x�/!�������7���D�z���g|�T�:���UK�벹�UŅ�j:�WmsH�d��Vh��w������4��0�U!-�E�^�ٕ��s���8!o�Ц7ѝ��TAM���')�e8"J ��AȊ���)v̱�@:N�0m�ߏG�g�y��
���D��a�$eܕ�)mi.A����g��k*�X�bj�t��=�2WNM��O���6�ŌÇ�"����}D��eIa���rP0�g�r�B�3� �^�-�_��5�I:��Zs�mOs���/�P�P�tg���%I�۔O����=��߆�����ʱ���el��W����|g�>�y�z��=����G7e �j�?�4��m�ݶ�i���a�TA=iؓE3)���v�ų���ѣ薠��;u��(���W�U�� �d�{�+��Z�G�S�ע���kђW����b��s&uM��ӱ!�D������f�^#�'���	�Me�S.�AJ%D�,�엮�s��8�O��7Һ!��P={)�����A�ڤ<��T��#y��R�6�"^,;���S&��a�2�k�/�5p4P*Ӱ �d�ܓ+ٔ�+�����aLܥ�vóN�����;	�%$z��7�a�����"� �i�ER� ��MqYۂ�i9���'`�e8���쇯w�e�ph�aL�.�_�a��c��7�,�v�㜔L���=���CΞ�ܿ�I������N� ���8B3)�&V���ї��&=U������˲w�Ov8}6���]�$iy4��������.Q�s<zs�xo����k�~t�?��2dɓ&L�L�6�������w���Y�=qx5�x �a�����d��㛠� �����bx�s=C��]���m�t�7g��Tsn5[��m�^qӥh��n��@88�@��]�v�
q{ q�\��p��b��L4��и�0��Bp@� �c��RX��:K��=v��q̓k�Pc
��-�Sn���y���<3�W��z��5StA��So�Ou�}�_>R�Hܖ��*�Fa�t^�q��Ƈ����F�"�f��1�O�?�m�������]|���y�
��;;�a����������Y��I�7L����=	.)&�NA3)؎���s>-��X���1���~���naOv��Id6ЎB�O�V_o��p�q����� �cn��N�Q�3�3ޜ���f�Y���uq�Zr	á��T�5H�j�Aާv�GŸa��Qp���a���� eo���z�=_0\��e�M<��.:�"\�!4��"�ta��ݧ�Ū�u�1i�_^�glE���w�q[Єw��,�ˊf�;a����]L�?�+�jy�
1�)�;Xu��X�%����BC��&.�{�`s�\O�	卼��2�zK;;)b��}�Է��@�{�>�׾NA�0�7	�Fi9jH�,� �D��!��{����C��ߠK���x0/7#<������o4~��*�C����N�����3Z�`�#�T=�;P�x�a"��2dɓ&L�2e��*�a@��~�?b�>��0�}`��I#�� �����7;�N��NHN�2B�%9̢���#	$k�zm��|�w��ɞPr[�da�P�{e��n�=�k|�7�e:d�ۮ!�l�!#�r��qh��ݤ��pB��*�PD��?2i���Mt�oɜ���|@~qS"=��7nn��z�?��k�B�n/�p�I9��o���b��"		��xxt�1xϞ��ѲtI��v��d�
!�/	x�6�[;`*ӐA�,�K�8���FftW,�����X:[���r�d8�d�U�f��&n��ӗ�>���֠��V)�,2@A�!n�:�pz��5���;�S5-M2����
Aȫ�,Z̝c���V�K��)����R#�y-������/���n6�����g�@��;�Y�0�zl�/9�� �h����������b{�2@���9�v
�ndɓ&L�2dɓ�(%�5O�9�	�z�\�b+pDˇ�$#2��
[�sef����� �d�τ819�smg3k�t��{�7�|��d$L�S�1{�����'"g��H�!�K�r&b�F��#X�>��'�cT:�p-��AZ��@L���F��[����u � 9A�:*K���w$�O+tnMZ8Yn��vW�4����f8o�!>u�yH�0���W�|��k��z���V����A@�,,�\
�gl��Ƽ��� �	�V���#�9*�Ge��:�vͩ�ub���3;���2�q���0�ȿ8|d&a� SL��D˻)�On~�h�rPIn
{Q��p=t��lA��C���N,j��d(��̓5���H��C �5�h�D���Kفwo[�ǯ���s��ƽ5����S�{��/�ۙ/_�0&�\��1���>��f�,��&�m؞еp�wx�_�豑�����HH{����i�]0�_�4�M4�L�}��"i5�,tI�L��!((������%�#��n�����U�|:�fPr��9�<l�gF�=?u~������)�u�	�%Z�l&�+>�ܨ���B'�B��:6�t�I$�w���ȐFr)�S �s_�v����K�na��y�.z��@�g l� �be;P ��������,� �,Tㇺ��{y]��|ޕx��;��Uy�|�j1�h�%����Yv��- �yB��
V=�r��/�k�flTh��E��<E�,d�j�X��B���KRqDS��C���e2
���y���/�W�� <�{uG�?��ـm #�e,h��˧q �����.��:k���#��v�����[���4Yؼ�>���M)��ןFM-�\���p���x��ť�/j:����g�+�|y`8�e�� ���s�ӈ�" J��˝�e��sr�Zi��i��h{>&F�����	�x`�'�]G���Ì&v��D%�b,ر�X����� �y{�@�Dٔ�pM��\C�$�[�\����(���ff��x˦p�(�'n�<r��CqzT�Nۘ�]%�d�-����ݱN�8����i���Ō��BQ���x符��u�q�W%�; ι���nLI�c2<���Ǎ�So߿I*�ǯ�����z�o�ǹ�k�2B�Mo�ɼ�٣��������Ӭ>]	I�x닣��;,�eR��,q��M�LM��D��Ie���,	�Ӱ �@L�b2���i����/�.�<E�c����$�]�l��h����Nb|��,d�S��}��Q.����#�������fq�����ͅ�&�M	�1��9���09�I�� �jPr�$��D u���b�k���{�I>��}��#ޮoJh��]��ۉ�����ݯ�r(kO�S�F [��2�Wv�%�ӡ߆Oq&e ��Qu����Fw;��P�HB�B�ñ^�RF+�m8�2z��ۺ|�#;ip ����AK$T,b �3��3b|쇦>�v�	��-ΰ	^W��y[��OnɈ:7 ��[G�H!kh��fPr�Ȓ�3/�@�۬ԯ��d{�����f^�l|��7���L�Fe3�fi���$���ַ��v��>�&y��}�ig��iKI���v{�Sm~Z'��YFGBS�x��s�s^�^�EF�� �<�P�$��|~��M4�M?`S�E��5+�;`����2tN$8 I�p�A���	J�{�����AZ��|�	M�9(vBeÝgg)6���;��w̗�&_�V<�#�ŪӐq2�S)��g�$�/��B���F��!I��L �.j�x���X���\�5�Y!����<����yl&�R�H�NJd�̿L��!(��fC3�0k�zPۛg�ݝ	�d��Kp>��@[�2B,�w)�����.��t:�p��A���j��sHbc*�9�*��'�G��l5&@wi-�;�����?����v��a�ED  y�>�Lo� ����I@�F@������ј���F(<�O���X�����c��LAN<Є���X�3�^�z�[8;��N֠�4�T��	�{����|�|�O/\<xj�'�ý\�皶�r�*�������û��:�ph� z�;n�Q3}:n��cׯ�b�^���ܡn�"--̙2dɓ~����(B	n��'j��~:�X[|��q����-T�˸ۈ����6y�c��1�!��4�~�#-�msA�M���ױE�Ȁv���1�@O��3(9%Ñ%��/O��7�#������x�5��E�A6\Ky0j!؃$W^��Guv��<������߻Q��jm�<KG�'6�y!�uŬ�Zl�ֶ/
��)��{}K��8�&,�L������ᓭ��S��$�G�{�fB�n�-����������b"���II�!d�O@W�����ON���NAM���R�7S��۽���	.\�c,���q����,�{v��<���"��-No��zg&k�"'��C'��v#�p���Y=(#7��ª�J�X�|A��kL�-;k&�J37M��s��O-��b2j�X~s-�߯����+�(��L?�be��.^��t��t�̖��Br3U��f�v�{��ys�7�ا��p�2T#O�4�M4�M:�Y���B�� 2��2@D��$-2�I��5�~���K!�ޮ��Z��#M����n�qi&T�A3)����{t_���8����f���\�M&#]v-Yqp�vW�}���9c��) �k�傪H ��]~�{�:qz�X�I��|�,�?E��Y� F0#p��VŵK�iL����v+��)����5���0�tb���ݩ�/ݳ��O<Z��=޴;4D_�/�t�m�S�ɹYL�1�o�Yć��8��/�ϲ�����jAܾ#=�����. �n�' �L�fW���f�9z����X��g�zL�ç�kZZ
i {޾�{<ΨH!V!�ͅ��^NU'	����U#0�'��I��e�绯�^�s�r[���.P�A����8OlHF�sW���8��GuMx,�73�����]��!�q��L�Y��K˰�����]x�&�����)Z�����;�g��G��[�v�/*l`��o�^S����j�k��No?{5z�y�gr0��i�k0ў�%Ln���O5�{>�N�����xG�����"�-3���<�����q^S|g9�&S��y9��!��vn�m9�Q��T��������;ۨ_)���G��+���F/c鑏s��/��۽�e>�{��n�� ��eo�p�#k�C��n����?wF���"��;*������<$����d���˺��3�}�ˏi�~7��ju�`�#�9�z%�E��j	�/h�{l݅k=�����u�Z�5٥� 7����>[����h��7q�I�(y��:=5����@���#^u�9��?l�O���F.��~	�=��� �n��{�!�Sۻ�B���]�ូE����������w�z��A:�W�SKs�K�sďt�*Z��;��������[�I�y�w�o�9�۝t���(�-}��鹻;�o>�un�ũ��?d>�9=[�P��=���z��/�͈nA
���C(c��3ݵ��� �s����8��|��vP5?���Ys�p"���Â*#vD�l�Q�x�^Z�J����,���<.$���E���I������-��KK!.(>ݼ��C)�����w��뮸뮺뎼x�������쏫&���fO1Δ7��I2@�EH1���׎�:뎺뮸�Ǐ>�}}}}����
 T	U>7HB`���$R�����뮺ۮ��:��Ǐ���|�7��Q�p�w\�9��*���y��K���t����$�#O����_��[u�]u�^<x�������d��wv4��ِ���$�t4c3E��<���y�9W]�J,���ok�/��,&�Ld�{�t��L �3���w2l˺�^u�κɳ��&��F'׾��Ҳ�{n2C&�廾�w߫��9�.]�~v�J(�v�`�{뇫�z�	��m��l�=���hm�2`LԈRH���Ym���ҎΕS1��;i�����:����[h�	����cӿ.�̡�3x�nx���W/������ĭE&�meR�Gh��ɷK\��3��1��O^���x_dae9��ݵ�EyCA����-�&nn���a:�5c��w^����utt��ގ:���>��C�"4�.�dY�	��cG�.�at.�V=a:"��_n�W��w���;��]�p�jqa0۲��Z�wN.1�!n��G�������N9��!��X�=]����n0k`�o7��1.rF��NS�˦��O���޺g���p���tY6.#A�n�7=�;����'q˸��ӻc��Fq����خ��>��=��nR��vӘȨLg:k�5�@�M6�p����R ڍ��b�\P-�&s���<:'�n�Qlm��qv]�,q$60���ۑ�n�p�m��׭o2�x[��۴:^un���	����l�m*����#ŷf��d�f�D�-��fm�`ڒ�kƆK
\����c0F�=a��]�-OU��ܧ nӸLZN��a�Ā�V�GK]s�Fq��T\[��X���Ę�ػQ�1����ګk@�ʂÏ"�^N����7����vG�c��s�9���6I⢷�V����u�v>�<5�U۱��ϰpUp������E.pqu�e��O;�����W[��Vnу���V0=���hM��7�3�0��ێ-�����Q��$�ôQ�o�MC�}g){;%p0bШ[P!L3mvs�#��)'����6�7d�5�sp�`�M�׵�WcM�B�65oi�'8�o;���8۲�^�l��f�U-:�UTm@�W�.���6�zٺAn[�ֳ�ef�e��'��Ã�ؓc��w�vu{�M=���ݲ���I���qt���܏˹�Z;0Ptp�Fg����G�)�VQq�iK��_"&�b���(F�-��Q�����ݭ�n��mo�2dɓ&L�2���QT�î=�ռ|����wi�X����.�-̮�J�q���lc-�Faͩ�r���l\�^��;����dĻ��i�1�M."kB����m+a#b�ңl����@�&��Q����u5�;���(p;��V^Ҕ�Y��3�ѓ��۝!W�h8��hζj�q� �|�帴w4�ܑ%кl#�}��v�ƜZ1o���Hʛ�2`������<��|�~�Z=H��iv�Σ�]*Ѯ&��h&�I	Y�x.R� ��?#���\&t&]ش��}�J���'��rW����3ؽ��C�]�
ӱ�����5H@#cfx�D�d�PKN�>�}��87��N/\�{�3���v�Zpً��a�q���<��Y*�|ۺs�ʥ5���$	ȡ�UY6��d�Ζ�k��!T��&P1�<�y��aM�������=���f4Wd�o^��g�o~;�1�E��SL�Jv-2��e�w\{�\��t�zEmhܥ���W�a�I3�BS�	���'�N{oO�1�']n���XRK��n����t����\q��(��RB.\�X����i�.��'�/v�Y���s^���9��iBb�V��TT�>���;0���z��E�c��&9n���o������}�xc*A8t#�o�����aCb�hP��^1߅y��ؗ_�ւ�i��i�_]�7N��Ol����`�"3�T����5�O�˨T�%;n��d�J�4�LD�[���ox� ��X̥�]u<�5�*ffy��?D����1��މ�޽/����2�xb��;�ByFZu�e)b�c̯J�\���:�pۑ�jyz�Tw�tW	�l�5� z	�zY�%�'�U;��az|�KXJL a�%��t����x��S�b�:�L1�2�k��~I���-8~�M7z�]/z�9�Gg"d�J�{P��gk�.Pv-�@oz�sͭ���A�z������/پY���^n�j�2�2���nV�T��a�7����H;�&��U�?R������[�2Bl�fƽ��z��g�[�j����g.o�?<K���o�_μM���T	:�"�[�2dɓ&L�7�8}��;��O�7�U�zlW
�3�3�Ӵ7��	�L�}�э�����us�_�L�Th��;t�뮦s�RΛ����T��>q���M2�g�jW^����������^|��dūVd3�J�1.+�^u��z�Xe�=.�.��%�E0�m� �ƽ�����DC���b(N�f�%Cuh�L3&L���Z����p�ݕ�}.�{ɨGH���J�4�3��MK.�*.kln����W�݇n��uʹ���&m��b1������K8i�jjx�Y���H3[*�ܮu_�/÷�6ۈoX&�BeC�����[.-�*�*���ݛ�{�*xVP��-��[=;CvP��/0��J����O9�E�3|���}z�<�+�l��~�8�h�N�0�r�x F��M���Ny���[����|x���M4�M(��gi�$M2��1i��b+=�>�[9/;�y�uʹ�]�mL &f�Q������o���\8�Q�+F���=:����]��Jt�s�����S��[D��B�oK�����Y��q���#���$<������ ��MT�U �s��f��B�[q�[��{EO���[M�⯪���GQp=H�A���۞o[S#�_��67����g��ܻ�X�/7]y�uʋt�HL��P�cR�jəۃ�K{p46k�(2�=_��f�ݯ+������w��4fFb��|�^�1��	bԪ��#&�XތCs�7u��h��y�&V�f8�ް"�Nݏ�,,G7����෯�_qz�{��wҴ��G���N����M�䣴n����l\kʥu*�/��>I�/8+r���!��m̙2dɓ&L��KXu_8~ϫ�FU+�<�g��'	�Z	)cA��ȍ�[+s6
������	����=�J�m9pڮa�6/ݞ��n���ۛu���d�������s�s&&��v2�.FY1tJJF�F�4���n��hC�����\]��\Z��J�{q �z��69PR°�LBV�)s+^&�)����Cpz~g�=3T���n���f�t�S�w:-��^Fw�v������mU�yl��
�f��(�nBl�&�0�:�a��kvH��bW̏�h6c��z��F��^x��{M֧�}���&��[�.&fg܅=�y;B��X���۴}��o�Fw-z�jf0�̆v�cf!���HU;?F���E�@�E�$������N�̝ml��	�gi�&c��9x�D�g�N=7�2P��s�w���<]r�DS=�����q��T��h��&m�0���y��39� ��g�4���;��F�|�3��]�2��U�"�n���ݶ���N�sRx	ixƊ	��g"�WKƭ9��h"�\�ު���1SP��ѨG�堦�U��{��</2t>g�\>��g��u���	�����*3����<1���p�y.�1�N�f�u4�"8����zv�x��x�n�y�f_q���?�[v35	�jW�k.�׏֚i��i����~��6Z�p��gT*��U�P��UT��;]��5����-2�(L�Ә�o*_ɹ;��ا��/��ԛ�홏�!dp/�0��֪q�)�4�S�z=������3̨��߷Ѵjx^S
�Cb���dl��ӳ{�ud�we��UL���\i��#����c7E�ҫ�r<+�32���T=��l�/�,OE�-A��)"�8PL �m�ۉ��z��I�z�@H��IFeV�˼V��U����aT�m��ժ�m��ͧ�
��9��W��Be	��e;E1=�8�w*9�)�q������5��d��ހ�f�Vׇ�Q���mp¼��m�gj����Ʀ�ry�K�Y�qM��6h��AP�@��T�Y3��>ޭd�С|
����蘺�������2� �J�>>y�ު����ɓ&L�2dɾM��`��_�J���?5D�CL��&W��
'�$���L���1|����;�볎�k. ��L�K]8�$�HU)�����>{�ؽB���3b�G�f�gd2��A}5*>�p̐r:�����8�)K-�(fe�.,�����ƅP�Xlqq��4����|�;�y��>v�T�G��J��������	����F��P�^��\6�5>~�?`g+V���R��{�x�mMJEx����'�t&1j�Yi =�$"��S)�}6���� ���u���S��g3כz��ݽR�m�V�z*�j)�V�+j�w]T���>~[���i��������)�pׯH���a�oge�z�;��YX�v,��x�L����z�ޛŔ�q���'�9r��@r�p��2dɓ&L�7�~�[HL��e	����3Z0];����E�fw_,�=)��������;~_l������v�s\�n�M�e�,��U
ha��Ç�IBt�$�\�g�:��7�ўő�T��8�b�/������2��� �A�2���e�,EL7
�����M+��/<����إ��ǤJ�� ��bm���|�<�."�Ǖ���Z'�=v��y)��̾�k3����l��T�Z��d�m�Ǩ�y�<�T+U��{�#b���r3�)�/��vI=9lfSLCkUH�MT�4�I�7s�Wk�U��@߫l�u��<��x�����>ǌe�2f�>S���������?�\���;������Շ��	�!NvV)��߇�i����~�������x�O��2dɓ&������6z�)F{��8�����8�zkوy�Y$«4�۰����kc]h���c�ZN6㭶���^@��2��89�6��֔�.�;7l�;'-��ojۍZН,�����.n�0�yB"��8�-����u�y���.���`og����vp9Ã�]{t���>�}ȼq�*JI���mAH6,���]�\�}�s����P��˼e�潾�W�y?v��쥮Fm�[
8d6���1�
,��cx!��L;�.�v�͕�(!'�!׼���}7�&Pg�k���h��-fmϢeT�����@L�i�hlmyB�����\���~I�r�������p���7r)���m6�'u2�]�mU߽Y�̱��ໞ�NՓ>���W����2�c2���mI�<;����� �+ԦSvgg{ƍ�k3����I����ۛ(fC�%4�L@��&\�H>�M>�Tbc73z.�w�5�W��sb��I�3�t���u޷&}�/���/'�+GV�u-Ʒ�Z�^��+f0���3��"A��8B��399p�zR��\��Y�1�|��ɲ�0�����iy�t�s��(E��{�{79���7��<v�u2������O�����B��%�
ˌ��K��G����K�R�{^or5�7���ɓ&wgggf��G&�@w}���;�me���VL��y'K�H;��n�~gi��rh.�d� �W7]�y��V���[j�:&`L�3 ]��꨷��!r�U^^K�����j�D_���m��g`N�c���ñ���ø;���gIlT���hg�Zˑ��>�b����G�����O��)�!�����v�Ӭ�+����/�Kùb`9�R��HI7^�4�|��*j��{Eo���<!��%Eq̮���5�J��!�S>z�}J���s�4�����ע�������[�ǲ�˹����{�M��&�!TZf�Z3o�?�q���Ep�Ѱm闦�5���Fޯ
���K����Z�5�-�>��� Im��yE�S���#}b�-�L]ܻ��2{��[�[�g���G�w]?�3��矰&�����q=�������׷V�yk�;�[����#���{���f�}�������^�o��t>���/l#u�'��B2W*+��F8��b{�u��c�?<}�7�}xI�=��Y��6�S�=���6�\]ۣw{�ؖ�r��s Є��P��X����G�Co`:,��=���93�J��rO�W���������Ō����_z�^�SR�^�l�Ж����ٿW�m��¯�p����gK�Y ��0���w�/����w�l�����Rg >.����q}h�'q2gfh=����M~��y�/�7��l�����}�f�?`��՜Z����C7xC�X�}XC=��\�݁�$�{���X��v{�F�6z{ޝ�v��",ɍ^����>9��q��p�����u����n����{�\>���'�0>{qL���`�=��=��RN����x��r�jɗ׳P�P4,;��m���8�\)'�w�{r��x7��<�_%�ݏ�v�����-�4]�<�^��ALtS8a����]h�wgLc�c�F�k�7j�r��I�`�^#��<2i��AǤ����n6���e��i��XC���o°en�H�`#l�	(6��3yf�`�E=ܣ��&P�̈��K���u		FH
��C����ׯ_���뮺�<x�������{e�7�ػ�#"�CD����s�)�y�o����뭺뮺�Ǐ<x�����{'�Po��Fae��Φ�ݺ��Ж#>�M������Ӯ�뮼x��Ǐ�����$$���r��1�$� �%>w1�wk�tC�iǏ����:�N�뮺��Ǐ7���o����_�"1`��.I�>:��s)����G]r���ܻ��R��4�ۦ����E���rRY�
$a�H�b�~���nI4$azn6 wnI��:�1	3{��P���A���#xܹ�e�] Q$�c4RC)	.n�s����(���������5��2�kt�bl29rLc�\$C/;���"���FFK���u���n�m��]��II�+[�'I��o���ͦv8�S+,@�������������j�o����w��=p�N�)>����kj�{({e�����z�v�E����F(��/c���C����� Z)��S)�ʊ���4u-JID�v*;��5�ۉ��j�c��'%��$�J3 ɿ���J�J��~_�;Iݥo�b��H�, �=C�$61��	�h�	�:j�Y��O�Rh�y߼��GM�N��W��t�9L�z�]���AR�\��@t�f`�i����LF�s���4��{U��`�}q�a9i�g	�;��5J��u{I�&p���>L�W�����R�˱[�Ko���e��T���U��]?X�?�"���1&`��\�N�di�O/M�]�-�_S���^?po�¸�'K�����/n���7̙2gv�n�m��s�=�'��_l�v��J�I�N��Q��϶������z�p���Ҷ)�j��>�����$ϐ.]���b���%v�/v�J�.x�4!���39~��M��~�|���ۚ�Z8=�}q��j��q1I�H�4��R��'�mF�6Be����9���Պ��Ж�������vx>�Rۯ�l�~g�=8���JL�u�w��Q~�X2��e��^��h��z������F�܃�Z�M2��1@�h�}m�3K{b=b�&�/���U�Ez�&v�틥�o�V¡8����Z�Wx:��[���<��݂��<���{��"(��hw;&�/7�z�1+��E!��G}���M��N�v@7��\2V��o�~}|i�m��۶�l9�}ڏ�0�Vn[sek,�A[�u�e˘֛;�����+aquqZ���.�p`��d�XN��;h���ɼ���)�#�٣q�AT��q��4;���LE�m��%���s-����/���Ĺt��Y2�5u��)��d7��b�ł{n�d�8��V�P�p�at��+�N$�,����\zQs�f�"Dk�{��ɺ��[������ؚ�5��W�ض8R n�#
�;\���j/���y����|�L�V+++�%�k�3��NMn`/J��Mn٪�S8���1�X���]�w���+pҾqg�,^UR.�Ѳ��~m���v}�p�S=Uy���Wq�79�<Ui��z��#��$n�nU;URg��/�����``�0ʆ�:I&���U,����TFɮ�@�@�}��s�E�n��"�N�Hy�̾���ۻ�N��ޞ�5xJ�4��=�M�p�L̦��l�����C�Xl�.�1��:Z�*Z�]��5�m�[-n�\!�����.�]�j���9�W�v��t�z�Xy�}8��I��kj�O�|�#�Nw��H����WF·�(vv�/�����h ���v,���O�?+�n]������?�ӽⱎ��\������l��l-��i�Ϸ�A�j²���(x�5��W�+�	�O�h�3�6����$�vZ�X]֖Y�����^�7|N>S���&yp*��	o2
a�D��.%�u�d��3�p��s��؇��_Y�)~�x�p^E��m�J�03(8�]/>�y�q[{gm�����$���)�wCL��Ì3&\����!,�Æ�Ʀ�B�niMr���y���^i�&�(���L�yP@�Kw������k����5@⎪�ۘp�Ȼ@]��Ȏ���"���ݭ�����﷏w�U�/��u �n�Ut�����s�������C!-E
��W������x���X ���~K܆����yt����f�x���.)�8g�e�WL;ٽ�l����&M󳳲dɞ���N��������+���N��dW�3���yJ��8��ޕ��4S����os��y__�D;kEP�X�#6�C^�mT�*�J&f�^Q�A^�s���(��_��m	��U�{~�����iq���;F�d�k��y8WHG��w�om���R�D�+��v��Uٔ7Σ�+�2��ۗ^�@?z���i)��@�����f=�q6J���5���*���&��1
&�ǮtMw�F�-��,m�ީ
������&��һ�#��]}ü#��_���i�T��@�wq��rtx>��8�p�������\|��h����S�k]�}��/؅ݸt�^����/��*�^Y|�˾c��q���6�)O��-���ܢ=��qv���G�*b4 ~y����md�9��w� _"�t���'�G�L���]�i���97*�4BS����e�r�7��m�Dx� N�ZŌ�8I�R䣾�x|�*Ï���m��i��=��^i0�a3uH}מּx��>gi_M���v�TE���͕,�fa��c��%`��,��4KF�v���p�n�ڻv��"K�[~|K�{1�od�L�3�j/�D�����������v���{�L˙@L�P=��9����W
���;��\�3޶Jm�<�Uu8F�s��t�W���h��T��Ѝ��;۳���)���]Uk2"�/��&vʐ�2��S�w�=�l�C<b�La*����/���v_Pu{��A�=��$�x�^e	�d�+���\�u�~G��c;�<�=���ބ@����x:�"oLG;��|�#qb.nՕ��;V�Qy��ȷ����u��yds��osm!�A�/��.�ގ�>�w���`��yF|���%��6�4�M�l�����̽u�c��k�)��Th�t�l�LEUi%��c�Ku�Ju\�r!���t�E�;U/�����+@��v#Ap<p�{n�Ԣ�#�(�Jn֮����,v-�u�ťKq<x{#V��=�2BC&6i��q(v4�{8%�FV�	�2��3.�9�Ǉ��:Wm��+^�5�c�%��Z�Lcm��?_���_�P~!>5cr1��^�����l罸/ =�S.������6��N�n̓*�)�6k�s����3�S;r�|��C.�.�툨���RJ�l�V6uՀ�Fo9�=T��qv�Q��&�ɔ��}�]��_�yi��9�I�|���~���Wj�x����4���	��#��mx�7��VfzTW�0�!�%�,��w��\�j�
���v-�*o7���Lb*�ewe��}���^A٠E�p��=hL��C�W�U-1�#��� ���=Q;��T�//+��Ɇ4w1h�]�y�v�ǧ�0����r��7ƷsP�� �Y�Q.�ԅ[]���|��Z���aR�L�3��혧����bfE���̟1�&Pi���f��3�E'��s�	�^��b�
�ziN ����]�S��4yPPlg�s�Y��{=�`|�X��ڙ��?�ko�2dɓ&wggg�K���e\������\E�{��Ïf	���v���JS�!M]; V�2�1VD(������A&�W�b����/.[�Sn;lL��\SP���R�P��!V���el��w�b��N>y��X�=϶�-����fa����UT�+�'k"�2w�wK_���o���|�cn]���L)�����9¡C����<v�r���vz�kijl܎+4�l�y�o�w�x�T�M��{���әs�g��~����_�}f"���3������w�	��VKN�����עw��y��Jy	��Z�/7lER�@z��S0�fWs�t��Fz�x�2�k�駥�K�16��=P��0��M7�9s�^�l����h�Ny�,�]������dɓ;���dɝ�P$�i��s�{�����&���ʯi��]�pp_�z �M1g�g������)�ӗs��)s���e�n�6]�e	��I +��C�j��־����K�׷�/g�[w����MW2��W7�<�g�j�Y�	f�xg<7e�TR����k�:������G�7�57c�$��p:�'��o���y�h�e"j��|��M2�	@H��������3Px��3�5���T�߯��ϸ����{Q���u�{v*���.��a1幏��ۤI1OUꘙ�oYZ�@�2����.��3|y�Ч�_��9_+cv�O^�;�{_)�{͇��lwZ��t�+�Q^��sS�.�[2fy�|�ؔ���;V���30{,:�/U�s�m��K����˞>�q]�5ݷ�*K�^�|�!}Nb�?S[|ɓ ���2d�-��y�����������:�0X3�˚���s7uM}�ٮ��JcuPTj~Ť�=ܼ���(�t��x"yIW�ܨ)'vw���S$��Bp��׍r�)�i��4�oUb��y��oZYz&��}Z<�ع�e��2�ey�G�����[z_5����e�߻ۑOs�2�&�p<�P�"O���v�ML��M-���y^�D��(��צs���wW�Չ���wb��S<����^w����x{I���y3TK?*Žzf}^޴��|����n�1q�w����i��Y0���Z�V��b��X�3���[�9=�WD ���&hb�O^���sPgǿ���R-���J��6"1X/�A��_�</D9ᒻ�_�}�9�d�v]�w&�c[sR^J���a�ɰS�+��=�Ƿsb�\�����:�%�p�{�̓�F���=�V�8h%rw��N=�>�7n��[	xu�w�׷��Ֆ��y�;"�r��$��׽�Cui]G���\�B�p;��_Agc��a���|1��8W�������n�=�v��W,>�f�K{Վ�r8�-Ӟ>[X]���n٦_Y�������ޕ������x��ޏ7�ۏh;�R��!�����>����]��K�s�sԼs݈��ӯ�s}.q���
 �C�x��!��^;6�={�b�p����H�x��=�Wo��|�qX��|u��w7y=\W�W<��ò��dm������%^FS�=Y���Q�\��h�ɻ���{�o��t%�1{W��{��S�����~�}}y_u��Z{Io��wL�o�t��:ez��k%�3�`�u^�3�;|}8��6���^�G}�7����
����Dy-�p���2�#}�s�2=�)w���?j�/e֧t#�sΒ[�l׳��&����/.��/��][ݻ�T��'ɜ`J8Y�L(��L0���Ĉ	����5OR�=��!'.=��$��f�+��<c��$l�3�ۛO�9坳c�Vs7[k/�����@=�w�ǚ�*r(���ʃB��}bX�BM̓F�Ɵ;��[,�L����y�l�1��>?_]i�]u�^<x��������7������A�>ur���*���ƻ�\MIoJ���=���������]i�]u�^<x���__]��[����4��2�W���^��l"H��HJ����>��>��u��뮺��Ǐ:�����h!U!QJaP��7ۣHi�!��/;�W�t��u��R��m�����_���]u�^<x���]}t�$���ILa$vy�±Q���Ҹc�[���Y �nW"�����U�0X�$��bA�$�ﺃ_M��RccEz�;ή���4m��}5¢�
�L�C �ںst7-�zsE�x4W,d&Y#�ٷ<q,H]v�*1x��x6��,L��&a��v62T�F4��1���7k�oM�m=u����cEI\�k���6�}�x�7
(Ɠ��"��e\������}y�w�� &L:(R���8�/暺#��w6^v@���5T�:��V�F�Vn�X�ہ	���ܥ��6�r׭;�x���MkG��n5�9)���F�ȏ�Ƨ�cb5����Z�Y�d�F�<��ݷ,j��S13W��a�ƴ����e;��->{ڞ	8���A��v����h��Fr�*XL�7Rt��ͮ���YQ	L�f�֓Dk��=af�2o<$��8�;0��,�i�U�pT�h]��fv&�]3L�<�ֶ�Ek�tQ�4��PѴlb@e��nVR�rv�7�-:�(�=Tc9��{m]��Ja�pݞ����f��4C��.�K��[ϗof�t��/i8�ë/S�G���Xx��X�l'KYk�W�u���Fh8�X�mj�Z-�hmEƼ�.���c!�UA�&�e�-�]4ti�����H�&�W�eq7
��	j,\��\s��]�R��D�ڴ���/1��P��6��9&[�a�;v+X̙��Fwk7�汇���t���Yه,/`�nɻt��^��3��]�F헮�\��4:�$�=�htnx��%�n6�\Z�Ě�[4H�y�X�:�CD5v�r�;u[kv;0n�0U��a���XF.�h��l����z����ZP���&n�m�m��V�C����ڽ��L�IB��`�m5p��G�@�U�d��h���mu�]�v�c�v*��02d�j���Hc&��Ѕ�˦a�����d�K��룍���n�`c�$}q˩�Q����7Y�u��on1s���Ί�&:�Gbq����p���t�f\t�k�lh��s����Ʉ�r��w\u��孪��i��ڋ���,^ V�XѲ�4e��q���e��� ݊�a.\#�;zvYx���j1r��n�k-�wM(J����s;����GG=�܍��\i[�o!>+�	3;*%WKy@��Yu�,J�X;�v��٦�y��Q�:[c*�CG,Ma��_��;���3�;;&L��g�_w�uD�B���\��G�g����/	cD3�̈́�m�!g�og�#��YY��8��*�Gn�����p��CRf���s�Zv��+��.4����'��y��/\Hm��-ꋞ^��V�����G=��<��'
+��i\6����y� �� �v�h3Q�t�ۖ�șm+��ћe��o��Z���y����"xw�}^�s�]�kj�����:�{��e"|HكY�*	��Zm����!�12�I�4vK���{ӛ��_���лD{.����O��~ζk����%���%��~��\��[Jk����&�B.���Q��{z�q��i�o*�P_Ǹ�]
�[ɶSkU=R��3c|'�%-��w0�3�*/�W"/fa�P�����UKoD_x�e��m��i��9�U�v��U��	�ݻ�3�c$�54�����L���d#	�����_s���~Qw��0z}^��|U6�W���u�y%S��'�!e3����c6��ԭ����+�ؗ5�]6��'����%�y�@�[&������T_�F�CHW�LX�}��v��4ˇP)6�����(�O��%��u����[@�3\�A��n<�Ž�>$�{��>�b��v��qCވ}m�;&LX��L�i{�6Sw�}?m��`�*毐�+>�3�=xJ�܇,�ii)���ǚK���"���zu܇� ��5Yc������O�m�2��������b}�]��^��.+��^�c����^�ql�  �Qb��x��g�jj�j�
�Yڪ��1#�7�k"-G^Q��>�ɛ�9�co�U( Uy���������~�u�)��ƚj�U�m��z�;/0��tWWC��'q����
�'�	�۽[�=3^��_/B`�g���"�ݹ�`[�����j�9�Ȉh)�te�~�̮\�����&[	b"@A�V�U�j�a�_ۓ�P&ff]��t�}o�TĽW�����&� @�~������(-9�\�f�-g�{(����~_�HیI�<��&k��.��C�K��1b�2b��/Ӓ�q��;�>̃쬗|��- �u��3�S�DV�P��k���L&�!�՛�353�Nf��$�L_�lD�G[Cb��rA���X]�jЪ����ج.���8���W��޾��� ']��
�g$hx�C�:�BJ!�w(<�<������9��+(P�b!�x%�b)&�X�N��=:�|�{gݰg+&�����6w���8PobjT7 C܃L��4��Qnh>�u��<�UZq�}�6�����9���6��Z���'�@���i�&j�&i������oq+� ��Xv�1O�}�ބ���Uz��f{O�
������fL�C�v_=���9Y0/��oGD�=q�Bg��o��~V4`� a|�hgu�B���M+���UT�y�rȡ8Ʊë�dT!�j@8���I�,�&M��&�;���i�2�`g���x˖��"�����^T�Wa-��)��;G;�S�Vp��?�D���.�Yu(5�4y���1Lc��L�GZ�4LK�7�����'���6�v����E$9x�uVǩ�+)�"X�BZi�U��ye�1��J0����ϣ*�`Wp{Mm��U�os�L�	�D�;o]߀�e�n���V��2�����=V34T���w��q
fmuή9V=~q�o`H$K8=�2�ޮ�1��i�©l���UG��&S;2�i��� Cͮe��~z��G>��ɠ;�մ��7p��i�s�q�D֚I�/;ݢ��Q���{������^�ZSQ�8v{�"�ޝ;���U���J&e@["�5����4��Qh:l����J#�o�� �d�2��i�ڨ���x~�!=�m�3�;�E ���YÌ�`5��[76����S��G �"�S��n�C�x�oBq �t���խ���$�{Z�9�v�]O�ss�܋Ӧ�e�&Y�%�Z���P#�]��ݗ=*�M����i�����Cv�A�-lf�I�;�I�C���l�ykJ��+V�������7hI�����+�Yx��q��]"����	����S~�F����jz�ҷ�xwZ�&s�W咳a�O��O�<�������(^�gl���hᙦ�ݗ��1g�B�4��Ymk���9,�{��v�^�:�֮�1��rqp�!H�T�N�?w��O��naSԚe�L��&M�S���qO�ӗw�VWEM{��2�%
�kvf1�4I"�����m���1��&�qT�y]�ѓ^z�%�!��$�������⼄��g�v�"�Sv$�x��<�M�b�٫=Bo���Wc>M:O}9�=�ӿ��?h}�����+�z�.͔�3�<qc� ��L�ȁ?�g�?f<��m�o�ͯ{�FUd�u��*n�鈱؆l��ȶ���m��׌ƿ�.��]�j�K�z�2��;��r�&{�����Q�~��ߧ�tmg��殃����Mt_c��4� �_���C�����2L� �2&@��-�4�{o��&��[�9�)�����R�P�S�uP����/2��Gt�v[_nd�x*he��3��\&N��i�j��]�ig%����D����o�/�*�����k�R�C�Y�*\ʙBfZ(��X�V�!2�m�޸�څ5�M�}]�Jvv����7?P�ﾗo���m���Λ��M���b�v��q�]�i>oK���0�������ߘ��9,��6�v%>���d޿Y�{�,��i��i�1��S�J"��o����هͿt���ʦ�L�vdǖ�̓�m�ymo�z���w�H+.o���C.f$���׳kmLս�{u�lff+�¿M,t�~9�N5E�~#�e�$�/ 2)��[��Ʃ��o$'7�U%^�:���M^y����h��U����Uw�9xP��M�@_;<�c+L��ħ��2�_��3+�w�]��5S�SYp.�h��vdB�V�����nz/%h����H[k#�U!�w-*��=h�!������u����V��Ĺ���`UظKC��:����$��6{Z�Cz��XL��{�&2�Uo�y�uxf�|6u4�&�vv�M�^z���b
�Sf=����dշY��nx��/Eu�9��������ѽu��F��z�-T�T����_k����.��q1Q��͕��2���ݸ�*�T��Hc�8�j|�X1�@D�CL�n��:T*��TY��(G}灾�����x��"l���g_�����=�H�^��y5�ڮq��ڣͼ�Sݽ�5xs�,Oڻ<�&�{y�A!�;D LX�o�&,@DY�-�V&�jf�g��T���_��ɡ{�9��]�Ū4�̦������������[�եA�n����c����X��	�k�b!���~�*I'��܈cv��=}�s��k3*����3��s�{�w}�LټN��$d�w3 L��Y��ђ��Jk�^.��z��`e�L���؞׊ܽ(14Y���Xx�� ��k�eL��n�f��A�p��w܁~9|o2��(j�'u���HUFX�*qqe�s@H��M2�U��m�N��e�wM���}�\�����F�([U8�UC�X^�=���|���='��G/G��ͩ��U5n�iC�zj=�=��G��=�2o�ؼ3c��wu��:`�������(��~{�9�c�
�ܢX@�1bŋ |Y�ͻ2��3����Ϩ��1�7"�PX�D�B8\]6nɩ��CW"�`�!x&�u�6�,��n8hK�:i4`�a��l�m`�`C�c�6,��ᮠ�ŎbsXd3YY�HKxLY\M�bZvz����ؤ6�e���.�Z�pѯm�$�֢��ء��N���`Sv�F,p9�4�mқ
폾C}���E��>����!�ɹ�N���������=�l���hGFKyA{@){p�-�/PNT�xu!K�.�
h�l��(L�ht��>����GF������o7S�&��p�g̞s���p�6���}��9==;��˪n�L;a�}/UF���j��}�;IS*d���
!�_`;�N㏪EͪO�X�.#���g�Be3׌��W��5_�8��=c|6��a��vW\/7V����uN#���Ż�seG�������/�%��*����fe-]�Ǜ%�	ol]�.�m�7�>xu^���	�p�IT��RR6�Yh��$�B�T�E
~g�S /1R�6�nRZ�77X½7Ľ
/De8�M!2��UCU g��mz'�˽+��U ���s7�&<�\_� ��w���<G+�[��9T���Ia���U��&�,��_K��˅�o<��+�@fL%O�1�c���r�L'c��f�2������_6�k�C�H��[�S�����8����+�i�|�:9��X2h'�M�����W�z����uS�KQ~�r�yt���Z�!�q��γ���U�r����6=��m���HL�1���1�Ë�#|�w/V�7����\Á:����R�]���t�"<F�М��!C�" D�(����,���4i�j!$<:Fnk�f��I�"�R�뙎}��1yu]ɱ��?Qz�7���'S{��i��i(Gw�0f�������նr�_b*���V����f�պ��$��斥;ƪ�R��1�_��*y��w����<���z�YH����|}��vp�pg�I�pÜ�/S����y�r{��h~ہ��[��{�y����d�ʲ*�\�Yo�(^6zX��I�����L�_8?Λ½�J�S苽�E��z�ٳ�k��|i)�r��M�������	�qK\yi���<��u'�)!�y���4o�Q�[����ɽt�������7�8c\��s���I����3��/�u�餏v�˶�N�L �"��ybݷ;�l����+�J��H�oj�y��܂F�Oy�Ì�y�g���-*��:j#��E�ޕL��[��}�<��9B�y���Ovycl7�f'�j�^��q���xg{h�{Z ��olȒ��>�ǜ��ޏ�3��v��ⵥy�}� ��M̘w��]���x��K���B�6�����nx�"!�O;����o(���f���;��3��K�{����Ex;����~å-�=���3�����U&�̑&s컴��M>� �s��;7wOYp�3|�Ή�ۥ���7>�~S��Q��{y�C�%����!���.n��sX��n{�-e�v?a��=���ü�n��g�Jy�Z�}��q��ǂ����k�ׄ��>~�ٺ���uC��Q>�weh�I��'o�������xc��N���Q ��lf`�)>������ySV��`��"�����=w���a�,�����z���_���W�ɬP���6�6�F"����-���zZ��b�!�۷��㯏�_���]u�^<x���]}wbQE�sQ�M���A~�BŊ'�p����I�����iǏ�__]~:�]u�]x��Ǐu��6��MF�r�-r]�Ǎ��M����{tcTt��7{ݻy�o����~:�]u�]x��Ǐu���2Tci��1��\� �Z��s&�F�W�RFI'�[mǯ��������뮺��Ǐ:��Ȁ|!$�A�FHF��4#$�G�q�D�x��^Fwt�\�x��ΤN\6a��%�W�~�$��W1Y6"�梌;$Ѱc%%+��ڹ�p�,mE%%�o���+���d����;�1��*�ͺ3}us�e�Dm��4BB��}�b��&lX�o��}wlTe�4TW�q�V�b��=~
y�fffo��/���Qü6�fb��k�����
g�Z�v�T�`U�/+L]G1�Ck�֮#s=��Ν�YU��h#��7s��
��mB	��	RD�tmn���C�3���9�/�]㕣ކq|�P���*��|
�O�}�;�Ý�q"��*5���Ɔ(N�܌�ŀ4�iy�r-�9���O?}�mW��v������y�+����(>���,���p�P�@ST��� ���z��sv�'��h��("}]��(n��^�S�h�SsM۶�;JZ�(L�z�yQ��WX����9�9�޷="`L���[���9�M�����B��8��/<u�a��/;}����GTr��eե�=.������!�[�i�@WE��,��7�����_-8r��~O��䨊�nbŋ,X\��m�g�k�������\aܙ�CYmW�ѓ�}u�]�k[T�Uu�cW����韏|;�����z��&;;���(�t=��^]%N,˔S�ߦ�U���2&q����kbqv��H��u�հ�=㕡ym\K��H�(8֦r����4t��J�=Ḛ�O�q�{<����*MO5����^��޸g8[�}��CZ��T5W��=~
'L�x�OyE�M?N���W5�a�Ꙏm��i��f�x�WS��ʂ��:���+ûM�{S������B�gwZ����������©5U3�?�&�}W���2���q||��[~CiL�&rpnK.\�R$�d+攡@��~��2�K��˙Wq�K;����o�t�=})�cRD��.Ӱ���b����,X��)�C��^]]f#��&͇Ds[�,�b��D���^��q�qS�l��p���"d��R�����⎻1�rQ����R�hz@�)�����n1b�u�PK���)qg =�1Y�g.��n�ح�e�=�&ɝ u���\\��]��ۯ���?C���n��'��j7b��A��)�ڈN�~��iS^�AwV6��g+}��t{a#��WT�4��mB�D&$n�V�pcn�mq���<쳼����q��|Ah�
��j���9F�����f�����msc� =�j�MT���G�{v�NE���t曬�O�]P�������9���-5@0	2ٲ�M)��2r_#=�v��d�������1\^(�����'fa�u��`����S
H1pDcN���i4�u=~�Ӕjo+»�z�ٍ����rv&А%	��\LH�[��Wv��C=�t���|~�Q����2L�!c�g�D���q�ޖ�	�!��(��� ��Uɺ�9v�� ���!��D�Y7W!-�e0���ӱ��$���%Q�%w�4�s���F�iq��4s����*�2��R��4'S�������0�:��z�F�tx�3��{��eV�����d���*��G�ȧtF��E��wr���^���a^�J����1�B}�����ߜ���WӴj�*���n̪�U��`��_buL�|�i]����	#I�1}4��.�P��>-� L�Jbޗڮ����f}8�aR�c�W�7����O?�+�M{��:��jb��T�I�[�%�e:y/p��w��6�.qNɪ���a�.-��T�������:�(@��w,�ÈsJI�8R<ᗮ�i�Y�u�$�1
�\�@+X�X�U!p4���7e�Mh�d�Gt]D{8E{b#h�]�A�P�3 ��A���o/{��w)���٪��d�fQhoL5�5Gy�^	mǎ�1ݟe�ݸ�UPԹ���ԍ
_ܮ<�?��w��*�|��	�_��+HW6w�+c�2oý�닷:ôdFo�*�>M�$�^n �bŋ$�7�t�<D;��������5W��ބ@$��z��Z�k�+�w/3�⶙��;�#s����'�ЭЀc�0�`C�T7��5�5U�4����^�͊ �1��,�������]L@4�NK9�f9S��s��q4����t�����5�`�,, ��­�F!�$�	&}!'��ᰀ����Hͬ���;&���c߷�
�=�䒑V���r,Fd5W�<�¹�xԌ��YS(eO������'���M�3K	�ʟU42�[i�)�T���^53���w�%&*��Ud��(���5����x&�r�N�R�nf˫��1��A�܆b��3�5W����3-t�1;�j�2{gV�{(��oC�5�Њ�E��-{
���$;z���%7��4ۤ0�$ iŖ��,�qu�S�s ,X�.p)0�S  &W1J���2���-�n����x��w��:�0��f$M<��������9�C�.�w������۠�Ok��۵$h�J[Qڗ�7%�������=0�*��0&�nV�y{�T�ep!,�\�m�b�n3�i)�K8��w���;�V�{�׽1Xg|j�/���CuL�Ḓ_�i��b&�-��M��0�|�@��2�4ݑi��K���{����w;U) ʆ�|��`��zHk�la��	�7�&sy���SY��s��7�%(g���b�Q�6qg6��5L��j�^�.�茦���O<�d������hm�i�Zg�K�1���q���O�{���u�Y�����ѣ��	wŨ�ѧ< >�
u���lx뽛������|��%}�1�bF9ޕ!��w�Vh3(�T���/�Ӄ�*�p��I�v�y^ݺ������Ȭ�eiw9O��ϛ�(�Gdsƙ�	��уL�q]�:�>�jER4��{EM
��0͈�qH���M�[/q� q��{Z�s�g��im�8f�f�[(�$Ä�I���qi[��$M2��Fv�Οk��.3g3u_"|[��y͉p9�#��~n�����^xG
#�ܯ��9�3�h!���\��Rkk-�w5�Y���14�+��m�~=�x� ���c��v�= *�\�?�9�t{=����X%s�l�b"y��o5T-t<�0�w�&�;��Sz�g�t{��fpi�A��s�{z��\�Se[C@�
�,E.�t��ͥ��!$�HH���ͳ�U�u�/�[i��Qi�
�fw(��qڽɦW�V��u�ǂ��a0�75���\��%V�j���Bik��T�I>���q��J��Ub#7����k��;�=%�mM���!���zohBT26���&9�Gw�j3�狵s��=S�F7߫�۫SkE��V�]�9��7���2�u�������i�i�A��*� �����/z�/Q��sQ�O峹Oi��rC�?��ual���=+r�(y���QWVb<�_*U��ԗi�@��ŋ,X�3xO�����@�jP=y�����-�\��":8v������S*�s}A���ujb��Fw%U�ωՎz���0�c	�s�o���L�ec��l�ˮ�-��}G�)5p��f�yi�T��p5?���MF@����BJ��H��=��V�����DԢ{�zW���mȑ�Y��I��O
��; ���${z��{N��E��}��Dy�Ť�*d	�wݝ��*�38q�>7� ��j��j����w޵��ZYk��W�6�e��6�n�3����~��q�kj}�B4v�P/�T+�����(���7$���5�3?��f��-����Q�{� ��
C�ꚛ�G.������Ia ����ŋ,@k�%6�T7٦�c������%���US9��r�Ӻw"�nc݋���tLv�UYB�^  ��U ��=����z���7��U�	�SL�X�V�$����Ӧ.f��|n�.����Be7�M��~���w�NN���B׈&΋ԛ[���΄�X�uʳ��!�% ^.�jA@Wf�G��CL�ZZ=u��c��������f�a�Yjej�aT���&>��P�ZsgEFwU���ɭ;N������.��K�[�1�"e	��U�^nwm�x���D�I%Rf����񛬸������n��}���<<��	�����i�=ih��/�ǌ�R��U�xU�4I�H-%y�����>��g/U��i��{����)/6����
U+�A �z����b�-� ,X��H[uR�L]��$KI����>�O�.ƥ6��\�f+�����I�`!����-ջ��?t���n��Q�֥l�l&m�h�Iǔ�%5�\\�b�`����Z��KV;U"�U ;0���G�O��嫹��5V)1��6���{�L�8�R�����:��uFZ���jk���Vj=|�������AڪL(�}"$�b*K/bhL��&t��9�I���6���~A'���Œ��L�<�aWv�yyt�i7�L�c@h���w�FƓ�z^A��="+x�}ѳ*n�뺭4�9P&m�u��]�ޞhI�I����q��ǀ��\v#�����7�v�y��?�������7�I���
��� �g�O�?�� ��낊5��,�
�#õj{��efژ�K-�Yj�ki�V��1��ɩ����3jjV���f�Ե�kf���55�c&3m���j��d�U+*�3V�Ɍ�kLcZ�b�m�2�1�i�ͫLjZ�Ɍ�i����c�Z�ɛm2jj�Ɍ��ұ��ʬʴŕY�Y�LYm��efږ2e���5�Ʀ�Ljj�&2f�5��f�������R�ژ���Xɚ�X�mJ�Zf��mMFV�YZ����eZVZҳj��jVZ�śT�֥e�+%f�1�mJ�Աe�+9j��֕�Ԭڥfڕ�T�-�Y�J�jV[R�mJ͵+5�YmJͪV[R��J�jVkR�ڕ��YmJ͵+6�YV��jU�����f�+-�Y�J��V[R�ڔ�BN����*�b	��YmJ͵+-�Y�JͪVm�Y�J�mJ�jVkR��+-�Y�J�Ԭ��eT�եY�J�jVV�ejVkR�j��ԬڥejVmR��JʩYZ��Ԭ�JͪVZ�fڕ�T�ڥo]ՖԬ���Ԭڥf�+6�YZ���Yj��ԫ*�f�+6Ԭڥf�+6�YZ��T��JͪU��Y���R�j���Y��j���VZ��YY��eYY�-�������m+-eeYYk+-�e��*̭��b
�H4�� ��
�b��"�(+�*�`"���
+wb ��*�`"���(����b����(��*� Т�(�+���b���"+���b����݀ڂBͪVkR�j��jV[R��+6�Y�J��ݫv�++R��+-�Y�J�j��T �1P��-�3U՛T��R�j�,�R�Z��Ԭ��f�+*םV괬֥em+5��J��fښ�6�Ym�5+i�Y�_�{_�W��u��_��P �*����b��W��?����~@~�������������?���B����/���?����?���?Y�������O� 
��?�D_����`~������O�������C��_���@��B��i���<����� �������J$���"��ږͪm6�ٶ����JR ��T��Q��ښ��KT�J�ZV�ZkSj�Z��������2�D("	H�ET�٫M�+R�֖Z�m5iTڥVj�R�6�զ��Z�jl���6�R֛6�j�ifڛi�JmSf�5f�%�2ڕ��3j�ͭJkSe�E�,�E���j-j-���Q�UE�A@T��"� jJ���)j�ե+S-��RmQV��L��ڙ�M5ii�M-�,�!	C�?��,���  E@$ �@P��}������~� }������?����"
��A��L��������ԇ���0��'���OT]ڇ������O ���@@U��C�t��?_�|0�@T���B �
����P��c

�
��a��'��,��pPg�?C��������s_�S��@|�^���?[������~�� ?P����C��Ѐ����a��C��j����3�������K��<,��K���~��=>�>|��O����C�Э�1����?�0����߇��i7��� �/�`P~sPZ����V�u�g��!�S���e5���@a\-� ?�s2}p!c��                                       >�                   �
         �     �}�)TEP��%"�J�(�JJQ%*RT�(UDU
�HR����))Q �HPT���TJ   �P�QRED�� <|���^t�s�2�{�{�*�z����U*��G�
壶[hy�fD-��zH�uTE;��ws�	WvP   � �

w�� p�|��K�x%G�� y�  [�ǒ���(=�p:T��D���E*���oc�(��-
 �   �  }�*JU�*�H�����B���}��y�֍�Jr�%�zI�{��B�v{�HW h����T��%ݺ{e{۠    {�  ��{���zܫ����*��=�(����
������Q@ܥU+:*���$n܁S���'�    �  �*RQB�U�EH�O*�`������Q-��T3�n���*��Ir�F��J�:J��[��$r�    ��� �]�r�VmUP;���R��p��
�-QD�wUPwB9���q*V��QW6��EP   �   �ꈄH�EI*E%U)T)W�(U��"�wu ��y��ћ8��Cx�U[�
n�
EN��(S��B"����ޒ����7wB�+w� �   �� =U�Ԫ� "�B������z<"��j��q�4�9EJ�=nfoz�q��Ԫ�o3@ 
  |   8}I@IH��*������#�^X{kx�D&� t�䊓� Y��`b�]ۀTN��@Gt�E�P�z�!J{�8    |  ��>mEu�[�8="\ꂽ�sԀ������gW�h�J�Q.��s�+�΢���zdw��ҋ 5OЙ�R�L@���~�%%Td4h4�j�LT�� &�i�T�EH��4i���JJ��@ j"�ЪPS@��?����}?ڄw�����$��������W�Ph���X��Q_Q�߫��I2���I �$� BI!!�� �$�ܐBI�$�BF@��BC�����W����j������g2V}[I���^��p���70i��0�U������[b���M���d��ͫߴ�XE
��d�kL�^��[�f����;A�uj�hy�kLx��ՔrniOD�c%B�(�E�&�ᆭZte�ѫܕM��k�{n�������ɱs#�%�t�m�5��Ի+!L��U����ͪ5X2��,�����(�q��Th蘶V��l	zr���^��ɰ���m�{u�����vdD2��7^'T���X3n�%���J��Deb�Mܪ�� `�Tj$W�rͭ/��n�-0���n��b��8�*~5�3.Ɣ*�H�(�q��1�%n�L�5��Z
�3wU��DU�Ku��0�;%�ܳ7�ȫ���H��m��s5���e^ԛ����!�W�lí�LG`ۼ���jI��u&�c.�=�z&Y�vs���*�I	�*X�4��zVijӥj���ډ�ڶV)y��VȂ��A�)f	ݐf<��d�L��w)^iF�#f���\�E��M!up�j��M��[UKh�[�v���$��])��e��te��sj!j�Ycej�5�9��w��j�ʫ`�ۨ[�q�Ϛ�{z�ʺ63���a�u�V�J*֬�3@�!�e��[���M���A�!J���e��͸r�����B�V�jܕv�%k4�W�F�g�U�o��Ւ�q�Zb�KYz�av ��5�f5�y�ySe�x�Ie�m��%�Rm*�yz+���1���̄�n��U�ȝ|Rx�iyf�(,����a�8�j�ňg�y��USX�M�ua�C��h�;
�,�Z��6�6ѳ%l�g�M���w��XW��<�h��mb��ة��s[��:��ۨ�T��e���n�-6��zFf,�����jӲ��r������f^�^�Z�����N�ޅ�ܬ�`Z�`�����Du��TUk7j����4�B�kv�m���9��dv6��3�t���@�a�Kwij�t�<�N��\�v�u�ԏs%m�v5@F+YR�i�5́iU�%�e�b�ݚU���.U�7ife�kn�qcǖ ��S�3����jy�ڶ��J�A��ݑ�@��r�"m�v6Yf���5X<q��Q麣T
�B�7�)�Y�
���+_\[ʧ��DCgn�i�C.��U�l��wi�Wws&K�i�,�1"�,�d��]ܓ$�}���ƕ����;6m5Y
�i�����κmڹ+����5/*dۺAjuChmf�j�6�\�)�����:��up�jػe	#4n��X��ut�+�)^�x/PF�Zb�{6�M�kM|Sge�%ϞVVV�V�����˧�������5����b̷�Y5�Χ��aJJ���U�]}��v���x�m+q%OU�0��k.��@��T2UQ��m�%J�*�q�6�ܙ��G	��a�)Zi V��xt	i�*Ր��XYD�eQ���QZ*�s[Z�����OI�m�.��r����������DVB�a�Y6#D�Ձ��*�)R����f͙�5r�^l�	��w(���6�u�Xd�2e[�����U�����),�p5*��(w��r�,f;�f���jԡC6;��;c6b"�Oeա�R���/1��Y�깖w6�LJu��Ԣ��[5"˭ӢL��뫶�0��2#�Q�{�m;[b�G3Fm왯p���$��w6`RB�۷F���z2�T�U�;wnY0�;�Bm
-���Y�s5,�6�l0��3M�f䷗�NU1R\w��Yl�1�ܧv��[Q��y.�Ĳ��ظ�sr��zXxu۬�o6%���L�F�[	�*]��:-"���n�UF8!�F�c��9V��$����J7�8e)�{�0]U�ݩm�V.)�DU{��3YjRNn1y���}X����K�SM����Z��,��[��Mͻn�{ݥ����i���u��)D�[����c��%bQ$]ަ���QhUH��۶S��\��+u�4%�uk;��CyK.�ß;SN*�ɧ(�_����^Y���
���r��(�lV9�qaB��Jm��m�YD*tQy���1au3!+���4kZ�P��,�����ӫw���
��"ʭy��������:�e7��G2ؼ�W�=6��2��#��0��XN�p�/F�`M����bZ�l�����=�u�]�Y�7�g$&+#�ͺP���q�#��@����9\�SU�,;[���p�!�ͩ�����k0c(;���m�J��عX	v�F�a;�Z�L����ݻ5bKCx�1��[�T�;v%S��m�4%�y	����Y�����!)3pVc
^-����j�^\�+�x)��B��E֡y;T�SK%��4j����og6�(vr�:�N�vqt3n��6����E���*`�o&�
���<�c�^S�o6�)��%�
��Vm�]������*����,�
�Z+M�4�+ڧcB�KR�*ÃVI��*�-2
�X@���w�����i�V^lɁGJG�e����թ��bZ���ot:���m�#alڪݙ*$�E��ZM�{2���V/,�Ǣ���y{�n�w�\�[5�bcd�F�䣹wr)q�%0��3U+��$���/k�/Xf5Y���Z��5-�rB��°�#qf��ݤ����K�a
��q�L���b�I��Up�J�<�ߕ�ӵ��cj��Dݱޫ�UGx�䈣6�c��n����rU�J�2�o��k��w���WL̉��;�mT�K4��5U�ɶ�*n�=�@"��O��;�+rL�꥚okj��I�`�W�쬲��N�W��d��ӫi�5��D�Ր���Ϣ�#5+e�r��C�-�Z�UFr�¶�a�Z�ćn�#�e��pH9tS����k��n����pw�V��P&^0�b)<ߖ��F�WDTR`�ڨ��7e�ӹy��e�%��Fu�yH�
�u�U��Ěs$vͻ*�b0U�0ۣ���u�渪�wt��%J�fSf[�U�a��h��O-�P�ML��8��--�4�V���5�4��-F����)�Y��ˬU{���Kc�P�U�0^,m�7���li㻗��(��c.e�ZSJ��{{�;M(j�sk4M���)<�U��X5���i��R���p`���{O�T��5/�M�h��I��ٗ/,��!$�9Sla�/or�Um�X��+L�Vԛ��۷N�V�(�[1�g*�����Ú]�.k2Y�1n:�]�N^J��R�k+�b�t��̳�R���"m�U�Gl���rl�ܘܛg&n[��V��+6��aw/v��~����k
�2�wp�:w7s#S,+U�M�T���:Քszʕ�k��6+FJ˕�e>�v�;��%��Vi�#kFA�kQ�7�����T�����Q�A�A����VF�֘z�k�{vq���C-�Ɗ)a:�Pʫ��#�6�xn\�{k��9�O��U�)�s�\[\�M�ZT�۶�A͂���m�A�[�PP���.c�y�5(�ʭ���EX�m�̙"̏V$N%���w�5৷��'{lØ2��U�o\ã�9v3w6\�X�G+1�S�*s)�nW��E,&�����+s`�nU�]�B���Q<Ӳ`�B�f[F�^��IN��uE�8�iҶ��h�0���ٕ�p^lĖh�n�ϵ޻��ّ�^�FM޵����jm�:;@��Sn�x�ݿ����p�M�k�K�TUY����w�u�6c�H�S�Q��3����t�]��(M�2�n�r��U�k�f�VF�f�ۢ��XV��	
Ňn���9�3yd���01lX�٣��Ƽ�YÖc)�7s-<�"UEU�r�:�n���o�֕9��ЕR�Q@�5���.�m�f����j�]�H�gmK���L�n��d��S�խՓ1�*䡫^�dZ��ґ���ݐEPa�D;��CX`��Aݐ�S*[c6峬��{ccn����ɥ�j���W�3��/%T��V���g%ֈ��wr�L���^ӳ��4�"�s4^�-�+q`��5ܰ�s*������!NFi��V�l*�w)��˱���N/����(ʹ�l����z�Y6�e�Hti��{5+��T��h�r�rn�&��[)�x�
��Ƀj�ddU^�݅���&�`j�%�ʔ��ݓ/7dUvl�Py�i������tu�y����y4���E��=��CV�h���W�J�P[���N��GsV]4VV����VUi;̭$:�J�d�ʏA��3n����R�1t���JuT�w�n+�Vv<����ۢ���Rӡ��
%�%��T�hԛgC̘*�/���.�nYr\us&1���v�ݽL�J#,^m\���ˇi#�iܭ��J��@�*BR��NYr�v�(��jR�6�T���C%U����{*�[UL��6�]�QJ!aҭ��ޭM�tl]����_0��W�v��iߋ
�%d�kF_��˱J�IU����/�h��t�u�qa�yu��AFU�LTY0R�/f�{�'�%�f�1|˺�27a�KN��Gz�y����״r�"�Na[p��IsKC{��AL�A$�v^�vʬq�{�P�pi:�Y�U���_jF��Sڽ���L1� T�kr�A�h��Y��fC����xj���H�l���ک���*G�(텶��wF���]�Q�wlPx��� УY�+2��\$�to{E�������f�cs0�v�V�?e�9��o3��L�Zv�"��[����wF�p�&kOT1�o���Uy����#F����IHUQ�(b<��LGB�;��*��\��ܘ�Z�EU�[�Z
ݽ�7.�7�N���u�6F��%r�x-fJ�۩�p��{��t7nh���f=�6HN��ջ���6�يLw�xB�t���"�]	�6TY��H;i"rn��y���B�g�2�Y�ڀ���[�>�Q᫪;�����O!8*̨��Y�{���S?�}TQX���u������\U�L��;�J8���Q7˴ssL�r��	OVQO%�kk)���c.Ѻ�#W=ѣ�VX���3b
Y����v�M3P�Scw%h��fd�0F��F�= ���w�n�Z�yO4���;E0���/\P!��ή`�eE�q�(g�lh6�VJhƎg�J4���^K��j�ڻڻ���R�[T�	^eEN�5����	[ň1�>SA�.�+^�6�T�/&���������v����V����[2��{���ɲ6N]J�Jδ�![���p����x�U鯦�'`�wk[�)ٱM|h�Zm�ۆ���Mލ��H�ie:ũUe<�m��ٻ(қ� �n�6l�Au�DamVZP�<Ԇ@Lʩ�2�M�Y�vѯ���t�lA�Y�p���#^C�����F;�x[ڔ������U}a���.�ݕ��q�������@8v� �йU-��B�恷���
{!�N�7#���
Zduin�1ih�n��̼s7/]�Z׶������c���bA*��Y��P,᫧$����b�j��m�̽�VSG�@^
��%���uYU:��Tk%��f��ٶ.*��lʕ�V��q�mm�n���V��9Qn�����N?��i��7U�UfT��]�J�f�͍гr���a�j�F��k]D�4�5��L˗��ߊ��\P-��6i�
�Ѻ��O+2T�F�$�\�ʳ�нZEYͩb�?��/1�T[��i�}m��Qݶ�0"e=?LµSyyVE��}�T�הn���uWٮ�fq��r��*&om���<���b�L��k�i�����`Kjc�r�yj��򶋰Nk����sjYES:f�4��.��WB�
NYTG&˰�cp�ڭ2�]�Rӌ��Qm`���e�g2%[7*�R��նf��cMT��56ͩ����R�s�D�F��63fJD��^�յw;�/N+Cs͂71G����[���U�<$Di�V��k7���vU+p�{�x�ͫ�,���y��J;�kt�����F;o.�3/X�QF�zk�&P�76�	d֛�E��6V����yJ�̱��A�u��[��?Ll,�����)dѭ��?9{�J\�B�KgttJ�`�F�a.�ó2����bB0v�t3qe�2�,bAՄ�Y�&�5kY��$��h��Kq&`��!�Cz*�V���yq	�MKv�m��Av0���2%�Щ�YWj�����K6�vo�`a[���M	Lm�`�b�g2V�V�_!�5��#����[���`lQ��֌H�/w[�7/8��WQ���S�h�+s.���[ǣwsPQ�݅�[�E���s��]�4U��]�zA��*�!#-�F
B	5]�P%e��iӚ4YѨ�H��Yw/���em�D�T4+��]����d��h�j�pn��ݕv]A�kuF�AJZ�d�(ff�4֖A���RK�G�ky���
ڣ[���ղ�S�����.�	��]V�>{�/5��۲L
�ƣe#�x���!�ːLj��&�b�2�<	�D�^�e�V��X2��ڼyڝi���O3Q�p�̦kN��T:EeBm��*M�۩S*�Y;R�k4S:70,E<�1�Ű�����v�̥z��C���+	�j�Ru�WkU�SȒ[5��V�����FR�x���Zr��u�w�(� c6�0<�L�y��0m[� eS$U���G�6�n�ie<$*7(���f�ۧE!���6��ەx��.����ͷ���
�����LB�����G��ϡ4Vk�,[�YD��@�L���ՇsE9���c�Ja���늜��շ�Pz��[Y�IV�m��/�vC�c����["��f$�Ӳ(st�tVJY{L]����WqiDP��	ҵ�p���u,cq�PU�bӚ����r���;���f~�-�����$�I�d 
 A 	�"�RHE"� �	"�RA@$�@R$�) RE�!X@�� @����` �,�H���a	��$�"��XABH(E��
�
Y$��$"�I�$Y$�,$��d���I� X
BAHE	� �d
BR ���B(����"�E��R RI� �Ad�, Ad
 �(BH�H@R)$�I��$PRE�B
B!�H���@BE��X@�����$P$P$��B�I"�H)$ �k��.����*�ꋺE$�E$I"�,�!�iI	� �����ֵ����O�ܼ�]����r��+[v�I]k��wf��ԌF�E��3�e3]tMTV���@�a�[N���{��Yf��{:�ò�#z��ћ�v޹V2���]'�'@���ծ�&v���_�No`'[pG�ER�+��=ը��U�UE�^t�!-�;Wf}�V=�P���������{!���	t]��z�㛬uN�P,ͪ������,k+
�X�cB�;��
�n�u1���㋋O+e���um��x:]��BCiMI�Y�����.��=��G5sq�/*ѕZ~۠��9�˭���n��%��5>��;���dћEٹ��Xً]����o6����Fk��<������E,�:�+��S�`�"�8SV��^3�`u�F5*����g]��V��ʮ]��n@�Z�Ѿ�,>����M�0�<̽�Ơw��5:�Z��ξ:�u�z�eo�X˱n��uiWdQ*Ն�\�cl���K���ڻQ�X&�κ!�g.V�o�.�^B5��fXW:��iv�+ )P���U���.P�p>���R�T���2����v�����Yt*����feYe�9-���щ��}U�{��K2�t��~t��U/��Nqe��͊�B�'b��u�K��љ�'R�4+e������Ы�����W�C�+v���ެ�/���.!�v�����t��島��:�T��1�ѷo�gi�}ןqv��]�T"��!��vZh^��e�UX��F��t�I�A��ޗ>�o�T�Ԥ��v�Hq�V)Q�9�U�����&�{�6��'vl���B��9��k���J�תgv{O��u��1�*����A�����Z�UO7���;O�ݾSN[��}�\iЕ�hu8��8込��N�,^����_vƻ!�B������*�={ː̬��\f�6[��;���o^kW׹5�t���Q╥�/H�{�o{O*����>�v�,�
���Fu��1�Y
�����ݥ�Z�1����ҵ����G��#�Փُ�*.ݺ�#Iw�-��+n�un�"����MC���To,tMb]Z�c�;�k3�쭊
����vffNX�N}.K���]�՛@��rx�mV��q�Ճ����+����]�������v��iH�^p����W�w�4��'��1x��x�,�aP���T���j��W��}Y�"�V!3�Kj�S�t�dؖ�ԉxm�N�C���[�؞b�yD+]J�b�|��F���x轼n��ҁ��b��5h�]%̥��M�n���咷s���g}/7B���u%�	�,P��1�A�����u
^ƻ�3����/miF�gnR�xʡw��n�۾ۓ+�[��gpӼrW�M�1�&�a��<���[��^�1n�V]��Z�Ŭ^�Æ�;�2�n2�5;����u�uB���_`�t}��+	�ɻ��̙w��.u����W�2nT®��k���d�:�p�#/
�H��Бܪ)��i�����ëM�9���;��{gL�im�k?l�=�k��ld�Y}{���5W+��\/�̦�s ���Od��b�-������&�,���ǝ_bܼ[ΐ�}�hrC�����y�!�5C[�{�]�+{�q}t{V�xI��^�.���4r��c�]�,\����򷡂�ҺU�ɳ$��I��]�%�Oour�8J���ʲ5�iϕ�yw�v��7>�3TYhe��Q�Ǔ&UWݷ2�,rnVV��E��a�8�w$K�{(I�6�si��;�=��hVa��]eiXX&em�cz��ۤ�b��Wi�g�,�򕙔�)���%"Ȫ�"��`�Q�ik���d�E�d��cZq�}B΋�إ\Deݲ�7*�_e��ˍ�f�g3�j�Y{��]Z`���ͽv����y:哪���1�-�˘�����|d��:���T�k�n!4ٍa;z/+G���a�d���$Э옍��D՚���7��h(����wۨwT��`��;v�����{\8'�d��W�TU�l�n��C���KdX�nc����W�V��7�X��y��9�֝��	|u�����{q�^��̗hS�����7&����,�6,�4�#z�͓U��w�U�B�.KWt��0�kwRV'�-�,ʪ����y)֗F�%mWoY7z��W��w��"�c�#~s�ko0�ܮ��|K��Zzq5dn�ݼ6+�(�Wכ��������+r��H�za����E�S�]v���2��t��;/�U+q�e�3/6���3D�+S�$�Dt"�����R�v�,<�"_]woR�o+'[�YyZwL�i�t��gJ�;9�.��s�:�k��yC�LXm�Og�Kp���!���l'��������K�X�%L�]Kre��kn5�j��8�S{�ʳ��a+�r�
 �:�f�~%^�b�����ܥsUr[bNԹԪ��i��Ω���[����x^��G�>�giұ�=v]pɔ��Q뼝���4We���uo���eu
����j1���.��d�[U�,H,�|��P���f�*ݮ�Iӧ[}�<����ӵk��^��7f��t4��ڮ��oM�`�l��%�"��ӎMJP;ʞ����{V�y�����4ȧV���`�i��n���O�a&iZ2�9<���'}�t_����k����UYJX�j�m�۠Nݮ1IUu]�Z���:�u˭c��ޝb�:v�������*�N��L'�+��&�іt�79wIJ��ΧfsU}{�wU�oU<ܹK���U�N]S��R}��;�.�U>�j����Z��}��R�X̐;�q�u�RҎ&bN���7Ĥ+�H��E���VY��m��pܥ�\�������q&�g#tZ����mڦ366�*�)�m���2L��)�H㠉j/ܡx�V���
��;q.H'�mU[T�]��e��9�������Բ�w�n�V]Y�&�ݢ��wfs��:�}�T	[����nT��2�eb"��و ��W��+uK�S��c�.�wf��|�a�8������ɢ�S���av	�j�3�ჶs�DȪ����:���2D�=}�p��V/iV@��IL��FV��Y�[���i��}6[z��	;��Z�_aXr��\5�
={w���Q-�n�Eͺړ�'�en^��7u֡��G�闔o8R��fѪ��G@v��Li�f���y:�:�Z��GhL�(�W��J^f�Rوvc�{so{���bj�����i��с�;���GkB�x-^༵�f�`u�w�*�V�)j\7���z��.;�[ӥ�lq�/��J��:�m��YPiW.�uCbػ2��ʤ�x��܆�i"eUm� �iH��J������i�C����keJ�=t�e���_en���9T�'�`:�9}���M���9wK��f�,8�5)[�vҽ+�Ъ��ܺ�>�}CETD��\�F�m�o��3T�}�t;��Xo���Oev���y�kB=�ns��TX�ԈE}c������-c��Kv&f���T.l��n�&V��Ǵj���h��]@�H����ʾ�޺�2�b+s0b_p�S����`��+��ӵÎ�iQ��dFȽ�]əJ���*��x%T	KŸ�c7�~�q��S���rӴ�0��d}�r�X7�[:#��ܖ�c}2m���h��֟vAN���P[&z�IӳyUZۧ��7��^�vL͛X142�8�˼���m֪h�VDqc{z��o\�uu'{��484�J|m�0��QU�j!��uq��Tk'k畁��$}Oz�sSab�u�{.[Z��8�b���]�20�L�.��Y�R��s��|�v�Q��ک���m�8�QXK�D˒.r�:I��Tj�S5�3)n�YTo���z�X���������N^h�<�`�j�jɻ�������C���Y�1�V����ar���Cf���7Bf�fd�O9a8,:'9>��nga0�����>{��!T�`�2=��a�ժ��n�ޭ0���%=�@��9�ӯ�޼v o�fK�wVj��[J�#;Z�i��0`'��ni͝�s�7V�8�\��E���ͪ4�q�S̄u�բ.{d�Aec]�k����1w;�w3d�R��:�E��b�o�Or[nV`��oE��8.�ӧ>�9�{�7�ʯ�p㫛��W{�m�e���nt�A��V_����srb�\ʇ.r��S�VԵn�{���}U��To/s�*�,�[5kJ�b������9�;2}�TF�f\�$��	�t���x�t��{��wrgo0C=�����L��;��c\��d�N�oՁ�E7E��ZSe��h_h���!;Ss4�2^�Ӱ��j�E�Ek]�Mm�u^=n�iDiW�F�"���!�%�3�f��^�{ڞ^ua�#1U�)�]�j�ж���0O5ܮ�w�v��^���l�ݫ�]��E���YX��;�P��Am,��}�}s���a�q2��v��j]�M�QjJ�o]	MVoxa	��K'�x�SpV�֍�pt:�b�7Q�;���o>��ݚՌ�=��'���p�S�ӵN��1�.õ�E�/]�j����Q�+����.\�;��ĥ��+4�=k6�����{痍�(���]�N�nknaQ��q�o��Vl�[.��f�\7*����Wb�]}�s�� �돪��h���V���η���`�cL���52�M�tw./�H�K]��q+�%���Tˆ�����S��!b\Z������O+��vE�.�lYX��\f��^+U��
�V��i�۔�R�!�ws���d�X��0=Ѻ�Z��T�ʷa��.�V���h�y�Z/yw�SN7��r��S�(���g���U�(�u��l������6[���X��9�b�B~�,AR�+��t�Vu��|i�Vm�Ў��GQ/�]�ptk���Z��S�k�w�TaVl*��|�K�Y+��U��"�YS��l����j�ݗ2�S�8���Q����%�M�
��SUȝ�޴�+3���NbmU���T��V�#���7]Ar�ݜp���n�fe��7]�]L��,���Y�U>��i�uh0��w���no&���nv�9��ݕNC
y��vm�ux�vu�ĆMt��2�nwyI�%e�5��A�.�K�Wc]v$s���k�ʙ85Lꮍ�D��V]�D�*�N��%��}TNRm��[Ǔ*Ԥ��3����K/6�mFbvBڦo��Wl�s�2a]#��3)�n!��;�md�ʪl<�;d����E����t��O�b�^gB(��O`��Wj�O�v��u+�t^Y�u��{��Q��`'p�՚�p�[֗�n��"�2z�-��mc� ���h�uw��$)]�ze�k�}�uJ�Rd"4��BS;��VSlr��^U-B�]�ƚ���'i�|:�{���SCYU�En�_Pި`۾�/��>�;�7v������3+�u3�9v-�{{V.ʂ�	���]��e�7tAѽ��2�rZ�R�|��;�1:�!�_>�μ]�v�nś4��L��G��&���Y����(��1[hf�p���*���ìD�fX��iaj�L�
|�����ɵX2����j��of�_��J���l�y0�N�w��m=�91>��on]������%�ZKrM�SE]��u{k'a��弊VL�~�i����ӝ��vR�&���;��[\���k���ثm�pj\Es������
��J�3�_Y+0�оya0�$����ݪ]��|,ʴ����v�C{3���첎i&ʫn������	C#-�$Vb�K���js+�ԬØ�T����ż�?�uX9��FM�f���"���+��x�FC��-+;W�_,�}[a�����{����6&j�ZOxu�a�*=�刷&�\!w.�P�}cT��\Kj��F�q}k��t��w2�g2�l��^�Z�s���iQ˕2#(n��姘=��[sj�K
^U�j�X{�k�ګ��"����f�,,g�H
.�Ս�^b�V�4��dy��G��5��mP��`��9oCxWғ�q�ݵ��K�뵩��1*���զ�nv^U˾쑋W��;�6v�,���b�r�q�̂΂�	$1B>�4^Z��+�v3qS�&���y�ePv6������y^��XɁ(�ud��HMӛw�,�V�R�ܾ�o��{v���픂�����g���>ǹ���W;U.��^;܇QAڸ�Y��oe�����Ǯ��� ��r�7Ѓ(<�Z:��H���ktuK��[�I�B����qo���_L�]VU�����j�f�]>(=��q���6�b�Y�s|ht����˫�ʅ�X���w؅�On���ͧT�^!��9��Z� ՛�sR#����]�<��w�C��_j�m�h��U�|���c��ܔ;����u���Y�3jƍ˱��͝R�Ɵ&�jX��m�]����?=��{m-�z�&'�T+^�uF�k���\O�^���K݋��׬<�l�h�k�IՋ��7W��f
�7U�7����ͩJȪ��Z��Ʈ����j���o��e5/�c��uU�B}�b�Ѯ�+�E���$V6��ŤYհ.�;���Sҧ��ü�1�z����4�8��;Ϸj�>ɧn�B��d�]\,�5��0��C4�zI������v�<WV�"]}��q;�2�[�S�O9�ۥ[գ]�wV^c����kvQ�̎��<7)�=l�$�yM�yFu.{[�MeM���H�X��ڬ�����G�ǖ��B�Q�'"��&5W�L�����5���R��e������f��u��p�Q�S�nQ��͍�9���"م�21LW���X������|�p�d*�њ3a�cl__�fмN�S�s6����	�w9MUf����|]
;y��ִj����ݴ8]1����(f0n�T����YH�On`/s�E�7�3�Z����B���7G9i
����b����o[�|~� ��D 9��ʭ��H�*���+)E0X��jG��ʱ�.��ʔjvm&B8J�`�:6:�[sG(��6N�i�iJԪ8�
�P%�i�u�2ֳqVꉅ�qX�5H�j�Ғ�B45KIl���䷭
���b��Vi@�<&������f�X�ec��6�^N�M��[Un�/j��Ll�����b��un���1�\M[h��*�v�pZ�MqZ�)�h�k��-f�f�+�
���-�c��J�S-[����
��͸���R��1V���śk1/Pn��U&crb�J��*��f[G3�j�c\����Z��,�ap�gF��aq�:m�e�1���`��h��b!WA�A�#����\2��� 9.hX7X��V̕e{6͕if�T)K����,�f��JZ�Լ��jPcpJ"ۢ���y�,Z孇�`07��f	�<�7�J�nڦ�����W`&���Z�l� ����Z�m.���d���t��J�s�\��͸j�4�����	��G-�&�l����)X�1d�vX�h��$J��BQA�-,�5��%�h��b)�"K��Q����빢D��t]�snn�z�c�`�|�b�����0m<�%��丣��3b����0�Ԗ�ī�B�Y��YYv��f�M��FX�#��kan�R
0�u�Z.R��\jW LJ❺�:���^B�����5���2�����:��R�Y1�tl˲l�$t�ƈ�hs](ʍ3
B���-f�f2)���c%]�p�� U�K�u!sK��&�hl7F�,®���	(�T�]�ɞ���4� M�I[\Xm۫|�L�)d�ue���s�Vl��v���X�4�딲�f@��mf��
ri�#�ch�P��T�LѮ���,��s����Y��X2�]u�vԪ����`�WR�Z0�tʗK��b8�H]��Khm�V`�	cʌ�^��pĐ��-K]�hA�6�܄n��5巪��љ�v�bZ�b�
%@�2�M��p�PVh��@�V�;4�+u֭ �w���!lYE��h�kq�E&e��XMh�-�],55T�m,H��M-0uv6�͂�j�[Vpf�H�&%r���%�M�h����gsٍ�8�LX���FQ�@����a��nl�s�m�Zqv�fܹ#J��]C˷yB��Wf4&�A#4�ESL��6�Ѐ8�Ç]&a4��PfL]6������F���6�e�2.���#ia�e!H�*7m��V�\͵c��F��a)�P�]B8Xk�"fñ���K���["$���!�G5m��Fi�#��nCh�&��T3�1HV��靖iR��ĚSl3-b[�q ��`����:�(֐�2�3�sTH�u`���4YV$
l6�lÌ��r�A!N�Y���l���R#-�ʑ��aW+�bhl���y�5�
�	���\�2��`@!�
@ TB��m��˫p\�J�B�C�����K��HD��.�[Tp0N���6gF��K���rKG�R�h50+��Sm��J\��������a`j=i����M1�d�������p��cB�M)۪��	X֋.�\�Z�M�Ҵ�����������t�$��[ ƴ�\ �TmHͳ%,e.]`�q��bJ�u[�-�3b�/��rU��]���M���/�mO<5����\���i��i�&�r@�`q�c1L����[h�kw]2#Xvq��X/.���G���s��ڷRj�Y�rF�Ń� �t�I@�anΕ�\-n��`$ٖ`ħZ��]e�1a��tu�t��)b�,c�^��˓T��L0�n�Q�!�3����\�3LD2<eq4�v��\��a���0��q��1�ԍ�h���,*�����ţu��0��--aF�%�PDu��nML���0M��h@�	�M1�BWV\����p�-���3e&�И�ڒ����luE �i���tm�Fl4X�bd�m��GT��v���X77;jjJ\F�5�X�<M,lF����[EfT!,4f�)2��.[6�(��c���c���f.Dl��W��2I�'�h�ȧ���D"Ʒ�Mx�0C K��(�J%S'Y�cT�[le#.�
�a0�l�T�.m���qW-J�m�\�1th��9b�yѫT��%��\ʃ-�U�#��A�R�Y���j�#��:�ͩ�h���&X��1�`��v[5��v� �[�6��6qNit�bصe�3[�]�LiC0uf�lћ@�-���uԅ,�z�e4�t����A�=\�J��
c���F��0TŚ°j�^c6�L��4��9!TKt��%+\Қ�G[KL�$�sS^��h�"<�uh&ځ��8%uB�۳l���\(���RSK��	��hk:��JV׶��u�..t�c�#Zv��w6M��e:��Z�i�4/��-!�QV`)c�F�jj�I�X��]/
�˪���-6�փ��UÑ�.Jkr��i3]f�0�+���^�FBk�P[˥���#�yϞM���(d,��1��d,sae�c*����0����	*XF�:�i�iE��5�CZ�cZ�CA�&�\j�r�P)B�F`�]dR;X�-�+=H����n�̋��&��eل���e��,)�Ĩ	�7sr�%l[��[�S
����e��L&�A�J��#�wk14���FC:�ڃ�JmVb�̇$3���:��⅖k3��i0f�kFK�S��!m���8�i��D����c@8q9u+�iE,�:�Gb��<�bP�5�y珞�B\cB��p�s#Vݦ�)4��3���Vf�W[��,�:�W�3��+K eBm�� �A��&M�mæh^x��p�h�[�����\�"-�кL̕&�Ј�$�\���k��J�B�M�k��έ)�4r��R١��,jÑ4,�cp�[-%���Um�F���+��	6k��tQ��itb�:��t�-�!���Ԏ��fj*���x�=�(-��j�,4Yp�\���xg��j�����M�6@���C����Қ�;v�K�����`:l��F�e$�B6.]�մ\�����tNm���L�[����������:[��6X�I�]�fv��i�֐ �h �P$3Q%���h��c1��%A5�In`��Q�Z��3;���tT5�PwjnP�@�AD���S4׮�H̒�����IYkF�i���DҀۆ[f�b��P�#X�eh�B�fh���mͤ|��3h���Z0mЂP�#r�fW4�l�nF�,Z��Ɩ^����lY��k���P����|�B���V�Q�4�מ�f�IX3��f����k��khM7�1�ƽu��Ɔ5t��ї�h��L��hB��kk3Z�@�+t��َ-HSB`,4m�Yt���WD����L�0�憄f4u��L%�LZ8���&@��`�Y��T�o2��bbG��l��d��5hF�Z&�d���tf�=��f۴5D�z-�KfP����&#en��
W	���l3B툩�3Y�RX�p*�ec�$H��-SjXi�����3Z�s]q�E��͗n�D�.�]�Cu�6E�H�B���˭@��lZ#3ipb�-��9�%�`�s��45�1�%�(ݣtV8���u�XT��D� l�4���eu
[q����-X$jj,!T��X�F@�QDf��z�!ر�us	i|g�_%� L!Ktu���l2�jBP��k�"�	�<Ѿy�X�F��Z�hv�^(P�!��r�<<�h�m�E%�tw;4,����6]&,ѣH�n�661br�$�% �qF$�B4l;kA�7���Ɇ��Yf"酮�ۮZ�5ZD� &7WE����6��8\h�ЖU��i�q�.fQՇM�۫xe���!��@�\�w�Fk�u%	-��D�eK��&�����ʱ�q4�F�X0%��4U+c�BXD&����GDl�J))��Sf�#��iEPt%�f�&l��iIe�ڮ]RWV�B�Pj��f��ջC0�X��X`��F��+����\����7:��0��3yk�&����aiv8�z�븥�1���:5)��2�L\ha&�0�3U�� ��Xn�4&�FQ!��[͸���͋a4oz���-i�Y��!e��K�L��Y�1���as,s�3�]�԰���kF�l�6P*�r��Yn���X��wb�SG�[�5h�V�9��	�щ�n�k�]zb�	mt"�0�r���R�[[�۴,ŉ��8��Ц��-ٱ������T�+z�h3Qɰ�-LX�$Rԅ��x���g0ĥ�l�iں]h׆�Ɔ��Z�l3M�ٵ�/(9�\�\�3RZ̩&�k��T�%Ŕ��%����d�Q��mPhۙ�D�,�f�A�,�Hۈ�Utd&�5�m��2WFۥ��:ܕ�HЅ�j�r+.TXS&I3�2��	燞Z_
K+��#��*7���<m�l�cfbf�آ�r�,BT�%�3[��v��5�ι��(ť��5�Ҙ�{5�����a�Wd+v�E0��g.��F2ݹ��p�h�T�ҍ�Bb�e�L b�A%��qձ��ek�e���n.5DLl���v+\e�5��1d3��Vb��Cm-�Rf�6ƕ� �\�ܰ¬�����ح	I��\��@����jeBVi�[��i�&�k��Tb�/8-6MF0��L���b�y����J]�.�b\�nَ�Z�A5Hqm�(��b1*��MI�M�m��n�F\	�.��k�jXa)�blbk֦���CV�Eօph��kGr%e��Ֆ�ָ�L�V���l�b�h�����,Ի�\���- ��q�B[4��Z2ǲ�	teYa��rb�yبӨ��h]5�%�-�b;2�^]ePڲ�4���E͕ڂX&)%��u,� �WZ��l��&����B5�ٍ2uf��uV
�X�3�+W3eX��F<df���1�Ƭ�a� �^����;�(�=���NจY�j�QÜGErP��,�)'%�!(	tٵ�u�E�j��(��JN��(:K�(#:�D�;���m���۩�i�C4�fr$G���C�[X�;��2��B,�'i��	9�a����:�6�G)gd���$�INJw�1DG���.%ڃ�А�8��g9Bbqr9�D��N;-#��P�C�ݥ��u�qf�H��;k(N�$ ��Z�r����P9�h�P�q������BJ���gvN����^��� �NIJ"N� q�mZs�:KkG8�I����C�#��%!NA)D^���A�s��$�r� $!  C��$�/�݇�4j�K��5iy�֡ �m��%�X ����`�aL�ua5&갅D�e��Xm� K���lB&ulK6�؏:���֗CZ��������8�y�c���ͭ�.ېf��[()@.�4����X�Fٗa��Գ"Ժ��\�j�&J\�mM�t4t�f� ��B��&�:��36��	���	���K����m��Ե�
�#��.�R�2���V�Q&�gB[
,)E����0��6@�:���4�]K���wh��AJu ��e��h��]+VV�m�`bYs��!6uh�A�pcZ۲���B
�[씱�����S[e������4[�E��4Ee�SK)f�P��@6�3���,X2�m�9]�ZF]v"�(m��;D-�XLLن�
�\[wUٚb�Y�2��W�`�]�ήPU��G �6��bfR�&�n[FXPevbZ�CC	-�l�\"�t�{�b��T�I�-t5� ]u3+\͌��M�H՗�gD��n�l�x.f̅ ��V�%��؃-�s��ClJR���n����a�����K7���S[�ڶ�̥ɑ4ac�V���1�{CJj�*ɗ�]�b��ei����p��Y�e)q��EU@,!F���lQ��uYh7%j0귎ٗ��bQq�t�mp�\��SE�����l�WL�%l���01Z\֭�ee)�5��LVfT�)��+�)[m�Ұ#	��r�C0�pb]��μ�f-�e��M�����[E�Q|�KHku%��J�j�44�pj�^7" Զ0*a�pP�%�-��d;1�`ZJ�䢕�ٵ�!i��l��<mH1J��b�JB��7u��[�b�&(lU�aX�mm���&KKQ�m��GZ<Xҝ��n��Ү��1c)(�Y�cA3�Dnsr-i�x�jk����Ch�]*��7f�ek�j�=e����W�s�`�i�mgI$�u �[�E
���+m�Ub)�YQ�/XY�Kan����Č:�N`RPK��)V�lb���c���,j�	d��Ճk*J�*���Y QHXR��%mhѢ4����n���YJ�H�ȕ[�BU�Yic"�[mK^T��ea�z�a����	H��qb]I@c��Cm5Rt`F��0p��W)F��^5���@��AA�(�@������\ޢ�&�J������R����W�1_7u��/�M
�Z�Js�X�ܤA#fS���Nc{َ���E
��� ̖m��jhnm�9@?(�~+ܾ{������ac�T��$�}�������K��D4F���/�$i�wm�����ݴ%���P=<������ts}^��V��/���S���7���]�Mn��M��h�����#>����F�G���PdY�O׭n�9�촩�o4W� O�QfOِ19��/���0��{����J&�Į���p;nٱx��CP�,��ҷ#�9��	��_�w��hw�����r���x-��ou�]x�v��y�L�C#� �m A��4F�ِ������a**#<-��8�~����j�ՖQ-p��+w�w�1�p���о�#��vͻ&�8�W���)��"����'�}���k{��H�+52���k�A�������hq�Ai��?�a����OmK�����������A�IK��o��� �(���v���e`�Ӕ�ٵ��黬1�/��w������M׈ |C����*mڼ�~����#wX`����_�^��U�k�bu��jrt��ϫv���/��+50;�����t'�A^���i��&+��ٔ
�b�Z��0	s[�v�S.���[�44�C�}��	���ݤA#M�}�;�yV��IS�����(W?L��[t�(�r�v����N�~K�*��Vv�b"�,{��@��܊��n��b����O�A����̋�db܃��������O�E��%�}z���ǽ���'�X�Ǭ,=w���9"�ڜ_^hw���&��!+i]�˦�=���w�����{v��+�J:Y��<�l+�}�ӓ���n���j�O�x���~���a��H�A��ɺ�!�H"qУ��A�o۹���c2b�I�m��7�"�d�d��֑Gٓ�	<���*��� �`�Г��^��ĺ�CU�<ע���V6��:?8�_M�3$L~"2���n�J"sJ�HGh�V���]�#u��3���l�ڋT�thآ����тo�A ��?�H��y]�����.��W���F���F�r�S�;<���H�H�dC@��j�n����ƃ����-���ݏ9��Y�C���9�A�	�(�&���������3�U�͉��F?J�2F0�Dr�+��,i�{�;�o{���}��Ƅs�ѧ3/QƓ3,z��է&ХV���E��#y]�NҚ��$�y?f�����z����m�/-'	;��:�F�b��D�SA�u9t����d�숩����vvpvMY�2�ҳX׬q4����;ّfV%�{���+�60�2E�C�I`��y�a��W�B5뗛����G!��;������"��&"H��**�[;���݌�i~���i��h0�v�6ـZ!m�`꒴lhvɑw.��]%���%�|�� ���P?(>!%B�_����e�m`8�HV���4�ݍ��2	�A�����d!�I0A� ,��������+y0A��k��vlW��Q��_o�Vj��F�����yy��܉�	~�$a�$LH�ɡ�O�~���f�6������d
�%?)���C��e�d�(�D������A;W��E[ab�x�.\��5����p�����?s�� �fflЌ�&FH�~N�ې�;m�W{��"���G{�}���j`@�g�_W�I�[G�Y��X�������:�{Bna�����Qf�f�j�Lt���#��P�����1�u����+Gb����鲡��߳�~��(GXfz�b\Q�.�)6�`�:�L;c���m(��5M:k�G1���9�F�cm�fbZ�fZl�*���X;:��[�J�R�m��XR�Jb����)*�(�V��Y�I]*�7 �7 �f4h��tf��4�vtݫj%������bL�Y��Px�q6Ф�R�tfшPy�AV��Ե��8�"Ց��ƛe��_�gϺ��,�+5�c�2�AbMIUb.m�e��@-�e�X����$Rc9����_vy�$Z$C_E�{ujػ2���89��Ӄd��O�dY�}902F�Ud����y�*�؝�n�D|@��W�m^潫��Ŗ��E�߈`�͟�S�z�(V�g��F��'������2F8��F ��`���=�W�dmOȍo&�oF?C�}$a�"dl����x��-�Vl��)��kV�ٔN��i�M��@�k��!Y�I������P�L�2��~�Fg*�s��g��C/r�7��m�Me��?ih��A�$O�	�:f*�b��u#��]\X	R3de�t�n��Te�6*7kɐ-�K��5�&���s�vr�q�H��I|��l얦{�ھ�;0g���uv�M�gܳL�32͹�z��7�~*~�|����W�Ê���]Z�w�u^����1�T��6���g79�p��=�6�ʬ�n�-�f��&�C���Yx4�l� �C0!=�ksb��XKX�4�� ��%��SQ���1<�?u@�}�L$_	b��!Uq��x����t��ݫt"���03|�H��!�$�0��Z[��Z�a�&D���gd�3�m����嚾��3K���s_p�~��"tI�~"$I���g^z�#� ��,Ksb��XKX�4�h6�~�6/���+}}�R_����f�'`��$��&\0b[�XK�ai���0�\��y���/y?�Έ3����"M��f�^�lcw��E��$Iro^\MX������L����6	� ���+m��*��c���j�vKw<4��ھ��n��������^����>��f~��#�������"����T�=q�f�
�ߥ���şqz�bN�[���J�wR9��\Z��j��2���F�U�>ۂ��'�s�UW�ȹ3�����v`,%�ps��glЋ�fe�34j3(*}����aezd�{٩�{����	#,y���z屍�-Ћs��� �^N͜�����c~7�?� ���#`�$A�	�P2E^���{��0Ƶw���n紅[;W�+u09��%�_#��w�^RwN��:����&�j�2P
�j*QT�\�9��!�k]6l�jU��~_�@m��)�1	�ַ���zoP��|�r����\�Jۭ���!q�Js�DL�ѡ�T#���N��7hĴ�ƃ��>6�[����W-�o�n�c�0� �j�IH6��bJ�Y���G�6;� �?E|d��$�eYv�j���G��%��m[;W��
���[T(����S�jq�Ý��v��?O�N��h��������i���@�kdQ�q�f~���Kil8�
�T;�#u@���]��i�4�ك-Ec:,ۢl�]-�Ra���e��<qt���;�fM�Nu�T\�ˢ<]�>��?J�~2D� Ig�]��2��ׅ��yH_]�c�z�%�[�[�_r���"�hә��F&4p��w.o��mP9X�D(���I/ie����n4q��ARQ��]�8���������|���x��"d#T�N����%�����/[�3Rq{���3�U|D���2	����|�=R�"]�=�i�D��1�����l(C��M��	�� �d��N�|��j�A_����+��&D�|%��D<��V���~���M�O�[��B1��� F�B�Jh���/
	�,���j�� � [5��)c�����ww��-��:�24�_���j��ε�v+�=`� CD$I��i����`�hW�����w�>Pa�d&�WֶE��%?x$�z.h^~�̃=J�*T��L��e:���,Z�V;w�,���h��;R��R��y<��2w����ߝ��:������L�}����W�Hк�����fP׳]�b�P"��w&�څ��1H=�'<�35v*���t;�6�RĻ3n�uH��s\֦T�f�F�`S U��7m.�F�P�me6����P��-��P�K��Ƴ	j;.Ĭ/li���8lḛ�bV�l�S��ݞ��͘GZ)�bf�{[c.�����Y�$W-u���\��FR�J�@��������<�&��m�LS=E�MtiW`�`ͱ���qi����^��Kx�h�H���|~IP���oʛ��b���Y��]�Ն`#�������~�[�$A��і�y�U^�{�8�Lgy�����%��}\��_O
���|$�uK�o�Z�퉐Ah�"�H�A���G=6�����.�WP�v����6�E	dG���� ��~�(]vu���\��K��'�g�B�)*���Z�[��uv�F9�	`^YZ<)̷��bc��O�	?I��� �E�{���1��v���T�l���Dr��}=@���`d�0~�_#��ç����a%�h�H2�u��cn�S;��D�F�9 m�3
T�.Ck�6g���0��c��%8A!S����l�0�2{��j���">t<uHdQ�畂$�����2"�1��X�/[W�zǕ(%*��Ʃ��{ڢ���L\.5ES���Ac�^݊K�Ue�K�����{��E�Yg>��FB�=ܫ8.eӥqCA�D|o]
�O��J��չ��Ai��3|�H�Ѓ�,��X��0����0O��a�H�����������=O0<�����n��ܤ�_O (�����0���BH������.���xj~�F��=z�*+B�COE�"�����ȵ�&f�V&A�O0��U�2�F?C�|8�z��޵#@n�6�����[�9���!�o�`����S��ޯ����Q<��WWB��K�2�]u��ˬ/a�W�e]YL�h��������w<�`@� �sWrN�i��ܤ�_O
����ܪ�ʢ��>�0�ҫ�"�H��������鶺c���Qw���U5Z2��=�A��Q���)��j����?m}@�}�Ld��.>?$����-�׍=���-L]ձ��ͺt���7�B`�A�ځSӐ�B�l[�g*�:�iІ��:p�|o��I[��7�(���Cկ���)�7��Y��Un���H�Sܣ[���4���+�;��w@՜�-�2�Z`��R,���\�e텕�m�����>���x�tn;�)eի�再�X9P]w�)_^�v�.Muǅv���i�/o�P�A�]Ɓ:0���X�N�m�w�w[��1ƥfn�5r�Y��X�_7�vu���`A7S��z���g�rUB�&���P���b�bA�
�m��ڬ����70w �r�2���:�Z�s�3`����4ow�3��J\Y[B�-�W�AWB��A�hu�UۛC����u�5�ۆ>�/���ѻ�9c8��_M��nc�uӢ���
e��]��+xfB����[��b�h�X�5�z,y��F�̞��[f]���5�IJZ7���UE"���Wb�m^�T��S�}Z*����
T�RLuݽ�R�ۙ�����/���s*���>{�fJ���	�32�:��d��Vv���*�����'z�m��.����"�;��/��4Gge�x��U��@��z�mI���G<.J��e6�8qc ���Cf�|�坪�V�%V�VR7��5a��6KA�W��+�V*�䶫�z�a���ۢE�ʌ0�V��ȊI̛{��WFO|l��Zj0�xxne�k�f�S�C2<�yW:)��L)�l��:�rRk���^e������v+bI�R������r��:�l���O���I����mg��{e'����l��nԼ��g`�":q6�{n�$��n���ړ���(�fwul{ל/[FY��I*8"m�E���ˈ�qf��''q;�'S�'NqrRzڎ�R��j:$�;7:���q.B(.)::,�I�:!Ӂ8�!��9�Ӥ2ٸ�,�$Ok"�N�8!��q!	���G̎s���C�M��IQ8NI�	q�R	JC�%	u��˱٥�i#l8�S��l4�ēN��2�͝kn��E��ӂbI�M%-㖡;�?/�$��4���YQ�����%$������P9�Y�����L��@�JH,9�Xl�����0������}f���$�.$��gyp�62RAB��9�6G�����v��Ux��Rk�G���0�����_v�M��
��#������^�_��<�X�H+�@���n��zᴂ�H�,�AH)yP)�) ���sP�Aa���r�$��������3�C%FR�@�ױs霚��s�|	�7������T��H;(�$������ Ss�3pd����r�G�����fY�)~K�]��Ě\Se�N�V��me�WG`Ky�LK��&��Е��#�պ�<�W�������nd�) �Q���i���
�]��>|s��}��o=�x�N��o��l�y�7��3ٯ�_�$����RAa^�5�����H)�#)yP)Ĥ�Ü�ݤ�@s��Ir�RAto5�t��������@���@�w�3c%$)w�m ��{�;�ٽko�/3��ZA^Py���!L5�nd�2�
��H,��W�e5�{��z����s��Ü�ᤂ���g,�l@���)}P)RAaG9�Ci��R9�4�`�$JKʁH����G/W���e_׫��u��:RAa�v���
B�����I �uہI ��9p�?2RAB��9f�
AH+��- ������?|kG5�[�����M����S�f��ƒ
��Yt@H��m���|	��|���<rҗt�~���4�R<2R��R'�G������^j��<.�s<�B�d���E^ԛ˔54g	�7VU��c�436���;�Y��s�u4�<�U����ӽ��z���K;�C�Y��|���z�$���O�H��Xs��۴������H;��^0) ��Ss�1���fr�Ϋ�s���}�����ZL��� �FF������@`nAa��|=߽M��ۧ���F�38���	k�*�:�˝�i��m�k��!�W�
���N$P�O����gu��)��I�) �S)��/������_^���Xs���v�R����_}|��c�=�Y���D) �0) ��ü��I ��C��H) �C�ZAH,9�\4�R
o?s�~��{y�ﰯt� �:4�^�,� ��{��a������9\�f��~����l�y�
Az��,II�w��6�XlaH�,�Nr�Y����sOi��O�bRAa���i �6@}�٤��R�TH)hÜ��L�%$(C���~���D��j6�{��^�{i9|�3Ф��I ��ܸi�̤���9f�m$�
H)�C���i��9�Y�؁I������u��OW��d�l
B�RAa^��Ci��
@�z�$��R� _u�{�}{�ߏƾ���) ��;p�AHzU�yf�RAw���i��s�I8�L;��i����P���m ��
H/�RZÜ��L�I��捤ƒ���~�z�ߪ��R�낈���Mn��2�Y��w}��'vE'�$Td��
H)����R9�4�pB�%��� ��l�k�2`����S~ˉ�o�tYGq���U�:���b:̱�L;X�!���\�fuN��'jɣU��U���3�Vh�d�_/� }���[D����&f�V.З2��f�5骭ke����/+�ƺ�+�L�X�[0Z�ص�2��\	�Fm� �9��A&����]����0-F��;V;F�l\�a���e�G4��E��%T�K�t)h�2�J]�J�Z�g �*˚.%�:�v��롲�5�9xQ-�j֗�0�1�9�:�$kv�����Yv���{���t �Ŭ�, &�]J����ZF��"�����Y�ljkV��?$����AH(��4�vQ
H-ہI. Ss�3c%$*!�rͤ={��w��7����3��B�
��H);�������?o�g������p�'FRA@���Ѵ����A_T
H)��.H.��9�Y�� RAH+ʁHZJH,;�_�����y�Rw,�M�I��KʁH�����ޮ�~5���I�9ۆ�
C�@}�Y���D) �j$� Ss�3W~�s���:�d�AB���Y���R
�RAH,9��i��) �W9�H) �*�tAH��n~#�JF����{�����Ym���|����(�٤��I �j!bJH,(�=�m ��
@�9f�
Ad��^T
@���Ü���AHv�U��oq����o�{;f�҈RAh�\
H)h��v�ld���!�rͤ���������\��z�W�ai%Sgnd�e$��s<j��,���i��i �T
H)�C���i��9�Y��@��ʌ����R��5��)��I��e׶���E��I��)~��|׻�y��N�~+�߹�s���J�>�,�Aܢ�Z�ہI-�s��i�d���s��i��_w��J�K�{J7�&A�PMQ��e��0.��L�� ��ڜ�m4�8�Q3v��E��g�gKoӂ�
O!L;�놙7I��ƒ
�]� ��9p�>�ev�}����ӻ��@�"���;��c��f��9%/�HpII�}�چ������M�RAH+ʁH��Xs�����U�r�$�B�
��W}��ϞV���,�.�ujno���$����?f�$�O;�6��K:�v����v!���"�v�b��^�ܙ�)�WJ9b��'q��;��a�g;�	 K��$�����L���
!���H,7����;��������fs�B�
�RAI�
a���L�I��Ѵ����A^T{Ms����~�����~*���l
@�z�&�
H,�d��@�-%$�5�aH�,�M�I �* WNﺕO�}����O����߹�s���P{�i ��Z+��
X�L9�\4ͲRA@�9f������������[�_�x���p�'��H(̳I�������R�s��k������3���k�����l�z RAe2R��RAH,?�M?W>��n�����AH(�Y���Y<�^T
@���Xs��۴��P9�Y���R��p) ��.c��{��s��) x7�#�|	�xt�׭�*���e���- �(<0����)���0���`Wǻ������!tY!�_M�,j&�4�f����.L�Y������9HQֵ�I1�֠ �F� ���0d��A�.��q~~5k(�~�$��_mݘ�i�!�p���~�?���H��~���O]xB�Ԙ@��#��"�]�������ׄ7?h37�(��غI! �7��A�`��Q�/��F36�ss;Љւ��⯻���&�!5�p�
=�P�(�=v�����h����B������wk6�=�/DҒi�����	���^-�]�4�y.�ؾ{#�(
�H����.�����[s@HF>r�u����M���d$�P ��gٵty�^#�Yɂ�y�ҫ�"��$a���k�����/vb��qNۙ��� �����)��Cܛg����F�b���*�t�j��[s1���i�zU��*��M����ٛ���g�>h`���<E"��#�w�ݓٔ/�;+�Dה��ڊd�9_�:0��U���&@��"n�7�W�C��I�	�r��4�X��Y���� �~<E"N�Vy�{�`?z�}�ɀA�0��W��F��֯h;����FSX�3��:A#O��РRSD���%����������e�0�~��"H���Xo齕���l_xJ_?q�E'����'�'W��`�ie�ܛY�����$b5��xWщn�bV3�,��r��]/Y�i�@?o���Tfw�4�e�h33C2D�����H�<�f�e��}~,<%︉;�����+�$L$A�ިt�ˡCi��E�JE�D&~i6�0lŶmT�[�u�LQ�(��V���;e��yg���ɠA�
?(��%B�Ӽc^��SX���^ ������t�E|C���lLH��D� �꠲���bO����L�=��*O�w�Z�x_M쯡lLvF�B��ye���
M�}�������2	�yKǓ���Gw�O���'/���FH� �`�

x���;���̈3�W��	*��y���*��q���$i�q�����=B�6�� ��I0�2D�+�$E�꭛C_�\������{��.j�7�{+�G�[��0��U|@�1�����W������V�����Uo䧕�ki���4�ⷄK7:7���i��q�y> ��\rm`}��������Ҋ������n���$���zX��(�]6�:WF�,�Q	�˥9��I�9�fha#�.�d6�l�.Ĺ�����x�/�Ƶ�:�i),0�[J���#M�f���Kvp���[�D��T䩆 ��[�j`�-uv.Z�m��Tk�Iu�4�$2$JlFZD��V͌a�f��j�m�hL�r�Nd[)��2�eB�X��,�˦�����Ϯ*Ь[p#.��CG4F;3u��R�v�Xƹs�V!�������,���0̑|Ȇ��9�f��{�"N�b�T-vb~�(�D� �g�B�2D�[�I{��]}�����_�����5�6e5��,�H`��РRS�kGA�X,�����A�	�PH�Hƌ_m><��e�w��Ec/�u�Џ�&A��]|@�0̑0D1��}t�f� ���
:������U�j�E��d$����B�t�eZ�[���#��ʅs�D��5�];����ce��w�Ļ����{�b)֢<�4i��Њc�s����Q�'���j)2b�2�kq��cCE�iLQ�9�J Qb��0�Ͳ�9���� ���}Ic�u��xu�2�_]}=_R�%�]ݫwu������(W�"�H�H��ɫ��ðj�NT�F�E��v���"D��#je�ћFZ
�]}H�oo/3���ԔF޵�_`�{Ƴ��1��Xj��ѷ�oe�M.�pY�������O A��1����|j��Y��NF������">]W��]�`������;ɐD��~�+����0=�6��{	��щ�d�k%��[��:Aǵ�Jp���lܠ�ڮʖ�п�'O�yYD�Կ<oC�J�5���lr��
u��93�7��^�_o��2D�$CDIfH��#cHF�e������+�:���`���d�Q�/��o��P��$j�`�X�&���)���5�[���%cTn�Ь!bL�����L���3��+�"���z=�)��V���
��Lr��s�`�D4F�2D�����;�����;10A�a�>w��z��3:_]}���:�`���?N�u�+_z�����ɐAh�"� �!�Uʨ��"�^�Ԧj��Ϋ<�0A��vK�z@ֺ���\��TЄe�a�ɴ-5�ņ�N�/�{��2�Nk�C]�Ԯ������7oۓ���X3c6�NGݑ@��d@))�R�P=�,d����0�6��_gb�l�	*n[ǥ��d��2�-ΐA~��������R�k��)��_$a�$@3�d��T���w���k9�=���/���A���%�_#���V�����D�) Ji��e�
iR�\#5��:l��m�:R���Dt�~�ψh�$��D5˧z.��X
��Ρ����^j���W� �{�`��0���+�@�"��k7�_��xX?l}��B�筽/EDb&R�� �0AIТ���7�?-ʡ�Q�F8�'w�20�2D�I�n�ˍ��o'�,��z��\5v|�;���N��l�0~�_#"���͘�����Ή�	�峽;�nj����$�i��`�;�z�}�VL�y�t��H�Y�Y��7;������٠l�9�W�`gn�7�D2,��8�1�|`쭽������J���|_�2�� ��=��5��P���H��#��Յer����[�:����訌Ca Z���0AiТ��hg��/_+D�h0��Ӣ*�B�3�l�:�n��F�3Q�%�1T�f6hM���{��{<�g��ED��ϝ���m����'s����^��7'6X!fȠޡ_$�0d��	�"��>�q��j>S����!�9l�N�+o<��w� 缀`�d�=`�q-a�ц�B�9"D��ҫ�"�f�B��7��訌Ca Z�?GNa�"dh$lS�^>!f$s�C ?a�O+ �cϝ���m���|�b���V���}nօ�{5���z�};�?��& �h$_I��u맺�!�j����+oX7��$�9�@0x�2D�"H��URU���5�Tl�ͫ��\/��T�Y{4��P�^oQ�aަ#����Fy�a��Q����S�	�]!]�&2�.�����WBl�����8(�R�"�y7�r������屪��͑_Y�Y$+흇k8�UJdɏF�R���pŏ���.��C+D�)_l�rooM�|ꊕ)�����rR5�ee�}��z��1�
��@��������At��j��k�>��T�2z������F�`�{4��w}wךcz-[+��-]�m�$��4��#;���h���w�='H��v��gu+�3o��ùa_N�_XU���gV��XN����x��l����fF+�r� �����|89��e��N�a㚝�8��[OY�ن�q\1��9�UK˫I|��Ӣc���ѧ��+�̳s�������D0bz/�jc�r��h#U�^�^(�����|#�(�e���h���J����ṧ�cj�0��Do2Q�������[&����zOWi�m"R;��.��9Tw�{X�,V�
��9���quWL��.��c;��G�Σ�'A��z��i�7��9OT��������{����耻�󡢄�X�4�[\*u�b��
�wo���fph�+UίeLZ��[�Ʈ��ߋ*�^�ڳǲ��ӽ���RH�^N�T�wgZ�o�#2Z�X;I.��<�h��3N
˺	+��3��dK'j�K���_�1Ƀ�O_���!��2���y���pO#0o#h������i���Y�5�8�RN%��f��+s��I6�$,���I�66�`� ����X�Q6��'	�n�6���%��2��Ⳮͷ$�A�A�|�m��$K�fm��y���C�r�!�NaFv�Hkl��;�٢��"QE'-�چ�K,�6[7k��r���N�汶���4wg:9)�l�R[`�98�,���#2��	�;r9m}�	�{h����m�I��"�=�yart��h��p�fnS�86ЛW��h1��$�$��m�����_<��I�ΐVݭ�ηN=�b�	�� f�����}�b�j1U�鳶Ŗ��%�U,1P����
X2ئHZ���`R��6b��M�fvB�I��a(+�Z.ٻ=[����2Ð��+/���>XŤ3�������R���"˘���˛H�DM�6���R�(���$1
M0ˣ-�j���2F�!��+�ڭn����`�"ǖ�a$�Z6bңx�l�Y�2�8isxu��`��۩(��C��
ĺ:�0V�Q�X[�V1֝�V��(lA�#ұ���e��h�m
U��5�7a�-��e�"m��T�H��mH8:�gk�TM�RTf�5�0�	�YG���;I�IQ���+�3i���ʞ6+��k)����(@RVm0\J�:�fQ�0���9ltT����P1�su�!G�MAU��E�p��	��!,q�U�r�s,� ��\���ˠZ&�c��u mk���.R���Ć2^]iIsnr�Vެc�E��e�)Ak�c��/f亸�f,
��m���iA�)�d�s�I�kx[��c��
Z[��)�A�CU�.,�ћ:;kHub	A�։���4�l��%�Z�b)5���`Mt��1�3-�n��,�ːY��D��m��6�����Q�S�Sk6C<7V��a5H�\K�c0#T��M.#*hBb�P&�%4fUθL�s�m��-lmWk���\a*஫iF=o84-�\�[RJ��靪�hJ�RˈE
S'(fԹ�de�
L3 ����H�q���\��iw\�:զ�at$�b⎉r�,4�u�қy�!uX�6 n��]��nM%.YS2�B�3f����e��j\;�h�BY�&ڗ3El�ƺ�TUH΍)�Keh�M2Cm��ˋ[�K��e5e��ٵ��)-uG�4Ќ`�Qʱ�5Hcv���l�XZ�*��d�Ż��3�	6��m�R��ld�y�||�v,.�ŨK�h�Y�`��eR�m�V;[��ĴI�A�lՔ9���in�"�]��q�Ds���t	�m6��$���y��n36�]��kP2g�����6p鴱ba�Q JE��(�H:Э��)���s��d�K�r��x8,sMc�n���I������#��7Sי�x[6���$�i--�L��V`m8bD�X���q��f�y͙j-]�cQu;2؀�ytHvg��tU��9�5jB�٭��+��ct�΁1QR�1pA��N:��m3'���/�ZdG+β� ��P��SXKve)!�F!Qd�ac����y���}�4��W���	*!筽/A�Acll�x�g;�\����<�2y0A"I�dKT,�k�·��-#��r��x_y_=�|�b���V�������w�q�aWr��}C�ff�@�?I�E��`�b��m�[�z�zN�m�k��$�0A����P2D�H����C����v�B��0��#䔊��������Hs�g�Z�>�V�ϏtL�D5�F&H� �E$J�j��ӌ�B��l?K����k���;���lL� �҅}$_Lיy��,�6�I�MQ4�H:PJ$M����fVh蝶�SJ�نc��\h٥�OO����}��_�H�!����zw�6�%�L�w�`���L]�f��u�G7� ���2D�#t{�ʜ�>��F�#�ݓr��51R��mQ��T'�Ur�pmz�7����
���b^���4��Ļ8e�Ƭg<م1�O��vn�즱p���j�����ﾪ���|D�@�W�㬚�e6� ]΂#L�a�d�̘������#7܃{�0A0�2D�I���O�9�uD��}˷{r���m��_w�
ؙl��,W��#����2����X�?z���{8�M�z���L�J�Ȅ���A�5����W+����a�~�(�/��h?K�2���<a�R^E�t��e4� ]ΐ4�S�E%4�Ko��)7���T-��B���"�0��˂�A���jݛ���ǭ��fa�<�oq����|���(��H��w=2��k�ӎv/�nM�u��l��� ������|d��"� �h����U���M{D3f��0S���eUX��J�Ȅ��7�A���H���V�^c���@;9?�"H�?J���O�MG��ދ��yRxU	9�=�l�U�������UT�yF����>v��(�:�T��8fr���}���#n֢�;��8}��ߢ"u��sF�̽!�A$�?�|1-k�pT�^�B� �t�=�L�����n{n��k�Է;�G�+"do�Vj�yg� �����v��F��w_۵t���y`�F�o�{۩��I��)�w�`�����Y�#G��}}��>'���5|��Kc�V�,�l�`M�0�fM!b�9�˘B�3����X<��!���(��G�%B�sֵÃ������=x�Hn.��,��̡_�~���I7���h�n��`���L�=���]����Z�Z����VE��`�,c�X�����]l3۩�@�D#�n��V�\�=�٩���ro#5Κ��l�gR�3.h��fT�F�|�)vs�)`�w��Ma���H��ӗk\8;a�� ]O�F�#}�w���j��m��}v:��}�T��l�S��VB�����;���yʦ�n�J�v�R�/lV��t�^UN=�~�Y�W��]}U��o� @�oz��߄<�L�ѡs"�	�P2Dm���֛_��A�n1+�̖}�K�S�_w�VD� ���~�>���Hĥ��*��f����	�SK��K���s�J(8��X�SL�Ж�R�R��m���� �["�))�@E�7�OoSw�8��AN��w�FV<w�X?x�$L$A��
� ��b>�F�M3�W>a���|V�
٬��c`�y��΂�/��0�2E�x����N��C4G\l: �&FH��!K������B�D{���K�z�G�;��@��2�#�W�I`�������P�@�W�P;�hHF>8��~�Iފqɼ����w���F��W_Ua-2�a��}@�"D���F��e��'��b��+j�̯-݇��0����<~��,� ��˦�1�p��G4z��9�h�Y�=x��ٙ]�^��+����~���*.���ʛ�w��e�2���i[��w��R"%�*dK�k�EC߀���7qR��S�4؅���̫fu��*a3rrĘ-bvN�1l��Al���ե�J;f�աi�c�u��4��L�t�V���]�FYFa��\���X�c���)-#�J+*^lCqٓM[c3hК��[m�R�k*-mT��[�5	��(5-�dݝAeԉ�.��n���]ՠ���407��p���J�&J �Wk\k�FRm3|���E?º�P��,a����JMH�&Y��Ńc`�(��T����顏?r�"�)���&fh�Ws��vW��qLS�}�z����d4�'�P�F��I"�C�c�T�ɽ�sB6���v~���1^��,rw�gy ψ�d�3\��B���	`P ���2F�W��0��铽{�a�����[�pj<�j�B\΂	`�nE����F	*�1��EU���=���������ܝ�+Μr<S�}ޠJ�L��#zN�wT1g-�43�Q�3F����E1��fh�̽�<ĂOB��^���jӗ�^�S�M�w��=� �@"d#��W��!��W���M�����t-��Jt\ìu`ڛ�5��*a�d�#�ֿ;�{rOMH���%!��ݒ�G�mYhK��7ɪ���J�����0�|�"I`�.]b��ߵ�:�x��*��zu�bp��&D�jc�yZA��wM���u�����*��Ъ��j�[�o�gU
�����i��ֵ�,����|>4~k'�� ��s��4�*�N��+u2�da���(Bqf�������<h�����& �xk^�k������W�%憹ɼ�������_"d$a��Bg�se�,]������	*�Yi���Q�VZ�tH�~���-�)^�zj�H��"H���d��z����޿`�wl����˒��;��V�`����U|D��<�Ň�oFL�Am�L�*N��bT":
Z�Ԛ�t��D�,%{V��qu4r�-��A?W�0�2D� �!���{b�x�5�M�w����/]�!`��9�����f��e�2��.�No(<�������t+�5���a5e��/|@���a�$D��w����x�#���	��20�2E�?���^��'����kOwNa�f�m/431���x�9R�/r��+��{��1��~z��۟{qm\R�h:��O����-�6���/b��O���M�� ���!�đ��0Gy���>Bx6�?/r;��D5Y��lY�方ɼ����9� �!��i�������_	b�2D�;#�0Z�Y���cc��:꫽��:*<��p�u3�0zs��T��e����
T����:)�F��i��	SQ"[X�]��,������7�6��=� ��H���F{�2Ob��mb�k��]�=�]��?j>ƾ�������F2E�"3�Z��J����*�,�ܘ �
��{f>�.i|�ވ)�`�g ��H���'lo���*�= �$�3����(E;v�[퐷3֓��G�X��~�@��2D� $�0�w^��k؂v� A6Eo��Ib�י'��T��X�Z��_,����os�#8Ol5���&n�Oj_!����%������y��S�]w-�ϓ���pw*��j�U�ڦ{��'(5b9�ї�7�H s5z�3=�Oٗ�1����(���!��Z����,��Ǐ6��2���7�
w��܃ �@�"H�x�l�GY��T��T����/R��6�T��٣�kZS!L�v���^���x���`�(W�I��fw��	���.K�;/[�俼��w��e��}�A�!���0&H�-�ŕfh��
�LG��1^켓�W�fm�)־�P%f�d	�ޔ�=/6���g2&$q��0̑2"�*�(_��2��_\�.���7y;���0�"�2DȒ �Ҁ�(X�많jΉ�A����
��#.{7�����W@���A��0��V�3�u��ȸ������$��d�0A��($W���~`̷r{)z�f�b�k��~+5?�;#�W�D�K�/t~�u��2xF;F�1��:ֱg/O�|�i�f��֌�����2n��z�bD�&U[�}�+ii�/4c�nM�%�S������$�����s5��n��t�HY��#��X:&Yn�ƌ�%B��,�+T\UQ�%1tX�&�+RcΕĔ��3lsy�.M/`bG�JJ����`�.�M�)��a4.]C#��AM�i��Y4��u5�������.��B�F*&j�Э���1(�m�T�F�2S�ex7m�Y�EA`�P�)sl{W]I�P�k4�B}���S�G,t��Ԗ�Ke�D������褩��M+#)]�0QBi���������2D�$CB�}�l���.W6�� �y���:o�w:�Ϸև� ����_XF�Ud��E�ò].����X,�菎�С;X���S��BN�H�[B�))�z���Sp�b\��(���`�{b�E$L$C�g&v��~�����Rꙛu�����(Vj`����RF�/���n��U�Y��l0g�0ACC5���W�O_rmM�Aox0~9܃^Ŋ�b]gf�3��nY�E�@%%?RJ�
�^�ĕ��Zt!�e��N��� _�@ �4�zy��/�>r���N�'��z0M%�:�ٞ.��0�qrƣl�]�Wh%xX۠��챮r4E'�������"��0AF?W����Wy����"�7��w3s�w4A��?x�$B�2D� �\�6�7����6ʅ,��#&�P-s.^�yyi�C;�vPSdɫ+(i_g^����ޝ�+�v熷W���w��V�b=<FfJ��)׿��}���]����޽YA~p�f9�~����� �Z[�r����ta��"�;�|đ���RF3���C�L��g���er�y��D�B3��L̿�bcI��4S��c3j�ʑ��Oڜ����_F�W��Wꙻg;��ޯ�j`�;ץ�S���(
����H�`�~�$a�d�m�^ձ�[�(�;�ב��51Ȝr<rr��(��b�^xq�)�.�M�a�SE�!k�L5-(R�Ym2f.2�@c�k����E�:w��|�پCO҅|d�UgL{��<�PZ@���d:�ˡ��P(��g����F�2D��Ý�њD�w�2��/_L�u��g9u����A͌3���V���������#�D��d��A"���OI���q�����M侵T�UY�&�a�[5Ns�uShâ����w3y'�9����<�x�	tR+0^�1e�1`���-�ߟU���%K�R�C���ŭ�8�ڸa�W�]�7X��dڅk���`L�GS���ꪣ�.�]�P�t��p�[Uv+�����,,�ҸͩU��d^]�|2�T{GR��>�&5(r�I���V��\�7_K�<�k�cF���G:s�YI=ʲƫ�]��N]����.��{�����X�.��Y����@�&�^�A��kC�lP���v����Jh䮬g��(.�1t������WѠ�S�ӷ.���g�8G�*�2��N̸]l��)�u���y���������Oo/3M��%�
�*��3K1�oFF�_8�nZ��JGr�L�`@ڏ���Ln�D�e;]�Qc0��'?��[��$s�p�b
��
�d5w��G^r�0�[�uy�{�񥽪�U��p�NUNYTj�ux+��lKW�:�K+���8�YG+yU�t�o&��ئsB%:�1�+oK�۬;y{*�um����W�1uU��j}C^�������z���t��%�ic��pgU�`��AMo
�od��􋬯�op���3'ηiC!�n��+eq/{餷w���A䦞�sؤ��98�	)�-`�M�ލ�|w��t��օ��#���cud��U�h���<�d��z��H(���FwTktl��8����o��ɖF�ڬ�mb���QY���]�F��Nx��4�'(��3��įqq;�nU5���}y�?iԡY��b��E�T�I[c�v��I&�GY�օ�L��NI��ߝ��f�I҂H�,V�df�8s�BS�q�i�qN!I�4�c�DI���V��H+-�</ka݈�rj�2K)�� [vu����h��h��f,��{^��gν{vtU��ؕ��m�m��-��6��ֱ�!i����G1�m�x�;f�)Æ֛;Ag2�re��l��`�m�d��7Z-�d��mm���knp�\�i������	��5��nv�	��mi��7aٵ�
}�u�h��&Ev�Nm9��gv�aMm��,�D����
2�mqe���[��(P�Ս4�K^�I������#t8w.,�"q��	��
:D���H�?J�X��|��v[�������P��R*n��ݍS�$Kh9�@#L����V�����c����%�A� ��FH���qб�j^L�z�x�ݳ����P ���#6 �?C�I�B��N����D�l:D�Ѥ�jT+��#��k�j�M��u��,\��]4X�]=��0!㯒S��yOo^C��ܖ*n�{��c:ɨw�^�G�C�'H�}<�#�
�H��q����j%����>ԤW�u��j�>I [@���A#Lw6����0\lۤ"M<��r�E"`�"���`�:/�4����3v�r���/5|�c�_#�"�[��t8� �j�mMHF>����z;�+�"�� �D#��t�f����R�'	Я�t3A��qV����=ӟ6�eSj@���T�b�ӽ����A+~�u�;6�ܭ;W|��ݵ�mP�>��}�<�ܽ3��3�̽D��4�Q����ǳ�+ۺ�v�Z�����Tw"[@������B�JhHE�L���������|-�V�)�kŚ�]u����.�;.�B��\f2�7���`y���
Jh��J�};�5�=��0z�;��K���b��љ���$I��CDӛ���GD�G�w�f�`��^V����;���ȋz+��"��E$]UІ����g�?wr���~�#�U��q�3#kV�L��2b%�w:'Z������"���١���~�,>��bO�����H��޼�:�T��y��z����B�+w]��:쯫��w0��&A"#Ħ�sSZ(A�ǖ���1�[��GC��nf����: �FH�D6�<Z׻�,\U�{��u'o�8��^����s��F�b4goG���1�#'Ǐ5�!��c!��xWuJ�{�������I! {��QM�bqR�C2�GX�)L u�Y��A6QTsc�������a)+���:eKH�F���u�LĒ���+�T��X�n�jgJ�9�g4&�%��g-r4�m�����)�S\��X�b�1�D�č�]�v#i5Tu��SK.1Yff,D�	�1(�ܰM�B����a��D%�	t�th�H�E���8�"V����Tp[�4~�|�_����v�:�s�CU��a+��5t�[�q��4P�B��l����N���"{�Ѩ3*Ts3F��Y�ln�����m��"�����kl�3��ލ�r�Li33SC̳H�3|یw�~��xC;_1��\�{}�?)7E�W`�^j���������ݍ�q�t(�~�RT(�2"�R�8��f�̛�C�����o!Y�`���2��P2D��#�����]�Yy�?�"�Xg�U�0�Z�����%Nb%�9�	���{Aw�o��($q��0�H�fFH����i���{��
�goqW^ٺw,��|�S�c�K�F�#w���,��>���JV
�6(K��ip�+F�h�l���Ƙ���F�����Yd��%���f�RS_HF�-Y���Bhz<����r9Q�p�i�O��''�H�?J����B��ܳ��ly���f����,�f(�b�[\H��1rݮ�fQ���q:k�!*���oNY��o��c�
nl�۷j�h�����������_�B.s�tkQ��1������I�Z��g.�2��88����� ���("d$b/n�@��]m{')��⏶f;�ޠAY��sc�G�$����X�y���5b��� �3���s��ȏ�{6�������\��7..�D��jd��Ҋ��zL�ѡ��+}�=w]�K�f���*s-�)΂�3 ��͡EH� ��{,D|9���T����R,�H릙���e��awe�҂�!n�K1�R:�����m�_~:D��$�Ax�֊;��9ܰ�|rf_�R��fj���0~ꯈ�?��A�~y�.���� �h�m��3[��m9�К�{�m��5�E|d�o.��U�Em��*��&"H������빗����3c/������*ĤW��E���o�A���Ǝ��3��K)\4��ǯe�;;���Zr}Us��  ��m���2T�()�R����a�"~"��-�;��"Ȅ�E��D4:���q�ٚ]�,z�f�Gl��<�b��?P�����|A�H�H��ͮ�?c�f�^͙�W�gAuw�(�	�d���ED��6�̾�.�S��J��Y���F�gB��ڭ�J�K0a��505RĦ�at��^�7�9z���e��V�ݾ�t�ُb3�����_m�Z�n�?,~a��O�4F&H��������˵aM�����#3�3K��B<Vj����~����Qi;;�\�;�0Aq�����&@����泵[���̏/o���Bhz=�j���j � �|E"d#�*����_+���7��"�?l}$�P�����F1\��t�� �8���&V>y3|*���|w��\d̕:����YT��6\���о��8U�����N�3p��wm	Z�T��]��{�yP��}}��x}�ni:��ަfY�Eħ3.�N^�u����"�B~X�{j�כ�?OP%f�A��W��#ñp^{k�.O{]V!����%F��РJ�͘a���+3m.��.*�t]a����}~o�8�J����0d��A��N������.��P�S��g)���H� ��J|AF�B�2E��d*��p~���p3����v�	��ǧu>JUJh'S�8�_v��d��uYɊ�V�5ϯ��W�E����d�z�D��ݼF_eͧ}����5|6E���)"+�+Z���H��%���ۗ��&���mzr�q��{���y�v�	(	"�H��Q�g҆�(m
�9���$W"QN�������)-���������;��X���=tf����kd]�3�^��gQ�w�/�X'r�휽޽�v����5b�Qdb�N��齝�u|M����w}����#KbXg��	Uj�u($��C
S.-v�;Fip�h�u�$��72:�J��K���k-L:=��13%.C1LP�����b<��j6�`R�V��0��	m9Ylz����X����^�t�w.�S`��L�uu�6�Z�I���Dkj�&�� T��B2lJ��d!o]jG��\3!�ك1�s�"Жki����ƒ��%���R3{�o���_�l9�-�5�ۡ��p��6�(�k�]�A"�E-Ů��j�{�t����RD$����F߲�Ӿ�f{��7��w�{/����!$BIUt<�dg���̐��5o�ϡ6=^�h<ߚjzIbkX&C��a�r�@{ܾ�H�����m��F=�랫kɼ�w��InD��ӟ��ʞ�H�T�m�{�\�1uJ&1���b���F{o��y����Y5���z���۴N�`P�I$�e��a�jq=�ױ�M�W��7��[��I�j�՟yW���_�#��e4j���&zض0��P��u�;љ�L*K��f�3���{�����yb8����J�zU&ӭ�:{���ָxqT�g-�%�$_M��|��ܑ�<�~5B���c�m��}���_S�}��7�l������s��ֱ,^�X�:��w%>8k��*��[����_@����}q�{.@�r')e�s��a��x��Y�v/��K������5{�$�l�	7h`����Wy��7S�+���=	�jK�|�����*)rt�[�\��|����oN�µ�p��)�}�!�68���ә%+��$_I�$��z�"y�4��^5��p���:�v3<E�݈I_I>]\e�T~
�'�뮷�`%\������#hŌP	��Yl؎���0�%A��~�W��I0	+ۏ��s�/%�>�[c�wLN<2�Э�x<��RR��CT߯|Aݭ��bٹO����˗2�������o��¼����2�n�����_	ܾ���}$����z��mSW1r�U��O)J8��[���mI\v�NP�.
�����c��b#s\�5d��a>�d������6]����o��<F/^`��b3��"�6)(	"�O�1�owƼpZ�����J>����p�{y�unt��N_p�U�q���q��R��J�x�T
qu��8�kN���p�nSߩ@6RR�X������ CѸ4s0�k2�:�4ŁkhJ]5q5P���T�h@M�E5E�
O����7�	"�*Z����^�����coݞ��XmzS��/��{�>�)"P������&�nl�{rw/Y��lץy��4�|�B2�ɓ��3Q��k��yI�P�d��)vnf��R�;��r��Jl����|��~��*\X� �K�%?D�,�dE�݌�;�|�!��d���z	2�1�Y6��Ǜ6)�3+���UƳwWt�w#ݳ�x;��T�h�ᵤn�Zo�μj�6��h��;w~�� ���q�Z���P�JIDLugB�U{f�����Y��cs�Ҽ�w�|���R�W~�Ǐ��u�g����L�%s`
\4̥�f�c��a̭F���3bD��|�&�����~(�$��/[ӱ�Z�p�nS�B���<���|��%���$LZ�}D�s�R-���oC1W�c"[�9�VH�R�֮:Ab�Ҫ��f��@I�!���9<�dԚ��]�c��*|�y�,r>�T�	"Rh�S��>�W�oyOP�/�z^w��ں>ʒw)�r�*���O�Ц��_9�	*I$�%I2+^�� ��� {-I���Ŭ���]���j���%�$��1�o�d�V�W����k�x�H�v]>����6t���V�EL���3sg^�_iՎ�e���f�
L�U����sh�vC��]^w<[0h����34��qh�fɫ���0��;,{^i��<j�<�Ԗ��$^���>�b�����T[��d�bHvV:���}`��R�\~�C�Gz\x��f,XO$e̍�K��#�O��M���r���(ww�]SF��F���{����;�0��2�uE����]�}y��ע��l[�c{+���̥��*����I.�s�c��:�,I�su����`�x��s��tw�3�O�UQ6s2U⥲���u�b�:n�+��:��@T��rj7��V�Ӓ��1�J|y�y�|�]�U�;pK�[V;3tU?��l�CL{"4et�3o��t&���nB��7���{��51*Ԇ_g3b��(��]�ʪw���b�ԌWh���N�5j�O�on�v«*�u[�駊��+�f+3+���wt�g���U�7Ju�F8hز�c��n���"ж��r��w�@�N�t��o��/eh��8s�h�q�NlV%M���4�����=gfz���k�W7N,���GY-�R��;�y�~��� 9�Bʣ�1.����f��䠉[1�w��ynH8E&��ƼW��n�Y}]�x������;j�z����M��[��d��U�˫����;׳��:��5���>����yZn���iesv�XٮY�Un�Ʋ�#�����	��ا�KiǷ����v���U��2�]dݽ�[���Wو�Q�<(E@��@Q�N[��f�m��a�y�h�n��e'dRV��Z�ش��M���vg�$�++)�[-kb0���m�Ճ�&�gGm��g[h;"2�+"��m ��,��H�gYͭ�۱nm���vy�m��,�m�۵�̎�ݐ�twe��m��`������k9':-;+Hӓ���;s�L9�g	�Z�f�m[ikE�ii�YB9�%gd�#�+v�iX�vp��$sZ���<��m�y�t�������Y�v��a8Lf�9)mݗ9��w�u��l4��3im�8��m�yݧ{ko���i�VZQť�͑�-05�I�gm����jf�30Ks�f��kVv�n�:�(K��n9��gR�������a�h�P`�f�mij�Uc�ە�KZ3+��Cj5��J�	m70%vƛJ��i嬲�
)e��k�����9]	z�ScK�����6��.�����9�)����Ѳ�#t�#x�m�����nX���Ĭ��2˜�Ż1��]JW&��n�Py�/F�[k��]favR!jq���%c���c1�Z4��LًcNu��h��]\$���մ`�"°!s�p�M�gvv���8��h��l�.�`(F;B�MkK¢���Ci�1iKP#gu�	�I�hWH;n�s�.�ikj���F8��[1kt�%��k�T�Rj�Ql��K6n���T#u�J�,�Q�bCX�e�Sfjm�Y��3U�m-�,�4�;F]�کub��L⒅u�	�g0���G.�z��x"�C�)�:Ǫ^4�Y{��iP]%���r��jk��n����x�L��h�٣�Y�l�jk���"�a�6���-ȓ*hF�n]�]��G4�a3Z[A�bH�u�6�ɓ �.G�vYfb��mv1�0ּV��tc
LLB��2��q�+/�5�5�]��!��h���MH#�ML����Ra��e�a��8sMƸ��K�Kri	����2%KE�)x�u�k,ל�2���͙-M��3�W;huI6΋CY��Z�Q�b�l��X[1R�e��,kf1�f�1�qA!5j���"�Z����55j+4*SL�Lr��pZ��n&��FR��jRj��6�`*����5��Y��%H6-�:�]WVa���6 �q��l �5a
9%���itl�Jb��l�u�)ƻ�e�e.BA�lL��n5�`�ڥM��J]*(FmN
�K�a,���&am�"F0l.��Y�Z3�UQm� J6훱��ie�R�����[]�nb��
��c@�6��55��[ !_2�S��LX8�]e��G��C�\�\e��1^MIms)�X����,1��r��ۖ�kf��9��O1FWE��c��L��ń�FT&2Fň��/[�M�F�n�\�n+�F9 �P�`c�&թJR��d�mˉ�Ub�a2�YQһE�A!�����X���Y�V�`&-#.h�˥.���S2�	lk5tI�MC�sl�2��c�7�y毀&M�J�u�.��YX�ũs�WZB����U3p-�bP�-��GF�aZ�c��_�?m	`�/;X��f5�v�f ��5����bm�2e�mc���?���?}�ωO�@k+ۋF�X��9�6h�����{bW��k~�%)@X�v�͕��\�z_��)���;�����j��JyIS'�<���/��PE�X��-�&��}���z��.��,��b�J�I$�:�)���ӭX��l�J�w�ţQ�)�/�[߯�<3��̀����I$�$��"��E��u|y�37����9�C�K��J>T�R�_p�[�/9��UIpj�t��(X��Lc��5:l][���H�
��3-���oP����/���\�{�k<��)��۫~4(��e�%}$RE%
;�H:�SԖ��;W)M�w�Ы-Pð�]�_ak���tm�f�kyh��wQ�7�^�>��^�U�ˋ8���� {�@�W�ţQ��	�a��K�	#	҅�RЛC$_I�W�I��w��dz���6�Bqicr�Ӆ�BQ	(	"�_F֞'��ދ�"U�g{�k<��)��SU��Mgw��f��)�%}$BIu]~*����'��ʫ�7��*h'P�Z+���J(��u;�U[�/��أT~o�-4M%���s�lS�֨]�&��0ܜ���}��}gχD���׺6���Ҷ�2퓲[�z���$�"�!,�����ײ��<��3���}������5���LWk��/�����zIbH���kU���H���W]EI(���U���2��<U��f����n1؉6�\K����SGj��L�2E�w-���%���Vh�Q�>�׷��*2���N��}�c���IN%)D���M돪W���$�����>�9�ג�t]�R�W���}o�CeI"�J�P��ש�{����yn-�;��,��lRW�M�R��[Y��<�_y�g�tM&sX�h#S�hdk�M�c*V]�SJ%�=\�?>��q��JBQ�O���Q������r<��a�4���7��	+龜5��s�,�|���mz�AzJN��&��?P��i��}�*R����;�}%	"�I6��Vv���Jי��GۋZ���Y"���/��;�x�:en��Bڟ�ܗKV�C��s'������	R=�c���=;���fm��q���b^Aً7�U/�m�=���]~[���'����mY����g�޽����+������|���$vL�URl�2�k�cQN�^X�=����IO�,�|�f�̃�+U��SN���m<Tu��JX�-43�f\�Sf˰3m����y���=��%�$AIw��3�Y�.�w�0�����r>�'P�!�!&ǆGS�}��Ŷ1C�~���T2���䰝���>I^l1�I�ܭy"����<RIx�:[u����>���X�E?4���{��>{��%	"؆+Ļ����� $�*��Y�5E�)n�h�,b#7�83�}@M��H����!$���<��w��u�׉�*CȦ�a=�9`���	]Vס;���rS���걌��-a�V9k��ts1�=�s3�T�Z���]�ݶH�)U�����ñk`�1Z�c�-e����WV���og/��T�>��UMYR����(P�Xô�&�
�j��Z�J�.��B#f�-�eҴ�q*��)��΅٘��,�6����X3t�p�w(冶���A�(�fe�#\�V���"�.Z��jɥZ��LM�%c	m9� K��Rk3���tcFGm
(ډe]A���[Sl�M�D�]S;&����KkrK�@�	P����ڗ9R;$�{�'�������ֱ�B܅z�v&�0l��n�ȝ4S4Je���L���|��%I�^z����,jX�1�{��j����}$_q��{�C��~�y�Y�3ֆ�	��p���s;�sd�&+�w���e��9���IXK@�j�2F�;�ڽI\�(bZ��8	$������N#dӻ�]�7�$��z����j�4�@ؑO%�u��ً���|$��%	%�b�@i�m��f����{H^������
�"T�٫7��������f5��H�Lh,�&��`li�6fd�f�D#M�4���)y��{yI	C��=Os�燱Cd���5g����_u��RI/�"���7�·w.j�wȭ��ͨa�釆����&�g�m;�a��g��=̓\��t�b�v
�YU���$���*�;�%I�n�v�<�|.|��9����=��y�V4����@I�*T�2
�&/��}%"��H�g�h�~���u�k�5\�T�;�!�/��$�H�YY��α�$�3��<~���<�xe��,'�[�c�⧼Ӯ����d�X� $�O�g8Ղ����ֽm=���mF4��{w�S%�-�/z�Wֈ68���ߐl6HE:��&�Ap��pR�5`kT�o1�v�é�54>}��ߦ}�%������"�ܹT��9��Ckad���#ZK�)$�ډ�ZՌ�kM�ڣq��V�y�	�XOBW!mI&]ث���3�4X뗶&�I,}$�95�O$�f�e���܊���f�s���5����7W��^�gV.��A������Ħ@FP�/qa9��}>����t��ډm{��BI$��zv1��.��Q�ݟ�R����|X�Z�]�@����r�H��X�/���j 2��t��w��ޛ��ߒ�a%)-����i�b�LقO<Im)�����[-������kFm\\��Xh�d�O�#�}r>���(�%!s~�E��^Wk�]�~�;]��[��|�-�@IBE $��Ȭ =3�įv�m;[��Fȵ��g<�W�l�H���;��Ʈ�>rq�IJJR����9���n���R�y�����`�I��zW!l�����~��f�ڥ���hg��%?6�ާv;����v߾�Y���=涻b�~��;�R�-�&[躳2�ۺS��č[��׳Mۣ�m�omը�k1ǂ�7Qu�r��t���z�~�]��p��$_IBIM�K��[�G卯�j�6i�����]���H����+ufM���ȓ����%�,��A2T#�tv.7.%E�38e��P�PݲPI��?z{�O~���ԉGەM���y��c���;p|��Z�_d��ܤ�XE[�X<���-�ۻ���*�ƌ7Y�(�<r�8���}��������$�$�iuU:��^j��a���q�3~W��KI��Y�ݺ��腵��Ml�)'�/v�~G�c���IO�7���l���C���$_	"�J]מ{���d�:ӻk`�*򼶉r�G��9�%?%�R[��q�#(�M"��ZC��t<;�.A��̼�d'��z�pjJ�&u�}t�E�ۏm5jkѝdA[]��{�nˌ�u��5����$ɯ�4�n�\ˢ[,�Tڑz�F@�îB�.�&����k`��Ծ>M��9��]H���\b��,*�#�X��c��7K��Fdt��n˷SA%.�.�7�8aay[t.��̓)Z����VۙBijF�;.9TIVV�X��n����yf�J�WZ�1Ukr���Ym�aP���PH�#k1z:�3ڑf��j[z���#4YG�uՔc�~��~FPk�5h�U�Τ&-�B:m�M����,���-S�{�?f���IO�����j3jʕM���>��V������	"H��������S�7����8����v���X�a����|�;��:�����럒R��[�w&�z|c۵ov�+�4K��+���lBJ�H�K����3|�y^�@I>}��zV��>\/��z���⣁\�T���o)"�J�H���yn�l	sZ/��#ూ�zb��K�Hدm�Ձ3����I��i2St�&@�R�34�%�Y�.�f�Գd��;U����?~n������ާT�*�a�[�W��[�b������X�/��Vйa^�y�����-N�ǭ�9��0�ko����z`ɒp�U]ᣙ_mk�r�0��W��7�[���SbEM�s���k�Fu���v�;]��߂�NX� �P͊E�Bz�v.Zv���fv�ϧP�)� �~��S��������bo�-�RRI{�R���{F±�]g��]�|�H�߯S��W�<P������e�|�f�(I�E����a����.^H6�3���׳Q��~[�脔�@���u�{}�M��B�H�p]H[��e���[��!U#)�l\�if��R�;��脑}%r�����{W������??N���pŸ�I+	@IH��O��u��������͟�oש��+ҚP����j~IF;Y�u�/Tz��y}%I�O�'K�1y~�kP4����^��;L�ܑ嘂B멾�wv�o,����nd��W$�W\�>ď�fl���v+^2̰R��*T���Rw*o_�33fQבb7q��8�kӻXe���l�Z�f��j(���)�#�#l)o2��νeiTS�����M��qW�*JB������H�U�ӫU�����s�أ� /er?ep�mb�۩�L���<�:�g-�Ȫ�[��/&��
ۼy��
��ï���|J��Ҹ�׹ۑ��(E�]�sfs�M�����}�.l�nT�N��܉7�`y�I��y��]�U*��&��L�.b��WAշ�S��3�Q��W�7:��Y�Y������y��*�7�hgъ'��,��{h�9���T:�M�w�1N��I�{t�ؐ�Y!��N�vVed�q�}�CQ�CR;\8��=�'j���d����)�.��6ٺ(M�O�
ƺ�N��V�9+U��}��jaT�m�
� l�q��̅���)u
�vyP����/�X��>�YO���:��å������0�24�f+���yB+Y��w���ǽ,|�;��Jk�`��)�ѫ�x+�s���tp2��7��a�v�`7�7�i��`ỐRf.�(�SrZ���C�xx��V�zy�"Y���ܺ�<���$�������C�X
�7��wS���R�z����*	����%�m�ΤVN�t7���1����Y}���}��R�'5�[������V��^q0�=OUf�|w�����L޿f�Z��~i�U4R�
�;f+mͺ1�țrDo�����.mklNͷe&ݡ�;���V&۶ݶC�2-ȸ�[����y��q��"��z�[d&��䈤��,���m�t�I�ZڎH8Mn�Y�vD$rv�l�[�6�"NfH��wd�
+0��,4 ����ބv����eEp	�[8B�Kn,�t���[k9f�;n��rF[[��Ym�v[�&�/������i�R(m͔�Գf�޽ IIJ�͵��ۜ����D �j	Έ�*m��8�ֹ8�@��$�p%��e����{O,a[�ӱ�2��%�I��|��ݘ�}����N�:N�9��mӻmY�Z)1��m��-�}�xAiٵ�m3Y��hQIvm��+-q�⓳�� '&ݐ��e���tVn�ͷ��ߏ�ϻg���f�������W�H��&<뛽���������N�\==�5���[fſ
JBA�f��!қ��y���JRI/�u~܍�%�kۇF��J|d�|�v�D$��Y_:�ƕT��Ac�eˬ��]��u���$˪��%�0�3F��]��}���/��'�6z̕��|�_�^od�5����T�I���"jIe�U��r�ջ�8rǅ�-�HNI������$���״3|��!%	%��}w�θ��/e�7'=)��v�G޷��)�(	)�C�h���_��=�_�I�}���d�L)˅�|�W^������`�N���G�V�lD�>��P��f�v`0aWʺ�j����0o$�?r��t#:���6`W�}�ӏo��n@IHJ>	E��X~o?�]��g{�kN౓��Z%)��)%�"W�X83!�N�|����_&��c�cYp�08�����3�ڷQ�4���`E�@��_!^���O��+�$@g���N�Ty7�ǚ$�2����ے�X~��{P���$����nmz�gg�9_���)Fm������Ԅ�{r_*e+�߻�}6!$@H}�w	�ts�U����]NdX�ᅚ>��p���_IA_�^��2�,��K�{�$B�wy��ܩ�n1�4z�K&"c�,�d��>��>�BlBH��HM�l������/\���%o��Q���u}����P���z(�4�]��)������yTk�
�k�S�ͭ���m�&���f[�6�l{X��ȫ���mK�ݜ�6,���~��L�MD�K�KeR,��iR��Z-�m{i�4�+�E4v҅��ńŅYacme�ڕeZ�&�����C@m`M;a3jCa�)�,[)V 0̵f�t��e�a0	Dk�m��]��Kz�]�K��6�.V��6��c:��Z�.������T�\j�\��D1��v �(�6b��)R�7Z�ꚤ#e-pAn&���:��/�������D��).�0Ҧ��P��S,�˴�J�V�9�����e�TQ`��e���$�^��V��s"ǅ�Z
��3�Q�Q�㐒��$���7q��<ˀ���~����T�7�ǚ>���))������A���jF�)BJG�)n�~l����w�d��5[p~u}����E$I�kٓ1W�wo�W8�~J!�=+wׯr���xd[�7۸;���˱{��I@I�)
����z�����;���T���^<�����J�HY!�U�G�~�0��V��1�u�#�����hiq5%T�F��k�_S�
�%*�@�n��_oW�E���7�=�J�a�����^��k�ڞ£��/�>|����}$_	���)
Q�[w��4��D�G]ٜ��m8Zw�N;�j�gXZ6���0T���v�;(^+^�vs�Y�9���o���@zw%�[�쬱Ga^�Y c����7��<x��֬I%!(	-������*�Y���x��[~�Zy�� 6�W�I'�ɻ��9�3b�d$�7Wy��*n���?�j3j�{���$�$�$�I-���X���k���{{���g�7z��$lw�Y<�O�|�����V(��T4�v�l-nƎ�u�����5Ah�ɠ�F��~��M�y|�/�܄�$VӼ�~��^�'�E�{�\V��V���n�'k�؄���I�Zqxz��nn/�{�7�=%C��U"���C:I���V+�~��	q	���	"���y�fxv��3�i�o������͆ҭ���X`�U���Cו��n��V�x�^�%��jD�R�JRM���IU
S�#�f<�X�zun�=�#��lL�.jޡ$_	"��P�s�ؙ�d ��N���"�{�?Z-;��hM̧�^�-����}�BH�� $�F�f/v��ͦ�w���p��{��VtBJ�O�|e�/���租��Ġ���б�Κ:���j֠�sP"�!����A$蔱���脒~	��kݼ�X�#���B�
����$����S܀�!%}����daq���y�׾V�\ǧW����i���6�$�I�"�q>���X���JD>�3�m��*Ind��W=�g��Tzt�3��JE$D�đ�|B��%� �y|;bJnn�׻y�
�ǖ�,�j��}{Y��V_��v��k9�Y}��P��������X�̲�ř�R�ڰ�2̪E��gu��N�C�ٙ#|�y�]��?w׽?g4��O�%!++�f�Dwh>����j�S��wy;߽q�q����>쩥�F���T��>�i�ET�˘M6�0�f�Tt��4������7,	+-���� ���3'��ֵ{9fC�ЍR��<�ڨ9�y��������l�r�u�)�������^Z9Gao՘�έ�I���c;Pݠ;h�ݰ7V,�^�3�^Ub󼖝���C3Pݭ��=7̫�	�|�έ���Sm��k,�r��~�[�����9��z����|7ww�Iaٞi�����׽鹳F���O�����|7v�qkj}k���Ov2z�ikB�v��[��J�sn7ٚMv嬳P�LSow���lq�j����9��S}�������X��W�����׿�ejb��j�J�%�b�ɭ�K+���Fq4u���+[8�@�ƮlgS�-3�2[��y��sC#�M�[���+�f����ƺ�&�.r�[&��+El�sr�lέe�B�B8X�L˥k�a*�&�ԃH����EPGV�f�*�k� 8���2U��3/Yjm5�"�c��G�����˯8f%�,QY���L[vYj��������g�Rx�&ݙI�Յ��Ra�:��+{�J=n�5�Z2�W�# � k�<3 zz�n˩�ܬT��Ӹ���n������[��fFfHo�2������_��C�]�����z*���պ;��8��:����_n���7B��nȪ��VnO{2�������O��un���7h	�[�����}�m�מ��\�g���WN��(D��}�w݊��gPݡ�[��T)��]���­u��Om\�>��H�����zT�Ii`*_2�ݠ��.��w.)�6�n4k�W\jLG*�u�a����f�g�dX��'�^+�Q���L9�!�����q��9�d}����d��=&ۘb�󣻏M�����{ʮ�wv����N�x�[zr���'޸.��o/�2F�!}F���g,!�n���/�ݮ��N�-�u1����4��z���}��A;�T����-�� fGٙ��-Ka�jٳ�>�zK�;E{����V���� ��?exmk4��{?f@s]�N�\ٚn�w	��UQ�fk�3��^`l�/5�Cv�un��J�`�c�;^J6\���O!�z ���fd�7Ws���ł�(�m&e�*����`�j���Vnb�	\:��.H�*bW{����� ������*�El?�v#E��8=�m><�۬f��^���rr�/[���o۲��b�}~��~��}�:����z�X���u|7u��t��=+E{ԍ����De׹AY��0��o��~fчA�pۦ���ϔ��Yrخ�am����*�2�5em����sR�HuG�"�U��T�QNw���wW�v�hR�,dY��8	�&�����V�֢��
e;��;~^Q��{_wP�����[��yujM���~��/_�+Gс��{.~��30o=7}~�v���U�¹QCM3�+x�݃A�˨���J�id���t���N�����7hn�ʤ�츈���^r����v�"�\]{+���g�n�7u~��>��˧�7���[֢���Zv#~�G��Nd�/NN�b�E��?��d̑�e�7�qW����z��J��Z��Z>�������d}����C]lu�_�pJ��q�ב�yuUz�_)˽yEM�t߮�qna ���R�{+�͸�5DZ�)��1Gs����wVuuc��k�][Z��7�ۛe�D%��ͤF��j떋Ua�[�]��}[����7hn��Vw�4)2���[���:5�� c�`��hgj�7fh�����9e�T4�EP*��4i�4E4R,�X��Դ
��"�u#��E|Yl�(RmQJ�G�;�n��2�k���~x�F��l`�a��O�߾�hffg�̍�xAm�3�0}�.��RvDj�Iʆ��d}�3M�UךV�_wPW_f��n����3ު4�ZA=|�{�����N�^���gn��������Y��Kp����{��O_�/#���Z �^�Z�wK�f&6}�n��v���7V�3J�doV���Q��VM'*߽��>���fx}|ɇ�c:�mf�ں8�uM;���v��n�*�����{VR	���N�p���ۥ��uu�[�v��|��H�YƉL��OTJM7|4]��{"���
v�\�!�Y�L#��y�_Tцn��ԥg�ŋ��Ӵ�:Z�L��gh԰���|��v+Y9pn�nм���K	��aoX��g2�k5K��'nR�]�=�Λ,��-\8�c�K��N�n땓j��0�=��NXX���)gP�f^V٣����X]��ۣ��ݝv�ꜷ���t�!VZF�!���qgl�3;�hi�-Yv�MY�`سTsu��s&T���V�˃��2;i����[$�g#��3W�sV��m�V2����|ڕlㇹ�����2]3���A��`�N����vY�$�iЦv�`�v��j�E���_L�ڴ7V>z����d�O�PS�[���ܒwU-EY�y�]�:�]��:V�v[vwWK7��JU������U��������u��\܎K�R[�E,���)V�\�mΈ��Rm�rL��nw�鏶%t�82�ʴ�<��uV`�L�c2VX'�F��[�3��G�(��z;w���u]�H��3mp����]��<�]
SI�ԗ,zm�ҩC)`uc.�tV���P���&���UMꗶ���wWY���� ��B~��B�[}�;����v�x��`|��{���6֠����
�S*ښd���<1�:�r1[J�nm��۩d��Ű�����zа���v��t�O����c-�M����[v�Vs�˼�:�k����n|�F����"1��S.��L��g��)GDgv�g(
�IptDs���H�P�s+I.��8�a)"��v�';���5��t"N9�X��s,��vią��$$�'m�
*"���%:)���l�9�3_���!��2�rJt�prG^vN@Ͻ�^a�罂98H�jqJ'$�N��9�Y�nYM��)��R�X�䜱��l�E:p�aR�-�㶬NQ���6�6�;t�3G�����m��e�96Β���zqt�2�9ҳa9!�C�Y�_n�r�;�t����Y8���pge�)%�c��ڱ�2��a'��ͯ��(s���qE��2vr�f�챶�;�we��m�*��W���::��E�AJD�m�3.��H����Skq/��L�ZS�����B�1`�e��.A��{T,6�K�e�Ҷ���
�6	���Ij���aR�3�f��5��fם�M2a��#��q�1Y��b���k���e��k�B]q0a�@����LR����X%L[,+]�<��u��hi]K2��5{Jj��6mɎWPvF�	Ej���s������B�j˲�XM���d�ad����]�³Tb�kn��b�X�Jn�ƃf�łT������tv�@\��#M�j�5��k��jMS]Ƥ�6�uB�e��-����e���7U1�f�B���[�ql��*X�<[5`e4���2��qx͋H��
�,cn�I��#�=c��2�z͛ZKuL��fL0�@��Б�-�f�Z<��T�]F�����,��]a1��4�`�ˈi��-����G�)�i�0ٷJL8�+X�؁l�6莶�芬�U("ۮ�&z��v�{SM�k�����̗��g.�V�#R�ڌb��]� ]a�L����֕k� %j�K�SZ�㛩tk�A�l��+Xj��휮�c��*/) �����-��\"�4���ٵ��,�hp�Y�hlڂ; H6���⚗	
�\��[��m1��K�֖�^;n^Z݋7 �x.�.��-�3���,����,��]U��6@�6��Zn��W%&�v���*��tr�lS#5��/Yv"3fd�od�*(] c_��J�I��\��(Y��f���VV��j2��d46�s[R t�F$kS7i�23bk��%΢%V^��3�Y�W	�Vl*E*��P�5�h�WB��j��u��a��8!#ZU�X銉�]Kv�Y��&�-�2ڂ�����0왍�]k�h�bֆ{6Ì)�#��li��"ga�&�m�D�]����1z���u�V`��b�����$�f�6����/:Đ��f��u#��J�`� &��-�&��B�YE,6�λU�X�A��i���g�Yy�v-�X�<�i6Ҷ�٫�Um��b��lpMCKE�8�@"�6����G��7\��e����X�Hb�][���\4�Ĵ^�"c��kf^me�Be��+����K�m����Q��ػ,z�M��+N0ٵ.Q�jJ�[�΃��\E�lDԹ�ZGe dn��k��[�l�S�������\՚@���e�7��}�Mi��z�yqV��sBa�fYj:]M�@�2h�B�Ql�)�Y�W~��$��@n�����j+b�tKN�h�8B���]K�Ϟ��333�23��"g��}����v��y���>��.Y?W�6D���d<>Ϡx��޴0�_L�@�"�%"	J;6<gvw�����-1��g����wdp6�Il��M�� ��Cɿv����s��#\})*ݹ��TOE,���q��}��>��]��r$N�_$_IC	FH��;�nA�o�]�՜���%��/��� ��"H�|�?I��x�XJ��N?��a�B�Y��ZA!cf�e�-�j``��6��D][�%�F��"H<��J,�R�Ω��1�z�8Z'w�UNN#���@P4��%�L�}�3�C�u~NҌ���{T�;���$�h�ڡ.��(��U�x�J���p,Փ�̏.;MD�:.I���w���y*��X����?/����V����Q=��?q��A>Q?u*J=Y�_P'm}Q�-���$BR$���JD�{���|�6���H����~f���@�_$a�
Q���l�6�_�>Y���H(�^��6b�Rp�ml�6�I��g&w���\Pg�M7�� �������1{<X��6�>N���AK�� �|�H�R+�I�w��)�w��Zao�}��D����P]m����u�ل��ۛ�Q�mҤE&<=y�0OmA�y�P ��K^���K��J������>�������#��"�%"2WϏ���i-�f�E�uD�A8�m��wpو/�S��w���$�'⒙P���
�����^�� ��0A $��2F/�;�ׯ���5Y.+IznV�$r��GL��[u)��s0��W=��뾪d���N�Th�_6\������r��r�;�P�G�<w�%.�"��;�f �� ��_%?�A	*#x�q��Ψ7z�FzD��?RR$5縻|�Sī�K|�'켚8��Ѝr&�e���Ѩ�T��U���4�W9�{�V��X�u�M���"�pE���7�'�A["JJh
R1:��#6f���o������f�J�ܹЎ75R��0�8e-p����]6W7][���}�y��HO���Jg�T)���v��4!0�?q��^6�	��{z>���
)Ă	J$�A�( �<�癢|�LGD/>����%J���_	�MsdI`��B�p}��a�w)|Ae/��/��?%7/\ۇ�}O��Q3�Z�צ�?�E�9�-���&e�2�W�C��;F���!9���*;w׫�&xЄÔ��c� �(��7;�ocg�-���[�ں����ۼ�c�Sp�)��3��䪞Qf�*��M[��O���.�_<;~�㫢7�}�=�V�쩙�~�e�f_�)����F���G��%io[�x��˗��	�d��$�})*�(����䧟�U΃[Qv��12���j��X�� �����%M��)vE������?{����~JM>;�j B���n�}@�{��;�ۛ<��|�H8�hBR^�@))�8_EO���;�G�#�D�~O�=�����B
S��� �(�:�
)A�S�xǜzg"C��<��+�H��%4BP:s�9�*o�k~�{�.ZJ�[������͑?�}"H�2R��|r�el�)�y� ��a��$~(�׼����f�8�lo
�F�.��d���۟��`��	��!(![k��1������*
�����)�^~�q��(�R�`� %N�Ŀ&<�mM_�_r�����4���x/ov�5i���*<4s:��Xދf�_���t��z�z/PQ٭!EQ=Zo/*ԫW��&��h�Te\�˱´F��0�M1�e2�q�hA��]���J���H�!n��4�R��
��K����l+�d�Ү��K�0�)Hk 0��s�Ykf�[h0�G�ڮ��0\,�M(��[2r�,9�Jq�HJ�.� ���<˥��
��
F��Y�s&]�4
�*8�]YIY�MpRU��b`�H�U`���[5�-�٬�U�c���4�˰��{�I��*K]KJj˖P@)�%������ �2����f-�E
M�)~��`�� ��2D�	@�^}���ܼK[���B��Y�����@{־ M�3%"	��#1��Tk�Q���5��F�����1s�|7g�� ��$��j�z��cs�������|A	H��?��|��*��A���r�S.j�Gθ�}�(�w
��H%(�%
pTu��w@�"M� �"C^{����Ŋq��\7�#��\����'y�������2Rd�� �$a�%W�q@\�EcB��w�l�=Q
b��n�P&� �Ȓ���������wF���,�i��V�0��V�#��aV&"փ0�]�"hT}#���'��X!)�JE���d��x&��q��:�E,�,g��Q��O��� �R�!%T	J }}����4�/��u��{�u�|�q%ܼ�Vv�Ź"g�Yu�z�wG':����1�j�4�[м7n�������T�G�����(��2�?5|�!�O�wt\���KR�����@���	z�G�]IKqO�{�0{�	�_ $�0d��+��j.Km�;��uQb]ףvz�6�H ��$��% %�"�H���.����yN�v�I	G�T;w��|2k�x&��iQ���AݲmO�0٣��ί�=)$�0L�D%7�ާ63g��ǵ�l�u�m�D<y�"�S����7z� �Z��$a@V��~�t3s�2�	�;*ª5uA����ٔ�	).�,���c,�M�&�{l`v���o�c,��B�Q'�@���ݎ���7Ȍ|7R}���>V�c��@d��}ɂ�"� ���0��]�����=��6��Khnｸ�NWQ�Mu�c� ��A���+�PF����c�7� �{B�/�I	@��� �"�ϵ��Y��W�s���4V�4|�Ǧ=���2�3C�rijᙦ��m�!����B�(����.wE�p7#@D�2���f�&�M�Ӽ�M��\}T���$��?�|�X!w�.�em?Da=�(��D�g���ڈSp��c�=@�y|Cv?C���������A D� A�M
R$�]�c��/�檅-۶�8et�ѧ\v8�|���qРR���o{׻>��/��i�|�I��jY3��[e��(	��L^#�h��Mu�����篬!�ݘ�ND�������nÜw��ԭ��Y!b��g��H��ޑ?�
����E����F?Fǁ�B�~Y�q=NOW�3Z�W�����yA|A��v��х뫗�[���W9�A	H���⒡���"ӷ�g�׍�3�*䰥�����A��)D�JQ ����R��D�p+�����P5?m��W)�3gG<P�o�23��2f��D_�ѫ��;v/�f�4�V��"�Vf^z�j4�vK��e�ར�~H���T��]<��2.[�y���W?}?}B�Q?~)D�R+�R��3
���7��ԛٞ�
mO)������%�H� �"���e7_~Z�aҦ��t,m����K����I����W1�ML�{���9�Ft ��䔊�����*谥���Ԥݸ��Q�%�G|AǴ+�$�
Q ��
�I8�k����_Ҕ���K^}����%��&���A����7�=����6�c3�ը{�w���"�H���ό���0tJ��)��6�i�;�8�� �� ���)H������c�t�v럺�p#6>��
�w۸��΄��
_�����Nl�<���wm���U�쯶Ld���A|d�=��w+�*�D����ވqt�cn�] �|�~��%�1}�����ݣ0Q4l5w�C'�r�H�f���H�IB��[,4Ѭ�^d��}��v��ٜ�Z�����?m�ק�R�<1��}vKX՘�� 1%��U��SJ�X,!�%Ԩ�b��Ģ�惥��;K�K��������x��6���6-� �d�9�M���5�����ds�-�]��y�7Xbʩp:����
X.��;-e��Mk452���0Q�ZVch�*���ǔ��ѱ+�v�u�wck�
�����65]UT�C:�� ��YkM5�!14�(���>�￳M�Y�b(˚��6�!c��J�Y�Vh�Q�V�N�(:$QI2��e}�_W��J_�����zcD�E�m>�'�q�xr��|'J��7r${�_R�$%2))���7��(X#:g��"�~��Nx_F+�|v8O�I�B�P�%S�\ph9�$R��t	 �"JJh��JF�{�5�RUk{Y�f�4�8� ��L����$�������frhdnf�Qs.�j,�R�ןwI�1k��O���J�A�E:�ψ��O���� �� ����0D�\��+֯�*���痛\7#��	ޝ� �mD�AiW�E�~)G���N��11%8ɂ��ۨhhR���c1��&��jG%��[*2h��YI�E/���7���FH� �_�^����\<j�p9�H�wyUFWz~��4��_IfJ_A���/�iV]�}����ѕ���|ą!����7U�	-]��!ܕ��s�k��N�3u�e\�\D�f��)���n^��af���[[��^��؟�W�wI�&2�}6����͠� ��_I��S��S�U���Oť4A	H�BS��BJ��c�p��c�Ԛt�̕c��N��D�ZT+�H ���кG��\�qr$��@��#W^���]\�j�p9�;S���"�0E���w0���)|A�H�2S��5x���0����#d��]��|6}_,���))��R3U���v���m�@�T�Q�ˠ�ASvX�	�ݭ�Sg,��,
0]t-M�ۙ�Q�Z|���~��P�9J~�IP�緎�vd��O4�qMy�ژ6�!�ܤQ[��H#���I����z�{�����5��}�`L���e�� �o&�c���؝�7$��nB�H?nĐBJ��H ��]+��@�K����8�c�^5�������j�A�z`ꭎ'˪*�����p���a����!�=��˳c�/���L7}WT.�għ��(_mR:�����&�B�rh���5��`1L�n��\��������������)���r��4P�2Bi/��J�<.�8ɵ%+ϯ�US;�9��x��{��T���D��Yw�f]WZ�:}�?3tR~���^w*��e�D+n���8�e12Қ��qc�헎v��v����L�ݱo�٦u���mi��.�S�F�"j�*��2TDC��r̖�?����f��̈́���uǏ0*�|6�W�핔�E[�����I1/J��F��).�a˔;"���u[�,�3�,�ϱ|�=�3��W�)T�}�셵�0����ͦ������X��f�W{����J=��j�ła([����-Bb�z��Η�Iw8��Ya@C��(�0����p{��|{;���/:7]0T�ګӣ7j<�dVT�-ݪrU�w�k�ks������W]Ub���v�g
(�VFkh݋Κ8I-9�LY�|���;;�va�_j�5��7��Z\�W)s,w�IU\螺���_?�����՗i,�����՟ioZ�|AýG�+r�6��X�6�7�m�}հhw5�Gv)�3�t���w\���
�O.���bU�gv^UR
��j��2��MYYR�]���[��ؼk+�d�ϥ��兛3UB�^��8����{@���rin����V�c����Nl�ϵ��U�uUT�Fh-�f���):Jӻ~�޴n������̔"�@���.�ä�h�N��C�n���N.�kh�8�H�̹�N���ס�[�*��j�)0���-����N�!�j#mG$�$���8K�ݔ�QDvs���GZ��qd�m�C���3q/,���Nva
%�b�s�:��%)m��ws�d#n��F�6Ӝ$;l�Div�S�0�B�-���'�qm�mg#�ģ���I@���ÔrB'���N<l��u��KkAD٬C���ٌ'F۸"���<*:3.�6����(I�2��NK5��pRA�Ւ�6��a`vA9e�w[bΎ2΋����"�% �hJ�ڼ�g�r����m������%?%�y��W{����r�$r���
~�:�7��;%��c� ډ�����r7�rQ�y��8#w����+)@��?�O�%'����OdDv���H���5�DI�o��[���m�������%@�m�zk_m�`e�3��*�Ǣ	Y!t{P$��1��.�݀��e��N��&Q�9���_�8���.�B�Q �J#�?op��g:�	�z6
Y�3�{pWH���D�I	H�AIM�Y\w�s�)1Y+�0��?��o��N��0��mq��Q$ҡ@��v��g�*f�3Q$w���K�?%?$��)H����~��Dga͵ٮ�V����] �q��c�?�����QJ>��}����;s!���ݱJQ"{��p��yy�
�|6_P%d	#�69��b�����ˋ�6���>A�
̲t��Xp�YD����s'��u}{y�.����@j�wDC�+,YN�<"%�ǰӊr8p��"J"�"`�$A$�'����Qz�GW%���q�XvkN�~8�H�`)�����&�5���ꥼst�8ԂA���62
��u��mQ�6ck�(���ٓ�������'� �$A}{��&U�f<��#��r�3]���A� F�}$C�� �)��=W������e��G*s����#�YH?�RS�f:n�*C58/� ��Hw�0A�%���1��^�1ʧ�{��n�r��0��mq��'e"ݱ�d�A2RI`�g}Y��=qw�nt	 ������?%"Fo�q=��%[���|%t���sDR�z���{��{'���:�(�%(��*R��6ōΙ���>șm[}�U"��u#��F�	���_%#}��p}N,�׺�}j�ɼdQ�Uֽk�;���)��(𢸵Ӿ��a?+JyͿ/Z2��sǹj��o���Z����u��85s4�e�.mtP�sWB�A�n���H�[Jh�d�cj�K�uQ	iƍ��T���ci�PP�Mn����&4� �u`�Fji�h�k�WT�֨�r�r�6��m�uH�p�M�ѻ8N6]i�+��S�U����%b����ܰҮ��%�1����Af��RB*��[�bh\p��qZ�,0ᖡcf�s٩٠pM��o�׿��uI�8��r��u&���m5���aJeLb�uC?��V~<��0��ف	L�BJ�o�ާ]]U���;;���z����Đ~���폤�$��%�n��ڢ���S��A�=��p"V;�^��W ��5��I	`�����o�����Q���lI���@�A)GP��Y
���Z��ʇ�^O������ ���))�!)�$�?g^^�R"����J$_I{��S���*����� ��>����߳��_3���H�#`��H�1)hRK�np�1/>��x-��U����J�4?c�$%"~IH��Oo�\�������z����Aaj�,ol��,n�̔���!٣�����sM�B�U�����Ѐ�����
(� ������F�ȥ^O���@��
j���E@�Gd	��t� � )ad��E�$�A�>t�VP�����l<�-F{N�s$������H�N���;�U�����%�·��y[m�{��Ғ�.<S{J�7T�a��3�ޑ@?o��=]U���;�Q$<R(��>��r�s��0|����`��D�� ȁ�����^�������*��_H?�h�1�	z~!%B�Q���k��"�˄.���~J'k]�q7�B�ey>W0Om�~�kh�����&��D�IBJJ~��I	7��{��ϼ���(W������R��F�N(�CJ��H&J��[���rf�^U���
uUE���^*��Uam�Y�0���j�\R�d�M��ȿ����l	 ���)�AJD�;�o��	m��|)�˷u
6~��F�=�\��%�}aq���eX"�Tk�Ώ/\���`�b~��ؗZ�{�1�N/NW���w�	yH݁%%3�=�]֬\	=��L�V��o�� ���!(�RT==�;��C�wK[�~��ġ���ca�����@�b�]�^Y6��Sop/U}��k�sc�ǍS�[Jq.l���x`�v=��~���y����i�A���%��*��r�� �Q �ڡE(�AJ$���@��1 �!������͐@JD�֟Ou���|+{������C�S��zn1{<'�n%���0���_)BJ����Q}�x��TO�}���cx�~��'�ʑ��	 ��"@))�(�u�������刢��C�N��Sa�	��ڙ�X�f"솀)-���a�Q�F~�����w2k�9����%"��y�c����x�68�^��.�4�Я����(�T+�In-���#���^�@�~珺��-���z+zA ���?�-��Wڇ}�!���ҾB%B�Q'�7�H8���儘\KW8�w�)�0OmA��FH��� D�!S�7���B7���!܉��s?�P����5��(�g�} ⏪{��TV'�1�o��+i8����.�֓����۽H�j�7(w&oX��"\'s�=F���U��^��N��Ƌ�x�>�\D{ڙ��jfPY�e�%=T��!yr7��f�S����&��[�}7���DI_!$bŢY��宻}o_��cj��cX��e�u@-���1���e@�Z)��ԩںa�~�}��'���x�Q$�H���q&7�j�'��j���X������y�ܨ�+���M�R����%4F�!�t՘zݙ�1H��~y��q�Ǆ6��qQ��U�Q�k����O��u�As�{B�� �� ���EVG��y{urM�����Y6�
���4�~!)�J~J,���9�، ���(؟��D��{�I��Z��R|��KP$��D�s�G��
�L����"$_/���� �"M��8�G��b���Y�P���6��}�Q ��P�R�����q��lz%���w�/,�ϤWL���U�9a��t\���l`���[���o6Mw�M�1*��6�.޼ҷ���Jx�m[J����}K�14��X�L%n��_���O��@"ƣ��w
��SE�mF�L�"�Kcs�HB�t��SE�`�aCJS�����iL�h�k	���#�2�V� �c7�V(*�f�ғ-IeС�a ��ǝ.�h�`T �(�kP�A�-uֶ]M���ca:�H\kb��E��a��a	]v�"��queJ)%�F�f��s ��h���������#�e5�y�qJ!Y9�15�Av�3c���b��Pl0�b���ᗟ�}�"uRS@��c~�O���C~��OEoH+:q��t�X� �@��J��H#�I��iFά�3^џ��~:�D����Lw��z���p�KP$��"AIOU/i[�{9��{4��!�"~"�~�A���X!)��X�Vk�9>��.��>�v��4��>����T+�H �% �0�YV|�d�� ��?�� ����w��t�TC~��O�o �V9�C�����������?ޣNeZ#�V#33F�2��7_�[�Չ��`��%���'���(P'�7h d��dA��T����]�4��XՕ3U�stf�.�^���j�̶��Au^"�Wj��4��	��g�͑ ���	*}N�>�M8-=���)�s^W���}=�@���d�D�����A F�����P�;�~��"�%��e���MXe�|�hݺ���]V��Â�rx�-Xio�C���h�f�^��=�m�Ѷ���}1o�Å�������DR3����w�oԦ��[�+� � ����-�5J�#>/bH �ĀAX�QJ$�R��o�����v_g���-�R��Vp�AJ�_H����H!)=�1�N��q�x��#�D��3��%B�n�o������F��qD�1Pn>`���O����9W�\L���̢�̲㙗�^�L��X�>��cW|��Q	�zm>��w��%|��0�og8�{z����Zz��-�7�m5p���W�pV�Gac�WhTh�gK��Nj�����BA�q	����Q ��H���x��[��O������{�Ε�k��U�� �)��̐2���@����t���0�ٟ�6Ew��o���]9/F��(�AƨW�(����8�/1��1��~2�HƨP?p���%4)��X0v.I�S��aܺ�"�X�u��b���ز=��d���%���&^��eŊJ6�C5��5�q�ϰ�Y��;�LX��d��}�}��'�Si����� c� ���$�QJ${B�͘w$���`�.��� J<%���zz����^w�	J�-M��/|w�ޅ��t�!�	%"A����)H�Z�+���k�C��|MT�>nK�ѱ��8�1�R�����Y�H�?)�U�1Mx�v�jG��\���-�R#5�]*�l�_����M/_?�7dH))�A	H���|�Gq�	���|+`J�%��:|�)�G��F���%B�)G�R�#�굼j���O�8���ow�'�����^w�8�I`IIM�w1����o�����H�Ȓ;���'� �"�$����[�{�}|�J������@�CG�ˌ}��D�� �K����D.�z'���¿f�v�� �b���"g^zgp=	��y>��~iM簃.�����ׅ���=F�/�
��;����u��	7�0d�y�f5^�^� ueNf���c�{ET�^���T���cd(ٻi����]����9�`�ʱ��@�9��z����阱9�k���xy��t�S���	=�%%?W�H�Of��~����)i}h�A4¦�y�r�������E�pv̭j�$�C��b�V}���z��=	�������J�	޷��=�n]����Gq�f��8�`G���c�)D�D�������n�y���u����&� ��H�]|�::"��W�����SD�D���D���_ǲB/�A���$�P)D��Q�n�Η>��Kơ�'��σ�u}� ��D��� �"A	L��K����s�eO�7dI�����U�oWh"�yy�w/��|A6�~"�]���1_tIQ ���(AJD����v��c�M쉧Yk�::#'��*����?cS_qȒ�?$�`�}�6�0B*���+x��I������f��>�G3�\�G�e�N6��X����U��쭥�;^�թ��VomX���tj���[���q
�)`9�����ө�-)j�e�H��+k�f[d�U��,�YFW՘#f%��[�IyGT�8G̾����C�`�\y_r��������/Eޱ��*�*���xɬ&xr�edN�`�ҷ�Sܳn��^^r��Db��S�R�˻��n*.V�J����f�J�N�ޝ�kdѶ����[X�T��K���Wg���{n�ө���)H��Dh":rp�i���}J��he�c��W�(��2��B�A7w.��[v/n�����iu��}�aE��D����l�vM�0`�![�Pb��La�ٳ����[��a8*<��]\����
y���������T3.B`�V�r���YT&���W�%o;<;��pU���؉���U��ރnv�e@Эc:R1�[M�����og����.�ëo;}���+��2�]���ֺ��Oz�K-�o=���B%�>8f�����T�:Yξ}�#�m�B_q2&�neZ���o4Y�QL�cCx��wdj�0�j���Z(e��ٻi��m�l��"�E:���|$��t�b��v��
&�ܸs�)��{J�9]T|4��
⊮�muV�<��Y:�ݰ�⨥�����c��]��K*��L������aKLI��++hv>ۚ���]�ƷW�A޽�\�m�Y6�n�/���CZ��5;̢�N.�p�Z�/��XQ��*��u��ʮ� �I<Rt��(�v�[h;;8��I�prZGI%���y��qq�JQr!� (D��s��̐��r,�&�ͫ;kS�Vۜt#����w��R���{o[\�ɘv֌��̣��wfE8�E6�m'Kf�q�ݜ�I�Eu����;�
[Zq�%�a���D$I�RDqqqkkM&-Y�g%%�f��&��^vm����'3DG%ÑRDgI'������"�'gvEәkj�pB:��D\A'%�	(�q�frw8w�P,�3�&����qȈ��¤�8��mNTqćya���G9�n�����YaAr)�� ����Yؕvؓ�(�����=3L�װغ`nq��M� R�Z�m{5ܚ�&m��Yv�DV���bD3
�p�t�ֽ�C�����H1���0�k�֗���ƘP�B���2�k�5&��h�5Mf���֧1H�i������B�0�ҹ�i�@v�Tm:h5K�M2v3�h�ԡK���af��Ûe\jL�ƌĳ@��v���q�`�ѩ��e�Q)cb�nsMoQ�bs�1�U@��+�b�5��h�1hR�sw[nJ@c�V� "멢�?��3;MhT	�����2�;g9�G����[��!̶����\�U*��3T®�V�F;LGEf�;0�5�4�f*�s1 Ƴ�lu��V�݉�HYi�h,2��H�Ņ�n��`�c\g8��1���t��C���Es1ZW;,�
gGTv��R���#c����u�Vв�� ^�����Y4���`k�@(�vX�ˊZ���l,��h��Y�u)�R8tl��װ�2� a֜�Kn�(�F'h)]�t�uΚ�k?К��q�W��*U9e^ĺ���λ,1�6m����1�����-�٠��8�����Ev΅R�.���h��6�4HY��u�Ќf���QZ[ź�aj�:�T\�1�C]�scMA���l��P���7[u�&���U�YR�M��b��R������4Д]s�Ą��	q�:�..i.��"�YR-�؈R�,�����c�02`�-��˚�g&�.���Vc�ؖZiP�䍷�F��Y0�+˶�2�*JGK�M��MțC��	����S��h^�U�8��������s�)3�^�Ű6H4-���k\Gc[\���f�%ʕ̠����B&�T[���
��a\b�s`Q%��nE�
`�-�y:���M	�ѡ6���np�����:T�k�l���k�\��W*�v(&������ؙبt�m�-�2����M�j8�K2�������8ԭ����0���5�5�9���@��Y�kqM/i�n�M��nt�1�3���W�6V��@*R��U�@���VG[�)�k	�0I�j&�eՋ9����J䈶ʭ
J�77�r� 3kf�GE�aBż8� ���Y[l�%�B�m��1��m,
ƭˌ�-�����l&4����Ui��R
�f�\��Pۛ�6��E�khJ��ŷb���u՗cLJ�F��&5IH������oѮS�tO%�"�cIN5cP���
2����\������$?{�����Qd�Oߩv��<Ms7n^[����ܭ\��Q�#��s�_�2�2�b))�G����[�cl:�}jT*{m�|H�
��u/��|A�I5B�P�h���>S�`I��v�BR$��_%"��z��-_I����x3��O��7;�~zD� � �"D�H�(����1ԴUŸ���ݡ@���
Q#�������[���S\(q@�-w����'_U��+�?Pj@K�H%%?RR'���=�TV�����;]
�w�ݤ��ͻ�}.8~6�A&�QJ$AJ� t�p�xĉf*ET� У��)Mi��g%�!����\�7l��70#��y��皀@�IMR�#;��;�2|���|=��Xs"*z#=��][ӿF��O�)�(���D�&���L%�7�zo�i��d:�z��7ߦ�Gʧx���-�F�մ+ɩ���My�u:���aw6��#b���y�]]w���6�+�M�JY*�ËQ$���sx�\�嗖�S\(�(?=��S��n��,�����!��N54A	H��J>IH�5��u����\���Uy�u/���mĐD����L��"H�г���&����`` �ȐZ�AJD����p�錗t�i>���?En�R#}56$���{|� �H��AG����z�~��[�^O�$�?[�վυ}��ޠ�ؾH�{��_�g۾�3s��U=��<6��ծ��V�sWmq�X��*��,V\fZ�M�~��o�� ��W�H���z�}�2�Ӻ���#���Y��+jc��ؒ)G�)
P$����7L�rq��c��7#!w�p͎��)��=��~�sD�@Kԩ8v&F˼!fz^�¯�4��ܫ��ʖelכ+�۹^ʛ�)f�`���������ŕ:U�Zt�Μ�T<s�s�i��5^f�P�.�U6��Si���jh��P�8�e��u+C7�W]n��@G��z�V�7|(�� K�
Jh��$%�[�"#|3�u,Gt�#�>IH�N���w��6����>����*�����x�s�h��S3.fQ���X9�z����1W"zw-63���9.��?�L�����$b<�^I^���K�.�_���� �Q�hƺhj�K������;V�un��.�&��[�痽�ۈ~����A�~u�{��.��y��PY��;l��	Gɩ�
R^��S��5����8ޏ��hUu-�c��2�ߝ���Đ^:
P}�W8���H!�?���	@��H�w_g�Ƅ�^�+���B����	�9��"HJ>��
)G�م_,�܏]o8�Akk��?�]V>��8�/<r��|� �}�.J��3�����������ُ,-|�����n#���VWu��гo����݂�n�ut�}���XxH��9鵇��y�� �����RS@��s�5����V�.�Y��M�}8~+c��c��� �
Q��w����~n��:���4�[`�z�l[�6�źlE֔h��/�|�v�����~IM�BR$d���3`�Jq�'�=�+��ݍ����U> �jD�1L�RU�Q���O�D���8R�Wh�}In'g<�Gp�f��Ӕ�'|(�?�$����~F���MȒ5̂��|A�%"HJ~��J��[��K�M���?�\�$ا���$B�B�Q �
Q ��
½:i���0��� �٢JD�T�w��-Ju	�o} ��5��aY��᠉��{��JD���"E"�)B{��7g+��&���8=�Qj�9OB��_5 H{"AIM
R�E���g�i�L��յ�	L�^i���(��γ�ӱ2�n�9uK�c���nX/��3'��J����6BR�1��,�+�B�K���X��uL0L���pؓe��͵Q&�,��ln���ecq�J;BR�+z��V�)�����mF�I�5؍k
�:�%��/��i��V�B�R�J����CW!�ơ����
V��]B�)�QYWj9�K{M�*Ym+�D6Ir���0�H�n,F`�mΘm:���k�Zb4\�l��).a��RQ��3z���`�'�&�iQ1�[����c1\�,ˍR˫�	f4�uz�/�����HI��!)�	*����}�.),f�@���C���;^G|A���O�D�$�0A��#d����Z��\���	�M��͎�ԷE<���<�r$��B�9�9�ԗo�'j���@:�䔋(�)E���u��c�Sy��8b:�^�Խ�G���
J~J I	���{{�^w�Ӛ�M�jG��%B���{�w�"�R�|�q��$	FY�oX�9���q�J�R�$�� �����Slh��N]j��::R�8y���	�sD'HJ~��IP�����oۭ�U�鄇�����T��A�{IHfh���[2m�Qa���0�nmW�~���@��t!?���(���(��M��ҵ�^���B�:{]E��k�H9�4A	H�� �"dD��iw�W���yiw�fg]�})�W�Ov�K�$=��;K�%��e�5�(%�o_w���k<ղ}=j{�G���QDe̤|lĿ髰h��.��㼨U:W��&&-Zqo�#� ��N��^���p0uD�C̪� %�����t�Fv�b��t�/61�C�-�����A>�����!)�JE R�����y�]�����_b���Oe+|�G1��c��_�P �@�$!��������%��|A��D���?$��!(�	O��UU��7��nР'��8���%�� �^Đ@�u�Qd��w��p�G�mg��*(Q7�h�IO��Q�)[w�ĺW]5vl�iMZ0i��5�l�+>�﯏�@��l�%4BP$b��p͎�
[�s�=�!'�-�*��F��
y6A� ��'�T(�H)D��G��蝥T��WD�K�ܕ�4psJ�9z5�~w�?-�?��!]����vC�9G)�Ο��d%"~)*�gkJ����Q���8~�n�i����&��1�{���S	���e%�u2j��:�
y��Yrm���W��w���5׽�go��y^Oz�����M�9�bA����J�I��R�g�E^VVנ	����X��\3c����l���k�"�f�.�G_`榴w�w����)2R��?�����߲��LTRr�=��ގ¯+N��~�@�m�yd��dCC��~���O�lpǈG�f�͎�Mq{*�wr6�,�iq�^t,��I�O��p@�g���PX_$b�R�c���<�kM���<�yʹ�Fk��"ۑ_��JQ�J�R�0\�󏗄��=k:~��"qSz�f�9S�s|+zA���~���%ڌ�Vq�j����q$$�QJ$JP�wz=���;3�c��8U��t�k�}@��VȐRSD�I	@ڮ���tΐR�5z~!%B��yn��D̊M��� �������v~���������KmU�C�j����b�n ����� �7ZZKLFR8ۤ�]��m�0\ڃ�]��ޒ�J�8�� �Ґ"H��d��H�2D�����~A�qH��K8gG9N)�sZ+{���)�A�9/	���s�֩�lN��M@�����]�Q�Sb��a,	�*��u�p�x�G3:SWIV��}M(����QJ>�
Q!�|�Op���-��]Am���Eo���?n�@͉�D�/��D�<����R���`��?�B�חk�L������	�R �?���^ھ,Čz���D�#$L�"=��fW̳[��c�帬v�V����9/O�$�QJ$o�-�E�ʌ[B�/bA�Gb����p���-��]�}�@#��������l����A))�
R$�Fg\��>���]
�����ɚ�S��� �V��-*
Q�P�|���6Mi��r�C.���I�=�U�U�VSN�T�V���/R��/���t�u*{0�eE�1Żg��ʫx���]���j��ז��y���9�U�p��X��GBm�:�eʭ3�w15B��Y�\F���i�Wpҥi\1�pǴ��R�٬-T���)Jn,vcv��Xe
Q��ͮ{]tn&��)&,��ʃF$4z��'5��)��\5�p�sa`��e��^�v��&p\��8`@u-i�����U2ZPe��+����K^#��ic@�`ѱ��Q��f�=O��z�t�`��n��lk�TΰÐ�Wm�4baYau�
Y�Yfsi%�K��o�~�"`��I��8^�4�+�Z+{�
���2'�m����|C�F�~)*�(�)D�E��<���'�tYQ#���p�R���M��}_j� ��D����7���nh��to��Y�:'�D ��!��{UO/�4:$�Q8�\v8+c���J>�R��V(G��U��n��04~�"J� �"BO�W�o�q���[������	��a��~�_)��٨0d�A2R$a�*�W��q�R[���
UO���l���HN>IL��bBsg{��k�����*��Z�˄T���1��a�VQ�Vҥ�Ckpl�_v��}zFe�}w���k�6$�
i&Oڨj�)���@�D�A(�R(� )���ew��c�����=D�K�$��O4��&וj�.M&�n�H����%��U����Uo���U�3���ެ��dy�0a�WC�Tg��S_~}!.���x�7�8�]h�������^���Ϧp�\=�{zC>q �u�Ғ�E(�~)FG?M�Y��}5�\"��YM��_�'Ҁ_NA$_IC�|���4+~q<*�(S�(�R'�T(	����:&b�Y�m��?蟈�˝_MS7���DI�@IB̑T���wB���xw#[�t�δN��~S@��D��'䔊[�s|����b,DW���'���G&�j
Bn��6qh�Q��j&�c[vF&�3Q�=;��G�5��@�~ ��o?<���d��YM��\(+�ځY7� A�o�I�s@��H!)�~IM۾b��`�Pt]fh�'ⓡ_	����uL�g1�ƣ��D�AIP�R��3�z�}q�_�`��� A �2DȒ��36$���!`���{�����ub%�W]����Cͬ�gnMڐ!`.��Z;Y�T�J�ս�i������B��ݚŲ*U�[��:��]glY�1���M2悔��Ď_b7�[�x�iBj���~��hY��e��Z�e���,���QWˬ������c�O_ӟ�]X��xM������D���k�-�;+*��۬^6�䷱�:\�U�F�S�+��c��[���4鳎Z���V��Vp�{Km�&��2�R��cu
���뭵��2�j��c�]��Z%&�
�uˎ�o+{W�����k�E�%=�;m�WAɄe�����gph�V�u��{J�V��&�φ�N5N���TI�d��H��!�8h�M�Q����|�-"�7����y	=s�VC��.Ɲ*0�ev]��RǛy\bL���"�{�D&��xr��UU��rUg]�^*��v6���x�s��G-���Ѷ����㌕�cڍ�(Y�۽�yN���(tZ;(?�Y6]�+�u�W-Y�z���2���Ρc��^L:�<���w.��_EK�ƭFG��J��.��KOnr�&AI�)+/&jYd;-;ݾ�Oi��P���r����87kk+j���}+��a�����qU���{F������dWL��y��1P�T�X��"�,�Kh�Y�m�W���dz���`Ų];���Q�v]`�bj�YI�c�:�.cW��������}\��5y]��*�]�+r�&z��(�pP���7AV�=��C[<����"����ro_%3�uFs�x��Y$��m�I �+>Y�RcjC����S�)��������i��P���;��.H$;&����L�:#�(ࣶ�fS1�ݻ��9�����; ��i��J�B̭���*"���m�[Z��9�$q�8���r���ls�ͻ����A8�F��BVv�Rt�Ns����HB�!�P%��e���p睨r�@�$��	�\s�%i���t�y�%&d�t�.�[v�GNr��2�[�+��A$$��� vn-��arwA܇E��t!6���q!��{�Ӈ�;,�m�Бܖw6)8���t�ZJ�����'���Y�����X�*��ߐ'.&"~A D�/���
Q �R��ɸ��#whQn>��M�y���Q7a7�]w�-@�GO�g7hy�^A��S��=�	/�	�&D�%;��q�&!�/���(L�M�1"h\f6��p ��BJE�A�(���O��O>M��MH{��H#0�ָ!+���d,`�u��[+�4��:(�'����h`�}( D�	����)����oc���G�p���wsj���n{_7�=}�A� ?u��J�|R� ��H"1�����tO.�@�D��tf7}�}��J�U�oF���	 ��H))Ϋ��6�c�Bԁy�]?)@I�H�E�xk����>��~��ʒ4=+|j8~9� ��P�R��Q$$�U�̝���O��s�� ��H�O�v�u,�(�\'xH&����;׊����yy�T�evfiz,���N�RSX��ww@l�7��4ǰ^]�+�	�k�˽�&�<��2��S������>���%��v���q�~=�B��U�1̫�9���[�ߟ�,�z��}�tgy^gm�1�_��7�epŨ NA|d���^�S���t�D뀦.%cI�Tp��9��Ѷ5��:kp8�2��@�.��[I&�>��}ݩ�A�"D�2F��{���"EJ����Q'��xL5g�V	�v�Gޫ\ʙ��hA̢ќ% Y���X��M)�^ȜT�Wa��P��V��Oخ~��'���qS`���l_�uG��J��I�Z�y1s�z����/޸M��R8�	!8RSD%HJd=ZCձ�ӳJ|A$~�~!%@����1+�V6��}�:$�龇Z(�D����}��@��H ��H))��$�U�_Hy܉v�����Q^*�p��H'����/}?�Z;̑���c�����fX��ȏC,�M�S�gQ�V��WF,�k9�a4��I젲d�W�Y�뵬�"Y�3Nn�d�U%=�Ք&�]
�L:�}Cs��^�0��-3eL�*kj�/%Ќ��!�Y�қL8��m�k�L@鄕JƸ���f�����!���4�1qf���Y�ZQ���u�]�f���җn�:�K\ZM��aL���l����ڬ����Y��$��uQTۇYJ�Lj⑆NL�:���\4ԍWX�r���(�B��K�m��ؘ]�i���[g��sm����h��^FX�f51���[v��6k2K��_��_��� �]_%%(�N�����BoF��eH�'�i���  �D����2 �$�H�c��:�.�߈Y&�X��������X��Q�o� A�`*i?���vV�*�o00GŸBS�J~����Wq��+�%��.���'%(�V넸q\��$����
)D� ;�{9ml�v$�R���9�dDc3�M�����(F��e���(�+�C7�4C�J~��I�D� �	�z����nI%�g|����{ݼ:b.�aV6��p �o�AңQ̫�1̯o��y����j�u3s��rm��g6��:Q��T
��k.meɪ*fts���A��JlR�1�y�Ւ�
Q���	}"|D�8���yG_5�� G�_!$a�)�J@��}*u؛]����x?G�p;�%�����x-,�l������k*�
��R�bU�$ga'"�t���?q[Fvʇw��*�ϝG�W8�~ ��K�5�dhzr-7�7x
� ���%'{=���V���D�ށ?ޟ��d%HĨW{f��^�<}�z�o�1^0�;>� �}�b�E(�)D���(�A�{&�x�)��)�BP'�K�S�t�"Ӯ�A�|Cdp�Tg)u�b���/�b% A��K�AH�2U{2=OƟ��gtI���uu��vA��ʋM���	������ ���ӏD��ׅ{�ݒB��8QH�:���A�m�m�a-v�30�Q#6�t�%�cl&G�ϲ�Y�C͉�A�܂"D�Dߧ�~�����y����V���J��$i�
8�O�R"H��J��U�~��4�ã=�{.t��R�����21:�O��� ��D��@��*v�������_r�D�X"ff�9�q�Ulµ��t/�YM��è��h�k��u�ݙԭrV��j�7��sr��jj�,������g�j��vM���ܿ1K��6���E�
�7�gz���A��H))��!)Jde�XCw>�/�f~����ޙ���2��h麪���6��>�}�.U#J޻,�ğ�D�IP�~)@�R$��gN���=T��z�g^p��&1?h��8�k�A] %$�5���99�wu�33�f#���=/�
�ղ�G�&04*k4@�b��4M�͖�q)�bf���O(��?wm
(��(�K��{҃�.�o���s�5����@������2 $�fH�d�u��)�b���"�Wy>�Y�{�K�������	��d���7�c�0v�|G�>��̲㙗��e��{[޷�>���^u�e�K&q?p���s_B�/O��
��Z͌�=�����#�hP9�?���Z^x����¹M��ޠ~��H���&S�7�aεr�=Q�M��Rk�J�����1�z��-�n�ת7l����T���c�����yS>���S8��q9SSÀ=�4F� ��
JhJ@I��D�&3�"���rOGV{��M��q�A���%_%?�f�'���~C�G���h\�Zef�rE�+D��J�(��it4�Xu[�������B
�
Jk��0��ݼ�%�^zq;�����{�e��K� ���_�W�H��H ��@!�ڍ;�W={��=q?	N1*v����¹M�ݮ	J�Ӑ@�L����k���\A|C��%�O�� ��O�)�{��cj0�vZ�/z�Si�|n8A�� �J�J/�	J$��}A%iu�{��R��[�?�4)	u����\{3щ�
q��O|F��t���y�0�����Т�}%(�RU�QKڦ������t/��ٝ�҃�
�7�v�P ��?�	����)Hp�q�Ȏ�����3莻ȷ�{�?[�<7صʒ�`���n�|Xy3,��H��}An7Y���oo�}�V7�{J�z�]���C��<x]V���$:�\ ��S�.`K@��-H*뚂��-el�R��&��<�p�ݝ�h��їWh'��5�a),&D���1�6��u���3�"�+���*ˁр���`�c�[�KB؂�4˷���/��Q�cA�c3Z��xio��4 c�K�	�lT4��itY��&�J��.�H��l��L8��mL:j ��\�k+Bэ֭�������1���qE(ۚq�LK2��#tFb�X�d��m�[�.�m�g�P?�g��:D���⒡_Nכ���U�M����GN;��ɡ�����O$P9����HIH��	#^�2z��?Wt�������\{3щ�
|$k�L�����q��5Z�J��=��E��� ���@�A�(��댬����\����r��
�7��p��@�!9R��dA"@��۶c���=���z ��?	����_Vכ��ޕ�M���� Ӊ ���]�(��F�;p��I�AdA|d��������A}X�����bwH&�M|A]"HQ|� I�������Q$q:ê)֢�w]h��dV[�e�XM�ff�;L�]���S��` �i��A�t+�I�JT�7�)��o�K|7k�_�{jȮ�=���=��$�t� � %���y��z$�A���+�\9g ��n�{�cշ:�;-88���ۆ�������UW��mĒ�f����ۢ�f#z���Ƨ�JP�/#���_o���h�K��i��q�N>���_���/�왙0WGݻt	́ ��H))�A�)��ѱ�}�����Ӌ�F6�S��)�t��}8�
(��t��Ov�G�yt(�Ă	J1Jv�zPs����������!���?L���ݬ��9�$�H�Dl��^U�K��������ޖ'�/����iĂ1)�(������[�q��Q��i4U
e1ں�]Bv.Q���k�W1β��b��:���>����~>��vȒ��!(
����p4��э��mLz��ϟ���rꟘ��Dw���$a�%"	��{m*��~Y�<^ĐJ��)���A��c��n�W�(/� w �H���ڿ%u��� F��ɂ�/��/��0{��?vU��,�ᛊ��w�]"�5�{1u�&�=��t���>ز^�]׮=P�S�b̚�.��+/t�f�:��Zv���6��ѓ���7;w���7�Z�n�vwG@4�AbU�Qd�I	*"����b������A�1~�� �G;�o;��s��mp��	�)�F�w����=��8{�H����(�%(�AIP�R�	���J�ĥ��~����}�����-�ݮ	yA��O�� ����=���[F��K�	P)�L�K	f�[m�d�
!�MZU�)h�nZ��טZנϢ5� �S@��$%3�IPښ{����]z'kO���X.o�3�,��EQ?��D���J�?]�<4��4K�cA�9�Fl��{y��e�zq���	�4A] $���_C�����m
7t�?��IfJ�+=�z��wK�v=��>��o����@ �"~)+�̲�3(�[ߚ�o^�n��=�,wO��	*�Ϸ�ty��C��q�}�Ӊ/�f)ꃤq�˞�U&��ש�	+�TjjF-��_��N�:��f������U��<������v�ʩaW	v���4\H�x4��Q�Kq ��
�(R�%%.�|;c�O��'��ׯ�Çz�z��H&�OԺD�BR'��J��������������5|#��oX��[�
Q��7-c��]�ؗE�]?������|$��_��J,�J'䩿���6�p����Px���{C�����jD��k��.&e3.w罼�|tM�˝�!Կv���b��xߖ�G|A�I�J�1�s�_����w�+�}���A)
Jh��RO�u����7��~�D�Z�V6�S�'��5�.� ��~?%�V ���/Vd����_XΌ1��H�
Q %\�^��f���|7k�P'�<�F�h=��}��{dO�%~))��H�_�٘���0�вB����Րe�d�x�x��/�5�ݤA;��H!$�r@!	'�� ����BJ$��@!	'��I?�H!$�D�BO�I �$��$��H!$�$�BN�I(�BI�I?� IN ��� �$���BI�d�BO�$�R@!	&I �$��1AY&SY$z��'Y�`P��3'� b�>�t��  @(    J �@  *�  �   ��@P�  
   
 � UPU
 
*� J(D�
�D U"��
P(P
( ��%"J�P
���x}UB�J)A(�����T"$*��D�%ET�(������$TJ�� PJ� ��R�RR��  U(�%DTR)P
� �zY�� �U� JA��N�t�&oA��@'g=�z%�*�0�!����P(P(� 5��22�a�]��|�`z��� ��<@ w�*��  ��� o{�<@@=�70@�	�o� ��"�IPJ�$*�"IJp !����lV;�r�ӓ��1� ]�)�Sѥ����`���J{�E,�.f��K��
E*
A� �}�����H�u �t������B�=��^l:5WzA��=9;� �A^���[��궬�J�*�  ��H�B	H*!T��<_U�g%���#��)�yR�B�vw����x@�]���g@	�J���@S����� PR�_  }��w������n�B�;��{�u�]��Ҹ�@�u%Bp=���-���B���Ow� �@QQS�   }�R���T�
�Q	DP|� n�螀��Ī�@Q�0 t�%EY�`!�]�9C��(2�R�J�^� ���(�5@�>   ����G h
wH�� �w�� ^�t��^�bv 8��UF� ��0h<@qzΏLC�B�RHK�  �
T�R���
�!;�7a��>�-�F���Tz4��S ]�Z�"����� �A\�#�
���� �/�  A���B��^�����
R��#�@bt �:������J% �=  bz{ |US��fJ�SM�ɐ�S�a���  =�M��@  M��*h  OT��  h�x��Ē�yOP �����O����A$�H����r��_xu��$��	*Q���$�		�J�ն�6�֭����նkV�j����� ���_�5�����(�e���ƕ/�?������(�7j9l��`LAb�Hh��F�DD3K�Hnm��Y-`�h^��{t�nL�1Y��8����//\�.�[Gm���j��l+8�k����ӕ����s��+8B^M�Tߕ�5hh�2�7��I���d�*����w5��][rdf�|��'wn��yk3e�V����}`�k��/Rǌ燖�8`̲PX�I�(��@�C%� �ݜB|ޠ�nh͠�V2<� cS-l7�X�/Xُ.yku�	�J��D�r��vc�*50V��t�(zK�	�cp����n�R�v���BAzE[��h`�K~��l�<7/0mn^�Zp�X�C7�UږP��	Vխ@
-�fS�W���i�-"@�է,i=r,5�k�Y�ܡ�����eLn1�2�P�h,�$n�ȳ4bN�0��V��R֥n��pe�&�d�:.�Q�{zwbI@ֱ��2�H�ܺ�쨁�Xʺԅ�兕n��$k2��&�����6m`D��7B��iQ�W�>Z8-�ؠ���{iԲ�˱�����$T����W�1��^� �~��	�H��6@��0i��9Y4fT%{`�2}�ɘ����u�4��nƓ(]�Ҩ��6�рh������K/ukhaSU[Y�i�r�T�2l�pa��nR���֯4�&ٶ�1�4����P�3s�/�V��U�\��h�X\���@TYxH1�q\���ǚ���d�f	V�"X0�,9�M��q��n�� ǃhn=˧xAF�+R`� [��6�n�#���S��fi�xu���)"�ef���� 铍MfڏoF�M�{���j�aqU�[��<(����*v+��˭[H�?�,��0i��_�W�e�F
qc1d�R�L�S�V1�6im��|j��I��8�-��m���*��8�y�`��l7n��N�2ڇ\HF�:�ջAn^�sp:ˁ�u{��P�09�������̖S�tK5f^;Z-����\7d���Y�JvnL��7#5u!l�m��s3+,ɂӠ,T*����,����[�G�݈��-�W3(�	�����+v��r�n�ѯ!����ag�5��Mզ�G��Z�l�ڛv��;��h�:1cw�cW�҆��MV�"�FZ�l������^R�.�&\�{-GK]��*�֙�����U���������cr�I"��V�]�1� ������Ι�� ���v��>�h�p�@ԕ�5Kl�p�ou���zȼkq����������SX��f�	4{��bD��������~5��@@�1<Wx����
�����`9���JB�����e�F,��hmm8j;�En��̀��@u��kW�*g���)Sn���Ke*��t֢�ʲ0-{�Z�e�%����E���T�u\Ź�f*�-�V�3[gN�Yى�P̺��L��(�.0m�R�)M�#oaR *�fSɺ��궀ɲ��u��yL+NX5��9��˺�#kY�Ϝ�t�i��A\{��k5�Y�K�4Y��lK�(�tjW{���#V@�ugp^��[V�4Q���f�P�d�M�4�1B�U�ƞ�dV���y�Kv��I� 2�W�l�k~�2-"j�U��WF=�����4-i�#��1�u�֭5���w/.��Pݕ U��+C%�YreV��O)�2�meջ���"@��mmn����S~{@8�cXo+s�Q�y "��WtƔ�VK���1:��K�H��y��*F�^�U����D���a̸�I!f**�B]��4��-A�;[yz	 &�X�܄�R�޹�V��J�a��
5�%�6��u��QЪb��̀��^⫗F�L=��n34),ꅪ�@Zn��XVP[��I]��U䌑���j$�����*�H�ɛ�a����+~��
�+,��H�IF�a��JiKu`����k�)��1up�6!��Y��oM��ILok#�+tMn�5r��I��m�P^�g5}y��xM��^U��CIX��R�X2�ʓokef��t�;�up[wt�[զ�����9y���9Ug��n�Ȫ2�kb]��T��唜����Ҏ'.E��md�3a6�`�ͨP�ȴ!��XXK+n�%2�;)�<��1Qe�٨7��,TBZ�#^l1*�U��%<���`�FK�Ӣ.+h��R9�Zf�'on���W��|6�+"ƥi;7g~���Kl<�m�$)�$�,������a�D�dW�7��):�Z<�Xʴ��JS���ѵ>�W��k鷏>�@4��ʺ*�|�Y j�H{q?mJN�$�lS�D��;c\b��h3Xwj������e�u�ڐ�WB�ʶ�h�m�y�FU�ڄ�a�.j�*$>T%f��RC]�Ib�s.2�p�F&N��W�F+�J=�cū4�չcMO��+YF�^��:T!�7i J�ђ]i"��閯@n���ޭ{[��P� u�6����v)�fQ�-\�L�^Xw�df��ѶVZc]�EY�W��Z���&����)�&��ݕ��AO-�])O���l�ӱ�t�۶غ����Z��G7.|��e�Ye��ZLܐ��,�8��Z.fm	ZMl�Z �6��۱u#�b�9�z[�nꓼ�i�P����r��N�N�6I��6,�8����&��,�`5V���Z�y[,t�F��9hk�9����KQ+ˆ���kQgN�չv$$�c#Qa{S(�kfi�xv��Q����XS)���,F�$yB��Dt��Ҹ��y"����b�ɬT��$nT�Y��I���!ֹم���zN�*�Z�m�O*��,�O%ݍq�85������sV�XwdVE�I� �:����&T
�Z��{ �����
J����ơ�T�c�����5�J�l7z#���=-�f�i�
�r=5����Q�L�%�p��))�ǉֺM���߅#Q�t�OI���w7m���sEZ�u�w��K�/j-`d"��v�'��,܆�ˏ^gv���A�^���Jx dt��8��5��ٲ!r�' ǹ3;I�W����p�6���ء�G��ʺ��**��֓��.���/,)��o2-ͱt��H(�pm'E�`YX��H�7t��0"�^Y5ޗib�	��3L�JxqF%L�* ��͙3C[.a܊�j׵-IW�Ht��d�E�ש�����bø�A3.�ʺ'E�o5Q8�-����^4-�ۻ���I�hTa ���kz��ع��*�6^C��	�)�Lz���X�pӔ�eOS���݆3ϙ�8�n���ə������� I�?ekēb��q�jM�˩-m��|�k�L������{��%�=Mׯ�YlR�E���j^�4'�Y6GVTr�Hk2�,䠯"��=x�^���Mk���*����.�� �n��1�n*jkt5�j0Z��E�b�)_��eg�X��:F��N]ڲؘ�m���9A-uk�*�񥈵��Ua�p"V{�LԽ�Wx�n�q]�ML5��Y��דi֝/C�Y#{�����첊�4& k��WW0R�`VJ�6�۳b���4�P��$kq�ET-j*��`׷/���Y42�
X�u�[2~j�ԖQQ�
9.����CFl�`ӻ���(�Zg1�D&&���LK�,���af!�;J�G
�N�VN�ɥ,�T�JF�[ٮ���pm�wP�S:��m^��B������,�j�]�3\����DAT��%��E��{�ڽ��\Z�Y5u�Դ
����t�#�Z%5W�E�Y&�k���@�Xr��F�ܿ�^dZ�^�^M�N� �"]��t�U�Vr�g��(��sj�M�շ���ރj)'1�bM���s*P�ka�l���47]�#�^��f�bX�JŔ�Io>4Y�+�-?j�A��v���5I^��xխ�֦�$�:��ݭ�i�M?^Q;����(���+.j�
��hn�����c�wP���묤lL�����z@����-nkٹZٺ��v�L�BVS[�S�̰]��cY�X30_��n��7+-�Fcwzp��BFAa L�F��C.%"�nŜ�(틔7O�Kl�x伇L�)�b�Eҡx)����r�a�N�Jk��-T�4KM�5+TAʰ��M��BmV;�h�lݢ�V�T���"��%��- t^���m�] ^��[�[3V͟1�EdR �9{m�ԝ������b"�7$�Oi:��YDq��m�&ٶp r�%��U�thՒ�i	��F�[E��'8%���<E���I	���ZQ��b���	�L�ĠR�5(G �[@Ց�ŷGt��L�Jؘ�yz��Y����*�9��Y[$;C �U���u��`S�	�5�rڔ)�9YJ�AIA��F��#�-6���Gb^��ť��A���N�Z�+,�t.�D�K�Q�&����2��xwN^څ��,�eʚ�ݩ��:�ǔ�T�:� E�`U��yH胓�!��Vc�	����bB��m�^�͓4�x[ٸ��`������e'����V��
�c+��YV���+�K�cjee:��ƍ8N1�
ӳ�Ucʴ)AW�7�n����6�+�>��j^p�A]ۻ8w+.�Ŕ���H��-nV�u育M�E��A Jp�(]ֲ��I���[̚	��Q���E����]I�/o[خ	�)���r�`˶�O^cY3h\=)����ÔQQI!��̙����M���K��囫���4a���jۈ�w�e�˘���k/��V;�i]�h��ې�w���7��CB�5�����j��<%�y����Xt�j�`����Ճpe���ov��lCu�SR�Ѻ�h�fP9��Q�8�-�ʴ`��y�V����ߝn��W�)� ٵ�a�:���m�a����10���^%��z��b�@�zI_�8����D���j:م�[6�Y2�����[%��7v����%��sأp�ow�z0�*�f��+��.S3��۫h
ڷ���9@�j
R�S�Z&�7�V즈��� ��U̘�'q�י�;�1�*^�gٖ��%��:�[{M���0-�W�%�n$u���ۢSgC�y�ҵ}����[�(P��+6N�Ӣ��@�-i���%lX�E�Y+�b�=�8��-�&Z6F6^�FVi6��u���f�V*Q��
5��ss~�5�TTRf����n{4� ���X�i&n���X��<�aA�ܢ��מ#I۶�ʩ�bЀD�X��z��X�e�;�槻�#t�
շ���%M� ���Z�3l U�#A���3)��&��ε�f��C[9**�aٮޒ��y-��d�P ��\�tTx��`Y��;����=s,X:��SǷ�SB".u�cD���A�w�
�p�%��ق[��G.�'v�]�I
� :`�?Eܨ"@Q�R��H�GL�0|E���J�k���2��|���Y��t@�6h���y �F��(��v��ײm���8tʈfch��f`��AkR8���4�3XX�X�17&b��J6 ]��@��Px�H�]a��� U�4J���t�2��.^�b2Ӣt_�McqY��ֹ�k��D�-��P�F��&l*��ݘ���Qa���L�hŔg���Ķ��-�M(I2��������%��,�i�*���TܩC�(V+�`9j�T���0"�U�.e�ĮSWb�K&��ˏ);��hR���[�%W�)Jْc%F�)j�JZ��H�F��uy.]mK^-�f��l��yCC'��zAcr����U��
�m�"�f��ŹH�f�L�a�:.�A�=�P��W�
�ʛT$�+L.9+N��{y0
L֓�� �Ʋ�,,�jUH2�n{�Jd��a�R��lȶ����	{�P="�.���$��Glw+K�/"��0����u���,�ܚ6f�m�i�թ�ej4��x��H�/�K�(�Rզ`���P�R��h�0��H�*����\�-�WiV��6����7l�67v}�uyX���\�B#nmk4l�7<��Љ��݁[��	Y�)�f�h�Q�ag���0)��BЙ �*1{I�Yw��6*X�W�iE��n])MVf�)e+�"o3]öA�u��S�9J^���V��A��������j�%�yy"��O��XSR�˼H�D-��0F��m>��(��1 c*�h�Y��mf�Gu�NFC�*��*�U�Q�"�Z�6˛w����c����C Q�����Z޻���.�1�ʺ�-�UnT���84�AA�`R�[ڏj,�i[��L��;�a	7��0!mHUd
�w1MY��-d4�;�]R�&ܠ��$�ǻ�$cn���Ǒ*g�nZC$��X�j��/c,�f�������
W����m�{Ѫ�hW2`ڠ$�k1e��J�+`�5��WM����M�q4�Y[�����c|2�i���z�2V�q)m�]r�nHYS0�ݧ��U�! �72�L{�r�C,��0�X���t�BU�fb2��Rk/J·A�S��V˲��#sR��&��)D�+�WE�xsh�h�hV;�˹F���w�虄7J�+lTn�ɥ�gTJ���l܋7+ �F��e�j�'�#���3Qn��/k^���3a5����)��M�m5i�i�)��72��l�c��< *�F̺tp�!��d����ۦq�*�KH���j�.* N����"�ϠE
ߦ^��\�%�]��Ɏ�g&�Q��)/4�@ I�X�-j�Q�Tm�j5����+Q�6�kQm[F�Q���mV-��cUk���E��j�V+X�kh�m��j�����+Xִ[F��-TZ��cmlUm����b�Ѫ�m���մmm�j���լ���h�cU��j��ت�Z��Սj"�ŵF��5�EZ����[U��E��jŶ���-�jت�����6�j����kQmQlmF��kU�*�5kTm�cm[Vѵh�h���Z�ڬkZ�ŴU���U�5�Ѷ�V��Z�[[_n���}�����|=t?�����u)��;S���2��L�7�esco�`(]v�,��$��U���l3E�ڜYAM"���ׁz�4G�F6H,�w���^U7S�ͺ��#���n�Ҧ���j��
Nճ2n�����x�%c���]�v�8��޳�#Y�*�+�:�q��B���QU��,���U�JI�r���[p;�#�����ޜnt'1� ���Ż��X4|D�Pu3�2���r���vҶ48�`���D=���^�H���S�.P���;�ZS݁�t�)��vs,FN�v}jD>�z��gx��˰��w3%���fP �s*�9b�om�(�ދ�JY���z����]������*���v3{[�K�2V�Yʓ�=�u8��@�j/>����Sn!�E��/��[��=�i+�������Aݚ�)W&�f�C��̂�C�Dk�������i��J��}��r»��	.����mp��3:�F���M=�g�kB�x=��h��I�t���.P�|̫�gG(Q����SB�!>��a�d'W���t�Uv+f�A��:�O��]%w	9��\����*Ц^�tBmM
�dE�0L�Aݡc��u�'�f��w2d�6������u��#�{�nI���]}S(ro�Oa���W/d��4��ԇ2�Z坜$�+�u=�F�ӵ�3�
F}x�m����VV�c}}�A�5}�X�����Q���g8��Ij�me���)���7�)YV�6�54lv"�
���td�έ��sm�udQ��4+��d�ʚ-.����{8c�j�U{c�EJ�|�C�tՐ��(n�G�{�I鵷�dX�%��#6�ut�M�ۍa�Z��p��ݔ��j��類 8tvfo�s���z���V�4,�!x&�_mW�򳫤m^4f�e�ƁM��՛�4�JدYTD8���5Z�k�X,�)��i�tOH�-IZ�{�>�6Ttq^���#ro_ƭ�d��q͡2pM��E1��Do�P���7־2�1,��^��E�����G�o�������Sv3g��z�.�V����3��L��hc��}�>���Rp����h�wr�!�7�����<�ي� ��"��aΉfԮ}PΥ���5�V��7S��Հ�8�P���Ҙ���.�����`��jd��r���	�KFٖ��U���� �F�x��h�\��CfJڔ�KQ+96����c6�]�dT��M[%��f�.f�-H:�F�w{5p]�b5��{jU��HC,��-#�vV�C�)pp[Yh�#��	�{++0�8f�y�Z����P��G���a.b��	I�wJ���qh�����#t�/5;T��g��X����Cb�,R�u0o'��-B�k�f����1�ѼF���v�b�X�쳄j������OD�y��VC�6�k?,�ա�|r�S's� ;�v��cmnR��n�!�؄�L��]|���-��c��F���H�q�qFإ˔CJf�����]��<<�m=��tT�+=S �?��)�8A̲r�v�N��(T4���4't��̹u̻	�qYn��e<!]wwå�s(Sn��V�'B��۔���BoA'Qh��y�ڬ���[9�Fmrh_^�4q[�[�8��˱��Zw\�N$�&�{�"T�FG�F�ʙ��:�m�����.t���yVE��D3���@31)Ju�Z�3{:DM���`6_-���D@�)�!��]�[ÐnU���Ce�I��=Ԙ�R7pܑX�C7�8n���+�O�	�;�Ջa���1c��=B�C�ټ)���&�N�x��H�8��Ӕ'(��ùy�`��m����z�ZD*Ǟ�/Y�L�t��9Nظ�`�.�҅M��gQ�0Y���\X8٧mt��n�7ל;��v��G-������SF��MV¬�ڌ]�WJ�@�o�IC`��VL�ޚ/Eދ;���ˢ�W^b��R�V�|�M*L�v��B���3��Ƴ���WB0c7���F��q�7�Y&U�L�ٽ�y1�g-.���L����ok�'mbB�%�M�R��j���V�ӓl��l�':�u\�p��	]�)e��*3w7kU�x�օbI�s���QѢƕ�3zf!�G�8&���/y�,��U��@���.��Oŵ�i�v�
�g����а�u.��W8��A9W�1�,D����TW��3s�Rdz�4N���H��!xr��[��W�\�{�j�\�kvz���KH���3��4�Y���$��ŧ�e�Rj�7��Q|3xb*����]�d���W�]�{$�Pi�[�w2ʺwӼD$NEs�Q��<�'���F�������EFZ[�zy���{���M�5��N�GY<9c6&G7ީ�!9�X^�޶l'��k3/V�y�G!�V�{���^õ��K+ś��;����l���Y�����;��w	Z�X`	l����$�^w3�I{�+���2�o��g͍�,^�����(�����ˆ��K�4�Z���H����g�p��oΒ��{��h��cCye����6�9h����,.�2﷬�De���2U��(`��/Ž�k �j�*rɼ&\�K/n,�����Vf��5��:.x38�ޤ�Ҧr��p�«B��R���q�eJ[�^í��EkY��h�f}�ݜ���
�g�K7R��а�Uc;Czu���V�!��WZN�����C��;h�L�\E��!��˗@��+�����ƣ�=5P���r�Ǜ��t1�2-�
ܖ.r�Zd�vS��5vS�4�������q�]`�XΫ���T�.9���������X2�v���^�i�+�R��9Ù\ܲ����I���Q���c��y@�����J���.�;S#ߍkOVm�/9�̓�&޺�[�d�o�#TGm��K^��p�%���.���#�j����/2pqL �5Soз58�s3��>@ܶ��z��m�R��Or�h���f�b��W�p��Pvk�l{�"�O�/_�̳~ߥ���Yʏ<ze]��T��o�vw�H�v<<���&�J����x��IY��8_�`���^lnV�4"���O^��<�h��!I`认�jW����w�'�8i�*
$V���v�]��m�T�S+��d�Wz7I�����x��j֋�;Y�8�#���{�m(	�wq�fݨ���u�&�[�=�pU��25�)'��j�LS�d�� |���g�����8w=�Lu����2���:zi. �ͥծ)Z,���J2]z���^Y��[C5��Ij���A(:ы:�=7,p�f�c\�֍DY0Kvr��xvR���]�D��}m���u֓�N��p�v^,tI��e�"N9�u��/]b�46wq٠"߷��V�t�2�,l�R�l+ ����[X]��J�:��DgV֩�0�����g)�6�@Ҝ�7����Gus�5s>Tc.ӆ�H���/|�CY�V�{�%�"�V+Df[ႃΆ[�)٧r�j�IVge��Ph�
8uc���;��0P#�Y���QJ!<��h%e
�t#]�]�-@	i�
�tȋ�n.�:�.�3j�nA�sG9�"�����YXM\''w��+f������YIˎГ��ʖ�f����/q�C��g�A3�Z��uL��^��Ȟ��q�Kc��ﯮt��d�`+ۼf��A�x���(�RS�_�/+;���+kOAR���V�dV�a7�����r��i���-j�Wt�̴)�Ǡ������! صi��U����!}�IGF��T�w�h�)�/�H�vd�6
#���ZGd�)���J��i"p��n��d/�����=W�_1A�Y�J�s�����~����v,z2
#�i[���і�FV^����E�ك���봕QV��tbe���N�M�cW-���N�Wi��LJ�/;���e��j��v6��l޽�>�w��m�&�$_q��������q�x��YBjt�ox]ňf
�ˬ�β_�!2T�N�s2��@A�+�rW�v-�����&�3f�m^��.��E{�K5�>��� L:g�Z(����0�Q�.�����>�5RK�ڽ�aR��&,R���fs�蠳^_ ��Y����Ƿ�����l	E��g�(��1�e�͙*W ���V�#n�	j"ҠDCo�*��j��ne��G`ia�֔^ZNd����w��p(.=�]x&Kq`d������Ð���Wb�]f�[W.�=�U���]�2��2ܣN��,vw�W˘���P���=ݫ+xWS=���oH��{.q�-�"fa�05���!���W�YOn�l�W����u=*�5���â�k����cM����,�&�F���0�p�n*��ӌ�z,�\w������	f��3�ٽ�u��z��=L:f��.�%կ��Qӳ����)\�2�����3��ZѺ:T@Ja v��-�Yy�!��7՚яo�à��m��צU!�<S$->*Ϸ,�x7�+Z���b`�D�GJȣP�NO������ØJ��9��S�
��r��'%�D��wk#� �g.|n՗�º{�<�N��ӗ�+�����˓R�ʞ+��t�ի3�n���wr��v�4Ր�賬�3��4�n��:0L�a]K�&��-��Ճt��K@��avi�!��/T� "�R�ڭ��vޕxO`j��U�U�n��K׭�&�R�%�iv�&�9�-w��+��o:�)N�JE��]�A��b���e��.s��a�,�P5QJ��U0�mJ�w�U�`9m��F�jn.���s�E���Z�<JtB��!��&�N�ޭ�%���5fF�5s7���I�����1���P��,�!N�B��j+����':�q�:�����ݼ,�}��bЄ��|�g5�A	%4>,X�S�+��lˬ�v�I;`̩� ��z��^�)v��z �9b��Mf�Wg�w�n���()��x#"��u/�Fn�
�]4��]�ؼF>{z'r���[�Txޕgt�7ҥa�0�ߤ���Hq�(�4(�yR�"ξ������v�I
Fu���]5xf�p�r-�����O?�«���.��@ڷ��v��ӋQ��x�6Ħq�*L��e<K�8���$�%�V��u�E�U�dIAYTӓv�P8*�ɒS��o�3a7�U<|�f�a�ꚧ�������z��L��*�J%
f��[[G횮T�Ks�l`�q�綆��{%iBΝ��*�4Q���^y�Ɔ/FP�����׀�@�l���}a���K��xX3��Y�à>w���9f����e]�C&��SxJB��^�����qxI��#�0��̭Ke�e��;0Xes��i�*���!TiܱsoR�y(^j��T3���s�8F�-�gtٰݧ;;
[LoE��9ٮ�6����\\�;��Gv
Ѝ�ݶ8�F�]λְ%D����{s�mىa��%�b��������E�����ц��if-���,�,������I6���������ח�e��[��s�םI�z�	ϷW��ڦQ��u�G����n7U��h���9��U-N� ^���ϻ���uq
Y�;a�E�ʝ35�������l��l{R���E��,]��U�(0�z��hV���*���(�x��-Ϧ^��X�b�m�x�I��f��&��w�ڗ�εh�K]���N��+�5QfD�o�+�Wa-M��WlQg�	%��2�0�e؃��"FI�k����t܀�8��Y�=a��4w]��8�,����}ih�B^����d�SvTIL�r���:��YkC�Y4��U�~7�=i{qi�i�6�0�XY���i!Ia�4m�x����h�q3r\��Ц������U`�����l�N��1�`0[F_���ˡs*|(fR�f]�7)���7ǯx�WM����-��<��Ĥ�J��$grz�I�o(zV�v�M�+���g�h]�}��&�Z=�~���n�ܛ:֙��nZk@B����PX��i�m�V�hn:���݋;�7ݭ����T�����泓%g�r��]�ۥ�6�������Q�9n;*�v�/��s�V�Cs�&;�(�ښ]]�����A�R�yI=݋nS�/��RnKG�7Β^�R��ĂI-�W���<1��)�hՇ0���V�p�e�٧�W�ʢ�(|&�+3�1wr��Z.���+s���~w����b���C
aK=�򔡄d[M]\�;���4��� �b������Kۡ�Q^�o�����u�㶆��w�v�pջoM[[y����BZy�]�/�!��o ��һr�[�Q�y�U��>rHs(SԽ&Bl��9Y���ͬq��V:�̞�ɯ����3T��q���Y�dfv�{�g����/ڥ�!W�ݵ�Y���gu'󳳡(ٝ.r�{�ƫ�8�&gXcKfs?JG(]VC�[9��[8k*�t⩸f�l�I ��m|�R���ҫ͂�����X��Җ�f:�h�U�"ZE)t'gt����BJh|�����oB�KKW\�mWg�H��`Tw������ȯ�X׽����f��2˫�fe�p��,�$��p�l`7z�U�����W�+��)T,�]�Vm!�EL���ŜSP�}Ј^�)��ʕ;]G�1�[z�����b]:{2��&l�'��D���й�����q'��C�&�W+E<�`;x/�y$�Z�Q�,��G5q1Y��@����N�#��<������uk�`�����wN����I.��5vV�)�����efc橛e��aѭ�!6!���-�f�5�6vfe7\�MV�u���Ԫ]�6h,\�v��	f"ӌ����_���H����)X�\1c�;SR��-V�SZ��⎍S���v�#,ւ��[K�l��8	�2�����T6��)�,��f��ս��xD9�Xې��XQaBi��G\+ױ2�&sYX���гF� (�R�!.��Ę�[�Q�I�ٔ�uf�����r��ͤ���"D*�Y�[LَV_��ߒ궅`˘����1W��B#ٸщ5����HXʸrr0�����\]f���*�Wˋ��.��Bml�X]H�`��d۽����a�R�`�!��YEp�Bஂ3kW��c<s��1h�Ж�]�΄%3].6�b�����`��BL��Y`t���hiI�-���&͉.fc
(�N���̻���f��ʆ�K)�i��c���VaofR����]R!Aj����V�S�h���F�1m�Xܗ�C4�쀍��Z��)�L���B��L�� 6�!P5�nâ���Pk��h������.��6JJ��iiY�F�3Gm��lF�"��B�����6��z����1�st�0Z��lfXE�l��J�;��(J4���gm���e�4�r�vCLL� VFP��`f����ͻilu�,�����b k4ت<�m�&���� �GE��uɠ�fX`���$��X�-ci�0%�)�]l[E�N`��K�l([B5���
<hf��0�!�lٌt[6"�t�1�ں�]�f@09�!���E��-�1KKe��B��`�QJ�������4�-w*��#�P�ur��,X,�]6�f��,�,�`���UJ�%.��˝e��桍r����@Me �%I�ѺR/!thXcMh����")[΢l�	�iaHgKe��M_����_r��Y��J��s)WU`d�����6�bS��Z@hE�F��b�n�Ԥ�M�k4�[�[����8*��s^.0����Z�3[Ʋ ݭk-sr�%@��	�YP��RW� �i46��bօMZڒm��U�g�q}���05�������Բ��B]�9�Kbie���A�����R	*R�.��u�]�:�i�h�!n-Z��k,��c3��+�!S���gm��l�SR]��2vʖ!6�u����cm0�F[)@[m8t�ټ���"Qt����W;K��%����67J��&ᠳR�l�1��wrl���r��.��Q�K�A�i��kr`��M�X�M�ilh� �le��&`Z�[�8@T�ڸ�W8u��=�h�su#LK4bE�Q1CHC,� �b��a]+���&�@�cu���aʜ�����m6A�V�j��Mn�庆)�h�5F=���-X�h��F[�/j��Y`�1
`�m5:M6�fրg��i�u;h�ٱQ�)qW���c��Y����g1��^����˜8Ne��,�-ւ70+�*�b鋰=������]56ġ.j�����F��v�˱�����]��M˕#�c`Z,��]X�
Jc�3FY{]���ne	l#6��W�ke�!�C�e[6ob$����� �!�HYa5��ۄ��!��ȷFR�4sl�IB1Ia���kj�a�{)
�s+,�p��k�)e�<ˑ��j��5236�֐����D-��E!�+4�v�R`��1�f�1%�)euc�,b�(�6�hm��h��t]@1b��x�bQ�J�<a��8AT���b�``�50gX*[��G�\�A��p2��KF-�f�K5P�������ݥ���*�G�:hi�`5u�]�u�	�LdB(�6���hǮ�p,��p�]Y����<GQ�u6�7Cֲ��b����+N�6&L���[���ֲ����]j�k�V�5jj���2hl�]e��R �@��R�ʎ�k��˥�/�%�{h�$^�j�mB�M ��tZ��l�`J�R�]&��;j�d�e�
iU&�b��]�ir�,c�3�0��s�\��7@eҮ��m9ʩKE�Ȏ���5[.W�]��^L�R���hK.��R 5pY��M ��E��`�L�]M�JjmhB������м*lS�2�,����+,"6Yv��6�Z�%�&<�b���	(@ͽ�rJ72�Gj�3`K
�tX,�����ŋln�:��uAJk]�Gj��Q�s=�����;`n&]�V^�2��3�f��f�qK
c;5v̫pH!u��c����)Y��̹:�\]��ڕ�����jJlWm�U�����d��a����](vlbےj� �n�Z�glX=j�sS&����5�,��2�M
��isy�L��f�5��#ui[��Cn!S$)���,��f�Ya���r�+ CAB�,�۠�ݶ�-vθk֡6����e�1r9��f�M+Yx���J���)�1#{h��T��u��a��,�+��M`ˆf]��3�HMn��d�WK���aΉau��R�jE�SE�WJ�h�^��E��A�&�ճZͦm����F�cf�P�+��D3�,Wh�MhCZ�B`"�L��pk�h��%|���s+���R�j��knD�X��Ѯ�	��T�M�3�0讃a��	�0*u���7KuټL�в���4lh8�&�u�1�8��bƖD�5=�O�����Ze)���T�
��{��=��Kb���h�6� �2��͸��5M�����5f�@����2g;bj�9�h�m�(&5�r�0�c�ׅ���&�b9�gUK�nr\a��!V鈽��:n���2h�ˀfwlijB�n*��G8qf�hsMt�[F����I�f5bTA�5�gj�ff;U�4�	�5�c9��t��Q�	R"FR�0-�L3k2�!����ɓ��j:�!�.�kMf]��ha�4�kY�#�z�tб��t��0�b�\�x�7���L�-6�ۋB�H�wR�Z�i.@�+�J$�%c,���&w9(�e@6�ML!����\�����\cL�ےԎ$*��[6`�XP�Hl�����B���z�%!���1���Z��1Iz�A;kP�"D[�����`3c���������^X0��ݫd�F�r��p�ko#��k��A�i��*�� �چ�caTK%ͳM-��d&nqc���YK�^��B��m0�5��#��%	W �Zc\i�me븙)L�r�P��Ֆ�c�f�:�f��m�����cF��c&��#t���j�(ٙs�]F�)6ò���a`���ִ��2h��YVB�3Ui+C#.�[..��a��i]��Yv�gJ�t�C;a(���ٷd�X�+�!q����L�e�%�Rb���v$��]m�+U���u֘V�X�.�⻴(CN52�`c*]�֥�g X0q�Ԁ�fi{P�*�e��e7^��I�YJgVTp�1��se��%-�{�-8��3kuv�Q�[�=���Ԉ8�Q�#�Rí�ַ�E�R�&�+�mX�M,�����(�է�|��-���[P����ʺ$Z�A�-��m�����`�B��̹�4�u��k��ҼCcRY���AՂKM�Q�
mfU���3���ITwiu�KqY
��%qB��]�G4�m\�����FՃ^Һ���e�
�;FWA-��F�Y@"q��&�CF�b�U���� iT���f�d�*�q&9�lXN,��M-l�j2�Mca��yN�Ra���mt�luC+YS]H[���j�.��SE-c(]ZLmEV�g�����e�x����Ȍ^ckW��)����+ѢSL������5���f$D�K\[�!Ť�,][B�A�Ca�ݝ
l*k4�e*尉1e!�	�֒���&�,�o���gXc4J7�Wiu15�4@V��^�؅.Ф�YA��fF-���WT���T���:1s@3,*�Dp�xMq���%4h.-\Xh�v��uQ��F�ki3&�K]�˃k��r	,|(�%�n;Z5�vu6,Q]�������Z(m.b$��:��2�b��p���6۪["�vY��R��y�)\lj����mڈf��-�ctSn!	l0��8����]Z�Q(\MaAVj)�-����)�8��V��Łv�H��q׭�+)��b�0�օ�Q���Y��1��� R�`�8�4BN� in�v]��8e�r�jMvҔvM�N�r�Ҏ+�]0�:��35̅��t	k�[
"��,z�ĩ&3�eL]�.�t,�
ڃJ�asMMو�`���\���mո�����ڑQ�K�F��R�9���5ڧc$m6��ܥaI��V��qz�[]Ԥ� Et�4�Z�v���b[Ih̍Kr�E�]:Z\�͍�h�A��8�u-s)X�-��X��%i`��Vk]u&�1���b[0�T� ��԰�X���zi����[2���u ��3�ć9�W�f C#�l*��K3v�s�����Gr�l�[2�i���uSJ͘��X�G��Y2�����E����Q�!,a��m�3��U�#��B��-><�i���-!l��D��#rn������V,֘�L��[��p��eb�0tWu+��Қ`b�D2]���n�CZ�))��4��j38b5�&2�Yv�%�nƦ�D�l[a�Gf��1*R����Q�3��[v�i�T���XQD��5�i�Թ�VVๆ��X9\P�%4�i��kH�kIi���!4��H����˥ �ةHXLK��i�o k[ő)k�u�F�TؕD%�jl��ER�f�vM�[�C5P����6�l��v��m�Rm�5F+��`0������k�GQ�d��k�K�^6`�� pq	� B9�"�Q�
e%lI0��h�bb`��NW�4�H��PX�E$�D	&h-&H���h�rHMD��(�H���Z,� 1��س43h,"%!�D��4�&$�0�H�QPj ���!%D&��rH�;��*�DDl��H�A�C؈�#@X����i���h�PʍQc�4m�wt���`�62i$�%B%0�J \�c%��&**�Ad�ۊ� 0R*C�#J$����$�2�Xa�64I(�cF(Œ��`���Ǜ������"cnxL�Y���ΰ�Ф�%xoX��[ZE�]�ڎ�t��T�k�`F	�-��;qvcҮ�E�&t�����{	l	y-4�1v�)ٚ�Ѳ�0�٠ʌֺ���Wb���C6�Q���M�[]r�,�v&	7Y��`����A+G(u�B9-��9Υ��&ל�i�v��5\��
uzcZ�v��
�Gn��14&\JZ�Zd������UЁ]#X�q��2�M��f����1/2�=p���6��,���핱 � V3Y��X볮a5�h ɂ����`�a�c4t���i�f�a�]2��e�(:����`��cZ����ey�Q����4l#ټ�`��M�os�Y�=���3tZ�fJ)�3.4d�htաEbR:���h��v�lH�%�E5�ac�K�:�ju�f�%0̒�%�#f�hjC-��H[n���S<R�Dmi&4�b�l6�,\٘Kh���UnM�/bP�r]��T&���)��p�sr�Ų�i�)5�W��y% T|B�J²�إ�͂MR��E*J�K��5�����!���;ȱ���ŕv�/K��j�*@5���"b:0������6m���
i��u��������,D�`G8F�6<���K���CMI���t�0��m��͕�e�v�/e�¥�2�9,ң������
í�vc����u�[�:v��f����:�-X2�b��F�u#�iwUQr��j��5��И	J[,�����%չ�j�@G:U	K+2ǊX�]qX���M[��������#+e�(5�����G0�-jT5�Nt�YV�(m�a���Ͱ%R	tk�v����=2ӊL��u�AˣXƱ�*�R�6��rmg�6�t��ƥJ�FbƵ.�����Jbn�[�1%��i�4���k�D%d�"���b�kj��a�5W0����^�vh1֫$�Gn��6^)i��(C���JXղ+)h����N��KD����XX<��X�RbP
�a �Nmx!K�XK�įV0e��am--��X�Jެd�(�-� K����[hA����DK
�kV�F�
P���Ґ�0m���hM�0T�R�
����?b?�jk���e�G6�$�&����D��#�5�0+R�v�m}���+��A|[�������3U#�_�U@Ǉ�*Ӥ?Z^�q��� ��Ń�+L�H��W[�nB#s.�-������cU�y'��?�j�#�_IZ<<֏Y��ˏ�y�|��X'��"H��$_X/����Y�g�RxX~�L(���g+ ��H��!���uT����{��X=��H��ν�=t�{1ڮ`̴8��ZnaU����O��VA�DI�$VH�I<���2K�C<�/fu�j��$�}��ՐGIb���$B��5 `DՔ��Z�]\ô&�&�x��i��1En��)6\�A��V_��{("��ŃW�	^�_��<,_vS
->���gK����A�/���,X2R ��Y�;�eC{���7��9VYW���U�/��ۆ/2*�^��Q��L��S�%��8o���>�ZV�1I�a��[���S�n�6� ��X�u���N��*�X��@-�ř"�B�r����a����NVD�%���s�]�����fo�C�U��OW|A7��݋-� �[��������{~�k�:�͊������+���{��T;���~�:{�
��Y�W�2%��b�t��u�[�����.�F���i>�m�#�m��z�����9�( [j�?6�y���W�n_���'�5�M����7Vh�1�j��)v�i�\U�bH���PԕS�Β4�ݚ���������P�[έ���W�rz��;k��7W�T��X����� F����@�^6\=G]��4��d�dl��^�ga\7{���-rد���@�l�Kt�m}������ �+�۱e�D[�#]�Mzׯ�Fj^�e5v�6���|3v�Z����^,�������^R�WH��4oM,:�b�>�X����t�m�wiY����Q�9C��Z%�gٻ䠃,�,�e#b�VA��!���9�+��^���@A�A6%�mغ����}=�)׼�K���o���"�qh]YY�3��H��m��-�D7A�9L�תn�I�`o�Ӯ���opO_;5�\�/ܬ�t!��-��x��]	
uF�B��V��۲��.+�
�e[��ʴ���E�e�����m�5]T�#[�e�@�t��e`�]�ٻ�A�2���Y���8���\_=k�mCh ~-�`���~3T����#b/���Z�×�m)�r�{�������ز�V������N�辒� A���ma��0J9���}�nvA^�����\%���v ��h0[����|r�w��{�;u Τ%�B��؍J�>��%����r����'ay�_���� xf�Rع9�
���s7)$��`-�T"�yr;��\vϔk,A��o�) �AF�oMnJ[�h��^����p��AmX ����=�I{�KR�ߟ��ѬY-��׋�����>�Y�ψ v��n�?7W���n��ҳ�B�"J�F���R�)�3j��sj�r��p�j\�b�s-�XH"�yL�������tS�O��^�N�4n�T�o08dS�ʼ��f��m�mؿ�t�?�Ʈ�����x�@�_R����E��w<�0b�8�PDl��m��և�1 ���H����/�n�����9�g��ٯC<g���u��o�~��_ź@��-�6�œ�<����
�B�u�}6������*��L��4Z��/ܬ���SW�eb�cH�A|G>����/�m���K]?t.m�����O��s�p�e���@/� ����h_����3w7��nV��	���5��l�uw��Cu1J����*
s��̴sڬ?[����:{Q�4������g����<l!JJ�	��Z��XW7m�][W@Ҁ��@8��i5ŜV#�2��2�Z�K ���юl�P	��>YY�<vmLl4L�
i�!�]-���sKfc�a ��1�;�l�����U�Yc\m[�ٖ�F�` Y�3is-[X�q���l=�����R�LBW��/*֚%Ҵ.4"\�*��c�h� ������n.Ήf��¹�xOŖ���a-Jq,��i$Ŗ�ą̴0�L0�h��^ت�dvH��B���x�D6���݋�*�ʬ��z/j�눼��n.Zr�w�Ń% ~n�!�vźK��l��p�<��dO
�ZO��
U����r�z������;���ã��G�w�/��ma�_6��� ��l�
�\ڮ���zMwn�%3/��Aܠ�lAڰA���0����U��}<���� ����/�xVy�Y.��_�Gu�}H-� һ���S��}��;Ծ!���[�Y7>�܉���Q "��Y��ύ��S�5<tU��E`�����_۰�f���eJy�Ӑ)��j͒�бf��ծ�;e���3Y*�3���4�8��SmV>|�{���Ї9�@��/���]�۷�p�,�������S�߶�#z� �j�!�6��mY=�3y�He��W��N)�RWZ�|�J�i�:*�j{�m��;�z*n��z��KQf���l�h���U=�L��0��)�5�����8Ѧ�VZ�`}�=\��;�%�FwX��*���na�b���hX1�_[A�_7Cܴ�Ve������+��eO|�辽�"5��6�Yn�G)#�n^���d��"8��vR ��/�޾�U���v�.`Ŝ,�@K�~50��2E[A�@�[j��f�����o����g3Gɕm)�?a�Wb��G��χ�O�4j�tUn�_aD��n�S���!?c/3e��v��:V�	5etv4����-t��+k=_PAyA��m` ��^��n�W�׉�;*`˗�d�"r�<��{���nŖ��t�#�s;�g{�z�'ǲ����Z�¶��[��p�Fe����"�J��K6��;/0=��M���_[h/�m/�m�]���<�g�ǶU`H:9k�:N��i1��%fPB��b<��õԞ��Ͻ�ڵ�{���@���h��s̼�dQU�6hv%^�ٽ􊱫R���7Ծ#'/���|��`�P��zeW�g�E�+!�
�=�y����o��,%���Kws�]S/�����`[�� �݋�V;Մkŉ�,���I�_eU�ջ{K�3-2��C��ՃW�n�����#��,`��M��d�;ifʵ�Ic��#&�R�vh�P��K�s�������NA�_݋���y�ʌ�G�]�{�I���׺,*^�F�z� ��"v��Dxއ�⿈. ��zi��ޝ��<XK� ۋ�t~�#*�0��ur��Ջ镠��@���݋-� ��s�w�]_?O[����-����,���}`����mX ��!�	����^�d)[j A�W�mؿ�yxoD��|���w\ ���=�R��	W�����kס�%v[:�
��P��F[��6�<�v���V���A��xk��]g#b�fMO�Ɲ�JffPP�d0��-�e�\AhWA���`|�����3ń�|��5�D6���݃�������������
]o��� ��J�uQa��5`���q]�"n��R
��c��[�. 7����HKu�Z�j%��{{����;J�u��("y}����־m�V���Z�Z��}X������1{/c�������=����"&�[���G�OZ��7t��`_��"h"�V-���j�w�.�)����B��Y�:����h"��ͻ[��=����R��eO��r�r��H{޿3�Ca��:�&s�z������c�R6�xY��ޠ��-�d�@��ͫ:��X�Q��^ؿ�vyn�R�|����� ��DM�,��up�7۩���C����j�J k��`4=�f��U�Ӯ�foW�bO2��t5����@��y�Y�3��^����|�'�8������[�1n#A-\�M.v�o�ׁ%pR2�]�[\j�$�e�#��&�թ��͚��]��
SV6a��6��0ub�����f����ZsB�i���"�q;1�3)�$�s٘3*���ť��rhh�� 0٪8 �ij�Pk��R��E����e]���r2ҺY�:j!L��������֩4љ�O��y�\� ��-�k�õ�Al����@�錦�W.ŚQE
��q��矘q����#��[j�-���{�suh-ɽ�S�B]�]�Y?i���W���A_/�mذ[��n� �k3'UQ=H@{�|A��W�Wb�
w���+�4f_X'2���6 �m}�SD9~��}9�q�H��+�@����ݏX�/֞hWJ�Q�^��_Q��n��DM�/�[��H�݋A:c˪ �����k�m=�{�7V�̛�u<t%��VV�qĩa�H�b�ؗ����[��� �݋-�;�G�<k���Z��o��g�^��uJl��Y�PD� �m������j&�����<ߧ߶���3a���	�y`CH!%S�2�
k-�uEғ�kL��|�����O���O�m��fyջ:���N�����d����X.R� Cm���� f4�-�Ypʬ7�x�"��)�r��dv�{�Q�ş:���9�����\�8�$B���6 ���
:��'����^���S�bĽ^�Ӕ�;{r���]���m �쨳�j�^���"�_"� A��b�-�[�מ+�*wGf߇�	����ڃFe��>��ڰCt�6�g�ɼ�>�ϻ�*�����4Cmc��I�ug�t��A��W�+���>�����R �t�m��	n�����]zdTCyg��.�̞縦�����AA|[vQ�z�g.���Y���&cC6����R�[��A�G\\JB���TE�I+�/s+� JDwD,�H�[���_��)����ڃF,�����_�K����`�=��;��[A_ ~-�kӼ��3�����nł3�/��
����4s}����4�'�H�����+C���y0�7+�,�t�E����pvo쮺9����c��l���e:�7��a�`�d�ܺ�JԢ���;�(������C[ӣ��r]n*�WI�L�������#mꋲ�*�FuN��e3Ks�-���ja�Y��m<W1F,Ù҅X��Kй�� $��Ŵ"���݃�����	Qݐ��7���d�K%�yR�2T��W���j�����vY��q��0����I[�F�hi�۽����#�+��y�a?f��	��O0V�ƭ7Ca%��֣ݗf�Ovpr�1Lѱ�ѵ�����k�݅�(�j�����WEҐ8wMe�U�F]�Xƾ�ED=��c[�X��<B��K%K��&m�6����B|y�,�}�H�dF�:���qէ��8zy�"^���Njܴ̋vbw�V�̰'WOia��N�y@SP5�ky����mQsY{�N��Yf�^U��(��5$�h���h�hZ�x��8o8w�fM�~�tC��ӐMW�J��e�F�$s���W6S��N���n��N��/�Wj�WZ�5/.ü�w�:Zx��@us,�����B-����m�5��k�c�,�k���IB�ڵk�|VQ�
mR%����+U��R��~𡪴��iS��҅ez�P���x0������Ɏ�9mq�GdS��{-!l��Z$��Ua��͏�T�a�	��cq-C���r4�r_]ly�iI��k��N��B�Yz��x����t�<���JzCi��[ ����uzyv����	N�}وP�rݭ�rj�&5�G��ZJM!3&"�d̪(ŋ�4hԕ$hК�cb�d(H���(�ѩ�-(DɌh���T��6(Ѵ�Eb6B�I���6�R$�A�ѨŊ-h�Lj6���4��6�1�jM%�i51d��b#Ick&+!��#[D�����HD(�A�mE�h�[�ƴmѲj*(�Aj
��1�kDIF�I�,RF5�21|O�����n�c�����	��� Ƃ!�ʹ,�K�/6*ݧ���~���c���|ڷv:S����yp�}w8�+X�qnR'+v������ŪZ*f����"����&z��r 7h��^��g����Uu���a�&i�-t�n�W3F�Y�݌�)M���m�������NI2��'��"���9���r�j\��>z*I�H>��ȇ(����s��|(�J��=�=���h�T�T�u���}ݹ�H*A_T�{�ힹpı�x˿-�>'W�W�P&ﾐW�L�ͭ��}w��v�S�K�*@���uux��{�x�p�I�Q�/wx�����sS&a���� �*�ui+;��پAG�&�ﭠ����t���iC��Ru*��X�Mv���i�]y�*I�N�^�[���U��
J_���R��	w�
��&UI�����3������Sٜ:Sո�h�إ��V��w#s�k��t;J@&������v}�
���j����LZ�}Z�ء�v͞'g�
�I2�s���m�^O*��$�]��n�s�Sƫ��d�5��}��NHf����_����~�E��oY�Oм�u��ez�H|�$_H*A[���#�L�n;���~�l�]z�t:���w3r��'�{��#�TxUz
�d���T�;��׼�#�_P>�duc�m�ޑ�+�Z{>���IN���q��LO\�_���~�nB����S�]�Ȥb+���
aӽx�)
���R�L߃Gr��씍��b�T.�n0M��;�ǧ�������O�e`u�8c��m�)ٜ!��[H�.�FTڽL�B��&�	�Wcv�fZd.[�A�e1���t#Qz���-��XJKf�Z�Z�IpM�:ݤ�f ��ѫ5K�BSC8���� ������B�L�6�1-t.F�\���f+e�[�Ɔ�tb�-V %�nv9�W,�n8p���==e�W&@�Wc0��k�65��M���X}��<܋nb��(Y�c
� ���`Ậ�e5�P�_O��~��߿;��wo��R��ۧ��e��O<���g��<)�����I�r�ʊ���v�mW>�W����gC��]�_<�7i-��ަ*���v��v�u�|���썂����Wc�i쪜$I2�Aa�~��ϒY�>������>�te��_��}'��W�C��$T�Q;�_�#��u�1��-��x��_��Rag�O������5��.�RU3�\/
�l`��k�.��$��Z]�7V,�TQG�Ͽ����}�>�eT���2W��ފWb:й23���U���IRp��Z2��������SW���Tk-,Ch���t�������|���u1�z!���ua[���1�VY`�5�C�e��}�d��o
������v~^��C��W���%p��+J]B9�*�L��CU$���
��c;{}��Z�{�#��k�]��v��}��M��2�� ��\�+��W;}�<MpN!�Ev�:*Ƒ�k�R�$����ˑ�«yo���{b.��O;�w��A+�"F3%�Fd =�&.��+��eD��&Ĳ�M+ۘiHG�.4CCJ�t�����4ꦱ��ZhCL̑G�A2 ��ay���w����UM_����7���B'���/��U�0�B�z��M>�%#�@K ��
hC�2JhG#�s�9=q���A�ƌ� s�}��>�Ϲ���Zy��zP�4!��Hг ��}���[�G��{%Mۀ�І03 �!�̡� th@����?b�)?/�m8	l�ӏ}�,c�؃���!��5wu
 o嵯��yjf/f�C�,vɗ�� l�Yػ������c�͵�A�u~e�ﻱ��Ɵ w�!��h/�
Z�B,fJ
`�љ 4��#�Q��9�Ț�����[(\M��"Z�JXfd�6j�=Q>��v+��L�B��R4"��sf����M�	hCC� %�fd�BA�s%����A���!������� ����xn�c�w��N� &`>hC`o="�d-2����W���V���t3��쐑V	B�U�6G �K��d�e���-mv��`mڒ��e���NzZ���)���"��� HІ0̄��}ߙ�O�k���ݗ�y��Lٞ:��?y�JhC/%����P��#@fB ��B�Ў^���٘�SB܄%,;{(
>����^���ϳb�� 6`>�@)hF_� 3 
��ߢ��w�>yцT %0�d)�h/�)�̔����@� �\�E���s���L�m�a�{�ʝ<���������SB�%�f@�,̔&�̄
.y����a��aˆs�M�+M̹B(h[�SB�@O+���O�k������k$>bJ���q�Q��>!,�>E/l�î@�����X���V�}�����f%��dѪ�a��+ܸf���IB��xQ۾<��͝��<��
��#��s~�%M� H��І���B�hC̐D�2 ��{/�{O#���B!��Ҁܞs|s�>��>͎�y��B0+�
Z̿���� K@�!����~��������>b��@�ؔv[�i@�����Ά��G!�Җ��2��m�K�$����/N�h3�
Z�҄J`�2PS4љ \��1��c��~��������]T�T����g{ �Mv����@P4d�i�� �hD���'�����Eh��Ѐ6���s�^�߾6��ov��H|��4�g`�e�(D�Y�(7�RN���Ww�s��@�� ���	hC`g�(T4!���3 4!���@8>ٞ�՜���}��_���{6;��b/��-ϲP�M2 ��1�d $fHSB9lݽ��U�,hC�J,oe&m�\��3�̊����N�@L�|����B*���IQ�E��^�$hCa���)4d R�̀RЌ̔"��� naϽ�>�/�B!7�����������gv����hCh3�
F�0���`�2PP�,� ��W��Y�Gg�G�Q�v�6
������X%��X��t���U�N�˪2	*���ӝIʨ������*ݱ׵pf������>��O�q�`�1լ�5�DN��,���KW��a�\�X��2:��d�[��6B�ۚ��mC�/l�llv�j`�R��C,m�!it7dG��3A�j�fm�
�ͳB.�k�Ȣ�îJ�x��˂��DrW���h�8eQ(�,�� ^���b�r�reGYL�]���u2����k�+jJ���GM��Y/,lL��kcY�������;V�6l��EΔ�gHR4�X�mXD�֓Wl��:r2���n����{���hCߤ#B̀$hCC̔}Wߌ�����6;��b�}>�}?w��w��t�bhC=��M��3$(hCCA����{=�>���D��� 7`k�>_�+�p��]Ei�Lɡ���RhC/d#B̀>��g|��s��<�|�v�(
��
X�
F�fd��d-l3!��d�>�M��w�x�}�g3���H|І�oa _Єq0Y�"2d���<�%��ж�@�ԡq4!�nA�� ��6�(
ھ�fV��ϳc�� 6 >hCL
���&����\󾯛�!B�`	�B ���i�̀Ry��K���j������v���,ϭ��q�����֟ "`>�4��vP�4"�г 	hCe�/o��}�s�S�D�y�\S�
sf*1�c6�%�-ˣj��@�E+��M�8Y��tSX�|�؄
�} ���B(hY���a�	�9�_y���9|�������g}�U�/� �~�
�I�}(D�]����2 %�/ %�����CB=ol��*�H�_}���G��5�A^Tg�a�8�75{T}h��3 ��*��+fnu�ˮ&����Z����]��<˯F�
�_�/�O=����C~�?$	�? 
��l=�J��u��q������@l@|��6� �hC�}B2 |��'{�}�9�#�0���>��І�{Ѐ%fJ(`�2PP0C3 �ϹQu�N�繴���:����V� &`>��҅Me�$hY��c̔�-���c�ٓf� �@/}�RM
� KB�2�{�^׿?���6_�y!�hCh7�
Z���;���#�vP�4n� ̀�B���B��2A4,����1�w뚝�B)�����������e���� 6 >�� ���}HE4,�BR0̄.�Y������m�T�� �HݡJ�3[���.5\�vMH��jQ��v	X�f��i�I=�y�h9���_�����ALƌ� ��{���Ti�u;��f.��;?}�����\�} ����%��fH�̀�B�̀R�<�w���u��>��|�RhW�BR0��@I��:��~l�79�1�w$>����0�%�3%�v.���F��@�@^@KB`o�P�hC3$#B̀$hCa������s��L��ܟF%�ǩ�B5vӌ��W���ˊ�v�M�DN_iy��TP�B�}Y�},%uj�ɒ��Ӹvx��t2c��b�����! ��7Ǽ�G��2������B܄+��!4,�BR0̄�3%��ŝ�{+���m��"Fw%6�� ��ߞ}\����������BU��F��}��=��j�ƅ����o� 3 :Жd��0��B)�f@��;���b;��`ÿBJ��U�����ɽ����ܐ�bK; ���"F3%̀��������ߧ��F�6Q8���i^0�X���͋K+	�-��q+���t�����ӠI?y�SB>�@����3%A�v�7��o�oc7�����������hC^ܡ�@Ml3!,3$(hC�@������rޠVJ`�ў�	]��<��\����������hC��*��KB̀7{��Zc�ߟ�����@S@_�%�/d��fd�г 	Ml���3k;����^���u�S�\�)���i���)hG�D�Y�()�љ ���U�+������M�B�Ҁ>��l32PG��F�=��/��^��؀�� �| a<�w����Ԯ���ŷ�m��PԒ=��b{�W�H*�fn��mc��]��ց`e�A�b휢y'q�Qȗٌ���2.��$��B?4/ߠ	M��0̐���̀R4#2�,̔��ƻ��I51ǈ� 3��{g�Di�w⷏�L�c�҅Mw��3 � 6��	u/$	1(,�ݡߒ���$�(ZR\3X�,�ьZii�̧WCI��ݬ�X���� 9�lzKB/�JM2 �І&������Y�7�r/7�3�w$>hFfg#b�����}ۨ��p�Ї�J#w���!�Fd �l̔*M��>�}�����7K�օ�%#}������oy��k��������B ��� 3 �O����B<0ϡ# ��B���HЇ�(3%F���U]��ðI��/���
թ���SɁ[��$#B̀%4!��(
2F�w)��f�W���.u����Pн�BR�fBy�s�<o��?�#a��ܐ�4!�p
SB$��N<7�j �vPb`�4o� fB���� /! f@���>g���';(
�������s������&�1��@)��� 3 �B�2d����7����ӆ�#'��MwQ��Yj����W�υ�X����7o/_���u�u����1��wG�� ���e�O0Ń��{4E�_$��[���g9s�\d��I��<殟1[���f�V6ީ5��飕�lG�hb�7^[vj��c��U���`v�ZCr�yG����g޲�YRв�{���	��Vf�^��Ϯ拟H�6��ٍ���+s�ڵf풢�@��KU'GK��3��4��G�ap��ћ�j�*�=�q�٩�U
�nB$[aX�ږ�2��Y�=�|�vu��`JR��f��-�T�J.���MѼĂK`zrUa4r���)�e�Ga��-�l����+S��ɸ�Rۆ�ne� �Z/��q�j+[cv�.���^
��`�\�	jʊ��jTTs�w:�F:��k�n������!>3�&#����RK���	<���\�nn]V|:)k6�}[����cs��R�+��w������6��:t��r��f��1m崃O,�:�E��pU�,j�H� ���6��i�����aM�u�׹����%[H$��I=Y�o�Y�����4Q��]��U)�(���X�,���e���,m�}�2�ǲVV�49��ӕc�=\��pD��)s��E�4KM���sv���Xȳ�n����@ۏ4�ku�Y͵����G\��,�F����]x����c��e�(��K:�wT�]>U���OZ	�z|OoR:h��5�FU����Z|���&��{ch���c�o)�Y����p�-�vfB��m���֍�X�%*�Fɓ�4lm�2�E�I�̍�QIlcc#��b,H���@cF���Q6M�b�(�bJ(�F5&*�#Q�h���1�X��cQ&�6,�`���(�1��"̲j5�hJ��ڍ�F��6�`����UAQ��� TIQ`�6(ѤƢ�XJ�F+I�2Y��w��|�C]��Cdo)K�Yrc Gi
A���-C�X0�ؤ2�XҸ�%phM�ku�+)`����$[o����up�Sc��c)��k�.���ar0Յ�a�k	Ya
�6�A�V��1n%9F�WXCb�6�խhJ�F]��1��Ьat��3��ju�e�ʺ6���X�[H�0��"C k��ii)��f���Y��L����.m���֒�l0k�j��T�e�����*YA�MTȐ�6�Y.25��"�J�s�у�`��m�����,ե�KLV,���5���1	i��Z��F�-��f�ʸ.��xb��t�ˢ���t����vM��&rXp�٪#Q���f�ճXf��[͢�H��A��P�[h�-�`.�A�& (�l`�3b�;t�&5(��\Q����¹� i��D�f�����4��p8���ե��vv��!�n%��,eh4��!��\XB�v71�J���u�4�r6���5��4GD\�1�l�c.#4he����.mE�hD���(�	w44 Vĕ)�{U�Z��;R��,�i��x'���'�@�.�n2�Ζ3f�T�*��o��[+a�[y���Z�h.v�v�,��A-�;+�N�f�h���M-Ku�i��d�ۥQlm�sHA3-����Z�kff	\�-��QԵ��k�����%��a*�k��r�݃0KK�`�[E��֚��׌����k0laY@!0�E`n	����g�*�,��[�K4uXQ%�-{mD�m�S02���h�f��BS%6R3�K�њ��u�mK^��X� �=�7$))/ZJ�\�ke�/�S��fDn��u.��v4+շY�L@��l͑{r�
&�Л7fXh!�� k����m�],]D�Ya������Pq�YSldfw -��V�w[wa���rf1�K�����T�Vj�h��#�xY[	Aie�ۮo�%!E�f���+���*�.�VJԙ�˂��R�ˬ ��Ӥ�������)u�3�����^��2����K-:mUk��)HD�o]Qv�j&�"�#y�%���:a��.�d�h���s����@c�Kz]t�V���1�4�Y� ��k�Җ�	J43�r9�lz�c�
.b,u�Y�80�xX묁+�R��f�W���Ѷ�c�KB��2�\�)BX �5ںh�7
��5An~��~�"O��С�HZCMc1#��ۡ��h˄����Pt��C�RC�R�\� І���K����@� {�}��:�8Ӟ��6��	���rw�y�\�U��hЇ� ��� KB̑yք1�� ��w>w_a�>�!h^�Z��	�>�M���ב���r�>bK.KB>�B$`�2P]Y��ڿ���M���hCݔ*�$)�fB��(
�Կ��QY�d{����lv����B��! e�(GF�� Jhd %�fd�4!�_be�뇝�Pw! i��#��AC6�� �}߲o�\�s�]F��3�B��zP��ψ�˙��;[3��
�JF�(
h�	hC`^@)hC��B(hY�q�w2�bL'a<�����~��6��\��B�e�)�҄K�����Y�޷ﱕ^���L:uR:��c�Q�5[%�51��8�;B�WEil�hF3l.1ـ�4!�3�(T{�@����3%P}^F���ϳc�� 6!�}���W��s>{ �4!���I�_��̄� ��@��� =��2����15��YO�|5��Ԉp�u[��>63<�o��D�i�;�IoB�ɐ�v!��o.��̈�b�ZV��~~��]�]�R��	 ���|5s�~�¿�����fq�����:����m��%��b��T�$Ry��kxsR��^����%��>�*�T�{���r��jU�!�I�7�C�4�ps����ӡ�C=^�w	�B�D�E_T�������Q�:k8WM�c�q��~^���ye9!�&m*G�d��_��ϲ!�YK�F�b;RP�J�mY�(U�p�[0��6�I15QT����Ǟ�v�H]»�]ۘ%T�X�2�*���w�Y���]/(|G�ە �}RL�����VM��d2j�33��6���,ه�����7z��{v��^;ImzE�]���.�"���V�x	�w�KC�����	N�8oG���E�JC1���ü�{���6�C�ݡkӓFV^���2'6wܩ�͎?N�q�o'�bI"��8s�NUH>$�:�;���e�U���V�y�=܄t7kỨn�۹71��\�%kT#秞����[�)@>���V`��g/Ŀ��W�fT��K4��X%
��WA��a2]�+2�a�@���
�eH)|1��/O,�g���]���'T�a��I$���=9��lt|>�>$����K�bw�>ܠ2V���3�l��r��U�_y�7wln�4of�؏zq}�kr�[���«_���Jƶ�KD/{ԁ��*d_���IgV"�R�W �!�DK%�c����%�ui��5�0�'+/��U�W^��W��������ĬV=[�fi�:�ӯ��褿sU����sQ9����	! s=�.�Iw�L�I��
>hC��Zq.���P�>����/�F+�E_H쓪�_;�7�@����6��h8����F�3�f��j�x]cn%s�
N��gۢARL��9��}7|{rNw�(�J�����Tg����I$UR#o�S��n!%���X)�$9:5\N�I��� �3�������)T��J��љ���ejQb�,@��}�R��R	؝f߷+uM~�W�*�[�wW�ߚ��ٚ�\w�0�
VXNK-݁����"��} �d6nl��Tm/f^�a�	�Q.)�k�[͡�[��6�g����vc�X��/b�\䆋�=�l��J�qԺ�v^#��0��x7�&d������Μ�B@o�����wt�H����QҲ�m�R�j�R��-ɦf�Z:L�s��Y��-,�l�-^ڮl�k�����piu� ,�2˥kv��EL��!fE�\���4֫���Bg#)\��
��-ݮ���{ކ)V�l���l�6�T+H�F���d�M�[�%sĬ��T�F1�5�au�1���Ua�=\m0�r�	�ٮ�2�T ds6�\Y\!�Q�B������K������:	�غ4bu͹�1���JH�Y@Pٴ�.���I��w��Cv�ݥj��mu/��W�����W�NwE �T�+'�O3к����{�mTo��{�{���n��9�~���R��I2�K.`�_��"��^�&'WԚ&���ݡ��n�>�}�VsY��{��=�:n�ڷmu/��L�3��
���s�2:��*h�H�Y��lQ����7�{^{�����Orx��!�[�;��o6��!��U��L�.u��!�i4���mA��Л@�f[��L�(�#*��
�)ɒ{�bGw���3Q+���]�8���C����v�&���`�,:2����G��۫o�ʛ��4V81�xl�^G�ץ<�c�kV[�K�����Ż�>�7�k�9�Q����`������ށ^�55܌k�1W��6����>�ۡ������u����ỻcwI�;�a+���vo�y.��z���(��ݯ���B������ �N!�tʐR=�bg�յ*�-D�qIz�{!n�սC���n�ۺ��iT<o�T}� j��E�+h5���g'��|$�U!�N�K(�p������)��sf��ͦv42��Es[���-�hԬ��RV���|}�۳BΓ}�8����o�N�5��϶��*�i����k�[�w���[�3;�c7x�}�H*L>��o����A_I2A�;�5}H���|wK�����4�T�j�DE�.�Mf<	����V��6w���FEm]OI����Q����{L��c����V���C��O�t|�H�A&-��eX�j�X��P}@n�>��٣�n>����=�@yP9����� �eT��$���I�D��݁�9����Y7�n/�h��V�H����0Է�\V����6�@.��!Pfu�50 M�� �&�m�}�v��R8tuv���W��rxy0LL+���oT��������z-٭��W�>�v�֗�M����7������+0�#����H>�eI�"	�'���ӻ�Sj���-Q�Z�6�hn��}6侴����U�� 7��
��pn��B�c�F�{��Z�L������T*����+9���܅���_6�F��c��cRҵH�ܵ��Py<o3o���2H��=�qD��q�nf�> Gs�\���I��I���b���T���^ts�'����7� ���S� ��<a���4H�qkl�G�KaL�mB6U)���3Y��	�xp�=�t}�>�H���v2�����g�R\�w,���}��~��H>���A�(�:���:��!+�� E��
�r>���-��T�=XE|�U?L�� �" WXC�<.E�甝��o+��ʐH*I�ef�S1�nJ��sW�v�N4��y�喨�}�ֆ{o�i����쯾oPݡ�_�Cu"���yKn���
���[���k���ը}O�I3�<��֍י�� O��lѽ�_��˱XŊ�h��ls
����v���L�;ۺ�{�]�#�����]���諭� ���a��b����ׇ�Ke�� �1m����Q�q]mi�JƉ�e��]��XkSj�Z3WhL�X3M`��h��m`��e%�]�l��d����F^tBh�e��,�Ԑ�/R ̗g!-Eݚ6ŹKU3EM�.L�P-(]�ae�LPՕk��f0�Y�]��mҭ��K�˭�5S��������۪R\�/إ�
d��\"L�%�����jf8���$��*�D��&ZG�l9ؤ�9�����yƯl�{��ݞ�R	&} ��2)�����6����w�\���F�൯�m�9P�uN~�������P��7h�e�"������hY�r�=���T�+�$�Îzl��y���>�e�w�C���=0oR�}�x;F5~?b�*�;����H/EK߆�;��"�u�Uu�k@n�ݯ��������ߞ��)wh����%��`9d�h�0�n�"B�,9n�`` ��Na���T���􂰟+����{x 2z���'8.T\qH۴������{�k|m�����T��}�,�ky'���iO��k%6�#�/�e2�5�fC2 ��kӡ�]�NSҳ�����>��n}.�ϻ��P�'���^�P��vT�IR1�ñk���m��v�������G�0�w��\t�#�P�|�pUI$V�>���ឃ1���v�V��A��0���U%��s��Z���`Q��dyU:C��*�V�㎒�]tm���K��OoR�-��yn�۽J���w�HQR���c��.f	�������m��Y�g712Z��vV\2�NL����+!�v_��y�͖ݫIUN]���� ��^T�K<
�>�s��=Pk�L-�9UT�����I=,cz��[xg�zeT��I K�B��ek���k�Yj��XSOy/@��S����%7@�]�1�72�[��.�x �2��Gv����iD�(.��.��en�c)�7F��)�����F�NṗXӏua�u��	Xf�Rg�^c+-[4����f8S�v�V�e�$u�r���)-���l�#��j�m����Nu�B�_|n�F��%cd�4���O>��yƇ�Hn[h�����T��u����#afy�7�G�t���6Da����ɭv���wF�WB���5db�%y�[y�g�"��ڭ&Q��+ǧשW���y�yT�ğ>��]����5�40���]�ǋ�h��9��eif!R�~t��"W���P��*υ�gL593�4��E3�q"�mn6;���uw�FhD
�i��Z�-:����vR<�̺���s���`��g$Q$�Ec��ػ+Y��������c�U�z,��-�46�,�Ze�����~ݺ��i���VfX�WS�AA�vrZ�ۺ���z�Ҥ8Ns%���a1S
�ɍ�G���ۑ�k*�gVwk*���t��B�A��z�.����5p$��w/T��J�66���QQ3	S�Ʃ���`6���:y�N����������W���GlX�(ɸ�;I��$y���\q�9���k�tݤ�w��Ae���gtw��o��k4�������a�!t;k�!�:ޥ����˫�FY����pǽR�$����p��IW5s2��\��+�zJpOj\Z
`6�b�H�b�4h�Ү;��6�Z�X��c�+b4F�sQ��r�lj5QDF���5+�������ۈPX��k�ѱ��r��X-���kr�lnsr��],U�˛��G.\����W+I��S��v�Lj�m�[F��N�lZ�r�IE[�X�f�!�?�����7���˿sa�Y?S�g�	I2�	�ױcXX�WA��ݯ�������c�F��gV��Ϳ?����U{ے	$�Lڋq=���o���x��5�� �꣢�M��yvwJ�Ǐ�6�	%b�$*��%Ԏ9�F��XV���0bD�]z��*1�eմkM�럾Ͻ$Ϭ����|S�\ޥ�Ok�mG�ʇ�}[�&��$���Q�U��[��=
G�L�]8�O��~�p�w>�I�Ҍ _VϺfS�[��&H>��e��K�yF���wNmc^� ������W��@��ޏb.Wp�I2�Ku�0���4��}B%2��s��{xL�m��5)�f�(�S�����&��/h�>+��2�Y�"V�jr]��ī|N��f&�K��ɹq��os�oo�u�	 �ݣޅ싻���݌O�,�UU��q�>�:�k�W\m}���Jl��r����,��_*��͍���BF�l�],��T�V[Z�VV[�[���2��ht#kv��]����=�UU-�8_��Y\3~�q�n����[�}V�M�*�Z����7����B��>�{���f�f�	|�ޭ���7_>h��u1�Y<T𧕚�k�W\��8*AU$ʓ�5��8I��,�`�'����ܶ�� ���]��jQ���ܧ�¤$�Hf�.�V��{R�T��8��\WNiᾯ��@n�Vڴye���PAϺ�����p21ͺi�����c[��9hx��x�a��v�y5N����_KU�ﾓ�}[v�y@\r1�������-�!I���ms�8�l��dՎ�٠ʚ"a�XE�)t�, ��Wf�m�L���54�,m�k�5�:��A��6��6��l(FD�t#���@��̶����fG���X3f ,t
&�U�W!i����8yoY�qu �Z��eXC�v&0�̪�j���mX6*˻ܖ6���>�o������jں���5��bș%<����Si
����Ѭ�
Ç0O��)�}$�}��L�#��N8��k���G�|*I�H*�h�Y<T���j|n��s�UZ}�	!�c����0���q�w�U �}Q�7n����;]�����s����OTB��T��ARL���׻�WA;s�<m�c��{�,�』V�ʂ�3�W���}E�I��I2Hgg;�^�� %{���k�����D>�$���_}�|����x��)6Minם��hs�d��[3�m�Ŗbb�,�a�Ywf�ɢI�ߺ<�IYZ��PvG�4�������H�}:�ݭ�@n��u�\.:�\*֦<�	��a���6�b��1f�@O)*��M�t5��/z^���S'W��Gl���p����7���%[��>��}�&�q�w˶Z��H�kv��^I��g����}$�IL7	�&�{�#Z�,^���t�)��O���������Z�ޥ�KwhM��4*�������V׼�{�Wp�eH*A$����S|��?veL�7�#����{��쪒C$��?7�����cM�˫�F���&��]�:���:�A�� �)F���%
��4n]����^��n�ݠ����u���Q��Ҍb����I�
�T�1�U37�{�5�s�/�����8�p�87��P�3A�7�������w����I$�e��R��Pm+{(V�r�����wu�Ǿ�g�%�J��:��~��/qBws���(�{}�AM��������W˳�=<�靖G읔��A��$���}Æe��QV�ǣ���������(�[�3�������U�k��C`�g� �xB��i>x�Sܒ�R�y�p�9�����7}��{ϭ�0�8)�g�j��*�*	��2��8���lMZ��5	�8��8�M7RO��o ܋�����~�M���u[]���|���db�>�2�EI2�A���iu����R{���'R�v�P�~��}M
���|���]��>�s���"��o�͠���@ɵ�[0��=_l����ww}��n��(>�A����{j��m�U��q�
4Bw�J����c�/˖�T�)��Z�et��V����_Z�jԗ���{Tu�Y�A+����4�������@�🾪�����{�T�I"�~ٯ?
����I�=\V�=�,~���A�I$��u��M�f����F����*�R�d��Ĭ6�v١Ɓ@5s��f���\VSϽ7�jސ�3�W�?j�s��d�~�xvݷ�xpS3�wӵd�7ww��ҪiK��{��^�u=+O��i�6�m�]�Q��m۬��{��n	oU�F�렁6�_źD5��]�J�R��Ո�6�����8�s�T���`��̪L̒Sn����5�*Ebt�%��fE����v�%�ڡ��_��űq;��_/� �6��-� ��D6�j��[�!���x�Zv��NsЍ�^����n�m��V�jy����(��ի��R[x�[����
Ws�E�4�2�P/}�o8ȣ��ג©�A=ӥrq����&�̟N�FO�I�}���m�zW:�-dr��=VDc���L]�ݜD�Gh���f�tUnSKM��Vb6�K�R�Z�],��aXJ�٪�[��Mj��8��%�#h��bC	��m.�����lذ�c��jZU(a.�mr馫j�Rfӌ�3vK�4�/ZͰWW9���)�՗J�m(�Z�%���&BB�&:�����=l��i]1T�W��+G@_����F�[t�^%q�	��N�mXPhU�k�Ͷ��V�q^��,/����4 �f�'�z��\�B�<s�pK���IF�'�aUg�C��5q8O��� �����h"� A �Ց��Y��S~*�N����qX�ʙ����j26���%�Y�<����3��
[�S�$�m���X�ZJV��%?.Ҡ��w��֬�ź@�[j�m����?ya׵UCA�޿�V[A�ÜL�{�뮒�X^}��ܤEv?=�[FQ��_���t�%���ڬ��tM� �)r�_+�2a��-�����]����X�[�?6����_��C����z��Ud�6�)�C���g�&u�5�b�V���f�솮]t|��=�H������Ѓժ���g�iPyz��Ⱥ��7�g-�����H��VFd�� ���F��c�n9��ʯ!r�J�	e�{�>�e�^�7V����\�f��?G%V}���e{)�^�Y��|La,�:г+r�UU}o~�c�A��A_�~A=�����X^}`��@�t�V}�廛�-�`w ���A=�X ��@�H�mI�C��Ot�͚�݆\�Ck�'=A|A���H���+������N��eڮ ���/�A}��W���o�iP{�]�־�m�9��a�HNȾn�� �Cn���ӡc {S��๷�J5acC�;�� 6�!�b�?6���$jX�ݿad;�TQF��B�TE�i��E��.�L&飠���9vn�A�X��������GJ� A��W�{�(���D�����z����%����H[Aۿ��t�!��>��p�f���_�w �[�;�5��j������W� ��[���J���i3�z )ڿ�":�AnŖ�[B��0P�5�l<@�&e\�h�$�=����Q�ɪ�흪vZ��Cv*�r֬�g��9��V������z˼4��9��}����LV�y��]%����N�"�����͠�t�"Vo�	ii�c���:�@�_"�V>��dG�x�)[Ck��"Ø={끺�޿k�r����m�-� ��@����iwpiɌ��[�㕒�"7яV	�\�z� ��`~־n��m�~{v��h|�aU�٠��M3�x� �"��ͅ�а:Œ�c��ڒ6,Q�f�x���#dB�n� �����¤��K��V4$��wnY�{��R��"N����-��ڲ0?<s'�uo`�^�?or����D|�a�"�hew�s� �/��nR�e�	\�{�%s�H3�tR܉��33%Q�[�po�~,��,V�uY���ob�ƴ��@6��eX���q���.m�%}�6��\*Ay=��X^k��p#�F��޿q�B��/g�{���k��Kaߍ:kb�[F��gwvA�klV&�4�]�j�����Z�.ȯ��汖k2���~���ԙ�J̎c�ɡ�2I�kǛJ��¯Q˖���y���q:\���q��K�͡�t#�e�گ|(9 ����cg��&Z��[5���2�0����KrQROM�iCyؑ�7d33�"���W�G
�ޣ�z�GWP�M�dk�����_7��n����Uݷ���*�����A�A_���E�G�cH�y�(n��32IC33{�r��@�k6��_A{�o���P ��
Aը뱾���Lr�"�b�t���_�A���s	����+>�馏׻��z�KR�]�G ˺�A���G��wF{J::���{�432IY�JcY�E̂�8<ٮ�D��r�:�⇏�k��1�bA�2IffU&�$�v��rL���v�/8k3չ�(W$��fޗY��bĕdKj��]�2Z�e�9�:7۾���ʘ0�~m÷�[m;�ʺU�M��x���c��e�9Nk/s�d�N)��6�\Ah�y�%�mqB�I�ù󧗥��CWCN�ㅎ�:��βu�e2s{i���{j��<wX 
���1h����9�N�ޑm�3��������p_,�R��l�4`��il~!M��Ò �c�6�/#�q��ь��3/�����#X}�����Vu;�ݮ��ɧ�u2��G߈���}����h�Ay�ӊy�����ȟd��"�].�$�vc�/�v��	��F��t���\�+B�,��F�/�e쮣O���gp�wR 4c��N�ק\��^oY�iu__]�Y���e���(�hǗ�.�a�.�sD僻�k��Nx�v7$�!���Tm�Z��̛.�	ڼ�t�d��0eLt��]僷$R]���[���N
T�6k{X��v�˻��Afp��m3���}|iq���Jȸ�2��u*v���oqG�X�zW8iKѳ�b����F�y��������o�Ύ�ؖ����\��ٕ��y��e��ے���}J��u��)Zj()d�7��@������hro�`�e���G!�I�}x�^�cH�Yj��U��ާd�:��
w�Ր(�鬭��7a�rܺ�q�Ь2�U�79].6�*jʚ'b�U�`66��6�V-Dh�\Ź9�Uwur�6��4\��' �s��;����h�[��p����湷-;��ŝ�����n[G5˛Q���wu�u����F]��2\�\�tI),[�k���.k.�-�k�ӕķ9���N⹤�[��鍹�E�r���;�9r��ۗ+���Rs��F�r�8봘���QN�w]st��V�s���r�F�-r�+.��5�5[�sQW9s�r�ط7����fb���v����!suB�u��<ib�127Q��jQ�x���&��ge S`+6ZȦ����l%um�P��u#�b%�
8[��YmhT�3-�̤r�(ن��y�EmL!��F�u 5�0X�aFn�6��&���Mr��֥�r+(bc���y��]�M��(�V4���7b�ԣ�����Uv���f˄0B�u-Rf���lt
�fʺ��uص�[��{<��#[-��%y)��Ka�K�1���:ba��f�]H6�Mv-���{"U�-p�K7�tQ	�c�i�#����A5y��cF�i��\dæ��^���A5�L����I-��б�ĮshH�iz�\K�{;@��ծ�8��k��a�5 m�v��V�m��a��H�%��K��V�LCZ,���6U�X`)0�4���.�.��*Jٍ�\ebؼ�ɦ�tM(Մ�+1#��
+��qB77�.���C�c��!����2�2�[�vbnSY����%p;7U�`��t����@�-�E(�-HK��c������� ��#�k�%-a�Xٷ0V�Un�-���R�e��b�f-1eY.�2�a"kYEZ6Wh	�[�.�5hj��t-�԰�[R9Sl(ai(�˃M�fx��1�U�HS���v�P����I�f9�+�U��-��JinJ�ĽVb�l#̷���-��Jeh\��J�ZE���:ƩLDu�5"=F��E�.�c01��H��]E��0�4vD�Ќm��s`Q���Sd�-��jR�Y�I���U��)�9�L�B�^.�杒b�-�-��	��`�b�1qM�1�M9D����Ɗ�%�K�@�sZ�)�ʲ��;;�1�ݵL��D�6jY��%6�B��.��U�Ҧ�װj�e 2��Tm���k)�\J��ǝ����Tk`SJkKuŘmv�6�h8:ذ
](�,2^����#�ы� gc1�p�k-����I��^X���� ������c�����eݝ�5��.��1��8����5؅"4 d Wmhf��w=����%n9r�+6�R\�� �*7LaS�����L,o:�v���-l��wk��II5�m���e4lG;.��������7�q4�Tv�\���m��`c�t����ꖔ�-(�KLaBaU7Z�m�6�ۆ�
�S������i����rc[	wc�A�L)�˸�V�PY[��4V��,�}}:X\_7^?6��e_�����W�W�\�<�"Ub;�e���[��r�M��m݂[��P.�+_{�+1zg�����8{n���k��Σ�b��7��������7r�O�P�&��ԁe �w�u��V������2�����Z/�/�r��9Y��,k2Ifd�Y�H�"F>w�3�I�|��mm��e^emz�=Y��)e]�+*��O5��_B�vWF���	n���A��NEl����U=��mIi[�V<�/��G�'}��#Z�HAzҪi��M~���\`cx.�6��t���1[i�����r��5���[��y>�$�?|�By��*�Bצ�_���`��}ow=�v�W��C�_���E�@�u�g��1�U���^q�_��{2>q؍o[�1�}�A�z��X�E,"9�0kY�T���.Y5����O[E"�ww�P��*�h�y���R ���0[�:�=Y�л)^��e�we�t]��s՞�c�����=)[@6�����p�Gj�()�Q�vy�5�_��[j��3��z�/�eP�F���!��v�p�Ay�d�u��K�+.��W����zǫ�ւ�C��mX!�|[���fy��1}G`)�Υ�=�e!�ʺ��	%�-��6����k��_]`ԕ���ĩ�n1E8���=���n6MrB��KpǓF��]]�C� �O���"wA=��36�.���;w\����3NC�wr���-� �ڰm ~-�_��&�ny����f���xZ�a�/��{�d���@�A�j�ƺ�:��R�=HA��d�E�@�����!����[[yU�+�����.�Q�m������ܫ���gX��g�i��R���o��5�c�p�//4[�w6�[y��ӯpb�3G�<]z!����l�,�K�mCn�������V"4��j��H�!�b�-��n����+��Σ0��}���[�yꙩS������8�H�t�۱`�Zl�Y��w-�<BtS�J=|=0�eH�x��DA|Cm|���ͼ�>�<C�+6E+��Avٳ:�UA���#"3a�V�D��%�eeu~�����YH�-� ��V�*�N�>���z!��!Q�I�U|�(	��ز� -�y7H2�^它�#zX��Ƀ³t%�Og
�Z�����Aւ-�-r�^���.�}Ά|vP	�b�n� ����m�����^��
�X �D��_Ŵn��k�wu��-E��;)~-�b�*�O�5Vt�ȆW	�P@��v�,`�[}�ҝ��Æ�e�vB�enr@j$o1��D�f�����M]�Fl��U+w��H��ivh��ژO��:�{�*��� Cnłt�-��m��W�w}ş�j}��;�S�{8T����y}kA|[� �҂]�kвt�0��Z4����4���X���Ll�b9�	r]iJ٘ʪݮ��6�� ��b�t� ����F\�z�؂·����zp���ވo>���$y�)�̚�u���=�H�^��ʼ��?dG:mdC+��\�e��z��T��w�2�d�!�o/�C�a������^��љL-]w�{��:����-��e_��y*��$�,��-������&.��b��K�@�ObꭕY�O���)5y$��R�2hc�$y�rJ!/޺.#����o��6�!����P@F�b�n���φ��'+��"R�H=���r�%�Uz��9E+�vne�V1�FԢ����CH[�iW�Y{���Qu#v=��Vf�F
M�X&��o���.���Z�߾=��P����˥u,,0)5`�hj���@�ܗ�Q!�,n�F��v���Hh�;i�TΖ���q	U��]pM�.��-��m,o��؅&B3�-����)	wms2AL�kMաԔ��N&8�)�[*���Y���^�r���ìcse� L��--�6v��6�Gh�1����P�006D��Hl|�}����Ytr�j���9չ9��4�����i1�JJ�ABŠ�5��3)C�o/��;=��|O,�7�L.��]6���f_���5��)�D��ɠe��t^C;�U�p"���:�9)|A�W���.���+}`��_7@6���|/}����#W� ������l������^�@��W��cEƩ]���$��Čeܒ˹���lh��\�����������i������SW_p7����i��n^��������_7� An�@6��돬��<�wr!�AW�"=}.ܬb

��D����m�>��?M���PEshlî�L�0����0Aԅ���U�q���5f��%R���`C�-��ں̬��� 옱��� �����k� �z�2ffUdJf���Gh�CJ\�4_��߷s4L2aڼ���U�:��N�j�[��� ����,�|���‭8��ͭj]�`]�՘E5{p�/|~��r�󎄊�-`�����?^��ƴn��>F�>gwΐߏ��P�m�e�@��Ə�ټ�U���#���s������ F�۱�h [��	I����]ur�j�A-�b���;�L99�b��E�;���~�� ͤA����?�|AmmХ>��T�T�n���=C����؆�\A���A�@�H�mN{Y\�����~��K~�+�{�nv��D:�e�k��.��M����`]�sZd���,�'�e��}����u�r\71�(z�X�m�J��4��pc�I)�{E'�$�2-�`��WՋjy^"�|{k�{�>���pS1�5lA� �� �/��L��f�/}��A Cͻ��!���?_۹Sė�)��c�[Y�nm�m��z�&��՛�c�2�YN�"�FfX��a��͜��w:e6l�()�cn�Z�n���o�.�o4���K�X����A��`����H~-�d6��r���<�g���B�~�����ṌAC���/)������d�/��H��m� ��-�����ň<W�fVy���kg���e���X��t���9�}�huW��!v�4Z�L�`˷+����Q+sa���ҷEn��ް��.!?y�'�x��+*�|��|@.�z�!���^z���b�ZA/��Am��ϐ%��m�Ho��i��������x_w@��b
��	yK�A�D6�s�d'����g=�y*�8ƞ{�C3 ��
^����a���@�������� ��7XA��]�,`�jͷ���VU����tV&��Sʈ�]8E�ۺ�A7�Xs�n�W�z�����c�n�$�/��M�U�M����k;��K�o=Ug��,��,�]:-:#嫇f��K��U���җ�qa�'�p�+{~�� �wZ�Cu��6�ۢ��h-�Q�9Y��W���lz�{PP��^R!��w�Y�b��~{�c��uZM��MV`Mnq˪8�J��#0��T�G�$���qC�"b�ˏ&1�nU/l�<Ȓ-�a{+<v	yX�t�ف�|�yc�*��G����n�!�v-����a�{�ʧ�^��xRo�$���sk��S����j�Aւ-Ҿë,����d{mY�}��m���HChRb
�,�������9ѓ�^�P���e|��y��[_7_y�6/��#7��ng$���] �U~��0K9�_3Y0:�&�s<C�I�N�ù_'���-���A|Cl7��f���C^���Y��������M������ A-��U�A��3��UV+�=���趚jyܞ��6-UiOT�c���g.����S��|�ꭌ���F�:�b���hRP��B�ҵ�ڗVpY�,��V*^eQfĺr��BSD	W3.��֌-�Q�ڳ)0��V6�@"Ijf\�sx�
�hbgk�ɥ�M�!x�GR�3Q��Tt�M���uPVuX[f�bj��i�Eŭ8vi�&m�ڣbYA���d&��7\�b��"eB ڣ�d�����D�)K[��X�l3�J�A��X��ͅ#X!��Ͼ~���v2���Qf-t�!��\$�IY��[M��(���V*��i�9�F���F2��)<�S�$�{�3����kX��4W7]L�Ѣ�*{rHͽ��Fd��!JfM3���<g�[�u[>t��r�^�����5�� �6�/�q���Uc"H�TA'��㲐 ������A����s��t��ϛ����y�S��?^r�Aւ��HAm�!��d�l�~o<{�[�gR �����,g{լA�~}��fR#i�Y�n��'s�[+��R܅���ɡ�̕��u�k�X�.�:�Vl�j�T8t�`�H~m�ΓͿUC@�|��vJF%` ]�6�f!1
���pA�Q��k���j�ٰ�5p̤A �m�����V����9��U׹r~��ؼ���,��ڂz�ڲH[������x��O/qj#-�4~1L��7�x��풬��0V��w�&v�-���n���U�WU�^�!���Azu�N�Յe7�{JD���a�'\,g{ՌA�~}`�2�_kA��\:�ʽ�
u���@�;9X!��"Ŷ���d����{��d��JhuC�6��-� ���j;����}Ҵ�!����w����F=�*z����W��Ű��_e\x�wq#�zi��Jy�JcY�E'��1M�>7�E��u�';���	�X ̯�ւ!�w����nݱ��,/��lW4tVK�GFc4�ņ�	Z`,�ȡK�a(�f�e������{��/�KmW�/i�,��Q�\��Ҭ�T!�yl��D6���|E�_;���.�G{�_���^�n��a1�i��O�\�ڬ־n�����
]�>�ՠ��{� Cm�@�@��xxN�1G�ջ�[4��b�=eaK]n�X�0u9�w{MiՉ���m���<���Vl�K��h���\&6ow:ƞ�]bhE�ю�	Ɏ�Ym�г+�=�.Q�=f=�eL��:۷�F�nP�V�C7�����]n�W�K�쫑�I�iD�q���i���Qt)��\qn����1��EK�:A�s�*�5s��eo,��L�%����7(�����W�F�Լ�MǹCO7�\.�ک�EOVԑ�)K���6��թ�dz��a�s�fZ��D駸���]"�
	{	���5R��i,�Tb��ĺ�c����i�{��y���%p� ���'f���M��m?��9��fv��pi�D.�WN�,�mzV��'K��Ȉ\�ԣh�� ���Zs��3�u�coi'�ͣ��pCpq����򺯠�2��S9�;`��Vi��� ۩�u�׆��D����Mڻ�k]��x���f楁@������xyB��<>�҉���z�40g�;����{M	K>���²�`��Tcr�c��tu���;���NfSS���qٯ(��)?y�0״M&W��1�9�t�Ƭ��q|��+�,�������ljs�q�{2m�B����mq%a����qg+�f��3�c�E0�l��@ԗX���|��N񵇸�b����4h����|M7�ߙŋjmE�s�����77�!�(�ܙ����U��h�	��к㩔�Ԁ��\9�=�Z��ޞ/ջ�ʋ�\�܍rܲ\�\��A	�X�Ո�飲��.k��N㛷v��������sn�v�˘�*�+��w];�wN�E���娸��\�)��U�(��݊M�.��A��5�l�%Ŋ:[t���.F�j.�ѱ\�拖�;�tű�7wG-�c\�\���n���Ƌ&��Kq�&�G:�L���F6��s��];9�*9�ȑ�h�PS��#;��XљN�`�����\��s@&f3��srî�(�,�ƌ�.sM"�*9�α%��s	�4�I��sc7D9\���6�9����bb�^Rk�����k���T��ѹD� �� ڿ��^i�X9}�%Q�\>@�{A��Y��ۮ�Z�:��|�|D���~-� ��!�U���~��b�O��Q�QN������j#�_������n���Vk�p��$��`�Һ�hF�5�U�V(V���f��E�m�eՊ0+������Eʬ�S���!tY�J�4ﴝ{�{ؘ���p�)����cp�}~� ��_��@�H�m���G�`���lW����%���Ij�\�7��ؿ�t����
�Ye��H@mm���6�����3�b���N����ğ���{ڬ�5��tm`!���n����/yP���J�A���Ý���]�bb��D{�U�x��I����+�̫[Cf�}=�w��&ܭ�'<F�~�^�e��յ���y��I9\֐��o�̃�G����w5���}_��-�[j��n��oğik�<mj�-z%��I�p\c*��P@��,�Hm��^�����Մ�>^�KtȻk4����BkcaF&"�)�f�E��@pJ�Ջ�h_G`��� ƀm���=�{u�=�S�1�R~���W)��]�Ⱦ}_x���@��C���c����W���Ds�����rl}~��ΰK�@�������U��5�^�:��u�`����|�m�>���V�.�vQ������\'ޠ�"H�n���"wb7��z��n:�g�����Om�i�2�i����M��!��c��i�H�Ȭ�@��"m�7�!Zͱ�(`�U�;��jg�y�����^R ��6���J���&Ӿ^��	r�Q�C*�-��/+���.�J�m_B��b��`����|\v���VLR�p.o��}�'��F�_�%�>�����q�;�C�Eݚ��ci�¹�M7kQ��	�F�ݭ�ؔ�t����SdrpgL��B��bY��-�&ʛ�Qn5������k��H\ZU׳1`����F[R��1�T�9���Y���m�`8�,�q�.B�ҍ3�;M/�&H�����.wL�I���r��� �b%�bٔUƌ���\�%����+%C:�!xƱ��Q��ڱ��En��_�ϯ��?��Լi]te����q0��gS��ص�iX2ҫ���~ɪ�E�u�~m��.�%Fu��<�����c)܃�x�m1F���,� A��!�b��DqW4e���l4�gu�+����h�_(C�u>�&���sܯ��n�v�=s�d���� Aޠmز� A��=�q�rؚ�,����K�ɍ�L�����D6����A|[�D���+���n�Oe�|2 ���ڰ+{��:����F.�}~����Ԓ������:@�$Aۻ�|Ct!�:��X�_j7���Ne-�,����oit���'=���A�/�͵��qqk���t�+t�VY��3,�&)0h]u�S]�GfŌ�bR.*�����>�������MwGۢ���^:Z'����3<kĚ�=ڽ�g=ȱ��$�}���+28�����N��ffa������t���To)v/j͂Ǐ��t�F��;�p[�vV���(��q�;����ᆬu���~6�*�ז���6�{�7w@��z8�|�sV+�=����p�0���>�*�h��#�m��uv ��gh���%�����6���沈�+����z�	�'�\~�r�Aւ-� ����k/��Į�؞�Y�Pd}��ua�����U�n+�m8N��`���x(�[��S���/���� t��_Xm|�T�X��^�(�
��Q�{�H2�
� A�� A%�-�!�%-�e�H�
���I]ZDT��KB\髰�)D؆uG'jt6��
!Jmt�����P_ۻ����b��ו)��Ryu�K*zz�-�> ��}HKm_�7A�/�ʵ�G%��=�C�H� �0�:����}�N�߻���1��$ffWc�{�z��ia+�����~m|�x�j!�9�}��3�ʫXj7�<���L�M��t������ܾ>��oy�܊O��ϑC�5<.�����Q��R�r�# ʌ*��� �����#�3 33�w����F�e�}�z ����A^X�o�{�S���U���A=��C�{����A�w��_0q�Ch/��� ��Yn�]�������8+<�9��E�o��V����]]V�o/�BtBn�(��w{�C�	S7J
�`��mb�P�k�ڑ�Q��.�,.���E��U�X����_[� t� ��V+�=��*�v�TaW!�P�s��Y;A�A��{����	n�#�a���>VG�nuX4�"=�w��B�7�{�)�so*�]p ���`~ւ��V�\X���E���P����:CnŖ���hN������;�&���W�k$C�<P���C3:�<�$y��}�.o�����A�|~m���uEI\ʐeFp@��PDP��5n�^eݵ���<`)�mQ�������=�NϤ� �GP���h��W��ۧC��DR�^��ډ��[�<֭��)U;Ԁ ��!�b�-���]!"�_��ǿ_��4~��+�����V�П���sܬ�!+��&�a�����Ϟ���eсD�+.�Ye����+4c���������ѷM���_F�l�'��/�d��?H�gܮ���{�r@t?{�1KG�3N�倃9���H��+��X#!~���sy���N�W�e{��xj�eFoX �P@��X�$L�����/�DI�Y����Q�?^�R ���ޏ+�Ҍ������ғ��N���F���)��ȒX��f>3��R�R����ދH2 ������~��{NH��u����
Ry��6�vK�������$�������� �sGz��4:�Q� ʌ*�����P_�!`��dB����f������@�{Z�͍�����4NT �wq{�q`�"s\��3@.ZA�\�NЬ�Zf��΄j�)��uW��������a�ap��,��]�3C�Uͼ��+��(�˓�Tۚ���lX:$�LmJͱ6�Qͻ�Xu��:�[�[pKV0t���!����W<�tY{b3'R���)����Σ�K��-*B��v#�5�bBх%��sX �.5����R탚C���̢B)M(�nҊ�\�gf؁mQJ��"\VQ���̷ItfUw��о����eu,K�
UטuI�E�0��˲#JcP�+0i����ɻ����%D���$��{o}r�Ra��\>#.�45ݍ��8��r�	�+I�%Cׇ�nm�;���?�y|��}��sL{�w��9 :-���C�"H��`��Z�X[��:�	���$�X2R �"�C�+r�{���u܎��1~T4��%�sh��vh����ԉ���	%�Fm����,X��o;�\���2�ˮ?o�Y��أU١��@����$�`�%2K�8��w��������1������~��W�PI$�Ҩޡʮ�V�n�i�ɩ��/h�ՠ0֗!n�w5m�ȍ�4h�J����Ku��d/n�P{ޥ�Lo����^����x��X�*��	=� �m>�_�w+ Ȃ"Iv	�+#m��_��������q���L�j�:�R&,�T�z�N~�T��ZYc�|-�J{��%gZ�"�W3�c���ﮖ�~���F�4S���u�siL��~����,�X�{6Rs�m#���VC�B�u"Ib��+ ɔ21�O;}΢����GW�������$��Rf��ݎ������j� ��>�$V{*�\o�����0�pr�>7o�)TP#���9}���$�I�~�D������+�u�>�yb��b��^���A�S}�����!`�H�d��,J�D��f�n2ئuڹ�e�n݂��#p.�g-�X�+]��+4)Y��B�~�/�"��!��>7f��=�~C2��Q���}�	&_�I,Y���d��#2��
�w}��D�;�B`�h�Y��4rS;k<���@(�2E�.�c
�H�Zw�Dve���X Ȁ�e�d��W��rǵ���1��V�h�u���,�byѻ�8����;�]�2�o� 9r��u�ڈ�I��m����v��Ż$��[�QnV)���{���,X2R���+I.���Z���<�^�[T0~�e�.r��A��86=�w{������V�v1عzG�7��h0F���������D�2V}v�*�,H��wG���ͥ�iq뎝O{Tayw�;� �/�"�dC�Vy�������C�X�Ø�,l�(R%���j�@�[T%`�k�%*�~O���������K��!창��ڞ�7+�{D��_
��Ľ�ac�����X"Iv	������VoRHC���A�3;NٳU��{ :<���g/���$a	�.b^���~���`?or��Kd�$��8{�{�[�t�-�:��Q�^��P�0$V"D"I`X"�V���F6��3�Dl�%����g5�{��N,Sq���������f�~5��ܤ���4}:	5	Ar��K��[�>�;�*+H�1�}9��s:�t�����(����񘳥���ʭrW�謉%�&JH�$B���O �{���횕���ϞE{�M	�6I���������r{q�?�����e6X�wƸ-����iL`��S*���7�����7y�o�J_2Eu��_w��ʙ�Q�^�+ܨ���`F��h#z!g_+�A$�`�"���OQOVne��~�9��۩�6"���P"��nX�%[�O>q�}ج��PD%�H�%��aU��Z`��z�������L�VA���>�����d���j�ͭi����A�#�Ծ?I��U�.w������U�	�@cg�=��G��>�__r�%�&H��( �#���k~_Z�,zsٽ�S�l	���W|&���Cq�)L�0����{����>�����{0��T�M�e�s����wvS7B@�D�U��Y`v)(f.�z��%�b�ȃkv��4CŹčfc7z
���V8����<�ČR��9.�|Z��Z{2��{�[uU�Ƶn��'�b�xE��^.���b�/c�V�:5G�AN���w]�����',�]F��Bn�)�i#rFE�<ti;��$ޑ��ه0�{���Ý�{�h�oOfͶ����o7mN
�gv�d��֞���ۦ� ����Z�G���h�Z�M��z,�t�su�Cb���GO��c�c2�z?�J�v=�G�k�˕k��5Rb�$*�D��Y'm�k�e��m�e�3��
�Cwt�%gÚ�^ w+�A��f_ϕr�oI�>:('Z�gi]l�;���f:βF��Tx'���ز���x^�^�����q� x��W�o���K�`��홺�&�+7�iz��Ү�?^�ݖF�!���7c}yOo1^���H�Ҋ����фP�ף��el㨡+3���˱�N�H�G]|�G{�f��)���]|Nr�j�hnj�;n���]{S������*;ي=��3Br�~�-x/�V�Hn�j���^S��&W`�bY�3�W��?�b��.�ơzqڗZ�ڴ"ɹ�[�����{�-����䦉wSX��Zҡ��^��_��Vv��S�!$�ܝ�B�y[�DA���-�_H�>�B��MGI�s�'�<���L��J־S ���Y��ꬠ0]f6��-V�)�7�l͊�p�_��t�Ngy�ˋ��1��B!�dBP)�]
�-��1ww8s��d�.���k�4D��wh��]1I�9��iΦh#��wt�:�ܱ���ݶ�FB"�]۴�b+���E�����9LƘf)��s�dѮna�˗$�QLɊ!��7wf����D��D�Q��wV�T��݁`��Q�w�.v���wgw(�������)L
�K��IP�.])�Ц�%�[(`�T���d�f����wRQE!r���S3��.�f�%&!�B�nW&X�$�a���hHdh�L��wu�R"#�\)��"�b��%$����H�0�����|�Vf2�ɶQQ��h�mq��m�n���@�i�U�f�Z��n#+��6A�;J��j�p�1WZ�J`��(��oX�#�ؖ&��53�Klz��!�Y2I��B���u��X����e�u6iX�9�4��SiX+�ޏ\�ͦB���k�gF�����6��������^�49i�	�X���3v�\����h٣,ٍD����[U�(�̨1�l,����P7b6���˖���7g,Ƣ-6��ᚻbQf�kŠ:=����@���e�Z,]]!6Tm��e*L�F0�ƃ�1�1�0�̚�"9�՚#�b۶�0	��.��fjZ� ���Ƭ nl*+K���ذֲ]���c�S���0p�Fm��(��Wh�lf��)�(���2���-v�K��bs�m��-.K�6���j-�pi�[�v���`6U,�.Fլ�$c@����reKi`RYa���64�R]�i[����[5sn�%(\��5��jF6% �B�e��1��{d����xa7kzc��*�إ�
��*����K�Qҫ0K��:k(Yto[@�;7F�z��� ̦+6��.�5�4�v`b#�ۮ�����$1��MI��I��Ț]bC�
f\��d�&�٩���D��d� ěe��iu����A�95ݓhR�'emr�s����M*^X鱋���d(�\0H2��A�ueЀ`s5�������JW ���1�"�f�u��C[nUV�1�xl֡�z˚���|Y�c����uq�5���VA*�\-XV�7�$l��lk*]f�ɗ��و&h��kT���.�lIe�DU���L���Z��p�5��꫸a�Y��\���f�l��0�[LXGX�Q��B����j�QҚ���d�6�n��u����1cYf��,�&e"�D�&��)-Hf:�eJK��0l��7\�(�8��#�M��!�4�d͹뒭��A�b�W���-.�6h��0�E�jF�����&8ڙѳ0�)6�gh�:�u�6�V�E��v��y�՚��U�Y�	
��A-�S��V���,ڵrBE����(	!T4�qQv��J�k�1�����)`6�\�aV�Rʜ�)S[�k�\�-�؅�T0;��*�M+R$VJ���|BWe#C3-eұ�M�n�c�C��m�P�9w\.���fuԬXf-�Z�	kY�.��M�HZ%"oD���>��;���- Ȃ�v��f����@|=��c���N+e{-��k.If�Ҥ�wh��1�wf�������w,ub�O�� ����U�.w���SsTayw����rŃ$I�9g�s_�v�s<8��X%�VA ��]�D�ǖ�)��ݐ�ž�n�xH-�D�u�{�� ��fJ_A�+G.��A�TVex����ze� ��� �gi��6m-�d���;�3��B�F�[�L��Sb7n�!�b��� �$VAIIYRJ��R��G#�櫮����$���U�;�2��H�dB�ŝ<�x��Bg��ݐ5lj��]�`n,p��1v��8�JXmJƵZ�\8t{�0?��$;�t���W����H4��y��,��Q�ǎ�U�>�u�X�T ��,)|A2E$�W}²��K�L�}����/m;�Ү�i�M�r�:��k�8-�4���x�{��{v=wx��� ��g=�7V���/o�=�ʌp/b��33�O�l�[�����`��V?8��wv8ppDŚ�7�˪���Ħ�6h��$�`)|AH���Q.k7�����{�I���1u�L��rř"���"H�H{�{kw8�����`���_��Ż���s^p�] �.!�7:��u�x�D�VD����Kd���`����;(n�{Ƴ����������`�("$�8����9�C��r���"�Y��i��W����Me�F��s[u���6.������r���% A2E`W��as�{�57uF.��Ʃ�l�Zf�����=2ł�+"I�X&H�Ja��P�Za5!�������K��w{k��B|��~��~�r�nX�%p��{��3`G:���,X?��X�$_IB�B��7�>��z����G������R��v[F��ۅ�7��w�>�r̥�t�0�<	 $���������]%�Dmȷ��`3��]�2>���n��X&g+9A$�/�$�����P�<O�{�{�,Ծ?I��S�;:���ΒgJ!x��|�e]fÛ��~I���(A�@�"�H�dA$���<�����=F�dOL�x�D.��G��_�}a�b���d���.r�~��͎J9���v��0\u��!]3��.�	l�]([��B�*ͅ��X'��s�X2Dn����~J�^��gu[�׍KMh�]��=�^t��#{��$�fJD\���;��AU3��v����ײ�e9׽�v���,fPD��,����)OT���T7�0�X1�A $�/�$�:�_,#ͫ���I��u��~4�!�u�@7���ܱfJ@�d��"Ibƿ;)݉tf!�8��$�������d~���n�^?s���,�=�]�����*��B��<���
;^�}����R��,˴���m
Ѵ���*n��T�Z3j��xx�m*Ow�P�bS�vhc7v��`�����=�*U�0М=�gx�1�&��`���rř"��2 瞲��M���\>��Ch��MJ����3B�&���%��V�*�J[u2��M1�JJ�>C����� �9D���K��e�1��2xҙ*m�Դ�>>�~�n/�7�,ΤA2E`�"��U����``��`��!���5��o8c���X&g/�8�"H<n�%������K��>_I�d���$PvPk9W1�Y�v�ﺝ�{�`��`�fPk�,"��/�Kv��"��m�䮑}��Dt�I�+��ѽ��xԼ�m�N���E�Q棼�o;�5��e"	��Ȓ]�d��Ib̑-�d=K�P�|�]�3o��U�d�b�!���qD�}rK	�,vE����a�vb���@G��v��҉����_���Ŕ���6��;���T���ګyճr�6���ԾA�b��MZJ�&ѪI�M�ct�6)3�L&�`Wf�(A�f�bY������T�ȱ�;5GA����h�	���k���ֹE3x�^D���`\eK�٩t��F^q���c-55��������9�Ք#�.&�ԛR�	��@�%&%Ib�C��i�7�N�)3M��f]XS��d8�6[��L����ْ�͈WJa¦�D��}�=�Q���)�f�g���f�5p�.Y�-[�Mڗ��Q�Y��HB��B>�,�H��X�g(�v+�.�7�`��,�,r�s�j��z�3��w-��wiP��٤��|�G�����L^g���x�Y��=�S���Џ]]\\����J���K��w �~�dH��J}$�`��D��גr�;��>�:����=�"�@�:��+ ��A$��d�,);G��i����teE|�|A��`Ծ �d��9L�دawq�S׸X ̠���w^����F��"�%�"�A�$��)a��U��IR�-�#]�*���n���+���H���mx�mg����K���0a�m�t���r��P��l�\&e�ټ�� ]Y���h���2���A��;�}$P�(/e��f�#7=�"�@�p8n)�X�X��5~|�#_]�$B�����3_U���K��Ӗ&k��eR�)v$*�!��u٣�x��t�t�W��;�G.z��'�x%ֺ��hve�Yd�pSW��7wod��z��Ǻ+���;�������>�U{��4j���VŽ�3;�C@"������P�$�/���V��IڵL&�e�W��v��W.�Lhu~��ݢ��H�=ݚf��%L�~_���T��b�r+��$B����G�=�E�L�ڬZn�y�{�8<݋��������A�ѫ� ��,��Q���l��ϷP3`٢��_�h"�,Y�+ �����t�!�w(� �j��iQ��,fe3n�ҹEE�vu�6L\Jҙ��g׿>�]�VD�E��%��^e�1�隆U���u��|�{�%�λ�6�O�"{��d��"�?a'<F�0g����Š��^!�}��.g�H�P)���}�� ��"H�l�m�A��n�Y�K�.Ed$�fJD��o�N�ҽYbY�=�5�Ջ#m�2V���g�{�x)�-.�7��2s�k�Ǳ)���\��!�YZ�Lm�c}3磳�\�ϱH�w~rV_��{�d�~]`�^�@�ܿ��@ Ȃ��%�	��t�<�[q���F�I�$�/���|�ڵyw �.�{뫫/�j뫐]��OЉ�nl�ξ@��K	��%�H��^��^����A���.gb����p�K謂�$�I��I����h�h�X�i(�E�A�\<�i6P)F��G6�D�ً��J�kr>������~ ��`�H��]{9��՗��^��/˅�+f���!r�C�ŏ�tV?H�I.�2E@7a��=�-]T���M�Å�J�r��#�U��g�_��[��҈]�8*kߟZ�G�݂\����d��"D;՛���.�뱘\�p��ʒ���u��}�C�E��,Y��#�=h��#1ز�����g=�N���b�`��~]������~�h�W+��Y6I<7�]��u|�x_H(e���Eo���N�3}AG�Z���q%��gxW���X��Y��7���֭Yi��}۫��D"Ib����"$��a���}��=J���<�v9��z5]��r�rX���2E����ߵh窭V*DհX:���4�NͶa���Mf�3݉t��6��U����[���F�X�d�Ȓ�|ו@�>���t<3���Xq0�=�\�C�5���4s�$B�2R��d��?[&�ݘ��7&���$V+���gV_�1���h�\/��H�׶�rꞕB���Cy_��D�"Iw�X�d�>�ռ����'�������A��b̔�"��_�8g�j�Lc�@vα`�������U5ԗy��:�?Q���ϻ���c����b���"�H����׎��B�>3b>�{���Ҳx��/(��H��A�	�R��k,���K�ܸX;:�Ѷ����c��|^��\���/NjwsC�U4�V2��XR�Cvhzka�ׯ|�Ԥkv����u���)n�3EΎ��m*5f��m"J���P-M�[U#K��G��*�\����]`�uM���Dw
�vDt��U-��)c4�m�k���D���u�1�(/R���Lʍ��en�Xq�46s�[p��&�J�^B��K\L�I�!)\4 S[a˕���#�1J�K�1l���X��mAqa�l#f��9�KfF:b�G` Y���L�a q�h�MpG}�xB�J{I6kIB��[0���a-&�sst��F�҂%R���U:8lL�ܟk}$�7v�3wM�Iׯ�u�_+�o���'��u�x��ز� ~�+��%�(/�o�VS޽��m���ՐD��^����ӎM����A}���DJ�?}�<�{O/�Iw�L|�@�X����"����;!z��du�����G�p�AyAo�X2E��L�7�{����Zψ#9���IbǕ�6W�y��d���p ��VE�y�;h�9�|�Z~n+I/��AD�Ń$UϽM�[�ЛC*v+�}�CQ@����VD�E��,N�p�z̽���=��ڸ�4���m�b���MYF0]���maXu�� ��\j.�2�}��7>y���{����s�������S�h�]���k��N�/��+ ��I��2E`�75纯�W�iR�K����ѠS«(�B�J:�� �s�he*Շ\NZ�:r���9g��=Mh�R�֠�0IFV���]��W��EaNjͯk��A�{e:�A7�VA�X�%k�ܧ����vg�_�=���%�2EdC-����-���1��E{�	}��?8��g���2W�н�*\���N���_�V|AH��9�Ε�Y㡎WҔ���^���w,ɞ�����SU�~�D���A�/����!��r���c�l_ܽ�oɉ�w�9����o9X �,Y�� �$T{އ�q��3��e��LM��AMa.e�PҊ3�r`�7]�X�)���U�Y	��i|'.��C��Y�+IAu�j�rx���bPV�T�+�(�3�4ւ|�k���?I/�+��~���#����>���}>2r>�L�3����4{W}`�}�k�W�آM�y�~
��fV}u=�A<�X Ȃ��%��H���U]�si��7�hy���,t��C�sw�e=��HgJ�B��)��jF��y��Y�8V��	m6z��O�h��+q��n��k&B_�3A��!m�hǂ'�(!
�4�L��O.��x�I��Up;�X*��dm��0�)��׀�_b��땇��,�90��9B��p��'���3C�:i��k:�9BS�}�`є4��6��8�̳t�S�T��
�=�a��mǻ�0�7�{�&��nmhl"��AO���N��0�t_j�K"�c��]�ݳJ��n�	-s+x;�aIՂ)k�Cik�Q�1���fUyy�y^TX&��80Âefn�7Fז��t�)9E�V��BU������<��N��}��9�$][XDu3o�����ݕy�,���ݾC�+y-���Q���]8�=���Κp,�ohv���sE�j�a���өp��[jU��#ף��`�v��ZK�Z�+��
��W>� Ǫ�/r����x�u�eK����t$*�NZ��!��1�Qg�m�Q��h�o�{x)Qc
�l�k�`�N�x�+P��^^��~��qP���֍ʃ�wt4�� �6��5�*:��q��gf�f⾰�,��߅Ys��x�'�]l[�d7X}cߜK�uRA.��r9�q���ٓ(䫱�_^ʽ� N��n���4z���Eg-�|�ʶ��|���m��D�ʾ�v{�|��t�ekK^��aʼ�WQ�if��v���7��μ-�V�Hge���k��y�s�R2fQB&F �wiݮ#L��D#�����.n��f$$��F��rI��s�A��de�'wL.n]�A���!s��9tF��DR1w\d�v�]�+�)S2As�1�.�@��"���I�4�wnI#�% ��Z�������Q��v܌�� �wj���I�)v�J"�wJ�� � �������K;�ѓ
"��P�I�Ț ��ЄA2�d4ِ��Q�A��&BT(�N��'.��))!�D�i 6wpdD\�ą9q�.rf�w\�c&�A�	�O�{�s�CǱ�sv\�r�A�X�% ~�/��t��3����fu�NV2 ���՞+�<`�z���ً�"��R(\�3\Yr�^��Ov%�{�43wd��xp_�Mr�����W]�C�'�*�r����]`�m���$V����>�nT�	�g��Yp0�U1f���� lS*�����Ze��L��]nt��a!��!�`D���"��cu�;s�f�.��!�xP�=i{޲�aw;��"�H��d��������8�}tA�n��ۂw��A[�,�U�\A$}b���(����y�?wr��/�%/� �^#�m������+�ʖf�j�`�m �����AP@$�є&��w;MB�'`���X���c6��O�����׼����CX�W�ۣ����T,��%�9�u��vjP�]a�	�Zx����Q������l]=���'	���Uk'�գ��S�c�~n+"Ib�2PD0"�L���K�����k<O�xAk�D��޿��d_$�I�~:(�����)[��V����HGHY��q,h�3[���t�R�ݢJF�"��J��or��b�w!��_/��X��L���)t''��z�X����0��G�_�w/�H���"�+"K���=�����_�9^�;��y>N��v�A��d$�+�+ʇZ>3�a��`�Ib�.P@����/�vR���i9Q�A�z�w��z�%�V. �K���Ń%"�u�Int�FQ����njgR �d��T9�n���^L3�����!{� ���d�`�$A$��$V2 $��CkN�k�}���r��k'�O�`n=�k��XG��������EeT�=c�G�sn���:�����$�A�=2�:�'�Y���T�ֳ����wk�8r���"Fx�U��H�kDPcg��A��Q"�EYW���\.�2�4�0�j�i��� [UК�Ym�)(�--1u�:A@�%��,�g	c.C�E��D-푬��k���ƘĶ�m�D�6?}��I���B�(ˠF1Ԥ�h��ZF2�n�n�1d)*ֲ�Pژ��ҺݭTh�W��1��]��%�+k�X��6�	`��hX�[�7\������:u��q$mݜ�t!���ub�1�fTu��&4~��O�AnX���}r ���ܿ
�y��ȩ�[�ĭ��=cfS��>��1��nX�Ib̔�$VE��j�����_/�NV+�P�ҷ:��k&��x:���`���<�V�5�	��X'z/��DI�$��������ד�~it����;_p7����`+��2E��E�un�R�s��Хm�s�_u��o�Lx�W�"�+w�^E`�mOR����n<�q2R���+ �,_�J*[5�zaWF�8~�+��)���>w���5ukh :�ř"��	��~]�o�]o����O�z}0$r�L6ܺ�K����Qbt6*km�Қ	!�(�tV5��vi�����ݪD	%��{��ʺ^����|Exs�:���x_�6r�r� �"�$�`�%E�F�KN�ގ�^Ed.Y�75��,���]��;{ׅ��;�巶a��a�t��������XWy�yDb*�q{��0T��o*w2�W�r��ru��o�^<���q+w���y�P�D��}���[4�A�m A���d����|d��Vj��!��6��>���U�d�X-oX?:F��fH���$@�yE]�zEcA�]�@�X��w�N���{{;_w����]c�p�np��m"3�X"Ib�J�K�uQ���W ����,��WY��0V�X%�V!�"Ib��!]�c>����]��[�,���hP���]"���80�)�&K���k�R�-�4��b�?��!��V!�b��� �d����d�ns��=�L�J��ח^�{_���G������$A$_I�7;���"!HϾ���%���'[�J}��nl;\A �yYG,X2S����l5��G7��;E�� �$�fH���ז�쨹;~�fQ	<6�7�j�M���s+)�b���.��͢r�y�/rR�q
��Y�~9��y9;���}3��m�7(�G+�9�_,���y8�����VA ��X���X����4gxEq�i�P��g����]��u��;.�������΂"��;�Lx�r�� w �K	�+"J${���� ����.����O�m͇k�'���IIX~�-�r��vk`�V��[p�˗rMu��s�k.M�D��u�4J��J�=��CO{����[�6�H�-�ۋnz��F
�C���ৗ���d7w��n�=ؖ�vhg4��7��ͼ�<f� �[��W�����+��Qg�墲����������9E����Y2Hͻ���Ҩ7d�3wh�͒�Wuu���C��{����z�M���>�_X�X����$�Vs��A�7��� A��Y��A �-�-�?z��Anu�\�`���g��F9!��[�;7_J�7H��绋�2ѻ:�u�L=x_*��ww0��]�U���el�^V�$�4:V�j�e��ny{<8�Gw���2R �"��,)!�����Ϗ�ފ�{Z���̾Ҹdy^���k�d�Ȓ�Ъ���������#A?4}B�Ю��":�3�%hl�*�0�h��S��s.�pQ��jJͺw{41�������\������~��k�6��c�k>�|�oV� ��>���d��E��0�������s���o'��.[�[S5�Pru��5YD��L���݋=)����,Y��?IR���Γ���,���ه���`��__�E�IA$�,_�oGXǧ˵�}���ǒ���7yͺ�1�W�|�YJ�;��-_ky��|�|�EdI.�J�$�_�H��3[��u���޼�.���.n���u�\�`��I��뻍F�B^�<�G�ܱ��Aj�|���n��t�����UPOx�M��wy��m�.�_Q�h��W��y��7$ˈ�c���n/'����K�f�%3���$�IRZci�geSA���]&T����I�d��H���X���er���ͅ���c	���6��[�a�7@�R:V�r�.�&\j���fR��Б�-f�,��ce�(mX��j�*̏,��f4�ь,	i��jl�Q�V"���
��ڌ�bS0Ҷ�f-5D4Sv̈́b:�Jl����C�8ut���}�سЎ.�,�n�)���;h[u�l�R�]4 �P�Q�iQVm̯����� N�\�A���4�2Ϲ��Y�u*-ep�l J�2Ń�+"I���/�r�)��Z�`lۿ��%�$/;�~I�7����ظ$�Y���4��W��dW�]����$�,��AD�
}W��κ�¼��u�\�`��	&_�Ib̔���vd0�` ��lY�H����gz��L������X ����l�twJ�[��f�>��"Iv2ED�	&=ݬk��{����wa��Fi��w^ɏj�����d%�2W��tf�_��[�_��+4���6�Y���h�n90�(�+i1x^��6h�f�$-�	k��~����i	C�{�ژ�R��)�.l��)�q�^�I#3ުL��(Ov%1�ݓ�]��g������߳T�^�+'�kh�eg7�@_�����V��d|hax���B��eO�-��k�zn�UV^�]m��V�1�r�?l��3�vz{ޜ�A�y���y@!��Y�%�y쮡�^��c��Dg�1���E��%�&��2s����GN�cwY��Ty��=4��v�{�#{�4�����f�q�uu��ǽ��q�b���d__^�����^S���
y�	sU�^��o��GgX����Y��FH�C�ŏ��9e������vO]����Y���`�{��K��A��,"�A��������6�.���$4)gJ��j�E0P���$��gk.д��J^c�y���}br�$���D�ŏz����N���Y��Up#�����y݃{�L�X�c��n�!�b�n��ٻ��w���a��d܅�YZ������栂��&� Ȁ�+Or�_�u�;���|�d�,+��WUz��^��י[I���6�*P��5�I��#M�n�ǹָ��Z�M�L�����1�R���݊PQ�<Cd����e���݋ox�gS'�\�b�t��Q���+*�}b�r+"J$�b��y�����yr���u��Ib�y�ۯy;ǽ�fz=U�O�+!֑\;�O]�I`��H����"�"H��$Sɋ�MP��~���y����|�V�}`�\�`��"$�/�$������:J���O{�ݢ��&�֘j�#�M`Gks)� �T��h�/m�X�[�Ͽ�>y��=�����]|���w�7�0^{�<��T}�
� �m� ��dA$B�2Dn�?\����o?r�Jv��vQE���<���g�����+ �$�fJ}i�FA!v����d7�,:��!�H�~��+Ӟ�:!K�����]wj"��͹���%3wj�[�Kv=1�ɒ׫ܒ���,�R����/�����,�\�z=�����l�f�X�MzTL�e4RS:И�5�Ɛ�Tl�RWV��w�6�Z=Oph��\��Q0�l�V�foQ�Q!y�7fh�W��rI�X "�����m׽��4s�����ؿ��i��[�~}�ޏUp��@�X�%"2D:��WQ�׺����u���B��	�8��m��W1	�����[�Q���h�p�9H3Q4��w,�A A��X2E`�"�>&�=��$:�4uu�>�����r&A�@72�2K��$VFW5����u�_@=9_�2���n]_�p��0,��yA|A�,Y�*�Y��N�w�ٗ��VA��K�K��<!��o������%�0z��{p��H��)	�+��%�U���ʛ�}B|A�b�:�YD��ݽ���PA^ްAsW�P���V�Ά��9������_ d��"Ib�JK)_�GU�A�E/;��}^�y�8?A�fw��A���-"�lη����kⵢ�v��v�r�Bk��Vj�m��o>�L&�w��<�r���.�v��A�q��ݥ���p���h� �����>��o=8�,�)q����Ge�R�Y�yr�r������(Ѱ�m�O6��G9;]N�ͻ�M|r�앮#�ଚ���s�um��kK�h�p��Y�����׈�Ş���2�u�6�U����5�ۼH�ƖN�-�Qw�����gm���m@�|k���^O#g�kT�y^ʸ�X[0t� ;��r����ڰ�>]���>�bZ�Z�"���.�r�qqg�.�8�^(G�����f��rk!¥/3~̶]�0���U|�&�V�E1G'N���m���%!r�<�`�2��hW�q�f������s�vf1���"V�����/��гh�.��r�L�v;}s*�d�I[ɂ��3�F��]��ͦ\ɓ��Ը�,�wu� A�;\���][n�ܼ��%-�]B����n!z�U�����:s�R��.�櫱�G�n����J�`�#sȸ��ZM�ҩ�'Ek��q��<�t�o%_U�����fuH�8�Ѧ�z�C8�-����*��&��pp4,Y�6�߲Q ����8�j^P��١�њQ�˱D+��]l�.�S���@n��yƙ��X�e�hP�?vF��Z�栽��:�].<��M*��|�%l(��y���.x�^)��n�x�7%�y(Kg3��gu͕���u	P�&���cυ�>�[m0uu+t޾�������&`�x`����b�$�D�I'#(MG.A�$!X2]���5ݻ�˃0����'uvb̌AD�H�]��I ��F%.�dX�8�I��3M
M��bJ1��A��- Q2"�攰61Cr�S ۗ,h����DX���A���&̩$ ��!%��7M#Sh$	��d�$���$(�$��Q%2BL��A4X�LmD�db`�
*2`+�)0`ғ	���%�������EA���ݹ��""�AA���Ԙ�fL�(iF,h�Fe�E��&ơ6Ѩ4A�HRh�`�X�`�͘h�%�N	�������WJ�`o
Q��M+��2FU��c���uf�k�q0�͜�2��b�n)�UZMal�@�� ��j@���Z$�j$��h2�&�2؉t��F�h�fZ�Z�e���Q�tst��*�jh�R�mE��@j��؎�-nn��R0�Q�&j.��1p]�ꢥ�Y5�s.Hn:�كisC]X132�ik4��$��ʥ;	��r�$q,�1S:Usx��d�pq�,���C��L�G�cJl�N���屦ׂ�p]e���q^���s�����	�mA-c�[�h�%ү--Ρ��K�����[m!
[޾#�.�pƏc����՗�ks-*68�Q���q����o�eĬ72�B��Xʘ���fjks6kQ-�!��[@�Ѻ�캀�.6���^��u�0a���v�amF&��Ô���;,���m"�3X �3j�z��]pK�2�\�Hg���LۛU�<
�#�ݵ,p�0XkCU�B6�aU�����Xd������F�f6��i��RƼKKoZ(��[�4��GP&��Z�ءx�lW5�8�m$�@�)K&ʂcL��&I�0�*Cj��tv��&����1q�4JL���XJ�Ͱ���V�6q����Ƨ3qv�YmH,�I��3�vh�	��hLeج5\����~*b|G��dV\��۞�t�S\�c2.����6�&,&AtƶVlDfM,�r�K����2<�A�Jf�^K)�d��i"����B�*jl;s���B�9œ5�f3h6�
�R#s�a���W8�.[n�/XMDX���HB�[�T��m�2͒��A6i�kHsn���Q�m^CBU���2gYz؀Q�Uay�m�d��&k�BͅA���2��CF�+��Q��3k(f6f"���;Fj�f��DP��\���)oZe���,�xq�̼�<�4G1�r�c.]e�rf�hP�.�<�6���]`*�̰]�e4�&�i����Q��6Z�@��Ka��=P��It4��YN����u�m�y9�8�d�Օ��5t l��A�Y��R����,p���c�fk��t�s�֊:�+y6��X��$�B�vl�m�0��U�p���BXe�j���nK�vsB]z���Uƌla+0͆�n,݇�f��-�cxx�h։^��v�Ii��R��ifdS��/7���	�����0k�&\�pF��a\����&�6�N���YVമ�+B���N��d�	&_�I,^g���ij�?vdĺL��~���+�����/�+"�D���o��yb��f׆�}�������;���ߧ��]A{z�/�X �"�#�'���ʭ�|@ٷ���/�YI,X2R���T<�=��8�{6��g����X%�Aޖ,��~��K��x�F��̅�n/��4$���$�-��2���٧�0}��>���ܯ�cǲ���W�K��Ib̑[��R�t;�"h/�j�%藗�}]��b��p/�_�dA$�%��H�[�O�J�X&�IZ4
K뻵.�2f�X�T�+4�Y��k�nf��LJƚd|����?��gu�%` �d��e�W��h���3p`�gX̐��N)��}C�G��"�A��"Ib����4���7��<�]�+ޖ!G2�ߠ({;�$֖��K����]lQ��\���I��9Rs7&�Q">�|:�ݩ2EKk�<��4{+�Z������4��2k���\Q]&Q�U�\�/�%u*�^�[0o��j��/�("#�XH���{��^��]���w��Wk��ΰ~/�_�DI.�2Kd�ݝ��cuD���_�ݱe�@�$W�{/����<�f��~�/("<���u�b��Ϲ�"u$��H��� �
��彑���}c6��+:n���~{���dW�D,�K�	�.{u�g{��ȿ�5�̭03V�]��*��̱��˲ifL ���\YM�RH]�U�^C��A�,X2EdA]u�ը��ʵ��+3���Sf���GN����{�Je�ԩ=ݢ��ı�dVFf�3멕:�rJG��X�˝WE���](4_��:� �U�,��<��D[w��q}r ���we3�|�I��Y�w&Dkx�aum�>�D�/hs����;�k �VJ���MJ \�E��/���o�x���L���!/�~��;��޳w���κaly�rd�_��\'r/��h2R �d�Ȓ_�1��잮�}�,_ǧ+ ���f�FM�7}��b��_j�3�3��x�r�G��_Ϲ��_ d�Ȓ!(]-�|sgU��i��){*�g�.�/��X%�:�2E`�(r��]���WƄ��((�'M�ŵ���5�Pc��ɜ�k������+G���#�W�9D���$B�����4�5y�KEn�>���=���Ge�J{�+��˺(z%�wen����G����wW�}�}o���en#&��ap0�;����"J�D�e`IZ��J��]v�����ѻ�R{�#{�'��<q;^��ݵt{��S�������#\B̑_�IA$��ۓ����t���`��D���$�`fz�\�Ϳ>�Z���R[���>��hC4�*����[�t��W�:���Y����?M2�-���g�&�T�]y�5*�����J�"�fi7�,��<�0��1(���<�I��3Fy�% A-���E�d��?I,Y�+D��ޠ�w��>�CW�J�FM��p1y�q}��H�"Iw�X&e6Vz�e�+	�"�Сa�ah�:a��qv��p�-�p]-�i-��1��X����u� �,X2R �"��pVF�N�EOU*����u{6ypD�?w��@�D����n���w�k.�d�u�Ƌh��z|��ۅ=�{�>Ȭ��b���W7L�ۼ��¨P35X#ٶ,��A|D�H������|�U>�yT��Ps�a���^wʆ<��̓�7v�'��R{���z�5���12�lX�$X�d�vF�\/ڇ|^P_��U�>�!��j� �܂I�d��2 ��Tl<��;�Rdֳ�Znb�w|�Qoa��.+ �,)��O=U�<��Kr��ٜ�e�F`��ŏ9}2��v�yk��e:� ���a�"�����E[��WE��z�I"I�U�݈��l�C�[)r6[��]K��3M1�J6�٥�f2Vm\h*��u��D�(��P7<�a�[t�)le�S��k�RG�W4k���K.����9k�e�R]-��
J�jX򥴴�-+�mnL�ױ���Z�Vg��5�X�޼L��3%#
j2��v�A�˨[^�VLb�hr�3��.����Иtd�����}}}�ZԚ1.�!�6׊)`Ա�h�X[2�f3Z��3f�&�B�O������@.�H����[[�a��;3�#v�i9I-9A|Dr��"d�&8��0S�J�dg�gg��e0A=ܼT�cb4�pj��~�8�"�H���nn+�_1]h"9�,ܬ��"$��"	��K��o:�����M��=��75}{%�J�"�$�c�ax���r��t\����"��(���9ھs�|2t��*�o�0;|���_�V	�+ �$����E,��u.�=�W�|�+/�����/( A�,XH��"��G��y,	��Vu].)�f5a�K��ePp��4���,;j���E��m͏��~���k��'���)���3w͞-�#�WP�+��խ ��lX.R���YK��O��7����G�bH�v��$����ֻx��iA�W�}�\��"Z�dZ�5�յ�������U�N�V�+��w�Oq{X���r��(��˴s�� ay�j��. ��9m*��y����%/�'dV?I,Y��"�"�9��q�����Y�Gg��������;�e��I���c �� V��k/�uʍX � �#{Ə�U�Ɗh��#ܠ��gK}��WWq� �3յⶔ��t��Y���2PD%�2Er>�Î�79��Q|��]X�y�@��C�39X ���$�/�"��t39$�O��օ�)ë��܆�.���ٝX�cQ�h�Ĭe��'� �y�듬_���"���s���e��v�з�b�>��oH�%�e ���2r����X�A�/�%lW㛐�l��t�4~��x��2c�Y�SL��fE����Ƭ��b̕��$���zւ5��`�(	"�/���}���un�����z�U��T�k&��1~�IB�`;Q��Х\0�*���̄o ,A��Vc�mF���*�Պ{�m�i=���̫>�u�^}��g}4��d�3wh��ݢ�݉���ϑU/{mg����x������Ex��ɾx����K�Um-s�깅����?8��!�"��$��f��?~���|���ѝ>�ak�}uY�Yl�/�%#��8�Uz�Τ�0-%��s4*����	rY�]SG3�4�M٤14!�tU���V�_��0����w�}c��ج�������8P����W��
�:���U���4�r��$�,%"2E��J����ٗ��ܠ;�ϲ���׏Q�tpۃB���h Fȅ�"�F'�5�O ��w��c��2 �"I_�	%�~uw������k3=��zny�OZ��^�7�rŃ%"	�+��"�X׈^����@u�dJ�k�U�����@�y����f����@�D��7��Jئo�e�}I#�H[vj��B/�v���P'enc�VG�dY�^��E+L�='{ےb�&r�5��({�#���X������[0`71X�=�My��g�ΖU\�O��^�=ݚc$C�j�����^:E/�\j�PJ�rUM��[�f]��G�u#���fa��f-4R*og��ɫ��A$�$�{={��ne��^��[\=��~7'��=k�z����?I�$�,���r�U��>�YD�޵וzġ�u�P1^}`�gj��	!=}�Tm������o�ma�_\�Ń%/� �{'��w�^�R��=sR�¸f����ްO�����X�$W�H�"Iw�R����wW�?�=� D�b��!g�s���̷��מ�k�&�VB"���a����A�� ����h�L��%�$Yx0/?sĲ��·z�S�W�t#=��@Ǔ��;W�"�$���}�x�Z�P|����d�f߮�K�#u��iR%�N�z����p7c��0=�Q��fL��/p����f�|��ZX�m��ok��^����ڣ~I�m��f�l�/�����䌥��4�ۅ�FMn��KF&l�s�t�ˮ��8�h�D��f��[XP��ȃ��X�R�*����Z67U,naZ��uаfs\:����T�1���qT��JJ�Z@�\A������&wP�{X��Yp���b�e0eF��fE�@�X�ix����״6`��3A#[��֗���OM�v3����`Q�v�ZV�4mUV���7mk ����n�E��'|Ր�_I_g�H�f.��WPT��T={�����qő�� �;_Ed"�"�Y�S�Q/%��=�}��!αnz�9�Oۏ���z\����Vn!`(n��+�HPz	�ڰFλ���2Kd���E^�Y��Q�;�t��w+�_?g��u��E&n���K&���(��zs�2o�T�X�%|��fWfu]��n�nw�>�9�{�wj�_�a��%�&H��� �N�b=�l1�z�X����}O7O%~��\A �5`��rř)|A2E�>�u��ۏ����,J�m������$��A�#X�����-����dPoD,�Ղt*ҺP^������k`��{±���I� �����H��%"2E�m�g�o��X�`�l�+�q�[�k}����/!��	�B�#n��;����Gw/f��/$[8���ez�އз��c�:���c1go+��A��A���>���"�ge�*�{�x ւ��!"�J�]�d��ܫޗ��ۯ=��m+�K��&y����`�H��YD*Ͻ�Tw�A���,��%T}}��:}�ۖ�c���g+#��+*p��l_��2R �d��"N4o�oSDl�[p�?T�~��GW��
���ΰ~>�}���H?H�x���=�l�w@{I�`��e�Ìf�M��қ((+6B뮘��F�\K�O>}�����X��("$���D�ōY~�]���4ak�y�:릔I�j���N4j��|AH��!�JyN�;�����F���d;�Wh����#��-@ǭ��g+��$@I+�Ȯ������_P�}�I,X2R?G-�]�Sq�k<��Fe�ua4�*%�N͜��S8
�N�pg��/"\d.�"o��Ϋ̻Zp��"ݬۘ�a�*��6���f�������K���˙�@���/'[b�npT�<�����I��oL��Tw���\À��x��i�48S~>ʌ����(H�D{şJT��P���E�"M��w�r�e�K���(۪E��ˊP��B�����r��b�u�r�*30�3)����=y,�� WT���;�F7:�<P����(u��%\#�[.
i���s��WFf�%���&)w���Y�<�Y�������4WYA����tb[��X�gq7Qh���3y��1�K�k&�^����眪�w��wG����#J��"s�vA��-Q��j�	���Z!n�b�R�r�˔x���(٧�[�Eom��UneQ�8g׾+Lu���0��Vv���85X���7�$� �S]g/��f�T��U��˲�wU��3��r,Y\m��+�j�]�'Q���J�=�gU�����*�K��j�%ֱ�q�CT�%�=��عen��P��P�yc�A�Q���tY�Y�F[qXPdX�:��ő�}.ǝ�E�q!~���[T�1��a�s0�'Wa�.����8*��2��ɷHz�f�����r��d���	:ݐ�p�w�o]�1	��Vjf��E��%O7��	� �4�l�
g)��$���%^]d�T-W� �V��Q�V��~ �O��	F���@Rcn�@��r1c���̤b��)5%l�I1l�$lɘs�I��D��h�sr幢�E%)�BE��LF�ƙ���h6�Q��h�Y,dۜ"9F��D�1A3�,E�PF�r,�T�AB�%���a�A�]�#m��#����L�4��\���f�����&F�%EAR��E24&�e�A�4Q�X�b,��w\�1�b�7-��QDQi!"(��h�hɂB�BHى��"�2�����Q��|A$I$ SN�Wu��؍A���8eD�}$Z���`�������ü��"N�/�"5o��_4��m+���q�x� A���T:,��}�:����M2P_d�,�]��`�0�S�������z��9մ��_�9}n $��d�-�\W;ĻZ�:a���\�U9�.GM�u!����H�ꄦ��"��%QWˌc|禓��)�ı�$Y���g�U�|����5�yUtw��+���͢����ݒS7v�)"�/��p��1q�:K��/�[�i��4ߺGJ���]�Ǌ� �,X2SN������z�|,�j�׷`���%����A �7*������c=ˬ��g<R��i36	���L��d��{}��f���?N�,��?$Y����eU��Um��s( ����]N����w�o:�.���i�M��������ڣ�]cRּ=�sA�/�X�[9.`tF+�U��C��ϫh�C�/3(LJ���r������� �E��B��y�'��B{��?V�%.i����R�C�1��ř)	�'��%��ҧ����_�y��������ݭΤ`�%�lX�$��	z����uZD�m�t�_����f!�س$_X��^>�LT����j<���ƔA�SwV����A� }.�"IIX"�E�����3���u����y�'B���]F���P_~�X�d�����n�m:�������^�M!�ݒY��I��Dsw���&��=6�&�ѺW�G�����C��I�Čc�١��H��s��D�v�����{���Aݱ���"z���ވ��v�51v��Z�{��u����FƑ�X���_�VA�+ �/�)�����oe%�b��t��5x_�-�`��A���-�k�ߐ��^��{kkZ�0��D��΃����{v����+.���F���c;�����v߼ooF�yN����,V�c��se�$KY�Lb%����FJe�������6l칄!y�6�1v���c.��4�f�X�Fm�*Ė�;���-�Y.pj&^�d�T�k	l�״�L�ZHLK���,e�1@]�q��Mi9-֐�l�Ժ�ئv�΅"��1�E��B�Jef�Cf�Q�h�Ўu��@5��<����lH\-نc�k��,��僱�R�c\�ع2Ҭ**�������X&MVD��%���,j۱�����+�I��B�^���]�3re����־�X�$_I6���":�&����T��>�VA�^����O�]����<��;W�A�}���*�r�E>�$kٳLkwh��ă{�^+E�T�u��^���Zo�����E�C�e ��X��X �DI.�W���~3{��q��#�]�D����=������_���A�̊�"�����se������Ş�@��ފȒ!fJd�,���qu߈�C�=I�g�<gܻU5��fr��r�I.�2K�.�^��{�D"��HػHXA�vA�������^]�@�a��0	s�V��2�*��=��ř(	"�œ�B�UU�|L/-u�Wm�<��N�� �D,����%:TP{}�~ԏ�[�V)�8^p�V�s�v&{E���{�@�ݽ��*�쵻z�hGk� ��oUc�7�(�f/A"�ݞW�C�ol���5^xj��}�ׯ�]q}���{���S�0��Yc;>Rm��Ib̑Y��?wv�ͮ�����mSP1�48����@�%�/�$�,�H����$��+> �$^���Tox�xc�`�y|,�����r�<��k$�o1����� D�ł�X ȂI���W�α����N2J�)��)\ ̊� �,Y������|KS��y����l
�e�����KYU��KT�k�mI�8����l�]\i��}�� �P__u�$ZD���b���Ew:��c�|,!U��w�:Q��k옂e望F��ݎ��vhj����ʚ���O|rR ��^b���[�U�������X'2� �,"Z��Ո�k��6����B�|��_$�%�C��|�����LS���e�ɵ�<Ͱf,�A�	꛱]��<#}H�ۿU�沶��S,:��-d�EQ��_��M�G��>�=�<O~�x�R�Fd2{~��'��$�_�J�"�$�,{�q1^�z�T�ڥs�ܯ�$���^�U�6H�ΚP0������#���<'K=��j�i:��92R �"��/�%_�T�1P�
�oW�4)�UW��#e���#C��X ���~��Ka�M�X\dʤ�Mn�a�[
(����*ElR���k�iT�������Ղ�	"�$�/�m('7\$5��OW��(��B�i�xѡ`Ԉ&H�$�,���?L�VL"�s�O�"���.��nc_s-(^hq���?8�I��<���v�g�E}�7f���C݉G�">��^|�J��ԋ�UW��#e��9��X�$_IC� �o-�Qr�z����/��XĖ�(&�\5��OWO�+"�$�Wl�j���z���D�n�m�;�|m��<�_���1(�e���(:;�A��m�o=<uX�����S��������&�%A�Ib̑�6h�B��K;%^M>��J�ڬ\@I2�"IbV���/e�w���>,L�Mm��hQų	��܆��,�69L��,V%cM>|��C����$'�ߘ�+�d��b�mqOҪ��r0`��ޑ�K�T,��������D���$V�U:�����4��]�@}�/.�v�y�
�y'��q�,�C�s^;�ʽs���R��z	�v�Owf�읒���msG�n��:�n�q�J�}CO}sI�f�,�ڥ���c���.�+�Z�+Z�A%�Ұ�d���k�~�U�����8X'2�fgU���wi�p=�X�r�%�`�"�A��N������S��!%���n��w�z���X"8��% &H�c�:�Ь�n���4d9^`�קɊhA�g����xm�m��_a���B+���H�ǣ
}eY���������5:��Gx��v;q�Ni�*FD��L���X�7VFQ-�Z�&V�.4ҩ�Fd�`54ҳ,���i=S�c۵Ŗh�6U��KX��5v�d����(�u���[cR�#]Ţٵc��d&�e]�+\�®3X`�Fe�5CMt��11j�!�[��&�m�̻�6̍�W�%�K]fѭl��Pf֙�3Pf
u��6δ���{�l_sb�h@�ѭ�,z&��aV�cF`5�v4U�3.��a?�_w���-��"5��9�g=�P0���&J��fޖ�p �A�]�D�����d����b���X^׮7Tşe A;"���4�OҪ�u0yb�ޡ�b�m-ݞ~��ɳ�rIC9�T0<�Y	L��2K.���V�^�.vp1���OW|A�Րc�,+��+��%ز<�����ޡ�7�b���dIAz�fpǛZ;9�Z��o��@3�X#�3�=N�֞e[�wG E�X�����+ ��~Kd����M�}��7�}����?uUc��`��`�s("%�2E`�"�z�v*�u;ߐ>�_���Vꋦ�Eԗ����R��Av�v�@��~�ÿ4�����Y~��$�I��v6�	��	z1������WFW����^ �v,�H��Ȓ]�������#�*Y��6����{�.H�����u�=u����ʼe�u��^�l��2�a)Tcx���̹On����O���s"�A���e�p������a[C��V!�I11D��[��3`3���^R��;��A�X����FH�k��� ��S�>�3��Ϊ��r0`��	̠�;%�H���$�,U��'�V���^�5�� D��H������M��Kэd���j��ld������n�3�����&� (/��/�����^�7��U�� ��}�2^։���@��C����!�"I_�Ib�;���*"���wi:�x�5z�ƌM� �.٘j�fm�l�b����TWU` �n5�|��(	"ϳ:�O]?J�ǵ����8/w�x�[���"�lY��� �!fH����?V���4�=�6����/�gk`������=_w����#�X2R>����UOZ�DͿ�%"Ib̑YD01|Q��*�D���\E1u^�92���l<Z�,��u����Zٸ�^�K�U��S���	��Ý���nA�~z����"��sw�����1ڨ�}`�;U�C�"$�/�$�fJDny�y��o��\�e�@�d�����<m�UVc��,�,�A�f��^����7��L���K�X&H���$�,��{z�5�����*G��v�O�эd���sV?s�,�_ d���v�"�_�������,X�
���:�*�ɜ72���nMcs�.���5�4�>���{��4!?{��H�dA}���nS����j�b���]|bz�=�@��"8��$�`�H����t��������n� ��Vg^i�v�X�Q��u�e ���fH�\�9s���p�@��`�y�`1���ݪMn�����[�yp�Ó4v�Bh�y'�� �}�Y���FH�$��o�{����0`;ʄ#;P���VD��Y���ON��c��b��{�Y}:��wX�����M<�a�;��=�����+(8I�����d�RxW� E�7=��Ao�����ۻ+�P�x��?>�,+��+"8��(�AoǷ��xجM��b�ļ�j�A����("�b̑_�I@�Q�h���	:*���!��X5�YB�m��0�D�Qu��V�������߆ՐD�"$�/��x����&N!�>w�z��b��J]�mY�&d����H��m�%��[Ǣ�S��Gr�||ڰGu���z���{�0�b�C��VA �r^��5=�o��j��|�2r�K�"��7n�œJ�\'������2�B9b�2E`�"�%����j�W�ݎըA�@ov}$��Aj��{���y'�� s_YܿC������㯕�D��d��"Ib��$>w���qz�Wj�{���]�-	�����K32U�|�$��$$ I���m�}���m�kkV���֭m᭵��mmj�[kkV��mmj��kkV��m��[o���ն��IX�$�$$ Iu$��om���m񶶵m���֭����@��䐐�%� �$�$$ I�(+$�k/���l�[�B,�������73�0    �                       π �u@ J@B� � @H(
(�   ���H��@B� ϾTT��R�(@�*�����T*P�TTJ�TUT��$
T�H�J�R��H��Uwg �RT��U^�U���;��j�W-J�"ܪZ�J���K���YUS9wU,�IY��)���(�N��Wɣ���Q)�)H��W6����	+���z��uQ+��+u
��qF��;�t�v�mWZ� 5E
.�}m$QEH!H��W�i�G��@�y�� ^�y @��҇�@��޵  �t� @h(U�-�p�{��'uy�{���j��:�  P{� wE���R���vi^z�t����,���J*7wR�Y�U!q�����R���Ԋ�0޵k���B�(�B�� >�"�TT�)
�W�UUf�*��\H�6:r�J�訬�"�2ݜ���UBi/f=�B[��.M(��]]�
 ��� ����QL�֩\}![��ky�:�^�r�\ڧZ�s��S�L�����$Uroc��y�Kg��C�ER�AE| ��PU���B�H(q�*��Edj��nfET�p�R1ʕ�z刁�����Uv܍H�Bo{
��H��0�R�QA| �u���ж�%SܕUgJf�	�I%ɑGZ�TR�J��t ]�d�$  S� <T���!R�T�)�Jwq�V�B�ʕu����aћU�r���D�̪�u)-�V�Pn�PPJ����(��\o}^f�M�UV}*��#T�6��6��3JKr!]ҫw�] �m �5K�    5=���h���1�0�2d 5O�dJUS�F�L   �L4�j�
����Ѡ� ##FL4�*D�$P�@   @�	=RIUS��	���# ��0$�A2RM '�OF�yM�L5=1��q��U�W��7_y M,��)�g�0��&je�3/�H�	�W��tJ?Y$� �?쒂LI B�HH�O�I H�#_����Q���d?՛I$�!@"R�H��$x�T�2E	�$H�MU���?�������䐁 y�^q+�~�3<i+�W���@� �����/��.�?�R���b��Gf���R��wP��!*L8�����p�˭���f��V��qm�J�M�Ś��Mꪬ�1��L6t�o-}o/j�*�ô�B$�����e���`ș��ɗmB[���d���U���f��KUF��ܳ��l���auX4]��;�*�ʪb����^�n;�eRϐ���mL��vc��Gj�����n]8�t:`�p�3��4�5�{[�z��E+�Tv\4�V�F ɫ�x!ԫ�u��S5�n�cv�AW{y�ޛ��fY�Csf,�uv��y�D6�#b�X�I,l]��[Oa��J(�9Uaf[���5�Ыٗ{��,�Ӕ�R���U2��F�#�g2��YX�ʓ�y%�B����wem�s*����4��ُ*��ͩ55(�MV�]�"8.�F��xsb:�V��ʛA4ܰf;�������%�K[󭛹WF�j�(�m��&a�b-9���v�U�7��Gt3k.-Q�ATѻ6� �MK;��j���/		�̪y2�Ud7xn�AI��Y����w�3)^d����r��C����6���[B��Ѫ��+\uv����V+��$�7r�U���ō�6����X��Ǖ�tn�U�%���Gk6tdǑ����{�_���ڧ,�k��eм��"&�Z���ma����Ъ;T�k6(<��^:a��2�5#��D��1�G�\��jh���N�P�R$#5T��[%\L�����Cz�#�HC�Zݩ�a����A&���˄P�c$ԡ�40�p̬�t
v�2�Z.�,�I�e�{��f��Zj=�$��YXؽ����q��r�n��e�1
y��r�v�##��ܛ���W��J�Z�)N@���Xn3lf��,�1|s
�	-����3C�ƦM�vQ����c5	T�&���yCE��EAx�`n�o"�OSXV��ŹmV�L{b�{A@ⷥ�4����dVY�T򭱦�)4�4�ud��9*�;�X���U���Ww/�s"�Ƙ{�H�HEn���n�ԉ���[�UUb�R��[CR�#��̳!Ta�4���8�CW��)Xp�df2lU�i]P�R���TTH��Н�d�tݭ
K��^T���1A7V�{��������4�2r�i�[�ůl͏7ޘ�L�L9�4mC(72�����]6,��z�A��wF����ذfL2��������sq���y�R2�S&<f���x懧k��Y��6��\���s��enM�ݛ�nd"K����;Uken�R5(�۷J�K���b�Ї�yݳ�F�&��u3e�ڹ4�5��8,�e[���w2��enm�ܱ�v�[�{�6)W�����
�!
�%�7G[�U��[zm��WI]�o뤲��G��~���R����m�U�Z��I�t˒��p����K��C������v�Ax�w��ِ��{��,���1�:�3D7����֦]�ٻǕ�-Fpe8���,a�C��B�j�%Yٕ�%f��4��R��'1�me�yg F�+���4�	Cv�-Ef�q�O6��cL"I��5��j:��q�K#Z`�b��5���Ǩ�[��b��b*n��Q\�m&`X�epV�)އwi��7�۬aŮ[���3U�H��6ne�D!R�2b�/+wf$�efm����L�t<��T*n��X�F�tE/B�;���a[z�Mk"�
miمARd��idz$���GY��N��KE��Z�����uwH�w5W@��
j�f#���R]���&��TZ��Y�ɭ��PF���wㄌo��7Lmm��K��$��5���&ZD��N��kr�gۂ�Uia̯��w2��kT�J�,���^��U�Fn�x�v�V�ʫ���-��h�"����&�ṋ9�ͻq�i�P�w�j�y����T��G˔jeAO1���:x�Mky/`ˍk�kY01C���X��U	"�2R�f�3�ه5�����4�ī���pJ%�75�yR���چ|��yxwt�\62��&s���C*���j��nըS�P˖40��3Y��D���ܸ+Bj�(^fUI6�5���6�rh�B��ڹ�,��e8�ݖ�mXy�[j�@����F�2�ν���L�W��+��7�Um6Mے��j�fŴދ�*����P�K(��yy5��I�N�=����:�Y�gƥ�ܖor�d���F;�T�((+h��R�� 䈱�5s�K��m�F�%ز��X�G�������d��`�j[�n;�MhE�����2��%}��]��ɔ�Uo*�̖��wf�So&f2��!��ck"'p�B�ˬ��#S���Պ
�D��
Cő��*�L5�v�9�Nh<�1ݭ�eͺ�MU]�o*�>Y&^�j�0j�R�+E`ʧ�NV8�!ԩBL��b�r�Պ�z��#�Ua�@�l�+J�p���\�-���U���	aM���/ݼ��2��wi�ٻk	ZE��f̣��]���WN�/ #Qo15f�Fq�Hc��n�(Wļ[�K�6H������k����6�TxF���<B�����wb�]P��V1�G렔͙��+D��x��m2�n�MWgY5M�t6�[���Y��oB�m��ք����Kb]I˖f��+ϴ-�Z�U��b���m�bL�Yƨj�z����%�7(<�9�Y�6R�������"�ٗ���R��qꥧ���WQ֫5J�:v��Wu���,J��n����c=wD^j��9�1��Z�Y{F�m<��b�m����f�b�l�B�^�:M��DX��iƶ�^n����WU��,F��#���UECxun}��ʍ�J��<bQI��:�.��7����ӹ�j�M���Xn���b��g2dl��V���찍���=��E��(Wm���/`�T�6P�	�V�%�$��֣b�I
tR�ث^ed��Q�3t9Ϝ�b	OZT�V+�hh���<��v�j���R���]jڦvm�5Uf�$��^��ݼ��Q'�B����^ܫ�f2ŵV�����vn,c]]�0���ܻ˼ɳ��V.
�`�}34��6��cof�WK��͵dn	WW���n�a�ͻv��h�T��n���-n����v�m�Ar���m�͚"[v�<��k�7Wl�uSW6�K7t��W��H�r�neUf��
���5y&n��̺�{r�hiY�X�a�0]K��GXk%�
v��z��yQV,6��VG�1صz�g�#2��
5�QJ�0�3ot��ǖ�� �j^L��nh7{z���.��][YN]v����Mњ��1K���)J*;W��Z��+H�#6)�£����SŨ��7�l%��r�#��:sN�m��n`�{��e3jj��x����V\mÈ`�t������($�D�7߷A�v�W�#��ݒM'�<�F��Ѵj��E�4�:�3I��Q���X�4S�x ��j�V�̙,T[Mi�o`�S
�(jٗSY�Ef��u��^d�&�.������o-�*\����nUft+i�Z+"��Y/�VY�pc.�1��h× xa"�\�]YG����5ʈs���Z�*Vm�9&�����PR*���u�%�Ƕŕg0�U4������ɒV�ͨ)�ɀ��+w$��=���yg;�dL�h�R˭��RL���t�i��GRe�zi�^7���"W�X�i!�����e%4Ѻr�V��W����8+.F�ゞ�ZN�͈mܫ��Bƽ��F!j�RX�^��MP�\$D͌t�
�K�D��
Cm��䳕�a����!*�t��H5�Q��vl�A^"]W�1����^�X];�
���R`�����!t/"���3r��d�/D<0�
m�K�+u�c��W*�7x	����l�EUX��Z�K2Ά]:�����sl{�ʷrƈ�pnU��k�ک�Sݬ��j�Ǫ�R�c�mX�)l�'5HN��Z2��l�7m[:�{E^��m�����"�t��naa��lY�;��5Z�nfZU56�j͝��3"ܪfQ�y��qV`�)�TmXYjeR�`yw���`�����X���hb�N=ʧ�&�C#E�۱t�N��$F��oX�����k�~�f�O�*���.��A^n�e�++mf=�V��b�e�;ňJOj�n���dm�rL�O
��3N��	�3~��Mb��̘-]��d��d,I��V}o�&������-��%f`r��U� �0�N'42�EX̷��|lnR�������pb���m�12#���O(bb�U��o��9���̪��T8v�t�m�ӏx^��m:.n��6�xr�b�Xd�LP�4�M�"�by��YS�*�;V˘���d�&*���A�o$r�����:��ޛ\�rEDDl��4�[ܯ�'�P ˷�,�TWV�f	�U;Z�ӭ���ӹ�M�人��VnY���KMGc1ƭR���Ʈ���KQ�N��k�2�e��m-8�U���v
N�:���9���i��Ӳtٸ�^�7A��&�u�������2��k�n�����L׈iǪ��W���n*ޒwM+�n(���X�f�;���2��v�M����*��k��:sU9jLї
��u��wt�eY�md��.�Vn�U��m潡V-=`֬����`1v��vT`�ٌޜ����$����P�h�Ve���q��^�۫���a���+j�j�Q㫤0��%u*j		�Sz)n�[t��@��W�b��іn�����[u.��Z�����Pͩ&��U7��0�k[25y�����V�n1jf��.XL�*�VnӴKbe�͓vΕ�-�R��;�XMD�0M�z����j�Uч{nժ�S3l���,t��0�
f���Q�XTD���(�K�rã����%87Vl�0Խ�M���t��������Rt)�Tj�	���e�N�[YcuM��B�(�����d"�f�YM˼£t`��X�5r��iͅ��W2TZ��U9��+.�ձ=u�X�na�(`�V�S��-%���]`�GM�k�)^ڋnR׻���E�j�C���+4[�v��Wa
�Wl�Cv����Ք�ݵt�n�S�m�«O�U�m2��%�n�ͩ�c(��][9$�v��-__V[�ٻ��[r�ج̷��1��`�G���&�E+�F���6d��1��c�E��1V6VÙz(5�f�h]=�;V֝�)��2e�P��f#�p6���ۺ��	�˅;3"�I��Ɋ��,y�N=�א�pQ���)m��{Z㧺��4ں�5M����H*K��&ب�ef)�`؝V�M�I<v����T�M��]��L�����S�Xi�G7/c�m�u3T�l�y�0e��,ʺi�;K����.���3STB��O.�����tu�r�A@�hYz��ah��{gN��l�
�Į`�
�2˪ܱx*��Mnit�S�V�\Wmi�I�nZ��,U���+��\�4�]Xoe��sZ4MޱeE:�]��U�iF=�>V�V���#Ъ9G"̭ˉ*vw+�ƍ+��M�2�2����6�nd+L	�ޛʙJ��4oS���ݳ��i�����^����.R쩲��G����u/6ī�*`b���w����*c�X��zɬ�d����?O�ϯ�?���~��Б>��\�Q���|�ϑ�*HC�@$Y$ŵ���lj�EV���m�6��6��5��X�ړmEkI�TZ�V�Z�ڶƵ��TV��b�l[cm��Xڶ6�*�ƭ�j��ح��6��j�m��mb֋lm��UF�m֣V���m�Z�kU�mE[TZ�-X�حV*�EUb�F���4kZƫ���b�֍j*ѭQ���lU�+V�m��֭��[Qm��jڋEkQ�X����յ�V5 �! (�����ǵ��oʽ��!$	 ��'3{�I �ya }�x}���$�ٱӚ���~���]�oxwu_,�>~U��wy[�$�x!��FZ���e��[��e.�G1\Qܺ�Vlc����R�@�x�WWc��Ҳ�J�b��d��	:t�݆Ѭ9*ͣ7D�x�����ziz������n�I��U���Cܩ�ܢE�+�ed�B�L��5hT����a��(k���몪8r�L�8���4Cu�hn�.��c�n�{����/���Ys�a�_UcH��%���2��5�%�e^ї&�N�P�sB�Y)���7*
����j{�)Rh[cMV\u����ou<�e�r��(��Z=�w��_6Ȇ�VB�Ut;����;pfu�.�NV��8[�Nv��U�_T��<ιK���vdig�a#Ճ�}/�m�a��eЪ��[{@Z��r�I���[[����*�nPkUKoU����t:,�Ī=5+&h@�rI�)O�QT�C{2ݴ�j����wD-(rC)*��#os2�_аz����m�Y�h���Y��L�g���-���W�n������p��Y�A;�M:�ybRcu�A'��e;<+�5t�W]����,��G�K4�M���feb�`=1A�BA�V*��ЧwR�'7+�-^:%����v�ۡ�Z�]F�����H�\u�ڌ��&s"�i�D�*�Q�����R$Y�e�/sS��\�em��nZ���V�{�߲]Yvf�.��� \A�����՟�}2J4���#B��:���Ԍp{���*
MX����-u���Ps��]��d���ƃ]m�Zr�����a�y	V�[g����ƭJ�Ҧ�
��p���	�#]����f�D#b����߲UU�fC}���&�;��^\ZC�ڗ�評v��n�ЋKTh"�M'�6�U7�{�1J�t��[H���<�nw.<۬����r�o��1.)�R�jE��ی����i0Ӫ٪�[*�]"�f�v�FKS�w��d�i�R�!ɇK.(��f	e���i�m��@�*�Ǟ���v��R!�0+m�hSX�R`�$�Q�HҬ�Jb��C�����r���Fi�
�l�:�V�y�)U��ү�j�vٲz�k���eԤEp��X�";w&�|�1�[=rgKV�r\��5�"s�,R��j�ј�ڋd�����w�f�Լ��/*�ՖؕFj&fz���0�wT�p�)�@�w�R��ja�̦�Mv�V�Zj�7�V�bT�7A�S0i��{z{	�T���ӕ�uq|EQ�8����W'W�QeQПF�u�˝|�)юu�Ng�y�+����U��]B2�BIM]NW�\�T,˺2�˰�e=}�uPT&��{�57���-`��&a��e���&f]��.�:S��A{p�{�)V����Y3j�)�.�R��k9
�&J�J���
տn�[�J�5Pˬ9ZZ�*UҔuQ=�{!JZ8��|�m��\�V4���H^��7��J:J�X��(_D35�`�}�%]^�ԃԡ��*8GW��TCR[n�}���pJWWkw���+xBnTδ�m�R�,4�J銆�ʕ����6��ht��@�'�tۗ���fp���;�h�˦��.�l�*+��Q�����t�.����m�L�eqV�'烢�iIY�Wv=�*1�`��Zt�e���i�WZÅ�y��=�[p����;�=bRs�%��X|/j�1��hS�!��s��8y�
���K4$��SD9�����*�:��BUˤ��u��+	�S�-��.G&d���f���k����/��.l��K>�V;(�n]�۬a:N��`�	�JNu�a�f*�{B���̐ojd��l>K#fj�)�(J�yN�����O�n)/N��rh��ʁ��'!E�s8�闕��j�zt�(��uMti@-̆���]#6u�W�r���b�I�]y�qν��m���۫�ख़�*%oj��8�V�st�5p�X����gm��.�?n	�6�,�첵S7.���o<�L���v�_�e[U���4>�ZNٮ�ὫuRq{t��<p�z�7w8*0gK�jg*��\��W;��u/3t��S� �=�֮�8nC�Q<Z�e�9eW��;߹ǽy�1t�V��u
!���_m`(Pz��������汖&��7z�Ww�B��q��g`9}���Ղ�,��K��x$¯���Թ,^7WN�onZPm���.����:\�L:�,m��	��2�_��Z�n;Q�H��V�#boj\�y1N��Rʅ�mX*�e��+(��Րq��ɇ�t��N�iEز��`��G�6���v��6�rAp�:����T֫�E'�wgl�Z���7��� �]��R�P���x��O�ݱ�bʭ8���(8(���+�7/e�0�Xi��+���gDAu�j���V�]�*��9��=9��(X�9[[���!��\+M��6ݐ��.�3٤��g.���5TN�Z�G�'N��
|wo/����n�غa�ή��A���6F�bĸ��|~�:�4��v,���k�#��x�Q.��뭔��U|�=��/��tw�*p��sf���u�����U*��]1�VeDԖ���]51gL�]^�z�Iw\]a����zO>���,�_tv�*��W�ﲕ*�q�X�&s��2���/�����jxޔ��ƥ�R�;��=�/n`"�/f�����12�70j�.��BV&�u�)�E�;({2ͧ{Pժ�JF�=�S!!r��Ur���̆*�:�������l�2�����x�Hw�y�퍧t���F답��Z�U����{j�b�Kb%���C���]�e�e�7�p��k>��Z����sc�x����6`50��VW0�*i8���3�h���޸�vM�z�q�ՙ�5ak��*�/���x%���N��ՓH��j�ET%suT5��:+lEU[ل�G�LĻ��S��{s����pR1��[Z$5�DiL��F֚�UE��rɖ2�Tm��ya1]n�b���3wl�ה*�裄˥"�EQs:���$�f�B4$�N���i��a^e����-5
��N��y�5x�*�n\uu9ݹֲ��BoP24�8��P�]��MD��UC.�s�-kp���|�u�ͮ��(�78)غ�٬cF�Ev�9��D����z��QU�u��W���d#Ʒy~�eVj�@��o)���7�k�ǲ���L��R�5�FNj?S�N�u�.�o�}VNW]e��H]BM�b���$�T����V&�)J{I�*�Єf��D�MV�7/)9T)T���R��n3g��h��:aUz���ڡ{�'8ff�?S:b5y�$��%�Ww^Bd]T�����E�d��'$��}�N\��,S��|�V��bZ?fb8)A��>WƟq��ǈ�}X!�)���RAW��Kn�|�!�t�E�	1�G3��UU�|�LX�Ѩ�X�u1��UN�;��o��s;����yx1�9��,��c�9Ղv�1F���&�q���s$@���9qU�"OZ2"NN�EL�z��[f�e ���,���.eWU�}���꿘�Wuݗx�f-���γ]K!���Ո��u[��w)*�]�
�8�X��&U��N��6��j�ܚ�&�T�]�ĩT��V-���5j�#�+��h�+v��K](�s�g����rѠb����N�)�J<9�{��k�Ԧ^Z�nV����gS�ůYWLF�L��Dz7`��\f.'�����"��P;��xE�XחWWJ_.�-	�/bw2��y�Kv덭 �O8쾰��`7_\ۆ�n�U�<�H�5
�2³A�`�h�S,g��fN�3UK�iw�}fdǬfu��ā9�G���=��Ki�����.PU�Vлv-�6��w�WcU�&�϶����ff�C�tJF���gt%�����N�d���A���T�ʰ�qY��N�/�*�D5��Kh�qٵvܼ��N1Z���	h[�Q�l�m�X	�p��e�V�gru�ޙjm�[�KY��d��^V���Ұj���֧#ݘt�95��(�F)�*�'LΪܕ��]���8�����G
�u���/U�����d�$2�;i��%����)
KR�nnU���2H���1�/շ���dX�2�=ҩ�-$)Y95�o��˥K�P-�X_k�w^-ͮ��s�E;q���A�fk�T��Sr�e����T�\��K'���2��78��A��Bn[�-�� ���Qh�YcyU/�p�3x���������&fvm�����v�b ��a�mF���qf�{s�!�ѻ�1��t�7D��6�r
�*,e!(eR�6��33�xa}�/R��u����ܴ�L�6�����Ѫ{}�*X��,[�ͯ�����b���[��X���J��<ͦ"f��1^���z]��/*�;a���"k�;�ќ�/��b�;�t�� +1P����n�Ɔ%98N�����Z����Y��Jn��f(V���ZDm��q�A�侫�>�7,��������݌a�ɜ�z�J����>26�m�W�]"���F�c��"�5��mS�D��4$�2��lYB�^2��c�v��ݚyb�I�/5^�NhP3{�&�&Z���rd�ޝ
�}n�
�r���.��m:#&de��B�D H�Lٖ��n`�ywW��֯;��p'm`�|�YI���wY��Ar1>X�r��N�sN���eR��:1j�6�4*��:�kۻ=K��P]�.�v�m�I��rK㗜��.��w�O�n$Z��|���9��Rӭ�����7�3�V�84�ed�F��`�CsqϏ:��`�<��:�QoG^A�+m�WF�vAf�Ũ�����Q���aéZ�'C/�F��6i�Ϟ�X,2!��Cv�d��.���e�(�޼{E2�)/YѸu���ȊZnPք�U77j�t�a�E�}l/�uv��J��<u��gf�
ݻ:�5>���u�Z[�R�O�]w�V��Y9ݘzl�x�%��-C+9[�̥�w�Y|ծ���V,�gs����RF�/���}�%�fwn\�W���I8����:��B�A�r�EéH�nh��MS�KU��&2n�ۑSU{žl�[���-]��U�3�*���jɛo<�{i:9�O����Q��G1W��)S�1�G�	��0i���QuQ�]BV�a}��b��vB-ΩR��\���*��̍̃,��S�z1�FE�r�EI{����u��GqرN'����z���v����P��]=˼�bhC���Q�r�j�ٳ{�Я��[1Y�$�T�d�%:�è�ю�Y����T��;��3m�X軦�ƛ��]Ȫ��V䧰q���F�Ʃvu�U\y�a�!������S)����iS���w�-*���,����- E�����	5�ݳE�;0g+�:���R����F �UckY{�P\Y�-�v�MЌ\�|���;.�])]{���сl���m.�v]e���Ó)d^N�ڪ��5L{�
4�h���֕������W�����n��{:�.c���/�%��-�V���L���ܼ�����bk�JԮ"�8{-L���z�=��e��q9��:7VI�*U�����+�������;r�n���(ܝ(7�x����w���S%�O��W]�Z�.�J��Ηu*��q&�`�1��1[/����� d_�!!8�"����B'=޴�x�9�m�)L��Bh�-�a�@�27��mn"�ĳFfW:�-�B%n�n�h8�.��V�450.U�!,]����j�l�����ɵ�\Cj��0P�b���f�9H�M.e �5kW���>U��*j�6ґڄ�Ka4[����2�A�cv�l�W8 �e��ec�4�������A�f�6c����eב�Ynlq��f� \��K�%3��P�Ff����׈it�&��0̻c��l�yΕ��I��-i,fף1X�`��ڡƺ���l��ĺ�h��M��(�	��I��]^2V���Fk�0�L�׈إɴ&�Z�0����9�(�^	
j2��8����:hᲖVہF�+�M���\�P�����#�4�!�B�Pn����]p4���h.!cs��Ii�(5nIb٩�f�F�j�v�-�$���ѹ8��S,���q^�\�"� �YL�9���鮅l��X���t2�f%,�CeLP�DC
�M�C(Ŷ,�U-�um�ŵK�.��R�mq��.t�+2�X9�4`c6\
V	r���ڥ���vQ��܌� �v�5a�#�B��jEX�����R]��S`�/hh����LvY.�w:�.��Kk���.c��\�͸rA��BS��-mM�-c��Q�;$�.4n�qL�R4M�a���%T�l�#�[Cum�`����P��j�+KYn���������Q�%Gm�.hʛmr��+)e�h�k3�ᣡ��Z��u[�a���<y�m�ȰrܠP��[J���3�::i�4NItQјD�f�5�]�Gb�6���m��A�%�l��� �p]
�з;�F��c[GM�5x�8MX	A��f����M�)��bk�\��VS�2�\PJ�:�v���v	���;5P��v���j�1�� lj�*�f4��3�k��e��k@Q�����ը%����
�=��\^�І#�GbAfi՛hQ�VR�ҥ�C ��
0�]�,.�C+�Yf��X�C���42MZ��a`5�I��� �c�ԙ���\V�g
ۙ���9�!T�Yi�iP�	@�0خ�n�lia)�M|�y �c����4o���ZV�6&I�����g3-���CcuPd��Klɵ8%S5k�I�[-��{X6�u�u9C[*U���Ƅ����H��3(!,������!�!iZ�+�fךE�jZ�W@ۂ�i�4�K(<=I�֭t�YjE�h͙MH�Z0�pme�
7a�dX]a-�&���]�0�5�tz��52�6���g0���	a��{-!-0�H��6٭@&�D��ѱ��m!�r/0�w�q�B�T�t��p����F01i��i���˝VkuQT��Յ��!�l�3m[b��&�ԩ)�^��	-u�f�i��Vl9�2���R1�Y��fq[&Jԕ���ofe �����Ca�7�L9��q ��hP�K�c��[��l����F2�����[�X\Ⲗ��sw�fW�Srm�R�$B���.��Ksz�p�P`����+�M	�fٮҐ��E,��pd,� K��Q�����5�m�Ş�< +h"�o�r^�T�7Z�P�M�c�1iŵ+[�]\�d��1H]�	F[x��q�At�Gy|�VS���J�4��/W<��:5�%�l.u��B�K.R��G]Z�ዶФ\JE+�af(��6hi�4�B˴���ƌ^�"�m���\��l��l��:�Ռ3��7`ЂR&�*�eR*&�l�SDŉ��6l��Mf%sZU�n��ٰ-nDV�L;-�P�*�:�p�60�2�%�A�4��@�f��h5%�731�2n0�����6�ܲ�Ֆ���؁pX ۮ��Ж�ֺ�V�Ò1Li4K�3&�-�QjL��^��h$i����3hƦ��M-B���6eZk1Rj*]k%-&��1SV*̙ΰDõ�N�h�R�j�ں,��t�)�r0�vfrv]�,�ķV,X�m�fX��h^%��]3�,�k.���]�h��.�%uԠ�ٍ.ctq�\KsT�嵸�w\'=ne+Xl��4[qn�Ќal��=��3���Օ2\���cR�m2J+)�-
A��!LRe�Z3JUZL�	���՚V�% S2h�7j:��+l3;[6�#�6��A�Y\�c,-�z�tuc5��䶖3Rh��$�st���yRY��6%� [[�˵\���ƃlfƻ��i��u���!5 ;��R妀\�l��NA�m��K�7l#�Q��ن�F�	�٠�q��7[6 -�<2R٥tqP�H�H���mΘ��f9(����؉e��T)L���s�����mD��ԂՅ4�[�.�f��.7lݻG����&̨%qv#6Ae����"S8���47Z��
B[��+�54Z����J0�2�b�Vi�tP�����f�ohۆ� �ns,K���Y�&D�n6&�Dl�X��$z��#�h����L�,����p6cj�1�7����&1p@�Q�[���!SM)���eKucM\��)n��Ys��hRb�����1#�����1\Zю`��L�Ba�^�TUͶ�D�d�kb�(��X5۩1P���K2�!�X�@	m���f�u��e�֎E�*FgM�늖;h�a*�]�5�+L�mD��"��/:c%pڶ�@y��ҝ\�����JJjUnTt����۩J��F���6����d4i�l��a��a6HfIk2"�U%�,�`#+�.�uV��P.K��\Pq��Z\���e��Ŵ�PQ�\6�DXcA��5]0˴�-ڭ��46���`#s�m�I�5b� ������`�q5�M�k�v�k��k\ʰ���&ȺkHZ�b)˜Xa�pqu{q����n���E�B��Z;h�AU\��Z������@1�������n�:�B5��ح���n���K
qb���]I��]���a4Bo&�X�c]���4԰ƽ�Du%*F2�(�Hn,���Cki2Օ���t�ƨf8����-�8I��є���F�)�P�56 e��1f,ԩ�tH:�-��R�u�Sd�A�-�1�v]���5s(�\v��f`���X1�� �#-�!z�.K��;X&mQcC̶�Ɉ��*B�4�\GL�J�k+�aW������h�@%�]��4D��.� ��sU��B��MU�1�018��+T����֤��6�c�s���6f�KUR#[f�ka�����+���a�U�����n-,c�#Z0��]&��](Y�-0�,����UڋF�&{�讪���dv��c\6�%!�$Xsi��D��&��e�Q5�T�[�<�%��h�X���f#��Si�q(�!�����6�F�����1�%	l�����f�Q6�ٔO/�����]rD*��N-M�8�LF3k^�\�����	��G	T�.�+��d�Vj�Q.X��.*@bfM5���lf�e*�%��K$+m�*J��T�b63k���\B�\k���h�X*B���j;1k[��R�N��H�]6Lᕖ���evnsJ�e Z�ܘ�b.�r�h�J�*�[Q,��j�/d����1�f�	��l	fsZ�A��eո,���ܹa!�u�6(�d��q�u���\!��L�̹]7k�Kuc+6�K�c�fF�9f{Z��|1�f4�(�-G;V��ͱ֕�Z1�X#6�\j�.h䆙���^&��2�Sf�6�.b�Sm��clkLWm�˴p�+�s�J��Z��\��Z�
�4h��E���F38�@�A�,]�-�q4j�
��ʻl�mc���@ate�����i�n`ڷ ]��Z����WV�l5�<b���*Ռ�,�]�Xႃ�pm.U�S�������h7b�)r�l���kS�J�+�#Y�.��F��gJ�Q��B6f`�ij��q�Y�u�Ԗ�胫k��U�Jd����l��+����h���P�iM3a�b�3B��G;:ܮʸPX]6v�f`�.U}��}E�'�l���t8�R�a%&XJaL!���[��|�c=܋��9N��G>W-~~�ڹ_�/wh���RS,���ru)j��i�[O�5��y�*卯���-r��f��S�RSj��X#-�V���ב��4h�����H^�qDl���͕:�m,�{�ĳ�w&$���XS����>|������.R|�+���~y�|����%�w|�~i��jR5B()���&sSM3)���P�E�a&1����K��5����6+Ϳ5x幾\�E�W-����*�b�����4U�5��Eʻ�I{�W��|����[y[�wh��yS�����$�m]�k�7��|߻�Ƽ��.Z湹�*�w���\�~���{��r�^U�p��t�W�V�wu�z����h�K�r����u�~��0X���
%b�bp$'�O/[�]� G�Չ�{M��h��D#����e��S�եR.�lą���e����[��)�V�Wg�-��V�Ԗ�Q�����4��۰=�5#ɩJKRb=[t3���f�A��Ħ����Qu�	��9	��YY��Q3��6ltt�SJ�)ZlF]��u�F��q�K��aJ�b�զ��7lZضÍ.��ּCS�eb���V*3&�ca�[V�Ia�XЫF8�a��Ѓ�]JT�G!�.��5�!�ۭ��m�MKh��cnZ��^ʵ�aZZ�tm3�Λ2�@i��kp­�&r�D6�`ʱ����t�ٱIf�e��!�:	1qy�:�[�9�+$e�qJ�/8Y�gL˘#�k���l�%�͋4��K�GF��T�V�h�6*ˋ���c��m��"3)��Af���\h�BU���m��N��Σ
[Iue(��l;t+�1����\�������gB���BĪ��k)�.��7���,�ɝp�H��=,i�L��܊�k�γi�a]&(����+lj���"۱�(���+�M���XĎ�(�҆�h����e���]n�kY^)���˔c�G!���\EMp\��4�LfC��:�+,��D%�0�ĵ�o0�; K��*S+f�-a�_ 7Ö�[�3A�sZƙ��T�������˪2�щR��if�:7kY�V4w�g��4ҩ6��u�-iPer*��ִ��]U�C+mvUy՛J�e�^Yk�V�(�Vm+qrl�#n�6��4��k����N��v�N��d�YZ/-��:Ѡ�o%���=R��-�6�),D��) *��E��m�X����BQ���V)[�QR�	A���[,�a �YK�R-�(1ZR=����Pj��ֵ[R�"�����~Efu�A���F��A̦�aEb���c��������;����޽O>g�3B�j[����eZ��<f5�i��i�x��f�J���{�E�ۋ�{�[���1�C��z�֞�-|��m|�ʬ?3^���;���_c�c@{Sh6�mz���O �s�љ�9�C��\�u��43���]m�Z�m|��6�o�C'h����N_\vt>�n�_���a�W�{��CK������H�j�
��ڳU���5k������in��Y��C;xV��D+V-4;�w76�m~���~w���3uRXsJə{ee�^2#����`���?+���[-���ܥS���B��J
?�]Hպ����>G�u����WUw\�|C�ک�8�,�jM�n�mS���1�����n�_ �O8ݍݝީ�g	����u��q�؎�c[���9���rӼ���\�@H��J���#���S	W#;��iNx:��W����nǷ_uGHUJ��J&h�34(�c��a�4Щ���Tm��J��V�#Ww~�tA�T�J��Z���ם����N��|�����A"�]o�sB=χ{n�^{��G�fǇ8�5�Vz���1Wex<�ݒđ�2�G����kz�q�!7Zs}n��Ϟ��V,CS"��Uۋ
�L�{k�����N5=q`tf�[�wnJz�(jě�d�Գ�����s| ƀ����I_,+}���y��$��2��{ӭյ�k&�����[��dn���ݡ'���eFD����n/;��$��/t��/��خ�����uVn�͑�j�v3Q	�L�k��U��͊	P�6����u}�%�(��K�]<��J��e�U����uO�@�RJE��+�����E�/+��J�ܭ~������k��S�p�k
�w��΍�BD$�.=�ST�Y�ۘ=1y���nO}"�I0	�V�c�:������������]<��K��=W�J�<�e<�F���0f�f,���/��d�ʅ*�Һ�+��kbl��Q�8I�3<֑)n�t�I �$�빷����c�꤮^(�n��kn�z������N�#���)e���5��W8�.s.��P�5U]���|�n�݃ܳwظ'q�?-"���^[�~��	��%�9�f����jq�7��pu�i.��ۯ���M��hvu�/�%	^��p��7��z�u�o��}�D$�"y��q��M`�n��x�Y�������l�+2VY�>5�+�ڤ@I+�$��B1]R��3Q��]1�ֽ����v����TW]a*��JY�-��D���t(�9������m�T�?qt�&+�dSj�Њ�u/��,l)vn��4�F�Q�jBQ�	��nJ"�Kk5���T)Tl��m����6n�1��A�q�yx�����ȵ!�9�+�U�eˣu�3�)	���G��C6g���y��'�(M��[6f���C�#e��"��;<K30d)\[�4#D��ah��cGf�2�ckns��v�]*��߿HM?mQ�k�1�]\����<�n�h�a*6.�ժ5t��w��ߢ�P�	.�KYn{�[�o�[Fj̅��wwl��͓���Wq�Afps��u1�N����}�REׇWn�G��[�{��BD$���8Sڜ�2��s��a�Z�%޼�o�I,I/���/�u��=�7�J����wV�V�y���u�5�:b�T����ݑ�Q������,J&g_iN����=�$���S�����
T(���]+&�ً6��F�t*m�B�WB�ꐥJ��ܒ�!"@�G���pu�%�A�����7�#�=�IR/z�ܼ=�ztMEs���@��*����m�����ڮT���"1�mDvMe̼X]�R�b��{��ܟc�٬v���Zn��b��]dV��>]��%	��<�u�K}��US��̞�|=�I+��
�!-(��]&��y8���3q{���u�%ޫ�^��[U�1�_n�%"D$�O�V��ܜ:n�͗׭ݷ���� ݀7wkվ����4?,F�#�-e���Y	W)J���ԙ�Ũ�;;��:t���ϹUT��޹�է�M�=���R!$�)��\4b��V��U�f����[���ZK��_n�=z4gV� �	$�$׶r۹Qp�c�z��P�Ͳl��0D���S�(�r�6vG�q�/To;MS��:O���j�tn�w�q��n�ˣv<J�J�Z0�ڡ��>�ϹUT��޹��H�Q8�:��l{"I$~L�z�=([�zK�u�����wwy3Qu�����z��A�m�f%j3j䱋-ɡ)��f�)����L���=(�v�݁�;����ۻk������V����|$���_���+�\����kz���v��o{۱�w`:�[uC{�H��	"�+u�w]�FQ͛�����U��۷��ݿQ��xQ}p�t{�N���t���m����ܗ�w�x�=�F����FEK�(���c���j�i�!�&qU�x�	�*��!�(k��\��.��T�	����C<��v] �{f�U;��^���/r�I@Ho�y��<OT��E*��Uh�$e`��1�-��ժ&��7wB�A*f�]����!$��7�)��u��3h��b+%�v��݌��D�S{>Nm�)������ގ����(fۧ���oI%	��2�&��ۮb��J"gy�'N��ؾ�)%	�/9�`��}��k�_�Dp�olOO:�]�7gP�S0r�p�jIRI$����V:�W�^�����v�Ny�]�^����32�Ӻ�x"M��n�i��\����.^�>���/fV��s���.��k\ͣj���1:�寝-S*�Ń(S���y���{v�l˦fj�qF��5`ɺ���pf-e0cF$�͘	%���a�VmX���`ǩ�vM�]����9s��@fԶ�b�!]���A�Lꃸ���eh�l]u˚L�&��b��aġ������0Ml�A��6�8+��Rf.~|��i~��li�v0*�[Eh�[���&���Ȋ��F��w�ǯ���n��煣S���o��̠�C^�.ޠ$���Xr�)�Fw-[��"b��$g���i.�Bw���,p��:�辑I+�:��^gJٱɖ��m[�������wwpd��)u*������;��w�޾������=R��U���%�$�"���m�w&b�I�/��֒�W�wcw����Ͽ���%����GG&�n��-<��T�i�r5�E�ZeF���}�5脒�EL��h�Wt��2Z�8�1�R�]�:˼��d��E1�{��+�Ȓq��
�uedƯ#U�|Y(Y�m]��VA�����Yߧk�{b��ұj�rl9.u��t�:���UN�[���H��/���
��
.���>�}$]��i�Zg��~�z���֒�]ǵ�����ݐ�״5��K=*9)��9g��Һ[�z�ݻ=2oȵ�2h�}"J�Mio���g �M��1-tjt��݀�wov�Wi=��Vk��O>�%���]�k�(����P#���l-s3���^�}�W��H���[Nq���uN��.Y˥�ȧ[}/��ݏn���^���.��|�H8\�j�|;u��j6�0���.�`n��wu/~�|}����#�N�Oe\�mOQ�PeI�D۵wbcf���u�t��p��!��Hc���v�,b��UJV�[�
�-H�V�!	�7t,�ҨlK��5w��&�M�T��7"�*[�1��E��؜J]�܍�6��z8 j�ʔ-;�*�!#�J��Ϊ:�v��dL�pvM�Qڔ
�q��X��Γ*uV�D�N�΢�o=��a�OPZ�	��V�\�nf��-�PfA(�{�C��̱N��� Gg[S\U��K�l���x�U4��%�I��-�zɽv��F�s� �:�h,ݧ��+/\:Q�P���PP�T�Y��f�e1t��J41�΋��ywf�'6)�U58�P��B�L\�ɜ��"�hw	��[��n)�M������!옜HjRl֪Hp�MW�>���f�����k/���t��w4�z�z�n�n#���i��g�Vn4����fwmuln'�G�5R�>�9«����?Ũ�4��ݓY�wc��eV]�-.OjU;x]�J���nl��S*����������z����7]f[�x���[���ڎ���%S�'1OM>Y�r���+�`��]�9l�ZB�B��:�wK��h��ڼUV�J�g�A��2����}D�m��a�ͮk�+��,"߿�	�FN�
�ꧬ-���#uX�)��D--���=e����	d��I�1$��;Sn��I;�߽�o-�ly���<��^�H�����	#zB�U%���y�n��~;�+{�7��+go,�N��:�`1ө�����N�kpkIII8$�P��nh6��6K�]���i���N途���IF�u���%1%:S���%J$�����%;��өI� 6���!z(��9�7,���n���qg�����,:��'qK��u���_������x`4�J�#b�t_5�ç��~k�v�>_/+��q�sc�߆���>�y���y�m��~��8����&e,c��k���{ǽ/1�y�T���9?v�������7R��a�.��1%3p���>�u{��7�o���$�"�6��*{���Gj}�P ���U7�z��u��}B<p�<D_�7�9���vƕ��>�47w>�N�F��I��'��t
An�B��J��8�������+����ϟtw�y��z�{^��d,�j���A�����1�)c��M�q���2��Ϡ�箅ؒ�֦��U.�N�m��3�1�U��¾-�̋ڠB੕֯Jt��.�/CV�aν��	>�A��s!�3���=x�p��@!d�����#�2��fH��66Q�H��εi��ݱq���%D]j�&�e�g5��s���s�Qd�@*�_6"ivjuc/�dU�#>�eW�����X��W��ҪL���֎�TGU���ѫ��+��7qE�ʂkB,��ǻ�~��\z���dY��D��C����گ��C�;�����^�$C�����!�D�}��l�"�ʢO/#A]�wfꪂ�V�h��fhU�u+�lQ�Ѻ(���f��3���Ȇ�W͡_*zqj'��ֱ2�${�D�>��̐N@ �F���t(����Vo6�J��N�e�AݏOG��i���[�ޡ@! ~�/��Y���ע���&ot�tkP�Q��r'�2=��Fd������.0FG�l{2C���9'8�&G	� v_]�5�j��F�|STCu@�Y�t(�ҷy1G����7�Uny��a�dT#��݊���>��#8��s�r^X�1-S�r�9g)�W.�s��7�>4�n�� �x:��K��tW���_=�ܩW%fI��>�-/�>	�ۻPRV�G!(�E�ns���-��%���"��F�V0n�Y��]v�ᥖnk"A��	����cl�U��2�65�Z�eQ�b�2��%"��6���&�sKe�����k{fQ��S9F�L7f��
��1�B���,ml�t;Fi�]`�40f�q���׹��"lMMn�D���偭㫔X����b%Z�;z����b@#�=�P ��&��6��q�@K���q�'�f����9{b|A���2	̉!�Eè����r����γl�9'6�&GvǤwH��<�s>�T��@����[TA�]��J{�������a�"���ۯ�t(��(�L����~_z������/Y�е�C�jP8>�D����5��j��uB8��n�[T-|��m+ۗ�"_dl>��k#�'�=#�D�p���ӆLɯYÛ��Aa��*��]���b�d,�Q�0���˛vfF\�2+�y��hC��ϗ�z���պ�90��S�|$9
���7X���|�ݪ���
,�~mQv��Wj	�sTaD�J�x-F��q;�R�"Vn�:��S��w��j.�o��_�N�)��L9֠%��ϣ�r$�B�W}���T#o$@Q�}�#��������=�sbک(Ž��Òsoq2<'�Q�z�B��[_7�6/w�Bݖ��I=� �Đr u�˔�Y٩��;�$f�)�Y�Br= �"�;�Y�j�?7B�dU֥~�X:�{=�u�Z��su�	t�τk�fE�=�|~����\��锪`�l�m*�rژj_˘ܥnj&��WuzЇ�Q? Ck�n�-������Nm�@�{U�ױت=7�$"�"H̙>����W��/��c�j�rn����s{x���Qr�7����z��j��B�;ʾ �_2,�[M�%��]k��^Py���t'��'ތ�{.��'�{Gb�+��3�"��R8$��(�9F
�%%_��l,���aε/��Ϡ�p$�D�|2<1���&�(��r���=�����gL� x�*OO9��YN��>3'ّl��B�}@�<��aOk���
�"��#W����t=w֔���/�<�R�h_#k��m��fb[�C0�]���]a���]i]��'5P��P,�~mVn5�з�aε.���U�m^��v�I�������Kj�Ƹ��E���O�����"5U��F'V�� p=�$�Y����hg�Qk�?�
�@�>�ڜQr�)���ҙ��N���H&ED_"_Pn�B!��ٮT.��jD�" �Dں�h-�rڀ�O�����=����.-Arc�T͋j��Dڪs���!!	l+��1TR�!�F�֑���H��c��_yt|?D�Mj�]j���kG1Y�i�噛ݗ^�V����N��L���wH��@>�I��+e��mi�t�����)|��T3d����vфnM���i���'�����C�޽_OW��MV�Vn��^@S#�v܍��=���b�!�Y�[_7YwhWŐ�ͪx�m#�z$�%�	�� � ȥ�w���Ψ_/��6���t<�t�˕��[L)�щյi��{bH�E��%�_�P�[�gu��e}��@k������^s&���E�^ԭ���=�Ϭ�_T�YKk�'�E�Yr�ȕ:0��ҵ���I���}g���dH#��'t��
����5��m�4BG���O{:���ޞ�C�Vܐb��L��JF�z��17���7�>y��t,,�ٳ:�8h��Z��fZ�1�4,���-r��B$����s�хcJ0bn��[5e4%��k(�n
:��QX�56ņ�)b8�)ti%��B�Q !��:f�����i3L[%��l�������2��1U%.�Ҏ!��n�`���c�x�$�j�m�6~|����M����%ڻ$��k���#�912Q.���2�^��\zFG���� �A�}�_no4�;�l&<��|Ȳ	m|�AB�9�ovϖG��Т���{�z�hs���Co2���=w��� wǹP!�(���أoy��q��Ǳ.�w����� D�(�C_"��]�	�l���m|�͡_�Lj�C��F'vզGOlH#,Wt�_��A ƨ����!�(���>�0��7���ؾ������IG�exO�d��E�y�	�d�TתbDUb�R�^)Fd6��iB#�Q%-��#s��=��w��zhz �گ>�3v%�1n�Ph��%m�8a��畸�eD֮�֪�Vk�ӎw)�k�[G�[�'�-��91`W�e֧J����ӧy�'�cd!� &gZ�Y�t���1W��H���p����ϧ��	�V�2�=��7i�����"|p����Ъ����B�?"t(��Ϧi8�ݯ���V���^�Hb���ǥG��>��>�(��16c���q�|���ȕ�Y���>;	8��6};�^)���j�Gu(Z��֪�5Pfm0�nD�:�q<�bwM�dp>��^�G��Y�|��<���f��U-�.ep�уe��,����T��i�3"���=����CϚH9�$dz=��R�{��z�!��Z{{Ĺ]1�
=gH�fG��>̉�����6g�a���z�s�w7b^�S�M_Y�zu
-�"�.��/��$B��@��_�-гJzw!ߛ���O��Б*�]S�q�)�s:��s_c8�K�_]_vQv{}��l�V�A2�S��~�6��5���:4��}�I��*�9�}ټ~��A��P,�~m|����a��qĂ0�<�n%M��m�v�/
"�B�P)�_�{U��Y��k��̂{�Z�n������f��w��,ߝ,\��3|��j�#��4og>�מ��?=}h[�]E�3	1W��L�F�0��L�i\�����K�AY����:Y�K�}��L�vb��L����4��p�[Tn��Ȋ���>AO��%bR�r��OP�ސAݏO�z�U�m�DL����EN(�3 O� �^Dz:N�\���Z��:��
��	�(����_���J{��{�d3�������'ѭ^9���]�v��	�/7���ILF���7a�dW��ܭ�Xf5�7��K%[�����.^�32�u��x��K(�X������94��_ySZ͌t�Z��j�ggᑞ��rR��_l�z�C6ؒ��7u�n�^ܙF�/���%J�z�����Mx�Q��ጮ�]\��Ns6���I����=~��@Nd,��kv��:�\�P޹G�Uv[G� �B��TAk�Cu�[_^o�#�uNwxu������Ծ7����{c��P�Ƞ��l
�����7B|s"A!� ���ܹ|�cUbi�ab;�K��BkU/Z��MD�u˫��7�\����EcV��w�\��_2Vصt��^ !Cu_<� ��A�,A�W�(�MmR�Y��χ������L�֪�v_NY��&�f�8fK~����.]�yI�2m�1_�+������|�нSl����чz�7���}>�j�n����e�}��w�i��"��d�����U��L�F>�H.=s���u�U`�X�6��,ňT�r�3p�+{i�b5G�X�5CU��tr����׮�pܾ���{ݲ^v�;�)t�J/��|�K�:ۗZĸM��&KkV;�����k�L�*e��7+fY}"��fM<�k����P�yVlYoi¶Y��;Ո+��W��K ���!eM�z�e,��־�*�wkUq%��X�$��N�>(��B���T��3$�-��f����ڇ�f[�����b�Ř�cзy;@ơ)�u3��!�̢
jr�eT���UF��`O\�:�r���x��1MY-�j�{I�K6�ݪɻ�p��lw(dk�Ꝿ\�%�v�*�y�*ѽLdT�V��Jl8�n�E�k#.]"&J���=K��y\����w��M��X��@�"�%"�!��[�'��䘚�F4�S�3�������_f4�̼}�V����o��[VEƊ��VeEͬ�u�;"v�ʩZ!�)Ne[R��(��{pֽ6���c��<��pjuUU��Y�r����ko��]��-��&6�]����jhvi�v���fe�\���Y�~��	��]�~�:����I%�M"����_��˟e�o����|�4WG��z����P$��N�1 :�N�^�1#T�>�JY��qbS��MC�mID�#\���˚wog���s�������!/7�&�m��sd��'qg�۳t���5�[�G���$�Ts�#r�~^F���^���_7��HlTZKz�c��v	�������U�����M}����w���-��M/ݷ1/u|������K���p5'+�˚���}�G�ys�q�A�R�Q���>�h�wv/���%���w��[ȼ�뼻����%]b�٬�$��"����������vt��aV�-�	q���V��)�����emzܧ�%�񸆕,#1	5��=n��2�ۘ�t1����Q�j;�kU�d���Xg:�mX���i	f�hČok�����%m�� b�E��j��6�j����'ܕ�$I��(U-H݌�Cd�0�t��Y�15�At�]i�K.%Ì+�H^-k.L":\���rWX�l�v�(�Sa�3��%����˫+�i����-L�P+
M�A�D���f�4Ŗ��q��Hb�X*�`����U�:�gQm�:�Q�[�skB���]l������Wl���lX4�(�A+C[FCSbc[hHДB#bH6�ݭ���ɌUX/7�uI��v�i���³K��XzU<��`M��6���K�4ʆ��P� �Y]���vv��[���u�0��f#^�@f�;M���DG+6m�
j��aeX��d�����vmkXl]�����,�0��c�R��E*Mb	����It���EQ�-����u� v	m�xk�G$�K	i�2�b�R2��vʷM��6T�V��P��%���n�Zk
�b[��&�*�Qcu����p[T��Y������ڮ-���,�)�ij$��H�ٺ1.I�%�4:�ts���XVB�R���(��S29v�D5�il��� ^(Bف��,Kˉ��.����T+��o2�»R��7�V�)PX;^t��x��n�yx����,n��k��R[\ZVM�i��2,�+X��`1˕��)!��g*�Ѡ��\�8����*A�!��輚��ZMe�L��]+�m�S&�.]�|�;��<�/5K!�a�gGh�K\�q�;��彥�YZ�l�X��Z�#X4��F4��nf��4h���l�0��rVcj��cs4[l���WA�kh�����Vd	����-�mhQ1�,FVf`�\M]�7g+aLWs�(%e�k �30�v����]�\�\E5�L���}���'���e�e�Ҫ�8�8��΄.��LL�@ˡ4��r������E�_Ƃ�{�w���{���\��"���ڏ3du>#2D�G��-�m�k��S�4�?{ʇT�V�T>-ι��	@�r'�2n<5�7Vbq�,]�E�RkV\֨)We�����X� <��wH���u��5�,f�b�KD�l�Z�8Dvu-�}���Hfp�|wc�3H@�S,�ڦB#.���t(�ڠ-Ȓ0��n�CN�1��D�Ow\k4�Ür1t�E��Ỉ�D�[��oh��C��`��1�&�2�0J�5�6z0���&J%�2��W���TI�3(O� �����p�Xg�"����<�����[TCt(�� �湔\b��ܾE�(ׇ�l3$&v��snR��bڥKU]��N�k�wT��Sj�own�)�R������ ^6|�^T-���X�I��o�<����mo���{$��=C	��)��T-	I��� �����k:��{\3�H)�n����@�ڤ��P����i ���p�AH,uL�RAH)���Z���qSyp���8�o�#����� �����R
_;`a �%0���R
n�H,-�$��0�&s�{��Ka��-���X˵ �,i �;@`�RHou$���}���{W�1\����,���
���(H)��o���x�RUJAH)7��i ����R���� ����i�d��B�q��j��i �l<�R9�{��ﺪߙ��H)��z�%2�y�B�
A``�ڐR
AM���RB�C	1�4�����n����z�cX�N��Yc���bPHD�)��Ms��O�Yђ�
���P�RAa\�ᄂ�SuJAH($� 	>�����f���|5��
C��o�;�/�k6�j���R
s��H,��L=�h`II
a�� ���$��H,����B�0%$��f���w��y)���
g��
Ap!�$�﹯}��_��s{��;T��JH)=�0$��½�ᄂ�SuK'��w�󜖐P))1��
Aa�T- �ꔂ�R
kT�m��ouH)���G�>��F(}�5�z�2>�C�Z�B����[�%�8�X��v�b/.���ِ�2��Տ�xxMγ�1��U[�<�>!Ă��i��2�y���`JH,
;V�R
AM�Ɋ ��B�
b Sm2�) ����U��d�=���=RAaZ��	&�ZH)�n�O��t���_6��<	�ހ{$�J�i �����C'w���{��P0j��P5���MT ֨k^o�pw�
Aa��- ��ǵ�w�����\�����FJH(RJO|�-	) ��څ����L�e$
JM�7���-����������ZOȦ�]!�P�R]�u!�sIQr�f�˙�_��:O_,�D�tXi ������i �����RA`m����w�k��{�y�=�
ot�a �c�{��;�
�B�
A`k5i �ߔqD���C	 �6�2��P����h`II���T���������AI�)���
A@�)=� |��,.�_6��<	�ހ>4H)���q�I+��0�Y�Ja��-����{�Q�����I��) ���a$JL=�B�
A`cui ���H)��C	3G(ƶW�*�ﾻ;{�������c%$���@ZAH,=��i �6�&�) �RRot�0�Aa��a�AH_����;w\���R
AN怴�͌���T-	) �6�Aa|߹��zk�~g�s�x�S{��$J��n�i �8w}�:���u��w����Sq3l��]�z���woM�7j�4+;�藚r��\R��W\k$�� $���H,��AO����
Ai�����X�
AC"JM��Xbow$�B��9���;����)=��^���r��=<ƹ����	!UPU$��S��- ��B��II
����XӬߞq���
����͠)Gv�"�@b�ۡj̆��Pﮅ�-���a �n�h����AH)7�3AH-!��0�S~�ϻ{�u�Ny���ڦz�I����{����]��R�jᄂ�X�Y2�H)7����
A`n�H-�$�=Ǖ�e���x
Aa�*�R
aۥ ��}�;�w��7�y�;
ot����L�n�i �0v�H,i ��@{X��w��RHs�$�@�ꔂ�P����ha%$�B�
LSuK%��
%&�@[�㽿Qӽ���|��Q�gG���H�3T��$���0�Y��L7����%$ꔂ��RAM�a �g�y<�3��n�i �3�ڐR
AO9@ZAH,7���ٿs\��;�u�Ny�@��K=d���$�����JH,7�1����sW�!�AI�
`v�d��H(���lyV�Xy�\$���H-�) �C�,$b2S�h^sX�6{��H,�R��}Ǽ;�~g�s�� ��A�%2�y���`JH,
;v�ƒ
ot1D���C	7�Ǘ�L�~y+֞�N���w�xWGY��e�QN�+y̸��,n���E��4��J�yfr#rX;	
��E���W������4r��5��d{Ji�V*P/��d	�fPͥ�h�����XBg�X��^�]�6�ӆ��m�F[�[,E疇[GF69$���kJ����f�dtQ�0W��:���V�q�-�c��9(��.�F�n��aqLb�Bh�cC9u��s�ja�����?.�SfT�k6��J�q�]sÜɝTD�~�Ow��o~׸���JMv��1RAa�T- ����R�l���II����<�xo���{����Aa��- �;���_;~@�R�R
AM�y`a ��B��JH,�) ���3�AH,7���`���w���AH)<��Q ��j�S~9���]kӞo�8��R�Y) �BJO|�- ���$���J������
����-����ú�Ä�����Rc�
Q��H)��P�4$����f	�`�Q�^��Wˎ�+i���7�D0�Y)����-	I�]�R�������R�i0�L�) ���|N��4��i ���\0�R`B��Y-��R
ot�0y�9��|���=�Aa��- �=*�j�H-�) ��Z��=�(��@�AH,5څ����<�RRAM�a �S)��P�RA`n�H) ��@g��~�o���5�R�v������������7�8��R�Y) �����II�{ۆ
L!L�,��H(�D�G���מ>��P�����
m
�aWU�v�aq1]�Jڴ
�61\��:O�Y>	:)��R�R
AO|�- �#%0���RAB�n�H,,��Ͻ�=��w�3�9�6�S{��$G��w�<��r�hJH,
�ڐX�AM��(��Z��H)��L�,��I ��@ZAH,>S��P��_��ÔBv]��#w8�U���PU���1�J��.RZ-�e���T6mD���ɵOu����a��H)>)��T�X�H(D� $����~_0����G�>�\$�U@�R�[`RAJ��	�Ja��-�>�-���{'�b�H) �yA�$Je0�j������wjA`X�AM��(��Z�ou$�s��]��{}s�s���ߺy����) ��JO|�-	) ���ᄂ�X�R
AH)�����Aa��- �;�z��(֠v�H/$����AfJa��-	) �L7t��1�o��ڭ���|�6�S{��$JL<�B�
A`cq�\���~) ��h��
AhC[�a �"07T���S{�-Ĕ�XQ��0�R`B��Y75�L��s�^�ͤ���5�w�|�:��+{�=�Aa��z8H)��� ����`a ���{�ZRAB��)�{�|Ǹ�;���ȨG:;R6�V�%���Y���u��d�M�\e~��N״H,�L<�B�0��X�R�H)���R��xQ���K�7s���>�	��RAC��s�k�^�k���P�RRAa^yp�AI��0=�R
A@�)7��
Aa��hp�RuJAn0) ��u�{�u���6�e ���L<�B�
A`v�H,3��vw���Fb���#��� |��)���Z"RA`W.Ԃ���AM��x��u�k<�� ��T- ��
`f�e���P����h`II��P���X�Y3RAH)�����3�r���V����̉�9b�#t�M�r�]��=z�p��ެ�O]�LV�)��KZܻ�{Q�ݓ1h�Q�������������Xk�
A`j�H-�
H)G��H,�%0�����P���R
ot�Ad߼�y~[�w�����q) �*r�H) �|�31D��!��0�S�{�}�V}��7�`v�H) ���- ����9�w�}�����*���R
y��i ����R���� ���ov0�L7�����g�R��e �9T�=�^k�g���μ��a�����a �S)��P���X�R
AH)���R�7��
;�m=�?�<��>��j�IVQ�{G��6Q�q�YN�F�(�r79�$��>Z����O�(CII�|�ZAI�)�����) ���`w��>�����z�p�Xk��
B��7�y|�q���U)�������H,��L9�B��JH,�)���S{�- �a��{�Z����;�^�����qH,��S��1� ��G��H�<��S����[�|D�FJH)9�h`II���	&��N�6�f�s���7��ZAH)����I����p�R�JAm�I7��0�L7����%$(a�� ��^�<�mts+g[��:���_�G�#v �(�,��a��-RA`r�H,i ��@cAH-!��0�S �L�,�d����5����c�x���
Aa�rᄂ���R�g�G� "݀�__6��g}�Vn?r�Xk��
A`j�H) $j=�)��֭�a�ӓ��E;D]�ٌ��ԍ��R_�x%�}d3B��WF�������{�R/���� �� e �ᒘ|yP�0��
�˥ ����bH,�2�ou@�RA`n�H,i ��@r�9�_����	ȟ}�G��-�g�Z����P#�
�����.��;��hñ��`ܺcm�Ԍ�����2*g)�\̵}�>}	��F9��X#O��z���U�'��nw��j)M�w-��>�E��fH��A�D�U�g�C�N����A=�.�%��5Ic�o��l��}���c1|��B�r�Ak�n�����<S�"�M;�?Y��x�v* �P�����f@�uc���Ü���m@�S�#��w�m���y���z�8���XО���/��Y�T-Р!*�ޗY>����t���%���l�=�$�*��~���ܳ��
]����hk&�Dc+v�7'��{��#����bVJ��vM�\֜j�<�&=�M�r^y����?	 +Wھ5��������'V/
�A�oR���j)���3v���7g��Rbn�A�#Ս�aZMk[[.��@3��Ř,��J�,�jn(�f�	q���He�fFۛ�Vj1����VY��U-�Y�ʹ�t.f�i�-+�6��V��"��5�s4�`��%r]�6�u�1���?B�e��яVcje��h!tC���Z7cF�Dʀ�Y���/ߡ�}^%��1�^��ơw��t��dp"��އ
N�d����(�IPE֪kY���Rr��;�+��Q�q��Ǡr޾�}]g�v7=�5��O*RkYs�7��ݖ:Jf�W�����^���C��}����{��f��F��QmQ�hG�P��I���>#2D�P���t������-^[��79p$�0|�|�C  �
 ��h���)�"�um>�tq��co�� � �>�n�w����w�j�H%F��%WaU�6�T�B����c�f�����o�|;߯�7Մ�����_���W'��:�^Q[����r$�TAk�m
-���y^�H���xi긝S|)>��h�U���Y+f�I�LI5:yq�"�@ٞ��J8R���V5}��s^�o��Mf�'ye��W��k^WIi&G���nD�!���z.�`y����؏��u�.:�Z:��q|��Vq#����Sך�e�s"H!/��7@Wź \�	�/�t)h �N|Ȣ	̉uK��9���c�k��}1[/���L��i��n�[TC? F`7p9����ɑ|����j�I2<A��TA�E����ګ}�%*���ϣ�e̬�a���L�W,�BcX8�{aHl����j�.������"NdI#�去�s�i�}"���4�\(�A�Cٟ�Y���n�Z+���=���Oll�w>�<�^�t-t�l�<A� �.�)�kOt_ܾDl�_F�g�!��h@��vo�B/�����+��(T�sd�,�\���]	��J���Bǹ�5���i���nі��.�CJy�����Ό�Hk����r�w[�@�&HKT����m>�K4k��vїpp�҉��2r#��`��qШ���0qO���iT�܏zd�m�xL���o�朥�E\�T���KՋTYZ�ۼ�U�C_����l��!�sxrr����y��b�r����ҫKY*�>Z����*��VO���U4�o�����7�<Yu]�%�Rs(�gd��w(��4��"��34��ռ�k��u7��,�C>';1G�{��=)��̥�{�Kt4��N���������93w����y&�N�
ᵘn�/z�s��;.�[��J^\Εxr���c	�A���v*鸯Rڭ���y�.Uִf����f���W �A*�Hd�K��,ܖ���nso�}�ә�5�yp�En�J��u���!�̩�S�9�)�+ M�Iºz�sP�uU��=�w1Gf��ˍ:��ҕ�X�5�u������nM���U�oNd\��/3]ut����ќ����k�r�ښ6Ny2gh��Y;Eu+�����dV���!�(��jWT�?@D�x�T�t��D��T����
UR�h����޺d������9n	�s]��κli�3��鍍���������_�w��7��#���%�ƣfX�mw9;�k�����w:�w=�����-A���\��I�������Q�%�,l[y���ۛ��f����r�S�PW;�U��W�F�P%O��<�7���!��W���	1st�#˘��b���3	�5�˭�XS�|5��'ZL��A�{AnD�!Kj�n��v��7P�5}M}��V�\KO5��� ���V�R�..σj|[�'�	̏Nd��w�S�4q�*�����5�k��l��$�_S_y�ȉW���h��Z��MՃT�5�b!��1ɰl-�is*ی���>��z�a=z��"q�O���/�֓ n�b�2��F�j��@��"�����:��,�A|�K���n�y�����{�y�B�Ѣs��( #�P �B�d ͨiQ����V�[��b��ӳ�z������P��?�
7�׋Tz��L���Cq�̑�B��l�'ZL� ��@��u�G+������sc���eS��:'*�fO�[;Q�W!�̱7q��FN�j�E��C�����3:=�HǞՉ�\��RkT\u�:�#��f����[M��i޺
�	�bH�Cu_6�zlJ>��ᬳv��g�E%!�3+�bħQ� *Iaku����?z����hNdOU'���z�뷃	H��p[o'��$Ȓ8@̩�dI�;�����D�	�r��hu���i28��$|܉���sy�Ix�g�܁'�Ct(��~k��%�)��ﻖM�9�y�u����&�w֬�Hc:8E��7#T�ّ=UϷ���[�n�(�@"�"&��Þ����F�G�7B�m|��Ci[����B9��p+�C���A=���_� �2/����sm5�d�U
�P��X�WhΣw�of`)8�����t@��XhV�*(V�
7tV�gK��`�J��ξu��S�t�;���6���J:4���6i����� *]�.�)�,�mɶ%mF����+f!)e&�%���-%�1P���Y�0��Y`�e͚�$.��_:�M�Z�
��(�i�A���2*Z�\:�(� @e���4
��mYZi�H�s��J���E	V�� {Mt6��+n[��������C��v��v�à���I����΋.WS.D�ES�$t���2,������-|-'z�m���1iQ$���+��G���;�K�U�
��K���8r�mc����A����$�AG&�X�˰5�>�Cs ��G�#�2�����ޗM.�92��[���g��y(����dI�$@�Zخ�h�� ��$�r<�UwJם���w�A2$�ٶ�]仼� D��n}�P ��G�2D�!S�Dh10�w�{�X��c9aS���U��f��8u���li�k�C2�4�6^�Q�Ѭ��	�13h&ƍ���γ���������̩��'7~���o\��dq�/��R��CA�-����g�� �ޖ*Md�흫$V
��P��d�ܺ��wo���|�{Q���P��l{���U��6k>iq�ַ+�j_� k�c�$lz�__�J���^��������\�+���A ��p�fFNĩ�ٶ�mo,ǌ5OZ�CH>6}��[�T�j��;��ӴMT1����f�^�6gd�8�5�����9fW�� A��/�Cg���mp�s:_bp�@}Yi���av�|'ّi�)5�.!�X�ژ�f�ʛ�[T�WZ}sJ*`&r�V��rQܼ�ˌH�*����>_����u�DxẢ
i�wv�T�X�b�HYכH��?Z���C_"���@��Z������r'-9|tbh�ii28��=-Ȑp�7z� �ukc��$�ͬ ���t.���OWW����U���v永��q����[�/I��[0ܛU'�S�E�g�z��꭭T'(UN$b�|�� '�Om��s���@�ڠA�W��Wͯ�A�ǚ����)�z��̊>̉�����T�S�=�}�����z�����7u�k�~�Ck=w��>Q�޽��z��� x�u
,��k|e�{�(�MW��Tn�4ۅ�ٱ4)P��˥�e��7)?yg�~:���s"|A��;��+m���^���3܋Yu��uo���!��n�B?6��Z���z7ǈ{��__woB���#�p��#��թ݂��r��N�k�Ck��7C��f�]Z�^�������4�}}�܉8|3"��$:0�kH�> �_Z�z�gJ���ٽ羯�TD��ǙE�+�T�u[�V�ʒ�;�yc�j����·���w��������T�|R��3w��c3�k���ٜq���x�{˼�]"|CS�"�ͪ ��
,�������ݰ��G)�7ˡRik��=G�A��s"H9�����y����_�o�� �s�Q�,2[��:#j��PJ6��ңWw��� �TAk�n���nFZs����V�H3�@m�75+9(�8���ڢ��_�&��բ��H(�8�6;]���=}��dHa�s�g���"C(�j�� � fC���D�Rƹ�T�NE��� ��(�� 7t���5�/��YG)�3$ft�>ڽ�;6L�;�-I��z�h�l� ��/'�8|#
-��Ք��������o�f������|�n�|Ct=�eSB���{�W�l`��{�h�`�~�ɪ��Q��ͣ%Ex3��ʫ:�����_+�ή��{�x}�e��L�mШ�a2�Sv�X5m��M4`�)6��/Ya0i�ݬf`n�c�J��Wm@f@w�k�ɯ3]Pq��S���Z-Q�ͭ1������B����5�ٌ���T��=N��.uH��Ҙ��]tT�R�&+]�RƱmB�if��eEα�CsZ�,�����&ԷG.nYh�c[��]�	)J�:����*k�����?{����MD�!�":S�����NB�����psd�/:_/�5����P �������u��mϛ�'�|�r���i3��=�ϰ��/������gW����[TA|;��hS�&:�a���f!�q��E�7B�-Т��M;Pz���ה��ϰ���dGuu��j�������ϣ�(v)Xɧؾ�L��|Cu@���<37��Zg��.8��η-�͆��>j�;��"�ͩ�;\�K�H��G�Z]c�A֘�h��M�b��D�t�Ve��~�g�C��_6��C��7�}G|:>�3���Ƹ�oi�X#���t+��
��A2=�8���gV)�Z������{F�KH��h9'Y�V���n�.˳�j��(���Q�y3	bgY۝�o���{�{۴,��D�����r��u9|$g�A�ّ؍��UL//�#ު�*3�!���B����[ݨ�{,_ikYA�$S�a�j�n�z���f��VР\TA|����ƏI\ע���=����#:c��_h�P��DڠAТ��7X*�`Ҷ$O;�׸�����]�Y��=�Ak���	s�������*�tI���3q���|	��BW3۳�K]*�g��/��?gz�s��{u���{,gikYD=}�5����e
<~�!�+�����k �.VtۏH=8��xt���z.�}y��@7��⟲Q��P�t�A�t(�������Թ��B��U�7�`���̪�7Xi�3.�2iKr-Ѩ��8�hU�q3J���P����y~{���������vۑw�M�@ �"ȀPk�С(e]߬n��_�_�
>�[�={O"ֲ;�{"Au�-<���u$Я���_6���~n��7Z�p�� �z3k�ce��oA���ƾ��������G_�~��i�Z"�F�c���]���v�܎b�-�a�ʢm�l���$Vϰ� �ȑ+�;i�w;MȻ�Ю|�����"A}A��́G2$�J�`�a�O�����tUv�ȷ�� �Ȓ9���BnY��f=�g�?�
�_�
�u\wy�}Fp�7͙�ngU,�JZ�q5�.:J}s�Ah]��3(P<@E�����w�gi�q�>�EK�	�[�Sbw�K�I0�6I7{dW(��Ε�5���t�nR��.ad�����0�+w��$�|��sʴNԡ5���M3BkY��k����}ꎟ+�Ή��Ty�;ǲ=>����נ}��>�_���!	���5(�h��Ml����ˣ�ށ��B}��׫ގc]�_���O��fz����R�x)*!��@�ye�kVX�*":�\g4lq�Ի݅�! A��)�um�|�r��wGA�(Fo˙�wt���s�ьԤ�.��ӑ�fL�2Z�����s��w���-�#�&�<�� ẢfH��
��������+"@#�g<]3��z*�}�����R���x�r.;�%"�Uh�V\t�W;w�2_y�bbb���3t܊�}g�F��d`!���{�����7��:f�x��%��>4�f�*Q�N��ﮫ/�O9�����.�a��'7Yw�̕�Z�������b^*ᝦ����S]u�E���ȶ^`;���ኜxiU�0�;u;x,9����gSC��L���n��]H2�Lѩ�Ӊ��h�����j�eGF�Wpf��H=��>&���8ei�{i�2��;ϑΥV�eiA�ep������va���oP�mɺ[:J����0�b�fX����`W�}�����]j:�Nq.�3�ٔ�eRIf�PQ��r�����hB��3p��Uf�Ub�gfE�Fy��WMbfn��&.�)��Y讍��s3*���F�)쮪��-��l�AN���
�Lϛ�LC�طX�`�t��hn��3��E�nLt��F�}KX����e�8[غ�'���Y����kԮ�@V�5M;NV���<�Y�Uc��[:��#��v9ך���ЦU����[�p>��N�Q^T;b�l��D�z�ۑ��9:&X�J��� ��TmT�m��+�N�5j�vj͇b�^�U�3]�%΢�n���)�Ϸ���Uj���.de��V�˭}��Y��	Y������G �h�ᕻV�0v-�k1�ޑrpQi�G�n�r���[��&I�f�|.IX��܄�~^l�ǫ��חM�n�BIs�9�����v���ï^q��	œ�B�	�Km��m���.ws���r#!WM�:s&L-������$�tn�J�c����O5Ћ�4˛�L�mҿw9�͘	��Dh�)�k�y�Rd)��rD�?wE|���)���R)�!@�I$N{�DJ��L��)!痃y�%���̚)r���_���Yue#��Ι��q�uL�4�e���inD�Y�.����iġ�[��[,0٨\!M�L�Z�Y�J��{Xf6�T���а�XG���[�A�!���5�`ئHfչ�{.�H����̂^�$�LL�Kl�txAt2CvK[��iu�
1]�/R��j�ѶR��^�q� ��c`Z�Un].�Vы&%�R:�a�[4�bk����v�3[�Eq)���ͣrB#,��t�:0����^W8�Ҙ�衁�� :�T%-�5���
�3C`)ssykq6bT����4��f��hX\�:M�]�y���b��2��6"g#3+n��p]CJ8K3��1[U,#aubµ�f�k�ԥ�6tHf�v�X�X��	�m�Wk�1�5je�fW�N�1�<�0�f2h���Z�
©mHe�JX1&�-�fkc�h�1�-j��3eĤ���jD\a���KpZZ�Xmq�vl�Ś�V�D*�b�$�J��\4�5%Y�1E�#P\���`bFњ�Ѯ���7��R��&eWⴖM���%u �n��8eb�Mu�:�@��B���: �cD3ui�c(nv�I�Gp���kCmr�*,�Cl¤�Έ k5��cA-#	����cx-Í�S�ôƐB�9�]�,�ZX4Ґ�H�\�R0K5��23U)k�`���˩�8$]�a�Q)pZ�Z���˶�{m ,�Քj��V�6�kIb���{D5��CMJ�u�]�`�q�w�y��V���iU�W0+.]���ҳEknV��Ӎ��X�E{4�uC[��	�Ʀ�����ݴr4G,v1��t�q�<�5k*���.#��;0-7a�JX(�ܰ�k..�[���Դ�kV�-ƚ*�R�0õ�EMWK����%]�e�AH�����W41TѥhR�ũyU�9���+s5���qk�qm�7k�!B1�Z�ʗ\ �$7d*0�X7qf`�c,V����3ci�e��}������4��$f��J�r�ң��P�R��ε5ݰ��A����D6�m �O>W�.9�����6)�\b�|�D���-��Ϩ����u�9�Z���Q�����WL��o^��A2$�z��������H��TAn� YNdZLw�W��i�M��7"��?"&�E�D�Ȇꁗ��<�vei����|Fd�={�0���GakQA<����6�����͡�~ْ$�A3w�6pI���^��霮����j�#W����5��oW)�ʚ5�Ȫ��:���Ĺ���Z�&�q��T�#s��>B��$��@�du��1>s7MH��"��x�N���WǢ�-|��[T��{�hV��~�dR�UZ���TԮ�řҫAˁ#_����¨OU웾���L[�/s���{��S���ﾏ+߮c�Kv������H �� "5�%���Cq�|+2D������	��Uͩ����W�	̉�G�e
��B�,�C݄��_^�
HG���YY��jE_	��@"Fl�4�(�y�^&A���РAmQ����{y;����w*y,ڮ���8M�H �P������4pz��|~D�VI��ꣵ��3valڔ؊,�+*��<��@�u�$��w�W�0��T���l7�E_	��E8���&�R�s�.:��!�֪�y��J��}�p:|E	�C���Dܵ"�� �g�3k�Ն�cϺ����̇*��ƾ��7WźO�ː�33�]o2O3�x������eP����|6&h4��V����+Y�s�O\��W6��"S�� �iZ��mf�v���� ���|��D�j�����c?Y�����.���W\]�`�Cŵ�©�[!��+��(�-� ��
���Ӯ�I�������z���R*�}g�;�(���_��kׂ����X��q��&p\�b��g�y��<��TE�%tL�.u������~u�>9�$�m��O,پ���8�����_/E�D���,��o(��2�Ԭ`1� ��������Y}�`��_6���|�!��G\X3��_B��m,�Y�����y������B� �>�A�ّ���̡ ��M �P ��F9�3$H�����[u�Z�#� �D��{.�]Iٺ����Uvz�Bn����*�;��Fh��rOq��
�]p���o��G���s|�|BC^veG�j���غb�E�އDň#�ț~�½g�M���Kj���Ck�n���Gm[j�ߣ��z��h�}�6fr��&��T�L�q�4���ʢm}Dx��@��B�d A-������=E�}"�n�:��� ��%lI#�Fd{2,�C��'���}�{ݵ=�r��H�_D��=�]�J܌Š��=��t�9�'�2=�ځ��K9V�[��½g�M��[T1|�&}�A� �%t�mWG���G9�1Ԇ:w���)H�����:����7��* ��n���_ Cu�o�=�L�O-j&ڽ�E���N=���@�ć��r��j�iR.��x�Wn,2�����&[D�/R�ڃ2�O�Z��s��s9x��78eÔ�eK:N��⪰!�é&z�Zۅ�.o#RSBW���z����͍�ym�����5	��f^*�$\m\\�j�&����SF�Xt4�����[oTA�j��n�1fʭ6�Y.i4Cc*�xm�f��lA1��.*
u{66]���f��� 0�4�%������҃�!�ƿ}���0��R2U�!���u6��f+5Q �A60�t���`~<~_5
������cY���^�M�4	zS���}x�@�t+��
,��ȟ�\#�lk��u���#��Ls�,OIJE�6} �"Ǎ�gN:��o)�����(����D7_W͡��,��F�w�R�ֶ.���Y�C ��Bs�"�>�.�|Jr^^l8�|�z�Q�Q�����|)���6��@m'B��ޯ����_2,��mP �B�d1�Β�f���c�Ϩ�������ّ�Y�[���S"銙1ʴ���%�;� V�Ev�v�q�K�k�L���׽{�{�D7U��v�v�+�Ƚ��d�����mP �=_B,�ڢ����#�`0r�����kVr�A��\\g�>��zqG��^�b�FU	Lmsn��K��;q2e�c\��&��붿 ��h)D���ܩ��_�q�VΐNdH����2��%�PW_iA9��7_2,�[H����ork���:k>���g��?";Wͯ�����Z������1|���|�
���6�zb���� �q$*;�+fs��1"|l� ��ٗ �>�Ȃ>9���X�<�7����Z�����k��-���u�n�eЫ3`c���ږōͦІe2�j/6L��bC�M���p�ov0~|��@E���{����v�P�𠽙/g
�8������C_ ChQmQ�B�ݳ'�CQ�'��{S��9�H�6�H!����s�Ȓ������C_c�G��=EZx���[ةd��hܭCq��;�9�5Ik���0��3U��Yݻ�iޝ���P��4l��~���sz�p�qoV��Wͯ����}_6���c��%�� �ș����y�0�E�H>6} ��"ͅ*F���I#��3 ImP ��7��v��
���ߜ��*;<�KH�A6�|A�8DNdg|���绣�z��G������2i��XbQ�t�&�5A���[�
�]�{�����\�Wŵ����[���[�z�e��e��w��Z�~!@?/��!AmP#m{<��]P�4" >���+ou�\��q�>�CP$�n��V"p���/���倆~���	!��n��o]��[�	->���(B��[U�!���$�W-�� ��������n�L�_]t�{����=~���d{V�8p,�ؾ|Ty��b��dO�q�B.z3�Z�Y��ں�1�dje�j2�T���J�jұ!���gxZ�O�ǰ�>̉ �H��Zyr"nOH�B�EΎ���[�el��Y�[�>9� �2=���uK��xA�uQ��uj���j`߭���[���H�Kv��ΰ���}�>�ʟfG�(���u�(I"8�n.�(y�0�u� ��
0��mP!��?")�Q���8�eB �z�K���3.�,} ��D�|���9s�@s3�E7�n�d_���/"M�0޿9����3<(�෨WŵD����Q��*�}��� F8��H�cr幯/����^j�']g+����P��Չ�YsO�7B�mK��"䖅���nV����W_=b��ŵ����Wź.��\���j0]gUݮ4zcmD�bru���wx-zi�D�m&^��dfK5ub��3*�%�efIM୊��x��g;"g�P��u����I
� h�4-����Kb�m��&�׋���6��6qĳD��3f�30޹Z,���j-��7��ѫ�1�cR	�&�3�Ë�[����Z [��3m����M��%�4���EsQ� �#\�I4��iXKY]�Lj�h��\�=�~q~��"~b�WZޱ�(��Rn��1�-�!Gm�����N������ �=,$��ջ�V���H{��%���(�r��Y�ꡭb�V&;���o^�s>!l���]��VpV�"8J����'|�I���O�� ���|����A�$Z�W[�{ƫ���x�ˏ#�fO��2}�P>.*�J�={��|G��dڡ�z&�y�s¶!��>�9T�����w!Ǡ3&}�A���\:�q3�n|q�k�H��j���D�|ȰA��D���ԓ���#3kk�f�-�y���Κ�ipjlQsg����~��k�k����N��W_9�
�Ǻ��ڲ_ F�}_6�@E�����H�.��<��i^d\X��.u��ߏx���5Y�b̲��9j����Z*���P���>�a'@�}���x	�>�� ��D����f�߄-���@�? F��mz�N�n쩐(�@���A�TAk�n�|�Y��g���SŹ$�;8n��G����B�d"/#ٗ ��C�d�Q�>��O�lO�-}��^���U��Ay����S�ҫ����c5.yۚLA��Z:Ֆ��b}�h�dO}ٛkxBP.�pϠS�'2$�G����l�^�ح��J] Y��R���lEu��Y�Uڕ2�'�~v��$���/&|}�"K�8�=ar)n�#�Y̗�v��B�Z�o�+����d72���Cm^D�4�F�:�����fz�-� �|�������B�
!Q���֨��R#�S�|gX4{��U�s�d|6��d�V�f�\
�:����Ȍ�UگOcK���Nۨ�t4k�<MG\#�wev��]P���%�ws���k��"4�z�lŴRZ/�^�����&��s}6AxĎ�fҖ��}x]n���J!�WO����k0_QE�f����i��N��7q���p,b�+��iu뙗R�Q��}{gp�m�:�͜��;�.V�t�c(KUb��&��Z&νu2ԥ�;�o���Ơ4�N�7���L)Sw'8�ĬDڤ^�V.��Op��l�,�8�h��;�u)X���%�����V�UGv���R��l��s)T�s�,�"ҫF��d�#pmd��Mν.A��e4�9�a�t��҇=B�a�pMd�W]���fA����%�p�{(�X��ffŖK*aKj	c3w�Gk1;�І�5x�qb"�Lͳ�+7�Qڙ׈UeH{h������V\[s:��%��QMH"�ܫ�""��:SR���e%Y���5��^����v��3)��Y�;��s�f�o:P��p`wv+�:rf���+�Ժۮ˷��R4���ؼ+ݗ�Ѽ�!)T��7�?O��l���诎����b]Cm���ױ�;��b�;�Y��:��+�J���K�v���}c�^����QX��J�QE�������9�]	@��A�\�LE&v�?��bk���f2��l�.�$��ݛy�@i)D!�ܮn�#C���dцBc�rFDbouv��vc�"�FC�SID �4��%��$�(K�v��:�A|�*F�Y�DJbF��3Ww##)S ��I2�ݒD$��p;��|��T̗�� �!����1QO�|���Þs�:�w߁��3��s/�܅����6�r���tq� �_�����_���3d�@��_Qw���Z5��Ⱦo>�K?"n���Y��hP��T��y�̷z�]t��mQ�����n���<�ֻM1R�cسXB���ir�A�v)q��ᕸa�5r�$�z�t ��}�P>̍�cRw�{��^w�f��et|~�ÑQ��!�(��������	���"J���3��GVj�;�֣��p��g�ڦ6�H�N�@ ��Qm}_5�͹�^t�Jm��~��_f����-�#����|[�@�	h��l������R$�}��gW9̽�6�j�����_Xf����r0�Q�e��5��$�ɺ��L��0�l7{ݻz��3��sP�$��F������D���d{20FG��6_�\�e����=�߸o��sa�\^ޡ_B ��[ڥ��xX��ش%�Q�df��d�Y�.Z�V��[��*�f�����a�/:[TAk������}���;�Wү��ui�/�j� 7B� "�x�g.7b�dG����GQ���1�-p�M�@!8�s0��
�b|UJ���s�U��&�r�Y��*���;y�%K�o3X\��դp �Q>!�	�� ��������|/5�~�A�E�z}��s��k�^+KFWO�"A��E�ysU_iU|~�B�!-���p�Z��-G�ۉݫ��y˄VH���>��fE�}��U&���A�U#J��1U��N�9wv{w�����;�L��btdH�eٛO�Qr��������'wy������.�c
�hp6d��C�e6��i%����2%[.��L7+eu�Ga���`%�&�����5����R�S�lSm�c���v�h̬Ho��<Ğ3FR�vt#c�[K4 �H�jՄ�&�qCP�4� ��\�ݜLa,ф��.l��f*��O��/*8[��H�F��nI���M-��b��T��#?$����Fd��̐J���ϐ^�5̈́x�(�yo_D���B��G���5�,c�Ro7�/��2m�*�g*P)�o�5�/v����A9����̦�P��ţ��S>D
6�H#2D��9��8�\ި�;��.9#O��<A�ͬ��7t:u�'ֱ�&A_z�>9�	���x��GV%� �� ���|Ãx;�o��U�֮�@�֬�28f����J���m���n�V'{�-� �|�n���Ұ+<��r����ņ>�ɳ��%q/=Y[�1���Ԑ���*�I���Ic�'�	̄�d�6�1�B���P���
9�@C_� ���٭c��_���F��,u?��yRI�~�\�W�PT��qj��κ�7�n��D.��te8" XS?��W�	ϧݰ'�#�sz��7�RĴ� �Q�}"A�5���ޚ��bw�X�eDu�-֪Ady�fn��TH�tf﹮s����<j����W͡@��������$���\���.9#7� �?����=�]z��!�TG����i�0����O��j�Ao9Vs���G� ���#��B ��e�#B�>?^�^�٣�\�5���XiQ�-�u�SDlf�*�lQf�]/O��qH��A�l��˚�-��bZQ�W^��J�t�ѯ�������E�Kk�^c��_���R����R�v��o��������{2 r�&�p�B��\���T5�\f�aF{��[�J���$��{�o�v��)K	TR�չ��a�Ý\j%̪���;h,F��}9��?��=�Y=Q�	�;�#����P�Y�[TCh!~��QP��'�=["K�G��m�\׶���Ŀ}@�cTayZ6�n+_BP��ݯ�ͪ �_2:��q����ތ��T����rFoO��<AND��t'����o�z�z������2��,�J+l��ynm��z�JUwj�Vj��s�3�������6S�7�[�iG9ܧ��VS��}B����_�
��Ȃ�z�6��D���"���tm��Z6�|�$8��m��Lq(����ʡG@�"��t(@@���|pv��+i�q<���oVg}����Yq֪^�RkWe�l�;��ԯVח|�@�k�n����l3�RԴ��Q��Q/����VT�8�N�h�u��,flCV�Y�M'����˄�I3C��,[��+�~>�^�u�TD{ښ�t�GZ��mVץ^��_!��?v�幛�K_L^#��n��Ю���Y�uE",]�Hp�a�6u�#�i-֘�4v�,2Ʈ_�����|�{�ȟD�JN7��H��!��íLq����ʐNd{k-%f���!l�>܁"+�:����q�lH>�in��Ӹ�����4e#���k"M�7g�nF��Mumn�Z6�|�'����>�+�����3����8�D��GiGd�}&2E�H ���[�r]���{U��ƅ���1��`�_n Ax��w��7a �{�(�Ȁ�����W{w�H��y��5�7��+�hkn��?i��xg��8�E�wFr�ysK�>x�v����Q���F�����0��FWZ��,T&�0�.���5�,ƅ�e�E\H��Ek6��,%	m65�4	�X�����,H/JĹ�7�m�Y�Y��:$J�\�A�W.���Ԣ�khGuf�u�kQ�\�ؚj1�$7K42�+�kI6�lf�h��h�[��m4p�Y��ߞ�'�1-%��F�%��-n�*�u-u����W&�_q�g�gK��[_3����?zw�T��D*����
+�Ԩ�_	,W����~��xw��c��" �Dġ�%_B��b�^�}��=�(ԃ�LrJ����A݉ ����z�B�]ӣv�����j[�N���X'{E���j�&�F+�7��} ��R'Ÿ�AP/:����7m-�'֣�)
:��E���(��_�?A��wީU���V�5��7&.B��p�>nD��D�0�'K��m\{HI!.�ѫIUݛF�Sl�!��2ͼ#��&�֛P��v�{~�o籲��qg�K�צV��}�[�u$��t�:k5+���%B�,�A�D6����6�\{������G�Y�X(�a�աg�q�^wkk�O�Wc5�A�g3��\ى̙��i�KJo���x��8�@�����v��KEoH>6��}Dfej���+�#�H>!	����|�iWRT�����7x�=��5�P �� ��[_P|�0{�3
� ��|Gr��t*��$�=���I- p7�$Z�薠��7�@,�&r��n�Y�Cu�k�b����;x�>���j���KElz�8�>�Ct+��
w�35r��eb4I
�H�u���F���&2���p��~�G��C�4=���V����#�������mC�z�<�����,���2Po{ӛ�WB|_H��w[ͭ��I!��A��l�M9v:�y��7V����M�m|���"��uڛ�*����H�#T�b溂�����FgU�+{&]�zoۚ)��o�ΒJ|em=Uv�7��1A����ëO��᷉h��H>6�O��#2=9�$��wSS�N�ڷ�VtYWH��D���ESav��5�P��H���{�Z�	�v(�}E����?�V� ɺ��[�E��!� ��Qw�P!�A-����o�}�<���iL6�S����fWe�+�İ�&Y�Y�����c�"m)��Z������Ƴ{���#{�\�]��h؉Ŗ� <E��Ϗ�$5��Ȓ
��%z7OGp��)D�آ*�]�U����u5�ӊ�ڳi�ޮX��V�%	�Yp���1Y��+��[�E��!�슈�!D3�8���}���vi"�j�'TH ���+o�r�ỉh���TG�-��V^,�c�U/:J���p�i�:�õx"+moΆ��8Q��ӽ�Ӵ*,^ĵ�C*�)DV�3Q���5�ˏ���M��Z&�e��{�[s��P.�V[�����o��!���Bw!_��dh��Mq���.����ҷj���fa5�e"(n7Z]�����z�O�����b#W�7B��I��d[��WMݽQ�嫵�y����P$2���������"��|�8n�X+zA+"O��f�����S� �`��cTm
2�%����=�g����7�|*��P?�D���X ����m�ơ��Df�����rr?c��T[�D [^G�I_^"�F���\Mj�D�j�]�������;��_��u��<j���"_P�?cr=��1u�a}��h�f��ohñDB7���x�T.�'N��.�f�N��0i��g���J�ֲ�=U7XC^���1��gob�(16J�]_<�o�+)<���9���
�N�lj�v�5YQi�l��-w$Xj5���t�Ak��x�jqX���ٷ2f��m�x�"�]S��)�q��>T���A�՝�#U4�p���MO�o3{s�����EK�ִ�Y*��^L���l�.&�D��=�7:�y"IrD�_v�Š��zKu)�ڮ�Lfn���)H��M9���z�[�귕Xp!���(^6����#[w�]I��Wi����ew����9��c�a��mVKĊ�T�Ȩy��[W��6�[�����P���֡�X��)���>�č�)+�ai�/o*����9�[��F��q��h�Ż��>������hѼ/��s'��J
�O��_d4�V�m�)΢����Sv㩔�!8ڣ�j��T�"�2�Dmmczȅw.��9��nz��J����ӡ�۹��&��V�gF9¸��ňl�C�SIѬ���Q��^�m�o9��Q7�6i�2݋s&66�a��J���V ��5ϯ�k:?���e�@L"�����t�s��2�H�mο�^�CI=�	�����K��K�r���Yy�y�I;��N�\2wu��T��p���.n&#��cb;���]0��r>[�fI@�a|�Ƅ�4���tc&a渤�۳{���u����M4�7wY(�#Qc=����w\�h������r�scE��w�p7���92�=t#ˬ�b�%��0DPb�.�]4��
�1!�{����4�{1�Dj�K�ѹ6M�y��qҶ,mj쑑���nt�]�1a�k���^u!-��H`�cNх�33[�H�E��ipD;m����t+sA�:20�uM���t�h�.:��z���Er,���е����&��E��<fAL�9
ظ�.֑Bb�U��m�6v4ٹ@ѹ�f�c��sR���[�#IGVݔu1��^c�՚1�H������p�6Ͱ����K�4.�[�XT�c�%`�hb�q�Ź�+��ZP��V6��$.Kf]R1��$.%�m%@���i��
8��d����q�Y�h�ڔ#I�-�Ɨ�*^[�X�p��f 6Z�F�¶f��mq�n�f{VP�f���4�a��H�b�b٩q)�Kl֎�S&4]`��vm�]2[j�Z4�%%�гv�Z�:�!AFQ�i�\h�QfiV�f�uZ��)6�5��4z릐�&u��7-4ٺ��p�
�;Z�����p�\��h�<��T]u��B�q��!l�r��C�� ���R�h�f���^�GK���0+��%��,g�q5�K�o!RZ�)Z!S@����,�	������R��C0w<�`V8�Zm��S�`�W_�h�)؍��`�Y���z��72�Ѳ�������2lYYS=Ky����W�l�k������p�-d�B.�t�,�Xy�r�Wl-#{Ya� �Hgh�[:�/,IMV�hj�`	]���F2��F,V�Z�3.p�ta���ɦ`)�vv��eLc#������(meB�*n�J�0��Ġ�2�͊L1հ��Jͦ�o�ӡ�<��UYIi�C�i�.դ�b�m�c�B$f�Ks:��d�b��<�s�nΚ ��[Ⱥ�R�gYm���e
�D֬]�[����V����Vl��4EH� <�;s���kĹ�@�e�8�++ZS3SXGQ@��X�V�#/4����6�:����~|�/鿆,v)��n�$[�Jƺ��ջK��r;B
����?�訃�B� "�>��볽��j��R�Xo��N�G�
3UC_"��|F3�+h�v�@��$�G���>��:��#�>7�> ���#WnD��,���<~@��
�@����K����Z2{��zD�`z���Q/�v'�fO��".�J;a^l{@��>�ّ=5�̷�癚��A���>�A��+���B!���_Qd n�ee\�zn�P�S�j��Σ�jx^G�@�C(Kj���y�[AP�I�"�6b�%f�ʳZ��5�1�rl��ߦ�=���ۛ_adr.{���%=��Pr	�*�]ի?x�F�Wź�L�|V�)�h�S�^�}��g��|s֠��k��
���TUH�I-61�h'[M��v�^�r����ۑ�c����ό���p���Aa!��2C���$p#���}���_6��]S�>��:���m�Ե<A �G�@��<~mP!��t��*c�`��(����5�=��>�3v�x� G��V2W���!u}9��e�@��ywc]����#�1�4��k�%����	@���(��K#ְ?v�e�%�Rtn���f���6�y��gc[u3-��ʓ��48�����"���+�5ߤ��.�������}������(�ͯ����-ұ4��	��#���t���=C��D�A�a�{-_g?_��>#�O8��?7B��ͩ;'W%��)��9��"��K�3ɞFo);b���@:�q}��e�5�#xwPF�y�4����AI^�� �
e�8���\��4�s�X�UpE�P����_���J <�Vd���KuSڊ�j{gUh�|o7���7��kWa����@����o�ߡt�۞�}S5`��A9����#�fG� Uw\A�T;��yO�M�5�1��Rh;-��i3WA��@�u��b���TC����kU1�^�j~��|�]o�u�ol�3��4�!���s#ή�`�8eO��ٟ�H���U=����#�A7�$�D�".[��e�ЍR�GJ���&�P-� ��߬��.n{��ϔ��&��ڠA��n���B�d G[��s-�Ť��/�گ9�3�s������Aw�`n�2荞���姆�k9MW4���ͻ�E³ ��M/jyJr����hlTc�q4e ���>���۫��_�P>9������_I�9��k�Y����ĵa�"A>�a�̎��5sř-��&֋uV���Rbc8KsM0J�	S`�n�\��z#�!�
�D�R������)��n�C/�H!S<e�i�Ad	�|Ct(D�k��uJ٧�X��e|A-�����s��C�<D!�!E��6��oc��>#\���	�eO� _8S�*š�]��mE1�j{��>}"�e	m|�B���cH�A�B�j�|p�����[�z�ƨ܉�I�[y��ۯ����� ��n����v.v�@9Q*�A�>�H��Ait��̏I�7z%�l���XV-}��ڡt��c�3���]u�ج#Ν9�ɘ�+��>W����콊�Μ��v����QIwB���GZ��f��H��� MB�k�;H)aW3[C0nÈE1KyYIX��q
JD΀B��A��Y�L8y�b��ݑE��i1�E�Fє�r4*�ř� ��- ���v ��X����hs��b��ƛ8�K5#0v�B6��3{M��.[����So_>�ϰBb��f�Mu"V��2[)���--�eQ*�]_	����B!��7B�n�T��������ʼ��iG�v���j�n��������=l^��	��$oks��rk�7�	�R/Pֲ�=ϗ����gkA�Q��j"���7B�g�k��	���U��;������	�#ޡE��@m���A�ҕ�� ��"#�_�PC��&�KW��f�}�����n��e�� �{U|m Ȳt(���\�65)�dE���S���YCT�܉>�#�fH��o��I6����Pb�4V�r�a��Uj.��oj��Y\U�\���=|��{�@#x�2$:����<�C�#zB������"�K�G� ȰChP-�"}�
�n�!tp�'�<��-�Zw��2�]הm,�.��#��^i�P���z�mN�wfc*�V!%.���0����|~�D�x�5O�q_KP��y}H��K\�t�^Ă:�@� [�_�|A,���R�xU�ӷպ��ɳ���������t(��9�u��O_A��B��}�x��a�w�]{�(�#�#��J�O�� ��ؠ~-� ��n����6=U>=���痽1W�ݚ�8�;�WŐ�%��7�>�i��?ho�]5 V%�#��a�+�F�5����Vj��ؾ��	��Fy|��_/Pq�V�9�^���	��xqkb �z<F�����
,�A-�#�����ձ�#�q.r�u1sτCP5p�i�_O�#M�<�5;vy9Pߕ7�Ќ�JZ���;�D��|.�V�p�M*3Xc0�ˊ��M��F��Vɬ�o=�ׯz
�g)���B�ޑ�<]����XG��j� w�P,��m|�}Cؔ������{k�y` ��^��{[��r��'�9P"G�[7�>8<r�O�����(� �ڢB�d1<I�f�����Q
|ܚ���j��|t�>�fFFG������P����n�����5/;�/���; 鱙m���Q~�JؐA�<3(O�d��k�6��xl׬�f�������"�t�~n$�2	��>X-�0���F�(��{jTt�@�
�/��fW�����f}*P�����_2,�k�����v�I���!���}�w�P-����Cw+�	�SR�\z�3�3$\����b�8Aƨ��&��yX1��,s�GrV4����ǩ����V�[��
�Sf��]5�u��w�X;�3���i��y�� �h�|B�ySZ͌t�GZ��ȟ���ѽ��Ӯ·��P��	y�/�������=�>��IR"U_,��&Jѽ�Y���LJ�Fk5��u��_"}!~�!���|[U�-���׻�.�7P� QJٮ��@�C���dY��X����쁸��A�{���n��f��N5@�H�0Ի�B�㖅�CِH�!��k���,J��:^��n��W��fG�fH}͊f�%�4�dH�ڙ��|"���p!��:;3�����!�����!|CuS|}��� c҅!�#�^�u�3^�|'"���(�Q��৽�R�&��嵲SH+�8&L���K��|����K6m8��uʸv�ބ���l�:����6�B�|>���4�k�����kXۢc2�"l5�2JLF�	ihۣ���.�l�SF6p�B
շ@f��a�sJ��e t\K@�]cm����L� ��mM�X���AL�[d�0�!rRiY��@&P%�B�����Zfєmn��g�m4��A]�\��`�L�O_gￔ�\Z�Q���*\�4�������al��s=bOv~K�|�ψ �2<�_3������C����[E�TO5wkVZi��U9X�.�:^E=���3\�D5.��B�-��z����ί���G�B��Wź@�;���	���[���Mz��P#��g�-��C�[�Y�A��F:u� ��KL��_3������ȑ��Y��$$N�.�O��$2���D�P!��}Jk����ƥ�.��@[�iG8�A8G�^E�'�������>%I��B�vs(��K���GrYB%U�TJ�WV��!���a��hH�]o�y}J5b{�N]���B9�Ak�!�	mP!� X��yki��y�[���1�ýʵlB3�T�
��!���)��vӡW3]��Rf+�WUs��W쏇�=��>lI� G�Ͼ���g��� �^D�	�g5+�s7�WB�#� ���m!��mf��m[�2�6ʯo�P؇����(�������+kۼ��l�\��p�!t�}�`V�g�3�F,C�ؒna���ܼb|��./��@�Fd�21)��4%��� C;�5��k��cT ��8���'�2Fѫ]
��E���ߒZ�����dyi3
�V�+���b�kD�9�j�J ��ĐCR �s"z��N�W>@[�+,�	w�]s�8�"nD��I"̟H>9� �Ó��}�DP!\ώ���qP�:Tb�0���yr�㗛k��%����G�P���j�̍�����ɔ���yqaD�u��>�zw7����ǖ6�a��~QnK�Ik��`���ʹ/3L{���k*ji,�4�����ϩK�QfQ��f:�Y�a�:N�n_,c��	�t��2�F��zM�Z�+3+R��J�\��UTa�T��{V��	�
(����<�3lU��긥`����XDe��Y��](�aP�i�����Uz�����׹�U��B�dŴ�����]0�e�3m�ܻR�,�/7�8�csc2q
�w)�U��*�����%�����e�U����ι�y(�Ke�Lq���)�[�Ýa̺Ćt뾸,T}���:n�KƊˇfk�D:�
�T���F��[�u.�y���M\��C���=74�U�������}8��)��n^t|���xCPc�}�˖Oi�vq���E[�U��ӛ�7.&�j-(���Y%��)��̍��bn�د/vo;5��k�F��a�W�Tc�+{�f��k�Z�ja�>E�h��r�5,�FP��mĪ�f���!�0tm�x[tm��'j�
8��j�q:�����ʡ܊�B�hQGH�x���]Nen�j��6�����]�lʤ�t�.
u��3��(3v�6���S��mM�9&��>ѥV	}f��J�)S:�e��fp�Ⱏ\A@?�{ۚΡ=�'����!E�m|�|�QIb7����{�X�ݮcc$JK79
�{�cL���ɑ36<��gݹ�-�ʹ=�fB��h�&C`6�H�f���)���)ݼ�-��&�g�sQ���v���s�\�I�cQEwsDU��m��Ƌr��`�*"2X��W���ܠ�u�_-��BEd����r�а�
 @��;޹�sN|�O�dߟ���z����֬�4�L���*kY<}�;(QQ��%������
]�M�A���QW2Z�LQ�TA,���j�#����������6��z��u�J�X� �����>#
 �ב�\��֬A�	H"U�j�Й"�Feu��u�[�t�Fl756\����B�)޴����,���#}��s|��	��mK�{�e��T1j��DO/��C? [_?1��ܳ!l�}�;hW.7k��P5uD!}�(���c9Z�:B7B�;��?B!��h$y���)�⽝����4�#���.&����ZkWs���0���hP;��̄�����{�wpMCǚ�G��i��>���M.�<Gk��qH�O7�UEEn\���-{dV�"�����ZJg��<��Z���$!z�=O=���l��CZ��kW���k[ϴn@�ЫAY����Z�װ<��a+F�q%�ρ>	n�Z���J�F�t
2�LK�<�hJ��4\U�������ɴ��u��ީ�K�7\��o:<��ffP�d�u���{�߇((��7O.��y�fn�Im6�o|+����'�V�xf{�.پȾ� �w�m~��noa�rmK�^@̂�.1o�%R�oz��`t/��7�]�a�A���zǬ��)b�$�#9�%������I��tiwQǹ-�(������W.�ᴕ����w�G�B�͎\}��dv���T^�$���}{��?�b@�<��\�-@�km	�[NKō��6�	L������m�v9h+%a(�!
�(��ݶ����k��$i�d��B��&�3me����V��H�h�:�*sne��	,Bź�[�ˬ�Z׭e�ٲ���Ԭz�u��$�(�,vIr)T�m������i��!5�2���y�c�CLL
ʮ	YHW[�V��+����ml�pw��=�+��|�1*����km�iV]r����5���8���JŽ����eh*n��_6���qZ�Ў���s����ݛ���A��m�5�V����m|7W͡�B�s���&��^Dd �NDXn��b�6�m�v��8��"���[o��:׳�dC|�i������G��wt��+.-�fL��B;u�d�.�B��ku�s�����;��ّ���ӻoS���sV�K��=�X�ի��_6�m�d�U;������<R�6�Z����X���WэZ��&k䷮�Y3J���J�V��L�Ã�\�����hV��?_t�{����{���jv{k<�fo��|�m��8u�WX�j�S��w�=�V�<2!�A��i��ni��5�>�[�6��3�}�����|;��]^q��{{��m|����)|����܍zr�0����a���p3 f#;ѽX��3�P�	�hMI�CA��.Wc����l-" �ƈ!�šb�������D��ղ�u�k��U��fN�a;qSB0W@nh6�iON�G��^���<d������6o��C�M�Y��5S�&��_6�n�B��Wl�56\�i)�7q�r�Z�6�١u�ݙ��3���t�5R$'�'{@�f`��U�լ�; pwb��Q]&�~�������;G�>6[�N@̏����޾/e^�Q�-h�t���y�fFdxffL�m�5T#��������l�}ؾ��k���giɊ��龤�;Q��a���E��DBP�L65�s���@8��Ƈ͡�b����=�zM�Y��\��q���������R������ȹI�p������^�ٕ��\�0��ր��p1@́�����uC�4���Yx�}�י�6o�ü�m|��y/A���C� �.b[�|x�|le�,�sy��6/+&e���NEe)�l�c�}�:�Y�h�U�tQ�;#�prQ�&���w��6���F�:4������}�]]�}�E�A�m�`����B��J&�b��E�.�23&��()�tκ.Z�UwWR}"k_6�m�'?wc�3۫WN*��Ѫ=����ds`�U�X/���.��a�}�zM�m{Pm�2��s�V�m|�ƾn��o�b��S}�U�{WWc��A��i����B�����|���}�μ�kپ�_���ux�ښ�M���=�%��۽�=��٘S��_�I�mkmׂ����IʥϪx��2z�S��y|���V�u7S����0�g���Y7X�����b�4߿��|PI�&\�� �p�6*R��[B��:��*�"X�i�-���j�Gf!.j��Wcb��5	L�YFl��4KsWhhB�=�(e�fn(�V8õ�Ij��L�B�D��7�����ÜX���
��6�h#e��Ep�xm���iJ���ņGd��nf�֍����X~stsfj;��Rj�ם�<�婡�5*:��vs�}��y��
Z��ck(r�\��1�U1���ͦ�k'qz˂�>_�M~�y<1�Z�p<�39qQQ�S2&���a�~�#�=��ļ�5ӂ���6������g��G�����g�^�2<c�]X�9�oz�v"��眾dM�a��b�a��pؓ������cX�pw�3=�jѐ�p[���0d�Jk4.�ճU�L�� �U���@��WIR������v���{�{�WG��/��	�6�@6�ߛ97z�b�웗/ٔ-D궾�t�\Is8d����;�_ˆ%���45���=�S68}= pk��>���꩝�����
FH��4���k�2 ��ʩ�Ig\�-����wFb�ڐ��el��g�Pƾ��%9�]�Mw�.�|1����Mߒ������́�{�o�����A]K9<���^@��@6[���۪�WJ��TBB�;q��5e�e���*h��al�}j�$j��?�r�>_6�lG�y�����7�T�H�;w��Wͷ6�ɜ���/��ʯw�^����h{[UJ��b�lL_V�� ���n��^�$�c�Z����N�x�9�!�x"�n#�Y����]X0����BV!��!�*T}F��r*�������ݭ}�*d�}�	ɴk�ИI�[���c{��hj{��zS��پ�Rۼ�U⾶��6�i�c6�%���b��Ɏ�m{ڗG�m{Pm|�vLʸ}����hR�v����{5�b���Q f�
]33r�y�z�w}{=z;2whL.����޾�bd��Xz%@Ǟ�������Wջcul@D����z\��پ�]���l�m�`n��M�����i���>���}ڗG����m|��)�y3.��M��w�Z�n��M<7ׯ�ҦN�7n�:n��ǁ x"�Mg0���z/gx��uu���[�+X{���PUsG;�3lU�]ة�+���7����M����O(󇝕����m-^�@w�h6��f�K��3=�*ZLƺ&ɛD2��WPu3p3�C;i���~��wϣף�mS�wu�3�j\���/��(k�z�M�����}}"���g+j���{f�9��O'o_x^@\�ѝ]xx�u���p33(f[订g��V�oSܭ��f���y����U�0J���Ou��y�{R����X��W�����<�ɴ_6��u{���&0J_�x�^�o:ܝ�k��6��Ü��C������[��3���w�����W�*�u3s.];A�9�*�ZsU�;�کbݩ��ʑ�ħ)V�Me��WM��{8Cj��O���|[��Õ��`l�k3h��9�kz�n�n�[�y�T����몒�X����mZq��"ކ���tʰ�ѫe%��-ٖ���y<��u�b�ڲM��l�nn�T��X���ߕ�L�.�.�CD��QpPǁ�r�T3�6\2�s&�lNJ��jۇS/D�]�͋�WR��U�b���2[�(L�F�T��ṱ��Cj�[W>�Uh]S��ʗW�3&�۶)�db�AP�Z����J0��9�ܙ���4�C�N'�s(�<�`�M��o#�io7.��i{g-����9&U�?^�Y�p�cV��5��}��M��F�]l;�ӱ�Yz��n%�N(�=�)�.r8/s%�'5�wU��l��X�͔f�7����G�s8�Y��&���^fmPs�����o��{M���Ձ���Zq3����N�ŏ9e�5�IJ�*;ӷ��F��.u��?�sh�]Bi�7,XT���L7g�\�����L���i�8����3i�*`�ר4���)L��n���5�t�{�g*��mbd^]ʃm�޸������ ��9yr�t2�"i�^��1�ΛRL�6���	,��M�]#m���wos�y�{��r�"��W������n~W�RX5����ݭ|�_-Ϛ頉�ێ�^}�k|�,W���>j���j�~k����my������E�}ۄ&���q��+�W���Z6}�ͣr�~k�������p���W��*J��B�s����W-�|��+b���_��ܷ�|��V6�Q~r�|�ɢ����ͮW�껺�.��@�wy�.����6�o5�F0�6M��F>k�:�*���y������6��ga����(]6B�m��9ձ�LA�h#\��[	��f�FZ0ֺ.�Ă�h�l�"D�l,�tڙĩXQ��$)u4�{$L��<t-C�[]Y��i���=�(�@p�W�Q.�3CJJ1���C@ضP�C���U��с.y���[f%�q�u�aRm۔���T�����ZC�b�][bVY��+4 �3�h�׈��i]��,��&Q,����*��'ha�Ż�K��]*"�4��/�Gd�6�u�m"�rԹP���v��;T6m؍u+s��-�hh�2�(E&f�gm�sWvteZM�6@YR�h��2#�A*kw2��ckf*:m��%c��mAƖ\e�1�4GB)��كb]�ٰ�8�ƶ���6�V,P���H{\�eC�5��U#��6Q����6���������-ڼ�ʺ-��&ƌpU�렛����&Y�n�H\5��/
E�a��l����Pc)-P�-�F��P���C�/����)3Z��.��\�����b	�^l�lֳU�*;PMz�	���2�iQ�T��Ͷ��)D6�	v�M��u���KhP�3�Kv���\�JWP(q5Zl���)�k�4&���K����b���II�m!�Y���F�����y֝��v�T��
˶\�Vf/We����Wd�ܐX$;�`s�6���#�x��e�*%�3q��b�qhm
 W�]���2��v�s1�T��.���A��U2F���je�riXc)�m�g1����Añ5vM[���j�Wlfffi�rK�s��Gf͝p671�5�1[XV5T�`^�F�驣2�e�4����tmm�lF޺������c������H�Ɠ8�vkmE�R!c7�	�fx�:�
��a�Z�������U�.�20pٗ6��Ճ��iq���C;��f��Ҁnf�,�$�A�5���1����0��i���g����t��t�� E�WGcE�᫳����fG�#����}�;m����ÓOz�\O�m|����]fvy{oP�S�dMwa�Fb���Q��t��=6���P�ffftʻ�Qɝe�֞J�|-��&�m��Էn%T*�o���G��칭m�\�t�9�S��������TQ�([B\�V�kz�y��� �{2��G�:�_�hyO߸�K/���l[.hdS$��߯;�|�4�r�مeU��P������~���7�[�O�ǯg��nN��ͽ�M�go����A��}��ޔ	��d])g�V�i��KT˴�/q�r]T��YB7.���z�B�}Y.��&�j�N,wx�vה�^�o��mj��<�f�"�3���n5nVdfG�&����k���]��ca�.��Z��ٙ�o��UzT,�{2���/g���'{�hGx�C��2��hm6�o2�SE���=�Bg+q�M�����n��}1���0L�C
RJ����Mf��A3Q��v�n�A]%J��� �|ݶ�����z��s{HkW*{�-_��m��}H����BCN�,-O�e���^'��rl���o}�d�E���s_6�_6��J�X�����Ț�v"�������ipWw�y�"ý-ި��m@��,7.��Y���"��h���-�Ŧ����.�̻�=!<A��f^U���%�6q]W�]�a�.��7�.�m8�_w ;�m6�m|��/s9m��Uf�uT������=�d{0P�1f�'����x�Ub�����K-�Y����5^��w���z�O^�3#f�����kU�"ulN���3�խ ���Ѻ�u���u>�y�xE��D;SrR�EI/�6�k�����d_t��i]C���VsNm�}y\c_6��εe��Z���_^���ʽi�]�p.3-�U�
��P8�,��N�Q��fq�A-�r-�m�iY����jix�P���2U_���M�y���!¯�����}�j��l<�װ�����9���n��TA4*��EXJ��41�`��[�]��RZ5Wf�]���~!�6�>s�޾O�������W�.��fe�����b�tSyB+Es麦�Z����sg���3L�ܿ�r�����h�=�ޜ�y�����6�m6�r.O�^RJ���r��������s��슕S���^�3W�b���i��'��j�kv�>�wm5�+��2��eI���k�x�$nq�i9�Щ"vҹ��kٺ�V�ڳ��#��y�gV*����}�W�y�=��Q��B�U�TnaR+a�����mcz��Y�.pƯ�2�t�q3��2�A�۴�Rm3��%�*��	\`\ʹЍ�����Em�f��4r��г	Ĥf�[ͻXཌZ�r�n�LP-����p�k-�uM΄�sEw�6��4�K����F0ʵ�cr\	Y��VZ���۱�؆�k)�pV�ḧ́�E�]��2�k�UaQWWv.����<�Pm ߗ����]��\���=��O
�{�m��}�l��J�U�jȁRC�z����z��2/�&��͏yԶ͏y|./j�6�A���E\��1�3x��v�Z��p@̏6�_�C졻��|�]�=w�1s{��G�==������i��I/���i����'�k�>�}�NA���z?z����4����n\͝Ƭ+�j�/[���l̵��j$��MK��<�d�]gZ-�[�i���5w�����{W��n�m��_���t'�6zք�����l��s����-�����7eb��P%qe�׬�`t�ڭ��3�2���s(�њ�ɯ����9�y��K�����K�-RW�_F�A�'M{�[��-��������2/����6ݺ@��i���K�d�y��ηv��\�4	ӻ��Ա1H������>��=^V�/_��jn.U}T�D<�W�Fe�c�ȹ�|A�6��6��6�tn]]F��L�#�;jv��$W;>�'��=�̀af�w\��/^'.x��b���M�`6��oED5�=y�������o��b�uY�s�0Z��1��ne��U1�U�]N�,h6�hm��{U,!oe}1�vF���~�O\>�g���1���j�lЫ8hy!4̪"�o��3n��.n{��õ�h7�Ƿm��h�{�����3ӳ{�"é'�}��޽n�� _6�i��ln��v�B��3v���.�{����ٔ30]�f��~�q�>|���+��kv!�ٯXǑ�b�Ѹ0m"TU*���`F�|ݶ��ܭ�]z��K��J�k|}k=���ڛM�_sXy��f:�`�J;��oaz�>��p35�ſYjj���������۾*�{�{�y}��b��m��K$oJ��փ�k�w+|r�}�K�g�Ʈ�%y��G�յv�������*���%s}EE��KC;�;d�3	��M�T�޹��^�2��}56�mۡ��q����b���+{�m��`p3#1�������2<ۙl�֛(ŭ���&:�8���0�s�S�f�����Y7\>}�{�3B�T����C� �m|�
u}焝��7�޹������P�g��Q��C�"�Z���32����g/!��̮X�^wxc@N@6�i�J��W�ؤ<���ȋIfۗζ�{o��z&��ٹ��.�{(��[��͠A�M|n�jz�V�/;9\;Y�^@K2�f�xV�X�&�*Y�j��Oy�	���߹�ۻ�qlT3�����z�U)����Z�]����ls��s:���D7RH�53F���C\Ch�1�CR[z�v�`��b�T�ڬGbY��cFkF;�b����)���^%n��&�ɉ�"˶�A4m"؛Bil���̧�m��K@n%�/9Y�S��dؗ6Һ)���G,v��
�[5f4��3�#0�Qs�j�7[)n+���>��M����AZ��3զ���Z�� ���\9�^}���-���9��t*�u�|?Djsu\���m|�m ��+�؇��7���;����gzb�|�s���(u.�;�m6�l5�W�GS��9����ﱠ7Sk���#�nDm\�ס۽U�hww\�μ�����Y�ݶ2���w&�m �n��*y�<�7 )X���u5)���p@m ��>U�
��YDsI�*�|�U�F��+b[)+�TQH�Wp��M��[�[��gKZ�(�Vr^6s�k��m	���>U<*=����j{��z6CI�.��STR�'�E�U��{U�:�����+�s]�R�Kݷ&��G=N5���Wb[�{�^���$���:�m��7���[�;�|��<�ͯ�M�Mm��;��w�;z�kzL�L_o��_6M�^ۿ$u�u��r�7���{Z��c_E�~���9����۶�ͽ[�Q���D
���;�\�����ɴ���=c7��Nmq����sf�1KR��[�
1���˝����2�ާ�wRR������������6�m6�����\_c^�;�,�{b��c_n���X��u!־|�m�b��м/�l�6U�)Q�L���Kn<�VU���]GV���׆]�Z�]��}|_[܁�im��,�Z��I��d�6Эw�[�{]���2��oR7ݛ��r�g����&LY/�N�dQo.κ�rJ�%9��{1��N�P�ǋ��n���s39>��K6WkN�^N��>ŋK��Cg.�}2��f�^7wv��{��8��U�J4��Wu
���
�̩�_dh��o�2_`�1,�ػE�=ؗKR�Vr��ƞ%]sOZ�Q��׶&&�W�썷+dK���n�Ʋah�:�j��R �\����)�*%���뿦c�ْ@��V���W-9�S.�#\Q%ι�m�ʬ�+'vnݞ?'��r<��Pj�����A]k�/e;��U��`v�彳\u���F�g^��2����r����p!Z;��.�+4-e�9�h�Q-�dee
��_!5�X*�v�#w�
PA˺�:S��X�L5L@��И�+v��7�,������>2S�-Ub�{����(n�Ԫ1��ݹbd�yӐ]����ǽNƳi�tld�փ�jeZ�[g�敚���������o�ӸԜɽKE/o��V�";��U[W���v��t��1UBȒ:�n��v���Ҡm��KB��e	-X~W����&׻�4r�������������Tl[������᯿v�o��6�=����{��mF�-��yt�~nm/ur�r~�ͼ�DE������s�}���_=��(��Ε�����m|�˜�so�����Be	mf��K��,�tni(>cEr���ݱ�I\����[Μ���hאk�*��\��j3�i�-;޾m�$oJ$�$��gyz�H�ҷ�%�wqd�J����ܤ�'Lw`:SƇH�<�)"I��h
L��2�ShR7Re.�IƳ��x٭�xS�Ӄàt�m��-����s��ך��E��EȽߞ�+����ݍ�s^U�S���'�\,E|��������)0���}�w�|���1�>��cSɴi�aVv^�dn�K�����e���IN��|6��1b�]O-�.�{��h�m7qA~ӵ46��V��&��l;��^G�Q����ܽ��M��iJ�XU(����J�Ԯ��<�����r�M��~�6/��m|�/�߯���I��>�
�[��{}�M�n�m`��?*�.+��>�+av��IN��|��̙�s]5W�v��D�m��A����[�k=~ػ#�����i���瞡�����@7']�W$���}�y6��1v�{�f媫V�Y�(�߮�y_��\��D^K&L>6dx�%��b�$4��O���]Y՜�ݫcv@6�o�iISɤ�����v�wRS�6���33��Jzo�EJnH��f�g�dEH&D�:3n�!�hm����a��d�꒣Wwy~y���_n���W,��T�o��݁$/����h6�m ���1�mWJX�g@�7]݊y-�v��yьkU/��\��`6�i���o�����C=�ݩ�gzbo������1<� �;��U��ӎ\_u(�{���ڦ�9�����������6����WVe����[6��^@�fF`�{� �z!o�2��uf{���T��| >��-}����:t�V��V�ث��҂�2�U�O+ec��� �s��u�UU��h�l\��Εc�)Rm��|�<���Yf�\쵅\�q�+����ͮ�3ln�)
�3ch���nqt�ej]��f;L�@�(K.��ԛ���y��ZY�L]vntIM�L�kM��[6����[h\2�J:W�%�Am�e��D]\X�V��hA�F�,n���o���]/i�JG,&�X�4�0�F�J�iU}j�$j��}��z݆�w��t�:�m��eKl*��p3#2dsf���k轵}O��{תvG��1���U�:��n�i��Q��\�אߤ���Y�����h�m_a���F��j��̀�l�ϧT�ͷ�۷�*y���gJ߽��A��{����N����u�V{תvG���M�ݭ7�߼�}��_���@��8�ite&q�ٛK�lG6X��9*ػ6������<�h�{���ӫۯ/�g��^Y2�l�b���͠BI�==��V��k�I�UN�%U1y�]Y�D����LcȠ(C�o�wM�_�d��:W�.˶�s���ҷk�GBrQ��E��};^m>q�ن��pY@&��Cbm6��ISg;�f���'�׹~���^��߃h}��_6�_7�v��N_�̯��W}�{V]:[��-��/6�{�������װ���X�A��!�{�Nr��	�o���M�����>,W�(L�ev����A��+p;d�JͰ�6�MF��V�j3#2t�u�N��F���q��+�uOY������6��7�l��%�]��o>�ի.�-�y˧Io�ar�Brm�a����Vץ](0�mU����L�%���U`��*�Y�i�����A_b�L\AYRܳ�!��˙�R��=\o��:�ɝ9������k�ǦQ�H����{�o�ev{թ�7�����ۭc5|���i��y�o�lt��t�zk����1�y6�o�^�YT �c���Pu�Ћ�-ъ+�Pv��ƕe,Yc0�F;�����O~��W23 c�69��-cͷ�h�t6*(�����6�M��:�5;Ϋګ*���	���Z�T[��29Fb� �)�����}56ݷʎ_������}{<1��,m�j�սH-��S�8��g�c��s��>|,y��;�F�[�woc=n�Qɚ��.�ܷe�Jv��N�͋�u%9�V�j5[J����C2d��fk����/�hsA�>m �o���&�<b'�ӫ���*-�gy�fd�������Ϟ��H �JڻX$�h�ػ9i��ɼ�%���ʆ���P������E��������^��}o}�zp��~_g/�M�5�w1Lt��+���{�Q�n�=�a��qKn��{�b�����Tѭ|�m ��~}*b�L�o���՝��c^�M��&b��%l��h{2������u����~W���Dh6�@6�k�м},�
rܰ�8=���V��;�v!�A���H���ǻ`bXU��;D\��գ"D���u���TTZ*杪�uUZ8���Nm'r���:^�l�ͺ����<U�Z\���;����BȏJ�� ]2cm	IqREiYkNv�Z	�l�����@��(˳,.͌`V2��¤����҄6m�=vɓI�F-������Kb�sRj�6��$B��(��m4�^�!�k V�\��X���ex������Ԏ4V�����R�f�q����1�LVA�e�&����VKk������޾�Y�^JU�);�U�/�{�����������Cm��Z���eJ@dN#�O)�wWj��X�^G��ft�T��O~��@�7`fG�,�k����Ps��S��N�b�� 6�멧�Ur����̎j�1M�r��y|/"��K�u��ΠdA��m �}�?J��>��7w�|��v��u��y�3#ْ���)n���V�슎��!��e�T�ź0� ��ٕ�*/cW;���&�����E���{�1����|���@6�m ��j�QD�XAK���gQ�S�sũI���������vt<;-[�,ѐc�]�v=t�^@.]��=��U��w+�w�����ھn���^L�U�ur�}���7���c0}�ю_73n����{�2�#ِ(���k����k+ِ3v�6-wt�y;�n/�W��� ��Pw!��A�>m��W�Ri���!\��y}�^@�ƾn����u�p�Q?*�j���IZ�5�-c�&�pRgP.X��K�7v*ͪ������|�m=���W��U�}<�EO׾�Y�4;�m6�O��x�wn���̔����[��|7�ɿ8���h6��C�۰v�xן�����G����U���TJ�F�fĸD�ijR��utsܪ�s;�7���5<G��ue��*�����ݭgc����m6��~z��v'��/}�o%Oo9�t�� ��S̿)���U�̏�4>m���4]�溸o;ܼ����1}�M��$���
��RB�ں4T#�ըK-̸,͡U�:5Q5F$EUU
�UNזG�̡��Xa�g��gc�}u���_,uؾm|���)�˰��gG��yV�Go9�u������圦�ؼT��G�#30�sP��n�.�N^Sz��	���n��rs������K����@6��{�ó��ֳ��5�N^�4��9Kgʫu�*or���?a�z�v��a��n�o�>brͿ��L�4e���5�ƥl��}v��w�m�k�*t�6�K��%�9�u��� >����篭�O�7��$)�B��M˲�钉E65Y�	f6Y�uF�Q�����>_f��_�:옳�����7�S�(m��}����mG���)�����t�a�O�{����s��X��Rxz����D��m|�hN\��t��7�e:��2<FdfG�#�|�5~�����ƽso��S���LY�nPz�-�w͠A�n�
�h�N��Y�m^[�=�3 ����?�����D���� ��mjڭ�_��v�� �~�*r@�!�@ 	A?�.����R��%�����~xQ�X`��6�)�Pi
�`�l�MY�$�`*J���$~�5�v����?3����$�X_��?�Y�g?fϾC˓���ٽc���\�t\88���vc|@�	�9;��w>>��0��}��O�NHH?��a%����\�m����?T�'���������d>�C�(��d�� ����a���
��I{���?�-(�����fG�?�V� ��_��D5��	�~��Q]���a��_�I��ТB�G�<a�.�X?}�Xd�� ��w��!�p�	̒�+?�]�7�a����x=?L�� �h�HW�k��>��/�i%��}h��\��(|����?�O��x~���������`e>? eI?8�*>��?|>5�	?��>��%��?,�<%A�O��}?3�t�!�$���?����$������!��~�B�O��|��y?o�=�I灐����?V�D@���$X?�}$�	 �����$O���I�h*O����W���O������54|�Tc�.X���#�|��HHc&jL���f� cÇ��4��:�9��rkT~�e�*��v`�<�K��� H�a�>���:���$ H����C������I�O����{������C��O���s�T~��3��{�O�����~��������&�>��c���"�����~�B�O�O�`3���������>�O��N� ��~�ɜ�̑�?l�h��B�o�_���@�F�C��`q����3tjy������2H@�	�Ys|>_��+��F'�r������Ψ"������2�P~�d��d	@'�D�������c�����~���� ��?}C=�}�}A�����I��Oα�|���	�2�9�}F���ܑN$c�H�