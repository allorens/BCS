BZh91AY&SY�-���E߀`qc���"� ����b@�                 �{m�ډUUUUMi��6�T[j������U��6iL��L�*-��سLX��*V`Y�$��kl 5EHE"�����kێJ�"Tٲh�����Vj��+Z-��j��(���j5��fk`(����M*��6Ŗ�Y"�L�z ѻ�V�����;Z�0� @ ;�*#�9�@8ٕprT]��p��U�K[SU��,���ͫKDA��-��խ�kl���f� � x4ڲɠ     �@�6�@:���lm���v�n۫Z���l�6��"�K��Oj�pt֢�m�]���k5������j�Iò�l]gjv�hl��v5m���fAlѫ�)JP���Q"�}����P��^(Q�K��oiZ�5@�=秮�
�A�Ǽ:ѥ��x�z4�o �ؐ.�m� om {��]4 4��ɩ-F��bbF�d��J��@pr��_m)&�[������{+ˋ�T 6�{��p�kwm�*���=� �%ϻ�GP��=H(�����(a{�Ϟ:�}�Ѵ��T�
D���T�(�|>�]�W�}�>�>�l���J���o'�7���Y}�z��E�*��R��燝 5�7^�]���'t�D����^�^�������J�EmZ����e[�Ҕ�(��<�ª����C�L�{�{���l�'{�݁"�={��t���<]��u���.��y(�'w��4�;��UP�.y=� �^����S,�0��[5Tҫ}�)R�� ���]������֗:�445h��i{��P; ��A z�m��AC�"�m��46Ɣo�JIR����P����m��ւ�� hݻ�  i؃ Sf]s�4�`r �;��KG��6��.ڕҥ��3Yk4�M[ϥ)JP|
 |�NP g�:h�cՀt9��Dn��|� ;/����H�t�@ �wS��7 �*��bua[dM32�Ԫ�x;� >��� �;��t �0��3�� �g��x�M:w �n�c�E�� k�\mj��,�f��2�&�>�J���(���l ��}ǀ�[^�ۡ�w�s��cח� ��a@k� �w�nށ��          ���*Q      ��ST  �  &FS�d�*      S�MRUz&�&&��%"2�� 2h� �  $��ҒI�MSښh�mL���2a����%W߭~�����s�^X�_���_�[����<`-Q繩�}�]��h9�E[US�~�DAW�~�����j�耈*��
�I'��U���EO�
/?��}���m�����0?&'���h#�4Ƙ���ٶ�������Ķ�m�l�F���al-��-���m[c���[cl-���alm������a��-���al-�����[M���a�6���al�-�0���[�[ah�6���alm���6��Sal-�l-���[�[6�Lalcm6���alm���i��������[��l4��[al-�l-���l-���al-���nB�-���al-�����L���ǌ-�����[1���[�[-���-��������[`[al-���l-��L-�������[
alm������al-�M��al-�l-��h�cl-���6��l�-�����[cl�[alc�6���6�l-���cl-��h�4��[al�6���M��[a���[�[8��Scl-���6��F�-�l-���6�1�Ͱ�q���cl-�������[al-�����[m�0����-�����[��al4��[al-���h���q������al����[e����[-�e��6��[al-����alm���`[f�i�S-��[a���[m����al-����ݴ�a�6��l-�����[��cl-��[cl-���[��[clm�����i���������a�[alm���6���al�clm����[2��a�q���6��m���:clK`[f��8�0�T�-�6�m�� �m���[`���)lT�!LF�#l�
[ 0ءlD� �-�`�Jb%��lA� �-�6�b��0؉lT� �6�K`-�R؉l�b%0؉lA� �m���`%���؃lD�"q���`�F؆؁l�
b-�R؃lT�
[-���`���#lA� �-���cl�"[-�<b�R؉l� m�[-��`�R؃l�"�8Ķ �-���b��ةl�,b��@�*[m���[`!lQ�Sb%��)l� m���Kb%�؏��	l�"[-���K`���	Lm���Kb��S��[-��Kb%�`1�6�Kb��RءlP�([-���4�`��B�)��-���bb��K`&��"[-���`%�؉l�*[4Ķ"[-��b%�ةl�[-����؉lP�"[-���b�؃l���4�K`��؉l� �-�F)l�
[-���Kb%�B؃l�ءl@�*i���`��	l�([ �V�)lP�"[-���b���)l�-���M1�)l� �-���`�6�b���lT�*[-���M0� � m��`l� �-�6�8�b�1R�)l� �m���K`F
�m����m�6�[b��`���+lQ��m����[`�lD�(�B�([1 �"���(��l�(��CL-��D�"i��Kb�lE6�F�$`�lm���@��x�bL@-���� [`!�!l)���� [m���[`�� �[`!lA-��`6�m�:`L -���� [v�`-�@� b!l-�&�hV؀[v�ثl-����m���LP-�� �"�v�� ��CLQ-��m��6�Al1-��-��6Ķ%���F[������#b[clm�l���-����-��Ķ6����q���������0�1�6�������6�����2������c�[����M�Ķ.ض�2���6�ؖ�d`[b[`[m�0-���6��6��%�-��-�l8�`S`[`[cl�`[bX���0�4������q���6���ؖ�����b[l-�l0-�la�[��lcl-�l6�al1-��-�lm�alJclm�lclx�cLK`[clm�lm���-��-�lclKe0����-��ČK`[������`[cl��6����`[���Lm�l`[���Lm�lm��-�cli�lb[��8����6�����Ƙ�����1�1�%��6�l-�l0-�lKf���-�lx��<e1���%��-�clKclcl8�������m���clcl�`[1�6���lm�l1�%���Kclm����1�6�؛cl`Sm6���8ĶF���:�jT}�@m�'N	����S��L��je	1��o��[�ζ��/eT+�����Vm]���f�s���!���j�15+�N�C	���"�K�Yo�c�m��2�'�3o��(3l���s�ަr�ۧ�e��ʭ���ޥ�t��۽G�QM�g1M5�n��{��-ݳ���=`b":6�Բ����]��qzWė��"����(�8-^Yb�uڊ�eb�i����v1c4)�yVHH�*z�6���b�e�аIE�Mk�5�
pe��f��ܶ�c�0fTͳ�-��S��2P�s\������T��@V͏5�Nef��{��"�T������I]՚C]:rf��(B&��J��������52�-����+��#R��2lU��*�i��2��g(JrὪV��x�7��Ғ��!���� �+Yv��o%U<�S��w���i�r��P��-[�^�u��ָJ�n�[&[��4
²[ק.)��h�vCV]�.�ɘ�h���j���$i��;�g+Y�Ћ�M��+1چ�Ud��2�] �F�6�Q�j�ܕ��iH�m^k���v��]�SDn:b��(ЇVC#�̸������0��V3Ma��ZZ��~U+a5���8�eKs["n�[��DX�^Խ���ܕ���Ч��e�{�0��b��5�#2�$�y{��m�K)�3��X�Z��2"��-���3�*�۹�J��U{"�D�[g
^|~�M�H���Z,�fΤ|�(]fJJ�[�ͩ��k�h�-L��
�#-lu�ߛ*5n ��l���r��0�T�)�7N��@v�C_Rl��X_^�ZR֮9�"�+P��m��GoM�/)cJXS`9y!�G�T*�C�����լ/�kt�}�Ϊԣ̳�"ޤ�<�VFh�F��n�Y���o��Il�Z2-�[�f$�hG$���bY��,�p^SFN尰�-���Vɑ���c�u�Y��)B�ǹ���oi[(��*�f	���SJ"��*�j8�V�V�ed����m��I��gM�hw�[&��B!�\('g5�چ��CRb�îV�SR��%��aN!U呥V勵�HeaC,,�Ӑ,�I/`�u`��Ljw[@b�q6�)�lc�7x����Ć!Y��V�ݫ��jF ���2�i�"��ؔ��fUG�K w�3m�J������r ���HF;�!��ڤh;��SvΘ�ŀ����&	[U*�z�\�kw�Ln���$Jwt��V��T�f��̼�k�'eU�T�&L-]ַ�����#�0�,�Bm#�Q'V�P�l���f����4b��n��ɫ/C.ՓCd���B�p�7g9;ө�V0h�旂�5���:��{�0��.:�V�u��͛�m����b�UyZ^�چ�'b%NZxtUd�V�۔[���-h4�b�N�d�`�^E�n�t�t\�#�y�1�V<ur����;f+�寞���lآ�(�Iu�\�����2[r��t,\�	���:/�rX��憌4Fh7 y/#���Ѥ�T��l��"3v�F�r�FQ��0*�7*c��WxE�����	+.R4��X��F`ɐ�H*NZyQ�X.�Xՙ,6�m�«)˻JL�R�>T��}�GV23Y,f�f��)'�o�$>�X1�+��Ո�H�(�3sj,��*��Ū&�;����˖2�ĝ�Q�Ǝ㷬1�e��#�XkK]YH�����I-N��1+7^,�	��g����(��3����2k��0��͊�8�sC��e@��7���3v��9gf�;���gQ
�
V��馑tLM-�f�K�Oe�ck��=��U�P�𳕻A����xҳ���c&EoB�j�U\�3�m����A���i�i�J�IPz�j&wM�ii�HsI�����~�{�X�ʽuPQ�T)��p�-B6$A)4ʧ-�	�ձl:���bc�r���uMBJ���%u��G15�ݴ�$�I�ԂF!O^��Yy>�Уi+R�����v�����ig3xw5G�<�z���"霷m�E���=Ke�˔��lk�5�̻,gW�n�Ϋ�^Am����6���M���t�)Fc1�f��z6ԋK�v�3D
v�C�bdR6wj啉�*����d��Э^�5�o"�N��i���hj��c��S���:{F���<�ɕ*L9��^ҭrK��SN$&�ڪ$,�3#{e�"�I�n^���)3UKkj�!��/K��k^ރ6J�-��j��aLf^\�j�.�����Q��CM�mދU���Mhx�䍉���2�	Z�p��bމR��$&i��[�oe����ZGN�V�5���]�a�Λ�I�uX��4Ղ����ֺ�\鿛�j�Q�E̼ԦV�!���6������<�ip�XH���<0���dQ;77i�$�,�J�6����@��4͓,SxZ���hn�&��,zm��UiY4�X�7���IL+vu���\-+���J��]�b}�!��fI�*�%��Z�k6Y�m�z��ޭ׆��%��tj��؋A���~�WZ~�A���	Z��
�jF�6�DVPb�ʒb�P�t3�m�<`�V��Su�4��)�ʸ]����@��ۦ�HFY�Q��T�*o��4lf�췹�gp�U*��x�Ƕ�1ZNnEk7`[R�;�U�{�C$:ի������ie���qܷ�/X�j�ږv�,̗�Ӫ,�ղ֔�i+T�.��:�z-�h�2e�4Vb9U��PaR�$X�,�m�5��-�Y�.�Qk5}�V��{�������眝��vl���«�g��tF�ꌴ�L���rbu�f���YP%��G���!���aX� �ٗ5:��[�sV�
�L�`+�F�{�l��%���m0��U�9Vs���'��'4���^4U$�Wb�� �ce�[Wah:��7��J@���`GU�D��O\�]��L#/ �Y���]k��@��-�w4^����:�]7kp�לx�u݀`��Ú
C���k)�kKUsyׁ�H�]�V�>oi�J�VM��h�I����r�[y	�XW+�v���aMU��Tq�7L����V�nަ�=��y���+�t:��E�T8���{�=,�d��.���Qַח�m͡h�
��U[�F����޽6[;n�^!eAut�K�Be�����1n����>���XZy���jhuZ��'R5���k��Kʆ����3.�%YYŪ�fa۴�r��cs4՗29{v���Q`��d�j�L�Ԍ�e'"�2;��N���bIt���x駠�nޝu�Ǭ�/5��i]m�X�%^6��t]fѡ)�Je���Z�#��0�'ո�E��Uncj�ې[��1��^�m]���B詠����,�.S96$!�9w#�{�=ɩ��J+1�� �͖�F�o{��|��[�8y6�~6&m����$�n�R�Y<��E���M�&^S9����!��1�`��)J<Gr�v,��q��"�9�$K�V*��w��\q�ʾ�)����r���V�]ǚ�z�BV��2�4����j�6�j� �z���:��r}z�Y&K��[�j���j����kUdV��S̉[��(H�\lYĉ�Bc;�MnM����x�e1}����yANr�3��a�gUw5���4$iD�������h�a84γ���0�ci6���7.l�"��E��yG���R�j�۹��W/Aěur�B�A+gvݻĄЮ�Yx��g+D�TCBq�.��CJ�3cKy��c˥�2b���b�˘݃���	.���fh�|��q߭Ӭ�Ī�,]�����+�y@]Y�(��o���X��Ғ��x�3m��rih�k%a�k���
P�ҷNdM	��l�(6�!��4/X�x����ӵ��qM�-S�i�:��I�1�����1{Z���١�b���M��R���J�g�Zդ�ʱ%0�O��oi1������ą�&�cz{X0�-�f�X-���n8��S6ԙ�l�[N�ӊ�.jqጵL��.֛����C���ʢ�`֖ZA��{⨂�P���T&re�Y�k#ҖK� �j�JD�L����Ȅ��=�y��$�CW�:[��n��VV}WZ�
��݀�-�~�"Д��j��q�6�7{s�&,���Ǵ�PJ�0���Y�E��2�����V�7d�tcyq�N!d�#���#2�^��K�����X�,)�z$��/e�'� �vl�N�ݸ*Q�ʲTl��2�Z.:SEI�����4�U�n\r�J9BIC5j�1���{y/)���vTSf��m�Ar����z�3w�cQ��-+.M7,��-m"YF���d����v�K�-z�ts=XX|PE�� ;�u�;�Α׈��oF��X��B�e�N蕥3�ֳBܘ3(��!9-�om c)hܥJ-�lTYq�������HdF<X����e��G(\j�R��7G��ct\����-�Odugl^%��%�u�f��%�����׎�i�ٙr]�$�RZ�Pf�!&*��Wh$4S����W+U7M^;�C#y<��91���]�)mQ�mV���j�`���v�!tA�3�^s5B�U�A	��ȵ��Ze;DdѤ�z1Eω��(2-Qv�c�Э����R�[E�����$Er"��&m�o*��Y�g�:� nն�[����G(��Gm��'TKѕ�Cn��r�+�����meX�*�̩��^K0i�S8h�*&3�ެ��fػݭ��巭!�:���[F��6*�U/O��4����i�)�ouQۃ+�e� aj��;�Պ�cth&��
î��]�N�٣4p��3!*��(LN�5��,3���m��{��ۨ�E������(/�Ma�y$�z��J�ٓoL��(��l�Kf��r(��ЛM����#�5��fyA0�eU��ޣ[c"���G-����--O,�3��c��Ӕ&�b����3+-<�	-��Pe��Պ�V�I%��ғF���7���:����&���K��y:�gYW���m#B�;��3lt�=��c�0�X�A�)����Jn����{b)�V�"��g2��N'Y���gM��efL	h��^*Ɋ�Y�U�Xm^�Un*��2�ɻ2<1Lc$T�]!M��o���.�wQ���Uk�D���U'Ҥ#*��7q�����Oh���)���/tT+Hݬ�[�W�J	�eGa,p�B��İ�~�vED�ԢI%i4�ē[�V�-H�iq��$b�E.��g)�r��WD�J�N��V��S�I��I4���UD:�[�@��'��T�9k� ��uZ1�=�q�Q{�$�+WK�v�)I.\��l[J��f��ňմ����w��ںUydQ�X�WI��%��]k�@m�k��GWbX�\�j�o���K�5v����,k���\�n-KA�W<�^&��&ե��R)J�g#�r�"4A����_Y;mH�W4�RE_dmƚ�qs]i�X�ӥx�]�X����A�K�eۼ�ا'��qkJ�j�KS��@�"ԉ�诒j�*�fK�D�t���س1G��Yj�X,�	u��/��<��b�����Q[H
�q(�j��]�b�ս��U���Ҥ�-��P3V�z���D��
�-!���X���Ҁ�N��y�5����v���m������MV���E'��TN��:��ꚩ���sF�⸒�f4� �]��5�9e��v�'g9UK!�W�BdܪF�R���2
喜N��Դɥ��Wh�F5�ڀ�"��@�&�rqPMVwy�5��.�q$�T�JZ�Wh�����uN�Zie$������ԒFւ�t�I�K��ēL��_)�p�J��^<��S�b���TbȺ�4�kT
�ִ�/+*b<��k9`;���JS�$�&CK���8��Xմ�rOU��n�Ij�I-��qX*��b �^��~�TbpJ�\3]�i{V�x������MN���ؒ���b���x��Uʹ0iq�b�X��Zk#���V�.H��\Q'�^v�ܷ��&�G�I��I%�&�k)Au皩.�4�]+�5ں���J'$RآLh�i5*�-e(
i!B�X�Ҝ��J$�4�%�(�+F*�ϝ@�/w����o��\Yf'ʮ�=��:���<W�bQ�ǷX�Q�����,�ie�=q�J׈@��)lSJ��E9r���5t�FCZ�[jbiZI-J����借$�%IjT�4iz+��IbT�t�ҥm0g���J*i%I4�X�4�e�r�X-e�)��I8�)�s`z��t�
�lf7ɥ����P��[��ry�꘩`��E�I	�3�X�$�]+��0bK�5ID��)6�DI��[GUj֪%�Ŵ�%��WI�ژ�+��]��[R�k�-P�����X�EqD��Z�V��5@^���ky%�\���[�Z�F��r4��R�f�J��Wkt�2�ĚQ8�+�y�j�\�S�kTK���#��,V����n'K5[Nե赩�iX>�iTZb|��iRȩ*��\]jZ<�\�b��$�S̻�m�.҉j�F�,H_8�j��O�b�]R��*�Ŗ���b<���g*�V+j�=�);F�`�l�ɲ]��ػ��tV�b�����kEt���=1���x�#��6���5J\����M��Z�#�z�.>��H;z��F����(�%NF.�AQ[��b�+��@�NE����bIR:��TW�5��.���m�JZmbV�E�'EiE�j[��q@P&)$�\�׮;I-����$��mf$����]�k�"{��,�%���f��%9u��)e���3$��q.J�y]�m}圭-��c��-SU�wT��RŻy��Uv��n%�ōNJ,�F����z�S��}����r�VA�8�.ӥ���ыi[��8,եIls�뛊�^#��Q%��ǔ<��PI��E�J?Yf��wW���f>�>3�=6�f37����$?�Ï�(��r;}>�!_Qp��}_�?��]��t�L�R�:Ű>�5 ���Y�'�,����=��Ň:�<s�݊���ݷ,}���!���yr�f4��_y[%�Gy�6�=}EO�2�)ꪼ��fޮ��*�5l����tF��6K�i�CIُUCaYЍ;zMB����@ǧu��A���܈�r��I�&��ê�P�4�|��KS�^�l-�V`���:�W��V�]^im�6N4���ɼ\���3�ԁ��D�B�H�ڂHVQ�jP凒�ُ&%R����]�/0@�H�K�����k�[-lm���!>�ח����c,MJ�7�O�����ͤcRe3F��&bW�4�/�Fg)����+]�PeUH������b�&�gle2�Ͱe).��^s٧�L�h���4� ��IX�G�Ш/nd����(m+�6�2���ur�S3��g��DVv���U�^
[�]L��ħ�Ζ�l<�so ]+Tb��5�kr��R�om�M�L�f���ŝ�9>Z�Bu�S<��Vڰ�����FW$�va�P��ڜ݋�W8؏y�=[�es�Y�������<��[�,�NǴ��u��2k���6��9u�K}��+U�ʾ��L��ˍ�Z��njCJ_d ^��	k�p1n�p$�ݽF�[��F�Ѡ������_[ڈ����U��{u�׵m��|�d�C�&6$_FD����qז7��mz��Z�]�yKƳ��v�F3;J�&6u����Br�����L⣽��(���Cw�Y]W�Rz/h�l��6�d���1e`�B��k��^���=�Q�y�zuܪ��3;����ť����M��Z0r��8��ܷ�klWK:%��ustT=˞ݟ.&�D�"��6�H�Z 1�{
���Ѩ�N���ׅ;�fI\s�ԏu�}�X�r�������'���MlXj�J]bw��.(ͅS���Be�ZC�+�54u�2tp-yG���L]��6��2n�(�[J`ə��k\��ZK^1�D����h�TKS���z�3{ɷF���{<|1S�\9F�ɔ�bv�p�,	
G���г)�*I��#�WG��v��FEm�7W&ve�3�5Z�汄"R+��k�ȨYw,jN�h�Ø���U��������ŚJ�r�o{��Nc��n�
w7K1S��f�
�Sd�Q�c����Ѕ���.��Y)�m^��)��8�*[!ȼ�� �L#�.��:=q%ܞ*����s���â�����r=8)3{���H��L��*�ou��w�̹�������A��}M�-U���;�G}�l���J0rW��E�.wSmԱ31��TUsǷ��������$���wZ]�L��g���lJt��/p1��y�%3E\��y��S%��]i֧����߷&��xI��&J�2�d�B�5�u�ٹ�[��9}aХǋ<�k�"ѽ�xYκd�$8�r�~�E���;Ay+9M�&l���4&+=W&2�S�)[�c�և�cj��S��
���X��A�4�ElqU�#54��4���-�|L���lZ�p���B4�s��Khӡ��������o��AY[� |�i�Y&el뀮��e�4	#�V�o=4��ΕC����C����A�z�⹑��쫢j� ���R��ݳ�:��Nh��}��3r��(��u@����,���*+ؿ�����&���o#+z-��K��,�.�EuFn��19���3�2�\�N�6�Y��s����	��ű���!���hK����N���n͍��8�L��`�����B5�v���5w2���HJ'�șd�m��3���h#�7L��{t�m�Җp�^�p�˭�GR�wS���A�s�+�'6p$is�W�ַ4+5�>��32���D�n��Hܼaū���ϲN�\�z�W^@��0n�êL��&w	�4���C���0�;&�r���қKk]kf1�*�c;BՓz�F*�4�:j�L�t`��=Lf�x�&"V6���.��3�`2��u����	@���1�ܦ��ۿ+���l��)օV��F��lQ�e*��e�@��\:��b,��X�O8v.���ڨJ�]k0���u��l����n�gFݷ����,���U^�!ȡIcy���7��C]N�����4:���e�t�n�=�(+�uwŽELj�n��*��6��V�0�vӭ>��(��^��e�a3�W(�Ԗ/�����X���z���{��Z�Y�l=+�"�v��;�hbPH����:���t��oF ��R7r���M1��g��%e��a�+���§��.�Y�Ѯr����iNL�nڵ��UY����T$_�r�ӏ���FBW)"c5� nv�V���!�F�T�Ύ���y{�ʱm��
O��;fF�>�z@���Vp7����z�\�x�Dҩ��u����]�_`�,ݣ���E�X��z�H�4�@�jf�E����{Jڱ��>��#/h�G_<{k5U^A�:�5X����hj}�H'��F�˽���1x�k��J�Z�����D!G�� ����׏�V��S�8Ò�lx$�c�4�2ͬ��β.����X��/��X���o�J�l=��o�#�s�{�om&���������ŵ�����*����.[t�e��8?$;3F�ţ,*�inі��IN�έ��}�5�K�7i�hZ;��\��\�/P�i�w��.��G��7�e	�]٪��l$�����x�ѻ+_3���W'qU�j�����5S֮lΑ��#]����	���W|#�y�YJ뷔To�K"����1��O���|����(�u��뙽ͨ/H��I"�WGs�#'ϛ%L0%[�	�Cr�k�K$��L�N�y�t\����cWԮ�2Y��݋2�!��΄▗b�N��Sa���4��T��ە�ȝպ�q�X��r3|�[Z�nNE-��Q�eq�[�����\��Y��s����f%��|!k��j�Pwn��1,��J����)a7,^��Fd���p�4����\9s�%|�o�Xs����n�Bz��3\����GnF����ܒvr�s��]�2���R���lJ5�S��'vfP�;*Q�b�+��3%��}������N�,���h[*t�ɛӪ�<�5���C@X$��	�rq#&�9�lM�.�co����Ff֚�0@�8���7�>O2���/!�%Q��vU�41�;��@�ke�E�+��K�ʳ(�v���lj�U���i��<�]�_7����]�,�_q���!uE��ї����N����4vl.�LPM�T�p��'HZ�(K̔��S䠰^_uc:!}npX;3��
�7�E�J�ɭvi�r%n��VR[�ݐʃ]�l�jK��&_XJ�D��TtUF�˭���w]�d�X�B3&�������g���hJcM\��o&ʊ^�"��k*�Q��T�tɺ��֫� v�JwZ�]�97֊�8)Ÿ�s2PH�n����zWJȎe�q�s��}4B����6�ȶG�\��S�[vZ�F�����;��fITs�*���ӵ�Sn[��m�2�WL��rn�T��xŚ\:�\uoaڧ�q�^�Mi����H'm�.V��Wޮ�u�����]c������R�`̎�.�iI�5ow��xK��@���`���WM���G��K�~�U:�E]g��͡��k�\�D~	\���{��u)�G8�9I�9���ԟUt�u����3�p����]@�7j�e�w����A�v��^�V��K�w����Q��e!�^t��P�'c˃R�+Xa��^NE��ǹ�C��rK�%ڰy�CGg4��\���u����WC�1�����eMvYY�7b%�s��<P�J��|6�����|���V)]4D�r�N,�FvQ=���	O[�o�c�!��3�[�Y�׳yQ=w����Ys/J�c���d9�(GI��dk ���G���μQ�]\|,"��LNwyU�3
�M`��#���I�ے<����}�I��-l�om4~�*[/+��iP[�ӹ�!B�=Aŋx$ĥJ8C�:Q����xQ��Y9R\�$˫TM�ꜻ�W�s�G!pIF[Ȯ���u��Y�'�kݍ�ő���3"���=¯*����yϪv�5>R:ceKwR�A�Mu�J.�<����NH��m��w�ֺÜ�(��6��Y��̰/�̝���*��;�Mb�
�cY���[2a�-u]BѸ�c�XZ6Լ��by�U�E�uN�ӎ�hCFݮ}ͪg���»��	!�6��ٸ�&����h�(͡ةԠ��q2�v� -���(�[T�1�a�l�`��!8��z��*'v�Z��WӕK*Ʒk:>m��v��h7C����m1��u��ʕ���I��7��y����\�k�g"��50t|H�Q����o\,�Y�Gh�|5mڗ�kl0�>�Q�IYvm�Z+V˖�Z��;��)K%v�2�)0�'�uJ���U��2�;��{]�]ܮn���ں�N�}�2�_P���qni��=�3�.�'(['�[ðq�>(;��2�ުe�7���R�dZ8R��4kw��_�sM,N=yK/�1�9Jm���Mu�7d;�Է�������1�<����ڽ�2��5�<X�%g{��\�xlM�J�Gsr2`�ﬕt��N���:�LA��5���zq�\���-�<�4�̜��o�#�X���^�WwK͹,��)P�s���Όmen��F;�:t�E&^�ض�S{	���վ�D����E�wx����+)�-I{���gf�\�3�+�0ς2o!E�-+��α��]�K0�;�U�q�]�r��y[(kMkgT��h�Ե��jn���$�H�&f�4�t�[�u��4��U��&�1ME� $ɛj�v`x͋H���}{x1\b#n<	G��j)N��a�������eX綒���ƻ��Mf�]b��8�ʉ���k�fq�΀K��M���[t�l$�Z7P텊�zr�q;�jI'k�1�)���h={��WikF<͐�n����YC3Z��V��q�i����h��'(�r�Ӂ�N��V��t�=�<t��dWG��#ܑZ7��D]Z�f�hd�����_N�nU����$��B�L�(<�%�f���tK�8	Se�'n����$]�1fI����pP���g[���aqϻ�T�\�8_=�"����%�Ճ�UQ}U�( �7��(�ߜ�{{	4Q�k���R��Q� τ�da�֏`#�n;����;	�n_+�yt"n�����2�D99L�����j �޻�ȩ��G��J�P��x]!�����PA3<�+s ��$F�&M�wT�@|��\�H&�"�U��BT=����C�'g�u��+WHnj��@~N��q������; � \;�p j�\C�@�|�Q�P=�|��n���y�	���r�p�5��������B{O�.�Y�N�y;���nT�z��DCػ��2{*�D�v��5�i����ȡ�nh�b��3�m=�D~3z������cS+��Cq������1�=|���x��?]J��yfᨪrs��'`��(@�T#���+�R�*"0

*~�����j��)�|�Պ[�w�~�������O����!���?+�-�ߙ8*��[�[��"���9q�=��I{�ws��%�;��(�uszf.�iXZXu�D����b�>+�����9����]u��t��Q��@i>��A�1�k�`��&�ujO�� k+�)h��/�9y�҅�܌IZKd��6��v�h��u��N�}�x:��s4{�5p,7�u,�sK�g{U�hի��\�����TGv��B�tG)t��3mN[-"w��]L��խ+��e��-򜓦�kN>�p{Ui�8Ni�OH��U�y�2���j�1@o�;\DIe9���N6��+X���7�4��۲k*��5F�e_op�X��h��նv���Y���u�d�ב;�|��Z�K��:�;dP��k�sA/Sõ���5�<���ꇎX�B�����$����L�+��%'9a1���MC��Ly���lJ�}p.�k���thM�!�7.�u#E؃-Nǝ�c�rigvV����-�<���c=G�Xǂ�B��U���b����+W<�#F3s��jf���Ҕ%�#�e��W�Q��,�(k����������f{��;v����m�i�8�8����8�8��q�q��q�N8�8��qێ8�<q�v�8�q�8㍸㎜q�v�8��q�q�q��i�q�|pq�q�q��8�8ӎ8�8���i�q�q��8㎜q�q�q��׏����__Zq�q��Zg����>Lf�&�u�¯���d�j���j��UNvD�]x������f"����=x8��^�����\�FCԕأ�h�EJV�ͺ����`��ު=8�.���nǷY��a?�lL��G4Ԯ7pQ
�16�T��@7,�C��]�-&�>��z�h��<<}|Ь��i�a�uve��{��!,��tP�6���gM/�*��R�{/m*²X�+����2���ʮ����j�rv͚̪�B�n�����W�;�J��0ي[�n;����- �9WGNV F�Emq��4�n1z�ivWo[5�ġ��x�#��s��	[�恇�.���f���u)�8:���]��>�
��1��k��o�	ɞ��wZ����hQ��԰`o�m�`i�S�|��q�;�LW���X�u�J�/w���\o'+	q�RSV��/!Z� rۙۧ�^���[�-K�stL%�ok�����-��.uY.!ˬ�C�6�  V$t
�X�1xȸ+���YU�S$�H%�gP�ʧ��{��C�]�p��8}�.u��
5���\��o;m��"�PC%0uz^���k	�*W3��_\m۷׏}}x�8�q�8�8�8�돭8�8�>��q�q��i�q�m�t�8�6�:q�|qƜq�q��q�N8�;q�q�8�q�m�i�q�q��8㎜q�q��q��8�>1�q�n8�<pq�}}}m������8�9��{<}��w��UmF��sR�4��' Ȭ�,G���� �N��_oc���Wt�S��ϒo@��Ȩ)c_
9/3i�a�c*��8��������,�fr%Z<��� <5c�҆��5iD�3���At>���d�9(l�KHdZЛ�K�g������w�Bq�d
�+��<�|�
� �x=U��K���8�!
F���t5���v�VY%
�.���7����yu3q���k���)��j#���d��ܶ6yxx��{�*T�x0�fV*
����5�=�n�+���:��0N��»����ۥ��h��[TL�Ͷ�<�#�诩��ç3��TwBf+��>ޙ����\t;�*K���D��d1kZ�k��|�_�ZP�"���l�V�:f��!����<�w9	"�o�>���}?kPeĆ;�v U��"7y�Ư+�.c�G����՞���`��_�9q��U�6� ���V�<�g��û�'���G������n��w�P�s�����f��T#��r@x� W���fI�W>�����$ȃ>�sr����9ݺ�� ��g�.1�S\�'��L�mCW�$�V�Uj�����.�{�.UyB���Ń�$1��ܵı�1TC�v��6e]JnYZh�Be�nv�l>���$�����wu�/nGpӣ��������W�������q�x�8��qӎ8�6�q�q�}pq�N8�8ێ8�8�>��q�q��i�q�q�q�q�q�x�8��q�8�;q�t�8㍸8�8��qǃ��8��q�x��8��qǎ;q�q�������>����q�88�9��粪\+	����%.���]�@ň��Fa. 2u}M��Oӕ��Y�;����$�@m�#���/m)La���v��2<=����#�4�&m�9�f�Y�<,���ɋ*�ֆ:b�$b�#��VL:.�"F_����Cn]ru+�K�i�皔��,u��,tާZ���	E#t:�m����c3{Re�V����`����p��xS�W(�7����ŉ�{��8��ۜ����)kZ(�M�XbJ�:�'|��4崙q�7�����]�\W�}8�H���]B��F]{�]��:��0���!����Mk(J9|�u��{�	���2������&��� ��U���G�b�X��v%v���JV�$�U]��s�
t,zl};/�h<�J��x�zJ����u��AN�s���p|8u��l�D>�6�ϳ�orI��-���BT�/S4d+-U��]yr��Y��*�%=gC���r�.���``ѣ�r�.P�Ў��K0��zGuk��c/�<��	��5��+�최X�B��SǺ��������CE��e,+]��^S����U�i%��B�X�ۺ�iX��Z��@A�K�ɗ
���y���ӟ"�fwm.�K5L��RW�Rv�[�Ǐ�;v����q�q��q�N8�;q�q�8ӎ8�8��q�q�}q�8�8��}pq�q�q��q�pq��q�}q�8�8㏎8ӎ8�8ێ8��q�n8�<pq�qǎ8��q�x�8���q�m�t�8�Z}}x�>����q��8�<f�z��=�^��f������u{u�_9,��N��(M��M��Q�2��5I�eIR][8/�Mrc��!aCu���t�R��8�L+A�9(on�Rګe1��S�.�ҬJ*��ii��zue�[VG��k9BÔ`�kN�d=wO)��K�w��X��\(��R_EێK`���q�gv#][����q��x��|̖x���qx�o�њ����B��:T���S�͗�ʷ8k�#W�:���k�W9_-Ե��|;6�b۬+�elx�Y�
ѧ#>�%��l<Fˋ(�4���y���!�6ڬ�3�d��W@��֝TM̧y�V5��;�,����+[�A7�q�x�^�샸o3y�k.��*�9�sV2vqV�]�̀�Nĩ�z����pe�V��{���\�j��"T0n���]�'7&3/x����e�J��;�N{0p ���1k;5�*6N�Y}!%�����L�UYmڣ�B�y{�
�mX�ځJ�X�޸�A�;@�3��g��i/X#�'�%��syƏe�TP���dzJ�{��3�����*R�c�����.�L�2Qǘ�կ:�{|֨ƚt����Ǐ����8�8㏎8ӎ8�8ێ8��q�n8�<q�q�q�qƜq�q��c�8�8�\q�q��i�q�|pq�q�qӎ8㍸�>��q�q�qӃ�8�8ێ8�pq�q�q�8�q�q��i�qӏ����G���px�8���=jMʺB�,�ْ̳M��]��ʼx ɲ��a�'w�+ZW����]�eV$�`ˬ�j�J��W���&>�\0�Wk�*��3R�!�8>��Kȯ�U�����D�ϖd�{�S-�!�ώd=Wܘ|.�Qw�]��Wkolm䥔��lH��+i���V�i�p�I�wN�%7��x����KY��;�dN��y�^��������7U��g��Dǯ�>�X�nc��8�����s��6���Y��{9p�n$~9}*�gc2�l�ǧ)S�Y�����q�d�g}�1����H%��Y�0���w�fؙݗ�=�K��iitD�0.m�9�Zoe��%�� yٻ�	�t@R����j����:N*O�_A�Ƞ��L�uxve	��@���u���A���1�LU����V���r���<��
M��$U[\<��T���m���L�iL=E��+_lx�Td�L�/z4/.�}0X��<���s5v���� 4qQ1�$p���A��9���t��[ڋq9���a��VrG�R}��}���ui��`�[7��KVb��t��w`uJ�w�^���+�����<|q�Ǐq���8�8���8�8��8�8��q�n8㎜q�q�q���8��qӎ8�6�q�8�:q�q��q�8�8㏮8�8�8��8�8��4�|q�q��hq�8�8㏮8ӎ8ӎ8�8��q�v����������8㏎8����w���qf�Rk3r�F���}�\�WZe�g�ϨN3m�Np�f�k�4�.��������u��&!N�X���m�����껠��4��ʙH���e�3^�j�glz�DT�ݠ]X���x� ^]]�V�嗻}:瑩7M9�s�*� \���ox�WO0�eD4Ko<�<͜o��[�p�SkEZ�Ĵ�����eҝ�q;��Bs�4ق�wsj�;�:����q�n����������xm�:��y�/2Q����3�!Srk�����s�Xt�jĸl�Aڦ+k���s���q��A]ēB��e��Օк}�t�k�
�V֖n��g�E������ȍ����BSC)B\.����y�x��,w��e-� Z8��K�%��W�V�P�&����<&�w�ľ��3N��������/o,I�o[8=�W��jo����:�\���hwpsm�@
�Y}��t\��I9�g16�db�_N�] �wT�6f<u^ҚE�U��+�m��9F��< 1(����Og��lݱ�d�&&qo11X�"�Rj�[]]
�*Q!��f��ϔ9�^-��a�'-�O7(_e
�c�|�,S��ckh�*��9��խav�e�m��b�7���T�5=��!��~n�wc�-���D�.E���ٳc"�']T�K��=��RKy����E�M�ě��N���Wc�=\;jwA's��9���AJ�wj�:�$5�w^���w1�KY����7�,�mݙ[�}X���	wl�4�f�Ws���W���Z+�@�gurSeTQq���V(;��HZ׍�P�1.�Y�Ƚ{��I���.���a�m,d�ڱ���$/#�-�+�2����|/z�.Zm�1����C�7fu5�*��WT�sx�q*;}O]��]�g	��M�u��4���:o�o]`��h��Ó^��X�����z����C�ĺf� ZY���RfL�Sr�Y
ޠ��1/iWu���2��,���J�EO��²Hƍ�/P|ؚ��Ln�{���-=��W4!�s��Q�8�l5�m��$`A�I����U��!�l��E6͎o!i��or�:�f�}(�����sC��i��3�v�ҥ�J��TUue�+o�Jơ�KqVe�*��0���}]Р��h#y`�Y!M�Љ����QŰ��;��۫�1$��q�Yum�N����t��q�t:aC����eL��f��2���(Ȑ_^t��v�םm;�h$�e��{\��i�Wʬ����������:��rn]L^a3�;@}	���e�ī(t�_.�YZ싷�����8�2ޔ3(����"d��\�Ϊ�+�r�tCt�%�]uj������FM�P����@�۲Ec�z�geC�i�9k�MOs_+���BN�V�\�d�<�!���ΑoX��LZn�zG֖��b�ךնB��ZLke	4�FmcT���N
�
���2m�*�{�ŗ�pݮ��K a��x6�1��M��n�����f̫�-���������5U�dH	X���c�u��A*���g�V�u�ZO����ٙ�,�n8
dS��Ƭ���9j�:[[�vgv�c76��ZL9�:�Ok\���lG��-�P�q8>�l��Wz.����J�J����8$w��2Y��Ҫ�C2�d���Hbxx��WE���R$��9x�'u�걓�XGN�Iۺ6M��(��s
�O�;L����v�v�n��S�IJ���!f�3��N��˷������;]�5͗��5��������^`�a��V,�ų����E��(p|�f�c�jQ�湏z+�r�� x�n�)�a�։ĬF�7u�K<2��kr��9/�*n�ӌ���WV;f�3Z�p4˟D��!9�"م਌=��tZ�-y*s2��K�n8Ve�>��s��r.��A��6��˚�z�<&�qLۗ.��vAy���Aw�ӵ�5�Ϸ,¬ܛ���9�y��o��1]���|����+T,^��|k��(_�L���æm�='�ݓeL��f��-��w
+��f��L���4o)H[�ה{]�䬷�jI�U0B��x2�*����T����I�瘜Πc�%sC;ռ��nqW��[�E�b^�����b6�v�L�f�����P�؇!�y�q��7Y��/p�ݬoRr���&�c�f��.����C�����_��������_����_� ����߲~_��ey���nh�Q�noIB�$�!H�l7)P���f�j?�@�'�&���\>i��l��0���D",0TM8�`�9�S`2R�@S.(� ��6�I��ÈȔh��"�4����H�Bl�ҒO4�ND��a& L!jK*��)��jB"���D E&�I
���FY�ƄI�4�:q�owW3�x#��<["CA&�B6�$��� ]Dě#��0��J*8�`Bh�$*��a	��B(`Q��a��PH�H'Q�H�'�!�Ą��K�8���FK��D~P���S(@�-#.! ~F4$LO4}#,��L���e0�eI��l��j)��X.8��3��U)q���A�a>+Є���n"Q�M�L2ɂ$Da0�"BԄ6ީJkȶ�R"'�)*�i�K'�b)��m|��>��a�,�@�(���CH��?^��3*��cp,��uVx��.��p%AƝ�����[S6t=�&hS`{yY��+�/��oH�I7a��N�z"�.feu��Ui4�� k&pS�l��x3L����~Y��Q�؜�Ԯ2�+i���ﰽj��NTX��%wY��_&e��q��l�E|Tw�*od+V[f�%����l;�>��ͮSq�Z�qΣ�ѻ;-����	�dXUq�t��Xh;E���YA
��y7'n
�uuǁ�Q�sT����ޚ��1�E��x�Dkn,Μl2�\�[��!��f��ܜ:��Z����l}1��k�
jOl��A�'�����%�ӌ_y�1#P��������:+p�bU�:sEm*�֦�̢_'b�VЈ��`��f�a���(��}��M������b��st�b��/�(KS���53V�XD�3M���K��˺ȂGr�˵���YΪ����e
��g�4*�v�ę§L��_7�XF�V��-����7�e���&��	S�b��XJ����4�r��	��H�1����ۉ����Ѝ��$�� �L5BaN�@:�Q&�
"S�����H��Q��bl�*A
	2�h�⑄�1�A C0ȣe@���x�y�Jf&e qGA�Jdm��	���d�D�&�N@�A*8I&�^��P>�D�	6",(��.��|Ci1x�P��#�~'��%(��H��m�h�Il�4����a�m�!��d��0)?4��&H�jz��h��1 �M��2"2��l�#�7!%H�."�q8�##^,��)x�$��M���q� �	ce��b2�e��2A��ap��L���	�����FSMP�LHJ0T��Pڂ�$��`��E!�.8�0�e�A!��$Kb0�H�U�p�M'1!�9Q4c�[�TC ��l�T �& b2&"F!�	 �aF�P)n(� ۴���b4�)�m�Ln(�1�Q�L'<��̸�:D�-������
p�̀�Ā�bAe$b
&��F�p$��0���"�J����e��ba��A�M���$�q$1�$QR�LC���m��*�D"d���a4cf(c�#��@ȈE��FR	!~@��p�"Cq��,�J$p(�%	aQ�ѕ(8�d��1	-���d���S�$B�E�DW�����1J�(��!
��&�I�a Y1(L�ِ"�EJ�D���8:�*��	2��#r"�>,���%zF�*�L�,@�b�	4c�@�a�Fʁ.Jp8��Ȑ�#d/0T�e�d�f'�$L%��2���Q&���D#i��HF��d#�'K��Ɗ��[�$�L"�Mǜ���Є�"ͷ�r�!�d")%�NLS��t���ݻv���1��L�B��2��%�L�%|�D�����3Kv�mHU���,��ʁۜ�HJYhD#�DA�5�i�Dj!$�j�[��o�v�۷o_��1��}��E���gv�J�,�!)��26���,�%�-�������#%������ItIUe��O4���<�i4n����ċ"�75I!,�s���,�������1"K��Ib[��ƞ>=z�۷n�_��1ә�d�&Y'm$F���)�i��������%�!kͿ]��}i._Igv-�k�ԋm�'n����M�w<KݲE6�E�I���V�oRh�RὥI!㡧���v�۷oG���>���vkD�$b܄5`� A�m0��gX�s֘���v��mR2\�[�h��w$�������;m��n�<z>�z�4�^�;C��toD����Lɶɐ��S=9�''i�I�$�O^��M�!�=�N�M�t:v���nݻ|z>������~Ź[CD�v�]\��C;N�d��b$i��9�ܒD�O	9�����2a&B���m%�&���B��_ݣ�]�N��x��h�M�������,$���I��w�ݲF�_:G
�HSm	��d��B$�\�o5٢v��&�
D�rI>ѷ�{m���E��K�nFY2F�n4P�� &�'��R���DH� (� ��c��D
ܞI3n����0�Ie�'�M2��c��WGWn�d46�t's���ջ���Q{�V_#1��Bw3շ���A8�Z�BO�,���DPE��F�%��m�e�a�Y'��8��8�
4L��H"p0A��~��\%�Lf<AR(c�BIjH�	��<Ze���D8�@�B��Y^f8������	�!mB$1��IA	D�����A���'M9�4�?d��)*I'�@ D�6AL&���P=�#���;gv��ݓ�䆣2n'ʹ�d��/��h�!+����~<���׫�GF�F������z�b�����g�W�����_�og�l�*�7�`ʋ��=���/ƥKȭ��������e/��:�U���:��{��7�z�j��^H�R{͑~�ץ������w��Ħ�\�o�"M�[�]-�it��&��CUTZ�SK�\+Q'�܁Ava���
����0�f��to����*�[|������0o]�ш�w�ィ=��)e'W�5%�YAN^�1]��sadk#�:�T�;�=��}��l�gVa���6����!y�<VJZث2�	R�{؅�{�Nb;�{�~>*��z�M��*��fy�����6��5����ڝxm�B��ؑ2�T��^�G�^y,��ag{/׏�v��+�F7�Uvj����\sy�t����@�]�mNq��y�V���L�;����T5j��ϠJg�}���8�=:�KU{�κ{g�yֻK�Kl`�*J�
w8f>g1�N�Ʈ�	����*��U��q� r�_�xv|�H�oԀ��[N���<��ub� ��5�{�Rc�q{eQ �m�� >3~�1����d@O�ꤶ,2���f����Њ�~{|�׬j���Z�-x׿O8���J�C.m٪����J+��
�8���+�Ln�΂��%=�F���|l��Z(�|w����Д��?Op��:�춝�H�����ո�N�t1�+���s��.��}+>���p9��gŪ���w�ٞ^�	(3��!-/ �-�� ���k|�M�4�ׯ5D��zTR��j�5e^N�o��������ӱy4��>���96����K�/��=~��W�]�u?S��L��N�z绶x�|�ϵ�F�垺\�94��� �������.o�XFn��[{;
Ҽ�kӀq�oo�fV�Ѡ��z�:�|Wp���p�=��
������F�u�,q����a�y���If�Ձ�(b������t�of��u1�e�7��ͬ��$�,hxx�z���� TŦ+��Nd��v�bX�<#�,��Zu�Y��O��mg���`l+��%�$�t,PJ����u�}�yd�|��5V��<f��kQ^���E���9z�k�-���xW.���j�H%Y=X�S踤�ya'V�I��;[�	e���e�eR^P�,�� �#7,6jS�r��o=\#��IJ>�[�w�FP��$Y�e�K��,�3�����xbT�sEvʫ�i|m�R�Yn�b�sӶ�~5/�HΌ�Z�"6W���{�>T�в��+��������L�{ꎎ�K�ٜ���b�p��E��C� ����3f3��7�mE���{�	�b�IM:�e�e�Rh�T�Am������a����}��=��R�,-Z�r�lg<؋䛧Z���I�'�eUp��z�z����2Z����ܺ>�+�I$<��lgp�{��Z>���f��!���ݭ��aYA�L�PӤY�� ���}�H�ݽ��j�������{u���ʾ�s+ph�̰����iAլNVBQ����T(8 �Q�r�f�<�-'�z��9�,�ކy�k�#r��y�Z����P�9��n�u�K���U}n�4;ֵ^��:��
WG=�}��@h^K��W��~��>G�OǷ{��E�g��٪ߨmPrJXZ�ҽ�!��J��f�+�5���|<lZ���j�^������e�61�ہo�1�Y��B'v̍7�NOf���%��TϷ8`�!�Wez^�3�ݮyN����iˮ��oA^��'~�>���hu�5;9>$�f�ʍ�Mb��Eb��/�|���� T8[B��UI)[�lx�"����_'�J9��=<���G\��u3O��� S��&�o��p����@���/?C�2�;��wl��n>�b�{k��;�xb�b��G�}=���u-�ueUÙ���)��X̭��:�.��AZ��Ð����u^��7$\L�GP�JP�OQ5�O�ٽ5��z�W�Y�Q>4�t���2d�5�A�5��L��T�E�q�#,�e��QG��{��%�2e��lAQ��f�pQ`�߈��H�$��8P%*E��_öP+Ǝ�!�X���[^Z��V��@8�]F�X����@����}�}ܴ|(݉F?�����0m���$��<���x1��-�7�47�J��x!��{�&�Z|,|>|[��`a�_ْ�iپK�9�p-��'��*F*��/�p���(�}C$VI9�|�n�E���v{x|�~�3٢�כ�b{�'�g�i��fu���r���.�>n�	O{4/�
�����fʥL�M?���<��B'����}ܡ�o�����!T�R�,�]g1�"�A��_z}3j�S{m�IG��t�ɛ����z�Q~�#0(Hc{7��}?%�S���>Xꣷ�~U�u`@kUԇ�������<�I�^�v�S&�K��j�ź�==���p�Kˣ�K�;*�7���gJȤ��[���&и8�������qP�V�찘x=�H]��t�깡V�e1B"���Fe{��fvY����r���>�����)m�G���K=ٜ(�a,E��p3�a��"�=������Y �.��;����y��i�g7Y�q꿄���>/R�h'K5��h>�6�$p�yԛ5G������8ǆܧ���y��UZ5���"��i�l�i�x	Z����0!��\)nIU��|L���n%pb�m�ƣ�sm�T;���!Y�M��"�c�˥�m4��:��=���?��T �4��S�o��)�UfF����($��Ue�����ɼO)�����H����o�cȁ&ҏ8��Y�Ƌ,�UP���S5�F��z�`�2�M��fA^�a�fo@Qn��V'*�(�]VQ9�H��P�,���zJv߲�q�<G(����������_w���}.ڮ�s}*�E*/Ss��zs���E��}+�+�������H����Y�1Mӿ���Ӂ��nߏ87�z�8��߱+͠��K&U�p�-2�`����w�Qp:������+H�f��v�G��3_k��{��{��x+{��rCR� \�u*��-�:�՛{�ѝ���%�����oU��� �G�@��>V�}�������;�-��]��!�%����!�P��,IX���`J5M�B��� ˢ���h����\�~��)���I�=.���x��7���;�;�b�g���Q��&��4z��iWD �)�+oR[�dG�eJ��-�fc�{}z#��sz{�=���h�t�aѠBB�+���i{�0�!��'���.���뜭��S�;Y�ޚ<\L�폪�*�P\;}�H����1��U��6V�V�-J��ǒ[d�x�o�>m�M�.������&�D������5k�i����/�V3�߱��q�q�N�,'[!%�*�Y�jNy�n��W�d�+>�2{5$
L��?2��1	9d�)�fB�/};�׫v�gэ�Z\��ڥ�>��m��v������G��N ���2��o*g
t۽IE�ziCUХ�{������M�}��=�6�o���o/i4�X�e4fc�O^n�"Q�̤���[qCoJ�B3����=#r��N��Iǽ�#�����;DG���=[C��y�OC�{۔�Ǐ�*���0_���!����Ɇ�.�o=>���P����;A��)��G�b���o����
��	Mi�Sj6��̞���`"�?І��`�_*y�]�z�~��K��޵г�yG|H9���8s>����뵲�6��*�W��*Ԇ@�п������]	�S�h�u>��K+<����3c���]m�Z[G 2J�J��ܑ[���m��{�)G�c��N|X�N��i,Wf��[�.��lSr�)�EbJ��Z�Z���.K�"�p5�S_)/��~{{�o׳����">5Q�_�Ytb�8�0�Ge���غ=��c��kU��^�}Eyy����t�Od�^H�uJQ}^����=ӗ��h�Z�b��d�vِ�'/rnS���Gj'7�v������0E���~=�>kwʺ7�<o��μ��%E�M/<�Z��P�3N}���s%8�3Lޫ˨;�P흢�z�|ZK�z�	�nҝL�ܾ�`���� x�򒚋R6�0Xl�䀟<Yf_`�|`��L�S��S1yx��HI���6�DF�2ߡ%��-�
A%��ŉfoB[�AUmJ�q�Q���
�u�r�P�d{����3���L��R<�i/e"˺;��)R��uc��Z	�+j��RL��+��[QV�@�յQ�5�D5o�����ޖ*O.��>���^�ײ<���0���ԵO��>���p0�_f^^�,fI���_۳��}��z��\�G0+��U@�-�)��NԤ�Pװ����l�ܦQ�Q���"�(�"q�S$$��˽D���iWy��Db�� A&z���S��ϵ�Z����噔=�,�6�@���^)����S�Rb�si�Ts�G�H���p���-�����nF��vW�?e����|`?o�:s��1�_^�x3���r��0��P�A-S0�͖�����j�K�����7Ф\#5Ja��b1�TI*�{�L�����
��g�������z�Z��V��k�ݺ� ��p�V�ʚ��^P�J?	k:G��]{�]t�[��냖у-�9�M�i�����Dl˚�b���̥��2j��;F��u�ݏ6�f�+��	!�F:�S|U|��{�>~#j�2^�������o��
5V}#�M|]��G�_9z�./��Vח�n��r���W���8�L�
�0ob��E[ѯw���[��7W{]z+����$�cJweJ��ڦ�������r������N!���JY ��xlSz�b�K' �n���1B���+9(�bN�n��kp3}�"3D�3�ZV��kT6]������g��e�]~���z��
�DP��v����*$Y�ܪ]�T7����:��/3y�qM�.�ui��d�]�U�όsk'�=ُ>��һ��5���-���#GG��G���To(����Y��	�o�3�G���ݼ���Ҳ8e8��,�A7>�ﴻw�k7���+�|��= ڢ	�3��^y�I�/�����瘁6�M;�f�n�c�Z������;���&)�����YQ�k�yC�^^Q��ȠM�
��ʓTo"���9� /2*�^i����j��Iٚ���[c��"�;�l(.��`|�Zɛ��4�͙6V��+�UqU)u����ۏU&��ƴj��l���b���u��n(9;%��9î�qP��ȇ	NSn�.��	6�^��R����knw`�#ȻS���B
����ِ*{$�ʕ���w�A+gwÛ"�,Q�J�#�`ήZj�n1��uۋ\����d��:���y��a�F.|��� ����f��Γ ����n&���cD�Ǳg(y^c9"y�3�M�fGqcQiJ;�"����单7�#�
P�Y!Ҳ�����;c��n�8;]Q�}���[��H�s��LC����f��w]�Q�ʐY��z9�X��M�VV����Ee�N�u�9Upq�1A�,<����M��c�Ӯ��>�r��+K!a��+�Aqe�)�{vD��뚺!�c�����`蝄���m0^��3���ljw�7nP�%Mwr�8�Wov�On:9�\��x�Tt����kR�W0SOM���s�nÂ.�"�H�e��$�C02D oqc���S^[D���(������n�G�tA��(Y��YZ�v%��V:��4[b*��΄�B�U=~D�	�T�H�٨��C��G�>a�1�Ľ@�Z3D���$�K��Z
���|4rXh23]�r�����Gc�en��Y����v�]�3���/MU'[�0�s�:p�2r�C�M#�2�[��]�,p�N���Z1gJ�}������0�hއ��;���(�hA΁Z�f�s0�u�����vC���f�T������x�}J��p�6�]5�ݮ?�{�l��.��6�2oT��+:�x'/���;s��S9G/��uU�l��]��w���,t��ٮ��W�\ݞr(!ͽ�b�NY3!�:��������F��ܵDU�;�>��ӕn�ۋ!��1��ID�w]Jo+���DwDY[6�ܝh�B�n�(�NL�����{h")����B��7��7jR਻*�J�7�c�\s>�&��}YDʺV
��Vbo� �o-R�½OK���� �ە����ۭ�%1�-�vɢ��e	`"Nx)�ڸn�y���jve��ݜ��G�YP����hΆl�5m4�e�)vU'юv�Erll5\��J��%]2��{n#�A!2XDB_��Q��tI̪M�,�~��<q�۷nݽ}c�Xƞ�����(^i>�t	��]��A�ѢL�0ɓ��Hj���n�=|v�۷oG�ׯXƜ��i�N��6��,!QNMP�,��132�R�%�5T�kTx����ǯ]�v�����]W���>�zԚ,,�����ؐ�~�}��$*��0J�8��t��o]�v�����׭4���k�fH�Qa2e&L�&XBe� Q �6��C�o^�v�۷o��׬zӞ�֗���^Y�;�!;6�F��DQb���W�뷏^�v�۷��׬c�I!{�܄����$�!�)D��C��-e�D䚤/�C�}��ݬ�ؒf�5���Ž�M������B-�6D$$$��k�D	I",D�E�L�2�OV݂"B �,D��d�Nc�DF�dv���"%)K^���YJ"�	����I(��G.�cNy�l�l6�a�A̼�zZ}ŷx��1D�ъՂ'^���b�Jx����zx���=1�>�ګ��C��ߕ�������>��p�@q��7����l`���5��$�]`6��g\�V���|��O���0Grp7��j=w#״�췂/a�4v�
l>�}`Җ�\[$Oqћ���ݻ�$ oK;&�sim��]X��T�dT�T�q@ǵ� #u��T��/9�����;��Hm>�N���MP7pQ�o�@T��Di��᜜{3\���VfMP�}7Y�{��D8(�� $U"�a�� Y$��<}����������p14�]�z������Z��oU�s�&�� �WnOe_K�M���0xsQ�!�ۀ�˧����p��»]���R��%:�S���:}J\�� :/
�ou��b�%�����#�E��6ۈ��R��\�U7�+�ݼ6�؁�x��~t´x���k��)�@_��}x% ��@�5���>x|&j�H	���DrA�>�*𾮀(� �ʞ��au�C�Xg����<�_�Ἔz���&�����L�s{��-�������ģ�MA[3���;�z�D?m�~�kb<7��x����°�1>`my^������u� F����y�`}�8 ]��������aJ�v�ܵ1wʕ[���b��Ȁm�(�x;E�vN��=�v�-��s����^kI�%�c���%%6��@����FJ�%u�v;���Kcgdif������s87��WS���}�C�2�C���﹞��˩�S�����߂"�>>��I�F$5���`0�D��\�t 7v��m�	�&o�4���:\�{� {ܭ\�K�*D�Y��z>��k"e����b%R�̖��t.ϒ�n ���L�=H�ގq>3;������y��Ǧ��{��C��_�'uD�R^W�����G�����9����[��:ڵ������ �]��(�4r<ʙ�����@E/7��v�,�f���t��@&�3Rf @e�����;b�{����4�2 �d}$���؀4�b.xVjƻ��@{1����7�� � y�7�`��4 > }�p���{O�����<��,u��<NΪ���Y�: i���y�������!���0,���Q��A��x�S�O��ո|ycIV3�� �~�tI!����5����q�����@8���U}dY��1�$���k˩]/�	8,`0��9vH1�V��ouK<PΜ>b�m��g���� 
����]Jsv/-(�3sI����5�:�?��3���{�
�^y�M;3�<�k�v3��YgdN���T�V״�*H�5�+s�3���')����C'5���{�W0��+^�}u"mVL>�=�.�ⳉ���Бz���U�.�Y�23N�x�Wu��;�1��.��Ĥ����UJ�߃1�1�5^�ٹ����p�R�6�$�Ye�*���n��	�A'H�2BX-��%4�m 
L �e&�0#	!�j��)�[��h��йd�������+�y�Z�m����y�$4@|m��V܀5s�5x�Rq5m��������˶��>�|;R� 纋�g�, _0�`/I ���
�I��O���ܭu#���N�}cHa�<��|$6u�[>�y�3�����@iƀ����a�ݠA|� L0J*�ut�u�N�F ~����N#t��uY+����%�+���(�Q|p��@���z�j3���3�3��� ��|>�7�{[�������[	���-z�S�
�C>��U����=w�4@���Q�*���>������@��w�R��S]�4�-H}�?u� ��O8�;}a����|6?a؟8�_���^Q���V�	�l����4�5i�@0��3�2�}�;��	 _	Ӷ�&���A��T��{����������EV�*g����)b"���-*��u�� �`�"}>�/�����b�(���n>6w�ϕ�>��CǄ	叾�1}����}���sܧ�m`$�J����BT d��Q�O��e��f�� mmL�clqy?}v����v>8�3�\���~׎U�GO=��$�$�.r��s�Ne��O4�KP���\}�|����[��U�$]٣�He^�;��Va��b�F���r�9힃9�GK��g<��۽�޹���?0c0c0eg3��u�g{��x�&�|򴗔<@7�N Mu	TQ����3�O}�c�
2ݴR�ܕ0���'���l57�y^N5A���a��$gG��yH�^�	�vo7��0ni*b��kG�tI�脗\2>>#��\�־^��g�{*���Ⱥp��q�}{}v�^�n@r)�v��W}��%�F�}����� +]�|8ȡ�|������o�h�M=={XJ��{�>��n��N~G��SM|1S�������3���Rn#��|�������C�W�'��&7uf�bM�@�j������=՗S�=u 3��{��0h��0@���u����[{���:����VU�?�,�aI�6���l%���[�v�D2Sӧ�x�'�wT�������sP	�Լ7�?�������hb��R͞¡mp���[���as�Qsz
���D�;Evzp���Ql�|�(�I�,*��M3�V�}�S���`m�6;������:�#�.p4������=	�i����s��u[x^�/~>
�qf��a�����|�ϛ�;���&��O�]���@],��������C[�tX虖���O�[pT�sQ�Bo�j��N���fS�V$6�z��͒�^��]�7�<����v[��qzW�1Y��7���j<'R�=��qӪgKshՋ�!��uo��	ڭ-�q����`����������^�{�]o� ,�? -O9)�d(#�ɏ0���w��_�W���:}>A�/�s�&T��"k�����v;�Ռ��6ۄ�a���G�[}cP$zƂ�߼א4�~ @����?� ��u��F�Ƶ�ͷu�b����i8}<��G��J,�Şk�	LA��]��s�d�q��TK��f��r��j�9��=���&O��~0�sX��n)�7�����@	��I�Ưx�g�GæjZ�C��_�?s�g�@sl��)z�����~O:���_�6�@w垘�����w]#�NT󭨋��s��8��[���f�%�{��Žgd�Y�079_�2�'�~�"Wx��a�!/Cg�>0��
���2Ϫ�>ηe�^�~VY�8~I���� ���?�8��ד�o�AY��gޯ?�|mj�J#�+dWI
���ynIx.'����n�9�������G�{岟�Z!���(򋚷h��ӓ�y٧{����tIz�Gdb�"5/E�:0�t��e�&^}R(���$PU[>F�n7�WMG�=g����M�5+�d�r���S3��;ĵ�\$�:��4͆/�w��#�0f�ޛ�����^��/�SśbZe-�-[�U����7��J/*=D��<IED�}}�(U )wS�3/1�!	t�Mʼ�{7Nj��aƪR��4�Ĺ�ҏ��O�=v9`���c�̳	���41�!\�l��ƷG3N�Ϛ�G}-��D�HR�%O�E�Uytas���>���*�;3��C��xS���O�O����xj>I�8�څ�\�wdR�]#/�>�ư�y�oM��l�:��K@�HD�6����d~�(�?1/-�̼=��o7�'����!J��Ai�ɵW���aǗ]�݊�#u�旹�xJl6�%�#=&H|<zȕiK��A��kR�L��w�[�=Ga��ۉ�5�K�Bv}����&��r����@�g},�V����c=�t;	8����EZ�V�l��Yy7�g�E�k�5�>�Òf�UE{M8����)]�sP�#(����>�)q�'�W���ړXز�z1?��������-\X\<���n��\Z����%��>�݅���+mĘ������̌6C� �bc��r"�_�3�o�MH�����
	91L���3@z@@�P�����I��9��T�V�p��+��E�)�̆pq�3�z����M���������rG�W�&(-������k��п$F��f�����	�e�.⮾�XO`�ׂCy�a����.6f9�#�R�T��f�2���g>}]��A'����i�E>Բ�S-�ު������g�D�,)��%�
@RF�뫿��]F�m��Q�>aAD$Sm�Am�p$�:m���3�t�����L�Ɖ:�͐I�k��]��<��Y��ڤ��&4��/�P�Έ�:���`߼_��x�|�vwY\)n��Oc�. c"N��t]*�y�t}C����_X�8j`5���4ƞ��y��Z�Uy��q�"��f{W�O}��g������MIA����õ��;�¢�wẃ.���xz���=�b�~y<)�?!�ʈK�GN��`��t" �W��&��ه>�Zݹ�"���-�`�������������2ů,k�A~u{�����hZ՛�6ۼ[f7a���V�ws�����z4�Ê%�J+��+uѡZK��5b86�����k�kn�HJ�ݨ�4mo��}0�{���B�A��ˍ������O#�b�p�v�d�}Z�5��l��{��H�Sn�5�K@f��Cq��?���v9�Yﶳrm>�<ѡ_$�� *:���q����5_�?����}9�@l��3�N�~������L�4x��j\"'mNڽ�@�gy�q� kv�z���u0���dNN��A���[H�jb�G� �����]{���\�X���^T������f��TM�K��m�Wr㚋��T1���P~�t�=M����G����-�M�̠�>Xӏ.�{�����iI3c\D����KT���+y���t��������=�*X� /�^3�9;���6Ԁ�Ǫ�S�x�o�����\��l>�*@��a9MA��k��M�i�'���t����;ˁ��\􇛝>�����I��绹�Y��e���[7z���ƒ�NQe8��Lcq��]�d��I(�5�\P��U}�t����L�=�m�N%"7�h;��#�[]�u@�ǽi�<�`��e���X��Q�΃�*o;��{T���Q�B��]'q�M�ơ5��k���}ߧ�V��[g�K�4,��]�������8�p�޿96��F���͊ �i�vƼ�i[5�M�A�y�obm��I.C�{�)�[���Y���Jv}���'Arx��|Q.�C<<gH�x��ugΪ4�D������p�Gz�i,���k��5,�g�İ�����Ys��A� �0g���}k�d��'r�K�ͷ&_��	$�}�^SC���ӳ���m�.��MH�׉�W�c4��6�n�Sf�����{ӬK&��r(�.��/���i5-�"n���F�;�_ʿSv�aK�Gy����q_3�qQ�/�D�C�K�c��ko�r��#7�׾Fػ4��4����6k�� �H���Z�^��H	/#so�����Sm�u+�k!/��iE}l>ze�o%�i�Vͧ���.�<��$pva�)ɼh��n� � �0�T���=�{v���B�Y��oǬR�;�5���g�ݑdG�����6�� �\[uG���M��!{���$ɓ��4�'���)�DxP�"9Li[a����^�QfݳɄSNos7A��/k�Pb��sp�@�6�x�mc31m��+�������V�si�m j��l7Sb�n�������`OM8����������z6�P��~b��&GwYѯ�6���n�Yn)�Ö�E$j�ػ�M��yT��0V?���\�7�R6_јP��q�}��u���#-�[V�dp��y�� �9��o^t=��e���u��@�
P������қ��4��6��7�Yї�׫�>=7�5��[�ޚ�#)o�K#/;�A����'Y��`��f��n�fy���؞w}��lޯ�S��C[k����E�c{���gPP��h�D�f�������ݮCvW{%��1:������|�T���Q�Nʿz #1§"�$��z����}��}RnIR	�%�w�>����S��E��{+��~?g�}0r �����J�@P揰'��no:}e���/��ƚ�{�g�
�@�[C"	n�]�y�� �!/.͈,s��mbNޅ���A-�^$�\� $���޷��f�6�և<�UdS�mq��#&����Ψ�q�v�_�C�`�``0`$�\ ���Vov�[p�����M"�5�e����ω�
3��u�R������5L�kT�\2w�L�9±	,&$a��_=��9�aA�j�B�~��}W0��h=��
�)��Φ]����������_	{�GN�(c>6��7*K?*���0{������I�F���d���5�㽂����a�V�h�"����b�TAK���f}��{\�*���Z�5e?!�r�����d[�5V㬀�^��eGCN��qB�i���8@�0��{�4�v+9g6k{ MO?(�g�����.�B��^���R��r��;���?]�f�@{q��=�qn����[��oz=���%�ꁦ&:p�����Ո�a�M�|-��R��끝#�	J��#"���^��dy�/�e�qҌn7�a��R~ڶ~��w-���{�L&ov�ǟ]����������D�AO������~��յp�dA�Vm��BPxy��Ŀ����Lz��kT706���;l  V[��=�{өF�(!+�� �Q���V~~��?��+6\�E9��@m�.�W07�+�r��f>�tl�X��I���*�Vl���8�uWʉ�8����u�����{�D��-�^���N��I�<���[v�~2�u�U����=��:7���j����I�{&��R"}Bu�f�o.��2-�U���#�/��P�v�,��׍����gR�SОZ6���n�Õ��x�q�DS�b�ͼ�7mݣ7+6���[���1i��Z�-6̺l�7}W� �_T�e�v��n��ܽ-����S�rV��){�h)M�rW�`kG���"֤�r�'��OB��y�E�.?�Rzf�ؗq[c��JV23�^�,��w�w�bV�4զ�!l�g�a��K�Pb�j�{�P]�U�k]]��[��MÜǒf���S��ɵ��[�OS�о��d�i��\t���h�v{��`\�k��l1)��ӳ��[m�W�	[��[8 �1��OD��Ď��j��F�\�֧<�T`��8f9A��Z����ӽ.���wJ��_)����ybQ�/2�)�j쿦թ(�7��YT�2'
��G�=X��t��W"Kf�<���Q4� �����Wn�&aE�b%�A�Z�6�6���:kq�Y~s/u.M�U�z�j
B�-O�GĠ'tT�(cyH�)�Շj��P�ZiӃ#׎A��02i��l�}߾�Zf�v�/<z$7�v�`M}A�u�����9��ї5��V�������QC�p�B���нap�t�|��v�H�Gz>t�%]>�7����e=�i��ay�����Rsg���+xI���m���e�r�dJ������r�O*)�g�l!QKo�&1�(W�ˇ�og���6ή���!p���c��MC.{��C%��cW4"�K�8��F�j)G]w�KŸ�{�j{�G�ٱ8e��c��e��S�4�z�D7���	���oL��+*���3ˑ�g��L�s�̮R�L�,l�}s!�U���x�cw��m:���
���ϣ���v�r�20C+n|l�l+��aoaͨ�(��6��3��'&�:)̢��+wnPޮ��}�v��\wD�����$�f'�b��+��qm&Гr���{��2w�I���NeJr�u�l��%�I����i��5��-�Ie5v�zV�[di��f�FQP�z�->̮�lڎ�}?�����b�>��>5�j�]8��� ??��SI�孷B��f�M��vm!w6�����A�ɮ��RM����sN�n��۹񣜔Ơ���99
����m��H����2y�D��$�D��D57o�c�۷�\v�۷oGׯX��2�U!"HH��H"�K�=$�a*1�K���a2�$![K�~����_/��z�۷nޏ�=cL�{
 �%�x���J�dQ�ϕ??7�ﻻ��*T�z�Q�XӦ6�m�nߒ�ߗ�U��R4�>&�\�m�ږ��
d�ʊ�ܹ�
�%B3��P�z�n��^���oGz�}��$�U��0��I�]�1T��)'�h�<�*z��:c��ǯ��x����Zc��>�$�>N����引�=�B��"|��D��� HI^��Lx�ǯ��x���~_�U���̒���B��t��E� ���a(�������$˜�y��h���k��H���T�&���6��e%D��D�"�$�T�Q�MD m�F���!�$��	���eH��Q�R��䈄�قB
 �"$���L�E��04�D�Q6�R�Q"f&ډa�a��"A	ۛY��܁�RWv�|�ӱnq�Ǣ`(�`Z�f�Ĭ��t�K:^+:<gB�\���3,0\Ah��l�K��a0�)���j4r� ��pb�%($LE�
a@P��򐀛-��H#2C���H��-�����$��A0Kg���(&�-��%�)F��^1����!	I1�%�H0��q����M!-IH�s�6[*�d~Gqhj�(`��H�:�hb��������!��R"�B�N
;����e=A
)�̍))���H�R	
K�@̍�K�^n6e���D��� �����|���� �Q�@��#�U��R| _��S8	`�ʟj�����8�8{�l�,����-��`\��y>��ށ󅉞L3�xQ����T͘�avO���Uo��5��mCڈ!W}�ޤ�>WKEeK����-}�<���{$��2�g��s����,��J<�"������l$���H��j������\��ݴ@dz94�]�I)�x��m{�gC��=�ZÁ�m W�^Lo��֦��	�,c=�߆�S �����=�,�ѣ+T؝�j���.v1����5����1a�ž��t�x���n'�V���f�TOu�_[�~��u�`�
+ԽD}�o�!���U�}�A�$�美fhI��N��R�~Ǩ�U23,[�<�;9uHX����7v��+�P�\
 V޾)�@�S������b��|ܺ�52�21;3�ûvf�a��-|:�7Jղ�w�z��O��Ƚ�8��	�6�f���mL�ѷ�U��hz��krQ��끝�v�o�3e9r�V��=Y/FP �g�(��j�0_o<����U�B]wKY�\�f!-̐sz�*�Y��E$��L�>����^l�1�L�_`�w�!�ݽe��\�Au�3�W:��_�+Q�)1�N�G���A�tT�w:��+��W�����/�s��o��	�1�qV� b! `Pˮ�y������J�k�Eu��<�A�ᑱkQ�[;醃_��y�h O^���J`�%������\���4�J`Y����n�����D��iG��-�#�_����&���ߖt�]��	`8�놭n#}<h��y9�%��(E_?[~�$cC��4�ni����ۯX7OxN��	��v���4Wd���N�>;��x���聅�1��%gfЋ��<4�p�};��n/;�-���IcW) gC��z�����I�������^&�;�&s���c�4��.cC(#�����{�C��o�E��w�]��O�/m|�hmT<	���v��$����׾��{��~��ejz*C�}qe���>|q����IM��ڋ�'bSL,��K� nn'�i���r���zP��@�v�	@�a����l5�5�����;Օ5��n>���Y<i�����c��5�kG�4����P�鮊wVI5��M T�ūc:i�vv����F�QɄ���X��!g-w�N/G�������כ�
��Z�&��NL�Ӈٗ��5�b��,Զ�6��+�I�fCMn�������kN�M��Op� i�R ��D#� �� y�z�n�����4��3�����Y�6V�μt�l]�]��+{���Q�enP�jͣ��v�ޔ���g��a��0Gq���b��(�` �Ξ���������J�^"�~��G*���|:-�(�N׍S7r$`l���Ե���X������ÑN��ֹ��FL=:��T����]nEt%�J�1�S]u5���t=�0!��MY�T4Y���ik��F�~0�#�c��Oi���p}vi�+����%�QK2����=vހ_Z%}ɐ�ڀ$�Y���Y�u���Y���@�߳Z��h�b��"|ه	�t�m���g*�������G�ﶶ�>��&L���G^Լ<�q��(�Mwׁ��i��5me��oQ�1�ȏcFâ��M����kJ�4y[���S��4��V��[X���W	"�Q�����A�Ā�\M����q������6\�u�θ��f��1u�ӷ�9+a���p�՛D��U�[8�h,Y����a��D�iMg)�	��,gq�S���s����� ғ�J:��¯�υ���9��:~:�\Q$�P ��.�Qt������k��V�o{��x>ǘ���9��mÅ�Y�8��c��e�:�6ϟ��[-��R��g*��i�̻�YN'�w!8�
�2����$�K �5v����K�X>c� WPQ�x��sy�ᩎ�f�u��ɸ&Z�Y"�a����[;&I!�A��6�fU��y`�� * �D �U �O�A���G�� L�ղ�8���?�23���3��&A'���D�b��~f�}��Uѳ�� q���J�)j��K����NKP�k+��J�������s�
��-��t�.:�A�#�zl��7l�L��@Tg�y�D���l�6G=��mg�ra&m�˂��B�}&����uՈ�՛�z��p�v+g��۞p��j6X�r���A�(�+v�G���4	04���i��$�=����ܨ��陋T\���Á`�z�[�<W����4�n�wcL)��ۖ؇s _ڇ������$�sj@�N��'3�Ə58�
���{�.x��t�Jh��mv\j���!�:�ǯ\�>}dI�eU�,BM,�Z�N왫�_�˞I�fZ"�j�hǑ�ܞ8Qއ�������fҊ�]�G��>W_���y�y��mi��%X���u^�j�Eyl�~�*hKC��w�1�5P�^/�ʱ��zZ�0��]6����MQ�����Nn+m��?~��_s~G�yѺO�'ָ�K�!=��B���Y6����4睝�J���L�s����=�m��>���$L[���tXG9D�v&w��	�*1ؕ��}�K=�ʻ��:���{C,c�:eu���]5���X�5�F�<3�՝�6���O�1�D������#PE=�k�z�jBhܚ�id���|�~Է�m^Ċ0��0�j0�rb,�h��E�e�b2RN?��O��FB ��/�%|#��;��-m+YoL�=��=���|%���|2�[�Pd�&��s��HȷA�n��#LO+��6�1���~�� �Ӎz(~�q�������̼�/ݎy��a���÷�r�>�=��mO�c��ig�F��/������z�tkҥ���Wz�Gw���1;�sَ���8;�6Ǖ��x���.�3�Ys�w	��!z��ǝ���⡪[K�(9Ѥ\��y��j�x���a �%'kosؚh�Zn��u��D�S���d�ѦL�!Ʋy��h�����/<7 I��	wN?Lu�''/f� =��@jw6xm���a&��$���d6tp�L��pN�}A�W�������ԕ�
��cQ'wb����z��}�=M~aj�\��D�����	��,���vO)�HG�� o�����<sly���8�͊Y�����(�$_ivأ��B����y����rx��ET1�q0���Ϭ6���Z������w��v�SPц:���)]���ng���,n����wuO�a�ɑ����t�H=[FecX1��z�k�X�2��Mg'ĂI ��0�DD!)=�D �P�N�ۖ8�x�<���b�)��N�OvV��i�S!��/���D�6y|}�CH1�C1J��Q0_������P�h��n�}U���m��W�"�q���?��&>c	E3x@�Y��^ޱ��[�
��~H|~D�,��9��z.�?:"=��f�=���֓Q�3��7�g�z�-]P�D�θwh��K�E���ӭ�S���v�p���"��F�q=z�r"ZUS�;ɣ�.z�O'�o	�vd�l�i>���\�Î�'��3J�����
���p;��I�c�G���iSP�ӷS[1�k��Y��r��|��%���m7^��R8azqq��,i˞u��5���WC()�ks��TD�u7�ԙ��r��U^w��H�ߋ%&�܊_�̷��+��0�P!��j�~o7Oli����&�h.��z�ln��|&����'�#N��V�+��}M^5Et���aަ��&B����;�����z4QL���-gy�����er�׮���
[�j�sm9����6��"��eb�n���{�X6�y��=�����_�����~T"��N>5��9
ܧ�k3ىV`ܬ���2Z^9��>i��Y�~���NӚ��K�����ƥ�%XGI�����
���5i.�5dH5��<3�dyn ���;t�/72����E�����	��sb�}v{�ݜ?����{�A��
|�CC4U��
!����}��˟>{S�'�}�y�Lx%#jz(��>����}atͩ���(@l5�5���'�#�*}\,тɨ���Cdb<1���@������Kr���/Y*�0�.�v���&ڡ��ƙ�/�M�tY���@��T��XE}�����虪u�̓�D3;Q�����b��E�7P��z�\?�7�ɖ�$�:��(������8��y�[)�z�7����؈LGĂ�!��g��ђ	*���v�;"x5��1BS���؇1w/�W�!��@C-ߢ�� O�$���.����G3x뮅�w�P�^��s�Y�_��ь}�TC�J`W�_�_?;Ů±�#�]�-�ʇ{�Ձ�$��!�cH��3��2��T���d�:6�~��a���?;��4�U(��#���A8��T�6|�.��C��v>�r{Z �v��i4Z����]�1���$�h�����te���9U~�G4�>s�n��"{���ӏ./G1U�w�Ø����zB����wl�7�i�%�ơ�ȉ�|9�!&OMt[��mӳ�\gj��hn�9�	�Gk�wk����q/1�v�����%ئI��!AYsy�o�c�.�צW]��O�
R+�Q��f��mґ�lz�>��<r��vrU��cGb)<�Y�ާ����K޹�Ԯe{3�
}UH1NA���((0`����w��M�׭?5�=�� �D_G��� dӱ���q����}��21̈́�����)��)fp�ya�xF�o�F�i������V׋d~��s|�6I����=S��=#O(���-y�
ާp�P��.�,�I$
~ߧ�������@��_�Tt�~>g|�􍜅a����.ژ��L�<�J&��]JY���`
�%�R��u�Ӱ���x^* �� �k��lp��SH��qI�7��.�t'�j���������q'�_�HOesz����0;�@��o0a�-�5G���`��8�E=H x<�q�t��_k@�G��i��3���Q�i� ������%�Xb桵Zq��`$��:�;S��؜8��h⾁�q�2,�M���l��m��V#Z�*�h��D	�A�	�.��>_i���	s�&�˹��bMA�s=<���/o��+��x�5�mBIq�6��0
�g0#z<ڎ����&��oC=�먮�\�$��o��%��Ӽ���mI$^�y<���Rv�4!Z�˻!�dq��΅��𢡊�6��WP�l�7�Te_:���� �ң�"�@=׏��C	����(!�
 �@$H$O�@�@xQ~V}�{��mrĜ4���88�1��o��Q�͊�� �-Íd�}Z�![�9�Π�>�"�(b���CH0DS;.�I�'���U��;���Rj�����?gu�X��q2`��DH. �`��h�<瓌�[ L� ܞ�~�	U%EZ���E �r���K��f�g?f�%���>�ҏ�'h�I���5�bޖ,q�iLևֱ7ͫڥ��{�$�/@�=/c)�����F��z)*ɒ�)�ЫOn�^n��m$ivI���zH8�=X�}(}hF?P�V*eŧq�u��2�k�{'��İ��|��T8a�}��߱���J% R�g��j0��{�AqG��?�Պ�Z�i�bv��q��t��ot	�ؓ�	TS��H4E{9����'�	 �$-���u�v�y�*Z3xxS���ai�e�Tr�𽊀��	���x[��0�Է�)�eko��>����'b��@�`;h�At��kF7v��H.����ȳ�'h�{��D��V%�<5�vG�@Q��.�=�}�s��>n;�<��7�{*Չ"���w������n��eP�SD��?{�@�d})��=�&����	�}#�G�y�l��u���йl�!��7�Bf2���T�Kz����=��-���a���g���>LxE�au� Q-V�A����*h˳y��L�%8�cWֻ~}S�w5Ѻ�n��O�b\��W=��;����*���+@�(}�;�n�2b34���Nѵ�A4a��H�:lb|��A
�LE��Gsz�º��zۅg3��Ͷ	��h�,r�<�"�r�R�ڲd2��:'�q�C�UQ�� C S�(`A�� $��`�l`
��Ϟ������y������Q�xs!�H"Kx�8��-}����ϩ��m��1y���ЄS���B�{���G��������9ǉ9���K����Z�?���Lul��a��-�{��I.@�]}�|��X�g�n���w���0@c�߆�V���\n~�������E��cYQ�ʃ{������	�0G�K8��g�2yv���ׯ��N�Ё9)�Z��#2�&����GsW���I��y��܄�k�E���u����{3��3�nO���=��y�����ߵ��č��?
��Q�}�	p�&`k��_=�8u�E���wӟ�x��B#
�DRE/�Oe������Og\mW���p9ew��$��Q�O�}�t(;�W���T<�)� �Ā�M�S��Tp�%/|�C��H�L*�')ȟ{�l b�h�>�8g�o��l�񓼜���y/�s�F���cq�#���i?��U"_���u"G+�v���ǇX3x0������Z&�1��`�	��rwA`Z��8��Ky�G�}����lĠ{�����v �_��{��xt=VJ��h۩&�;_�fn��N�u�
&�MoFu<E���m��`��sڸ��;����y�ø]6b+wj���ζL�`�y3Ɩ��T.�QS�O�M��syv��ɾ���jo���[�H���o[k3C���R���p#X{B�I��9��>�Z0�N�^-�ض���b�xٔ��V�,4��$�ɉ孾�n�{[���#[1N]u�֎�FԽ�u�E��Sր����1T�C��v���q����yتn�H�dq�un�ڳ���l�Qn��Ǣ����q����R�+v��I��}��e[
#�LE}��l��<�{6��v+6���cl�h�9��ar�Eb�l���U�C��o���o�f��͈�4%��f�[c,v��^�L
��UV���	KLdü�vv��Գ������f��Z�f;�J���	��fs�β�]���Ѣ�;���.>	u�散�6md�'�oC+�@m��K���.�\�)n̺4��on,ê��u�U\�u��6�i7ch��u� �MǈY�O��aV]aKs,����y9����o��\�D�w�V�q�l�B w{=WY��y������<�L�������*��T<�9<Ne���{r��/U�PG�HR^Z�d�m����b@��E�� �'�@}�IH��!�D�͚f�BZ(z��yV����?R���nׂ��;i�t��U�x���$�훺�[��ֳ���>W0�Vp7��eΫ5a�Ds�h���yt�uG�;��͓.����L�m��b�n�1��Z�v�-F��놠�oj\���U�/Y��Nu�D%7۫�un��촔�aI�/j�YW9,�Cg��'���r�-
ӓ��-A`��Y��}���}U{(z��{iڝK�<��zj����s�n^c���m��LgUq��)/�MT[v�kq_lhK1���S:� zL����F��9i�{�u�(�iis�О>;�	�HnV�̚�DoW�yM���F�v�m
6;r��>퇶��-�������`5��K��;��>�;AӻF\�c�V�	��.��Ȍ����9̙�"L�n�0�ך�l-"�3��<�x�]�r��\]�M�9�
�r�f�Z"���xp�����ݜ��Z��=Y)����(!�;��z.�A�Z��6��=�����&�ǰp%�5�V�h����5�R�lM�V\��^`��\�x�ZT��1$�ۓmb=-�j��UӅ�����"�{�F��N�,NѴT�����/�*y����V�1�o__x����=i������j����c5.h�p�T�$��4��i��z��<z=q�L{�����eT��J ��fNH�
�!&�QRq�:c��^�6��ǏGz�{���]����{E��ȰD���L��3#2{�Xӧm=z���o<pqǭ1��u���%���rfK��D�$z�Ȥ�"<\����ׯ�^>=x��Ǐ�8��8�ڌ.W�L�P%AdD�6��jZ�e�%D���j������~�|m�Ǐ����;��Y$�UTUp�)!a���H���D�|q(O�!Q��4D��3Չ:/m���f�aJ��K�(���ȫ'&���r�UHZ@"�se�	H�X������R�4�
8P?Q�"���A9JfA��!;�I�sv�	 ����sV�m9��7gRY��N7.�y�"����q��V'Ɣm���.�YD�"����	C�
 �0 �D� ���畇�0@�HJ����5_6�cY��G�@��x�֍����(N����aUÜ���$6���o7z��<�O�G��]T��kW3xEW*i��!	��4yU�TZ�ϳ��݈w����ʌ�/�֒c�^�v��	k�eBo�����/c��ɱ��M_]Kо^�v�5�*uG���E�$ǲ��`���v��=�A���ng�;ӽ/���u�Z� ��p�M(�9=t}լ^S�i#cv���D{X�7��k\O���׋���D
��r��-���������W;�_���Ac��5xG����^2ueES(
�b��_�fӇ}�z������yC���u���8C�QQ]I�/�>�.3Z϶��ѯ0H
��]KFVٓB��'P�季�����sV��#�s,c����dǘpXa���s��^�c����~�R����ѬQ&r#���H�~A5g���Co�Lhx�׌'܋u2�=,�έ��p\��]�2��o]2&�@�)�����}_�>V��]lI��~�N:��]A�qǶ�j��ϙҦ�ƞ�L�:���w0���*g7��l��˹�9��TA(��3���2���=��<�ӯi��{msZ`��PqWU�o/�*%�\�(�A@ܧ���z����}F�r���U���_b���`�CN��
�b���C+Y�{�k��0h�i����h�
����J����_��3~���:=�$�vv����'�Gz���@f��3y�V���x�\�"\uܳ�c33v�5M��F�i�;m�6��� ���X��Ib��A�����J�,��t�f���������Sek�J�"��م���V��WU�gw�o�z�	?�H-!�]-R>I��4η���4K"8���$�y�W�^#V��M�q����0㴦�8-%�_���I�8��#;�����_�WY�3�[� �<����3Ee�S��'�.	z�R��<`x[39��§��ѧ���O-=w]Y-k/[o@un&�n+��ƕ�d@M��l*KQZH1>o3'� t�7)�ot�rv9�ut3i���kY�������ϨcX[O����wE\w8���C��G=kA/�Ď�Y��Y_>*���C��Mw=.���}��7,�/3z��g�7m_Iy�P��j m<�m������}������ڟ7sn�+�A���"��o�{���%�/�^����ΌМ�U������:�:��N-֩Җ��M��껽�>��i���7X+�1q
�����i�3��'^�6�U5�.N���Ҕ�ߖQ$n�뙕z�W��^�����r*�a��"Ȩ�1P �C�P���t0���ʚ���NHTv�q)#�g�}2oӅiE�2���`4a��̑7�^>P1"���3EF�!(�@)���%/������	�����+y�͋�ŭ?��aDY�ƶ�k`e�w�����<���LD���6�0�^���%ho��>���g�O �������O}^:��q��|"Z��.�����ג��Y��|�O�g�Gg�Ӥ��z]w���:����_����BX��iΗ	�T�m-�lX�#<����;f�<��A����� >������Q"k�z
0�� �6�^�b--�v�Mγ��=<���ٖvF�㡖@�y(�O4��~r��;�dp#H�ו!��"|�";!���΋��3Z���)0���՟PS��E����~C���%�NSq{hM�=�z�3;J���/����RO2�yd�A����Ƹ`��9�4D����y ��w�e[S��A�!�m�ဒ�Q��${��'���ȥ޸���R��^�H4�a{����n}O$��\̇1Ňj��o��6���0O���JǊ��Js�A��5ż=�+�f�J��>���H��R�'ti�<���K�C����8[�K�����
�B;w�+������>tS�C�l�|���B��c]g8�ѓ#��z��/T��ũC*:ޖ��hvG��K� �<| �`��"P�T�Ȉx�  ��3�W����>�b|9�E(`glx@�u�������r{�TxȆ����1$�-C<�뇞�׍v��� �W0!��o���i��*8�l;ɶ<���q&Ϥt��Y�T�lFv�pՀ��!�P�o� @���T)ab��$�>!�����ߐ=+���|������.�ioQ'����8�6���ߝ��Ç�'���~缊,�j7:u�q�����ٳ���O�o�7��0-�W��W��������g��6:��%�B<��R/[e�7�����f<�rDY�M�`m�7?�5�crto�W�vυe��4��g��,dbp�c&������{_��
�W'�p;��~\���.մ�v��WN-���\ a:�8	���5R�gCY��@�i/-��:��I������t3c���8]������b[X��o����гe��n/�.�����^��nmq=V�]�k3p��-I� �F��߯|y����AT����D?�l�k�F��iߗ�׆�N�U�.bU��*Р�i=���7;�䐾׹���!�2ñK��)M��hg��'ל�e��Pt�^�dH���ؓ�ܐ� ������^j�y�+sUmwH��${[qczp4���꼥 9�Z��n]���;x0�Nll@<<��I���Et0E�X0��C
�������iv��W7QsP����>�N�l/��k�6@�{���lH>}�Y=HN��Q.��"-f��� 8Q��۵��r��v».� �٥����чlL/bY�sL�cQ�c�l�~���f���ߣ	}�WR'�Gu܎�v��k`A���n� �b��tt�����"�`.���϶�퉳�D�������NT���N�6{9�j�+gl!����1���$� �ps_�qY%`���a�Nd��8��������i/ǧ�ѻ�.0ճ[w�/R��+�b��=��|�"�O~������������9����k�a#g�	��VP$���؅j�s����&q�Z��z�����Eמm�5��O��D�κ�tbte}ރ�F57n0I8�Be��~�z��ݦL5�D�����
�*��G�/����"��,?]n�:P#���s)�7��^t�{�y������=���3�da�]����~��
� Mݡύd~�X~�p�k�u�Gqw�'��H$�+�+�]�1�_0H�����ߍ��R:�;ґ���κL&�}���2�����Z%x�����z�i'	���s�~�\e�Bh/k�{�(�rz������F΂:�U�I�@�1ʳt�ʫ��v'|�rU�5a�����O��$���$A�� �������^����ֹ�z���SY�H%��]K \�A�FkH~p�S�s9��8i[���m��{ّ���Eb佖�%��x}
���<���ԉSf��@du���㶳���L��R7MG	����|D��\,��ډ��^�4����Xt�1�!�U��\�U�S(__Q�8.�A~y}�|�V7�_�	XE"��A8r���`߱�!�a��V�Ɏ�E�"��2�U�._G���A<k�^�A	�ψ��j�wk�g7M�K{��A5wT��!�*c|{{�G{WV� ��N�b���my�!(�0�IT�$M]C;^19���W�'ǴD������	�[O0�unx����[i���Mlz$�]��N��ݤJ�c��ww�d+Άn%c�k��|)�lW�<EE����[�j|�D���@�!�qV���x���^�� �5	� ѹ���°K�d������L^KkuuS{��<+Z1�wy�4�C0�q�B��^R���q9>/���g��H'
a\*��b綻�Ǎ��0��h��'re�:y��<?vˣv,��1w#��D�.`!�N.3�,�n���t��n�X��S�"���W�6�*yq�k����Wp溛��gR�=�o+�޷�3�y����a�+�R��`��J v#��˂4�\�2�F�-���?m�^��B�i�@�ڞI�H��B8�i��(�$�HRR�(���iM�>�}�=�B�����Y���7X���m3��=��`�Fǵ�˲�]5Yh�������w+�Xu�O���1~Lyg|�~��d\��f�
Rn�hc�����`�p�|�㗱\;)�4�G6�#M�HE���)��M@��TZm�%ţt�׼Ö�֝i�ڻ	��q��6U�wx��`�h>�|�[+i֏>?�]�&����S�ع��\!��e�k�2,���S���M;�q�o�W�sֵVv:r��Ѭ �i��O4��s�+v
s�=�p��G����4����948r�Ꜧ>��S]�Z�,�
��;���L��ė�;=&<�0�ӅF������L�N��gR���7rƶ{T�����i��@,�uH�mű#K��G��W/M>��,CnsGdt�h��γ �1,C9.�0H3�-��/��ǞP���O�2M\|��z"if��p� 7n��c$����f�f<~g�Uy�cCyP+�"�⁴hcX.H���S'l<�K^z����ڲ�L����e���3F���׹�nu�1jژ�T��� 6�����Μ�uI&���x��(�Eٮ��7�����u�mc�彷�:�ʹ�۷{.�0}��<4�؅���1�2��̔O��`	
`�*��  ��<G��ym_v+��s�����3\��M>?~a{}~�/�>2���N�T㶺�w"����rE:�����Wa���+����=m���� 9�yK��_O�HB%��0���������B��;��i󿗷]��k(�p�>�+�ȯ�qnӸ������f`Y5z���|/TA����b��']gF$c����I@���7,F�@��O�հՖ���>��C!`y�#)���
+��s�RQb ��=y�窟��w6��t��g}�Kl�;���q$f�=�{+بt�G4\\y��d�no���[ߌ�.C���3��B]Ѷ��x��q ����� ��ZVCߘiw������A���4~Q�!�]��%=�7t��g��n�ށX���~�I!��?�/��ϔ�����B���JX'h�֯ݰ(ķx���@1K��,��B�L3<<Y;/;P��0a��.�8�E�j͵��-��~��~���~���v�p��%v�ZU���л7�|����i�e]��)u������Lk��u���(�Rod]8F��k��;�k���"��z�"ږs� #�jK��݈�t��>������lN�y�:Gv���%�bA���oʳW�	Z�ҧ��H0D�`�0pG�_bVg}/5�翈��/��]y��������F�[��qc�:��^��-^p��Y��n99x;+�p��	5 a�>�<՝�U����٬#�"���rK�d�hm~���0���9k��� �ʸ�t��#�O�����Q�ar��E7͠�݃R�.a:�7~/���=I_:H}��_Po��Do��黯�g��TC��Vu�X뺷s���M�� ��� l�0v���S�?��mA��xJ�p|��1����(C*�M��.�����s��Fzn��]�s��Y-��"$��FR?y��R���è~���ѽ�y�[�@������j�#�>��;�|�-ڍ�A;���г�y��fRmP����bL�n7�p.%�ڟm��M��'��׽$/Mx��sR+'�lb�ߪoMwU�S�aR��|���!����Ʒn_���}>�!>W烪�e��5&l�<Χ&�Σ|�0b��;T�ib?3<rz1����*�X�p90�@2N�wկs&g��[�[ʛth�g�dV;m5g7Y�C܌ǮWVii�s��}�fL@R�S9�P'<Ȝ5�Uћ*����^NU<�! �9Yލk7Z�λ���(��e�Q:S���z��ￊ�P�`$�!A���]��y��s�����O�"���p��$�S]�~6}Ii�H�Z�||���w�u��沛�6z.��ݖB��(�a"�{�r�帅��P��� ۤwP	>&�:hu�:�B����B����`T�$�I��k��������ϵ4�0��:�Kx��:C�6(�����6/!3�!��v�[N�?���C<7����������԰mK0Mc��&ޞ�&�7i�xB��*����j��ug�@$�7e�1{����/��m(�άJ�N�)���m%����:o����aB�����v�Ǝ��1Pwm�����æ9�h�O��^�?+���MC�����_�����*y!�v��'D+G)�k�ѯM��:#O�?NH)�tȞ�Nt	ÓŸǥ���my����5yx�נ�&��\z����a	�ZF ��iML���$ӺV�cÛb�q1�� 8�SxDh�t���Aq<���J��>[�]t*|*�)�ޯ{��x&�������r��� ����4���؞um�����u�E��7͐����d��o��j��%,<^��c��7ou\ڿ<wϨRѐN����5��S[Ea،�Vn�,�c�:��b�7x������cu�-͛y�%�q:��y�Z;�'$&9�"~��������j�ߝov*���ճz���T��MY7j��{}�e�-�Z�/�8�t;�l͚g�]5_C��������l%�����w�:9�iȒl�j"P�o�����욏=����ä�N���iZ��ݝ`8볮ݬ�^��س���|�L�,�{/L�j!�iR�#ح]���VDa�dF�Ζܵm��:�$��C�U��'���w��؍�ݎÑͣX��_�3=����29�7خ��8�N��sm�-�S�7ü�7�׻�X�t�t��/&�M*U:ɱ.��xI0q�+x'(]������}�`���ۍ�H�6l5�v�ңǐS�{����ҕb�ܮ�Tm@j��BV���_Ӫ�-��*�*, ����Ptݭgab��[x�(Y#�{���+3p���_b��Y��,X��c*u�,kYxN��Z�~�s�Q����?�'N��8A���S�i]'����Z���w�(��߆BYuo�k���oa���di(T}n�a����D���3�_�ո���CD��'�M��9�QOm!�WQ�����I��C�Wj�R>�e�(�FYy�s!r�<��åR��&�J�op�)�J��3���q��7��]�P�znۀ��r������Z�Z{qR�Ǔ�ͪ"��-Ƿ�+l�U��tUl�+\]܇C��MPم��T�ao(#���7���Q3�<h-�W}t5�/�Z'.|����b�&-V��t�}�7e�9�]��tz�y:)b��刽��j������lf�9�Oj�)ꍢ.�v]S�	\3��
=7zA+�Ҥ1�4�s\9��"[ä��N>a\�<�k�C;�vv���9�ɝ�;���r90�{���E����i�7s�Uv<���క�#��uH�-s׆����|��ʗy�ޣ<�.��#6{�F�u�i��貓�*��#U��a��"�m�Ơ��;�O�������G���tֈ���3���ፌ���\:t-��t�Z��=r��д�D� �9�����#��C������h����#��
D?[�Gk�V�4�!)2�-�:)IҡT޽~���Ɵ__^>6���z�'��~$��]"*�|�Q
ze��ǹd�e"�D��c�O}|}x��Ǐ�^�i������)"HP����I4&�ETv��z؄%�c�M��ׯx���ǯZi�?B���Ӣ&�I"(��]�$"��9�%!D.�z�n�<t����m�x�z��M_�c��DHV�D��k��'�U	��$Xɐ��*$|z�N�>:z�����<pz��M=�TH����%}�32���>V�%گk�*Dc=���C׬iӷ�O�^<|m���ǯZ���>����}�t�bS4�!*O[	�h�?�羼�	�,E���~i7��b�䉫��'��$T��*�3B��� {�g�d
�Rwn@*�!D�fm�h�6Ÿ)=i5)���J��� %����AJ'���n	"JhƂ`6R6���M�_��2�%Ke��h �h�A6'��$�!8�!(��1 Po��f���j�4���fG��O��Ō��z_+�O3t��0F�:�e��R9�>l!t;���0Ka�E�
l`2Ԍ��!��h��8`S��!3HBT�H&10S�!�!��	��$3<|�.D�i"�sȘ�F�bB�!1BD��I��a$�E$#��QDYa���	26!��(�����$ ZA�.(���-(c0�Ti��h9>%��bL��i��H�����7��ܔV�[���C��:@(b�`0`�졊�"��<�]��D�d�$$p6[�k���d£���-��=p���m�Z�y4TE��j(�q@��&�d���v����J�%{�����~.� ��^�b��^� �i�%	�{͉/���/�g-��r{fLێH���	^wC��� h2+j��l��ɢ�b���c��^����MdY����^~�1�+.���c1��R���K��6�Jq�q���M{���;�a�
�)pKO�����_+Q+�W�~�ߤ�}��t���WB4����4��6�=�v�C��`$��r	�s�����w�U]�<�����3Z�f�t1�=����m�15��C�8V�.�xd[�MD�&|���un��,c��~L���LU�K�5q�'9�Ե��}�0�sӆ�\{r$��X��8p� �����h��4x���M<����m�>sx��9U!dj�x��t�έ�k0��Y�������&"=����3�K[C�!���8�i�&W���Ⱦ��f�uh��p�8sw4+qѱ`k����֚��Ӝ�ϚU�����i�����_��w"걺ܮ�,�4�dc9��U*��H`�hai�\�c+sں��*'�P{�ו6��Pu�c|�"b~��j�r��R�t�8!7rj�_Cn�LYۑ�y�;g�{,�͗��m��:O�:Gg��N@��!)A�z��k���b�@��Fr�a�Ŷ�	���lk��S��HXW���:n��NGL���k�7za���1��Jm��þ�u㚪Z���p��yՙ�=�D!2����%Ǣ���[��<Z��%?�ϥH���5�n�v�Y��v��?ٿD�����k	ߘ�߄6���Vy�@n��]y��O���o.�̴����1�g���BdeŻ9�`q�3�����Y��� i~hNC�D5}YM�>�Ƶ4I��5���y���1ړ�=����5����tU5�v3LǶ�_ͭ	0������?S�]�ٹG��F��ڐג^NL�I"�Q=~c/�د���)H���>�/.���ǋQ��K���Cb��DU�98��Q���<Ü,7�Y�a�ѭ�tK��8�[��@�#k;v&!CTή����|u�=�"s/��<��~�������k���YB�q���a,7���� �DQ�o��f��k������|֜���q��O��4�L�0���m]��vAfe�y�V�fk��d��\��j"��y�V��m�ӱ�8$��x@��{7��wa؎=T�Is:��ޔ���ޮ����6��+�V���vJ΄��UF�����{�<G�##$(h�>}�����׳���~<�{3�q��j�"�f�ݭ^����fN���N�ްv�)��P��?q�_}=���4�ƭzj'Xׄ���)�X��e���O^o���❳`ˮ���+y�y���b�%^�:��� �����;�}�׳~��eٔ�:=��s�@��zsƼ̥��±�+�@ݡdgy���]���J!��ofV�K�di��m4`h5Fe"�K���yk�ʄ�m;���1CP��o`41>ߚ|��EJ��h�!Aq3v�,�8Ɩ��o�#G�-E�l�6z0��p�Gr�[`ˮ��۷���]����\���fA�*��5q��J�0
2^��N+�i���n��7��}ޒ���f[0��<�|ps
�{X��Qw�u>�dzk�<�[�c���ƾ��F�q��FL��x�|f�uK�%H��!���;-z�f���|����l��ަ�6 �x�i<Cz�&R7.A����c�r���j0�.(��43?]�vt{4�YV�~-Q#/U۝���ZO���d��"K������놯@H{���4�4�T�c�h
8~��_>���ra�%� �ydlJ�r@ާf�iA+L�F�k�5��I�CӮٛ��gX�58Nze=�Z?��x�$ ����|�d7�y�����x�Ab����[���v6�%�����+��@��+���#�F�B��;]n<<�޳�;0��f���R���7�w=[M��'���g���v[�vL?olNN�!cc�i%�L�4Ӧv�A-�����
ׇ5�o������~,Vl��G���ja{�.���2���1U�����f�w嘍��$��Ìx���{c�)�;��Z�
�m�4�ZÀ����g{CdY���lf;z�k:	"�?�� ������F��az8W@��D�wԙ�_8��s��p���>�N��he hno|�\�ރ��}�u��8/��,���//E�w����?'���Y�}~z!#�"��M��v���B^n�#/ʃѐ�}���$�4�Yw{����h�츶�L�v>�n��,��$_Þ����������ɋ #)��WE��0�@���:�]Qw�W��}������Y��}�kq�c�O���	��m��|����W�ф�4iss���L�]4fQuշ�9��R�nC1��dfd��%l�C+pA�R��͜�0�q䬋5��6�d`�b
õua�tO\!�MS��q�7���/�Ϡ>�1������ȏ|�Ri|p�	�2�(�㑷$����û��5$2 B>nHc�l),�)���!i@��~�4H���kB%i Pm�P<餓h��B
�^<��F@�����i��ژC�����k�N�F�T�X�g���~��\C���sΜ�S{,n���݉ק��[��iaO�An��V�r����o;n��P`��k��o����uK�?#g'���x$���Ѓ��Z���k�*���&����T��]0!{�Yx���V]�f:f�;�P%v���r�1����p�W�M����$�o�A��	�S��W$�*;r�"w�ل	�e�Kx�(�R����^%ܑ����yڅY��uL�^�g����Gc�Kk�E��B�J%d!<��xv����:�mO�xWMo��`��y���4�7Ij�H?gF\��ܙ�Þ\� \�U.��ۮ+C{��A8��s�J{�&H�vpЊt餅4AI�IE������i�li�\�4gE�i���qN3��ǎ�f������pų&�����g��@&;7�r+�A�=��_�;�Lߞ�a���a���Q�
��6�wj�C�f�3A�'�2~���H�������v�W#]�X*!ugZ�Q��o��m�^9뎏�JOٴ�*�L9�-�h%�:A|N�R�W�ܑ\�}r�zy�c�f�F�:���`���<�F,0b�gbP�
��5���I�(����lM`CG7>jobL��s�{;��Az������+�m&C'��5ϳ����Iv6� <��sX���8��M*a�4&ƊO�Y��_��{��)
g٭L�b�朷�� ;_0�<��>�{���4`L�����XB?r�'�e1��y��+�$��<዇ڌ)�Ry��&�)���tRm���EVW�0�>oh����F��q���g�q�͋:\��]��)�Ч�O	�����y UM��X�p/Q#�~��,i\4�wM��լ�#G��a��0�ʂ�&�*���)@�Ŀ75��5�<1�B^c�.yG���ȓt� ���ه�|����]yp��p��Tn�RO򱈔;���lQa��A�~!6�2㹠�6��m�嗺����ԇ�vP�����sx�)�ؿ����<���(��������:��{����/:����tU5R��歀cۘ��3�'S�!�����71wf���b�]%��屌����������ꃛ���~����W3ؚ���<�b�����Ơ]�OZ;R���>��>p(�.��v���G-�r!�`-챻:��r�7�E+���rJ�nb�)^»���Ϧ�kU�yց���<����Ń0M��|��}~�s��ƲM��N��si�R+�WM��ܘX�N}��L��Y
#�X��h1J���K�{���z^ɖdwW�p�0�h֎k�JG�W#)\
5���v����n俐���|l��,����nƆL�u
�٭��йF��BZ�j��[y���s�L�t���fŤ���tM\ލlָn<j=q/�n�	���o��j�z�.tAf�>>�
n0� ��n���nԽ͌���XJ�I��bn֩8b��&B�}x�	�����y�sW��5,Ly(­�W���X��R��P�?��^�w�C,����{iK��T6{����>���au��L	`��	�j�(�K���"���M�dx�ު�c�u�xp`|�y�_���0�e��Fw��ކ�G'qCƒ�goP�la;w���s&�C�)}���0��P���S�I���]�4�� Р�\�8Z�4OOӥ�WAMץ��s��P�hv�����-;�|G�>��q9{��]S��L�o��ܯ�#.�����v�o)�=QLkP̥�ƌ�ԋ��F�܄g��.�}Y�,ٻ�b���p�����j]��	Mv�]����%GݗC%�morMm���,�;�ij���#�e���|�|�3�=�	�bA��bC��|H����wKP��~f�t����v�:�%X�
sW�ߔj��6F�R=�U���Z&���j��,Q@���zQ��������si~�ҕ��Ⱥ��x ��#������lr���,��]�-�dm0�k�8r������"�ju4r U��^�3��������/�sX	M�ßY���!�2I�٘34���a��2X�$�)�9��x���co�� ��ǝ�@���<�1�w��I���F�d���w]�z�f����Z̸���قioͭ��$!hoC��a���m�ؖ�r|�����9��6VѺy�15�+��Z�q��g{�n��{�1�=ߎ�`f����@ь`y���w%�ςr^���ı���ۛY}��g��4�s��]l'��1�h��a�XT�p�~lM�3�"Σ��Oh$؛�G=�x�w��v<�Ƀ��"Δu���Q�l�;�;֫��T�e􊎛m�/�Ul���o/���-嘅���{M�z��@�+��\�ח�<Bώ���}?
�m�t�V��BHUM�(�ۺ޴6�����o�YW�o�oxJ�ԬcګwOîE��K�{���F];�J�.3czx�k%أ��M��Ϋ�����1R�ʫ�<�k|����n���0�1 �x����}�V�e"�d��f�l��d|�;R�����:-�4&�QG��
n �I8�M�̐"�()���ÐH$>0�P+[f`[��c�i���h=q����G�1�y�; u�O�i�=��L�(��Zٜ�H���|p�v�x��,;i����߫��p��Df�w�=�gm)������(��Y#��`8\(�.�?0�/�A�Y՞���mx�	��4u�[ͼugk�d"����n/J2���5Q���}�퇘\��7�WG��3��-M���8m���dp����{�Þ�F�թ2��N-�[���{.���v��ٝ.z⟭��8b�.�d�`B�	�5ڗ>�M�y�ͬL;sM�$�>�I��sS�l�	K����ס�sn�i�0-#5\m'-��&��p�^�������	���(��X���ܿO}���3�%�\��O�M+�m�\lY�x��[ƌ뱷n$����߈����"~�O%v�TC�c�O<ÌS���zm;Y���2L��Y��ؑ��3���ܪQ��e�>d��ʚ� A�����~����'�<ܧK2߸��ACm�Vuo��G��U��	$���4�R>���,����P2�zfPZl��V��b��p��zr��r�7U�I_�ٛ�J�/�zڎ�u�m9S4�_qW��&o�(ۊ��`�6���Zޑu�������O���H01�,��h]M�M�4["'q�ݠ�O@�F�Y�`>!贗�<vˆnS.��8�5�Ur�Ѓ!u���9-i�)n���xw8�Ω�����ǛT��3��u�f?>st=�����=}�@l�m-@�Ͻ��[HX��"�S5n_;�܅�M�o(_�G"��̍��o��o�A�<�2)��i�{ϪTp���2�*�ݞ�F8N�'��X3����z��c�@�g/���ӳj$�25-G{a�b��k�TFl�-�~m>�51f0�k��y�g:{�=m:����Z�`{WNg
�>2Tc<@.�֙������q�Dz�^O�J�m5��"���;�Vf�O��,�˻��9�q5������=�gKq��q���}1|Q7@��-h��ݎ�2�fp����Y�$�OG��rP��8A������}�W��<�=�%~]���m]���j�r����^:"�e��P���%���:���c�&��{��;9����f�ɞ��b����2Ǭ1mdV�ΟE��d����%��2�S.�]�����Rq��e��81sٜ�੯f'{�F;#+l��C$-�uv�r�
�;�^���Y8��O8u�2�W5��9e5��gH\�{ �q���D޺ǩ����4hx������6���YiU �
Ώ�j��|�� z��2��v�|���U��5���A��&;��&
קGv�o2�d��!�s1����z�`�\��M��R�*.V���w���8Ӡu�X��l9Kj�[8T��������T���N��Ĉ̩w:[[a�;gU��3����.�'@ȪSCTS���Ԛ+�8���7nM�}/��!e�j�KB�u8a�nԩjVZ�		��x�#��uؚ��w�]7}!�%EjBp�2欮��KT�ԭ)\�^*�V&K1�Z%�<@�t��֪-�L�����f���x�3��o^G;n�3kn7���x�����\��/�	�5���u)u���R�� �Ù8�]��M� ��8��e��n���]�8?>j��$ܴx��u+o�U�3a]��r�'7�+x�ժ�WZ�8�q3
-�Iy�>�OO
]eo�a�����um��������_S�ҳ6���3�9��!�	�{a4�&�m�R�* �!�dk@��D5���6cpBM�����*�z��_.4�K�MW[l!Z�EJ��kI
�rzJ�v㐯���	��T�h�� ���TX���*6�L3B�j�%�w	RQ�<�(^�p�0�-z�R���Z]�\�w��e^S����|/#����w@uə�<S�2z%yti�������6bv��х�RV����j`�ܗ�
��#n�v��g�1[��G
y�rڛ�����N*[�k�9:��J��N��WbO���BFNZ`;���%o-�Ӂv�.���ҥ:�ܠ�^v^�(��.�kK�75�7��"�Y�7�J�&S6%�_��X$�9w�=�b��u�8��Gd��2;�WkP7�fc_L�v��]kbJ���o�Ow��%�Y�Ռ�ܡҹ�SM ț�R�Ғ�l�PY]�b�)�;h�fN߮�b�u�&e�qP�/��V+A�@�N���/����+��n��M��(jkl�����n�à����Uqr�:cYu1T�Mu�
@��8t��c]EJx����3���ՖN�Gp,�Y�k�;$�)������.��:�g_-�8��������x���˽�M��fM�Z77��P��A��O]�i�췳VIǣ<�:� ���5��ط���n�3Z�����|�3�r�����Y�&{aY�m��s�o�b-���Qr��͒J'��ɢ�6�w Z#��$�U0�K~1�M�t������<}�z�Nv�dw(!;
�,�_"<\��
� DI	$�zƝ;x��׏x��z��N�l�?v� ���)��i�k����B�D�L˖""!��:t����Ǐx��z��M9��/�Iu� ��y�f�""r�c1s䎞'���C����N��x���=z�����GkJs(ɔf��N^]��"�nF��H}��^�_��������x���=iά���UQ���iG��Y�g����h��$�! HHHHu�N�=v������=�c֞�dd�#'eA���e������,HJ�"���UZ��Sםً
t��Ǧ�����;d�&)B��dڒ��rz�Ac�i(�����~i��HB��'�ŉ=m��t�g�TA;M�"C�//!x��ˠ��ln�!+����q
ʩ�%lӫ.�f��hZ��VW.{�ܣ���0�2P�5[Ta=V�e2��&���#S�ڟ���1�K��X�It[�z���Y�/�����9�����c��OL����p��e�.�2�Ib15�����םi�'%�ie�t-p�p�)|�7`��6��,����ϫ[��� %;��8���R��/6kes��=M���Z9�O� }�}�H��ʼ����={�U��/�5B��v��JA���f߾�p�`���`��_��^%�<��e�Ǔ6�JEt�M�@�W6�A���[s�2m�������7��//�$��F�0L�3O4�P8���͏o�/9q�=��Ucf�n�1�"��G�Csه`8�Ë�̆3��0;v6���sf?
w��������Vr����ܡ/�.�F�cCXh6a��iMb���.\�J��\�ں�ZD��[�;��6zq�����T96�)�`��"��%t�a�v���D���&ը�*�e��潑����>�1�Qe���<�<�,O�bx�k��g�zH:���ݴr��-0B����>'2����^�1�Mhv�C}�|��s����U��w���bXv�t��^���·d�k�U�bL�ׯ:J�7]ewn�6ze4�H�Ѭ��h9}u!-�������#�<A O��{�n=����%��o��x@�����$��f����S�OS�@	�!�����1�z%�wB�U��ǃM@�ẛdS�����5�K�*[h�[�l��G�Z�e�+�pd:���t�f�f�+�$�	��U�$�G�1�T�����( _���r��c)�����U^�|b:fv�^r��Ȕ�G[C5l����o�X{燾X�U4].�����I�eg[]����dK��ӝ1��x�%Z�]���ɖ��,�?L�7էh���ʸ�`�魰HH>�P����]$/�X��~����w�?���%��f"��Ŝ��Cu�����B�x0t�\����}�������lYӛ�or"M���+�o��b)��=L�8��C��>�TY#%.��c2����Gm��o#s!�����/${e�Ӳ�vH.O�LwX�Z����iL$b�us�j���mMp�OO<�f��7�Bz4��0�rH/a�ܚm��=}���U���~2�.*\�;A��؁����u���z�C؆͆�4uN����V] ԝ�{�
D���#�t{��F�ͦ��nQ�)o�u���39�PZe��}�p�r�nO翃ď�<A$x��b���6�P���"A�[�T��s�g0�%E�!q*�!��_��� ������!�&�I"[�$
����~�����C�nrTj�/��(�8n���no�=ͅ�1��*�G+ݤ#E[d6ߙw�B*{#���8b�{�K7��3����I�m?X 5B�g���~gn����=D�Y�>9�aS��:��T�rMp�J���tPn�9��Tߟ��p��1=����ݱ���m�)��c�]���m=w����6��3�o5�A��x�i�z��V[�4�B��3��/Og��'�Gr �Ŗ��<S�톶j�4Q����6����ҡ�W�\m�jI�?1^�~x�/d@����x���<q��a�ח|����I��M�/jf���Ҩ�I����L�FK�V�/���AO�~�����%�,��-/�r�kZ^��e�l-�I%���}I��~߬uXІ}�:�Ok8��g3&cr�t�1���њ��ԃ��{�\Ϻ%��b��b��@�/��eY�������B?�v�7̪՚�{w�/�
��Uc3'1�s��6<v��V2y����$�"��{��>o\�,
nc�(�A��n�;9@��n�٦��k��ɡ�}q	��=��4�� ��Z�f�w�aa��X�BW���y�r����˝���iC��[>V���N3S�FK��=m� ���W���~w@\��=�]Ϧ�`+O�~�/R�.��[��^�O�{�@���/-�<.SD���3��3�X�o����g#bI�p$�o7/�W�{y��
5��e���N(��WN	F��Byʾ�շJ��c���!*�%�0�~��T�S���K�NI;��2�ӶqM�`����[�������Kc��\�Clț����t�̏8oDCa
e�M�TPH�J��M�zۏ����s�os�zn��uϐ��ƙú��-�N1��?z��`�n�t�"x�/SѰ'W@W}
}��稍z��Xbl�b.����ǲ
��3=��l����ƽ�.+(�bY̖�����wx�sX��^֘��9C��U����\~��	O����=�C��h�pBe���b��7x�뽼�mUe��d��Nz�,Ɋ��Ư{aܤ�>�z��u"Y�p�+6�Z4���{ɯ�*�����gS��fS�Ľ���_�5z��|����2�����q��0��V��P�{�%�>�8��N6)�g#}b\����(��Q-Mk��c�IP��Jn������i���ZDE��+$��l�Ľ�=f%�U&r^q?vP�����aK�YCV��g���Y�m��g䙱����SWL�w<>k��uV�ɛ��r0j��]*2;�e3��b�RdT���%�����ş>f�fK���������Z=K����+������q��BT_\Ҁ��$g����S)�CZ�B� �������p/5�f6F�D�L�IqsT��O��z�-!ؤ��1Y���ж���,����u�'R���z�7[<�7`����4���uzy�䕏d��	��uf����jzT�UL��8��Tn���<���h���kp���B��{_��-�
�˕:�������f���m��"e�bџ�D���뛪��鰺���)���`ڬ�����=D;6������h$����/C|�;��(��y�D�W<��d��DdE�)�8sb��d��T�޴�����y���CG�#ɠ�]��R���d}^4����ѯ�Q�^j�{�C�K�GY��'N>��X�y�ϖ��5c;\=�n^s*�-R�L��ͬz�=r�X1�r\I��I����ߧn�E���6����05c��\:�����GR���S���)�y.��� �T��w��k٨�a۬��M�?g@�Ǉ��]1������>���o�{�3���f�����_����{~��Uҗ�ȹ�>��^v������5صW�^�K�5�7����Z�'���׎hM��\2Q�YM���=��SG�z�e����,;���y�V^`�"��|N5"����W�{�wra�x>�ba �A~�6#�x�v���*��:�T���VU"م�g�w����JPdNB�������ك��Ml^��P�$̎��l$�%Gٿ��|=�.����ׯ�b�=�ך�����/�m�4K+�Q�>�swWm�O�/�'$;$)k�3cy�����q�Y������Þ۝�NU���<�Dx��G�� �Z\�	'�E �B!6#&G!RR9�:ۿr8����i31"A0��G�Ȉ�J�A��L�C	 AD�&5%�d�P��}���N����!�[��\}j�,�6�`HW~�Ʊ����!c�~��3ƫԷgw�b$?`�#7(�|I�Zex�-�j�T� ��5�m:�7v�dC��}��Y�L�l��� �R�=	���<�aܶ�.��7Ys��6o���z2�x�]/�X��t�h5H�D�]\Ñ,P�r]��D=k������t�W�_ofק�=׶��ܧ����:晌��c]{͒ws;'���E�	�Q�{9F.A��uӛ���������rЬ�Z�m^O����}�<�6�F���&0ξ4>�T���8y�]��y��I���~v�Ⱦꌽ����K^�������EiH޶oO��2��!u����T'n������)��hbhs8S�X�2.sv�l�j)]h�0u���ԋ�K��z��#�R+���C<�1���hƣ�3蠂=��IA������,��}2�Vu[���7�3sm��6�tӴ�y�������Ń:jP�j:�w��>|��Ӽ�;����q�������R��ën�x�f�O_su�Ͻ���Z�j���zb
����ٰ��pgc͕�řO����٩f�೻L�4���V��#l�C_+�m�Uı-Q��0�A��彏'p��忟�r�۝N���? ��s��
=kIqw-��vo��hZn�������\��?�kwf`��V]۬aH��m�$b�c�dC�Y��Ng��-x10'�a��,{��!˝_���	�XIƙ�-7Ŷ�e2��y����첞������,��w0��v�/)@���m`继j���ު��6%�Mٞ5�h�n�³^����;���YxV:]>�	O@�q�F�jz�5J���a[�f3gtã���6m��i5��}۝�Ńvk;��7>�8�ך�-K��Y���JG��U��Oensտi{�9a�O݂?y�`���҂Y�R��ᅟ=fx�&�M�C��p���Q���Fo-Ja��a�pvkhDj�c�uk���%plS����/~߼9��~��A��7�Z��ݗ#>LG�nC
��a�o��7�֧n�����cз�"�'/1�9�$[Ͷ|gg��z������@����Z��*6�^En�i�w�ޜ�ja�a�Q9�R�XqXC�l;��}�$qY0�����RܮB��l���Ѹ���4��l�s�w�>r�-!ɲ�/k{uK�$��,Y�6C�3�,�30�1���U>ˇ
H��F ��E/4�n�Rn�s�;Q}7oT �=KdU�ҷ7� Z�Z��c@ذޭ扩�譆���b1m?oe�oݨ�u�hl�.x�U�S���i���Zʛ���f{�6�$ޑ�>5]�k�R�'{�܄���<L�N��Zg.Y�ʽ���>G����N�<���~D�Q��}��f���2�gl����򥧵*.�ϫe���~����P���O���nËZ)q�n�̈Y��ї\�PX��JU��삏�}0ĉ�6lc6�i��r��oI�
 YDx@�]Caoz�vΌ,2�j实���t��у��dn�<$|�Ǧ*�g�~���q�~g���{��0a�$��k@�j�Į:�u���>�|���i�C6#�!�w�ţ��{Pj�i�n%4�����\��N��AwR�� �\�45�1]D,w�5PIn�ir�ga���ܝ���_���ZՉW^�K�<���՞�����~R���doT�x�Se����n�g���U����r�N��Uwx��)/⽡Ud��=83��-�k���3����>�Ƙi}]����_.]�� �+��Y��9��z�y�?6��7[�ȷ��7�(��֓��ۺ�a�_����}l�k�FI"�;�.�%TP��q��9��ܞ�m(�q��K�k�'M��m��P�V���'{�!����`7$Xr#�F�+�J�,��EF��	>�}��s��<�1�.{�9�O��>��H�[`4������D��-#�ɷ.�[�n�`�w��RAfم:,X�K�+�TSm�}֩�'Hٜ�찟j�*���Q>�����V<���\���\��έ�B'�y��
�+{��ְ���D����bC��ƺu��pͲC�eC�`��&�ھkzU8�u��맻N����)�N4�^bȬwc��np���s��a:����������Hf�k�j�C�y]�jF�[m�Nahc���S��K	WEXk&�Dq9&u����nbK�솯uvl6es�l9�H���gkH��r�b������������	�}U�kuRh�im\���Ȋ|���7(S9n���w�@k������>ime�k~�ՂŲP�Ef[�I n��5��sm+T3.eP�sF=B�;�-�����/�Ry%��W�*%N�P-۝/p�J�n�3�bOvÏ0H�Ĩ��7�r{4UU��-j=���A;/�S�Ml�-�ǈ����y-l�����J*�1z�p�<��4�"E7{Dvu僄q�1���z���w�5�ox���g>b��c�X�G4�ޮ|�6�+���8����[��x�cW�28?~��4��lRŞF�K�F��c�͖- �xX�Cw�������P"p��פ�Ym~��_A�䧭�es1�+�7r��){�-kvZ����J���d��K �;89D��lۖ���5Z�)ms��V;a��m���"	�nl��{zĖ��x_d��
���d�ά*�|�dty!�wy�$�6dΙ�'�M��e�,�Ketٶ����h����z�ɘvD���P����`��w��/9����eJ���%�Τ8Z�W�K��'Cj�Q�3Z��vp���ÓH���N�"�M 6.�k�Q|�T�^oZ̖�Y�P�48���!�y��w���I�5&��r]-7j��P�իlM�h�.�SP"a�iMZ��5d�Lv.���Y�tr"=�..n+����7�t���p�A
�m�db���gK�C[����Yv&+���V{�<6�v��z�YA#+H���\-����؝<���?�d���-9���
�:�xiI|b�u�Z.�1����A[t���"���7�����ܣ,:��2���i�/)Z���%��f��n8�pb�����,^�A}�y�F^r�i��*F�@��	5�f��t7%�t(E{X`�$��M�"�$=wRԈ�PX�Sޘ�L�~F�LzY��}���㍻}x���ozǭ=��$��!)`��M�}d�BG��,'զx�">�ۯ_/�����Ǐ��z8��Zz��*J�H�6�E #2"3;TD�"�Bl��(I�$�=jԄ$��I:�ӧ��z�����=�c֞��%2���9U	_6���$�T����l/i�)Q2dC&���o��_/����۶�=z=zǭ;s�r��jB\�HBٓ}�N[9$,�BA�T�D�$��}i۷Ǯݻv��ǣ׬zӏw*H�2�I�ԒD$�����Md)jH_mӭu�n�>6�۷m�|z8��Zs�[<I����B"şRh�*�RB�6�R"x�)Q�BA�F����$`�����2�˖�djk����E@�O�e�D��*g��:�TX^\�e���R~ږL��kfT������_Q��f���q,�M8(�5��}�w|a�' ����WJJ�$T"LQ&I�#	F���[d�Mĉ1��RY$�ى2�"B㉘�����H��m��#���	Jt2�mu�j�5�^7��v�Nf�V�:on@L���ȩ�m���{�=�ť���U�)9�_'N���;wm�Nݶ�w	���т"�d����C4�m�Ez(��E$D~(�L���LG �D�i�}m���2�e3J�F0ہ��bm�"���( a���f[$Yq ڑ���"�I"�m�D�^���L�!	EUQ1�ҠӅ4�q��A�7q�Fӻm�m�e�����צ+>H�Kr5�a�Zh��e"	����b��|���q$}l�-7��-B$���H�
�@�eF�d�FY,jzc��C}3c!�S��u��8�Z���2����[2����z>��zܞ��Y���a���n�&���eK^����Ǔ����yپ�cm��&46rq{,�b8��P��~���\������Zuз��5Kߨi�;�P��_P���X������.�h�Ba��6o2��m��
z:�G��n��+��f��y��2�I�c�	��kl�K��U�1 �4#S��t�[�ϧ�����������p�]�����e��H.����5v��bR|�g+�Dٻ���u�4�9���ж��yj���P��Ȃ&)���#���-bX�d��g�	o<@r��R�B����."�Ǯƫ��lÙ{�J���s{U݌���Nܾ�6�HX�Ff��t{{2;�_�6|X���b����oS�����X֫Zh�*���]�3�w��}.�e�;u�\�/�wvF6����B�ns��).��[8��Ԗ�fA�v,�g���M۶�Ndn�s�1��+/�]ŜjV�1\��>�^[�=����G'�J2:��[���2B�}��{�f���,Օ����P$�G.݋����O.�����E�K��Hwm��J��-Z@�ŭ��w�[q}$�x��WV�iylK��K-;ͯb���To��P�#�6NǶ���P��좌C[�n��=1�z�}���4潌ؠ(�\���Jc������q�nۃoT�ޛ��hC}�-�޿��A�8�C�>d���e��g��7M�eO' ���Af��J���G����!�u�J��eU��:��ۘX"�܊����	'�@��\��4��A�XY�mi�A�ϩ�ĉ�~�w=D�׌~}v�������Ҕy�#9H�������c6�K{~���q������� ��0X��LLn'�f�8ѧ;����([.��?��Y���6;Wa=
���D3(oy�~Yt!���s-~�uRttG�����^^�^>$���O�C�v��[��@�mH�	�pg�:�.���K�`���`�S����`�q[lS���4?WҀ� {��=���kv�ĭ7F��߅�wH������ْ�K0-�^��n6���@��W[M�u��b�p�����鮞ᤓ�
�� ��P�OK�ROm�-�gY��]t�.�9f-S�]y:�5DB2Kd�i�1�/]�F�9�N#�sWW�<syJ�����r�m�k�{`�I�j�-��$�b���"���4���m�Xdq��E�_� �́\#T6���WYF��U��w�<�Ը�!�SA�U���6�g^=�/V�/�3T!�����!���>�m�bIIF�w]��%;+jͧ]�8rҖ�^�P&�D�zc�����V�3ln���D8�ՙ~�2����=�qU]���~��S�������C����>�nk�NKc��p�_�=Y[Bc��jjuR�5��n�?��6
�F�b�V�$�ǶN�اC ۬	�42��ȸ�jw���V$��h9st(�ku�=ʫ��W�6����|;ݗ�b��r����zn�6>��lM4;�{�o�}(q�| ���#�<�U�{I׍9��ӑP�p���þ�o�9��"��� �>h{�Nu㑎S�K(����5�5��+Z<꼣��Ov"a�}c�dS[�,�]�q��34"!�31xo@�����v��<�V���eO��<[�<LLn57��n�T��;������.1'�E����ߡ��Pe�j���u�䶄���yt2ah�7cϓ;�)e�$b��4m��	��8�>˯�U�0���ޅ�̖��wL���D>�P�}{���s8;�%�k�����bS]��6���m�4-Ww
���-�n������4�l'_wU��z���[fD���[i�^ebO�s�\ڀ B
��.T���?�գ�Ѳ�j)S��	��wv��G�+�cp*Ok�l���깪sH7P�V�mU�zH*˖l[���2Y�F^�k	�ʧ�2ܺ&��<񊙝|֦Z|;#5<{:2KN�O�B*z�1��VQs��sל=t{4/��p7�L��M$/}�n��w�<i <H�?#�2�,6ӂ	j�ڋ���B�g������Ӹ�(6am�5"�!b"�oѴ#%�P
��KnF\Q�(D�JHdF�>(2�������Q��w�1X
�=�]!�Ǯ��t�7�7&l��hF�\��?��G�gH�-6���\/wi-�E٫�Wܻ����e6�?{}]�{"�����ծ+�T��>oj�%8I\&�4d?0����x�e �(_��	 㞲#$0�u)����{֜�a���mm��L�r<��/g�-��і�N�6R5��@`�沍wp���\�M69�
�S�}�]���!�;\k\�ɾ�`����;ﺎ)es2.���9�P�F�Ooa:#�b�W�q�ks;���ul��#'2�U�!!�]��5��%+~2a�	4/���?0.ͣ�t��_{EH�B9L�m���}߅��N��ߤ~��� ~�oS���_����ޟkKK�osR(U;6�s2-p��zr}����_� {�X2�F?f5�Ec�JS�L�f�׊�p|&�Mՠ�:驪x�<{s!�A�7cvH%�� ҉piN+��9.�k+_^�<�f��d\"���%������V�`�iQ��[�6+�W2B������<nCֺyg��T�weE���Ueq~z���l�F7(O���٬\]�n�խ/�H.މ]��!�	h� ���r��T�F�Vl����iZ�=aOZ��eɺ�wWOM��T�6`WQf%���Jk���L&ޮ/J3�Jٴ����Bcz=�t��������%ٳ̎]E��V�g�S��u�B�5�n��B#����lu�z�6W�ƪ�#*Iw��+���7'+�Y��Z����q}�ˠm��	5V���Ͽt*0�4�[�H1H9.1��2��-�����%��xw��+�ݩȻ:,3���~d��2���Y�P+}���٤.�v�5g"�Z)e�<�OW�7� ��yT�O�M?d}Z�*�W �0���C��縋{��������`M88����K����X{��oE�Y�^���?()\�yr���߯S&��'����$�՞�ٞ�����Ur��R��ű��6F�P��^`��;f�pʂ�1Z��eW�fѮ�\��O����<�M����H�?���_  �r��{�vN%e_6|ElK"�s�5l�\��ƆΏfH�c�mO�9��x0��!f$���[k����@UV�%�z;C�:V^Q �c&�z�kI��<���+4{���,�c��raX~p�'�.�(>h��P�$U
�>���x��믔�G�3)��l����ky���^�~\�GQH�P)D�6�:���\�\����K`��ig�-�^�M��+�1Mm�&)��*�s⁵
=��ř�g���Fhމ��ڔ�x�����g�nǛ�����%5Z���SJϲ.b��b��],f�[q�󁻭܌D@w��n<�f�/b����%���=���g��yX����.;� ����:�w�Tj�W�X�.7G�k�vk�wrs/������@H��\�ƞ!��l�<�w�u2����̖�L삆^���OkG�*-0�q�Ne�W�+>�����6҂pەʅ��B �a����fD�Q�jV�e�c��]�[X�4R��^D;�FXn�4wZ�,��:�0w`�'+s;}��" �x$<P�y�[Eh�l�r�Q{��A��$��S|O��Sݛ���;bb��7� �;ɶ�Q��JP�z���ӋD�?�m��f}���#q�Ń�k��zDU�
~��&B��
�T�r䘇��'��Qo�qv��.b��N�6���f__��p!�-򧢝kK��8a���u�6A���}���A�UآT���uz���9!x�)�W�8}����Z�y�MA�ݖ��Rz!��eUCP�R*�$˵�o�
ְ���ޭ �����k��V�v�W������7=N��-`k�dN���nGWf�uL�zS���\+vV���-�5ꤊ��z�5ͣb�����hbʚ�NJ��{!6���{���ە�9�fP��Y����yR���qH=��-]�g�E�+hEc���wVW���nU�GBQ�V�Lϥ�1Y�~7��O�iq�;�[��������ڍP�N��c�b���/{�˅�|[zΎ��L�t2�qc���إ�wW��zƉd-0��N���Nݝs/��@]n���v�'����!IoC�գ�s�w|�[�[�j�J����"�A��?ܑ�|Q���;3?b�Udk��	D��I>-�Q ��N0����F#%"\�/ �$�v��$��J�=@x5^m��g�M�+���k$=����9��wkT�@�F m�{$m��@���S��M?u���6  �R�O=�ê/��\��59�|�'���u?���m�ړ���j%X�ɧ����Ɩ��g���˕�e��qPs��c����g����ђڄ��	���*��Į.�+  �G����cq������~������	�>�}�}w�� fc홽jC�zm��!����&�� ����%�37kUǢ����-FO#��*:!dxx�P��#�ٱ�՞�o�����^�b�' DgM�IN���!�4< �vxvz�z�����za5��#u��sȞDB�l2!�jB�1g��Ѯqg�4H���/l�g�n[����Y
3ǯ^����.�������k[�b�7�v��J���#K5��!��r�m�� �)6e�!b�I�W�^3	n�`��瀄V���Y�Rʾ��,K�o�1���;�<H$x�U�7�iK��� .�,'G�63���e�8-mZ;U4U5?D���>��=�C�M����>��� N���/�&t�Hs�g��s�f������ݧ؇�����6f�t ��y���m��
���v)f�= ̹�����O��,�������7f�����w�T�����b�u4ߩU������۽�%��՘eT)n�'s�ȸ�w>���s�N�TޣEH>��;���� �'�Ld>�]�s��&cͪ�6�m�0��'� �0}���1�����W@��/T����ɉ{{�+;q�q���oh��a���+�H�$�3@]xw��?����`�-�[��^������9ڲ���)j��ͧ�M�g<�����,J��渎���ff����;ٳ��:#���SX�;��UΓM/8��>=[���M�+lt�Lͥ��t�z� N�,�НC�6��$Œ)]5F�X�X�)����K1om��s�8he�l	2�0���(���fͧSp����Q��ً����B���Ǹ�T4[Jڝ��,:��אX�����Oao���vN;w�&K)U[
�0�J�����>��^yw��Y�φxݣ�K�r�m�/8d�}�쀄Ű��s`9�{+g3wY�8��KXFjҔy9+���j3�=]Z�姴g=+�ؠ�$��^���U�GK���hj�,!3A3 4"PY��x���lHe�J�s]�a��WV(��)�y"ݳ[�؇E3�4��;�, ���"���6����N��bEf�r^�R�p]=���oK+L��Ki;)�%��ڷs���`UJ�w��q.ʆYr�jGzn�%�q*]ͤ�E6[v�;���ke�u�t��\��	�����[���0<��4Yu��w7i�ӡ�V��$��6N!ͣww��%Ǻt%�pl�dn����:	 R�a-�F�^�1����։�3�;�Yyȴ�p��q:�k�Ɠ�B;�c�8�W9jd���T#9��Y�v%�ME�Q�U�m1��(���Q��*�"/ F.s��uj���r��q�c)kQ�P_]_���hZ��p�*�C�f����=�H9�4X�
��u̜��or��X�G
6���M�N�g�u�/hځ�/�^��.��s����'����=/-�b+L�����3����ڬ�P��1��;���D�s]2M9K%dMb�q���7�,���ucf��<�Xv:�uw�;��qV�
sj�X7�mv	Q=���F�+�UQUˮL;�Y���h��#��1�g���V�d��unt.��Rx�:X��7����I; �0�7�U��&�]z;^��u�n���a�B��%�݅��aSꋓY�o%ʷnVf�a��u��I�\i��+r�sGd`�l��<<9T9*��1
ؘ��&إ��-e`���aZ2�}�Ye�Sw��mQ�}w�Ox�^����i���H�u.X����6T��t�z�u@�u�����Zbc=x6k-���ċ�	�y��Țgf'Y��� ލ�.�Q��ãJ��{sk������eݸ1�k�L/2�<��ܡͪoJK�j��D�s���ujg`���i����u��Mr�.x�U)Uu<��ٛ�o��n�����:7�d�_F��ӽ���.WBW�_ff�J���9M�{94�B�QN:���47[(˾��6ޞ*GW���Y��i��9�1}�	i 	�@��X��L�Dz�d������<Hx���)��""~߷^�6��۷n�z�8��Zs�I!=����R-��t�3v�!g�d������
�$�nt���nݻv�����=i�o��#���	J�]�2j�*�$���	�ۧN޽v�۷m�}�c֝���f�i�/�"B��ˢBTB�����!�R��CZt���nݻv������Α�̴���$#��f�(�"$Fd�4�!;o4�N�ۧn�=v�۷m�=�c�'� �R��2�OK�r��$��Ib)a����N�I�=i�O>;v�۶�^�^����_�T�@���,\���GƗ�
��������BB$AX[y�9nJd�?w�2E�e-�����B_�]�x�B"	P��^By�%�$$?Rd�t�.vȗܵ�z
T�M���",��v�D����~w�^�9���Mђ�5�c��YxVPdn�g�+2༼pG4,�4QY�լ�m8�F���C�΀����bŴlF����͖^�`��ߘmW�^����Kf��;_<�5B쾢�[d%� N�y,�j���0�o�\�P��i�5tս�h��u�.�*pk7�� A��t���٬jű�yڪ�P�=E��p����qK�Uc��*\M1����|��f]�'Y?eÿ�����6X�w ��O!g�.��(*6V�뒘`���wa؊D^�Ᏸ��اmB�������m�}��
�nH���'Չ� 탶�]�Ά�/7	^������z�P|��	lstFLN��9�#���u��|yu����x̃� 4��-au�X��<�]Jwk+\������:�yR뉹-^��,{}w~/[�4�#��X�g8�$�敷���Q-γO���iyW��M瞫)�*���b<�i&�sY��-�.Ɵ?����Kι��U��&��V��UO�Sؠ3<ﯕ��[�(���eX6ӛ���W��=��1_��}c����V�J%��jof�Ӄ�P�{l�<͛�u�hoyj�<�!�o��)F�Y�,�y��#��
4U���2����k-p]�w�f��������R��꽬�}���ɠ�L7!{���r���~���Ntwe��luq����5���|-���q<紱�j"�3�9�{�î�J��h��3Q���:���^�ѩli�����Q�{��]g{k�����X�ǧ sc�Y�ϝ��&n�K�]��G-l��U�<� 饌��Ʌъ�h�dG�+C6d9�K�CV�X�s��;��-^ ��#��k;�q{o�a�_�k��t�	a�^篭f�)��N���O��y��J�Nl�:K�Aբ�S�M�ÆU@m��οH�,o�ey�vy]u���~:�ֱ�N��*�nU�M�!�y�<����i��$�_`�Z�y�g}{�jw��1{��.���U�ãŪ�	r����g}N�;�[��arb��M�<�8t�;8�F���;���K�=ǋ��d�s�*)RM[E�ؼ�������u`��=;��W��	O�ų\��c�ųvc3TS�,�#ݒJ64�'�ڕ�e�G���O��`�^4��]p���x�=�P�{�jG�M4
E��_�k����"�Q)(〙�ɷ��6ۑ��:y�r�������gH�0RdBA?zv1[��5���͖[�E����[��s����ROM�{�S���3���?�w��{��8Lk��-���X��y�5�&)��u���S�3a�;d����M��߬��]�8+���@޸.M��~��z�S6��x���@�H7f�~���� ������{�Ake;�pN��{����I;_NT\Wf;��98ɌgJ�UO8Jq�m�Ǎ7�Q��ќ�����{���M����j5�܀�Glݍ�捜p{���{��׿f�}���Gu�>w�~}��[�w���m}�����\�9���H�ݿ�	����~��!^B4�P( �@�����d��Z�V(��y�����9�X�����Ww��еc�-zt){���l�����|�����+8�v�U���]������7�p��Nb�t�A��뻛�&H�oM���$�����/׾�jJO�ռ^JB�3Z$�e�h�����nJ�(�7�m2��̸�JZo5�8�>{.E,wI���
Ğ��ށN������T�853�}�k;:��UW��䫗����y0n�0���jz�{�-f��Եh���r�s[�Śͽ�]��0���18$j�����O������x:մ�OU��]��7��Z��7�c�l��y�NW�&z�w��tb�<9�-kF$�<۫�A�2�`��J��
Wo *����l��ZW];>c��@C�C��(x���n�I�I���0͚�':�qq]w���#�"T�Dۈ �$_S;p.��=����/�4C�7�r��g�AGn���̺���=?G�[�u`��O9���X�q����*kn�/��}�jU�T�*>���"�i�lUķe�v"�z�)�]o{�]İ,���Kz�(�ޙzi���K����7%匕��F�����[1�݉9���"�����/R-�O����e���)&&�7��X�M��Rʺ]�|�a0�:֤8g8���.BJZ\m,�;��5����ڭ<��
��^��]g,���h_�>D<T>�}��4|ٿ\z�}^�FHKzzn� �O�"�32��,�1���o�!<�3�� ���7��m�@��]����ݮ>�8�ٖ��:h���ܖ�"��������u@Wչ�B�2��]^�L�%$�ӳWpޞ���n�}poY���DnZ��3��9�DĞ˺���wN��>g,	,��'��͞�\�Y{������*8�0���e/g�'M�ػ�kJZ��]@;{ҝ�i��A���f�������v=�.�<��7�;���wQ�eZ'n{��۪I��m��p*:��fel��7ʚ�h���⫧�J����ڌ��}h1q��1��3A�=�l��0b���}�-�)�g�Y$��<���F.��"���^��U�hY�ߞ�𾟍��To�m�*��w0�g�r�j�ۣJnP�t���!��
���0v��9L�.MU��n�_�a�5�<J^�U[��a$4�Ɉ@K9.��D��e�R"DI�γ��Y^!E���->l�w���}�K�����ؤݝ��b�}xy�m9�@�IS�<�A���C��{��ߧ���$
�em�XZ�{�A���å�k��^�v�ԣR7���e*��j�g�������ڙ��a+oO��~��э�L���Q<$^�f�XTu�j� �A�z��9�� �2�b�/+V���-�ٻoX��96��vlb[}P�^l鮞�8�[HmI�r�T�mF(����Ϲ�0v啖�)�,�	Ok�Tup�%�W� ��)b��-imS.z3~^����������Pa�D�_&ż9{�ˬe/=���*�Q�w'<�q��v���{c����؉i��{ɸub���lx��vg����;�
�\��ND��׻���P�ov'��}��y+3`FM1���N[n�֑l�X9�,�r��8�[�}3j{��;@��S�ƣ��gBq!�ݱ12c��������ʢT,��.�Wwe� �M���UC��=J���v�-�s����
+����:}�n�F�:�Equ�|�;E@G/�W�̑���ˢ�L��� <O�^:a��@�.
 ��t�Ѧ�$�=���N��JYB2$l�f	#>)$槓y�M�ri�;l;m��cO_�1e�³��ݯ:J*:��{�`eK���ؽhN����/�C_S��ͻ��8(-����N�{�u]0;W�q�����kݭ�ŭ��
�M��Nt��Ӎ�.��=��ٵ�674o]�j<���-Ӱm����F�P߀*w����gM��3���Uد�ͼ�o�05{q,�d�h*���A�����u��w�m�����BX��W�g�"*��i6���\Û���VA���!t
m$���U���͘�R�9��:A}���5#��<O��7��<8Yӗ�,��ܨ�I�a�7b���"]��d:Q.ʎ�H��HPa$�l�
����z��g�:k�����v����!V泑�ّ=�,�Af��+�=�SF���L��x��Y�]�XN����P��<S�=;������+��ʻ��!c&I@�,$kZc��Ƴ:��mXO]�`:
� m����gP�'��dNnoo__(x�:�&Aӗ��@5�\������U��8j�4V�Ӆ<Ů`���7_���3x��͙/y��n����eѯ�r��2jD�����6�׷	�V��DG:{�<��?vu����.��ʹ�-?˗hO��d��َ�Q��⳰;u�շo}+^�لU�ڕ��KT{c�=�w�Uʊ�f>dR�V8�=S��"֋þ`(3���_�cO(�����oM4SQ�i
�׹�=6��gǫ,0-�pW*��m�ٍ�]r���=rT�S&������;��X�r�|�����6���[^�Z�/��(��h"	,^ǣ�����}���0V�#�����xx�����u������0��7�x�1��clH 	�nL*�O2cL�3�i^��'����eW��1��s�`����2�ν{kHh���>1��,�s�̀Ϲ�M��(�������L#���ZQ�gĹ��~��[gV:�iȡ�Zs�[st>}k�j�n!��6$�D#����^��Ag�'[R�ݏ�踚���gc���5hgP�l��n�.�F�|3@�����m�
���>�|H��Ŗ����'��p)�ly�ƽz^���!��	��P(ϵP%�����}���~�/)C�e�ŔY�6&I�|b���<?jy�T�Xsu�%�O$���]G�-jt�/���)�\>�?OX�f�+*��\`������R�V@ �Qf'/o�K��T�@��ޖ��;Q���ݡއd���u���AA����6������ m5�q4й����ݙ^K�:j=��ُ
��[��v�U��#�nVņO��8)�lv�Yi�&K�Gv�6��{�w7�.m}�~�;�?��������'Yڝ���<?l;�y���Yn������m�Ce����d��[Յ��3\�/��h��[�ُ/�kEu�uj]�븬V���a�2�l�3$��5�z�imay�ta�}Q�&��V�����H�����¾��~;�)5�����10�\*��ՓM��n������G��9�l�,<f�%
�t;�t��7�Y}��d��V��K��9Ңp�K�]�n�Nᓝ���2����i�3E��Gt�V+��~ {����jE�[t����QQgh=����7_q�fi�k���sCtdf�#�i��NeRQ����Z�ί6w}��֫d�s;T�O�$q0�!�AE�n�5�n>���(PUX�',9�����r+ˌV{���M0��lA���0��*�tW�%����7:��P��H`ؾ�^�}Nт��Ǔy�lp�L�/������T̩g58�x�$�x�!8.��ogEj�f|c*Z�z_xw67-�����^�.��D�1z��Xu����x_�+#'f���4�͇��W��@nʀ3��V����Q���4���yֱ�E�٤�]B���l��ЏlC6l�2�/9�."�\t���e�vwQ�Y�VE��t�$��fѨ�wXR�:)��N%{y�݋�%gײ���"�B�	��[�ޅ=�2��K]��8�B�;��
�]7���PfZNh��^l
[0���:ua�uǇy��T���Wq�j���r ^-��<�]��V=�)J�H����u�>�_U�kP{S��u�	n��r��"޾�KX �����F>u��QR��j����ݺloD�P;�.�����y����CV�VF�e��V���Y���[��7��*̕[�e�h��:wj��n�_F-[��kh0bOdrG7�K�R��V���\�Ӣ�de�l=�l�ȝm=U���u�7����0�;������q�ȍU�b�$�ʰk�9]:gKܣ�n�oVn��V���~�G(1�����Ub�y�*����,mMpVXR�-�3&��A�K��`ʽ6M�}YP�M���}�)�c�tu�Rk��}1���7Aa���7����k�����͸�^��VK0�+K62a�rS�+����m��*q]6��
L��]�Y��w DVd���"��/*�V
�H��hhy�����qnXPv�.Ni�$ԥ���n�t�q��j��-ҫp���Ůy�ns0���7���ϭ�I������;�'�ƫ>�(
�T�盲B#h�M�Gi3(�~߽äR[�E��C�'��a
����� �-�;UH.A"y���� I?"�1xE��#�Jy�}��R�.�2�$]V��u�
}/Kl�T y�����=]����G�2�6V��˗}6LKyr�I'�C�\�ݽY*N�Q�O[G^g|��⦨����s�%B�����O��ZQ�أ���o�R����!�������2�Jn�+%�����WH�t�K֦�(a��)��o8z�XG�]�Km�d�J��3�NnM��7XX��Jw%��8*u��*fb�YRu�a�2K�2b51�Y���st\y�,�eW[&�c[z"FM"`wQmwePj\�|T{6���!곲Y��2#��<��lG���%܁5�c�ܕzP�V���o.�t5E�i�.�pʉn��Q=����D��v�vn9Ns/�8����]d\w���L�ܼ=rd��&�K�����Œ�{\�lX���(缲�e����	�	y��*b�2�q�g�[[n�YlL-Ϯ�ͮ숽�����]��Ѩh��t�R�q�h��P���ڭ��*2ods(E�L�˕튤U��ţm�\�3��<8.�V���YɊ���N��h��<Z�g7W�+��\K��H�A�ʬ�#�o�I @�5�e�$)DK�FK�@$>�t���nݻv����J������!i��=}З�y@HHB��HIqq�;m��ݻv�^��fU%oA�H{��3���;_�	/o�]�Rȏԟ�/�4����v��o�=cr3U�[����f�;Y�oI�L��"I�[�i�o�v�۷���~_�W��$���Y
D��A"Y�0�*���Ο:��q��6��۷nݾ�=�crH�$��nK�&Oow�'�ם��� Td���4�޻v�۷��=c0����RBBD�*+�s���<��n�/Zj�"���N��h�,�戰��Q"�m%<d���I��y��M�����5������D%�I��	 ���}.��,��a#yқ��٧I���9am� ���$�*�����	Ƥ�'q��BI	G� �@���f�,B�d��^�c	d�،$��"Ch��B�2Ka�BAFL!���"av��]���B���k�;Gf���X�F�ܧ���l����'Gh�6�;��j<��W��4��I6�H��H� �!B�����h9>���!P$�	��#��&H�P��p9�$�!�X�F�& ����B�A6�p�P$`���M$�C*��
b��Q(|�j D��P�	I�a��FF�Hr6�r"����
Hف�B4�%����D1�T�è�ȠȨ�M}��%��)���M8�'�E�@� {���#�(�I/�㛈B1<I ��A!$c�H@���"	�Z%���Xe�Z$ �wg�H$�Q��O,p�VHQ����JbA��z��=ة��M�Vn6�]R�_;]{V�ۻ	u�㚃���0R�FS{RV��5\�?&���̳mSN ���O�o;�Wf��Hd�����ql�v��V�-�xɝ���z�\ֳ,���n�ߎ��������o>"�Dտ��_�%��/���@��j}wʰl{$�&�[ZLM�V�w	�5y]����^�b���|�0���uѲ䂫�2ϻ���s�|�Q}��\t�o|m�j#sǋ��Z��g��Ǌev��;��֬)c�أ@q���1�5���ϼ:5�ƍ����0n�$Q�O�E��6�*CHX���Fky!cV��R^�<c?3r��U]�V>>��sT�y�Ջr� ��1fČL#QP5Q�JKG�?��D�Ml2�"�)7��w<;Q4f+�r�*�^S�y�"{Siؿ��������3�]�p�����&;��.��`g���ad=���ɼÃ���>(|qxK2g�����Ȇ��of�U?;zv�r�?�f4T�>s�I˭��ڌ������X��@�s�;z�*¨���pc�d��&��ӫ��M7qkں�L�2�h������D�p�I��X�BQ��tD�.m���j��|����=9nL*�`�5{�@4{��lQ����ݫ��}��b�O���Gw>۞�ŝ���G����9U���y����*��5��K^l�����0���[u�]˖��ܨ�eL�ԋ����n�͙����gbCi�E0��NHJ���?�^u2���w6�;�n�(���l)f��U�_v"#0�9s�Aݵ���r�װ&���c�M\�Mř�ۏ"��ï\M��^�q�%�:)��^߲7g���GDf�WI)FJY�:�(�F���&��u��c�g����TI�{�٢)���~6����^��kqFh�h�n[�Lf,k�=�G��Uy7��*	�+J½k�r��/3Z���#�`L̡����l��ήj4��$��R�Dښ{9�wfn��b��O�+{d��U���x��f����t�W�vv��2��m˛[;.7tkX��n��D�}K�8]�.���^qjD�9�sN�ƃkJ�I��/#�W ƴTu���Ƈ�͛����	%��9R,]mH�lz40�R����>y+�#X̻%�r����87A�{��v�,J,&���o���>�LVv��i��	V�P�D@H*@d��}�K�r]9���s��;�鍙}�꺅2xVЮ���z.��Y��%�lpfF�S<?j9����iy�[I���Gg��	R�UL�vz(v��I�FU�B;�����ރ���{���$�f����Ҷ;�̘�ǉ�
�ʺ��}O�||	�=�u��D����~�dw�zq�,�}>��u�|������oOK�V�K�Ȗ�#0���sg��x�v_�[���CG��(>L<�k�mּy�Qܽ�x��*�\ǈ��WJu�b	���]��Sͬ��
9$�	�0���7C�0�]��H3q����4]f�f6����M*9Rk�:�ɠs��tv�Ue�<<<�y��^��R�Q�srH��Kȱ�ʡ��9��'���]����=�͵/�f(m�����A���L�l��q�,��q57WWX�ZG.���D�((�������m��|��F�]*ee�0]؀q�ż��s��͞U(?z7�ٳx��--�җHAdj��7����ӱ��s�vvLp1=~������mwPܗ�O���[!{E�:|��^��T�-R+����Ql����J��+�)F�x�L׺�}y�)��S�)N^Q��5�w�\���4��C?�^G�_@:���zʙ�u��os�/�vg��o�5gd8��|�>9�]Ծ�g���%'�S�J��W�vR�u��ꜟ\�J`g��;���W� �{���Ŋ|�>��x���;Uj���YN�1,�N��h���_����+i~�w�V�p]�.�眕36H.�R�#'gPb��U��7\��o���'��V��<a��<V�ny���d��.jQ��w�bd0���K�ǥe3��d���'w��z�]�+�p��e�? =�<��AH"c�E"�d��!����k�~@�*�i"����QF�B$H � p�c�hv����Mxbm�����|�^͊��</<�{�Wew<=��-��%�x�4�]]�,�p��9��y�jf<��Y,�d����P���g�,�n��J�wu�;l�՝x��B5+�MʜV$��j��q�ǈnz��f��S���]�ڦ�oC���.-�ֲ����v:#yK��CdH;�}��݅�ݘ�V �M���-]>7@`�d�1A�'T�v�KO�-���^�j�����]Y��wb�Ut�执��
�i�}���	��^5�1`[7�����[�Y����9�Ϯq�%
~��{�M0��z0Ӭވ����z���g&͓1Y&����f�|p�X7�V�L��5
@KT=~}�.���?u ��*9�Z{�ꑗ9��lX�M�1����u�Q~�l���{�=z�;�`0�S�9OZ�ۛ��:"��Ų,n,�Р��w+�y��O?7O;=�rŻcer�BB�ǘ��м=�}{Z���w��7�+��H3��wp�1]�W^�R�[���b%���Τ�g�.����,�ia��Q�t�W ���D!'2��/��χs4f~bt� pt�|д�~��s��w��v��:��鳱�ݙ�yV;�j��9�X�`jN��Uuݭ
{��?{mp�i��J�C`�|��W�X �I�1!<����t�m&�k�6�3����`W��'�3S�Hܱ�k�AҼc2����X����7���6z����#�}�/7O�יkiyj��M�;<��8Gủ�fq�pL�CY�zF;3��u#�5��ս>���E"� �A�H@�f.���گ7�|��uT�]y�=�k"e�v�a�!ު�D�Y%+����3�1uJ�은'�GX��Ŝ3>y�hm���Π!��9Q҅o
Ɨ�T��'ў��M嫠3�ѯ�r�8�ڽy�ۖ��¾^[b�#&-�*��͞C���;���}V2;77�{s*nL΍�Ӊ}vv�k��SZ�̣�OL7�ټ�ea���kI���4�v��U�%��-�+k��S��;��m���,p�V>��@�+��J���ڑNz�مf]�\�[^r����0�t�p ��KB�V���*6��n�����!j�PŘ���Y{Ngz�Zo�}��
��c}��c��{pb��v=S�3w��;!�FcӘ�����-7w=%��.'��sl�׫=ϋc�C��
~��-���;�[c��=�!��WTNs��Tmo���po��N�6��;����;�A��(�	?ʹ�I~����W��3��o�-�����6�Tͯ���U(Ѫ����c��3ձY/K����vU�:ϩο�Ėg�2�Z1�y��Ӡ��9 ��{֚^+��TP�%�k�`H�E�i��[Е�mj�y�jז��Z�I�tMk�)����;@H���h��Ӝ �F5Q����F���q�'��l>��3���]�t���Z���V�����7��Kz�1獓oL��8���݃�%����B�-�(:����a�z�Ӛʮ<�]Hۙ����>�v57 ��[�v��B���A|�y��P��.O6����a{�sc���:�*gX)�Yj���
�V�՗V.:�Qu���;����h#�<��	{�����:�Vo��{�=id*P��U����"fm(u: De�\n6yϥ[�3"�m�s�wf�\�WL�*��lA�L�-mɁ[;y:�UͰ3L���4�`v�5�啁�w��_?]����.����s�g�h���/}�V�~K�}��OEz��g�;}~�P1f۷*��M7ս��sv�FUU���=��a�smaP�mv,�;�~GK�V�T���dB��C]��^��]8��]��+��)�6::;����ǧ�@��e4�SyY{���ց`�=:jD��z��%�9z�TM�w���OM�O�G��Ҟ��橭���n2��x�z�ݾh@ܸ8���Ŏ�&ZAl$����W}�^�w���rB������-��8�?��kZ�}֪��[�k����NE�����38t��8����N��YM��k���,cUcvJ]�ҤS:Ό�Xv-��P_E'7\����H��Q�����=�c8tw�cjVt�\Ô��C��'Zc���tn���7��Z�����#RӐ�|P0����?a�t}͖�&$R
B�r��#N(_�f'@�R13��
>�"b&[p����+{��I@/#z�0��:�d�D�̮��ԛr�Ջ�k���-ud6��6�9����;<�/g�\!�������uv,��r���ư�y���v{p{�����Pl2�wZ6�PGL	^zeu(�Z�W�V�f(3f_y��34����^�=��&.Ul���K5��e,��1�,V?5&ÕV�y���妼wQ�]�!��ژ��������Qϋ�0�/�^��U�Jh��Yz�� ı$3j�� '�{�]7�>��f�m�3_�gbە�e�U�pQ�-��E��2j0�W9�Qk+�hk.�|�Y�B���a
!��$�TIL"�$��ڇ��2�=�2��6�_M���UB���MoO�C$��R�=��K��w���\r=wz� ^G�=Yz�WΧ�>�S�oC�an׮W�k$�����aom�/!�NLb;���'��s��T��f��QfQu��S�p���t��lȖ˴�̏s�W��ӄ��];*����>n��s1NYKK1�#��d���X#�>���*�؋(�����sט7�j���Qz��l��uռR��Y��ރ5��xg'�|�Bob-�T���B���Վ+������%�4��߲���8{��sJ�`g[7��z���KnE=ol�Gt�
m�ͭ�	�y��`yL�p-�={K����xM��9�}��zb�W_��� �_`O�����s��T���du�k������npq�9B���������潐ٶԔ�<��K���7j��TK`��ƛ�6�-3��6�fL	��������e��az�s��'J�䡝���W��pLێ�Ł��-�5�wP����s5W�a�$�ަ�Cj��ƗzZ�ۍ�O9�v�~��.��7H��}l�	��Ϳ���3#zAm�������_���UEz��V�����6�F��.N�ft��:Y�z���VP��(�ʺx^3�$��{��5j�5�je�J��k��a�^r�����6`�GV�\�	�����E���ת����أ�6�����Rǽ
����3�Â��gh�~L�Wh(6�@��Ȱ�%ȀF�����bc[���ѱfeH�u\��9uKn��K{���y�f�����r�jf�CEn�+f�
XN������ܑr�4��2����)�IP)�Pk��;Y�g�V2Qr�H���kw�g�nY�1����.P��½�r����x�'���k��I��лMj�zk��Z���1���8=��p�n�V>U�/+X;(M��wj��ˮ���^6Vԝ1d�ɜ�z��:�G�l���"wp-�ǯ:���Y����^ S��cZ�ȭ���8aoz�r�6�|���kq�f�lh��;�+t�I�����\c̆����.%��9 �i�1�]��V�U�g-���ӹ����+�&�e����:f0u�Ep��t�S$�}��r�m��ӹW�p�����Z�qbǷ�rcJ��,��NKUGS�z%!Lo��V�u�i��l���l[�(B��̷Zº����klD�#��"x!D@u ��1:��M#�r�i�h:ʞ$�P�el!�x�h��	�-�>����I��'61 U;C��\U������XwwPC2n>�bo2��ͦ2^:
J������V�="d�Y�ۿ�y{
��Y?�YީOl�L��s�c����|]��ܧ�0�+h�ђ�
��^�5�
���^[��[ӷ���:�V*7�!�-�%���z0�S/���8��4��\�"Y�snS�e|�)����*��碴ч&�eH���N��VTn�3����Q��C:��]s�m�ۚ��p"�Δ�������nĩ ������5>4a�,��ȐA�%a$q��;wz��%��q��[��Eg5j����J�C^W��Mv�u6�a<�"�o��ֳn^[Mv3Q���b����w��T���}�tCEi���z�D�����v$�&]�G���y����V�\{����^`ݢe^cW��u��Q�o7wX���D��t�Y��	�;�S*x���[��J.W}E��ut1�'"lcڱ6��c.��EN��"�"6�-,�C]�i�Ptu0�j˧�\\�=�����2L����go�L��jY,�Yf���ڼU��n�\q9��엽������6���%	9ea�9��R�Q�B���[�J�7ȩD�R�2r:|cN�x�nݻ||z��\_s��HH�*)"̐����6e��Ғf��6E�APe8�N�<z�۷n޾=i�e�~|O�m�E��B|�f����mm<[�d�O7�sΏ5_�u�o��ݻv���֘��ǳڠ���tK��V�,=�v���w4��:G�r�t�OXӦ�}v�۷o_Zc�������U25ʦ�m{���'|XS��;i뮒��)=cN�=z�۷n�����߇ͬ}șK;�zb%��D'�7Ihw���m�I�_�޽k���SZ��u�ӧov�۷o_���~ߓ���9��{��~nA'�rz���e,����9���eN�o"��NWi�{w\���Dy�Xb�ͤ���]ܝ�OVT�a'��m2\�)��6�6�'/,��2$��O$�r#�$f��e��Pte�f��;ޜ���ך/����rG���I�Ι9&JI2!3���kWY���J��!%����YqX6����ɚ�s8��C����J�Z�1y�v��Ρ��^m�<?P �<����<�y��a�zY�}�~����:��߭`�k���Ƈ{V��5>O��C��U7�=��Sң��Tj=�q4��3�[�<dV|�qF;�u�������k�{2���v���s[���� ^�S]�E׽�"��'n{�#�w;�.�\�p��]sff��b"�UM1�!	�Y�!����̣ �����q�}jw<�l��`�٩��>�Kvkk1k�����Sd�X���]���d�[���x�;hJ����]�n{f.	�od����խ��.����}�A�����K.g����%��uyx�S�i��b轡n���֏T��==��������*�nh��i�̧�e�si�Qv��'��8��=Iu�dS������0�D��z��f#��{���L�[#���K��B�Y�x�1��.�J?gk�Dz�7��ջ�E%w�3��*4�DB40I�Ȇ
��+@�ǹ�k��E�νja��ʭ��g�2�l)��Xx���f�*�\��kc���T�;z����j�@��>��wI�M��nrL�_VgK���k��m������O�N���g"�]�}�5V;��f�-�`�i'I�����c�X��3}�`�����$��3U���vn��c��A�"^���'A}q4&>5P��\�_C���6'*w�5��O�R�����qd8��>��v�v�8�Q��^��{��;u�l�^�^����ޝ~����4�9����Ӷz��OIU0Ft-�l[��u\e��k(m�z�F`�����ͣVd�o?�9#��'����-@���5�֔��ԅ�c�^,��8�<�H/2���q=sB<�vr�u����W���}��E&�۸�]�>���q�tǶP#J�ܔ�l�S�.��# <���M&t�[��k��E��$����՚5׉\kP��-kcI��$��(Ӛ��q)���$@_PN�Ǔ0�R��8�JP��Sru�\�&�Td����FM.`5ϛ�t*����A�k~r��V�+S[6��'<�`�����ϕ��@!	D�p�(
	�~LDG���Q*H�@0	0�$�QY�	���󏷡.ʮ��S�
�E�Fofx���'�u�� �j��]M���C��ܾ�ܟw�5'���Sڱ4#����U��V!~�oV��7��V��9۩��[#=�xe�Ԡy�h�Une���΁�/�X��k��a՗�p+�\ײ��׆Q�V��=.Y��ր}b Μ�(�*�>K�
7��t6LGuЕ\�w�1�<V�̓��s`����k2����Dt��Z��<�X�%��f9L��;8A�h�	l5��z�XP	�����g�(ɫ��|� M U����$�8�/Q���L�[��;�v�!E��P_Q�_ū���/+���1<��l;���kԠf�U�w=�|�2�8��ܒ�dX ӹ��V�����E�S�^�5s�ctn�rǯ��\ڗڐ�O�2k�s[Q�{f�	c�	�;a���!�z�zf4�`90ra���Xi�^���f�r�
�W�]�J�diU��e�a�!���ح�����[���Kܧ9���p$zH� x��Y���ڌস�^h�CZ��6����9�V(�j�{�3ܣvs�np$�rU�5z��e�T	�\4T!��z,��[5\޴�n�a��������#�r���K��I�C-̣�m�*;��7-�3�m���%g]#�Y�����̞�XM�I��㩻^#0�eP{��ܹ�׎N���y�F�f4T;�:��t+��e���s��C��M���<��	�䝖wLc{��_��/�v1������ڣs��)��D
��m��Ƌ��7 ���-l�u�{v�N^"�m��(�Hnn�V����g��t�Κ��붊��&��Vǟ:<��շ�$�"�s-5rяWH4�ެ�^��Ɓ�aǀ�T�=�/� z���E�ӉEK�R��l�a��.z����Y8�,�x��`]e���m
��D�L�w�	�Z�oj��M�N�=����	�I[�❦v�c�8��csK�"V���F���y{�d��T��q닩�;���yϩ��٩׻b��<�y"��v��b��0ͨ�]߫��Cf����ޏ&��mG;L'zś]~�m�UC��3q����6��q�<��<(�׋�n��V�靷ؓ���L�x�{�\� �3��kɇ����X�O�{����l�2�(��9T�R���D2�+�g���P����.a_;��=�/�`�5' .���R��כ1�IuTX]l����z�X�,aJ�2��LF��?���5�������û�P��8�Z��T�s��Yޱ���Դ��f������՞�nC_����V.H��v�U�j7ii��n��H�I>#������5��яٲ��WqQ�]���M%ِ�p[��ַ���J�I ��w�����y�K����-�����`if�Qa��w�G0z��h�r��*.���M �~W��sIL�c7�;����G��ę��
+�P�e������9:Q;�͵|�XֽR�9�R�C�������W�Ҿf�e�΅����+>B�uTF�k�ֱ�&r�>� �$&1�s�S��W��v�iEs9g%���{  ��a�7��E3��b�p]��U�\-����WT媉Ԗg�j���ʆ�[�J�U���ͱ=�r�n�Z�@$�����W��0�J��b���i��Z�ϷXd"�I���Po7"(4w�q�p�XÕ	�QW2�N�ˇ N��*xt!+K�+�[r�[����o5��S��� /G�}b�d��P댙�����\�X�kN����>��Ə)�)�`�=۾ؚ���cz���TOU��\��]�]��ѻFX֝�=1�y��4Xg�\]-J[]Mz{u�h�ߓ��F�j�,��5�5L�<�Rwܜn�m��,�@m���sUP�2��O�ij���WG���K�L�D��et���jr ٪e��Ehm8��o!*:��63���Q{h���u�WP�m���Z7K)�Zj�}I��FΘ���MrMU���â;�������"�}(�ԏk�1�y��YҨ�(��oV]�ݝvp!�����"�Z���<�K��+���w�dP�2!�!`�P-�٣E�����]�y�]��$J���&���S@�tQ��q#�
y?3Q6��H��ʡ#`�Q�$�
?���mK?����̯��g����L	��p�bV�-��/2�.���L�k˴����M9W.�C��M����s�u(�W�it��_7�ؽ/�����]�����8��.�ֻ�n)C�A݉����6����􃇩�'���O]�΁�W1�⫢=ٮ#�@˾���[�f`�Mh���aSo�n5�����{��׺b0���ށ*�Ƙ�묙��x*��v���y2��),���ٛ.����|����9���n��#[cy��m�^Q��H\��.K���u(���ϱ55��o3f��w,�AK׈>,�K�0~"u�y��5�[��k�<Y�k$P��M6ј󉟐]��3z�ǚ����M	m�U�|sCp�?��������bӒ����	_�W���|�GZhȶd�olv��O���H����5R�i�B�wTG�q�G�H����53Z����ܼљ-R}Σ �܌��w �G!��&�]����g���B`�n�df2�·�|���
������_��쟂}�J�K	orXoAz�9��b�z��K`�0�qE�)�;��ZH7h�vMcs;�Z Xv��i!zn��y����C2��A��3�c��!�A�[3S��	��)PJ�\~��U}߷"v4w�׷����~��~tY��3'e��#��Ֆc����O��{�4V����FT(���]Mbh�@%�4�oN|�mj���k��Ѩ{�%}�ў� -U�Un;g[R��\q�8`$sx���lCjo6A�I�p���������gnOgW7�r���+_�'����gY>�ݷ�1G�m�[p���w
ν����]�\R�s���Wv�;�i����[���<���'�z�7�*�w�.84�Yl���2.�#
1�c3�,�4%����X�<�[�T[zqD�YeSWo:�в�BP����ޛ�9����4�뭏L�Ńn]�x��<�77���S6]�|'���!�8D#�6�*Cy)�� .·Q��@MV\ي���(ѩ�W�Xc���0�0��0�6#/*���<A��#܌���0l7:������s�졏b=�u(u2�CZ�������K�ú�	�w�%~�����x�(ؓ��ط����|��8k�|�۹�����}B��}s?H;ۊ��
lV��(�ʎ9I�c��^*䗌Oݔ+lO=���O�o`��{�UNc1@��MGBY���)��໒Awz����z@�f�$}���7{�r������Yؤ��{އ�2V�<����ſ�s�+��Z�ڍ���
HJ�c�h�R{��ԍ�캧�<��)}|ۖ~�WUT�s��<%#�ƒN��;����o 3.w��Шew\�󝒷]nN� �6��
'�Q:��RA$J!��E˂H�9�:�7,ϖ�TVq�~�����<OG7�
į+:;f���J�z��/y�~/��':�ڬPȸG�`��o�a�*��h�C�Gd��,^x�Q���2�:�Hǜ�y �e)�dy4	@]̭�ȧ���=|������Y�oy�4ev�@C�R���VY����h�<�m����v�4�J@fg�J[+Q[�0�{k.��$��8�ݮ�\Z>J=��S���am�w���s��;�*߽�:nYF	��p�1)��1;��X���R�$�&o���:(P�:3�6��Je(�� ���W���1�I��La�>�����豊gU7l�=�5fN�?T���e�-�C�1�º����$$�T����U�4Yv�хJҒ�2BG�8ټ�X��U7��m�����+���횈z]s�;��+��
�FCd8�� ^�U���P���T�
�U3W�K�\L����D�t]��7/N48�H�d�L��q�Mss}��k�h���d��/Xc�
���_l�xH>���(�fy�[�a���B���NQ��^��/P�ȇ����'|�r���d�����گ��.�F#���K#'��w��O�����f����8�(��/��?ҕT� *%�F�� �0`´9P��Z���B0��"� ��  @B VF �B�*�Y��"�*���`(�"���@B(��D����	����)�pvElQR��	�TU@�B @B
�@B
�@B(
@B**@B  �B��B�@`!U !A ! !  !T ! !  !�(�DTETAQQQ �D@��@��A��U !D��T`!�@!�A�� !HARA��`!A�A
@`!AT��D`! +H!! DZ�i��@`!D��@`!D��*�B�HA��`!A���� `!A����� Qs���D�PYPHI����?���>�����������3�?�/�O�ƺs��Z��������` ��C����O�PA�� "
����c�����?8�ڟ�g�!�AW�?�}߉�N�$�~��O��?�Ov~_�~A�%W�Т���QYX@�DFD@U��E�Y@VD �  !DU� $ DVE�TaY@FE!a@X���d�E� X�d�`�XEDX0Q`E1��X$���+d�ab�@XE�Q�1E,U�E�V@X,�Q��D��adE�Vd  E�E� @V	 YbDHad�E�@�dU�E�dE�E�DE$�@V#YX�U��E��FDX@X�d $Q���1V@X�`DXEXFDX	YbDXDXVU�E�`�ccaX �V�V �FVV,���!c`�X�@�cX �X@X�X@1V 1E�AX�
�Y`D� �I`��V$� @��A`�EE���EYdX$PY$D AU�I Q�* F� �P�������QQR@DP�@d$�a�+�?����������?#�ξ�]�A���~��a���?�)� �{a���6~��U�����]u�'�U��_؇����}�Z��ua[O��iA��C���h((?�+�q>�G#�a�6�Y�C�~���_�<I ��y��}����>�� >O��A���Ђ ��~��@D~�}p?Ca"~��~ J��?��?���:��<����*�."y��� ~a�?G�4������� ���A��j-O�s�\��
C�O�����)��MՁ�F��0(���1�{�UE%*AJ��@�!"R���QP�*��
�*(J�J$��U)Q*�UDQ B��AR�$P��D�T�(UU�D�I$�Q)R$PR�*�T�*�)"�J��T����B�U$A��%JJ�}�T��@���HJ��U������Q%(�������P	%$AH��T*J����P�*�*E*�QTQU�J
E� �V�B�eVU�5�֩"�5��J�*U��5� ť�V�����l�������j�*��m��5R�J�آ��ԥ��A@"�RUIU���� �t(P�C�����B�F����lhP���t+u�֔�R�+X�i%-��*�U�)d�[(�m��ն6�h�Zjͦ�[V�4�+ckj����UB"B�J*��J�U� �R���iiX�V�ҕ6�X���2�w����#dmkB��ֵ�VH	��hUZmE����F�f���U)B�"�J�  l;Z�dVj��I{�9�QZ�
6�kV�U+R���Z$UT�6�U���P6hUU[j��Z�
�kDR���!D�ERE/  iڨ)T1iP�mKEdT)K
�UT�ԶQ�,�T�����U$��eR��j4�U
��SL�U
����UR.  g6��4Z֬�&�FM0�i@he
M���4�0  3U`@!� в���
E%*J��UREQ��  &�РFV  4F�  �� � ���6E�4��L �UaX
��0@i*�DI�"�
�   �  CLU ���Q��� �jh �L@dj�@PiV !�2��۩v�0ЪJ�H$�   Z� ���04@F�(  �0 �iS h Z�� jҲ� �� E�@%�0 
�H��AP�JUJ �� n 
 ج �0  6E�  2��  -l�  �M� (&�� 
R�  f�h i��)��*R�@ �{FRT�� db*��2M=U�d ���R�  )�!�   BR!<��  3R�dSf1iE�
���R�<+چ�40��Y�(h�.�ڱ��諭������=��栨������(*"��PTE�AQ�Q T�/��?���9�_��Ҷ�T�+2��P��A�w@^�li5�*Q�'����fe-�c9Oq�.n6�`���Ɇ6��4h'
ӁS�r,�r��YV�5�p�YZ�b��g���73a����I�-
Q͎��"R'�p��k�$�m�N͂ܥV7R�fڱ�v*0n^�&0��^Tc!����&-�6U�[4�p;Ɛ[B�����Vɩ E�fm�J�W2࠭νfhCU#�A�'�����-��q�n`Ñ8 E�k2aDݏj�DT�G1�-ЩHXn�F]Z:F����e�J��W�[7�[�i`u��J��*� 7x�H�Z˕�N)�k92׊-���`�2�`kSE�K^4�[Po��أ��������Њ���nϔHnw
ܶ������z-��K%ƛ�tȂ��YD*�
�ȭ
�䛂�dʠn�#�"B�t/7Z�[w�56����Yb�W���hb�
�Ӻ>j�oXCVi�E3����4h����8�<��:�I�	@.�d���aD��0c�i��-|4�^l!A��В�,�U���[OjهD�J�� ��e�%-��"�-���N
��a�Z�Z���ud�˹��A�u�Je
$�K��cQ�+R��[!3K�*�]l�2����`�L�h��������jÀ\���u#PZ:ղfiԲ�;��`�vq\ٮ�&%��YQd�����se��}(�6��MU��cN�&
ȫV��6$���;O)0Nn1��J�\�{2�"�bަ\�U���V*͔ ��8)i�e2����$z)�	+%o��A����p=�%v�Q[��wVf<�4�e#,D����� cy1 N��A�]��Z%��O-�b�����P�\{`�JP��$��\6P" *�K�BB�4=�ӫ6a�,�[Qn�YLoKLK�wEGJ��s7Q���U�n�ی<{@�W�'C*G�m]޴]lϬ���R9$�ߎ$��óq��T���㷖4ތj����O/mą�m	�L�/-aP��;�-���m5�5�-�)*�wd���5X-on��BW	{�sZ��S�Ff���FA�@�Z�e�JL
�v���c]����r2���w^3An����=������ױJ��u�l��EM�X�"��a&Θ�� N$oqY�.�ূ�����ͨ�Ƴt�P)�֐��ۅ�͊L�iM�n�ڰPF)[nKص��5���Y�첪�r�e|T�HEEd����	��U���{m]O�)�A���)7U�h&��z�iɋFL�����o0��H�9M�oM�N�]6�ʭD24�q5N�*MXn���U����tHO�2�u��o[��_ٹgaV����z� ���7��N��u�d�m�� ��n�EM��fC,�1m�ؽ	��r)Zܲ�v�h�l:ځ�W+SZWJ�N[R��vP��]=��Ī4F���;a���j�X�����D"�.��d⡥-�Nbԩ�Mj��]��#2�� �Y��7u֜�"�Gn@,Vm]�-X��[��9b+�fF�l�y%ݩ�sx�����ɮ3e}�)�e��`u�6��<����U���`k��ӓ,a�n졭n@��VK�>U�RJ
�h�ɺwX@�u�hi�',��X�J��7�.	3[Z*h�H�܂R)eAu 0�d�[.�!ѷ'%��l��	 �%[FT"�����'��Qx��N7+(K# T��Z�&�.ev/��0�c�q%Fh��%˂5���O�m�J�ZM;�v�h���8騵Cpi�Z�NIa�C0+��
�kL)f,v����GwS�Z�:�ݦ�J��H���,�D�D5��U�5ݛ5nŝ$�m,̗��A�(l�@X�q3�~B�P���� p֕�(���FLՑvov���93cL^�mV�ԻQ+(M��x����BʔH�V�ڳP�K��kݿ��! �Ay��Y`
6�GAh�CU Ѭ�/aojI�Y��5�`K�-9@�դ��Mؽaei�n�Fp��eS,av�XZ�vk����lj��nR)��%� �A��`���1\5�)��a�X�ڀ��S/X4G�bM����hڅմN���,�g�DjQ�S�w�fa����"�.�R!��ne )m�Z얅]���<EjL]]��k�t�ȯJUb轩d&��n���
��,�'6��4�m�z�鎘�+Nc�Ɋ�U�^J�4nSĎkѴtm'GV-�k)Jyy�H�]f0��ҽ�.��C�&��|FV6c���;iQ�f�@y{I���9.Χ-�� F���9�#,����Y�Q[Ӹ�0�-&��o`Xv�)8
�WL�F ��:񬎵/$á���n�,�:�ArأY�����R�D-©���t�޽Z�ElGrYŲȔB9T���ɦ�e^�h�#Lu����;YJ-�4��Q��� �/.,,z�[����x�%��Q�V`'t9��V͊E`�q�VX)��0-!���X,�(�CPV7��m^�[	���n�c]�����]Ԧ�wRV��n���^⿌�N]X�*K!��#�[A�``ѕ�y�"F��Ѩ��ٔ�S�2ndD5R��������� �J�쭥)ة�kJ��Nꭶ�ƍ��˗z��[D�V��(�� �&l��6�Ami4by�n��25#���P���l��Z������I0��Y�b�T�Ne)7
ū
B$��g�ok t*Z��]Cl9WO*�f����*3$�劶)�3Q�n��a�{!��D�^աDh8"-dF�IV�Ǌm�yR�֑��˶�-9:ڽ.�<.�,YpRղ
���]��̥���k�@^�W�Z)$�3IF��LP�^��\�Da�8��n�r�i`�me�PR4E@u8ѵ�Qܸ�������2���i� �b�W�J����V�L��j��@���e�Zjʧ0V���0b9��EK[{5ZKd�S*,7yѸ��`��!̠���x�5>�nѹM��ƕhݩ&j&��"�Z�I� �̣� �k$[��.ir�Ct/F$v�1�����m�/P̣ZPʋ]JA_G7Mj�����e+b	������d��9z�
?mU�����͛R�k�T��y�i7�%���p�;�SIN$IKkn�U�͠a�EҌ���-�.t�ҏ,m:�"��V��/kcY��-a�^�~!a��ɻa�7p��RY,��Y�ʃ�RYoE7.�S����)Ȣdk����YJ��V1ސ4;�Y��贰�A7`��:��B�:�J����/ww#g4�l�R��+y�,��� �3k�q�T5�+J��o6񫊏�T�$M��F雳��.XA:�5b:t�x1�*�~�[W�3K��E�Fj���x�ʗ%)Z������*���H��{m*X��Yk�B̺5�m�5�����gȡZ����o�G�dlB%jaJ����S�{���m��n�ڔ��I��b���gcU��]�&�BR�Ԇ�Z�vHA��1N��F��;Z��x�hҧ�Ith�X��k�*q2�
��h�)V+uҷP��E+�4*
㺱����b�������Gei���XN�V�{�1#�`2�۫�6%��?��}d\Y����,��2c��ڒi��>�9i���!{��'�`f� ��r���Į�w��!BVӦް�M't�q���.ɣ�bz/猭�BG�N��5�T7G[jY�ٸ�n%D�6��7si�ii ���T�t�j� K+�e�邳FYG�v0���U*:Oi��c���"l*�4�j�V�V7�ک�sv�zO+UEN' �?@��U�Q���z՘.�I\gs2]I��ޖ�X�A6�"6���֩x
�^��Љ�`ٓ]n0�������n�Gz��Ga�jhPT��yxwY�`v��n�'aۛ%��ԲI���fT�rgkA�Κ�I�R(��m�`7FX�.��5m*��jƤ�X#z�bK&"���
�BuQi5O^���6i1�V[�Y��mJ�����ۧ�*Мp���W���7����"�n�*�Ѷ���e��A����4�׏l��wR{��B�ăd�tl��^\ յ,�$Cj)�V;�x�4����nݥ���UWi���݈��hU�ǭ��I,FĚ4l�jmp%%e�L�[��d�X���B�f���9��"F]��aC��(R�w�^�'J	�i�V^bӡ�TE����ot�6�W��m!����RT���@�EV� ���^@����p�й����{Q���VdpԚ��C#R�	��Ki�3/imӱe�S��j��LA�nn�nŬ���E�M�p��+�V��Mۇ�Pyh�Iu6�� 2,����ZR�k3��WǙ$Êh��h2���3S�T�{)�GV
�DY,ʧ&5+9qX�dY��,�.�j�`���-�����F�]	�3Z���{R%H_�@���ea[[�1U�n�:[QSWOQ��|�o@N�C�pY�h�"E7���lZIZ"�]�R�r�b�U�� ��� �P(P�n�֠i}l�GoI/�R��QD�p��%���[E���;�r��Rκu%��#f��T��+C��(<��c�m�����Uݼ�ڗ-��8]g�aNDVF��M�6K[tÊnٍ3��IF���2)��,�����f��t�b�j�%eBC��Mۖ �*�[)Jt�
9/oKsr�ּ���i��44�<��fe��.��*`S6�.£,VEct*�����c{2v�i:Wl+w�m��@�W[Sw&ƉAұb����//�Z2��r��(�j�E,�f�m�Q�PNh��6R ����i`��<�Ѣί����O��r�4���6�vP�o;iֺ4�4���yn\�ST(a�kc�����N`��TL`�z���P\���f�Zb)c9��tK��t�J�eb���9@���)2R�Œ��Qܩ#vpë%��njԲ�4&�!��s��;Z�����*�#(U��A�ئ'ί16��MZ3QOu�w,�]�� �=������Yr�@7U��iؙ�M�*�ʵP)W�YVIEe�Y E�i�W���RH�&,�Oӭp1v�B��lɶe	,���SǱb�`mw/l,-�h�9z4I�X��}�(�S��- ��:fjy=��t�T��͟cۨȅ���t�2��yQ�[��^\-H�]o��w����i�e(@���ŏ7�C$���J7�9j�D�D0d�ckoYD�#�7a��f�/
NHɽ����lҼoF���N�@J����aŰc[B�h��O�Z��A٧!F]��s5��9!���Z@*;�uz���:�H��ə�Հ��ں�2�VS��'K�PLX�R���{���C��օE-$�P��@l8�<#4�M�ħhv5B��]�b�BHk����[bm[?�^�-&����+/)�@%��H7[�sb�(�����J"D�8�S���U��H�â�nX�Vwn��=��jt����H�ip�ɮ ��Aֆ�Ĉ��-�/��Ax������4(�0��gKw0��N���̭hVHެm[� �	B�a��{).,����Mâi�l�Y�L3(�v�0�*#j�T�ز�wq=%-�Ze����ה7)�)�����ؑ�����`dڼ�r�(\�&�m9�D詵��D�����1�T֫vf8RM\�����Z�m��"Hf%&+{���Z1�n�R�zfō��B���3�;U@��Ww�܃i�1Q�*;�(�ະZ�`��P�OpiؐM9��X�ƞ+ơ0ؙxn�=��Ib7������R������� Ua�!�I&�t	F%����N���"9i)��w��~�^%lb�w���Pe���n���ˎ��b�:4�nn�(�0�L<���Y�]m���4��<�.c7���qHӿ��+Zs�kf�TM�ô��JZ�H��m!X�77>�r���5Mc�`��ʗ�LF�x��d��-�n�֋m]b�aT������Lv���wS�K�fCY�GSz�f�*tΕ�t�j嗐<B��r��qKt&��D
8�7hf!�l��#m�h[Y�7%D�M��An��F�א	�=����L��`��jKE�3n���n��T�A��ɍYz8��lV�(eոe^��v5,�5��ˢ,Zu�,�3U��eZ5j;@�1�D�w$ij2r�SZK�idsp���&�@l��@��b��ۧ�6K��y�a�FU��l��>��YwaT��q������I
P�xp��XHE`X���28憁�x�N����z��HTz���.�R����6n�-�(��ҥ�f��ڒ1��ص꿆�L��l�m%W�(�(��F�r]M5v��Q��{70�
Ѻw���e8������6�J��i���ba ���D�-V��Z^1��9t����W 9(�� �j9��-ޚ�1���n����4�Z���=Y1V���7�smjP�v��k�]��\Gp48�a�4Z�
��%�v^E�c��l&�]�b�cѻ�2���R���[h ��д�$��G�"Ұ���{-RF(��=�NX8���,3o2S��`۳�^GP��׷*u�a�*;&��2���RX,�ĭ��v�9�
��(v��jV��h˴��	i"1�˗�e�yBS�+pq���`j��v���)"���M���/Ch�ƄK�XN��`�o5�T��/�+]����#�Գ�������3K0<��i�������>���ja�ì\*>�����ȝ;c)�:�×��X(k�p���EC��Ъ�G��LS�k��ui(��2�u�2ȷc���QDp�9
��4�=�����rg{O"BV�;D*��Wk�V�{a���4�i���S.N���૟N�&�08��v)�֊�4a?�eZ}�)wa�q2p�8�f�' Q�O ��2�R�������u}Z�΃��M`k4Wiuv�@~$GH_>Ħ\����' "��a4�b$��Tq^�Ѽ97�:���e�M5��g��N�WQ�h ���=P}�v��8��ܪh6�g-ͼF�1s�B�]��{Le���z2��VP;�kg0QLG��;��Cymf�b0n��:��)�IK6Y7X ��'h��/�c�|^;�6�L��]���Ēyhj�V�"�3;W	n|e��>�w^��}Si�{�L�S(.�˜����H,�;�E[J5�V��p���5gmU�����)���� R]�Q���
}��s@�ך�62�O�̵����X{謲	�+��H��	첖��ب-خgW^anVBn�S�@�e�|�gLڄ[�ԲE���\B�zQ;(-�{0�F0���"&���^�Y;s��0���'�Y:˷RoQ�?ps��#�Dt��}F�Ե�VgP�i7|�w0��k�G�X��۫l8f%�y]�d�x��s� �͗��Ԫ���.�-�	qQn�"�L��f�ug�`��j���/�$-T��
�v��Yc��C��������׳dm$z�C����P�
=Ar�:e����uܺQi<�R��Ͱ�K��N��D�H��ګ&���9��b��4=���[���o�\=�B5۹��ʂ�֌��
h]��OT��oi�u�ۗͮ��ŏp4b�m��6��X�`�Q�QFt�Q�ԛ������%ӫ[�s�ǹ�Lm�_wwI�OSB��N�:��u��Z�j�7��/:I���L�A�Zf7���;SY�1ڬ/�Gܘ�}�^��o.WF	]��\����xǌ�s�@�ǵ�^�\�h��C��P9v�)����w;i�|]-�6Y$_�خ�����*�<y\L,��'��0�3JV�x^|�B��u�h1u+KӬ��=��Jh�˵��;4���U�����r��+��6ru���s/���Ǣk�ے���x��)"�޹�J�X�]bgok"�X��Ovy��Ac5�^�{�g4��nr�]�zimoc����5������Υ��&�n.��|�;�e+�Ҷ����Dr�jO��˛����S��כ��l�k�z��9�.&D>N��FR&����̖�Sٺcy���|0;KM�^�ۡ���vM�Wre��u�TA�3Fiiγ�7��|�ɛ��rn��Ju�[�� �U��Ԭ:\E`�F��Mz��	WA ���R���h���y�E�"]��],�|���9ؔ���[\WN�T�̇�7ɪb��5�]���en���C�
�Y��j��|���!�ۆ�H��3�@T�iXƍp�#������V�Lq=L�U�n��N�U}�B�]�D�����[��F���C���%�]�
�<��0c����zhM��x��4sx޻*��<�c}]N�:�`�֑/ڪݝ�W.R{������>˓��i�"=&ӽ����#��S�g�s�wj���̇nЗ�kcl�B�*�o���p}��m��R��=�Β.��*}9�y'�
DWwm��8�#��	j��m�/Nf��Gm����b��;:�[���w�\ ���ܐͲ���tF�[Xa2��I]@���-) ��j�;%d��7f�������N��jݼޗܪ�R�z���rVe�IS�p����58�����b뷛���K�6�o^�U�.j0lh�{��: �*G(u�����Z�-�+-Ѳ'&`ox��^Ea����gϢ��GZ��k��YcDUh�ND���z�{2Rnf��x���|�)1,��o��a�#�k*�yN����ڰw�]�� �F��J}���l��s��)�K�k�.O��o@nc���*ڝe����{:r�$-�=�"��g���@��e�JW"˺t���<P�laǹ*<:���	�^�9M�F�]]��\�wI.ay1�=�.�f���A����kr�9k�՝���b7	LQ�7zn��m=z��BڊgNvFh�evƴ�_ A4�!���ucX�2֝�I�a�e�Ɓ���BZ��B�f�Q.���)���s1̍����u[=�mf�6�,�I��V�&�72�l��y�C_R��L�;���H�vݗI��U��h�ԙ�W���*�s�]개}χo+,�J9s 
���k*��I���!&��{�M��vf�-��b�g<,��Q�^҈:�1�91����m�p�*-�|����fW�s4f�oE��������E�^wv��JF�*9W|�ٛ��:�GJ�ލ0Pe�¸��⫪eīDڠ�t'��T���e�ߗ	3v����#��S �}2+�S�4y��[[l��v�Ֆ��A՝���h�_����,݌�LWH�Y+L�I��+�v7���o�x{�l�\%2�o��+���WSF-�7�3���Q���������q��`at}f���ք�r�V��\@�	dl��Ϊ��]��I�X��Bj�y|�P8t�j�;��]���_Q.��ʙ`>쫭�%A���"�M:��ÔN��4��C����E���p�*���wc�J��Q���2s	��n�<gm�m��1�,=Kuj,5�׷eY�&�```��G�t0�7t�#�h�M�#�(7F���A@���`u�c��69�Q�9FX�7�wَ�m�*��K趁]�"�մ�G�kILq���ʩO����f���!�α՘�>jc3F�tF�ǝ���y�<�v���Yj��b�-�� ޔ�+�vb��f>�9� ;��-犕,_�N�Y9�+YE^��W±P\K�����MiŽ�c�ɝ�u��D��k�=����9�߻�	WJ����.�`���̉��L.�n:̕���S�^����5�Y�N�d닶�Y��_-c�ae�FȠI%�ĀU��\�˜Z�q���h�%#����!�05�\-��ؽ--�8�ju_vT�V�3q�wn�<3z�Ӻ��b��TށY3�T�	r��Ԥ׽X�cukq��}�'X��V-�Y�:��F�.�b���Th��'�b�Hm��޾W7�J5�K������ޮT�kHEB5��g*w�Z ���T��hX����O��< 9q$k`6;evۗo:e-/�¡٦b}}>�f�2��ΏN(�F&��i�"�ǲi�u*y�R��P���}�J�+�us�+�Yf�'��o"k����h���g�i�p��[�ILr���~�u�A�����ٮ
�5�ʫ�|V��.�t��6e�T˸�=�>	�s)U�\h�����[[�$q��#SX�Fp|��/�^u ��GԲ��uLÃl�N�'_8�6U�E�«kuI�l(�+(X5}i!/l)]�L����o��Nhs��*>���Jf����ɛf�Vd�d݅&��Ȕi,�Sz.��E-g]�U�G�u�Du�,�>�àm&5�ovsE�����R�}�v^[�M'����)��0�E��j��m��ȸ6񝑔.���ݷWOsjA�Pk���t˻O{�Z�Z��}��z��wML�����sY�
	3zsŽ�Mʛ�9�֚=��w/��n�X�me�!o<ZM]!F�S50;��h�SP��h���y�O��'��������[j̝�$�N�/���WIn��HYu�-'u��hn���w����ɦ%k�uO p��R���P��7�k=��p��j�^����tɪ�"�V�F���9��*H3�w6��BqP�nfo>�K]�V����v/�Y���q*I���n�C����3j�1C���s1]�<�E�L�ܰvT�ԯngZ����j����B��y�c��r���7�6ļa�)r�˩	l�=8Rho�6�۱ÐN��k6[�}�p��S��/:��:6��sT�ؽy�d���]������<e��T��#�jlү�휣{9,w>	Iv֤���}DK8
s�B��B��ٹ�7t ���Z�Ƙ�5K�X\!���I�:���O�#F�ME�����Pr�9R�굔l�x't�	�{&�5��۹.��(n���̚j>�`a����D���A�zn���yA�l�36\G�3dX�i�R��U�M���ft�4U-|���˻�ְ��,��i	��f?�gf:���ĺ���g5!�!.,���D���]0��߮q�}{�u��Y�®� w����Alb:�u�d������VL���ORT��(_-�� �P��f]ZX�=���5�+u;J�6��Vb��CB �(yμ[�2˺���������Xq�-������R��w,�N3��pӴ���G��z��]�����ͽ�}���ζ�tv�D}\�<Q̲̙����*d��صY��ʙ\{V�R���3�&��������0V`�"��PH4�oh����E�~ w&ə����B3���l��R�凂[kg1f���5W��� U���hV<b���R�؟;��5`ͨ��y�;E�&͚��N��Կ�^XN���Gk����&�o¡�|��(
N�)r]�#9o����u�%J��WT%v"��sn�4�W6
�Ky�{��WC�8x�͖���[�2a�*���7X�s-���p9[����4w�y����z+�ռ%�qq�Mu���;U�0���Y&��:�w;�y�+�iCE�|�������S2��E�m�k��|:���5fT��������f���į��y�5%s{*>2�^�i�C�'v��/ybq3�zw��<�Վ��Ū��Tw֪N4RچX�v���;}BI���8��SEu��Df��y0�H"��z�ud��7zuJ�0��=M��'L�ő]��uKn���1��O�Q�l-��m�٧3�n���e-slb�]�P^%��i�i�+9�\9�Tu������9-|�K���̧f�)�5�v0 �]5}i�Z��%�4g�w�H�%lיf�E�/u��R����.�>���_H�������+���p���_(�s`��e��j�Ҵ'��"�}x���|��O�b�C��`:���8A��6�X�rP��;
)�|�z*wW;g��{�r�u/+���e�Eǻ����U�U�yy��6pN�R�b��vuąܚ�����{u���1V�	�7h9;�H%EW(��\֜����t����%r�}O���w�C�*ow/k�� �y�+�c����R�}M_.��ŽB�l�+7�z�]q�r;�X���ٛ);�c��0gv��-fpT���;l�8��[]ҁnڱRFd-9��,́%y짽j��A�q�op�</]���o,��']���]&�k%����ua*���)`�H(�8��Ȏ�H�R�d��9ɫh^Q�`R�M��w�/]m��]b�O+����+�s�N���t٦WAB�q�i�>˂7��V���f�}�-s�+�O��ɗ�B��ArS!nՃ_>��J����)�M�J�v��yc�;��3�9��9�I��
�"�ƪtj����=�΂��C��Ù8Cʄ�q��XZxC,���{��#JfӪ�c`��\n\����ww6ڜ��K�ѳL+�{.��p-ݼ���W�\\~p쏖x��o�,�{;��Ï�	�˙z���K\��>��[��	 �^�{�t�n�ѯ�ou�9|�ޯ���u�je�͇%!�E���$5Gݼ�8^����Q��0run-8;c��u:S�l�/�BOP��e�j����6��Ӆ:��q�R�8*u
�uj܊��e��S 9�]k��ޭ���wr��4a�I���/UM4ks�_*Hݫ������g\瘥By�i��V��|�"�1Ў�"���9�����O���k�V�ՎU�5N�Ht �ҶjB��3Q���4+�]��2vJ�� =;t(�t�?vVI���<�aZX嘤)�j5�n��Ύ��g[�{�y�hW�*�:�eބ3(�b�F�Cvr���A�U��&5l�+Jc ���9��j&����`��K��}|$W��Ɯ"Wi��j)l��|S,C�]M�X���M{2�3�^>�>М�D4�Ӻ�,;�W�.<-��1
�E#@�+��u�N�s��J��!��;�s��^�9��Zm]�go�8��c����3v�����7��Ҏ�3�Nn�!��e=�ڪ������@z��}�]*��oT�۹V���Zv���叭���+h���
��[�2sw�F�����f���:y+cz7��c�:���Y��ҏ_�js����y��!�ܷ}``��S������.P;V�j�S3�y}Ov�-��L��=kI�v�����<z�̴p�K, �j�kM��w����I��@d"��YP�Κn�R�(vc<�}:��I:�#b�vd�6E�(����M�T�0��:�Im��ZW�VF�F�guκ���l�|����2��Cy(�,���,�C0��w�}Q�nI.�CQa7}����eN)`�M��V�B�"|t���(0$dt�m�N��c�W��*jQS"�����!vbL7�9+3Ou;���8�]7�3����s�Z�t��3.�hI\��ɯ��>�W'[��1���S���]�z���H�%u
�Yu�:֍�%Ž�9
κ���� }؞�}]mg�ڐT�#�l[̬�ZI!���2�g��-�u�D��'m�ǝ�Z.�q�Asb�hm��ӔVdV�Vl����g��毆��\aͬϺu��ھK�9��a5���1����]�n�}��5U������*"���{�����z�{ﯾ�}��/v?aU��B���[3[�L��5j4�k���Z�5����n�|:O(c��I{΃6d�w��{�}��K/��c��Ʒ���LЗ*L�IݔhEe�#+sT��{c���3D�����9�Эց�O�h7�NW!Ԍ����ck99����`]�۴n�^n�[� i�@�S������
5�\8s.u]ƪ�Zv��#��V�gXQ���� �U��#]�D��K����Sh��jٸj1�2�v��	Y@�nh����э�*�}ø����l�`�Gz�7��M�+�i-�.���8�BwH��5ut�;|��dU���J0.;0�q��_>Mˣ}�1ۘ�uw�u�
}u��Vt��8U��,#�u�v�&y�dd�c
�˅��XS)|�׊�i�Cy���0mvZ
��{NQ�([��'c��}�E�9�VV�J�q�cZ�-㔺���GE�m!Oy���U������RK#�[;Y2�+_�}F��)r�oD�U��c��(sܺ	nԡi�i��ؕ�����j�9�Տ�b��C[�Gi_Yhep�޻����K�̇�徔��&�T%l�����h&�+�)@̊��9@(��M�ƣ0��si��d�+�Uiv
��f=����S0�<�m䏞�T��֋����۽���8���pX�k���\���W��B�hpR�6;¾����t�U!v�^>{)��,v��tک����j�Ki��XL�����g�$��Hw��MP��v�t����!Ŕ�Ě��ʰ
(ne@2���`o@�ʺA���T2�[X���uuC�C:���f7������y�V'�J��ԥ��n�dA�.[w�R���I�gl�U�Y�A�|˭v+�Q﷮���a��#ȁ['v]���K6�]DM��gҘt8��U���h��+x���[l����ߝ��Luv����_m�h�-u�ގ����{���.G��e���+Z�O m��\V�`��أ��&�Z�d�U�WP���lk����f��,�:kF-S��k'A�*��
����V�ޝ�> cFcĩ�|�1�n�z��v�vv��T2RoUJ�C��]�m�7qM�9�|/�Ah���'�Ge��S������p�3,c̼��� �
}C�az�*��!}�lT��p����c0Jevmq��r�ZtGC�j���2ȽU�Ib'xi����~���1�i���ue�Hj��G>�ﺋ���t9���$��Y����sr�Nd�O�+��0�+�ɡX0v5e^Y�<�h�t�^T�՗�r��.\�Gl,�NfW%ǗV.ə��uf����'I��k��n\�E$Vn�/E��9�����b��f I���f��C-j�l�*�|6�Ԋy k�&��J�\�5���1��R������Ch�<�K�Jc
ā1�~��Ϗx�@��<�N�c5hְRw;
���g�*�KFl�6��1H�ʍ�u��:����P�B��3n_�ɋ�k���R��7	�/aq�������{�9�$h���m�����jս�v��s�=Ӌ���xEU��+xsYRgP�	�e[�D�y:j�A���U�q�F�m&&�]g,���N�u.�J���X�u��V<`hzhY����]5�N��Mk����hndn�֘��j��nwY_ �i�]Lh�Y]V�u��w������4�(R�u�ЏCHve�7�mr�}���+�I<Yk�ƗwEr��{�8��e�ʸ�Τ/�{]�.���+����\~{v����i�e?�B�<gg.�}:�+\�to��º> �������׆��]�{�H����V�釹���D'BZ�lm\;$��ڻ��J�:�=[����h8r��k�dwP[������z��TN��,u]���u:dH��M=�W���ν�UffX��W�lWV�&�]ց�[�ώ��۔���X���B�v�V�"=�yiut�u��s*W�	=¹�|iRz^)w��%�eulEJ�@qM�li��ϗ f�9�q�f���n,ͬԯ��,8��.��K���C��NP�&�)El�p/����8���k�7Q�EW$���"��\�����6��tcY˩#<�㘩X�P5�C�_;��}��7��0��Y�8@�8:��O5�ʵ�����<-�K-<G0l��WA%]�B�<�����ܕʐ4S3��\���Qq���|=�E�=Տ��I�n�iWwk����;r!���á�!� �}���[�յ]v&Y�����7Fs�"H4snml��I�nr�)��z/��=�qw�tF:um��1�hPYc,w#��Æb�X(���á�8c�x�c�B>XY���Iժmr�˳-9k�1�ӷz��@2�s����qI\�X4�-:�$(��e�%G�y�__]�uR��Q��յ+��n��s�X�4h*��W�W�c/BX�-���N�]�ͥϖ=�NN�3@Z�e�7i�,��5�wT�Õ��7��Fа��]�9�c�&�(7ǳpf�\�:๗¢X�v@-��<e��/p��9�`,.ؔu��٤+g)1�ή�������pM��=Wf�.��0�d��,H�Et&�/�/�)ejg��SB�nu��7�N�9"bx�H��>k'9�s��U�{��Y��&bW9^�F�����5��
/f�鼳�[--
*;H��u����j��`�W�����C��GZ&���eL�<ӓ96�M]�1��1,{F���U�
��Wϫ��t `���.�=�u-������kH������u39��NV5���J�]�sM/�ٴ���8.^Y�P�_9�5�v�3��Jc�`+��O9�2��w��ڤ/I����b�Z����ta��y��������ϝp2L���;�B��]�mބ�<[Ǧ��E�L�]1X6���"8�^���]v3�N�];ӯ:�+xSL�;v�7�z2��£�s&g]�����J�eY&�� ��Z�ZWG2=��;UBWb�U���FqǕn�o.�\G��Nn��f�G��V�_B>-1b���-���"%mڐN��u���u��a7N4�=fK(:��/� X�)���i�N�Ÿ�E��&]�\�on�n�QK;j�V#�]b��6��4���MԾ�ӢNM� :�f��w�A��Ƿ���nɔ�\�4D�;5���	��́�r�ː�����p�n�n�	�i*�o`0�έw�캖�TA:�X2�j�<�0EajS�s3)�v�nn��]�f��:�H��b7�;M��7��i��ޘ*Vw[ם�It���ds`�/�{�xQ0�}t�e���sǸ��RDfG���83_8��5؅�y�z�ҽ.�������1��g���i]�u,���}f��í��3�J�P�}�k g�V6t�t ��J��7˴���	؊�33�(uṊa�W������O^
�7���>��;F�k�	1�2HGG;���;�ku�vr'/��̙���#McGm�M�v�v�����*�n�Φ����b��PK�T���i�/��%S����
6�w#� \7�������ޛF�`�N�G�
l`��"l͌	�%��T��-dy�vl1��G�Rl�[gw���|��$��ls������(�����ۻn��a�8wMO�"��@@�w7�{}x�%�����[�X
�]�J �)����C��'B�O�Y�Gm;�ت�j5��z��_v�����Cr�p�[Q
�':�<�ε���n�X��2V=�)��UT�K���0�Y��;	C����0P/z�KD(��;yۀǺ�:�x�[�,�A��I��:+w+#7��,ZY�]JAT����8I�ÿ a�V(NN2t[�UI��T�Xp�Wu�0g�L�C&����v�� �wC7/n�E �ڽW��M}M�⯵pѦ���� ��)]KU{�¢Wq�-ͦ�+�ȱV�0@��kF�Um�[��1`�Fv��2喙�qjp\p$�hV�p̛{x�cz����O��i��.;JU��:���S���9�Y���Y��y.�����u�P�_-�f5����-iQm��՝�����a���q��Z�q�F�����;m�z't�.�Q��r�Aw��[ﲞr�7ǺŘ�g��t&��=9���9��đ��H
�v}��s�Ww ��B9�U�c�V��
*x6r ��.:��˳�vb��ѱ`�Aj�O��J�v�=Π�ayM,�5����B����P�fcd�o$d�Or��-���+c�t��-N���U�e��e
�E������9!&v��zf�3F�u��
N�h�u�JY1��u9�[9N�\��T�[_kT5h�5�]�+9z�"�`R����ڱ\�ޫ���u8�\�2���T�5%��ݭ� A��Յ�)��4�W@ʥ��M��rC��8���sb�6�N�w������d��%���d]���h�Ԏ_�Mv�ocS6��Ꝙ_Q��n6F��r�'v�Eml��W_v:G�VX��6KyW�I�"�С�Y��<U<���O����cln��޽�`�̇{)6���M���Q�Tid�T�'�6�乺�Q�����uFt�s+a8m̼��Ձ��;Ճ�*j�
�����8����1�q�[�H:�?�1`ǵ��:�T���[3���Ժ���w����9�_c���^T�WՄG��K)Mk;J٬qŒ�N䀣�W��,p��QױW:�9>ޚ'v��uJ�� �処�tS.*��������4#��,W{����J;=�Ԯ�oz���D`�h��A��9���G�[<�eo��Z����T�+=���gP�y�\��*�Z5glk%�l��b�s3 u��+��NxFZgq&^a��Z��P��qb][�h�}�`Rr/]A�sr��]�*ظ6;��qT�A:���]Y��Y|p:&Jv�I�mSđҩS�@��>Z��L7#J�m��v�;��k�3�q��t�Ig۽�t'<:FΤLqY���6�b>���YO��)��aY�Yԛc���n�KSF
#���є�W L�KK���J)�%H�k{����]�ȮջoF(�VV��E\��wR�<	��u� C.�n���jr�@a���vܚ��M�m˻z�伙�U�7βnT��~Qa�	`Vg.���
z�����s}�n��ŷM>�}���[��$̑U=] �(����_��{�Ӹ>T@EРV���b�w84�n������*�NGzYJ�l�}k0)9v�!�l�:���U�+V%Y����c��f/�vP�Z&�;\���������_m�%�l��O��ut�;��a�mq�[	v�弘�pc�)�nن�a���u��
��.ǜ)i�����l��1�Dn
a��tq���BlCZKn��%��;����Ƣ=/qm����{8�o5A��떀����d��F��4lus��$tv^�R?��U�;���ռ.Y0���j��T�r�2� ��Cl�-`�-=�[̱��=Y�v�	�d����\�%_K�n���[�a&�����s��.�+ܼk{M7��K�ilz[�{UǃU����ZM;/��5�j���9�:��Ѣ�G6_(h���\(e�!��	E�D�����o�a�BmWj�܊�($h���v� �YK �-��qұ��xt��E���a�
��Z����7Ox��zTV���.vtg�-�Lյ3i]Վ�����,��K�9�[��C�bn�o^�ם�Y�c˾���'9[Z��U�Q�.�a���L_9љ�v�	)r*��{w���(� `ڙq���2�`�����5���FISiQL�����&:}����.��x��2l�]���WfV3�7\fΤ�]n$�v# o��ӛ{������l^�Web��]�q�E�\Z�W��6���vx_Ў�{�z�����p�s�;���
wZM�:��`q�{�&�C	]����jO��t9dj^^�"2^�z���k��p�娫2��47�=�O*�6�����|i�Xc��7�]�R�ܮ+lI��ZP3k�M'6e����2�ti�S+��t��_�ELw���7���U����/1ʗ�6�w�K �v_SL����`8S����=N��z-���w	z	�)��M��ۋhiԪ;��K���zMc��`��93�����p��ݎ��q����h��݉��9e�Z3_S���n������K5��VN��@�r��a3x�U��Ԭ�G�	Y���)��;r�<�X�T8*�WW�l�Bvhw"R�u+�+-�F��oi����_F^BRKy�=� �i.�����5��ņ�m�������9u2�l�lR�ˆ_ْ8�ͮ�&�:i���u3a��67�^��X��q�P钬ҽK����]-v�Z�g;H�z�Q��O����Xs������d�$8��t�+�9zy�a����7�^�ٖ�p���\�	�\hw7�U�M�:[��pw7Ork��⼵B��"�O,�]��1/[�d!���8��9W����<ҩm�iTo���4��ӑe+=XV��*S�e�+�A����<˳1�{���oa�.	�ț��1)���m"�X3;'�VJ6.�r\���n�Q�J/�Z注�k���� ���-��JЬ>Îon�B��3,��U��2��92�i��t�S�Xu�?uj�G뮍��7�O�XH�tBE����� �����M�ES��]�О�CN輺��xR2j|�۵1 ��,�z�\|�V��p�Ie{�	.L����ՠ�^�s�H��T_ġ���2���P���(���fH�
��S4�v�(�$b�/�1���������Qt��m�ڣ����������7��Q6���ըV����u��t9�Daq�z�.X5�x�MH��B��B�%8��USww����ھGb�m�2n�M�*|s���b�{�A���-�AX��W�Tb��2^�W�.��a��g&V)�^��i%7Y����9FU�|�go"�u#���F��feK����Q-�ڜ7��,<5s��q6�:�q�Ԙ��P�8��aCq
s(#:�9�լ�˱�-B�����4:X�_3R�#mݗ���.�gmK\��O�Ւ�{��5|�Lǣz5�2S�U���`��G�����hZ�"T�>��l��or���IP�iX7�����]{#]Ck�yE8[����l
�*���y�˷XC&-!ʇ�c�wc ��vp��[�	��@�\�QR�s���v6���nQ��v��'.�K�]���;YE�������M���+���OYO��Am�wtx��'7es@i��}��-t,V�pKY7P�j#�����3�M���uv�`u;�em�2m�����Q�=/NIQBZ]�6�5y��6�L���:];m����iwMM�ٓg��byV���i^�Cas}]�3s���ͧ�'9y�G|�Μ0�wv[8`�܋�����EͶF�MUF�nc@�'��
*�4�J
�d��!䜢
��4Ѣ��m��R�8Mͤ+F*5Hcm�b��r��71�1m�Q<�F�C��к5� ���塦��&��V�"�m�cRR����)t�'�U��\�j��r)9k@[:�5�����. 9�r�h
�8`�8�9�E5�h�lK��X�F*ūF4m����@m�V�0��<��G 4��T��	����L�����t��b�9���rf"h����R���u˛(*9��M%h����4-��[lG9�C��Ǝ\�AKZm�DE�ri14RG2��8��v�RkEv��}��)b)o`�9����i�*՝�4*+��E;N��1��t���v�N��k����o9r��T��i�᜝9+{f˪��mL/2�4�,�1,B��w�.�ᔈw�b�u�y������,nk���O�.�i{h��5�6��w�UL���M��P�=����]�6
���?F�m��v Syw�2�y�N�s /t~EM����g�?3��԰��������Cy���m�p(^@��T<i���x;�[ ��&n!@z"��s����j�����g����u-��W�`�〯[�1s��1Y��O�^]�z��,��qJ�������hO���&*\2sC�+7�b������w*#������_��m����>I�����	`I`Y��.�,�q�2� /��~ R����<T���Mؼt�N��wKm�9��w`:���8|�Yվ��uV����ʳ�4?�u�`lP\�pP���0sW��l��U�h�L�Sq�F��~U�־Y�x�v��� !�"�;5v��V�3����a�6*ƌpԹZ��خ�^�=Ur��C�}��iu�f� uSϰ��M���Ӵ�҆��*��Hl��3��du�z;��'$a�xp��t�*P�u��֙ӥ�u��ڲ�^dD�|�y�U��Xw: �m䒻�p�cxl�1	�]e��>��Z�:���B�Vb�.�8��� 1�n��n>yA��wgP�f�;��];{#%�&���*�Ԧ�[g|1��\m��1���t+�T�gP��&����*��,��ƥk���ߣ�Wvp{��p��-F���Ƚ�fp�o!�F��R�˺k�Eӻ6|���_5^'m٬��ܪ��A�÷~�X85�w��� ,g���w�C�m*5����4H@̴��+g�PUgZ~�����v,�ܱ���^eB�����w]z�aG���������vb��ј@"'!����0aO�0�-���U`�cb��8��e&�u��/��~���0���#3;_Cj�պt@g@��97Ʊ-|_G%YUJ�W����&��Zٷ����D��'O�{(z0o�� J�h��S����b��~>�7X�r��a�!��+M ��L��L�Q6�o 7@/�݄�{���an�?t�o98c�����e$+�W ߱��]~��߆���5�}��6+�]�����
f{�}��߳ӯE����&3�y��6�ƒʰ���)X� �/��^;k�����\\ek�Q��D��*�-W�,������Y~���E������=;��R2ҵ{(/��v�@?�<,bM[d|�c�<����\��IK��簦벳��%�>Y�6�U��ü�l��{s�mG}43����/�K�F97�����/���q����V�M.p���\�@��n���Z+�*�^*���V�JW�e�,m�����3y]��:��.�{�Ô}f�w�#,��+'�"?�9�KK<�Q"�a���W�5g���sfr4!�<��$�iZɛ��x�y�����i�PWq>��l���}G����6�)<&�6.�9��t������ʓH�L�ڏZ~�����)��'7 YGa�ڎ�(�%ݎ�	�d��>���*�	��pw���>�WU�w���\����$�J�
P�b$�����|j�Ίt6��p	qoV�
�F�b1�~�Ͻ���
L?j̲�xf7�	wE\<q>��ڟ��j-_X�j��S���]ܯb����<�_��%�j�P>ХL{C�&��S�3�:U�q �y^��ts����
R��L�[�Z
ĵ��$�i*�7i��+hO�>;�����Y�^�`��6��%�����d�߻8���(���ǃҒǪ�^:�{ʫ��JN�'�@��.�D�f٪�E��3�' ��+^�P�����[���]�F�䶗���R*)��՘
ˑ��]u{����
���7;^ai��M�V�7�WuF[�n7.=-y]fʬ�ydb�������0�g
e�;�K��`1�����oiZN��9[����Y���̰�[�aɈ�5���Ԗ~s;	��;����k^�zV�"�+�ۻc_���>��7VxW������������pҩ�y�:ۄ���į`���ܸO�>:AC=k̕����V(٤�m�)U���گ�Gc�7�%xL��5T��ڹ�}�7�g��qTc�n ۃ�ռX8~)	�٣s�&��^�b�}�V��Cʟ��� M�k�F�?��pJ��HՉ����<�cx+ؼ��h�G؎����uwnm���[����*�~T2�q���uk~�jUq,�m:���42`����0��g׸�� }�[�|/-S�����\ �,xE}���VO�"5�
2Ϧ��D�+}�{��9	�PU��7F;�Aį��@�߱!��Ɍ���|߬��*��ɞ��~[嗾�&�����h��>R��Nʯ9�N��Y#x��xo��\)�ra%MY`�?%jO\�����Z��=|8Mv2��ȭ�^���'�v�X�ꮡ{�}B���^���Hț�7U�M�ά��7�)c<�A�N��љ&}Ӭ��~3�=�]Э������I�_�j_>e�f�aӽ�WX�Sv���R�o;����f�U�{��� Ҕ�D�L6�v.�T��`��/6���t� ����fg%�8��ϲ�5{RF�7�;x.7L9Z1�)r�O�l���`S��@;r�B�%�@��X�D[/Ϟv<����z��q*S�[�<�_����%���E�#�Uy��ۺx���v�Q�hfu6�k$�✳��+@���$O~���k>o��WJ�+��a�/�I���[�3Ph��{�z��pQɹ�Ei��xy�ȇ	U�>��9�h���Ǿ��g���6�ӓZ2�Y g�nJU�_e� W��p����́/H_lx̵+=
�r���n��Ww}с���(�\5׊�|r����J��5c� (�t|�'��5�kV{ΒιO@���C�7���0)�d�^E]V�|~d��mz���S
�����ګ�e��/7'&�;;+�O�DK~Nb�[T�ó3��$N�D��)+F,�����Yx���z{�+٫U�S�?{�������u�+���0� v��7R6�.��K~�G�)�7P���8)�����-O�=o�N�Dyױ�h�'�ȷ���ېu�)���z�bٙ
"ƪ���f^ �"8�MA��fs
'B{S��j�/�d]~��RV��F�<��	���;M8���	"�ٍ�c}��l$2� [���O��n�}Xv�X�-Pq�}�j]n�en�h�c��Ƀ��/!gaX~����^��\ ���o�Fd���0u��Sb��#/ژY�fa�W�A�ʼ�����^x0��$HU���Vz�����¯)�eR2�Ϧ��Ӣ�L����1��ZeN����>�c#�<�X;��}�t�ZX~��ʫ5:y�K���r�����|��^��.z��ĻF=7�4|��i[HQ��禞��b'�����(�a�SB��ce\x��G�M�6���l�]�����韽�����:�{Sꄨ��K�y,<� ѭ�R�q�P��2���_O�z=���Sx��O�f��J����QǊ�F��?6/�Kˈۺ�����	Wh.�/�U������Z<6c6�o��^c:�����>�2��3��^�U�+i
��x��ț`�z�����c�z�ЯQbsK/ܺ���Xz��0���D�#,9`1�ٖ���m��g��/��d��2N�H��a����#�:�����3l�������<j����fU���ٗb)/OQWԧ*M�S�觯mp��Ձ���VI"�Cz��&v���{�>����/N��a��]4ڹw��m�p��l��Ķ�^��Jb�z͇̈́��̬�':r�0��/�� ns�ɹ��t�����l�}GnK[}�bcp}�g0��̭aן�j��P����P���`:���.��lT�^��ghy��ۅ$�R���oO|�V�Z��<3���L��:�ư�N1��;�
5����g�$�;���m�'�(ػ5ҭW��倦����ǃ�R<C�U�}�Y�mNH�7I0���
�E�d�n����Ԕ$�N��טU��񤲕����ʼ�s$��Y�M����:�j7!L��JJ3�-�*�׺��>@m�\�s���ō���s��<�4I��Q�u8�P�Wy����D���p{#����k�"2�W?S��ѱNs
�}$�un9��زn��^~���,�W�-�ߘ���\N����ԼE<���~��L\�C~.݃�/�6��\s}x]�ܚ!tT����w�jB����{W}���M4�ބA���9���pCI����{�K��������zK���P�k�D�o�m��
�>y�Wh��[�x�fۙ��:�>c�Y7�્c�y��R�U���?z���2�.�c^+9֊çrbu��s�yV+9�c��L�ܙͰ�����
}����z�9ص��O�����fOa�1��Y�u RV�C����f}�ΙČ�S��M;޾j��_(r��p ��ԙ�\��͗��5V�*�x#�u��(b�0���!U��6]�dͽ���2����m�.hj^0]�s@9I[�}Z�����%Wz\�%lO�_āܼOƲ�����Ӈ��iewv}��{�ܾK8&�U#�~q��.a�V�����s�3�:���ā�r}^��g9خ�}�բ��k5���*K�y��ݨc��SV+NCǧ��s|�5�8:��,3Z���w���̟A(�{f�C���	s�Lh�L#�D#���Z4țxk��a��W4ގg�g{�;��8z*Z+%��:B�/���>xm��3���vd�!����=c#��N���f��ox:����$�gf/MG�U"�]�����������7W=����~;/=�٠c��͍F ��E:揎�S�Y�7�+��ߑxj�j��;�4�*��ļ͕�s���Ý-�<*vfaKd�~��so�WP��2�U�dQ��j�.�(s��O1���p�y��6	!>��ۇ�1��C�/�{ON��7M�PW�`���O�hy`k;����G3;�b���@���3T�O ��n�a�򡸻<�}n�JYd�Oݗm��a5�����s5v�:�b�V顓��*�^��}u4�/���v3>8֭|���8v{���G):�m���+�+vҡ+C��m.��칕�+�:�����X��]���4�yb�`�M�ղ��ܥ3�]�w��Ws���V�*��Yj��'ecC�m)�1�ܹ�.�Ok'ʱ�*e�$v��y���J�}��5��½�Ѩ+_�����B�W�*���u�>�8ӻ~����F�������:�����h����m�^�o�F���}S�:VH�.�^�j\*R��e[�%V����߷o�ݹ5�~��k�;Ћ�*hǑ�7��`?s����+��'�
�	ay^�d�~�)]������ن�U�xn�/
u��x;���@R�k�N��r��gP�ۻ�!��]��)N�TE��؊��5^�Z_��#���-�
���Շ�]�{���&�ٙ��xu�Wꍱqy�g?��/q������|���x����yƻh_?y�:�51��e{*���Ŝ����i������b�<"��LxX9��1G�Z:;��>��#�U�]��_�T������}���m�7�5�w���\�̱da6��^���\�ա�;0+���{� u:z "_p����d`g����c�U�{�4��m�'��ᤥ�wWފ�*��9�b�Ԙ��/��:�[�;��4֞��ej�xl��&�!e���t�XS9o�y�*�6-X��\�C����B0��_A�ye���n���:XW���We��u��˶�j3��t�1����Q�L
���wZϰRw��|��d��*fc?P�Z�αpS���"�`]�Y`��$ϐ˧���k=%�����^��ݜ�*P'Ӳ�
��:"X�	�T-�r�^T�NЁ"Lk����Ip�2�c�:�~�q�ᖐ�jǅ<倧o�UX�+È5W]x������{��b�:�'o����}� �O�G�厴eU�x|.�
˪�^p���=���tG�G��^7W�*����^͚ك��U���@��c���^�q�2� /����g<���
�=)�3/ۋzu�i^�}���1�Y�C���v����[K5���^T�D�z��~o�)�jeN4�����^�w��n��h�yX�v��H���sU�1%��=R���%�>W�7,|�=��-\5'C�v�,0澕Zc'��:;+��|e.�b���]{�)���ܞ�v��筋+�K��{�q���w�{#�y����Tº�M��쳚r����W%������EO��s]@����=ƶ=�V���r���> X����<K�i.�%��r1G�N�x�Gc��k��*l[|��,�9G�Z�ƺ�{J�S�n��aP�N�s��}S���Ďr�֘�YyW����I�m�����SY@�`Yw�Y��?3+� Ց'L��1�����GZ����,l=�=;���ˢu9J[��<4�(��2���� ��,,r2�]�1AJGy���v�t�α�����bp��*L��!�#�&v�ս�s�8��|���ټ�C]f�K\�\u.)έ��/��:�⭥Maٻ3���Ь鏲��0FM�$cnʾy�D���s�v�uRNRP�빽R�u�W��%p�S��Xmm'����s���c'��,т�$�Jd�fn��+��(S.�(�����6�
�+�[+8��L���o��M��ٖ�Pb�n`��Uop=�2�@��M�Nu(5)�ևQ{�����o�vO3��.������Qgr]��g8+�`����4xh\�0p����L�0��̈́i�j�ec�+�̧ٷ��(&�˹�#��
�ofg16���l��O��5��`4�s'Nw]��)��,rjTt�ۼ��N7��* )�̷Y!v�6�ջ(^k�^i[Fw����U�ۜ�q,���2��QH*��W>�1����q��|���;�gr���O��Շ4B^c]��k;�h-�@�"F#s��|%:��}$}}d�y׶�3�p����)���������m���Cc���WW�}7TEr��R�eݷ�P�uӼW\�Ʃ�w�;L3[t�&���bn�=y7#="��b���m�)0w��׼/�����
�"1G��}���Rh:E�9�.�	��%�v{���=���	�/�Ө�݈e�'E��s�VϦ���3{���L�4@m!��e�Ɇ��Yϲ	�y��ԛK]]	uy]��.�����kO�Q�yYt��)�&�5�U��WV�:�o��&q��17kz�[ُ�:o���̳�7��e��I\�iwYGs���:�拘(����)	A���T�\)/-��z�H�`)V�S�a��¬�bq��)��t+r jc黣E����Uw7x�\�b�u��a��L�����F
�\�w�����ۛ������IV0)i��׮蛂^�Y܏U�ވ 7�O���}ZA:��72Q��$�F�r#%�k�/�!���ɑ[�̆$�.'�	�_:gl�ګ�9M���c�6
�h��8Joz�G{]/��Ju�:�Pr��1��Yy}Փ#1ӷ����sgf9�]l�L�\x)�ՙã�t{2��w�!j��c�}�$ov����w*v���9`�i�&����[Ckcg��tf��#���֗*=�����V�ن�5�v,Ҍ�a렳�P��hq�:�Q绢L�����-��.��J��j1�2�Rˇ��:��sS���]��enȲ���} �m:�f��y���C��j��v)�����Fۍ���N�=K�
K���̬uϪ��OVt�����\Nwj��H�^N�ϖN5�z]�w2�x P�| �4�@ry�W!�p�TPփCF��k!ADAK$H�+4Q�sJy���nnM��r��t�KBPSUE4U��X�Z��<�F�Th5N'DN��QS�'Fֵ;%�lW&����ri��R�v4UX�KM;FA�Uh6#%<��1QQQE�Sc6J)i(�
��6�m�&"�4����#CE�#0P�t�-��퍬�j���9kX�i
g`�#��\ܹ:M&ؠ�ڍ:б148����'��i+m���4�j��F����6�����<���J4ht�m�M��Z9&�j�E1��e�k���nsK�u�4U�i���9����' 4&$�j֍:��R�O7X������D�(o"����3FY���t��q���w҇v�Ӳ`��ֹ�r�m�Z��y��՝3G�w_U�޿��s��說c�J����y<��`����������q�?Z��<��w�A��>A�A�&���8@{̟�|~��C�<���a����yD_�����~�>�9{�|���Έ��1A�9P�{�4?`��]�\�C��]?S�{�=�|�������>\�ϼ�T�I�~����8�Wr��s�?G����n��OP}�������ff>��N�	s��<�����!�	w�׬u?א�^ӛ���h��<��h�캯�߿:�z�I�󮓗�d9�|�Ph=�^Ho��]4�AA�o����-R��������>�>����s��7Ԥ׻{�B�_G��y'wP��#����?.O��q�4w	T���9�C�~�^`=�A�Ԝ����u.�>^߽pcK�޸�S�t:z9�4y��{�ܽB�:`�L�Z�<�/�}r��5�����|�y��c��^�T���������e�C��O[BS��׹{���+l�C�{<��_�^�`+A�|���;�Ѥ;?���s�� �0&������U_��	����?@�=w8u ?F�A�>�~��S��|���:�Kȡ�4a����9�k콿���A�;���Ork��%?=����r��9�u!^�1]p~�7���~rr���<z�}@._����9@wC�<�������X�;����6��|��������)��^A�~��u�4r����i=�ts�p`�����*KD�50�0qVP�gT�5�+7�A��]K����t��wНT�?|����;�	����������P�����t|���\��~�~�������? ������{ �u�i���(��#�)� ��������f����{��@~�^g���:z����u�ύ��t�'��w���?e�|�?c��_�*_��{��:y/�����C�?C����O���	O�ލ���;1S�@Qm}��+\q��Ջ�������]{�B!��<�Hk�
�|��A��/[Z{�`��|��{��M� ��k�7�8���������u�?Kϧ^�A��h�����i�2�\����u��O�]8eC�[.���V��}�+�ʉ�����ݍ���\�����4m��W�kY�ԙ��Ouwk��U����,��	�w_k�m<N��lVodB�v�qr��W1��� ��R�x��AȻ�fp�z�kh�)�������1Y���]�7�;�k��_�){D`�쳙���U!T�W�c����BW��^F��ʟ�켄�d��Gp��>�n�'�c��_��Hs�����=����R�?���#�Hw�=�^ɠ���y���\��ug�X��o68ч�|n����ݞ|�i~��|��.���r���nBy������_�xy"s�?��М�_�y.�e~C��pݏ9{�B>��>��}@~��+�h;}��K�r|�����? >ƗO<���<��4|~��z��t���A�>A���O���!��G?�� ���#�+��1^}�
�7�y���{[����w�0tC��L@���-�F1@����W��/^c�J^�ࣩz��C�|�΃�H���>�j������� 4h>����� ��wQ�>A��}GM|�RU�Q�^X�e���~�����x�'��t���������'���>@y�w���v'p�����Η�y�9��:O/.�?�z���.��*��C���~�����BV����70��銘��q��s�>���w�?��]u�{��=A�=G�a�BP{�|�����9/Ϲ��
}���>��u�4{��y/pF����|N�@h|���Ri5�_f��~����}�~��럾3�^o�1��ݟg��_�B�M}D}U�� ��U.5�����O�?������� �u��p���-�4?�h��-/��?�}�����i{>y�Os��<��7ߺ��~��s	��ފ��z�ν�R�{��� �����A���������P��Z���?��r-�k�:�����CO���u~���u	_~�������_p��.�~W�1�L��G���q�{��x���?GPrF�_;���>A�9�\h���}��Y�����s�?Iʞ���̞GP{�G��l�@y�h��h}�_O�}����$OL|g�?B�����4!���8ѝ׻�������B��ѡ���~uBP�ߝq?���%i��&���?G%��w�_����{�~���%���z���������h+����������U|�UxQ7ޞ������n������4J�z�0K"gor)=���e���S3K�C#�O�ɢ�~�jFs�p�u*��;�k���O�Z�]�w���n���R��,��f��+��+��Y��s�[}K�x}D�UDW߾��u&�^�e�<��:�A��/�8�S��{�8��T�O;�u<�`��C��9�܆�ײ~���}�?G��	O��>]C�u����T�cC�;��)��4����v�J�z>����LA����o�|��O�ry?/�yټ�Ӫ}�t{�C����>�>����=O��u=I�{ù9>�#�\��B��5�}��>_d4�9��-�,�"�'�E&��s��_�c�->K�e��^��c�<���������x���{�������/uL4��P����>���7��1=����V�ve_��)��\�R����B����>�ʏ>�,C��Y�>���AԶS�ݎ@6��L�y�}9�>�����h{5p>�ǅ?����9�<�Z��m5y�~���A�&z���R�]��O�A�����wD��%~2����x��s�o�_.�m�ykl���:�F_|==��{������^�(�A�eyϩ};����z�*��7�7[�i���z^�uul�!^�<�u^�k-���)z�`�����c��O��V���t���i�m�n ��3�E߲�,T�T/s�;�
��Ӆ�GNJ�0)���e�X]��,0�0�_xo�N�p�?����46�T�Z�tE��z2<>�-���G�:��n��Y������<��咬�ԋ��Ps�;�H�t�F_fpꂍ�P2�x�W<���f��j�	r5�����j���$c����V�>��a��v�]�����γ�|��G��~��(8㙣�(\��T�؝��uNص�H���K��U����ݼ�����>�b�3����;x��c�pux������DI��nmz�yˀ��4[����Q��Y뺟M�g&�������X��xW��{�iv���$:��hhw��d�gMge�!�U�#ں� 7گ%*�/�Ր+�L���d�l��7�y���mf�2�4���0]V� 5�=�J���_xn�xݴzRm~�]��[<�=n�D���v�)��]z�>�|����
dU�d����;��Y6\��2������_'
|	��OTB���h�b+qE�J�ɸj�L�D���l-wU���1N�����2�@�]7�v2��������Ɉ+,�6j}Ge���+[�S�J��l�C�\9�f V]��� �S��[�|=���F6��NS������/����n���ym,A=���q�2� /��������L�ӻ�������3��b�Oa���1�w!�V�����K5����FA��b���*�oӮ�����B<6ߏc�PZU���ǥG�V6R�ox"\��R�p^3��2�M�5~9�	������$�%�+�Z;�Y粥s�t;8�̰���OC�w!K��*� �X	M���^���Ԣ^̙����H*���*V���N�{U���?�K���d��IW���7ی��n48q6 ;+�h4y���J��9	��������D��E�z��J๩:��2sR�Le�uƿ��ԫ�
�-ͷ����SՍ�O=�'֦�Mh�����>X�ex/�~�#��}tҺ��(�X�!
�UgS�eZ�@;���'���k;�i~�gM�_g�j�[i��=-|�|�����:�����p����V~�>'�z��,j�������>�X8*
+�#z�����ե��p����{%����~2��#Ɵ�j��O�3m~iZ �c�#�sقSdy*����j���%�b���5�����1_<�@?�$/s<%b�\2Z��B���g��;���g:_z��l0<��M�M����b�06{�u<�Q�i�uޥ�4�A߻�	�Z�S����^X��Fx�?9�<���îy�ѯ�XKr�p��}�+0���ؿ5$�P��@�h�M��~��ҭA��,x:��oS'��<��y5�3|���2XB�ԬCGTB5���w-�3"��+'+q�|9��m{(�Fe�%������F�W!ڧ>S��������oV^��k���A<u�Ϋ��b��T��t�c��H�eS�تsC��LGoWm��
N�b�n
�8�<�Ϙ��47@v�R�Gܶۓ�l^X!��yH5�;�r��#l��]��֦�]�K�5֐�}]}_?Xh']�N��粽��fO�]��x�pB��v���{���覰�񃉬m),(b���\�V(�D�3��f��^/�ݳo�kޅ�z
g��s5㺣��Xv�����r^û��Sグ*�s8p_ԽJ�]���:y�x����/=�+1�(�O�lV�yoόIҵ�7R��+�C�P�q�L`vjG�{��I�q��|�݃����Lɜa>�ݩ
�Y�����etu��9J59�V֟->D�26�F�N����+4��,S�aBɮQ.��q�HK��g��t�K�{��"���k�>oG��c�d��|��U�)h�A?z�٤rp?,κ��TI���{���&^(��6hyӝ�*rW�n��ND
#C�e�R��Ɲ-_k9�P��~�K|�����'�����;=�~ߧ�@c�h^894�թc	[�̤/�&u\�}�\�|���r��^ox/�ɎM�ǎ�88b����}�m{ڊM���a��{�_v%��wJ�S��k=�ӷ��u�����Sh�����[lh=v���é�u�����͂�p�i`����S��[�k��L,+Ҿ��G�<�%��&��u�u���n�+>���1����m���I���C��̇&�nykM��)�+]6�{����j�w��ŃҒǪ�E�6وDٖc5*�x	ٵ���T�\H��>򥢲U��P��A���mU^u���\C kt6�z]�Rr�������F6gn%��V1Q5]��Qj����?mK�Q�¼�p�)�������:�w���|1|<)ڀޟl{ƃ _���E:揎�P�Z�o2W&��K��c+���T&�ǻ+�6�7����30�\�Vju��e��Sj�6��������z9�.9�=]mᕇG�O�5G�^u�U�_;|��Y0W�&=^�i����S�Y2�v��c���	�w<2���P;2��g��+��|��_ڻ<�z�y.Q�V�s��gnx^;�6IF����3�~`Vq���|.��0��}1�앯��.�x�`�61.�{�{���S���9�Ơ����V6Uy�0�� �W�/�
�X��i׽���X3��8$�8���]Y�[�U�fD����=j�Q�խ���!6ٹNf�[G� �h�Si��๛�%�j��s椽��or�N���']\�u��v��h�2:l�����omnl��&�lwl*��R��ݦ����L��do�>����}'��"�m��7��O1�\��{^|�����JF���}K��r��F��c���ͪ��'Z��M��s��yɇ[�k-���)z�`��`V�c��v-�1`i·Ԟ��%�u�x��N���M���}�ag+����;�\B{�.��/m>;g0)��l�Y^�{��͔��|����������fz���ʗ銈��ہ-��������%�P�Nv�z�V�����jte�Ub�
XA{�}����ͱr�>�b�3��qݪO~��W�w<���u�M�.v�t�@CU��U{���J�K�eb����F0���@����λ�5���N���aļ��T�S˸3������R̻�������W5� +֐�>�u�\�������Yu:¿W�l�r�ꎏ 5�� .w��_p��x��]��*���<�T�ۧ`���L��&�U�kʯ=2����H�[�M�	�2�}�`�j��T'vT���~�(�p>�l�Ɩ100:c���l��4D����)mS��Kʙ�B�3��0��}肹�G\4r�[g��KFż6�=�{0+-3��_G2AW�ҧ��ܘ���XH��
�>9PU������ÛPE�ɽ�#]wYЌ���2�[���T>mp7GT�e���oS�9 ��fapvmx���s4!w\+���}G�m�o��Bh�?W�/q�IcїEY�ҭX�X
��fS�r�����S�HD���ndF=k���~��Ь<�{�v*{��d��K��^����Ņe��𣇀�O���{��C�:�*�cŨ��e����J����"�nݏt���0�U��T�:�����'�	@��Y��fa�2�ƫ(<�=��������}��	�����>b>��f]Q?q���_s9\G��i��.r��d�0�W�ÜB�2�f����ގGb�bv5w������={�+��̺R���xoU��K���YD���;>��Z�%����������[ˇ�~^���'n`a53H��7�M���˸��*�R�����l�E���Γ�r�X5���eu��z����m��X���5�*U��R���Λ����ݭR�G�^�ύ�x��a!3�o!�@�U�<?4/�Kͪ3�w���\U���;s�>��U��sk�!I�x\&v\�7>�)-�*�#Ɲ���R�)g��yu�� �<Oo��m�M�Ww<�kf^����ۗ��U)�[%O�^e'Q�[�՚����S%=�����x�u�}����ʛDqˋ�cw_S� �u��x�F8�۰�����R!d�����Y� ��DiS�k�v�o#c�ѣ��ꏋ�kX�1�+��G�&+2�Y0د�VO����ƃ�^DJ�Cǃ��Ҕ�!9#v[u�;/n}�Ƨ�2�iU�ݍ�T�~��]�xvY�۹�FC�T@j��m�����:���b N�v1A�i��`�Og�j�r6�t�F/�>�*��ܨG�2q[��P��s� ?��k@&�K�IX=fG<%֦O#ʧ����w����d���S"�_g��/��%��|��JI��:.�t��{�倧��J�ڠ��ÉF�R�)�p�&���
��
�g��꽰��2ud��^�,̟^a�u��S5X)�j��f���_Θ|R� ����G�4�׺��>@m��<h\�	W�fSk� O{�,��Tm�_���2��^�Xz����:�~½�@�X�u�3ł��Ê;\m��vٝ9ʾ=��Ds�¥U���g��Ox^g:��{9N����,�o}�Ϥ�5��ܷ<W^��F�A�^�`��B-�:���2�/i�ԅc�^ojன�X=�5S7]��]JnKO�����&;EE��Cl�I.��7�w^���1B�w�fwWV7T����t�u���읕m�Yzq��|p������\��y��7"��)�L�tVT��ڌN��ѵ6
qV6X�8̆,��*�B�Y
��;�s�Cw[�:��V�Ju�y����f�@s��ܶ1�F;��5e�f�>��2�O0T���B%��.�+K�շ1⫼�Y's������� ��x4�r_%V����OFv;�̱�h���E��]+������BC����r��W>���ӓ����9���4;7�\3��
���-��mv�"v@���'{�7���CuJ6H���zKγzRƵ�k*����Z��]���hH�1u�Tގ�r7�;ī$��F�s^^|�4����]ʃ;H�5�t
VWf
�^Tǔ�P�6�жA��U>g+�u�ïihi.s2�9Ν��nLۡ;�I�9q"s&\!�N<��7cH�(�zk���K�f���j�p��7��f��f3���´�+)UF76$x3�\!u�9����d녪���7e[R���su�w�P��q�)�U�6�e�m�<n�k�L͙#ݨ٥ˤ����K��+������b>�v\ۻ�e.W��@j�������4+U_^<u��N��D4NN����[*�k����I�7E��,u_K�1ݝ۲�Yz���I7�O�Ȧv����.��ӥ$�`�"��Ηۨ�Q�N̜��=� �@���Wkt��=�
��N�����K�[���f�`�"yJ�b6��:uʧ����Knd�n���k.��_]��DU����#���!�2e�蒂Һ��y��2���/�w�!7��r��>�%�h�*�74hc�hЦ4k|�sc�CB��',voi�/K*Ŗ�����ɼA֡���E�Q��b���pj'���Ӥ^;}�kZw�q��Gy�Ay�TG�ڨ�7c'J������)V̕�oE E<����+���/B�,.
,B#&�o)�"4G�s}n��rIrL��^n�+�c.m+���[ՠD��˛�>�,LT.���[VTYdhm�[9|�X{@Ԃ���S�4�_E�D�C�ؕ�{�Y/�4s���n��Vy':_t��I:�R������-3h�m� �t6�V�h���( �<� *J�hM�Ǵ'Qʕ���4�7�.�T�vo#ub�r
�߁�,�[�>�I���Z��;�i�/xr*�S�鲳Tч�>�S#[K��a�\K�3K^_evK�+��,�ޠ�qZ�86��栭)�*�|e�),Gk""%���U�4�O%-��v;�J�ypV햜�"���m�\�A��2�
�[��b���c�
y�b2$ⵃYw�L�lt<k�A���o7A�xMk���6�nL��Yk��z���ԝ�G"�ҕk�������Iշq�y�:�	��/bA�ʹF��u|.�]]Ձw��}�/1�.\��g��SAI8Ű�cVͲh61I���6[e*���X�浥�:M�֝�qbUNٶ
��@[h(�TC��H蠣N-]sp�l�rs�Er�S�F�lV-TDhŤ�sj��i�Ps�����s����b(��ca�:i1SDT�cl6ۜᵹ͂�7[c��TPEO!�ιb
֠�����5�˗5�F��᫒k��m�͹�m��s��#����[mgI��)�sl�b4ӣUV��m�6��4���*��-��ђ�#mQ6�d��1V�j(�q�`�U���(Ѵf#lV��l�VcQTR[m�$���&b�5��ꬶ&H#�u݅�K3M�:d��l'�;k�7B���mXM�q�|:�(Ґ踻	ۻp�I:���1J�Ȭџ�}_}�׫g�{�Pe,��xVJ��?Oe*��N<�����P��)�%N��\� Q4�6=F3>�����\&���
]|]ߥLMΘ�Bu/��U׋EJ
��p	qo4��4X��"���m����j,����۞�/���>^�Y��D��� �K@�S��7SV!���~z-׻�e�@�̫�3�Y]��H��T���_1.��j�-By��V莕VP�;�˞_BOy屙����D�8VL\�!�l7�c7]t�c��\khu9�F�ݣ抧׵�Iz5I�����*U��x����sb�n�//(KP<t�F�L#c@l�n�{,%�:tb~WUw�۴K��s�ϼ�xVZ@AuY���9uc�m
�ׯnz!�Ki{��:.�d���$*Xh��3�n���R�.&��=Q&�{2��8�FV��ڠ�d�\�^�o����y��֝� 7�{�f����0�	ck�O��U{����ӏ1*����P�==��,�*]�� ڢ�>�C.fa�n��ȕ�so�
�W˨p~SU/��ԦpMI����@nڠsj����=��� ���~[�g%R�L�T_
ΝZ����X�x��(BW�����C�c�ugyP�yR�z�"��c7Nw�����������H�a��7�V�l1��Nғz�D�V��7�u�y1��w�ا0���?��>����Z��F2k�u����+�������;�5�L��9`
c[ʹ���V�+зst����V��Dd��q,dX�\���O��̾C<�i�7T����5��["��R�4+�c^�㫫Q�X�{�d��Sr����a�L:�@_Lh{%k��W��۷w���x�U��ӛ��ڮr�q+l��=�A[��� ��_�� +���zw%��Z��ۧ�Ւh�S��J�?���]{�}�W�ѷ^�")�;�W���Q�F�lL,�}R��7�K���ISF�X�#
;.\��e=;1�1 ���x����j���afv3�޶f]�DtX��҂�z�%z��C�`����iۜ�NPCe�r��/B~:�!m�>˲@�Ō�~�d��@�V�
v�oUn��մ�dx}��[>��K֢��$��4()�P>e���BtS�!�Ka�s���E�;>�s�װ������Hּ�ߟ�l^�/��ʨL�{���mY��ڥ�r��1�|��A]��Y��U�����J����Q��zsqnV�K�0J'���^����Lp��׵�j��&���iTJۢ��ɍr�j�u��d�J7�����G(�4�]:z���l󌛋c� ���7/��Lj�#3�Q��]�s�;�(QWG
�p��Ɲ��g}{�U_}�Sw��,<Wx�OT�D�HۅP�CŔ��W��Cܥ[l�j�Z��۱|6�Qz���A(^�f��'�����ȹ��Z,"�.fv�ˊ�n��-��Ϋ}~���s=~s�7�G3Uos65l_���qά���W0���ʞ�7Y=WlZo�=���}��z����7�4|2�x�������7�S3��gٕz��n0�K�T�1	�ﬗ�n�S�G��c��4J���~��\<����`�zr�;��=Qo���]��ߏy�r��6riE#�H�\;~�kaý>M�����Y��>�_�ˏ�����9���:"�ۼ{䏯ԁ�N�J/U:����X�c����{
��k<�7}���8(��o�r�����b����1A�l�Rz��~yv�����ףD��y*TH�-�~[0�@����|�ٳ��ֽ��?���v��k��n�I�}���ݻ�A��k�����F�G�w.ۘ�p�Uyb����kV�eҕ��\���IA�����}wac@.րo����k�Z � 4�M�e1�:��VaY4/H=��M2Η�%u=���rS �0�������8Vl�U�}��~ٜ<�^�_��d�l���k+}���Dt��Y�=��}͘_�����+�.�y�[��y�:�Wz�շ>�)S�]:�|�wo�U�5��YN�➨pB�/kk���2ߴd��	9ع�Jm�D]k.p�ze��~Z�}��ձ7�΄�ﮧeY�������]�������!R9兽y���2�)k��y[�t�#7��|�5*dedi��Y�R�y�㐲�*�%��I(�ޙ���5��d6A�Wq�fL���<�Z{9[��z����Zy=�ע����&�~��o����u�S�f�熻��}�z�H��o�מz;���,1�m8�U�6��Ao$�N#��A�B�iؚP�_�n�۵r ��DT!�ͷ-�ʪ��Ungٸ��l㸕t)��1�w+�|�p31}`VYj���5{&���#L�=9�ק<pCD)�c��;�u�h�w��k֊גl�J�AX8E1��{��X|�	�x-u4zVf�>��S���8Tq--Ŵ��a�i�1+c+t�Hq�c�!0�V��������o5���:w�b��5G�DGʣ���-f����K�)���u�������ڍ�Wg���
��h+�V�^��o��������j�eǽ���oF<
r�,uWH�HG*Ř-�o!��j�w@ؼ���r�k�:����m1寪w����R+z��+O��g:z��S���!Ҭ��{&�B����-~�&y-/�����w�zƮ�j{_w�~��W�go݇�򔪞�P�������^hy���o��U���H-̈́��=���^��	B���/�U��2n�no�$Z��dZ��q�J��q?_�^�i���r�-BU�
�^z"1���~t�Is�v�����^oG�fS�{��.��ݵ��:�ۻ=���`���_l�o6(w��f��m��{�T[���7�'j�0�M�8j�Ѕ0������D��-��!������n�&��g�)����z�A�����-�u��-X�ڂ^��E�*X�d��[n&z���(��öХ��,|�"�w=�ޔ�GGdA��W2j��-g	f����)tM��/hZ�?l��y|;��de�9���9%ƤoX{�Wo,[��	1~����ꪜ���v3%tyz6�X1H������댨�Zy���?_eh쮍_V@���D�4��H~�F��F k���n��J���3��.��ʜ���9�������Խ����לCv~�c�I�q���HUe{���~��g����^���zp'|��ћ�bf7ԪK+���n�U��hQ�Џp�3�}f�����+�k��>�X��~�ÙW[������hPac����P/
/#ɣ]��%��R���m���]R��h+���ԪgV���%�2ފ]ۛܟu�a�j�T?5��F\����������W�~u��NV�Ñg�W��x�����ί|�Q�o�ڼ����%���:��#>����� ���r���ЋjyOȭA��t��8��|��^�E<��ϖ�)}>ރ^<x�6��~�$}���C��ڡţ�;��C�$>�k`5c�������I�O4���ɻ�Kב�˴N\�5:�o�9���IpJ����̊��e�ũ��-(�l���;O\�1�NN�M�>�{�%l{%�>�n{���N�����i����E7��u�.��yfm��B�8^Ȇ�o:�-7|�������>�����nq]��~�[�QZ����?�M�jtj��oi����^�l��ii�W����w����T�SΔ�{���S�s�߄^ظ�k�'N.�t����W��A��v�'��G:�G�i�B�l]{<��e��{�窣ԯ:e˦���jXE�{PV�	�>�J�zƿbLһ���ۡ�T��Ww��E/���+�^�)�+Q/kov�c+���ݼSs�o�5|q���ɷ�B���K���,�{J�(\hP�9s�R�0�W��N2�M]Ȥ�zU��=�\�¡
W���/z�,h�M��j� ��y���
13�Q��p���ůf+��,�*�Y��*�D��r�%�Y�Wo�^�~�#��[��Ț��QI5R�eC��چ�V���S���~D%�F��y��z+��I�
�
L�K��Q}ɗZ[��{�Ul(_*�KG|���h؋���tє�~f+���S{]��u�vQ[��u'bv�8U+���� ²��SݽKx�]�:0I4�<�}Fa\@�I�۪��Iيj��di���>�>���ƽ��-��B�����,�<�j!��j��q��m�e���z4ς�`׋7&���q�m��'I�?N�wyw�������k�T�� ;���0nW��N]�Z����;���{�����_s>|��~R�p�~�,?}ğr:nK���{N�7�m����f>pl�������%v�׊o���чT���S�׵V��;;~#���^F���#ۗ����TԟUi�Ԫ��b�~�W%Di鬪�r������pת(�)�a�{u��7���M�ӵ	�x����]�^KCáCRm��;�ռ�E�j'jQ�cs�ߙ�_�Z���.>u^����c������  ���Uf��z�Nh���������PӺH��0��+)U��58���/*�yzɩ�T���PY+�k���'���:sn�U�ܶ	[O)�W3C�7Qg.GՑ����愸���kp�n�]��5����YЎ=m����R4)dڻC_��<Lxv�Py���Hq��ׯ�d�z8�R��n�U-���[Ԃ��ӛ�4ї�K�(����tD}}D����v��c������+�B��{2|�<9U皻�97;օQׇ i{Í#���zS�J�쭭C��Y�~x<ꤲ���'Y�[������:�^n�<rR�^[�.V�߻o��{n�/��p�v_�O7�[r�뽂�����q���� ~N_d����jgk"�y���/=�@���>���Õ�r1ǃ{��/0��ㆡ�;�@i+��냽=R��}K��#�iz���P��՟��|}+��k����ʹ�I��կL�����>y�
���n��/�Q�1z]�j,S�[��e�P�g����7Q^��j��%q�J��9��#H^�>���%���X����c��^����q���<^m/k��מ��7I��p"��V5U���|����%�ޤ����h7Q�G�z�ʓA��_�p��)s�=����39�aU\�^���짽��6���c��|3�5+��az	�`�n�U�)�zL�H)Q�G/oөw|g3�7����f��]D���o����nϨ���Oj����ʵ�P���v4b�؃5�j]��.�Dƒ쮽�$EW����d�9�.��(��>�">�k�d���~��ڋ	��<��1=��n=V���J�x��q�$����'�D���Շ�����M�;�6�|�˩g{}�wA�KܪI������G�}޵+��p�|�g@�>饾߇�ߧ���8�ѕۺ<t�����p�a�]0�a��jBk{pV��%3M�ޛ��'��*�&��Fs�}o�ꆜ*��H�C[�5�^}V�]�Jy�m��ݐ�����:jŀ�'>0��JhW�\m7q&"��-T�r|��*�v+6�7�}����޼�6/�/9:�_��t�CT��/�Gs b�k�c���=�Ս�5�,b򱔻��L�tK0��t�u��p�+֟�zªy�~}�y���/\a�w}�?H?b���h��?b�d����>i�9OҬ�f{��︀�GT[�~G���R�1��L�j��Z����Z��GЄ�v�Ѿ��9֫33��([���W>3X醉T�Z��C�#jFk�lc��]I��f��|�t.�������#wJ�Q��j�j��)gPz;:�Z�/v��g��O_%f�줁Z�Ñ�h:E0V���qڑ��$2��g��3Y[X7���n�Nɇ��f�a�x��/��!���n�)[�yxV[N��ّ�Fm��`2�+��w��N4͑��t���ԃ��f��d�K����I�rɗP<.���"t��VVh�.nD郁oS�>c��*QVq�1�X2��d9jnF'}�ŵ��e�*�D
�]1�_m�)�!���}�����l��M�f-S#�Ðo@��k`�z"�:�VD{F,�ë�ԡRT��@���H�i|�V�ݓ�n�j�[7���5.�9��u�uJ�9�1��A��0.��)�/�\7O7�J\���Ыǣ�\��KFP��e�HY1en��,@�Tn�\�q(24�FGٵ���4ֲ¾7�ֶ��씥�q��׹��1��y>��̭��eb�L�Iѩ����أ�s2�������30��h�Z]�.��I����÷d�gL,�wR鬚��p*g��&Z������]$��Uf2��Fb�ֳ�����S�X�m|��(p��T�u�|:�5)���ռ��&�4����I����R<��n&r�S��8�t8��t{4P9ew��W�1B�������!�Y	����{+Θ�v���QʘF(�<R��WT�(r�6��u�+�3���or�,�٭�4��K1U�zi��*�h!$��u�[޼��c#U�����
觯�oJ�t��X�M��I����okGq��1����ls��PA;��ۂ�=�Me�F+O\��Ay2Y5��v�tei��16$��Ǳq]�2�v�rԛ���&�gaov���Qv�߸4M�
�D0�Qn�����<���.��<�Y��k�C�ռ���}#�{$,�Սb@�:;��+�sw����^T����?i���u
S���z1>�V�6�r�g:��k�<6��V�GR��{K'<l�Ƥq������T�Ȭ'�+��\6��f��ڛ@�GZ�o),(RV�S۬�.�ֲ��&�Y���}�%#h�+C��ۿ%��Ǯ������88��#i�,�N�;�s
Oe%ݼQ�����i%�s6��C�yn�Rh\α�����|ė�lrE�{�W[O�3��7]%#��
���Ŧn�}�#���Ӏ:�o�O��J�D�\dڄ�����1�W̬��FlJ}S��ڗ{]Y�[��9�l� ����طWg)�;ܮaQުg9�6�+9����c���%�M�_�44�D�j�)`�-h*�5gF��ih�j�mIMD[���5����h����!��*(��`��ΰE��H�����N(�b"��ZڍT�Fق*(�h����ثFcd,ઝ��V�!�6qS51A���E�A1DQlb

����lӵb66�QQLѠ�U�F�U$LƝ3E�V1�F	�UTӢ���EPZ�T��gZ�j���j�"�
*

b*��m: ��gXմ�U1�Llh&�����k��m��*��l��j��`��F�EU���(���Fmh�4�LU���&�Z��h�&�����ÿ߹���?���=�XT�B�D/�g�}�F/s-���X���|d�n|���'&,�$�>��R�jEa��U}��E�)<�VjoW�N�7ϓ��U�6���*5Q��?R3uu/c��5�|2G�|V.�QTTc�' Rz��5�y+�d�o�����zk.��[ۙ��,�qGq��N����G��Z�*x�Ŷ�ӯ�O�%q�x�r
W�p�FR�1���3X�Qcu߂U�F/^�J{W�y>o��w|��.��.H�OL3���O���{Ρ���}γ��ɝ݊0��7y�V&�V���B��F��n)�Y��+���X�Kj"�+v�x�Kko1�:[���j��aS����/o�ի��xuy���C�[Tw���w��[R&&���g��=YY��ޤ��8�;�j,+��}�5y�s�uYh�Tx�%�O.j�P����1��������W��S�Euܥ�˳/ճ�#y��n8R�<����ˍUP�|���jSBS��7s\|k�z*<h,$�2��|��ų��<��pN�r�%p_�Rڛ�l-�/����u]�oi����	W[�h@� `��o��g��m�o�� ok��oˉʊ�z%��ҷk����������uFk�m%�1b�OPٲ�}h��=��H�=b�.��U}��|y�����S��rYK��y��l�|r�J9�F�k0p*	�Ex�Ѫ�w|�|h�w�����S�P��y�-`��/F�F4K0=!���'�$*cO��k+��2z����#K�H���c)w��k%��륾����Yg���Wɩt�{}�D��������4�3b�ݵ��F��M��C.���a+�n*#|��~����^�G�qmv0}�լZ��B[%��M�U�g1E��1����BT�˼X�N�{�� fz̾�7̷��خ{����\���gk����s�O�v���$���$�(!5x��Ԩ��4'��r��C�\5�{��!q�N�s~������]ၾR�y!�a��8���׾K�+~n�`Td�\�^j=IW�Nǽ^�������i{}��9g_�|��(wW3SMeo��N��C�ikS��;V�ᙼL6�j�1M,M�ͽ ��!�"dJ�����-U7�blg�
�C!�1;s�Y~�ڥnG¶���-���;qkg3��H��1�N����lݺ�C)��h��RwUp.Ta����;���m��cۥ�.Z|�,�0v��@@��Vem�J��WG��G����e�V�Y�D:j��-ڏ'��ƽA�ui�����¿AӵA��3;��}Y�'U#;�ֆצ�6���z��k�^j�awI\1�+���52c�/o���>Z�O�KԷ�r'�ހ�u�M����R>�"<��F�u|�ܭ7j�XA?��*�cW�aok&��U}�m�Ћ��[x3mٺ���m�wK|����n��:#D��1��1V�����U���6l��cv*(m%����m+q9T'
���X�V�{P�̇��u�����g��a�\�o�=�h���t4�p��-9�e��u>�^�O��u���&��zrQY�{�W��[�Z�����]S� k��QqUKfv4�����|9.)b^����=��ǍC��_7�y��dP��U(�ohU��nS>�c�ib~(��]KϪ����G����k���ww��A��Q�����_�F��_�<��b׭��m������2�'
���cT7�	���ce�
�����){v�Ĝ��˩��c�8_x��u�S�R�u�.8�h(��}�Y@����Dx+m�YL���z� w�V��um���_�"�uW�>o�mT̥\�1ҡ�;�}/E�z��t¨���+��J�����Ј^>��WI�>t<Kո�A��~�<׷|]W7��ŷ};��TB6�Y���O�{�m��u��ǹL �p�i��so��q�w�Bus�ȷ9�k�x=���N��h���{~�=�4��_C����� Zz.W�)�B�زl���-*�3���9�Zӳ��M��-���H<�@���6{=������|{��e�C�á�'�ރ~>�[��@�I^����#���e{��+һ�xúe��7^�HT�~[����މ+�%��gly�U$uǜ$�J��w'�8F]ح"[�n
�[��΅�b`w�eo������i�q>�����v�SB����3�T�V������pd*������<�P2vV�K�g0[�60_8��q]9����|���u���]XwqJZ�������}X2�;,J���3��W8=�v���U�G��FWr�i��Ԯ��p�5��u.�n%���d;i�MW��Jt]Wq�
-���=�f"�հv₷f��A��W�}�U^��օ==�j~�Cc>����2���=[�ޡ�]�k��	ئ����ؽ⟫��)�v�~��c�13��F#D�	ĵ���T�a5�J�͹�~A^�~�y���=���;�/�_y�A�ź�*�/|UX�^Q�u�[`X/�%^�<�Ԉ<���s!�����8��y�}Y]O;�-�Bp��=��̝^������^ef���������:}��#7�@�[gkm�A�~�V{�Ua@���cQq��7�ό�CW�{�w��Uno�����c�Y��#~�{�=��~^���S�j�v�'�o�{��y���T��tuբ6��y%܉�~����D6�]��Ƙ���SæO���:EoA˯%[P�-"�E/H<�$�(;l�@Tl�4��#��wO�n�=�u�������m㞏{��8ׂ�3�W������*�򸨺�*�ڋ���I��J[��*��x��I����w�-�zÊ����p����6u/h�M�ޱPǣ��O��e-�	��u*�`r�ݯ�0I5�x�P�v��\� ��]t�=�Z�Y���j�;+{z�ʎ]�Gﾏ��>&��Κ����~~��������c�׏W�Q��κui�$R�>�K'`��ץEV��k�Ս[�_3���������)���T�%g+-I�e��X5y��9�/1^�T��T%W�,�#\�&+rjf���S���%,7��-�'�r��g��}��j@�;�=����_[B%O҆��!
��7���澧������n�T�����W�9�R\��"�_��x�8VDk�U�h��L�����oر����
)eI=r*�cS����k���=��~��o��|��;��s����85\�^eI���Uu��pwm�~B�� g���{�	.�s�;oN��.To}�����Ju�x,z���-Pe{/�Y�S6^9�Ϻ,]�Ir��S�\,�w�r��:�?j���TBO���^A��Psɜ��l	/^�8-p}k�;(/#Rǹt�񠼲��v��9(^1=�1j��84p5�:6me*;�U���WsS��)JUػDV��WܺN�O~wCLh9�釫h*y��Kzξo0nR ��t��Φic1iX������:��`X2�b�?}U��WϞ{�����������S�/Ӫu˷�X*���Ƣ��%U����*yS����o�7���W���Ш��G�_��}�AS��h3�ks��_:[,��s�:���=��iorD�}=��M3�Y}^�rp��ת{r�����o{>�s��s�P��l�Y�n���LīPN�¥�����`��x����m>�f1�W�Mތ��a-�/g�nxD�J�k\�|5�u��=�h��=$}=�j�2��^ͪ~�h4���*��kR���x;]�XP}	��7��6���;��{� e^i�����/٣�(���O!O��m,����7����߶�ɖDQ�=>'L/<T��O�6�\�]D �/s�+�mA�β�N�es��+���7���od8�UD�j��[�ȅt�V�{@,g%��/�^��YVY���:�X3�т����i޷H�n�EjDgaF1L��H`����^���֦:��ڔj_|����n!|���ä%�^cx���ӑIٕ���x�)�jq�k]fwu�#:�>�2p�O�W��}�{j߶�����x�y�.�T��q�����d4�@P���,��9�t��j� ������X���13�J�K0��t��(t~�I^�����)�zx���,�X������19�~�ƊP���F�(�F��E���ڜ��Gj����׷�7堥Խ�O�Tά~>�!�x,��2
QM�E,��{oc�u�r����T=�p�_�/uu.ڦ<�z������UX��������~��+��%p�m���F����F�!�(����r7ʌ_��CT~ըT*x�ŵp�7k��)
��n=����J��'ap\����hݯ�-W��G��[���t���}�n!�
,Uhih�R��=j���P��\��u��'�z��Rܴ�)���M'�pكCT�P��f�؊�����2�����ǫ��9�Ǿ.�v����8����ۀ�G��:���qݩ�����5̻��OuK������b�3d�����y�;H��S/!��[�U��&��,A�#;~�ȵ0��뾱ϔG4ʃV���u�+8b��Qu�0�*T#�6����������[hG6��;p�
���tg�U}U_=�k\�k��L���lc
�%(ͅ��Ѻ�?^��"LvVn�X���!���hP�����%���cVz#7���?U�D�qX>���2�I;bUc]�� cU�}P��O,E%1�CU�`��im'!$F�]f��7��(��{2�U��~���DZhPN=��T�V���q�YFyg����-d��=|Q�8��V?\�:ey���p�
�W�y޼'MS���pg	�y�k�Vz�<ߍ"��`��z:���C��w]��h�[��~���g[?z�ny`ذ�x���?;���=�w����ke$�ga��F�gCYul7��aZ��4뵥G�)��tH>�Ō��g�)�R�>~��O����(	[]�>��`����k��q�t��(�}Bv�wyt����w+l�<��S�D�4`�嚀��?9���Q����АlC���b���ŕ��>Λ��4b�x��sے[ۢ�GL����%�x��o��9>Ό/�ͣ��<� ��х��y�&����S����cM�Z7E�Ib_&�{Mt� �(�w$�]��?�}_}��99H��uԎ��h��������G�f��D$���M�z;�3��\R^園^N����6渆[��c"��s��a����G�kէi'J1	�����T�b��"��G�-���*�F�����E}u�������E��#�w��#��zy`y�59K{\���Ymí�p��;�^Uu����c�~��X�V0���8֕Dy���1�w��+��J�P�q�r�Y �	�����L�R9�N֪�A���������5c�?;�k�]0�a"��o7��"�	ovpC�O�g�L��|��{[^��TK��%W�,�P�m(��1&𧾑�;�OpW;�PT�+ig�<�����*ϼ��aڔР�j��n�Q����x��w�z�t�] ���-��i�1��fA�V��㾠�t��76��M��EE�z3	SQ�^��0�y�_����y����ZI��O��-���Cx��K�Y�������H��hSMӘ���՚��,u��VD�ɭ�6�/��CZ��I����+3dۋ��$`5����2o�iAg@��.���gI�5	]>�8�)fl3�bp`w�`|�;�wGk5q����6�I� 99��U>7����j���I�{wGj[��ύ[
���:ڲ���[�����ٓ+��4o�T�0����҅un�P��0M����j&t��8��M�.�t�+_Q�u4���ZWJ�J��헙̳3����K3�µ3�N!������yJ��E�/LjЀPyu�m�b'��](3��cy)u�����2��i�M �p�SP�Siax�O+�G3�Q�L: X+	�b/��o@�%ӕqu7O�gV��x
�o����-���"��h>�cU���P�bLGT�v
���3�K"���Wu�4k�r�1�� I�II*W!����{��t\��y\#�3-ҩ�u3hP���V뽽	�8K�1��y��Y�� :H9�X�H�]&�������k
���s��HS��S�)��Y[��%�k--��<�oQS:>:�>��\ �w�e���|��g�]���q1[��ד�R��}+�0�ugܺN���Hb7�����Wv⿯��wm�7R�]��5�����߭k�#z#}	�2��j�m�l�gW1�t[ux�Ґ(6,����g�ݣ`S����}�� h���wr�̀��S�x������_n=�v�G+�Eh�ֳ�]�Ka���9=j�Bpvm�G����G]��wޮۼ���nҽO#jӭ�|C����x��Yu�����r�M���z+1ਪ�,�v����b{
cNBH�L�9x�PR9�l��^��'��]BE�c�;�c�8�)G���]9j�Vkp@F��<O�����w)%�)��� 
_5g;iҷׅ����UЦ�X����F�l�tx��=�+c\+-�P>�ѹT�!ϴN�t&�ofS)U�}��jVC3�l��4f�����Z�V�8�X�e�F�
�!�z*�8ӬW�1��L��@O-� ވ_q�_j�4��/of�u��f_5y:�4�68v�i���9,u'���fe:Ӷ.�f:��
+���ݔ��e c�|��E�"iRWδ���m3��\r�k��[J^�Ω���u�����Yz���΋.����4�Hue쏭���k8�2\�.2�N������mj�+uWnQ=�x'	ᥔ9>��Kn�v�إa�%N��]g|^�A�����BL�-h6Ç{7��ENA��i6�C�An�Z���b��Bމ�k\�y�RԲ�w�N�c�<WWv�Dn�a�f���y}7����X�i;O�q^B�Ŧ�$��Ժ�7�j�U�p�=�B��2A����,"��K;Gd� րCo���9�����Պ�#|:l�gLe�R�鉀2�IOyu����v�p�)�!���E�f���L��|���&he���Փ�巐����P��0I��lkUM0hѣR�b�*��3IEES[hֶ�TDDE4�1V�
�5�`�F"��d������։�t:
"kcPC����'l�SZ�m�cUTT�L�M$DQEU4��Q��������"��������(�f��٪1�ES4��PQEj������FjF�F��cl��Q[j���ikAZ
��fht`���"���4F�4�E��4�bhb�&�b�6�EQX�h�"�t�AMDUD�TEKE1LV�TQ����:��ڱQ����h�4�hc%E13�U5PQ5APAIDE:L��j*�j*��J���};8��ŧ�W+���]�,�#ʂ2<�l)|��9m�y�r��6�eN��ܷ�w�!��*�R\ 	������>��=��m��爊�eoX��X 뗾�&�_�s�b�;g|�	zaS���c�ޙ��~�����;B�� 5��3��995KǶ�k�؄�έ[�J�S���Ѡߕ�z>yMh�
$���p^��Sm�\P#}��p�8�����R�o�;�8��n�϶2�笭�� }U9_3U첧��|{X�!{~]K��-�}B�OEC]�~`���;~���5�|�O�\�W%}��n{/gǸ��m�Ŏ󧮳oU��Wks��\4֋��4&�ܮ9γ��p?{Uoqs�b��o^e�#R���H�y���O�E*��_@u��L/W��R�z6�2�>�㨆��OX��)��羚i�~���{�\jk׍��ju��+�jUg*ݽ�W�c�Y�ߛw�t��* A���5�{��I�zzI���+Գ���P�x�o���4��N�;�>�':�r#��,�@�ȟ`�_g)��MW(�vgK�#iE�ŕ�u�q��9��]��ӐA�K���W"��\����}��]uƭκ*e�]�-�`��45�Ұ�H, �T�9M�㔰��M�؛j���k��#x�7
T����""��������m�����Z#Y�:<�B:��<<�^�u¦i_=�w��M�e�R������5L=���FTa���饹�)��������.����O�$�}m��w����'�E�����1�<rr�X4�`�XŒǎǆ����%d�M9�?Q��I¸u>T�A�h���u�y�,�N<�r������8C�#^�1�Y�$��᥻�k*���mvߤi�<w�7�a�z���m�8�<�q���y#�V����a:a���gׅj�RYX����dn8�{}_�w�r�91@��iF/0�ݠ.���@����؞���o\u���Qo���ib~Z
]K�O�L�o�;|��qF�/!/&JQ9J%Kې��'x���*�{l�k�^���Ӟ�@{��t≕���5Hjx��<�Y���2u���c�$��o�2����j�|��S�1yM�W�h�Q0G>��۬���YV�;PBa���̶��L4Ut�������x�̬9�6�+UQ��^�S�N�=kaq>��
���tv뭼���u��f�Kΰ5I}@���-s�֤�!�T|*�{�����?}_U}^=�V�N#o��u��<���*!S�l�[���Y���'()�QH[�b�D��[�}�n�t��<GO;��nON�ow�x�_�����ם7�1�\�^\����W1�[�kN��;�~��Ϧ�]��6��j}�Xv߷�n�=4/�a�y��uǫ&M���t9ʜoٹ���Y>rh��;�s��qc|�7�l-��J�6��<���kLς�3�p�+ɴ]V�"�-�G��W��C�F���Ɇ���"彪���c���Y��=�\�VqOU�eSo����m�wz���H�CU#_����[�z�+ҼƳ^�qق�'Vd:�9g�õ�����w��r��{W���VN�O�Ӄ���+w��j�AՏ�*��NɈ���J3q{�����z���@z��:�7�1�UY��Qar��w���~'YC��u�E�ez���ƫw�lK*�Ԁ��խ���#>�K� G\}��)�w�e�r:P�KTFs�x�Mk�Y{QսeӅ�d}.㪷	9��U(���sr���n;p��4=4��,!zB�DV�/Hm]󴳹��;�]�����+��>&���ﾌ�Fc�����˸?B�A
�t���O�ׇ1�_z��v2�T�Z��f��w��aL�G����[�Qv�س}���T^ŬO�8�͡�[��k���u�vi=G�>�(ǝ�����D7�Md�.��G���0�{�y$�ws���]G�?R�o�[	4���v=�}�Yt���ۍ�:z��ҭ����>��k�;X����P�T�\Bx��#<���|��Ӯ@�qO��hy+���krB�=8�ݯ۟^�H����k^<:�o<�Y��2[v���~�yk�6����MdY�R����S��M�T�
�+[S��if�jٹX�2�P�6�+�⾺�5��Ϋ��O_�**��j+��ݿ�ܫn|�gA��&5ca��8b��f�'|�=̜���H��T�%�G�ߧ?q^��x�f����
�?W���֌��<�vJz鸶utf�*w�\�ẉ�sb?,��ҩ,y^~��]�K��t���h)<{ݣã8�p��(���������r�-/%%��<%P���7�S�H�u����nd6n�F�d1�R!�][�뷩̫�v�_>vF������n���b�Y�Y�E��˸�[��5����ڃ����e��]}%��P��7v�3TU�W(C�N/��E�x�yp��Ҭ���P0�JhB������j��K͜�����}��삮WG^��~{K4�	��d��j��͑�ۦ�VO/K9M?M�q�\�O��>i܈�{����{~���vm�5�0�Қ�<�Fl�6����� ��e��UC&�H%�~�����4pf�odH�S��*0����"���`p��U߼��*ҽ�П{R�Kc��Vk���j�ڏ����ͯy/b��ɧְ�!�/t� M�	Mm{;���G���(��F�qI?+U�K�8��G����B���&׽�$T	P�l��cH^�]K����Yg�E�i�s:?{O_w�a+���Rg��>��#}�y+��g(��Q��Np�.���K|�+��!G�hY���ƠZ5l�fե��c��jj���ȟQ���mե2cx�Ù��P�z���,�7���^)
��.�H��4���e�Πo��6k��ƵM�4!Jc���m����U��w.�l�����z@��g��>����""���o�����N�cA
Z�@�{-/N�AU�u���p>���4z_� ��y9_L ��w�w.Ϋ~[�V���ѣ%zۂ�(Y�Y#U/d�8�U�CőWM�Xko��G��y8�������w��V��A�I�9!C�¨�V{��G{�h�MI�5^�/K�Q��<*5g�I�:��Y�k���_s��[�}��>D��Ty�-s�1��ծ�
����k�Tg���n���Cn��cVz2�E7�sKs2%2�T�}짯�:���G�_sVϾ��̈́��'
�ܘ�X��2���~�98b*���9�mk�.RW��7K�9y�v�ƺ��6�n૦cD�� |��y9~ϗ��-/F�{s-�C�v{�,1�)е��Cu\������y(��|G%]S�l�}@g�/#��c��DmR��,�pbڜ��x,�#�1{ffT�<����{�$�=��T�M��͊ި���J�ooK��bG������RӴ�x��C��*~��z�&�A֟A,>�]���	^��V����wPp>��!���Y���0\��k4Hn��o76��x�΀�r6b�~�>��5��U��;T�)�^5����,K�a��_<����պ7:����t��ެ����!�}Y��k�w���g�Z�������~ΧO�.YZT�����^qt�+5y��V�����8}��^q��5�7I�7�͚�����S�
�?jM<
�Z�=h�[C�\?v�
�V��(��]<���j��Y�s�Z�*xڵ퇾���γ�XEn���\�l�){��?[�cUE����*�*?^�KJj��8xe9�[x���W21����P�����i��Gw���}��G=>4c:��q�9N�G�=����euv�0�xh���qQu�Z[�I��x`5���F�[�Z��X^ի���?y����l����]^����&���h��`�?#5[$bI8ި��ڋPݔa�:���
|�-�(�:��~w��
.�z�8�J]�w!����t��$N1�-35TG]�t.V�N�@
�l�z2`U��=v����]�)9��wm][�s��6g^�U��M�w��l����vTJR뗐e�|$�&e[f���+�y�T�O�op)���ՎJeoK�`�*(�W}�}�x|�S�mU��`��R1��|1�����Z�8�Y!P�*Ox�G��7�_Gݥ��_s5݇)�V)�y���?y�����7��#F�4ק��u;�o�YW��-���g���H�X�q*��e�䟵ƺ�n�e�E��c.�Y�T�� �􁏠�^�"��a.�L�yE���N� ǛP����y�>0�n�\������ُ�+�G��~v/��Ӳ��=)Tyz�iCe�g�_F�m�q���z@y��ɇ�o��M�!�A|���`KZ�8�&�*=�#J��n+|��~�4�����~�/x�kwC+�dIw3�<�w{Uc�uq�#��b�'�����z���X/�����K_�vw#����\5����!{iuN�c�i��ӧ����V��^[���z��^�4w�>���w�\?{MeQ�CH]�G���?��v���>��Y�N�糺Rm�W�1������_�Y�	[���em�t�ti��c;��
�)v%�UD���q��e����zv.@Os���+sN���P��j�-zP�մ�z$C��jGW�t�a�IO�R�����Z@�
�����33�,�1d��
����l��>��מ�m�X|*=Z���y�?<��H\mdk"��v�����7Jt��/^��S|}�_w=�6q�|Ͻ^ݮ\�dU��ւ �����������^>74{�綍%Z�k�'����n��)\NJU��X={�{�C�{��~sS��z*ߎ�-��P����Ʊź(�E~ģ�#w�����]צ�7�v���.f���?#sKp�&b+�U�����(k^ ![��w.Y=�M=x8�޾��
|�-����T*Q��_F�Q��йӢ��;��F,݉Y��A��	S������Z~�*ų�w;G#n^5�nB�ʯ�cU|5ï�������� �`y��\�#�اfH�l�*.מ��Tz&��1��y���.
��c\���O W��+�����t8�,���㰻�n�~�%A��:l�SG!� ͱ{YrR�T�Hо@Y��pgn6�ձ�̱�1�*��`Mg��T������>
�b��'#|E�n%���YCZߢ�E���3C�3�{5!�G���o�Dj���֯� �I��[;���C����&��Q�w���4�r7z�˾`^�|��,:��d�s�
�3��}���RΗ�z�q����BJK���UL���L^����+u/W!����pZ��ɣ�v���0!���_�#�~]K�O�eN�Qӊ�]4��4�v��e_�����v�V߅鎫�g*�kB���]�y%hFJ��Z��:Q��Y�8�C|�?�qs�\�#}�=�}1��F���#���h�{�}=bNթ��y�>ܝ8ms��>����]�����ȵɠb��w��k�{�����8���~}�Gϣ_q����5n�o��e�`�j���IB�����A��o"��]XKo�ז�Ǔ�_эz�:nMLN��6�RNݪw�8�u��	S
����q_]&*--��Z�{����~�k+&������n���ʱ��q8�Ϣa"�Jo�B~��4�Ԡnn+���)�x�����+���v�5�<�b�Cn!�j���c�O޹K�E�� yO�fM
�����7x�s���Z��z:��p����"%?�6�>�8����;ڑ�O��|�p^>�+�7)�γ;���Zn7��b������F�ww����9��g"�-���gm�l��f�F����1^[٘z�R�,�������S�V:���@�_��^�=}��d��NG-۫�����:#�s`'0���R��\aN)����I��/(��!2���;KJ��K��u�j�x���aq}���-�K������5���;x2�ȝN(�L��U�I��`8_5�yg<k��{t����1���ʲ�I9����)We�?���`#� [����^b'��ew��\�tRyQL‾r����M�2�Yk^���0R`__�u��N��]�̭uʣ�޳�U����>�}��������2�*� �����ǪکV)�@&�7@_R���[���(�^���V�hW>�qm*:��A۪����f�|��5��7IE�0\ِ	���++o8� �Mw;WE>��i�O^3Ð�����u���D��V,�g����Ҭ-t۵j�(�]`��R�T�S+�y7�$#^&��&�u�v��s�ܷ�u_uY��"��jM����l�ej@d:�b�CѺ0�p��
V�uw{���K�3�������N5�wXg1����)���<!�t6���Q�U�)�@�9���`��wBL�(@�,�@	@>�u���e�֐�c�-��V�#eM���XEo�m�v���u��62�Uތt���@�nd!�|���6Il;��Y2�^D�B��4�W*��7��	 &f<�J���[Z�eu�����\Y�ѓ5�Wƪ������hi\�Vpb�H��:�����CX�ysW58%���.�́|�}]�֠6�;}���M�lːm��{}�/�q�zCv{���Į�x�*�hK��,y�L��t�ԍ���[-�L�x�1b�9�0ҨႵ}��W}5��U}����O��;�"[�����}; �\f4�\�(]��������	v�z��7�q���0�]�ğk�Z(�]��!��('��:/)1-b6oϿǸ�|���>SYX7*����
i�wZ��$h	&v�p���l�� Lf|9��^R��"{���{f��hM<��.��t��5ʮf�Z7)J��6eu_7aǨ��	fn9Ƭ�E�֥�Mn��w0
�O�P��İ��#GN����7Cw�ulҕ�Cӱ�VoF�+:�$j�'(�[3����:�nn��gEEhd���j�4�5zX�u��C�x��j�����f�p�4��#Um�xX��QA�7���Ņ�	�[�͓{�cL�LLC7���d,���m��}�)��Q31w�4R[h��l�RѶ���
����i�"�v�Q%�F�CTE-D�u2P1�j"�bZ�
�m&�l����)�-`������UiѣMLQQLi4��A.��SD�SAN�KDl��4Dհb���]&���LZIS5LAUMPDUiMl�%��ETɶ"*�*$��

j�6�E�m�������CF�X�Z�jBb�
5��Tɤ��	���Zh�Ӣ�h)
��$*�M5���"B��$#`�DS�1!T�Q.�)�i�L�ΩѪJ*�))���Z

!��i�


6�-USU4�Ik$Q%5CMD��4��Q��
-�ѿ��vf�ep�Z��45�C�]@r�<�.����� �*�|G��HJͮ�p����\Q� �u���Dw��DD_�=�N�����&������	8U��i9��KW1����ˇT2�cP��;}��63�q�|r�u�!_�xo�r��K����H��Z����g�2���ĭ�-=�>z��P<}��ʙ}�OY?+q�e�!�/�4�z'E��ũ��N���B��9���`�b�13�J�D�&�yi'�L=�2���9E�Հ5KY�'��31\f���P#ŷQ�c�����������r	��Mz~�ܯHW���~E'�K�y;���R�x6�3��m׾����]E��Ь�^B:�u���sr����y�o�F��S،\�t�|]/ko��*v�N��<Z��%q��{��G��,��Ğ�2yb�c����eyыը\~�r�}�W1-B�P̼ؽ�p�j��eC�e�^�G��D�#�Ʃ��ە����ow�'����'��Q��{5�=b����gJ|���	΍�p��R�C�^݆+��=lwI��a����]�����-HR�ͫ���r]HvuX;{Kį4�v5���޸sl\ǽ�y�5d�����7��1@�;Pe�o_PG�\���f��+��0s�U�<�g�GWD}��c�N��
����>[]���?s����{�+s��b��
xǦ�>k�3��C���w=���������:`�t�x�N�V=����{�3A|���yz�FN��¸���齮����\����B'�����zA�k��{�?N���JYwO-}b�B���R-�~ɚ\�z�OSF�Ը����X�.���m���j���������A�
Э
��eS��ޗIe%�'{ꂣf�����U}�U����8�)4�"n�7f}�*Χ�
�B��z�
Y^�\^{oy9޿^|:-C�g��3v;�g��۽��/}G���](J�R�dyXy�r�زA���W�W-H�'�F�,�R�16R�
�CtǕo�7���3A�zq/-��OMa"�KɁ�X�u��]�'��F�p���9����Ѐ��P�c�G���9+H�)��b��N�or�>�0�L*B����75+I�V�UI�~Y�4{s�3��-ɹ\�Ǽ�A[.��E[�f>)��H�.so��a��&;���R�j�O$Ǌc��Y�����z�[�:.���wE��p�TĳՅu݂j�É!��PO����>�P^~2�������o�T����w�w���4�GG���>� 5�>މy������G��f��Խ�Բ�P������x�%��o�;�o�v�Z}���;%Q�؆��s��Ɛ��K�v�ǖ�P�ӂ�I̗�mi��F��wO(35<���zN��J�e�J�P)-1TXz��(wU���7R�Myg�&G��p��M��:��r�o���~��H\md������ש�Ocov�p�k/<��Mם�K�$����r/z�M�嵒P/�\�sٻ�x�j>3�42��j�Oz�9�>�R����w��+��K�(��YC�c���ԑ�}��*�;�t������:y罅�#Wa"@z
��~-ZŖN���/I�}�DP3�w�d���dz���`���}#z2{�ԯ^���wվ�F	隗�we��u\D�t89�)�Ͻu3����H�3˱��t ��gZ�4 G�q�"��+�fnb��grS�?f0��K6B�r���y��+)e����!{�̥3�[��.wj�G��+�μk�	�+{f>�����.�L����ݺ�����n�G�]}t��+k*�mIa��wgva�~��� n�@��2�u�M[��&ʩ�����GP��ߊ�x6��~�F*�U����E��J��s���*�(�2���z�dTs�f�U'���j�/ޮ���}���D�?����BW��g/m���r�����Fz�����(��d1�5� �4��G|t���T���/=�VW�ö`��������Nzi]�Mƪ���x��_uT��3�rB����y����'���q��Ա�;P�̨��Ux\G���i���WWM�"s��-�'�s�L��x�(�WzAuC���o�
:=��0;��$��W����3�}C�]̎hﻲnx�;w�Y�뭻���'�S��eϮ=޳�㟨N�Ω9>Y�br�^�q���\y��91ϐ�Y=�x�0����O�3n�y����q�ޢ������zBϺ�NW���2+e�ξxR�x��-��H������g���nkV��ԪX��nD!P�H"-�o7�D	`�UL�]ҭ���U|f^�g��[��]�W-��Y����.y�뾿֪���%�gm	=vd���6�uZޚm��ֹӥ஭|��*T��-3|61�����ف	�`<Xɕ�����/~�὆�`S���!cj4�K���po9������4��Cs2�+��z墖��=�̛���A�y���h��x�k�1.ѹ�k�7p��F���V�f[����+�W���޹������	r��-m�Hd1ҽyݝ*d`ҧ�����d�o��J�-�\�UK�D�5ĩ��R5>��2'(�p�h�ه���w�-'��+/F�ԗ����c��}���]Nxa���؟X�>��v؞�e�`�uᥞ��oϹ�]��g�D䙥SQY�r%Ҭ]�d�bx:�̳7�C����0@r�q�s;Q}���xys�ɥ87G_�Ô,�d�W��l����}Hņxi��L�������&o�RZ`��= E��c�h^xѵ������l�K��Ec��D#�t�B�.uJㅞ�w��dþ�7�ͭ�V4�ߴ5W��=��7{~5�#�-W������>�U%�B�(S�2��*�����b�f/�}�x�waU<A_�L��O�M�u�A\j{*��D{+���~ ת
�Wt��8O(��-xw�渼��['�WL�J���!�pO�q��{ߡG�n���e+Ƀ׋)�"�<�]",*��k���hZ�]�����,\GmW��#�דq�(��������l(?�Ͼi�竻5����5��{��wA����cqd��]��ue`�K[��|����DKH����K�ľ�T���y�xtja�}��3�8wb�%�M�'Sʋ]<�z����-N�вC�£I>�\�RL��W%Nf�5����y���ȣ~���j�8��z89����w�%x�q{�P+;,��9��H	��݉�j��?FR�e�i�y)�wc'����f|���m9�1	�t��:�!ud���y����R�����تG��$���\}�`/U@�on���/8̧{F\�x���&)ɿ����nܩ�.K�AW����9���;НM3p�����\ɋmd�S�����]\�	��6uyA�v7L�k��_�������|^+��v��L�j�2��#隋�q��7�m�O�&�LӭOw�eT�zT��I����u��|@���0;%=�Y�pXr=��z�g���kϷ���dWB��Ln��^��<��T>����k�sp=%�(�=��F.��\��8����~֎�9����y�X7z�^��/�3����B7�33��o"���y09����v���FCS��9=��������\�i�n ��"�zF�w�/�w^^]or3t�uvO��쁗+��D��f��̮���ygF@���a�ޑҰ���zTe��q��'@�fΚ������Mk��ȹ��B�r;�Mc�zÇ�D��{S:���(�.|Zf�\y6���p�U�ZK�SA��gd����b���W�"L'�����q�nMN��.������f�w3J���w�õ\�G�(w���b�����F���C�� w�~�����>=+�Pw����.�AK����֖yӮ�ѥ��/o��<5������ڙ(_ό�T1u3_s���8)߉��=����k�ρ4#n@��8:3�]�/Pq�&2���pCU]=�/*dW����Ϳ�1��V����:����.U�S^��~%�h���H>*g"6��M����O�����5;MULr�PQ���ܒ�yՅXw�tϽ��OE�q�!��1��i̘F���쮙�����������d���l9��:��ؚV����������m��q���=��\G���^�Lϫu��C��ͻ�:�.셻��u����XniO�f�s��s��4z�R�s���u��`>�q��SOO����n`X�p�Xq�B�h�%#2Wy�Ю�>ѐ�����,�Q���O�,���f����n0�3��dҏv�0��s�묹���U\΍��2�;��q��6�nf�ȃ��*�L�/��OU�.1�oU��d�d�<��7-�m9���n����v��!��t�̺�{	*g�*�G��ٵ�g[Yt~a=�xՙBdX���(+R��*�MM�˵���
�f��A$�w��°t��;8�J��hq�Ju+X��0��:��ɽ϶`bi�Vں?הw?gW��2<�B�����heI�e>w6�d,t�M�p ]p�t_�zK���'�O|:��'xC���˭�kki�h�������w�������a,7<��j��$�^ޥ;}]q�p�`y���ԫ�=������/OHe���L�7<u�����7������spx��?uL�Ӊ^s>�z�����^�H]S=��7�<�o�3�OP3�;�̜�h��a�W�P����1{�����c/�D�gzC���e����K�>����LĶ2���b/��9�#���}�FMER���/�A_���U1q 6�L���5���"n
����\7ѷS;_^;x6�k'K}�����K�[sǇ�U�ַjj;C(Ǉ\l��=s�S5ϲ�*'�߉��{�f
�8^�EG�N߲|����}�=���~��>�h5��E>2���9���� �5��N���%q�*���c>芫��dx׼#��OE��k�S��WuҨ��������_���|wW.�E]����TК�N�c�l�\<�z����x�ә�x��'8NG.��,�z�����稥`uɡ�;�Փp�
:=�z�W�í�9q�{��p东���|X���,������1{�_hJ�.�a�c��@N�w��NɥLn��XԊ�UeWQ�w,�m����hV�۱*�<�W7�S��E�u��lVf_u�؂���q�u���7:�	`��hV}I���z&��N��GY���;l�~�;�:���du؜�uz�>�}:4�>��j���7g��_��$��6��������z� ��/����|z�:�Q�<fw�a�j^=�=�y��'�z�x���Ҥ�t��)b��=�!	�ƭ�E���_z�ϽIM�!��g��/7����]��rظ�u���yO��]Ҟ��S�(]y��T{=���+#�U�OF�'SL�e�U\z&���3q�S��hm��]$/Y�[w���~�7��N+5]=�����#��0���f��\�Ӕ�O��ț��'6����.���;~���^N�V�X�{Ð�C���N��8��[
��7:��]�s"E���S�S�`;]��ﻺ�� ���=� ����#��fj�0���`��~_z�e�W��<��?����qS������Շ.�v�z�U[tb���F�=2�TS5�L�*�����:�P�}�������.�������z��=;�%�R<M/BxJ��Wݙ3j&v-�$C�>�+�ueuu��V�"�IP�ݤf.v�s��[W�
���u��	�*R�����a.��X+��옩��7�K�H�R��p̳ĉ����i�SM�:��5`��O��`��*�о�b8��_v_K����T�Y.��U9ֹ`�F��a^��1��8f�����ª�g��
�`aq=�Uf������^�y��*<�U�m9��T�>��P{�dv�|8B7j/���ͬt�V�ɤ8vT��L�C��A���޸~��d� �T>
�����>E�B2�1~�r�n7���J�U��yW<�'˨pzn���m�Ƀ��,x��|?��_��@zʍ�;ԅs��u�q�א���w��r�ټ���k�z����V�O�#��9�!Ԅ���fo��M���S�w���4)�
��֞�16�����ʏvY�����������������~���E�,�z;�ht�{ؿq��^ў��3>�<�_Iϛ���T���:!,����~�ܑ�Us�CWv��XEx�Q��Y��	���2��ї>����MS�n�;k�]F�;%��xsO�(�4�r�F�*Wi��b�F��������oL^ҸhZ��W/o���2�׳�;T�>�Y�D<ve��gy^�r!���ۙ�!̿�EL���2&��f����?o�U��{�����Ѿ��B�x==�xw�ί���ny�˱q]L��WS�:ʻ�Um�υ~���X�(_cu}*�Ϝ���{Ƭ���=H��#o&)�Y��:��p�w)�Rf�M�(滤�����Y��z̅���˫7H��^G�]Y�E��$V�K�����lRH�,��q�8�XѸ;���
����9�n���J��[ԇ%	���m7����t�����
k_Y�+b���<]��hއ��[S7zz»������b����f����u1�����gL�e��>#���}a<83a�3� ��O�Wu��})��4)�x�su��?�E��wA�z��]�Ώ'i�%�Xi�W�����s��t:�kka��'Q%����W����G:�m��l}��)7յgm�h���SjU��nRy���96~\]�Ӊ� ��N��\(�X3�� ۭ���w0N5�w�7�E�qMlĹ��B�Q���En�br�����bf^���z�s2��-j�l�X��.Fb ��/�7��%��.���>�槼!�LV_ʛ.�G.����u��7�싾7�.~�Ξs�V)��᤮�K#�
��s:&v�\�k�MܴK�pinst���P�����p��$��Eݕ��fi	�����n,�]
�����_]�	�|4�S�*��v�z�N�ݶ�c��R�q�SI���`��\"��jѮ�^��a�w�XƦs�¬�ɨ*�۪N�1��(h�hVer�xo�����[:�V-
�Yz�Gu�4���9�j���z���p��<������:s���y�塍����Q}Ni	�ׇDd�M��D�Af��vN7}-�C��[f%�խ��+6��\ �VEy�\�][|�v�ctS$���Jެ�;OVfM(���n*녷��5�$�/)�x���v�l7R�	J��+6��ݽ˟����%�Z���a�W��u_.��@hT���#�ܹ��ܧ>37Y]�0�v*l����d�N�/�T7+��q��|��,�z�h�F\*���+ꅷ����[V_[���˃��-�\.�5���:�;elTh!R
�]ݚU`��7~�
�Fӧc6.H�Z��N����*Rs�鼹X�G�9�I'vZ�-�Z�e̳վ�t�y���Ab��R3�|ӫ�k�۹���l�u�cZbjvo%0�Nd�d�#w#�]wn��V,�IQ�/�Njy��b�x/����3��X�^ed
�)&��Dh��c�D�L2�ຜ+�\�[�6�rX�N�uֺ뫑�~�LT<�}�k�eۛ}}ʕ��3 �ʜ*GT�.��]G�Ķ�4��	�ɟv�W���qA��T�4��*��Vs1q��S0�B�����bonsF�ӫr����/����Xgo�{x�s�WXTk�^�5,v/�u����ۡ�̥�!J^f�&��Ӫm�����Y�.���S�ྌ7����j'�m��Ds��U������B07�U��+����'�Qŭ)�����%GL_ns\����u=���E
�@S@h4N�UTQITIT%������i:"ZR����(u�*��Ѥ��b`���)���[�M.�:t%4USlfh6��S��l�dhbi)�Z� ��j"�O�4�B�6��3D�Q�qPD�Q\�čIAAEM���AT�E5M��h���(U��4�TDI4�D��UTP�:MUPQ��H��JZ����h��֎IZ�"��*�(��Z)�5E0lj�������֔��R��h�6tƒ �f��H���T�PKDZtU4�K@PDt-m��4IDDO-PDSE�R�DECE-5�RU1-P�ADkMQ�DD��@P�� "����Rp��z�V���б\ήu	t8&�W�y�W��b;S.��u�����gq��T�lN���G�#$���C�0��j��Z_��3>��㔜���@�خ>w3�^G;�c�\efNt��S]��j3Z\���W���ѳq��o���w>��Zr���ϽĠsu\餷rc�����VH�߭��F/q����ף���1<=#v��~q���p}�4*���VC�3ڽ7P[��r ��񸌸1�x��D �{�a௷������[�77Y0'����^y(�2N
�fv�����}͟��������R�\ �;D˰jv��^w��>�μF�\]B��fS��cjf��q���ɪ�=����E�BcӒ󪴔W=�g�;&�*T�U5
�8�|��P�WOC�3����`���'�N�������i��
�AE��v<;}�Oh�Gd�t��뎛�e�M?W7��s���w1_r@Vж�]��?{h�͌����t�}���*��Yi�Y��j���s�	���/S#���}@��	wS���( ���#���~�~x�3�Ǿ��ۇ��V<��v��LϪ5���3|���ㇼ��{�S������GL��4�)æ�*+�ۻcY�\�-Q�L5���I��1�%zrt2������
W�u�\����I_��yg��TU#��Ϸ��3���s��$�9W�R�f:�e����ڊB�|@5�{�>�?o��۫��ю�r��V,��Z U���C�K���B����'e����=^�z�����r�;��S����β�n���^�X>�>���ܿ]dR����	o���<�B
#;�e��>���ɚ���o�'��Q���r��[�z���{��wsHrePϞ�:U}�<5�mL��Rʪɕ£�PG��g�1�-�-��:+�g���ϴܷ�Nn}��x=�AJ���e!wA�SY���zf��Z�\,��)����ɞ���3��[
��1i�Sq�����ꎐk��YW�*8�\.@�f�q=�����뙸�-xzZ�z�7�tPN�<�ۖ��nw�����>P���隞�~��<*�2Ѹ�3-�γS�;�̜�h��=P�U��:|>�+�_x�x�*�J�c�����u��}�>�uL���89�)�Ͻu3����D�C0U��]������R���C�H�U| ��2���2i���U�x����ǳcs������*8\��G6;]+�w����+F�9J���4�#��!���3*9�q7�<�͸Ĥ��q@�њ�	Xd��Ǖ�"�����o�!��Λ��qrr�Y6&��
E�^mf����ng1L=��oZ6d��"J�^U� �X�k����o���گdJ�qڸZ]\�j���Υô#���}w����:��+5z�ۗ����x��g�է�=�j���{�#��xu�>����R(���W�����3�>t;���`���Ѭl���K�w]6�K��:�=��ѽ�-���G�]�dׇ3�sq��̡�}Q���p�=��|4�m9�*��A}���vt�|8�3q��'�T��0�������5Z=��_�:L��z�Y¢<ϸ�m�wB��+�}e�k[��<�u33�ͱ7�N��r�����/g�;�Rr|����F:�zw0ss�ly��C��V��g�o�_��O�E�&m��3�����D.V�ϼ0�=����1�d0����Qĕ����=O�_�JA�i2�OMO�T�ۺLYW����������c�2��}*�f,ʎhr��3��~��^>�%1q��]����*o�V�+*[jtJ3����MZ~�V��w��v�|�F�v�ͳ�B�{j�M�eL�2�b��\�3���#]$R�
���\���B�J�O���G�y������^������y�8)�;a�tΏ������
2���{�ڵ�(�T���)u������}��)V�!��er����J�{����c��!G#��3L���v���d5|��j�No[�*Ki�ww����r(�\nv������}�7�����<s�U��2o���2����mwv��Kվ�M��lv��{)Ӟx��q٧�z(�ʃ����T"��A���Ïԯ7<�e֕lX�=��_�Q�}]���-��;�fj�S!NG<�ǌ/o�����]���'����z�T�.ժS���t�}�[=d���c���n�g�=w�f���'w�{����y�j{�q��ە�騼~�B���Ϥ����t��
�q��Ξ�_wG�U����<}�=��r��v��y=R�D��𨚇T7	7Y�1~��~�U��]a��k�������˙��ݘ�{!s�=S�Ϙ��3_7}fM���Y��d*��{+��� }��D��/�D��7z.���#˜�$xt{�Ϙ��Og��n9`�&�P����������0��e�ܩZ֭Ӏ���&#k���3Cޣô���w�&��<F�gǠ���[}>��f�&�����t3�^�g��hs'��y��&�*o�Fه����8"㟦�GU�ֽ'"bn�~�8�U����Wbs�w�a��3�b6����3'��M�]�����Q�vQ����:j=�&C����{j@rІ����Ob�t4Ο�nv}� ��M��;��1'�ݛ��g4-`��V��<Z��gYu�9(Np�E�2���򋬭t���>Ē��³W��]mbt��zA���ѩ.|��,.*5|\�S�n�/R��,��8�GB~�z0���X��`����7O�\g���.}oU�}��r}��}��==ތ��Ğh������ӟk��n;�T��rXY�q�5߲�`)��	�\3Ir�۵(ulw�u�ڎ�4�u=�ж����دӛ�A���3N�f��ӑH�f���ؤ�y�Ȩ�UѼs��eEW��9Z{�����nݵ�gVu��º�,��*�[�WS�ys�5<�[�^������+����+���wDo��ё�g¾}}q؇��s�=%�����ǤN��n����19�{��u>���2p[�&��
�ke��6eqЊbx�fvEI�����޻ϟ���7gn��C��S1^Bb\��˺��ݕs�e���x~u�t�O�/�2���Z��ٰX.�nw�{�0OT�ﻳ �E��q6�W1q�fWi����W׏�pd �{�&
ޓ�ގ����~F&�=U��^��M.z:T��|t̻�U2i�M���e�G�\�h��`�/ü4�qO��gʰ)側��Ɏ��1��vС_&fW���y���θ��]
@'X�Ev���O�O�V�� �@��5f�G)v{yU5#pu�wߟ��Z��F�=-��-܂����R�y�m!~wCՑx6ْhV�sz�M�t�떧=���w{�`���Z�ýn`�V���ތu�h$~�6�cŪ�KR����(M�>*Nh�I,��z8�@���R��SP��>�8(~W}=�S5��o���E����'߇�k+�s٪o<��tuMtuS�~=��= ��9�]q�h˨������^q�ד����l��9�z׻bH6׏��qfP��Y�x״t�ׅ���7��L#LL�Y�-�Gar�<J��=��Y��e�ST;��Y7U���=���g�b�~0ד[���\mt����ʍ�ePw��\l:�[�VBx��n�����|E��魛��CF�ǫ���u�9Q�r�>��q)�wS9��ǽ��r�]�E-y&�����L��*,g��\>n��r٥7ޣ-����CUW2b�Y_�z$���mw�<ow��g��]�B�T2�:Ulp]�d�͕(�����у)vzO��s��?�3��^�7�~��'���M�w�����|1�CE�U���m�}��3ko=Է����qڙ[�]~���x&n2��n#a_�Y<�|�S�;G�?m�Y��s�b���O��V�{���t;�ꎸ�-�D���O�kʙ�FYh����en�6x��F�,�ޏ^ �_�tw,;��/���H5���񧉱r��N-�ԃr��8m�W������z���*�ڻ� �y��b�7�xk�[�"�V�ua�a�h���X
�Qf�Hx�)��A��tf��Y�B���l�\�:v(z�k��������ڝvE��Y�߿���T���\<��2ٿ2���5>�����-����C��l�^���M"=ëan��j��gF�*v�[��	؞�q��3l�D�9��sq�1����}Q�~��{w=Fȍ���ܽ[A���׵<J��d\�2��,M[��&�*�Z(�_w�1��-Ⱦ�׬�L�}���*o�E�ؗ7\;�����'���u�S5��Ӽ��V<�}��~Gg�����ng���?���������ɓ���g�*>|eq��Ow<��Շ0��j�W��@��MK�>ګ��dx׼!�������S���:��*��> �Uo�C�	 v���q�V��?��۷0�6�X<.+��y�O[5�� ����y�w:�ǘ��}=�q��O�)�9�n;iIb�r�C�Ϲࣣ�z�W���3��{����F�24z%O;��aC�f��>���i��4۾��*99��z�C�'|.:JW�br�'��U\�>����%������d�1q�3�vD�z5�Jq3�v{��Ͻ����([���ק#�X9*}s8ӟ�k����P2��B*�jyc�7��3�)i�k���R����o�Δ����Zw�`����w�B)�Y�:�%*�o۾U�8	��>B�T��}M,c����˹Rr�y|��Y�&��'}�[�o�h�h�#����k%o�]��}�-6n-�(����-o�����O��'�y����k��5nNE�|���>p�G�Jŵ��U,h��]�w����S5��~o	L\F�v}W-��nj3��6��u�K�w�y�z�׼p=�
�eOq������T��蹗�UǢj/�.f��b�	r�ȍ���N�������^���Pz����7��fம�UYa�)�}T�S>��r���dM�|J��M<�3�i�z��xtQG��ʇqΒ����g����ݹ�����"=�(�[�������7������ԇ9�iC�W�K��:-�q�{��~�!x��O��m��Su��J�۵��(����s/.5����M�?�j�n�[���<�v�z�	�#�[����X��%��h,!���^K�R�.�?x��u'P��OnEz��k���4.1���oЏҼ
��W�
�q}�w�/T+,̮o2&j,�q7
!��B��֏��}��:����*���ȩ�K���ӛZ��1���W���d�3κ��Dp�A���T=�eqī���=��*�p�o��.�Q�0�K�G�-r�%���+B��ށ�j����
���q��J���ә��]O�>���I�ݾ��c���ݝ1����Lan�wk)�&b��gR%�팝�t�m"w�=KO<��bI�4u;B�p/*Չ�͎.��f*=�u�d��uGE�&fG
�s��ԟ}�hMW��������W����M�V����k"i!�g:��p��MG��;N㔋bg�z�����W޼��<t�s��T��zJ˽@z�:��]n�^�z���y�8=�3�7�̢�&��q���ox�:�x�gn�{��q�/{���ʞ����q~$Z��0~�D�*�����7/�?m9�?Bw]&����_O��
W�+�r���>��t'�,E��M-�x���`�������e;��.}oU�����=��=��%�׼7w�ʟGnҕ��SL�rXYW3Q�� ���:W^w����ߦsw4U2g��}�דp�a{"ݹ��_�>��,�ڙ�q��]�fpWl��U}g��˿M6��#�K�0g��l�w����h���-������7#Φ]���e�
��c��ocFok����y3a�&���7/a����z=��/��F�S#��z�ttw����z}<X��2��wS�;O�' [�'0��������\t%*���_���=�؎���5��Ʉ�d�������C�*�:ơl0����K[�t:-r�f8q�層2g&� 轥LR/�m���X�o:��e��%��>r�V�wQ��6dp3|�i�q�xƞ�r����]ko�*�<����k挕���qQ<��C�<����{�z��g�ד4�\�F���୮"]]��訿z;���Q;�=��
ٕr�L�Q<��g{�*g}x��@���a�[�̺N���ҏfrHߥ��b�2��*�W�v\�E��37�+��p�m��TE�X![}��j�����G�{/��+	��V��G\3�<�̞]S=s�S5���C��T����SmOf\z��v�'�X������95����s�
���"G�}ph���few��d	C�{�/c|��u�;����g��T�[�3��^�����t�GNF��q7���q��v��	g�{����]ߊY<f5<&�#8z���w����9��ׅ���7��P,L�oet�z�m�^�Y�_�S����RV�"�j��P��VM���&�y���{p�=��_���i����.��JdS��Q�.�膝f�̿hܿ�\�mK�4c=J|P��F;܃q���N�Y��`�a�5��V�q18�Dq=>���)��tzq���v���U(gY2��u��w�.>i��F*ݬ��*(ʍ@U;��M޾R��K��ƕ��cTL�) i՜#�u �sܻV��`��[֩ ��=�-ᫀ�N���2+��;V[�jK{;rچ�)�*��HDg�{�ӚAκ��MR�����p55����Q�Z��_r�w���������*&��qb��SBѬ)�F�W�dgB�-�N*wNK�X4`�vb�Mu�鱋5J��]Z�,䶇>%�ST�6s(Q{	��Em�C/l��;oe��OK�f�Ȑ&(�\;�9Z��$Z\�ie$a5��,�v�f�`�Z�As��8[�;�xUpQ*�j�,9E��-��.��{k�\f:�a�<�*���>�۽ƍ*����f�pWm#B�^K�9�'��+���Bs#j��ӧ|b�oRD��=l7�`�����=iYA�mbF�>9�2�N�
��zS�8���(���6�X�\�����ލ��3)��\�Bݏ*fgJ�h-�xJ�G��Ø��� ^�]�+�B�{.�ǈ� @�Fj�.pr�7)�N>f��$���+��r�4�|�u� ?>aCV����2�[�{�ut%���^o,}�_S֘9s����фw3�cd��X;(��E�q�BJ��V��9���.6y]dQ���h��TH*.�Qʆ�1�4b9��G�+�]��/]s�]]�r)�����S�eMT=�seC�r��N�b��w�]Ȼ
��̧�W8�@�u��λ��aN�μ��,;Me�ypi�2�!��*r��y�]'Y�aaSsb✻�i�޹���X�l��&wnT�:��h"��K1kT4�Qu��-j�mQ6�=��`r
�@�<m��&C�[���-2�	�M
�(5IgMFa��-��b�>8���#�F�vU뱼���%��e���:�ԕuJ�e݈�L)�-mZ���%f�4�Jߥ�8_g�M&�!\�@�ǧ{A�u֥���5|��T��;Wd�Cq)���8�4��8�F����M��=��+�W��,}��d�	�CZ�6��O9c�����<R%V��//������SC8W*��i���\�QD�H�k[i��E 3O	�ܼ��|0���jB�Q��,��O���Q霟�t��pч���M��{}b�^��oR��9t�s,�P�HN�s�_)�����f�������c���mDG��T��s\�)\��<L�5�54wg����3���\�S+��A�v+\�ewm�<�+�67�VYD^}+��m�B��
�f[��8-��u��A����3v�o���[yCC���N>�� H���Bn���#ыy�f�442�4]d;,I��G}��2�k����v�uf@�o���x�
���r���m��H��(3[��.���,G�g4bH��\��69Xԩ�+&���8�rv���EM�����
�sYun��*�΁o�x�$�k̜\x�HrJ�Q�O��Ve��.-M=K�4�+ݺ~�>��>�*���
h(���a��T�-%QTEPK@U$C@LEF��A��G!�s��6�Z �)�1@QCQSCsbJ�9�CE��a�����$AM�"�
b
i��C�18�$)�g�mb�4���ڊ
ӈ4b�� ��	H��PQ!0�Q���T,T�*��[�+Fe(��%&�����npvƩH�(�f���(
J*-�A��BfJ* ���h)
�H饨�bF��)(�Ѧ�i�����
M$�\���F�[	���lQD�Ӣ�1�l�����a*�l�5����
h�0DD�4�PV���墒�()�m�<��cSA�1����h�)h�4h�Hh���(����E%4DZ3U��T�f

98�B�m�catUP%U�RST%Q�t�k`16ˢ�B".lRu�����}믺���6p��ML��[Ձ��Y��ӑ2���f��`=ʻޙԸ�P�{2__`e�ܮ޸��:�t֢�Eo����"y����L�Ѡ�w�sHrePO	��j��ʇ�ݹ�Bj�-��T�^��1/_9��뽙��^q��sxKC�M�w���;�����Pi�^����1��U��F�
���pfe�~�~���x&o,��a\F�a4T���C]���Ƽz���S�z�eW��o�U�!N3XC��lT_U8��EQ���T��h���#+t9e��SQC������ٺ��⥼�u��{)�O�����l��L�zr:�O��]π���y;�s�s/�]��һ��Ϻ����8�F�w3���Fg��4y�����	��R;w��L���^K��s�uW��+�k� x*5�GY�R�Ȳ��U�vX���U�M�U2�WxO��!��in��ԢW��w�΍��ڼ��9�}>�szd�zz���uJ�tOTOmL����w�`E�񾱩MșfC���l��ۛ=�9:G���o�]>�h4��EC�+�yW�*�s�g�Pι��fJ��iw���g� L�&G#�Uw��xC�����vA�s��w]+bkS�Yg	�,��2.�2gv���]�T_���ן�[�x4�4/��h��g{�A�7t᎚��Ra�-��`�~y[�v�����P�c�
+齇���RIM�"��f��Y)	 ]��i�>#e�z&�]�QW��d\���&;�Q(�]�jJ�Å�c�<��oÅ��Z	���({��v�W�p�#�U�x>}4=�(��ϼ=��}�L�}�}~��1���rx\v�z���Փq�U���5훖�/�*���c/��z�4⎺�KC�}��B��fg!q�p�t��+����@k���%�����>��g���{�ꜻ�j�U�o�'�b��}�dOf��Q���g>����>��F��C��Ԝ�����o���K.� ��/����߱��g ���4�{mt��ɪro�t��k6����eiW�r	=~U:#{�*��Gg:��6��g�a)��	r�6�[��%_aDd�M��r��j��.WAT����p����d9��2&���{,�/�%�CqGfʔ{�7�H�a�mx�7�>�R�zV��������}A���QĹ���g<u�D��h�l��5�Vx�bRu+	�f5q�{}q�a~��������s�4�:�p�h_��[oٞ��������޻�7�x�J��׆�~�K{\k�_���|���f��T�R6��^�{�5Q�b�Zh�#Ζ����j~�~�xu>� �D��'7�5�w�`��t�g�{9���/3e�#[|ph��Ű[KE_�y��Ψ;��zm.��[|�l�	a��N5��o�QV�M6��T{�]͸��-��8#�g!;o]�:qv��p{*��)�l�*���T��G&:���s�L��7Cߎa���7�����M2�]N������Ӟǌ󓶡\����C��1g��^�>���������.r���x�N��@��R��oo^�^}9d!�wvdL��5�T9&�5��z���2^����9ƞ��%�;��s��<g�A�3!�=�{��Y�d�]7�T�}�c�\Bș�B��J��U�y��`�C�J��$p�ø���yW7�Q�K�pz	���w�^�Q�^̞��ї\�U�����ׇL��Ȅ13�Ǹ(�٫�Us\��T7G�ŏN�heΨIxO̞��ֿMg��Ou�ʞ+����a��̘�N�k�=�bn��9��Tx�r�̕>�vnmLx�%�3B:��џ3���[�������>� 3ڈ�y���_��ru*�Q��3S׷5��3��FtW���y^�+�/�5U����ф����@w��<3��iY�߆Ax����ܞ6%uέ>����ܩ�[4�v�,��9,,���&k�A��1��k*�`�a�΅[�B����V���+ �2}Ό���.=���\�Bhs��j��EӋ���v$�����'�S�2�޳�x�s�7�xr���S��Е{u�)={ǖ�*�T�vPÖ�2Z	o�t){}���rƥ�F�<%��\r՚�)��α��~V��^���k����0��[�=6{�o>ީa\rW3oS/M�"�z-Α���~��ʍ�,�:r�'�]$/�_qͳ޻X=/��_w�n���!���y�˱C�W�3�{b� s���t��=w��}���~�T�����7��[
��7.�Un����mF�xS���H��sā���o�S��ؿ������Q������n���<¸ͭ�d����qЎ{�.2%G U�r��Zv2���˙=߲*n;����<�ǌ/s�]��o����υ��}�z��#�J.S�7��{àx썾O:g��]�M��D�3ȿ�L��9��z��/�c�ӗ<�(��������`��(v>��K,���2��\ȫ}be^�nw���:�D�S���ͣ^�;���F�tB���`FDv}�(.+��WT�_�]L��+��Md��͙[��Y��g�m����[�����|;���s�
��֪��/*!���ϥ�L�5���wj�~�UO1���3�����V۝Ͻ^�?]b���+-:���ҿ	�!�A�����+�N��n���8��LU�ո��X(<��J���*m9.�W�fQ1f�s��EI��W:��R�=	--���;�������^����{��ZoԆq�W٫Wu����r�v�66��[���%��l Sc���mwI���[�]sذK/��^��k-Q�3ը�XJ���WC~̘����A��~i�=i�������o��	�br'��L���BQ7�|�S,��7+���Y7�5���8<���ꆣ���@g�ŷ���]<��y�Z�����gS3-
@�u�.��ےvv�8��Gc����{�}�H����f&�y^��H����^���ީ���`�m�O��}�}9����te��>��U����/��ٚ׳=S摾3/3.a>��R�%�����!ɕC!�|,�W���w���q.:���o;a���2�e�Ы)K=U�>�O�o�� hr�M�w�ݹɶ��oK�Pjt��^�`�o}j�M�֋�5�.��:P��U2�R�L�^��3q�Wx[
���	�����To��k���e{����v*�TϪ;��:s�r]���2��O{U�O�������e�n0��b&����Fj��Oy����:���莩��쾻�2�GZ;�-��Y�W{ٓ��(�"}�;R��!��_��ΣxU��;���/���6ộ�w�{,�[�dM����`�6��DE��l�	o�4����W�S\�֯��'���>�t<�?mܓUw3o{����V�/P�3u���'(�%P�j����X��Lӆ��[�e�fZ����7�!��.����	Rc٭<�E��¥�bs�#��� ����ˏ�*���إn����+/8_;�3]�ݿNd��`��TomG_��HO�����zD����zD�i��ں��ԞRC�S�ڻ�ߨ���V�Sq���Ȑ�T*��OR1p8��AG�z�k��p귣*,+�[QEڅv:dt'_���ϒo�~y��b������5�����3�]پ��51d��ݎ�S��Lgp�����u�~er��G_�Z~�������>.zqzݳ�N|���q5,�z;Ԉw�S��\��L�.�C�շ��P��U�	�{&�0�\k��0�{|����{�����O�ӓ��+�;����}�t���J�[Fr�7�HS�3 1x�U�j����sʯ�s>F�8�T'S&�7�N���k�4�3��z.A3,n7��[��Т��7�lG�o�?Uq"֯�`��R�/z\k���L�2籗�*<��m15���ֲ��9�m����F:x��.0�A�/n6�ni5NN��>ʪ
.;�=��;���X���{";����U1p���]�f��?7��.#	r�6�[f��<;"�6c{�&d2t��4�̐��u�� �p�t2/M����aKg��s�9����c�2U�@�F�MT�[����G��n�Lc}G*a�ށ(M{�z���FuN��;([�Qa�$��/k���Z�;���T�+��ݺ��VP+k�Ŧ]KZ}���v;��a�q��4ͺ.e�q蚾칛�)��;���,̨�\���gP�et�e!�:w����쎮���URø�2پ%L�7O�7ˮxU��B�g��_d��1��W}�#y�P�u$.<�c=�}5�n���}\C�-��R�+��\
�o��f�3���D�wǝ�s>�l)7�������#�[3�w�����ڣ���lӗk��n��X�C�f�q�K܏]����&�i���=Q�[=�F.<4�5xU`<r�O����]�{��T��ِj���@��/q��R��o琌��"f�;��.m/W�7�.f��di��A^Vo�rW��灌2t�!�*��"f�g��T9�j�_�z��̯^é�ȃ� ��;�Τ�l�Ղ;eK2==�v�B�3+�ધ�d�2+�}bn�wC��O`G2��r�ncIr�#���:#�@�BB�]ӝD���3�;��;U�}�5�pzR7����>����7���o��~�ϼr�o�pW��;]qց�&n=Ǹ_�v�zk�*�c����L�MY�w��%%�\Fo�$��z��D�$g�Oa��<����-�i��l��v6:q&�^�%���Z��id5�H�F����>�s��S�J�V�94�EA�Ƴp=ëJ�9�`�/d���@�Lb釩�p����ZA�k���wxD�ӕ���\��6��ҧw��.
�_V۟dz��;������q���W��N|;8������=���\糎�a�[������:;$��gY�Ng�Ӿö/����ў��3>��m��ݡ����2�I�N�����~�e�?zih2e=�-��.0�p����o&;j��^㘯�=첷"�z0�	s��Og5nNE���ێz}d���ۛG ���3ﱿdmK|=�U=��c�SY+Hヸ�/�}��w��j��E�s��~���.�2Zf���[9ck{3c�\:��̈́�������dM�l�`,>�a��]���zG#�,���M�a=ם.ǇC6�#U�+rzd1�Ϸ���T+����p6�˨�U�#�K�^fg����gd�k���=W������]=��<�@u�zF2R]f	��qݬX8�a�v�u���6����+�����F��2߫��O���r�댻�ٸ=޼�Z�=�{d���g=�km���<S�n�e�]��鋉��S���&ev����U��k����d7[_���Y}jrΥ�2�Y��d�
/��8�0Ղ@#����6����X� Q�Zʛ9on���Gz�0�{������y��.��D���Y"���F����P�YJQ�7k
��������mGG��[���1:W���}cpV�=5Ɛ��K2�L��}�3_[�M��FXC��\�����mz�]�c�n	�}w߿N#���- <ȇ�A���euL�39�s��z-���U�}�������i�
x����ޯO(���ǧ�����FD4 ����=<���L�E���]����2������cF����*���?�67��>.gOTt�br��#`F4�z(��/����j}V�ٓ׀��px�l5������1���a�o��SW(����vV��N�c�|��q�f��P|*p�w*ɸ����<g���׷�U����/x�u\s�+�����YS3�T�\o���5��������~��rW������t�a���¤՗��]Q�-�\xtJb�I����S'��`�;��0�c�����ޣ-��gL*�g'|��-���r7��&j1�d�	�1a<���Xw�y7�O&U��|.
�q�g*�w�V�.U�;�SC�tk��B�������3W��' �p��f����-���)mnk䥂�/?FM{s9���}7��˵^�֝L�)�D|�)0wz>8e���1�{&K��#Y\�Ƿ�3^䑖�M��Zy��p�b��I�Wv*4�$��II�5vw�S2�,W:)kZ�|
N�ky&��N_�t������6�z��|pv���\<��#r;�����ۧ� uS_��>���R�{ǥ{Փ�gxX���=|cs�H�{���V��z s�p�q����!΋�Q�"Z/�%������5�L�2�@�B��A�~*U_�hqU��%wu���gtZgg�{�g��N�g���8�2ٸ�3:��Y��o�\����c}�U��)G���{��V�P���Y=/���S�dO3<:V]�5��rc�}ԙ�K�㟅���u�_�2G!�2 x7��i�R�Ȳ��WuГ]��_�XV0c�N��Sc�D�R7���~9������b,_��9���2��ai�ŋ��������W���q����z�f��H��Ry 	R��׺;#�'H����z�k���4�ש��VEi�T�>�|�id�+���3���SݟKˉ��`Q�\G#�Uw���?Y��Y�Ϭ��&4\�+8�j(�l���ɽuA	�x;~�}w;Aة>��3w�����]~���2W����z���z?������+��.��s����3%S��D�	����r�B�;�Y7�Q���2��W��٢��@�x��K���_oJp���k;����֨k^>���J�\��w��:��r�����N[�����C�R�	�Lk�β�4b���p��=�S�ĖSuj�&lb"_>Rr�JNhs0j�pV��7��1��r��u��Y�Nw;M�[��hr/+(>8
w�e�$�����:�����.s_eAz��	Hѻ�d���]�]�;S�WS�EIn���1_Z}�a٣��q�L��b��en�]e��1����ٽbJ�����.�8�����cC\p�v�d��6����x�uvQm%��_�;�Y]ˀ�1�!�䘔�D�B�׸|E�%QHp�-!��	ڰ;u��t4�ۣX;�g>G���G%���ƴ�T�C���8��v3C&����n.o!���@ʲ����u0:�"U6���gdA(T�8�9v��� �l�N�i4#�p��p�A��wf��fZv�jg�� �&_P�.m�b�����jn��Ճ�&�n�$ۍ�w
�ڇ�
��ջ}��Z/e������s���O(��w=�S�^ʽ����G��N	�͎51�m��n���>�/+��.Q�-�ΉA&�fnZp�mt�&��eЇ��9�[�.���<][UP�5s�\���s4��b^��CFJ�y����J�I�|Ҽ�r�l��e%4��7L��ND-T�h.��&b����l�wa�˥��x�:�}�)	���*/"�#��cZ�;��w[ȕ�����QWr��w��5Y|���h@�:߯�D�Q�h�.*pm����g�-�Y�v>+MZ3f-�ebɫUi=���ť5*7m��U}���w.@� ��"�&h�Em�$t�y+�+����M�Go�p/��CJ���rL6x�����Z���uN��^(���w�&
����K���+�u�̽]��"M��S�L��6�g�o��Ş���r�Z@@��YF���ukZOb��л�t��NՊ�]M#i;�1a��H�"2��ڛ�E�9��p�%q���Ca&��ۏ+n���ۭ|�bĠ��yq�<��r*;�ڒ��5�ULޙt�>�$��i��/uw���r_��[�@��V�-b��&���+D��}}b
�>���)ؑ�D���9����3�鮋7���K�'�:l� P��<Rjݲv������d7�B�� f�{��Sx�[f���-��3�՜V��o���=.d3j�؝B=�e:��*��i/SR2.u����W��TB�_-�hޡK�]͗Dϛ1�W0Q����tq�a����"�MKy����)��*rô �94��)Œ�m��r�*�m�om>1���q��	y:qw����m�	�:w:���]�R�QL%U@P�QE*ETU1TQCQ�E&��U��@6��b��*i�4LAH��CTQ��
.*(��h*�
(+I���C�8ER�R��0�M$C3G6�+A��)b�-b�lR�J��@V�HQEISIi�jɠ�
((�� ����"�ZB��B��AZ
�LE!QIAAMSHQAMiӠ�ѷ9��%i�ST�ZLQSI[aփ��bH���%�91h4�h]�4$HDRQCm�C���Jb��@X���SBPQLM4���Ѫ��@\Ê��9�i"R&��)654DU:CZ֒�*��b�:JR$���tPŠ�Hld���&9��u��߿�w��}�����Gw� >8���hp��|����ư�{E�����v��~��QN�zk�X�w���>uk�ۜ�c1�%�?������������'��u2qug	��xf�s��Ϸ)w�0��S�<%�{anU�f������z[�W�1��}O�ǘ�g�'�k����ͻ=�gw=V����**�^��Ko�WF��(tw��ld�zBȎ����3xO��9�I����M��+���\߹֦�s��v��o��7��m�ػC"��3L�V��%��bX�U7��t���^��}�i�����])��}.�s���9��*�"j���j��p�T��ݯ3�Σ<pw��gѶ\�e �Y�[�>����I�(�H���Ne3�s�|�:��i�`*�����^���V�k'c6��nT5�!��9�A��v[�9���1���*0�l�d�cǯ=�Zê�D�B�����v��ld[���g�>��W��T+>���8v���3<����̰v� �3�ΐ
n�����@�~���ڋ�NL�+l�=�vx(�3;�����������[btNw�=���}��6��&Q��p��������<�Cь�����`��h~UG�f?�V��7�9��/�}2\ז;��W�u�!dqW*}[�Pc+^�8��@tki����f�%���R�V"�,����!�릴_>�邥f�n�j�#��Zt� ����u��m�ngu
��S����q����F����	es�0�B��7�/6�IC�~������2'�S�o3�ĢG#��Wp�vx�G�s�ޯjw�X��yY�����O���Ѵ��Q�%�B�(Wό��
�{�@yS<����A������cW���*�����Tx? k��B��(��>3#������M�����2k��b���&�#㯱�y��n��q|��|������Nˉ�����?u�U����fB��~�!~�H��O(��@S���q���;#�&�.<���Ƈ2U;��=�bb�Nt�]��E�����u�+l��{�����Ϗ�����gU��Md �e����+oW�q�-{���s3ܻ/d��W�r78�{�P���M=�~���_�������@?�;,��m��޻^�P7ʋ���u���MS���甧l>PT��%�,䠸�\�u�̫.(���?�+Z�YY��h���LdF���n����4q����)W���A��fK����EJ��;�>՞�+��c��wOEx�f�]��0�f����oζ��|����-����F&_Q�)�=C�=��V*��x�}�\S:8F��>��>�m��7_��˫�jw�����G*'�]�p�]�ˋ���)h�-�e�;��e>���Y�7�ws����٧�U���e���%V��.�u,�v��W$�7O3�YMvU�zޤ%m��������	���1b48P�k��b���{���uߦo��oa\{Փݐ�!���NܮI��#;�m9���힚�~����t�%�uX����~��������-����^��Sr���{��j�n�=
{�A�fz�;-�T�up�~����G��}7�ד��C��A�\l��M=���P�Us�;ϫ���[L��H�a�L��&+��"o�g��3���g9ƧܰL��Gک^{̡���g�&
�rzix��g�����e_v\�[��3j�0��z:�Z2�kލ����wѷS>Y�G�?џ@B�0�z�.3'��3�v\�eڻ��3랧�=�D�W=�>�9��Gxx�ק��9�׋�}.{Ъj|�b���O��=�.�̟w���Z��ꝅfg����e��yUm����W�;#�'����z���k�:N�}��U �TX�TV�����9Ƨj�j�b��x��c����x��,
<�N���~y2��sgv�R����3O�[3-�G_ݵ����ɾy�{�p��[pp\g^�wt�=+�g�qNM�WSc�wiw�-_V�m�L����°������Sn+��D<ܖ)]g<@�T��˜�{��T6Y���f�__Q]^S��R��C#���Xz:����)���������HY~��h���6���Y��L����u���]�jq䝟\:�s���=S�������W�����Y �����I���T��2�.�N1�>�9��2�ݞ�|p!u����ŋՙ�W�:��BȎ�ɚ���o	�1�reh2��]�B�T1�|��Y���dR����|���p�f�]�������FA��a-��r��9�_��l�<}������&��UV�����Z��C���讱l��{���5{O��e�����x�3dӣ�&�ov?4=ޚ��w:siusG�ou��N|�K�y�e�q�T�y{�94u���E���b��K���*���};�wGJ��t_ɝ�~����u=ǅCQ�e��&S�\l
ĝ�����-����ə�g+b=Q�*/v�����X����d~��;�y�"���ub4��]%v�����\7�fs���9�/��������(W�>��̧P�$�`�wJ����'mB8L���&���Bٺ��۩����߈��g�n}!�T*��Zz��E�C+@�E{/�@+N�y�L�S���3^]G�5:em��U��n4D�]�a����n�k����y�˲���i��*U�D�����v��|�`��=���7xr�.��s8jQ=�pN��o�W3'+���A�XA�&/�q��s-s�e���k\ˈ$ơ{Bf�L�SG�C�������ިt����/-��멚���Ry�����W^���"���z�k��ۣ:�g{`����3Xk*���uO�.4Jf�5ò%eD�� ���r;�U]�{>�xC��Wh�K�٣�][�oB
����t禕�)�D�P�\G\wUO�c9W<�'˨}qշ�n_g-N��N%��u|ⲷ�{����t���z��H�R.O��W���VO;�ȭ�a����붚�Oو��Z�kܴ~_�U��^?]��~��o{�r~\o����N����5�Ď�\�����-SyK� '�?P��t�]T&��/�'�b��3>f��^��?b���>�)O��s����lvno޸y���<,��zBλ�˰gф���y�K���>m�Qʹi�f�y��fyMOBj�M�S|C�Q��P��튦-��λ��E�~o�%1�o}���9S���TI�Y�>���\n}�ih{m����[�C�uCQ�K4Yٖ��2'��&=��`
����ׄ&�e��=
ϴ^���=.�]$5�C�=��f�=}}8��1�Le���:h�i��(I�@��eZYb~+�5�Gx�ːJ�����u�b��͡g�j�`�37E=���Sݜ�IJˮ+��}�0��>�H!�#b�J�`�
�N�N��U-F��#�x�	�G��i�-:v�k~9���>�2�N9��ț�6���*3r��˩!>G0�Ov_[�f��9EϽ��g�Z�
��*�d>��� w\G]T���Nd�aI�=��ٻPǏhS�Fb��5�c�&��(!�s.Hm�辪���_x�R�=w3��NL�+o�!�n����S~��Vf4��y��y��i�᪐G#��q�����*%����<�U3�j�١x�N�gj~=vjk��W<y����%�<�}�4���+��Q�q�"H���Q4��#pMTy�ǯH�����g1]X�9�-VQ����\m)�ҩ=4�����Ws�<;*f��Q�]�`�K�&3w;��33��ѱ����垈�~�y��*<;�|Qr�#�}����OOl����κ�ɨ�]�����������"�iN��d�ǎW���a�纣�E�3����]�nfW���͕SN9��y<������_���/�?����y��i��~��'���ΰ�/�U!15��OBt�b����O�X�~�J���h>^$Z��z:s�v����3�zۉ����2�Wd9K�Tˣ�#�z�Pc��z�����d��+�Yh�,u�P�Vz��9���\��z;5۠��uq��c�
��9���R,5�"�8w�.��آ[Թ$��슌��A��Ci��>3tp�wwl!�&�wB=
~4l��w8I�GWLɏs�rs�{��ܫ%�o{
p�駣!�V��Q��ܲs}?{��)�����?�'��s����#2��6�����W5��&��xvs��S��f��튦,��´�=l���}�񦗞��f\>�����.0�+�i.^�S��0��,xg��W���TY�W�U&���s�qb̾�k��2��WLշ�a���-�Ƚʆ�+����������_�_u��/e:���\�:�xmǺ�]��e�3�:��7�C��al+�s�q	�B=z�)��O��v����uah�	Ө|���s��[*�^��wS냴�2p[�'0�V����o�t�^ũUR�s�肩��΄W����W6��\<�<Ǆ/�뺟H�ʹ�ێ�z���n��F�37'���D����N�sp|y�����L��fA���1q7⹏2�ǳ�x�o���8��n�^�ݻ�82 l{�c�o���(Tiu�F��fU>˙�]Fe�|��`.�Z��}���>�nV��39�#=�T`~� ��I��A�̮uL��Y�4%�������M�.��Q6�QeJ�o�����vk֒:Iy��w�Sd(���x��]*�Y�����O#u�܋D�"�e���!:��"t�rP���9�<h��w]�1��q��U6b�ő�ީ^��'�:�.㮂
o�j��{��ȏ�k�ρ>�<��~�G��|���{�wz�`���[&�L��K_�����;����g�O��vA�s5��O��]�Q����,��S�q�TOx����k­w�&.9x
����;Qپ5�sｆ�����=��O��ď!�ɳ�]2~�U�3oL�%��voVO�g϶�m����L���B�<j�=���k��̸ҽ�suUѝ��Ǚ�󸍮��Tk�������w�ߵ[��+�r��z ��+���㌸�>~D�,V��U��Ɲ�&�1���'��z%0��'���g؝&}G�O�遼�&������*TU⩞��o��{��$+����}�� �ф����	��h2���sHrePP���tOM�~{q���tayc��q���Dv��1n����+�L��?	�H9���K��	���E-{s]�>�5=�����{E�yTr�8CQ�z���e5U�&��9Ap7��@>���7�����!w�C�*V��o���uuá����e�qĨ��q;n��T��oh���_㫗�"�/��QɑSH	G=ɾ�z`Һ�dr��y�v��X���A���1�K&/���7$'U%}V2�>Y'.�ԕ�4aM�n���$��x\����؎%�	��ʷ��ΔW9ih��y�����m-��l.c`�2��)M6xLo}Y��L��g���XwC�������Ow��g8�wXjZ �k��G�/#���?g���^���5:;��}����|*/�P����}#n���y�b^t�wB��\orƔ�>���X�dOC���"���z~.Ұv6PC_�Q���R�23��VҿI�q��֗��ze?���յv�Fe�_���3�n�7���Ȑ�*MC,=c�q��O��^������7���멚�u�Lک<����]{���'H���i�y�������;H��4MGU����S��$s �\A��;�k����O�3����F�[�����g �ޮ�5
�n!���������}�ʹ�^d�˨|��#,om{umip�q�z�=�J��NfL*��D�	���nk�GY�ܫ%��f�~ܷ�&���y�����ߩ*�/��<���WVxXz�����)�'��!"��R�w�s�^�X�c:����/��'ta�9>YUӕ���'�c�N3��מt%�������t�Q����g}Č��]9�j�ͬt�pQ�jg�\?]�5��Lk��v��4n:T�w�9)b�v�R�<4�Y�*^AC�58���Pb��x1%�����;�#`[��\���-V��gBy�mi��9��O����5��}'X*����sBO?���U~�8������ʿ'*#<n0�1xO ��e*�| ��~�K�ƸJ�T�硢��S�|p�+���aY�L\:8�9�~��^'�Yp�mvmٻ��璴�8;�R�MKak79�Z_<�=g����#�w��S+�G���w�2rhW	�X�w��*'��.g(w��^�t������}5z���i�8e�3:3�+�7Yѧګ}����O�V���5>��2&���o6���C�]I�<�c#�tM:�!%���=�^�H\������b�zN���U>���ND�
N��n#7j���)���o�D�$�����+߼����N �:�I�uL�9�=������Ϫ��ӓ�-����C���>w�GA�-�yBJ�|(�X�6z%������J��.8�S�*dݻ�+�����U]	Y�G?���ԧ�vr�}L����F��<m��.�����~�Q4�k�Y5P���mmC�w��V�ⴼǳ<w]U����:#ü^ӟMGʤ��\E
��eu�T��<���}fO������X�k���ҋ0 �7�٣N�FkGu7�D;ۂE]{�R����:m�S6��;�iȣU�T�K�#oME±��`���fr�
A%�ƕ�p�hNU�-�U��2`s����j��T���I�m�})����@Q���c�;9����[]�q���eg����YW��	D�.�^j�5��z�n˩tF��0�t9g&$Q_�]�`��H5v�F�^9K�v6��b[���8������o�Z.���PfTرV-�W��Obǲ#�ĬkM��x�K.��a{O�eÃ���R���笆�[�K��I�� �n\+5��K��r��W�ϙ�v��m�FiĤB f2�"�jV�
T����+$~�;e��w��tBf����E.�k�$%u[�xQɇ���p�n�"�5Bo���qG˶�I"ul�S�(`z+��e�:�9aTn���l^��#+���k45Ju�r��:6�N��C2�]��h;HU�I�n�������q�r�J�W\���8n�}���tH��q�����mq����ƚ��Ŵ��l�>z{��H�njNĻ疴g-\c/rtn���Cu�ʣv`�'p;5�%Q��gG�>�(l��ڦku)5�ӝ�<|��v�A�mZ��fLu����DfZ�o�����܇9"fl�Q�3�J�Pu�a�S�庖�-�V�����B,���Щ�þR� f���ao,r��7x��m��K��޳�>M����uf
.���wD�mu�_<������!C}r�Z��ZNJz"�z.*�;��1>�e�nw^A�dp2*�i�_I�.ỻPeU�S�*Y]5I`v�S�r���ن6��u�$�NRj��04�{i}���#�u�4�˃(���E���l�$��*Wp�y �l�v;�+.t���v�������ju�3�a-�wf\-P,uwo��t�K��YW\+3xہ�D���V�>jΪ�L]Ծ��n�M�O�����'#�f�8r���R�sqщ̦6��."c��5ڝ���I0�ܨ&�)�]Kp�l��EɨH�C�=i,oe�+�qb��������u�؎Y5���	N���e��@�k!ǵ/e��C@;���7����YOw"�03Ի��M�v�k�����`��w���I��Qs���0�����sOَ�6�*�������͚�ψ��3��n��t�6�8'l����;������*�j�ܸ��@e/��}�B��n��P޷���־�ڲ�0Nc�a^*Q*�'X�vcwصM]mF��]���u	�}�ecxj�ĺ3����ۼ���Qe#j�5gn�Ŏ>5|��-%l��yDa������A󐷕�������F�*�yp��Ӱ ��Ye�֚�qVԕ��H�H�J��qWtx�64�
<K^�]f`i0s��p�*Gc�ٻ����c�Z�i<�2�ұ��
��#Q6�}�K����2�%w�=�4��WF��Gj9�Ȼ�������
�C�*�6�:b+�6T�t�
*CC�����UD1�MAN�!1A�uG1�Ѥ�i�������"�93�a�8��-�U��Д5PQAG#� ��(������������)�X9�C��ht��S�
b
�*���p����T<�HPkT	��KT�Rr�m����Z4r9�A�C�y<��hI�j9)�����`�J���Q�M4�hnF.l�W!tri4��(A��C��"��t3H
4����A�ѧ�hN@EG--9��DrW���1r��4�����*�i75��󯻟{�����j��n�]�ShM`�[5��)�:�4�ٴ�9�K-��f=\�W:ͫ�;� 8>o�u���D���*◝5V;O��w���jw�Į�e2+���P�T+�s��æf�v��5��q�*=�e��j��,��=	�73(w�>=+`�d�Õ���<	�3��;8�������?r�˽�[��C�E�ڪ�5}޼��YD������շ��U{Gdx�ׅǙ�q�s=3��Z�n�k���x�,��n�x�y�����3�w��uO�~����q�;�{����������n-F��\�.���z��̔�M��v��β}��?d��8f�UƎ�1y-E;��}��z�ٞ���_��e="\��ץI���޾�:�)��!����S�U��b�*��=��v6�?atz��Fr�A����=+�i.]ƺ�\��OOD�~��O�����U����;qz����N�'S4�8әzr)L�_<ț�i���e�9f�v�_��J����>��V�j��m��s�ܩ�f��,���;�O�U�:�L�:N����T�񭨟j�w`ܥ��(�X]�Gwmv���g¾�C+�s>��^*�^�]��ix.f�Rr�MG�&���B?
�{��jL�hs���ɞ<s@�e
�����n�K�ǈZ�#����1 �7ۓ�w\�R����ouf	x����fj�X�B��u�V1���@�;9�w]B�5����š���N;u��M�m�Z.ŕQu��:fŞ��ܞ�+���x�gW�33ݔ�*'��5���c���.�vB��nV8�rμ]Z}�=��=����%˭;�����,q�n�e���ϭ���2���*Yʥ��/�R��pc�y�Ã>�;���oI鯗�!ct��Lʮ�s>����+�/3˷���8�M��2���W+��3}W�X�h�v=
��� �\fW2�>㧫���s�Y3����}�)m]
o�&�X��+��{�vN���'���q��<��UB���lkɸh3�A+��}=�3=�I`��#�u[�s�^����7��9+�H�quC�lk�]H�9��}����_/S<n;�O��w�&/�^���('_����pz�k�;~u=VME{z���$������s��iL���&j7��f��#���}C�Ͼ��=��86��FM�f�P��%�.�Z����J���ϻOL�{�u2c��p9�=������>�6{�]��_w/G�]�wW�qU��G:Ȝ��{�n#	��q)��=�S&)�q��I����{'� U�²U͙�H\ڻ���k����z�9%e+Q�N�*#��z�Yҙ���v�
��/$�ի^%Tk2 l�p�+��a7��vX��팁�z��칆�NVܛZ$�f�[ܰѷ�tb�Q��P�g���o`W�Wϭv�������/���o"�O�,뼙����o	�1xO&vD����ɾآp'�)�����]��3T9q�,�Q����8<�ڙ�-�S�rߦj����a��sE���X�y�Wzw�\��>�Z=�q��Tv��F�wEu��]L��W����	���djfc�9��N��5〡�0ܤ:*j�v��ϨO�����Q�0��Om1�EO�yu>����~nnx����`�r��n�7��<�g'�-�M�W�i�ṕ	���G�٦��xt�|�/��S�;�̜�h����E��;�[}B�zF�f���ȶ�}]g�__z��4��	�7Z�3<�:�Ͻu3����ӑ5�����mG�Q��B��d.�͜{�I�:'���t�3��vX��U�HFe��n��m���^;�7��gb\��>����}��^K��OA�GLv��,��ؗ�s,�"g��4P�T�ev��g�N�)ލ�j���fn�Ej����;]]>�F�R������5=��g�s�(��9lUY������?;*y�o"��n'�pQ.�n��kH�!GbV��ցU�/f@�1���c�B���wFa�כBD��.�)-	�IJ��P�(��2��|��;��`�b�Ti�+:^�h������Ȭ��N�	���y��w[�JXC�y�vnq�Ӎ{�~��3yl�^�=*���Ȑ����P���>��7RBzu�g�;JUVu�F��y�x�}5����ٮM�~�=�L5S}w}���!�&�m9<;l�����K��̍��g#��z�E�a�^�h�\g^�vx�x߃���'ԝL�\o�����{�-.c ���N����,�M.�����G���U�ʌuz��1q�g�������&�9�oX���]�'�,&]�y��q���P�~>�;H[�br���f�1�|���_}#6���b��&{n6���j����s��\m���(B�J.��#f������5�u|�<j���{��'P���)���b��nk;i��yNxuR��G��7��gi�	fM�s�^v9L�8=q�6��ϲ��a.Z�z]ƺHjg�덧>��<��M�ȶ�}yS��z|Xň�b��[7�T�Z>�g*��7m�7�F��ʇ.���=�>��oX�k՗������c��~w��ϣ��q#�̶,zJcs��}puߧ2$[
M��st��׵�յ��68ja��PP3oE��ݎU}8]�ڄ�uZ�����wk�����`�5Ij^��O�g0�1��=Tn+)+~)wY����v<���u�y�M���[�!(@6a�:Fs��{U��>l�i��J�q�UVzN(Sx�� ��ϯDWy$I%��J��~�	 ���OϽu�V�
r8��/�
��빟_ud��[���<�P\8���$�o5T��F�L�@�F*<4�g�_z�S<��T���;=����}���<�k@d��>H�uh��W��J���K��X4�ieq�(�ʿ�fD�[���^Aq����k=W�;�ו��q��!�fW�����s�U%�j�/���
�{�@YS/���ә�/3��,t���TV)��d�G]�5:�}�W�p�=��Tx? j=P�R��7�¡���`ݱ����b�O�%�\�L���Umt�D���N�x9�M}��N��#��m���D��]�f�{X��u%O���}�������m��>�W�vG�Mxy��)S�p}Cy��A\���]q5�i�Z_���ʏ���8"��ktd3��>wbr�:�GN�'8*��RF�����t���U���g���*f{��.�`i�d�j��(x枌���z�ۢ*��Nh�
�.Ǔ�J�����Y��}���fS�%�{��M'~w]���nT���;u����3��@T���4N�.�H#����w+������/Nz��g���Tp?"�Ngl"<	�ԮL|��5������9JɵfG�5�R��S��aIG�͊5����;���R�֚W�'¥�/�b9�O�O�
���6����.�w�8�l���G��b�=-������ɚ���n0��=+�F���뼛��a{"�㞝�n�l73u�V,��kN��M�>a�L��ٔ��ɞ�~Ȝ���[�f�v�\{���Y}��yd��ԅ`�E�꾾�,�=�y�˱����wS�:��7���7���<f�\2�g��x��q��HD�mw��8wgd?M�GL���������U�i�d���ŝ ��{��8�-�W'�OD3�u�ml��=�epЊ���췑Sq�\.xA�< )~���Q<i��u���c�WmM����xY���}#���;�͟b��l��C�/�@�}]��"}0�LbгҾ�q5���JU�v��L��T���}P#ƭ� >�D�x+zOMB�.=,�=3+��!\���V�/=��7��X:dr}bf�Pa\�s�7�u3��{��v��a���(<2�o�)f�>��B��P��_K���~<A�y`�7�c��{=�9��? FK�UO�폚���Sy���{W�T���"F��B�WOg��k�]��'���V����z�=�yX�i����y���6��e����R�NDuU�����R���9Â��49Ձ���է��n�Y�ن�<�����bʞLQ���p3�6�M���>�*�]A�3D�7)&�5 ��{�:iYve��/��1�/V\�k��g(XV,�b�M_K�ٸ��`�ߟ�'k��#=Q5�Ǎ�q��Z�fL_.�mPhgTv;���}۱<�{���+����Xk����m9��13[�]3ki�������ɸ��2��.��6p�"����t�l�A��׷��V.=�g�mt��Y��N��Ȇ{��oVK"��oػ;�+n�x�mX�~Sb{'�O��u׳��P��c��7���ǃ�Lh9�ީ��L'�:�u��<3ܵ{�pv�;S��h!q�Pa�u��w�8�\��=I��[4¶m��f���n���:�{�Ҩgл�x[�Q���X�#��i��eU\ʋ�~xm2#��oȜ��\t����n[��Ro��t{���Tu�#R�m�Eu��UL�ȥ~��cˎ4c�\vN[��j���Bg��h7��Wny��R��Cs�S>������cҽV=�#8Ioap�>�1�ٷl���s����u>�<�s7�Z���y[���ޤ�C<�����R���Qc���%�j�D�عEm�Ŗ�}�>ew�P3�ݗr�h���T>���1��l@����8V��o��������60��J}|ue�Eo�(�O܂������Ӧ6��L!w��d��3c���-ǭN����w+5�Oj���1W���h�V��x<-oU�{z����뿳�n�p�e���P��M�Q��xoEL�������f��Q�����jfh�N|�We��Yݺl��1�����_Uqp�O7�1�멟_udߢE�-�@y��׵�~��=��gp�k��©M�=�H�|fUC�6��$32�p��=ѷS;Qx��T�c=�`�z_2�5"꯭*欑ɆdG�����!�ힺ�뀙�Ry�&���z����dyVw������������������3��2����ۉ����4��Gv�K��;`��	I���m�e�s.��Wh� �ާ=5򻮛D�&�~�#�����\�H��4�{}�t�^!�=ʀG�շ����z������Fә��}}9 g	�^V�z��)��[q����Ʒ��X;�Փq��tx32�l:�3�շ�N�����'ԝL�&��Oss�ڬ;��j&�dz[�ӝC;����3���z.@�?V+}�tYt��q���\y��/����¸��(�=�>���;;o��P��:����Ǌ��H��^�!�b���[E��>��H��Ħ;>�g�OMO�5NMӮ|r�܎�,튦�/=��a���κ�n��UŇ�*oK�ކ����a��Կ�ٷ\r	X���]�E�},�0�W����x6T�TO�]w�T�˺X�)t��s�p��@Z�7{x�w��f���0Ŗ����h�`<��Ч�u�m���q�|�t�f ��e�9/�s��_��7��0+�jZY����SC}�T�
�=<�O\0���=�l�w�9��l���+���ԩL�*'�O����e1�9h-���5�B�Y�[��s�9c��d��tMcW]�c<n�Bڠ�Ͳe��[7ĩ��)�\y�7�]>�6��nT;]I	[q��n�0�qoy�{E ۃ������x�q�je��coC]d�M0��=ȼ�7~�~�7��t�F�ļ�~�6���tWKE��.1���;�fk�uL�< s
<`�{����}}���U^��Bb��-�}����=�vx(ı�ǡ��.㽙����3jB��E)�{��D٨]YԽl/mf�ޙ����Y�b/F��:r��:ix�8�����&i_
��%詓^��I��4��9�	�y�z���=��:�>�s�R\��(Wό��
�{�����\_��P� �æG'�&�{,�$T�x�W�p��\EG���P�R��(�U��c�>Q{�Pn3ϱ7�5� ��U^��쫛��d�.���ʭ��Õ���Õ����W�g��z3������FLҫ�ꙴ8��5 {���fSp\�.nk�eE����+�\Bށ�]Δ���0��RI�:�R�Č���.u���Iղ�8΂�=�޷3o	��!dlL�v���Gh��h=�R��+o�}��x�e�wHɊ@*��9Y�~CT���NE˞�t�G�5ܯ'��F�gGV�O������+�?kn*���o��)?�V�t�p�]D�iy�&���9��7��q�5�	��a݉��gg�$�W셎<{�Jn����xz����;��=��i�Ʉ�Jg���o�����M=_?W+uuN/ޯ)�J��z6�
Ʋ���O���2���eϷz�v.K��w<�;3�_r��������)"{gu(�9,,�������d�TճҸdi.]뫚��0�߻zk��T=�&�ۙ~K|'�&�/�s�hp]�d�әzs�g�5���D����ᗹP�ҝܜ!��P�s�z��wv�hw�o�����V��[<v�?0=����͡y�-��%FC��߂�Ķ�L{Е�n�T�mu���7<��B��ё�3�]��Hݫ��n�߉��r��6�x���j��^3�g�_�I��/��ͭ�gk�S���=�pf�W��xA���2�Л�	\��C��~�w둋޷��e{�����4(3�<�9�������}�|+��DW���+�UDW(*"��AQ�eDW�*
���TE������AQ����+��
���
��PTE~"
����*"��AQ�UDW��_𠨊����+�AQ���
�2�ͭ�`���������>�����+�t���IJD"T�J�I%UR�}��H�UT*��(���R����>�*J�E ��)T�AB��TJ���"^ �[fAY�M�m�5�1�����wt�.�(\ p�ͦB� [�: �ƕ@�{�Me��)kRR�a�V�pwZ�F�6�:�۠6��sn�Gv ��5M �a@�	@�� 9� .�P9ڀ30:.w(��Q�s3�;`� ��� n� �(݀�w.hh�傁�p�@V��ED�p�ڶؔ��%T��m��4[2���mjةJ�@pĺ���MXXT��-hiUBSl���P \�;H���k5��­���U��Ej�J�K�6�m��ViZ�f؅�T�֤��0�&��l� c�ٵU�Y����Tlh�l��m�(m�'z� @ "c!�)E@�� # !� O$�� 4     ����*4 #F��4ɠ 5O��JUT�S �     D�Bh�4h	�F�h&OQ���56ԂM$��U51Hm�� M2`F8r�ˏ*J�P�-�*��kg�[c<���*oUT��(�;�8���P: U*�Ĉ���S��?6~g�C��f�v@cn���
@�ހ
���j�$FA-E1�юzk{�g����m�
�*eA�mJV���R'�e.�F�I۟QM;��|R۹�V�+_+c,��{B����RӐцżo�jbwxZ:ֱ�x&śAʟYд3s@�����&'J��V����
����kb�:X��iE��e4�&[0�syʪ�.���&��ⱌ��⸴�wt��VK�ô��G��z�q��@��J��+e��J:��RK�����:h�ۚ�އ���˩p��<@G##&l�ڔ&h������c�t���5l�����)���A����4��.�y�n�v:��:��n���S9���cP���%c�MbЌ@
�N�]����@�7Hf����.�&�����k)iH���Q(�3a$�;CU�^���ۭ�^+�Yn�sB�*�F+��=� ݣcS5r��Uw7<Zf�w�A�)�7n�vDl-S�HO^�Wt�T�dٗOtR�NJ�o3)��k��(�]pr���9*
�l`��G ���-���ڣ�m��fx�]˭Ւ�C:�hz-M���Օ�3��֊j�ʁ���&P�rY�����._��QZ�ә�BƄY��@+mQ��H�1��Z�`�Bj�A�^�(���ht?���2�ʄ�n�U[���m:��4T(��Ccͷ�XuYUuvii�	{Gkpʙ"Tq�^�`�A�:�`�+�&m&����TõgI�w
���T�e�O	h�N+n��Al��H��3E�Rx����.��zH{��Ug�r�Eڤr����V--��m��]���&ܗr�����NbUX��B�hda}���8ۓT
l��[$�K!Q5u��T�*�2^�d�?g��[�% �'q��ٌ�7�)�i��p��[�Ȱn�9��6�-X6½ne4B�W��m��x.�h���0�s,L����wJB�V���i6����L9*^ո�J�T�Jݠm�FPL�j��]�kō�(�ͣ4۬�m	(�mZ�I[���ᢚS~�yv	���*�+J�������Ν�᠖�,cM���K�`e�sZ��,,��蜬İ���X�i�"2T+)Ĳn���X�U������tBiɎ��avJ��2�TyH��X�-hl	�6��W��P�Y0Ġ5y������z�ęu�c�py��lU�i+��cte�'�p l軭��'B�#YW��y��]R�SE�%^�9�qk��)��X�(kaF\������Nh�Ch��;������H�dա���R�{T�CY��y)�F�PޠM7�p}eØN��E��I��j,�g0�H)�`u4� 6r�Ji&K:��۷vVgP��ӽx��T.	��*.�(��1U@����2)ج��ٝ��C�P&��w��@�]:vN���=ݙDV����
Y���1�w�u�V�mj���f�[V�ޤ��#uin�,)�C�q]ĩ��J�n���75Jt��S�pS�͚��1Z���?�5�z���ۙsWա���^��b(`�A���E���
�"CF�1ڑ�^ݛr<h��.��-ڴ�Ťg٦�����gmڰU1����Q��)���4�u��h�j�
;2<�j��{V1<[ٗ�ǈ];����L�sLsZ٠n,���",��K���]^`�@ǵV]���m[�@'M�\W��2��f���5��d�[B�hU����8쉰���@�n�fb��S��r]Ì�1*:�; ϖ�Y]4f6���Ѻ:nnPy�@M�������deU��ZY)�:�IT{�:�[�wYS�(�d��c����� �cV����4J ��
8��q�9�M�zh�2"�_m0Su�ʸ��6^�OX5j�ipSsD9��)H@GB���؝k6���nM�9��P��D�b�t�Wu�� aV���IڨW/j8Y��"n�Ɏ���[�>=�am�k�(!L����pH�`��FmE�Zme��U=����Ն��#h��-�:Je���$f�C>�T��ɖ��,�����j���b�9AP���*l-�V��*wV�Q�Q��3VQ�YN��:2[e؎�BZ���Ͱʱ�PIj3i
�yd�In
��v*��T����dzsK7��D�}�F��5{���B�m#4TD"��������M�6�sE�Kf `ZХY�c�`�h�8�-�kB��^^�BRۤ5jd�:�4��f�Ӳ�]1�b?
Ǹ@���y�`ư+X�a�u�x�t^깉�Z1����1��1��+
�5b���;��6��	kL�N�wA�3	�]��e�w��v�B��f���fm�
8K�O� �!;�Alml���f3�M�4�MZ�1Q��=�ܗ����� �)b�Tq��7�E��#)��ph�y��hxT�phw��".a�ǌ޴aљm�a��
���~U�L���jpYV���{�����6X0�oYԞl���Su&�e\	�H��IȦ�bI��w(YJ(b�Sdu��el����!��"��W6��t�K����q�{F��Jڶ���4�M��ț([5r�3Yv ����6�����MZ�[��;�:֍�p�`�L�p;ܶ̓0�!��X��PT¥!dS���ωBWL���5���z�B�K@�V�Nћ�'��?�������n������H�����)���D�W�/��l`���D��0�.R'v��K�ₗ5�-��-�݆�{'m0�L]g{��E_.����i<,�'��1ݛ�;07ڱ�S���X��u�`��o �Ia��Mh��0�l�Fq4	�:W,�;�4 ��y��TkT�jO��j잫��>�Pպx�/�÷�.�T'�`h��^�p��7��t]��}q�;��wJ�9/%�0vC4���p`cx��7k)�f<ζd�1em�,ʙӝ���\:VUT��5�<-�*&�"�����+��ChE��g�oC]i��O4�0lՅ*�\.�w�b�k
R�py��W���{3E��S��$]r�I�/*�)h�1p5��O��i;�K��ʫ�j����hͧu�ZV��}�J���k��l�ӥU^�6�wtX|`]�r)ʺ�pmd��V���	��B�4�g;�j	ۖ+:<�S(�[l򲲺��cr����g�yl������v�O��c�*VS4Y�/z��$���ڳx��R���'	b+۽-�������ӝ��8/����Cyq�����#9�y��B��Ks�cPc�:]'��z��n����;oV�&�4t���VU��{xHDf.x]\�Ů���{�_5G��ç�B�h;Nn�����&�a���kTT����Q�e)P'F�snV�.��0�`Q�36�gz%#��RI��y!7�D��c�4]�,�%.�4t����uh�-���Y
�����9��g|h�Wr�b�������f��#P���O�N�pM��r�u��R�+��32-Ϲ��&JN<�aծ������R:�G��u�=�g'j�NgK�Z�c/
�d�N횭�r�:��/g�M��O�B��V�l��އʠ�����^��r��=d���;,v R�c�7�z��e3P�t����jС�W����s��(�Q�Uz��قB�a%q��,ފ�pJw��@Q�w��s��y�F�x�n��9�0�-$j:c�kZ�YϥĦ���B���:�o�m�-;1�lVh�3h��{p���DK&l��'	�3
BQ�Rc2����z�V0E�.5�+�\��moN�r�����|���e��z莩�RJ��R��-}���K`�r:�;N����뺇�X�dk:r׵�vft*�O�%u��#f��d�>79qB��-�q��<*�|����#���6��+�4��.w�24�`۩�"�3wD�ԁ�[k@��(`��C�3��]��m�7L56it��2���|�OV�(���]�uXu^`eqmug5���g���y����	�K��N��ф�������_!k�^�&�Ka}87�w��d��걲vN%w%��Qޔ\:s�5�SReczpʐ�&��uiĮ�c�V�=۳�mFK���,�¨��I��V�qem�:
@��8���:�Ѣְ�y��c_M&b�|�����;��Ǜ��;�׌,U�Vfj	��͇�	����wV=Ka�I������9��p����r�ߋ�p��t��z�l�k-d��N���c��/�J��	�L'�=܁U�E(�(�w�i�e���[i)�3Z�n{f����܂�����U���+�ő̰��]>}h܏�z�[�L�d{����#ٵw,�9f�ܾQ�㜌غ�__Yp�[�N���u�Q���{��8�q��9�w
)�4䐬=�01$o��kz�\�tɩ�w�GL�N�tWf�1�.�9g_>�+���dGd��#�v��6^����.'j��4�H�-Ԝ�֧��tF����E�sh�jYי��S{Ky%fw0Ȫ���'�E�Ҹ)n_`G�f�wL3N�,.�2>jӻ�9��K��O�
OcY�"�=ӧ[�^ ̭P3t\!��tz*��w��g�޺X�Գ�,��N�2��N�u'�ur��T6mu-�g���m7H��w��$X�H�8E5Ciѥۨ��k�V��!yj!wrn�����wln�_�!�������]vQ��F�fPILd�ep�
��I�״��w �9
�婮�}	��߻��Cb�9����R�m��F�Y$�� ��@�Y��j�<2Tt��_�r�]�jʛ{:��_m�^���>��b��Cz¹VS]b]�$��S7�j�}�^
�x�j�l�,Rz���#]�7:	��jS�ew[Z�$�iN�.0�6L��h.��MY�D�j��kV��ߕ-��#�{��"g4��J�,"}�@�oKW�6���*ZgIXo��*\�`f�n��-�b�g�m��ǵuk,���֏��P5�vY��`�Y�!�>�	PV��-h��.��u�r��v`��z���F!kF�pMz�*>��N>W.�	yd����m[�-�>]����H��9��{�$.�Љ�z��3K;/�e����2��Y�k̛ǵ���fہ�JR�NY�,>.Nu�[���ػ���t��}�J�;����ے�}3 �
�+y����x�GdP��
���}tv�iNs�SyJ_}�Ĝ��zge��Xqok��N�m��]�w�^=4U�i�J��͖-"�;	�k��X�����wV�΄��0wb��{�2�m�n�=� �V0E�F9��R���aJYF�*C#!\`����j�0�D��˃"򂀢��!����TU5���#�gTEN���f�z-:.o�r��7�3���MXUmW$2�o]P�M��Ь�r6�wjm�Ue�W-#7�tY�ve��Ct�Z
T��W*dg�kz��9N��.³HU�[�mR��8��ol��Lak�FYL�+[Xw�51S�*ݡ�S۬oZȬ��A@lp=���n��}��4��N��X��0Mwϴ&3�7m�W{�v�b���dۅD�a�,,"�%��n��
����6���׻��}��u�|�Z��,/��ݾöo�X��dE���F��I�PǝS����U���yQ�F5�w�'5Ǌ�
�2�rl�B";E�-G�
��a�
�ӕ���w�d�p�ۂ�*.�
ufsyt��yŖ`���fsZ�7a^$��3(��K;\��e����
U��?�֧mrW%,�;iWMtm��l�>k�sY�s�j)����u�bK��ogLѽ��e����P�u�3��}��"��jU�*��tT(�M�Qb��v�ʃ,���u��Ĺ�ಪ�a�t���s�^5�p̏�ѕ��'t6���t:�ʜ�Z[w��<m-A.���+y��/]4j_1d(��#p	C3f7YϘ��R���8�+��L%�p�/cjg}3�o׹J��O��C������wh#�BԾ�KvH�]�X}�d�Vj
}�m0� 6i���j�wM`ӡ|�9�^��Ox����j�wе�����5F(t�'UY��s�`�`�&+9V��n��|���mb��)�і�,�߹��vC�b# {/��.�F��8{�1dc�&�,��{)�<��8s��쵝��3����h�4�tpբ{;���sP�k�ja��5�In�7�Q��@����ܔ2Xg�;������Ur��asku��,Τ����9��7��K��W�J�$胥�e:�8����jt�0h52�ơP�"��ImZ� �w�M�[Y��݃-T�e+[�1w�f�;6.Z�k�xK�1��)�8������H��-��٢�^�-Ə1}��C�WU$��+Ky�f�,O����Q�v�

�$s�@��W��}5)���n��q��{I��S��VcD�<5Pv7V��~z{2��Cf�p̘�Ma=�2$�N��7����r��.b�+�V�����9��V�fW}}{,^�8J�1l���S���;Fw7ZDj���Pߥ �S�Ȝ�˶L�bӽ�|ۡ�F�T��x`��r��
�oU���-��I=�N;�Ҹ�:J��r��fN���ݑ-�j�Y��dNP�%��6p%��7A�Ebr���7n��PC���}�<��'Ɔ����CI��DùPe^��ռq��9g�^�R=YH>��� X��a�F�r]����ѽ/G��H��<B��at)��6��tA�P������V�6l�h�n��PΕ�4�]��f�l�ve�Qdv�G�;���B�#;�J���3"&�Cc8���~�2�>{\�w���E�׽!�昘6�D���SŮ��w��K.��du_�KE�a%���4��6m�Uu(�Z�M���!��C�e�ղ��ڋ�|E�Qf��묹Cbָ֓�t�uGnV�.��P����U��`�h�O��Mrנ��TWko��J�n�C-��0����#iyqޝg��M���7&�0�*-���)3Fށ\���h=��#e�W�����7�kw/�j��U�ŕ����
p�i�ء�5�3��.%��N��>{Gj^��sk9���X�<I��8�O(��m�4��#�BB���vP:;���ٛ���G��=s(W.)?�$2+�n��� ]N��M�\f�9[
�F���V�a٠�Lֳ3�c!�T�<:���Hn	���a.��v�k^��AQ�0Wd���܎���O�B���M�QK쾐i�v/�?]<�ܰ�Q��X��vu��L�/���ui����p�v*�7��bc�[�ۊ�*��AV�A�[#M��5p&�Я�bj��I��񮮇��\_dF�DN�u+���l�3��F4z;�{���/���»��y�T�緡�d*�+��5��/lQUˀ;����T ɋE=x8���=��Ú�W]�2aRj"�BePWUեk+�<��K����+v�iGj�Ԧ�]����Kw\{!�l�i�:R��[�
�1*/C�fVJk���Kn�^�nZ�cU:���K�C�h�A�PS%m���*ʹ#E|�+�p�"�vJ���yS��W�e"ıKk���t,�b���#�R�έ0R��CJ��'�[vdl�"�w.2�;���*z�1hY��PV�#&lL0Խ%}�	�\&hՀn2Λբugk�q����ͷ�a�m�f�{;��o��:`�+:v��9�l�]	�wz�t0��P��q�Q���3��I����}�����V���6m�ؙ�#�+C�i�=���K���n(�&�%��e
�x�`��r���WQ�㧩k�_V�M��q�7����wMbSg�Zm�9�N�};�Ô�^;�:�tl�O!��!&�-5f��p�&�J�%�֢�ה�NnÛ�!oH�~��gdr�Kˋu�vj��*�Ҳ�92��|i���tUV*��G���	���GgM&��EDT�	O��L�6Y6����U���.:����\ou��6I�ᶦ�r�u}�1*�wM��\�h~�OTT�uh�[�]���9���U$�pXrj\9v/�b�8��f���f���ccA�c���u���Ծ;����?ۡ�.N�S7�7r��Gt�MJ;aj�s�6�ɦ�!���AS�2�hR�ֲY�X��9���	6'�)g+y�-4���mg_l�۹�����x����B@~lNuN��<��h�ta���ٛu����(p1t�Iv�)��Wd����X�3b�1��D꼍����#9�1&ٕ����h`k�������r���������4��x1 �GŲV�) ��311�c��qQp��Q[��9(�ZY��(���\4R�31ј�ס�-+�TU�F(-Ŏ.Q�:��U��-�-��n$�2�*����u��&�:�.
&��M��pS%uLr�-�Ҭ�r�.��]kgYMj�ԥ�]%�F�3Lҫ4��3]a����Օ���+�J�-���n�[[��Km�R���u����5k�\�e¢�����]k0�`�qsH��T���nb�nbY�kEO!���|�ﹾ��������:���"�;����#|��K{������(�й�>���a��*am2jи���We�[���UZ��Ho!o�����!s\^�R�q��X�I��d�u�;�쓛�C�m_�嘕��O��b@��}�u���m�����`Z���U')/�YN�9}[f�w!���"󇋫��~=٘E���4�0/<�G�v�)�Sh����m�����нM�����.�ev�׭sP��Q���vϠu)���
q��iZ�MF�nKϗ��A��շJ|UEO�6vWF��Τ�U�K��w{$��-j�1n�P��i������#��"��-�Qz��ZH��Q�8�,�{��j����e�c�YxH��i�b���osy��u�
4��q��rԡ>����f盩��J�MeҌ�t��"���2vp�Kμw8'�d��Ns�XpLs:�>H��He ��.p����rn�wY������~/�cnx.�ʠ��}��w�ކ�k;8;���S�igA�x�r���3�������c}+��mdt����rzriI��X�ޗB׼���vY/H������
���t.]cu���������\���l.[�U�Q�]}�6:{��}CwS��lkb7q�yˠ%���&c�s��Q�_S������
�"�5?�+�ʇV0
�5��e+�9���ݍr�W����fB���w�޴P1u!���!�k)����aSci�|;���o��µ�Bߩ�v%p��[�x��ƻ�:�.z4������k�q�*���޿Vؖя���Y^�<�y��+^�5[��e)���J�&���d��Y�����滛\����T��X�E�	g�̣n��B��۰�XiW-4�MCe�=�eGw��4}o7�{��8�X�	����ׂ��J�7N��<�C�nS��!�U��Cљ�6�n�´Έ�Bi�j�َ��Q�മ�<�&�̓ה=|�h�z\MW-�WS.�.x��7�e�Hw!u��i�Qn\c>ވ��4�P�U����D����cB���>1wt�[�b�ՙ�����̄���Bnw=�-�R��5q���]n��&�ݱ�wt&��K[�.�ZC���aCچ:�ۨ���\t��;i#�u0ثo��E�UV�+����{ ;��v�v=���Tm_,�t�qZo1褳
�m�c}}��u����n��z����9%؏s�/vQ��;���y�]�:�J���������ڦN3�V%�l�K���:W*z�ĭ�%'��.��VE:mp�|�1!7j�����d�`l����}.��ő��d����8�i]ٞz�#�NN�jm.�s��멿;݌�:Y�p�E�p���$_<lnŏ�����e�����C��^x�.u�^$�;ٛx��^F1�o{}�]�/-�wܫM��4����C|����b�h�-Z���IFI��j�jem-��<�9�܍a�v8 ��
��������l��O�0�fy�l��u;�,��b2�a݄�fOg(;�l��8��!0ZRj1QA��� �3��H{uf�@��np��2缞h����7�<ng��F]�n�Ruc|J@&�pɵ�����!�҂�W�7M�!\��3s��Qz_�R���֙��'�k�� }z���e�y�w��#fq}ӷ�<��t���z1D��8�ڭ�㞺�Y�%���t ��N�}���y��Y��R��[բ=�ܚ�Q�/v��@a��đ���&ĈaT̻{3Jsx�SѮdӕty�`c�na�̈��pN������[��hą�T���>Y~������%y��m�a�pE�x2jT�X���R��Z����0�!�	�击�L�ހ<�O5
H�ս���ZJ����fULX�Z2�-�G����<w��q��HcBy�z=5W���'#2ףG�v��p��v�Uz5)A{��ׯb�Rnk׋�����������t�����
��Z�{U6�h\,�S�SS	��m�j1g3�N�5�*��2z�Z{K���s}z~�w�'�ß��G��]�k��}�����Rxtq�Z��]��q�wΒ����	Wf�h��]���V����<a��G�6���R7���Nmg\�=� U����-��ۍ�4�ur�S���vs�9�x�9���3­���5��
#6:B�r��@�n�'jrcͺw�����W�ש�>7Vw*��9���uׯxu�2D:YC��f���^�{r�!���dM�S��j*��]А�Â����z�.�
��
�Ywk R,��G�;KC��yZ�:�4����D�0�jA5[A���U٫�>�+��酂@/�gb`�v3Tm9�r+˄Po:$�U��wW��f��̩hX�j3r��mRG Ceӥ��Kp�zQ��{��*�b�	��U>�L^0��L�3	�#Ug5UI����r�&2���UEo���cX4.��zm�Е1m[+t���]%N:�,�Ni�;M�����m]��)�t
���h�ef
�S�41Zb�EyiHI��9�̶���g�mfD�#˷yxBi]3Q�"��iZ���������i���d$m���[9����}iE�T�3;j���Z��Z�Lu��N�-����У�Y��уKEJ���L\[�k2�V�Ն`��\���\��0L-F#-�\�F 8�V����aU�.	UWIF�e���ئZ#A�Օ�Ӭ���rܥj�5.SYb�Ri,r��Ʃ����]&$X�*�I�W1�Ƞ�cY5u���Db*E�:���z��������}U�6g��dub=�IO#V�������9f�j�Q��� Դ[����j��%P�ۥEu��Ϧz�J�����S�mN������n��Ϝ�N��)��/"���ǘg��$�A��`o�"ν���G����{���qvX���e��hq�]��ޯjeb���2;%P��o�"��Y�n�cs�6��lcG2ɮ���v�b>���̄�R��{��7-5�Z���W�{�T�~��j��5���`�o]�����d����`��IO���ix@��i�<���S;6!�9~��~7P��ݾ&�|���_UM\VHt��Р0���%(F��T�,]�g�Ψ��v�,��Umt[���,鸐�2��:u`vf"oH<jU�2]�ǽ�wfK�Л���[����t`ʏ���*��k�`\K�\g�S�3vqk�����R��Ȑ9��z�5"a3da�k��Ӟ��\�]��t�BՁ�O5��	8�d2z�W�$7�}�w�s��Q���UL�6�kX���ֆ &߭��	1
����'I']����5������ z�q�a���=@=WB�US8��76Q4�^-���̦g5޺<8����;a�E���	���8��M��հ6�{�����$� c	�H(��L���d6�i=Ha�H^o����������;C�����,	4���!�&��B��C��C�C/��W<��:Cn�o OP��l���$+l!�	:dSL!�Q t�~��|~�;��
�7��C,�`q��!�+xl�Ҋ�ր�Z�V�d�!�'>z���W�(w̘N��\7 ���Z٪�bK\�g�;���=2�9^�uwR��0<@ԉ�հ�p�8�'��Tä!��`v�d>d;�4�Кd3�a!��N2Caߺ���{���<�8�&�v��CiY ���ע�E*�A� T�)���� �N�=��|���IP+	4�z!�'H��5��:�� ��!6vy�ϻ��������4[$1v��$��;`v�m:d��� $�g��4�}6k���g�*^!x�-ⵋ�H{l4�1'�C�VkT�������s������>d�!�:B? t�u���]�!m�'�&$�`}����;�������@����͡Ձ�I�)=Ht�C$�c hϼ߽vHd���z��Мd6�<a�T!�9�hC��%@4��b�����~�VC�$��	*s���$�2(u� �'���=a�$�޻�o/���ē�d4��H9P3�X� ���Ή��d(����W��Y9Ot��u�VB�iO�Mԧ&.���������f���q����~�ټ�q��7i��t���Μ�t��Hw�$:݁�H| 0i��*�/����y�����[�ChCC�Hs�x�H�R��Har
��[Fejc+cx!��A&0<Bz�>C�t�`^Sl!��I�!�RH]R|�{��o�xI��Hks���#x��3��)��T�4�*I��s�oϼ��Hx�ڭ �l��A�(\3�bb)�@���n�i!�$:��p޳��͒�a
�x��FhC��I�BqI:Bm��x�߷ogٿ��^�
��P2|�dP�l��v��I8�@;d�P�@ߞy����w��q>`z�wI3��$�@4��V��"쉔�)h&"��L�4�^k�n��^���0P'�H^!�z8Z�����&Ǌ���\[���o�u�����I����VT�R����s����>���y�f���ނSR��.��b�]��/rv�m0���g!��ы'�C�SF���ra�1Qy=�!{�ᵮ�g�0���jo�\��z����'�}=J�m�-5wƼ�"ǈ2[�h��j�;=0v5<���n��7�[o��bڐ�/-h�>.���{�j�Du�M�ԋ~YEu�NӮ���3]��������ȗ�;���J���t
#n^i!�<�WIew;��<�#-�,3�d�î�K8<�CW/�#�M7`_�����~\*ǥ�6�ޣ��qy�����[�k�����mb���V����]"	�4�� ǅ�O!����jl�H�ճ�����C&��c4/F��4sf��呶���^UQ��Ӧ8���"c�s6k�ua>}��|Y��l��Ϧ��7�Q��}���q?'�f����a/�e]�p�=�8u˟1����LըAU�Pꝳջ�'$ŀ�(ҁwOߪ���{�5��:�0>��gd(�m&�M�A.,O[��+���c����t�|�9���{k^0��(úͩ�s����٬�p�F� gE�u���eU	z�̼w.P����e�Rl�=�7obV�����=���ۼY#�;[Pnunz�+2Þ02;���h�`>S!�U��v,
�x�ƍ��oֹ	�`���J�uIyݹ]�t��QA��X�hC�W����խ9�!l�랽\bf�����(�f��[��ˈW�ͽ�%3V囧��N�|Y���ڷ���-�W�#��I�L�n�dv��[~Y{����ݡY7��\��Z����SX�*ͨ�>����9ǽ��v����=�~��6���VcWm����qMcW�-����y
8�����)h�|h�'�,NK����+G��<5�@չ��=�m^~n*��0�uq���c��O�h�2���JC1�c��n��Ϭ@Zj�UpY�"wgivm�Y��qR*�P5O��}W�ر�.��š�l��C�ZLTc��UV��3�QO������o<$+��w����H�v2��.��3�F�l�f�u�}�P�W		��#f�2�-c)�s�q45�LgS\��k��CS=��d5;LC`���Y�ac��wT�To5�4��X7*�;*�F���P+�2���)aJ��Wp��Y����ObѤ_s��Y'w[j:��`�;+��سB��;HI�V���t�hV'�������O���j6�r�WU��4F*���i��Yd	t�r��GC�����U��sT���*..vRj1�mDL.�p����#��2���^.×�`���;tk�]�/�%�Tx����p��n�\��j������c�B���q��$m�vrʧ�QF�!x]�/��wV����X��Il]Q��3���H��,E�	Z�):m\fT����Z�X�T��T�c���fCr�
<���A�?�[B�n�x��s�R�!���C�j�da�Q	ʺ$$P���ZYB�Xm�Ï*��0�%uD��Ñ�ɥ	3��h$#%�V�mVR������<.�&S�fʔ��*3Q��H5�G�
�*� kk���wO)�9�iЯI,�@�^R�����Xpi`9Y��!�?|�B"ǉx��p�EZ����TL���j"
�QE�H���b��p�Tf�r�eTDFh��UEEm*�ņZb*��Ƣ#��mV���cKj��*1V�*X��Z��UV""+1EQX-J"�(��6�(�a�EQ�V[TE-��F)�E�Q��TE�XĶ�lZ�	B�����{�:6�V��[��,{
2��mF�śĭ��""=�o�1e�����*N����=^ؼ��U�4�>Iw��r�-u��1%�P���).�z��Ȱ�Z���^���<|{b�r��E�{Ҕd��9���Ǯ�N+X}_�y��J�^e�V.g��GV�Z�blj�e���.a��;4`�^��|�C��p��aeF�J�˾����K�z���-�����zn�,�9Q(q̒�Sꇶ�Fe��z�6��j=�$�ie��C8�YϬ:�SI���j^j5Tm��Qn,�wa��r�k�����{�^��t�C֎�F�wy:�ޏGZ��GwaH�T�;�I4j��̠6��v��혔�5� ���xGV��=W�+��8�&ݰ�¢�Gk�9�3��A�u�9�a��Vs��6&/����.I�36�=�_�����43�qr�O�{�.��Y�u�o�Rf�r�3Tn%������W��D{Ѽ�^�_1��μ9�!O�w#�9i���kk��c��h}��J|<�e��a�l�cWƐ��a�
n��gC��l�D.�,����Qam:;�d�ǖ��*И�"�9�H�J,��p�����B�#������:h�䇱Gt�ΒL�f YB��ЄB)�=V>�|��O���g��'OOSZ�'L���st���K=�zy��q֫������xΩ��7�^�+����h���6흾���O1+e��5؟�v4�Lgv�޻����ɖ�*�J9"���^�3�5��#n7.3�rѽ������|�9?����!dT���9�����.U�h#Uq���x{�;Ǧz&��i�/iۼ�u�h�a��-0����(�j�zг���;Cj��y��<�n� wS�fh(ٍ}�+�i��U����
G�{��hH���㔀���-��5W^�3��|���҇9���{ST����+ь��8h��g�����\���b���ڕ�5ax�C+(U�ڬ��[̿Y�w���Q�R�L!��0����c}:��	�p�p�~���!��E�p��i1u��pqY��D��΀U�塟u{g}�:w�.��=�xHA-�ZZ�q��}4N���u�� �����=5��k��&��.r��B�0�!��p}༏��^��ψ3��qβP� E�NLd�l��1�!�)�px��a�k�7��Wo�n	ܾs���y��{M>&w��n�2���z͎�}���S<���6|�����CuQ�5�~�ϻ#�;9�
X>(@���҇|�/x[N����?�$|t�p��Ɉx�6�ν�͵ء�_@k�x���!$x���5����˥��XtD+Uo;?Qj�Ԃ��<�z��MR�������Z������Yix�D�z�Ap5�-��:j�(����]��*`w�B6�����8�?�Bs�{�l��wO^������|O�t��^��"�1!�0�䅜u
FTd�[���=j�6�{v�NP�u�~k!�dBwz5�>��F��|����#Z�F��8���9!�!���MU���<����[R�W��?q���F<�F_;4Ci�,�[K6���|9fj�OSCǏj�n�ͯwo9s9�yq�G7�lӧ��/bc��Q���}-�Ƣ���6Q��"y�v���_�ń���v�0!� !"F�/�Y�ΰr�m���v%�u����'|���C���j��*�9q�0ያ��G/���z!�sv��;"jt������5X?a|LmG��>��>���g�u�=_o���םU��x���0�C)f(|Y��.��h�������"4��C��B�a�!�g}}[�r_b�T_���(�,�4,�8E0W
��ٝ��!t��0ߕ�HSC�����;w��ޭ��/��q��Z�]�3�Ɛ���C�~�0���CЅHxf�}D;Tp�������j
[!q:E�Qdf��l��|~Ćyq����xç���a{Nz���A.�M�t��'1�*��.%v��oj7\��k]Bqee_i�Dh�=SU��.+YJ�����W�a;h��kT-R�'�Y�z#ވ�=�=�F}O_!��w�ä�j��|�>��u�뺲h�E؅yag����!��E�����n��Ά�_/��hq8��׈�dY�K8n�X�愐��"W�$��!��l��������6�^C
HNB���'�I��ƹ^/Ֆ��`�Da$C�@�C�}gbY����~訏8B��r�/��5)��z=~T�fx���q�DCD����?g�t��Ln.>?.���ɝ��*f)�W����M��l��qj��Մ3�ᯱ	�0R=�}�&�ׇ1.`�̄L� ����MX�[�~�{ވ�fkG����LdB�}/��Qh� ��+8�X�؆E���v|p�/T����]��X�������헾�7jϠo�y�A�*��������e��_n��[^��>he�6s�+�ƈ�9������B��H�aߺ��'�:m�OM��٪,� F���	�<t�Ō=R��slWy���s�"���O�D���?bF�ٽ��Yqx(� "r���T~�Y^}��v{	�\D�w��� Q�C�����o�|�Jយ�8&b���܂���W�x��������*���'�f�GurU=�}�D6�iڟ�FR�~����<F$�R��;�r��#�e.4}��� ��Ф!${󬐳�O��^_+��d=V5B�eZ��+��@�e���T�+6F����;&u��aO�}	T)�E�T:ㆢ���~hW���k�1}�f$(�0��Y���}�15ٳ��;|G��/���!���d6�ҽ��(�B�y�`��g�U��XF��T��jJ��Y�� 3DjC}�a �0�7E�����8��C���p��D/|����F2k-��ޜ3+�^QS�1_oGW �>ͺ�K5��Ϟ������]7�8I��٢�10`����D���jN�̢
̶k�v�������G���w]%����ݏ��ks�o_cYz��De�n��un*�����԰Z�nr��N7�l���� T���B� 	`��]��)[��9Ri5�lI�ˣ;S䘙L��If��w����*7�p�f��7 x���
��Ƿ��n#���nU�����a�]6�r���Գ�
�i���o5@IՌ�l����[A�Q6Z}��G��'w�l�YB��W���Rf�[_kT�Ŧ��w��U���G��a�C��#LR��37#7�f8�X�2(�mV�N�&��TR��k1��h^�T*�ƥ�H�r�XE�˙V<��Z����2�3�C�e�bISxdCX2�A$f����e�j��zSE��YK.��#p�MHE��BP���d\&�7l��L�y������:ϱ��n^_��$�I��J�**���%`�����[j-������E)j
�[h�,N8���m�PZ
(��m��h�m�+Zֵ[h%-���%kEF��J�Qj(��)F�j*��-mX�"1QDb�(�Pb,j��ƩEDU"�j�ED-�*�J"l��e*1f0R�,J��",?$� ��w�8<�ڥ����֑�p�`�Cqi��DDz"կT1Q��^���I�[ǧ�o/M��n�|�|�;O�yY�!�~�G�}l�`��Y��XsӞ�Y�|I�����Z�"K������ؾ���6��4x�W/;׾�/�"�j��Z�3�����@��#bb�wg�ؽQ$B!�Xl�|���]s��2�T�N���4��s�q���cb��cU^�PG�CZ��e�f5�4.��}h��w��t�Ѩ��K<B�`�M�,���Ѝg{�1LVG�"�5�H"�˪ç�u����Ն���� ����gl��5i�5�Y�j�zts�.�Γؒ=(�ʋ���]b*[}<��m�BY�����|z��3o7�/���p��z������C3-��X#y|b�XXA��LQf"�?B!־�T�Wݏ۹��/��9l.�hqa�J���K�u�n~T~�{�"�2���6���(��=�{1��,���ɡDY�]�|r�-`8h�6<s�1�ŖC"~g����z:#H��wy�'�WK�Q�/�^ ���B��'O��l��(Q���j��ܡ��g�Y$I^���`i%�����ڹ|���
>?@a�Hd{�,�S7�[���xj����	٥{��GFT��,O#��G��{�u����z½}f�on��a�����r㭒�b�u�/ˈ�(sa�,�MLd�0�#h�.^Ƿ�˟_e�*���2��$x��i��u�Ú �(<bjΜ!�EGb�1�c>Y�}u��כ�1£�F
�;�g�@ֱ�s��!�ܕ�5��0�_'Խ�+P��W���Y�^-�� �a�9tBϥc�<:9u#x����ч�p��a�0�Lþ~����+�8��,!�^� ���ԃ!P�������2���qÄ�McyY�B�|G����R��]R��aW����3��޾75��޵�.��v���|%Gw�fL��#i]������@7�=����:J�:���~#LcVR�q�B|�.�a��9��':��m<_7e��q8�Y�~��ȋ�C��7Q�z��]�y�|�J�Y؃�c�E�F�9=�v���o���ӧ��#�Y��g��?(�]��^?�-0���֡�z!#� �q�(0�~�Za;�+���ո~ ����.�qa�+CB��5w���_Q������#փ�ӆ��|2k�}�1ix����B�E4����DɃ����ab"7x���m��g���qt���>*����-�|gd=Ʒ�7�ĀO}߾��fS��{����=ꮜ~{k�=��vg�ߛ�e�56�ߔ��'5C!6��'M�.�gr�ݖD"G�E$&!g��ZlݺU���#~�vh�Da�b�%^���g�
�@ٳ�(�E2��VI����ޖ(�����~������G�����;'�x�^����Ějr�Y��"�Ȗ�S���\E
̠�gUx." ���`@B�L�}=�p��${�����{�Z�����3�^������zk�Q�\��a�w�ڶ!yX�o|�'��i��9�n��m�' i��0�f*<�n�;,��}3�|�3X��J�{�Jv�Yv+d�WW19�;��	{�s�zΞ?e�	��Л��F6o�Vh���;���:A�/ǩ�D?�f� ie!��Gz��!��!�c�ۧ:���h�<zf�y�����V��Äe�䆴0�,<72R����v�ޫcOȆs-���v��/�׎��`�h0�C������E�6Bq�����k�k���0�A||��l��,$.���꫷��0��G�͌>?+L��gH�ʷ}�E�c��B4@����� ���6�뻳s��ѫ��H�Y�W+,�T��=��e�ߊv]��bzR�)ي��KGfة�|>ɪiR�S��1_s��
��Ewm?!�y� t�e��O���p�;%�g��Ao�=�Gb�<\D$��m�Ӥ$��ӓ��bR� ���Dy���v���t~��b���>#M(�����l]S��ֈ,�c�3ǈ�Ay���	#��:�9*���Jcqqlx���`�Gr��n�/�Q�1|0��C-_,!�!�� ~��̛����E/�UP6Gz1"���P��]~�^��gج�-��/�+&:�v|�r0�4��e#AT�n�D��$�����_(Bp�w2���`�ƫٻ�=�/�`:�������k���r�Մ�4hᦾ�B�C����ioOI7E��-U�GD;U?9�"�]ޖFe�*\�K��{".����]1�+6��:E�1wFs�?o��4�R^/W��d�^����?+������qf��/�C�B^1�����fgT�~ʿK廽���`v���)�Z�K�x�;�˾�_
�ʼ�?#GO�<��5�&�<S��7��d�,�W[`@&�,"�'�ث�ڄ��ր�ֈü��<AWfK4ɴ<F�b�59Cܾ��!�W���#֮�Iᾊ��.�z`X�{��m��L9���v�FtR�Q���سj旴�rp~}$!�|��<4���������ͽ�n����;�۲�������	��7����Ȭ�=hR�g���(�g��Xp����ӆk�[���/W�}��5̈́F>uPg�cur�|��Su0}yp]lǭ���KB>�ǟ�\�W�<CC̑�(z��;Q#M�^���b���a�!�ȉ_����.�T~����=t����x��4A�t�8q�=��R�҃�OM)�p��A�B��<l����2�e��:E����t~��]hl�]�5��k�����Yv7)��ö3Y��n���)�o�d����](�a����ĳV��舎�������ؿ Y�M���"������W��"#@o�j�NX��lb!�FR�x��_���24F$��#P��<�p�/R�>��û�#uQM<|p��x�\���o�K�{Ϸ���E�(�`�>6F���x��X����fѲ�jl��)�dvг"{�ǽU'����q�<B/Ul��+��(B���w��x�Q�-##�g5BH��]k�c��G���/�z�D"�li�e�3�eV������,�Q� �Y�ȧ@b�X�t/��c���`� 4�f�%e*��]�,�c�2�[]����n��K��9���x�Uפ�hp��6�FE���]*�rM�Z���ڈ�
Pܚˋӆ��TT��8���|������D˸6�:��P����h.�)5�x�4���9�l�(�E\ KI�9����Y��o�})$)������܌Q�J+O-�w�Q�ΥvvcR�b���%��b�VQ*>�*j�M�s
�}��u�sCkf9X�������8���h�^�3kڼ\���|8,�(�	�*�f�u+��^`�+v��v�e)Y���W�=���	/.Z��ٻx����ا[�s,p�ZS�%ET�ڻ��h0���Ì\��tc��+#L;�+����L�=!��3sV�]Q�N�Æ�5t�7��sz��X�͢�X&`��БY�lcˏ/L��r�����C�;��KKW
`��b�hV����9�c�ȵ]���8�lm���v���\�঵�mN$^��ǌ���ǟbf�ڽ��\���E ��6�Z�'<*�Y]��*`+�K���OP"t�����g�������b�Q�Z�AUYK%`�DF%՘E�bJ��j)`[%AQRڋ�F1LJ*�V�J�)PYB�1*`�,Z�"���V����V�X�mJ��-kX�Uk*[j�m,�
��1U���Uek*X�,QTXVH��F�0X��B�
�TPk(�U�J�+
��A �	{�u|�uh۩���-v�<�w��h��~��DF����z�-Н?��:�#ƭ
��Iv��/p_z�o&{k
4I�TGb���3�@�L�0��'�%8�,�a�Hz��!��p�r��QKz�Gu������ay�{흽����!A��̞߬�Fu��/���1�1��� "�';{��	�a�o�N�G��J;	�*����>"�|�h�BD�*SӞ@8�*��'�k��
>?@E:��::�6{G�m1"���\�h���ׯ����3u��F4š�&kˈx��afW�/s��'�����;�p�h=�+Ԯi���O�q`l΁�JEwئ��
�:��� e<�eN����~UW��\�>�N�g|�����ɴ?��2Ђ�$x�>0�`�OqK^8~��;}y׆�xR����=LL_*+�F�e�Q�CK������?j_f7g�x���էgN�fF'!�VI��l��$$���N/Ü��2ʾ��onfT|�N���j�o����k�~��6������Ej�:K⚽���<�NOK��U^;Q���šȕЂ��OLd�!���y>:Ww,���5ּl�C<GDO�C�p_ׇ���֝�۞��*����dw�{r���yN�YM����j�Et�������9��{��y��&�����Y��'o��m�t~�_q��+ˢ��"x���W���!�P���h�.?Y�7k�]��cƉ"�'-�(�����)���M�xR�0�<p�?KXa=�u�v�"�t�H!��_CfV8jՑ�H�}�j��Bh�!dY@�O�0�5����%]^G�(�Ç��0�3$441�B<טݑ̕�� �Bg����B�<t�Dbw�^^�o�h��dq`�a� �/��g�V:�xuh���%����k��ܓ������M�������f���l������:��DDCz��者`�C4|B�Q$B7PÃ��{�
ϡ9ٷ����փ<U�g�0���͙�N��L�o��
B�Q��v�"@��C��Y�$a�<y[�@w&~��Y�Us���؆�AY~C��B0�iJU��]O_��M����D{��@^�[���ɽS���O�nj����J��6���<�h�X���z�Wk�"|h�H�,�y�<����VWgm�u(3�yB���:~�c6vUݼ�e���G�W֬�h". 	��f07ע�9��@���Ǩם�ô�P����|::H��Ԥ�uK�Lԁ���-<��G�ڹ�}�.�y]91ݷ
b����~3W�����}o�o�É�֮���^^Ӯ�o���6�:]���6t�����A�qۍ�f��#*��xZ�t�ExO�!�E�,¹0�d <ϔ|q�=~B�\[Ak�4ED	�7�w\}�u��۴yW����;t��x헻:�Α����Q��x�!�CH�� Y���Lߎ�@�<pٳ���.#����*������1��`0G�u&��~��o7��r�4����։�.,j'���1	Ig_�9����Vq\:HM��Q�y�KwF�p�`�Ώ���i��;:����UU=�_�H >6C�!�~B�
s�9ӓ��[׹
������5��"j���
0�fo�����*/bq�5<��a�x�G�~��MP��Jx�G��{y�äaH"!�tk(��^��!����]OA=��d(}��ي�9����<�OuN;y�A{u�d�w�ol7�������i�"!��E w" ��t�����ev���q�\Y�g�"*b�(W�y�F5f�ys���9���=lw�B,�9H y�Ŭ&vɤ(�ϒ7Ւ¸S0�CT'6� ��y����b�ʗ��їRJ�O���q�_���+<	p̮�4;nU��b��s􂶲���2�G$�Z���ڥҠ὏��N��~#m�(������������zCt���V�!�h�ᜰ�~��7l�r�P�W<��_tXE�*!G���<��b�M�:-G�%���E�G��d��rٽ^��`,�c~�T#��1;5>��R��
�|p���Ʌ�Ŭ�9dB�2� PhC�y�%�̢<G�7�]+7�mS �Ǝ�3�,���n�G��#��m�kiVs���7���ۑ����ő�L<Q���~�ZaW�`��ߏ q^�� �z�#�}(+4r,���z���@�z���Mn��8nn\�m4P*�;��SZ���([�GWvw-v�}�7i5}1��a���3�������)���&�����Ζl���0��᯹����U�e�dIq��L-S�A�1��l�4P�e���^�p�?C��6D4~���6��v}��z�����_���(D?Q!�B�*�.:�W��pä7�"͑F$��s�d�$��chs��
�@��v��?,���sN�;�g�}W<�8'��۴:繦_)�,������#��jk�؆���C�f�m�^���{�jC˘}�I9����A�m_\�qzj���K��ܗ���4�WdU���N�Ky<�������W*�Ѱ-�'k�U8��������zǇ�FF�#��B�Y�5����խ]Ro�g&y
<D$�6W�����>��C��=_x��}`�l��=�*{e�.���A��~VFR
������}v�Qd3M:{q���x�x��h��N��G(���C��4p�5j�2]<������.�P�x6�K\�͋{{R�T��Xن9"7'�m�˃���-�
ԋ��VFvB�]��g
.gglRVSΐ���(�[�ω3�|�2@{"w�6�v�o�%	[*�Z���e�G3W��#fw�}����Rm�׻5�u��~��+;�@�sn����v����եt�.��.E(ҩ[F�y��ܳ\��g*�B/y(����6��ꬉ-f_<�u��ht[�!@Yu"�JyZ��c���F�M&ua�w�֊u!�n�ؤ#�
� Nd�<����Z������gQ�h&�l�-=�*����]�.h�3����G�G"���f�)���T���
�1d��y�:=�Ū��M��nU�Js�Ƃd7��ݥU2��调�H��i�����z�q55`ګ��#��r�q�l��N���S��+	M��p:m��g'gX�t�2���橪^�}�+�ۧXG&t��f�o��R�-�f�Y�9/f�t�z �����4ߗ`���h��y�:�cS�lYW��1�4Hyd���9���R�Z���'I���#U���B�ݏ0p�\�4�W[���w%�ob���&[��T�w���W�N��}0�	GM�/��k���>��c�^�9I0Un��qվ-*Ք��m$]o3]6;��v�1E���:�َ]*�!�DӬC��⌼���X0�	rR{N�Q�m1����<C��� �xN�._!5��W��1�@ChFkY��78*)#l���w6wA�N>�΢��(�|��v��&-u�!���=]�6���(�\�
�[g*	��]fd��m� D��"��j����-^v�D�x���z�����ݪHsk�3���0��N��������W[�m��v �����p��i:�7��ǘ��d�X�(}}�F���Zт"1D6�QQĨ��d�E�G(U*�5�@*U-*E��"��b,X��*KhT�j"ł��̫S��AY�W"���#RU*X�P"�ʑbc`����2ьQ*�*���KKR��(�2-�,b)1
�T��.UX�F �Ŋ��I�����q��o3w�3qybO�j���i�s���"3��/�#Ѭr|q����}����`\�6�0J�:�ٕfg/pA��ǰ�����9�;fЕg�`��ھ��v8bW1��S�m�ق&�1=Nc�ٮT��������Ä��͞�c�J\`@{#Q����+p�
�IW��t��dg|���N�9�>�%sX/:�O���oĐs�Z5s_9���3�j�8��K�},˻�N�;"�5���9t�����Nz�x_���?Ի�eSw"��ߛ��B^{d��u�sg�h�트\f��rg]�gk�sz���O�ĕ\Ƽ�U-�F�Z)eT��W1<��d��P�w ��p��t�2�׾+�Tpj��:y�7;�NYj1.�3�%9�z�W]�#��q	#�IV�aS�lp�ٚ��
%�TM��.�/;���3DzߕMɣB�_]ze�l������֥I�Ya�}s�w!����h��0�Jm�m`�;j,}���m�Ts�#uDu��3eކ�����GV�'�n5�=�"S����a���a�*E>�Js�N�[��n�#Z�W��'O{6{�:A	8��w��C-�]ƤN��:�W��I�.�G#��v�Nwb-Y��Ԓ�HzTd��ԩ���X�~��g�:!�v�2���1r��H��Y�Ȳ>�- ���x����1��C��	������쪯��9�/w#fû�����Ϋ�>Q��%nX�&"��.���}%��bǡ�T�X�C��:[�1q�����N�r{\���Ӕ~\�w?��9�D�!���;)�L^U]%F50ҫ�7��]TnQ��fs��|yV��!�m���zvū��OU�¶"�7�侄z�,T7q�\��i�o��ݹM�3�h�j=2ڥ
���T9u;�Vn�_���u��ȵ�FՊ����A%ρ���u�.��M��]�a�!�W�g
�tG�rd]s�-a��%m5��k:�s��������-��6���b�����@�->����)��_����M�}��b~���I��a��T���(]��`�K��Y~R�������qIh��l���5�^ �Ļz�h����BJn���{�(W��N��U���gi���������-:����/@��Vp,��K�#е��'�2���ј�B�j�? �u�a��2���0Y�e�t���ė\#m^쇦u��;ie��[��+&��Ԃs#W{�:���V=�i�ێco=��[Ы�I=ʛ?P�&�}ˉLVu7i<����3j�I�kk"�0n�.,��/653�w�ys�F[RC��L7���t=%�yˠBc�S3Ԃ�w[���:��Wm�yH�I���w)��Z�@خ��Z�4�Ӓ�5�O�s���k�����&צ������p�ǰI�ߌ�5�b��n"��ѓԊ��鞛Bv�ձ����Q�l�7yH6Xw�
��L�
cV�ȗ}����[�YUY��4�<�ݒ�Wa�>R+��a���ɤP��}9��f���݇�wTEѵ>�}׽b;�;�u��< �g[+�nv;Ǳ0UBp�d:��
�B�gik5���Y�_�\�����*ݗ#N��mw�}:^��c�Z�i����1^^�I��۬O��eE�d�k�n/Z����5h\�u1�f��;�sx�1�[�uȧ�b]f�ja��D��Z}9�h��6r�����(��Ya���l�<^���_d���E*��Q¤&�����ټ��YU�)~u�ߓ��y,�/<�n�R.�P�>�#�6�`n��tU�m�݈b ���r���3{ò��,J��w�1t
�Gs�%�G������ �Z>4�����H�EVy�N�x$f��k��u��mn`Pu홶	�&�#70IV�����[Zqe�����Q/�Z7��6:k�[+����"
l�׻�?ncT��'�?dˬ�P��{�������ǆ/q�:�y�_w_+
����^ޑ	���S� 88P�v{�q˯b,igSwu���� {܂�J'���{tX=gus�P��׫�#f`,K�!٫興��i�������
6jK�)��r��%�D�*5��oA93�x�fo+pѮ1�+��R@d	��At����+|���|=�ǹ!+g#UY��
�-�l�	�A�ؔf��p�,8���K�ɢ��\�곞�������V��s��;�U��qδ ]��l��އ�pV��bϒg΍�����뮊��B��4@���1�7/��3���c�ʸ����#�M��8���>n�n�[�w��7b�-�o7	:9�CFUgolz����w�[��ͷ�c�۠�͚���"��B;ۖ	w��xd�;��"x�_
i�.=�qظ�ީ�vF�3�F�ѬT�Pn����w��ň�$C7�!oX`�&Z�7�;)S��5}畩c��e��
����m�Z��+�����nm:U���J���4��1�Ed�O�U�q��O���雋&F��mrU�p5���&�MNh��3S�ذ^��41+�.�P(sc�0��ڱ&�C1	��*�q�	,�r�1Y�VN`�v	5j$R3�����$��V�Us
�X��>�V0�RH`�eg��Zr��#�B_�*Z��7U+���G ��r�	e<U@��Ӷ�h�H�+�WFە�+�rP�,j�J��Q���E\���/����D�����:ȭBj�P8-�Cd�VL ��0�\�2��2Ҙda\�p��T�ER5��Sp��]и,���y�� G�~ DjbL`�T
.\qPP�Qd�1��Eq(+��E"��������*�F�J�1"�(�X������
�h�+E*,���h*/VQ�c\��b7[|���|�[|ޝ�\;�ڳv�di�|/��ţO�[Wb�y�,jiv�R�7�q�2J9�_U}�M�MD?�2.,B��ɫ��Goqe�a�`�����8a��hN*lp��7�o�x���v�ɶ,�G���N��b����[J����(*�Ӽ�c��5وX��M�ʷZ�ܨ@�wV(E��o�b�dk�6�b�aR�.S���^t���wݸ,�n���V��M���u�gp؆��x3�Ī�7&y��7y$�cL�W�#_��|=)+�B��1�#���Q�V���c�]Ѫ�zqf�x�`d�ap#���Gm6�q�p��Y�y$E3G�v�:����Y�&L�קf��0oz��u��/ͺ�a��4�Y�!���Į��%�����cn&߲�\����YC���KF� u���v㎪z��m�B�k��v�jΕ}w&~��M[�L֋r�#ev���}G���L�1qzyn�_D{�rj���}yF�q���_V��ٛ�ngBذ���nٌ��V�zҝ���qm( �}��vV�Vq�~ގ���X�LT���~LR�λRɪG0��Z᥈(�R\6w����X���4*C\���u��U(��D��ZD��O%cK���������~=~/�c���F�bJ�ۄA5�����q����x�m_s�('��婨;�s����Z6��{�deG�>+-K+s�b�~g<Au~\�^�l�������֎�r�;��ܕ�p�c���F�~��9ϒ�8�Tj��t�+������w��æL4*G�_i��RFnM�:���fPJ�F�N$Y�׃��7ٌN��hv&�%k�[fssl�Ȥ�Fm��ެZ�K�w���z��ns��+72c������մ������>�C�������й��ޖ6��������iSʧ:��9C��p��2���㔹�8q�D#]��FPYE:A1��=�y==<L[,�J��k���ß^�י����ػ ���A��Ff�O�_.�`a)Ƈ���j{���k^���UԶݒ��QMWf����{GM�ؤ�����&;ƶ���m\���}�1L��䯀��lL���{ٕtۙ��s��Y��$$�O�Z�V:�jH-�"���_u`�C��+��Z��*�����[�p�8ވ�	���:�����n�y:�s�>nt�ʳ�ʧJ��U�D�z�M��B�E�9��w�뛤;�='�>khœ�y�X�x�t��)^-�N�m��L�@���v�e!Ɉ�v�uqg	�OyӁmu�Wj׏�?yul��!�mn4Z;��K)�cue�r�)	�h�Ѿ�Ւ��v  �8��#����3��Lp׀@j:Rlw��r��=ջv������K��
tǯ�}������st�����H`�Z���0�����x��/B�8y�t�7�_˵�w�q��Y�+%�˸��Y���D% ��n�ح�z��پS�R2u�>�Ί��.Euy�/��\勋[�e�<�������Y�8^�:�nM�2�$�^���ҧ˂�$8�oV�P�yk�eB
�@����9˗=�g7���k�L���.��3������^���9Y�(�ԓ��_!��g�zz%�L1�+���_3��ԑH{U�P�Y�X���n�E]r���Pg{�j�(�1n�y2��캫���9]��p�h�*���8��j�!��zuӯ>���WP�z@5&��x$p�M�NΓ�$�͘'6�ϊݛ=���\sx���Y-^��'u������$�'�9�=��"<�MT(�/a�ڮ�p�ۻf�C������3'���M�P�p��gNm�.1φ���>����{�o\I���]�������Y{��JJA����>�y�B� �ph��Ko�R�B�x`3kP�8�I#��Cu���78��=��/*�0���Cȴ��:�ˆn�d|��cNL�m�.˾��r��0on����z�w��w^��+��6݂mb4F8B��'�U�i�xFSі��W��^��拃R��z���}�ޅ*:c�L�Wv�*�f�4#��#'*:��q�1J�o	lCڇ��r!7��S]�IG>ݙ�y֒�9*g���~M4yA��I�S�E'\1��@_C[pP��H���: @�eP�0%��?]��p'�}{�g��6�ݜ���VLԊӳ++7u�Jp�x��7��M��GiT9����EĦ�a��u8�Ykw*U�yj�p���qN�3n�ը��R�6s��Վc�c2P棣^>���DY�{n;ֳ��,du	��r��?������ܽ�ڃ��mn�^�AЮ����p��m�j�X�@�Gs[Z7��Ic�5��wr���,�w��T�-�����q�[��+[ۖp|g7��}�����ܛV�p�{�z�0`��fsm	3�^��X��w^-��]�nn�-}��i(�M��:����ȑ���1L�B��G-;!�a�
�"5h�Ne��s][n���c���A
h���A�`�i�[2��%	NA�h��&}�X6i��Ռ>�,(�'�d�X�F��P�LBL�;\���̠ZĔ�Ȓ��,X�L-,�эճQ�rTh9h�V]�7bꪬ�AА^�l����i�72|��Rg�R��U,%E,���Meh�X9��P"�Y�����fCeU�Q������Zt�c�l5q����A�R8rΐëvF/٦��C���:J(��J�(i3 ,�m�h���9�VW��)���eeU�E�Y`�-XҶ�q�-��mk����&ben1qS�jܥAeAT�n%aP��*����tj�e[\�b�2��\qL�-ZJ������-��s3�U��-��kZ�VKiK���_&�goPTdp�Gz�=4�h��'L�'t�� ��q�7G�nkhc�����栜���dw����1��ct�`T��s#"cB��9��+n��n��˒�f���I�U�S�δ��cVn�)��c;��X�����4�n�ey�҈����9���P[\M!L$���ޜ�����{Y2z��_k���RZt��;r�u�X��=�[Z���D��^]�ـ�Ɩ�8���W���#Y�M��C��]�{8��ΝW_t�Oٖ�k���
�1�*��.�s�'u��[~�ͪ��2���묂���ތ��cr����^���g;\�z<�c)_�c�D����
��i��r���^k3:���4fkX=R.��uҷpg^�B3�7yv�C�T�R�!���˳���u��$c��i%1�SӐ�1Q�i� Q���E��Z	A;�e����NG�G.�:�]�S�����4gϺ�h��Y	f�[[�m,x�Ţ��j�tmd�%K������VP�8�q�=��j�^V�W���5�:�ȷ`�0{�N�Nn<��i�=1��b��1t��y�v�}i.��=ב-u�{��΃;i�΁K��^�A܇���Y���8�^k�L{[�����G��\���~R�*j�ՍkЖ�{��ŪA���:�\_X�w=\F��M��j�@��oNtvx�ܼG�E�uP�hT�%�L<���S/9'�����a�t.�{-�b�������V��ތ�Zf���,���Tj)E�������B4��VgӊU�-���ڪ�N�c/Uʊ.�<�PZ�4c�B͗��q���=y���T){75X�|]�u�t��B��h3� u(�z��bߖt��胊h)����Wo5N��vU���vXg8JfV_){���c͜\���W%�����J�yE\5o�ε��H�OF�3o��;�\�Y�q�/h���$ݡFhW���C�w�Lss��{cJ�ˊ��Tu��R����Bg7��]��x���7J=�ʐS�U�⽬�|]���@�;�[E�gV���z\�w�����vh9��YV4�_��wQq���0��-PK9�>�^��V�ĎɊ�>�%�f����W����N��E$�e�G��z�r|���4;۹����e.��ٜZ۶�y\'2��'�92��Z>���P�b�ɳ1n7����\���84�I����n��-�vc2ywYF�zWvFZ̧-pQw���v�. E��"���lG'�+��q��*2s2��6���i�t��F{[���.��.��Ո1%NJ��R��C׸Nx�ާ�U�	�_L�[@֜��Wv�-��������R9����k��}/>�Mc�V�f�Ѥ����m\/�$|����P{sKˤ�%T��򣂻L��[�<�ޫ!kA�� �b���/rf�b4�-B����}�p2��,+}�%V�N���$v�Y�7������u]9�D�;�0��u��]�1�GVS2�Yٕ�VZ�8a��˻^��i��J�`�\K-�����Y�U�Oj������G;\ھY{s(��yb�E=�����w�4�J6w�$�~�e���`)"�$� �KeҜ���)$�FQ�q�\J5fP���Ιi���V�E�Uճn���Ԇ��7PRӂ���t��l��� <vJT rU��U�[H��՝�{��gY`D֪|^O;��hW�����>��F�x�i����9��M��a
#p]�I�h�>����z-	����vytR�j�rx�<�NQ�����]�����9�������7e��T�hM��<x<��\Mv��;k-��A��B���|���n<+�����MhY�M+���,�ܪ�������+�bІ���m�u�j	������/7���/W>�;ڎ�� "�{�q2�|�"67C���!�μj�^'��;z��ef��f��#1,�� j'�6m�,��!���Y��$�a)V���[Z�c�{���s��t����ݻܭU({<�9g��4Nm�f����<W-	У�0e�P��;|����.��-;����X�x�0J�v�V��<��;���,�����nk(�*!����+'��՚�nɰ5�m\�� $t����+s�k��]:Β}a����۞�=�U��&�1����ʮ�+��~�r�Ӡ5��������IZ�rb|��v�	ڳrg�Q�M�����&6��%[:��{EYi+��eԥ6 �u)��{�ӓ�$���ve��f��܂åt����������6�})�ۓ�u��ʁ�U��g	��T��Y�r[�`!E<�=��X}�a1g�7��uEB�U�k�5;��H�
����;}5�
��k`�~Yo��	[��G��v�|�L\9�&�L+3IڋPYh������5P"Yd�β_d��:�+�>����8畦1E#W2�L;�v���T���k7]Yׅ;��лq�zûd5�iܭ��׀�kF���q=�q[w{��iE��1��uV��IE����M�X,b�2�YU�!�#vZ
`b�Ie�[�"[4��aV��X��L�`<e'�s~2Q�[
����Ka¡�Jٕf凁e2)��-�l�p@P�cb��(�[v�A�CY:/Blc�QLk8{����~΄Fյ�+-�c�,0L0�r���aZݙ��*j���Ȫ-E*t���Ymb�KE�Q��2��Tup��ak+f�enV��"�"j�LL�ZV�fdh���31&e�\��M!c2�ӥ���R���S9W�-�M*ѱ�3ꕘ�KZ��bMi�bb�]%t�.\* BlQ�?S/�wv���})n�!o��ʜm6����m���]��n5wD�s�E��	ît���N�+��-�<o�^�����T�#p��x��T�wy�!��W��el�Ʈ���5-�U�=s�5I5zz�SfkO_�!w˺�M1��Dgkc3|��u�!��f>�0
{�e��!�����t�j�	��ȉI�kƐ+
qZ�#PpR�0�w�G�S������q�L"�u�΍���Myds{�Z�H%ho1�ۖ��Έ��5�(�1�&�����>�đ���\�.cB;���a<���A^LLV�\u�l�p^R��ڂMG�&%�w���n�Uu��Z����l�v��~��Ɲ�)9-��q�2'7��/r22:WT�w!Vw!��U�{~�;��w��{_���Z�)�K���M�׶t���)���B���D���[vs=�=��A4?��C�o���������e��g�nf�M�Tlǭ�k���rGy��~N,�|��u"�wo<j:}��%�Sq!���Yv��2�Du��.Ğ3� ʐK��s\9�$S���Y\��gFW���m��S��߉ˡ���7��ml��U������@�vI5�]��-G@��۶o�����e�m�qQ
k㞃�/J]��Ε�n�{{�展Wj����Z�ێQ���k��T�sJ�غ����8~���K�:7V"�+^e>�[�i�eNS݋x��޸z;rt ����%�%�v�b�����}����1�"ᔴ�R����=�9l�Ӥ� P���Jbj�n}���>1b7�����Ε\U�d�FU�!�f��{����z< .V,��������{�J�
��2�]P���y
������n:�I��Z��;��7u1v��^[�,��n�nC�'#|���~��|���ܱW��h���R����Q$�	�s�b�=�ՈQ�c�c�cx�P�ם-���O��ˀ���[y���+��>!WI9��{wv�F"�^�`���^�u��&�D�8q�'K��mc��b����Opƾ4��������)�Y0���U�[�)�W]�5I�v�B���۱��p�]���qoRK���n����������{+����������IS��*��:[9roe��G�ǼW�z욡YO8)��*�YgW+���)�V�bWb���<"ߣ�{�ꛤ�XRǕ+;BO_Y!�M��պU�Pp!#ꭚ5�\�[=����!��Y��@����o��.�Q
2�H)
�P�7�B��{�z�7��SWee�{�|��\ڼ��IKU��Ӷ�1{��]OĞ7]:*C
ܤNN�ƈ�2�^�2# ���e�ʥQC�y�.�I��'�� �����
z����j���};3{Su�;�2��+>lt��{)����N�Q�{�5���7���<q��sR,<���_�n�b�:�^�%
�p����x�uxh�n���Q��ԀL��9�[�u�èk�o{z�0{�r�f�s��t���'U`&��U����l\L�y���OJؚ�KU��{\S��!_�c'����u�|8���b\`�#7�1��\�2�:�MD`Ն�!B�S;�rɫ�Ǌ4"�E+�9Q�Zi"Zb2ܦО@Wt�޷
����ӥ� ǝ��'~�-��㗰a	��+�|�����Ҿ�l��]��`�;�:�hVݰ�0M��Ti�V�,!�cs8����Z/Od���BG��}��wr��/�=5V�������j>�V�GG�yv�[V=(��r$=#0��o	����z24sZ}zV;ܩ�b�/�-�B��aV��Ym�X��'��~�KO�X�45`>��������^ڛ��v�ء�Խ{/���Z��{�>����ݩ�V �R�hb��wJE�~��o��/`Ț�l������kt�g�v�I�B��^uGVu���)Foq9�����fw��3�_��[MT�o"��������ֹ��Wi����P`��~ɟl˗���/-��u�x��}n�ܵ6);��uUٽ��,��[Q���}�s���5�3sT��$�#�*-���ۛ��SQ�AR�"-��<��[,NPS[]=���&B1[oG���G��w�S���iٌM�d��pgc���[dJ�B���x춝�T6�8^�Vmr�he_Q?h�P����(�&o3%[��e�zM]O7���P��]�H��1 �Hț/v�`E�(��^��z��7�k���1��Y��%��7㯌�\��¯{_Cz��ׯnp�Zn���]���v�� E�À/n7[�.��{2�X�@������j��J}�(�sC7��Et�ٷ����в������;w��uf+�Y�t�+�'`�joL�x��$��:�M|7F���嬜�(b\������ηV�X�Q-t:��.FE�7�����!�}BU�.�ȸ_�0�z�3��r�2�rCj��h�r�vj��|-v��W����L���i�2]Ys"چ��3x(F_۴�j���p8&E���٣��J��6h�2��"��3����yͥL c�v�%��t[���/PZn�����"d���@o��V��wupی�zt�T���e��՘��r٬��t���CǸ���<ul��*8����a�)b�;jS�yeJ��K�zjƤ�Q�Uärؖ�S*UߒxOKk<��c�TtZ��-��˧meU�-���Xi*�-
���噕��e��c�Wk,�t�,p����*.*r���4�,J[KX�.e\2�L�na��Z�L��S4k3%Dr�s*-�h�er��QT�+qrՃ��.�b#���5����Fe��Q�n�1r֣���i�(iLs��U���8V�2�h�L�5K��F��ޞKܟN�+�GJc�uܽȹ�Z]�3�S�;��EN:����v��6��ycZ�ިҾެ��y=��ׇǣۉ0(�sk @o�p3��(
|.��S�U��[��˓�S��#5�?s;�ȓ�3/������0!u�A�28B���l�2����Q�/������,�zy��Vy���r��'����"�E��tSŚ�DeF6�el�u�֗ׄ���M.���Q��qj���.�'.v7��lX���1訅�����:�G{�E�C���M ewg�n�K������u1���k!����\�
��]S���9�/��/�Q�3���Om"�6l��(������⢞ߝ���.�J��"��+n����{���4��O-�B�-]�8W1Y�����T�[��K��]=n�4��$��+�uz\���/��綳�|6Tw}�-��Bd��dފc=;���>I���jeM=��N�d���f`b���y��(=��aВ�Aq�Jヲ�����vt�ܳ���I�R-�
,=�wX�n�	yuc�2��>=�-؞8B>��	BaӀ*>���fjq�ʮ��=���Y�5SVpg*#���s�bļA��_�����)�U"KN��Q�u���ޏ�jnJc�*}�wa�[s=�q�Nt�N�}J�nH9EXp[�hv��fw_/�R�W����]���?8O�K�sp�|�ל�q����|-ʬ�S��A\¯y��穭�K#ݯ��͢=�gN'}�u��r}�GT����`e'k2uv=7�S�dֽ�K��֖[��Ҷ���)̓��z�Q�!f����z�,-eS�i̽k:3�x��
*����1�!ɡH�WTpa횚�N���_F=U0곾#ƞ8���+s�Ֆ���2Jް}{���ݨ$�m�� &��w�<���r�7��� ;V��0xj�L}��t7�t���"҇�VM��֮�MϪ�Μ�T��8h�]��!Z5�����]�S�fR�		�]V�������n�g@t�j
���V�!�J�?Mc-�9��$�r�P�*d'pP�q{�k�k���fl�;(R�'\����ٜc}�^�mz.�-��x;����L:v{X�T�2����3f:����rJX��0&(E9�0_Y�&�wo-J9�F�y����*=H��|s.�Vf|}����;�n�;.��/d]��MY���DBnmã|�GC�a�$�cYӟJ�~7o+��^�/��]���I��nܿ6%�J�ɍ���f���n�t�WL�s7{}���v���\R)D����}��%�)�����>^��)c0�>��4�ݼ��ݢ�	�u�Ǖ+�뇤�����`7|S�#F��'�B��9X�FN�ʻ)�班�3�/M��sf���!�x��HMB��Q
`�򓳝A`[�8�2�TQ�R�mw&ʹ���ܜo�3�C<�rߵ@��(��>/v��e%�u�먯�jE9ӷu�%&�=�<����,S3���8zw}���Waѵd��g�҂�f�����u0�Y҇X���8l�)y��hb�@d�U�\j�n�&�RYbw��᧍_E<����Z^�r�D1r� ɧB�e��dO�Ǭr����ǒN�n����d�H{���I���rEh}aN�*���jg�A�ר�h3۳+_�YB*���].�v�h�0.
[^5ȟd�*�Y�-h�ǳ�P�Hݬޥ}����zL���y�ιw�t�����R{��szE�Ϋ�'���]B,���I�˖ ��}�����(��d�����\�7����sV���;�+��Q�mo+���3�k�?�L%���`��"�Ȱ�#�eHV��\��&�^��F*4�-nm��r�\�Sݏ$*�;�� �cU	�m��W]��EO:�ْ̹�:�R\z��pP�[����MWb���>O�|qi��j.�L�W���^�#+wf��d`���dM�|J�W�}Y=�޸��ީ�*�n�q7��n��Ә�ӛ�w��e$x�  &t<�;�R��dɏ��m��e���ɸ������*:
�h8�֨ǣ�;Uu���ퟜ�C����0��iZ����I$ �YC��*����J:
�*jڇ�#����ˢ���6S]���h�:��ہ�� *(��+ڶ�|�Ֆ(�KP�m	xb���_uQ�]��Z�wֈ�������i7��Ϧ9���5v�:��Ҹߍ�S�ƶ���/�̠e�k�Sk&a� �˕vr�M��US�M��צ�t�3� ���(
*~�
����qFD���5����Ɓ�?����<�P���?���w�yn{�%�TEL�`yS�W��2A��_a���MH{Z�&�o�t�'�����k)�\!��;�x��d�n�u^�0�+�A�?,DT�^l�m+M�=��	tTEK>�P밆���)��Jcu2�J���s �.����OTEM� �q1ޜ�嶾�����v��,���m���y=��4<�
̼\~�6��UR���eW�{Sv:���]����=���
Uش�@����˸�Gc�It��z�l�պ�P�1���=�F�S��@�Ϗ�H���fۦy�s�!�%�O<�;�.ʽ�������{�vФ���2l�y9�
j\}�¨���ՒB0}�V��@�1�2TT�[�'G�I�O�a�5�=3���V��~w�NĪ� �bR��E�[:��,����P��v�ΜQQ%���>Ls=��q��}�G�������s���	PN�p�j3�t�I��^�z��dOZz�=&��ßi�[���"�*t��8N2x�(Q^�O���"�*Q|��fmO��<�8j}/w�bs&׀57��bb�T���P�
�gU;�A���xk�_�hG������}Fu2t���w]S��ĸi�qⒻ��c	���9�wpc��v�˖)ϙp��b\^�C|(
*L�a��y>�#�ˏ-������M�m���ݘh���^��խ�&����]�������H�
&#��