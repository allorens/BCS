BZh91AY&SY-1�8;!_�pyc����߰����`���*B*
��E@)JQ!ABgaK�l����U[f�Ҷ$*�L�b����ݻ����7���xPP� `} R� �@�T(U �ۀ$=�Y���}�|��u��N����\ ���*^�c��}�ٗ����3���144�`�!x ^+�k,�M�Ѻx���X��ow}�ϫ���`)��=���ow.��{û�>��>چ��V��֌��ʛ����/o��N�xb���Rӷ�w{��:`�T7=7y���/��ھ�t�D��zosWjkE�<���
)|�����^�w��m�.��ǧ:}�{��z��m|s�����:�}wjݩ����ֺk� ��#o� ONŵ5���7��i��]ݼyׯw��;��񶻹��o}����O�u��*l�u      �     ��  �����0� � �0`OBD%J�F �L�  �i��%*F���     �#= �%J�F &�i�2i�4bI *D ��=��G��0i�x��(@�U(M�S�&&�ɉ�d�&��R�! H$�� 2*��H$����A>ϵ���!@�s�< )�-D�ac��+��@S ��Q�Q�A� ��uB����?�3�ެ�DD�#�TH���B��%	*I'��@��t�I$��mU �C��o��'����߷��A,~bl�o�p�Z1?l���9�(�	!�|�!�d���:,1���ƌ�8�0o�?`b`N�tc���,&�
"؋����jL&P~e����*����%��.��xSR��)����ŽJ�e�@X�41઒��$�����["Z|�臠,KUl�r�B�&���XQ�r�vU6���Z�6�����޻TYKE)=!�d��vS�T1�1�̃(��NM1ln0_�$X�!�X�@�$��Hr$E��
��D
"�43%��MF&��1J�.+�C��`�1�黎�,P2ɍ`�a}�j�ނ.9`��)��5h��- ̤m�v	�-ehZ�[�!������`�H0��0�A��Z�v�U�R�k���K}Z)�h�cB$`�"�`KN`cU�,N�	��0����f炅�c#��,@v$8?!d��0�!����[�]��U�d"*EHR"j	��ű�=��p���'E����h������.[%����_K��:�Dr�D���}7K�J�ј��+�#F�`�,c�^�SQ�ΰEH��D�NP�.�3���3D��2H�N1� �����H�`�1s��us�oQջJ���Yv�b'VV������������Z�0�l�no��d�d�%�dn
ñV"��Aփ��$݂+E1!Z��^��V�^h
�T��1���n�#io"�k�4`��ɫ�	�L��l���v]�Wm����h�f���@�7��{�N���F�͇m��ubWL��i�Lٚ5b�LT��]4��I�4�$�$���K�ԕt��/--{�;��d��������=-�%����
V�X�%��!���r��*��5F��t8���^���3��gp�[���IW� Х��W���=����ޕ:�;n����b���CCKOC�>�/�!��ޏ�V���	�V@��t�h�N�G��V%��\YCId��)i��).�H>����C�A���7��G�R��"���Va�³�)�ׅk�`�%���4]�K		�M�ͬK"�qI8�����J��Ԕ(��d�'J�J�I���HzSgu��^iY��Ě�[�{��3X�L:�q0,�#xF��n���2!ha�<d��ޖ���M��"��Mh�K��%�L���4��+z�m$�7%HooDj���ݗ\X#,h47��+[/5�Y8ZԷM�ҳA�H�4g�p�.ʫ��6��6L�荍�f�%��.;'JZsK�I���6wN��%#�I�3�7e�bp���U�m��Nm��J�%D��-QKKƔQ}����H:�Ӳ��qmC%���t��z��]"�K�f��G7c��ٶn�CN'��af�A�xb�t[�����$�c�V���j��46��{x:�g�سti�)��K|o&[͑�s@���l�4(3�b��7N��9G4�3����8��I�#F�K�ݛ�l�:���t0-[l������*��/4y��<·�3x5�	���7�����f��᥎RN0���+Y�eS;:4H���
D*��;��gq�l�7gFY��cҞI�Ԕ	D��I8���e�!�!�C����\�[c����e�ݦ��Z�Mh�I�њ8�K�Ki,��(h�E�V����:�&�-�p��Y���+�����_GEX�T�CG.lXh�.N��7!N@�0���vSNl���U�v��We-Uf͏85��*u���2LU$Ŷ��)
�Mo��i/cEK�&�6��)@���0\�z�qKEQ�������)l�pz�n�1�-�̌��$�%�Dd�7,a4YSVX��$�e�_��2O��We����e����a�"���c�5H���q��}Ji��J������k��;�[V�@�L��%�m*�R�^,cIPh������b(�E!>a�B�!���2���D ���v�N����f^��-��ʡ�A(c$����'F��&���3��ɋk[ǣ��64�\���C��a�!�cj	֒�����౰X�iZ��[$�tA�$Чi-�*CK�̿3�$�H���Ȁ�N��zSR��)��J��ŽJ���i)�c(�w	;��j�����)���*�臠j��w:6�x�jl��X�Lk�����M�xϘCcH`K>�Ȁt(iyA �b���bF3�20[22	9t��K�����0E�BA���pN�%����#x�T,���Շ���MhuU�j5\j�hձ����>?��0� �LY1*���Z$�l{�Y�K?)$����_)�fۈv=��m-{[<(g��
x+�Y �/�:k	<B�ƞ�-~�~NE�>�z���_9$IX�	
�������P��f���'x��'�&I"0��ى�d��3���2$�(��������������r��S��5�d���&�����X���@�J��p���×2|4���2r�|�x>	�'�=����ӃO;$ݔ邍oF �Yd�3$q�,��.�Ϯ�O�t�q�G��O�C���ɣ$��&e��م���Cǻ�g��#�$C��!��<�V�sg_yoB�YǑF�#�>�y����w�ݽ2S������ɜ<��с�Y$����g���F���aSZ�s�5TQ]{��'L1��I�����'�s}��5�Ν�;G�ӻ���a߽5�����I�f�3������>:S�!Å:S�Hi�>��`��l�o�߹=�O�
�f�Z|0�< BA����%t��\�˩�'�"�<`�ʨ�WK��W��3J���y�p� :Y� �T�$�}w�����>�f���3�(�J(����i���0�
�/M�<��/�3��ț��O�g>�  aD��<h��Iې��1�|�f�3�d�N���\���O�W5�2ɞL� ( >8P`}�_]W��>:-7�+/*��EaQv�d�Ԓh��d	�:j�,�\q�e3�{v-o����!�
0M'W5wxb��>r�w�Hv��(�n�p �D�>���v|(I�Tߥӂ�8B�ܭv��|��e�ښ섁W���ۢ�d��F?���G�jl�%��=76Y�w.�}�>/�2Y����`Sվٷ��vM:et����<��Jv\Y��Ɍ�3y}5����I��$��"ʬ09R0�|�Q�	!@=١������O��8t��!:�:|t������[)D�.��/7��9�L;|�k�M��/鷵Qב�ʉ�,	,g�Se�P����<8wnty��$�t�
2'�٪]��ӊ��J6Y�S�B}ف�>��?\�of��@=�Q��Q�J�4i�J�I0��A���t���Ӧ��-{�6ï��7c!C�}�����N������W⛺�˽SG�A����oc��c�>���}N=��{df�G�'���l��
s�{�n�f6,5g��!�b�{�8`�;?.NV�
Rv9>�^HΒɑ���)���3fs3%ޜO�N��b�5yT��������iD�rໃ�&��NF�eg8�F0(8vn-���1qzwlɣ�wkO���%��C���s\��8:��q��rҡ �,~�]���I�̳rg$ndӄ�Y�,�rz[�m���x�t�3h'%�������$�����}Qd�7���V����,�΋LmGd�*�:YO��M�]v�0��f�E��ۻ��<@�7ݛ+�U��u�>p�4���`��ij`�&)�9�k6������&�:y㜰�@M7lc���;7|<<)��4���OW�r@O��%8.�N���<짤<}[�I���Y��3�4��f��QӥLi�:`�&��;����DT�s���`2�,�Ye���џ� +�U���#N���J+�6t���I$`"��#ر�ى��*b��0x;��NKJ�(�GN���:x���8Y.�ʌ������ͲO[�ۧ*{w��IҖ�<pұ{Ԓ�v�f�nf*���d��@�]�b�xm�m����n��������:h����:4.0:W73':hp�'93���'��080	|v��y�!�Q]�D5�:3xViV\8��Gih�z����>3~�K@߆yw�a'�e��9v3��)t�\z�_"�����e\Xv�.�7&ǔ5g	:Ҋ1��p�15um����D��O8$�vt��\��B�P�(�V�{S$.���::U�h�����0��ΥYvi��5 #�ZN�*�&��**�N	C�x^=4��I#�����u~1����������3�s"Xx��|&�?mw3;}�ؖ�;�v�xf$���P�"���ӛ�d1i϶D�4���b�>>O|� �>�8O~�#��<Y�1�^Z�Q���p�[� (��	*`{�4/	+�����
8H�.�5�]'{2E�H cQ��h��Y�%�i����*�}S�!t���_��D���^��'��DFy�$���ل�$��ĺf�҉i[�����b�a'�xX��%(�G�	Io�?�>���~rB��|����!�OR���>���!�$|�'�h�c�}��g����T���V�M!��Tv$\(�	[&(H�jt��x*T,��}��&`r4k�����i�2kչ��w�sLI�x�^�}��p��JkOA�C�>�(�N;ʷI%�vU��F�S��%jrZd��B@MEɪ���(��]��!�%��`#���DSP���T�e���B����녦��X��&�:��Iki�b�p֠b��*n�`�b#�T!�y�ӛ�D�
�}Q�-��X(�9��,�U�RJ�y	��q��Q�gn�Nк�ެb+˙����I�nXBZ%���E�lZ�d���^~�D�ƻ:�q�(H��������sv<�5�+4�f�FW�!�M)�̚'�V�x�R�jmq>���ڶԘ�^��]��FR���)�X(�V'B^G����>5�D�E��c�?_����]�jM���L�b�1bM6�cX��
�-�%εED�US5%���[�--	.��Չ�/�YRVt�bc#T��u�L�9Q�;d�y���M�E`^�C��M�(�Aj��B��L���Gs4A�՗*z�W{��Ƶ׽O�wMu�)��������Z�N�E��$yD�E����NIgH�����7���L�Hn^�F�sY�1���}a>�5��Qg9^��ƀ���G�?�������B�I�����>H?o����;_���cf���r�n�m�ۻ��m�i�ܶۦ�m��6[m����m���޲��[m��������o-��z�m��6�m�m�a�ۦۖKm�m�v�no��^D��5AR��H� ��o7gF�mӆ�0�&ۻ��m�e�ۦۖ�r�n�i��x�m��l6�m��m��=����r�n�i��x�m��l6�n�p�m�M�!��r�m�m�-�� �� H����(��(T
�H��-@^۬�ݍӭ��6�m������m���m�m�m�m�m��m�l��m�e��m�������۶�m��0�m����m���6�}�{�[o{�������QZHj�e ���wr��x�usm�{6�6ꮪ�m�e��m��m�m�m�M�-��ݶ�6�v�M���^�m�m�m�M�-��ݶ[m��-��m��m�ݶ��m�n2@���O��$�  �<r�����p�o^&�n[���m�m��m�a����m�ݶ�ܶۦ�r�n�m�m������oYm�ݶ�ܶۦ�m��0�p�m�!��m�{4�m��< � 	�G� 6�fmh������m�uUR���۶�m�ް�m���m���p�m�m�m�M���Ø�m���oYm�ݶ�ܶۦm�m�~m�m��m6�z�G�m�--�*
Z��g���"��$��/�?���}��W�� � }A�?�W�?��o��z��o�i�m6�l�͛6ڻm�M6m��Ǉo�>+f͛6�l|�n�m�m�m�m��+f͛6ڻ;;Uvt�[m�M��o[m�ͽx�Jٳ�f�i��m�m�m�m�|��6��<xӦ�m���+o�|���6����m6�lV�y�~w��{���W���N���)\�]T�7�X�C��Q�XF!	�Ggj
��G�Ҵ��&� \�v����i�D!р:R��W����,��!gMRM�y��݆��ҶX�G:D�̲���q�K���m��j�V�L�ڶ�uv&�5n5�+�g���ha�/������k5њk3�nչu�W!�˫�+
��"]�\�͋I�&DIEڒ��6����J�誨��g��a�������l���A�Ĕ�	��j�@��cR}g���uA�Һ�29ʢ(!Zcp�����Vcj���(:ǳ!�p����歉a��[H�GL�q�2��l⌵����2+K�2�Hƙ�`�m���E���v�DESc._�aϧ9����wVǕ������QGc���P��X��l���x.Mz�Q�Jz��Q<fl���:X���G&5k�hr�ų:��f���]��D�.Ҷ�ִ��V��f&���^֐�=�!�6ʭ��R�X!�J����d�ъ�R(K��SJ�]ݭ�Ůn7DT�Bp�C�ґ@�S-(M�]�j�F�'/D2콓XB͋��:Sl:��[d�U�ݠ��%.���3o`���T�	�^��mn���*%���B��i���7K��!���k-I�Bj�iO�/��v�F�ή�2��\R�t��+aPGWj6[�,��Զ�F*�E�M�ôַ���u��gɱ}��.)�5ˬl��A�UZ�B��km�Ͷ�ܜ��1�޻�e�U��u�,]��	��\����<�Ĳ��[v�guz�b���V�&��f���CW�͵�*��\ZE�)q v��n�${!mA��b��M7��X,��.�&�Q8����X"ֹ�؛��+v�ĨF�HZ����[�����f��.�n\a�sB�4� �eMf!J5��|��L\�)�+���F����6U2�HE�V�&�ـQM7/��qes���-ѹ ̨�*�l&ó4f�:�;f�Yjӵ�2���!3�V���f�2���Ѱ��#����v6i.��%��6J�	0m��$�������� �Bݵ�#{m�bovʖ�@Q�+uٔqY�6�}�zE�����2۩e9V�I��ѥh�f^ɐ��뵼��&,�0Z�t�1k6��k0J�MaN#U��f�Q��n<{J�g��fa�,nڌImT3�	މ�k��[u��c,����Q�z�i���JY�Bǋ!u�θ��A㾛>��4c4D7[�7(e�j��龫|M�*d��K�`l�ia#Z�u��	yi	`Lդ�XF_��K��[5z��ܳAn��1&&�n`Չ���b�,k�f[#j�aLD��,`}��C�{��fg����y)�{��ff{}�<���'���fg�7���%OwwL��o�� �J#���陙������J#����]u�\{�q	(>z��xp�1P�-_����AP�畢�۪'�ۼ���vz���+.������4�t!��撄�6&�@��+e�@a*�Wn�9�i(�$M���L%K5
�	l.�e�}��'�l����m)S<�3���c.�	at,�P
�f,3avdk7[-���bYf�(i��Z��l��P����uoݦz틄TճI��S�����Bv��!Lm�F���KU:,�Y�t�,It��
��Z���'I=�ͱ�[e�%��� %H�%���r�� YT�#H��=eeK-��z�W��5�t��e���Qꖕ���.
=�uU�H9$x���/V����m���jۜ\�EN;(0\��؄�p�f��t_UTID}nĢp6(0ƕUۮ�e���[^�X�;���� d�k���)6���T�}a.��y����Q6�C� ���i\�Aq��6ؚ��M��!�k�>c����UWr��WTr6�IG!bp���il�;qQQ��[��+����ןy��Q7�z�R�EEZi�x�^�
���B�֛l��i.��h���62`�.a�����L\�[��t�tvv�iU]�AԳVU��~����ג�HVĽ��U�.�k�FȚ8�M��r���}>�UO�D�&Li�Ƴ��>@FEc���J�骓OR%�V��n��o�6�Ǉ�l0ƕU��w~���s �:��)�
�*(�!�S��쓲x���0]D�jY1hWUo-�ܗb[w�F��̰���n�Ҙ�^1�#C�6�Ыۦ�e%kf�ʺh�t�H�6.%��)�Q.�m�QؽݭX�8ܳd��2��a�fmb$&�Y��b%��MnI�x��L�p�7Aʄ�-&�F�T���
㓸��W
��m�֧� �i��z|�iU]��3{�Z�Z�zO%b7K���.[�/B5�V8�#�Mws5s^��ι��>���\[{��B�ƲB����;ݘ8QFG��a�*������V�Ygzm��#��q|]�\"��S���^���X�	���^��vwcU@��E#�w��KL@�ҡ9�S��k���}�����^�B�}�`���&�n4�]@ &LF..��������E�e�����,�4��/�x�O"�	�����e�ʾ��]Ź���m�[����<�s}�m��7��گ��޻m����Bi�$-S���\�������ݖ�d���c���.��|�e��qj�,��OL{e�Kp�jU]PU]*�]e4�4��4i��D������M)����Zǩ�Q��ttn��S7���up�i��2�M�t��t�@�cv/ژ�VS��9�$rw<Y��UAq������O!��=���[x�;�,� �4H�cQ	������c���ڳ2�3׍���v|�XY����zcm�MZ����
֢�┧�Wa�����4����Ēp�t�
i;����mK�ъF�1I3���F_2I��r�u���eguZ�d��1��]E�X�^�3�rߋ�lz�<gNe�.������8�x�c�v����.8��V�-�x��-Ux�*�����Ut�\,���x��Y\d��q�Vߙ��*�>������q����]��{��W��ūū�qX�-_W�W�j�/kⳋ�/�q\zͪ�ϗ�ⶼ_���x�W�
�j�j��.:c�ݼg�e�x��(1���p\��P�N���p�KG���C���΅'��s�.Q��Q<HN���]��4|���.'6�uq��3My�϶�~�_y���o*��9>qNk%rp��vr�s-f7���q��_�?����)����`F����C��> .#�}�L�����G���fg�ww��@�{��ffxgw �@<;��ffxgwx%x.����J �����x���i��Ǌ�FM[�^:u���断Z�l�U%�,�oz�ڭ"�j,J��cqA��OV5�-�w�n<�-&�>Y�����h��Q@[fu5�U��^�[`�pޭb�UB�08[]��&�%�ٱ
*�H	Z'�=Sz0�;6@^�ja5�!�'�U���1�*�4�K$W��d��&Ktvz�Xi�����__{n3Zk���]�Y�*իV�,d��LW��$e��$b\�Y�)�:�2fg��Lm�U�@!!w"X�@�d��4C&���u�`�������wF�jP��O�ˌ�~���2��_1tDlѫ�9N��w�S�q�u'X�M�=r�؛�B>.Rh��R����W�Q4"H\U�8��kw���V�u����D�����ţ5�g @�����2��B�T��M�iLA۱�1 ��Q��^�5�Υ�]�uȄ4W@���	�Bj4m	����)�f�$4�'����tΎ�U�k�kܗ2����JL��]D}�)�/1p�N&JA�DxE}�����s����"�"p�bx�e"�+����)$V���E�Ȕ�_�1>��5+Ne���5%?6��`(�k��0O���<jc�G�6�4ӣӏ�����Ǌ�kb�5�ЀU�Y�#�� R#� 8,��4DnY�&͚�j?��!�PX��Y��:I#�B�<h �8�����븑��߫!j�+���V��q�YD�(��ccʤ�0&��$�����܁
<�0if�c��M�~Y�<�����֕Z��a4'H%��m�6j��0D��y%��K��{[�x�H��.\V�d�K�{XH�E�+1Zc�/��U�^d�jիQ����N��ڪ��,Y��<�+����;��UZ7t��L�ItIL1%�f/9����4Kj��5<O�*Ε횕'����c�3f��g��X �@m٫(\�T�_+Vc������������)p�d�j�J�� ���/�s���iٳ��a�+Ltc�|�Y���Z��D��v�oRI������l>�&ר�l�L�2Q��������x:K*hUچ�A�Q�(�*��%��^���������.J�O0]WMD�����YcJ����F0�� �n�ے�f�n@)�R��.r�dc�#�7�v5��)�%S��o2w$�t;y���Xz��Y�8��Y�֟4ӣÏ���1я<|����Y�|;��K�����גv�I9�q�qF�`C��BV=l[|����^�OliT�o��1��We	�m
m+�5AKw4�U����Ё�����t�K>�q�O�u�j� X|�	ԃ���H��I�#�j��ip�M �A�Y�d"�zU1�t�H3��	��=�<�P��l�p64/�c<��zǺZ�OD��Ѝ؋�{c2 A���s2-K���l���lѦ�ٳBp���,X�d��Xi�1��<m�\�Y��+]���U�U#h�d���S����07c裵�Ǎj]��̙��]��-D�(��&�D���D㲇o}�T�wI�>`�$�"e�f&
�;ry�7c�5���u͛���+�,��s�8� ��0c���&B�I)<�u ��,K1M�d��W�&�6���t��?:������1'Vw,mƘ�����aZi�ti��,�dnY&�՚���j�H�z��S=���R7,F��#�&����g&i<RPf> �H�	�Ò
d�*�Z��1InI""F���q	(a�	H��pҘ"_x�]�N=#!��X�# ��D��/�n��3��.64Y,��0�la�B�P7��o{�hЖ�l��>tҮ�2',?<~c�G��+
�Lc�L��P-j-#XQ�JM16D���i�vA$w�/�,�KZz�'dB��j�%�ӂ�J:[�)�HDz\�7$,��r���8M%Sn5�R"i�d�h>�!JZM�,�6�CQ�F�gYHI�����b9Lr��I�:�ц{$%���K莓I�����
��	��%(�:x���-���k�g�3��1Ƙ��\Z�/+^1ƻq��/�3K����[W��r�W��⸵x�\^�WKUū?-i�U^*�Ìg��x�+��Ǻ�c��l��[gj�t��^-W%��W�m�'x���UW�W�j��L�_�1�/k�g�j���qf׋�^:m���UºZ�Z�S���2)���`\���XZ8.�Â5�E��s�\5h�gck�������x��q��iƂ@�7�Nő��E"��f��d;�z�A���0v��`@�P	����ueE�12�<��j!F�Ʒ��S՗5І���(��D�g��9��>HR���U蹌D�6��DĘͪ����
����J+fA�=�6�̍�$me��XM�	U6������v�~��C�$(
��S�K��������	��|���K���}���>u�6���R4���N�&O�����tf:���g���D�ݕUU�{�	D�ݕUU�{�Q�wweUUp�ȦxwwvUUW|�D��9UUßm�4 āa|���Q4�J.b��9�X:T[���6�M0�n�b��B�vH�H1�fX޲ۨ$٩���
��~}�Kp�EeaB���uvȒك^&��MpU2�+��2��L��X[��V�v3�Q�RĲ��hfY�m�P���a6v�0�n.yh�6�	qu�ph�n��:8��]�2nl�S�v��d���Z[l�M�!Ȝ�ZG{�{�kh��a%��[j���b�6�Y�2�@��150�r��/Xv�����L>,��e�Y`jٵ��{C����p�6�qև�N��3[��pz�ã���b$,�Lo;Oa�.l�o�Cz���4d��L_B���:`Pv��[�hi��gs��P�侰�5Lϓ`X3Mm�P�*�[i�:�T�TUa�sc��M`��.�&@�q�f�T,l�ݰ&�r�^b\M(��8�W��0�����rZ���U)�l�Jj��
Le�@�z�5��O�coN�+
�LMT�����6^ɮ��P�K|�h�n�ӎ�8�!XY���{R�T��,�e��4x�,�����<t�7��W F�g[��{֒� �VN���ƓI~��)���VEdP�b����j#����� <橏�2�;�����G�%��引�&���\����7>q{�f��κ|���so���gǏ�i�1ѧ��:$�f9�@����K�bܘ����&�J�񤧏���3�y� ݄ɑ��������3���Em������\����A�.x�a� ƙ�(S\�/�3��2���ҘD�aX0�=s	�,2i�l|����aZi�ti���� _����NkȮ���f.y8�O%�r!=��B���;p^\�gX�M�%"�&:�K�J��Hz/�[�6�J,<V6Q�H[Č���$�J9R\��0�����I�t6�B>{URYv�CF�%� [�Z� +�;�*�/8�l�t�yӹӑ~~z��8�XV�bj��o��cmT1F�P��z�����cCt ı:hƶ�k�*i��X껚Ra�4�aB�\�PbF�,�Yx�1�A�]���ʘа��S�}>�/�N)b��;#��7.�կ��D6�d B�=U��CIb�N1.��k�,� u�T�T�[���b�����R��u�V@�m�����"�	qq�☢K� W�@//��nm�,�o~�z����+
�&��E���O�^�m���Z�=- V�:�@,|x�mS�^JڱY
�U�h{����:���1|ҝ��J���>w!i.a^�u�l�L�ߞ쁧V#�,�.Y�>�Iz�~���A��J�B�vRe0��{��[]6����^�ɦ�L%RN��׽�3���F7?1���v��<x�+��O���OH�d���S5$�u44�\���X��"�#��s�/��K����Tp�T5)�)R�B��Y	ŝIS��x� y�����_ŌO,��DyA]��%� X�>����������ˋ������i)�dZ���O_N�c�gn�~q����aX����;�MC�6	�IĚ���/��"��H������0Ưx^Zp�Q���PaUc��O�������@�Ɖ�*���!|�%=a�7z]эI'��%���/$��a'��!c �FƋ4���Jt]�f��t���ⰬV��<z��κ:�ޠϾ_l���0�J���������}IM�5��+K�3�
�-�lQ�(	�VUw.�m+%4UE�:�gE*�EiHGM��#�L�e��jJ�u-��f
�m�����R�vI#j]3�2���~��R�Dl�_J|�6�9$��RF%�g�-�S��LU%>_gz�$�"�v���ʪ$���z�!���G��x�����g�±Z:4�������:v��_4��73�]/zӹ��w�oZ-�V��g���~KB�xW
��.�����`���K�cbaj�<�IW���L�H�L�r�(�/�K@X�L�$�3|��x�n�\7�<�㔧&K(X���*���x�/O��=���\g�c�3���i���������q�q{,��\i����W��Ҫ���-^-V����Uū?-��WL⫌8�q\^���q���q�]���|�z�K���e��qj�m�d�U��昺!�M(�0O��<GƊ�+�����x����̶��-W�ij�j�N+�ӌq|z毬��и4t!���X<Z��V4.��8Ŏ<Z9G���:WM3�[��5���W��-��b��?Q*6�[Bh��z�"���q��hge����B�S:MOccPs}�B)u�]�D����1e8$���������W�N<ʮ���L@ė.�qƳ�]:]�gx�-׉r�Y�n/[�7�\���ڵ��p��TIn�[�� ~�*��?�*�����wwNUUp�ȭ<;��r���>Ei���ӕU\9�+O���ϑZxwwt�UW}���,��BhQT!E��]�� ܉��	�f����0�8��@�.��\ɴ�zM6z�J��2IEZ���FJ(���:uﲖ"@&^&-x͡3�����ZG\�=�T�7��ɧ����]��3h�z���|�w99�6����aTB��B�L𖡆4x��I.�-�v�X�n`�a��̀�oA����ZD#l(&�mH8�o!��ެ��=��Sm�Z��\��+~��R�C��'s�=m��N��{����b�.�ɤt����p�UѠ2��`�:v�*UL&5�)��l�ѓ��#׊±Zt���_5z-�{YOt����GC�?�=(�j�p׎�����n��S�h���(�I����bhT���Fm	�����
�+,�=��_�q�gL���$*[���7G�&\4�0�ľ��	B����9s��!$&S#�9o���"�����r>�ۍ5$L�p+�S��L�QR���^�����1�{վO#�?4��Ǌ±Zt�����������j'Tʵ2��?Re����J2#�F��N��9>����#S��X�{rX3	&�72�:�����$�	�W1%�jJ}��l`� ���7İ
fҔ��,"7�����kHK��0T�h�� P�_��,Q�^.5wBX�[�':ܠ�1���6�[�3ܝ�MQ�|�޲����T��yd�IkQs�͉�97o8j�w]\c�u9�����v>q�Wjk_�^tzx��<���M���5��j�fr�拫�k2#;x��[<��|\���*���5��+�7VjZ%��u[�d�9�VV��zv�Is�@�3)	89s�J1��x��O1s_�t09�醶��:N�����E�0�!A
!cd!c%hs�-Dʧ���|�L�k4�1���(�h��	L�rM'�G��.�
.��sE�P�^(�J�B�[��G%�� 	��SsQ�����,x��]0�$�\���s�XK�	�]<��n�Qӝ�o���S׮��>h��ڦ��_!
./�~�d^V��6;�V-b���	�����8�L`T��7dl����In1T�_k�3�Χ2����-�;L������;=���Ŀ��<L�/䳓)��gn�Z0�\�q�O��O`�M�C;(�s��C8rA�Re��I��:d���ڰ�V����]�z�\��l���o.���e�&A,JJ��J�5��M�U6�f�Ϊ�$dy7ce6I��j�jY�6.����[pB�M�j[��y`��Ɯ_u���a��Me\�r8���	����ag��D0�1	~I&R=����tܹr�W�h�Ƭ�㻦��v���Z�����J����'�>N�;��܄�XAهTH�䐑�H��D  Y�8�>�Vq}2<1�?i��i�fw?8�GgnՀ���
./�>��G��b �,��%:����=/��ŬQTX��j������od0���K�}4�4��{;�_m�{69��T��f�S��`y�F��7��.+�9#�J	Dle��)b�gs��'�>vtz�XV+��Zx������2�۴��Rq(S�nyw�!�-��G������n�}���G���D��:�;"�A���N^vU�;h��������Z�hL�4�u)��H�Qp4��{�5Icȯ�Ox���ڰ�V�*��\얁o�/�U�l�̦��BeǅxʪH��^�h������\%ה����yoN�]�= �g�`4g{����9V��6�O�L�.�+�K�cCI���>7��J�}~g3��}_\��]����Ε�3�3����W��/���4�����\^+�������*�eV�W���ګL�v���U�V�e�x��_�Lq\^���q�+�⸻q�.��;f�@� G�#�B<�Dy����Hh���.L�+��<C���U�q��cj��9m�q̶�f/��������,���x�<^[�papa0Ѡ�0��аJ&����q-	�	�������"���/"Q+ʔ�y'���6�^0�vM�Y�B����W'0�-��x�T��?n�K���������(����\%�qY�״ݘ֙,-ـA�(7:栯I�U
����Q���˳o9���n���d��[*݊��tk��s�o�O/]fF���/����o/��z�8x8��D{��Z�m����(!ۊUb����.PIE4:���sw�\��/o���{��r��wrKq��ʪ���,=ǻ��*��w$���Ꜫ�ܒ��{��r��v
,@�H �����5yҀ�V��
b�9��^M=�tɽ�c�k��`�o�3�]n+j]���B��f�!�K�.�t�m�-4�Z�5�hH1k,j��cIsn;a@@�U
��_%|x�I�\�Z�K%(X�i��F��Us��J�c�ޡ|M���+��IS:�B�� �p֎��r�M50^�X�Q�p�&+][Hk���a������b�Z{��MJ�M�B��!Z������e�T��J�X����!�U�*��Hגdr*�a�X��k�%�q�3�ՠl��!6in�]�BV�T]�`��L�o=k�JR,��S���(-z}�� �]���URV�ƀ�i��X�B�S�N7����2e���ON7}˒H^&K� ���Io;�G"�Nڠ�]-N<rެ�:ʑ0�m�M�F�,�!@&�ĪQqo�����;�n�KԱqY.�S�.p���,���6�pL'�a89N&��ٰ�I$���-��	�uAw
����lh
���jI���@ߣE�]Kɤ�$����n+�$��q���rK�ӹ7U��ŭf��&o������cæ�1�?=�0�%I����&��T@����7�<J$���p�WJy�7�����'��=�qE�Ma�� 1�~���ێ�+sW1/�_&�8&�.�$�MP��׈p�;�;���2�Ɣ�!r餤䐙C&{�ϞWN��;a�W�M<c��;֤���'�eKM��I	����nj�ǣ��Ff�	��C�4�Ô�b���H2u͊M�1)ϰV�+��28*���x�@�t���s<�/{ڪ׽�x�/�<s@Y�z�ⴜ��8va�\#Ny�æ���`H�asz�!+<��T�q���d�8�3�(��RJ�A7���ׯ�V�r���f����9��{�o,���P�F�-�rżRE�>Z��j�:e��d������5!=�ɶ��RO�_M%�{
-6N&
e�cE<��h,ޝ<L�.�2�l�ˋ������ȜBꘌ��J�#��z�(�&ˍ�����v-�]�#3����q�7�ٖܽ�=t��۶@�"����}�UU3%	Jt 3Ć���b�#%9=��
a��}�T�'��,�7�۝\����Ïc:��K���s�^���~��6�ged�*����/	]Kz�)�kį4K�]�f�<�_�gj��G%%=]�xw�܁#��fEWJ�թ��B�����^xrdbQ1�H��M���eI1z���*�Ha\��	|!E�y���{3__�@g˥R1�e�n�i�㉘܋y���.���R�ad��J�T@Ӝ��kNL�h�>��0��<W`I�K7olf��մU�s��s���m<���6
r��S*���I<�ӳɤ����o����+�V<v���81��1L�Q2���o��)y1j��P�4CNWT_��c��j6��n���-ʔT������.���L�m<�l�,]����q4�L����4b�3UTUWŊ�	gZ�5nJ��-xi.\�s�2$4l����b�Uc�o�̼ű��_;
8*5�"r�W��dU�/*F^$*D̛TB�$��`ΐr�:�t!���2#���M�r�t��/]�����jι�1��AWmQ7J채N�Aw8�M{�W

*�.��{Y*I	�t�e;:��)f�z]��>27�S)AQ�Y�g�m��_2r�:��ˎ41���c�уNw�g���'�ь����d,x�`�p�A�V�X��n�ֱn.Yo��ӭKQAIԜ����Wo'22���{I�õ�ˣ���s�m�SD+��Y4�M��Í�6�i�-+��U�*��t��-�ǪZ̎S�5�g�wIƃ>'�8�����c!8Hx���L�x�����ͼ�z~gLc�e^4�q�\/�3�����z^+�1�U�6��b�׵�mU[Z��b����W�V1�m��j�U^+��N58���v�W�\q\]�q�x�8��E�ūūūŕ�������1W�x�~Y�z_���?1�~x��qv�W��v�4歫ū��UW�W�8����y}q��e�|�oW�����^���8�-q�8�z��6\d�LpLA9!D��@=�8)��Ԍ+PUy��}(���yFi���{�N닭�(4� P2.�P�|��5`�7�wE��ʟ����_+�$�w
��S#Ư}��D.��ɋ�>b$���/��.�]���H�ж҃�o7�r��ܒ��˻��*�wrJ�w.����+=ܻ��r��w%q�˻��*�wrWܻ��r�����ƍ�v������x�}�W%B��8m>���\&��ᴺ��7��ԕ߂I޾x�t��X5�^7��7��������,P�2�J=�.p����y��Np�Pu]����[�Me�`���&�%𥉉z:�w������;6�1^��a�t�!L�ٗ3�V2~ ��^�}��k*Z����K�3�S�H� 7"(����F�/��s��%�D�.��xB\�i�L�!�&zMg6î�zH�o��l�􄄅�_���K<�t�S�Xhx�V�0��٤�B���.C��,�{�� #�t�I�ӂw^�rm�>�o�%oM����b�M�k���e0�WhZ�k�"j�%�i�Ţ��4�8:�c.��,�Yq�,o1Q8���m��.�~/*ʗnu��UUX&=�/����B�<(�#��%7�qx�#�SnM���ڪÈ�<�z]�P��I!�n�2��;�4�9h��	�"�[�ː.�|y�Ӈ�.C'�LQ��5^�EV�4�:K��9������Id�A�ϺjT��t�W/�Տ����%����8�C�2�O)^�z/�A&e�=���?,���/73�$���u�BgڔM%ú�����k���$�e�̕�/	��%�|=
N&<MZ����,/�#��<�?0�����+�M�;K>o��CF	4
��ݦ�^���À�d��!	`�{��߰��4HJ�!C����gn�`�p�wg�<Rt��e�K�����\]W�M|�r�-�ωZ�b��,��Ƿ4\t�=$!t��=�W6M:n��x�Lq�g�+�|�Ǌ���g���Zk��-c@J����~8$pr鄸z�#�Dڊ#�<2��U����S��:�!l���e3�t�ƛ90���/L؄��n%i�ø�|�r�2E�$�̜�Wrl��0 C^�	�/�o���L�]h�u�t�t���H�m��}I.PWZ���#B�Q5x��l9%FY6!��Y�q*v�F����Xi�[�nN�ո�l�җ�J�ml�YM���o�W��Y魹�4�|��1�����B�S�m���=�����i�m$-��\-`� �qIe8�qNd�[�Ӷ���K�ֶº�
��#�	��w����ˉN�Gn���ܳ�ϟ���+�z��_+&�cW�%��g2����K��X ��㎞���I��)�=n������ET�����}����3�>�>��|mc�=���	UV�i�y�)�&-�ISFO��)�ڕڼUc�>�Z��� *��Μ�.e�y$�=��y~ %��ۿ��Y(v��ębu��s�����#�E�%Þ�d��-|�X�G)�\�.��$�c�&
r�M&0���Bk��hY�D��N"�Գ�6㣥:=R�W��x�n�!�a�&J���M�p�h۪"���-�\8m�lJ�w S��y7��`�ɾ�wwİS��l.�ģ-��y��:K΅��+���I��e.Git�^��8p'�	k��b>R������#V0��t�#KW�4֜e^ūÌ����qx�Y���v����j�U[Z���|c1j�Ug�.���V�1W����x�׊�������_��?e�W���q\-^-\q�x��2Wx����v���1�L���ҿ/���������qv�W���X�[W�W��ūm�-�d��.�g���s-q�;|�-q���n�5뼾3�r�/����xap!��1�0xhX9`�PR8(��G@(���0Z�ݨ��Rb;���rp�~�����q��_K�5�6p�y:v3�\�j�h�������Ғ"6��1	�9�v�
�V
ٱe�Tb��	�������7/r��'��*�KưRۨVL�b�ԶR6���I��4�n�.�&�5C�e�3��x6�;"���=�"NEJ��ۛ��W��꼯�E�Q�v:��٩R����S�\;�+]���UYUø����U9\;�*]���3�9r�K��:fb��ʗwtt����b��@`4$-B�Mq\b=�?+)%��L֔5�KMf������gOa@�E��[u�+e���#
����6Lڌ�����,[R��e�õ�7f�&���Y�-Ò� 6:Yu�C]��B$6��dp�k@֢kGRk[��Um�K�:�Cҗ8�kw4ct���[ B���96�ڙ��e-ΆH�&� (�)L���V�"�T.=��{y�%2CM�R��R��k^-��6��ĶVZ���Lh�1M�M�V7:�^��$�At$jM �QX��a�����b�$�\�XݠU�I��cq`;�̈́�B;F1�,�j�i�P�1z���-���t��n��̡�B�ݘ4�3�Q{���ɩe<h68xY^�Q�*�b���0%�y ��q?�̲a�*�j!M��G���C�R>7z4Pڝ��]�j�x�<���c餺pq/j
����p��a-�>�r����b��S�.\.�ӳM��[�R�`��4�A&���[�-���i9c��sVoL�t�W�CɾGo�ҝ�)]��V<u���l��4��b��^\_���cS00�tRy��Ɍ�6��D�0�L%����d�HGL5�����uMZ��������^�&�.� "����FpĹ�[�wL���%����HZ���⾯N����[-yP*ŭi�|����ҝ��e.g�3и�\\�@u�&6�&�M�a�w.�M���5���@�s�a��s���tэ�g@����!��F���Z�P�]��*mb�q:��n�*xx�v��x�ޗ9|�U�V�]>��Q�B�}Y������L4�"��ʺ Tҭ�%�K�4&�]��d!\,z�E�R�6���A�!F��j(+*l@
�$�*@�uɷI�����$7�BM��l�M�N^�Nl�UJ�p�ZK�J,�"`�s�s[�5�U�rĕ{N�˖�$���7�M��JM����1���鄒Tԍ8�����q�Ț9!�<xٓF9�!�J2t�ȶO9,a����D�}PBT(��`ƶ[)�L$/F�oAr]���{�Y���!^}�(��3)O�����7J�ci�UU�0?b�y1e�h��ܐ�Gt�j����)��H<c�J��)]��5׽b�(�2,<K���V䝪%��,B7J�j ^���_�Mn	&�OD���
�E����іD�U}�1�3��ҁ�I֞�i��hT�2����ɫ�S�|MPv+.`��ْ�I�(���>=�Gwf�-���d�+�ӝ���W��+3*��Ң����s�l�dh���ѣY[�YTe���'*�����H����0aճdU���m��#�iJ�ڙ4m^�#`Q��U���qœW�t<�@��S-L�Z�VuH�5�#(�a5]XeMX�5iPI+[
�!��#�d�@A*1��K�L��H�D�nGD��-9���قd�-��q&�܍�4����Kb�,q1+����V��i�>P��\Ff����@���`�d�]�6�����sDH�%2� Ȥ�"�."�X?YU��[b%�vYNJ�55u/��T�Sq[@- ��g9�	�oBn�üK!H�8B��A�朦��)�,�KUZ����#�X���)8M�wI���6��#�ǌHC�o[��v��L�lZA��>�UTWn���v��x���+�<c��f��4��4u�D;k��V����U�n��q��.u�[@u���]
���v�t��aY��cηJMƛ; $���t�wۧ�|�{��b�	�����f��S3��+�<@G�ͤpJ�Ya��ı�HNߘ�kKr٧�\���g��.2g<�w�$��&9��+Ȍ�S�������Nͩ]��=���u����J��U�.%=#$�`p��a�!�eUJ%�s�ec�'�SԺq9����s�VU�����o����g�
plFT�3�O?a-�2~Q/Ǐ��i��׎;|�m�l�Jٳf�m��V�q�|x�_���i[6ڶ��ݱ��m�m�ͽvێ��¸q�����ӧ�q�N8��{W��m��+fͦͪ��lm�M�z�oZz�o�i���;m��6���1�;m�o�>v۶�h��l�E:W�v-�UN�q�&1Q��XD�t@�f��,�,P^���"�\ q\1Y
�!a�7R�ő��jZ jn^Ȗ��8@� !n`�k��Q�c�w��`���L��(���p����f!�#�f��bT�i��=;�K�:1b�g�b��,�(2V�z<z�I �#�}�)#w3��ޕ���L^T��]��|U�$����ʸ�j?��P�v���[��yR�����yR��陙���yR��陙���yR��陙���˔.���c `1 d�/S ��DpO���k�!p���:0�"m�D�
3� ^�/z1J�Gk�KCLk��;���K&Ε�0X�xy)�ӆ�	E�$rV�/;;�RJ#�]J7�e�c���T��U�3���*��z�*���&��Y�=cXL��/$!N�����AIGH9���/�q�%�]�c��y�Yݒ�Gd!��S��A�9���O�#b���+y6C/Znm�F3IR���9|d�v�:q���J�U^1�o{�翺���w���T�[#��Nw�����,��G㑫-�Z�q��qZ)D�v�ZE4���mf��uڒ��Z�S
T�B�Mؔ_q6��:�,Q�9����G
$��1t���\<v��%��Mq�$'S�I�=������Նdՙ���4�(�<Y�~����ZkwK�p�0C&K���ڪ�cƺ��w|'��ߎ��hc��v��wc�.w#M���}�N���}ͅ�5�ѱ��#	��Q]y�h�a��:z���UEXp��Î����V��Ŭ��WԚ,i�,D��X���\�P�L�֓lK�����Ӧ�楦�q�o�<v;=R�B�����R�V�o�e��"#Ȏ�TJ2�05�%9,L$j��d�w�y�uF��6:�6���^��2�$���z��3�v�Y٧�$��S���gGJ�ճ��x�vj�X��۔�N��R�[ ��UR�tgŒ�d���.�:ݢ�����5�H�$6�1���'	�٦<}�L����CVr�,�Ƥ�/
r`0���o�)��U:n����:��6���ڕڪ�cɷ|��M/T�I@z66�9�"�ՊOj��!k���Z�i2��KF(�Zh�g�-W��7uU�0��<�LV"8^�֢�*�Ӓ15�����v̥��{~.\�t���QT�Ad�t�qڸ�.��ҍ{QCo�"�aQ#��ȼ��.��h<>m��)mQ[#)�i,�ź�]8�/�ə	v볦L���U�?:ˎoWX�?M���k&���^�:H�l�L��b��$�IP��l%�'Znh�I����R�c�[P�R���)��[��n`�˝�9ٙ$�N.)���]aFL��ڕڪ�cƟ^��W���{�g�}�UT�#r͋X��r�P�vi8��>�Σܐh 7�OM��&
L��5�[6��{��׹�)��hWS.�v�#���)�ݒHg�K�ѷ)]���<a�d��y��!x��`�IF8N9.�ɴ�����x�<�~�/�2��i�4���\��r�D)޶0m|�&y�ȋ�V��'��M�M�J���Τt�h��B��sOy�pԖ*���є��iפ=�:<8�jt+O�8Ǎ�x�׍�|�m���f�6m���m�i������ä���fΛm[m�nշm����6��m+f͛iU��Ǉ��N����v�>q�6�獴��>M�V��m6ۦݶ���z�o�i���;m��6���6���6����m�M����c����%�;��E�@j���+f���9T*��!G*�al�bbkJsث��vlSq��z_B�)}�D¸�V�P��R�ē�l!*�H@�34jPD��w�KP�(-�1	�e���Tjcr����n��&(��/��} �h� O�<���+�{�|�Su��"Dl^>�Ǽ8O6&�M@Q�����/��_+��33?gø����33�ø�����33�ø�����33�ø�����33�ø�����33�í�ׯͩ]���<#�������2PaiF&/�k�wT�^�9��C��tE�vvKu��HJglM�^׆Qp��Ź�RB��4�m�%5�r�c5���k�����d�駩+,���6hVj�����ؚQ��V��צ���ͨ��
��M��Ԧͅ�T��`%�ڊ�+u��my��M�cZ3����T�]�CB��a��70%���>��Jrk.%Vf�����v%�B�����5	
[�,Ŗ��Y,q��ٖ���T��ae	��]aQ���'<z���
v�)���R�7:͝f)�CU����R-8��h5UU��$eB#�Fڱ�k9���gP��d�-�j�]�`ۤ��D�RY.�6H�3��?g��^#=��Z�M�H5!4U�Wk��9
PQԘ�/L�r�~�T���>v�vx�v���qׄ���i忒�:t�~���ų
�#�s^�nf�V�&����Ƌ�4p��5�%�f�b�Je<M���l�v�/N����:�4��C��+�U\MqX�n�� е,�#2��}�@���{�[d�Ɂ�cVK���ZZ�5�b��]R���7@0^sͷ�Xw0����=oX�cvy�$!xe�Ļ�'[̴��K:l�& ��J�U^1��fW.[X���;�i-Í�."wfMr��0�Q`�ZT��$�>�k��|��G�v;E4#�`��U�l%�T2Y�Թd�g;�/ĺeѧ��iҒ�n�q����lԄ��\coGg�Wj��}�}w����e�/e��UU�\�*Ǉ�����*4:^��D-Yj9��8t	t�1��W��F��v���v��b�.�V6;��LD�
jT�R�I�>K�K2䱧��,ݻ��7���z{�SwI��t�,a#@p��QQ��[A�����UP�;&hV��i�K'[|��i����}�Ui�m��R�UW�}��	��쪅URm).i�a݊i��M[����S�9�Ncv��Ib>4���)��sV> O$�4�LB$Tw~:�ٗ��%2����ыK��U�[�QZ�>i�=�)]�d�9��X�cF��\͓fwEUe.Y6�i����bk�mҊ����흲���LvT'U�/qj��EW���T��I���O8x��nZ��ܛ���㻤޵d�A��-}��Tt&et�4�lD��Ѯ�d�X�Ҏ��)]���5�{sS+X���u��jU���k[�%&�iMА�c��72 � �T/���{��
�����p_���bo��3|��6�4�6g��_�oj$��S���m���?j;�n;O81�m�<���P�5+����1�.n\����I�L��N��.��I���P1�1i�X�#�mFV�ݶ���[S��0B�͐lͥ��5&�k���n�ёX:Հ��ּ��|]4X�G�$�	qӔ�[[	�.N&9$�0�v�Ka���&���۩���Ȏ�Z���lل!���i�a:ٲwf�HHBgΘ�o���Wj���d�=�MF�#)�v�����tݜ%�=y9��D�Z����3�^���KC������k� B�U}Sܿ��u��KN�J�"u���V��~�{�w�{��=v��J%B�d�N���1�$��Tu�J���^�|��o^��붜i�+lV͛6�6�N�6ۇΕ������I�Æ͛m�6�m۳om�m�m��V͛6mѶ;q^;Wk��N8㏜c����W�Um�cm�m�M�m���[m�lx�M�����t���6��ϛ|��m�i��b�k.��뙓p.ʧj����,��vj�]���Pb�$=PNҙJ�Ě��eT�f���D��D��w�nn���˽քHA&���43Ff�m�33/9�{��ff{9�{��ff{9�{��ff{9�{��ff{9�{��fg�{̼�׏XǮ�j��]��Ǻ���r]!��*�pd��p�幹)�Ow�b�Fk�	���PC�����ٛ���-B�T�bv>��}����ue�?Pt��ƴ��q������v��J�UYHC �C�t�1ĺY��2Z��*����n'������1J*OD闤,cG�d2�N&\nСHF�g�i�x�p�b��=b=ޡ����盝X���oo��M1���/��B�rzпG�6���N�mv�i�B�7V��Բ��لq��(3M��#i.t.lU��m�-tR:�1#��J�YZc��M�K�\2ӥ�q��S�hl�\��!sMK����R�-̦L��Y1y	�&�=�lM�9祏h�|y��a8ʳ��7s>7����K<���AG"M�sh�qU�>��c�1����ޟ)^)]��M��G	�W�\䌔;LB{�Z�uL�� B;�Ƹ����8�3P>���CR�V���3qkW����^�w��5Ox	J����L��h�*{8d�zɾ�6���hý~�a��2�z�vx�x�t�q�㚰��9<J6�B�v��,������O��NI�����U4FZ�h@�MĲCvl���x69��$g껊+�f*�<��{�����<q��;c*�l+�Uv��<�J6�<i��Mn�8����&�jB)D�59As:�#2!?�|�|�$�Y��؞sp3:y��i*�#���ܖۼ�[.���t�8`����SM&����u�T,��~���P�{�3��wSkĳxUʹt��R��]\0���k�K��m���Yp%��[���Ĺ��te���qA�\�Ip6� I��Bň^�Es�v㴣�:L�CP�{��ÚM�$/Bp�:�< ���RDR����.��/��@�H�4`�P2g~��d|�m|����1Ҫ�k�
�(��q)$M�$L�>e8�N1+r�	$��)��v��,]��fss�>�6�VzJ�e6��RC[�4W&8襑8�μ��G�5�������w�b9������(�M5Ī]M*
.B�cצ����n.a"u=�/W�W@�P�0nX�(�c n-�J8�����0<��}�M&�v�m=�/]�΋�p�=��S��e2x�����1Ҫ�^��O�Ǜ�2�К>�p\�w=��Lhj)�R��r8�s��gq��U�W�S&/`�llbi\'}p��&1uZ�Q�nY+�펖2�?h?�?���A��I>�$�I$��UTID?1����@��C�)o��ݓM-Wʈz�"Db�,O�����,�����V*�b�{�@�$�X�"�)�%"�"�R,�R(*JRLARPT��RX�IPRXE�X0X(�EkXF�TTPQbRRX��D�d�$�Q(�Q`��Qd(��P��QE�`��Q`Q`QHQHQd�I(�J��)"QD��%!E�QHQQY$�����b�"�QbJ,��QbJ(�*j��d��R1!E�E�QDQdQQY$��(�
IAEDQd��QdT��EHQREAI,
,�����RJ,XŕcL`�2��4ŚYW�ť�I,�eQeQh�B���P��(�E�X��,RJ��FE�YE�,��Ie(��Z,P�X��$���X�eKYB���Т�X��,Qe(���Qh���eQe$��YE��Qb��X��Qb�(��X��Qb�)%�,��P�E�YE�X�����(��YE�(����YE�X��Qb��QE���P�E�YE�X��(�,Qb�(�E�X��Qi%�X��,Qb�YE��(�I*P��(�E�,T������*YR�%�*T�RʕR��eQe(��YE�YE��(��(�E�YE�(��(��YE�,��Qb�(�X#IB�,��QeQb��E��E�,�eH1 ��`ă1 1�K,�EK�K�E��D��)e(����)b�)e�R�X��X����)%�X��K��)e,RK)E,��YE�X�Y��)R�K)e,Qb�e,���)b�R�,�XeHdR�YK�KYK��Z-(��YK)%�ZYE)b�KK)%�-Z-���J�YD�YKE���JYD����K(,QT�Ib�)b�X�R�,R�b�)b�)%��R�e*�KX�Z���)b�K�J��(�Y(�J��,R�b�D�J�,R�Kd���b���U�b�VR�H�R���R�Y)b�UX�U*�,U*ʪ�eR����R�UYUR*����Z�b�V)b�JX�ZY,2�*E�)�"�%"�
E#S$�!a%ARXE"�(ְ��XJE%"�H�B�D�X�"�)"�,5RgxFD)I)HR*IH�JED�X��d�"���#���?���د�.4%	����>p����(�#���H& Cѯ�b�����������M��o�|�~�������}f;���c����f����Fa��8J?��~	������\��~(֏��S����R�,��_n�S��EU�����^�`~����?G���E �P���X"���hS,���'��_�?�}�x�������������=�~w�����ȇ� ?�"��ϭO���}�Ұ�>�����O�v-B�
��Mh��II����׊4�5�g;�P>�:�/�Rf;�[.�Ĵ��'�~mO�[��?Dm��� ʊQ,��
��D���b"#�Te���(( 4]��!M3S�7�So����\=����q��E� ��ERI�	$��ʈ����"�����D��'��8}�[��hx�1�?��~G9>��P�x��+�a��_�C����_��?Wؐ"��%'���Y~��@�Y������ߕ�?w�c��.��ܜA����������0�&�	�π���@?�诛�����~�G�P�qTO�~�q��Y��_��? s����!� � �����EU�x�_�~&?���h��}���|�ɲ�\>)�;X��?�(TP�Z��ÿ�n��Հ���~"� � @`X?��`\C�%��)(���4?o��&���ި��m@�d��\'��'c�A?�x  )J`��?��pF}}���*����0�"��I��W�j������_������>'��W�0��]�}���
O�~����3���$D��������~���K���|�C���'�/���0��&���A���?�-�G~���J|�������o�q�� �H���@����7.A�z��.�� �xCj�?��������_��ģ��c�n� �m����TL��H����$�Q?b|Ϙ?1�%-����a���?���6�>�}�E���рȥ�����M�|������>� AA@.�?X�耟Pn	��Р�0��ҡ˿����������>�\��߁����?�*�0����N�.�p� Zc�p