BZh91AY&SY�(����߀@q����� ����bB�|      �k&�"T��l�U���f�Zi������%l҉ �m�*�Ul��BKkM2*��(�QJֶ5Z���i�ي*kT֦�>�-��em��[iXmUeE��j���-����5U&���0�Z�*AkL�cɐ���b��jSZ�-�f�(PP���в�����d͵mmm��۶(6�d�g �v�Vli��+R���mjƛ+#km�KY�&��T��VKhZ�1%IV��-��6�55Cm,j�o7vm��VkUjx   h���V�b�r.�Vv�u�A��:�kR�]�����c;�mf��ٗu�m:;,�Z�v�n'JI+��c\�-�.�fV�R&֭��fm0-o   ^�� ;��P 7;7   wrp�4:��\t �-Ӏ�@L�  48���z z��PN�`��4��)�J�hZ!�6������  ��zPt�x{� �����(��ˀ�@�]� ���q��@�/.� h}��j��  Wp ��XUT�Ql��T�2����  -�
��8�xhtz:;^�zz�]���� =]�8 �����P=���z7� ��� ��\4  ��6����6-f�!m`��x �x  e`)��qg@�����()Dܸ �ۍ�A�:t�84A]»�� :YE��3�P ���j,��!mcmm6�d�a� 7y@A�1݇ �p  +nۃ� �n �;��@;v͸ 5ӡ�����r��)�;u� t g�-��eh�F��[Z�m�x  ]�v` ��S: 
�p h4m  Ӯ��ѻ�p :a� mu� ;�� t(�� ���حSj�6յ�MV�!x   ��( ��w8�@6�E�� :�6L  st�hA�� ݜ
 %�@���[em62�j�M���&��x   v��@t�j P�,��w@;����ꀺ� ( d� 5�:���uIv�,�Z��kb�b�  �� �����.  wu� K4 �8 �-�8(h���P:�  F�@
>�    �!*CS eJT�0 d0� Oh��)@ ɀ	�d�L�����J��@   O�S��4     �!3I�@���4Q��J�mIEM���42�4F�����X�5��u�^�\#���2��ek�8^��*�0��W�p�^��bW"�T��QU� *��*~� ��?�?�dETW�@����#����O��*��f���@*��>����+���o�������L��f2���&`s�L�e�L�f2���!���L�09�̦`s���l��G29�3+�0��̦a3)�L�fC09��fa3)�L�f2���&a3ÙL�fS2���a3)�LØ&0��̦a3)�L�fS0̹�3)��fS2���a�3)���2��̦e3�$�a&S2���e3��f10��̦e3	��fS09�d̦a3)�L�fS29�̆e�L�a3	�L�f2�̆a3fa3)�L�f2���&e3	�3�fS2���&`3!�L�f	�2��a3	��f2�̤ٔd̫�&�#�s�eE�`̪9�ʁ2�E�#�s*.d̢9�W0(�Ef3
eQ�"9�G2 �2��E�aQ�(e̢9�2��Uʃ�I�G2��T\�+�Ds�a�"9�S2��Ds �d� 9�0��L���s �a`P̪9�0"�\���s"a̨9�0�2�� \���s"�eQ�9�0&dD�Us.e̪9�0�\��C2��(a 3
�@�+�s"��D�s
,�&d���0(�W2(� 3 $�+�@s�\���&L�fS0��̆e3	�L�f2f2�̆a3	��fC2��̆d3)��f2��̆a3La3)�29�̎dsd�L�f2���&a3	�L�2f0���e�f09�a�`s)���29�0̦ds�L���0�L8a�:0V�;1�nU"iH�J���b���)� z�m�T��A����>S����w`6Gutٶ��WN=�V�wj7��fK��z�����9�س����c5%����W���M�bd ^>5��n�|7\�A�b͆�Rlo�A��_[��n�Ә����f�sQ�Q�� <k�QRXko�W����'�V�tn�T���%�X�[���ǔ���B�n���T{�+;(K�JIEPU��5��� jв�J]a$���k .�i�ڬj�V5�m֊�ʼ̽#Z h����Ɋ�c&ܚ��ܸܮ�B�0�*�K�uio���ȵ�h�ՈC�b��N���t�
�i�tDp��*#�ٙp����V���;���0�A�7yV�����@;Fn]2mn��$�2<�pdϊhH�Vफ6�mKXtb�;Qd!f �G����P#i�#v�
��줢X��mJ;42���k0<`<4����)��B7vj�z�=��j�֫u�j^��3�d�*�R�)�t�<���>���t�z�4�Kur戠{6�&a�x"�k��ҭg0A��=F s����:"����7@m��a����S~�f����
�Z��p�bכ�O#����**��)���S-R��N`r`��x���r�e�F*���gx��j���	3��r-j��-�mMSt7c*]���b�1������]5	���Qh�x6�'�bOwU ��wr�ZL�Af���D�Q�r�+!�
�n�S�7�;�4�7G���x����X���}o*a�|�u��eX�*;�� t�S2����r�KlM� ��t��3^aZ���.� ob�S�!�cS���CK�)&Kmh�ժ����[3˙zޡ��b�+���֝fb�A��ac�-��;�x�(7hD�7a"ûd���qΈ�5i#V����\�wQ!�Db9W�QQz�s[N��l��cv2�/�A��-���Y��ṬgB@���p7�(����ewi�@i�7��h�)�*�<]����MQTv�L-vƆ�I&���)�-A��W�s73t��T� (��:��٬��Ch�Ǥkd;gR�C,���+$�[Ya�PSI�I)�C����(Y
֜��*��^-�{ /#{W� 5[y���E����&���F�[ :6p�(�2fZLY��f:��K�1SWV�,[.�{b8�7���Xx2�T��+���Z(��%��+��L��h��s*36���,�U�f�����(.M�a�!&d3�l��R��q$�ˤ��p�� ʶ��Z�W5:���!��(]\��j�[ŗi��"�1g
kke34����)e6F#�-���u���N^$�mk���������i��ы�Z���*O�:|x�>�a�kN�&���"e��]w�z�@>��:�t�D���L���g6�*V�8��-K��r+{�@��hi��t4F+�Ju��`��P����H����ǵkr�:�f�:�@�g0����ae�Z2^6kJg΢�-��F��zN7K�DZ�Yr�	P,T�Ў�Zԉ4)l	=t5fޥ{�F��Dp�F#�'�����G�r8�h����eZ�pʵ��kV8�6�V���2��l�l�zu��ѸZ�� n����*m�.�72ҭ�2��k�̛Y�z�wXhĭ�a5���Ř(�&�?����u����(ml��1b���76\�	xr�,eP\BA�}Y|�n&2������2�U�mJk#;)�̥�
ǰB�mb���/&cۄOr�@�B�X�*Bbz��P4�i��b�d�����b=Ѣ�X!�%�V�q�Mi�Ne-y�{Z@H�y���2����T�YY�i�՗���>�����W�I���l��tU�߹*f�S�;A@�n� okks��x�e�ؕF���@"Z��2VA2��~�j�)'(R���D.h���wqTB%p/�"�^�(Y��5�k�x\��҉<��1�KʲP6v��w4Ƌe֮ͭ|�x�Fe3,Z3K?F�V'�����Z�R�ia*Q%����f�j
��u��[�FF�Y�g����F:�q�(7ڑ�Kg�x%	H�,9�M$w#��u�p�B���8��5:F��ͩt�c���)�V�9�w�=��'m֥\�absL�u�Mg�nYݻ�riԆ��I��J�+��^�&$���U�&��L�w{ �^�S\ƌյ�Mfj���gf#Q�Qd��y.Z͐٨����?Z`F�D*�ɶ���{N��f����!̃�M�]��0lĦiݺ�X�
iL�@��H��nk�V7)���l��;�*:f�k$U��&�PThŗV�Lմ����œNe�I��,M�U�o�*��u�3Lj�nR`��
"�EBѹj�ʹ�D�K� ���U�f-��3�(����0LB<����4���9����
.J�6��U��,�M��4+
�]��������e�DH��+
;�q�Sn�W{"q/)���Al���<B�A��E=��2�S(�R�i�c�#��C��	f+��ؚ����rVhtwG+i ��˩�y3�4hԷ���̭��n�]:ڸ���Fm�pʄ�Kg���M<�Ȓ&�:���F�U�M�k����u��RnZT�q���7����F��v���QYsY݈懻VRf��w�c���c�F��W���nV�q����� �����I2Xmk����V�[�!k(��k.�T@�TBV���*�m�)�A4��k/Iѥ@���m�:��R�=�cCס{V��n�@;�0;��rm���H���2�ռ�l�e�F�+i���$���`@�W �Ȣk3`����Ц���f�Cw��4X���V!-�\zt�Cij�̳ID�`"�7{[h�@��K��<k(ddˡN�֚��1Xp�)�@+(�x��ɫD��yWD-5��0�ō"l���V�j/���j����772Q�<,�B���%��T&�a�N�Uv��6��X�1D
A
�X�ɗn恔Cc1V�su�S�3)<�mcف�V��	��p$�˺���$�x*-��{�e�*���v2�� �Kt�)�[Ø�c[���rlL���4^&��B�f�m�a�����4t^Jt/eiP*�
n�R�[�)V=r��T]�bA�j�B���桧(Yt�i&� �8�8�C��G��ɷ�L�����Lf)c*�L��ETF��s����[�� 9��z�k'�urMݓa$(�P:��%��e出#�$  T�@�9ô`5��B��DC���ie�"X��m�J:��(�R��������@��+e�4�m�9y��`�3#�Spa�=5��ȅY�6A�[�׸t#5�kR㗪33c7D�m�1D=�Q����	��nb�hf�s[�3&�^M4�k�_9�^��4#vF���tMff��ouE���!À���� x#���E$�7���%!�P��	s6B�d7�¥P�F��i��-��T�T��a��r=��!C�҂���ȍ��/�I��k\�0��ڭʦ�kh+�I�z�Ya�N�#Ĥ���`���`���H���܉�(�\��X���CEY
cA��!U�ݕ�z���ƬwbX$��-� ��Ϧ�of��]J��weiYq�záQ3e%W#���8t�n�ا�Ҡ��b�Qct��]b$܂�{�3+pZq�c4��[�aX�^�����+h��Jri n8důw8�x�N������f����R���oD��H�ⵍ�I���KSɦ���ahq�s%�;M�j8�ܥ�e#�n�`�t)�R�E�¢��T��Re�!z^��DF3$�kt�ѐ= mf<K`Su����`�Y!��/P��ޑuӯ;��\V.�n��hlq�^��+QɊ�ਠE�����c*:��;�Y�I�uqhnb�NV������nE�3����t�J��[�PS/L P��SEmݡB��cb�F��j5GL̺�\�tr@�9�W�	xwY*��V+f��X(e��.L:i�1թ��F�ë0u�N�in[�rXvml%2�aHW�}-�v�Bf�b�;
F/ I���ᗠ�V7�%��+cL*�ZC1Mف�*wYC2��ز�L����j#�݃)[�lSt�KN�e���j%����u%\Z4��~�/�MU��e�W%bG�1<���e��|��c��N�I���eK���K�6uJ��9���Ѵ���{�ήh��9O8�O��vt�c��T�0�	��i���f�B3ܕ�0&�
��R�yGEJ���9�elE=v .�h��Rdջ�1��,U�R4F�v7"ի���P�T��orIN�L�hF�V2���V��5����ܑ��wT�~Pk�Y�yc][��t���⠃���h/kqU�֝u�Q �A4eQ��IV�ƛ��r�drI��Vj�C�$k[%^�u�e��	B^E���Hj�I� ˵TN*��P0O���Ϧ\in���c�qb97�Ԥ�����pT n���6�L1
x7dP�X�͙z"�.��+#�k\�-������aæ%{*�`��p�)V^�,̛�=ĉ���� X����k�"	+&\Tw��sm���U�v[hF��4��0[sMj�?���,�c��%ꎱb�/w-k˳=�P�1��u�7d/p�,�E��Ε�I;��s,���c�"ڮ��&���ϵ�@	^�� R��{cv�棩0C������G����5�yԯ�d����#�R��x�*�m1�H%`Y3sJ��n�ي�ۊ�$�X�D��M�	2h� T�r�kZɴ�U�pڭ�Y�^&ZMѽQ�Se�4C�E��t>U���5mL����Nl��2TJ�E� Eق��X�c����]m7����Yx�q��b��v��
��$�� ��cQ��-Y�j�{7V\z.dn��fV�{�y����{(��k.3�<�92����f�n
����}vN�RNKLJ��ui�:W��Cf=cφ�Y4f��ݐ�3!)����If����&��؍�R��;Z��!X@���'�~�Yy{��T��X��OT�U/��2���Y-�dS8��f�]Pa�M�)�3U�a����3JM�VSVM�����Z���R��ei��Z�=�F�m[;[��S6�	��K
ݨE�����h��x�QAp�.��M��G-:T�`A%a߳����ő^P*:4'&����#`j�`L���Ou˄��W�,��:M0\��ը�kz��v�CeT���I�[�#u���*�aV�T��
�;)�ҽ̈j[r�K#�Pn���-Q��t^=4��G�&5V�94��Y��6���3%lȕEkڛ1�,m,� ��s��.�v������M���+���KfD�n�ŎED��U����Fa��"�@YhT�6H�a�K9mIf��KA"�3�����Q�:���D ��q_�д�2�I�܆�2��F8���Nڒ�
�b;L�KY�Z�����ݻ�N��*�K�d�pCm,�ӗ�0����-��J��Ki�MS ��9;|�^����n	N��pS2����C��'+��(��7t5�-V�^˰������+
gN�[n�njSMW&��ܽ/VQ��ux�[1�&��
�wa��q�L�l,5*�r�R��;���(�*{5b�Dp�ku�R�y�1��+4
�7�GMn����呖�gFR����[�Tj`�u�WC�-JI�,`e���e�����ȁ�R� �b�HI�LX�"����3f�ujV�2U����kLw�V;�(�R�m �Mnl�n�Z�ӕ#T��m�#���&�V[����f�@bP��v�2fƞF�=�E��U���L��R���ME�m�.�P�F��w[d�2�n��q�J�� "��>`�z�u��Օm��_*�Ǔ��'}�j��gD�bUaP�HI����uf�fʫ���ZF�ڐSMdZ"�A�$�26�i�ol*(+��6t��5�*�q��ʬEh��[Ǖ��6�\���H�bu�bY	T�)n��h�Yܡ;�y@+[i��#�0O���.�K$�"=�lK��B<N�R2w_�_ Q�<Ļj���c|oHHͶ�,-�����Ո�z��O^�u�4E��:Ć+��d��&�9�Z��2И�n�¥��ʏ#1U���Zta�0�Ŷ�V�Z5ol��zQ����(JsZ�e^4\f­]��f#eT�+cin��i��� Ҕ��U�^7���V��S���м���`�J'#ǀ��4�V3F�
\QϹZ<+���7e�E��'!�_A42tV��8�Au�6qA}]��;3s��wȵz�]��N�*�X2*,�c[ף���%-;�g���I�t�}��Yt6���c4�J�b�.p��7o���[�q�3~�G�j�#r�AK��PAA�Ä�\H��`�*��s/��2���J�P"az%mC�IW�ߦ��;j`��p��cY��s�D��P�!tyY��-q����(*��gf]δj&�)�v܌����Q���;����u��.�%.̦��0�~���F+4���d~wTBTT%��ͳ=K��,�UKu$��,Q�Ƞق[�]�YĻ���7(̦�9��=�E�V;�hP����
	u�T�CEfp�,PX��J����Ä9��2���YiՇ�N
I�Gmh�
��;�)��3}��`ݰ�1C��KuV����\o]��8����Ƞݵ�P.�%��*v)���V��8h<������-ȨP��>m)K6����y��}]�V�/[��߿=��>)�����ҡz�4�{�fAφ���%!O�Xqr�J�k{;�S[N6���ʝ5;j�Hk�R���ޓ�[�&��8c�Jn����T���]ovns���C5�J�ʓT{Y��-
�%�)K��<]Kb�AR9���r�u�̬c���R5u'c�Ѹ�ܽ=�y�a���od��e�5�_9Yt�c�om3�\ ���ll/�R�́�W���ñ��{��E��ԇ�S%��ҭ��o*���J#n����1"]�.¸TV��s���i�ֻ:
m�V 'S|MZGs��k��7��3:��N�'�rt�eA8m����* q��Rƚ�v�֔�6�!����_+���s@�+]��.��<-`���- imֽ�g?��Fa�^D�
Nr��T�.܊ڦ̾j�!j���%9�7Z'<xh>&^EM��}�sq�}4k�����+�;%v��!��7c��jX56�ѻ:8V�sf=�:+*U��V#�Jz����}�<Md��nݥ]O(��+�P蛻����szwma&�ú�*ϻ��]�ip�/�4��[�o=~G��L�{ks09ᛪOHk ��ZQ�Tdbʖ��v��=r�UWË�>ș�lcł_I��.2�u<����gat��^�I9Fs�)WT"����q�3��K5��2�Z����̳�������F+�=���y�Q�q��ar���T��W3�s�%�!�{�oT�� �5��[�݋�x��9�4�.�M���j�tB�O�\�Ł�ɝi�3�#�%��jGf�Kt�%������C��4�_r���k��5�+��me:���K��&�;@�AzT�b��h��u�5w)�yԺ��9L�m��-�4Y��0i�J�K}�}]5��R�݌zurU��&�TJ��;��pK��#Zs��ė�v1��K.S�\�l[-b��^L�Z���h����'�������]���7
�Wv��-Lf֩�bչ��I���J�v���VޥK���w��C(n��u�]�GK��o6����\����]n�I!���kR�2���`�F���t��m\�����v\L �=��螻P�f�	���jW{DP�S{O�"ؔýɞt�HAG6zZp��t�5��e��iW#���
"�1�.�
ZV:κ��]���Wsk��o|٥;k����۝\��ƙ
�,]��\�k��sl�C�p��O����}�$��{�u'�ƽ���q�ƐMx�+�uUѦ�cFm�§"Wg!���Rj�I��]�ydL���r�S��
�j˶i�F�tUס,�J��M������U��I;y������ݬ�A͠;�h���M��Y.��_b��Q�[�`
/D;qaڽٷ�*��:gf�s�~.��~(v�
�%��Ϗ6�h�.fs˥tyD��6���|�گ���q����*wI�n�&�Лx�ҭ���5�\��Vs�{u%�C�87r��.V���cڹ>!l+@�2uud2Ίc(���-�2����TK���a�ʮ�dpa��2�̘��&)�=�*�c',�6���F�Z�{$�42Yw�%�ʾ�k�&�ʸD�W�B��nɡ�e�ed6m`�n%5�Ö{�Z�K�tj
����d�5-n�7O�QržǪ��wҵ��+��Y������I:��d��3����� ���=*g�w���nhc�9@ucB�+/zi� p��m����U�p��dym;���r���ٔu9��L�QPe[է:	�A�y�if�(`��Z�����4�u���]�-�u��E�uHe��@�e�"�p:f�b� zyD�E7�5_j�Zq%�rj��t�s����fo&�Ĵ�w.�ՒN�wj�<�.̣�puֱG0d�{wR�)&f�z��ؙ/�t���z��U%���{٘����*��0wVFX+ݘP�3��P���lg!�(�,�.�7Ҳ�%p�z�,{���,�ȫ��J�y��#��uv��8�ñ�.�=&
���e׽oZ�K&�nQ��>
ۼh�}ӊI��u��������:S�[[���X�:b6�� ��۶�ξ��D���*�mP�(4��J4����K���i�Y��^_M����$dGr��B��l��"�:5S��]l+ag7 h����`����T���
�/t W�N�9O����Hb.���Z���*s�t�t@́Vέ�1M9���7���^8o{������Xv��Xb)����5z{s���>��9���F��)qsө'
¯�3��yb�_s���*9%X��kM�#hgX�wm�?������/��-�(߅NEl���iG2���b!BE�L���Y�]� ���iYBK�����XX�GP�gj
�P|{���C�ɍEN`ˢG_*{�_S��^�Z�k�K�N����a*�d�SzČ�]��`���>{Q��)dǶͭf�FK��x���7���f�qN)[���U׏���h���/-^��`�,����K8��}
�:�� "*�û]H�*�RP`��֫���cc���GF�9��ʺ�ou�e^.��6�(v0�0^��6�u�d��X�3q*4�3Yп4����ӛ���Q�B��tRG���Զt ���c6�@�T`--���m+��w+�R���
���^e���	jBj�sZvQ�ݮ����R�k�ڭ*]O���&�Sz2�ˉ򭝆k��q��κx�Z�Jm�Cw)�']��R�0��@��P��^R�&��v$%HL!4 U�hWk����]9��Η.#y%�r��<,c qrqò�q�ی���DQ��:�]���%��=\Ʋ-1��g:鈮h�̩Ji�'�tz�ˑ��+�mg'�=�}�w��D�]C�ۡ0��K�dz��o�s�݄��5V-�3�g-Ӷ4ed��r7�s�gk��0-l"]�w]�������},+��K�����A�|�m󓛓��ݮ���4��{>�jR8��h�%\���	}%��vs�P��nҔ(q���!���K7�����,��q��7��5�K��&�7՘����S!�`VNUkwnd�~De�%�+h$�c�*iX�,Q��v;�(�:,P�ND������P��P��K�yu�C�-0��4�J���ݹ�-�
+����c`���|4�K/��
m�q�®�vy��)1� ���Bz��k41&wJ�X�N��}�/^��-�d�D�s� �;�ݔ�Ӕ/oc��fa��Zv��T�l���c-��:�1�W��(P�œ1R�M}�J3=�L�]�����,sh�u`��"�(�;�Kl�RvCڮ�rY#��B.�gu��C!SY��v���K27Z�4.�͢-nJ�v����Rw"]�s�A䉑�~�4#yz�����y��V��
=Ɗ�m��8���˻��rY���[��q����8�k�ٽ���pS% 5�m�r<v�`��X�Ezq��e���[5h�u1�VJ��fӜn=�:�J��ݏ �n̛V�^h�k���3B�Y�9<17|�q��u��93E���w%�%]Viv����urX*L�w%9�̳}5;w6�jEw6�1L^�S�Y���gaAۧ�èL�L7��Ba��<��Yř�2���kMIZjK%��s�6Cu�3���BŌ�۴;*g1�S�H�}���Lv&G�ي��ݖXDҰ)qҵ��3s��o�
�����?Gſ����^Q°j�3�a��kd��A&뀘+��>T皖|���wRB��;$m>�j�Z�/F].Q�1�U1�]�L����3v_N�p�[y@N��J�)Qۦo�h�J5��w-%ߜFr�GYLӋ�/�X�y1�B�qO_��j
���Hd���ɬ��r�����h�儉k@;C�!�/��g��g#��pzޒ�o�/��ה)SX�=j�Xř�F��
���4�������[d�]��1閜�cY�kM������!��Ϙ�kX��L���wя��W�;^.*��q�Ge��ԧ��4&��lǅ�nTa;'�U���UV]<[%3:�^��9�i MYv\�	��+�]��S�XC�c�E)V�ٖ+��.����S��%$�����X5�ʱλw]�����6�^p]��*:�K#m��G����Yv:oG/{&�Ȝˮ��1Vr*��DMfA��Ք/Z(n�nea�[N�+�����W��ۚ��I���䚡��Y+���PF�a���_�ھ��WS�S�r�oYӪUc:s�Z��Z���n����'��.$�K��6������$X���1�rRμ��ۑ�c���JE�*�ZJm�
bFQ��]b���qK+3o�e���^������j�hR�Q٣�V��-di�ͻ�#�Μ�w0.��1��s����N[���
�諷�P�Mn�C���%V�n�+�}�zҡǺ�2�c�o_v`���"^��$DլC�|����:�]���bF���=�T�a�n�!	�+��A�`����]#��}Hl��.���5ڲ2�hY~����ƺBsSڤ�Ve�i`�Ⅻ�]�ɔ���R�4�JH�a8�����AV1Za�F&c�_f�U��T�w�(�!��N��K\��@�&��%�f��R�,luo��s=��u��.�H�тT]x��tkc�p)�;�jOq��wO���1u�fT0n ,��b�^�ړj[�A�[�l	��e�]^\���K]}Պ�AW�b�3��(��>�}]��	��_L.����h�^�8U�Z-ۨ�;o��s.kKDH��-�g]f�1Ȉߡ����tK�YlecI��l�ɖ:�:�#��ɒ����ƅ�\���.z�>n�����f�W ���P�+;�>�����-$��y�;�V@��b�C,M��ZV�Qr<v���fN�A��ŢwZ<i0�$�[�O�s�0�+[�7Ғ�h��K�����0�م��
b@
�Z�t�������8.Ź4
�xE���ݜ�K[�fLy�.��J[N>J���Cn�%*��h��n�cV��ዜ�xUt.q�3�
{Ntk�2_�%��G��-�iҚ4��
V��ʮ��Zf��sc�uX��:��G�QV��앗��*�Y&��Y52�If��\ܧw��ʺS̹PW���A��ж�^�)��1J�uB��P�>�SVwli�P�-�zi�Fc�h��PlGrR�:�c��*�[W�fc��a7���k��:�G�U���w�#V���3��ד��ԳTКG�w#�iX�a7��pt�=��	9H�u�)R��#��G�ʹѫ5ݑ�k�����g�4K*�id�޷l��fnޚW8f3h�}ދ�l5�N�XIP�����*ևcĂ�;���x�9�ce�U����D�����{6�Auҏ�����)d�ӑ ���M΂�c\���ok�y��0���X{��%\o�
�V��u��ș���ޠ�#���u8�af�F2�V�+TK�B�r��ۻDǔ�"'`��ʓ{W�ڻM�p��k�U��d�9{m�h����m�Ӭ(�hV��T�꺎+��w@	�f�a�Lٌ({B����\u��*N��X�k�w�����ogF���CH��$�կ�������F��hͳ���·�Ȅ�Ԗ��%l;F���Nbi2���C�RE�vg׋v^��V�_��l:Rb��Ї���Q���V�<(�i�qLq�0u���ݾ���=앝#8�B'']�]���V<60 ��X���/������ܴ��u݊=9`]vv�2��5���9k^2ќf���|n8�Y��-Z,]	�"ch��K*�K�^fd<K����k�M+W�an��Ր�kU� �j�Z�T��m�N�E�v�܎�Q�%M�-��c���0WD�]�/D�m�;2�ᱚ��*�{�V'
���9�����)f�{{�����;i�V�.|��½�n��`{�p�l���S�l,�>����bS��6�Y�H-�c9��g��`z��fVd든�S�^[�/\ȷ�:��d�\��<@���Ĳ]+u8Zvk��Ym"���#WX���R:�5���fWe�Z�_\�������c�+B�0Ie.Qe	Çٷ��[���HΣV�2:�bݦh�������y1;x�&1�(���e�Y�֗�5PK�C�7Wv�e��tG��Jˌ���ƥ�k����aH���V���.�
*^ֺ��<w}���?-��C�5y�)d�T�S/�L���I�n�=%c"�:�o�����D���m�VŖo��xrhHC��n�(4��1��*fܚ�]��\h�I��J �8�&d�m�u;/z�%��%N̎��F��Hy�\Z]�u���8r�H�k��ʛ�l�M��uѹ�*�4�!NHӒI$o�U�pl�'㴮�TX�}F^��6��P�\�O��ܹ*�{b�Rʅ�;m����P#��pR胤/,����[P�����n�U��L6�d�Ѕ�1�q5MR5��~��:>��QUW��+	���-	t��$A��_\�Ey��3!KO
��q�)������M���4��M��C � $P
RH�P��"��� ��*tn�t��X�`8$�GѼ�I�[K���� ��[�SU��
;7�)��\i��a
�@�٘ka��)h��Q�m����Z&��B�5b�UI@`��⺚�L�
V�.�*���{C`9t���w�Zִ[8���� Q]�O�Z�
�[4�/�f��a�""�����5�a;mm�ӳ�D��yn[����B�����N0f��Ɲu�h���hƫ^��-m���h�Ĳ��pȬ��evW �MvM���	S{' ���RNVCIQ]uc�[�F�9������*�WW*ݖ{x���Ы��w\i9G_V$��\�`��V�U�Y<��oK����{��M<�M�iTgTS���Ԗ��0հt�/���ֆ�֝���Ӝ ��,%��@u���|�i�SE�<��d��1��E�}&�u��]��^��f���)���Z�T���w6�.�\t-���X{�����)Fe�DI�L�p��M�|��s�Y�#�b!���{�Y(^Ԭ�6�س4)��j�n�ﱧn��7.���-QkV�¹���5Ybe�п��-96���/��Kjќ;�]F�V�= t��f�ϰ�oegWgb鼷c�JSE��FP":ۆqۧg�����9s�s�Vۢ�K��d�t�hYV�]׶-DV����ɦ�[�|�e-�f��(��Z�4>ͮ�yv4E��&�׵jW)�":��D2�m2�/�V�#�C��M�[K��8Yf��+96
���<�s��5�h����x�]ƒ���FlpY�]˕�̰",Դ�:Uw���t���f�a�|��2�V0��t�L��wI8gq(�Q<��d���͠�Q������e>s/k5����|��/����}>�G�o<x����<x��Ǐ><<x��Ǐ<x<x���<x����x��Ǐ>�<x���Ǐ<}�x���Ǐ<x�}��o�����Ǐ>�<x�<x������Ǐ<x����Ǐ<x����<|x��<x����Ǐ�<x����Ǐ=<x��Ǐ���Ǐ<y�}�w�����Ls �n��Vs�B��;���蘱,=f��<�8x^wx�!ZLO:Z�o#B�Pp�{;��ǲ⡍A����w:���"����c�e����V�;�۹Ê�����2�'3`�r�-	pn���1C]�W87y��b���j�^I;�����h�����rԊ�m]ݺ*�vC�
T��9�k3t���srW[���v��-�e;
ZO�ko]�W[��Ru��l���b3�Z��^��j�hl�y��J�HB�*�1���e����D��Uî[�tx��������f�}�2��B^e����^��={��2�p�
��D�����}�JO%��:�#�U{5��b��r���Qh���5�ڨ�U���q�����F�#ȧbZ�,c��vrf�9����9���n��n}��F�t��Ʒ��>�J�؂ed�jv�Zz����[:�6H!^Z�j��S`��Ucd;�Uk�%�C�-�955I ��7;
�OT��<�77�\�hT�g�v�m1܎�K���k���K�a�֦�q�*��6��,,^H���7����>�A��0d?�lbTos���v޳�.�pR�A�VD��m�*������2�tջe;lf�f�^���):��@�=B�e����5�V��6�����jSj�z�}���������x��Ǐ<~<x�<x����ǏO<x����Ǐ�<x���Ǐ<}�x��<x����ǌ��Ǐ<x���<x��Ǐ���}��o��<|x�<x����Ǐ�<x����Ǐ=�x���Ǐ<x�x�<x��Ǐ<g�<x��Ǐ��Ǐ<x�x���Ǐ<x�x��Ƿ�[���]yu����e���-p�5�}MI�@ɩ�a�r�An�<S�Ö[V��9��lu��54��[�c$�m+�,j�5#D�*l�ޒ�L�5\����
�����sX�.�[;8��s��gbܩ���U6���ӲC�tc|*�=j*u9Ҩo;dwp쌭��΁��t�˕]��3����o�eV��)�]3B���:m�׶�.ݛ��]Vg&�-���p�-v&0�}X�n��ބVad�����E�AB�d��[��<�3hH�զ�n��k��U��;Qu�Wˍ�	u��,L��s$E���B&�C9x*b���l:֦ݙ�7��iF�T�օ�Z�͹N�$WH��W#�y_S����Rw�I\����|;������_t���6��F�h��i���2��Fl���e E`�_jg�%���]5���R�;����ld����Ћ�r�]nm�:+�Wv��2��'���$w,�p�ɒ0�\��5��ũ��2���O���ܿ���n��SersF�Xc��§	�����r��c�h��v(�ߍV� 7a��t1�Ln�5��H����J�
hm���P����ӫE�x�%�\q����:gt���^�E�I����z��+��ѕ�7�z��pu����X��E�)-^u-�6m��3i�_8��<z�v�y�������2���WKq�8q��$��e��@v�!r�ы`�o�j3F��Uѵ��*)�-��ݦ�v�=0Q�/�?Nۭ�9\gĝ=��En��f��#.Xt�Mc
�n���γs2p�F�K�Vf��>�)S	u:s:���GQ=�^�32��5|գ�:�Skz�+��Z4��O�Wc0e7{L�7Z);��S�W�h�9Y�]C��ಱ��']�[Y���\�+�N��[�FR�������v�7��Z�37N�<��Vv����T:DQ^_U�Moc�.��]��Eb��@L�4�`�^���D�x�hl]R��j��G�w�d��X]z�@ ��Y�)�r��Y��e��^R�����������Wc��6N�GU)��0.�9�f��t�V��.�E�F>�y~��䠪�J�Z8�xhB��X�M��t�.�G�.�62-�Br�Θ� Ҫ�X�x�=����B�c%��mbT%��5�_
�ݡR� �Sz��MNN�`�ܱB��2Z�|��F�lO~�N3�m�N����=�/{RڧK��ͦ���;�C��<�����nk#m��z������5��ڂt�J���J�n2���S&�}{��J]Xs/�d��o9WP��5�U ��Jg*��d�\))_c��b�Jѽ�ˉ�9�8 ��x����ٚ�\	ܹ8t���x]w܌7ǵZ���aQ�#�W�j�eB8W��&7^mFjv�z�u�ZҨ@õ�\�r�㭆�(�(K�j�^���$�K8jI�A��.��]��vM�}ܕ���+��-���3W��J���`��y���@ovA�Pb�T���b��Cm`{f6ԭI�5�页��`��S� �Tu(I��:{��w�*�eH�dx��"j�K�����eu��O:�`C-����1��pV�BL��u��[�X�B�A�&�yl�_#ǅE�ɚf�c#���n�ץ3ɚEu�g�'Ăjv*1��q�����u��%�_H�w;s�s�գRL�k�Ȟb��7�����*c�ۤ��,��GX�R��EEB��f��P�Sb=��D0��MP+lj�+���eۙ�h}�T�'��]��D��gM�-[���.�ܩWJ[u�(��0I48`��Y#�e��C],<7Ld��m^�eA�.S�Ѿ��`nX�i�� �������Z�f�p��BM�ۚh���^8�஭�ہ�C��90�Z�EYQ�F�`�����ޚ3�9f7Gv�Vw��"�j�#��-pƸ�a��0:Ʀ��à�ղ�-��l-"#+L AI���$���/n���kZ�B�Ki+�Ɂ�w�P��iC0oJ�-�T
:6z��'f>��.���TQC�{�Q��WV�k2d���L��[�π��Z�B^����5P�M�0��0QZ ��;��J�&�j��s���ӥ*WR�DunԩAp]�um1yצF���ed�(�5�C�kq	O^��G�-[��;��GAI۬j�+3�����
�ƪƦ(�(�oM��k�)׃^�J���n�ynҙ�rI�n�v�+��\��%U�"4�[0�X�d�tpֵC�~>vgf�l�2a-
�]b��]���f�C>J��XMr���,�ŷ]y��K�l<���M�/r�r��8�,�J��$V�賩���+j�L5�5a̻!�&�8h�E�DX������_-��rj�fr�f�.�^栧-������Q�W�gj^nj�ۑۭ
�I��5,�(�\k�%MQ���a;tb�[O��v �ٖ���]'�;W	M��9�����b��.{'a���ϡ�Յ$f;lKB�H=����0��F����g���\�y$��Uv▵b�������᠂}��DfC�eh�B�r�p�����>����rV�8�J�ے�ur���
*$���d��\�[k��鬍��U��yiD��}�Y{ڳk;�id- ��x��Uƙz�;.qO���h-�.�ͭ�p<�Ri�"}%f�j`O�+U�}���);���.���sF:DŠ��f�yi��$ݥ|�fX]��;f�/������/�Q��ִf-�.۫�T��]���giZM���u��ǻ��9��M ��]$��{C^$�)�:;q-emѻ��2�pz&�Ǳ���PM⦯Gi����ۆ0Z;W�(UL7Zs���(�b�����X��Y��%��f���B]E����A48�x֧��!��T��v�^l�o8#W�:�l�= �7o1��;��D�d�R���L��P��0PႲu󨑛ԗ ���ں���B�{r��r�Շ��V�$r�6��j��2L�J!���X��XW\^����:l��g[awi�]IX2�5��M���3����n�
���ҙ[M3Еx��Y��+���rDee� �Yu�u1����י2@ݷ�ߘ�m,�V9�LՇ2u�Ԑȋ�/u��������p�+���*��M^#6�Úӑ�Ys��U����E�`[g"9��[�޷з��M�{���YJ�t�4�|��]a���ޱT�W5����ˍ����,'���.!���Am��r����545�� �����nǪ�$�Ηq�wY�+�ҦԩP�N��$�5��&��v�!��V;k=�'j��H�W�J���N�:]�8M�F0�a�d|���U���sjY��3Ѽ�+����G�I�.ї�3���N�gIGۥ�E�I#ح�c�,��r���DZ;�]!-*ۊ�Һ=��q=����^3Q���vN�=n��U�Qё�Y�@m@�hQ��vcK\�������o]A�z�J�����Woa�+��m����7����q���O�:!P��w��-�e��q�*�+)+�i
٘U�ׇ0AZ�]��K�y�������46n��mNy�D�n�eJe��Va��<����/:�6�ԇK6jj�9[ _˘Fҗ�[�P�ձ�r�_;�b��f�񀵮�����Z-C5-AP���nl����wf>O���bTw7e.⥕�l��־���*�&9��'�쫛W��	�ː�+I.�*�d�v2�kݙe�o���΀��H�R��,��Y��іa����(���hWmeI�:���I50�3_+��ź��T<�{�����Y�d
b܍�n�[��R�&��fU�Se�B�a�)���^j�f%9e>�7l��q"�����Hl3�j��D�6���:�҆p�'HG����
�Tx5��[�wz���\UӤ�H��v�����P!;�yK`'~�T�t��x��&�V��$��s�(q\�=�o��|�v\�\�
���׶�����7LP�6e>��+-MzK4�M+��cq��}�����9B�}҅j��}�-%
��ʴ[�_V)�LYÆ�<B�[\6-�a��ve�Qn>yU�����k�����g+��G�� r���Af�����Ue��t�̢��i.����ѩFf��Ma��Y��Cv�����և*�@�S�o�:9��� a����h;�n��o�e�h��;/
��s%�WV�b�ܬ���, �s���Zg2$�Ҵ��F�X��Yec�a���eƸ�iT�Eu���,�K6ݺ�F��X�\B�[i�{�We&,ְhd�͋.���Y�z�8��|ª|8��)��ӆ3��Ŏoe02*͛�_*��(���6A��V�H8�[�V:Z6����5�՝d=ϻ�&��k�����To�#�]:QR�ح���-�x�U}�'�&ڡխ����Őb�x��8�ow������H`�L$�NU���?M[W/\��]��\�i�Wb)���}��J�c�m�7�T=��p?i4�A�N���JХ+��4�6����ӊ-]�W�}{�::����b+�K��+0��6�gҾ�0�^�]����Z+Nzۘ-���g�_s�NOh
֕��� ���
�N��w@.W�"[�� ��%��0��}���T��E5Ք]��X�'��x����v�)�c0�&��ӕ-��
�뎻·���ȳ���gu�S%��\�"��}�����c����^�[��@�Jۂ�4�d*ázۮ�9�|���z�]Ytl�,��	��)��{a}�?�`Γ1�&�Ua��:"w�Q���&�^��[0�L}�8s#�wj�y�6�m�p�C�F���"Y��&r���"��;�#�;
����/rh
V����w0,��B�����9=-,��1��jC%��B[֐Ҥ��ӯ̘�\�_RU�Z-,5/���ü�x#g5=J�雋�w�Z�u�8����Ҫ�SA�	�g{��u:/�p9&v;cu�g�����-=��3�U��K�w� ���s��\�'V�ҭ��9��-`����)���d��n�UN�LeЅ]���Tl$�f9��nK�}�ǝ*
�����(X:��V��\�/)��3_[�
f�a�ŭ�;�a	�]i71EN�D����-�r%��-W��0�g�Y��[B���\���$�����1,`��FC[�����ƣ]�-e�q��(ݙ.��h�0\����1\r�$���L��7�*��؃��_^�=���-w
Ki����I��"hM+H�+h�a;�A�e�B�e+&?�����nM�{�I�V�&m`Ed1�R��2������V;p�t��MD����6��z"�[)�N�4�yOY1u��
�rfWb��f�Z���R�f��,@�ʵX�o0PJY'u���%5# v��u'�*����n��k^,��Oaf��x@Z�xR���@F�Y��[�M҂!��Χ&n@TY�9��e���쾫ʲ��Ip�}܃%'u+0'�:�/"�%�N�7�p�IoYCX.󓨫�¯m,��W�B�Z��:b��i�.ϕJޅ�6�O�J���T�ݚK��Q���i+Z����\t2��[�u
��]Ft��mY{���a���k4��Zgb�1�E��{
�W�6�'
���[��&�s�� k=��,2`O����;+��ѯiV�EѭQ1�|;fwX�
&jǴ�L�g�V`LcS�;�UYטD�s���Boa��Ieܩ\��$nMvno8��X�����>$�?h��1���(ĩz6�3w��Nu��m���g���X�������8N����-�A���V�����+�<�T[��kr�wL�������2):K�n(��C:�!yU��Pn�@� ��<�5%j�ͤk:D�{-�[�ń�*ВսVo�6��V��ɫ.2֚�e�ѿ�(�B/�@$ٺ
��]B��w�T�T� ��@!R�Hj*A@�'O�]���*i��%T�SADDDTW��z��h�����(&��"j��5S>�=����������~>�<g�&�
*�j���䙉��<�4�4D%4�P�::���
b"("h�"
g����?������~><g��1AEQPU%QQU_-LEUO��T�M0TA]lU$U�KLAC��TQ3QTHD5DEK5E��ATPQ54P��Q��QTP�-��f���b
%���" �mIEST�D�ST��E$ET�%��MS��*�%�"{�EVޮ�"J)"��"����$�%5Qz�m����5��D3Q%4�PDEA0EK�U	K,�%�owA�i��QQؘ�q���h���1�c�雫u��#�%X������Q�5�+j	�Fq��֡���ڧ�K��׭�t��u�L،�kNڴQQ	����ZΊ�l�:����v�����V0�Qm�kgm�*���U���i��ml΄�����֥-�;[MmHb������_S�w_{�;�m�)#{PB�fWtǳ��r�+Q�%�b��O��m�!�v�p
=�7H�կe&:��p����*�:���C��CY|(��w���Ts�\�_#��lUC2dz�i,)�3��s��������� �a=Dɡl��-� ���	�^j�[�vi�S��#��V��(�c��Z�Ɓ$�sƞ��6�z�7����6e���vبb�~�՝x�>�u)s�Jg��c��\#P�l�����=��;����ʄf,���Q���=�%<.���r�]�ԺL���󏤃ӼF��g[g�z|���S�([h;uY�f��{Ԧ�g�mn�+=���F�f��ρ�;D�N� �>�d�ʂ@3Wr毄�[N|��V'm��=)�����OL�ssO�-�̺��[Ue����:�c:� P�,%�m��鸡�vԎ}��{d9�sv��L���ޝع�:!4gz�ƽy)�k�F�ښ���·�G^���=�5�fHe��K���� ��������:`t.8��#��ku�N�rn.�����${؝�/o�5V�2��&�w������ٓqւ0EQ%Α)����oX�e������MZ�ә��!�$��n��U�ѯ����x��� 	�;A�����9}PE]�m����[}'��}/q��=��xn�qpޙ:.�	oa�9��s]b*�14�/l��U����4I�.\ݼn�07�R���������IP+�u��m�7�v��#����"��^���	�w���V�� �cy�s¥�x�� �k6��Wme��l�"�Uj���S���6�aM�W��֐3l�μ=�}��1ǋ��;��EG����i�>���6M{&3x�.AqDɣ�q&g-�\����>�\�jV
?!�z⦙�N[^�*�+�����߻#�=^��n��*����{wW���\��ޟC�j���m���ɂ`
�D���Fe�#�z�ܶ ܿf��{��x=C�x�>^�]9�gP��k�F��/���z��w�>Τi����e�yzh����lv�;�;��5�E�Z���1�Fƃ���5p������e��6g�v�$�SX�|�u����|����Y��������s;۰n/��~���DѲ<�ˉ�S�.��3��9m3Kvϊ���X�\F���oUұ��6֮��ȕ����8"m��]��t}N3G[�}�Jfɡ|[}7�}�W4t���Km�w3��h�Y[U��e� �݈/�H�-
�F����f�ޛ�+��I�rs,�KA�m��)��t~@o-�ܺFXt�U���~���kn������ߋm�A�c�u�T�w=L��(�,���)�S�T+>���y���g\U��sj�/��������S�\�����}~K���z�kȍcڷ���NįL�y�����h��[l_�K�V}\�\秭眽�� ¥�tߡ�L^�N�xyK�L)��޺�ހ��%As�͕�\�Ϣ�����Az[�qk �>�B�:�R^8������oҷ�>����e5k�`�h�P�B@�!m-�]S2WQ>��u�K*����ާkq�-�^S������5 ��Ɛ//��l���\xX%��l�?w:��8��O76�<b��}���s�4��|O���rF��im�8*��2�cM2)ޜU*�r�*�g�[���Fm6�'��Eq]t����KCL[�����K:�s�X����Q.dN�1���%v���y��hfBf��mN��f��})Z�{�t��q;M���2�m��`0�B:�#j�_��f��7����S�����i�^Z`�=D�n��U��k�[3o2��.�N��;u�.����p�;�Hxg������!v>#�Eq<�4�{����g?e#�B*��U�U�u�S�����{	�uL���F]�fn+��k1:_sM4E��^���\�Gn_�N9��;s�9]�Z�iZ��P�VO����r���1v7 mm�¸�D�^���Ѝ���_U�9=qb�<���T�G�B�W��O��@.�m~����9ޘ�&'7��N��u���6��K��������ex���
_]JO*�<�麆���!�=��
�>na�@?u��ϧ(q���U�]���[>0�&Z���;RC�z��υE��}�E�ޓ����Ԙ��Q�!��xU�z���	N��ٙ��ol9�['��X!5�@��y�!T�,ȁ����M�L�TC����ٛ'!���T>�hc:�Ͼ����V� U�Q!���n�"_��%�(V�$�Ҧ���/����z�^km�Su
Y)��C�L9��]ڭ3%KVC�M곡P�>*�
f�K\���t*	�VWդ�)W�|�/^�?_�]˹��3 U.���k�n��v�EX�����2Y���E��3��������3=�k�]��v�?)V晉�W�T㾝G�����������5�x���b�3�ޔ��d���!b�?g��}:�����m�*�%ru�MNC��Vtn�?L�75R@�����\��;�A����h͖ ��OV1�í��+�}��?΋����;�	��@L�����I�G����cK��&st�����I3�O�ӑ6�c*��	[�=ZwX�tx0׽�>-[J��䞞����'sG>ɂ-�?��o�ح��oFla�ڹ����Ј}��L����+u7]y��w���k��ُ�.��n�A:ƹ��^p�{���YY���� ���<O��mw��2/��G}^��Svd6���[��R�į���9d70YUdcXGD����ցW��>�S[��BM��^^u
��Ϣ����6R�s���P�-�	��B��}+��o:tGk[b��Ʊ ,b�r�>�l��E<� /��y��r��r�a"'t��'CL�_����^�ck�q�>�޶��b���]<���՘���2/Q����O�A.}���&ϭ����:o��o�G�0�$����3��A5���7�p��3p�����r�
~|�e_���dt������h��~�U�'��>�����#����$�ʋ�8I�c�s�d�k
,iy-�O{�e)��${^�W)][u,|��.�������Q^����C��9݌�5�7�舘�L���Z�v����w��U��*)�۬	rT�s�KA⠖fl`���Wclz��j�;éM��'ݵ���N�>�_.�TjQ6woqJr,�*9{��x�N��}�t��߃�k��]�3޻�xG� yIe2�h��.�D�����/ѹsp�2�=\��w���uܞ!���-Z�ٽl�2�g>�
��7W��O����iRr���^�n�x�5��I-�=�iWeȯ��u*fCl���|����e{c�yqP����LAh�?�7l�&	L����u.�����:q��<r%H3�u8v+)�0�ΖbH;�ԡ�N���@���[)]g`������"�â�.ܔ�j�w�S�O����9��/S~��%R��EM3�࿯��{XpIX��og�g�+��ޮ\hoa�OK����q2j�>�챿M3�j��}E���ތ
}��|�����g�xh �䁯M��������|�G�	����[~��Þ�iz���ETϋ��'��왙~����y��~0�6�31o�q����������4d
͓WŢ��ϏQ�`1�%��[��ej��[�ߘ�3�|9
��+��TG���������w��I�u��l��Q�}�"񻝄��n���ec״%�>qs�o�)u���r��=^r����ߊ��K>?\�%9�)z*����.Z]~��v����w��_J�*��pq�5Ŵ��A����*����_��(��>>��xD�{Օ;
�o?z	�T嵲cڨ�ڳL^Fd��^���}i���pe���6~��T�0��O���pŭ AW7*V��R�+tZ���V��\�=ONc��
9.J�!b���h�M/�|.n���7�s;7��O�.DdUv�7�fK� ����#9N�K�b�Y���幂u�v�S�_fD�x�K��Q������K9��se9rD'�Q�N�]XWK�4L4��Nm�C`�<�`���z�G��nJ�x��X��e�W���I+���P��MҎ�L@���z��2��V���K�ޫ�7���'a��T{���6�'��wv�L�U���K�W�$�q���&i�Dono�Sٻ$���c����)�U�؏	�ʾ�{����+�a��ox��]�rT8�Ԓ[�ޱ+ȿo�j��?�ܾ�13�K�*C���m�����,㝘^	�`����y���4jd�w�����Mn^V����խ� �鐿P��ϼ!��"�Zl��9�sƾ�{:a��u{���!��%����j��2�J��+��JyT^{K���x}���� {3�wr�n�U��v����oS�q�}�݁vczx����KM��vcb�Z�e�S���c�tchR�	⬔����1��3!�`r��J������T�3���1��e#_7��D�QV��ğ%0"��^�'�v�y66Uv�E�;.s����E�au��6V�6����W>֌���RZ���6�m��.jR��t��T��,��W��HӍ �>�_�<u�q!����n�z�s�K�b�D?q?9���5ⲼJ{t~_JLT7�<�x�J{�0lD�L�]gIn���>���&0����[	Y�& a0���O|_ޣ���(RLW����ig��x��x�X�L��=6fY�:��bl���2��g��[P	2/"��Gtq��a��c"s��<g��7}��z*>ߙ���b��3�x}U���.�:��4��0J�O2.^f�u�v{�����A�TLO[�k����tњ�D�r*�>��ϫ��=�cG���N�8v��ߤ��^�k��������z�.Go��
��ν�зeӴy��V�G�'��/vߨ�X���{�:r�W��ȣ�hAۢ���XZ���m��Z�9p���FX�)�El��ZVFpN�e�;E[������ �˛;RwcH>���;S��w;����SY˱����u䠠x�̮�d�W�Ra�bV_�ƟIu J�gsK��]��'f:��u�d�t "T���+��Rk�2���2��ŕ��}<(dޡ;ݚz��X��6�{=�!��쁉��9��]�3��g)�$\��`V��5lȉ�r�r�\N��ޛ �o��25�!��0�R���M���=LV�ëR�F�ٷ�SZ���OD�����HKl�:�>�."�F�4�:���3�y+��g�3GZ���J�{J�~gޑ{��{,5h�.�z�3��sX�U��딧f?"���~�z�~�74����~��+�)2�`�&g�^;����d �\����y�x�`w�#.DgP������9JˑײϹv��{����Ě�[L`o�h�q�z݃a�g��̓�>���G�U����'ֽ���+)�W�~��~yQ��\ϩөy�L�b�+�;SN�m���Y���(+�k��� wDv
�A�7}.�N�����>��ߕ��~���K�ƕ�Y��i�k�j��Nwe=��I\{DJ�5���1�c���"�n��D�֝D�m�H�澂�߲(ND��)��]A�v%�Myduuv�uJQ�p�CG]��:H�Y=�U�K�T�FTSW�b��x�ǷKr�>�^:c	I�E�B�z�9�J��[g'm�,����e7q:�Q��M�b�����n3.k�1cZ�,��p��3��
S�n�0>��v��R�2��2<�i��K}v����P*�j�]���D�8�uG�r�X1��T�� ��\j���Kh�N�6wZ��N��V,��I��-&��jd��q�<]�+�i����X�9B+&SR�c+lu�@�0I�ygT�����*�y���izu:z���ya#4���o%��T2Ǳ�{����`�R�����r�Z���y�4�U��9^퍫f��Y��з�GQ H�e�K	M)�9�ԃ�!N5BL�З*�j]F�N\��[zmO*�$��.[�l����&���Z�o�pEЮ���.�w��2'�7g�6tu]�]eb�w_fL�
�h[xu�
������lx����#�WE$�[�	M_o3�׉*�E�/s��ѦlՕ�T������R��`��p`��ɂY:���dڰ��m�$p�*r�����虲�T=]�����W0�!���N���ZԶ�E�ӂ�G#ԩhhVөJs�:%+k�\���[�k��NbP;p_Z��f��-��������K��q���0���!�*�G�"�R�lj��O.��d�aue]� �+᪃1V�Z��.�����&�h��Y�Z��9F�7��7���n!,�WAA2��v���mv�'v5�֎�Ps�c��D��.���6��#���e�`��͖�*մ�û��k-ͼ�lv�I����*#4
��h��5�[y͜m���o#yJ>Ɨ]�.Ү�x/�Łe��Ʈ��Z0����n�q�7L�\�1fܜ��N�Jy�Uʅ���oY�|P��A�[I�R�V	�K+���To&�GQZ���:F���z_I��D�w��v#pw�!pq,�!�qJ��h�x.�I�eâ�46�co1�֫�� /N�t�"1�#f�ԙ�o8�I��+ IK7�R�v��$r�wΗ�|����k�tP��*�êl+]�P���r�-�;R��F��[]Z�<+o6�1N�w��vi�6�ʳ��p�iҳږ1�>1�����.t����w��α��{�3�;��x9:�Q��"�/��`�,]ձ:�<��`+�ާ4i�=����C]`�;+���Gq���}ADn�6P[Ix�tO�^�AX�h��aa��7���8����"�<}ϡq��=YKM��ʬ�����h���-����%[h�aƵQ���yֺ�*Kd֫1�Ӟ��'մZ֭�Tm��Z���D��SA>=��������~?���������A�lQURV�kcZ�i�c:v�lD
/6�b9�WY-�V�ƃ�u�m���l��}>�������~?�����>�(���C�#m4yў��H�
()�m�c�h���:�J�b"h����������∪�*{���
�������%&*��(��h�h��N'l1PRD�Rk�������"��$�6�h�PQ!���4�D�4i1RUwj!�� O���
%N�Z(���uD�AE��Au�MPD�JQI��Mz�%T PR��0R�ݪ��j�h
�����.������h�&�*�����f�((������+�*�� *������KW�W��TxX�eњ��B��NO��$�Hι:瑄6��	`m�����6�F^���j���άֿ3W����OX�R`�c�V?��_U�P~͜ol�Ґ{)��	H�4� (��M�c��#:uʇZ_e�N�By�=�����gkm.sոwdkvnf��,%u��(.��⓶s�3������1��xeG����/��X���Sªwy>8?}�%��A�����^anS9�z"KG����W=L�<2�DT*�붛KȌ�O)�`�K��i�"v��w�QR�݌�|ͭ�z*#���\�!�������K��'"ڭ�6;�P3�-����5l�2��t����j�s��̜��E�=�Ѭ]�7��Ĳ/a%4ʥ84����n�,#�c����\l�y�&nzۡ�m�-�7S$=�>�� XW�����p�'�0%�$i5����O�ê��*5t��oS�C�-�2��Y���@��}�`���'z�$��S��t����sGb��J�yBM:�ٮ�Ngz<����SAa�C�mLpm�^�5��K�ل�^�dNV��A/��Qb��˸���)���4x{4�u@~K�^�!��i�#�L<2ס;�7_���k]�E��x�8l��)�{g?d<��4�	�kj^f.�mU�%h�2nu�|�r���GJ��F:ͰA'�hX��n"u����6��x�A7��AK̄Q\� �:Tխ��H�/�N�jkeH�+Ghڍ���rxmw8߶��2�y���F����S!�.%�_�P��;�t��v�R���
Ɩ�>`���'�dN��="��<ꋾ��+w��ٝ�j���cy���GQO�}W�U��Y�R"�������dk�[f��L�VzfS�
�]���/��3(y��Dc���S�B&��c�c��VߍW4����;u�0gC�=���Ҧ�����f)�����C�"��vokczE�^ԓ�~Nf�W����sP/���}!�wh3�`�����P�9�PC��ΰF3���1��~��V��}��2'�Iv#��v��C�HTaOK.a���Ms���t-��7`C��qn9�7�,U9�v�Y��2&����3P|�C��Ⰶ�{1��c�Hm�uT��<_�T7�Dʬ�]/�pT�˃���G
���ף*yՒ_�^����tG���KPp���?��R�d�ey�sgYP�ΞAp)��'$���7^�_X�hO�Xʊ��u�NP�mǇR�jЂ~ka�j<%�y.�g/��ٔ�9.�� 3 �gE��f��;co]�C�ˌ��v[���Y0���:!Z�9E'V1*�Ҩ��5+�i�p��1��߿)�e�_v\�@�\�%�+�hn�Ķ&���Vnp���SS�A�_/��فf=��˗=��v����۩FH�}�Ԯ�e� �׺��owKWs�^j�I�:`b4<�jLm����FG��^��7Q���-��u'g2����<���i�_�u�4Z�m���%3�B�8���B`�Z`S��SlX��Y'�b%9��W�TS�oD4��0&D��w��8��
�-��9�k�^�cZD8�1�[,�4�Ϻ��oQ�.g�2b�80s�/[&mk֙�=���.�d6\
�o'ې+�!��r���#�)�2�|i�g^���po&rs��΄���4�2�X�6.h�f5ٵ�}~p�Ѓ��0�7sЗ��n�Ŭ���5ƺ����
��Q��Ves�U��^l� ���7���C�K�ל8�,7v�ke�����l��ڇ�=�-�������zw�Y��N?����X^#%����,�=ۿ����޸`Ԛ�	s��#�hL��vk��"�ׅ�̜q�_�k��2���@���6�2�[�N^Z��sD{Zý�Ph3G�?���@|.hL3,���q���J���5�c�;N�Z�U8:�5��^�J���zf�0d=0\D���3\
�Τ��y������ba�'U�.�9�E��M�u�i/3X�zVB�p*_�ݳ�"|�<'��0�o=;��dh�o�)�(A��2\�2�ކ�����+�U;c�ȡ7ko�
ƛP��PV^�:�$+���m(W�z��w�+N��P����Xg��n��G�Q|��2���|: +���q���TpT�Ҡ�ފ�}�k�qtF��H7�Mj+̀l�
뻶!�׫�� ���-2H�fo\�a�?pt�xXi�#.��T:&�׶<� !\07l�RM8^f��U7!쫋�SQm����؍w��Z�}s�%�y�S槹}n1`C����ҹ�����y�w:�6_-�Zݳ0P��C�����/sQ�J�Xj�Gy�N��,�R����7�#�K�7�1Sf_R��m�H{K�9V�M0G0ӂa4�G<�lc%bv�����%6X�!2oU�"��d�m�\���ٹ7���.%f���g��u���\8�"+��+�^�`$&���k���BcƖ�L'C^�����e:=���LP��w�9�^��xOV������|�A��=| @�QB/aM>(��l���oC�<z"��܀/Ⱥ��ƼQ���������֏H0͓�.|р�'�=.&�$q���|��ī+�f�0�~�~�R :��5{��0�h���w`��C�2��v�^���s�!����8@	�8���>NN��k��^��->��%�5�K�5'�5C����k��_�o��Ͼ�j4_���"���h�R����:�0��v	�&2�Gs�Gj@W����x7�{���\��(s%(0�NӅ#D�g�e	YzySS�D�5r�E�f\^z-������YR��gT�zz[�)+*[Y.�;希����r���2��[N��g9�[��ۙMr�F��ξ�Km�L#�E�U��5֪�����>��¾���W��[�Z�qM,��� ����8t��ꘖ�S�Z�L����J�a'����r�ʼ�}d�_��]uǂ�H��]pQr����(r��U�e��L?�Ͷ�Y�l�hmG�S������nCǌS4W��m�ʑ�Ǣ`i��c޳8���3�<C���:�\�nqјс��*����C���CŚ���Pv��'6Ǥ�x v��=�D[��ptMz"|���/�j^3�(�gt�afS�"���>/��oz��Bv����H}���OT4��޶��EC�C7.#�ĕW�A�=����K����&��'�zǣ���4��� �5X�8����o).����˖-}�v����{�V�o#	g�塈.�Dde9������W%L�ge*
�|�fqnv�����W�ߒ��B���Jg͊��|p8W��P��H��j����kϧ�1y�V6��p��-9L�fo=��s|�{8���ѡ���������ј�oV�^���t����%�Ϣ'�H{r&��Sl���%�2�b����pAV�50�?�1,��H�2�F�[�[��:-�=[ۼH01^(�UsUU[Z1���$n�3�Ţٌ���F��W�`_k�L��"��{��n/v���/��` �	t���W��Y6f���X+\��O�A+2�a���E��`�ʟ�mK��z�Uy>�Z��`;�Ե��2�m�fs�& o���y������;��5P��5۳\?y�Xg�g	Y��ވ��9w��B]3�Lk�Ml�q��ȸu�^���ME�vXؗ�C����BF��kP��ʹ&e6e���Aw�e'�I���k�9�{V�5D��Y�v?f��{%�]Q���E��p"�9�jc�l��5��K�,�n�E�?!>4�{�A�给ɥ��'���N�9��W��a ��"�'ֈ`��4C�-z}4݃�)ƪ��L�!)qL��?LO �����^��q�?���5��&H^Ղ��@C`t�~����k�u�0���L���0�������&�
^�oIo&��`�Ʌn2�0��#j�wf��`�70����k�L7:&"�vF�m�cI���k{.���:|�R)hs%�:�L�c/��o��x�~�hW�`���ߙ�tf���Q��΅�[�B���.����b6��' �����0��;4�E�7���1�Sզsca�PC���3��� �GJg��s�`c%Cv�^Fv\f��q�b�lVĭ�7������Ɣ<u�X��y���%�m����zk�'vG�^_P�O�:���w|oQ^�ߍe2��4~G�	{�ns��)=�z1�G��X���j]��j�{5��<��`@�k�ڂ���1�D�Qլ�u��bJ,ޏ�� �%�5�'J�5���m!}�:�L^�+�"���-؏X�bl̽T�b�כ��vc�<�	y�hgv�{��� �?�·$�ȊW�<��"m�����&]��o�i���l�w�`0%��c{�d^�5r����*�	�tGR��᳏%��%��8��!��%�CPH׫Z,f�˵�hO������7D���
y)��ƍ�~� ��j��
'$f�TV5���u�Nm@�4�V3юoccd�C�pͳ�uE�/F�f�)׉�=�J�o��N�'�X�xd���2ok_,��u�R�
�RXKo�d�ź�)�Qh�=7}�����z��t$F��(2-�R�<�^�7	�����t�?x9oo�
Ne)�ODM��,�;�;sP����=��.9�-��-�����ސ_Ū�A�C��)��bE�iޥI��k�,a�	����\���M�q���s�W:�޶�� AƘr�xLx�"�����ޙ�lg*�z�d�u�����<w��L���y{�["�ع�n��M�fng���p�݀!���B};|7���
6��8ař��1|P��-��6�V߳���P�*z%�W(�����o���#�@�`э�ӊa��ѫ�r���l;����Z�~�4/�o[
�*�
�cVַ�����>\�'���ێ�C����¤�T�i���7ckz�f�o�R�,� +Y��گ^�cj+]H��bvhk@��qqv������r��ͧ���Yޑb�:L<�R�R�2�u��v�L����И�pٝ7a߉��%V�'�/��*�Ȭ�� ���m���J����{X�,㟛���ޛ�"�6��+^ʂ\�j#�`�+{��\:D��k�C�T"�U�^��5�'��!f"���A��19�0�پ�a�Y�Pp�����v��-��6V3Ɯt<yݢ_���my׏@��3��5C�.�4&�no�L%�'[���+�$M+�W�f���G�)��y�ݯ^�F�PS��j�����W��w��KK�<���e���݁w{��0�۫��� ^E���^*>���>D[.x���f�\Ge;]�`�ơ��!�r�Ed�{j/�5�^A!���J�!���O�2�7C�:;@���n�u6W����o�������ב�Q�5o��ەR��J�:�(,�o�Q�yK��^��d��<M�χ�X|2c�htS< �4��c�q����2Q�͡��M��BeuL��u���mއ=_.wRԽ��C^��W^��g�`1m!8��B`$&��CM�mئ�ó)����kT�
��{���(��9�	LT"�]�6s[m�>�㼆�t��	�Bt��3���L]�͊���/N���lz1I0՚O�/�w.��u �����]��řv�b��&h�k���;�%��ZM���¨^�ϳ��%�*����@��ђg�wK��+U�
������c�)����b*�V�*��cA��L�O���������   v���\�!�����>�wL��Ĳ.���LhO�7��1e�#��a�ׅ�Z��śh����cm��pP�4��u�.�dމh_Rw�y.�h�R��n�c����4��6��S�Lf&�D֖�*��,�d3&�B9�L� N�s�fc�ѵ�S��ܝ�V���XJP]�����n�\4���������x��waɃ�֐ ����T���	�`���Y�h�LY�CN�Gz�鹃ف��������z��7 8�Û�t�LR�^���S�Z�X�kq���^�5۲*M�s�:B�1EοsԺWҮ�ht[�!�8������?X�v�� ����?�֓`�<{#��i1�2���ϧ���z�׌Xgc=�����z٢�0óg?싡ζ{���a�J����0ҫl��E��x������v��zA�ū�C���.�q��!��|z��ٙD{;���Hx�V�%�-��������$={�Cy��OT0��J�Fb�b�]�w�6̐���Cڸ�}�\2O��z��z7�CZ}��L�}�J�dN�2i8q�|��S�����Ӿ������)��3��O������O-��\NY�%��׷�ez��<2�~yB��׳���UӁݹQ���Rx[(u��ι�R�q�6،G]��P;Ɏ�}�7s(�v-3��N������>��o��W9� '�z���&(^R�{w7��כxiזx�	��a`��I�::�lMO����i\�3lI�Qv���ʸ�Т��/A��a�@��6->��V�S�-��â����U���{9tCH��٥��\�vd=�1�D���2�&�Ji=���Fc׭����k��PR6tD�˽��z�ڳ��X;2[B#����n��Y=\�� ��|bY[�H�2��F�U��;��<�Dp
��� o�b�s�Ҵ�WҐ��x[r��| !��y����b%9�g�H�4���ϷІ�W��]5mf�(���޷���{W@P-�4�6צ82��`��K���F�r�:���(�g=>�M$�9i��T�����z�O����"=D&���ٽ�j/xT�O��M��x���p��Z]=G���OZ�)�jM>^D	��?`a�Ϙ(֘r9���-z�4ݴ�5�U�jd�4l����l_-���3+�}�c����?{��
�c;4~`��0쟍q��h��)�v95Pu
�M�Ge[]�IO͈���
��+�[���CA�y�����P>������Vٹ��x�뽐�T1N�\����^42��w6��+�f�K��U�y�j4��B�ٙ�>V�K{I���#�C:�/rY�.���3C�-䢅KF-�2[s�`���S4NїI�,A����I��:��HՌ��"�J|'m��o�`��Њ�.�xro�V����� i J|t�rUx0��f��Qք7ثmgu�Еa)�ʓM6���mX��ܙ-�)������h�'x��(`���P.kx�������o]h��Ɩ�E~�^E�p�3�,b���j=��?܊g_79� �r�ʟ_,��j�]���)�VV��U�[/�I���;�І�g<|�T��&s�|�b�0�	ٶՇ�3��;����Sm�y�] �kR���o���au�W��szt�n֊ƁU��,֌lh�Mꙗׁ��T}.�<�mgi��Y.Jn�mԱ(	�dn����l���9�W	�j�q&�^�,���wq�w���B�z�K*Ţ��a��5@�5p�ŗ)��)�����Ȝ�3S᷊���=�����3b������w̡x^��Q!h�iā���mLdur5���W#��"[y�
���8ta�P�a{N��{�:�.����vve�	�6o��ܬ$G$����}�K9%Ym��'���:c�@�-\�r�s7����W"��8ޝ��Cb��>`2�\�S��N�N���٤�������cpP�@�tq�z��|�?ޕ�J��#�;a�F��ehҗʹ`b�nʺ�9	� ������vP�[vNQ�쾡&JS�h�oN�9y�k�0Ѧ���o��]ĵ���@^L����6wj�FY261��W�W��<V�¬�:�j��*��W�י��ѳ��Хom8���P��&9uo��㯫�!�0sz�JC5��s�'+�d��7�O@�/9x�+;�L_P��4D����G��Da-�Fd����;�©WCG7���@L�*Vgjj���f�՛��#��&���6_!P��Vkr�:����R��lEX�����L����Me�"�g.��s"N��ZL���l4˭����9݅S-��ի@�#�hIiC����k{;n�eW���s�i��[�B�XX����PW�T+kW�O���x�;]��(jV��+gb$ �s'��Nn\;�2V��X!C��fƵi�_}� ����Kpj�������C
���s;��u[eJ�3���Wǁ�)]^�t�����OxD�f���'��:�<�va}�\#�B��C,�� �0��SG��b���Q$�3q,��&F��;T
�t7͉�*�*v�ON�Q9�$�ۮ�	ұ����˹�f]�y��zLJyιt.P@��(�4�(�(�R�!mNMv��@~R+n �,;
�!����z=lm��Q���{*�)��*��i(��j�4T�i

)�I����|~�>>>>?�����<H��U'MEKJQET�RQQ5@�������Ǐ������������|9���*��&�h�9:8jh��;�HUQ�4U1E,�E4D4Ĵ����*)iJ(5���B��
CC������]Grj$�@�CU#��-�G!4-	5B]lAUDAB�F���i� ������e��@�5EQM4=��H���uSL�Q%	CKAAAKM40E{%S@A!QP�E.��A��CTWrw	�%=ɪJM 	�P{@B�V��D�����]���r�V,v��mgS�i�31w��q�J\�e�����F+ia)VәN�]|=����9���y��c�����y�����{�zB�uWR�]�`���;k�xf���еa̖A�k,{���g�o���G�Uά�)�X�������!�kSVY��9�}i��X�f�m�}�#k��o�'�Nf�W���h�����Q�k��o[�?W�>�*g��w���;F�c�ql�{v�k�a�;�h�l�4�w��@釋l�ܛq;C![$i�m����8���"a'W1m����>���zL#�v�TV�~�f��g��z�� �9v�Ɵ�qvWҵ�%e|����*�SE_�(?'u�w���(]�o.��rY�l/u �}Z��	7��fB�A,����z͜e�)�>zw�X00��g�ꋕN�o*Z��{�l
�f�����M�;��>���	c^K�����eEÜ�֎��r��:��A��8��צ%;O��g��d�羈A���)���J�QaM�]��h�|U:S�ׅ��V��Z;-`*�-\�uh��F{p0:�U��9���'.�m8�;�|�o6y�k�d�s�HI�.-�-�ȶ�]8މ/����e��Y�i��>���R�}��&`���/�R$�m�6�
��c6"a���kU�����J�ٕ]�msٗ\����.�r�ҴU^�κ$�R�j�4�-v)�,�*=�a8�vlqr�=��[��9���t�A�����W�H���˯�"3��A�r�������N{뿧����x��%���7�3e��-��@AƿC���L9Ҍ��ن�ys��?h�BX��;H�)��)�E�.9�4�/�i�f�}~�_c����z65���K��ڎ��t%�k�ƅ+�I�U�\��-\��T:�]�
�z���C�Zf ��R��W�L�saCB`��}iz�����f�I�|Uk��M��a!=��8�se�=%q���[��*p���z󷚋��^n�cB`ke�H��d㎰_�k��2�bۃT�MA:2��Tr�
�Ė�{�zi�>f�69��s����kVrT��f|�p��.�6Z�w�=��].�i� ����0�j�<�w���x!0�L�9�0|�Ɂ�T�s�fV�A;OF�^%�z|�9瞼�v<��0�C��ju�|d,�_��Oh�����bI�eS0�ڗVbޘ(�-��i�a�-<�@$?�˥�|tE��xc��	�g9~�I�gE���|Ԇ�<�|��v�>	��{k��>��C�P��9�%r�"_�K�O�}�J��^B��A�E~���f�x�@��S�����d'���9�붙��!1�A&��/.嶠������u�;��Ȓh���C�ʕn��Uw�3Cjf���5*���AS�9�����fQ眐�*A��6�f�3)Z������}���W������{�ͷ�
&ap��`<2��/��Ur'�>����}���D��!s�;2��B�f�e�S�K��u^�L��9`�eY�(��VR�x�ix�\�ڸUm�sX~"S` ��"]m]7>~���a~��KM��O��k�*ాg��<�T,_Ɵ��}5{�t�c���������t"��f��؇<I~�L�	�"�F�c���xOV�>��Ŵ'H>�M���������oq�C�}W\�/��z �<�y��[����:�y���?���X�2�h�\{-�6��EnQ�׭��<潜$J�:��E�y��E�ئ41u;u���v�Km������hyQ��s>���7M�F����������jm?2N[�����#�\*b���[�w���H��0�/2��I�hLJuBL��	�d�2�tS�m
�V9�a��F���A���yl��������;n����O:V��ix1��5f>���{?�v�*`NF��~�sO����y��t�z�Q_Rb���۱�c��̩��z���>�X��-M���M[,S��ȤV�H�5e=f,LO�>�����am�w�m�<�^gC�`�|��5}�9��*��Qp�º)����nE�Z�;��b�d�`�u��t7C[� Ycy���K0�������~�y�=�y��p<=��)�mP�����:�n��ێ4�ߙGS�īկA(-+�ZC����@fp0��=��4��ka?X9n���t^�.�퇼��{(�X/��Šv׉���lZ��;��z��3��'U�װ>0�S���/�^�ҽ�ٳ�!�z	\ZOT3���7 ���Xg{?*���KF�VU&
�_����i�z�����ui�Φi��,ҋ��&�a�lZsk��͝wylleZX*�pa����kC����ʫՍ05����9�kg{��ff{e3B�3��1�����؁�o�ǫxT:E;��$z�"����m���F�F�gκs8��RU��!6o�J�҉O�J�����[ռ��#a��T,�]1���^����RXy�l{Xp��\���A8��%���#6����q���L��n{�UM���
ok���;�f����S��.	he�<�>x�Js~�S����}/pĬʓ�fi����,��WG�@0-��f�������f��q#z�$��S�}XIʺl������` �S����oz����ј��u|������y'��s�\�|�1+ԞL�P�L���	P]��c��r��e� S�Yw�����5RdC�l\4A�F���jgw]bݍ�����}�%�O�+˱}K����5
�;���+�F�B�@@�!x
4(�W]um�(����A�r���{��5T�9��̢�5b˶?�C�A�9�hLpm�{<�^��K�ݗ��vuU�˒�-0�L^����@��0�������:��`�LY��f�u�Q[U1�Gf�4,��(�ֻK���5�Ƣ��_='�q��ݨlc;�6�y��`���,���Nni�k������B�R{��,pGu[^�$��b2m��W>��ͪǷ	W�b��=^��X��Fx~w��!a�ö�cԻk��B�,8�V�O�o �@k�_�?�q�OR`�"�&�¹�9A;\ߡ�/hr�C��vֲ��'���C:�pm9�aŜvB��s'��m�SSX��֠��᝼����ڰ-10���`c%[�^Fv�����v�sU}����(f��dK�q���u{J�3����钽�� �j�	�L$��-���z��rr�Ž
�Z��y������;�'�.v���F\��c�bz/"m�4J�t�w�XP&@"1��ЁG9N��[l�cr���5s��ͭi;x8�rnjK$����=f�2��1�={���O+*0��w��z��;�{I,��u8���ի;}E!ᯣ&�u��s��֞�̬2۵�`J��;V�I+���G�w�P�gi�Ǉ3^���Qg����e��2�c��s�7�u���⏑Cy����nVtǛ#xz2P�<�f�O���[}� ��{�@����YEU3�6ٞZNt�t���v������"��**۽`���c��r����V�ю���Ͷ�Ie�<S����̍y��a�%��Aqub%8������M�0��e�|���Ī<ԭ��m9cbT��{�&x^�`Y{N5��Uq��7��ȸt���Y�H��xI���$��-v�y�1�����n����*nU��F�0��Шt�zA|k�H8�Co�_S5�ν�@�].���,���/ۺ��5�X��&*�?8�e�8����,�׃�[�	��64Ð��f����8��0/�j�'y[o��o茔�|��Y�0��F����������aT��	�N�8�9�{7,ͬ�B�H�/<�9H��i0��+���r�����ǽ�[�8���"��Ϧ�;�=�;�Ѳ��ˠ��d�����@���/:꧍70\Q����aV�y��WZ+�uj���jܙ;�B�7�?C�B�����|�����)LlK@����jÙ8���V�k1θ�|Y�v�o[����@��sg�Ƈs&<�F�5���ve��Xc],�k�ʍ�����Gw�HŘbܸ.�
q,ٺ�o��i���GWd�i�i(�7;1B:����Y�nX���&��ׯi2�V��e5Z;�u��{�����6Y��`�	"g*i.�b�͸*�d]N����X�7��75��Df�g| ����q�x���< ��-7����zP��5�?ء�r��nj���Ɂ���xm�3����K�3[[w�؇'�9��6����l�e&�%ٷ�30��-�`��^�<��lr�u�ji�����g6èy�L+�Qm�vY���,���Cגh7.�l:"�P�xcՕ)�'ؚ�wM�����S��fM�Oz�ۻ�y���}sג�7�g͚Jh��ا�R����_0mS�̽�k���:aa�s�����{��j���UKcR�!s�tnnsk�ɟ34c�9��h���%���.b��{b��!	��C��q�_.�-�ԥ`w�4��k�S>�}�
��FG1�F��>R3�aw�;��p�L�G��~4�qҺ���y�/\q��7�*��Kru�t*���rB�LT"�]���z��	�� ���- ��a���V�A�v�ǂ�z p�|����N��bi�u�cݞ(�a�â���1�Wm��J͏Vt��d$d3k�a��n�!�.�/���ʥX\ʹ�.�nX�m\�SNi5Ng��zo��og�^�a��3gVǢ.�����y��Ko����Ay�*�F�}����"�q�ܠ,p���j��X-[|�;J����;w����/�I�}� ʔvЇx���p���aWS�WjY�w25��}?��9� ^~z����~~~i�兏�hiD����!]K���~=�f��wV�t=Z�O�ݙ������3=\gm��1�ڕ��j.%ߵ��݁��֑#[�bK�����r+[����E��W�}<�nk�u%�?n������Adi/����!å�G�í~�1-�D��e�<�����Ӎ��(N�k
�ekߊ�^��+�iWr͵�l��0n���첊v�=q�l�&�&��vf�ȩȦ��1�N����3�ǠM�^����yu�j��O2�"��Oa���U���q�?��T�Db��x߻Ϩ��q�KϏ���-S�^"Ls�SK/j�s�IA;Q��D�tý!%����=�{�+���7�XCN�z	\Z�<W3u&��ƟvT�-�#"*�Ȑ�p�|���M>�؞��[ѽ�^nj��LӚ��Z �P��m�F�T���ˡ���w ^M��_0�ǖ���)�@���P�@���V6��\�]�/�Y�e�Wt��%8i�{`�$,�`Z�;A�6q=cռ*"��`qm�`Ћ���0��.����{y��Lj���՘ܳv:Q�]*����m�@��H̕����7�JF�2m����i�E N�=f�M%�K����*Z�:�p�y9p����'""�֊������:�-2�R��9H�ʈ�Y[��q���3V֗L�&��=.�,�71)���� <�^q����Ǽ<=�7B,T�S/W}�Z�z������lr�5�����`y���o���".:�ް�s:�dqi��Д4D�� f���9�"��[W�� ���d_3L��Ɠ_Dv>3lՑ��T��d�U*\��{3��[���2B��f�r�g���&�O=��(��T��H�9l���J�H�WnTv����-̽'Z�t����so>a�`�"��zS�6��S�},�_Aw�F�w��vM�܈ٓX�ݖ׺�ڷ^� �E_�Ú��LYz|�>����@D&�~�/g����]�=7<$� ����N� �ct=j9W�H%�jM#��`y��q8����|��e�x3������TsM\�8��lf�k]���Ad�c/A(�v�(�q�b]�=���#�l����4^���m�~��
��;k�BdN��OH��궻�����#&�UG�ʪFVŻ��?k�\�&ٺb��S4oV��3ᐠ�{��ͯ��]���ȥ�s%�S��{�}\fKNլ�H�]�L՚���z�C��`�2g�!1i����.���ȍ���r	��,Sq�vQ����0F�@��3T���w�Ư�����i�f�ϣ���F�Oݵ��f�H�vZ�̈�ҪX��9^��=�;n�#�=%��
K�&�W�3���Xٶ��%�0,�>[[{ȫB���suz޷�X�s��=U�91�}�xx
��{���p< ����ccv�?��\Ÿ[����6q#��s;G��D��701�����t��7u{,�B��"W�Ms�x�v- ��q'DYz�x;��-��D�N�X`�蜃����Rӯ���輳BkzQv�%8�5{��i��5��y��M�$T<�0&m�OBK�����u�s`V�<�2牨�����t��B�Id����=��T2��{�]��)�r�m��n��[�	q�w<�1�L܂r^i����(�s�ϥ��W"�l��h&��$�%+�����|���W���3?�`O�D��1�\:�=�-{��Eʞp�b.zd��R�%�s��a���k�SWvN5��so��$Ao@Pd\:N�{,�$_Jn^w�H�>����y�v֊}�9ȴۥ:�i*�	TS�z�˰��г�N����i��s��Kp��rm~E���ߩ|̃|��n�2�qx	��7H��W���w�xa>����	�8q�e�5ͱ�~B`Xoc^�@�[�7Nݓ=o)�E�"�ʥ�^��́�ˬ��J���qq:�u�s�=GEX-[��[C��:n�e��Wx^�pV�$:�T�fbV�HZ�����U��3o�`���;8���{������n�3U�H�_wc�.GY�M�M^T�F�h�g$B�ɹ2�y����j�TM5��n�Ff��0��Dp����|V��q\%�)W:3�
Lu��8��W.R�-[�,�;�&�S�V6P%�i�i�<fM��z�0f�����WI�������Jv�3�u�NvJ���V��7;xӌ�O]���ۂ�ynwFk�Xk�5��LF B����L���Z�O�,�6��da�ʺ�|�"��O��ɚ�D�5�;(�w�"r��S+���9�0�}��f��Ó������W�Q�ȺM�7 :�S����U����ұX����d̵�ܥ�H�&����F��Dʎ=�w�e���qݴn~y��߮L��hj�]�Y�r����J�����c�P��|LӰ���JeS|���+h`����B��q �9��S�(��y4B��}��B��wZ {��p� �ѧ��z��(��1��m[W�p�@`���B��S��=MY��
�$��&��n2�!����+'Z1f;��W��wNu�G^���D�O!��.�����u]4�w^L��R̬t9��� �G�]�������a���.gzsJ(5��l����	,���w�zḎ�kiQV��`���$E#2w�LR�R�T�Zm���@ �+WaSmr��h�����ҵ��Vwх��\ʷW����$Mq��˾�DH[��A+v���.�,�����uou�*b������� R���lVd�9�3�H����'��NJ�?���J0�f���c�]LXW$��ER!�	��n�[+]���%�#I�r��:�r���;mAҎ���Z|�m�j�ߣ`��p
��;21/o�0��N�c���2���C�:P׌�ݱ7��v�ʕ�����z������]Վ�x�WA��baKZv,�ws;N�Rd�*��5��X���Q�/\Tz��Z��]�}S�m-h*��Q�5��VG��YOݧ��:�n�º�_v]r�26u���_.��n���N+�|DU���c{u|E{gf�xH���σ�Wӫ�o��[��s��ci���:�����5���է�1)gFh�i�N��csL�gf�s�:;�&V;�n�Q�qK����cX�h�e�ci]V�5P;d�����]SUZܨ*ʮ���VN�d(B�0�ۺv�TI:UxP���ٽ������P���F���b��gOiV���Bsݙ��)u
6�DF�ouʃ�啭PK�c4�x��e�5��Cv�*70%���F�9r��k�vm��-��%ā�VPB��K��1�f}��zrӥ�Cz�@����\��C�E	ر��}��)j�)*���tM%5Mx�|}>�������r�i��"b�i~X�(h�)��J@��6����������������������)(b�JZh	�h(��AA�hJ�����B i�i&��JN�EPP��ECA���IHPPD�1	C �"P�R�P5M��$AC�T�1RQHRQIE y=Bu-	EATĴ4P�EBD���EPEE!@e-+@�@P�@��P�i" JR��B���J���KmAJ�wV�.2�q����f�%��f��V��~��r�e���e]��6�_B�����ˁ��M+�Z�@-}���W��}����� xz�����Ұ�~Hq�ݐnO��_���;��
�2��W(��RX�-�a6���#i\fӤ/�ϙ
 C�`ɗ���rxh�Y<hY�9��/����]<�g�kP�c]�PND!�{�
�p��U�[�ɡA��
*���W���0&U遭�z�Z�2q�:Y!�:�-�8c�Ykb.w�o�At"��E{�W��m@s�w���`�y��F�4��s�R̺��M��@�L��Ú����;>f���[/N򠭗Mc��ӔMKsqe�Pg=ϸ�����;�TM�m1O����L3uY���4�&�E�^���_{~m
�u=����U�2��4tK3��7��Xd%xQ�y���ov��Ⱦy��z���TG.�iD[-�ш��D��pk�8��L��%��ͣ\G����|�p��Ƕ�f����$<�}s�P�.�U>z'�g�c�~�#��U�<뭃u��\�I��ė�5�ה}t�֍�\��rzMs�*���N�]�/�Pk���<��o<�ڈ�=�����)������Z?~�!��w{C�����/�f��/�����`�1Օh�J�G�E��U������_���}7� ���:e�&�(!���)[SG�N]�y��w`�N��}��q��|t�X��'Er��~�0�p�W:C����]nn��G]����~?��� !V�.i�n.lf6#��<L�ʭ�¦�e�zw_iᶞ������S�����ޗX+0OHW�W�7����LW�x��<��2e6U}���hc�o�p�?�JT�J	�����o�0�e��?C����
�פ5J�k<K"�<�ģ)�kθ3����4x������[�z	ٷ �,z�A��	j�����(�ac�J.��)�u�A�����a��<�a?7����vB�*�π6Avlk���L� _o�i;��YUѰ�R�}Yn��/�Wp�9OL�Bc^�%ߚ��w�v�}�S��@`鵦8C{�cO��S��|nF���������nsC]F^�Gs��t;��@����ېB�:|t{��:�3�۲�!��4�ʦ����M}<����l���������3��ʹP�~�룯g�(�%�զn�v���;3e��t�9����GS�gӏD�4��,ƌXgc����M*V��{HfB�@x���y��{�d�"�C�^�/ş��G�H�%�j��Ny3?�Aﵷ��r�%;�.�{GJF�Mx�x�ι�>rԇY����r]c���k��xv�<��n��
A'/1JXI_�9�;�\n����$���Ɗ�+�m �sr��/�<�nQZ�5w*l���(=M�T*��Rg>�t3{��]=�~�?����UG�{���߿E���67�b�v%�89a���*��/��oz���6��4�A!�H,�l.xZ�D�M��@�Ɇ��O����dAii�3Agkd�<%�ލ��ְ�w�Elz�(��Dl2��LҵN��|�R\�ux��~P��������~b�~x�|�O.�2��Av���K��)f�e4�q�jH�SC�����V��"���HY�߯���VO1�_��g�rf��^m*n+��Bl^��&�Ji=���z3�y������G�9U�FZ�0�ᅻ���=��b2�k� �W(�E�0��WIj�.�M�tDj����=ܸٟ�?C��&*۬]k�j�L�	O����'I��Nv��������{�j�A��{Rkk�vIj|��TK	�qmP��l?U��_Iw��5�d&��Vlu������tr�tEs��7H�Cs7���1e�>G�C�c�	��86�_�U�.�;m��ޮj.�t�M�M��Z~Y�R	z�o�u��i����4[,kX��
+��/ �7��^��V9[(������=��B��k�7�N��.��]�t]0�)`��={���e࿚¾����F�����2��=J-w�o`���C,�ף�}[w(����K�Nuͬʀ%sWN��b�h�/R�R密6��c�]���,��z��T��B�|!����3o�M�7�s]�6Qx��5��O�����8�;�{c�o~��OU�Y�F�R�(2��!ݘ�����n���k�oJNZ��ɷ�W?g�v��o̩X���~����x^��1[�5ӟ8}�r^a۽С�K��O�MW�2Xuݓ1!��>��{�x`�ڒ�ĶC�Z�W�1��T1��?��R!}�P�:�_��X�e3Y�t2�>H����D�<��y�V�u����k�|�����mx��j�~娽�q������"ac���v�[E�n��Cb�G^��Of���Y�����^�.Ť��	��\��x����)�|��hᑌ�k���6<��S�����ff�c8iY��cYS���b���%ڼ�d�#.�o�}���+ ����`^6D�g�Ұb��9�=Ŷ'�5s�Y��>9	7�k�o3JZ�\��3��5�w�t7x�)э�|Qd�I��B���K�:������!��D\teE[.r�p;(�PY���3.4�e���������_�;gK�WW���k�2���.�dՓ��D&�2�Cj�4~�Ό�ථ3���%�r��e^q�+\��{�1��7�wOl��.�b�l~��-��9#|�]�0��#���EV+B�,ͻmn<��{����PbVu��14ør	�۳�N�.�S���7y��֮}�bk�F��N�L2$=��Z�y���ý��x�����U�8©~���xM
��QaMK�q�uEë|g�彡A�u0����f�v�4$��[�#v;��������ADb���&��J�ג���]��0��Шt���t��X�����LQ���E�ِ́��z]���e��&�PLP0'��QT�l�|����p��q�]u��m�蠹�9	�	�����2�_v��RS��e%�,c�Qh���+�D��ۉ���0.������������J~�Oo&^�4��_�\�y*�J�y0v�άg������qe�Ç�3���耛��4�+�AR)s�X��ܕYk{n1�����U5J�0��v�b�١@�������#[0^��Z5AR&Aܫk��+�pR}��I�zbG0��'Z�=�~�88�3������j��Fk$<������s|�7���:��k�C��R��@��^�9��x�`>t������O�<�f�]}b�QK?�8���v��E�/���7k��i:"����]ݷh*�@�B��?70�m�~jn�|�t�いj��	ݎ-G�BS�_V��j�Nޥԯ�܍�K�8vv�:$�t�ޝ9�>h�o!S1%kWk6�����!
�wk�g�Bz[�:Q���r�`&��vvwt��o6;����+��y����W��r&s�}��F��[�ǟE�q?���!�W����fo\� �~Ne˥��i.U���c��b��^��l���O�tg��3�Df00+ӻ)=�j/���k��[o����Uk-��v�gwf?��őCwg̮6�5��<��x �Ut~4n���X']d�`��*��N�Tb�Y�L�|��Es�}�fW�g�%u���8�nb��lS<!64��i�Ŝ�� ��k����V�g�~�������r��U�B����Ӻ�Xe�C`���Q����4ɔ�?�~��w�]����^ϸ5r��JdY�Р����3��V���z��xO9B���-��ά-��:�z��;�`qM��L	��@"o�zF��N��K"�?8�c~(�a�P������U��ާ�~�N{r��S�`�4���b!0�z�!�o��W�]���E�S "��TK4b3��zT+���=��^vU���d@����(f֘"t8-���B��4��Wd/>5�-��ƫ�[��C��g�|��R]��8�x�aҼ�|��`�4:]KG$~?�����?U�h}ݗ,p���ph+%@4@�0����U�R�=�~%���8W��'6�u�+��Y�� ��F��%��˔�<��,�	�s�eY�
8����(qկ�U���A9���F嶦�2����r������aM�u__P���ܙJ�y��{��|o8�lu�#��9� �vC.�G�4(��;�a-�=�.��p�����sV��sשd�j�zp��PB5���3�UFU�u���`ݹ@LK,��M�V ����ײ�׌<���eu۟u�G�*�%���H>��C�����Б^aؾ��6��gM���1�Q��a�z�<L�Q7,�uZa�1�/�76����e��fq�
�B
y��|/bW���o$;d��E��x����;:��&y&Y�XV��^�{�^^�m�C�C��r��h|.&%M��K�:W����Vɂ����0"l��}�k��-�R֌�h�MT1m��y���Aiid�}�:O~��z���=N���)��!,��i��,y+��R]��E'��6��5���C �4��r�۫j��;_"�.c���?Ԛ�iso�#��m����M�,�d�9���t�wP�F[n����i=}��*y��)�6ۡ�38�Q^��D����ɨZSI�t[=�3���7��M	ʉ���Gg�$���x6?��&\�C��h*��?B	�Q,�ߒ3L�E��~�F��ܙn3_����֙)`;p
7�N�j踵����W�%u��\{iWqж�t5|��97�E��P���XU��'� ��;�Amǉ��Ni��Բ�����"���3��]39^�"�9r
�]7�޽K[/�gY���w�{�8��x �Hv����\)n� �dkX/�����dOٲ0]|$7�y�%:u�3cѩUO�T}Y��E�n������H�jgo]�����\����۞���E��U�[�,Y��us��,K;}؊�+t�5���5b˶?�s��SB=o"n�2�cL�-��=n]F����A�2N��]��&�~OI�H%�Qi^Fi��K�:B�K���yڛ���X��+��Ap�<6k����۬Vs�n׆x ,��e�u�`�_�H0�o�9����xB���S��_��Hm}�2']P��
n���m{Г���&�l+�4�2I����gM���{���7��ݶ�Y�̤t0g���<C�y�;k��.��7���s%�����W����`q߾�����l��mq�t��<yLZa���xp�d�Y�B4V�::�:��m���8-�i�\�4¼�@�b��p�-��;��<3ǴG3��|�&�c��V��EX-B3u�>,�琖�]�]�b�\by؃��ZI����������.���b�l]���5DClW�,3K��IVd棪.�wM�oi$��}{D�����0.�#�>�}Z�g%}%t ���s��y�� �O2�{b��'�H���hb�,*xx1�t]bJ�(̲�:ԫǫ"���6�[F`�Ȼs�'9p�x�/�����������rH��X�Z��Dŧ똶�u{�輳BkzIv��� �Ț��ִ�^m�)����z�f��#���v�\	�,G0���^&���m_��:Aƃ��_��-�i�g�.��s��3;7���l�Ϯ���,#�ُ,"*;쨫j����vO�Z��]�R3��9f>�҆vֳ�����>oL,��fp��g�	�q���i]:ɟs�)!��	,�N�<�����t�Q}��P�r�����8����g��AA�u0���F�s���N�_�����YY'.�dQR��},:��c�B���9�f鐢�n��P3-I��Pm]�
�����z�R�*S./1V�Qr��/�\�;�0x�.;�o���4N����"�s�q�2�{*Jz�r�d]&��75j-#�u;�̫�~�Z�kF�.x�㬗^w,����ppu݈n�%�?P�4(��E�Z��ԮQyz%!�����ޗ�S�����j"��≮�a��T(�r���/^��ƅ��8�����p��9B�x��ƨu��������p5H;�L֘׮a,B/�fu����7���-=Jd��$��s�Tŷ]�t��эAr*"X�˓*C��!J�M̄�Qg
x�]�gRp܂����k�Bŵ7܋��F!�y͑�[���+.�X&��?n��_������A���wa�w����+�a!=��ty������`��� �c5���jxMF�y<�m���:�o3�X㢠���Q��Z2��ϕ
�>}Z���v����¯Zn.���Bx���d�óVi0�s�%!�Bٛu�r�i��5-�yŗ�^�9�"]�{��U#-;ZyޗU�A���mՉ�mN�6]�s��
ė�a���q���tE�޾�jH��ռ�?OB��������<������3Ǿyހx?'7"�̊����N7of<�Bv^���؛xc[�v�
��\=�$�5��ןc־6��!�3�7�T�M־A�8ȷC��h�k�o����^��h��<,:� ���5��P��f%�\�Fl�������n��fP�`%G�=oN0���s�,��&Ɵ`�,ʻ{6�S�u���=2A�'�nƶ��ږ��D���!2�ZT)=��g��u�k�<4�{g`9❠��IF3Z��Y�C\Jo?W�#ͼ*��C_(-΄&<���,!��n�
��,�V'Y�G�?>���a�[YM�{}fo��ͭ����DwJ��H��Mu�m&�w����/E�릍���ZdjV���ɮ��^�s�i����[�NF��2������uwkO(�!Y<�v�-��>ݹ`�G�m)�]p,n�V6
�|�b�!��8Ij}'��j���R9�nZ��ݼ{����`�Gu�+nR�U�1%�Y܄�[@S��H�9A���/k%���r�k���p�f�`t�wôҗ�JK]m"y�ʽ��n�آVm��,�-I[N�k6QRb����Ek3\p�KZj�9e�x�.���g�V+{R����������I��١l�8|5Kl��)���b�l�]Y��{e�Eats���>�BUǺ�X��]�]F��0t%y,
h�aV�R^w^���au�B}y��a���s��}��1N�L5{#Q)��5�$�e����%CK8��Tu��S���GQ��f�h�N���uy�Ltu�lb��
�T/,� fLQi�R�����u�쑂r.&��/��=��Z���ْ��7r9����}��R��R땊��c� 4�4ki7���4^� �R[��,͜�����2�n�p�}ԍz�r�]-��)�PiPʔ�����hS��;��V�pI�ą��]f:�c�ٓG�%�.kL�
��J��,iir��L˼|d�](,��y�_>�S$��H��fiМLf�vB�jl[�r��(��ä�&���X4��Y-�[Z1n6�a0�d���S��H�,��u��N!)�����BVl�ն�2��S����ЗrHc��N��[���y"ŗ�p���WP��pt�N.�����n!�ړC�:�I�y�`��aOxtx��c�l�"=�x���l�"�8�q�/�ձ���1oS��e<4厲LT��]���6�ζe�l�k��nK�C��ywn���j}m*I%�y� �|&�w-�1
hQu����x���T��:�ˮ]D-��f�Ԝ�e���vEScNU�}�P�-�s'n���N���tT9\�#7����m=��	�[��S��L<b�1�C�����NS�E�VCw�(�.E)���$���z\��Y1a�{3���ת�ޱLZɍ)ً%���CU*�1Yil�n���fØ�5D�.RÍ�.�b�;B	OB�kfF) .�[��v�`�y}�u7[}>#d}.�	}-=n��.'ݤ��ٖlqh:��KF�vJ���L^G$ޠ�ۛ��)�,,Wcf2���)��XWr}��VVS��}#��uE@k��듨���vV>Z��r�P+��
��XjN�"��d�=S�.2,t6�왔�8*���04��3� �5f+����D�0F&���ԖP7�����͔���Iݸ�-n�T{��C/w	�%�,���XK|��Q7p���(��@ɖ��CqZ��'b��ܺ4����j�vE:�Q�I��������Z��aҔ;f�hB�" �i(�`�~?O�Ǐ���||||||~�_�d(J�)���:�)
S�����CDg3��<x������������yȥ�"h��~�i(JhJ��	H{�u�M'���P�D�!���ר�S�I����w���.���h^� �1E)m�)M�$&��ԁGQT%�P��R%1UБ�ZR��i:�V��RSA�3QE�h）���+HQIO�4�A@Jf���J�(`�l4�V�t:)tP's�)�&�"�J����q)C����P�79�[������l,���Ҷr�9�&'9�q���&��д�WY��\�]"�*v�-ߎ� �[�;�W���^o�߁��p��9�3���[Ŀ徻����<_�|�'��/�z@ޙI��d]yby;:��}��iU�ז���N�)`���{��L[��֏H�f�t�s����D����>�(�a
�] ū��)����Ŕ��(��=.�4��6�zhAC64�����ީp���Уds�����QTo���f"�)#���,ŧ�%�j���^N%�=��XG�:mi8F�G*{}�Y�˧�:��}��*�L9�J�h�2��;�ҩ��di���s�B��&��Z�,5�^`�\��l�v�[+��kW��Х�z� +��<��f�������|�k�а�4oV�����<��;s�H�f�y�6��&6G7��џN9/���T�1�M=I��;By�)�ņvR�fpB���Cξ�K�}���{�p/���1{�0�as���Ƌ��U�ȯN�d�AݎtK� 円���E�/x�Xޠ�(;�]6�t��������B�E�2����$�6�-�;P�+� AiiC ��{d�'�(k�,��5#�/��UZ�?��jң����M(���:�S{(��R��=n���y$X".*�+���R��:�,�9B����^��.��}YB��ʌ9�f��2�dcc�>.��uev�wYa[�-� 7�l�rj�t��I�]�c>����֥n�u��_�*��������f�����WA
��p�y6��<��>זx#�Z��p��d�l�6���)y|��2����I�.-���S6��A���PH���8�i�qmv1�N�j�[���m
wVkF�yq�Fg%�Q^��%6��3F'�eN��M�0Q����ؽ�cL�`Cˇ��xc�Y�H06���,�kw��� �*��ދ����˝Cl�؉��4������8֍l�|s)�âUa�~.�%y�ʳ�_3&"�H"E��x�cN��Y���o��ټ�Lxk-/X�DO9�5H�)MMѹ<���ty���	K6И��f��*iAÄ�ߩ��r��IA#��[:�'��i'�c�6�y�E��s�_|�}�4[!x���a�dڊ�z���3t6�MzPl��<�^�j�i�	�#���?"�q@���Ԍ�	�?MFX.�i�Vs(�����?����!иf�*���z%���5���P���<��]'�~�|w���`�"�2k#�߅�v�����}y�=�vOƀ�����)��OU�����i�oWb�&b&,�����y�JW�˴�n@��������T��JlC�G�ͺ�ߌ��K��ڕX|�Eߞ�	���$�n̅����f[��3��i�s	�b�[zU�Y�s�ǥ���|��d|]�սV��nႻ9����o1|za�/���1n��v3�~j�H?�v�^-�M5G�:���`�B��=�� �?U阹Dn��΂�>����������;�X�`ϡ���ŝ���K�|U�x#^[(�^��}ݶD��87��i�-��xK��k�r5�Pw��|#��4(-���P�N��Z��Q�ev���-��h6��;'ś�5�h�P�.Ť~c�쾋y��CdK�uu��Z��� W[��:fa	e�b�DLsM��wg�//�N���N2�ö�|kN@XO	)�k�^�&s2G(����cA�N����^�}]c6��-�����A��Rڐ�2v�sUP���xG4pW��j�����.�<UWL�Ʋe_��U���4��r^i�ڞO�$�uˌ���w��+�طG Kmxլ����2���\���29�B��L��������6�_o�v9w��u�s�r�*�Ia-���������kK�H�_�γ{��,���D{��u�?����U�9��ܲ.�D� ��R�<\R�l�	�dX_�<����q���Ҟ�����{qe��aӶW��^��v��������Zsm�ؼ�>�ϭ>����0!��À��aj����ۧMv����l#1cn)�_A����ք�Ƣ�j�v-G�0��J7�e�V���0`���m��]������l�[,�4�nwj[�ԦE�&�t�/�)̂D���*uў'!��V`z��F5�K���i����`�7�%��m�)��)�E�09���6���H��'�~��Ԥ�gHT���<>�Rmg�^�<������z���BxУxi0�0��k�	S�%�Gu6�Op�T�zr�ӵ��C���}v���1w	�~���n��OjS>����*��N~oQ��]E���e%]k	Ov�8CGE
���B���|��� ���9��Z��/n����8��Z�9/L���;bu�s�w���y�λ;�L)��~ɨ��uttٛsbղ���óng�h���JA!�Mc߹C�� MKsP��dl�`�CZ��)G������XO�ʵEVR�R)m���h�fö�vQ`K�}&�^���4Nө�Q�Я3��~�
�����޸:|H_��j+���*��|^򯾣�:j�#�f�29�� 2��K��lk�m����	�"ˇ̄�f���uo���[�����CC�4UsX<s��bcx]bYqE�EH.���%fr��v�9��� �3v��f�E3��뗘�E0~�}�q�y�yA�7������l\�7%毎��X�9Zi��^�Ѯ����0ҏ����rR�ţs�*�|H��B���}C��fɼލx0��F0=Aᖨ��@���y���W�}�����~���+�g���IĈ��.ˆ�攽����pj��f;.�j�7s0�ۦ�� �	�̩fP�iQ�Czq��\�1��g�!6�gm��Ӕ�SU*�n�:�D��yu�|�euK/�^�R*��R{���z3}oP���x�nk��+f2�Y�/V�d0-/:��"������ʎm�B�Yx��(LEP���܉�a&8�mc��,�xz�v�nq��},-�L�0Ǒn8EoW�f̒��s��r`(��O�<7.j@�~���s�_Z$f�	��.Ct��"U�.��C�ұu��"�tA�@iz`�T���,�;*0i�S�mxw�A;65�8Bn�=�	��:�z�1���,����"����qT,��z���XJ��.����]�v�}b���Х�hR�F;��*߲v%�������**�*zy�j�r��3�Uz#��XWC��di/N=��ZUd��{�6�]�&�������jdA3�'�J׿r�^��\q��Y��߿h��
?���"t�����=KVF�4)�y'Am:�*��h�c�Y&u�&���X�̰�:��On'��X�P��˱}��9�&=��K��9q�*�0mv�z�&T�����R�;�GL�3x��%�����e��7�ǴN�r�[��y�4
�#�ȇmt�L;6��gM���I�O���ϧ��l#z����ͧ��s�Y
�`l���R*��E�/�����.��o$;d��/��HA�Z��9S��1�uz��Z�o~}L[�;��tK�y,#C�q1*l��^��[C"U˧lL�n�l4Ov��76�oA!��Z�MCI}����~��g� ���2�r9��E�9c��rm~��O�4l/߫v����i���&�V%]+��p��I�(P�i`ʇ.�O�����j����_����э>���75>���m���m�������9!�"Ӯ�5��^E��ƕ㥥b�+�7э��D�t+�:��Kף#��V�J�����&�	A�U�4��pl1԰�uM5���ދ���L�ט\.���z�ɕhT_]׽E~��E���=Q҂q�M���!�Uލ
��O7S�Ji��Q��b#��s�:zkw�!�Xd�]�*a0R/��!�$K���=i�n_�Ok��'��xNH�"��H�kk�<��ȸu]@0-�JY�	�����;f�vlKv��"��I�]򯳲�A8�Ѭ]�$4eN�\F�9�:��mR�`�Z9� ����J���ʥg*�:���ɫ�
��ق�c_�t6�;gn��D/v���2�mQl4�FJ�����w�Q��w�[����I��<�f�x7!�,�f�y�N�I��Rr�7H�X��s�]�����84N�'���wR{��r!7C�m�/g���¥��c��Zv��_5@��a�B|e1w5��Q��_��b�\���N�C��Oy��Y����`a�^+�$kt������	��d��Ǳ�o��и�v�������wfOǄȝu�/�k��P����z��F��Z�p���ͪ��x��UH��f��`��C�r�a�]�%�_&oM�LNTWl*2�4[�ڋ�(��{	t����h/���ݮ��73��~�>�Yw��{�!��kk���d�S;��H�C:�pl'3L(qe]���+�Շ�>7D��
����b���=ٓ6����dLbss�n�m>���q4��^�.Ť��q �/��y�����nsV�UA����ua�4P0�Ŀ[�m�V7g�yf�����H&��W#.ϱ�;��Y-������{?!zz˲�k�J�E ���`��j�/Q��ͭe��pm�mm�k�T��z�g\�q��+��5+P\�W*�0e�=4����;6b`}u�P/��N�Z���i71�9�I��VnW�[S������Х�8;���sE�@��\�}��]��0i.m�^�&	ԙs�j:9A#�"v>Q�ʗ��|>�{����y ��j�(��O:��WX�7�_��_�H�*7n��p}7qWn�%�5��������p�7�9�>�sn!�y~�ϗa�=��Z?KT_��)?�4���m0*T3_�n�
�m,���2Ǳ�*ҧ�R�U�)��N7"��f���ؽ��|���+W?9�}�B��-zac��^��}	��tBd���s��AP�%8�ȶ�"�vZ��"ۚ�i4j��o/Xp-����}C)��h�����Re����%��q��J�aR���eE�o��Mn�]uo$^��<o� 4��-���/�K�4�=�%=�d]W�Wv�|�څlOG!,��H]�<��^=4�c��sץ�t�la�·+�D޻.ҦN�=Α܍<2���)��F���^O.������`�T�>���%�kW6L��!��6]�wP+�8�����̦�c�f��KӇ�	�4���gI�hVf0��b�Zxu
6�L� ^��̜pOB��T�)~j�i�M\����aEDI��w�e.���A/�E�v��-q��P��k��)Ң�O� z
ǚ
�ʴ�\|ՠ_5Zn:!��z�3VA�4̑�0*��,j?R�@T����&ݜ��0����>c��G�/$/W%]�Q���3��c�M���Ƽ�c��F���ethW���t
�SM����}���ZN�&��`���j���ȼ�vcu��o���o̺_Ց��V�R��_j�J���~)���,M�'��xa��S�ǈ�a <F[��3$��핪K	�/@q�nׇE�B~���<��fb�U���^��<;Ϲ��<0 V��ό�gる6?}��
UW��ߞ���NZ4�]5њD�u�Cq�m<#}���s���(>",���F����{iL�ϗ��ɱf^�짓���=�yj��u�Bȸ5�ʟBm�as��ihg��  踻���6�-��w[�c����t�.#�Ka{�����b���X[���~K�h�Ղ�Enϟ�l5D���K��5L�kQr�=�d0l[L8�yc��7��֣��	��T)=�;Asݼf]��*�Fl�ˣKs#�h��xeO��Ŵ�8���@D.��|���B���s�JS�1y��uM�E[�G�nf
4�K���̳���m�%{��Zɧ��L�E��D���ze'Q�1�څk�f���8]!ڹ��j�n��&y��.cX\�>	�ׯK�e>��_��;��񿁇*~�-'��F�v`"��'��v�M|n�9��X�IV��3��MXyŕ��]z��{-*ۦ׫�n�>GY�B�@��f��Zv�&Xo��-���m�:6_"�pզG�fY��F����yGᵾ�晜m�/7��da��t�����<��8Ԣ����.��r|�C�/�,
�=W�o��4�a��N���^�bܷU
��>�w�*z�����ؔc��.���h��,#�\9��ۜJ�Vs_h4����H�'g�sg+��	Uu��5�%C��8���9�y���2�]7ݚ�ՌC�r�ט(�8}�5t�i�\�
d��L0{yJײ���{�r(�tZ8�9uOԳ�{ͪLօŰv����(�h���.�X�f�y�6��r�����eZF�8���w�X���/�����4��gn���G@xBwml/�K�|�z�C�l#�g����4�u^Y!�8w�c�4�x����W��v�����!�Y��nac���E�`�Q�̱A�2�Wm��w� �m��!����������qh@$�1m������ճ�5���Vt�{��)C;Su/V�ov� ^Y�iނ��K(!@��`��x�?A�2�a8��齃�t�C�*� ��WR
V�ʆ��M|�\����f�rn�������1�B�y5�� ����xktL�-�+U���V��e�Ү��ܹ��SR��84�@ҵ�|o�/��R�(���"����_/j�����Bw��G(�5;p���qlݝ��+T���A5�!it��aWg��3�wZ7�n��R����WM���Y��r,9�1r])�ã�J�c�Vwj�q��p��fPb�F庑X5�|^�6��F���+2m0���M�V��2s�/�e;$�іa�'hJ��1����ק>�vN1���32�b����f�Y�WY�_B�T3Vߐ�{�ٞ�P�X6觛�V�I�GV۹����w� �N�rO�U�X��P�ٜ�噺�Z*�]�N([�^��ST[ٙh �٦oB�%Au,jU���g�Ha��{K�wg�M��p�R��Hm��mkV%k���F�1�7��]�t�W��Wc:\��[is���9���*�l�K�# �'���'c��X����='�"�3��X����Aά����L��W �,�~��8����y��8I��#�%<u�t�J0tǳ�r����>����&��f�O;k-�	k'I�6�]֫7�Qg��=��aal�C����zu��8G������E�A�� ���@�o���=jݗ �yW G�; �"��&n�e���s0ϸ�0�sl�%��E���S�.�%�U4wV��[2yv�	aj�B&t��u�E�Vg)'�>��Q���F,m��� �KZ��J�-���Ь��e�[�Q�J+Ȯ����c��[�!̫9�!��E-9��SB⑬�MWY��'u�F���M�6�qZ�m	�ܵw;�Ãt��&o��0W<�J�q�`�sn�uLp�pDQX����&�f���jB��W'�N�s�x�y�Y���f��gQ�I�1�W�\��0�y��i�4��
}:�q�z�i��{�g*���,*Gy�5�i�
�E��{�\�:$���HK��eugvR�����lil����(���kOu��U.�7�s]śL|�ݙ��.��Ǚ�c�E�lE�#��̪��ӫW6����y�L��[�DB���;i;����饎����A��,����Ph!\ֻs��n�Z�B��?7����Al2�|��u���$��H;�������6�b����:��:�Y�d�1qk]�G����:+�v��;Y[�2�-�M���R���&W��\��ɀg]1����t��ۛ9mY�֝ᓭFX�K_1�Y.`l��}�9�dt�xbeP���崳�N��K����Ŏ��r����f614��c7�*�g(��J ��i��f����+0ɥ���
���n�ʺ��˥�"w��z���c篞�|/�?9���+lP�]/�HiSHR	yd���ՠ�Ng9���~?^>>?>>>>>?_8��aѪM|��T$�,u�R�$I��Y������Ǐ�������������f
�	ԽV�����4%)CI�ѤӠqh�QF��]tz���=GQud4�IF�)
CN�K��k���%�l��C��E:M- b�U���lP:�;�κ�A��D�Z�OSF�3����RU#Ɉ
�kM&�N��N����Z׫J���֩��F���ox5GPh
{�1=M	M�Ѣ�M�6
K-�����R�)���
�(xPO��cZ��pcՔ������ՋxA�çq��\���3�����E�X<V��s6��ݢ�B��Ϫ�U_�*�I)�ާ7�ML����a�����"��>S6��Q^�<�C7�4X�(2i�^�Srs/=]a��,��ؼʺ��េ��H� D��px=��
�����jR$jOS".�{��c�N�Ȗ�{(�2��Ъ�|j�t��{w�LN5z�K�eL&
�\3-\�.z�i�E9�pKg5�ܲO�"S�H�)MLz7$v=C�hh��ʩa�y�;��oX=��2� �6V�0��N㷩RO��&*ۤQ*y�7�1@>@>h|6���\.s���`�`�C�ƽ1��E�OB�0S>�,��}���|�G4�4��]e]×�Mi��ul'�>��f�5�C��&k��Kv�*^�+�(,����R�e�?X�z6_aA������eA�^,�YR�O�W�9.옧�	q<�S�)��z����c�!�����y�i�;���¹�yUH����`�C�y���ץ��-v�؜{G�m����=������Ʋǰ9t���nl����ۮ���M�Ϡ{�
bX�'��?�i̙���fb�=�F�[��:W鶙���	��]e�u��f����vKX�Z�� U$�����Q�5�B-ֻ}��1aG���2%Z����.������/�g2�B����@���1n��3N��w����/�����\�1,��hl8ٯ�l|�E鱷})86�L(rh�Ozmڋ�9j�/a�G<3ޑQ��;>#�{}w�c��� ���"��v�K�� �B��N���n�=�o��/>q����P��3���SD/aB���CA��`�؝wG�^Y�5�(�RRj�����4����F�\/%�u���^��������	�"�Y�W��_71`U�/ޣ[w����n����_�����yC���*�C&�s��<'�}�`�����P��#~�O�J�hy����\�0mmT�lj~k;'�,�,h%լ���e�T9����(>�\J8�ޞ���Bl�Jy�{vu��FGs׺ �M�k�	�0��%s�8T��ǂtV�����~t����97�o�&���尤uLf�H��E�&�ވL��xNx�A:��S�[x�c�2J�,�ي�-\�zC[W��'�, �U��f!��"G�ʤ�Ʋb�1�I��Fu!%�
���9�ȪݨM�A�+��ᅌ�d�Y�'$L�}Y_p{#����=���L���H|���E��-㕧͡Jpy�d˾\�N���+e�MYʖU)ўz7+w�;'Ç9H��2-��Vnn(d��/ph��p�;9Ҡ���r"�4R1��y�wU��b��Je�BN�����-��������(��¾�~S��Ź���O6[�.,{��ک�i�}��54� �c�peς]7H�4(����6�m�4����.�1�3����7(�����e��3����`�i���p�y�s",I��\�P��{�ƪ��#l�q|T��5���`�{mi� c�Ccjܫ�&�V�	�J�jT0N6)�	���z�jǃ�8≮aK_
�/l�����`�_6�r��DV�,6�Y�Mj�fX��&���aٲ�VW0-Y�P7�t����HV�J�=�U�ӗJ�Me�pV״6P�t-�3�!����h��#-���{�v̽TX�ArN))�D��Y�Ы�n�h�[�"|��U�-��,a���'���ݦa��{�����f_d�F�#�sBFG��C���ۯ��^��h@��1��I�掄�ۏO�vq�p�F�7<�3�1nYQ�7��9�=�>�w���B�5��t�L\<��>�s�:��0czqj�׾-�Yp�V�sؚ�*�a����B�:�2+2���뇠3V
Q[����r��	�U�˂\'�r"_"�0�/��Mу�4�D�KC�y�)nH��e=�hd���:�!B5�p���t��t���k���9b4^vV��E�n�D��U�T�5s�����K1�s|A�O��r�����
���{}�u��͚g��{����:r5풌�c�#��M�)	��"S�ܑɭBy�g��Vc�OD>B�t-�����C`�э8�Z� "%ux�>��Qb�!6�Q)�\�8Չ�V���6A�}~T��E/F�Ob�Ӏ�p�.�X����9~���7ƽ0r��T(J窨�5��9؍>xm�Hs�5�&�خqA����q�3l�c�^�!�6��k��Ĕ�%�w�����1�λ�yN�o*�]ycغ�-�b�������P�2XV��7�֠��Ι�t6�a �!�hR�1W;���U���-9k�M�j���A8��v�y����ެ��5Fa��<�,6�LZ���Ȏi�<s��a�C9e%I�V��+�P�zY�um)l��Ӣ/�t�Bg�)`c�:��xmX'hS'�a��R��%�_1���ؗ־�K����!ڟ�@]Գ1lH��`��~/0�ٛ-�:)�˄¡ѡ�i�˗۵n�EΑu~Hϧ�rq 3�f��A��F�f���h!�wnlN��w��}�9�-=�(�_b����L��m�*���ۦW/���Q�\;�c4���Q�}�1w��j�K��%��b���
6j-��ohJ�a9��:�Χ^Kʖ	s�n�p�R^��*��6�:fI(�#9���Փ�F�)^����C����M�Zh����4�>�R�܃�����3��@ܮ�Oh�nj�C�kü|�@�踨WKj��͊+�ڕ�s>}W�A�+z��5�|8�I��>�n�鋇5�,�Xi�1GM�By�C ,lc;��%�ލ�ע������%���PB�Iwy��ku2��9vf��:��Ó��<��}hj���Ә��s轌�8��n;1�T��mޭb�
��El���8�@	��=G�ώ��2nQ�.��E�EǦ�J�X`eEzB�%6�u�L�K��l�m0�#�`kd0�z�,�z*W�,�=Ve��@��YyI��I��lOp���li�����/�t�'Q���Ƚ���+�B�G[�sS:|��xOٯ7��J��|ucq1��T×�D�{=���~1�ߊ��S	Mmb7$Od\:����)��ɶǭ��g��h�9�����ρ�L3�����e'.鸠�7�T�n&,�L���|<.���+D��og/:|�B�}Z�L�Y�&ޯ��H��d��(���0L$s7����%���q3�6��e[c��\+(u��5���0�v�T]�SA��'��"���/U0=XbMA�z���Fv_J,^*�쬨p��Ybr�W��c�eMT�Z�۲������[6�=[a(�ܤ�<��䮟Q��'�i7b�W�������ʫ�$S�fK�4�u@~��-�kL9!ߙkН���"z̮xE�m��^vsy`�Zἄ�ˮP��c�,��wёl�"�h�\���@�u[�em?%��M�6U���z�+jA)��k��̀�}����w���
gvmf>!����;1t^	#Y�0`�YoQ��0��r�4/m�K�I��T��=&#ϖڨ�����Af����-��<��V62��E�]��ox
I��P��_&�{K�6�_��P�0����~Vm`����X��@���}�0��C
�ʕ=�I�r#B�:*/�yڙ�Ӽ���;)�_���ol�0#_�i�q�"&z�֜�ǵ�_X��%�Q�|��0��}���b�8�7��ol�Ʈ|�o�C3�<&P�aql��xU�z�ٳ���%�*�o�B~�~�]!��CspChH�l��S,����x�؇�zaf֭5�36҇�;�\�RKʢ��wBO�~;4����]4��5h�~�@g����X)n}%��P���ķ!��/�ӄ���ʟE���{]��s�h#w��,��߶tZ0w�0,X���3�&W�-��	g� �bZ�C@mV7���z��[���MPi�ۮ�Cv��pf�i�T�o\ɷN�#Ci�T��}�j@X��t	㾼j�����Sl��|*�<+���]���D��e���vw��k8�f&�ӽXş\��D ��BeiH�
u��=����2�_$�ư̂�W{�����y�{�ld�R��`���}}%���$�c}4�न *�����)�q̰U��i�.04��;��!�Añ�¶Y�4�ޑ>ޕ@&X�LVb`� Τ���vT�j��[��hP�a�p���H́ �#}��	�G<��ʅ���&x���S8�=U��s�X΍:�1M��7@M8��m��p��}"q��؆��.��r��<�Yξ��}su
9�i���\��kr�|��F��gw��t4P��t?[�[��A������6����h[Qxh/jw�;'_%�-�c)]h��\Y�xhP��Ӱ��"�kʽ���PP�L��� 㢛����z�еa̜qD��{*	{e/�^m;�s��4�4�>[���{|���)���V��Я�K��x��ó+�VW0M���C.�ǾP'(�1�*n��s�[[F�52�3^��3�C3����0�y�2߯��<�C�^�,:)k���J�#D;�����Am,�x�\�q&��'pZӀ���fxJ�|B5�}#����곾�]O��9�x��p���Q�8W	��u����L[�NR �7�k�@_�k6�ׯ&��kd�7| ���E:��^=}9��K����O�n������}��֞���j^�;.ӯC�����c^����?Wʎ�>$/��e(�~�W���&�E����'y3n-�}�ܕ�Q�8�*���y���V��P�9�v���2�f8�7�+:��]A��xWaN��R�NE����֛�(<�_A/^J�!^Dך�%�g��T�S�<�8Ԯ�+�֘��yç�{B���b�h�K�B�{R���!s�;2�,�o1���6-�EE��q�������R�Yi�g�[E���A{��d�N԰�<�%6p*E��,T):\Y�z9�����"b�o-~�ӯ0���aU3_��Ɛ����P]~>#
���BfqY`����-��h��N%��w=��y�j�U}��֦t��{w�-�"2`$�=| ����wνM�j_�t�fs��x�@�u�{�L�1E��!�eJ{��
�DA`��и����X�O�7/���^�b�܀�6E���EL9L)0A�-��#��ܵp���M�8�.�l�"��J|���%3��z`cnz�zŦ���wEOC�����PX׵Iw�'ڳ�)W����?m'����L�b񽵩e���2u�ha�<�KS�c:��k�Y��z�=Fuk&H@�y��b�P�^��Ak�Йr9[���[&��W9��-���(�h���جִpW�6��B��H�',��^��bW&+a��>��y��ox���,�d�������}k�P��a�^�YB�Reվ7J�T$jOzN6��w蚑 yo���"�x�8F�2ã�:��xlY;B�TwU���+^	s�_���z:.v�Ej˩�]u���R]�펌`�|�C�q�1�����wc�7����w=�<�Gn9L�f�;!=���3����c�NܳO��;M6��_R��h�Ϗ�����l9MN����'��/d;l��y?t;�ks�S��c�J$]V�O�8T�Q]�m�闕�N�~�� "rQxlnW�;:��4��$=q>yI�l�}�>u�Dx��-��j��-	�W˲�XΆЬ)���kr}��Y{�����3N�^dae9Aw�
��^���{�gk��a����P�U0U�k*�^�X���\��y�ױ�y)f�rn�������o��d�	e᝻A�/i�Ũc�:�t�w��ڼ,:.���L	ܨ�=��-�ԕ�Kެ�h���i�g��j$� �����[ռ��f��,.D@<���SZ�d���g3yP�xԠ�x�� �=�#4.�2���] %���GG�)�,��TS��g&X�6������Q7Κ�!�xRy�QfW�9�����B99�΍�j;�U�cPF�}�� ��H�w��I�^"b���Rε���t��K+yj��B<�o7���Ѳz*��)���rߛ}�)�����+
�
�o�C����=�ă�]؈����M�u
�۳Z�L2oD��q+�P�UL���O�
�Li#I��<7$O�d\:z4f6��Sb�K��-ٸ�F��/! ��Ft�O��e V�0W���7��O�!1W��5�J�a͝�/Aa*����L�ȋZ��\"-�K��<�l#��D&����7�$�|��m�,��(�����$�[��+�lbLr�\�y�a#����[~Z���~ҳ����D������ef"_�'x0�F^�#[��y(�t��0�;�d[ �10m�O�sס�y��ȞuX�13e��s��Ӧ�ub�r�����k��ͅs�
�FW�-ݚ1�3���C�9�3=��R�۶�i�l����-j�P�-̖@�k,{�.�Q���ϖ�Їm����s
��h���-�Y5a^���ngbܟD�ɾ�Yғ�,0�����ͥ��xԆС�@U:���P�a�/K�<h������~oC�w������F�]�q�nc_U��~�<�z���JJ�B�.Z�`�����#����F&+�Gk9r�cj����\&���M�]O��aE :N�	vNf� #q9k+����s�M���t ���v}Հf|�E7��%���l�Ԯ�˳�)j�7��2s��p���!�{�\�$�V��zvn+ǎ�s��W\���4�57ы�5k���)�_6)�7p�fJ��+�s2ܠ�a����K7�*�2.X���m���fJ�Pa�#߁.�� ;R���*(�G�]���J�>ɿ4x
�9�pU��A�]�	j��-N��Z���*YVk���x�-��a�UFXL���V�8�o�䮗e�9ve�iOS�n��Ỵ�R]w�U�*9]��� *���'7VXv��)hT�a܈����A>��;�횁�4:f�\��|s���s���l%oV���U S--��A�M��B�5��&'x��rv��0T���1g��u��*�'�sy�xl\�ǻ���4�ǥ_n�]m��N ꢷu
�YL�2p�N�}�况�:�`�V$q���V;��G�KY�^��%�$Ƥ�h�Q؇�I��B��f���ֵ�D���*<+����x�Nֹ"�����H�R�]��@�5��t�Ӌ3$J��fv�5cD3FiL����t �lc�D���䅪��nJ����'���0r��:rk��[t���̧���1i�a��ˋ��d���c��v��i��8�3$I�p�"s��I[�V��Z,��	"5���Cʫ�*��Ч�Oh�]���ʎT�1���3����'�>;/�t�f@��'K�<\��j���m���&��9k6nuM�6$ʹAo��ͫ��8��s��6^��k��h�b�*��N��HU�7������h,�R���.K ��	Q���3**fH�m�՝=zU��!A�U��gn���������ԝ��<B�
'oC)j�����d���u��Ǧc�ѻ��oJ�h�e 0��SmǊm�7$�����i$��<\������������Ѱ�]A��;����u�1S�h���ޞ�.LW�X������C[7l-[N��f�Z��*�m2)�$��3��6�6�Z.�ӻqBQ�`�8��[���ow(:@u80$�=;�ՙ$�=�;b;;| ��%|�qB�#Sm9�[�Oi��Ǻܺ�����X�ʗXGI�_f�����8�q|;��:��к5�Q�d���Ԥ��x;b�aʗ�̱���1�7j>�8H���9Ns4�9S���\�=շ@"F�g�q��Os�I@r������/[������W�����	c�,�,������l<��r��]V�A�(%qm=J�e
n蔴3u!�D\�1T��'�v��hFL�E`��U�][�8C�8�-w�6��Z����aN�cu%�$oO�4i�K���U)�ti )�DB
TCi
MGmʢ^i!���D-
W�1URw��,TTCI���h�u���ϏO���������������x�c�5��y�ui�]g�w�$�Q�i���s9����x������������x}��i&�j�I��$;��4Qԝua�cm,AI��:�]tP�bu�ӭ�h���޻��M%L$Iu�RT�Q�و�������Jj�)�m�ڴh���:���E�JRPD4�cZJoV�Βb��i�%ֆ��IV,3%Dv��4�l=�6��T�t���ѝ��ݢ��5��-uMm���:�JS���h��DE�U��Dui(��LM:�"�Z�$�GV�����(h������j��*�AVF�����ƻ�c�:��nw;�V���Y'�-�>>Ňo�)��jL�w�^R��ԓ�&=�%s�:Νq��ɠ(�vE*v@�����7f���ǑA�C��`�;����k�h���*����т��۫�S��n�pDy��o�~��f���uV�_W{���]qPߞ�� �FER�!�-�{ʷ�]d�v5��#]�Fݼ�ʙ-�!�vA�A,��ԑ�בO�\����x�`Xd�P��yS�4��o�(Uol".�ʊ�<�>���YX�]Z�F;H���467d�Y��]M�}x��М��?�1��c��� �X��*��R�T�_0�=���I['v�dսmb؇���p�Y�ky9�v&v��ºkk�`u�)�JB�U�����C���Xz�&�T�����ht�MƏ'�;��e����:'̀oR��٣l���g�C��i��Ek�4)�+�����	̀��b#�k��']!���{!Zk��N���0���c9��X��&�\�6�Ms�װ��G��2�e-��֦������7-�B��oUn��X�s��,kB`jJxw������A���1]��M�BR]���.��޿>WW
�y���h�K������B�5ݳt�e�lX�zvdq��%:��M۽*ܸ�@��)
�4+{�|�Oi��.���( �.�EA31^�ǚW�\Y�3���̤��"�����C'���x7��� rҊ�t��m��@�I�^[��SƁ�vN8��*�
�y�ڷ���O�]/�K���w��^�xC^�鰳t��?2�&�ޙ�9��(���eA/l����8��[G�,�y�![SS���g#c�D���ʤVW0MC9*�.��F�v�f޻Zd��Dr��܄��Rū�`az�{�L�g�`>�L+���s�<���qͶ�u�Lڦsל����L�D��Q���z&dH:"��)П|^]�X0 p|�v���TH�є�[NC�k:��im�;��a�-�sd.�4qpCp9����-��^��6 `J����!���cj�����m%��d"��X�ۏ���-W�K�J�!A^i���t��:RN�K-x��fW���?@T��AYC��r'�5z��Kc.P��R̠hy):��9��e�ʺg�؜�ͣ�����1P����k�g`���1�0X+nXW	�yHL��ހ���)�3��ٽ����۩;�(�f=��Ot��;@ Ųaw	W�i�y�����[T��&��ĝQ�@餭e�u�3;��sKC���I9����GE�{��A�S1��r;����ctw*���ի����Þ�؊�@��G2�3���:���$���ӏ.q�`��:��Y�!�����R�9�W�I��GZ�߽���{������.s�c��,}�b6s������{���2%�tTn܋���E�$Wlh��֗��A	nW�wL��Ĳ/atS �I��~�X�'Ң�p���̀�@�ɛ#���]�ǕjX^��6^�/�;Ϸ���ʥY��41u.i�hw�7ݖ�us):ǎE�I��Z�0NDk��7�B��������='�%��R]���f��bn2�
ێ�S)0�a��-�*X!<��69�5�ܧ����2��kUR�x�uu��:�6y�x]��Izp�7 <#Xt��G�2�����S�)����N��?Ï����gvJS����yI�^��A��l��e掮���������C�e�<;6&X�&b����E���ֱB0��c�Q��}:�_�N�z����ۧ`38���h!�{���E
Ȩ�o��յ�	v/�/d;d�{?�=~���
�s
�%w)��J�	X��*Z��;�8ɉU�Kœ��@�
��㢋�K�%C6��t�l�C׸�$�K��,.��͸�Tݩ�������[�c�e��Pm�����K�0*p�y�%��b�>YJ3ﳆq>4��ѼK�����ȴOJTtX��F��'��Q����>�u��V�\�)�n1�e��W.����-�Nc`~���cS������y�o0��m^����GQ�{��������4�RAd�Ľ�ѿvׯ/��szK@%��v�U�$��':��,x^Vj�p�"������,BibǙ��9�&���B�1�%,��l��wC4=���q�â�^hh�t7+���r;A�f�'�{gS�)�,8���������S6�(�2�y�P��XP����\�n� ����2�&�j$�%ӌ+ǣ1������P.lD��<�23�1@�Kh�"x:��{Xmd�sWD�W(�E�%4��^
:��=���S۹17����UQUm�&�E��bS�u�>�a���
���N�yGI����^H�kk�nH�#����D"�zq���yl�[��qR�7!�~��],�M�q#z�$�b~n�Gg3b��Q
�Df����U���e�1z���j�IW�� �M��0^Ȓ����({���o������Vov��H�YOZ�)�0�H�==�qQ��0�a�mgb9����ֽz����[�Y`�f�[�e�B�s��<�Lo<!�!1�����'q�<Cû?�-���u��y�MĦ���˼|��n�z��٘R1��s��k\ٴ��i!st���C�c[	��d����,u�Kʻi�H*7A�$��M�P�Ý*®�'T��T�+A3]�7�gJH.رٝĲ��o��	:��&�ƟZ�Wf"���۾˰;C	�7����c�V�jk/�dSf��jނ�!k��ͅs�򪑔6-ݛ�I��;�J��b����N�eI����z��z����"��2Xu�e�c�O��kg>XH��.L᧪�0Цi���p��Ab���ς]���ChgJN
n�a��5���W4&�ؘ~a~ ���ޮ�v�3��2���`�B�p��;E��+~�&d���#;
�1%��Y�23S���6e=��xn�hdll8��-={g26D����F���Ǿςpg�֯�G~�7��+����!�wf����v�� ܺ�[R~�m��k	�"�G���������&�;v��Y�tN4��Hdzjb7�Hca9��/&�W@�t��N��j#�%5]qP�/��{̀�wi�dS��Y1RJ[]�6���~s�­3�p�'��Z3~�4��P�(�B:�D`�O�-�b��+䌞�0uR����N��D>V�%&!�.�%Țg1s��HG�xEj��)+�֚g�~����WE���d�u����a�(���w+g^v[�*�V�&�� �k
����z�\9��N���^��Js"�%w(��w5��
�{��gzP�N(ݱ{��([;�P�u��[n݉:��j�[d���y��oxB+wl�	��g�>��=ŰU���nH��D\�!V�[�7�b �����2������d��A�
�66ƻ�;����K��v�αQ�� i��v~�RQ�hrV�\HmK6���3��@���;�������
c�D�=��ޜ��,xQy���Wt��Iڼ;3��b�S��^c3��d�XbQ�GM�R#��g���r�k��*ݟh9ßE袱�.i`��$�To5�0t��p��~ł�Ҡ�ܞՔ8�R걏z���Z�2��#�A����;�<�ƨx�*�VJ�H�[LFr����Ԝƫ��ӄ�\��6}ذѰ��Z0#�/�%��!E��d6{u��n�W�;���,s@�;W����v@�2�k��D����`�K��Jy�(T���KF���p�$���:*5��@��C�"%��=�V%55T3�C��y�k~�Kpu�ƺ�4$B�K�����	��ټ�B����S��g��[����w�0*�QX����B�_^
w�d���4�������:�� v�p���a���BY�&6s^�f��m����님��͐�����o{�t�ϥ���^��՝b6���m�"&�Ϲ#Nri��%�DQL���=���r1N�/K�ر��ɡ5�s娮�AHWdL�����~鯲��G5!��~�X��Z����0���FD�*�h����q=��LS�+��=Pz����sSNdU��pM˒ .�
�Ƕ`�h�պ�D__�p��6Gt�O_�)Q����D��gX#4�*����om?\��"�V��G��M-���=�_�����Шv��qh!�'X�4�j�j�0��j=0Ox��N�@a��˚��7uFK�j�f�Onv3���y9��mf;���貚=EkΚ:��t��r�	nۊ��{�UFc� yLbm���Ə7��S�w_+�J1��nc��j�k����ٴ������0ހ�oLl�~��wW�(z�yG��=d��qİ�/����R,���� ����`�;/$B�zWQ�/2G�ü>%LI���S}�7P"�Q�?%��dN���i�_Jo#�"���ؖ2��u3t��&mlUܕI�yଟz��=�ӌ�o,�-�u7�d�/�;����x|k/4;��~om Q5������\mW��pG��w��v�R,�p�Q�i����3�(>��n�u�NQ<vE��표�4s^㊤֭�W#�v�)�m�]��zD��O�z�P/�>�k�����#�D��	��;���Z�p	��-`:��5XhĤE�_�W8�=�!%1�p�:r�yq���(������_~��P�Y���I,��47U���H�M۴�һdՆ���y��e��꘧R0	g���'T�D���]��إ�]�'76u�afl����A#�#6�.�@,�P7cc����gZ(Kk1wl�n��+d��#���%ঔt����d�ә �Ĵ��iq�P������
V����P+��]���A%*�t�۹�n���*a�m;4BW�״����p�)�-��_8=�]#@�oP��_~�]����W��(�¬��*5̂]
����Qe��P�)�qN~��]l���r��>Si:P�}�']O/&�����|6ߡ��+܌(j#P+%{���d�dmh���qt�֞���TJ��ԫV���8p���kn
Y�����w~��hP���q��C��g��4y �`?�lUbJ�����'�q����̗+��(��ţ��R�θ����f�Ρ�{8q���v�|�x���m׎�CE�P���:=}
Ev�GZ;[��UUm�rA�Fa��~e��Z��zg:���,���������������~svx��Ȯ:��f��I_�x	�>[\��p�{��i��pӖ_{j���A��Ty��7��Kt�P��@�c;k0�&�p��j>|,wgE���+g�y�k@�4���x���$��졝dՙ�0����5yo����R����/��	�ei̾K��)�ɻ��aH\��]��龙Uw�!����9�꺣�U���w����:�}=�ز!`I�^���):$ߺ��C:��	K�"�����g��c�]�f^N��;f'��%14�@��t[���Q���=����H���G8	�i���Tx�^�qV�ڻʃF(S<(*��-�O"��]��t�-�hV�m`t6����W4��˪]kk�׀5�u[�CTW�;y=,���U��K��tЅ'F[ժM�-
�tV��4����^�W��R̜��/��j�� 7��y�n��75R�M *��f�s�Jτ�®U�S��6�v��e�1�2�I��6U{&*Gr[�A4���dz��c��0}�;	8�s��h�η�i����߄,�j1t���u�#Bɒ1�ϭw͙Yt��b�o����H٧�4�B���+xEj�b��ڔKE]��0WKngJ:W���R�7�N�vd	� ��)���
�J��n��pؗ;����G:EXn�%q�6����� FW�.�M��1�1&�p�f7Qy��ccj��낳ڥq�b��==!�8a1"�f�u�D�jh0�f��k�Ы�A�o@�3�/���K��R5�x��?�T���p62�E�jd��v����C�a�u�h)��3�^��U��ʽk��*�N��'kV�z��Be��;�P�ý���h��yɹ��Y#ϛݘGj��ʼ۬f٤�<�p�J^�Kh�K�NN��j�k�7qIjf�sEQ���+�0*,�s�m�@�Q��2��4�9mi��7�tp,�X=�Ldn��Vs�.��73I����l�jJ���#}W�d+í����ۻO�.M�ט��9 %����F6K>��r�Lʓ4��`�����QK�8����r��uJpQ��V7o��;%h
��Y6F��;8j:�Ý�s�dWX,�X�
�rc^��ގsQ�@Xd�'}>�*챻¹��˪�{e�.��98��5���cLWX��P�Q�y%�C���9	�*�R�FO�˺`Ǒ�k�n`���3�cю�0�v2�2J�5��a�[�x�W(�0VV�d;���9bN��Ck�cE�ڃ�چn�|�f=�Z�9��l��b���͵3^��]�l���tV��w�t�#�)����(��--�1�Sn�aȷ�"W��׵�־+�pK���hh�Wt+MԮɚ/$ۑ�l6�w^n�vt� ��
|�s�,�]O3�ۡ�yV���D�a�m|�1	��wq��/���� E �7⍾����@nhm��p�U5��
������F�����mP�qX'Q��ru�0UҗDC�{>��AOK�7|M�]�MQv���"�r���z��j�<�<�|�<P
t7.	��N�R�5�y �Ռ��BF�)�l��onՋ.Jd4�*�U�� �>����wrTI���Oz��8x�v�=��n�����\T�]ź_]/'e�����yR�P��K���:�.^ΐDF�{ٕ��R�uqͫ��h�{P����W�*P��J�O{*�L�q^�<�3J�}8�]q���K)�N�-L�?�PЯ_��}�1}S�z�A��t��qV��ߣ�sh#���CU+�n�2ff�p̬3#�YEI0U]8O*7X��Ri=�s�{�ڠ-��>��%�щ��pH�l���Bݭ��m�;)�-f���"��sD�k����8Ӗ���Ւ�C�'.�U�x9Бe)L:��c�Wl2�|��/U���t�H 	P����vv��w����o(���	ǳ���u3XŤKӓe�E)!�f�LI�d�Ɲ����۹��"z�����Gg0�(�x3�Pԁ�5Шȅή�E���m'iP��ܗ�0Ȯs���� y�ӱ�%\��#m���=ٯvrqҫ�0쥦�����G��:Y�*��خ=�@d�|��jƥ)]�:�Գ(���{Z�`A�х�9��1��G9�Q�XVV98�f��Uhʝ+u֐�)���JJe��s��V��Ԓ�A�EU�]������ԖᷱT1)ʚ��n9-K�OFN�k�,c�ֶ���6'JBZ]|�r��-ǽ,޽ �;B(�� я(��M=��� ���n��|���Ѡ��l�EF������
	����c�3��oo������������Ñ�)"to�]=BDkCE%�����j"&���Ѡ���z�����������������������y��}�UC�RܴUD�ƛ�THh����S�)f�tPUTD��P�u�SgUN�5EDKQU�)M���"��j(�؂�����"�*
��-�ITDVا�&:��EPMET�MS{��8���f�j����Nb�+��&�����F�f���R�1DAUDUHI4kEE��QETAMRL��DIG[E155;mj)���)�"�h�5�b��5]lDT�Q�h�:R���������զ�cQMUM4Uu"b�`�d��f&�����AQu�
��*�b.��4UATkAE'��Q@(xU
(
��kZ�.���.y��f oz����"����3SY�$�p�����qU��tHw$�#��{X�T��]z�=} �o7�~2'�,�%oݵ'�рv���^�G4 ��z&F*p�5I��獕���pw5R�ۍ͞���Ę���V{�ぢop-�x��K�����;r�C�<�^�Y͑[ˉ��ov����h���'���ыp+p���og6)��W��km���	�H�ǘ����V3*SGOw5��;��be�ދ��Z�ѷ��7v �DD�FH�{���vM̎�2�����z�QO�����P�a��עc��.V�� �.���tc�X?uA��{�j���1�^Z��u�ԅPF��+q*�dM�1���"·�޽�g7�~���yzҕ@B�v��UC�l���n|�U�-j�wW+O=A�.	ml���#T.�R�@T�w��� S8��RF:�3�6]f��P��E$�z�h�ҧzRE���Ӳ\����N�y7��qsw��]~T�ɃF�)�@�ڗ{aI��� ��I�Č�OT]��4��wn1Ee�e��|78�z A�v-����='�R�씎32��q���J�w��wzK������m]k*tQ,��GZ]ï6��(����-h �x���4]vl��/7�x>�_p0�M�/@���ugP�
���)%�c��Y�Eg����ş��7��;N�
3(j��}��������O�V��I�O�V��4u6��Ѯ�5-����Z�O����8mR�'[m�t��w)�g,�L���mW�q��ov����ؐN��i�t��L�`S�>��7)�ͽ��q�j�\���ۜ^��qY�P��d7�r���|�k�8�3�O;������3���::�?�! ��pX�~Z;f�9^'���Co8t�h�\_�w�S��(�*{g��S����~G����|&�o�ʮA[{t��i=Qw�ڎ�c�qA�;>Q�5��{Ko"��;���F�-q9��SO?@���W����?��>�@}^��Yri��]tF�KZ变O�+�v���Ķ
�S�Ng�,�:  �5W陸�Ȑ�o~(9ي�w~1���jQ�����9�6�]�oPR�>�,?;�FR�X�xg��92�j=��]�Z��E�8%�ܬ�4��2΂�N:�]�Jv�J�_GOfM�O5�}#ʹ.٫��)�qS�r�P���\��S�z]]��ݔ� P#�����������eܑ-��$;�WƳ���M�Ii��]2���׬#~o:O�,�_C�Sj��#�U!���.c,z��W��pUj���z<}��oYQ�7!�;�������Z.Z���<�)�͑��\���]��.�^:������l�s;��T���M���p���5�5�x=C���(�ָ�!���g�S��F��{*�@Ąy��<�NR/y�oJJ�G>L�ǈ�T�Ì���ڶG�{�����,Bَ�
�W{r2�^:y��ph�is٬C��0q��[��8���I,c�-�B����]$t43lA���Tׅ�Ui�a��{�\u�H�%�+��gme�[�n+�L�b�޳��V�{�̇w�\��K�uƪ�u^�*in�2�
��ae�	qӊ���{|d�+qܦ3ۓ��K\�$�}Y˺x�l��T���Z�wn0�ڠ��A�A�ִM�Mͼ�e#Z��\wT�ք�%c��ѫ��D��Q�8P�;��%�j���ec)}¨*��(R��=��vVP�Z�&EC��$��w������*c�es�x�]���lajx�j�C�������=��9����'$�oj�ِfC��yy�<݈���o�\m��i�I�ing6���V7k<V>7�_����8�Y���U����*�Zq1K���wg�;��፞-�G�t9��0C: n�l�	�Y��q���k�P�ߺ#0��yf3{<�y�$#����=f`_�!d��5�*&3��k�l��.�D�����$7v�W˄
�Z���LJ���&ﮥRnl�1�.(n5T+6z�L\��m�4qI���g-�d��@�����Dшxd\���g:��ߡe�^�]#��t9"s�N��m��ו�l� ���/�Dע[4�6}^�Q�����iU�2>�\X5{߰��c���O�$�zH|��GЎgH�ą��sT��so��7h���@�r��t
4x��J�-���s9�#�u/S��O,N�Fo��k-���+Oe�G���<&<���;�I��0�	�Pv�;GI��sm�ױc�er0Sx��h�1g���И���޽����֕�֥����0v�*ʧ����U��$��l���BQ�j�{��y������`?DJX�LW�A�I�M�O��\m�t���Xup�6�]���e�f{�V�v��|`)�&C��&���J���T���a�Q�1��Get��^S>���;!�ި^�S��l�N�ʅ��g{i�64&[9�k���noZ[� �m��8f�a��	��B�zLM*��QUzE?�:���.w�L�8޾>8M+U�v�Ͳ:��o�G3��~iV+���$4S�e˷Om��j4˦�j��;�a�F��z�~�w���{�t�߿$�ra�<`vU��a�L�ݒ	����6�z�vr'S�������J��^ >?�)y�ռC�xf��w�ǚ :)J	Dh==[y���0�'�D<���ϣb1礦6��o����/�#$=VUs��8��s���I�el�b��8��<BP�rk�1�+.���dc7�b�&Z�2��hE�����츺��K�7�c��N�-f�M��s���ÿ�������4/ ���M,��ŏ�m��Y�t{l��^��v�L�m�8��-[�kGh7��c�웻�jw	W��y�oT�=�]�]��o���/7��0t�n�e�"�w�+��kf��sNz���-��m.�.W�&�aa���ۚN�v_��T�*��u������ȫd�e�r�3�ɍ��t�_Kh�݌-������d�P�zɂ�"�����:��M3�
� ؙ�-zؖ�:!��}��B=[�F����il�+���m�cE���w��C�#��s�q�C�]^�:=\
�ћ<���)E_���ZhMd��\�;n�j�oj����D��lx59;pY"5l���R�ȵ:�g�U���Y8{_a�H��%>4��S�ͼ��Ӱr�;���:T�P�'{��λ>w�h�<�N������7=�?G�-�L�f���c�[S%��*W�6r_v�{��(��T�3rR}�7��M����˼���6*K�)�]�Y�h?-�݊�h*r�= ���u�P'B�=��Ǚ�GC)��,��G�vJgcp�l�t��$@[׻�}}h�5ƛǂ;�&;�i
�iV��c�����5�{G�]3���S=a�^��2n�.�6�Hv�Ә�]|�W��J�ͤ��Զu���Z�n����՛����r����ox�Ϸ� E8j� x�4�D�����o7�r�D�������%�0o�@W��O�Q��͗����9�H=3ۚ;��T�d5�����³N��62�N6G���O�q!��s3嗌8�[U���jǾԁ�*?�"/�cߐw�]�$�`W��S�T3N���Ѻ�ȍ�=�@;���B@�Z*�N�9�KŎ��U#&D�����j�ޖ��cغP]�8rBGZ �F�:٢�,L�Eo�v��{Om/X6/�`�^Jdl�*����׹ ��t�v��fP4��&�+�'���:��P챐��'���d�ʑ��T!t�|�������%\����f\~�����~To���^��'
<؏3��;]�fx�|�޼���}��H�2�n:���p �H@~
��"��Z��H���t�[\�w����x��=<uq4u�=��A�9]x�C�U���plx��z�~ȹum��l�]Z��	+��td�J��{u�iܬ⎟l��#����V�������z#;ף~�ՈN����]x�>_v���3;)�W���w#۷��-ךs�\��o	]�;y�������o0�������bѪt��c��Ə
ߏyM��4�zζHeH�n��-8�����pXD�Tw��7"P
 ��3g��B�?-y񴌥�˱�2�k�Y��D�Z��c��Xg!��~Α�Dj����J��S
�'���a�� .�M�EA-yL_�>�&}b��v+&�5���.�}9��u_�����5��Gd�9THec���P݈��+N�s�3��3K�o]9wY��s��7z���v���힐��C>�g��u]Qڒ��4S�&nl���.&rIny��4q5�;�g٭ˉ|:(�S�C: �y���H���]X3���6�Eڀ/,��{� O��Lѯj��heՌ�ߐ�ssQ#Diw`;�?�lPă݁�b\VVݯOa�U�GJVD��\��O@��;��e����3�ܡRσ�P��Q�"l����f��	�4�l�Pf�s���`�ێ��}�G����7ك�\��� �����4� ��W��V���H����+������`z*��_���=��Z{w����E��#�0w�&Ѝ�R��AY��Ύ�j<�7�͋rV;̮&��7Q�W��5�ۻ�{�7��و���"Zr��������X��-��bTO[�d��J���&����N�j��'��O4��B�s�HEoyn�^��ϵ;PI�}��{�̯�x�#^I)Y�Ǽ��<v�wc��̑k��ɨ��3ߨ�����*F���u���<��d�M�d��>֋�67+cu��v^^#��sg*{�j�,i~9>��A�-;/V�\q�)�Ͳ{������*�B���fzޱ��(#��^&#���z��UB��R�h��xӍ�4'��c��w���d��x�`r�ޯD"8�X�7���J��-a��1�+��o8�g��v���^M ���`�lͦ�
��"��%���s�	F���I��<sr�	�`*�6����������&�Ӂ�_�u���5>f�<v����hgk��M֧�~���R��� ��7Ƴ��&P���V0� ����+�Cͬݲ��=�xҹI*��wp�����'D|/�b/��LήIQA=�w�r:e�+tP�)!i�e����ӝ�N��,#i�cv�������tp�g%� Î��Ο�uӥ΃��8�nU�3�umx/7��N�ͳ2�Ŕ-�MX^�Lh'�u�&#݂�@�nq�y��)x�y��]U�+�8ǃ��y�w4��>�Ǎ�D�I�<��l�=s�],U�O�
���i��A`=%>���֏{՚�ϯ|�C�װ�� ���^��2�}v�(wG�J�MD�H���]L���g���oM7D�fj�C��2��]mWKni��>��4����E���`�[���A���Y�&�JS��n�%�������=s���2ky����tƂ��|�y�S�P��B*�C̡��Y5���)R�|/�����Ɯ>�(�V���IYxElv��;M��5j]j[u�3��;M<E��cO�^pj���WuŠf�%�QLГ;e����fىK��Op�ɺ�^*͑m���A��pY"5l���в��_�֭`�sC�Q����ԇ�c�u+�ɗo;�)n��b9�b؈�f�m�O&�W�����/������;tJp���k_#"`=u�����u��;�E�W��2�'r��%��>ٴ���=�6�m�z�'I����2�}.��'k vh���r�X��~���>�\j�j��%ջk���k���Wȕr�s���L�g���<��}�V�0�sKi���@;��$Xh�DmءZ��t�X�q1��-'�Xr�E[.�U�g��E�a��*ы�Q3�v����{�u6[�e��r��{�˻�f��Z��]�;�[��_e���^��E�L�	�:�$�h}@$kSK��u�'R֙u���]��9�f�=
*0gBy}Cv�R�]���f���`f�5���i=;�q���rk
du�S��r�����y�̓�Ow!��wvQÁ[������Oe�W\�Ҫ�p�4A��3l*ղ�ޗ|b]G�� �G7(���>@���Qe_1&��8����Vd�ƅ�*<�y�r&�S K �v>�q��JJ�����uY�f�*.(U�	_J�|q��k"0�wv�J���_`��2j��R��"����K�-�:r{I㹈�a'm�AY�l����]r8�;�����"n2���c]�܎�2�#'<��$�쥹�8ug%Sv�8�;w��/�J�p�[B��{)�@2Y�ы2�����B"�L&�1ԫ��X;#�Ni���V�@9�/6���N�J:�R�VdO'�Hu!�c`��m1�V<Tc�_3�u�B��=��F7�������uQVgQY�X����{rh��ui�u5���alж��F���p��>�c.�]J�֗jK��[�6  =泟522�:K�4��yFp���Z�Aә[�P����u�����@�x�s�Ž�%@�	S��Ź�kh�mq��Q,0�:�[��e�C��J���{�)Q#��D��Z��&;/\>��������eb
ԩSr�,l'IFs�}�>X�q�u�%eck���y.;�U�L���w>�ȼ��W��t,K���G��d\�ʭxu[y�.�̷\�ᱣ��V��ࢨD�@���K����*y��*��G���[��\�G5*�,��þy9bt��g�2�Ub�ә��\�i3n�@��`��ڲ�lE�0���suU����@KLխÝ��sϞ�!d���T�J6�D�3J��YM��>k��� �����4�w��9-�;1!cjmJ��N����C����;�Gfj�6��Z�o́)4���)y��0�#���ג��|���tm�D�b�%sf��nּb94�+�\ba�����H�zg]n�cb�	��n�]�jA��urh�������IU2��^cT&8�$A�y>)n�x�4nuk�.w�,Jﺬ�=Nq���,`	υn�3�V.G�a���ny�w"B�����osym�����B�$)*4=I6�ӌ��#)%P��HH��m��K*��p����h$(+	@ �]W6(�ͪ���ITEA��OS���50̕��Q,L�}���o������W��������������h��)h�&�(��**"��"Ѣ�ւ��<ɡ�����z~�_O��������~??_�J�������5STԓ����h�
Ѡ��H�1�DSITF�H�������QAEETLDQPTMUPTyfb�"�JJJ�(�����Xh�1%EM��N�DQLEET�T4SA31ԙ��S4QL��T�D�5U4��TAբh�� � ��ECT5TƝ@UD�EDEUEDQ5Eub���U�w��Z��N�S3T�SA��1AEEPu�SQT�QITT�S%U^�T�&�j�����b
�.�z�f���H����(�	�j�b"�H��D�M 
[ }���hc.��f�Ǌ`������pV3�HƩ���b���]�4�SjJg�c��MEj3��10M(On�r��� ~�v�����^����s�������VQ25�F{[m�w�P~ܥ�����D�6L4��o�%�P����ɵ��Lq�ʜʫ����Q�<�c�0�@G���������OK�Ү䶊&�ODV��>'�ٜz��fb���5\�6��:'�v+��\
ΥA�l�b�T��ж��7�-=�=�����l�FPj"S>����o�g����=��o6��]{׏9K����W�o}	z�_G�s���xp�uf���f{}���]��������0�ط��}�1wq]�?9���W�a��C ��TUɫ9�;J�7O'{�v��hrY�lt���62Z����	L�&�jM��G���s��"%Nׯp�CZ>&�H�nm��e-�n��׍�ָ�DIС`ۏ=��Y[s^���.�84�Q�Nڣه��q:�)��j�<���'�h��]�n׬f���3`�o�Y���Mv�ƮQ}����<���qG��ȵj7���\��t)�f��C��4OrWyw��>.
���Gq��0mX��[c,�6�f>vl@��N�@Gc64�8��Ѳ�Ͽ}_ʂN/d})����}6!��\ �|�&v}��T9J4����+� jׄ;Nw�9�V?Q�Ϋ��*���9��T��p��Ӯ���}ډ��ަ���8��ۻ$�W$T��{n�H� �H@~
=85F���1�8��z۶ Ŀn�zo���<h6�O��u��|ۯ��\ �-��z��-�:s�*c\�#Ȟ���EJ�r��bֶv�=���f��x��
{*w2��'��t��T�f�oKs�;|���Fhݫ�KBd�[z�V����;A���mfT �9���b��]]u^�J��������[��q=;��n�}n��NXH�0eU�KϺx�ߖm�'1�i����ۣm�Ǳ�uJ� ���۾��7b8�+N%N��;{����v�O5�RM٠��pu<������W��ܒ�I9�iMk9�N��,�u�H���G�Jd�N�4n��y�{����7Ɗ�V�,2��mu
��ެ[�{'I�$�E������ �բ�wo9<q8��|�WK�Ǣ�6&Y�%��{��]��T�=1�-�"Z�;����z_i�9;���C�l}jOGN�i�q/:(�S��;S�s��Yh:�n^(÷����1�HԈ��{�@3��t[��b��v�6����xG�-B�H� =�������yp���#��
�V��Ԛ��:�tI�;10���-@�+���ߑ�r��)�}+Z��~�����  �|����V�q��0��@�[~����}֠�k��pWa���� -� �.��Sb^��E�F���9�|���oU��@A�Twh�?Sx[�	G�+}Y�CE��J��'��s9����5�J�xF�J\��kq�p��g1�²�#�e�Ί�uA(B�V��l$o�"��3�?����:*\�S��t��g:�K���83���c�y��n�J�-��J��W�����Iu�$7�'&��^���~�
�Ln����_%�W<�T��lNE�M~ҹ�I.�i�֏,���BOP����TG,N�[�Ɵ9
�d@	0TQ�s��9e��I�J�Փ�p����L�vM�����8�ݓeq5cvE8��b�7�9�9nh���#����J�}��8�y�\���y��鮶͢���Ԫ�e=�v6@a���\w�
�8�����x}���}�C%�k#&$��ґ���x�,�o��X>[f�|Wdv+{�er�ȑ�>:=� v�q�r!��������ݻ�s9��|HO:�|.��kOb��Q�M�C9#A����9�����l4pc�>j�v��9[mQ}T�ڷ��v>�J����>�i�X���&��+�k�̯��6v�����R�Ѽ]pZ<5[Ҩg����L�g=6�����{�<$L�#����9P���*��Q|��f�[C�[ �(B�JZ������B3�^�)����OT�{����=y�G�u���U���O��;�H�ܚ��a���ء�s��o�l6�ރ�v��� ���.ƛ�R.i���<���#�^�of�5�L�iO!����B�RT-)U��{[�3�L	�[��n��\Ǚ�F.���p� OMOk��Tn��S�l�0�����lh\��<O�nB��=%Ǒf�2� ���T�,��]UB,�85K�
\z�����q���k
&�8�n�`��09����l��l���b�̆AEdw
�]�66N�U�@�>���}i{�z_��85/j��xG�a|���T.$�����zAr����et+�y��݈/R��\yG��T W#�\��ޔ����j�Ճ�eO�b�`���#�l_����9o�gQ�Elp>Z,��\Z3g�e�Įh����7\W����vls�ɶS�����n^�������Y�`�w2;5��ם�:��$L�-�������~X%;���,����Dw�"��O˜�D��@g<�wdS�m�z0ok*z�F�2o�"`п�IwH`�'η��t���*C��Wr[ްRW.��nFR}����`��B��f�5�"A{ǜn���ο
.��[�^��d��ح����%����w7�w�5�/L�1i��΂0��\z��O�Q�/�7;�Ձ
��n!n���ܺGE��Pg����;�)�#/+��f6���]q�_��;7��}�A��2�|1�]Q��,��8|hD�6���{����L�Qǽ7�'�s�Jm��7d�9�.
�r�ȝ*�6�Z��^���b�ǖZ�㵱*���z�N!���fG�]mf˓���V�D�x�:۝b|��ow]�;,�A��V�|d��;y�Y�����7���+�����LzH�=��7�z��n�R�7�ht��͌�p,td�%��!�R:����(��:,��@�H7���&Ѱ��ͥ�LQvڋ��sQs�:Z/8���� P[t���qd�ɍ�����"�t�v���9���9�����Eѹ��hځB�.j�����\��0�b��-�N�cl����!�#��ת�ͳ��?S��G�����C�U�H؋�D7��^8+Oy/����"�����=£P�t�?���ssj0]�{�S���kK%[��-�\h6�q��	� 6c���.�,�EOEK��\�6`܉� ��Y5��m�����V���b��=;#���͇ݸ�J+^���&Ƹ�G�1�z#�c�z�Ɗ�&�#S⻵cx6�sfo'i��gӭ�b����7��Q�*��W����J�t$���v
���۰�Ə\v��,6=r�̡S�v]��u�/4ٱY����#.�Z�n��E����\�X�ܖ��3Z;k:���G[6��B��j�2�$(M[����Z;N����vWyy���͞�=NP���G���A�������F��uB��%V����� �Y}\�%��Lt6�?$.�ɦ�ћ ��������T�ǴU��V;)��y}�]s�3zt�*�)�졛!��͢��w��K�@`���1S6���]tk�����<[ah�ݤ�a�3��:�s8��
v5���&���-�ь�6_��#�tf���H=;ͦx����Fz��CKѤq�M�V�\Ѿ~�6��q��y扡��//�w��u��O�?<����r�lK����}�"GD�0dh�ov��M]^G�<��u�a�Ҳ:Җ8���y����798��t��O^	G��z�M��d��\���:e��狗��G�w���i=qQ.���L�ǬA�a��yv�g�,��:�,e��km�P�#���dנ��$t���wo'7�3��u��N&�[)�F���\�3D=�G>7+�fݠy�]3A]e�M*��X�ge�e��R7/$��	L��;*�L�:�����Y/m=�\��:�^l�����7.Vpt�t���C�> �0���s8Q!�4#��,�B�zf�7��a̓�u1��e��.�g]��#^I)���|�M��U۠S�u2S۽ׇo[KUv��^pO�gA�B��ly�)y�L���l��PO�W=������v�=W`;�C����2��#`V�U���+���*x�mD[S�b�wK�����'��UnKޭ��0�.8#����\g���UY\�ǩ�Ll���mW��Z��쪭�#2�(g������yܷ�?5�3�.�7Hw�<�s���^�w�]�s�0��^q3}S�r��.׷�{7c^�ك��n����=�C�u+�;#o���'�0�Z���y�xd:6��t�+D8�.���H��Y�.}ݽ�� l1�q��N9֫���:d�4%�r��2UmWX��&��-� �x;�;��.t��q7*�1�p.4Y�<*4"��m����7�=}�`��#�)�5�r���ҟ�2�Js��c���^���C6��WJ��aѦ�p�R�`��9~������uEQ+=����?0t��U��tH��g�G�+�5W���;.���1,�pN���^�#��F�1y��2N�o5䎂3M.͓;V�Dg=0�, (K}�����d���ͥ��Nl"�A,����ּ�H���!e� .6���w�9i��������%�v�Wןq�'O&�^Z��x�j���=ܛ��ك$ �Ou����s`���R�P���%���/c�ө�g(LE[k�3{�,���O�+�tT���Q��+){������4Ϸ�GK�oR�PO�4u�F�"�l�
����,�i�B
F�]^K���RZ2�����X��=���\J�p;����Dz���JJ��4��[4�X*�C��z�tu7l���A��Z���s8h��gT��\qlmm�f�l��]�:�t-��@ �qC����s��1��}�����ƍ[�� \_��)~�ػ	uw�]�q�����{�s�<�i���>ha}���£�p�%]��2�r$�~��^#�z�g��D���N�] ��ea�!>�L�3>��	�:Idm�νW����s�h����:eGf� O�YU�.�v���;����N�^߽;��EN�Ț�V�M���.����A (c�F��]&:�;Nn��K�;8���U��6�smw,��`��+p�{��3l�o}��{k���g�Pg����Α�ce6���X�(��
��f�&�昁�xob�[�)=�a>}	�`8ղ e���ܧZߟ�������G���������O��c��r�l�W�ʖ`�b�Q��2��������}���Wk��$��ǅ�l73IƄ�<5��K�wnq��ȗ�fo}���8�v�}�H�,`� �dlS�P;�
�3�X��bz�oX�R��߮�>�K��ז�O4��#�k�zR6)�C^n>�_��]��N��CU_<7�*��$$OZD�\�6��VT���وS�)���'���w1ޤ��_�+}ow2�5�N'k�H[C�
E(�}�z���r�P�h�>?Zw��~��ُ��\`a��5�<!v�dk�ue�=4�5�����6l*����Hn�7��vgV\)n� �sS��<}�C�Y�te��j~��]�{�@5�z�ۜd���]�ф+1[Y&_QE>�;��p].�t)]KݛO�(]�yĚ;+�0]N`�����W�u�7Qw����&u��j�l�B]�M"Qv��Yp�wdV@&v/��F�8ܖ��m�Q���`@��v{+Q��x3���=Un)(C�*~��V�����6���r�ie-���J��Ns�eM�z�9x]���l��A�}H��1W��g'
�9U��PQ�\l�2��PI�Zro	h�Pt�\�!�='BVY�x�|/�W�OS��aZ�-�Ԥ��Ǵ�M0c�ښb7��A�F��l��A���8:���M�f_�ʙ�ʇ9���ߢw�]ۡ�����u�C��.�ړ����:�AW�/i��d��bw��քbm��WƠ5j�Ε)ƽ	�9�tۭ�mu�W\|UB'!�R�<6�1 �ܙ|b�Ƿ��o{��N�P�sC���*p����-n�H�c#�TX��.��U諝򡾥�Z8P�^��pSQ7����%WPdJ,Z�2N�"��S�d�ѧz��ϥ
j�$=i׸t�/�ۃ[�+sv���"�k%��70%\�V���+(K�usZ�ER`˭�g�և��&�C�u�L���m�>�֦ ��N�`�7	j���{ת
�@w"j�mT;�VXN�O]�EY-㹗�0 1ʛ��X%}zE�y`N�Z��m71��}]�JJ
�ae®�EB�ά\�b��F�5(�t؛��V�@c[[����mWU���������;��b'\r����lnN/`��|���L9X����b�]p 5�lU�vd?op`m�o�s�E���E��D�p]�A�4Qh��� �U�4��@��TY
nw:K,�mw$TC*�u�v�w�v��E��Q���7��BϦ)aU�j�_�g�>%��F�K�&H��9)�+x,����S���A.uw�<5���}��W���(�pY�A��%�l ak(U��ڐ}�E���fol���<�4�q�"��vV�px\�Ms;�x��/4�١.��ʻCH�Λju����	���]*��C�P8I�4�Z�hz���QU��.�Sp�x�[%�9p&c�Τ�ܭ�}'EAvШ�j��l>U�_U�
��ɀB �l����R�V�r��J��w&LGG}{�:�S��|헺�dG��؊VN���"��붹�5-����q�B���Ú��*n�ʱ]s�:���P�xd�Z���T�oya$j���ר�1�RʺG�^�ڔ�
�nX�g�i�oLr���q.�g�*Ô3�'$&96��ҭ��a�E��v�d�O�����U����&\����%�Sp�}���e�yS(��-��ų+��i�g�*ph��o�]�ٕX�]n�^�꽒��rp��PFFe�E =�LE%33�i��1EPT�j�:ؠ�����5���O���������>��5MAEE1U,�D��QEAQy&�*"�(����}?_o������~������(������&����آ��IMP��MZ�ITIU�TP��Du�G@Y���w�UMLDwj����A%�&)��)"���(&��
Hi��(��*b������ �������54S4�Q��S5L�TRLTQ��TE��DE]Z������zN�x1AST�5RA]Ɗ�%��"*��-4�ADUM0U5Q��=13LETMSHMU]
j��h*������������j��
h(��0R�CI�QCE4�M$DEUKE�� �*��uj7#4���9��&�N1��>�O��nR[\ �f��*�FTf�V���1,P�r�L��V�߿}_ٞ	�~p�m<_#���W��4EU>��u>\@7�*c�5��WB:��r4����m�)s-ᑤq�<M����x��@��S�3��"�A�]>�Z��jh��p��r��-mkd��9����e:SGY���_���;ZF҈[B7�O=�対6���+�}6_�`�ݮ���Z�8�<[Z➙��� ��������1���:귒ڹ�h�cvglG���٘#�|�u�o�50q�# xl��y�E��՛K�'7 w>����	��D��y.�;��l������s�b$�u&��Q-ϯd�:"��d����Urn��1�v���1�i��qG;�ٍ�J�TE�I%�͊!��:�]��}g�GH�m<K��G��l���u9٣[��8z���Q�T �/4�gh����$O�"�if��=���\�u_;�W�>�~q�e�S��7{B�����a8��Y �23��9hӚ����H�T;/9����a֮ʝ�2l����F�f���軉$�7.����f���ԙ�>O	�Us�o+��������7���O�b�z��tU��`֤>gʽWT/2=�$:�����9����n���}��wa
��5�n��`�è�S�"n�z��:�{���fޟ�9;�oxB��u=�jM �kI�*%��g+�c��;}���E��C+���b�#��V��1s���'��`����駋�[ zoW=����kw�;�8��P��>��=[���k����RK��|�#r�b2pe՘gW[�[�W�X�x\���j,3�� ?��t*��I\`)ǽ���͎h���=OopX��.�!��a!�/���ѷ�(��\L��T��{^�,�j1&9J�,�xwOHa��� �n�к=\g���*]a�1�+9�4�s)�t��N|z���vlL)h�m�H`��odBO�������m�٠��-w{r�O��*;������`�-������Ug�w�':ͧui��ȇ�1a�s��[rFIv1���#2��Zuj�oS��;I�`=����ܱ�L�r�TOlTٴٸt��0��o����jN�|*���v�gW'n�ku�g)�,Ѻ��v�<�1q)J�,u6��e�/y��wM
�MZ!U����^��q���`g�<񜇡.�=F���˛+�/{��H�M��[.o�Tu�;35�,같	`;1�q�o�VrZlF��1r	��Σ�v��3��31�.6T�FPj20s@�<2��(�k�V#$���ݍ�,Ym�isݵX:����6+uS��b�Ψ��7������y��22�����~��͘qh�ǚ�Z��Ẃy5�>��W\��q�L�ڹ�4>��jѹO=��>9|"kW�J��D��Z��}v��J�귙�ȼa�ѱ�M+����^Ȭ���]�AN]���/-H��3�� �bU[�^�+��/t92�:��w
��B��|��aB��Z�[�I����~˫��5{�]����0ίY�3ә��wFy��.�Ao�-B�JKQ���Όᵩt��dF�뽖�i�@VQ��p"w��K��[~�ij��p2(z�	���9�`�U6�6��ћ.�a�N����v�u�1��<l�����k.�$*9�������g;�c�F��Y��5#���CN�!5���K|\+f���GrSi�g^f��OK����9_�t��NTuA5Q���;]͞����gAdv��a��<{��vl�S�?�*�9+jx(�	n��싍]3�����,w5���e.2���bl���[m���T���bi��uU���*���=B�����V�3�I�Q�������o
Q�%���:��'P}���m�u�ymVbE,�wn������Z��4�i�h��E	�UtȈ��	�g�o%�o��SrCW�yY9�.�g�٪"�:��b9�c��"�.�Yԛ��v+��_Mqnjna�N:�k0�98��%&Ў����h>/	1�~�.�O�z"T���VL;?B׉����O��BM�>Ѳ;E��k�Ձ�³Wr�hKH���q�~�g1w
�H}��{�"x�2���^7�Yb����[�Ջ���/wn;��rZ��ayK�jLwo
T��˘��S�NQ`�Qݘ�w�m�@�̊=y����C|�޽d��w�v�s��.�@�n��4;ɽ�^ڣ
QAP���x:U�ܥ9ioX�켃�1+�Q[�]�,R� ɗ�ŏ�ӂ���9=^�1m>̡���j"���hL�	���v���j��/7��ە�rn��QCD�v�����{��Z$�4��s�fr��9�]���tl^��,�����&}�8�s�Ey?���yY׋PΖ#�g߮.�dK~�#�U P����v�mY�|������2�;�#���JUB�;w��M3���:+�^v;��3�F�7E�p�T!��h ����^�l���*y��uӭ7 � ���u������*:��w"�����hҒ�uƃy��]@�3��s9�x+�=����D�_#��V�U�h���\�b	>�q�Z�[/,�kϳ�LeoCV=$.��ep<�7�!l�7���L����`��<���Y��B���y=ɘ�=D,�9��۽�ͯx��"1O�gź�:�5(���=ױ3;÷���n��H
�'i�z�ހ�1�[�-N�x���O{xE[K��F4����}�T�[󺵙�б�a��1@aH�G��]:�c��U�ӆ��,�ܞ:@����wz9I�yD[;�v�KAu���/��������EO���ޘ3�J�(�tm� ����o^Il��y���qmW���UF�l�v�ٺ����op]s�<D]�3�%�;��1�=���#�v<+�c%u _eW&�c���Pc���Y�{�흫
ڳ��=V���Ÿg�4!jT3[`_Y�����j28����<FZ絍9�ρ�H�OR�#��i�9Cתl�7���:	DL";\�o��3x^Nu1�/g�6mΊyL�/�ϖ�����h��b۰A�,���΁Dm�	��W��ס���PJ�OTM���<�q�M�Oz����V�1(���mIK���xsC8A\X)e8�ͱ��%���&x*����V#�I}
�rt_�L��UG� ����c�����^�]e���&��K��Fh�դMmym{\���4]���i�-p��%]v �J����gy�̧�M��[���?�֎/z3�#c�"�A�xi�46�ݡ7����I_*�#��I~>���{;M�֊Ƶ��c"K&ALʞZ�7G(���Δr�qWw����~��*�� !�(*�t���KF������񗓱@�Frf�xrt{�א�"�����;�ڴ���.��n��O��͕�c�4L�E:(�����/:Ok�T��qR2e5S�l���#ΗH�#kL+|Z|/���f}���Z�k�nT��6�==!��L
�~�Eq������E���.�e��rX�Gy�Q�h�8y������<�|�_V���m�-��ˆ�WE�����cϷ����rW�ҕn��=�:X?��9��N��殮��GX�Y3:@�4���ڲ��u(�U��Xl���'vҡ�>�P��s=e�8���	�N7`8U7�tg%%���{�H�I����b��G)�>�u+�vUb��eC8�`��x�5����k��Md��׋t��qj�;o��<�7�Vރ#���f®�EZ8��1�hW�̹�3c��~���:�k�Qǚ
�5��}|�0��I�f���/��{�$C��7wL�]�xP�㼍f���a���ߦ w������
������U�਋0�f�!�֧"��<0M��n2��7W��!����y\����o����.'s����O!G�����6-���O1ҥ�5o.��)�v��W;�{�7�Q�S�����9x�˄���`���w��5՗���{Nq���K`�O9;B&�^�G�{˳� ��oc^R����cy�J~�RO;�ٹiE���R�Tdg���ZR�uN;������V&��8��~#�N�ȷ�?ޭ�-B@��"�U�\J=�݄f�爱P>��x�T��	����4���Hʖ��%\��=��%�_K}�ڭ���ggM����z������Z�ְ7L����]5z̒��ح��2�<u��h�1�ӳ��
�H��dZݞ�����jp����ڦ�'{���f}�rD,ٽ�6Sh�+b��<�"�{Rl�R5 �wc�N��D�7w�c�z:�yB11^w�1���qʠJ14����6���u�=�F�3i��`c��>����;Ӫ��K�Q�%iD�KS܇�f�¹��V�و��_�T��FϘp�8�S~�]�T?�?=��/�0��}���	���(�P̬�I�A�]D�	������Lm˙��k�R`���cU�u�|2���[e�4�{J���U1Ј�.�v��a�K�tH�Bx�vں|+h��;�@����j^��ͭ�X-�nw3jE�P��ub*�ϻ��z<��6vb䑻Ө�+����3��k�v!(֤@���'v3��D�������a�+���ܑ��+��A�����Z�LR��"uF�c�]�V�|F`Ƚ�;�8���V
3�O�2|�T����Wmk�M��3������GSP�z�葺I��E��v�NcO.�oq���{Z1��xt��g��L�.ѿD�^��z�C��m��h�����U����ۖUw���,₸�Iv�M�8���o��Ld������8��z�'�ѝ�KA��.n� ���u����j�|m��%�eNo��/OK��9Ua/�=��U]2�Ϋu U��)�ZPb���z��N�e9�Gi�J�7F��b�����<*�j�{."}�
��V��r�]ޭM��]����c"pRU���<��T����6�O�׵u�����N�Ǟ���l�|���C����w��oD����)<7j�w�@����圕!S�z]u�Hj63
ŵi��4��J9-pV����_s��[�30^��5&iq=Ŧ�W3��B���<����[hVmKR)ۓ)��dq7�"P��u��z�s��-B�>���g\�jh�%MT�X�[[�*������ݺ��"^�r[���#SvzG�b���U���&c_t������ �'h��%�[��~��;v���q�6��&�C����gi��1��.ۗC�Vc��W�6A;�(i@UQ�L fy��6`��pQ���%ߋS�=F�kb�j[5j�er��s;��N�m��0}�(��ɠ�γ6�b�e���ә�丶��ɻz�/'l��Pc]R��qa�����g`���A��/'-�SX��>VЄR���XqR~��Žήm޺%�(�����)�M���v�pQ�0�xOF��ةN]19�S'���,Y�kM�F�i썷2�=�,Ǩtۙ�����s]��5u^����Q��y�����ه�f8W�0�ƸHC�I�6�}�aC�H&�V��}��uUEgԠ�����є_�Hc�dU`�>�{�̋2��@!�eV@�!�a�a�d@!�a�a�eXe`@�@!�`a@�U�!�a�aV �D ` � !�eXeX` �P!�`a@�!�aV �!�a�`a@�U�U�P!�e@�U�D ` � !�aX`@�D!�a�@��C�
a�a�a�a�a�&FQ�E�A�A�E�A���E���a�a�a�a�a�a�a�fP}��{� a {� d `@d@e a `@`@�8@ P @PP��� d@`d 	�� !� !� !� !� !�@6L4ʀ� L��4�!0�20"2�]t=4Ȉ*�LL�!4�(ʈ�0)10�2L��0�4�&ˈdW�*C Ȅ0!�P!�aXa���VVV� !�a�a@� C�2�0 C
�*�(��������~���B� �� �'��9���1��vT���������;Cg���G�$�?/�Z��>}����Q��O�܂(
��QX�������bs��O@�w�����ˬ7q<�Q 	�0�LC��A/P'�Xr�$F�QDX�@
 �� � �d�E�  A( D� $�$, ) C( JȀ�  J�	" @� �
 H���@��� ,(H�� HB�,�@B�*� D�R�G��������O�PDAiA�@(
�G�o���_��.���u
��F=�EQY�N<��6��	�X?@���:������S�Ј��������_�>H*���UE����DP���z���+��������=�F���7�='�=���:�;DUEn�>����*���)���Hr;�5e�n6�'�P{�ETW����ETW��~��?o�v���<�	��Hd��GO�5�%���"�+d�Q0|�~ɐ?�;�|�������'>��"(
������P��[�~�P�O��d�Mf�Ij���f�A@��̟\��|�笨�I@kR$���UH�$�U*�*����5Z�@�T)H6j�U)(!D�	SF֢*I���BRkHʪ��T\�M��i��cl�UF�%l-��!���T���0�e-����T��iU���ckcm�V�,mdh-m����-!V�TZ�m#m�v���S�K����m��j��mf��l*�M*��h��¥�kT6�4���A)�ZV��f�cQ�m�,ڲ�ڵ�kV�h͵V�kղ��5Zh�R���M�kaJ��   3��ԫA�L,5m�۬�m@R�-f���*��7M�U(�,�/����\�M����սw[�Wr�Ҕc���޻�B��m�f��dݍ�Й��   �g���"�H�фꛏO��O�TdiZ�Mtn����x�bو�[��6eZ�w}���%��ڟn��4zt��ӵmAm�VۖvѶ��U��J��2Yv�T56��糃��c\�(��k5��f�6�l>   ^ХimV�w�ެ��
�mdu`�fTi�ݫ��2Փf��9M[T�bwr�/VuuJZ��+Cb1T.���e�VP��F���Z�mmU̫f(�V�Ɩ��fի'| ��֣����vR�چ���;w5�mv���5֩���]GT�5lE($���QCEN�փւ���w3T�4��j�PkZo� sx=U��f����HѴiUB���l{u�f���5�3{�J
Qt;��6h#vpAtQZ1�2R�E�Je��BmF�cg� {�PH�����]�v� N�aM�8t�9ٵQ[4�c�۠m�:��45<��TG, 
;ݩ
�i��YA���Mi��5�ٗ| ���V���x�Ά�֎�i��4۳uZEUY��ǧ���{`�S�Gv�;s��zk�t.w��Қ���.= (�dFl[���d׻��4i�  -π�P��u�Gxz {�z�kl�/]�裡T��=(GB<��z �V  z���@�:�+@<�um�^u���Z͚�d[L�k5�,�   ]�  ׼@馀��8� 
^�t �����x =-�U�t ��^���v77j
 w���w[�q���)�-�՘Ֆ�XՓ)�!�   a���Р�e�z ;�g� ���=��==�� ����p U���z@�m��ҽ s�w=�k� �)�̪R� 4 E=�	)*��h�B)���2��z��Q�&@E?��� &�jm�%T�L�Ѡ`��)6UR  �O���F�ߑ���?o۽�7�~�g��~B�>�������;S�g��{ݹv��@<�m�յm����V�����Z�����ֶ�m[m�������/�<����z�鄿��)���<���h����j���AGwuxq�k	�*j/[ה�xE`�2�;Ěp�I&�F� �l���!��`��9'�x�#K�� U�m���������ᧃ[��e��CA��&n�����G��7&��4�/�^M�ǌ��S�j��Y�*l�2���EZ0Kt���<��3�ܵ��X�e�Q	��K&yB0 OK+X��tK�aÆ��P��|Ĺ*��t��M�Ksu�Z�Y��L7V�V��b[�(�R�oV�L�I�����9u�Q���=�F�2�m�{\-H�^�룷{�:��t+[����������X0-��NStnM�67+1�J��"��'/f����݂�r)����-��J��Ws&��c5
tm���b�ct���G[wY�WP5�i��Bh���؉h�W�c�i��4^ �1�^D�0ިie=�l�Z�I�+����i549%�M�\��1)e���Ǘ�6IJ5�)C
TJ^61���kChY��/��X{�V�VK�A�6I�Z��p���U�$�u���Ƣ�}a�Œ��Nj�ԗX���n#H
���v5�	<݆�).�s���C��HnZ�t���`�MՓ��^*��4ԤUG��
�	H�� "6��l�S7i��O<�qA�3�k#�"��؎&�6Fpw�[����L�tdT4�tf;�qѳ��{Ki8�T�fV@�QUu5K�i�m<ȞY�7e�i �h(�
���r�U�.�ՂL�B�J�z^f�qjU�j�>ŏKN���ii�[�e!Ib8YuM*�7D�`���q]f�P談Fհ�r�+5�6Gxd��5�2����,X��ub�����U�b��f�<�/��|�jO>�,�uRYkQ���4�m�(�}�7t��>�3Z�R�.��W`V娶�<�\�t
Y�ܱ%�6��⺏6@�U�i����
.�Xuy�@V���gf&���䈹�ݷ%���Z��.U�ř�z�F�ظ�6P�pY�9L��YwKcZ�%q4�-պ�%���9Lq����q�Vvc�j�[�F2QX�����ь�+AI:�/-�h����n;�NE��lKD�*���N�,
f�I]b��]貀:��-VCJ0�����4��Ę{BCF^Ἤ��@�1�M�V�FZ"ч/�e�Zպ
��${����t�X+#X�ӹ�ì�
Cv����Y�3n�j�ث��R�n=s㻙r;��#��h4IrC�̩��u+&��z��%eE�x��SU�X��r�{M)t5��-S���V�kU#�!!3������@V���m&؊Hp�pS�Wb襱��TŖ�X�em�Fq^X�u��q��ܢ�V`֫V`Z�ӹ�	�"�@)*L/��Xlj֨��,U�'���5F�B
�fG{-�AF�m舼�
&*�*V3)�:��T��Y��iʽ[5i)�r ��KBlqnL�KS߅ԅ��
�[;Y	�W��SR�ЪV�r�5�e�q<t����J��w�v��v
p�1�a2�,���y�X�Ӹ�����9j(�^[mRדoS���Z+[m��m�"��fP�6��h��;��37]��L�"��ٶ��B��3,��Gm�弗�
�
�>�#N��V�z�I����E9�凒&�{��B�w�;�+`�D^+Ҝ&�U%�ս׳OH��sF:V�ȶ���+e;��Et���L8�h�橡���n"e<Q�[	a�����nȉI�����s,ސ��,�w��� Ќ��7������r�z�֭�z�g���R��Z[r��u$V<AK+ڈ���5��`��������%hnX�:y�Mt��9���5�pM��EA�Zj7b��Aܰev�1�ⲭ�M$)k�A�6�V+u���h[�D�2Fb�*�ݖ��%�rFf�ͳB���6�ͭR��Z�n����-��r�vؗ�����Su�B`⡹�B2����_a�C[̭���]8�+mQg���5ǎQ�%P�j��-}m�K�Lj��S!x�q�iP���7K̰�������:R8������Ln�-��(Խ-�{YL<;s.C��SFJ�F��2ӡ�j�ҥ)Vm[1�2��Q�R����,nm�GLX�m���׌�gkc��iܘT�H�pɵ���k�FPV@�cȐ�6Ӭ��.F_@� n����i����eb[���K�/11WZ�:�#̩���X9���n�$n��L�l^�9���ӑ9�ظ���Y��L�+�ęc'�Z�Z�b
�.Z]dP�Ѥc���N��.�U��܉\�Ԥ;O(旻�b)�ao�w�ެ9�h�[�6V�0�Cq$�M�0���(e�*j�n�4�P�޼S.��(;�����}n5M�A2���<��4����( w�YW�pCؽ�g����^�P���
9M���Sj�y�X&�T�bFk;GI��1o�;�80�w�b�4h3Ɍjզ����[R-�Z��oJ��B���9,;��� r]⎶��uWnn��ӊ�hz�ɰFἥj�#sQoK��
���J�4�+ُMj�xp�CY�CJM��	l/]��]��·N�Y��ׯC͙�bt$80�V.�P�J�%,���e�]Y�ɸf7"V��9���n�^�[X['sK)���c4�iT#��EQ��*�df�A�WQ�&�)͋)(���x��9�V�E��6e��V۠��Ӄ��*̣�+�]�x5fB�h�eM��DY�5[1$M	id,�TvUƞ�L�x�Ta��!I!�C���c˷�@9�ㅀ��t.m��qM�yI$\�p�v�VJ�	��KWM]LH2"�ϱ�u3�\�V �.�e{22�Ţ�)�����p�������Kӡ+��QsV�%�Ot\%,K̛,#�#�ј�Ce�:hU��U�Z��O��[�eB���ÅЪ[G%<�,�:3e�Kl���M�JhgU�L=t_�T�#.�cv��HZa�CY�r+�wVܧk�����#,E�v�(�8l�W���M��t����!�兑:P�Wg)�<[��VKtEf���e�V�۶��Cn���N�ͩ4��xV"CW�D��?7x�LJ��s CX']�2��M�4cH5��2GW�-���4�(�����E�y�t���������w��IsA�Җ��/[��[�jz��fW����l�W��8O'�$R	%�85�w���n܎ r���q�̏a-�Xx�%�ʖj��&4ֲ���0����V#��"(H�O%Xն���2
1Sec8����*4a�=����a[�yb�݁(b� �.S���(,�Xm'����7n�d)R3�&s���֝�5ֱ�1�iW5�-�j����$�a����.庥ti@�I���[�0\ɹJ�̦Bof:��h�XQ�٧�<W#���v�m��#5v�u�ު�Hm*̈́�1+�6"��Ze���˚���ڱ1�"�4���)�0cv�:�W��4^�t�'	@ʰ�ku2����b��h#,�V/�O1�S��#U�Ln[�^�ͻQ^ə*�&�~J,��� &2n��T��{\
T�X]��.MK2Z��-Y����9�� �g-`X^G
�[gT�2���T�e&[���/M��#���9q�Ɏ�z��q]�4I%�軽���SJ謱�ى$G7[E,�k[�ŲUҼ�BfK�	�5̗��TU��/�*4�
� `����Nn��6(UJ�MnA��d8f���&�m�,;V Օ�h�y�nؘ�D.}�VO�,C��-��Q�j�(j;�N�ؐ��i6����
�u����Ơ�A¬P���e]� �.�1*VU,вX�kl����,ԥ���@l2�յ���"�X��
.���"���N�֝2L.ӷ*�$3I�D,EШ���Z,��lT�oA���^1j�bo;��-iZ��ܣ�{�mG�&Pk�Ұ�h�7b��.�u �d<n���1ʘ�J�k�[��f�3�iՙ�j�2�n�^��X<{p܃Ӝ�rɞr�c�[7��N��t�ʶ�P�b:�bH�f
ݘ�C�ñ2M�5��Y1L�ۦ n=�V�Vt��q�V<nP��J&�nؚ�V!��[8Ⲗ(�:{N2aYu����X!׍P�RI�a�w!Q���$�$�,z�#�d"�&��������1}����!��5����Y56�jO�1^'�uD�c�i�8�-��p��!��	>�=����y�]�"K*3��9x��Ӛ�;���݂7o7$�(\km�&*[eD��4dy�2�e����� �+7>,<�+	�$Y��A��%I	��\W��d���ww�	���w��,�x��vc�4�`i곈n=�n�ӧt�g�j�[H���!i�ҭ]B�G��䀼'T�Q�j� ����U1�ZV3K�Q������)��n#��WT���&��n��A���ڻ�Q���I�cR�ONN^i�h(���}u���˺�#
��{�cC%;�s��i\�q[�ZU�޳�P���(+������r��Gv������v247113cѸi[e��5jG7;�e(R)�s����Z*@�j��w��ꍄ�u�����ۄf��hd7z�h],؞���b�D��%a`e��/E�.�Wrҋ �Y����6�&��*v�"q}��Se,�� Z[�Dbn�+��2��ޯ�@�GfV�Z!�m���k�EVݝV$� ����w��TE��,e`��@a�6v�_T.tep���#ͦ���vա1GMQ�Y���x����r�tȩA!��-!��̦���;�p+t�JT�[ݼ e=��'�2S(n�MP;K&g�\���,%��p�9X�5)�cU^ �z%�ʡ��d�k"�(�����Q�2��&�F�D��/Vkn��֐��W�k�-@�f�Vm^��I ��z�W>��C3kV��#(QF�Q
Z��o^���X����Thn�ǒԁ�%S�^�����yWX�E���A�&�-��t]�n�f��+�F٬WW0��4-�H
q�h1]D&Gǯ���oM���lp�W��uT4�2�Ӎ��3,�t���+]�/�j_����,xKa�*��n��eՌ���S1b��nDf3�(�ؚ�S(K�ɱ��ָv+��[�-ˤ�R{�v�j���S�Q4n���w�R�0����#�v=P�&�sM۠j��N����TU�kK�J#ah���9E��z� #!ݬue}eSZ�=�y���L VGR`KK �J��,��I�v�J{�ˑ�6�v�����P�����p�4X���SJC�������K���pmB��9�斲�1ݩM��咶��$iS��˻X%J[��S{X6�=NTn+!�vf��r�E*�w��,%V�YE�HT4�̆��2�r��vd�Hѵ�HZ@6��\
��h<�Y��R�V��7.a�*���x	HP�`A��p釻��D�L��L�daք�sB dWk	mc�fV���卷H���UH�����\�hap#$N����;��Rg�m hR�Y����,@̳L��4c�$B*F6��hX�㧲f���Z�&.qHQ�vU�/@*��P�*E����	IM.LxP�7Y����(Rm+��*n ;��%-:7��r/P�9R0���hF��#m�[[���[q�
(���mk�˼�-+r�VGތ�с=���&�͋��-Wx555�p�r%�����ʟr*�&��nY�J�U��N��b<�f	�F�z�&&,T����n�X�b�PSi�CK]W�*�$7UX�34e0�E뗤T:ۻ�Yf��d�pP�XF��b�I�mVh:�q&$�ESu�*͍�W��ԓVSC.ةOVf]Ҋ�`Bج����Į[���R�����1�v�.%7V�A曥!��-@�Mϯ�@h�4�B���Mc[�֔rV�S���ntp��c��Ь��.�G����8�̫n m��@n%e�����o�1:V��̰��W)֭��l4˧��J����*[��@B(=���Д�:H�=�.���єqݫpRDYX�wg�b��%w�n�FYZ)Y��2�!��e�[�����I��k�FN!If=@cԛ4j�Ӧ�[��	A���f'�*y
����ߍM�R��ٷ��F]PK����+-�������`Tt��B�xtX��V���F�L¯e�m�N�w��l*��2�2Nr��L�v�M�8p\���~fڹ�ͺ:EC�'0�,��jR4D5nRj[��DH�Z�5��Ų�2�Rݙh6qb��H9�����Ko��N�
�2\�	�t���f�,���Wz�`Vi�2Ҩ���3OhSZv�	R'dXŶ�����!�J)�(Rq<9S!�(I`ؐb�4���u5�q%>�LA75ov�<q��j�J��kr�cR�,����Yګ+u��VTɘض��i�$En�=XUd�B<�r�<fj6���[B��WYQ�׶��ib6Ͳ��dt¡H�xI�a�yǜ��c&��D����tr�!�yC�6�5�P�T�'����H0+0k���j��#fA,ñT��ۺ�Uf� �\��5)���*0qL���q[:��PM���Alԫ5 ��HB.���\�[G��Z&G�mYq�C0`H^�Ʉ]ә�������i�M*ej�(�R�ox~�>S��S�s��[n+v��,Y��$[s��oZ�콾�����<�τy9��0_+Tpp���1P��i��곔��܄N����I�=bۡ���CbҖ6����D�3��Ѷ��rta<�.-����q�3OX�؈Lܥ�y�"����ڛ�`e1yu%s����[,/�������Л�mѵu���{
O�q�\M���(�&k�C$t��k�J�ː��Et�l�W.5}�38,��z�d�}LIT��J��4��m#S�>�����R�네�{�w\�3}I�)���$��≡�J�Yi}�.��ˋ�ś���↺.{n�+Әe�c8֯!��bѹa
�v���͏nX�'���dq'$�ќ9ђz����ج�����]D�8z���*'&WVJﯭ�d��έ1O-��r�hKw�N�r]�a=+[<Z��BK��H����5�����������:,]�/�;�b)�9���6_E|<�뉪��2��LA�Z�^'�gT�P��=D΋��쥔���F�0wo�����}c�4e�)֡5ݓ�s7�mx�J���%��D=�{�8��(�*�Ҷ&YWR3D�fց���@2"��{]���սs0W���n{�z��v���B�ٱ,�oI���NP7�J�n=Ŝ9�v��]]M�(�Y� :���7�އk�s��/���b�/�v�:�o�v��ދ�g���Y�gNw
P:�<u*��u�v*o5�ck�xv�W֡��׺��A�Uۗت�\\�uD��$�v��Y�����W���"��h%��F���u��u�]��"��v��;��y��L��g���l�w��ږ�ƶ�_e"nS�� o�-.t�
nK���l��Ӝ�t�jfW `���^X���9�Ȯ����L�6�,:�)�w8�����; yS�_�n�Hҝ��SE5G`���mծ\��t�:��W�e��཈{K��I�t��w�%��wX���S�6]H6g!�5�B��/�d�{T�|�i\x�O{`��
A�;��ǵ����Ξ\����XT�;O��g�v�s1�\$��u�N�ea�ّ�ǹM�ʘZ͝p�!�1k�_ڴέ΄��C:����u`dJwj7�<�,��۩�k8X��AcH�0r|8�"��<�}}�X,D�*�,1��u���D�����ڏ�'���M�k�Ź�^������-�"�*�:�m�2�uiDՙ�i
O�Ե��i	�@��2��k�Þ.t~���h��y24��:��P�<ڢ3�v=���ud��U�z�ϛ��&�n��S]e�v����E��KF�Bo�9�V-d-&
CP�#����a�4WF��=��M��l'�<i@ٜ��	���p%������z3ʃYWY���`ײ��������(z��~ɸ{2�!G��EKv�d�>��*��]�]�Ѽ��8��%�w@��kƬEH*��:���.���ɊWl�ӄ0a��8�x\:�w�5%q������ڻ�)�-��M�&�Ԡ����wm�A�lx�d�6r��Ua�z�A|�,��Gdպ�]S�Y�0x	n�6q�$�3�]�P�ʝ�W��?	/�W+����}GoXa�Z�1� 7�L����er�V��Ƭ�ֲm�n�2N����ݵ|�}��uy�H!~���廷a�/GV޵�^�/ד}=^����<z�Ղ9�6_t����XaN;���1;�۴9(ݜuS�A�^�);�A���?�;{N��[X��ҳ2�̓ ���r.��-B�7,R�,�I���($�ɱ������r�Ә��p0+�I�W\����϶r�;�P"�vf�p}w�h[�	��VB��)=+gv*��L�BXm�Ч��F`�w�ھ�����V��ɹ�^#���W	mA�=�ut];\^Ъ��.up�Uξ	�F���1m��6��l�A��S�j���_}�g#ʢ�/i)\E����7#�a�]*��^�ŬA/�%�m-9M�¦[l�4�t����I#�[z��\\�lݸ)�{�gi�/��|�xI���
X�'x��}�Cl2ӻRdc)�uaL�+�[Y��l�2�Q(v+u��߯z��5�-����7r�gy��k�[>4���v��\`����z�jE���e�\�\&[����r
�'�J�þ5��=U[H��I@-��ti�)([{�t���r�F�vC���;�ǥ���:����% ��;'����,�=�-��8E�}7-I׬᳚�J(h?���%B�1���}�-X�o��p�Wִ���l�|�cW�,�M-/:Bo���z`Je>=�5���N��1�n^�&�����i��#b�F�Ӿ׳M�� ���滂����vig��d
:J��"�m@�:#�r��3�b;p!C��Q5��*h�q�q�>
��Z*�`4N��$�cR�֊��-�V��i����y�'x6�p=����e���?f��M���좀s�-Rk	|d�TKH� S����H��vԥ$ݑ�Zf�r�:N�fcH�L�b�Bk��l��b�s�]�V����lw���kڽ�u�Y/i�jS3��|e��s�ZR�7p1[�Qz�2�w�f ���4B'`���EKݧ�f�}J-`wr� \[�0���<K�Î�L��|y��c�y�ⴃ����jm��}�����I��dDG6�;۹O�ۛ��5zn�&P�eA�zq�_��=�U��l
���p[c�h��0���!��Y�+KD.���rʉg�%<��)R4��:�w1�i��ne |�����ZS$�SV(�@6���/&P�|u�<��U�OFE=��Nw���� �j�^���{��m��ҙ���EE��^�K۷�0���3�v��-���@SՄ��v�� ��{���]�w;i�CS����B����Z ���"���]Nh�^�g������տP�WCg�*����Q�oZ����.�l}V/U�5��J�����I�nwʛ�OPb��{�6�6Z��t�"��Ό�y�-K�:"���3szqs��wK���7Fv��!�إ����E�f�U�9Tޚ������6i^��k �e��7\S�zsy�3�xܧ��l]�w:��`&;{G,E�upofP�ǔ�V,ha���f���ϡ��9�a��ë{N炮˷�mmsj��p=E���1��c(�i�{�$�:P�I�ŏ ��W2���7m�F�ݥXNz�2ge�Tn_�c����r�p%�4��A^�l!��8�㖿���N�:���d�+�ca��j���#ȵ�5��8��o�gw(W �Q9�y:�ݳ� �������,��_(A�O�e�#j�e��`�_���"^�?5=���:oNʴ�4��|d<�Ei��=��ݧZf�t��ܷ����o��u���VCX'��g3|�V��6��h쮊�ʝ㾁ٟ#۴q6o+2�6{�9v���c c�#�P���T�Mm���$�[kZ�f��u�a�C|��_3Aq�77�1���}�Kb�m��D�4p;y|���á���Ի-`<sy�/nȿ��1t����#`���f�l�̖����h�d0�8�0�8b`麳�E�f��>�[!c�Xh�ӵ2l�����ֻ1�|�����a�	��w���X����;2\U����Zz��@kUe�&�I��3��8����i� ^ޗ)��U9{��Vή�~a�^\�t�b���u����A�Ӌ�=�3v8A��ʋ΃�i�+v:���)�{�R�Gf��v��d}+q��%pf�X��u�v8{�BH��l� E�۹�n����Y��ڛt���ˡ��k9ǆ�m��U��c��mp�������(\TD)y[�A]ʱ�*C{�QR��k��Lc�<;�/|:b�I_5��#6�`�z{��zggb�d������Nև=�������uÓ�U���swkN�W�
����r�~-}�+:|,�V�г�oo\���]9	oII��ĺ�M�g�8���v_e�_A{�.���I��`9�H��4�h�i�D���¶�C����Ŏ�j��6	�����CH�ua5i����aa�� �_S�XPW$���v�:�I�VT�;�H:����>Y�3MY��tRT�룂-��ޔhG����_I�܃�.���4|i^�v%�ìލI��� �5�+/��=����N,��Xs��%��̤�QV�t.�3ƛ�.�雱k&�f��M��t_v�	,j��W'��(4�l�L�' ��Qcs*ƅ���<@��6�4yfiy�G%�t��S�N�J8����p[XЦ2����eе�����J��ֽ��S�d���[x���<�p�%�5�UQ�Q��p��JFTF9��x��2�����VH�}��&�Qm��r���g����7�2�)�	����-���]֥8(� ��e[�i7ɑ[�,#w��y�gZ4�{J]@��C�x�ʛ�� $���,>�I��4����)����=h��n4⻻��ٮ2�{���mCA7�1;�Θ�w�V�6$Z*��8ŭ��s1��+y>c��ư�jNRˮ�n:v�6E�(���j�t&Ĳy^'����hb*����
���{7M�Xeվ|�>dӃPBV C��³h�7U/�˓ܯ�^|���+!��,�n���z'w�U"j�z�-�`�9�� ��ڞ����*�����$6�D7����H�{,���� ���`�|�f���9�z��u{�4h&�t�&œŹ�+[�nj��IK��]X��Q�_\���Rq܆n�i*"�-ގ�.wm� iqwHWTy�p��BⱁuFٮ{�糖�s*���
�[ϖSBӨMH�4fǑ�t���N�ô����X���hQގ�e5g���	��̩�ԫ�C���=�)4hR�@�`�e��憠�V����}}�ֻ߄�YH��8q�0��n;y�]x�}�d�.��(wcgeJU�<ލQ̮P��m�eAٺ�7�_xOm��m���_�ήF֜�^��^�!������fiA �{k9fh��+������w��� �M-׺�X*�5/�s�m:��Jݓ��ݰe%�@Wޝ����1��u�-���Ù���;HK�0�^��'H������Lf<������whWVw4����+��Sz�ަ��Ys5���ɻwƅ$����z�������r�θ�pk0�L�P�9JN�>Ӻh�tz�a���7<4��+[��Fe�P�F'INܞT�������,���Ĉf�{�"@�io@M
4͌�9n��6!��"&4�u�=���Z�<�ur
��� .�x�`��b�g��9�M�s�����`�3Ep�v�}e����\Sl�;���N*�չZ���������{;��i�޿�Vl<>:��l�w��w���9S#�_'8�H1�u�I��#�S�ș�9�hZ�ݣ��ק�o{s �}u�6���$�mׄc:g	�d�Gu6{���E��|D��=c�P⊤qǱ�����LSn��j�n�+,�7�������?U���xmI��S<؂���9e��}��N�cΧ�A�zѠ�K��l�s�ݪ��bze�Q��)Y/��n$������,�g6ן��Q�p�:�n�I}�R�
�AK�E��N(�O����pҡ��;��U7j�K4���P�p�5�+���]�+
��Ɩ��6�ы%�g{u;
��Wx�g�@���-^% �a^S����2�8�+_.�{X��|����dLK�ӷZՄ8�ns��L�F��� �%��Vn��ηc������r/C�ϻ��Ե�gA ����[]�%C%��(22��J7t"�!5&X&����2'�z>�P�͙S�SK�����Tk���U�rJ��SI粥_]�nX���(���f�/��/�3m��zD�<�Z��v�*I�k��J�(��կ]*v�<�_���meY����.e��U�#�u������Iܬ4�
�s㡬�!-��k�ݟs��L:Ͷ�oM�0y��zˀ�?U>�=����0c���`8�:�Me�V��i]�t���G�W�0K+yc�;�Y�Ҹ(�5Ӹ�WZ@�Or��5��M�[��ZB�Ht!'M�A������R�0�G���1+`Q;G��L�M�r��s������Ӛme��a%��������ݵ}�CO��^�`V�Ο��Ƿ�{��{pV0�7��g��R�m�-�ڛ�QyC��P�+��0K˸� � �p�I7�{ĺM���(��\�ǫW��t�z�2��D��	,��ȝےi�×7䖬��	=����n1ω��x~ޠ7Zo�����G6r�U�I
��{�+�";��B��$PAm��/s&�2�j\��K+��U�;!%�̫�q�T���R�ej�Zx�BR�g�q:xQk;����.���1�;��r4�٤�q!�%���#�I)��������mOM��H���
�V:�ԯ#���Ȅ�vVu��N_ks���^$�.���8e�l;��:��YWe,g��˄ ���E�cmæ`2�l�
��;'�i^��m��������;�%��)9�UE�R��l=v�k�$��㹅Qeq�e�F�๜���'n��5�V��zf5n��y��Y�P��oR.��$s��Y%��ܬ8�n�E��y�%�v��cF9��p��[Y�����9�f�)}}zy��[P�+����2�p���E���׃��Gv�^��_r�_x{�����������}��_F~g�*<�M]Y�Ъ��_F�-4RW��k
��0�Vn3YE;�w��_t��k,_\	���5^�U٢n����N��B:v��N��p�θ�o���N�l�%IY�U���]JKyic�gm������$r9�!E�B�S'��y�i�yktշE*	aTwǰ�4�(�+z��P���!WP��5:�*-��f���3w�!��V�L�,��V�v�A����\�n�����)�Wk���N�B�ˮ�0�Q�65�i���\��a��V�3�`繰) ���k�%�b�X�q��+eI�5M��Mm橊�v-��J�i8���T�s[�՗��K2����Q�כ;~�z���{p����\�_9ݎj�	�\,ZC7W���_U�����P"����K���u��Q�@z5Չ�+ 侼1���Uq��iqYaT��5�ŝ�%�a��V[�s/Jz����2�yp?w�z�; �������˴Sm剙���v4�͒<=�i-!(<n�"�޵��燡�lpSy)�����s5P���^ۃ��Ê�rE,O�>����]�E`�NC����֗+��@Қm�v��
E�tf}����m����c����UtN�»E��
���($�gk����i�̮������iݮ�K˜���H]h㹸�#�Y�Ahi�ݣ��7�����^o[ڼ0*V��y.��Ȉ�Nr�(�$z�,"�v`�ڴl_R��H%��/9�奲����|��wc��������F�:a�B"lV�^qCP�v32��|[)���.���u'Xl�H����u2�>���P��9�y����[7�n��G�P����n�ߥ:A�N���t8�J��
tw1���81Z2t�q*E|�c��'��w:ʫ*��tD�����yٗ���kB���� {��'��^5�BVcʺ����o��D�YҏoL��ݴ�W��n�u��ޓo��e��T�	��P�?"�n
�|�@-&�ٮ�֩�Yvu�p�7�:56�,�]�U�f�E"I�]���B�.�g5���:����6�=h�L�1�Q�Dd��:J�a��o�9�m�]�H����k��7���n����f�E�T�XFT�%�9��~�x/�y
��Ӣ�VW+�=�f�eJya��lԦK�f�7A��׼K�%	[��9ʙ�+���.�<��n�ӚF����^H��)\�\�F{�xd=�R�ֵV[u%�V0�����n�t(*��x���[��J���!\W*�΢�l�T�E�U��o�g.�xh㻷u�G\;���b��-�]�4�}�|#���߬�i�R,s�6��[�*��XLCL��hز"�r+bƪ��nԿ���������R���a�SVr��`�j�<��#���i_\9W�[O(5�8�R	/� �w�QH���<��"�c��ɜh������}��B^�(
DRK1�HSz7��Gb��n�؊��6��H�U�|.�e���9"��v{���VU�V�WG�#�Dl}5l:cA+�ӻ<���L5y�CJ�z�;n�jFC������t2���s��g ��+�k��L!i�-`EV���b=��%8��S6q�V�s%V�RR��=ξkk�XU�y��!2��3)��e�Of����Y�w�OI�����0���tM�Ԭu�c��ڊ}�i����Мz��6@f�oCAR�	h���f�u�'s��Vs���N��N��$k]�SN6�yX�0R0��Jl �i�V-3V�`�,����k�>s=��V�^��=r���l�����Y�N;\q74G}��e�V�h���ky� esJ�է��;x�w{d�q����t�w;�&����50��T��-z*��8�-��5g)TP�gIFM�v{&F����?�)��x�LQ�{p�v�!������m�ӏ2�'�ٔ|gv�7jQ�K�X9jʹ��RZ��r6U�M�
�M�C:�pZ��U���<��6� �)�~�S�jR���,	w����z/6
�\@'-�������nf���5*u_'Wve!݄E��{�ȠS��~Y�۴v��{�j4�S�h�=L?]K���&�h��txL��;ɢ�j�̚n�=����ˆ��$���d,���'fL7��N���ͥxf�i(��dɷw�����ou�rx�A�>����1Y[|ٖ_c����xr�d�}31�{J�j q�nR�r^|��S��{C�ZMOt�׶80V&�@���qۭPu���N�u1k��veF�8�'e#U�Ӧ��݈rړ ׮Q�ݾ�2ܵ����/9�C��~���q�-�:�\�8t�ٮ�@�k�9è�����#R�i l�Eg(��]t���i��i+>Ef�8o=�g����w���E���.y���S�fU�ԣo��fVd�a\2u��99Ljb�'O.n͉\XJRH���rz�x3��W�J��s���̖��<%^�o�,�ċD��\s4w,.��@�؁��j���ܴ�����٩Q����j־�U�3��%�����F�μŵt�?�n�m<A��(s�\���[�iS8ҽ��Q�C�z���b�2�1^E�x�o&/��3#� ���I�q��T�lj,S�bÍw��{e9 (�ڝ�;��hCYd���D�lc�7�Co]� [[��wD'jz.�]�ݫ���M��!�*VA}Ϟ	�b1�k�n���ʬ��Uȶ6��
׋n�$�,T.�ҹi�Ie��=���f��e�dTSu��M�b�cu�er�0A�I�Ry{�
M��Y���'�p{:�]�T/�\�Wj���	uw���v��M.���z�s)�3
墐���S5O<w������#N�﷉�n2n�v��~��4o���7��{&ݠ����F��qf9���.���El������Z`9���}�A�M�^U��W�rJ�M�]��O:&V�,>[k�Q�Yw8l�[{4��d@��t��l����tS)SB�-�J��Y���xr����)ou;�ӨuvI�kh������n�v���9_QX!-꼓�.Z��NK9\�%�������m�o6b��n�(�K��^h�.�Dr�D��œ׶]�!z��*Θ�iԈ�>i����=͋j�u��3J��U��=��F����og[��;Nvv�C9�)�W������i���F�i۶�b/�X�t�Y�b8GQ���yPa��v�Yv��ڻ&��G}�ʻ��u�%��Sk> �}��ul�ԑ�܇�%9��� ���x�Jx@�v�6��U]�C�h����Y�:`�j�vm��e L�Z7�Vkp�b=P�7�駃HL���e�A�3;�d�!l�c��-��ZZ5��K' A����wV�g���	����Y��2�7Qq�X"��^57��ú��Z�n��Hɯ�/�O^�M��jb�z[<�۬�Gq'�*��b��n-�p����;�/@�4#ɥt�,�rڡk�*y�ts��.�ގ63���0
���E�<��׺��38�f�O��H 9��(���A����m�<o+�����x��pa�R�n�q�a��t��f���Q�%d�2C��x��z�4�	tSo'֫�=;�,r7�Ǉ�*��\B�(f�o"��@^{4���c�0=-��99��:T:Q�[� ]O.�H���+�:�im�
�k�Lۧ��bf��V���Tx[�ʳ�z�8U�Q�)��[cz�-1M5�W7�=�!�H>Z;�/fZ�[|�Г4�u-�v0��jqfU�ms(1�:�c�|h���PY�ٶ�I�`��;�*�m�N��zR�&����]}Ѝ�O/	�_nz�������P��7�����A���i9�a�D�X��jX���\��n_A1����{k�y�.�0BX"����S\���i���zFҔ�l\͵ה�6w�D�����8b��/P��`��_���G}��aČ��K��d��c�CѢ��W*��T��"6:Z/�B���mS+�nO������qFۄk��_5����Y)|�,ʵ��sY]o(p���Ġyf�Ŗ�!��{9��9)��2k�Y�r�wk8��
D����^ɜ8wo�j������^��;�]�0�N`�問3�LV�Rr�ƙɡ���_*�f�Rq�,sK,_-}uyZJ�e��ө� �st�)yA�!K��6λ��r�V�KQ٢b�k.�,�x���m��e�U]խ5��NK�/���|���k�C[�˝ε0'\_�;/n��d��M�� -8Ժ�:c���[G����B��]��L��k};f�&l)��M�Xs�Zp ��lB�u��P�ݽ���a�Œ��_;��%Wڰ�7dA��;��{�Ș� ]ʱw�agۇT���o�PwkA���򛵚s/ܭZ�]�#[u�9>��e@�4�֤׼�s, ����}|p�ך3��^�^ԃ.�7KP᷽�4��R��Ð���e�0�ݹ�+L�'jщ`��xu��4B���\�'�Z �d��Ol�^8(�c���4���~y��
�R۱;Qӌ�ٶ)PX��e���iʴjЫMI�L*��<%����u��X\6]�y�ێ���g*g2{�M}�ފ��>����#Y�,Ւg%ӈ�'_n�z��\뷡�U�M�/nV����#D7H�G<s�ۆ�}W5�Gal=B���2yt3����׫ h�x�"ձ��H\�-�׮j5��랦�����Q׈�i������ulˇ�.L��ʛ��h���Ҵ � n��u���l=Yl��͡���K+�w�x��6����統3�fڎ���j���Y������5�mwY��
����:\������<��h��q�-��W��b�b��ݧ�	�5�j��'�b����h���`���2vr���1����{��G�Ĭ��e�����do#q-'..��'3����jҊyP�}11�]����*W�6�'�Ō}�є즵��b
�����85tY��=���]�釕�fΠ�Mހ��><:�U�Wcu}i�v��{j��Ո��o�����S�JNH����,�!��u��������s��|���s�WP.�	� �	���C[}x⍋aq�9Q�Y��8�Z�Ofs�.� ��~��D��g�v�����K�b nե�,�_Ū�kB*(q�fu3�8���H&fֲ)bw�K�o,Z���d҆88��bCNn*���f�����b��)��&:�2�í!X��璹�B��.'�B%E�[�/؃v�Ŷ<�����`:u��-ij��H.�C��Hԫ�!tDM�� ǎ�s��.�b�uh�c�>��>�`ۺ�]yB�sዢ7;X�U�Jzv����e��*\��(�RIA���yv0�ĝچ��W��j�/\�
+�D��8�S�.�x�:XZ��y�ZY�t�..��qvH�=�[�k|�����O}�c*�[T)�u�mռ讌�@N�YrYK���&�&7��1��uܨ�;�>�:r\���	�>���N*f�u�n.-��6���f�s�����5(���[�p�:��e����9��ݭi%���Q}�0�R��ժ�m�ԟv�y�}�۸ȥ�{�JN�h=}}Y�*6���|����쑖��^��J�ԕ�c%	X�p�T�rD�*��"/�Rsft�{�h�N��=�+%`�b32�;.D(Xե7��P���xS��/��ڻ�\N�Z���.�OI�u̳���)r9N�;�B�I�\Ug{u,��{��r�� �o4^v���Ҧ��k��'�c���i���gJj���]�S��%���H�� �l̷�0�3�T���C�]���"iX��OxZ��,d��/1�[��wBM��N�4���]t���1�$�ի�w��k0�;�VuoYLt��l2]gB\���V��sW)\�M��tx[l�T2��³�\����]ۜ�z�Fs���[�G'ƕ�#���m��JZ2�차c�}��H��:�z��Aq�������mXnbr�-:�٤�=Z1��C��N8L�e��,.+s�z	Rѝn�2���v+���Q٢�q̈́����NQŗ����g�u��D�K�啵C�Zv�<�)����g{7q%��|B�/|-邋��ڇ�RjpjB��ʆR��(�[O t�YWV��=ֲ���젟_A[pQϢf�F��6c�׉`�9�kN�3��G�֧�hؾ����`���!4��=��6[��i~���p��˦�B��l�3��&�e�K��&`@nkS:��~d�IǬh��V�[�4ͱ����je]�t"�h�!��z�r?WA<<�uX�0��m������9_"�F��v��M��	tʱ�P�.��*@J���Z56FuMP�Cq�ΈZK��@�܏:#���zB�T�8���4�]]z�h�w2����&d���*��ǵ�m�9v�m7
զiK�[�گ�ݱ[�֚��9p�p(57Ď��k�ԩBӸ)k�Y�`��T��\�׮�&��quL��\jcx|�ãm!��>��_3Kb;(x�"����[��� ����\�V�t�Ri�*U���{��Y��U:!Q�҆=��Q%h,���������
��d�;D�;�ڳx� `�zlVmf�D�=B�O�	R�!_+nneڬ�q�L�!9�[�U�Rع���c]v�C�������+�Jq�r�e��Uv����Օ/Y$�?aR�uT+� < �������zT�BCe
��=hm�����:���}J^#[M*�w�b]3�ݕ+gW0�S�A�I�7�5�e� .�[���v:�h��T��Lf��4�L�n����2�u9�����b�Zݨ�N&$��a�zP{���g2�/f_ow�S�IN�$_m�|�i���J�4=��e#�f�)F�T�N�*��km�3ۋ�D!W�P���WQ�|J]��iu�۠� ����{��t�:ѩ̋���뀽��	�A�V{=���Ɔ��g�#���!B�3}�Zv��/���܈6�)�/NF���,eAݻF9L�jX��UX ��b7��,8؊	�Fo��/��{`����|���,�UaS8����Fj���=nb���e�r��cj��J�j�R֜�8_Z��'��Y�\�p�u���`�<R,SR�)������v����ڤ��p��)��&��n��#a�xz�r�%qQ:5�|�K��+Z:i��o�S>��k"+�^S�T1�s�Έ�:�;h�7c/��㹺ƪʙ.�)��g�]3/�I픅�j��I�����۠������L�j���B��q�BtŌ�U- �bM�@	AI�ftk_d�����3�ɬnK)کd+܃�N]�W���O�#��VC4�{�f��qg[8l\}Gx�w�]�	2��3�0`ġM30�0I�$61FɢC$�����	�i2A%���)�1""LFdE"a�BDw]��w;]�Ɣ�2�'8�P�%��h� `�r#�u� k)�������c&ņ��1�	$Ě��d�L�JLnU�#b�s�dfȍݹb��Y��!���!�2��S�f���;��TE3&ęݮA.�A;�	)���(n됚Y�wk���Fs���9J��CJ1BX&6fwqhɍˤ�b+��@��0��@��J(a	��̋���5����Wu��,�:��E&���H�I"51�۳wv��2Ar�2Ph���1!,RH�ȉ�f�c��fI�$6Wu�X��ӺBJ�ؔ�>0}�g�{�>�
.'�l�z<��wl�{I4�ʉ���h��-6	b.H;]��L�D���S"jU����"��f�p�J�1W�Bsy��U_��t�@����J�c�(W��V�{����!�'8m{�xl�Ա�i��,\�����?���v6��O���:A�)^��Lt@�ޛ^�o�޸��Q�WOmߴ6��y�f���VC��\vFO��qx:�q<PE"�a������KgH������^̯!V6+��S�z����"�٠4�FQ�T-X���X�S��^�%Ǉ�#�I�ͧ[�`q��;�S9�R����|�J�ma�h����2m��Z���-���VP���B���y��Y� �oN:Zw�N���׷Kw=�[9�W�3�&�ny����׈QC�t��+�8+�ƅj���q���LP�)���z�q'9�[�![y�!�^���ޑn[�s��4$�4eW��<4� Ď�V{�����mtì���O/��v��E�T�s�et+t�!�NЙQ�}A_�eP��Q�XE;���tZ篪��Q,�o�r�e����6�PQ�y)��=@�<i�]ˍV��O��yi��:�4Jz�Puu+A���2vZ��";IAZF�a��>�Yˈ���(K�7��<hv�ٚ�~>BrF��~�|U/pP�үJ��kx�i嫭g�V�ؤkd��k}�^��Z4)L�`�)��;&*ĉ��ՍE�'$�7E��pUF���uIV��E�ё�.+�ƞ�d��T�
�"��@p1ӕ�R�L�x���lC�9ٍr�1/�l��\�����N�:j��;�Q�����h0to���kQ����ߴ��ߨ�*|ȡ1��ҥ�z������t�ף�}���q.VAڛ:(�?~ys?�Z���x��J�����D]�̡�m�fϼv�us�ב����.e��_�rf)�����k�=C�s|�S���;ŝ_/�c��5�8��]�""�ۻP�CT��R�s%y��Ba�L�)����5Q��0�#�#�G%@�.
���kQ�᳻��r�R����ԇ�u]�����MnP���Q�x0������r�d[��ҕ-�����yo5�2FB`��E{�V�/v\;;G!��v�*U��|(��}kOf�B��W�P�4��Y��J��*��Jj�M,���j"(n:,#,��O����vm�7��НY˨{�/�w,��	̅V�t{��EVK�N�"87���:��q<Ȫ�v6i���;�XzkG�tc���;t��y����
Μ����5y}FL�CBƳ@#;��O8�h��kE��y�{�������AHa8{������ͳx� �J���j�v�]/:�\�$;¥�d;��-{hd�ҥ缳�z>�=��O��Z4��:.%�A�[o��Z@h�ٖ!J��ׂ��/�5��� �)��G^G�\>�t���P�Ma:<�%��4����/]�\�
��GG�qZ��T7����TB+������ק���E8�q��f,9ո�&��S�]�-�F�`(bgiE��:S�d���N�z��J3q�y5a�x)�g�"�(軠�ёؔƆ�����$��bD�"�ZV����K��e4Fk���\t7H���m7qW�U%8���p�'���&B �ZM�̬�B�tW�>�%��|wΓ�1��;��ͯk�济'ո�gY�O�H�z@�D�ҭ�pV���Ƃފ�N5�t/|2_u�(n��/�N@L�yY6�^pQ|�<�{T�h;�E:�{�k�ٙ���]``�MپTc�[PFP���ߓ��Ysl���DR�D�f����o�v#�bs=�$������KUpC�4u�w��f�2=�#\�Ѣ��X����5�݋<��Vx3��2K5��-�fiM���u�/L��Br��Q�7'BB�/�y�{�h�{�MDu��K�=�8V�R�=�x�ˍS	��'�������fH_t5&ۣͮ�/��Ajn~낫^���ٞ�i����tG1b{�5뽛�2�����ٝ��c˗�o=5�ub|�z�f�]�E���,\C��ܸ�hs�+�S��z�t�K�V]�r~-谝b�?^6>��HMu�$>�g�5Y�����j���!�ƛ��&{b9n�^��L?�ƅ;<M�`�Tst��������3�ɞ>���m�2����3	�a�%��JG��쾎$j��uCЪ?���N��>���'�*A��B��'�:��Uzgd��4��N���y�^��[��Dds&��Q��	}�|�T-�E���G�kݜ2��M#T�*R��g��#6ӷ�;�]HGv��KW�a�����I���W旅�z�C��}>�r�&R:�w]���i#EǓ�%nn*��&�D@r�3����q�E�J�T�Kw��ćx�!l��q�u3<�3y����w��Z��p��FG���e#���Y����*xmc�j�����M��7ypW{�{w�1u�n��D�����0���v���}<%MM?7xY^y4�r�f:�nE�1�tM�y���Lx�(N�dfD�8;ç��adc�,mo2�-R�SK޲�OV��\�78�sz���0���N�T5���F�������k٩V�ta�1Mֳ�3�t�;�h]�,�Z�ӛ��Dr��sO`F�Q;��Rv�	�@ڶ��X�V�߹ Em�m =]����Z>�QɎz_l��\���!�eoOF��;l�&��Y"�hM�;n�٨��J4�LX�E���s�{��m8W}�ه&����8����=�]N"ڲ�-��T���l��ol�;��@���4ǂUyGa�G�uL��N�_NބxO��P�2^e�k���׻��n.Vv��f;�#ޓ�j�Շ	�@��a��iun��d�PP7��m�y�WE+�N�Q}8Da�����ݛ׏j�B���Q^"�������W���?vF����S��Z:����������9���m��L�ޗ�b0�(a����ٜ��7.:�d�W��8��g�o�s�<andJV�X˚D�cz[63�_�L��_��\��T���hE����C9�2�;�u��DU��HC���u=G�2ou(��`q��;��s��	U�w*�B�ʝ8T<t"^\����W""u�Ux/�v��vc\��k��ρ���K��ه�KPv�ߡ5sG�/5��F�����n^�m�	`��K���͚FK�<����)�2����<ɨWuN�xUm��s�Nɔ$��u�c6;� ����i�Ѿ�m�u$�O6�u��y���]m-�E.�/Y��*��]��V+��l��!��Q:Ye��{;�c��ҽq ����x׫UD%�3{d�c���b�ٽң\T���Cu�����z�t�s��m�2E��-�uEs���|hiAF����pd�J ��r�V�9�m��8yc�Ȱ*q�+&��ɮ	9ip
���"x��/,�y8b{f�M=��d�����Q4�����/NG�1�}aE�3l��F�#�7홆�Q�4�=�t����������۪H�_HH豽��J�#�o%G���
J.m�;��ffouo ���C�P�Ej��i!����:���Kj�p�eF瓮�lcv�ݝ�viu����[#?ABWCu�'�ʺ��#a��:�V��FG&�B�/��W{"dsrǻ���F��_��]�v+H��[N��+�Ս��\��otvPQbc32��Eⶪ.�b>��|�y��P� U\��T� D&sǧ�V�EIL���nڑ���kr�Z���/�˯�ڡ0��MM�G<���"�8HG��J�^�t�]���w)��'�.Ys��pWV���B��V�^�:�4\��G���� �S���¶��
�TQ�x�`_k�Y��q�F�$p�T�M����V�GݠөyQ�y�vR��Cu����ͭ��'A����F���Wp�pNކ�IL���Sm���OU@ˌt�|��[�͐�����uZC}>rhr�n�����8zG��a͔�]���B�"FC���gZ�$_�eC�����S�:�E��}^�y�i�ܚ�/4���E�:N�� ���!�AG ��Q��8PY�,s��>��G��嬝<|�K�{�ߖ�e��/�
������EV$����#�
�N�-N���>^�oF��}l\�K)�/gںl6��_�����"a��d�:��2���@h�e�h[��7��:���x�Ԧ_k���n�Vg����IOC���U!���|�{�X�8{�Ot�!���*�D"��r�X���Q|Tt���0t:�T�l�U�d��*0=�6+����^|��S^��ǯ�å��#�j��f�6�X���:������^HRfm��*����ʻL��t}:u�b|�xX��~�J��Љ��/Y���usv5Cٞf9u�9��D{{�"AJ���+g��y�g��5/��������b�Ƅ�K�P�X���((u+���Y�z��>�]����Ԕ�Db�\t������BGU���,FƋ��r+�br�x����v)�<	�dq�V�u�ǤE��byX��ԅ�V�}�@�:�t�;�E"�FL{�w��/\w��\��{��I��@[>g�u\��w|+���vX�<����<L!��S�]:p��>ٷg./�5Rf���}n��y�T���'�֏j��A3�7u�3���찟�F��9�n7����[���.m��Ȋ
m�:k�ds���D4���E+&�jrfUAD(�q���Ε���l�L���vh�r��*4�2L��GF4n�7.L�u�;��i2�>ꂬ���2,K�����U�wuqe��	�姆����[k1�U�r4��q�U�f�˕ٛ
�����>�xJ���(w�W�h��K�.s�_�2��m�˘�q�=Z�B��x�`��3�땯qD�nU)�Ꮵ��ڱ���8N���{�/	����]	��΋y ���Td3����ƥ�^���WRd�%�l+�t���'��E�VyT�e���㲽�l�<�8j��|���R\}���;�yYy3#�iK~G�w���3�5�=���:}��g���[�:�q���"��7,�ND�E�cs�V	�j�V|s�ͺ�[�u99��b�uj�]W#A�ۤEҡ��h�Ȳ<Z�r�R�F�ε���|/�ٕ�������4�CŃn��kt���vyܜgމC*ជ�g#������ ��KP㸟2�opGU�+�� �^V�B��X#�a�*�^�g1ǳ�f����~��aҁ~N[=���00BNl©D6��ܝ���\����(Р+.��������>���]�}��?VW�5}%�^v��Mߎ� �����`K��B�EF�R3�a�
��G���lE-�.�Ic^�aX���$��jw/x�r�dm�u����c[���O>@����:�s:W��C(\'9�=��b콶�U̸�6
�㴦bp���X�V��`���ƞ�3�D�O/�%���2f׊k��o��X��Ƃޮ���N�#	�-s# &�uT�B
d�gd��2��1ج,��\E/D/���axׄ��:r����amYg"�*��^#V�}=[�N깱
���fT�		�Oa6������P�*0�C�sR�j�����e��;�8��y��+��Dk�/�'k�f�yB���ӂ�q�C2^�{n1DGۻ�zj�aNۨ���,G3��n\F���FYx}���|����鱌t�J,J
�CMe#s��V�W��w�.�E_��ĭ�BQ��'*xy���2�9����J�v+%SO��<���6�?k.�nX�[�+sjn��*���s������K��b���ե�B�=��������D/E2]�K��X%�k��c��Nx�Nzãmt���,t�]�G��o���_�����D�r�FO�e$=x�Z@cJs� yo��hr��T;�ҙ��j�aL��_6+�\����4�iD��-O`B�>�p-S8;���V�5�V��Mϯ_���S�7�7�U�vr�DuF�~�E�^o�����>�ez��8_�'f5�	f�Szp"k�z�U��;�L*B�*˕�V$��</r~�7�(~�7�!�Ot���UD�J�@v����l���~�[�ѽ���R�R'��[�P�v_���~��-��0�f�eW��`!���@ш�^�7{6�ժ��acO�<�1�l��8���8H��$�	�HZ����7~�Kon�W.,�l���������<�2��i�o�(�3l�n
41��V���o	-�u�_[�,J��
T�۟X�l�v��E�ё|��G|9�i��q�.����I����t ��@u
� �j��p�����Fz[V����q1�=�i:��ݐY�@H�v�^��ʰ�3s���@���P�f�WI�M�b��Ɂ�F�M�;���Ұ?D����(�k8@��L�{I�LZ�ьP�0���=}x������x�Y7��\�c� E\����)'���wNL��������$�������8��i�if�j���VW5�f����ow2��W�x��c�(c�����9���e��_S���*�V�.���S)[;W��<��n���H��u;��
a��R7�ἐש�W.!G;|�y>쾝I�OL�w9*���﬇�ǜd��`�=�:#:=Qu�Yל7p��=}b;�q��3,�� ��X'D���{��i݋����w=�ໆ+³�/�e���k���V*6#]p l8ν�w�R�0������'�&㓻n��Q�wxt���q��'��"W?�Z	��y�'V��Y[KV[�Tǩ8��n'�h$FP�������s�~k.Y;`>;O��*V�8��썖ԬL��E1��� b�I-S�3^m�B�К��l�Vx-8�w7ӱ�O#��(�0��K<���sKU��̔r�[Z�ˌWv�G%�l'�+�[��2��T�����.�a�z^�X~Kyvj��Y���*�`M��\�?<���w�2�i�e��6; �u���ӎڌ��
�tt,�j�⸽g�p�%����>fh�p-�9`��<
HTЭ�b"1rpW�Zޙ;�}2�2k/@����VTZ�Պ�[��mL�2;�儰=�Ҳj㮬C���ێRN�0�65�5���L�	qs���:�tT�g�Z��lM|����h��1U��N��[[+�\�U���wn�|�ά�{"�]Q����MW$&���ޮ�[�{H[�H�I^�fp�v񝜄t���+jv]��k>`kK.$1�;����F�_��垻<�z���{�Ǔ����=��;���+^�$�)M�7��*�=��P�=�X�!+�򜵎Ǣ[�شe����6��6�[w�I���1㷶g\�7�78��X���������9W`�b7�ByԧB�`��O��W^`�$���_Pz*��	]�?�|�S�R݉Y6��+�;Y�O�Pv�U����0�|sZ�ҭ7�������tەLa{s$�WqF��E83��z�hOL�Wn痼_���A
����#H���p����3����f�������u�y�k���5�	�"E$�>���TI��/t]��k�'��WZ�9����o�h�+�z�r�X���u�����~]���.w/���a9y��4'Y&x��x�J"����+xֹ����:��p�X�51�^�`⁌#�Eη����F�M���v���=Cr�:Ǚ4����+������y�J&=\-� W�9kqI��#} �63itZ�w+�'��A�%�$&Q�F�FK�$M��%JTI�b���a4�#(P�wt�DnZ�)��fQc	����9r&jI$�0А���"Gu�k�FѲAQ�$��i#!0��Ah�%DcD̂I��\�H@3,hb%)+E�nW�#����E&r�B�F��BD��'9�#3%�HX
��AD�	b�4j,Hf��")d�,Qd�	@)�hуr�d���"$(�$���I)9qBd��f�Aw\3��`�s��b���Wur5s� (�b������6�H��wn(BL�%;��%#	1ns$�1.둀�0 > �>����lK�<O\5��ύ�6Hga9h)�'����^v�ݒ�"�*����_4,��0���;Do�6#�����h��m�Ѽk��ӵ��^-�/�׈�_�޷�W�����E������������& �dzb t{��=�*�ξ6���ṷ*�\���|���r�����YQ��o�����,^�?�x������~+�x�����^��ۻ��~>�kF��ם��o��������ϝ^9�y�Z��ׯ�_潯�{^-���x��^/�������T͇��MO
�ղ�%YJ�-����_o���V>�M�m���ϫ�6�;}[��{[깹����|�[�\��|����sx�ݽ/ž==4im�|_W��y��^��^��������d �O��N~W���Zj�標�Jc���=0@c�'>�� Q�?�|��{Z}���z[ҹ����篝o��x������;�ms\��_���-�oj�~�������x�[��x���6�U �G�0 p�/~�})�S�}�R���鹽6忟}������O��[����p���Dy���ǂe{`d�6�wϟ}_�~?������׭���Ҽow��6��77�������ߋƯ�7�}�=���w���qP�y?�K��j��w�_{�j�����_���7�nU�]/��^7�n_�ߞW�{�x gt�T8 ���`���x���N�������_W�d�8��@�o�DG��:A���ڵ�mSB��U��%:����n�ֹ���ƽ/K~/���x�W�x���~y�zZ񣟭~�ŧ�6Ȩ��G�0�1�x��@�w���ͻ����mE�����=z����W�/�Tg�f~~OR]&�Zc�3��w��>=4o���/M�-�������^��o�ߋ�{W������o����ţ|W�x���^փ{�� 
��]T�L�} L	��S& �cK�*���ݝ�����d���\L `��\C>�0=1�T� xG�X���޸ (@�|��c�M���������������o��ſ�߽��zo�~�o~u���ѿ������>����/�*1�]���~߿�����߃b+��W�����^�v���2�>���H�}|��&~�Y��}�?N-��u�����O�_�����so����������6�������ob ��( ���x���(�뺜��ZV����	�2P�����U��YwK���6�W"�a,I�uԒ��{~rb#�_�|��c^T'z�eq�8&��:�4#�Vm7Q�*.fUʻ��)����c��H0X��\&�ռ�T.x�tⴭ-#��cҝv��=]��z�����*i����}_zȪ>��xDg���=�$zbc���v��[����|m�v����9�|k��o������^���׋������_�E��v綿��W��w��\�������X'�.iA{}�uo��=��=_��|����^��^6��5�߾���P=P�{H����y� p�>���8 (��'!G�� t
�~��P�������7��ݏ�}�">�!�1{W-�\�Wη��x��o|\�5�w�_���-�{�z|m��<��*�Q�=�x�lyG�`pS���s~�����}�7�/�����_�)��z�t庖@�8��	��[ſ^=���~7���o�����^-������/��O���{�>-��m��\�7���ϝo���<�֍����E��r����|C�Q��٧����h�|G���b��$}�����/k+�ͼ^~_�}Z��+�����/>u�oM�^y�x��*����w[��E��}��ίm�m�u�7ux���0>������/�f�}]R�o�F���}����U���W��>���ƾ+������\��}m��Ͼ��^���xF���@�@<`e}>�x�����6��ε�w�^�z^-���ߛμh>#�o�=م7>��~���eL�Kƾ5�_u�[�}^+�n����x�>�L ��@�#� Zj��������=-��[�~W�|���[�^>���kگ��r��/o��[�w�S�>�#�D��Q7-��J�z���R>���zW�i��j7��ߍ�W�_�/So���=������[����[�~�[����=�g��F<.=P&�E��6��Ƽ{W���>�oJ�������
����5�'^]�!^�xϹy�E�zm��}��o�v�|�{��W����y���W�O~����{��7����}m������+�������W��� c��쁖G��`s�{ğ{��zo_9ȼ�#UT�N#��>��H�>:j�@���>a������^5��5�w~�KF�_�~w�/���h��]}[����x������>���Д���{��8#n���T} ��o�gT$��~������<+.�V�D��D4�_ig](���l�R��ZY�i�]�d�ǖS6�q'b8f��f[���x�	g�~q�M�yΔ�`��}�zK�,�,�n����2B7�����)R�4�_-O8��~�������>����=�w��1�|y��szm��ޟ�O�߾W���+��׵�����������~�w�Z������y��_��h�������}�S� >��#��k�C��`9���j*�9�ڬ�<#� L�YJ=��_W5��ׯZ�}~��o���/j��{o�����V�W����/��k�~7��-�{^M�nom~����w���x{���L8�D�$��
�<yǊ��[Ơ������zM/�!�p�DH�!�SC�>�/����Ϋ���ߟ�=_����|���|}[���/>��k����������" (��ZG�0 @�FG�1�x� �����&=�����h��
䌿y@�@.<>$T
��=�x������Z������o}�|/J�y����||����b�U��|����:�o��ο}��m�|k������hߋ�59�h�B"D}7F=�^muY�cu��߽������nx׵x���W,���y������k��y����}W?7��G�_#�t�� Ǽ�Y�� Tz�r�������ƍ�s���4_W��>� ����|�1"8|�|o;7�:g��޳�?}p��G�UX��PUh�-���W�{oM�^5����k����;�:�U�<�?�{U�s~{��UB�zc�<nn ��1������D}l���#�>���+��U��
5���K/���{�<c�=����x��o�����E��������~+��Z�������^7��o;x��x�k����zZ������^->v��}xޛ���
=�P����3�C����n�V���=p@���O:����&��1L1�� �Gўs" �"��2<��m�o��~_~�_��j-��:�{m���j��wm�/K�z�o���
$8��@���͝�I}��7G��W_z z�c��ʺ<�(��P��ѽ�����Z����x��u��C�xl(�
$��}�{� 	\߭�������-�|^7������?@ ���<b*���A�O�w1!���m��ۗ�}��hܱ�(
Ǉ��b#�R 0<�( >R=H�s���|��~+꾯����~+��7������ʽ~�����U�i�[�#L`�}􈈱ю�ۃi��B���ތf��	�3M�s�%^��kʙ���:� nΆp�0!j4wYX���J��q�In�7��CNŏ�E��ͽ�H
�K��V3�%�KF`�c�^G .*���5ׯ���/5¼��'�{������'�5+���W��Y���}y֠]���ͼo�~v��J�n?ݯ}������^�u�����zom����������?���@�yJ�b#�Dlz�U�=� Y�����V��k���k���4oƾ/D��q�x����|s�Ws'����} �W��-=v�+���=-��_n��zZ7ߝ�������;��n�������y����߿�W�_&>�*��">b �/��E >�!?iR�<^[����Y \l{�t�}��y�7��ݷ���ţ~6�������A^��׋|���+�v��Z���Z��y��o��h��|��k��+���������k��~��~->ur��ρG�yبՊ�ܴr{eʪ�qC�DG#�r���?X���>u#�>��DD&d[�soן{�v��n_������F���v������{���!"D_�c�>�1�
�o�2�J��O��j{��V$�a���ء{�:�'w�<:�Ϭ�²}�d�}�ؕ��b��|l�jio���Qb���q�:��<s�[7��W�����<�݃״3J�Ph�6v9�ki+:�\a#�!�Ȍ��u9G�$�D��R��jÄS���ܛ]����z��:���k�\��g��\>��N'fS\�8�!DH�V����}c6��-_+K�y�@�P�̓�[-ř#�wX��Gs�ഺy�����^ں�U��ϖ=�6z�3V0,����-��5��xa��ϻm����NH�+��W���L�>��<X�Ŷ�����1�Z������Y�b�Xe������s| ���W%޿I�}:������i9���'(,�J^�Ý�
��+�c�lkI�Me�Z�s�n;y���ݞ[�؋V�)9sI���;'�D���67r��9��[3����}��#���]��� ��꡿qt��|����ȟy������ɥ\pq�\��^ޱ$qοp�E]r'�X�iu�C	����s�9��6�PQ�f�x �e=�D�ҭ�V:�+4%V" ��DÕ��}c��3�ۯL6z.9c���<�!Y��((e@���ww�C�1L�%X�"��B"5�3�AI� �}9�T�룣%�`:�Q��ܝ�7j`=�q�Ӗ�j�/u�:n�#��0!uz'I���Y��`�����v���xn�y9�[l��{��L�p��@6�b/���YHƓ%m:6�jnFL��!�I��������C�j�`.�Ry)�W| ���W��g�4z|kK�q�c�v�̰m���zmE1S�����O��ک���L�6���y~ݴfQ A\&WBg_qgc�Zwң��*^VS�qY��]yag�w|Fy��ɫr���힪��p>R�<�_����7
���V�
�s4��WZ�$^�vv�C�R��ys�DE0���~��PP��L���Ѩ�ǇmhPX�z_
��q^�g��H��[8�b�Q�φe�Kk�ʯR��]d�
��Vȣ��*>��3`b�;o�����!Ϫ���=M"[�;�ɜ��uQ��3U���)�r.�k�ĝ� �0��s*mR�K_#����s{y2��o3}��������b ��g�V��[��6���Ԣ#-�q��*[�N��r\)B��L+	ds+��͹�Ϣ'r��g�̅WY��fOx��Z��xzt{^��{'\��C�[f-Ӡ�9��ںl&���E�j�Z4���	�r��Z�Wi.�G]OK�n�[��H���b��Y49L�w^q�9��Յ���m�FOV1�8j�*���hMEEz5�S/�O9�F��R�eD"��[<����Q|Cs�ї�����kq�2`>v�>�J¼Z�J��+�T¾�������Hz���|��\� $6����t�qa�y$�Q�=Ć|��͑���ס��xX^J>��X]���S��VR�C�0����x"�Q� �B$�I�̬
}�0��uݐ�7
��6�&넱<�8������'J�^
d���ƾ^�xXJ�c�����Z�>A�Gq��3^[�^�9:H�s�8�`����^pQ�I᨞�cٚ4�Kv�Y>jb�,b�ϕ^�r����Jrm=p/W�36��F��R˰�V
We�#S<o@��i�r��+PcA�bF�_��n��(Ƨ��tqi����p�	�;vy�ޯ��6�;w��0�<���=U�M�qd���%�	|��֎�k!�$DE@0����e�q�e˭Ѵ�t8�i��M� ��qME˰+��Ñ�.T�t0xb����Z�����4�Wa��dzW���(sN��r��L�3O2�v�i-\ʕ�W
%��u�_c���v��/Yr���d����H�*�����f�r�=��zb�	u�UK��h���f�]�c��b@Ýu辐�����Q�R�؁�q��ͻ̩��3���a�E�BX����Z�B��&����2�c�V������9}i��oe
�
*��o6ոș/	�.��Н���(r^���J�4CLT�Fè�יID)�qΕV��S%2�5a�U4�d�Tj=a�~��[��Dd����d��DBخjVe�y��9�KE�	}��Msԩ�u�6�d�����"'�Rʍ��p�Vo�y�!<��!�� �@V��tW��V旅�8��������Õ�r/h�S1zǶ�T��k�g�*��u�mq��>��Z�"{��*���*�
"��g0p���@�j�6,#�z�ܻ��Ў���h���{���X+1
m$Q��YLZ���'��N�mH�-G�s�"�C�qf*����k���.d�_E��M�{͚#bAwU�utRs<y}U�{`�W=�,�	X4�9<�}�=�xD�k1]\���Q����Qo�ߞ��uЅ���ĕFG��Q��lr;D��̨6��;-O[�l,���>�r��9�F�:�Zq�����؃D�S���%jUͬ����xqMUz�^�up�ⶬU�e�q�!�i����mٌ�S�Fl3=�6%�\`��RZ�Y���$���x�CGi}��; ��0����22r^N�"x��5�g������ۻ,{�H�|��b12yt�J!Ŏ.9)��W.�
0����R��c&#n�a�G<�� �ϫՋ]'�r9*�U�����8<��������Џml��N}����О{�b]���u"^e�k��N@�qD�z��e�
��N
!�O0������Ni^vL�e,t�x��ݫmF6��f!���ix���gу����Mx��'{c��R��k,ѕE���ԤlP�����X]=�~�~Co���y�r���^��.��}KՍ��	�oɈ9<v}B2|�Mӌ��\OҙΥ^�)�����s+G;�z���=5_KQ�/��X�a��Hp},����s5av����QM��V�?^�yŘX��]�5��jxC�Ug&��4^��ܭd����|Z\��^1�������][ɽ�Cv�^�uuKH�a��g��R���3{��jƹ"]{�v�մ����}U�����W�Ƌ���8H�8r#'F���:<M���<�uׅ��J�\����9�j�'z�S��Ow�;��zȽ�k��vʮ
�W��n'fS\��\�z'����Kۥ�դ{����Z�����{t�y]�3ơ�܌��N�P�@���w���	�y��׽Q/�֮���1X�7=�)��u]7%e�u���@�>V��$�0�C#��ge�A�4AE���,������c��zTa뭎pp��`���r��`�b���D��C�f�RJ>:Dq�=M+|s��/�>Q�-���m��&��9��z��p�{�S|��J X@�:����]uI�v��E�ё|��Gy�i�op=���{��;�Ӛ�H>e�*�:]m3Y@yP5�HtN�U�i\)������?�}}сq%x�>D����`{䝃��gԈ�g�`B�t�~�u�o�iߑ���aV�]���/$}�U XY�V�AJ�����&�U�-b�� �:<��&7Ҷ���FI�v�7K���x����]�ؽ\+�|�.�Z��u��n;���<
���U�����9�m�x۠��� $�~�ܗYS�� �;�vܤI�V��>���*\����u)�ev���$�@߯I�8n��lY3AEO,��ľ�� ��޳|����n���)r�iPrkɺ�/:q�h���T�׺mL��8��ws#��Z�Z�nL�����I�r��J�~I���3JdѴ�Dsf/@�I���cC�K�׼3��U����5��~v���᮳˯,$�V����@[� �>�Z*;�,3�x;�b�����]̳��@d-!�ȯu��F�P�;G!����',!Z[ǟq^+��64�\��b�Y��{~�n i�v>�Vƫr��_`��=wl���=��x�/�߽~��*vƙg`�/\���w��C.�b�t�wo��Xh���@�1�f)�Ѫ2�*bz��zL(����K��)ϵt��`pk+��$�Y=J����bd�2�������)�3�Ґ7�,B�e���2��yƯ9��PQ�:rN�4�/��`Zc��`�+�;[y����L��Ψ$R��VJ���V�e`v�ہ=)�yyO0�S�����Y�G��x�8��\�k�+$~|��L'U}���z��O}�,��I�N���<C2�	�x]�K�f�u��1g�c����Ʃ%�x�`�a#[3�@���*N�v6F��޽�tt�(p�Zݝ\�,���E�����W�,W:��HҏSwWȻ�S�^�Jt����Ne)-�v��(�����jme���n9���ʕ�r��do�-��z�����r���nɶ���(}�c�W3��z��&��wԓ�\�k�-�+����\��֟���.��;�����ݺ�!�xEQb�B�n�/��^f̋�`S6e�8�'g1�`c[�L������Uܙt�=��
��7f�'��N���\y�w	���	Dި;S�mo�����(y�\�;n��,Q�Ĉ4p;&9���g� $,a��G,QK3��i��ͥ��Dl_s�6��FΛ	2�,�����Y}��N��`��</j�r�^{3 �)o��AOvW;�E;�,e̍`�Z/8 ��Ik����l�w�V�X�/P�6��9�M�~B�h�y���3;��&��y�`���¸��%So�G��)K� �/9�z��YѮ��A�Ck�Dr�ݸ0\J�è�r9}}�����Us��5�k��a�nM��hΨ�j�ВTWSC�ߪ���[��}�ټ�z �"A�Ҁ�M,���j�\{Sw ���ʤe�Kzv�w��}�1#�]�2k�S�޲a}h�/:��1��<�����z��Ua��z�,ۉelm�|9���9D�����3�o�X�	yƝe%5���:�A:�Չ�ٹ��������<FP���rě7?��׽�y���i�om5�&�N��U�V5Oi!e��E��-7R�3�&���D���Lݳccu��9��j��E@,n+o�1]��-ɠ^�5:ZZ%�|�%2�v�z�c�|=ϳ���l�1�ӱ逽{A�RZ|si�`�0D|� �Q,�;�Mnl�ۍ�c����_j�z�f�o��`�qΉ��X2�m)��G�}M�2P��v�{�[s1;�us9,��.�ԓAdf�Ō��{�ݲ��5:s��`�Qԯ{�Q����AN�YV����]Q��ʣ��;8l��9��l:kS�PY���N���li=u���]��˖6�q���>�o�Z�H!v���y\$������b܆���|!�2U�������-�J'o2�Ƹ8���}H�0gw˵cB���V�p&+�G2V��Э�w	�p3�^!��V)uM݇瞨D�A�;<t����퇐��}�B@��aM[m��8��T:t�_q�\Os�|�����rp�U�{�������w`�t�ױ5s�7WNU:`��	-HOI�:��v�D�<�K�u5(v�����W)^�j����A���m3\on�j��VԾz��7`�H[�(�w԰٩x�����5L��������F�2�0�D�Di@����,A�Bb�#`B��A$��0@���Dhڈ�H��$�ř3�"�	�D�Hd���H�.��	���s$!�Ҙ��q�&����$�k Y#d�M�#s��]�^9F��"� cIDMEx�fr�F`LɊ4Y� �#Eѓ3&̮�k��
,��r 
4lR���d�L���MA�iRC9!��b�(�"󮢐�&D�2D�D(׋t�\�:����)�&#!������`�Y&F)-k���4�H�E$!�BQH3bPj2\�*CRJB�v\Z,�}�e{�.���wg *3r�j����K���W\!Q���B�tuNki��r�8m~��=�xu�7VÚǆ!���;��ߏ҃�}�	:�P;���]�6]	v�gE@��"0)Sy3.ӆ'sc���"�1����8h7n�ȹ,�xoI��BS��s*����S�����q������v$�C��U�㺝tq7�DF3�x'U�O� ?}55i���9{����Vc��T���VdO�[�^��"�������&�b.]\AL����d�s����eޭ>ek�D�^����#0�L؍�#9u:=��t=��{�ގ�����}�����0�v�fɆ.�k�d$:n!��q�ExgJ�~�ta�s�RE{�vh��zfI�4Q~��#�Q^���i��%��g�C��]��>����p����_�b󱪋�ܨ|\B�L��ts�$k��v�N1j�e�~k���ظW�M=�2�Ԧ5#�+L�\?GVJ���k�e�5Z����Z�B�q2�;�Q�uϫ��!���C��>X��У�s*](��<��ڷ�\��8�e�}�`�����]F11"��߽
V�R��njv�Vܢ�����f���7���l�b�"��5J��_*����|�;L�䯽�r2��^�s[����v���qu=���eT��<OT�x'u�rcD�,��es�ӎrf�A��25v�UG,�2,�k�_����9#f���G��~5�u�U����2�T�<�%���z�W�η�C�Y���L�v��~�Շ��=�Z.��e%�؍sՄ��]R�[ǁ��� 8� Jw����"�F�!�`�M��^�`�b�V�+�t
��SK,�Vi���z ����lӗ�qO�\��4ܺ�y8E���(�]gDU�`��A��[�Pl�W�h�X�懎�+{׷N��c�w��X��/�D-����%]t,�d�i$�3�D>!f��cd�i���#���L����l���*�s�dm㨅�������D�����w�}/��k�μ�>�� I��뚅Ǖ�b�q�x�;N
�e�=��h��Oҝ@��pmy]������@C~�H_��:�tT�и������DEih�E��\���)ų��H��Y("O�������Z�";�LGʼ.P��Ӗ��{_��)���'��8���.J=]��)¯	R�Mq�'A#�=dt��&�Eq^Υ=�-�ffa�,Q}��Ԫ�l,u���Q��7v���|/9�1�Of2�7��Ӫ�"M乭R�H8��^�R�I��m�����d7�:��u�=���y���ʨ��G�嗏��X��;˅iOv�SO�l�p��.�Ex��w������{��WMgRUN�2�(�>�ҦK�r�5����Jt�D�z���d����u35J=7K]�qS�����%���@�;�یmUѸ�bW����Fj2�x}K'��|��xu婚F�OL�t�.%(�R��g��n��L?�+f�ns��4T����=ix�겗v�v��Ɲл����|���Z0�@ RJg:�y��6+�Z9݃�w$��UH��1�I��u SV/K�.��H�k�*�t����:<Mʽ|��]x_�oҨz�/ѬŖ�4���+'OcSN��W��o+b�DD]׌�|Tg�'fS\��k�{�#�3�Kg���p]9�y�W,�`uM���{t�o+�����e��TDl��񑈤���Z�☊Ǧ���1^�)��)��uR�mg#��E�l�G�s����]��v��5N�4�{�H�5��ij�8�zpi󇗎�dXt��䬾��)V0p��uOg�w�9� I�RX�b�Y�NȎ48�TM4���a���>��[C� �!��9�h�U�j���t,�pcv���'&���[+��ɂ`�N�U�T�+sjF���}s��>��νQ�^��\�q����Uh�OZ������W*�|����w�/��v�+n�0|�+7��v�ܩ2�T��Y�~�������e,��j_Z�;��e����J��=CJ}���3�ۯM�FE���H��s��['w��k��r�I�m�����RQ��PTv;�WzW
w�z4��E	����k8�}{�m)���wc�tأL��DB3�0!uz'I<��S�'kN��.���ix�ʛ���w����V�n�"�8�Dכu�%��0!��姎ɂed���������9=:��:���_�P\��XJ����y�>�/ ,o�*��Z�%������L�]���C��&�����ޕ��O�ͩ
�2h�u�!�F1~�����x���@*	���/a`��>�����!i�ז������;x�ÜW�Z�4��2z�?R��`�fi�5��|X�Tk�l=�𚕘�zUfǃuta����o����&]7�pW����G������b ݏ�XHW���c����#�u�EoŜ�z���ɸ�~�T_��r��Frct߷��hIZ�Nd�����O��`Z�9\Ǘ�XaS7��U��YE�$9��������5+�X;j���g�~���.�Y׽:�Zf
c�H?vZ��9�r+��j�H������efJ�x��]2���.�����*�z1��D��׳�]���m�/D�Qks)B�4�$���U�U}�������$!DG��Y���l�s�]-��涺/:rH�Qd�a�W-���]Ά٬�,T�u\g�	fX�d�ɮr�}�y~q��n�AF���O�s��=�W�9���/�=1i|N�0�O�^�S��4�}����a��6ܶU�r%�e��ٷ������}����E�q��/���ע}�?>W֩������]5�z�e��%vh���2嫸t���j��ٺ��'A�'�� x�i͑���pn�?�R��ўTg�i����ĳo�t!�sz�q�p�v�<���z<7�G��7K��F�d�u��s-���zJG-�^QC�b[��e]>;��Gy�@X�<�$y:� �B�>�s�3W���;�ʧ���=�Ƽ���\�$p���/+ ��"��f�N��g7��_f��l�1{�hC|tS�Ñ�#e3q�e]n���t�d�@���H���*c���Ew(-�]�1sl��� �fCC��Lw��a�`r{E�ײ^્���k�"<��}��3oE�J]��l��4�h�M��sA#��h����42�ؗ[�"�e�\e�&�o���w% �k����{`(f�e��݃� X���+y�y��a�M`Jw���R��\���,'�� ��O���b����n���x3չ�t�{}�hސ1}
�>ezx�b����4�v��)r��(���gU{\ϗ���_h�廊�\C����^� k��7�N�#��6>��bA�\�f�C��Ι�G���9[�����ˁ�k�f���S�c�Tíq�O��۠`������|��Ru���A�r��}M*�V'׫�7�j�dxM5NG����s���-��� "�m�����&*�A���&t�e"Q�� O���ԙL�\Tj;iu����(�A���[��f�	֛��8k��&ix[	}���6#\ǵ]V%�t�.�Vr�<xf���^+lm¦?Z�az���x���a�׮�߂���<%4�)������ǻ���V������lx�k�/�5���ԥv��n[<�z�d_��Q�" ly3fz��nd����j\��7�+�{Ԧ	u��]������g��2��B���	W]=%�%A𣍨W�zl@�=�i��.�h�	�3�^z��D��iJ��0���QM�Q�����A�W&��;noK���O$�g�x�4���� ƭ�U�<B�0b��vW���M�x��Y���<��w*�bp�k�Ƈ�'��p�8#-�Qu=�\�X2C��Ȱ�9˅��u��o=����b
F+��N�����bي��z8�mA+{��������jrڝ~����CR��8�9��o��S�	��;
f c���lF�����*
��]�o��,�V$��F4�A)�_��z�B�Kz�;�m�ZZ.oe�p��/x)O�W��u�=��'�I�\����7ژ�|�������� �k�����}7��Mv��=��1�+�ׄ�J�5�T��#����(I�rf/P�.]k���T�wNv��~\�Ë���9�d��.#^z+���c�'DXp�͉���crk-=�3Ӫˢd�e��r�q��WDc199q^y��/�}���Ӟ~a[�X������h�}��k`��>-JF�{9_'w�:�tla�P2W��
N�xy�w�_`+x��p�+C�7.:�'΄�8Ω\N�ҙy֯Ȑ�خe9Q�aی�����fsE�y�@���ypl�҉D(cBʜ��z9c:�F�Vl`�5	�j�!]dvp��:�,�U��rN�¹����@]�*�!^�����y�P��^WA&m��)Lu��5�.�$9+�M\��&�D�hxWq�y�%$����	�s^�.�[x��1^�8��9ijwU�-��=d0�v>�7%8{Def����'gf�ˍ-����7���#Cn	Vs���*���ac3w9a�W"�>�꽃��НSe:�fo+�����,���Ăv����7���+sZ���]�<�۾���C�~[&1��yNX���䬿��ܶh� 1Y�_g]��y����X9��U�e���I�iAF����qt����,c��T�®�8�����/��G����
L��K�	�>����>�;"8׸�TM��9�a��4���%x@�w�ق3�9��@j>@�(� 4�xl�4
#n��T��x;7�Y�	v���LP�#���1��d��!@BIGDDf�3����'�%uѠ�#����״�d���ɵq��<����Tn']�߱�M�Q�|�B=!o���u�s���e=���cUX-%�(�
G&X�ȡɫQ��D��8�D�m��X���D���!Tm��:�DL9ׂ��k,ɣO:tn�gj���E.QC/�PrSs�Z�L�W�r\^�[�/�W{�+�*��g�A�ƁS�[9�-��~ޕ��O����	�Y)�F����v�`)���my�k.0���eqY�AA��H�5��l��ْ��-��.�T=4z5���e���;ٗ�׹7.��F����U��*nUɞ�6n��m�Ԟ���PZfV�@�U�ס��X�)��M:\W����-;��ga�ri�d���꯾����&�v=�F���U	:kN�6�Sy��~������]ya`I��-]S�0����y�mj����`�y�a���0y�@�]̫9]^R����� *Sy��䙛��h-X�^�10z��n����8Կ/�ߏf�B�4��r�	
�[���~�&�&Uq��^�a�]�����qh�9�Ο9���}���˺���d��2cPr`*���>q�NwP��tՏ|�������Љ��:l�ϵt�j����yӒB`����Ur9�wW'�J�$��bg���:�g�%��	e�\�2��yƯ9����R]ۘ���=ȐxU�^u��/U��&"M*'�:	`����[�Y�l���U(6Q�3B�c�;!��4pk�q ~�~g��%�ᵯ�g���pik�+$~|���0���Y.�;�z:-��/BQ{���ˡӌ���j��V2@Q�$� eD�&,!q��2�'��jJ���Ө+G��oT\�q���D/k���\t4ݻ"�Q�!
xp�Oc �T�wM_��/-o,�u��sQhVV��<�]f���A��]���5�پsg!�}3.4�d��bݥvn���iVs�e�PȬ�G"���y�{%�
> �i!v�������<l�H���:�T��õ[;�=�e�ek�L_e���ؗ��k�;&�f�Q?y��tPZ��X��tB�|s��tq7�DFP.��D�32^++�N��ԥ,�QJ�" �R�؂��ȟ.+z'���F��w7��b�U���S��Y�Ӽ��$����&îh�(	����#��.�b�3A�{�<��*�^v�#Ι��wZ��ɛ�/$� ��c`#�.�U��5�t�W���ޮ�*Oh�j�@��蓮��Om���I�6����*4�2N(�}� � t�6���i���N���K[���#c��CN���E�9�n\A5�@���XC�7k*CW����-#�5��w����hҢ�ܸ��FB���9U8��1�����X����M!R�k�>O\$�1�r����샖�hz�{\~�M���2/�ҙͥNC�Xj��4v���Ծy��W�����L��[�G3��^�'к���Gm�-�<o�7�Xx�i2���j��[_u�9��_��xυ8j��#f�\-���Iy��cڰ��*��޼.𷄪=�@R�����wV��[N9Ն]Fx�t�|N��{�ps��go�4�W�.���U�N��s��Gr4Rg��K0�u�'�h�3tmo���;lv��xJ�̋�8n��ڜ�Ղ:��:Os���Esא��.�Lگ�E��Ϲ�e��{t��4�[�[x��ʻ�rZ/4F�2E�u���K�R�v� v�I�D�y����tr����t.�F�d\��.5#�Q����t
Dp�v��ob����xg6Gp�3xehb�w��F]�w�$a]12����U�,T0�'5���xb�r�^�^c�X)�u�z]���Є�{��tXLUx�4��K��!}�W�c�OmY
󌈪9�Ӟvz��h�pcAJ�冧g�ý�������^�R���8�j�,��wv��T�y�o�����MvĘ���W]�U�EIĩ��!u�
*�Wҡa#���ps�І�*V�F���	��2��.)/��X�k-��=��c���{g`����9�٠GB$�+B[M��|�2^��u"�$[�]�ۛ�@֛��^�,��6b��V�m���4ā��V��ûs9� 
�LV�n����u��|��ꤻ�F��=&Hl�i4�4k/;�=pVe�*�cn�28�>�7����CG��X��&x��8��ҧ�6j��l:�U��Ty��SF����1&���y:�P��|T��B�c�f��veR��a|k���|8��7����#4�p�� TҊ��q�p�z�f��m��(2�a�Y���=��;-G�#���-!^�"� ]�.�կ׍q��4a��ף�1�!�v�8ڗ`i�7�`2��$2-�SmO�zj=��Z�F�=g;�gCy{-Y���"�L���۶��Wf$��&0���m�+q�$7AXӒ�_IP{�kf�G��8㬽"�����0tnR�ڊHOY̪���cV�n�����J:je�Ou#�Do9k 1n�4���w�'��ʐ·P�hT��Q&1�%��.��$������|<��gC��/�ՈB,��P��h�4,��t�
�*�.p��H�m�[ƕft�]A]AGp>��8��n ��ɼ	����aY4v�w;����:���P[������﵋xZ�Wu�0��g�h
�'%�@��n�]YʘO�.�vF�V��Xn�Ub��{sz:X[4TX3,]��e�� �w�e���=o��L^��Zw%��;�v�0Ñ��6��)�/un:�`rɻv���R�.^�mַTQ0���-�縇����
=�O�p�c�x�_b�o����`���yN�w�E�Z�]�XG>@�` 5�2�a�x����ɝ
��_��u
�8#BD��5n�(����*Wd��r��E�I9�È6�"-����ˍ^j��ܮC�cx�<�32'�3l����Ϥ@��@ D�HT�J�c��o�FlFM��(��d�#H��&�!�C������	����),Q�H6"ѷ+r�b6�I���l�5Q��b�j�@�UwtT&�J-���IX$�b5��sEEPQ�2E�IQ�h�͸l�ՃX��6ɍnW4T��i2I������EW.�mF�b��3Eɢ*LTlP�76��lTe  ������ټв��Wj�>���`��A��2�rlԖ>�HX���4o���1��콡h�)b�Y4�p���Y����x#ˢ� �7����9��C`��x�i�a����Rm�;VgJ�2�W�UB+���q�v)ZLvZ��Q����E{t�_���g��C�2/���R�@��>L�3ԣ74�,+�ƫ���k0�/��G�;n��-��bC��u��N���Sк2J5�x��芞m�Y5J�Og[L�σ��
2�y}v
"Vϴ�O{��#lc������co�����Pr)V��x�UR��[ 	kԏ �yU![�Vy��y��>K�t�ʼ7�yY48--M>��#�轒a��§ڐ"�m�_�鄫�!3�6:oWGg�;l��pNv��-��Qr%�ǩ�R��{('�'��#Ǒ"��b ���-��^�2nGL�[�M$�}>u�8��^����q�,�E�U�u�*U	��T���ȅmV~���w��Ң��µB7S霞DN)��ޣ
��>楒סˈב^��N��(�aa����q�g���Z���{�L��bS��=D8ɬ�w/Z�UьD69J�g��Y�n� �Vפ>J���]�452�o*����U'-kai����?�3ZS;�8S�D���e���u�]5�@�Ob�M
�M���u��_[\Hx�E��R�/s��c�;K�<C*�ږ���5�ܺ6�k���&�oi���⧌��������u�5u���>�6�,6���9�=��e;�/��ޜ��Q��P6�^=DJVm��G�r_.Ҟ��p���`��:Q��L�L������^|nkɋ�F58��Q��T�4!���߸Q�F��U�\<�Z�ҩ�g�H��7/_ �����/��	��ıuK�M�j�{1@�N�r.��Q����]�b��נ�ߜNʃ �����wr�W�_?T��0{M(����<��FT�Xl7��c{jxݖJVg����!9��;y� �.��u��k�p/d�R�����:������]�1��zkqNY�o\)ܒN��O�H|kHB
+UP]��Ӛ|��v"�*q���^�������^�]L���`A�D��I�z"��)%`ڐx׸�TKJ���|iBqQY��ɣ[�Wl9�x|���X�<����0=@O ����>�_X�L�v��f��ҡ�K۸U;����tob��������(
�T�xEیeߪ�h	�Қ��;j,P�j9ScBRe��S�����ܽ!]w\��'��C�$Μ�-�i��(�i�Xl!��;�4@P�!޳�����A]��Gx�k9�NFEw�;1�i��]�C�H1n��yk�8NJ�4���-����J[ܦ�O�_UW�Urk��q��\�U8��Jj�`C���:�&���:o3���.��$sQw���Kc071��n�T�F`(�~����u����ը��"|���؋����B�m-2F.���Qt}�b��':����X޿8�(���%7=�t�#b�����6����[�<��Yz����]Q���v=�lޕ��_��	��2h��#4�9���l������fxcb�j�IZ��f��P*\:=��쥶ⴅ��]ya�»&�)�C�F���$*��a)�V�;`7{f��3���"�-�V9�k�l=�����䰧2,�Q+]qi���9���n:T�Ρx��[G��f��� ��g�V������t2�B���N�F��/�x���n"(^�,#,��󑁩��9��^��������v��[e��0�7&��R�U!�X6�����L�2x�8��|���u:��ϵtߛU�,��9j�=Ǖ�'�/Fx=�v�ѯ3��Im�Ec��)U#b�@h�ٖ!_�e�\�2�^_޸���˿4����TĮ����7�^��w�"
�R��;[wg�fuevp�4e�`��>��&\�lU�V��@m4�sas�[ՓQD�1��6��1�.�o�y��ԋ@�6-:���5z�է�����v��@�'���g�3#�)����<=��T̍-��Щ?_�Z�p<$��ts	`�M/j�Oy�i�b�]Y���ڍ���x�S\cro��bA��×��̎�㢏�pP>��Z1�����P���m�ۥsVK�s����FC�G8&�>«�(���z��"q1�``D:��c+�8�r�B�y01����}��r/���,.LLxf��������귏R��$DJ��N�o5�WKv:,t��]M�r"2�tTOB��ˋ�����5�J���QG���`ߠ�/2'ˍ.����F����2�Ln��un��ч�����-�OX�ʱ�fI�Q�ڥ@Wx�T�a�v1w���[�����K��۽{�:��p���}u���S������}Z�<k��\B�����iګ�uT��xk�OQU9�a=�$P'f���aH���� h�w(b�>���wβ��lz�V`����2���Œ�=�zu+s���3|s̍�Bn$f�uѬ��uALE髄�`�f���Q��� ��\�l:��;��n�M�WWwS��>��gX-��s��d!W;�$C�X~���]�����'C= ���΄[־�|u8��ίo�Ѧ{i!cO˯;�`p{��;��x����*~�� ��7k�d�<�������+��_-a�9�d�ѥ�*�M��̲��`����]�Z�~����g+[Js�/k��2�-��g���hP��G�-�9��z&��L}���z/����+I
|ӵ2��Lʳ8&�)�dqqo�ˍ�OԴ��=ih�XssشIA�B�#˫*�:�{q8}7�+/v�H�2�]���=�\��l>�ϝ	
�\bI��Ȼ`��7P�zeu�qX�X�z�V0U��U
؍������Js'ri��/�Ĵ��濱�.�ӟJ��^0�c8&��*�
�����.��ġV��̓�iP��}b��ҥ�@���0��8[�Ȉ58e��V�Я���J������}		�wmk����=���r%����$��B.�9�t�*![�q�=L���og�gЖ�B|MΛ\�~�s>Ki��fL���t)�P��bgR��㮠|���GӘ�ѓ��c�C\���WF�8c���b��Cv�0�X�	o$w-�o;I�]گcz�N�Օ7��4��H����Z�d��`��̞�fŴ�Q��t���H���.�w_�UW��E
O�/ow��i�9�A7A�9��)쾛��'�o��ɉм����#*{7���v�ƹ��;�V!ؕ(��נ�Jl_
�E�E�q�'�K�&�����}S�8j ���(�޿�]q���!�k��H��]�[ً֟k��U40�c]�f��B��l�!�Y=��l�}NƯ��uB洳(e-}��[{6�N�ְ�t��ŋ�f���fS��{3%�vn��:D[��>[U����}����Gi�L�v��}�g��O��}S�?m��y>�~|.�Q�/��5��,�,��Ǎ�G�͸��N�ύ{3�F��F~����j$-��ZZ8��u�>�z�a{=�E�F�㓣��>�J#�n���n�y�������&u��F��%Ww�FTrb\��	v�j��x�v�9�U���bvd�5�UX�K��K���*�vq��a�	hCb�f�Ŭ�i����g�cY��j���j��7�}��,����׉@;ucЎ��{�c�:�;�\4/�bXqʁ��
�oxG�M��<�M�kiO�=�{�t�mK��f��]�V�f���� ̋x���I��"��`�/�P+V�W����}�;� �ב[tuo�㊽�g30��<�EÐ�#d��%*ړ�=3�4��Y.��G���e	]of���ɭkֹm�ͷ~����lwD�K��M�ԭb�#o�(|���#�jC���S�Ͷ��	t��]���%��DfT�m:�-w*�yb}��s�V�{�V�-���u�*�tܛ��w���Ӝ��y!m�a�-�\�DrT�eM �C^�j)7����BJ��y�%��.���#���5+rk7�.Q�˙M�4!��l�*��3�Rk��eT�GW�*:��4����|;���ɝq��B��b�9���y�+�S]Oƪ�����eY�^�,�o�y�7�[��v�-R���Wy���u�Xr���m7�Z��k������U/3d.�;�HOp2hj��f鍡�xٲ�ie��Ӎ��	�)Y���6�dXJ��Pv�Xr��\/�V���Ia�E5e��+�&[��^�w|�n.�A�g��>��~y:�mu[�2m��r�^J�w���'�Y�;;��<< �p����](���w�oyKլk��x⩤�KKD���@F|U��p�m���)Z伌��$V4�)���z{�{�C^�j$�uj�\�]�p��;�:�]�$͜0�oaB{��曌������uM`Q�tMm���|���=p�D�=^�A������������LOdQܚ�g�K"^��Vv�V�l�� �%�	�!-=[�5�g7f����K�[Z�T����pK,6�9O!V�.¨V�l��ʄ����r�m�\����j�;�S�ﳟCYx���w������ ���,��-�������y_]J���[X�`�3�z�F7-����|�h�]y������}���_L7�=�Y�IDC��P�n�8���=�ϫ��}��Kb�-wq˩oFW&�ýlJ7T�-�E���a��Lj�`�3w(��x�߃�>�̺�ao}�J*��,���,s���9[;Wif��1�}Om�vB�^⁹����ۢ�3� �ݻ��hǤ�W����x��!�}Xv
Å�	ѹς�\�O�f��z�<���tG���_}�܉i�;>+��Gۏ�SH��ѰAO���̱�-���+h��Pu)hݶX�������v!X��D�u#� ��V��}�fu�x547G�����k��Ѿ�>���8���ޅ�F�1#�lŭ�w��S�=^�����;2go��Ģrj�\�M�9m���9�5ى��\F��׳w���?E�y�<��w=�nV>e�-a͹G5���au��&{�G-�3���#&-���M��+#3����w=]η^��؞{��]1s�wN03�|�ϵ�����np�c}��oW%~ȝآ�ܹ�t�,�y�;����֚�sެ����q�/�ϥ�4ՠ3�6�n�V��XqQ��'ϵ(�Im���	�3��
q�@sNY���ih�
����Z�)��:�.�4�W���-k,&ڰ��W�a�NDdRT����B���9�X"ga1Q<vL��ܡ��9z�x}X`��OT�JL�)�s�tխ��څt�D�E_D�޷YO���X����R�Z�%Æ��I���:��^טv���ROK�sKBr���@��E�ِ3LԱ�i\D��N%U�/���V�q�xة��i�ٴ�Z�v���0�^5���U��\Fw>�5e,�N��܎u�%�U�UI�W]P�*GRw��klai��&#hwU^�F'�/mSܽV"����/p�F�V:���-����1��W:�7�{4��Yu������B]*
�w��=���:������3����gtS���$���!7��9��)H��y����4&�$�6�YNNr�p܎͋�M!�0�F�݉
��(�z:�m���,�{�L���	O&�3Z\�R�5�iÿCc±*F�Sn]aT�.����+�{r�Z��Y��z�ͪ���hb��Nd��ݕ/vU}wva�����j��W����)mb�N�'#���Q�ݬ>|�Wg��{^�O�~��V^UY3s�Bs���J�E&�����L�&f7/<]��5+,Kݵ׉�Ɍ7n�53w4���?��x����&�ڞ)���C�^�rwQ�^�(�W�YZb����軺a�;�f�hH]�3nМ�\{A(���O
�l��B�hQm����Ӝ6n��s6�/R��d�垻n/�/�vz�[ë;q�IϘ�{�ݹ(g/��g:�8�-��Q�b��xCH��Q٧|�J���<�X���֧d�W4VZQ��h�[]�����T9�r����v(�Z�,��N[z��gsD6�v\CO���wry�>��D�봢�v�Q٪��i�"���.�w�y+pjf��I��γ1f)��������K��z�9v,p�O19Ѽ�D;�j�;�er���։�B[��45 ���F�ea�׸�k{�%9w�,�{ћ�o��#6$8��n�	3F�Q����K���򚌠:�_v[�W����p׷XC���Qk*ec�r��:�E�c]X�n#�a�3ݦzp����U���f��U���H�;�]NY�վmjL�!ŎK7Zxeu�\��V;�/ۦ��F7uuꂘy�)W}c�o���4��p�158Jm�� ��'^�H��cA����T���R�k�di�l�յu ��$%j�B�h�VxHe\�dl�	�� �<�V�v�ov��s���VJ�9a5ذ�S)ϲ��-���m$��P�|��U�;VH�W8tk��6���c����}�۩3f>�]�����9ƛ�D��/~�F`]KuQ�Gi��ؓh���еj��n*/*�i	k6O������m�:�����_q��ܷ�u�r��7�:�aђnQ˭�龶U�W�9�u��!쑎�YV6�x֪:�`�ѵ�v�7t���{iVh<~��ȅ�o��5�0�ʼCb��V]�a<]=�G����ܜ�U��'�Ւ��q�"��'�g}��Nӷr���V]�ѹ��w��L�46rtXU���.@�r{Ɵ!��ʊ��)Cj�$1fvlje�_Rul�+t�7X��{}����`�M��p�e5�P�����۲�ik�;LIepz��J�n2֨�+8��r�TR
�K�[�#�}W�;3��ECn'Q��ar�Ďh��/�[�Է��u�J�6X��C��U����E�o��A��D��1�O�`���N��t{���z0_:)�6�Pc�P�E�����u�����>����%g��/��C�j`�T�,<{g\������r[θ���G(�n���cy�̷bMt�X��[<�)��
YR��Ɣ부����Y����r���_M?�-�>�MZU�S ���-�k�oT{lCYH�ZaȎ�����e�v�4$��Es6zi�7��]��B� {S��;7,�b��s�R���L;6�* kol�*b&�j����Mg�4�*Ҕkj�vm��`���,�.�b�0XڶJs��{��������߭&�"+2��&�W��h�b62c��Ԙ�V��D`
R1��&�%�0Q�F��#l��I��F���3T�h����BV1bf�-�H؊-E�r�IF�� �L�cQ��-�.]�ҘDb7�guͮ��FL悇v7(�L�ݹ�]"�&��ة.t��.m�Nv�
-��њ�����6.�4m�\�����e�hյ����r��[5y����B���M�}y�fC��&x�5W�aHܮ���n�O��u��I��\ާz6��G���*�ܜ��/��w�����5�c;HSF�fG<�fH4��5��gN��W֢�����ӵ2�y�|�v���7�.�Q�m�r��5���gp�QX�N�[�P�J4�M�K�'۷�)�(���WV��9���6̢WW�\��	s����an9&�;o���x)��7�{B��wޗ݆�(��V�l��*%�ep=]���n���������k{.Y35EQ��^@M��1�A݀e�z���GW�iu��.zނ.&T��3�����	R|�����|����>�//��&m;�1�Yo�Y�Ѧ�s���vk�-�nR�EB�;��\�j�����e���3R��5;�}���u�V��{�m���$iZ��/�,qo����|,��]�9u�^��[P�BnŞ�K��2��!���#&M���r'�5�q�%23�3�j�ʼ����qEl:�S���]m�25=
%�D9�ss�{Z���7���N+���2Oa �M�S[r���zd��7��Ph#��{�i��,�tQs"��nn�c���}�ܛ�i��y\p���<wj2�njV�f󠷣(%��M�5�1W�Wt����vo�W�rSW�5�=�����jOc��M���sfe�*�U�X�1}I*���~����Юuщ�1	�Ǣ9#���y��B*�-'��=��yZv�mg[N�,a�6�my��׆~�?
�Tͣf����Ww���~z�4T�6�����g܋Ō&-�]y���5aK^Rf�G�3ؘ��mv���W�n3�y��>�iߔ�����j�����V۔�[pN�Z��O�}8]�>��(�u'�m�	��j��n��S�Y����
���g-��Ɍ�q�
�Aީs>}c
C
q���o��qZ�6a��疸ϵ��=A��x'�����Wpb2��M邁,_s��-ٵ�	C�5�o����{l���#a��D�P̺���k�ܕ���H�մVS3��?L�n0��#8��0�6﹁�ز�*<:�4�m������K�j�l��y�`�����b������]�(��s!0������u���}�44�O{n�X��s��&k�|�'�F�
^�aE�B�rN����y�(�xI]�;+�T17��a���am&�ߊ���l�u�?�YC�����7y1]P�ʖ��Xi��au}A�l�������8l�w0��^Gy7��b�Z�h��B�ہ<�5U��틉���9�{�u�.O���,G7v8�[٣�J5��^�5�iW6�n�c̽�~�̊�O)�9�aO�auF�`E���z�bu絇��	�������ͷ��;P���WJ;�1�ek��F����u��cz6)���.rOC��T�4�lc�X��6D-�����{�n{fxw���f����q��SKsA�6���k�y�IJ};;�u��6�]Q�%]ק^��ܶ��Y���9�n�ޖ
�{�Q�y�w`���T��Fb6�Y~�N�{I�]�W��-��b�%�� ��r�o��y;�XJE�̝Uͬ����{A����֍�l���М2��
�B�&Ll�pG�v�Tvu�w�z���8A����L�}�:T��H"I�,��0A��Ͼ%�9x�@�n������S�I�Pu
ڳ'�Jf'ǵ�۾��g��ػ�<�Ψ�����U�Rg�j����= ���\�,O���׵�>�oŵ�-}i^m���b�^ ���
�S8��B����1�R��Ofo���휪q�G�ۖ���O�u��]m�IWSl������i�<⯫˰����oF�w#fU�x�:�oǴBW�/�QZ�R�-���kh&�Ļt���hٻ�CKǚ/3�KA�rﮭ��R� ��aoT��=0Ԣ�����5���յj���:�n�S��B����7�P���w�r�:�j�K{��t��Npʞx��wiv0�ͫl[^|��[�j5�;�W��m�$����A��etD�槙��W��{�^�M�S�r�p]>��,����ř��9��g%K��X;�ób��A���;P�T��(�c���>�Sn'fx��{����&��t���r��rb�M���,dǬ]L�$.��m6����D��1y6�R��*S��]�S���[�Y��"��V���KC�*���[|�w�m�M>�+�a
�.�ѾYβ�n2���y�6��4餞A�zȫSٵY�i9�$y-s�8hCc±^��&���W��
��!�#�Kܠ;�坯mT���O�f��qCo�֡�pi�xo#���y�Y�ҩ�[�=])Q��,D;s�v��-�
��߻XSV�m'�A���O�2ˢb�����9����3}�8g��]zz.�!��7�u>����ˆ�]im	��7Kmz;W��G�,�ɩ�bOte�5�;
e�v�G*ݰ��t�d�B�(��m-/��׽�3�%��,H�J(i���u�v����e�N��Y0�}�R�I�����8��<!����W$�睷��^K�*x�;6b'��yg7�Q�"k]�ʣ���=���V�s�Ϲ�ڿy�ņ��{��h����{[���U�y\)�؍����`ɓ����F7�qB������l�Ţ�V2��[�X7{�9e<�4�R��kfɈ���[9�:K���}�,��X�-�G��8no7��WO��OW����.�+��W�S�J0pCk���IM�wzKX��WS�L��ނ�4 D���t�#�&�x�=��/>�v��r��m�6݁
|���wC���\�ч3����ru������h�󕵸����t���S��T�ovV�N�U��Jbeĵ#�݁�v'�7�5�{��=�n��b�s�_l�v����m/E�+ײ#����V����ތ�M+��\	3՘U�D��Y׷/j��Io2h|�f�:~������7�yoFPK�ץ�F0��qf��ř��b�q���U��0|�1��{�L��9E����ޢ�sʦ��q)���\�]����U~6��o���{�2�.���ޭ���.�V��sM�@7�C^\t����9q��Jc.'�yk�d�r�t���n��c��^�Zà-�]y�ݚA�z�J'W�{��$BM�S^�V��.+)Oj�zWfyY��Or�k-�=g޼��\A�M�5��<�[`�iԍ���c �r�����Ȫ�{`�1:���LD�l!��uA���z�7�1����A.���c[������������h�K�X�@S%:����J����/~����*��o�������@��ȝ	ė��}�G�@����xI���|;�p�VG#:x(��76:^k�|�F\o��oԍ���
��%̃�>�C��5��n���kt�>���c;R�:oo�V��x�D�7�B{*�>���4,���S���#{��Ln�в�U��[m��O(��ۇ�b62'�t�%�&��NrML�'U{j��JtM�0���&��*�z*;R7l��}q5+3�*�Y�D5�o��*[5���Mm�au[�\�m����ؽ�	K�{c�^����#�W�R��@��b�޻ъ�H�:�!�tuV:*�c�=,�0����Vj�L6���^Af��}Ow_�vq�m�m<��x̹�aOL.�� �3��y0"T��vhY(��{T靥�����j�Wą+��<�6�����C"'j�f�y���:Ly29v��Q(�^�5��Ad�x�L�CN�&uݼ/}ʴN�\�R:���.�oi;�Gk�y����Y�s�[�P lp�{:<�w�&B�\�j@m:���)}*��ws�C�L�����z����/m�N�
L6\�2/�P���O4�lc��F&u�9g%,�x�q�x��;xz�w�����x�$�V0�lm�o�e
U����]w���\#��j�L�B溩Y��8��r�{Yܜ�-a���x&!D��/C���s�|'�{�����Y�ڴ�k��Nv�}���zϏ���?�5�ٹ�_��h�NNx�����g��~B�;�_5�=��:���z�Xs)�s�{�����ɣ��3(�����WZbڪ�R�fk�h�1'Gm�ר��su���g�7�0��\���*Uk1w
U#u6n��b���;���Z�n8-M�;m9�W����3X5w,u%LI��ȇ'��v$��m U-T�io/��yc}��'����ku�������o�m+��!lF��	)9������y���,�삐�R˶�/E��`y]�HP����ԨQ�4	X���=�\�����DT9�5�;���p��y�|Cc��T���F��LK�O����\�/;<e��<�c�e]�P+4�|(c����g�Y�vo��k�M¦Z�Yc�v�k�ۛlL,^ސP1�#�k]&j��;��eE���Ԝʗ㼲�ƻ �3jی�t��B����ƜD).*d���7*���K_m��AּO2��+��9Q;˲3�,��y���Y��b
R�s��P[є&�o��v��o;d��f�>��I�=��P.�pohGA ��+npf��2��4}ᱍ]m:�o�<�5ښw�!���.'�Ѳ �Q� �ɡ<�s�os�~mTެ���r#U�gn��Ǵ���~<0��:�<��}��[��wV�#�\�Sʟdu#m8��<�[`=a�[B5;��f���-p�[�/3�pP�S'��ˊot��+�E1�����r�ֱ�k���<�4j�(̠<����}������׵�!�Rby�%�fr+=��<m�O>��kf�)�"A5���wT=�3�b7��R���p�5��0"lf���5�#��m��;�g*kxkB�QbY�oi�gXp[ngX��?����e��3��83�jG�knh/��.4E��0�ur�G�c=��,�޲Qַ�j���e��N�/PO��ݸO0�Y\�<nڹ��������!~q�0�"�(�i�A�.Mn��]}��������j�����]���z��=[H5`iad7�7�]�k+�M\aNT�չ����cin��x���v�lF�<�A�^��e�-t���H�i>�� ��'o���ؽ��o�:Ol������=F���#�c~�#]�l�����ok�is{�5k����i��1���5|z�g���ZNȞ@���:��y_��
���X�vk�o�)�n���*	�9y�EM�Lum#�����}��q]����pT�9<��{���(��(��Ώ��K6�}�P)lP���9u-���ҿC�n�08�m�]7����_��xo�ҝ�S�%ne�7�-���36�K�(vM�o�9��ӻ�	÷ET�|:�ڃ΄uϊ�4%�K/��f����r$nR>� o���&��+�B��y2v�����w����T���6�Ѣb�;v�ih��7�ք	|�=]K�(VP��IP{�g���٥=�ɩ_ 1�]��������Q�4F�"��;�<���[�f�OA9ٶ�W���~���C�-v�:5mar9c�A����uwc��R=�x���V��*�s���Z��oi�}�|yF�_X��x�9�:�X_e;�>�U!�IڻB��n�:���!�U������Z(���P�ќ�����B9b����uNB�38{U��Ю��av��F�oS����;pWgi�/x*:��^���)��ީ�s0���W>{���M�V
kh��3h�ki��'��`�7����aG⼠�I�,���t6�.��\�t&nj��Ma�;R/���Ǹ���S�+5�#5��N�󣺧�-��w��_A���W���%��mԞ�HG`�ᥢ]=��7�e��0�+��^j@6�H���r��֑��*�3��/���қۓ-��w<�.<<h�+�X����MH�Rw�$��Yn\u	Ɋ�F��<Q�w�զ���Si𵶦R#��2�9[d�76�YO���aD=}�l(�	�!v1�>��.#)�װ� �s�]���yyC�a���4e���h:�a���_�>��( �Q7o��s�v 2_n�һ�[��16�m�Qv���L�`N־�qt�#��4�m��G'U�{���֗m`� &���T�̆F���Ze���7�K�x�n��ծ���%�f⏬���L�f�^��T�H�*�7���A;���Q8����Xb�W3l�3)��=j�C\;�	�U�v"�lHVb�� 쥷R����z�l ���S�-�SVQ���&y�l�V����*' ��Fо��:����)c'J�J�\w�]����Q�X�U:U���WHN6P��wh1o�튻�B;��=F��s7��N1���dp�!k�yJ)ҳ���L�їjW`w�g�Ox�5Ӳ4�7�R���r��wx\��CzPCo�)9�����(<�ӝv�}����M��1V����+����ڹ�#�1�}��*��/z�D�����5�����.貄6�O]^��(4�v���߻��k��c��MW�ŧn���N�k��-gT7����7���w[7n�t�7je���U�	@V���]
0<��-�Yw<5ba�9�,�Ba�v�;z,e`c��Ѳ�O�;���-���;u�C Ԍ�F� �zi����y8��ht�W�JCL�Yg`|袲©��u���n��1� x�O�*T�1�Vm3 �f8 ��8B�_wM7{h��6�vsܦ'�et�17��/����]]K��1e�Y	x��ťd(�բ��"
�\m�f���	�Z��4w��&MUzi*t޵����
�bj�v/@ޮTz�s�WbΚ}GV�e菞t�}��>�G�,X���hC!�].���;��WeAFѨ�J-&66��ܤ�ݍ�Di�×s�3�st��K��wX��v�;���0wu�Dgv�YMv�$R�5˖�W.���JMs��nk���ѩ5�n�sd�K\�8�r�h9��,\H��
���;�5�]�nYݍt.]"����;ͮX����.�u��nl�r�M��+r��;�wv.s�$�`{�"A�v�2Rua64*Mu�ά4w����â.�tG���w��k�{+�5�wo��Յܵ4x�G�3Ƶ�dS���I��ɑ��B��T�N%�10!X���O(ًZ$U�g���T֕3ҩ��-��WM�I����m���<�׆$k������fz�/�R�u�}e{k<���?E'��u���^�ZÛs���{�6U@�͚kN�����Oב��z36��ȼ�н��L����������D��s+n/����71�
��q�@s�x��s��q�0�>�|�\��CJ �ʅ���X����k����5ij��-�qʰ�����8���e�։�[n�����Pi77�{3S�Y�v�8�b5J�'g�愵s�{�ĩ����	\l��Q��K,��<�W���S�xe_�iG���L���o��:G���r�Z�z[���ag&��W�$kSHlX.�"�t]LKq>yr�$��]P�Rٯ�Xj�adl"����jX��([��gf��A���u�Z\uֻ�K`�FQ�8o\{\�o�7���pvH�_@d��TT��/z�1�D�ɬV���'e�,��00D9�}��}Ũ<�˂ȧΠ8&�V^�Ϋ�>W�jܫ��]�����em�����qP�/oI@�	8�	u�]~T�kž�)K���t��K.��\3hZq��.��aO{z|D��B}w�r��pl�e���_wd۳�VΤíi��?&�h:�4�#�W�`�}7�;o���Wg�|s�[�μ��+ܹ��7���V!؟)G��<���bV�=Չ�6�[�3,��%<�������4�ߙc�X'�ыێXԙ��ʪ9KC�w�Dv�B���̱-d��[]�]��M,a�y�5��*pv{�zo��G�L��/>��GΎǜ�\��I�h�R���M���*��O�����{x�����ݞ@����Ϧե��!9�t�zi��m0����I���~���g��I���Ѻ���_�17������m�g���m�;��QLo!#-�je7��W79��{�Vr�FeoK2�-v$C�}-�y��JX��j��,����ל�&��r��i��*3t�7�B2%�"-�##�3�k���|��Ŏ)�[#�t��.�{Ի��%h�)���罵}0����k�]8^�t�E篃Y5A�gp�H^Lq�Ѝhʦ�%��ee�S�T�Ia��1�zuu���k�&{�j�:aW;^�ޞ8�����s�q��]J����V4�W�-���:K�u�h��L�[=����6�e����au[�R�ė��
Z�pc�K���A�i��E_\��\w6��=Y;�˾V"�J؍�����Nza �T�X]��W��%�	��cPolch|���� ^ޒ��wD�v�~3�7�7�o2��
�ݱ���O��,k��ζ�*]$&��`�ӹ���Fd;H35*jwb9����m+�z�<Ȧ�ߝS��fצ-���u�71tR�"�dF󛗫,G$���>��;�E ���
Q�i]E��oj���h�Q�A�6,��	[�C7���s�ޗ�t����Æf�}!���^��J��ǒ�����{~�psX'�/��'��?.���'�+'^�φדh{�V�7W�p4{oB�Y�z@��)��^�,�]�jԶ����U�
٘�[p�-X���oz�^���ojgydg��I�C5a�-
���c�Yֳze�C[�9� m0RR:/��{��[0a.��)�����R��v�E礞�����xb}�8Z܇l�^��^� �����r��)畧oroXi�ߖ�����Uvn����Z����	��$�hZ�j��������:����g��{���^8�� ��K�rZ/�Q˳+��gW�BkX�{^{#/9	��~
e�sŽ᪷o˷�(s�4w`SP��3�k���w�Nc��j+#�7,�/���Q���Y����Vd, �{�M'�G��M~P���Ŵ8�7��M{��,z�iz���e�D���7{%l˞D9�ߝv�:��b69�T$��@���sC�W%�q<}{6�խ`in*�o,&�[��ʾ��T�F�+w#������ɋW���:���3�7��V�:�}��NSޔ�]�oe������p��z����w@I=�]ARل��<k�k��-�kvk&��	B�\*̛�xzA��;N��k񠎖�6�:Cg'N���BX>�{���f�Hܹ}�C�4M9���l^r����c=��޻��s*�٨�[�P�7�����8�����=�,�[��{�U2���e���X���^��O:R��	]����߫ٲxOb���q]���>�����妐��:-r���<e��ϲ�~Q�u�j߻k������j�Nr˩����<3���
K�/y+��y���.ᆞ
�4�)�]@F�'0�4���w=���{�5g�w�m�4!ۇhؕJ$u#�9��k�^�R�P�g!��2)���}O�ڑá�����8��5�C5щ�-h�<r2�#5P<�jrfe�k2u������V+IԬa�y�#y��0l�3�ܕ��r�~�����Z�I7������˪��߹K�Xsnb�fa���sUn��rw��:���b���#�.U^����=��{��ۋ�͐�r��1���-t�t���|H:�ih��ۇ	뎐B�Lf�I;����d泳�FX�ߺCS�j�������B��%�T�儭��R�guc�;�[��NS��)��.�u\j��5�iկ	<�ŵ��xvꧥ�0�w}��
�s;�6+��,.�����7�dX	|n%�^Y;�|��O5�2��9��.�\��ڋ�|/�����G���!���ʌ��u��m��Q}Z��~��sM�t��U۩ڽ��N;��\�lE��ˢ�$�h�7��5��t���+ւYm���\��U��*�u��MY\���zb-��>��	/��T�*R�io,c��[A4�n�{2�ӽ�3�Y�*���\)�؇T>F��J�ғơ�6��W'yv���=�;�-T�o۝A�lL,^ބ+Г��We.R�(�co{�c�e^�Uc�R�k-���WmM���᝙d�X��H�AإIhm�������Ϭ��u�8�7�_�ߓ�������
�L�*�:�R�s9*X�O,��z2�sW�;�jt3�Q�(�C�*��e���vfl��主�s�ץ�M�� �C��T�Ӈl������&���|�oj�+�����(B7GV�2�Nb��[jg�0���
�q��
�n6ਁ�B��7Ҿ��c�_�	+��>������m��b���/��;���M=��l���'T�p�hKQƼ����+'Y��}�cR&��D?��V���X�wբ�a�T�롂"�!uput8�;�����7$Z�g���5������}mY�m��K~���}'2��{���)�}��C��,��k
m�9�oj��׵�Ho�Fb�6���o�t$}[*����d�燵d^�_"U�Q�����¾7�]����wwC[�j�(���b��`�k�$�S�#���fw�k�k�}�m�C��ia�-�T��&k:�p����:Q[�}]�_�M�:��r��N��~W���4s�-�ZjY�4룝xr �s��	_��V0��޺o�D�W���8oJ�fW3��!�s7��"�_	�s�MH�J᥼ѹ7!��}�a굳G�e��c��[���W���� -��B�>Fz+�<gi�z,�>Ƕ95����/��큨5��am[��۱
|��'��7D�f�X�cor��6��Ou��>�-�_,k�c6����+P���x�'�*y�X�ҜI/��9&e%�h��o@r�ذS��^�M]�H�<���0/瓧���ͻp�~]�)����*�[�e�ەm{�½��k�`�R�؝�0s��ޞ{{�ґ�*�)N�\@�i<�B*�om����۫�eЬ���WuM�,�$�v�~�]K_l6��z�݊�e:�=j��1յ�WUqu��c��׳��>)�Е�.9%���W�o���Pˋ<X��=���m^3zOZx���F��Z䭹��t�Is��ؘ����m��ݛX�;#��b�R��ኁ�:���ӽ�Y����<·=[:�J�̞`g:���&ƻ�3t5���E���=���zܳ{���O9c/��������a'Z��*��ʡ�ָ�k��SS��(E��Yt��d�r�T������c�s��X��k���*�x�#�݌�ج�t�7��=C�>��>b��/��@8߾��u���k�
܇��Yqz�����;���$������ӷ-�޸����(�Mű�]�ky��c1gl���}������)�d*�Aޠ%�PH5������C,�r�*R�;�[�yG��-Ł��w�ֽ�|��g�3�jY���� 9ŋEݻ�Q>�Ÿv��)E��t��O����r���Y����.��-x��v�H�8pf�-b�Þ%!���.�z�Z�	m�J�*bK
w_[�&���3VK�8��m����k{;Э����:�>ᆇ[��W9;��hf�6�Uu�n([��6��'�U��*r#4���>���f��V��FL�'�̞���-7�5��Y�4�n�dY�&3Z��j��;��*�X45!s���R�a'lsƻ5�ڷѝ;`��!
��eε8�u��Q���@�[��v'Ɓo�����)"#.�d�We�6���u2�-E��eD.��RدB�w����sQ�H���0�F���)�7ou�:�y2)7��t�aH�]Q�AO��ndg>�r!S��9��iFuS�v��Q�ϙ���aӇ��R���ڃ=�Wjbf��<�}$�̙����7�k������^m�w
��]�r���-�n�3:a��B�1]���cumx.�V�����4b6��*r����w���[���2�*@�C�^�BЏ;�<��Xd��R��������H�\�//���ǽR}��oP>�q�N�b��*�\�vK�r�3��&6;Eoe^݁�sv�;�f��Z����ڗ3����Rv� 3V+��B���s�su	u�]z��υ�=NT#t�y�o�y�)<��^5;<���^��[�R*sn�ᓞf-b�ͻ~)n� ꖳ�3�����9Z?)�/;�ՔP~;�g�yQ{k ��&����^�k�=��Dy�v�D=|�Q[|4����{\X�N���w�k�j�~��C<�!o8̠
����T��K�.��p̝�7��Յ8曅�M�]����ô)�q��G9�k�4w�_�m�����_a!�{�R������ߊ��{15����UELI��Y��:�ݳ.V�j��o/���agf��3�Ϡ��-���Nk�9O��A����Q*����uC�Kf�Ry�'xj|;]��u�ܚж����7M�T)�ЅGw����zL^��i���޴�sO`Gr�y8V�q1�@[q��.�Q{z|CIگ�'�B�xd��2.Ώ�c����sܗQ'[�x���#ζ-�m���xR�ۧK8�B	�0��x��d��Uz��m��O?&���d {3,؄0zֵ���ǉ��^��O.�g_p�{�*Lq�ko���P����U�vf��� r����$�t�v4�٦&鹪G���|.��wh��qp�ⲵ�e��{ð;b��ʇmm]>���st�k�suv�C�g[İZ}�
m�;�[z)�ӭз�ҧ�+�"\�bZ�����[f(�� ��W�;Cf�Zː�g4c��5���L�� �¸�%�;'�Œ�r�-�"Ƽ�Bڹt�"�!�{s�T{��c�A{/vཀ�
��� �)���ye4�N�X� ��-��u[��v�Z��&۶0i��hM���N�'ͫ@��F�6�e/a�r�>�./�z�7���**�Q�3�͏b/��Oݗ&Y��E�$<�͂t����Ok2���i)m�ۙ��Q]�7q�͵/	�+��x� �j��cmp�Rø�)5�}�mr���:�m
9��Fk��Xv����eޮ�':;�ǉ:��C�sm�\���-�6g`�`I�U�N�ڽ���;` "�"��������Խ2P�g(mt�%��5|��^�D�gL��'��0.���]E�%rά�`QS\����2˼�l�}kq�nM���J@/B��b�Ǵ�`�){h��ӅqY�����\r��p�dPy�)�)e�Vz���T�Ґ��sn+�
�֪ĥ˲����&@7:l/3n=�u��:�g�p	�plu9�̶�:����u�JS}�Θ�,���@pr�ܺ���l΂�nS9�3�P!���Q^�Y�?A+���ɲ�m�LȝA#��D�J���CɶV��*����g�$��X�݄���92�֘�������ؕ�끼�Gkz�|2�f`{kcȟb^�� �rq月k��EK=�7sпK��݇
��n;|��S`����ռw�*�z\�,s6�ǰ1�·6��$�xt��8Ʈs�}p��o�Z��O5v��3po/#pi]�4)K�ڸ>����.�I����i#�v>W�>=y˔��d��8��9їk�n��k>�m��t
�(�t�b�W|�09i� ʲ��W-�,OE���g�j[�8�@���yםy�-����\h|�K9.j�ήb�(Me��@���OV�$��«i���f։rۆ�P�VC}ѓ{�Ž�bCWրV8��ڒ�ds:��e�ҰM���|B8�U���	�0d��,�렸����i�m`�e� ���Z����e7�+T�+	�"�4%θ�Ž�o|�R���-�aX.l<�ks��p��YI�$9�ML��`�u���2�˽0�Y�+7�S�u����n��=,Dq=��2���2��p�)�SR7daX�_v"�\�MWlvfgҹ��F7�M�ޥ<L �D "�x���ksn�W#'wss�5&��sk�1d5�h��Ѯ\�5wu�Γ���Fe�\�颹sF�sF��v���C�r��ݦEp܊4��j4RW4��\�����nɮ�عs�j71t�.Wwnr��-&B�u��\���7+���7wh�r���3��.��*�pѹ].S�r7Gv(��+���;��\�:�6�.��sn��9r�7M�p��Q��E$��	ӕ����r�.],st����nE�4A�_Q}@��_Q������\T�Z��q����K�l�5�uM�(cw��5�n�u
��V"�ն��У\x�ŵ�|F�0*���E�:�+������owX4��i3�n6��sHt���V�a=���۵����'���ދ寜7��C�:�wR'��7��"��d�;v�����+һ&���.P龩�sN�-�Yǣ&wjA�*�8�Wt���� ��V4�O,K�~^��ۈ��)�pV��Ec۫ǋj�z��Fdk��q��Q�"�s�������Nƨz�u���O9���зH�^�޸�Oz2����]z�T��\����Q{���YJ+7����.��ֹ���mh�{�̨)�8���]t�=X�� �^���IN2�r춝�2��8����^��6�Z��i�������z�s�,�;|�/O�~"�RѰ��|m�����ał��k��K:��@WGur �s�6�J��V0�Sxu�N��C/U�yc6Jh��TCx���:�5Ȯ5��T�ceU����M��R�w�M	�x�P�2�=X��I��^����1:��aB��Ӱ�����A�%�r�d��`����m\A� ��g!]�(�:�b�-p�8��I\�&,=�U�iq�%�/P��;;���DFl�R��K7C�B�'�8�k�������o�:Ol�A
s/����K�}o�U4�(Y���jkv���6���7��5�1���g9��*�oIB&���U�ȍp�m�	�j!�L0#7�]7`:}4[����mzی�.��"�[�N^ɹ��H�h��k:^�~��DU��S������e��C�{���[q��v�1�R������vl'<��蠟{Bs��~F��*[ќ�J�g�57��T�͝�Տ.T?^�H�g{�R���	[�^��v��l+Y������ܡ5繉w�3:��;�"��f�N�n|V�Оy!ĉf^�{������{OdȽQ���v�,N%61�4��1<��-mz�Ťa�19W|_i-�9FJ���N��ubI�r�ж�m�^�O6K��ݒPʶn��%��N�w����VX�9��JV++��/"9�v��R��FF�9-�t(3qz^O:�S�5~�	2��m��胐�+T/����Ӹ�:6m����=�vx���^��6�Nv,�!��yF�+�,�\
�8l��L�����O���"�s�[�o��w�r�k�uCU5�-�n,v�rw��ۍ���fP-�f:�������3��Ɲ��^E�z�Y��F����ګv�m�7�4����C�zr�8����M�87v�d"���B�����v�CX��mwX�Y�v��e�F��K��A�)*�!Ô*��WSC��I�����o�b���hV�ls�A�5�\(�F�3x��Jak��T�W᥸�a�����t��*�u��Vŵ�xn�Z��ŗޱ�^������^���{z�Yx��	���6ނ��
�о2]��j��K�\FH<.�����R٠Ry|��/1҈U$jw�7�ڙ[j+.s���H����%�B9�ߣ�W�'�����㾔��Zg;k�u*��L.���B]#AS�\W�[!k��\�GMk%�8�ĭ��P��1o$4��k����}���C'yh��}�[�ة�����q�9��QȲ�l9�O\y�����3�a_U�SO���3�	����v�m��1V����n����ɽH�+�t��l\Q{X�'�y�D�Z���jN�޷�dW�oL�F���`4{ڔ�B�EC݀=s���õg*���[є�i7���v�!R����P;�<�Jy�\�3�t�۞�RL���y43���p���Mi��lk��5���ծ�˵�J�٫��;թە��,FwT+�WfX�ogug.�I9�l)Iǳ4�7JX�9ՓnV��Wi��7�=r����7����K��;<��(��>�D%�S͂_�2�����yn��Җ���߭.���h���uv�����oK���B鼜�6e�Xi�Y樿2�����8ח,8���aD�Ob*��k�k:����'�ϝ�)���t?{�!���
z�C�j!�g.��zy���Q
b�ʝ0��d'��R��v��yv����2�^_���c��so�n`�T��'PJ�l�YJ(Z	e��������G`�AL�Pl�Jz�
��v�.�z�l^E}=�&�*9�6�]�N�� ~�U�>�v���Ĉ=�*3O��f�B�6�xM����Ww�8<+w\�ĨGi@39�7+>rw��X��u	/d�4'�/Mn޾͌Cvc�ݪv�S��?;��뗝�UlF�JDF;�mS�aZ�z[�����%�f�����wX��o۝�`��~��+b:|W�#	wz���
�˫����8'e��v�!;��Ж1�-�o�)�n�H^ޟ$�%˻6魺N�b�b=������O��[�L^p��*]#^F�����4i����mt�f�oSEC�j��{�Iw�c9�A7N�ʈQ��݃�u`�Ul<�(�0���>;�j^���-����_���b�W�5i�^�Jo���&�x���F܂��J��N�(t�T�4���TIS(oTGne�ӌuc��X�f	���k�����;�ȕ����3�z�i�������z���^�]B���}΀Ui�K�f�F���Y;_����_���c�~�]o�����6A� ���g�ו�����q�:�Z�GJ������g.6X<h������EP��ь�+J�W���)sXk�J�m�8��u �۷�{�o��@)�1ط:�s�-`-b�P��R����[�	_�P������]�Ɩb��=��Ĭ_m���G��n�b��h�y&)�7A����F���.���&���S^m"��Oz�k�?u��ٽ�i���n3m\5&^�n+�^�wpv���i�q�qşO�P>�a]���\]�p.p99'��;H�g���k!�UI����_�i��g
�e�I����x�ku���>.0�>����%qBpϏ�U �Fӈ�N�SΜ�t��[�Cm���wϲpl����������_=�	��&aa�;P��W�TYj�>�nț�����T��>��6��9ޞvW��7"V_]ꑷs��5y�zag�e��*���rx��Z��������\��z]?�)�g��}9�1���(JG���P�B�����e�K�^�+���>�%�+ub�R��s\�V��9������^@6
4����S�۲�q]���yu��}kB~����qc��8��
-���q�Fw����ӻFCTA�ћ�]h��.�5 � k�=�. �}9�@�C���"[V�Ay���:�&7 ��x�{�ӕr�fS�e�[���%�|'I���[F����GL$��F��}P�`��Z?\&\�Nut��!n�XZ;�/�oyQ�L����=���xbpq=�P��v�x�)�͡/���y-���j��fs�#X���G�GZs��E�ì�Z���F�Z/v��!��#BjI�oR�tu�7n�QκO��d{����ֻS{˓�����D�N��wQ
e���!"4��/k�̦}��6W~;���T|�����1�5s�c�o[�6�x0�)��J'�A�L����)?(p��5;i�fމ���x���S�o_��]wF���4n!7@kBd_�e�d��0�M�4��O�+�u���G^f�2�'R��{��f�-7��!'w�1k�tn1�o�n�f�K�-��	�r����ZJ��Ȣ�����}�I��;��םw��s��\�s��u`��q�b0�]F�z붳�:��.�f��������[YOM�J��u�}~j�ϕS�c����=�������x��`le�=�ִ����«��j�ϝ���VW -M'���F��59�5tv�d�!Ϻ�);��֧<Δ%�R��vOX���be�f:\��˙��{(R�V9ş/(�5�\l�q��|�2��������k؅��:.�I;_L�o��[�ٽ�.�W��f���"�yLO9έuadit��t~9�r��j��S|w�{�Qw��z��o����ڷ�2��ù0��w]�b�@������N+�C[SB7�&.�Rs�֔����8��u�nk�਎��U��e�qM��p̮v-g�iM���]�*;	�O�o5qA�2���|:�R^�:��r��S�y��Z�WZ��rN_l����c�ʱ�_�.�_ѷu<o���_�;cF}�!���j�㷛���L�l�7��o<c��E$�A��E�r�O]LK�V�E�����蚱��3����V�����XGo����8�Y����T�"Ku��+�=
�F���Hqx��ܭ1�W~q�����Ӕ��7\4�nH����jd�� ]!�7�J�
�A��g�F7ۺ⧹����M�޷�/��c*�. ��-�A~�&��E���O$O����u9�(�9L~=�X{�=3�Щ8������G��rn�Ĳ�KBl5ą�*v}CTy��)zi�f��R���V����)��J��rCKj��杚6ܸ�*��[t�Ӧ���.��nx�Y�]�J�#�DJ�(z~[{ۯ��wS��5w��wt.�S.���0܎sB�=B�?R@y��b���(��0�0�u:���������Y��c��7Ֆ��qט��t��u`��^�yR2�<O��9	�;����2��5h9ǶA��j��D�-v��2�Թ����:��!�/��Ek3\�kq�X7�v�YF�]u��B�wk'`��yvQ&nK���xJ�ٻ)�|wR�� �:�=�4������#����s"�F'�r[]�t_2�z�c+J�]�,ˈ�V7��N�o��iǧ�g����{hd:�~'����5u��٢�NIˈ�`���ea���Z묩�"z��|}u���&�5=���.�.�x�i2��>��V�vS�x?d�ů���5����6�m��]��4�S�2���t|."��]9��X੃��2�ϝ�gr����d,��Q���}�;Fu�ޙ�D���yٔ2�t�qS/�֪��l��
P"�)ቺl���"�[�Zb|d�~��C�����Pz�Wr��!4�&j�!q3�on�X�e�Y����?7���oM��s�Nfvh����:<��pݠ���++���Q�GI=Fa@�Q��d_]�e?F�o��֣{q��Ԛ�qG�]���KS��� ��>�=7v���T��5%!*`�rX􋾻U�/�3���T�vM��[늸���S���'#�n1�#�N���2
5�F��f�#�i[��Wnb�΀�qT��`�38��p���dJv��/6�,��v!7pv�ݳC��I1ը箉�k������<]ԑ�c����M�:ϲ t��oY��u����8\�%"w�'A��Fho��c��A{q��v�,F&�A�>xug��.����i��,�br�#��q��M���z��e����q��-��V�ǥe�o�����;؍r2���.Qe$�zqGk/ �)c�.�za�ܭ�e#n��/�J���:��PJ�z�b�m:7Ew���u ����a����~�IH���矽�׸�z�O���<�T`�N�A���N�2�/**V׼ds9[��[n��6ˡJ�⪳'��j�~t�n�^|�ЭyR}���i�������sQ�Oދ=���Q�/��7�~�������@:7��,_霸�`񨃒�E���q������Hv��c����x�TfڸjL�1���s+�k����՚w�m�T`��������Y����>�V�fy��C����EJ�O�=Ԁ�cYb�O.���7V7eϣ��Q�r\rO�X���g��W2��x�xW�C��k��P���B(N��\���Dh�i�8�_g�X�<|�6�i�O��ݓ:v�'�Vs�;P�"�W�TZ&C
�rחфMD�:��1�5��F���|�P\��7%e�ީ\�'M}'��=P���4�˘��'qӝ�q�z�5�	�v����K���C/�w��;T��J��Y+�B����@w�IgF��&#^vlO��F�)yo}xֻ:]	j�׳]Nط�CL�Y,�5�8�\����!�ʺ��sH�3�VOU������㾺�y�_�Q�.K��w��;��%����E�4dѻ���.��3��ח)�<���Gd��=��z�t���+�ӻG�=ӌ.���o��Kow���a'�b8����L�`�ꙶ���g�8�]d���.=��^U�� A]NM	^�4�k{�C�t=�1c̺J+�&y��v-��c�:�K�b_B�l�/�%ȗY�n���)Ep�ң��ř +Ϯ*n���]�	�Tg��s��O1fZ�*V.vZ�,@J'>�2����증mN�st�]�,�Z�&��薻�:�S��ɽ��ޙ0

�ؤ�u@�Ӷ�fA��2i��Q�(��E����D�����@	Lټ1���`�� ��N�y0m1�[�3y�d�E�=�]Iɶ��3q�޳A�\���@\��}���,����#�6�h��=���4���R�VL�Z�7�����F��v]j`*��̤p���L�b�>�=�U���O�'P�0���p����q׋zF��g��&64һ{���S�;j	��X��eh2�+�1 h��2���������B�E�����{(���:b!et�<g���R��@�*Yb�A��ޮ��{{���;R�S��������nX�mu ��C��q��D�V�����������}��<�ũj5;,ye^�Z�;�-ɾ�˸r�#2Ʉ��sK,c��2���M���|)� �k��)���ZH4��ab^mHK�ɫN,U�q����CjN��F�9�[�$����T=�x�O{t��ϡ쮢��1OeU���rv��B/c��F�P>�q�O��/ky�����8�;���M�L��yolS�%xN.+���nh�k��ɕ+������܈��N궢�ș8��r�[.�t�2F<���c�]��'.��ln��/��FC�f����ˏ'�&�w����w9Y��+���ΧJ|d��i���^5юCB��=Fv'"
SPUm#2��ŻU��wI.��]v�7q��uۿ+l�QRk�sپ%�,���)������q ��W�N�m��N�e]�r��R���=��ݓU��-A5�1��%,g8um 7�0��cX�����:��`�ћ�ѐgْϣ����5����V�]c"ٜS�	=s�[�c�X�йZӧ,m�Q4+(C�E��S�jPr���.}֮\N�ǴDx���xVu���N.�2��4�G�-�X������9n�U��3�f�;�s��S4�旋Z�o�F���4�ɚ��]�Ѻ|��,�%|U�7=2��Oz5�����d����'E�a�{i����7Y����>���Ԡ� 0�G�DQ�9t\(�+�;:�w:N�Ѻ]�s�͹�'ur���Wq��w\�wn�A�4�s�rPsu��t��wN���'u�ܸ���2n�r�7.W8*w[��twv���B\�Msn�ݻ��7e��ݹB���]sA��F�rH���s��]�Ign���ܳ�$���Ns�;��7u�v��39s�s%ݸ�Q���uIc���X*r��]�I��t�Ĺ����w\��v�s��]v���ܮ\����I��#'wu�r�p���]�T9Ė5�Q�v]�\��s]����%$ˮ�˪�7wY.빸2�ȹ�Q�SEa�6̊7wE@W���� ����k�ʷ7{�ko�H��{.{.�V���{���$Z+���^�8��o*����.[X��<�۶m�,/^�]��v�19|0g�/�3�,WT�w�V��jT�z5�ei���>�Z��/��Fw�FxQ��C&g.�L֎͍up��ql	P05��t��n�Uķ|<2#���:�����>��]��Eu��[�u���=N������Kd�'�N`�C���%�hd�lm���dW��۽R��Ƿ+ӤK����t�ؗ���<H+��3O��Pn��60.�T�Dl֖L��&y��e�h��N>p"m7^�v�&���(A�΃�be�}F�;A�n령ۮ�mҤ}N;���Ty��G�u���:`<�*�+�T���N�Jg��{�ڲ�x�ѥ5�L�)�)Q����nD6���/JdѸ���!��^L�HeJ.#1�
y��r��ռD.�h[8���z����KM�����I�酮%�X�@;m߬��=�T����Gc'��x~���Y]ƭ�pz"�V���H;ͻ�c>�Or1k��S�ySw�E�ߎ_Y�u�R����=0A:[Vea�s!U�ta�O����5����< s?z~w��2sQ�R�K�����ou-#N�ϡ�J�!aq�t�[��
��6�F�Iw1��i��J�	�R�N��n�J[Jů�l�i�S��:�t! 厧�
��7
�����gX�$C=�8�o���/���R��!�f�n���M*�S����9\�*Ck ����~��gS���*�M�--�\<Ley��^z��ߪe�J�ߓN�}9(OO]�VN}W/ 3V��M�u1���Uó������v����+ڎ��&F���\���A/x�۞���̸
�]2o�R�{���}q��Z�I�w�I�	��j�/��o%�ə���A?�ti{�G��R������e��r��v��U�\ĸ���f��t�r��XH)�e�0���S��j�x�:��U����t���#�~�s(���9(��Oe���Y�;>%�GI=FPq"�.R��캉w
�h�JN�3�{�8|}���κyt��.���*�|m�w>%�D@ި�0��I�y��P��/��
9e�ַ:mNMӉq;�F���Bu�I���#�N�	��2T�q .���"e*�\k[�=%Y���W:���@��}�S���*=|��r����~���~�V�ڙ%
�ƾ���!c+^J���dz�݁��qΘ������-�&3~K��L�%�͢SF�
Sh�(6�:8?T��O9����I��\NJ�m�r-��F��a~�������I1u+exp������a;��ݫ�{z.��sXT�w�qms}��l=��Aj��vs��}f�n-�ئ^�9L;Kcy7�[ǥ��+���m���k��-I��@�{!�����*\�ͱՂ��Q�S��u-=�Hm�U�ʍ�r�k�e�7��;Ԧ�)o��v�����d�N�d�lf
��OMg۴��.��Cwt=��JLX���xVb��[
���(���Ƽ��,��0�a��9���i}��cG<Z7�����٧W�/C�U=9]j�XS���Ջ���~�O�	�>�B���1N�J�vw⎫Z�+��l�7��Fm�cU?�Θ��5u�r��,��a�k3�s�I���������a�%ﲗ@RqJ�M���㞙P3�T>�<�'!\�{"W��;�>s>���Lb�������wU�4u�3�*΅qR��IRN�e�*�7�2��wM��}q���}�`�[�Vk�0ƭ��߬�R�e�T���g�lW:�^D�g���8tǘ�v|6�:<�f�OZ���87�������{�g��� �C��R�e#c��觏\e"B*�s���dWW��_�TKg��y�S��W:9��#���3
 }0�(�G�{�߭s�V�̉�����]���,LD�\ ��Lo+)ڕ[���Zb�38Ed:��;�x��7�8�t��;5vр+J6��;{j�B-<�.���U���Ҝ\��]̥N\��:%'�*
��a\ �:�-�����Ƨ=��y+����qW<���9N� ��>�=mݰ��|�� o'T��Z,�=�w��z�~��Դx���|z![늿�[��N3�S#��=t�ћS �,!^���e�/��+�WT0L��#�<@-�����o�� ���F�u�Ώ�wI������d6y�=]y94����4�O�|�H3�<�hJ:�h�aZ޲=q˭�2 ��Y�w�Ni�,]���zļY�S'>�m@u*H˓�"d/������F�����k������+��w.�����A�wS%�3,8U���x�w��Zo�/**V׼s�<ϩ�����Zv׶���ɭ��c����pm��6��W	�K�Fhf���,��������^��z5�h�r����(�E��Ҹ��o���x�-t���	���b���i`��z�]�nWK#�ov��A��Z�V�ߎ��l�o�n��͵p�T��n'Y�:�>q���O�oW��P�bկ�-�C����g��A���f0����WS�|$��s:P�k!�UI���Q��ڠ��]�i���O}VʿUyL��j�E_'�p���<�R�/��j퐥�Mȯ���4�i�4pN��=���p,�j5(���[�,��P�b~<�$<�T����n�e��v�ݭ�6�Xw9��a��)ٶ�=�R��������������U�>��fpБKC�{y?���O��(��?qd���YB_.�k��U �"�_g+@��q(uFM�fd��.��+�J7�}�ҋյ<lY�����xh��)s<v���k&��sO����r�Դ0k�KvE��M���0Ӫ�Ǌ���kjc��'��+�Hc(ق�J��lI�H�~�{�zC�.:�K6��������y�e�>�o�>v��ϥe�P,���'Ƽ��k�Lc��KJ���:�\EL�,e��F��j�U�V��!���#��>�[�9�e��{����f���o�U*tp@�Q��l���ˤ˧<+�[���q��;1KTX�����ǳ���g�w&�.���@r
[$\ϧ3���]p��Kj��ѫ���l��V;�NgZ˿>	���'�8eӨ��F���N�<�h��ʻ+ݿ�p\��q#����{8�F��l�h9����x�n�iL���BF�;$LJ�tT��;Y�ϼ�;����8�w���*=%���p� 1?���R�mL迌�e;�oA���lV=g�GWB��-���+��M�*���Y�Z��JO[��^���
ú*I*���Gq�m��`�v˒��%ލK�k�G�V}��A�G;�3�=/�C��T�],�p.�E�6��KUq�O�.�����{e>�d�����������3*��N����}G�_��=�xڻ�kҙ4nt�&E�y2^fUH틨��Η��:�x̌:5�8:�{������ݥ��]~�Y	;�1�\S�x�@:&�H�۞��7u��T�R��귈����qœ�&G��mK��U��n�6�Ξ�{`M�)T��,^�c�y�o��,Z�������B������u.��q{
�N�J��';�[9��CڧzCT���:��rmp��ȼ��O�faa��*�_қ����C���Ek�N��4��Y��7'��WN|���s�������:���;�C��������~����Uq�.G�f\x�d�r���Cˆ�c����k؅���tv'�ѕ�7�U_�k�I��L��	�qS/�.�P*n!k�>��q��/���g�������q�P�l8<���7�(��3���v��2�����ӥ9X�'LxyÞݤ�;��*w�Q�~5���}��汘x.J(i'�e?@=Ā�];�u�Z�6�U�� ���mFI���e�vq��?R `������pߪx�vr{"~&ryx�7w��߳�I����A�9�gL��B��6�\��k����,r\�\Z��->?"fHz�\�۰YC�mXͦƼ��� �˼��E��l�=h�o)����D�<�>^��z5��ۈ�\�t���B"�0�\�I�'��s��.���	�t-���q7�g�9O��:��ctG�)ݡ7�*x Hd����}5*�V���/t8Z��������Q�N�*����~�i��.���S$�o��z����ѹ�<z�=R�9$LO��������@�L��xTz�K�ɿ��ĳ�8�y��Gb��G_<�W��6H�;= ��c�}.u�N{ƽҼ{\��ڪ0�vh�dv>Ľމ΁�][�a���Ơg��FEF˳$�N�Ʌ�^��w��>��zk#v���XȱQ�$���6/w9E^_��s��7	� ����RF�'�L-�>񎸧^�Z_q���"��۟1�g^W�с�m���j��ϖ���c�
vrڱu�HˏJ'� �L�z�lIܚ͡�质�y��F��'t�/�<�m*c�U?�Θ��]D���}�-d䜿�X>>�4��sbڿ��=K�Y����N�x��~�}p�$�2�ϕ�G����vs��_D�-^g�:��w}�o��u`~鴁��)��A���NX:�5�Kgi�����:��z�Mq����H#j�|U.u�s���[�3��ͤZ'V�����"DB�&�!1t�6��ݯ����&+[X�����N
u�����P��RZ��p<�_�L��>�%�����ȗ�u�J��u*��������V����e��[>�^;�����{�v�Յ{%Ǳ��3�L�kL���J+��+O�i~���+"����ysۀN�<���R��χ8�G���Ug�]�n,�Pf ���3�on�Co��g{���sVЍq�����l�<��ӏ��/)C�%�g�*���H?*��|���:���9]vB
��9�v
7�ֶ�"R���5;��@-7�>�=mݰ��U|��7CJ�0�N�{����=�� n�/�4�{P�u�z
�g���㷍��uhγ�*���s���=j��P8��u����xfq���oW�N�1��m9��EI����N�̗�}�v��4���1u��І�z����A")ڀs���/{ޟv<��|Y��%�U�R���2�퉘�bwT��FB��{���T��OfUT��gM)�ڕS��Aǹ]ж�2^C2���
��'U ��(������s���x�I���������y����h,�8zd|F�R]��K�>�q��fv&��偊�nN:�e=�z�/��� tU������BAW�����]��jT�}Ԯ�vZ�����a�(�eN�R�%������#:9Ҽ����hQ�헓�'e�q�{=S>���x����7����mUѵ�@:��큥�3C.#_�A��d�@8��w�ۋ�ފ��R�*�;B2]��7[=�#�)|o�׶y?����F��!:߮��~��}L��A���q��������8�t�l����])i:wJeDf�\<�T��n'Y���;tw��&���U�f����8���|g�ϧİ�=>
�r�������H
�5��|���	���\��ʚ��{W���K8���V7r5���ו><9�½��qN����]a~�}�NO�{9T㛀>P�o%��KV }�:l�|�{Ky*���Q�)p2z�����vNwS�yc�~�R�{��	��_�-���M��!�0�;�nD����#h�'O��9vLaZ��qc��w}��ԗ���p%��F�O�<�2���p�N;T��Ҳ�,��S��uٯH�Q�,�^r	8�����u2���}tQ�V��\jV��k��ӑ�!�}p�:�GN��Bu��j{m珠P:z L�bO@���Ge�g��W-�����)
��>�U��Hq8�DВ2�	��ߙ9��ki���L��B�wv#�����z�g)�����Ń7�$"�ت`G'��dy��|qv_���L[u��-9�Wf�*֮�(yFQ��Ņ\�M#�6G�V�g�\	ٞ��I�F;s��]����ۖ5�v^[�(�m�`���΢�8�����مJ>������ s�������|8;1,T��]��niQ~�=�;C[�x��n��˧Q>�d��@]�N�<�h�����Nz�s���ڧH��^{�d`i5han����D�&��[�q4�\�\!#pvH��WC�-M9��=�N�;)Q���?m�f�!Q넺�M��:`8S`zR���ΏrQ��.��K=7�t�C��y��mX9偣��ҼWsۆڪ�н)�F�M������J���t���k��̗s�tv�
rԭ;������O���l6���\S��x��LR��b��G:��z�b}���6��Y*�$5b6����pN�zN����/d��g�o<��w�G_x��ó3֡���r��u`��߅���~Y;�d/�'t�9?q�T��;]p>���Xk����j�^ j�CS�#�>r���q��\.=�R2�Y>�!��~Tߢ�3K��j�_V9�y��4^����'r<i�+9+#��nJwQ��Δ,�5N����Ĩ� Dfɪ7�_�+�Xg[�ݬ�p*�Q��A9,����k��n���2(wy��틊зN��5�I	
v�]�nKeۗ��^��i���pu�s-\��d���z,��&�E�3b�^����F�f��N>����u���ֵ۲����:9����{���0�O��Zڧ;�
�K�/�M١ub�X���zX��i�
�F�j�W@����P��h9�xXU�ҥC^Z
��S�L7BA��9^
�]�A�юː��+-��AN��PWn��r]e6I=���1��|w��1҉].��u�*xJ&�kA��Ӎ�6漺��<�F��}��ܰ����;��1�i%��s/j.��F��D����ѵ�����E��ͣ��V>�C��w�ҵ)����a!vn�n���v,�I����jX�Ti	�����8/!�Ɵ����{�k!�=���ʰv�q��ߘ	��x��H�5�F�=�*��P��ݴ�{-���L�۫���0�"+ٽeS�I��g:�%���og�Pe�9����_Mȶ��Ӷ�6��̘5�Ņq��̨������o&�C(�����U�Js)V;�*�Wz!��K�۱=��^]7I��|LBP\���u���n�J������XﳫUmG�^:�/^�n��+� �2���8e��ڙ��v���*�n=ww���:��5 �&�ه�7�t�ͮ#��}hb���6� 	���R��lyRK+iĹ^�l�`�Hi	@r��9]�2H���F����3��:ç�|��"�������j�T7=���*�N������R�3��\G+V��E��C�Jz�7(P'K�Z�g*a���ȜYwA�٠�3���\r�-V���&N�.��3���=��%�<kt�}�_Y1�p��Bj9�mwq���ED.�9�7SǢ�f���bs7�Z 2b��͎���x@�6u����;"<ۻ�Y�݌Tj�Ƀ��dҹ0D3���2�����p\*lNTYQ�ڃ�>ܣ[s*�����C���ztSpc�ҡy��nZ��C�qA���Z������KU;k� N��7Dwf{���e���糍�-�*����V���t�)�_��j��Z;��)�s-ڱ�_\�|���v"?a1Bf��=��H�a	�{1q���wY	�ɻ/�=�,ˎj�����pP������.n(�-̭�|K��Up�)�[�U/�uaNZFpˠ0�ďx��bb���-y��;^Xu��Hg��b���.����6�t�P�0�٢���>��e:E!(�U��H��|�������*���!�sr֒!�X�Lr�zh���J�F��5X�\C�Զ�g�Ȃ}X5��0y�g
֩������R�d�ڛ��Y�ƍ�!��_��W���[�?r�i:gH<�y�<��1��|�4Ȧ�j���_uM��T��@�� R��&�܊��nv�D�s����]�f� �����b���A������$�H�	��؈����Ac��I��b�q&�i��0�0D��+��']fI$d�,(�B�DLk���L�t�!F��s&��bI��B�@ɠd�ZI4i�����E� �7З:G:��f-�`�,K#&�;�3,A��#LB,��2!Jad)����u����Jnn�˒9�w\��@ĉ��0RC�;���f��g8�2f�e�ь3��+�a0JY6�2#H�D��wn�_����������X��#�ZG݊w;4Ƶ���.���w����D[-֢�2ž��V=�O�zS�I>f�l�s�w�u���_��=0�S��Fܸ	%�]��Ȧ_��$uþ��ƽ�Ni�滩e�Ǻck{��J!ԛ"�$�_L�u&t9%�Ǣ�P*V����.�7��/�2�ޡ�h?o8�eїڮ}]��zⱝ�F��o�� �(�BOO��JW�X������Ȳ&�t�ձ\�4v�.5���mv�WqMc0��rQ�GI<
q#��]9�P\������{�G�E�^v����b��ԯ�"�4{�k���ñ۸y�_" oT|f ��9�ߜƯ+߄�ߩ�Q�hn��aTr7O�&���8c���S�&ے1ӻBmL�5@�{��[C�qR�2���7�sJ�0;��P���xT{���f�R.�xM߀.i���nz�Ou^S(�j�>^�*���I͛��D�:�RV��)��[£֗[�i��Y�.q��.���8�gB�T+��1�.m�:�Nό�5c�GY��s�5~�Zo�����
�{ŻD�^���k��gƎ�B5�"�ç�2MY=B2C�/Wһ���T��n������&�mN�3
U$�ue���d�eSCyn�c�̌��?z����-1^`��~��ÒOVo9����>y��;�h���W�~;g;��S9�ՉD�*"�=9G�b{r�{�jm�n�Ѐ�g��FP�9SԝG���HWm���|�]Z`�wg��+�B�����c��ǵ�з�A��7,��<,\k�H5,���L-���¸��l#��pf�7�ߟ�*g{:gR���7��e!�2�\-t�sAO�[ڱ�s"�҉�	��ܜ���h���@r)�q[O��L���l�ٶ��UT�Ns�9��WQ:�/F�����\��;�5~�=��n���&^����Օ^ $Oɕ���y
��,�C��{!��%���������	���*���L���9�X�'GeK��%H}8J{�[�9�e�ܢ[�S��/��ܜ�$ֽ����?��ԋߋ��2	D~�є2҆T��:�"����b�JjUof�dV׸v�zV��!�峪�G݅�"-��f��=�C��2����Gޔ���++�O���![�!c��O������y�o���"VW�$�H�'��(�e�������hʄ��]UV��R��̆���:i���G��a�6J���O<�B�tf=��*� ̹8�:�lg���X\r������AS���'#�o�<�"{�6� �g`�W�}lz�JA���k�
�����ahgȢr���=�{B{�h�e��-v�}��YGM9*�P��c�J�tS�Ś��#���>���m�j�lU|%M}.1�ʮ���Q�]��ڍX8kWs!�z:dw��L�%�8c	x����c?���a�Uޗ�@P��8
g�p+�-��;H�Ay��H+�ѷQBj��o�eb�t�{�pv����I!o@�"d��qJu��S�;���q�������߅�m��2ލw����J��2B�Q5eI�&9�Nን���Q]髾}/��O�=��G6��o��}O���U��}UC~橒�`y�W:�#����;���χ�����;���vZ�#��fT/�� �WF�y��;`ih���x�z����v'6�Nm摽k��,�N)׼n+���>6���9;�9��@:7Ȇ�,��4ݘy�lv�~�3�_�e<���:ǧ��e1�ZO���)���뇊���g7̭�1�}0�E���3��r�.yg����~���pͣ8n8����2����^����'��9�(�5��ｔ�]�����fd��.#n���W��j!xm�N�E��~2W�OȡqY5�u*�|��Ky�S3����9�r���A駌E:l�C���-�Z�����ĥfC��;��@쯱Wu��7��(���j��,_��6��$�F��3��	}�n[� r��a�;ڶOV�Wq"[�w����W&��؝;A��%ۧ�%��L uX�GF���0p�u�U�:"�;wٴ%ZsVU��R^]שX��c��&�`E^E:V�q�w�����m߹Ti�,��[)��<��w��*���Ɔȴ�����[#�0y%�f���M;���>�ۣ+��p%���it�s�9�g��}9�1�+/�Xz�о�ՉW��h)tM;��K��T�R�E��Fժ�W��9���9r���sM����2{�����U�٬���65
��,t�0Sî�2ݺ�W���RٟO���ʁ�t�wc9�]�^|��H����>�wh��rQ�� oW�@s ��E�O>��P�~�A͛��;�]7�rՌu+cͶ59�������u�fK4�W�x�>��uq!E�T����r�c�8�c�:����|��sĵ�D�n�÷q5�s=p���.�F����x�t|o�yI����.�ޢ��_��p�
�\%���h:`<�*�*R��>��d����ѥۿL���Tਕ��WR����+M�=�xڻ�qҙ4m7@kfÚ�����vn�����z}�]1Ǧ�䡷�u=㱴���ݗ���l6���${Y�F��K��w̮X$�������Jc��ż�={�a�,Wf)�6�/u�j~	 �'��9��ZY�*p��6��*+;ٸ6*w+�=z�Ce� ��B�c
hӆ��^��A�R� �m�#�JF�����h[��W�2fF�;V����n֞|�W����g��?w������OT�]c�ि��ZN�F� �u�
1Kr&[�����_��*�����{����<�Ճ�u���^T�O�s�xº�zyצʉ\�<��8{��[mn#z���1ʩރ����uc��϶�_�*F_K'���X(��M<�=�Y��)�:UZn"�S'�Ɛ�9+"��t����j���p�~����>ּnvD���]��S�����}1ΝW��P92�+�L����^���u���]9X�n��L��aͷa��Ib��I;Q(*:�L����U�ֺ��9`�c������0H���:�a�X��G~o�.��p��;�Aڃ(�S����)Ŋ�W�*yL+�WVfzA��\+ش �C�=��A�M\=�SX�<%�t��e"
D��������׷'nc���%�A����(n�s�|uƺ;x����8�Y@@�w�a@gr76sG�e.���v�8�KD�'Qy0��{Q/�o����M�7Dz��p�J�_H��%��evD�?,v�]J����8V,����("l���g�n�NV;1Y�ea>y%ڍvT�a�F]�}���瞶����(�J��}�Lv�;Yyq+M>�s�l��l�n����ܢ��w\�Y7�|K��2Z]�9��}��;��?�20����@�/J́�����N�!���'� >��Q%^gzni.�zY_�"pyܲ�������k�p{�f����]nM�	��Y���=}��ƒ3�~K���1��f��❛�3�V��C��9��u-7Έgs�a�^#'=S㔯��~�}B�э�Th���ׁTdW�.̓Q�����1R����T���ƞ��� �[��iex��U`йUPp��:���v�煋�_�A��OPɅ�'�1��6�څ��q��h~����Ώ�|wu!�o��dr�zs它5F:��gڱ�s"�҉��D�*���sk�ǣp���W���T��>9�L�Ҧ̼'T���uLO��f�C=1yfbظr��)Fͱ�S����&^���\VUx�<�ㄨ��*�L�|�u�܋�4\��̠�ż�z��េ`��g�`a��Zڼ�}qR��]J��s�(�T�tJ�i�y���sqF�F�s�A��u��x}j�vy�z�{�gN�e��fP�JK�>R�Y�]]~)�;����r_������7^��)�\�T�:�PX�
�TZtha\�u���)>�[R[��rڸ>uq{�N�pk��Zx��\�)��>��2|�y�itooV�;��bҨP�MD9��[�{�6:8u�V�[G��w�58e�K5���F��hf���/�(t����d;�p��1.�J7gI;Pf4g�XƩ̉C��1����#�>���S��ybin�3��l�<������Ҳ�,%�$�����j7�Ļ�҆'�B>8�9"���
6�m�\D�o�#���s΀Zn1���~����|}J�/�O��ۢj��H�@N�7 �z�VV��[���{ǡ9:y��X(�z��;�E���0����Qy�I �%Z�)���W�˫�dJv��1�=ܯ���kͳ�����~���k���ۇwlиS%��!u��&O>��Y����N �>l�^�;�YL�q��a��Qe|\�%C��
T���eI�&B��Oa��F�PBjbgK����Q�?t�>^�q�\��9���|�2[������܃��^>Q���T�r|�����ʇ)���lG�p��w=�3��]^t��;`ix�����^bK5�`���S�n���ˀ|;9t�tΟ�����{a'�V�����Bv�n�Ig6}�[}�c�d�I�ٶ�;_*; ���?@ς�j�j.PG�ò����%�r��OQ�s���J,I�z�]j��D�"
tE��`bv�K��N�ޡXp�V����t���3�@�C�GY��pڗ�^(��xVv�U�V��b��㒤�S0 n�xop��'���Ug1+��Fׇ_���+)�_]-'Nn�f�;�y�i��L��P���t�{m�����w��._�����9����w�[�C����;�j�?[�K䂌E˺�h��2qƏL�_�}�[ucw5��U���"�ݳ!�?"�Ed֙V���P~�R��^�}���������E�u4��t��S�<w��\.=ީ�Yd�Y�X}
`�Ъo'^gC�#l�����MPag�-�R���<�d;�nDJ��k�R7g����
�-����O��p�+�xˠ�Q���:刖_:����8<�2���p�N;T���yY��Tߪ�{Ԋ��c8J�:	;Q3�H]P�*e)c/��*�ЯF�oNF��+�7!uj�?F�l嫖����5���F�7��'����-)��R��n�T��P)v����C�-�q�����o��\��n����0��rQ���d0
[$\ϧ6E�J�"��x��e_��׃=�Hhq)�C"Ͷ7Нn�q���n�m(��D�'I������
��(�_�PØo�f������R�8E�6��VV�;�(��$���5�Sb�UD/�Y�p�d}o��!��纏u��#��ฦk�Y����I�ٜL���jԥgX�{f����x�@�jr�æ�z��ݹKx��oWm�Y��]��դ����z��ɺNʏ����P������MZ��Zp"nu�-㸚S.g�7sMW9݋�h5^3�ǩH�.I�.�E2j3��$&3a.�F�7\�����i�;U�wm9���=%�..o�P�3;�q�^�
ڔϨ���Zn;��<]TͯJd�Q��=���=��U�=�s���bd[���Q����%�l?EJӱ{o�����W�Gd�U:.5V�cQW��8�qJ��9P��߬�q�L�?�FHj�ml;��;�n��͹�J(w�S��]Q^{�=u���ۿ2����C��F��v���,*��>fl�us�x�#�ݭF*���S��h��qS���=��ĩ�UN�s�})��\$~[*�SaO����ʌ������wC��+����g�=�4������7%�ǻe�j�v}�ǯ�UB��'^��6$ڽ���n��n�Ш�o��)�����X�d�9L���}]Pf�m�ݓ�{(�X{�.=�����9'F��'j&x*�3�I?)\����+]8*Eۖs1{��xMf;Ѵ�pn��&���uY��ޢ�:Xֱ�t���a���K��Ԓ�?K��٣���/6�a:^�9#�̺[,�)��r��E%�>���Э��R�ܵ�-�uw0�u� �pŅ�5�9Nh:�M�o�a3�����eż�[v�S7;y�p��;ò���Ug�{�Q�$��P���p�ۺt��G�>�w�e���]+���8�s�4j�(f9}˪���a���x���\D�H��C��qqJC��\n�C��d��u�(\���!�SG����_���n���%�D@��x�)I�U}����84�qw0���}q%��^S㾄�F�q����v��Bo�Cⷭ��&5z�ѽ���� ٨$�h7�+Ḱ�����G����D9��Nr�7�6��]6����}�O�?�����L��I?Α����R��{>)��&3R�r}1�sU�J2~����_�%�`1h߼5]қD���;7f9��*u��a�G����7�#Τ�H�ӫ���B��0�N�n\y�U���5Q;C$>��@K[{	W�����c���My/q����Ƥ��\/:�ۖ��B��H5�d���\C�>�U]��&��5eό'�*~7s�W{��ћYLlr�zr���:��g!���]�/+�3�s�ڿ~��deo�]�"lGy)V������N���ٷƦ��nֺ0*e���'׹|�\lĪ;�)n�1F',��R�N�2f�������n���x�����活�/������{��ek� �xh�\9܍��ڗ\Q�2�%���-���=-Z����7.� v���y�xkX�@K�B�l:p(�"�y�����M��Ɯ�xR%�z����R�Ґ�Q���
�H�MgXlV+�h�,Z�r١h�v�����vb���l�5,5����#�X�����8��w���s����ᭁR����sԪ��Z�y3X��t���j�Sz�zoV���v��e{��T���������s�x|Ob3jB-�ʬ���&���x��kr����`�Or8�Ӹd��Z�FN���h��@l�NSg(wNМ�)sz\�,�bx2�=حúQ|!X�]Ձ�5+���b�5-�% ����:E��_���M����Q�H�rҭ
�U��8���,Ι����]iq�n���51�k[���G�,a��ܫ�^�_}���Kf�Z��0��y����~���SMw�&S��U'/,�r�x�%�]���3��n������V�=ڭ"�cħBG�l׀v�ֹ)ۇT׮XFV�˻�!�����T�r]x� ��=�x�V�+61�4��+�����
��ͪ��W�(<��O:�'1�$�:$Ъ�4>��6K� �v��a�a���+K�G�WT��IV����S:�&���d�}�P]n��Մ���f>�jpM`S��B���fc=z��9#��>Hs�t,�z�'�lo�DSj2���X�o���J��I�"H�Om)�;��Yz�e�]3�� �b�1� +��ru���vx��M��T������ϴ���5b�AZ����>�;; ye#[�����3����<�W�C5m(��qv+u+�XC�Q��(���z��)���5P̫Z���кE���u���&n�����m��#�y�k�	ٳ8��qq~�u��z��4�<=	�\4\�㽖��Gd�R��L)5Y3����ř�xeǴ�	k�F��XO9�V�V�R��h]܃�iV:|�ͧ&s���qK�E��A�cڼ�=Α-�uť_�}��w`+Q���J�ٱ� ojc�a,�O�"ҭ�Jg��{U��'Yy����$V\�{X
h̫| [���s�+�)�����ai����������a�֙ZϏ({�50�h\�ni���k7k�dU2�:7�`v�"F���L���*�ܾ�JĥK�f��o4+���b��kS���Y{\8�Rf-1[6U�.�[gQ;��[�,��)cd0��j
+b��k&���;]�Iu�܊ج�&�z�`bv�d̕3x�v7}��!0S)*�`�%�!IB�u����j����7��tS�j����n@N߿_�~|���{�w�b�!�!�]�wF$�#�L`�* ��urd˻�#(b�c\�6J&�!'8�nh�F��cF�	�)�P�$�$2�0��e���J1L�B��Ɗd"F�IY@)wk�j$�@��Ц�JLj)$ �F �� i�&2$0�IE1��T�#&MM2b�")͌�B9�%��
�# ��&�K�1&��]���f`K3D�LP�2K9�$A�,@PFM("LE#!D,JDI�-%AF%I��H�i�(���F��u�bB]�ɣ	���4I��`�f0]�����v�X��k��F aΤ�Ղ������g����Elΰ,=]M��RN��m�d�L�]֫���.b]}�n�з�52o���þ�@;�:�)�u2��85K�߳��ю���y��T5u���pZ��ݿW�O�`򻷡�d�����v
�u�ZD�d���ʁ�����&���_���F{�2��Og�G���a%�j+M��Ņ��;ix[	h�M~g��1���^�^� �+z�����f�\��<D;����y:�1��>+�,��P�J2��3�8^,��������qgv��L��!�N�<�x?w�Vq��w�Q���'h�&G;S3��v��>���S-S:�����b��>���g�Kg��@-�N�zs�Y\@�(�����<ES�o�J��&~2,D��te|Vz��,ڵ�R��c���r<���QȞ�]z���̬���۵���6O" �$ !)���;k��|���\�}�>*q��J����%3�z�>�Y�XGw��������2
5iꉐ���3�8Ǣ<��ro��y55��yX�Fz��{�|�}�n!7pu�S4=�J5RB��m2y�кS���=��}�X�v�ܕk|�LCI�Э�ck��x�f�oޡS��2^\�֦t�	�D;k;I=b����*�XIL�7i>�oDb�l�w�=��A���z�u�x��K��wkkk;�Rg��F۸c�탵ǂ;���#�F�嬓YI23�=V����c����v�#��[g�[�,�s����d
�R�����;bf9�	�1��[��ɮ�1�;�g�vR�#;&���v�Y[}wB�橒���*������D�H{���)��TY̨��*��Q�}W�\-7�s�c!�WFם �Ӷ�����^N	�:��Y��u�[�p�r޹�UA��1��K��ޭ���w�K�~Ϳ\vrwzqk����W~��zn��L�@]��ByǷr��~���`��X��+�������t��n3o�=��K��)����F�f=�{�w�=wpv�&i���8�8�R_���X=>�����~'�W�u��zr�S�~�Ur���!uI��U{��%V7sU��\ϏNg��%�C�lD�ا�ֆ�J�fn�4^�����#Ƙʐ#~�i��N�<�xg�y:��:o���z���~�뽏j�Q4Y�P����r�j�>�nȿ)M��S��7%e���|��{��w��~��E.E���%�9�za�|onT	Ej���]?���G��}'º�U�:�D|N���ț���xe���7z<;��ŋ��+�5|��'N�E�Z�C��݊��}T`��S��;>i��F��� �A>'� e<���3X2���fM=��Ipz��Ik=W$��;ހ�ٙN�r�dX���'4�rn�r6�'�z�c�ܴ|��:	:J�>�RJS�'���
�i[�U*NV!��e�SK-�)��L3�1���Mc/�Q��2��<@-)᝗I�f���������7�;�Ԝ�b���`my���r<v��>��wh��%������-�*���5+Q���j�N?��	k�:%�h{L{���o�>7N���#%�8���V9��.�pn[΋ނ��sN����`ꄭoaɫCuĸf�'a�^�;�T@7�W[�³}�]�S4�����tn(�>����s7��*=p�[�i��^L�ÜuyO`�Q��ծ�L������s(5�> ���=8*Vׅ]Jg�n=Ҵ�?T>��wE߅a;�1��]�M�b�oI���#_�f�2�:~ٓAHeM|mxl��ѮÂUd����n�i
��X=�;v�=|Z�e+��p�{]ޘǮ)Ѹ�r����o�/�p�id��]��/�Ï����F�h�z��F]4M�ަ�f��1���FB�C���s@��1����^Tᱥ�&�>U���4~����s��h\��a�8�m�{��}�Q��~�����4cQX��b��N,�w�xW�e�j�=t]�f���B�Ser����N�R��ܾ�p�����{s\*wGbjup&�p*���&?jC����hD�e� �.�]^�,ل⺟�u�}�� �cV�}�w��s��W����O�eH�Ys���w]�&�VGl���*e�{#Ɛ9*#c��nO��j�MN���o'�{F��'���9���rJ\�<<K��gj:��U�t�ٗ\x�d�9L���9��{s����^��wN'O�m���O؅���t]�v�&x::�L�"�As~}5	H���������_^���-��"�s��ΕC�SzR=�(�E�v��$��*z�i������o���ћ/���U��s�4f�t���#�M\=ϔ�3 \�i$�A�JM������q٪��3D��s��>�����k4P):��5�h��5���s���n���rY�~�0����7qx�8�� pf2��&��{0uB�y>���_ �^�4�F�q���-t���UrW�,�;���	6�W�ܙ {�Z�
��>P���1��rv�ޖ��v��.���k��I�j��}x��^�߀=4��L��uI]6vH�N�T��{Კ����kAaW����ˢJ�����Kk�f~/��2�n�8�vo��{�i�c�pvk�+�n�\�r�p:99�����`�g�^��wy�.[�c$��0����a�ea�����V,R����|��%����y��������.��M��y,��mb�3;-#�`��<�g ��K�k �6��*vl��;�Հ����9��z2F)�S��s)�)�;/����D+���_4��l�p�.<]'G���[َ�lh���LU[���^.gg���i��W������Z��o��v��P�s 祓��ȟf���M�G���	�wN��q�/K�w[/�Ϳ[ʩ��Z�3W����oj�@l$D�a��}���Z���8���>�C��|n*ex�qL߫��������LsS���@����ɜ���8�=���Y9'/e����
�%ς����S̞9��9��μ#Ց+B���%�`���w�jO�]�����r|}q2�P����K��q*��.��)�U�z*�z�sP��V�u@p���l��cy�X�Z�������ˌ�3��Ez�I|��;���>�뺂+4��<]�E�ä=�'M��u��S|c~]�hi'{�>���\<��h�[��K���ϫ��L�7����,�>�-߆DyĶ}� /'\�����O��=e�5���V�zۤl�ץ���c�>��j>�R��uwyh�t�(bOE�n����d�שI��	P�R*n炭z4:�u�:�OyWdpV�h}6�חN&��1}�ɑ�6��i���v��}���P��`9�P���j�sU������*]6����g	;FCHyF[+=j���}b�%+~9�5;�t�r<�0�T4���{2�|ȿeW�?��]) oMI@HJ�@�;�h-*����[�㸜N����7��i��최y�x��'dz�Z2�Dt��d0���ȁҸ�.��B�={�sn�m���Fy����g�&�w]U3CЦJ5�$.��D���B�9��n�=������Ԭ�#�5�dz�u����9�s��b�z*���ʓ�&c��nN�`�th�0�o��.���*��)�j��L;�\����5L���� +�Q�wp�����A|GNaUޅ�[�2����AYQ_D�׼s�-U��M�s�c>mUѿ�� �:`x�����|"�\��>�~����̩�K'�H�N��q^���wg�*k��������S'�����ׯ
��ۤ'r9�X�/�9q���0���x��V��~㾀A ��yu����E��{'c��ٿN8�SO�1�̯}��k����|1\?�����;��Z)�� }���nPۚ�ٸ�<����{]@/����]C\{��8��%��9|�n���ݎ�J|�m���~��[��ܼ��N��WQ�^t�+ZX���.u��k��E'�9�ŽAN������l���<�n�WWB;�����;��N��c��u��&�F� +��C
�<��*�q܄���{��"���:mN�!��}���3r�����d�c�
���<g�Ժ�G� +9Z\u4��t��w\=�"�p��ީҮ\������|j�F��k��Fv��*�7Z��4��tGG���|�}���1���Xފ�[����Ǽ9Mm�>�z�;��N��)3�
���mʁ(�-Wp�9xq���Ø�`�g^T����x\O\���p��^_��.��z�ˈ�*Ǫe�]TQ�+Ub�`]��`�^� �(]�{��B+�ǜ�v��}p��2�����#�`���)��Fs���v�Q=�~>Qץ�n���Dr����x����\S�F@�(��� =��z�w�U��kP��˺RC��Ns#���]p��-�C>/6��Bu�M�w��۸�	E��r9�E�Ss\s3P�L@R�O����Tn(�+�:�+[�G�&� ��)�87���־�d�mn��އ54�\d�L�##�H�{N��QZ}V7�/���P��}Ex?���
SW�D��\P߇��lXmM.�y��j[|�'F�'�o�Sun�r�;�Fl�|�c���!ϴ�kL�:f��Y8�	n��&{r���:>yք�]śމV�~�D�i[�JV�aV��W�ex�m�6:�r~`�����f��|���Q;kk���� L���`:���y-���V��U5���Y��n#��ø�;��P�a�����{E�O2h��>�j�^��ɨ�zk㒆�8�Ox�_�m�S�5
m*�{�.�����{��߮;!�w�2��F�ʀv�����g�Ol�]W��N2�=[�U৙�Ӕh8���w7k��ͻ�c��\t-t9�y���~.#�*p�F�N��Gt%�'Mg�&��_\c�V|6�	�1�YOM��x{� 2�SS���s���!���v#�D�V#qi~�:iFۘVQ9�#�4Z�M����HY�Y.Sr]L{�[ҳ^s=[z����^o���y��T��Y}�4s�<<J��v��"�W�����.�L���]��������>�[�:G,�:{�n\r=���w!�b��}'E��'I���je���j�Tߧ�u(̐���ܫvm�����:�+�>n[=�;Wr
��p�x�7{$�(	�C�[����A�3�+$�m��9p}w]Nr;X��'lh�P��A���܅5���rQ�GI=gv�7��3��y�sjB��4�\f�	�:�2��U���u`�]�
�T����yR�YD���pX�����v���Ɠj������8���?�w
���w�*�֚�����j� �)�8$�y�.,I��e�ӵxOv���Sk����t�K����(�I�}}uZ��(\����4{�k����:�|m�w��7��Jf��fU�:]��Fc��I�����Ǔ�-����|w�'Z4�68G��t�f�W��z�suX'ĝ��鯉 �J��/�ٞ�A�o�P�	�m���2fc����fJ>H���yA�~�~����.i��%�WO���p��Z|=�e3�bS����bo�����3��RR+IE�s���#XB�D��;7f9���R�Y�/����I��&�I�kƽӾ/��D;�����;4o���א�`�t�fI�Y<0�۷�OW}��� ����2�9֯�"+e���Ԇ�u߂�N:����w�čw2c��(Ca��=��g<�hX��c�� O�ceO���z_{���q�~�9L�Z�3W��)ٹ�#�ET�*��WxK�h<����D{�b����W����Jf�m[��n�y�m����S9���]/��Q;p�٢�Y9'.6X:v�� �a�L�ڙ_��b4y]&�iw���i�Y�銆����u#��k�fނ&��wj�bY�[����°�u(h:	K��]BG��:ܡթ�3�=��ǉ�u�M���;��:��Cٵ�K�{K�YۣE�Qv�s<�+N��6�*�n�L3u�|n��T��w�2qƸښ�����<ڨ���{�a���M�ļ-��t��3���@G�)Ak
:��t_�����@w���T�pp
t��Ս�^�/V��?��C2}��#O3��L��O�)U��!Nt�qS<��s���d5�.�#����t��w\�U�b�z���=
��#;�\y�'��fU!qS/�����,�4�~���G� �:A���>�*�@qS��oi�۱�IF��K��L)�*�ʅkn(�O���H��(�QK+wW��8�ϭT�f�᫶@6J�R ޚ����U��;q��.9
�\Uh��5,�U�n��u�}�F��/㳌��5#�o�=t�ћ�2
5�F���%:@)�˳�c��c�G����z���>��r��c ��h�ϼM��ۻ�h"J>�X� �s�5�Vd�z��`<�L�R�+������#���C}e���*>�b4N�ב�C��t����3�}?�蛲*s�ѱE���j��.VaŷU1^橒�3.#T�������U�m��ժֶ��V���j����kU�m��Z�km�ֵZ���5�ֶ��V�Z��Z�km�:�k[o�֫Z�|�V���j����V����j����V�Z�ҵZ�����ֶ��Z�km�n�Z���Z�km���
�2��s�[B�������>�����f��;Ϫ�
�� eM i�5MM[UI!"��R��%(�I�RUs��W��c[f-h���D�hm�m�6ѶlŰ�����j���V���KdJ�[(�p�zI��),�[T��,�eM�ͪ$�1�mk6�Ԧm%[[H�PmJcVԲ����4i���2�{`��u����4itlvw[�V&��J4�;6��UkuM%J��w���,�[U+� �u�ֶ�5R��M�Z��v�� t�@ �   3��
 ���  ��Ӓ�닠/f�+��3sqI�Q��Q����gk����;�k�m�'�nn]v���N�̨���P���Gv:4����Ƕh۷qR�MSh��I]l뮨d*������L@���ܳA@A5C�Q[jS�]�Y�� �sX������t��*��VçC���@���δ���՝(]c�ܭڝ:�w:D���l�W7q��Q� =݃֨Wv��5lv�Ѧ��Y[u�Z;��FjƺU5��
(.���
������T�n���5$-f�wF�J��{@�{��������s�M78�@��tw3C�� �9��j�M[�e�5]]�s�صE�.���� r���ݺʫTv���j�.���E��A�]iF�-��ݩ�WM��.��+3�]�ۼ ���U�j�S��\�3v��;���6��tbv륭Fv̻��ۊ��v�T;9ږ��� 殪/u�uٷ7'l����ҝ���ɡ�Sk6cT�;j�Wct4�      ��JEP� �  S�R��FL �d0"��	T�	�� M4�h14� T�A��J�`   4"��<��M�h�� i�h R@��0�	�jz�G��M���f�א�S�(|D��2`�,
�l�+�Ĕˋ��AC���4�~@(����6PP_�PP�&���YUD7��s��?ſ����v��h=Rh$SuPABL ;� dM$������ ((q	�~�>��}��#����?_�v �(w����q���>f0l~�/0t��9�Λ�F~��}�Hk���=���������N�s}��~p�sw�+8��h�:8���1����N�fj��Tv��P�vx�ϋ�fVc�,������K��6J�ʸp�P��C��(�c�[�YjMtb
 \�n��V�5��'.�x2 �mʚJҙQa	+J�y�Rg�d5v�d5�,�:�sRǈ]�Yd��2���GF+I�U��Z5x""�a�l�n����m��S����mHJ�{G�5��jl�ZJz4e��J�[�h�O"�p�8�)yYW�j�אP�H�aג ���C{A�=���Zu`�5@ٓN�âq]��U\[[w�vH�ûT��Z��%�34-�,b��Z�����T�8��M�,I���P�:VV�3,ӖZC{��ԣGul��
18uPѺ��ukZ4.*�̛R(��ku5�1Ǫn�B�h�1E��r9��-f�[ȍ��l�q-+)J����;L<��B��:{O,��UѼ����kʙ�QZ5�3]F�d[�����C-٣�^�Rj���]ᗎ�y��4j�1ᆭ��ɰ+�"�Z�f�Bx��L�d7X^lJ^ɌL��-�V谰�T��24V ��ӕfM��É̸�&S¨Icp`���f��-��Τ��{�~�]0�k�"y��e��j+r_�w8��yd-8�J�`�5��թ��ӷ"��ؓi+z�	a��<�_�%JV�2�%;�Z�45��;l��$^�X�k��ن��2LY���scO0�cR�ف�&ʶ5�O��������ZCE�={�N�V��w��Y���9;�rYכ�k�� ���El;m�Y�c0ØNC�*�l0�{34��5�$suakV�/�>̗��M�?�ξKR+��*�mWXV�_ʆZ��%��� ��y�ݒ�ݽ���Y��t����<�eދ��8%ŕ7��L�v&��y��ט�ՍdqaHSٗ2V��n��t��hM�v��+)�RsM4lCM)�oȃz�%W+��9��F,m���^�����(P�b�7�i9�3v n�Ex
���������;�D�Z(Ս�D�c�66��4��J�1:j'�VʁeB��1�1:�?
8�l�B7H�K)s����Z���Ҧ�T��N��.]�4<�q�w0�B�G/i��E0�P��5�:��؝�]ޥk#Մ�(*JaA����-!���Hl����*�%|� ����X��2��u������[0!�j�=C>�����y��f���n�M �t���B�)"yX���͊�}g7HѲ�hE���m1�������˕b���<��Ab���ؓ�D9H� w��tL��K3f���Ƞ���U�� ˔����ncH�{K/�%5�sr1n	���� -xT��Į�4��g8�E�I���k�T���E�ܭH�31T�g~��bsn�YyRcJ��P��7:t͗�i�m�+J쌳R�E��ۗN���JK��ۛ�z�c�r[�D���-���P4�
-��~��ݖX��J�2a��6j�I9�:Ի�\��I+��Am:�nՍ����R��o2�%�T�3l�6�(�Q/JJ�[�i`i q��H��!�y%�:�L9��6�Q��A�b��K���cU!Ȏ�쥈���xp�j�[���7Ij�'���߬�2��Uqاy��E32�i��:j"f�ڋ2�z��"��e����˼�-������Z��7��a$�[y��G�V���ܦ[��"oP	�K&�m6��m�L)fe�	V�g]0t�)�z�F�N�U�mq�w���t:���M`�J)�m�֜ƺYD1���L�P����P�,`;���2�x�2%0 ٻwN���U��L����WG)��R[Z�&#�� �P�k!Û����i�+r���?]̫�����jld�Ȳ�ڬxY��	�(f���	�*S:p�V��ŗX�F�zL��{W6�{ZY�F*)�ӰßJI,b�R7�q-��+
Gaӳ����b��M��X��i��jEVf[�(姥�.LG,2)�>Q�Cj�]QV���v���oi#Y��R�X7S!�#H�"�{ WcR�2�S#��c�%�N�-c�jj�xXWI9g7	v��N���KQ�zS�V��e%h<���ۚ��e�+4�CVYaCy5�0�=*�)�$<3k.�Mf[���Fn�d�n�U�cS9���R� -�ÀR�ɲa��R��<^C��R��WLJ	2��hݔB����C5�#�t��E��e�]�$�)�2�j�Q�Rl˫H�13k̓&݃&�l�Q���쿋�,XiH�*��U�G*�9���s�|�o6��0���.�/�A�*��k/,��`�)����ymAMKJ�'I���XE�W�ak+&�����uѲr������6幙� SI6m����C�KwI��z[�;xh�փ��"G#7[H�yga���!ˌ��Z h�(�x��]�6rh�0��I���Y�#R���2
�K;�����Y�����Ic��іE(� r�(��Q�k���9����Ӊ%z�uhmd.�i��l��ʂ�U��ʲ��5D�Y%�5ao>�7�t�&[`e�ƕ�D�l�׎��)3Eԧ0B$�v4�K\���-QF
6�aô����՚�D�Cn���֌��i
8��B��C~˕�lS�3�{x�ۺsm��&�i��b��,$���S[1T�mn�a��xcrZWX-��ۋv�;����K%Y�:d�Pnf����-e3�	v�	�zE	�N�EL�nv�a,ݐ^�X$5a\h�w*]����=�����ʴ0���E�%Y�T�
[6�ń�V�v.�ѢY��üa�m�1)�O�Zڶ.�dC �4n���#'4�8˕�@�f�͜�dh�r���+����h��F��Z�@�yt�,�/�h�S�F�n�(bɸ��ejN����&`���1[�h6�օ���j2"�4&�F���V㧢�mǭ��
V����������a���ڴ �������T��s.cАq�9�S�U�/�3��q�i`±X���ܙ.B2�5oS:쪻W��	�;ٴ���8ɰ�Ɓ5�0�sH��$
���P[I����$��٥���lXT���> ��z���L�&��=�|�u<�����e@��&�z)XV��{l�Yt)�)<t�)P2Qμ���+�$j��[�7�7uUm4vU'`+�l㼒�ˣ�_e��{�k0$)L˂*�f����X�[9su#��Dc2�b]�X��c&�*��G	��TT`��Q�mAr�n��
�X,�)I�m�0k��؛MP��մj�=���Ē��3u
[��)j�H�Ҭ6�X¹��L/h�Ճ�Q�A��j�f��ŕ�i�� �(�~6��sUy
s�7Y�cj,,�E$�,�NT�Yqd��ެ�O*��:WB<�����������J!��p���.��l�7K&;�V%2��³LUX{�7m#N7u(��n�A�ӡ��٩7w/F��&��@�(��l۠��"��m���I�&��*عcLKg���I�̵��LѨ�y��=%\��,����a�c-X�v��0�&.�&�� �=J���%n�a���*�}��S�v�A�U���iV��Y)��	���V��i=9�����j�[#ieZ�����X��b�Z��j�˗i[����ԫ�L�I�w�WM��R�[in"��ѵ��L֭��A�a�ջWXz�#G-3R6�*(�ݲ[��f���X�Y�v��{��� &{blp^��F��W��ՍRv
H�-ӫ4]��JQ�����%�j�V�w��9��Y�M�?���a��%bf�ph�
yS��(rՠ�(`�#єq�j�>bf���f�p)��c^@�=E`:騡��T��+�-ݓG�b�r�Dī��5���h˄�s%ld3&���73o(�Udz��t�¦�� E=j��pZ�Z�٪- ����Iy��,'4ܐ��wQk�#�Wq���*��]i������M��݇����WYt����\P�����v��K/A�@����,hχ� �߈O�~�����? ���u�R����>������b}E���m��g�xtu������mk���        �w
7w3                                                                                                      ���讛�����d�ш���Bu��h� �s��(�H�к�b����V�q^�&nfnG��%u+����V�VZR�!^[y�8+0���ɫ�G��O�e�bh:�w�	}7�K�_[�N��{���Vu(s�JN���^������{/��cM4����O:#l�S�quvZU��a���F��ֲ&�%�=!�]�D�jI�^����r��ԁ�:vk�v�ud`�.���f���;cWe�f���TZ7���9zaVz�7�jAWZk&θl���Fػ�6[�r�a��:,S�%��s��5+R�c��o��w�F�TP�%"�I>;S$C2�9�"+��w+(��]�^v�ܐ]Y�mP�uo�����٩�k�g,�������7F�����m�d#����f�E;��l4��������(:�V�*�)�ʆQ?;�0 M#O
�M�׮S��H��z,�r�]�ݓ��"�&K��h��0*���
VC��]��W��-:y��E5�,O��{-�W:h$�n�bZ�l=�	���F�l*[�k�2�QjLDgX�-�^DQVj��.��
J}�3"n�7�N�ML�B-U}�U�&C��P9����y%>��+�d�[G�wk`"�DV^��Лc�H����zL�w�5e�����FV�R��j�gv��:��vt�&l���KH#ς�����!&�b�����w�:�>�K���
��Ҍ��+�����=�BW6�Kj*8�'2��OaS2	*�E��&�BԭMEًbZhKŖ�Eţ6QjbR�ݝ�NƲ7>��	��v�G��z
)��qޞ��k��>sari���ei1���b3mR=[��Ml��)ԷݖZ�Uz6h��+���詌Z��@��Y����F��<
����}h�;+SR
B�j�Bֱ��Syp96(M�RȽ���]���h���>X���6�p�1�̜FÁ�
��	3�Q�5},i,�#��E���}�{�TwX����]�o'02�L��]G�(�t�S/h�O
��Yҭ���K��zE��L�%Tz�j=��I�>������Vk��n���z�C�r�z�ϣ2d����%]ą���̫ѻ��,k��<�ud�Vr�4��m&�rɝ�Cl�3��.ť�RU29�a��>sL��2H��νԪ��ג�>�&���&�du��j�SK,Q߲�HƷI�lLf��b�T�����'n���V�8eQm	A�u�\Y���c��6��CQ��'l_#C�F�������t�h�X�r�]�%�Δ.*p�>��B-u.�흷�4��<tTG2%6�zs~����:iʎӅ`��e�;;�� ��+En���xN�/Ɖ.�sk
yl� P�h��ڂ����
ЏǓ�5�X"+HAiW����]���i��)�I�)YS����v��v�HSq�2!��5i��[H0t���UY,��.i��勴�hC�r�i�ە�o�J�����ꤲ`"c��/(HKcӍ�ԋZU�􅢶S�YqV�3c�eG�����\����鉚V����;��P��{P�a�s�ѳ�:�&�V��֙��>�M#1�x_}uq�����$��«�o��8prE�:�3;f�Wҭ����<������&����@�c���Ď;�1��DS�PN=\�*��6"���T�;��U���H�֝<Y�)�+j�ۥ�K�]�٪��Ͱ�x���<�{#���'%���\�SwX�K�㕮el�v�6k�W�)��q���-X�:�'Wh�i�\t�;���E+��w��EH���p�7����sP�p�u���i෼��W�a]'ܬ��n��B�`�Y��~�`_b;DjvZ/�]ܒr낏�����3�ճ��ao�٤��VL�蜂[,OP�VYs4oV>'(A�J���)\f��&�����9�G�h&^��j�<��y\�����X�MI�����{v}�n,�t)c�jJZ�Y��Q]���z�Ty�EsgE샹o,��E���:�M��{y|���l�S�u���X�;S�÷;r�hX1S�Hq�]�F"&8�><�����%��}�FZ���:�AMs89a�O^駶�a�Eu,+v��p*씐Ö��j@��Y��5�LAjȪ��m�g(xIu��S%�Jɂ�䘬��K�s�N���1mrZo��k��qw�������*aSl����ZLÙ��� �:yX[�Ֆ֑c���U�8��-�j��3Y'�<�R��=��Lh��.���ln��<��u�q]�m�+����w9$�s\
��%dմ!��\�.:�f�a�#�v_��x�v,�6]
V��\&�}�/+l���Rh�6�4�ozþ�ή�I�f+�pS�ϻN��5c��}��f�iwB�@��)�r��Q]Q&�F���1�g��ǯ]�˘���a.�z�4�.�]wqλ�%�O� �=)aZ�HMv�)ukȆܲ�Z�iN��T�&�֫8.���I�(7�!|Aw�"gwu��m��v�*vA�w���S�i O]��E:�	oN�]'����m+�K�+et�/ha�a�n���w(ڗ�,�0�EQp�/M�ъn�^1n��ցz���ˁޮ�z�5YMa�w���+.��mB���-_K� ���b0k��; ��>��%�]�S��/����,�M��f����!K�"\呂��~�fǚNӶ�b���	ym
8*Az�Zd낪���m�ȕ��=˥H^���mT=G��.U��{����B� ���oN�r�~x�N�{w��8�9�G~��X�W?Ux���r�m3�ff=,�v�!�rRۦ3��jV!o�Nu:@��^w�`�u�-־^�{��@�����n�����%A
����f�m(�ogE%��CF7l�#v=�
���{��l�w(�o�
3�Uec,5��}��t}�xm+:�i��A[y@�+v���5���5;�QGYp�&;�Q�����&���kv��q6��x2��rCo�O�K6|R3�-�ͭKiĀ���е��\��㭹|���u��]z�&��%��;�Q7:���3e���Q�q�uwv3]��O8�%zq�2�����H�.�A{d��U��VG&���M��%�e2-��jp9��F��v�N���hu�߭!N<W���uX�Z�8mC^���W
)��wc��%�Σ`�W�e�&C;3o�Ĝ]�(���2�Zn���Iy�Ӥ�&Ҡ���L�+>ɜ�ux��Č����::��6!N�q<�D��� 9���v��T띅J����^�<�X�C˫q#è{�
���,j�P3�J]�d�����ʶ�K�V�*W0p�9�D6��sݥ���X��/��l{�B��&�Ktm�'.I��t.��Ant�lD�緲��M��dI�Ǻ�__S�H�	̶���a'�]\=Xx��@�כ�z;8b�rZ��F�9z��`�y�5a&p�H��]�vb�%�5X�}�}e��Π�$�4�m���m��f��;P��(٤��:�":���_*Tf�#U�����N���%�]=�t���cs��	����j΂έ}��N�o��󱛹:�$Z��\ajWgJ(eM��#d�k5�R�z�%��Ҏj��b�v��JCne���q���������&�HEm|&������b�;���r�v�:�%�J��c��K%�g��֠�G�h�kv`=��2�6+%�"�P4�����0�8�ɭCv�+^�n�0x�x-}�l���k|��j�\R[\��SOwKv�������>X�\�i���r��3R�&�(7��	�9�|`z�سiɧ+zM̕z��%���U���ENR�B�tL��.s+{F&��;3@                    �c4�ot0b��4��f�sd��o������f��                                             ;@z.���Λ��J�.���}!Uy��:U��^������}�����g��7~�~Y�~���o���@Qz����tQC��z�O;��&Ȉ���?2{;�/�����wַ���ۯ�<�)�y�ϩ�9i`V�<��ͫCpsk/�Q�(=`��Qa�^���[t����.�b�.
�m@Q��OK��0,�2�bh��U�Vzݬ�Q��ʏ�MX0���v������˧f�[@Xq0�iQ
���%;�՝Pb��u
�R�@^��ǹC��\�R��͗Rc��xn�"��#9\�����j�9e�%Z՜G�kJ3�d]s	�g�W&X�����j<�{ZrZj2�f�K��&%��ji]O2�iEv���Q�O�Ս�1"SǛ\ec��N
��?,�!YJ���v�e˥m9�>1wV�ϭ#�w6	a����L��b�;���'��ٓH�|�T�8Z��I��<�'9�{�ߕ�U��B���ղ�:3c�];���E|ѷ����"d�B���ڶ咘Ӝ�m�R�+}�/i��6��W�K��n���r�)�ʬ�+Wc�r�e�J^���5ԡe�J�8_8c�b�K�R���]8Ø7E�<m-0�l#��U����Z�H�A�;�׏�m�β�Y
�Q�/)C�Vှሊt HWl��w��I�ut��hAհ�"ׂ�N*�-ټ�	@p/�k�i��>�"e��/t�6��W�Zg�"U��H��͝-`!9jO>6-<�A�U-�p�y���'U�f��.�}$�(�\f�%^���+����X#-ݰ�=o�ᮬV4��`�i6�N�^��N2��qCH=�L�ҧ]q5he+<� �}�U'���]����)����c�of�n��n��nn������nq֞T')����b��RP�u|T�[���-7�� j^m�eX�
�]U]��N�2m��Ge�� m�ueoE,����ϩ]�[� ��Q�sz��%/�����<�0]�E��V�b<V��ST\,��g2� j��
A��I�t��gˑt!������nژ$�2��sq��Vd̓�#�s8�V��Jk��J���"�ǫI:�BxU
�0����3*���n�fP��X��U�WM�H6���n�n޷��G���L��B��6����ul�����٫����	���JǓm��{o%�.�<�04��/m/��_-�W��+Ɖ�X�at45oz�phwg.=��v՚�;}�"��	S@���E�C�Cgv�Qvf�L����1*.-ATL��{F�#����(F��M������
�,��/YӃf�	y��yg�c��-�e�ٷWA/��@:uD�vȮo����\�.�h�v���c���L�	�����"������q�Յ-˼�K3r�N�}��w.��ڴ��S�ҩE�cGr=��Pu\)�Ḧ�3&��H��In�%]��H�e�N.%�Sڵ��rˠ ����Uz&�#�bru3�����	��L��xu��x\��hc�usW	��I���aS�)M0N��V���gEs��e�k���P:��*�Tz��+�!Y�oi��D�/8��w�T��m0���U�}�R�E[I����c���k	l>T"��!�6�{��݃s����oYP^��ZA���u��kV��r�@��U�F�u���[W�b�=�ku���TYW��C��m�t2�����v5��0.�8ç�	閚��00(f�ڟ_ݬ����-Q�	s����뉠�l�zM�Q,�e��q�&m��n>����շ�Gp�k��mܓr�wt�D�N��VY}��M&�北��2��ُeX��k�JYٖi��g+bt�M��ÂCKor7��N�m �[T��M��j�� 2�p7���w��`��Z���������J��6�b#Q�a�h�-�}�݌��A����+��[�Q�V�b`����05��Hy�*<p�z�p�\cF�����+�����Œ��.��G����̬X�е���T���[Q2m�s�;㪖�@���Gh��YL�SD�/I�q��w��ؗ3�����o��h=8^L��.�Z~(�G�4ܰӣ�c��#�g�kR�&Gu���+X���جa8�9fF�w�t#U�o>S�P�и��:T�0����m]v���Wxe�,ɦ���R5Z�8���Y4���ag<��]�QP뢞�hU�O����ۣ�e�r���t/�iO�G���2vUѼ&;9���!
���e���[�g�ڮ��nE���!=�vt��J�W�)Z���x��x�ueV����b��fw��&IV9�۬��W�����#`�G-�S1WS�WuGSb��ޜg��~�*�N��[2�
X�<�� 4�>�$��N�J&����ŝ���D:�Ɵkhp��61Sk�;W��/�l�(t��^�	u�*|�9Vv��l��GY�J�D]7��
��U�S�V`����g�^^��7�q2B�P�W	�艾�
��Tr�8��9�cG��;P%��Xh���
Q��vXp��D�j�6��6�B�ۛ6��I�3�#˝a)�x�Ve���n��۴Z�]��ئiZ��{Y[|���'3vAWt��[��\}���H;��h֎�y�ˢ��eCV+t�O�1-�f�\Fb�9�N#�h��2��*�h#Z�1Ib��K�qi�:��
�g���gYT;�}1i�A,(`�b�����)\]-i�	�Ԋ	"���*iL��!9���$��H���(�3/]5�J���Ic���O�!�Xh_��h"��{Ǯ�{�$=/��U;Yjc;lٖ�񵒯:\�e��y�IKg+wk�
����QG*!��-um�#��䘮-�ʛ�f�+������F�#۳c������g���/�ǥ�eL�8��,�5��$���� ���c;��ںoD�֛��>�i>�DMM展��w�ͣ���Ol:�i���dE��J�6ȧہy����^%;���g�t��spD�9f�JK۶9*t[̎�Ff� � o/E���Y�hϝ�u�ɏl˴���٠���@[�aQ�ݔo�L�K��}v��6�� �3�T�Nw% +b�viܔn�*��A��q��$�Z��I	��*��t���.�K��[�0�9m����C٭	�(N�MA�]NJ�8�& =��L��iF0�3��Sw�_WSgL��9Ve� ����h�/2��_K�[X%Q&���s��1GF����Wb�Uӗ�]�eu͜#I�E�����o�]�������E'����y�R��5ݎ�N����팎i]|X���k�ksW#N���K�e�ݖ`��ճR�%r{j�]hAށ��a�7���a�Wrɗ�\KODċsa:udB�A-ݩ0��,R���{s�\��b�$�k����v���'�M�׌ZUջQ��FH����zz�N�Υ��Qlԓ�{)4^�X��¸���Z"\�#�]]�rmL�[-�θY�������Q����G(Uc{Y��,��2�q6M�`��xM
��9Z�W%osXe�{�n��ys3%�5\-ַ�d�bt�r-�۬-�]�MJՍ�@ar�쉘���
'U�H�LX��k9��޳Άf*7�{r�;�c8Àp=�C��WY�Ѵz0���h衲;{	����k,�4c�k��4E�X5�R�9շ�cޗ�����W����wX%��{7t&I76�wI���.�s]��o3A��瘾���`��mf'k@�b�O��53�2F���ls�Vh�^І��+��t`�̚�Q��HOu���r��6gy��3C�g�:����#���՗�~��l��ac8���.����iR�BQ3�����L��Kmܾ9��O��F�T��w`�[Y0��2��fs.ykʃsS#>E�=��EѮG�j��WV:�3���*tgn��W�u�ʃ��̀�[y>d��Z��L�����UN��,���~�,ӮF��i�i��v��av*�B'�D�̦��&��{��7�CV�)v� ����iL��g>[����g^@-훫����y�*��B�+��IbUl�ϒ��sml[����m
Me���* qSG<�+.����vi�N�`���t��-�HS|�gFz�B���hI�\6�pΡF��p����A"���jhB$�����=�	�m���w��^w�}��       t�u�T���<цQ�����k��Ak81��F.ҡQk4rr��p.��|r�=�%YIa1��ǲ��+���X:s~<f6H�8��\�f�o`sZ)m�kÿ��Kϟ1dj���R�3R��.���$�-PE<�Mofw��d#�����ʚ�U�,i�����N+��Y�iӋ*����4�`R*�c��iΙ*�������%pl�ǹE)�u躗�w^�\C�V�ޠ��&�v�ޒ���J�(Pb�q>���|�oV��.! %�C�is=n�{�d��=��8z��w{S�M&�5��>ر�|m_5vm�c���rSeX��!L�ù��	��SN+�-��V�2�ke+��(���xS���V�꧉g5"Oiq�S�NMa�&��!�k3�⟷t7x��8��  ��;�r��"RER��k�:�2�C&��2B����)
i�0��))u$:�����p��h�2��ԇ��T�K�#� ��HSM.�&@R��E
dKWCEm�����7�$��N ɪ�����5 d ���������M�W�f�3>׈Ű��q�k�c��8��U��h=+���x%��㌼�6ˆ��]��)+_����}�]�CX�V;�F�s?��[����f=C�A<vYV�>.�5�{��u{+EJ$2|�'x�����||Fv.F��6��K�b���O��*���C�hó�C�����(!��{���S�y4�#����pB�X����*����<쏅�P�m$����cY�S�Kr����a�W�-��{}rf{�g7W��M6�����{�~#Sy�v���ŏ�%��vK-�6j��;�/S�� t���u�:=��΢�7k���	���w�0�?��x�z�7�a�c�ƕv�X��=<�O�)jP�� �m�#˞6e��:�oe_f��Ϙ��0��r}dۆ�Q��������w>�[<��̵O��1u2������Q,{Ր}h�^�i=�1P�E���Zq%��ޥ=M��³Kbn|�6���p�c���C}�������?����m�|�߉ÎN�~�y�Tf��rx�Ij��c�#j�A�n;+�u5�"�r��lϚ8bf���<���`+t��v��_��<�N�^�q��s�V��X^�/g��+4�1�NE^�+�*0�"̕;k\�uQ��{��4�mnz�M�l���>������S}��ǌ���Ȧzs��o;~�WWGA�ZT�܁ws�P��L'Ig<�x�1��K��3C�ĳFR\љk�i<bu9:� �L�o����*t@���M.�G'{��w2�����A�u��Me����O��M�h�\�JƧ�,�vg޺*�,kW<��G׳����x�JK{'6^YQ���e-f�2�b(�<���M^�y���V|c�7ί�Soj՜$S>f_V`"K�m�ML���a�'`���j�R+���i3ֲ�V��8 ��kޞ���Y��x�'�]A��K;˺z� ��L@��S[�H���z�ڗuAX�U:p��S�*�^B��V׶����9�<�~�+U¯��>��v�u��^�4;�A�T�m�:���4��л-,�Oi%$�r:$[(����W�=��8f��{�e���������U����3���'4��٭G+s����6��Os���-��>�I����׎ꋡEZ�}X��� F?z�A�y�Z����ح�[�s59�H��x�)��rڎ�/[��=)i��7����є�u�[���p�o���G`x�[�݋�OR���P�ku�g��M�s�$��5�F�&�k�ΚeY�S,�ب���ت��0��I<��.��L��)cy;�k���5�q���(T��c�	����{)�ɾ�C��k��}����ݯ�0�8)�׋��(��]o��ڤӿ(W*���^����DFl;79e��9��Iǝ�U��ʀ�XC.N;6�̭��H#�U�T�y�2Ԝ�rH��[�Q��C�J������T�]�/7y�bgǽ�~O�p��]r1^(v���o�\��5�[oc���b�U{{�WIk&���E��X.�/�߼���p�������!���?1=���lO��p�z��]���H:[�jX}�E�~#�'��VM����Vvw yu�-&M�SN�F3��;6����㹛�7�R�_��/O�=:ݬ׋k7u�Yǝ0����7K�>kL���u�A��g8��������R����6qT�
�+��{�),��~�	�%\��;r�]�.���'���{��Ѿ2��_�Z���֑��e3�Q���}μ/o�>O��`��N��ޣ�V2ӆL�7�$-�(��M��A�ƳY�S�Kr�op�������%�D��ٓJ�M�\���l��\E��!ی�0J�-{]���gh�)ޞ�'��k�BX�=�:�8��
�ԌI�mOx�s�}>:$�J�B���m)���^&eWgd4�����*�{Xq}s`�ѻ���%7�㔡\N��Ů���!�ڹ|[KދnO/9�X��јy�@�����K��=$���F7�{�&��xz\�ǥ�%᫭9�!���7�VT������9�Ao�C����	g�Xp�x�D���{Ȧ:���F�v�^m5飞[�>&D-a����)V����KMKITWn�vsW'��j�J�''!㈐��0E�[{�ĵ){�"�������e��KWZ���(���F�#�%��g*ә�F�ͯ�fA\%x�����z��LYU�A�hjmO�������������Ev�;���6�O[X����o�p���AI��	�j�������Mz6�ݛ�8�zz=��Ӗ_�lf�d�*�ƨ��8�)��|}�W��z�9��.��xlP�{wv����\-Qk��xM�����C�rdy̥y��	
��D�5��52�d$����~���z��.����9M��ְ��4�*��PQz��g/}���Y���K�ݯC����ԡnB��G�q����xvvW�0�@��9u�;E?Ne4�Xαr�A��w4a�0�x�z�`��wg	�PĤ�������e�Cŭ���kٰ�^z�;�n�bΛ'e�wʅ�ªk�D���臆���]��6j|d׸ݲ����;�ҔqY�~oޫ�g1g��VU�]5��/9��݅TpmOfri�A:F���9����;{ڏ����xuOz������}nQ�u�\�ef��:Z��[+D�6c�&��C�m,�v�pz]�
'i������#[�Z3��kk,Z�"<����*������lON��y�{�)��˃�eω�NB��O���g�.��7���IK�`\94@�0��`֘�Qd��{�U�<���߰dr1ks���N<��(V�9�zj�ԩ�0fl�e	����VSl%���+��n��u{���Ӻ�"��Yf)=P�"�}�Z�L��ݹ�����p�9�W�����i\�*k�Ϊ\��9�W�T�c��Ug{Ȫкdl�N�s�x���� �S$�[��Es�8nYJ���d�D��Zdb.�U�ɫ~�F#y����]�5��E�V�_�9��
��ӮR�\6��,�7C\��;����\�X.�!WEϰou<к��r"V�t��de�ñ�g>{<󕬩5k5ܨ���jΟb���������C��/0h��D���j�)�����wQ
�
��u^�=e�u�$)���)��)�JXb苖ga�i�n�*��qꚴ���rt;{F��8W��a(�얲Z�tFc�Hg�+�-���wܛ��m�@���!�/�!=��R�@�	�w*r9Z�Sl�>����?Iy�4�R�����&�Em���]�m.��{�u���d��޹������~�͜kb~����}���ٻ2h*�|�bfY��T˰��a���O�e�����j앤���S;XtyI�iL���>�A��:?:5����-��r��ftFzL��H�6���Tfeڤ��:��'�}��W/j�<�ۘ&Q�� wb�X�O�x�~�?���ï3}F���b[jS5�����:Ά몴=�I�[�*��EL$�w-7�%�9Q�k�WU���5W/�m��^}������_t�j��owW�N䠰L����*B��B�o�)JM՞[P��
��0�ٲt�}BUc�H.gp`���mU>,1��-��6�U�4�]������S	�>*�nNEh���9�ͱY\����Q���,��pr��8xr�+��=��zm�g�uj��nb�������g,�Y1v2�.(�R�7��G�a|沼�(�2Ƈ�D��Bl�@��Z*�ۿ��l�����M�u�G�`>@��d���(�i���ǆD:�^͂�vظ�X�l��Vgr�D3���ʄ�=�[պ)�a�J#��a�:��"mS��x��ݕ�2���ʔ������!����,H�]�E.���OT�٣�obz�*U�JB[H�;���WcS��Y�.�7�|�T�N���M��v�o�z�A����        �{�j��nKa�y���ɕq�y�����%ؓ�ۓI����x�Qɀ�ivf��w!�@�:O�:�{&_iJlӊ<�{{�9Mi��k�#���S!�ƪh�`0�j�m�q�eXR靲xA�E$�>�
��!b�8h[8�=���]�fjtZF��7iC&ۓ��j�;W�0�/E�+�c=v����5NeK��dh�Z��5��%5��)>�B�J͔��R����>7��+r�T���un#	��vlvv`�s��=�0��6�^p���?JK�AL�.ÅC��Eδ�{��]�k"ZU)�{j[���D�C
a�8J�*�u�]��K����]#���x��
ѓL]5�,�-b�V4^Qi��ڃS�K��Nq)w���y�#��SY��ck��]���ٚ�w�p��  ���tu!TS��HSEq�BP�����I�5@дR�F�9 RġJP�@�!I�5�d��,E"�F�M�u*P\b�SA��4�F@P�H�j2���� �*"fB�59�dy(d�H���)�(uI3N��j�0(j�#3)JZ��W���2h���~�k�Q�Vq���mDc%�	l�;V�%:��?8�Ɗ�΁�#>la 3��ו�]��d��KV���v�;X��u���>^~��<�Oo1ɮ����C9�c9���߸���Fs���!��:}h���.����O�6B/,BI~Dr��|��?[z֏6R�Y�_�g����t��aLW�UoUÂ��G<���Ag�*CEЮVr��ռ���/{�f{˒��j�MqL�w��5ᭉ��C嶮�#��H�ꤲ]�ȗ���'�GoR_�S�k:Op^*1��G�u�o��y����t�DvA[�����=OU�8*e_�o��hB��?L��Y�B�A�^� �8;Novp�Z�i�&�hۻ)!���́��3��]��Y+��<�p�dK���� �l�P]m$UJ���	�	��_������{���K]?l�{Y��
����VRRKC��2o�,���w�v���8&���-�pؚ˜��kyw���f���eє�r�"��b�ƫ�o�~K>*w�%�V�-�%���ryb4�S]��5��[{������]�@�#��m�N���Yy�[鏌$)~+���Y�Ss,��o_��ߪ��VK伬f ��N��n�����o��d9^k" =��~���B�뫡r�~_4di}�14�fi�����1Y��ir_7��K�_Z�Qp����uL�,���Y�x������h�S���yh�W޴o��fnd���)^������'���4 �� ���M��{�t���vqB���b��v�aR%��{�N�f�����!#."��k� .^!���La#����җ�ߝv�~��x��w{뭍����>�Y~g�^�"Ϻ��ݤ�8=�(�[����I5�V�҃�x�y�k���[�P��8��\H��*\{V��ҫ]�������w�
��:� �M}�M|��_B辞*�ņ�oy�\���V!�{����sNC�����C6��]kM����F����⏥���+�>�:8bޞ�NH�v�~���_z�Y��y�8�F�=��"o҉���a{�۰I۟<��*j�-��J��躐R����V	�`�_�^�g���|�S�%���T��b�������[�6��Y��ovlW ��os�36��M�W纮V���=hh��a�R���n�pS�z.7������zG!�jϙ-OJ��O{5��Ms=:���w��ݡ�l�4z{-��:�Z�KaYP���VO穦���u��W���5�km��=�9�=|�J�:���z��$|��Wb=�sq�존%o)��W�9=�<����5y�^�k�ά��ͻ���Ng�0`�]�@�L�!B����fR�/���ة�����M�1Oe7�(�M��uq׻���Ͻ����FJo!ԔB�u�HR�ɷir �Z_v�8�#̼F��z�Ѷװ�k�8����s���|=C��S�xB���w��N�6��B��J�߮�)�v�崯[��i}��bw���3�:�\q��o|�|��N$�h}8�7��v7�w��6:��@�8y"k�v��
��%ӿz�������;�]��k\��~�ߨ�jB��^�׬�a��m�)ܧV��.�y��&�:��z��^��Ciz��Ҩ-��+"���Oe��]6��sJ�[ja�p#0����fՊ�}�S���o��Z|���w`JP�d�o��,�덼��z�I S�
ʪ���E<�z�<�=��,��>=�|����ߌ���N����<���q5+����.�:���ѽ��;ۮ����]���e�����x<Y+���=B{*u�4Jw/�=�Q��'��u��}���������|7��y��}��}��]�\iS�h����6���@��c��]����}g=��{�g��=HQ��q&�p���7:Ǹ}��WW�/�x������3����>�n{��ö�	�g�.���Sk�<��=9�y��7��^���=��6���G~��w�7�^{�=BRҜI�g[�vs�m�u�}��o!H�ǽb�W�m`u/0;y�ܾ�����m�0�˱���p�ǒ��'p�^k�~7��8�λ��=��|�%:�l�}��^!�7=��Ѷ��o)AܽK�By#�Y�̉�� {��u�:�x�N���^�`� |��3��z���߼O,��w��}��@����u#u����^﷼�ߧ��{�����G e��{���Ss�:�$)t���/Q�=��m'�H���<�o<���������|����:�7���G���5)��)�B��ސ�u�u&K̆�b�/r��퀜���'��{k��Z�%��fa.Lˣ�5�<����fq�b�toZ��-��{C�W�����%��y_��e��!�td����38�k�fU��4޿� �oy�����~�����=�B��qJ�SN�GR{/r�N@�IAܧs�� w��^a�\�7���h7�}��ͽ��v߾���^��]� w��������6����7�+7ǸN�<���J���@��|������5�^��}q��/w�x�=HP&[G�>�pm��R{!��ShC�89��W#\a�	���
N��~�ߞ�ۏ|���}��+�m��һ��;�Hm����b��x�G�y��N��B��m�*qϜy�f{�;y�]s�g��pjN��^�7��}��v�l\��8���Cl�#���I���������;u�~��|��ꇐ{�&�v�g�=����<��x{��^������dö�=J�ʞ랼��ν�y������N�O u��>A�8��5�K����P�����Z���0�=N�6�Hs��y޺םuǞ��~�j}z�;����B;��'r�y�ԯ2u�K�ď��\�ܼ�x���۾7����z��<���2G���R�:��'P����B��d�^��S�|�����:��]��v��6�o�6ֻ�y�����tr�f-+�`�������/6α<��M�qO%��%;��6�a|�^��\��q��;�k/6�m����ؗ�Bd×x�,^�-��"�<���*�J�6�ƅ��<'�H�{�������gq�sפK"�+!jR�gkb�c�nK����46
�?{�ff�3[�7���� mm��.�q+�|��J��`�Na�{��x����]@�%������Mvrg|�םw����<��<��ꧻ��þ؇2=�w��;K��
s�)�;s�pd���:�����N�{��n���\m������j^�a=�����s�0��^c��M�R���A�u�:����� �O%�-�|��ݼ;���߾:���%�8���v��^%6�ew��}b������5#���;�0��6��g7�~>K�2g������;{%�C��G�z�m��/1ĝB�;�����C�5��XjD�J�;�:����kk��;�}��8�ӯt�#��Z^��6�����k5[B��b���w��n{���Jw	�^yts�y�[m�>��}%H�)I�FH��%}��KKݼ@����:�Ԟ�>bG�;o�H�{��m���{<^�r=��Mw�{!I�%'r�� w/;b����/�J��<�8�G�=C��u�|���q�����~��Ԧ�i7����B���v��{��_%�8�\J�/{��/��x������dO,����?�D4�#�s��yoy'~b�Ӯ1�B��8���y��w=��M��d}����_u�ғ_��h;�,�W;�꣭�в�)�7ZyD�`���:�$λw��5����{�i���p~�#®�R�,���6��S	��}�<;�35��]�Ϝ��*�Ј-"�]oם���#�B�9J�-`s)��q����'RuB�cܽH���Ծ\C�)���ߞ��79�7ۏ{����d=}ŠJm�o�� Q䇐���C���B�m��'rl{�PRuK����q���u�;���_�j^%�]�v�5օ5�'1�>��X.�(�<��q!u�'r����%��0C�:��{�Z�}��=�y�>�zqq+Ԟ��̾H�w�̾J�ך�M���G'Py!�gr������N�)��|̻�/}�}{�]�)Խ�ϯx��A��H�@oq#�Yԯr�q��/3�[iS�iN$�0N��B��N���3�Ow�}�;�z�=3�}�ۜe�_. ��Xoq#Ժ����#�v<��@�Zҙ�p��.��.<�<�~���z�ԄJ�'3�X@���w/�b��R�''�r:9Ë�mb�@��`��P�}������k�<�{��2�?|I����\��Y��VR��?cA�aTV��FZbv��=�֣��:Z3m0�n.g��~s���Ӡh�Ff�^����^~����}v�\^����EBio;5�.W��譬��/��"tsy�$x�ZiPJ��g��On�LC�b̊��I4�L�6�4�VPKzDC�G��C$
@�~;����>^,�W�߬�V��ܠ{�=�B�ě���R׮��u��J�|,�I}+��qȂ��	ʙj�X����O=>k�YַR�u�����ֳjKU�6U�c3�`������gu�:�r�����91��Ԥ!��\�=F�[��meqg.j�ɕ�7�w&��㽰�G�p4���q�Cmx	��JƽZ�{��~���i�m�o_���q$��/}Y1V�,Գ�㔸�{��8�7k�V���������n{y���tf�<���v�����+�/N2���b�����~���s�UiwW���"�L�Q��	煮[ԗgeF"��qAZ�#mL���$F7�&��}�}���
 ZTAPJ
T(P�B�i��iJ��J�����y�:��-����{�Ь�ݶ�a\w2�f<�����qN\��כ>v��'��bȺ���Tb��_����?
lUע��_%Sm�m�(���ݾ</���Ng���f�� (VjiG��W{�&�M����y2n�3J���^�iW �x;��k~�T쏞�v&�=����T���y/nl��t�Tq�߫)�o)m���R^y����簗~�vP9����v��[+��P�W<o+��������^�׉k��OWiUN?#�`�x���~xi����ך�̩jz}5B�]��7�W��`�՗ZI���3sz��#���X���	��f�=\�Em^I�sMI&���wenk�䰔�Hw_K�Rw�ٙr�3.D�߻m�rX��龔�r�e�tv���oU�y�ދk�v�j��D��Yըu��P�nB�u�����{.��*s�!V��Ѫ�[4f���!�L��m�6��t����p���)ԛ�04��:�3s]�4�N�ˬ٧��1�����a*�,��.�N�0r�%��i�y�kv�Q�%����ڈ \�ׄ�oge��Sú��姖���\� 4���S�ٮ�� ��W�=9kj�}����#���z�ǡ앸��-rw�\/���f��=#J�r�E�ͮCW�T+P&u�V't=�^����cs>��yt3�"8/�G�D�dlo���]Z�w��+�6;{����7ݚ���	/�        :e���n$w�l�j6�זx�=�9i�|��^^Bu�S�zR�P4�cߒ��U����	��a�O8J���^%�沗)(�4�s���b��ϳ��1ˋ�e���n��"�*��xN庰�:7G�!���h��
�\qUܠf�G�����1�{;"s[K��/O���nf�����#�噚��.������`�o*e��N�R�ڠ�+��go���TtFG�"��/i�e#W-�zs���}7|W���ˡ�{�z�.˃4��D�Z���zQ�=:�������"�+�������(v5}$��.]#��da�;=i�k.,��.�	�uyF3���m3�j��n5������iZ���mJG�Zk]p1s��\Ӫ�͓����٥u;��źF�&ܣ(/3t ��   �4 ��~]�|�椡���*�CRj
�
 ���P|K�J��JbR�7�M�Cm`�QBQ���r����� J��]F�d!���1A[��j�7�w�\FH|G��R���s9 �d�&�s���m��D4��c�|� G��6��W�����8ߩ�|̬v����>��E�c���ޛf�c���;s��fo7�]�!䐿]՟c�W�B���>�.�:kN�d�����iK0�.�gkOJ��R���4��9���ͽ����T��B�&B�]�kᎿDc��<��ۄx��s^r�k�b�Y��|���ݴ��tr�-$&�mY~�ݑc�sǳ��m�ۚ�9��FrDM�&y�)�A�Cאi{�D:��TL��ڹr��im��?.A���^7j�o9`��욃Y7S�%=�gS\���<F�t]��jy.�ԧ�r���/E��~��ǁ]Eo���J��H�z�G��3�v���%�4��o�kXw�{/N[{?O���T�>�xJ�02�įz*�\��94Gѻ�L�E}_UWު6�!5@���P����LMKvʦ%ufOK�W�^.e��a6�VoN���[l!��N�޻�H��t�;)FkC1'We�NgU��Ҵ�=��PR�Q��Z�%�� +���͠#��@&e�[�,}3�W�/8	ulߢ�&E/{�� t��n�3�,�^�1�)Oce����%���	��l�;��Sc��nq5B��g&�m{�M�����z7��4�o%=�N�k��ԓ�e�]I��<�I{�nz��v�׸�jX�>�HZ���xuAs@�p#����Ux�v\��ǫ�E� 8CU���/�{�ۊ���l� 6�3#《K���Cf��UM*�L�H^��b<���o3{�f[��	����锕�>��FX�t:׋�i�]�w���y��ڂ%<u�s����CoG^�����a�B��P�V�Q^��%�t^�b��2��C`��s�"�t��sz;����(?���*�yxey\~l1~�d��w?C�OV���[�L���U0[K�P��������<�?d�QRNfLq��0�[�5.��s6mH�3Y<I�ѫ�S>��.��3jjU{�*ɽ�������r���J�X��{�R��Z,����:ri��BW�ӻ<����f*�L��!��}Xf�(n�`ؓ����xvc�]ܕ�."rC*�љ�"�u�S;�}�U[�1�} �����������Z���n��I�p4����y�J�$P�DF�ɫ�K��Eu��K۬yX�������B��-�ݖK'o&���{ZL��Z�E�����G�/Yp�9ax�U�3�/�|L ��.�dB�{i�t3���GG8��z���o��\Q�a��i��e-�9�R��/�`m�`��"�x�T�i���?ky�\r�'�W�W�n�{�����cޙO*)�^���+8���]n��}��mOx���;v2��s~|\��p%�~$�eC�'?e�W`���jәԩ�p��t����[n�Ŏ:=���k� �7�ɻr$s��[xEL�{5I���F�1q��_&د}U_U}��m����/�U+��	�=���]6�I n{�l���{�+��ͣ�Jt��++3;�o�)��!&��7k�;%����D����Le�w"�e_C(��t'�����M���ӐE�d�h7h#՝-�3-�E�^��Ĥ���2�Hay�V��$W)�+T(���Y͏{}�k�~���/5W��5����Xs�|��%�T��\S}u�Tw|D9���U*�s/ޥ*����=ʥ�hf�/|D��ǘ�W<����9�g�".�w�fe���ҋۀ�x�˳l_�$`�Q�ne{7�룝��5���ԃ�
�e'0�4&�>�[��I�~-[��V+��e+�9X�L�-�Ab�9I_�������r8'2�y�ھ0�|A�wU���
�h�&��~Y\�])�Oy��Y�1r�,\�y����ɵ�Mq�!�l�J���ϔ�Yqq�u=����.��v�{^k��S��Q	��+��7x�Q���x�w{ٳ���/Q�X�<�Sߎ����5ߟeSb�jE^h�.��D�q��Ф���Y]nk�+�6{f�Q�&[$`��oA��Zd�9�-�j�r$�H}S�eF*�_m/t5�+浛˻uٞ�s4�eXʕ���~YE�9��F����UW��n ka���ž"٥�-b$Y�Η��0,����]؞rk��7Ҙ L�"��"ݵ6\^8`�:���0�71a�@`v}�������@���떮�.�wa���AX�Êޯi������O���ggb�o9�� �Kx�}���no���r�I�eZ�{ʯj�=Q�v���������<�3Xc~�>��7��{n��f���G9�����Z��'�^h����KhAY-��4�[HdY�-/z�dZ���WA8=�[f�r�G&sv�<BJw�mv�h���Ss�W�Z��K�fV�܊~�m�|�}�eR{x���w�+�*M�2�A�*F:=T���X}��W�9c6�w�ۦh{t|���&�G���U����RG.jfd��~2�1t zEl fIwS:`��s-|�p8!�k�����RX���[�}Ͱ�4���T������F� ���m�e�N/�:�ͯ{��VvtYTJ���`I�W�g[ D�WT�ͪ��>�5�ˑy��rLs��Wr6���i[�*ʸ��W�&����
��r��h�lm����v؀�\�v'9�Ԅ�7���d3�Z|�qR�ԑΨ�Nua�N%�e{�MN�.����8o�"��p�a��޻���=�:ѻ�3v�^��'�g�v����*�~�WXZ�b��Mɬ����2�y��7	�;��J��n2��׻k(R5������Q�veS�Z7ј�h%���2���[4�[µޥ��]��;j�D�Z���1I�>�wN�[�]����=���"�-Թ���s8C�󦖨�Ilu(7��h��|B3�2SNU����HˁJ��ڙC���/Z�/Š�f�vU^�{d_-�p�g����oƢ��t��SAy�Nͥ�&�])���{r�M��o��Z%�z���&Q��ko����$�g�ɯ#��.��Eu�F��������t':����S��Tb�H��yǋ�K+;����DJ��yvN��M���S)k�a���X���1]aݬ�r�W���ǉ:7mt���+1Do�6��
ˈn�V���j�S�i�7��a/HR�����W���*�$ݢCt�A7Tk�}_WД���>l��RPpUF�L��y%��{����ׇ����2�<�hu��tM��Jo��V�c��k죅Y�o��n���?Zr�>d��:�2kv{�ݓ#��]���Ņޤ�/OK�C�kK�yϷś�KZ[-՚�jn��$ᔞr�kE�Ԣ��Z5u�Ow!6jZ46'�g��v�Y��(E��wָL=^�2��Īίnfа1l�|e*�&�n-�F�F�\�[�=�,��Ÿ���Z�=�skvon��5�{���� m ܐ]����i��o��]�Ŏ����S�QS��� �� ��\��Ve�Z-@$��*J�\��Ӓ���΢�ab��=}R�`t�{wF�cL+ˁ���j�+�4��ԺO{>�X�\{�y�f���:����Yζ'��ה�I,�����		��� d�Cf���љp�]-�{V%�P�m�Vl�9*�5� �q<1P5i��ϳwC�{�eĊET¡9�(����kWDA��o�f��k9��3��UD]s}��K�*6��l�������*9t��M�ױnu�_�4����%��@�����؁�\Y���]I�˗]�v30�H���6jM|�gPԻdm��"$g'h�3��s��J�f�l�{�����U�
d5�|5c�����-�7�e��5{"gml�k	�{�ҦR�NQ�Q�o~6�u��6~ϡ9��\�y��         t�ނ���:f��3�J��3�J���Vξ�8�uuF�St�b��Z���m\K`���t��_>�N���u.'cT�ʉR��5���X� q(�o]5�j��WL��9k ��:A���D5�N=W����.IY#�+'Һ�MI{y(�y�������NFV z�����%�
7��@*��U�VyZ�����|�3y�m	dZ�Xw�iܼ�r�K�X(�t���R�.�)����2��:9+{��.�F�Ыոkn%�vneFfƺ"R�T���o;�Sdc�$�tG~xe���P�v�0��J�c��5^��s��1�ڤ��8�GXW]������RC;�\�#jv�	�u�ù�hy�0xf5�Rm�D�}���h]^@y(8��Ȫn��h�0۬1I�O����.ň�8���mg   q� ����w.%��vfS?�k��CS�Dd��&�(0�CRѩ����qɦ
d�31����[la�U�9�E��r+Q��`dfe�E����ط��������lp�F0e�@��fdeV���mq�� ���2��QM� ��Q�γZ�%w�oqeQM;�Y����o�	6��r�L������kh���2̬�ɥ�� !@�"���U0�/X2or����i���N����E�=0QQD�/bH�ӛ"��r��{�~f���Z!":Ǯ�צI�hRuq����v	��][,�dLnآ��V��mQ�
nV�3/�FT��{��{�"���Rw->����*���gYP"���:��˾�I�+���T��c�g`Ut
�ڡw�7+װ���o�(��T��V�'�{���'$�-{4U�M(ڽ���������Ir��jHjL����2�;U�<U�Om���L��H�X�|��b��Ϲ-}�uv�*��;ި=��s�Nn!������o��>�fM�׆.��Byk6���r������X1틘,�Ǉ�L�<�}�R�Ɏm��7��k�Ƭ8����f$�*��ĴMW���}��7�%ޞ���$�vX*�?�g+�o�v�槧�>'���\�)ĝuu.�ĳZx������u�u&*�+SWS�ڼ[� uFs��kW6��wJ�n�
J�s��?I蘱��!��<�����aө]�mv�i��P����nK�nf͚�1��3�[�4&�lE�VϷ���=�>�9	t��y�K;�)��x�Z���`6z��i6�a7i�m���^�S���������]��.���V�kg�L`�;��y�����K4�3������}y0k�}DI�!�t�:���޶N1{�����4<fз�j2pt2u�!��`��r�O+S��1D��i=x5�e�hoo����R�����
TO���C�f���%��yX���i̭i�۵��K>�ʃ
���m?�I��+��{��}����'�x����=(tg�>7�ϳ*0�����yC���r5���Y�t����%��R��U�]=bj疪�Ilu2�}�H{r'�xܙ;�G��<*����쵢L����$�м/J�ra��(NY�ή_����i�f��'\�S����9&u8�Ji��K7�7����^އф�Aj�m���Tg[�����0q$���Ŭ[����#��P@"���^h1eǇ��r���Z���Nچ��%��7�� 3y����$"g~�ʝ���-mR煜�}�E}��&����E��r���l���uv7��������1N���Yӑ`c-��c�t��Jח�(�Y�IkՉTK6��^�ǽ=Y�-�4-�=k��`U�ʴo0p�8r�J�#f��c#N�k�w���rB;�ܯ?6w�[���5��,�"��z�vw{��|7;�r�i�!��O�)�����w����{;�CXA��K��Z�J8�Q�rOz҅M1J��b\}��)�6D/�C��,1��*�����җ\(��v���/�l���}��iLic��Z4��8�^��!�Ѯ�ՅI���e&=�h]+M����ݗ�]vɎ=��5����=���ȏ��j���V�J6��d��"n�Ee(��7�rG��3�!��҆���V��侶�w����2�˴�M����^��:}yfM���A!�$e��vh���ʛ;�0�!������	�M}��sT8h�#o�����'�G��wv������6C�D{��D�r��>�Z���%���#o����𻩵دxe���l���[�G%]zK�n��h�W���<��ե�CW��-[�>��F-3=G��3�x4D#ۏ�ǂ!nm0�����B�c�*���y����i>��+�|a���㼡�}_n�&�&��#(#�D���س��w<r[���
�W�O8N$V�7��/,ZK:�����]�whƘ�a��N͍RT[���;����i�뻂�"m����[[�N)/�\'��,Z����/Q6A�{��|�o1��$�Ƿ�5�$:�8#�ܫ�R*�!�R %�0[q/���l��v0��+Op�H�,�j�[ �c:� 2O�/��/�=�9j����tĆt ����=k�Q'M�r������>���)|���
l�%�`���Ŭ�m�)y.5�ŗ��=��Pޮ�zp87�a�ㅖ֙J��,ցz��UBj!7���n���b<�F�wp�ѣ���g��c��Zg��r-�2*su$��*��.Y(ONΣ�)l_A~�K��S)\r��I�,���EG��������\d�*؇�Q�n��s$�'Wo�r��/�d�>A���^:k-ѫVe8}{�=U{'��=���5�c�;)�k���E��;͏*.��Z�7)k�sA$��*XU1G�(�v�Hƻ;�^6�РkF�u��49HE�'O��ݷWn�"9M��%Eof�Y���e���`�{��\^#��iωkt��v�����]�7l4CZ��vT;���6�+��>?H�hs���OE�V�c����<65E�Bֶ�@&]�vS������h�<�ֽ�����V�W�%�˫龞�'}�	q�s��x�KL���!0l�!�C��uI=p$Y�Ka����CpS���4�Zv��j�}�T�ҲnϛC�?�0��a"l�F���d�����NדԒ7A���:|7:���֡c[f���B�V��/|;{s=<v#����L���'�=����^v��h�.����j�O:�F�YA8C�/��DC�:p��@����2�ϱ均�אɥZ��C�c��g�� peR�B;��3����_n�9�_P���`��fIl�p�ڗm�hO!-�lI�i�]�R����v�,�̈�mfEƎ')	й�D������=�}�y���h���:lcBκg�1h���c1�����{���ܼZC^m"0ҋO�o��V��Q"���b��OnN���45q����Ɨ!0h~$�U��(�<��I�e^ox<����ҍ�<�&/���!�4��T����ޮ�"�N�����-�7�L��T��#mXm���qw���knIۃ�Rj����+"P�4� �q�Ʈ=jZ�N'ݾ�S=$n�[�];���Xb����<X���S<��	Ǝ�7�;�����+1Ѱ@Қ�U�C�Cu���z��f�0*�oJ�7�NVz�Ӯ��)G��/MAk.����M9��Y�.l�u�z?_sFŦ��\FlbA��g��p����G��T8�]��'���jݷ��B������;}\��=����Z&B����J[�u!��sh*�2O寰͸���/W��DV�@gH���dfh!�J�룜�|xח�7�Ð��:н��Pڧ�7��B��C�PH���D�\gڂ��w�h��G��ӽ�'��B���x�>$��MC=l��[ZX����\M�ϭ������<Ĝ�DI+c�-�>�	����$Ey1i�>U2M��{͑rdd��^�a����ǭAY�ZSܶ�o�`�|�:�d?���!
ӡF�	�p4=ٟv�s����n�{�'(���I��@0�x�&EE�>���T_�ٽ�Z�,.��W����=A�	�L5���׆��{�S=�{ޔC8I�l�^�� �K��E�^�3Q>/�J�ܑ�Nk�ΟC���h��ay�V8k61a�/����Ɉ�hg�T=��0|���u�e�n��5sN.�o7/�����AvLyѱA����vܝ��Ȅ�ޟZ8�s�DwWԫ��L�&a�����}S�E�z�U�b�qe~���i��\��گlZ�p��%��5�r�܀����z��5�78�F�� H�8���9�F�N��9�'�����O1gڸ�9�y_=�ġRW��n9]V�B!��H�;�=�d,�O"�����V���J��P������rF�0�P���K��<w�Z�_��f��l�g32I�>c����I�p�HĆ=1���oe-^	���DW��D���8�:|�	B�Ai��x�'�$#hj"���h�+����-�ۇG�L�4l�Aג���^���zpY�u
´ᇈ:g��Ń�lHx�t/:�6��ݞ�
׷�M����p�&x�x�96>��[4��io_���XW@�eZ ��4$�����N+jʨ�]t�x���d�[�Ӵ�+�Q�>��6����G����J�оH>d�V�u�V��r���{��vW:�ii{٦:��@��r�.��`w��c�=$���s�k���\�����.Z��Ke�z���(������}'1SDH�R��}��qK��Lj�D}����r�<�8�sU�n��/a�ݰV��u�Q�Q�.��wC��bJ�1���4��i��
�h\�\^��jcoz͛��uu�R�OA]�f��v�K&�����kD�Fp��
jW^�bOxk�-=K�ق��F��.��\�뙔�W(����˄4�� �E�)'5=3]^�;z�[6mY����ki\�Ս����x��R�Pwo�άx��Zx��SR�N��LэC���(� ys����Z�Wo/���^�  �  �  ����-^<�ٙ�U����\kx�#0���h�ff#*s�F�qV�v����n#�h�!��s8�&섔9)h�szf�.^�!��|�f�Y���Z��+���7���ٖɼ��z�V$�,��B���Z&U��j7-����Rp��NWr��V�Hv2��U��4䣊
5��Q�ed��{�����?;)�/*��^�����n�q\v���j�艙ygG<�k;#6�ۮ��$�"�T�k���{�W|�EvNf2�Bڋ�F��O0��,,Q���ёS��ed�z�q�-b�1(8��b-�Zx7r�s�U�b]��}I�Z��Q�;��}����70'L����L��g��	��6;�$�/~�^Q�j%&�饠���5���\c���dna<�.N%)$���$�����g��jb���ڢ����Ffm8\o�oojw*Ԛ�MZր��a�m�հkZ�I���f�dd��4dZ͵����:�Xo�SN�lh����փPeZ��e�q��v��Z1ի3kmf�k-NM4m��4f�h�4[ٴbQE�[�Ѭ3+28�Z�,�|�(���fmY�Y��U.��D�Q��k2�edXdW�Ñ���Q:�32*��6͵�m5��Tm�����j�e��[[N��#+00���UV�Q���m��Fc�do�o�)��؇�J$�	��������u������l�s��ۼ{��D�}sy��!]Z�m�T�tXo���RI v�w�̩�oߪn�oe�-��[%->�L�;�[�Y=F���yS��wqV|7��Hdx鴡n��^C�I�
�!��k���;��>�|�J���/`�O�;�8�����٣͞��=&��{]��6"�s�{��BEx�.1���J�I��7�J��r�F�yeu�.�
v��ZZMS��+��C]��Ir@��
����ԋ7�N��+���C��C0�)��6����a4Bu��Ӳç���y2�Ap.�ղ��{{o5D���-��8���m����	���8�^�N7�L+ڬ(����]{��Bb�C�!��J��Z���Lm(I�2�03��oE����
�"yQ�W�k\a$�5��yZ�M���>[��^~�|yޤ#�)r���ZNr�%LZ�;�#�n���Գt���[$G,*ĽF�t����i�SWV�I�bM�˔����$��ʮ�����"�G�-i��GM���m�+��{�;�2%=阅\G���C�K�ş兟�ȑ��G����Vb���{�_g��cj���HVRp�":�h#"���t�����o	Iᯈ��W�Hڳ�kC.7�Ϫ�ŝ,{�ooo���x	̝�F^~!�}x�Kҍ�E��|:�^M��Y8�w�,D�,^-!�6�A�^����2=<������uU��EC��:�O�@^."y�e5�K����u��6�ݺe�l�!�k�H+���/��b$]k�b�^,��헞������q����^C�dD�\wU�{V;��T����U��z�5q�lq�&�lC�0�Y��=��iD'-�A��U�-��N�]yNEo+�[��\�]�w##FY��.�[g'�B�i(l�N��AdR�=�v;Z=�2gI3����YQB�����\c~����F�����
��2=>5���&���mb~��Q���cn���;@�
j�@��j�2��kG�<�:w�v��[���<kW�ys����D�7������z��8��o�'ۮ�ǧ��Ƅ�r�\Fo1-,?�q!Z��D%)#]��̷SNVD'�Wr8��tFl2�O��R�9D��%Y���p�#�H�������Y�;�R�O�[*1��6%�*�K��.�����P��aю#}Oirs9��ٽz�t��}I���Nh�I;���o��[����4x�)�<%�s6���Ƙ��A#DC"$f��hj6��9�k�Cu��Bw���Y'(�
��L��x�k��g4����;�0����5ni��c]�-�
���4�e��f�͡�N�D�����|�f�.�E�7�F
���v��Z������ߛ�֮�!�PO?�����W�0�xޢc	8II�x;,J���w2��0��B�����8'0����Td�O����7�ν$�v�>4E�N��+��<�,��c"wB�~��*��jc�vO���ɇ���=��b��Ç������U�}��ԛj)���Z�"�.����O]��-1u��gK���b�_o�î}��bF�cC�;[6���Xt���ܶ32�,��d������:�c��}�Zޖ��@�>�xneyy*�Y�+��������Jk5j���ǽ��r�g�\����ը;�B�g��R�j���^|}b������fE��j��N��z^nt��j�U��p0�fO�ٔ����cϏ�}�2nL��W̗���&�^����u���޼J-�	����B�3��/h֮�8Nwn���C�{+���p�H��������{0�h����B\p���~��>���D���Y&-=�R���M�_Y�U}��ߍ^r�U����F����B!��f������,3�?w�7�Ix�g���������4��=���Vi���~��{��|�L
�٥v��������g!0��%��}�ǻ�0�?#��"le�1;@��jO	<Q~�Ռ�bRQ�s�6�<л��9M�NؾW�.$� ��>�c޽�{ӻ�}�ė��ʡ[mZ�5����)�km�3�&���1{:{�)��er�<=O����;)b⠹�8�.�܊Oj���1���1o�K[�ld�LCQYܛ_nabTs�ւG�������^�������[4s�3P�C�=8��^�7-O.=f���Ն+�î�m�Z�M}���r��2w7B���HiN��5m7�G�̍�+1���]�*�	6Y��,��]d�ԈN�����U1k������-�{��G�<�Q>8�r	��.$��Xͪ�I�k�u8��d�V�Ov��U[�C�4�Ѥ���>5�Z���k��w�M[�;ý���2pi��+��FC	6����^����$�!�{d�}��^��3O]�V���{Pָ��&�Jr<����Ҟ�z{꭛'pJ��c����i�ڇ5�����P�yL�\����G|��+h<|.~k=u����l'T�^�����L;N��a�>'x��Ǫ�����E��5�L3�YA��e��͞��}�a�h��w+ƃ�m1j�0y�uf{ݫ���5�g(F�O��0�\�C���f
f�b���um�Ǯ�{�OF�c�#N�$��i!�`^������4]�=��^	3�o.�+W]�]\��o(qU���>���y�>tk��J�-����U�G7=c�0���W*�7/��I�>o�^�}�����ꗪ(Mo7�t��y��8�{�]L<O�Y��^�/I뉇�S\��ؑ���k�ƮK��wa�,���A�|Q�C�Bb&���kor�ґ��}�����ܽ�{�y+����B���݌���=�W�
�-[�X��QW�}	�9沩���%�y�FIGj�ڐZ�������~#ƍڴ���x�x��->,�qA��ϸ,ڒ����ǲ1�t�=��}�f���T�yCu���&=�M���c�=�MS�Ǎb�i�����_��o{�d/�ѣ�3{�ё9�\��P��x�P��w��ݝC�|2�&��&�����u�]d�\�(:u{�8�jS���}��^2���f���V{Ӻ�zy�(�{D%眍�1.����hCSI���&K� #���jx�M-��T�n�_S<2��֬l��;9�p�;|#U	����
'��q�*��7S[��쁹@ag�:w�����Z���!�L� �Oæ(C��Ho�t��T�-ѭi�yޞZ<���L�����I'd'�ҹgr�_�΢�\�D��D;Sj�=�(5q22C�/R���B����K����z{��p�U�C�4�Cs@�l���463�FJVb��h"�VW�����7��\�Luq��`<sQ0���]�y��鄉�g-�����8וyg�s	��x�L��ǁ�>���L>�>!��j&���+�G��\[�!�7�h��ڞ�h���]
#���^�`_`�0~k���W._^��9��e���#��N"Z�Jgi�E	�=(aļa��O�q�7�=��qCgԍxcGj�oy���X�~UK��������n#[�.��7�&���ǓnI�OwI�{(oKӡkw���<I���j�u��'1/7a�h}�G3c�*�@l�μ��Z�E�k*8�4��o
�@H�g���h�����4��-:d�,���2���Dq����0��}�)PHB�a�$��V��a�-��OX��k���2o{G�vqa�֋��K�4#\�㼬ȴ_�W��z)� �{}\�z*���e�.�Z�wf��n��?��׳����Ϊ��?j弨�m���IB�s}���V5�IS.���u�>�y���/0F	B%Z�[�}�W}�7�:w�`~���P琬�>:||s�ח��q��g�w��B}�Ð3�P�����F��<Fan�g�{��Y�Ǝ{�ӹ�>�d����� �c��;���
`u���y˗糶
)dC��(^Ə���J����)� <���3�/s����=��2L�\#�+�\D�"�0v7���W���geZ��rl����7���ܥV6Ad9vUr�w[��$��?-$�����W����*Z�rw�~��ݶ�K�Y>-sv��v���󳧆f�VsT+W=O��^.�z�)[Lq&|��c���d��r��~�2�Z���1e�d��1��M��0�9��p�P�Tw��ݴג��J�:oƈ�	�r�,��0;hK��L7,��N&�zIW����@v@��V,�~�vGŌ+v��XԯW�퍷[���ٶn�xS�D�=�|j/�V�K�>�:�l�p�C|3+�i�z0H�M���%o
��-�o��E󕎝��|'m�x��9v��.0�M�g#�A�� �Ƶ�/I������K�"\�nZ�`\]j����FT6�+��{�2A=+ԅ(�h��k�f�|}��M��#G��0'�׼�_�4��utf�N�,�3�E����M`Vzbpvm'+4#5AjK�O��)mh;��q�ՁVs�����j�b��Es��s]Y�J���m�4��e[�uk����C�l���\C��&#YX�-�Y,�(��*�`Ɋ��p|�Ѻ֟1"^u�\Q��ꕐ�T�Iѥ��CnX��[�yXn�����I�4e���V���p����������7��-��C���2�����d�PVn#�m�{d�A8������8��3K+��)>���İqQȨ�2SZ�S�qB>.8���yia��U��4+������kG'^�9-��PmK?vD@i�����̎|E'�+#�9M��[]/N�Mnػ�h�Ñ��gW���wL��i�	�h��~�q�����<M^xuE���>"��5��wO�QIs�L83���ߩ����B         ��b�F��j�����nE�.J��{cU^��f�,+�4>Ut���<>4�0�xu���!�۲��î
i�k[kQ���y�M�]f��h��4�C�2�+���P�p�sf�ف\i�G������U,��Ƕ��á�,H*l&g\���w��tUu{�&_.�C"�'JAH�X����CEpIZ�]7�tރ��EUl��]��dܬP*�W5C�H]f�����N@�;�G�x��ض7�8���DL��d���vӣ�����D�Fv�*
�d&���6]��+q�قR�;����U��k�HU��B:H[��֦�WJ�gX�#9:��\[0�nti�ݖ�%\��]��<�I�M��`�w��dO��"	>2�ɿ.ZVs�Z���������ӳ��7x��   ���C��W���a^NE�y&�e�mkVDdffZ����Y޵���QZ�)����i�fmk��5eok[�ؘ�md<leE��ma59a�2��H��m���"��d�A�5��ѭ�u��EPU�LQo�14�FDż9:�\F�Qma����(���
h��ńM��oj�'$֬��H�1�Ձ����F��335EM��PUAI$W��i;�?鹺�{�Q������s {��y>x�
�f��@����d�,����`Ԍ�������>2ז꽯j��e|�#�ǖҍzEo�N��`#O-/#o�%���CDq�xТm]�w��C�C+MY�y�����Q��w����K�h�yx����0̦m�=�c��Y�<4��x��#�L$ԓ���#�/�u�=�?%���q~��E{�0P���&S\��iYӬ��QBս��b�m�T0��T��c�|��8M��Bҭ�o���
։u<�.�ئ�ױO�qP��.P�/ʁ�5)�ݵO�t����<|"�㔑�⤆r�P�ʡ�M�؇����v��OxYIxj��V;��˵iuc�Ņb>2�����g��ݧ&�qyD�P��m�Y�5ɵg��T�k�9��dC3��Gk�,r�ZC�%� �� ��O;f0��}Pׁ��wG���UH!��^X)�
��ܔL�]|���..�A��&k���i-�����y�K�;�%��I�oHcщZ籏դi���¡�B+�W�o��M��ݘ%�Ux����|e��W���r�Fs�\F�b�V�k��JI,ש	+�_VfQ��~'%��[�!�Q3�z��i�g�hg$p{�=I��r&j��5x�̹t{�{��?{PƳ����|�æ(C�c�!��I
�C��Xz�6w�/O�vP��\YG�C�z�b"I�	�&GUr���N��kR��ϯYE��=C�ia���4�J�j?]��	���)ǧ��P�!��<;s9qr�Zt(�{���KrQ��}�����O��2�0:I��������#��DH�Gi�hU����k�E��g �=^>Fy`�7��%T8צ�bCB&�fN�<�P�ClG΁˫
Af���>�&�k�d��`����zuF6w!m�ט䃗 ��8I��T��VW*u�z�J����M�;�feΞ���k'�c#�2��N2���vƜT�}9P���1]uv� l�l�/��aP���s=A}V�\ǱB�2D���vw��|a���B�_'�yh��Uޔ(bļj/�<E����<��$���e��q^�
���R��9oybm4':����:{�����k㘡,[��Pó��_{_ˍt�ȥw������$�YWNT;��ZS�]ڢ&��������^tp\���ʭ�����V��8N$p��.|}tĤ3۲}"ߺg~Œ�w�I5V2��c�c5�8�8�+L$�͘��&��|^e��{��.���<�;��I��K	0�t�lGW���[{}��ׄ~"�/8v���x�o:����*���U��b����c�N���E`QJK�m��,�W�m�W�{�^Z͜3bus苝�#�@�'+��jf�Ӷ�a13{UXƼ=��W^�_��@e�4��oy�Z ��qP���RDs�쏪��|t������9^���TE]��#]�S@�^>m������������2�p���ht_W�w}�Hf�!y(w���75�'hL{�Q��|���I�x:g�F.�<I�9#�5�(�aӔ������6}9��ߥH �AW;�Ĝ�[�թ��:1V�er�qY��d���z���R�'e;J�L�Оo�2.b���E�͓�|`pMy
E�}J�rf�LhC���Uo��]� 9��{���l�l���j"9Myfi��]�|4�>�2կ+>�,:Wʒ�P��!��q}�03��V��u0un�?�}tщ��Lt��'g��ƌ<e'�%�Q	Y��ȶݼ�dZ�CwF�+��B�>�b������3��E�+2��Ԙsy��(��%:㳺�6��J�%�&�7b� ϙ��]�V��8�5�$�ذ�Ų0�Ha&��x�(+f�)7ݢn�y?z�]�"��թ׈�B�NXFh\aa"l�9m՞�[����+��x�Z}��*�3���S6��Ta�گ�.'�i����E�����!Hx�q���룳[�=~��=�;���;�S>�0��-�9�ڳ�0+M�tn��2+�A�:B�T����>��%��!�㮼hQ6��;�L�&�^}��������;���	�M�'��x��0�<��Yۛ�:��#k��y!z�ic6�jP�ӗ�Ɲ�����w�+ˏ�_$T@�|a�<�a�5�K�z��RZ�'Y:w�"�k�R_�R��1�c�Bn2CP�~�7���d�ǃT�c���l�˹�s�G��%�,튲���v���{H�Q���=wr�krk����@�n�!צJ����ƚ�U�y����"��>��`p*m�_<�ރ|����Y���ޘ����ג�ށ�;�6a�H�Uk����<l�5�GG�j_?e��ӅP�F%�^>�-B8тե�-�^��Շ%��dD��)��Rݛ�|"a��<���ظ��ڳ��ڪT�B�˄�+tH�u��j�yޮu�t7f���^���}��7�G�9��5EG�� Gʘ�XɬP�=_s�6=4U�M��lh&Ƅ��{r���I�;�2�(C���ci�b^<}v���~~49f�7Iʍ�ں�FCbbGOM�->�0v�\}E=I|��3W�A�R��;��t,�ތe/D3[GbF�i��u�T߅/v-t�l�	��ޣJbó����q�I�y`��a$���z�$�|R>ؼ��|�ָ��Y��\�Kx�uu�����ݤ.$�X�z�9�J�vvV�EW3ъ�2�u�����^�OF'3yŗzU�H��f�h�B!���q�g�!�؁4s�B��B(dd�ҵ*h�}m��o��~Vv��Ɓ�N�ǩ`�Cǫ\<D"x9o�E���9�{��(z���^�����o��KϏ���[��~�^��{���K>�H׌�h�k_j����֥����OS�����$+��q*2x���d3/Y8ʆ�_ ��L�!��C�k7ݾ��G����K��r�YP���s=K���=���Wv�=Oo�ϫ'�-r�#;r�G���ޔ(bļj/�%��u%t��"-{�4Q�bc��-2�f�#ا[��\�(��:g�S�^���h{�"���aB:����ش�Nb�}�|bu�5�W�}<e������"F�}�?��_66.X}d��ƭSM��j�8��ݕ��qrF�SY���]Dh-�7SK&�(v���O����<�k��>9\�Z�h�Q��Hm��5�y���U����S���)�.5���;�~�{����yCk/>4>>�b:|���@;�'�p���ԓN�vKy	�����V�i$����A,2�ي����{d��g)��~!U�ۧ<���rj���w[�y3[ero�U����[�Y<��\EZ�|�F��� Hk:aԪ�]�5;��cnZYMOD'����it2^!��ұb����mI�q/Fl�Ɓz�몡5W���������2�ns���^�{���|�C��M|aZP全.���ϕ�yP�.�_I<
JϾ�yw!�L;����H�%�&��V�mC�ܞ0���د|���hC�	3Q��IR����;�+�U���|�9I��fV�+W�>5�c��hv+�-m[�+��t�%�f"!��ׯ�c��$��k2����n���u-�KY�����+���$��l�Y
�h	�U[V3!�6�;#�:���s�r�0�Ç�"ڇ
;J�y
0ld�)�a���7TM��:��R�
>Y.�	j�&���2���i�]�Q3�tV�lV||$xs
�"a���z�><N��������96e��d��ҝ(N���&Jvh��a���Qx�/�oT����w���n�z�CZV��(�Zd�<��h��I���!�G�K��5j���A��9i��-"l��Ӊ�>��7��h��GNZ�>�o���+����0ɼ��<_��	��a'�VsƇ�����>���13j_V�_�VM�-"�HZ�>V�x���s��(^׵`N�;S��k~����aֻ��<a��lH���CDu�^�J�_h�(v��dB�û����%*���K��n�Æ�-�.�m<�"�)6C�뼨����WTB��먷�I"��qk�"��8v4�Xf�v}��њ.L>��d�JzL�!�[��%�4a��?��=��mo_�����3�;GW�8�D�x���QZ �W4e��oػ���r9��Uk��ƹ"�0mq��~���Et�fn��1Z�9����2!�UJ�<A_c��/��0�R����H��k��5���_'��0�ԅz9Ӳ���&�9�	��׊�Փ���D�\@_M.���Q*�˭^��r�K����8A��ت^>J>�-B8ѣIN�<Z�
��"#��9��듸D�{��b��<畑�{���� B�4����<>��������"��|M[����[5��<��ރڴ+5#^��;C��qu\�]�[#�G8��ŧ���`b��B��>G}YOĸ��Җ����*�z�v܌˥�����.��
��-5��;7�k�N]X;��"����vP�zI�{/[���ޖ����k/ۉ��"�r�kvT g��R�R;��yB��j,���?%HݹZ��S�J�4"A
�$��@3���/$:㽡�ڷ�Y}u��D�`}I��ķXC�V	��f��r[JP=1f�c=9�d������>k���iZ�\�sH����E�k�q��qk5+ޥ��A�E��T��WK&�r���>8xV�w,#w[�A�8U���₍�و��U]N,p�ԻIXn��>�w��0�͂�,�Y��oYz��-,�����Y�禝\�q l�^���������.ɘn�lg&{33s���SEiJ8,��7V�)��E+�n�˴6���s��	/�f�K�z����*�en����C}��s+�=bMܭ�����'p��)q}!.v�P�x�]�w�������         ����f6l��3�k��xy��&�&�,�ͻ���]s��ws)b��s��t�Pz\D�D�wY���9L�����Q�{9�$*Q�Wٯ*�*J��з��Z�h��XD�B|Ȉ����u�W}�7͕�B&�(wt���^�P� l�6L#lr�^s�F�o�+�f� �X����c�uk���t�&��WK�\s5ID��S���w�ې.���*.7\����M�s1�c96BX�w2ib���;B�f� ��#6�D����������[����4��q=�gb�s%�8kR����v��fܲ�-In]�Fw7��[j�u t%}.հp��s-6�����jܽ�4Ev_qhnb�6��0�����|[n�{�r�U��VI�7��U���l�p  q�wz]����0��(��X��(��(��5E�cla��f�"�&#3(��XQ�230���*&�mi��2�"��h�S�A�j�c�h�j�2Z�)"k35�4��ֲj�*��3�32�
����uUq�ư�F4F����o�*J�(���ES�2��,*�aRj5:�ՕQDEET��T��Z�&ɷ�Z�"������Y�dA3��3QUDY9%D5ٔU.N��:�0ɲp��kk
��E%$EDPE�D�hA �I/�TܣW�y��i��[�J�Nmv摍w�lqi{��K�.�TiF�4��韛-�K4ײ���G]뮰Dq@�_��������^������~��*���5)�<��x�CORD,�L��Z3ގ�m�͓���g��1��ԑȑ��IH���J�n��Y���S!��Xry�wˏ
L��{�"�$���9vGW�=�~�	��8p��H���Ƅ�F|�
/.��Ż rw��Z�=V������'_1�x�(��p��۰�ּ����>�8���J�U�����߽\C(�=�,�9���'��PH��H�#���V�b�O�_+���f8��[����	�{.��&"x���5���o ��Op�����J��x��(W�~�����]�|�>�&W��o׹�^�g�%N��h�h������C��UǮ�"
-]�)jN7����Qm��Y꾈V����v"/L�ϭl�N�n�9.f9�Np��y��\!?ݳO����Ǉ�<ű��y���g*�C%㞺�����N� q��e|=�Ʊi��2����g��bښ1]�+�T�0=٣O���J�����z���=K��s+�V�@��_�ߥi�?�+�5��/�'�-h����>$��jՌx��\q	��;���.���Y�^��5y�AcG>'�u1)p66^�=]�'��R�ؽ}�!�U�[U��'Zaw����5����R-� �2��uK�*���][�
�fS Z�]�N��$�L�Rt��|����Q���DKU|G�Xf��p����/D\��H�ЉX������\oW���b��|^���z-�}w��>:|x��hx�ʡ5P�(�Wq�Ǘ�7��ы���4�Lɦj����Xq�R�/L��9w[f�j���t�����ѵ\8���$� ��L�(ޚP�n�f%��խEU؆̔ :]�������X�4V��D�M:��׍�r��ia(w��/�wCoY��o��C���A圇��>'�܇�:r$gk$Qf8�&�{���V�N�c���K��!�	:L[��m%Jj'���_�C���'�Cﲍ�˖�e���K�%��L���_*e��U�@��&l^��}���J13�-��!Gb'D�!�*�����xe�����C|#�T��P��).6E�v!0kf����x���\τ��.����ݔ�-	C�P�	��P;��}3P]���̈́%uLt+�:GJ�E�>;�sT���F8�u�V-Y�7t�фdCs_b��z�CI���&Bi�rnN�e�~�9�N_��֡����k��P�g����^��փ��64b��&S����:��]�o����Ȭ�+�����s����r�3y+��=��I,��Ⱥ��(!Pn�2�m�R�%C�b<�;;~����	�n�F���*u�S�߲G*�\~͖�l!ڦ�TI}�;��o��0��H!{�/R��>�~"f�>h��t���X_������$~�4�҄�~�Hw����n��p0�"���)sAa݌=���C�q�+Ƈ�V�7Q�{{���^��Fa��&}_F;��O"wy���?a��s0�Ŧ��{^�NMK�4�Ñ$���q!�	#/ZHO9��o��w���:��%�˥�~#�
抈��Yb�y����QI�M��G��27��WDCcʩWǈ+(�!�5��^]�H2}̐�1Ѧ/⠖������\����8�ia�M��*]�c���_Z�/�FE������TJ������K��ڀSzQ%�-�J��e��˾����c;��b�`���e���V��ƒ�H��#�m�Ռ"���I��7��0':L�7߾����N�#�c��u,��د�<l�V�Z8��U��e���o7��;�=���X��D��<畑�{Xm[����v�l��ڄХ�a=��z�4���щC\�cƵi{%l=Չ���v���~4B'��Ux������c���a�S�5�gd]U���ؽ�zy�'J��g���c(=�KǏ��%�٘��{u+�����Q\K*�J}z�brGA��
z�!/<�m5��誼���t��.��A;��g�F2��jH��8tß#�����f�=;�
�C޷I
���a�
L�y�P��a$�w雾���;���xe[�Zp��T9	=�(5�e��g�+os 7�u��C'U�C�d��"�e�x�)���M�°'�Z+XkdT�q6Yhu*�W�R���8mJ[���������KܙR`�����7q�C�wm'��/a]�
�6]�؜�|y��K��ǯ�o��r%F�^V��0����ߩ�C~_TA*����Qʆw�������}�q�:^"F��*��ļ��^Uּ3Z���|Q��3�ì����W#��Oc��D�0�Z9�]�f;��d�7Cq[C֬�y��|��J�U�Wi?:^y�P�VڮVj9�h�y�d��dc��u�W��J���^	甇�"ڀ��2zd_��\�᝾��j����+{7�i�:��w�L��W���D��P�Y������#�Y��qBmi�P��W\�n�	�Z�.9�bG���n�7gNR���܅�ĖsV���F�^�N����z|;��g����0��8��P��\}�ĝ�����o$����~Uk��~�j���fmV�	�酀9�&����3J�
�}�Od��Y��n')�f[4�h9���K����6#ki��|Ff��k�`��dvc��xv��y�}������~f1f H�z�����=�z�����!�r߳�b6��ꓞ�I�ĕ������CԼE�uY�p|'��15O�ý����ޞ< H�M��!�y.=z�w�V�������/+yrA(����a�\u�&��CE#j���Z*��W�Wy��a*8Q�!��i���aI�}M���}%w�����w1{6��^7y/W1�҅�4z��(���	ϼyέ���1��P�W�U�I0A�4��^#�R�;vu�^����'�����)�<hm�6h�T*k�
�3�":�%]݆��tW�Խʣ�W���ǏԔ6Q�-��!F���H�e莽$�Hi������1	�9�I������t�9C[H�ty�+NW�7e�f��ۄ����W_��$x{��~%�V}w��2&1qqw���u�v�Q�n��T +pfT��v|�6��!6�������;X��ޏ�����W�C�x��C+[ꬰrL�Q�~s�R�}���?]5F'yw{v�/�.���(T��wk>��Z��^,�c�-�/UH�	-+KJ�X�7����&՞�1�)�K�b�����x�j���1U����l��x�M� �r<�I+��~"�$r�uǮͦy�w���=���)���#	B�B����<�H��������P�qp�W���:#^r<<i0^�E�4�B{J/kڋ����}3��cx�#�j<u��S�;ؑ+����u-K(X��Ey�Aj�������?���g����Oo4aci��3_�t�m���2��Ι�,�\xޖ��"D/T-!���U��V��4�|���0YaY�-Z�u�Et��jg0��wu�Z4�k�X{'t[�2��7WvGnD(�%�BXw�7�uk7�=q��|���@F�R�������U�?x�h�*�hJޞ��ވ�(]��V-��O��d*�B��ȇ|�����q����}��R��#�k��-���T��2�2��T?<8�S���w	�d'�d=�KO���Շ�RG�Gx�!�U�ˬh��S�7�=�೤g��!�A�u,��+4x�bեև�m�5~����¼<��~z|p��"a���b���[�dD|�L�J�������.`��u�z�:-�щZ�c5�+��>�ٓ���~��J��8���FK�|f({�Y��Wn]��xVQ�����:�����#�Hf=�J���9��NCL�ᚓf��'�|�D2Y>:cBrG4��P�ĐFw�Nc�	�Wό��B�ipd=��L0�T�֥�����^7O���;=L�$��(���h���Tʅ�fËm�B�t��b`�i������8��d�wx-���[k���,�61��!��/�:a����Kݾ���ଏ�c�IL��#�a������=H�9���޵MOI��$��\���}���4x�*hX�'��5�F�ڋd�z�wc�d����Tx���s��q1|ǩGS�S���}������7�����#py4���������;����Ξ⍖4(^�y�t�$m�>�.��|iAxk�𣙫&gz�u{q�^�	��x�#�B2x�\C!���g>��x@���f�m����V��'0�FO���8�c�=�>�\�g��O�P�QgNm�ݾ�8�2�����@�Q�m�R6]Le��3�qĸ��"�]i����>8tȑ����[�&��o��..^.ݙ2�dނ���N&�÷wWR��V(�L9���4��y���&IzJԤ��V�=X�#�eީ[ ��wl��	����sT�8,f��q�Fɽ��A,k��L��"uh�N@�)F�7�����w�zZ�D�.�k�0}�M��d���*v�E9�X�ⲊT�ϱU�].��fJ�%��t0.xT��W����;�;]�A��+�<���t���D��e��[{YG�9���d
p�2�[�6�<dޕۓ+�v�\�uK�!K]�Bt<���Z�D\ښ�H��6,Y<�;�rM��JxT)'�vd�<�"E�w��W1�2&��%�xfJ�c�x�h@ݚ'0e�o2(����K�pF[��t*��v�;S*���,��L�yr���B��<�\�^'����0����.��4�କ4t��%�31R��~Ap9�n��[�
�w>�uݠ�nI         ׍�zj����Aj�&j�Rv�Მ#�wu�](*���	GH�l��Y�p])���h�,���9�e�,�W��ho>2�w�[�4�\Ku��f�������ƦA֜� ��\����кʍ�v�"d��ج�Z�����4+(<�e���1��/�՜�	�3Z۱ۉ�EF�7��]˼�0�V��n�e�Hm�%oS����0ح��Oa��PD�OK�M<;���gMNAE�V�P�\4�W�M/\�����ƺ�>2(z�^keE��i�gZY�=�YPn	n�Et}Za�I�h���٬������f��m��)�mv�3m_Lуu�J�b��T�I��fU�M�(c��uj�mQ�2�6�i��Sׄ�R�G1s���0pS�������'5�	��������� ���{���߬	����ǩ�Q@f�Q��U�eY`\�M�e�i�h�)�$�����em�hi+�uh��-Q����E�VaL�YcEQYE1�m�Q[gL*h7�"�h2 �u&C�E,M%%4U݅E'��dfe����0�
���2Ƞ)��5&��f�g��͑U5��$TnYdUAE\F53T�IC[fUQk��2�j�
6֓Ee�omD�!�d�A[��!Fc�ABd�AM�F5#K�`m��@哭�DQ�afAKC��U:�uh�!��)3|5P�&M��"hhh���|0m�
iM�0���7��� ��&�r-XPOĂ@'�A ��n���웓�'wM����r�������(���n��8`��5���L*z��,�A\�V��P�J��s�"�y�������c���M0�f1f��~|n���t�"��!�1��<I�{~5ǭM�=ᕪ/u,N��s��y
��B��F�(|����u�y�4����}"��:֪Z&��S�QbYj���
�k���q�G�x�H�C�=�Ut6�9�k
3)n��ŋU�ڟx�އ��Kă�yC�߈�yC���x�a�P�fGt(7�ҽ�Z�"�`����f�Ak��/_��
Ҹ�$�[����ۛ8k0�(�����ŀx���_�q��c1<�;�5���I!�ts�S���`B#N�NF�a�Sd[���Q݈A��K�ț�r%)i�L�;�\����H�d�<߽��lRe�~��*}٬v�M�Oy˷�v�p����Xe��[�Y/t9hR�����4�h�:�&�X�FR����-ȓꏞ��-�C�C��@��}���Pƾ���v�⸅\i'([��	�T�)���/{Ϡ��W�+y|a�n�Z�ڡX5���,���3H#�y�[L1p��q�����Ds�D�׮m�R�����[��I�]�R�<h�3�f&��$3�6��H�^<j�����LlCˤ�8��s�ߟ�f졔�_�CiP�/L�������:�Y��NmSV�@�G����w�Sf�#��mP��������`Tzl�k��WK���w�r�V���K6gw�D��S'T=��MBOjpZ���ڮ�8�֦Ľ9t���r�����jr��bPm�+���e~<|���͝�7c�*����p%H^��m yz��yi����v����Bvض�gt��y�.2���DI�eқ\1c{Q��(b�z䙚���zș�־r��qX|�f�2&=�ɤ�א�y��b� ϙ�:�r�������� VF�D��wABǵ�����N�����e'�a��g��a�a��i$ל#O��*��ӻ�5�hQ�G�y",r��#b�xo2Oo��S������h��KHIq�CL�m
>><l$ ���n��w{����$��KK�L��*�6�T<���^ʐ0���vg���~8���y�E'�n�!����W�Wv��Q�/����{��x�#$f�Ѧ0b���]u|���E]�=��<B�Q�2"k��ȇ4x�${�w��8r�%e���;m�XGU�ŎB�P�O`s ��a�^b
l�{e��Z9��P�Z�:{�ύ�2D��p���B*�����e�=fH`��H:�vԔ�L�����c�R�|��K�Gƨ\�9h�w��6*�f`ɼ�����k�jPsvb�F|k�F�3���gKq�7��yR�I$a������협�S�5�;�N;J�m��]Y*2��rM��6���V�"�C'>#*2]k�1a�� �{d��t�f>4Gz��_NbXXc?B8�3mbGNՕ�W���Ze�W�7�dW���u}���Є��T=E0��h��t�~�x�����v-#C��n��B⮌jH�H��u�˻���a���"u8��f:���~���{E�(%����"��4I;���&Jx|G�
��^{HW�O�7=�p�#��[��/R���;X�C���{ C�R�n�E{rl��l�a����CbpcA�L��_*wZo�/�L�m�������GK�^:D$�H��[DYç�]Z+����E֌2��R]�i}�9�@K�n;�)Z����jbyy3�O�}��_�)�&�/v`�C��=�w��Ԧ�[�hk}-�����$����.BB2e�a�⫌���|l�J�L/c����.���7v���GjD˗	CIlT�Q�3�<�<_(��v�+��9��7��{����-���Ǭ҅Z���2�Rױ��mď*[�n��	����(bġ��?W1u��gM{��[5���񽹻�#�o�����2x��+�`�� ��{��+�ӝ�������{>��X��D�wJ��u�(�54�N��{�]z	�e��x��k��`\��Ƌ�5ٕN�^I���7�Ly�p���U���Z���m@{2S�rt�q6�>Hy���c�w����hn)�o�o/�&Bܗ�y�^
���h�k��X��^/�B��_��ܱ}Yǉt!t�HwQ[�5��9��sEռF�$O��=�Yz)�R�0sW/�Z� �����W�]�zgb�;��k��}���t�({V5�j�+B�&th֚G�u��ְR������O�{�x��4,���0�a5�|x�Bb����z�����8���c��>~4<��!��dd��a'L�=��^�b�9��K"c.�JRӓ-��#ZZv$o]c4/l�nf�����|h���uWB���uI�
Ɵ"�`)}Өf�)�OE����n��1
k�M[�dv�T��+�뺹[����^.���t�
�(�c���gmQ�7�����pﭢq���+&�Ձ��D��mB) WGmܬ���{��S��jE��|CNxT�h��4�<�sea��.gOo�Wr|5ig���lg�Z�����x=�f�������U�Һ����X�cٕ�/KܐU�*|3K�ˮ@�Toi�-�m;	Y��WSN�ɐ���w�;Y�7�n�l����H?-29YOZi�H���D�uo��3�jH�{�Kt���pխ0�Y�75��X�����[��ݿ{��q�,.ze�	�]�l�����m�c�.}��wcX�1/C�x��$+S�.b$��|����J�]��0���2OxU>ޠ<n�7��gH�҄�{�Z��֍7��̋�~����\v_V�\�^Ue༢�Fd!�o<}�}'�`�}��b��������r�R�0�B�0�r�m{����DQ�u�4+6|w��1�H��%�a���&�70�fU���wL[G�BmÔ�H���><p$2"D:r�z��t�H~w�$,K��O$/�(~��Q���{N�
����xK,�0�OxD�4��Դ�]uB�W�*�3�
k��Roh`��`��z�,���r����L�� �����Zٹ�BGR�Ur= �a*
�e�����ާR��[�"�?���8B���y�q�3P���7B�awהO�+���rj�':ؗ�i�N
����<�k�;�˭L�w��|�h�\���0}�Z�f��cމ�tN�{��V�p����z��Y�Ƽ�.�����2y�` '�"�zOf{�P��O�-M3��v�3q��9�p�J9�e)�x���L&�Zrֲ����m�£��!�玷��\K�y���obO9�6�p�Nׁ
*�O4_�7=���5��7R�x����˺yV�j̆5c^�{�w�3��W�B�ۜ�Έ�ې h-ݏ�Ġo*�����f����=����3}����p�Ek�Y���o<t�{�`��:�i� ��B��l��sn+t�\���5��'����_�ҟ�6�gE���~�v-�D�/I{se�_]�Du�ij���U�����i)�V����N��-`�E(���?9G�ս����y:���c*�Es>>�t����-���z���ιS	��^$wO�v��l��B�~�ߣ:r�j�]������M�������^����Y4�
\k�Tʞϐ6FyLI�zU�T���R�ؘ�V^ޭ{��U��5ʻ'u+��'G��M�L�,�~Ǎ{�
~�Z��E�/���^��/��IWO���נ�iž�ݼu�r�
+��_K��f�EC�Mj㰍v^d?gJW�Wn$:�w&K�|+B�]�)��C��� U�9$E�%���xc*��ri�;;>d[5�X,ݾ��)��I:�-��d�v�kzZ�;)�m�K;y"�;cg6��b�U�a��]��}"_���$�gn<�kܾ�;Xl
[�_.�nI��$�J�����}if�K~�Vz�i�@�D��JxW�,���zUБ[%k�/2�G ��[�uG�D��r�9;¸-��?D�z��6J�[PH8*o�����ɣJ+ފ����,�3B�w���;VC\#L��L��ģSaM�#�Sb�}��ï��|̝��Z���8�'6�&�����Bz�u"ya���*"��oz�V��!T��.K��b4:@y�t aK�1�W�׈k=�N��Q�du]�5�RY0=����4�|p�w<���ģӗ;q1�o�<�w�b6��G���R�[���4.C���}�n�q>���: ���8jt:j��ܮ 2�u�O�y�,W$�Ve]^�/��BWS��)$+���iށU��d
޴�m�I��t��a��яGfո�6��|�h�j��W�Vj���9iQ��ڲ4��U��wz�_f���)�������"A��!y2�w
RVp�=����3h������4{au�3�J�L��c�H��̩�T�(-�Z{�4X�7E�
��Ȫ�9��Ph��rf��ڶM�*%0���	�+ni�Y�h��Z�%��d��G�89`�̭��A�Y@��z:i�����TQ�}�        =�T�ӓ$���u��WHv҈*�Z�F�5�rG���e�l�Ò���Ec�m�gr�Ш՜�w4��-5�m�s 4�m�@�=L��תR�r�oD� $4�N&`Q�i����0��kV֞9Dm�Se�bib�wI�U-DGXİ�(T��'�F�N�(v�m��d�����E�@<�7��-�d-�e����q��D�C�\uU�q$n?cܶ}r��OB�\��eX��*Y�s��K~�9M�9�s����=�N��&���ĸ���b���%=ں���)%��y���#1�Ĭľ=�/n�P���L`3����fe(Փfpܫ"���V�yI�3�re �$�+b��%��!`uo�r�E4<�;sP\q#*|�:���*��ԄN�K��,;8��8��   4�`�YT�����4P0KLM�&��!�i��(����uӒPD]c��R��r��)i)�3�\�՛�d%�:��+,�#!�
(�A�

SRAT�Y��tJA�P��ӫ#�2F��h)�S�R��BPTMRR�� ����&�b��v�X����yȠ"]�$�*�iJ�
b6�B�FMM�HĔPD�T��Z�¡
(u�I[�4�m���8��@Jڝ����0��m0�M.t7�CT�݈�6���	��ŵq;OY6�h��f����W��P�I��ݮ��n�-�ԶmZ�F���M�ݗ��Z͝
�����9 �&f���t��
μ���e�����V�h�<ק�>̫�may�VV�^K
��>s��=}r��~M�"���F��q�Id�<e�*V�B���h��.)z�ۏ(p����:\�����(sWzOR��oz�� ��l_/ ����xZ�*?z�>��ZN���dx�e��I��$}�6�(z����4�9�c���]א��D:H_#��]eI��[�&^�����S�/"�'6�c��=aX���ٹ��k�S�ʸ�fŊ�� ��&�9�����k��m���%��}x�w���ܨ�5�5Uڞ��OY�5cw��x}�O�!����c���;\(�E���闪�}و��7f��t��t-���}��G"<ڞ��Q�H[8�z�N���^��T{�=�w�af�/��%f�e�Y�� M��K�3D����Y��(4��3���f���"K�a?FdML��VC)��ym��TR��D�� 3��07[�5�-�VM��s]ҷ�%�V�Rj9��=�B��'[o��1֓ܵ!�U�}��e�KB�m��=:��a|M˽��h�����c4�Gطu�r�/ye�6io���d�� �5&֔�*�S�d���0(5d�VK��i����1I�Ig��"~sՉ�+W���4�
���S���(���<�7d�Խ���f��CU<@��E���櫷��5ۜ�	�k��{C�m�ŗ=!���®��'��uwV�\�P1�\۵��{��RG����\�Y��g�d�bЉ��৻[
{*Y`�Wn�s���1+����J�����[�{w�mL3�>��$l��T'�̃�E�Ӭ`�?;^
M;�3&������Az*J����Ro�;ɳҋ��Q�^=����K�)��/c:׌�+NeO-��==؈��������h84�583����r�m�z+,���͜�e��S�Ѽ"$B����%aj��P��3��Ξi)LΝN�j]%�鹛6�S�fF�3�´��$�uy��1vc�#^�����Q~JU�I�D���WgdKh�J�Y=m��V��bI�M�^�'60UK9PS�6��m׷�Ҽ����=�V{�Ŕ�����)�8ϗ/I%��U��{�k�+����I���v�Y��Π"ƻ��]��<�oA���s=�Gd�y�jzټO}�����Ӟ�EzJz�����Rvq[p�)�Q�qf��B�M�f�,K#�R!���o*(Oy*p����o��l����`��R��_o1._�m0ۻ=>�������kf�g48��Q�-��&e'K
��Ҋܾu;6�]�]��ejAt�\�/��ޗ���UE"K�:T�g5$�7aD�y���x���m��z��X�&�&�y�h���y3����ϲ�7Lw�p����Ԑ���{���F�X9�蟶UL�Y��Î��β�V�o^���*���)si����Rl�[�&��]Ad[K�z��[�E�����4��v��b蔙77vҳ��
��8BgI��IVu�l���DY��{r���ڦ����s[k�n�ii�73�A���O��Q�yD
���]\�_n=��l�~�|��w�&]?|����]�j�7\���BƢw�⮵�e2�vRx�S̛Ît�e�h+����J=�`u�"�8U�0�sl��2ܭ�WLJ�G�\��x�{���|�)M���~���zN����ڱ���B#S�T�Lɭ���3��o�ňp{g�}��}u�q���t2/�á���ML�.w�9*����kצ�?^ ǽȓ�%�*W���}j��u��j�!�oENs8j��&	aCc�k����b'E3��5�Ի0���
�����T�׎#�P�5$��]GB�0SYy����ik{�z�4Xk���he'q�e��[T�lj1�}HpW����e���.�!��H�һk%Y=
�G���a�{��~7�O������T������h�#6I���Rܵ|ܘ�N���<w댴de9#ۋ�e�Ș��i��7���n�����ԝo������e�P�>|\À����uh&�^�E�Q�Z���S�kn�K�����G+Y�9v�6�g1�X��6�e�&��ˬI_V򖲰��Z�yM�1���|�Yk�M��O7�弓u\��u`^�8�t�sޕ�O���b�v�^�cymV5�åvƼ����_Ş��c�5u�fi���F�P�f�6y�;_�S�b�mf֞{%�x4I�M9��21�t����^h�u�w���/��ڼ�P<��g��k9q$!��ʞ{�}G2�0���G�����������d��_wCNL�Ѧ�:'-���C�L�q�pg�ռp��ue��#����F�{vWd�ҝ�ۏȍ�*A��G+Q�{�ߏ��sҰ�/ޙ�*y�����sCkunL��9@b��/+%�]~�F%��*vj����"��)g1�
�O{5/�Yt�Y�&6e=gT]�G(nW��<]I��eJ�o!���:������KxLr�\6Dϫp�Q���&֛����w�����u��Nlb*���=�mjTܷ{w@�Ojt���צ��v{y\_[�sڜ��w�0N�f�L�C�eV���>�=������W:-W֕+�ÍNv�۫W��L��W�]�d�̏7�Q�w��[J��k�{em�;r��C�r��M��ީ�2w���K�8�g�\*ӗ��M.n~m�c�q�1R�N��i�b�X�����rϰ�}&ȥ?#L
��௽�j������-�h?^n���z?X\T2H/�}�;��>�-�Kuմ�|��vp��轚疪�O��99�N��H��[e�?%5�y��b)�[�h����^�G�ם�ozj�o�)D�;��V�ߝ��}��
^�!���[�g�$땪c�ʙ�q�ui�7��Q��<V�n�8��}Đ~�lw�ٺI�qt*��4����mdU<[��nDdt��O'Q�:�Q��7�V�9/TY���AY�j�h���<�T�+�k|�ĥk�^�oH,��ي�zgneӡ΅�Nkm�&c�~m�U{Lٺ�}<]�(�؜��:e���<Z��+:sf}�t��Kr�Z�=S����zy\(�o�t�L���f׆��^�������	�?�Y�1 we7�hXlCN��z��3���S�l�QP�����ʫ�����׽A�����o�|���}�Vi�p�2��N����{㼃e��Yw;�P��*G�K�5-�e���]<���_G�M0E�-V�ؽ�����*+s=c�W=���Whܬ�8Z�v�l���=��)����Kj7�Z��"� ����I}:�h�CR�y��3!Rt���9R��;C����Ayը��<�W)�zZkFdu�� �!���[�ܻkr pW�:D������`	�$[�Yb����G&�-L#ۼ]����hX�M�EcN.���͡!f�5�!w3��U�ֽkv��j	���+�����ӵ�t��1�Ğn aw���N���m��*���c�E�ş��\lC��IYk=[�I���O:U|@ř\�K%u��*Ȣ:~*P���L��(m�Z��.���q����e�a�R���ʱ��!IXf��uɳskZ_g$WEu�Sx�S.�uֹT@;n�<�����˳״�����U����-`�en}�7q�m�[�(��9���Yc�o}uڥ&�*����g���O��7�$o1X�7��ۯ��g�N �       �KC6ڳ8�Ӷ�M.�����EU�rVv�Ӊ�V�Ӏ���548���[�D�]�4�#d�ErcQ�F���9�Wh���l�>�|��Q�5gk��A��������
�y~qzavmݖ%���(-�\�MO��g9>Y'h|�vLY��B���2���˘B�q��w�i���+�3fP;��&#��n�����P*v��+4���%����ȭ��4���;v��%����|B�7|9Z���)[1㼍ApL�f�؞�Jۺ��1"�HͼgKY�nԭ�p�8���-����kV=[��ޛ�}+�g1G}6�-����Y�m�6�=)�Ȭ3�M`;/>,�h��e&�H{���ru����QX$1�����-\���,F��"Nw�]^�  ��������]�ݽ/�n$��i����"��ȡ�R��H�j
R��(uk7��:�(�L�)M�rB����*�������kR�����FYoT�4�CB���"]B��ME-)����혺��H��!�񬨁7���%	@�P�1CI��%4T�c�2 ��Z� O��w���8s�\���+,��d�R�ls15�+X)���NH���5��\v��3�?6g�L��w�SM��Z��M������]lWo��M�h�z�T���t���h�Z�9\��=���*`�������%]@�G�
�%�L��f�9���yZ�n�oe��f�%�Ú�U����5x�z�p-j�s?[�����k�����(b��O9]�؏�����T*1�j\�˺��$�*�>-�މG�	�n��Lӽ�p'�) ��eo1S��?q9���o9F�Y�"�3>F���Ou{
����T\���ܺ�챋P�{�+6N��?0�~l�%KG\ܰ�Tn�.���Rޏ��7i#�S�/e��8�X7����)T7YNB��a���6_L��r&�"T�N�*4f�)u	�5��7��[�<�ܥ%{f�yx��g͊"�c��D��v�h�=�:�O��(�/{p�v~�-hc=o4��j�[�zU��?x�A7�YV���2����j9�A�硫�'	U��@��7lF�ݹM/1@g����cy��[��&ɍ$��m�Qܡ��fzg�TEI���Y<X��uS��o��"�:��!nLL��eb�ۜw�u��kL�y8���n�ئ�]s6n.��קM��sҶ<��K	]�k�V�k�9EG�]��t�p�zBt+�O=Lͷ��xXk{M^֚K�r��b����±���}:�v^f����}�J6��Q�(nъ��u(!3+4ڝI#�L7��������F0A�=oI��2"L��H�.�sVٱ�K9pS��Mj{R^���q��0�{��-?h��J��&H��N��s��
��Ϸw��xH��8��k��x7�'�����6��Z�]��w�W9��&�ܾ�g5d��B�W�m6����^�j3�,.7��4�V�ni��������H���7��`��[ى�|׽%׵�Y�j�}�W�N)��!WC�m���U��G��[^Pz
z^�{G��^G\���{ΞA֞��k�w����nݰM!���9��g�1����#�-�+�&h2�R�)\��aV�f�骺s�L�"�����˞��W�����fn}=��_�Ξ�ާo;D�����
o���^��֌�Ύ?Q^<U�A�u���S�yɫ}J:F�_�;�{_d}-TH���\𳝶�;���}0����S)a�U�ک����ɝ�V�����v���'���[yyw��/>+0��<������zΦ��s����;�q��Y�fq�+�.(�\�^��EO(��"�}��U�]c��a��X���8q5��f�diޛ�Yάkq�8�Y��Fӂmޥ��4����-f�	IYW��<��j�!���=�t\ n+�9��|�2��f�y���{_t*.�Nu��dU���o���Z���u��'j��;���N���D�봆�w��S;�6�/������oԝ���tǓ�>�젹�~���{�~x�o��{j9R{��k�U輑�̇w�\�������u[�1��=��h�����OSk,W��%]�����=2���_�˞��o'�BP�v��R�q��i�]��&��܂�%l�5�s�^\��fSy��ؽ	s�ow����P��٬�������v��m.MƬTý5��爢|�υxĳ�{O�wz��º-KqT�-����J��h�w�k~$;J�=�B@�dn���2�}2]]��N����b���A��2JB�:8ʽ�X����yH�bv��؍-[a��Ug5	Dy$f�ިnʝg�R���m%:�tms���n�IЬ�IOi�E������=����>��y�n��ښ~Κv���K����=$>��k{��z�\����S�^؁�_�D<��[�˘�|׵��o.�J0什W�|���Z�B���'�=ԊѸj��v��){�g���y����ŭVz߃�K�>�^~��V���!����_^c���WC��H{�L����|A�nsk�y�W����W)�Mg�
�U�^���0˕��5xx�i=�����.��F���.uCխb*�K�HW��]��ݪIn<6S@ԛ�%ҥ��-_oY,_K���NqIhN�MR&\l���^�U�mo�2�W��֮�L��BSY�3��^�~���UC�����9����ǘ�ըCrʍ����0�|��?%�PZ�e�R*��rz���R�ai���jVy�@%�J~�z	�x��3+YϢ��H�},Ԫ�hl��}=��|¯%t
�ٷ�T��uV��6N�$jLGT��O�%D��Չgf�ʢj�-	�\}l����Jma��X��;p�a>�z�uLO����RfЀ�0��E�2�x�j{Պw���.�fg5yE�e�uόrP�`��L�\�ai����5���tލ+�����}��*�Y�
��a�)��v4���֝c6�)Y��+yo�7Q�o�ܶ`�H��$]��r&T/�ˏ��	ڪkޫP�G�!�]�5�on)�S/��̡p�#U��o��hğ�G�j������u���3�>�륞��n����+j
�M_9�*�rhy0�ϑ��l��황��.���w��P���zg)�i��y�;P����3Ґ�"7&5`��>ᴫ4R�?b�j&4�R���ᾃ[�=��mB�4��,�՗~��0��6瞬��g}��g��tJL�=�)����a�����z,�nuM�ϭ�V���^L�wS��P�j��E�*ږ�)|���H%�t9�o��C�e\�����t4k��[�Vm�p�����S5e�{�3L��>�����ۈ"ˬm��g�p�֛e��=*�Ԫ{ڒ��94-�=h�$�^Sכ^��45�]n�K7�zN3N����R�X���"� ��O��[{����Y�PD�9��'�.��EY�
��V׶���,��lS͎�_q�tڞ��Y��X��pC��բ�ɞ^���� W�_*+d��˾���I�9M�4/�9�6�? ����lTZk�y�������O�5�=lS�&��mdr�Á\"�2�rIv���G=����������_;Z��T4�|+EÖ��-f��	A���A�_�y���-t'�]po-l��M�7$T4����Y"Y��XǡFo���!!�7:3�*hhog<X��kB������l��t^�k)�ӫ�?f�G#�ZE����	sLn����nOU˨k٨Tn��]f����4L�J辞"��V�ou��ͱn�LrŚ�گ
:�&�Z%6�vS[�*SU�%�p���yq>��G� &��	0�ߟ�3����ֆ�6��2W��l���wP�0O��0>d�<��t�ھd.�ژz!�[��I�b��O*�z���}]�2���̯z�r�������\��k���~@���^dSUM?�, D5a��P ���10{U=�?�$O�&�Z8Ӯs��M�3���6?�a߃o�;�"(���b�(@��P� �����94����o��|,q	�')�A����9|�C��1s���J����C_+��������?�������<�a����>��4�`������?��p��ӯ�GA�~�r��� �h=�7w��9�AP��<�g��k�}�� X^@>�DAC��^UQ�!��Rb��������������ˀh��s���u���}����>���a�~�PAC��u?�?�A��C��h9�JhT������?��C�MĻ��75
g�v�3?\+�O�~P~?0�Ns���:��G:?��b� �F�>0�޳F��m��� ��~�I�[*��B�8���>9������rl'������c���ڪ(}�<�T�}g!�!���}&� ~��?�	�f�o����w�?��[�SG��p��������?O�?=\� ��p�}�8��(o��,�i�?�O�����B}��G����0������09�_y�����>��>������G@ ����?0�������?PAC��%�����`����>7��p�4Dh��>ބ�s�䀨(A֪(x��;s�@�65�}F�۳���az�:7L>F���-*�
 }:�) ��4辜�:�\�*
��b�<�
}G�.�m�vy��q����8J�Ï�BC�'o o��Ӡ���`��AC�A�ϰ�O�z)���*�
�~��/�B���?@�a���������|	��R�>����S��a�/����4_3��z{��'�O�#��>�6���:M����A�����I�`~�3?��:K�*�
��p���G��C��|����~_����~`:>B~��ςs�r�:H��h_v�|��?��~�ψ8O�O?3�_e|~��I��x3�߀|�U5���}bp�}�������g����y#��������>9�xϫ�q6@��#����}00" ���eGO�����;�O����7��}�0DAC�_����;�p�w݃�o�p/L�����٭np��)� O�#��
~^�>��_���"�(Hn�U� 