BZh91AY&SYme���_�py����߰����aU~xL   �(         /`   ���   � rtPIv�H��l�Ph �]su�
 :  �f{�{� �@&�4h� ��  P   	@     a�   �l�����{F�7y��.�{�mzd��yݛθ��{޻+nJ�� ��������ݍ���]��{�Ӿ�۟{}�����|�_]o��2>�}�S�{�|�ݻ�v����f{�����h���T��: �}������� �ݾl�ӞǠ:]�J�{d��������z��[QM�vAw��x�mXm���w�)}�{�Pw}� k�:;�<����\Zwuڷg�-����䞦�i�wu�ɺ�� S������  B��;n�ݸ�ۥ�g\���9;�ɹ�l���mݙ��f��Kx(��:@��=ݗs:��p��k�K�۝:gg �wQm�w�{�m�6\wS������@!�� �\j��wr�{��W��)������ճ:[wuu.{��^���n����Bq�����nۨ�7@;]�mї6$n����k{)�6d۳�n��$op  .f�e�a�fQ�KHá��\�Yjl���9��ԜoB�B�Fn��6�i�x��s5��kiܷJv/y������gtUݹ$                  *	H%	QP�            !*zA��R��C�2hш  �214�J���	�� A��JmD&R�H��h4� �4�0*j�"m(О��=@4ЌM2hCA�&� &�D�hL�z�m!�2�d �jR�Q��&L@0 	������W�(�F������LUir��a������(�Y� ��PA ҡ��6�˙�����q��|;�m�>���g;u�>��}u���{���~8�垣�m��jJcvM��6���1��9�ʾ=�wcm��coV����$�*���$�GpO�����v蟏����~��Ӄy7���O���t�}+
���xK�����u����t��'S��-.�I�od8U	&����eɯ�'�bG���͖�=8M���I;��͛8�S��V�BUnK��N�{ ���Ţoy%�6#"o��"c�l�����'Q+�I��aZ�S|�4�S�:��ڮ�%���ådJ#��s��"'[��"{����J�� �ܤK��-����Jӫetٷ����':DN��-�N��+H�J6�&DGޕ�t���r�DF�V�]J��y)�%"/%x�\���H��U�2�cy+��J#��ʈ��J��jj"S�H�ur���nV�=��7{��8�R'Rx��Z�<����"{Vl�S��V�,��Ҏ:��w*�ǒ���SY��"m�O:���Xtw�ZtܤM��tN>���<�RYͲ�Z�JD�r�=��6c��z��ӑ,�l޼��d���'��^�ʡ�-J\��;�-�n������FӺ����:%���Νg�ɱ��r#S���jY�t���MXx�� ���74�j��m��k5`�t���"�1��|���X{&�Zo��&�D}<�Dug���O}(Cy*��U�"X�U%�I,� �βN뺑�;"9�*�ʫ%�ġ�K�T�C;��:�� 9!�#��]�����J�R�q.�����	�'`��\ ��sr�d��1��w��u�=��F;����Z��E��k�]�s�G;�s���G�q���ۋ�G9���}�w��wؿI����w3��.��۝��M��R�KrR��W�=[�RC�����ʳ�꽓�U��~j��=����7D�"vc;+]���F�����&2��34gqL�9&�K�'����M��R&�'��0sW��J�
�Ğ��LOt�="u�=�-�*�Q�	�:��#�WI��ٸn$H��KLĖ>)�7�x'(��<�e����d&��ݤ�tMўH��K��Ii���<�{]�!g4��D�=�����I�;�ɿ���'4�OYmɉ��$�{$�7�;�O2LH[$��2{b{l���2{	�����I��h��5�$.�=�&ĩ�5㳒k{��8���-����F�I�N���e�^�,JL�	+�I����&$3I�LN	�d���y ��4�%�䎓�V�I��f�I|�)��|�0�:QzO2D��nD���ɪ`��'M�8��ON�8�,oġ;�0�	��(M�*�"]�-�(IH�ĉ��'D�bD��p�FB"M���	H�-0I,�����ҍĈ��DE<P��u9{��!,H�K�c�DÅu"'���hBx9I=�H�����x�<�<t���3	�a[H�^H�JO+[NN��xt���DK�D���I!�:"]��Q�pH�ĚL�:l���<$DL':0H�Sd��&y'��=��&�������'y'���.B:�l��R';dM���&����(NA1�(�(��I��'���
a��'��L=e��!f�A�gdIB>��.�{"xC��<U��c�,�zz��s�r�ja�p�d.�<����r��Ʀܳܝ
;'Pr$+�׎��P�#����������i������ ���ׄn'��cɫ:�N��F�T�ٮ�é��i��]i�Wv��^J���W�]�ٚ�ʐD}ڈ啘#�IEX�&̢�&�K�����Գ,�S_��N��6Ϗ�ʟzV%����S��þjxߥ�楒�sH�&��tk�xG�Q5}��dJ$jvvt��ٹ��^���˒��#s�4�7�����DX�7�=�A��x�!�ꈋ,�jʨ���H'e��;����R�J�<;jY�H���㜈����*"Wbxۺ�`�"8H�)�FUDF�Q�R��jp���id'jX�2�x�54�$�c�DGĈ�I�J�-�I^�DE����	�55�M'���B3��DNm�D+���G{����#2�'����o&��Tã��Do�8[;��p�擃��D[��qjP�=槈=�OwR�gj";ʈ��P(�&��"�J�Q�jt��t�&ɳgMȏgM7���D�D�%%�������ɧC��9D6�Sgh�>�F�G6�@��K���D�e	����G��">��mIc�gE��{��<>�T&�j`�����F��^�x��W���΅zj		p7C���D�G&l��!�,�!5���i��f��5��j=�n�F��Q2�TQ�8\�<;�:#���JL=Ƨ��k�K=iI�*tN�S�5f��D��ji��s[E�m�A����n�Zއ\��;��F朚Y��ߦ����ʨ�un�{���<�����'9/���P�>��aWb͘N�a�<nG|+�>�J���n�/�Vv�d���G������Q��ܿ5!q��jz�F�cQyQe�������t�ٚ�릎:?t^ϗ���8];�KW�5j�{5}��=#rG=R��{S]�Of�K��jvn�����a��NI��`�=�K�Լ�؇rz�S�Q���{.���:]5:^�F�jk���J�S�*��K�ԫ�W'c��J�z���=��ި�p��:w��S��7=����.xrk�ɕQ�%Wd�jT��w�OwQ�ߪ>�R�Ժ�z��^�er�rU�A�B�9ʘHHY zNɺ�Tyʏ7Sc7Q��ȳ�S�ʮNS�#TS����ܮ�8^���$DrI��G��+��u����9����Q��i/#�(߷)�Do%i�Ԯ	���<�R"�W��ȉ���eY�2DNxfJ�a҉�DN;���Jjk4ԤM����Qw+��+N����_%lN>��Ŕ�9�V�O%"Q��"^2�غ�twr��etٷQ��"wuSJ�c�M:������<�".�a�w�ZtܤM��tN>��Ŕ�9�V����Rp��H��U�1�ç�74�OS+d׵�'Jd�ײ	�^�g�TsH�*ܕ�;��l�u,��8<�9�}�ܪOɘ�a×�^;'�����O1,�6oV$7��pA*��5��uMV�Y��bt�r�f�+���N�x{��.v���O'�9z��tju���c�XX��I��D�ʪL��[ ��A�Ӳ"W�ȎD�x�S,��gnlw���7UI�n#�-�t��$=�rCzoR�r��Y��ri.��ֹ�9�8'���dVJ}9�O��n8=�o��wQ���o]���\��ŽE��Q{�ٮ�9ߣ��9ڟ7{�^ܪw+{{+�e7<ܤ�z�Ta�r;�&n_e�r9;s�rMɒz���=
;�{���p��L_��;r�wpN��jYێN�';�p�䁽\�v/�g9�q|��9�o�g!�F���$�ΚN6�o��Ȣ��a��G�����
r}r��䣓�dg����b�_Y�~�)a҄�Đ�J�Z��G(�Q;;?�ޜ}Uuh�E�����z�{���[�SZ��˒O���㹿�����榾򶾧=Y�b$ݝ�'W���V�]�&��-����#�Ӻ"UU���bAϷ�ߋ��yq3�Ս5V�[��5.f��5���KvWɕeIg��3|4��I����q��.l����'�}Mt�U��9����N&Ƹ<6�.�[�}O��{�\��MZC�QD��_�i>��.ޫF�<��+R��.��{s�>Y��j���On�鋘�>�O����*M����Z���ؗ9�w��kDU��q�=���j�WSM���qD#��;g�%��uz~Z}���9�����?�٤S��{&���,�rl�ww��YV|��S�.���?�߹�W�+^R^&����N�v�r׳�WV(<\��S�Εƻ}����{�����O�SvdY�y�j����i}{S��{��s:���O����>g��E��Þ�N}�nq		)ĥ�����Č�/�����U��&s����N�~]�Ν����Oo���=�l�ss!�ϻ���[��8n�ʾ�7��*����Nr���vyx�vX�,����ϑ�o�_gf�;>��;�
����7x��</9*�{���z,�3ʨ�k��-O�b��R��6l��}G�<"������h��n�s���?��Z��9�4�xE����+��Ν[��#�f��G���A��r����ܓ;ř��7��%�ywy�|����)��ּ�7�w��W''V}э_ͯ�͟/-Z�������v5SW���Ij��IU�4�VT�Z����j�:y暆�k��cIj���3�uq�}��y=^�1,�Ȫ�ժ���w��l5	|���\Mjj�z�g[;V����%W�ċ2$��˲F\��g:��g3�%�"��8M5%3�M��T䑟Mrk[.��c��vs�*|QuURQT��%
��U���K�-ӮdYWUj��(��
,�.���:�*���|�8�|�k�gËʣ=�v��b�"%d�2�8�5����m⼜Y՟_�Q<�|}��91��1�y���g<̽CX�^�sX#����g��K
�x)�Σr-YQ��W��<�ƚ7���<�b�3Q�Oc�p*����.�(h/�qz9F�n�)Ф̫�>���g����װ��5�V�!y���Y��8�9
�5�7\-1d�����{Y�BE�x��;�r��2�!� �4X#h�ĉ���̫�fr��Q�|F�L8`b��I���ˆ���4�˞݅�2�>�C��o"jw8���pY���e�(��_���ˣ��3�[�� =8��%�u�L�g8�7�����063��9ÏK�?���P���p�Ӄ��/vB����*D}�z��I0�ά/P��{�#���-e���B��/N�_�E�2��҃���L<��3�xaSQ����x��:��>��F��Bg0�
��+G�nv��{B/OŔ5�XUP�<�~9�̋<�����Y�y�,�1|�%g-&�|93�f��JQƞ𻹜X�]e���5ydDl�c�Y���F+��qm�>YՍ��B�ĳ�֑�7�ݵ�u��ѩ�0�Z��9��A�^�2�M���L>Q�Ǵ�^5��X�=�s�5dY�y��_-�>X��Y��5D?��:&��o���T���nT��fY�>�\\�*����W+���GS�5��o��"k=wH�i=�\��g�C�	�_��]��֝�jϦ�*����ʖ����<����(��� �g�G�ʢ�tg���+�bZ���|X���r#��D�h_8��\;�垻�L���:|�Z��}3�7�L�=�i�o�^�۰���z��ʲxmX�>���߅�~�{��9*ϓ�Y]rēC��y���$�Z�_:����oQ��󇷮�ŋV|��oë{�(��˞��;7��{�K�(��A�"|����A���ܵg=�?�C�?z�^�C�{*?�s7_�:h7)�'����؅�~:�ܣuA����l/���3ۺ�쯻�}ՕΉ�7c���{z�op~x�yyg[��)����j_,���S�x��j� ���dXZ������)|�E�s��,~X��9�v��Z�P�kG}uf����z�����^��V|���E�	�u�ש)���ȢĽ���Y���]��}Ƴ�;������j�.1�qcIc_x|W=����jFG��C���];�v9��X�:����NG7�3�{��_v_b����K����\B�՞IcUf�������.2H��f{Z���ˎg#&㉈p�v��õ�ᒣ���j<���#���Kdu1��8�y�����úh�u72S���ԩ+,u��擬x���y��s�:��G���"ȍzL�(�&����?#����=�1�\�nR�*�:��RW�E��G�q�q`�r���cY�hǫ�/t�a{7��U=�:1q˘�#��v��Օy��4�^y��>,�Ʋ �3$������dj7E\vǱ��ӄK-(�׍eG՞���3z�}����=�*/^��-g���4o�z��MY��<ĳ/6o,C��x���ő`�q`E�c�Ƕ瑾C�Ks����/��5��3�{^$s�:��u3��if�,/.Nd��mx�$myA��k5��o�qdGc<,�A|Ǩ;ߋ���tNmWҲVC8����7�=��X�.q��G&>,���r��!�'�,3�d{GP�MB�M@���n9��}����^|���wnDf���b՛��7�4�si���k.��*�zgt����=3���O1��sԑ�FN,9�#f?"n㙰�랣GxN=����ĳ�Qx�Ώ�mE�XM�H��f�nv��w�y��L�Ǉ�b��a�y�PWI�q��%���7�|X���o�~f�:νe�e�y���F��!��?��o!sVy�<��g>y+ϖDFͬ��[���My����qG��!.<��]��C\�E�Z_�{���p��>o�udDo:�4�X�ߘ�gdFDj-x��;�{+OL�4�׳����aLԇ{GE��<� �|N����>�t�ӝy���Kh��2�
��A�o��y������g��/�=YYQe/۞G7Ṛ����՜@������"Y��X�u�"_"��cF�;Y�<��g�YŚ���|�Ip�ğ���>K�=}����![�Y�l�ǟ7����{��{49=��~]ݗ�{�qug�L����wܽÍh9��/�}�^뽗�5�O��q!���<�T��Tg�s���)��|�k��:����V �T���f�F�_���9�~\��>γ��7vV䬜G�qS���Ps�xZq���4��qbX�\t��$�x�䗋��꫻�pU�����p~���+�����QH߻
����;���9�v���C�g!um��WJ��%W]�^�q�Iw�x��}�C����nW�)����nr�Ob�,,k�N���g��}��Ȧ�%x��t�^��~��s���s����H}>�o�������|!�ɼ�:��/:����;,�;�7�&�7�����/+/$�M�Ջ�zy(���ս7U�gW������޻��]�}}���$]����v���@�lNe�Y������s~���l��?i�|�M����.��J���+�{vs�g!Nw���W��+w��l�g����g�;�yo#V� �����s{�WZ���z�D�޵�Mr5�2v�ߺ�ݜs����g~�Nw��{:.��;���F�N���竾���.�׏�;[��|���=��|����~�,����z�j����~�}�Q!�ѷ����x�n�?_��Ϸ_�N,�-N:7��Rɻ]������]�y�^/9�r��z��s�޾{�����3w�y���{�{m˦�����,���a	���t�U���v~57�J�_RGL"R�J�I9��V�ҕ&45[O��U�"I(����z���uQʢC�+]��	�/����䭊�]��YY���T�����ĺ���ȝ."��q*�ܮ�͑L"�Ucʸ���z�K[j'�K$Xe�<�NiJ����)��Z��%NB;m�I2�ڗ�U2�%\���KFE�b_��;��D:�"ʏ��X��b+uZ�&)v�b�bMd���=�1�DE�RBCZ�%���-X:�v�H*�����*����w"�Ōd�n�'o���	I��"1!�ߡ1
�"�"6�]{fђ�Y{�зr1*�7r�"��ƪ��TPR<�:�r�6�ƭ��U	�,��Q	eI4�.����񥪢��BI4�im�)i�9�
��x�%��`Tst%CmFu���I
�l�%G�S^���j��ēn2G����r;�ԩɑ�bK�U�*1'�����%UHJ��yLw%��?�ת�	R�ҙ��7ks$�H���Th�jS-�N����]�*��"n��_�R�H�ly�*�$��h�s4��Mʔ1�&ͩ�5�iU��E|a"|�בl�	;nD$2��\XԘ�j����ui[�K��yݐ`���f9]����%m��]%��-��"B�kM��V�ڮ"VLv�T6�!qbb��)��qʭe)-�Kbs	�^p�I�1�1+i-t��B%cX�P�v6�O ����$�!��
.UU�����]�v!%�0\�)���7]��b*Mn˂���u�;y.W:�C2m�Y#%a��Z!s�eAΌ���p�ǫ����s07K�u�0�W�Ja��+��<�ê��w�H�ء���\Qy�7)W4�� ��\����U���S�qM��j!b%]'`�$Gp�tFT�E�5�`u[�<��f�C���q���D�*�I�{\�����H	&�딕�T�*��w�MA�Y9Eq1D3�pC0D3 77$S�y�.�]�ֹp�s�O�������4Vk� DI~�d���@?E?��~srJ���W�GI��O����_�����G�3@k��ATT�5�S�_������;U_*�U|��U��W��U_<iW��*��*��*���UW���UmiU_+�W��Uv����U\EUUEUW���ګ�W�UqUmiU�Ջ�oj�U��*�|��W��Ux��U��Z7��iKi�dM�b�MV�VD
��:�lP�M,�(�bY�V�f�L�7-��r�:��(��گW��U^��U_+�U|��W��Uڪ�Wj��iX�kU\X���UqUUU\b��Wj��^*�U|�*�o�^*��UUb��W��U_,UUX���ڴ�u�v��kJ�����1TU��U|�՚
4h�Z4D֩��VC�5mF��m5f��KX���dc$	HIA{����j���UW���UUU\b��W���^*�Uz��U��W��ڪ�ZUV�*��*���U[ZUW��Uz��]����UmU�k\Uz��]���UU�*�{ڨ������UqUUU\b�Z�։	jZ�BkC����)BZ�Q�g�k_���z����gʪ�*��.�W��U\X������UmiUV֕U�UW��Uz��U���W�UqUUU\b���*��v��U괪�����U^��V�U�U���U�UmWj��]����Umb��,]��F�T�,)���un�ܜ����Y�թ�s�:��MLnFȂ�dE��TP*"��*	Sl�l��(�q�
mM[;M���;C�v��ը�������~v��6��������7_g�y�����O�~�������?i��?y�K!��gH""'�Dĝ �"P��,D��g��< �Abl��M���'��%�`�X��`�%��"&xN�(L"p����YH%&�O	���dN��8'8'l�"'DDL�"t� ��<"`�"a�0�0�ӂp�Bl�6A�&�A0d�@�BpH'��Yg�,Dĝ �"P��,D���6AAA:@�H>�0�o��j���,+8mn$X���Q���dB�,F;G�JU H�X�Q�
���WRHIU�FT<�$tX���B��bn��e+���U5��U
V� �ɖ��q��\r2�g�22ɴB����ZYk���X�U�!ē�ev(�B��UdIDZ�R�����Z�)JJ�+cP��BX�[V\���Ȥuq���p��e�?�-�c�8��*$��b�D�d*��B�2��CPR�jQ�1�Qb+�Ɔ���׎$�(m��A�P�JAAe�$7pE�i�!In��hbeD�b��2,���qL�cʋq������"	T�K$���D(�pY
��%��&F�U�&�lB#v�et�II���>|�N��U�U�Qx�R������-�Mdt�����
K��D���Z��vc#u���܈�����ej��Q��1G#�24�#!�\�eRJ*���&(8��JFe�ㄦ�ȮBۈcvy�<��Y�52�c@�A$w�TPD�%�4H�Ae�(XX���v�K�!!�eC�ɒ�c$J$�42��J�� Q4(�H-� K��IR�E�Ke(��,�Y��
�Fێ[�X(8XWT,��Tt#�A�d��R�(�F�y$�Q�&Q̑F�KJAb�2��nbC))H,�BE-!!j�.!*�h��HA�L�e�F��"�,xD8��XVD9�x�GYb�������P���!Y%&VV&V4�HVeeV��V���E#��)qe���v�h��`�1dcRcTT��C&E�;I1܊<�I�`�)�Dʁb��l�	��Q��u!�T��pX��:1,i���6De)1*�Ʈ<qa\R$��Q�QL$�d
�t� ��Ȉ��,��+FKfD8&Ҋ�A�7�"�:-��)���22��T9�"���rBH�E,�T�+�>�l3q6;F�K�-���<�"�т�+pb�ETE��ZR�b"e��ǍdEy ��E�UFJB�F4���%�d,.4\M�И$=!�j�H�+R%BbE���R�U`� �-E�B�����D"��a��R�+!�F�.�,�لaJ]�FIi�E��*b$)2	�@�2��(A���9<E,(8$�%��SlB��ī�lLt�!L��!+R��D�����6����X�1 �IErBQ�Q���U�������Q���*,X2�)2X�ʞ(���G/,�2���IWdmmW��a"�����)G��!2�n[e(��BD��d�40E��[6QJɕ��b���1��A��AJ�hB
�U�R�DŔ�DmT!�2�r�(�DQ���Ul�c§u�������Y���3�q�I!�JZI[��m̵<�K��b�:��8Z���9S�6܅n��r����r�STn��۪H�`�X��NX)eV�X�w�GU�%�2Vӵ�Ej��:D�Q)QK��VݒWJc��MKkU�IK]M�HI�v��B�',���Z�U�*�"�"Gc�J7]����pV�)1ى�QS������!��c��R�ڔ�`��VEb*��(��T�Z�V̌�1(Z� �TQ(��,�6�"�K����Q)ll�lUJ�Ǖ"d����T�MHݔN	�DY$�Y�iui]q�cN�[VRJ�n9ehV�]J6��+Tsu1��J��r�$D;+U��L�r16ة�:�R��$��%&F�n�ԡ\�HI��UGI�%�b��J1&۩��M�����Q�q�J�� �eJb�ۺݚ�%J�*��e���r��傕�*�\�s*�--�e�"�vZ��\V�,J�\J\�㩥c���e(��pU�BU
6*�i�kJF�lUG���Q4��V�4��nY%�9!%���D������1�OZj% ���G�m�H���Z�J:�T��VG\C��j�n1�%�V+��4Z��J�-�r���F�����X�#�%�(�LU�75;[�F'\��9
R
��,ld�j�Ei��J9%Mq:k[ �e��5 �G#��H��+�-q��HV�%-�n��R�V5i)�j(�\ȮY&4���Ƭ�V7Ui�8$"+�ǒ�b�G���o���|����Uy�s�}�kF�j*��������s�s�kZ���(�������Ѡ�U�UUQU�9�9�ִ�P||C��kem-o6��:�N�Ï:�8�"���=���������e�[�&6�^[��[ĭr:�R�A(A��	�����\��EZ���b�*GR�$�)lU�Eb�P�dꄲIP���j,�8䖕�8�����H�V�Y��ʊ�5i
&�B�1�QE�����a�m�9,���ʫ4�LD �	�GUŔ�	��J�����
�H�R$)I���(�R�h�1!U�YnLub#�-("J,�V�LLC)Q#.B*�[J�.1�Eu)D�h=�����LIc� ��D!YJ�Q�h!�dhz[��!���V�N��)b�Wi6mOu�I$���Gc���GiŖH%��umIB����	���UM��%�%KZ��bI)Y"#�R�Gl)!2*Il��6�2�!5*���EKT��mj�I+ ���ڊ*��ZZ앺��|����KZ���.=�ԫ��$��c���ȶ�y���xu����:�1��8x������:s�s�;���*��!:x����l6��;V���N���;69
r{{�}˫τ������V���=�9��i�j'6��΍�I?߄�UBæ����a���H����`d��+�G�&,���,�ףn2���Gq!������4g2FX�E�L骪ᓭ�	7�~l)t��Ԕ���]eY��Ee��VQUdv���e����U[���ρ��d<f��At��Ԇ�!��f�~��D�8`�t���8C������׭j9D�x5$�Hq��Ш=4�Z�_��@��G��:��yQ:;-��D3 u8h4�$������&3A��iГ#�w뫱6C��#n��n��e��a���-ݪ�dD��IHUm�AZߒ\3�������1'���A"�_t�C$;�8!�����h��2�>e�\iky�0L:$,L0��6x;tj��".6fTUkȱ�����I$|�t�#QI���	����d�Ӈ>��z�	�Vϸ��1��a�97ǡ�2���C�r���F|w��%%(�x�u�i���Jn�32e�Ao\6j00��LCG:�8tx��F�#�����o}sr_]�S��8`�y�9�%[������V�Z�q���<�6�-�Æ	�0L:$,L0��6s7�R��$�]Ʀ��$��>f�ŗ1��f�g�{(��u*b�t���AdҷZX���Y'ϣ#����L�{	}h�&�qV�Ql���#9��_��ԩ�#�)Hއv8rS^>$�Ql�V���ܝ�0>:m++⠕��&���+ԉ�H$�U������.�a�.2�N�����&	�0�x�3����Z�+ώň]7P��Ս:�]&w��]u�ÈE��ɪ4����X��q>��mNҕ���w��9�II!w�!�;���]�w}o�����m��w��}���vr�{��k���f�[�{4�|�v���#�V�����e��͛�(�};��?������}V�Oo9��}��x��ta�����<�''ާ^�)��rx�>�����b �9+ej&a\?}�C���r��	4BqN�$��`
�e��d�~��Ѳ��Y����7��i-�*鏦х֘6��4�p��%�HZ$!$���@����W���+��m�,�!�x�vy���I+G9��m=�W�F}�M�#���HM�4�HA�v:�C�^�0#�p�p�0���8�ۺ4�����C�:xO��`�,�a�,�p����e��?������>�$�G�s�:�4�A0��^��hh�\8}�ǈ�͆I%96���3N�̏� _�'d	�x4w��1UM�'�p�i����g����ĐYE\����y���$N5l�;�<C�ֻ�v�n��HB�b��g�9��6[C��Q8jT컗,�큼��h꼭�e�u�^e��y��D�0OA0�xލ�MԪ��>t��n��H0��.lԒI<�_4���411P�g�*>�f�3(�wT)$�ס
����49��kD�H��2N8��"T���8��y�Q���X��Y����؈&����J�qbX=oT��M�m�l�,���nA�ϣ
)�D�T3��d�s�+��G��	h��)"+�BC�epK��IO���Qke�+iխ��yםx��>>!�e���gYf26�t�+C�I$�pV��x����eǦsD�C����Ƌ��Ɖ!U��!=��z�V��Ӽ)¹�����՚6�q>ڔ:4l��~�m�3��xb�M�Le�e?fiLF���=F���U+��Iթ��d9M��1d8pJ�*�q7e2.�2p3$fG�\�6���!��6Y�����&	��&B������ވ|�M�h5e�(R�:͂�Ʌ����Lќ8n�{i�[!Mc!��b�"!�ֺ(��:��AS�=n̊7SQ۽\����$�&\�8����[�{����|��{j�_��r��{s0y�g%����E�;̘s�>ʼR��F����M��!��e ���.k��N)Zo�6C���jJ��H�i��M��>�|�����	Ù�}y75�EC+�WHV��I1�e_*<u�}�$ڭի;����ɢ��\�'CY$��ì�(J��׏W�o��Y�e)�g��68���B��E��#�c���M�Ù�Z���ܦݐ�$'ż�fܓ>%�,*pv���>Չ����tܣ�M�Jb<���Fl�gŝik[o<�:�n#κ�6��k�^�p�+Sk[�$�,?,�oߝ��j�:+�'kǫ�=R��ֈ�FE�V}X�U}I�� �X�Sx�9��:e!&1Fg�Dn��2�L���>zA<G�k-�iI��$;���=��$�[��g��W�^4G�ϲ��K�!���$�
ɟ�n60!F�,�r�'�!���<���b�'��l	����$�	?g�����<y�<_��t��Y-"ش�X��[[�^$��Z-��$���y6���F�*-"�$B�"��؉rTZU�	�-4�i�Ki��	h�ثF�1V�KG�u-E��y�m1V�N�����i䴴���u8���-6�,���m�KKKO%��ҭ�-[�i�KE��ٴ�i�-�[�r[KJ�i3'����d���̘�ylZ[�ZZZض��Y-�2�Y���Z�<ť��k�ܞǎ\���<m�0�I��[8�����0�h�[����+��Ia���ZU�Ii��l0�q"ثO6é�똝u�KO-���lE�il���[[�^$Zy--��$mlm$g؋��q�'�T���ǪKִ�!�l�,��E8P�q�*��O��s99G�i�5����}(W�'8����M_z��/�6������_{���s~���\sm��+f�}�z�l�/��w;Ӈ��Bk�]�s#��y��݄���w�i���z�����3��t�ۚ����5b����M�9Xq���џ#�s��s��������j�/j���>�jӽ�ޞ�~���H����}�w�ш˾s�;_k��֝������п̻�����ø=ݕ��]~�W_��~9����������}��ѭo333�b��"������hֲ�33>�*��*�{��@љ��fg�g�O�U�U����uu�Yu�V��y強�많�!��U�n�QQZ�EA�~�����۩��Hh�Gw\��!�<�<����a��*W{!&���B���)�J����?#�fh��I���dH@���x492@|�$��p0A6X��dhL�BQ�L�tٍsS[�$��zegu,�G��s3���J4�)��z����}⪪��YCc�!C��d�d������aDE.����7��Met�;�
�}�I�&$�b�n��`큑ܠ,!���vV.��� e���i�	������\��6!P6m��Y~i��m�뎸��Z��x��ꍩE�Pv��.r1�*+BB�IH��e@4| :&��Ú!@���!�ʐj� ll���YC1�d�����?
�	L�"��zn�j�nz�8C���
Zb'�g[�)l�ԃ�(d�<V%�g:�wV�V�!"^�4���5l���dV11���zC�	��_J3R]��A� a~��T��c�I�JR�JBe���x�?���1�R���d�(-���GĒB�rВ��%"b�����> j�*HB	^*&:�7��I�����(l��!�cªC�Y0�6�V��K[�o<��,����å���ܩ��o+{Ӳ��Y�)r����	�oeL�Μr�
uH�^p胇	ڴ��H�^461,*�:ӭ��i�Z�Yc�0Kn\e�8��EEEhH{E�J�4]���3E�~!ϑ�s�ڞ�̻�s9څM�U��W��kmt�t�(#����Cxu�<p��?{�~�N���Ư����{<�����ou	Û�9�3{/��/���n�KÕ���+f�t8�p�fH�N��Z:A�SDy��E=��A,aL1�t(�<s
!Ǉ#��ɋ�u��o(�NC+���je�B�!�<0�$��ZtP�A<�D0�/��1��a���k��-�o,��|@k�Ie����p�;��ϙ���W�R*)>��"F_%7P�{�Ɉ.�2A00n�F���ʺpy����l�(�G���8 `�Z��.ehzg�����?A,�PL����®�m(���
���Q?�����7M6��sy%[�K��������b�MzLX聴�KH����ٶT��^v�VU�)ڎT��ZG�~eƟ�~m�`�%�$>!�� S�8s��{e�.��մ���$(�B����06E}Q�J���kȒU�H�m弸z��x�H�ɼ�h���iY�i7$�V��ן�d�a�@l`����d�cl�wA��d��nn4�O_9R�m��mGC���\*x|н JE*w�eU�{*�2f�`�
�d���e�;����2!��Yg%�\�J+!��=�]QU��Wzc�!Rh���U�L���44&���EP��!A�*b~`]𓃁0A��y�H�G��,��e���>n��Ack(^HE��06���e1Y�+*�h�H��,�:~��D�,�!��Q�g�� 1=.ʻi�s!ߑQQPHQ�$�+ĒI&�+����Q�X,�F῜«�r�� �� �*�5�IMI5K ��l��t2#D�Ғ!^7AX��ʔ:
D���TRB��\�]�<��9���yJ=4�z���xhXM�h�@��od�#wp,��F��5
g��.��F�t���UYfdƱ������F�P2$�!J�`pJ0��*���Dj�A��j&����R�q���
�LXA<��(S#��b�c׍L�Y��Xm%�[���ق#3���AftF�:�b��$&����HH��CGjL&F�qf��
��f�Al���#��BJN�c-��O�ve�>y�Y�O��<"&�e�?��@�aQ�BPX���7XcBWϕ쳜EEEA rU^�H \��*� @4C�$<�X�3�Kapa�!@���k����M,��1��d�1y�s�����,�f��h�6BH]���t]ф��({ �bTSCU�(4Dw�>��#Be쐻1L�3���ZaSw����Q�n&t�N�oN�84�s�CQ47E�uA!��h�~1!��gy��RDD�88&F�Bg̤��F��ܚh	�c�U�&�$uG����`ah���1�H& h����l�C{(������7$�,�փ�	OA�C���Z$����<c�-#�~e���?��"YbC��8j������ӛ���gή��������>5�����yrw������`{�v�7���h�����/����V?�Qwe�eۃd�Y!�z�5�:E�ϵ�ͷ��?t�&��!���{��P���zV3��(�ﺬ��g*������@��/u���zo�y��/�[���|3.�1w�҇0�V��gVO��_;���է\^nH�(���{=/�����=�.f��v7|�Ư]1��7HJ[Zt���%��! 0��͍�,G�Ä����J�pτg�L<d���C�n3���{1��m]z�����y!�v�lC��i	�I	�0��=Y7���<2�4Y�4�d�:ƀ`�!F���Ɲk,Т�sS�p�^��v�	��4^��B�Dz�!S���3����\��q���0;R�նrͧ���8n���
�)�5��sZc�!��`��!A�ˌG�$Qҧ�v�6��V��U��F�=�8�}=ne7�-7&S���1Թ��������!k|���y�^y�yu��\ePy��A��p&M�***	 ����0ca������dś$���C�o�)O��>
!ʰ�#!UL!Zte��?}�w��ףN�mUWDCD~=�FG#�9*����B܍S=�X�j�껧o^4؛ o	Pe��ޖf�XS�@��F�U�5��$�X#�}����F�&���t����~�ǉ����+�a�eXT6�*��:p|�� �#�s�5�6���������f�
�0����C�vތWǟ2ڵQ�⢴�^�
�8A,��l�N���D�qǑ�Vî2n����*���0�AB0=$.$&"�����I�5JZR:��U�FS���xԕ(f Y^h0t��}��2SC�ɋ@��m�����h9�>,Ch�l:45�)W�"���M��[���^p�QV1��������	>��RY�8}�|��S SCr�(<�-�� �Gó�%G��<`v	kc������|@�A�
,8�ѓ�^$���i����쥢)���������P��I�eÒ��m���,�!9�3VDeľh'NWy�05��m<M�Bc!��000S��{KOJ�d�d��l0p��ύ��>?��"YbC�x��yj���1A,夷'�Ȩ��$�*5��x4�k>�W~yYuR�-B��aQ�b�+T��P� wǟ�9�UY4߆$���48�:0M��"i7�9��k�����&��#��0�foF��=�$d�Ω�fM��d�c�;�ax��V7U�$���p��h��?u�>����ȕ��y���0=:�N���01����	;��O��N�z�lq�,b���|��Û���)�EED�ϰc1��@0�CѰٸPӓM���6Gd<GQ���i�����&����F��� �OĹ?��<>>���W�!�-��-�M��Ky�����b��[O&�IiD��%ԓ�~H��$'�x���l�C��)��i�"Z4���LU��Ű�U��հ��eo2���M�����i�i��u�4�"ZZ[+a�-�6Ţ�����1����-[�>�ť�un�i��yl<�-��nKcR[���i-4��L$[����شZqlZش�la,���[y�q���O%��l-ѭ����Љ��)l��<�$[,�0�i$�L%�E�N�[Ʃ�qq��U�o�<9�o	����Zy�N��q'��ii����lZ[+̶-6���$��Z[�6�[J�e-"Y�1%ԛċH�dZD��]F����"4��c�OW����}7��\n_����'��&�>�����|slJ�ȋ���ޞ�M�V�����>���y�|Իr���U�kۻ���^�߻��4�����I�����ߟ�'_rF���ҳ�>�n��Q�x���u��zr�4G��F���uq�s�G�G;�iyi���Yó�~/qo�}�uM����>�7�N:�#M��B{�Ty�r_g�Wn�{�������\_svl���.�5㽲Ǟ�wR�B��y$���=��g�ˣ���t�D��!sygu�^��zp�e�Fp������P��N�<����)���/�?��9�Ӝ��jrs������U�Ӵ�t�糼�~�&���{��gD����9f�����ƪKI���.7�����ջ����g.�9��U4G�g����n|�;�g�û���!��}m���≩�+$bc[-U3cR��HH[dxD�A�8�vJ(⤵��Ih�F�uX�m�U\m[��Ŗ�5bn*;�`ܕ���Q�e�d,��Z6"�kV��Yl���9%�ٓ�{��^ 97˙�Nϵ!�  _����}��}>��qw���&���fg�}�}�}��}�h���o�37���}o�}������W{�߲k39����V���ﾾ����s�_`C�����.��klDL�a�,��7F���X�ՙUi�$*���Ҕ+iYm�D�-���%W-N����&Z�jJ�J�m"%���2%X�!x\R��e�����H!���TĐ�F��8�$O,� �B�b�S�F�1�a`��^ABK0�ܩu��B��&Adb`��D����� �
A��R$2EI(�N��,!�NR1�l�Z*��#c%�2�B��H'��B1�B�(�&1Iq��Q�AP��2��LB,ARW�cE�V$���1���HD1����BQ�I��U^-+�"5��I��J�DQB���G�Tj��Y�QH�
HĥS-�)+%��q�ʭ��6�ehC��bC(���Jڣm7k.)l����F!��R���Uh�[�q	�C�UQJ&봪�)m��Km��*,����*��T����`�q"�36N,c�@���_��쀤�������ݬ�����G���KC�����3/d�n���W�&d=F�ܰB����D��"#�����qZqL�կ>}�9���\�{M�����vT�잟}|�߰�!6�Ig��@&��&Ŷa�]� ``a��D��QS��-Z5����8�+kN�4��{J��U��^��Df�єVj*��A�7M�o��s���c�f�XQPl���P��h�C�H�!Ġ���h��N����·YeO��C�$]l>+�_bJ:���P��]p�!1�#Љ��w���eT��ﻸ�4��� 1k(x4P�VJ����D�-��ǫ������LF|$31xa߾�t�*�췞�1Grn��[��ZY�B@j��]�C
�&�,�N�Y���~D�ĆBϋ r���;�/,qe�ti�'ьc��@�����nG�B�󭡲K�bd�{��&ݰ� �)�/2d�� d`oD��B��%�/�e��2�&�����%�y��i�$&��u�2@�l��s�8Ԑ��
m��(�E0t�h�B6YA�����w�%onGiT4&%��� `�cx��`�bV�4����� pJ1&(o�(/�q9�JPZ�D�G�C�:<�>Dă�̄$�D,J F�0`p�q�8�щ�,q𑠢X�:5Ny&l4�������I'O��4�a��F�Y:h���;a�6�6Y,�g�:x��D�ĆBϋ w�6K%�r�r�"6�Y�YPqD�T]s�k��9�1��{�'�+E�E��I�ܶ49�(�e�����M8u$�@��O���$���TT�!�����;�o䉊��Ε kXS1YAeP�Ιl22��XS�@��9��C'*��x�\�W��v��U���"4�s�&���;�b;�h��!'NAn���� b��9���f�X`�	�LC!6R�_��څFxE1�3 4�J���ִ4͙��y�}�Ԧ��RjVa:li��t���ؒ5U�Y��tF�(�H4BB�5{�U�nƃA�.�����+V;���p;Q���Q��Ǚ[+~|����μ�,�!����Y�M}��*T�R�@�	���	��4x�\i��P��v�졢B	d60+T3y�!ǃCch�٠���@X��)�@i/�*�����AUTE�&�ϘC��9�p�]��nHB��"��p~dH�h��ӷ��ݙ|om�: b�T���=����ģ��D
!U�KB��5�l�[�0O�)���
���&�&A�78�oirX�r2l� �t1oL:���Ɇ��S�V+,.�V�"���n����� i��[�,4>vT��&N�0G0q��BfP������e�u��^y�ߛ[�"%�$0�|Y���c7�z:�V��#m�'���p���
��T���m�&�����}��HnzDWc��q��!EF�~U4�M4�1��D�M��t�|B��=��S�]8�/�.󘪩t���E>9ϼ��̷MNHg�{au�w�/��A{�t������� �.���:�:S�w�~�M9�9����v��O��	��w}���[v���̮Hq�׳�<e���Ƿ��ުO���˛��
j�(B�����1�5�}!x��YV|�d�%C��D�I,տW�afF+w�X�ճ�2�H�(r�h1��.�C�@��xՉ8ac�9�(���f�l�}ƛ6`�U=QXp���V�nq����`�	����a[T12��#�wc�Ǐ��D�\Y4< R�"�,4�Ҍ����!��zt��sG��svY�KY³:�����	���� ��ܡALlBs�s�F�x�l�ˡ�x_��������%]|�x���X1K���tpx���9�I��!긆���Oej��Xn����i��e�_�|����L�a>,���gМ�9�$�-���=i��i��#��jKC&Z>#�T[��F��i� `�N��F[~���@P b��_#�:i���
�y�l��Ʊ�m�GX4Iв}Rx鑥�G�Ly�GD1a�4Z�ad{¬�2��W
�C�ﮊ`+B�3묇ò�'
Y�Y2R�t�l������������{�ᡕ�@	}���!)�.�1��{�[�F7
��~{�Z�T6Tx�� 6@�1�(ؑ���T���4@4�Pl�`x�g]hmX�~V�����<ˑ"|��@d��"�C���S����+�e���:��>~~mo<�Ν8p���p�{����Ic_NF1�i�b��	$����_�C�74�&�!���:D�PQז:>(l��C(2@��� ��m�T?d��,v���D������w�0:P��h���L7c�9��AF����\d���Q&������$�^fa���׫�J`J�5���-0�`��@)��R�&ɢZ)��q�ҭ��9uZ��l~�~?2]��E:�m���|:0�N���G%<�m�$��:+�'aue��l�#g�<0tǝgbFn�z+�H��@k�C�"�$���#0P����G�X�� с�c������$n͎�(���W�uM����O��??6��u�qǑ�QŖ�x�d�DDb�Z�9]��j-M1�c P���+ el=*J�'��9"s��T� 4i�a����Iy�Fl]A������r:s�_����8�n�\{���y�m�ٰ��CA��Z �`��������]4�.��䌆0<�!�y���S��F�fd�,pE�&�Sd9�B��$��c@tq��;�RV"�0��W�ͶHB��f���a���i���u�*T;Jn�#�o]ۚX�I�?NB:l�e�f`�x���4`��F�}�0����+�{++�J�V��XHɦ���ӌ��������"%�$0�|��}7~�*Is&����Ĺ��!��v���@GNE�����kNA�eN+�v�0h�I�.����M4�@���5����}�}8~�'\�i=.�8�t�D\�g<���!���DV��ϊ[ٴb��{������oς���]��馓��̼��Ī������uͧ��&S������_����O�D�k�y~��tI������#�rfpC�6BC����!-4�n3��1]�M_���6�:ʱ��屌h�"���2�V�"�t`p>-���<���(��V	r�?��y@�s7���WV#6�}0VС�!,I$���Ν6�f*����"0�^U�J�"�P�c@T!��8:��$�l6E4p��*���*�#(0�47d��S�����&�9PH0�:(A��4A��X������e�y����mߚ�[�V�0Al�iV¾�W���iC�Hё��ǋ�O`[�
5f�\+���'A*�!��N��K[�嶵���<��<xGO�"W��J�RЈ˔�M[Fb��V_J>qji��i�b���2�xC~�J(�V�m��cwM�r��9"�cĎ�F�8S�1(���(1~��,��UWw�#Lz{�ƌ�$ӳ.�l�!cDl,��%��cp�(�ql��2}�T�Ώ��O�4�M\��rN�P0@���3�,����ۼZ`�q{����e�T�� ���[c\��0���2��k�
�!Zi����я4��U�+�] �ÏB3xRuF�(tRc�F�낔��H@���>`��c�YZ\2�n�'HM$7��	pl7��A�)���rh��Z:&�	�pг�âx�%�2ش�-�--�%�~k)�#���2������1�-�KĞKKy��0��mL�ԗ�H�.Iid�H���Fҭ4�i���ZW�l0զ�N%Zu-[���V�Ka��ŧ䷘~F��~K~ao�Zyo3��4�"ZZ����ضضX��ZZ{�����O"�aii�ZZ-�-RO-�I�#�^&��׍	�x�&��+ŊO2b�Ɩť�b��[+KN>c	e�ii��im�d���Z\��e����4O���O�"Yōx]#�+�xUxq/�q<):Q"H��Z2�L�[����t����:�gX��u�->OIo��ZE�k��ٴ��ش��%�<����a���iK�/��rH��lGY�-"6��?$L�I,h�D�9_�_��o���LH@��q3�vS�G��{�u���_�˿-p�M�r��|�r��ܾ�
Wz��S����v����|�o^7���e�_~|��V_i��]�ܼ�I���Eˣ��;~�w/�U��P�>�Br}�Y�%��v.�;���l����u�����.���vN.�n19ֽ)�u���No�n�gn�Q�ʙ9O�?2��~�����}�}��ﹽ��&�fo33Ｍ*��g�O���������f}��v��~����o{�ٙ������U|�������Xa8a�u�����<�<���.�311�0������`],�]#$�L6�4E݆��\��F#9�GZ�N,_gI�|��l���䁎��<n�)�d 4P��cc��JL��ￓ�p: �G 3ز,��]�?T{�����4v�Qs��HM�ߌ?#fз�GY��iF7�8j2H=9�u$����ړM�#�����P
��ލ������-�����Z�;X�u͎���2b mԌ�v�8p@��1LѦ��D-�e��0I	q�L�q��d��Dn�vbx>*��Hך���jpa����zL1�BBB�*%iͤʱR���֔���4����-����^y�yu[<V�eIX[lnQ���b��$%A���=(�Ƈٲ���tMe��6�,��.G�n�NL��/ݨpk('�r�H%3���;/�cX(sGG��x��`l��
C��4Q��S	%O顮,Nġ���m��{�Q���CE0��?c�c���L;ltD����5�"�xr>44=�?b��E��hYU�YNW�^��
ٱ��ۀ��<49�N'ō�Z#C!�_���d0|��y��J|a�u�Zy�V�oͭo:"%�����cE�!�&����Θ�޾}�j���Ș��SM#;hlc���/C�utߠ�s�渳�gI�Q�#�Y����mb�����1�.39o�~�QQZR?f��ᮼ���+���;����;��t����(���!��/��o�S��=Ә�Cd���zN���&�Q�k٬�4�9fck�s�U���i���=ܼ�{톮n��^n��x��o_�}#�ygI���;�E�rc[��7�P�<"X���B�h$!�[=hh�銹=�����k�~"4�gs�,x:p4��1À����$�!��orუ�f��#G̒ r;4:�N~������g��Bq��S��z4X샬�l0DΟ�7���Ĩ]�f�s�	.�,�U��m�ɀ������ADx���ʾq�n����"w���@�+�!7l:��|�
QB�ޙ�?�p�`��Ő!��!���%C���LЏ����+�<V���gJd��(�̼�O<���Z�y�yӮ��o�%fF*r�U�͢���$5�Ȣ��zll��#�5��#G8��V�4pm0�Δ��Ҋ�W�����B}8��b6=!�$�Q����hy�O��L �rBB�f�{���e;�&^�
!���46p89��L��8��5��cbȡ�D�x,�i�U��7j�59F���!�0X��Cv@(�e���s�F��R�r~�>�vUl���t�x�,r�b��F9Dv[�O��S�2�aF�r`4=Z�!��[e�m��ŭn��yӮ��Ǵ���8����e��7���_]�7�j/�QQQZ�ݏ�o�N�K%�B��3�,����|�F�!��[pxhqA)ۚ6hhi`$I5�L�X%~�kc�r~$$>�|h�F���B�!�<3�#�B�\2���$8o�(�We��>�gGWk4��һT3�����C�^CH�0꾩[|�6�wU�ad�W�i��W�X%���ؕ�����{��[p���~!e<#z$��۱�Ec�AX[	Cac�f%�*��t�o$�$%��d���KC�͎�*�>G��̶��ŭn��yӮ��{��:�"�S8�b�5�E%�DE�&[^�1�6�T�Cc���	2|K���G��Hgd�Fm����4L{����f#�4D�{ƒ������H��iw���|#����gC�Q`6xf��]'[p���0A�[W�V4��Y�f!�>eV�c��)۞#������Ir��Ruy��81�thp�`�Υ���H解����R��0�(�?�[ez6s��UV�;|�#�ݦ��e9h@�M#o�y��-���ַV��<���:~)����S_�-֪)#�A���ia'Gƶ�i
:���kkujY�9���
�y#TOu����|�����$/�ݟG������c��ZF�t���^��w�9�8s̈��q�������}�sO�f�{�2��Z��9��{[�.�vwe�d�{q���NF��7��w�#����Nu"؏��"rs��B�����^J��/(���2�.�Xd�<vU��g����:t:C%fL�˟�=�L���,��7d�Hh�I69ZZ����3�����h�xk��������h�
Y��@���!d4��� �%_�X�m�IU�a4�2��6�$F�Ԝ�.7|D�C#P,����|HB8�p�Fl�e��e�����a�~e�����ߜZ���y�����:w�GE�y�T�-�Kb\�,�$g��**+BB�=p�$ٛ�!�2�ܑ4sD\K���1�	|}�xFԅ��z�[h��4٭r@�Ƈ'}�2B6Bgpa<�����̄��!Ξن��J�W�U��i=YmW��~i��#W����8H�F�]qm��Df������7�r6��F!D�-�}�N���ۧ!D>서��GO::-�BB�٬3���5�n��4�_CA��~[.��~mo�ŭo-�q�<xGF^l�zZ���ÜAŻ��?��**+BA�7V��	���Bh�3&r���(�g�;]��`�G+V�R���R�����"Wx��%r6h�XA��u�#��c�]�c*%ˣ��J����N��X���oO��l��zk��B�q%�u�l��p?���xt�~ls͑�lI�P]=aQ'�]l!*���H(��h�2+Sl*������[y�2d㌰�?2�ߛ~-kyo<�F�9�uEA�F|��9��ÚLQR��k��**+BA�+��4�d�h�6r�4=6�+B��N4���>���"[>^H|&K��d�ZCd ���;7RU��6uWu��a\V\W��d�zf��O�|ɫ?$L�|q��1�ʲu.�*�r����_}^�����6=l�0C�ɣ�I�'d6B�Q!}�2J}�.5*��g� �.R����C� x��d�!��>N���4��:��c���l�f-�KKu�K��i-#,Z[̶-���qy��尵�Ku��LnKci_&RȲ,�.�%ZDY���Eɖ+�i���+V�~~a�~F�e��a�O�]~a�Zy�հ������ly*��a�o1o1��i,�����Ŧ��6��-�'ԉh��Zi-�%���b��'����ъ��'�4O�<L��'�	���ilZZZ��ش����0�/b�����/�b��y�G�ż�rxt|;%a��,��<K�'����Ú^^K�xrN)RJ��L���Z0�l6��KB�0�y��c��:�u�[M-��Ka��[��Kqy���akċu��LnKch�2�J�,��"�6�Y[-"2���$FQ����;��_�>7�>�u=}���V�3z{I�������*kDA[[w�ɩ8S�kkX��U�9�_:K�������O���;G1�(���9�Dt����6�李Ü������i)x_nz��i�?."i�x�/O�{͎��4Bo��}Ȏj{��`��݋OXM+�q&j��\����i�'���w�TQ�!q�B�~����Ӫ��v���ZB�Ϩ��Q܅g4[q΍�5�/l�C�W�-�mf�%��gD���u�;��;f�/K�_s�����T�s�ܝ�����H�}�|l�3����)��Z��}��M�oZ���;u��Y}o}�r�}3^��O��1w�⓳�:�?JC�B��K�Z���V7��\C�i��"匢j�8���e�n���y�2��+���Y^��C69�We|w�5.��9k����m�b�2�@NT*ܑԔ�%�#I��*Q$B�Ҽ�Kd7�~���9"��Vy�}q���U|�/���w339��}�]�������>�ffs3>���^�K�{�}�����}�^*�V��w����0�Xu֝e��mkqk[�y�8�����VU�N�S��tCj�H�d�\n�
�qb�1�2�TE�mrA�"X��U����dPDAi"h�;+%���7[r1��!�tbcI�!bqbm��Jב�V�1Kؠ�h�J�;	5�¶�X�ŒwZ�piZ�ХȄǍ�!KqU`�Hʢ��lU�k%!q�e�!QeD�!2�!^6X�*Ɉt!B���Y ��aFH�DA
c�A�L��d1�Щ
�� Фx�&bB���"�	Z":T2�5�.(D���� Ƅ2e(J)GI��Z5�umQ�V�!8Z�6A�%�)T�ED(��(ԅ$��bN�Q��)\pm��J8�bȢi)H�,t�Pq���$��6��D���I��q�V
�ڵ�
,j��&�K+nE��&�&X�1��.E\��:Ҡ�u�*���$pDPU�mPH��!H�N����x��C\QQQZ/4n.ɿ;�c�>8���2Օ����yӟ�B���R�;<�8I��SB��}�_Rm��J�����s��yԗȷ�H��ƈ�O�t�i�wT֓�P�9Zܞ+�XDF	���yk)�à�v1��4Ɂ�D`�I5W�K�d��������1���7��ŷ�6�+��ȵ^���
;(!	M�8x��&N�l�e�����9�`����p��s�VT�rdDA���|�oY'��x�V5/I��*0�S�;	�D��x��QL�c�a���ƌ:����AaÅ�hɃE�u�ַ�����F��gR��`�s�s�y0����QQQZ(�F�w�N���M��x���Z&P�9��E��L�"hRB�[�uZW~����Iلƍ#"��v02tt6����Q�C����*����:쌆FáaMA�A��g%J�w��S(A��mu���d��:zi�1pQ�pʗ��ᐞ2|9NC�������_��*�$q�����z�ҾiY6/�2|�u"E�Zw眬�nV����a�m��q���Z����C�Dp�����D���6&;M{�**+BBW�0j���Xݹ������i��Տ$D��i:���
E�	b�r�޾$����e��ـ��CNvI����O�@�<}�y=��5��){�s�EÆ��p�Z��i	8��=�~ �ϼ��{A�rI=L^���ǅ+5�����J��_mV��|�>�>٤G��[V�U��H���֓J[����K��ܦ�������	�����%Uq��)BE�+mW�~W+�FZF_�il�-��~qk[�[�8q�m�9��,�1*_p̨6�IU!a.�Z���Б���Vt򭬦%K��h�u���z���A�$�3��e�:��8N�ѓ���"�C�<�s9��`w��F�D0�O6^��B�m��'D��1*2:Q%��m���l�N����w��&��F��J2�B�X�c ���>�������W8�v�R9I�����7[�ѧ'���O68*HZhr@]Wu�ϼ�y�����ce�mi��ikm�帵���8�-ʴ�CrI-��}�#�!(� �q�^E&R��%ȆWĂ�R\�k�r�Fڑ'-��+YR�Z�T��Y��������$%s������׫��H#�$wX��G�3��1#��{.���T)�ސ��O�N����������k9�w+���;7�+��ou�Vw|��h`�lx��o�:����b�b���~�򣏽&#{<w�{�T��O�l+"�h`�46�����l����/�r��O;0x/%dvh!7� �f���(�v�G�
!����c�;C�p60�ͅ��Y����'��Bs�.��4�1�T�[����O㧼o��[���i��3����f}L�??��w#CD4����YSrF�*P�#pj'��N'�V�����N4�Ͷ������������vZ�3D�eTd��.a�-� 5�a�a�*җCN�O�	#{��J�^1��C�3��!��g�T͖����.�2���!�C�����\�V����;�*�zѶrO�l,��fhɗ������1������\M��hc��CR8C�.p������&�v�!��*�rMd�Wݐ��<��O�2u���ȯ�W�&�>C��;������r��م��N�6�ߜZ����qf���9&�	y�XY4�޽ޢ���$0�S�*F�jxc����_c:̻v���,�>F�!'��ɵf�GS��!�`�a��u��T��yXm]T<n�|mW��a �Yv����Ջl��VW�	�:t�>��.B� q˝p�Xhsn���GL�Æ�K�P�&S���z�!��N��8V@���R���V��dz�vP���ȁ���8�?C:�5��<�V2p��i��[N���?8����8�6�4������E�l�����f�����EU%��vI
e:.��Y���!�%;���荼�Y����Zɫ���EȮ�.ď?�w#�����Sf�jM�˾c�cdD���b+j�u���A	NeaDfn��'�g�֧�4��-ỳ�0@ g�U4��I79��BL�\~6aއc=���H��-+&GZy����m�������F�[˝I����������o��F��ƙNO�WjE[o����wD9Dk')��#�IsVܼ3d���"���1
�����ph���	�q��r)oN�*+�w�a�C�㷢(s���L�7x�;,<m8>�=J^�����_�z�wގ��8X^��Z;�t���[i�rj���>>��;J�z٨U9]���f�˚�6|q=YiV~�b�:8�>�ѦHO���Ɉ!�p��q�@t:66�ʃL��o�L@� xTK&CuH�9'd���9����s�J�uYGu%��ʺss�uD�gLA����w�4G����؜#�W!'��{�7tv�"��JQ��Y���.��f�!;tVi���ڔ����*���0���4��i�o6��Z���t�Ä8&̄�[@HU0)�\
�谓��TTV��ҿl�8�|d2C�^�J��c$���6=�Z!�E�<�Ę�,��i+R-ŞlϸQ�UUk!���t����<;,!�u�`��������������겧�C�!�Թk@��O4~N�G��946Bx�I$8��>x<�mB2�dt�8U�Yҟ� ��Y���,]Wz<����Sl�l��.4�O�?���J6""X�f� �����"%��t�B � ��E\��6'N��<%��a�	�`�&	�Y��N"xL,�DM���~KZ�i�Z2�V�O<�<,�a� ��pN0�H"'O�'�H"'D���t�-��p��bIBlJ�al-�,��,��[2�<C�A�0�ŖY��K6 �K�lO�""X�:'N'�<|��Ǎ,���q�����F���λ�s��Mw]�9L�]��:�x���߻��N)�q�[a�����:{�,���'���9|�R��W�{ߎ��"�~���������)T��z�CGW�:{��s_����w���Uot\=��=;�+#`�В{�9�x�&�Q�/����*�A�d�ϷNS���7��{�*D�/Ǚ:};լ�F���y����=;�i�L�a��.����/7��5�A	�w�.��Uvzz��m���}�%�ӹ�}����r���W�����s333��}�W��U����>�ffgs>���^���>�>�fff{>�j��^*��>�>٬0�a�Np�V�qk[�[�8�8�o�3�e���**+BBk�����:q�QG;#	#84Cm�<�����2i��Yǣj@�0h�I$�y�-u�o|U�i�+ʭ[J�ߑ<uV�ybK��L�bgYcU���G]�E�.�Y����`�=�^����ʓX0Q3��c_����BNC����Ӗ�3Y�񕆈��x��!�Nd�~d���~~�#(�夵ni�����cǳ�t��!���:206�$aa�Ϛy��<��-kyk:p��fq�V�&fda%1�5�qN:.��|&���EEEhH}�f�}19TH�"����	���o_��xi�����_��C�a�=�O��d�BˈV����;�(��f�'J}����2!�����.�j������ev�#�j���s_�5��a�ٲ�d����gR�Y��l!�$[�!��d$Ւ@�,����s,��a�}YoD�0��~ƌ�_+xWm�m����Zmؚ��,�D<��""4ϵ_Vh�WU�#�8�柚[��q�ŭo-o8����o5����y�oxV�r3Qb|tN҈���.pS���B�Г�X
H���ڱ[=�EEEhH?_f�xNd�s[��g�j�ӿN�K1��""p�35���{=�g���^�;8gzsm[/�Þ��}�o�uVG���K����㗜5m����o89�M���=�F�ȕ�L��Lcı�/ɬ��{�#�t�,��������TJ�(�y�����������]��2�����t ����0RW��f\2�C�����s���{�K�w��-��K��{����lh�}D�A��.�\>��Y��C1C Q����}���oF���nP����t4����[&;m��v�AB�ک�YK���	��/�Ŝ��n�����P��N$=L�ka��:'�e��N��[�Z�Z�q��8i�Ω(�ՉX
�oތm��К��^+��� ��ܔ(2q�XhWC���/��2�C,b|l���I	����V0[t^��j�;��I�D����C��M�!��;lSx��:J��I���߂��B3�v� di�|�r�d�d��mg�4���qU6��4�C�0?s�
��lш�I�އ��5��&ǟ6��&��&Q0p4F�?Hω	V�Z���u�m��2�ƝZ�~qŭo-o8�����U����CҮ�w�Q���(�2��"��U%6�9�>�c�Ԩhx�������N�0Y����#���ö�����b�CI܇��t3�%�C�?�Ø�q!آ�����m�2����:�nѮ�&���f��l���e�F��8���� <�AG �챣~6B=#'zٻi��O6-糫��p������ǼN�IR��p��C�N��h9��d��y�2��Z�~qŭo-o8����"�b_��jWѨ4��"�~�TTV��[+(�hΗ����>4�G�n�B��&��89T�R��!�F��Xӆp�78����zy˰�gI	g�X�FǣA�q������~��6L�8h2�h�i7�'��r9*h|<�d�I���^�^ɮݹHg�{|��?a��ɧC��,�Z�1"��5U��W쯏[F�a�߰h�HC<ӽ����FM�m<���8����qa���|i;�I�&�R�:�8kb8����ia��s�C�wz�UuZ;m�F6��#�cu"�YDJ��EEEhM�zo���ڿj���N��/��uN3��':JL�=���9���×�����K�u�Lw���i�ߖ���Ӿ��e>Os�W֧��Z�5�0�����x/��(������`QT��Y�Op5����Gn-�u�m������U�RT�ѧ+����~���.�WVɤ��W��r�6�~W+�]d�ߟDۉ&�4�d����g�m~._�@��V��e�
,ï�i�>;�D�QXJ�>�U�z�[Uu�L���|A�[#wrF�������2����N�fHB��4x�x�!	ɓ�ϗ\���Vj���0��|��yn?8�ַ���q�q��Ï4S�i��I���"���Q���{GL6> -��޳L�K�1���Nz��!D%yJ�o�y�*��2lv�a�R�6�X$�$������Qc�܏��&3�(���O$w#K��~�����_�)2�z
�e#���J�������oƗ3�Ib^ό�OóA�Ócc��S�I჎I�>�7��q������[H�8��h<�4q�e��e�<����-kyky�Gn�3SV�1�/��**+B>����~��5)�v�8�Lg�2���>�~U�LXAb̭P���]��T�3�#�8q���!q\��;ס	���%�*�;+1!gL�x��ݽ:9�1�>��=h��FG�̆L�l�m�2�9Z%V��r��D$�ړ�IT~$������]2d��M�͛?�Β�6
g��ܨ�>aŲ�֟�[�qŭo-o:tGFp���0X�yIFD��ie���r�[��&������a�ԕ:����I�z��V�0F_���<~2|�IU$��a!�X���a��mĂd��-�A���5�[���E����-�i�?G-ˁ��?�|�قNA�l������u��Mw)��?>���I��R7&F̃oX�c�a�AIA�܏L;fC���eUx~���R�|���B#��3F��믚e��N8~ �"&�DD�K(A��<"`�����(ACb ��Q�8&����Ǆ�0L<abX��`�%�"t؈�,K:P�D���b"a�HP�>:|||ukZ�|��O>y��<�-��=$DN��"lA��"X�`�,O	����BlJ�� �"B%	�#��g�p�]m�Z�[�<y����xD����6P� � ��D!D>:r�P����i�A������r~���ھ�~*|�-���
ɽ�Mϓ�9'��齣ԑc\����A�|�_wT���z.'��k����4w��q(p\�ɟs��h}ˢ�k��:��E$���L9��j�E�!Hn	�����ru�����e��Eύ��$�!Q�A�l�4�9�%9w'���jC>�J#Fow<�O(^}�;�|Ē��};�]��ɾẹ��*�g[� p��m���e#bQkdN�c�#s�\硄���W����L���P}*I����'�:�-��m�?�W>���";���G�_��LM����mB��򏄍�jh��K?��_}��v4��ؚj6Z[SV7���Q4�a^9j+gwRڙ�hVԔ��I"c��R�"NU�����Wj��!�\�H�TWv�m�k�hU[kq*D����P���AV��U!DݱH�W����9�I]�{��\�ʛ�7���Ux����;Ϸ����Ͼڪ�W��yϻϷ����Ͼڪ�W��y�}Ϩ����g�mUz��]��>�գ!�a��4�qn8����qa���q��PJZ��kS55�mV1d����]�H,I����3s$DQEZ�L��u�b��m��\K��8��PQe����&rݧL��\�´챌L�A9H�TZV�G���ZF��1�ڥ)rdT����$:'Y	
�B1Y��Yn�eYr���A��f�c��(��1d�q1U#�eH���
J2�A�+�Z�M�H�"�-��T�J' ؋:Y�DK,L���MX�!�\e!
: V��<y%�� �T�BH(Z�Fe�7K0�wq����kc���iFV$��!	���1Y�-�Z��jժb�lm�Q�]�RV���Q)e��D*�eb��(춴Yq�(�͏f�ⲍ�V*��\jѩ��A�:�V�YQC-ĥU��%-q�j*BD"Ʀ;m ��Z��թ�
US$q��4֨��d�o��**+Bd�W������x�n�1���<Y���\7֏l�Q:�%:M�Rfl�.ٯ��e\=K}/w��p��]we���b�<t���wާP��7��$���<^n����\�~����q���yR��*[��ttޯ�������{i�����;����<��:[��i�|Oņ�#�z�Q=;Ӕ0��	���}[�/x��l��v%������H�K��~,���B]�����t=��ڹ�߈=��>tBB��������Ό8nt8Ul�g��W��~�\Q�65v3��>��
)�������1��h���m�e�β�m:��~m}�����n8�0�{��1.ocA���B$���Ow���s�˺�\k.O������])�BD�Q
��X�D���CGN��؉H�W���!���J�W��r�EgA!�~<�7�|�Po\���.\�/{���ĳp��d<?d��Ý�� `�l5�f�L`����`�I�� LE��������d!j�-�F��:�N��m-���[�[�|'�,��x��L�o����z�P�N�**+CY�s���ۘ¶r?��ǃ�[p>�$e	�q��!n�?[&Mg�+�gO�:2S>�:&d����������ߞ�"��M�/��\B�������zc |@�}0z��,����;�`0^�X�L��l�����k��_M�|yɀ�0�&�Tt��d,�5��<���װ��ZRkzq��X���0<�ó�C��΍���A�4QӅ�m��-��������n8�0�>��BFQ��
�pb�óQQZ����ΒFp���N;YJx�q	!��	�e]<gA��|���sm��|���ʖ����$,�JXE����K��]�w$�C��D�S���e�I��AG���08���`N�CF-2jk�$����~�%��G��z��ߩ�M4��79��\0[����=Lx6��'F�l2x�^�=R��çD�ѳ���nS�FQ�y��ӯ-�������n��0�n�ﺹ�e�����q�]�J0m�j��(����'<���k��T��[q��#�"�ax��/�����o��{\��WI�.�{�ʿVt��~�ߤ�����zǴ��b�:l(s��}E�s�6�{S	(��d�t�!�8��c힣	Z��/�5��/}��&�ھ^��S��r�������ntbl�</������Ϗp���ۤ��u˿���`���N9}��P������|�<0y�C�͏96���2!}�E3��fP���o��H%'���J��`qg��I�G�˳a��CZV��ja��=�/�#�L~��Ǆh���5a�ބ>8�m-�d��qq\<���Cᖍ��u��ĕ��?qa�̭�ߞyŭ�����u�q�ҫ�'2���T��ʐ� ����j**+B��N�Lw�>�\���zJ>���F����΂�r<$���TW,���x3�M����Āz_a�R!��U�OWM�xV����U���*M���r�~�I��.IS5���ZCe��S�L�0���e�Rx�T	.�i�vFCo���1��K�?q���16U��Cg(C���=��$:Q<l��r��#��ʹ�0댶�ku���[�[����=Ϛ}�-r=�EEEhM��Wwkv-�	D�g�U\���;�\>&F�ܟ�Λ���v���!�F�t+�P���K�����	+��J��ȴz6�S�W���`�;��Nh6|Q��v|0��=��L�r`����P����<g�������|�P�Ӆ1T�ㅯ���	*O�ʐ?���{}?x!i��cï�#�c�!���e�[~~~q�n�ռ��㮣�9��%��i�j�e�+�66��К����V�H��e@k�
�xbǜ8cp��?0�x�S�Y0��D�c0>����p����/�w�㒌	C*U>�q*�!���](�*��N	Z~�߁Snd��/�j{�|)�=�����1UU�[E�t<��9��x��p>��*t��R�8��?Y��%U���v�N�]|㛦Ќ��4���m��康V���B�<5��ʞ2}U˲�s\�Wgj#��^��jb��E2wy]W�yӝ.J��W�r%�x�QQQZ�o���������������|3�u��!Y��gq=��Ό\��^|p�{~;zs`w^?��o��9�_�R���V{m{:N��y�g����Ư|�0�z�|�]K�=�;��9d!��CQ۳D��C:c3����!0�����t�C�σͽf d)�%DI;Zo�m���c�4�Q�`e���6R|�(�N˯�JцK1�Q�F�dzg0�}���E���'�C&�T�r�0L�:m�Y$y�����G�hc����o�ܺ��Wbܶ
��|j��Ba;�݅�]��_j��Ul��[-��uŭ�康��󎺎0٧؈H�ico(2��TTV��n��P���X�h��x�C���[������M4����f|���8c����5�S���I�%BI
"�jSy����	�z=]�m�z+��l��C��Iy��e���X27�JlG��F�����&��b�]�\�FS��d��P�l>���õ�:G�;��Y��t=^~�xl��+e��i֚a���<��<��<�,�H'N��e��"%�<C��AA�"%p�"lM��<%�ɂa��0L�0L舛,K:P�D���b%�I�B�؋�yŭk[�qm-�-��e����"#�%��H"'�<"&2YbxN�8m�l�	BQHAA	A�ؐD��Y��0���VZ�k[Kx�o<��<�|��Xx��Ǐ<ydZ"!���$�\+/'7������D����E���?�\�n�IӖ�w���˥7�OI�O��Uo���m�ۛy{}ߢ��m������v�-�����d���{/;�~�G��m"�/c�c�B����w�;|a�-�&�y^o��WϹse�n���yN�y�;�~���{O���ظ�������s�Y�_n[��Br��3���ߦ�u&Jͳ������~�U|��^s���Vfffe��*��v������333/�U_+�W��9��3332���U�Uy�kWr����u:˭:�qkun-�ǎ�>>!��!_e����'�ش�I̸Yyo~��H3���s�<k��������ЕVp�jrV��ä��c�u�BC��ɻ���^b˞Ց�LT����W�[:H����ю�8dw��IR����k�鱅�O'y��<$��3�[��2�:���8:��{����q+���5}7]�W�0�b�̺��-�ŭո����x����ө���E?H�����yj�Ƥ=7���s��TTV�6<����`��oï�o�M�$�T�o�?%�l��K&a��d;O�p�p�GE[�G!����!�:�|`�l-�bf|UD�<�dd0|p,�Ev��m����{$�΍�&����ɹ��q��>���3���D��6x!���K��hfǁa����^��v��f���~�~#+l��l~Ke��������[�[�:��S���ͼ����q9��Ip���5P#��$�[W�&;8�+c7\8:K"��ě�v�)j-�.�m���6������'�K�g/n�_���ph�~��)�>9�Ga�����}ct��~�)��(���ӝG���n��B߽�o�����t����Q�2�ѯ��g{ݪ�z�Ͱ����������v������Z�Q/V��x�%u���O�3�9�>��˞�~5g����k�K�{���Ҵt�;Z�+U��=	�����^��X�]z�to	�^S۰��?S�e8q�n�4���U�2׼����?[�X����Q�yŰ���FG�}a��'I���J�U�x�(�N���yל~[�mo-o8��N/lET�"��k�/&���f^��QQZ;E=�$$�;��Md���RBI��l��X�f�C�?d�I&��qbI	��^����1���	����ú���}$�h�聸��B�S#��ͩ�=;G�VL'G�`\�ptnx�ś�:�������.c�+Ą�	u����� �
J�m�}�!n��%A�c���8��J�{��!�$$<r�8lm�	�cu��+ki�~�M�mcIl�����[�[�-o8�>�SW:�X�ԽN�h����0�L��F�T%J'�[��m��Ak�q~w6��)�M}��2pt::>��'aoIõ��}����5�%އW�B$V��l�k�p��WJ-OК�*⸕��ß����A�#��C�m��a�8�ǯGÀŅ�FI@��x-�I\8��&�;��tt94<�
2C�q6�m?<��[�[�-o8�x|/`��O�m�[֚i!U�\�b**+D>>)+��0p<h���d�2$2��ɰ�A�]�Dj�\�~拦$���5�};mU?j�����x��̄L���Q���Bȟ#������}��.Y���|2���;�y����.C��a�֜���ƹByX�y���י�o,���N���]j{�6�2e�m��l�4����ukq��ucix����Ύ3��b%�K[��h�DqZQ-cQ�(�-J1ciK^F�2 J&*ƒu�$'mƉ�!ĩD\����m�+	Geu�kgs�TTV�����>_�t��ܷ\�Ǯ^a�u���K��c�d��bf��۝��Y���rp�C�{6l�Ş!�K�z�=��^����a9��3��{3��պ����o��h�I��#ec3���~!����aG��IrL�4^�1���̑������j��e]#������8_�[��~�OM�1~#���80=�&G���x�>^ϵV4l�����;4���d���֬�Bj�n��Ր�������Ӈ7I�-�?�6{��%��\3N�A��h���4��~q�n�n<��㮣��:zjN��qe��EEJ�L�9vd����m�:�V"�����pz��ѡ�^����U����.^pB���¿��BM�#N�����A�m���!���_a	���� H8�S�*IbrB�Ŭ���sV�9�W��`&��[cpc�24�\2�Ή��<
p�#��I���a�	WgÄ5���/������`t1���̐���q���~q�n�n<��㮡��W����iŒ��Ae/6V�j%-�9����clm��-�m�WU�0|�)d����sNi�a��?�����I"J�+��Y�<D{��DK9S�RϿ�G��J^s��/9æL�z��8Ǥ�#�,�I�+J���ڰ06;v6lkAb�beq��*���'��P=�e"1�����y�'�I��%vr���}M�~acil�����[�[�-o8��?��%��cD�UH��I_ұ�*+E��0��UѲ��_Հ�&��7����s��,���ZNY�Q����Rj�Q��p�Q��&�*G_���yf)���mW�>WM��W�ݏN�ph!!�ej��NOj����"p)D�1(�I	Z}����Rk�p>zi�hpS�0: R�{�h�{ǋٓ-��T{�U�i��m3�8��Kiy�y�'DDL�"A8""&��:'D鲁AA�F͈�b'DO	�0�0قab&	�`�&���Bĳ��P��,�JI�����,DD�>,����x����0D{""&	��H"'�<"`�%�'�ǎ�}��(J# ɤAI�JbA����,�Ǐ<�Ͱ��疷�Z���|��K<x�6P� � �?����/��'���.ϯ}�mg/Oל�۩�X�}h�P���������-O��z�uM}���w���g��};����/�o����ڵ����U�;��|��$6��Qr�EՐ]8S�LJl�������>�>�n�Ud�����ӲM�kέNs�\�d�}�8��;���d�rv�s�m�aHpo~�uv�}�1��iy4D؊��9��xY��M�*�OC���rP�2��_:5�znW�TJ�g�G�I��6w޿"��'Mc~|(��	ш�QDj$�rvpP���̺���l�g{���*�fu+�7{��߯>{�}ϡwS���y�s2绕�_o��w�s{��NR}��{�z[8�G;�?���|�v�D�ш����5͓c��1��CM)�DyZ�8BH���T5�J��7X�U�i+b��֊}F�D����i����Ah=&��C}Z��Ǳ8Rٍ�)29�?ƻv�qս��̺��=�kͿc�EU[ZUy�s��陙���}UmiU�9�}������>�������>�����g�UV֕���k^��]G]e�]i�V�[�x��ǎ�>>!���z��r�Z�$]^!X�,&G�u�4�HQDU���'"�+YIFVĥQ(2Q̄u�L��m��x+a*l�M�n*�#vA����!DC�P��P���M�	IjW�.R�x[e��B�[uB�V�M�m�ݎ$V(�	�ABTH�$�W(�c�+�C�v�H�ldN�:�K![,h)]1�RB,�Z���+i\xʢe(�آ"d�		2�"�fB(1�~ۓsjtm��e�FP�K H5��FU�ҊR�*�R�0�AB)(� ���2��Q��ʞXG(ĕ��&���-�c�4\q��]���FDB�T"�R�nV�)#-e*��YS.UD���i!�Z�p�T�Zl�����1!L���D�I�YR�J&ㄖ�6H��P��d��ȑJ5k���cQ�	-!Q`�#C�V5FW��/�k�f�??��jm��r�[�3�e����孞���l��׵��!e�������t�G]�Oa	ݔU�N�a!������s/{�͉�ǣ=ē�9KM��M���wy�I��sךw���c�a+�I"�V�.|J�`t6l����$�ܿ?)�;����u�|;%Z~��&�1�{�˺(.�}�3�.]���!�=$��,�7D�î��[0�ztO���2g&�m���04`v94���J8�R!�p��p�t�l�Q��vh��L����s�8<����4˳â��87a��t�g�\iן�qkukm��um�V4qͩdj-�M4$%��=10������\.�~5]aZWr�/�x4����a��l�%�z�we/6>c�C��$>�0�=
�F��#�'u&��ve�x�������͟:������b�F�QD-d�V���
B��%Lϳ��8j}}�$��U��#�ٴ�����$'$��9���)fΟ<3���������(���6٪�90�d�:�.�����ykuk|����>��S�_+טʅ��ۈ.�BBBXl��s(���>��1잞��:hc���Τ�8��>p[#����w������'|;]!J���^`���0��ɇ�p,�q�!6pd���Kf��Ƈ�׏�q�In��x���ɖ7+a���F�S�xvy#��C>���U�a��n���>4�8�-��O��m�庵���󎺎���.�U��X�1�M��		
%=:>ɰ��ǪPUV����xύ���V6���LD�+�V�c:G�R:�������O�{RB�,�4�'a��ä�I'^���Б�^"��e��1�s���F��0<�!!�F�/,	�F>�h�Q8XC��A�;
p;;�6l�kt�e���k�����93&͗]���|�?:��/�8��Z������um��y���~����Q:��I��r��x�Hh㘩Hh�[��8p��/9��y�'�		#�"O�U���i2T��tn��*�UN�/nş�����~��{�f܇[�5ϼ�\&w�O}�<�(|3�d'Kwǩ=�2=��=�@�~�!ô�Dо��_�Ǿ�p�������gK���=��}��rw�z�k��ߵBm��i^�6��׫ܕ?4�e�-�)G���ߤ���Ba�6��9���FO�~�ĳ/�yi�l7��A"�J��
��pM� t:1�|�PA���}$���:���?_4��tn�T���Tj	�B~͖�8��(i�܇�ð��B�#U�b��t��~[.2�Oο6������ky�]G[e�|���/7�>�G	Iaǵ���!!!,>��SB	#[M�-<�$�0aɡ��}�X�MY	$V�q_G�+�����Vg�9�Ͼ�U�Sӣ���3����j9�A/��$��J�g���6�j�2�!�
��ޏ�a
d)W�
eJ)��=,���5~T�H�0��/V�D�x���2������:�����U.U�������$�#�m�_2�N�<��������um�\��b0�U��&!J���_4$$%�D����^4O�&�H{�!B�'�Gd���K�m��&�T̄H��qX>h���'$�O�����{�{)2$;Z>��')Hi���?b3�ץ~1���G�J �8;X�u��8�N�����O��
�B�~�H|�뾱>=�*����������u�.��N?-��խ��[�:�:�/���fy�5�̻ؑ"Jim=XW�]�Y�4�~1b��:˛������tvһdH�s*��Ԉ)v]�sa?	^��N��cAECm���͏��Ci���
�Je��A�\|А:.���A�V��l-��wWp������ó>,! �;�d�QS�C�����$BD�X�FC����:�l�����&��e[/�m���ֵ�����󎺎��jL�<�-�l��bU���%�9W�E*F�(.Z��Gj�-�Z<��BkZU*5,�V�rYM��脄����u~}�����ᳳ�n��d��]9�'���*�'+�g���f��GI����	�R^B<��}��O��M{���{8�s��J�.E���Z}��9�Q�΍���+VG`�v.���A�!.�J�l=ƝvNj�y9�(i��,I*������.��,�K�fׇ*�h��߉]`���HN��!��`�~�ӑ�~�\F0��!�y�δ��BnI7���f�k��ڒ�7M���gզղV�$�EY���j��#�2�-����������[�:�:�+�=�be��^�"D��>�m���,}��G%|O;^bY��~�rE��*�4'(�_�IU��Ch��?8_h���I1��9�7����$�ueF�f����#\��/�\l4hvxt��|��6���!X2������J�R��,���Z��
_ٕ3��2l2��v��~CF�t�:pç���0H""tDD�<P�"P��,A0D�,���B�A!blCf��lD��<�b&�0L�0LDL,�Yg���(D�"&	dDJ ��'�N�"%��8'ç,��-��mk[��y�<��fDG�xG$L��xL<p��7�P�؛ �H �&�H��؍H�NYe�Yb&	��D�b'�||`�	�O��ae�<x���"�-i���������$~F�{{ܧy��WS:��|�M\�R��<���ҋ��}�}���}��>��>�E�g�|Y�>��o)�ךuz��w�;��-�>N6/�5eָ|�����U�
i�����ēM��~��
zp�p���d{}f��}ʤH��]9�u�?{{���}��Y��q��(��%���J�ƙ�%s�|���!��W^|�5�Ϡ����/vq^������(�ތ��p�U�Ķ�.���+>�ΜN�G>����o�誫kJ�9�q�������UUq��9�q�������UUq��9�q�������UUq��9�k֮���ˬ�Ӯ���n�o-��㮣�2�s�"Jy]��Gðprn~
\�k�o3C��g��GN���`
�uU�D��\��l��U85�Zc���{��#o��n� ��6�,����� ��#:|�,=���F��+��e�S��~L^�R�Mh�ڻ�,p��<p�,��(0�0:�r{&�ggݚr����F�e�^i��[�ukyo�󎺎��]��s�F������JW_�I FA?�����Ƭ�rF��]�5M�öUks����S�$������V�$8F0�`���?bǥ^��G���	/���6Pg}����J�\���B.,�?����J�B�>�IO^0�J>�y�HI��9��� Jr��W��4V$�1#/X>tg�W�����#���.���mo-խ�[�:�:�.�W#=����^mn���AK��h��{0�����wh�d-s��5o�Z��l��c���-�j<��$�@�Vw�M�gG��]����t���������gM�;i��o5h���/��q��w��gh�ҷ���ȝeO��[�N��ݼ�����s��~�N��H���%�����p�{�z�=ޝ�\�itwE-Ʃ��{ǌ���<�:<���H�4b�k�;́g�O��۟@��`}��'�E�hR�iu+��{6p<t������Aᢨt����:k��s��b*JF�a�		f���(t}q�d�u]��YM���6a�Z�|�m:��kyn�o-��q�Q�|τ��[�����SV��9�@�1�>ԒI���X8L�����5`Y56��$$X"y�?:k�9*���������e`o}Z�O*��=�!��@�t��T��j�)�}�Z���/�iw���n�O`������:'ӡ��MUO;}(�d>hx8~6Ѭ$��7�/8%x��UXE��u�+�V�Zl�H�̿2�O:����ukyo�󎺎���j>vT��[����MIq���H�s��ޢH��r{�.�[��ƫ��q�Ն��BI���6�NS���;���Iei*_E��	8H��Vc �1�>��vAیIu&$L�������z`��;�(������[��M@υ��$V�w��q!��G�]o:h�(��/�y�^y���V���o8�댱��1�e�s�z��]ܒI�V��c^)�T&��'��ajB{�Ǵtύ��kyt��q�ǿ	h�$���/�����#�'|���'
`���ۮ{x��74L�:��fI:6/&t�ߵ����(}��4\�Rٳs��M%�a�m�!�*L@�F-QAPp$����R�f�c�����̭�Z[��[�<���]������>�;d��u���u4E�Q�1Q
j$���G�aFT�q`�$]�[\�s$��%,���-|�I#ݝ��3��<�C�w�m��L�p���C۫0�;/X^�޷vCewdO@Ol);��Å��d����e׫s����T_}�f����.���Ԡ��9��66�J���9�_T<�������&H#��K%��/�O�6�6����|�!$󱭼064QMtza��V�D�m����.�|S=����t����W�4�ϭ5?i�R�=�f���~t6�l�=�P`���lWǿW�A!#�&��m�XޫZܮ�:u(tuқ����6d��l�����ߞq����qm��W[,E�*�Vfe��I!7XE+u�{��K��u8�;���$�Wkn?���!Xొ����B��)ֱ�>ɱ�m��c@�i�+BԷ��e]�����!�T䞮pC�|v�NA��[�~݅������A`�����g������tϪ��G�1	06��í��Zv}���|:6O��x�nH&�$��Ļ�ٳ猰��2�-��m��yo-�V��l��K��9+�i(�KX�Ãʪ�\ ^<J����Yi77��$�D=F��D��B��+�d���ˉ#m�*���QhԲ���KFO�-0:NWjW�4W��x�ɣա����+3&&D��k1۹VF��􄀝K$.��o
���?����^x=P�*N>��'�����̿��VrLՅl�|��-K�T���������o�X���g$�Z
�[���̺˭8��ky��弶Y��:p�ǯ�䡱�[In�M[ޤ����#�������a<TO��C�잔�w�c�O����J�waXWM	n%��Y��h����i����O�sؘ`���ѭ�U��|?F�8i����Brb��@�m�U
ۇFI<8�����c��}m������R����J��M��.'�~m��^�Ϝ�k�cK�k�0%�4Ѻ A$Qh�	���|bҘ8�m� t�bX�FH���t�ؚ�iZ�KDE�&--&�E��&��4DE�AD������"&"&�"i�H�&���i����ii$�ΦnI�$�4-"$���4�D��i�	���I��&֖�-&�E��k%��I&�KM�����$��4��i&�I��H���kLZhI-"M"Z덝d��K$�I-�M��L�Ki4�id�hI-"M"M$�kKH�H�I!$�k$�H�I!$�I���ZD�I%�ɴ�I-$�i$��I4�4�HI-"m4�I&��BI	���M$�I$$�:��I$�I	$��ml�BI	$$��m	$�$�$$��m4�2D�I$�HM���HI!$��I!$��HKd�I!$��HI6�Y,���-&�Zm$�I�KK%�	&֒ME����l�$ZZD�M,��ZD�M,�K$�KM�"Ih��%���$������I��Y-,�����i��i%�"i%��I����I��Q"�($���%��Ih��KI-,�&�Ӧ�4�M,�K$�k"i%��h���"iih� ��[I&���ZZD�M$M!-6��"��$��֑$ZZD�4Ŵ�ZbhM5i����hu3q��i��i�i��	�4�D�I4�M4M1i�M4��MM4KD�MLM,D�4��4�Mi��i�C��4hѣ[�����M���L!��6F��l�f�fF�F�#FC��24m�#LF�F����٣CC�8�vu���JZM��gn��M��h�4i�44i�44b44:��؍#L#XF�F�dh�5�F�h�l�#9�ѿ�g�f#[25�#[b4b45���g3di�m�[����#CF�hr3�F�h����h���F��X#CC�\3��44i���fѭ�i�5�F��G5��u6phѴkai�4���k#9�4h�ѭ��Ѧ�ّ�ѣdi�mlkh[l��!��3hY�1�f�����X!6ЃBas��4��m��m	�&�&d&�ɲ�Ml�̚6�ͦ̚����X�[4���8��k2hi����i�����,&�ɬ&�Ma44�i��hɠ�,i�&�&�hi�&�����&�&ɲk2k	�&���Mm�M���d:ɸ�i4&�kM&�MƓBl�I�4�ɤ�MM4�!4�ɤ�hM&�i4�d�i��M4�i5��l��q��Bi4�I��&��$�k&�M4M4�4�I��4�I�КM4�5�Ți�КM&�i4�d�m4�I�4���i�ȚI��&�ki��M	�&�i4&�Bi4&�I�i�КI�4�I�6I�4�i����i����"i����&�hM4�4��M4�I�4��Zh�-4�I�4�i��M;�ƴ�d�&�i��i	�hkB�h�DH�-m&��DE�4X��,��E��"�hȉ�DD���4d�E��-E�4HɢȴZ,��Ț$Z2Ț$-D�"�d;u��l��h�4�F�B�#-�E�CZ$Z$Z,��Ț$e��H�,��dMFZ���B"FZ�E-DFYBhY��"�i�D�dZ��h�"$Z-	c��FZ-	�h-B�MZ
CZ&�4i�45�hMh�MM	�"h��ɡ4i�Bhi�Mhֆ�	��4m4&�4&���\n��\3�	�Mh�hM�E4kBh�F�F�kCZ�BѭZ�h֍�ѭ��h�B!h�Z�D�h���m����#-�Bh�De�Ј��h��h�hDe��&��1h��1h����SZ"ki���������D֓o2�x����S�2~X�zд�����8���f���c��6դ;�c�W䙯�����_�s_���k���������HT3�:��������X ��h�?�������c����g���k"PNP��g�&�_��>���eh��g)�?�5���`֓�a��g�{��(��E@�T���<O�o���CwM�ۇ�67��=3|��m�����v���v���X��?ؐ�?ҤJ]E}������'����n��|z}�����=�������ed�{��<���æ�}��>ϟ�)?���ȸX-���ީ������I���E�F�~�èi�?r���L����XLG,l$�������?�Ra�$T��*X�*�  ��q�4���RR����v�����1�6�Y�I��f�33�v}�h�ۄ2�@C�(���g���bV��<m������M��x9	��&3f�ClnBY���Z6�r ܇#fc���aBF��Ov���}ͽ@T?��-xM�_�o �g�B�#���� T8��?�?����t�a��O�����Յ�l_�����{7����5� -?�h�����f���N?ܯ����i�?������:7���z`�V������>��?^���Y�޹<|��7�{N{q�o�z��y�&�f�l6��Y�Y�M�W����x�����N�z?��ݵ(�W~3N���m�����ߥ����?�l�S�2�JG�:C��_��r��������6
Y���(����_��"G߀0��Ȱ%-�2ATB� 1-���l �BX��Ţ�#A)(b�)
�ٰ[�"�|����7�����8�r�y(O���x�?�=A )�����}����^�o�o-���uݷ���G��=�{�>�7n����g�>/?���{[���M�����#g��9�u���N�>�{ϵ��s�7іmϧ:ςo�s}�no�n(
���a%��J�5�����9�p�MYZ���mM[V��Z�5jիV�EQZ��e�(�V�SV���j�څjQE�j�Z�SQYX�[V���F��L�L�+5em�e2����ڊ
�b��V(+�

ؠ�V+�
�2���b�AL�b�X�V+��b�X�V+�jj�b�X�V+��b�F�V+��mL�jQ�jjڊ�(Օ��)Z��J�VԬ��J�Z�)L����ڲ��+(��S(�QJ��R��mJ�+(�R�)�)B������Z�ڙYJ�JP�eb���++++++++(R�������������������������++(5
�M�VՕ�+++VQJ�Օ��emYZ��VV����[V���VjV++SP��)Z�յj�j�)�����ej�)���V+j��+j��e
�������+++V����YYYZ��eej���Օ���+V��YYZ����b�5j�+(�[V��Vի++j��jՊ�e�jڊ+jյjڵmYYJՊ�VQYEj�j��eV+R��J��R����5mZ�j�b�X�V)�V+�mX���V+�X�XV+f��b�X����
��5
�5eb�[+�
ƭ���m���l�V+�����5j¶��e2�2�5e2�J)Z���52��e���j�[+5
)Z���B����YYYMY���Q�Vj���VS)���m[V�V�Z�V�jիQYYESV���e�ڊjԭEjիe
�E
(�ڵ(���S)�j�յ�5���(���YE�Օ�j
�b��V+�mX�PVPPPV+�5b�[QX�V(Պ�b�[+��b�X�V+��b�X���b�X����b�X�V+��b�V��ڶ�MZ��VV+S+R��j)�SV��Z�Z��X��5ej�jڲ���V��QB�څ5mEl�J�j�jjS+R������թ��P���)[V(��MB����P��(�QEՊ���ee5eemYYYZ�����ejڲ�ڵ+j����+++(VVP�YB��+++�eemEP��MML�b�LV�j�QX�P�Se6S+je2�l�PV��)��VVթ��j)����e
�L�X�Z����+5
�ڂ�Z�[��b�AAX�PV+��b�S+��b�X�V+��b�X�R�X�V+��eb�X�V+j+��b�[VV+��R�(յf����VP��
V��J�VQZ��e(R�(R�J�VՔVQYE��)�VV6���mJ�+(����(R�(R����V�����B�)B���ն�����eee+++j�)YY[VVVP��YYYYYJ���ڕ��Ք+jն�յejjjR�ԬR���e)�Z��������ԭL�MJ��P�������w���>�����m��~��O��q�Q�����	��������ƨ��V����$Ę(�1dP���?Ű��7�Ha �?C��������|d�J��g�`l�8[���2�* h�~��j��JH��7������������?�����~�� �H���ّ+J6��9�q��;��?���or̍���Ƴ~=����2�O�����:O��G�O�L-C��ƗO��Sm�xo���?�����l�?p�7v�f��ǧ���"�(H6��n�