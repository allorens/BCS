BZh91AY&SY�PR�H_�@qg���c� ����bJ�}@    Ϩ(�)>��F�U��lBk��P����`�*&�U���RMaRхH
Km
���&[�6
���	m`[a�]6KYU�-eT�$�қV&��)�
�Z�+d�l�T�e��Flm�m6����ekM�cF�iYm�A�ْE[Z����ާ��#-�.7:���m����0�ڴ̴���Ւ��\�k6�յkmR��ZT�-ijm��b�M6�l���lE�31f6���jj�3m���9v��ef��   �}�������:�Zhj�Y���v�wjɻ*%*����4:wf�h���v�A�MC�n��wmPPX��[Yj�-2�Y�)��Z�   <P�� sN(W`9�\� 'V  P�d� ؘ�vr�� �� ������n� (:֟{��+YP��(,��b��  ��:  	갠 =c[� ���^������)�0�� Tz;�� ������t ���y�t ��lE�+6���ѭ��l��  "x4�A���� ס}u�x �7���RB�=w�  �}����}:�_|���@_u�< z�ß}�� Փ�  :/�li�-��lMT�cHZ6��  �<� j9�  ��x�:M�>��� ϻOxz�����@�Pm�=��m{^�=(
z�G���+�K� �=�mM[L��km�TV��  o  ֵ�՞� {ݳ��ց�5�����xw ��� ����a@��N�  r�� �9��@��P�ژ���f�M�[U[o   t�u���ܪ�t ���GKN8�� v�M���u�jܚ�Ы�wK� ��@�E����b�kU5KV��   n� �k��C�����u` �ۨ( �0���l�@(��wZ ���� s�U��b�hV�m�X�mb�M��   ;�����] �� �i��h���Pk����u�h��� ��p�Y� ���Ym����K,ڵ��G�  �  {][� 7Q�  ]ڸ��` �Ӏ���  ]K���@ w� }�  	H$L�)J�d�b`@�2i� j��b���L��� ��d�2E=��*� �    ��4%*��4  �  �=T� �L�O!��z�@��ѦA	)OP$���M2z@��=@ � t���o���Ƹ�q�L[z�t8�1�5�j_[��q7i7I�qY�(�D�KcS��+�E eT?�W�!� TW����{���A��?o�9���QTV��j������
�����$�H��APW�����/�}?���?�dO�P�<`O��<eOS��<ey�\�2�2�'�/�� x0��!� x�0���x�x�L�� x�2���x�2'��� xəC�@�@�<d_�@�<dO	��<`�W�@��<`C��x�0��2�2�2���x�0�/�"x�2��	�x��2����(x�L��	�*��2�/�� x������_�_�@�<aS��<`|f`O�@�<dOS��|`�<e��|`�2�� xɘC���<dOC�T�<es�xȜʞ0���� 0��
x��0��)� 0+2*�0��0 >2*�2>2">2>0��"#� #���
��
!�"	� ���(�x�3*	�(	� !� ��*	� 	� ��)� 	� 	� ���D�S�@DOOPOOAy�_@L�
x¢xȢx�
x�*x�����2�2�9�A��� <d|aD<eQ̂�ʠxȪs)�"��
�� ����(�2�����<eO� ��<e|a|bd�@��<aO__C�1� x�Ȟ0'�)�(x�2'�	�"x�2$�2'���*x��2'�	�"xό�Ȟ0��'�GA�����/���u���X�����䶂��-�	
qe+��j�Yxm ^��=�[���e�[������r�n���D�*V��!����Mۣ��Ie���:T���`�Ek��a�,!��ZՉ���L���S~�U^���wu�5��g��C4�櫶���$[x370=�c�*:�k�kf���ͷ�]Y��PL��J�M�m[�a䖕j�07!�X� u��a��k�U퉠e�A�k:߶=r޻�F�XY���@-�nB`�˙���� y�ks+��!ȵ����`[�`�-�VwL�2�7����e����6͝���Y*=[4q�eަ�nY"�L�7�rՑ3#�%���sփ�t	)�22��gA�6�5/$�pJ�)�����(��Ʀش��t��yX6�`���+a�l��
�ޢ�W&MԻ66h�I�U���
��t�w��f��1
f��ԫ]��8�� V��YGF7T�ٮ�I�T�j�^)�/�G2o����D�{���X0�S��cg&�3B���=��g/�`�w�<�O�trj�[ U�M�����XhYB��6��TB�d2�Q��]��Mح��m"��s3&P1
��J�Xh�S��F3eJ�JXTosp����|�O �Z����a��7DR7L��7��sp�#���ڬt��h��{�=I66���Iq=v��NW<	4;:��t���ԯX�hKa�żV L����M嚺5�da��C��V�R�ة�E�M9.�5)m�	5�Ȉ��5r�ì�Q�yX�J8��L�	v���4�;�!�X�ݴ��7wE`�Ĥw��*!���
Bک�@��?	*��pl؅iQCm�l��B)�U����N�S�[>�]��R��ȃ��I�:�oM�4�d7�B��ap]^j�� Ϟ�(`�V<	���SL*GC��Jb��j�'�:F��u����hU�겱ֈo.�;X2h�E��n���Dl��gb�H�SQMnQv���f�Z�\��`m�����eXb����A���Z�by6�n-Nu��E�꼱`ei��Z�d��u(KA��w����2�إmh�a�p�v��e6�)Y.a�-����Y����������ED�����h������#Eǁ
�/ƙ{��Y�j VE��j�j0�.n�X�Z�؊)l�?�5�Aڌ�"�L��ٵ�W��A��4�]WJ��D�M�u���{��[�[�hE;�&�0e��j�V�b��ͨ��`Ǳ��KEa���+;�A+v���,�$���Mjv�(���z�0T���B��ږ75V��EnЉ�)õ1L`]�2"YN:"�֝��5��M0WV��
�C,Z��;y9
Q��LyM�Щ��/ipVAw��2V�YSj`tث�[������K���sE��;�n@`�m����f�w1asNlI��׭�Ļf$���$&��d5E*� � �UB((�@]�r�
L�C7D�\�B!Dև �Y�U�q]0)M٨G�5��E��p���Cs�nn���nK�u�2�n�u�A9HE�]��ah܆c����4E�v2n��S�՛��WX�PJ�g*����oq��;�S�*Qx(�)[Pխ�*չk1��"�5���h`�V�"�6j���4�!u��1ӭ8�9��Bz�,:��m�U�W��ؙ�3v ���Ci�M#�9k�ʁ���Z��E�N�2]�nv��r��ӡ<ul��4qcf;��nA�3��ՙy>-ʄ<�#I�XV����;��\T����E�nآk0��Oi|Tq��tյ�`�M>�b�5�c�0�8̐L ��*�Y�W���5S7JL��RWA͢���^�j�`!�m�Zv�;u�I��ni���6K�8��o.�9r����T�h�l"���`�\CM��e<��ɵ��ށ�k��a�
P�x�[Y����OЋ+Jh�Dݡ�P��c�l�d�����6���i�0(��"B	U>ţe6���%]�-XNc��,XՁ�V���ͤv��@�h�m\E���nX�Z%bg%�p��Y���L��nX���
n��d�,�0��-�.�46���i�[� *�q�������p;�V撲e����l��@�L+;����Q��(<
���]B�3sC�NVϠkXaJ{��5�c�0d�RE*�pƚ�m��e2si;�,'E��1�n��45�����3�z	��-����ݼE��Wacx�4X�o�Y��Z�hJ�n �C6�虺K�]�.���pRu��R�E���ۘ1h��Ery٫�2S8ݣ�`�j��N;����0����3s-htm1]�9�W��b�zDBL������:�)���4LbMʓiRhYCkb0�m �V��c%#��2� ����>�ٛ Ւ�M�N�]��M��;�H-궆�D�]��.�*W�f���X�J�J�b����M��:4fV
��g�p�8E55�crk2���)m�e���V�l���	2��r2@U�!([ afűf��Wt�x��+cuf�3�ވ�k3�k^��5pPu�-l�sspօ�t%Kt�t�E�V�*�&���%��)gҤC�ZK
�cƠ٥na�\�p�-�)�6�������H4���ՍY߰'W��v�ҿ������v%DF��bS�J�U����;R^�@�sv,Qb�>���
���H� *�P&M�OnQ�s%!0i��F3������͙B9�Rܛ���S��y�x���̓f*ݼ;[{����0n��##���ǒe;�ӯt㩻R8��&�dwV,�44��ee
�3B�n�N����预�]m4$T��or��Mdt������^��˵N!�)�<w��ڬl�DR3��[ɤ^�cY�V�6ti�fۃ-� �6���cJ�3�;h/뉭�ҳab�ލN����Q���L�AԉfY���R����6�<ub�&��L\͗�)޽'3	t �:N�טf�ף.
�,E�e����H��Q�^h�܇=5w���|���lnD�4.a'+umm%��Sy��X�g3A�X6�ڶ��(�!� Q�0(��ulIA��kb����x5j��2*؏h} zy0��<r�M��@ԡ��FLo3/RE�ؒ��o/m�r�S�V��:3*Q7M�&9Y�l=���	WO7fe�њ��jlF�v��(��0P6P.��neV�Y�(��,��R��<ɷY�vNr��4�5�]�Jƌ��F]�� ����� "8������V�F
ܚK	�?7ob�ѫN�@〈$Â��߶��r�ZqV��b��vo#(<VM�������@�d6�;T�@��.лx�g`Ѧ��k�M��Y�m,��7ؗC5i�����۩�\�[v�ZG0#{�r�Fef�OA9��$�`�"�� ��1Lj�:ݬ���N��U�y��cjn

��(պ8�T�3Ӹ e
�.��q�1�O��
��N���`�����j<J5㭒Íc��aE�6���i�-�[̹Ln��~Ƒ�N�Z��5��SP]b#p����2e�fa�crQg"
EX����V6 ��MA[���IV=��ǓE�����~�� �,��Rh�ڗ1i��KZ��u"e�j��$�Z$cE�cE��&d�b�խ�i�4�V7Z��eL�y�[R�[0�@�����Z� �(4=Ba_=Qǥ�߲�U�s�lY
��fY�Sz�L���yfͽ�N�F�U�\�W�a�ӯ�1L�ME@	�d��5ͬ����ݶMK���:�O��K!���JJ��cF:ɡ�U  ��q�ne݀],�VU�x!�X6�yF�XԴ�長�`z�xm�Zo2����"�Z-����@ rXr��X4�^�jC�V+:l/��#�I�$�.�j̿�]�4v]	��sI�cٶ�X��jU73�.dV0��Yl��d�Du�(]�TVct�$U�ud���TC/V�l�F�l�r  i��ks*��)��y"��f���m(�Ö��vB����+T�%\�6�FԽ���>
B���#˷1�YI���B�;�%f�b�6.����޷�:	�RBc���^)��Ml�@�Z��gH&���ˀU�hkv�8���]�̓bU�=�K�j�]�Y�q��ǌDf1�4��f�2�J� 3u�
ұ�uh���ՆS�rS��6��֪��A5�3�Y7�k�s�B�)�#m����M[�r�@�R�n�7c�s1�m�66kʄ�+��R�Kyy�m��w��j*�� �H��S�{sUu�K9qڈ�n2]^�R�z��f���ה�7v��!��7������'0��w�
g�-P�zj:��tHXi�f����I��nfm��^A�
�z)!A;�h�NS�[��(��dNJ@1��=Ź�]J)�ik6����˨KXEf��� ���z54�/�1b�i�s�$mE��:��ܘ��GV���p�本�`�X�Gi��6�w %�8�^�١�Z,���5|�ko��e���8j��V�%�'*3u��g�0|��.����v�b�roǠ�k.����n�B��֮�Q�Vw.����;�s�#6Y��O���-9�ͅ*Z�u��\���[�ݷ�̟`�C*�BE�8���޷�d�����̰ι.]��3�&-Jt7u#�E[���m��J�y�6���� cۙ{��(կ��#*��QXH��p�UF�q`����0f�
�y�+ˬ�q[!��uj%�E1�v�L:��LՋ�vCwB�Q��J**�xv�H+b�L�G[�f�&�=�؎�@��T�oҁ�ced�+	�"�U�w�lH5 �Zi[-�ɚ���5��t�V�����ڳ�Ξy�TK�4m��VGQ���3��m�(!/5��^�q������{Vov��C@X��shkp�*��ct1�t`ڛ���� �<�ӅG2�MŘ䂎E�a�̥nF��[yYR�4�Lʎ�����{.kYlj�&�̭�DX������ �t��Z�P�T�dm�Q[yh�ۦ)��Kj��+cE��^��J"�?A�j��p�ݚ-���5HL�X�n��v��h���t�mXYl|�E&�˦�k2a"n��3	j���>>ӯ6�=R-�S@E+l-Ӥ66�b��#!�T3('R���cnY�J��4\��IctY;�YL]�(�3zi�aۥL�% �˰�8T��Aܨr��0*&�/3p`"��"�ekv%i���1\܂�[շ4��0�E�����6i�5�q� V�
2�f��>M��Z����p6aR	PP*� 0:j�v״0�JD�j�ʆ�%� �MЧ�k����b֕%�%n�k��u�,Rb��ڙq�.d�I���oH�u�:5>�ӣWR:4`�{���)�X�l�I��x^Z��'��fcq)[ &��f<�X7tL�˽7��m��to樲��@S;vCgB!Ib@2E�]5&Pٓd���B��i���C6a�ؚWH�l��Ĵiɵ@��:��e��o[�u�G:7��/���rXYK1����(ig&iFi2ef6Xp���������"��4�qYЍ�F���C4#>8�B�bXN�Z��]�L�R��&�Bkw��Z��o(�[yqᙢcj9��=���&�;�%٦�1{�h��;�:����A�f��XU���±�]�P{��2�4��y��-M� ��mB�/�t����q_aޥ��+f ��Utc�r�)�ٔkjbGNV�a�a���	��t������uc)�=n����b�-��k������++��/`٫๚#���!�]��V����if�	��)��܊�M���8�c�2mKe�u*%K[�.�=�-��U��Wۘ���-ӥ"\����W�(�t��.�F���o.T{�V�F���%��O/4��<�"ȽD]�ޤ��&��o�M��ƻ��+26���nj-d ��5d��v&�L�����X�����?��,:	��ʕ���&7
������l���!�Д�9k4���V���X�m�:/oM���Ʉ[�h��wɷ`ɟ+������{5-�6���W��Y�Ý4f���45�o����]㠙l}�n���5��A#�Z��:2΂�aoi��YX����Vv@˛��ʸ�!U�ED��I�4鼴�
&��{��O�hnޔ�OU��D�X�Ptqb��{�a��vd����u�p���H�:q;�60I�]��6�c�YU��&i�Nf�u��j���V��kB��St��.���1�84�LD^0M(�,м���z�A#5��cB�3v��r�E��2oKD
��z�ce$��8sb©466p�*�	��V�փ�mMq�1�R�����z�,Ǳ�. ��V�Zե���ܳ/b�M�	1j(��/�R����CE2qDbț�7��4%��Ғ�&��-�2�U�v�g�i;�Q e`��ԭ�V��k
�������$C��!P�)��p�k�(�+�QF��x��a{!���&^��·F��aU�@���s;Ɏ�x��Rq��ʥ�� q� �2����!��]���w�!�6�N�b��@��:� i��̴f�X��s%���M���PA��ev�[�s��fĶ�ُ3P�
�0ͱ=C`��!�D"�bל�uh��kT*q<�2�F����0H�o��kș4�;E�sV���[h��ǿlJm��8��,(�H�&�$N-L�8���ę邐��D�5ă�<L�u�	�z0���ctnX׋�+,V3\Y8N��c<*����|V�M�D�.��x~�15|�l�v=���~�9�c�x��/�,~���5��9ڲj�3�U�m�pp����nd.[�&���Cp�H�Ɂ�[�aj����r����콚�V�W�cR�,����%�/���}!�$���uT\�`��,nK�I�����8(��g"�lbN8�Sķ�NwF��[Z�0�2n�RR�^��b�P��у�O���md�f)��A��w��GPEt8IF�(0)���oJ�'Dw��H{!��z�X��E�bY���|�o�΢1hM�VҢ�-�$}��A1T�:ժ����0�����2��\��rě����ҵ�W'{{�r�<Gr⩕\k)
�Э�7TQXB��8��H4����¹�*�)JO��p[ճ���[-8�eN�SU	yKw�_h�x9�#�nAi-X�e���\�=Xt6�U3�a&������Aڼ� Z�ѱk��V|q��IWenk�������bL��Lvnr�����:��qWw;�l졼�gˇ[i�|����p;Y/+E����cQ��]Vgb����=1c��(R�+�*kji{�<;@��y���� ��Ty��D:'N�Y��eW3p7t��ki�u�K5�wIf�����1h����z�4��9.G��wtLK&X��*�$;bѝ�V��y��eUƲk��i&.�-�8^^�����!/��	��UʸIO2�砚=�T]:#]����ɝ�m 4�'{[
�U,�A]`��}���w7\� �e�
�s�wg1�� �-l�t�	T�ɕ���uB���{B�MN��6��/���z��;��O'f�Ec�OlAf���L�/W�V���VW>��I3Xȱ�uȮ�Ze��P\�ýf�Q�~�H�t]�R-�V��j�fuD�5*�tt�J+{��jg9�(!(�P�Ծ���	���;�,0�e��캵l�u�Xզ�DR�"2\�-�t��w�2�hX���G�ri�j\��gMzhvު[[ۊTO��o1�QN�ly�f֨���p��%��r,�	����֍J��Y�%#�qm�F�7�_x3�^͋&�Ͱ�(1A���nS��u8���sx`7�Y�a��poPi7�U�V�4�H���U�Z﫚z�����������Aۇ$�zɣ�i�d��-ݜ%ۤSa�����VjPu6���:X�䘯�lp/1�f!m���U���2��k-�wêv>��߶\�)��h]d���t�_MB��szv@�.�K@T 9�'xmO7+8(��t�����L��z�/���mu��ѽ:+��b>��\��Y���΢��,%;H��ծ@e�Z�c��k8�Oiؕ��1U��؅�|���'PUݶԡY;�������wq� 7�I����dJ警��Bn[OH1��V72h�<�lν�h�o�;����G�oj��7+��c�[�)�����
q�|w�is�Sj�umU.[��r=�X3��ۻ6v���B��A��z^f�U[�o���[d�T�Ĭ/S��5 �*؝���'`S��&P����{i���;EIh��g�-�����z�ض�%o����,6��k%ի77p�m.��W7M�z�j7zIx�D�5���*VN�L��L�W;:��P�|�q��>܍��9�=�b�1�t����a�RR��j��|�'mn�`����r ���մ��<��T}*U��|�����W�v��� {��Zy6� WIW�9_
㖟'�L��ѷoY�YAv����U	��KQ� ��j�6�
^��k*}��MoFe�OqHD����I%��x:���o�u�K���f��L�c�*���{1���Ǳ���3`�ɛ� x����Ck�g",Ǘ�a���MY'����뺹�G)��a3���:;��&�d�7��uǖ���KQ怫�A�6�4+4�鐄N4�jj����:�^ۙz֞Q�n��K[��v���]���"Q3-hb<<DT'o�ҝ(��£+/z�\T���%f"��1R�٭!��^��i�Q|)=.��7q���f_[w���
�m�f����.���͛MCH$�]:���w��#�pLј�l��͒�Q�Q�pҮ�of�!�u]O�l���Ɋ�f�mj꼇��ِ���4.3֛O��NԮ��x���h�^��UG�_�;���ҺĵF�p"^�x�[}{T���(�Z�n!�����
T�3����uf�]�Xӱ�p+:�VvZ�v����؏u:�9|7����XBKˀ��*�>3s9���Z��6v^#{�*�-�z����0Y�fʐD��iv�E�Ov�q%�T�,Í;�������we?VI��.�}[�3
4Ͷ�#�b�G{���x�c�յn�0���R�
E�.^��f1�1	CJ-��ٕ"�E����m,��TKaq*V|��y�}.l'�kN��D��u���9|����`�n��֓=G7ks��Ҝ�5Z��F�|���jdǯCΞ�|cl֕��2,��݉���t"Nm�}JS�`����<�G;I�UiP17�5B��z�vS��/�x��G��W�>4r��q�<���n�ӟlV����XRЮ͂��
9�����ٜ��s6W%���խ*r�0J�>�},؂|S</HH	l��롔��촭���ts��	�4[ֆ;b�/]����T�(7.�ץn�:V��%�9��LbΫ����b��nI�,Хc�q�`%Vk�+���O��v�f���]�[��̫�	�QŖ���ݻ�N֎%�����B똉V���.�Y�su3q��!�C.�RC�+��HF�twi.t�ҧ�g"�»���si���fk�r#�������[�����w��B�~�3�L���[�-]�^`J<ْ��ӛ�45T��"��4%���+x�s�����n��̞�NhK��u��>�X������>��'*�쨇8��b[Bd;�u���M�ш�4Id�hcHwB��frky%!iv��bл-�S+uhr��-�q�\�� �K���Ү�]4�a]��V[ֳM_.�X$�jE��١.��|���N�WbS�U�����:��GP�уF�]\��НZtn��Ú����i&wE���."Ɓ��]�[p']�gU�� Y�٤�CAp�7[C�B�ա��Y�.m�F�im����ubЩ֭⠆mC�\����U��N]6<��w8o��`��Ճ���e�֞��-��kN�:�Ac�(��f���3�:����%���N�je��Ѥ��|��Z�R�b�X"����9r��<|����f�\��'�GvJ��/XZ�y���ܛB,s$!	�Uq�օj��p��ih���P�О�ŋ/+��g? 5y�KV�>�YBf�/^�tC{^I�t�,^<,	�h2;��G+����R;y�}u̢.�a"p,�X'��*Y�)�j�7:֞2���tR����r��^L'�U�7�[�u+ޔ/1+X��sF&71¢W�(r�WZ�0���}b��gc�4���FŷFjΙ����@�`=���+b%n�q �CۓW`��R����Iwe�&L�$���)�)�i�EC=z�T��T�u���n9��͋��B�n`SU)��`�kkDA9&1����h=
خ4k.v[ v�n������LAn���o�}O��5��Q\��S�Pͫ:���4��1Cx�T/	����s�uŻ�����8:4�4 ��(6����"��n<�3)����m��h�{N[��8D��X9+�Y��浠i���6*��M�W� ��,w��[�����h��`�ÞG|HL���_3����m<�QgY�E�m��m�*�#�s�#f˷}��6왴�^@&�3B�1��gk�-�m���Sz�op��H8�d�k�h�i)�yaRund�pE:���Z������������)G��
G)h��m��c��(4ۺz��9{��쾃�AyuVμ��+��Ji���)g.r���6sid�C�H�df��:�M�&��MdIT��X\�# X�.AS|������s�(L�oF3���.�Z3R
���,P�ݽt���!�����:���Ft�u�U�i�T�F��iC���U�|W�`j��/��t�J�pޱԇ�d��T��'�,�.W�$�2f�H\/U�]#�*/2'�Hn��Os6.���u�Ī�T�Z3�.�`Nn���j�t_@��,�7l7�d���8�e-m��΋�ٱ_m�]I�{�L=X1�o�=WZ�Ѡp�[�q�6f��tQ6��)��0^���N�*M���ꛀ�����pn�ym^mȳm��@�1��5�6nk��F��TR7zĔ�Y�jᕇAV�f��'(���I�uܦ�D��Ʀ[Qp0����
ʺ[�4~�M��D��4��J;��ؚ
�3�Uw�'�ϫ�p��X�2�W@����	��)�8�Q}n�P�tir��ޖ����BQ�T��I��uf�V�Q����
��t/�������yyS���3��Q��]-�	��:�i8�Y;^r�H<}]{����a�㱌��O2�� !1�]H�0j�}Il��v��)�E@�a.�=`��-�@���ͮ�4/P���0�+ ��������D�J#+�N'�7�k� �n�^=�%����+�C1vl�#�4[	6m:��P���{��R�8��A��y��ݜ{���
�pD�2Q�ޱ.텥�A�'��j�0FZ��b*�q�
ږ�wT�U��[>�j!��v*�W�I-Ř��f��.�i-0x"s�oRS_0���V�7u����AQ���K\���d��*֡�abg�P�Q��3wN�iQ/0"�s�<f	���Ύ��x��Ե��S�&�}������ApU�[�B}69��+�i�ئx���ۖ^]Ӱ3zS��/4H�t��M��rgNٶ\�=g5�����t*��x���h'v^3��;�V�R����s��0��|�n�dy9�`�J��l�9�՚�I(Ќ��*�GB��cUeY�[e��aUS���	�+Z��)�57�2�o2ul���dF5z�;�\���n๠3Y��c�7�$��6^�5k�l���V)��J{�:e���QB&��o�n����n�GV��1�tu����!ER� ���$a���|x"�!W[����w�1t��SЖ�2�`���ݻ{�:����'fb�
k�t�۷7����Ç�˘�|X�r�M]ĵ����,�c�U����@�|jF)8�Z�ң�=�BT56}�1[�I4>�FV�㒠�[+�F�Z�]lS<�{�7r[D�O	J��Z�r^��P����Gtc"=S�U.Pe����Գm��e8)�]����X���"��1�TLr#&�1U�[ԝ<��RJ��[Ƨgɛ�#V8s��Ys%�t���g����.�-���J粕�Ⳙ�n������)����T7��6�l�\r�e*5��U#t�'#k3ܡ�[��K쵩�ۛYCQ�oo�
R��z�vs[�_-n���Mt���k����Y��}�\-�Q�j�Li:�iJ��2�D������8�Z����w�W��ʕ|�����ܵd���v��Q�T��dN}��9�V�P���m��˦��J7T|\�H�iNU��W�C�����D+���(p��t��7�㥻��)g�:��+gu�94��1��g7FC.�vL�n��-��Qopp�����Yvf:+�C��β̺׷��ѹ�ѭ�[���E�<��5]�-�+x:���Ѿhͧ2X�X��7�
'[[Wܴ����˪�l-K�E�ܬ�wyl<=��$��**��&9*�f�����|�F~�Ԗw�?���ÆF�ꛀ�9y�äJ ������CWL^&{�<�?�b���l�1ݓ��
غT6Q@��eA���geЦO�b�M����m�6Ub1����x��k��AI%g1�>3fQ��)���|;� 7:-��&��2N���Q��2��:��;0%˗v�����2��j˹v���nZ�\��yv�}~��g������}�j]��"�+
�T�E���
�1�Ü�[:�Eְ]T�mdU��7Db9�eΣ�b��A�YJdL�Twk��t��ؙ,�{�\�{���4+ny�y��1j��:���o�⣲U��-�=N���m���n�mTlkɄaڊ+��[eS�BvH�oe2�4d�	���B��-�#��o�|��GT��C��jT8�Xk\��n��a��w���%�sԖ�q��m�1�n����k�H8��Y&��+%#Ҁ\�l��t�������57�Vk��B��9��_ 
|�e�������}}���Ӥ9�]���	�5ou��@Y�ɛ��֫�&?{�r�W��q�Lo��o[؛����,���˯p��8d|�f�;�h��Ul���:$�=/h�9M��%d<�7��[n�K�C�t���J��ٙ@
�/1���u����|�_]��Ӷ�ɯ3���}��V��v��lA�#i�Z&mi�7�n�oT3`9��8*�lp�$�K0�Bl5�;�[�-�":�8�&e�BS�ut؜P�n��b�/��%��;h�*�|�K�͚�����z�w����j-��Í���.��|(����t�\���aMX��x�a��(!�n�:e��@��
#A��ڢ
I��Z.ݜ��,?5�|�b��^n�/����8�Q�T��$@��i�d�j�� Q���lp6j)4k�Tn�\����s����w�^A����c$E�����yy�|��<�:�ZիY�Z��kpZ֬��(�����v=�DQP	�]5���٥O������}���ǐwuZ�ݽ�l_�מtV3b���g���/(%����Y���wهeB(2>�
�[y�X�Y���ᖃ�����VF B�L=�M�:���jkUm'�#��P�[W�Q�)hѪ��5�nⳢ����,Hu@r��	̦5I��[ĉ��@*���.aY
�xq�NR��bA ���9�d|�r�#ǳk��Z�kZ�"�v9j�D��C&�ssR�̰��b�+J�3y"�8J*����n���1��HR�֊�K$h�ڸ��)U�+#4sV��wY�?��ݰ�"�A/z��r�N�����d���k��F��3����h��;Q��\�݂���7��e�N���P�,WL���"���nr�W�*�L"r���ݳ/m�� ��>�Sͤ++IҽK�]��<�';g�6�%>�4q�F�wz���\E^�%"�����µ�B:��kNa��f�(.*��'��:XHC�\+��	:����(YT��x��(�8Q�ӎa���J��-X�t(�O�մ��5/�cF��f�u��a�%Im�n�9���Ģ��j� /^�݌�&�sV�k��ۆ>��-$|�ČICsCE�׎Π��x+�Gp���G!����0��D��Q��2��)4=���oGev��Iʵg�{M��o�6�9�u�(۴,A`p��K��s-�*�ϥ�١�αl�����/Mܹp��wLc1�c�1��1�c��1��6c��c�1�1�c�1�wW�@��㢕�5L�|��N��X�u�%
�t�L�D���O]����uN�Nw7�,gkO�&�f��2�Em���_Iw1���Yئ
}�_>Va3Vf�����ٺ�R�M&�.��:���ZK5����tʑ�9�%[Z�1�7��	w�����G���Q���
�a���oFe�h�[LإnW���0�i^KS�-60��:lZ8˻��Е�A��Y� m��@�/U�O5��ӕ��;i��W��r>���OB��T��ܘ�ܥk�|k'c�}�cH����K��|��1�����UdE�ٙ�Oos{�L��3a�f�Eֳ.����>��5�%,C����p��ʶ�Zn��m�9��s!n.ove�\���Sk&��/��b��n+2A�U��簕�e7÷�l!���b��b�h�8�F5�� &�Z�����
sٖS��zp̎��}�r�p�����=��Up*�0�����X�V��������N!kf�,��� �BVfE2�^��v�����9E�4i")Z
�󯞚��: ���>�
Ů�څ�/m��7T҂�Ar���.l�66+e�*S*�f�77aY6�z�=�B�AuWu�D��a+q2�a���F���Z��}(2�V����7��Am�ŗ��d����XhT��X0�����W�1Y��\4���n]���U�/�3���Lq�e��1���LcLc�1��Ƙ�1�l�;`�1�fΘ�1��1�X�6cǾ����;��y���V�tW_#�q�d��Q���^�ih;Jk�{��]1�U�E�O	��YwWb��:�Ff]�&P��;1��Y�Gv��s�ۀ�"����Q�� -�fR[�o@@�7����!����K�핆���< �z�^��R��)�������/@U�)�Pi��_���U\ļ�y`[*���bc
�Y|�.���\y�]2;��`żbZ�u��)Գ��!�h�
V�U��Y��l͚�֊���g�+m���B�	<J��;ee C7i�T}O��R�	�\���J���_ۄ"s���h�]}�^�!`dӗl���[2�.p�8vV,�`;��_*-�;��P�����&�,&���h�TwD[��y�����������ú���,me�.gkנ2��6�o̸P��3���يH�{t��|�ݖ2���6�2�-˾���̌0�5�1��m
P�M��܀Xx��I�3�.	���7�>�a�;�g)y%�<Nŗ���0/���_5d���Ύ
��]q���8FL/B�HĔJ�M4��4ט�2V]K���\�4R��Y6RlD�R�ц�{C��y�S��9��--#yeo+T�99��Ѻ�e�����)�ɹ5����4����3�ntӍ�>�3t1���V��:v�I:9Z��۔��ұ<;��VU/��ÇLc�9c�8c�9c��c�<1�1��ݻf1�c��1��1�X�1�[w�j���]��#-�'���f�j�om"x�W�3�u�(]��A]�VΕ|���.[oB[�Aam�
�ճ:Q�&A�}����S�e������
����Ӆ��xֳ[�]�lx�e��}�[�,RKOq��W�y#��A"�͒e��BZޕ���du��6Z���gvH)ýu�\h��X�U�UʱYv��t����uqb;���_fÝ������C��]rV�w��v�,
�.�Y	����M�Y��;��|��M�K���m��aR�&�f.UdC3��WLC�u+D�в7{,ꨩ��1;Lm�F��u�,Q���Ѓ�P�޼�A�ٹa�Z�k�ޜW���&T=�6*����Z��򂮣Lf��}k�]�4Y3a"N����<Q�f��8��7-|��ÇL���^μ#��̭�uoV�L,�՝���
,gK�9K��{α�T8h���ôn^�!�
��]��3����������G+�\&�ֲ-�0��,�\3H�i^�Ap�B��Yܬ����ňDr�m���ߪ��ƭL��NӀ��&n�������B;�^0��[n�b��$p�ŭ�X��n�F��Y�u����٠�X:e�M�uX��n��I�=r̰gw���w��=�F�/'6[�i`)Z�{��l ����g���VN������Cӆ���}�/��:v��c�1�cv1�c��c�1�nݻvc�1�vƘ�1�c1������[z'V�o�q���V�V[h�Mlt`YMmz��2X˲a���Ff�Z���FydѴ��p;�UN��I��	��[� zc��V#b��Ӂ�/�s��{K_8�^�Tp5�A�u6��W�f:�����X��AC�4�7R^uV���Mޑ��R5/�wgA����o[2L#M�$�R�9`U���[�BԮ�ޙau'�>�΍�D�LGSB�r��$:;[X��d�e9`�ǔ�����[n��t����,��B1���RQb�Ȫ=<�uV�Y�T9X�Q��yD��YDN;��,�O6ɇr ��U���hD�͠���pV2�
�W4]�\S�L�1q�؂Ȋ|8�>�F������_<�\JagEs&�U`7pue��ɻB��V��;=c���Ϧ,�Ϯ�9�;A�k�N�D�5>�؍-�ȍƃD4�=���p���jv��$�����|�CSQ22 �9�,|�YzG1;�Uy�H��G��O��O۷������83!7H�kN��:a���n�x]_mIuG�w_>0��P���[��LdVY���`؆t����]�jv��n���!��s��*�.-���iI�� b��Re�/n�oJ��Il�c:@y��gU�<��w�@�}A�=����Qw���l���ʵ��@�� �Q����'fֵ�nUu�urV�7�x�!2�U���t� tUI���I6�������4/ �[����ymM)of0����j�E֡�ZX���"sp�p�L��s��B�w(���n1>��k↭�+���凘�)7 ��!��*��4B�h�1�� �*����[X%�^�Ƕ1-w�Lix�ZۓMZ����� �Hڷي��TlZp��W<��u�XL`^�[�B��ٹ�f�KetdR���g�>�Ln4�PZ�r��-V��ymR�ٗ�d׷]ZX%�N�'3���oA���7&�F������%u���
�<�0�ϡ��j�>J>�moV>�H��ZL7����Š�T#|Q��U��1�\Y�P���;�sQI^��7*.�D7+b��nh����=��*%lx�ԛ�JQ ��e�BY��1[u�����,��q� ��P�Ç�)U��qڝT��٥P8���RdG���
n�z.����1��P�l�m�6+��.��1�����m����e�CG�n��M��2w_0@Vu�S	���]ӞGҩ��&8��]�u�w$i�R���.Cj�L���,�wM&��8�uJ�$*���D���{�brO�M��|��$��Y��LEX��Y���
,育Y�ܶ*]�{Ws9�&�hfG�MPx6i�b3[B`1�zGQσ�LAۏ�mM)ݮ���h�;>�:n���O�X�Æ,���mt��*��є�Ttq+8�C�Wn,�vc����znT�g^	�6�sw;��)4�����T��q;=ڇ��[=��p�h���Ay/V:v����e˄��;`��(�l�b�6>�dV2���v��[}X�=x��a����o�%�{���O�H\���%�И���ug��j+{�1�صOS�y���\��+�(p��@[m�X��k���/��])(� ܕ��d%����o�Ci��B�"d���e<Rf�����k/��X}A��$��waZ�}�SC=٭��`��1Ihp.V�Z)/�9N��f�Z��0�i��w�B�eI��}\1��5Fu�Y���ۉP�4G���J��ԙK3�q��a��{u��e2V�;�/S������Mە,�*�/�<$`\�vq��{[7b�4H�r���	1W�U�*`�ԻO�ݺ��
㋄�k*��㕪�]�u h�a&�oV��S������v�̯����cB��]7:m�nG!�3^����d�68!�1�>�K��.m�޽燻r�Um�v耕Eiح$Dkq���ðv}��/�g�t�b��J�b�����%N��{Hp��g��u��Sk�Zu�ڲrKl��\tɱ��-'��r����
�j�0̎eG"�78��x�taʆ��ZGE[��]�4$ �;x��r�K���}	<F6�)���s�!�R�P�6�2����0��<Ok�д�J�� �4��:��)=�v`J�#�w�y�7&e��[�0���R+ң�Y��y��Qi+2�%<d�/���$s�خ��nC&\����.Sq��+�&�])�3� 1�f��P�9]Z��q<����A6��1��mèsB��&�A�&9:�/��z,�0�1>��ieA�,�9�p�I[
�K��k6�Ɨ�h?(��պ�;BYI����aR�(M����ի(�7Z�O��rA�f�pdN��^��������
�+���U�mu�ɌY�X�!�0�R�e�NH�bޘ9�!�7}��o[�����9�
��k��R�s��5��b� T��D iI����/��*�ަ:��A��k���m_K�Y�r������4;-�'���ܝ`�q{fH��������L�ك1��:\D�U���aa�{wΛn�e�rI۫4�4m�x���{�@d:�ZYэ�7q�L���r��P��	N�Ăֺ�Z)
%��'vs�E��(��у�d�z�XU7{7���*�RNP����k�5�����&^��*�>=��`/4 �,�Z�0(�4 �2h�EoB5���W|z-��
]3{Q����µ����`I�<s�:xm,�v[OWP<wt��Vv�b�tP� �&���2��M�����7"%�*v�={��6*�Ǐb��l-��1Z�{5|�3wR�X9��`�`2>�
�4�3������/
��w2��t��X�����wa9�+��4���r���i��¨M��}�+6��̧�Ʋ�%�1�Rw�Q��iw�^V�mk��d5:PNuH��4h��p�!�Lժ��A0�u]x�L�!�/Z:�:Ԇ�aˬ�Y�yt�`�vM�ӛ'0�'�ۄJ�o�i�!cM�!�8ӱq�{.r����nNd<��R��r<�r�k�������X2�+nq��R˗H�΃Cr��l��F,��&Vn�r�x&p\�1$^XbB)h�ԫC]h�N���[��v���Om��Tq��&5��ɵ_KsQT�����;:�<�#�ѝ�c�P	�˭ぐӕ�J�+d@K���U�1W=]�M��յ1KoH��(���ǹ���x����������a��@��8�"Z�\nƚmX�sq�unP3�t���� �4e.n�%1�LK�.},�)�2�
��V(��d0�wj�"��o�[�ݾ��5�h�h,�gqk�=Յ����v0(\T��1�3ɏ~ohK��/;�n�}:�D��;h	`vJhJ)N�Vq�irc���W<͋���8^����W\w@����UӖb��\Ĺ%�*WK��}�g}E��!�nPw˞�b��xk�9�8��3*�s��1Y��5o���h�N�n�a�w�2w*\̫3p�`�z堹ǨQtI�u`�v���pA
J�ҍ���z5��~<���̌�;��"��Y,Z���;�����bԖ� �ée1ҷ!��4����_X}�N�oO���nT)��.�P�
�F)��_X%�^�Y��`��3+�w0�X�s��ύήΒ�Erqڅ@o5�:Ƒ�󽓡�yï]rW�T�,�W�qI���F��0�#Ph�t;x)��_:u�>�l����a�� ��R��0Z�y��f�kiU�Hf���g	`���K�G�Y����S3���Nu��u�Ф�`��]O���CX��7Q�	�kY�}m�;*c�؆R����qa�-�G�H��-�l�*�W-`�R\T�pɣ[3���aX�=eSw>M�2�0N@z������6��0i�N�VMŪ\��r&���µqZ�٦��i������Qp��Lr��{�Y����,]�cf�z��9�8�p��RH#ٷa�O!�j�	/y���L)U�7`6�V�\�& ,ƹ1Qo#�Cu�\s��n�hjJ0��۸u/���"*��X�o��&�M�J�pw[ԏ�~C�;���7z��޸ݭ$�u�}���QTW�*��_����~�zJx�����x�z��U�U��tM20K�AM4��� �Il:`0W���"���M�[{رF/��-X�ss7:gY�smkoek�'To͖jV�U�jU��`�{ԝ��j�����p9��v�b@:�Zfe��T����Q��ޕm�Ó��<{U�KY���"sz��G�ne��!�g�,$]IB+(�-:��3\�2Uݞ;��w1��64�ǽ��_rpl��0^�]�UdS8��u5�^�.�4��bC��K..�mw*�K�Z�M�;Z�V��K�Vw����pk ؽ�8x���q��H���p����sh��|�Ja9��ꏮ�O��C���}�	j�D���	]��r	�D]4���f��.�ҽ��1���ko@+1^���y_և��H>���z�������6�T Pm�w5�4z�h1���s&�Q����U�<��*��0*PO�^�h��Y��/�0E�6'7%5�rj�u��FgmL]�V�J]��==ݹ2�,k�`�S�Й|"L0w�q�̨8c� �2彴L�&'���"ɽ��ؾ��X2��e�����qR�7�̨�����Ӟ��)*'m�Y�wh�_9����4����5).f�{2gwa�vҝqU����n�U�\$�7�|^�m�ڭ�j�:���t�^h{���m���c�-�A3;��ӏ\�1vt2���ih9���F2&ꕤM5�Gҟ:ݼ�[���0�}9#��8�:��Rgh�u}Yb���B�e�j�h�H �f�F�a��1�2��4IME(�Ƙa�A�	4�c��h&��h���	M"h�H��A�&�%�R��h"�R_:H 	dSF��*4G��|��P�u�i(5��Z��!v�تK�`�����;a�Q3Q�gm$����8��������ޒkmk@i-cF�5Al陊&�CF���AQS�vl�Ѷ�w:�'>������(-��cX���::B����t��:h��RU�DE��vk�}}}}}OB�Ζ�ڻ`(��%!v5ƶɧGA�,�w]Z
)��m�^�g>�������66���5�릨(h��"M�1j�C�]cM�b��n
��ErE%4�1kN����lWOl�
��qDm�v���EZ�4�ڛ�\Qݠ赊퀪:��v�Kf�vˢ&b�������۶��ã�P���=h��TM:��wd��=ݎ*m��:-��K�+�����u�.!�F��]�]Vb�۶H��D�5BF�]�\LD�b�JJ4��GTD�5�����m�:-�)f��"�4��:�Ѧ!��gF����]���T]c��m-�E1|��oX�I.�ݝX�䯎��;�8���9Lᔕ!�B�0̝�Z}j�i9kE�l,��+�r�bf�[DT쏷j��5�>Yik�N��PU�W-LH��������Yت��V@�p��ۖ�j���7h�ؠ���㓟A���H���*��!:�x��${L�}��Y��	�ͯ���ot7���5�;�]���٧/�B�f$��R��n�#��'�\��-��}��m|A>�3�	��=�w~8�?L�[��ߦ��n�UF����V�+z�ls��{A���6dt�c�>�ߩcϫt�	u�}�\����EfmU��a�^W��pLN�ig��y3�:�>힖�%�[h��$�}r5����Ѧ���2ݷ�v��6v$WQ��� �>�0��cd�7��.<�y�����|g��b"�=.�o�7�b����h�JU��aķgf��8=�^7���@l�,M�����I�~h{p'Źȳ��2r�Y|�?�a����sXޟk��;�_;o�W^�ƻɓ@��Ru�`�3��$^�OƧ��Ѣ�pw�;:�_Q��.BZl+z��:�e %���,�<<�mK�1���y�
vX&�����T�8.(�UDX�Z2�oI.���k��Њu�q{YI�zE��7u:+P衳{J�Q�
��٪^�_G����s��,�=/�(1(�=,]
�6
ƿFz��wA�.���s�+��e[Ճ�y��D2`z*X���C����o���<�Ǜ{�pVf����i	�W�����AbFb�#���u�z�K�5��ޙ�f���.����1xy�K��=��������J5���FZ2Ŷ�$W����p�Y�ɢ���6���w^� ɻ�'��(��dq�c�=��B�Fuט�������Wc7�����&I����G�^f��;�s��k�]K/�Ϝp%T�����Z3��~��������Xrk݄��ހ�ۭ/��d��{�+�mbu�\�_�a�A[��'�些��ꔼ=*�lͪ�rtc��zz{)b��:�׼����
>��i��b�͚�0B/X�h6I6<�#_��sn{��������y�F���1oI�D5��n^�.��u�-�Ǧ�à�xk;��7z=]�g;#��UVH��#U��B��(B���n=�V��ꦌٓ�34�2�y���n���L�|1�����6�:���#��p!�+�2��^�nS}&8�Ԥނ�����# V5����gc��m��l>xF�J����[�73�dJfU_���b�V����ŏ���z^}��|'���yZ��YS{cΪ�m�:���A���9��?o�2g�N�
{��?]��ƈ9��]�ĉ�>X>�j,w>�T~��>_�/Lx���7$o��݆�+:���8�\��o_��m'	�"��c{$[�M��:0zXWP��E,#k=:�k�=:b�Ӽ>�Y"��������(�}%���4T�b�<v�!&��ط�����|m�o����:v"�\���%�;)�����y�`=M�O7��u.���~�o��-����ݰ${�^����|��8��y�>�=���b �����8n�p��i�{�}8��S2�V6�a�4��o;4y�՜���_��Į�Y^�BD��3�_z���Y�)��ZƋkLŔ��q������(�x����[F�9�n9�q혂�L�%6�/kx[7�x�:��؛�4��C��.�+��m�v#��"�69�.�elrA����{.<�:�m�nJ�.�T��e�ߩ[R�GpLu�i�dQ����W74�B� �h��.���n�&yQ'������~��ޒhY�&:0�\��s5l�; ��}��թg6Η9�o�{y�� ��.�>���	����C�	�z��3��o���3Ӗ��έ���N���8h�-�c�)��I_�=��_�����7^��9<����B˽�
Zl.><�\��~�)|�'�u��=���!��j����\{��t�dXç���`l�l�Ϯw�[��1�÷�|t^�Cr�7\b��I�r�'m�^C��N����Jb����GE���ٞʒO��~I�;�$������C�e�[I���#N;G0k�5'�����t77���}�;��#���'���w�I�}7ϗn�r�s�ԟ`��g�^���i�6OzW����1}�uUv���ܞ�f����L�^���`0գ��d������g�7�<�n���שxJ/�M��Rȴ�D.ݒ��ǜ� �%�%�*�s����d�B$B�Mrq+U�<��(��7��v��3�]�6Q/7���G��`�5/wgQTpd �T6m�y#�Y�B� Q��t~b�t���������
)�vռ�$�Z���Q�*wv{ڡw}X*����tG��x6�6cl;��"��6�mN�.{��v�m)좵��^��f�C}����
�p�~-�ɠ"j��g���tq�������i2�f7��N�`�~= ��=�ޟ`x�:E[����yڪFA����Hm��1=9Qqs�r�aA���{Z}�t�����K��<��l����Ѝ��b��(�Nv��g���c���q�+���!�9V�G�*!�C�]�=�A8�6�=C�	�_9tƽ���-f[�*�28Iifw�{����ll��p��8k����I��vZ�a�V�Eyx�j�9s>�|Xl�eͷ������b��<���X�vA����W��g��'��ɟY����^� ����f}�Q�벫of�B��s0�݈��ܣW�,�sU4�$O�S^<����M��V�ѱlȺ�GW6�$T��e�_Xr�7t��N�!8fH&C�]áTq��C������z������':p�j��j���F�>�����F��x��n�5��ޕ���&yzzL�箁�/����Q�����l���d�G��<=3�[�OK��n]���w2����+̢��q�|�x�fHʆ���pl�Ni�{�=�V���� u��O\�C���^�X��>��ͪg�a�z�b義�I^y��뼯�N]9D����Ρ�ͬ��`��}G�%=�/���J��A7�}k~�=�~������S�3�)�.�C&=/�t|"4�β����:�����P��~��A,%�$T��!���z�	wIU�]/�=)[����QxA�������ve��m�Y.,�$�@�x��=,�bV�E�P�c���r�R�����/7�z�����E��v�=誸 �捯y��A����>�����; =F�l�Ǳ�����ףx�z�7�<�kU�5���%s=�g�j�op�=������m�ř�\J+OjA] ����}r��2�iӟJ	����Ķ�Zshmu�Vr�-��֠��Q���v�����޺B��f��X2��FuӀ:9�9�����|��#7�^�L�<��}�z���Qg��F{Ew�t�g�	^��xf�}���LK���'3�����p�ڹ�{R�mbu�냏�=���\_�;t6ҳ��P-h2��7飸y������v�׫�ym�+��u+���L^�q|��z��v3��=��k�a<��C���y3���@�M�NdO�:Iط���c��q,_�9dE�͓B���}�v(���2b��x��R�/9����{�2R���P���	�����~{�z^�<M��̩�T���;�x�>���1t�>	����MO/�3��j�s{��a�qu�s�L�z�����ў#�c�P\��(/F��:�kg����2��N��rx�˛���5|Y^hv)�����=4>#�O^���L�2�q1�H�_f���=27�nGtoh��u�o��F��!�D�_y�Qf�R$j[���L5U�ݾ,�d��wC���G��V�y�W�p���JE���Y'Ff�����NL3�u������WOJm���M��j��Fv�>&����1c����C���AXF輭yN��1H�:��*'�J��v��t�K�:o蹗.�Ϥ�D6�
}.j(�`j�<"�l��D Ho�����-����) ����;~.���w��}X�_`K��!��|��D�n������Hɞ�'�:�$��1gc&���j��̢'P��ez##���#�֡�݂�!X��� ��d
1��m���E�?P�A��E�*of�/z���O��=�{7���A=g��h�L��ؗ7V�т˜7}^k���7�у�>�9u1a�yO��{�	�z�<j��Q�{ţxdd�Y���H�Fǃ#,hX[S�3��g��Oo���3���R�w�4�&k�>�t�xWi���;A����]�\�d�kcr{2n^'�xz�J������c�N���i���ߞ�L�^\_q��%
:�1�o|�vK\�v$"� LQ�u������h=X_^_��C�^�o�G�sl.�NO{8��`����i1����G�k��&���G(���XW�uϫVB�H��.��r(�u�qS����*i�u��>��OvI�K�kl%�;�.n�Ӥ�8uح^ӯ����g�'�	����+�����-t�uy<���4��I����O��O��s�>���y_ܽ�.�C�� O��z����{�˼�� ��F����57�}��
��D��|�9-����m�ϒ��\Mp�3�H���K�g֪,����H+�9�;!R�Z~����nί�+��"PC�(�{}^�����09pz���v��RY�r�xRھ�vm��>{^�6+����:ǣ�n�|6ac�h���Q^Z�m���ʭo������1�|�L��p�c�e��y��b�����O3<��]��(���O��'��= ��<�;�8In���{|�V���=��Lxx������y�-x{=ݓ}���6c"ã|'�W��tԔc5���w"=}dף#F�5�x���Fv��4��#g�߮�>@���Fֶu�rw����"
 w��!�]����WiH�ó�r=�!�Z��<��ڴu��˄ ,vor޴-��Ȱ9E�.�.��Me�6 �b;v�&� UL�0�{�HE �5���wtݝQƌszU0�����c6��m���� m�O�O����x$ʮ��������y��ȋᘭ�#�����8��B	�et�=X�g�lj����S��~�x�����U9�ǁ�ϤC�~n��X�uma?x5�X���xK�:[�x�kɑg�dv�Kp�_�x�|�d��n������͸��������z:z��;ٞnzL���@�����Ԇع�<���P�H3��#%��I�"��OKϷ��߳����Ƹ2�O��髽!9cF�e}C��.���FN=F����NW�MF��*�ds����=�=��6�o���F,�`�.�����J�mQ����9yC6��O�{���oZ&M,}|Ģ���mt������K_C�ǏϹ!�s|j	�߫���.�C&=-�C��������G��cA�����65��u��B��������b�!�����|���HV(-ˮ���=�����0��ޙY���j���Z�K{ô�NtF�<ۣf��!Pft�7k91�S�6]�T�Vz�U�ȓ��q���p�9#A���L�*h7���b̍�� 
t��O�w�N����LW����Z�Q�!G��b
���hlۇ:<v�8�Yy37jV�t��9yp��c�X�d�i^"���t�~��n`\�2jX�r����n�c���	�G��޶�wk�9���;aw1{m�ux�]`��ɚɲ�k��1�1��G�Ҵi��ڮ��PK��q��[����l�A����d���n��x���z��7��`ꠝ�6N	n�u�A�Ҥ��"����Pp[���`�p<Q�ep=���v�K[{�$�#z��v���Zst�������*Q-hRyT�j�����Db��n�r�L�h����)d#Z�W��]��̈���6TV��E�<���k��Z��}������[K���
��gyҤ��y�u�PIt����ǜ�m��'p�] :�h0�F�K������t��"�����t ��eE�u���i���֙@��u"C��5yo�SM��V�R]iZ雍5H�o!��e�]�M�pԾ���ۼ�P��^��BStv뢾�r�(�RL�}z��o��%��.���+�`ۄ���!6��y�+�a�jn�q$U�T�vun��cو�V(��\*�*�����7�t���|���r媊����m�]a���Y�C��%{�nH�U�8�SԎ]u{�͊�=yKsU�!��Rl�+����Cx�h��>YAm;��9V%7�ɰ0[ʭ����1eɐ�ij]1�W6�fs�X&-˃Ly�`�5�9�9].(,\��3iV��H=�'f�6�g(�-��{� -#�p�\�����2�������b���̺�[�4�њ6r��\�]nn
�tm��-j�b��^�[cY��V�'ZB6m@+�eqk-n�8����wҊ��L�}��ʮ܇�6Sq�{;�l�y���wumLkd"�Bب��E��;���-ϔ5�j��)b���rQK��4�-�컠2��El��'�5���Ėp;/�͸.�9�^�Ν䲦����s��|]��k*�F��^�r�n4s��q;���5�]nV��\rR���y���_v=u(�[���Mk�SV���˕+U�;�HK�Q��V�b5]��s�����^Y{]�7�ŷ�m�7����f٩5�k��	w��,2� ��ir�����kk�b���\���޽(%�a�.�e��oJ<��l��X^�&$���u^��7/wD�Km�o��|� ��|ʘ4����d2�k6�n˝X۝f�_V�"��qjo���+ی�p�,qݷe�n1/u�Z�s�q�JsN=���\�����?_��%�Z�Uk]le֍m�
(�j�������j���";�vz�N�֊O���>��.=娊�� ���-olABRQ��n��AѨ�IED�뒨�ю�s�������lFؘ����j�l`�G��#1Dy[V�Dt��m���i�}~___`���:||��"t4b����֎����b���3y�n٣^N��c�cmLu���������>��v���:����c����wn�w]�v�� ��OcDwf�ݠ��kF��"ɋ���y㷞y������WU٨��ݱ��n�b��p^F/#W���"���]�Xݸ���;k���2�-��F���mw�����{��y�+yƫq���\��Sյu��m�G�.�碶:�Wm5U�U��������LQ���Z��y�Tǝ�Ѵq1Z�Ku��lfv���v駘�7s�熈ӯ<�݃���7o<;��-�]��#��ō�j��b8�ל�xy�W%1Q��������;kG]���ݒ�*n���]]�n"�4Ĕ�U�6����<�ɧU��n��5������w@�{�A׻*�z�	˷�>�&�9f0������{�1�Gݲ�Q���BU�c��tʇ��Z4�'���~�� ��y�۶j����N�2�M�v#L�8#Iꆟ�o�}o@Ց9�]TϺV����z	 ��)=_�����r_#ޓ3�ul�4W��H���PB���p�/&Ӟa{q�e����~��[���*yg��1��.[d���&��Ϲm�u&
ٷ�A�{rq�g~�萝�]:��eU�Ƃ6���&�U��ιS �P�g�C���ʬ`���zcx�MJBö��+���1����\�$$�Ъ��yޙ��^��Ϡp W�>�u񢮢'�$<��n���N��M�ؚ:y[/:�5�/��H�2���m6g�;Z��l��H��x�%D�f�8źa�T��ٓ�kxDq�_4�$Z����9w��%�Ml�Q͡�.WG��Zd�$�:�s;�4Af�QjY�L �#�]��Iw�e'��NP�x-�a�K�};];�'��%��-�6!^j����� �ۢc�l��5��K��M��!��~Zy^MX�l!X��#�1Y����;2 �nXf�H`?K�
C��r9ó�ױ��Mל���a���3��/���j����l�]��h�S�^�Z̖���B�O��L��y���{;9��J�V�mJE�O�6��[S�j�X(ge1���ޗ�~{�5��{�B�x3Y(��$lS��˿�;m��j9��&�[�:!a��v�/��)54�g�|�ݾ�zz��m�G5C�9.Z�ƠK�@���@Ccü�������
�VjE1��{�j��V����d�ƞ��}`	0i�񫺥�h+��P�)��p���C�WS��������^dŊ���N�d��gu,�0���X�Ǥz���sQ}�����:0�����kR�1����U��wo
�lc��_�4#�$��df�qg���b���r��w��k���`�x�9��v�gB�S;E��H���oӲ5���A���H�f��v-�c�� o���]�K6n�V�y��<�飔��
�b��5������}��%��������ב�&_-̋Gd⦔?v�A�P�o��~�L��eySt�S�ˤ���Rq|�n�����p�������h��]���0C&�%����Q�g�ٶU�l��sӼz���m�ȇ���0~O� ��)v^䴙�9ӐC�hA�u+�!>��� ��@�4
��z9�m���{�6�@A@��IX�K,�^����Sp:\rbK����}���2���F�+UE�5*�i�m�e�G����u}]b㼽�PkC�@��.����֌9�m��g:�82L�Bk:�.�jwc��Gs~�����"9���ś���ѥ;�7i���Pܖ�tB��`���<�S��o�Dӑ�z�5�F�}cfA�;!w��ޝĬ%�~�~o�#ؤv�|�x��MNOb:k��Dsz2:Y�K�{r]�vAnm~�ɼ���u��U��ơ,�g�*�*:�l��n�6�}Ы��p1�C�L9��ۃ`��v��J�,�x	�N�zY�ӓx[q�Ok:T�7-&��GM��|���չb�B9�s�e EL9�C,Ɲ���wL=m�4B|(�	��[�It���摊V|��,�F �_߁��>!�9��Y���&�Lf�:��_�xaG�0�%s�P�r�͔ޒƑڈ�N���x��O �TC[R�������NS�7!�4�*)9�YB͇2u�߸�,(Q�nc7J�����\�����Z���Urj����q�
篍��	ړ�-0 ���G6�j�i�,q�ǥk߁PK�X��B��q�m�[,|W�O;�r��ˆy�����;.�kݷ�,9�JT��H��a�u��1C���nsg��ԑs!�*b�zs���Lw�8�	� <F���r]�IՁ�,�8{�e�����.�.�ή�����v��30�I�Ƽ:����.���3�0��yO�j1�Cr1�L����F��m�Z���g6�Ր�׽P��ޔf�+�#���=RW���j���y�ir)EZ-
w�n����'9T�F-�ԫ�ș��L<�qt��ӝ�e� e���?�)�m�}ݗ��������tx�dqf�0V`�x#��2G�A�ʽ�6�C��d!]��S���nk��*/����f�s�ME��e�#s ��45fA�����4���MC�.WE3���d����Ż3����C�p�q%�j1�X��ln�c�;  �eȓ��q>���1������/8��i�r��L�4A`1�C��q�8g(ن���D���!2�g�S�]b	�Jt�n��7�5����[-��i	Đ�e	�����أ�@~BS�e[�W�];�^ �.�v��+��L���#�׏C_q���HqmN�|�L���Ë9eD4�v�]����_��2�W9�5�YC��L��FS
s\S���k��3d�&�3y�Ƈ5�^
����c�;�j��GdRp�R���eKy��^<ǭ�W����y�ޢ`��~[��u��$� �X�Ʀn��B��4��S������_��Ƃ�0����\:q3�q0��S���2��~�A�y�z���Ƒ�YP��꺤�-XNл�2���Q�Wp��7x��7�񕟝�+m�w��x�P���<�fd��b&W{[�g;�% ���e��,^:6ޭ����CZd�F���
�ǯhƂ�gf/b�]/;��iY���Rڌo6��Vi�hN��Zr.Y2�mTM ����e�A���� >�2�����@{�l�A����7hw�W���^�='+�k,:<���`N�6�����&
��{�J�lط̣D�77��wG������*�;@�0P������[��g��q�s��n]<ڋ)�WJ��=͗;Z���2��ϧ��g��v嘷����Ln�ΈE�9���<b��\H#����"�m���̞����}jKx�[���qgz8�zN��-C�C���%�<��:o��C�2�""d=���Y��\�D�\����~84��cx;N�$={�@"@'�|_E��b+�0��%K"&5�*m(���|ܷDh��@k:�--�9l�=�'�'����H��#�j���d��4YA
�2aÞ8��:ٞ�D��uv�����o k�<ZZPM>���6&���@nL�W�%L�geTۻ����5J%�6ͪoe�=��mg>���J��-�48����{G�X�+�^�ke�2K�C�2ӽ-1աsZt�ɨZSI�*��_�׏@[ռ�o������%�Ȉ�!�"i3�A���Dw�BB�h��N8�2O�H�2���k���ơ�l����s����7�r�}�wSR���l���z�
��,7����$�ޔ;0���Y��JM�{<ѵ�xLG8�^�a���|�Y��7���ߟ\��eI�OP����d˷�CRw��F�7ݏW+���#ڍ��t�=��N�ep�v.�q�T�'D»{�q�z��Ov��=.ͨL&V4�}+������y6�NW@�\
4�����@|��QY�̶��{̇jB�C5�#�Y�?]p�lp@ޣI> b)T�(��ȃP���*��Wh�}z�m^��u������a�r!6И��"�y���y3������Z~L�_����w=:U�`���"]��*��z�a6��坈�����i�����֡�(�5�t�^y�X�;��en<y�u,�@l��$O&�Z�B���L��~3��6?�{^����+[ƔQ��9��X�`%?5�2m���>�S,�Cb�ٶ}�r��n/Yv˚���f[iײ�����BՇR�u1����[�շ&+��_l?�C�u���s��m�9����kwY��-"؞5ߟtg*��4��~e�5l8���^u��[��,I1�&w3nZ�3��|gd0�b`���ld�ޠ��{��#G��q�bѣO=����{򌮁o{	��/�uzn'�	�(;O�\sLL ����s��f��Y}��g������[8�A�av�j�`�uꇚ9�^f�k>�C��۹d7v���pѭS��U��ϰ>lP�m��ח!Qc�<{��g1���^fm��(x�͐�� �KtwU3֛�oH�W>Ӑ���W�Xj5fm:�c��"o��w�ѫ�%��U|���6t�?�0���d;g��&a��Z��O� ������i/�r���U����ȵ�H��eu�	����h�f�6�.+�!MA,��3���6���K��`�����&,T8�gfP�#[oFw�V��z'��NE�At�X렜�P%�]6Ϡ�[�W���5p���͛��e�VNN��{��^�\m	�Ms�x�E��61����2��򜣩X�S%��ڋl}�p�����a˥��9�$AoGA�k�0���r]�H�����LO~1�X	�Y�B��@��=�w}�5N1��ȶ���|oD�#a��e��}{����T�H�z*9������/l�ZOB����:l� �Ѹ�lxG�!�!�O�0�H��L��'"�rHs70(錎.��J׫&@�E��9�4��W�������>p���"�}t;QRH�Ȕ�螋�w�ܯuu
����%s�W���^l 4چ�٠vC�Ϝ>6��|�t�-���]_o[�R��)�8*)9�YB��̝qw�Qa@�ph��u�'���N��P�*�չ�X���e���ǝi h=ݝ�gu��R|{sljA���;�<K&»�긯�1>�G�Or���̾���	[Lz��QY�{]�r=�ǵ��+�u�ܱ���⚆1�؎]�F�L�R܌��m_D�L�j����]�����|y�<��Su �����!���9�uH���4-X��:���`��ʎa��K���=3Y���b;_�^ǰ�l�38ls �9�טe�;h��)P6.�Ǫ��Ԫm��*/�3wD�]i�����t.Z�9�dK�p07���m�@ɼ�n�6��n��n���U��mN֬`�D�j�v�z�3�q��?�3��k˼	���C�|a�ˆ��v˞mT�״�0�{O�h��A!�2=��.�D����}YG�
eΩе?$Gu�I����_8^�ek��^=��ƴ��(<5� �VHB���5�˦�z�V�!OR-m9���]��S:#F�qQu5��cOE�5���B׳��*Y�(ߒ��y\"�F��30˅;˶�~Gk�l>銇T: �x�G64����C��i�8�e;R���Bk�q��^5m�(���jA���tz�`W������߇p��΄w��Ol�A{k	Đ�S!#��COb�h5�B��h[��\f^'�.kI�K���_��L��i*�ߣf��q���0�L����#�4dy��溻i(>ݯUвUqS�x�f�UҮ�&}R���B̹�u���؎5��s�(Ż�`���>\�e������c��f���e3�T+nۮb��Hva����Y��//T�k��V�}n�{��($��,�*�T���w��V�GI5>�I:����`����`<;�9�Ð�\ Gð���)�x�K"� n�e^(�a^~/�:#�h�m�����ӯ?F���]������R�1� Gg�����E��R���L��z���1���p��&��W��e8W=g���f�C/?5	��z`&���2��$�yWS�Qx��T4I��w�)sv�a�9��.�2{}B�:`>�P:mg��ݓ�t�lb�Nȫ'<��߱Ao��#UK���4nv̢͓HD�k��:/n<v<G��`}�<���h��m]2Z�:S�.d��3�u�th�Ӽ�%^���*�Y���?a44x�`�DH�^B#��T�X��6Fq�S*c�SV�i��ن�E��i���l����ϧ��棷 0K�gb\3h�`<h�]ss1�m"n*�ln�v���N��Ӏ�n�f��K���I^������+ǃ��1��k�]��YfOWmF�Vګe�u��-�=ۉ*l�k޺$�gv���L��D�%�T�x��62Ι��3%���.��c�кUĳ�}h`(���!�z��^=��ݻ���+ݓE�������zP���[�����ʜpYx֌�
��HZ�;��Xi!���K�+{-<UЊփ��%�=�U<VH$M�j-����lƔ�a�bcȽ7+�e��o1G{��<�y,75�]��,�������4KA�n_݊����έ��y��y��7�*w{���2�L?��/f���xi��!4��&�Nl	����D[.J@f�h��#�!��Rd�o	������V�-^8r��l�|i�����,���E��2=<+ҫ#9��#����]��������:؆A�ZQ)��[xE�з�x/m����B%���	�6(����/�I�|d!B3�f�A8�1,��H�2�Mw���9�<�{w[���'4�"}99R�.l�q�*��� ��xO����~�N��xNH]"�e57�i�Z�ųv*��?foCRq����cP�e���e����Io;�2��1���(���Z�oEK��GV�a̰�p>G�g�"�@@����1��jk�~3=���ؿ0�o���C? a��G>Z/!'�E�r��>�"�{(~�X,�B k�<�f��G�ٖ��_&�3��[P�<�4dct=q�����2B倏�~�U��)���_(���/6��Xhڷ���Ѯ�S��"���c^�I��tu<�R3̮a�p\n��}˻�V�ZQK�[���{���Z��V�q�X�� �ˌ�㶇,�C[�ST�r��w�y�F�Te����8�yc��(D�7�y�<�u�u}���U�T��Ž�5�����'t��Î��Z%^0i<ꥏ
����4�P���M��v����U���%^��}��NȖ��c���B��KEf����oh���c{��.ʧ�Yy�7B\�3�S�:�mM�sq��3����V��.������d�7'S�ē�}t6��+/�6�����>}����g�]���om兀�kZ8nRo^�'ی����GJ���q6`U�.��;��R���onu�*���W!ɔ>4ށʸ�[fam��z�j�Z�b�nvG�mkΪg�NHzT;TM�~��ʜ8k0r%}7����&6M��unP/�5ғ�y��Jݤ�v�j=׶���I�A��fs}Ց�ܧ�����ک����9���KCڜ�^� q��$\�׸!��L�cU��4�b�o0�'j�y�h�D���tF��� k:�'E��o1�[��3�sh����%�Ô.�R��Ex���NR�g�":��%hښ`���:�H��-�jve���P�Ut&�B��]��f���QI.��j�*n�Nv�
Z�Ř���2�����DR���7u�tq��4��ځlaTá���oQ�TDϊ7�h����f��N�Jv���P�̏�;GK圆�I�1�}Ɲ)�4�Ǻ�7Z�Kwz�o ����ɽ����Xӗ"w�
��dz�j�84���P�g�J���M��T�LһH3�簰��i��U��?n��fz��ԟ(z�m$�z�����;D�c�����A:�>1͝��o[ӝ}��0��uzK�X�.u^��y�>�)���s�Q���^(y���sN�l�}�2>5��f���T���w��U6TNF�+s+.Ӣ�V>���:3�cCW?�H]�3'�����z�A|Vm�y�G���c~1;b�V���P�[\��[h����W�^��[}�Y�oX��������v5U�Y�>�.�����78�a\�X"�s��t2:�NO0��/������t��L|�B&��׈h�Є�⥚�
�´���q,��-�\�a�ɼ
����n�qݒa�Lg@S�|�-j�G;�9շd�,�2��|P�eDB��Z��U��AOm��#�ʏyGx[:�5�*ร��tk6� �ڴň(��� �i�u��7k%ˠ�tV|)<٩�����Vti�co��|Nh���Zs.
:���&C��S{)Z�ŻݥP�w!�B3�2�743��{�wl]:��O.��� �-a�ߓ�賱b�G����Mۼl:��}��ohΔR>4���9"��CZ;L�HX�/��w�t�f՗Cc�9��V����|�M��9ݬ=z�D��VK|T� ٹ�ĩ{��������'sۊH�We�݃vV��<��xF��5��wy�����=�g��+Ɍ�cT�Tv�����bj��]�fO'q� 5L������{Rh�E5���T&�4S]��幍������Ǘ�Y5Zg������A�i�M{�я,y����z�h�F�:���0���������{y��m�]��!m���g�<��F�N�GwtQT풓`�_____`�p[>[͠�w5�OF��kb����ւ����m��Y�Gk=n��u@h�]�w]Ath�N���4]�ɪb֍];j(֢h�է5���b.��h�F���.�"���ݷ`�'E5F��۱���O"���	Ѥ���k1]�mA�����;���\L�kl�7\�v4;h��͌y�c%u�:���[Q�Ru�1uѮ��:<�����vv�PkF��1�u[��H ��+���<����0 ��{��M�a��yڟ������օ�X^\uL��V�MJ���j�1�(�Ø6;w�����*�EY3Ϻ�1��Ëy��v��?�O� ������ `��r���-�+fݙ��2�wf�����(~�^�˃�L:��5�?�Nt���0���:�;pI�,X&F�,I1�P��A�7��S���P�ѯ	}��Ba���#4��D�sm�d�EN�W��)�\�]Y�]�[�@�Y�a�k;<����-�0�͉��%~ޠ��s�F�.���몛�ΥZˋ��Rv�B�9�H�`"���o
�D����E�6D�N�zq��lpwO��˲�F3�1���UV���>���h@.���)�A�L�[kR|�x;]��`0&P>�a/����53S�A��i��qy��c�s�k�w��
(����E�z͛eY��Ϲ��=`��"��Iq=�2�wc഻�y�k�
7#6��V0zO�g@���K�]X�F:�������eꩤМ9�V���PfV8"q�C�v�i�d����X�8ǽI�#"QU�rSL����!s6������aE�3��ހ�L��L$� nK�	����2Of"S��y���=�-��~sv!�]�qw6�}��k�8މ1� �a�e5����^��W�(�=TIkM�[��d�ud�l��xnѤ^��s��A��Kj%���/n�TV�����c���w��}����>I���G�:�\c)wgLp����]��:U:��o>zy�3v��Q���nVZ��V���A�KDc�����}�����_P��a��o���FP��|\���(�Y+�I���76^���O�  ��_��O���}�� �x��!�YY��΅�^�4� �IOV'�C"��摋�F����&Q�=__߁��jOM]��2�W�̍�G�9pi�R�ҥR�p�a6J疳P��Q��#�$'�vh�����o��V�kO��Lp�	ړ���@,y�+��u̝qvOy[��]<�eN���O�w�A�c+n��)�c��t%�q�����������dRej���S���6˭�7z�q��J�\>Ȏl�b��Dy��lsH�����-�Û��@��XMd�C�s�]KF��p�G:J�(#R����0���dȗ~��t��m�FC�N��Y���g�v�6l�nAj�¼�Iv��]����"�zcã����C�ydh�/e���5N�q���3-�<ͫ���)���L�1�<i�x?'2�=0�tE��xc�`39��@���bZ����n�V�~�)�n�O�Q�����3! ���*�!�Dך�e�o�S���_��w[U��}9�	��lQ؅�ȟ)�Ց��]_��^,�];�;�i�L��V��u%9�Y5���b��7i`�^��C��t�I*����RV�_:��l�GA�s�Ђb����at]%y��l�+ػ��K�*>ϫ��}C����y���i3�SY�i�h�~�b��s�����{��j�r���.R����%�"O�ҳ2)�9:�\�ڵ0ј����v�U���R������iqi�8�_�j[���� ��GB���n�G���W{�Cq�����h��0�>�2ׅ.ѯؾ�Ģ��c�E"�ËA��V�Ȍm�x.tq��5) *b2o����z��y-�$Ʈ�D<�CM췍*ٹ��h�BA}������A.Qx�E��L��L)�+�P{�����ϱk#��2�re�]��vo8��5;�΀�A��@���]�vEL,r#�I<��L��P�@�S��<!69=��^���ۋ�פ�A�׃��֘B9��n�2$�N��8���'��)Ė4!XS�F��ƛ���S�l!�Ѐ�L�Ƅ���T[�D���,m��Z	Te����G�\����L3���c*|+h$��1ip�� �û���p�_�ӳM���je0���$ꕗ�TN֭`��'\�%�\Ҏi�r�쾠f}0P����s��g�~� ?A�z��� ��/��y���9o�'"�*�����c�Í�u;���MKWHN3tL���)N�fZ��r�N���i�"U��6���U���Z��^��P�V��d}]�
�NY���FRrr�?N��C��
����csX���I���z�D��i�j��7���	(.ӆ%ֲv��gt�JS�u���j��3�߅�l`z��<�ʀ5��z��0�S
�x�˥�Á�u�yN��L:~�7d3l��E���ŠvW�,[=�!ة�����������������<(��;��2����4���- ��CT�!�$��ٗ�x��/Yn�R-���T=�Ȗq������!��E�G�;ϝ��9�n�h��%�uQu�.�Whҙ�2�҅���4]Ls��p����_J\�����(�}�&�\n%��������ߗ�7{�6�ku3Z��Bӈ��O�;a�oN'�cռ.�.�Se�%�.==ڜ�V��&Y��]�?F��XBLW���,q�5Ji=�]8�{i���-��P0�����1S�;|��-a���t�dp�#sP~��/���,L������9�<b�f�v3Vy��X��gbyٲ�1����&�O=�뼡��9!t�eEMm5۷Q�Q��A�nإL����p3[9P͸&82��v
o�����I��NP���ф�R�́��G\66#�wW^��T�\/ꛩ��2�f��N.�+%�Xۙ�5��<� �-��t����Y¬3�������3@��]�;0������"�,v�ť�A`y�aH��Ae�٭d�u�(_w��k�I�ɠ�n.2]c�|���?�"L�L#0��x \����C�=��V���m	�1����}�}6�PB=D&�}�΢�OxT�v�~gw��,��|�PD����t�,�X�%��ܺi�������C�Gզ�?i���4�[|�T���b��W5��E��zF����'�q�=�:5��y��n��F�Ɯ��+V�oKqmy��B��U"��X�{ғ�X�d�̨�yT�6P���f�"��E����ue_�����Ϟ��.���P��C�P�aԦA�k,{z}[~�\����a,�Z�io;�u�(T0gY�z�r�!���=�ha4#�$��df�W��7/�wdI}�������Tq~��������ig&s]ݚ�����i0�͉��oH~~s�LM�*c��ռ����t�m.�dK�i��J��g��
�Z� P�>��=�z@BN�zq��	�U�NSx�m�廛�[�����f��K��/΃XD�6757�ay��CdS����!%��ise(��7�WO��y�wԱ�]	��VY������ ���)ó*�y��e����>�Z�*���.��P-L�o]~�I�g9�hUs��dq̔�����NŨ��vՒ.0K�Rߘ2��p��B|��E(�i
��Z6(�uT��ɿҿ/ï������RJ����3�`6\N�r<]n,����]�WC&U�V��=�����}��I�Y�Y�ZD�O�勔�\���~�ݳX\M�*�9�@��Z�;'�P%�x��g�c��e�u�5J|�B���[W�3�h0.lD�S��4βj�d.z~�c�����#B��<��-pF_M�O���n0֍���z�+�� H�ޏ(2�t&v��v�#�SsP0\JgO����u�"�����].���6,WE8���`q��q�A�i�H8�C)��nr�sK�Y�ﵸSq#b:5�;Q�8ڼ^b���)9\d���1z�[�	�܁AƑB~�|�v�"U5䗉��͆Q�P.�큞�V1];OeJOV)�E��+�X��à�F �պ�'��/�X����S�5&6����K�s@ҡF�L*�rW<�Y�E��RX�;P�Bxwf޲+�/v%)l��_��˧�~d�q7'���uf��,ۙ:��RX]<�n�kӹT�S��T�μ./���� �ȊG�u2�u+=Bc]R9��ȥΥk����zV�Uls��y����]����;t2=�a�LR��0v�:L��6��Ja��j��WHU�{	ArU����mwh�q����gtWc㳷�q�
��r{��J��[a
F�����[Ov��֙����gk�қH��3-RgL��ء�욂�ǉ���띍�u���͕�lu���H�Z�U/��{M�.�l���'\��������� �
�P }���������?o�|���?�5�S�E���<��{�|dK������^#���ş^YY-�[�͛s̝��,�f21e�$�P�.ݏ@q����-�����yy�חxH�v�;{�f:ӶgM�^��W;�k�
�6��a��m>z�M��PiG�A�ʇD���sht�۵C��<& ��U�E�B�B0ZX�xf�'���֑�������{̅��y�cc��+sp��E�e옸u]� `��,9N�$�	�Ʈ�ʖƯ.R��A���tDW��:��~u$ngH��8���XئxBll�q�8�+�-��a�xէ�m��Zb:�ٛB�����ѡI�J�w�zw^�=[�SO����L �`����<�綧C�{��D!��2ɞf$Bc��JueI`����]�M��m�'�|w�$8�1�>�HЭ�Ȟ��[��C��B�>�锝`/Ⱥ�7E2�i0����2a;+����EE	|՜�9Ƣ��2�ܰ)�K��"�H�B�����(�a�aK�)� ���ڵ<���������[�z�jC_x:=���K��07ӎW0����Sr����XD��u�|��W;Rz�t��g(ZʘL�U
��wC\e��Y�F��-�˖�a�jnoT��i�������J�8�ov�N�m#��t*L��_K���S��HL� @�% ��矿����_��})����6<y��@@�64�8Bn�����У�S�� ⮗���OhZ�2�iu���wj iB̘tń;�p��#�6��}���ނ��z�{��5��ϛ���!�������8Lb�����#]Mҡ���9�K��p��:C�C�Z�S�M��`��S,j�=�q��nz9�1nB4�0'�c���R�R��o!u,�=��ɂ��o��_�g��ug�7��L����|zd#a�Y�LxAT��(�|�3�ǡ�g��C1�b�;0�ڦ�mu�̎�ܵ�و�wAװE��)��L2�U>��<~�iʰ��z���L[)r�qT#Q��ɛ������C������/���&�ݬ`�#L��Fκ�|�`��u1gus���na���F�W�"��lK<{D&��!�ZD=�OS�x�s��4�w0���\ZeF[���02\.ak˶�`÷��דi�sͼ4��<z�sKH�Bi����&��^*.
M��C��WY�
!�f�V�-]L�keV��ԎPz͜O@`pϕ0Ք*\���;WP����~�}xw�c�#hFҡ���Zr<~���B�E�b�GoQИK]����9�o��e������2��35��h��W%�j����+'Q���J�m0��#�g㥇�W:���X��1=�#�i(p9w.�E�Y���ݠ���ϝUW�?�����Ȋ��'�~W����������־o*q�)zO�Ԙa�دH}��f{��ɪ~��	���.����8��ҍŷ��:�����E�;f�C���K/7T�<�`������QN&���Fi��)�����|eOK��g��SHI��}Ռ��c�H���vl�0X)�i_A����'�)���w�3�i�?>�׻�tv�Sc!s�O�p�� �5��R͵1���K�R��q#z�$��4����}�5���>A�T��Ԍav���za�!b6��m�{<�^^Z�]ٷx6�F�ejl�/I��%�Qi�7(�a��ȃWp*q���!�������U5Q:k�J�m%�VM7^�k[��R5�=�A>;盨�;�>3�3!�;p��mn�뻲��
q�;[���I͚�L\��[�oJO�x��y�R�B�ʥ��T�[�:|�Y߮�:[U�T�`@p�����D;)��n}�;ML�6y��c�^�3�����*�/(��L�v���B�FzP�`�����Bb���_s��}�3���I��Fi��f������Lu�̹QŇ/���ee����燳�G�� ӥ�2ьAmr�E/>w\�W�AS5(��v�lX�ζ �ZX��j\�)܏:�UbA�(hP>��tʘ�����ٯ�M]�oE�l���R�۹D�!�J?��~|������������G��P��)2 ̊Ь�4�*����o{�Z�{��}�d'?=����ܶ���xg�h�gh��&9���Xޠ��c	��M�G0˛��\�S��D�.�.�/�;�1���z/��x46D����F��i���(�����a歫#V��1Ƣ���>�3���+L��T[ �����^~��`��i*A�N��<ޜ��#ss�l~�e�sW>���Z�#�t�+���=fͲ��l�����k�G���ݰZ�W��@2�d#D.p'���LK���-��WA	��� �ӈc�uc<���c!R5�!�[�/eEÛṗ8��Jq�1<�#T�&���� ���):�{wtSLTm�r��n���#"���Ǫ-���7.ld[<�-�Pf<�uP���;p������P๦'1v��C��̼O.n�^Q]_�4-Z�)�ߣf�O�"�g0�oH�cY� ��:���P���B�k�3ٰ��'O��7�T�HQ��g�x	���%>���76^��[�	r��cY�ʬ�ڸ���QǄ�)��y���WƝ������6Ⱥ���8���:�M�r�_G�xa�B�\�^�5qB����*�c+ts���;���W�	�u�x���^�n��B�`�����:=����i��D�;��)���#kã�f{؁�����V6h�	/�ll4��%wtqQ�o^���f�����!�(&�gw��sd�%� �Ai[y��%"�ˠ��mua�:�Tk�T����oe��*:=8p�l�]�s�҄T;��:���m���ۥ�	¹��P�hf������m�Z�r�o���*ږV�}���jkHS\�;���j�!�����YT:�h��2�Txc���Zs�?�I����Ӫ&u����F�l{��č��y歺�ƅ�C7�O�5����C�
�H����E�3)Hbp�1d��)��S�'V�Q���=�O���� n�l^���k2&��¯�U��1o��'[�*VP�uL��}����y�F��YJ�m��^���f��{d=7p�uP�65�U�u��i�h�Y�u��x*|Θ����SH�'e\؅0�ҹ�����"��J���V�8Kʬ��<k`��]1Q�����C��r�jD�n�m�%Nn�������!%�v�h���6����e-U[I�r��p�,=����J�]����L5�g
o�\B�A�������ƛ����b���²�iVau�����ݹ"p�脩J����{bMd�4�%��m�ˎ
ɨ����N��d�`سFΪ.�A�$��mz١h��fM�GI�����=5;�I��9\J�c����fvޜR�: �u��T̺�%��Ƴ��䙙y�,Y�]�4�,i�
p	��Ce1T�-�I�Y�w��L�<yϲ'��[�}yS�7V�K,Ѭ1��ݧf��y��s5�9.(�-fвq5&��Qmma�ۮ�]�=���&&�uJ��s,�˧���2ԥY��C�'�E�-�h]c��x�;R(v�K�D�3b�w�R�OgX��ަ9�v�Zj���됾
!Mk��Dsy`O-��άv�,:~7���Tx �yr�dLc��N�r���S9��Y���K2���n�˚Tc{cK��-ގoe'R�&����.і�3p�X7��d2�'s��T����Yv=�zJ�X�x�RD����9rR�]�lN.��銆��}�l͊�D�%M�wF�H�	�a���xfn�ũ��6D��m��ݒ�g=z��oNI@�%lO2�]k[/I0gP�Cx&9҆=Mo*(	dt�������a�,=&f6��l��O�R �ki�Lh�;�ma��x�M�ʨ4��m�s-�A�sn���&C][�b���mG�,���4v����V��XZ�g]��u�ؔ��7�����o{7�T�s��>�];6��6\ewU��k��5� �.f7�ϳ!X��M��C��YH�P�j�Ⱥ��gv5AAM�A�Z�7k��:��;�vz-�۰ִQ�Evڻ������>#���1h�GGE����\[n6�wc���5t����=՞��h�ݧ�___W���G�N�裮�շ]wY��`֚���Eݞ��T�3ϯ������	�[����SGA��Q����[7j�u��4m��v�][Vy�����>;���ڳv�ki�q��Uӈ.�V�f�έۋd�7F�����vѴu�E��V횩�����)�SQ��-����b�j�tj�'�����{h�鸜[mX�9�8��(�mb�#mN�buWc�tb���SA�l]�֝[����V�Ah�l�q�u�wDX�ɶ�Q`���[����V7튝������q��VpuݬF5��%Qv5vӍZՊb55��~ �C��י��U[:_��*t�l]5=�꒮W*��,�C}�+kTV$��8�ʦn��m_�#2�mQ�VWϦ�������ﯯ��2 ғ P	@R�0!@)2!@�>�{�{�	e;�:���k'؆���y/��hQ���
�����"�TsrGjd-͚f�<3eV�k'��n��L>��~e�M�qz��V��f�s'\Y*K��c&�0Ƚ�3C�J���R��t?/L���"�~ڠ]N�u���&TjG6��T-[�Z�L&�8�˛�ASF֭�IG��	Q�:��B���Q��ܢ)~>X��潣x�ǩ���u;��3i��-*��˦��q�i�����,�j��.��ƈL3���͆�F��]��um=!;.�9��,݇$�����q�n���:/�Ѝ�⟾���:��s�����!�C�c��z1�l�1;��;ّe�4�$���
<i��I��(#�̤Y}d�"�53nS��\g��l	��O�2R{��Ƕ��֜�$<5� �W	A��9�ٔ3Wa���Cn�y���?[�Fϋ�k(����
�D�%&r�e7�[r����r��)޻1u�m�wK4���֗e
6	�����	���46)��F	��xa�cT�.�2q���]fA^C�8m��\�����S�L]9�ڵY[`i��}Q�J!f��J�U��oN;�,�"��XbqaL֯�6���4�.M���lʾ��CV�I�z^��M�9G�%׭��4�R�vd��"�I����2��－y
ě����nZ{��{��Z(�����+@R�0�-(� %4ЈR�B����ￛ��u��_��M��	��&BeV�
W2����=�^ǫxi�=�� ��S�/�0˜`Ye�I���51u��C�B��Vt�7!	��N��,P
J�w7�Z��	�[��u�k�(�X�w:��v@c���G<�M�H�I��,��n�e^(�aO�\ᷗ\���Ű���������f)��B�l����ק=7W���W�]�vEL/�J.�x�[T�ӧ�4�Ljj$�Ր��ߥ���mxp��0͌�8Bn�0wa�'p�w^8���wa��e�S�54=�(��@�&TI���]���a�2mj�5��$���,C�����,�V�OgZzgcq^Ԩ�ը�s7J�s��ť��8q�t&P���3��d���l��8��z��v����J��r�Z�T�/t�����}�
<�С�ƍ�]��v{�ݛ�yo�7�P�͎Yz;,}Ίc�U&7�Q���=��g��ܳ1a��������>Of�'���A�B`<P��0�9�v�V�m��䠐�=)�g�<��"�Z��to�o��TN����B����!��y>��ۮ��ܑ��յ�����(�zֈ�L�	��P�m��ͺ��G
��kr��0�\o�w�.�9�I/��)�P암��]��Qջ�˰�*�/�.��jf��;������������J��
B��H!� �U� )P(U�R��P�h{���e�腶��!}A�(;�akk|2�;l�K�ИO�>�=se�^��>&���٦	W~��y��pku�)o`�NݙL���#�E��lEC�ȖxAii�6Igld�@��ǳ��9�=�ʴ��=������f���
e.�y�/�y��.+���*�ha�&||�=�vu�l��_Ee�݉~�>8��fq�q*��� ʔ[d��Y�����t	o;`aL�&�4��R�3fe��M�it!G�קk|��;��Jl�2b-)��z-���x�-z/S�#A�<1KޭNݫ�N���S+�\?f�#Db�jЂq^��=�#4�£I�+/H�j���fu���E���3�T��6?�LfʘL�4�'��y��%:O�"S��y��͸�y�'c]�C��E����<��hs�= 80�m0��=˂�`��:g�]Q��ױ���2�]M6��0���8h���(�.�y�Ek�s�]���� ����jc�l��-1���O#9omC��l.�)v�,��/C�Z~X�%�����L$��!��`�ZǸ����퐕/�s��2j���a������֕���d,s�U�W1ʷ���l$.�|)vn�y��)�֑�h���=t5{u6g��
�H�%v���Κ:���`+�鼗����4�C;�fS�6�W��uZF"n!�N�429#_χ����H$ȴ �J��"Ъߟ��{���~�����>�1���E�ʔ�vq�j9�P�#X��Q����5μ�!r�E"����q^��VrXue�;�!H0z�vns�:�W:�R)��6ՃzR~k��d�͊S�U2͙���镳˞��.��C�R�9��'�C��/]S�~}��hZ��K�1���q�����nu���/6�e^�h���q��MjѡHT��_�Q���}K����K�V�q�tV���-X��E�,^9)��o�<	7E�(֡��X/!c���d���~GFV���%��~t�A)��^�.ŧ�c���@��Mϼ�'�k~���x�ӄQ�m3�jKJ�RY�L�g֭���	3忮�sL��@��A�0��ԟ�)��υ;��T�񪺝��i���X{`��["�&�|�bڋ��}(1k�Pb�[>�w�e����_��v��[�[(1���! g����yٿW������'���ըǁ�<��oU���6�=�X��Y#���?�ʣ�R|k-��i�:ɟsX�(��uB���ׂْ.�-��(��M�D ��3~F,SC��͠�z�=�[�����v��!D򛻸�lgQ�d�n����2��m`�d՚2��B�`�د7��r�
����M�ԛr��>�N�~~�����a�($"I��P��)
�*eJU����H�P)F���<=�b��N$C�5`55�]�rT(�UE�5�8����� �����d��'bv^��5�왞�;+�n�(mE���M���)�FE"��qo�L3ݑm
�q��c� ���-�۪�ܬ���7x�v��4��v�)�g	��@��4�����n8�͈�/�j쪼�W��B�sSy�%�_v�ʒ��r�d]`/�4ӳ\��6�;��I�4>eVn7^h���L�.����]��xhO��hQ���L*�J疫7(��*Kn��+�Q*p�w t7̅���:|�񗛛�D�^��ά�P�`9���l�	Ul%ڨ�sm��d�"a��S\�J��	�Z��nX0b[���0&4:�smG��$�2���x���6�;K��`㢠���*9���'Z��;�8a���F��>,�j��Y�Sb�wnF���b�F�u�2ĕa�Mc�a�r��R��z��^�9�dK��vD��d7��׾�n5�J��sy�~�7N�N&���.�^�T�4�h��1ʠ><����2~�� D���ަ�_�U����2�ʹEsWsEq4�n�f�S/c[��W��vb�;W��G����鄛zm��x����x_��2�ở�0o��w�����'5V�;RT��� ᷵ɓ�i?H�V.�*��X�8�x�+fd������B4�-5J3(�!�4#H(�+@4@�R�@REL�D�������ߧ�_�_��"\G�B�yO�+ѷ8��K0�Ȳ�^� ��TB=0ۘ�8��#3{����B</���_gt�H2/�;�t"�j/��c[1���Aw�[qg��;���>d	�BF�Ϛ�%��1p�X̥���G��N�H��;X/�<�0d�ʺcn��֊m�c��֡��GA�fP�a*<����g�b�μ��魬C��#��A���s��E�qYzpr9KBMK�`�M�`&FҡI�We�zw^��LK�_~�e�N�w�K���N��T��ʎLD���>�S�A�	Ll�N���1
J�w7�C_q�=����HuJ���W��O���9� *��_��D�|k�t�N��K&�e�ߜM��U�`��e�+����ν��`ܸm���s�@���& �\�%�n��"U_Qw��]0�U(��vT�ؤwU�v"��5��%�_��6:
4[L���!7W�n��hQ�4��nK>E��0��Okuș����tYt�
��t~n	Ļ�;�C�@`鵤��S�0�3���ٯ~���ٔJ��wmj!��7Z�Z<k5#��B��Pe	Z���h�;x�E^b�c��4ܺ���.M�����j�&m�g�@�UV�UҎVjZ:�,�8sT�Ds&v��+9|�����P쿻��w�����5���I8ű���u��HB4�UP�"L�JL*�L�#J	HCT��@�����g~���g)ݙ�ݝ�y߀_h]�Uz��}�Z�K�p[Sݰ���!��ã�f�F�"��^�m�6�����&��I���6Ö��^*�e�<?[@f�w��B��u�fO�{-cA��G�2�b+�D;M"2�r#qM��*����������5x�f8KD9�jiعWH�k��^z@\l�� ��<��{��:~�7d3l�}(�~����x�l���������ެ-m�ۗD��X@��\H�Se�N�k���c#v����NL�����Y�Ps���� �o�P�Y�--(d�C�$��=�elSp�b�u�sNlFB,܄��v����,%�F=��~7���R�~����ߴ{���s=m�S���e]?DǢ����hEv0�g�.�����9A�b��ǫx]]�#��3��l��թ����e��b�Ӕ%V0*5����%6_A�P��{Uӌ=[�-N�J+3ԍ�`њKFj�x.���x��`f�q�<��dB1W5?B	�1,�ߒ3MI���q����~�3A�JL�aY�"�7˅z+�ȩC�����-�&[�Xd�� �x+��=�{��&5>�CT	Jt���X���W��p�ޫ�p�Pq��k(���<*�p}q�̩�� V�N�R��c���݋�5�CVwa�ٓ/s����I�)JA�A�I�i�J�X�F` ������7	RBL�ُ�M�i��t�On��
HQ%ٲ�0�.ƀF�<����=Q���Y��� �2�v��,PMmq�<�"���8�a��҆m�1��d;�Q�V+i�C�sr��1�w��k�I���V�0�<��_#ϳ�a��K������P����ە�z5Hb��:ԟ��?��/C�Zrp�	}E�w�L$��-���rl$�#)��VG^����{	Ĉxe�Ch�7_��s]��^k֤kI��
��~(�0z�{����)z�g�F���.CZ�̟�uP�u`Ԋc^�k�zRp9�b2m��J|�pT��Wx�425��f��n��}����7�v�E�uCs�{�е`:�Á}eoSou;=�v��痻�^�S��>��m���������<!	�H����;�s���O}���{���ngOc��r�aC�@9^�p��>^2�����e~^���$�<r_!Lk�5�F���ͺ~�"X�ݠ��ث��+�Iv;�ǌs����W��H��y�:bb��x��3=�-7�`���pw&��C2��<hݝ����ԟ=c�)�����]
�^����5��1o۸�q�瑩 &�P0�Z�0��[�\�=���{B7�.�����Q�����K����<����jnM�j/6�j�j���
 (Ba!����o���a�3xz��+h�^,B7?x2-�L+}����s��@̵L�M�{ŝ��dwD1�ִ��y������Qj=��iww��֚K(��4!��8���7kZFH8�rb�VJ@�8Ϣ.)<fٴ���]��X�lgNZ]�
`t���z`�p	�Ȭj����t�ޑ�D跹P��#"����X�Xg���^��[���t�b$��x�mQ���!s���[���������]��&FK�fe��].�N�g�*���jQp��3��-���'b�EZ4D;���8iv!�-���$���F��UE8�S8cz���֌���	
1�%pb���*��*��[���Hp��A��R͡�^�v�wQ��<^g�W�[���QT�����xaպ-<EK>��g5���`�8�Au/��%�_v�)�yM�.���sb恸)�q�h���K�9���+�N�^C������"��z��]F��I�Q�\��,ܢ�6wKh�R�Nbvɞ�jk�a��MS�x� �x(T��Y�x�{�����:��v��h{F��We;�,�ѥ���;	ky�]��Y�>�f4-R�j|�N�����]ef\7w|95��^���m�\�3�:�WZ��\��&�і�X�%RUW�u0ċ�5V�*�����d�%�c�s�����J� ���i	�$bTi���i!��T��O=��߿����y�������)�U�\��{��<k�Cku0}ni&=09�uK=&��J.\��s�[ta��<��8v��EA/m`J�a+hN�sدDut��s�O$�ssĊ�ֽR�H��pζ^���l4�a�XR�m�Mc�v��5-�PzE���̙^j���6����+$I��~˶�G[�ra��2��2�9#�Y�p�ƽ4]���v�i������^�a�\2�[��}u�yw���L��������G=�L�=�^4�$? T�#�V{w/���ݴ�vFMW�-�tM�1�ׁ@�B,�|�I�ME��X��>̂_�����ٞ��*��{��L\��VH"���[�l鋇T:)�, Xt�H����&��**բ����vtB���ȵ�Z�v��l ʖe
6����H���5�g�!64��,��;N���\��)��;����쀽�ˬNԷ5t)���L�����׹n���m1,[O����D����V8�ٮ��[ǚS���{+�4��f�!1��)Օ%�j�]�ɼt k���T�R-��2��ckm괣Oo�6��X\o��71���f-=�y-��.m�W�3�.!$�<�]f��D#���B�5%Y��.��/�&�ck!��D.��X��^���{ ���ᗇ���WBo��.�w_=�>!����w��
죣�!��x�Gv�k�3��e.��ť׫����Vr=z+�+*`]�_P(��*<�-'Ci;duvb뷮����� 0s����vsO&`Jݷi�2f1[��][��u(�Kb5��nB�l$/5�6���)����]��D�ۙ�(�;XZ�v�]p�Ćr����ηvHAc{s�m*�|-�d�$D��ٯ8���I����smh�Ec[�M{��vhh$$�����mՆc���۱��,kW,�l�԰J:`O,�w�2^'s�s�	RS�H���StT-(#�v����s{��������ge�#��Se�VϱX��uQ�
�U�IԨ;��aZR��5s��j�q�-�(�w��7�G��M�9ï�}j�&�^��j�:�9\.�a{o7
�������1��WWv7�N���Bi�wk&� �T箮i0���Է8���Q�/g9��aJ��[y9�u����]�
8�k�����"�e֚q^�EͶ�ր#7x�7n����P����З�.=��9k� �zT9[�7���xƸ���{�� &�oN��}�02m�]�s������q��X�F��X�VPT��˳3��O����Z����bZ�̾,c�;�%��pul��$��!�����mb
����*su�]�0⭬�k�����y�����;�TƇ�x7�mf��8�l�]�Jp�̎�#!�;���ޛ��h��y����,���F	8��.g4���o�*�r��W��Zߖiϑ�B�ܬ9|���{��ۡޒ�;�Z��CFmZ}n�6-5*��~�o�u��Q��</���0�F\��{+�]�znQ�;h���8b�P�v�i�Q�gf��)��0�yp̖2v
����x��EF�r��\�E(R�$��*�r�ӝ�.و�c�'&��ڗ\շ�����ǭ�˲U�+���䝀A�[�RY�[b�^bA�Ei��o��c��e�Z�C�;�P�}K'c��Y5����z5�K��j�t#��fc��j��r���Cx��3W9,�����7�xN�3�!�:�c3� ���̢Ь<ɢ� o�R����2^öw8�����a���_��,ii&�:#gŅN����.-��:uCُ0��7�J�5���Y����[��H��J���O����Y�����͓h�ՂHo%�f���|���&ff���F����L��ڢ�\�[�ʹq���h%�p=!�;f�ޚ���.�ǻr�b���P=eG%�Yv	b�4n�a@
��,�i"N��(�	) 
v�gj:8�m�N�-E�����۸2E���b��*-�nջg�ϯ���CO�i�QQov��+M�tq4G��m�Z�8�`�1��;�����������b-j4bu��kT�kDɈؾ:�8�`ű��荵TM�Ϗ�����Y�X�b�l�mX�6hu�km����Y�tW]A>�������5Z�Q�`�ѭ���(��Fu�X*m���666
36cg�6*��6�ѣI�"5��ڭ��M�ێ��V����UMFۻtkQMb6�鮬ckV��l�ݺ�n6���눺���8��Q�]�[h�qv�����kQ��������1������v�U]8"`���lu���յ�Q��v�1��[V�wQuj�h��`�֍m��cq���E�Ef�mk:��ŌgZ�w��Od�mZ��mo����r��6؃�����J�׽��`���Ի	�d��֞���`�PM��Pv�2�l̉as���K��
�\C�&r2��go��8��a-��aNUƼ�߃o�ޟ|w�h���A���I�J����@�U�hR�P��)P>{����_b�j��/��'�.�~kw�[Az�""�	�_Hƽ���/Ⱥ����ie��&;���Ha���m�zȠ�s	���H�f�	��!�/��T/��ϻ"��!V�����m����4t5�:�{E☝��1��b��p��=4 ��Dp��vv�5�i���jUG]�3�y�bī��Y�O�`�,kˤ��PN%���aÝ��֘pmn�
B�K���!�/��^z4�9�/m԰-X�л�2�-Gs��#��di/Nc���B5��xn9Z'0�������5�$�2랢���*�9t�r���sJ:�}�7,�F-���x��iǆ�����h0e��X��>�b��#!�q�:)�AuI��Q��c��{XE���;|띙��^����Qv��m^Ȱ��z}!�P�f��wh���;��vC6Ⱦ�_��c����X7�j���?ˤx]X�����y	�JH\�lV!�Kýpr��>"T�{���g���1���;sv�'ڙ�������$��i�[�@���A�p;��R�J��у�⢒���_��������W�T+4>l��@�&u�z+;�O�������8vj6��T꽸�0�s Zۗ\�8�-F����qp���U$ZoDa3���-����1V�}k��RQ�t�0�U���B?"��k8��#�.�Å7�|��������� h�(����a�e(B�R�`��xy�xV�M��:��u��>�C�F�f���׊�W���)?4S�%�ʷ�++�Q�����'w?s��� �Yz|�MO�^��3�AqTͶ��E�-����6����v��
�;4^H��	�s�L=���_�]�=Rk%s�^��D���(7y=�U4�OE�3-B�CV�dԪ�J!�q�ۡ�S�/t��8�+"�V�!�O3s��.1,���.ɖ�&�c�W.��f�8�͚�+WMn���:y���c��vl�LƐD��<�AL��׳.�w0rH�΅-�9�ܻ�9K�S*(ҟ=��d�6�C�x��(f�~�/�k�H��eB��aCtӸgmN��VIw<MI��NP�x-�a�^&0�y�<�!��BG�kZ�lK"�gtgQި�
Z��n@Z��^�.�rt�{�Z~X�A/��w �i����Ge��_�]Y���u�wXZaq�>�� \T<7S��Kv�8�5ؓ���(���I��t
s���g��9��?^�߭ݡ�ga��:�o��C�~5�B�ՃR)�&����'�16���Q��{�;|�e��uW�Up%T��@�~�.���ֳ�ì���P���& �=3���ۼ����F?�n�J�ϩl˨�0�nV�=ͮ�-���q�r�\2�|��6�'j��@�|#�R֬�o�R(%��y�����?Y`�	�	��)V��(h
�Cߏߏ�����?S6M/}{2����n��}����C�y��~�n}��д��)�v<����{m5�rcMK�y�	tO�`J�i�����ε
��R�M��*�#�<n�a���w�Q,�G<'��c=�Ѯ�GY�.=�{�@9D�sP/�� ^ø�v}��xq5��S�����}P�N�L��P~|9�B����C�v��w�K�Fx?�(��:���^�z���wgG`�E221�&19�ON6���>ݽ�h�4�x�k �֯ ���H���kw���$�Ue��L�[��Ư\�w�H|aa�-�{W>���֜P�q^91b�e��A���a���ܘ�C����9������c��~��t�D>��
7 ��X�A	��8���VL�MEkV���7KF:�X��g�z���<����W�Q�J+²�uH.��u�"i���xY�����Y�t.�ӏ~&):�dJS<�X�E�a}s��Y�D�Y���p��-PPV�&�t�x�%�
�vBVO75?Bd������4-X
�����a����fjs�R���/��{p���Ҳ����g=�G�1�s}��h]�ݜ���{r���:h�/r?�Ҵ��
������)^A�:��L��x* ��]��`��>&^h�4�d��PNOoE�Wіf�������Py��ON��R8p]�[{��b�i�U�S{����t4�M
SH�P	J%"������������?'~&��p�m��f��/z]���&X^b��J}+�b:l��1�jw�6������c�4�Ѓ�\:���#�o�K*�4��0S֎Sl��/��y���E1��T�#��7ٰ�'�@����Ð��	�:�
6L*��\�һ*�i�;�Mܹ���P�wN��P;)�v����vn�|{��l�����Kq|ꊏt+7t,���;�;Y�v��TL���ũQa@Z��3*u���}njp���`!��@`���$�c�m߈<B��ח#P�(gu7�R��б�~�BTs	hN�{�ÿs��<ͧ��-7�/.f��&����v[�%�7aJ��˦����^��L��pz����x�f�R��^�5[�k��5��X���տX��$������\e۱��2�cX%�Q��f�!���BƄ2�����y"�L�`ө�C�>0�ۜd{��p̋/�A!ꚥ�
�VAr������Xm��m��ڽ�6�ʶ6�$!\H��I�ME��^�kPetmh7�ˣG���h��-̑�
ly�/f0oHFXߦR�6�Ư%[��9�Q=g��暉e��uɋ���T9���]��%�3�pi鱓8@�.s�۾rhP���ۚl��#C�-�u��A�̜���]1J��M[���>-�C��J]��(����  �����)12!0 ҋB ����YP�OS.�ys��6���"gͷN��b��tS<`���I����|�s��Mv<	��!l��e�KRj[��]�vd|e
)I�ͬ:q�F���BW�_��tl��O������nK;�d1N6�l�soA�/��ʭ~t��v:�ܷC�~�/e�mm�����;9�M�k喸��S���^!�sk��ߋħEA`�G@s2	�|�Sl%�+�w�} ���mSWM���B_�8�[�+z��K�/���u����$�kk�qk�l^M��YFF�th�^@c�/¿q�}C�ӪD��]𱓻�m�K���׵���&'Tc����]���,k�9���r�䃥6�����R�:گÍ{o�j�5{���H��%�JX���Y�O�`�,h.��IĻ�;����Y�j��L�_Lf�K���Kv�-JbS�0��'f��*��Q��eO�s�q�KӇ���1�c���}y݋�=(w�)0��y��}�;4ڬOR��P�a>�|is�z/x�_����{���!u�������,=��]j�����BF%���=��Iǫ�s3xI�k+�dt�]��ki�[��>#��}��wo{>�S��r�\��땒L�B�/o�a[���.�73���� ���G�9�v�0w�כ]�m�� >ox7�xy��{���o7�=��<]�m�N�����T��8y��ϡ�����ݲ�Ϸ�L�I��������uS�PSU�������Yg\˾��ؗ���u�zs�S��T�/�v�C�y��Wn�h���n�4�8�zN��-���þ�円���T�{���m���B��cM�d>)�l+��1U&!�D=x�@"Iꆒ�-� lEC��,�9hjC �;n��S��o�Yj��t'b��.���w3Gd��R2a�Ƚ�O~�tR7N���-�w�^y����b���Rͩ����Dde9����7&q�ǒ�m;2>�8������ޜ�Cw���Vdܪ�"wlP��_{˵ࡳ�k��88ƌS���ܪ�	\�W�x�M�aLE�4����y�6)�wװN�8m�+A�3���m���<B��P���r��ث��b:N//v��P���
b��G-�E�.m���,R�I������l������]�϶* �H�謭S���a/3+,�X�h1������������E2��&���j|��U�����������
ﱅ5Z�m�e��G��l쭕��&,�Yr���H��$@#9���r�`c�9#]�z�pj�;�s�}���>	�����{��-�6 u�	������o�p\�۵���k3�/�t4w���2|�S�{2�c�L�����������
̉0�KJC����~y���~�k�a���v
}jy�Hԩ'.򜡰'�[\�y�����}�4[���p�U����W��z���A�3�5k߆.��Λ��='ғ�%�yL��)���m0j'8���[S#+��~�A��.X�vC�X��^���M��u���@�P5��G���ݎ��L�;9�Sj�g3p�P�!z�]� ��v� ��y쟍�B�՚�L\����I��ӷ`fP����u=���P���q�
��|�-��$z�P�O�Q�H�?�f���w�=m�/ۜ�yd�v=��
�l&8��V��7%���GP�n���73׈�ŝ������&7cˑ=����^��ޡ��I��23L(q
���+������(��A{K��o�m��M{=�qٸ�\�D�'�P5�oP~|9�'x�j���q�wtE��sͼ�ҺVn���5ǭ�p�چ;�A�4`Q�"&:�ON6ۜ�Fe�f+L��@��B|�c$�d'��V�oe�;.	q�����k^&Ж3 �-P��l�y�j�����֜P�qG!-�wB�r�]��w��j/����V~����Tõ�r�#=�]�z�.V�89��8��cr-r�@���7 �?���.��(�q�î����s۳��+�D�dsr�V���f�c�q���[z�J?+k{Qvjn�n��n�7�F�ޟ?'��߾����
i�f �������NJA�&�Xo�zq��f۫#��О�Ӽv���4BN����ne��NEc̼Y��I��Tp��\9헗A	��	bWM�鎷��z�8.3���\fLO;r@�U����U����[3rVɣ�o�9�c�yN�����U�?tX<ͣ�Q`)����r{�����nؽ}��������	�]�d��òsh~$�b%:��V��qw�ٶ;��6����3��of���`�U�?C�����f�����Gu*L���X�I�� �mfp��g�����~}�r��O�|k�!?W���0Ǆ�ׯ�;OeIO\��Q�㹤l<��s�mn��WDK#��*f������.�p��C���/)�t����A�)���D:޾���-�h�i�����j8������{m
~(�;	��3��G�~^����6��d���/�ܪ��C�d�@d
TXZ��3!0�`����W����
����(R�z}�癫Juf��۸8Y���!1Z�R�R��б��%�G���Z�!�L�,Pޢ��^>$.V��f��Y��9�.��,E�҇ud�aҘ�[���U�"�kWs��/�9�vv��*,g^H}�-�hL������͙3qk�Z���
s-N�RN���T\�{szR��:�eQ-�uh\����t�n���u����Uc5�|�W������~��/�'� L���	�t�Ekw�o�b��D*`��v��a��
T�]5�~�ӕƥ����.�!�`�Q��1gWks���(T�w��`<!�y�6߮r]�uc�Y�p��$�Wv�w۪�=@�j�(�ؾ�n%K ��l��-��u��0&F���ПE�����Ho�g^��M�&�������ϔ�Pu���!���O�U/o�����`L��Yq"3%'�zǦ��#6[ndN�]�'�i��ƻβ �xc�Ar��|��i�WL\:��g�XE�I��<�34��5���]�S�ClҮu�-[br����T�׳��A��B����ދa�1P潱L�2�X��fj�ɝ�=��O��5������x=�����D���)	�ZT)=�]�.�N��V_D��T4^
��3Wk�!����Ӊ/�&B{+�4��O5?!)���N���1��P\#g��1�u��^�3�?����ɼz��	�[�zC�h�����| 7ƽ#�e'Y��ɭ1��E��w���[���\�����)��!W��|j̍~:4c� 0�¿qC�;`U
�=s�-�B��N�{�n�[m3(3��2���'Mi��Q
������stf�;B���jD�Kz�C)�8h���2a�ٳ�orSe�,e�E��f�3v+�Ƶ����l���%T�/�9�y�9@���Ĝ��6�&�����6�oFd,>�>��I��J���������?;�c�&w��_}�js���^)�f�Cux�S�n���m(f֑G7g(]�j�8��*ۛ�<'�P�+��B��qGz����1>������a��w��}�j�n�,�ù{�k����^��h	�O�0X�'h]��F^�Gs��J�s�q͠�:����f6^�S�d*�.X(�u�;4ڬOQkep�c
�ҵ�r^��>��Ȋ���|��k��õ�3J�E�u#d0l#�=x�6����q�۝6�ʔĆQ��.��Z �]�:�=�������]�:��r�hņv3������y�����t����Pi�l.���o�ᱚ��k��(������vqy���NZ:�;�xA��*l��Y�`����u������%�4��M3�����	\Z	ꆐ_E��b*��΃���E���c���>��8R�P���Eײ�uiѸ��+�K@���0a����ٴ��y����F�T�g�s/U��,��3��- `Q�"22�ߦ��Ϲm�J���vPeB���Q�����4�^��p�Z�=h�%�cPUnvf�yJ����έ�b���9���.��P:|G
Df�����h�ȋ�:�,vk�wks�f�C+yKh�)�l� �#H���g+��ǜ% Z��Ӗ���iǲ�`�i]��U�f�;[��|���,B�c�O��l� �����s+�s�u��I��q��S���[A��n
n�	 R*���h�s�_��e]�fa%��v�kO�H	�������* e	[aL��t8�f\���ЙO;��qт�B��)�y ��*o<�Q��rEE�R��ym8ζx�>�ٽ*�\�R=�����e�!4j���1NXs�6����҆�*a�8U��Cl�.��2�Y�m���Хg|��k�;К�u���l�1Mu�V��G-.�g�>��ofvVˉЛ/3���t<��w�svvոe��	�]J:��&]F@X�So�ej�ٚl�-�DϷ$n1�ٸ�:ci:G�iaL��U:�opU����=�	Q��u>���T�|1�=�]���z�Uz�x�,E��^%��`����`Z���[�g1b�@�Ԩ�typ6>�4;ΘpФR�ґ=��/[u��!�;��� }i��apoIx�x�]w'r�oKo ��ȅ�l`s�+��pr�M��F{���f�GI�ʑogn7N�
ʈU�t�m:.�gP�s�5+M�豖�J�U�=p�i��?-o&��_I�5��Z�|s��Ϯ�w��m"�p����G�
�M���2�k��j�m�d��.i�HK�ɵ�l���5wDCzR�֑ٖC�*�\ĳi�{����<�����P���-�T�9���I�p�Z�"��"�r��ڨ�wP��5�C猬o�#��o�t�η�<�A�n�A�t���^.vµ��}Wj��T���T���_]ude� ��,�ʳ{�7yé��Wor}�����8֛<S;mL�Ek���x�8��[Ek�0ӂ�lu�`2�I����|0N�[֯T�N������=�U<$�CT�wB�ُ����W�Y�i#V@1�^u�rf`\j��c�F���3��Yظ\/wV��b���&"G���͗޼��"���\��2�nwR�j
\�Or�����}�����q*��؍�ͥoV1�������w��b�m��kRsx��Q!�4r��K�I�]a�}|��ЊsD]�y]�-l�eu��c�R�cA��m1�$Zt��\s���!�*��,1��WJ��dA�ǴtwK�ͮj���W�vd�"�}Ȯ<z��̋O:U�:��S[r.�*�w8��$*[��,�P��M��gƷh�î���5���.�D���l �����^s�KQ3[�����.a�j�f>W$h9�ݼ�/4��s��U�gwp4?_^$i�R"��(#�D*#�qT\kY�n�g�E�u�h���5==�gcd����_=�[��Q�b��m���wbۺ�j�#m�w�t�[�U;�ZӠ�]�ݶ�ܓ�ϯ����5����n�E�u��k�lE��V�"ѫN��h1U7\��`���ϯ����Ǻ�o�4�AGF�q��M;kcv�UM,M���;�6M�5�'fƎۮ���9�������35�G�ӫ�q�-�V��v�m��U[b�Ltf���cűֵ�V��5tb�m����k�V���Śi�����v1T�d�b&�-8��%WX����n؍���j�WFz����v�;��cu����mEv�Ϋ����.�buSQ�۝�cm4[;�M�=��RU� �5��b�Gv�kGF�Q�+�u��8�X���b#��ERV-7mwmU4UF� ѭ���N6`��qjmb���؋b��v1u��u��]��X�Tֱ�m�V5h�� ��n��?��������R�;H�h�����ՔШ�G����SUcZ8�4��Rġ��Ve�ÙY
9.�9)�ڎ_ ?}@|+� � � ���y*C+�V_���WH�x[@���D\zz�V0J5�ټD���(2gt�m��n1t2.�Fq��x��z���-��
H���DCϵl�+�1W9���h��Sb�=�<�s��,S�Fi��F�]�u�5{gO4�� H02B�.�T�`�k�脬Ӵسَ�#�1V�k�<s���Juk�S*�F�[X���lz�Y��@0�mq�4R�k؇x�͌T�T70�)�%�b��,�a��]%�N�I��NVy�s�f�U��Laz���͋ �m�9|���X/`�d���p}��iN}�K���tڪܢ����A/@j-#���,6`q1y=�����+`��4l0�`�01�"�p���mt�u��\�`��V�kvu9�/a�E��b�P˟�?����u���������<ò~=2'�i�Ơ�Uv�����~"�7�繱�{�3�M���Ъe�+b�ٶ}���n`@�Di��̎;~�ix5�)v_/6���n�7:P}���c�Ǹ���Ě�^��Mjg��Q�.Q��+�mH���������O���S�u�2']Lw:�\,f��X۟wp}W������9\#�Q��VH���Wiy�vp���Eެ�P;�lrX��$��A�R�Irp����\�r�Յ�k�k5�n��Zѹ�6�օ2:	PM��?�h�����������a&dG�������+U6�i���'a�Nk֕u����Y���sW���,Z���xg������[<����ߴwp�%~��X�궆�8;h?<�Ρ5�h�;����1��^<#1��70��Z�����qp���)�B�K�!�p�}:�=8�np��fY�h�2K���X����*z�=�W
|kO���::���N#�{�d^&��ٻZӊ�ۮ���.Y���Jk5�Lܮl������3�͛eY���K�z���'�A�6(���}�dX]���g��?pߠ8�k�r�-@�5⺱��c��^�����A@��\f�P�mmŲ6]v����쀾�ɨFGs��ʲ8�'K�Jg�K%�8��뜗W���m|��b5MN"ۻf�B��
Y���m�v�����2N]�:�=W�TS����a8�gpK2��l:��[�w�Z������rC��2�V�7�{��#��&X�LU�sȤ�4��#n^��;p�9A��f�xa��"1���^�sϯ�K+�.��ʒ���O3����|�l�B�_v:͑&R����)):��_F�_ᠫ5�U�c�L�tS��&�f����n^P)k)HL6�cl�XaE./N���p�jz�P��Q=k��C�(e5��f�|��u�!������ze�P�)2�͓�r�Sn���?/��<?���2L�ȉ�|���,�:�b9ó��#�sϟx	����G�l:	�a�=_����R�{���G��3\�<֨������2�yj��(%�;0�Bxwf��BÔh��B�������x���~��-�9��j�r�����닰J�½k�>�����Ǵ�ߧ��`�+F��m�z��L�O�Y�{��Á��B�n�2m{�еaԭq�t�{A/mr��Jm��+��|��V��a������H�A������|g���e���,9�
T��Mc�)��V�U,Y�To;)��*�wv�x#�нu�a�OH�x(D&�N����������c��~#T��)��ý�]�/�I�q�t�0;D[�ΟZ� `L�L�u=z��s��wS0�h|�yt���&��S:���q��4��i:"�s�<1�����Yq>��I�ҧ=J[����C��)� 4ƴ�G �����B��5�˦�z�]��S>,7���䔷vͥ���P���/�f�٫����&��B�:�2+2(Q��p��8�����W��/�G=>����'#u��v���*]�O����8]j�ġ���!SwFf�#/�#����5k�^PU���t��
�R�\����l.�9sA�U�8XC�ܽI�k:�V�DE����/5ДGfm%`��X?>io]}��}��������fe	��}���T3�b&��cZD8��v1��ږ�8���<6&=P]%"]0�vP���iw3��ֻ��s*���q�ۯ�ǆ��1���2a	�";��Cv(�����6ħGj�zb�WB㏰�P.��C��߲Mֳ��h�:8�y-�:A�	�� �Ƽ_�q�x��9B;p^-�η�1(�b�1�)��#�,�l���>�HP͓��s��9Cs�$%.2a�[����+�����.�r�E��tS*z����Ni��6��l�;66e�w?��1��oTv�-Jc�1����I�UU��f-?5��.��^N%��}2��7���5�ծ~�Ԙ=64�"uzby��,V�.�*��Z��3t�w=,������s6r�ss��k�Ds,z9���M����V%X.��~*	{�$7�.���9E�l�E�Ωf>;@�_L4E�|��f��Y��4�y�L�
�����,#�����..i�in� ��q��1چc�,3��`3?�h�]�5�zv?v���tg��3`h.��Rd�z�(,=g�m:v�|W� �u,c^K����e|h՝��NJt:�se�y�.��В�V!��E�x�VY��0�诱հRuLѓ����k�/�f�(w�1�SKpq맮A���{V�`�;���r'�s��>�y����o7��.��(~j�����߃픟���^���^b�'DS��Ǟ�x9a����Y颶E�)�v�S�;��c#6���t�!�Ë@ ��l/���툨~��,���uAo�w�����sK`��B���{9�S���h�4P�X�YA
ɇ����N����\�<�1�¡�Y��)��T��#Z|A��Nnj}<�7&q�rTͶvPeB�����y��K-,ل�����u�1�Q���k�E;ǰ8��Ƚ���J�`��v+��Bk{��s��x�Ǘ�������.{J����]v���9����2��0D���@$<�V�"�q79E�C�n�l�������:�5�x��I���VMw获���ΞE�;ą$lIvl��^tE�\���]7D��R�ִ����9w���)�FSStu�3c�0�X:=b��{ؗu+f�n�n�,��E�f0�7gd�>���$�4�ሤ�ct�5�+\a`[ ��o��
T��.���g���a��B9��1��@��j/~¥�E�mO�ϭA��%� �s0L[O��X�.���_Qv'�8���-d�>��V����Y���w�����9^⋓��W\����U��ELfY��5�b�w�s�0,�wq���\H�ي�`f.Kz�̺��xm8�dʔ�J��o��u��4JVj�F�fu�":�o����������y��y����g�IC������q��,"�)kL91ߙs��ɦ��U�v�/2���Py�3 �fjȻ��P�wHsT:a'���8�;��ga�����}S�OL��ZjE1��ʬS1o�A�v�O\g*���m��͉\�~k��y�S�
�Y��-ݛu�5�G�~/0���"0I�W���f�ؗᥥ���f�Ja��1���O�nMsI}�~�4Y��
���ߦ[�o�C
o��m�no�C�-za��q�rQq�23M�kZڳ�E�c���`�4;s���.��nḃB%��P1��|��aW�x9�G���2�{�9=��X��)�4�-ۭì����t<ٵ�X�o���8�6}���&*||��>Jy��|���͋��;U��ҳxǞw*�v�7/m��
���P�*�[�0�`��Ⱦ	��WXݭn�ݺ�޵K�q�����82��72(�0��e�`c:r��@X�8!'����A�OEt�SqY������BLV5q��Y�A��LJٶs�o�^ʋ�5p��o���͡�vUP�;,z�r��&�3�ՙ�Xܺ��O�m���]����.c����Q�Uq�����]�b�0�f�Y�fJD�@֢s��4R�Jp����u�Gnuk*I�c��*��nb@����������z�Z$=	B4�]%Ҽ���469#X��(d<z~����`�`�`<=4�Ce)9%gSW4;C4C4`�-.+�`���K��Z�dv�A����):���+UE�5-�ƯuE���f�7�r�u+wk�n�Å�����_�],�&R����kxi���EˈL��)�FE%3��C��۹�g�b��z�"͹
�+Qm
�q�cH}���!���Y�4���H�I��6���&�N��
����ԡ��-&�����O6�`AƘr�8#� ��,��ӳ�v	�*�6Ru���bu�����9�Ax�QiAl���w�~y󇶀C��>�!�=�B��I�����o�E��Dw�P�[�=�XJ%s�PnQy����v������f�w�`������ҡ��L$�T	��m�n#Zi�^K�U�,���(�<�Z��3b�kׄHC���je,�{_�_�X����� ��O�M�="9�;UL�n���+�{��Ombz9���:Ɔ�ջ��;v�o;�u�g���>��7���s^��e�;h��0�@�.�ǿq�i�^��I�P1�{��7&�]�T���^�dj.�Q���	�����vd�$������o1�ׯ+�j���UL��xyoMj�N�g /C���׌��dp)�v��?.6�k�^�Z�Ь|p~r/��kٻ%����5}�Au��I��#��}f�u懨DZq=�Z'l�6cN�-�:ӬwRVV�9��a�)M�}���f
$��f������y���a�� E.���h�]N߀.�c�\fb]��ǜS9|��N�0&|8F�B|`�Ql�}��/0"���Ddo3af�`��x�C׊�;��2�tE�����466�%��2£f^L��k,�m�U�����-y�>��A�vAҸj&��.2�5t�îyg�o��UG,mU�fx�w����Z.�ؚ�jW�ʖ��P?�P2�J�8zzq��b�f�N��F���հ�lS<[@�0�}#����%bv�t���%6�*AeV�
Oy��q�Wʩ�Gj��ެ�8�qHrޝׯz���S�_�����K�?���k�x�7b�m�Jc��	ee��M���\hl�|��έ���,PR�w�ɼz��	��
l	��0O7�9C�T#M�54tk���2����"�k�=%�kθA����։�DCy8\���^c^��#2rn/S�G*oZ����S��9�>r��C]��;�׏8z���\��Wn���aW|!3[(�	�	����P��S��9i��=�NZ�Ab�y��$u��R����;~��3b�3&cÍ�W#v���N��[����z��<Tk%�r��Y�n��_�O���0�'+��j��f�[o�cqu�Gn8-���9.vRg�] �z�ZƲ�p��NI�`!��\��\Ik�#/i�v���U���"x���)��	��M��>�ɉ.�`�-d� �F^��q=�jT�]��s�]g�ֳ!��C+zp�/�8�Dk,:=í~��mQ�Z�!	VS��ҵ�0e��O=ks��D��p�~���Uѫ��1}0P�!�s��g�`�f�4�M��:L,����>�)�-�;Z���7B��;>�z�3��v��1a����Ap��:�_q��LDk��igE?z��!�N9C�C1�-JO��1�3�qh�8�zwDS���GD��A��#Y#ׯ�2��s�<�D��{�5��&�ͬa#L��$��i/��m�b*��ix��mj*�hB{�c<��Z�m��OE�����7p�4vA`xPB�2a�����
�6��s'n�]��Xwй�^}O,�,Aid�{{�;5>�ODnL�R��V�ˢ�'�Adv��ʛ���T�kQ����[>���..�8�ʘ(T�(~�_~\��6�񔴿���ᣂ��[�z�~�ԏ=��qR�!�bQ:���W�E���o����(���@$;�6(��<�3Yr⯞2�,Wy����[HN�nM͌n4A��ֱn�"�m�n��q�Yu�huu�\"gC�he��r�P�� �ebU
¸�4&������i�Ӎ���U%J[�cy���Qb-"Wd׼x��Psn}�ik�N����F�#`�E�9��/�����
����*���A�Ơ^��y��x��c��/�v2�Nv��].ͫ�	���#���\���'�)��t�e@i5���W5��çM(K��u���K5��}b���Gt��!��K�R/����2��1����H��,km�/UF=I��O���]�����l!#�C�ۘ�� ^�5¡ۅ�mOC�Z~Y�Y�@f��ixW�AWhD�_4�zi���z`u��i�s�ge�ck���g*�
��mOv�ٜ��gOk�] ���YN'��>9=xM_��?	�P2U��/�ݰ�Δ�غCƐ��tM.7f�!��Ѧ��d��FM��)� �e�+b�ٶv3���~/�j�Ut�SDu�l�����N�T2sKUL�0�c�����Ě�-����#a�>��&!�s�ܸ�]��g��ܝ��bz�����T#��$��bXo�p��m�c���dY\�ܡSY�f''���_�8��ρ����	�&9_�hk%c:����C��v�2�[��/cX���ʧ���"�ff?�N&���I)�.F��L�:I��w.}ٙE�YW����5b-Z�ģ<�g����˚�Y��4�(�c�l���42Lq��u�F�@��KJ�ka������f�Ź�wL��ec*!�l�k�.�>�#�7Z��mn�0��QX��U��&��4��m��<�f�:"Cu>m@�F�Z����.�p�� ��I�k>�ʎ�1�a��K����� B�f%ـ���`�6�w"��q��ؤ������­o�Z#�����+�gj6�8�#}XN�"�K�s[襺�D2].U�;e��Jc-Nxl��j����2��!����8A|v��ˆ�ӹhK���|���W�;�v}��WRZyZ��V���p���`8���r��]ٓ�n<Idj������P$LY�i>��3�_8��WiE]xv�cS��u�zP`u��˕�,���ѹS�j�$�F_T�p�m���o��2B�.��M��kN��4��2���M܎�
:��!d�E���[���]0�V�+2�o]�ս����l��v�@�ũ�0���7��ۮ���[r��B��pפ�{l.�֤�X��o~.�����W)�� �Ե'���֛%����I��/j��)\�c��?|^�u�&�pr�[���{�9�Z�F(3 �%���]�Ho<xU������p��Q]�m��h��d�B�)�^^�z�L���/���rj1�(�
�@��VA�f����clc{�������Emw��|��7��r.rv>��nQ�Ӹe�n�m"�Ԛ�#�P��׼����I�E^�AT�}��
i��Juy ��bտ�����'�d}�Mc�T��Éu���c/D=�f\�[��杝�F	�7���h�*^��{���B���γ���	�ͩ,n�%�z��gbݵ.1�8G_;���&�vL��[�Z��|P�s���oh4���v:݆1��}Y0*�l)�St١�ޣ���ߗF����n���q�,���=�{ �mn{m�
��Ix+��k,�ӝ����>�S.֍�up�{9�@�K+�wpH�b���{�I��ٞ��I?2���h���ۺb�L��n���@�↶w+ngF�Ƶ�w�_�jWr�[f��.g%��'��le�����_Эsw(�\�X�*�]�V.�l�6�����5b�����Y��J�u�����t�;�z�z���7ok�>ס���Ι�)�e�
Q�h�,Q�*���u��c;�K3�[�KPnLt�ݍm�v�>�6�:kZ�K������,��]N%��U�.`6�@1��+1�|U��	��w�of`�KE��UCp,���'W-��6jA7�2�z5]����_��V�:�	�I�L�I���Zm�T�U�B񪹘�id�-��w8cx��Ç7�u>����&�ˠAN�7wǟUo��+u�gى�5KC?8�\U]qsݮz�؝��������i4�����~__�LQV��X�=n��N�m-�I�n��"��'�lm���RWv�U9��������X����lf���klmI��mb���v�b*Ӫ/{[h�
��h��i�}}}}~/k�'F*�h,٢��1{��v�5�Tn�5u�[RlV���y������v��Ѱ{tv�1Z����A�M�V����I���f�DA]�1��j��ۢ�&1���ګlv:7m8��u�ws�F��;��Żkh����ݻQ���UW]�����u��ն�1������(�u�n��&�����wY�*�N��f-��uh�ͭFKgU�����tQ�5QQkZ��ƒ�ډ��V�`��6���u��m؋PT�j�"mlhы���GZ��đVΦ�D펝�lh�l7g��`�(��D4wnf6�س��c���Pݭ��MQ�b�b��`�j��/���4bU��I�� n9���0��
w��I��zࡍ��2�j9�m�!���.��(h���M;�0����CV��p[	�ml�̛\:n�n�(XL�I����I��j��C�_>��O��t
�U�"��m����ts����aZG��\��m��vd�!�wk��;�)�xl�ߘ��y3�.�d5N1C��i�ִ��O6E;�~�C����
�?x�q�}�VAl��˅[���/Y���9Z�l��3��l�,qL�'�zw�`���I�+�t�-�"�7Xa�j���6���D�'"��t�Z��	�Z�,J�u;>��2��G�Xj�3.�?&�K�$�����f��x�����T�|uϯЃ,~/)�M
W�TXS-�����2$=���6jM����Ƴ�#�Р�5��Nې��;%73s�I��N���k����B���zü���j��b�.ȶ�^���>1� �؆Vl�pi��i��&O��ѡp����:��C[,�	�\x�6#���w�xa>܀��p�'��<!���W�Қ�I��L�� �e�.'ܥ����V��賀�nn��=�����p�*��#�9f
��뵭ޒ.��tDf�"'�VS���(�*,*�rW<� \��`�,h�u�
����G4pooR'�XAV�ٖ/?t����ǔ}[rc���~����xiy�j\�����E߶���G�֍^��N,,�}�7�������ծCwڭ��Uʯ�n^�JpޮZ���԰6�IA�oWV֐��#�g�
��i*��V_+�w�v����˛�n8k�Dh[j)93r(���J�ƷJ�Z�K�>ӷ=�v�9��~�t�d�~�2���"݃Bnj[*zG6���ԭq�t,~��$�6J�a�^��԰y���Z^U��p���S-|�[�0��f�F�3����-�Ûp�M#�.��O�n��t�oyIxWo�b��{��B���<)Ɂ��ǴBax�����T2N�,��y����Y��ǣYɶ�i{�x�e�]���3t=1��-���˼ydh�.���>00^��bb�s)F�젟�����SZi�f=��0<��za���e@tM�1�׀��5��}�W�J�sq�fv8A�\�5�m{������� �%��5��m:m3}0��L"z�ob����u�wg^��=�θ�E��x�ƞ�#*[���PY�(�TyÁ1�zLմ�=���#|>����|f*WE3Ǿ͍��q�����	�=��)������)�!��R~�1s}<��d\!��9B��Vk�M<5��;A-�'_!�C;+�VE�%SA2����q�J���vɥ}���֢�7��`t9���j���o
)JSv벝y����:<s[�r��	�g�����}b�%!f:����i�ly�+v�\��*�]I_�\�q�x��B2��Ⱥ�ќ�"���<��mpU5-�cz�8����������WYD"�D�0��5�'��W�T�	��J�vd�=k�:y�������P�ڭ����v�7)l>��p�}>C��N��d]s�.*}��t�q|)��6��w��D���*1B���<�iץ�c+GO��ߢ(wE�L,RK�n�eAoP��Y�6�zo5Vڜ}��sp����`�9e`Lm�ΡJ�N�E�S��^��qPX��0��Z00\s�z⪹+�b�����e���A��ƑF���u[S�0��.�	Te�֣X�K�Ȏ�4����a�b��*�w�x�%`�H6"���a�tz�Z�ڴ	�ʠ��S���5�X�K^M�Z6�o:	G�{�@
�Y�^�>�C#�H!���E��h��8~�~q����sݣ�d�|䶡��`XF����u��s�f�9�3�H�ϣ�<!��5V͚�"�3uCj���:P����}�}$������U!�S�}�E�[)��^� 
�뒆�ެ���c���"��p"%M��;����#cm.H}��I�C*�v��n�H{��ʹ]���
��o���O�����0�m���fˠwMNޱ���9cq�!��B�b˷ ��W��7k¤�Ok��"p�/*��n�,$�t9�b�llj��3H�;l��mUY/\YI1c����6�?����u�M�.:�Wb�tv�g(��|��;��[��>��g�4@��E�i�z�x�{��3�f��%�����f3��-��Іk9�Ep˵0��?�.
�K�a�z�*��ɯ�>�ɜjԕ3���q�S�v��tD��p�6i�`Y�Pz͛OC���w�aŴ��q�Sl	��-=\9�mN��E.x0�������l���ɫ֢K��u���]���~5������F���Wd��$�@_	󧙹�N�}4����eaQ�T�����Ξ@��u�Ć����Sgi�������Bc�n�@ᝒy��$�D�I@�\Q���#�C��{գ|�'�ࣧ��N����������D?[p���q�*@I��&*ۤQR7��V��5x��y��V�NF�z|�<l[�"mLpm��^jO���}���x�3�`�ʮ�Z�t(k�1ϗ��a摴vi�s�`�B�XF�����!�s���Z���M҇o@��&[/KB���1b��4,�La���M��xwh���>`�a�q�u�D��6��lj���9��3Y��\��>Gi�g,\I�R�ܰX��~Ca�~�zO��ERm���ʲy��KW�]��_b+Aj\4��S�}RۜS!�)SZ[��v�I°���#��ɷ}��Ca�غs8d�.�p�7��f�}~^�����V`-D㞘ڣ�c]�JN*�O��?~��ɪ�MP�K���6_T�#�շыxpS�@L6�/^]�W���졉��y�w��2ע�t��B�i�A�;B�v����sdM�w�N�~�֘2��
�Za�o=;_k8�ꓴ���23L+�;�9>&+����F���ݾf��n	?__�G�!ѣ���=b���^@L�l��>ÝC��v�����b��a�v_2�����c��hz/��u;����*.ߌ���}�����F�B�;oe'ٙ���	t���b_ZӁ\�o��fq��y�����<��6od�K*���uc�]?kZ�ZgE�r+�b�\ �
2of�P�ΞG=;Ń.%�D�vqֶ��kr�1K�!ֽ0Q91���+b��oAO�ga��P%�{�^��k*5h�wMA:pB������\�d,
tD��a�dώ����e�б�0�PX�Q����6^�͸��M�sN�m����q�ֱ�ی��{g��szf��I�r�SsS�!��į���{4=�P�ј�h�*;��Ġ�4+P���6������[ov����nZ��opV.�*���on#����9�ղ£.k�NTV6K �X�pɯ*���ιZG`��<]�QR���-SHT�pr#�r9��d�=rl��b2����� 7"�:�N7�C�G��H�2�z�Y�4��2/�ע�UU�=҄��ϱsB	�J�<�OEq�A�+�����	́#}��L9�I���2��Ve���ɮ��c<�[;M=y�T��)�u��O�sH�;5��]�0zl=�� ڿ��s��4�%��w����j:�ˤ����aPrW<���_�P[��{n��$�lVQ��l���L����;��Ј�=mEs��(0u�X%QaV�y�إZ�K�k_B�W:�d�Tm���y�V�Зs0�	��dk.�"�:��+�Jײ����� 6��SP�&�us�k��x��m�ҙ4��08�fpF�4�|O"2�W��s�R�`��	`L��"���2ѵ�yג�9\�[�����^�9����?�YK!刏ߏ��`�[u�>�)766K��nKU�.��2���8̉b���KG�$����lX�n�#���j1���.�%�Wc�ʂǗ���XJ���$�"
���]`�Ռޛ��P��������V=���d
��B⫘������Z0�]��b+z)
28��]>a]�S�5�$����o��ft�<O3;/�[a��3!����4.�[;�&�C������ujW>ϮU�vk\�&D�N�򆕛��oZ����FQW����rgꯏ����0o�s�y��V�p�5¯��і���kNd� ���HB����q��&����vkX_2~�e�z�Y�`�a;��q%�j�nT�5.R%lA�A�,���.M�"}q�3&�-��e�w>4�;,�S��0���I��T�}��:�l�k<A�����t�Xڹ��3�dX[7!�XA��s�?B�4�<Kw2掍3��@���&�<�)*�ϵs��=4��@�#5ڕ�ʓ6��pܙ��#����GT�鄔��yl�{�U��-���=���LL�0����~g.����q�j�jު��'L�$7I����˶���s��FL�퍽��Ԛ���vU��}]��^�0SP6�'z����|���v�`Du�>�h	���)G���h;�9=�C9mW��-�"mq��#6d��������6�M0s��(q�Ì8�/������T\X��9�"O�=���!���]�_��m:4çB
�u��H�X#B<�^a��O[�`#n'�]g,v��J��r�9X.×�unT	��e�ǹ}��S��6V�{�ݹ���ʝ{����F���˯��|��w	��sb�����v�Ę�5Q;[��#�Q5�����g��#��q��;4Ta١c ,�͙t4OVd�N��Y��+�t��!�=��}ݓ6C���q+���Y�^x.W��k�<?zmzc��-�w���$�a��V ���zt�>�v��X��'��Q�6:�a<7���>��mk�2WV��m�I�{��q�Юn)w��(���2���%�b�tvT3�*�u3�NJ����l��ٗs>�g�b����"zz��fS�p؝qoA�R�6x�L��w���1iQG@ͥr��Z��lw/9c ���b��r6;t)HY^PSJ:G�@�䋚sB�U�����^V<E�ݝ�4ݬ�_ː��v�����
�2���S� �^�u��'���\O]�}z�jzY��v�c\[����n;H��I[I�QU0SՕm���skCV�����\r�':���}�>KWU��C�F����<�[wk[�K3�,�87E݋��,��C���q��\{z�f��z�)MṴj�n�=7�wB�h�.����Mr�r"4��W��on�QV���:f���_of��vg\��8n�if��>�{W��^�!t��M�E�6�$��q��r��m�Z���"f���c�T�3���N]���+^jleٵ�e��s�Lή�K��i�ֶgd����p��#z��ؘ1�����3�T��^¼yL�]J1�?s��,�v��!����g`����/"�3�`ŝͽ-�Q�
y'*��Jin�W���"u����VgF�n[MSn��Ugo�peBkڠS�� n*T䮦:��� ��2�o��\I��v�yޣ�4G��p�XMF��k��z��rc�M3�\3���Q������G{y;A�t3�����WP���w7���\�f��wfs���Os����xq烢�K�y���	K�Z+o��34�l���o^𚼈��ͩY8A�$?��$灋mP�2��7ܸB��#�1_����uZ�;h�\7���\��%ǅ�ys�ܛԕwR��9	S�ZoJ8foS�Ѯ����[��|�W�|"�����Y��;&�ٵ�nSE�`�r\�$n؎[���ۓ��U�� D��GF�I�����b���K�>�=��r��l�ꉥTs-;������Y+z�`�m~��j#�[M]bٓ���H�F<�R�,����K(vg�T� �V}馫n���b�~���Px�ўu7�4F@w"��B1t��׸��t�dv��O1U��< k����,4��8At[���mm6���]������֬<������c}����Ԣ�r:�ݑu����!M�>��Q7.�i�l$��~4`�߇:E_<���l���N[Ә���T�(��3H���wg:ǶG�*�sG��-P����6.m�v{��j��]u/�owY;}����^{�.�֧��*���h�4]�w�J�v�;��WQ��jL����K/<�W�,kZ�fR�f�3g���˕Z�1^����L=3;<�LV����EK�&�3c�5��.|�]�Rp�_�j��  �\�/0���-��&��v�v�;�u��L\	Z54��r�83���7�4��oU%��2X�����s��#���'��wf�oX�_RnS2�IGMeC���O�˾�9u
H�I�s�+ދ3���=Ȭ�-
�{"xs��Q4�UgR�fnzA����Y��s�[L5�3P�\�굶�a�;��T�.Q���{Kr�X���`P#�.�0�����;b�KG^ʂ�RG�=�:]��.��G�\�uYyFR����ܵ�d�6�X��;�j]�E8l���1������է{`ųvbE��/�����R(4����d�ޡ�J����__a�N�}U�Z|��O�*�gv�0�"�-7Q�G�^5�])ں���rq��NvEB�v�ئ`�v�,gE�)��M���4+�Ln}ԯ�3Z
�^���0��ǝ��}; ��m�@Q�Lf�z���ą$�����um���Jb��a�/ *�\��9ɝ�v��&��6�(�U1�q�fi.�Ƹ�&�X[@7he��֠)��9�u�:ɻ�]�m����J�V��J� �"ˤ�u�G_t��e��-���b�~�IME$$:�r���{��{o�MN�����(٥QSv�Wj������¨.��X��7Tr�f*��v���3�OEz�Nu|D{ע������V�j�1F�u����XR�M�;L�bU�TN�����]K���;��Β�8"Ql-���Y$�:&���Nk.-ё���+h=O�1��T�M�KkU��e`V���:[�ٽ)Mhmu�E�hñlP��o��v�ŷ,�#�� ]��`��i@�I�2�k^�'�Xn�9ݴ��b���}o��
5��Y����hV`��K�O{Rg0��Z����;���G{��f�d6V�,���d�z�A>��^҆�w�zT���w*#����9e���]�����7�R���<�r�k�j�=��r���f!-���ܵ�k��N5+S|��}dY�s��ѷ����3GNp�E,h�,=��v���L9�Do\��{��'����\�h���#ݷ!dl�ґ�c&?'W���7�d��rK�O����U�o�\ȥ�9TX�-u6��U��7R���#�n��B �.�Xn��e�:��{MQc��x��P�B�VS;�I��,��:o���+���u���/4	��r�P���މ�o5c�]=n��u�	�;v ���X�+����t�D.h��Og;K9�g$���+ʫ���E�{��a��w{��9�7�C�O�xj���§�cu ���ǜ+�ג^���_>��)	�I�:���ڃԵ;�dMB��ƺ����<U�,����x�8.�(����s2�͖L�Loe88�n������';������o�~)��Z�mCT��f;mbݺ"⣧����V�j�Z&b�4SZ4�����j;pg�����������F��Z��D�[uv��0�f8��v4��a��uۺ"
�Q��s���y�������}��Mi�*�����Km��u�m��EVƪJӚ�5E]�:-ݣ�Ů�F�tu�N�3ϯ�����5W��5��vk��v1լ��s�*4n��uEQZƌv5�F�Gq�����h��y������1D���c�W�qZ#�����l;o յtuFƊ��tI�D�jzM^y�UU��lVѺ5u��)��ADT���)��i��o6��j)�u�V�A���ɪ�؈�;c�Ͷ�[�wc��)����Zf(��QEEETlcV؎�]��(�6,ZƛF��84DUD5���Z�DM�9�4=��!�
��EM�������I���Ψ�ӂ���I����*��GV�Ti4ӎ��I�c�ws�i�ڈ�n�=q�R�.ƚ�QX�l���ۮ��E�|�|wy��~~}��ݰ<��62�5܌w]��M�)�vVkλ{
:2!�I'ᮔ6�EF�\Ǒ�x�8�g�|��{��{�g��]"���r��9�ɉDx9A*{g
����S�M2�X�;�e����f��ލ�Ttc�����]=[���}_�kU���2Uxo�܄�(�.0F��u���=>�o���ݚbDr:m���_n��ѥ:���ó-�gw	�$�x@ח�hw�i��gn'�S $tF����n{7w1��zQ�$�&)�_�n�_���uPs��]�\n)��@��5������!j+lACk����m�6�nE�c�R}������N��Ⱥ���>C�UFF3v�[S�T���Q$�L@�ѶO.UV�*V�䁛W"���[:��lHx��y����_G.%����,�,HZ]��Z����\�i�2�[Ď́�9��|�yr���Gl0z(���ҤwJH���d�x�~���ubr��X.��k���o|z{�wf��ӏ��P$9��4��;ɘF%Gʦ:�����~��b�2�^R��jॄT�6���p��.��u�fğ%���"���0�\�G;��u�:�z����G豈�y��LtR;m�$�<X��BEC����u6i�vy+�mҧ�f�a6��w&A��ܽ̽-ϯ�PY6G�S���dƭ��4S[�GW=���&��i�����=ݼ]�yE���WC����O�d��� �Q#�g�?��5��X��q�6�añ�!���zcgU<Z��q
�Sm�i�讎~���V�g(����?��>�O�7|�ȇ#�cf�瞎������p��B2�Q�+d7a����q�;#�7n�T>>��F�fMR}͎��>>�g֟Ɠ_���ރ�ܥ��-�cg�^5�O�Ԇ��i�U��B�f�b�
��e�����N�D�c-T���cU3N�b/�� ]ˑt)N�?H�g�Bw�R�7�����u�;0������w��'U-XG�r���rY�t@AU��JO�q�2�N`j��e��s&��`�׸�s��N'.�U�(6I(g��CCx���6�&�^��7�d�h���q;R���<'N�:i�ϱ�k���\��c5�u�?a�:Z����;U�p�Se����z�Dp������b�y������?�h/;f�:a㹨Dp�ֽd�q��m"����R.�l4�7gly�H��h��չ�]�lc�==��,��Q��m��\Ӛog�U�Q�p��ݽ����,�:5ijY������)$o��\�����������5��{�gw�%��,��NE�%��ơ���ڑ�rt�Kk �כ��Zc_oC>�̬}��ۧ3�P�t�y�(�mR/y�zRL(6��W8��t��uYt:7v��W�a�������w�����2e���kc�̵n����^&�6�l�vJ�;��r���2ڛ\w��ucը��[�z6珲rz�g�|:�l�rF(������k�bŁ~Q��>򎮺�&߄Qu�Zb��,M�䦖�{�J�R6v�2��T����~<7W�1G�.��?�{$nT䮠�VW��UA��|�
�-3�*r�3/0
�N!��8��7B��(��:4{�|D�$o_SuiB��|b�ÈI�_o�;�{*27N!��d���T�n�v3�#B�p78v�v���D�"3]�"U
4
����p,��u013xb9Y�+{Gn�7���C�>bC�#Q��o���z��eo�9�����yf�ޤp���SE��������2�f�́o��uE�F���wQ�j�ჼ�S��o����7.<����9�d3�G�sΟ<$&��B�����[O��=Dg(̴t�
#kߤQj���i,�y�jvx/�*Q��m����	��<M�]��!�;2
�$��͋�V���:#�)��aUc�n�R,�3
�����dY��Y�;`Ȣ��+���*��R�/&h���z>����&!�a�7
T����B��ax"�vs.e���ݲ���.{ӸA�����L���8���t�����kk����CVꗺȭ�{	�x�]�Y��QRc�P{�;��GfH�I�!6~���Fmb����/v�>�G=���a�T��|�;!��ϳ#"fC�FLmC����pd��5����sF�;��6+l㱺ؓ.6�KsX���D*�墌��r�SR��`�3�&ù
�4CtF��MU�Z:�B9ko�Ǹ�g*]:-���d1��D�nt�ݬ���XP�A�z�(�J�l�429.r+绽Q�æ���*r��hrU{T�7��/ҷ���s��t_��<��Y�`�8�½�@���f;/��8�&�"Wo7��t�g�[k���i���>Ϙ�ǲ}R�v��fR�6��ew.D]�7C�[���ɷ��''{d�6M:B��O��!��0K�;V��Ҡ�e�����Z�*޴�O?~�_���jXPbT��n%G��\�y�=�V��N�Ck�8�P˦��`ލ��f��� !����ti�ٝ齉���b3��٭�1��ǳEor�q�'�u���=�m̎��TBJ�>c4��&������������H27q��I�(�$�pL��S��>I퉳Z4Ɩn����L�lDjC�R#*�n�fI��H�:K�-�5|h�T�w	���T����8@!&��~���z����\���UUF%�w��T��m�vن�'��q�y�^�h�Ȏ�q�(U`��dp��/fͫ�1�S�z7ڲXr�i"�ի�o��.$	���0Y��<���&�0��4�tb��3\!z@*ތ�.Ɩ��ڃZ�!�OY9&��BN5���U^�2�1l��3;Xص�H������Q�6� �?q/4�[<ȻȺ��/��˙���]ܒ��w������s"��q�k�1�95w�ga�'�-�,�	z`ØO��,�7 ����R���JJ���F�(�e����N_l��б��C��W�/�wBK������#�O��d��a�hF��gg��y#�~]��g[(�-͞K���n��W��~:���Hs}�z��o��M�T�����?�>���ol�ΓVSA��^�Y�X��8{vGn�����ػ�)��FN���0�� ?�`�X��wF���XĪ��u6�kA����0��s�}�vA���M����<7�0k���kN��@[,��5�F�z爌��=J��[EQR��X����e�;�ga������K�T�$nuV�v�o)�c��O�U�L�al�������vĥ:����Iu������lt�Ԫ�\c^L}n)-I��ء��[)u�=[[�N<Z��	w8�M��z�b�\�sC���]��[ͷǔ���d��rT��U������ɇ���=��`$Z���g����[��D�:��m�琸'B��B�v~��~�_~�o���n6�.��y��oF����L�RJ�"o;��w@����AP`<+5S�1+��tyf$i$T�v�Nf(��B��ޱ�v��`$��}�*��:�j!Ю���y�<�{�׸�$���'M,S�n�����y*K�K�J�lS��K8��&��H���o�_x����T�YZW�h$�O��2M�Eiͥ>��Q���΋ӱ��R�Q�#�qTȍ��.2O���(�㶨ג�9�q=v�+��#��l�������V���Ӫ����jW��T��JzFv��kk<q�z	��T��l��t*D"�n7��R47�{h�Q������;�o
H�j��t��1�d��Ы�M�}{̲�}=&�VS�t��|� �@k�����f>� ��_������j�E�_��;V��X/ι��,�>ݛ�G-;��'� �olR�ףsu��Z�0i8e�*=��v��:A��(8��������Y�+)i��D�S�	4=���+;3k�k>��8b[)K�%v������I�Am��v@��;��P�<��zǭ4������������?W�Q8G�ԇ�������R�9�%��*z�Ǝ��>�H�'�4�����D���bW�{{���G0gs�m����8��J����V����D�T���N��'i޵�2���s��S�k��a�Fz{'pҠ���;�	�wP�}A�N��R]�x�HZސ�}��!sv#���E���i���0E�q���h��G���1�v̎��:����5WT_$��ؽ���a�NCgO<���i�7 �h��+}WĽp���q�B#� R�t�D�I٘�[��U%3�G�/����,	�#���i�6-�F��_�����\�i��<��$��=�4M]P�Ⱦ$wa�V���+%����5���z�&0�"��r�6Y�@q��z�M��~\���QRoxv~�����"
�t��'���.����$rS�J<�u����2�;ȈVts��4mI.�j��j�aԸ�w8;h��{q�1�U
9�U�ef��"t�u��m��)��O�os̨2�Q��r̉�#��m���u�7)�+Zާ�]|�ڂ!S��W�s�b_�����`�=b7	�h�b��*l·+oSe�!�MVY ��P��Tv�z=5-H�\��a|*u��;&/s���փ�G��[�xJ�EH1Ʃ��r�vfH��%{���ܜ�f�:�g'
�8�(���'�"�Ҥ�lm�S�÷��`�k��*�U暻$Q{7"حR���u�U�W�b�� ��-C;K��UX���Bp(#���0�:��5󄞎.�2���͡�M㚫��'A�GfC�v5�<�;���ޭ�(�o��	ڢQ:��7j�����p�{�ͨ����z%��r3`0��gO+��\�X�Wjf_&�g]����	��C�u+�жF�Sv�G5���)�L�Lֲ��ۻn�l�D�k4���CF�.��i������|l1�C��4C"}t�]M���w9�]6��(�i��ZF��;���
$[[sF������D��9�CG��X���J�1��ĳ�L<Ր�^���mf�̫+V�ɣ�*T�;��	a�۫b[Dj�ݻ9��Z3����L��Ԏ7�����N3��m�{�]>��q�2D�-���v	�m�i,��36No�|ݶ�D����iW�e�7����l��D� �~�ɵ.���?����� �Ϩ������&��C�SWF���b!��<��M��	�yA=�--�?Հrق^�~�,w@A(w��3���
e�<[���i��]h.!HWfR�i�婹�2�:���s��Y<4�Zv:�����Z;��4s��8�Uhʥ=}�����W���s��`~��I=�/z������8H�� �P�y*��Wc���ִ=CDgd<�7n^s�mAZ���������RV^��x�L+� [̾5{xn}���Nf��.�]RA��Q��ٱ�h�H��2]�=83M��<��ݑg��A���,� �#�]��ʫI�Æz�H����M���2n~z���Q�n��9�f긫y<�g�4<F��:��ڭ�%\T]�u�̎�*Q i�fjO�L���B��S�����p��`�)�G��k;8��s�?z��>�!b�Z7z�_����HW%�dGˋ��Q�q���e��닂�c��;�[�:	v2t7��%Mzr�,�����M�5���ʪ�����/�X+u��U���m+y�c;1ƅч#�C�uV�;݊�y��8��(��:�X2�[���&�vw*�/It�l$���;��P��_ic �t�G%�Ϭ����/�3w+��#�\�� �MR�0���9���՛��GҖuŷ̷*�8A,>�kl�0�q�8��퍬P1uk�.��j��,W]KU ͒����yu+��MTB��f�g7q�����JK�q�_J#��#�՛����PS�4���.�B˙g��Wj�)����
�r�k�E 4��f����㋳*p��:�u�|��-�V]��_c�e�\j�EY��H�d>C�l�=�-��Aw�0a!#�� tɃ�靁C��cT�O�auY��(>��l�t���[�z�� ��f7�[�w�wm1���3q�M��p9���՞�s�O��Q�
��նdYݫU��m�C�l��H�!-B^St�sT-�ݙ�/�jKI18�����͒;�iˮ��6�c��bGg6����i�7W��B�eY�$�t������Ɖ7�K�>��Ȁ-�uN�q/F��ږ̌mH�pGx��87̔�s˨+���w75n
c7"�:��bof-�.nT�8jP!3}t������E�`̣�wS�{�m�-��ۀ1x��h�`*��]Ø��յ�D���������[S�����nu���k�[)J����f���⬧Z�5�{
�/~�췸�;b���髩��CbdL�lg@Ia�
����<Ah�R8t��,uШz�ĭ�X폞�դ�j�9TmA��^IiI:�ir(:�b1V�g)5jʍav,6���d�r=��%��o8G�͚	4q	�ӊ���.��JA2\�*Rꚦ��Ȳ����:[�k��Ư�PK3�i.��+z�^���z]��x�M�2rS.�z�:��{z�Y�&�2�!
���\X놚Q�����9t;Zcy��Ԫ6����)MJ�c�<ܜ����Ϊbj���*�D��:,-@�q� i�����G4��(1�T7����<T�
��y(pج�/N�1^1w�f�^�24��R�Y%҈Q�Ʋ�n�o�a��Cu�qܮ��C�éb.p�Lj�ݭ���S�f��H}��XN!}�mm�z��Wu�I�t��뼼!.�]�v"�e�tǮw9�1,��Wg;�V1NXb�.���u�;vW;��J��ˏZ�ںTv�T�qL��s���s�H4��!�]Q�8K�,�S���O�S@�5�^Ѡ���&�v2U�ŵ��E[Z("7q���)�n�m���lU:�IT�����__J���/lUA�lwn�lTDX٣X�Z
�F����l����� �ֳT�SDĝ�X�*	ϯ�����٦�)��Ɖ*�(��4m-PDb��.���SF���4V�Z	�����Zh�& �ѣE��� ��&K��TT�&�T�4v1!�X ��TA�������������ذ����=���w`����Z7gLQE�;��k�ښ�N(�X"j����T�m���*�d:{cE�h�Fֈ���SQ�v�T��5E5Z��T�*�4h��i�����Ѷ)�Qu�(.��{*(�sQQF�	Eֈ�4P���N�TTLQ:�]u5V���F��kERQZ�l[DQF�
58�C�+=g���z�j
�Ս�t��th��e��-��lSA��֘�j���}��f����d�]fS��������꾇K�=�30���{��
�t���->���꒎λ�"o;��M��'�fs��n <�<(�B��ńH���M��NZ��ǩ.�ד/5V�����iV�+���'[l��d��X#5{��Wl�t����ړ2�Ƞ�m�����Z���h��,;��y�l��t�n��ޖ�*.OP�= ?u*R��D�P��e��Rw�Bm�?v�W߷��'A ߏ�k�y�����N��l�o��ԧ+�s��X֤�DlM�al������|���})��5�c����2���o��zg�ͷ�s�f�j���S</�\��8��l;� �	,ꎈ�J�[o���-��i��*�pe��O�E���:�3�D7� ��$d3�=���J�u�mI���ڧ��w�3�2;��wh>�Eb/����rYŎ�AA���ܗ��~��ޭaWZ}�N=�$$u�g��Em������ao����#�����=��~��0�r��ظ�<B�PSJ;���ז͚T�J���W�����eAY`+��?]n���g#�p3���Mw���co���:A�j�Ֆ$]B����Z0�m@�.����NyqGգ4s<��8��TJ�ǅ��zH���'u�iq�?6��Wőd�M	u�o�D�F��p�Ȧ ��Zm��/�`��iՀ=���
�}*a�� ���һ�Ӈ����F�mˌ��#U���p 'S�!����;HmH�x�{�[��mwxC��[�}�R(��~���*..<�~)�A�썫f>��Ԉ؎�~b�ͱ�x�Ga:��a�ُm.��-�^�E������\����\�E:�}ڮEm����K��>ŭl��^�@w7@a��Ai"�WYgH�1�=?k����~D��1���2:���$`��]�Y��4h��w�{i{엾���;�#o�X.[�:��ѧ'*��S�[����@���4w]g��� ��ߛ�.�=���+\���VCK�C��ci�#.����u��N��φ���g���tW��ez5��Ù�p������͗3�|1xˠ8���1��du1��9��p�q�mf�d�Qc��o�Uj�4���?�47%�o�������dʏ��Rd���·5��ݼ�TLmo.���-|eAC,������mZ<�*���ll�c�=+q�u�Βq�Sq��V>MB�W5:c ؽp�I�WV��w>��
�ݺ~��ޯ+8�X��}>�$��>��w��p�^;H��g(�LwT��a
{�,�p�:|�@sW�cufZ�{ŁDa�x嶹�̽qKs.�Ƽ�>>Wc���2"�P����fG��9�]�G�hI\"sk-�,EfE9�sw�c�Wc�j�t5aP*��S�g��rY���qm\9���_/Q��?5�{Τ���u�� �,A����-gy5���H�z�MD�KLOh� ��MxΪ�v��#�� ��� i9�AL~�v��TF�w�[\p"��Z�F�^����Mr�n[���,�,��KFY����U���FZ`n�F��(t-+����T�-|6��`�Z�7�>�A�q�}6+T���h뒫T�65��j-����vX�˻�ꅗ{~8�|?n�w�g�_%޻Q�S����<ӵ#C��.i�7��|1)��MYB 1鰡��I,
�y�;�:��pg.\���
�GG��9╒){6�ٜ:���=�Rv�F3�cy�0X&&�[ҮRǎw�X�^�DN�U��Jhfi���+�k�X5J�;x��5ݝf85���:n����O��\������Lr=]3��3f}g���*7q��:ni�ǫã����H�QR�d��K�`���l��]"3�G\��ͱ������� �����ҽ�Q5w�]~��'��?�������۳�9�>W矃xm�z��Ie�z^�y�zw�'Nea�'��U�ss�u[4X���p�6)C³Q��@�o���'�u����<��_8|��I�ߟ��[����}�Z�</�����9m�ć$��_����uNm�C&��X�Ǘ���p��,�zJE]nM�{7`�C�4�}<�A�e�?_&2v�+Fn��/)H觏l5�A(G��5�	��x'�}qsG���5��^ҏv�ɕ٤�v6��SsNz���N�3�{��܎oC?(!º�d8�k���JR��j�%́V�q�����������NWrE�C�W�TՅyy3I	�1�/(0�jL�9iwi�9�2ڙ%ͫ�he V��If��gQ����*+�����O-+���R�|xة���b[P-�Y����q��g�kn-�ѹM��]a��S*v����
 V����y���#b�� 5:�<�)0�����6�'��Ꝭ��+��>��1��w�⫁[�OJJ��4�g��51�y����v�R��l�ӭa�m�[u���ћ<��oP���#��^�P�k�|�M���>���M� C��Dg�u��W��S�f9SV�]�<7�C�u�$
&|��O�����WS��ᲭDĬ
63v�ZTm��F���P%�K9��wd]&�_���~ݺU4��׳�w�D��I� ��ҥ���Җ�(����`\�'��x�<����jֹ������E�v���ܝ��Y��t������P�8���wi�}w³��Cc�cڙ�!3���3�'p���=^��̈́�*l������|n_r�,��S�(���k�����<+5�Vko^>���L栢P=�iI]���V���(LB�޼�+��enA���p�ڱ��7}��1C,����SW�)���L�Q����I�[+����P!�w4����t%�c�=��Ot�j�?�jg^�gT��U�wZ�r��9-�^�7�����yz3q�;�3!�h
���H��e%$:�0�-��Ny�z�s��!���r4X������m��g���=(;�u�Uk+��q3:�J>���#����|MGsiH�d�ܲ�9yo��YNdDX;���vA)@{�sz^��.!eqAO�(�;K$�z"�v�8!�q��!�qꈹ�����f��.���ы�7`+�%
����1�9r���"�/�av�ϵ[�m ����H�n���W>8C�xL��	�{0�`V�(�����O~�����~�t�F�]H@��N��n�;�(f�tt7Kk"��́�)YsƆ��uu�-��6�/�N�2s���ꌾ��Zj;DI�:٭�s���yR�a>��Z����R�K;jj ��S�j�,t��O��O����'O^�������������{�����mC����K�A`3����JΥ��!�v����3������ Ɣ�~�S�z��y��{^_Yvl�([�Ex�>��3J-��.go0Õn!n�*�e0���@��6��	4�#R�]��˼�O)�w��r{7�P��_^ks��0^���;�`��;3��I�W�ؘ��o���a���"{�y%R�J�GH�S�y���p��t�H�5�V ��3�)�r�{�����ksO��U�[ �����{|�C�B/�Y��'!uS��g��k��oqc��rc�	���g�1���ᣙ�,�N��0�Vj�7ղ9ev��m|�"5$�o7G��f���/xOC~c}�k֮��u#h*1�ʅ7�gGpR��x �}z�dn��C�.;ņ�F���[kDB��FG9�[�=����� ��	�����U����hu��p��푓���c���}Y&u[����f;DM��k�ض���g_
����R�U�n����r�4��O~6�vӿm::�7�� ��{|v�ͽ$1#.��俍�z���;y�/��A�8z�N�%�߳l�c��������~p_Y�����O��u����m[xn��L��}�/��Þ��w搭�PVxd�����7w���a���z��pRa�o���s�}�c\�sf=I@q%������S��{D+=۽���ѵ��!�O
��춤�����&8�0{�RاY�̋䦉g|�Y�۽{��Q
@�6h�[ۮ�΀E_������l�u�S۷}|֏3��t���2��mi���-뒨j�����L����֫�S��n����vXc���~�u����*8�����1�dM�v�C��(��L��J���5�����l�F(��[{�m݁�^9�3;�}��=��aV�7�$m�r3`0�o��V�7q�M�Fܴ��^\޻�E&�����Z���R�+����Rݛ���EM�����ťpVo�8� ?1��^��"Yt�1r7�g݆�x�c�4ғS����U����C/H����L���Ƈ#�uqr�U��u.��jLׂ�ƿ��3Z ��������~�	���$���J�(�+V�t�{z��%����^�ı�)��Il�
��6�|g��ؤۘ�PK��r"���p�z��xZ~�AT��/$w��U���$	L�=;w�ݢb���X�.��*q��_n�5������[O,���5mt�,]��F��4!�+s�N�놁 h�S�q�͛�Fu��&�Z#����ʹ6�9ﮰtbϐ���6���v��H���H����&gwC�w� ����>]6�6Ŏ�A��U\h�=3yx�N9ݗ~��7�s��m��)
��]�"���ӝ��*����id빵=�i�g�8O�,ޡ3�WE#D��g�V��K��/ZV`�8"i�..ݶ�X�-�]�Ob�nAjtt�W��@���9;(N��v��˽�����14�?�+��d�Jp"<+_���RVxE󳱻cwvy��8��r�?WK]9��>�����?*��N�k[��6e��r�5�sR]E+�d,ݟw_Hb����y��l�ջ��dHK�u�����5�$V+�E�btw�j�=$p�z��:wCe�C�����.�T��GM̨����+�Or��Q��ww��O���cU�m��p�Up���7��)��%5�A\Xe�e�MKˠa���,�r�ub&�^K�h��?Gz�2mN&Ve,l՝�!c�G��������f�$@���g˓�
�������{
�"�����ny�ml젹��";u�)��k�����zEGu�-,�Gi�Yޝ&A ����Y̻���I���o�X)*����L]刳�4�]��y���6�!�F}�7$f뎵a�h�5�yNB��x��n9�����T�UohF�n���s"�G�d����<ܶu'�tX9��boLp}���X܃ѳ��/��A�]����f�q)��#����f��9�6K��rsǂ���x�dlS��3�Ю+_r�c{5B����Yܣ�ڮu���.�KC��&��%�+)Ww�"�e� `j^ӛ�Z����CU�"T�ǼҐ���m*i��H.�������hm�z���Y�+�c�y��Du�1o���,�rAM(��u�6crjڮ���Æ��+ʴ�>�;8@�
���V�����&����B�op~U��I��v�u[�l�@.r)�Y�����q��b]5Ri��t��\�擜�U,�8��M�7�F��';�û^��Ŷs%qL*����C��D>����]XZ���U�&��95�U�1��yLk���>T4pU��5d��u�[��P���n��]��gqn����=fZxgSo��(�F�g��gTW��`�}f����J8�uy���f�ݒ��:�d�Rऎm��0v������WQ���f})L}ӷ�����.�L�\n�y"�������N������̣�\����@Sk7��P֖� ���B�����[T:�,�M�J*mV���l�}�����U���:�ս]Yض���:S@<�Iz%ɑV*<f��#��[�%k`���C.����zhL�:�*�Q�f�������ȬrH_u��Ewe�R��� W;r�Rc��S��J귔o�d��j�s�!uCo�ӽg��\Ԭ�
洎Cf�)C(�F���|y��?t�Ppy���YB�2��o0a��y35�n}q��K� �9����0S8/+'���#ܙq�Q|���X�rv��X�-��\�R���k��ʡyB8�0���|�8&<m2{I���V"3Z�*,�F﫜P�����.q͍;WW�sf:;K7�ΤN�ݕ�$�cja�2�xl ���<����f����j��d:',�%���ɕB��!��Q�wM�(�7�e��[c�:�.m�8-���5����gD�[N�Lݜ�����Iη�si�)f���G�f���Bw�����{��K�q��:��%����UN�&���.�m�;���'�<��Fj�zR��Ȕ��V"��a9�y¶h��u��n�{.y���5y]�qS����gи����s�Ӯ
֝���>#7r�T]�g�q_]�ji�d��V��ѵZG[{�ۼ8�uERt����F�U��K�K׫O@�56J���927P�X���5��K����I"���0꺕�+q��
^Q��;������ޅ&�"5@M�� }S���mw ^�A���U�|h�9l핶8��H�R��7�rQ��I�j�[M��6�P�����������2\�5�7��C7s �%^����e&����-�H��	�x�ƪ�h\�񋷖��7��9)�cl&k3m�@����������=�.�n��L���Z�0e�ŷ/����g5�(>��7Jq����e�º�7�t:ˑaE�>R�ʵ�c\m�h̖΃L���WgT���.�f^���ηB�G��wtNg�zʻ�Y=�qr.gm� �LN�V�	�t��b�'O��j�-�6c����Jx�8P�Lp�鸺��C�u���70\�_��;.�����Wd�yʟ�.V%�\�Nɔ:J�t�Jn\Goj:��2�v>���U�Ȑ��S즮*̎a�����Ir[7S�N��t�'T!P��T4�E5�ӯ��:kQ�-6؊��"�n�v6�b"*s������ET^�&��MSTi�����A����c6�t�$�.']i�>�����ϲ[4�mu��)�5l衣�b����Eti.ƺ�5UcBj�>������Q@S4AUE^��-V�b�-:�E��j".�h�j�4�____C��ϰ�C�h���cR�l)�X4� ��q:(+Z�Cvt�uE4�TSN�I�[bj�Z�C�QE43MV�CI��kZtb+u�a֩��SCAD�tUA���b(����N�*t�#Z�������։�lm��bh������ִ��h&�
h�δh"tj�l�`3Rth�H��FJ����tPV�l]`�f���)�bժJi)-�Qi&�U���,Ege��F#�f(��c�kl&��~~{�������ح������=`k_a�(�G7����k����Qn⊷�nf�r5cuT�U�:�n�-n������(�mo��f��Y�x&���US�O���ip ppO�8��/��Sx�Dt��dU�n�Ih�\u������lǁ�Ͻ= )���5z��@M ���l)�ָ/#d�5ʗ$۾�����ɷ�k�s�ՋA~�hA��;!��>�[���|�@�[\�F(��ܶL�ص' ���f��5;�-�O�^�@�wG�q؍Y�h�-��+�sV�z�ǃ����z!��v����FN��0���Of�ep���p�9��k=���z��(��T�[/h6������8��EQ	��-\�����Ŀk4���	���ɍ��Nّ��C8��B�r��dm����+�5x7@G%˸u��1�B���QE�p�#����V\LՈ��� ���h�{Y�{P��F�Ne��4�$A�v�j���/2cI5;X��DP����M�*�@����R�<xQԻ7c��-��K[n$�ͽ��v�f2R�r'����g2�H��)Y����
�.�Ȁ�;7�Dj°���N7���P����b�U.��2w �+>��˼Ԥ���s)��C�?_{��"�4P��[0�و�j�2�{���a�?5E>B��4�\C�M�74G�'dj�]B���L�X6y���r��S�lK�I���&8L�n� � ړA.֓��\�P��+�惿	�%\�}z�z�dp~���ǫÊ2s$׌�o:%�<�@@���c���G�<L���U@����a�v@mI �$Q\c�S�)r�'�"�Z��N�f�5,��#�ՋC;��:8Nw{v���_��7R�Z�N���9�)�)�w����h�Ce:��A`
�6+L��,��r�ڥq�ŷ����P|����8OAv��K��e>;=,1�	VH~�к �3�|�	�GI�S�7O�W;L���d�7����|0~�|v�@}[ճ%4��<��gH��۞�~�����(��b�+u�j�(�}Y��Z�l���_�f����i���[�1C1���=�%�O�Ar��!g"(h�G�	��C��{��HMzM����,i�S��[:�ێ�^%j�F'^��m��ގ�]��.���Q/�^�O�7"�e�\Ё��������d hd�F��P��2f	�����j��E��_���Tj��^Z��Ǻ������ݾkJ��<Xmwlj�ճyݍ�+�m���YG�e�u�.w�dv,1�\'���d`Y�՚����(<�PaC�T2��,��j�C��<[�9l���}���s7v+����r1[�@賏
���{�ve�vf�w�xr-f�g���Qy���́~B�IX�����+"����UV�����w`y��l�=ɦ�<��P�A)����u����U��S�&.G\\��%�u*��K�����ӝ���1.��V�һ��=3���(Э�Q�nё g���%C�i¥j{ ��]�s`H���F�Z1���rR��g:��&��ȉ���]!�:�z|�!\ ꇐ�9v����y�s"l��W;Lc�L�1�,��d�G�|q��/����5N˿5Ìx��z�ӽӠ��[�Г���|�j�w�д��t���r�� �=m����oQ9OX�@�#Y)�V��l��_��/<{�7e릱��v3�և���W3�)�B��g�v^$��1[�뺇!5���'y}#R���%G�?��P��^����n���ɞ<_�?G
�X���Em	࣭��N�;M�<A�1��M��d�*��&Vn����-�
p����m�\��8�6��̞�=�T�v��h �؝9�.�%o>�#'[m�r7p���9C�#��p�,�����8��Ay<����x�big<��6�A�~���q��u��D�?gks��@��%�T�����Q��-�
&����wŌ�f�[��|$7ױ�:��8�,1���nu*V�vr�~�x�QM�v��+rC�U��ч��̓[�!����}�[U�J�1��tf�m���&�27�n{�dGh����-����y�Y�!F����m��:-Vct,��t�'�����,Ϻ)�r�~��#7�:���Od��:�R�(߻n�����X�%�VR��Ns8��po;�"�&y���sV]��.���J*�c0�EcÈ�|�Z�
�$x��F��QGP�xpP�ܡ��im!�vXO,�:�䳵�҈��x�ڑ� l-�9_7�Ff8q굕�f=>:�J�z��U�Iu�WN��,α��*�ii4��-�DʝM����-�p������r2t�'�:K�OEb�ļ�ͫ�Y��k��[��8���P�2Y/o�����M
2��VQ:���s��s��y6�����ysN�� ���Ԟ�5,x�v�F��f�mT�n�&%�{F��T2�t`;W��M6zt�S��=V34)��ת�Ffc��W��[��}!�'��%I��[euө���R�?(��WѝKMGl�te�/KGt����xk�R��_P��f8��b��M���^rb;x�:H���Z�=�J�R��ֶ;��1ٱ��Y���_b���;���u�ޱ�vzz���[���S�&��f�.�.}fmD^��\gfuGK�G\���Iל��k�3S�ne�kp��1BJ�R3e�z�Fl���`t�2���图�,
w���ɧϰ��q�õ��(cg�YN�K(���4�տz���q��p2
E��Oq$V���0�ꡚf���k�/�A+v�7ek�q����1x1��7����]q;W�s'Oq������h�*QŁt�"�vPۛ����]Cs�O�y�[���|�q>kѶb����h�cި��kVl��6��^�deb��c����&:A�2:��k٪�*P��'��/Ygv�;�3��nb,K���TZ�o�tY��1�y����E��l�MX��n�j���h��Zg�ouh��2�|IQ�C�Qyr�F��=��Dd�<���O�C
 !Fݢ�77��-8����&5oq4�XH���Da�7��+$��w�U�π�I�`؉�����-���]�7o���D;�p�Rk�v��׾��s:X&�A`���LUu������������VqU�-�+���FuU��	�s_��ϵ+yۙ����$�{cg�לo�{l추�gK�EH1Ʃ�#q��"􇌖i9L�
�����v��C�#�X8V��7a#`s�U��MJ]]_,xs����ef>n�-��c��ǫ�����M��N��*H7�JJ���<��W��gS��;v-{8�:��2p�*�+���ZI�)i�fM� ���J�T�؍K�H�ޱ\m�pj���&IA[N���$R'S'_�
Wb�F��j�bĕ7v��F���{E���R-cϹ{�Kw+t���b�K��F�i�^�-�J�3W1������ݨ����ˣΎm�v{�N5�¡0jX?�!��z��+1�}�5�3��kK�EF�]�w�H�;#�5�,�����.ǘs5'��Ow�Ɇ۞��-e�c�q�V��B����`�l���mQ�̹ŗ{'P���仴�A��Z�x�R�\���Z�7�n�;k2:��sn�	��ǜ��7#/��R5�]7CA����q��e������1;]^���87�N�222��ј2=Z���$8�8��LŘ�U]�~�t�gn#pOH�n����e�I�x����b���kǫr�$�1�ϵ1����m��D��G���}|�10�w|��Imn�Ng5�gm9�佧`fr��L�h.�����)�� P�m�΋���K;��[\L�[��m���P��)�e�4���M/;K�oH?p�ҍ�_���I�A[e�
I2U
v�#:y�h����U^���vv�s��-y�p=��6kt����,^��Cmi�ݜ��R�y!|o*�eXR�8a���mG#}ُ����||�f��1�2���Xqj�o%�ה��ܑ�oF'�v�.<���h5�(CD�BN#"3�WZRU�JR�����x�a)���H!���f��7���m�Y7 :"a;Kr
F�E����%}�q��;�Ն��u~��|i;�	��>M����(^�f����;J��lp��}�@�q��g��=�t�F��*��f���B�f��ٴK�'66������ wO~�H�n�!f�&ΆMީ���e��2�������4T�Hͥ*�-&�kbF�:�L�/����e)��a�o ��|릹���wK�+!���T�'��8�Q+�f֗�V�<��92�B��y��/<�<�"`��퍝U�*_�䷴��D�[C����<e�,���4Ed�j����r8�TF`m����h�v����۵�v�q�77��k9�7n��lM�W�\&UBޤ!
�Vgg�j/�����֕O�<j�r����qF����m��o��c��szJ�o�nT�J� [���X5�1����2�F*,�:�3	֯9���TJWvl�j����(�t䎦�mnkx��9?h;B=�cy��9���3�1Q�Ƌfkәz�oRv�R������}�Io ��&�?3_��#�=5y%�����^i��'��a��N�;-<�5�E,c���;�>�j7ܛ�e�w]��Z0N?u���l�X#������}��K�J%�%n3(��'`�/�xF�7kh8��}N�����>Ԑ�ց�M�?��q�ujMW:N��n☁yF@�^~�p,]Ǭ��E��.1�+U���2�y�=��D�`�0�N�گ��\ә��*�B�r$�թER����z|��ϗ��C�fޢČT	��#*���;W#o�&U�H�\'�E�Z��*�s��M�f��Њ̄ygpԏ3� �J�EU?T]B�,��
<%<VM�,�&N�V�u�D{�F��-��hҒ�\N����=�{ߨ�3��!7�љt���(L5s���;tpu
�K���ޝ��uB�����]�g;����p�<�&�t���(,k�P�������g��jm�8��Z��E�)��fU��ZP���;�&e�x�|��N�K4S�(|of_Sp�)�prr�j��_�������m����ѶJ��K��>��^=W)<&�w���;.��������f�����r��;˧�'�����M�g>uU�gz��u�a+˱���mhf�v�\gfut156�c��t���^�:yR�1BR��FH�`�<�f��a�F�8������+9Q����sÛٮJ�u^��uP�� f�m�G�|��\D��-ێ�pNo�:մ[ v���s����d�'lϺ����@W	��d��2ѹm"F��յJV;�Y���+5ñ�os����v�̥���{�V��r��C�K����i��d<�$��Ƴ1���u	jw�r�z�o�t[���p�B`=�Os`fb���Դ����ى�����l�;,����6�md�pr�r��7��}^�>9C�� �
����A�@���q������ޜs�7���řB`A}��xC`p��!*�@�"0��
!(@¢2 �w�'��3$40�<�.Pq #��*���VD ��  aUf�@PB���+�f& �f&A �&�a	���a�&	�@&f	��&f&� �E�LLL�3110(�L����y���Abfbe@	�� �� !��E ��  e@	�$ @<�U�A� 0��2��2   @ʪ�ʪ�ʪ�ʪ����0  
�*�  @ȡ*�Ȱ2��8`P��D6G*��?�O��3��W�J*(�
 � ��'���~�ë_�7���r}���k��zӫ��K>uc�6���>8�Ǩ�b��+#ڞ����Q����UQ_���_��Jȟ���C�C��Xw)��������9y0�B���I����i����%�}	�;j�WpP��������!(ʈ� P���"�������� � "B��J ,���  B �  @ *� H������*�$��!�EĪ�� B H�q��M��_��'��`�"- �P �U*@׸�^B_�����J����L+����Bzv *��OK'�OV>��E����ǈ��Oèrv�5QTW$�S�>]A�y���"*����������/����~��O� 陋Q_�!,��~ ])�j�I�K|289�Pr%���UEk�c�;��?�OQTW)��-a5��7�vtOO#�19'�{��J�ԟ�4� UEx���ܪ*�����N�U��>U�C�{����̤�(w�¨�+��E.�#dO4���It��� ��9�/�?���
����d���~A[W���WfC��,�P���e5���Qp>��� ?�s2}p$z�w�J��{5B�P��*�D���J�mJ
��*QUUi�UE����T�)%Q�TBTR
)��$*H���)Id�cX���[I-�_\��T�m�[m*��)���)lkm�Zm�-�6�ն��
ڶ�E���ȵZ���kkzzr�c.�ujQ��D
�[����6M�,�SlMY�im�-��B��55�UZbM��UڛWl��͝s�mWp�v�b�m�طr[,]���kIVfj��"��.Ԗ����Պ�j��   ����zL���ݵ��umv�w�z�OGkhuw�.�ՇK{7�kAփ��U��)CE��Z���駭N�=xWw�=ݣq��r��4ޞM˰�����M�ʴ��kh�(�[�VZ�   9�(P�2$m�-ԷP�B�
(s��Q"B�cl4*�症�CCC��Ӷ��7=��.���7�]�;۵{����;�gt�7����ڡ�;���zt�nz�z�^��^�dڴ#l�y
uNɋb�Xπ   �}��ݵ4�]���[zh+��ܷ]�л40�Ǯ�+͋yQpх�v��w�ޠ�=i��Ǔ4��GI�y�ۚ�zힶ��x�s��۱���q;�z��Zk�ҭX�iVŶ�c`کZ�   G��u�z��5F���+^�{��x=]����u��6�.�=�=��C׻/t�uM.��-�[u@�k�tT�����+��\7X�ih�[Y�*�)V��l�M���   ;���ˣ6�f�ww��4�SN����V�{umΚ͛ۻR�	ƴ:�uʭn�t'N�Z�]5���Q]hP�R��f�iR����Ov��   ��h�Ǽk�;wS�!���љ���v�"�:�۱]�����@i�k�uUPR�㮨.�ݴ�km*��m�,��*�#E��  ��c1���}��+g�o	5����t:�e4 %��T����� P�i� [	���P ,@��ڳ�u�u�Q�&ke�Uo�  wx  �  ;�Ӏ 3�  �um�  q��A@ ��8 At�  �Nh� � ����� �u�[{\w`[Zzܙ�]����  �  �� Ձ� 	�8 @�/�@ {��p  �w  4���� 5� n��  wvա,��lh��-m�e����   =π P>�'( �W@��V  ��ƀ jn��Pۃ�  �� (;s  �s� _ E? 2��'�  ���)P  ��D�)F  )�CIJT   E?jR�� e*
�  f������Q?���q��?�=û��_rH�"͈ �Qm�?f����h�鯾�諭���=�y����M��1��clm����m�cm����1��M��1�q���?ǿ�?��wʒU©ݟ��Q���Xf��⣶n쥲�S�V�-̻�������SwI����^��E�����*ʍ,ie��� 7+�k-���y�٩���e�	�-v��R���̼�`�f��I�E��2�ĬJhۦ�b4�.�^IJ��q����.�-͖�څ˄�,(ӡ8Uz�ö�ßpT�����M,�ZH�Vf�`[�f�X�JGw�6���ˤ�Ӷ�����2�
��S�GWb����2D���P���n���w����I*�e5�U��{[v3��d`U	��:.*9!$1��q���y>eX�"�dk�4�9%��yv�� L��Mm6�yp��|u��ei�2�?i5�N��v�Y"���pX�R�h--�S����vʺPP�b;�؁:���!A,2��6�<�G4�m�hϧ�X �@��5y[Rɬee�xN�Tr��-�GC;�Y�(�#IT{�(Y֨Ji*�4�L�<ر�b�V�c��דs$Sj����*�a�]67r��1;��%��wup�7(]��[���T2���2�$�&�t s`2��V�I�R�)n���3)%��:OȘ���*�É�4�v�'�íԃu�D�h����Z)Ϊ\�D�ͲcrޒY��gV�����6:L[7x�c&,inSsZ�go[�.�UM���*V��yZ�">���r�t`�Y)oy ��.��hU�J��kdU�RJm!�F�Ɠ��d�7A�:�M�c�D9@.f��m;�S`�f�ҏ*�כ�V ���Bv�Ym�v�2^:�1b5D�R�EK���Ģ�����lQb���f1�ެĩ�f��DRI������ �k�oV`�ODh�u�&%h�n�How5$$�p{B	5�VMک�X%���]����bI%yn��`Y�N�Qo�t�B�Y��Q�7x&�wa,��Tݡ����31��������J5�6@�TƜ���x�����g��!���nQ�Es&�(u]�*f.�#�Օ+�A������C�7C�E�GV��JV�۸0[P�f��+n���N*��Q�9���u� 72�՜���u"�oE��zJ�VƠ�^�kvec���8l��R�b�Ɇd���t՛;2�a��S)@��/M�Lع3.��3akv�P��:�/Y����+N� �ǷvK�Bn+��7@����	R6�,Ձ&�r�$R����2�6ު���쿰G���m鳁���e�Zx�X) �X�*��6VĘ0(�����kCB��i�/FCr�KBf!�P�Xv�n�82@����*�pU�;�A ��&�ńc�o&�Өn���L�� �Q@^YY��YR��DV�$����a3:MZ���6�e�w��e]���A�p�n�'�^G��qV�%������kM�7Z�.XT�<��
�Ue
Y��v*�eQT�
-Y7r^�D�{M�(`���MLR��ȁm,�N��aa��.�C0z�w��GN9�'"�[�JŨ��Җ�r�4tk6�4m���f(�8��ʼ�v�3x�
� ۑ��7c��(G7��-m�th�K t�A���R��SC�l6��!V�T��Ğ��i��f�/+od���c
� F��Z��T$�-n�B�b�5n5k4�R:��h��`5�-�Fm��En�n�Tr2���IM[.�⬼��6����U�pB+R�d�;ڋq���QI<ܠPX���1+*'�T��]�Ǖ�e�[�o���(�Cv�bE�A��WW��r:v���J�,�$`ތT�D�4j���A��x��ti%6���]+:Ptq��Ӭ�#R�&��z�,��U��ة��l���T����nRS\6�v�ù�J��f*g��;�Ŝ�*b���1nAJۚ�`#]�gR�7q�z΃�DP8ތ����wR4�'s348�z��ì�J�6��Q�)�w�:o׏��tq-v����Z�H��q��)��`4�CK��Z�I	ML��]�PϦC��� ���n1E�$r��u�/盈V���b`�6�*19����v�ƅ�ۄ�Y���-�t�vi��aj��#h֕uͫ���st�#�g@�(ӫ̽FfVX*+���\��`iQ�S͹q���:^�Y�CB�&A.�1Z��(�KyNnˢN�n�V2�7�Z>λi�P���6R��YvN=���	��ܫg5T��6��u���jV�*iBl�F��M��ZPTo\Me<�@8+7b���������b�5��+���bY��m��H�@w��-<X.�b�Y��Q��*�[YH$UC,`7��,�����P-;�b*iĒ��=k���T�y(���5a�@�Jd��S5��Ϯݔ�JȬ�e4p��Oʠl��sU�ksD�غP���ÏT��C�݂�����k�]��y.ں����
pL�[�f��f�Vι�o-Jq4V���Nn�³a�t��0|I2d�I��^޺��P�d]j�"3M!b�r-޶��J��Uk.�7$V��g(�����sb<G7"�ԑ����-�K*GjQ�!�(:���`��ir;��5d�ȩ�,m��a[J\�	۰�R���M"�9�Ͱ%2��{B��a'tm8�;����5Gh��Y2����[F1!�Y�	N� l�x^�� ��(��m�q�o+^�(�{�F;�t�	b4Zr<�6�@eLD2�P@�������M�wn�oV�.�ͅm+b���F�/I�$��Nج�zŌ�.≠� Ńm�D�@L݀%�G*|�#%����ȞZI�e�DbX����F��#h'Zn��J�Ab�]PB�ǖTwL6�c���;��t��a�V�V��V��k#�Õ��h�s&E��F��Q<�Z��a�)m�VUm�v˘E�ugײ,�SX�p1�*ʭ���"*T���U���&�:o-�p�xҳZ�4�{	XX�~T"����CCn无eh�P	m��U�:E���ʷ���u�Ba0�J[X�md[�*�Ρ�ѯ0�	���ZW�O���,Cy�b@���,ϲʍ�U�:����1�y�[�'uD�e��]�-���V�{5�ԩ�wF�K�v�t��4��J����ݭN�i��9V�H�q]�\��+����.c��=��}�[Z(ְ��L�2��ť�)�(�{�,�w&����H��f��@ɦ�BK�g+M�ť6fJr�b
h��c~�),����"�U]������F�S[s�^��Cwt-]mϵ�,����u)�1� �`S6�l�j���E*�`;d�Ȍ���@ʔ�
q�,�X3u�5��l����2�v6�0���Of������@��p���j+�LeK���'�[V�u�^���\����P�Qdh�ɛZA˔�F<cb�/JH���Ypw�X�b���䩇�V�R��0ZK\u)��U�;d�v�)�p���:�:��J�,5(n^�\ڬ7���nC��!S)�0�B��%�L����={��CP�kj󵷅���X�	�%�C!3k3t+B�x�d�^X�@i�G$ش�׏E �*�b����}��B����u�*ʣt#6� Sxs~�5Q�ë(%�u�\)1��� #�A�S2��)�S�9@;l�9�LħM��3V��)^��n�1��(&�Ͷ���.ɚ�G�wU0[CRE*
F�)D�Ĥ�����`w0|5���ߊuu�,�a 5�2a0ϤA��5OfUک�W���sqm:"���V�CZ���zK�Y�N锔�����a>2�B�%��=���,Fӎ��N�oH�,���z�E��v�ₔmau�<�D���4��R�TձDF^0�O$�*��5�	���Xǆ�lçhJC�c�(�(PvV7%]�n;&�S"t�i�X\�]'�2��`i�Uw���$Zu��P�_S1�w[Z6�DM5�E�%Z�����kf�V�C�m�z9�5j]���;]4��Д�Z� E=�㼂��k7H����aВ8�hӄ�k5���zP����fA���i��3n�[1J�켘Ecq�lT/,v�JT�R�WJ��0��l��X�&��O�B��y�q]K��G�X�b`ʹ)n6��׵ov�dt�ݝ'6���vɘ�Y��IІ�K ,�v(E�J��:�y[���L'+EK*��!f1���%&)p��uc���yγ2�v��Z4�6�
���>s)�]қԐ[�E���'��-�P���-K�$�+s3U��BH�a��*�/)��ibl%��*�ô-Y�[��L��@^]�2��:�T�z����P�{�1�	J��J�(��MJnVVYw�"��IVP^Z[UJK
��Ļ��˫� �)S�j���!�[����ǵqL�V�;b��A
�5���&enj�d��N`$�_X B[m�3�t�F 	Y��<U�e1p�S9�RTP�2�k�D�]��h�oe*:�]��q�+M[�ݻ
����D���NWm}깄+��pS�s3)�L�R�$�r�`�����j���ɲ�u��xɨ�����p�aI������.^�[hH�A��3m���`X6�RG�+��|�$JJ`�svܤ��:����;���i#n���Lq�.�A�tF��m 3,��j�Ѭ�Ѻ�Io0�h��ڴ�)r�Fнg��e�b�%�y��� ���Õ4

SE�D�X�.퓤���ldغi�K%���v�QݴĆ,#+ ��J��-'�e档7-j�t5M��?�U)`˹p��6�Ǚ�@ŷ[�X��*�F��X���Gp��4.��rKʳ�Vsv�Y��m��1m��6���2^���e�(&�L)�ʰ�I+e��i�ܡ%5�㫗�u�7��Fc4pf�30	��	 �E]B��&еy[5�H�rɓ*rnj�Pn�$��[����:2CKv�Z�Њ���%c�D��XN��*����(�[����m5*<�MǛڍ-��7��j�^f�觏q��XtT� ]��F(� �.���gN�c��7-{��sZ��.%��0B�����b��,b�b]jB�k/(f��@�h�سKV^��flʣ-	blhD�Ya�j�F坢���n�����(b�m���i�*eYf4)�/�h��|sAXi�iꅹ��,��^���N��Y�E��?c
w�]h
La�!\���+.�^*e�G��D�=�8�F�$�N,uv��W��X��V����u�3u㶍"ܓ	��&D^�h�"����*CV�#>xI@H���i���[6F�$-�?K�-�2�^���]$&&�N;ƶ���t&�dT�b)�	ީ�%-�Ze�
8��k�����;l�¦�9�InowEs�:Еȥ�l؂�4[�܊�d�O�4�/dR�d2��v�]e�" n�'s@d�ȱ��`�]�n�+�2�Ր��k$��#GM��Xn�2K���K�bݽu�4hY��f���M�JTY{�N$�ʺl�52��̡R����*[y�U��,��ԩ[xv��E-`Z\��t\�x�;��9fb4�-ѵS�Z*�Ƌ���k{�����]
�Z�X�j<Y�C�HS�x�n�q�;����Y���cK()V,�9M(�Ȁ�c-��Ik#.,�MG���ɥ�!��X�Mb��B�-�C%�nϦ�t�m���2e+f�ob������Ҡ�FU�Q�<�t�7�00GF60�,�Ͱ��|T5�Fd��53���]��V�-�L�ں˩�����"�� hcݺ�Mi�-\H�د.m�at����b����xL�B��Y-٣y�.#5�0=����U�Jh�i�	2Xȯj�KC� ��b�f��7N�hM�h³\�9C-�����Xʕ�R�����Y#�6��Kv���)�*�q"������dS���0-�Փ=��"�iP�c���pEb���8Z�yn�:���M67YC7V;����ʉG���d;y�6���{�T:�OlZ�!�ɂ��2�ӌ��� �cv ��h@l�A�^�qͻ�x�8�}���ĬnR��1hQ(����@-�+^f��������Ѵ��ͤ$Ǹ��ݒTf$���h\ӹJ��GZ�*���0n�Z3�դV���H+�5���!����'�^� ݖ�Z�!DS��2ҟeI�!n��SAb�Ab���`	�͗S�q�pVXµ�{L
��,�ܸr�C1mAR�jm�0��Q؜���j�-aI�+)��ZwoCZ�(���FX�:5�5&e�G��:ެ����w1����yof��(։�l��}��P�Y���됃,�*�]IG&f�p�a��Y�E:�,\Ƣ������V<(�B�m^��K�1��(J̖�<u*����ˎ�ԑ���	���մ��.A��%K���+��͘�K`�d��u�-���,,��Tr���MGV�%	�3o2'J4�g6���i"�9�-;�nG��
a��P��v;uqf|NM�`EO�xjy��'r��t- �Y��SX���6\'[�
m��h��BM7��M�%�ĩ��4�+����K3�t!ISV/@�Ȏ�bn�V�c��F�t�J�����Hhv1Zۥ�*�-"G�)ܣe���E.��;X�Sg`�$l��TPMS�"٪��I�RXS�Kci#������嫛�!(b�ⳛe=�)J����[��\G^�%"\SmnJpE�)ӳ�b���3ս8I�i�}�Ӄ���K��s��8�IR��(�B(�nc���2�m=���֯,k���PH��C��
��X�9�zd��u-����q���zhuw��gl�N<��
R�Rv����]�_j-�/$�gZ��v�6W���hvP���LH��/]�[	��N�7���#�R���5yC8���S,��Rq9[���:��%�����%]]�%��ٷڜ#:\l���Yy�Q��sZ�7�Vc�T6��J�J�+=|�_]*���9S�ɢ
����V�=�<�R�Ɓ���"u4��td�=v{`멏��@���n�⻧�i�wڝ:�VP�J��B*}ϤؾC��p
�mf6R-��L�z��B[����;�Vc�j�!�X��S\榓�i%4������H�ݛ��nQ8��u�����o5��}��s��b�X�f����]G�k�ݗ,����N����pѥc;�.aY�]O#�����n1
pj҅u�b��?{��-���%��l�I����i�`m�r�m+����ˉSk�=dt���6GgIҞJE�S+�`˧�<ڝ}�O$�%e ���Ȗ:�u��rª�:HP���#V�Ҳ�b-����R�ԏG�����O@z�;B[Y���\HKK:f6%�U/T��#��-�ƣ�x��C�M�V�4�H��1k+nũ���h4]�@��+�S��9�n"�I1F��N�h�C���Nh]w���XT9.��C��
�M{W�b�lN]\�0�m)����2�NP���Ι�<i%��z�Xβ0����!�}���W`��G\��ͼ�L�|�����./�. �u]MT��c��Q�Φ�Z��宦Hn�n<|#Տ�IsED��M���ǒ��k�&��u�o]�s�n����pW\H�i�d�;z���U�ɼ���7�VL�GV�p��h��#1��ֆ�� '�%��i��%�4�ZJ]��2�r��;�h�M5�iW`�1ٮ��A#W�`�x�ls��ӆ�	c�'����S�M̦�|,C�\%�J��n�(�*.�yU����h����r��U��/xŵ*��
��[e��ʵC�..�A�s4�:v���O�`���+ҟU���Wd�{c��͎�`�ށ8���sΎ�ٹ��y�U�ѻ砶$�\�m�)x������)<��kOh�� �vE�g�tݑr�T���U1�-�^ˍ>};� V%�ЇI���O/8��9��Hk�L���Q6�pp�%@e,�O�5�F�� ���j���B�`����0��SQ��՗\++r�d�D8�Ej6�Պ�5�y��L�v�Ά&�*aZ9���h�,b�j��|ΠO;�D��a��WJ�����	�7~0I�H�[*�n*;�gRے�a	�2�����M}.��q�pYHNuke0�Xj���U��7I��He���掻[f����$*G��֔*�J���tɜ�䝭GR�z+`�C��&��8R�/;3��Y��&��r5/*�!v�����W�u;Xm�]R��t;䁏+5F3+/�Q��{W�����$�Ͱ@�X7�Bt��18�-��:��̋&I���4i�I�0P��f �:} 64�Ž-,:�ni�]QobL5�`��{Q��o0�K�Zx)�r���y �W۴;j>�W�Ԁ�K�.muѷ���� 7	���f�\$��� �WaKq��9�
�6��P�-J����W��ek�7Ӗ�i�4l�a���ͦ%\�s4J��w��t���$*�ls�.qEk��{g6�]b���]NT}�]�_$xn2��"�g@�&8�9Wx:Hs!.�㕗�,��Ջ*�
w�+�����V�h��Q�w����EG�G�i>ذ�.OaAZs��SY���L�2��BF]IM@HZ��Ma<��Y����C�R�Aݺ��18�2���p:�}$���M��9�A{\e>^waS@n'����L�������wP.G�5w��qZ�[�"Y��Ú��R{�*7On�)��=W�]]W�V'O�}��`f�|5)'�6�T�1f���I3n�u��]�C�=N���m[���Y�Jա��lF<E��'K�闧um'NR�ҮR4�9ΏsUmS.F��[��g.�¢���%V7��pPf]Z����\W�Ү�%k�K�YʒĂg�A����%㕷�C4P�g�m^��o�K�&V�=կi�Һ�^u�������Bk�6���1,o��
_qq�㝐uh{H�\�f"��.��sBp�ϸ���+5Ρweᢸ��ľ��Z��]���mYb�t�9�KE�^8S���H�����s���1d�=��Q(����NY��r�,,��'f][l����@�uڠ+))إ'o�ݩ&�
K2��Ў�.����O�]�\��kh%s�YI�L�gjނ�5����-��E��9Z�ʒ(��3j��ta�]�䕋m�:]HǱ㴎ffX�ի\^�S�p�rGea⛢������6<�D���*��]�&��sq�i�]Xo��5>�wwb�x�9�_Ϡ�0�Y��S�ua�[Vr��؏AhQu^���ݾ#cHC���VH(̝79��.�ʔa�_,���	v�V�
�+
��d�b�I܂��������j5��ݸ�՞�g�-���-]�6���T��ޓ�/E?�V5R���b�n��'�Q���m��*Q;3���b�����'�,py��fM�>�w9�%��=����N��n_���c5��t��JMP��'twR�18��ue�.=��3f�;�P5-]��	oj�0��oU�ݷ�j={�;mғ�R�\��zP7.6�Y�3nۻ���£j�:�����E�S�b�2ig��Y#�y�Q9;���C/����IOjm^`�ϊ��>��ӥ�R��ӱ��l 0b}�*�:]������R3P[��W������J��]�.ׇ-yki0�!ΚV�[ܺ�vQ|P����@�⵴5�y$'�_:U�:�Μ�s��0Wshk ��JZ��3[��6��K#�\�B[<AS4p�;Cm-��Ȝ֊{4ʵdFY9��T���t��բ�Dv�����#m�^��z�u��b��w5�}�G�խ\y�έ��Cv�s�F�ܬ�B���e1
J�0	L��O�N�O��Z�2�t�	���ǵi�v��u��ۮO��}_a���+�[oE��fL�pT���:�Xu��b*`:��k�S �-ゑ�ס�	+3mU˂rK �j����W��.K"n����h�)�ciEu\C�SX&hb�u�7z\9���L�ݒYhk��Z\/��]r�)�i�����j�B�V���[*�������_tY�8�9�'qq+����z�}q�p���U�_آ8�{��P�9f��1J58:�<>��Gj�}YS��l������HD�]�:�٣"��YG�бvA`�+S~�6��B��yu�*V3(Ҍ���9sk
˛c�����v$EZW!��+xc�4�����$bq'�5�ʈY�2����t�]�
g��< _m������Ϋ[*�;u��%α4>��N�'%2�S:%vp�.2��P3m����*ˎ���r|�͋[F�b�ѽ;6�_Iϯ]	Hw�㠌ꑼ�aa܋��Mk����W:R��>2p��a�ô�f��w�&��� ��ŝ�u4�1�WJ7J�k+�+��팄gG42�\_%��̘�X��k̭�1s�G�iZ����I��l�:�L��'�@��ȳy�]]E�J��n���-������LWe�l�*�);+9��Y((�ٝL�ڙ�F�Z��EF��et-|/{~�Zݡ̳c/N��%�\ۨ6�.�r�jx�3��]�x����^J��%Ȯr��Z��TQ��>h���|Z�;��X��)(�:7�[����J���]ݔh����(zi�Я�LKڜ��5�{bp�lh|'0
֬
J:��5囗�i���0�@�(%����jP�Y٬�!�$��������[���@�JR�Z�:�W}���u�G�Y�� ̬�j^me������mP�.�96fhX{z���
-N�-�w*d��y8�l�;��̈.q�X+,h�R]\�����V}�Rux"U�E)��f��.�X��;y�=7,u��G% *R��
㥦�w8�]#K;k;ih��+�Q�zrV~<����9�+������o��9�%���ucg����p®/��nC��^$5���dDnv-��n�8*t� |�wV��=	yWiʭ kK�L-��i�һH�u�`��V�Y�2:R�T���ٮ���[��\�D�&�mk�I���k��;�,���ͳ��!.�\�q�۽\8�E>��[[�3�t9��彀�b�	f�k]���]�a�b��Mӥ+VY���M\��8V�r:�`��o ���V�	��

1��Y�+o���5�NPo��NS��}�����K:�x(1v+��v.�,�g)7k3�쎁���Q���*7w̮::�=�=��fJ�m�\��Eyx*Ay/.V^�Ɏ*ѫ�\�gG��;�n5/u�l����,V.�|��M�x�Ŧ�T����RR��%��J<ڼ���v:ҕ��:�&3,����iW).�$�$D����H6�Q����*l�I�`��,�l.�e��+N�W��5.�C� 8D�a>��H@�:S���a�{"ĕ9SX��~�L��0��vU�_]�����}�e(�Hl�T:�%Xr�׮�2��V���֊������v�Ć����QT3��R�m�2m\e��JJ")����c�N�Oӱ��a"��@�̹Y��i����W$8KԣC�ց����z��I\.��4_|���o8��QGC���!1ɐBJ��v.��b�WGl�Z��Y`���J������M���V.��#צ޻o띗�MՋN����&��w٤�����q����_��i�6��;��`�N���[o2R=Z]+XV�5Gn�v��m����e#��([����5//�`]�bY�ab���R���f�Z{OyD�eL�ו̫8�d\5����
b�رbv��[0�n]���8j7�w���n�&.i1^�V�����=���ӈ�8(Ӑ'x@���W@M��J�z�[h��\�Y���C]Xu���ঌ�viơ�W��$\�B���lzV�K'�G+ݬ��aOF��.=������p�Evt7�/�8U��Ӧ�\�0ӹM��������=��@4�Vg��ev��L�V>��g6à�# �٥��G��m\ʛ��w�5ga��JU�@���|'P����J�dg^�i��ؑ�6���@�t�v�)Ԁ
�����]���}�kÏ|vR͖JyN���.k���g�.1����^_=�|�-աx�P��ų���fA���X��� ��tIh��<;��mi�s7n�QO6����������dZNĺ�/��ob�j����ހ�eZ����#h5o7���>Yv�U6M�$�:�5�X=��+��L�os�۝}*�ϱ��б�B�9�Ů���3����LޙA�z�3�C�-�n�D��P��X���U嚌F���d��\եm`v��Hn�9 ~�z����涹�y&o��B�Qո��EKk�`5k�|B��t��1��+���VPã�^�Մu�"�������S�)$(��y��qSF�4�v-�[�f=�\{~��J���	�}9�[𤰖�	K���V��ClC|ogG1�^ݛ��ka��ki,���(��.֎��0���vwr�;v�^=! �u޽���pj*yP�t%`��Ӯ����B����y[��ƙ.�BW�eţZnP��$�U����da�/�-8]ݴ�v�$�f4ťb�gR2�>͗\����Ops�UTf!V�K�r`��y|B�]���oj�ysDYx(N�M�*���0v3���0�O�9ڀ*�]�36��h����f�`
�_*)�L\X�/6;/wf:G:�f�6 f�`k��`��nY}�>��X�� �7rϘ�t:˄���$*��j
��Ԍ%���7dg�B����� ���5K�0���̭�ڧ.��Z�n��5�,��W�����r��t�����L�d�ƴJd�J�p�e�{����V�s�]%���e:�������gedjI;�j�[���ْ��8׼u�v{��t)[Y;NT�X�9+(V��\	J8��O��p����5��U7�7�gm���6�*u˹���K�� ��#P�Mn�:�V.���h�J�/+T�h��L83'<��{ ;:�IDAo�'Vu�#�c�hj��PZ �lW%��v�����kA�}��t�)�l^^�]�rǉi&?�����ڶ8Ց�<RQxU��+��Ն�f��)p�Hi�(:��W�$:A����H3�V�u�]J��2IV��|���댣���,Ca�y�-�nՕ�-���!�Tz���0[�,�N��:^����ᗦdR%ɺz���^X��Qǩ^G1	�L<�n����^o.Opӵi531u��� ;#�*Q{�)X�[��瓂�Rr<mn���Dɏ���m����t�:�%Y{��RL�j�'��
R�p����|�n���]�ۭ�閙T��wE��[���+)�l�� �.�v
� �R�L�b^Sy�J4�޼K�G�:�W�d�ۀe8��Oo7[y��/���ٍ�]��i[<Tt�i���^����	���[��i�[�{I��9�Zk3xu������R��Fԫ5���ƀ]�]��r׻�׍��Ie �#�u#�q�� ���vܨ���u��U� f$�fS���Y���l�D�cM����w9�W�}�}��W�G����菣����5?e�¥�VF���Ip<�M�!&�ǝ�0���!�|�YgHZ˓E|0Ւ<ڍ���C��0�V���h�*76.�KqX�(Mu�-57������Gӛܢ�=��E�t���B�b�*[���X�O]n���b�,W;w���9!ʠ
峡Zt�vFs�*%6��Ix�z�ڗ�X�Q3�4W.�B�NG�V��1��)]�b�l����̰��]��k:�au��{�>[cp���Rb�m_%��Wi
����YzY��e=R�����M��g1����X��@��u�cr�v�mY��n������)���J`�us��3�J�U�*��b��X��Õ���R0ᗧ����*�]�콜�Sm������l�3���n�Ë�1s��wݪ�f�$����E�/4�����Ie�2B�+]�w#ٌ�=c�V\�ֺ�l%R���t�ʻ`'���MyRNZ7�7q���8����(�@����I�>��|:U��nni�>V�m}�pe{9��+�ָ�Xh�mm%E���2i��
���wn���Pq�S�1;�Lr%*�6��w\{���@��lu����
w�H��[h�(qV��L�<z�q�mޚ�}�W�2fM�opj^W5C�L.�6�R�R�n��`��n$Qt+eegS˸6��������&d�j�{|�;��akk!β]��R�H۝�;Yʅ��/jZ)#�9,S��B�L�h��Ϧ$��ZŽ�#g�Q;�\Kl�M�aߜ���/����PJ�j���ٌ��v.`a6m�3i�1GR�Ok[�w
�˂՞�٪�1(�˷j�j�''�;�f�W�r]���E�.�C����X��t�ۋ���sZ$���N>�&Ҵ�Ǖ6���Y����gS�\ʙ�>�����ff��:]��T���7�O��V�!�_!%��D��}���=�]�CC��G�A�����+�
k��t��M��_"��H�B���e�ķR�!-���'B�YSuw�evkj r��K�7��jv剕��]��2]�)��B�ŻS+&w
JK�٢.�y�,u
ꂆc���5�i����U}u�T��=R�u�W�jR�tS����/c�-��5�xI�J2�`�5�#1/�+��{S��P�Wh�Xf�]�X�c+u��Z�l��5�S��sn��DZf�������b�:��s�F̕�����e��}a+�r..���:]ں.��[��gU=k���im�JР.��$)du{���[�P�:������%j������!����F�b�U�VɈ�j4C�]����K4�`�;�&��.��Fee,wU����l�K��
�5]���ܨ^�VU�D���1�;M_j�ta�Z�kpbz�ʷu�9�|�u(=W-��7����>!!�O��7tw�rM��r��vI�1K9V�ĻQ�X�;.Eyj�]�%�Z�l���Ť��y�oTƸ�n�l�U#�/M�Fk�|T����ۅK�Gx�G�t�rp�4�bh��{F�X��m��ۏRk.Ƽ7�&>�7���rը�3o�"��ù�Ion�m-�@��	������5< �����_�5f�uZ(�:z.{x�;o�&f5w2p�Q���-p�Mht7v�U�'B`0;�>����Dl���55Zn�ҝu+DnkF%�V�g1gn�V#�T�Ig��v���D��-�ɷl��^>�P�+�d΍����q���RMi����Z��w�r�)쏃�/�� ���3��91�������B�
��v�k.H��7�G��)�ֳ��B��bN.G:�x�qq]Y�kd�
Z��Z���@S������E�㽫��3Sv^g��u��L�.^���A�+OnR���)�P�Y�y�I���b�tVڣC��'��7|',2�Z�殀�J�m,�T̫�]����'�3�r��r�2n
#�Ɋ��Ȅ�b<îή�̆�5���v(>͊�V�;uj���#s�Ȓ����&����kw�"f6�)51ح֣��"�h�J�.U"Jt[�-�9�')J�1����µ�ϰw+C��a.8{,�m,J�`��MC�ELP�z����2ƹ�`�|6e�	>�g���H�R��G-� '9<�]e�z�; h��(.K�f3�2�tV,��gZ,A�Q�vrQ�/G��bC�s+Q)�X��`)L�6F	�,E���sU���V�U�w6�z�CT��k{/�)�BV�u���
����ӄ�eᮕ2/���#븀,��j�ۨ���V]A%aX���z�JK~"@p�>�y@�*��!���΢�>,;�,����v%�����jRX#��%L���z���`��<���\�;N�*���xe��E�J=�n��@<�����3jw@�\�4��VMy��B�2�<I��B�:c�^���ے�h�����p@��x�bā� ��k�F��k�eg6E���Xm3m�`4+R��4a��a5�4*v<N��v��vK��U��'(�Z�� ӭE�9ʗ(n@��=ȺLξkS�M�Ԁ�VS�fӺ!�C�F3%2�q��C�� ��F)8Y��=��Ĳ��S[�Kv�ʽ�1��q^�р�3V�;\�����9����Mr���ǈ��n�;펤�h�����P#k�㒤��:��2�BV��ewn�N��S h�S* /��F��j��[�MA hT��Km���\�WB��rK�T���bcy�����Z	5��B,��ݜ8nA;/h<�t�[�[]i�03��n�j����b�+�M�9��T�l}�D/z�c��h:-�>g��}�ؗǺ��c�a�ǫ�Thl����]/��Q����`�Ln��m��s��X-�I����O@!��@�cA2�:5�]�f�Y���wx��,n�J�<j�N��j�h����j��BȥZ�+:��i5jܺĪ�d�m+�qJ�~���vFA=���Tu�4Թav�x�-Ib���q�e��x6��^v&�j��k�U��-��D��u%�GUe�&�b��"��=E*��5H��G�H�m���;l<�:at�E��9��5�jw+uD�]�y!	i��-$.�\��6No\K^�9��������Zo8�i��%jp�ɹm]�95���o&�*t���T�]�*�&�k��A6Y\2NmV�Z�̻I�4�{����3]"ڵ�D�<Jt��;�כn�
�7�@����L��kY�)f��p��K��f��I`9{�0��iCk�hѡW�S���ʝ��2WS���O��$m����2�<��:*qN]�+�s�Cfv\�wo-�(>E�7U���h��[�ʒ-���3==w-�J�NF?��&��ZGqZ�����kY�(F"P+HX2 ��/���Շe�^��ʻvWq�M8�5N��}uoE�7�V�U� v#�Ld�Bp�Qn��MQ�s�s5� ��
��t_><	��fS���y�k�pqX'��WV��uMw3�����q�N3��v�i�@b�".i&1n����т���iA���kH]6f�J�$N�[�� �P[�x�#�����+�\E�K7�S�"�m 1D:r�Y������:�PY�l7I�Y��N��-���wu,���{����/�\���^�������2�bj:$�r��Դdg�	:�9]�fs�%E�-�Y�*u�T"��^��P*:�q䷹k���edU�g��D�����cǘ��9b�5��]lJ��;ԯP.NJC�vb�/�J�6 [��[̔N1��9��O7;��C\]���CYѵ���7�]u�:��*4�[��9�s�Z:
�z�a�˳�T��D4ӳ������NQi�j6q뾹�%�%�%C�Z���{��)����N����c�-��ٓP�u�J��[��╴�����=3\M\����rY���3�Uݐ m-��"$9��EK hF�S��42�S˽�:�#1إ��V��ʙzl,-0�]j��e��|�X�M�*N���Eu;5��Y���dfi���iY����Y'fHF��e�����*�协�N��C�~�f>����6�C@�ѥx�;n�V:�[h�\�\������[ɝ֘l������鸧>��A��L�|��o��tBh����$�������Y�7')��\`�yw4���m�-QAo���۔��7vX���VƎ���"{�"�av����t����g)X�K�m.Z�Tu��+{C�uY��H����)�N�"%�%kUz�ON���<�m2+++���f�cF-d�֞�$9S�����	S��$v�O+LϢ��V�F�]�cH<�q�ٌA4*t���ڀ�598���i��j��i�)�.f����R��S�Y��5fli�6B��V��A��*�d��=�+�!-}N�7�;��&
�c�=oz�����7.�V���!��p�S��٩7S��4
�ܨ���U�лg
���
���M�Cz���T��/����@; �(@�+&G�%&�;-;��K��X�zjZ]Nho��1��<q�{����+�%>�:������sz��u &3�O�;����a�*����]�����Ť"�����k����u��j���9'��E,wopڶ

��[�����97�'a˦�[�Z��t:M͜��Ї@ż���(��"�Ǳ�&8�[��u�qr�˖�"�&S�K��_C:2A!$��Nm=훬G�.]�.��P�y�Gn�ud�v|ҝ-��7kr�*�N�SY+�����s�V���8W���rĤؐb�G�뾽��qF�d��pD��>�ޒyKP�-�t�߮COy��GF��Rh
mM&��q�(v�n�����s�b�'���Pݢ�-�Zs��˄�)�i�ww�n;�t�e��|H,��Sy�x����6d�d�S]�;��"�t�"�
�e��zn��P�o��#��϶������&S�(�初�/A��w�;JXC
����+���O"U��}e��Ty���,�ty�<��G[�y�׵���x^ r��I�uvd�c���2v����X��ݚ�[�5Y��i]�i�\K�O�\�sPV��Fۼ��q]t{I$���t�wK�y���󄰍:�����o,�{�7rM�B�w[�n�g>�aZ��J��&���"-󓔜.��nHCU#���i������S��Է��r8�tv"���bwo��r���%O��W�.ZRJ �9z�hqK����t�H��|�.N� xnC��ۏB֘�΍�|�.�α���Ů��������7*'��$��0R����7�A�6{��/��R(ua��+�k_Nī%�5���V+HZ���.F�v����x���̪x8��Ca���{p�)fA��x�f@�X�Vd��P���X2��|�a�y�z�B]Đ����e �F�cV�y��Ѽ�*���o0*S�`]������I��'O)¦����=��4�.��l�Q�-Z�^9���8Rg�	K��,�K�ht��gr��̂�W@�e�7�������B�����R�W���ޢz�*z���0��m7����N�ޡű�Vм6�j�%� ����M���ܒAl3���#��Zk:*й�Ɩ]����5��Hz`:��.���Z���fc�]"�u>��]�?6�O�\�")hc9Ү�t(-����|Z^��
�] ��gk3GYKt	]J��>ݻp�kqR���t �����`T�w��P�}�'u�wY�8ӡ��>L�x��9�v~����;X"��wQ��=dY�ҙ�ٙJ1=얶]�ӥR�@u��/��v�29��.�Х�����p�f���r��W,��A������k��u&)�]�α:����K&�b�<�<���Z��(^3c^���*�s^�AޅHe���:�����iE]l�_H��v������O9L ���A�a�ڔT����n��%��h8/g�N�K�Txm��<a-��JY��X�#k��lR򯺥t%7+^��3,��8��;u �\d�&�y%��f�k/�g����3�ۗY}X����S$$Ղ'Q�oi�o��)3��^�;�Myu��D8[��\�o��
Ynmdc�^i�\��n�](��3*:�Fr

g��Cr���}�M"����oIN���Rf���ua�Î��Ui�[�X���"��^N�lB��yp���Y��R�V�����nNz*0�϶-�ͺ(F�ś�Ϲ��0&i����M9bKRť�/��G�+ܭWN��o:Ȳ�q��ń�f���Ne�Y*�.5��.e_m��р�s�R�:!iO2��(d}l��c��B"��l����[�V��yܑ-K���
�;�m,�.�{q�
h���4����K����F�jY��Q4tun��;]�87V� ��66#R�\ױ`I�6$#c]�`���Dt��Lײr��oUf��l1�u����hx$�H�f�7�4T	H��=�R_�p�z፫���r�}��-�Wb�5��NFL�lb��'%mЖ�!�]v��\���-�8���ZI]����ecu��Ӿ��Y"`�4��*�*s/Mj4��Xӟ$�W��<��A<̢2��V�Ԥ��9��&����\�!Gi��J�t{�-���X�τ|V�Ա�h�Ux�̆��ƺR\��,���v�W���^���y��ݵ��xU�x1hb�(:���������A���*�gm[�N� D�'FYM;��0�ǀ�
�����<��9�H��v���_��S/�g����������v������\�	�e�]޻5�
���}����ڜ�E8M�1\�Mm1ol���*���V9��嘜W]��E�a$'{[$&��+�㿕qT$'XT��"]�1�.�Z�����k�9db�b�.���D���^��K@�G_��̡�^3,��ؽȫg'�ړSr��C-�mm	��%#FwfT�p���ֆ�B���k�+���Q���#�KV�e�;$�=O�S&:��H��q�YėztT�Nn��c��w*�\s��T���E:BAլ3��krZ�{m񪢥���"�N��6�4e�;	Z�ѽےL���W��xm�4kN�A�X�e	 �rB��ғ�N�)Z��\[}��T� ���"�@T��m��� �C8m��*���oGB�`R��f�l�>�fK�0�T�|�\knҤl��ً�#����#��_ZHv�-J�[/.Ԇ��U�N��Db�G7���Ut�!��<�з�]6��E��ޥ"�b�K�"�	Z_�m���bo�xc8Y�:��Դu���Vw�R'x�^�a�̴��I��Y��:�{���łe�	9x���S���z��N��D�.��h��)��m��*��;PγG��F�����,�Fs���gL�͙�U��5 ��LjQQ��2�ڕ��c�2�����+�y���Q`2��PĎ�o���T��l*�V�>�A&��wTẢE�<�
Q�$�Q8mP�[��D+�Ws	�1B$P�MDMd�����P-DȻ7W)Ti릝2*���MT�΅�t����h��d�+n���2��Ua����]�A�0�=�皡]�W(��䈩VD�F�eyIX��j�E����(,T4K�9�N�QPW�sջe!{��4�AL ��%ii%��㇂�AZ�X ����3I��r=�T��"ê�4Z�L���"$D��N�
%f�$�����d�Xs1�sK)*�2�MT30��憖�n�D�Ct�ڢU��F�DwqB�1�JʔL�h�Q,�i��H�"�s�j�Fʣ���wD�C��t��'q�<�3$���)��S#2#F�����hherB�"��l�f�^�+��0�Ҷj��y^NiO[y�NJ��ʽ��p����R;x{78�H���:)�f�֖,�8���]�3���Yt�\�.H$�nm.OZV~�<�2��	����&�w�.�5}���}�LW9�R�yb�*�4l��6h�k�_1� "��h0��%߉x����$w�}
�k��m�Y)��\>��wJ�����y���`!}L���J���[yAg^���s�o�.���¢ἣuʽY�����s�t�/���B���.#���٩��ڌҾdZ,�фeDףNz&\�&�=��-�u+{��6��Ձ� ��۹�\0�uN�ϝN��	Վ�u��U���+��w,|���76\>p��l����/�0����i��;�[�l�+��M�y\�W9��w��˥�Ϧ�ΗY-ٟ�L�Abx�ժ�K8���D����O)�X`+�Kc�|ô�轑�9��mL�˖I�G3�U}Rkб��rs����H�V�t^�Iy��og�\�\&b�*cr.tu} �1<P$�}2�����0��t�Gl)ab�%ҟ���R),_˱#�,x����V��@���,��� �����q��a��{X���I��NSθ���f#LM��¥@�j�
a�%ϲ�o��t]��1�RbR�q�^�҉��*�;eq9sb�|�g�MG�;�]gA��\N��C6Gӷ�tx�@�����l*{r>�㙵����x�vJ\e𩕅�n��9;X�G{�.Ӹ~p�V��M�Ƌg����H�9e�/��W
�A��PN6��~+/O9˧>�r���D��]��ҡ-�ʮN�h�m_�졹���q7��0Y�2�ޙ�{=��Ξ��(9บ_)Ϩ����vuArj���"~b�'}iz���r���\�]��ʰ��T���;$��9�\�z�+���Z5�Ó��l���6i���sT?��j��V��rO>�B~(��G�����B�w;Da��ei��P ���b���K�$R��M����b�:a�f
߇��mL?�̶�,S.zU����U�����Z�.N��/�O�M}mu���>°�4UB�t�q�k��,�gE�Qp������vN�R�3���401qΟdf�AY���o�k1*A�#�]K����Ȱ"�Ϸ!�m�Lv�b3:�K/�^d��NBu������꫃�}(�M�P��k��ﭴ��.'v��,����V���x;$M%7�د�a���d����QZ���!	�e���x���X̳!�T�DЗ�e�qF=�|�	�TDG����������	¬���v�'�\�7y��(]��'���l��\ܵ8�+9���ߦ��V������-�L�NZ:R�<h\`�׆��}�sh�_�����8*��c�����L��2�.�����|n��U�7�z�+�7[qϴ�"�wSQ:(�}+��������'�A�����i��u��.���v��D�o�f;�d��B3�0�{k�iT��0xm9l��ۿ��V��0��"����^M���ڵ��(8�tѧrQ�LP5��k�(Z���GjW�ͳ�|(G�8Y23Ǽ-���8x���!�$����:K8H��,`��ь�#�9���X�&z&N��f�➷г��(��O�a����i6�Vd@U�
���n[��ny���նzr��|�R)���zBW�U5,9�I�+��n���|���9ќ��ݯ/W:�+O٩s���������AyX
n��؃0�A�lJ��r���ƭ��q�>P��tNVB��R�`����1����h�Asl�
lSH�P� ��6,��X��P��.�Q<�n(H���aƩzu9�Ӟ&*9�f��1�LTdj��LL~�S-X����LB�Ϟ�dXF-�Vre��x�9��뼌sM�������N�6%)R����
w����C4�9�)���"nf6��څ�����r�7�BE��x��'R�٫V9�V8s�=\�7��1k���T��'������N��f�[��\�w���lŌ�t��AІ֫�����E��i�`ѱ�'=����OQΤV��r��R�>�4��ZG���f
�m��׆��~}�c�Ɨ�OP��+f�7)SԶE��F$5wR"��<N@���r,���r�ӵOs�H�z�i�g��g�͚5ћ����d�D|����{j��F�=a�?_����"Ƀj���&�J0�QKFe��2S�Ik�֪k�dČGzW�\5Y��Eٌ�N��C*����eps���`��hf�ҡ�t�Zj��)�C�l�|k�n�7z�\i�t���⥝�SE��q�������WLw��Z|�vF�__C��L�uS���q���ivdM�e�Ǝr��h��0!�3��!A���[>���G�5����/x�U��7~ж���q4;�����N9x��W��(l����O�(�?a�L r��}��N緽���?M`{NtDd����ɐ�=�#�!ʼ+)�ͮ��2�t�6c���D�ni	�R�76��5���K����7�U�۰����;��5i����(�y�]����s�� ��}BJ��MM
"����ү�@�L�'�B��i�0p�Uy6�l��s)��[i�� CG���Jp�1'Z� ��I�B�F��[�o��%$�_��Ȇ��)�#[vF3(�G@x�#g��-#1�4�EG=*zH�دP�ay����`
ґE�`�����T̊�6aʩ���(��3-yy�3v.]���	!��B�mT!�K���W.��-�,��]��1
�D�4�g4��ږZ������:��c�/T�MU��oR����>��y�d��9`k*y2A[5�o��|��5����D�h�c/�*f�gi�:�,�\�"��������]���z\��M�vM�sj'd�c�_�E��F����ӿ�}ht��3�i|\G)�M�u]R�m�s�����+���ؑ�꺠���˃Geȁ��n��k>�q�	�^s�Guq(��vڿ��3L\sq\��wpz�j3M#��(��>��9J��0g��0��{^p�k��M�gS��cS�b1��=�Վ��z�m\Γ���f51u�+�7 e83&s(U\���U ����̌V��.Sgr!]}�\ع�Ggms��S�J�=�A�8�w$I�?`�����y��+)v��l*�l���B��m�!Nj��n�$������X=�����{$O����%��0����1U��H8�9]W��^}0T̝��k�jMC��(wiU'"r���8��#3zgk�}O��Hp�>*�P�)⾊�I7�e}I�NO7,�l����SmE�,T*�c��|��3�Z�N��3ŕ���5�X��X��&вY��bb��Ysq�ZR6vˁ�8<��pً�*cMN�c��ș@L@}P��Q�7)e��$꼫t��u����\��\�BjV��s������=�7�rCe��� 报��6v�gy^�ckl�Q���"�����]�v9��ג��NaT*L+Ą��]�,k�������-$i-����Nx`�m_�졸�w��/pl�J�m�n2vP�ŷ�R�ަhq�E	�(��~Ǉ^�1�
cDj�#&� ��1w.C9l�`�[��W ��V�oĈ�d�F��+iѾ�H�bW�јƭNP��=�p���>ux�d��H�0�X
g�W�\Oʨ�.���=���x�%͕9g*�3YS�FEʽIJ7�\%�&�$t,�dѸm��:��$�q����'�W��
/��y,�8�.w׎�̽���TU$�'�̷A�����Os����)G��r𑽦���L���e� ����2�;Lܙ��9��-�N�q�]�>��S[+rҦ�P�z���̝��q�r���f�q�;�'��z/���R�������73��ot��t�7��S7*/���5�~ri��q�{f�8�3����m����o4c�<��7Y�PL�S���L_۲��١���O�2#S��,�u����5g{�I�ϭ:Od��_=�3�s;����C�δ ��Pţ,�3��3�k�F1����[S��~�W�U2��|�L<(�#��D ]k�H�9��Q�sG�suy��]+'ھ�j�墽-hꬋ�<LJ��ڎ�uH�t�4[��y �I9;��*�5�&����y0��1�Σ�@p;�S �m����7������ŗ���U�:�@�z��ѥ���=	�eg����f+L���R���Ǳ9�ͣZG�yEACp�%�B����(�폵Ô-D:��{��~C=�wΧ�&��Ĕ!Y`:��%0���#���Pz��(g��w/�8�#����h���ts�������ꅣ�}^������=&���S��뉹n�R6�����"'�2S�Z�Օ��k���R�T�X����.�T3tW�����K1;����6�+S��%a�\3�����__i�>o�>�:&B�`�:�b�I��ۊ6�ǜa���f?�V�`�b�A�䬲�&5r�S�`B�N�Nyq�T��'{�@vW� ��f[ k�x|hɈ�n3�_ɚ�	�Jy:�4��rni�gާ8G����{+p��ԯ�M�� �l���,Vײ���5o|y["�9zpw�zx������'1�����Kς��SH��9f9�b�Ne,uV)�O��`��Ǵ��K�q�ԇ9�Rc�th�s����.+eْz�f�+E;��;z���m�S��ľ��N:zo �CkU��_�;��L�s�	���oqۿb�y�yT���͝�{���\Lt1W��[���r�\!�u1�D��/�S�V�f�Uc^�9v2>�Nΐ-_z�����ʘu.��0a��w��7j�VW�eLb�Y���u��Kv��[rLFj���H�/��F�Uߣ�\򅣹�Q�!��e�~@+/�G���Lh�����Bp�k�dČGz!5u�U�n]��\��˙C6ŉIgLb��bkBvy�y���%��.1"�Ը���N]��9�	���W��
P+K�Mz,,bޫ�ʷ�@D�+UE��]�m�]^ϸ�PO���Mde̦GeJq�A
�Y���፠���4�k!��B
���h�5w��70R%t��F�K�D�ӹgh���������)��FoI�c�;Uq�b磖����B�X�X���A���K��x���{"�p}�@
���&��]9ر���)\�f ��?6d�|.�Re��R]��U��^��@��A�s�P�y��mڋ�����DM�¹8�<�~�{�u���}w���i�n��C���/ ��L)�>��q�� ;��do%�mɎ �h�L1�*>��f6l	�\U���+B����q7���˘c������"���O�T�!���7�{v�{��.�(s̍�����<#ƣWȔ���ѱx�Q�?z���W�L9�3%���Cvk�nJ���,���/�L1�������˭�0����ŢU��S��P�{��"@���7*��6�͡s	؞�t93eq���A�U!�{3�橒�5�8� �ʖ
w�%�j�I���Ja��D�6��{**_V�sl���_F���4k#=�og�4�w[N�V��� 1M�K�j�:?��.���UY�H�+���Vx���+e�<��#�Xn��m�ϵG��m���c$�C7s��N�Ws�5:��	�n���wb���k��	�e�]t=I5GUN�:�a��0�j`Nx�^M�N���Ti�	���m�j��<�.ul����f�+�Z�U!����|�r�c�^��O��a�o�߈_0o�k|ҵ<ƾ�[xp끓򉶶���=ս$۶y�5v�d����m*��L����s+~�j��i��F�
�S�;=��a��<�͕=Tè`�m�H�����sݕ��]C�u:�cuc�9�#��͍��.'66妻5)E�0`0��!qB��kԪ��	��i�
ӿ��l�j�ʼC��T�o`�~����W:3ngO��6��\�k�#��)>qT���l �B&+\��]Ϟ�YY)��!\���b߲�ܰ��J$?]�>�^g(!(h>޽��b7��+	{��,n�L+�.�ae�lźT���h�L\q@���!��qkl74;�n��p�֑��1bt���P�[�̆^�~cj�\!d�*��x�A����tc�{�+Ȼ�S���h�x������P[<0_=v��FQ,}����Nl����H����]j�eE��2�a�"�g��؀��bs�Kj���e�N�$W�}����eن3ff�9d՝�K����U�X��`l���N�{�eŃr�c#|'`���<F٢�U-�A�u�B�1+2�#��N6���i�h�FX��r*7�= Zh�&#X���mS�)�՗|'3O�/�X����FBؚ���hU��ooFm�bb�y4t2�ݓy+�;قU�L�J�L�mk�"[�yͬ!≍��ui.������NRϗN�d#�)� *�� T7d2����#�:��J�p	B��j=L�d�%="�Y�En)�ʿ��
�}��] +���|Pܥ[�v�]e�ލo�s2�³y�:�Mv��ǩ�Н%E�,��y@�;��/�z{$�>ܓ�:!�TqH��<��dnv�tt���^�4�1,JR�Am4�]�^A�cP�63�����
��62L��.�N�q>��"�^^w��vZ�Q&q���L-?4�˻���k�/�+�����u�X�_k�n㎏h�d'���.�Q�XsAi��Gsk�t&�����nK�2R��!�)E[l�wf		�[����|yk)R�b�|��`g:���J>m�s����Տ�%��6���d��|N5R��$��X���p��mFA�����sL�ݱ�.�p�aN�Av��b�@�Gځ�f���:��x��=�1g�QA�7��5��۸�Q��R?D�p���ݘ-]�*`�jY�핖�	�i���zZ�2r��qZ�9�w�G8\ܾ����`u=r]^�f�jS{�|ұθ���H':=�)-�w��Mz�Fut?,���35o t��`�Z��o2VL5́ڞWEN;�����Z�ݿ�O[��+��{�!|�n���r�*8b�.��i��M�l���Su��60��lco
�*��ޤ̪k�e�B7F���Auo�j�89Ԓێmâ:·-�	806Y���K	ŧI����=[����P��B4ۊn9����8�YN�oU�z"d��[9ݚD0��ru���733��i�}����:���_s��6�4H�W�6\̓�\�����</U�V�g�k��[�a/J��q���-��:�Gw�g/�#�m�B�FY<�=L�A��]/�Y�4!x�/�k���D��dyې�i�h�wL%<�n�E�&��c��4i�75���C�E]3zQGQ���}���V�J�ik&����*|��q�����5�����/�ͽ��;2�Nэ=���q��̚��q���.�]��6Γt&�)K�RYkv��ݦ�c�s��V�E���,��Q��8�m��y�Gf��m&M��V�}��.�I�,e8��70��St�)E$c,�V�ԗj�v�Egi���rҊE�rUg��T?>��Е��� s!�hK�yL�'�Q�w�����/��7G��ˤ���So�\H��zY�Y�^��#�g��|>�����y�ZM+M�N�H�	r�LYRG��AzV�������w4�RW*�V
'(p�*�z�T�{�亷w	�Y^�B�D�e��j��HԬ�O<���"c�qwv���U��$�!Rj!&D���=K]ź���J��U��A�b\��(�L�u��n��T���¨�RD�]�KQ�tW'=L��Ew$���y�Ve*%���P�0��B�B$b]̯H2��%.YZ���H�����S�N�沅2�Ԕ�����e�U-K���p�=f�\�+32�дJ�T��*���K��:�h���3CUNd��!.��l��;�u��*�E�YD�(P��st�u��1fS�$M���U"�9�͢{���D��m\T�����Y+�� �eu�ʊ���y�vm]֝)*QS*�R�QSH�DIt--K�F�
�!BSS78�.��e����B���K�ZW�*̌��dJ>S7�0]ָ;5pR�էRġ��}�=�-�J��H����������)S�}�ɅS���}C�|B��N��C�Q����Ʌ�������P�?�z�xT��~���?x<�q�������@�I<�>���Ӿ�H<z��(��O�nɛ?l�SPX��) +��yi7�'�'y����]�ڭ����=&xO=a�ߞr�<�r��~�ϝ����F'x�>��ǔ���ro�`�}O�9=����{�aW~M7����~������p�?t�y�?}HU1_P��h��<;s������]���~M�~�)�!:v����oHI;�cxC��X�o^y���s���~Nw���
�\x��{O(&��~���ʈ��5�a���Dh�DG�#ܻ�}C�ޏ��x����Uǭ����7�'��F��'>]����m�<��I����7��P��:_ܜ�����0����xO=;x@���珞�~�w�*�c�'���~^�>#�|E}��������<x7�{}&�����ﶝ�7��{�緤�]�ǽ������ra|��E��w���m�����O_pz}�}�$}�{�M�D�+�av�E,�բ�kv��8���ǌG����0�z�xW;H���}v�y���x��<>ݹ9P����xM�	�����ς��N��|���ߟi�0��ߟ�m���#�>���X�#����+��/.-z��^��g�C�>�ُ��##G�b(G�"@z���9�'�=�;��aW}p����L?c��/����y����������&�����{���ˁM�UY���~
�©����k�K�����H���Dh�#��|�1C�|D}�8��cۏ
�]��ޓ�yC�k�o�s����?���Ǆ��;�?;�
�����n�;�o�rs폤�"!�#�#�"w���������;���X�X��#�Dz!���?}���[���a��;{O���뷔�	�~���w�|v�z��!���ù]���M���o�_׭����S<�=�<� ��G�P�(1#��g�GS��{�{���zWe>����[.��o�i�����~[���}��ߏ���0�~v�Ǯ���L>�۽o��=+��N�C���ӷ�����z�{C��ܜ �>����<"}��cW�z��Y�[�����;S����phB;y�W�W9ĸ���c�A��^�#e�.��{b���|2�Y�/�n7y�w�JE�K�jIҌy+.niݺ��en6�_�\��l-��3�T�a�:�(2>F����T7gS��I��Ճ���odӪ���"l��G�>�E��?|�B>�2ܟ]�ѹ�.�}����S
o���������]'���'>����~O�9>��1�)��|�/������1G�H�>�D����;oG��6*'W�����o.'i���:���L���������i�;z��׍��M�<|�<8�x?�}�����S|M��S
�L�����m�7=�d�=.�3k��~���C�
~(<�&�BC��7~��rs�!����'�q���ɹ	<�?��8������og��|��� xK�ݷ�N��;���o�/���D}1ή���ng�g�w�U�D iޞM�?�p��N���>~���S�aw����㟨ro4
��㧓�e�y���7�۷'!�]Ɲ���}�����S�;^O￼���@�>��'�b* �{y[����ӏ�﷤��<�n=��ǔ���ܝ����HO�~q�<}�N���x�m�����'N���_�Q��L(wG߰yw�k�{��}O�9?&�w}�q���ͼ�=�Ⱥ��k���G�G��<8��|���rS
?~�x~���;}����e������x�<�������~v�������$ܟ�c�xv����2xv��ם����i������/+����+��5��>�D��|�����r�^�e��xw�?;��o}��rraw�C�ߞ7�~w�9���ɾ!&��������O���q'��'��&�/'�1�����]Q���2>��јS\��������վ'�;H�8v������v?!�-�����&���|=���<��N�������.�_'��}q�=8��������Ei���s����-�9Uu~�g��|<G����ܜ��@s���~��W����Vﱽ!ɇϏ���U��ӽx��}O)�������{�I��>ݼ�}x=&�P�G߿�m�=y�N������m��#�ц�Pƫ�J���1��c�}Q���o�;ÿ����q�����?�����9>8_�����ǲ�Ǵ=�Ʌ9?&��Ǥ9����c��$��>8�>|��������>7�ߚ�>\Ύʃ���S�7z�vS��]E�Y}��T�V�5��C�� ��LAW�_���-q�E&t�?
�眕����ف��@����%�p�*���Y`tzJ�Mu�2���:G|.o�a���Uؒ�Ҵ���+!�0*��i��tҌЉ��n/}�G� G�m�Rv�����x���N�>�|￸<8]��C�yO)�Ǉ��Aɾ�'!���w���~w'�����aw�ÿ��ߝ�v�w����o�,F�������S9�~U���e������oHRq�x����nܛ�����)�~�|N����	��I�����n�o��8v�N����<&������A�X��&<"+L}|��W���Q�;�%���}�G�c�#�E���G��s�!��w�»(������zL?����7�|&��'{|����w�����=&O����ǟ���E��� �G��1�"G�h����M�˟�`*�ٙ�h?�b>B �G���\
o�y�x~�yN��M�>;x����~8��ڣ}}o}��]��T�nM�����G�޸.���r|w�y��90��{OG�ݽ'�>�ɇ�y��Һ�q]�<V�������>b>"G��"G�l��L�S�~�X���'zq䣼[۷&���<Ǉo������v����=���ޝ������˅���|���~O.>��ޏ���~O��|w��w��[��W�ytg�Tc�#�G�M �C�raO!����þ��=�r���{|n��~���x;��o(Rw��xq�>?�ǣ�w�$¿-����`�">���}_}�>���|an�v��xU[�W��������)�����~���i������7�<�w�bw��c���;�s����}q��9��=xL*좝G���&�.�H���1HC�\ň� �|~�}�x�������-v��7�R���HW� �����}��C�|�Q�ە��=~�I���������7!?���)�\
o�F|�rw�ǝ;U���xOa���ڠ�Q���ߝ�M�׿���'~��/V�3}{Зw�>�1>���n�ɉ���O��������'�?xğ�� _��ߓO��w���<PI��z�����;ӿ!�-�ۓxO�cü;]N�XP䝾=�������nF��y���[IfǢ�E��}��=��ߏ}�}O��>���.b ���!"5������B���������zC۹�]�O�p���?w�<�����G���v�"�vx8w"�/��-ہJ`���S����2�تN�/Z�*c�H.��0ʟ�^��C0b�m� {�+�Q��׆yL�#}OB�R��]E�سq�gs!]C�Ѕ)���r0�pv��d!"���9�cS�UԪGF�H�[�Vb�C3&�A�z�/��㓟.�������0��
}NM�H��;����xw�i����x�:w��_x�~B�m~�ە����}��ߐ�F$��S||��}Nq�������D�-��.���F��R�(^����(�>�yOhyL>-��;ÿ>s�Eo	�0������7��_;�q�����;Ϯ�������.�����'�o^�}����ߐ�����xW ]�aX�n�N������B#E����v߂��ÿ;U����y�0�ӵG�?>���C����A��������w�'���>>��ǔ���9ǿ69]�4�8�=���a�� �mr'���gE�z���(��~��V��ɽ���s�k� y?~�	�!$��������.��!���y��t�����rs��y�r��S�ry��M��bw���?;����>�O=ݘ�P a��r*)g�O������w�}C����xWН���oHyL?#z>}��z~;r�ߟ�\N$��v���ݏ(I�������=&���ӷ���I����'��N���T8UeG�¿~n����2I��[_�,��>`� ��z�`�!t�џB˯�����H����E��������Ǵ����W2������5Ńe�W���)6&�y�>�^�4�kD�8&5������ΤF�Y9�P�(u:�d|�X��8���"�Q5��N��JNܐ�f��3 fQ�C����k�R�/ '��i����	f'f6���ysJF՞�܏�^�;k�愇��C>W�	��x[9X�'S9��AL�����bڇ�=��Hqғ��yLB���7m�_>���s�h.���=��ev1�'�iǳYS��� }�x�|�W�Z�OZk��gR𴛆�5�w0�kU_GS/�9x��q�ݔ�-4cL�2�2��V5�k��;c�6�j��|Ogt��7�����2�R��ݾR82�y��9ecͣ�f������y�IsjR \G�Gv�����µ�1n�1���h�I��fJ& ���林q�e�~�v?���-5��C���XN��_��9�9��6��� J+A�x�F��-�7uH��s���	�&N�����fR��H��9봎�9z�2X�W"���sGncY�v��*OP@}Pd!i"�g���tG}��-��u��U}RБO�Vu�oVVK��:n���}\hqU����i|��f�Z�=��1v��0Xy��6T�;x��Κ�κDņ,"ju�;u�`�@��_"����.:峫<��)�lo�i����3�aIp���3L���o�O踟�#�]Q��#	��WC����#{a����Y��/Cu;�]Cj�W�'�4m�@s�268�t�;;�Hޕ��Oou>��4�
{��B����Ӫ�95\���%����jܨo��l��l�m�*5u�jz��U�C@yP�R_�V:5�8����ݔ�ߣ�>��\�#4p�!_��t�'\w�"g5r���EYܲ�tn�a���-;Sj�����7&˕/�M�Z�R�܍^)�n��^P�-\V����%��|�6&p��3����y�ծDb^�avv�[���RP�;.H�m,�y�Eϋ��?�QV��:l{�� ��+�5���͝���FaH�� �#/��i*�s�KR�\*�OQ��த�=��=�wrp�}��rU����Ks��P��*U񳀒�;�S�D�Xv�D����  ���6eס;R���hS���b�"�i�ω�.��,�u,���+��1�*r/n�B�����f�fT`�ɦ�2�^_�+�����B�Λ����c��8�y�v�ۄ���eqS<�/��@�Z�����/�r�Y����P���zc���&\]׋�c��҂�S�J��5_L�w���SF�l}k�Hf;
�����:����h���|U���c��|I�KJa��;J�]A�o9J�i���%9���'�7����5�a�5���C�r2���D8Uu�h]��9����m��^K��`ߜ��I,������WO��:4�f ��	�2T�q #�QJ�.��S��M��Nn��ݓ������c�_Trt�؆�w6�7z��F�]�ӗ!k���(&1#��g2>
�u�9�b����)m��B�ЗbZ��K.Nk���Ȏ�,ĶU��wj����5i�WG�ٝ�ά�"إ��dw���-��ɫ"� �ױ9�q��vnJڙ+�Y���k�}�]�F��#v��k�Y_����y3�=�@V��]e#ÿPw�5���tn��ŗ6�x�`�$H]�G��l���u��M���31]
la	H�Q�+MƧRÞ&+�vh�Cs����;�y�!b�J���&�8�>�ǐ�����|}t%��S���Ww�7��gl�+�G3���� Iz���%�,=���^&V�n��/,�8�W���<�Le��p'�Nz�&=Ѹ*�|ǋ��,.�ʘ��+t�=Tw]u���<�@#��M�QJm:=����R�����Ő{�v{C�?=:5�A���u*Ѣ��cc����Z6n֋��'�L�L�%�#~�j��ʦ��N��&��}7��/$iʇ�%��#���BgG��A��(��1�2��w^�|q�J������[�k����׸�q_(j;��|��D�ԇ��3�zhs���(D��V=�c6��������)����s�R�F����3?AQ�iHn��>���b�*sE�o�{ӽ}^B����{�qa^qt�{#���n�s�'��u+3����
4�9�0v�+��d��5� ��W�,�Jrǖ���Y���o:S��N�Z˫Ra�B*}�Ea�L^�]ɡ�� �gnj*��"WBnղG-2Xwaڛz�}U�}���V�w����Ʌ^�@vN���6��/�h��$�+�!�Te#�g��;1#�J�[�(\�̃E��?��؎r��t�x���U_*�h���@��JĮ�|��:�>�:��"C1̬sC8�&�$�;�Asv���ڶ쌷4�ҙE��W+�Mn՝���W�k!|���Ap�O�g+��U�o�k��d#ƴ$�A��mH����@6�y-��Fu�=:_��}�CQ
����������e��9u0�k���}�wg(V�QUv
Y���aQ)ƚ�%Ө��2�퉘�aL4�Eݮ��������N_ed���+^ř/��Y�g����7
�����f��OK=�/�t�#ˮv:�57���w�%+��%����km���@��`ip�hhv~���c��7������Ѥ���oj< ��x��Uc��S�He.ܧ�{u����xh}��.��Y3�a�X�V�M���k.������Z;�%���Or2Y��L�ү��=1q��s+�Tɋ���]M�v�f�[e˴w�F��N�]HT�^�5i��0c���U�%`f�S��h��vf�Fe�X�VV�Vʛ�1�5��8����*D;�]������Fe$������\�x����'sM�z4VR}O�j�GsmOt��4)�'n�A�>��UU}�����&�l l��b���d�W9G�����HƮs*�Rs��y�y,�SA\�X�ڽ�'|�^�T�F ̣0�p�U�a#���iLE��WS��2�V�X�^�ޛ���7��r?H=䠛1�X�=Я�#��xV��G�,xFTS����g1v>���v)�S�~���]_L[�G�aaD�W�_�2�80>RbR��x1������*ˈ������ӃD0��1�6b�t��ț�p�P$��jl��rtչ�*(�^���@���;�	���9�2�柘�}P��.�N;��۾�������g� I�%�NF����*�g"�����]�v9�����=�Wz���E��ַ���r�:�U�r��6�DHD�K�B[����[W�F�ݢ��V?
���N�=�S6-�U�M�wM��~��`#1�@J�N�κ�Q�8*�E!7I�62�����ڝ�t��hgźD��N�ۭ�㸚0Y��~H��&%m:;W����2,H.Vư���Z�Bj!��r���燐,}c��u�
�j�1^7��V;Ʋ=�x���*hͤ�=�f7`�nWa����ɽ�b�q����v7��ik���o�ֹ��r*�n��i@X������2�$�]lK�r^��hq�ȍ�諭��޾&[Z]��kѪ�CZ3�T94���C4�,!�OʩI�����!2��qc���͏����"�US��S�h�t�7���ک'�4[r��C�2J�f&���gL�k^]�;�՜^��Å�驇��,�ʣ����U��ĝ�1��~rjܨpN܅��Qܷqq���R1Qh�3���>�1�^a�;�JL�����o���f�f7f�{���V&��N!:�m}o�͜aT�����6+���}n�m� s�a�k���sg���m`�6����;�[�؞�?i��8	��G��׷�,�+�ܔa�)���OcCg�E�)��v.�}{�����y��"�i�]�^8������1�d�k��F�LBF�f\�N�Ԧ_l<��A��utܝt�`L���;�!��J+�0�	���鋊�@��Z��it�f.�Br�Y��ۻ���O6�ѷ;ʧJU�;�i��Kb9/#�����}�2��P:�1�}�!�芌�]��26nq��Y���%���L֫xm.�����'o	�y5�ly��!���޸+6*��n���
kv����O=�z������\s�*;Bl�i�oV�e���[R훛�u���C�l�O0�+�CjmF���,c�_^e�P�����;Ï�@.*��fmȟR**�N�Q��;y��
�hU˳Sb�0�{��=�ml�B�:�V�^fJ�n毄��Բ���7���:`w��u�ZYkqvf>ʊ蚸����Y�e�:6Z�x�h�;�R31#O���w���N��u��(��9���c��%g+�[�&�]�w� ���k)�3˞fQ���n����R�B��S3/Lꜣ���8	��1%�i+����r^���u�8"29W��q�)wK�f1���rY���)h��XD�Y�6`�� �o������'v_tpA�	'�H��q��M�`�9��ϗ�Ž�Т�����MF_X6�&�z�l�ܝ���@���t�;�pFp��u�}V�R�⧴�^9ku�+<z/6F��+�[��otn0K��n*Uo���k�J/Ma�6�r�(�L"w�
t����
�A[�i�6�<w�,��<6����5ZAf]Ak+a,���֗:ٖ�3ho�N1�QwF�j�N6���8VhQBq�{�@&h�zc����D������ai�և �M����ɘ���w%� �"1�T��L��gP�u�EF-��!^)��{���=��]s$.ڬ�}�褍�2n^�S����[��#�K���g8J�>I']���^�+9=�V=˸V=�W�V�����/e�|�#d?�-��-��$T�Lˡ�Z�U{YW���z�S�L��9h�qajFG��������3�r�5+W�:���#���C����	_[��N��[5��B41^;�iq�j�f%oO:E�k4� �b\�y��gt��ok�`��<��W��W^�Pe�����Cd� <��E�9��E.�S>Z�b���i�����Ț��z�]ӏ�����y��ky�3w'gK7{�ȩG*�]���]kE"vz+2��m��B����u�>Cr��5��B;nԂ9�7	���]ʄ�x���SN*]��TZ�f�_ʶ�E��g��S��J�Bu�m��e�	��jL�ߘU�f̐�Cuu��#w�Pr�<sU�{��޾��ld�r� �L���b�]���_,�Z���wW�n�����₷ˡ@�$�S�'0�fuZ����}�r�e+�&9�%���%1ar�۫�__xwW�|����#WQO-t2�N],eKKv����|31��6)�}9Q�w�v&��p�7���6�ŔD�-h�6JӞԠ)%ƕh��0uux�an�&�juٙ1��<֛b� A��q`�bwT�Rָ9a�f�È��*�A+�
)D���Qjea��]����9�j%�vb��]۞P�*�,�"���H��t�J���Z���ȳb%�P���͘r5�]�<��Q,䬋2C��xZ�
�PU�VjYT��i�+2K��Rf�K5,��(ww
��T��J��$iV--V�-
E4�Q��S�j)�Z��#���R����QC�F�	*�U���\�1t�v���xV���
 R�fL�UR���#�֦���$�-�tLH�jeReJ��B�J*�B���A3-E�r�Jjb�(d��eCM*�l̺R���ib%�U
�ic���Ju���-T�,��J�(�R��E)IbZ�QjT�.I⩗CR4�"��IJ9�QfR#�M�DU�8�$#�!���"�ȪL4�=k�˨�QK�]K՘X�H���,�3�V"T��5U���4�ǟ�.�={����'��5>�{Rr��*���5���i^��N-r��Kλ���R�H��S���v<zF��_��諭7tu�j�j�W�p��1#�I�W �	���Ѫ>�}��]~���:tsc�����K����yצ9S�P⁘��t��7Z��y�:Ζ�,Iu��쫞N /��K��nㅗt��s�IX� �uHMB�)8@iP��7�9\.�
��z�=Q8BZ���1*�g+�9�|�C���!��;�n��͈3
d�ǭ�n��;˔����^�Q4}D�r,V|���:S7x������'1��.m����٥b۵3��C��BU�m�0���w��x/*�Aп���b�7�Ԇ�	��4����5FL�v�[Kx�BQ��2MGOW�'�٬��m_L�;� X���V�+�ַ�܆k���Q��zjR���`z�+�X�l}���A���OT@Ʌ�wOś��҄>y/Iv�TU[��&_n�S�!6�xs�b9k��qb��
:�FM�69�;�
~y��L�D�$�Ӻʫ����SF�-���c ��r�4Ts�����f���8`�m_�bB���ٛ�~��=Bׂ�3]$����Z����6�Sm�r��].��c\�sxs"x������+��`7���{���'w�n5K�����?o^.C��#y)�	��V,����,�xd��u�Z�J��|:D��P}�}��|��ԬM�����J93�jg�(�و��|�k�d����&��^��q�n_{�Si�^Y=���
���8p���4��T_1貵.�MCȦX*�g���w'z�(;��C\�x	���M^5�#����6�����B���b*'UViuag�]|�	��0��#Q�X/E$\+��cϨ�3Y5������*�����7_2ǅv�g��e�귔[X��L���G���r�k/=I=~���&-�;��'��
ĝ���GV��O��ǝ�Zo֮�qEi��T��9��:i����\���Lu�+�����^U�J�]z�f��6:�0�Ti���ǩ5q7���ๆ;N' Fշde�摔_7��3�xȻ]��D<�e��|+�2�C�3�F.����c �ґϋ��/ �-]�ʙPr��)k��҇��D�졨���Lk�^+ेe��*#�[\u�gJ3�&�Wp:�����G�Mo�{^9�K�W�3r��	T��S�����i]l|=�U3W2��f�'�ܴ��g����v�T% �p�{�t|�����hE�6�����.=�"FB������#謠-fVFPxVc��� 8��fwN�v�}���ɳ*����X�e�j;?�*�\+�/�"����j[R�6��ץ3�_�}_W���y%M��8ڱ���k/�䩒��偮'�9�#B'��ZC��Y�]��пdM/:�wһ�w3�n�!��ښ��c !M�K�jŏY�/��1��i�Uk�ޣ~�W1;w��Ȭ����6P7P��V�7|�^T���֕a�<���p]�A�+:�W#C.x(���M�q�O��Ҽu���Ի�#Z������i��Ӝ�2�j:2_-�S	@�|Y1�s�
�r��pd�gR�q��3�T���gKr�9X���4�(��:�ݜ�o+E�0�0�ϊsXn�Po�j���{�F�'��K	s��M	�z{O�ٝ�����@��gmT�sB�<JVg��<jo�[w��Uljv�α\��5C�`L���Ss����B�L[�G�an�$�C�P�-)F�y�'��:����&5�}�]��.���h�^;��[�LnM֎�l��C�û�����)�R�UO?�x	��Q�2�1<`#	�+|s��t^�٪]m�ç�'��~�\T|�{GҔ��)��2h\q��Ԧ�Ӥmμ�P�F5�9�k����+�tn�)j�^p5��7ws`��t]s�{�c���2��n�`n�u��)&�=Zn��$)��r�gJ��+3�㯥f(�T����zy�3�G�>��� e�N�:�>����l5
L��<��H�x������E����iS�ʢѰ���W#�^�z�H��5��?���s�4x�D	�Wi#I�S�ৄV'\4T̨ZX�
�'k/k"2�Z�s��A��S��2�P��S����!�����K ��5��ŞT;���d�S����ͫ@7(�P���mցp��M|`���D	ks��
{��)K��w<�SU�
5�Q�L9=	��^3L����&j:Q?gw5���DW�e������xԲ��ϲ���I��Q��\n9=���Q"�O2h�n�~�����G'��c%��E�I�;�}c�A����쾋|7���S{j?���
u^����t(y�$�j��)�u�G�)�ϯl��͞��]bc�
��ZL^��f�+{[=
Z~�ۀmv&�o��6�ak��w�o���8¨8	��m��G+���s(���pv�j�42�|ߦ2��"�c���*w��Ln�M_[i>��ݿ���ꏹ��a8;�Q@��A�x��:6������NoTV��x�����M��Q�v~\����8N����V�{��K��Ub�Ycju��Aك�uk���).��LN���9ہ-[���N���Jp%�[W�:��l�ӫy��bX��&9:��+���L�|
Ӿ�#菾��B@o-e��`$�%4�jȿ��Cd�C��t�j�CW<:3�$ĆO�.o�Z��R�Y�Q�ꙺ�h�.�J�ȭp��aY|a-��j���}	.���=���&�#�N������:���� ��N�W����ea�����G]9��L�UWS0���Iv�����q�GDj)�]�P��s��G�|�����_�Q�X��w��!��y�M�tt����㯽�^�E_�Ψ1P(|I��@�HuGʺ��t}.¤�~h���X��~�J3+D����,��k"�s��p�*U(���I0�H�hUÝ.:�x�=��5�3s
�C��nㅗt����A	��1���'�$y@ �H�w����7���~s�`��\�Q��T~�^.5�')�l�s`�Л��rJφsg�i[JR^�ݒ ��8�*�h
�����($�E�]�=�����6�t��b����Y����r�.@8s|Ht`��3��F��-��W�v���C������E+�W�z���ht��)�p�{���(�>��h���k��#vzy���7]\M��#�� ,�d2.�o3Ȭ!�8�Չs�kQm���○����|�.�4��L(帪1�:��= ����e�c���ec!��"���ί�_}�}T[���'�S(���LF��Qq�ђx"w���CV<���N�>>�:��h��C��{rf�kyM�w��u�
g��-f��K'�L.�;��s�xs�8��"󐜡W�Ֆ!'	Z,ed�|ꘅ�C5��b�ҙ��u"*0�r�gCG�B���n���&�P|�^,�S�v��x*�j�����1�un���`��z��O��W�Z���Hv��&�x��*����2�(�و�j��*��Y;��j��{.��x�T���K�ެ)��X�>G�y�K��K��/��Y�pz]xG"�`�`��.�GowrR2l������!����$����6�O�w֕VF�V�՚�����xΤ�m���u1	�g�)��g8�B�F������\.�R�W�s(����9"4h�Wm؇�iN�>���޿���Z%дauP�'�_V���R©	�j�����Ez(�gd[���Ei���O2�� v[$c�U�$�ކ��"�������Xŉ&�_D�=m�ud
�u	}99ԭ�t��Vg a���g��8U�2`<xn��Wc��5i
�.�B+O�qI4��d�hL�+b�ld��v�:(鍪��w/k������Z�J;q��VE5�cT
P\5(N,�ʻ�_W�}�Ϯ�K�Q`���`)�_i�ʼUcx�&�&�X�!�c��rmE�dfܬ��z��|�lU��UԢ<^[�&"R����C�3J��òS��a7�#[��y�%���.z�(�6`ۇU���4Es�j!#=��:�ܡ�ò������F༂��^sw��CC��vY)��k蟕*���*N�1��D`�=v�T�x�-\$����m�)G���!�?W5L���^B��)~�ra�����eD�YC�����bm܎���Ћ�s\_���ݨb:5=�3��]����|ܰ4��-��v~���ݒ�f��&���"��]�����2�=ǉ���
�.�ϗ^�n:�=�.t�q���	��F��cs�vIɵ[�/�͸1�P�?3rż��E�7s�Zٿo�.��������9g���S1{�u���,N��ZϾ��8��C^��N'&I�I����M*����b�����9��rޝʌ��g��3��j��7�q�3QU�
�<��e߭���{"��%���n���+1�ɧ������y�i�9����5]��kjn�ֲ��65�p{F��ۢc�V���.�y�}��4Dz3�o����[���*j�v�Y���%X�ަ2�.':���##�:h�{&��-��;������ǨI�I�X!�u�dur���Sgq]}�m���S����J��b~'D(�m������,[[�kg}�]�=Fq��uƨ!��e7=�<�!_����o�Q�XXQ%^�A
g���ޯx1!�b?���c�}�W=>��W.�Yx�0�K�u��k[8Eyk5�=�^6�G�ƀu3�>�r�-����	��r��#��_�O�j�`Ncʕū]m�y�m�~Q����N3-�W�^S Ҙ]=�n#Il���o��?�g���J�#���=����<�Sم�#O\d��S�B}��� ���H�J{��ÔI\����y��wyKQ�zJJ���e�븛��.!O��	�(M�)Љ��uq�g �O����S�����eﮈ�T���"b�1a_Cn�x�&��f��~�+N�Q{#�k�l~�8����딏V}	_�V�j6Ҩrju��%�8:p3%��{��]����E���7�=��?x��<�G��;j���!Zz#����U)d�&���dƺ����~[�z�<F�w��X粦����U��k��+�k�����w��z(�|�lm��":2t��A�#�ƃ:�ʒ�ev��z㴙��}]Z֏���KIl��0%�QAL5p3�Z��,&8��w���C�l�����@�Տ�}��}�	��H%{�H��9�$�zE�#~Xu=��[lXаl��s��\(�7�ZҺ������4������P+jMZv���� �m�{B��^��>�1I=<��~)�w1�-�zP������\�#5��j��|�b��$C>�XlW`�A�룖f̶oU��'FM��:P0g��Xr�c��u�뙎fFaߟu}QwR.���EC+����f���<~
v�߼�T�%��������E��6NG�~��i��ep�Μ�	�O-�ni"˷�������.����T��h�."Yd�)����5�ƒ���[#��W_.�"������&0�@�Ф��ʁ1��˾��9���r�� :����ůZ�se8�{��X�Qf� �p
�v���kg8*=�lDu���G��^~��4|�c����Gi5p� ͳ�@�&8�L���	�WB����k�]���n"s ӭ��"��9ܴaF�u�`�.�a,χ��J^�l���۷�ы�@*�Hf��Cޙ�}Y����W�:B�/b"�HW�����U<���#\�z�eGO7�]v�H5���sv�R��nV^�[��&;�Z��úS�ݭ��d��KV����eF*+R�\O�=H�o87�D}��D=�ͮ�P���|�Vd_p����n%���>;��'�/]R_)��lU��L�r�oyҾQ`0�����F�1*�g:3�e9��_
�9�`)��%LVS��v�i�;9.�jl�[/���J�Qq�/�[6\i�c+�[����I]4q�W�ɭ�t�^�߁S��J�f;����2����1�V���C�c���n�%��:�BdÍ֬�L�c�.4�2F�6�����s�ӵ���E�R�q�0����5�%!72�����h��e�N�58>���H5���0��N��wY�5١�IY/{��x��G�$��`��9̱��f�%�MD'0l�G.�*�{8�\ƾ��վ����)T+��H�1�,dFt�wk���!�5�h󩃝����تh�`�}�o�U���t�p�
��8�eV����J9f"~�j��*��Y1#ډ�\��W�����aw��!��X2�#�/�K�0���^g��z-'��.�(UPG�vB�X�6��BMf}ntG���-y:�0���� *R;p��4�.9;�.����b���.t,���*���ٿd*#0�.u���vͺmb����T�T}J�0�9a��b÷L����7�=�Vz�(o#W��ZK6�F�H��ԛ{�$�Xu�_XI3"9�
-j�sy��3:�ޤ��k��ϳ]#Z�4z���E�VHU]@K���ܰ1y���{�n���'pD#t"�� dƑ�!&�u�L���|�u�rl;N����y[H�*�7Z��E���76��+����D6�`6��%�r�j�v��Qn/�f������,��r��A��VK�͇����/I2v.�O�Ӳbg�l�2�_d�8�
y͍ �|ӷ�X�O�ym�{N7��N�G���Xv��t����B+(�q��jr]���O��1�f^�;ʐ��P,����� F�ih˗�*�=�$�t�:ҭ��J^�Wne ��+G�ֈ������r:^�h�V��rE2N��>\�%{u5f9J�n�:��V�*�Z��Ѩ�Й�NS��2&�
�H�y�{\z��<6�����m#�=c���1��b҅N(�� k��uX��Vŕ��7���5�H��s��Ne�|�� �Y���j
��ŷ�Gn��\�/v�2:��j���uA{ڎӫpV鋪�츶��L�j�z'7�D`ahq�CJ�g:�ĥ,��uү��H�|�u����E�{�.o��5�;�'�z���sQW^� qӗ�^(�R�)�������ɨ�o{�T���eBI��qߺ���cr�d�]K9qt`�t{n�Z�s�d��dD�	f�_+��4��:�\�P:�4�� @[tt]�Ӥ��3]r+��z�rř݆g�wa��<d��*l]�^��g7�-����jF���n����VmNzz���1�фR���]� ���w�ql�mV�<;5����X��`�%�lZ�1w�9y���ާ� ��Q>�I�]۽h���l����η4��A��6�����g�=}�@�AV;q;4����!��w�
�R��-ʏq��Ĥ�{}ZaB����i�.7�X�2z<8l�B-��6|-N�#��f�`̨�;�ê�Φ�� #�	%Fa���9W.��kp(�诹	��6���%F]#���PX�Ւ��f�J�V>M*lK�ކ���-GS:�}Rv��䱺�-n����ʳ�\�rSE�\k�k+E��Bu���Xm\��o����8U�ݵ�Y{��H���/6J�[��拾C��3�X�N��[�ѫ8���b�G7��l�WE�e�ۯ�,T�j�Fa�+Z)6*��웷W+Um;�a�]e��(w!V|*�ƁG�9�����1mga;G���û@ϑ���m5p���
#���YbK��*�\�wr�S*B��er5(��w�+��"���F�wH�"9%��QE��*uQ"+����9z�U!H�%#9�Z*�gJ��e(�H]�t�"�R8Ql��JC��%J*Z����"
.�EF��VWS�I ibDJ��h\��UvDA�RMd�T�eI�s4�g5�t�bl��4-�GE+IhT�Y&J��2�U4VEr�+$�"S"JĊkIkLΡ)�d��DY�˴��E25�vD�� Ť�hIrDḪesbYmT+��%��%��M�.*'K,�Ե�Pr�²�%,�����E�G:F��igR�,�+$�MR�d�)�T�TSD�9L�8J��:�%QI͡�5"�"������0�����y�;�>U���ڔ���n��e���/3��-J��g$\�m�K]	M�yr����k�Z�e�DC���UUT2�-�O���Q�F�&{q�ۈn���`�t+¤tWt
���^�[�q���HGP��Ԍt�,R2�c�=_ �9B�͗:��	�!�̲�%�|�O��!���;�]w�i�.�bJ'r�ȑ�1�SWb��|&�r΄���jPu���3	1�}}R]׷VS#;{T�W\O��Q� �+b��2��R��#¢��w�'�"��������ߵV����� �B�0�h����V7���%D��3v��g�6���uR�gmA]���.$'�FY ���"�y��]���һǅ`᰺Ύ	���ً�4\����5��sK��-�Rk�<�OyQ������#��DW1��'�c6�C�Ψ;����Sk�����r���AmYg	�D�'��J�j8ʓ�f9��1�t94���O�#���<p��1;�ÜkW!��~��j�/ 9`kυ}`'0D\qD�D!iz�K�/��~��ly��R�������
��CZ��ګ�p1��健�[V#�~�����)�b=r�53E2Pk����U"��J������h��OH)�>X�Z�2q�q��Yή\҃3��:�]�3+���� y$���|6�q�yؤ�'d��N1oi�Ԯ�u��+� +W,܎�*;n�*�OH�:�h���;t,b~������7��k"�zcD�s?��^�r�X�3�v#�ƍ�B;����:��!�vi<�[�7m*��rX����ڣPT�	��տ�o�0䋼f�NJ��|W�Vooo�q����w���p�E��L"�5��u9G�r�e�Ԁ��=�k�ni�#M���ڸ��=P�7S��7V;�#��1F�T鿑�3(�!��U�a�ZH���~k0�ԫ�m���ŵi�
ӿ���:�~�-��[�S���,�������lN:qW��N�U�#\�W*.!����"���!�1
��7m�K��j���zȘ*��dW�[��8����$>1�@(�bWp�9xT����f.q��N�s!�%݅����g������@L@}P��Q�.�`#P4/��{��>g��ӑ]�n�}ӎj�{�X��p��&�W �<z  ��:̭2���V��M��7����rZ�xZ{��N����h���i댖>�k�v��(�#���k���R��s֡NH	zp�兒�#��«X�+�hʖS{#!C�KXa#��Ĭ�Y�\���v��rh5B��$������w�|��+7t��si���s�r�����peE�]i�v�@u�2�#�9���9ُ6�H��X�sc�}�DGVc����$	���CFKj���eNwI�n�����g�� %I��˩�.���YyЏ"2j��s;p*�W���ɫCt��XD�6�@v�$@f7e��U)��e(_n��Fl�Cf�n��̨ۆ�=%|����� h��,�I��&��d5��rL���b �l��%m`����gh��S���ڨ�K'�4M+u6�Ă�n�>@����]�x<��]i&��B�q��������G�ڏt1�*޽N�U�%?96ʀs���V�!j�XU��ƽ���57�1^�d5�<���˱=N�pci�����){><�����|P�7(gޫlW=�G��i�ze�.R݌��� X�m� Wێ��FY�g�f���G�_λw,nӸJC�	�#[�7���V3�y�ժ��%8�@@
��B���6NC��t�&��\5���JL�L�u�)�u�|�/�tY,a*�;1����1ٗ �'��V�Ϡ[UP�ұzn�]J��sՋ�;��/7�V�d�z�X��hr��� kKf�L�x)�w�BlqV!X��6�(�"m���I�+����K��6�"�L��U��
m�W�O鲶���ά1�"KT�*qd�5+�]�P:��ҥ姽���_���������'�ՓY?~��Z:.�h=uBgB���_L\Er�LTbu�.�6^*wO2l�����{= ����2�ۿ�D�̡E��d��@�����ݗ#.���ͺ8�v�"n,�|>�P��,v�M\>�6���'�,��P
���*��N�<�w��*Kʴy�:�\JF��[ϡ�����V�e�2��6ȺTL�~�~֖�Vo���Rr���@P!�o *��F'�r��>��w~�8!7Y�@c���[A�_M�̹�\H�����5b�1���P'�⻧���#��l����1՛
�.4GVfӟ���Sb
$��_�v��*~,V�ˌ��Pw<uMv|�W���qyd���#~�;�[;����䴦��^�ͰU�`Ҿ�f;ֺ��)Y
�v�{��3�z�k�&&�W-�o�$[��Rb��vh�b1��T\V�Y�<LcW����.��m���oD��6D��n�^#l�ᵪ��-'wB�`)���`P�����H5��'�d�i̼�)Y��~�E"~�//ޕ�z9��CG�mѺ��Ҏ
��ʿ?1���GD 4��iѠ�4�dL�n���!�\���v��ޥe�f]����Y6C�*J�횰�t��X+GkB0���S3�./j��h��ӷW-,���f������U���9��/uT�Ǝ��WJ�����ed�G:�"ֺ�d�`�LČ뺑��7�ќ[X�5}��XL�َ��h�Q��8�{���b	/	��LCG#���.����(p�������DvLh�l��b��M�S=�Qó|�CRgYD����˭���5�\��2�p�_�q�yЫ�X'��x�a/��/3�.C�=�̠7loN�et���9�����Bݒ��q�6{>5�7o��Q��`��R:+���V�M/
�ަ捛W�Ԛ��ʔ�Ў�G���.��HE�-��u��}s�R�F�����cۺX�����:1%��lgm�S-��A�WI]�Z�	�C/ ��;�鸚�g�Ҽ;�)�����e��~�v�e��}w��+O�*xs�r��ǀDw���2�W��#�Q�}.tu;��,�|����!ʼ)���Ɍ�U&�&�X�!�c��n��.��I��;��oU�΢-��e��#�����J�p�ftpA�+���++j�5?e5q0��A<u��lm��R�lD��"�aD�[���g�̵�!�am`�
�G_����H�	�qO���r�0&��ǖ뻥(�1r�c;�GI���F�4������L��C6�"�[��(�`:�@�ׯ��˵�'��Ͼ������E�J{�m�X�A7ţ�1�*!7Pr�S2*�F�U$W1���3�1��xd��{�)�zR޸����i�*9���|[VYω�D���*�Γ�r;�z~;D�k<�.���GKw�@�gI�9�%���\�/��~��j�/����N���( 'G��x]nr���]����hM��8a��ۄ5<}���c�4ۍp�;�1���:{Z�9���{�2�K�5���o>��+Uoxꮞ�g9�߹j ?���sx���^�3����w)x;�m�5X��i�q}'x�w�2�T�|�������J9��t6�m*�u�fW�9�f*���9�h��R�Y�
��m*��v.�2��W_���ޯ���!w�U��,�ɠ�6����V�g�̥�����_��v�S$[1��kՇ��$֏u��GFKWړ�pu�{���*uCWe��cb���>v�����S�2�)�=�}z��'R�ts{i�\����%앢�
̌>�}�*�%oM�.����=���5m�^ d68g��I���#�z$x���4YY�Q[����J%�#�4��ܫ;�%��uZ�\(�%�޾b\lڻ�ο}}�G�-d^���z�Q�E �N`u�I}Q:�*�J��io���[T�]]�]bg[�p�O&�E�f�P���0T�II�uQ)Q�I�Xװ=D��b����h���^�v�@��7�����b�������X+�)�e.z����:��j74�=�����q�V��r�r�H�5�C�B�]v�_ǀ2��;�f��G.������7�e��;չ	�l^ח��#����|ZR���E�&�{�->Y�@o\��\� -U�.9ɤ�|�v�|�ȧl��ʥp޸:��x3"�jjs8�|\�GR��N����9��|�.1��H6I[e%4��v�4�(p�cp�j�ɨ��w-��<w�����3�319;6�9�Tȗ�ղ�,{�!UN|/��=~)��v��f�u/�&.�Y�sj�kS��m.��Z��}m@��<��]���:-v@�U>mq��RH�zS�+�b�������eqR���l��;mAM5�I��+r���7�ZҬmb<�I��L�C{�<��S��ǹP������
.��.h���1��څj����Y�y�]uB�6�v)��;a7BuQ{8����(Ͷ0�0}��}�W�p�R�0�V���6�#��Z�_(�n�d�A>��}��bz�0n)�A/K�3�(EiN�zv������q�Wl�M �����X��zf���|"��D��D��^�
�i��:�֚퉛>>��b�d-:�5'�.�R���vQw �T���hp�b�����T	�(a?u�Ȝƣu.�Ny���Ҳ� ���`��|��R�Ϻ{%�fb.z�Y'��u%#t?�G<�M��y<�⺦����+�ϼ�Ֆ�Z�S�FJ��붛�MA�>��5�=���Yq�����:E<_�k������]�����/W\E*
�-4Ryq�ϗ��W���EC�DL[�:�*�{�z�2_Ǡ��V��`[��'ƾ-�\o�>OtU�2��d��z�k���5u�OO��|�t<	����"y]�s�W�{�_��u�� ��C��5�Rc1v�3��s��W��
K���<<��V͡)V�
<�)]�[��A%����9oP���1e�������q�Q}R���ٲ-�;��y�����3��0�3!�:�+�LU/Prss7�!F���(���T9t�ןϾ�����l��oWC�=슇L�!Lt�.
}5K�r'��۬���sA1*�ɺ���ØvøF�JH�DΠu�Z��m:U+��hn��"�Bjs�[�R}SQ�15��
�5��l�Z�z��f`���VE<ڇ�۞�v���[Z��$�j!c�4ہ��UDk�&5��׻��~SBr5]cxZ�o����fW�O=}����ܬ|��Z��E���qk��7C��f�I�y�j�>ђ/�@�u6��%`ʎ��r��^���"�Ol����[���kkBo�*�_��xfQ�[���DI���b�������S���l�}7#.��{W{�W�禚A��̢�`�9_	P����l
�fSs�$���j�F>9�����U۷�7�^�	��ʮw��W�ؕ��#�յ��飙�����Ψנ��h,��o�[�Ӫ�/+ |��=qFٕ�=>́�"�ן_Fo�/!��H��Tۓ:&xn� �X{LJ�B�\!趛ʭ9��^�|=o"��Yh�6b��uJ\Q6œA� ��x�����M��[u!�]�օi�v̺�j��&*Ɠ��oxc=�6tn���調	WJ����@4�$�T�qWIR���\=e�8[I��kx�+y	
�̇n'w��j�h+�T������%-4Ryq�ۈ�gnf�C5p�=ۭj�B"�����3�<5'K����p�ͷ[S=�/[%f�fϻ�Wb^��qw���p�B%���4+�!�H�N�1�j7w�9�wY �Ɲ(��;7�w�d�)62��2�S!*��s��̬��������G>㕮%_c㜹�kBa�W����C�]P3�����E�if)o�[����].ٽ��#Z.�o�k�a����rGs��.��|zV�jl[:��/s/�Kj�umF���U4�������df(X󌾳���psS��};��
�şח;�E��ymnU��'\�&����a�I>Y�6^��}�LL��L�΍f��-��m�U��Jy}V�Su���W"���<5���;��Sn��Ʊ�q�E�Е��
z�����U�k]-cn�v�Q��ҋ��V6�/�ȡ/�hu��
;]�+X���d&�ib[�Ѽ�ŷ�lR"V�%�� N9G:R�au����{%�Y�M\����S'���jU�du�,���E)v�$��R�MB��۷��*G����{��Wp�X�<�1��-�x�h�Uf�������%G��/�7��]^�%�FRQ��{CopQ�M��iU� ���9nj�d���q�5jh��J�*�-�a���R�r��_l]7��'���;�	\+�M��ȹnvP��r˔_Iqak��Y���S�h���c��wb��uf�v�����#�+�S�&��C��P̙��¥��u���{��a�b��W:��U�K�9Qb�.�ɘX�(�/MA/��Ϙ:��X�%;Wm��\r�1��J[E�W��z��k�L��Ы)���ё&v�k_R�L�QU^���f]Ǵr�a��1���k���n�����KF٩d�:-��
?À�X�YY·*^r<���7�����mk���Y��L���\K)����/����V��Q\-�n^�W��t�w)Y`9+n��Ǖ��F3�s���)6,�א��܂�&��K�L�l;XеQtk����m�O,�֓b�A�ޖ��N����.!Q�F�^PڵϮ��nЭ�=
��{}B�.�8�N����BW�'g-���b���h�f� v�:̅s&���e0���\�t��͚{v�s����itiӃ��qZ�mM�'W'S�N'}[}Bї}q',d��4��d����wR���oNS���A��:']+��R�v4&��,����w]�<�3�b���.�bvf�)J09����c)�.:Tƴ����hS�kV�71mj�������{<
��g�'�����|R�j�;�VTے��2�,�m��F��:ytW%0�z�W�h��{���78uax��{��U �;K����x<�������bwU���*���I!�ͧ�F�g��E]Ay�S�ukx�w0Waf��U9WH^�mkϢ�ڷ��9�{�۶��z�����}�>�}q�}�Lk	�V��X����o�����X{]5�C%fu)̪E��ΗrT�f���tT�I5&<�����Z�5v�5;ԙ���vW#����g�x�4}�k�$q�ӛ�\��Ж�Y��m��ِ��V���:�9�91����sk]�Ӣne˷;��ah%���(�xةJ$Mؽ#9���SP�͏6��7��g�]�Ia�=Q�(�]*��˙(q�b}�Ѥ��}V�P���J1�е+�Q��n�9+�Ef_I���x�lU*]I��Ž[S�uk����:C��4�$j��,b��"��Y{��"չ�T,���u]��A����.+�K�o�*J/�!|�Y9(�L+�W9Dh���Õ�QDJ�a�A	R�B�.d�g%(�Uf�G9UQ�t����dV�Q�(���:��TAZ�U�%AU��9�VaF�t.�G:a˕h����U�Ȉ��dh��J�Mi(��r�p��T(��
��\�3�sd�Ur�j�t"�kX\�9T8�;(���!&�9$Y)H�Q\#09L�D����]՞�:�8�A'�۝*P�-I͹�"�'t���,��+�zVS�zF�KC��Z�UH�R�Փ�d��'D�W��չ�#�\�I#�XsD�'E��u�ZI�QaC�����n!�G#9HAz��̣��Z���҂��u"�ZF!Ù�Y"IF����Td!'1*�Q殮r�Uy�OP���D����k�݁I��'v��!'�
���@��9TJk��G��EG��V���IS��d�d��Q ��h��;��%���v�r(kU�B�*vf�L���k�J/��p�h��L����4�d�gV�t�+*+*ξY�����1R�Q�ޘ���3�p��k>�C�j�5z�e�bʽ�cث(g���h�tW�9��mW��v�Sa�-�n�o��՗g+�̨*�/մ{�>��{4��[�,Q�2��=Z��ö�Lim{���W3��߳��fG'�0_8*�j�\�N�KAk�ca�o����)_@
v��#f�T���!L+Ոt}������Bewq�P{�z_���i�++)�0?!<�0����i���� ��#�'�c�3�0����c��M���s�aK=\��oz���h�0;yٔh686�v��b�;�j@�S��F�-�_<k�\f����r�

{��0�d��Uyzܾ���UȎ��]p�^'�Iz�!=�V�ʇ,�Ȅ����b�P�Gk��yDf1��]Ӳ�g�����;Ш�{�Y$�Ϳ
;ΐE����8��s(�f�@)3=�TWS��o@D�})W6>F��p�}��V���˂I��r��;��2��|�	���7���r��.�-ĵ��*�w[�2I1[�հ%��S��r��[�k�i=Yk������菾�#�l���|���ӥT�h���GR��N����\�|]5�yUm��v�$�t�N�L9c��	�WA[�o�V�r�N��[_i����FdI���f���	��k�o5��t�[A۩�ʉŮ���&�3� cg�f�|�I�ɭsuֵÚ�j�yU��}�E������NV�c�ع�[��ut����ە��^�-q�f�_8��4��~���,�*q�{[���yz��{���|��K� ��t��Q��śY�o���lj~�T=��ݟ�Br���!1ۅD��B�Zlc�\~3[=x��=5ޗg$z��=*�{�m���P�F�c�d�5c�Ț��.�6����X�1w)��sҲ� ��_��C��Ye���y�LgbkWHƳ�b�w�3C�`k-6��'�k{h�Rf
�Cӌ��'׎���7���a�h�WY��B���:�CMM�Ǿz�_�:�m�	�Q�s��V\�rrˀ�<,��&f[w(H˱C�����r5�S{˚=Z/hױ�c����X�%����\�:�Ɲo�N,���G}|J�N`s��˧t�PciY������䆔�1�����9R��|�{k������Έ4�@�������D��������]q0�BCz����KM�U�����S�z���ˆ��W�ysj1Eդ� \_������V�k!gtb|h���by�t����t́�y�Z�x����̄7���Ȇ#��O:3��W]X��b�V	W�5��S]v7�Q��D)���h	���K�pru��kU��M�z��qO䷦�|�����;�P~����ek[�ޫ��!EJ�MrP�*ͧ�r��˨o�k�bi���&5��ȵ�2��`����m�-���Q���ԝӋ��ㆹ���6�m5�Z쎱l�Gd��
�xK�{I��������%fTO-}�w=ܛ{��������v�뤏�?9u��͓��� �N�Kyշ���;Z��Q����A��̿:����Ú��d1gme1�B�A�sm��,F���x��^�0�l]L'���Xy�r��y����,C(y�N�����cm^Ȍc�L˫�'�ϫgV�rΕ5a&����%,��o������Ԕ:�8�.u��v�1݇ȼ���Z��~��������Z�P����Cj��v����P|�����,f�o���U��g��^� �f�j��2��u��5�5�Yvr�xf:=j��זPC������i��q^�}����u�1_G$ؿ�7�{3~~��J��o(�5�������xӼ�tl�s�NO*�P���R�����_=��g���s��I`���m���9�'��v�R�����=Z�p�4����M����{ܕ�o���PɄ�b}���UW""Oj~�E׸�g�ǈo!�ҏ�h���&;>�&��wFQ�I�������!O'��ӓv;�NF�q|�����{��f����Q�B���CKF�Ma#4�	����q/ZU�ә��i\z�|`��c*�������\����쁗k�lꞯ�ʞ���u��Tr桾h&*22c�n}����U�㚨T��v��&��Y;��&,��bFr4(�Ǐ��W�@��6Ի܄��k����>Y�y1{�&=:d���i�H����WP����t`ך���Y�5�v+�"U(5�B�C��M��:jL�a6����ט6��loRn�\9�8_r%*��~�������6�L�Q۞s�ޚ��v�����_C}S�0����q\;d�t9{}ԯ��es��C��6�̸��{�u<|ک�X�K����X�6I�կ��0�3����Ww��{\ކ2���e3�)��;�rt�i^��qO?�P��;'�\��}�L���2���\C�����.{ժ�65w1fs��%�k#�w��r�jXO��I�	l���ǹr�8*�F���e�|-�>��iڙM�u���͇�՗g*9��7�@f��n�z^bP��'�U����)�g�܂\��4��{���x�dq�<�M�������r��\�DN�J��Q����oq�iV���}5�*紪>����{��kڄ��2���Z�$�.>��H���V�'E�s7If����O��{pkz��pQ�yͳ'���W)�>v=jwMía�D�.'�(�Uv~����5s��*�uXo*��a��ѵl�>�C�e�15"�Rd/k*c3h��'W�VnC��}[tb;�V�:�,�3��4���Ô��9��nb��[ �5�X��e�[i�밷���>����������H�������m�z���8��U���󿌣A�mW�T�R��#��\%ٹM*�q-�-�\sƻ#\fն2��B��ﻆ^l>;�H�ݶ�cK7�c���/�Bδ�]�;ո�����Ye�C����S|����g��
<�j6�=��V.9ɥhN�#��Q0z����n���Z�����C@[龥�7ܝF�v�K��q�O+B3xg;�b]�yc��#�Oh{���t�W@�R���]yz��[�v�e�Q�n�[s}�nꕜ��n5�9Z��:E��O>�̈�Hn�X��2'Z��V*q��_j�V������m@��<��]�u[����{ej�K��?[�'�u���F��u��c��/���]{r����S��_�ע��^(_�'p���nu�YT.p������?mK� ��?�LJg2�G3{nZ�1�8�N�x�a'/�]�LzȖ���m���A�4���+̦��4_9�L;�PN�i�e��wܪ7>�x^җ���a�ʔC���[�l*u��0�!�uKt�2��0��ݘ��Z�*��A{�c��DG�]\8���l�^�.��C2����D��D��^|���ZlM<YW�ݰ�����"�8|�������1�P9e��=�~���_A��E+ ��T�*�g.��m���C�����<W�s����AB<�J>w��G&B2��>�wS�5��}n��;��z���P�hP�$��2+w�w���!%2u��Q�i����Y�'�j��m@鍭O`�7˹ҋ\�tTk�+�:�KMAI��ƻ5�m<㊡�"�n��Wb|��N�P���cԨH�|���ub|C}�����U;�+`Lf��y��갨,�o�r����%!�Rѡs�����֘bf3mi�������:��ff�1��g��
M�S�g�B���h5G�]3�%]J��V�n�e�M��Q�.;��}Ϝ�o���w�7���P3�z�պ�U ܥ�>�	㫄A9�'E�����=V��1����ܹ���=F�۷w���^�~��K�e[QR�͈L�v�ݵ(�!jV�K����U4~�w�']j��\{�87�2������]2&B�KI=w�H��d���=���Ԩ��O�gm^���u�MG4��n5�	�/a�Tk��A�q���OC���@��y��^��Ska'S_,p����^��V�7��)�)�6يE�z;��{�3D�ʞZ�;��M��r�����@}�øX6�k�Ggr�}ܳIAl_:���}BV��Ory��b��a���n���?'��m������d9�ꏮ�ge+Xꑟ����oY�x�L����P�Z�M��֮��u�Y̐���n���4֘���o����s9��J�wz;cc�l_Λ�=����+�����PR�g7����A�Y�Q:���=_YHR��/����o�{&�<c��V��)T�9��\�Q�H'�Dw�R���q���zˌp����Q��+.��[�3�X��As���72���e\���heGQ.�̭�����cs%9�t�E�bW.�B�Y�����k!C���-v����]*�{n\��X�ǜy�s�*ԡ��u����w��49��;;��&��ӵ@md�C���Iۜ����*��ۅp�أT��UF�f�/F�1�,�8F?�_W��]�?/{�Q��v��\/aJT(w|�/�a��%q�X�{U�"�����R�)$}�i=�+}��f�[c+�(�!O}�&CKC�۴|�3���qsվ��G<��Ҹ��R��BleC�f
zBP{\@��A��{w�h]�y�{z:��z���9sJ|:As7���H��͆��u59�6�+���5t�gy5�t�T�4ø�0��W��Q��Ʒ�Ĩ��y���"����IE�=vکUF����|�3mTfK�Mk؍%힭�9*�2�j�\�T2��Ë^��o'�Rם���	����s���uu�-p��;p��G;7_k0-�@�U{�j/)��R���-/9�"�I�.���2��q�dk����څvn�P̨)�2���`�����ýo�go3�v[M�
!֮��v�oeQ�&�c9��P�����M��&�U��C���o)c����M.=5�B�x�kz`l�_�����Y;Ճ���S-ԏm�NV��l�X�%��L>v�����-����t�7yY1w{�q�,����R�O"��WśkV��
Rl9w���J�����o��k�捌��T���fW�	J��1ېmT���݇��%��j�n-[ܭ岭�[��\;�����Q.xꄰ�m�7�"yn���S�⦍��ݩH4���mÜ��w+
�/�@�G�U�Bet�3ȕ��z��Q��KZR7m�h痍���I����b*��=Dzq�~��-���_d�z��o4�H�r���k���Qgվq��6��*u�Gv{�Ge���T�h]_r��%�5����5���ͨ��TC��v(���{yNҰnΗ�#g[]�#%��KE�imf|�}���Ұ�V�О��ڜZ����[~T������4_��,�ʧM����a�e͈k�d��]]`���竂�kn�fg�� h%k����=ɨ֎�B�5���0D]��Z�U�L�ւ�\k�q�P��6AN6�۝��{O�e�m�xV2tԵ�%s]�ִc��*@�MC��9�vO5�MJ��;,�ς[�T;�BZ�;Pvར����"C�C������Ǫ B���>�v��q�嗒������Z��-"nfKûoz�Ӊ��sFT��
%6�N�;/u�.t��|�6�@ÖӀ퇔�F�<\�)]D|�a��'y����slu��I�V\���B�	���V�d�Y�5�3vb|�zS����Gge��y��\��	äW��8[������SE7f�d;�W��U�J���|�4Bp�w��p�('�#��Pu�sQ �軰��,f�s���Wn�����\�;@Ҏ���~ڵ��Y1�-Y����QoIyF�4���1�%V&�x�䐢�CV1wt[�)�MJ�C��Qt0)�L��j0�%],C�p�u%� �x^�ԇWi��M�aC$��A���J�
�j}�/�rv-�?[�F�ul��i�d��uo��8�)�6�Y�mp��c���V�K&#Z+3i6h�CS�O8"¶s����vN�4���Vn�� ���v}�YvU"lN�"���F�7z+�����\q5GW�(����e��)�6Fέx"K�i�9c;y�(�I�`� �f���Q1�am�pJCAk2v�t�
�ķ(�T";Y��9��;	��]�J��Wev��������%��v�+��`#m�fm�i���\�pۼ�l�&#Qd�/C��ӡ `=�}X��qd;d쮒'�WR��r�o��:;������g�C�2$���}��8�E����b�u(�um�9��ڻu���aT�5�%�1J�4�{�>���ѓ��V[ݼ�"��ݮt��ͫ��T@T�+(�ow���nj���b\fn3F�k�>'�&�d�Ju\����5o�\)��຤�Q��0*���tsV*^�d�6�ĩ�k��Š�6{y]��
�ý�etMa�r���ZB���5W��EV�,�D�$z�wqo4j���]�Fat7i�d�W|�8й���
u�:s2۩
U��B �}C�L3�8��D�yB�(%&;s��6��͢��kEk#��g��xh�$�Dt��f�H�F���J�CѲ(3Ywȹ}d�9���$H�!�f���T���nYNaU㓃B���HG`�ؓ�����^7�e����LZ��,���������S��P%�+0TN�d�]�P��q���`�;&��T)c�:�q�{D��-��Ʀ�wq��hy(yf\�WK}7y���Z)��a&�`s�=R	.2��a���X��,��vε��ixr���$��<�ucCW�P���R�O���5�)�5̸ݒȧ���Kp΍������N�����v��ongtة>�A-�5|��]�]�C�\�F����A<\�(X��̱��WI�8�R�\w�-|
�*��+�e �Y��ӱT6g�����q������ʊ�a�RL���J-�6E!%����!�\�ڹ���:.�]�7D�UN�h��!�*�X��D��8b�t!]ܧ(�i�B�%�(�UUB�TQj��T�"!�\���JQZ�j�Ҳ��yݺ�D\.�)k0��QRK�**L)-��X���T"
�j��\�I˅Ҩ��+��RE("E�,�"���s#�NlՔ\��P,��]5JBB�\�sR4�(kгTDa(jy.�r�*+�R����%2�JE[4�L�(�a W,�Nq:vT�ӄVd'C���Ω�d����T\�r#faj\
��=S���shHTr�	��(�Vi�3�g���J�U)a�D��l�VU\�D"�Q�+�:
�[=�8�U�u�#΅����H��(�!qK(&�Uk"���I��*�P�K�n����Z�.�ȥK��L��W)(��{v5��<3	��s{�PtYy���ԁ����c�P#J���R�������W5�ϧn+��MB�bk��k�k]��tZ��;mS���D�}���ҩ�qsu�%b��[Q�դ��sm@��<�tkXޭ��3�<�oh��M�	*�Y�<�n�k���s��\sY���ܨ�*ĺ9=��=CQ��2�9��ͽ�)�T��)�o�vg���ӶV��9��BЖ�X��Cw=�SH#[�l�9e�x#�Vg�߸�� �{˖F,z¨`j�n��N�g}�/W�<�zU�=)�_��^�o;��`WWugZ��s����qsErM�C�����<]�u��r�zx��ݱ�_9;#���S�g$q�R��د������I�و�� b��Ztļ���[y؟�]�����ڢ���I7����jOl�P�7��\�?L�,�]��5S�@t���P]u�KHIێx�dk��LS;$��~�ss�ʝٖ7�<����5.�U5²K4� 9ˆgJ���ګ�tdV�-�����g Q�^9�6B��izM6����[��V�5��!�o-Zop
�˃��}}�DN��s]mk�{K���*YR��x�T�|�F�_f.����U_U�aqO)O�N����J_	A�k<��g���<��=���'�i�Kcw�^����p�o�,x2!��~�?WOTU{K�eL��"g��f��o+���<�Q	��,�ȅ1ҕ�M��TV����v�;���58����^��Z�o�9M�h;a�#p��s`zl��3�S��6y�pr�j&����wڙu�}S\�ی|���[w���;,��jh[�-T���e�7�n��U�'3бm�ڌ�.���m�Аt����ÖB�%_�dkَ���ʓ��z痧06S�q:�޳�3�9`�_�sgs&$�{o>��~������v�l�-9�1'z�)$���湥ZUӎ���5�Fs��NѾ���=�"np��U}��#D-�]���.��m'�e61֭]��^祤���hr"w?�t�!��� 3ze��we$�X�adV���i����}�~�+�U�dW�%暇,�Q>Wu�����.�x���u}]��OtI&�ї:�wI�<;���/��t��&�,�����%ƹ�)(�twz�֮�H�fWSM媛�菾�x;,�5�̝���@���£�0�*9&��:onv����t\U��Wlvƕ�(�|:�@-ԗ�:�+�3����B��/����g�v�.q��W��s��(Z��ʦ�n+��_N�*⒥��硬1\. ���E��F3�Bח�
��rkN'�~�h>U%.����R�2N���lt^�YQٯ��{��o-�|2��_
1�>���&4$��Yxo!�m]J��Y��j@�S�wQ��u�������8�S�w
$gO,�bg_t���,�o�sؗ"�W�w�C��NY@+�I�fj�!��w<��%�5O���7Q��r桭	�h+�����I�ѩ;'���+/N�@�V^����7��u�P�T�4à7���ٵ����o��[RY�W@Ŕ=����?v?��Ow��!�/�OocQ�r�X��v�&]�ރMM�m46��V��;S{�V�;H��'Tl�q*�W��%4�$R�n(��k�/�t��s���q�jƛ�ѩ˫5�a���[�5�3��Ol��t^��Spq�EǮX���%(�7e(���ʃ�34z"��gy��uL��)��ۍwL�5���Q/�^eD���7>n�|c4Ѹ7Io9Ty��_ss�)�<q���s�u�E�φbo.tս�$�{�5I����\�p�^�N9�r7�檣Wj�v�O�R
\�9����}{��,f�M�����je63�Z�ۭۈ}�^#=`c��H��Km?G���ݔf�P�e^�eY���V8�)�&>{{��v��/���lr��M�y�TgY�c�*����;��Ɩ�cc�a��ݶH�:������}i��}��<��wb+@���S�/k��A���K�{�����9���!�莜&�\:OD�u��@l�P`>U����<^v��nv�TK�5��{z᪈�)>[f��C�#��5��w�cf��nv���T1�&Χ�襦��󝵪���T�K>��pV�Bߣ�ۣ��Sv�q`���*��3]�U�)Q���++���/��f��%��-����/���,{+(:�5���F�����m�Ok3�4�!º�ز�pZ瑹��)\��M��S��XJ]\�X5ĳj�>�+)t�[ϩ���w������J�g��G=��k3෪1>�����q	��kg�d�P+v`�y��&4FG��
�_7t 5E�#�Љ��ўs�w�n苲����ޱrs�"zm{���|�Ȩ��(�{��nzWf�&1c��vc�c$���u=�8Kzj!���̽p�2�1��@.~S���DD��V��Y��Vm8�[Q�������1)���\ƺ"c�فke	��[X��6��/Ż��o��}����٭�_'�Z��2�I�5��Պ���z�ө�+9������e�Uo�ګ����C'\1�*�&� E�Z����y�S�F���9H�F����ϣ-�D��br���P��s�X�����T8�Ԃ5�m����#X7�^�p�"V���IZ���>c>u��]�^��<&w�;�\��>������h�P�ю���t�Pi�%"�47���h�e�*ݠ
H��<&��R��w�@ד�@D)����ɭ���(��P�������W���������@�ř��L�Y���eRT�u������U�`�E�3�VA]y�����p��Q����ڝ�T<	�|ӇM�­ݶ�W��v��vb9�$�ejmI��G�4�O,O�#9�.P��N���<e��\:yFrw,�khn&V��D*M׺zV �E���[�Tx�N$�c��F8Z�y��e�ո�4�gWcP���`l��L�OH{�����mhW��Ź�[�\�`v�u�V"��|q�Pߞ����b�O5����d�)��i��V�s/�`�Qt޼�vT�l3K�h@J\3����/Q�]�IWqoU�߱��U$�)��h��X`��yN��B��J���%[�CCE������2=���}�������o��H&*�?u#��v_t�KĖB�&��v��P�����G������^�T�G4�Cn1�W5$vj͛�e���hz�U/(��y������UI�]��P� �Q��)�^Ɇ�Tʚ��2K*ˇl�\yD�VA�췜�Ȟ'������r���Hn�QP�l�:��
�dV�Ӑ���N�^~,=mT��H�����8n��wh�q��J�ѭeu
�Ϩ/���u�[� ��*�<'f�.�[,=5��\I�p3��*��'���Zځ�%��N�}��F㰡\���P��N��S�]�^Ex�;�MCg>{r�����ٹ��Atỽ;V�ਜ਼Zڡ�>�]p�^�r|�F�P��_;F��`�G��8�H9�3"��d6���X�N!V�/�|�Sc>u;WzC^�� ��l��e^��C3�C�r�� �.߰��Lo$طM��io���$Ԟ�r�n�z'!�W�����Aق�Tꄮ4�XH+[jm`�,�r���Tp�
��ta��ڟ�٘�Lr�D��:¬J��iouZ� 4:�n�n�S�k�.z�y�kz$w 6 (0�D��q�uy��۰��\��kU(�ﻳr�C[x�m��+�����g��Z,o^��J*�;^�T�s+�s����o;}��f�b��)HW>�����O'<�0�46��gѹt��y���%i":�0��M=��5\��k�t��w��3q��춄+���P�Yfb�R��q#өN���\�F9�����c����_6�����Q��H
��!��uru���m˫�2���䜾�V��	�����9v�M+�_��ؽr̕r;<�7׷֟���!C6��������%6��o6�7�ä���%ă,�u�Iut�	C�Zev��P4��j;#V��^��^�^�ս�A��٫S[�25�5�u�q*@;� s��-̃|�9l��}|C@�s�.��s{�n!.���5-���κ"v0���u��8��,�z2F�j�7���Wec�������մ5;���f�X������-�5Y�弥n&�v�߷[��u�9{4�ϵ����J�4Tq�N�4�}�ty������v/�b.c�e��_e�v�Z��ns 1Sں�l�U(��Y��bO.��B���"nr�Ko~�*�� e�=MY���i�(\m)�ջ7��Gv)���`�;_N�{��{���L�Ey��U�{b�E7��y��/k�_!jp��r�Eu8);�����sm�lR���V��g��a��t;>��v�Y��w��SYuqCq	LI6�c�hGTf_ʿ�@%+�+�w6��R��I�Ӎ�	���Wj[����ryw�zm������@+��`�'�����1iZ�c��@\qݴ�4�OWp�|�<�[t�7 \e�g�C�v����m�O<;���U��[��놪-�ʄ�m�J�`{i��<��{�'�?l�{��ЯD�S	i	;�k��ڷ�m%%��.�����u;�����1�"H�N���}A��t�]9����*v��c{��V	�s@/U/���$c��Ϻ3��cG�Z|���.1��'��9��v�n�c�l�6��77ԻV�L�{��>ܨ��p���ִun��Ϝ�o�a��"T�1�l�.`eb�)D�

:2U-X\�7Rv�)�{Q���o�j�~�ޥ�6�^��k{�siW��v�������^j�SKRu_,p��7��q��̌WLNQ7cbrGR�^��N�f4�IBd���}����#4dM9�����h����<h]jx\T���ڵc�F���f��MͷM.���l�N>kB�t�*�uN瘮�u�!��x���f5i���I��s�-s����Η��f'Sc�C��*��ݖ��~Jyu��^�(Z�\R����J�L�̗/[Xo)U���G;j�m��y��#-�Q]W���4��;<%���U��5˳np����Z�H�/�Z<.�,��S��K���v$l9��]��O3o>�^�C�U���{���ir���v���puF;�GV�G4ݺnvF����!�Ԗ��c�F{H�J�W��r��N��uC��v�<e�&�\:yFp��ڃ���sh��kQ(ӊ@)�����TmQ�i���e�c���o@Tp�:�۬o�����)�#����{��\WPu�����};#F��>/�>�Y�I;��O��^���{;������"�6�&s���X�\I�`3�\��_Ƿz�
�nBy�m��(�#���~2`�����xC���&�"���+j�^t�\I�UmM1�}{-÷Z�S��p[Mmp�w�f�rw��GC��\�-��hв�e�)���j�,cY{c��3/��!h��#
�|3"�,o5l|d��_,]J�q}������$�[V�q�)�������w|���Zrm����}�l��#�B2uwM�M֊u/�4�҄L�b��)G6�� �4Sȯ�i�
��#�'PFQm�@���(��͇�ZT$�]l��ӚB�[��3����X�+��K^�J����n��n��F�(.� �+���P��կZ������`�i�*��Σ���q'|FX���&<4���ђ����4�uJ��H99L��5yV�S�ͻ3-W�n�g��܅2��I�V낔7�8��S4/2��g��-{���;�� u��q�����%�"@-7�]Y`�8��J�@�WY�l���Q��/T�Z4@jQǵۆ�:��ү^M��ޭ ^T�J
��V�1��J�hn;u��m�
�c�Xl�S;��Ӌc)M��s��B����PǙ�'R}��CjL�Nۻ4�a඄j�+]E�a<c���L���2����R��gv�i� 	#(�E��{a!��u�5��P�ĝᦗ!��m��v�rԡ�K�7�nLq��L��.0�2�w���a�'��v�V++^��Km3?�9��}˔� J�Rd��.n�-Uً)hVJ��Nl=
��m�i���b���B�Iʝ�O�:�=���U�7-����M�v�pjK��\&�\��ջX�ެa�moE�F�	A��[u�[y%
��	7�Bko�X�����j�3cG8ͼ�Yʵe�0L�u���B]
א�Xs@�@h��&��j^s�U�����9�@Q��W�i��l�����r�9��'$����ZEo!�f_$z����+S����uW,8���X���A��wa�0P�c��:6�g7��Mݬ�ڊ��ևp�鯬��+bq�g^�8mv.�!�!�8�2�7��,�Z|A�Y��B�Bѓ�-��u��b��T�F�p���}���U7��k��݃%���]#��bTC;�k�:�����R���:�e�"u�)gf��wa�B��\�j*�шZi��^�$n���"/�v�n��p�2]���$�ǏD��k��+S��*�qNa�c\q�!�Z��v��4$ ]�s���-�ݦA�}�;kgL�UGY-�Q(����/QMԎ��2�⻾<��zk��B$)O�;PWM��j�M�ЖC�<[՗�N�Nw2Rˋ;7;kj�k֜�4~9rA��԰>yv%LB��p��53�q�ާ��yS���)�A&�$N#2C{�L:�uIqԙ�իØ��k������ghm��Na�E���֪.
+5�-�+(�]���7u�Ԃͅk�l^�~�h����[���q={T�a7�¤�(P�D !G.��.u�W{{���.���*M=�tI&Q�Ur�Dʈ�5*I�A%�DQ��a�J�$���Y&BjDU��9!DQTW��iԐ�"��FBW9��d%TJȳ
*��0�R�:r����W#�&T�\�]�*"�9(����U�й����9n㙖�]tp�U�����AE�J=��r�R���RdW�ąi���bҢ4Y�EW<��'tIe�Tz�Y%�I�tOS2�Zt��;��
5=.G�"u
#V^$E��],��"��,$Q*���r�M��z�*rD�3�{���;*8��%UȪ#��B��n�ETQEW"��EWn�����w3���ǿws��9���3����5����[bkN���@�xbҭ}�im<�R�S�p�1`������܈�r�(ݷ%8��T�+����=�N���I��t�\t���X�S��W����� g����ln���5�?���q?*A�n���{]���8��P�z�ork��z�}�}SQ��n1ې�28�b����8�k���l��m̿J��ѵ�}
�G�|�wx��՝(�9����dg��M�Y��ި{�3�^}��ʵ���H�����ޏ�7��)=�R�^E����%�^��}����*����Z�nÞ�eU��U�pz�5�5pO�InO>S/o������6��u�w0W�	�������8�w�Z{k��r��:�E�iڙM��֮��I�24�+��ę�^�v��pv��E�T�	P����G$ؿ�7�{2V'l��"�h�v�!���|���:;U�t{7�U���U�Rm#o4�3�����1�B��]taM8�yU����f�Dv!�N�riն)�S�5vIӧ�e
*�Wv�ck[����	�]ȱY)ř�'N������͟et�sT�g>YN,�'n�d�Od�Qb����(�u���.���'bι�m==$<�̳ձ&��rx��ݶf%��y��R_T���c˴���r��%����?v�����"���w��h��S�)��:y�p��\N�i;��m�c��o��RU�����uFWvgwq����D�^�a�<��E><[��o�!8ͫlc+���p����r�!�K�Dd��
R!�HǻA���ߌ��Cڦ��pϓc.��:�d��E4�+��Ш��2T'#A��f�6�=Ȁ��kM�o6�|�}��rs9�傒�淊��Öo�;@��i�-s]K�w�Q��ĺ�T�a�3s�yU�f��������2b�Q�w0V�|o�RwJ+67��%o3=+���W�����n��5SK��g��t��*�����B�ѹ8�]*e����+^j��W���-p�E�޵�eʭ��o
\b�ze3���6�5}�(լѐ �ؖ��h��yЫ�X�-�ܫ/j�Ӕ�����ʮ�ܫ�6�����`�}�y(M�<��F�X}f��M����r�g̸�0s�,�󸰡�]���T��s��}tYV.]gcQ>{.N-h��u:���s�؜k��uCܫF�B4���E ���Q��3(�ͽ؁+^r���|�L�G��r���]-Ԫ��&�m��˳u�fV<�^�e������ ~��(KD4���q��oG�w��?F��������f�;���������G\(3�F:Z�*x�&�!�j��۷�=Y�wc��7*��>��Ҳ���N��m{�E��u�j��lW�X�z��{��Ҁ��_p�{|�<��{�*U�Α�/�,*�J�}�ۈ�e�8[I����zvNv[���bq=��6�
q�S� .���]Aԥ�$׮3a�v��K����)�`������;�(�	�_�p���/��7��W���E旜'u<Գ�MۈKtW���QȄB��)h�+�d@[�8eT�{:b��S�U"nE�'jgP�q)�^~��#�����k:h���!�Qqe��×�Sٜ��v��02�Mۉ�| 3M�����Թ�7�5F����^�Ȩ��4�6��%����J��Y(n:��Q^�49l�Of:&fo.VsJq�y\z�@y��m�T;faх�ƃ��E���e:��%sHK&�-q���1�ڎ\�|;a��\O�.����X'�SY@b��C'qs΍�7{57ݵ���˦���䘚mƻ
�u�惸�&
W�T�ԩ��J�[T*��2�ڸ�[�i$�Z�
[p2y�We�V�f(�:��R��D�?{A�9��oOn�F_�V�=���ͽ�C[�f���`��N���yU�f���úe�P�ù�OI�Ѵ�����9�LC��nd���l�l�]�AS��C�y�bUnS���lw��h\3FC������ld:���k����ts9�ʂ��B%�
HL�̎V��'\��@���£�
b��[�U۶�*��;3r�Bc��!�J��j4_8*��$���p��+��*��o�s�U��c6���B���IMA��3�m�v����]�;�zt�d�;3�)k}��� ��mKj�ަ+O��N�)7���c��-�XulPE/,������\z��Gf�Fe
]ww1P�ܦ5aV�����Z�Tb�*c�3���U�[����UF2qm�K��a�s��>���{O_�\[��D���{��o/5��V��eu�.rSW�����(��x0;��te��Ϭ��eȌ{�s`�]��Lc��G0��J���z��3��\�0;�y�Q�D���չY����u��A��NwQ�to�8��leC�g�B�ﻦ�U4��'p�"�;���#h6s�0-�]��4��J��M��,�Ȅp=\gjUȶ�;��v0�-)��|�j#�� �p���n0�|����� ��ӧ�'�6����D������u�}SQ���G=+g��Q�&n�����C�p1g��tb�<���(��<��7��t�[�FQ���Ĥˎ�5�6�]������:`Z�}S����{m�j��8���7��w��W*�x���z���x�5�d���u�.�m�iV��Ĵ.�-�4��3g�w,�ξʤ�f����[�%m3ugK�=�6ri�J�X��P�tx<G#Xv�U�c����*C��ʯ�K��.*�K�}{��B�騴��yiSJ�E	��L�Nļ'�{O3���Pik�5���"�jX�Ѹ/���q'�Nr
����75��\������k>�7{��.}i��{2��ӓWd/���pډ�ʉ:�^r���)��s�:�ļ��{���Rn�o���7}T^؎e^�e���V8�]��8�6��pcdun�o����9������U����TN�J��=QR\��UZR��Գ���^޿S��~~Zu]SZr���s ��ꀃ1�3q�Tmv.k$�����Z��^6��t�٤�n ����OQ��}8bp�R޿�9����;+��4�Iϗ'��Q����-��0;���;�\%�8���MQ_uqq���8�[�P[��mj�\f�[c��\�lw]X�-~}�n�9�I�����Y�oTb}����[��3B�xg��'��cD��n���%��yK#��Ό�|��+ՆCX���=W�j��9��;���,�:����w���ń*FY� ���������U��l�W�e��a=�YJީ2��rLz�î�}[���2;1�C�]=}���ԃ��rs[��=
�h�ĥY�Y���
Uq��(z�IZ[#���;@��;�yo\����b�y�fg�%6
�=q��Nz�b��u��z�"Z�9��]ٲ�|��*��(��6w��rn��9l�tJP^ls�Y�zϒ����C���[>�4o�����Tq�̚��g��9(r��2��ݪ�8�\����*>����:'WR����yp���1���^�y�`��e��3�z�\�d��='��)�m�U�'�=1��Z:KӂW�I��Lz�n�xb�ydg��Az^�z�{�����U�eQ����w��ט��s6t"s=�N��w�VW��u��j� �����31�V�G���7��۳Ͳ?v��^��a�۹c)�Op54�A}P�+*���2�^@q������Q�w���yڱ��:K�'���]9�n�Y綆�r{�|Js/|g�ת�����4��}��~�qg%}������������q�~/>�+��^�bѾ<.�I=Q2��jrb|%I�Tȹ��;�c=b�S)�Kr���	��x������~�x��[��g�o�|�a�K���gv�j��*c�/��/%���9]��t�#ꇎ�g%��X���F�R��7�,�z�}@��Tw5b}Kl�/�;]к�Ds,V]l6ѩo���_WS`�D��h��\eD������SR�a���Ζ�Q�J�sl��o+�h�&�lǵ5�VQ׮\�� ����+O	*S=k(�t�X�~���7}!�~Uw���pl/	ܬίb����'M|ω*��`�J]>U0}��p�q-��b�יY���>3U&rEPv�w|�X������.\��%�D@�À�':ex�����~W�j���=�י+�^���e/�~�M�g�Do�X�Ir� 75���1-�q�Z>����T����Y;5�u��*>]ƣW�M�}9��;��փq�z��Nx�9�Z"KgOI�G�rz�gn��N|+=b���ϼn7��u�j�F�ޟ"|r�|O�́�i�*g���搨��t<�b���!*�}���D��4.+=K��%O�?L�(����߬Ѹ���;��.J��ΖD�����_?(?O'�,�ƪ�V��1F���g��	�4��o�a��UA=�Sn�2.XO�7t��]�ok}������H��4X������J����]�z�M����ԯÅ��߇_T:n�}�0"2� Z�5�kԏ�t<O�X�kߡV������<6�����������*��×Mu�����u�@b�piP�����r���^.�y��Q��F&G3�������9r&7�-��.�z�q�Ɋ������R�p e5��a�\qc�h�Zr�鎆�Q=K4[�������y�9��ۋ�z�Е)�GW+\4\�b3ؒU���m*��U^�r!z����wPu�_Y9'.:X:v��xj�C���*��!�퐶����L���F����q�u4�|O��<���$��������ى!?G�Z�?f>�b>�s��d�^>'�t	RJ�fX
�K�q	���9����ΕF�X�I��a2���zU%�p����ω���x�]L��!�����z|�J����)0:��ѹ�qw��r]�ȷ�6�T>ʔn"ω<?�*������]AWIe�Y>���P�#��V���'��uC�+�P�~�=�&炱rQ�E�U�O�C�[+�]��)������
���}��^o�}+o��r<�}@>7�R6�S��U���I`L�����\�����fը}���|�X�g�U�޴���?H�מ����f�s �JEz���`Կ]���9,�If�2=)�|e���:�֩�~��a�u�G�a/ި8�Y��fG��9'���_�����ژ�p2SSBպ^=�χ�|�F�j���ϧ-)��詺�.݉��l�z
K�r��יt��Y�l��i�o²ĵ���������~�X3�]Y�vT�{�iL kd2�����`�S�Fj�ǽB]��耻�wP�[�X-�|q�ۭ�cʹ]ge󽧦����9�)��Jp���(���D����w$/C��}Q4��OX���=�*_W���o��Lz��G���(��-�'���g�ս��S�'���j��0
��Oh2�Ϣ_V���^=y��6H�)����v�h���$����=ګ�p����޿���X��T���[ �|n�q^���������<�=��͑8�s�����'/��m���O�h�Ͻ@z�箠��]��g8�QX�M�6<)���N&�~�z��,��������x�ݶ�=����2�R�{޻��������gW~�5�hGv���ˮ�go�J�k�����<iФܜ\�s:X7<�<3�T��}u̬����5�Sf���K�(��v�Y��w3��'0W��/�ɭ7�@yf�`V'k�F;~���=�����
��%#�e�]xw�{iS��
��r����5�T�Q���P�	7�..:�`���1��rDm�/�Nw���������9\+��R6��xԕ�QUC�|����w�Ƴf6�H��%�q�}��O��}�����G�ׇdM��X��OTL��_��An*}�7 ^�`ї�)���������/�&�bM��c��;�im�;7qX|�/�b;ⶤ�$�
%�p���nT�fc]��8�^팙�:qF$dn�Ҹ���Z��`�����׸���6�;7�/--3q8��5�������w+��+B�Je�N��q�%����1#iS�9����*���e��Z�i�؅*;���aE���̼�v��"������W����Ɓ崻D������6����mIǛ<+u�C���ٲ�fyt���Ǜe��.�[����f! :�t��w<�4��`J�]q��c��W:��*ԗ���ƽ��zj��s���u��is{i�I
���*���b�wC����b�;K#�V�Nװ��v�!r$�>���LXj��<���3�Iu|��Ҳv����^E��u���P�BW[F�k����+*T37��9�d�|]\�0TF��g5���d�&��me=��X�u�c$�w�v	�fB�'�t�뱢�(3`u�ԯ��y�>'�[]vI;�f6�!�KB��̻�X3���z6^w<YCE�\z�e��ZOH�Ͷ�-�F��F*ã�s�g;-�% حQ�1�{�mI�g ��˹K��A��%�tdZA���A�[N�����v<3�ѷ\�u���k)���C�B�c�Z�I���S(r�;-�ׇ7���|wU���L9����#sJO;u ����uC�Jm-�ڵ����v[{�U��9��x�6�8�0�k8����M9����J�nMǔep�]\췚(0cM�ڔ�N��� <�5}2�lg�H[�{w�o�D�z���u�1a*�!���o5L�+�Ʈɳ�p�&��n�lN,�W8ވ5�F���Z,�)|l�ݲ�{*`ށ�
VU:�*�)f�����^G]�/_f�EL�p�u��7���^F��]�9ۊ=��&ޫ�{�V���/�9ə���Үc��N�oxA)���!�MC�;��U�QJ����em�g=���I�zh�9JJ72u�M��F�7��2[(���W.T�K�f3�j���`ڼti!l[����{��^�C]�1՗�u��'a�-F'���������O��S��h�m�٩8��C�*\l9܊�̧ݷw�`�[����]�-�}S1���*u:�0Ap �X�E�E��Η��Х��P(�J��"���n�qY�Ya���[�)��Z�̩3*�X�S�:�69ܯ�U�XUľ=[x�AP�2.��q:�i��d�rmfX�<���-4��N'��+����c�N�M�?i��BҙY:���0�D����cqIY4�Қ���Q�WVX����NN�ЬvPX�U�Sm��]�ޭ���xD��hA�/�Z_2�Ծ�B����Q�xa�VJ��1>��y�����Owy?�s񽔫֑EE�]rN�w7iL��Ԑ\\�Y��� ���v��d�s��r�)̥%�3�ru��Q�sɔ8T(�.�N���%�p���Oq�Y!g�e�#\�W�r�*���.z���P�Ua��7B�
�
!�ܼ�QՓ�"�h����ەҢ3R�\�nE	�u�˅�#��9R�痠�d�P8�y�c�gfa��Q��c���;������78�U��.�Y��Ĩ.P�dk����J��c�'���-v������]i�EW�D�:�\�=��;���AAAT9Xu4��t=f�ḻ��9�K5
�5ZD�%��u��������r�z�eJ��RXX��y�&�7	��rB):�U�!�z�Y)�E��秙��#,��	QE�Y�w���(�{-�V��!�	J��y�ws���m�o(/�t���/���)��ݮ�{�4�(��qs�<L��((���'���X���R�#�U7V&�i߸���/�Do�x����i������d��FG���Gf����m��&��7��,dk���z���}�CFB���;�{=ꃑh�����5v�<���\�j<��<[�"���;�<ƿZ3�y�}�lv<ܞ��U$��~Z�y�>�+���^��	g>D@n+��z�G�cSֲF����r�Od\g��^rW���\�W��&���Z�=q4�}2��Č���6�Z=V6�`ޯ1w
�ڃ���->����^W�6��@� z� �C�~uNL��Y<(̿*pj�Kg��۹#�����n�ONq�>�>���Q�������^&���z��dT*8��M}����p�G��l���B;�3��qR�迫}���oS�q�.7�c!���F�3���~��^ӣ=�;Qsz�jL͟D"���J�֏I��I���Lz�n�xb�yddk��s��<�yE1~�RV�5���=��b�y�8t"s4�/P��ⲽ�K�65[ Tny_��񙹯J�+(�,m��39���ׇ�b�n�ʾ���2�cV�����{����7×�]�Q���_Dn� �K��߽x�%�~���C��+t��K?�f��#igì��=�'�������8.\��|�OhJm��15C�v��MgT�t"j�$�oNϖ��7K��B�X�>[(e�Ⱦ,��f��T;�ʭ7S/īݮ�Y$+�o�����-`%��rW���;��Ӑ��}綅꜓������K�YQ�V�#Vc����k�Vz�ΕY�tˀ�ᾯ~r�}��~/>���ȅ��.#T�}$�+��SY���Ϫ����h�@�c�S<�.+��}���>����)�}�N��i9��
��<�5�u3�ڏK3g���π��h�u*��E��̷4'���G���77����T$�������^�~�ͣ(�s�|IU��) K�c�����/�oף4B�ѵj�d�Ϸ=��ԽXs��=p���6��;�rY�D@���q7�+��Qȓ>򩆽�q�r���Q�����J��0��#��É��z�ۏU15�K��sP}$L�\
T�K|�u�7�%��I�.�N�Q��o���O�����>��>��n=�^�zs�Y$�D��^�f��Y�����o[�#ӽZ+�R:7��x�M_��{��O�}Ӿ'��Qi�s�Wu�߼T�|!x��)b�Q�7E捾ꓺ��@?[ ��.�������s_0��n�'���X�A�ޣ�u�7����P�W �5Bm��Wb<�S.c����[���3�N�˝{4%��^��Y��	��Ȏ���eE����ѭ���]�Ԓ�q��F�_�����߫.6��*9��z��wF-7�4}����t�a���c��槣}	^�R=�2O��Q=C&=��a����dV��ޖ5G;�g���LX�H<���Vs]�KS�����b㽕 ��>%T�}t���n��R��l%~;��0���J�F�ֶ�V��X�5T��ޡ�K>�^���j���*F^�'``^:wj�Օ�}#w�{޵5���̃��:��4K>��}����ϴ�^��#���ۜ.NI��`��]��������V�f�����FI�O�@���q�=��t|�/���^u��9�:��k=��~훍��/�9��2�T	�u.���N���̰�^����}S�N��w��a.5��)ŏ��{��T�qe���g�*�,]L��ty}V�O��h�1��2����%�����R����+���[s(�����f�T��L�n+������)�ǖ;����;;��n���g=��?SҦ炸%E�U|f	>U��e*�U;��]���r������"��Z��仅u~�I{�ӭ�!��l�d���('�E�r�z��%,�;�uB3�IO��.�Mjf�KPY-��`��%�7q�i��Sޗ6�Ԛ!�66�@��z��
sr��tJU�������IB�Nz}]��O�{/H��HJ�3ʈ��S�H�H`5�T:���7�]�{������������ğz�#��{O��F��������3_9�Y����R����#����/�,ϧ���[���e�߃�F��C�%��1�g[g~���&߽pw2}�����s�tyᑤ�*L'�DO�W��T�x���׾W#m5~yQ�]��f�8�$��n�~�Q�+��@�=�&az��b�_W��d��yʘ���w#�=��#<lWNSd��/Vj�P�r�P��� ���R��C�g�QR��NV�����1����	����M)Б�]��?:�7��P�#޿���{V/��T�J|J���ߎ�S�-���J��'=�}4�ӈ������b~�Gz���L^ˠ�����`��BBu�_�|��wb�_s��XwYLm����7���vڸ�>�	�)x��]�����?��_�Q�ǣtu�IS�g99��=P6t;�����W�܈�L
������T��c�\��,W���I�v�2����*n쳱�؝pK�ۢp<��TF��0���.f�܋S�9�Xl����{�֗rxgp��gE�P{�>��U{w69��z�I
�| W��1�u�+�.A(ݤ���ս�Z"@�;��]��81M��ONl�P�)����|��A��ܝ�?A���q�֛ۘG��٘yB|��t�r��/�/������[����۴������u�����!�r=�.5eO%.�0���z��W�����@7��OI�ݿ���r;+ږ*��w���y��冽�Còr�R�w,�ą�UC���S'�U���}�+=x}�t����wp��>�i�t�������ׇd�pV���,{�u����7m���׏��Tz��WQ멟t��E���qMՉ�i߸���z\o�x��y\>ȃ6���֗�>�E�nE�����9��ϲu|�r���-�5�����}�Z1{}m�vd)q��z��}�>s��គ��c��(҂Ud��I�L�9݈x+���C�O��̨S9���-�T\���Kz��y��&��z���z�X%���0{Ӵ_\�}�G<�!t�W�#'=ڝ�w�1�O���}�D� zp2n=�V���D���}2��ٿ���2��Gq?�@��b��׼nFD�nt$���kˮ7�j5�^����R����>�
uNL�B�O
�2�W��EM�W�n1� E��ȻTp)S�����3ݏ��:x�v�޿�^�9�ԧx�o؃����BKs079�
+)j�7)��^�G��躣�q����9Ҭ]R��f����݆-&�v���M�ҍ��]��5�wat֧�޽��S<���������6v�,�A��~о�~�g����=��h�����@uB���.�L����?322�q��wԃ��/�Ps�\T�:/����y���}߮ь}�Q� �n�sõ��~�S�27��%#Ώ�Xg��U&<�mhw�O��N���<�n�xg��告���5�zs:�Q�;䵼J.|3%�>~�_��X��q�~�����$�E��>2�u9z�vuh5����׉�']�;yծ�X�*����������s˩���'0vQ�wYU���c_����7��[^����B5�
�7dZ�M��u�rt����B�NI닟��L�+J�&�1�ޓ��y.;յL�)p93�7��{�_��~�\?>U����Ʃ�<1�z�)�F-1P�Ԣ�I^�AЙ���L�L]w�/�4�>�q���9����dz�Ǹ^[�;��%�}Yس�<��ϰΚ� ��`H>E���K�"�Qf⛫q����#��6+2�90��uؼ���{�X�����\>���.J5����~"E�M�]A��|${/^+U�qn�o�o���@�ȕm�0���[V��u¸�-�h��_���ʾ�rƁ�.��YND(9���fm �����bw����Rx�I��spо�N9Z����N��Yt�)����zU�R��|+���dZ�BmvRT���.R�;0S+����z2u��W���70��G�T�V��i�l�8z!Өv.K5�"�0�Yn����ex��]G��x��j��N����*>}��n}�ay^G������$g}�%�\�B ��H}t�gGY�3��^��Gdo�}�:�����h�m��l��Ӝ}��Z�� �M��|�Ih���Vߕ��Yꑉo#iB���*H�ޤ*�]4xv�/���#Q֚�Q���>/����s`n�GO���=�����\��=Ǌ�30�q���nV�ޗ����#����f��>������^[����Ȩr��(2{`d��>�����>�u�7��Lw:�6��GM�#��Ypf�I^�CВ��x����h�}���Ī���N�q��7J_)���x��y�)Ѹ{�9w����C����|�W�}�5�}x��ЫU͜����!��;�����m�v��0)�#��*�קƧY:r7��n;m_���i<�Q�NDs����s����9q��ӷ���ͱ�H�moNg{�Y�!6ng��S%���V/;�dI��d���̬���%�w���v����Ѿ.`r�F�ִH�rQN��M3�b���ڜ�����h��D��)år�2��-��e���R�iXb��W>޻Zh[�8���-Dz�ɊSb&�t�r�v����Oz�0쭝t1��ۇ�K�e��w4���N}/)㌺K�c�2�d��D��Y.��4�yNF̰�w�m:~>�>�ۗ�6��+
����%��~���VT��R����2*g��s��ϸ��<�>�9����	����ej��P}a{����������R��`uA�~4eST�F뮠��_�>��{Gz���&o�#xoVk��;���~�=�&炱rQA�V�f	>Uv���ǌ��e�n��^yi�E��(�y��ܷ~ӑ�<�7��q�TF�:�
%dB���}&0�|=�D�|�r����:@�q�#��V9�uG�}�H�Nx�;��=��������f]�Ϸ��T���YX��}������#���O�����x�� 瑽j��~��dg[gO�@߾���:��l���� ����	��Z�߾��2+�\�B,:�}r6㒶+^��h��l���{�3��l��x�d
���|W����0Ӫ^��7T�{���Tǣ�uh�m?PZ�MR�H�w�X��u��M׉�}��7��w?]�5
Yle�B�����:��\�y	��s\��bٷF�,-:�������Q;��u[�w���m�~��4�,�WT�O����_ݍN�z�];�3{���b�*ֳ����(���bQS</wu�fkԮ��_mb VK:W[ժ��F����y^����Jżų	YRuY��]˿(5~��^�q�{�~�:�6����޿��Ջ�;�R)�*���܏��c&����7&�+'�T�z++��l�)���=�u���/� z��]A�����P.�z��ޞ
��_%oA���VSp�����ޗ�}��<�ϴ�B~�^/{�p{�J�u|*k;z���d)�>�?~���s�p�3����χ��l�w9GEԪ�N�`Tny�xd:���>��֧=���5<�D{l��Cw��z�m�ΝE��;��X�+N�^`~��b����<�=�G,��ګʆ����+�����g������*x�Y�)��q^�Fc�����D��/v�=z�*���2!������_��<�ԇ����P�*F�\�O�+Ư7(x#Gī���;�!v-:���E�(ϼn+����5��y�q�{N{�����Ǽ�#��ó��Q)�,j��g��$ދ����Q��Oඣ��9��WE�����CN�ǼG�Ӟ!����p��eC�kK�vw3�c��Ӑ(>��ʌ�$)^3q�[,dk�����Bo�����|k����_��7Tt������fX���Z�7u��,dk����~ʨ�S�wX�!^UH�Ͳ�5$�Y3�&u1A�x�� �b�α�!1n

pf�m'C��6�}B���\�w�M"��j���%k��}�r�F�L=_v]�v�e��u�U����gQX���PŻ��U�/��pv�T�;%��A*��ž�/�^s��W�և|����g��c��+y{^��=��;_��������z�j��" 7_	�bbW����r��{ۧ��캓Y7�;�������*�ۑ���v�z�>χ�&���h�TK'�= ��=$h�pW�.&�fQ���#��_�D���q��3Q�ڿQ~��|ǫ��|`ꜙE��e�ʯިR.WG���3J�}x}�};բ����Y��/���\{"=�wF���4o�{�{�~�{��Ao��7#ޔ^7�y9��S}5������ԭ:'_W���|o���o�\a>�W�秧�)��潚ͤ�/R5�_��l�3�3��%E�|�և'�poԝq=��ǻj�xj����&/j�����}<�ɺ���@���Pq2��d�����a�O��Z�QQ��R<�3ܒUŰ��hg��|���/��c��yu!q��#.�wA�g �T2�e
���2-淋����T���f�@^tB��In�5t��/=�5��|O��=�7}�fxz�¥�(K<�j*'"Ӌ���^zsѾ���XJHv�1��{ܚ�b��*z�͸V�	�ޝP��Ȏ ^;�B�Ƙy�a��+��eq7o�>�=��1�d�}/�sڊp�h��b��OK����$����P���ɘAEm�@��:�a�湶�vW
E���^�k팆U�P��c��d���qgf�WE�����n�Ž�m\��/E	���X�9��*Cs��Ƒs��܈!'2*���}p�Bd0���#@�r���J�\�M��ƘX7�g2w�E��0����
]8[��.&U�v·o3�V��Wꚶ�i�2�fnv�
1,!�q�/6ٌ��D�%����n+��DZ���h�0�c4�t�<rn�u�)��ɺ.&�L�M����ř�NՄ\<��g��\w5xm�(K�mÆWY�Iޗ˓�6ә\��Y�-v6����q�Ӌ�f]Yv��S��A£+�^�,�:"��m��C]Y�l|�5Q�f�5;	�X��$Y;2V-e�8�)��u�<�w][��pd�&��n�1̔O��T�n��Y�;u*R��D�E��^�����i׶y]-�1���g���W�;���9|
���+%۳�{(��u��VXdA��[Gx*"2y����OG�m}sEp9A�Y�m*��\Q-+�8��`f�,�:u���j������`V��KM�T/��F���q7[�6Jzh��@��rb�d˚��(�P1\|��F�i��m
���f�P�k[���;�k������A���ipX�s���y�8�	����J}إA�m����x����e��j�7z��q��$u;�d��6L�Z��4u����(Z�l��S#�v��4���S�'<J�+���h��8Z�zM�q<N^�����%����,+ˬ���Q#����,9�̻.��ʷ˶�r1y���véػC�*��e����pŠ钞A�:;���*�mK�����+\��{e�fd�m�H�y�ouV��@V�n\�V��1(�r�T�*�����/��n�̫[,�a�^�D\#�ϓ[��֞�9x�ٹ�����S1M̺O��)gX+�r���^�@ۭ�u��20k�-�W�v�����b�`n�񹽸�����rl�J��C~5x��S���5�̨�T,�Z��J�)i��A,����8���5{z(
��<��]����]�}2ȤM�Nmҁ�;�rB�K9OM�D������g,1a��Dh�Z��N�]���FOX=��޹�ӣ�Y&r	ǚ�F�M��Z�_Rv��=�+zuq �m$��j�Pʑ�0Y�;��;ݨ�e�ne�S�#5Ԅ��[j��cM��VƴN����r;w�b�w���1mE��X�J�,�ykp�9�4�g.�*I$5^�1��츪^+�j�s&Vqɨ���CW���+0. �; u3nލ���/B��z�Q
g�W]�a�ݘ��8t��%�Q9@R�t���[\�D�!2p��0;�꣒����Am4��1*ww8�y.�R��/V�#�E�rU���V��r�wB�,��!�4#��<�NWw\�*7us��)�Ф�\wp�LNRB���A:�$��
��y��w]�=�IʯE�{���wKr,�s�B
wEģ�uetw��X{�m��D�n���-ԭs"q�]e�{��1��+	�<��(��*�*Q�wRt�Z"�j���2���N����jEQUh�.aB{��5w.���\�+����Usgr�	���9n��Aȹ���YN�K�ĕ�jEs���� ����T��Q��"�^m\�=���8n�a'B���w%�J=)�M:{��Y��B@M�VH|�J����x��%�Y�-�ˁ�ܙy�Us����a��ʍwY��6R��8��ӝ��MT�f�T����s,���\3�3��o���y���o�����������uQʙy��gv��TSrtz-�%���xzI���@��ޫ8���O�������w�'��Q+ke���~�`�6̣�I��& "ĕ+ƕ�e�ubn9��8��Q8�O��<[~}Q^���T<zߝǻ"ߌ;�rQ�|ITe�?�"���o��������bFN�c��Wʒ���A�����=�2��0�xN*a?��f�ʾ3 nx���'.��u_�yw{t�BcQ���+����!��y�~�M�{�F�z���2\�Ȁ���_��g����ǗϖlW�<��h��1��h�m��l���x��փo޽��~3�WI�k�9�qn.����I�>58���>�!V��<;~F_��������ǽ>D��N��o�Gy���3^O�$ַ�M!���*��30�c�g�ho�X�q�R����~��Wta;����^��ǜ��e�>J}�Q�Q>�$���`��(���N���[��F"�}Gїr��j�8e���}�e!�u|²Y��3�j:4T$W���mt�ͬ2�$��D*䴳��wޗ�yvV)@2	����S�%?��sS.���t�d��czHB�<˕sc����e-��wט�����lvgP�5��M�ym]з���oޟ z��4X��T��Ĩ�`�J�[�gn$�-�'$�
}��-��c��m��b�W��ޡ�K#}x~ڱq2�e���ڈ�������S��v�唽��H٩ZN��T�����c�h���c��4"�l{j����K�=x_���Y�[D9Ŵү`:l���*t+���q�J7r\
��q�u4�|NǮy�����}�aċ>��6�w�[h�d΋�):v�|2	ಧ�t\t<�6e��K�i���;K���c��󣱝Ϲ)�/��n�=��cU���{�A�2�ē�g\�V�MU�wέ[3l���)�尫�q����]!��7�)vT�qe�x~9�LI)����S��޶����~�ܱa��{A�9��P���c�rnx+%�E�U�O����EڰWv�^ދ��U:�,�S}q7�Kw�+�yο���q�TF�|�w �+�Iȃ�Tbs�3����Z� 6�����xx�sCx���q7>��r �s�q��z�=�#No����������m���f�)n��L�Y��������^�qn*��s��^sJ�r��-Ov&)�y��N:�Z�.���M��/gȅ͗
���K���]�}2���wLL�~�W[,$��He� ��gtWY���!{���{�6�77���=�yoc��?��AF�pG�>�."[�㌿6�W��!�/�ف��l��>"d�U�{��vO�������E9��D*�n�u?I^SAS��9����\���g�b�ؽ�k��U�ޡ�kTQ�%z<j2;uP��e�J���S:^��7O�+�uߖ��U��z�ǒ����?*��|K����@w?]�5�O@!��>ʎ��ǡx�i����M���EɿZ2���ﻮ=�����#�uto羠{��4��b��eH(���|R���Wν�
B<�a�s�]*�7[>������7�yp���8����`��/nX�?�/�s���vwa�z����)�|jK
4��VW�����<r7���m��c��q�O�K��=[/�
�ʡt����Ao�b(_����>;;q3���:�NQ�q�J���F�`Tny�xzF��{{Wey�{ӹ^�}�+��Y�c�>�F/�̩�p�'v��<��X�ɭ2\��>��SLI��yZ��vR�#�߯�箽�Υ�����*xݟ���xA醀�pzbxП�b�c�UVH{�%�M��v�)�}�כ!��>��j ��(v�7sE�U�ʺ���rf��+�c:�Z�6�OzH�A�`+�]��z�>ĥ{����ѷ�����Q�GH���l���_$��\*��aQ#��Άw5GM���+?^�W:��j�,tGC�M�l{+��}Hxj���*F�\�OI�
]���c�p�Υ]м8{h��7Q�:��P=��<�����I�{�o�=�9�^�u�[��EM,��f��G�9�X$�|�j��EL�>j�t�X�i߸�zG��#�va[���b���֮���3h��f�Aʌ�$)^3|e��k���+ޤ&�}�CDϹzU^ǋ�&��+�7�u��a��H���Ps�T�;�rY�P@J�2�}$gL�9�x/�$ΉbH���j�(��=-+c���ߟ����z�鸏W�&��,�"t'���=G��ny�޺��S��9�zp�z��q�Y#E�	��ޔO��Ӂ�q�z���뉧3�`�l���H�I��f�sl}(x�Զ=f����W*�x�6��n�Hd@�x���
��93��*�$��EÎ�Z>�T�5>�p{�3��s���EM�gl����㟶���;�7��^&���z��,u��C��b��k��zG�gnd�Lq鯎Ka�u+N��}~�/J�w�>o�hßWk� 7,)�(�*�J�P���e(�`�j�ۙ�*����L>�I���`O��@�]k�a»;wif�} �N�����U6��Gg|�΅��WY�j�Zk��*Ձ�3����\7B9��r�	dK��l�ؠ��e�s�Y���#-H��2kه�T���{β����||J�0֍������q=�,{��g]S��8��K�l���CT�FF�P^�ޚ���Xws6t2s��wL;��������"D�+�����IWF��iW =��WᎫ�����/�47ODyu!{�R2��wA�e��+=s?~B����p.��[��'�9��Y����M�
JnJ�u�rt���C8ܝ��=Ǒ����,�x5{�{I�~���L,�uH�Et�g:g�o���G��vǲ�����h,����,S�>��ǉh^C�FzrJ���x�d@���|�/��@�}��z|��G��f/q��K�>����z�*�/�
��v|f��=�Q�H<����T�r-eo�����ӿ-q��h�{<���p���U���~w����Ê%GĕFX
D�%.�y���r�#y.���r'=���H������^��+c�CO{e	���(�Qp���Fa�O���p���{כ�y����ze��߼j9~U�}�g��y~�J�z���SP�K��t���t��Jh��Gᫌ�1��i-�g���h�40[��]ӣ�vfLiIqܢ���v.�d�Vs�ƤqUƫ2␃�\���7�8ؽ�2���(vb�M׊���ٷ��Q��)n3sD>�9,��e��*xV�C�r�]������J��Yc�b/�]KI��R�Q����"b%�@�q������h�m�~��Nq���mh6���;hCI�]�r�x߂�k���$�>�R�o��A~�)T�tj�e����j:�������O�>=��;� G��T���i���d���5�B���f�V
�=�B�.7������)|�UvS��&�r�f�U�^vh���{>�"�}fI��Y=C&X�a����u�7��Z���s�]����&�/H�}�w�^�����W��O�=y��z|J��d��;��v&���fM{��߭��Jw�-��Å�m���^Gz��,�^�߶�\,ʑ�,�k���.w�v;�8����>-�;���7�zN��/����c��q8�Q�O:�9�C����˅	��}�ךW�rw�����C�ʭ7�+ģg%����q������;�e]f�x�/8��[XҚ>�~�F��L�NN���2��qS�:.:S��,q�߁�A7�/��"�y��z}tpu���J�w���Y�Օ<hx���@�.*g��s���o�3餤�gd������TM���K���9Aj^��S�l޶�|�vn�� 	�J�nh���K�q��Z���Vڏ.��� �tTFzVM� iV�VŦ�w��� M��Ps��k�3�\t��9:����q�k��ڋ�,�94����O:�
܈_W.X�g�o���q�cq����]!�ό����R��Yd��A�L>����O����Q[���WPv��,B�}�ё��w#}@>�~�=�"nx+�\�iIO۫�V[��w���\z*�*�=qF}��Z���qM��ܷ~Ӌ�<�7��y�Dmêa�_�W~�r�^�կ5d�s�O����o��^F����?+���޴���?H��n�S��>�D��:�v����C���f�� �P��UO�����_���GZ�5K��cW�����������v����W�Ps�U�"�s%�&��D�^SB�V�x��s����؍�ޫ�Tھ��Z����?C}h1�}�g� �q��<j2C�Q5�2��������Q���s���k_h�L���zw����w�w#���wB�y׉�|=>}��`�r|��� �|{�&�u��q�G͈�~z�cg`uQgp��Q�*9���=�WF���u~��>�j�����Q��vu﫶J�^�j���׾�1ޣ� Tf{G������s��v�D>��9�9����t�d�)vI+"o^_oN�)#��֝G��
x�����Sk�v+���j����q��*�-}B˻U��n"�n���]���z��N�Vr��ޞ8�m���]@�4Z�%�]��I%�o���y�[�UЗo5�[�(�P���{�����VL�`�_���Ⲽ6���x�oK��Q����*��I9މ�,�'K�%Bcم�z�~�Yǣ�ٜ7�>;:O��Áɹ8:�W�w5S�V��;�n�W��W�k�cЪ����޺�VC�X���F.72�M����	�,N��pv�	�<��.��_��Ѿ��ߌ�O��_޺��:�$��=js9�!��2����X��M����}�g�Ӓ��L�'@7�j�+�-�Jnu�+��"+և�dD�p��eH�dXK�`l��-�_�Q�$�����v��)��\��wp�z}�{�����Ǽ�=n�;3N��z)Y|�:�ڡ{���r���I�`O�ʡ�-χE����ubZu�+���s�'b���%�_v�Ĭxa~����f�w�6
4���FX����e��w]�W�HMW)wvөθ~�v2--n�}�ǣ�U��uF{�n=T�;�rY���#ž�/�W�����Aȭ����D�y���ﻺ��}�L3��c������z���z�X%�D@n��1�Dw9l�>���^�08z,ӵ��U!�����'9�����:��f��1�E����DL8��)�{فP[ ���C��q���6����.�vErP\�f��P,Y����t�)o{�қ���S�N.1�%���(KZ
!�ݜb� ʻ�%��yI�k��o���yd��^ʞo�F����z�>ȁ��ɿ{ՠ_��_9�L���ٛz��%��fR�!�|T�3�J���6oz�����5pڿQ~��}� ���"����z����\�y&}�ı_A�����%�h�����r����n=�Ux��^&��i������vn�,�=T+�s&�a���Jp=8�JӢ��}~��O������_�#xi�^D��zֵ盫Ԍy��7�z\��{f�����U@Ɇ�mhwS�:."��'�]�>����ҭ�k�`&�\�a��U���:�����[�{���b��TΰK�az�Ni�����z���e{n�
�ׇ�ki�� +q���U��g_�x�^���e����wn���]��{e�j�hz6���G\VUi��e2V}����ݑ*�ܗS�{�� �<����0y���~�Z����O8��%;1Ҧx�VʀƇE�d�jS;��+D����7U��
��,�5�ϳ��NI�E��z��C����"�|�.+���z�<���8�q9��t�OQ������=�ʖ��^]�C�����R���[7O'�a�#l�FR�����Ty@��o�,ף]��ذ�u8�ꆄRe��}4O�QT�q{�w�m]c5�i����zR��Z=[�;n�sJ����l� �Z���zr|�p�4F,�ȧH��6v����n�݆o�#�e�$��� y3�K�-e[��=<��5�G=~Zԉ�`�%և��z���u?;�p5���F��%T`H)/�㢣��}�ZJ��S䮠��<�"���z2���ߣ�CO\G���7�C�%�D@�ǕX>}޶��;9���T|S�&�g��v��u�TJ���!�^W���Ѥ������T��V��i�ϯ�ޮ�_�F��h� �<Gh�a�j+�h�m��l�Nq���mh=h�̥��=]���H_���3Nd��������"~��
�WM����5&��zn�u�TM���V���5{k�TJ>=;�V@�`�"�zk�3��}.{ƅ�V:\o#�>)_���j��a'+w�s}ޑ~�.�����>����:�����&�OF}�}�+�koG��xu��Öt+�J�	Z�k7:���c!�]�{��}����,w�d>'��|�1�f�z�MnVOw��1���Zo�R���_�������#��CƖ��<��b�eH͏���y|"��w�0�����21!i�i4�o�p��P=n�6��`'d��.�-��H�g8C���ͷ�C7��T�f;��ʐ쭩Z���iҲ�dfwG���[���c���V�d,�\�{1+\5�߀Ÿj���b	՘��/�ov��%I,���]u<&:�[Gcw];'+E�iv�ɽ%�\�"e���j�{ż>Hճ�KZ>s/w=Y������k��"���л�7N]��kpk�������)��-�|q���X����e�pc&���� `$YkUc�����V`�j�c�Hk:��[yb"�sr�"��ymӓ��X����d�`�q��<W�spf�2rΩ[�⠺'PS/>BQu{:n��/��޳��{hZ�-��f��B�+x��^�8 �ҧ>�b�#̨�+׌��{l�Ѱ*����$@��y� ���R���Vci+3�[D��;E�bh]�Jl���&�t6vj����}��p�p�*[����n�>�*�В��΀�S��Yg.��D4��),�[��N�M�7co̦{hu4�M-h���4���3zs_\�'�;��ۈf�1�#�A�]0=j��,��%�L���f�5�������� �Cڟm�=�^��,)P��z�s����ZM�#���g&t�.���;�2��]OX�ʂ�2���HC>��`�Oo1����iT�@�R\n�lK��vS̳�8'y;)TӝR��Ɋ�pΪ汝\~ZCѿq���\�M�J&
����}WH��,cB�8�f�������l���v�V���Hw:�fR'9�sz�T�{Ã��&���yv6A��K�-f���Q]y�έW��A.�����S��u&�y�:�j������U8%�܅��m�Gm��%u������սvs�ÊG9�f���:��-�Rl;TF��0�왲�i�9�
U�	�'qռ�ՙJv�c�H�rI���%�Bu7P,�yp�c���$hť�H�v�g(��j�B���Ks+��΍;�F�!�Cn�Wd0�9�!%�����YX�LGo|�r��@b�Qcs����m�/2U�;�>Nً�=R�r�du�SV��*��=�T�j�t�0��s�ke��t'֞��*��x�'E|�+P���BB�w�k�Gm�]ӝ�@,���א�ڙ�J⡘Y�7Wω�@���o,٭j�9��ӱ��!i���1�I\�]_."��^�]��C����5��%5wꝒъ��1+��z�1�<��2��a�1�}Y`���5�@ո������	�!��}I�N�U���M�U��=��'͔���|����)�K��.kW��oMz�γYs�c�\�-���j-]�h!Y�x>�G"�yԯ����q��h��LQ���u��7���wvt�]p��%��DLm��;oN�n5�]wJ�r�����P�$[�]u[��fF�l��;���7��Q�Kj4D$��&EÞ�p��*���xGIȝIu(�t�u�;�t���2C�
��k�45�q,\�u=\(�n���(�z'ww̹D肞���E.��u�#�9�#��(ᣞ�\�$;��T��n����AVl)W]T+�<�)hY��D��gN�zz��9���a竞nr��sP,�Vzyu�rY�Naf3і�{�%�'pU/']�W/E�2s�9�+��5)P�ܴ�2�<�jy'��ut�N%����I�W7\��wt�:������ii�͊*.D�N㸫u$��:y$:���qKU$0�H��2�wid�D&ȔM
Śx�G�Ћ�*&\�ʧ	=���R�yf�����S���B
zJIPE��VID��V�3%K+�TR��,�VQZ��5��hT��rԒ�K
�s��D�HIe�(IdF��Q��9��%ZHR-r[�Do>1�gR;���Ka�sJ�Fh� ��w��������N"�fV?�r�v�f�՗Ӆ'NrT���Ł+��kB���I_�'����;�u�Ѹ�S�'NF�~7�j���I��js�������Kz/�ǜ\)�����=��r԰t헄x�y�\o�^%;.}��=��ix���!�uT!Eǐ���_sJG��y;���;�t]��ߗ��ۙc+�3�\T���4�yN��N�!�~
݃k����-�#�r=u��v�;�޽f/VT��R�,e@3ŋ���/w٢[n|-th1W��k|�H�w��X�F�^\g����C�{�g���d�0��Qز�=Fa��Ph���zxlv.�޴3�c�3��+�PU�Yb��X�O���7���c�TM�p.J3�_zh�#�[�`߹�	=�3
�{�:�ϙYj�������ND/H��HJ��s�:�8/Ȳv�,Z�~}�ޖ�X@O ���X�|e����V9�~Ws�ZG"�<Webߴ����;7s|�Xb��{����f�̂�(!Q>�s��~,n��7�R
�)�����ї{��3}Zc�{���O?z�����E9��B���Q%yMNW�۬�una�߹�ʉA/��
W�:e�f��0l�ϕX/��j��%쟽��`�G�[��ym�����*ﻅ�Uԇ:k/H:wP�i{��b5�5�)�bQ�����E���-�]�s=�5��ߠޣd���`��������kU.�H��N�d��d�U���}���+�»��g>��}���%�L\Nbx'\	�^��`�%3�C���.v����f�t}Nyt�9���T�=�qμO���g���`�R|���ten2k�?����-1qe~ɦ@���^�h�����utn��u~��>�j±���Q�	v�2=s��-C��)D�������?��Q���M���U�5\��z�}��Z���X��@n�]�W7�/�y�Xc�3{�K9,(ӡ�φuK�t�����vڸ�;���N�WA7��K:�ԌzqK����=q����fp�������~�:�S�t]J���˼dL�V���$�ql%�!uO��v=u̧须��z�m�Ν�Y;�ü�X݇�U�W;�q����gsק�.��di�F/[�߯��޺��:�7O{�H^���Y�)G�9�`֙��v��8R��(�˨���;΀�Ȏ5B���"��n{c�^s�C�T�pŀ?f��������˝���D�H�E�$�_I~5UG��3�n�\�Ʒw���W�O�܍�u��$�Q�E�s|Z��z�Ѫ�JPW���
��"WC`܇����J�t��[|�=�5*L�-Kʎ4u�l-v��V�<'Mt�3�;Ո��@�9����H&�/4�w��O��-�^���(����!��k�{W�S�\�IN<p��5��M]�-�jx/@6K�S�Iꉖ��w�L�>j�-�	؆���;�Ʃ�3���o���ˤx��W��_@6
5��|e�!J��-�25�w�Km�q)�w@�ZT�n{��W_	��}�z�=냷�a���|��� ����V���)
�Ԉg����?��k�z�}�CB��y�}�lv��w��A��G��_3%���Ǥ����FJ�ܵ�Y��&=�m�떋��:�w�d��~v�z�>���ɿ{ՠ\{=q9t'�e�F�I���b�ϒ>ݙ�#�䉟uz����VDr�~7�f�o�����ޤ����|���DO���7i�O����U�f���xW�f_��8*"_V������Y�J_~ʏ{ʪ�N멣J��E�{���:�h�9z��doZE�x��.�~X=mv�}�}[)�&�:�`�w`:��^���Fy�v�gϽ�7�� ��e���3����a�����T�N�W~Z��{�Z�������q-)A{��G�/W�FDk��{���UǺ�X��eN���ݸ3�+}�0�D�̿^ѹ�:=���!ʙYB�7f�f�b�]�RC%�&�3�+�s,��9�v��V���&ky��z�ڷr�q�ۈ��x��;f�)�Hp��G@���[z��o+�lk<��R�X+�,��_Q�_7�sU����ƺ��?�91��7�sʼ:�_3:�KůM����s*F{�#칕�-܎�R�A��!za�VUi���x�����vE��ܜwQ��t�S��W>�q���jYI��zrO]�%����=P��(�WK��s���x������y�.��fJ�K�C�}�H�M�<�7}�v1z�$��$�L��3��>S�s�\���~�w�O&s��]>�nr�5#}��3���8�>�^�Q�Qo�fQ�H;�X�>E���KǔM��V���Ͻb�6�H��;�B}����1����[��a��b�P��*��2��-�@w�+�ۥR�H��M�wP]�M�	-��dB�י[�z�����ӨqD�b}���w�	�Qp��.�2�f ��9�L����3Q�޿+���yb��~�O�=�#y����,��׸�\�;�'��%MC ��"e��o��}��r7Ѩ��M��z[%�i��3:rEO�=���z�{Հ{�M��$����l��"b_�
�t������#Q��@�5v��k�b]�k�j(F`,��ߜ��'�t2/0�H�Z /<U�D^Vw�^�ʿ��x���wà᣹��� lζ���b�2B���;kq��m@����ڣJ�}-��e����s(��5ͽ�Ƨ���l�}�s��l�ޤ��C-����#��s���Ϗ�<O�̲̀BE��30�p:�T���c���:L{�Z��}!Fʵ���>iT�p������*=���@u���%��2�צ�_����+��f���OM�lx�7^C����5Ds���~����:��z|���.#�� �O�Y��o���t���-���R0�S��qJ}��~J�8\v�߆B�W��}�4�}x��B��8���@;�j}����5zE�O��pwj=u��nK�t�j���J�:����Q�M0�=5U�c£6�I�g%���{ی;7&����/�}:�Uq����Q\��Ǡ�ª��Dԁj���[Ӿ�:O��x����%�w��i̙�k�t��2�P���Q�%��˭�W�O*��v/+V=�o�Go�N_��z��=��\w{ՌYS������� �:=^�	ڽ�5�'f�+{�X���>��Q���Fz=,b~�x���]!��3|b�eJ7Y'�N:���^l�Dt���m������s'uTR�����p�3���_��Ǹ�M�U�p�v�o�������9&:.�6�1ѭ��t���5��;�_L�B�.��?"�2��V��b^9ʽ^�.��DdHٺ�� ����Pd�#2a��֌v�6��$ҹ�R&�ԦsX�C�^a�(J͹��{A�5A���.׵mc㧴��u���wW~~�a�P1����F[+>�w��뉹n���y�do���
e�m;�]�M�t�嫅x��R�%�) yI�u�x�Z��#�S򸛉��#W����p3g�o/�����9��H���YG����25
ETO�����_��9�m��G�Q���>��3}�j�o�?D���a�u�t�wI����n=U�"��f�T�q�FD��4�n�b���t�����p������\���W��yY�6�kƣ TC�Q5˓�&a{���QՏ�Zp�}�y����������q:�^��;��{�:�>���������ȴ��o�������N��g���25/*�w�V�g�#���~���y�Ѹ{����_��䢧�+����or7��o5!z���*A��K%W���;8�w����w�R��v�\,O�h�w�7�:c�c���K;�`]BwPv��^L��,jK
�·9>���<r7�����N(���T�Q�<�IV�~��ʦ��g��)x��T_~�{���ٜ6����χ�:������1�Q����O@F�!��˛`S�aP�"v��ҮϚ���Mr��J�fC��4�e˖&�n�+ȫ���Ƚ��- Z��F�JۭKR���Xz��e@���cW`��E�<�z��O5��T�&H�}�lN����)��*
]Xv,��]�W�})��&4'�>���l1�T���:�/���vG��1�s:vd���a�\xo�1�W"�Gu�n��=�xz�i�TYi�X�������׼{!�!�r=�/VT�wy�i����@7�ǽ�G��^�0��A�T;��T��w��L�V�=����|<�W���B���wg,���eH눹�'�}'� �� ��+��,�uP�z}��{����^���Rs��#��j��mϾwԇg�u�X6J���z�X<���s�j�qMՉr9ĸ�t��v�/C٭,�,��V���;�#�;�<u}�W��_|��( yQ��R�f㌶X�͙�������R~J5 s�Ͼ��bo�����h�zF���޸;q�aع,��	Q�.����/{9Ѕ��v#��îgǮH�ޙ���x�X�\4z'�v�g[�?Wq7�\7���L�g`�L��&s&ȼ���@���Q12�*7r�}�G;ֲF����>�"}�NO�����������~���3�.���o��DϺ�F�\�z�+��}�j9�^���H;��W�fl]��� ��D�6|.��͕��]�v�7�C��j˷D���#C�*�A�wl��q�*'h��G<n�w0e��S��	k���qG�"*���[ŽC$W�w�r5�j�4;,>��Q���+f.wv�[�'�`T��sR[�� o���>�(�tw�e���N
��բ����Yĥ�����?6�X�̛�8�S��꣼Z&���P�s#c��d�zt��=8�JӢ�+__��h��\�rѨ>��9U�G�Gu��^�W{�G�g��<�YGc���7�y�U��ya��\po�ݯp�����OdwS�����呑�Az^�ޫ\{�E���S�C'2��3�h�E��+}��2yj�z*�%#
ⲗ�J��V���~gլʇ�^/��q�.�=��*��{��8߹%z�#x�s=aᯋUⲫM���+D�bnȸU)�8�WO��o�����F��o���`����.5NI��(m�L�4g��~�F�\3�GL����8Ĉ
n'W�FU�{��yG]Bez+�㻿m�w����"L%��	A릗�UuU΁r�����vzB���M���@��>>ӑ����q�ό�G��7nH=FX �0��"���}��q�F9�y�m���-e7�W�X�~������}A���q��3~0��F��%Gzm�f�r�����:d�b��JR�~�	��.�-�:��M̤�(�X�')��)
*3`�Х�L�;�:���X��]��j#ۂ#;�d�㳪>���^U��ܦ
�r��G�R9�U��K0��D�	y��:6�[��|��&��su7�4��{#�n״
�%ꛏ+�>�o8H���z2�����P���Bt�s�#Q�{�~�}9�][�J��F�ޣ1�W����ex���9��q7�,C �+�����|�g�Ƽ3�;�0y^�w�p����L�4����"e��n8�Gۡ�r7��O���ĕwB�J]ټ���6����{Հw��f�s$�D�Ξ�&"_�
�t�����\4ۥvy�U��W=��Kk�����'��<O�:�)�2E"�H&��Ղ�%�x���v�EE�o���x�P&�69b��o��T��w�R=�*�1���h߽>����"�}fI��d��}�6+�p�O%g�aN�~�+��ީl�K��wS|��1������M���y�
�xR<\fMX[�=�^�j�����9��1��0��K��xhܬ�B�W��ޡ�K#}x��/�8N�993������C̩q��ڀp&n�C���#f��:u��m_���i4�g��>Z��5v�j�P�f9���Pv�ݹ�Y�7���ӡ��>��*��L����d|��>���sC��m�j���/7o�u޵�.{Rz��Xd8-�sc���T����/t�Xw�pA�#:Ѵ���V`��fjx�:�e�꺜xDz8�[3YQd���ܼ[|��4U9��S�u�b8
����M<�6Z��6��O~�r#�b�������?V��5��w�<�ϟ��Y�z�Ɯɝ��͉�2	��Q���SUG�K6�n��rwѹ��}
g���w�n���s�]{Ǳڸ��z���Օ<n"ωJ����	��sY#+qi�w��FǪe3t�_M������S��^�Y�=���]�(�F��U�lz�/{�=D��3�D�B�����u�RYb3�^���'���@z�������(�^��w�VJε�B��'��UA�p&�C��,u�s�>7�7�r��NB�9�E����Y��|1j�����Q:��6J� )�����x�-����#�O��Sm(d:~p�\Z�h����q�^���3޲6�4�ә� "�}DL�\����v��C�؜��\�>T}�Hq����:�;ӺM�z��Ǫ�dW�d�P�a��DO]>fiE�z�ǎ#�4<�i#��{|�Ft&����>��<m�׍F@t�'>FXꏽ�k�M���mПo.*J�[�
Y���;T�wEy��^�sC���9�d�X�(�}��G�}������co������M��1����l�[m�cm�v�`���v�`���[m�cm�v�`����m�cm�ݶ�1����l���l�}�m�km�m�m�cm��m�cm�v�`���6�`���v�`��������v�`���m�m��1AY&SY�+�� ��Y�`P��3'� bH��Ǫ�(�RTPUUU%()U(�""R%BI*����UJADEEA@$����R�����H���UJU��"�(	UzV���R�(��R
�$JTR)T��R�U)]���*�P*J���D��H*!ASX=�	"U$����TTJ��Rm�A�*RD�"PDU$�U)$�!骐(�"��*U"*RUDP�T�)J-4�EQ'x  ���ML�p ��FHT)b�´�MU���m@�L0SAe`�CH0(	��٪��	U@J���!N�  �4��Ef5 QV�ƨ�n�9�4  �Ѣ�M�  Q@÷th�F� 9��:4QE\9�Q@@h�Վ�(��(��t*W���%Sf�
%O^   ��(�E�m�UV�al�kkA�hl-h��@cV��Q�,j� ���+ Z�!��%{$@	�  ;�(U�`�Q�V(=
��Y�QT*�h:u`��*f����%��� ).�h �4����-ݥ�T�DIE)*�<   1ª�(�� t��T��7en�1� ��.���*��Jj �M c��S�j��:����ԥR����ڥl��(�EM�  u���mZV�+��C�E1��@4	łT4ZF�sh�Z����R��A��kP(�k
3l@�ػ��ҩAt�P�!		EU"+�  k���j�v�R�4;q��m��Y��u�Ӯ[n�u��i��imVU���(қ0��ƀh�V*�i�i�g%�N�C��$Km�T �R�k$x   ���f�P��ݶ�R�C��iV�Khɍ ���v�b�Ѡ��)��@:�mt��+l�,�êkZfP4m��a*�����JI	lj�   ��i@P��i��4�n�b�SZh����
#:��# �t�ڳZ(ݎ�b�m�l��`Ҭi�����҂�H
 ����QC�  -v�����+MR��e2�
��mY����E�@d:ږ�@Q�F���@��hV��[4���a�`o ��&eRR�@ �{FR�  ��Ȇ�z� )� ���@ �� T�L��i*z4ʨJ��)�W"�Z�TFRX2�S4W
:*�~��L��k��u�o��k�$�	'5��B�	! �����	!I��IO�H@�2�HH[���������m�yy��A�T�h�.i���yz�ڼn���)n�P|,C{�T�L���j<Z�d�J�5Y@!�JU�f�Զ#��5�Ӕ�\�d� ��ҧK\Q K��J�d�t��jV���G4)N����UM3n郹�dʀ�NQ���n�z��QՂ\�lxi��3�Y�k�B�n�	�f�ܥ��%��'Nە��*�J�炮����Qh-�ԛ)
��К��`��6��/n"tP�LO�w��ҍ;w������h#^�٤���B���7^�ҭ/XM��D]h��w��u� �GExD٩�G촣.��ŗ{W�1���E۽���j��e�ZA�T���:�ae2d�ޓF*�w��ْ�mf�P	����K2�o�;�3Pci���b=R�̱X+ Fˉݚ�M�jˎ�J��J��/f�u1��}9���T�҉�l`cHY۬v���Ȯ�#��Y�$����h`%-5i�r�n�{�*)���9t!���2�S��D$+]G{�;ɭ�:I"�p7#��)0��n7lJ,8s�û��B)2��am�amH񷺦hl�`��F�{%�a鬆C��_ �y���2�Exe��������7�̧��UtK5�TYLz�YEVD��c.��U�t��XV��L�*�[�v�*P�Dݗ��)ڻ��;y �2��/C@hp3b��w��2�o@$�N'��"��yx���ڰҥh+3!�h�1�W��j����b�i\�5-]*���k\b���EG�+:���̢�����;@<������˄p��X�i�m�:�2�2����Z�*2�R��c��5U�9�v��c����P���դL(�GU��dm�[���2VؗL�,�6T�5X�4���l�V�C4�����
�oj[�J)p3M�Z�e˽�([U ���e��@ʸZ��Y�"��g1�j�9���@�kQwYj����vB�$Ұ�T��E�����{��"ME����!��P��]C[��@^,�6���e�hazͪw�e;���wI�x�[TS"��2��+��ll�cU��A@86������6��u��إ�[%�j�`4�h��2��n���.V\HIW$�8�p̼R�陘�٬�-8Q��ղQ���� �\���]ؓ�J�_��E,�Q̠ʥ	ٺ����T�4� ����C��[P��Uq���¥��fRZ��4��n�)jv�ie^�Wz�W�{t� -E��j���I��KF�j����n��̱D��Mᙱ����XýB���n�R+LIQ{�m�H�i��d q�̨Hj��l͸,�������2�1�p�b���Bp�n��`��V�JJR�c"�m�sU�&=&̙2K�M؛[�E��$6�
Zӥh]��E��T���bJe�՛-^Ӹ��;5���)�@n����M[��VZh#)�HJ����&���ٶ�_XL&MG�mnə�(ܣٔS�F�JU��km��A�w[I�iݍx)�2��WyN����[E�i o\�k[ �k�/���;��[7#e�FT�L9Q�VUK�u�w5j�RS��--��2���e�ʋU���7k��.wbQ�1�uZDZ��0���5x���i�kb	��r��޺E �� ���Z�`��72�^���q�̼q�e~�rQZ�,ҙk.��?*t�ڠ�V��]���5	X�-:`��I��ۍ��Rۅ��m�#Q�$dn��v&�m��L����+q�-���D����cIC�&2U��-�G��Pmfꛆ�2�9��p�:�d�.P�o5��L���׺.����%8YRUʄ^�:��(U5�Gw0̐N[�voֱV@h�!�OjXTa� `lr]�U��L�EZJk�v�ۉҬg30If'�f�K;�X�(ųrf�[�K�uݴ��#Y�E�E�F�*bl)f���MZ��d,TkZْ����\�iu�1n���n�ߡp��h�%��i`N��S�	��ݠ,�%N�!=��ī%�{�6��D�F����i��,T�
�Zʏ][ֈK�7Q�X����\�m�7A�4j�j��U����m����ٻR�w�Bn���r��̡��x�[����B-���~�V%I�=5+q-յ�=�l0([���˹tE��#b�B���$"��{��[�L�X�6�R��U�a)�����Z�m�����n�n��Uz��yܽ��G0Y���VsQ^5-Vkw,�FP�b��A��Wz�Ʃ�Ʀ(Ru`l8���
��U��2��b��r�V���A͇5�lhz����3h����3�{����Q���/�N��l�=_�0*�ӭ�
���\�T�z��JʸK^�K���u�y*�vh�b��QKB�Q��j�`2�Qȡ�V&��K\y� ����^:lPݚ^)wx���33!�)=L�k6]�m��{V��7�� �����^ِ���ùB�ݲ&r(�`w�����X"�7��V���S.T��Q����W����z��wP��n�>�VC�އ&X6��u�R�Mf]���(oU�(i�w!Q���v��tZ�b�M�Zr��O�m5���rc4���0W�D��TL��`L�2�В��WF��(&���R"��B��d���q�W-����w��y�d;�؉H�����@�l	T�y��2�V��fKNj�kOh&$�Z�l��kd٬1
эKͶ��h�,��Aoƞk���fL{��j��:dmk�D�f�֛���H܊�ۍl��7�p&;�+[�bL҂a��i�{%^ẚ���q�a�//�q���A���4S3YƂ�xu����B�k���`� x%z�%n�K��9�9q�@	x��j�:ak4��rw��bKc�$ 6�X%,5��cѹ���(���[&�B��V�ӛ��J#�e�ڈ6��Ғ򎺹�mH�Ҽ�1��ي���%� 4�@ڭ���Ә$�P�qh�u�k�^��l@Q�[@�F�إ-0E��,���l�6A�G�)�PjE��:1�i�eLϢ���A���l�ɴv����6J؝*B,ՈGI�dկfZ����I���b�*P^5z����V/JbbӔ�Kj�@�8��M��@�@ZJ�]nҴ����ѡb�T�B�S�ǆŌ:ڢ�7��F��a3�҃>�Z�b��+F�:�w�� C�-�ww�|NV��]wYVS���[��Ѣ"��V��*��fē՘~8kZ��0Dee�f�n�����U3v���Ą9$�,�XW�jf%OU��L<mދw�(곓��*V"X*]�yl��̫PTӪ�Tuᑛ�ʛI0p�M��(R�"x(Q��-c�
$e=�J;hc�m�4���%d7>2zL�����j����+�2���F��ͣR:�f�#)���F�j��m�t��M���J�X��e�K7M8�ٵƘF�͵��M�ql�ߕ���fR,�v�������FA[�4w%8M�#&��H�(��0CH+&�X�H��P�\٨x�
�wEd�l"�Є�2���:��'N�U�6��x3i�c�ig#��<���Z�)XveH+stG`�k���"�#N=̢�qݣ�6���v�%�YDC�E{��^JY��U���:��x�ɼ�.�P�Z�'�:� �ڗG�|ŌNַ`˩zU�ywm��j�[�WW*��#YN�^��.g֨�V���ӥ��X�;NGC�E
͛�9w&��,m=JP�hY��g"z�L`��%Hb����MQvRwp�xfQu��H�X���(�0v��7'�U�"�X�j�mJ�+�m�
U�������R;�a�e���r���#��KPMϖ�,�e�`�V�<�J�2E�fY��C-��LUN���ͽ��U��B�ثH�=i���`�7S�䷫B����n��b +�)��n��,U5�V�TN��`-[y���S��lf8�[c���(��>F�Q��S�Afh��rݦ�M�4�f^�2ӛ�[�*�ſ&��6����GInZ�;�dY�u��U����MkyN�H5X�а�芼IdP���[	�C���7��D�;�����K.�;���"�HmE����ad�_:���HM��֝h*�M�+���zե��4�چ]�IpaY{a� �&�^�p�޴͝�Z����NfP?	�䖆�Ɩf����VځV�L�D���F�(�Y��,i��^��y6k/ujQ�ˉT�iEʳ�NT��4TTo#�J���U�ڋ\4������ʻ�:�M��h��@�z��E�ot6FS2=Q3�u�@c7i��)�m=�u�{tTsuZ��*f4J���Y�6�4�a��е���\�f�H�e�/Q0­�la��Nm�z�)��M^��Яͫ����}���Z�s2��1���jת�x�9drZrXc��s�,�6�y/�N��[6�P����Peѵ����9��ٌ�q���kb��u��-�d��,a�˼��7,KL*�$L֋�1�Y�[q��ج�4�Z�n+�Ӈ]
�	ң�1
�BV'%�E:�6n�kwq
ơjX%a��ħ�(Nb���F�a��ݵ�dHP�/P���q^�+jk;�X�*��pa�w"�>��4�9�
7u���Y��j�`H_^ݝ ᓳ3.�D�!����9sBDG���Ir��7b۲p��J�^�ו��V]��b[m��vȮ��3�oX�EM!g]b�F��%eǱL4]+�C~&˔���+5�Or�9�fև�X�ƪ8C�®�kZѠ,c&� Ji2P�����(��~��;�0�DU������]�B`�0
7E�j-ϒ�K5��U���2�����u�(����D��4��X��JYp�ث՛��)�4�zZ.P�C�hˉ=�6���-mӒ�N��߉�Z�7x�YلlX�cTň��7Jˤ���S��<��.��YA�Q���Y� FB�X��0�.��h�6���mH�!U0Fo0��xh�
�.��40?�1���X�.`I-�}�j��T�+l ��H����ܫƚ��9E���.���n�A�6�'n�d�:kL�@^���]��ec��IP7R�^��հT��+� ���2���Ń.�L�x�E�-�)�$2 �^�����>d�7oVa��-m��Y�J��;��vA�cUj�e&�6�q��c��Uma�*T�<إ,�,���Ee�]��Kխ���)咴ZP�M�[�	f��l���č=iIM�*�����X��ϯEH�?�+�5V^0���<kt��řS+T�[�����.�:��n�VGQ9*cCs-:ll����p��Je�{�AhL��x���mX�K��^���\�X�g1D��Q��Ch���L�{&�,o��-%wL���j��m\�!FS�����@�@��Z^��J��%yl�v����ܩ�⛖7U���2�\C�aT�nՙ��ƎR��oɗiGgw�Ȯ�eh(��#�Z�.2��U��f��7*Z��1�řY�Ƭ�i�x�
�aq�zA��
h��[(���$u��Ab�=�*�Le��Y�s䖻�u�8ӻl飲�<n��VeG��N��ԺSn�U�f�sK@5�	�X��Z�Q�eL��)�!m���Wf����+��	ws�SW�Sٸ��ف��2V�h�f�X�>�&J��nm&5���^����Y'Z�0�N��+vC�⮺nLܦ*��$Z���+Gv��3�$u �ihY�j���V[�L�cr���+�ui�JRq�(,�dz+lR��{z�q)m�KE���Tsh,�Lz�b����4�n�u���H�va!U="����1�e�Y��ȣs$T��8˼tp�vZA���@M�fixU*;0�
��0�С���)e��V7(�:����`<�wbZ�뷘.��qЀ��;��Q�G�R���-mKcZ��m-���"p96
�	�TҪ�,��m�Y��C[C�۳�n�<<1R遪��^I�!�M���n�C(f+�6s[[{��M��	��z�Y�m��0�)�wke�J���zՄ7JD�X%E5���� z����1��IK�,ޟ��W��e �R�F/���+�-��F�,oV��"�OuT��1WZ�3�в�ocku-���.�9u�B�r�'�\3~����3T[fj��m�d0�l�%@U����Iށ��gpǬ���a��*b#�tX�H�){�����I��ԭ hˬ���7(RVi���\��r���(�W]k��#��׋X)Cv���n���!0;��T�e�V���
�(͍�	�dW��˱�W2]����5�<'2�	˥1S��ӗ�O1����G+S�1YEܢ�Ib�/A�M���Z`G��x$��&^��V�0�rP9[%\�N+�l�{b4�51Bjr��S>���f���>Z3.��VK��
��>�l�Z�j���i舝�-�KL�.De""�`d�!༫b�����ً4bӚ��|�j9s�¤�ҭիf
Э�n��R݌^ӥKZPk���Vt+(���42_K�(�� ��+1�.�,:�r0���n�(M,KG)�B4��K{u y�����mj��7/0!��*��ĭ���>Bk��Q:L�����q����Z��m]^b�f^`@������G�u#Xٝ;7��u�"5���;��.v�j&��ؗN<�.���qV�S�y+��Z���#�ˋ#Yz��if3��K5��k��hv5N͙N�;��\/�ID�׽ǶS�g{�6�閲�0�#�ɱ�K��;�x�{�gA�j/����Q�q50D�z(��W+(��Yǖ̮�0��ή���l���ŗD� ���)K�O"�:#J��x�����+o!��?t��gV�A��v+�r�zT�X�u��!4ȳ�t�EY�{%wò���U��2����\��%�q\ow��7P��X�*�����×-��\Yi��q�)���A)f��0�5�RSץn�\�԰ft�����󊇵�VJ��d�;���xR�o����'ع0�o-ۖ�b�+�����s��+�0��O4<�*%B&-oM�p��`�`b]�zv��#��M����9]0�vS_i�w*�2�.
��D�Op������d2��i�'�FI��aP�웬��i�!*X���Jٱa����m
�n�_^޶��hΓ�]����]q��gm�&���G���p�8��s����,���^��@оKE�����2�������axf:
����{�:�K	-�\������)k��\pԦ�F�7�����l}������L
��%��凱 
��qQ��u�q��9y��������+�� �wp�\5�<��Ǔ��1k��|Y���ns��Y��^�����:u)V��WYt)w"�(떣��g2��f��{��2�I_=q�rV���W�����]<��r�C�"��[͑�6������x$���ԕ/���t���ޭ�dD���s��Na��T�)�[j�YE:p�Pua��.��_/.���_.����Hvp$��'�[2�m��\��▫qԝ�uR�囔"�������sڂfKk�V�v��c}}���BygpF<�^n�AN�.��e���_2�+TUM��Zյ��ӅL�96N�ձ��*�}�DICyQwn-�3J��wz��|�7�����E���wz9մ�a�VB�颰_q��~p.u:�xwkW:��	&�����x�9�/1����`� Z�6L麫�v쬁r��F���l��Z�5���7��u&r�;Ԇ���� �y=[���o���ʓ�f�j��nW0�wa�lkՀ�9X٧wo�<H�G�#��왧Ijڝ�w5Q�ª�r���I���rBh���b�n2pzˣF_r��*�3ۜ�W��n+� 'l�G�P��;/+���'t7Y��i����W��Ι)���e�I�$��䷷�����v��G���o$ev˾����ù���c�qkxnc��s�����ohvZ`n�x-�^��H�"�]���q�2]��I@z\
�K��{��3/�������|���{|����9X�4Ȳx0][Y�Rd��J.�5��۷��WR�B��W,���
$��`�Q�ل*�J��ER�7zvC$;9V%�M� y�tE�]�+����Vk	5-.���4��j��U�VY�ػm���H��M7^qwjͼ��;[O!�����!���V�Y���rY���Z�[@��#�C����սco��X�8�[�M��YIh����(���,�:0��w� �v_�&B�^�`�V�7��s=0����Z�V�D(��JG7�M6K�0HNj�&ҡ�n��l��)�7�5�s��[$�Yw��=�@��:�KmI�����ܝ�<}bZ��t��B�W:�ԥu$�%��k�*Zǋu)�2#o|અ����F�·_S9),�c1�'c��ˢ�N�$sr��_��[���6ys� �m�����u3�ە��i�X�lP�2�q��-��|�;0`�׮����;	��Y�u��mb�SmK��;6�ok��=)\Ut�4[��&F�������L�]/�E��
�a�φ�ظ����GEu�nE�R�
tu�-��ݦ��;Q�v�y�7�\��v�|�vҼ�[�H����,n��K ��d{;��ܓ��T�κ�Pc���&ͥ>`�%F
��;q%��#�u�=ا&b=��	�e<�E��fA���R����n.�ׄxWUr�R��R�v.CTZ��i�^�j��I���Jꚙ&�� :�y�]�waT��ɨ��Z����$޽n�T���Z�N���X����h��Q3f����*�غG{d��?t�hjZ[��P�u�pٙ��ή磢�\�kl'ovPLu��r��á�:1��=C�2��*��T�%�o���N�e�r�M�8���\��v���ZO���y%hn����ejS�P��A�ك2 K�����}3�a.	|�	��J4��� �v�s<p�2��,r���� ��*C;+)	������J�q���C�����C�l�f�J�]�^�|�'X�z��z�u�7�����rI9��ut=:��4���v���1+�77��#�tӖ�>����(���%4h�&�]�a����v�����γ�v=�\���#�+�kb$��=u�nl�c7ot�����A�Գ/dQ�8�L9��N��#���,�Xl�]˦�;�lL��D�]N#k5�tݻy�-�9Q+�	��nV,�c�3�<�gt*�͋�[N<�MF���Q�ꕺn��X�Ҿ������(}�Xܫ�������ºd��Ի�Y��斶���V�e�W�l��-FZ�4^�Okr���K�(��ҳXG8WK�I���+_e-T�;��->�:&�0;D���勚@�Ӽuя��I�˭���O��B%nƆ�ۃ�[�u�7�C��k��Kμ@2�Ku��l�+癿9�.��n�P,#7��p:��9k��>ndt4B��]�ڠ�+�|�]�fU澕�Xo��������,���ᣇ.��y�9�MƶQN�=u�>�yˊ�ms��oa��t��p[�d�&J���ܺ�\�u1��U'��r%w%��{��v$�)����!��{|9N���J�LMwGDK�Z�	֝b
;�o���Fd��N�p��l�FX�9HY�"��3�|��7.��J��΀���)�7��n�H2���A���u����A��Q���P�]�A$�;T;���*8���3��oZ�c���L��r,V��t\�2����_�آ,��\����HV��1������9�f�$���	s�	%���Z�0��4	�*Z ��U�{r�T��O;��o68��o8!׷��w��ᠱ�S:MG���$����car�Cg,L�>'���sy���N�|�q�~�\�)vR��$Ь����aR��ܧ�=�y�;K�ݑYc�d�i�ܸ��M��yk�:ka���u��q�1up9VJ@fr�i���N�J��,X�:Ю���^o*|q�m[��GE �����A�߄��x@rn��W�f��K�2Z	Id�9Z��gԳ��miH3:Mq�1���A�1���6ԝO���YLTOj]uu���Z��j,Iݳ	u�S��L�,�^�5��"��X Ȼ��u�"c{�o����S�����d���t��,R�o�۲_<;��a{���u�����m��ۥ�rի����먎c��h(���rU�٢�&��h�{-���^��z�<^���`�cC��ܭ��m+=T�Kя3M�A��T�u�e��\�:(<<��nm���ؔ=�P����
�@���{}�\աص�g'n_Sњ���A#[M�/Dh��docIr����`r���2���e#��M"&�yaԭ�,'��m^�Cvw�q�ݬ��?j���N� �c2m\��.a칽��s���$��D�aH���Qm��!����̶z�+]�)V�)K�e�\���Y�G� �Y�3�נ����*:T�U�����uv}���"]K\�MUǟv���hGK�&A�����z���<��b�]:���E%�8b�b��c��5G��ѭ�|�_R;�k9���.��Ur�w��,AΝ.ס�}�늭�����A���s�*$*GIt�.}YL-��s��S��H)��u�9����ϱ�gk3Z�c�7`���`+�Y%1�f!����84S��=86���z@`]��7n���y<b�bE�,S7iP6x��zظ�f�;.	Xێ����j�Nn�u�Clv�E*�vQ�P�6��6������nZi��XL�
&��q���M�M'�������$h������k�k\C��βBV]woMQQ��H����Vws�zl�c`���VY�8W]cj����/��ۦ���v#���NѢ�M��ZW�W��(�p�)⬱(��yʷw>�c�	���3�F�mʑm��[ɣ�v�3��4�{3m+LX�7.��Ӿ��ι��c��j��u"§b�={��V�2j���]�b��;G�8�C=׻p�RL;/m��C�R��T���[���w8pt�[�eenLhnj�ٮ�$�mk8Tj����m��fМ�8���df���2��=n�:�f𫑪�����Aӭ ��7��Ӫ�I۽Kw;�4�Ϳ5�~�+�)4�1X֬�K&�}����)���V ��(:T�љn���b��,�����ou�=�"�J���a��F����YwO�2oXRv7Ou��<	S.�싺z���"+&���.��h�n�9�z�p�*f�=x)��`R��L�����TE��LB]�K�	e��*㬲��)��~��W�Өj���2�TGy�y�hY�*_lCV���+j��6�V�eO�I�ͦ����c<6pԭ��D���L�y�`�કfr��jк�����H����J���*@��\.\x�V�<yds�H�V��x+��z�op���Y�`�n֑���3�5�9e)�6劗b��Sw��b֮dꕢ
�|‭7�����K�Ӷ�WXޔ37�	n�șU!�m�Yӄ�kn�Nq�y�u�����x���Ѓ��z�(��]j�DI��յ����+5��
�M��Ir��w �-�Mj۱M��\����Mt��DTF�P:��,����.7��gc�r���9sK�;�����YL�f�a��+K2S�k�n�gc��c��$ae�����uGmj��j�����|�Op�[a�D���x�]�jk�<vGJVL!��=��#�
���W왔�QƟ
;G�|jU՗�V�n�p��ڑ�M�u��W��1]>���'ur�4dI�$�X��W�9o	%�/�X��΂t�+����1��D���Zھ��|-D�uJ��	��(Y�>Iy}˺��3x��v��9�j�c�)m�����6���8 VC����� 5\-R��vtyN^��"���\'d�z��;.�'���O�9	{-;�����N��8�"��uա
+���
�Y}�߀�[o��e��unʼ�v�w��.�d|�����A�:�Ep,��a$�4v�|Ҭ�ђ�́q������+���Aru��C�u���Kvg�K��ow�3�ϲ�H�Ыwt9A,	���vι�������eHې�a�#������q�ns�P9��ɛ\ c3r�珲�3S��dI@!>W�ϻ#���M	W�5��m�5+rhRfj9�]�%չ:ھ5z��KN�z��2YќGz$�&N�Po<�$���@y��2u?��9���}�����ط^BT�����VeZl�,9�'T�.�L�w�ً���{���	��6U�p���}wۡ�>U/h)Ne�a���e�8D�2�����b��9i�asP��"y�U6��=ȧ�j�걵x��U�}ﻅ��}���,�Qe�WD>7z�N�+�啒^�̾��ʖy�읳t���q�F������dV��×F/'m�^8rI�F�n§I1D��sn �[�j�*W3{�U=��:<<��yώ��1*}����an����ө�{��K�(��*}� �|��Ò�|���`KA �+���`O7�N"����P��z��F������J�ݤƎk���kwqUгK;�h�m[�X�%��Ԝ����80J��7��k�K�t�P�Βn���H�5ط���3����W��3yi��l�d�:MW�@[��k$��0�/H!�����
�7m7����wl�7�?7Z(��z����뫣���,B��}t8>�y:lޒ����R_N��NX��,ޒ�Wiz>�X��aX���E� nn�P�Ӱm��ln\��\�ڽ�����g�`�_;]"x�toQ!Ι\ٸ�7�R��;��a�6��[�NN�z�,V�[R�-e+dKl�;�Y�Ft��E"F]栃��_W\�.���	b�Nr���Q�(��
�#�����\yRl}i�_mu���5��9�3\n���㷪m�1�s�2��%������n������ԏwų�Sw�7���̱�K���>�	���*Я��=���wS�G�����;��W�M#�[�y;;�_^|��)�J��,����@*�d�2�8��)X�Z��������X]��a��
2���C�A�'-� ��{���:����qҼ��#e>�j8\�f��Uh�}ӌ���se���þ��'m{�VmL:0.��u�f��o3����ϻ�·�q�)�vӹ^��B�r���nٗ+���ق�A9�SpwP��.��S֘��=*��{On<�h�������@e���s��G�=�i.�]H�����޾���܄ �	!I�y��4��"i��Y_�E��)�u�5�&� ���v���w��w^�ւ!Ca�]ٹ��S�����kT��,�7.�]DO���C�f�MQx�*�;Y���� ��ms�)7�V!
��g�������p��
ޭZ���K�#T�=����w]��J��KD�)��`̷2 s��u(�3��܀�����b�9�8�wkN����^�m�}�e���۫ɝЧ}R9y���/����"�q Մ��hQv��{��c)jĈ�;�`p��0e��֝B.����o�n�j�7+�vmL%	��QI��1S8�S�d��W�P��v��+Yw��Mֹ+͝�1`?f�nDh����R��Y��Y[����c�I$lf���j���_R�/㉥2]�!i�^v֛I�9I�F���<�%v�}t}ʹ�?J�Ņ�mE�{y��&�KN�A�ߴt߱�Jn��f����^,Ը��%
�_Qs��'�������5�E��'%OE �45mp�.����|���Cw`�}�^�����X߱�/pgԀNǇ�7���>��MX.,�|�3LV����Dv�M*M��ܸu���wf���L�񘯆��4�vw�.��3��d����n\R�wr��w{-R���Z]����mC�Թׂ��3��;KJ�ϴ&��M�h,��RoQ5���]q*�M1jP����ʑB�;�n��*�8	Ӷ�+��h,ڲ����o�X�s������ař8��n�#��[]��cn��xR�yq8 =�e�̌S2�ʚ�v�F-����4^�J�C��v5��+���J,��[�.)J(^\ꌬ2��YrUe���R�˹��st��Q:R�B^�T�Л��#�6��szT���JO;R9�:����b�r�:���x���b��o_)�i�lI\7P�n\��)�x����1����;	7�b���w^f���r�i@q�pȸ�T�����:��\/uj6l�|���	�CZ� �Ȏ3���=�mv]j;P_���=S+M,� r���ڛ��V%l�5��2=��v+���W
�z9�p�a�������M�PR��uЮOs7e��}@��+�M�g�dܸ@�R�y��z�3ZL̼d�{t�+��b��Jw��"2A���\��O�]otZ�N�!W��p��G�oT� ��'PXE��(�R���@�|���<��.�(j]�Kg�n����%;�F}�erv�N� "��VN�ݞ�V�j@��]m6q`a�1r�vI��ƳWS��3�tT��g��u&E��)�a�/Ji���eŌVQ�ws�EӨ1}��޾9ZF�5G��"�^Ά�ü(N/8eE�^����3s)L8�Jge\���圢�^��-SnG�s�lb��������x�W�'q"D�&��jm-��V�K��IF�R�pP�X*��z��ݦC���VH��cs�����ۮ�r����Ug�oh���+��䩝[q4%�u����}��.sN�_:!&U����]�2��y���֞L:�˚���p\���Ơ�K0%��*��D}z�|3����J�ր��r��WkvXx^K�0u.���7E�P���Ǘ��VeJv��6�@�{ơ��#x%C��Wªb��3N*��N�=����G���]3 R��Z(cxw���J�>�b�+��/p��R�$�TkM��C7oxɹvz�)J���$\���l]��W�� 9͌�����e��F���CՃ�>�X������\�w]Λ��g��I�Y�:a��sv��Lpi$����G׆���򅕒���㓰v��P�2��P4�:K�y��af�נ��W�ғ<E9O�[�����UǥU�2��]q|����9�V�	cE}��=�(,i��iQ�����Z��U��(�f�q��̳B�D�e-	�E�$s��ku����P�=��e�^�f�>�3V����X�|�.Y��f:o;� /a-�U;�弹�:qczDĮ���{�sF u�VWs�w5�Ԇ�)�7��Wc�|��ۂ�+��]�vYtpbsu�gq�Hw3��2_nWWB�6�'Ւ��Y��H��	�),�}�X&ڬPF��(��=��ʖ����',�9+3P��hjǁ���_T��w���Q�j�7k/-�����YP��u(�P]�ǃr/��G7�P/�غ��M	n㺾�>U^���&2�ih[w毝���aEʶ�pD_!�9N�1�m�6�MԚ��u�־��N����M��q_<<'v�x�1r^(�b�'�uz\/�)\E�U��4�W�u]�q�΢��!.J��υd<�{b�N|��*��ݍ�+�&=*5��Tނ�we8s9�l�H��ƻ���gs�K�6sW) n��M�/�������/�c�`��b��v���VK.r�4s̰w*Vʘ3^�/���DU�}�U�j��,[�a�C�uf,�bW�mZ'���sU9�2������k���D]+�,n}:�|�T�}Hҩ����Z�+7��V��Dݑ��#��^jF�M��]�t��͜iZ�V��Yb��9N�>�`���1��'G(e,3z��S�ۓ�ۭ�b��=`>XRP�,.���%1�@˲HM��\�s������w)7��[|��tU)�&o|"J�^���ѝ�#@��^Y����y>�4�Xs/l��8�m�y��
�W���6�J�8�X�0G�5Tu�m���:���,�v�^���ʹS��ʝO��.��<�%�g(_^�����m1�ut�P��Gp�5X%<�Gi)
X�)�1痸�������"�����L�M��r�0��i�G�J�v�r�9&�YK2�>�ۃ�R!��f�qx��b� t����Y8�1�w�m���@s���

��5h]y�~Y��,��E�uݨ��20Ois� ��p,Z�gV��AT�_#�sV�O�7ϒ<]7Qt��ɯ7�P��AT�s��h�I^�Uy���7��IFv�L��^uJH�k�Y٘�J���6T:�i�\N��w�R�$qnp����;������]ʳ2T�&��R�������vS�|�_9@��al�+D�wy]]�Ⅲ4�������h�����=W΅��G��v��.�B���*�Y��5�تV����[p�;5���Ѵq��,���y��ÇY��JGU�A-Ҡ�AIcT�,�f�AI�	���2J-`��;h	OC�Pm����s]�]�N��2ns �Zu��u�{��F���p����P�Zp2���B�*L���Qc�+��buoSx �G�����빎m(��7Υ_tꛔ�ؽWZEj��gR�S ��5�1�uu6��Q�vq�����|�u�B�� �vN;�ӄ����:��=�� ���,�m*E�K�졻�edpZ�
F�.����	N��S�����s��B��cn��wT�`D����Ӻm�ݣ�j2�w����\)a���evsfJ��V�+HOU.�d�Vr��[�mf�m��[���XXL��ݜ�� �[W�e�0WS��o�������w�j��+!���W}����u�{C}Š��n�x�M�b���������5D�8\����>G~�y��;+*%�7��ul d[��5w��U7)��T˼��1{����/h�w-ߐ�p�V_+KD�5�]Gm�,)^:�ԧQ][�`��t���Ku��5s�Wк�R�hpb��u}k ��#7�@]��Pˆ�+t*|;�ؕ�j��g��R��飘EQ'����w��Y��)���
<d.�fఓ�X��e@�v8殒�#wO].�e!z6��x�����\�0�՛�S�0���ތ.�\�bD��f9�VC�o�aiS��N�͂Q�����:��<Üz<Ҿ��6�R�j�h愘r���	�@��.�d!ŽV���4t�J��;vV͑�Q�l{�t����n��P��`�&�d^��{��]YxäNP�5:6/��ǭREL��W��ܫ�Hf�t��tj��j�kxP�맍-��t��~w���(�It/[�;NW]u)+i^-�Gd�[N]�}��Z��x+�;,Z����@/��͟17e��k|%oe1���v�C�ݎz�i��0U��v�~�2P֭ب z�0�2۲,c��s�5mᒘy�z��	gT�Lb�+�"���׶�wN���[��Ý��.�.��WZ6'�Ӈ��T�WR1�u�Tw�NU)�iKj�7�.���]�H�u�2GԤ�Cz`?M�ok�lu>��%<�DkIl�������ԧ�v���n�%�VӜpYk�%0{�Ehw�2��^�jM��lv�k��K�5���%=�*�1&��#M�+;'A�6�{��wFZ�B�݋�-����x&X:�B���s�5RqP���C��攇�0���K2�bsH�`؋g�&�ټ+�0�5��u�����5Y�$A:��>����B4�|nv�e�b��A���(5ֻ6j�lК�k��sy�����6�ੱxwz�QcO(d��z*�[y5���F�EP�&>gr�S�t� ވ�/z:9�B�E����G2�R���vE$�e��Y+�J�i�xh=��d<�DV^e���1:� �Ux�v)ϖ��p�X�^�d������+
�T�7�U����!p.b�f�έ8�) �ݽ� 
U��ٱk]]�M��q�V���e8��[�%�0&��_P�Q��*��1����1�%u�%+\�����K�K��ޞI�4,/l�C3��zLU���&��N����j��Q�J�\�u���9����T�gWm���c�;���D���x�S���G�.S��pƢ��N��"[��W �k5un��Uj`���b�,�����w	ɭ�:��A�.&T����S��R�ww�ӈ\m"o�i��Dv�r72����R�f�f�Y,u�������3ba��2�	��H�C�YG���ַ1�ړ�=���Vދ��nf#c�uќCp<w�S�L�ش咎u5l�r�XY�"�N��V�p�N<����&P�+�T��Yj�Y`b�4y�xs�Ke��z�{�
��f�ǻ�o���-�� ��[�P�`cnܫp �Õ�b����x��,��Y�\��`"�Iع/r���6U޳m6T��5f�rN�ċ�8���U��)М���y�{�iԝ���[��1��HҀVڬ��Ef�����>����ʳ�qU�ՙV�>س�I�YP�k���,�E'6/��z�=&�I[��5�Y��2���y\>���O�=D�N]s<FD�.C�7o,��U�YY�~�YMJ��sWCU�i�����;ɼе���]�ԭ8Ժ[wF`�D^f�/��8S@�*C�긨����B�Z��a��KW���P2kWC4��mR�w��r��L�|���2p�4-E�s�Υ�}HG8t
��S�j׼E33\"��\澜�WR����U��m�����hh��C���3�vd�4�,�#�����Io�eۅ�i��g�N-:u����t�%�2^Aa�T�!ȱN�Y��E��ޏ�]�B�I�.0lk�Sb�n�WD���=)�eʵ����;�s.H#�o`h]f_q���6��hB�ͻ4F�EƦ(��89��z�{|o]�"f����I͖$<���hH�A�s�*�hɩa��(P�1�s5�dHQ��8NA9Y�r�I�k��iQO���N�d�R�$ n�Ŏ[g�֪Z��wz5��8F��[�E+�����հ]Z:��Զ��#��e���]N��������������C���f���ۧA�S/}`��i���|܆ ��� ���/:Ue�,Cl��ga[WV��E�]�g$���* of��1W4�z���������y*oѦ�W�Պ���yo�$�eܝAgV.�g��9xl8���!�f�wLJ�p:ffr��i��"�n�}��ƀ�vn�3J6�,돬\q;l�D�E֚6B:E[��'o9CW@g_|�	�f�a��qp�r��_��J˗�s�7������ݾX`��ƨn����cٟXC6�εo�a�ڈkE�:�H�ǆ��2u�q���*a����<N�ǫg!i�|ԧY� ���Z�L�.[³�3.T�������Ӱv#L�HY*��5��)�^p�ċn�g_1��ڷD�+�˚C��$���7l��Q��]���k�rp�����Lܫ�WK�m��J8�뺬��Mە�v:�rt;S[G�-�.�!Ǫ�v�u������k�.��k�;���1��d�b����	�pM��]��7CT��v91pU���x��|�g �j���ox�u`�j�Ĭ�v:�Ir�$�ª4	�K�3�D��7z�]��@�@�H�-��2�No]�h���͸A�ft�.3�ݎE�[۫��mmҵ�\�1:u`������|�pۉ���u��Nr�8�����`���nay�]5�Rւ���w��c2�ڔzJt���M�-�  �Wod�k�^��N����ab����q���;1�vf����K.�v�mCW�GsV�>7�t̭ʶ�e��P*���b�N�S\lc�5T�eg6�^�Xs�b����dq��p6�q*��ԫwt.�ɳ��Z����/$�J!�dΗ��>�Hr���_iݚ�kڧ��u�2�;!S`=�n�oM��(]�y�{b� �r3��WV�X�]�j�8�\L��`&��Y}���B+޳Q�3fr�k2+ō�CJ43o�I�	
�:qf�l����k��R���l�"k62m�����7���G�F�����_W�O6Ȍ�����pkj��k|/VV�墢ȫ(�����C;{�M�Pq�oLcS��T{���:�)8�}����)٬�GeoYC���xﳵ�}ڬf�0��iJ�.8�$�(Q�ar�T�#@�BSG&�q����x��7�'m��BZ��cU2L�;��D�;�K�{J���ٮ�< �y���Ը˧���Vq�+s:�]�Q@�23ո�U���wk�>A���@��p�:=�����)����7�*�,4�D&ܚx��y���
͆���[-
���;N�:�f�"(T\s3p��Aܕ�z�*�A�W�K�/8�sl?wH�v�B8i�Qѭ�<���(�2�l�[^��Ҕ��V;<��,s������㫧���]r7��ӭ}GN�/�����mP��u'2gἠ@�;�㮇�h��Z*����1K�k���e�G���3��5<�)�żD�m�mr{Y��^)��
��*2��F-�:�h��^O��o(���u631]�m��w�f�X�Kլ�o �<��]s�L��Gp;���.���t��w���:T5e�n�t�>u�s�����=��K���7E
��ݒ��}-��H�8�H�e�z���G�<7Y��I�jMW����X��G\�+�ݶR��4���+s{�|~��괮�I�����.S��՜�y۽�k�����O��?�����0�DH�*�**�F�r��V(�8Z��UƩ����ZV)3.
2ZR(,�Ɍ����ą���f2ň
cm%Q�G1�,S2��U�TƌTEb��e�ȫ1�Qk*
�
*����Ȫ,�Xٍb�fPX1E&�IX�`�*�kZ3D��,Um�V0���\l�QL�X�dm���1��e!��e�"+U���T�"�r�b�b,V�b�T�Q�kEZ%Dr�b[TZ#s�h�eW1s
T�KJ[e�VQ�U`��dm%`�YRTX�a�#(��4�DaZ+�"Ŗ�amQH�[m85%�TX*ʕ"�JV��\dƋ9E*E��R����$Q@�&����o�_usP�)�묩�jhg�Z�ek���{��)�q:��B����ʙ@�܁J�wO�igv��
�����M�s�sݙf��?Ɔo)f���B|�0�*ױ�5��I�__g�(c��e����vp:&j�9NI�B�+�w����P���CY\��U��9��d���w�l�˸]�K� Ͼ�I�g�����(^EV�8����%Q�l{D���!�[\�����U��af()H��]������E�鑙�0R���j�i�a�OR�&�"��z�o8��9u�r!m���:zx�#t5��W�&s�>��^d�E��<CzPԸk�®;!ѻ�;!kyl���u�^{�-��)����<%�W�/3!�;�ؠ)m�uk}T��%������z�Ҷ�S� W�p�+�޼���ǆ�|�+��ǥ\|2c�˽�՞��e�F�[-����$�#��qA�9��>c��!��|`�[���9�ہ�I�b-$Z�O�b��>:dK�\d���;�����ul�C�Wc��e���^��R1	����i�uW��]B��.���k6�1:���K3z��k1zx�yL_8��8B37#<+��{�j���lw:�T�'Gs[�Ԫ�(��c�;��䵂��������2��X���G�rһ�"�T��%�fV1`�]P�YLh�gq��HOFl�u�p�����&*ⳋ�K']�����.�b�ݥd�`�jG+��������[�~�%pt�6;�e�V��,��a����ˡ�0m�zi᝼�m�	!��wl�VV�i4A�"�U\f]Qu��XYȦ��Iw��s;"��ߏ�?u�P��f��"�n�j�ԋ
���(&e��췪�M���g[3}��٥�r�E�o��tս��?\kؼ�ڄ�%Rǒ���S/�q��Ռ��1߻x;��d�Kl�Ӂ<�;��Y�Y�.�䞷��C��~��'*��n���Q1~�����I��
�gS�zK���ƿ)��̩kǄP�#.����%�����{�4{X}KwI��HƔ+)8����_��Ƚ��MgIb�9Y~+��H|��;�Ϋ]�=�<������uF�T8V��G�y��<.�}���Y���db�),�b��=jtB�s}B7E�R>:˸^%�r$Y�͜��}{E&U��r �=H�˫:SA܎�)��,'(0\Y��1ҏ+ܻ��X��]�+Ge��R����֏�/�X0��5>�楝�YCT4�z�U���y���s����^���v��OP8�����!6s�{��5�sF��O{���$i��ئ+����{��a�۔�X-T�꭬��m���CZ�C�$��pR������ͥ��۸�o�Α��4_+��;/y��,z�|���u�G�u2�}0��I�oJ�u��vu��KD��{�n!��%�;y��~���:��cF3�����<�W/0_{����f�,��L�w؆ᗣ�t4�{�Y��YxWE�Pտe�E�`�;t�N�������{��S����R_���w^8z��>����Sj�Ԭd(_
�gQj,�S!Ř��lr�>��o�Ly��&�j��C�=���Y�7�J�KM5�UWR����T$��3{��r���{�˗���'p��V���\���4=ɛh4�Չy)
��qg����G)��FWW.�kص�,��� i{.匓�+�����S�	��_ʈ�_%�uZz���
?(����o�+���j�.j�S����&����V^Gxq�(;R�;��^�뽷s8��uٙ�@� D �0v)�9�_Zg>��j�S��RƑns���OK~Ys9I/П�˹�Fq��o(�g݆���R$�_XPq_�ƃ���uD�6>R��8M*��_� �|��_� �t}d+\�V+:�cQ�2
�e�x�DsS�z�8r��QZ�-�:k�6�{/���ͭ~��81��!=��ЭI�B���Wu %�5�OE٫��[��J�7�N֡�����k"Ȅ�l*�]oX�^!�_n�˛�<�Ps�h�p=}T^C�XP�))4�du/��lX��+�9��OxSyi�G��G�J��w���x��/X��`�lL��D�ī=�� �S;�[��g��9&�Jv�|�;�5�zU%�C�.�9�H�6B���t��I��h�ʞh�A����s�����vl�۴�+N�[��rU���j�f4L�2N�#�*į-��}�f"w�rz��
�mj>���T�����X�m�k�nV�N.*�\���#�bz����i�^+r]S殽�l��-Zچ�&g�7¡L��U{]����:[G���kK��x>���;���E�3���Zpx;�p�%�sS:�Eͻ���\D7S'��U�g�IK��x�M��L��#�{��VڣXUVl�Ғ��O'0��y9�Ǘ/n{÷n�;���c�e�v�19V��oW�.�臨`�VZ�8R�ꑶ|��G{�k1[��\�;Zd�_T�p����S����n�= �z1��j Fz����WnT��AVm��	�&S���uo`��5�k1�0�ed{t�	l^V͐�[�}D�h=��zo�ze..ҾDݾaK"�K�,��-[�p�˓~82��<�u�QP�j����ͼB��]�-�<U���n7iwpJ��8�%c�|ٱ�$��%\�0����:���������6��;0`;<�*WX�7�o�	_\�u�A��F/.%z�Z��'��n�vv���b��hs�O�.���x���<w��e-����=�Ht���;��]D/��'�x!ү��C+Ӣ���Uv�����8ʿ>�7�\�՟\�K�vB�x�]:�]S�Z/s:wyt���s��J�|]G�E]�%h�.m��PvM/o�.ؿY�~
tcʼxř��}����w��,9��TŸ;E����wpWu_�S��mh}�R��A�N�&PO}J?��~��7�4�:�-�z僗]Ӽ�^5�c2C�����v4L����W�1�ou�ӍOeDռ��kڻ9�|�z��.vg��^P�v;=�{������F��k� дN��2���Qk�g�ݡ��T{{��������?j��@�R�N��7kHلi�k�3��M��D�͔{�A\�Y2WZ��	��W%�`��×l���H^�p��P�,��`c�n����sIn0��z�U৸ؾ�:�s��OS����>1���M���7��~�ګ�~�6�7�u�~�~�i��=�F�������{Y]�>�F����-��.{!�C:�]Sw}�ڤū�s��o���P^v�v�����;}2z�¼{�5c�^�7�����k�Q���D��[=��s�3��]�I=��<|뺠~Ǻ��j�����az���1���1!��O|��m3��o����_�?^�\�xN>��;�Ŋ;����u�l���-9XW�9T{��6��@�us��'<϶�%����x�@�N��T�x{+�e����C�2�/��m[��ϞN�q�L2��B�e�sgQ�<��N��t�W�N���Ǫ���/3p.�����/�_V��6v�E�Ir>�վ�r�ld�"L8h/Ga���N�6�t�fU�Y��V�uX�)vr�`n����e��k`K'u��^Y��^nb->��xw")��Mg\�{��(c����X�X�Է��l�]EmmZ|���}�fU�8ch%��Y��:�ޡJ�є���X����R��)f�͐�Y?)�g���|��]y}��/s��L�65�4�I�n���3�zږ�����-xv�۫�:���1��h�=�]Gd��a=��}{~���oňb���p+�K:�'�3���?uN�Ÿ���|���q��2�N����[���\$�羽w��>�{�{��瞜��Ա�q�ў�^n���a�7�������Y�3��Ͷ0k�a��cӂ?m���]	O�:�O8��	^gݰ,��[�*z�nE�37���������>�J{ ���hl���U���^���[k]��Q��/��`�r�r�i�B`�n�y�|;��O�s�����L����h\ͯ3�ϩeF/������%��W������o'Ҷ�|y��I5�鞛�+9�S������b���d��V�M�<���;�14G:`.?w��}��
����]Oj�����f��b=I�!vj���9�Ś�M �l�s��6�E�;(M�F;�P��<�/%��3Q�aX{�G��/>xx����Oj�x*V驻Q���ݚ�p��]�ciZ�yn>*�7l!;�{�.�%���ym���r
�m�6<Ğ�A*��q�f=3�	gZ;L[�;��s�3|��ݓ����u�WX\߃�3�
~ޭy;/ qܒ�x�}���zQz}������XC�}}N�t�����s\�tjǚ~�=�-�N&{���%�x%|��>��/���g�s�[���ς���}��7<���"��r�����d��.�O��:�w�8&)�{'�V;�<��'�ޟwF�)q�U��h�^���ח03��{<�]��
\��f(Ͷ��<�2����h�<��b��a����;������Sڂ�v���n�e9B�=��ot��z"�����7���~B7�k}.h�[���^�����ͱ��Կ]=����S��6@��s�5�税Y�fiHdN��U�[��$:��}�?]l��=<�>N[�[�}R��P�`G�6g�x(Xu;�H�;G����ܼPcI��7R�0�En�N�"�m��כA�m(ݵA�hJP�ZY����^��>�wo�N��\+�aM�B���8$�Y�K|�J{K�F�I��'A�]_�)�ٶ�`!ud�W�2崝�;�Vz�?^�<�����ҷ�Õ�o�*�HN~��h�K�~j��W�=ڙ�{W��|}ލUqM���J�*۴9]�����<����C�+ݴ�i�=f��zӗ3��`q��	�7���i�ܻ������^m:�n���������cq�Ӌ��M�C�bz�S�O_q�����Ǚ�|s���-wPu|/�7�$�A+�f���g�m�KQ�٫/��7����Gk��l�j.�6l{�y�~��Q�J�ߵƽ��z��K �s$zYֈ����`!ί���75��Vz��Ym�>q��s˩�\�t_������I_X�kFu]�s���s�o��&t�%� ����Lڒ��他;!k<F%�:-����Ν�3��'�d�^J;�"��%��slLW�+��4l���~v�J��K�V�+4h	�e��!n����^tO���2��7�kd�y�ժ�4N������X��^��Ok76�U��)�:&E���ܷխ��\,�lСo�ĳ-^8-(\�sd�ܔx��	\3�ܶ��N�	�':��Y���k.�{yK̏>�:�����m��e7+՚yw�qmCw��X=���8����s�c��f{�6�Vk2��~}x lOϚ=6	�+�q���~}�f���fg�.��Y�A�:z�sw�zU�]+k����z�-^�l�½~Ծ;ڎ�Q���?a���|�=;6�f��A�q�3��{O_��A�n�n�*�b�x��^�g:����oo��d��9{�y�ld~�W��XU�S?+�A��O�@��-��˼j�_���/�,'/�#�Ms�Or�W�Y�k�y�n���
��CL�?|��h�{��l��y�i΄a�zi�'�2�-3u�z6��+:Z���w��;Ke�Lu��6���ϥyp����*�}�</��=&�>�s�-��;G����%�E�}ښ�,_a��-PY���T��lB��+6�cȥ���I5i����k4�e ��kM�Y�����luLYq��sv��&YO�-Px�]Ku�*�3s+%"D�8����u�wS�l��wYڍ)ە0jw,�����'e�J���kk���b[ȟhF���u��z��1:��T'�a����$�BO1ݢ��(���s5�k�(�.�`ڬV�'���z���ƣQ�u�p���y��ҭ��|:��x�Cy��ts��k6�f��s����`pݳY�V�v��]p 
�5��&e���-Q���#\�"�O��'P{��>φ�nh��$�=��żB�0
�GoEM&<��)�!��!k{��`���G6��(�q�j�QS�h������{���*�%��wr�#ɡ�J.���跴�ewl(F�+�S��x#�M�%]��r#m�Wl�dj���&�5��qf�U���u����U$R��2� }���Ǣ�6̥��̭�qX�Q��	ͷ<��G��}�ݴm�d�Z��.�U׭�;;R�3�t�j�J�֡22h�����L'5�d��NS�$�+�+5�>ĳ�4��R�Pd\b)�#\��"�i���]t�Z�Ġ��c鶪܃��skM,�(@S"XPê=�*���hk���;cQ��.���Q��^�g/���wa}F�gk����|��;�����r����=k8��VN�o	HJս�pNk�q΢�,�r-6⫢�/aB��D�]])�DJ�{4�X��-М"{��ő.t���h��F�x�kY��{7���f�.�X�i&޲�J��(֩-����޵҉}��L;�Z	�iF��p<:�k]�W��ΰ�.E:{���Ԭ�OK(7fm��f�ڏ��=v�(�-뜪-v��W�r�V�֋��WS���'��]@�D�W;?s2'��\E��m�[�
7��
�ʘ?$�j�%���R��
Eg �xZ6�s���H)����Xe��Ӫu-�5${Wٕ䆤�4	z";Pf�T���C;���3NT��p�.�J�z�!��g������w��o����RF�d������P�Ǝ9e8�嗋��r�N���jU��;�<<s8�Հ�*ۮIX�g�
��NA)��6�)�jN�é���-�k���JnO���N�eK��?]�Ó�-��jp'��G9���kR� �h>e9g�4ԼgVw-�!caZ���d׵���C0ElZc�����v.�|..���ɨ6�{[�+m����@*���H91����;��g��r��� ��솞�����m�d^Kf��.�o�ҥt�چ��1�=�L������ux,
ؠ��Ε�;oG%�G8���Sy#� Wcs���Ӥ�&Kj��PU����r�͵�a��$�͠ˊ�r�g�׻��s^��\�?�IH��	c��T�CQ`�+eATX�0�X����S��PL�T�
�DV6�+*�̪#mEUQa����Z��*

�B����Ĺe��*e)�UKh,����Qd�Z�@\�Ec
���1�k1Lj�j�S-�Q����H�(���P*J-��C��V�R������T*�̣KR���%�Zʂ�Y�Vآ�0Q�9V孥����cm�F��QƊl�� �*+dPQKLs-1�e���#�-��*Fҵ�Q�+"�̮$YFUT�,W2�AAE�kb���c����1m�i�q!�0U�ԕE[TR�5fa�� ��faKq�Qb �\��+J�-��ʸ���f\+Q�dXb8։e����331i����bP�32�\��8�Qk�b�h��Qkp��4���TcJ"���Q���c%����p���*u�1�s�([���5� ^�l�8q�k���qh��:��;y���C:>��L�;�������Tc���b;����9��>�u��ņ>:�r����JO��x��������������5�;/w,�J"�'R��^F+/��=���w�_W�7y����75U��|f�WAn�x��%~ҽ+���� �a=;� ��'����y�W��~���͔�2��͜q����_m����(k<h':�S����=^|��1�VQ���	����WAO`lV����םt ��6�,\~x�t�>vYW���s}�>���Q�9�V�Ÿ��|�<����/��Ok�rs�v���ק��پ��0oDi�
�����ӓ��nzm�i��s:JkJ���lc���r���6��{,>�c�\��q�yA`�]�֗�����7�z�M�2��ԝ��\Y7�������:�*v+345�C"U�l�z�x),�:{�,�'�q�yֈ7	�̕7U��"�e�v�m���'n�I�#��a�L7�n�U��=ok�]��J�f��F�������K��E�,��f�
BΎ#j�R�[}�+
Zz��Ψ������{�S�����SZJ�жY~>�|)��;d��Ǝq.�G'��#�zs�+z���H����ޔͧ��5��B�6z���f�y��|���co��4��I��L��Vr�M;z�;;���u�3t�u��>g͡��63�C�M9�8�xN>�۵gG��oE��x�gl�6�:'�>�R��Y�?`aۚ���g�Lۖu�U��W�gי�[ì@������w�����s�O�Տ'e�f�ī۩뎚�iɇ�6�_o(r��@_S�y��(�y��Pl��3|C���{:�Os��S��yxu���Cx�K��qu��M�j��]��>�d+wq�-��K�ȥ�$�՟\�r�tN��B�Ԟ����(��	Eyw���\�tg�j�WN�����8+E�6��#�u����|<�8�K�ϖ"[;kX�q��ߋh�����^Z;�xSJ��H�s}[('�fg�p59�y���mt���x3���ڷ��ٰ��ƪ�����J�uV�]����fml*�%ι�mwɔ�w�g��9dQ�>���U�5��wr+%9\E�������g��T��]߶#C��DƸ;�ÃΓ^t�^�N�����\紫9����~��c��loDh�*�.B���J���o_y4�z��w�ʹ�t�/��G�6湧�@��KI���٫������+xe�����n�O:�����a��[ݙ�<ˇ}�K{����A'�sf�L{�{{=���]���\y��+/���*vT�:�þ���>v���ӗ�3ds��<�����gҕʮ�[$��畾�&�@�gl���,'.`�;�9�s6ng��nw
�O��޼b�4�E���פּ+C��pl�7,:�0�i�B�t��ś�ɶ�X�|��!�y��`ŰР�l��bOg��.M�����~bz]���Ly$/K;A��>,P;K�3.Yc7^�w�:|iU�魥��U�<AiޘI�qս��d>�z2��%`��m��h��}�ޛ�򣝘XUU�Z]n�L_r"��Wu�d���ԑ��Vi[:w*��$��q��(.��6����_+Lu�N��!�\Wcz�7w�Q��Ծ���c9�!�A��,M>~<ǹ�Τ��=�,�:#x���5�}O��6o���uk=Z���U��>���Os˩��n�����	��w3�NFs�)bb{Ϸ�>w��i���z���I��K��r]�a�ȶ�/�*Cʱ@߇tUgL	�U���R��[�ʏ�U�Ϝ��T��?Y�B����^�W���>�n�A�J�&k�S��͏YtǷ�������8m�vZ�뛎�gs+�ls�A�Q�?������}O��?e'6�����a�N2���i<d�f��>gY<C�gY&%a��>���l~������#�?���P�'PX9̂�=J�S��'���Ld�a����$���E��X��&�S�2q�ה4�&�q"o�k�;�ڞw�&~���~�#O�q����T:o�u�T��'�,���8�l�y�p��l��׿��d�VJ�s�	��N��,:�x���?o��Ͼ�g���~�~�����L'C���i��>I�2�L�A|�0�hu>è,&����'�>�<I�M����r��d�޳i'P4����M�q9�y���u�%.��lן�^o��Y��!��̆gO(i'�O�_a�i��P<=�I�:���z�OP��2u4�6�y�Y8�	���:���=��M�o�ޏ0�����V�C��>x�r|�ݳ���Л38W
�1����@�����J`Ef^���U�e
w]�Rf�j���*e^\��Uצ�o
o��iى�z�4�_Z���h=��0jn��\V^�z�k�7����N��1V0�Vr���>�����n}���c'�NRm�?2|�2�m�d�k,�$�+?j�Ru	���2q��>�6�:����N���N��'��}ì�v�k�{߆��ϻ�����~��=d��;�2N2O]~�+&�����?$�52��?2u+8�|§���I��d�&���T�I�T׼��I�����=�߶s`%�gxH�����}����veu���w�|�0����'���|�qњ�+��C�VN���d=O̜J��m���Aa>O���8�Ԭ�k����߯u��{��~߼���E'�4ʝ9̐Y6Ü�_�N��s2u��>d��9$��&����'ɬ�IRm!��=ed��hu����I�8�֯����;�޺��5�kϏ��}�''�s�Y>J��{�8����}���5�|�'?$�l�$�'f�d'�&��d+$�~�쒤�C���+'Xx}�^���߼��7�w��|~��hq��vad�$�~Շ�$멟`q������2q����}�I?�m���O̞s���<I�Ý�N&�5�2���ݙ��E�g7���浭��~�*
�,���
�u'YD��O�7l��ᯰ>d�C��O��}������3�<a��~�����?7~��8D?o�u�����k��$��'N���N!�z�T&MߒVN�d�e�I�(�q�i�ky��q�rÌ1���8}�:�6�)V~ύ������W��g�y��^�*)�O<I���a>f�>b�ku�jw��q��IR��N0��%d�e':���j~��d�y����� =���G�~��U��e~�U���~��0��Xvs�xÌ��;p��Ğ�y9܂��M��P�rC�m�]��'Rk�d�*I�w�+'ψ�d�&߾�he����'���o���+��Q���˲-
s?Cwo�x�n��:|DF$�5�q�3AFƒն8��T}\j7{8�����<>�uj���ф��黠�v�*�h�t8 5��+�IkƸ
�8ӵ�wx̱VmM(vv�]z�mc�c����0l'�e۫͏��{���|���'��B�I�=�u�bV��a��h�ri'R9܂�=Af���'�9��I8���2K�q��N� }��sϻ?U�|��|���߷�>����a='{a�M��y���Ou&��6�̜C�gY&%a�sxu�c����N �4s�=I�M�a��p��i?Ou��	�O5�E�������o3���}�+�I��Y>�q52Ì�����N2�O��I�ó�i��_7�$�a�}�PY&'�9�Y>J�k���6�����5O+�����~�����@�'N���N2k�2J��l�'�XORi��a6Χ�?0�	��i�N��Ow�I�d��z�I�a��p�i�m���0|��yy���{ח_}��'�Y���d۴��́�O�>������'�d����XM�I�h�8�=J��Xu�O���~I�}�m�u�)뙗E��|���o<�9_7�a8��;��l�I��2sv��2u���{�2�O]N�$�� x��c!�YY����,�$�*X���G�t�w�]���*w��}t�����I�
�X)6ɴ���0'ue:��'Xn��Y>}a;����������u�m�3Y%d���J�d}�K���"�����x�̅�;�[�'�x�C����qC��%`kϰ��q+5<�P:��w�;��u���ì�}I�'���'��5�d�a8�L�IXm��^w�ˇ^:y�ǜ�ߺ[�����I�T��c&ӹLI:���8��'γ�8���)d��{ܐY:��gwa1���=vɦNsnI:�'9���Sw9�{���uޯ�7�IY&ӧ?d�����0�:��Hm�u*Vi8��ى&��C����y/0<d�'_P�}�	��g��>g�GԘh�}�W�}���]���z��{m�Ȁ9�v^�@�J7��g�ק�#��>���o��r�V1��r��8�����ӫ#�%�x)z�𳓪[�������.�'�t����T@-��A��4.*����MG���S����>U�]��7�� Q����0��~�N�L�y���i���J�����'R~-��d�k$�'�3�	�hϰ>d��C�y��z��k���^�%��mw�{ߜ���i��G�~�����'��$�q�Ě|��!>f�59�E�q��IPP�nϐ��J��2��2|�a8���Շ��8���^u���~������O�Y|�]}.��vN�O^!�gp�'�'ϝ�:ɦ�y��M2|����N��Mu���C��J�$ɻĕ�䬟����|l��7�߁�����x\~�������ꇹa:�G���&����>d�z���4����i��0�wa�&�Y����Cl����u'?RVV��x�]3�PS/
���W�H��m|r��OY>&����C��'Y:���!^2i���I1��w'Xu�p�1��)��z��v�Rx�j���}Su�9�@��#�J���u�"��O{��d��I����=�C��d?k�Y<d����u�L9���&2��sy:Œb~�0�'R��Y�s��߱WT.f�u^��\��� x��!t�rB��������q�Y.�����'��:��a�I��k�d�!�k�=gY<aĞ�� m4��o���*���y��xsڷ���>�#﨏�:~�J���i'=J�}��6����$�'��d��	�|���'��,8�<z���4��'�y���N��G�{�������zh������I�$�Ӛ�O��Aa6�{̝I�VC^w'�8ɽ�=;�l�2h�Y�I�M�z�M�u4e	��&�S,�$��-_��^������{��;�_��?0�	ٮ���'Y<u�m�u�z��$�g0�i�z��'Rq����'Y6���y�z��|9�IY=`~��z�O̜Os�> ~���Z��,Z���PPa��
ڵ���Z��..���6f�����7���j�ND��vWLy�Pܲ��W*q2"��� '��m�=άAk���vT���� ��1l�E�(�ܓ�#.a=����*Tuf�e�-��U���|g���M�u�+F����{�|�y:�7����2~O�(m$�*~Շ�L��`|��MO>�6�:�<޲�:��O�'Xl�2u��l'�;�:���ׯ���G~�򷿽"��c����JɌ�(z�����k,�������>a>B������f:�!�>�)8�ĩ�9��a����_�'_����������g��{��u����_����q�$��d�k$�$����C���+'�ÈV�1'�ˌ�hu5�è,'��}��N2�4{̂��������������}���pOӮ��ݪ�1�t�6å� ��M��9��'_�4wY
�6����VH~��d�Ť6�Rq�ˌ'�8���:��'γ�����	�c��_��=J��lt� ���z�Μ�H(C]�~d�'�N��M$����q>d��a*I�~���V,&Ct�
��
Chq���}���!� ��`��i^�]�]�|��s���}'�'��!�'}��2q���=7�:��	�i�Ěd�'ƻ��8�������ɳ��V�~���T��2?}��~���#$ʲlw�n�Ͻ�����'?'C$���5C�O��k�̜ݐ�ì���g0�'�&�ϰ�Ԟ$���I��'�?'��Hu��h�I�;y��7����������׿|?��	ӷĕ'��*�:�������&���u�I����!]�u�N$�x�ɝ�L:�9�nO̟0��O��߈��̀O�}�K�W�
�S�f���}	�I���������J�$���%I�+'��&�:�t~��@�~<�O�u��=7�!^2i�'�&'Xs�G߈��rS@F�{U�L��1������1Ht9�AC��Af�9�:��4w�?2N��<�*V���"�����&�=8ì�d=��`x�'��~�: 3���� f��v���`��a�]���v��yp>�;#H��(��ql�v�	�,��V,1~�{�W�7tM�nvj�ĉ>�zv��_�R�,�|\���P��o.|]��D�;Yi��}�Wcs���������e^��\6����;��+R��<n5�W�9y�U�"��~��!��qC�������;`��'�Xr��=d�9�?2N0��d��sF�E��X���I������8�{��sxw��9�߷��~��t>|I�M��>�&�8���:�|¡��a�IS��p�'�,s���M�����
M�~�^��u�_y��|~�����?}�����0����7�᯻�&���hi��O��Y�M��Ow�@�i��/��a&����Aa=C~��q*�٤�$�������?};+����������Ы<�?��o�ӌ�2z����'�=a<O���$�����L�b���Y&��'P_7�$����'SL�l��a�N%@� ������>�����?���� -�������{���'{��Ld���i=jƠMe��8ɤ�Y�I�V~����C�'Y<�ɴ8�Ԭ�ް'u̝M2OY���Χ��������kߺi���S�N2o�N�|�:�=u��Jɦ��������P���N��Y��4�Y'����u�S�p�'q�9��~������s{��W��<a�;���N��Y8��y�m����?Y6�|��d���š�+'Xqd=O̜Me1�m��P��]�_u�<|�.Q�e%��_�����R�;9�I�O�S^s$N��>�~I:��fN���'̝��OY>�N0�&�k$�6��hz���)?K`m�q9�s����������o�ޜd���v~��?2M���q��X=��d��{������>v����w��i��鐜g̚��m?��T�#�o�О����_���U����,;l�i���|���j����>o�8���Ce���d�=7܁�����~d��'5@��M$����'�A�ަ�q� �-q�-S��E�i��V�E���]�:1��"�thګ�<#�.\N���|���;�tz��7j۰��(�[���\�;-��=F�N��M<�'PY2�[VQo8�R�J�+t��zd[���^njP��*n?���_n�O.W�i>�T��%AB�m
��
�8��zRO�u?j��d�g鯰>d�A�0�v���'Y=a5�g^2x�g��'k�j����ܫ�D_�����~��<�$�~d�<�Y'P����6�%d�VO2��N$����q�i���q$�5<�C�1���<>�d�x���$~��g��w�������~�����nd�OP<9�'Y�O����`N��Mw��qӚ�*V7N0��%d�e':���j~��d�~�y����P�	��^U�*������t���g�a��s�xì��v����=@��r
�6��w�!�6����IԞ�̒�I0��
���d�&�;hZz{�T�������X����	�4��N����
�&�{��I�Xl��u�XOɮw&�q!���(q��k��'�?sY?$�I���%��8��Y����ߕ�Sv.x�W����e��OM<MOl8��C�י<}d�{��>f�:���βLJ��7�PY&?����8������'6����������ત���U߿^�����Y�N2w�d��$۠ݑa��'FXu�x��<��'Ƽ���'�8��~d�L�b�7�$�a�}�PY&'��0~?|�G���c[�܂]���ںط��>Jç{�z��M���N2{�%t�l�M�a<}I�h�a6Χ�?0�	��z��:��8o̓�4��ò��i���μx]4����ާNM�M!��a�'R�<��8ɷi=�w m��O�o!<`{�'�d����XM�I�k,�$�*~ՇXq��ņ$�@��.oO�e�~��>���!�M ��Bq'�k9�Y���<��d��'�w�:��i=�l'����+'��)>k'�B��:��g'�S�~�<��ӏsS6y�����m�OXe�v� ����j��F�a����z�慫w�n���gUJ5|�G�>�]Ӻ���)����iEY1��U�1��_We�Ŕ����n�z�G�ɘn�=�s2u'�s��Y/m�Ŗ��q/4mX��Ծ(а�� �;��o(�ٙ/;E����v�\�D�H$�>f:�)<�|�P���G���6��G�r�k+3��v�n�'��r�EJ��T�6r^"jM!1[AKR�4���]3fm��j���(�Ӯo��x��� ����غhn��WD��^m��Qy.\�a�yS�*�;����T�Z�F����ʶ�cJʶ	�B;j��q����t�|.��
�Ӆ�.l|	����%&7JW�Y!���]���um��n�9}���,h#�J�|;&�0$ic"ƙ��IQ���86|�d����#w��䮄��0vrS,
o_K�.`Ldt���u��M��/i���`��Nԕ�W�����2������]��o���Z]���v(��7�8� ��.*E�η�Y����]���=Z��-�j�@�qj��:��Nhiץp�����X/�y������=H�������n���[=M��
}z�ζ����6�<�r��54P��J��7D{����^P��5r����!����l�|-�P���R:֕�9�����ug��$�G {\�OV��x�����d(5	�Z���7�AA�R���U��NU�Z��@˷�b}�ϯ*v�r�S��y{�ql�c��X�ܸ�J���l����<����n�G1��ޕ-x�rp�S+��۔_bo�[yL/��`�g@��56t���z���C��n�,���4ld���y���g3M�K��*�%o���V�AE2�]d|@���,��y�,L����"i)�T���2i�e�c���U�@'k&~��!��;�Y�A�����u֣�AB�qQ�^��$,1�]��V(GG�}y�����[ŏB۬�5�����+\��An�4h�����w.ϵnM|��	�, _w�9}�q7t�cv����sB&��Ɗ���j��W(���q��u��ו19�J�'%b�ξJ���2�ЗX�o,������6�bF�A>��I�,o�6}�'�L�Fa1�K���o���VL<C��4��Y�z��K�n�0F�s��١;�g�e[Ɨ%���:��9&���֞�n=��G��ݜ�ں�J'�K:�oS�З�{E^0�T�����9T1N�^a�{zO+{SV欭i��|��x^��އ�h��J� ���%��"�WF��J���������ʡ�y��P2�T�.e�A;}e���73櫣���ha�N��7j�Ʒ��j�j��-G��`B�$	���0�����m}�-\�z�\�$����!�Pq�ހ�h��s��L�F}�eוާ/4�|��;����u�<��ȹ���U�P�P�Vʶ��AIDPU�FiX�Y�F�-B�p*`���*���j�+[*Im�R�QFƔm�%H��X[pB�mT���"�JS�+���0�mZ�eee�`"���(�Ȉ�m-q�--�ŭ��J+X���U**�%F�-B�V�J��)iVեAjT��R���B҅J1ZՀ�)Q�P��Kh�U-B�
�Q���6Ԣ	�V1
؉mRҕF嫔̢�#m�V�FV���m�*V�-[YF�%����*����Q%DT��iV2�RڍJZ�QDQmQJ�[m���k�ŪZU��ZVQ�*�UQm�Ah��˃TR��R�)iQ�ЫD�e��4mcm�.1TF�JZ"�X֕KDc-�LjDnXfE����ڱ��E�k-Z�#mZ[R�a�U
U�9�#eR�#L�V#m(5}������v	}1MNKk�ż )$ ˥��J�zN�4N�X�i0]��B��P�s��M�0��Ho���|˼��6O&�υ�	}��k=I�9`����Y�(O�u��f�N��/�u�����:��x��y�u�z�3Y%d���J�d}����߱�u���G'zot�����w.2OP�1�RO?o>d�V����'�G��
P��d��I�^a�N>����ߜ�z��G5�q����o�CX�5&���{����1�����C���VO|�L�>C�'FSM��k���I�>�q��Xy�Xu���{� �u�ܝ݄�O�*�__���KI�����~�7J0j|/���I�ğ~���i߿d���ŧT�A`�6�Y:��1��'_�|��'Ό�!�N{d<��2q���{7�x�nT[wV��	���X��y�x����.G\&�D-���Xs��vڴz����o��e��اk��dyy3��xd-�.}h9�*�`�=�V��t�[�.�7�����K�I/��w,:�Z�k֏��c����3��J�����v��w9�K���^	&����~�/Wdi9WJn���Le�:�����'�.����� 2��x^m��v��T��=7��J����+D�6��Q��{����`o�_Ǚ�9k�RVjvʃ׈��1]�O���;2u�'�#�uv�rq��wț�C��Ê�}�{:�����:��i����t`��z�`W|��>m��DQ�)v�s�݄�
ȹ8v�4�4��9#��u4E|���ځTƴ����r՘T��R��_}T.��׍љ��s3M���ҙ�a�cE�5��|����v�\����r=	��tߴ�������gh_�Y�ו�zy�܎�k���prv��/bS������o�8͌��}&���x쿗z��pw-��%5�K��>���y��={ ϶�XN_�8��s��=���_HV�b�uն{�{�D�2x�v�{F��F,gk�i�N\��w��{�Y�{Nl\��s�+9^�L�?8�Z63�f�c�S�����i*��O�f�v�f�����]7�gG�g��]A�|��dx:��f���;��Mb�b��zL���Ǧu�gh::<Xñ�S���%����CI5�~1��s27�1sy�	�ْ���腼X����W�Q^��t���s��UE��ǣ�ʻzgs���yx.G��\�춈c���B�<�tC���P=��j}*����5_�����y�Y�t#X0�f��)r�s�᳇wҦc���u�mv��b��N�� 
D�}V�+��[�۹�,f�+�6&+�Q�b��i78�x���z��m��񋩬GSApIܫ!�T � �֢�M�ќy��s�j>�}����k��T����߯����n�v'x�K������
�ln)��&�x֭�{DA��K�U���<㳛�i��j��}Ґ���QV!�ٍ���{]\�V:�Z�7�;���UE�)sw�������۹��x�㑔�lv�M��-�2���ԣ���{���<��|_�`����/c�rذ��g�ӾÏD���lXY��N�n��no����zq���89����_���q��뜣� ^�|��m�@g^^��=�S~��`y�r_xɞ��7��Iu]W^�G��Ӽ&��0�y�^|z�)��W�b�_�OWow����aS3��}�y������ y�z�{ơ�^�?%�LX��m�C��39qtN�e�nN�y�3�s�&���2z�Tn�q�|��O�}l*� R�1e��r|�T=���e{+��y~遏�[W�<·�p7���d�>�3z� ��,f�ӕ ��a{�9�p�;�`n>ů{+HL�+�X�ڔ9h�oo�O��E�N�"������tٳ���WW-��؜"�,^����w���%�v����Nt�\~���|�1�^������B��;��<��g����'Iљ�\���B����D�vi����u�}�j���-���Cѝ��7����=����]6����c&�L0��� u8@��9�I��;��]��3�͠f����Kdx��7e;�����=�l�h�5�+�Ϭ!Ҁ�.��Mϋ�����:@x�L�=��T�$�׋}\f�x;#Y�>��j�'`ck��魼���[�I���z/7 �_������&A�+Y�@':�S����W�ܬ��6��[�y���>�.�kj[�}?g�
�rM������@��u���˿v�^���^��s/�<��[�y:�-��b3�I�5�T����Y���\�*�}����AK�����{�f�E�äa�~0C�E���^/t�u�l��X5��pg.�ػ	�A�����\�Co���{/�,h?-�Z�호n��t�'s��3,�*Ē��]��L�2��L˶�|닣�MN�����ѻ+<�롌n��y��\�h�b���t}W�-���U�U6��>��I_W~��\��|�K����L~��c_�>�0y�܋������ga�WC�f�&���e�n�~ߎ�Ul{�=����`v�0@O�7��s��zk4�u���瓟Mi+k�(r���##���Ӽy7
�Q�7�mC@��c6ܴ��#�rk�}3}(�gv�OWE�˲.��x�����ic�{�p��$7����\�ӽ�I��=7��*2�8r����p��f}���o�zX­���bP�tϋ�����e��Őo(;g�XS�}���|d<���`T�<��1'��A*��Gn��Jzre�e�Cc���չ!{a��������	��]\z<�^9�Tq�J�h���{��:ys|�)���w�ô��՗;�S����0����E����U�����ps�VL�/λ�n��0�{:­�|�|Ϸ�"ߏ���V�c�j�t���YxE��{hۼ9Z��Eͤ{�ze��Y��.��2��8�����wS�U!�س�p�=!̙m,�07�cr��b�۵B�/����*ٻ�i�u�O�H�xh��f�/��X�×�s�l[����߇�����{�g����q���[{����/;R�$���.�A�7쩌���<;|=,o��p�*��w�v�o'�v���`R�Ϣ��8+E�4g`�y�|=\s��Ꮔ�[��u��30�u�н�I�wc���G�*]K�Ɇu�wz���f�G&��@��m��&h��'��}y����0oDI��m{w�RN������q�3�{����	�V�����S�����oZ�ln>��}���o�U�9���`�{�*�w�Nu������}��v�����z�9�N��Wl���y/�����ɏw�M���c�;+��������H�]^nuq��U����Ӝ��dq��o��]'�rR��BPu�8v�{��+`^w.�p!Z#v�p}��.q���=��U�W�0���5� ��wv�R��@[��ᱜ6{�s��%�)p����+�f��	���OGk�QŻ����%b�7V4��\��^� �X�)D�r.�NP[ʸb����y��O)��Ν�XT�G�>Ѳ��N�[�\��r�.�d��ʈ;�sX��.ˮ-�P��9��)��Y�1}�o���� ������ӭ�����&:����s:�;<*�l�e����R����ɱ��V���n=3�Y���>,Q��%���Jʽ���ۇ��OgMk'�Y�<s}�J���>���$�Y�tF�귌�v���{)�mI���<(�V����:v��{_�z9���)���C��ȉ^�T��?ft&DpᠶB9��_t���N���3|.K��K,r��e{*�s�y��rX��YY�As꿩�f��8�n<R���n=��{ɾ��O��vֈ��0J��x�O}��s�,�r}}��%J�75ً��L���Y>sdTŸ;E��ۙR�xLʕk6����M�ui�z���&���}�����{[�Ÿ��ϝ'�vw�f�LT����o.�l�����A/ח�7�oN7����s�N�[�j�v]Ͳ�b�6�կe/=l%\�0��d���VA����],�UΟ#\��F�RtFi�A��º.0�4�zQ(2�����oN���[غ������oZ�n5�v�tfRw�+�F���H���X���Z�]ʝ�K=������|>s��v�8
�}��睄��\�y�o��k�>�l8���;K��L����%�����;��}H����[�����VǽK���K�^�F��ѫ�C'��N���t��qO�����ۿW���Yգ;\9飺���c�Xۈ���M�f��>��o�OZ�}�?��ȝ/�W,d��k&�[Q�5�=rZ��������ӽʹ곴�w��7W�g��:6�	��g�Hy�J�ۍ�bCc ���:cS�N9�]�����k�R�^ѝ��R�=�f��S��͛��$݂0.v�Ϥ����*~!�Dw�d{����;x�#p�;%�9о�����=��-�e�9;���j-,��S���[��f{�D-�ϯ�:U�u��MϾ/3\���Y����7�+f�Ϧ-~��پy/oλ��n��a߂�փ��7�s*{�hK����*�-����G��>mh����4��� �� �+-K��4�j�t�Hf>����Ƹ	��@U��[B�4�+�;�j�{�Rʷ��[�}E�&ҀV��\My(;�j�#���߯�.۵e&�V�N�[]�����%�Z������e�z'Ni��߻��R󙕚�Rl���k<i9�V{�fo��U�<�Vk����7ytϽ]�mG.>S�xh�m��Է���[<�ל^�1�=�3��^׮>2��#�J�-����,F}�c�w��k�[�z٢2�޿S���v��������ވ��{�`g؉�{�*�H�������R}f߅�.�����6���c���K;�f���.�:��Ͻ���'����<�	�>2ۣ��=��Hm%���>�xi���Ϸ���a^�t����o�ޛ�[��=e�����ug�9��up<�����϶ܰ��g�ǳ\�K�O�����8���s�g�tVn��7Y�N��haV��88{�ƥM ��d�k��g����!��/YG�����2w����'��� ���xį���7C�O��:.�MW�d�S�1��.��v+�U"��6�ʸ�*�O�:�o�.j�N�5��gl�㸁��RB���(k��[W��[U��ռ],�&��S��J
7G =�Q͔5W���R�|��;l�#1�R]��k��}�)SP7�g���]�� �[����ћ�|�;ް�1�O�Z�T����y�=��+�wu�&K��z���N�3>zg\����(��������^����T��n���;-����*{z�瓲�������Ō���<�u�q���A�*�_���ι? �������ܜ���w�:݆�q�!1{";�+{7�j��un�����~�9�KΆVI+j\�(=�.��տJ�^u{���`�p��uS�͉���s���諽�
�����ν~�l1��&�X���d�%|7�a{+i��o�z2����?e�t�|#��g��H}o����m�S�wP��:�ʡ̡�u�����h�Yk}�=�Uy�u�F4)э��b�W5�a�T~���GۀY�P�����կ�կ�f�k�{��*�s�u�KW�=���՞5��w�i��ܵ��[<�v}�5��;�]��X׎kE53f���,P�0P�4����oV�ż�j�n5��bGH�ٳ~�ilWv�f��ʇ�S<1����Gl�M����aV�U����Bө������C҆�q��iE�JO��[/��nY1�<���FS����	���vW�YL��7L΁�u36o��{���}S,�˳ ���&�� �Õnۧ�5��P�4��Z�ӣ��DU��˙Se`k;�fn�Jw���r���B�^	����ռ�ou��wN�u�T�a�Y��7�m���v�V�	CJ*��ѥ7���%�E�w�tb�wwԱ�V�Z���
'"��Yudq	]؝�J���y��i��=Ú���V[��,�9�س�KJ��sWi=�0�c����x/��"���r�&L��y��d�ʳ�{���u���MX��V�a��ɚ�X�E*�,�Gs�=K�Vq:�e���[N�]W�]Z����΀���ܽy6�r�.��ZI��RȜȭU�E�C<C����T�Z��n�M�9J�n��+���Q��.:\�
���Θ�w>�ZJ��x��a�8�ᦪ�ݖn�R{Ӛﻲ�WB�Ĝ��8�Ax����{�9'�Ӓ]���]��vMa�uz�)+S�mݭI��ZV���z�� �(lT�V���d}|�Q3)��;����4��wZ���g:�l�e��W[����"F.���ń�	�3-�u˺��ji��5��:��{78�n��2L\��m8���P�q����Uue���ziڸ�Xz�����Jٹ�r������8Q���tɊ�|oU)������qJ��$�tNW�m�4�n_uY$ɻ�1Y�� ��h�3�R����EB�p�]1����xL�����1��7���[?���6�U��}/w�x�X//��̼���9R���q�@�k��T�
�O�'F;�I�Ԝu��HY�2�u:��v~���i�bhL�
��]�]�/U��hbuE(X{���8_Tlm��og��#*IE�Z���h�þ�/�6�f��!���zt��Gl�0Q������l��*����Yt���bC8	G1����-s�rct�����c�����JyV�H��|�fMr�gA�K��ťڢ��Pu��A�G�B�
U��	^�.���<��pN"�bx��e�"p�R�`j
s���b]�5n�*��^sYJ[��6�vrW*�#TR�@��� _L�|���kF��7�o�G%gf-RY���[5ә��(T�Α��Ky֓�|5f�:\�J�R2�v��,6006�^px�k(��Yx4��}I�RL'�.5�rş�Y{RwϷ#F�%�G�����yn�C}��#�����{#��=�{��ۼ��e�	\� ���H�Qj#
��.Uc��j�����2�cHԫq��F[*[km�*�U+�\m����-�R��elU1��2�-�aUV�����[bԩmm���-��A��������F��0F(bjVW�(�91������ԣ-��Te�2�TnRcȥ����Ak
2���m*(ҭe�Z��ګ-*Ɍ�i�ʖ�V�Tb��q�֤�.+%VT���J�+�qX�1aFfS�KQbсiAk�e�,�X�7(��L`��L��,F���T��r�-�X`�m�+"��RT(�Yb��Ƶ�A[jfP�ĶU`�Zʨ-B��j*��
�mPYF�A�,[l��
�iX֢Q(�UE*T��`ۖ�E�����B�E(�h��j[me"*�b�
���FӢ.\����я��]]+�1��A0����r�dʝ�]%�Pn�޴p����7�p����y�UB�o��|>�����Y;a�pc���/k��^�޸0��c�3�߽�o_^˹Bb��W�~��F�YGr�e���W��l`��i�9~�#���z2��V�>9����=E4����1=��x��^wjx���h�{;\86ܴ��F����Z�{���n=��ѷ;}3fⳝ�3���������w]���A0��J��\~�4��Y��9	��?nz�>̝�~P��K�R���w��1(\�0��Ǧt��tv�>/���MXf�Ac�`�=���,����㛰G3y�	�ـHX�v�tA�����N�AWD��~#v}}R�G����ι�yyr<��װ��9>�U��'����7Q�ϸ!�������f��#�׆�񼙮w��{ݎ�λa�vB�x���t��lN�q�kq�3��v}w7�N���uV��m��ڈ�r�m*�j�X��f
�"�(:��5�E�>�����ܷۻim��7�nn�Vܮ䗼�,5�E�-;[����-(���)�UN�r݆�M��w\qFޛ��Y��.��4_*��������s�^~�e<�ܾ��0JvN���I�sc��׳.�||��=��)���t]ȁ"�/�hr{Dʖ�e}ò��Q��&���������פ�vOl白����%�n��gΓ�Ï���c/{ld��醫ø�t��*�;��\��8�����1��A����<��L^e{^�����~�6f�+�x�;�V{�2��������'fo���&��� �x�{oo]����߇/o�{6=�+_�O�s4�g�Je0����;��o���9��=�7���\�y������߂{+0֥U��9��}�g��'/�6G�>��o����}�3k������s��\k�r\�x����;ǡ��ܷS�|\~����*��;��������7�ΧD�pt/�6<ć �I�s�zYs��ڠFu�~u��(�Y�nfS��u�}Z�Z�o�-������Yk���Җ�v��+�b�Ud�xy�5�e�Rs�r`�W�԰����b��m��՜֜�%�TT�ò�홱�>4���"-ɰ+����'z��>ɑ�����UW�}�q����������C����J��>w'�`���X$�o^��Jh���ެ��~،������;G��hs���]�����M_�u�*Z�]���Rޔ��?{ն���Gv&BQ��>��C��~�����7��xay��}NYo{K�@:G����g]����a<��=���w��x��J�^OJs��ݧ�(�O6��K�9/�
�lK����w;҅y=��+��f�w�Ɍ�K�˵zz��y����r�����X�m˩&�=z���ޒx�ⱓ&�	Ϋ����)�b=$�rذ�~=;�;���+�l�)]?>�^�aɢ_�R��r�L��z�#��8u���5�S�ʌ��h��u��ߦ���)�m����r���r�:�&>�@ќ��z�^�gs�5�������cӑ�oog�޽=v���|� �n�X��W��h��=zv"�ǻ�1V�][ݖ�C֪�NC�H@�f�	�F[��ݾ�s����*v�ɹ6򮲶$�rQ���'s��{�:9wSa�ϯ�JV`��w�q+"ֱ��u�Lԥm��A�h�����u�*�����m:O+C�������<$�Hw;*�ߞ;c6�:J�9���jy͚֥y���w����7<��ﺸCf	�_[����m�i��{�\z�Z�^��:�D���c�o�<�z�9o<�l.��B�F/88|���\;:I5����M� �c���ݮ��4m���Z�w+~U:�]I{FWd��gx�*���5�3ͳ�>�ݫ;G�K]L�~�\y��I��{G�%c��ۅ�l\�Em�f=3�Y�����b�;%���&A73�nTQQy�~��JZ�R�X��XN��ؘv��Ŋ<�:�T3�}�ߧJcx���X����o�)}��Nyy2<���<��6�3����q���Z׸�S���tϓδ7��������ϔ��_�I/�.K�6jr�Yq{ٳu�Z�EβW��4N�������c��b���Dw6N�~�Zn;"�wq_ǎ����<�Ľ��{�$f�Z�r;��e�����JA��I��X���S^]L�Yf��zz1��Xttp�J���+��b7�|xS�U���;E-�.f��:ܜ���!�혰V�ݣ\�a%���6�F�o�nuB���}U�W�a�z#���l7��:�tM�=�����H˦=�Z8�F���;�L�yZ�b�h���t��z%�Os�:��y��,�k����s�^ɺk�)��`o����G���Jp�8�G�X���1��?g�����[N����}��3\�o�U�q��ǧgk�_���q�\V=��f%8�{}�-���_����~�y��V^H��9��ǻ'��y�J#f�^q�i�����z�?�0z�A�m�	��GI)���6z.�)��}�L��<>���������Dc;\>�����1SA���{t���gt��=�9�"�����َ�<R��z�kV��\BS��F���;^s���с���t�\~�oε�>�����x��v�'XבʻͿ{��<��g�ߠs��%ɳ�s�xN>�v���Ŏ�0x-RYa�z,�>�O;Nc��}D��_K���dUE��׳)Żs�P}H�����\�qz��9�I��pK��en4�[i疰.���7/��A<���i4��Fe�{T���}ه�e��eX��@[;�N�qyӹ�4�ee?~�� �~�:w�^v��>K6��<���o�	Bf�f�d���g}�i����C��Y}3��2 ��Ihs�}N���v�8k�b{�]H�蘹m�n����%<�8%�Ch�5�is�F�ʞ�_=�d��N�ZK�g;���69Mo��Wmm@�\���
�k��K���v�_�딡�<��_O?f�`�������nx��v�3~U���C|�L�ve�$��\U�z����z���e؉�}�iN�y� 7���a�ȃ��+�8)����˳a���a�}����벓�����Q����\�>7��h޾���0RS�"�I���(��$�tؙw����ݓ�5%�H��]�a)�ٿr�_G]	r^�C�C���,మm�ōy-�X��z��W�1������)+�8�f�m>��X|�\LpT���f'�wک߷��ۂ�Ļ�ЯQIR��p=�n���cӱ�a�^-k�<�9�v1[Vx�f�0��չ�1�mR'��C��6k�h�]3��D�ḷRXl�5(�}�X�92R x��v�Y�s���C3-)�М_#ԩ���:c
���|�t�+v�����;.�T�WR�=����}������W�w5����8#��������N��;���A���)�E�{)�>��lܵm��:%�2R�1W�_p�ۏfkN���3���a�\���f}N�->�/T�^}��,JL(ۡ1Ғ�|&�ۏ�f:Vؕ�ٰ��gR�h�p!���J&��+w;!�N\�ᩖu�Fo¬ޒ;}r�V�k���f�j��Zo�UT2���M�:&B��J1_�N���t�Cܗ�[��O=<�`y�$�rP8��P[P��\]J��S�86z�ձ���oi:N��+�*���l)��Zf8*r�����*#I<�Z�Aqv�&]9sW���G��;�;��x��Z���ʕ���ޙ�}�g���{�Aڹ���.�"�<D�\�e
//�f�40���5멃]G��8���z�?�����zrNߗ��W���d�����'A_����Z/oގssF��=��g���`�0s�R��?EB���*b�R���L��ǋۨ�=c}�>�cUi4�«�VF���Y��i��Qps����X��ʕ�:���[�(N{e��v��#Ƃ�*�~iˑ����t�6�>��={���z$�^�W<�K�Y��s����
�w9�wa{ڀb��t8��
.Y����n�:Y������K��V͓�a���f�.�(p:8����zu��k݈wb]Cj~�����5l�S���n7c��h������N���3�OϭE�zU%�C[����m��U�f=0z~�H��J^W�v&��(q���<�kդ���Z�v.*�'�4����l��~x�]�xx˼��)x]�Wr޻�S�v֌�(�!](=+=��Z|�����nI&V_�\��)�n�&t���������Y�w�^�؇�r��%VHk�m�\ʋ�^�o.ͺ·ݫ�$��}��v(=�卋�Zpy�ie_��n�:��F.��g�*Zz�W �t�s��Nb�_��Ĺ˃�M���Z�aşS��|%B�Muj���s�:���F���pt=�ۣ�B05�u�U�mg�ե^K&���a'�陁ܼ9O�g�IZ�����u��Z��u��VZ�F�M#�Oi�t��|)Ďy��/J$t�IU=]5N�G�_�Nm3��ֲeC2��!ai���y��:S~gDG�3y�K�7�pk;f�_��Zl?z|��d�������Q��H�˴x�L��"y"9���+i(C�����pI7�
��5��jY*�÷;
!WtMǁ;+�6���5���-v%�Ł43l�'Iǎ6�r��ټ��C��H���J��`JՇ]t��Xt(3��墓�ɡ����Msj�͵�a�7x0HoW���| 
��#�6e>��
�c�M�fw�fNv(�^ܬn>}�dhu�
���  3w��$�1�k~�yƋ10���:���5春5	9�b��rfŏы.���p��I�~��[���^J���"�
__�ݨ�C昩��Ɋ�H��G��:4%��Y�&���PL%̴�ґi]:���z��w�u�����ʙp�(W+E�S��n�<����7��ɥ��:�JO|��CY]�q����Y�C��<�v{��X�d���.�����*)���SD낟"a'D3݄�v4T�E�ͪ�t�o��:-j��O4_l-���κ.{k��@h؊�!��`���
�x�U�Y9���D��ab=�7�[���g���o���C�c�}
��1��agTv���͸g���@�t�7��x8U��(.�q��l����5�0��lpX����J�]˚�\}�f�����|�&u��}[Hv����\������Uq������x�!Sw�B��C{Z���a�\M<��q����TS6$=�11��,��Ƙ�� z�\]���֛���^�H�{�	��P+9�9t��ޱ*�_-.P��U����yH-K��Z���x��=�J�mÅ���n��A����H<;���S�}U߇�|���M�1�*�I;c���T�|u�.���4/EB���Đ��S�k�����xϠ�ه:�3���[�뇼+-aTWKցhj�TG/�����{�{���4퇾�pǢ�k�f[������8&�y\Z�GO-5Ϫ��UXT{��|¡��>�p���xP�Q���ъgޖL6����C���>&��ؗ�M��*[ �\��ԓ�t�b��km$+,{���q��l���r�w�g��;o��M�S\x���SW�=]�-@/Ծ�/�fc�'��@���S..7�Ny�fKcY]��N��7{�])��4H���:y(|��yB��2�S2<KT}EY;���0%��!�r����۵G�L�z�:�U
j�/���p����s�C)��L�z/]��R��]qwcg���i�P�#�eù���( �p�#�>b�]Y7��1}1�D������{e&� ��Q���?Evˁ3��v�˳|�#���f�҆�� D������T�+7��*�����l�HOj����&Nfp��\�ɽuǷ��f24�P�=9�󤒲nL��6V�Џ&Y�t��DT.�
N:�ҵ�J�J)�b�lߔ��ma䂡�9�0�v���aN��ɓDư�l�쥹I���WW5�}X؈��9���T���At}�[�I�\�ŝyMFx�N������;�[�v\�E'e�<S �6��N�ke���#�vW_S\�-ZɌ�"�J�cX6�=���D<�7��e=�Z�V4�=������x\�IP�A�mc�iۨtS�5q!���]�pSkdi*���F�(��p>�;:�j�.&rK]�kL����W|�w,R9�\�ۢ68��m�}���}��z�Y��#0=��7w����b�Y��d�![�u�-J8=|F�+�w>�7�����гj�i�R�GF|ۨ�H��ꊑFr��sV�n�ͩ��N�Ou�E�t����ew΀��&�� �j�ʇ��>�%��J��V�rժ�+7��I��n:��1#�Ǩg[�;��@)���ڥ\J�2��������A�����k�J�Z��	��%q	ܫ����(|�i�E�lӳ�����ⰳ|��u5�r�ī.�V��3~����zC��m�[�89�1I»�@;�Xi���Ǐ-���'�:k�)��6��Or�m�V�;��u\�G�8��7Ik�{C�fn�.݁�R�Ю��T�e6fZMbԞNBν�*�5'N`�J\��G����������2������Tuw"gv$;���� Ծ�����I����=�JW[�s�Ө�Қ�0˷H*3���8�SN w9�ͩ����K�7*h��D Qi�yg�ng���5�#X�Z�#�uo�D�l�;���qu��d(��CmiWkm�=�ԡ�cwQ�5֪�0�.F�h*��\D���怼�,n[��p�Q1wee����b��҇D�_P����W�:�$����N��&,��sjV45d̕����%k�^ee��R�����=}��;/�n�|��k>�}ϩRÙ��n_P(��GիzF�7ˋ�ô�jh#M5ݒ�S<���+{�d{ՠʺ��DG%dP{AW&MBW��c��Ve--�@�WR�ycy�\v.�b�u�&;�ǵ.
�biwS��ׁe�T��7�i:��ʥ��?e��N	��x�*B�2���wE�5>G��GV̮{�i�d���@K�3�)7*���INn��5�Ag1��n�V�E�N�̸��m*Kj�)����z��i@!˻�=c6�6Mj�Kq���_^�99��B�c�\t=[X���*��.hh�a���E�P/������lf��(x*���6SS,Jb�$(j���A�;u�ٝ����+�8��}]�]\�L��]
soF���{��5���(�Ww��������oWVo֐_c
�j�����[b*��Q�6ڵ�V�[V��ihU�l���Q"�
!U��Q-����"�
Ȉ�2�*T�-b�����,D�,m��X"���X�8�����mJfS-F��,�b,+%,��elr��ňƔ�+
р��TX1W-���RX�X[Uj�nDX��UDX��iZ���Z�(���--։l��
�őAUk%b�E�kE�(5���E-mcR�QUQ���+l�A�Y*6�jV��������U��*�YR�6�hƶ��ZU�U��Z�UE��YZ�*�6�UJ�Q-��EUAb"�R�"�h�m*�H�"�P���[J��Bڲ�l�*��"*���TE�m*1���b֣0`�-��""¶�ej-j�+l�TeEADm�TjUZ��U�Z(�QT�YX1D�[n��x����:.	�}I��A$ff���5w<|a�cה��Ť��&�9VH�ݬK��ﴹ����
�9K�����vh�w ��w/�aκ�n��,Ն{��3z`��9L��탮Qk�KGIܹ^���~�9jv{q����΢F �7����zg�ߺ�Z�zQ>pP;ʲ�+�{�^��ߏ��iN�+}S��iG(�*)b��O�	��`� �q�ǆm�F��㰔���5����)o̗�I"s��+�V�χgX���{�#,��X2���b>Rg��J�Klw�8L/�t�G���⳧<��sҫ,���b%V`Lt�/םY3�+��+2��ޙ�r�+]%t<8f�L�fe;����^���s,a�U�⨳�o�!����ݓ#k3U5r�I7�� 9��k�2Vˇ�o��&Y�t��)�5����[�x�O���L9�K�Z9yoW�j�����'P��r���;>�����N4^�����T�	y(o��Eqz˲ө=����`�wm&��罅�N�v�Uw��԰?�¬*�fg��81��l򷣬W���v�E�Y�f�^c�Օ��,c�����=]l�R�e��h���Og���
�Xc�ymo��v��%�]�V3����ʌ��k�@���p�jH�_aj�e;꽅 �*�� -����w|���Zd���| ����\K�,���=·�z������=(;V&R4�"�����[�g�(t�d��y�ۇ��u��,�=�5yO\:�)cHs�`�2[垞�s'��na�k�ȒY�%vv�����`T�7c�W�(��!A��*��3�`�0k��^y���*b�r��`�|(�i���c��@q�F=K�%�%��}Y���V�Pfd������Z�}U�\���m��Fյ��*�e �P�A�;+K�%�?>���+C�^���9=�ޥ!�����J$x�K��P~�Z,����]/-��pN)v��>��x����#f]�]��ǻEG;	���m�d��j��M�������UQ<1�9�3��Z����΁���9�Pz�r�p>�q�8���}����x�]��L�6�E��B5�k�Yᗜ3��0C�+�A���x�zz�����^���ҬYgi�j��'{�X�z
��gR�u�wp�"�nË9�6(Ys���]^�;��q��˶ކI�vy]\��h���M[��Py�3Ad�߇��K��"�>x�i��OkqZb�ɤS7!Y�gg���U�-����S�%�>�#���^qk.�J�}�ޜ���<����2Rڹ���m��Kv��v�:��>��S���ϥ�@���ﾤ��ӻ�
]�xg�aU�-2`�2�y`.�sU��	<<陁ܼ�Vq��7�Ѕ^r�ˡi��8K�x�j��Cj��+�>�<*��L_
q#�b�J�6�k��y�&vx]w���__�����{L�ֵ-Bi/!�x�f�#ir(l𻇍7���6�ݾ~�F���W�xL��Ƒb=�����̤z��h�P	i���AT��{�Ϋ]���S���x*Lg Յ���L6Nx(�sb��.=l��0�K�������l̬�D�?8�����š����~N��>��';�]=P�����y*��OfgCޚ^��a�H=ԢVS3I�cǕ�l��ֺ�lsއB��}�)��]ߧ���>m�
0\�ŀv
Ì��Gk��9M�k��D/�"/�U��0��4�s�U�zS�ϧ<N����;��E��<������Z�/~���{�܃<=]p�1{��T��c���Խꃺ��N(^J���=G�z��!��&��<�|�X֯m�����g8+WQ�J��r�g53�$!j��IHk/�w����b�G���Q�[��o�v�Y@z���x�M~���_N,̩�n���V�3k�>��, ��2�^�m��Kҵ> u`��ءB��ٻ1��,�yߣ�����{�}����e�y&��א�{ݞ�GJdf邓ۆ�����ԣ�|h�<M!�N������r���Y\|�{*�;Ƚ��]�g��I�+�����ά�<GK��чɏ@�ܭ�����Äa�<��*�G����ۙ߳��6W����-����Nt��{7+�����!��s��o�i	������/%�`b�m]i�;,Acy�1!�(�����\~�"��YBv��ԯ	�J(���8�[�A��(�5��X'ޛ]���w��c~�q����g��Nf(w���ꙵ��-
�ԽhXN������v.��T��ν�M�Icק�W��3�������8&���|^
�G������˫�\�vN��^v3P
T4���Q-tb��d���R���8��˱���]��5��&[1u/#`�2$��TF�m��9ձ��k;������캝�/>Q�f��nѡ�H�`�şPL�uD�hw˲�mo����Eib+������,	�`��4z�1��ei8��'A�2�1X�v��y�_�xk�Zux��=�5y�m>xBF��-���6�6�ϬAUx�>� w�M6�-a>�ɡ�t�E���=l��� ��Z�WH�5�5��ޱ�⾥3����}_}L����V�fuܰ�-����sh�W%��^P�e�4��F��$5��.���-�M�'��qa�r]���t+Em
w�x����K��pyY��)���/"�ѣ&�������
3��o�feF�a��&\;��H�h���RND�V�V�}XÝ����wٍ]˱�N�Ě�>��Q�+"�\��(C�&]�|>%�m���s���2��Ѥp�4v�hu����"^����{A�����PR���d^��"{!=UѾ�ѳ� S���.�x��j�D��AP�w���5�G�8��c^K�Sr����LD�Ə�hN�k粲'G�M�mS���8�ğ���li��'ܙ$o�e�����j��T֋��	�=��h�����hw�$����o�^����=Z6�G��|����D�*�2���N��+0&^
�m�E�1��񽁮(Z��B��p�ئ}�ļs��z�k�F�}2�Y�5�#b�Ub��g7�6��^�&�JO������潈U�����+�����2��6�����"��C�~�;�3b�1:w˔��J�wҚ��Z)�VC���ft�;�$(D,��&�`�j*�:�b蠆2�ܨ^N�p�"��j��|>��g��AK(��U��>�d��(U����G�YL��r���[�}�0�;��O`���y�X�k�8�AVlVz�M-4��U\frɡ}P���l����M�~�%:�O�]{��2�����!��^K�:����~lt\��D�*��z���Y[��٦��1����|��ʹ7���V��Y���%�p$�Q.-��i�<�;�$&�ߌcv|�t���Z��\��Y��L�i� E!�A-�+$��M>�^��q�����l���=p�Х�!�y���o�zz�ɔL;0�4Vy��n�7쵂w��.�I&�����f�3�������K� �"�~N)kx\�x�[Sf��z�����_R�j��Cև2^�^vǤ�\O>ׯa5��Pf̘��>�T���O���w���Nxq0��T72�T:R/�W,vP�0�H�6����΄m�϶w�=�sʓ�z�ᣮ���G������?��́�LJ.9��f�+��[�ծǇ���˃��T�t��_��A�l�k��U��<�p�V�㪳�ߪeKO���ޏyi*�C�6)��0����gt���1eS��g>wf\r���X '� �]�j����ܵ�[揵w[-�a^��}�ג��d~��j���7�E[��B4N��2M��;T'�zאx8V���٣��=<0�W{7}��w~B	��r��n)�:e���4o�<G����Ϛŵ�1Z�|z{+�wKw�=�����T˰2�������nWbcۖ6!"��<崽2���,i�UuV��e眞ƳJ�D���*��I�J������=T9���z	P���M�k�״r�z�W�9���yM���+�����ZV�vM_
�v!&ǝ37�h�W�;������s<��`�[���	yn��k�0Q�v0�T)[��α��5�K6q�[�$�S+fIKυm�����'����߄f��jWKP��h3��ȡ���BVה�~��0��G8u(<�37�0�`d��X�o�y��	��\�G���6/pó�||{;'l�W���$���ؙ\�6Y��0�o��Qɕ���S.e#�>�x�T~��;O:ٙ[��ωm,F! �<u!���:�L�r���9�{��e�������+�`RZ�������Vg8T��[a]��]J�� Y���w''^�`e^�/���ږ46���C��[�ɞZX��X��{�Y�["��m�K����&w@�փ�Sb�k0H8E\Z�1>\�LݷL�YB����=^a���|�^����c�M<\v�y&��LƲ����ش�ڗT��g^���E����	��3;�]Ô�x����v!G���`���9Α�_˗�8߆��D/�"/�P�?rˌj�nx��j��[=���
>D����$4k5ĵ�^��x����9o�Vq��=�7�S��)[`M�'���=�ϥ[D��&��!���w���
�+���e��r�;�r�>L���t���z`�a�CF�P�nCOR�����Dc���]M�9ӫ�AU���!v�S\/������<o����;�rO��]�1�agR��C�curo���%|@���JT�\/�\L��nd2���^���tϫzj��׼�va�1xK__ �Y[�4�<ҏ��t��\2�����ǃ�"m�.�}ES��6�IҖ�rK�=:�(d�g7R�%�QDQAO�n�c�
#�u�t��n�z)�l�¨�<x�%7-���aΔ;�`;��3ju����¨���{�����l��x4k���)�uyN��x�y�yb�k��l7�L�(�-_=�K)�CN�ͦ'h�f~{�j����:�'P��76��t��/sw��}�r}���IB0O[��c}F�'�f�,Teg�p���Z�ڍ��Z��)���������"������ c3|�CS��x�|}�B����r��',x��Xu�q}�e���L�|/�W}�XD2����y��F�>f�G�A��!��iX��=,�o榜��]�Wc����|�# ��l���v�=ea��� �mU�#pV�qX�M^�e�#�KX��q�ݘ�+���	���N|�����wh�$X�+��(&e�6��`]��kGQ�o{3s*�h{d[�y�K�ޛ�}���X"j�h��;�}����]L��L�M)��;,�j{Lt�+�#�8��K�,J��0_�ޓC��m�
�:�/q��=w��j��=�x�y���{�h�O^���]43����L���֘a�G�\;��H��HcƟ��7󇈻�`���Y���b۪�w\��)5��<��?|"�g pS<"�g�u��=o���L�ڰ����2��/������&o�"_y2*��`����J�͹O3�̋��'������/�4u0�n��l�ļU��eM�=�g�_���P�GG���V�i�('8*޻�6��ٹ�h;�y�[d�AȮD���0ю���u-|.Ef�����/��.���A����B?p�J�������ֵ���>V�T��1�u'l8�z����3���Z7徰o˔���W=�����|������)�������7�CN3�}��P��ǕK��U�șu���z.���_<��g��i��~u	"Ù}�zJ�]}Bp�do��e��`[ꊐi/I���ge�Zm�!g�q��i�?v^��P�Ӏyǈ����X:W��y�GN�VY��6<t�[t�/�v�2�/-u��X)�%�@�֦}�l��b��/��w�L���O�H�{7Ջ�q�7CC݁1��/ES$�e����<�ϩ��r��K~Y���붧DՇ����~��	�\+

�n#��X�KG��}OW�7�D�W�11��;���v���[�W��Ca�{��ǹ
�9 |�%䡰��y�*��\�/>�r$Qױ�S�����7�1O��=c��n!�Ys�iy�X�a�� 3����,b���r��u�=t�����[�����^��;ÌJ�̤h:��t�	T]2�����ڸ
y\Yэ��fT>o�,i��	��,��������?�C{��nT��k���4�  p�BƒR��o<�ks�h씟�bb<s7t��;�n��z����vف�ݣơ���l�v��[2��fL2��7�CP�Y�=3xv�E�W��Yw\�Au���c4ͺ:fSvŖ���9ٛ[LJ=�6G�V`�x�|���s��ޚG
����t�m,�����Z8����j�^˳@B�}�I]O/^��r,6��TSU Lh�[P��A��[��쒷*Ѿ̻R��]��V��<�P��|�J�E\y��t4^E��8ۈq��L���g��8L����{�4�fs	��"��m �g*�]����샻�2Z�(�`fegcvA5䨜.F��ʘo1��z��$��>�;��]ѿ[�4�;��"���jԏ>Yc"��҃0�n��'�kc5:en���W+���KJ�;��0�����4�G� tݽ�bT��h���U��k����º��ֈ�` PJ��3o��g�����"���:������T�z��b��=�Sׂ��XvQ�9���ٜ�*-y�c�9ۘ�ͫ�1��R�G$8QW�gʝ)�� ��vK�iZ<�9�6�
B,��ՙ@�ܱ��`�����WI��ǔ�nV�7��*�o�:�mnm���;����Sh�2�ZfScN�3��p��@���������lXŦtY�,Rbݵ��5ɪ��䚠_IZ��s_Y(ԩ�b��c&��������V)�`�����f��w���aAw{�f�;�w+��,ހ&��Z�R�gGאn6x�
�[�ve_4� l򐫣�B�l�D�����Z�k4=;��/�sXhM���;�<�:;��^�#ә������$��rU7�c4���/p&�wCY+W7IF��t^1�	��L�F�'���Ի��{6� Mn�)���5ɭT��e㭘���)�͉�ث������^H�R�͹���'+���+5"�u���������O���:��(��eޚ��{��M��8q�[�-�$����!}����*K.��_Vi�tT�����v��cq�H����Je%Z�E�z�v��eR�_Dom��eu�|:�5�޲{����SOq��������w(��-6��+&u�ܼy5%�;U!�t��-kň=]�ֵ��"�m�"]qg�9�5ĨU���"����Q�J�ͻֵ��)8EI�6��4yXy��
pU�^ڌ0yIj�NJ���by7Һ9j��cZopvt�چ1b�7�Q�@��n����D�pFOr�*ou9�[�l��h�[�V��Sn9vI�υn�mT�W�v:�×>v�jQ z�n]!�ݰ�e�"
-���[��K8���VB"��dY��i��}��0�T��\y-���o���Ϧ�M�#�����D#�����U�yd���<�>�)�\�|}��t�����oS|��0�>D�-����5([ET��UcR��eR�4J�-�ڒ��JŢ)Z�J��Z�Z��"��iZRڵ�EJ�EUF#ZեAmF�*R�+jKj�ҫmJ%k(�-�QTm��جcXU�++%�UQ����QDAEU*X ��VUm�B�b���%��QV�h,V����T��Q�QE�ZJ( Ŷʕ��d�R#JTb����U��mEEX"���T-��B�AU�F�V�(--UYZ��b��DkQ��#F��e(�UdV��*��jT�RU�TUт��VF�j
�j�������U,A������",AmUDX«Qb�	Z�֥eU�TJ��-*��m�"�m��,E��D�%�X����*
��"�J,[J���s[_.k2�]
�1��b��|�����4HY���v�F1����l&�������G[��iU�9k�2�����,��}����'�"I�ż !A�y�Xy���3 �0k�A�*�ʘ��@��+Ӯ����t��lp��.xm�C�f�@=a.�����}�F�cK���ڝä���m\9��o:��7��ѵ�9؜�eCbe$��"���R���T�,������>��잭nt����R-,��v�Ϝ�G��%/+�uҶ�6���^Z//��[C��N��;�[s'4_k��z���fX����5ЍnS$؎����zא|���joRf�A�~㓫ym=�{KS�ظnV�~L鏪G�E���X#����xJ��i�r��_��� o��L�ii�q�;s>ܮ�ǆ午H�ty�i`����\�N��ȴUP���ĭvQ8`�H���g>K�	O/	�z����
s0h7���oҪ�3��wǻlߩ��\a�)����y�no�a�e:ү�B�T���	=�9o�A�y�4���h��gҧ^	��^��z_�e��6_°R�Ѷ}),qu
Ojvj3�*��kb�8�:�T��-���O�U�H�dw�h�U��'���-E�K��?*��m���J��%u	�H,��۹�Fq/�=���\/�Ju7��X8�Sf>l�+1����V�,�[�v��v� [DA�#n��LB�lS��w!�[+��\?���	������hui�M�X=/�v	���#5�KP�WKP��h3dm.����l�nx_�sh�C�;��O��J���l�e��4�����S��H��v�����3&zWf�/����Uap3����ܼ/��es�sVg���&9࣓+{��)���+�k����~�^�z���&��R��B� �������&��4���,I�=�Oz�h՗:cW"��K������G��3�j8!-~�|����6G�{�\j��Pk���KU��4(MC�����0����hQ�r�,�(7t�s�ZWN�wUh�XFo����s=]6��Gڠ=k*e��g�4t��%�^}&�g��Z<�as��vqf�{�ӗdX��n?_�|"畃�H�R(\*�%��Q0������Mzȸ�y�K�J9k�u`U�`HCY��G��s�F`ޘ)=�h�P�m�OR���ʛ�׬:�w/UA�p�����3��C��{)��y��]�f�c���]f��ǯS����j���|:nB��3f�F�;λayF�뺱�̓�I�*�ʴ4�='f��j��EnW�wa�i1��۹�ؼy���e]8��Ĝ�j)e��u&m�/p�K�W�$��E�S1Z�r��P9rS�4��*]t��������}U���*�[�������6�ώ��YɊ��X=��{n�g]���;ًSt��=�N��[�T�����SҼ��lg�-�d8�v��[O�F:�|C��6�+#����`���a|�{�τ�`IvG�;�������ڤ�^V��Qn�;Q�b14��&��zoz���X^:���,���s0��(w�q�ݩ�L쬴|X*,vs��%�(�l�8��h!�>���+G\>��i�c���<pM�;����iYR�ڛ����['Α�>^5��"�CH�*
-��:1L�L6���R���*-u�1���'�\q�g�]�0����iDo�ȰUP�UDm���+>�E5^y�@c��/5�;^v�:���.,��D����v�}�H�eqqg�2��vo��;;�G�C�Y�Ie��ݨc\rs�7���R��C�2Hn���(l.�^P�fJ��)D'>�x�{[��i8'����gpWL�ƤXt����<'�̓`��#�TJ�e���=��]_f��/g�ym��iϸ���	J����*
>��E�M��Ԯ~�P�C����y�
�,|M����Z9:�Y��Z���r|�Sz#��6��q�Q ���������=}������;�9Di���u��v��e�+�8<����{�Y����P�.R�=%�C������5Q�0�Z�L�w���
]-��7�\��$�2����~����E�+�
6��?��p&tJ�lZ׋&�~��Ŏ�ލ���!|>�W��5*�������_����H�]�
hP2l�!� ����tb�r��s.���l�H�Ф�>��~�;5V�ା�<<��׽�s<j������PPt��ە�.���P��X�"sP����*�+�N>�3�_�4Au/��-���u�i�}x���2�L&���$X~;�ª�c��3kƾkB�Yci����ue����g:��"�V;k���������6t�q�>�C�[Ҵ�vvQ��b��3&��<�s	eӒ��̧cVP�x_��@�-��K^:�/V5�#|�4���/�*�{��K�!�a�~	�'�K�	u=J�7ȵ��+�d'j��U�ٻ���x����f~�!�f���bX���O��| ���O�V���^�8�ޗ������}�([Ŋ-�3����d��~�]��MDZ7W�=�yFf��ٳ)�v�^�7�}50��[Nt��'A&�2�oh�;��ޮ������8���FK�C*q:ZT��uג��wi��\�}�U����_q���B`.[�њ�ʹ��uPK�H�WU�����e����@z��f����o��0>;��2N�n!���ƻ�L4:�ӻ�U��z��4�Y��U�I��3�����L�%�^S����d���{�σ�y�JZG�;�>w\�D"B�z�ݷ ��F�x�
�}j��j3*6��"Ü��3%<X�����]�5�����KӾd��(���&�_�������IR`�e^ �B�]��������znc�r7��yLg<�0�5ғI&GR�!��~_*}��5S+�x��4�@��}.��h�"�8�Z0IbrϾ�* ��}�|�c��K]3��j�s�9>��p�7OM����3���&a��l#�%/+yvw�$͎
y]J����[�=ӧ��M�>���x�=Yިt�O�.����ՇB4M�)�n:G��ʱ0�� �u��]Q�Qʆk��H7Q����
Ҟ��g7�qqV\���#�bz�t����Di]<�;㵥t%�cJT�%d�[a'N�����iJ�R7y��p;����Ս��S��G�q�ZgN��$|A�j���oz���	��-v	������y�X�J�[�f<9��4+bSV���JA�+,]���*�>�Ӻ�/5�v-��쏨�l�Ƒ:�#���ż%xdK��*��c=����֘���P�y�i{��)U��^3v;���6����%�<lr�˫�p�%�dK�<|3���B}�h�T��J{H��/ך{����f���>k˷� |�ˈ�yH!�Ƴ��UN���d���c����x=��#�����z����9O��w��0w�e�+qՊ^�2��_^��������ٝ����`�+ZG<�8�z\ ��'Q�3^��ʇ�*��o�O��Д���G��f�F�J��W�<NU�./��s���Y}�{K��T^?]�*,���7%z�1r�*��w�DsV.]��W<ii���l�a���Q�2��^݆K���t��}X�]E�Ϩ�t���u�&��J#`�0�A.�6�Ν���U��l�v���b�Q�{���2����n{��Glt��t�V*�� Y�4�����e�KH�z)���g��<�ǳ�U��r�W��S���LY��A��s�ZN�/q�⍺	��G���&�����M%�e������z�Δ�+'�1�r�L�5ܱO�����Sɫ;�A�l3V�\41#����Zw:򶲅�"O��rDF�,i�`�c������nbKX)XV�b�M��-�+kλ��n݌�!��i[��v����"��g,1��T˅�Ev��P��*K#�IerU]�����,noo�[z���~~SMp��޺0�P��*��p'��a���x8[z�Ax ۾}�8T�.���+�D�n����=5�[ޘ)[܍Y�"���৩oh��t�R�����GJ�f��������!�Y>��^qp���.�Oޔ5.��I�\�^���f��穳����ë>o	�{�p�0T�A~�aˋ���x{*k�}@_4 C���_��Nsvu�� s���sƁ��\ ��eוּ�u��1Vv+����k���[�Y���9��mC���-����]��<�2�z9���+�[�!Y6XG�c�6�������m�_0_"-Iy��AVx��"X�2��;҃�z;�ՠOu������9�7����},���K(�Z��а��WA�h���L���)��	r�����ce�n՞F��{��+�h�(Ȱ��^�c>�H��Mu*�G��X�X=0�l59CL�������7;��5�s�Qj�q��q�rUg��o_V��F[���ر.g���
s2e��<��o�3�u�I᭾�0H#qkۂwR3!Épy��zf��:�5Sˬ+�%�ù�ӥ��B՛G�P��'��Pi__�>"�{8S�g*�֛��_�̓P�?~4=��J��q!����Ih�i
�K_2���MG��۸�	j�zD�?(גׁ��͂�#��aݭV��b�\\YA3,c�,+�[pf�,qѩ�Szfw!\�[��k~..7�Ny�~�|׭z �BH��h�(���yg=P���Y����>����+R��p��G_�}0O���=<�	�^��τ:t"��������wV�7�62�ϵ${AB���t��%�C:K��g�x5S�7��.�5��cd��Gs�ӄ�[�M��6I(U�qu��|����^)5�:Lo�+"�]�^�O�<��D���X��zKY9���>3ZC����8V�G�YO/w�E��0RZ�x������S7i�ǳՏ(��� 9�tZђZ:e�C��V}5P!����?.�X�k��1Lk�ԗ�L��)��-=�T�భ��l��!����	]h����yT��W�i�2�@V{<v&����~�.ؗ���<c�d���$��̷�xGN��!<=~��j>v�
f��LU��s@��rr��ub��;��:����RAMňX2t�g��i�֯~��ꅇ�T�������]�[�g�-�ҝx��]��Hm�S#֎���+�*	'W3�h�/�Z%,���&�}��.�f�P��������\���-u���ƌg�951���/0O��Ћ�Uvr����[`�e��CI���ُ�Yx*�)CV��ȯ����ܶfS��O���=�[�=J8�sޮ|�;����j��o,:�	���3�Ixa.��S�5�.jbL�guے��Ϋ��t�Ly����^�u�	��Ϫ���J�Ϫ��YU\eJ'�_
��蚙Z�g�V����}�vN�Q�<�:���]�3cZ�m��Q>JD�Ql
U��s��L�:���۞�y�l�^�䎰��ޔL��w��	C�Ó�w,�hu�Di��$�}���s��r��M��zբ���v��r�=p�{�M[��+>ӥ�~U̿���}^&��Z�<^�s'���-�g�(s����8)���ʇ��"9�޳�=-�e������ߡ��8����{E��Y�v&�R$�#��Pq_ټ�<�3ڧ�I�_���A�9;���i�u�>��9?s��F�v[�l��C,�s�&��2:��ڢ��T�G{��S0�7قk�T����e�i]�!�7��6@J~��O;��?N��Y╱������Yw��#W��#W�G`z�ǯ�[*���C�Й,\\�[��Eݻ�����ԩ�}7r=F%�`@b=��Z�xu�{�a���p��n����-�{T1���ǋ����%��&
�(��C��^�[T<e�
-�}s}�w�<�>���z]$�0�2��$`;%/+���y޴�7�O.�������5�:G�}|�d�]�4/+=���ܦ-�TW>�M_΄h�d��4E��׵]�{�7.��R��}@��_s+��&��6M\4�pT��n(s���%j��%�n�WGv�����+���	Yb����2U%��*��!�۰���Lx�ӓ6]�Pg�Ŭwf�k�Ġ}뇻C���0�]����Kpȗ%������Z+�x�M<s�z�O��>��*n`ؘ�{���t�^��.��k�V=	�[�jt>��6��{�n�8w��u�Ϟ�,��n��N^���A��z{f���h�ţl�ʽS���u�ǐ���CU�RV�p&�:<�H�z\"�s�@�~�.3Z�L�y].B,+nw���I��7|�	^�,�=K�R��,���T3vY1䱦Oo�xƣT>:t����&�j��k�|��F��x����>�﹘ɩ�&_j}�]_oaO7hWd�(�\�s��Z��[lJ�̣X5Z���\(Y�gY)��wup���(me��kX��q���V�Q�Ҽw�o�K�	W�n��c�7+�{�Ogf1��}mnq�%p�]YW���X��������tvu���_�4��>
n�Ybe�dyX�������(pZ�v���˙Y.T�7�j�o!ts:>���l�x���!4֣��A��}�K�������7�dZf:K��(�ak+��mݍ�. ���*p�H]��K]�L�:}��'w ��A�/R�k�����/8��4�wn"'F��޵q�盶{�N kQqm��ʺX�ƺ�uz����>��o;�b���%A����u��:��[Yg�psk�C���ȴ&��n���E:��ͅY�"8&�����^pH���*���^fos��la	�>���ht�,u�]�*ꀗ�M��0��-2��U�2ɦ��n#��y��㹃$Zz�Eܒ)Fp���K�t�P�y񮛯�����]� ��V�Z�d�3jQ8�,�e�o��5Ӑ5��}����U�i����i�=`wo���:��9E��{L�Jɺn*渻��[y�RO+tՋ��d�{���������CC���:�Z��7P�����������r}��Z ����Ɋ+[[]3ltJ�|��-/�%�g���,�.�`��=gWP	�Q֫���I=(] �{��$�cT{8���!>zV�ۺ���n1������D�y|������y�ؤ�2B��]B��s���t��v3nnە��]��V�mM��Β<��t>���6���+����U� �%������JQړl�kr�hYIX��v�%���^7+��3л�\����u`Ȫ�8���*�{`���/�\���j�tI�ndiB��c7�)���Y皀Y���<�e5�P�I��(R�ĩ�y�,8_S�����]���Zڼ�d�U�2nP)`�tsۨ���ьV�x�u�T�\:�Чh:o5�.��{���+3�=�P���v2�,c���U���g;��ͤ�2��w�}��c85k�VQ>�J�F��i��z�+��cj_u-��,������2sic�U���mVQ�58��ÝA���՞�0����u���/'����,�ۛq���t�ZO�u�I�vkg�clI�
eє���q`����Uss��+@p/2��Zo&����%�\��i�{ڹfuw�ً�`�E�[��e���:�4Fa�jg�q	͛_n�D%S �y��Cz�{���NN�Y����k6n�.ҍ�#�9t����2��wg���r���:���y���q��Sx��k|ORz��O��>��X�J֕Y�"�D���hX�*���E���m�6�b1",m
�"��UBذ���TQ�Ԩ��UQ�D���E��TkUeU�M3QEDciX��m��J�b�[+"�)��X���Ub��,Z�U1DF"�2ة�b�����R�J�E+"�,F��Q+*1�\��0UD��-��+jZ�
*EQT��+`��X�*(,r�m(�J��(��F���V�@DE�dJ�Ubڰ�ł*�QDKV�b
 ��*�UH�c,DQA�DUH�ԷE��U��kE�����((���eZPTU�F�*�QX�5�!l*���m*PR�*ҌU�4h�e��j�V4��D�T��--����6[J�a��`��6�AZ�UX�D�R�m�DUJ
T�TE��*��l����X�j%j�¥e�FEm����x�oE\\�To�W� �M�I@�Ϸ���{�v�c��r�#�tt�
ĭ/��j�Y����q�]�=�^�N��Y�v����;�;�|N��	q�H�j�]��\񥚰�7�0�ld炎�)��~^�̯;^��6�̬u��y2��bY�ht� ��8��b�c�|B��M^h��ev��/#Ӗ>�!$��b��P�����<)��\�D�f5�PL�ƃ���ɞ�}���T������+�k�2�s�ܬ�ᒦ!F���邃��Z��-+�P��R��nٌ��ǳ˯�����9��w#��r�
�p����	BZ�s��b����_O8{-����cʼ[J/�}wǯ�~���I�`޺3>S.M�>G>Pè���w1��nי�wK��vClh��巷r!c�ݞ�G:df��K��j�4X&�*�8�6���:��f�8�cJIh�f�7���/���:��ν)x�;8�4綠���RvM%��â�<��{����0p�7��c��
��j��
�^����Ղ#*b��y���#'Z���>n��}���1�豭K��ӷ��Yk���m5�ǟ��m�=����:ʖ�p�Y����9�e1=K��W#Ct.�V�!��b��r�ĠQ�軹O�p�J͙����d�(�4[�ӆn��%�2i2,��l{�Y�H��p�T��V�
���:�f���wA6a��� �9[-5��}��"ǄL�G=���>���*���;�����ԯ	��VO���Kycq�]��k���{'Vf��P-!�o��
����Ln[39�w�,=C��ݩ�L�W�̯Lk{�ߘ���!�B|H�h��P��Z%�s��-f�f];��.P«۸.z�хL��s���������&L�Nގ�24:8��3�h��u!���V<��za0�������y���]5_�?Z�W[�N(g�	���hg��������F��t���앤���U<���_��G(�`d}�Ї��AC����v�Z�E�qqg�PN�Cs7�6:y�����]�ٽ4�^ŵ��'��Бiy9�ܮk-?�Aڱ"J������(T�Dr;k�$���Y��R��踞s�
�G]R�L8�k�OL�92��8s��ط��{�ν���A醱+��P�z�u�P�J���C�>S3ǙR׏��D�r�������;*�d����\�L"�"�z�r��dLCn��#��_#I��A�yO�zl<(�yʲ�ٿ�rފ�.�}6Zwח��8oN���e�А"�>jwv�0(���OwTv�u���4�-�|»WQ�=e�]�j9���\pO3w�$`�r��Lq�v�&�+k]ЋGl\ק+V�����hQb��%h���e_T��RV����m�k�ƠlU�0�̻0��C#�"�ˮ���f�/�z�Ypgk��_��`o���vHכ��J|�2*�L�(������w?R�:�h�g/���n��
��X�^��[��龽w�~;�֙��.���
ܰ����K
�O�z�#�v�GKbw�iTwjK����O=G�T�Vm��+Z��LG�C�_ϦV<�E��[ҽo,�bk>��z]�����&�y��ܐ�_�k���1�x�e��u�����׶��eym6:�����,٨W�N�Ȇ���b&`Li7���/ꎸ��l<v(6���b�����L򜹊��I>���]���(93����]�>�Xw�1��>ļ0��OR���U�M��^�J,�u�Ê�n�Ϛ>l��׮���ޯ��\��p�7��iZi`\q%����S����S3&�{��W=�*�0?Q=�y�'P��~[�3mzK<h�	3؂���,P�[�Kw#���h����s1k�>��g�T�9�P�Y�D�'y���5�'�X&l'k}���i�m��.t�6��
�rleU�⭵}x���[����P.и��}W�u4\E`6�P~�Y�_��Ӓ�i��b$�6�h'���m%s5X|zF��0��D�85h�W�)ګ�'�`��Y
wхYAX*�ѴU�au���or��U���t�G՛���Q��-}�h[����:�����ɷ��Vy�<��J�y��!��?k��+_���H�wh���)�P�����8)�����{�4�s���>�%�W}e�x��S��=�\�h�/�
+��<�3ڧ��4�?��G�����s�.

�b������*e#�&�}T��VC;@fŜ[1��Wۋ���\zS�^^�u[Y����x�mh�%��C�ҀY�}�W,vS<�l��i]�c�uL��0��S�-5�7��W�P�Ī`�H�6�����y޴�=:���b��N���t�Z�}mׂ��.׎��1`ޗEX}0���%��'Dx-L���uw�=�S��G��ܴ!PԬhq�m&V�
Ҟ�ઙ�G�����hߜx���Քp���ٺ��n��}��ȥn�p��-����ᒒ�~��)�L��L�#�|�����Ɉ0t�-�w_�S�T{}M)��g�e�<o��m��gY̖��zys��L�:��~TQ���"'�xj~���.:�a��SV�l�7���̆>Q�=��ݲ�?f7�tD�{��[�
YD�c*v^�Xͩ��3Z�������=�d-�qvv!<O�V�1��n'��NAE�)��7V��b�t�3MwS�(;v �X<��j�g�x����X��>X)���B�by�=�C�_��<||��Xe�±���H��E�2�!ݝw�A1~�K��9�L�����z�.�Ol���6X���䂧�CR�J�����9�m\��_�L��G �"X=.��5;զ�kY�ʇ��v��rr�wx���.B/o�:��T5�@x�&ZV��f�l�fJa���W��پc:����Wͣ7Y^j|��v��-5���i�X�v;>�x��XY�����k����^Z�>G�s����J�މƠ�S/&Z<eO4�<
���y �]1�>+��+��l�w���uH�M?�{����QOI[�����J%U3Ϩ&EN�8��1��q�7޷�x8�\�C昩���~]��!G.Tœa�hs�ZNq�>�gxp������άf��_�f��h�X[Q����Wlﾔ%�.T"ıB(P]�+�p��ɬ�� 
�`�/���z���A�k��Ta����Um�OQv���lz��X����grů7z�;�h�嗋7������ܦk)��������(
+h�����uK�9֌B�a<;LXz�iG�4:��� ���.V�9g�ňg*����r�F�Xf��z+u�؉��O1X��:�����PZV�ٻ��8X�`�МbE���܈y�^EÝu�.x��g�6�3��~Y��+7���g��SR�v����o������w:��s�h����)(o<�E���-s��jRF,/9ll�����T���Q^�U�Ê����G7NOp��X�}9�=C||C�(z}�1��J�\����{�p�����u�e�����צ�������\��e�v^��IvF��wC��c��8��cM��d�l�����u��K��;ȷh����T�(,��K�m�3��3�t��������y�+T����}�쬴|otյ�����ϫD��i��m�e�N�(}�t�T�C{�9pz���0x���e�z=)FF�G��K��Uh��P�\�K���fm�.B�R�o���'zT8�_4=��C۟L�x�+���x��xϒZ=)�+n^Z�����c'zx��겇���)��V2>�k���f}�Xd\�CmݭV��.+��<�\��X��o^J������45��q�j���X���r®{��X�n�&G��,r`�o�X�ë[F��#
R��m��";�}���;���R�,|9o�����fT�W(������o�x��#X���+���Iٽ�|���B.
�9鏝�����M�/>�a�O-ͭ2.9:�֋���k�4%��"D�v��_�����Tc�H.��-'^=��2�e4��t�ʹ��8{��k���*����ޮ�k5N�W<�צi�\@�3Q+��v}B��ιJ��]43�ƿ)���Tŧ��m1�N-]=ٜ�co�4dǣ'�l��s��H�iWaڽ���Rk3���j�a"������Z>��j���;beه>~4�p�f#�<ԧ���U��+��5�;�[漶|���Z�`�Zу�-6&]Á����H��l|7��➜�j�!6b�u�/<����ۄ�Q���[A�+ӄ�r���"8�D!�m��u�nk�X zha��r�y3}�m:��},��P�:]w��:�Z�n��M�6�A�ӥ�-i�jP�f�}J5>�u�ݗ�c�l��8�*�zm��ϫ]ze�w�~P��el؆	Y��O���i��U����|��̊��yڮ����z�9�w�Z�;Ó�ʁ��s�ymf�V�i[�j��F��\�sU�g1����������*�j�z�½}ի{�n���L,��Ɗ��	���[{-�ܜ�ne�bsP38r5�2oN\\���6/n�D�t�����-��U�P��1@o�%����o���v��k���VZ[JmT:����_
�M7ם��9�:8��+K��S�s2.��C>�=���Y��J�ʭ6�
��W�R�9��u��0tlꚀ�V}�F!'P��.[��fƵ�h;�T���"{�y�;�Ae�N�y�l��i���٘)܉	�҉��w��	C�ÀN5ܥ�;/�JO쬪���z�����KJ�'Zr�qy�Ӵ�
r�2��e�oռ��~�<s-���1�����ɬ�	�2����@����\�Aw]I�)����ï~Si�0�7g�L{;��T�$�o��o�>��s���0�<�$�#��PqX��a�3�Sc�2/{�o���c��I���� R��w��~X�L]�.2ށ���$�F�p͋h��Sz���o��s|�ݭ���i�����0?Ev<q�6�g�X��`�ne$����
�!�{+�^�)��G]g�����
	�I�,oK��桅��]�p9D�bJo��z�x��+Bp�%�:�l�i�2�Z<���{��J��BɫW�w(u*ɯ��[��j��dY+�^���x	=
*XW�F�x�����!ZV���LQ:{�h�Q��w+c��ɱ��5��4�T��o�c&�1曌gn�
�ʩ�Y��lŏ�`�� �J(sv�3@^V{���R����ɭt#D�$�$xX3�w�#}.c3��2/����!^2��Ʒ�I��i�)�
��G��7���-Ly��{�6�ܱ�4�s�g#>=�jX;D+v��Vط���^R\/Ҫ��/$�k�1��<�}��w��:���M�s���S;�,i��L:=�Z�]��U2�ߏ��mV�Yc��ju;7�mC��\��p�vI˱��i\�{��u��f���Cs�W�{�Q�}i���z��T�OY5pSh��Icn��)��<\�����=�z�בY����e<,ў�IJ�\��G�K��D��	Ď�1R%���S�@�~�/��k[��&k
�ږ/���{͝�VZ��źm`my	���|{�_B+Ys���&^Ka�(�w)Y]xxv����5$5���]��֚��\C���J�˝����7�л�k��۫V���I�>s��eoz��y2��bY�k�(���A.�]H<wu�*�qb�#��kY����ӏ@��Y��(�K�A�~�Dd��u �m��ѐ'��_P�:;���;���!�y��hVw{;B
v<���,R$ x����p3 ��ҹ���;�ek�X�U^`qq
2���@e`ygA}ݖ���3#��ᤛ��l�� .i#���˘;<4͇t��ΔJꙍ��[Pկ{VL�w@^�qJ�ࡏk�)�:җXt�+5{%LB�}r�,a�h�e&1������%|	{���Y?N!��;]1��Ev��%-��P��e�E9.��U�o����-�cӲ�B������{.����ޚ�g#�K�hxy������2�4K�{�6�ff�&��сC�o�����hK�]�t�-���~��\�o7ґ=�x!�a@�.ɞ�Z��e�0g͊z�����f�#�;�h�V��p�2�.]�_���[�L��c����;��>�����%�\�9��:�Y>:76�E��VL
������|2�vD�����Ki�a�^c/Fu�(�J�-�7<�4�5�	�Ǚ{�d<�I��ݵ}��'��iϖ�嫇J��8p?*���u����K�7<�2�G1����Z܎��mn��GrD1S]ݜݯ�2mA�`��%�]���w"��*��K�1�ļ�m�er*�0;E���Zn�x�X�%g�Y��.9yz|���̻�� )�0��A�qk̦pR��֫� eVJc CyЦ�2fog9�3`�nJ�|��\��K�@�k:]I԰n<�c��g@�x�i�K=�m�K�1e�GOx�i.��KUb�]���Cozu'�e)5wE`��l��c�6D�uxss��	Ρ`��"���
�n<r����e�s%�#5�|�Y�Բ�����	b6I���Y�r�,�Ā46�&h=(lȅ�q��Xa����o�6�;�����M� Kz�<�.K��w�߹sb�9&�wo��E���!�D���1(�KEu��V&�n㵙
S�J�2��cud�^��ѷ�Qt�`���շ�6��L�;q�8��ŝ�FY�o,�ړ��ݨ�N ���S��6_G��X�3e�5e�Se����n���<�1�.�"�54$3oL'�*���\xjFsc:,��gM�,��1R�Ք*�Ҝbk�l�٤�m���s渋���&eqwL�2֨~��4�Q�ω9�%`u��dmm���d��7`�ԛ�E�����*	��J/e��@=���d�+p�$%���5�4l�<0�95o�r����������<s^2�G���e��2�+�ݢX��z`��z��ps�"��j��J��u0*c�
Y�]k���ݖ���s>Q] ��Y�UO�}�yr��j�-��4歶hp�!Ҙ��|�s��WkQ��C�͆�`��j�Uf�c%����fF6�ȫ���5h��Wm&������$eqNқ�wQ5�Yd}�����V�.��n�ή�O$���nW2p������eu-�8J��֚MX�'<�K�=ˬ��]���^B�� <�>m�^�}�65s;�ڡ��۴������՛�;�-�j�n���5�`YO��+�U��@�.v�<�M��m�3[�.���v�s%wY�y�F��Z��F�`w3��Ӻڋ���e�;Ք�Q�X�1�Xx,�<��}׊�}�,���������Uy`�a�qֻ�qGAjR��D�K�[x�ӻi���cv��S�Ta�¾�ir���n�]�]j#i�j�<�X�3��%v��k�ܲ�,�Z�!�b@"x��㝉F-��9}�{��Q{;Kq}����PO6]	��+�#�ob��s�x���.�nê�,�d�p{�f,�N�Nf��}�A[�-�'iROi֌��P��m%�S<�/�޺ՈC,O!
�E�O�o4��u�kJ��j�4M�S�(�4���,�"�$��L��*�c�Xnþ�a������gi�	�x����o1r�N���fG�f�n�&���y���] m(u��9�ܐ����\N��2��t�J�%��,�R5��'&7lR歺m����c�������r�S��L�����{�4�#��������ύ��Z"*�*V�-D��m��h�֢���ūb%�EH��J�h�UDiEV*Dm,���D���)me���6����DUEEE�(�
�UQDUQ�Ԫ�,�`Z�D���F��*��J�IZ%QA�D�֊#�ՙJ+��ֱT�X��f\-�*�aQZ�Q"�*QU��TeJ�J4R�V"\�b0G`�\n32�ƫb�Q���Z,b�����cQU�J�j+"��DF1�ma�"e�\��h1`��D��e�L��5*�(�DDX��
��P�EU\h��Q��lb�)�������*��h�KmaUm))Y�Fʷ�*�,�֖��X娋1*9��Yb1i[m���(�E��\Ģ8%m�cimTX�F+iY�̨�1(�\����m�20��#\j5��T�0F�1U��nem�R�ё�30,Gh��̲����5Qc����c�P�cV�ĸ\��j-Bա\��Ue111D�kS9�,c�Q+I�S�e,X���TjF�ff	�[Lr��V��xfg�����j�1�6T^4�ѩ��&���J�;'��]���ۘ���ޔ��B'��n���5�w�j՝C�.�LMɸ��2W3;��.�FE�]�?H�4�<�KU�(�h���L���<�&��m��n�����.dK�gm+<�kV��E��럧�\,���k�f��*7T�e��]�y7��o	�eΨqԾhN(g�	��eq��Mq�$���Ŝ���Y�;���ֺֻ�^�:�����M[����K^0�Y��E�45�-^�u"������ًUA$�oM�o:��PP^.�;�2���1<�6�9��%�^�胵q&�!]O?u�����O1�������(S2�R��#IwVwEt�8�k�=38����D,i�WMc�-�5�A��Q+���B��ꔡ�It�Βƴ<J��n�J�n�g�eL�9$:��^�.�l��̓d�����N.�a�w+�lI�y�Nϲ��[���S�5V*���ɵ�G��CY��(���ϔ0�2�ß?D2:�,��i��X�%���:t�4_l!Z��h�K�5�hr�a��(��JG�f]��,S��O�̜h���(sfXǍ�Ѥ��DZ��{V�N 
���p�.o^j�#�L0�D�.�%][lnݶ��:��B�LF3��nAt���F�G�~�j>W�]mۉ�"��U��QVJ��e_>�H��z���滰��9��Y)����r�͛j��ޜ�mᚆ�g�*��1As���+�hVr|.��C��l�Pٕ�f�9<���v���P��U�o��fM<-}�<e��	��I�oJ�^x�Y�b)ȚYә�r֜�;�(�4h�R��mY㶤^�u�ݗ�`u�%ڜ�b�ajeK]��w)�{�n������lC�0&:%~2/:�p����P��b�M�՞ӌZΎ#���'[k�V��}���Yu��X�����LtK�C�\X�wηup��������|�G�$�q:�l�u�L�Ϻ|'�CY��=),� E�6�؂�xm�e�k�A~�h\�9Ș��:1_�:���]���mu@�#+s|ka��d�ڗb^Tz
U�r���ȑ���"d�;�ߥk�WoX����t�vHN��<8�,��0I�N
U��Ӵ�r��)�{e��{��Dv��z����Wz0^�+�r	BZ���ۻ@�<C�\�A{�֙�M��u����T�|%ڱ�nx}�!���xLٕ�{Z�R}��Q��4(���)��j�Q���j�]z�S�"n�Vj8��o	�ڏn�P�Z����9�Rշ�e�Jvm�R�-XrV��u�b�U�:^rG��뻓b��7(k����4��{`U��j�\º�u:�1���\����R�sd�����+޶re�4O4�?q}�
+��8�����.u�&}�&���w�,?d�5�)y��T/�E-m�L�}0T70�=i$��B[� ��z'U�͆o�	���8����A���S&Pá�6�`X��邡�2�W��hWH]�2{��w�̸F��ł�KEb7���;MaޕI3=>2탎Q#���R�"������=}�k�]��g���L��d�虍��k�|7O��f��]v�V1�v�^`����C����T��:����؝t��l�O��Y�~uy*��)�
��G���wh/=�S�W��:�^�}���=J:Do޿X�"���f&	��^4��V�ɮ�\x'�^��]w{.Çq�_U���,o,���w��5K�z�~�w/`w�H<CfS:�(�{��]�m���U���>ܮ"�nË>�3��P���C��)���^Rnw9�9�N��/OӹI��d��}9���.����G�NU���B]��`�]��oe�{��к�z�Z���!���l@P������ɫ5���ތ� `����&^�������z[�M�b�C��[�YiQ�~�A����X��&��4� ʁ6&�غ{��,��F��ێ��/��kFTF��չ�w���^�y��Q�¬R��F��K^��[�N$s�1R%����v	������C����I\�V�a��j	��`���XZh3�$�J�ʨ��J��C7e��e/�)�'l6�s��5q�[n�T����ƣR�=�K�x��M@I�$s\.]���*���z���������T��>>�;'����[ޯ	2�L�x�(��J"|�_^����uܣ�S�o߶9��\B+�~_�R����j{�{�T#+>���;)�I�(�c�w[h�4������N�y޲� p�|hu�<��:��1S/�r�W�J���Zߦ
��E�u�S���@�'�%u���{}�vu��g���YS.��؄���J�'����u��� E���Cx�K�댼p����\/9�^kCҨ�ҽ��4F�9��Ӣlz��b&>9�>�*���(O�WI��υ܈_��=�F2*�p�%��m�>ohR�~�fi�a�]�Ͻ̌e�8h�^!�Y�xm�}u��`a�RA�^:��y�-�ۂ�����hc���X��r ��7�Gp����lM�{rc/h�����@���Y���
*ԺӮi��v)L�w׵h=H4F"�\My�������'B)n�u�	[�I�zzS��+7�뿻���/���Jc�s��g���%�k�±�1��E��Y���ɏ�P���,_�ѹ�+&����A�,�&W�ng�:������ ����U�z��ZQ��~c���Y�g������Q�[N�+*��Zm���zdG�v^��]���q�=�շcd��^��A�ߟB����I�u�5jW�."�#���Ey¬�|t���n[39�w�w�����;ݽs�����v3�wu=ړ�p�G��WR�B�t9X����.�S-K�����>�v*�ַ��&�9K�P�:�<f����)FF�p/��U���U��e*���qCw\sV�X �m'�	f���59C�:��N4=��*���m&���ȼ|��3��n�a�D��7��R�+9��b����XdX�hk�Z��V�\�W(;��0�Fׁ�zgԨ��9��s��P�}��ȸ��9�̮k18��6���>��GG&9���W�һ�y�����]����̱�Җ1�#N'��}]3N3�0`�6���	��i���oMߦ�����=f1W�\�qЕ�U��q٢��cA�� �Q�w��wݎwr^���X����=�'.���Ƭz�������C>4u	�:�t���/Ufa�[ǜ�����r��
Զ%����j���G�P̿z�^�4��S�s5�ݓ�蹟�%
�T(��Ik��3��)C�zK���ƺ��6hsf��*����.[.{��;A�o�ɗ�����l��K��I�ׂ�>W��r*>v��Ϯ�פe���//A�0Qq\A���������o��"��xg��̗������^s=�ާ�U���Ys햚�ޘ)+ʄU�3."ׇIh�2��b�Y�q^Lyft�J��U{�`8l������<^��֡Ϸ��W�
ܰ���y�Kå[ɷc�D��9f���{O#�[��{�l�@^4��1�S��g���^4y�>�M_��H�̆���6t�>����=^�8&̮�5�	�&d^u��P�/����^�=W�ǃנ�ZsV4h[�x�S�����}2�����
�_��ΰ���R|.�%!~�7��5}��<���5X�-��N�-,�������e��V⨾��S*�Դ��.gE.y���17B��uQ`�C����|�[�����Ra��g���}L��+n�ON�Fr]���T9�ѮM���L�d^$݁���*W-�DLĐV�_^�Fl�˵]�t>Z��[�;;j�C�H�s����1³�7f���윆���;Z��)�kHYY�K=����,�h�w����]ٽ����k��I`�O�紸 �j��ы���L�z�c65� �A���!QM�B�>˕��oU��Y�e�\^\�/>�r$pl'��(�y'y���5�V����~�\��f��xhu�Di��P	lQ��Ӵ�}N\�৮�}�ɶ�|�^�c����	̏�ǡ��{���Sh�]�(���K��(P�ԙߩ������[�?m���/y�췵��)cH��?zτ�����d������Α&���Р�0`j�{�m��{��{�T������)y���~X$����22@�i)4��:���Ď׏�ӵ^s�*�"Y"�/�]��:�=}S&PîQ��$�9K
�ݚ�����Rm]<���Hz�V�vA�/v���VXޗIXj^.�."F�4ƞ���ߝfK�kt��ZjL�ܤ�:8)�㛢�3@^V{���R�ޗEX}0��6��zg��z��f��$�$r �L�^A��+|��I�Z|+J{G���dx}�2�ͮ�ؔ+�23���VlEÎ߅����NT���ٗ:e�m�1	ݖ$ꢔLD%�����tn��ͩӊ�=�l8��\����]������;��+�ΝN)�w��9�s�e�ж�v��\:���;���K��.� �m�ҧ�_F���8��,��=v��}�-��f�%��-��LҦe��#����gs���짉�}�cb� V�[ѡ]+^�S��ao��E�do�W��p�7��*�o�lw#��z������\Dm�q'.Ǵ	P��O;� u�l���V�wxA�۝{�E�Pm:�U�q`�J�vM�R#����N�f&�s<8��|��!�{����u�Q�.�`�ċG�y�..����jD���E���gr��u��.0O^���kՙ�f}!�jZ��VZ���u'b��w�c-+�Хߠ�͙s(����&�X��	���>5�&R=*��妠$��9��v9}�>��oӴ���{<n�`rç2�6�f��g{�h�ё���K!ݔZ6=ٽ��U��a���Q���ØT���qD#����[�P��.�4<�y�J��u����Y�R㚥ȫ�BZ��k�N�ּ*e��nVj��*br�LU��z4�E�ه�͋�t��:-�}�+
�(�q�ۡ�=P\����<9�ɊRY��E�5jI���+�1Ϫ$�E�9��x����A��<�ֶ�Gv�<�dGuαB�p��t�qL�:�ͭ�,�8��.Z��ig,c]��%,������*5�Ksx0�>�E^.�~kB��=�v3��6�J]3�Ev�ҫ�}qW���,�����+���r�l ���yj��K�'���z�E/5���J����秄7���S�C'�*���اȘa��TD6BX�]�t�-���<�ȃ9�j��h�c�&���S��67�)=�՞��L
z��4Qg9A�3+t]3�Kb��l��������|����4W����,+��Ȱ��:a:osn���ֳ�xE�z��{#���f���k�eq�m�1���P��_��7<�4�zW���ZaD��h�N�fk�}]�p�q�|~�������%��">��d�dn;��xU�p{<�7g4E�'[]��,p����?R�.�dyW�r+¬�pyiq,ܶ`A:ɜv�-�a��t�D�o:�����=�xVZ>7��WR�B�t9X��
�K����&x�]�'�9��g�m@�z����K8޿�_����C7�U��
T8����{Up��6��̗��ru�����	ٷƃ�,B��}y�p)]2>A����6�쳣���K�x:8�ҍ��s���N��L��)	��l�`�7siE՜	�($Q�+t%�40nѥ;�1�&	�
J�C�8��$~�=}6C��`<�!�^)]����~m4�-K����L&jr�K��{�c<g���G��a��%]-s,�J�7{f��{��*���uDK��(3qO/Db�#얽�0�Y�`�ȹf��c龾���o�������i�2,�fX���v���[�Z��Nw��O_5�WE�q���K���zL�:}�h�P]L��P�f&��1�#N&t�_d�w֑��/����=���rCǌ~��9��p�� ���J�.k��3�u�P示h{I*�����W��[V;����LZ|"��u� 8u ������q��/�c7�[�/bc����Jv��`p�ݵ�8kC������
��0��2�Á��4dv-�1M�E(��y�~uw��������Y�޵f��IXr�nf0\E�Z:ne�09c1g�Nr�*�t�x�cK���D�5��IP��{s��èu�w�R]�
ܰ��+�j^�Ƨn�:��|�n���Uy�j}�v�}���0uxi�yT�I�Z�<6�o\�4ՏmwL&��]��g��{��ݸ����m�~�yM�F9�Y�P������rXd>�ҖEպ�j�k��[��G�p�����ʍϏs^!>*}���_t�f�ҷ���>w�:Nd�;&iG���'Gs;�n��t� ��9絹CP@�HV�Ms2TN�|-X�5;��{����#�nw���j�-��X����˹ڥ�w=3\���7�Kpp\)*��°Cϵ��[�`�\x%.�z��R���P4AkB�sR!a��V��`�(���zmV��<��	��Pn���"P����̢	5��+��Su��8(��aӢon^`�$ĵ��Y�Q��b� ��ߴ���}[��S�1��'h)T|7����62�q�ڲ]5}2�u���Q�c�Ыc3�`��ܬ��w����)69��_�k���1�pYь:��e;��c�H𳦻4$����ӻ��vž�{Fc%��j�d�{�WFr�_v]����(j)���'.����dm�w(;��u������+똨�}=K��V�u+AQ�S���[��X�FE�{Nl:탸,�j�8u�0��c?@5PYX4%�t+G�G�����}i�sp\Kst��Jt�O�����G#j�hϵcG����������ɭ��*�i|����=b��9*��aЇv+�¯�;Kphҷs�����Ƅ�J�I���@[��Go�@�헫Js�'���*�l�7��9��˕�Vu��v�M��ƴ��:�n��sr�(GLgN��qx���}��\�bE,�2�&������Tv�e��K�F�i{IrՆ%i;�.�g�5�<�1�<���fb7i��bRY���WYj5D�m�)�Ϋ�����w8�Q��j��ɤiR��7��u�*ĭhr��W����[�e��T��1Asd#��Y.�Gu�:'M�w�)m\u��iP�%*�o�(�ʊVQ�ͨ]�iQʰ��7�~�}Ԛ˗.�d����e���"
��m�G����,֑��N���`1`���#��;f��=[4v^�Q�j���']fO��ޥg���ТM澱X��wʷ"$�t�+P�bT��>T��wp�T� �@�m��K�s��9ܣ�pM�΢�n���
�}�h��<N�J��A滜�FR�͚�]X�}'nb�|Wv�r�9�xTE%݇)�:}Ӥ�,ʜ{��O2��w�o���l����|��U�
�f�]�)@�8���*5Hw2ժ;x�c��D�m^mnp��(].x�%L����ՙ�t-s���2.���i��~G{�U	�
	x�̢��_�CP���^�'�*<z+9iB��t�[�Ԫ�	���^�A�) Z���/Uʼ�۠m���9*�^u��Cx��۔ܡk�b�c��+��W�c��K�&�wQ����B8w���k�YI�~5��?{�Ks���&��A	fTs0�%h̴+��e*hT�E
���⣃A\��*V�1�Ō��a����[cˆKYW�r��2¶7-��pQj�m�,r�DE�T�1�X�VEUL�Lq�e�m�m�-K��Fq��-̈".%R�++m�`�*,F���af!F#�W-m3(��sb�Rص���R�TW1b#��clLmj��SV�-�+�U[h��LLh�\eť31LE���2ыZ6�h�%�s2�D�U+�Zܶ�p�Dmm�%2�-Ab̥�؊���2����ċl�!Z�b��)m��T�b(Ŵ�.d2�`�r�r�ڦR�#X��Q��B��b4�3��j��Z�B֊EE+ER-��q������f
�K[ElUKm��*\�`�Rb)m�֑F�5�b�fS9me��+EV��Q+P�*"��+����#"��h�%*)\E��h�Ɉ��"��������l *��h�\V�Y1�;��P�'Q"VM��k1��_���C���u�@�mEU�Dz�5�'UΌ�:Fv�q������]��U;��pb�R��R�4�|x��U��GyL׉�r�Ro;;���Zh���Z3�E��U=���g��6��/=����2�=��]3�c���;��]�a�m1�rىԵ�5Փ]�7�/O�L5�b�&:RXϭ1����-�*]�{�;c8��*����b�)���fC��oW��u����ʳxEy�*���x���Ԕ�x�|��$�<�����	������F!&�p-���3cZ�?o�+L��ϥ�vnH��r>����+���J��.��w"G`Bb�(�y'y�ZƷMU���S^i�!���C�Qh%�0IئҮ/.��pS�5yO\#���uו+ښz?W���ɟ9��Yy��(;V&R;`6��WP��J�R���G���Z�N�ò?	���w'�@z�סKC��,̕ر�q��K2a�y�I�G֞���mP���4�4hZ�����{TRX�aK� ���%L]~290/U�v<P߱:L�k�݊F����W��)S��.�ᐫ�N;Z1���Ƕ�	��}�3T��6Al>W�� P�g�t��K[������6�����:�ѫ� �j@��S��H���
��P5��R�j� FP.ɣ�\=h����7ֶ3��4;����ǕZM/�P���h�Y��k��g�A�� ����aߜ�kD�&��u\l�/rw����e�X��C���/�`�\EX�dm/E#����oK��5/�`��l���G�_��ߏ���a"��VF��m�|mYk�E�\8���[���o�d+��z�wE����W���\}7��$�t���X�޵��{=�W->S��𐗚����^��WեG����%��O��_-[^�U�w�10@�>���JN�f%ǙK��Ö�^�ω�oD���gFş��)�����v�cO:a�K�o^��LK��5���r��y(1�7�>̀�nWm�qe9�7�T-+�ܴ?m��|r�Vz��7��=�#>�e�����-X�����������fw�����-�/Y�mӨb[���]]���c|��'���t�x�"��J��]�J�tь���լ���s�T�mzv���r�\yl�PNX��W���4&T<�� t��ړb������e�o��}*��-��G�Ż�V��[Ag�̖��5��(a���y��P���)etH�k���_
��l%����@\]��;�ou�α,`�;��KMd3s�ߕ�݀�K_j[}�Nw^k����r�o�����=��;m�E�EtO3����w��u<�8��^�F�e#���G�Ҡ>�.!�DsG�Sm��O8��sZ����+ݍ,��7e����[ީg��ё�����G�{]��o�Y���n��+�|���^q��A,�A�v��u枮3Ps��ؽ��X.`�Y��L���8��w��<�?y�-�9K�X\dX(&E_������íxT���ܬ�ᒦ!E���427^f龦28��֧�	s-�"��P�˸z��yԎ���kL�\~�2�N��vp�~w�=��n���B[�I
�Y�J�-s��5�^��\3�擮l�*g�J�<��O&�Q��LL�}[D�pS�L0�$D,<&��»����m�܈E_H����/97�/���wg]爥or5g��7�pSԣ�}�+4Y�4�k�!�X�����{]��{z���4�x���=�t�ޖ9,��=���>[�	�csnV�nOX���T�]+Pm��-0�z�L�_���Z�J�,>���Ɩ�^k�ev�wx�j���C�ب����h�v�}��^�!�ⱪ�%�gG���ɱ��vdh�c�͐O��;y^!=���蓭R\��V��u'��[�����N���b�:��;�
�W�1R	)���Y/�2��uq�V%љG��޾�(��!,Y���t5�-c���Z%�M��r��k�}�[X=�:�<��w7U뷛~��X�d�os�ۘ�oҕ�щQ~��8�F;Dx�jDw�"����I�a�{�.�w8���}N�;�:Xz�z;�բ{�WH��M\X)m�Z�����}�w½0�������v��3L��l3/�w9C�Rŉ^�v2����FF�p/D�� 1;�T��������d�	�R��B4Ұ<��}��mNP���C�N4=�3グ�w�9�ܶ��5X:I�U^���W��eUB�";���A��yz#��v�0�Y�Pd_��e����6���;ƇuR�>]H�`�2$2�QlS�������"㓝���7Bߓ~��S�/{v�<L�K�!�v�����@O&^�B���Җ1�#N|�^�1�0b{V��18�O�9}m��~�^&^{��x�:�-f�V)s]�)���r�.�[��i�JU�zӮzo�z���ƿ3<{�����(o��2���K6l��\R..�SnX��z�4�`e1�J4�x�z�ܫ�8�>��b��i]������㽃]�Za���Ӿ�+P��� �׵�vZ�tj�j7=�>�n̰�ҒB��#v�_k8lK�Zjj�(!��m1#�7���ov�f��ݻ�iti�CSS����%\�د;wb�Ǉ(hh�&6x'��:Ll9Y~������;beه�"�o{��,�5܃x��)x�E�x�d�^#��^t�m���=�8�q�8	->��V{{����b������y<D�!�9ҡ����6�/z]%c\�,0|�^nf{��uW�UH1���Q�<�n]Á���Ϻ��i��&8*r߬�ى�jǂ�Zu�aU#�g��'o̚��E��zW������ּ�$sU�Kp�^<vԊ�-��Q���to<�0�����^;Cv��.�eym6�;�rݟ���㘼	��m1��Bok�v�j��ݕ�@�]�8Y�Pgۖ�N����^�y�Vy�y�ބ�?f"kT�"��;�#��T��U��x�
� 7�E���+w3!=)�B�>�=��oEN�WWc����;�f����E����UUqu(�_
��:�l���d�?g ���5���� ��/��t�@oP�՟%�X+���J���v^S�;DLl�P�wk쳝\Om���+��Z��V\.k̲�a�˨k�ZkE{�nm#�z6�2�Q3z8�:��&F����ln*�.�[5j���V�����u*`�u��Ɣf�)����_o�[n'[Β:���R�Li�Uh�j��u��e�E�^�6��ν�W����u�v��hqDi'�`�Kb�J��N�9N\՚{���+��us�����߼G�rɡs׼���<��JՉ��ۻ@��0I�P���w�:ڹ��I���}�^�3��_&g��z�׿)cH����Y�)��=l�OY0��@s�I:�=�]��f�snv��]@�Ռ�X�L��`T�5���~*�T��r��`�_*�ޣ���OJ�p��l�0OR�W�V��X3��q~�5��=��t��x�mo�cd���;��t�rac��j|&
�`<��s�_�T�"�������v�ý*�桅��xv��r?[{��{.y�?$�G��Η���>�5ᱎ��m&��D��Z�t;��<B�{ׅS�η�EO��&�q�Hi�l�[ʱ0�� �o��T[��{�c�"Yd�Na���#+<����8��}p>q�=񘞥����v��Vط�����[t#W�|��{��Tv���P��ۘ!�]j7,z! ^;�-����},i�r�a�r�s���5����&�����FP|(b��jʸL��m^)� 1�sަ��]$��yD��	���w�=��IR�d�)�T���sj��Tޖ�g;Rd�ftٗ�^���'6�ݎ�Z[�� ��Jg��FWZPXu��-�o� +��.���*:!�� �/fs�U3�^:�]�xnW�,�`�J��dwr{.ǝ�	����U�i���VY��O��П'0="9�|a'6陔����$�ﮟ�8��z�Mi�Up���y?���J��)��jg�/�����	Ď0�K����ʰ���~�L-�"	^�'�u��ֵ�eC��rJ�I�*��U˰�̘f�W��)r�^�U��M�3%0�{}��S����.��`-5���{������L�k�:ۗ�Gb����Zl�=�d�Nx(��ݵ~�.=y���=��v�e����X��=<6>A�n�,��+ƪ��q�����S��˘;;�g���<��o�L�������J�S1�#���v����N�ֽ�L�ܫ�k4�~�ZI�g�w!Y~��B�e7t��Αi_��x.���ay֎�Q��R��/��n�s�=��e����gˋ�˕��yi!_k5�_�댺�{~�� �V����#i�7s�ޠ��;W`+��J�����@�VϺ�i����"�g>�E]�s�,N�`v���e1���K�q��hN�d�s~����]�*R�x��۽D��r��e�(�K���\�������׼H`�~���y�)�/z��E☡p�h��D�ϧ�U
�u�^m-��ӌY��̫򷖞���9��5�$��=E�_�X�޷��2�Â����:h��r8�zAk����>�J>{v��5^��W ���j�<�[Ξ!�oK�k�°�c�+�b{nժ�m�`�Ѿҋ1.��_���ɜ< �5�(/�^�}qpu�����ؠ=�{A�1�S��K���x��p���z��C���{�2�������-�T�X���:��-�����7VUj��^�ֶz�i���rw�W���+-�۲��B��'��0����n�����d����Nf��a���wTͨu�Z>6���
[h�/e�+�/2����s�blP"cנ�i�1`���r��u,x������|Z�G�ҡ���zF�f�gv�����^�y�m\�CH�\(;\�J�������:��	��}3�o���/$W1��FOP��`~�.D��4]Qu��Y�g"����Y\��<� ��~�#�)ܯBU|���4�[;�N�G��>�ZVs��T7�\T�Ӵ9{H��:v�/���y\�A��Z�ɍ� ��T���w����N:Vp�հ"���UA\^��	�	��5���`��h�s���{[F땋6���"��ܹ�ƹ��LQ١��ݭV����+��̼we�;�g�年$Zp���q������S|�����\�ؼ.��H�.�:y(�S-�߲�R��#M����yc�=�Q�oo��צ�a��<�8���X�k5�\�`)��>�uI�s�]�w��jN�7ut��mSC[��fx���Tŧ�(o�Ϧ\;2�v�n����`��z3��(7{1��.�j�9\��l��`�0Q��dA�T��
�����]�Hܭyt�+џf����g#�
�����jS���g5a~z�Y�z`���*V�c�Z𕞝\=j;�ںl����c˽87Ԭ�Hŏ&�xg��%�ϵV��3|�7�X]`��>�h���E�cv0�z,&����#~�>���4��eZV��&o�}��
��ob+�wwe�)Y����қU�N݊���c��3k�5�	wz���o t��{�w_���^���5K<��K�ǻ/L�P�Ӄ�2,�/-���V�0�4����^�n���W;ޤ�{�)􇻺ru��h�����ZB8WP�[u�.�d���z1��#�ĥ	����ܠ\:���5ϝ�W��^��c*d@�.��2�d|6m�a�w1&�̧�p)L.�|�#kA��"�`������J�v�ݜ�ˡ�)����J���qB��_[|�@�-���b��\OV	���^�x�~�}m0n�z�0�Q�7*��$Υ��
�΢�I�����|�[�0��Xݬ��g���^	��	V����*��^"�D�>1%����{K�	��x:1	:�&�m�^Z6״�O>����)�CcZ�m��U���_��]V^}J��.��w"G �(O,��|�r{�S���StM��C~�5��]�&j��A.I�N�4
U��Ӵϰ�ud�-�_�����|�cv|�t��������_�X��\��Dc�lФ8�%�C^]�Q�C�{�p>��;d���IsW��ì�#�s��g��ߖzz�̞�a�0�%ӗi�6:����\ລ���_�
���q�<��(�L���~P�,��.�}�!¶��S�z]c�z�W88@�#~�o��!T��Vgk6,��5�k0uz,��L��~�&{�j����>X����t;TCs)%])傥qU3Gmz)��5�7��D��(��{6ߗُTK�Ee���t��������"��erٗ�7h����Uf��C���>K��NS�WB��S����
cj��+��%�+7[����ug6����}�eM2�L�˛�2f���ܷ�}��h�4]ͩS��7�BW>]�U�$Av-�������B��>�6�#e�ҥ�2GL����C�[�r�#�4'��7_�|q�P�R�[���f���w]��Z�{F���x�*Vg_o\U$ ��ck�̳�
��K����W{����&q�)v����l���r�q�+��s���&T߀��==j���V08`�:�h��E 7f*��u[�7�+��T@��\�{֮�K[����4p�� WL}P���%�`"m: f������WgD�]+�dꛐ�7��ʫ@�@�l5�f�]\�����m�6��ІÈ\��.�r�Z�.�?�4D�{3N;i�%n���ژ����-�(L�B����/9L<l۸�j�λE^�
�#�ޭ���`S��m���#��ݑ� �h�sL�R<�A)V.�9Z�'��6�>�s�騸��-�6�5,	[G�:_mw	��.JԯNQ�B��6&�\����&� ;1ӊ�ޟ
Z�˝�����}�O��Þ�������lT�w�w7��]vr�V�b[N�f���aǘ�i?5A2�L(]s'̋��.�y-�I�,>����y��)�;�>⊚6[{��2��C�Y¹�ޘqQr��NVg���ze��P�|6rXݙ�(��cT���P�762:Ȯ���O�J*{���o2rtjky�A.���bb�9�*������:J�:�R�3v����/��Ov�:�g+3:��{��T��D,vy/�k�ï(ςc����4#��_:Nɸ_|YŜ~�[�Ȯ�:�N����+����Ύ0��y!��~^r�w�ȟ��C�c����[��^�
c���"��������O+��ѝn�ܮh&��` �M;��f�����Ef�4�z/�U�#�R�����y���l.9�}%6�0���0d41���;nmX����IՐ}`ټ�ͬ�r58�Y�(�4�cU�wh��M�)�15������-�fc纇]<���/UgZ�ܻ�ma���Z���[��wV�������6;m���U�H�ud���*�|�Y����Awu�u�ISڝ�}�	rp�阅�{�|��w�e8��	��)`ɭ��1�P#Fw����n���Э*���th[���_F_r�kk/8T�"�+Z=��/��r��
kA��D�j�L�bv�I:/[�FX��Թ$�{�e�����s^�B�y���9\�2���c��� �;
�l�����3�*��s�]�iF,�ک:�`����f��Ӈp�
�[�~���hO9U�֜&�.K�"�f�`:Y��_48�݃����¢����T�V"�85-�1��"6���#��fQS-�,�D���.�[B��T-��G-��Ɋ�&5dX*#T���E��f�����D1�m�R�"�LIX���l���!�*�s`�UZZ[@P\�0\j�lYUYZԭ,
��aYX�1�D�q&&2�R�b+UQDT�Yb��X(��c-�)kj�)Z���Z1�U�kZ��q
0X�2��ڪ�r�G
�H�ʕ�Ŏ6)Y1��̤���h�*���*�Q�,Ƣ��塔2�Le��L�ee�V���X%V��PY�khV&P��	J�q�WQAm�-�fa�AF��`e�B�B�*���3r��Kj#��ƪ���qp�1b��
"��-Yr�B����Qq̬�*,b��0eQU��x9�����p�ݟ[m�+R�7���^����7�\쭬8��eq�_�5��IXDR�ݦ�Bl.�z�o*�*����~�xh�uL��#�Ȗ/WF��$�mYk�E��u�8����󠈫��p�N�)��j�7�E>�Mjf4M�i�n:G�ʱ0w�y�+|�\���:$6��Ԫ~͒�zo�[N��w�����Zq8�����yǈ�3�e{���n�%Vط\��d.��__>��9�~�.ҭ�4��y%pXu����=��)�ޞ�{�%�T�qX��Uɗ��6m0�����Uv�ʦu,��2���=T:%��y�y/\����	�=�+����y=�7J��K��V=\�U9��{K�"�h��n����,oz���v_���N��᷌������IL��HEA�̺8��)�B�S��0��<HQo��tg�#��¶ҟ7l�u;�.����]2��+-rJ�:�E�j�u4A������{��e�"��y�fo�a2�X�|��j�|j5�L�zĻG��5���pX���g��:���TH��[�sƖ�,�pل�y9ࣟL��W��S/>-'5��5�]9:��x0wKN��Sڞٛ�<��í��^t���N�&��+W����)�x���Bf����>����tMN]do����\��opuNai�Pek�U�N��{v���[��>Q�ae�9������˩����鸮&qo>&}%/#`�a �/�u �Kh_�!�Pz
�)����G�NV�P�b��7��=�MA0�6:�C�(���cX(&E_�\zm`N��/}O/�ל<<��`��!M�d�9�b��z����LR�C�@�:E�b�B� o�]^�#�D����G(*Ўx���:�Ξ-�ڥL�z�}�C-p8.T"��(Kyi!CY�J��x.��t�^�5������Jv��+l	��1LP�U�N|����TD.�C�VD����F�z�qwr�;���j�׍p鑘7�
V�jȔ�:৩GH�B�E�Nfg:�{zW<b�����,�k�u��W����Qs�Q-pP\�c,�pI�.�O!�{���m���Uy�Y��[8�X��銡���L��nd3~ξ��G�X�s'm�f����֚��.ՍjP��L~-b5��-��X���*���:��2s�Z9G
▐<�{C���K�7 �[e��|�OV�Ϧu֭:�Ev#ʮ�Iy���g����������u��4!9�^M#�; Z�vкs�E0�\gݓ�L��x9�r��*�mf�<���R�RS���9#�_G.�d�R�g]J<]��d��u��:u�a�ٺ��d$A�*Ĺm�/X�����\��c���鳾�
��ƙm,�r٘)�þ����g���Z�C�*�7�'�>G�W��JM����:���W������kh38S��|�X���kV��Xt\��>w�/Ԓ|����|ͥ���w�J:1E�za0�jr� u/��q��ְ��t�ƅ�н�lc��xϫx�[J#�E�U�e�˩����M^(�yd���Tᛞ���F�­8��f����j��R,Y\\YA3,c��5���Qw��Z���-,OǃB�}���7s���q�b��jD�H�j�6��y�
fX�iK������6n^���Y�tG���S��Q�:}����z�,��TH��"�V�;�է���2녿W���J���C���=�b�衾G&\;2�gA�H#r�+������,>�y)�\�EQ�1�V`����;;���|"�z�g��^w%�/r{��]{g��it{V�4�Ș��;.�Zf�_���Qf��Iw�T"���=i�3�,����3�6(N�"�����@�8���^-C�jJ�J¯8l{���9:�pKo:�\��5@:���&L�7ζ����늢�[=�i짶�h�'��u�:8�%�$wkt�v%ݶq� �{��:�GTqU|⧖���wW��Hi����E��L���8��KGM�]ÏԼ�"E�|Y���K�˼�;5V��>��D�����e��^jk�:~�AO��k�[ҏ+�p�&eV�/:<�\LpT�Yᨗ�ɏ|�elqu��/�vS�����6�o��ۜ�?v83kƚЄ�X�Kf9���Iw�����,����|�5M7��T:��=yj�zh�㔐|�}4��w�|�c�3��^�^����-{����}�8��]�G�]q����Փ]�7�L�>=���/��oz��{6�^��Ct4=]�1�,g�%�	u<(P�9ȵS!�a�̇�t���w���h����>�'����{#p
a��g�RX�KG�?0S�^ H.��E�~u���Jy�$�܆�<����sWo͛�h4�Չy)
��qyr켧r$Y܏e4��<������螰1����ß=59g�tP�
��z������.h���q*'
��'����
��o�_P��]%�?m��߯yYy��(;W2��wh@!��#�-p�|s,Q�K�09N�ג�[�-
9�wv�����`,ۂ�n�-é�ҡR\�u�c��jh^B������
����߈�b�g>��Ţ�CSpJ(�������.h��(U��,�O��=��{�2oBzm��T�"�.s���&��P��e��s�n�2��aKE�9��|'��,�re�پ�\�=��y٬1l�c��4�!H�8�o��i���-{^:&��nE�Ap�s\z��WK畳v�{��ŗa3�H�:M$�K�3�3b��Թ_m.,����c<��J�V�w���=�03�kG4�ft�玔p>�L�c���מ�'���c��^>�=F�ӆ��p��t��K<%S\�G�����a��x;֒f�৕����T�v�}�w���{�et�f���֑��������j�1�o�2M��X*��޵��S�ٓl*��]|���-��۫���mM��L�����h�����,���յ����$�>w���2w]�֍8
�=KO�iL��U�!Or����:|�4����p�j�;�j����<ɒD��x�l{Եr]��UC�dP��f@}�\DT:.�3�a3�H�=I��W��B^7g����O=Zw�aY��c��.X��Oi{�O���e[=r�1���ד/̝����Wz�ͫ�JK_<��O��b�f)�=Ƴ��o,!��";�n�X��i�t�V��\ژ!1�_d����"YO��}1^��o����ѻ]Ԥ]4v���}gR��N꩕��(��R���8gH�s�]gFfR�p�����ׂx5-�8�ɉ�;�VZ�8�j���SK�)���]۾�aO^���7ݡ�$_��JK�[��'������{����Yk����f�I�ѵ��TB��&%�>�ۮ�^�G_���f�f/�4É���ƣY2��l�d��66^U�ծ����I�\K�q$6����+�4�j���l�a���Qɕ����
e�[��i@AZ�v��Q�7֏��>�>+�$��0Wmd��P�\9������E�Gi^:z�R�j�w7z��R�	��P�wH�J$�1��d_���yC���yv�P;��v��3��^~l�guf�jZj)jL�����:E�t�y��=~��w�1��{�t��=]4��9�>;��yp�j��(e�ʄ\�B_�夅k5�X�\eݣ3oJ���� ��=^��jb�i�)�˘��SD낟#�(aەDCo	�8Ý�/x���ص�]�R��^]������h�L���0R�����Lr�a3�s# �S�����Q��f[`Kp*�'���1��SV2���,C�Ś������F����*`LAJ����T�`����=K���\z�l������r��Ȧsk\�X����K�ni�=p�vP�{ٳhb@�$�.ڼ{\:���I�ǻ ��uP \��C:��j��Sj�_�nY@��L�{�=�t���%�బ=��ï��&��3���uoe���w�۽���O�=P_��xe��^7���_�{%�/;Iu�h�ir��D=����7��=+�rBb��76���m ������cҮ>�������]�Q'&	;�_?�2e�����q�3��|�OV��3��iԪ.������c5�<Y}�;���W�A��q���>������uh��w]���U{E��=�|����ޑ��4П-��eh���4�X�fX�s�>�ҳ�5[Z�_ʞݐ������t��d��<`Ƽ{V�x)P�.��ֹ���:1E��L,�P�Υ�C�]�t�W��[܊�V^���3��<�,�+��҈�+��%�h��:������E5{e�Ug�7��Sky���M����C�ř�XdJ(o��Z�.�X�����	�����a�LD������Թ��e��ݠό���7��5�^0�W"P�_\��S/>)���`ˤ{y���;B<�!4�]��*̍'
s��[qu�ʠG;1mɹB�L1�b��s!㬵�Ce���<����i�d��F�jKCN5��{Xw+�%@����J���Uۦ��O`��2]��P���Z�b��wv������촞g6���M�q3�2�ﾮ���՟�3�L�hX!���TKq���Mv�R7`��nNՙʚ�B�y*R��%�C����=��LZ}7�˨}�OY,��Y
�a�<)�wםM��0q�C���)8������^�I���`�9Y~�+����Vxe�����"G�fwo&��˳��H�+ah��4��]�:뵟3})nT"�V܈�J7=��Oϳ�7F-���.���^S>�$a�͜�P���nx�C�B��ƺySZ�~ҫu���)'��+�j^��W�w�����xi�U.&8tP/�gdNo�dg|�����׍C�p}0��;��}��/v8�ͯ�Є�X�u�w`�����:��"�W�,�s��u� ����x�OX�]����(�N�y�OA'��6�YF��OVg��j�2�"����A�rٙ�;����5�#ڝ>��^x��y;�UM�3熼lz��m4�Ԯ8_
΢�X)��s2�)�ĝ^����躛�h��{��St����u������	ˌ��v�_������2�~OQX�nY�>�^L���3]��2�g��o��nuV��*h�3�)h��J�oU�Y�c��eKn�io&HV$2ͩ�fR�3��inJ�ޣ�d���%_.�&=ï�:�r�+'Ԙp=�Y�T��RKG��Y7�BO������|hє�w����)�^�L�z�3Cܙ���T�&���Z��H�>~lw]��YV-�ە<�R�f�qP�A��}���ޕ5t�C�#N%�0l%�J��?�a:�P�rF��fy�>��m2���fW�K�د;\�^U̺�Dc�l���XɈ�B��H.��Ğ.����
n���P���4�s��g�����yoY�{m��=,���[u�;zw̜1�hu"M���(8���=L���R`��+}|7��a/*n�9�?w��2c8s��T7��H��hBZ������Ycc�b6���+zt�w�+GH�ǎ|�Z0Ibr�2�KbG�(���U26����Z�R�/n���[�1o�j�뤭�axe��H�\G.�������)�u+���R�>��Uu�����jx�x����C��O��+�L&�3&�4�1�s�*�ϻּ������˚EJά��ELi�q<�MGse;o��\�i<ʽ�NO}���}i�8q��!u��q7g����7}�����M,�Cx+�X=�0�u������=�\���j��Ofm&{9����V���9^��֤v�7�Y&��eF2�t�����'0�sʰ�]������twK[C:^D,g��5�+qB�Ҹ>�8�-w�q�!��q;���>���;r�3����jД93o"{s>���Ǿܱ血���r�R�Vf.-{�3�����lWϲ�����,xƱTΥy*~����qmP�xe��E�X���Э�E�>��~O�}r��`b�߬�k�V=�������T���V$^��M����J8�a�L��r�O5-��A�ڼ'�`�VZ��)���LT�)͓�%��d��3^�X=aNH�1N%����=M�}8׹dL����!kƃ6��F�E;����7�9�El�`�be��3�6a2�Kaς{}��>5ɔ�O�pw��A���v��'��Mx�.!���]˱�\��3���&9࣓+{���|#7[��m������f���҈�q��8�.��oɎ�Øu��U�Ξ�\���d!-'��$ˇ���u����-Z4i�7oۺ��3����{��$ I?���$�b��$��	!I`IO�H@��B���IO�H@����$��B��`IO�H@�r��$�$�	'�	!I��IO�H@�xB��@�$����$��IO`IO�����)���0X�;�/�),����������0$/�c�ٛM��Օ�y��:�k#�b�{��m5+6�`.��6������{`�hd�-N#���ֻp�uӼW�W�-�Ҫ���ifХ�Ŷ�r�owm������/s{m�m.YI��o3�k�i�h-�3�^��mm�Z����x�$��ҷ���7����l+�
{�  � ��h�F�&�   44� "��Ĕ�T0 & �L  "��	U(       ���	T�0 �&   �0�PI"d��i��L#F!� Q&@A��&��z�)����y�4��/> "���I�Ut?x��
&�U�O�d Aj!��}	�X?S�I�Uq�:�
 ,L& 9\�� Ua�L0" ������;Y�Gӟ��;�D�P��M >f�$%_�;9>7h��`]���o��#��c��NE���r�B�MU���j�f�D�{r�����LeA�k���\�)_̲K���W�Zb]B��j�l���U��j���Íb���V�v���B�í�)�N����9LJ���=��.�L�$ɹ�L��n 1��V��3�\tR��(E�@j�)=�.�m���0������KA[α������/�ؔ���ML@ʼ�r��Ƶ����E ��9�(طZ�(�t7w#!�pAYn�ֶwK��k*�a���(a�Ce��EE@I�K��Ӵ��Ӭ�;8��� �l=MV�Vdܥ8F�3v��S�[���ajm]%�uq�V���U��Yo/"�zEp�-��H]桐�)��n��EJ*�&S�E
�4�[̨ɭ�w(�d.HL�]<PO`nkJ�ב�r���
3���o�-TV��B�����t3M�Z���q%�,��a�uX,��c+�++r�P9��6Yn�:ֵ��]����؝�UM���Q�Uj�F�I��ZZ����쩅�,���4%�m�B�i�F	���lFof�°-��#�r�_�i��r��`�^�Wv�6�U��)S��[0�w
����@��)j�ve͙�IK
���fEw����܂���!�n�:!���*�� �&U����1(����P��C�m^�~G���(FvcV��&dpc-j���e�,l�F���4l�l��ێg�E�M���m�q@*`�䵹�2e1���г��%�4D�lf(��n%���c�|�;&'(�Q�h\� ��6�D!����[���[�-��������X�A�@��;�ͮ�»6�}j.�+���;�$�G+3{���똥.�]:�v[����퓣���8'W�f�{ \ށv#�_mD���/$4� T��˦��2�ײ.��>�`	]M:���Gi�G�w`z�Q��L}�C��쇷��탔����������8�(�I��s��E�J�Ƿ���g��͂�jǊ�bN��ڜy�$��0fO{`{3x�xE+V�}@��C�<����;9!�n�6)����X�9��<��L��p�{E�Sv兪g�2��s�$|1%˂]Q>�cѓm铊�,�;�;2M2m�)��׹}�b5'<�ȡ�İWX���:���x3����R���wtZwqJSMg���sib�rmmw�o�[�v]BGV�S� utn��Çtଢ`��l��ޫ�qv
���Vޘ&�}��ko�,Z�qO��%��ж�����x���
\��
]�s��S;�k�v̆Z��"�d[{+�3�����ER�s��6��#��������}Y4++�r����
w�MQշ�FoU{�\�h�OD���ެʽ����WW0����
��	rwq	g.t� �z���˦��T1(ĕ�5wI�+�*��$�����y���G�K���1�M��r�e2)�+�V�P�V��f��d��Abm�����\�Wh�y��#�5���O�����ҫ��}�n_.���R��;�`p�;���)���N1o�W&���8A��$�a��Õ�C[��S��{���;a�eq����6� *��$Dm�ST�\S"-�K��T�+�%u�>��~?�7|�O�p�?����y�Y�0eje[���j�8s3(v!e�;Hv����D�X2`�V5V��;`~I_���_�+�%`_"cj.��,����*��
��1/�|��`N��]7���o.�_��^@ٵ��e�p�"l&�++(l�Y�c�+ކ;��i��L��Ey_2�n{�桫1�R޻
0x 3;x3��Mc���L���/U����ۆ�p������4ݡ���U�;��v�J���`i�.���npz��h�Ŷ q偹}/F�e����)4��.�U���''�`C����o��݀B��

�./j�\|�_ee��-�,�N���^��]d)�����1\7
�׬�6=w�eB��˳(E�g�B�*����)j�B-7�Y����9�a�����7�%$��r�u��¹a��\��� ���tiM��)�
8:�v�o����i�(Q`قP��ۯG"i��P�/��
@�#HP��p�?Tf�l��XƵ�f*�Sq��sZba	(~��!	�uۣh��wI �E�&ද2�͘�+jAaW2.��PE
ֆ��T*���3r]�!�y�r�5����<W�[dm�`-��u#U���J�]hW
��WZw���� 3К:J�1+v:�¬��FQd���G/�j=؆80����Q�c��4��TػmuBL݌pŃ��+n��2z&0t.Y�x��륊zhpVj��_!cQ��h'�G��,A�Q��!���J�|��vl�a���p�����Y���Kd��<�� SoC:�H��I�&�5iZeZ�jZ�ʵ0�:.�D��@W��jC��aS�͈Jg���۞�+o1�j
��⋫�Ȭ�⇵��$�tft�/�[��(�p-��tS�tL!�g�x��DZ�T�BJ���t�1�&$��} ���P�P(}A)J�d�PX,ň�ъ�"�x>�ǽ׸޺��㙱���߾�
ʯ^��U.��.UuL��`���VYz�= �R�9�d��)����m���� ��N��O�MI1O�}�H�0��f��VĀsd�FP.t:/5g�wDÔ�J�p�̪�]m�A�#v���c���{p{��`r� ,��t�M�k� B��"�b��������#�6�aV��J�p\��K���n�'��+�9��zM�}�&.|Ţzp��񵠘"�|��Cj
"��}kb�y��c]u����,�cB�g��PW�6�X�E6����jD�3j�*����8<z��ng:��4���0��r�ߘ6ɔˇl�e+���q��_l㗏�.N0�&�PS7:ɧ�L0¡X=��i�ԕ��NXaȘ�3�bVL ��ɇ.��M!��p�&��>��*��F����e)M�mp�s\���Ă��6��5�>fL�`�ĩ�s;px�v�S׉�',�N�nXW�z��s'I\�Re��w�p�Ei+�=B����kt+Vm�<�S.�,2�AB���6�|f]�~���8���>�>hU��n��'^H��wG���xV��CU³J|��§����]��9Ǻ���f3N�m&0+��,�.�e۶
��=|�z��N�����ƌM�ӜR�ɔ�.����@Qx�=�-g��2��Q�� ��n�+5�ץ3�����b\~�v�{ݭ�:F��~��ߥ&�x��IY��m�3)0��;��t���{}L�ӧ��LZ���>��!��iD6������R
u�u�����)��+%C��t�L*q��k�a0̲�6�*<�u?3����oL|���_{�`��6�Ns8ŕ�:���`�iP<}N�� a�����x�r���(a�M�_SR��=p���5���&�Ru�p�y�}gq>�)���3��e�$,6��~�3Ϝ}���6�^�4�>G�-fSCѬ֩�Y4�&��0�t�����5�8�9L$��p
Ak<H����(`��Q��T㔃�z��a��x�C,�<M�WHi�+�:��=�ӣ���`]�=M�2|��b�}��t�3o�!���M"@
ݱ��\�R�]!�H^�vI\�)�|��3v�@����G&[�Λ��ͭŎu!E��ص �7W;Z�=�ewҰ;�����L%,�ȸ�]��)�z������������NR�����i�+����˝�	��vr�Ԟ{0�T��R�^�IȢ����J^fgZ�R��%6B�ĈSSe^M�������  `,��+ �QTX����DPQ��ɞc����_~9�x��+��T��f.0q*a�a��L��z�L9t�r�̒��{���g�2����<憓	�>+����븗��1��ȡ���r�_5Nw8m8�t�_�����n�;��׎�r�����3�s?-����*2��:R8�Z����&�z�����4ʭO�p�o ̇L��h����5e��SęL!�����M�a��)]��9�;�4�g�0�&MP�yK�t�jý�fx�S��;��mRe
��Df�\ �Z{��,ڝ�JT����J�di���l2��C�g�@ņCP.߰�s�R�ZGu��)�A��Zۍ��`�&n���ds�(���X�捁��x�*nnI�V}Q���|J�}$�|�d"ȴ�D��Q�mO��ɗCT�iTm�=R�7}OS��Vؿ2t�7�?^�AJfx𗛮S ����`�`cO�.�x�
A�.��6Y*3'*�>Z�+�;��Bu����7'Y�tÀ?�
.u��U�8��%�5����`�DF�cC��k9ݟA��Q+v!��nmR~�t:�i�sgb�*�˓n��Y3u>NqR��h`^Ke�t8 ����e`���y����j���G`���B[�Z08�U̻�U�{�ɨ�z~�(�QE��&v'���A��^�t�9`�k�wD���%c�|A9��!S�v������Q���oy�g��CW��6\�#���g�Fr��@�e��~�z���8efU��ѐ����e˖,��0Z���<���幙55v���@��բꔤ�ŦV؍�{��M����*�P����i;U�D������;i�F���"#\#���>4�Nۇ9WNf�u
�dĉ�<�<=�ӯd��t�����]Ե���5�=X�Q��LB�ب0��Y[I\�m���1V�<�%�q�c�n{C��uǹ�v�˽s�_.۬�:u�����]�B��
�5:�Y��bl�'-�ff��XR�IT�*�bLk^]�Ǽ����2�
PF �j�PF�T`�
���ȉU�*�a͞����~_/�P`��x�5�we|�S�ӓ#w3� $��!�'�$���P*c���p!\���L�Pp�H��k���Bg�����A�,��$$��BL$���Hq�HT��Ľt��;�+-X4��y��ޔ ����W�����@�	8�38fod����zi�/�ƞ}�#�[N���u&�����X��d��b�]/u��ܲ)���gٟ��c��XZ�Ϸ=�@Yu%�#/;�xk���Ğpݕ���^Q����q�{�0z�+��.���d�ҔjϚ�n�s��-�qe������l��Su;���舿��GI�����yH�|FP���N�T!v�o:��md��J;�����陋��'D���e+%+L3x�$D'��G�Hޱ�#��v�1+�;���.ח�9��
�j�Jc��
�}��(a����+�c�y[M�U�G���7]���8�D�F�n�s�lgV@/1{S�������;��J������������<C�f�����4��y[ݞ�\�]�A/m�V>k��=�����=V�޽ˮ����#��h�{..=��jOu{}r�VS�n.��K�����o�\8Xbh�Xׯ{.�����͛��ӹ�z.�'�"�������#�����,G����;b�V��o��.���S0�*�1��?���\$m�rs6:����A>�z�U�m���xQS4���gc!
K�u.��+eF�zThˮ=Qs1���f�j�ܩ�΢�o>/���Q�}��WK=C�GdF<^cbc13ib�PQJS����V2'
�7IU���2f@ 3 �"���U"����D@���ջkv�,�7���X���k(��=~�4!��뗂!�lz�Uu:�	��F+aU�T�"�M�g6��l�g��쾓�)�ա/a֯�� K?N^Xv\I��
�N�{�d>��ъ�r������u���y4�=OS��K&�ۉ
V��h��U>+4���:y��뛧Mc?y�߹=���K�b#�G�0}Y�5����y���Z�9���"�-�h8�f�K�e�3dl�����N����{��{w#�I��uw��9y*��+ȼ}Q���we{���\�\���73��u��v�o$U�W�o���zu�6]�N��c����4��ihS(����;������R�<�$��O����ֹ�G?}�?�oW�p��v��P��V^̣�����h���W�-C<���ӪӨj�V�U�m<���e\��33���k��6�0�ءj��k���r�}߹��ȑ�dLZ��5z��W%��/���ǻ%�Lqb����fw�.f�̛s��7{T8�f��f:�-�H+��y�"��dϯN��Hk�Q��&��&��ox���H�>0�x�~4#�K]Vj�}L���M������0�^���#��O��a�4��x����j��5�G����c��L�v�쎻���j�m[X�<�֗h��[�ٍ�i�k�*��+�l�b=bPQM�#�R�R.D����#(��)�;^�t���]ML��I�eaJ&J��R�U�E=#e�H͖��2��u�.wv7d���9���]��.����Y\��{��d��Q`�DDTQb�b<� �ɜ�J�+*���3�Q�d�S�L~~���^ ƄI۵�[���ϼ�I��}�gG6Q��Mm�Yw�Snd?�q=�g�{E��ǛrfP�WJw����~�����O� �Kڤ5�\8�� ���:����|U1Q����ߣ�ç�����Ѹ�K���]��^�%�I�W�_Q��s5����:R>��P�_�-��mx��E�6�U~Y�桾�2����/���H��n������܌�����͏�ud_���%�z�<���	�6Q����;=�[l�T���<H��ޭ�Z�u�\��yڵ`�37�OH����N�T|��3��X�M��35�����m�מPq!v�"-؆�'�Ǎ�N�=�w�댬����fgp��I̺/�ޮ����k����@�r�΃'��Mѣz�Ņ�r}�j�GZ��Yu�7�\���X��{��sf�yt���<o/ ��8n5|�~L�������^}��KU
�/|Ŋk={[���Ib�ʩ��fff��t����
X��=ϛ_Ѫ�,[:5An�~�u�������g����+��xw�fÑ��E����{�%)�D��r_$� ���N��u��G�:����O�_&�F��r�<r�;���كw��$���RV(�y����ȣ�'��g�&/����Ur�L]&��̏��RS7kե/"�z��z��X�3˫ʟ�(�Z��:`���Dkv*܊P�m�2�e�t���o����.t#6��`�+l:�O3�o��2��j�5|D�r����c�� yA��ě��X��3sgl\��ɫ���4s�{ɫalnk�I��UxpO�S�"��<L�K)+0���J��c���;Ώ<7��'��ʖՕ�ը"�-,��j���H�|�f��hս־nNU�_ݛ�g������I�l_��v�az�G���÷C�i-T�B��̯�t���/!�t7����'��L��̹/_7���s�ꪢh0�Z6'���ȢA��Fa��� ��]Z![����L)�RɎAD9&��s�U�l]%��r�'��ı�����=�(Ȁ�2b`~��rF��[���M�um�[G �-ճ~*������-ڜw��4�g����6�諭��Xxq�i�I���ِӹP�+�Ȯ�Hq�s.f,!y�i�������W�U�Wg��ul�qjw��g>h����@pT{�:l�˗�f\����ű���>D}���v�(}��^�2s��
b�#jW� ����z��G��7�Ϭ��=����%��{sf���(�L��:���ᘚ4E�`�Q(����X3f� =ģ��a�Q�ws��1b�x�y��g��(C�4$���駳(K�3kv�˰����6�h =2��?v��<>�����ryӶ>����f'�*"Nơ��y�/@z��m�^�B^���-�לޖ�=�xJY��K�CI�Q�M�{��V��ĉYyW=�7���N�+�q��Vm>����{���}�I�J�j��e,�yGsȡg��9=��qh��]�f��j���fw�T��\�A�o  EX��� ����+,�S2�<��1u�y�bhO~:��]�	L� +:��ys��+�Y6*u��[��h���3������J�.���]�gj<p<�Df�
U&���������b2,)����~�ԍ�)k�W�Ni�˫d��	/yN<�Yg��s�r_+ə��rЍG�ѝN>ј-��\Z@Ay�H7*��H�(t�������5�w>�7�mwIP�+Y*
�R�RTX�E@m �X�e
�#�B��g��I5j��=�e�1Cue3c������^4{u���P��c�vg���)��&d��ޥ�i�g�+ƪ;3sV�C�IA�w�n�w�t������._�"�d��c@�a���� 0�.F���Vkp�%C��8t��P��|��7R��(��_���>�J=���a�=��/�w�fV3��^q�������)�P#��z��:f�J;��>|j�	�y�'�E5:W��zU�^.fvRL�@O��վto�{��]�K�&��4��B�̓	HW%���v����.�xx�Y4l����6�|�J��W�mP��[I�����N�yMP�o<�pLK��S.��~���y�^�"��u_МA*��ע��d�J^$<&�k��:��*�\V�2�3]�g�X���-�+G�WOR��?0�YM]�@C���i��K6<��t�t74�Q�I��ڬ�ܿsn�a�|��ݽu�}��b����c�<�/l�fβ%���Ӎ����c�ow#�盝�Y<o�X�?3�v�X@�??'���Gh*�~g�r��@@�hڿtX��
�;���v����v!���6�^2��<�BW]<�}��l�>²�H_�ʸ:\-И]r�}iQ���{b�uU�1u罂s|�2���Vݤ���a�@m܇�8��9�5^1+u!�L[c�]�5�}�pd���KP�\ !��g\	�l��%5��VԌ�����.���=�Օ��`��F�֠{�#t:�/�r�yMP��"*�{N9m�f�����LOqܬz���z�4d���n�ƛA ��B�����xJ�
���t-l��� M�<<�/�d�v�#��*�P{���M�e��'XG���T~�T�E �V�Y*"�������KF�֊��A��m���"!RQUQB����O?8�2�a��l�`�ٹƬq�d�w�ҥ	KQb.N�~���RL�=�显����~�����s�Qf�{%��t@�F���wB����h=�Y��Cֈ�Wz`��Cιg#���6
3�K}2�V���4ee���ҜѰ;�����<}t��m�}B���쎗��!�U�M߂�=y$�&m��0��.��gyc]:(��=^����@����q��� WK�A]!��؄4E�1���~h�=Cf���b�ߤeU���.�zϳJ.N�p��w��l�꾦Bá!�_��x��W�n��Ki$x1;�eHl+f���J�w�m�O-�왳�t�q�d=�P��|��:g�}�=pV�[
��R��!�A��6O�N�ȼ��=��������ŕ�]�}�x����u�M<Y,���������23�D�%U��A��p<U��+��v�����4Km�Q���;�h�˃���O�䕡�Es���.�o���9�jW����h�=�jsf5W/U��/bm�I5�c�\�ۧg=E�{� Vek-m���&�V�®�̿:��ʳ��au�ɦ�6Vn�����I]\S,��i�;�b���4 ���@x�*ڼֆ��U5���tR'���w-�1��/��6��'�ҷiMQd��ԇ+r�Z������m�9�i!ꏤ͘#4��oy|+F�75��]\Q�t�f�Ü��,�\������J�)*��)��Rh�2A��ov��Ge��֊�K����\x���
���x����Ĳ��V g�t�O���c��D�f�c�#���!��Dkb0T�U#j�#"�X��ڵ+H��l%�E�EQAE�eH�`����k
�V*[l-��-�*V�ѣ,Am��ն� ����m,QV�{�s����ݫ� �c��2!��k)��C��=��Cw~ie_�V�D��=-ݤ!�6[�R�wE`�{�"��7�s�E5�/w��O����fc�#�t�D�^<�ȕ>�t��km�7oYC�I�Fֻ�IL��-����0=S����hl�v�Oa��l��Q�M�N�hhP6���s�I
���C�k����~��-��'N�$�?���Do���`ha��������\5� �c����G�P�j`��S&q��ϕ���k�6��;7�����䮇>�"��:ö+�0Ј}+ТGj\K��}ݺ��g���(�|UBl�'#O�ѷ����o�9L|��D�p��Zͦ�:��6砻�:��U�V[�u>#PT{�%xa4�L؞a�.��Ѩx�E��'e���<�sȦ���We���5����ĬS ݮ�z)F��m�H��al�^S-S���uH���B=p���V�9�c �h�^;x}���ؕ�(I�B�V^/c�pR����c�iKW:>04����SFĹz���Z��TH�K����X�F6��`z�~� ymo(���+�[��ϖ��z�����8f]�{�ܦ�N�����YCp�:�`����P?bMHuƮ���K��3$f�x�>���a�-K��++���f�44��8^��#L�{CtZ�Dz�Cu�f�̼����L�YՅ��Nַ�-��l���)O������Ҵ��-��,ď=��6T�7��dT��}�6�ﺦ���QV+vm����5�q�W+���'tR���9N}܎wZ@I(�p�ʙ0#N�N3P�f�(���IV"!Z*�,U��ѥaZ�m-�m�e�R+V*����#@ f ��	�5i�ݺr_z��w� 3X͊G��_m�<��_��kpmx��_Sv���ZS��$�Y�%M^>�cqR-��t�=LT�z��1.i\��+.��d,,g��(įr�>9+���e�R�d�����&^�egӷ�8\N
�ZƬ���1ߘ��N�G�;o��cY+8&@���1����.{�c�����C�3�O��K�J�I��r��{9������^�E\ol+u�q���F]{��̾�������~L�Ҭ��������nv�E/g� �s[�{�+t"�XR"���K3�Ǎ�n���E��O�K��$�k�V,��������cY*��S���;,�*ǡ��_���Q�������^w��\�ъzt�x	��)��9[�� *��(�j��W�U~�M������xS���?f�F�;px�cF��u�K\^�����-BJ�t��<�O�nrne���F/�6�OEk����u�Vg�|��1����Q >��b �pZ^�pPaN4�#У����7S��k�}��N-��웝��S]�`xfd,a�mpxv�"���e�)c8��k:';�ߖ���r_>}��w�u?,��r������������G����阊�6��󦽉x腤X��F���LqU���Ej��|ǯ���~�������O�J�TV"�I�B"�̜��D��\�P4����3�md���1����<�T���
P2H��|�$��* -3�B+!!h%t�&�Q)�5�� Xl��!��ؤ" /����B�y�������fP�Ҵs�4�J�7�
�C�����U���HazSLR���# �A�"�=E�-�\2@_��ǖZW���hs(�/�a�/�"V�?�:ӄ� �Jۃ���O����h=S��tkNH�'I�(�����D��@��i��B�HP�����m�d# =�ڐ!?�j3>�]KF��\/~��5��D�Ay�"��\�Q@T� D�W��W(�C�)r�& ��A��
 �X��r��Bm�p�&�����o,���L��DѺ�����s�~���� �N�"=ܥ�l -����Q_ �?$%���{��<S�M|BT@[re�!Cx{e�����>�.VO���4u!(J`�z�����7Rt�]�X�Sf!ᮚ!�_����L�!D�$$c�Ýb��ie��cB ����L ��CX(��"��(������2�{`yA) o����'J��dbXdWYd<й��"p���C�J4#l�(^5�"��bP���p���Ȧ�Rޔ ����0h=7�}�fKa�h�pJ��
��=\��!��Qb�G~��ǫ`�!}��y���5��wA^\w���>G<#qҧ>|^���<=fԧ�~�_�H��n�m7F�X��&I���)n�D�����E��vg�9x�]�h�������L�D�SîB�-�t�-p%���v�Z��Ȅ��7�xw{�h`�*n#_�5�Qx�!�
�2�#8,S\�ԺbAۀI̓^�vf�I	��t^w�X*�!��f;aQ@_�O:y�Cp���7�����ӱEzP�q]�p����[����W���JX�� � �>$�r�Ds����w$S�	nsP