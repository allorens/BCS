BZh91AY&SYV�ƭs�_�py����߰����  `�^�       �����H   �     4�b&�       �P�� 灈>�p()�>�
         w �d��;�p7I�w=oF��G�1�f�w��U����t��T�z[��öл��S���B���pS��uﻩU�d |� �{@S�QF�p����
�����v�0��v�Kf�i�{�x�ol�5W�爴�g��\�n�C�S�oz/Q�sw�Ҿ�8�m�|@#� Q��U��wm���=�m�[�]�V�0u͆��oz�f=;:-�ю�̭V�n��kϧϱ�i3n�|��@���,{���[VX���ٻ�l-ۃ�������G�%�	<�:=ۣ]�c�z�m����_j]`l�U�o �   �oU�2��֚���֍-�Y���v	�U��z��7����FmL���xWy=�������@     �hi@b
)R� �D�� (   U?HѽR�(��h `&���S��%T@L &�!� �2`	M��%J�Ѧ�C F�1MDT��&�& &��M11$�&B ���'�0��zSC���e=OSR'��R��0   #&F G3�D:m*�*%RB����ma,u��׽�q�' ,Xҿ��"�T C���J'�B   ��A*��?O�k��籧�GVo��9DI#	_�EEP[�楡�Ԡ�$���U@r}��b����p$$�7�b�(&b�G���<�>5���3ؖƗ����I�p�˒��s�M��ZN3z5��MW	��b"�'~ΒYu+wzLA�I��o�&��sBu�);G5���`��+���+aZ*$K�I��:��:<)�5�X&�&a�H�:����$�^�q�q#��L�}�ԝL�����^�5�W��h_N��2��I�/Z�Z)܂o�rq&���>�I,�H'Y!���M�)���d�����}d��6ɸC��2}�Hv�s���d9%����Chm!�:�xM��!�oRM2hMi"bp��#�2N�I�`��$DĆbC>N"b%��J��	�H�ɾ���L��tH���E�L��'XL;�16a�$��4%�"s�&�:= ���Y,ѧd�5���6�����I�vO�3d�lD�"w8J/�D�X&�N�"h�!	�0�ݓ�~�$��h���$�"Yi"%"#��j$����C��Dĳ6lrbGD�2aC�D�ZDKĘp�H�Bp7I9Ĉ���8`�p�,�|��Y�������4Wճh�h�,��H"'t�:=�(~K�br���E��ԔA2$١�&	�DD�l��BDNi"wfbM�}������6t��6o��Ӷ#!�I���
DݤH�$��}�Л�1�,ѡ(�g�!>M�siؕ�4��'&��1:j���&�&�#ȋډ̉�8�+���p��MY݈�ggjpu8a���Ì�L�h�����'GS�#�^�NnY��N�Q�s�
��5,p�1���f�4;�#r��Y�3�����2��p��l�j�5eM���Zq:�N�9�EoGm+��R�?X�&����"#˨�t��0G�N��h��EPMDn<����8.T�'�_�R�0�ǻu=��:s��mK��ƥ��Üjt���g�k�9%�YV#��G�D��h���p��ir�q�TN����]���lA���Z��	%�g�n|�9U��(�����M3�#*�#����	s�>GUQ��DdN���H=�".�'�"<ʈ���U(GQ�D�L0�*UDG�����Br56A��d�S�;ʉ¸��I�C�d��""�aej"<�DE�D�kR���A��pӪ�?tk�c����5(�'Ȏ�Q{R�fTD�ږA���S�D�$�*"q�K!�O�j�"��a��Bs�K ��8i�J�Q�TM�EB�O�j�"��̨�͵,���?&I�h�f�F�#�Q/�D�"p�ғ�:��y49>~;[�C+��'�̯�M����9M�RZ�4ޖ��;��Q�T7Q�����+�.TL�J���
��8%����G����ú���dB����sZ��O�#�4f��!�J��x4���gC�gC3���0nh��=��L�W��òt��*%��j1��9��
��"t�8R^%'r������"p���{=�^�=��C���p�C�YE���ugt���՝�;�^��.�gqT7����#<����3;��@_�骎�Q��lyڎ]G�WG�	�9ĉ�U���W��d^��sY�k�1����=A�A�9���.c=z�p���~gW'��x�����"��x��3Y�I�V�v��ݕ��ֆ��t����}T�-'�,=���{����j����K��=�8s��{�Ӡ��@�!���Gq���'Y�,$�oS��<�c�����jp�K�q���+�C���\���>�1{+=���fyu�u��g��1�0��sG�1p�O��8��e`�=P{dg�_���i�̋a����k�2�|Ǝy��b�[�B6[=��׸{��f���9��52���钌�0�%ᣈ��N�4�l���W�&	8=�&�FM_��>�!�0�骳C�tE�V96�(��&DN������lM��+d����;R���I�����YVhu8�;b&�Id��"Z�ᣯ�,u�_pF�Q��5rW����jUTDy���jV�ӹH�w)w+���D�e"_Y]4u�"=�VC[��#�D�5)�J}>Ϛ���r�8�R���%|��R&��V&�JDˑ�I�ze}_;�����9���1�ac����eY�O��JD�r�����|ԤM;�{:��J��\����H��X�y)k)8oL���r�4�R'1��F?L/�{Ϝ���Z'���S$Gr	rRt�~ãQ̕�;|�dM�	�>�f��r�E�CȜ69,N�����g�J��jD�M��G'dN�+D���B���n�J�DZ���5_W��F����PE�&c+��0G2V�]���'(� �#��r#�J��K�gJL1�W��49��j�0{$��A����4;�.Djp�Șk�Uq���Y"P�J��T�f�w�:�?'2A�|�H=�r�d�y���v'aϋ���7�\�N��a�z�šڍ���-�K~�߻zk^]뫽�]b��Cد��3�\�U/�\�N��vh��򯴶�ۏ�o�������C�OS�\:��{�p��<��7�c��X��i��0Y���/�~[�ن��߸j������ P�y`�0{�t~Ny�:6�PVc[J�i��n��
����F�	��z���Me3~<�s�`��K���t�:�W��W�8�ƿ��ܙ���������~�cc��
S�rH8s��ߓbS����&d��2�.v@�����{���;f^��72璉���8���<�}wY
}�����6tg�	G��#��]�l���zޞƐi�醖�s�2I4�F=!3�'<��}�h�C�a�|�9>[�>����r%���q2d����[{�DyKu����wqg?nrg?{q���Q��gx�i��g��f�>d��~]z%��p|�0�g	��|�b\��_�]2q�1��X,����f�����2jfsy��l��{$̿Nw�np�9�ʄT��E!O	N:<C{;���(�W�^������L�9��ֳ��p�]��rza������0�zl�BogC�I���^𿯧7���J~ͯ�9��&�8a��g����B˘��s{������| �NI�[��-����3���~�3��g��G?o2�S�����p��K�N���'���K/��^X�laS��J �|�\��lgM���f�Og`a�2K{)���Ӣ]�n����l�4�B�s6L��ϓ0�zp��n{�S�^���������.M��l>!�˼��ri�sl�BMyü���70Y��|�t��v�h�p�qk�`B=lK5�8p���)��ɚh�?F0��� ����h�����pi�raç�	sϞL0�JA�p�B�<x�d�n�4�Hp��nw���ڥ�ǹ��hC��OgM@��⎌�8B��w�i�A�(Y��Q�C�0rO�  a@�ZZ00��0���)�<x��ܚ}��i���~�c>R�����I�>Zh��O�C�r1.!�&k!��r�2���d��.�k�G4!�Y��O�,�F���~|~83�$KkŖEI?
���?ޚ|�D�>��k�u���8��u�Ӵ/��7Ye��:;����
T9�Ǫk���n����K������ 8��8�5��ѫ�ϖ/�u��bkQ�ܳ� �^�@)��ȓ�X�.D�26�D�/�ϼ��a����H�m��P0��+��h����5�Ѹ�֞@��Q������eѹ��I���{�9���>���eoq�u�k��_3���>cJ�>Y$T 4��o˷��s]>T�[��_O�:Cm2޽a�=C5XC��0�hc�Ĺ^/g�:}�J����rC�������-O�R��d��e��ӽ���g@���pK=(�~��=?4��g�}��Y΁.O���Ӿ��W���������5����n���$>T� `Nl�vfl��ά�۪��3%�]����g��L:���:}�xx���}���������'�\��օ���95�e��޹�bw�ɓ	Q��N�rP$0�R�9$9߭��:8��g7��}�o�a
p�јiW�M7�Z��^�Q�6�m�H3��)��>�4f��w8`�H1퐤36x�C�\�Ӿ��g��4��֎rS�Ws�:a*�i�9(c��8�[�DL!�@�&U|;�; ��O���w��2+������A��D��{K��Dv1��x;���;��S�xof�0�0��w�2zpJ��/=��q6�(2  ���.vCpc � 2&Rs�iFkN3�0�4�ǈ|�pf8iM4�L0��Yӣ���t�a*o)8a�d�)��!�ӇL:u��Ft�(�p�~׆�3N@e8x�9#��|���>�tӯҚt�ë[�{�N��G㵙��k٫͛������>L�7���0�vqG�!�8}�����p����4�iR���SQ�vh`�
p�3�iCO�2�6l�HC
B�!ҁ�>^)��\�d �	��d�M4'f�p������/f7�Zp��i���nf����|�9)͞�y�Xz�(���wѐ�p�:�J���t;����O�1�ש�v��'����t�2a�o���dӣ�)�{��������:�x��4ӧ=�㛓D�����`��i�/�U�Y���gy�|�i���.�C�t���3#!���M�������:%�����I��Ж��D�zr���|�<�m�v�-���^:>�s�Hu�S����gO�0o0�zz��Ü�͖N��������%�uo6f9�'ށ�׬�|s�4g\�s�9����\2_f��5�x��8���f��.�=O� x�N�^��j���$q�ɹ͕�s���aTۗ����ɛ��U�~2�
i���f��4�������vk�0�w*�t"���l�_���{?l�{9�l��gO�}��
���tg��(Θ$��gɳe ݁Jxw�|�|�'�v�p�'��Ç㙲��xc:g��M�?s4Y�)���-��!��`����F���M=;>_�pzp�g2y4ù�W����&p�t�3�f�1kj?)ÇL��(�׆��994�a��))����p�.={:0͙?H:w��Q�J�}��)��5����\pPw�XmƟ&WpI�9��?O<���x�2[d��c����U�gboVz�ɼ������v �Fa��شζ�1�]>oD;�?OLj��Bgm�t�ﹰ0�:Zy��	-�	/Q�9��$������H�l4i޷��]�*�M�X�#�� ���	���3�YB�����!��r:�U&44�������t�U�莛�S�n��Q	E��Z�5�I�K�K�e9X�Aŗ��˺���N�Q�Sl��җcF��r*j�ݎfR��$5�.�3r`��ؾL�VX�M�7I���UID�Fk5�b���Mj�[aQ~�k
|�mx�S����M��.p�̺��Yy���u����2�����L���3�Y>��;eg�L����#�c���nϡE�?WLm����EZ.ń�I�>ƚ���%#�P��};1����}��b�$�] ��#�Դ ��Ե��15K�>���e�C/Ш��@�pLJc���> u�|G%�**�L}#�:�2��cvf8cx2VV&c��,���B,�&I��N8cu5��Ȁ�}յ �����:Z�@>PE�u!آ����?�m`��l)Y#���"�B ��P
��Gb��&�*��А���m���l�K����w�!zj�3��c5 ��J�Biu����m�a ,j�C�l�� ���c�ר -$)�u � /�f�Y	Đ�U�Q�&��N�:���$-��a�2K.��'�@� mM�O{�8�N�!5Ti"6�RB�P�%�ԁԇZx��4�(a�M'%��w�����HOa;Y�X+� QA^<m�hC~<�]����̅�;�{�W��O����K�'(�Q���!��H~b���6�K�\e������U\b��WJ��[X���UqZUW�Uq���UqU�UҪ�V�v�U\ZYUUUUZUW�Ҫ�X������0�`����R@RDE!)$�"�"��� ,�F�D`�P ��x�{���ꪫ�Uqګj*���U�]��Ux��U�Wj���Ux�*��]*�*��Uv��*��iWJ��,��UWt��Uv�ګ�V�t�w��������U5��4BE*�b�k�� ȫ�"	�AHH�B D �A`� dE��W���{���U⮕W��U^+J���z�����Ux��U�U[Uڪڮ�V�v��U�*��t�*��]���"��UmU^+�U^�*��t��Ҫڮ}����>�>�W� #"��	�0d��}$�~	�W��=Z�{���*��t����U�]��UmZUW���եU]*+�W��եUW��եU�]�UW�t��EUx��9�t��եUUEUUEUUEUW��w��l�����\dc	ʨ�H�P�����

B :���Tj�T$* �PFA��� 5����(8�aa-��IuJIL�ʈX����:ǵQTdH�w���|����/ ��w�q�X�50v��;�'��lL:"`�&	�0DDç��B&�N��:A	B&���B&�dKBlM�� �$,DD�8P�"P��"&"ȉÆı6&�	�(J ��� ��>M�FH��8!ba�(�Bh�p�DD����� ��"%��0D�:X�l�!�A�<x�şv�X���C)�1��\,pU�+-�UA9$h���B���>����b��:�\�9dmX�Q:���Q�Q�5(�Q8Ֆ�(TG`Eceh!J8�rB�Q�B�KRd-uKb�e���V4�-�6�jH�J��%��e��ՕV�M��b�'\�)dIR3��f1�XI��ReRGH۲�4(��Q6�lV�?��V���ԪH+eV7T�'h4R��d���;U����!��߂T55)[dC��Y\�X&"�+k�lq��b�u&�`+c%$��CLl����ࢌ���"Cea�$U��X�V�7%��φ� r� �Ϛ���-�ʨ�]�$�-ND6'ej�Uu6��$@KU�p�Ȥ-�EW��8D첄�:���L"u���c��텬�W��+����E�qX���6���[+�N�aTj�����>�6F�pu�����;U��d��ь�QWktw��]M��;Ij����g��V&�l��>��F�eQVT� v��mUX䶅��5b�M�A���|J?�(�p�
���;��2���ӅF���T�WS���--�����j�5j�Z�Mϫ���T�ڣ��n��brYm���cnJ�C*��
儌MZG~����R64"K[T�+[U�F�F&ϝD���etln�(��� *�m:�q�k%� �JV}�4F5�H�~m���d��v��+l�억U��
�[QU ;��N�V�mi�F�Q�FJ�pN8����@bAa ��$%��%"XF�m�Ece �J�N�e���M��$���������G,���DD��j��cpD"�lc�-���!DX�h;Z�:9� ��)hʪ�Z�AA#��j�Q�5K,�F:R��P#��m��Vݮ��m��A
"�ڎ�ʏ�i�����ma%D+������8�mJ:�(�_É�eQ�$�r�O�kP����j�\c�N|�6I �m���/զ�+vE�ص�P��%cMD��"��FՅ���h���5�f��ߪ+m�0�@�?��UK)a]v9e���T�W�v҅-���i�*��19~�
����YU�:��:�Ȝ��r
�+SHRTՕ����VI���rEAT��pi�#MQ��R�b�P�A;BF:�I�#��(��pQ�H����&���X�e�,���
��Z�hj��b�6�T�2Ϛ�ϔg�IU,��+��9#�2�USn�Q��R|�#�5
��>q�$) |��_�>���|��%qJ@��j��#�B��%AQ6GH@���-mB�
8����p(�p,*>hdl��4�EU%����q�㭪��i��6�M9#�1DA�]�W�n|B����j��J��	����V\�b��)��(�hbh��Јw�9#m�km�28�}*#�E\+l>B(�jN!KSN2!aEE%�B�mM�W-$R4���6����\��,%UQ��i�*�:TՎ0crZ��V�Z���"�'�Z�V��pj_����e�}eGZ�
	�(խO�����@��(��W��pS�J�m�"%��*�t	�C>eR�Q�܍ߝ�b,�:�m��G��j*�+ej�Z�$�9ej�_��"�B��>E��B�:����ȑT�D�j�G>���=��ʊ�wwv����{����EU���|}���{����**�������x���{�TU[����(Ue*�8ێ8�lc[�qn�:C��?�y+��3�֊8e��b�%�D49~$�Q�7*"i��l�qW*4O���X㊍4�S�$j�d�N1�X*����)�VA��lp��&K,r+Y1���u�-b(4C3*��Z]��.e1pp[���W$	U���#m�	ډ9�@�%����V�Ģp+T��n�	 ݄�3��0���\��[jJۅR�,�!�ʜu�~�`�����&LM����v�Q�(�+������ڪ�bq���(���h:��bG~��i��m�t���QDUZq9!M:Ƙ��P ϗ�5{��]��|�^s�{������,79ǌ�7;��qr�����)�}�s�7�M��f�|�����9��.�{������9v˶,V��x�r�nHI[>�WhJ���Ɉ57��֋��L����救�@��d83�x<X]4ܙƊ��sFC�Z�r%��4y�;��p���˱��4l�R��u���IO������|���έո��٢�\ىVkJ����4]F���M�CX) H��]|\�$���$$��6l;��d�*�3��8sX�{^L$�SoB��&M�)�j���rX0c���h�	�F�z*���GO�0��[�un�źu�q��S���a1u2R���˨��J��������������&����ܱ y-�����M�V�A�j2x�ᤩ�V�d;S%�aQ�0+��q���dKL�����3���E13�-�����92YF�糽m*���f�`U�,i6I�ָ@��Tsu	6p�Ɗ5��aΞ,ه�	�`��٢��Y̜�b��9�UMæf֩44t����UA��$��Bn컗-<��lr8�.��Y�U(�F2�G3�w�lFP��Ϫ-T<d�rh�w0g)��S�&|��*!Ӱ�C���ʅ�0l�gD��0L�a�5���֕
�	h�S>��[�P��>�6�34�b�O�0n��@8�:H�  ��ۼr����y����H�V}r���\����ݺ��5�l<y�ǼOc¹�����s6�����Rr���z|o[�G�=�^���X�	V#&K���)0�p2T e�\��	��}�bH��u_E��6\73:Ud���*�n�F�,�w���\0��'�Os�<,�b�L��϶x��60ѫ�x�M�fAu|Wŗm�qa�I�L%kZW�iZDs��o�=Z�[�un��00�8h�$��&�u�ŒI kF�Q�MMI�g&d�S'5��+�0��/-��W��F�4h���_L
�i �B{=9���t�	P8n���N�O>Ұi�*�q�4G���\ȷw�2�FQ�&j�=^8a��*����5*D��袍á��ز�x�Kz㭭պ�V��:�8�pYh]UP��]UU,�L�:2v4�Oh�I��f�	a�UF,�/p�ɸQG
:v`��^Q!\�h�&�V6���we��:jz�e��I�{��<�MJ&d�������4f�s�~uǕ��W�W\Fֶ1���V���R����Է$qE,��: m��L��
5Ӽ����TR����2���޾�ٺ�)�VQ�.vLK,ȕ
��0�9�ܝ��/%ΰ��0f	��v{����=jB�a����:p��8t�0L�`a�:p�S�n�����7\���&j�����7��dN���/�B���u� \�Uɕ��ޫp���__T�;��P�{��KֹkM9Y܆���3W���35��7\�Ի/�����]��v�b��j�������j������~0�sS3;�r��ĸYP&$���FcV�CC���%lrh���K]���t)��
���G��ƌ�}Ń7_A��3�F����!�n���f��VY����_�u�8?���,L)(N�aӂ`�&	�00�4Yy�ؔ]
��&��x�fMM�X�}߯˟h\Y��9�mxז�re��Ld�3pQ�$�6��tN&�钡��%g����s�5�����V�m�Q��`��7�����L3��Ur���Ub{E�#
����U1�p؞!�!��^#}�Ui��q�WS�ub4����b�bZc�c�ɉ�c�&>jӮ5��ZLLLx�1�6�&&&&1�8��|��k�x�����'�m��1�-�F#�j�7&5�bV'��Lk��D�bb_�j��k�6֓	��k������c4���S]�kk����R��FS^0Qk�>.��f���RЏ�_ȢxPg�%yS�<'�x#�����Z:ƞ#��ԭ%���X�Lm�f�X�h�5��1�Ʊ1�X�Lklk�Ԙ�LLt��)tx�	��|)�bxS'�Sm1"V�$��VѤ�bz�(��e�}��w�gwϑ�.��������|���n`.��r!d�5O��>A���d�;��6מyy����=׋���]��ːr'1�!cjp�Znd�>����䷾y�����}�nf닕g��6C\2����M�/m����z�v��YT��������]�{��|}��z{~���Ϗ7w����U��37����̻��}��*��2fff^e�33=��}��Q�oͶ�a��	�tO"C�6Qw*������&��UT5Vb	��Ȉ�̀(Pȉ
��,I(NA�;\�M2�4�pOP�&!�P#ꚁ����ĸ�Ȇ���*C8�4���"`aB����������3%�+��e�V�h��1gq
��00��.JC�C��7�����D�2M��B�%w=�&�(rh�cKP<!�r�������sB��Z���n�I�� ��®b�P��Hj��U*����c[u�[u�,��p�����UUQ��F	I����f�/�R0jJ�v'~�NCEq��.(&�9�J�4��/I~��>ԙ�޴^�6���Qd%l��)��;�L*�>���J(�!Q!����w+P�QGXnQA��ꔔ�K��d�]"n�0؇A#5
18Q%��P�*R����	F	H`��B�2C+%K��'�MtcP�d���Ќ���tHi���63Ph���cuo�[�qn������3��<X���kdָ->�Ͱ��ᘒ��BJrH]8��4�5�����g[�@1H���^���m�A~ռ�޻����ә̻�z��������=vKs��~Z�~�����>�^���8sR��ٹ����3w}b��q\�ۜ<:��;��*y����wB.��k^k�=U�{������p�d]�٘�3l7&�A� �p`m)]�+i-�5U++��M	Y�`h̨gc �y�	h��6��"����p(L$B�JL�Љ��dXܸ"``�``&>6<���93�̗�'��%B)�-�5H�H`�Qd��X�bJ$}��9u�1ƟSu�))|�3"�y��Nu�ު�v`3;62pI�*JI��6hC\Y��B�FC"f ��|x��,|��պ���-�^8��מ5j-�6j^f����UBUz�T�d�����p��ª�A��:0���j�I�L�`�D(�0lc��,��pa�;��c ���� �r����eB��$���'i.�t���(Kf�����8�2!����n���mK�qM���"�PCL��v�����D9L�j�!�r���_�5G��Cj�¤�����!���8\0d�b���L��Q���M�6i�6�>uk[�t�i�=_ =*O�e���G��UTJ'.M\���00�'�Q�IߕF��tCJ��P �Jf	55�������K�dy�d:�1e��HYƂɊ���/.JF���2��ǿ�-�b���=��W�2[%���G��F<	ai�)�R��$0��Q<��H��g�"NMB���'�!V�6!�$0 �jD�r��b%C�C1Ho=e"UT9���[p@�d�P(&�m��2լ�H�(����q72q6?�V���N���\z��z��$.y6[��i;֧/j��%C��D.]I�i��"\MA���XH�V	`?�K�M@����Ij�����_�U�W�v���P;�8%��Ix��m,MO� lB��	c�4Z�RD0 %�{�m���5v6J�A9�,H`�(ȗ��%ϊ�(��$���M�ݥU�oPȝY� ���5D�O��X�"f`M�B��F�a� �����E���j�yE�h��*�
:05�,M�O��wY��0<!�Cƨ%����2%�$6Y�|�lc�V���N�Ɲq��~Iq��?��ɼ��aJ:8��֔��������ٓ �ʝ���yUUD?�[�/��G�������������w�W7{�Μ�E�1�uvNc�v��wreӬ�E�c�8�\�B�y�����{��u�y�^__�}rs�����00��r&3G�.���4�Į��lڽ5sP�E(TB8(�@�Yd�Ic%��P�R�ƀ�(���S��16�J��RQ�n�]�]U�����
AC�E칄6!�$�T
��'aAu���N�M�2���L[@܉P7N.[%"� ��a.L�@��)&eQ�ʃ�4���QȊ����~�KgL�mN��b�51�0�\�(3xa�0S<T�`*M ,���r�e��[o�m�|�έkqn�u�:pÓ�>�Lu�&��/C�r�*�����b�ɓR�o�Q��`����eMA�!e��埪P�ҳb�+����/!�8��q�P�0%�Fh�[���b�>�1u������ɡ��Pj�����tY���q5e& 2TO��A�*�1,C�?4ՇfS�P�NC0��<XX�`B�B\�zK6@�@ʩ�& �#>��15�p�l�D)�d��N7�40�����淶���_��;^j�??:��6�>uk[�t��\z�n�y*�)R��UT@�[k�	+�o��^�b2QS,<y�f���X�ÅC(ϊ��X�D������J�����j�f`C����!�H�jo�C!m*�0nz�nT��K�b|}D���j`�Y�ql�i)�v�E��*}P��|!Ȅ��5�|Yu(�����Zc7=��T�ڱ�2��V��
f��T������kMk��O)�u[���ž|��N����M�w�T٦�WyڥUT@�C�?D���ǆ��ly�,a����%��]T�U'ueА3�-]��#r���J!�s>��4!� b*3�Z��9Ŕ[��	l8QR)���W������Q;\��d�,s2`ڨ�˚4¹����fkBW���H����V���7B�JC�
A�Fx��IP�؉L�/}�YwM҇LR�I�q:)܆��B��H�)�N'��1�Q���u�1�L~[�-�Ĵ��u-1-�b[�uƽcQ111�bcmb111-0�ZLLF�����SX��|��k�|���8�4|���M��������+DČk1�&&'�զ6֓	�k�5����Ϟ|��'�|��4��k�|�G�i�bcּ��`OJx�|WŭD|*�����D�,�)�����x��i��u�<G��b=M%�\k��51�f�5�-�'�l~�i�DcX��Lklk�1-11-cM�����1"bDeI2�����wSM1"bDm����OQ���^���yg����ۨ�^�T�f.Π]��{�/3�����/&�3[�Փs�|m�?v�s�۾�o<�g}�g/�����q{�>�b�kb6dm�$ִ�W�Ver?&TM�qK���1�t��7:�ȿ�����.~�x�8��W��_���Y6�����ܻ˯���
�@i�(w{��fw��;�a�|����qL^+�y���K�{�k۵�)%���3��!�&)��x�.Ey֬9_6<�VJ;�."[�uسq�ey�X�ӑw<Mc~����+�� 3[u��kA ���V�ݶ�XXF���0��&7��K2`��"�"�%`�_ʅ�R_��Qǟ�]��Vfo[�����Zs�go���_s�����gY����������s{���{�*�Պ�ܻ�����������}˻�{��,��1�uk[�t��z�&ڞ^�ԑ�*n�ʔ�[]���ԍ�+#q�dv��SP�_��}~��G��b��n�DD"Q�mUF*����T�
�	��ӑ�IB��Ea��A[
I$hi�q;!j��� vU[���K"$������`R��dQD�q��#%eD�l,���T�u?��"uW�}'͸�Hꃴ��ڨ)>j�
��q[+�_�$����
��d�)U���L�6ܮ"H"
Y�<[]z`�V��,�O�jҸ'-�hiKU�-%DD��RR([T���
+J�u�GA��+#���! ���*��Q:�Mƥq�&Z:�C�+�%T >�_�N��*�H�'�&�m$�jTA��8Օ�)D�&ӯ��apdrb��uUUD!�����w_����sܻ���9����rC�`ܓyy-{��|�r�b�A����r.�w=�=�;̹ū���}}��>l���s��L��;�^��E���}�%���6ݸ�f,f��ȟ�<}(�J�����`�;,��q�L3�Khh��tD8$C�	���1u
C�Z����D62%�:b�1��y0������D;:ł��%�gڄ=��d0̰��`�����`�J��E��M��k�e~*�Y��g%��O��FbYy.,�,0jPOC.2~�%C�g�;�f�h�o��u���&%@��T��ȝ.T�A�-HhǄ60�v�|;��RQ�e7�V�����c�|�խn::C�������+�UUQ!�%CpL2)i���4S�I�	�����x��p1�TpB"9RyU$I!.�KG*1����z&��TsU���$:Y��' �BX���
�aIсX(,�2`O�(�ɓMJ��2�W�_F���C;z�c�����M�%OFN'F`�����FJ��7ȗ�w8̞���e�ʨ#,
�v!w#Qօ�,fҟ�ƨ��1�<�m-�����|a��`a�:x���ַ$�\��4^�����J�J洗�UUH�|�7*Z*n\:'�`���QDd-ʕ����c2��F	�C1&��A�����`�0���\:!ʇ�
���
٩e� N�*��\+��+Y2b�sIu[������2˔�\Y�D5���H�=���hΠ��z!����U(00ІhX�83�Cƪ�9�������]��FЩ��g��*��!S��'��DU����t�:J����w��T�Mk��j�E��L���Q��:�(�/U'�Ty
�4�'���1�o\c�c�X���N��1ǫ��L�i<�^<�-,����UUH� v�(��r�`CM�(QT!������Z�SP����[s4��I �{30�3Ӳ�`�v�,�>j�0 ��\f�(.��}e�&ɸ �b�CXn*�@���YC	�+�fL�!��B�P���P���r��e!P�l.	i1E5Cta�(�&�I��2���e4U��
�G�I\�2k%Y�C0�d᷾ �S����NV�Wulq�V��>bص��N��1ǵ�W�i?�Ԫ?g��p/L�3wF�˘��W3�dH���F�$b����o	�qUUH���K���6k_�̝�{�B�ͷ��ɳ��,����OvUݧ�����t�^b��^�����L��ԍ�W�:�qf+w�ױb�6^n���곩\s6Y�z��;��L���_���+��J�!p�*Xz!��aTT&L��A�,
`𹂌C[C�o�֤�÷j[;
�_��\-�I����u�6Ŗ������4]C*�n��*k�VqX����(�C�;���Pـ.t�\N0̌0Y��Y����3���:Q���%Y���,�nDi�0��@B����+�qz0m��V���,<�9
� ������4��žzۯ���l[��!���+���nK�qUUH�(��S��:a� Sފ�9Ȧ�P��af� �sp�,B�9{sm��wv�9�S�f����{�[��3|�;���J��b(����FGF��CNa���v~��|6U6JJ5Ja��7wv�]���2oY �H]�O�F��3K�t2\%�a���\7(�\��l�!d�%�!��QF�%�gݫ�Ðو��+\LN�	U�gƜq�|����8�N��6Ǯ\�D����⪪��L�DK��J����oo�pıȅ�F%�,�3bS�auv o�I�YVp��ٺ��U�s0�A�sehk!��:Qþ�g�������޸���G>���z����#����U���s>�����f�؝��Y�S%�6 UT�4]v��p�4!���+���(��&����R�U��\�ꌥUg��-��e��ĸ;J������u��u�����c��Ӥ8l���5���|����%~kd��3}��C��a``���6Qp��E�A�A�f��hMD�}+��kً2�"֮&�xEW���J�d��UJ�(�P������5|���a�.�B�py�/ gP�nh�)���r�J�0�z�8��r̅�����C�x��8����r�.`C@�feB��E�`���r���!g�3,�8N���d�z�y�]?V��f���|��8���<x���C�C�q�js��,F�X���1��=�r���p�J��򪪐;����D�^ϻ��u�cVV~������n�^�}�/=���ǎN�w�c��j���{���;�n��ԇZ�ȳ^�\<.�~�s�{�k�޻�k_+�%�G擷[�(R�8T(����S��\35�&�l�(�Pv0�TLN��rf6LYUp����5�{�_����=e�T���I+#S��.��i��,4�K�1.�,3�rw�Jvղ��F�u����-=��f/e�\��Q���b3S"�^y��cyTV�˖��t���>=��}D:e��R�FQ?�$Μu�m�c屌q��um�T���>�?���E�VH�Q���ʪ�Jפj�ĩ�i6!+կ�&�|�j����B?b�Nh�C{r�30���n�j��*d�`#s����},�c��E
��>��4d4�2fWN90,=��V�b�&>��ơ�.�� ʖXr����h��cl�&�A��I�Qa�������6ȩU�
�Z]p�O�_�����J�8����Q�i[b�1�L[X��KcLcM%����Kb�u8��$LLc^1�Lm�LLF%�q4���5�bV=k�bb1:��$�5rM���ܘ�|����ɡ��b�P�?P�����>��y���洘cX��1�Lm�11:'�����Uk�>,�t�*`|7���(<]/��xYBxU�B8g���b||T�+��u���'�j�G��|�UOJM�������+��x|v�.����jxǌN&��&/S5%���{kSG�ЙE�1<(�U�F%ɦ��Dz��Ĭ�{@M�S}}��s;��o�q��eÊ���e'�z���Z�k��m���Hnyrw��w{VMY.�!��i3d�BI��.�w;�չ�\=�֞�u��Y�)�@���ж�fK�����\�W�G޵m���o�W�k̺+��~���5�Vw?��Պ���߽�yt��X�~�����yҪ�b��������J��i[�.���l�,���1�[���Q��=�5�kZֵ�7�QĽ�jJ�E6hƨ��>5I�9KP;8d5�T�=0e��+�s�5�����BL+�Ӕa����C���t��h�b.e�p�����+�{RٟTK<t�F���szZ0�P�B�UE�	��
hbM�XGQ�s%&���h�rY����R�M1�of���8HW04A�.�v�3�f�c-���c�:�8�Ƶ�n�W|����(���4T���tN��՚Oբ�:3ߥ��?D�0���U��&.��/�?��0�z��M���6Pb5�W����t`@I��"��G�NER1��.n��B���P����<c���Z4��Hפ��x����w^���<ۙO�mǮ:����c�:�8�Ǐ7��ޓ{�s���BŮ�ܲ�x�Y��-Fq1����-q��Oʪ�@�jp�9﷒���m^�җ�����-3�����랖w��v9����=�t��}�N[�kqM�'(�o����s=����r��j�L}��{���d�8$��g��/�v�+��>{��K6d7��ΎB��<V!�����Wֽ���=>3�����·��o�n�.�f�Z��
�-Qt,�Wf��/1!����UVT�fJ�-&�A'~����.��_���#�Q�H��[���e|��ٍr�[�t9����}fxvOU_:�����>|�X�1�,����ڕ��(j?{�iUT���OF��Q��������k�����~����������*�Z/O��5�+��c�_��2�&r�f�ɸ`��o}��9���'�`F�jY�,�p3&
��?��}�n\��?���Y����n��3�4!���4��W�x��>~[lu�8��[�X�ևM��}�\-qkV�i��UZHn�Tf7�>�2���3�с2T5��L	��2jf<q�jh��7�!s12'=���b�ئ#}�n�������ŋj�®.lB��w�E�v:jV �7:Q�bbgE�����2Vz���~d�q5�Y�
9�\��
<ok�l�>��]������k��D�O,��cv\��*��8qo��qo���:Ŗ�u���j�ˋSz�I��*3`Ȉ�3�1d�t'�8`���i�2F��ퟦ[	�g�;Xz���J0%�'afa�Č̉�9!�៌�G��2%�fA�88a�(��J��M??�y"���f�9�`Й�f�.��[a���y��Y_���4ۏ\[�|�0�Ǐ0��$0᫪��}��w'ղ�j|(5�j��4۷��E�ܹ���2��ʪ�$9��x��m?e|K�zU㛹y�;�L��r������{/*��h�;&u���N��B�m|�m����wn>c��2z��H��/����?li6t��M����!�`{%��5p,�>>�4'(_���F��٪&���3��Ahߎ����VX�C�x�����`��Bv	̮K5��D�ٚ,L� ����>ƍ���r@Y��<�J��6.m�/Ĳo��4���5��b̽V��p�94tȆ=gи_oh����͸���ű�c�YkC��w����V�Yzѐ�K=ߕUZHJ?~��К5]2��D!z�%J%CMh=�zl4&�������5.d��7"&��"""|3����e*��(�b,>���;�+�pM�躤���f[�]���LB�vu�D�_f!X�j���>��VrٓʹO��������O�=~c���<x��"C}B��kUG�j�UU��7$��5�0�I���!�>AI��%s�f4h�B%��5�$���_�Ä!V�}Q�j�����;��ک$W�y(�T!������D���jN��Ðtz���J<J8�=��!S�U�в��!6�*���d�nq2nlq8��c�]:�8����y�=?L59t$�6ٜh2���r��I���h��T�v�C��FQtt��'��V�j�r/����dc"�?�������K��||�郳e�7�S:���h6&$��{�j�zQ�јp8x�ȶhO�R��N�s#7G5�$�$4	*�,õYf���G��V�f���BW�=˭4���r��ɲ���M=F��q��"Ӊ�8Ǝ��Q�hŴ�F4ŵ�hĶ5�b-�-��1mbڴ�z�N�&'�������5��m1"b1��=c�����bb1֭�cV����ܘ�zƟ���=Lz�i1#���c�bc�J��|d�<Q�Z��}��+�Z��Kkli��ܘ��=y�~1��Ƌ>'Ĳ|X�<���%���BG�p(υ�D��,��GÁ�M��Ʊ*�k�OY��FK++��[_��'����j&&4�&5��bbc��F'���1m9�5�1��~O�0����O
<<R3��'��<�M~�xwO����ycF/�6��O��2?4��q��/�nAks��.eu�hfi��=i��oyˋq�tkNuye9|�-/ڇ��F���M;���v���'����+�{n^�v��W��{��[r�jc�z�w��jVƻ���N�7*ٺ�x}k��N�n��fz���l��xP��1�6���Z)���tr�_�}�-�]#�v���/9޾���}�9���ř�fT#>q�9���rY��Q0cM��jG=�6�n��-��I���c���ᨇ ��+u6�uȭq�,T���«
Gc!P��7r+�=�,�u��?'��K�~+J�����{���W�ҷ~��{����U�i[�]߽�{�v�ڴ�߮��鳥�t���O<'�������4h��#sUx]�I��HV4��V�mV�7]��48��e�Ѷ��*�9�#���2�G�O��UT+u���cH'jc��'(��%q:���QH"�ۭ��$*��FZ[��#��]�j'J$��@jT%Q�II]����++�u:�H�u���A^Ea>����*m�H��Z�P"c�ƥ�D��\mDX�WYu6AE>-H )�2AH�M�E-�B'SuأQT�6:�u��AVT��**�v�XYr�X��%j+cEÍ�N"Xېj&ܖ}[��d1n*0�3�.7sI2�nū!%8M&�iu�x\�2*�)H�q���?���[L��!ER�6�pe�8�P*NJ�V�ȗ��Iw������;9��mֶs�3���g&�}'��ڞZG�sy�2�����Ӫcws���s���QF.��U9��y�ݨ}���w��F���66��T|~LN!�(OC�N�|UC ��R�D�T��h���Gv��pɃ�錙Ff,��2}���2ͰJ��UQ�UL���b'��CD�$���'qV���w}�F&���^g�R���;7���A��s�#�kY$�x����>u�>qlbض1�N��?/;'<��%o�=��ϭ!�D�f��UZHt�nIS(��ي�8�M�h�>��I�RlL��v�WJ1Ew��9Okﲬ0�P��P���&&�a�b'��{�2j�}��m�Q���OIh�vY��w0��ð�z`�<Q�VQs'�CP�6�B���C�BC(�{qSG�~���#�_8��c�c�X�]:�8�C����oe�o���$,}X�J?;FQ�*ą�՝f�M&T��\,��p�lwNIHM+B*�>QD/�PZDH�]Q���C휜9�gs&����;�;�L�NLBı9�la�������B���l��H��tPJw[,��ㆍ��1����+�37?q���[|�1lq�uӮ������d��T-j�.����@���m�Qu��}�7v���0���Ѵ�ć5ؼc�K���㇫�r8k�p�"h��>62�!��LA=9�Mh�==��	�kRsE	��j	g!�R}�F�P�{�j4%�Æag0'o��Sm<N��[+o�-o�8��-�>>:t:t�Q�j��y/���n��I�'�o^�<{���$��!)I!�`�3�UUi!ϻ�=�����?m|��ӍV9ï7����q����w.���5Yo^��Gw�k|��M��3N5�v��4�\S�\��1�]����s�����h{�V�l�/���>���Ƹ\ ���k���,���T2���>�rd��p��u�`�Ksp�0�x%%��-J��Yw{�3C3#E��(O�E�]�%��ù�Z0w�C�"p�>7�h��Fl�8k^����n즕�>Ҩ��gq�/RTl؜2ӶR�2�u�����K�V�Ԍz��|�_8��[::C���<�Q�R�f1��L2����@Л�T֪����nF/]V�E�ȝ��UT0j�:����l�EY̗�����A״���غm�#ڮ�MĄ����d!,�q�K���q[M�>7�f>,A���ff
7�4\�1�\�B3��?SL[��|��-�[ź��Hp���sӺr�"kZ��*������z}��o�N��E�!���g��0��j����6'aA��!9��ƣ�e���7^�6����o�}��K7���&M&#�I����+atM�z�h�~>Xޮ.��6	����]�Ϩ�=FS>�4`D�C%C3&}p.�K�ILOړU�״��q��&1ű�c�ӡӤ8l��Yd���IJ�UU��Q�5U�9W����ޢώn�>9E��L,�o_pԞ��H���I�Zۑ�.�xʮ�g+F���,�ۄ�|OpH@�C��ȘC�ы,�%	���UZ��7�CS�;9FNf�9�F�C�"Y���e4$>�K.��w[*���̛63�/��3מ�z�1�c�c�-�WR����5%�5�~�*7l��@�1P Y�Y$�&u3*��U�?6�m����"���ɜ�}cŞ[wxt�s��Kx�]�1r=����K�l٘���^�t;�^qrw��J�1b�r>b�e��մ9!5�Tƭ���&but@,O��u,�*	Eyh�6|G��G�e땅�5�t����S�33&��i�%4�;���QWG��(O�3d�U��f�߇�L	�%�V���ɑ0h����L���:|�!�|�p�# ���Ե����15��8zh�4{%	P����5�V��7����=���~c�_8��[�]u�u�~֠�W��($�	���UZHv�s�j��e��9t�܈���`�'`am*�3��!f��bQb|m�@��X�U�V�^=]9w����B��a�'Ol�mU�w<�/�Q��I�m�ӏZx��Ϻ�����jW(��Ш0�c����]U�r̙2};Æ{5�|��~b�ckqn-պ�D�0L�0D�0���P���:hA�6"X��tE�6&�؛4&� ���0L(N�D�"lDN�&�,M�f����ؚ��vO���P �X�b%�ki�c��=E�q����:�㦏$b"pD�8"&8X�l�AL �%	�?���|?&�sy�ƞ�G�]�����ۗ�"��<��ߞ�4��y��N5ә�u��o"�>��j�J��ߧ9����y�3Ӝ�������!�r�s�꽐&����]�����,��֩Ź$�W�=��^��&��5�Sӎ�m��*��ފ��}�{���o��������mZV�~����{�ګj�[��߽�{���[U��߮��{����ڮ��~�߳=��یu�1�c뮺�D��f����$#�=��k55m��8�eJ��3���z��vYj�MQtk�ǘ��9F���C@�!f�^y�/��"}C�<%6;�������q�����M�CSY2!S�"�,4|p���^$�2&�f>>����6sj��!�x�f".S��]��>�t�m��q�V��c㮺���u��(��5"̶C{⪫I	��}62��
�˿ɲÀ�*�"J,D���>���q�qV⋫�[n�Y������Dxo%	�2��a�F~C4n��}l���Qh�*�f`�5�EP��Fx��W��k55�����x�C[�a�P�G{S��Ѝ�`˥����U�P�P��g~�LB�.�Ÿ��1���[��u�t��_C��6;�ϻ�c��}���ky�n�Qu�Ƹ��ۏ9��e��.Bc�X�^����Cgw�Ͼ�xO�,�����o��n�]��O'9�ܝޙ�έ|��q����=������L|l�+�����Z���FԜ�/��_Wj�/=w|ӛM�f��fQ��i���o˒�6���j���s$�]>���:&�;>(	���D��MU`�ri� ȉ���`�����]�}5��>��6"����a����Ĵ�E����r�Q���OXl����T��l��kZ�ߟ�?1m��1����Ν:C�p�ɰ�Kn+ 2������2�:r}G����p�d;�r��Q�xHY���B�(Ѽl�%��c��2&6�����k*�Ap��8+���3�ϴ���9%ҋ;ϔ�)�B&%���0�ĥ����dnO��_�ef5.>.��(�6d�6��]no��=��(�*F�!�4X�F��F�3�k_k�~�8���c���-�[n�:C�p؅��N�V��z�����w�&����$8gUE:�$ȗ��pѢ�P���5���ɓb(����z���tW�ǅ��Ʉ8e9��ѕ���4;2|��N�f!S�^2&�v\,�]�>����X�܈�i�i�+�d�n7����'F9k�J*~ϝ�_��{O\~|�|��1�c4p��8Q�|�f���Shy��s���$;G�ԁ��%}F���Hq�����������<`��t��-r���v~�RfU����+��#�ھ�����kG'��97f!�C����A�0������M��H�I�X~A9[?Qt~;���8����W���Օ�֛m���6���x�a��/[���i�����j(=�H���uJ#��6H�F��n�G��UV��w��u����y	'x�׶/f�^��ӫ����>(d���9�ݾ��Ũ��'���ɩ��;nr��a
�^���i�4L���^w�s��wA�ӃO�ӟ'Ϸ��l�Y�%��OMC&�����2i6 �!��>��L�br!eo�j���]/�J,n��9)7v˗VssuK8xl�0Pb'��QF�t�i(�R%]Ye�3<b}�f7cǎ�&������4���^>Z�cn��[��]ui�*�\%$*J޺��Н�E�t5���5A�!Sf�(�=g�� �/��3����wwk����7��9>����P��O����Q}��~�	%Ed,���pXG,��j�k�G��@�	Ҍ.�a���Y�w��1(�ܔ|}��O�,bR�S�m��u��m�>b�ſ:t���6�`��ْ�V�⪫Bl�=�UZ:&���>W���4%'h�t��+�ȜM�OQ�u�U�
�`a�S~��N�Ӈ�pOq�B��fO�e*�[�U��}�G�C��B���2bD�)����OԺ��)�z��ͱ�X�-�[�]ui��\Ԓ��U!#!�n-ꪫBrU5 C�7�Q�ɟk���ZC�a�;�O04|��̱Z�\��I-��ߚs�M/�x�`��P�z�P�D��Q��4��CA�4j}܇Œq6<���8�ۍ�~����:h��ϸ�h׌cWG+��԰��7�ᰇǫ�I�ɺ8f+*�p��8t���hɂ�2||d����pN��0�0L�tDH"&��"A6��:hA�6'DL4"&"lM	�6hMFH��:"C�� ��0D���`��؛4%�f͉�(J'd�>A����b'�Q�D��6x�u�1���ձ׌1��1�Ǆ���pDL7�X�h�AA(�K<`zNQ=��V>�x�k��s���8��)��YO�f<�[s6BM9^Κ�.v�NM�:.�GԳ�2����_����cfsw��>jq�^\?5t������k:�wdWs"ڰ��s���o�9ܡ�=��C��ܗ���:L�1P'wwDoF��澬��˹һ;}W-�1��ޝ�����L^����������o9�Nf3��_��/9��ȏ}��<5�����rm\3�m5=֡]$$W�b�"�F�nTՊ_�+�;o���hu�8�UG��Ym�N�����6�M��B��;h�n�[#��D;ћ�]T�s�}Wj�[���~���{޵]��n�~�{����Z��t�w�_��{���Wj�ۻ�_�gN8p����x���8[�j��j���]�������Dr���
�ea��'Y���H����F�2H1FJ�Uq6ȕT�ҵU�n��\�U��(ₑ�X����H�%��l8�,R_�uD_��(�+��B�-'���J�>��Ui#ER���Gm��2�jImm���i��r|�cn��u���G	U���(�p(K-�}i�R5�K,-�4[Q�݃�mZDAZZ��$�#r�*&�jX���F�C!�%�r?�S"��l�A�����,�wf�����T[�,�7�-ɋ�4:�Y��&R��p�O�޶�m��U��~����~��{��735j�����z�w�v��Hu�P{n���;p]{�f��������U���:��{	�^[��'r����wP�uy���"���_l��㜘�0�gǍK�.����Ї�������ʡ+#��b�ʢ�x�tV�;U��ij��#՗^�=~_���ʇ/y�N�j�{��	��^Dԑc�����!��в�(;��"{�(���6�n�l[����:Ӌk�d�QL\�%
=�}�r�rS�UV�0�M�g	e�,f��2��QB�(	��w~��ǆ��+��� [O|B?I����O������Cg�(�|�Ji�8�۩]Ѧ+��.�\qb`@�6G	�[p�ild�'����j<T(���q�a��C�P�ڨ�ʓ�m�F:��co�������:C�p���r�O7�UV�sO�m�3/.�/;DM�ߤT������oMSm㕺�G���)�|1T�r9R�Pa��϶����2j浬�2��t�c�X'+���3d̰K@ɒ���C�!�,���Ua��]��˽oZ��3Zӷ���_[���Zej�!�z��|�ͱn-n��[�]ui���EA2˅6X��c]*��&������FY�PY�v�j��Kݍ��ʨb��Dd�E�<p.C�CQ<T�f	�3��2\������}F�U�M_z��q��6j�U=ArrL���x���h3C��}�[�i��o�7L���׮?:�ͱ����:h�aGB�OzJֵ���zk7]̃���D]�tϊc����]�~�ʪ�	�����f�r��Zf�ܯ��ϳ����m�u�u�d����n�Yǿ���3��ꄻ�P�^�rc�C�������1�t=�vf���>儚,�^o�s��p���3c��1&St�r�ӑ0�NR���=�t��[�,���0\���,�NW޿�qMQtO����p�(&��eOC�>�!g�E�Rl�鹐ف�J�a�2�0[+woj���/������#J��j<y�km���6�1n��[�uiƫ^O$���y(2�V�J��	6X�(��ჳ�5�B�92ve�s;I����=�\fa�^����}(U����e�w���}��̺�Ys�4t�z����s��k�x���/Ux��V���>>6@�+��j��e~i����c�-n��[�.��u5��ߏ�I�1�	���ު��'5$�R	��h��������_������ݍ�&�eM��>*f�27iO��.�a�(�Y1��	F��OIɐOósP�>���;��US?�v!�s���`Q�!^�.캺-�pى����D�zY֏)�=r����O��ϛ[�>[�|Ÿ��Q֜krm��ĸْI[$7�*��$��՚,�V�W)��4c�j�>��>���n�ί�2�s�?={��%��&fb�s��`�������He�����g����v�13�����}p�0�]gY��kWe��}GL Ci�çG1�6t�Y�eT3���5��i���Ri�u�<�>q�ͱ�&	��tц�����\�ܛ���"���&�L�.��F���r�t�]��3#[�y|m�|��М��i��w���6O��U:��c��7�.�|⦭�;�7������,s\gp]�Ъg/M������S��}����Y�t�{�gKf��2���yU����}k7�^۷v���c��*bn}"vzt��{N	[��~zh�d�<�FG2�h��|j��֊�����}��6�G�p8eW��eUp�a�B�\���hꈜ�K��'�56x���Ѫ]�<Pd٣I�ʫm|˪-��K��zC"c�d����������Ŷ����Ÿ��Q֜������VBcT�Yo7�UV��~�XxЙf���]'���Ǭ�j`U3�&�Q{P�g���k;8$̒�w�,��t���LM����e|J��I��lo�k��]��t���v����ej�.�1�FfϬ5 �w�8��t�'A?z�8F~��qź���m��N,�&	�`�&	�`���ΉӅ�����pHhA(M�"'D��blM�D ���:P��H"&�8"`���,M��L�IBt�����萀�	ki��[m-Ÿ�սzǌ-�u�z�1kun4�֋Z���1�Ǆ��0L8h�,�B � �"QBg35��go��\d�M/������r��M����{��;��w���oŪ�rC�7;VL�د^�����˼>�p�a/���
Sˋ^��{ս�n�;��_w)�s���ߺ���\�%G���υ�Ź��+�9����Ű����'+7ׯåWm����{����q]*�n���z��{����:Uv�������{��եWm����YӇN�8p�㧄�<x��Ν!��⪫F�5'�&f6�^4J;7՟�摛ڪ� �!�h���0nL��&�|�(1�^�c)B>?72[2��=�����O�k�G�ӟr��NK�����.�w�CA�8|�كS0��ٳA��U:�mhѩ����G3E�>���2̘.|�~~G��]b�b�|�V�-ǎ���$�:4v��J2�gy�UV�Ȑ�E��.�'2#�P؆~}A���6�I���t?eH����|�2lp3�4Pf&�4���A�2�ˡa���+�{�鲃Pٓ���������}���9�k�sm��c����G^�$�r|��2���z�����(�����TM��bf����>m�q��[�-ǎ��� 筃/�$ƶ]*ݙ%l�"$�Z8�M�ϭ�$�nq��m�����C^.*D����~�-��&>��Fw{�Nm��?����V�h�^�t�V|s�L�~��槻^�I��G[3�>�{��{tX��e�O�_���?h�f�P�f��O~�#F��#�����,���(���13
���@����84cr�������*�>��;{*��\��J�&2\����HdԹ�Q.�"��뱇����T��ȗu|&Z˿ձ�	����ׯ[km�\b�[�:�:�$�xE��2倣�!v�;�*���(��E�N�U�ȁ�}`��fL�jPfr�M2��R����ȷ�*�eM��C���,�oh, ���>~>>�L|-���Sa����m��Egn1wwue[=��˨s�j�XYً����p�Gg#�nab�W^>|��|�lu�-ձ�q㮡��ۋ#����%f�UZ=J��Ð��oh�F�d�45��g�>���A���s�o^����g{���ȟ��퍥�mbk
���3�2�|��K�J�LL�5��4�8l/�g��}�g:�]z�fe�w�4k]��2�h7h��[Y���2����u�1���[�c8YӤ:<��+���P.k���ͻ��j���|����W6^��k�On�S8��U�f&��gy7��h7�;����1��I-�uC�%t{͆��&�w��nP]��tc�-�j�h���5ᗇ��;K~�6�b�6������1n<u�u�/!��v`\ܱ=�&�z�+�/�q�M�9����X�`�ې)U�m���ӛ�^x��׍2�uM�v�{�f��>�y�"�,Ƿdi�.-�jùdÔ�9������Cw�u5��:�����;��v�rn�N<Ң��~>�7�/(�WK�b��88�d�p�ݜ�gC�R3>|uV2*��h��9�2Y^���xfv1��:��{��p�>��.��r�͟CP�C��ʪ�J*��UdVB2O��.���t,�t�,]�1li�1�kuŭվb�x�:<�_��߱̈�⪫D���7�.d�Tu��7�p=`G{6V���C%�ǻ��e�*����;�;�E��OR�<��C�<fnt>��#���ʵ�֊~mU�+�f��{���%Wq���%þ!�Cг0�Wª�t϶5�����u�c|�V�-ǎ��G�k�;.��̘�6�e�L.���UUZ/�����G[��玚!���i���Cq��2��oWzfMCQ
��Ս\�z��.�WKB_�QL��V��(�����G�:~~��1��u��8r�u��2�4p�	fwcI$��8��[�Ao(�6���!�sTr�G�����Ξ8x�çǎ�,��8V���SIJ�r����?K!��]W(�~�]w7���s|eۺ�ݸm�zVk9�3�����s�W�M0��S��9\��0��9�$?gh�r�q~uw}F��MB�1�G��C3�������[���4zh���9�p�c'��e{��C���׵��]m���c�x㍭�tL��&	�tL0�,��%"lDDDN�%DJB"p�:""tN	��X�l٢� ��Ȉ��p�H'DK4"pD�0N	blM�6P�;dM��ԟ �
IE"%	b'
�p�Bl�G�0�<x�ǄL�"A6"%��X�1�6��c�M0��, ��Bh��sO�����/��UL��|���qa��Z||�DѺl������s�/{�؁�������C�Of4��_n�ºth�����G�{�'�Ys�7���j³;��]�k���b�,���ޝg\��('�my�q��j�^O��n)��yܠ�zq��d̜h�6��Ν�R�������7W��:�^�=��1�ofׇ)�d�*�oMǝ�G9�/a��e�Sox�u����I��)�Ϸ�s��޴��Z��3-�8�S"��ԣ�V얐���R�ۅ�%��̑�&|P�I"n�2����8�>*pr�+	�8������y8s>����L�rs���J�ۻ����{����uiU�ww�ǽ�{���եWm���{����{�ZU[����l�g<p�㧄��t��uqE�2�G#$-n�+��(��~vB?�N��+a�v�F줣�Kk�D�>��G�|J�EU?��u9- �"DM�-U��+RDZ���7�V5iI�B|�w��V��*�q��P��k�%+��dڄmDӨ�X����X�r��*b�ђ�4�m��'\�K[
�ʲZ��deN:Q��Y(�r1B��m@A~���D���X��[>�b�3�譥��ϥv i�K�vW'�
�l����-R��2��t#�$�5dj8�c�AYYW3ō�+p����mV)A5�t���F�$14;%�(H�6�U��&F+c�.۲`�ȋ�	`��������#�֪�F{��m�g߭��/zssw��\w�����ʮp�*�|w�;��X����z��]�Cd��\*����L�s/ڵI"���=��=���n�Meg��`�4^ʤ��f����ds.f�c$`��{�T�m7�"lm�Y�2�1*s�á��u��n@��ȚF��v_��rc�:�Vg�������SV��^�X��Oϟ�u�V�����G]G\x�[��e�LU.aj�Y�U��ؗJ�3�5_�=�������LcH�u�c���+��zjn����'zL.��C�VàinJ��h��l�EX��U���Q?��	
���ͪ.O�@���El�8p���s���H�m�~Z�m����������8l�\｜b�~�H�U��UXv�T��M�(��nWP�Ý��+���x�S�O0�2�5�Ғ@Ţ���\�^K�\�L�w���y{왆(�=9�=�3�]���
�a��O@��#����ג�o��%���� �M �=�=>�h2p�o�q�1ŭխ�8�����?F�RනBQ�*�,��&B�3��^ߒjO@@AN��$�eŘ�)/(���}|.v���2|(ޡ��3���(��ؚ�b�0
UV�e-���j�Y�w4��B�#�"���a+��˙�U���96��i�v�)t�]c�սm�ku�-լ��8pN,�<g��R�F
J�\��Z�q��-L+�,� |�s�����jr����������]����g8H��^n�1���8e+�R�Je�Gm�ܱu���(��*8��^)�x��1v$Y7]ջ�p���\�qlr4h����<�f���c�Mr8)���rB�g_UE��˒�����y�'���Q��_�OՆ��Y����骱�,��fYY�|1h��b_Yf7���um���>[�[��G]G[,͚�j�m�Baƶ����ـ�fa��¥G���~��wwEU�|���z�a�������0vÐ�6bYB}���8nG�����8��m�]�~m�22����{�_�BU۩)M%�Od�������=DG�~!���-�9�箺�m�c�t�ӧ���z�SS*��˽*�7�L+UB�}S'�a���i����kKP��w&�a��8e~�r���C��|~�6_W�L�-�^�X�M�U����ǵ'B�\�(2NA���rMfCX�0m]I���iV'|v��j����^���0�o��ŶŸ������Q�9����8E�C��|���G�-��������X�����~�}�{Z�r�ӫK���#���v��
���R�<��hۦ�9$NSOijCT{�v�~x"�"V�~�� ��7�l�c��૦$�*�E��S!���I�*�p�&����<z�6�n-n�n�quqE�4s1T*S��@q�]�p4SX�ݺ��MS,owb�l�B��B��#{� ��~�s���ܩ�����p��:����δE��繽=�~��5���Q��(�^��<4����}��_.b�8��y��-j��p��o�erb�~'��Y���=1�eK�T�E1,Ĩ!p���͛��n�Ǖɇbص�qG*��]n�{Azܐ{{�ѥ��G�Wժ���p&o��Tn��4l����n�n��u�uǌ���m�U*�����=ɘY�O����ziafC���7t�U]��R��,=2`���_l>�U_I�p��`Εsf'O��A�=��U\b��JO7t�SiW���'C�&�T�;	U��J���w^�W�i˧�W���8�z�m�a��8���&	�`�&	�"&��"!B&�DD�:AM�"lDK:"`���؛,�I�"A�DL�"5"#rA��,KblКd�(J,�C�I�X'�AH�:W$���cK8�1�c���'
DJ�N��"`�<m���Ѧa�YkE���QL���V�ғ{NM���y�Y���:f�-���^׶i+�����lȩ��P��9�{��m��sxs�Q]��m�x߸��Eʽ`���2k�b�}�_gj�8�q��rκh�2��}��٫��ݠ<���-�=zM��b���N�g7�{�ַ9�Y�����_�:�=�#ϳ���Q��ߌ����U���_{����{��U���_{����{��U���_{����{��U���|l�g<p�㧄�:p�8pN,�1�U���P�V*l�o������T�B��}4^�*��f��vv;�o�=���30h97av���I�yvg
�5��T53��}��E79���`;�郐�l=U���_G3&*�^r����z�tl}�ZG]b�m�qkuku�#����t����ꃹߑwCauXz�ט�_r���7ź�ﯶ-��u���K�hˏ*WO��E�n����j��bD�0�3���&�����fדv�'·�~�vfLɄ�)3��7�~�we�pkJ�WC�<�VT�8�x�����ط�V�_8���]\Q~W���Ñƍ��3"�|µ���(Ќ.Sw.6�Z�ϙ�<R��W�>��[��s_{%{�ֳ?)�����׳ՙU�糦UoS8���sz���z��<s���3�7�5�o��JI�oC�h�d�r]ct?vs�]s-��Skhް�7|~�Z�&�ѓ��l>>f0x҈���r�x�nn��i��W�*װ��WPg!FM�Æ��r	��p7t����G�p�<��*Ki}u~��U�-��p�j�2O������W��z��'9M-�ۍ�돖�ӧ��Âp�g�zj��EmUa�DY�a��0`52�ޮ�tU)uq�}Ȗ���MBQ�Q��{�RG�VF2p����
�(9��Qi�*�������J�V�F&W�2/��sx;*fYea�����"09�@[�O�GejK�7��>�r�ׯ��ێ�������Q�;�T֪������I$�ܕ�Y���>�9U���x�X�4WmL*l��d4p�'���{�7���^r-�h��K�N��G<b�F'
���zdE�,�M�vg���eS^۬a�]cQN�S���:����u�i�[�?:���-n�n�quq�y�?My'��jvT�UȪ�4 >ߚ���U����9�����̛���+w��J�c���I��&�]8|z��D�ڪf��\��Mc��Ƀ����6\9��2|Tf�Y�{'%������a�EoP_��6\
f;�ۯ+���kn��c�-�V�����Ht�>�U��s��VoeB�e�9UC��K>x��l�n�2,4�U�$��V"4|� ������߯���>v��=��Θy�����pM��=�`�o5�;�{����x���p/=��L�n�w6J�K�qՒ�]�F�z�;^�X�T����[��,-�����G��{P�x���VUl�v�I�ly�]�rXm�5e"%r	ٹ��L�9�c�t0��c��}VW*���zx�y��:��n�~��7�۬���8�@�%�D�T|'M���i�"I/��v�~m�፾|�康�8lM�,����p�����`���Pkk��,�tg�)�j�߻��r|����{,ٙ�s%�5UTqQ{�0�����TK�BՑ��+cN��2u�үN��>��zJQx>����Gxh�W�a�k��̹~x��H���8���[�qo���٢��{)!�K��P�8hd��Ix�YΊ�k��V�VSR�`e����.\�wf��FC��x��fQ��d0���!'	ܶ�����,�\�y�Js�y�����f	�x���T��.b���Cr�C�nh�����St�u{^�LWV�n�m�-��㧎>�!�e���[ �)�r����`�{��l�̣�ˣ�0{�~n]��U�T����pĖm�%P�62�wM�JJ,	K��bN��att�G�:��$�$�5\�p:Q�����ˆN8]d4M��.����?Yܒ$"I�$�$�I�*�4Q󽏬�C�5��ނOhq�ر8PPQ��!���v���_Bͮ�f"�(2*�(!āPHČ�0A��Ĩ$�A�(1	 �$b�`��1#1#�b0H�$b�""2%(`���A�H�$`� ���I""D�b�`��1 ��$`��`�b"�A�F"�� �b ��H�"�!$dA�B  �D �!"#�A���0A"bA�H�"$$bH��`�`�`�b"0H�$�F#�DI����0ADF"�� ��`����Db"1�ă0D�"1H0A� �DF �"#���DQ�DF �1F$"�"##A#"0F1 �Db"0H�!�#Db"1Ȍ���A"�	%0DF" �"$��"$���"� �F���"	��DD`����F�����$�#�2#�"#��Ȉ"$"#DDb""0DH1"#A""#D)$��""0DDF	�"#""" $DF�Ȉ��#""0DDF�D�#�""0DF$�dDF��$b ���1 �Č����F	DF$`�#D`�`���A�"1!I%1�F0F" �D#D"#Db`��F$ 1"#����1�Db0DF ��A�#D���DH1F�$DE*)D�DE!�V�H!H%U �TT�QPE* F`Q�HT�)PJ��R��R��*@"��-�� �?�!U���U*  0�Av`��-� 0�U�%UJ� �J!D�������B��R	T��A �*	UDJ�)�Ĩ-"� �� @!JAUUA)PEJi
�D��R�*���DXV�D��	EAH"�U ���"�U ��B�EJT��� �H"�!H"� AP@�R�� �H%UA(A)P%QQ*��JTD � `� �2D	D#� � �
�P1A��c%2�J�5H"����!
��BR	HD%!JB HT�$% �B�B�B JAJ�!)BT!�J�D"�JB! � Ȃ! ��2 ���JAT�B��D%T"��D*R!JB!�P�J�B�DD"�"w`%T"	P�D% �%B����J�B!)B2 �2 �2 �"A�P��!	HD"��FDdA`�1A�B2 �"	HB��*R��!A�A�0B �A�A�A�B0B��BUB!*��JB�	HB�	U�aI)�A�`�0AD��"�(DDDȂ ȁ�"��
�JB!*	HD%T�T�!�"���J@�	P�%B!*BB*�	P�%B�HB��%!��BT�����T"*�	P�% �����B��JB���HB��J�!*��@��BT!	HD%BT)*	BT*@�H� 1A�AA� ĈEA�P���%!JAT�!	H!	HD��PD"�J�BT"�"��J�����R)BT	P�	HJ�BR�T"�D%B ���D	P�%B ��RT	
�
J@�ʔP!!D## ���0@`��0B0B��GQF	��%!R�%!IPJ@��J@��JA*�������DD�`�`��!!!!a��F!!�x5z�`$`F!��`�b
 ��"$	��bH� ����F	���0A�$�F#��$JDD�%!)��B��e��ŋ��H�9
�}�8lAI E#Pd� Ć�I:>��k���N{O��M�=�hZ�T��<�Wݞa_�������[�0e���B�9�� P�����N:�?N7��'�o~�y�s�п��~7Għ�g�?���
��C�ͮ� x�����S�DO�`�@E(�@��~Q9��`��ww~C �D�NV_�	����;�A����\;�<!�**���'�z�?,	 J�4R�ۚQ���n�ye�$Y�ޚ!��bRR|���x+M]�Κ�!��<a��Ýλ!��K1��~���m��*�!\�X����Y,#H��A��*!���*h*�H�"(� �}-3N5��M�=V2q߂c��G����AT�5�R�(
�`F�� (+ B�� (��Q�����`�&GW�3���:�]4�zGn �G "��x���R>������� @PN��։d:Z����_j���wR??���~A�]��/�>���d(�7p7"�È�n����s~���<M�'P��@zG�	���Y�ܯ����p>�|B	�y���"�����P"��ٟ�����lo��8MC��75	��Z2���TD���7�,��#�6v�(4��d�d�*aC]��I)(��Jh{2�Y����V6#h7,���K��Mb��QU@iLմ������wh�eQT����Ђ�Jt�z�*�������:������2Y"��:�S�}	��#����3�r@�)����bl�t���<�WC�PRz�����j��@t����x���9���r>1��8�~!�=%���A��B��;F�nK�(�7;j��<$�˰�q �-����X=L�[��7p۰p�����҇48��2�v/C�c�(l}��=#�>~�!��n���^�H�K�aF�����.@yq^�EA?�+����4 �Q��r9N�sUA:��mt���r���):��N��>yz����;qM?����ܑN$�q�@