BZh91AY&SYs����߀py����߰����a�      CF�   ����@�Z(�Y%A�mm( gf �@P m�������`�      P   ��  <֫g���]�=��e{�v۫]v釪{�{��=v�7�y�v��,z��i���z��W����zӅ:��m=7�:��3@f�����r�(6w  많�^벜]\��)����;Ǟ^�w�yV�q6륢Ξ����w;���J�9��l�j��͞��M�9���m�uÝ�j��rwwm���v��C��PF� >�{նz�2�u͜�������s�g[�[v��Y��n�ww-x8F���Sk+\�j��n�����3�[�l��ۺ�;�s���z g` ��vl�ڷr�w;�#�.�k��nunwt�q���]�vׁ������]�g^��^���]ۮ���k+\�]ݹu+������ ������{k���a��{�r���k��x��ݾ��xm}建k���4�^�u�nn��YtK�R׽��@                 *	$  �         @P%S�4�R�H 0&�`di���%0��UMQ�F	�  i�0 Sj IT��0  FFi�  MR$M=R2L�0�� `A���5R�L@h	��iO�D=�~�PMD��T�2Ɉ 20������e7
�r�-?h����;a�� �����PAڀ�~B"?�_���X �i�����?�����������}��'�9?�G�B ?��@in���J�P�$����?8/H�
�����@PM�>���1��������?�6M)�'�c�ӌBKz[�4K���1L���4^�&�jͺ�K�ܘ�ܓ���d����Y�y ��/�$4�;g)���d��'0�d���N�/��6$d�!h��I<4];7'��i��8�!�g�l���ɴ�IZH��P���"t�w�%&����u!ߓ��':�GR��J1��"ȝ)�"WG�);�w�>Mٌ%�:�,w�pp�� �a,H�&�&��d�F��丑�H�9�P�ԝ8u�>�͒��7�r�"/	E��%j�J����&'Rt�ݒ�P��D��DLN�&bV�"R"=,�Q"'6���QpKDN��9��ȑ4;�N��"Z'N�'�LM���$D�Iâq�8Y���3��Ei"%q"%a�h���������	pDٚH�9�P������S
�H�ԟ'bK4;��8$DN�|!C��%��$N�N��M����u(R��f��8�e��G�4C�h���:"RW�8F�f�M�+�	։P�!>��>h��D�tS��H�7GN'L��&�A���IF��"<ʉ��8�+�����L��s���������:q�S!tA�F����7���a!��6�ؔ��g>����:�`�f�4V����;�:�<!߳��N�pY��uR�V�%Օ7��E��q12�Q��Sh�J�G�?X�&��F"#˨�p����E$�8M�(&�7/b#��pཀྵ��~�K4�g�T�'��p��+i�50�M����{�S吿���[�*#��JK*�U$42^�]��W;��D��0���"<��&5>L��$Dr"q��P?m��pA��6[4Y�.DG������"5���bP��V�s�G5Q�"ev�t�j|�UDL�b7���Ħ�l��"8H���@���u�0Ќ�,MjM��Jrp��������'(��DG��������DG�Q�ja���N�O��f�܈��Q�S��>MA�TD{uGNH��S��mO�$����Dyʈ�ʉºM]O�wU���ߞ��CmN�+�&5R�	�r�#��2|�UD��*&��Ѧ�K*ڟ,�����Į�r������D�5,N�ә8o�H2d��	y+<�y����k�G�	ѓbx~�s|(L�s�e��\��hѡ�s
Ћ���,�����M�,F�QC�ȉ�58_f�u�gݣP�J� �mO��
�A:I!��d;#�=�vC}����9{0��{��<�<�D��n��t�0jpF�S/�elG|��5̴��%"QӬ�&+2��42Q.s�O�ϖV��pu6L2X�c�C^f�|�ޤ�����^a��sL��ʶT=r������+ǲ'�,�e�I,��,�l���։�Y��=ͳ���~�=�<�7&#�lk�}��ލi�խ�֭����D�U���=J����d��;�J�j�������*n%Nm(��]E�v�\���C����tԻ��ޣ��ɪ�c̩�g�����rw��:�77�f�|k�Z�ԃ�_P�<�#�9��.MH���q�n9�_Q���7�R�S|�پ5�'�&UN�\��ު���Q�yʏ"f�*\j]K�K��Mi�d{>{&UJ��W%GrdoU�r�Ɇm��9�P�&kU/%g*�:��:Ha!�98oSU�N�v�v{�['�/�f٩2ON�����\�E&���鈎�%�#"sf�%	�dх8W�!8D�%g*P�$y�������Y�4q/\��C�`����WbQ�tj"c�H�������r�A�4&��%"v��1��벾~�U�D�8�I6A�Dy-epя�,u�_#؎M�_D��Dy�_#�&��H�"#����T���r�8�R"�W���Б�H�c0��D�g̲��6�R#�(y���5)N�"&H�����\��r?=��j�*���H�YI�ze}_;���%"s��4u�t��J��eY�O�]8ܭ	�r�Gu���5)N�"q�".�t��%|��Mf�X�y)--e&�%}_;���%"s��4u�t�M	���'kr�O���,�H��Ioj�&��L��n�R��_bp�t�N���{�j_�+�0o%X��V6[8\��jDjl�"=�'f�&m��}��B���?9*	���i�(��DnlM�)��Έ�+���{+��5�����4:���{�IcR��ʬ���H�U&�	�+{$�t��[ Բ�F���ȝ+���J�F2H#ߦT����~錃�K�ʐu!ϑ샟Lə����مMdL��_��o�7�'!���z��<�q����F����c�M�јo�{�\�_j({Q}�ٯr9��=��,�񋻋��F����q�\Y\�+vJ�q���̹�ǲ�\��R�ԧs�Y����V�T����d��N;��g���j��9���h���%d�=5�{��e�[ئt�~W�SS���J�l玩95tMCF�I�T����y>]g��K��9��G;&l�K�6왣�;'4[�s�q:$�G��	fQ[
�Q"N��Hbw�0xS�kf�}%���3���A&���i���ę�+���)1��U����?J�����)��w�ʩ����2�g��XR��R��3�c��`�İ��p�����:��ʰOdjz��yŜA5��}9�-�w�C�|���~�F�$��*�D�f͟��ϵ��Y�u��r7	�N����of�#+k��Q5:=GE�j����9�^a�S���T\�m�ى��>��l��&���\<��>���W���TJyr;كS|M�eY��t�Z滦w����G�-������)d���Φ-�R�W*��}È:�v_S��|V��1�Y|���e����f���F;�T5P?�qd�|���o=�wbv��ͷ�ԙ������k����WVe9�N�_�{���8�G�N�����w��5��^�]��~Iv��?w��ԯe߹���5so�f��֣n��e���U�_��ܖ,��s��gy����~�Q�Y�Y�����sL��r֬��\�V_�v����i����|�':��>�w�y��w{�s��y�g5���}˪��UF.v�O���'Q�~��d���q-�����-���R9�-�;���<�,�Ս�<��.���_�r�-_(�_r}�y�^�N?o�<�|������^�H����u_���2��^��˽}]]�,��N*���ۼ�qD�{38�{=�Ns��G��q�������Ԛ�,���N��ݓy���1�NϤ�2��5�Vu�����m�\��i�Ӌ�+$? ���y?.$���3V��������3x��mT�8����I5��H����^\I%Qj���7{��OG{N�,7d���o��X�w�L��m�7��ө��QAU��~Uj��V~Yަ�I-��;y��.$��ݯ�������&�i*��qx�F����UR_]��Uũ�ME����y��$�_���z}K�����i/-]Ԭ�̩���90=�Mo��KN��U-A�������M�K6Rj.�f�휷��a��b����Iq���mf_p��J>#m F�4|�w�Y鮴B|뇮A�}�n�h�S��8 h�dl�o2Q���Y��i<��yg!������x���+���ʈ,�H�,ﴘ}�/�6%�<=�Ū�!�h��+���!6���:A�Vd�yϞgz8�p���N����L��*���8�	���"�������3Tc5o�a{h��4kg's������؄�93�	G�Yx��Y��X���>YU�m7m}���Z����nj0���f�];����s�n���j�oi���y<��ҵ	ֹ+�sMIZG��j>VcX,��x�D?p��5��P-yVs���B�4Gz��O�\��y5���2�^��'ad�!��%v��vo��t�4<K�I�D���������r�O���L�M��,�7�#ҬA8��V�;)������̆���D�O:\�ʐ��o�>�������n��ۏ���������j9e���9���v&\'�k��L��ס}k�%�׶;k�~M��Jej�Z�ֲ�ݵ�yM�f�*��,硯�������{p�������e0��h�pD}ƙU�v�v>�%w��JƎy~ֲw�?������ϴ��ʱ���WM�$Ȳ�i׍�ϧK垃�ĳ�8�*=B<:��>��͙�8�h���-Y ������9�R�+Q�*E�yn;��l}-d�V���X�&q�J�^<�,�uVr����t�ŝYV5��8�,�5f���Ȋ!�}[XE���"���q�<č�����>�4��>��4Q�����Ŗ�-���F�7�A����s��_p��X��p��S�n<�#�h��+����rWao�Y�Z�k�n�G��;�q�c��q��3��YŝG�ȱ,�>xn���+Nv�a�VM��js��V����Z>C��s6�Ƅ��:����:���Lk_-��E�Q���Y�漋�,�C�/�m����;&�s����	�{�>Gz�#N��D�)�4v���ϦM�DN<���o^r��h�Ƴ�*��
����5�;��cB�8�/Ɲ���������I���I��qa���VqeX�U��N ��^L�Ds��s�7>:��cD�Y>7�:Ǩ������g~�Y7��c�݇_3��H�c�)3�~�*�#�2�!�/�w�D�F.��ݹ�=�((�՞EG"9���=�ig��{T�ۜd�����g�?!�	��N<�s5db�5\�Nz�!I凑��,���2r��? ��:�}�8�P�ga6�Xw�Y�X�C\Mk���n�b&缚�g�=My�S+!zh��6��5�����?Q�4^U�O����=G�?#c;����.���lC,�:�_v��yG�^�q�ʎ|���CI���hU�YVU��|=�nTg_K��9�YZ��pw��C:���^A�L�A!�k��<5��J���yC?Sq�Y�b&#�����Q��Q:���V��y��65Vym�'��>i�TO'�W��e�~��|��u�Ǘ���+�ڮg~����[��Ԯd�f�4�����*��k_��]�)�_������1����W���Oʗ-�����Wت��٬����H�|M��ս�=[�V���y//���l�˗��%g9w�q��c�{����Moo��{{�ޭ�R��ʟz��N���N���vض��Ǽsds�ά�����p���󫳝��ux��۝��?o}�:l}�f�w������z���V��٩����N���^��h���p�^��������[�������{=��헼�Riio�s���z��5�'l����oD��Ӎ�ɽ|��+�_��{�s�d���^͝�.�5�M~�Cyۯ��W�U$���׻�i��w��j����j}���M�vy��)�a�ےˊo5?���9}���?%��<��M�y7g^�s��{98zz�7����~��e���K[���䜤��ƻH4�eG���M��n�����:#���Z��9H��>˾�Wb���m�|=d�{ϧ��~��_�/�h����?�ћ�*ͨ'-�qj�*F�ݒ��uc�YW��=�²!ן�^F%�H-qJ��R� Ғ��Ȫ�H����" "İK�[��2��-����1J���F܋5���C��\���W�v��W��d6C+|v8�,V[n[qV�Ҳ��ȒH��lQR�K>����j����Ȓ�"q�JnFD��D^Z�дr3�M�gcmj�]��,����ΧF��q��Z������j����&�ZK]�L�dL��u;\�ѷ0s9=974_����1HI�FI����w�qpE�	rAeydrB	��������J���e�����[1U {��������y��92���917�8ƍ��I�NmV�1=)%�W��*�,9*�96I��Q�iWZ+*Q@7a쒺��&��h�3����^l'#���&�,�2,�Ǜ����K[o�^�Y��Z#DJ�V��*eIe�Ⱥ����k�a�J��\-
8U�3UHז�,��Sj���et�	ɻ��X�DF͹J�z�wy1"lJ)�Ff�ԕ
E�z�31	z�$��t�I�n+�h��Ud��U�\<���8�A�W`-eF�@��aD�T�u��i���0�9�5**rh�"a��S�"T]D�8Mf�/�Pԑp�`d_xj���,�f򙛣��35�h.W3;�B{�<�g���)�+��+��\��;;x(*r;����<������p�*��P>u+���P��1L��E���̳��8�g�.X�U�R�5�j"��/6�T���b75�7Qy�G1�g[��ƿ�!�����_��� ���������?�^$-'�?��?���?3��~ � ��P��i$���o��,g_����w��j�j�Uv�ڮ�W�Uz����UW����J��WJ�j�UҪ�UqiUګjҪ���S�*��b���UU�*��*�UV�����U⮖�@H'��� HlԓfK7�x��Sr�4�ͨ(ՙ�����@���m+�gUx��UqiU^+�U�]�J�⴪�*�Ux�UW����������i]"���*��t��U�i֩QUUU�UqWJ��]*�t��Uv�ڪڮ�i�ω>��Vj��ڶ�cj���O����Wl⪯X���Ҫ��*��ҫ�V�V�v����]*�*��UUV�v�*������*�q]*�ZҪ�Ux����U�]����U^+�U\ZUUťWa����Vjƭ��1LQS��ǈQ$=�{���yU괪�+J���U^���-*���J�������Wj���Ux�Uq]*�UmZUWUU�u��n�U�UUťUW�UUťUUEUUX��Ջ��C1Y�D����pE*!QU�� 3�
��*�qF�"���E��EL�c��юC��[)[W��_����**������??�_���c_� �S�~y�G�~Sg�8~��6a��:'D�'DDN�pK ��"lDDN��H%��D����4p؛4&� �%��"tN��D�:'DN��%��6&�	�(�8!�!�A%�DD�bX�:lCf��҈aDD����DJ�L:"tL,K6 �AA�4&��B%��c�P빕���%�cu=���_3,��1vH��%�z�ؕ*��֬��䍶+U�+GF���ME+�E ��ubc���(����b*H�*cR�J8�L�TҨ���E��v �cʫI�2�1���b��V��n$�K�N+��L�(:���C��F������JA8�,nL��	�:��jlq1n��R�ձ���Qq�� �h�QV���C�kQ%qYEF�Ƞ�ʥ�
VH)[���qBD���M�蝊�HJݒ�%�5$����4�ٜ�$ۑD.e"U��EIe�D�e��H�Hq�7Y+v"��9�H���jĨ��z��v����;:ފYR�*�+H��Q�q�h��Ԋ*�$B�+UZLR��`�O⸅Y��q9r)��f��f��p��j�Sn�X��"������mb���َR�b�m6"KkK$�9[Jª�^�J�9�1ڪ���7�D��*RWA�[�A��JB�D8݄�q��*ۮ��ESU!�J��^>.m	F��ժH�e���iQ��26H�Q"�)e�d��x�ƪ��ZF!���\o �B�+cc��;�	�Z2#F(��qcFcDPf,�Y�D�,.R����X����\1B�hA�(L�AE�YLv��Aep�&&�Ab+&)c%�Z��YLHYd��k�c�8����u���R4p�f���sD�O CaP�q5�e���,��IX�RBBb�)2��y�!V�CV2�L��ĉE! �����d�1R��YI�*���!hv�*1�d��1�Y$��pw=3FjYH"�5k��T�̈́�2Ҳ�V�T�FVZ�	(��x�Y&2R�2B�	
��Bc�"1�D�Qq��4] �!�X��%
n��&A1
�Z���KHQQ��&'h�����++�n�3.1��؈*��i��fJ6�e���V�"Bc���"2d
YT"R���찺�Q3)�ɂe4��!�b<�� �ɔ�	F��x�8Q�b�h#  �,1V��%XОtF��b%�2:;pcc �!�+�O" �2�����
Ad.!�!�v�"��"�TKm�Y��8�F!sEŸ�W�K+�)d�Q��8�q�-�,Ep�24�Yc��?n�|H�M�IK�D�N*�VU�H���UU4 ��ۖD�"��ZWSv�	e�M��e���Qʜ�Z2�[&&ʕ�m���u��F�&�J��U��1�b�~U*Y�J�+j�'��k*�ڱKc�SjD�KV*�嶴[��[M����W)\�Z��u���nWD����Z(�X(KS��V	��"��:�H�6�8!���h��Ru��bR��e�E�
V�FE<�z�Z���GUˑT������%��b��R�����Ԡ�i���'
�����Ӯ	�7Fڏ�MK.�RQ8؅1���W�0R'H�x�i,�!j�m�h�����R����&��==�7llLtjڒqRW[!$����Y�4T���1��m*D�cTi�m��:�nEmDn������&��J�(�XƢ���ક�9��X�T�XB�$�a�KV����lT�I�Ǵ����-Ę�r�J)85XU,�NBQ$G*MB:*"H
8܂���vT�����k�B7�r��MEm�u�3tIq]m�kC�8�+��Wd�Tz���k��}=�g��Ȫ�wwj���>��{����yEU���W��}��O{����(��wwj�>>��{����uV�������UaG[u�uխםyǞӄ8��7���G���J*G��j���K�	(�4(��pV2dIA�c��!r�I2�A���tPrQȥv:���7+�'��V݄mج��T�TC$�ؖ$����HI��8�$�5�Q�-����cto+�P��K��"\e�L�d���e��A�	-Ȩ�P�4PA�X�1�h�y�e�(�G� ��H�ZH0xR�
�׎Ҕc(�<�T�,DPc �,���Q����c�Zj�X�P�6U$L��mQ5D�Q�%e������%$�Tu��2�#	eY��5%r¦7&U �;�+%j!TM1�:ے$�bīHv1X5Ru�q27i&F�%��G	[�jX���Q"=I$��E:}�.�_��l�����9���n��Qpy�F��+�{��.�F����Q��[�%����fh��l�ƻ�nT���W��<�[3"}$���a��y�U����Tqۄ�b�����ǟVϘKIKU�W�:�(�-�˃Ҏ;�?��Qw���J^D�5��gx<-q��;`ǿ/��4x��Ǐ��Ǐ��ӄ8I��DGRd���\�ܒH�v;3�h�8q'�U괍Ą���f�WU��'�љ�̂8sC)L֗�&���*ˋ�0ߞp�'�?�o�o1��^kP]IQE���[>�b�����뒠kEv�wr2Ⱝ)�i������Z���u�^q�N��6�mS���p��+1����2I%:�0R�XCE2o���0��fWa�^���Z>+@82�����"����c��C�N�WJjU6����ª����yF7y��t�$	��1U��F�� �K�	+\��'2Y�!��FV�a�O23.#�)�}�L�iJx���]yםyǝ:�8�-�;_fc�2�krI#������:#��E�z�Y.hŦ�qE<�#�����2CN@�� H�١��Ҷ���V�j��f��o��*�nu$s�OV�=U��ayռ`��:&	���p�÷͗+7U�q���d�V�q�#+a�[��54]����!�1�RI%�_:�U��I�K�^o:u�ɡ�x�A�t�Ho��EшgNy�/C������v��k�Q�[zx�[cƻ���J7����j:gs���ď���+w�p��P��[lo;Y��޿y��]ه� BD*�уG!|$��m]�V}��֭|�I�9Vn���tABw�8�ֻV�5.!&�D�Ϲ���fo��*I�o6�i�]yםyǝ:�8�;�����-�5��7r�X���JGCƋ!\�UZz</�@�kc��I
���#$����%�h4�����"�Ֆ�u�k�m�I��<B�W�f���Ą�mI:(��Z�ߊ���X�a"��B��qfұ��h��8cW�q��y�^u�^q�N��6�dHd��b20�J�I$��4zo�m�����_����0X#��aB���HTd���7G�~Ƴ���6���o�C\!!K��XG�4�Nt�2}�a���>���\k�Cc\F���-~4ϱmU�L<x����m��[έםyǝ:�8�-�޽WP�d�H�uc���D��y4gTtCjeR�(L��%s�����_�#�=��<�0`��V����"Ad�5�C]+���Aup�:�������a��~���iXTG�e]V�6���u�^u�t��8C��^�o�Pq���Z"�c�L�#4X�C��r��mvſ6s{�C��Ƒ���("	��M9XՓ�$�W#��4��}���y{��r��4�����;�tᆹv��e:pV��Sc�&}�M4��]�w��Y��~{�V�;��{��k�u����}+�~�ѫ�{~�ͱʬH�m|��n�č���č�����n)و�>�\cFM�d�V���>�s��'BA������sC�Mӹ:���lҐ8lh��ŉ�1��3�M#�v;u��!�1�e1a�9GsFK�s4�V�����:�uםyלyӮ���4g3�n5	D��H�4�kӻ�b���pd.I���#�bJ��O��"�Bꌹ0?i���	�Ҟ9$�8�F�Hf����T�6_�i�&��L-f(��\]HW��e����rA���S�8��}�����) ���e3���d)��O�c�Z??0�Z8�ka���cIo0��Z�qKO-�O-�?�<�~m�#�~O̱���ͱiiii��a-�[�ţ䴴�6ŧ�o1iV�[o1�-�'�Z|�����,Ţ�1�יl[�Zm-x�M��Y--x�[6�m�KKy���ao0��lZm-�*�Im0�l|����aķ��D�E����E�E�F�*�e��ҭ6��Y�>%p�֏���0���	<gF�c�ik��ٴu<�6��lZ[,Z�-���N�-<���wmlmFd�"�*>[x�c	WRE�h�rTuJ�Z->E�b�[h�Z>[F�0[�	T����=_�$�����lY_W)�$��uu�Yδ�VE=���S��������w�[�}���Mz3�������%U>�}꠽�6��ۧcu/�����7sW�S�Wo�s���gǻ��;�x�o'���r%(��K��vx�	����F��Y�Η5�F�jd{��wC,��w]�u�w��j˨a��8�Ǜ������\����O�Wz{�o{��i欗��o[�O� c�}��~��Uw��o��og��׽�{��QU����몫���ww~�߽����z�Wy������]���������n�㎺���8�����0�5�Qi22[���UUSA����I�Ȭ"�����"���e�b����������$pٱ�Sm�R��]q����T}���z;�`��u��d��*�/�w�'9���M94�7$��7���� ��7��C�={n7�ۇd;&Y���(�PCV8,�B[
�%��; ӆ��7��d��= � ��:A�i�]&�u��Ƌ��s�u�Ns��I3�i�����~�6p0�K�mc���9UjD�l!�ˢ�0i!YJ� �R�N���ߖ��:ۧ��||#�:S����X���6��m����$�M��	��G֖%A8�(���>4&b3EN��F�����FUTs$�q\07��1@`2�dqH�d��A������iș2�l,M�ӪtA;Y¹P��F��b�V�G�0��bd���bi�D�$ a`�IPE�b�t���2����f#j��#�1G��LI�zɗD�@����� ��v8��1!��"71%*J+-����yoμ��<��||#�:S�$�K��(��H��R��\��H��*J��+���jH��R�m>"b���q,�U�-�d�UU�o����7��7��5y�a�9��5>ӧ�M�}��.jgo{�Hw�z18p������<v7��ͽ[懽�~���T��{��,���^~���n�G�M���s�;�駔���V�#N8yhr:�j8���t�2�T)��y�o��s�mI'*��F��L���Һn��m�0�_�
�a]��Ec#������a�gl8����̛�!�J`�C@� /G�xG���5:��RlqvP���#%�0�Q�CaC��!C��0h@�C��4A��,8{��~��I��7�t��ȿIH�V�? �G#���2��``4�A�ၧ%�B��#�Z��]�᳧ͭ�矝yלyӫy�Yq����ws;����UU��B�2�0tx�de��[ե�� �0>t�v0�
�!̑� O���#�)�f,��,fH�I8�w��(���F#DE��:9h41�+$�gJ00B#�:#���NX�d9=�=42��e(|ق���"Ӷ�a���1�~��d�c�CL�|�E�U�d)�ć��ݱsB@2c�AȆpZ�����ڡ�)�>��V��1l�Y��J��(a �� Y�5���2��r���� ��_䈈µQ�4ד���6i��1���?8Y���K~u�q�N��î2��n�y��k3-�s���UZJ&�$OйG�dXýřd ��4-�P䁄��4����-d�����!CP+b5ECBQ�� 1xt�qzGM̎�kn5�cEåJ4@����Z��1$nf���c4�#uVY\��Ft�%�¡ 2/wH��n�h4Ѹy�FA��m�0��0A2�4�Hg.`2�<6S�&��,���C态�0(Nn�Cd\�>:�3pl�}R$��+�Rj`�(!䉰�����J��SC(�?T=������U��[<��~~���<��_�u�ϜkU�{g�7��*�jV��I�#Õ5�UU-QZFHNGPf�)KVpHX��M�K�p����ڕ�\�C��{T�c��)��Ըمs_h��˧#�¾���[FQ�]J�}����6C�+�:�i�?*�9�*R!j��L���$A�䱳-`��HB���͔ �a���ǪU����E�d,Z �`�b����]^4���D�O9Ta�>d�D�u�&�~hS�$ ��@h���(���+- ����2@�Ai�	q2CCxa�D��������ǎ:|t��x��g���O{�����������?s���"��4k��(��B�'5	�x�*k�q�2��m��99c��n�UTC>���]�r�g"Y���+Rk8q��v�p�Fh̓'��-.戆i��9���Ä��;׭�>-�Nl.=�o9��+wR�����5=�jf��EU}#�(��(�4�E�$C�by�9��]l�)����7Q_C�>���-*9)�b�,S4Ƙ�	�7�0A�$����7pLʄ�����YEiciL���)��&DLeo{���G5�d�{�O4�9���j�����CC9��0��F*�i�NWh���~Vz�ز���Lݹh� �!�6f0aa���H.�O~�ߵA�����ea���X&3V�Ƈx�	WE�U�8�AJ X�OJ1gePS�`rА��J��-�V�����<�Νul:R�/�&6n$�Xʪo��4��UU*k�~�`J|��H�s�DfUG08������8�����$��i��7=�e��,00�pCE�mɃi���LEa|a�>f���&�>�i#�He�cDm�Pќz��3�v���sBY��q!�L4G3�~>Nv�(6��vSN��xa��p�%A!���(��O�kn�L�k��C�;A�WU��W����En�1�&�՗Q[Bm*`�3���F�ے�!	0��pI~~yo-o�μ��<��Vî0ÇC�%{�]{Q��
_5n*������FEH�0�B��T(ʀ�8�D�tA��0� ߹\δoRQ����2B2��d�Du����8�4����b��2ãm	�49&����A����{fʆ��J�c�>���*]ݕ�/�~����OX\# �a���M0r��`����0�Z�3f��0t���LcG��$!`|�h��x@8��A�9����`z1�����R�II����M��`�x�O'�	 ������SWɊ���	O�>m����מyǝ:��ǎ��Q�5js���˻����ڻ�mt��9��򪪈W��<��L��pX�D!_��paFrRl����>
M�(qC8 ��t�~R+,toCMQc��^��^2=���D$"�*�ZV{��LL���S��s�La<9q<M�Cd;�����u��2%��ɚ2B�
pjN\�.�����iacϛO�D�ls��D�A��D��DK�����0ђ)�����rCe�i"�&�$!a��K�Iq-��>?VTω�>4Q��~p�O��a�V�N��ŤKKG�ŧ�Ǔ�1�؉iii��im�iiii���a�?&�i>~c�i�?'�~q�"��ah�ثM�l}%��Zi���KH�--��KKN�������-�0�KK��������~g������Ǆ���d���d�Ƅ���|K%|K%|X�E%�E���I%�J���"�	Ĵ�ZU�hZq-+��V�a���|�=�]c�l�[��-�y�M���fZE�il�2ش�ش��%���o0�mlmL��E�u$��6�ċw-"ZDmFҭ>E�b�[F�h�l-��|_��=�Y��.~��3X�G/.r��^�Ӑi$���I��\Q�p���	w��Gy����yGk,�{Wc]��=��hɶ��+�%~������~q$�Ěe�4.�'�!9��wv�q���w�Wz������s������
���3�O��#io���s�i��ɽ>�����Y��N�<��J�9ʶ��L��Jh�S��V�J�.G�������=H�t��TsX���������!��2k���K�s-���w��f�6ZK٫���b����y8GՓ�O���k+�LV�7�V�%��$�D4�A��R�Ek+s*����&n,YF7U��Gj�Y�"J�pU6V��H<r~�xl#^�w��Y�~�C��(������������Y�������{��,���s{���{˥U��}�]���y=�o����,U�.���y��㎺����8�]G��:|����T!*��v�H<E�4�(�D�Tq�M���Х��R��,�["�rT@YJ�C�PDw6&&�-L@�X�KrbqZZ��lC�RBP�B�D�Щ�!+�EYI1�J���ǋ%��J�3I%#%#,"�ǔ�*�*
1(,�F<A1��C˓**�s �!�c�����ZV͔A����Ҽ���H���W&X�*���I�UV:�4��k���;��kU7q"�RX+]��N�&(��e��QYLm���$�N6��8"$��T#u[h���r�ʩ"d��N��T��_s�ytg�nd��s��j�ɽ�o�^n
>���-E!���%_���ǁbC�k�ݍ�w�x�<���j��k����������'�w��Y�D�8X�n^a3����Ɔ�ES"M:"� ��?vU|�M7n`lr9�Ş�85���p��z;��:1�6RC�!*��>�TІ�7��Z�l��V��!�����tl`}��2����F�d2d��F�4̾l2@�FA���s|b�gC�jP�H�B���բ�+F�K&�!�K<%]����}���%qK�3��I�_-��{�+QPn�Ɉf+,|���scz~,���(��p��ǎ��[�8�]G���by>������J��Rt�I5��Ҫ��W�0る�B��ƀ�4��n(:1����<m�!0m[�w����U=XV�u�Օ��0hh{�8�&C�<v7�����l��e!8 ����	c��bч�*3�
Bܟ5�Jh��i�?��ir�BJ�t9���>��I�e�4�|xň���L�bE�cCD ���h���cm�f����u�qOe�_Q�+
~ّ��U���8��ׇ�y$�����S�:��??-康�q�Ӥ8|pÃ��Vd����.�U��Y�$�UT�}_���*@�h���?�>r���C#2ؐq���6�\;T�ի�*{���G����7���� ��aٖ�jRn�2�*U�	�'��_1!!P�fg2������T�Ȓ z!_NU=�SM�
,�m�>b��ŋ︒5�����2���Z�ꑶ|��S���L�>����0�{��Jj����!ᡶ�9�P�DʘAe�)�#2!�X�W[|�έ�տ<��q�N��-����h���̹�/�yUUH�⌅S��n���L,��
1��t�˷�%a#�~���IZ���}���m��9�l�w�x~l|a��Ɗ�MB�0Mm���[��UG.�PӇE��,�m��Zz�)�P�G��C
d�Ä��uHH�����]W�땸����=���QD
�ECo�9>x�����5o�V^W�QS��D�W� �%!卐0�2��:t��LS �q����1�44��mZc�a�ז������q�N��O�Jt��e�Ϳ(rf�S�8R\Ջ�p��җ��ӗmb���j51Yx�=�;jn�Fթ(��&�|�c�yUUH޻���K���;�7w��_'a��II�:Cy¶f	P�ݏl�|ћ�t�J��p�{�����#;ל;y��c�I��o�{�x%�D!�h��	���7�;j��k-�-�)�ph$8d�9lu<��-�X㕲mP�0���i�
������J��Fb�����%Ƈ#���.����RB�R3��� ���i�<f��`�$R���I�#���E�k'Z<D�n�п5�T���ӈn���8�Yit��6�]��,�k��앣�+̼�����Ya�y������O�u�ku�����t�<a��Fʗ���v'$�z�y~UURU����Q�d�I�}MZ<��3�c;��2B��� �s�P:x�Ft)�Fi�%JQ���0a�����FfXJ4�4{Ci�dr⌁�W����#!����|M>�~�C[՛���H����jߞ4d�-�CL����)����eɜ�ɚ��C�bm��g8��yki�k~[������N��ώU�t��b�0��UT�|g	˲��X٣�ϑ��Q��)p�[%2_͖����!���������CǡDf��h~��'jiD�Г 1�C����]y3�|bd;�&~�b�8N�������L8Bxh�N8g��0�t����}W��xx $���E���}u	L�Gܢg��xǚo�T�;��O��?8�ߞZ���:�8�+j�"~��x-��P���,���m��b�0�F@��HgfL� n�L�q�)C��?	��������u�Hp�,���3�B��:|����k61:t���ɮ������d{�Iֵ�VnT��愯���X��ƨ߉�m�	����E�����h�h�IUn��:w�2k�(�x k��h~o��M���-ŭ��n-Ӯ�����>F��})��Ga�8!,X��1$�J��H�y �A�ܑ%��UUR^���d���h�Y����wI�4L���,��?�Bs�3ᗇ��y#���;�]!�=�ݥ�_��-�2�1�\)S3Z��w�:��߽��~ާ�����of7!FQω����B͆���e�x��܏�h-�C�I������çc1&5�$�\�ul��Κ��Oz���2�!��\G.�-T��T�W��]}Yl��5���2M󎝢���ѿ2ޞ::4�a��єN�_�	���~_����u/�<#��$r(7�g�E�1���g88c�=�X�4l�����gO:��źu�q�V�o~�ڴ����һ�K�M�ָ���W{�?}P�S���4�Ѡ�Y����y_��?�>��x;7b� �"#P�ڄ$�68r����svl!ц�%Yd>C��ʹh!F)�C\͔��	�^�$:~��lY"�$������*٭F+|ի��~��|�6�w���mʏ��b����L�6GQi�~[�0��Z|�O-�"��a�i���e��|�"m-lelZ[l----<���KKF�o���ӌZ-�K�ylzI���<��yq�����/�v�^T����el�Z--��U�䶘�Yx�ŦR���^e��I�G�ŧ���l~6'�Ą���hL���|["є[,a"[�0�*&RI-"-$Za-:����S�u6��OĮ���&���<0�'�q-y�ť�ť��m3��lE�kę[�M��K{�'���b��a���i2�R^%J�Z".J�"��a�H�#�Z->J��W�ah�ZW֘Z-8�k����߽����i�*���T$3(��]o��3�v�9�W/~���עꍧῧ�⏈�O��^.<޾}W�7�s�[��m�z웾��ϸŻ���s�J��>�D}>��X������G�ό�w\�tȊ�n���}w2+㳚9��F:�^���[7,_sy�p���_(Xek�[�����	? _��_�����������{�ⴭ��w�{��Uⴭ��w�{���U�i[���]���:㎺�n:����ź:C��:V��UU n�ʵ�T��QŒ���1�������F��׺ƛ���J��J��U�ϙoX~:h�	I���֊H=������#��_�Y\�ƴh�DTcƑX[��0�ur�C�]0�}�ɔk���Α�����ˏ�r�O7(�!���TJ��gFq�9��T}��Q��Zq��ێ���n-Ӯ����fLcޱ�j��5Y,����^�*��u��ej���*&U�q�O���W�M��A���F�O�?��4(����i�f�Wr��z[/i�j�~�h�]��&�9s�62;��x��N��@�	o�e8l���BFiBdH��i�ޫ�D3F�,�����P�[�\+��BA��P�*����難�2ӎ�-��Z�Z���:�8�,q|�ĕϘ�k��f�A�"�Q`Qg�t�Σ�^{�����^�kmMʏo���:�k�Z�-��7��ʪ�@�g���|��No������.�wޗ�쓅G�G�;�6N�cΛ:iu�e�uۢ�sy�������N.y�~|�����{ۥWδY%]ǲ6�A���Bdw��]ܘ�W��~��+G�t�=�6�#���R$�]}\}[��q\�����b;�I��^䛫|�M&ُ��+w��9)��Y2�6x�:={���~�!R�d߃��c�'p`��n��߱b@�Ԕ=��!I]21��!��n�l��uo??8���ZַV����M��V"��JƧUUT�����r�|Fp����)��zW��LF:���6��8�����}ZoJ�Ch��i��rO~2Hd~9n�ID2n�828z�0td0tS�}���	���N�wtQM�d�`hk�[��R˨	�U��a�w.f�VӤ�~��Ee[J�(�th���|��̝(��gO�ukukZ�[ǞG[em�e��v��Z��%��k<�����"EĜ��h�W�n[��uSL4�e��d��~8�F�k�I42z�cɧ�@(ΙiC�C�$rB4�0�U]Y'��:p�&�{E;�t6bP�p���M&�J�O��)�L���'�$C9w�7+�״�1�h�������g)��i�>�0a�CA�!/�'=	��0yW0�,����y��խkuoy�,�{-��Zf��UU Jk�:S���ع����Jc3�C�o�Kk�����a��o{+��)&���ݖXA�E=׆Nc�� S�ِ��g����;�L�8��T��G��B�e��p[�	�ѨJ`ْ��͆C
o5_zJɍ"�n�������է^i�~uŭ��kuoym�k�sx��k_q���i�:��)(�"74UK4X�כTo{ÑԌ�t�p�,n%�vM\��|���{��2�߾̛��|��M�/D�(�~�Z�rn����'�<R|2��ۤ<u�.t�>�8x�v��3�U8L7��^��^U��3[�+�\��>uN��l8RQ8�/|,�M3��W$������1����H(�Pm��#���n��4P|������g���Μqo~m�Yh�s;�.lqY$�,�l`�8�#m��Y��Ř<rN���ɡ�C��/�
�n�{5d'�u���t�Ĉ�:kt2J���]rBB���<}�$%MF�0�<,@����K��YD�O�~����:��[�[�x���l��و�d��H,�zܹ��UUH��U�8Q����>��:�M�93�_2h0>�e2�R�� �c�̼7�&0p�l����Λ�N��p��q$#�7?��7>�/�vȭd��&�%N�H"$��
��g�u~Eb60��~&	�6;-Py�l-�������wl���_����GO��8��������<�:�,���L���c/%�UUH��b��_O��yɂ�^o��?�z���Ӧ�h�TN6?,�<�m��[��xL��>=?t�1\�q���P����!&v.�ss�� �0�������a������醆h�N@��dr��Z0CsLa$���n��a�&>DB*��[ο�^u�8�����Z�t��L�}ǎI�/�!�)$aէ�͸�ĎbIV�`h7��UU��_'J�|9q����m���ad!�ϮəU�0��!�������ñ�`�0hR�.Gْh��Hq�W7٥}Z����G�S�iZ{䟰�Q�b9��5�UJQ�$�9���S�{(���=��6Bw�<7t��!�=���
e��3̝��Y�Z�F�p��
<G����0����-8�[E����b�b�c��|�[lZf������M��KE�Ţ�䴴�ZZy-�2�G�Ǒ��ZnKb�[%���ؒ���k̶2�---x�[+O%��9^%[��[^&���o1h��obF��Kch�lm-�I��Τ��KgWY~f��L"��ˤ�U^T�T���S�e�-u�&��:���ah�Q�'�\�J+�C�t�/�+Ş'��Z�:��b%����b�b��n/3�-<��Io0�nKa�i2�E�d��"�"ȴ�i�iXa�Ɇ'�\�`�l-KE����/�����{�ԟ�yϸ.�)�v����_9v�$���jF���Uf�K;�ids��Ǻ�����������齝�u/z�v�k���ܐ�fǸq2�G)nu������'�+�`��>9�>��pӌ�3d�_�.�8C�g�Ӈ�i!����"��_V3��^����J�"��}I�z����4�Q�4E$6P���z�-d�a��h�ޜ7\��}��u;��I�w���ܟ����sښ��9�t�j�#=����y�!yy�������U�[GSu'j�ȩ!��48���޲!I�)�	��D?]+.����.��zۮ�m��#��*�jm퉥D��YebN9i&�����S�Z����:ڴ��9w~���.�[V���������j���n�˿{����U�]-߹w�{�æt�æ<[�qkuӮ��2��5�>���$���ēQ�XX��aVR+rW���Zpv[T�F�����E�H4�-D��&���!dJ�q:JW�R!+���TѤ�P��Tx��%r"WP�)i(�Q��!K�ѐD�Ie$��*CA)J�Q��E(�q�x��pE���񍪲Q�I��Rܷ���"�R�Q`�rq��b��hWˌDEb��$nڬV�QMH�
�5cq�A��Q���F�qX'S��$I�A�Uu���vV���I��)UU�+�Y��ĭ����$��֢-#n,�XX��Opr�(���Ěw�����C����{���ɦ9�X��Y=/�W�o�sF�9����!�_H]���>C8_p��s���O���8���J��.��!>ޯ'd�y~Gٯ��8rW���owÍ�e��_��s�1G�V��p|g~��n�+Cֆ��Q�%�s�����V�����X�>��xzM�1��ɂvsc������"Vkj��S~�`�� �����pш����~qJVn���8}X���'�L�D�!󫩊�G����v~��k�ա�Y[��u�^~ykun�u�q�^ӸZg��.�\�W���~UUi!ev��}�	�G��i��aXi��H�VZ?O.��N0rp�)��l��`�v�y���BW�0g�(�id�drs����5%p�e��T]vWO�#�%%�El8ws�����%�D!\t�f�n{)�M�4�^J��jI�ڮ�YZ��}���L'�ێ���yż���Vx�x���Ao��Bbi�As�m�ꩢ�$ё��3�$:B�Cs�!�4	bգ1�2�gٹJx'}�'�8tG�W�zT���dPRBt��e8*�T��c�E��njM8!Z(}���!��n�$��h�}"p�	I~3Ʈ�nJ��ܒl�G�o��"�9����v� F���b�*V��N���y�^[�[�uӮ��2��s�1r��2B����C)6Y_W(3��8�C�:��۱�0C���ަ,.��8zCѧ�Z�d���`��ӡ�ԯ �%BZd)�P�<�������8gD1�|����K��6y�gç�fp�
rr�!�5�xQ��衲����G'��p�#�ͼ��o-n��N��4����Y&n�xN^9nϖ�M9���v�I��Σ�N���N׼�X�rG�y2̐��}�I�w��_�{���o/kf�w��w|#�C�Mt�{����S��,���N��eF��yԾO����ݳ�{V�F���f<^�9l��q�nzI���ړ��H¸l�鶕���r����Wƪ��Hpi+�Ń]�h�H�����v��V|~�P�n!>
9f��ދ
!���J�}�\�i�f�W��������p���?eQ~v��qT�S�L�p��צ�̐BJ0B��w���\�*	;ui���q�2p���Ν6y�疵��]Ge��=��&sLf]�UU��������V~!�%}U��ʭ^�x����e�w.�L�@�����M �Y�a�E����4h��p�����e�!h��h���aL�X���l����˹,!2[(��c?��||g�� �C9�|Lg��0�1���S����k�U�W�ߙ[θ��?<���ǃǄt��/���d#h�z/{�UV���d�̹�HI7K��'�$��)��C�l�%�X46k΍�D-�f�?�2C��$!�2�-�9���p���c������t�ͅ�&�[���>i>z��(�>(lm�e�G�zz}�\:U�~K% �R��"w��?�ܫ�!$K䲶B@!ս�Q�N�I�c��������~[�Z�uӮ��������.�6���C���(a��f�\��8�&��g,%L`�����
T8H��[!x�Y�����p�J���X6��z�t�d#���|ѓGQ����:l���6C��I!��)�Z���I]�O"�[�7j���_#*�eȑKk�����D1�t��dvx���V�ۯ<����uӮ���׾�X���h�{��p�62��mx�np���m�51qSuq4�iŎq��n�Z^�3���|���A�r'l��5&{�gb��ۏ:�q��7�5��O4�E��"<r�5/�oW=���𧗡�v���o��.ﮫ����N�u����N=��M�a�;���|@�={��t��s{�������x~�md��x(��ip�f{�2��A���^�	���0�	!���0g�Z��>B�>lt�9(�*��J��l���t�g�,K��q>wv����'ܭ����/=�|�#���+L��fd�+�h�x�����4|�ߞZ�m�]GXq�X�kI+8�PU�1�K���
���Q@ճY�UV��~���$#X�A����I�s	Q���g�P�9O��V��h�`�<�WO!�7!a�8L ��š����=q�����Ҵ�_t��ƓS�H{׌I��DH��u�S���]�n�k_T�k�F�i9��̐�8�Vg�?<��~[�:�:�J:"tN�pЂ"&�J�"Y�H"hD؈� �'K6&�؛4&� ���DD�"p�,��'DDL,K�؛4Ɇ�bQe��|��BtL8hL��Ye��mխ�ֵ����ǞG���'K:Y�ĳe � �	E2P�blD�:pO��g�ʯ�ν�Na9f���J˫ޞj�{�ٚ�[e<��mf�Ԯ��y��o$�����_�w���o�n�g��$Ν�%_:�'{���D}�q�e��y�����_:����|&���o�_3i��w��zn����-g��h�Z�}��;r�3UA	�Mֵ�޸�+Zl��5�{����t�w�{�=�y�]��n��~���{ͪ�WKw~����{�mWj�ۻ�/�����m�[�[�[ͺ��6��]�s�UUi!�����!	$�}�I�C$�S��!����[�*t�Ǜ����:#��1��;]�����\�h�wi_��8zQO��>tK���q�0C hyj4�3\Du�'����^~w�P�F�0s�ǜ$��,����n�l�Uu��[��oͿ<�����u�Q�m�>�NƥI$���S�C2��UV�rJ��x?z� ��E�!�0�aN�0Q�|0�|D�����.ԕ��t���J��8�HZ��}L��}U[mX]~�8�ɟ�9�fg=U��^	��^�TVK�2�3D�����*L�a�aɉ�V^W+.+^9�lI���{ª�8�|}�ْ|35���]u�ο6�ߟ�Z�m�]GXq�>�~���L������7G��������U\;,LӰ9%��m^eKM�n_<���C��4G=Y��������}/[��9��e9�빭t�t�:/���������p�xD:w��~��(��1��t�-V&�Sz/����I�}�=��]��}}�>�q7>}<�XH������Zv�aG���������+�#��o#�I:a��b�M�Y�~�'܎ߌ�p���"#�����w���^v�����TW�h�v��~7E�ć�!0��&�E5Tm��6B���i��nvQ��c<x?�m7s[��X�R�$��ӥ�2h��&��
����%�q�Ɵ�u���<����N��:Æ�;�n[`��U	�uUU��-�dΚ�A��ԗ^�pcB6H>ٜ�o%��vm�}��]�2f��Q�FǏ�Ɨ4=0t�%�8����t9y�7��T�~�q��[Q%K����8d>��f������������!�$��YQ��XD8�D}�h][+y�ߛqտ<��Ӯ����l�>Ĥ�!��}2S�rꤦIF�cW�UV�������
��~<����!��f���28!��!��8C�ڦA��,�t���!�|6�B{9Z�	W���}����x�3|%�S��92��W�	�`�,>m��$Ӭ��3&:���q�L�����Đ���X�d�nӄd�ǝmמ[�[�:��6�W䞒�I�$�;�*����^�2�V�H�bW0o4�g���?6}��A����#�}�.��d��JJ�C�S�=8C�ǝs�T�����!��U�[l#uT�2z9"M`��������YTH�W>i�&qrU�!���h�w�|�����i�V|��yܟqki孷^Z�Z�i�^�8B��F��ޥ�G֕��e]v�pz�	Y���K���V�&6Y+$��%��5�UV�{���=����p�w��XtNu���QқN�sf��\�Q6'�;�p6oz3��5q'4~zJ{�U)�;���#�{k~�wt�`2���3����+T!ʋm�o���]qXm��$ړq�i�⸈��>�ի�i���G!K�S"n�Bl�zl�~���<pY��АѢZ0ؐ���i"]������$��~p�;��r�D�V�o�͸���Z�u�]GXq�W�{�5���ə�i5�z��I�*����R���aXa��kuw1-�ܢ�� p���ǌ���%=�2|1�D80�Z��e��YH��7UP���f�O]�t�5O����'Џя�Ի�%gT�p�Y����#���r�4KUoV��~:�0ELoֻa�=^|���#m_G�p��Ǝ<x����ƞ<#�:p�M	�{-]�J�Ҵ��*���]~�w"^���!����QQˉSc�y�Mp�5R���P[̲}����DeK��I�C���/���r�RB�9�`�d���o���u%�\�S�m����00<i�֕�b1WY��o��5���<�[y��疷�i�Q�m�ޭF,įssf�����QP��Ij�oG�mUZH|V+��6S��k��V����F�BI9�������/C��,�d��{Glt7���#�n���֙���OBQ+�8aC'͜<ݤ!���pܔU�\��7�c�_u�Hx�~9E�l�&2���#�٭���u��n<����:""t�0Æ�HlD؈��&� ��b"`���e��&���f��4""`��� ��,��'DD��%��6&�	���4l�2|��A>AD�:lp�yǟ8���[�x�[+y疷��-h����<��:�o<��K� � �"%"lЖX�8&:Y��\��Uϻm�y���']H�;6��V���\�N�wW'aG�]�b^pK�7�S��߭�x?�RI����Ϥ�?��^^ƹӳ���s\�]jsf%�����K��৹D��Ru�1z��u:�ӛ7�6���͐��߈u�er�hw�����y:.>��({�X��˫�}嗀<x�>�A{����d�8�`��D+i������K81�ɣw ���x;��TOP�z��%�p����m�F��ug%�.т�_w�[:����Cn�����rF�%+���5�qK��:����vѕ�A��K�t؉7�֣I	�ҡT��+bM��v�VH��N��X�,��$�����wx�㽷�|��9�}>���ww����{���t��������y�Uv�����{����]*�n��~�����m��kZ����:�:Í���O�2)$n�,�YmR5G\v!HU\��*���ƋP�lj�ز�
��ۑ�D��:��TD6�+$ySBı�G$n���T��."8WBRZ�I�q�	�"V �4
�-�&$�˕ҍ�,�����aI�<C� ���F��F�%GFK1��$"�n�,��lJȬP�Z,�pq"`�*,����2Bl���rC%!^H𢑺�q��h�$�IG%m
4J:+��6V�#v��X�!�T�8E�D㤖���!#ʫH�)Ub%+V��:��¼�M��IE-cM�D�J� ��XYL�e���qn�"a���dɾ*����0Y����p�w��ϯ��p�&��O'{�V�}�<Tu��:-4�=3F�wa}M���&��tz4;��Yq��_3i�s}�b;�ӕog7�񻷷�m��d��!��JI虚~|��	93�1�M�9�Гf����240c���9u��6���U�8��/������v�-]?!���!n�hHG�f�����G������8C74B>eJ�.�]%������L���4�ܲ�wZF�uƞmտ:�����]GX8l�@[�_A�J�M���[��9�����$����J��'�\!32o<��U(�⦙���.��O?"e�w���}\لC�<FV���W��%�)�X|h~-����#�Ӻ8B�m9U���H�5�����]J]�^0d�φݓ��� ��3�H#��7�N�oH{��5�����?:����[�>u�:'�u�tIطg9�UV���$�Jѡ�C�ǃkÃft0��4QD"l��m��4q�x��i0����K��S}v�"
����ǁ�!���i�.C�$������Y�t<h�}�փ	���6]P�}�����zusM8���������5���A@`i�>:t��Z�yky�]ua��}�i��q��>�f���(fkw����$>��'�h!�A�i� ׶�����-��M1ܳp>�j�;~�i�ǂ�P�.���4v���ᇹ�����T[O=��H�r�S3M��u�Oh�ó�DVjڬ?+&�%[�rL[e��6�W�ƏӖ��R���V��<���[�2�xgN���%���#���s��jh�5˔�N!Q�/3���rNA�an��wĚT�����ڪ�&�g��������g9��w�f�v���y�?�����G/9ϡD_{�;/����W9�9�Ji+�[��j�Uk��VM�XS�w�<��3SWx�����߈�o}��I=:p����S��&喊���z�lĘ����e�T��̑�Y�y
�|^B�x��E$�G�h�,,�c�
=��Y���`h�Q�|i�Id������J��R�ǣ �t���c6��,��c��z�������4朁'<�Tʯ�,�ӧ�GN�<x������<#�:p�cph�Ue#,h��^�UZ+����W�ϻ���$'k��2m�Z�¢/f��dn��Æ��N�
6����r^�@�t�H�HMFp(�w�ʕ���<<r�3�L�#�u��������M��������nX��2?������0��@���Y%3�zV�~y�V�<��[�2�xgN�j����)j#J�$�d(��UV���YeܑD��K�L�HI�p0��]v�}9A��&���OA��^�:{���ɫ��G$'
�ŶJ���I.,Im���/�x*Vf���h|�8�$ǌ�`q.�4s�t�����!!��i^1&2|���M>W��lҼ�����:�^~[�2��6X��	1���q������ОB���2��t6} `��9*��So��O�L���L�gC�##�:FX��d��}��V�t,�3�f�;yn�5\k�p�����	E��@z�t�㠎	�C�E��ѱ�a�9*}*����?ڏ<���N��������y�<xG�t�����"|��M�K����鷧H83���&F���o��y�>�LQ�����":�*䒻�5��ߕUZ��&殽os�kM���7�;h�ɾ�菡�s�|<���{�<A:p�O|h�OtGQ��r�_s��w��X�tk�Ϝ���𘻽�_�(��uR�e_ �y�2�?�9ե���\0le��`��&��l��+�s$J6j�}^��?�H��h��\�[:?Q�C�|F�a\�H��K�Ε�U��ç{*A)g���B��BƘE��	\�%}ೡ
�v�JҘ~��m?>[o8����[�2�xgN��i�XA	8HfW�2�7�UV�6�?l?W�����g��iD�y��M�m�a>ɝ(�:qbY����C%3���9�QIA��`�eÜtT>uj��[��DH�Vȷɜ�3�C�N�sM��&n�k�́�ßPhzS��d���+C��/�!F��J}C�/�<���S�������D��tN���0L,��M���0ЂhDК,LDN��6`�%�6hMAB"&�hA��(���0�ı,M��BhJ:&4h�YD�DJ��<�<ˍ<�m2�Σ�[��u�x���ֶ������D���� � �"%&�BY�0LF�7����{�fE���o���z�9~��M�d���=��=4������/���N��x{�m�i��ߟ1u�]�Oӻ��xo۾��5���q��W��O{/=�w�qS�:�ל�_6����sa;��'���).���]l�V�k����t�s3:Ҫ����=�{�����V�������{��J�www�{����yťU���}�Qf8ێ-ŭז��e�Q�9&�o�$�{⪫F�D��r�C?N͒VF��]^+E��8��q�ʺY�`v�Y_U]J����������B	�nFi��������������V���4�!�<d���&J:	��D�#§��W�&�!�S�-խ�n8��?-�u�u�N]^1�<�A4��Ŀ#V�A�yf�n�-��Y��UU���C������'^m�h�j��'�I�d�k:~$�VA%�ժ�8�z&���e�����tl,�[�$���z^����՝VݭD�T�f���9$�JB:���\��S4ہ�R�n�X?Bh�n��͎��e�|���an���-ז��!��<3�v�n;�u�?�H�[�C] �ǉ����֚#8谙1�����q�F��ܒ~��U�����Ɩ�ПFxii:'C�����_;�n��g3ꕧ�Փ�Ո������I��������f�W��� p��^u>	U+�C�m����0$vh�p氶s!���|���G�]�H��$���Ɲ�Ez9�|�Ӌ6BVG @�Dya;x��hݶ�H�2
�����4�X�aC�E��r���<i����:����:�-�������U�y*�Sp���������������F��)0�Q��s!�yg*��|���z8�����>)�h40t|:�`�����Eŵ�����6��ª�<p�Z�	ʨ��͒\%r?+c�n�����@��ӳf<uԐ�����+j�G��u�x�Wն�i�q�_�yky�]uc��W�}5���a���Gj��,�"�0�~!$�=_鸒F����2��>5և�
��G%w�6	ﺖ��7ĸ4&��~�	�2L	��A#���>�y���@�z�����;��^��JWEt�l�Y����M3�|���Z�qoμ���.���e���"I9.�M�UU�+��:~�/Ѥ��?��Y�����G�4�j�D�Y.]�4&�8���e����C�����B�6�NE���N��v�$l����W�~:T����|t�U�u���f��]4�׫��;گ+m-XZ�_<��n|�uo�q�\q�y�������5u=bӸ�m+���Kfe��!YLF�����(3k����>'��*wͶ�o��=���C���G؜���Y��ѫ|H.���g�B�8S��!�.���g�1;fs�+9G��ɜ/;���d|�7Wn��w�>�u_�8�)nC��8�*��!�*���>i<ꮾ�����9%s2	m�hLa�s����Fm��RE�{�&�8t�����F��%!z	P��o۷:Cݮ��®�fx���d!$V�����#���*�*^㪘t���q$|V�̶�m���\~[�<����M�e珥��1�j�ܶ󊪭�[l+֙��R@*S+���a��B�gړ�f��:�Dr����i\-�����]��<Z��u�]��<��@z'�36�7�>y��Y�I�b�7����2Y�����c����$�J��X��#�t���m�Vv�]?[N�:��μ�quc��\�"4�|Ʀmb��֖Q�vđ��UU��V���&�.	�2e�^\�G?)�hG��C�!�C���a�5��d<�|l0p�N�ê��OIr�ݲGJ�;ZK����*��9Lb��p�}I4��yM��$0����!��{�I�w�")�^dI�Ua�V?<j�7Ï;�8�+�O8�qŭמun#���p�,s���YmJ��*��M��0�h��m�iq����W����FH�A#�p��z~f�O�������C�b�4Pô�'�+iE������a��ɔ� �l2v�N5�a�,ϦN�I���M��*9G���i��u���`�:`�YB"P��0D�0�H"h���6&��'؛bl�_2|��6""'D ���lN��0�blM�6P����}�!�CP� ��'��0O�q��-�y�uk[Ky�y�� ��0O	�ǏY�Ś(�xAA(M6&�L8"z�+9:,=7WWu9N��rϧ���wȼ�q'�.,{��×b��ӊ<Y���U��~S}��ߝ�͕���K�7�N��u���Ur�:��Mz�ߴ��߈Wt�牦Q�T�n�A������\ӻ�-ë�;���o� ��t�M
{��ivg34n��ݛ5�!�1�nwf2��Q���^�z���(ܴJ�g�ҕ���"pc �v)�o�=6�p����&�%y���r���)��m}�w\�Y���2�I��e��/~�;��9*��'��\���o���WԢk҈p��UW#OD�1�E�7)��"c�[�D�mM�dku������9�j'8���V���I��GX&]�d&^1�cy�:�uz2��.SM�=�o5?�~��{���*��������{����Un���{����{�X��wwo��{����U[�ֵ�]���m������:��QӤ8C�%?7��8�Q�d���%�NF2X��qƘJ���mUJ�,E��Z1i%U%����4�Wdm2,��8:$,U�)JK2��V�����u\NX�]�n�*�Z�i%��	2�P�XR��
(Q;F
HǊ����T1ҏǈPI(�^&D2�1Ac�hW�yT�<��A��"y1lqb���!0��*��E)+PtEeA)�U��W �ʅDX�DY\ǐyb�iK-O-r�d@�c���$TU�c��$8�n��`�I�5A�U�v7U�TB���h�)�J���i¸K�q6'�bJ�Q��If�Y.G	���Ӫ��H�72F�M¨�n���1awr���UZ8W62��%��?'�����]�����h��3�q;�N��9�V�Xvq�b�����#�qrw�Z�$TRG��Y�Ǵ�'zo"ޕk���q�mc��=[?F��$#$�����	ʓ�V��f����hf���;SNQ�����^pt��~&��!���*�z8bw\�ǹ�%��ـɠӁ���]r{����a����D����>����>����.�\W>S՟����$�P��!��"pN�"x������8(r�;��j�4��ۼm��f��f�n|aC#����z�vd5�{���eʪ���N�C��ex`-|�3���J�d7a)�P{�MZ�U]VϮH@�m�$Y�	���3e�>��v: cC`�uZ��[�S���t�.�J���[�<��-�^yո�����n���p�1���)D��_$�X6q���R���R]�c怇�N$�N~l>�4����0vt�f�G�|i���n�Ǣ"dx�x�i�<�dB��*5^+j��9�6�ٗ��c���cfR���<V�T6�}������2I-��?p�Bgǀ�C��3�6+
ϻxy�mռ��:�έ�u�:C�'"V	Z6�r�V=�IH�4���#�̍	6>�d;~���V�lq+ �����7v��m�ɲ�仟f����C�C���,�L�RXt��vH�6�ve��2Y��nB�Қ��C�C�O���z�hHy��g�2ωܡ̙ZPӒ����S�үI:�2�-���u�[��댶��o������/7b�Ej��8����I�c�#{��ڻ�kR���8Y����I$��^w�7w)���={�m��6VQ\��Ӽ>�L�����������B}F���9�(3��5;������ȷ���]�>�g����|�&����FR#�ټ�7u�kT���{?�F9�0G/�c��a��N��oJ}���c�FNy�ۡ�Q%��S��m�k0��?�̌��1�O��(�	�?�&�r��)0DJH�X��q}S֙��G\~yǖ��:���Dx��!��}��*v��K��I$��v����������Os[��Q$��V����5��͉X�F���+�t�!H�h�*`n{�!�꺎L��sv�s��eN����
�d��K�b�r�f�����?l��<��~[�yמun#���2��g�q���"�T	��$���J���)+F�Ҳ��38Ε�F�r�C��qM+��fJ��`��;
̚�������'�*Q�f{��e�ղ�K�^�1]WZ/u�,�W�7\��_���<ҝ2�b`�:A��(0��
��H�ۻ���F���p�8x��uż��:��Q�m��w����5M���Q��K�����'iu����"#�+��*��T�惿�]cNHq��s p4��TĬ��tiӳ��06>0��Ð�z��R��}�����T:Q�*�ǁ]�S��a��y� B��*op>�Yd���pNd�Q�a�)e�j��T��U�b��k|��y�'DN�0�N�醎�7��q��y�=~V���B@�!����;ÒA����=��Ǣw�b��56Ě��X�ϒI,6u������r-�Ӥ��$��o??p���.r.#�'K����g��|�qw���4챾�/>�a�^�i０�*'��뜙V����bE�L�X�W
�x.��e�p5;;��g�u烮GM�d����<@Ff��,E�6��^��Xo�U�ôE{o��u���&�%g\\�'>c�Ã�N�Ή$�s$�'�����1��Jp`ݔ��Ky�^Zߝqo:�ζ����!Ý������H���$�XS<L
g�hs&~?����=�5c�_�)Y\��1����&o|��~6W�(x?:��H$-�i�C��D�?��$�1F9��e3�7!�=���i�Ž֗S̭�VUs\Sg�����t:|=>��6Z���m��>yպ�:�:��	��"%�AH"hDD�N���X�blM�(HA��""tN �D؈�:&�abX�&�١4%NQ� ��YDu%�bpM�lК<a㮢ֵ����6�Ǟy���"`���x���x�E���"ABh�"lM�`��We�n��Ui��\��i�o��9�9�'a�ҷ�.���璮����tX�Ƚ0]���Q�6���O�k���wy�p�ӽU���~��\w�������}L����u:.���1df��{��ڎ'�;g{8�p^���S�<���_�s˫���J'��D��=�dwȚ�9��{'��5��ؼ;_;��4]v�%���]��y�T5�+g$5\̼���Z�H�n�ޝ�x�f���/����Un�������{��X��wwk�{����yEU���_{����{�*�����_[u�uո��y�[Y�Q�����I%��k�Ҕp���	y�}��W�T�>�����]q[�$Uꅘw��^*�?�eķ��AHё������Un��IgF�.��re�����2��4w��<���1�s͸6a�W&c�$�*���6���U���2�Ͷ��\[μ����?/R�.߹�_�G�\���s�I"|�ن&R0,}��*}%p?a��H� �L�G���D��.���#���3z�4v�k�t�ۅ�b��ç��J<Xl1z�zP���A�Q��kx�f��锄�$�p����2?&����,#�jWU��
�a^��Z���iź��:�ζ����2ۿ>����/�̍j!����E	
�u�Ж�rf�Y����TnWB6�QKl��$�|x<_�s\�c�}�w}j�8<�a�=�u ���ph�d�|#K�k;x\�����ſ|�~�>�}�6̹w�����>
O��dZ�z��>�<�ߦk͑�V��]mX��}Z]l�q��s��ã�����p=h;��MW���'O�'r��8��jb���ղ\DN����Һ��?���R^]I19�?>��f2��eʌ�d�������^[�8�μ��댶��^����eUnP5�J+�I"Pѡ�]1�n��=u��p�BFAI���(�ܺ����oG=�������H@������3�>��J$�,�2���?ԶׄPY+�e�Y�ϲ=^��;�~c�����a�}�
��1}���V�y�]m�^q��^y�ߎ��9�Ϥ�|CMD�C�I,�ߓTJm��/��f�E$p��#�ɂ�����mٻ�]��"V�G|�o ��H�!Ŝ�gg�R"'%il����Y�I2�1W�u���L�]�ܔd���&M��k!��X$U�웭ש6p�:Fߜu���:�ζ����2�}_��@��Yb�e����Ie,���#s�U��:wN}#�Q�\>�y�F�Kfܽ�ֵ3l���x���������RG�re�ٴ���F>s���h��6|C��fZm���c��Rlz>rdѡ���n2:�)�Ӧ�4x��N�礳�#��۵�Ӿ�,75��cd�9�q[I��P�@qJ��t�9�cFm��r4��尭���I,�s��4�s�X�����x6;����}�F c>:S�=j�o*0h��~!�G�x�z�OwY�Nw���n���M�̚x��[:�zO���W
�]��<�!d�&�┲=��q��ʺ�[5���Er)%���Nt��*�$�M���>�ڧ�[htѝ3������~4�i���Kcn��>_�t�.�/9.���ǁ�.蛝�!=��6=��V�I$&���酼�o�?8�u�~:�8�-�g8��s$�3�4��{Ej���&^GŜK9
=f�I	�4��Ʀ=vy�.·h��G��#0��iK+�\>ioWk'V��-u�D��s�îG˒Wͬ�z����\�%~��=>�Nx0��'Gf���$�Q �?�!���j�Q��>i��帷�yǖu�q�[m�;1�E?,��	���H���Ig��Vn��<v��6�3x��8�J���C�-���)7�"�A}v�W�c��6CvH˶w~!�O�y[r�o?T�`ʭz}t���'�g��>��ZzCu�-간��� �.��O��?*"�W�����:&	��0ᣅCYF�]�[ު��5�$���n��k�\�������~�&n�M#B�~�*C����S���cu�������������>���f���>���G0����d��L=0�2[�uE�S�:��6��2�I$vp0ɗ�_�������$�)e|ꪫUf�a�'��]��������A'�?�vNSMqQ�2��~ť0��o����VjƏ_�K$�h�e-,�E�h��M-�$�F��$�"4�$��D�$�"&�"I4h�DI&��4DM&���$��M2�$��I��X�KY�$���$���&ZZD�id��X�4�M$��M$�Y2��%���$���KKDI--�D���4��%��&�K�8�-)$Ѧ��h�--2$"��%�i%�ZD�M,�K$��G:�n��Z-&�BI	�BI$�$�HI2HI!,�I!$��$�$$�BI4�!&�BI	%�L��4�4�i%�L���d��$�L��$$�H�H�G��N�8��d�BY&�2iiim&�I;��	$$��I�F�ZId�i%���"M"M"Z-2H��%�KD�&M$��KD�$�,��Ii$�D�$�II&�M$��KII&�ZI��MZ"ZDi-$�Iiid��mĴ�i%��,K,���I"Ii&M$����X�I�Iid�%��I-2H�$��i%�Y-"Ii%��L�"KK$�KK#D�i%���D�-$�I4�DI�I-$��D��Gn4���KD$�id�%��$��F�%��ZI�$ZIi$�I���B""D��"ih��4I&�KKI�i��DI��D$�4����Җ�$q6�Z&�--"e��ih�Iidɢ�KKH�h����M$��I-$��id�d�I&�M&��Qi��M���Id�!,�K$��ZD�dKH�K%�CG#p��4-�cBcB�ІІ���lж�	�гd#d!���l!6�[4s����1	��4&�̄̄�Ba����Τ��u6�L!B�!l��ж!6ИG��ЛhX!`��B�2Ѝ�����7�2d-�,!�LA6�m�[4&!B̄�Bbdd!�fB�!3Bb�:�pHi��89�4д&���BB�X��� �,�вBB4$-	�YB��D(Z5�5�#���D�""ȑdB$k"D�h��-��YD"D"ȄH�!4�D�D�E�M�""ȑ�H��,��h��$H�4�E�"D��4h��"h���8M"h���"!&�dH�B"&������hD"4H�DM�"""��"4���!&��4L�����"�M�D"dM�"��$Z"(�"�4H�H�$M5�ȶE��-&��Z��"�h�ME�m���,���h�&�	�"h�	B"ȴZ	�E�Ț��#M���["h�h�4�4Z,��E�Ț$kF�(����"�Z��"�"�dZ$MF�-�dM"h�&D�h�DH�ZBО�74DHZ-��ME��dM	h�-��E�#H��BhZ-	�Z-4-�FZF�A4i�4i��BhH� �D�К�s��F��4v�ᦄѦ��MдM	�M�d&�К	��4kBhMb��h"-Bдe�hZ5�h�E�4-	�&�д&�;�u�Bд(�D�ЈM�!4"B �4Bh�D&�"!4&�FD&�BhDF��4D"	�h�M�MD�д-bF�&��g4&�hM�4Z,�h�5�Z&��4kAh�&�E�4I��h�M$�i����M�ii4�h�5��D�ZZe��Z&�K#M���d�ZF��{���s{[ώ|\�4)�����?[# lY�b�����|Σ�>���k��5�}���i�����?�Y�N�o���N7����
"/�7�l3�����ŧQ����h����w�M�G�_��X~U�����psZ?�������5������:�� ������.W���� �P~��	���{m�����1p��'�?�1����w���a��)w�a�F��C'�����!��~�� ~��**���)�����FH?������lK�� ���"�?���ą�zs���D������i�k��\�ħ����!&��c�XLG2�@?�S���u�'�F�AP��e��Y�v���:mͳ�����fڶ|��Y@	 @��H$t����Q*��M�?�[��'�(��&���:��"F�
$����`ƴZ66�H��PfYR_������t�(����b��N<7��`�������[���ߠO��+�I����I�TDY�����N:�� ���~���B��O��Z����������gd�����!�!���������@�D�n��`�H?�|���?��~U�?���~��cg����TU�K�`�gW�?r����_��O�N����!�!���3��ި������+���5�v'��h���!�������|��m���6#f�2���ӕ��HC߀0���G�)o�*���%��h���2.D���iE`h%%��SG��{��(�O1G��L�N)r��П@��������p��������?��ut���?�eO�b3��o��O�Z��?���������2X����#��~wS����/����������T�2��#�����Q�����EP��O��6Y�dD���˷����P��YYYZ��������eeej���Օ�++VVVV��YMYYZ����b��jVQZ��[V��VSVVP���Y[SVV�mZ��[V�Jյ��j�j�VQJ�+jejՊ�V�V��5j+)��jՊ�b�X�V(Vj�b��V+��b���m��X�V+���MYX�V)�+��b�[
Q��FV+j��VՊ�+5mXV)�eb���5+QZ���e2�YEmL��Vjղ�J�e6�Y[VڍEeemL�[(VV��څe2�AMEm[QZ�jիV�Z�ڊ)�VQZ���mEjjը�Z�f�V��VڶV�QF���jjڲ�E5b�V�e5eSR��B��X��Eb��X���()�l�V+jj�V+j�X�V+55b�X�V+��b���b�X�V+(�V(Պ�b�X�V+�Պ�b�V���څ5ej��jյj(�Z�j�+(���
յjڊe)[V��YMYEjje)���QX�E�(����QYE��VVVVQB�e(�MYYZ��5j+QJ�E
(R�VQEej��QYYYYYYY[Vյee5mYYE2���������SV�����څee
�Ք�ՔSV��Օ�eeeQMEejj�e(�յ2����V���Q�P��(V��QYB��+(V+jj�B�5(VP����)�emY[(Sj�Z�QYE�����mL���Z�[Vj�Y[j
ڊV�VPV+ڊ�b��X�Ք��b�[��b�X�V(+��[V+j��b�X�V+��b�F�V+��b�X�V)���b�X��)Z�jڙEe��el�(V��5+Q[R��e(R�+e)�VVQ[VQJ�+(�Q[SQL��mEe�VQYEmJ��J�Jj++j�VR����B��ԡJ�5m�+(R���������Y[VVVP�V���YYJ����++++)B����Q�)B���+VVVV��YZ�j�b�mYZ��ej�j(�[V��ej(P���5jڵ
ښ�S(S(��S)MML��V�L��JbBE�<�ˇ�y����?B���D\���?�I�O�N?�?Xy��Q`~����c�TS��� ��E�,����?��<��E�3�z��J�0�<%?�)��ἃ����S*��:O�%�̒S!��� !��Kj��?+�>�������~��|��H���fB��`�~��������等��mf�z����"?���ht���8"'�OԆ��7����Mjm���������O�~x�BؕJT�~I����H�
p�`