BZh91AY&SYT���߀pyc����������`�8��     @
   c�     
� �@Z ]� @�  ���   ��wu^�v���Yu��(� �]�ﯾʺ�c{��v۳y�H{=�  ���}=9n����������Tˀ���Mh��C]�k�`c��v�]&8 ̀w�5�ol��x����f�ռ2����|���D�������A�u��8� � ����/�v��h�� �n+������Zh�{�Z��p  I���7���-W]	�>�3{��`M���vΰ$_^�H�(        7���       4�~��UJ4�	�&  ��d�HI*TF �& ` F�#ɄE�I�e14&���(�	��6����
��@*�OA2=��#11@H�J�#4�0	�@��&�L�&&��zI�5*��@ɑ�0 	��ɉ�}�����7�|B*�o���dTU����"*�y܀����Ni���	�OvĔ���m�6�n�����s�.U�{���ѷ���R����ٟ��-��͛�ϖ�/�|����=�{4��M�,�s}��ēy7���p{\��l���m�	�mcm�m�m��^5�<պ8%��3��ȋF<5ƚ��D�y�S/#�����g�ŭhCF���M�m[n���`ލ��j%��t�7d8-��x�tLEC���d��LDb!�6���!����1��v�L���kuƃ+k[��Ѯ6�b*>��kw*a\cy-<��Y��T[z"1����9�^)x6��g���~dE��[~n�P�uP7s
��4,j�4xs��wn���8�%�S�!��F�񭼆d8f����^��5��",v7Ÿ���,��Ӛe�. �\�Q0�n��q�Z���*}M����d[��`� �	�7�O\F?E��r[���K<�m��l1l<l�p�k�e���j��qT�Ω��ܖ�(בn"�q�ُ*!�C�ű���!���C�z��[-�X�"i�6��Բm¶*h���F��q~���p7����[��œ�p�F�x9�ŏ0q��ߛ�zc��ccLq��v\E��i����[���lM��CQ���:��cwn*�ŷ���7����q�2�X��c�lt�_��)�(�F��f�4w���p�������t�cl��\�`�.3[��c�5ƃ��D��C�/&b�7O�ōZ>������j��Cd81���@:�[��:!�C����z�"C��:���8��2^�XK�!Ŷ+o#�vꌗ1�8�q�����mk��s�Ӹ�v�f �[�[�G
eο(�U~p��b�qY�d8����!\�U:B�b�8G�I	���hnؼ'Í���'�,D<!����W�C�����O�G� P8S��]���&#��E��R�¬F=Z�b�r�y�bѧ���5�hSokR#\q����C[�[�r���8�E��1���#��aŞq~����-�Kz��#��x��kG�԰g���^'t��N-Qn(���<-����5Y�,
�qx8�u1�j��
m��8G��m�6؞6��b��(lT��
�q�����E�)�"�{?8�h�88�ZІ��k��J��c�*5�^�,��V����j٦���৪G���'�V����yP�P��%;I�Kԗ��IX���	�	���?-NT�NDЫ�_�&}cv��M�Z�Z��V�T!Ou��d�PRr��А����L���js+�&,�<�:[����,^>�kLT�B�N��k�lQ�B^�إ�%�i���B��
�LX�VС1bv�z��1_�Ŕ'����{i�-� X�R��QlLZ/"ԣ��(�P!m'�D&���]�oӃo��WK�:=6cWq9��}�?C�_d��7��<��?c�f�"7^��kf˄SoUk��R�̹�+�:�[��DP�����wpɈ���<�D֋w�Y#yJ�O0��N�T��6�W�N1C���j�z��s�gڳSkuh��C�>�����P��S����[b`�Th�խƞx^���D(߳��3�(3��H�l����e��n����Dc{S�ˑ��������w��6I�����>����
��Uwp7�]!cZ*j�9�8�Sj�y��8�%�M�%ﵷ�?|co!��<P���5�����8�{�r|�M9m�9�[2�eˊ���M���לT�"��_ȧ�]&l�.� <����Q�1�1�[���e�ޡ��)2\LDa�eC���!��Ǫ�y�6S����Pݨך��7lW��:����h����!���C�C1�"�[n��qN	��z�*b��ﵹ�Q.#]F8�C�!���p�zݷUbm����Ń�wn��nzc�w�����n�l��o)~��p���1�\��sC�X�1��nKpc��/c~lo[�I��o���y���r��~���b�:��B�2�f�G����K��'=L��m�k2iy��`rG�J��]ll����p:��oNai�ۍQ�`�)����Ŋ.YMR�<#v�ˤ��!Et��oؒ��Q���R�>�Ks��G>�8�uga|��[�qڴi��nac'���Y{�7̈��%G/a9�,�W��l�wO}�-�g�T��ɓ���^�<�.x�F,�/̿4�O�޲��e��.��s$��V���t���������!U��TJs�!���Y:��j�p]�79��'�9���	�o4��إ�$���0��U!�Nz��Ÿ��S{H�7��-g�I��zAK�[�?��H�֎�"���#���g��3͓�8��'�7t��L�d��o�{s����;�������/i�R5�g�3�h��
i�cO�'4i����G���y�ﴞ�{��q�C���m��S�e7[u
9��G'�W8����k�y�Y8�h��<���
�=9�]�q	��=��t9Q"hw=���u�wx�9r̬[�ۓ��9���Ν�8O���V�f/n&s�棾C�x�u��k�D����I�������:����>��g��k�lU�VJm���×����i~���>������|6IS�2�p?�(?�Uh�h�����Ű���x�S��Ni	�}�Ԝ����ʡ7{r�7n}Ҝy�[�Ȅ���aȬȢ&�Yu�4���v��見�g�Q8��������q�i_-=��q��?��N��p��\�t���i	�~��)�&o�*���z��,���eh~q������}���i`�zqL�>�t[�v��[Kr��&�����Ig�&rY��û�9��>�6�v��;>�ҏ�u�_$�e�LQ���������sN�rg�j[�I_��^o��{Է��#���zRgw�ÊQrv�B���A�|F�Bq�Rb��y�_/A~|X�G�ٗ':mO������Y=I7����}������J�(�u�}q��G��4uuwZ;�a�7�p�]X�U��X��G>�Q/��(�YE����"�>2q���y�C�5r�Ǒ��d7�u��B�R�!y�|���H���X�uE^�ܕ��=�ߺ�qǑ�qG}d5i6BK�lO�C�'�R����Ӹ�:�Ǒ��^�sF�Y�K�p�R{��Q���	�;ޚB���h���d�`�G՟#�ˉ|Ks�}�/3I-����g��/����%�$�W54��*�r%�3���P�l].��ruz�U��g��T�]�5q�|��_;���:�?��}"�i)�9����'�"P������-��|�4�-����j_tuF�\�?t}�3�ﵿ�b6.V��NlK��J[ω�z����챮�g����#�{�!���$��v�����D��.�f�-U{S�s���5��1^�8���/��"��iD�˳����ĺ?oEY6��K����D&�j�9���V����Ur������E��um������N�*?_�U�N��ip�Ϻ��>o�Ǡ�q-�)q��SG��=�P�Y?=�z8���ӞϏ(M<�\�o�׺�̷�Ov?���9e���P踷[�;�^��:�[��%k��k�n��^m��&��6n��5w����~�"��?�6�}��nXn�H�z����}~����|n���m�w��z&���Ww�����^�l����ɼ���_�<�xʭmƳ���#�j/1k��V�������4�_��NK�o	t�*���r���bG
�6+9�՜D\���2�����z'��I����α|̂�{�g��>3)I�O�	xo�d�E�2gY|�m�=z!��lR'G�oQ�7��i�����{�>�I��=���3E�s���Fr���/�'�~��C��	�a�_~lN!�h����~?��RI?�c���z�g?˞&ӎ՞����2�W�T��������j}�Nab���j�|�T�����z�mO��I9{�N�ξ����Q��M.sm�[�$S\DԪ�+7���gY4{�����%U�)�R{�W��_��N�-i>�p�9\;}�#�}�9�؛G�)ͲN�]n�\��Wm��sD�yi�dU��gz��H+*;ν���'{�wus�zj��;��uc�N<��x�Ik��Z�k:N����Z�k޷�]ͷ�\�ڙ,��B�>��h����_5����ŭ�V��G�̻ܷ>ܪ��ݖ��`��r�X1Y���D����$/�FA�����?�����C�ǳ5dNJ;Ul��a�f�Q1eń�x�HHI�.�&�ZPX�Bo"�$K�R���J-S8�4���k����*NOi5�"!�UJ��ֵ�m	#�ۗ50��In҉: �8�4�J����N!��Ľ��1�.`��&'��R|�r�T����ʓ�屷e��-⑸3�A�,V�!WebE��ګhX�k)[z'i��*X�]�rJ�]�_{s�=��P�j29ig��n�r��J=��"N�&ڵO�5�׵����%
�NT�W�K�NF�q�����-htD���RA_���<����mC�5,z򤩮Li�"�)�m���?H���\����ҊG*s��nO���Iq2%���4؀�V��gSJ3�F���]m ]eFdX�a���eQ֔N�M'|H1uD�<r�鞹T�^S�5��Ґ�[�dq�'"M�%��^nq�u?�:n�U��(�T$�q'0C+)`�6�춅G�U섪�BȂH�j��o�ܨih��p��i�'[vd�'��٦�X�*,�������,�(�+�E�����n��E]����e�7�*Q�u��(�4�I�$�ɂfNUѧ�Å��;{��;��ڢ"��s��	�r��/��IZ�P��w��I����P�D ��=}��m��w�x�fJ � �  �   � 0  ` � x ,A32�     @0 ,  i�o���6����������� �<઩��< H@   �` h@0 4   � HB	�� �  �`   ���� _/�K�1 � $���0  ��� �  X ��b 
 ��́  x , � h� �����I|��wwwp T��    �< H@ �� " ��2g�  @� �   ��%���m$�� `h�	���    �� ,  P�	 (@@ ����   �<  � ����$����T��@  �   � 0  � 
 � `x  �3*@ #F `0 ,  H f��i���&�i��G���2�v�x��L|ݿ����_`%J�A�?%�~�~���8p�q���u֜:��\u����:l��Q�^:Ӯ��N�ۏ]uǎ�뎺ߩ�Zw�˪S���N�:�8u�]u�8p��ÇN�:u�T����Zuz��7�/{����G<�]h�4z�{&��X�1�j�B�YK�d�;�3Q�%�X���
�8B��򲌅!QH2��q2�yb�!JAk)H1�g���ʍD�S�R����D����bN�9"��Q*�؈Q�2Q�H�RCVL���.<�C#@���(�j��1N�,$4�Qb��bY�M�X�!b"�B���S-T1�C�8�(�m�`���r��PT���¢j �H1�lL*+`�r����(���d��	�bn�&6\X8*5���
��!
+,��E�Z��[m*�*5�M&lI&�4\n���Z�����D�1X�()M�i-h�(��NJ�ɅI�,���ծ!���Ұq���� �6Seѥ�S�lU��m��Q*&�<�U[�;u[b,ɒ����6�H+u7��Z���NF�!\I�Z����%j*;cB��D7�M�8�?~��#s~~����m��EjN6���J"2�'*�b��U��<��Z�&��i�չ+L��[kl�U6��ku��*�H�K.R�l����E�V��)*o*Pw�-�hD5�$�M�*�H�� �kMXH��ő֣�q�%�";)UԩX��$�N��u��"h�G(���1�Erd�n'%+i��(�R��'�Qb�ke���@��K%�u�uʭ�,o1ʒEDjA��
ȕ+���t��ȑ6����L��1(��˲��;��}�˫��9|��/����{�h���K���9$���wu]�>O����}�u��Wqϛ���1�c4�E6��m~��򕸌�e��m�$d�DL� ���t�)U��*B���D0BP��1���:ZƱ����)�"2�8��DU�J��ǫEKUl�������*�Q��������Jڪq!T㎅���b��J�1�ȁ �(�\[!	�k��m�I�a���A�蚁 lwL���4Hɕ�pw?g�L��<�ˁ|�嵖�Z7D\B!$#mE#i��)��7a����(0g�3��������y��� L��x��3ЊBB��
gY��M���[ީ;�k�oY��|��:�0a����qJI	icm����Ł�����Ƈ�o��ˁ�衃Q8CCE�>�"J7�D�p�E�����]i���t�﮴���-D�oٌ��qh��@5�o����FB���1=z�t�uLF����2QM�֙h���x������Uuu�ۢoE�|�%�|�V�vB�ӥ(ƕc�/c���\�zb�{�Qe�������M׏s��7s|nog��_&�D#!��b0dä44��p�g��u�qV�m�mܰ��7�%q�Q��:l�m�oV�q(�M��#��F�"�� �RR��\IZ���-�R���b3�c����iG�l�NG�`s��v6�d�th::�j��K�"4ӱΆp	�ŧRIP��:l�!�:���{;F	��e�O�˗9���^ޒR�������x�|lu{
jj�E��9��F��i1�������m�,5�֩B:�U���g!�OB6=y�����O�7����Nj䝛�V����.��ǫ���o��疛��d&[u�n�ΪYZ�b�V0Z%O\M��L�3>�e�c3ح3���&��ڪ*��0��I��nF�(�f1�S,�Sh�L�i��I�7�5��Z�o���}r]ۋ8�}���i��6��I�D.|�wRH:kjXǔ�<uÇ�*��{�I��������ӄ44q11���$�*��[���W�P�����:���J�q��n�+����o����#I�2Ȭ�*1<�
\�ر�B[��B2��	#Q[AF�h�I��s��س�|�1�MK��6�^r�ScT���Cn*s�FI"�F�DL���r�n~� ����0Rח%���\��m��w(�k�Á�;b�g	��I�6Y��ҧJ�#A��C�&G"c���ײ������H�$�(�"}�14�3s�:X��=y�zu�Ʊg�)���*�Dh��OR%�:��H��ZD�D�E�2JN���J|�&�h���-)�ZZc�i�m�[JRZDYH��-1iI�ZZnM�2[j��j��:�Z�:����-j�U7Rմ�j�.L�l�g)d���Y--N3jU�K|���e"\�"�ԑH��i��'��$E�%�%�%���J���i-ڭ�q-�����������,~K�o���-�.j��G�y�y{��],-��o��i�n���wS��������הz,�wˢr��/έ��C���Is�ɝd~ӝ//��滽g��O?��k�UU׫`s;�ﳞ}ߧ�����u��WqϟwO>뻺��>���˻���C���~�����>���]��]۲��X<�4eH���-���R��)J�M47�*�� 84j�8:0h�O^������7�m�]�3��i�Xa�������ߩGd�D�$�6XB!��A�A<0^���֛��=�7麙ɷ�����N�w����=��[�mkY�M@8����88J͒��!,�8�����yum�wkw)JR�@�CtJ�n[J�w�E��'�8���c�,���+��	bUSwW�{r�s�`n	�ǲ�NP&�߀��������0lo���Z�5���ɗ7�<3�~��6g�t2Q	d�q���S�3&ީ	++%!+R��C�N���J���E�*���(,�6���iKKU��V�r9	U��					`&,�� 1�A�cG2bQm$�G1�c�&*���dō�"�$���q����ogF����fE�-���SB^^9� ������x4��|4�rpr6�]�5���u�T�\��TD�����z�����y���U;�}��B�����(�wf�ʅR���|�žw�w���\o��۰\`��.�X� vPGZKP��TVAX�4/�}�]~����[��O�����]����*�U[0;��o���H�6ǰ��1�3���#*z��e�g�[�)�_y���|^zR���6ї�X�Mt<>Ԓt��Z��6Ǯ[�j�6�п1����q���$�����%l�I��C:<˦��p�S��t4L�x��������G� ����M���?&�,ڑ�8�޲ѳl�0�	�
F��9�`�����^I�m�sv�09��q��c7����n�N��VԻ�8!��0<��#C���T��l����i�'F�[|<�P��p=q`g-�zƀ�T:��>]��4p(�1�!���������C����$�,�������6���;�-��`��WP��Ӛ.q)�,LLT�y
�0ַqL��i!`:���(��E��I�*A��'L�8vݸ�VP<��+a���$���5�U6;�Z���7l���.!a[���b�����9��LHc�b�����h�$\C��dn�����1)y�����q��X=!��E���Ϗ`41��jUZ*��ip8�<=k����d<87��F�۹����a������N�4���T%;��L��49\�
�]��5�$Ł�4����*�o���B(�z4��І(�%�>,�h4WL�n.
�Ŕ�0��&0	��~�x怭��`YM��^:j6�����4�q1�5��b"⪨����[,	+�;�+:�[ϭzo����7N�}n�j�
A�c۠)�M�����Co����UJ��"/�g#,�O�u�^6�S��챆��|�ƺ@>m���󗛫�������L������lb�|�����8��a��
����س��-�>borجg.$�$��:�Np(Aٯ22�.@��x32�|O��Q4H`��6�8�:��өԉ��Z�-jfIl����>O�I�c��-��mE����S����c)�%�h�j�jܛ^d����ҭ�N��J��Zuj�[�z���Kgi��Ĵ�-�RY�ZD�,���ٴ���Zm-�u$KLG�"&�IH����h�iiV>R�>DO�(�+h��Z2�i�iV�L���Lu-8S�oZcm���q�!���{��^�yi�] �D�a���\��O'�_G�8�O1�[Y|3t�]#��$覈���i�����>�Q/�1~;�/{���F�.��s�MZ�u�;��)	3��ػ�k��;7�sb�:�����3�>iJ�NR��T�YY��g����1m�w���C�E+�촌=�ys�R�:�ߥ��u9�_��9<ͨ��m)]����$�q�H�~��V�����Ҫ՝�����t�&,����c=��&�~�W��#_<sdPX�������ks���U"��g����DȁM���=b7k �V�kc�\eHK���"�ޯ�Í�-�F��e���h�rF�4V"ؔrJ�"U���V�a5�gɋ��mT��v�ަh������z���;�?>���˻���C������>���˻���C���˻��寻��Z�{���ܗwt��4ʔ�--���~�6�l�ALbC�ȫ`�<yI(ЂX��FE�ʙ	�Bb���8<�D&Y���d�J�,A*�H(KYA�hV�v��㊥J�ؘ�+%V�� �8\�Y5�$Iҕ�[���r)-I!8���ȪX� �Hv���UU�M�n�c���B:1JL��h�Y��*?��n�5q���4j��KI�i�l���P<f�C H���2Bsyt��\��`PGc��������vO���ث-���]��H@4>�b�ߜHM!�a �l`�`\�vʺl���Gz�J�)�q&5����T���[/��OЕz�����`lm��y�5�<m
���V���>��) ���qe���R[5%@���� W��K
B[/5w�y�q��'���h�6�k}��H�������T����ӳ��:Y����J:��r˜�A81��p�-A�o�狠-�>�6�j�fv�B]]*eؕr�J�`[����ޟQSC��^�|�(�Xq �v>r�)�R|�3ba!������r�c{cV�:F�R���̼6y~�����ou��w�Q+~;m~����!��ۗup�섐��Ǯ���۬P�����xZ�pf2I��8c�ȗ��(x��Ӑ25N.�*T���i�����gƱ�Α�*R�[�^6�Zr�/���"Q�/3D����9ur���5I�q�5�wx�
��R�,I)�#�V%*u$B*)�-ɩ�>6�+� ���M�i)cQ�E"+,J6V����ϬsM��/:��۞�:�
S��nE���Otx4?6�Z|�l��C��C|���C�j���8x�m��~u�NW'9W�^x��G���x�ݏP�[O�:d�B�C�ύ�`4'!�c"|O��o>��wsm�$���J�_)�J+�@��C�����?r=<�7^k����k���� ݨ�mpXՉ%s��ǛC�� t8^*��J�Rɗ0y�����z���I
Ƈ�M�(��!C�k��g��:������V����UT|829��hk9�Ħ帆1HLLF�	MqЎ��(mB�#��~B�z0r7H|׈J�� Δ�b�}�Fxc����0�,��e�g�	� �4�+d��~���Cަ�B��*BGՔr�v�hxm�b^i���X��`�iHs�	�v�UU(��p9��4��:��G�P��.���8xE#/���i�r1Ԉ��J�BѹZEj�1
��"X�s)2��ݦ�V�rѶE
�TCQt�[���h�.A��4���jm�M�J��M5VˌYT�ю��FB�3��囟$s:e������P���)�Z�>��<����tq���2�W&{dݏ2H3a��mRz�G�v�$�* ���$_1��ۀ�q��We�nF޼`�kAo��0PB�S�!��(p8/�]��8"cx��� ��z��=ve��sl$a�;_5$<�A�C�,u��7ٻ������o�������q����.X���i������z��湿[��KC>hz���Ч��~6G�T�-"x�X��ĉ�ţiԈ�DuN�Ғ��Z���|�O���|����-�mV�Lm2��%�Z�&)"ZD�Ŧ-�x�[j\��ͥ��v��n�iԴ��Է�\�U�S�E�Ĵ�/)Q,�E���%�T�V������Y�e-"Z"x���DZD�D�D������2�g�D�򏔭���>O�M+�Ų�E�χ�G��D��x��|�sa��uI�>��d\ۏw��q)��<Ĩ��ۛ�ˌ7=�.�d�������յ��i'������hJ�w������S�~����$�c�_��7����K���k��{��r]���Yww�ܵ�wwUe��wr����U�w}�˒���Z׻����˻�e��4���A���T���v�FIk���:�@�a��������l'J�]Y"9"pbM��w?3:eB�Cv���L�xp?4�!_4>()��sV�D�0��a���R2�2�Ǐ�h�s�i����)>�dx0tp���N���ֺȊݪF�Ges?�>���fv��Ŝ�$����0C@�=��\������Hm��sC�P~`��!,p���Md�A
!�%�t�H���ƋF!��K�4��֠��Y-5�F���"��7R�+
G4�S��28;U�ȤvA�#+>�MB���
ɑ�HNVLQ��n��U�x��(Y#&Gt��9z=l�9�v�;ƍ����r�9��Z�yo�o�[���gN����?n\<�p�h�D7��|U��w]�v�θ�9��|�U����m��˘;��A��FQ�Q����F��e�������a���Ǿ�[� �#�68pD:@t9X�4q�:�Ǻ�1U*cA�(A��P�x�$��sF�~4�;~��`l����\+׈S��"���q���n��)O��r$V�u��ǭ����-i�u�{�m��w����_��Zݜouu��o�M����9�9r�D���֦�nGM,~lx1t;��6�;32f�4�ܒǌ�<�۳�R:��u�^�bA=�y��&q8!c��$���m�������s��O�,V���B�g�x�VwsC�����vwƪ�T�,rw�� �tq���:�]�$��~vXh22�����Ѓ�ޑH��\S�6m�߸�Jm3^b�Y*�E,�@�Ð�T�Wɕ�H�l��r=)�1��1���2�lN̘�%�H��Ң�I�G�����|<w��� �<�iq�s-��YH����S%D�Ki�=�g�N
��;��"a����
2HLp�����p���24�˷#C����?F���;>��L�����+��ή\�q-��[�����-�����E���Q�m�������x���"��b�V��<�i2�÷�h P��lyDe����W�ݏ��,:}���CY�)���=#�%r�ƛ�261�ER���noz��_7�z7���)�l\:�94Q������q�o��g^C9�g����	CC�ca��|��0L����ɹ��#?	|1��85BLs*b��UX�ͅ�qA��e��r�S�0'�[~|>�f�= 2��|��!p�ltPۃ��?
#�=uCf��J�J�I�yY�=?�sz�������C<7Aӡ���4r�3�J��I�7>7���w�x�md��a!�0����<<��9lp&�OCBͺt��/!	<��'G�7V��]W��t�ʗ�/ڼ9�%�K�ߓ��������H��h���Zc��>q_&��O���b�nԵ:�WRq6�]I�%�����%�-1i���W��ꖖ���-�\��iի�n+��ږ�I�j�-2��TK%�d�Zuj�*�����ȍ��$�����>)|I��/�O�F�)$��U%�.�Z��-<K|��r|�S�T�#�|��)�z�z����؉�S�G�s������3���$��)�ԑ>�6�)r��D�Q�nT�ׄ5����,hC��H[�ka�\D��rR�Q���Q���q�-rYQ>\R����%͜���7��Z�ڞ�boe�n��m��g:������zH��dcXNE��.�7�u�ɒ�a���퍨�9'��h��5>M4���;�]��ȒV��5u�NX-{ӆ�EJn�S��Zc[�r]G���LE*�K?~�_>�z/ͪ�]��Ï<u9HI$�H~Y^�<C>��N=/`Ć�DԮ�'�TA�ڭ9\�,c��/5��u�O\l���n1J�&���N'D�#,��j^�[u�C\N]Ѥef�(4W���s�_ݙ����8�k�������������˻��ƻ����.ﻻ������k���Z׻�������e���]i�}���TB"�4�YF!�-!���	h��A�lK)yQ�#���'Z�WUF��\����РZ��24�Tp�dX��b�eqH%��U"r��")j�Q��)��"�E�;(�%vRD���
�h࢘�$�C8g�G�o����*~<��p�����~շǽ,7����`ef��rB��%�f]!�3��W�1��e��^��f�#X����r��:����8;zl�B�l�&Nt>_�ѨH���$��ra������
�p�69l29|��h4��G���J�R?{����#���x�*�=9���0�3��04���{H�c,|(ʑ��1�f����[�[5 ÉS���Vв���0m
��kC��#�i�R����Έ.~uÍA�%���iU�S1l�K�u�ŋF�Q�A��8�C�|ǹ�v�.�[���V鲟6y�����ic����ϰ���#Jq���NT�fIQ)�k�8��l��v6�e���V]�q�g�|zߵ:NU%�v������oy٣��|��(Ѡ>��$���@B�t�Z&�c�P������#*i�э�yN��D����Y�X����g�[[[D�%�e���V�f�:�ER�+J����f�1,���@��`�0C���+\�Hdx�7��;g�c��N����xo[���p�\BO��4m-�����TIU^p} 6����8xr�8�j��A��r\�u���yo;������Qm�9�'CE�G�����w�6@�:Ox%�aD_e4���FX7�[>r����C�Bء�^2��fY�g)Fb��㏎���'QᾹ-U������*��|����o�G��UWO4�mN��ٷ^p���5�-�c��qCao�i���c����gi�Djf�U�G�,����q���V�r�T��ݼZ{>��gF��Յ�w���3����z�4��#�xӃfڹ~y)Y��1����V�&�����|��J��t�!Yc��L�K>6;)�,9�~UK>���������/;���^˳�����/����҈uM>ll�x�1�ןr���<���՟y���R7�U"�
�ز=�ee˓�ڬ�B�Ⱥ�Pʶ��1������KF"n�(Җ��R�q�6�|��P�37��C��:�*J4dpF>�$�|���Cgç��G��j���"�׍��}������+xd;y�~j;$�
R6��,l�7�R]9�43S�#�m�3et��V�|4t��0�i��I$1�h�������)�1��G-�ж�t��KH���n3gE�t����˖�[-R$���L�x���~�ӡ�����)}�x�T�TO�	�D�z�-"|���DGR#�$�DN��I�uJ�#��>N��)�q�-1iթ�z��E.��i)�i�����m*ӏW���KT[��:��Z���]M��i䖪x�O�%)j�d��e��KTZ�-��:��:�JLRDu"u�":�$Gɵ+��Z"Z-J�1i�ZZ4�-=-X�Zuju�S-u��|*ދVRZ�h��?_��|k1��zy�������s)��w�̘�iP�=�+	V��w1��B=��O��=�O��B��U_8 [���J�/=Oz�U��ҫܷ:�n�8�k�����.������ꪬ�������ﻺ���˾�]���UYw��˻���-)SKll������1��G���:����xzh�F�"������C�I.)�Z쥟��#L�,�fq�OOK-��$s��C�BO�����]�Zv����޺s���1X�x|e�êG�z�cf�c$��S�w�칒��� �mΆ�T#CbhLmc~�)N�9�|�ieU�ԣ3T�Z0񹡱�ÁM��L;xtp9~��4v����oy�y0���L����ɓa�p��� �p�����Q�jHD����Me��k]�v�42��
�l�1f�47*U�(�1
�,��34x��$�J5��Q,RѺB��m�#Tj8,�Ι��C������t��p1>�B̰ˊ���7`cYk�}i�ռ��ID�\[����5]�t�u\�492e��G���o��S�66m��Q��3�)0�t.F5���;�S�w�c��Z��G���!�˓����[[�
�Y$=Ϥ	29��,�P��g���RI.Y%N�Ԫ�+�BHIf���9������Hȣ����!(��p��"�6(�J:p���]�t͙6,q#��C�� �6�����#C��:��4I-mF�H�O�c�Ins.c�];c�f�}ʔIGͻ�x��v<9U?n�{k}Z����|��������>S�6�z[o�C�"�2|��!�̫ �Q�<i��g���/�H�t�rL�ܻ�I ���Cg� �0�{�`�wƋ�lp?4�{�Lw�����3��Q8���ٶ�c�3�0��e����LDRH	IJl�G�Z6s�ebk+"L��"˔�l�()������^�ݩ�2B����<fKX���ce)2��c얧+*qe��T�����o:>��I.�fU�2ڔ�����:a�М>	 ��4:(�úpeH�~`<Ԇ��j�6��U%T������$��;rJC&�8pxfKJ0Ce:h����=Idj(Jк�|XᵣJ���ht!�ݞw�Ld��6GF�p4u0&�S��	��yf�<~pg�Q�~�R�z�|�V꫾\��e�ǽ��~p;~�F&���nBjQD��L�tE��pB8w�������_���09r\���׭��G�!J%oF
%X���cg�h���[�41!��ن�0~���p��B���Hl�㦇A=
�*�-*��ݍ= I�CP����ߦ��*�1����ޖ�\�-VU��*���KH��3��!��xpl98�}�yf��2���2�6f@��!p`�ˣy3�(h�	���"''SjW'��|�)Ԉ�Y�IԒuX���u��)�x�#�i��|�eO��Z�G�i��Ԉ��-!-"ZD�-X�Z2�[J���qV�r���U����ի�n������KW���ĶUKR%��%���ZR���U�>DN�9RD�"mH��N�N�&>#�KG��jD��[*�-%��KR�թhA~��XJ>���ǟ�Ì�硹W�
�K�r�:��ޜG)�F1����ZO�	D�h�.e*N	�)K��&�nܙqR�m�&2���k9�4<�Y�܂�Ȩ��a~F�G��`�]�	�$QN���X�4Q�b ��M���ݩ������������po���'(s7r�Ɉ�" �RbVQ�(�,~c:�8��ǝk��*gi2���v&��c�2��_�MO�s���ɼ3�;��	!=UZ��SF��oܧ3���Ǟ�#��\Ӥ�}��;v,]�5lMV��s����\���ß.��jB:�kƍu8�%$M�B"M��+Sb�LM��u���}�.n�-|m����51-�)B��R�qEl�3���U5�U��6�Ncuԗ���&��j�I"!��G��?/�Y��w|uw>��������UU�������ff�����q�US�������ff�����w��)�P�r��p��i�TT�Ը�2�ܥ�(��CMvK���PzZAB�h�,ȊXL�5FQ�Ar�#�D"�QB��\�-,Z&"�������1$ˊ�A�T�1��d�R�F�ZD�*q27h��$���A6X�U�J�y*��9�VEH:��IFM���"�y�2[���$4Xڊ��*�I��CV�P�<��W�15s��L�H��8�*����z⛨Q��m�扢���� Qf���c@q���� PC/8��ve$�]r�N%:�.N�w���ouI�p��qKi�Dm��$yUY�Sp�FE�T���Cc�%8z}�ڱO��n�s7���jy��`�A��9�z�*�Kz��2���}�(��g��'.n"�Ͽ!�s�צǃ���G#cD��Qjmm�DFٹ��b�U1�Xɖ��J4��S����C�r�/:ΫdI\�6����A�RjC�âS���\�����F0ӑ�Pm�����̉)$���nC��xgƜB85�8�3&_�1���fh�m��)e���K.�JB�-�K+)��8CY ����&��G�N7��H�Kie�#TT�v=�X�����&λu��zI!�o�å�SO�F%��+GT㍛Dm�k���m�*���E$�[il$�c!A;*RB��W�r��uir*���W%�:R��14 E6�һSq��I8��(�"$@��3�7�9�����L3ѣl<.N�G)�j�B>|�������Q�G��{|zޭ�9��W-�ry듎s�!雝?a��.��?LE���T��͢6ֱI0��UL��d�(��C���A8���7��MT�fknCO��m��I$>t!�CǍ���h����U�؉����_r��!���:`�G����N�i��6lŚ}��>
4CE>4Nl�q�`�ʫ4-��#48���t�@�b2�Q%*���|7��tߧ��m�k9HI��er���9<6S�ݰ�+��v~�ׯU}ow�z�Nޗ��O#?�xg�9f�E�zo�ޙ��\�@<U��؄Q�F�ȆH���u3�)�ٵ˷^�"m�?a�sm�9�a� \t9r�!�/�E��C�t�F���em�ED��m�a���=0XQ�(ɳA��ny���$��c!LQEnd6M��!	���>QTC�dE��p�Tu�kT�jT�3-��f561�T���حi
%cl������2�6�:g�I}�������p�W��a���3��:M���۳�oص��ύ.7�7q�O$��8�{��^�1&ޘ�3m���!���4^F	%����M��(lك����c�7Ue�.��}^�D�8�-��Ƣ��E����~�M��iwW��Ρ<ӑ��I&2��=e�8z�>:�Î��Nq�o�����ks�Ɲe:t�#�T묺��Zu��=u�q֜u�\z�N�ˬ��T�ӧN�z�u�ZY�Ӈ�p�Å�t��u�T���)B��P�OR��+�ޥn��C�!Ykvv���O��<���ɼ�E�g}>V�*̕kލ�*���ݿ{ym�躵\~���=h����|O�$������*�%�U�&8��G�;ﶏNIJȨ�q�:���5s�i=ϻ��fo��{�wuL��wt�twuT��wt�twuT��wt�twuT��ww��;���4f���kB(e1f� �̐h~��c�����wC���q�
�K���}��o�]t?A�ѡ�=���MS��!���4,���t��IJ��f#-��;��%�����7�Z��_�A��7�2�:}Cco���r���3����l�U(�]��\�r�l�u��g�09=w8b�Έ:�:3O�����^g�R*��A�9�N��K�)��5g+��q:��x1E^h�d���8C�"�p�M��*�hJeRK
%r�-���X���E����#�s��;EV��cA�Ñ��s~o�p����L��4����d04����������6IE�K��)�$.yԗ�8y$��L�肊z�SO[7�{�b爒�3�6c�ֈ�t��	$������h1����v���|C`�>``~^���(���j�����m�I%���>%�0� Q$��w�޺�5ܚ�;�N�6S��O[l��rnb���Blp0F����vp9ͽ./�#���H�m��i��Ѷ��櫶]Uݚ	�z<
�!'���y��x:N���γ|i���˴4Sh�M��ft���3�|��U*�4�:J���ͽc HJZ�a�Ν|����$26hpX����\�v�>hz4��c�B�C�����u��qM�ٲ����k�S�Z(BV�l.+�&��y]J����X���:D,ID�B� �cA2�8��fǲ�Tc#vZ\0��c.Y��1�B,lph�
�E�����u��q�y�5���{�n�o{������;$���t�'�&���g�]�>r���v�2��L,��t�d����� l��Q�(�A�Ԟ�Ӂ����Ct|�??�����	���65��d y���[΂��gn�=J�V�N�vZ�����;�뛳�׎�ǋO�߈
2Ce6h4���ъ;d|��;��e�#<�0h:]�4�QTS!�cϾlz|ns9q!+�!b�G$�*�Cc�X��䪔d804/GoZ��lv���[�,>
<CE8h4'J��<uiq��m���7RYV("c?�B��i���Ea�8t8�k�$�Zk>p=]z+�/�ny^�(Ґs�L��1	��q�ۈ�f�M��8p��N�=q����Z��Է�n���8t������]x�N�ۇ���:�8�Yi֙u�T��i:t�N��]um����Ç,���]E:����B!P�j国o�*���U��9�,������>ѱ�e&>AG)�Q�Q(i�r��I�8ϝDؠ������4'�&�҇�3�#�=��9f&I�]Lg�(4mG��N���)�EJ�H�BW�H�B�Vv��W�<�W,�h�=��\�j�k��c���V�:n��1�[���"�	,�Rw\8ia�s'�4B�Bj�u�^���s�djRM��)t�1�Tq�%�j~�c��^;����1������w��_$��֕�>#��H�8�E5Ǿ�o�x�Gǌ���	�͏�����(�6ؘ�_Gع|����o�l�}���K�Z�\bR�$R	(O{�E����d
��G.ֵ��dr�U��n��(9�E�vB�HK���R:գƒQF��)zU��UK��71U�����S��~���S3������꩙���wtwuT��ww����US=�����wUT�gw{���*��P�5J?�>=���Rba� (��H�1R���Bd���QԊQ��!wG���� $PoB��bIĜ-�ժ;��9��Q$��*A7)��Wka��k��m�Y�ʒpYV*ǈh�J�QAK��(�Y`�Ȥ�5Tm<m�`�DB
���m�!2f��bCr�J��a.@��Hc϶�����am�C!�	Oǋ$�ް>㒥ITW^��/L�����zI!�%�	h�Q�%�a��?S>2�C�:C%8h4L��!F�;`�쐋M�q�$�6���%�v:s��l��R�����Rq�,�xá����B�g�Ǝx��Hs������F���l�uT��X-����N9 HF���r4�o�r��;뾺���\檚�Ϟ:nyݥ;կ[�*���������xo�k�{��p4l��+#��:�3S#E>G�q�͗����X�^���4'��!I�p`�q)1hHiIh���>X��L�K]>x��뭤��Ǔ��:�p���xi�g3��oռ(���:�f�E�w#IB8#�t,C�D�[��T��D�5�[)�Q1�Z�
�X�5"�W�&B�u�jIJ�K`�`���eB6���+#W\�KUUs���׶��n���zR���/�w���ǚ����ʺ���|=C�����ٷxXs`��(�[�P�Ē �w?Q�������á�l((�x٠ӼӐ�uZ���v�"Ha�CM�(�\�z���	$��CĠם-w�7��u��su��-J�o\ܷ�.�.]Mt�a�پU��	�c��D���YC�o�i�?3�?��Û�L�Y��x9���I�������J���B_ɯ=v��V��r��R��w�z4=�����p�{��,v����D}�b!��Z�)�mO]49g�>j��/#9�@�X����%�o<�Ӯ��ԝ:��sm����k�����0��h�l:��cN�N�Zl9��I\� �dtrMԕ4`>q�N|0XPQ�(��A����IA I��Dw���#`�n�
,#Y�b���{u�[�H*V�1�j�9���!�Ժ�OZ#��j㑤Fq�5�6�����"	H;e�,&(Ֆ��j�4%(��dt��Q���^����]�Lbb��?;O4�c5�}m�W,�]vFCa9|m��p�����\fp��^g���K7T�c�M¹%���6�g��Ó?�����D�N9�<x�� ��Ӂ�W�dg�<�����#UI��d=~q|�2=t���W���缮�[��k��L���4-`�4x������~�dU֛�^�sn[�"�zn1%��œ)��q�GCQ��{N�����=uN8q�t�눵���ZZ���˫q���:zu!B/!
P�(T�+Z�
�I8�=m֝�d�R:t�Ӯ:�:ˮ����8S8p�e�:u�T�Y�u�Su뮸�֎����N�o�Ɠ]���ŭUo�Y;�ߋ�����Os���s,�a���s�p\��������#cg�u6~�-N�7s�����KtVq��}�����)\�G&MfL�ow����US=�����wUT�gw{������{;����=UU=�����ֵ�.�wWwye�E<G�Z�6�Ą�>��pv6:l3C�b�9hv,�+�/�-q%+$I��!w8��7n\�G����m�_����[|<fK�aHF�PPQ�(ѣA����hw���gI��l��(�Z���?�m������s�tvI!���wr����X�I$�n�v�m�{�����Ӊxo�ɕs�B����׉#ڕ�0�(ǎ�0`�#�8|p9����$7�:����G���ȿ��r�����ywG���ckRM�%S�aԖ�e�K\z�ulN�V�0t^1H�&k�&D+a%TD���M6��*��3�F�C��tۆ�l���9�i�Y�:8k!!�0?���o#����$��JS�w��Ӧ�[�}����NqĄ��R	~4��S��y�K;�g��4��i�նm��L^tƞPպ�㗛�,x�<1���v�	$&�C�������ʩ.�,�#�i�1�4΃Bs����߼o������99˜�8�o_2��[>:0`�"������eP$የ�		�xp8`���UT%kM�i�08NG,*��僎Fr4pwk�ӵ��i�ɳ���
>v��O7��*(�Q�-�L��q�2��q��{F$|�FO�e+���ڢ���w���ی!^#!3���x�9����v�lr�=��4���7��޷ݝ� �*iy�sW�׎]�,((�t�d�yθ��)Rb�q'	�Ջd�أT�����8�����Ѿv4�#�H1�ft �o;�u΅C��EV�F�Q��X$]���R�I`�% �(��\�EN��U��2�2�@�:H�$J�Qf���3���\���C��
��=�:�C␎����1���eHT�h�	mYwE���$hq̌����L�~:�w(�D|3���r�թ��S/�B�_��g;�BI+r�9̡����2�C��m��#$m�2p;a���{�$m+\6�2`�&L\�]U�'I$m��|��$܈���0�I�1�TQM��[F���W'�[�Cc��Ɔ�p���BI ��v���e�R�7��"�?	�9m�i�˟����;2t��y���ؕ���(3���CH~��k8���b�L�׈8g1��> �I����Ys��0]�#P�*���c�2؞��x������HQ��� �������ou�m��G��`���RA��W�UJ��[m����7�[�[y�zV+�����uҵ��6��3mř�<7�����sN�:�vyD�Ro�ן}3vƛXh	��M��M��M��m�F�kn��b����n�M��h�X�hu��	b
�ebA#Z!4:�kM���&�	�hM
BRSL$�$�ZB��g!4(MhZ!���h[B�hZ��D&���g6BhP���&�B4,C�pΡ4(MЈMhX��:�9Сb��hMs����ѝ#8д&�B�&��hM	�k�!hMBhZBh�!�7�4,BКB4&��	�hMBhX�д-MB4�M4�MbkMi�L֚i�Mbi���M4֚4�i���M4�ZkZki�L�Mi�5��4i���X�i��M4�Zh�M5��4�Zf��M5��kM4֚�D�L��3�M54Ѧ�i�M4�&i���Mi�MM4i���7�7�֚4֚��M4�&��4��i���&�i��h�M3M5��5����Y4�M5��i�4�X�i�DD�4MmDh�MD�h������h�X���hDQh�(MY
(։!מ�"�BȴH�ZE���Z-&���M"D�4B&�"�5�4MM&�M#I��H�i	4�D$�i�I�$�4��BM$�bX���I���Y6M!&�HI����d�	4��M(jM!&�$ҊZ�SnM��"i$�i	id�M!&���%!6M&��HI�%��M6Y&�I����BM6Y&�I��4�I4�l��M&��I�"e�bI4��BM&I6M(����I��dDI��Ki$ӭ�q�h��F�I��I�w�i4��M!&��$�&�i4�BZY&�Kd��4��!�$�d�I�"d�Y,�&�HK$�M&KK%�d��6�&KHI&�&ɤ��	%��d���-��d��4�Y&�$����I�M��M�e�##4e��-�FXh�6L[m�M�mchu��ʹ�l�h�6��6�d��4�3M��M��M��c��1���M���k3M�m6��M��6��� ,�O����5�b��T�j�7���cddPQ0Qda �$yB�&���\��8kӏͯbp��WQ��g����p�s���
'�^:�8{Ñ�d�{V�Ǧ��5Y?��4�!����y��H}a�;g��M8p���7�r0��r�N'P��>~�����{�x��|�*f�<��?�[��g4�Y�����	�~9���@���?����%]��@��x�S��r����x�ϏF���} 
��Oq���H>򀉢cP(���	Y�<	!��`��m���D�S�NF`-j7�]xn���N#�>=q���4L�I�# ��O����6�G��C�f y���4@�D�0Q@�TP��B-f�ؠ"t��nk�O��2��uE����tg,�j�	�f�BѶ�P���l�	���M�I�@D��1o!6Ww��G��y;|*'κ��S����+�?^&x��$:�I��oS���h��
�<Ԇ ��Bz��K��^�o��?����sM�(w���G�>������h�b��H���!����ޏ��q��c�{� ��־x)����Y��}��o����CE���=q C,�} 
��ЬW�z�?�ޭ�z<0:�ŝC���.�1�~l �ȟ��]�IHN>�2I0�h�qED�@b`>N��&��%��&G*R�+U���D�TD�uxmOC�L�_nˠ�f��� �`�(��A4�t�����;x�C�U��	��g��=`<�A;���������?�s0?mKڰ��v��8���*�����ϐ����?����N#�T��ΥO�`����,�,յb����B�[+++(R�P�����������������(PV�Z���
ej��ի++eee
��eje��B����յe�
յ(P��B���5b�������+P��Z�V��B��5l�YZ��������B�
j�F�B�B�VP��B�6�P�B��ee
+
����6�YYZ�
mYB�P���)�
�mB�P��(P��B�ښ�P�ee
(Օ��(P���������el�������)�+QYYB�
���ի+(V���YYB��XS+5552��)�j�څmY[VV�+j�ڲ�������+j�ڲ�����+j�յemY[VR�Y[VVՕ�j�ڲ����++j�ڲ����jڲ��[P���+j�ښ�ڲ�����j�ڲ����VՕ�emYB�����+j�j++j�ڲ���ڲ����B����+j�յeeejյ5mB������������Y[V�VV���X���(VV�Պ�+(VV�+j�ڲ���5
5�e�mF������VյmYF����5jj5Q[SSSV+VV�SSV�Օ��j�ղ�ej�)�jejի+SSSVՕ�5ej��իV�Z�����ը��)�QYB��(������QB������Ք�(SQB���յjj
e5jՕ�SV+ej��)�j+ej��+jSVVVV��L�M[�B�
e5e
(Vڅeel�M�(SVP�X�B���
eb�ee
ejmB��M�V�jښ��P�L�B�H�H����	����~4�"u(�s9�+��:ϙ8>ӱx�����z��H��°��� ĎI$�&\�$WC�q}P}f�z7W�����1ܡ�	O��3�\7�p���2 ���{O2�^f�R�
���@z�U¹�Lp�n�����9��q�đ��P�Bs'�p�=��~�:ǾA��	� ����O#a�N�2��{�WW�mf�Nӽ�xh?���wgȇƖ�h0)Ϣo���H�

���