BZh91AY&SY=�d��X߀`qc���"� ����bD��          ���:Ҥ+lP(  � H � $   (R���� ���P@    �ˬ�-��(�hk@�
*L�%��4ZͰ+TX4ѩ�F�Tŀ
�me�"�2T��=� #���[\  Wf�ttkMP� ������s�*4  �Ka��	`mm P���k�+-l�(С� h�JD4  >zR�  rءJ�e4j��P�� �%6���P�a���m�T
�B*P�XM�m�d@hw��y�mZ�!Z���T� o��t��oy�{a��*ԥw���v]��T�Wqu{oV�]
�ܯx�=I�ާ����C�^���{�E����v�}�E} >��w�4ѡH�͵�ѐ �Ҕ�����>�N�q�zA�m=�ΩEKǯ}��}uh ۶�}��j������@���/�zQ�z���{���=}�tm'�x= el=��秠[+V�V�֖�Zѻ�J� [۾;;�IR6��ﾀ O}�7�[@
�^��Ҿ�V��O��YW��ޮ�(hƟw�N�F��}�A�mm��n(\�wj�s��B�@��  ����P�T�`��}F��g��Fj�m��J����vkB���'�:zr��U��u��t�::.��R��iGB�M���Q�Ҕ�k�x=�P��F��6����ScQ��*����AJ�m�W��
�Ps�L��ڻ�m玎��S���h� ۅu%�l��<�U����t���˥V�{�ATtoNҶF��M-��6X�c�UJ�����E7\wn�b���[;%���U�"�����A*�3�	���� 7D� wnt�W
�ѥ�Z6ŵ �Y���P8|�5r�uAA��p
�n4�ສ����\��5�\��s��4X��H�}�����ö4��'l��
Al���Ҫ�z�ѫb��T�K����B���q@릮�U������vK�����:5[���P�:�4�X�P�4�Eh�H��|�R� =��Ekk�3��h�2��]\ִnun� �i�{ҁ���۩T�]�u��8( ��Ƹ���π 

�*�B

* ��2�J       ���*16� #  L ��AJU#    jx@��%	��b IꔐeU dѠ 4  I5�$�*~#Q=�Q��4b4���?/����~����w?��4�RE��$��f5��|7������=�W��(�
���t� "�ܪ�*������J ��A?��<����x��B ��$�}hT U�*T Q|����~����1-�lK`��6Ķ%�0-�lKb[ؖ�Lm�LbF�Kb[ؖĶ�-�lKb[0�%1-�lK`���m�����m�l[b[�4�`�LK`�ض��alK`�-�lb�ض0-�[��-�[ �`��6���-�lK`[4Ķ1-�lKb[�6��:e�i�l`�ؖ��%�-���c�6Ħ%�-�lK`��%�-�lb[�6���#-�lb[ؖ��%�m�i-�lb[ؖĶ�m�lt��4Ķ%�-�lKb[�6Ķ1��-�lK`��%�-�l��Ķ%�-�l`��6�`[�`��6Ķ�-�0�%�4���-�lb[ؖ�aL��m�l`[�6Ķ6�0m�l`��6Ķ�-�b[�6Ķ%�-�l`�2ؖ���-�lK`�ض���&�����m�lc`���m�[؅�m��Ŷ6Ķ�-�lb[ؖ�0-�LKb[�Ķ�-�lb[M�-���-�lb[2ؖĶ%�-�lK`[ؖĶi��)�l`�ؖĶ%�-�l#b[�Ķ�-�lb[a�ƘF�-�lm�l`��Ķ��`Sؖ��%���-�lb[)�lbi�%��"6��(�b�l����F�(�[`�lTm�-�Vة��[`�lm����(6�F�	l#K`lm���Q�6���b�lm�`�l)�-�Q�*6�� � b�lDm����ب�b�l@m���T�(���*�`	�)li�-�Q�*����blAm���0Q� ��Fب�`#lm�-�-�`#lm����
6�F؂�`%�P�Am��Q� ��F�� [b�lآF(6��(�`�lDm����*��F��LU-�0A�
6�F� �b�lm�-�E��-��(��Fب�F؊�؊��`�[ب�[b�lm����F ��Fؠ� [b�lAm���E�"�Č@m�-�E� ��(��*6� �"�����[b�lQm���@-�l�U���F�"�[b [[b�+li���E�1� ��Lm�lQm�� #[`�[آ�[`�[ [` [��
����m�l�4�b[LKb�ضŶ-��6���-�m�lKb�Ŷ�b��!lB�4���%�m�lb[ؖ�LK`SؖĶ%�-�l`�mb[ؖĶ�-�lKb[��0-�LKb[ؖĶ%�-�l�`[�Ķ�-�lKb[��IlM1-�lK`[ض����F�-�lb[�Ķ�1�%�-�l[b��6ŶF1��-�lb��6����b��6Ķ%�-�lm�b��6Ķ�-�lK`����m�lKb[ضŶ�lb��6��-�m�l#ؖŶ�m�l`�Ħ�-�lK`��6���1-�lb[�6Ķ���?�5����@���]���MMT��yM3���X�#jf�^���Li1e�Y��n��UW&��p�[i���8BB���aSͷ�2��]Ʈ8)d�d�J����wEe��+`U�$�u��;�n��fe�	X]�C �f�FX�u�L�2�j�+��Eܐ�R% �׉'ۭ��X%f��eU'q��i4�0�t���-6���"C96��"Mk[���*^��y�ֲ��Un*u{7*�\����a�-�3i�Pc��YW�i&�9$"{nÂd�/a5���*nȲ᥉�.��T-�[Wj�� ����6�6j�R�,���T�Ӷƹ�3��̡3�����HMխ���tfZ��N��#*Q���
�NYL�j�۹�5�Mb���͜��a�2�UUR���V6�iXLͻ5R�k;��Q�m�/6T��5m,U��
i��7eJ��tf�i�N��p�jW;z���)�QP#l�7y�()�dw7+�D�{�0Hvfu��Sm�u.L��{M�m�[7!ڪ��\�3JA6`ՙ�{�6;/�(#�rL*�/�[��4��C;�Y%SV��2Q�������N�ͱn��r�<�]!e�7f��0�[2qқf!M�]���n�X���̽�]�saYY�k�ܥ������U�bU�Tɖ*�n��Q�J�7'	ʹd�f$ע�'cV�x	ĵl��A۬�j���r���t���n�'5(�Jq�a[����P��u�N0�=G"�ct�tU�JY;�Ô��{v�kV�)��x�#Lا�.��Vѻ�J�� �ݯ`)�AYǷ�*)��j���>�6�ӏ%��7g��nӠ��YFf�4��fdA7��i�9�U�$Yl6B���S�%=���4A�uJma���UIe�kj�U4�aV�1���2h��\;Rg��WV�S�":p^J�nRPC{U.{j�6�ܺ��EQ�֕G��7	eX��.l�d��L����`����sl2q���s7"�[C2G�6dT��j�HJ�Ԅ�f��B����3d�!fq�l՚W3��(�(0�'cj�UjS7j� R�YčÒ�6w̄�4ٚ�ク0�A�6�/4(X}�r���]Լˌ�JVv�O��`m�E,5S������RT!N�p�{�V�6d)��
{��׭�5���*�n�wr�
�V�����f�Яe���\.�+�I7�B��J�x�fe�	!����Ȳne��ҩ����ԕݬ.��Ԧ��n�T$�¹s��
�D�:�d*�n�-YyU0�f���ǥ�4��U���k;�"6\%��f�;�L��&��@�Iͻ�tn���2�浌�b�%Z�H������X��I���c;1�
֍�z�p��ڕYn��ʳh^<�t�Vb�-�C2n[Mђ��o�j�4�9$1#x���i�G�����I=�Ln/^�)ˡ�'�u��n�k�dB�9��/b{h��C
�Ņ\��n�GN�l�����[HƯ+7Y��A]�%1FҊɣ.����0]�Q�n�n@��N��-V9�֊2�9uw����e��^t�ҹ�Dkw0^�	LJ̔ ����Y����30f���ȫ^Jl-���E�yx��v��܉QZޡ��J��SE���URS{��jZ&T�j�F����e�d��gґU���9�v)��[�0ȱ�jĻ��e��ڑ���J_Dlm�6=�i�VjxS31��z�*�d�R6e�H�cSױn���A�*�6�+�����©��'k;B�RD��oH��b5�����wul�X�8@�j�5xVixs�D�
�+P�y��j�t��ӗBV��ú����d��56Fi��P[��qx���ks|���䤐˂��m�yIK�ܕ.-U��=8�I�'�J��IY*�mn8���2�Z�WE���4c!mr��qe8n�/*��e�/jC�Ty�W�v�ӹP��y7�&���)Nf�e�N�)�D��`��^ѓ�ou�;R�,zS�I�fKۼ�jAk�V�&�5+���e��F½N�62��ʕ�W=f�Mҋq��.M�iɑ)�i��J��a�"n��Y1�ͺ˷T�r�ԧy��BSw0���l�(�b0�0�CN���6��RFS�r��&\P�W��r�u�&r%)��=׬��r�ҝc7@�]��(�Qf�t��7r�fm�Yx��jŔ�9^5Y�t�av�i��'"+1�'3���J��������QǬ��.�	�;yV�m̱Uu�Q�*i8�1E��m��(D��QA����`�{Bl�
a^^�Ya֦�x���XQY
V�dJ�ǆ�i�Q�3C���5k��^�KY� þ�d�÷R�44�V�v%����CkVi�Vʘd�ө=�c*�S�"����)a���ǻ�g����i"�1�gEh�e���f(��w`�h��5hВ�U����(L��F���Vl�u��be-�Y�����[R�Q��U��7oJA#J�.#[i��d�7�(,m�2�K	f���L(�Y9&^\���v�	���'��nֱ�y�5��e�I�F^��jdah�Nhj��D����%]���5orA�]��t)fˣ�*EXso3)֤���6�^C�y�m�.[��{l]7HҨ�Vʤ��y5˖`�Y	u��wsC�kW^���2�(��*.fjlۄ]Z�(4�[��dPS6�Vڪ��=�+#�Z6�]3�u�;�vc����!��2��y�*�5I*9�U�n+�wX�E�$(�C#톳U�L42��)L��Q�U^b��`/LNY8F(8(�V���r
O(ڬٮ��͢4�}��."���T��ԙX1d��j˴5�l�J�#����E?]��]]սd`�*���ҩ�*��V���碸�I�K�AӅ`��A����&	��F ¬f;ђ�\�V��A�[q���Y�(��鲭�����J8�na�ދw0b8,��%ħx�\y�n�X��h��1
�Kh�hֻ��=�li��F�������)�7]��Xmd��oj��`�&�-*�ŬG�����DF��R��	��n��M`�ڬ�mG�P�:�-���2cU���w���hw*�&�;��sw���jm�	6�B7��Y֦!�LLSn��by�zMfȨNCKM0w��M�ܤ%` �(��8U��ˉ6-�٪Z`�{2�����EՂ�+�36�ͫ��"T�L-D���B��%�l͈1 �tf'��$���Ian��]By����wlC�)_�S� �~��u���:�9U�R�:����yV�l���Ŋ��8�M��{/i�j8`U$�D9�7H��ė(�`�*O�r����t���f�V�J�0��^�!��K[/1�]0�2���)�V����T_vE���֜���T0伥^�����7���Y9�w��kI�Ժ�%�2��[�vL�a[���	�J�%y�LͧJ���i�d�����;�Fh��ȶ��i���+CwB��JJ�T[.��e��f�P�M!�9���1�4�@�AK��ju�+7���S�Z�h�����.].�HLwUy�do+dRm���Q��n�K"fm�ʍ-���+&�*����^lp��
��THg��K	��a4E v9{{���Q�j�(m�x4ӎ-��%!�JܬB��Yq�[��Ҙ�a&UH�Xr�FK)v�l�Ӷ0Z�O�z5�7��杽�J�����[V��V�-���⤌������QV�n�&B��V�K���`�v���4�K`�R�8�"S�ٰ�T�ۣ�r�5DY�oL��\v'D0���y�KU�"�OpԪw9��7Y��j��C���q��ۺ�l�Р���Y�P���˪��Zp]@�3e�%U���z�c*�X�k����*�5�t�J�o.���d�b����zQ�5d����̱k�۽�Y8��ލQX^ح
�7/%a���
��ǘ����I���c�\�%�8�k�:�V�q
�P&�����IŉE���tp��2�ۃ���«-#�қX�/kS�H��[D�omm�j!��:�.���aS.��59�JNr���ƫF�0Ż��PUX�Z�7h-&�
z\RǗ-){5�mm�mai�1p�+���,Ym8�M܈��+�.��U4�Th����9U�h�T�.G3p�r��V�F��~.���E��JA��%�Fn�F</���\�7z�kJ՜�T�/0!���K/T7uz��E��{B�L�.��6`�G�����L��w�[&�www&Vx�X��F�l�Į:����d�u�w1�Z�̫��I�R�(֩UV؈��U��iI�
��Y ��U�,V��M�3�Ǻj����lD1�X���˺yk!�8���RJ�4�BY�J���ex�T�f	im��[�OY�WV�n�X���5���tR{-�y[�&#�&I�5)���u;�s%+�UtiЛ�y�� �Ի8�]��[��n�i��'�L;��ӑA�Jӓ-�[������Xr�}����T�œpnneJ/M�Uj��J7�*�K+)�"�Ns�e�
�H�,������&2o-�6�Ռ׋u�ڂ�^�q����/)��`�Y��sr�=��,�c���t)�uTwI�Ց[$8%Y�j�@�;�Ȫ�g��n��4RSIM��]��N��wKD�V�˓nXEJ�3�z�����ů}���Pl�m���ɴp����'r��0��-�3t�ݫ�J���4�B9#>o.�����Uf^fZ��4/qn�P5��K]Ga�+j'WN� ���[Wzr����.��vA7��` �w���u�I������˩�ҷ�i-�*��AvwU�,eژ%j����kv�3�t!Q�z��6tB	�r ����S3`�s)fF�G��2�9l�6�k`�]��YUuxB��&m���ֵ!�G��-�"�e�J\Y{0��^Uo�9k�ڈSfh�n{1�3�Dl.\;HQ�32�O&���2F$��x	�q����l�X�BB��5cw�D�wc+X�,�q孼)^�.l�7�bږ.�rE���l�:�'R�3qbŗ"W�"
F�dKw�c0������buA��n#Yw�t�1fZ���P*��eQ�P�~5+v*	��+`Gճhڬʶ�̈́.ʢ����Sʥ7fN^88!��,JØC.��R���&
�`;vM�{$�r�ɛ�V��Ube���F��F��yt.�0�%��X`����8g#1V�r���%svPE���ЉrU�7uN�ч6���X�%���WH�w�j�2�BD(���A��V�KS7H�.�{K.�e�[��Smm�zvi�y�^*9�̗ya*��)&QH[RnAe3QnC�)+	��h��a�2��0ܶ��D���2�SUU�&){$i/QE���X��-b���Iؼ�o%[S/�f�����`F�8���s�X���e$LL`�ef�m�M�	)b�D��t��pG����3�@PӉ��!�wn9Y[��̩i��Kt���8�u��Qf�WU��aΈٳPHݯ%���-S�-Uq��Bvmēdd�fj׎���$fwNAGEV��R��G+%V�PL����ˊ�J����Z/&��'�k1����6����̵̖7�$���	Wa
�0��N�QВ������5Ƃ�1�LY9E96�,X4�kQ�P`O^��פ�W&��v�kbI+hd�ک%Q)Ǧ��G,n-
��iЈiɆ��/6�:�Tz��\���x�w#I5�j�'w,�܃]a��V�J*�R��k����J�Xa�js��eՙ�S:+QƝ��L�f���0�ٗ��u6U�˶
��
=��㷻��b5�0�&�N5!فTXt��6+2}i���B�r�b����˅���o2�-�b2��S%��{A&[,7���Ҏ�7[ ��M�9cRܲvlj�F��f�^UbS{+/M�%4�u�*�v��;�{��e�Ś��KR�]i%v�4-(�j�������ڔ���ҀШ��#}�mKZ
��,J��F,J$�dwu���C��گi0M���]#IEI0i�yN6�FӤ�X1�J�Ȳ���47/8�{X�-v�%j�mNR"�,�Ţ�Z]��X�T��QdO3��%K	�O������Z�i7�|~�[�K����u_Ցn��Nv-�*P)$�j�dGU'j8���,T���I��jM$�)L�Z��
=i��*J��Q-T���J���{���k�ڽ--\��M$M<�4�'*򮥹��DƖq�.ҋRx�8e��F*�ydWj�gJũ4� �m��&�ւ��*�A�`���@�k5Y���Vm^Ե1`�V�v�K�j�E)��Km�L��X�ؕ�����ҵi*L���n�:��TW�ﻶ]]�L�Q�j��U�\�ե�j���U�bI���- ��R��V���e���t��	���Q�:�����W��_,I4Aض:��W��u>CzȗS�v��Tx���T�ux�U��:j;$��m~ե-HJRdn'>E�L��Z�~J�iR=���f+HK�;j��ަ;���w%��w���eN���*z޾��m��n�eRR�a �"���Ʈ�S+��j�����,Z������k5-2��N����lR)��`�'�RZ,�S1RUVe�=����r��T'uZH.�Im[��V�H,�u�E�C�}g��Z(l�_R6V��.�&,h��z�A�҈'���w+���]���8�Kz)nC-m�;�E�dR ����Y�C�p\�~J#�䦠Τ��J^R�jr��IH���Ղ��XD�K%��D�QN%D�[T�.��yu)�b�R ��	�Ï-^.���\��Zr��j��Ԥ�^���\�E��)��)4��V��"ċT�౧+�J�j�Ȩ�N�㻫ճxK�@�}R���V��P�iR�W���Fu'�rMv)K.�@cV��-^�e@TZ��Aت*�"-e���o,�9w+��ؔe������g>��~P?��zT/_���<'���Ͽ g��l�i�HL���\�H�Z�e�6u'�	��,����Rֽ9 ��Ր��c0k�pb�{��xJ�*��Y���}P%׹��{�P$2%�k[�w�P+%�iS�"2��l�D�"v��/Z�`�)[,;ۆ�l�4��i�:���D��D�h�t"km�H�h्nL��m'���s�=��y��x�nλ��Ni�����'k�X�ǖ\]L���9�NŴ�Г���/�&ቛ�p���o�+�}Vt\�`���:�Z�5YR���f*�+p�j���\�:��:oq�Q0��2il���R$v���*�i73)̦���ˁT�k�O�E&�N��%�RA���/L�٥nW�Iw[���͝���z��R.�ݛ�f�P����ٗ/_3Ɔ�M�ɔr�w�b�R�ǅҖ�gvk
wr�%��ikO.Q�8o9bH-������(�\�od�GȰ�F�(D�S�9�f��e�c&��ݓ�.űB8�MR�k�I����).�S���͝á�{����7�9���T�5�V�="m�f�WA�7��ȭ�8��aux0�%MA�SV��瑤2%N����G��W�fl��ޱtaڪ����t{oL��/������T8=z��1��2���0`�NMk�4v��<��d�uor���7۽e���l���;R��r��7*�Ȓ��꭛��5ven<A��3�IJ�D+R�,YM�B����&]�r���iM�����kO/iQ�Yjj���т��=Os_0WG]Bq�s��N���ț�X2�T3RPI*K5+���m���8Em�*ܪ���n����K��L��2������E� �M�)�.�^^ڬ>�q1Y�w{�N��إV�i��c#��Yk�-����thЮ��vE�Z�^���Uh/)r�޵4/=�i�4���}6-myܮ�d�z!��/;tV��r��ˆR필��u�j#��<��_Fۋ$�K6�iR7�l�9�v��۾�Q�u��C]r�KiC�{�n��V^[	lά׻�:�r���n�{dH*�a#��kX2��݈�ՉsB��n�iT��3���nE�9{b�4ҧ�u>F�s�9m+Օ
y��uxdx�sG��i���mb�k�rV��R�P��.c.l�q��7��8̵�pn<Ye��n�=��O�j��Ώ^�FcH�V����n�d$��Ω$J,y�x�!���V��C֘�T6�t�ǳ&iAsŝ���w��M�'�Hk2�;wx�Y��	9&p���6��Et��]�H>9��e�AY[�7���GʟM�[z�]^7criHe�ۄ���
\��_fu��.=n̢�rx��bm��\<�N�M&�V3Mj�Z&�H��b�o=�ɹ|(�;eN�}�D­���+;��̈́!G,�N�FjX�,��DԍSX��b�^���OI͹��u�H��$�Jzlѧ;76+ �W5q���Zܒ��e���Ji̭�bFi���1�C�Et�}�7\�:��Keؾ=�t�e��˟Wh��F$��^Ţ���0Ѝ�F���.$otW-����e������wu����୚�&�"��%P�{�K�^�=�T��_N�T�͜�囆�5����Q�j�gCy�D��	���
J��5.�7X���n��b˃:��K����G�ƠAy�&��ބ��4=&�!�҂��PZi֜Ү�\T��fY���z�Yr�(���<*�4�
���`��++قUoj�)Vj��vl���	�k2=�^��C�1`��t�Ie��dfe���j�`��qb��v�e"1*��͌v�ï�*�2�)4��1�`�(=�۬�;�w�����a��UFcCl;�]ז�f�C: �ɒ6kp�E�����^�"(�)�;Rʝ�-z���)�ҶF̺�Anٰ�3&a}�B��,�|$��P&���uI��T��e��K�x�	��5oL�׬MZ�X�1�|�\�=.�,b�q"��Ͱ��-u��!�el5�$�K�d�UMؓ�{x�:��U���گ�F�:ò��[EҮ�W˕�U]�ut�I�/T��[��4��x�~�H��UK\5�˧�[X.5L
f�5�*��m�9N����;:*��rk���b�B�5��!)�0VB�I��6�9w�D�\�&�b�oE&hOL�UMd�G���δ2�ێ�a�Y`�a̩	�e�vH��+��\T��.��:�_���/wjss����Yx%����Y�'i�j��L��W�˃���Ia�V��'���uʍ;���g^��q[Е�Vt��:E���'L(M*�v�{T8ݚy� ��A�Wou�g-Yz�6�����1��QZ!��C+d��[[��UJ����S�b���hSȓz�$�J(ȶ��-��`�U�2_
v�tgA�j��u���`3K�a��u��f45�<}�Iܕt��RӼ�Ǯ�ƷT�)�D�l���0���U���u&;*��dl*�J�\�٘Q�G.�ʌy�$��i7����u)�ʏ9nѱoni5z"��c.cK�#63U&^Lc���j���V��!��k�8��)]�8�in8��ͥ������c��UTQ���nnE*,�x�[��w��	<�
n��������{[�ՃO�K|�a*����̝�uf�t��	�j������"���pf:#
ׄ�1�zeR�'H�J��'lB�U�4��jëxQ"ޫ26wo��8�Bf��bQ�6�퍲�KhLɬ��6�C\X���O���R�T��|���+S�f]ޥV��Y;2&�ɩ6�q�nZM��ju3���7�@W�oiK��S8��Ǣ�"��ԍ(�+h��7-b��k����b�Z����oK�fm++2��/h����Va����ss�C�4n�B�+*`�kjR��ټ��h�-=N�aʆ�*��S6�JR��E�h���*l]���fiۻ�̣��p�peZ�7X�z�B���ͥm�7�2���J^eacQ͓Rn���cf�p�=m�;�Ĺe�q��O���uΫ�*$#5Ċ񖥸�UC���Z��=R��nV�%׳�NI��t�PYsZ�V��j�m�:X�U0ْ]��2�UT�4�_JHA&dd�9mE�|��*�b�X���j27w�����-�Q$�J�[��5>�V����`K���-�x��v�7n�\:�%[DK��5N�fq�Z6�(�*\;�����%3 ጉWS��5�<b�L���Y�sL4M����@�1����s!�<>hM�Fc9Ib�������-�9u���X�2�}�����.�	�6g-+��W"g��u��3��T����u���n��j5j�j��ν&�[Pٚ�-��RXw�Wp7����6rh�2��5���(l��x1�3O]�[�؆�����ܬ&�v���*vu���^}�|�<��3$]�z�;47<SAj�f��U\�ފ0ۉg�NU�]�[�+�����bɳj�(�:����J��+V�ţ��H���oITz#]�7yx�YY�o�dfXq��Y�5���ԳRL�9a=��Nk�.U�Vn��z�X�΍��C�pm^+�4�A���)U� ް�g%⑚�h�a@r� ���Sֲ��U���m�)c���]�R�E*���x�{'iĵ3�T�ȃdԖ�V���0ͼޒ��i������>�w��V��nQ}�qAdG���v�J�]��f��n�`������5l� �D�Fl�Rt���X���DR�XEFw�����T�Vb��L�%^XP�=�a�xŮ�!<����b�����W;�b��HҊAR��~2���5�!��ᲯM���>x7YR\���]N͝Ï!:��Z���qIS�z���G�Q��yvS�X*��Q��4+46��͸���.�`�Z^�=%Z����������]�'=8��W�H�� �An�fURi�u9�Ļ:_-{�<�w���b�2�6u��Q3�8�gu=5�vN���!����DV�gM��6�d=�a3yfN�U���l�xv�;{1*
������!�C,�����@Y��-�q�^�b�eV5d*��	�b�.�e�j��gJ�K���X٤�Ƕ�aއsVh�]&�UH�׃g�`�h�Vf��@�ȕU�vT�Q��Wg&B�����\�޶�j�c+�uwP�3�.�ka�7�Q���z�Rb�0����'aV)z�[�OZ�WJ�j�=�:VT��Mr��IvM�����@����Q;ws�-�C Da������mT�
޳]��ag�Cb!<���$ݠ��7�\���ܺ'�����T�������;A�N�X6nUjʖ����F8D�-�fm����]�,��gf�eQ���f�-fgO#���V̴]�U��;1���ؚ��kCY{O,�^��,�:ۣbŴ"֠U�����I���Z3{Q��Wڮ�a�˫�������YΟ���U���.�R��	�v9�'fʊ��y�������5>ͭf��\�wѼ�]%�?��NhQj��;{�{Ƴ�ff��a�k��Y�Cg4^�0�S���U�fZ�@�E�h,�r�8�XA_[ɻw���.q]=}b��']Ն���[E���Lj9*f��æū�e%h�r�B�5���h�K3"\�MS��Uٽ�ٺv�9��U�בG1w���^_hX��O�t��s��;���oX�g�!��o���)��ɤ)r������׸RG"`�WX��
ex�\�ؼ
�Ӿ/�o	V�L؃�m<R����Ĭ�5Lemb���lS8��GX�6pZGCM��D�o7T����@ﶊ��z`g/����Z)��T�Ո�iVT7�0n_WR�jk�_@�X�eN��X�7M��v���r�_b31uj�m�ΥU��l�0Z��}h��|��$�_*�U��蛩[	��$�q�ɓ��ʍׅ'jC���]���K	$��4�����fCP�uӲo��n�k-��P֮V���]�Q�t��hN���9FT�VX�9�F�(�F�����o)m�]��2Xک)c���]�H��^��n��'v��3q��^'[�wN�����:�iޞ@�u#�V�f�eL�^�x�eW;�s�ӽד�;���m&���7S�����'R^�sx�m��C+M�T�wȡm�M\�8&�$�� ��u#.eL3�-�:2aa��Ղ��$s:��䈹gI�z��&]كI����α�RV��v�ګ���V��b�+dfm�̼d�xF-I���gnZ9�n�Bn��9�Y�9Z^ښ��L�(n=����#u5����h���dHG|�s�	[b�`�.��!��ﯟ��-�\�b�e��s/�ݶ��J�5��;g��U�*�-}p�h9S�
��#��ND@�Rq�׎�O�Ws��1R mǓ��"�x���tJ�e�Ö�SC4:���n�rbו������U�u��v�a�o�Jt�F��!��V�#[T�v����T
��I5��gX���=H�J�]�=���C�ּ��Z�Gg/q'¶��%����8�->y���6%6�;e�9��k�IF�f������%k��K�D
4cr�eUoL�eZ��7�O%�'���(�2�6*P�ݦV�K�L����xĕ��^ơ��p&v{�o�磺KG���˺��u{����guI��d�S���fT肳]K.���n�R����R�o �2����OCS7�ۻ�Z/V��b�5�j˸�VT�a�ٸ�\��E��ų�K���磕�k��X�>*�/��+(AI�w�-+0�.�/Ef�!�9��rӡ[IHՏD�d4�"$�Py3aJ�Qj�����:Z娳����j2��f�]�Ǳ�evh��jlC+�ru
�#D��e%�sBY3�*X�s8�JY����z)���5R��Gk�3&��1UZӕHٝ��7,9p�5Y�i��t�T~��4�9�ױn�dvB���^���[E���E7�J�7/kh&����T��T��N�V��o�=�uK��!��5��C̬��/HiH<V������P#����@nG��'S���E�ϲ����R@{�A y�U|;u�ZG�#��G��]��$ � h�N�I�n��E�v�8� �.���
"����#Z��;SQʁ�N"E]�@��#rSb!.�H#�ՄκX��a��A$՘��>�z���;��D��-?�F��?cm0q]6���Xc�U��GĀL��m��(��Q�hB�UK�d��/nP8��xR�K]� |Ydm�{��h����ȳFϽdʴ�I��~g�c�H�%��%�堒>�̞�n��b���Ϥe��<�@���}���a�t�U�?u�]/xuQE���f"�y�r�����#�>Wz����=y��S
��8�!
�e&Ԓk�2�/ 5#��Z�)���wUz�'����H�&�Pa�$�KVI��{l�#H��7�r�D� 5
�!z��e݆���I��� A����DQC�ϴ'������4dPPG�����o�������	r�x�z��^�楧����Ë(��=��J���v;��oTU\�9v,SZGN����G��j�Q�ɕOr�XR�|f��m���)m��0�Xy0� ]^�x���&ݚMܾ�aǜ���R��^%O���*��22cƣK���ר��嫍��e���b���K�Bw�c۾�p��c��$�ЭB�z�G������*m�v^>�J��Mv۷x"��6-9P��Ɋp��Z�O��H�Tf�*i=�!{Ӎ	�nB���!��f�C;*�k�צb�O�&
ՙQ(*еC�n�K�ú�Z����������aul��4ٌ-}���팚,���լ��5���;f32&�c�᢮SAF��gkE-����UF�@�mꡞxiZ�F(��i�<�a��3�|pv$*CZ�k�)�F�����Ў�UwMDn�ò����֮�[2^A3U�r�Y���Ԫ4h��j�����BAՋ��\Ȕ;ۂ������J!uLw{4����'��&���|*bA�Urn�M�c��z�tjy�TP״e�m�U��T������*�=Y6�[:d�$ƈ�P��Lن�[2��ksB�q�����2�S[A&6�+w�R�6���o�q��8�>�㎜q�8�8��8ӎ8�8���88�<pq�q�q�q�q�q�q�q�_____]>��8��8��q�\qƜq�q�n8�q�qӎ8�q��}q�8�8ێ8㏎8�6�8��8ӎ8�8����<�[c��\N7�ӏC,�`�
|�ǁ_n;�\�Y6^�=��Y���J���R�f�h�u�gU�r�:�1y#@�`��.E���uW;�hd̪l��s(N��/Muf��
�-˰lk4���%*ۧ��{�Qg��8���;U�Q�tz��S�F��$K	�����eW^�V`�r-��t{'e�uS
�.ʆ�K('QjJ�X�>�ww���Qd'*ZV�]7B�]Z��)�E�i��/\5���A�:�M-�.��6�f�]���a��e��n3����f�Q��d�;��gJB�H�r���J�gJ��T��+RK�x�b��-v$��C��������.0���"�N�LΣ5�	4:�����©��ӕpnr���}uvn+�����䭨;ݜ��a�/b��.��tlV�N�ֆ��k�,�����*���\7�J}1�rS޾���2�f��|�$6���s�p�fX�}��C���i���:��LRh�:V�lh٩�gt�h��p��Sr��X��8ҽ�`�.��Ņ�y��a�Xh�fn�,)'bv&��Z;������`��dr.�y[�ѴQt�Md� a$�ʜ8gN��aF�;�b�k,��x��O�fjJS��� a��{��i��6��88�8�;qƜq�q��qӎ8�>8�6�8��q�\qƜq�q�n8�q�qǎ<c�8�8�������㏮8�q�|q�m�q��q�|q�t�8㏮8�8��q�q�q��t�8�>��㍶�8ێ8㏎{���^>WIXS��&S�4K������^�׮�7��)��G9����ʸ�/US����i�%�=K�p�h�Tڌb�ro�����`�ķ�c6:Z�a�>͕6\���GFD�%y��K��<�l��w
f񳒌ɝ��<�����֫�2�u4���pR�P@�3q�8.&p�U���V�F�[:�����M��R��]o��'j�A��LF<��[v`&$,��C^RnL��PI^K�e�)�Y����Mi����0mX��yx�e��B݊�2�кùZxj��+��T���Hhٻ��kg�Mk�xK�EҬV�Z�Q]��e�e�f�����3�Mn]H�Ŋ�39m�
N/#U��81*U��PĥfH��m*��d��rk/���c)����M�H��mI`��7Q�z�˩��*��N�d�
���4���Z�`��B� ��*#[37'��E[�C��K��l�P�i�b]>��:�,j�Ժ�{"Fo/B��.�WY[ʬ�c��X���즫e�v�"h��ٓ+j������;�N�����`���6�Y���5uz�ҒrEVpekk��]�=�i[�Q����ޝ�	Mp# �v�O<}=��g�����{q�q�qۃ�8�8�c�8�8�i�q�q�q�q�q�q�8�8��8�q�n�o����8�c�8�8�i�q�qێ4�8㏎8㍸�8�8��q�q�q��q�qێ4�8㏎8㍸���U_9~猗［�� W�ۛ�c1����n&U�����(X!m��iC�r�Ơ��F�k�p��f��c����7�s)@Ǘ���(���QN�J�z���x6�R��k�3���C��n��w�)�Hs_Qr�.�`=ptz�Z�9^�P�D%��� �8��X[�]\��;ni��N�������$�4��8�X�����g�֡]P�{��P�{7Z���B�b�V]oj��kM�j��N���S��רղL�|I�r��Iu����+t���A��7j��C��HP���v�]��m٫��N<�{�Ɂ��� ��Ԡf�F�L�%/h�b8�e��V�FB�
.-i�q�SoB�6���J� Vj�l��I����T^tv]cV���9ʎ.c��ý�A\��ۼw��ʛx��]����ڷ�ņ%_s�w��쥞2��W��5��B6�u�٧#�W���c�l��'Jn�j���Wdr�I��FRJ��fERǧ^�i���b���I��,q0S��Ͱ�1Ie�?V<�֍LJě��;wͼ�~vO�K�{uY�ğ�8x���ś,�Nڶ�cWH{�l�\�іqKjt#�[� i}דVsܲs�ԦܦF.2v��A�T�﮺���FtD$���T���4�D�wۅ��}��_�����}�8�n8�>8�q�n8ӎ<pq�q�q�q�q�n8ӎ8�>8�6�8㏎8㍸�8㏮;v�ݻ}q�x�q�q�x��8�8���8�>�㎜q�m�q��c�8�8��c�8�8��q����������P�3/)F��geR>r�B�~kv�ݝ/c.m��9^&ِ�s%cJ���*	��e�p\���(l=�:�^��9�Z�eL<v!Ĥ��𪜘�Z�4l���va��%����H���NBS(�rZ� S��|�v�b�R_1���a�6�U�e���-�z��� `��ؚ�Fv!�2f�WIUӇ�ǐR�o�Z+rX�^�����jab��f*��Q@��;Z��Q&�29�93Z����Ix�2��2��[�"�٥�Ê�WW�Ve�Ҭ^�QZ1C�S�m�mll7��XP0�I0DA�&��
���@�<5��#[EmẨ�7fa�{N�](7a���S%��5ۀ�wa[�
�	�O�c��v�E巩uG�j�Î��ݘ�5Mu��:�c4#k8a���;�9��ɚ+sE�7: �2�cpթ�@�`��8p�wϫ���%�X�pTx�om��
�{���LJ'`�ɹ����n\
��< �j�Z%�<�������C��k"�̳O�ەW���
�[(� 8�{r�Zك�f����w"��Jz�e��B��)e[�J�p3��#�ה P�f�/C�SU�؝ܲg���T��}o��.�VX)
ز�+y����=�r���YܶݬM�M�dS�MS	��WӴ�;�c���|���Y2K���bg��}R�+�J���86-h]m:�@zCڭ����h�@��uCY/��ݝ���қM�y6������7�� *�$��AK�����T���P脖X-�]Wdn���v�s�K&���w
,��=�Ch��:S��{b��V�z48�|Q�`�w��S�:� T�'���8�>��TgU���F����Fqq�}�����]�T��i�����]��(�a��+) r�mV<k��2��
s�� CR�%��W��Rn7JMZ;��(��v)����v%��&��勹��7'1� �`'�e��9t�N&�E1��Ӟ���Ӭ[����V��^<UYy2ee�3ԫM�	v�A��:�KtÔH&�c��4�U��M�Y�i�q��: S�fو�྾!f��{9��=��b⮱�,@��Y(��^�8��g�a'�Z[FTlj��P���걲B������qv�����B2���@��н����+4g���^n<�v��ۂ[wf�*�:VSid�Ȩ�[ml�mE� ���d{�]5'�pWZsm�1���S.���'�e#�	���*��Jl��cÔ��v�|"�f\�v�kJ%'U�#B������76�(j���W{�^�ۧT`Q�es��LA�6�8N=��hV�h`K�U�|�Wf���DC�W���o�eN��Pg����v��N{�m*�u��"K�+7 n��O�.i��v
��2��P(��ӷZ`��sE[{ǒ������21��4�R��)mTӽ�@Jl&��l����Za��+˃��iv��bY�l���	ޚ����49��W�]��e�ɔ���:�:@�W$ގ��ޕF(���f�V:�ٍY%U��P0ۺ}�dS��3b��5Yc�]�on�n*�N���K��Mi�����d+.�*�\f����y��̣k��0މ��_���bB������pf�l�\�����h̫��X)xZV �[�C�:EP7�q��R�[�al �w!� r�Iɤ�Zn�M��Iɘx1R�"��
�X�;N �{��/w*�&,=/+�29V�����;Z��N^�OR��.��Q�
X����_:�`��(�z��UC�W/>uJT}wa1\:�T�i;�<%���D1�t\ڮa�Hڵ��o[&��r�y齍3y�nʗ��KR�F�겘B�(KGmea� m+Fv��H�͍o�se�.�:��x�����#��&�ݞ>y��<,;�Hb3eX�F9J'�6�-�sl����l��M��.�L���],-�`�\��L8K���X�d�i"R0Y���o^��*76�A̓��Ѯ�Og���L�[׬է:J[�!���݉��UJ�F�⍃�a:������%���8��[U�)�m耳pFe�J����9�a�@z�]�ZM����r�t�%JNpK۪FI9[!ݼup6��oݍo���h�#ç89������WZPg4�^E�����Sx��4���NMۡ�+��:<ڄ�:m�['��R9�]�k"5$SR������Wsu�֓��ͽ��Tw���eu�q8�q��zn�pT7+��&�5�)���,���w�kɒ�2�9l�nê�mmDO�n�oK��]`5����]!��3F�,JG�TT�Ju;h�����m�7�8C"��L`m�H�[2���uǝ�]cy��Ź3&%�.ѕ[Xe5N�>B�n��v[��7j��=6l���usq�inmGBa�mK�h��[%�V`D�k��(�2^�Or!^��"eXp��KQ贪W-䦢yI�Z�Ҭ]��jí[,-B�)JT��U�v��L2SśB8�J˝A�A�٬ήE�ԃj���MV`����)�t"B6��yZ��)��ƪ't���^�m��Y�NuC�L�g34���+�������]a^4w����P͠˗H��"�b,��l�7n��ugee�=�xrJ����v�v�W�,���G;r��`��52'ݝHW
����LoIc�SU�嫁Ko��Uvkt�.���"�;��Gk�P�ُQV�"���R9��])�&ЇKZ���7P��S��"�)��Yn�Tњzۋl�l�ۄ;���ޡ2V�sEv*�q�Cc�nP�9�w��.Ab�X�D%A��[�K*�Ǐ�hf�ȵ��I�;�v�D����y�Sr��gV�����v�}�\�xjՊcq�mY��Z�.l�*vs31kmT��;��p�[�۫]����e9	R��V�7��ʨ�Ն�2�,����AD��3�+��l��c���;';95�9˻Y�,��n� �[�e��Y|�f�;e��+ƼA�sv���GlJ�#�7Fn6EK��-�.�������f��$�\�����f�����Suu�r�5۽e���Z�[��뎭;���@�}/�Cu6)w��%U������c�ɡ�LVr�O�Š2
�p���٬�T��;��^V���5������mBa�I�
ǎ�8�i��svVE��mA�,V٬'nq��bܪ�6�hz�l�;#$@9c+e���0�m��V�SZr�]�#��n}Jo0�묋���t�)9rk7�(�(;iU��sU'v�������ە%�*2piM���KV��Zr���svi7�+Rh����j���R%%č�'%/:`���u[�sz�!�fj!jG�QU��!c̴�k>���l��/r�������؅Y{M��y!'�~�Al3�tΘwE:��:�U,֍�ӊ��U�KO�z�_k���0AJ�:(�{��B�aw;�[�M��/{=�5�\�,��a7z�э�9�n�PF�ݵ'�ܕ�j����Z���7�^�k�Y��Aa|��[Ã*���9r����~4%k�&�5o��ͳ7�@�#{�k�R�;jNT�z�BWj�U�L����h�%���X�i�}6��絇y��j�b{wu|�M����@��,4����tn��^����+��sn��f�8i׋�j�dQհ��e#������ж�4�]'�i�v]t�H�<�}\r�PTE[N�sܾy'n�+��J���¡oV���Qi��H�oZ���м��Y�f��P �m�ѓ�XF�I�ST��r"���D+츙j�:��:�b�ѩη����K���x6:�s*�e�q�G'�aٲ�����^f.ܫ��N1��elyݓB�˶��14��NI�ӭeͳ�"��=����h��������@_������?��~�ܿx�W��'�W�F��_�FB�i�\0HP!&��H�����)Q(0�j)	6Y�I/OO�R7l5V�J���'!�|[L�a�^Bx���p�Č( ��Y�b���ayҪ���U#�4�@�6L.�
�*���T�GKTBદ�R`-"�	H�) 3�2IL�	N$D�:�MQ�J����RBKW��dg㈩U�K�f#�[GY��U��%Ff�\D�wU���5,��1d�776jC�Ǻ^`g�������#+.��Yl���{{�^i�#��B��n�e��̽�E��lQ+Q2Х'# �v���7������+�H;�%�lu^T�pl�K�a������gR8���	�f����8�Yٺ����[��UHƕ�t�i`͍b�R��1�Y�p�t�+���2Tю]\u;[��'��
ڠ�4�KwbM�OfU��$Q�N�s�TkF�����ᝁcy�Ṩ��nɵ��v)Q�>γmfj �k;�yJb��XD���q#T�(���E�Jz-����(i�`�����qm���e�7̵d]:�)�cӖe�/4ũM��%�\���Hb���Ҷ& �n�K�+	�8s��P��1[O\5c�j���y�m[�+��N�yY�Z��9�n�`���):޽
�?9ut���*�Z��U��R��fjf����[�4!�n��X��Gt����{F>��iR��2�^���T2��zkJdPX�j��ͥ�d��컽H���G5UL�iW`��c+��w�Nׯ����ਉxł���x�C�����-��'��0�`$"$!���'��gL�Q
��-���H#���n8ӈ�cFl�p��"2�p�F[Z[�/��RaH�"&�Q&d �����T�1"�1"bCA�")�ș2�P�d2P���-OF�)�(�f�D�6�aHU2E1$(��G��,@�D�6.�e���A���2a1	^P�ɒy1l�i�6����#I�"�A�X���E��M�P!@b�$$��%(�G)Jڦ)�K�(I0�A�bh7`�!�H����!4���`5!JB�R"dH�"p�G��ʌF�M'�H�i�`-��i�d�A���򈒂0��H$�a2�!4b-2��Co����y�q�t��܏4�$�㳜����e"1�R2i����\v�۷n�\q�a4"I~81��	1'�t����F4AZB��8ێ8�۷nݻv��;��Й)9sRE�M�\��`�����:z����nݻv�۷�� b�o��n^9��;d&��\|���ιݮcvn���\�s\�r�uC#��o��u��nݻv�۷�X�zBvJ%Jh�o~]��М��Dmˋ�ƺn��	�q۔b��wu�ӻڹmxܮU;�Qsmwu�0K�ΝkE�n�a�S���W"�\�N�k��X�wu�uPf؄������-�Q%����V1�^6�����DѼ��<�ͬ�wfgw]�]�������.�ے+��+��;��wvf��<�/)ܮ�ܚ�������s��ݷ#�.��Чw.)nN�nE)�(��B[� �swv��su�j��]t�����V޹w���`t�wmӥ����oN�{���,Ecb}]�袙X�n������"�Z�nQ��d�$�M,���Ĉ�yv�C�W"�}�1�ۭ�sIP��{�Ј�A�<LM���J�Z@B'�%#�"
��h�X,���i��;!�br�̔6���0�rܼ8���IĒz2�d�]c�)��E;3I�x�e\�t�p�5��Ih!� �ψ^`(Ip<�$A$Il�6)�D���A�`�3
2̈2$F��7!$	���M�� >�>쨳���ǡi�ț���S��՗�{���A��r�ߩ��!RȲcr�����M�b�䤆��U�k��7���	�tv+�ҥ�;ys����Z����J�c���B��������;�����3��a�=�rõ�p�^D�ɔ��ۿwJ����oB��3����^���bM ��p��e� o�����5(o�Oo�3������
�ek�h��c���jӀE���q��{[��9��<y����f���N�.�`uO��QP��=�#M*o4j��)n�%� �:��a瘟9�.WrWک�H;��A�r���s�}۱��qyU�꺤�`��{v�@�� ���P %U��u�G
��a-���v$���tdv^�aA�¸Ne.�6�#Tb�P��;}�3����Q�ݞ��U����,��4<zn!�٨�U���y����ge�TU��UB�_\�t'�����5I$fF��Q0���O4Le1�q0n��0�1{��u��������5g��*�D��@I�t9�
]���GR;�����3�Fێ�ϑ��xN�ɚ�Gmzk��ot�Κ�V�b�J��Q3[+g�<�֜s޿r�৊-��|Hm
�A�Q�[���{8��*��m��g���xŨ0���ہ{FbTqY�5E�i��I"v�ᡍ���r��X��}��M;|1�8�H@�ƞ������Tl$/����V�y���|:�'����Ε��Vr��1�L`)�J������eKU���A��r0]u�x�C���Z*��~�IWW���/v�Ύ�ԻTw��nz�i�9�䢟wQo=����5�m?z;��ݽ���9�fc}|�.v��*�� s���VZV��l�z�1.�W0#TGް���&�|�ڊ��2�T�.{(����5�d=yk����e�ꓨ瑹����|�l��U[�cJ$��~�V9�HJ����zz�swZ���idM������o�{X���2ఽ	��1g�J��A`r�����N��\�K�\�7W�]̂�s��3�~Q���CT&���3�*N�a�\�����${�;�ꓽmvK0�+�ىn$�	T�wTzd䒳
�ar�s�2�N�A�Ȟkj�_�-���� �����yP7�����zS5$da�Z՜���&ˁ4&J��p&�ãL㰰B����:���]:V�HEoJ�rw��^��mc]>X��_��o���~��، �I
���
q"fw�l���{zr�W�dbοM8E�/E�!;�h�^<�no��݋�wP�n�7�����)���K�^�f�tB�[J�j�|I��r���ft(�j�2*�.��ՠ����m�j��z8�c�H�0!�R�[��.ˊ+�������t:�3��ْ7�����/s#f�b	]}�D��ʉ��*�¾�I`�|zd��GF}7�o;�T�����\�?]��U�i���k���%�ت�W��U!Q�gxE
�F+F&d�!�o3p�j�,*�֍��O�w`x:X����~����}�/�@���v�ò�S�[vz��T�b����J5s�t�����y4/"GsE��d��v���:(�0L�|�Ek�8�ő;˻��v�B-��[�����C:y�B���yBl�X���їݐ�ϭ�y�v{����e��ٺ�w�z�����	��;~���	|�Vy���'�RF�=�;���R�uj��[W�����|��h遚7��\�{+��Js����AA��jF-�s�\>Nhpfw�4'�J�
+#��W�}��BlN=�������{��:[�������e�ói�a�\�8N�z�[��}r�Zy�Ӏ>o0u���B��[fh���MN����:�}C7�#��*�y�N]�!�N'[��2�+�-g���4v�nnA�r9m������i��4������e��e�$+��������Q4ɋ�v3Vp������u��m�˜0��ް����%�Y�Q5�{��)�ˊH-��lli�����m��33̆��W^E�u�h��>��zaY�Ъ�w��7z�.�\��\�pN�
�1���U}���͟*��5�̨�êm��|)��y@�K ���Es^��P`�U^��3\�������.a��Mg�H6�^�1R�����/ϻ��;A�;W\J��j�d^%!�r�5�ϳ���9�dѨ��p>�;�$��f���WWFM��`]���P;yU�Ak���iۜ�0
u�mt�,��(�k��3��_`ܩ�����ZVq2(�.v��/�]�x�؉��%�P�2����GJ��;EsE�h�*��û��9v��Q܀���%�pk��.�֣�) c��t "9�O=^*��a��Օ��Q|��Κ��Hs0"�5}o��B�p؁�k���Rr/�=�>�Ph��W�F=����zp.��>�2-���X�pE��/����=�UN&�&ә�]�>���gK:+����go��3��s���-�A��0���_S��������4�9hHq�x-�@tV���ӎ��wZZig�w9r��|yY���IĢ�DM�ro!4�Z;�n��GM��/�L��['J[�^qu�T���;仛��.�A(T"��U%;�Jo1Ow�K��q�k<���qs�O{�_���9JE�wi�5�UdDrrF�#/hMo]WT�������م՞7qsېx��n���~�	��27 �Z���~R{n�./33�YR���7-"��w�QB��Τ���
�L�۽}�p�9%k���i$E�N�0�h�vЊ��U�,�틜,����y�9��W����h�v�:M�y��>VK�j���|Vd��/OC{a�;FON5b�-y�ͷXR�gڼ��ӊ{jǾ���cUX�Ky�%��Ԩ��
e�~�9G�
U���ako�ׯ��Զ7������s}p������� )�1�0�ynד���t�~Íϔ|��n�tTyǖ��(����5*�U׹���O�1�ɞJP�8RL�eg��2p��X�\(D�&L�Q^�Y��j$����Y���yL-��2�J��|E7p��=�w��e��^[���pɝM6s��E�? )iƒ6����wS�kv���`�W��"7'��W�e,
��:ښ�$���^ �e]�����ί8��n���H�P��F���NL;��]6�WL[l9c�9|�M>��n���0J�ry`����O]N�f$b�ܺ�����ľ���Ĩ��W�Ȅ���O��:R�7���aiC��[8(�:��Ĉp#dGv)�Y*�9Ӆt��]Ж��u��׹�k�K�83��4#}��U,8� g�Ѱ0���m�(TO<�KTP�F�u�Ӫ�;���!�Hzj*�ت=3>2J���'8pT�����<+��^���Շ:�M�����
�H|�
;3gD�n����VQ�=�=��H�S�U�3����*G(b���N����u6�gEai}[z��z�mgni��������ܬw�'��kB;���(�݊c�
ιI]�P-�Z���������2K�(�%-47z���Ps����m��8���D]�X�M5�_\r9;���d�a�{	�a(ٍ�nܓ�ŝo��u+i=YM%&Ŵ[6�]n�Nو��<"n�U)�1����l��~*���60=�LґG�&ț����Of;��<*LX�19�"�jt�3��榻�UP��Z�)��v��+S�`8��eGR�@����튉��H��*7$h�̧l�j��.Epլ6�Ü���(m;�������WPA�Q��c7��w	�����>F1�^ʹ��8a� �0�ݻh���+��m�8��y��s��(OeW�ۯe(�JR$�׼zf�P"��O+�8�_m�ID�r���y�z��k���m%�z�܏h$d�Ꭳ��*	Ww8]�!_*{��+��"�,��j�2k{�c=f{��>�V�'��q"D{��;��S�cydW@�5g��kPk��qX2�=^�+� }�=z1�\��s�,[���9:�̕u8�iM!S�%Vm��;S�x��;
v�
��c�pSu��"���q�vz�������B�D��R����B]�l�@g�2iS��FŸ��b��',s��ty��v���F����]n5��W����v��9 �T4��g�s�[L��j�י5�p�k	[�Sdy7M=��m4
���k���>n�g�X1!4!O�1�R�Y�e%F��㯱fq:e�{r=��;�m��s���#�%z�t<-�+tL��]���:/�U���%z��K.�k�>o0u�6U�W��w���R�K�{��	�׾��a�`��p'[ n����F�*��NA�ТU!����Tb�^�ףf�vU5j�UH{�K��j�r��d\u���A�S48lX���U�Pb���D[|M���c�3���;0ˏ6��'����/[ ֫��Y8�wt�w����e�P�|3�_�����b-(DL:[Y���q�ҍ��껔@�:��Yû��^[��<��n�77r���cz�'���wk<�2�$�u�}��lm����WJGE�Q�Q)ծ�,�c;Y'��b�qnv��V�`��E�Ę2���-xr�ډT���,�A���j*5c��8�UV���n���t���@ӚLf�j���i���b�z��if��Z.r.�B���Պ�k!E�\�E"�Z��1���r^�����8��jqu>�9k.x�5�����G&��HP;��sX���z���]]�c��z߶,1%�K��V�3'NHy���Stؤb����ٵ��'o�u��Sn������@3^�øC�3sURq�f�i�@w���RΓ��O9gs�<��:wڦ
3���"��gTwQ}ӵ�\&`p�0Y��<�����l�=��-U�l�ޛ���kz7��|x�@����l��@G/�׵��UuI(��|��͞�Ը�t��٪���~�~^C/���}o}j݉<��];�����l�S=j�s�܋9^U��(C�']�C���u��&����P�d�a��3�6�^_9d���r�>g�C�;��=�g�c����M�|����;j���1�h�3eJ��t��s-��	ᨍ蓴ԛe�E�w�z���5�ݽi%&���+e��ʻSh;5DZ��6:�]�A�v5�-�������uΫ_mj��2W^՗��1�g3��0[J��ރ:�e��������¨�{�sp�J2��(l�jIxM�7�7s(��M;z�Ԩ�C���7uײ��y*t��}�Oh�5����q�F��s�o%9���Za����)Xx,�x7��.�+����q�۫��v�,A�L��w�x�r�����3F��HcZԵ�_^�D�jAG��e^ξ�)�SJl=�I�����uO��U�6��{h�i���*��hغyoH��.�����<%�^��K{R��i��]rcn�m����	��wT�b/�vr�.��Ty�1+��f�:ֈT�_Vn�"�-@�Iͭ�U��b:u1x�m���BS8�#/�Qy��N�vU��Jg]b�b��K>ݽ�k�Q��,Tֻ��g��_@���ͫ.8o3q�ևG��뙘�d�6�UO]=�� �ֽw�0�Ob�}��:���D�1A;6�d��ݩ��E]�j]tF�+z�4]���):���T�9�Z�eh��.�6a�*n�f��*�H���juk�^7�>��7�=�0�a�:I����"�9���w�Wv�C�xFjn�<N{����O�~_;����|��u�4�ʗ���g+��h��v�����JOƧ$a70���f�n4Dj���'��R
0hl�#A�T
��W�nf�2m��]��l�.��Rl�9��+$��*�����\��1i&��ˋk�/-jf��j��n����l��x�f��q�8t�-M�ob����*��p�sI,��������8�s�&^�ix1�femWn����i����AL˶�°D��Ɖ-:�$��#�Q39��ãJQ]�N�f�Y;�o)�*�[���!����ϗ�L��B������'v�4�{N�;�p`���8�;�V��U�b���o9��� ��<�X�]�W��>[)�c�4:��V���:�kQ��h��V��I)؝�u�i⡇P�0&w5�r;X5�m*��ee��s65�X.L"،a�ʇBn��K�����;WݚqD2��m�fFF�=Rö�I�Pg:����N�{�hS۶"����u�Bo\�u�S5}Ls�Ш������6]���鐶h�'	sN���{�H7 ����'T--��t+.�;2,ڪ�6Ćo+#����]�����D�>��J)�Td�h�k6������K�m�DDx~�͢��E9J�TI	$�ӷo^�v�۷n<x�ǣ�Y!;��v�Oer5�.�o��Q�ٚ!$ �#�Ǯ8�۷nݻv���|�����M%�ƅYF�We�L�Q��=n���ׯ^�v�۷nݽz8dd	��.q���łg���baDQ���"m��"�o^�z���nݻv�����$��F5�JH����A%�`�Ѩ����I�X�ۖ(�RFA���]��<u�Xŏ�����*'��Q$�������YO;Z�c/���(�l�6M�X��4F���y�26$��{m�&�DE� 4Ġ�h����I�A!R�.ilT�E��]���P�ݲ���Nɝ,�����*�¶-)�j'���}k<�nM�73���z^r�{'_X�0#�\�<�gw�dR�G��Q�o�ׁ�|�s3�� o##�or��=A�N�X Q���ܺd��I��Ծ���~��4&>;�&���u���Z�)^W�)��yհ
�q�ku@3���<�7m����<,��\?�
>�x�X9�5n�__�|���jU�]�C*�S��[U�H~������Tbm��:�c��x��3�{�Sy� ��Xd\��J{ov��5'�����$t+�Y;:%8^�."�[ax��/#>�XW�i5��f�[�=v`�sb%�.}��P<�G��.P�P>>n��r^w� a|e�1�+z%�r�K �t�/��� vi�yQx��v�!P�4��n��T���^�,ŏ� Ql�xX�Q���2o��]%Ǽ�&5>N�~�����t\�.�Mw��{�k�i+�Å8�Q�|�7X��
w'��$oV��ꈦ*�t�Q*y�1�p!�hovf\C��W��� �a�h� ��$#�Di'����c�a��~e�ŧ���so�/1:����=�mG8>�u4��0����`!����7�l:���=��x�L]o�b����oJY5�H���p�y����eQ4`�e^:��Wd&��.%l,��eDK����W3gaTzO��E�s7�NK���3]&�[���X�;��]r��m��S�R�cl����޻�{��Ɇ`���g��lbF	=��}3�y��^e����	8_�gw�aad�0u� C&3����.%��Ѵ��W~��J�ǆ�2i�_;9�t�[���=C�����4��D'W��޾_�>�.Ԑ=;�{fOy{����!����`����;5�@\_����.����q�#��d4/�X�o�:�����\!�{[[!m��\������&oi'�������w��O�sn��{�Tf��c~l�'����=�cύ����a!�&߮`&�������^���N�$�r숸�c0�J�to/��>àW�W�x�(�#� )?�r�"c��+�K�:�@�>M����k�&u�V��)l�w����3���'fd3�A� 8܀� ���-�s�>��D��<� ["�����N�n�b�N�����FP���|��h`RY$5y#>/)��0}񱰢'�t�K��@G�I���)K�9�������{�|���3�`_�a�j ƒ��p�y��u
b�dz| ��}!��*�CJv5��W��D�ၬ���O:��kH�ƌ��>e����sbA|������f���O��׬%^��)�Nc��}Kzv�힉&6�]L̮Qө�C�uo�VR�]V��^��Q���1�����`8~4�#א��,�Q��>t+FJ�3��*i$��5�M��q�z������&�Pər�������ga�i��xު���g���RS������zrUd�.o%�e�/�;�[\��w(��r��&b&�� V��zg�E8�����X)�g�{+�g�M�z"[ɕ��*�%8���mꙃ

�l�^���'����/�m�!����8�pd��4��'��7eRc��	d�v�jz����{�����6GX^ .2�x��A�+�������2� �{�$�sS�8n!�R6����Lr��Y=�6H+����cN�������~��גߵ�)w�@�a (��0���]7P�&/��Mn��� ��� �y��ϼ�i	���4P�}��@�3��0���<�yO�n����eu���.hz7*��&��aMM���^Н|:E��qv	T[��c/�����MY�9R@01'�k��M+h�O\;Qu�<43ϝ��[�Lxct���R����a\zV���Z�K�n@�[4��57�u(����c������/�|@�ag�4O�랯ޟ����p/�i�#�	ʭ*N��+�+K�)��x�8�&&�bf�%��`S$�S�!�{G� �'�����v`���ǟ"�&ob��=
��!�p�� n<Ӏ�������"@���!��� TD����)�C����Eʨ��|�6��
��v�P�"��{3�F���wD�8�l�?Ck���N����Vb4/��;���2!��A��M-� ���gR�|[Ưa�f���7BP��n[6s/{���M�8^�k��fe�rĬ-0��.L��9���||||@o0��7��,O��Y�/wE09�z]>omA��%�0�D�b��� |�"�|.8�S�s5��Q�\��<<5�-R��^Y��[���3 /@���F��}q�髦-�>ז}Ur�˽xB���������>#o���P�	�H���Pe�:/>������}�Ȏ��IFk����o��ϰ��(�`��}~2D�}� }�>c7��`��vL�&W�J�'�3GS�r�8҉��z�w8x�u���n�	Ĕ@�v�,N2olȀw<�|�<Ͼ��� �8�g?6	jʫdkDq����K�d��`(T�c0ENc��L��S۸"}�2/���'�f���~�g�8����>��x �?�yoL����/`.�cE0ny���ПX8/�X"m���[0�qW1�˻v�/{ã��:=L3�:���):a�a7�-g�x��������S������w:�)c���N<����S�}"M{��?����K�zO̓���[����'�j�eѤL�Yxy4+�����<�N�ǰ4&'��*t�ay�PY��޵�8%^��ْ�a��D��г����QJ5NL8�ZzUI���ڻ�A�eɯ�EV�Gg*ٔF��L(B��Y��Uj� f��V�*$#���Om���E�g4��j�;x1����-g��OmbUB�-:T��Ô�,�ع�Z������x��������p�����z�ةz��[}n��c	������s�A~>��>�GX���ݮaCyH^}'q�n�ڪCWT?x{���>��yI�����|��sD%&���h��c@����|��{���K��R�5�A`G�<���r�����z0�wC�
�@�܏P�>�\'�c���
z��O��q��� ���a]�*>��	P�W���z �v}F�ic�{�{htx�^s�3=���� 8��8�~�&�"�^���F�g�p�0B_���>d�l!�]�h�v}]پ��҄{<g�UY>�tuZ�w{��ե.��l`X�iiɓ0��^��[��w>�֡W�����է�D�'n���ܴ��J ����[�����a�����Ɍ?��[�N�R�C[���t���o\E��4ج���d4���k]�u�~`1��� �Q�_� P�}&��}_C#9��;+^�Ub�C�c�0K��g�&�j ��}�Ր��g�Pp�OB &���-�r@<穛6��0�qj�i/[���({���mi����%�y5�������?0߾�V�i���^
E� �9������υ�Y/Eke���gx��Ybv܈���*n��q2�a�͝wU�p�KVX��Vku'�١�R.u�O�-5�F��˛:̆��y�p^l��T�&�&om9�m*���g�s�V�t�5P.�'�ܹ�ۗ�~l�-�`F���)�B$�P��󙘢{��N*;�a��O��	ߘ��x.IH�)@50��vع��u����SF�r����ql�U�[~A�����vAoCԩ'��N[�۠Q���s.�92أ3:8k�  y��t�xضb6�����CV�2���>�v�n*�c?`�Y������F�]��yۭ�Sȣ�	�ng�9�x`<��v_O�
Q�-Rrq�Dp� �2��ۡ�1���|�'���e��(��~����/����{}
��S���WU����=��؄]�`.��%8�-t�x�ڹ�*��������p�#�6 j�2$^��Ŀ���i{�a�g�g>���p��H��
���b;9�����v���4�F8�w��$���������Ѽ=����l�& M�Ϯ����7�vgB���/�M0�-��k�|_��ŉ\ �Y�
ar������M�G˥Ԯ�j@�h�Z�{Y�	����Ə_Y�[�%��0�̦4g!���ߤٗx��]���~E� ������r�D�om�� �M|���Mj}��	S��IgʮuJ��1X�-y?a�Wyq�w��%UT:�z�9�MBl�meʻ�2%��cw:���t]�IJOz�4+c��f经�++,�8�W���q��ܶ�t�N�r���Ԝa@�eνƲ�v��M�'	�{k0�h��Uj���oƊi��F�A#h�B�<>|��o[��~y���p��Z�tZ����[�'
T��!�o�(�3��ƴ�sE<��>e��6�y~�ec��:�%\��%}��T]��^�/·!LU�6����{,�|��f>��G�g�t�K��Ч`�����kɔ��<���a���m��؎�A8�P%�]6�7��ێ1M�c��#"���#ue�!/{�-�*��8��`L �� ���@ac�ރ�����nȕ
u�%�츶�f��f!mR���|����:g*�n�V�5��/�eL ���p�PllwM��oDJua%^Wb��Jjȴ���������1���h�0����a�`>��_@v�3��s\іk0Үy(gG���G�~��AF��D�[�!�c�} :O��9�[�d�g����='��ph+�����wT��`��X9�4ӳ\�S��?_��<0��hN[���f8�ϔ�ӳ:��ۺ[<��k�vhf�����-Bo
�rW<�7)�Z�
�Ƃ�P�^`���� ><��h�
Tj���\�:�[�@� ����n�sL�=~����U��4�1�XEt �	��t���A��M#�]��$u��w}:�{/+z��ˑ ���Fem�5%��-[���������SՓ��p͚��)b�����CV�Q��f��0Uk�LX��"/-`���._���r0���5�����s�<�3^s�_о?L�d#M*SM)Ҧ��n�5Q���Z�c{ӷ=���K����|� �L��8�c-���O�����Jײ��%�*�a8�[{v�L���\[+{wR@`�����p؞�<��]�0M��P�z&�6Le�q��T�Y�7�b\7�I@��\&g�K�s;!����p��<�o��E����͒��`wZ�*s75i �=���/�O^J��L�C��W�K]��a�>H����Eʻ��w�����8��$Br�ם���!��;`T�T0���O�;g	�#M<,�S��p�Hhj�L�'����omV伶nG��@B��Џ3������N&��vGX���yx�����#<���C�,�S��K�����?@�s����#{�\O�����3�kr�o�/�=�,�ͩS���~z�c_�q��0�d�d���&�0%�(�*m.�����[��q� M����=�n�(�j�<:Y��-���G�7�{�A��j�Ƚ�@yD̜l��������I9�e�b6s����@��x[&E��Iطs����6��تw/C��F��Ů�/jn`�
&���kJ*�um|�s�Rvs�5Sd�]f�{�+:9����{�(�.�F����iqPsc3�ʊ��2�����eMԬoJN��15�c3q���T��g������ZՔU�D1e0Ո����Ǥ��J��)�Z�iT���"�(H� �(�3^w��d����;3E�<�|��x3��9�X����6R�a@T0�p�6�e>��Ǧ�Kd�nđ�����Ùz�0vJ��7���U(��Ϟ�U���(a~�4�!�k���O�0�u]�0��6��:[��70t�0����l�q�9����-?5��.��0Z��KԾ�'����lBŅ2r<$4x������l�<'U1�5��C�Y[&��k�Qu�Fă~�h~�n���;:ͭ� >���/�̀OO~�؀�����"�~��ͩ�,�ѻ\�Įz�mzği٭O�(��_��\��*�����+��'��}I��G��mZ��i�u�VMb�����6�'���s��ӕ����n9P(��+G@xB/W��x����ը[[n?� Gү�B#h������A�6{=�8Xh���������[���?Ӹoq�bY� \���E��Z�s�ȯT^Gt=07��A�G�f8�R�l�'%Ov�S�d��!��8v@���!� �ץ�ގ����4&��t8}�gO����)ۈSbV��pj��J���kh1�O��Yw��޺B��[B1P8n>�]�[�׏m&.���5�^�=�}f�v�e�:�#���r��ު��r�UǼ�n�Ē� �y���eQ��]�.���G�8mp���^W�_H���~�T��F�{v�\��Sv�m[�V*��0��h�)ʪ���;�����/,D���$2�(�>P^SuG1S�皏E2�dm�K��A�շ����qx+:q�j����i���Τt�w,8� ����)E�&z��2Q2$>iXr3��>�C0A+��M�F߳k�KZxO�.��8��8�oUl"K�?����H��Qc�E�v�fQ_"ݞπ�\�w@�8�5���S���=��8Ul�hЦ�m���s�:ض�x�5���w���
p�=�T��a����s�]ZR��#)����#���F����C��s8�t�=��K�x
���>���j5��Hܞ�;�R/��&*ۤR�'�[�SL-�_3�Fj�@�mOD�;ַ�dU�{r_Ϧ5�z��^��Cud�(�t��-�徇����R�m�d՞l&�
�^e�P�>/��
 c�ws���^.�	�c�<����?�P�WA����_�j��T7�**ks�������w:lw^񭝂��p웎�xrb���k���d�T�͒�!�E�s]��)�Z���cVW����u����
� J����s�<��]���Bh�&E�M��T���ۢ�F�V,k4�	�/��5�C��u*��b9Q���J���v��rZ#$�ӄM(4�n��1�1�.ۧBn�A&�%-Y�0pW:��3�fr���V��ڣt�=:��P�:�㜴��nodf ��c6Z7�f��ާL�Ijg^��@�zl�9�H%�gB5��]䤠�/�/JTQS6�;}٪]G\���6;�NntF�-���QE�T�/+-Yf]\���xysC#]�j.��lgM��N���Ua�w9WU��%����>�Ϝ�mEƑJ3R��4lc�+6�n0(I�!��t�x����{��]�\ ����j��r]�Ъ<���m���s\�N���D�*���TF���Vۗ�8�Z0*JK3sH��D9�<F��	3pN�gv���¹��Tir�u��!�U\nY�S����:y|���\�۪3+�4ʶ��ZG
�6�A�3W��YY�_�v呹�h����uT�ɐ�W}�J���V��m^],+����¢	��>S!�YRvХr�S��w�#pÇ�ZV���7���eyE��X�u	Uƺ�lhІ��ש=��X���rg2F�I0v6�-���LDb*�BԥFk0��n��]U:!Vb�:M�w*�9��f7��Y���]*>5Eke��y��)�HX��y���F?b^k�:7R�*�;���r��":T�_i,�v۬G�˼�L�6�ͪj��e��Ҡ�����SJ�Q��x��[��ɩT���e�q{6Xܖ�4C��)\ϝ���\޻B�Є$�����5�v:�*��{]{\��	uGSA�.FN�ʖԃ���dIs���,%�ڳ�,2��ڻ�Ҫ�q�s�k-,�^d��2�;�-b��qfpoL����\�MK����i^�,Hp�ZN��w���ek=�����x۳�{�.4җ;qs�6��Zu$�Z�h7wҕk��M�"�2��lq5P�㑂�ȪoX��wt�N��(f�8�u��̧/���pn��F�P���$�U9���;Z8I����{���h�2�aW�T7{wׯ���3"����B}̋�B���j�vvʫ�
R��܁�.�0�W��_D3 ��+���{NU��[-m��������M'2>`��ycZqcw3x�s	�߳\�Qm&��S��+�t�f�wY�)U�X�����wr��8;Y˻�%�&M�γ����+.��]v�en�.��)��.���n�e��yG�z:E+�8v3cWBg��11^���m�#�u��VDn(z����U���֒��[}���̈b�EH�/\��!:��Z���z���U$
8��tH��n�P�(G.aZ�����S�'	�h��T�(��lw/��"H����MF
�6$��F�å�����|x��<x����7��߾�Iwqh(!4��dh��Z%)$�c�N8�^�x��Ǐ�z���FQ1�m�c&J���,h�����q�;z��Ǐ<z��D	!$�I�`"흖53�Q��Fݛ���{����޼x��Ǐ�z"���	Md��F��n�#"X�H�J���5��$-����KdDX�h�1�/�5�A�Tb�o��3cb���E)��D*5�ȣzn�k�TZ�+%FH�}v�b�^wlclQAl�b��"�F�6)�$A�z���P`�6	#`�R�����j�RJq�H8�D��h(��!��Q��nw
�\�U^!`��myeg>ZA�W���bf�i�$�H<�[J���Гh�-i�r{7.�UdB�F�(��"*F�h6,ȡmY@��'J�I4M�/4Y�(�؄�_�4E4�5!ѩzn�UU	Z�T�W�*~4*�Y�ݻm�՛�kZ���B�J�$EIP�@���anD�2�c돷0��۠�@�T�b	�Sĕ�n�%L��D+���9?��A�w�d�pC��?)7����Ft3,Ϭ<0���>�`oW��O����^Ng��X���z�'�db�q,�w=4¸���4��M�y�T��[����V=2���5��BY�=��gt޶���d��}f���w�ZQ�eR�	��p{S�2��v�;7	�|�}<6�B����q����a�_v0�-����T�L�v���.A͸C�-M���P87â�Zz�m����>�@a4����9�ȋS\�g	]����Z�k�m>���A�T�������;{,���Y_��*I���GY�i�DUԐ���|vp�ˠ!�=0}pV��m��@��u�N��	b�M��1��@���G�����zү�J����S�O����';9z�^t������t6��]��i������H����F��dC��z�s#Q��)�x�ގ�"�L$�7<�&�5��Bn��xN��Gg3+&8�r�hk�qO�l܋h7����SxBN*�SQ́��qY��2-ٟ�(�����[e��r�Ն��Ḝ|z���/07I%
��؜6b'\�y6�t������`�C��U�uZQ9�e�tv"Q؈;�k�(�P�Z�t����̽G���sR�#7�[������9����vC�*
$�����F�Zi���*"��,���*2 ����js_��s�}���9���"���Ckο{����������s��:��F�'���\�6!}�"�}U��S-u��g��%�7G�.�$��?z Bs���g2ϕ;f;4�/U��V�Ժl��+�q�i����.��7(��Ƽ��0Y�q}���u�+u��]sm��7Y�=�~v`���>�y/��*�1�5Ms�0�V��c6����^�Y�/ogPS
)��à��p���ץ�{�7�70otݳO�ȥ^~�.+�JװT���U�U�u9���I��,�r�5;��0D��x�_�����fT���^�C�z�.\�Z;��8h[��#^r{t�	�J�4���b�o����g��Ap�?�De�C��b�ݶ5��˓5nT�ÌJz&��t_���s	�^�tS��`o�_�
���L���/���սw�G�dMt�z�G�NQ��n���׷���X�p�D�b�-硔�al������r#����|^��-�=1YH��fo�'�+7�tg�O�� �`���a�*a������m�g{��ݵ�[X6�ge&�Ս��hf��;�+{v���*��Y�D�יJ!n����3lL7�#{��1����X�G���A-u�n��hJP�]���^Z�eL1�!�Sh�9\ɛ��}"~�J"i���Uj ���B�� $�(�*H �y�ϟ3ٯ�;�򷪹���5�!��b�h�0~�R)�-R-���x�9C�KwN�O�����}9x�/��a:k�k�Zs�0�����4 �kd�&<�=��Sg��l≓�Ԭ�y�>����'ʠ����JTQ�����m%ĵ���c��p!M��M���2zm��Au��nd��)]��f*�e~R���Y����߾w2�ļ,��g�mNכf2��'��Hr�t�S�͙����� U��c��������9�eL���n��g3�ij}"N�C�F�����ݏ淔�~#�_}U)���zE�1t��c����,st�N�y�N��&hZN���p��P}m�	�o��M{��8�_�w����Q����k�]��noQۓ���4y���������֘���x.�c�k^�"�qT`�Le�$W�3:�9�n����������'��-�K�{r<�aß��ֿP�a�6J�~�C����DHg.��Ҧ�b��f"��F��~�sN�Cb�l�`0b9ĀC�y�a��Լ�҅І��_��E+u�)J�pb�[A��Q�Q�RvL�G��=ӎlL	��f���㋉9FmȻhD����l)ꢜ!�k
�qm�c�E��6sZJ��g�e�[�Y%YSgE�7Qg[�PA��d�����3Z7��#�x{���~�B�h
i�P)����Q��U�Z���UX��<���u�����j�l�=K���;�q��3�ǯ�v��y�3�N�f}�TV�aɜ1�%Na-��
�Ї��Իk��e}��:�ŷ������1H��"	��g�����\r��ڪ�co�'�E^�A�B�OŪ��j�"���er�2�����7�A�c�ʾ�8V���#��0����%���4�q��@>uu1u�"]�B�g�J�kϦ�tμ�ɕ�R���S��sb���L�ee���}��Y�#��)G����252k��-H�-�ӝr����ʒ�`Z�9A�f�'Ʀu���Ëh��E�.=/(F�Fʓ��^.Q��[f]�vcj��I��j�5Q)��Fcз�x/l�a�agL/�7/V����m�/Do#r͙֑��%�r�K"J6���<Iݑt�f�o5�p^��1s����� s�8���+ h���]���^��[�O��<h�hu۷w=&�#G�!
0îo?�80-�AR&�)��
F��8��qj�r�k�c��驷��쩈K�I��3�N�#m��6j�{D��lP���`�BUS�"�[{ ����Ŋާh2�S�"���)!�}�VK��ҮT[J��^h�NN���{%�)��n��J%�w>�vj�n���*��T�T��L��KߗeF�j�מ}*	��)��V�iV���	iT��lmVZ�ح��cZ�@�	��ٜ�9J1�)?��<Ǭ�.)�T��rӪO�_��a�OW��CO�����|�#�v[睵0͑MB;�r��I5�u��E륉�Û49Çt��Q��G8�vZ�Z�,�a�a7d����0�,l@�Ъ̞x�P�A1������� �;�Ƕv{e���E��bs��}����m�j��@�����<%��n�k��IŮ�/%\�T���n�1�2V�^s���9xs��y�8����׎���?�е"�B6��Gg�~���@uX���I�7����g���A�O�z�<T�=9\:���ަA^��^�����D,���/a'İ>��;"N��nku%Ff��҈��}g��~Ŧ�+	ɕ����m ���V�b`&K 6 ��d�����m���F����|L=�H~��0�]�`�?~�A���mz�*j��_g�rC
�ݮR�X�0Q��j�׆l���J#���o���Rz/6���0�����5��f�,�����u��Ϫ)���N(n�-Ed�֓��`ױl��l��%�ݯR���5��ܮ�l:��mbٸr4��I����ISW�+�»�T��Za�]�V	�dӶ4C�+yD�w,P���}�=�`�6y��F��-�u�1M�m�K���y�Jj����K�RĽ{F��Z�b�ccQ[A�L��p���,~����TE�$F4Ң�KZ�v�[r�-����m�@ ��y��E3�:9�>�]��zq�nm�oAO�}�B	�Z�,���Ƙ�qՉF�Ne�ą�K[[.U�fO0n��K�!@>S�g񞵅�|֬�,jҡJ��l��1Uv2���[!���]Qp�Ol�8BoB��>��"�p�>���z\M�/v�͝6ʛ;w]W;�e�;�!IN-�-���B�Ӎ�l�'�y�ː�呌CTc�c�>aGҖ9���l�c�Y+�E'+����s���"{1������˞#y|�?��;Oe#�vu
�C\���e�:���Ⱥ�x����GQ���^��c�KD�N֭aq3]Y|�Hj[���D�|>l�8�G���
���H��d�yj�r��
r�gL0^O�,D��z��4r�d���\0~m������]`�#��x���*�]�J��\������n�-f�3���	iw\�9�����8P���YhʑJ���^��X(����T��<��,U-�����˪4��sM{��Ә!p~'��ƘY�-�Ef�`��y6Le�۸z�u�<���l���N�b����q#�-�ry��+���W���y�7:u۵HS!kx�ۊ���D���o�*G:��o|�f�UF��u"�nҊ��g�	�PQ.#8M��F�3*wTʭ�}NUn�I����[�s2I� ��~��i��1���hT�"�H$��`"*�o>g�u>,��sZ ��=5�`���hsq�/���z��9�<p0���nH��k�b/��SWb��t���m�V�t/wI;�D��tE1��-���;�@ǃ�nV�ǻ�3�g�&�Bi�
Qy���$;�e�;�{���l��u�f��*$�u9R�H*�a̸����*��N���<4��`����\����
�7�r3�B�S��8��M�mU�Y���,����BC��
�+�q?�Tc�T�ǽ���l����U���>Nnn��1��C�+=���� ć5�L�D�<�
%����|d�d�c�-�ر7�FmEN`ͤ�ٶ��ds*ҡI�J�y�ޚiᥩ�� b�Bq-wT;�f1j[�߳Q������Fܘ��6�x/$�w�BgU���Ǡ5�=5�Ё��e����=.������%:���y�Q��(��sıNBئ4Q�|��G����˘N��n޻\��Ģ�kf1;�/X��L9�C$���Qt�̀��.�3�,{غ� cX�ޞ��B�[Z�qQ����JN���n�#�_fgK�7^���S�}Ma�m_1T�ۅ:�zj�A ��?
� ��}����C8��N�7*3�b�=��,J¥�T�����Ք����3>u�L���$�D=�s6l�Uj*��j���B�h��v��&���Q�R*�"���Ù�:|3�7W>�����}3^�?-�0l�H�C��8��=��?4�C���*�����;�{�����7j
X��������uy9��мE��ĭ�D!��^�U.���lRT;��@�^��ېS0�a�ã�:��xlY�mB��jb���[�!m�їE�q�P�T�/a\
�z��N��2�f�T�g�S������L�E�;����G���!̭�Q�cQ����K������r��L;��q�y鎗T���!Б�0���%۟)�%۝_D'Ǥ��<z�����\&��Q����-�ʆ<��ۯߡ�k�L$c�ʞ�1aH9�I�/��d���l!�\���;��
�M*�k��r�������9��b*c�=��h"��]2O8�s'���t�۰s}N�v�Tg�䍎i��-5�N7�Pb�w�G4��}a�)���xz��余uN���uI�uC�X�v�nB����$r��l�ucs���#�S�-�â��Ϯ~��[���b��'���"=|ZD:Aѷ9IĹN��1�2Uǵ��/�C��H%e�Yb��ZeE����l1�G�H/��K��	#�T]�e��[�Qu�UA")�H�A.I�T2�����DD���gd��;3�eδn�J�Qwwd�( !��B�iU��P*#ij H�"��(��� A;��y|��y�n���:�7F*Ҫ�,�9�)1$����lc��øh^��ȟs��#ڈ��cT�ɨZ�OA.�`y��=oV�^�˾N;�1/��O��e�}x;��1^��* o?c�J1��p.+LK$���+Tj���=�Y6�*���K��Em�l�6�����I��1��B �!�V1�S���1/��]%[�[>�]�tګ��4n�����na��+�<�d�g�9���m�C���u�I�Z����~���[�z��篔5h؆��.1�1���� 7��׏[�@ǡȄ�Sm×�5A1�٧	s�l��� �b��{l�^F-?$�9�iv%�{��4/c���ZD9�:dP��,%��L�r��t'�Z���B�Y��,�La�Iz	r�;� �;�=������U��ɢ���#zZ��t!�2$��0%�cv��z
p}k}��X�*�2\Qǂ��"&�?���4ITx�|�LO��
�~��ٵ�>	^��;b�5���0�Ѭ���	��o��������)!1]uJVwI����	��d?
��<cX|�"�&̌�^�@8��M0h2��baU&5M��iX���$�C���s�w�������Ŏdz��%��F����_�q��g[ꥸ�gGN���Gs�;P���%Đ�fꎿ��Y��iZ�9F�ڜ0�����V�w=�٨Ү�f�YJ7�8Z���_���5���|�W����Mk��@dV?f�J ���* ���
���*({�f�����!�js!G�u����5q��8\�����7��X��+ߗ��P|����Z�D�斗Иg`�����8�`RP� -E�5�cA�� C�������LLrxY̟w��j�DI����cN�.�=]C6RzK�!�Q�0�M��Zk����a���Ř�����3#��?��b��m�q���d�ԑ�Pwئ\�����h,���L��V�b�`nױv�¢�.��h�	>5��	�Z�,�%�3�Z�A�� ��8�թ��\9^�Y1P�^��X�����b�o�:�?*��.�����1���ۚtԱٓ�L�.����Y��ܺ�(�9g�\�(f8G!��I�[�0�P�;1�y�}��R�j���S:��o*�\��>����L4vŴ*&��)�q"�T)�q4?D���]�&�� nx�4��<��)��q�^~��zw�xa#2���(m��Q���*`XǶ��;;�nSmLQ}��L�ŕxs�-8yGf���'+cj��w�lܿ���sɾ���f�w��j'�3���]*�3vv���*eK�p�*�ImfAZ��.�aGpηv-V��.f�o(@��U�$I�9�3��Ug�_j���ɳ�:T��p�3�SA���{-��o��h��곗�%�	���h���ݩ�B�jTGa�;	f�6���j�w���e�W�6��*n�XP��WEF�&���#�N�wJ��Ú4�6�M�J��0-׵VĆ�\#]�Dn�Cif��ӎ�sB����9ۨ�Kh�P�۫6��ǱK�;j$��d��(�q^��y))i\ƺТ�si�mӍ�Ft*�N�H�*�3.�72r3lZ�!�&U�sd����h�ŋ��/�H)��Z^���oOVD{o���)Y��d�˖Aؙca��WEiuxʀh��
��5*�����ް��y�۞�n-e��.ͫ�%^�檩c:fa[����i��V�ضA3*��e�Ħ���R�%�8�]!��M��kfݕa]ԍ
k$ фj0���0���6��1ޮsn�ǎk��k��{]uo�a�����D�Z)Ȫf?6�\{��޴�\�Ѫ	�XԽ�N�.V�Q�Ƅn��ku�D�x�2��9�Dj�4,�\��$��wv��A������-�]�,O�|�j�u�o*�Fh�;K��ɼ��$���zd�_��ыO��抴�������>9R$M��ۺ��ÆD��ݣ/,���t�4޸eӱ�2��o�m�lI[�47��Wp:/z+f����S��*�_fcC�V��)͝�j�E]95TjKen�n��`�n5A���Bm:�z*�"��Z��\Ol��y��UM��F�e��-v�PKZ!D�ѫo�c��;&]vK�T�g"�(s*Y��%����.�2�7pܳ�b7mu�nnB��."�����OάD$�~MWN�T�g�gFc���Ѵ�
�a�;���*#J����B}|�-s{�o4Vq�u����ִ����uܗ���[�!-u�uk�ET��Kcr���Lw�KVҺ�ν��qɂ^�sf��)ƣN��N���`�tZxڟ%L:�o��6\\®]�\!�!F9<��1zh�lgY��R'eӱ9�I<�힣z�h�����b[{���Ldig&2^ ��_�Su���o�K�˨���9ջ]h�O���E�j(43*e��tiٵ���0��e|�N#�}aE�:����5�(',4��S3HP�nlfK��6��um�D��}��&$���N�}wh��j"�+{BZ�l��Ŵ,m����wyEC{���r�ƩE��S[�ᙃ&�v�,mݛ��aI���h���jUl�\]���S���/�Aj��,�� �j����Y��-hٱ<�G�y���*���!�0;�QA�J/�F�P^�(�|R@��ZcN�8�뷯<x��߻���V���DZ�_�7,ƣcl���$���H2B�q�qǏ^<x��Ǐ^�: $��!"H,!���mF+�o{����{��׏<x��ׯ:��H�"ȡ�r���W7�U�0h�RH��jH�*	��qێ�x��Ǐ<x��Ӭ$E��T ���%�Q���r� ��j61�v�4l�7�M\ܧ��MD��W �h����(d�h�#I��5H��z��Mэ�wu�+!F*4F�эF-:j,llBX�ͫ�E�,�H�H��[���^��c��Q�ƽu�
H��
��$��"��w��&y��sq�lm%$��p�5<u����m�3�qqL�nn,۪�^D�2�Ҧv����+����|޹���<~�Z�"�hU���Tݺ�ͭ��k � fqbsRq�7�Ä��~A���>�}.D�_Ra]�y�o\��T+�����؈��<��s:؎T��Rf�v���2:I���}]��ñ��Fx�v;�_�gOQu�WV��)rc����F<^�
c��O�M+�#H�80�*`c+0%`~�.�]��I�V�b�?2���R��uʉ�|>[j09ٖ�\x�"���� ���v�}����0���W�$�6 di{�C~v���*��4;$q��I��:ňL&Fh���
[��y(�B�|�f;8%��\B�]wH���$v	G��s���]f#���*���=�>�𳲤�����{��q0�^�<����f*�/ w:.81z]��UHɵu̫�Χ�����IJ;��?|&��	<4��SSX��<��{��B
�n`v�O�3��_մ�4����<�z�*c�� ���}�
���E���*��[G�nS�s�ܯv��[�J�AP��Y��$\�C�������aAiG8�%��m�y�����}��wXt��1lr�mH��d�ٲ+*�����97n�&�[y���\Tvh4��of6>-H:jE�ӻ�_B-j�X���j��X���vgT��l]�'w8Uw3��u �U��鵽��^w�޷ӾzO���٠Zi�iRn�nj���[�m�ڍ��_��fH��������� ��ZT���l��p�I����K?%�?��ح�g��[Y�hW-�`h��/�Jjމ.��I`��B}w;U��L�����T8v�����+-���!-������H�>��2���<K�E1��&��"��
-f/b,@YFqn f�c�� B �Ƒ�����vI��oEL/�J+������e;Tk՜�$[�w�io�噃c�O���^"c��!6И	�o�I��P�E���R�K��Z�-5T�E�&)�u#s�`'�3`������XD6����!�9��9����yə�I����G����9�F�xͥc��8�������k���p�_�j�mՇV�-&�z��cf�2%�}�\�桼e[ߊ�^��
MT��l[�����%��(au<���=�[��G�'R�N5�|��W��}~�^Wzt�c�
���*�u�Z\T����w|��'��v~P5�92,�-�v�ׯ�}R��Ƞ����u�X�.(%��^��b��ۧ���j�5e�8�G׼L;�N��ݘt�|x꼴'I����:�_#��f���ouubZ�7��#��������Yܮ���s��׉K��9�Vڀ�\"���I�Cv�"e�3�� �����P�QG%���AƳf�!�nFUܗ.���~4�@#M(�M"TF4ЍD��	I$@����z��Z�{;[����l�w����F��@S
�n��>'�G�������C� \<(��%ϵ��;@���L�7���nGVT������݇��~ߨ�)^��鮡��I�n���Q��!P�+w^vz
�����5���^���!(��	nA4�:���*����E1a�rF|?0ջ�����؜/�r�C��-����W�br42��H܇ѝ�O`k�:�dS�-���ג�D����A�଻��Ű�B�ϼ���0�&>��.�`u�~�ב2�\�õI���*������@���,.b{ )�:�6 �↘�I��)�W�Ъǚ���t�4+���R�[��y�=����u,�u�d��`z����&�q�(�Ľ�����I獞��� !�eWh��)�T��/��?W? ��xٞ��A<��-!m�C���\����T���7����G+�@��:�	7��sW��1����ئ���	"XBm��٫��(�K�Qu�s��r>k�l/��iW�1�I��E<�ii��a��s1l0'�Ǖ�r��iUo�f�@~���-��9��GRA:5EXHd�[�b�E��u���Z�7�)�)&�.W�K�#�4�<C��V,O
������Y�7�N�쥸$����'R�q�[�ԣ�K�{9*;�^Q5y���מֲrߤO�Q�F4�%4�njWn�ە��lUb����)SF�
q�<2��"[j�P�ҹ��La�~��'�pY�񭝇sm�QPf\��k���V�J`�]�6��~�£�F�s]�JN(Z�n1*���U!��:I�����?-��zqC��D?Z �a�A�;�E�_[&̊U���B��N��$Ǥz,�`�9�ǂ�;k��f�Q��Z��Ph�D/'�|t���|}ƼŲ\�]��*"���ަ�^�#p���X~�D0ci��,(�L�~���,/[���"�nN�n��vڡ\bS�v�a�@8"�����"a� ���^}�P-S4t*T/��{��>{$�8`��}1f�9�r��#(f�.��|���.Ҟ����9��l��غ�xU�*�#`ՍCM��$Ey�;�Xs�d�Gllz�,[8#��L�,břXBm�YD��o�¾_�J��h*xՅ��k1Q
��w�-�T$�ݭ�A9�Ye�Xes7l����v�V3�\,q71P�[��P.E���1;~6�̋���y��(vd}d��E ��(^�zh�F�8��v�T�c����Ut�k�נ�]����r�:hCܥ�g����]�2��j��m�I��Y�U���$�2c ���7�F�bӆ��˱��N\�#�N�2}ߞrMl�g<��y�gҙ?�h*i��iT*o��y���_�k��W���+�_.!>۫+T��P�_�A	-�
*Ez�ԓ����[Eq�5�M���[����G;�u�IP5
Jqo�l3r-�WN7�5�'I�t�A�Lh�-����>��0;�Je�:HL�7H��
*�?Es�w�xa9�5٢�`Y��{VX��Z\h�̄?'����ϣC)�چ�ڞOc�S"�<Ӌ�F��睎v�HE��Ì�lK0A�ם�F��f}���¨�� ��j���	��{��Zr��*�e�񦶵�ٸ��y�)`��;�J7��!�t[f �z�K��+�k���%�XwS6�p����WX7M3��R�(u�a �����]���1}���a���c~��6���`SE?6�����$ݕ���b���F���>@*?E�~�枯w�i��C��+�l7���v7]�0eX/kU_gM9�ųﲾ/����3f�`��PQ�1м4�@�c�Y�B���<1�p���� lm�eάL0��ݚ�,�q6k��'n��"�=��t2l��AuǪ�nq�4=v�g|ދ�\VUŘ0��yp��˜Z&B��ܳ���5`�Z8���U
6��W5n�X���!�zgi���e��p�1���`�����4�Gm�r��E2E)n�4����e�7A��Q@~^���� ��R�����j2 �a��t��	N�w�B�FI�y�zT��?]�e;�� !�H�w�`�i��]ҧ��&0�F���	k���Mě~��28l��w�S?}
�8E���n5W��O�8$E���_&R�w�TJ�|��g�ϧ�,������G0�']����L��a4�e�GYf�ܬmە9ֆ�s�b����3� �6a�t��HtX��4I0o�O��y���,+f)U����BN2Ƒ�q"U�2*��R{��@�ݽ4��eo�H@�5�K۶�i|�]��
Ц�@W#d{C@����[�)��),:?X�_��R�ӑJrk�۵�x�Kk[��ފs��>me�y댺���ِ�3�͙E�{�%�u�,J�,q�o;ͅ�t^�u���2����9Ì�dc�a���pc+��0�7��������vu�k�R��{��zjֵ�P�
8r�����<��z���^�	�lȓC��8���+g�P��~T�!t_Ê]O�V�V�䠱��L?5y8���>����Y�>���tUړn�I����|#;�S=����,��tI�mS;ZX�,����uW�� ��$:c!�N�;��q(��j��k�)��%�n�F^�mb�����dX�U�Z��*�Э�AI�y+��éeK�rgNQ5ێ������,;����qE�Q6�b���>���ٻuWnݹ�nݮ��f���^ʱBҼCtgP��)�	�R��A$s�Q�����{�.b��f0���up5�����tXu�0��uaa�T��W�=�F��v���7:�l��:��{A/s^�o��F�ȶ#`0hk詍�o$����с�y���*`�`�n�u3�hb;9�[����b@;r(��ΰ�Q�����y[$w�v�*3��"	wml/�]���`���[�<�p^Y���gDh�e���-/$�_W��hF7{�М;�x�;���K�*l���%@d����{,�������,��;ZA�OS���o�P�D����~>;�I�Kսr1�[��9)E����Ǘ���PͿ/��r8f�l@�r��8��!��H�<��a@��5�W��8V����qՁoP�|y�=2� ����'p�$7QS�W�9]�ӯ��l�@2)ޑ��qg5��K�xt[��
yD~��(�� ض�*���$Jk��Pd�-D��%ӌ(��Yx��gRK���ֲg?��0]z�]���-�p���5lkC��i�d��R��:<q�=�k4��{���6$�ݑ�%[���1qR�Z�1��ؔ���!�.�b��[T��+eDn���;�>�i��b^���	�=�.�M+�S�s`��ʃO��NLr�[��a�M�Ф���:J�^�.�c|��ẹ|�������饦�A F������?�����f!���������_���mbO�i# >������Ej/¡cόBb_&����k�̚|�6ڨ�;˥�{zB���O)����#��gG��m"�#%�peK�%�.,���|#s�����P���k��D&*ۤR���(wK�Qs�NS -}L|����H�ƞ'�D��N�]��}��j�޶�u����>�>u/b�q;��|�Ai�-#Nİ���l92[���Nԃh�̄>�D<1�1-�/U
�}+�'�d&0�T�I{ �;�Axw#�Xָ�׾�ք���9�B��<o��A"��1��\n��)8�]<^l+�P�U�A�Bb�#N��r�R���(���r ����_�f	�>Q`Ta�}A|w�$���4ӥ�늨N�V��|s�xg+�;ֽK�u�r�^�h4v��� P�11�?�U.��E�^m[��%��q��"�"F�h���@߁ܤB�2:��Zx�<P����~��B�
^��}/E���9�>�K���	l��g�B��ƅ1%�#��d��\�j��Xi~"Vs�Z��'�E��x�16g#�y��R[��2��ե�fefI��S�#NFޜ�d�0���T�6�oV�G؊��fM�t�5�҈�U&8Y��2�5�M��r*���%�խA�od���e<Qk%U5;���vl�u��_�/<������?��33.��܁�ٞ�H���=6W�=]u	��E�(�2\�\�E�kb{/9"$��f�F'#�L�ld����J��L��·g>W-�OS���q�r81j+$�Hפ9[H��
�L����c���8�p1�=;�N*��AOB1�4\�sl��R��1�uB	�⋼�欼�����!-�aU8�D�q75���	�?!uaϔ�~D�S���XkC���	���x���EVU$�������p�||����i��fƩs��50i-�P�eLbv�^�u٧��7\��+��pA⛘	�c���$�l#��S�~�aӑm
�q��"'��<W3��ă��C��O���Y�f��Lps�,������:�;ݼ0a�ND��:�Y0��b
�!�<怘�g���5�2�yP�}RK��\<ah�-#��ѩ���|��\U���sN&�%��E� u?%G�"��A�ɿ/��a�޾�¯���;7(�ST��N�6�m������;�S^C��R�4;�$Q�ݡ2u=K�uRdu�qq_�Z̽�w�_�Az��n��&�����'(�����{rG���U;����s�o-��2bof�땹��ؐ}q@g�� ��#���՗)�T:�UԤ5�F.��y���q将�P��sD˄��q˱ne�HZl�y��Y��}�_���cT<�{�+�|;�ϗ�nmi����"���[
"}p7��S���n����ԇqo]��V-�~��F�0Q���ygJ�lg��m�P�x/�ڇ2܈	� ��8��G��Ɯ�)����P|wh�e��3�-��a�"�;����3�Ǿ0'	���\��Xh4H�z�k��D�eZ�������t�[��n����-"ݚ�Q��_N�f{�r�҅��g�΋��x�~#P�yuO.����}�����2[��:�.^o5Ă^�����1�����]ݯ���;!DE��<S�~��|Q���T>u���̵ڲ�_zIzl�/x�"6mҞ���y5:��Q�^k|�R�/�5����'
fM'�. �چ�eD�
LV>�?�1�*2��*����	�~ȶ�����bf*��3��o�
��&�ᄮ�QW[�I�i4'���̟>j���d&T-*��vP�z3�iᮝ��9ܶ����[���]��x:)Sr�K�͵>A���u����o/D���%<�5�EP��t�>���x ��I�".�ͮ�f�-�2���ȣ�Mb`�3qm��b��L�7T�X0��p#!b�!-v)�3��ˣ�p���]t_>�2.Euu56��$�"�l[�thՙԈ{�w�p� z^�M�Fgk�k0�6	D�{I3+)�t�^��K�����Kz3���k�{���2��ܸ,��\����w6zu�K��I�ժ�a���2y�n��яx[륷���B�k7��"��x&1����6��bm�2&��S#:�"
�5�T�Zb���72�h��X�S�X�f��[d;�e�۪��۳�2ޞ4�Ó&KI7cxZz�uG�2J�F�-�ի9�6��ȣJ�L̔���qf�9F�PAnl:�YE^#7s�(��Sv����n���d#5�>��$�R����+CD�`99l�T���+z�]�)��5G3ok�Rz�K��6��]Ek�L�+�̥v.*�&v��抾��,�R,�\�`���*�������F�R�!Z�ER�{c&ej���{�5�|�)4鶅b=xܮ1�RP����9rU#�,L���ז�m^;��THJ�c{���n8ܭ�u�=��Dc5�K�(�wش���v\��V�v�3#�6�sj��������\v2p�j�#�e�S}G��$.Բgn�����u�[*�c��W�'o<���WM��?&V]�DѮn�v��Xq�mu�#!�}
�*���NC{�& ���V̖Vm���ot��C�CսRgl�*���QY �̧M�T�4�i�u�n�$�L�EaZ��"�亱\���D_>K��T"mX��W�lb���5����e_q�͵�)m�+�0�@�J�_��r$e�PJ�6'�N�e	x|y�}���U4�Ni��V�n��XBR�;	�z ��7Ngh�mv��U[Ʊ��46"8K��)Қ��x^wXK*�P�ͼ�Q�W�p�&��MĪB��v	�tM5�&�8����7KuқK\�wed��%�2�j�/�ҳ��H�X�Tm-��^J9kPF7X�(8�,V�}�X�w��v�oI�ו�5�6��$�m	Z��)��.)�a�z6���P��2R��[s'^#�kK{ڝ.�Х�s_�e��a5�v��GBB8��v-Ͷ�*��x��S����U;�x(����٠섉A��4t��Y����t�|k��:[�����
���T4�^���l��Z��ǡb��y�n���X�z�ǜ����QZ᫫�s�r���A��[�f��u暾�\���~%td]���"�����V��̭3r��C�3��7���Vd�31nX�u��.��W�����U���?}�֫%��_�sr��{Ma3�O�p�T��5]ۻ��9�l
��v��E�}U6f�NkP��W�S"Qc���}Z��]�M��"	u�+('
e�-�KIF�)�d��� ��nkF��jMQc[�r��FIq�i��q�;~�<x��߻��{ml��7VB�T�m��Ʊ�����8�<v��Ǐ<z���B�X�����),TW�t�"5M1�q�n<v��Ǐ<z��-
"���lH��H, Ȱ� �֝4�8�=x��Ǐ�v'b�I H�����b��Tc[�sR��6F���k����ƍ`�"�ݹ���h��cb���梪,UXڢ�u\�9�睨��h��ssl�[��j�ۚ��ŴQ��\�MEEm�DlcA�$xF՛�a��LF�D �aE�	2���e&��I�a��I���=sr�'uw������`�Ө�U˒fK{��,%3�W9�Vq��oM-����sZH.	$�1��N5j��l������aF�a�|��Q�m9ME>"D�8��H�EJ��$"ZD����#>�)�i����;�9���ޥ�o���2_srY�$pV#y��?��_����x[G?t�8���4Z�T�Uq�>髇����_�̸�3����Y�E{�}/�Sx��PL|ť��6��.���L={z(�a^ݠ���>k���՟8��%����t�??_j�:u� I"����	���6о�'�t�pg�'i�6��m�d8ݸ�u���m?2N[+�.�4�KGlx>Ϛ=�dcW��F�8a��(��v��#7G���}S	���*��%F���w=,��%�� ܎�D�#�U��1��ً����5KX����uS���ޗR#v����A.��s�>�*���dg�os&���۱���L�
`r���b9��-�WE1��CG>��1�>&9�7"��Ju�6�ۼ����h )�3������z7�>U��!ln�~�m��!�{"��y��aK�9��6�!���4/������($t��B��Se�_*!��6�xKA��;�*�a���S�)�=.���!�y�<EL�G�#��(@��.9���&I�g��=�1�0YP���5כS���=�b+���"g�kz�4ᣐW���Q���d���|��>]�N�-��\[#a�U]��U��tg7�\�����u��ܤ�M�(c�1�l�2ռ]wSs���h�����{���>]��}�g>�W�YB������tO�]}P]��Cb�I�.(��J	�ݯ�;���سpcE���׍/�1�OM-ڔ��+ά��z��kK2�-�Z���}�H�Xl����.�{�ݘ��0pZ��"�� Ű&�|����cL�ɭD��+�Y�{�m��O�e�gN���9��=o�&�ṅ8����an�s�YH�:��Aq��|��M���r�yG����s	^1��o�l����H0 '�p�/W�;���S��^��&n[�=�B�>��<ӎ� ��V��b�����;��{���`���UH���%{�T�Tw���l���5OC��IN]Ͻ��-�)P*��5x����x�<�o@���y�K\iW�b:�)n�!�Oe
��QX��f;���I�sNq��vi�s��s��Jb��"K��|�,`��+ʀ���'�Mu���I=(�]��*��犵!1�)���|wmu��;./x�:?�[�ʝ��3�����􏩃�<����U
��CV�ݮj�zRq^������}_PYe5[K����gMRz�`GZ�Jt��
�vK�O�]mL�U�;h�CuU��#���3^�G��;-Wa��95��DV

6�&���/'U]�;����sՅ����1�k��.�e�ɲ���4�!1��0K.cς� �`����
Vv���z�;�g^�w��c���ACAZk��Z��D~_�W�T���� �I���
5.��C1�:�O^4��.i.��(��^u�a��DeNd��_�]�Z�"��scۉ����Γ,�е�9�P8ý|$m�ܴ�F���6&1B4�L;Hw�Q�C�EU�t�c�ex��ǂn5�.a��͉��z`��#�J�=9B��V	���f�mvM|��� �|$��M����S����y��+t�ǣ�^���t;����#zbi�V��}�Z*W��C3��$E�k{b_%�Ϫ��Y���6�҇}u��}$���I�3������z��0-������q��'�T���
��z�m�S�I����]{��D����&�Dv�/|���'�az�j��s��5��FP��Y�8_��\���CD��л������Y����T&T�B�ʮaM@�L5=����Y³�R�Q��}c��!x�ͶPY��B��+�;V�λUό,*�li�s�DIui*B�QOm�!�u�fE���c�0mV���y"�����p��"��k^ռ��͋�2����r�R��i�n���Ļ���R��S�aE��L�~����=X��Eq�J�T�`�7*�]^[��VѦ/e�����h$�kS^:���U.�^D�٭��ҫo�,z��:�>>>>>>#ʧN�;�C�`�I��J>�	�&��Y+�t�O^+�ӳ�ۢ��J{I�(r�{٣��k�j��!�~�L9��C-��l���P�q�d]g<	�{�3��Q�M���޽[�l��,����咔}��F+���2���D}�~�p<��̉��M�}]�5\�Җ8��y�L݇���M6TӯoBiM��0�'���k#h��-H~;��S����t��ȭN1L�O�Ofs�9iq��Qak��W�XGp騆A8Eף<O�'� M�Y�4��n�-�2+((N(�Fr��9/maTsK7��N��ۿO@`��#�˶�˚J'`���n�f��4k�C�eȩ�	�R��Ǧ���`M��'L{�G�w��з_H0Ȯk�����A�
0",Ba� �-��'�vk�RX`�%�a�����<^���WU���5�,����9���H�o��b��d!U,���D��r����q=ֳ��Y����2�E���~#��F}����N�=C(��͘�����\@J%��Z� <c@��O
B�i/��s3�4��e+��z�T�4w�R��u�[9ؘ�P���g���2�ӽZs�TWm���{z ��슦B���3�Hݭ6�Z^�v��1
��ͽr���Xp2�gz^�V��͊U��.^i�˭��ݺ���Ej�!�1�fnw\߼��5w�ᙪ��Z��R��MN�]���n�l�]c���������0z���t�yזx#�@A���@{���(!O�@6o��pb��y������d[V� ܼ����\�s�5[6F]J�����3�C�f�݈�=�h��b�g`���wl�X½5	,_l�ʭ*�Į�z��3�g6jr_TP�m�#�\|�����4����;�ψjOC�x�-��pJK�ҟʅ�Z���WU��&!�^⾵e�/Q�V��͏��>��c6L��98~7[|��\����N��ƻ��:�[f���p�Qңy�@��ИcH��fh)��vI�[��3c�ح�|��3c���rӞ�`�MͲ�xn�gh"�N[]�ký4 �/���UL|��N�ʣ�Tr�Y�#;�C6qV����1�~�����PX����q-�C��0t�s�Oz;�&�W�uv��5Z�G!� A���K~��^/��.�-򷇯Z�c	H��e�9��}�^ i�,]Ph�Q� 'c�&��cG�F�My�:�0���2%���0��p�s�r^��+� *�"7�J1lZ�F���YR:�U����)
6'rM
UV�s�J�	�O��kfՇt��Y�r��X#�iQ���;���F�4+���2�풻�A�U��m2�y�aгvm��{����3��L������$~1�c�9�s^��7	�{���p�:O0�e��-�
��K���}���J�h��f!m���ݟ����L�܉(K�v�f�A�F/�����;q3�l����J9�9�K����[G;-�C/g(���M�@u�����sB���$~�OR����d��pH5Qt���K^HvՑ&�l��/-�C��(4"��,�S�h���"L��ZV��<�}���]m�-P��]Qɖ�3�ҡ9��Xp��E.�2/MoK�ɨ�������bq�|H��Ý��[	'-�t���ssОE=4�P��2�T���f${����KhrKbe<L��tb�sP%��ŴXw݈��O=�'Eϸ\Bj�2.޵\��P�O\e�܇;y'3�,�~��5���<T-�A���2�:�*Q��؂��J�"�Եʼ�cHOo,iW�JL��m�5s�:z��d��0;ҢS���a�;��eti����|��u;I�Cb-����9디K[\i5���f�2.s�� ��D%>8ϟ����~v�����)�2�	�G�@��s�hΔ�W�"z"D�Yy^�x�u�W��kb�[����$14��]���ʖ�v�I�{��c���<�YY� �M]V���k�Ok�930�wT��^�Lv��N��gx������`�8�ݩ�5k�ca�^X_�rzy��I�>�N�_��g���s�;Ӯ�+�[��\�Ѽ��f%f�sKG	^N�!��Lhf��/{ja�ױ̡���y<�sg(`�)�O$R̩̙��*�l?���~"F��0xl�D��Jh�>A ��<Pd&0�Q����T�o&mN�Y�}Q��Ч�vý�~w��8�"w}
�@��h�k�oJ>P1�PX���eE��[���1����R=��C+]���<�ු�G���Q-Xŗ�K'�>�A����v�`����{?=^U�C�M+����5�RD�!�hp�8Bb���=@���\[)"vi�&��0-Y�N:�Ǥ
`H|n�&���\q^�bfD{"LN	��)�*�m��k�0�H O:�T�Dc�^�?�񑜽K�=�0t��D����Cg����!�Y諉��<��d=�:8�5=Х�@f>�w"		�B��+���I� ֤��Z�9�\���� a�itqh�R��M�{	��`0& �V/8R�
��`)��@)���u�>˜���E��^�qm1��W�,��4�!��Ni� �]���#o���Ä�$"4���s꩚��e��&��c��&�݂֬SO�D>��>
��:/G�ID���ΝSpL�A
�b�Y=f�q^Sr��+bo:4I}���79���f�Km�+3pن����wՌ�� �o7�����d�%�$�I8r�>��c@tgO5����PQ�`g��0�"Q�v�՜��D�;f��c~�?Gj�}dLpO^�YR]X�F8c�1P�3y� �a���q��^F�
.�Y�����j	����~d9���^t&41*��0�;qluE�ȫ�3:[ٍ��;Mԫ���S� [���%���7`���&T()@�,b��7��up	�1_V��5ݬ��ժn/��]����}e�&�*}nY��۲�1�pY!�$���L�����oN�#�Y�t�ǆ�wf�K�\3���&!��q�o��"�g��a��E�,v5:���V��+�3�ԃ18��qE4�����۸nx��qm_�.z�M�`GWJa#'n�,�(ԛ4Iw<�<�=s��,[Ը�0L��"�~��w�Ms�e�7�y�	j:8�/�T��v���,�8�ZK��p-?O1������Hc�GMt(��@ ��DFsn���&3�_P�LP�	�E�)�~�N3q�Z�9/LUO��Rܝjp���؁���ν��*��lӆ.�Ú0��
�*�o\V�R+>�C�y�Y�B�˨�й��A��[���-�Ꮭ�$�J����	��oA�MC.vK�8�Y��A��;{BI�wq��f�4�o!�wJIfY�����Իży�
¨������;�h�7�}��:CX�ɈUw)� ��,���½��;��!5�2;��w&��q�i�o�9��`��_�j�]a��ݔ4,�C;����>!��[�#'�����l������s�%�܁��)��m�ޓ��<�5|��w�X��+��L~�Fϼw�A�jB�a��dl�`�qM�gaU��Z�v��۷�u��1�D1��ۯ�ݓ��0&P�.$E�O6����.�4>Ys��2�<��4e������B�x�p)�^�礯=^_*W�E[	�t�9�2_���0�ip�='o�JU�,2���/[&��өq^���lyCٟ�k����wW\#1�ʳE�)�Y)�46?q��K]�v)�[�!#	�{n42c�3xBk��BeBҡI�u�1׹��f�"�R�/v��"O�Ƙ3�e���� #*|CT����Cz7ԡg��`�fh\�f�`>��k+"���Ս椐�����ݏ�1�_�8�d�F�C�$����(a�oD-r��8i���0�;,��6��S"��7GEs�
�?�i
�|����.xy�T�~�.�P�� ��^��Q.�'0�>2�yݡ�9��3;cr&Ҝ�Q�)v֨�QZ��(w�h_q�#
Ɉr���ob,��$�}�8(�$��F�Mz�#ā�L����j�W�&>�]�٫��ܘ55�S����:�4V�������$:ꤗ�ubѫ��uó�����c=�w̬�����WǙ�7\a~�R���<SY�8�[����k�ȊiV��_ ���uqP�v�죽���o��}q�q�o��[C��S���-?2NX����,!��`>�hܤӦ�ZLI�� ��I}$3�N��N���	�0��{����EQ��j5�PJ�sס0�mj/n�{�tZY��Z=݅����AP\F~������g�X�-g_�`�R��lA1QW(��v��T�ڊl� ����ŰRa��!�'�X4wB�/�?$ˆJ:�9���X=:��\�N7��eL��R������o�w�Wz+�+�?�Q~�F�h�P5�>T"3��Љ��kj,���x�ZX"��j#
B{�j����~��������Xh�N��x��~��3��,Κ�v��ԿW���e�ٛ�{�@2;�~:.ߵ*k�2�D��ame�HgT	�إ�M��)z�dY�l���홦j���Ac���C�����X���̜��]���I�N�X�il�a`{�6>s���L��yH��!�6��}؄G��6c�s��[s�F9����e�0Rμ����G��^գ��i�N��N�/��H������UH�$��YyD��HH����e��#0���i"�18�n$�w
emx0���Ú���Mコ][�Ʈ���k���u�j��!��Yrj2��mnV�������O�X���r��y��-��w{(�Lh�q�P밭�su��urَ����2�J�G�vǺ,n�i=�j��^j����7j�ɺ��wJl�����}I�En#U����x����m�6�J��9���9�j�����n��-v�t��o�g��� �.#�dZF͊�ElԞ�@ϖ�ѽ 8ӧ��2�X;�V��Uzv'.�f��!(�����Z�+wmJ�n�x3�j��N���`��[O
ӯ���1nޘ�!+��n����h�V�|v�,�9e��"ƫ���K��Z\k��]�.�ત�J�)�w��w4�n��]n��wv��_��U#�o�KGk��γ�Ӣ�>}kAj1v8L�1���԰���)1�Y4u1�-TE$��5�0$�V��J��r4�+9d�1!�\D�8�5��]��|/.t����,mU#:�<�����M=v)\���yά�m��gy��U���u�����I^�Nb3$*�oQյQc�V�d�lm��>������������a<r�i�Oڕ"��Ϛ��1#����2*�T�Li��P�qQ�� ]iM������e��M����\H�E�F��@� ��G3h�����ڌ��L��������I�s0Du�ͪ�9�����úev]�T	-��n����"1�Rv�W�ZQ�%Js��s8*w]��2��l���u�;�Vf�ʸ���əkir�ࡻ�ظ��8�G���2���V�|�K�;�v�&V��X/o*�8�[`�ZlF-�"�Q6���b8�H�kL������v�ͬ�yQ�:�R�XUKړ���qN�m��-Eobt��/���b�%�n�D��eV��7�(D3����C��8�qk��]N��f_��XRa�(�8Z�zg�2��.R�BK�QŞ-,ލ_u���yѫ��C��a����{���R��륶��"��j���Wf�N��֋�Z!���P��1:��K	��MC(�n���!R1��:NN#+V�x�S/������"�xV9Ǒ*�B�2�N�-�u�"(S���L��\Oo1�m��	��`&�zq�vM��:�gJ���p7�*MXm���`�̩�R�S3�\V�D(y^��ӅR�m�k��Z2������
�j2���L�"t�0�2��'���e�K5-�,9��/Cע�K�^��,�иoE�al�fj�N�[���/s{j�C��I�.������w�^����6�I�bD�$IdY�4����q��n<x��Ǯ	 ������h���U;7n�7��{��x��׏<x���H��H$�k箵x5�V~�r�Ʒ�4���qǏ;z��Ǐ�bdKPEk���Θ�TV)�=tێ8�Ǐ�x��ǮE#E͵͌[��Ǎb����o�+\�Qgup��ѓTk�r���~6捱���*,m�c}:_[�z���65���S�hذR&,�*.lk\-�I��ۖ���_K�F�K\�9�*�p�*�"=�<�B#�=�2u��Ý�j��pfu�-x٦�I"�Zw	FcbŽ.����-�W�̇L��c[t.�{�p���c�07�7���B����b�hB�� 2�z!G��,����!5i�1����T���m%�����y�f8b�gu��y/^�wd���ޚ`�	u�6�cOw;�ʉ<�;�6Sp9�D��o<6@�4���i�r��)(��(|���������)��Č{�=���� B��Ad^�"K��R)�i5���U7c�:���@1miL5D�o]v���Vڹ��(/C��"��t�I�;�RO��&*ۤR���mt9��P��x��R��B̖h��e���f��y��zz�/��-��M�ј�?�H����M�E��6"Y�OP,�H�vo[!خ���3���Ӭ$ �(3�_B4�ڟ&w/g�To�����õ�[�{A�+�7�V1�S�p����"��D}�f�$��l�=�a���g>��Ɓ��&~[J����lR�RvH�M�ߔ����Uj���0��?�wf.��6:��]�W�{�󡺄�0t��:;��:�A�JۯG�
�W�
Ё\��gE/�r�Տm!*��3F&]�b�~����I��\�Mչ��h{n��j��z��fgnk1|�>Ěu_O����j���q�P�謝[Ɍ�a���״�Ln����d��շ����Վ������^�ߧ2�[�ҳ*�d���SLcÜcq�Yޣm���:���V'6�@8��Ð���ܴ�F��� fD�I�.�W��R]j0��3�
t���R�i��Af�t!�0t�t�$u�[0^\TE�m�hp��0�Tj�mܖѡ�����\X4	i��<וL�X6=WFD�ץ'o� �r��T�w��n?J����9k�~�w�^��0(_	dH�,���N}T���r���^p��Q�n�~�0Yܒ�I� `/i��ȟ8~���.b�����"�#�D����}9?F�}f��M� ����QX�@�c���s{��S%�]j',A��動�ܯ�ق~�t?4k�kO�!V�3���J�+��"�n��B>�Eh��s�o~���|�<�ʐ�cy��h�P�3��黟z"S�	*�^�}l��.������斉�fw���l]�����֍����E�q*X< �O�����T���>.������k�x�C�ջRT�0g>�]4\
�i�8�c9a�~���h�5h&�=��`
�
����I����k�[W��g�Q�9J�9<c�ڡ��pZ��,h�7zVN
�@Ƙ6
s������ؠ��E�"�J�	�d��,Ӛ_�-���fhHK���`�oN�*Ci�53N֚M�b��Z�	i��A��<*�TD�`���������?1����ݢ�f�Ge�I:`��a��;���Q���Ě���_F�@jvki8Ə'!�<1n�2'�����=19��Ѣ�k�0���xk9r��*3����a)��u{"1�f�`�bh�3;��**���8��t�f	gy*,ֺg�{�ԫ�8�^�i������} ���
��ȓ��Q�����GW�*a ��h�3��q�Z�⠗�R��B۝j�~,13��j�Ո�N�(G�C#���L�S�q��P�z&ߍ��&�4���ܺ��v���9�Ύ�)���Χ�3>��D��ba���vk�R{�9��M,�p�蜞ї�y3Qu��
����ˮ`�Ո>�	�b�j~VE0)�g��섋��\b���J�硻5kGl/�@ �h{��*��ĸ�Ts��ABM�H�Py������8q�|���}'��g�ΣY_0�hq�����%q!_OZ��Z�htv���R�0?�TK���۬����.4+�
�oU�,���[��2��4�L�Z�����Rt` �T��ַ�5Ǝ}s4�Ub�![Ԃ����dw!j��1+�Щ�OS9/��L���[�/������'���/^<}��c�ʾ3o9тJ뽺�I$d+	����M���]��;{i�t�uVB`����w��I�h����c�z������������õ�kڣ]�:����-ًا`iN|���G2�iP��%vP���Y}v�Ps��������o����i.%�b<1��H�u�`E��JusMPۜܐ��sN�w]�j����?w#�ߦ���1Ѕ=��amI�|������t�1�]�7T&�[��5�y�F����[��nOau�m�FS�(��=��z��q ���P]J��I���~�K���}�C�3���1E��Qu͞�cڍCc��3׷zgLG��tʡʭj�x7!Qߚ~T~*�D��}14�l�ޗ�qiAcK���Rq-�ݦEnX�N�~|���}�!��,ץ	�^���@T��z��Ñj5�PIz�/s���`���tAC�7�w@N�x�~��x��Ȟ�~U4���~A/F��VB����`� �r/�1.������l�j�n�C��GVH'�����7�	���0M������6��Ki�gpM:�[��4݋���2���Tp �ȑ�A��^�����O��|�Zs�B#�f<Z��X�����-^[i�f~�rf�s
�F�]]��RE49�%����S'Vj���$��^n�Z��lx
�Y�4�I-��f����D;p�:êMUD�dw������&kE�ܯ���:�Ѻ6���w��s�*��c�g�{��|���"��پ��������=- wt;��;C�Ǩ$oK�x�����&[�j#4�;<��݈���?�Hj�}V�@͂^����l/�n=Cb.����bw0X�.�c���fk!b��q}
�u����Rͮ!�}�����N����L]c굛Y{X�㈵X���Ά�0�gd9Žŗ;������Yj���NS�+���ݡ6�]*&�: �����s�l��"��Ëh��%�EǦB�`N{'ˈ�����(�d(�d�]t𕼠4������o1�|���n��(���Kw��@M�J��^,�/����dE�qCz%�{ �4���Ъ�;o�|�ΞE=�DO�	�~�� f+t��g�Ō2\P^��y1	�{%Մ�S �I���#�.s�,m��U��U���Wo3�{I��:�L8�Tk#r{=0;�έ�1	�V��)Ɩ�52O���k�fM3�ذ9��k����B�0�
��C^}����f/=ja�~d^��O��9����D�����>�H~ta`֓�q�9:3��%��������I��"���|	�˚�8�~�2"e�t���Ĝو�ǌ�OT�v�KK�v۠��d\��l����oYיq
'4��I_#�N9��0O~��� ��ouv_>;v�q����J��S!��Z@�!�zDD2ס=�@^�}�.�qxPE��C���g
�#5;g��gBO^O��ük�;���\�ɺ{����FY��$������ov�����ȶ����Z��(�'>C�Z. Y �#��f��> �VHkw6h�;�Ó��6��Ee4��������*���n�C�8���+��0l��G֭�h��V��ۓ���3�㭏M0�D�&��u9Z����ɍ+=Ok��f�}�{�M2�H����H��q�\��Vj�\����/K��lw���_��}��~����+#S���,f�2sw�nJwil�ZG��ț��Ʀl�˙��5����g�j���L,����@K_z�	��?^��+
\�ME?��[Ŕ&����9�4�TW��A�RY(5FCM��*�Ξy��=`���D{��
Χ��F�t�����>E �����i��������͸�y�;�����	�)�n���
S>��a�l�.�k1a�FZ�6.@X���Ӛ[<g;v�B�7�0Q@ͫ��Y�;/�P�%��u-Lܜ�����g��D0o ���<����n5��wuB�Q[t��7�wu�#��/4ND�C�)fȍ˭�m��V��3~axr�tB�5zx�~��� >"N���1��[����^��D���V�'�HEU!�@���G6p8�70D�[�΂ƭ*�Us
j=��C�-���ݳ�LK.�<΅�M�^������ T��t�Ͻ)Մ��y0�Jܪ��T+0p���n�kz��"T[B��>�����9r�X�!����o�G�d�c��Bn�gO���b�n�u���L����;�ݼ0�p�{m�:O���z`�m�CD�EBu��Mjn�������:�M��3�O���=f�mu��3߂��MW���h��b$�n�꫽��4�!x�v��P�'����^�PX��P�Sø����6�:mr��ot&6�7�V���hSW:Y�>?�N�������لz�O1���k�/��6��z@��`����KL�Uc�
�X�O>�>k`��ƀ��f�~�.+�J�)�ze/�ۉ֪nzB=����X�K ��D?�A0O���'�xA�F�ϡ����9�jĤh���c��P%a���[;3�O/�����lW��6��n	����e��9�e��-�ˈ��;T0��ګ�>˥%�������ܘ�y�U�i�l�2����t>ܓ\H�V��4T�C�xsv��!����X�u͛)��z�Fi֫��8ڼf�S�M����өE�Z���b\�vS$��')�\ݘ)ȓ���$w�����{������[A,��gC2ǠLDS��w�ZK�/.�c�5��.����=�l.������[�3;��$-.(2z�!�8�ϧ��8Z�׊xn��́q�˃T��n~n*ی|���D��Q��8f}N{袯c��J�!^�k�o���~��a��Q�l6���&���ޜ���E�-�P'�T���C,��ZUtP������l+`c�В���Y�~Ű��g����:m�9��dz�oCJk���A2�J�'6f�9J�a�{��y6En�{�9�G�K?%�2;��W��j��w	-�q�t��O��3h�X;h�;��m�bd3�,��/���&�&�/ɳuW+���kb0��~X���e��A�w�U�(�1G&:4v���@o��%�{]ƼQ���ר��̘����x�Ba���z{`�qfZ���7*��OY���I���E�{�)�b�F�D@�T�u[���Ͼ�w�
bW�|Z�w���7�'g)C��@���W��g�s`J-�.��Iıv�:Y�]��u~���oUBT����x�&b�q�R�'C�s���Q�t�L,��}[/!�S���3�*�y���P��ocдS�i�CC�S�U��.���'��N��o!�C�W�Ãs��k����5�.�s���>>>o}��8�9�Ȼ�7���h���֘����<Ú��л╩{��K1��w7���7��.�uq���fJ=.��ѐ�r�B9��=p�_��تd\}t��O��N�c����5,�m~ȕ�tc�1����׾(��~/~�L6�i��v�5��S+�7B�n(�ߕY0����EI���3���P�8"a�T"%BxO�;���l��))j\©}��4����S�0���wѯǧ�h�#�^��%+c�3����>&���0�p;�[H��\�Be�]�/�v�Cd_U���t_}Š���с��FL��ߢ�0~���<���`/|��
!��c;sr|�oF�|⮺��͚���G ����e*��,;y��ؠ�OB���O��&Ė��0!�-9���z�֥B�d�G����?+��d�i^�Y:Φy�w��څ�F�1�0oN8S�X�j���;hj�_Iz;!7H1d-D�K��i��p+��V�^���7�F����2/cӟ}*T|���VfQn�-n�f�]��k!����L�[Q��fv�e�B�������&����ܽ�[����(l�*.V�ǔ/�{� H���I�oh�n�b����:��sQM;n�K�"q�n�r�$�J�����/k��_Ia�So��Ȧpw�3�G�h��Ɓ�����3����w�߷�#�8o5�%�{N�'�3%&D�Q����l����A���ArL��5�b�ݸ�0�@���p�Pq��Ľ����ґLk��I��X�l�]�P�)�/�0cۑ��?;�ޏ˴p �+��qȼ��� ɢ�7��:�Q��t8�w_�ZO��N���"�S�9��r�&���q�8u��b�48��g�G�1�r!6���>�%�iL4�ߙ%��r��n]=&33ˁ��3۞CqM9�6�0����԰���H�8��D,4�ګӜ�-���
��
����зI��l�e@��u�bA��A:W~L����H���e�N�=c'aY+trчY�+��X\J�[�4ڐ��z�o�B���oRX�?��6̈�~�FKn���9@>o0u��c��t�7���7so���-�1���	r� �mΥ�ݲwă��:OU��-��a��zp�n���gЙx�3��#�}�/���}=C�?Y�j0���}�]�&�Pm �D����%�&��Mjx��Y�KI���%_��7Q�����]��3�A�To]g];�l�����U��'
�A"�*ݚ�Fb�ĭT�JW��!�7zȖuJ�խ@�S[J*��y�m#lf���q�Z��xcJ�;~�ֽe՘s���S��C�4��[^dJ/*Ε*��h��1b#*4�F<H�jɋ7%ʈY�b*K�ǮkHV�W�1�j=Uב���o��6�E���jݞ�.��Ǩ57�v/	~��[3q�(L�҉~S��Y�\���xn��Ӭ�q���3�H�'1Uic[vs�K���:!{�j���*��w6�5m����3`7���[��#�C����wF����y	�1,��&%�ɸE3w�i֬�%�G[zdݬN�,e�h�D�ݗ5���c���ܢy�:Q��AnZgv�-i���+��o'`�jN�����֯2V&lÛ�J�r�v�^m-�4*�ۜɥ��N�s={F��3�c|�s��Wg��/v�ưv�zB�r�]کKz�D^��;y�V�\&WY�TDu�JrJ9��
��;��i䴬�,��5����MK�CӤaa3>Y�F�t[�U��z��"�e��b���>�(��j�͗�.�Ҽ�]�dmfϡk+�egĪIA�ȬP�cU��{�(�g�\wxL��Đ��g\v-�b�\S����鶍����.�AJ�Q�eu"M"s���Sr��j���6RV��\�%�X�\'H]��az�u�CF�uѵebfԒ����nn�Ъ9c�;�E)%-���F���[:*�֙wly~ۤ�j�	'a�N�l�5%��t֘���a%���Ӛz�٩2�c�E�U���l��gY������3XN���N�q�Em��n%\�jFH�Z�'p�.���uװ��k��]ڃj��U�Zbf[؂��mn]�FU$]"�m�n���^K�v�^ն�k��j��Q��1nė.���ZL$ns^�������5+յ�K4��y�
�7�)���Y�-0�����r�mE�!2�v\5:݊qgEf�B#n�%q��'�=N��gsJX�+*�ݍĝ�u���fK+ax�K���kԵ�8�9�TBѭ�8�F�;��J��TS�K�]1�v���%�u[�f�7��4�pB�2v*¦e�R.���c�������9^��\i�ʳAd��"�<w'�N�x�]W��VcY����\w�S�+zUT3�w��2�������%샐�Fv�;g؄岄�Wk����s�^�Nv�JW+���u]�S
���)��"�qu�:R�1]��0��R�����n��uW��)�4��
<j��f�U�mc%F�xݧU�w�J5�{l��Z�ڬR�Q�V��]�9U�W!t4�;2gܒ��W�گo9[�4Jĭ(�n:��j��82m�P?KL
�RO2S@�A�^$������}�{�57�N: ;��"ȗ�V�9&�`��ݿ7��}�Ǐ<x����Ǐ\C�:���P�}��o�M�**6��U1��6��x�㷯<x��Y;-�����͹�HH��I Sz��8�Ǐ�x��Ǯ&A;@�ȴ@�h����cS����Kż�q�����q�<x��Ǐ=qs�5�C[�\�A�k��Kǈۑk�W�l��]��#'.mt���b�6�o��yعQDR;�V6ܥM�U�)��E��\�nW*"#c������x�����F����[����m��Yg��HD�&��.&�A%� f#pB��� �Pl�Q��L�73**�sC�������a�;�v�jT5�W��Ox��eḾ�{�����ɰ�-V)�eK�I$Q�C$�G�'@�R��`e@}񍒓-3�����T����%�]Be�TB�J0�O/~����^^@///-���R���*ز&���;��������'��z�����+�W��,�i�����~�t�� ќ���R�j�� ���JbE�c5��G;�ٜ;��].�3��0e0(�ݣ^��Ѳ�sΎ��K_�K��YȫU��*��jU�,�����u��|�XSBS��n���U��ml�-���3*�t#yPO���=D�c��j�s#3���󚇥3kD0#s�+O���u���c��S�}M��&�U@�f��J�l�f�e�=̈́�n9�m���Jpq*����zү��_�>�h��������%���e���-�J�!E�#�l���s>mGH�vN��Qx7�+Pm�#��v@j�9����ן7�7��0�]���]88��fB��O��o���~�9�-��M(m�\({v��a\�"�{��]��a�d�U^���J%n����*+��7
��G���澷4�Ez��Xf�D�R�6�vc�-E�kmPkSYvtnԜ�c��ׄ����m�5�0F����jUm�p&���n��� u亮b��L�;��I�U�IX�	�:�E�؇Li�+���z".�����W����$�<|||||}}]n�7�18y�~L��.��5]˕Z�0�wM�{���חi~�b����ba^����Ra^��9�}f{ʄR4����IOv�GxkM��>n��(K�a$&g�g��������;�����w���ݙ*C�Q�DU��҇q*t���H�cz/����4+g����J���W�v���㶻I�����S�I��.;�kpv���i�QjY���&�wY4��֞�-Pr� �	U���2I"Gc�[ձ/��1�ɷ��陁�W6o��A��J�M��-.����Nnw9�e�E��ÐRr<�	���)��S��zVo���#&�����a���~뇧���L~�����/�xt�|Ͼ�e�Ϡ=�O֔�^�UY�%9Ǆ��Y���` �i}��KZ{Y)g�^֟X�N��l��
a���E�U�k�<gH�ۗ����ё���"Ws6��au�J����m�Tc�u�smU�bէS�k3#RW�T@p	��(xnWc,������*�c��ކ1��#',���mQ��Eȫv����2�5�^9���ڙ;�
x�����珏������+����u��be�"&�C��4�U�E7��!�˸�e���#�<��qЍ�"iÉ��3Oww�.�T-:9�g��x������E�:�����ي���sb�g�J wgZ{���_*EX�>����tk��q�ѥ�z.��P���]v�O�w��q瑦��"d./�6-��4�+{��H��o���}�W�F܈��P��z�PSx��Y�Ni5/��3s�NOu���5��v�RT������yC\]����ۤ��k,������߄p�͎@�uE^�*�����7�G?���y��FhoG��q��q%�KrOzN��M��S��z�t��ͣ��K" FP��g���䯹f���}Xy��7v؟c���8��pH��:��0���)arh`�"i<TYSb�k���L�ů�t��2y�q��2�EKH�u�NT���|�8��Kee�O�P���op�h��b+:.n'�b��<<g)U�!E截��A;���Ś{Z�,qߝq$,�SQo�ʻ�{��t�����Ī��g!z�	�RZo�y��|wbZ�M���珏�����eӾ��n�C	���;�z"���>������j6Dk4�'%���(}=���]����o<�����!
�n::�}Aj[�*�R}O�/Z�k+`���Nu%^H�f�˦S���@7�B<���i��?�y.0�i���u��I
�u��Ҏ�v�x�d��z�M�2�?\���-+����'sŷ"��1�UC:I�IJ���|r��:�ԭ�a9AO-,��sj"�f�;��&�숵�" �����mh�D�4QTt�<�KC��Vw| ����u̽�܋��y�f���w9��$}�D��>I�ԇ屒��J��k�����E�R1�낸Bَ��Rz����i7��(?l���}�Es5VL.��ӝ��ϼ��y�k�4�Cx��b�;�I8��{�/��u����\�2O=⻥v<0���k���@u�D��zb?ǂ����d���m��6�K|u�r��]��"!"�x�t�֯��h)��VeM�e�x�]LWw۞�}Į���v*�r�aX��l���3i�3p�[���o��{���[�{P��ǻsqH������]3m�m����v�o��$�~�������뷟g�9���cs���dM �ܥSU-?�O!��\��0T�v:Q���Ϟo��1���.�Ǫ�Ӣ�ޤ�lm__�/�C_��������F?9�����e^�����ʼޱ>)�w�7��]���Nݴ����'����-yS5]�9��3!��K�@���gTk�JU����뇀�ޭ�R.�q���Ͱ����C-��@3���;,�: `��H�(�+�ae�`��f��jM,P���U�p�#�nYK=��440�b�v��✋�LY���ςI	��?��_,���V������T�:Y�`�܇���E���;B�lN�\ ��uQܮ�p�[ի���]�B���}Q��65�wu���X�T��!�GH��T�d�3{ǩO��2��R��Q�ftf����Nm�.ȩ��Db��}�7�R/���l]�9�)����0�W4x$n��|�zE�9���L���޲�c�	�׹k��c�t<1��C����ɶuN!V�=Y{C��c�Ue3E���m�Լ�8��՜�3��jGM;������t�#t�t���S�U���;P��ޏG���� ^�7���S�	����=#r�Ϻ�$Xt�����
������fro��r����M�-$ozJS��co�T�Fbn�1UPգFډ�W��s��p^���нX��z�R*���.m���@"ׯ�Ơ;$�>��x��4�עǀ��oK����>�*���(��N�U���V��@��QNױq����*D%]�{��;�	V�y� ���z�����`��t��?�a���#�O�<_Ԩ=qoi�{��z�O7nd��a,re�]ϑ����/\D��Y��?�ހ��8U{�ޥ�i8m���4��h�����9ùL��;uy��}�h}�4���4c���H�e�V�>c0����S�A ̀K��'�M���@�#E��>��EFΜVӺK�n��>\s�sqz���I#�6x�ח�h;���X��}�C���7�U�m'�(�mbԍ�NM��Մ�̇{;��N��	S%S�z���Ӌ��p[�N�Z޲�6�m��˧�$Pk$�ۅUu˭T����bj���,1ߎ�*jRȈ5��K:�w�6%kno�Ua�M's��b��=P����o7����d#�:�X:=�2s~5*���g�����>�祦���cyw��f�啎��i�dǞ�=F��&V�����Q��[�t���R��W����"��E�Y�ce��������,J�q���B*���m֙��=��g��%����no�un�x�7&�<x�RC��^�*r�+6�ZJc�o"�}n�ǉ�$GRYv�w��~�g��#�]�6��D�F-��� ��ޓԨ�炩l�<Uy��\��nx	:�-�SѾ�;���F3��"�\����N_a�����X��6��N	���V�na}�>�-5��y�p�}[]P�v'�U�yޥ��%��aK�bïuv�\�f���Jo��ǚ��H�w*c�f�<���g��P�3��,#�L���t��q�^��a}�ޯP��"!"�m��WѨ��?-�&�5N�ϕec�	��9���E�f1�EGP�.Õm)�ڭ
����6��j��1�ᔹT���[�twj;;j�ehՃ�K���{��|2��D �2IsL8�E�svd��j7��8���9*��A���{���:�"l�7����y�9���;p=���#�����rj(U'«(]�����8�q�yޯ"K����=�NpM_E�olKn�o)�{|9e;���R�>�~��#�/L|�7D@�'��t�ϣp��nӀ�������) k���>U%N���S�BRy7��j�:���7;=��[E�� �k����YY�Z'�Z���{�:A����qK�Uɸ�����㶻e���[u�O>L���Fqj�e=�S�>��![��p�=많�.�H2��+�İ46F͎E拾�[ـ�6�$q�6��2��q@�Gc8gO!���i^秗����9Ga�n��O���{J
iO����hL{2}sNdVy�V�wa�u�m���t�D�ԥgoX���!�4�Z�.�*�U��m�aɲ��K��=3������#�/�(�f�����׎D����my���-P*eHm�T�}{��;)(z����?in���=�����՘m�X�C�a�&[��g\�8���*l݉Q�z���e��kwn�'9��f(<J��Xչ�a���hªӤ�$\�`�ޗ�L�g\���l���Qw�q��q{����������ޑ��UV|8LZZ�;Υ�e��6k���==3�m=�N u�t�?%||����|��>�Nt6��
�a����W��-���+����vNbu?��u�������sQ�C6�z�'�Y���g�ᔃ�`a����Y��`pm�x�$a޻#�&k�^k�1Ew.����mpo��,-`�ҕP��ٵ1y�;Rz{Y�3�����S~tl��I
[�i�����>����C:��>���3Dƾv1��/P�f�-7qFT��;Mڲ��w\�9Xp�7Lb/���U�U���a�ϘW����?�pߦ�"�.�1�4H�P��Z��w���y�5}1�GHe�^x����B�~)�;>ܮ��ϲ�R�Ȋ:�]�HǺ�w�P��>��4�Q#��^#{=u%`���t�R�}�n�1̷r^�ky+H�@�Z<V_sӜ��?��(������gV"���>t�T���ஜϹaۈQo�畘��/"�i��C��k�9���AA��0J�|�v�{�� "ؒi �G��U��,m�xSɹ��x�#N?+��	���}�]4f؍ɓF��-�n&Mɪ�qٽ�[�K47�x����|}�U���ǉ�:XZ�����wg8Y	p��R4��e���B�gz�Á�N�R2�Ne�:��y����zw���gg2'j3S��lew	����p۳�?�V����F<�0#7����q<)9�9�'dݞ��׋��뷻]4�&��.��BQY��Y���^"I�v"���:��`)9�dy���jgXey�WV@�n��VIs�4$��4����/���{��I��F��ާy�e�7����>�65����uz�ut�ei;�Fp4f��`c�:F�z�I��J����סq����3�r�R���E�O�r��f�nP�$GtQ��U�_yE�#a+��T4���{^��6ZN�yص{rC���^��W�G���r�]�+ʷf�ܾ?dt��a酧d�:�=��9/|���wgfv��oH���/T�������z�g+=����^dH��9|��D�+�ARx0+/o��b����v��oi��>�=ӋjY,��_%2�4jeU܋O�����Z�%7F�[׭�]$��+`s��]�W+vS�V��JwZՈj��'/Iy�(Ȓ��L��Pd֡ev+D�D�~k7f4f��T�DKĄ�q�Ջe�Ax�B��XUP��3^aں!�+N_WZ�4jaɳ}6�v�e��*P񱏰��n�7v#��j�#|��7�b�zR�9
)K	�5��R]�3�:):o�m��`j�ayr��q���7J��
�4Z͂�I�!%����)����6($��=ۯ�\���գ��n�����<u8�L�2�ܚD�' ��.��#;+A� �7��H�B_M��%Wz����<Ԥ�"s�s�u"��r.r�4Q��X��]܅I�ލ�Қ�Mf� �ɱ�".e[v~n��#����]��δIFW�詢g,6��H��ﲭy����ܷ�{&<.�wN�}ë0��܅�Ks����dM�y�/�#g-�ٸ���8f�H�A+��{E�$��d�q\�!�<k�����q�TiP�ED-�ޣ�Q�`+2�jR�����4G%�nʗ˅�h<]OEvm%�C굍�^vP���/G]�F Vp;�z�<�NcU�j����vs.S��xp�˪��ŷa�N�5fU�:I�������Di�qZ�YGH�ȷm�:��-@^��e9��p)"@�"�*l,��˨0ꫪ; �jn]���a%p�N���V�`��}�h�5{�8֨r!P��A��ҥn|��s��!�ɕ�[h������)0J��[��u���Ou����[�3��}��J�R6c&����#xX��7z޸�.8��.t]�3M,�zi��U�]ug+ ��n_X1{����j�H��x�B�mJ]�V#��u�v�E�vuu�������靌�۲��}ɎL��uݽ05s�$�r�:�ݻ�����]���5�3"ؚ״����=9ǰ�`���o
��wz�G��,��Wٰ�*q���
j��M��Z�n�5���v\�WŌ#ٍ��;9M�=-���e=�k.h����nv�A�gL<;�+�,@w��Y%q��_Q�Vf��
lS�y-����2�a�\ڻl[�sn��نO��ДMY���6�80���n�����n�.ξ�"�L{/�E�!=s�2A*�,�"ءN�	y0t�s�m�y!�1���WLȖ�'bV%Y�v�xl�Ğ��Q�4�I�2_%0����bhw�+���&�e�0e�7�.C$��/M�N�C\�݄�[t��T��V96h:�q�/e�ҩ�����[mF�y�Np��E��M5G�tܕn�_okҲLj� ��GQ~z|4�	D|H (��ԑJ��RH�� �:v�ׯ^�x��׏<z���bTHB��CZ�FE�UET	�B�CLi���q�<x��׏=s�	ڨ�������w'wg.n9�H�%PSO^���x���o^<x���>wb�r�\�~qxܽu��PBUFI1����q�<x���7��߻���IE�PX��������"�'׻�W�Ss��5EL��Wu��p�����%�+�v	/�u_�r����co:�3���!�pG77-���1��yݛ�"	ݹ0�g+���I�Ŋ&19:�b���M\�T�D�H��Nb�$�<H �>$�^����9��ҚxYѕ�W�%{���d�������Ǵ�6�N66*�U�eڔ�e0��u;,/w����z=�H��*�� �s��狭�^A�|2#��U�ح^�z�8 NW̰�敮�op'[~��~�v`�h@C�H��ߪ�sV�.�{S�������[��X_��7��2-������wLv�Ӭ�^���]藿)OyX�	�v�~�ߩp����Xf:�ju1���cmGt���vvwP���-�z��dD��]���D֘]9���A|+~��̎�QK��u��U<�P(��MU=!�cҽ-���8�}���W�+��]�Pb/-H���i��<��1���ih�kTܰZ�f9�pfQv9�#r�^��g�J��u�ul���r��/=Ү��Y���7�&{oG�h�3�	PJT!T��G��dk�p��s{4�fn����9��0^wDO( �ϑ9�x*��1ˊ�kxڏ��m��u�$R���bU����ȖV���a� ��]�Q�fbYT���3�VKb,�튯V�f��}�G����:w��$FR�JSз2)l\M>�'���H��<��m��4��:�T�l6�]#��t#�;�k=��������{�1 ���p�]���r�S�l�W�T���&mnڶ�{nk�S��P���GfAd��}#���ϣX�:��>S~	���Y�":'w7��N�m��l�b���:�+�0Y�l;���u}��pF}Z9XIU|�αL|���OM�wdk��i�q�J`�������1�;��*�v�U���z����@q+@���8��.l��e-���G*��+o'gS7i�-84�ɗ����r���yzW\!�4��Y:���63����qB�#��{>��?r���ߑ��}��GT���I�3��2�a����ÐG(x6hE�>�m筮��稖-�DE	���<�FoFp���|�d3��G�~)W���&�/+�Ӷ��XZ�N�M��p~�t��$�o���<��K���>L
��F��ڧ���ܬ�ҍ�}���E3o���WqE̎�vb�&Nqu]�����ìېS�/x'��ɺ�7F���t�������u�ٱ��/odI�M*
u�k�un^)�w�n�;�Z�Eckq�љ�1��9��!�mo��������k�{�g��e��aTn9�*���&eA���{��A�6�$q�ٶ�]2�i�f')�k��b��9|Ӳ�լݯl՟TP���>�$�=�Օnf��n���M[Y���م�!�xU�p��MQ���JbY���x��Hm�0����3����3�P�z�@�Nja��G#�ϫ�Oh��
��6���j�1�����d��}��� �:P�pS����wJ>Mr��Z��&���:o�������O;�σf<�tY��p�t�)�f^��>U��y=Ӂcf+�\�r��k[0vJ���n�3��GN����L��wغ���Y����؝8�rF(ܻ |.϶מ��t�4��O;��l����L}����;�D�_�����t�E��@o"��EKHfl��o���n�2C3j\o����#����mхb�\iqگx�U��O�zs5sh���+�:
N��Q���{��ZEL��Fo6nt�%El9�~�(��MY;4��O�9�\ɽ��\�����__�S#Q��y>��UTgBܖ��ԲuRt�4̙CJg$�^Ui�*W[�SUgE\�./js�`[ս���߼||||||�&�����{*�1��y{���G}dQ���	/���
���
��Z�u=#xW�����He!��Ǡ'gU�"=�+�\_v!3AI��:�-����z��7��������C�w��;��Sղqj����&�sH�9u�}���38g�;��" ӭ���v:*��3��f:��w�-6g[�BO�N�� y�4{�(�Hͥ#:�n��M���9"ݶ�٬�H��pH�^�U�B_�I}�U�c�y��Z��ё�ϙ*�w��8��)ۄ�Sϵ���Gz�X�]��ߎ ׌��)����sj~�:�sZw�Ȣ �=���u[յ3�A�d%���z�1������Fw9���Ἅj	㺒I��-nTx�V��!{oa[���(��/SY��Ww��)����65�)Xn�%q~j�3���۞~���lȳ�=!�ˆo�#�n��&DnԞCo�$�����c^���L%3��ZK/'!T�"4i��E-��ٰa��<%Rq[�P�7��V����N�ġ���*UԠ��ȡ���s1M��xf]�{��8e��-T~��������V7����11�F|~����b��ϯ�>��.m�vzXc�M݋�â22�7|�(%�C��_lMj7�K�D�&���ET�+o�+ݶC���q�s���0��U)z=]��w.Uk�<dwm�ѫd����K�1��`�o@a��O��Y����ݺ\1�j��vh��{<)�!���X�\�����ȇ�����:�~�:�G�!����n~+�� m���i����Ժ��2"A~xwrN�'9�03I�M����VY����KĽ{zI ���Ӧ������UE��;FL��==�
���wf�ŀQM� ϳrt�~��o�qw���|Q�)��F3����Ca�k͡��^�JDN�`ݜ֪�g��l8y�H�B�;�8����Bd(ٓ��P1�BP��]��������R9�C�j(�U������n���|��/�]��}�*��Iӽ;�����$,-
5��J���62F���8�o����X5y��ҩ�Eڬ6�7��U�ӄA��1����%މݧ�o2�;wE�7�z=�G���>��tO!�"�[�ݭ!�o��̍�t*�4�*Ҟu�kS���5������ttE@�7����u����9V·m{�q��٘�B*]�%|���dD#�b��0n�I����9Dq)T"���e��W��T�[<�~����'B���dF��'z�&�sz
�ǼQV�=���g�ʼ�7����P��a{�]E���%~�H��s�&:P���=�ß�jݮ!�p�`�@	�������i���{���*�wo�`�wc{Q����%f�w�c}ʢ`�n	}ǧB�0����k�����W؉�P��u���4s���sk��i�ѡ3��O�:ê�"����t"ugumGe�;�����V�+�Z��<�gMu��}�I",�ip���ݛ��Q
���Ka���7�7ݝ��Cj��e�����6�}�ڷ�ز,)�:8��V��R�>�]V(���tg���d$AH�d���:��)<��S�{6Q�@�m��b��>w���-S*�'��DzC��ЂAf�nY���۱�m�V:�Z���1�շ�P1a�$Se{�������>ެ�@�!9O������8Z"���f�;Q���1^I$��@�W����H�渶����R݀r֯����⍵j�ƺ潈�[�Ct􊙐���Cx�<�U��J}b�WWD��� ����,VEYw�<�R3�������~�;��~��{1��E9�+[k��>��V�|?[��as��㽎�v�čTU"�s04t	������s��]���������4�ڛ�Q�P7l���[b��ݡ��r�dlz���r
��J
|)G����K����je�J	Y��w��Xj���lG�Y��ۋ~��Oy%*����g9璘��̶��ڹ�Ump5��50�xVh�����
�ߺ���_>.�g�|m�D�`�5YT��]:���p(
3�En����릇�	L��f�C�o�񳸆����(f[1�Ѭ.��4�����Yqcn��n��y86w�������/�>���V74b�VMP�E�I��z`�o)��Â�C�8��Q��T-��G.6�S��
��Nmdc��xJV�Z�"�O^r�j�j:7W�M<�f�/f�وݍ�7{���o7����i�����H�m�r�2�����l�,��7@kC��N.�2^H�DAo\���W��ϫ�^��Wt�.ǀ]�m�z�����Z��oswt�co�s7�0�[w�՛�H��b�+p����?�8����[����_�G$
���ۊ2�>���v��q�L(ĉ�nU}��꿵M+佂W��H���|�.I��jZ����Gnl$��R�qӕ!�xC�)�u�p��0���g����@�p�o7gv��{={T���+y�hϚ�];M��>C�P#_  ��U}��g絏s<V3���������J�[v�A��FۇY:Kl�`��V:`=���p��nq.�����K�VR�<"\dۙh�N��mc�R���f��{�竓��r��{o��>���a7�v~1��dB���F���b���U�Zk����&ۑd�ZRBX�Q*�,��PN��i�ʙ�z��hѕIg5���AD݇X2�t�i�#���B�DO\�He�ٹ0�
y���6]C�p4�P�\B�7.BT���f=�1#����f��n��ֈI��D��k �qb;���7���"��W��p����y��w��짪��藉>{#�3��)���膍�i����"�^u��T
e���}�#��O�{vhc��]U�@Y��V�q=�}+F�s�b+}�3`�k"�I�2Wm���s8N4-�zڪ�Tڷ��\;�0k���fѵ�϶��c��[�k�������ʸ�5�"au蠸��z;�t�E����瓞��䬗�ʸ�*��v�y��ʩ��Q=�j����"
�=�[=w܊�a�2�k�"%��[:��Ld��K�`�>�*���:�o���v+0���U�fׅ�����f��(��.o>��?����I@��t�sK��*�v�UAon*�=4���e<������ vd1�b�52�*8�SmG��8i�,[ג5���y��zb�-��gZ5�FLã7��ٓ&8-�̕�}St<�=w�����YY}�D�Jډ$q��*��0��o-]�r�cIJV��4k�[��aS˫o!ҒۈÐIX��� ��דH�T]�za������z=�s<N��,�@Ί����2H7$�`�>��nf�VSڷ+bz�Ǝ��iC���ioH�S�6���D�>�͉�y��W�7��&E�f^@������:#�Yj_?M*��.B}�^O���v�}h��ؖ�NM��s��|6|w=���Q8������.�bd^g	N��I�/�9lMɜ�Z�'B�]����yfni���
qA~����s��]��١��k����9{:�ґ�UB�k��54�j���L����쿯z�f�nmi __�4�A���	�KL!���1����%\JN����L����*��Fa<��m���X]���t��}���G��D�9]�z}Ǐy=������׈-�u�?�e��8��Ö������6g��r�)��ŏw�j�#:o�g]�������A8bLwl�A���Æ�w<��}��Ɯ砙�L_v����	T�u�TÛg��]ۚ:�:J�Jn.��]=��M�b�M	�F�wj�ܠn��{zk9]�J��J��ނ�R�:Yٞ^yG�C��g!��5�C�bIN��e+:e��Q37@�"7Lù���ؚ�g)h7V�ԪB�(��]g(iC���@�( ٗ���Ix8���s�x��뗋8!t�]�Y����2�/ p�����ŭy1u��R����tR�qq�s���,�#!�^Z��4��܋�t�a���bȴA�[��c�SI�Zn��gj����a=��;X7����Ӛ�t��Ö*�R�M�U&k>�j.����QiꨧK�X	SV��0L�uY&�S���l��{�NW��"���o��wa�#�n�i����g�E,�{����f�r�\[̒'=)$ BP��
	٣p��$�Żd�7�ћ�L��VFh|:���K�������ʆ���K��ZK����v|�;�Z2��*��0+X��9���7
ttփ�|�7��\8*9ژ�.]�v[xY�k�de����UꈬѯM��N7�`J6���(�h�:�i�!s�mi5�Jvr0b�����Z	B�Ǭްʠ[�u����z�ˀ�6�6�ڢS<5N�7 ��V��Sq�(����U��jtU����i0u�մ�YS���݇��E��A��N�ԏ53*�S�S�(�MV%��,�����1YA�.��4kY���]�e�1�V��K�+.���)��QbYN�7���e�$E٭��Ia�bw0\7��w��!�N�\g\v��"�fu2�%,ղm�]Gs:�gD�g���cS;�@�8�1/(�u�\��w�9��j�7eM����鏰�a����RΫL��,�O0N��b��SAb���{��Eu ��mW��]�֗F�S���hP����b�t��P�s��j�aʂ��H��J�ۧ!��vR�B�Bx1�NwH��%��%ғ%cT�t�m�p2u��ǉpK&i7�+��Z��wO�"�-[@���eα�y�����R&t�e;Ѝ�U���ŻZ�d����e9F�N!`ܮ���nٷ��sA�*�w�r]p����l��9@���yqv�OMj��$Q��9�����L#y2�r��Xv��9N'�n�������H�^�ΘF��t�:R�^`R ;�V��\�m���o	�{�biq��� ���V�lE�u�Fj���թ�d^˔9T�N��«5U� K�Tm�"��(C��H�p]5x��Ts)�aqM��F�h��e$yX�6i����2����6�n��Gd���ݦ��<+�T�{J�gom�8�L$�d��C��P*��)�Dm]]b���^.��!�$%D�����rӂ�u�Uڿ����匑nnX�(б�$$cO�^>=x�۷n߳�o���/�@F0h�E�2k�7��Jo7��|�[�{�v�۷�ݸ��d		D�FI$�&Ti���F #�z����v���n޽{��(�Ye��(Nk�;x�wv�sQ�FjQ$�1��޾>��۷n�^��7�����B�6h���x��0���H��_17�����˷��LJlh	Jn�fA/�`�Yww$ι뮔���OϮ��܂PH�;��r�M#�B�ss��2o]�4"LO\����L�w"L@e��-2E
M�df �¯N"����߮������ÓŁ2'EDY��Qj(�l�P�IRPA�X�o���h���Sl�)��U*�%	}B�[���i��$�`.R��3\�Z/֐[ٛ�Y�z+-?�(i8H(��M�#I�L�"�l"�~Q��R1�Pa�P�LB�qB�A�K�L�Q�1D�5A`%�LI��p���1�c�]�����z�9��w�F-Y����ۦ�3��7%0doG�nWrG���Y02�c���+����`;����+�����9G�yZ��TR�@�Z_�KvU�y4ϸί�����`���]Us�U�&�\���~��ռ�p(�������7�����z��y��*02�/-�X+�K����=�g(���]�Y�$ϻ�nwgj��N��ԦCg�\+�Ղ��/�:��O�����s�ZK�^5w<���Q�k�2�m�,���-)�n+k�p�ۤD�p����������7�4æ����o������}�!e�Ԓؼ�$T��
.雥��o+O�!����t{��n+K��rK.g����}䫾�"(�O�[��L�����`Va�*k4��!_� ����m\����u-|����qw&t*�v��AaUw��Ɣю�N�yv�w�>x&�&���i�9��z���5�lf	²�Xf�T+Mr.�C	ܕ[�O,��IZL$�5��G]�;}[��� �j��j�Y�Zw�wpc��TO0���r�R���ޜN�[�wV�8[2�U>�s�"GL37��2{�|||||@�Į�KΫˍ�����O���U^���"�����:	�$�6Z�wjzE�{��n=�S;4sX,��*��'	�_�LVq�>�T.�YYr��p�����Ĝ�J�*�?\u�zC�L�#�>�b{��U�>�ߥ�R��>N�)Κ���x���㫨�21��U��[�{�P��<M^nխ��z��衰�Ɨ%	o�5�}-To�A§(qI��wѦ�rw��1��2�k�vx�5K��ǂ��I��,�]�ѽ7Sx���T�TL�j�~ �w��g��M����H��b��"BV��[�|˃1�;��٪�l�7���,��2��V�vώl��MQ�+���'E긎��~���Gp��
��/@4�U�?v
Ǹ$<�:�;�Ю>���B7��%��s��Hc+������3��`�Y�S��a�Ȧe'k������]�E�6n�ت��ٮqT�u�#aW,s�t�d�Q%�Ę��w�9`��
�|ȶ]�b�޺(�&e�e9�QRS;���s"�1M��Vq-��u�ݫ��[Fm�+Q��Y��ø�}k߼|||||}����T��9�
��.��q�gp�)��l�".~z6���n1W��-A��S��=>}�[�^yE��o�j[�u�܎��:��r|~-�d�'���lh������=ު,/*�����*Ȕ��2�P#�毁U���V�V����Ӹ������Ku��u5o*��D��V+������3��}�����+�)h�zפ\�O3���v�v{|�L�g���<$}�,U�/�<�V�)m����a��駏M32�(/�J]�}�|T�/1��{�Ta�_��K�sƨ>Z��u#�ْ(f�t�
�3���DE�9���T�w-w��q�H�"�n�>r��H�̞J�7��I9�.Wզ=��5�����<�O���ճʆ�\o\�*<ڽ6�������+Gʁ�!���_p=��(���@�<�en��a3N*pS�كu��oh���#.��҅��d1�*��+-�kr'��2�A�v�ӳQ��a9�{��\��"�Wh<�����vj2�S6p-
x�oS�V2%`݋E:C���+m�\�#RI�ْ�=U�%=�Wg#�mh)�������z=�)���T��t����)!�*���B!)z+���0y*sQ��$G�Зor�V�?�FǺY�/� #}����1[[x�[?Vglۭ���"uWJ޳]+���y����bv��~���ϸ1VJQ���
����8�=A�M�z���d�c�d��*!�'�Ӂ؈��j�i�B�VZ/��'|H7<{w<�f|��{v��HՏH
�\��!��x76"����x�Ȓ2��r6������긾2��ysi�N�礮3²�v��xj)	�tc�wLYs�C�׻�wji��tSǶ�w@!)����~���:�ܓ6�%���J�n ���sݏ�>�y4硩
�K;��`�5���)�λ��*��=L;9c�6���+J]}��&�歧ͱ��v�������wYsY��x�:�ga��U�]'������d)S�f:8��&��l�剉�i;w�]"6z�d�ox�ޮhh[>Eޗ_ZN꒩�KQ�%}ov��P⤼B�{�hJ�Rrh��hⵗ4�ެ���	�U��),ݧ}ױȝ���D����������X�}Uȇ��'wf.�Ks�*i�eCedRq�2�U^��MV9�N�9F�Y��1mg��jYc���K�I�^|��_ƲI<�u]��c��G�iK��s���*x�[(��<8�U�y�4uuژ�/р�ͩK��E��2�Ϭ΃
�˰��hn�� ����:�M,���o�'m�"�=�=��6���d���!l��}�ZǇ� ���44�n��lF��:h�(����^�x�`��C�e���og%�v�e�7]c/�n}ɳƫ�o�R^��M3�v�F����"������-b^WyT�zt����֒��&���\�-�y�&��c`���J)�?G�p��
�z���|L#���}gs}q�Q�/)��e��0�����5��!��t5 �����`+�� m?r�n�����5�EoObA���p�=� =���]��	^�k������¥��o�r4��3^Ц�
���O���M�O@�=Obm�mK���\4��-��jT�p�,��9� ��T���,�JP�B4��dh;��3��Q���GER�U�V�ZQ�e��Ǹ�.�\-��Qݧ�IX����y9�t�^����������{Zz�a��ڤ�04��g"�d�K������|)=V��V��B�\�&�����u~��X����f�)�^elȏS[z����+Q����Y���!B�T��H�!gS^K�����F�)�N�G�R{��Nm/#C��`ܑ���M��+�iAH�$��M�	���HR�b��E���7=�>��N4f���=�5L/��m�|��G9����v��Nr��p�ԈF�E��9ɳcwcgev�0�:s\7�rY�*�$UP~��R4�l�w�?
�9<�a�9f���8Q�@s��!T��<h6ɞ:�獞m����R*�7Ay�[��
��'O�y�|���&���2��Z֜��]����k&Ϣ�9~���^��:�5lGT�ߧj�L�.y�Q���v:u����S49:k�ʂ�M��;�V$|>�Əq���IEҽ�iKS�om���hyZ��^fe�7��2��b j�HI���=Y�����������jRٳa�wN�s���3{
���;�7}�A�IT���E�D'��G���+ɧ���aO��|�Oo��tT��Su�zpo%4�z+&��`���du�3x�*F[=df��pQ}�{ԡ��rmDD�&�-�J���4���F��r�cXP}�����8�z�kC<vuJ�����9��Gy����t}˩؍�Z��	zP��|�Y��)iI$�s��J���c�jl�
��k=��^^��-�BA��=��u�!�J�7U�-v�I�s&��7�m�օ�U�Go8o��4�@��Q�9)��t�_6��Q�][��F����i<�X��'ss�*���"a9�z��ղ��+VףH�Πt�o<���=T�zn�r���3{|nH�{� I�R�6�k}Q.L�� ��'� ��P���ɀ��n����pQA%����\�����zƧ�EfР��.w!�0�*������|˨����s�0�	�������
*IW{�籱�T	h�l��k������ʄbݵ��:�h�Ư��s6ˮ��0f�j�$�swAΝ3NE�p��bq6�j�����w���V�����~�������xF��qά7B�V�y۶It{z%$�y:ޒmOe��;2f�iv-�U/5[Φ�>�>�Z�"�� ��rR��jܷk�,\kg�{��a�V@&��X	�C��������|����CL�7��	X�6�:;������wi���'�^��\h[
�3�
1�6Ѫ�a�rQ��6'Cl�ܡ�i���I�$�:T3������~\j#T�<�,�fΊ�j�����؃��}��U��6wJ�����؃f�a~�H�@���a��~�ΧV��vu���H�Gwz����Dѵ]ml�t	�4sUqx�ڴ·X�aX\]@�J}z�� W{h{�m`"������}ӰÈ�gNUh����4Lp>�@��a8�Ce�%>����ZW@7_p��Zt myW����Θu�EѤ��;��,�����k�1�]<���S�'�ٯ~^���,��/�"�-5��N��\{`��K�̬��Ӻb楷Ivr��݇�r�7�\�R>��j�d�{i�3vl.��Nt*�B�`Fi���0��;a�y��]�/6-.]�f>z�a�{�k�Mb��td��{��������c�60Mu����\9�(n��A�nq9�Y���5r�hY�Q ��r3��c�g��׌ť1+�G����SЈ�%��X��C�Z�4�9�3`n�%w&�m݊3-�=Ϻv�%�n��X��u.{]�˵��J:��|� &J�_�slDt��^P�azke�j��!s�.by:�SQ��:.%S�����u���C�ӯp1�1UO��+",�#�gB\H�QU�<�D�_grݗ�:6��cL�i�>X&��N��;���Q��-��M\�ͪ�\�{��y���k�Rǟ�@P��4\���x���U �U`ђGg_J]��[v��b�A4d1�d58A(G-�F���\���=Á�x0x��۳+w"�x~����ܜ���
�1�	�m���T�@�ù����K7J`-�F�T7�ˢ��Nڜn���3�ƈ�&�^�T~�҄/���y���Ap�܁�Cn�ש�>E���PT�pK[wrv���)3(ڭ�G����S�����	�y ����O���#�g"�,�7��&]�{�v�墔�M�gi��c��,����j����8L�����y��o\c�<X�Ǥ��u�&���䶁D�T������T7bN�1rGZ�+���`�dq��e�AlW͸����p7_�������_~����h�j����13�,���2�fDq�4���.��&�(;�h9J�Y\���zɰ��a� j4ic�X���kD6>��nپܱ:��G�N娟g$�- Κ�G�yo?{�|��+��1Ļ�����羮Ѫ*�E)WsS�y�D����Z'o/Z�C(�����u&���V�$�`��2K�oT(R*�-Jv�\i	i͵m��퉡ޫ��\#`[q�g���Mw�MZ�c�|�J�P=�U+�9Wk�v��o{�Fa8�v�m �fH4�C�����>��&Ό�f��tF�+U�J�ͦ��q$v���4�����PM�$P���r����b�a���~z쫨��@9�K4��0�����5q�z�唨ţ��\#X����^:h�׏)�is9��u�s���=7ѕhoBkT�ɋ7iH���*�+t��B܇���ؤ���w�ظ�����QQ
�K/�
]�`�Ӕ�v/�x�B�i�_ �Y�u��V�r��[�'":���ҩ��}�����i���v�Ee.��l9��7H�TtLǮ2�*IA#��N���vr��$��c�8�{�rP��қQgIˌ۰����ŵ���W1�jIM<\�*#4*ͽ3I	�;��J;�lk�K驢m֥�&��zƐ��n�ZzL�������g
Vx��8�9p�4V*ӳ��i,I��-e�a�4K���38P��������5�+�7G��9'na�k ���h廣~��y�^+�݄e��@�Zz���V]��YV��4�/U\�We˴Uf4�r�j^-t;�V�o:��UC۵�#3���,�/X��hE�38�-�%���P��B���+kJ�O��b��{+�Gk���fV�tz��+[�����ő:�*m	�5޺؍ebe]�I���Z���F.񹡈l۷�U ��~R3cV&T*��gnm��g)u�wiTȜc��+I9�b7	��X\�"��a��P2T�崙UX⎔�DUG]�s���g���bW��3�Ԙ�M̚n��[���BX��oP���>�D)��7ػg��s5&��S'�܌�D�u��'C��J���[_q��u��9E��	��(P0f�F∖$�/B�#�s�UR�̲�b�p�՗�j�k��Wn���R��
��zmuJ��^���;Xf��������&;�A�lp��1J�X�.�`�?ZME�N����R��T6J2q�RJ�,�c{$�1WEs�:v,T��]�z��2���;v���u=Uظ]ͭٙ��L�wz�`W�R���]	*�.��]΢#(vM��f�hu�fΣ�:�rqi۸ҡ�M nu�<�[���%)C+*3^T�F�d��zVJ�M��e�[3��:�1e��ǰY�aokW4t�Vk;�{��M��1J�e���a{�;�����&�|0���*;Unu��+=O3Nu'�D�;�|҄�R�M����u� �$E���Gp�eХHr콊���J��U_2 "���h�oV�-ܸ���^[<؅�wt�7�&��e�B`@�ZɄ���al�d�ۉ͘O(n�Y���x������wh�Z��s�W}W���o+���c����b$mim�]�/�C���6y�E�Q�C{��;�ʵ�Yx)���O��B\��+`�
{�΄4�Xۜ�6���y�Mb�U�]В����� ���(�7�V�*�w:<���i�n�$�Y��5e�}>��ׇ�D�*�i�}1b��Y��Wvm��*i�@U0��G;���ATՒ��wlf��Q�Ls��F��k5I$�A �A	�C�Ћ���`$��fI��jv���ێݻv�����׺�D�2TbB	� �F��CIjf��o�����۷nݻz����I!	#�u��Df$���9v���H��i�޷��|�{۷nݻv��ׯzFI$d�$$Ԡ_��"E$�H�DD��7��&�a�׮޾��۷nݾ�q��ǅT�*`�&�3$i����=5�(�oJ� (JE�t���[�rIJ����>�JJFAj����l2��܅�ۘ�,)������1�
1��/�nQ&#XP�t���2M�\$ɼ�K2�̦x�'��2|v@�#"0��)��,�����&�� �|I �H�gf�9�.�z�j�"�\mkrt�9����aٕ�5��H�p�h��l}�K���T�p���h�a�}��z=�@�=w.�r{�/W��h��H���q�N�i�n�-�S;�p���p�ֱv'��}��w�_vr�f��%�ݓcZ@�:Є��iF��Nc�m��v/�ix��ֶOd�2p�`���1,��_vm7)�n�X�����������������Q_ug|�/�β"�"b����/e�z�"%�úw��; 5ǖ1��`ζ�U�߾�����]�x�nc�����WCi���6%0m����=��b�j�%���=&a�h��ө��^���Nx�<F��co�I���5��4N����Y���^ƹ`�����럟u���3'ε��:u ��p���q��z@�XU�WG�׳��6�$9�7�m�6=�i��u���gm���M<�T=f�l��7�����q�C^��gUɿh%2C�ً�ܴn��&f���1�::��~O+l�!Od=$нn�P�Ÿ�nN �1�C�U���HS����&U$�u�����r��Ŕ̓c*�z4���In�8�,lV�z�D)p�R�a�b��L�+"$/|z=�G�y4��O��u����~����:�������j_���1�)��Z�^Kv�O�&��� VWj�Y������OJ�+Ϸ=n'�o,��X؇������v}l���Y^��OkI��qNikC�Ön����[];K��=$���\�g#�Pu����D���p��)�l�{l�^�y��i��U7�p��6�䟯�I.s���7���ؽk��Zy�u��~ѦR�2���ѷ1�V�]x�vrRJ>--�ց�57��z8אyڝn o\�ሺ�[�z��}R���G�H�K�s_a}�_z\¯p�.�J�/�H�VzQ�~Ow�f5��:������Nl��"��-��Yޑ���"
�.�X��t�r�����F]����k��*�ŏ��2���̐F�#7j����q#�R��
�)c#�������Ԡ��T�RD�=1O��l�溄}�%;��L0�@�HRgw(0s/�M��\;�*���0�\�^�#��U[a@��L�T4M�Z�q��{"�R'&��M(M�Ӕ�&dĚ��R��> G������q&�[uj�syۥ�UD��$n7�1�S�,�Ռ���&�f�Dxc��&w��T�q��VW��R�*�;��9��^ʥ�(�"f����G��yp���4���H��~���2Gv��"�t�=\-�:�A��8r<�� %)��������А[՟e]�S���>�=��En��������j'�f��k?�����ݝY�}�X������C=FbཚZ
�5�0f��g@�!e�+5<�\^�<v���~�Y�k�Cp�ɩ����S�x��=��J�3u���a�떃��oՓ}Rh����@�c�gc�籧#�9~W
}س{E�-4�z���P��Q��u�6����Q��U�B\����	cảʠ[��[m_�E1q��.��gᶲ.�
ȊY�vs��JUoY�1շ�t�%J��~��D��w=޷�g��0q�	����]	qng�ꉬ�ۈ�"��R���x���]mǎ��鱪���1Js-%��
�U�:pAH�����Ƶ>���?�B"��ܾ����f�R�+p��.��1��ܗ))w(����.�n�E��Nd��f/[aN[��C�����z=�ݺ�.�{6����j�.C;��1����~pn<���ˑvl^��;7���s�ټW��ҁ�ifp��ZEJpYi���1�!Ёn� �g$�:���	5�ڼ��ϦV��D��@n�f4��� 4�4�5Ί�S��ﴖ'>�1��S�f�⊃q�����8��5��B3/nYⓋ���u�����d��_W��^k��)g��+=i�a�4K�z�h��:�t*����D��y�s�ņ.���r}-a�d��V,v�E�͆�F��X���`�[�1!�d ��!�=��x��FM���=I�}<wV�fY��'F��ٻ:[����vݢ��5^��	�4/jh�5Na�G�Wd��w}�+��\WWњ�����]�EvY%ʿL��O�&G�����d��C)�P�nn&:2�|Y"��k�d�ݼ��D�q.3��g"a�4
��s6E#cZ(���U�������ҧԉsXj�Ds������q[Ҹk뎻�o�n���Ɏõ%�Y�ޔ{4�27T0=�;C�קּN<B�k7�Sf���5joa�S�ػ�Z���k2�ߞ>>>>>>r������Kfd����.�p����ݽ�S��=�OA#�\i�ڼ�b>�+M�W_Q�YOy#q��x���Qad��3��W��:�3.�
+>����ju���I���+i��P`�T
�ޘ���ڦ�5�-`�,l\�6�p9�! zuW�R�B��v�G+u5l�9����k��5��e�"ڄ����#���/��<Nk��Oy"����t�K�Kc*x�^���怙^B�����/�	-�\k]��]@�21���7$�{�F3 R^r7�8l
u��z�gr�R䚽���-�;t���8<��/:�#���`�ޅ�F��.2:�|��\�Z�0�P|�t���W�^�y�]s��m� 5�o�29�#U��
v>���W�s�O�e!L2�|7 �1@ҏ�����#6��;c�u�S���a�oj!�V�hɻ0��Z	�gUܘ�	nc�,�U����{����Y��7o�]v�j>mJ�� w�
�S�]o��{��^V���]�Ϣ;�unސUo�MuR�.����qW�3;�,n��5MZٺ� ��;��*Vߦ0#�9}�9��Wr��C'~�E��E�v��8l,�z�5KfDC�2/+��u+�PG�v_)����n����; �\����9O0�A4�l�:03o�Р����J����H��5����w����~�\���!u���8ע�I�Nz���g�r���MlH�&R ����6cZ*&���5w��Q���t0@B���n!��b+&j��b\TY�;O���Eu��s�E]h�݈f�X���_�`�k�����D=T�z,�%�t��Tu]�s�c?��$���S�Oe��ȸ�:Z�ӻ3�r�[	%��i���f�����o����� �	<)5UQ��駉��M+<*��=�[��K!'͔3Ү��.�gI"Px�y��d��/UQ�`<)�w���9M�cb/V	e�l�;0��V�����b[ȍ��y1��^��l�T5��xaH>�+(Br�B9R�"��n'���.�1OH�{��}|�w���P���-9�*^�J���#J�^��&�����vR,�E=ZY��ڱ���ޭ�ݩ7�e;V��%����t�}!��v���J�\I�I�G��������w��5����J0���%�V�{���NBM�
K��~�M�R�ԍ�����QS��3g�������z�f�k��c��F"!��,5��I�,�2!t
0E�O�*��o6ہ�]���\s֕����̀��0j��BW�埩>�μ���q�&��GdVoUoV��Y�+����{-���u��۪�Ǌ{O�K�2fDN{i𯚻�����+h����͝��7J/FfZ�~��;G2��c#�E����P%���A��qu�h�٭�ӡ5�/��c8:R�Q��Aw���}"U�T���'�f�&�Y��&�Y%@�ǭ��T������<*4"�>d`[eXg3�Ѭ��Ӱ�N5���(��W�^�r��,���WW�%o��e3�U-<�3�5�{�k��k4�	R������d�U��ó�@1v�Տ��3)*V������lܩ�4�A�b��י����2��ݴ�D�	���:
{I����pemɜ�L��Tq�ԩj.�X!�4o`#&�Ii:�5ڞV��5י��nVo6�<�B\�����j�^��������K.;A:(]n/A��m0���_1
J�(���o����;1�J���IB����@�FE_�׸+ө!}@K���΢�ǳ��o����:Bי�u@ۛ�]
�
Y�#��I�;�CD�5���9���:�s�B9w;�3T�9H�6�U0����ޚϴĥ:-4h�݊Z�F�H'��0I���n>H��	{$F����G����ԝ�;��"���Q�L�8��"�7I��{���>� �u��5D8��������S������S�}�Z�+8��R�ev.m`��0�����|�g���O���^��<�l��Qݷ�0o.y���wdڙ�n�Q�������b#�=�����=v"1O�fwf�y**��fハWkv�SVN��oޓ=K�p�� ��vL'�fg�Z �yi��褾bf��7(�)�v2n7�W�v�c5�
�(:�(�k�%wu��U��e�-���i�@O��'���8��C�<�7N�6j����P7w.��D	ku���iҹ�w�Q#QlʊvfFf�nB6޺|,g�xuOƎ����4ϕPKOMt��d��q�<���`�Ԝ,��>�����o�$�?_e-�>��y�'�s�9맨3���xG���>囉�F�Ȧ���:d�v\/]�B�b�\��wzA���y`�*�ﯢ�.�����.o��~�G�>W�6N���^� q�ޝW��S	��Ԝާ�#�C3����Ar�w�5S>�u��^�>�h�`pMo:���V��U�@��#��6Z���z����V�*�`����B^�+��D-�Z�{��ʁ�,D��hdE�~<�HeTT6U�m|��L)y{"�U�R���c;.��ĵ��o:�P��K��
�C�vd훌aI�E�1/�^ג��BEU����L,�r���xa�=r��3=�O����؜@)���i�L��'�����v�(v�_�yZ	ʏ4^veK��}Ʊ��C|u�E��!)�ެ�l6� i:��Y�-(Zڊ��sX[e&�I��H�9	&�D�S7ut���2�W��������k���J�o5%�OT�Ę)�峗X���\�^@ٝ��!�K���kXʤ����]��f���]9�v�SQNc)<Vw.0�Brc�9t�y���m�c��7V�Ap���o�'�G���w�F�����8�b�:��Fv ��ș1K������hgl��S���u]" ��9�:���HC�/S+��q������Q�4��{�p�\g+$������8�W��q�~\�/��:�{��X���꫰���3UY��#�M3*�����ļ���w�	=^v;� �!��XCv�ݎ��` ���0������q:�{�����W�x�}U�'��e�+��w�}��p�O�W�R��̺vh��}��J��]ޣ�޵;��r'ל�Ⱦ܎z~�D�(��2N,�~�kN�����>���ސT[�5�I�o��&��1>��L������/��?©�(�
��* ��������Q��*���>���Ͷ���j��m536�j2�J��j2�1c6��f��1��֌��ɛ2�1f̶�Q���YmS3mK&L�fK&V�d�Zً&ki�k1��TƦ�L�3U�f�MI��fjU��m���j2�L�ckM�c&Ue�i���2���&[l�1���Y�fk,���&L�i�ʶY�mYXɒ�Zjm3m�1f���Vf٩�J�m1c-�ƥVVm�bʴ����+6��eZeMM�,YkK�m54ͭ+5���ҳ[J�[J�ZVj�S3kJ�ZVVҲ��$"�
@[��eel���������������[+5eY�����VVV��YY[+6��[+-ef�U���[+5eel�Օ�ee�Vj̔}׃`7� �`�
��Z�YU�VU���l� ��1U4�B 
� �T��U+5�R��T��@ 0D@5� �DU����R�֪VV�JͭT���J�Z�Y�� 0��@ 1P�J͵T�����کX�� ���kZ+y�����֥eZVkR�mJ�jVU�e�5��H4@b��$(��J�ZVZҳm�,���Q5� ���R�&mib͵++i�KjVkiY��56��V�ZcSV�,եfڕ�Աek+5iYmJ��jS-k���ty�{>��� H�� �b��]���{��pk������������w�p{���kA�ؚ��?��/�����QW���?o��#�h��/�`� ��8���@b�O�/���������� ��y�����G��4�
�zl?G�a�br�����~�D�{�k-i�V�+iSkF֛eZi����)�MR�%�+5���KRڕR�*j�٫KYmKR֚�iZ�Zjj�Zmi��i[-i�kMl��ҵ6���HE"	b�"	`YV�eZkMZm-iTզ�kK*�l��ʴ�[J��3kJm����֤�SSZ�V�֥MjSV��M���֓kF�lʬ�"(�"���T+���mZ�����*��Zf�I�I��U�kEZRڒ�%�J���Z�BD�K���%������O�
Z��kh�Uj���?��~�����'����>�@Z҃���_�O���؟���?�?=�HC�����?���@_���D���?�T U��@_�C� �X}�*�-}�:�"� ��
�J�k�OF�:P@�_����#����
��C�������
��m$���������/��?pA��X~��҈ �����_�" *��}��hXK)?���4~ JO�P1��à� ��8,��B ���{?$��
,ո�mz�L�����/�>0(:�h��-O����o���4���1AY&SYZ)c& +�Y�pP��3'� b?;�>|U��Q*�֖��)$�H�(����
��HEQ!P � 
%)PR�(T�����*DUT�JR�*�R��
P!@*�T� �*IRUU%PT��B��Q PѢJ��TT�@��"�iQH$�RHRZ�f��$*�@�*/�u�l�����h$UV�!%EJ��D�J�TJĩDJ��PDA� ���D�*����B�ȶŭ�    �UO/wWv�٤���u;�
�
�7w;�D�v�u��2�;�Yڶ���v�Ӧٔ�����n�[P�ݭm��ݵp��ږ��m.`i�vڹ�KJuH�*R����k�   �{
(PС����ٽ��lHP�F�wO.�B�+CB����v��7m��ݗcK��l���͝�\ks�n�WF��Q���[�t��lksN��YNk�]��Ϊ�Q
P(�P�
�:jx  �{�j��;�g#Z���t����wd�Ƴ�7::b�wn�v�ڕlX��u�:7]�:؆���Ns���ԧ\�+���������;��k�Y�R)PUERQQU� ���k�\�+:Ѷƕ92�˭r�:���w3[q�ĝ��G&V�Q���u�v�;��۬���wUnZ���Q4\��R�T
 ��!H^ �N�K��p���l�#l�����'4қnj�f���n�ZWjӸ[8��n:��v��k���tlkK�L�Ys!$�%D��VڶEUT^ m\6��5n�nl�]����sZ�gU�V�.j�1G[ZmgT�h�ε7Q��+v�须��50(�Իwk��s��I@T�*]�l��P����:UR�Rg: %�j� 0R�"��r� ��SrI[t���8����t�t���Wr�B*�)
�d�  ���P*����R�P��M�V��*s���R�K�A@���5¹R��`$�S�-�
;�)�9���P.p� ��R* TR�P)T�  �ޔ h�P�e

p�Z�w*��hSuG�4)K�.U"6C u@��F�(QE���]QEYq�U��K��$$�"RD�x   ���:�@\�`4u[�TN�3��U�����QÝ��n�r �V�����n@*���p�P E?!3%J�1 ��a%%P��Oz� )� ��)��h� �=��	R�0 #'��	���  l��u�&c�����@{D��B�C��T@� d{"����@�$�̉�@|>�������=��jޕj�j�U���_�kZ��mkZ��[Z�٭UU_}�m����u	P����?�� PU�J�֑˹F���4�+��)��NQtm
L%L�����QVD,�;F�7dvް�ݫ̼�t��E�mB�論�2K�J�R�%��J1Pc���v%JP�/(YL=oUwBm��a���I�ZƲ��EЀ���z��Iv�e��;���0�"9@[Kw��ʜwO��ӳ��%JMh�ȗ�����/wb���1�[�T�ٛq�R�`'OYH+���IS7���a�i-���fY�Bԣd)���n��%�61a�h�t�է�M�*ˎ�J:ͫ����N��x�e���B��4]%�ebwG2�i�-�G�i)	�bX�UX�]GM�Ĥ�v������-QV$b+�D�ٟCe̬N��QPYH\���skfe����%��[O-+Q�EfT�P�B�c�Ց-@�������@b�iT]�)����Lee�Kh���/sF�ݣ��$��4l� �:�\�<�;D
���`�CN�W3i��N���m'�:H@����8�nJ�zq�Z�6"�V8��M�[�˺@��RH�/2�A�bj]����3�x��� i���V�Ƿ��"q���v�$^[Ѧ��E(bC)&�a�F��`f�#��2mKǭ�13N�֊���RvƦ�a��{u�
�	H� u�%d+t���"�Yvh��"EBH�,�'A�ԫ8lP:רf�Z7)* �oS.����kU��c�Xi��Nm�V�hyO@��tм�43R]�%nޤ�i3�ؽ92+bK-+���1+v+��Te��� ��m�rM,M�uspª�&�T�7�oi�J��[���0e���Vf��u�Sn�5V��[�#�6)�b����1!' �N%�f�2 ��EHa8�ء](C�2�H�Պ��*,��P��[&��8�י7�� �-:n�M֠pv-��
m,Qɹl�Zw���V�-�G2��"i�eM�Xd�m`���И\y�'vU���0�#2[���D�aP�d�o�U%�nPGta�Fe���Xd�ƅ'�2����ܣ#�+Q�	��V�����fګX�kSB$j[۔��D	�둷@�v�m�ƍ�r@Wwi�FI�0d{�k�"�0��Q��w*F�5�$�@pe���"9md���6nI(�%KQ0�:��W��Ҧ�X.�����EP��c.�����D�(�vvg Vj��a4�-��݃�VP��T�
ҙD�7,3je�m͘V16+�YSL�l�+٦��rt9�Q���K7�@ �((&�-�Y�7	*Py���^�[���x���SE��n����E�DǇ1��fM��I#��vu�Zs"M)p�3t�!�g-^�;Y�
'o5��M9"-��0ʺr$�Ek0R����5:�5�s%Z�d|wm�#Y��` �sA!V�TmD�� a��Z���@��]fY�w5ݸ��5L�	ʎ��J�@��Oh�ڔ�!n����J�r��#n�Qñ�k�P����d�'�ؽ�ő�aF-Gf�r`�
.^Kq]�gi�۽��8nd��h��N�4��0-�t0�r�����Z+[ʓr����&�l��`��:n�Rk��ҩHbŎ;!ݭ�	j;pG�i���fQ6��D����<�.f�h圛��V����3kAm�Z����[N6�Qd8�n��S٬+��l-���F<�����kA���ì(�kN��b�fc����Gf����V�arFΕVO�LRՋ�h|G	F��uYՐj	:���v>t
����Gha`h$�7+n˗
Z�Jf��VӼD�)�;�f��/��r��'H������@7q��wjU��8�;��f;0��V�I��}1������-�����I4�q�������Z� 3.�̵�lj���=lj��hø1���6�]��2�ߝX0ݶ�zwii
=�!PU��ayDQ�5*��$-����j�U�+m\�BK6�!�T2�`�%�b�[�u�*��&��0c�iۃUw�,f2�%{�t�!�c�	�u4^��u�1Y��ס�а������ �^b8��Fhv+DWzڔU�����i��eYZ�F�V���6�"�J̙�\˥�Ut�t�ۡ�&dp-�[��'Z�a�4m����V��[!%h��]�X�N�;6��4�j�*a�%X�_`
f�b�?��*�,n *6����C1�����أ[b��*�L4���D�װ���$�6�uv��`�K&ǕwSn6��|SL�E���`p�U
�3t��Mab���QqFZ�ge !��<XV�D��"�����!��l\l�^6jMj%l$RJ*�����^�'0�����{.�(���l,���!T���@;���1I�ոd��V1�e�A�����j3P-;����o����=.�����[6؟%{�v��iM&�ٓ1�ӎ<�ԛ1�:Q��ñ�h�o
m�-P��M�ec��[ԳyJ�xēU!PB)��At�dr­�c\�F�U4]��JD��ו ��U�+���Nf1F�a�<�ī����(Ʉ�4�qD�vS�*M�u����5�5ͬm�/J��ջ'CZU�aű�Df��o�b�=�i�4����7iǘ×���6��^�s6�`�5(�F�[r	w"�	ID�g��b��))��lT�ފk!ڰI�bt*o̱�^۶��B�5�^�� nm�Ijȷ�P��2���nH��R�u�V�TJ,ڻǛ2ܖV�6}fӈb%�V� �Gc�����'��m��3k0�"�`�%A$�+��Po��� Y˧Lu�v�܁AhZd�=��k�M�A��;���Nn�r�4�g�������j(�jэ�{��N;f�,���XN���յ�Vj2�b����˹2<�-\�l��X U�`�ЯfR�S)6$pسy�,�$j�E^���/&�0�� ��T�$��/Z�L��!-�+T���u3��(�(*|��J�-&���Y�р����>�2!�M
�ڔ&�0��m�����ڷ@�LBhս7��zpํ�)	�Һ �x���n[1'���,c�ն��wU2v&Vl��@��]9M"X;�œ;�I��Ī����F^�W[�	��t�eq7�p�;)�*�%k+F�I�7�--ЯC4ىT��F�cXH��'��r�k�]k��0V����L�7CTŒn�9��h%�7+Uܧ� oI�qɨ���&�[_��)�OzƢ��c�2��JJ��a��+]RB�E���^�"�Ɏ����ƶ�"��%k6��ps0,a�����eQ�6#ƛ�v@,�
�r�Xl�6񚡥�����k5͍
� �̌L���ǙcZk6�S(�F�F��O�t�,u�v�湼��h͡9;X+�as	{��-[�0�Bԣ!�!4��::	��CM��`�u�ަQ�]SK��)
�n�����iܶԗM�>[/1�4^��C��h+�,@Fc�7AJ�2�շ��;1��2ֈ�ձhcxQ`Y�IR�z4Li4+2����IR k���:,\���k5a��1C j��0���Ƥ���w���ڛ�J-֊�-���bX�"���v�J� �X�\��[$��N�k����VL��.��eڙ3FL��4�R�Pa<��f���mXo$ #t��`��,�X�m<ZB]�����y�1�iJ{)�6�2RaMĖk�t4,Q�Y�ö�Muu S�P��PM��EX�O	yxˁ�I1Vhؽ �uϪ/�-��TG!��[� te��3gQx��E�,Qk)�dU�(�ͬ�Z�J��nҗV1VQ�hiR���Y��+jdb(9��V�\o0�Uv��R�7�i!G.��hV�m��k^��f�\U FN���J�����Dhj7��i��QHK6
��T�u��Ѭ������̠��n�Ke:��wZ�D�ex5Gr�J�,h7�F���w�`& sf��9��)��In�6E��t1*ό�X:B�A�Y��א5(el�[�h����((�DU0��1�X�GY`3VjZ cĮ�h,���]l�0��@`,R�z��b�wzw���^�́���īBꬅV\HM	�f��j<�6�E�zYT�`��Z��ײ�����M�.�1���)R�oH����.Ժ
����w�%��h�x�Y#]F�H1�%�L����yXt�L��:��B��͹r�r�7zE�bd��JP��3*mgk3&|M�]���{&����ӥ�De1���eyT
��n�J�m-����%u.U�b�f�M+�܌8H ni5����$J���B�p�
�.�c6ٸ�J����]�Ph�˵�RP���֧XՈ�wv�$���73k&��c�F�9t��uЍ鹔�LźCQ�n��c�utm��M�V��ej��FZN��@i5x�T�Q�)mm�z�:ĚSP�V ]�8F�xu]�'�ި�(�E���8��i�T�`ܬ��7%���B��74��a!vc�&��:fJ@�ፄ�RTo�(cQz��fb���U���˽&�tڈһ��S'1k�WR��Q�FÐ���A��i2|�5�L���p��±��S�HJ�5H`���;E4VV�4�#)�ǵ�
��B4�̎FQ�v!��I+�v��[	��P'a8��tj��b0�x�ȷ$F�f$,��CA�Mѡ����1S���/^�Ń6K�͠��j�c�o^K� ���%��f��u��ܴe2�P
����L	ՕY�#�F��jOD�%f�6""*:��͘�nX�p=JhR��xwv��d[E��Sn��2����'Q�z&�Q��,��ܗi<��b��+A�4f�����vi�"�a	(M�K#����NS�Ȥ�C>պ,Њ�^�O䣫�nV�In�����.�wt�5Eǒ��V��k�[H��Zg	zAä[Ū�bZ�ɻME��IK�a�^U�ġXrP�̥sL�ňwH+%m`�$ǅ�v�Ӻ��B�=z��{-B�����R03K��`Gi������yYm0�'�e<��s)\e��i��Xj��hM�ū�a���2怍��Dd�M��l�hfԆV�-Vة�]hCW	�J��E����������h`%�W���=%nE�$�j�V�ò��4�L�a� Ǳ*�K�̕���j�\ʕ�� �t���dժ������n��.)�v�;'$-a��4.�ݺT�*���m%LY�C�r���'���6��I���QU�4��&�@Pl��*��V�J�`�aªVB]l˽u*d,��t�) ��u����̩�qm<pH�6�҅�(�FrQYQ8C��A	���Rvm3���vsn�M�`�dE�f�U��E�+
�|�kٙҴɭ�����>X !�bP�Ǖ�f�Yj5*D��`��2�S�h7�8��e|�5PA�"�W�hYBv�dzݺi�R)�+n���/�B�#3r��K�	+/j�&�� V7�*J*��"�%J�B�E��`��;4��F�Jm�̈́p%Fћ��V4;ڏ��r۽#(~X]�K,�9Qm�QkM�,�53%�Ѧ*��`���;y[�Q�z�Զ�H��&�)F�E|��v��R���)�7-�ִ(���X�,Z��ov��'ؙ�1�e���tz���Ĥ�-H�LϬ+�ΕPEn��q�YwL�o~�qlr-���Nd_\b�5����˶�q��J�f��.�:��� tnQl�z��ڊ僸P.�����z*&6�XQ]=����u(˧��@P�b�ʝi�N��LJK�Bnh�w�BE$��SU�[�M<�X��ñ����Y��鷆R�l�����)v��ӋP͊;t�{|��r�-�t�BImklb�S榊Z�$�m�8��A�>!B��#*?�f:ŻY���i$�]���y�W�=�P�\�M�6���,yv�f
�oDx~�TH�N�Z�n�Ę�A;�v�-Č�Y���x,�!�b��d�E,U��X�e`e7t�](�uaX��o��\;��s #.VṲ���n�o��N�O&�e�|.��[�*o ��)Q; ����`<-T�N�^"�V3%-5�J�&@al�D�ݩE���9{b��������I�(T�c �;%��Y-[��� ��1b�l���u�l��4���]<Vel��� ��? N�D�H��)kkV���*ʔB�~@]��P]i����P;Z�w$�m�
Q��֜�.n�p�v)(l��/w!@3vQy.�h���+iD�3CM��r�U�� �홴r���j�^������n�;�bN�YmU�hx16r�#�e���/St�E�z�7xּߑ�T-�-��B����iE�1U5l&�d9vc��T�ܘ�bK2���n�V��XHkw�����ZXe��B�˨&8-Z��,9�wBV^��E������C.�v�E6�enƚD'
9���t)9�F�jbX6�Z�h
cy����"J����iG�*��Z�ff ,���N����-�FB����#)�k+q:�Өr��ʲ*�+�(Z8��%ZU�����2f���%�ۤk\�2���m1h��9LY%C{�� ���) ��jř[�]Q4#Jn�a�;��3Y ��� (��70�����p�5S:�`��YP`,�l��R�o#��,��w���%a�Ԇ�`����Y�ɖ�n���:jSm�.�(�e�I�[�jb(�K�GtoU�n�Q��n=[X�qd,&D��/>��4��q�Y�{w�{�Nt�^j<̻��;;o}��tӒ�N	�mN�M��G'B:���9Z�8c�ih���ΝNh��t��Prښ��^��C�����E�l
��ux�n�i��8�� k��%��_d좭���U�\
R�
��)u���e�ؗd���T|i��w�Uͨ���l)�Y)��q�����֋\�O��cE֎����*�S�sׅf��Z9e)DQ�0�Ws
3{���w�	1�S��]���v�ۦ���h�,<��]�����(m%m>�1-v��X#՜
��9�2��v:��B2B���;�9�0�.�/Z|;+�d�b�v^u�;]��$�6��D�ɠ���p�E���N�S&Е�oj�[����jٯ#���Y���p>��;�ө��L�K)â�a��}�yؾ,u�#�8,��EA�5�f����-"�����lzn��)ջ�,�_)�:����л<Rbޣ��_Y�cv�D��y�-m�5as�Νb2+�ʰ����W�i���<�zyD�>�v	3ٹ��tF�2���#I�YH��F4�G��&��N����)������y`
Pnpr[X\����Pz�*�z8�O�ڡ|�EW�6���G��n��2����/�qd�+���i�f�S�pσ�lit���g�W[��8�2v}�)@�e<��}�Cx���\���Db�֋JPο�͍�K��TB%�T��]��E���wל�n���J��o����S�ٮ�Af����1�/��%^U�ގ�b4�1�7�Jop[��S�����tm�(������Ϯɗ}��Q��Q;ekr��+�]�u��vQ�l�r���0N�ꃍY�5絸0#G�k��wڱm�LH;Y4����j���������}ᙖr���<����ă���Tޕ5�d��oA]�2jb�[�@��� ��u�5��r�r�Tn>͠�jMY�k���3h�f�6��q�3���:��qľ�:;��CFhE�k�mw$s�|���"�%��|�����k��F���EaV���f�f]d��5��������|���2���ŇxQ�v���qޜ5��/J�jv�c���Ʃ���3c}�-�b��M�ǶZ��I�V�]�������ԃ����7�H�F�*Qu]ۻ��K�5��o!z����R�����.���<vp/$�S�=�
�*�M6ū�$3�����lD��Y����nk�L�Q�X�f���N2n@�͢x+�yX^+����NKP��=O��do���
�U�������[Xl(ܙ���N�U��Y��k�%b@e
��!��2�m$Ƥ���.L�DEϱ��_]����X�`��ȵPV�P��I�]�F��h Z�b���Y�a�2|��S�f[t=V�*� �Oǅ�5ٝI� ��w��z{T5Ld.5��fk)^s�"���|�j�L7�8V!!�ӕg�Pk1汋^&�����5pm�jؚ�X�n�`�K�I7�"�
�f�wN���o�p�c�Ӻ�����<QV��g��=�-DV�]yh��f�����{]��N�nVT��:T��NW���{��v��	��vkL�@��v���J�r�L",y�9t�S.�F���b��M2u%a(8��U�����ٹ�nf�J�.�L�"cA����
�_9}lS��\�6�ar�>��S_+�}gs�u��"'sH���`jԄ�KQ{"f�B^N��]�]���(�ڗ`P�-PDu��r��i�����u�8 �&.8I���:�]Z��U`�x!�Ū��jv�@��+J�V֋1����KxU])D��F�_S��ɓ��A��'!!�ʼp���R�V ��Z��S^�S��0�U��h�i͵v�鹋;��-����Jq掿�[��ѫ|�!g�;;�sb̊����fp��	��]:���fB��E8�zh�5�"��!�z�t�ɣ\��M�4^ʈ�	����f�{��sr�y�������y������bSJ\�tTē�R�/q�p9[t�.�b����<{��?b�҇��/CV{)��A�s��x�}(V�ɱ\��A�����[�`��}�+7��:zu�85�ǃ[��,;�D�BՖ,��D��EG�U�^gWEGC�6�k)c�e�a���@b��ǆ��q��k�v�����Y�Lopmwc6&�w��wL�ׁRe�3
�r��\SڋH8�f�=�lRP-��"�n������=n%+^�b����-ѡWzk�kI��y�`���4�W<V�܎�1�H��/���{�G���ѨuZ���o���wq|��9�(��f�q�}S�����ot�2^�.=���J�2j���/��Wot�t�Paj�WU�p�3��:���~�:�V��Z�*������td�@6��7��oy�Á��[Z�s8�Uz���Q\Uq��Q� �*�m>T��_�z�0�,�2�5��=���g�`Ҏ�3霴^m��grN���-FĵE��XT�vk���*k�#n�K�2L��I}+^�)��a�T�K��S问vAG Z,��W\�Y3`SLJ���*My���+��7�A�ndz�㜵��ĺu�"�V<��/El�n�v�7���s�t�ƶ��V("�.��vݥ�
�_ﲖ�ĮTF���Ը��P�s&f^MfD�]��nB�*O-�^�A�A+����f�g9z컗 ��fwSb���ӌ���e\wvfM:]�O'E�d�U���z�8�j��-�o���w�cܢ�Ӵ�yXp�������|�
�X0�N4\I�>쬣zC������3$�͘%^�D����NV�f[j E`�Sw���@U�}6 ޮ��rE������D��VZ���>�`s9|�K�����Y�sQ�M_;�=t�+9X�����/����mR��:�s����G��l�E"�7��mwL�}j�g��z�"�Sa������F�y��3���Vr)��Eͽ�&;ҊWIR�`��D���X2ċsU��������X���X��|�̼A����.к�{q��N�Y�g(�n���؛�jn�=|�}�5,��㲻' �څVS�s�����_`���mt躵�+�^`t�$sz�z�w�Ռu�͓D���<�����v�Ƣ�*bS���W�T��G"0�EB�����W�]f���sC�l͝y��]�Jv�H�R�{���I���1yp���ͼq-51����ِ!���胸��o!�x>=�`�kR���D�[˲�#/-"B]+��a|��/��Tу-uՇ/q@�4��v>-�v�����tɭ5���}�RS�˧����૤KM�`�S�j৐pfeK�	4�)^2������9������7}}q�\_vV�]�[��[N�]}�^B��#��(Y�y�C����XY�s����_��5����+��^˵8��Sw��X֎���Κ��L��Q���X��*w:��]k�قc&��˄}V��olY�v�g'k|�`̥�	�m�h�l�W�;�RwR�b����_�-�����]D���2C]�6nb��2�v���|3/Z<��rRk%Nrw_�tw+h��֓wr�w9�(����}�n�g��p�P�N���m�2�;9Dah�6��B�i}�3d=��#ʀ�3�t�U݉�˜V����|�<�+t^�l���d1�w>$��}4WV.�|7U;�VU�n��r5ͭ�Ș��m��i<�]=���G8Tx��Om�#����
Сɜۇ6��ί�����v����������1����6�8l��ee�ɧ-�E�ScVۃw��r�ä���&�ed#ny�� ��Ỹ�q7��@��kE�Ǥg4/�2�EsV�Z�1��N7�oVP�j���	�U���0ʿ�������g���f��oo���oT�85��U�y1�y�*K�����f�أJ�AUy�&^]�z����K$��"�*�nm)��nN[��Qr�[cY4�����E66:�]�L�kngK+t��e��t�\.����3q�������qT�!��ƅ1g����#�2��JaQ���h�$���|�u���Pse�n����*��³ �⵱��'t�5���5����lɘ�)"G\E����&�1��v�wa͊��	�fp�$��ٕ�t���T	
"��4��ʺ��P���L�K=̇%t�9�T�Q�>�~�5sֽyL[���n�;��.'�Ȋ�S�Ȳ���`/��|��5o]E�5'��q*Ȣ�]�;��q��z���=l����u��kSC|�ܗk�AG{�{�F��*�5�eݞa [�y-����l�:ۮ�]�{B����{�mGj�q�E��v
2�I���N��#Ċ|��މ�φ;�t�H�k��|kv���H����o@[����.[�;���`^r�C	�-�X��wN\���֤-3ݲ��}K�]7p�6x�P�m�oO�:ѥNDd/.�[���!�]����v�Z�ŧ����o�	7��u��/Sź:�x��LD�Qx�T�1c�MjU�s���B�攝�%��jҡ��I�c�J����n�YcUJ���5z��dU�yO�i�Į�k���Z���N��*r��좗H�溒k��g^��s�ţ,�+��0g*'���SX��N�vμ�v#��q�Δl4n�vu���+���L����
�ukk��{��K�%Y�|Z�o�@�����������P5]�2���=bֽ�(u�s�s8��_S��nM[�)ȝqW���� ]#HgZq�X;W�$k3Gϒ	���lUqׯ��*�^^@�Z꘥&.q���3�C���eW���*��43��PVc���f9�nㅺA�F}ӫ��� ��v��[��K6�۔�K�{���aG����]�\��AԴad��cR��w2���l��o��hm�܁����hʍ��l��ܖ	I�p�N"��vEt�1�^4�Y�^ZY�`�n�����g��V�yt�ƫ�nV.��R�}�ԕ��;7ᴞC2��%���J�ߐ�:��Q�"��(e�.�ϧiQ�� ����W���u������K�����#�@�'R��d`f �)���o�{�\z	{:4����𭸱\���kk"��ۆ���wꡋAWJ}�=��$C9l8,qL�r�;��}v�5�hdj�getW�m�e�t��ep�����M�@v�T\\{8f�I[�c��-��1�DB4�V�:�m�� �l�.�/.WPnU��XG4\�Y
��l��z�W
�5ݕ�fmܼ�Sa�0j̷p��+F�j-R����[��U��SZiڮ	�<8�
�	՗�������|���h4�Y7��/z���
�=��u��1��[��1���0�nN�%n����)�ul�%n
�єH�[I�+��wp��܎`F�z	wY�Ҽ��Au K;YT�`������L̜�c��rC�K�se�5����}f��p����%qˀz��Ƴ��b�]ȼ���9��\�z��������4�a�[�;�%X���HQmp|��7κ��5X��c��*�X��Sy�j���m��ەZ�k�-C�t.�J5ݩ��k�̓�"s-w$(�&x�6J���.=����Ө�x��h�8�7cW�kor�{�w_S#X4�h/��&.V6�kk��rEV�s!q ��b���s�x�7�e�핲�`l���x�"���V�-3���6��+�;�b��*W*㦰�qk{^�9d��6��,U}dgF�a%�Kʹz�g
@3+/�	 �kt�B��wkEռ�{����a;|c��.W]�9c[I�#�����)*��h�T�Y�l�fXM� �He�u��X���D R���l�D�y�m���:o��D��*{�]Kܔ(<�@؊��_��r����:�Z8��9=����s��op���)�k_]�%�sq�wv�\"��� �z�%�\�s�cta�]�4��V���Z�����!�M>�·;�!�z-S���o(,����$3��:�Y�J�u��F�y"��]Z�u�*��7��c��s	��1��� �.��0R�8gW^��YM�gG.��/�.7�qr���[��@�Wx{��KGs��̓�\�tk+y��<��uG#�����m�4�&AJ��֓+��y��:Mi<�oL�H�|��ķ'fL�$m��6�u�� n&��N��9��b�P�$����6n�'�X�-�6��Ɍ�!�4!�M����s���^\�Jom��3[}�ABݎ��l�s����fVw_4���r�u�
�z��B�G�[�<�L��;쬴���;�����d*�fDo@�!ʵ�]fS�����SwW�$��`{70+�۩Ywa�P��bj����g]��d������NUp�;M�KIn.��]9��vĶ�p�}�%�w'v��7,%5�P2�RZ��iZ���n����4f�7{����b�Y�ۏ�����.�����J�7M�@�����wv��m4�dpoS6�"͆��[b��d�.E�w���AnE�`�ٷ;tW�e���1�Dj�v�W	�N�����v�&.�[ʖ�ޢ�ej؄���=���C�fc���e�KvR���a�]�bTN�5����nȭS� ;���oO��S}��q�*BEf`éf�oN�䓿K��]�AI�e�=�q�k�ʚ'PO��u*T�2Ү˗�����7��+�p�X]ϟ=v(�j^�[�!m�k/ f;f֮ť������'v�g�;yٝz��ڛ�&��:�5/$|�(�!*��լu�t�4Iv��b�S,u�����ݢ�@gU���t��p��c��ǽ����r���ٖ���ua+�j���n�6�No�H�<�*s����5��69�]�S������������M�{��G�   }����������:I�>��83p*�P�4bp��E*W4<mDr*ݥ��j&脒�x�X+ S-)-�o���-,:�<�;G6��nd�jl��\խ�ަn��DZAt����ڝ���:2r�Y3�n�m�x鉡3
-�`�������6��ua ��Ն�qv��M��;R��X�8��ź=�!��W`�,�J�#9n��v1u��]u���6*⭅��d�%L=9r���.�r�,o�.ؔ���l����u�Ԭ�*ڸ�+(�x�x� 9\��Rha��ҭ��h����xY��l�C&���<���h��i:R7$V��hH�ˉk��˹M�o��vayN�7g�q�zO��Lh�cZ���������������<O!:���om0���f��f��ggS�����vYK�3Rh��� ��di�V�\(ڡ{<ŝ������xۥdغLvQ�i��M;Vĺv:VU&Vz(�:�f��֎�_=s���$}�Nm�X�L�x���A"���|�
b���n���G0<�Ul�i�T�T�Z=53j���Y�b�q,t�B88~#����%U9 �M�^m�m	o�wI�T|�u�K��ğbˣa�c��u�WT�+4�]�6�
",k���s���Z{n٢�D9<n�]2j�"�5��z9Qծ�]��B'e=Fi��ݺ���9�bL��h�f�`Xx��R���	/)䳁��%�A�N��b�,�#�9�K+zS��|WY2�`�n�ݹxn�,���}�nc��¬8���UP.���#\����g��u(�:n�Gp��V�Go[X��h�[V�c�Z��ٹM��a���1:A\Wd���I*7P�Uڕ��Z[����6�����J�Ø�C��I���f�ǂWź��%LV�fq#*,a�|(�o[�%T��kJ2���&G�o�D=����V����	��`�T�{�o8W$�R�E��ح��d�t�r{�_eZUL�Z.�]&��=��-V-
DO<]�4s���IKfgu̬��R�&��]�Xf�0�}��+����6�"��Ǝ����>G�ؖX��J�սяMre��R�S,|��J�jK�9!X����1���K)ے��A䡴歷�����}}��,�G�l���do 7J��}k��K�^�Y��9���l�ʊ'흢�����Ѱ6�x�(�ji��+r�4�$����m�T%iA(bSe�e�̶
�ʣN�lLN�f��M��RZw��\���kDeиkPȻX����N�Pj�T�7���-#yw�`-`��p�Ɂ!@�5`�q�R(��ó7��X��C͹#��N�H���B�h�j�˪��_>����k�>��/�h�M�Ur�!+yYe�Yj�z��;���EL����+S���g���ݗְ�{������#i�`�v:x�e�VI�y{C���C]	���J!��#5��\Lݽl��.��gf��i���h��c��	�Le�`͡�jF���7��H�$ݪwoHup���c��
�7�9�t6�Q��É�#�a�$��� 2f�b�W�4=�!VQ�w8�;�"��q>���Ru|N������=��@lgA٫^����E8ù��9@�� ;Otaz��/	tu���i�'�]���P�t�vV���㥗Cp�;Hn1k���j�R�(A��3�8ִ�
ڧ�6_U����ÊvչL��O��Cu%}�+6%�f�f � ��)^�G�$냂4љ{�j�e9da��-���`vZzs��i5C3����HE��u�!�4�de��
���%��gm�'�eK�r�'We��AR��y�����=�R�V@M��ń��"�D�	6�Y�J�ݴa��]��X�r���*���co;�(1�����{��te���D�����o�`�+A��N�YmL���)�Y!Nq{��7R�s����a�n�Y��r-��h5�l�aR�2M�Ah�4��-Ɗ�MĬ��g���A��v�VG��Lv �ej�tf��	X�]Nvp��o|���)o�7/;d8ī�ŕd�k%]@�zd���-���o���s�>+��{�b ^n��̈J�\� v4C�������ve����:�3NhT�+i��T�5,�x�5zDCj���W+�E��jv�.�]��j<T&\qP��4f1:,`�x��@�
N[C�3v_vt̃r��d9D���L�&��|�6S#�aMܚ�g+��ҷa�f�V��GH�]!h�o;�����g B�Ґ���k�9Sܬ�K���Y�*����Kw.�ט��x+��ss�m���[]Y@�����Jp���.����K��H�e�{@<i��d������|l�����6Y1"(9&e�]���6Y1uB�Ɵ�Fq����~b]tL�uT��z6��M��dւ����<Q��#�6pR��[���U�ݧ�u��GU���H0���]H8�i���ΧP3��n�k�Q��7G�+�i��62�_][�#곺�v
�j��}�`�)�f�sg+���:c ���u�e�[���j��h"˄�9I�&���v�i�5м�3:�5t�i�^�p�iq��1�v:�-d��N��&��9��	R�a�FM����3	f�
٪Z��쓶	��L��}pPAj�o3f�����Ը��o�U��:d4z�\0vX����ĺa��z����ev@�=_5��ڼt��͊����|���ʼ��S��N��#�EkujB��JWW��E�pӸ��z+ GS�h���8[��"���{W�+K�\0>ح�/@�ͦz*��U��8�V��Uy��Wo�|��tɡ�Ϭ��`�	(%��_j�ǝMfMS
��s�ח�[�ԧ��1���^p@��]�!�����U�u�B�z�rlT��w���d���L�޷$��*6*��b�7Gs��.��X��7�cP�wk:����6� +1'��t�A��oh�ŻwK�ۻ����3mpA���^kT����	�<���{�z]<,+(D+���� rF�Y�!���HQ�5��K܂a�Kr\EХ��h�-��;�Lʼ�-�G����\���i&�^S�3)R8ɫG�n�uyMӬӯyw3���F��|5���� ��:MFX*J��x��J͕�Ki�IQ��
7��,Z�s*�\tc�#�v��+׌�il\c���R�T�nC��hS.l7V��`�j�]�"��Ry�3�l]�3��u��o�l*��&�v�P}�P�\*<Uw�9.�j��&��([L(-�*rEm�EQۺ��n� �w�-���K�m^� �Ё�n4AWg]� �+D�H��:� ���¹]ڗ���G
��F����l�e�/s��b�`S7�MdF5R�	3m
ѧ��Wu��[	9�:���Aݖ��&�rɋ. ;V�� n�X��-�eS��]�M���PAIX�1:9�����%�͓�����e�S�:�:Z�윙yz�	�:7��a����U��Vb6�,����%x&�
���J���W�Wf�*(�Ҝ�Kz�o��i1I3QbP�y�ZUv-���-�]�.ԍh���E��kaL3d�`�0� ��3�Vqۃ2��u�}̈*�5>��7�R���m
\%gfR:�ip3y,��k,�!�w7˼�VP��#`����i�LS@47@ụ#ǍAU�ԩ�J��4��v�o-�_9�C+D�U�Z��9��E+��X��w�*�B��E�X��2�4�m�xE!��I���bޕ�B�{@�y�`�4�3@��]�jp���(���5jQ�=�@Y������{&X����N��1;��n�9qo*�]f���ʷ5A���v��f}���k8s�O@�"�)g%�o���S���I�r�Yr��FT�O�RJՓbL�hhrem㩻	�kH"��ٔ�m�O&`O��:�Y�=�@����"���˩������v9J�͍` /) �s�]�y�LgN���r(6��KV�[}�̌0�Y*�8����C��W�|݁X@��Ѵ��t�<iز�R�G��x��#7tF#���i	�<Ӄف��g
���K�b�]%\0#���ֺ��al��^�(I%r�f1�Ħ��*W�X�\n)q�wgKXJ�ët'w�i��ujK/y�(J�����Nӈ@{{wY��̽��4�x�w�^R�s�5�	�]|�;v��t�n�`� �h�����-[Pb����<��}���1��V& �"�Z��Dn��%ΆP �W��ܵVq��ma�L��Cy�1VGSJ+Y�����������i��A�����I�LD�a��ŷGj.�f���� 85�� s��;6[��r5�J�7�!��)1��ژo���5s��'����������ݾ[�ۮ%k8��ՓG��s�T������[�]YP����?)t�6�� E9m$*#���r�SR��p��v��"kzP���Q�g7������y���0Y���݃����q!��a`�A�f�mH*`H�&�IJ$�@Yxɜ�n$E�"s��쫆ۼ&���GDXo	YN[)]��-��y&d;��H�z�*õ�и��6�:	�r
�I
�j�F��f��,Q�'k�NؕŌ�HW"�ީ�K���!�����u�kY�]�� ��̠Xvp�x�j�J��,ص���I�7�U�n�	�<�g&�N��&W!K!�����n,�6Y+Wr$��e�������@���Ӥ�19��*���Nm`�����������ڴ++�[]E��1�b��qs@TV�v7:���<Z�vu �V�J��n�cKkP�6�j����:�M<����� n��� q�܎����Va��.��WM�XQ&M�*����s釫Qdk�}�Rk���T�-��p|5U���\�lA�"��jv�F935غ��ɊpU�bZ�{�Y�M����M)S۩�:w��Y: �9۴�E �fSr�1[��ǗI�t�l�y��wJH彡*N�ݑ�'��wa]Ȇ�Dɱ�np9Q��`J���zHH�-	KU:*��8'�n�jz�(��wt-�w
�K�i��uo��2�:����v��K.� �`���N��Zr�Xlwu+�7V�����4U��}��Q�(�[Nm�1#52��ܴ]g}������r��d�뾍�wv�=;�܊=R�J��<��{��f�[;i�7t�:�Hq'�<ݭ!�Ư����V�Cc���!�`"�{%��1	Ctfm�ؔ{h�YwMp�K��7/����u����TCR�Wd�%��Pd(�ia���3[y�T�mj7��m��mQ���ڰhR*�N�CE-9Ճ�V,�C��Wܯ]��-(���ǁ[Ӷ����k�x��/�:q��!ClI�ݘ/�ڋ�N�t�+R���w���Ґ���z���:����̻�i��u�l|���]�^�Ci�2�g�-�A��cXj��AGL
݈�azjiڡmZ�Č�1B;fV#0�"�nq�N�6�SqG�i�0S��H��h:7nG�:$CbӁl���|�um��P]\�W����m �Pm%�f��g���j�R����hڱ��}f��'��d��,�G]�#6 "H�B�ܸm�
9�t#r�pҵ42̎(�s��ҝ�|���Z�+U�*�3*Խ�YZ4���B�
h@>�C�Y��PX��GEZ�q���ht�3��(��k�af���-���U`c�xm����:~�v*V=e��Ǎ-(�Ŕ.�K����V.����Ϲo]q{/5N��
��F�&�ވb
D��ب��+����Cv�DT��er�ܨ����;�=��>�����;��]7�(��?XD�ұ�ݕ�oX�wPو�Z
c)�J���.�
�Znޢ�`�vVV��ݼ�:�%3�3�Oǝ5�Zd-)v���ԊV�Z�J��l�r�w{��Μ�<��X�Ӣ��_��+6���}h����ՍL%�L�%�1��ݘ��U�ɺ,^�n-V�[���|5��S���]�F�R�e5�Z.$.�iR㮮cG%�����dZle\{ԟ#���|��	�;1�����c�w6�6F�ܴ�Xm�61G]��u���J�omX�W��.�efW 1WjNv��f�ɘd�.��B�v�21��)��7�}[�wg0ܐR�[��3V�oZa���Qug����@-yћ�i\"eB����dI�p���2�����B��|�<4�����Y$�B� g��v�lU�sz������{������h���WA�<y7u:Vp4����ŉ�s(P�s^������Jܔ�j�Z�����ªYzՉj�J��c����'���=I]¤�l+��b�,��ʶ��X���Ӷ>(�E[f��#�b���]�Go+lWa�;Bi8��Z�m�����V�^r����I2�D����A��M[�χ->;}mY7����6� �����m�0�缪�n�/��e�6�5��r}%u�#��
+hU��Ƥ먓�ƕG�U6U�CfȜ��Q��BlU��Z�N�:��ɥ��Pl�g���V*�^�-儌�����˚�|�q���R�peu^���Su�Tn��TM��M �^GBJ	��ml�xY�m� b:,U�ӕ�P5�t�8�ݳ�(�\�c�)}���;eR��c����;ВT5�R�}%�ڱ����m�΍�J��px;Q]�aHd�]m
_;�}�}_W���������s����&���!���o$��4h��g ���fv��C��@(*y5�pn�F�t��ý�����m[w�]��hw`��rח�������5Q ���Hf8Տ�n���fdł�A�f�P/�;�"��K�S5w�Q�Ճ/1��w_��دK|h���lB����2�ȩ���u[�o Tcp�{G�!YJ9ٕf]fG�+w"��"���OF�7M� {w��ܫ�o261��K�MN�_t�ѴdKANԽw�ѥ��[X1�-�8J�K��3�uanto�]wz����B�>���[.��7hv��^�=� ��ү�4���O+�(��[P����EZo(�:�Oe��kj�gaj���:�w�NNQM�en���W�e��X�[Ȑ�9�Q��@�fZ�Ɨt&���
�6�;�M��[�tQG`�h�aR�����m���Ȯp����L9�V�(yvh��/��!�&�p�ܸ������f�9���X��rqZc[l%09����gc���KrQ�3x(���Ξ+'�>�*��ȴ\YI��q�&\��#�L�Yv��N����L΍���4�YA��Ѥ�����7	W�K���li"I�
ȆL��Q�/FeN��4��£���j�uM���!�V76���os��Ņ�D�Ml˅ޑ&;��ub�9֜��>��� ���e�!YRf�L$$H��C!!%F!bLeL,��qĹ�1D�)	6$���ɢiF�!R�I����a��M�S4T��dhdF"!	2f��%�ѰT�Lh�$�H��"LH��ĕ#J-D�f30,b"(�4�s��!X��9r��$��)�RY6%�2R(&��F�fR�D�#	4�6�� ��d�22Q��d�s���E4	H79�����,�"#����4���P�!d��"b�`҉$�����Q��J��R[&1f"J-4�Ib�%F1%�!�DŔ���*4��`��D2A�����a2hL�	 ��L�j(+I�F"H�h�#�M�fgI�����F*4[6L!�F %'�ݸvO>���}���j�!�t6���2�R�B뻩�98�I��D�s�cs��\]�k`v.����� x\�.���bn	�N��;��+�v�tV|9�f|�p���h���+wRBi�B��,�����gFT��/--K���6١�f��u�z���,z޼�)���pT
�<7]��#S�kd���EP������
���3�bRQ�
Ќ\6�v�Z5[��au�[�*(�m��'�=�z�(�jL�1G��e��z���5��:^9Ǩ�0=>�������*�9�y�K*��%�'�,	��(UT��S���}���꧌b�0P��*�9}-k�2�;ʉ��4�*8@�9
�t�p"ǀ��45��t<�_��?�MƿV��t�СY����Ju�%�dX��'2|W���|x--��6 �D	�U��g���lzر���>Y��kW+�>�˸����O�v�����.�Ȝz�5�<�.^R�z��SR�^�^ϴ-b�L��T�z!eh����	9�`
���O�CE:G�x�������񾦻Ԕ��=�'��N�����%�8S>e�O��iIL�!�A�[уat��A�p�� U�;s�}`l|��5��C+�1f�G0�	�vgn����Z���,��&o� �'v��Չ��7���oR������sP[v���;.���c��N2�t�GIY6h�Wc��YX͙�h�RH/�%��'-�o4�z�2��aU���"ǅ���s��#ߧGިn������]D�\8fw�ݱX[/o3�m4��4�
��w��³o�wl��
���7[�ߛ�:o�4��%�š6�	5�ᮆl#�0p�=�$�� #��7* C#SV�w:� Ǉ��V0�6]�ÁV��ʗ��˰;��g�aA�������c=�2��[ym�:I�Bp�R7itq�*���Yo�V���u���X��Lө�B�0�pVSu/NQ�+��V���=�^>���bU)�L�)�f����|�������m��=�p
bk���{Wwk��y�4�s��:(����n\��k��Di��酖�C��]}�ػU�-�ץ���C��,��^<=&����q�[�@�qXs��G��xNpU�q}cv�w��澂�AH�(GC��[jFŁ�t�3�����)Y�e��x��=~s{�2�|���>������{�"���o�ث�}��9�^� w ��m��+�g�8���X�R�,�4/�V1��Cv�um���G�EW��{��Wsp�xt\h,��l��J�����mwU�\ 8�V�e�վcpN%ܐ+#>Z:��j9�G�aI�ʂڜ��l�gT7ZgTǼ�8t�ƌ��j�K]3��{.���eyk�\!0KK���֯%�
�aڳ�7�P��W��7Tfz��k�d)����b3'��\��v΋�h�89A,^�I�������O\�����Ǩ�x��Puˣi�e{�j�˅1zS(D���A�2����&��ڍ�Ӳ�DE��SR�Ϣ-MW��yÔ,04��ڸ{�5���TY9�p�͊syx:��D�=� U@ߏүN�x����©c���ы�9��cA�١2�}���L�=S��R�\[� ����(*=���s�����N|��4R���[hy Z��Sz����/� X�(K����  ����E��6U�t�C�K��>���r.�ܭٺ����.q`����Q���TQuʑ<�{T�@�7�E:G��^/�>¼�Le1i�s��_�X0���>��4C�m�� ��42UD�$��oM���\�8���q�}}�Jz��D�C�d �qC/��������G�= >�(Pޘ���s[���&�Trh��R���Ľ��P�����s��7@�=�|��e5�n�KK�N�s�H����^��?�C1K�Mp�{Ye$̉�b
�qh�V�\6���yg�u\��s���j�V �����gR�z��,�ڲ���k�ƃ���w��ʃf�����=?n;�������l��g�)�{�|4����WnGFU��D`u��h�?e.We������G	��HX�3L||���4V�C3׃B���*�����	���ѻCe�3h�t�P�Qg�^��,쨵�N��~����y���/Ω����1"�˨�{����M+5�9�l�e@�u�p��3W�w U·<R��@<^��}t�>#�Q5�e��N:~��'��D*�f;����py��}��.ǣ��|*�o�xs���M������;�Ѻ���ur���(�r,��<<�1U�#����{�® ���Yb�*u��"���Co,s쌦�9
=�5Zh@��韌�1q2��)yU�v���u�^�_���4�jH�=�3���ߣ:��<}�I:�����k�=��ixo���~�V��J�o�=�T�廦�U�Ÿ��(bu��rU�@�����<;�����t�P��յ%�T��q�eu��#�\�=�Z�AK��%`�r}`�Q�����ǋ[�zl�]��_N]��]J�N�L�Cc��>F�`��4v�����}[��;�b����A�L�z-sVQj��݉��Ε�qSV��� ��e_(yo%��&[�ο#50���{$F[tE�S�Ex9���*�d��U ��^��hz���j��d�F�w�3L��U�1=��Cj笿���S��ҵ��P�m�=@
�h��\���gf�)���LJ|����l|�jv�-�,���MCn���6�*����qc8�f�c�T����LfW�1 �8��+MG�Q��B��7:KC��g�ӫ����r�j[Ko��Q�9��֨����O��j�v�e
��*�N��=j��N��[��t/YK�FgPվ�:o%��}�3C,��1���P>p?�<7�[5�kG1��W��V��޽u~�Wo�M��"�Wx^�ѱ�
�}�6.Vy�J +F�l���b=gu�څj.=�� h��w��K�O�Uv����>Լw���U�+<�5o�^!O��Ve�Cݛ��m��f�K�ɹk�w��k�v>��������ue�B�3,�òB�-?+��r2�cGۅ�U�x�9`Í�b�k ������ӌo/��s����ד�[­�3�k�W&ļ��	4���v�\u`s��+]ea�9!�Z4H���m;;-d�R�Zr�q��n�H@~w��|��ޣ��l�6Ж��q�hv��y���ce� n_st���s���V9}S]̥װ�����U��j�Z}�<#�5��U���^���2ewE���{�<B�����pX�5�)��2�*<PsUksC�zܮ!�F4�f��e������1���}��c8I�ct�8�0;4F�_,�a^��Xܜ���&��$=��Ϊpg��n�-S蕗��Z�hԪgA']%�!�uҚCEޙ�p#<�!k�CT�P�/�1(�{]�>�rx}~C*WZ��.0ؔV��A>�#��qG/YN��-�}`���T�|z���bƿ:�/\�;��na�LeԲ��/V��5
��U�4�� ӽ��<)Um��b|��}(t�ї^�� ����n����n��Ꞿ����)��@��	��
�&<��0�r�3SV���k1�ck*rVy���x��y�'ݚ�ӥ A6����0��y�3�{Ne��������>�
�<.ZcV���^�0�����ݰg7<�O��]_���i�{� �����U���m���Y����v�AƩL�6��5��k ��q��:���)�<O����B\��=,d�������(������:WT	o*��6�w��N�J}��ا�S���`ב����iR2��*j�+uL�}�
jݎ/��6��΃k��+y� K�CVu��|�(��:��9h#��jiZ��Gy�Z��Z��;��VN�zidc\(וwx�~�ϔ�n\���eƺ@���s��N�������hj�"C����5������6�%}���]�@!�O*�rW�)��=0k�ʽ�՘�=>�@�b����^F���[���G\&����;}=�4D���e���>���u�{�k��u:P�M�w@�=k��ԇ
Nq;)W M���dU����s��Yo˛F��֣�w�ˣ���f�yk�]d��bgY_�2�%f� vv��"��,/�qMiK	�`"�1ֲ=
��2W/
̕ޕ���3�~����:	`�$A���u���9&3;9f�����p�r62��!�OF�����k�9T�뼸R��u؝/����}Ϥ��=G׃}J���`iy��|���u:hB�号�!��G�ڸ{�SX��O�k�J<�{ں'{oP�F��t����\$�o����19��ԽƮ<�3�3^줩Q��G�.ˉ[4��ލ-�0d�:��cSƄ|3d"�Oǹ�ϗq������JqwJЖ���aP��6�_e����Ԙ�A��=y�\v'RGa�g�׿]�#�P���#M�	0={��:�v�q���@����c��2�(v�����]�-������N�n��,�	U��=�'����3��������Ũ%�I[�U\���N��o4��b��}"!Ò����6� !?��@��Jgk�WiK݃�v'3���G�x�x�y'��֜{����r�H$�1�N������3kľV�}Ƕtx3���F�{�Q�m���s6�W^/ �)��y�H=H�Ц���oM`\��t�Ҕ���\L!�L���8&L(�I�g��G���x�
�둭�l%⩇��R���G���`����D�~4!�㿘���E��k����t@�u�'�X©�߲������Fl�zPd|<	G]y�o����.�|૞=-��K.�/k#�<�Ҹ
:nhoJ���L}0N(5~��ok���t��������#[Vi*kg|�o��e`p&K�\y�tM�{��Ba� ��{�.6\͟��0_'ȏ���J/���G����k�)Y�!��5���OS�:qc\�]VgZ�nf(5u�ӱ)��~?���r��ڦWc����4/��x�|\5�*��k<l-<��Q)`U�U�R�:����xmsc^����*��ݻ��g=��lp53�SWlAN�Xm�/�]�k�Y?1ˍBc(�ֲl�� 2��d8T����� v0]�'_1C���(��$���:��=r����ֺf�*!/�[G��%�C�������*τ|����8��Zc�xU��:��r��}N�=j��R��E���oAF�32?(
�?v�V���1����c�_�}�b�ԫ��	xoqP=�ǼW�����уڶZ�@���'h��C�
AH�詖5@�m��v˴:��C����(/�'�@,76��C���a�+>R �5'@�����a"�?h�0���"�R�A#�s5��=q;+��/LOO�E������#O?�1} ��2(Cr���R�ܞO&����f@��㘖��o%�LǄ;sr����UT�=^�ݻ�&�q��9�׊�/||
�4/�sz����Q��x���o �����4'��0�G�r��N���u?}�?39"=҂��E�=���\Dnm�����7:K��)�.�|�<���.���@qLw>qk���Q>�>;:]�B�"��\)Vg�p��_eZ�f2�Wc����W�\E�,��T]��3��;P~�1eG5���Gl�<m�-�pE\�0`��3��m�>�b����V�� }6{_��z���y����Д!�t�%o�m)V�?�<���c�ܔ�9��qZ�ȭ�^��쮣\ki-SY�Ճ����� ��2�� G ;�S��}�����E��ƺ�=vP�����LΨ�PF١q���r�c@��uB�g�Ĥ> V���k�5۬�ޭe�Q^Im��x��{��w��.}_^H�"���_b]�1�B��|`�����PYЯҸ��:T�(6SW��>��K�;!>�6ԓ��7�qc�W��M�[6����H`�Ђ۳�yu-�����@]�Z ���Ӊُ����8�f���׷i��O4���ے*^g�eWt<u���t^�~��ۢ��������mZ��� ����+��w�q~�>���}پ�����=2��>�tln�ZI����4k�6���\|޸�����
2kί#���U_x��v��fRǶ%e�Z�hč�ɜCڄ�N�~�4(�V�R֬S����C�2��u��t����eCj�S>e���$.U!��a���{w�N���{ʣJ��ժ�j
E��5㴎k��n=:>�sC�Q�E�܊�r@g�N�@�Ftx ���jwT
����R������"�r�&>�|����I�=0���=�"�8�M��6��,�x��H7�ݧoA�ž�*��#p_]��U:�H��Ts*mčҷD7��XUH�wcK�.Y��Z��t��p����n��
̩FwN�uS���MZ�`rz��;{ ���+>#Vڭ�9�9�ސ{؈��\9��.F|-by�%_ ը���\�2w<ٙ�,�a�KRY�3\���K	���V[��X�Sk*R����x�N\`���we�e0��}�gb�.f0a�,]�J�v��]6�E�E�,� s�m�5�\p�Wn��!�h�M�o/q�o8�J��@A8�7�H�Z�I��f�yj�Ѐ:�*,�ien��7�2��}�����n�|�]O�&��L�S��&
���J�3��Y�	v�2밖h��\��:9V6v�e����F������>��"�+�]���Pڀ��u
�4�T�X�}c�K��:n�d�\,Z(^���M�-��\Ug	`�j>���� �ʋ�ҷC��ҵ>�+b�۽@�[Ȣ��)�,1����{H��Pv�ui��q��4C&7'#�^o|��U��.�3��o��LN�K�J�y�ؽ�xS�|��ʂ�0z�WH�;�L�F�ล]1.��y7��Q�(�C���B�u��0^����+��k��5�aE\�y#o���d�Z�KO�w�������
ȕ�Hni�-��3htk��шb��U��n�at(��LHz6C����t]a�ob�ט��-�1"��p�n�Wt�w3�O�j�d�v�
ʔT2͆����hٵ�.�O�M`����+(�,������w��uS��Xzx^ҷ�IX��Ɩ۾g-K;�`yl��`'2�s�`%f�]U�i�`�a��q�9w,:šv���@ഩp����{g!���g=�Y��j��W����m�q=�Tl�}h�p�� ��%����U���6v|F���݇;F�[\vH�1Bދ駆!������b�t��7��|��0:&"ugDɄ�1�&��>[�������:���Ewb�׶Y������	��+;�쬹�)�l���r��dp����V�<�9��U��Wb�<�9X���1������u��h;Z�$��� ܫSt��k�83��}ܤq��P�9�[�Yk!����q���:�:bu4�9Op4�!ykm5����d�����0EsG!	G��n	l��ޕ����r���(JZ;�eS��&��of�gUF���j��L(�,Q��ǚf/���q���������t�X�k�FRS����6��q���8؋�g��M���]��i�˵*!�	ī�7���-�W�R5��JPU���W��Sa�z@��3���.�Y�����v3�GN��KSk{4�X�]m�܃��a�ze��*�pL�,gXsB�!<Äk{J�3]J�.���2L}]�� ������`&1����hCb��#0����$*
4c$E@"1��L�i�́���HDh�0Td3"���	3����(I"R2�b�b�&3!�&�aJ(���E�hH�iA"شNsWJ,�H�%�i4`!"b�"i��h��26"�b���QŠ�[�$���6(�	�b*��HLE���%Ʀd�J4�2$\��@F���I�� *K)$�$h2TD%$2�%�CbI1��$j4d�1�1��ɔR�F�1�R%!2(���8��B�@��Q@��)79�5IbA4FƄ,@Dh�i(�jSb���	,�i�lD�-��0����E1cE��IH}T(^���7Q��4(���ȗp��/���0��p�yi���N��fHop�ٸ�s�V=Xs[�(����-<]0s�Z][ճ3�U�����/�\�^���h/_~���]/�ޯܮ�͍���^�r�W7�~�ͽ*��]r��ny�~����/�ڷ��}���}_|Ǉ�}����?X��w����u�.F��t	����>�qo���n�^����k�6�9������n��]��w͸�����]
��߾�z�殹�_Λ�������t���+������[��\�kA�[��~{���Bysr�1c�ye�\��`���E���]��vۦޯ<��龶�\�,����6�\�����-�\\n�����-q�W������o��=�7M�6���M���CQ�w\����x�=r��(.Z���=�.�>�~{��:���� 8��|W���W�_�����z����~�����j�W�����-�]=6���m��5������zU���7޹��j��ow�:��ks�zm�v�n��h@">v&���٭rs�|�|c�q��|���Ϳ���������o��o9�m��Κ�}������_/߼��׶��Z=���{_�j��u�67���_|꽪����{��^���ۨ e��m}.BO"*�����ޅ^���+��^����_�s�c|m�_˒����ۋ�[��񷋡_�qo���o�z���-q�6���[x��-��w��sn;\[���Uث��t��bأ�gǮC���V'3��}�W�O/��_�^ץ�.��}�ջn.��+��/����Z��t���t�����k/��W��W���۝s|W��7�_����{����Qo���_z���>�>�7��)��<^�eld��wы������ή��n���׿�w��F��η��{W����}�v���W�˥�~W����_kA��|����+�z����x��O�{�| :�����oy�fA�K�{�f�����m�W��yz�ݽsW���}b�[����������ޕ}\���ε�ޛ�n5���[���ͽ7Cow�]-�t��s�=��Wm�o���\�o��h�[��˄X�,}�$}�,{�,�<�:so��_~s����Wk�}j��ln7ǝu�v�Ww���{�}�t����]zZ�nr��+�qi�����U�o͸���:��/��:o���{ꯋ�M����o�� p�fwEy���n:_dշ#K�i�WnS��b�K�{?d~��}	m�2�����3k:�쫅�N[����/_b���J6�gP�J�"����
�ó�>�O��/��T�N��t�kkf۸�&�t��������F�q�Hue��iU���B�ŧu�΢��$��k�����k�#�S���kG��/w�m�������ݵx��~?u]�9�_ۯ���^5��oK���εv�/�~_<��~^֊�o���B"G��i��#�(G������i��R�k���_���}b�H��p��W�s��W�w���o��]sW忟V��}��o���?w��W�{�֋��V���� �C�ECs}��Dh���#u�����xl�v�-?T}Q��=�����+���>��+���q�U�q�5�nu���n�~\]������t�]+����}����|m�^�?_�u��>#�|Gޅ�����D}5-�ev�[����m����@�����'�#���=~��{o��x}�{]��~]-���_W��띭?�����s��ޕqq^�\�7m��6鷽띥����+�>� �|"�g�=�ЗW���q՚�*�.�}� }c����.��ߝ7Ƽ��W�].?�}]|�]-�q�s�k���Z�vߪ��U��6���W�ܺn6�9���sQ���uц�E��1����1>��}b�����gzs�5�}���>�>��D��]Q�^֊����v����t�������ǋ�n�u�u/M�:����^6�����^��:ׯ|�ź^�r�vۧ_�k�_yzm��oϮ���6�ۃK��珞���y�8�e����Aj�z��X��#�;�K|_WJ��>s�9�����ҽn|�Z7�z������5�t���λ[긷���םU߾[�]?/���W�Ƹ�_��z_6�W��w���Kzv�����[>�3�0�ǖ�뾑�.��zW��o��{m�^�����[��n=\��.}����ۋ~o-���U�\��������zn�KG�����^/mt�.���έڢ+����]oKO|�� ױe�����tݙ���oH���J����u���z��5��]-꿮su��{WKO]������q����˵�o�����抿.>6���W��ހgw/�p�1�����O�z�R�g�a�]�קU�Rʼq>c�?n=��u�kF��=}�֟9^���z���|{n�mt�����Z7���|��o�����/���w�k�ܮ,x���]�����s�=��{mگˌ��?H����w�01uk��px,�"�v�MLƹ��;XF���U�جsmgr�;hG-S����w�5���h���p��YC����١�3SzMfq��z�K�]L0�����Ӭ%ۋ4'-��YW���҅\���-�z{q���ݻzW���#�-���ߝz�\�ˍ�n/�v���y�Z�oM�7��S�/Mv��_�u]����_Z�\�^�k�⾷K��_˵�~}�s|oM�_˦��st5������58.:�M9K�3^`���>�|�	����� @1�R_����U���;�+�p����ҽ+Ź�?���5�����[�����ݷ�_>���W:����]j�o�z�r0DV����ös�>R�𼉛������n���˦�=s��Mt�˥WCb+�߿;���i�6�}��{�}~[�\\�ﭼn���m���έ�zZ�{�~�^�r�+�O9s�/m���5�D`�#�H��r'|�,_�������򯋎��.Ƣ�[�|����Z��n�Ϳ>�����os����}}\Z
���]���+��9}�x��W�_[���[��ѿ����ok�!#���bgY�q��+������v���]7���|�,|^/]s]��q��\���J�.;^6�q������}��}�C�|Dp��͗^���z������.�����V�o�L���a��T�«�O�e��-�_�}��|W�����������ޚ��k���k���]Oܷ�u�]]������{�r�׏��k����\[��m��.��\W���o��ox}���_��S�l��ws��{i{;��6��o�������������z�x�>��־+��Z�~9�zq����������K��o�W\�h6"�\�������������J�m뾮�p���?}/ۊSVWO��Y�Ղ�#Dt��>��o^rߕ��?�u]󗍺��{�^�qq~m�������oJ�.>��=u_���[�y��v�۵��j�~�m���6���^��WM��9�7W�"ўN��'���e�y�=7�0`|������Z��7���KϿ?wo��hޗ����վ.�{�����[��}W_7���I ��# P~��� 	�c돝z@�~c�DC�1C�|h��"�W1"���c�^�R�"�!�#��
6̌|�;��q �����zE����.�]U��}NԾwjo5:nǂ��c�xė����Du��ia��;�딦a�Hd�T�5�x y�{��'|5⭠A�D���� �nvamj�Ȭ���et�K�����jSz_GVv��NP�قa��hrH�*f������:���g]���,�h�:�W�X}WD
�T��bbS�^(�ݽ�@��x�OI��*SM7�3ӧ�׾Gn��^�.S��=gI#�h (@��2��ĳ����/���XyM�q�5y��q^��*D�X�DX�t���?34�}�kU.׌ϙ�O�u�[ia��Z]�7Cތ3�=n���<�T7,-#�\x��0��a��[Y��V�**Ӽ��򥚭ox��VVdu�w��v�`y��� V{�	u��L�`џ�6Ό[lC��n#����[-`�����e��^b������1[�g��X�v4�\����Х�f7a9�C�~�.2�R������؋>�6ԓ����8��\wc�r���^��Ě�2px��+�C�WfYU�U
�<8��T�x�� ���A��o1�h��)�%;��v��=�{~�O����@s#>7lT#ך]S��~ S%��Ǫί_�i�F��]�Ѵ�DM��\9����!ÿ���w�Ƴ��:�q��{MA�w�)���P�W<�o^�Ef�>��1v-�khx�^�v
^�����Iu�N�bb�o���ڥ�� ��x������j�u�ʵ��u�cWs:�i�|:�{��ݭ�38�~�-�g��&�c1>��c��_D���7p�郸Y��<���#�lݣNU�A��ty7�(X�A�t^*�7�]Q��	�Pل���-vM���Hh$�|� ���� ��JYo���'+�[����о���F%��v���rx}���m\0��\xؔn&��;qe���~D)A�G��P똒cYϕ��h�X���KJ�q���eU��o�T�N�Gj.<65�}�@�2�@� ��S��9�C>���9��}�����/Z���R%�WMѦ~L�g!�T{����Wc�ܔ�Bi���*n�g��2G5~�o�)_�Z&�u�n�pȐ��i�$a��m�+NeJq�d�R��7[c.w~��5��iT9)��Z��"ыa;��sw�W���,��3�£3�m��z�T�J�8�l���_n�_R[R+�R�4m7@kb|���5Շ[1�>-zع��6���凅xX�,]g�K�v�f��:��U"+�~�(wO7��SM)�oUM����kT�xY���2<b�ć��\%������Z5���a�����_�5�6B����d���H�ݲ�E���*4hn3�C���{���ԠY�4l��o��E�np�a��T����p�83ʐ��ٵ��m�J�@�����8�����f�l�&!�2	a��9n�Ba<�Dꣲ���XՏ$��MU�n�҄�k9���?�W�}r� �63=�P�Ά�+ƿe׏��&�?c[#h)��pZkc�}WHlSoڐ�׃��yi�2#���<��t��e@�4Z�}�N�7�M�wmz�������7érokC����L��� �[���ڪ�cϛ���dW��V�������:�m�8f5���v���I�xf �y���1�9�o���2}�³'�ޕ���3�jZ:i�U�t��d����rj��&pe�T�ً�r�>�c|��:�eѴ岼��
����»�����wP���xyxuz�L��;D:+���B�:K^�M�f���m�OG��r�q�[����������N��ry����C��㤞e`
����U��KF��Ko�׃�p[i�m�3lf�o�*�csH�܄p!�����?@�T�j�1�R�r���g�
�g��%�l��R���vmE9�pŕt��7Df����BSIyp ����:�ԗu����Z�;뇻R��Va�A�E����')�|!�g�8;܌<�@:A'a�Rw'q`mO�sُ}Vy�o�P�}>y!>��G��ξ&u�3����Ωʽ�R r7�z���|��莴^�˕"$�X̡�"�u��zwX�Q^ϕ�:q�F�e��lb�{ݛZ�=Ԑ]�H���Y����ñ,��g�ǝ|Zj��j��_[�tX���I,��;���K6ͬ�<eLG�K��'t�7����*�V�G��hb˛D�|�x
N�ŃӺPZ��ُ���eez�#�A�E߆8-U�8m�v{��k#�-�����L�̋k�79ӓ`�hoD���[�j46g�B�
v�bU.^���s���m�<d����m�ծ������;�g�
�4!g:8!��҃#�Y�H�u�^����콽�i�w��n�K����j�_(�Уf�����@_L�*;��6�k��դTv	f�G)۷[�/�N*aU����s'�$z���������p��hL:�9DB'����.vWlqܺ9�+"�+J�|�i6n +��Z{��/��%��_;�	f�QP���=�8�9��n�����!�S�<�ǣ��|h]s���j
�T�cy��bk|]wG�AJy��]���8
��?&)�C��i�m��� ���W-f/+�¶.��yb���mj���H^��u��a�5Q��������O����ô�J^�a��9�C���{��.�������Ie��7�GW	7���9��坱�x%F�o���S!Z��2�Oi��I�۷G2�8y�7��.�[G-e�Hv�uҏ,E��:�b�%)'m�}zf� 9�c��j!�f�1,�Uhhz3M�cm;>���nn�mF[��)���������i��
��~�F��N��PzaH)�дs�3_���_v��=g�_��}�3~t�<�C\��z2nJ� ���FHQ���עd��������(�|���&P�FX^#�ۄ\���=+|�#��k�g\��@�V	�$T;]To]�6��9���!�.笽�
��.�s3�~����p�+�zP���[D
�@��5dДa��Pڍ�-N�AAmYd��g��'c���^�u�}��k���W��H��Tt��-��I���[�d m���3����ݕ�G���3ʙ.`y�@/��>�St�ޙ%�;uN�i��f�>���L��V-��F��+�%WFǑ`�nX_���\x��uJ�~zF4�zd���wni/A;�і��=��*3��'�at����VxX�����1�H| ��^���qId\�	O2��GM��~��ï�s�T����?s+�Q�~���M�Z��&	 ���"�����iނ;b� +]�Xʣ�9������㚙פ.�\��R�3���)�S�Үpy��;OL�o�1І�:3��]3n�w9��l�WYs��Ί�uc���`�o_r�R2ԽY��#���Πĉ��)F�:׵������.'f�ݓ�܉���قC����r㤾?X��t�b%>�6��}Y�����_|��~�ez�jt���{��Q�
���v���{O�ve>^:��M砏IΆX]=��v�)��.m)�k2�����Y�dP۔���u��E�r1�:j)Hi[�Z��F�v�P[��o�� N�nk>~�#n]h���5��^�#�� �_pC&�Vq��� ���s~�z�b��
f�*�^�.���N��l�jX�^�媶�\Q�I�6�����ghfgi�,��LuҚCW�P�n�F|�?d2�^��m\1cf_ۘ�2!u�������.�D���H"I�&�JbI�e+U�7�� �Oe�#=b��7��%pe�^��eԣj�΁ a׳P��^�{g;��	�:z��;�N�w��H��l���t��'ptȔ~�'0Y@@�Q�Q�`V=�vy�,��
o��ӜRr`
=���u�A�P۬����Az4�M|H�����.��xM6@�3���
� 8��lnp�Y�g�ð�\t�(�ݫB�:���6� �;���*a��ک�;f���8�B	����n�[MU����i(�C\�R��o9Mr��C����]���\��°��c'B1��x��'/y����ؘ����ļˈ�|>����:;���o�D����GX�C���� �Lx8��߁����5��r�\�=��!�-<R����p�M�j�YC���%�#QL�;�n��������2��ޙyי����8��gEx`�.[g��5
��yN����H��~�(wO6�S���\���9ksjf��.�Qf!a�T-W�V9�k�l?�+�&|m�:��o��¡�Pb�,�j��XWL�͈���GA����g;��Θ&�9�6Fڑ�WѰ���Gk��"m�s�vi����3<\����3Y�Z�y�Ŀ�a9�⫬��?�V,\ǘ��ݯ�i�z��mf�=Y]wc���}ۨtE��{��u��C:�E�Z#b�� q5���W�>7O�k�`֊�����@ڈ%&3]k#�*����K��B���QН[ҢJ�������&:#	X�M/j����TmW�ʳ΃��%�FӖ��;W�aB��K�
�?0�����G�LX)q�=Dep�W	Ik�UK�4��[��]1�ǜ:C�#��:�m)x�:K�=��A��^[������zn�txշSIW�,�!��]E5N��}�4	L��&����d!gnK�b祚�b�����V�5��i1ʔ��Z&�I7:nڋ�h5��q�;��J��5A,��-�mF2)Gxd�]p�cn��!v13�2+�t�[���#��1"q]]�yj��-�c9F�Rt+4k"L��ʈ/�:�>��7]�|g;���w���+�@ї��W�J�2�%�9�V�I�u���;��R�Qj,��T�0�SN�E�r�]{t�5R��*3Uػ�
X�yUc"�Uúڂ�+Fp9�GFވ$�k 5F��c]�ɶ��8WS�*u0;HX�ӊ�m��X�V��G�ّqO��2��-��6�;���ˊ�KY@�'����t@�3%'���&k���8s�ۅV���b����s�E��4�l"�i��mu�BQ�-�F�s�_;��S�p��v�EnN�p�4��!s�o] X�)X�ջ�f�沅$����Ψ��dbz�ט��a��� %( 9���|r�RtiA��woZ5v�t%|�aVn�{n�LЀ9�$k3����&~F*̊Y�PCy�-Od�bɵ�}��F��a˭ₕ��(���755�*}���i���ӫ��ZW[�P�����]��}���S��f�$�ۖӾ���p�I�5gh)%���l҉#7M��ШT�7�e.jW�ws�Q�Z��H2�v��%����)]��P$�U��	��c���1D��k�c3
]4)�k�΢��8�ۋ����}$v�2��qn�Y�.Q�<`՚���yZo 괝:ڔr��0w�d�򓙐����s�)Krta�D�kf�N�Fw�r�A"�p7�^�"��u�X�M�h=���w�{���<e�f��Z��n����_A�����ux�mu
]v,��Z"�I������؈���������-��[	H�K���Z"˴��v;��+���E[�֦V�l�qͫ%R��c�;q����L:;��m��,.)YwK'|��U{����moa�\�[�l4f.SmΎ���ǔQ,�#E�wH���`J����p�\0���|�=���qZUr�e��s]F}�L�wc&_!z~[z�<�'7|����7H-�fκȰ��v�ቨv�
?�\3m�~@ݢh^#*m���o��3��Z6��
5j�;����&��Gf��eվC���DF�c��V�Ʉ���z',�u5�N�}�f�Ĺ]tɻ�G1�U��e��N̾s3��}�{��BC˫�#՝ft5e���rGv�j����-��7c�I��� Z�ҡe^��L:�vا�vUi���Ě��6�̼�tPe�I?��"��-s�fvMV�6���}$QRK�%e��h	�}�;;���)�Vi�V.��]r��Ct��*L,M�L.�N +v�r�-����@}@}@
@}@V�n���P�6#A�Di"�
LbKh�c&N9��-�F�DV��R1���b̌i��� $QEb��%JF
4��$���L"2�\+�#���܆��EDDRDqn0�AI��F�ň��QTF"�RQ���e�0E�E�&�,2�n0Lƌb,QI��	H3LDEA�Q����$�12H�d�#ZJJ,b6(�cQ�9�b),H�QEF&IB&���c�M�FF�l�s�qA�d�� �> ��@G�i�Ā�M8vj�򚏵�;*8�]Z���(��tL.�/zhTj�c�Hδ!�� d;��z��7�Q#j����[v��q�������5"��|>6Ȯ���Fp	�^�.�aN�j��P�Ѳ�Q��B�\�<o������O�8��������0#�#��2,D���#��6��r���r�k������CZrxԲU�Ә��o�9�=E�Bi:�r�  ��f{>�ၽ��I��ٕ~��j����f��q:H���CD?M��&쌺~pQr�O�w������@�2j���Jr^=�zc�,�V�G�1��%k5�/lϚR��㽑Z� '3-j�$i$-�M�1!1���(e�1�������G��Y:��ڌ��S�_>.�[�%p҅7T3�Z�t����Ӷ��vy�@��#/����XM�y%�{s���21�>�>��ҫ����=V�=��Wl	���D-u�*Q�2s��'s3ީ%	m\��V!c��$l�_���p��B�`�BGa�v�ֻ�x�d�-�Y���u#�":��(N������:(>K�m�{�w���D~�$�<:�0���S+֨��c��ɗ)f�B�]��y@�m*��p�ck����k�{$�)��ݝ�eZ��r�[k	�z1Zu�m�8)�3��ؓ4bۮ�I��F%��tusl�6�⶝�uj�ݝ�I����^I�M����v3m��L���UU}UU�{W�\���~�,W1f0�N��X|�ܓ7�#DO�3��>:��j���"�VC�L�Ȭ`��5�k2Z�r�J3b>CڧՇ�]�G��^{�B��w�aŽ-%�d狳L����o��/���(T���(<-�1MrvLz&8��O����^Pz�S,��m.C۔���h{��1I���B �,;V���1���4����^a�g+��Ӆ�Yާ��#a��������֦�5��:v0��~�v��
�lfE�k�]��+�&h�L��}��{���c��e����C}󬿜a�+!Hy]�r��pGs�)s���w�L�=�6>��hL�e3\U̡�7�a���7Jx�G}��?�k�c���E�G�#/�$C��d��@�Έ��`~t���Bs#4�=&��V5�����*��YUfb�$��ـ@Ɉ^M	F�f����Q��Wt���)ξx�ým��g�"��[ޟW��sO�ϵ";�8<���<<����I�՛�^x�8�]��3������r̷2gڠ�ˋބ,���[����YQc̅Ӡ��u���;`V ]2��dΨ�D+�҅p�;1j����f��3�Wl�9�CX�-e�^<�����S��y#C�&f�ef����|�������N�$d�?@�s�6�Ip��S"�
�����?3*��}�U��.֯*s��`�>X�>�I8�J�z�Ը��^�=	*�6<�Sr����������C��A�����5��)�2�8ț�mE�{�ٕL֓��!�
ٙ�	��09���Z��þB�YD��pź�_��[��!���k�t��Gs��h��Ɯ��y��x/��w���!��mwxE�\=���Vr��0����K��K��b%>�6�q�g:;u���ç������V����<�^�2͉�G�U�P�i�����|�ug�z�ukQJ�߸p?eet�̸��sI����1�H^�cy} 5<�Y~�w���ύݻ�~�-�w�lZ�{
꽌�	��ѫb &XsUksN����������۝$騉).���Ae_��ͩN7�u��Lc5��Y��U0���@Tx��v��b�g�}mUg3/�,�B�{��y�rR��aN�I�$k�rH��,j7��(=��,gLqq_3�CCw(lF�K.v.3;w1�/+`��n����r�9p�mZ��cP�ϲ'��W��yGtm���v�U��>�3���@�G�Н@��*NͻM�ڿ&R�?��k=Ǉk�AC�.Wu:TQ���ս:�����d�� ��9���Ӄ��X��=��I}�y:T�(����������gI���V�~���Y�jH �΃PJb�cY�j����c��׎�-�4�.��.���$�o5׃���|Y����`eԲ��~~9:�j��u����8�Wb�i@��.�����c<�n������,�"T$,�4+�(m�g^�4t/z�����ˀI�@;�F<<M|۬���&�Ȑ��i�F �[2R�MU�.��v[�"~�1�!�j%or�<��N:V�Q��WA�5'�F�/\��KR:8p}��'���K�Ф�����b~P��H��)�F�7@k�5�E���������Zc^/U�S��K�l�)w��-v�.W]wzFi��II/�4hO(��{{垫�P?�m���y� :�����U�f�fç��(�ֶ��o��~&���N��E3"��3�D�q�!,�SJ��0M�}���5Ѫ��8X6�~y�ܡ�H�?z%y ��!管��#U=rё�/=�k�Q�J�c��_�}|�%��p�QZQخ���pڽ�K)�2���֏�����DZB+<�����yh����Rc>;���Q�-N+$s슯9Z��:l�K�ru�yrs��V�i^�7��]v�ս��m�g�K]�Yi)ب�OoD���}��>�W�g��ct�G�Il���`״�*HtEl��ܗ�u��_gZȧ�Z"��\]��>�7c�#�G�<x�(�ʷϒ�H��W���_�"E�,�R�b�l���!����ˠͫ���Tief�Qy9�����N��N[KڪS��G�m��D���r�T�-�>Bߧs��{�n���UO�o.�c�A�Exk�+�K^�M�o+�������⩃��^�����#ipP�|ڸ{�R�����$�8�i���I-�������e��:�VNؠ�������>��t��,����s�N�>��Pt{�L�<�ouzw��ŎO�-f�~��+D��~ә�23L�*Ǒ௼��@�O:�	->/Ot�m�r�_(�i!�ɼ:��6�+���RE�b!�l�n�˧V ��y��a�� �(��Nd� ARV=�^���aTj�h����f�+v����ԹZ������žZ����xX��I���E�;#�aF�2gx������4k��zu�X�@���^{0+�X���x�SoJ �Z�/j�<�Wme�h�*th��1Q��ɫ�{-7�}[*Dp
T�e��v�y�Kx6xWL�C/����{ٷ�C^d��uj�������ܭg�:������sv��a7����/0�\i�X���U��'Y��O���G���A|7���/3�r_k����ub.^��p���rdߚT/ц~A�%wB�e��?yx������to�vP��h�?,�$�N�ZpҶ*x����Iǵ�k�c�a��ћɊ߻<ǋ�9b����L/�	��a��|��8��u�o����m������:��AƵ:�b}��}����$zǎם��o"){x&�l&�
""��ˎ�ҳH�f��f��k�f��"x�韜�j��s���޺��<�Ҝ>�L�E�l�<%x���Q��!�X8�z>u��y���e/U�y4c�h{��QN���+ޙ��y`Zg ��W	@��uNhEJ��ǌ�� gR�۸7����c�Ih�X^��ê{�?�,���<!w�#��[��Ҫ���SK�t�^�3�de9+�y�Zj|S��A��X�-ǝ0�]|�uW�B�6
4��t���#s!�,ՄO)�����x+=�N�g`\��v[>d3� o��m!�o'ެ-"N8}�]u\��󄠻l9wDք�r�3�#�d�y��'��d]�V�m%�2)��j�T�i���0]:����kv�p���g�������U���������Z/gA��<5!0e�=���P����\Њ�Ws]�����G0G1�כֵ�������d{�$���`�`�X�`h�j(Δϗ�\U�2���j�ai���+����0�X�����V���a��!O�4��/�s�B��EeP�� c�q�r��!����B%D��>�sݝ8���8^���j��V��M��Z���1)��Ӄ�G�;|dY����.��΃-]��8]��=���f�E)2��ѳ$%�Ӂɯ��14��'��~��!^&�U�֊{��b�\�P��%�,5DX	�z�:7�Izo�Q���ڂ���':ְ��Q�N��<Phl	��]t07uR5�yl�<ZG�05�9)�SǳT2��eѻY2T(s�),�l+�Y��>fa�
�A]7}&����3>��
�^�b��Jؑz�}a����;�]�
���j�}��j���:bxie��^b�?V�	�6���h�-�=:�M����BbFt���__L#�$r�h)|~k��r�p
��n�mq�ү^s�I�ݛ�&���kf��o�8/L����Q�e�fW��{O
�>^V��P��Ƕߓ�Z�: u꡴]�xM.p]����LK�����8����H��CR`�L���W�P�ޞUW��ɪ��~�2��x2�#�x�}y�azv7E�S�+�
�I��wW^\�.�J1�Wr�-^�}�vm�{�W߾���菵-jї����x�i���/���H��f��ઈ@s#>7��7uKBE�#-{*��of]x���H�) #� =��[�ȇ�b4��৞�}�Q� �)��q�8X�h�G�	��U�/�3��I����j4����.���~A;N���Lg�V^���/��4��$G|��O/�n"cq��dh��,j6�J3Q����k������
��A�[v���Q���ݕPq3xb����D��ՠ�}ܪ4�|g�Ƿ�߇p��cp����L%"��rr~���둇l�Oަ��c.��P@�PV��� /���jv
��uc/-T�s�T� �������+s�=��7����ބ�5���	��Kՙ%���N=���o�®f�ˀ�� �/լǠ1��ju�n�s�"B ��ۻU)�ku��f�����J��l�xO�N�B��UJnt�:�`��F,	N��L�V��iJ���ݚ�*�+0���Gq�r���fa�/w���ډ�d�ߓt��.����*���/ҝ#깗���fqĥaԇ��f謋��D����9�jm�%�v�Ժ�u��u:܄��_)�j�҆.�� ���VR������t�O�B��]��B{똩�ʐ���Ye�s�� $��#e5��:
k��bܮ��TV��~��>�����ΑQ�L�� ~���U��ת����%.[g��P<�]�5�6��U".~�;6���Ǡ��w���Y��q�f{m��]�V��Х|�y{��k�9V�%<�\s�ؔa/(��#��V\8z�	� }�7qXo_��9�	x!�ؠ�F��H�6rݖ}ʥ�P�Z�|9���(3����*��s��~������6�+�~��Gm*��l��C7�����s���{'^�����+Ua�>�vR� ���uͺ��U�{��u��@gZ�}R��	�#\5j�z�ގ<Z$�_L�(͡��+3 v
 ��8�p��C.!K�=1[ymF�^3#�W�<�����X ������旵T��C�j�6U�tQ�'�"�5�e^;누�2�u�N�ޗ�Fۿ���9�r�K3����6�;;��l�+e@؎ƢێAu]���{q�u8�א�pX�j��3�1���.��ޜ��ܲ�<�-[����<��s�-���eǜ<�����w,�_j�����:��,�XP����G�1��[�I��m��ew"�V��]���	�N�,�9Ll�7� �Z]ю�7NL�Y�T�m��[�4N������x{��[�9�O	ܔ'5\ե�a�t�v.��y�ō�0���)�����E������泻��;�I^���sPRݰ��6/���K�i9.їN=x�)�X�adHM�����1YM+f��	�s���bp��� �5���)� �˓j鋝3k9�{1���V��8�
�3/D�I{��Ey^��=�]ϕ�\���#���-]���eG/��҂��Dz�o�����(�^ba�n<��N.']��/j\��G;�|y�hn������o����~P��|:{�=��B�1#:�����Ҫ+CL�]�o��u����M�]^9�u�M���ҫ����6��)}|#>N2o�뽈f�*�Ck��rc,s��]LN�h<�	��y����x�~z�w�\���Ձk�unL�J'<fu�(��7�jZ��i�3]{C&sEl��7�E���r�>�|]�M�o�/j�X�+Khq���B^g�\v*��+Ns�k�{n�/-U�&a��سKƋ���M+�9��qeɇIW[o���c�^:����qC(c�L�3zM/�ǘ�ϔ|��F׷�Bn��b��x�t��dc�l剘3/"C��8�ܦL��f��J���Bjnp�m�z [�� {h��gu�Avh^M<R+��7(��Yr�.;��Zl�n��}�u\�ftM���[��;��e�1T�x���9��ڄ[�0��s�.�H!(� ym���V�%&�ݮ���|�Ko�e�Xw��IB����.T�j,|֞հ���l��u;��-�d_N��-uU��&.��\]�*#7�J��2�7�4�>���]sj`���g)�jv���A�%#�r`���#�@N&�_p��R�c�ιs$�0~���vP#L؊u\�-J�^gFr�Q���!�0�Wbn@�w烋j�A7��L TX�7�b�ֳy`��u�ֱ��0���C}{�S�R�ql�2�4�������������F\��ܰӬP�Qǂ'����o-�L	��Ŋ��]����dw����k�&at�X<X�a�f�.摲�!���.���
v��|p3�|b��X��P���b�Z�8�t��Z[7n��3HѪ��r\�(]wt��*#�@��WR������ú̠w*�kDi�x�ys�$N�3,��V$�l��[Z�3ܤ�,�9�V�����6�{�m�{$6EO&������k��eg7�u��8�EȮ���7��%`ӛz�}חJ�Ff����˺p�j��	��2��R]�&�f�>꿊Ը�CrXV��X�ɽ6�CC�X�fi�U���tyԯ(� �)��u�n�uԬ[�n�˼[�S�]�,$am]L�(�=]I_Y��x����r��H�g'�xve�[��#��1����[����`!�|Ca�4Z�2��LU��)c�̼��±+bܓ���g4�����:}N���K�xa;f�'Hq�s
#�O+c��T�fwMc�0@(�I��e/���0��\ƅuf���gd��f�T���]f_s���W�H�G�t���}�<�PIŜ�ٝ-(Ɇb����p���e�ƨӏ�L�:��^����C��<�r/+;�I�F��ju�?)(�'�w��� >�Pd�bZ}�6�J޵ԕB<;�ʝ-�ݬ�ls��/3og`�9q�']w;��h;��������Br�VZ��n�6�<�d�V�X2��|O!+e�;�m6r��k��1jW��FHL��&N��|[O��Ęa�9��	1�(�X�!)q2�����R ��V��c�I�c�W����V���m*,lLQ�)�78�M��ܩMf�=� �*Y�����f�L��w�*�&��r҄��O�<Ǯ�h�Hv[�&ʻQ����ƴ��Dc��Ӯ��]�qȗd��P����1d�A!AȢL�,�ԤV*}���ƒL@�0XK%&)1�ES,F�h�,\r�!�-��!�5���1��b�b�Jh�Mh,S-,Qb�&��(�WƤ�9���Ѣ+E�F�D&RH#��6,�Z-@�`��+6-g9��i5Xf���ƫ��ʊ�(���QBQ���h��sP�QTm���Pd�"-Z��8�r���8��:�O'C	��c]1��=��L|�,>,�O2T��.m@�pY,�R�w<l_2�n"�(��C���\.�g>��������|}����R����צd���]_��7p�@�:^Z�]]�)nj���̭Wˍ��yS}�<$VvwO��{r��7��kӷZ��5K�ᠠVR=^y��f�z���k�uW��0���Z�6����_�}��YU@׃eЩ�����7�xM���$�!'��[����Y~p���c6ܚǮ�n	�����Ǉk��f#=_*9Dv�C����Z��K}��ǂ��&c�3���k~H�������d?\#����
c�s�_<��Ƈ�݊���;�ܓަ�-�s��v{�]g�À�}�.���y����U�[oO�x;)�s=���c��W��%�0�
�ߢ�sniL������o��
�
������=I�Tr�}	k�M�w�n<���NبSnj4��&ڧKs/�n{xԤ{�]\��r�z����C^�J�/�i����2㥇r�����+�\��V�ocV�'2�ţB�R<+.�u)YB�8�G�lPy�v�4r�B-���)��*��am��u����C�@hGS_kʶ��
��=��qt���kM��V�O�{34Y� O+��}��*�ov�A�`��fE�kG����B��ɉ�Õ'+к�u�q�<�W�\����9fۇ*ځ��ՉBl/2��4U9�ݗ��.�z�2�De�ؾ��<ڝp�tԮ�g�{ι�κr�-�Θ���zy�G{���tL�*����� Cz���S�z#���T��w�i���ڎ��C�{1�[O�˯��h��bj[���M[����pᑯ��/��z��y�U�R��5{�C���|9uzn��>��m��}.x��|1|Ή��s�|�����y�N���(S��z�ed��V�� 1���R^�J�U�Z�.-BO~M���Zx�����5���c�C����?l��
����	6�=:�ʚ�o��8k�J���Q�M���
�=�幸�����@S>��ȓ��q��;�-j��o��eK�3�G�����_?i�D7M�Qk�H�	D�׳*��f���&��,����l�͞��dn�\���*�˹%u��?���K��k��߄�q�J��-��Y���#%�efu�)�[⦾l��r�ɕ���a3�֩�{��G3�٦���oabN�d��\w��˩��w�]�D}�}�Z�am���]��l�׻a[��y����.������`����j��S���<j�����^���^n'};���x߾�����S%:}�fRL�{��@*"���ٲ^]�y~	F�r��dp������4P��<N�ʙX���z���H�R������wֳ<9�kO���^�Cx�L�m�[������'6�r�v!Rw�;�S�!�<}<ͻ�ܴ��c�7���}�`3��{�ZΗ|(1|#$C�B�'�:����`��c}y�k��7�V��o�J�Zn���Χ5|"�+��\��N`��f�Eμaj�U��lz��ק��(���=�9~y�N�>�������*�J�wl�ƪBO�Դ&�1 �Vv�N8J^-n�1�&)�M^7;�o$Zә=�xe���ƪ�x���tvXFO�ug�zz�gsuW,o�L��O�i�9\}�h<m��1u����xc�[m���F9�Bˈ�7v�e]u��6L�#���T۳�r�33�۸`��@�ܦw��]�����] ��q��x��mp���ѷO���V7���4��h��J�����#���X��}_� �et���J���Sݹ�U���9��t��]^�������Q�{�1_��b������Ğۭye^�k%�h?������Q��F&��C�G�\�)��C^���eCi���e-d���̟BOә��NA���J��3����ϩeV���m����b�i^B�����a�^������u���AKv·����-�����*-�d�Z璖u�[e�tK���X�E��y�ސ�/�U��xDeP^B[J���Ehs���?��O0{je��t�=����{;�
�V����V��a�ݯ%�qx��$-�����'nk�S.j4��1H;}*w����Kn7�v5���܌���2�ð�y�B7�\Lk�:�g(sK�iu�O_M.v3mL�ϲ9ն���7z����k�����i�|(<�iv���������(eAթ�f䌳"�浧Z�"v�1�ew]j.�hκ�v�(!]�V�K��Gm�a��op��Uy]ǯ�9ݹ�[��d�%c���� t�{O���tkO���+�Q� �ʇU�*�\eżCBy`�'|���_�M���0p?�b߱��Z��=��?W�O��>�=��P�7D9ɽ�rz�X�ШD������O8h�)��ɞu��:���l3�M��S�8+��'��z*1o�>>�g�ҿJ'�aŵ���]@��:��KX��[�����P���+��}Nn��m|v�;5MKS��=)�Բݍ��<���L����kJ㾩��_-����2�ͯ��N��cv���"\����\t׺�6fv�R���1X��H���Z���{r��mBkӷ�h%o�Θ {��N�m�g�rqԨ��R����y�^�6��Zyj}�2�u�&}�}���꽢�2�<�A�y��N��/wQ,Vgu��t�m��6��Z��©W�p��)��忆�U/���#tHiV	�<ye�B�r�N�7�!�R�~Q�;ąm�+x��R�e��T�������L?_8��Ƽ�*���"Il&c�$�<��AA�%�u�s=�>s
,���ъ��K(��W{�[������ȵ��)1.��7���iq>�C4���;�*DÕ�˙E�gD����T�.)�G�k-m�n�Q��v��G�=Δ�!���sl�:�$oﾈ��x��'�eW}6�'��ʗL��d��~[?�5��ұ���~*���CI��9S~CZM+�w���S�sJe�ik��6�b�I�ǵU�5.>�o���w4*���|���7v�ħl#NP
��2�3����
X���,N����|����:��pwp��2�ZHځ�B\^P;=��9�P���,V�u�q���޷��3��m��%C1G*w�_d����}W����U�U���ͩ�<�MV�E�;�Rf�#�9�w�L��S����g��ϻ�s��ZH�L7�鮴��O~+���P��k��Z��.ߝ�̿O���}�����]}�GjDvl
������=�zyi�塕��h����.�[���z�|קv�o�=Z��RJ'�4�@�qT��D�[C�7�G��Z���{q/s/�x�l���-zءg����x���X�q��q����%�DD�mSah���	��!1l}OP_u��Ĝ�_���Z<,o{�4.������Ƙ���7�!�ιv������q���'i�B�z]�Fm�8Hw5�${7� N\hom�>w�˯�_W�-�{�yU�KT��1�D��F���F�'i���I�TiSi�g3����
Gm��q˸�fAQ��J!\��&���>۞SWo+����;)n���k��뭟7q,��Z��}�*J��z��PPZ�&O8u��=A���/t~��Y��q�Z��۱gқ�Ef��C~�w93W. j��ɢ���V�=�y����TK�j����T�7#+�n.��^)��te��0c�w�on���}����ws�x��n̺"�^E�����}̡B[5+=뀜�*�Z�z�vǺȄ�,V��8�C��vi�Պj���(,s藾���ٌ$�d3�J���X]��k^f9�)�{�;Z�X�|(Hή��E�n:bw���z2duQ]_1i�O0���A���T�᳃��ZΖ��bo�`{b�o���jv��i�;�k�H��Y��V��������b��\+7I}'b�^T�+U&�u�ز�5�z*a�������u�/�Wu�h�;��k�SZ��.kWc��g�'�گ��ؠ���o;�gw$�'�#�,eV��ٴ7d��G�Ԟާou����>է�9�����}��{��U{@�����1�D}��`�չ�g_/-	�>�	��ɝqC7���zm�]�t�W��=<���T���W�����s����z��)�q)x��ړ[w���|�G�C�W�kÖ"'�{Nz���z�A�S�Н�=�E^vpx�5:�b!�<Z���˩�۽|&��U�]���7&�8�ۃ�~ή���g�' ��Z=��ʪaְ��m��3{���.��X���M+tӳ�"e=���/֩_E)j��]��^�8YM��ޭ�e�P�0r2�&��l{[��߱�D˓�;�R�E;k����TE�����e�·츘�>��W�����dL�_I^���%��@V�=�b���X����"���z7f.��$���>1�%���afF�1\Ҹf�N��r��n*�3N�7�M��S��)\Ln��>P��_�R ԒgQd�N�M���hA��+T�މ�R�0�u$���+�r�W��o;BiPP֓���
�l�y���:W&�&M6E8����͘]�y�h�B����R5�>��n���S���ҩ�2y֡��V���vz�����u�Q
;��y���׷'n/PN����t��t���Əg�]���>���KR��`�k�����ci-���&���
��uۗ���K�/|��ظ>��=���+�ߖk��z��}_n�|:pwp���]�獉~S��C�Kl8�vWWc����"����啫Os����^�������~��3ׅn�K�kU�'V�g�%��-�V��կ�.w�{���&�y�Y�2۽�|?:�ίK���Ck��뚖�Ӟ���)u��YAli������^m�L�S�>5�cer���o���C�_�maŵ�^�З���U����d����s��wc�z���`��(*��z s��N'�z�w��2�_w���NxN����tMf�t����믶^!��v�ԗ��V�e���y��0��X2���
��o��BC_\]V��(�,f7�Z��M�ռ���6kܡ��s}�K�<,O��Zr�陇�L�q�5�]��T/�"�a޶w�ͽ�f��"��z9Z��|���|Ytk{H�Q�>�6/+Es�����6����sK�A8�3��^W��U}�)_�{��|;]>���{z����k)snpHUk�2߃�q�M�x3�$�R^���'we���\J�s�����E���}~5O�>ݱ�]|��' ��U'S�yf��2�gM���}ݫ_�&s�{�4+z�O-�����6H����ɨ�K+�n���[5�Z�(��8f��y�]��yq[2u�r~�c:�ma�E[��{.�V�t���c}�֦���;�m�c�sJe�in3}g͚��M�"�T:�)��W���-�r�M�v�;M	ޮ��1Gt8�ꎬ��`ѵI�Q��"��vܠ'��z������(kމ�z���\U^��[{��w��(ԛ2{�����ju���~x�h}��:o'0��W���ǃg����5|(�_�[�Cz��Bu�A�p��[��)M���^�Ǜ����Y��B�dKc��5	DO������+�a�v���`2�F��˕�n��hK����Lj�_R/Jx�f�R�i�I>�D+��J���5kN�H�M='KwbrnD�����jl�r�]�J�|uZ��,[;���;�u����+v�r!�ګ�����u��S��1��V��k�nDv�V�+�ű<�2w�jn#�oe�G����]8�%v�T��^��T��t;�]��\���q��\
U�!v�JJD3���{F�+�;[{ˮ\��C���9T�R�����N�f��2т�)�B��
�J�I�F�ơɇ����w��+��/.�WT7��kTk��a�OR�I���:۰4��s.��E ��{x�ݔD�+��^� � ������Һ�7%���$[����yԱ/��vdZ��J� e�XJ�C ���֍�Kl7���� ��FV��0����������Dhq��r�(�4�z0oF��T��˭<��1uMߡ���T1�V�D>�ގ�:�c��r�-�@QG��u��ӶKsY��b��`�dU������u�T�5ϣ�q�fޙ����.�LZ㾣Y2��Ce�^蔢W�l�ν�5��EKr�y�N�ː&�$fd`��Ϩ;��܎V�%(��M�:r�iu�����U��:��N�*IZv�U�7;er�������������4U����*�3*��L+J�卽]�P�U��$��C.�;}��QnG��{C���*u�يkh����jwup�VR��Y��?fa��[��	(�ZfNݧV1qo���/v��\ck�����p9@��j�q&[���'���V���m�.�b�v�ݮ���d͜�k"/��W���Q��5d"PҺ�r�Z9WB_��^�4{��#{�"�溙{J�i��Tc��Ԙ���
�R�]��2&�R��-X�Rh�o.����X+�.���^�~Xͩ�ѝ%\��{�"l�T%1�-/8R�c�&���˴,Lwq������Y;{���Z����a��SJxn+���pь�:�ӣ��x�؁.>j�޶�j
̨hZ�呥��K7xb�V��U�e��{8��ף��Ye,�Ό�LW�&6^0&�P��J7B�֧;.��:���@G/��J�Fr� ���0;OU��x�s�8������ư�d�M�W��WS�G�<�x�v�(�r���fp�P�\��V�֦���֠�:�-^�&��]\���,Nu�������A�{w�Q����f٩JY8������"��Y��v�`duh*�u��Z(
Җ	G���dX󲤧�貉�)In�+GƲ�v�/G-CI�v��&<Œ�Ժ�Y�XV4/�IIK(Ƨj��vt�2�^:��ೋt7OUٖ���9p����9*�mp�$�ьNi�Υ�fb�s]�WE�J��TR�V�]�7:�삫�T�1�b*4BVM�QE��Q���QjKDZ)��h-Ib,F�$k��Ʊ���h��HF5F�*1F�F�mM��65I�m��$b#AX�٘�$�HA�m
5%&ƌ����X�iDDV�+�*�X��lju��ޟ�{����o8��h��e֚e�C� �s#�i�W%^G�-㕄-�i���;�`�������Zm"u��f����C)�[/�<��|3�������U;B�Ch�?Cz��噛�g�{���Co<�
�ό��f�zx�g�O�j�X�+KGx{/�^9�N��/%�.�Ft����?vy�^��9���v!r8�ym��:cY�|r�Azt��tv(|1Ɔ/7;��u��{.뭰�5������ζ��T̵��T{P9Ωk�Q��d�x\M�I��.S�iP��f��]\�O��$��9NqgM�s*��ӍI�%�ȈW*k�����ݽ��k���{a�\y�������>n�YK@L:\��~�o N�s܉�zu�~��+�YS��sή�߯���]˺�]C~��������Bg�d���zӞ����>�@��]����]�hO-;���م�Cr���&�F���clLsޯ���`U��x�;���Fm#4L�j��������qW��N�)��`�N�Z��(����j��Э	��L����]��vX>��h�~���k��+�z���[�to3�m�jQM@�VJ��oMR�)��Wr���ȋ���B�g<'8>�p�F-p�j�4��$���`�=��rcv'3;�KɃ��i���zd�������=�����vh"�~�Sͻ�'��g,�Z'����t��O'_i�c_�'K�i�Z�����l�雓	�~�n<J!/��c���N8��Nw>��\�[�_ҹ�uj�Ϻq	�-��)�q{=Z��fr���+��Z���bo�d�{j�w<�ӊ..&�����چ`S��,�Zx�O]�*�i��_gS��;"b�C���Z�ud��Z瀆�	��:ᯞ���dθ����;'��>�N&x������N-u9�Ţq���n�U�	�u:�ה^�y
g\\B��@a{���X�gZL��G˴�u\�+�?Xssط:�5uL������΅�P�`S}ͥ+��s?v�����{�I���G��k��B�G��d��R��h��^W9caް��&��ε�U���wZ�������V����0��\9�Z���͐�XG��;0i����o�e��i�t��%��в�VMJ�XH��%
�@�z��kg�
�jtN���r����LT^�]�^���y�3Μ�"M�����g+���m�f�Bʬ�|�����a�f�H7XF���̋� ��Z��wY5}3��V�X��8k��)���O�X�*����*V��U���4�Ĵ8Bx������յ�W�;γ�m��!�ܻ�	�۫��)3�7�]ɮ=���#�Lv�N�>��+㻙Q��n�޴�䆌wfI���J�W�v��`�$�_j�(��'�ad��M(��}n���}���V�X�Q۽��cfN�ˁd��Bv��vLᗶ��N�i��O1)͓�*���&������D)�'�v���))I;���'y��n.*�F��Wt�ک���z���gz�Hή�0���B�\l����=�jR<un��9{X��wuJ�t������0v.l�پۑs�QK`�ც����h�_g����i�N{Y���g�ݔ|��d����nj�F)V�c��ީ�hN�k��5{Y3Ϊ��A��׷�����jis�M!�v�����n�;*m#faƧe7����$�/\<��!w�N��"��+*�7�l��g�"�A�A�om�%t�����<�^+ݹ�h��#X����҇:Oj9�2�[��mu�t�u4�����W��YS���8�~���z�]��{V�j���7�:zu�㎧�Պ��=I<���z���4�{W��~�ih����˜`��8|��K����܃��%x�Kڙ��=����.�.ͯ��d�Ս�*ߵ��ѽ�W7��9����K�z��_�]�{9��x���9����
��k3B���� �Q%�}.5W��q���8k����KO�^�A�s�-�J�z��vfm-�T�s(:Ӆ�/�=W�;�oc5�䜠���wY������y���F�іU/��tCI}'S�����^E��C����K�3��^�_=���.R��_j�1��Tײ��Cd�7��l�i*ʛŚ��W�_[�ˎ|]���I:�Ϸ$�7�.�o�s���=��sՊr?_�D�w�_���Шm�+�snj˛��4�H�%�ݸ-��i{j{7�%��	�v�𽮗qbe2������ڻ)��6�σ�zQ��==���Cx�+S�]�Ϝ7���Ofq��+1=�͕ɂi]�\,�Iv����c
NT��c��U|c��'I��ۭ:���*&VVVo̆�(T��ײӾ��sB���)���Ѹ{�s�v��N9ƭ<�w ��}X�'ZF����i���}���~W	*���Ė�W׏K��Nc�ݬ/���5�k��H�ݵ�Z���C���Jf�Uݗ�3E�傟%�*{���.��Ҿ���i�R�2b�����v�]b����Y�CƓA�jʸ9f�p#�=&(��.�ٕ٢m.�KG
����::���-��!N�ؾ�_Ot4�Mu�����}�v���S�_p�7����ҟj��7[�dT�=��������Og
l��?��fs�Z1RC±Smr���G�2%ɉ=��5��!:;��hw������ɬ�.��������~��;�h�s�{ӣ5i�A�C#���綧��5�:��B�����=�R��M��q�w2��~�.@=;��%�U��,�r���c��}c���yaJh�2=�t괫
Ͳ�1�-������l��*sK���k���R�n����
���,���A�n*q�ׇD�a�j>So5aC�'�.<*���؃��	0���#OBĻ[�oDN����V�f�m|���YФ�N�����7��L���B�v��>h��>n2�Š!�CtTN1=ۊ;�z3Z�fW	9�@ek����]��/�^x}M�v2˨_j�6�]�c�)��fcuF��.�~ӛ'|�j
[�[��y��=᎗��	���I�f�����}��y�'}�TjiXw�û�O:�[Tr.�זF����hp7L��<���`'�R�ް��-Z�r��~��ד�R���y!l;a\#q1	�ӟi��s}8�9OZp��r�o ������	�U5�I���c�n'�qq���
��f�"�|R��v(櫥�9�v��y�=z����f�C_���-gK�/�^Z���g�'���aL���աuG�GOV=hN=�ꚕ�y=t6�t�����SWR�ICڹB�v0����b�	b��!�5�s�{Қ���:�{:�d��{�Ž�/J0򒎩�Ս��F�+l���6�ً��h������ �ʶ��m�:N��m9�����:`��6l$>[�85:�_���N�r�gf˻�s�c�}���F���Ӽ,B����ɫ�-���T���x�Hަ+�-��:<z-Y7��{����8m�5�R��F'���έ����n��yo��S�-C���R�5x�g�V���Xsk=�uz����B��n�[�n�C�x��R�\*y��~U�vhn�AW �/O���r_�����
V_������oo�Z���Md���s>��Z�٣�"'c򎇏�+�l�
�'D��(��[��8k��)��հ2�Kɔ��G��;�V�e[a�l� pj4F�I�j��)O���k<�}-5֪O`V��^�{8Ϫ��_k���O��RW�)����oqiV~9=�2��gh	t^>��*K>�T�d��%0���������1B����[�G:v��+m�˲����~<*g���f�S%W�!m|#{%c��m3S�+q��9����|��a��;At �ޮ�6g�1��Z�s��H�S/��>���l��p�ͫյ�ʺQ��DgSk��9�3hlӌ�c~G<{�d�au9 �mۧ����F��e����{�u.q���ݷ�i����fU���(��xt*��� p�!ĝՏ9�a���P�cP�YS\S%��_P��yW�ǹ����m^�#sC�Kjk�I�Ž�����nLn2��F�ö����]�9^*9�q5�/N��U4���|یh����ǵ�v3�.�m?fnH��rJ5�6ck�G�"���|�f����^�����}���_aps3��\�}�cڞ�7_��]v!�k��p�:Bj��G8���Z����O�,��nv�f8�q�,��vz�����Chd�oMs�Td9��c��f��:z&ް�Dҵ�↥�Ns/］�~����sχ��Zì����7uy��������h����Ko}.�.!���<�N�EXݗ{�׭ǔ�Ħ�B\�����qC��gD�nwK��+�=�t6}�5��)��z��9
=�3�`'����%F�Y)\an�#���yZ��\b�\���ӻ��ނ\��v���x���l���z�H��B�;�n��Sr���ܜ:���+^���{5��7��*y]�����uk���f�D0�N]Z��␛�A�ǡ�����R�)Щ^D����b*��rj�����3���VG]�����gjRW>gr�`���Q�ڐ�s)�j\s{�An.r���%�3��gk���r�)���~e/�dA�#tL�DI���)�m�S�*��ֲ��r�'놼���eE�<\���t��0c!(�g�τW�����Q��V�M]�f������7�=�ύ����:�}�n��DK]h�w����&�R^�����54��h6�0�d	�Pۅ-y4o#!ë�K�3>���5+=5����
��)�}��B��!l�5��i�k3�qu$+�r*�ɋ�1؄Z��/��r�z�]������کΜ��c��+�Ή[��D����-|��];_]�.�N6��}(=}u�L��ҋO%��Y)�S�%[<p��_wK__U������<�mT�tm��ԅ<��cy�&V�0ә�~��^<^�#yT�_m�A��Y�5N*�u�g_K�By�_=k�k&u����3�/���^+��ޣ�p�O����f�& ���+b�ݞā\���x1��Ab��->�-t<�6�/V���,�j�Pa_���i	�oF��]��G-�SF�t5�ݰ	z��1�m®�J��|:�=��5��Y�t�]ݖ�%htŮ��o�c\���/w�Z�u�Wu���B���qz�]Ft�3��{<�*����>7�P���~�%��r���\���`�H�x���:;,C�3�E��t�W��km%]ˏ�w��^f�-�^���d����*5b�i��v�*�{��=JG,�]��_Oo]|��P�}*���C�_I�F�F�v`ĜY��f��*���w:õ�ᶹ�����QX�'"F�^ �Z��[y�έ��7^+^��)��k}�8����St݌�Ȩ�O��z�f*7����P"6ā��B6�\���5v>��wE�����:�i�T�ݍ�,�u�%"0��`/527�F��:�Ś���"�9�{��}�*��ٽ�:��L�摯���D�.Z���o!��I��y0�;a�#q?'l>S�֑��c�G���ٖ|p�����εq�O\��@e,��)����ަX{����a�1���\�Ɵ���
�l1�gL}�hu�.�۝aqt8V�
8˧Y-�]��vD{��� �U�����=��f
�q:�u��#��t���N��g0��^��V�Dn�q����.�b��2u�wVb�C2'��{���:�y]Lv��\��)�/�݃N33�\�vi<�tr2��릱I
�;�B����Y��m��belٶ�❊8�h���PD�61�#�ü�.{�Е�_hȕ�9���c��h��(��;v"t��nN��@T�͊+N�C��C����E\�n����
[7���ZҒKM�X��1��]Z���,�����1*�w>��h�M*fef�6M�#]1�v7AW=�+]��)����͇\��vV��wf��uly� �pԴ�C�KS��k#+o1���n�m�-�o���:��]�s��X��>�;��"q�_ {'V�BWD�Wn����ѯ�d�z��/�N;�� ޙJ螑F�6oX��qb�3J�Tw��j�mۺ4Yt��»��XM�g^
Tέ��)�4��ѝX���P����J}���i��y��.)	W�����E��¦]"�K|)n��o+��1�d�yk9�
�췵�`B���9�]��=��S�nװ�9�g����9n#+hRx�HTgumN��-��1��V�O�}cp�p�8Y��	�N��WV��]BIJ�%�J瀚)�ib�dA{�91�v���E�x���vѭ��8�T���.gSy`cw��ݼ�|������D[�*Vu��7i��խ	Amdo�,#O�Wl�VWC���d��c���k�a����{)����ᫎ��T��0+n�ȝ"�o
2����^$c.�Kd`�l_�V;T*���/K�t��v���£ʚ�nM�q�Nl�М���qm6O��|�6�g��7�H�����^��Жf�:���!�����ȫ��v6oXq�2��5���bZ��i�9W+�Y8Q{��`ǚ]mlL.O0�_��:�d��}AY�Nﺞ=�������gf���})&��PѮ�Z덽,��Y��p�+p�����u��I�wPTj����a{l��٦�\u�W��p���d��[fS8��]�Kc)�&����W�����v�Z�2�/�m�+n��^�]�梲U�_
U�z;ԇ��J��x��yn���l��k�w+v���}7�miz����f=������zmeugj9�w�!$�>u�ٓh�e�q�ów�Q��M�t5�\�V*�Р��[j���}O������S�ub�Mv����CS��� �-C{/��Guv4���{RI�8��H�؉h��:q�ә4o=�x."�6���Q�V���cZS���w��I�LX��y�F�k���
[:T�F��g�c�|�ˮ{����I�)S����4����p	w	Ը����rrL��5�wٚ�uKWJ���q�w}|����#b���4D[EhѣV���6��f��T`�2ڒ�A���f���D���,Ah1�&��h�J(��h�1�}k�qq�j-Ʈ5,cqTg�+����T������Q��8�Tk�8X�� L<�}K�Zau��pj8������=�����r����u����:ٝ��W|�=���htd��'?��&ns���M��"ℙ�����8;�_P�B@�'��������;��܆e�]���]��	�r��?<Uՙ�V�(wp�C:Z�M��4v������60l��Cz��mO>��~	��Y��;=^Ny��xܮ.��t9w����Q�ǩ�̞�K��g��^߰�mg(h=����L����Fᓔh(9;�5w�SM�b�y��+6Jr�˷!=q�.�g��8Ɏ�%�]��o.\�2����CS�j�X�+KG��X��f���y�3	�G��^��KX"��\j���<�oʾ�Y;qV7h���|X���=V����2-7=�۳4�Qz���*/Pnw���:����5r�������)���ДO��}�%�+VE)[qܰ>��|6��޺/4p�Cr�fn��5��ꁙ&�{�!�P��JDn��k\�ޫ8v��Ϥ#V���J�-�Y��Sg
ɽ�z��J��"*o"�(������j�J;|:��wJ[����KQ+Ԗ'��!���=��i{���3�E�c_�b�a�u��13v�0���VU����!5|rμŚ*�7�4F�_΁k8iËl��5�_E������b;uIր����{.ëQ۔0��|�ۉ�g?OG����t�'%��g�0�J$b{6k�׀�a+��4�5N�97o���7�x<���K�k�2V�� F�f&��U_�V�g�sO���T����}�֭j��v�b��'nk�S.j#H[z�]iۖbw�;�=�<R��9�P��H�B[SQ�0ḷ�#q)���嬋d��^�W�6��[9�摬��o˔�����C_���6���G��s�R�ڌ�6�y�bFmA��u�y�'W��7��{X���(y&�3��Wg����6���/�d�����\4���:��I;=�`��í���}�3�����{��˦�|!��1��j\l���=����{]��k�}p����>?L��~������R���8�+J�o��i�=r�i�Qk}�8j��+@�{�\c���{	�a؞Ӛk�p������K�u�Ь�#G� 5-���x�E��Nn:���W���|k�����޽��%�s��V�\�e�����m�$C�ל5m�e�C�gG6Ɣ:�g��SX
�����L��bn��Q�bȶ����k�F�K���A�܄2{8T)m��e�y��wc̟!��{��1��ɣH���rS;p<�;��mK��Q7�[�|�z���!�C��pz�k���֕Ꙗ�>��j=�7�#�.��6�v���T�w1���oa�k��}r�r->~��29N6���w2����v���pzq�9����}�:S���k��0Gg<�_í�6��Go��6/��bH<�����fo�/2ঘJ}��m�Ŗ�y��=���.Rσ������<�*���o�Z����2�V��Xy?o�;��W�7�=�{���dK�iL������c���Ŭ��~S���_K���-��Q��a�ô)��E����y�9�x����.�?�������g����nhT���އp.�����=�ط��	]��ml!��V�4vܡ;�Pz�]����7���V���c�0�D���_�N8����e퍫$G��f/�K,x�ؿg#�TK=��0s���gh�+t�J��
<�]���^a���թ\�%G���'�����Y�)�ý)^�{R;bڎť!�y6���,>��o�r�מ������-���];_B�B.��#����vZ�ׄ����g��if�9e�*�DZ�о�������;�V���͉vg�<Iz��-��*v�O�'���gP}<m񿷕N����U��^�u�V�����zC�Sq��n��|wϠ���O��H�~j��wF,/w�-��[e-��b��ؾ��Q[��u#:^��OQ���}��͜y$�q'��o���y��{�9ATc_��x|q��^��Q_S�vdΘ��x-�yg���]��s��6g�j�,��s(t�|j��!:3d0�~Kc9�;�u�n�����{r��S��S�n�꛰�܍��g���Zj�Ĳ��ԭ����/ki�ؽ�l�ޗ}{Y3M
>��㋠@��ț�p+�`jd=x�ziJ~��Ʒ�c�O(�{}�o=�By�s�ND��#+���:
�k,0h>��rD��f=QF�Z�����j�T|;��*�\�ۺJ'1�[�;�ƴ��ȯ6�3a_=��v@�Wϩ�7P�V�f���{��˽�|2�LA�5�k��A������F�+Qޭ���#�s0�k/j='���dT�Fkٸ��w�$%����Cy�J����F��N��9��`���q�%���a	D��,��`Z�ݛY��׫�����y���䊜������v�)������0٩Y�Bc2u�i�$iMcƧvFH��Rᷡ�@vôn'��iϴ��2��2O���[�Wcy���]�O|�Ȼ��7qJ�މ_sq�Ѹ���������~� ������aã�Z?c���M<jOnr�vN�hgKB�1:E�����鷙��v��羳嶓܉nr�/�V�<j��3�Ûr����	����n���bs<Ea�v_�zmZ]���r��w��Z���Vmq���d
���_����({���f�[[���8m�?�jZ�s��WE��X6ӧ�o��{\zg[��[��ט�T���;B/#�n���
"m߮��L�Ny������]b,֎N�����S�bl^���ƪo9�M��K�#��Y� �Ŭ֢,+燇>�x�V��p�8�5,�{�^w��R��.���t����'7�����6�rz�#W��wv��,˪۫�uL�v�ԧZ_.�L��+�bec�����9�է1���u�s�m�PU��=2x:��������|h���!:;9�Ή�A���oK��>��5�d���S6��br�)kv <���@)T��/U¹\i�x�^�y���y�2c��·/��<�v�ɚp2ʭ�����I�j��)��d�^B����S���3a��y���䩻eR�T��?@J&\��^�5��g�\	���a��ֿu�zX[�НXW�v~���f	�ŲD�ż��suR��>�ʗ�z�i/�f���>��t�|�J����
�^���:�vn{�j�D����oC��l�L'nk�2�+u��u�mF�3�#Q�!LS��=�P{�^B����Ra�qoQ��471�l��"s�V�S��n���)둗Ϸvg�;��*�N���l
�Ņ��$>��2H�{�o���^o��L&@F�ջ��k��h�ᚐw�e���_������T�Zڣ�y�=7��V���ˠ�	J�Gݙ4��;�4�ѫ�w�3����]���21~�7ړӤ�yx�S�A�兇��nη���Mxi��(<ڃ�ڇZ��:����O'Ұmݱ�6T���nrv��Pl�}wå
����pe!|#v8oP���bI��X���_h<�����Iw��k�9g;�y��s��.�l�=��k�R&6%,W��-�ղ����k��R��ɜ�Cg�hoM����R�\6�����.)6�V�Q���-��f���h����/�-�s^�|߷/1ҵ{��c�E�j�!^,�:���|��Ĺ��T-����oV�>��zLL	׃��5jⵍ���I����&K��v�y��t���b�VzJ�_m���d�Vײ5k�I����+ڬg�܈��٦7\���+9�nJ�����i����}^�~���߼�3^���O>�y�_�\�$���o[],�[�Û�q�yf������>�����W�=���f���!�`�.�B��x<�ۃ@���nHԯJ���*�e�ѹ��G�|3�Vww�JIW����3C׹�TWE�������;lɖ�V�g�$g����Lh$�)
�JݏJ���=�q�fZ��{�N�Ѻ��AQѲ�_��L�����ȭbnnw6�?�:���9����|��m+�o7���9Q<�؜�󊰎�s�tqtM�}w?@��k&�c���[����M+�w��SC�����9n��n�W3���������ky�����u�36qӂk};���BQz���n�F\����{����8x��C�:^y�:�f�?:�a��*����n1�3�q蟵ەp)�@�u;�W���ZS��T�;��v%k������ff��߇J��DZ���eW��l�[{�O|Iٽ�ܹ��X��%�Bu�O�~�5[_^O]���x�|N����p0��Q��ld�t&"_|q�Po��򵫨Q�>33��ޞ>��/����[�9�����ed���-���8���\ߗQ�-}3��b����T��������}�������)��!�7�8����A��ת?oTzhv�6�L��a���\��"m#��c2��w�S�B�'ل�U"�v/Dz���\�����ģ �@�R�5���R�63�8;�4����y��넦fMnS��L�.eC�����<]�q�s��|�Ac�����=���G"jSh�qݯl���W��=�)�;�^����_CV���Y�]� "������X���q�V��\M�I�&��KO/��SyŜ~�w2��w;������1��*��s+]�+�5�߯5�󅍧�S��e�q�ST�8���� ����ۂO��7���������(>�����Ӝ�Y�ö)��te@g����bkٸ'|�k���V�#V���g�
ݭ^�z�v�(<HeDJ�i9.�_50#!(��Յ���s&�Z���-�J��]��2�~���M�El�)�����]1}雜�����E�G�s�u��K��a�Z�7�����7	�����Gk��&E��p��٧���^]�^�{��)Y��+��զ���BF;s��V�=����S�X��^���9O\��V�g)��g;�E��s�z�9�'�ھ�,Ǒ�M�&p��V˻�x���b=��T1P�+"-�HN�yZ�������w;s�\3k�����
ҫ��kr@��� p���fsoq�Wo��}6,�`[�ڬms���ˎ*��i3_�#����txXᳰ�X���=����֝�&-�RwAWa�؋���m	��W�Bj��e���Óg�����P����z�g�8��usO@������J���u�_H��'�׻:�:t�tdy�f߾oӏ�{�^k{�b?Eih�^\�!=sg�AtDQ>\�����x���=�~��R�six�g��}�nE��?yL�K�<�wL�Յ�%s^�o�9��=���o�>���Y'�nO�okƕ�f��;���nԞ�'��粃:+6;�7�������x��0+�
hR|�8<��S*'�dv��蠦wM%>�n�CDi�gD������`쎞����5��N�O����kѬF5>4�$�3O*�qe�T���~yqW-�aؽ|2�����krum��^0��Fu ��y�#/��zϤ�r NjN����ِC��,��z��)�*W���N��WD����!�;~�2zi���Bxۂu l70=M]�i�'���̾�����M�2���R(�j�S��n��(�����;�S�N�j:�\h�b�܅4��F�F����oǪș%�{@���s�Q�����)�I�sf��kh�gs|�c{�_��\��v]G����.�c��)r�V�_F�n�-\z�
��vһ1����;��-]e���%;��ԍ������x�*�:�NdMPN�Rz��@��t7n�����%���W7\�rS�1�H\��/OE0���e�*V&�6��' o(l(oJ��mD�
�W�t�Z�[p���2+0�w��rL���5R��zV�`�R`ɮ�`�++��m��ml�C��ne��ת���l��
�L�`�r��u�w��l�ǵv4��aou�� ��a<̩���ʹ��4��1�痉<ҫX���X�열����x�n�6�Ynp��j�>�t�Z:���,�|��(P�%h+��>��7������E��X�;-����5���t�-��hko�Jk�\����^�[Ҟ2�!B��R�&�H��ʓJN�+gW;��bL@�"�fP�{V�us�l��(��>a҅�0e����Y��.�k[t	�m�=u��]7�;�nt��r��Ķ�j�焢P��we���ֹ��8ֺd��yt���G���i�A���:�.��ϟ^'8[�j��*��a�MZ��!YY���[��)�o諤��]��b�j*ӊ�ǣ�'_ԉ�]4��54����Vg'�αCb�kB]P�=����\���#�Mi�wy�� λ�B�]�2k,�m��n��I��5��SA���]�bV ���2PI�Yz�wV�V\+ؗ��+즃C3�E-F(�Ӫ�Z�Wx�).��'�T<@�Q'J�n�ӌۻ���(���_ph��}[MT��-�	�֊���:�nD�d��I\9Q�Z�[�Y{��lj�
a�.�n��?f��j�l�̦](��#{D�]�dK�w^,[8Lt�qܶc�6K.:t@��b��涻^g-F�7(���R���a����Ӭ�Ne@ug];� ��ݎ{��q�=.s�\���ܣ9^�j��4�GlY��i�`82��w_S��^�AHяkH�V��:
�m��u���
Es�kQm+Ш�"�e_��*�^�h$�9���9�jo;�W+�-��D�G�X�:�&;D�/�&�`ڱ�[�Z'u{�M�/c
������_R/%>]K�pf<=z�n�[4��ei�c�뺣��*W)����S����{`���ُ���{�v��p�Xn�L:k��;g\���uAp̷n�wE���Q�W��p�$l,ٔƲ�ʲ��$�z�ݾ6W��t��-�wwD,9��.y�El�L��$�K����E.����pyt��*ˉ��t�Lv��5���$]�ƙ:�	(z���t�;�D���fJۧ��;]ԩ��k{�R���g%p㺧{�Ϩ
��
�h�Y1�i"�Ӝ�q�9�9[�Nr��sq��h��Ƹ�(��"�[�\E�9�n5��q�sEqq��pXM�!��#C��9̀��h�Y!�\qmq���1�k�s���n1b$ы`��qs���*�р$ɰ��q��q�� (�@b���9�" ����8\���>��֗Άa����Q5;善qk`�����Ycgv���$���>�఻Y�iK�5의(��,e"g��K�9s����_������w��ő�'�]�1�y^�6�Ͻ�P����f(rJx֩1ڟ�f\��0�r�����k��׳B✶s��W�6�v����>,K�y���!�~��{6�чφecu,h���G�d�eD��qu�-d��KKU�Ŷ��\Bn���ç��u����Z�����߄�z�;���Q@��FT�y>�Q|r�*[�^��ʑb�����M��w뼮Z^�c��00�C3C.>ތ���fU�a�r�/+�_zϰ�s'�$��͉���?,��.g�x�Uac���k��LN�;����3w�F����8׫�y=�B�z~n���ݛ�D��g�լ�z�i�'�K����N��Y��}ư��'.g�V��4�x7=y�8~f�1�\����}s����C���z����\R���1�~��m|x�{�yh���,^G��&s��քN��PNU�]1�L	�v��]�u]�+>����:�^�pqg�_/<�p���O!�T�DY�)W�G�Fq���At�v�ZQ��g�B{�}�^q=9>A���s�b*(�R:~�{{��|�M��O�e^���� �7��ͮ��b���#�躴��Wm��D��,�����I4����q���n��j���gj�9q	[d]]f����m�ѵ��Rr��Jv�%��x��R��eg�����v��T��գ�<�
�$��%�FUC�3��3=�a��	�ޅ^t�ʮ����v��8��P��Z��yh?����IU�L�9T;��nbR�w�׫ga��a)��^=�4�\-��>ޑ���#�w��c��ށ��,�8 &��a��N9Q27׹��9^LI)9�~u��t����m���;q�냓�L��ީ�;�Ф�vaS�B��
��>r�AR���,jέr�;�m���ݝq:O��}a�O��V:]=aD�N�OF���� 5B@�%:�7^��@�j�f��.�l{��H�08�{v�`E�N:�B�}��=U`��?D۪��@��؂c���f;Whw��Ď7��VR�\m�58���u�I죞R�|:���k�w]p9���'��ٱ_K��W�K�r*ڜ	��N�<��)xkTw_�7��wF��&��wu����F�"�W�˦�h�Q��eE��y<2e���Nt�J*<r�Vu����g��8vx/#O���롗�Cٽ���� �z.���Bɗ�ۯ�s]"�=�d&��Y��
2��05E0mڠ�;*W��r�fPѸ�	�q�P����@ҥ���u�P��Յ�b�O�r�]c��Ʀ��{­��Y�wMҺ7y���:/�fI�o];���H�����`�6_�/�qԧl�O%��ǐ��q��٫��g�3���+�q����7��Ǯ�*{8�H���Y�ڢn��װ����]��]�K�A�'\�owӱ�Z���跞J3ٜû��+��;���n��>�:�M+7_�)�&<��3���U:�S�f��<��/<��"=2�=�}����/9֣��R�غ�g�Fq�L����9�ժ\nH̭õժ+�[��,�Q�Ը�dw�;���j�w˳�g9�Z�J%��ΆtF?/7���ꉩF�{:��oU�bQ�D-������Q��S��+��v'5�^��L��$����fb��X��u�.':���迪z�]T���?MX��x(ގ�3�gPgn;��o��g�"������f��P3%Ϗ��(�@E#�S(.v��}x=�k�Y��*��.�w{�ex25C>�t��y[Q���T�l�	ј�[�*���a鯖v�UĶ�����_[�ױ{kܙ֧�}Dl�S�>���� s��F����/OTzd�8	�eY�}X�G��u��<p�`�T�[zݒ�o4G��ofA�.���\���E�zc
{�셣"��I8|�ҫ056rtq,5�Mw
�f�\SD��,��ʔ6�C/��ӌI������>��O��혷C�K̥���2-���j��^ŪuI�ؕ�������u��|f��T�.Ij@|R��x���v�F�:�ᷪ�;|pg�������O"x�O��bl}^�C����!��{C�x�uV3�H񪞡���4.+e���5��C�����}f��wO@�bb�zE�)G�[Q���'FT�hׄT��8�=��O��L�>ܻ�a.���u�����:l#�ע�j.GR�fiM��F���j/C��td�EH�؜��+�0����L`�����g���uW)ߔ��/z�yF],��f���=9,w�FV��PߵmAq�5�7ht��d?����{e�T�����]����׻G}�U�O��u�q�3±go�_ϽYF����t&y�}7C�ҳ��2O��_�b���4K=�"�N�+���=7��C3%٭<��{�M��3��]j��:���李�4}�r\��l�l�X
���j�\`y�_qY���w^3�*�
ϟR�|�9���9t�/����'��rW&�/aw y1�»��s��cֲٙ��uZ�JV�K�휈��u�����L�0gN�(@��r��{h(�
V݋�m��<������\6����9S�H�˧�ko_�^t�.�׻�L���x��J��q�)og�������7���O�ve���\�8R};�C#wFh���S��-�@��N/5�ig�Wm->���_�:�)L�J}�s�������/� ���{p�Ԏ(^���D5h->�YH?�K,"K�1�&*�te�3��,}tz��j���VQy�q~����==�wN�3���T����ށ��.܀��N�?������u����0�4���������*�������H÷�2�ٛ}T'�Âu oNlh~��P�D����]{g�p9�xW��4�kC�K�lǺ}���ǧp�����r���s3,��h�]����kj쎬p̎"�H�ZsB�x�
�m��5|��Vx�������@�����~�5�h�ۑ\�x	̭謓*�|�Hj�혩�qZɫ��c��!�m]�M��¶'`f�͖�޽C֫<�hTXǮB~��h�<�ڐ{%������:���נ��~�P+����;=i��m����_��2=�oF\
]^3*� ��;���t^�x)�����::i���w������]w������bsc��m��3w�@h�x+8��9;szb���b|�Z��hOd`b�ڹ�1pݞ�W�.����Է�Ls[(��K6�*���K��c�>z��7�jͬ�Ζ�����(���gϜǚhn��Ki��tG\O��GJ=K/�ܸ&��Xv�xU�k�ttc�p ���շP�:�aƪ�����2��n��৸�7S5��I���>�\s�xN~�Y��w��������Wtz��P�8c��(�_��n(������^�:Է��9z���+�v��VY>��k���n�ȡ�q�n\N��S=��'2����f|r)��)���1W.�4��N���
���d�u=r��o��]�ii�,����3�u����T8/Dat����B��	��v�9��v75�(=讴8o�e�o�]�IF�$�j��tg���&V��Zg0}��LyVj���X��<,��,_Lx����}\��^Z�g$�P$�p�H6��;B�˾g����高��OW��н5�սw��ޑ���gH��������l�K6��������ɶgug%"k���z �b�g�O��`��n���󭣜��ۏw\��fVss�qً"�v6���De�N������=��r��X�Yף���������}��Z���a6 �F��*uF�����S{SS���D�WVѺ/Og�L5P���{�]u��^�-���Ӏ����\"A[��t��J�����W�R�0ڇ�VoS�}�w��*�ܮz�ԛ4�)�ΰ�Ὧ�����`�+��@.=����ϟYƲN�����x�B]/CsN�њt�l��Y�$'T�.��D,�8�<���练;�2�������ĿG�ǉ��+��'��MIyM}�I�4	�3��^F��T�|NL_mm)S>��r��O^�#�{��wu {�:����޾��T�D)��l�ب����5���/�֓>�W��>��aXk��J���_F�;����5C/z�K�éϠ��Y$�ch������oEO��u�HU�Oa��W��K�ч��_�X;}�C.7�a�/���]�̼��'�X��MtLv\|2�m�R�࿫�	ˌ�:�����S�p��P]>Κ�;~��N8mmixjat�-!s����9�&XΘ&ھ��#�ϰ����^��z�VA Տ���Rc�����f�_��V/���߫�����n����{�M+4�F3���w(��Ml�{��az�8��8���Nwe ���/��[EQ�P�L���B��G�
=��0�i�*�"�ys��,n�=�.=Y޸�+�j�w�.�1��((�$�K��^�t�v�F�NmO(�F�x\��bQ��q~�OT
�Ϭ��/�q��[����7ea�]{ć]Rw�O��9��[4sJxF�����pcZ��f
��ٓd��~��eC���O��Vgo|��X���A�U2%X=�ck���ys����i_�����b�*< ���-���C&"&�4˭r�a�s����X+�f����' ����:��&�u����`�?�>�RU<��2n>��z:��gPgn;�C�Fl��?Pz��Z�,!�F�<XD��3�L�"���n*e�����>��{\�u�K R���}7�iz�6���[8'�*u��7�	������R�0������U�J�����Eu�9��;��F���#6+�؛��S�l�9�4�ź�Qe����>��l��Cy���=�*}M���x�Vp�� ����.fd���� w����;��=�7�rz�uN#�= �+4L=���Ǒ<_ǧ�O16?'�b�&����7�x��C���"9"�z�T��4.)��X_�}�D;��T��7��Q��O�g�Pc�����ة�ə��h
��deʣ�𹄠�����,��x�����B]wB�u���ei��!��²���W��5�=�V�8ʈC9ѓ��dv/+�_#�}�E���l;�G���;=siFs����g�w�<U?*����J��󶡼�mAq�4�+_��S>�p�^B�~l�Й��u���Y3�0�VR�;�e���6�YC+�t3�(�}���8n��oMbFs�vA¶^��.}ζ��6��î�������nVh콨G��D�^	O�\ay��n�p�o���Z��2+�$4��l�f��1�{���w��������U]��:��9R�,b����Z6�ٸ6n�y�}7�8�]�⋛{э�=zz(��@Ŝ�9ɕ�=8��we�^U�k�9���O����8��uC�k`�f�i�=g����Ȋ�M�`uѫ�q��]}�du��w�׌Ƹ� V	��7�}��R�-���r�O�|g�����yd2�d����Lu���wӹ�gfr�q%Vin�S��e_���^,Q�N�d{JutW�gt�J}ϝ(��yT0Ŋ��2.
p*_/9q����rg{]�}��is�A����f�Iu�����l�(.=ՏW`�-�k��J�gJZ/&�+��w�}�G9�Fu ��v*���wýg�[ �bN���>��@�����r]Y�2�gм��t�_>��Ϥa�wQ��f_Ϫ���0:*�m�T�z�f�-[�ꦸ�����R�@zvmh~�}m��{\�=;��uD�~���#[;f���Q�:��O	��uӧ�RF��$��MS��8-��d;�{k�����������9�|σ3tu�և��;�h �575��M*���=o��q���.����ۮ��͒�t撓Z��*(\�xcF��7If;3�O�<5c��+P�q>�w7�1ˮ�S�y?Dnr֭a�q�X���iz5�;��S��s���2��eG�����
3S�Y;��߄����*�+Q�Lv�NQ	�^Fc�ʿ��G���1�C�j�4��~���m۞	�{˙7�<���9�z�TB�_Q�FI�4r�Sخ��x���Y�O�`w"o(��\��a�c�����GgP]��a�����hE�3;BGa�r�y]�Y�3Ϣ�Uu�f��i����z//�S�¡�PF��LN���m���L��� Q@��k�1�hwq4��m���Ք�\T�'��������*��0�D��uW	�G��{�����a��~�]��|�z��펐��p58N�t�T��	���2X�ۆ5U'�u׬�����7K��?��������g�� ��񗜋�2��2���.r�@꽍��|Y�x�s�!�{ܓ����t��)�{t������?3����F��Xʡ�/x`�>��f꯲3=j:���V�MdGz�r�u��|�-��.���$�_D��*a�<��d`ݳ�LVo���p��E���K�_�|�˿Lx��������_���IwP$��g@Q��;Wظ�����Q���X�!b������]1vp^�oZ���q�z~D.9g��	���(�eNzm`�uȎ��N�����@V�g���γYYu S�/U���ߚΛ�E�)j�L�}���� 1-?
�u1�tt�+3f�V;�m;�7�F��C���d��ԑ�Mc�gV�S����>7k)98��Le(^�Դ"Ā�,ңV2�,HwM�w�s�t��Ԩ��$(o_wR�iD�WSǎs[I�>x���v0�5��e���-��Y�]��:����Kޣ��b���;����V7��٭&t�ͭ�qK*�r��m�n�	dro��Ø���K��"��w�JZ\��0��2,N����{��5J{���,h�HT�&�=�pX���Qa�ع�����N�j�_ҵ���|AiÂ�ӟWoX��[�V��;���O'�=���t��(� ���=��S����6�+�uv�U�g�����d�l�u!ܕ*�I��]�iu��PȯkQP��ԭS��̧r
�� �Hː��]$�B�t��V�J�`��=����W��a<�$��8�.�^��'e!-Ll�H]m��0G.����,bl�)�w��=�)MSe*-��բ��幆�<lgB7xU�X�S��ũ!*�ϝlN��Yǘ�g|L��{���*�*�B�)��f�|XT�Q5cʄ��{M�<+u�c2�̵���@�NJJZa**=T�bέu���ʀ�֬]tt�,�Á��(��Pr˸�ݎZC���.yڮ�CV��[�]�غ��&��:�g\r����3W]X]w����s�|���,Z�>7b�\	L�N��-J�����ʙ�]�nf���2&�N�����͎Y�n^�K��oc�Rk7Ӟ":N����5t���>�eլ}��ԃ�Gv��;�Z��x�Z��i���b���7���r�w!roZ�f؆dJ}���v�A�|Zs"�ˬ]�9Ŏ+��m���ȭy���34^ȩ's�z�m��n�r M��٬�7�m�Ft�k��cqi=g��j�,0:9�6�>��c2�L�w��ƱT��:�d�4�#��fӵ|7O*ZsS�}Z�3�`��.���jn�
�Y���NNZ���'1[�����Ӌð���gPVs�ę����-����y.��R!t�*��r�ߚ�C8�M�<�$g
��� ��˳�L��he(R�R���Y�j���Q��uh�j��q��m5�eXk���X����n��mwB����rR0m]vo׬��.��$ݖ�0.Dk��T!%��ү3�`����Q�l>���vԘ���Q�C/�%�G}�X)U�� �ԥ�@�)�դ$�E�Z��͑4��͘%�F�٘�.<瓘�4�@������]����	H�����i�;o�ﾝ���
"�9�Ƹ���+�\�cQ�%������n.s��$���C�\�������s���q�dĘ���q���+\[�A&L���E%L�M7'5��(cmd��$0A0#	�5��8��%�����d�&s��,A%I���ɒ
4d-��&	�C�9�F�s�(�&&�(s�4�9r�9D���愙�r�q�$%8�E����v����_#�Y�X�F��އ��n��Qv��p�����v<���c��/s����AV�j�]k��_v�b��y��}�5`��_��sf.*U.>��i�����^q�v+��g�z0ؖwy>Ι����o�C����6����b�e>�?:�E�C�?u-/I���u��p�5ʤ��>Ac���8CS6|4��3�6@W)�cYף������m��k�}zo�jFU]��Jgo2zw��۸�u5,�"U@�0WVѐ����Գ|C�=�5B������lu�yvW8�^'�=.8�{��0O������L�ѿ�f��7��(=�����d{���xnw�Q�Tu���}ԁ�|:����޾�U�LZ�<��́(׎��b��S}�Z��u���Q����n����U%�4n#���D3T2��a����s���EՇS��a�
s���q����zסP��*��{�����Eu��.����i�u���Ŋ�U-��BoЌ�0N
#09q�
}g��	��%�˿=��}{�L�Vn��jb�,؁��={�3=����w\V��;��=0M�|d{P7du&���M��,���c�A��ٴd����Y��ʺ�;M��C�̥S��r�E����Z��0e�����(�
�i�me{x�rڙ/�:��h4F*�]X�J�}C�����t{jʆv��;�o��*�{������d[т�.Z��i�V�R�Y����Yd=W�Zyu�tv��Y�����c�*=�6{�}~wJ-��&e�C�4��w����gz��U=[��V6�z@~�6zW��p֧#�)��h\Fs���s�P���Q�C_A���v���I�d�Ny��v�FTat�+�W]Cgz:��c�[�~�h�1[$���^���P���@X9I�"�΍��호����Cٮ/GL��<z��Oq]N��|漎R򧏛O��_C���zphw�υ\�>��_��X��H_�S�ϟ����}�=�Lg��3��=
�(���P�)�i�l���,�>��W�k�jx�$�3�"EA�l�T����(\C�׃ة>5u����~��+������0������7�<n�1�r Ҹ��X옧ڈ��$�����rk�xN���w�pa+��F�U18��zm�9�F���@��5u}0DX-tn��������	�Y����l�7����X���|f��T�-T��lW���2�:���sG_��^�A��^S�n-���y
j��}<��8�ɚ���ď)�������דB��b͹xqX�Q�n$AJ����H0�p�j;pe_5$6m�r�����sw��kGQ��s��/=��>���ѥ���{M�yc3���&�4N���x�$�w��[J�P��t<����@��qE��d5g�����R��՗�.�kef�ޅR���z��s&3(F*�;9�D��*��YY��j��jo���=;���{�(_���E�!�tLw��x��ʢ��s��T����N{_�d��j�1��]�x�L�
�ە�[��7�=�:�� ��7��e@޺2V|.a��'0Þ��Ϩ�=��ckO�X���?]xZۭ��5�}3�:#Wi��j�h)�l��]��oH'���b�G`M{M�nCJ���W�z��_��G�f�/m�*�xJs�x�̱Y���f��k��c���7�vT�Y�rJ���C{�ʬ7G�(�Vr��I��§]�wz�u.�F�ΟeN�v�>SǸz��ǣO2w�P�|&p;�tpK#��F�.�V����u��~���W�zo�὎n}(�=̥��N�=:X���FY��ڰ��+Ɏ�p�I��x�[����'L����<L����F/��.��D��f9�*��R9U<���a�s��&��M-Yc���\�b��9�����lv�C������e]��?U��-��!���5|X����r�;�ݓE�\��暻�u�B����)��]�9�g�K"s��2��y*K5��^`{����Aϼ��d��e��%m��²�9�׵	s��wu�(��wE;�1��[x�Ǜ\Υ�s�#ʕ3�kKgҷ@�E���Z1�ݍ٧�g�_]Bw��+��8�:�zo�T���nKߜ����<�3Q��	�i�{uM������tN�tg�i�/<���$T>ⴾ#�/���}]V��>���U�3���M�Q�j�J��O�"dL���(W�鯡fֆ_Sft�o�s����q9Y�;���(B~�lњw��^r�1�)òHJ�����Nw�{�x*Y�C�M_<{��"6�*�뛛��q��ފs�-%�qA�C��\�y�lɎ�9F*%�u�-d��K_-VC,؉��tmv�>���U���P�R�|:x�|�ǀ}P=�}EO"2�6^�a��("����al�z<��5�-������] ۚ����遅�d{��.�2�����'�ʳ��+�ts�N��x��g�#�{öU]:c7�X_g�G���LN��롶��L��Q[펝�����]����2�|��] ���5g|k+j�=�>�\}�U·���Qwÿl���8<�]Z��GE�$V��0nl���7AKF�ω����?cR�b:z����
�=��I��NF�F)^_Q���dd;c9!OG<��Y����SN��]�1<��ո��a��Q���Ǎ�g�n�+;���	�VG�ي�;_.�îoF:���Θe=X�o-�2Y�+�[h�Xi��s��U��C��lP�<\U���0�X��0������i�o�,��4���d��L	�X���� r�`g����D�:�F��6��0�fݷ��/w�lz���ǽkb�ݔ��,�����y-4�	��7%l���	{{ta����t�w��/WZ7��-��A/��Q���AS�=۫3��3��v��l���Qp;�ٞF����gH�����3�xa~�	���.�r�%{/0X��}���U����D�g��zE>[��晫�����^�Ft�v�\=�Mgڿ4_�X�G����O�d1��C(�1u2�K�>�D�h`�'�m���:FZ�m�tUQ���ĜA�{ˠ�Vݣ��Y�����-�+㲹Mx6�Yף����#Qw�U�5������X���r�&�z��>^Bo��jY�D@j�H&
��7E���	��>#�N�waݟ^�t���,{u���=�>�����_\K���H�-$i�ؼ�-M2�H��{��c\��ͧ"��B�*:�W�m�R�:���f�u�����-L�R����tܜ��mѵ hM!,�}h�;i�ٍ=r��viG��&�j�Lvk3��+Y��^͌2�Td�Q�I�6u���jh�ۯ =��|��;�A2��9o	���Gb��3'j9ڕk��悍�z�txU�%�K���3�2w�t��{�M�q`�����g>�����wtnK�h�wP�f�e�P�m�޵��=�o9I9_Xʹ�7<64�YR�����[���د�.��	�Eu�K�w�Bv���F��r��vR��Ю�C
�V�y�-W�1�����pJ~XNJć^UXc"5Wo�Ӹ����k���y���}��9~Bl��;��x�-�2=�&쎤װ���Z�Y����t}�f��M׻GFUu�>�u˧��۲���_ќ�_Kv�̠���VWפ�Q����#���ξ�{�:h����{yY��qg�=��H/.�B��u�W����]	�e�F�x5�O�=N�_7�~�eW#�z���
�5:\z��q�W�����[
3�e�4Zj�vew�)	$�D��po���S�9	ͽ���|�/�z���w��:�]C���q7_�o�$�oaS�ު7�<i�Aރ:�-/�H]T�r��u�����t��A!�=�P��ֲ�՛�=���kn��q���K7�(��΁0
D�=-����y���q}]7^u��K����3H��{�Si8�M�W�Y�eWs�>��6�v_X��_k�Ǻ�S�v��O.�oYӮ��u_V&�+��k���c��_ul������{\���qtZBe��r����[�)+�	�ܫ�{��Vs���<�5�g~��wk���z��(O��w_\w�o�x�2 'Pf6 n@����n�o��'��s�\�g2�����f�qW�y��w�pa+��u�]v��C�鿙 s��F��.�r�k�K˱؎���ӈ��	�ҳD����>���=� �Vo�����6�K�ڂGg�r�A�@un���@�f�'��{~�_��*�j���>�i>,�_���B��SW��D_y3]�h	��d���GI!o�Ӽh]t�5���F�Q�wF.}f��BN����X��T½7�|^�o�!?(0��P�B�y�#��Ȝd)��>efK_-��`۽�:2�2�ձ��o}��tn������ފ�oFT�%g¤vP��#�/+�H��fhj�"���7�v؟w������c�J��{�8���ٹ���FV��P�yA6����7hs��N`���#�V��R�Zz�q8o�y[\5US�|�p\}��V�;}���E����t�rV���D�����#k�OA��mת��D�q�����8��@R����.�.�F����[��vph�^*w�Z����=��_ Vmb{�z��5w�G���5���}�ƌ(:\��ЊڎT(��n���u���eqc��d�bN=c'�3���t�7\�9l�����J;��WZ,��Z9�����:�kM�Ә�W!��������x]����8#r9M�`,�{�]k�C���>**{���/���Y�V��W�j���쥥�d�pe�T@3�����n)�eF��.��8r�.칺��"����\�b���u!��5�žyu��P�|eSS)��	��DT��ufu�=z�(o}���c��|������lv�|�)ᾩf�D�l�a���ǾO�}���9��g�e����ˊ���ﰮ#��@X{��R2��F��� k�л�u����
��j�TJ�D{�mB6{Ƃ3��_�惹n�!�Ⱗ�0ﻨ�OM31^}G�Y^s�l��������c�`d��
�/M,�����1�}�̎8��>���~����Vh��S����?����	���z���`��x���V�B�jV�
��PrJ��Ǥf�<��{owşK�<���y���R���&;h}�Bؼ�{nU��<���;G����Y�<C������:}~|h8���!�u�kL��1�C��v{��g�G�眷n~�viHۨja=W�����e���k��M�Y�d�W��`���i�\�`�x�*�L.&sӠD%ml�g]��o�_ټ�]��K����E���d�6LVj�n�sO�uJ|o:PNZ�0{{�Y��,K��$W|�ū�	'����k���yly�WF�y�U��|�`��}�p)ux̨�Nzc{f�ƭ�u��d��c&��9gp����WN�1��/��Q�T�9��CnPɛ�]���c=׻��_@Q�U��A���2pm׫�]Oa8n0�7��UMv�'�K��j�V��]�k�w��R��{�\�����s�5�ˤY�:���1O��9+�T���x_5��zh]�M�����^��s귞|}���c=YdP�;����ݙ�O��Rr��9�K��+\ŝW����g�az����{ށ�U�ҳ��7O�����H�E��@��Q�C��:Y����ԃ#�[��K\41N��:���0�Q��wMdw��)�C�(�Yh>~�
��t���nR��{S՜�&}y���^�+¼��qE�\n�0����}�8�{���3�xa~�	�����IW�K�x�6���8�9�	>�b�C��et��ORg��L�7]�G���3��b�{7£��S�Te�s�{��O�)�nW�t	
P09�����|��\�h`�����)�=�k�J1+�Q�]㊂|@<P�+����^�/[ݼ㇫��?&��r^��wZ/)A�(!Zfq��5�fJM9�>�3>[�i���,*VE�A6ov��e
�6�W�-޴�*�洫H�gO8���UC��,��R�_gV<���uf�d���e��^�NS���u���<����	ѐ6d�r�_���:�p0:C��j�5Oڼ�`N��ˢ����c:!�n�~�:n���\��s�D@j��+�h���IoF@��^��Oh,�΋����ŷ��҉�:|7�Հ_���D�:��FIh�#M?9Pw��Ǒ6�jC]nO]����_�P���*�����@�\ �bl��ꯪc�%�V򗫎��
`*<]OA��:�dT�r������m��+���7��������w'�MT	��%�<i[�,��6�)���l<����S��W�d�8��]U�=讣y�%�q�k4����}y��j�eƺfβ	[���T�ߦ����0��_���U��V	�+���	�������3�ј�j�Κ�9~Bl���t�g�	��=�"n��	�i��8x���+�J��v��M�෈�����W^��O�MJs{ku��z��n��#�@�P��vxgH5T�Vpy]���G����'o+����SҸ��kS�ݔ�]���NQ�>%��+>�~�h����v/�0�\x� �D�cl�Չ֭�h�;Sk>�l�U��R����f�*�t{r��X-# �=r�j��۵m�<�옫B.���(�3j|qmpt��,��v4�S���!��� v�%��]��[���Kx:[��*��R�qFyk���7.+ܱg��8�=@*��qn�>�˩�k1�-\�-�f�).�q���DD?V�9�]m�I�㤊6:ct�m+�B��N�4R�K�w�JC/1
�=�v��b��v����tw��Y�
�����E|�h���9��:
� ��K	�T���7����ݤ��@g�u��/�<�w�!���}�PZ���f�S����0[*��ӆe776ww9k��CB��2�L�P�*ՈC�5���&�N�gj�G�k���� �#�n7z��s��sP��q�S�9B��7p+��;r�)�株�G��`=nZ���7Ш���s#w���xv�@-쨕]��� jL�Lڌ�'�
]�r̰�Pz�']���uH��nvې�.r=ٶ�=�_�7�2�z���/7�;�c��#�͵�ٝ��M�bGPm7��9/ښ���Φ�vn�ۈV�-�I�	 +Pe�B�U�Y�WZzƱv�[�Ud�;������n\M�첢�M˷4��KVрw��i�����+Z.�θ�����'h��p3���9��ʻ�\�x!���a��\�t�1�&�`�un~2�ހB9�F�ƀ�r�vۓ9e9V�+nQ�c�
5t�Wi��^a 
Mf�t70������X�ݝܢB�q�on��1G�)�TZ�8둵V�o$�ݎ"�R:Yz��spd��&�d��Wf����
-3���=)
�y�V+�]46���YہU�8\�gv�Ψ��HZ��r���)��[�a���CO�$��e G�
�DpuY-1�L��w�5
\�)扶XF�o:���@��>��\)v&�X��Q��ֺrmf%�Qo9�(w]���]dUˎ�h �e^qn�[ͅ�:��aoq5�^��2��,eY���b���=�C"\E�̧:<e�[�Hu�y��;�,>�;-b�������3�Zs�f�BX�ͺʳQρ�aW�Y(ح�B�Wؘr�UR1�5̣�5�Kub�kwd��v�	֦�"����_s�[m����s���߯w뀕�=�0��.N��C�I"�h�]�+�p�j�+�*g!�uu�v���1Ʋ��*�w[��E���.�OP�:�z�A��*�۸ܔ(�5�zr�w4�>��^�s�əl�T�ܘ �ÑZ��:���g#�^�x���b��qut硱u-�k�Y����ٯ;W� 6��\�x�G0=���L��C=��W�ĘWQ	e�!-���w�PR�-(�a���yd��[Deͬ��}6O;�*��N���ߥ��3�����u���뿕�@������HcNr7"I���#LFS%�	�L�8���d�!�H���9˂DfLT��Hn..r� ��2H��#7)J�7$&�Fe�q�4�8��rJL�0�r�6e9�2Pɰ�&��Zf&D�	��"&���Q8��$�h�K#��q4fLf���� HHdSJ"R"�ɦ��1q����IDl�L���AXIY�����DC����RI�a1s�2!�&���@���L\[�����.�73��13��D���f! �q��%"���C��d����ĘD�3A�C&A}�_�>|���Χ��ѢM�̨����0,�9�9�E��ZDи��t�c�[��3���!�n�$*`�}�؋-n-�I�S��_���]C��U�G@h���0����>W�C�:�[C3|������2�/u����n���y$���
�Ύ����1t�'/L�kOT
�>�Ǩ���;÷5���|�WJ]�[~���~5�;ex�� ��΁?ȱq*�������A��c�p�<׻;��	�a΍ۦ�#y��t8�s��_9��ᾩf�D�Pg@�"EA�l�L��l��e��2}~��o�9=�C�i���B�ef�*�)	�w_\w����zf6�n�Ψ��V)�w�0�vr��e�s��g+�	��cۊ�my��w#��i7�6�ؗ�3Ӱ�����������<��f�YS��Eׄ��K4T;���>=>��re`6�� ���3|��Q;�y8z;@럢:?[GuO�P��*���t�_,�P�U�T>�D��ǧ�O^�~.���F����H�^�F�ʣ�)���mX,��t�5����Q�Wtbk|���r�YB#ʧ/5�	O�����3_�Pag�3��yqR=������\5��*�C����̿#7���:��KO$��i.ԏE�r�[,�R�4�m5/p��R�'��N��#��f��yt�^���"����s<4pǬD�����)�+���3fl�Kz�I�c���Sm�������W"��ݱ�����̦?m��v���Ρ�=ǀ9���z=03{�d�0�Ķ+Ʒ��=�Vd��6���C;��8�њ����
�u��j]����*��GNK����;j�ڂ��c{}�]%���3|9�cq�+�{��Zn�a8oq��/m�}
�����=�,Vy��s�VQ��}޽�E:�s����M��|��L���J>���w�M. y�V��;��$�Г/ޡ�~˷�W�����*x?����:�OQ�S��n#W�]��]k�^:c��<��^5ٗ:������C1��U��N� e�T:X���o�rW&�'v���Q[%�N.Q���wU�E�|+��]�z�����b�|��I[c��2�������=���{�T���t4�Z�a{�������߯�ѝ�sѝ@=�;
�u���cSƇ$�F��`i�\?{�����@��.+��i��Aqv�Q[��B��}��q��e�u��@���ۻ�"L�c�y
��:� }=���
S7FQz|��qWݤC7�a|G�p~��cE����[뉧r���s�ۻ�\�qw} MU�l^(X6I�_���w Yx�<�-����
���cw��䓈����Eu���n�Z�ɒv�|�̳���K}#uۼ��ޡ���HB����^�Kޕ���M=�b�/������階��n^ƪ��3ت�鿔��n�@�҅h/M|�kC����{��|�w��"|έ�;�{+<��U��ӻfE��Y��IA|
�4."�����T�l�u�,K"���D�Gc˓�xtA��x�����ƣ�_TS�=GI!��b����m۔���:ӊ(�^�뺏f��9��%�B���n���<�3q�)�z�R�_Q�d�DmL.�@ZU�[�}3�=O�T��_]��)��ʇ�k�pmMQ^��t���2=�ї�W�ʼ�n��ɟ_�*:��G���;�U�o�=���4�5���]w��HEǺ��ꑕ������{��p��Ѫ�(�@���^�����f����T�Yox-����ɷ!װegtn{1s���p�˧ߋ����ߒ��,�5l��>_�� �e��u��zFM�
�Oۗ>י����8�zW���,��;����ݙ��y.+�Xe�9]E�;�.hk��x���ۯ;k�z����u�}�Hg<�E}gĥfa���@���(��3��~YB���H�X*���n��&hyY��Nt�i�Jf,��47�H{.~hk���{� .:S]p@	^�P5�}~͛$ݻN��S+�V9ڦC&)\��++�u�����u6y
f�7���9��8Uk�X�$�1�ZWJ���[�&v��P�q�U������+�'K�k;�×���u����Az�Q�����w�!�&�h��v�o�=��@L�=�a���+�Αǳ���}\���yh<���R�Wut���zf����w��pI�L�D��C����&}?M3W��a��/O�:C;9{=S�/���eV@������3�U��W�F�Â`�J�nb�e>�|��ޚ�x����/?^~j�"�S�:�4cz{��;q��.+�ه�z������d�vW)�@,l�X�f\��gf�og�����蔺�����t����M���n������.��8�����c;�1�:���7�a:���8Z|��(�@��d���X�{�n����FIh��u��nX���#5�N��-���ʎ�	����/�P<�up9�)�!�:���#ځXn�����^�R(��>95Ob�T��ѫ=e�]C�6���<��Ѹ��7�a�,/b�z�zp<Z[����a��L#�܌���\X]kЬ�7{N�n�,##4�蚾�E��餜���.����.b�BU�g��eu��k��s����E���g��}�\o�\7n�Q1��[�cҶ��	�*m
�\)�����t�PѾ�)h��4�x��n�rF��"gT��nw,�pKԝqu�SM1Ƭ+�ۉ�
���:���= �u#��<f��zA*�za�X��Np���:�<8�	���\��>�������/.;��.��<gg\V�}��� �{`�r���w^���4��;P��7���}PW�lDJ}��ƥ�p^����MJr7��g_����9�f��~^~��w�<�8�\��TŘ�_q;�e0ǓVE��\G�Wj{�:5B�/9��[>�s��w��|.�D?t�#z&W�ʇS�F���r8:�r�N�����:���wJr;'��l���y����3��<���`V�'I��NG`S<�.�����q~��=P+�>�Ǩ�z�D����M�ɾ�^�v��
��k3h�;�L�RATg@�y/�HL�Nv-�8;B"\�]�o1X�<>wS�!�b���`_�q��P�1ү�y���:I�g@�R$T�ʽ�ЯDމ��^�Al�����y��Wu����ޡ�_��@ٯz�C�F5>5�o d`�����C�������ru�1�W�*)�-� �#�;�F�{��ۊ�&�}U=.h��G��}[��+�{AS���8$T٧χ,w8�m�nfS̫=�z�|�[J��U�����n�n�=�:��r>��>��{!J�F��87t�#2� �NNS�^���	�֦0Ƴ��bq��J�%af����\��v�(����Qëzv��M����<H�/j|���D	���f��'���ǧ�{�A���^ @�쩭�ap���}�H�F�T��%)�@��+�/N�����W�m��'��80����H����S���>�k�76����mL�Ս���C+�a�/�7|�u�c���!V���뭿c�>�G��}f��O@��3Q�� .��9�Pr�s�up�]>���PG�`�PϡLg��~�W<����K��\<�Sq�<����<-_g�;_EH�vG����ҕo��>H�����q�UӦ=������q��v{��]~����k!�e���J��NHQ��e9�q^������a|j//m�*�xO����䗡c�c���`F���A�U��>H�M��u3��zn:�J���3�$=�P��+|b��e��UZV�z���Z|�����K��ʼ�|kg��r9M�a`*���k�Ś��h]���*���`w�mu�+#������b��{t��ωJ�2Ǩ����#S��oDZ�Q���d��x{5L{���f\KKL<|��S�,��˾�Iu���0.�u��F3d�ռ�o��Uu8mvd3�?�t�yS��mYC
Cx��δ]�_*V�#���&���ѩ��r��3|�0ܝ1+(^��]A6�npj��󜳜0>��·�������}]�z"����9�F-�ˮ>��*��r5�Lz;oڌ*�:Z�Ee�U��g�Ǫ��B�������3��<���[�β�~�o�Y�Q%����sy٨�ybr'� W�7���T����ꉨ������9��3���H����}���� �ǵǫ�!k���'ݒ �5'@���t�o�(�>^츫�[���.}�i�}#Ƞ���V��b~��pon�b�*�5��O�Âu2����@��B��K6�?}=�� ����;+ᆟ'�w�[�u��l����r����"�UK7�!���M������Z�r�e��<���S�''���į�ܨ�m�����qW󩮣jd��M�{]G�:0}0=�������W��Mx�[�D ��Pԥ�����gz���=p+�޾�p�����9e<�;��q�H�zm����6��j[�|=�6����:���/�����p%�Q���D�h��nȜ�W�fk���l��l����W�^��\?j�/��#ȿ)���d	Y���#�*��t�9��j~�{������5��_���hʀ�K����4��r�ܒ�F�)����2<����=��ǒ�ģ�����VY��,�u]��&i�V�Sr� ��x���``�\�¯y�N��Mn-�Գ?�L�-'����x�kåX<�~�u�f���(U�P�>d���B���S�.w�[6���{:��o��c��L��O�L�
�d�wS�8%��#%���c'Ox]�էvi���|6=ig��<�Y�������{�3��Zw�p��a߄�,O��j U���~����<�OK�Sc�ց
�w�y�wt����w�)�3��"���ݯ��go7�!��"n}�z2���Օ\n����eP�9|�.鬈�W^���8k�R���YQ��ں��� m^^F�L�t�I^4e�+�<����ߞ�0�z�_�r}���>�����쩉)}n��||k*|��dܞ�����&t	�U�*e��=)�fY���a��/OF��S�&�^ugGV�3�m��g�y�	e�=�3�L(�wH�w�8>W	���hϼH���E]��u��y\�1��s���O�/w\���f�z��� 'Pd�[ Q�\��p�y��wc7�%z����α}��c�/���>y^���,�i��^�P��Ob���.���d]V�sK��5� �����v܈v[�z��.�Oʽ>xi^�9�u��n�V5���2��#�2��r���6��b��r��O���\��>/�RV�e�:�v�Y'$�e��.���C
v�Z8�L�/�y��������p��_*���q��S��)����O����f��->vǏu"{ç��}�X�=��M����ڎ&R�qX�b�q���M��2o�H���x����wj�:{�`����w���G����Pt�Nj��oPx�p8���${�������{��f�w�P��e�|M���97l�m۫� +�j�[t0��N�:��<��������W��⫨{m��u�u��M��o��n<5�<g��4����롗��6/zA*4�Y�����p�G���')�Z�u�9�t$�����{�&�}�wI����<�&�a��UQ*���$hqs׌f�G�OWO�Q½�\5U;�}	�.�r��;�a���y��	�]��Ԟ�F�F�y�a��_�擔-tDH{�Cg�|cΫ��9�H/B�:":��6F/��;>�=Ĕ�$T�mҪT*ʁ� {5�g�:�l�u���[������۬��d�Ίn�x�}/�Z;�iD��&t;��SNC5&��au3@�(�>�q�}.��(�̱>z;n^,V�1�ά���BX�>2�v)Z離���5;(�^La���-&cS�38��7�G[��w\tMA]�.�FZ���UN��R*�t�J{%I%訷,Ѽ3���z�6��V�w��֠A�+�]�v'�l=ͯ���?���z:�;-M^�]+3�$_��y$�C*�����ݙJO7zz�Ύk�'��*����~Q�({�C���W�˩F�$��:�<�q�2�
��K��l�ʏ�S;���(�]�{����uD{�����;�}R*5N�^Mo����yyi�߹B^#ŵ�Oq�o�\QmZ���ﻪ3M���#n+�؛G����5ݚ��Pց�非� 3�3�@�)��0�P�!>�ϏO��9��E_���k�F~���w/?U�R����?��h�r���~Zr������EC�M_���z-z��Ղ�[}�K>��_���8��׈��ב�\��5��yo��gl�k��g��OJ����<�ͺ��d�������7�E�O@�bb�!�)w���1ʠNق���1z�b��T�e�y웽����^�c1߂���y�:��x��\V�xZ�Ό����]��)�q���=���g��fc,��.��WN��/ac��q���V��#�hm���}Iӏ�:޿�d�"`鋵�T�s��,����i!%�P�J�-&��@��0\�gU���Yܸ�U�����=����4�ͺ����>9�u�}Bq�e����D��O�恻2�HԾ�BdV;��7��fꦶJh����3e�i�I�"��R}X2�Zӥ+�j޼V�=��m�B�������7�dKN�|���E.
�^	�\���M*̇�����)r�F�(���u
��u��*iۜ2J�Z0֡��*��*FFt�{V�!чa���v��07G�[:B��Wk��1�,ut�6.��y���5�3�g!�r��W�x��!v_^�V��t�;���3�s���9�a���YM��[�{�}d�2�v��:�[Z�X��M��2��Os�������*�kX�/o���oN��݃v������[P��fm0e��qU��g ���j��+>B��꙲|����Rv��^�jX
�J�}�EB��Ţ��Ȯ�Hsz��>����4�0�%�yٵ�{��ݎo.��TŠ��5��
�NF^�짖��P����c�UrasI�|.���<��66���S̠Ʋ̳5�M�;[5�W�����ʇ����V��+��93
��Y;�#����b��wJki�8q���~��>�7O���<h�]���d��8-5��ެ�Uٖ�'ӯ8wMδy]���U	��@�*o=� k��P�zT�72�E��'��~����̭��x�v7�dSWhը	�/"Z�yK�qi.��8�p#i���=Ct@�!� |.��X.V
4���YΥ���f��r;}�	����Cn2BZS�M�.�m%��gd�݆�7���W1HЎ����E����&^f��Z�.���L�I�[�jr��՚��'�1d����f�r�t.3�c�
I;-�c����!>�y ��Nc7u�Q��p�r���sc�jF@�3�����Vk���#h����Dg.��L��'k����u�an[YZ���rn�H0�/w�n��޴�Y�A��ق*�fj�n�o��E��A�J&o��n�v�[Իl9�'�k
���7�y�g+�]��	(�NT$�J��,YYh���g� �;0+���'�Q)�g���td�d�@@��ͨj`��d{�T-��)Y|/8�rj��q���kb��!l���k�m�����^��ڕWL*Ֆq�&P��]���\x���>W��I��bǙ{R��L^.>5�hc��u����:�ح�닆Lz�sE�����a>��Bk�:P7W%N���Y����tm��s�0
KF���BƊ�ܘ�Qy`X�n�)�Ƕ�<r#�<�}y����rJܻ��n�WkJC�kȨE�tY�����FR��#,։����wf����p�i�;%��See=(��x�p�ptﲇ:�y���n�cNБV%Ǥ!%��;���sq ]'e̚
1S{y�\�C�;RgdX4.U�h#�q�حc��L��>���C2!)$D#"�c�ddă$L�#A$l(���)�d#&h��e6fF$�"#D!!	1B`0h!0a�I��)9��B����%d�0������1�`�`�I#�hH�"A4�f�D�J�R� �D�&CF#a0ɚ$ƌȌ�Y,�!79r4���D$�%�� '�i��6D&�%�@R(�",�8�0�3%*1!$
BI$��!`" �h&��&�2JL`�4113I"`�����e�D�(�4�h��C$f@�4a,h�a��#	�!!� (ؠ���4�S!#�Xm���e��h=�о��X��W�;RZ�I`���2Nk7Ԇ� �o0�F�I�y��s�ܫ$x6���\�},V���mo|�@��]ק����
��A��kR��&����Uu��Ƥ�e���o��%�-!�.����N�����?�3��o�l�e�េ��M,4;�a3�$^��5&S V��d.���u�ŞJ���.�>�����NCۓf�L���
⧨��G)߰�9�T(#W���X3-ßW@�]{����_�~���u��_���Q	εV ����	�S=���>����)�����a�*<�_	}��ayl{�W�w���N/���jR�̧���U_l�f�p�K+�S;�谺���a�4�_���{�z#:���u��\�Pq�2��Y��T���!�$�AD��:`獩���c�� =����t�s�����Q���;���u�W��]���
}%ې�:����JF��\|��qW-�	ϸ�3���6�lxt�+ү�W��o���v�dd��/���)�2���`/��������މ��V���Yvyَ��_�'c��'/��2/�UR͢T$�}��x��`�U4\H��U��Q��*
�ʝ��eJ���F"!��mI�Σ�镔�W�(N���K�F5Z,����Q(��/6r���j5�e>�W��+e�=���n·3�f����*��n�Og	4IY��[IF�������s��9yC �9��.q�����ћ�C���1�=��A��&����y���3�l�1�B'�~k+��߇b)R���qd��JKU�	o]��q=�<w���O�p*z��%#�EP����]�먩�Xl�g����sTS���}��i�GQt"��ǜ����g����#�^'!�����k}����~�ǐ�e��z}z��<���ъ�L�y�	���י>���wC/�t2f�] Q1����W]\2�^��7�0���W�l���/6qo`�{��f3N��v�p�����k�q��􃓗?��8=o��qJ�X�������{+�m���o�r��'׼|�k�Y�{�/;�t�n�dsQ>ð�{��
���c���'V�v}Eܞ<��E®]�u\ξ���ӡ�=�G�Y�*lz�\�dN��Mt<gjҪ�u�Q��t}�.��S�]hFZ�1{zuq�o#izґ�����	<jO#Pfc�=�B���[U������>��R��#�{ٞ���'��b�U��t0���Z�֋��yY�8�j��dB�۵��K.����S.��tY.��Қ��2e�����E�g_q��7��m���Ef9d�z-�M�T2�V[���uu���7�9���R���TF�wY�<]<M��I�A.~𾕗�i���r�%T΁1�C���a	�,���Ҩ^��f;���ǳ�:��~>�u���X�t�9pڸ{�k8��τ�l��|g@�
P09��%q��6�������z�� r{*cã�u�s��;~���f�z��Âucd�ET��eG���쫎Ֆ��z��]
�c�e�h}\3�s	�w\3�0}�������8c͞�Z�.Җf�
}u�-��a�ͲO� �_�M�u`=��I��_%\*����Nm����u}rz̓�n	BR���Әa�՚*�����z uG�VD������9��3sۆ�1�8>īT�$�f,	�^�AOx�4,��3<�Wv�"�-���#v���v&����4^97�8�hg�3��q��O�F�'qAo��a~6�o��+q]�^qHf�3��1����N�qpo��C.7�a������le`wS�pq����mˌ��W��ug�����WT����vyG�?J�6���,5�y�&^z`�=�hx��춪�?��s�:Z�I�	^��5�8]��5j�;Y@�F�t�T�A�ҝ$�����q���]EuntΘ�Ul�\z�B���5Ӭc�k���	�]�7��!c[ݕ�����58��9[>�����ڮ�x����*��&`���x��V�|�7�C�~O�]K�࿷�������]�ӊ�t�·~J�5|^��;a�\I��0�k�8�Ϗ���N�e Ǘ+�SԸ�|�kS�޵���<�z��,�yU��]lx�=n|JL��;0��FD���x�_F@Tj�\j�(h�V0���Պ�+efyƳ���7}��g9��B*�e�_	����S�9�Bɮ)<ܽ=�y���콏*���Z�<z�q�:㮣����]+3�ԐP1�"��R�����=�ynB�p�5�k��jh<]\,,��c=���w�sX!���o�t��ȃ#��[|$wKB��F�x�<��M�L�����([�׃����u{����ۙ�z8��>^�
��:`A~2(D���gx�Ȏ���Ag�ݯ@w<�/��3Mǻ����3�!�Gj��M�o0�r�Oj���D ��0��*�C%3��0��ه���}��y����ظz`꼙��Y���g��fк�񞙙,b�-M� l��_T�<3��54T=�w�V�pƘ*���DQn�� M�y�<�Y�³gz�h�%�v.&䕮���"�Eĥ��n-��acr����h$�9>Xs�u*�&�[����a�c��؇Jw-����a<���LÖ�[���w/����6�{�(�@�1�lD3���Þ�����ܩ>�l����_��8�;����k�o�2CW�ڰY�4$m�U�,]wy��{����Ty.��j�_ɾ�/�zs�Yz��#��;fRw�s޸ /�c��}�N�E)xk^�U�
�:GT�t.��7�P]*ix]�<�I�3J��N7×�n�E��>�1l\/�ӡB���_ݞQ��Tt���hn�Ų��;ۓ�S�!�3Ǥ.�Ԡ�B��r=�&��<�f��]e��g�u9����	y3ne{aV�ў��&�=�w7�Z6�D2�=�<n9������O׽�s3�+^^�n�d��eמ��b��/ޑ�|�� �K�9�6n�ȩ�NF�S�n)tǶm��2o�h�%�w�ĭ��q���Q�ָ���`�:��z�~ۥ��d�Q����8E~f������j#��Z�z�{�r�r���=B!=�W�X��ayl{�X�\>yt/�:I�LL��{��M@�`��G��V����qE���wA��=����g3�/�����u����N��=OܭN���s����i�E���6L�X"w�ӕq��%����Wq0��f����P���-^=6o Yd�Yn�݃�ڎ�CtV���J��GJ4ǝ�]Vl�Fr�p��p�:]���,WqJZkd���V.*YWn/F���ˆI�ˑ�FR7S,..��%}�q�=�ïP,OG�`^���;�>���̴�Ϥ�Ðs_I�$)�1�# �\U��)�-�L+B��xfv_f*�b��y���÷}de�U�p�|'��{2��|��03V�@5�_m�>��J8{�����{\�=����u��Y@���
�g�M����ݾ~�^��΀a�F�,����+<|z|���P��?PU�)^GI1��f�k�=&_Y�\J��"�W}חN��E<����ԵYIo]��<�t�ކn<�m�d�e�̹��G���Wu�G��%�S�^���}W�����a�5E<�W�|����͸NR�.<���!]�2�W�פ��il<���!�᱅��ɔkʧ~&T���Rw��yu}�w��\�W�Ԣ�<��j�� �@�adWW����+��c �����ǧ�rz��=4�/���d1��[�Ǳ/B�G�����􃓄� dਓ����_#����1>%+��u�,U��j�82����c�ـ��ۍ>��3�0�s���뭌v��y������s��þ>=\�G
��>Ne�����<�vz����=�;���t��f�]��v�yAὣ8��֕�{�;���Fg�x��](
�ۆ5R�`�yg�{ex�畲6��ɻ�#��i�A��[c���Ȗe�E��S~�v���z�Wk��>�	.�B��{t�8�̭����:�"�B���3�f�ʇtꑖ@�� +�NWt��S�ֆ�N+$v�=��#=�������](��N�'����Q�FC���{U��OP�!��Ģ���ϧ�r}нy�{=�%Ho�^ZUmEJ' ߇*�qS)L\EWRg��L�O��Lw���3|=�1e�m�#�a�����Q�����τ�mIѝ@�@<�����lcQy�}��[>�^�v��Q�Lxw˳���G�(�+���\c��}S��p@N��{:���㦫��n˯v� x湮�xm,��B�hx�u���[�߻����q6�jx�}'�禩��͎3�W|$	-P�=����՛d1��;c�{ռ{ t��o����3��}�@����q/[p'�;�=T��N�La���G�ݱ;�m�v���>�@�!ɞ[���vLffl�rc��tYnৎx�����/a2��:��K���Ob��d˧Gڅe08p���>�:�Q��gu*�d�����6��[D���䳒1�9��*��M��&�VEF�h�ʯ1�Xr�`�X ��g5��VZ��z�Y[�`j�@�Cn~j�$}�|u@׵�5��3+����P�Ov��4j������c7�ؽ�]�s
d��}�����ޡ�*W�R��
4��K����Ղ���>����rxc�ș�8�r>}N�=�U"(u�.F�����롗�C���o�X���և���z�ջ����(��Y=�d�Z����C5{��ǔ��\g������&^z`�p3H��zfvd�Wf]����Rq��'0�]z�7Np����QyY]j]W������Y/��+����T7��Q�aݧ2��N��P]���_�ax��ng�B�uFS O�+��eqg�-����W��1��w���>���/ە��|գ�Y.��e�6��Vf8G����,@n�(��������mH�=��ɘ�qS���g��s�(/��QD�~:�L�r�VB�p�t����잇��(�au�ˬ��>}=�z#�\v��y}/q�� ��<(�w���zǪ�mW�e�,+�<��/��Q���p�=ѝA���q���b0���T�p�$�H��z�� ������I��8D��Jw��)Kn]�!d�Y��fCS6�呛r�s�]��]���
�f�Q��gm��1���ʔ��ԭSy��xA{��f>�έI��G����yW�N6Y�>���u�'c�^
2L�կ�d0�n�
zA��$�z�x.v�ç׃���;�#�W� ���z���ß�Md]�I�3�E����f_ � yD }=Ƃ�f���myA~�Gs���8�;�uJXn�=S��NCq���3�+nД�g�a�sRF���@�/��M,ݸe�6N7xH��r��M%��/W�xx��i��ˊ�3:��Ū�Ԁ��B�*^��ۤ��5�W���J����vFH�n�g���'��O�/�k�>��CUu�L�Ս���Az/1%s�ޞ���o2V=��6W���_�F:�v�")7�x����3��5��,��稥3�c�K<�}�&����jk�$xM���ì����R޼uT�C�l�1�7�|�HǞ^�ީTbpL���	�=T�d�EH��M�2vm�G�}�EŵK��o�i}�Q�?*���$���3�߯'2ns%u(��B��q�"�5�%T�ѿ�ZI�Y�zɳVw�
���jK�tѮ�)o����V��<�C���K�9~�q�w��m���6n��ś�&���,��o�~��?mx>�84@[x�[�̥�+qY4��g8�R������X0��O�z��w��I����;��O+y��b^��G(uf��i}u]ˬf����sٸ��D�F�'�����M tX���2Ք�Z�b����=��������WW�����6_�c��8��C1�U�пK�9uɳt&xz�J��pV�ho8U��Y����=�'s��ڮ����[⺮�3c����HвR�����&8z��o�����VMq�r8���C������?B�<׼u�-�c�W�w����2�����u[����s������F���a��=����g=�×����+�,qK8��^^!��g�\ẹ�"�*�3`�P�<*�b_������vM��7"xoe��]�w=�<+rtgD:����l�K� �N�0�4:{����89��V����9,�c���7��������Rp��{��ˊ�_�O��pB.�d�����
ʩt�U&��ӝA-����f� ��l����i|w	Q����|d[��e@�� lA�!'*�$�Lׇ�Ս�����x	f�a>���Vx�6�؎���u5¾�μ��;`��#��<K�VѺ/rj�a���ZN�Wɺ�\>~=�}�����km����km�����m�붵�m����m���ֵ��mk[o��k[o󶵭m��Vֵ����ֵ���[Z���U��m�m�k[nm�k[o{mkZ��[Z���յ�m�ҭ�km�*�ֶ�歭km�͵�km�mkZ���d�Md��c�	�~�Ad����v@�������^��P@  I*�*TA@�P)@(R�*�P*�@Bx 8�DU@	T�B�"@�P�QIBDD
J���U)*�(�%AL����$�T
�U J(HTB��J��(���P
���T
T� q��)��f��0���ZPhT�dJTkk@ �@����AN�J���B��DZĸwV      �   Հ   n�   �+�.HtJES3%R�� �UŪ@�Rl�i�R��b5H�#�I`�I�����KU��Z�AB4�*���1�b�6խZ�Um�I�ZյQ�j֓aUZ��dF��klST���5����Y��b����*AfȐ"n �ꩫQj�MR���m,���cm�-�aZ%6ʄڰ�F�f�SU��V�hkfh�kR�ZƥTdR�7 �SQm��Kc�*�P��)�E��@��*Ea��-jlf���+J���kI*����P�-�ݶգM�m�U�6��KM�5[f�Ca-Q�dtj��5 ����I-jV�]��RJ���hTA� 6�jٶU�aV�I��35JԵ*�Z`�A�
�m��d�SL�R�T�(�����b�T� qs&��f���H�m�l�f�[6j�CMSL��h�B� ��H*n ;�Ɓ�ZRѤ)UTCj2�j���,�"�Z��6���5���R�@ � S��ҩR* ��� LF@�{C
R�Th#C 0�4 L$@�	��ij1���3 ڐ�~%I � � �  sLL�4a0LM0	�C`F&� �j6�4  @�}������k}�v~߻���nw�����2��{�!!���0�9I���Id$���t�$"�a��V���b�Xl�����e~/������
���QQ#	"QeDj�D$#eD^*���
��eH��e��1�`S��n�O��I�8$�%�K�{����J0r�]���6gN�R�+e�cAEA"����}Z�Ե��s�c�UgD����"��[F�f�L�P�E�n�p)p��:;�f�tGpi��w���Kc^�u[��iԞ�?�Z��o��&�׶��R�
����X
+v�:�S(4liV�Ej���;�����B�kq�tJ�h2%ɳXDY�z>��XR�4fn��Z���2TU��Pwz��A ,�Y�����q�cU1m����Uѽ_%�V���t!�y�A= R��������*­� �$�ժ�����Wc�X�o�ŵ����cv��p�ye6_�s���JY{țWu�:�*���@IyY&^*V�H��N�(e�$r��)�zv���}a'%���`��m���^Z���*}�8��ެۥڝ+:q�M�h3��w
C%F���۲������ѭ468S�:p	W6<��H�H�Ʋ�lѡ[���wJ�)�2��V\����l��U��,� ��bͦC֙�7ZM]�ӗ�)�h�R�{r��su:q�7t����Ł�7�x
�l2��Ӏ���okhb����qԌ�d��e+W2��$����b9�օhY���B�f�C(9&�k cl�A�sUf�̫�6Xs.�)�-����9OM�+6���f@�H���j��
��v��2�H�tp.dcZ�/S%�W��Sg�EJ��n��Ǆ�368���g]�6*ɧ�$O�X���6����� j�	�3\"dg5�Z$� � �jܻ���2чTʽ���=�v֓^���I�T�YR����2�[����B�-�Ǝnn-�s-6�����0�K��C4^fI��w�iћ[� P�9g[0¡q롏-V���k�-��.��	vnSŢ�wF���r�d��u@�M����m;;-�fÊ����(̭�D��4r��c%��&���@;�[�5H�=F�j�9���3y,�t��.�0f�I%B�.������1!w��N�˗����̗�L8#���7��G �̽M�*�`�`���Ɖx3KWK��z�Zj�����*�&Z�Kd�BY� 7ik���7C.��U����v]�a�v�R{4VԶГoV(-<��ܴ�����یl��@�MKu��Kwu<�sQ$��D=��vV����b9$�+P�v��IMiY�Ȗ�A�^R� KJyTȬ�fn./F�A�J��A�X���RB/r�[ۚ!H]�@僧
�!�X�ݭPe=.��$�F�U#�I�X+E;.H�ѫ/Yv��FU�qSYJh���hRҬ��"�vr�����]oP֎��9A���.��D��T��hQ����/���QT۵a�@��pKLcgi��J�v�;�5�,���N���hv:�����MZvz�b��\Zz��4E�$V`�2�ռ���V�q(��[m!��A���&�R�F�2�u��X1�G;�}�|���$R���F�)�-j�U���oP0�L�5sF$���@��ܠhW���81̦H��x��UԐ��'-�Eɖ��mV7nP��/p�u��R��_ΫY����X��ln�����.���ݺ9��Ҵ��v񃁷�X"���xj�2	�Dj��ֳ�t��bU��"Q��vaڱY�j�R�(^n�11px�%�S����B�"�K�ImM�ܱh^"��� �bXrA�g-�v�OZQսu��|���D�n��4�IR<wZt,-̵��e�L�Q�Tv��@����dDu�ֵ�[��hF볟-���ʰ霥�����X��[�����[d�:�,^_���ˬ\ PM� ���2�u�3�X��Z�c6�|v����k)jƕ��72��d¡v��c�i�R���p�M���T�[[��� օVɚ���]i,d��)��E+���g�̛#<iS�i*�F
X�VhD��&��N��f�kV�u4y���К���o�;�Rj%*v�P%�ko��m�2�T�[�����j7�meX���۶��7t
�Ӈ5�Y�b�i�@GR���e�`���ݽ�����U��Q*�Ę/*,՘5*֥�r����[%����ͺ���~t���X��`rYg�,�Ȍ)m#���"��5�Ue���s�t�Y��j9�s>%P�+[r�B�FI����[Bѻ��Saٔ��������V�ݽ�Ctݴ����4��13kr����������Q"�JRӶJn��m���v~�K���j�ѹ�3ED�5�I�����]�P���:77%ڀ��t+[z�H�2���Mз��J]6=ղ;ir&t�d�n�A�cՅ�ӛ��,ߘ����6�n9Pҥu#��	���m-�Z^
� V��;:�p��Yx�;�3���&�.$/�Chl�l]���bjm��V�I>y�Ыk6Kk.�[t����+��b���;W���	��>��&������{��J���5x���6K��ei�VҠr�*�%&��j�(e�^媕
���4����G(1���fC7]������L�a']��7-�����Z�7������6٧*�X4E�����Ȑz��+���J�)1e���D�Xv�_PF�fh!\A���Un��*�H�pڑ�V-���"J����2^@���/!���wnW�M�Г4��r��n��TfnVX8u��fF��N�Uu%^;o!ͲN�
�U蔳YNKK�l��dʳo)T���
C+^�-���z��-s-�3���W���ts��ux���j�1��8��]
�LfO����Ůn=�E�"��1��ְ�$V�JЦ%k#V�y{Xnj��̙5Rǋ/dYV\5;]�鬛n�[��7��%�H!��*��Mn����,������
ׄ�3�R0ۭ�hg�f�pTF��]x��J�ýB#K+ c)���p+� �EYp��h��֣��0!l�1��ђ����*�*Z�Ylfu^r��
w�7h��������+{���p�m���Cm�wCv=[�B�i&ܺ�_�XSI���	5d�J{�qo�u(��U��(e�q�jZe��m)��[5I�Gm�B`e��ln���umU��X��֪\��+��$Σ�%�]�Lz��%���zU4�b�-Do$���(�����-o�05�"i�.�ef�U�+�Bo �3-nm�5�d�Jށ�[D��� e��)y�F��%J�c�Z����u�I�\��03Y@�ڃ]Ӷ)P;vq䣱������5V���I.�!��iv���'/��h�y��m�	��0��.T�GQ1<d#�K�Yˢ%��H������b�4w(�\�X8h]��@���G-�K�Zw(��`lRY�����7��ᨦUX��%o�5�SX�X61�W-����	���n�Y�l�e���ŏ�i�7�6�l��V�ǖkR�J�4�P@�����*��c�ÙW�������[��(�#1���Q�:bL怩�R�vt訔w��V�Ƿ�V+f����m��e&���y�J�K�Z��ս+N��L�ݑI��ٹ�͇�-.\�5�z���ke1�y�kS͵��@��p��Cs&ʊ+�U�1^%{1&I�nJMg1j��]�[�p�����h�\nνu�U �hb|�un[��U-3���ӷ �L�]�J���*e�.���K����H#!*��;Hi�Y�l��u%��`e�l@�u��6�="��Z��C�8pa�M$wh��+I��Ixq
����F���̍�ܨ���+N�vT�kY���^�ʵ� �w0��2T�e�2����)03j�U����h�C{�pl���ol�t�i��Gi�v*U�yJ�,L���m�ƪ�+QUu�]�ʱ���;����B�@]ʚK���f+�I�ՙY%b���/�vW
���;`�$m)w hQ��V�|n��0��a��MaI���k��6��%+d;��.�.������D�I�j5{J����;5yv�V�ƭ�h=ӹ�-��{X�w���	+*��^�jZƾF���:�潩j�Y�z�7b��w��L���)������*jՎ���gCU��5�f�+��As�j dI�j���q�ʽ�hˏ1n7x�n��hi4�b�(h�+^˗�X��{�3%X�N����M�,j��[V�4�)5ui ���i�7J��)��f��ĳF�׷f��h�%��G���r��u�KW$H�y[�h[�����l�WQ[�0ե��[D�G,VP�m��tEN��X�U���8[m�$����caHd�p�o:��dhm[���`]U[ZҒ�+w�%\�0�8��Aȍ
JR6tۍɷZ�
�o0��
��7h[���X������{@V��5����W�B��J��o�,�F�I�G��Ӷ�S���a�]W���⒥�U����u�(S;Z8oσ�M2��z=�W��                                                                                                                 �                                     7��$>��V#I{��ucΣ� R@�t�����-r�����|o���J\Z�Q;��<�m<۷�NΗ1�O/WR� 
j�mZ�{��U�]:Zڮ�ԥ����{��5�R�;��G뎷0fȳ�]
�%鸇eJ�^K�q�6�뮥����@[V��z��NȬ�����rq�7ڰ�>W1Y�t7�\�4��鲠mM�X�ū�����r-���VuZ��X��q��.+VU�k lF�k$��9��;��I�A����U�*��R�-���J�7��fZ2q�s��k�K]�:#����.��ۇ_$�Aa�����2
ޡ��R6�{xtdYy����^���g��Z�30����:N�l��k�ЎӜ��d���(��蚷��q@_C��zFv�Mj�t6�׌�L1�HeӮ�r�(��Nē�=5in#B��iǞ�]�{���bj�AN
�[�7Y�_Z7\��ި�sV��nC��tm]uc۶�}������er����kgk!��¼�]���u���)�jf��;�)�����T���2�閵�g�'��-���,�y����׽5$�H$���]ұK��l*J�M4s��r0��G<��}��qC�^��V�g�X����ȫ��U�56t��)gWXi�`�����V����K���^�wh�Lш�qQ���ǈ1�$�> ��Z�y����JGS�4 ���z�5A1
҆�ݦ�-��D�
ܠR�͐�*ڙb� ��Wςv�^^NV���ҹ:��M�<��\�����i���םEń2yv3����u#iln��M���i\��1nupņ�V��)Sqe�vX ��{��?�� �ר5de)g:�U�Y��_:N-���.Y����*��*���S(gpڰl�����:��-ˠ�P������Zѩ�2��:>�k"�{�<q)-���M�7��zb�L��X�lgF�U��Z��'�Gtv�Qӄ�瀹\:6bì�]��u�A�3�g�@B�7�Z�e�.Si�t���:r�d�kf%��j�Y��* xR˝y(Eg�
���v,�.�!�G�㦱ǷL4�~s�й��]�qr�
g/��>��tkvAN��б�|��F�Jؗ4;CE�u��'���b�VeFh ����*'��#U���Էʥ�صŨO��Uo.yu����3�LˤgY�'g�V����"�y�wMdмG�j�MÕ3a�-����j3aئ�>X����$��e���X��ì�\�N�.��ˬ;\B��]%Iӗݜ�KT�hGq�>0ը"�̡wGF�����VgT��� c�V%��hItlH�SW�;�v���H�40	}XOa�B��J�14R�I��l� 8�$�7Æe�,R�l�[x�d��d|�âHO*έ̖p! *��6 t�fJ����M9+.�d��Wf���!�8+E��6�Yf�Hp�Yʹ֝��s�$[��P�:HB�*k��9y�~{�:床�ת5���H�N1�^Wc
nj��*Ŋ5"b)��	��.&���@,"
�/,ӂ��ɷ9e�(����e����wl�เH6�^�&'p+���%t+�꬛Et�E�ʗm�ҳ�%��.�l_UB��T2�Hr�X��_g[M7��h�槙�����c�YM�K�Z��y(��d�(�����y��::F���v�c�#���R��z�Ѱ��ܭ.�weTqu���/�u캅H��L!L]��^��V́I�ɴ�,��08nZ�:�9K%��eiٹR4"��fF���4�W�﷘�\8��c<�j���V5��%w�E�ݼQȃg.�<�2�X �P�-j�o�m(cńsʷu�u:��ј,Muʂ�%�D+pg*Y� �fX2]�����
MN��Z6�##�𚇌YY�jz
o^[n7��â�n^-s%	����9u�|up�e��PǠ.U5R��u���[�ۛ�6F;έ|�/��A��Y�*�k�� �l����α�Ǝ)��Ʌ�ij�"�)�L��0���t�X��36UԽ��B�0Z�l�SԲ.�na/��U��d4;�^vyYW�ھ��-�}�#�RIM]�kF𳱩��>Ψ��8���5PTb:;�
�uk����L`^��m�1�<�wnML&��r�\��l���Wdw'''���[\&I׃��.��V�@��N��-��E�l�܆R���@��<A`����ֽ�V��je���V��Y�e�pi����q�3�����zŢ��]t��t)��6��N��^l�X�Ն
�="ԯc�c�s�ujٶ�T�\6r<v��ͺ�����mJ#^�=�6tf6���4w6=��%��"����w�:�n7�8�\���;�b�P7fk��5���n����v"7�K�j�&JD��]J�(�k]g�vV��v'H��"̜b�C�9Kd��/���u2`��=���j�v����Bt
6�w[���`�K���Ŧ�賅�v�c@�F�P'��%�:�����J�x�'��]� z�IHe"�;��=�ڽd�÷���Z�s�Z���R`����Y�_u��۴���R$����s�[�J�-M�V`6��+k7]q8^\;}���0�c��u0�pýv+M�j2-�\:f2̾Mu�ʏ�D��J��f�s:��j�J�b�:��ӡb@Λא�;��.���{[Isu�͞��{�h4A��v�Cp� �,N��/&X������X�[]9��H��ʇ�ZZql�K����δ���.p����iz���]2���9F�%�+�ʳ�M���)�ϻUm�Ԥ�Tz�*o/��ͭ����r�R�I��[�s��U���L����;���J'��ˇz�dp/�
t�	���b��IW`_;g ˆk�j�廥3ɚ��<'��iS׸�+��d᝖ѐ��*�B�9��L��n� G[�i+vm��ֳ1�	͚�U!Uy՗m��\��nE)��r�Yҭ�h�h�Z�يG�Uh��C]�����Q?��jvX��췠V��VQ����d�c'w�a<�b�5�7�(�CX���m�yͬ�ث6��qnFD�q%@
�;/Vfa�r��#�}ˏ�	3u�tY������ėXU��;9�K�v۶�"�\������;{�#y�Pȇ�JY\'�{�1Y����4r�SG$�F�u�.ıΎ�:��MS���,1E�8��f����&�ڵCE��ke��/�y��CF�\鄻���o!g{��mdNY�/�v���3v���9.WH��l���/��j����z�p;8	����;�k�ᒻ��:�_jr��}�ˤZ%��Mb�㆜���a���".����޸�և�r��3A����oW.���bj"���EdSuu]l9��N]ғ1��-J��6����-6S#�rͥ ړl�s-�4±gQ�e�:e
6bZ��QJk*r���;��r̬�{���Q|�p�+�Ƶ�K�ou�ՙ��q�9� �9,�;ҙ�l��Y��q[ �2��\��@�uP����T�g�����z-L�c:I7F��5�4�Y�V��U2���iެ9�a���7�[z����7�n���N��V-�ix��_9i62d^]�C�7P�ˈ�͈�WM�A����C$�Wp*��������:հ�_���6�3M"*�u�;�.͒����3��m�V�����"ΊK�ʁ_V�C�rq�a�;lK��e�嘁un�,b�W��2:Z3{
f��9d���Wg'�g��]J�<�{ �{W{�{�� ���)���s�[.�6-�[�D�d��`��R�DT{6OP�hmk� ��u��DRŹ��"l8M���M��˾�	��6j�2��t�n��«02���s.㗕���G9,	�Y���j�[�}��	�x�&����(-���~Ԟ6��o�M'7/a��*^jU|�k�j"��E
�zVU��D�纯AZ*W!㚺�ϖ]vR�O�5C ����zmۼ=�໵\���>\q[yR\�[�1r�����|�������)k]��b�Y�����nf��n<�S|�ր���b�ֱF�,n�����n�Lw)l�*Ծ��6cP(���c����,�iI�ԗ Nl�s��J�� �Bޡ�f�h��7"��ܤWN��Q�\Լ�ɘ���������7���N!Վ��(.n�cfv��:,W0�E�T�v����P�1�iN+3L�T�c"��d！                   � �   �iM�:I�:8�nyP �H@              s��9�s����_�~�'�O�������F?�BI!�)�ՌD��j�H�H׫j��܅�I!���8}�c���{͵�X����Y8�����Ib��������J��T�&
�Ƕ����B>����0��9�5�\�8EiT�Fb���d�z�,�vLxݬ�B2����8�9B�-8Gc.��,�z2��j�䌔'wU��a|��J"-i�z�8�*���S��ʹj�R���q]vd��%+ic52(W�u�������R��a�E�yE�Ѥr�5h�:��ki�5�c��mM^JV������*�̓`�: �wi�yK:j�]ֈ2w�y�bf7*�A �,-�C��9630�}`c7��xa�Fӻz��w%�������Ln]n2���xm�ḣ��AYƾǔ�[oJܔu�!�NL���{C9"���o����2JQ�S�H�^Jx3��p9�����b�|OZ����NU��ȴV��7"���H��^���|pel�[��x5��(:VRyGrAԬ��/�MvM*�12d��v>f�SŐX(Kpm$TN^]��~Â���(�����N0X�H�S�Y�ˬ�;F��	B��J�r�+f����|��#K����pWLv.�S�Xh陳jP�Y�u���R��Еi�L�Ҧ_lu��.��*ҥ�F+��5κ�j�8)��0d�˃En�[��D�|��{n�b\v�[c�9|tB"յ��� �W̙�v������a���Y�Ĕ��M��e�2m���E(�)��[Qm�Ysv
����L��eքT����6�5wBv$;`������s5 �j���u�z��-Q�n� iN�	z�=���ކ��	t�]K���a�D��H	�%�p�p�V
��]Wۇv�&�E01V��K� K.�䓔�㖬����F�v[9K�]�*��ʻ�wl�!!��Jʱ� ��&2���4�o {9���'��N�[�-J#a�&`�`���9�%��H�<�U�;^�|�1��FZ%N�?�N�3�;�:9j}v(��t�Wi���}�w>�4-�ٳax���&.�\9�i<S�h��RН�bk�ު���Yu�|���b]�
=W�3{Vv��ƱFۛ���%�9M*gHZ.�f��h�ج��೪݄��ݠEZ�jB��@F�s�2_���u5v���M���N.?��Yxy�dЖ
	k��nZ��	]�h�]��gVVl�/�b��w������]hZ:�S��4. ��yD�E[WcO�����X�݊|�d\*aȫ{2��i)X�/9R���S��ţg�D}�/�٬���%�ʺ�����M�d����[	�Hݙ*S�ݺ�m�&ىǹh���{�WwY!b�,V��g[5 Ǽ\V3UJɕ�]]6�[D�ú���������1�N]e+9#����+�Vq��`͡E�:i�@��ͫ�*���{)����p :,�I�{z�3E�.��D��2K�)��\xn��j���c�7�M�;��Kv����zU�q���Z)�li�\P<Vs�*�L<�7�쨠�~�&Y)I#ʔ�G²��芼�bn�A7ai��R$P#s����]�8��Y�e�`�d���
.;�7Y˶�=��42��^-�`�Dur��Ē�r�"�C4ݡZ����T�3r� �����۴�B����2��h�M�Δ4�pvJ̱��j��Y���-��o�*��FhoQ�ĩ���K�></nU�͡�Ѯ��7T��ؚ�q����;I����sP#}�Y�U��$J����gr4�R����ǽwN�Z�P���]��լ�L�q�-W-4��F<5r�Kw.wL�T&�b��k+����M5��8w\t�� �[\㧱��R4�{�Ei��e��B��SEX�]'[ٜt�Txn^�pG��Ò�Mc��� Z��6P� ����nMu���H�p��
F�g)\��
r�*N�K���Gn����n���ؾ�D�E�F��gM��YXxM7��p�d땬�"i���7�e�-���'�zs�d�F�s�;���9ff�s^d'���B#VP�˭�0�c/@n�m;�%�G[��Z+v�t�ssEZ���X�mZ��"r�H�G&�˅P�Yi������,�wi3��M���E2�nv�T^��n;��R�Z_�ݗR��S��#8cO��X����\Eo�3��[�k��SM%�X�b�v�6V�F�o03s,fN��WAI��֙�Fs��s�Zjʒ�뻏"$N�N�o�%i�8��;X�ɻ��X'{3���&��%Go3t[&b����t�H�ݕ� ��dJ�3DޡAf����Sy�U�2�Py��}]w)�9�a�(0�nQ���	���rT��`��z����(+�������ln�s���B�	x��5'�-������VYg.=-�B���çk���m��b�Z�J�De�f^�w��X��+�`R���,�,*���L�@I���t�r�P�G��S�0�@':c�<_�3r�6>{�ކ�i���r���f��3x�����S�WN:����.7t4�����,������#�P(�4��� +���Z�3M��@ �i�ّǅ���$�Zh��ڠ�%�6ږ���;R*T|�����BĹ(]�����|)�Mܩ��k�h��ݾv38Ϟ��)�]y�^���ƅ-;����cڻ�]X5+�TﶧDibl��O��c>��u���sz�P��Yˠ����NN��`�Ӓ��;y�5E����5,��SeEU�X�嵴�\f��d���X��ӦZ�f�t��i��U�|���\CC�u��XŜED�S��2��a�:��E�7+-$�AO���w�C���ݼ9Mb��V��	H��2��#���z�'LMrwC�1���ƍWN`��DuE�|ӭ�e��b������4$#��ꎲ���r�-�.|�f�[��Y8.&®jY�S�/S��D7 T�>pX�����Yǟp�-Z�v���I"E(,˲54b�Ϸ�qr���瓜�[պ0[r^��%���í�\���ja�au��Y���b\�k���j��S�QV�ͩsw\��Yn�{�-�	)��3e�>��՚2%�^d�d�Nf�C�%֧Ӻ9�z���pM*KLf�:�]vK5)�G,<��p:K�@�!Ö��bӫ��ʇ�T�M6]�vΣY�R=��I�����f`��2�)Yj��y]&���H�WZ�%��}�C�P�F��j&%݇�i�J;�d��d���n��\N!{�ٳ���^�]�;�щ&�R�=Q���WdR{�A��d2͆Nڝީ,-E���8�:tqa�t���nƓr؀��U�z��[���yu��T�ȷDY99�҇�����o:��ܶ��d̬� #yՍ�V�Țv�wԜ����1��A���a���Z�QgS̄#f�]ϯ)�4��0���Au���^8�ov����rD֫R�ʼ]tr�T�!J���v��n���(���!�Q�h�A�moFXLug��d�Z0)֨��m:A�C��L�fÓ4�M����"�]ŷ�i�ǪB�y�����Y�d��73o��O\�.�l�դ���N����m᭛I.r.�(k�mǍ枷��;�e�7lB�ftn�7¥�y��P+]��y}$?Ly�,��S-Ch����D�q �G.��8�!��J�Q�����j��T�8)�,��41\,Avq*�5�cfi#]�
5)6V��gr��uL�&Weadh3x��s����u�(�)d楑���w� &'c�엔+��v���+Gu��6��F0�i���m�5O�����ƽ�G{u*|�<+�(R� ��gF^�[a9.�
yf����@��2�=���9$�_d�@bq.,+�m�g$��9C.Լx3FV��t�,�s��j"s*�Ћ��@ 4u-�%uսJ��Zeu�4�TR0Tٖ�t�F��37M��HUZ�&T��*��̻i�h��.6S�E<��\��]�0PO�m��ݗ���k��L���َ�;8> qf�b��Q�{(U�z�% ��A�
z��F=�/#Q(�����u�]RN��^ź�`�E�:u`Q8!�SZ���X����>���յ�����J��K����u��u�1(�Y݊��f��k�nT҆tc/v�v:�T�3CŦ���=���cvu��:�*c`Ys5��Gj���!<���,�j��[�aA�xa���z��U��j��f��)��>�dSE�V��B�f]��r���j��+"d.���m(u�,�VT�EVq������Y�R��ޖ��	v:D'^K�!Q�.�]2z�I�p�2�TG���ڎ�b�d�7B���e�3�Ze�յ7HI�)U���t(`��h!$��A�l|�����            -����镛"	Ҭ���z�c5��Hѽ��ҕb��/���ٳ�4�w�XaIx��Ӄ����ޫ��,[���<�kM������4�-}He.t��� %*Uv���]�з��d���Ym��⿹��<��Wl@����ym�Ɠ�o7hXVTl��ֆ A-w�3�����d3�V�}�|V�P�����|�6����}Ʈ�\Z� 	��S���̟dV�Ө�\�m�6`�@�Lخ��L��R��p�O7��V�mujSgDqG�՜ؔm:os�q�O{'^�T�t��	H���V�Y.�J,�NΏe.$��j��f��Ji�Q���;齌@�K3O���X,z��-Z�s�K����s���6�n���1�L,�����7>V�!�3f�%M`�l���O5v��2�<����DTj^z�8    �3?]��l�H )$6�%1a��Hq�$�/�%2N$4�$��!L����E PE�Y"Ȣ�H�%�%0��Q
,����T�JdR!B$�� u�Hi	C	HJb	!
H�Ł �E$P��E �IL,�I,��`,��Dd���	v��K2@�I���"�܇uU�M{�Ƶ���k3���������[��nt/��c�n��N�J��U��E�o>����8��}_�U(V�gb8�|h�WH׿q�^�#�Ϟ5z�vS����A|W)�Һ{����icؖ}��b��Ba�~����*$�X�����K�~���y��/!��Ԝ2�}�?*I�ޛA�Rܠ��;ʛ��*z|�p�/�v_�oOT�J�`rbNt�\{ݐ}Y男 ����x�{7��x4{s��;�8�|�V��E�&˩P���R��0��o�b�� ڧ�+��2&�秺�������S����]Wq�w���ϓ�q����a�Np�T�I�Q�[>�=�����A[�c��X��f9��V2�4���̡8y�jUoM�2�t��!���>Up��j�ð�G���wN�������.���ܒf��ͺu�%)�4A���_�9�5W���(�n��X�{)��kf�^o��xQ�{1�+���!tw���c�������;Β{��v\x���׭�G#�A}���ᶷ���e��δ�m�xك�Ǵkxﭻ��q�)�����kh*ZO���=�!�JZֽu�fT����=��{�L4j�~sW���}[Q,q>�v��Z�6�W�'+�p��]�ۚ��w!��j� ����r��m�V����Q���;�N1�'+��g����e��T
���ĉ��y���ɹ�׆H��u�����G�w���Gǎ���NO]��;Ҁ��K�oG�q=~�ât'��劊�콊�.�r��oy)Y6���4�6a�S�����ߞ�Z�~������u���7K�Z�(���9n\�s�R�y���!`�U�l�wn���2��^G���Gחf�b�Wx������{���7=����\����K�ܚV�6�TS��y�9���neZ�Q
�%1�i�f˾�5T5�q�_#<��	�'��Z����W]Lg��e��oOg;oO!^9�!�D��.j{��]����Z�$۪w��<��-=��{�+�c/KI{h��z�z�~3m�wgk$F��&��D������=I
]��(�_���԰�۔�zˬ��TE�y͏w^_T	G�3๠udĦ���3�j��Ŝ.!�]��`��Y]�r_���=�n���$)�xeH�v��)%1,o!o3s����/6Vs�\{'e�ͧ�L� ����+�9�뚈=���wC=<\��w���sv��u�'txeV2�Xz����3�����0��
u&RD���\lfln'�g7���w��~,���J��禲rl�����$��~��e5��?[���p2�W#�|k�ڳ��sP�Q�ײ������i���;���Z��P�j- �)_�Gz���0�EK��9��Z�(�&��M���il�7�����=����ѹ�1��7�*';�����3x�Xi�5�hC����#�oopg���g�W/xE��.���-߻W��K���:7v=�wE_��
�\gH��^�dOy�UP�N�D�٨�c�C8�;/�:�|�q�p��wJ���\�D(�����;�+���Tb����G��)M�ܷq�"��<6�&`�ޮ�{[�t�vu�$+�P��_y���UL��y����cw�o�yzcag��β���bxۘ���C�y���������>��Y��p���1�y��*L��̢�����\����mz�ҡ�u'��f���w�b=�(����t�"%���%���-I�u�8�c%�s��a93�{�U/�){�!�zT8d�Ě_���/���l�b�=�ys3�ӂ�.�~�<|�;�������z�w��c��q�Z9�<ܘ��_\{�8��z݌#�Q>�Ŵ�˓E�����\�B=��p�B�s6v�����7�bʇH�[�O>\�7n�5�y�"��]���\2�.�7�Yb�D��bf�nVo+��
�)F�m�b������{���ߦ��|�����J�O��O2&�]�]b�9�i����{;ƭ�;�<}�e�9���=L�Nռim��>~���:Ij��=�jx���W�u���k�ayV�Y�p����B_�)��D�J1j=�{�E%
��b���[���P�Hr�+~����'�6^\H������14�'L�Fh/(�T>�ѝ�RЀ�K2��������mª��zWѭ�yN�)��S�֟��ܪ��}q0Wϥ_���edF�A�l��ʷ�Oh�SP��k�g���F�Xwv����	sz*K���a������N��0U�B,;����"���Ĥ̫�_ajbuv�]7��r[&>��R7)N^��c8i�$j���]��{��:�^�݃m8����Fq=��{�/*��H�Ƽ���k|IϬW�rѷL���C�7L�������[��5ݺ͏>u*b�91"�O��:=~8�6����e�]�x�S�õ�s�U�{������sݏ.�YK�cu����n��x�J/��gz�:���Pη��Nj�'����i����coُi�:O�&+�=y��fzw.����ۏb~==��c���j�����S�Mp��[��k�O<��	�;�M��nW{6=�;��ۃ�c��ʲ�b9�v�D���YlR�x0��г�kP��Vs&>n0�4�����/Z���C���#�ۼ�W��lj�jƾfh|^�RE�Ոd�Xb�#�B�9�|��Mϊ����hg�R�1:���!��G�����n��=��������T�=��y��5R�x_����s�A}�әI
]��E,�N8kW�j֚��l*{���PR�&'�~L�s=qnv�cFW#�/8L�z>]@��2��N�)�w\���{N_�i�aO��<�g9�>9��Rrs(!H:ß������s��S�輼��<��u�Tָ��ǩ��*ששn|��|�e۲;�SX�޵����>n�*���t�*�;��w��ۮ����ɾa�pS�E�~��-;�w5a�q���J�j��6�˳4ݕg`#��o;3�ºU�sb�o��s��ZTvnU+�W:h�"F�9�7����%�9��hR�Y�81�����ϋ��F�O�r�T_D��>|qh>�J95����#͛�f�r4���N��{���2���}^����������<�\ى��v��eoQx����Ӕ�g��f�U�{��>S�͟Y��E���kܝuu�k�i���׫�(#g4�I������=9���oի������3{ч�N�[�X���L��E����$X�T���g�Y����f��=����f����x�B]ѣ��q\�^b|���n�Q�W��p>��+X_{�`��H �	) ��l�'k/kw/�CI6�S8�6���S �j�&��0n5{������a���2ϓ��P��x���#Wl⹜C#^W2��Ҹ�	*�e�c�A�̌;鎆	�A�?�يxUŭ�sV�.1;�6擒�����(9^
|��8���.5N�3a����+�á�6�~�9y?=]FOw�<� ��nPh�3w��}J��p�#q�{�94��x��T
DǽՓN����c�sǉ��Խ||&J�REZS�ǿ9���m��Qykd5�2h��ޥ^�,�K�K�r1�쌍u��{��`yS�6�V:$dۼ��yr#cڿd/O�d^,����ܟ��0c�v��<�.����U��(-v��X^o�����i��z_Oswr��hֹ��ɳ'�z�0�����i�{2,�(fc<3��KA��J�ubN�Z�p �~E�Kf�έ�;���YB�F�sz�MwSh�&[R��:!B���[�Y�<�$F%�X��a�&�e�̤QŦ�v�� ��:�+	����AH_%��3��{�fU�z���&f��[9���+U(U�G�էfW<��ef��V��V�]�P���Z�q�R�K�w1P�dz�2�ﻄ�Ѣz��T����D������Va�	�d�ӻCon���J�Pu�\�SW<�i�y�k�ՂB)�ձN��%y�-�,�vKFw��9�mLܭ;�,�R(�]�r��4��3��9�ŕ�cd����F�T�V��-!4z�$o&�f�s�l�}���qCW�ir��٬J\���H�oX��C���0XnL�{�P����
�;�U덌D��o4��;V����r	���zc����s/�NɊ�P�����w2ы3�+Cu5P�'��p͗���r�Gi��w���q��ls���Aې���_�N���=�            "Z��Ԝ�[��6�^=K��Yn�T9T״�2�R4*jK�U+z����N�[�/�J�ʖ��W���"�h-Y�ӭ�<���][�[���;+��܅�lB�~*��\�-����V),}X�9��F>�V��-Vp���`�}��ąf�v��:���>�}���QY�ѯ��%�-#��8�^��xu59M��]u���[�Xヱ��6�A�����^��=Re�x�#��v�Z��R�x�n�zo�W��yM �K��s�T��;x�h܏�m&��t'��r�-U�M�9+y�X��:#w�^}
�x[S4U�L���Nx�����t��.�X��cn3Jj����[s����U�[��<A�{FW.��(�1�Үa<��d�wt�l�7���/+�[��bfme.��M�w��X����&2%.IY7��g��    ~�+�d"�H�CL&�Y�

	,�AAg�@�,�H*�D@�)X)��]$���,��H*���$R�!t�0�.0�,�S!$�!H)0�0$�0�J��P�� �
��Y	fHRE$��P���X�]�5��>��[W���wz!��8����5�¦�0� Nw:���Z�|�!QB�?V�����o��K����[ތO^Dw!�����v%��wr7�Ϥ�6�4/�'����q���_�����O�^B�W��_�����~o*��zgz�)��Jq5�ڊ�V����t3 ���fsgޟ�]��T��ߑ0����={9q�מ�Ɨ�o�k�U����QȎ'`�e����[�'9y�pz�n2�˚�	rϊ���u��s�N�9N๳��|߱W�ۭ�˨���91&�n�ޑ{Ҹ�����S=����v:
�:�T�r,��O�o�o�Ӗ�A�;��n����k�=�пi�z�!��;��j*<�]�{��8k�/-���\�9Ѧ�[W+�:�;�� ���YK5b*�L0�ɽn�.u�����I�؞R�� 5d[���J�D����_�4H�Q�1�mb���ʞ���^��U]��Ϣ���{�R[�N1��i�����U��d�������/'���ֺ��ne��#�=��n~�4�Q��w�+�g���Zv)�� 5��\������!��C�>\�/�1�yϒ��w�{4O�;��_�r��m�G�J�!=�s�U�U�������"�'=rlj��L��25�[�y����Z�����3�.�]�U]'�1~ݾ��[��[w���i*O�{y~�����L�81�&V�s�����b�~��������?�.U�8'��듺���� ��������f���7rb���j�c�����K�D�C�紆�Z���c;���Hꔷ����N���Pk͝ZV�ym�}�t�qCl����{��>���#+Z�����/���;���ؕ����k%Aw��3������3�^,��M�)�Z�Y>-x��siy�3�+�"�k�7�O�4n8�-�hv)e�=������]!W�e��Z.�����h?v5��
�q�ȫJKQ츑�U3ϫ�Q[��m�k��f{T{�x��n=���^�T#=�v��Ȫq�,�+)�NwI����͊�$�s�p�T^˔�>��i�RRi���=���u�\��ed�Y��>�0�y�$�c۽W=�^��W7m{w�;�c��,�e��a�'Y6�zW}p�Hb�J@-�!�4��W'�`�m/P�`X�Hy�oX֯��-^���x�~[Ҹ;s`j"�����{��2R5"�����<Vw��5���^�s�����p��AYu�1R\�t��ϐ��S��jn�^�l��Oe���lf�U������u�zn��BN$Ӷfk��̗��&�s���q�R,��)!����a�u%2M��ڻ����nc�V{�s�סvN��:ɷ(gT@�L�a8ɫ��|�c�	��&Ru�g���,���:�2ar��L�{���k��c�����K0�2��'�T<��Ԃ��8ɶ�@��^r�;Bɴ����&Yt�d!�痐�=q�o|��{�=|g�;�H��@�N�q�CM2N'�T4��B���$˶��	�y	���]$��'�Lq��_z���o|ߏY&�w��=IL�'*,�l��	�%��y��t<���g'�e�&U)	�f�ϱ����Ƶ�s���a�1A6�Y)�q�۷�����$�M0/TN2i���0���Y�	�C�)�!���a��߭���o�{{��2K%2`i����hY<z�2N0�ݻy,�w��&�P.Z��M�i1j	�R�r�1�_^�9��E�m[W�}�c�,�d8�S)0��N2`{�C���dǨ�����Y�$�*E���P6��V��zk=�9�s[�zC��P�)8��Y	��$�CI8�)4�a���u��}�Y-�[�%�9�%8d�����}������H�æ���I�\�����.��L�2p�]!�PC��6�P���t�d�N00ɶNY�9�Sڶ+���\y�l9\|77"����V�X�KP^��-�{m�eyKi���8x�%.��r�o��e�^F��.P��M8J͗��U�[;��������l�u>z�Re��D��sTC�K�Y��%�Re2q� qn�fIv^f��m$��6���[�߽�cƙ,���=ʁ�N2\�,I�{D�fIt&,�d�e&�T���:�q�'�'X
[I8�������}����q��@���&]���d�'Y:��$��Q&XdP�B̅���i�OPd���s3��J}�o��9���,�S�(��M�I8�[�Ğt�bj�y&]�u���U���A�Ri��*��M��߻�o�=Μϯ����1A�����I�O!��Hq��/�<�6�$Ӷ�I�̞�6��	䆪�Y0�,�מ��c����@�`z�� i)��'�Z�l�B\�<���gU!�N��m$�'�2��I��&q�e��g��S�s�{:�.�ć�S�S!�
I�$�I��ڒ���̞z�`�2m��`���_��i'Y1z��'������/k^�:Id�&��k�!=��B�Ctm��C��چ�I8�0�O9d5*�<��Ũ�Gg�m[����s�ϵ�׎0�@��&�t'��2q2N��vćQ��Y8�Ԛd�j�	�M��T<� ��INY�M��{�o��`u&\����՚6�yL
d:ͲC���Y[�)'M�XS&�����d���z��&���ϻ��~_8�_7G�?_w���U���d᠃����h���|/޻8�]�j��,^H�K}�&z
̓����ڄ��s�@P���e�
Eg��������8�큧��UU���g[�}�.�Y�*IN����alԜd��R�B�u2f�$�)$�M�ۗ���5DY4�W�ky�v��w���ɶM2m)	��컄��{4���JJa�T �1S�$/ʂ�RM��I�R�{����ݿu�w�=%�$�}ڑI�(�m&��O2��N0�ꁆ]��� ��N2JM���C�Y�
�i�w�V���ν�x����9�I)���%��M�).逡��a�Y�-FS�'m��C�1bL!�I��ox���-��\�|q��B�4��N00��OO{W�Y��夤��~T�L9`))��Cl&�FYt�s�&P�!��)���Y�=�랷�!��,�]&�!����O>I�8ɩ�X�(ϬM6I<�3D�`Z�q�e)2�U�Z���׵��>�Haک:�P���N���1�<ɷ�'��q'����|sv$���,&kԆv/�Wu�5w������f��z��Ikא�@�(�a���i'P�jq�q��G:���0�'Y6��L��=y!���v�8���g^�y��S	�{�If�I<����I-z�עi�Y6���u3ک'Xq:ɴ��=�$˴��:�6�k=�{��0�߹p�d1Te2K�CL:�Jd��N�P�`y��'���C��aɊ<�u&O�c��	N�ߌR/�uhha�%vp����d!��)+'�O�e���^��C��~~[��t�E?_O�1X_������Z������cdj��'���s6��}$�8�����k|��I��'�>��2Ì�I�����T���K�P:��$�N&}RY P�&��2U6��P�۪�h�+ؾy�{ m��[r�q&�0�oڄ�.��`ŭ!d&�U8� ��`^��m'��q�u����Ź��}�o�׃,�x��PN�ä0Z�y����>B-Rm<�u�z �&��I�7��B�N��[�8�L�Lgx5��N=��u�{��%2u=��*��f�&�j�I�hf�$5f�!:����e�JBm2Rdk|���n���{��l�]�-�$���U	�L�K0�d�d�Ci'����HL�P!�Pd��E�C�:��6��d�}�����wǠI�۷�����L�@��@�N7M^�Kb��RN!�ԇ��x�S)z��$�h�!ąt���o6����Z�k�P�ש��-�,�4���/%�'�R,�n�I&R]�j�!��|�.b�a<���� P��\ޞ[6�������I)=�0�m!s���2c��2k����I:��d��T:��L9L��HT�O!6�>N���k���!�I�2���q ��u��e�u���$�&�]d�d��ZJI:��I�,�C��6��v�o�v��_�{��	�y.�/�(i!�h�(y��T��i�`,�7P:�ǩ1�(Iz�I����'���b�-�[ǩz.��'\�i�tW�3p�����Y�U�^);|Ve~o��݇q{����g*����إL���rrL����Et\΅y*�\;����c�s~�����	�I$	-�w��|��B�'I���	k�Y��%�@e2�Bi��m
d�fY�M��=F�8��):�u&���R�~�s��Bq��v��d����*����@�Ik���C��Hq���P�a�5F����d�j��5�Z��}+Y����d�'Y>LԚ`m&\�����q)	�.r�2˰/T�<�=P:�X�C��k�4�l0�:�^��}���m�w��|i�$��Y4�a�a�'Y6�<�q!�J@4��`f����y,�lÌ��s}ֳ�M<�c:����S'\3��P4��G!��i�	������:�i��qp�d1TE��U�`,�,6ǷW���:�����oĳ$�L:��C�q�l�p��D!t˦���I��'Y�y�ū]s��:���sC��I�ﮑ�mf�v�ƴ�c+���W��[&K��ڵ�����ߖ7*����Mm�_y�ǁ孙c�}���)gU���6�3�7"hF�Zn0=Փ�'<��.�30���k���\%�����?[�4�,�(�y\2�Z�FdA�]��J�`&~|b-�_:}n�Ij����?�z�f�uMJ�i��8&U�`�U��\��)���o��T����g�ϗ�~�H !$�$!k��y����M��{�N�A,�z�ֻJv��gf�1�]����:��:�TǇ&$u�ن��1g�rO��V;o����:z�|RET�r4� �>pG�s�^R��=�Q�����we=��׽E��w���+��VE�x΍U�m��5�����?#����ǵ�����A+��u<��+��L��6�����]�/�븞�Ct����J�����Vo�Q�'���O
6o6���v���&�|�׶G�$<���<7y�^K�1ԗ4��]�⺭���	3B��{ƽ��[�|�t��An��޽s5��&���g}|��'˘�b��u��T���K�(�Y։�U��r��_�!a�K|�Wc��0�9w�m�-��v'y�o�添�淃�I$�R��) �H��� ��a�E�
H�"��((�(�Qa���yޘ���om�՜TLk*��M���g�'Ȱ�mwqjxZ~W˼�I\��
:U�^ý�1�:'�09��{�n�o�uL9�H��:��uy9p��߱xI��ٮ��/h�I܈�{d�uI�x�r�=�d�#��܂�Ǒ=	o'=ң6^�ś��h���>1�~�7x�Q~�x�]�/s:<���D�E,���zյ��~"�Ma%���޿cގ'Ⴝ��݊^c��i���6�܁��]�jz���9��l,-X�ߔ{.q��^Yt�[�U���+\-���qZ�X��Ǵ��+$��&=wC�@�����u�z*�f�5[�'[0�I��ӋQ�����Җ�d���)��V��>)w3�9�qR�������y*T�։����y���fC�U�B` ���gX������z>�S*���ژy���vd�K2�*�d�W�C�w����-���RS{Xl�(Tٻ�s ���ټ���P��F��(d�Zt]IY݃�V!	���lƅN���v��,��sT}��k}�pUwo�Һ�۵>�Yp��r�M=̕/�14��%oVu�3S��WvJy`tu�T6z�,Э�XF��ܣM����N��֭�L�"�jR��ԧ�nk��hp��`d�R7��������+B�P�,6]
����=���]^p�u&����p,���Op7������h�G��K�C�vp���Pl2�i�+�n��C��C1JWt�
dF��z�	q�J���j�~���+�G��            �F^���w�GUb����/k��e�Rb���q�vt������l��&�J��4ǁۜź��7S1LN�=؝�)�:,w��G�+۱�3iaV�^�s�X�M��Wt��fr�Pl��h�]װ��&�P���y#�`p}��q47eYf5��x�pPh�YV��-)�E���Z^�+�/1q��_^��m� ��wpro����[�,+ł�QBa	!��L�Mh���[=�2qb���N�u0':����6����CC|�w(�(B���-w^��EۺɃTvV�����(%p���k,�W^Y���
������ZC'rD3�ZכB�ʻ�٦�;O��B1�)�Nmv�����ũS���sR��*�
"�=o@��짩m�[���i�]b��gH�}ǥ��.�^ݰ!A8�����޾��~�T�-]�z��  �s��9�[��O�O2�������(��HR"�$�K$�B�"$)$��@j�AB����O�,��R�$�$�
`�,�S)���Y"���d�d���d��R�&%�$�E	
BS�� �̀R�
AJ�$QVHR@�/k,$�dHE�F,!d��R,Y9�@<g:�~c��U�x�N$��/wz,�*)�q���f����!�"V_q�tg''��������k����/�����)����N~^����V���_��Ҋ�H����kJ�>>k��g	�3�ח�y )[�m�Iʞ}j/N��.�Ѕy<��s,�i�r�cM���{�!u[=���bM�J�P�v���ho�;٬�c�O��s�ljr�^���<�$��gk����e�����0�,��Lk�|���iwE齏��ݡ�k��g����E/�˳����߸�	k�~�O��/Б�<k��n9�'����a�*�m�5~s�<>5n��|�E�;�*ys��D�]�AG�56z�z����	�;%��z�O�vY�k�%[Kn7��u��#���R�
��0���1X�\�q�|�Q�����[�Ԩer�V0|p)6Z�KI���GR������k´(����"������>u�,!�����	��n{��[���c�{��}5�7

	��V��=���Em[����eyvf���E���pcw2�oE���ʋ׽�'fq^���f�TW� �ߛ�ߋ������ڷ:�y8�� �y�}^���=㣹5��'�>�f���n(�����gm�f��W����]iO�eƘʲ*��a�u��@��=�#�W�0~�9��Oo���^�x�yq�}7��OԼV�9�9�n���e�K{�����9&�����5S��s�]tFr��Lr�^�ɖ�
f04:ufa�KKR��t2�՘��4R�U������}�F�8���<̔��?3b���RvUq���.�Bp	ok�#��L�͑쮅��2�k��"">�"{���-.|bQo��q�3̢��gu�Cb��O��=Y�?�?Nr�i�T��}�q��ff�uN)F�F�򘥝T���ǽ��;�=����͸��!�9�j�K�~MYj`��wQ��#���W%n���Rc���A6�-��\�"(��&�����fV�͗j����B�?^W%@�k�z�FB/�/�/�]{�z�#GDq�>�v'�"3)�9�q츞Vʋ�{D-���GKG�y��5���u��<����O*�C|��W�e����;�w�=��sYq�j��q=��EDSՙ	�N*��9�,F�t�Ask�l��t�Wi�8��Wc�;��o=�h��K�@� ��^�<b���w��o`k�m��K������&.���}���b$S��������9���9m`�|���j�������N��1���}xs^��_��ӣ&׷���X4�9�&ﾷ}���bW���{��%�I�3{U�ܛ�~���o 8!��/P��ɏcsu����r���=��gy�H�\�{K"N�^�'\uh�܋`2�&��Eo������+�����6ʄ��I��r�/~l����a�)I������_.L"bs'+)KZ~��=٨�M�Սq����3����+�U��}����P�I��=~��9���}�]���*��9��;���|�޻�y���3YM����Uc*.����]�&:��LImn�꾄�z�`�X���266�ܼ4��M1ͣ���Û�Wi��Ge:qW磌ꪬ�xS7�	?|��P[�����]��bi׹�����X�9i����[];,w���iz>���Z�I'#��Sj�Lp�w���qUY��T�`��q�ތ+�h�m���yӯ�n�-��幊o����}U�y���=�����N��OJ~�̷@�XfiU�\l�������*bo���&���b�)�I��e���ތ��Ѿ��{�t�|�'�O�ǐ�6�zy�H\Ul�y�=H&sw����0]�Ž��v����NUe�粣��C)I��g|xҗ�w*�[��"�A�˥��T�n5�&x����M۞	B���Cw!�+̊K�42co^��;Iu �Ջ�ͱ8�i���Ҹʝ����w�ޫ��2P���1�r�)���4>/o�f��U_}��Q�种l�E��|�~���(��eO�9|���'�~p�穻�j==��*�2��	٬ؚeW��s��8��[&*;
��ל����{�54��G��U������]�T�nA��{µ�����N{�_>�^��l4��;y\�=�^O�r�{[o(p�+zpl� Z��!GT��q���ގ��>n��ye��Cz��.E%&5�q�⤕�ֻ�h��{����Tsg?'��U%��Fc��ڇ���ot�b�^��Yz�E�ط���Ka�8��6������i�^�z���K��S�#,� �F��N���x;�:Bv�Vъ�Ÿ9l�B�Y�q�����雗c��;��0)�a���Z	m�8��������s����{R{�E���ȝD[�K�Y���ݴ�ʎ�����ƪ"FF�i������T]q�0��ڌK�m���ta���1��㻫���X�i/)s�*�r�z�}����u=�4��i�.�j&5Y����4k{b��m�!{Y�9�F'�/��r�i�ԨE���z+:������;�g!�T�>�5�(��׏I����r��	��R��j��t�2gV���fw^5�1T�5S�B�ԙN��U-2�k8(����W��MƵhX�Wm�>!˞��(�/�T�,.�����F���ënھ����r��/�\PJ�]s�+����9j�pM0��5ѤwWU�w1��� �{�����C�fw�B��mogҝ-~�#����M��Vw�%yObھ���S��������վ��;��S��_G��Y2�-z6������V���W{z���y|�;������F����-�{{0�3��*����:w��OYNZ���'o*Y���"��g���1?5ڢ�~��.{�_f��Ƹ���7Ο5������Ũ��[���~��»�*T�|����J���ֻ�c�k+�{���ǟ4�܉2�[&�?�~�:]~}��򷜱n���퉌�*B�[�4*v���;�3k=��R�2�����V�=��X'#�aO}6� ]$oi��$㵫�e5�cAօh�$r��e��
��s������u�ԬTT�{zu�c#�չX{�P	�����kse�i
2'����ꪡ�=#sϣ���7�2bX��EI̧.��(�w�S���R?d�g-2+k�e�ȓ�Ȃ�c)7^���S�|�N9�o�o�3U��9]^;,*m:�]}�&�Rz��U�R�\GoF��s������/�\���RIO
�ex!�-����>�?`�6��e�v7݃O�\F��W�q��)䋙N�����.�6�E_{{��Nה�O#��)�3�̧[��`�3���u���x�^(�ykyq�i׮3'2�z��skb���W�y��Uqz�:Ϧ9S�%�mǅN*��8Hq���1��-�b��<\)�Z�,�ko����wF�q)�^(љ��L`KS��=�F c4KU���ɉ.����;�uvӹ��R��vaq#�VNJ��Mu>��\ZB{����G�(mHc���?UU}��)I���ߟu��(
 q��������vfu��{=.��tK����O�P���x3�V
��pI*���z�����+r�
rLf����?\&H���Ǎ9�X5�����3�W�� B���l���ɔtkyH�e�x/��U���C=�̾�

�N�M�.8-ߓ^����=}U�/)�+�:D��|���Vܲ�f[��TKYq2\z�vk��"*e*���r�k����8׳���� _�ly6�c�^CBʬ.��s��uV��D�fv���)��X5�.&�M]N�Q�-��x5�?A��o.wo�TO�ؤ�G�V7�0�+sȚ5r���1��5���閪��=[�EU��:��܈��Lu��~�{�������B�j��T_Q�^s,���\���2�7��u��%��Y�b��3������(�Ө�:qAO;�h($��r������4���!E;�q
�=7�͔/��4�h�Y5�=��MK':�fG��v\wR�5�����)����fn���wJjH�Ԓrq��N�R�⊆���R��Ɂۇ�®��"M���gM��[���:��JBZB���hu��>D�F�5hU�&JzyК�Q$c��s&��v)��U`��D����0�[���!Q�HJ�#@9�K�q]��[�eی�d�
q������VGuضoj=��m!F<5�����0^jȈ/_&a��й�#�4�I(^�k��1v�:s 0ス��Gׂ�Ln��rr�HN���O�HW��]Ү��z��N|��P��Q�M�a�x����Zk�	S.<�|��WnuC�6�lt�v��&��;���e�w����e�F�d'��i�e�a���^�/^�!���R�_�ŗ��            ɛ�3��HN�1�gap�2T�8G�k_W3��OfYxjd��!�1+��+�(Vҹ�k��6��k�D���P/����W�L��`�%�r�%�ӥ�NmɅ�Ά���@��|��sb�����%���#U+�48��cmCG/�@�}x�؏��rsE�k��}|�\��H`��)���Q�.�����R�ɬƯ]+�ﷳk.ң�����]���O>]}��1�^��{s#�L���x7��p2�V;�'sP6�$��	ٮ�c��~A;��t�,F�+��lD/A}%ޠ�t�U�)�ɜ(c����M�ہgStmB���N1�݊Ի:+R�0�'Z")�m�6��QT�lIB�����`���٘�H�»^c�ӕN؆_f�n��X���ujR�9[9֥Y�[���CV��y�Q�B��g��� � ?�{�OЗaI� �� ���:��E�Y<Ɇd�ń��2y�RE�R�ʪ�QBȳL)!�t�����@�C�0 �%��UVE"�Yz�����I4�Ȣ��R�U�H",a�S �E�BR��*�1n�H��W�}���/�r�pYF���I��!�6L��zzTπn>L`ߦ�>43�n'�c�/�}_WԎ��zyfZk?��B����b5u�j^����'ټЦ),ҳ�/�b����􌾣[$�����u1�����L��v.�����z�yZ<&���P��0F	^����u�	���h��������dW�\+����LK#M�G�~|,hM�\�v%ؘ��M^˟D2�'Ϭ�������wQ�+e�X+�~�^�U>L��S2��ʟe�H�'�nu���~SC|/٦-�E��w�\�Z;W�j�������L*��2����U��(���.�Y�~�`[9���݊��W������d�Pi��מ���m������yh�QxT��Ò�e��S��_{9��x�}[�F�![���� A��Z�q<&�/�5��{�=Y˔�=k��oL��*�,ۣ�ʟo�����f]��_o[y��ؓ%�y�P|Q;��/%���6�HP��'o{�[:��z����֊��J<�-nL#������ڞ�`�X#Gb\8V��h-616�u{\���J��ܷ8eQN�
�A-��h�T�`U�Xh��ۋf�����d�o�e/vΦC�U�q��j�&]4\9���M����W���o�ݐ
�����yԗ)�3Ʀ�T�'�˅.T��T�E>�G^���<<�@h~R*�����D�vc���q=��)��k�W�yNm#�`�5u�e����
�Dt?���������QO.q����k;W�}"�C(P\�~��}d�Ǯ�n�fJ*��7���_����\*J�c��ڬ_��\
��{�i��Oq�V�T�j쏏���O.��<=�^G��= B�r�M*^�/�j�wfϽ��^K�w*�Z��5�5����z{�/���n+�.!��Jӊ������t�y�u�%�	�~\����ox[-��68��ͩ���]܂K�	36�^���>�B�Ud�?}DFW�m��F�����Z8 ��ګD7޷U��Yz�ހ�۝���^�^G�>��,e�.
`V�b�A�G%�hBc�]��ݽ��ǫ�6Ug�&[u\*�
����b�VG��ܕ>Ǽm��ҟ��|'��{��?p99��H��hυpض��L�}����� tP�
��;)�A{�+x��(�$td�OI=�];�ҵ�����9����J�J��nzjZ���y��ڼ�h>�f_ۈ�|�Rip�F�k>6���<U�����nw/�k[omN�F>��yG,�Z�q<*�p���q �,{�zY�Ѩ���]6T�&�ڏ[�{�Yh��K�kG�Fr[�ǲo��!@�r<�P�h�Y�nT����=�����-�oy	�Z[F��:&�s�D�5_Vv*��n���X�M=�١�Id�*z��,+�5�m�m���E�k�B��͔�uҡ�@Ԭ��R��9��������~�,��`�M,xQ���k�ʭV8:�`�5ε	iG�+d�y��t��i�v�J�b��rT� X��v^�j�o��Ul�s.�k6�����\��*��I�Lr��?}��������s���%"�d֋4R� Ⱦ5��t̻�[�d��o;�x��i�.�`���_Ϋ�(
 ��Y��
OP8m��X��}�g��t���Kz�a�+-�9�WM��u9��&��cqdV_{�~je��7ē��j�������[��Oi����X���y��[�8^>W��=f��;����#yYH���R�j1���\�:+t׬�z&M8H���J#||1�t�'l��~��21���ϝL��/�JK��E@s8,W;[HժU��o�pV)~k��1��V�hu��4o}�����%�z�PW\������c�][�����!�����{�0u΄_�*.s�;����"v������]���_�;�B���m�'b�ӭ�~��'����Q;XT1?�5�t���@/P(R�89���Z%j�u�26ϚU����ثa8�dw��N��j����</�x`g�bDV�C""��ͷ� 9�;w��UΕ�����ߗ��5
�I���EFI�_c�o\e���u�~���f��u�1�����J�B\�S9��;1�������*�qQ�|uW;Z��,p�`��u
�^�׮�i���2�s��?���s�*��
�G�}L���|2���~�yȽ�������wY?0T;U��og����P�F�Q�~|�n��e�z@�,�F�u�����^س�����U1��]��P�=�d��G�C��wy���ߗ�'��_��"=++���X6�Q"�H ���啙�F>�ΠXc:��b�.����Df�v	��bÕ��l��ڗ�w.�v��h<i��gE�R��,%�VPL2d[���_}S��lft���Ԭ���9x������~����t�7��5�y�֒�w��lo6Ҭ�ܷ֬}�[����U���X)w������T��A��I��Wuj烸����^������v&�B�3<�^�A����`8�]�.�R�vm6<��=~0׵�v���V(��N�<WXtxV":8�.�񥼍��$�p�}ӆ��==���xz�#��~�<*��p#�h�Ŭ4U����4�I�l�������8�T�١���Z\8g*�T�w�*j�������;�� R��'��0�צ�J�4EZx� F*fk~��sl����� `~Lւ8`�DÆu�A��Y����zw^��V�[����p�A�4��<
��ue�+���2�\]���yg�6��g��]j��)wW�K�]s�f&����(�ۀ�׻�d�*�&��ES�W㊈ev�	��K����_W��c��p�ϹT9 ���Lݏ�UwW!e��5��Le7xb~kƠ�g������^$w�C�\*O���ڬ:�au�&�ޟ,��8�^����W�K���`�G�����蟼�{f�{7��r3�+�y``�\��GPu�g�m�a��4��AX�O{�՗^��Z �P�eq`��c: �5���[���~�H�Y���O#��s�U
�s益vf^�U�$05���SS��vdc}�{��o�X���eVx�<-��?�
��&B�uM˩��|��7���,�����S>����3'4r!P�һgZ�#I�ҩ~�yKk���	|�d�WRդu#�tv�4z�ᓸ��_{��N
�¼1S��S6m:����Ѭ�ySʞ	��o�W���;(�4!*�J�
��̣�����u�W#Vj�cJ�v��cO�f��F<I>�7%��N]�+)p{&YF��#׮��#p��=q��%㧌�?}�}����f��Dht|�R'�
�q�U`x�Y�tM�W���y��c��*ԫ0r��Ô�`�<*�p����A��{Ӭ���{�(z&0:���V�<��R����Y�Iݗ[t��x���է������N5���
5������O��Y�;g��ε�d�L?{d�rŽ�5�W��k�郆q�D�G�H.Fe�o���k��ү+Y�&���HV-�>����f�G7�YQ�OїX�`��QV�7����δ�W�8O���l� "������V�^�hJ���𫘴pT��,*�>��m�l&�{n0�U���y=��)��LT�	���.����J�����'��!{�2ܢ�d��Z�)��Na��]7���
�t���Pc�%���B�t��eͣK���Yfe'�4fS�Pjȶ�E�K����۽���N�@��ή���n�d��d�hv����"�9��Va;�5~�>��yw��~��zG�I'��ϊ�����۞��q���a�S�^½
v�V*[�.�����o֥�L��jћ����K^N���-�xH��>Ǝ�U�U��z&Md������:sq|EW�y���|T��, �pi<=�ɬ��#Ww��L��(IO�eq{��쬢�������0nf��Dz��VC�'�<1z�ױ�gNFLd㉫�q.N�!P�Q�9e��|�u��o=�pMz��ޗ���lz���W��Rh�%a|Hф�[��=�Sl�H��w%͏Th��'^c��3�x�[ʍ�xX� ֠8wЗ��د���j�P��$+ԯ�l�l�O�Qڮf�x����n��̞~��3�C��Ds��8Q�:���B�7mX���M����S�l�o���&{"����] ������a������j���q�م��9�p#�.]����/$��4��t��J"�)�Gp��%�-Ǳc����E�9��W_��a�oƽ������4�hp�Tz2�㞲�<Ѹ*�&�~-/|��TX�p�P�Q��2�p(h�W����+��&�chFnNʙy}'�ԩ�w/��R���>pq�mֶ�ꫯB��K�F3j
�v*_ o�qW���+yx;��;���Ĺ�ӛ�9�Z WR������PB�3��wK��O|�M�����z�z�����! b�65�$5�U���o�]��r��g�x9��m�Ǯm"��2�纝WL�L��+���]{Bc��t��#������7p��uѫgn�DU��P��^'��Nf�фέ�h[�����*���s�j����t� ������5ܧo�ٽ�G��pT��6]��}g­��:�C��M`è��2���Ǣ$x ~9�a�i���)�8����y4��<ۧ\��[��vG�X?C�4��ɤu�צƅ9���B��Yi>-V�ަ���z%�{t�Dr�����|���Q�W�
�{3{#�!���Q�g�2Cݮ�K,�j��5�5��̌9���+��`_�os�,�q��޲W)f��īq��x�����J��f���U�sk^�4�j��GV�B����;8����i�ʼ���8'��L\6��=�\o����ȡ{��<ќ�j�B��jZ�e��:�٨:{,���O��R�roU��mN:��\�I5(��dne�X��J����R�T�(dxs�@��f v��W��նR��N]�ެ�`�4����9��l7�1�j��8 ��R�Y�G�t�i�V2v�`
�s�e�#%V��`[�b:�nbZ�:�H�ۦ���V�;�v�x�0�m��"\�`�w���A�-��ɎR{3�������OE��S��+hI�            w�E�gG	�X�ܐ�6�J�
!��`���y�/y���,۩�S�;�{:����T�q�]��k�Un��r�f-k��o&ؕÍ�vw
���yq-{��{|�g�B��M�Xkt���v☯>&�K�Qh;���H������">��{i��t7����^�,�Q��D��bH��ŝ�V@oCOt�zS�Y|��ƞ�9�
�ٶ��ڛ�<$e��ӻr�D��t�p�Y�3�0]Zz�R��p�؀��0
���o9���pBԹW��uʱAU��1�V�S��i�ݫ��	������h'���Q�v�'���*�Yt���2����&���v>9 �·m�ym�ʙ�F���j��ҹ��.N��Z+y�y��m�7�>�rc��.����'B=��^TR�[J��
0G��$�ȩ֔㭝8�kVu�� @ ��GLGM3(RB��� �L)����Qb���*��U������
��$5jU�����VS��XL3(e��*,"�% R,a!��F*,�Tg��Z�4�$Qb+ ��2�F����4����K�*��b1X���P�����+�)���|�u��V׷ksW�2tK��N��s��gs[�OiM�qw2PT)��:s���7���S�{�V*މ�m�*ڎ�-i�vhx��vO��L�s�z=#{��&v\e��܆��+F'Gl�)�P�u5Ui�j����gcp�T���L����FB@hG���h�hu�0ხ]ep�޻+�^�~�4��b�z�O�9qz٭������	B�:/�����v��]y�؈��P[�UqkU��i�r�C*9�fh}F��5T��LS݄S'����ă����W
��X���l��4v��_����0���u�7�/�	rL�ةF���aMQ-�?y�{��Ձ̍�Z���d��Q<�T���D�Nny�/r����iL��Y�o}S�8J���ɲXY@a��j�|րj�U��y����=VF�I�(��\VWA�֚��> ����<k�$4��~��oT�\��j��,�]��y,�ǌ�3��;U�
��r��}vE���wN���ۼ亁��y��S.����/ Z�[�.;����4��<�wE�=C�s�r���N�5�_�C��nI�°"`Th���Bu�׋��ޫ�t�+"��3��ַ�Nh���^��K���4쐱�:7�'���1�8<¸R�5�Vgg�.nd��Ľ
Mky>�0ͺ���ښ�����3fӫ:;<��<�0����=�;��54��_��`=�#C>X)�Kx<;)��nY��,�*lM��>�֫�@�<'%Y�P�.��O��J�o	z�i��U���(��H��YVB�'��- w��{�x׺�BF5�u�7�q��zJ���٬0��ʹ|��yB�c��!|����}����\׺���O�~^�:�����F�PZ%*�'����W��߹��HTۂ��d����nۮ+r��&�����Ҷf�FZY�/�]��]���Q���:���ݾ\굔���x���� X0���׀�wJ���Bv�F52���'��)2ܙ�B�or���S�B?���L��?�{>��ڣїJ��`��9-���~�n�c+�������՟����>�u�b���e�T Wڲ]mr�w�/�(�zI�]z�d-=�rb�
^������M}E�<o�k�Y���Ռ��ݫ@����<�d�R�)�Y�_Ź�3�Q�NckRN�Ӣ��H^�%���{�=3Hm�������W�U����6�\��|y��@�U�r����� ���=zVKU��L����WJ�q^~�ʜ��D,:43GE.�\�5��
�w�J_�s��. ��fqí��.=W7�Uηވp 	[��K���9gïܲ��t]��H�����Sڧ�En)T�5�Y���[�|1կ/ov�߹�=蒛.6`�ߪ��N�%Tu�y+iU�C۝��~���U���Ȧ��x��)\��վO�M�F�,w�g˝-U�E�|��a�ޝs#9)v���H�/f�>L������[{��֢����O�P����z
��|'�~5O���|��x`g�bDV��A�o��|��s��K^F�-JgG��W�sʀ�4e��}�J�PzJ����q�R�=��g�T�m�h�>�lv
\:��W|^]�_��$0���h��^w��G��S�q�YСC*͎fԪ.S����ssގ��J��]�<o��JyZ>*�S9��zi��k�ll�j�����n:b�:�8~�����5<���(\~Mrt�x��繞�LW��~��
,u�F��U%��R��[��n3�<�=O�^{O���j�{�� �o��.��>yx_�Ϲ�LO��|��HR�K�.��=2�{)��Ϯ�j�®��~	�U��:�.{6Uz�ʎn���*ówf߀��)]z��<��G0W$i���f{&�6� �Η�)�=�]�̼���8�U�w��Z���ה�m��;�n���bJI�	�˩�\�E>�'[�*���V�nl�x[Q�8��4��'��X��U�8�_�/��A��8889�)=�[���_U�Y�����ߍ̕�[�
f/�S�P����]ސ��B��I�ׇr|���={�R�}ˆz�_�:jr.���$�J*-S�j�J��{A���H�yZ� ��|n]گ��
J�鯾.��3���]2�vb	ªa�䫖��uf�f�:4=���n�k�ױ���%`� X��ҫ�0[��tv���SI'E�|�%������6 ZGZ�+:���8��"����r��W7=��|�g3���roق���X�R�4x_w�'�͚{FYt&}��'0��#��B�X���[y���kD�?vO��]9�(ֶ����Ok�N*i�j�bA�|�:�\*q��W�X[���!���]|ğoW[ڋ�k�]ǲM����|�t@�fŎh�d�ұ�nL�T�%X�e��u)�<����1U�]Sf��2F%*:���U{�k����iڂ�_�
������|XÙ]()���3;�٧g����~�󩜿\2py�pT�xA��1�<k{:�$nF��[�<����e[� m�x+��K7��)ަ�	O-���������2�:�T�g���=��  #D�`W��
Ԥ���%�<����`��}�*P��P���:+ ,�^�O��'ٹ��J�z��J��q�-���巏�������8�L�/3����T(ׂ������2���.�!R���ە�D{�����Q�Q�v��W����f�w5�Lj�v��4����5�'�S���-T�}��"4��c�V5S^6�f]r���j��q!�j}P��`�T��U�5YB��Z�zR\)2���=�rZ�g�ه���"��Ѫ��^
���/*|emg1pu�1�ꡧI,ś'E�V��M�-�=l�7��+9^u�QCj���I�	�)j�5�(�^��"*��A%�M~�����\��T̊\j.�CDY��9���^���_l���ALS�-��-h"x��Z��Į*y*�A�/:�&��e��}yi��W��;b��ǅf�k\6V�=�~H�l��۾���G�C�d���ТU�
݊�x�O�sh�m�Ip���p����0ٺ {E�:�
xp���\�6��IJ��s�7׍���2�L�z���ou�t*�(�Y�C��%ի�.�<(���˿<WX�SA��N�W����@��}2Ts����>XN��T���׽0��iKP�6@���|�z�Ʒ��x���D{�'� �0�ٸ�����L�r��O�۟}$���Z�&�B�3�����0_�h˪�s��C����}��x�F~���#�v{�1̮������!���7����DR�s��i�S���d�G��31C���3.�z���k"w�}��3n��"h��Z�-���+��z}��P���{޶�=ز�%p���C4�xthth�^�\��z&Md�Ϯ���{	7��.���*s����=�Dq �I��h�XYs����~���g�Q�+�K������]����-M��x��ɖ��^_�U���
�l]:�qp
W)䭥B���)�_��7������4�ǣ��,�_*%W>�����{������8��j��W-!����<q�L����9��3W�w&0��.យS�H��Lw�����*��ej�iÓ�{�7kw�y��g�}S.`����I��ʼ�hT�0���
�����6zT�Wq֢b�;c�+��Ҫ�V�����}�H�5c�]��u὿R�,ڸ�e���u�8r]N~}F��Ud7�_uZ;%��'�;� ��h��Đ3�N�O9�VV^�����V,J.Z���ݠ�W��^���[�y���V�Y6�kj7ϧ9��H�f=
]L=�c��+�̙�4��}㫟������V(�s�c�ʋ<Z4=�P{����ߟ����������3ԭ�8 Q�"�~����~_L��J�����^
��>�!a���.��jk�!^�ú\�:��YY��zf��v��ʩ}5U�7� /�a�cx��R�U�����`[��RN��^�ksʧ�u~T��m���d�0t�R*/��ON>����3��鞥:�m����T;�F�O)��t����DJW��W��i���`+��c�S>�bYC���$tsK�
�4�E�	M����xh`�U�}z*~F�����
��KG�\��R).z��ۺ4F�Qs0�2]���*�;��x�ACǯʬ�ｋ1�ve�＠&�x F<��� )�4`���r\�P�MD���0�ݫ{i�R'.�6.����!F��W��M��3:���j)}��Bx9�Xږ��n�Vn�4���{�e�ߩK�`ǒ����XJ��s�qO��#q�������-8 �<|MA��� `���p#�FZ:��F���3����K;4��ſ[�R�Ł�ڏ|��jJ�������w����#?.(?~*�4��)۽���]����NQs6C�_l��z)4�1Sǟ�j�bA�|�n���:����n���Ԕy߾q���ܾ�@�W+�]�ł� �`^�!���e��X>���hƠ`���z��ʽ�[��g�򞇐��Ԃ�sN�*GUhd�,:��Ã���Mhڤǝ){�YׂA�PJ�u�dB޸��^�+�5����$ z��[
���ɗr�Ż'�d�m,��S��S��,���t�̓*C�#=1���E�L:�n��R��ַ�M˖�f�|Lw��:Y'S5{������e��!vv����I��bئ�s,�{k��`��w|�G����^E쫲ǮVNq��ޓ�;�Q\��=g��G[o.ł�iAAр�{{���8�s ܀Xf�?0�R�:ei�D�rV�c#-��a���gR�L8�m�V��I�p�ܼϥ��t"J��Y�0nP��w����+bM����5�eC�m����|6�}��k"�j�>{�Ȗ6�!��f\���=/�a�%.�aTq��[%��h�l���7u���[�N�a_�Bkpv�9�\��J|�����7WZn;�RF�y{zn	K�Sw/��M����.�)��(T�H�\4�]����\��y����������0��)j
Z옪�m�k���� ������b�T�9��<�8���Wh��e0�8�Mv�i�\�-꺖=@��̝W�k��M��e��X�Q(�YL.�5��X�N/��0z�z�����7�Y��M0            ��(#s�R�6cʹ��U��p���&O⥐�p{����+�w�4��y%�f!���jE0���)�rk��*uZwJ���̮ɪ�L�5�-�>���U2�eh��<���,��!�6f�2�T���w�	�)^��{���Y�ͭ��,V ���Uܕ��ʃONޫ�NU�O]��eah�����!Dqf-�-��V�]@��T��|^.g(5aU�V؛��,��[0��ݨ,�9Djxn��P\��gYٶ��js�!�v'�0�����a�u�4f:�!ڵ�s��i��V�'N4%Mv�N��1S�*�l�@����AV�������I��W���ba@�i4J��}�\���n�\ŷ|{�aÄ���#�ڿ�!���]r�r���r��,�i�v�4��U�1��e�D�wQ�f�Lһ9��1)�e"�o
�7.��   ��1bfdQ��F�R�Jb������RQTUWXR��)�)��UU�YL�JAi��2R,�)PR,���XIve���h+7����`Rݕj��.]��RF�)��נ�H(�,F���*5��4--Uj�1z#jR�)QF���(d��g^��v�;X�gl�(�^�Ĺ��vL�b���t����^^�Y1�q��J�?�ރ5�7s��i#��
���k���Q>%a�1�3w$�o�����i�[�@U��ht+�'��3fӫ:;<����ۺ�j����.�{Ne����?�N�y���"4?��
M.*���׍��7��ߕ�1����ko2�wu/��о�0j��ËV»e�w����}��2���P�����4���Eƣ���f�ۓ�|�Uq�A���
�5�BE��B΂�J�ր�GuUME���wh9���
gŸ�R���ꈽ~%MI�:Q.b�\ͯY+¯�+F��A�J���R���s1��GR�m����"��S�}'�/�>����=�#���ì�@�
VC�cj�V-�l��Y7��s;A��6�/�+�T�8=e������hU�LVZ�1Xc�{�h1y��lwt�U7mXꆟ�f�u����h�cF�yJ��T{��e|��Z4�6�ϐ��lZ̃-Vi���4t��:tN:Z�7
|�C��U
o0a�1����e���Ryp:5^L){i���2��bDey4�q]�ŕ3{D�WH���>E����^èV[�s���6_���M�?:S���w]s9��m�O�9S��A
��r-����X�������|2�`�E�|@�>�~�����s�0��]��5���[h<�Bã@���j��Dɬ���h�G[s�}:�f䦎��FP���z!� '������6$�i��)q��-\�v����RŢ���(�@Vh `�ʀ�fx�5oww������,���W��(R��ßشsJ�-][R��+Dȧ�Ԍ�|�W����o�UNɂ&�M��zfR�c��������4z�"*�F5h��H`������������`�[�W��y�
�hvO��ۤ��
	��7o�nZ�`��� R�U�d��M�bѕ��3sh����$�nNz*��p�����(t��G.5j+�3y���Ww���t������[Lҿ*ۭV�@�zR��j��黾|�����	���j�(�Y�n�&����|!�q7<���+�������P��O+G�G�8T%�[���r���ޙ��
Z���i!�U��{�����J}WyoE#�͡uO�&aL;��;:E���yTظl���n�+�z����
��Y5�K�_p�7�:�	�m���[�ll�/��������>	8X�ˇ�U��+�8��f��B����]f�r!��ʲ5�E�q�zM�1|����!�*�^�^��-�~g6�u��?u}y�=g;�S�f���A��8�8:��DV���{��M�|s�]võ�_�(|���ãP�_m�"�QJu�׉9Ef*v����G8K��;����S�W
�m�y`SBW �� M9��3�X��y0�tD�E�G�ǲ�@F���V��A��-����ep���n����?x�=�a�5~:N���<��d��<<,`A"���$���|�ijǣl�*�Q6�g�n��^&�_X�WD��8t]el̏�~5���~96�Ѳ�72�ꎳ-q�vhxߍزq���NH@!�5���4;��-�Z:;uC<k6W��5w]���l��4�������0;�O��֍8�y����7��ylL@�ޯ�xR�^���*��܌5{FY���6�˿w�?����O	��::�@�5�։Z`����=����-�26��,�4
>Y�_���j�}�_-��¦e5��2^�n��7���bY�:,�\h�U������۸J��;g����Լv���P^�"j89�pT�x:�GP�0yW�q�6���5��ܞ��6�*c��9�N��a�v@�9�Ζ�j�ڷ{�8��N1��-q�n�n��͒����0����<R�`���ޱS�vZ�5o�T!��I��u�)�ob���w*k@Jg�VE�f��H=�Ǜ�2��l�\�dzao\z1[�{T�;���f������z���=��q$@x����^%Z��,7ٮ�W:��'}�>-�Wy�El�yS.�h��"*.�-���巏������C�����}2�ު#���{��+F|+��
�b���|&B�R�\z�^�c�b��Z������n}�1h���K�ht+�'��6�����D�j�ٳ;3�]/�:i��>5�oy��$h�傑<2�Ս���-����eU�C�:-��i�`���f`S���]-X=��K�g��x8���d�_�X��@���� r�T����M�����Y����2Ϫ��
B�g�f�P���*�:�/�i����/s��RA��F6Q�nU�Ëq�]��T-�,/2�s{���W(�C�ޣ�3p�:3 ��I�+%\�;�ms��dq�R�qS���Z���I}?}\^��ꎈ���r�x���:6��?��>�����+���<��B����.H��Z����`�SQu�K@U��
���[x�A�㷔��{��H�� {N	��;^��(�����Ɯ��%�mC����;I�j��t���eq�[��ԃ�[,�ٽ��H��k����=R֊s��
����;�Vx�ꂔ��By�+�~�-�^|�j2JW�Z)�;Z ����5`��q�VU7�]�i��1��Õ?���z��.Ig}�$�c�>*7�Ш���=��&�a������y��X:�<o������V�Q��˷��w����ʭ��YC+5�����Up��\�\�EX��6=�u*u��#�]'Ns�r�k��hh �X4�>��جy^��ޱ,�Q&{Ŕj��Z��ͺq��Uٞ8�ol$Y0s�W��,N:���+�hYɢ�U��3�lv=ys1��4�MP�ʂƧ�ms��R�|_ꯂR�v������f"*�r�È��:(i��@U� x<�ի�{}�b�/7���Ⴅ�Sʼ+��+hp�:;���,+i������p�)�z.�S�{�M�o����W�
_4-��Չ�í����n�X��0�+}X�Dѫ��8:>uu�sʀU���M�����I^{���C¬ pu��T7�A�PC��WLѥ~u��V�f=��������lԳ^�/��L�h:�D!T�GUyז�G�j����Ej��Ѷح!Uל�{3]f��I�Q���{}�����f�w�E<Y��(��C����{]b{:Aq
o�\��\2��ڡ2�U�;�G���E��b�YƐ����O���rv��p��+�7�\8��Ȫ�1m\_�7�8������G�b��N��|A�w[Kk�$�O+�Z�@d�v޺��@!����wzs'�+�S,�el7S����mL��"���B��1�����k1IDr.,��� �%$�V��a���
�;�@�E�
���M(��'���w�o��=\�iq
��zh�H�E�+x����eE#�T�(3�T�e"!�N�>�ʨwi��86# ��w��v{}t�ZЙ��p�~�#��NTá]2�к6���������f
�X����ר}�ý�IS�swP��{�A����y�2���3)*�.���O�پ?A��+J�۲_��!z�`�5W���`�o�ժ��\|��6��)=ٝ�c)^�4�U��0�BY�_<N�n:ҽs=��½�tP��<8U�Ծwqq���1\ʛ����x�mK�;3���Ly�k(Hk�t>�y�����*;��4�{���~8 #�c����Y�<%u�L��A�`�	]y���{�9�#V񪹑rY��B�⎇vlN�	���Rb�ѭ%5��k�7���%����\q;:���G��9���"�߯����3"�����jV�X��ɘ�k���̿�)�~�s��U�h�MX��]EX���М�����fL�s�*�bǫܬ;�.�C��^4+R��]Qc	�7�ŲON2�G�靫��j�Dŀ5���Bx�?s���m]߆����zrc�5����t�P�R���`���e���71`Z�k'1�$���R�+��ގ�]Qq�o]����ӟUL��s�J3r}�m��mJ��H�����F���}x�W�&�T=�3�����+�&��"��ee��\Gfڝ�?���γ�h�C�j�[ƅ�"�`�B�hU�U��ץ��t��85�з�^�y���P���
� :+�;��.��u~�����y����� a�Ѷ�@�Bu{e�G ���n��X�ܬ����vm�rM��C`)ׄ$��|��+fB:�p���B��k��q�wAWWkȘq����W�I�['Ѥ%���t�5�)f���#C&�t_�Ӈ/Ooz���g���J�Z&Ʊa�j�H>5r
�'�����f|0f�\�\�F������v=o<t�M���p�g���#�oS?p>5���Ƽ4	)�it]��f��@�o�����`p����*��h"ٯ�&8q���}��pj�����T9�X�$v���6΅T�u�b�_��{��osUc�i��񾵣�5CP�<T��6�jg�>����j�B��L�U|�1W����{��|�ث;Q/����T=�����)��&�R��X��n���~#����kСQ=������Z)i)���r�*�Fi�Ϩ��y�V���Ҁ�[��+dC^ݳvk��ځm�a:��ө�����7���h�=��P��1��n)/�������Cl��؃�����Z�*�,8N�!�K�U�lR7K����d�bX6�="¢�]���:���h�s�����zp���VS��f��̣'�y�)��S�Ke���WZNt۴�'���1�]�C{)dx��O9oL���m)Tf@&#�t��O�&7�Hb&.�t�kz޾���C\�����A2�=4����<���!���9�G#�S1d�� �+���Q�*����l�oh1���V�'��x4D�O��ʊ.'s#gsV�W� 7/bvAI��2R�6<��h�7�F�5��v�:֧Z�:q��y�r^!ա��.�(V��"�bC�.;��uuZ��rB��LK�R���V��!�n�6Łh�_U��D�ْ��q�6���%�٧ q-�؂,�e�TY�<\]'ֳ��O��6���@             �f�G��`����Kt��l�PPa�Co�9|l�6J-��]խw;�0(Z���Y��V�w-/j}O��*�*rp�eȶ*Ҥ{�:���J�цL�Y�,��FF���v��F� y�����*b�V������&��#1*�-+f�]�&�xڮz2�_s�B>1���.�ܫW;!r�.�z��%�Lo��b*��40�ذ��T�=	���$�~8e�d�)�;��� �ӯ���$�ϊ�v�k8���s2�f;t���Ņn\+B�F�� ��.Kx���ro,�2ס[!�7�i��]N����;n1a`p�SN��@U�Zf��gj4��zμ}��ZF�h(���;||����W��-9 ���4�su���﷞��Zsi��h�; q�r�m�L���C��5��L+C���ݲ��}+�'o|O�2�ڀ  ;��Ī�4���,�)3b���]��d��I)�(��H���^��X�Pr��x�/�
H��U�����M��Z�ZE��UH�U�R�@7�L��ؤ�URQJ��R���P���ښE��M R�X����-hSLU��TřJ�JQ����R*2��,sRT���ܤ,��Z�B*
S)JՉdEj������V�N�;8��ow����S{5��X6�޶��Ϻ<ҳ~�R�.�?�}7�����Lt��F˟��9�OǇ��ƶ�8Ci�g��5����W�v��ʕ���]wwF������b��j����e�~��T񛪕e���D*�X���{h'2=���әX-m�xV���rr�R���PU��f�A֐ �87/��}����j{��։jͻ��]
�b�BبuR�����d����&,P�5/�Z)�Ǫ��p�R���tu<������Օb�^� u�v�xEkE���߉���S}u���6f�\ʍ�������^x�D��.����OJ���NT����ݻ37�P���Ь � 8ezg�
ˌ]�b[����va����2ﹶl��5Y1��4�&ʙ��E��$p�L�������By�a��d�V�qR��W9^e�n	�Ŕ�hҕ{�#Y� ʕD%����}��wawE�!`��N�fT�j$Mn���h�sl�6tPfD��#P=�NO�}���9�y���k�ǯʢ�[B����鮆�L8%�kT�r(9&����{�o4e��>V�bA���/�����g��4ͷ�A(�y[��q38�K�3�ل+�Jem��o���L��Ȭ�A�߿>�:�5���&�W�ԡ�H^"�bi�$�w�HJ�h�}g<7V�+�X/�x;�)`uq������yUܿ1�YO��ʬ���wwvU�f���}q�=Xv.�܅1����4\�.����n��;M/eK^>̯!��
�0��f����,���R��#l����xT��)���^�b�&8��u�J�z�}dP��^'�������+B�Ã�#FP��N���k�Qxhc�k|M	Zla5�nx*_?#f��v~�Tma�g������z�Y�+�F%kj���ʲ7Q�Ia�uC"�Z���09�L>�[�3Y�%��\���&��-�}�nW-a����Һf�#�1��W��=��e�C-�
w��3�TSۺwF�t��76�,�n�nk@;+oƱ�ĳ�Udӯ��k��1kA�d
A/�jDZ�v�Is�����ء��1�$�Ɓ�*���L�T�������������	�dܹr�W>�3���
U溃�<�ʉ�Ճ���Wlo��XEzP�>Ϙ����g\u�r��u1ڪ]f˰�G�SMg��*�됚�����I�T��5��-�n	��$b.Z�1�����ϣ_W�'�b�NUzE^�t�rrN��կMm��S��t�����Ҽ���p`ʦ�a�[����4a��EOI�}r�^ܿU��qz	�k�R���J�]�._v�n��A�j����X89�{%V᫧���èR:s�՗q>�M��z�X.�~��}�{[�oج�A�o1��MO��m��upջz����d͛5j��a��;��X8e�sn��Y�,����D{��:J�R��z�l٘�|D5��c��-��fʂ�q�l�!���ޤ��7��
���[U7.�@D�~B�������S��a�N�4_">��Q���������R���2L������&
�pi�KH ��X>��O��pg�i˳;��⛧&����۟u\��+l�NeۀZ�@��J�K��?@.];HኽVx+>�T�H��
�ì
	u�4�s�u��ԭxa?DS:>��:��T��ES$u�"�zg0[���ۼЬ�d�%����8P?U�)2�����9��S��t��~>`�u"0�'Fδ�*��M(*f��iH���/��ww���h�`�5�+�n�:�	i�Mx+:��*��Ť�
��E�7�!4���˲��&�b������n�*�ᬛN���p�]���g��^'H����AG��2���e��G&eJI-��F���|%�1���\l���)��}�HVj}ʔ5	��tuX(v�}�F�]���+����g��������;��1��-v�d���n�����SŢ�:�������^�Eh�L���ea��G�Mz\�L�o�6<�f��d��G��r�+�~ʵ��fW�篋|k�
��V8}��1�����o�N�wHR���+�G%��s������x[�k�E<�;�(���s�#�;ҲZ�G����3,�-��P�Jz�:ܿF��v\���O���&�˳�۞u�h��ވh �"����oC,w�*�h�Սxze��k�:��*T��D�آOvcZ��|:}���T �%�.ׅ&hB���5��Tź$�ɩ��^J�ʾ�A^��[���s]�c�4���8��Zȳ˩�����ʹ���;Iv��@}��^^��牠e�Z;���j���a�;E�#R�t�婢�:y�(nF�R�V��Q���>iW��oD��f�/>�w��ܳw7���Bi�U�"�ƭ�.������<d>��ÑI�f���CT9պ�:�����u�8�t��\w�WL��-�������\�~��P�J�ʗ��J�� }�f�Ct�t*�"l<� �{��Zڞ�^	�a՚��X��Tõt����6��UϦ>���~�E�o�5���S(`�>f�		�QU���]*b�9���)+)�����6��B੘��jz)�������B/��9ʩ���{�_k��R���V�W���<�[�&y��������)�x)|\�}A`�to��s'�K�:�疤�ѺXc��ݎ��f�|������ tX_Tj�{�U�s-�ԯ:/=��е���ׁU�5L�P��I!evx �mi��/y��5��r�������X�\�Ɔܢ!��cu���9��^kf`d���G������fY��@����/m�w
�^�qpo�]�6�݅?zn ����W���R�~Tr_������������֟�F���u��P!��F �,��i���~N+��w"�#^ヅ{Ʒ{[�h�e46�ו���A����J��x��Pjì(y�����Xh��搫��;��3 8���?vw�g�
��R��}�q���ઁ0� S�g��V�ga����ͩ����T�W5c���0�%V4�[���#�}׹����V��̡pװ�2�
�=Bi���do_n���y�C^���_h�^:.���VjԈ�j��>�%�d�C;>���+�UF�Z)WB���ʌU�^�Q�%��);��'�Y`.w#н\��ů��З��I�1ǴE��b��	P��1�8v�1K�u(̑pWk4J�7Ӊ�����'=�cD��8�icE��ÿau'D%���GH��dv��V.9�ʘ��8۸�-����5J��� D�2kkq;]ӊ��[�gt�:=�Ѓ°U�^>�+��UGR���[U�og	�P�{��|25E .�XT8<���U�jޯ_��?'R[��T��7�.�x"6��{��*^>�-�/��O|j/;�7ɾ�\ul�G,Ͻ*c��n*���r����T�v��)��5^�,UZԅޢ°b�F�.�[1{�Ʉ�F����'m���u�|>�˃��Ţ�:�Z:���?���v'+U�z#���U��_�֬_!Nrsn��n=�Wnׁ�yI5+��[5��ZmS�����- V��B��/۬��y�Ħshf]{e�0ӈ�j�#�����9w�)ҲY��{8���^���s����Aiݭ�*vڱ��3V��Q�ur�[y0�j����ihu)��﾿^sc}'�cbL�+d'�ϑL肸���PpѴ8w��^�1{���s�wk�e$�.�u���zs����W��(Z�^	�ۢ;�oڮ'!n��]�wN
Ɏ�hZn��Y�>�|�Yj{u���K�3�q�G���׈�x<5�i�F�#��^4y�~��:��>~�ʕ�������wb���m��7q�T��e�;����#w}#�졂Z`ܵD+z�V��뢄��ĳ����' ��{ɿO����� �.�mX�ث0�E^��p_�CިI�Ng�)Xg�Sy>������~&/��Or�ʼ4,���oz<��L�zu��۩�WS����fӯ%�͋��i��ș�of����2�R�mͤ���N�{W:���їj�Opw�w���ëg>�����m���[so��ёq-v����ܷ���nr��z����
Ef땽���e�3,m�Ձ�6�ʏY��e
�'�����G<�%�L.��Ҷ^_��`hSGw/i<��+�LITM���jm׋�W^֬��64vߝu#�>�4WJ�腶s����%<����\%����,���߮��N<��wN��L��'=��Ƽ���A���|*١�^�\.��ޗR�_f��n���DfƓX0�*�Q��'l��n�"�����P�=\�z4�w��s$|�8���"�ƈ�	7d��L�=�9��H��mP	��P�<*P�5�U3�$��ڬ�>z�2�q��=�y��j�k�q�W���G#=�8L�~���g�ON��p�u�YԢaJ+g�3�Q>��ff��fT8�X�������Tz(`��+v� �EV+j��َ��>�*Sx�	��[?(�y7P�h�lՓ+We6y�v/w5�Wr���]>�J�oWE�
T��	���k�7�)!|��N��ϊ�����6�m[��ݨ3+�¶��f�6]�@�=�(0܉���n
Z͢�:�E��W5������dS+r+W��T`��}�Lsz=&���H��zd�1��q�,�t9 ��ɤ�W����R�KbQ��un;�4�[�� (�i����:Կ��vZ��%n�xX�&��W'Ҹ����L���C#_Z��P�TO_#W�TI���9���v����u٨'�jSz[c��K��0?���Q�wh�k^���}���8�6-T��ܤӉ��n�S�^�L����6>i�}9w.
���&`s����y�z�WnR��I�G.mQ\�w1�J�$��n�Z<��B�ekGmڝMLw��Db��:�bh���9+�̀.����fWv8�|��!.�y����:�8Y��Ka�bt*R��'#�         	$�H	"��,,�eN Ν�v���̐��7b�q�@�x�StA�Ճ>4%Ydi,��"q,LbYׇ����7�w��|*Ь�`e\Gj�e.|%�o t;�bvi��1�ecF�Tt2rݻJ�����w��ve9�3p��!$2�r6��$��|�YR��:����V���\��[u������fY�6ƴA�CI��Su�v��z7P�m���p��2�
=��%9ƻ���{tdu��Ť��CXv���5ݦ�@!]�k]��f�Ⱥt*����X[�B����s����+�7i[�h��\���1b` cū=%��n+ڗ���ȑV���VWP�N,E#��G��E�2�"A������h/�fQ������&��Տ��u�oV1�7c����P�4����G�5��}��;�2�q��h���P�3�y� $ �����D"����R�V1cƞ�0oR��R�V
*Ū�Z���TX���+j)i����X�X���,Ң�-3�)��*JX�M����F��TU
L�1V�J�0�Ei��R("���QX�ILP�����5T"0X�(J�L$�ER#"�b��T�PDX(��X�DQAb��
�8�A�K�B�X�UQQ#0�X�IL5FTs�罽U��Zͬ���`Y:��%���I�T����R�/=�3��T\$��Q�Gՙ��C��Ih��T���LK?�:�
�9h��v�:מ/6��|̯�z�g�-�� �]����4��@��5�¼�oԫm��l�o\�F�پ|%o/g�o�
Tw����|;��ܽ9^~H�&��g�!V8&s��O|�L�UPT��4B@W�>(-Oy[�����+��vz��W�������@S���U���uU�'����F���>��X=g���x~T����u�{I�����􋏰ד;B�
"4P��Y垵a#��&���s\�ޜ�*nja�[�}(��Y���]RU�\�T�M�}i����}���|��C������+EX�t_�����ѿ$��������u/TVuX��q���@��k��0/�k� S�R��C���!���k+@�)�����0�����@��E'0�"�%����
����j٭�n�yC]ݓ�.��Cϴ7�b��f�r����{����̞��¦L�����J�B���X���+Q�]+w܌����L�|Oɿ�x|0?D���-UZ�^�"w.���{���Dȥ.���y{P�<#��4E?�X�/���XÚ����oV̸�\9�Y-��ئ��WwG�k��*��]yI�W�t��xkէ½���+��� ���u�6���7_o���Lz�>�*�*U<���x{Ʃ\L{5 ޓ������Y���x:�P��`�����=[q'&v�}=V��^����,]����t�k�89��*�[���F�Vb����0�j���~#��`SEC�0jVS�c3^b���֝�G�hc��|�
���|MLu�
}�pwೊ�s�f���7s�˔��2	�]Ր4]��������m���Ρ5�gk�^���H�@R@�Mew�8�̼X��Y*�
�����N�iǨr���rOs�㸯.\`�~�Tu�W���dkB�*ѵ�痒?fwl}���
�X~�|v�A{�*�wJ�R���>įU��RGWs�/k>���0]%~�Z�|�8Ԝ۷xc�A)&p^��t33�n��vR#�}g��	R�h��,�=�S�+�{=�u~�<��P�mr�Ғ����x=$^Ta��Z��o�ۛ�XB w���ԅ{h�$Xs~oE1��uC���y�k�nqo��:)ڻ��.�7�,�;j�� h��I���Eu�hKU5�_�s{�N4Q�@/��p����Ga-&��}�y�<�{���VlV8��}^4�����hu�*��>Kr��O�{�(߆��]�[�߭��1�`w�!46%�<V��þ�.��t��Ew�W��R+j
�V!�㳓��c�=s�޸{�o�zƱ�f�;�s�^�
���Yօ	��pɍX"�*��\����{��~�g���Q:+�
?�b���<<*���S�V<]ה���Q�ܜ��=WF�mo��[��Т	5~u��������x���+�\�t)%�}:��jA.`�٨ݢ~Sr.�o������v�[gmJ�d��+�W��B%�Nv��v��K;V(��b,�S�?��]~�\�����zVKL�t��k"Hfj"7�f����orU �b�_�oD�&���Ώ?�=)��>�S���%�ϳpCoee�*ff�n�]�@nSV<�鈊��\�3N�,s�¸���bJ�?}��72�e�ǽ��
T�W�UyѮeu!���o����`�\�y�U�j�t�6ϝ��9��S�����<�5�㙕���d�U�>
���#FEm�me#We��b�e�E{�^���Tv֕�`��b�l�E���I\�9�F`��L`m�׮�&���v[��nH�qnZ�Y��´kq��Yut^��Wm����f�������7}�S��@h�9p�Z��è��U��y���&jW6�w<�!^^U�3P1S�R�T��|@t+��G�q�;V�kp��O�E:ۇ�n=��قWF^I�q�֢aKaY.���zk�תyZ<4W˲�ЙC��f�]ϫ�&bIf��}��oJ�mz }�.�Cx]Q�AQ�3���5��.7/��g����ꎗ񶥔Ký�ժ2ɭ����SU��}��Ez��K~��9��a?MWYA�w�WF�q����Q���[��rU�-_V����~fUu�'5Z��Cy�����o���ɮU�t�X����Z���n���;�):�y�j�vޱ'�K��UZ<M�BǼh�
�u`��������K�S���Zp������)���hv�gL�{;tl�
<�������Onc}�Aޡ���+;���5�r���tSiU��gI�s �m�23���w�S���ǣi
x�к�T(Q����O ��z���T;/��#���=��F����4�����],����(����!G�y�x#u���qC���/�ך�cEXE��D�7��xjL�OB�T�&$�u�Ū��j�:�}6�d����X< �T��:��?���V�*��ǅ`|�q�%=��C+Շ�� h�~L։H�`~��+��h*�
�2/!��s|ST=P�*�TUo�+56����Z_��-��u��OO5=�W�t��*C��u���,>c��F�w<�+��gx&�V�_�������l��~G#^qݺ}�>�����=��[�Qʨ\����X$ڧȺ�^��Y��f+|h�T���13���R�P�)�r6�N�3�si��r8�1HP�X"��LTz�@L8�	��;#��{"��<����*����~o�7�o��+���E�^��;e^K�P�T<b��3���&���Wq�O��>Ez�ƛ{��EqU�C<�wONr��"]��l���b�k�9��Ƶ�ӻ��}�[]��Ρ3o�u���|R����������now�϶�i�����H�??�����g��y����qOzzU4=��1��&'����ä��^K<��xgX��޲�B^�����YF��;)'�y��bɚ�{;������k�~T��pG<&{�QQ��Tq��h����x����䜇�RH����@������]�H��W�w����z"U�OWo��ї��Yq)�a'�p����d�H��0��f���/�^���2�Wm�;��*{M�)��F��w��/�Zӑ��W����PE
p7q�z-g�uUns�8w��{�1Eh��^�gv�V<���hKɼ�}f;�+��N�ck/}Ŧ�K��J��N�8f��������p�ˢ��3�{#�9���:�|���i_"���y9���o�9�F��i��i��V�B�O�b{7��{�[6�,�aN;�s�.n:4���]^�4���C�@��k���FB�������;l�#����������揭z���זU�� �|8�_Dլ�#�^����P����*�LCCewoNV��U��Τ�}~i������Z�/��H�˚Gsf�7h���%㧌�?y_kM�����F���J������dT�Z#3���3�����S��� }�[౜���k��A����_��Ŀ��9�c*{�u�yз&�w{�S�kS��+9��J�?Z6�4qU�ȣ��ٝ"~;ޮٛ�6PU�~t��rT������1ď�YZ��틴�ee(�y�H��%w/\����g^vt?ToF��/jZ�s#��7�S�~��x��q13���],�kɶf��O�$��q���J���G�k���������a������S@�v�����D���C^ih��^��ůp͖|z�:�hB��j�Y� �����G���}]n���;Fc���[�Ӛz� �U�:-��dT�7��-��j,�9�q)ś���'Q��W���&��x����P�~����U��ފԺ��H�^�H����w7��}ȌͥYc~z����8�������������$�og��9<�]�Y��Z��	�m{L����'Ȯk��iv*Ή�ۈ�I��k��|N�S]��7��=IfPc�"p�vb���s��rX�{z`�φ��W*=�'/��E����=���V���Uͨ��7�Rc�L�4{b^���^��_�rn'����n��x�/�(����A�s�-f�V1�{�.�՛9߼-���e�wi�7c=ʵ[��ں�GN���'\�0���i���ކv�+�om̥��W��<�ZWd��(�B�����oy��aB��ah,vd�*�7�Yui�%r�e�\W+�����N��Шp�J�G�OoA��$�1^a�:]��t��Y.��M�M��2;�>�7���N��)��z�
���)�8�'ov/��V������ވ����;!+��i1ֶ�v4�X�>!a>ީ.�r���QZ�39x!�4����N��>콽���b�0N�w����*�z��D�֧(�)c��zͲΗ���b38M�-�g��}aKi'��EmR�S��/g9�7�Z��
��-�9v���n�S�У��֒ʕr�J�
��˫��+��4������cTt��GoR���E���:�����+N�tG*��Հm��v����c�r�z�+������
3��-���s��{��6�`�M7��b.�T�H           �iA%�C����)��je�f^��)L�JZ!ᣛ�n˃��v��Y�&�or�4�'��?.�w�/:� ߴ������#J��{nޭI��v�J��=҃DFt__nrT����B+���p��iW;�����|��)J	�X��:��h�|k%&hM���s5�-n	�0N��+����t� ��ċǶ.��˩fA9�8�ʄ��݌��:o(]�V$5u�{N%]i���q*�v�}�O�l�E��!�h��J��sf�1�S�s�]���[c����x�71 [�)�\�u�T��B}��N�S:�3kx�4�٩��3^�5���Ǉ^IA����ZVP����D����݃=���Õ9 \{������wІ<խ�s�\nZVKFWV�,U��\U������j��P�`�jʜj�I;�I��R���$S[k����   .�'ꢙ%�r�J��*���"(��BȢ�ݪ���UL%
�;iX�"����"�Q,Xe
 ��X�b���Ub�(1bE���&U+-A�"�1X��ȰTbŔ��(��((dQDK���EoR�UT�H^�TH�)�ȌX�*��^2 ��0�a�,X�b2("��Fb�DX`R�TE�"2(,�,���*�ұ1��`��U�@o@��p�R��T�"�IB���,EE>���[H�4=X��,��܇��Ś3i�j�ڳ��7��D-ʀ�n=��&��x>p9i��J����|�o��	F���˻}�zr+�Ч�Ǔ{��h�O+�5iec~������R��£@��߼�=;y������EG�^�����}��{��3'bW�<_��8R�9��J�����Y�S���G��'xy�)z�ټ� U���U	ۜ7�}�޷�� Fu8����Ƽ�lUl�g�V��.=���K���Ϥ�9�����yuA��V�~��b����ŉ9��:�`��ꞹ���>+���k9�]������/}&'
��]�R��5Ɩ!J�6���/U��Ј#�����`y/+�Y4Vl4Z�;�;������?v��5m��U΄XS5��Tt�����W�x��M�J�=����?���~����3�C���s��&�0�Sѱ4c���e�8q��+"-n5ns���;>��j�2x�9�g_����]�Am>�׽�Z��{g/$�Љ��h��{ןraꥶs�{,�g��
��	�}@��ХM�Ҙ�F��Q��}浢�/t��m�G;.8�RRd��^���w��Nض��^��cuъ41v\���������FoeA���x�0�|�6D���ѩO{��M�ys���ya�Z�VsV��/2���Q��w��!z�=k������q��Q}�$�'m;/=&�w)�:�e��NѦ��<�.�A�WR��1�h��nh����)͹a�]���5�$��۠6\�ӈ���nX,{{W���*���T����]e���ew5�N�y�a�N�i�����zz����q+��y�1#�6�N�p���oV�ZLv�O��VذKާ>�?W������oL�U�y��{��؏�z0Y�
����o�9��&2����[���3ܸT����>���{:�s������vKr1۾�c��,�לw��$��Ч0!���R�gVFs9%^�z��J����6�p}�㨞ׂ�z�kl��eS>�Rw��Y��ky*{^�VQ�K�	+9���Kٗ4u�ֱ����v��Ցx@��;�Zޥ$G;��u'i�1V�׏'$[�ޏ75�핥��J��%�W��%�3.�h*=��;���A���5/$ne��;{h �:�#��	��\e~�W�ƫ����ݞ���d_I�����C�e�oo�Дy��x�L���mrk��q�yI<k��yk�x��cGOG�s��(q�.6q��b~.QW޵�}���fr�U�-1��N��|uD�C���K��z;s�}�nU�,Գ�+�.p 15~վI��ľ�{G�@pC�=��^��o��z���1R��wb'>�H�+��Ê�~m3/wq���Qت�{~Y	���zJ��P�{�F,�S��/�`~��9���|��W�׸P��Ў-��JdtRw��$��[�vrAtx��۰>�R��16�/�̜�3Nu_c���&�i��'}�d�&�*pra6��*����}��mI�<M���.7*%���ȝ�Q-�l,�_{�	�6Ѵ�h�ԯơ�ݘ�|F�ʼ����_m�W����s7{])��.���k�կ�.᩼:��(Q��Z����~�5^���s;<��t<U����lvҭ9nc�e߲���/r�+��WFRu.y!�wb��":<�,`?c���~�O��S��Ǡj�߼�MK�=g�k��mc�%�j�׵^�`|���wY纼�n��:ћ��gʭ*�\H��үK��`����
��y�S��s]��$�o�����r�*exmۭ'RF�"\k���b��*��+՟�B'3�:��}ݣ&r��ޣZ��㱏�
�ni:��Ja�s�-&��yۻ+B-����WrԎ㽯��R�LN��ٸ�Ǣ�{ڲh�K�򷾩�&?��9LJZ��U|�
���{�S�TK�m=��qbI�;��]���{��kޚ;�\*%�gT�h1F����.h�9��M�Jp}0�%�5{��ǀצ�
�Ǔ�{������~
z�z���[xל�}�w�wޞ+M�'�i�WM×å$�����Ofs��z_9�w�|fz����j�_f�OsF1<��iދx�N�|qej�����*a�)�tg/B�ؒ�k���.w?V7ӗe�oA�坛ƹ�E/�Vb�g���db�����@�n3L�^>܂isD�-�����&k�h��2M�"��:`��cB�:���vjk�^'u�����%�2���d� �с�0o����.��q.�����ý���QQ�cke�?_j�M:�<��dɼ����f��U-��z��{}�O�%�N�U�|�m{M���Ud=͟i��<v�.<-p'��iM⪉��ِ�6��E��̿pſrw<�s�蝚�I�ss6��	�zl��oR��{�ngB�s`^`:�}ɲ9Η<�:���5��y��ٯۯ��1�Cq�1�_)�ژ�����y���x�~ۛev�^���1���F�9o4��*Ƶ$܉� |�`r��Ӻ��{����h��{�����TN�sEq66eo*�	;؞�/6&�����KN#P�L#J����3B]̲���S5C���q�ɴ��&��ޙ7Q�܉`1i
27�ؓ��sv�ۍ6&��muGR�����k��cq��{rM�k>�}���	�Ѷ��G� �Q��_ԟ�dG���:&<��N�1ZN&���W��#�R����պ���4��v�kR+�?��77c):���};S|�^�$�w��u�9ꐚ�Dt�<��	�>��Ӄ��yA���V��RwH<����4���{T��τc�s�tT{]������V�罽��k���e�ދm�9<w�j���[:����>�~����z-����=T�^`}	�q;Uឰ��bC�V5
%>˵���L;ȴ��r
���$yP����w�ɏ$i��B��ᓨ�o*ӡ�ވmI�I"��w�Ơ����Eӟ��^S�D��RM�"�u-�8!ϼ縿�s���9/ޅw��l^΁�d�}�9�'�]�.׌+�|��<}��a*(��7���F����q�^���F�w\��S|������S��򚾜��߻a�����\��+�4�t��˸���s�g_����Q�\Mt%��=�<��9�e�(4w�2��ػ¶]������|���!�
�Ď��x1��
��յi��d���2�.W\��J�+�5�JlM+����|�W��׎
N���N��c��ų��|}"���d��*]���輄t/_���>�wY+iw��d�́M!�ַ�]*�ܗrf��w���\��|T�5,���צ��l�9��=3TRp�?g�.b����P�Tߧ����;*����&+xל�z0�ϓ�U.]��y��!pGk���]�^��追�ě�L+Gy�4��O}���TIΌ�zw]ܸ�[�ݼ�.{��v>�?m��*�� �/6"0�=%I�^��?b^������Nz�ۯW�*��M���^���dk��@�۸J�.�2a�9��5�	��C�BE��G^�k��s=[~	'�۳8�9�<N�ܳ��[뚉3ܸ�pb�z.�>^���)�s���B9Lgc��[�o��>��������]��q����P�P|q��e6.����bK��	���j�G7{y��l��7L�Ʋ2`�'5A;�N���W
�յ�v��	��r����5y.�\����M%�eq����u7�v�-�Go_;o�mv:���]����3�ȃ����Ś��[w�Ȥ�灵-PD�uު�K�ce�yԜ�1��$���4�9|�a�G�b/'�*V�������0�%[n�UJ����X�7�4�9t�(�J�^S�e�
�9u��++�^nrs�gG7G����K�pp�l��sLs�no�����kѬ�s����+i[(�*u�ހS�Ŵ����g�m�3������Z�j7��t)ӽ�k�sx�87Pum���9/��{���d�X�%f�=x�ɭ[�j1���\� ��.�ku�7���͙��IN"ys]Ӊ�D��[Ǧ!���]�W��u�9�tյ`��F��rV�2�Ȭ
�ha�pi�R�^��k.�ྜྷ��lM�>�U܎@            ,�z}w�%��:�0@��[Y�-��n�T르���0�+���w�X��Yy5�sܩ�ź��茩��S�IM��J�i{�a���}��75�
U;�ΰ�e��`��י륖J��ƕ��r��u�J�Ԕ��kݙ��;�Y��
p�ӥ:���R�7� �/8����Z;RX).��cn�2bһ#\�S��=Q�襱w�muA�)î�
��j�ҎV�� �N@+�ξ�c�㴘��̡h-x��_`ϻ�X��YIĦ�ٯhc�Sj�1"���S1�gu�)s�&�9Ջ���zR�N؛�T�n�gu�k����3D�k�[9]���C��Ma��I��a���(H��J!�5<��] 32Գ�y�<nM���Y. ��>ը��z�&J�i������E\�s�}����O �V����   ���
'��>����&b�

(m(H�T`�B�Ғ,�H��j S&
H)��*���d��)�X� �#��)�"�I`��aHB�� �Z����E!�*A`,�C,��)����"�) �J�mj� �i��!vņI,�UF�H��T�).�j�
cz��,�ِ1z�P�� �2I�J�3�˷��V���AfWfCô*8�4�Rfe���쮧��Q�G�a�C���Om��`S���e������Aو�>���P[��{ӽ^`_A�Tj���0��Kr��ڥ�|����0~�8�/^��#�����+���	g{(��0��_��f�v]��¾���f�S��WT�x�̧�]���q(����>���lB���y}���w�~�i���]sǹ��=�����W��9���1�����Oj���2��g������Qۏo�Cه���|�|%�<�����+'K��\��X�ո�oc�.N���5#gl�wMz��7�.q'u<��7��������w�nHg,ʬ�W�����t�s=�^G�T�~��g�O�+���4V��{�&.�Z�����H0u�E:�E����foI���N�t���ΡN�l?&:�ۅ��\ٻ�cru���=��W;�j�bV������w7�k����g*Ⱥ/>�{=��Zg�ܳz��<���	{k;2�\�/���LS��������_�@N�8��;\P_"�A���S���*#�1^;>��ό9a��Afȵ�����^��V{�5�~��2²��C�U�z�ڛ	��k��gܛ��*z���}�k'KGr���!?�r)�P�Z�g�U��^�x�;.ɂ��̾���QhIO���r��/)l��]��g/; ~Z�^��_���Hr��k?_{wg)��u�rl��'*���ю���2�BT���ӗB���Q3����������U\sf�9Ŭ~��%%
�ܦ)���yWݧ^`�Zk�\.�t-S:'���lm��揋�etX����=���i�[�uy^\Ӊe�P�Z�i|@�'����ٛ�f�L��{w�/��F�yy�O��Us��{�ӽ�?R����zom&b�|��������>��W[�םԛ~��y��m�����?o��g_��*/.��-������+^�CL���mo���T�My�,�%�+��{Ƨ����;W4�c�gu-��a�P��߭AK�gscw�_z��k�������n'8'���F�k|�p<�-�눗���b�8�FVG�JQ�U��^ဎ���M�w]�y��]M�ܺݏ��'�RfW}��C�TB���Hv���7�ёv+ݬ<�7��V����q�3R	ˣ��e>U���l[,a��� �ڟ��*=�w�=�0uJ�d���ju���$�{ܛ�׻S�>U�_&$n�e����c�BY�&����ӂ[^.�Hoʘ��	��J��[�ʄ�Z�~����Ւs�ٟ�~��k���p�\�lìܼm���&[����Ʊk���b���Q��n	8�Ѵ��&M�LV>��y��C���(��՘	~s���ys�)W��OoE�u]�k�׆�y y��f煝��LS}*$�FZ�2�H�f�=T#\��+�v>�C~����PV)��Ǩ
RC[Ǳ+��{�x�yJ��H���[��F׽GƉP9��8�bR֬�\
�>[��Z�f�6uJSU*������9Ys �o[��B榅�l.����7��(&䮻
�Vb�R��[d�ۯW=�I��>�Z3jڝ��ŉC��թ�~���Kas��K}�Lpѿ{�G^�j#��s����{�6�x'V��[��);�9.=�g� gW�t����z��^��e't;
��j��oS��?e��=ݹ�rsV�~5ݔ�nH#��f{�zM[��]�η��Tǂ�z�n��dҢ�A�s��������k��E(x2�y��RĆ�%f�
�"���]�-P茟L-.|��d'��&��_z�(�I����O�.?^�y���^�ק���^=��J�[u���Zx�ś�5�s��b�,�^�Wb��g�͔�����i�n&o~�0��]L
��|j�����w���e&����@̓u:�n�^d���Ԭ��-뚷��nd^#[��~�5W�e?!�����=�s��_0�8�=�ow7������u�>�Yq��j2&{m���%�����&}��j���z�/�8K��·��G��%�{|���K�/Q[�)��3����W.�`���Qb�8��������s
�}��s|�g*ȫ��gg�j�W��t�9�I�PRo�ى��/���M�����Wm)�ţ;)�s}Ք��B&2udm�����ex;��x��̌��^��rr�
A�y��w�mOM7ի��Gۜ����Xd�Ї�|zE]՗W0�%�S8��N��,�33bW�8Gc�M�� �)2�8s�0p�@�yj[�-S8b�ȑ[{�jC��7��L�Pe��:�{�����9���U���V!��M/z��r�S݉�d߹D|��w�V>�t(U"�e�mu��/���<������/}����Q	%8��C|�ܡ����ػ]���	��3�)coQ��"*u�*����h{w��t��q�]��|�gy%&���{��"�XzZ�6�]�|M��ᑾճ�=��ꉵj����Ѩ�}~�{�����Q��^i����n�R9֧�Zoj��-/nU�G͂y���#z"S�>+������^��7VN�R���6e,cW�-=�|s�V_q=s��W���*v1���2鄆]'��M��2�Eh�"��ue<u8��ʬ��q7e)zn%�؉��6+zR�e�뗳�km������Q�Z&���� ���KWc�_t��`n"\�z��դ����)�����¯���vz������1�+YZY����Ic���777�w!�G�Jf�SZz��9���1��f�]������w�a��S��s��5߬����v��v���z�5�����L�$6�]\}gy|��=��Mr���go�!��Љ��@�{����9M�G�Oݧ�s+U��l�J�7a6;Uif�U�{Z����k���_G��Q�b�,.���*nkM�@�4��zW�x�1S���QQ�e�E)?v��&�^=�ѝ�(��_��f�-����D�k�]J[]�5�yiYg#L�YW�b�x�U�;�qs����y�B��	��=�ijz�WP���V�9˶�rq.�X4gJ���򕡅f�#Rqdx��e�Nkx���e5��Fne��p̭*�ynF��#L{����jo�9l~4��Ҫ�N~�08�,M���7ؕ���
�yϹ�'���ҍ��b����Ê����K�������~X���W�eOF'��U��=��||3�r����Xf��������])��^�kN��}��P���� ������{6x�*�1�y'��]V�����ň�p`�I�-�>�/fV�M�zG��M�� 9�=c2�����n����vs.�y�&G��V���_:F�}�]���pU���M�{X�1_A-�+y �Y��R�{�V+�c�t��9T�1��~ߪYy���<�^�s�i�OR13�ri�nk�5�Ⱥ��RD�IG���B2cLG�\�� �5�W�t�ɽUM��O�A���G��y(��"kXFK�Vv8�J�Ϸ���fj�3�ֆ5ŗ
�����]\�3�+�/F`}ɫ��g�+Op��~�R��&����μ疰�`"����RyA�R��Y��vW�e?!�M��a��OOE�C��^6�x�7��yۑ��>��.�J}�Y�F����R��lf8
�{�q��[��;��~���y����k�-nH�숵���=罏�T&r�߇��cag�:�u�G1?b����@Ù>�7q6��!�y⋰c�W�1�o:���~��'�>����O�E4��(UO�$B/Vr��$B=��j"H�l0�yʊT��0.X��\-��^B�k�C�\�&2_�u8��R �D��I
��$H,�H�U@O���e1Z*i+4䉤�|�� ����S���1�ZKk�|����!�J�՝Us}-�V\�l=���͆��e)y���:0Qy�J/�ƌ��4�;,g�io6Q39�I��
�`�a��503�$�����8�_��&�}d��0넒!"��@HG������vGG��9#j�A�I�dOZ<�Y��sO�u?i�bu�$�g_�D#C�#�o�Γ�IJPٌ���*�t����
Fr�/ֹ�db�ԏr�W��~a�j�I(ǟ���J�m��sӑL����$��� �>�*v$�y���R��_B%�	!��lKI'��x%K�bmY��k�1���6���'����"H�n�"d�UT�pdq��c���i9��yůJ����jLNc�Q�n����<C�61{NO�Y���׬��7v%KID#)i*k^)�;�#��9��d���1��.��i3#�ط���.�ӮUb��ğy�sh=���d��]�g��3s��I�aԩ(�:=�����ۊh��к��~��DYR֑��HE��"H�}�ԟ)��_U�ZUYj{R��i�SF1bF�!䌛�@����=�ETQI�^]\�IG͢n�Y���EI��b��H��2�����+\*2�4��@����B$-$�eO�KRZ��3����U���e$B5˞�K���#�GL���
�v���I(�8��Ry����Z�������2oE��'	6��W��V�Y=ɯ�G�x�_�9�a��4�>߹i	"��7���[�Ux"�Y�Ez�$�E���˴�%���1��l>�����FټK�#�ݞ�g��FpT�S���)E�z�ŹC� �ݩ���ܤkQ���j����^3MMf�;��7e!$B/�Ԏ�evF}W7[�,U)�̲�ƣv�sl����(ڳ>���F(�)�Gn��T$��IRO)y�.;�#U:k�wy7�^�f�I"�'K�7�&I���:���+"�4�s����^����*�(�;"��9lmDپg?���)�^pf�