BZh91AY&SY�]٩߀`qc���"� ����b_�R��� Q(�                                     � �x �A�  F  `,  �        (   @  P�( � �P o�J�
JT�A*$T�(��Q ��A$�P�*�*�B���$����RR� �R�*��
*�:P  t���RH��@ >���*lB��6
*�D�t��Q��Sv:$n�#u$ZpiYb
w}޵� U |����hziͨ r���
gn�l<�� <���������	V�P��^���`w����wP�h E�� �|R�(*$��)�%R�������z�y������)����Pn��Ǝ@tsc�΅���gxP�#����
   .�T ��	z;��y�U���^{�����{:ձ��-��m� �=� ��u�4y q��   �M�� r"IB%(�O�&z ww@d��x�C���t y�E*�= 9#����=�l(S�yE8 sc�;�  �(;���p�{�=^�2���C �@z{�@{��
z�z�*XA�a� n����ǐ�� � }R  ��P�$�QQ��Tm��6<@;�v�:�<����T=8 Dg������p�ǐ 2*�nzz�x� yڞ �  |�� x}��N� <�{�0��� ���� g��+�� �9݀r2 `  |�P �U �H����aJ�n���@2�݀:2 b�)'m�c�@ �K��8��n H�A�
  {�@ }�>�@n*U. m�@7`:�pG��8��G ,ƀn�uF���P �  ��*R @    O��IR�      4�j����  �  &F6J�4�S(      $�IH��� �4  �� "D�DJ@	����'�Ʉd��i�I�}�������#W�N��������;;�m뿈*��� U�T>��������İTW��?���3���vmS��UQX�RI$�j*����T��EP���ߣ��	�0]��f��]�vj��[�Wf�e���]�]��-vmv�S�LJ`�	LR��1N�BvZ��ٵٮ�e��]��-vU�k��f��]e�`��)�S�	LB�%1
Y�vj��k��f��]��-vY�٫�We�ʻ-vX�	LB��i�i�S�!L[���]��5vk�L���k�We]��-vj��ͮ�]��5vU�k��e��]�1i�S�	LR��1Jb�ͮ�Uٵ�k�[��f�eWf��vZ쫲�ʻ5vZ��٫�̻5vU�ٳ5vj��٫��ͮ�vfZ쫲��]��5vZ��k��ݖ�5vU٫���]�vj쫳Wf���fU�Wf��]�T�B1)��LEJ��)L6��V��kmvZ�[We�i��LQJbԄJb�S��4�BHDV��4�T� �HAQ� �1E)�)�Unʫq-j�	�m�*4�����D�"�0Zݚ�vU[��[��쵩� ���4�� �1)�#L`�0P# ��������� �0 i�)RE)����LDb��� 4��
�1i�LTb T�#R��4���0Ti�#LDZb��	LEZb�S�4�A�"�1U)��LT`!L��"HAA� -0Di�LEb1�Lb�Ԅb��� 5�kvm�vU���emnͤi��LDb����1U)��b*S�"
S���! R���D��֙����]��q-mvV��We]��*��n4�L��1
b�)�S�-+]�]��vZ��٫��ͮ�]��-vT��k��e��]��6�6�5vjgf�e��]��5vj��k��gf�-vj���٫�We��]�eL�ٵ�k�Wf��]��5vZ�e��]��5vj���B�1���T{��0�������z����6��ǝ�	ئ���V�ۼh��G
��E=R�4]�8�w��ۜ7N:�Z9/)��uG�_n�Ho>W�"����:�y=�V�9ot*s
��(�-�B-�.u�<�պO�i���l,�1�#�V���>\\ �1��8U�;�ou�i��3�8N=e��}�'7f*��	P��I�7� �Ǭ,�k;���C�M���k=$����wd���{�u�1JcCp)�I��a�[���m��ͅ��Æ#���nJ�R��:>p�օZCp��ƶ��h���u|@�.�뮞&p��m����9�&u�&��x4��"��{p�{ga,l(�s�F��7ۻ��p��d�`��'+��]o( �E���=at�w��`�m���6�.�q����Yn����EW*4�ք�-�.9�㚅�;�ob��,����&kd[Q��PjX ]�R�&vT�0�M�1�[Y�p�7���zI�a/dX�t�w4^��)=��Ν��(KH�ݚ����]<�9�A���ˏ���tg����n���7�;6����Rov��I��D&��vB�$��od��=;7{���{:�����-�=8gn��g&5=ЫR�T#����'6�'7�Gw��"�,��)�,�\��q�ɒ�}�}��rMũ��݋J�K�vۣwbՐ��B�Z'JHZ�͜ksu�v�Q�I�h��8^d0��qyr�{��dZ������+h��@��@�Y5e�S��6��&�l|��U�=I��-�9����[��z�y:�M.��!�
!�2���Ps�|�������xv�U��EЇgvt������I��5��<��:��9l<d�2�o��K�=�<�úp�p��[<��"M+����e'-
Ǆ[7�Ѝ�ǲK՚�kz���X�5�c��,S�A����E�6����2\�&M�7�	b�2��d�Rwy�����Fq�m�9<[ۃ���wl�f�9��A4�ۚ�#�X����M{e��n���[,�-�����3Z�yk�;���T�,�U�߷��9�e�� %-��_��z�Z�
<��{
�{ҋ�Kon�WI����g"Y��fۀ�gmx�雏�O	���OF27��KOl�%$�]{75I�!��u����gr�v�4�ݠ��A;��V]���8���ܵ�xb�tj�f(tͦ��z�NX6'�r��sa���6D̀=0� �źٺU+��w������3LI��9�f�0s{�Ɣ�M�6H���V��pQY�M�%�Wx�Nw��ߟW�p��t�ٶ~�v��ӠϷ�S	�:�hz�;�uv%l�c��g
�l��P���X����-G�:�b{S0�V��8��}9��!��rb�❏✏vrL�K�g�����`�Lѽa�8�����cwu��3��N��>�O�b�ɪӝۡ�t�#�<Oq\&�QI͕�Lx������t��n�а���s��ɴ2����;�$�E�#����FT9h�o5Խg,��alZ�R���[M;Z��M8�w���J|N��L.�0���y�e�t�pq��n쳜�CH�s^�+[��As录��"�g1���6�S�<�wx���i�j����Nkt�ٛ������@�K6�ta�(�3�M���v��rޯ��9��j48bh�z^7���'*#�F�}m�&��s�T�q��A)�O�r=�Ѧg	��]��<"oϻ{�sa�hF�0�y]����,���A�ʥ�4e��r�}/|�o�F����[�� ��wV]�A�N���n��ʒ��2;�LD�0��Ĕ��)^����9g&{!��;I�o�j��]+��3��s�����L٧tm7��Zh��&��d��m�֚����������Ͱ��503��p��.oC�����;�H�E���{I��
=�x�g7�F��u�n�np"�X~L��X�KԤ�!4�=��6B-��+w��f�v\��i�;����Y�$14M��pZsEx�[��7��0�z:���=�v\��o>����$�۱�j=��$G�̭7RR��-0;��-X9�8v��� J��X�ݍ���̊h�Lls����ڏ� ̔��6a�O�=��~��� ���mn�1̼�a�;v�j&jܓq�ln�n���7@�k�Ǩ��-�/w3�����,�$��ǬƱ�Y�0N����rߖZΆ�3w�7o�R��3�N��r��� +��u�;a�ŤE��6[� �Va�3�����a˳�+��S�Y�!���7zf��gt9�:;] ��;�������<��y�@�ú��F<�vn��×ئ웻��h4��;�4�w��m�0��>ܽ��
��=A��ܹJ �1�\)P���[�Xd�4���8�"�����m*�p���.�3�MQ��E�;��G8j�0�h����म�gvv���a�^KHrw��G><sGuMh�yn(qp��h�v��|u���ݺhW��u�ж��S��-n�#�̵�2��CS�v��:_4��Op�7n�w�|�γ�����\�@_6�[��F��3�4�Gr��-g/G
�����JYݕw�%J�y�횧*�`z��`m�ܤ�|R�&���_R��^Njo���ȸ�Ά�ٸ�Nۖ�ѝ.�P/�B�O���v�c1�$�rp�T��ޱ��uKK�-	օK��w]ӛ:E�z"ڙV�l��B-�R	_o`L�r����I���t�-|�q���3A�0WWO^%��!���y �J���v��GykD�\{p�'�FsM�U�����W�M\Edqi��7�d��L�5�&�x��`N�G/h�bz�G�8m�q�RYÇ-ѿ�wm�{X9$0�]7��#ƴ<�^�5a#R�c�Ì&�q�ӽ�
F��Σ	õ���f��8p�F��1>�����K�okǝ�r���FtٷX��g%�YĽK��0�'���JUpoP�DCn�ӳ l�+�Go˱E�,��8Bw���۵f�sh	co��w�@�uLӠ��ڒ�q��:�K�P� �/9�m������L<x�..H,�L땀pVq�Q����NÃ�o%�x�N�9V#C�4�yό��:w��HҸ镍Ӌt�9eY,c��+;��Y,�U��d=~����gA�v{؈��������&�[+է�~���5�s��w{\
�@�=�Hf�	��ܛ���pq���f���k���L<=�.��)}� /L�����6@�Rf.%��S:5sl�t.� S	���]�3��+I��F�O\�4R����;�V�ݴD��79���A5���%LG��/N�x���.�F	�;{��l�*�e\6�0���Ym��,as����}s�s3J(���.�jA�7�3��؏VU�<�Tɹ�e�Cj�o�m�����ͤ��z��f��m�78G���q�h����[��B�O�䚆Y�r>�ga�{��=�����jm;����ߔ��q[��;t�|���*��Z���ه�W�n��ݧ����٠B�I���6u�7^1���l*��;қP���z��f����^}N����'��A��Q޼r�^�ž&}֥��8�c{�oN�o+h=�������+3Ojg�b�B9wq���0ԏ:<*��)���x��B�a�Z�g׵�Ε]�N"4���=HO"�ʸ���%�f��)%5v�:;9�7$��-ª���[��3�l��Yk[Xl�x���u����^�׫��y������Y���o����|���ln}LX&Q��7�S'�ӠL�k�;��r���a��x�Ҁ��U�ܧ5A��]:�:��92:%>�ԕ�^?��җD4�����rԴۮ����9'q�l�[{��Ќ=`꬞��Mr߇H@�.�6c��/-]L��a��哻N������^B��tM��>$8�oQ�5�'�Y݊�Z� )v�2��}%�=�j}�K��H��.{��G'r8{93��)VWd�P;������'�he�y�.M�k�-�y6.��mN�fn#�m��:�?p��"����tO%򰡫7\;��[�����X+�\'Cm4sb=;��oj�� ;�Z�M�sg4�vꦤ�n���gA3d#l����8����|]��R(���c`Y���z��f^�@�x5��Z' ����hܬt�ݺ��� ;��¦�<w:v�xbz�`!���y�{0�s|qgu�:��0�5vNF�p-�n�:J��nn@�wT�أ7���.��D�d8{N%�y���y ���I��4�]�Z*E�k�oZ�1�.wN-�j<�ǯ�w�l;�����!lg���qh����n�b�ܭTz�%>x���YӮ�8w6���%�m���z��[���=ݽ�p���4i'Q;��7,��&W��г�\�t���i��˵ϡ�FNe�#��KM����,�>�����3���R�XsS� W,B�+�\P�gn���:�To{v��A���%�:����8A��	���-��.�]8p@�@8h�O��ڦ��I���sxzĠpy�fU&�6$�
��tgu2���/�%K�`��gc$�+���3n�X���l|���ۙ��F+�sJ����x��	ݷ5%�NȢ+���A��M���7*����B���4Ӽ4;p�+)�G,�J���܇�b�˭��'�_7О]ܐk�����m��,�Ѡ
���+7�Tq@C	�:����c�FH�wJ<(X���.q|��YR��8�ֳT/����~��4.�͕ٽ�s�����^ͭ"��������5n�D,�������bwC��!'q�34��7�����`��2�����I���:S`q���8))՝ۓwV���;����X9�4r����|��Xt17�#x��v�=�80���K����=a�̻zw98(|'Bl۠s=�j�� "�s��z���9�m$�y�8��u
$ݹ&���e���#&0�5�����u�"�ԇR��u�v������<;��^WF���VoZܹ�(�ݍV�r,���u�F^��q������Y�d�� ���6<�휹��_f�j�p�l��;m��Nq�7P}j���9nJ�������7�vA��y��ۆ��g8k�4�t]�]�oNwֈ�5{t�&�E�� ��3;c(�[�b��[{D�X�4.}Cl��t�ͼ��G%�
.��J ��4�*�uN��, ��*�@�9N4�4q�{g��݉��Y��(]�I�܂��1e�E{��5pR�en՜���N�k۫w��4JIl�������Sv���-��q.�7w��N�U�RYۏI�No\y!瀷]sgD��Y��j�cJz̖L�_>�dg��0�}��o��\r�;'Gm�ء�$�t����J��{5M9&�gi	���*��s�,����o��:�>�oZ-��p'��<z)��wRM
��g��v�K1�4�C�\�<�kbMC�]N� b���8m[�'��z7M3�gM��,��Ȫ�o�����m]�-��U�q˖��b��с&��&�93���'�Ӳ|�q�N��G74�ݛ����i建�����'4�Q�$z�o
K�΃�ǰ���M�cZr��Pʋ�梭���w4v��u�%d{c��QE�=���Zuc3'q�.i��6j�qZ��q�2`�z��_N�h1���$�+ч�3�F�V^�Y�����l��oS����Y	���!�����"\r�0���T� Ku�	b��FF��T�k��������^e���M<߷��74m�ϻ��d@߽��Y\~�(#����l��wO>ee7^��Ԯi��%�A���ڲ1L5�Gc"�#��\�"
����۫^��8ݓ�l�VQGP����{����ŜƧ��(Bz��$�|ޭ�Y����u�Tn�Qē^ ���Pv�}k�~��#p�n��"�P5��R��2e�M�s��I�}Pycܫ���=Ҋez1n�{�za<hU�Rص�ذo-6�wR\�lt\흍���p��j+�-���Lu��p�˳Z�AFvNz�e�Y�'J�m���^0�ٜ)G[�[�쎱��� ����WS�����%K-�����-;p��YJ��G���[�2i��pj��63�N��'�Bm-��������K$���x/�駤�j'I�8&4<�&�e�����^��3�c?�q�q2���s��3K�|K'Id�p%˧w5��~}�1ZZ!g�妽d,�b-�^��ݗ'�J,����^��c&���<I1�`$�����2���Y�_"2��E�Χw-�:ws��'N��ϳ�v���|_Y��!��U��q�|��V���.�O����8���z2_gz,�$����M!&i�Y��/�������u;F8�+���'����2[<�p�%O�^�t�G�7�v��l�法q�]oe�8�I�7F�x�����v���Hc��.�,�D�g5���I�6w_�R{��埉��{3O�zt�֥{H��4�K�"�8,=�]%�t�XV�a8)�n��FF��������B~[e��t�Ųpl��!<e.	�I8��pH��;������D�5�$�c�a��a�~��x �Bcv��SW)١�Y������^�#�������������<Ҡ�@��dƶ��Qm���m�EmQF�h�Z-U��ګ�-������TZ6��mmk�Ŷ���5Q�h�[F�[mcm�5[F���ƶ6ՋmZ�[F�5mb�[-m�j�kh�Ūضգj�m����Ѫƪ�mQj��Qm��h����b��lmQZ�-��[b�k�����-���Q��Qb��+j��V-�mh�[kc[X�kcmlV�-E��mkcm����Z�*����mTkm�k�X�ѵ�-�V�j*�����|[O绕��Ж�_Wt}(�7աQ%P��Ț̾��:���yQ��}��T�����gv�T�nu�Cފ�Rr��\���B�<4��E#�oySH(���i2�é�7�w����&=��xw�w�ld�j:���I[�Ө��L���TjT'�7���ހމ'�5�%'�bO-�$��"u�z�;�.����{�w�S�������Qf�z��PnrPș��뾋N�/�P�Z֋j�ȅ��L��x�����C��� ����!>���)���>��D����������W�w�ֆ���;���Z/g%�w�pV����c�'c����z�Mз����~�6+=T���$�BT����֊~z1+�q��ո����Ѻ�t�Ƃ{�q��7ۭ�f���;�G���3�Z����'o k�IK�<^�y�4��V��;7�7�_��Ԏכ�0�s�{�_a#ў�3T�����J�O����h=�T��,��i�M�ξ��h��P� �\�ur��9����tW��՜7�����z@�[�i�u޽���׈$)����.]�<~B��������Ճg}轱�Yɝ��f�3ڗ���=�{��m�~�U���6��3A/�=���;=��[d _{V��k��
���1�!��8��}���a����T�٧��ڶ��J��ݛ��C� �b��5�T�+�S��v�=�r��P�p��:K��G6C:�˓�:����<��XOo��o���Ӽ�p,��zy�}���+��9��������1@2zw۸F�ϻ/�/Qb�=�����s{����@���}|�u�+=p�l����ܰ_;�)��s�>'�fǜ��S�\����^m�I�Fp���!˘�j�I�`*�1M��
�aǴ�����5�^�5ȯ	�����&/0;�9j�.k�m�g�~W������>�´oes^�w��o�^��̚���'(�r8���n<x����㧏<m�Ǐ<{x��O<x���<x��Ǐ<<x��Ǐo<m�Ǐ:x��ǏO<x��Ǐq�{{{x���<x��Ǐ<<x��Ǐ;xǏ<x���Ǐx��ǎ�<x���Ǐx��Ǐ8��ƞ<x��ǎ<<x��Ǐ;xǏ<}���|�]����
�$�����Z�^�d�{�{V^/cZ���^\qޛ0�����\�����'���z��уȍ����μb,<����Ό�T�ZPi���Uz�)�1���s���8h5{'��.�7=���ܒy�f�#��m����ן��r`�{ҽ=f%�)��t��}�x��oM�l�2�yA�W����
˖%��^�B���g���n����1�$�s[��-���P����=��.I���g�5Y�mr�7wg\,���-~=y!oWVh�z��DBMY���v�li��L����ޚ����{=�O�׽n5d[�qnt7��Y�`���L��:�gz�4���tp7#�pD�Y��w�U��o��tzzz<y����,|��7&PRSf��dI/�(�{���cB�a�O��7�뇺��w}�_@8v۵�^`��F<� �zw�=1� A:n-��g�Q��A�
ֲ��T��ПIu��>Q���pH��y����u�z�9�y<�u�ܼ��}��^M����$� �5������}�`�>�ޯ�wo?s����2����l�%3�����+ӇV�/�2xy�S<<��`�4Y�7�x��,��M\;5��1a��
.����,��1�����=��_�Ǐ<x����Ǐ<x���<x��Ǐ�<x�Ǐ<t��Ǐ�<x�<x������<x��Ǐ<x��ǎ8�8��<x�Ǐ<x���ǎ�<x�㧏<x���ƞ<x��ǎ<<x��Ǐx�<x���Ǐx��Ǐ=�x�<x��Ǟ�g����{<��g�o'"ai��&i�W&�E�̃Qb��,�t���q�ǫ�zO{����-מĉ^Y�v��s��sk��ܠ����[o�O\Z<ߦ�x�����'�/�Z꽡g?;rw�<ak�����޾߽H�1s�w�F@�t� �r�6Y�wr�榥����x�{ω��z��ne\u9�Y�Nc�;����鳌����%[F��Ҥ�IZ_���ac�=���b+��{��ݘi9:f���y���K���'ٻc½�?Q�n-�^���������*�Gb�6�C{n{q��8!��C��Y|.��0���\��>�@s���3	Ϥ�s����z�������|Զ��G�:��vyp���Q��Q�;�&�zD�QA�3�=�����b����0Z	wăwzp3��k��q""��U���b�gf�m�g
�q��Bf������F;� 0�`^K�n��s�]�	׬=i��z��'�W�7 1��E�"��}�����;�RH}��N���}o��9x�[(\G��_ۺb"�8z��d:�_c�<n����a��;+���x}�o���z���9#��no�E�$��w|��5���g�uY'w%�|���׍�2!���oj�}�)�a��1�;]�Tjz���g���z��<����gF��S3�	��|�8��0uW�`���q]]"�u���u��cl��8/y3���1l�=�mc}o�Շ{۬1��S���V�Kq��	�JN�.���2ݏ7F�ͦ�Ww��c:&�w��ݢ�����;�����઩p2��˽��=vh{w|�?��{�����N��iK��쳻���xvna��Oj����7�f9�˄4k�w��^���m�+�0���x�c	��V�Oq�vm��嫼�|��
5�;;{Zo4=�~�mIe��Q�i8s\^��E��'��5˗6����=^_M��u�Fo��i�v��*��^	��/�ONszz��{~���Kw��W��e
@s��{{=�É��U�A�����۰Tb�����[��� ����<l��~%�F��8q^�ԫ�u �+����o������1��Ƿ�>Wu��U��o�~.���ͺ��f+=�4�-�m�b~��ι�d��%�/�=�|f{o�(�R��|_�P�i��n�u>Ⱦ�xiݾ�˺R��F�σ�H���㯤��w�R*��Ȁ�@
7�����Wû3�{��;�tx{�R�Ͻ�-��n�/�4�t�eO�6ufo����͡���R�^��7�nC���q����6��ۢ�p
��oA�x��j�9B8`����]fO
�����݊���=N����<�˦
�ǹ~/{�,��+�WS�����&��=�z4&v�;�Lz`�}%W}��Z'vwJ�ͬ�`����� {��=	QȳN���p�f�'N�����Pi�P:�����Wy��E��M��%�n�M�4���½�^^������G��������]�Nw�_eڰ��{�<����v�H~-"s�*�&ws�T?!B��{�~����O{{>����{f�6���V�	'��A�yB�>�5eB�>�SίF���Nn���}�C-�B�yx/<�6����'"�{;��@��2�^"t�-^~����9M��3��?E��Kĭ�-xw�[9�v�;j�4���wf�L�G ;���ntS�xy�٪y��mOvh���vT�
�:=^�u�\o�}Z�E����۽;;NunP��ﷶ��8	��n��)����4��6���Of1��u��E��8Ix� kd�18�ẓ�jg޲e�-�,S��-� �v��w=���R"�����ᬜ�/Jx�Gq��M��Ͳ���ga��Z�76��6(����8O��ý���:�v����^��j�OW�`]r���o��La����d�'*�緧�y1ˮ��7�� �%{�D/t��4%�Xλ��w�^ٻ�X�oó������/c��*��E;�Ox�n��n�7�#�s�#�ӛ��׀�2���*��%��ݡ���s!'����XyC�����a�1�a��L�wٶ���Q��a�k�=x�m�Ӄ�y�0��&��������	JXB^h�5�;�F��y�^v�/�*!���pf���{��zJHf�}������ӹ1�0ʃ�͢�Y9��/Qc�K�/���a�س��g�*�eP�K��c��q���h�}�wJb�sT�]���m�Þx��y�d��wF�]\_O;y�=�k��RǷ׸�;{`͘K�J����Kor"O�쵎����ΚG��|���Y��W:���'����}����vY��L�9��̤H�
զ�.������9���E�����O:*Q����ym�ֻF���v�KGgd���J��X�0��uN� �8Ȝ��}����@�̼�:Ԏ�g�.p�`]��uI�2�΂��ܽ�s���v>T<��	�99��W�c�$��so+�gO@��ٳ���wu|�Mq�q��_��}�վ>I`��f%�}�k�g
B	-k���.�z�vqO})��{���u��52�r��w��}��g��1o��M8����{s����~�=�oHw<
����������]'S,�������sqj�ߢ�L�I9���w=�쉰;�9 ���9�������,��J�3��������o���d���`��5��v�y�/���������Vj�W���H��̀w�`��.<q��_��������(x.�S�9�4��b~�1�<y�ؘ����
B�z(̾��f�O_�g��Fu:�-w�2�^�q�~n?<�;�S�ծ��8��\�Ӱ��/nY��Ƭa���c��vl��Ȍ��#��{�L�V����FW�E���=M�PA��C|�(��'��^�뽸�� �� �n����`6VF�IM�䖡oF��F4��X8j�M�k{{϶����̛�%�qHO�\�VZ�#�5�ힽ��^�|���nq��i�C��o�݇;�/���g\�k���puw�=�~k6j�C�K�����5�#̬3=�ʿs{�ߊ�q�E��8;ܹ������Vޙ�Q�`�Ny�<{ۯOs���om�v��4��m�=�;�'��Qo�I�M�D�%�����y��_o{�|�b|;S��s�/jo5���<��W${�5�X�J�;ۭX�^>9g6rj�g�o���b�/��):�}jjS&�� �F�d=���^	d������u���}잷Y[���O_M��,��B�û��-%��Vg��݅{�G]�ٳ�v�Tc=�7��_�x��BY���|#Q���ƾ��{�ǵ��qM�w=�&�8��{�����3{�T�>o�bs=�C��&Kw�����{۷w��p^4D��
�����s��Oe�mS��.��ob�nw�=x?rCU�2�Ď�x{7(v�^�q�ީ�r/p�����~~��,��2��2��/��r,��A��l8�l�]��7�}����� {�Ŭ��g�ɽ���x��j*�9�N�ɱ��/އ�$^\���U�{�BG�������Uܽ�a����l�$��#��^�����{s��~��^�*��������9�����</��g<��w�O���j��@Xb�n��vdA���[��"K���;����wp9�X�r��L�*�p;�a���4x�T����,�<n(����;�fX8���;RVp
d(5!��/
X�u����-�&�`�ߺy��.�<���p9�4�����2����G}�ś��(=�.+�}k[��7��x3�\U���6f��,��ۗu�m�Y�1��79��sʾ�!�����tؼ��<�gzR�燴ڤIa�!��}|m�7�'Ƃ��i�<�՞���~֕狎%�h�h�V���1�3��(·�c�gy{q ���1@��C�"!�M �:j�w���`#�X���D�_{�(Wx�:t׿}�c@�˂<���ػl۹�kȧ�r�k9yd>>��	+[؀�.�������,�biB:4 ;ܩ�K�o:.l�eЅ���4�����{\���zg�L�m�ܡ,m�G>��(h�	��sZ��������=~�l�˭0��P��%�������k���;u}S纨�w�����Ǝ���d��藭߼�.�+sY�}�����x�6t�+���g_�l ��J����y�)/'s����<��>E�:y�q���і`x������}�0ǉ�[n9ugn���=��{�zd搱B��0���b^�:���u�R-�E��ܷ�rx����}�/�o��닺��4e��b�GoU�M$� ɕ�s�Ot�݃'c(��Z4!���u[$۰��p�3�A���:��"ӁXK;�ڼ}7����w�~�+vY��ל ��&D�������zr�2���]9������o�����+l��ٷ��:���/x���\A���Qf��������zF4{�M�I8Q�����A�����TF~�g��\�Ju}�����x�H�ðL���LO�xdTy}u[��\-G�ස<�ᘴ�~����{��o7|1��r�cgjy��J���_mƲ��V�2>���}:�g�^���LR�p�`VE�E�˃JN��f�(`)M�X�nù�����Z������{|%���s+$�[��;������ �f�׈��������rck��|���v<-.���xy1�=��l7Qlk)���dA�G��pno��	��/�������O�v��^�/��&��G�{�d��C�jp��n�.bQF+�{Us׺�:�<Fo���u{Gf-/pE����ct�7ޕ�o���:W#�3��u ���b]�D6*Ħ�TfV	��!v����Ț�>��c��x+���Y·=���6��9N�}<]��W�yM��ȟh=���+�z�5x��ҳ��ݧ��
���ì)�׍�d�Ób(P��r�H�̽�ö���ݺ;�x���������f�`\:�'0ý|���e�������}l��Xa�yp�O/b���,�bqr+FOM`_�}6'���"�V�T��簢���&�fj!�����0_��&�pҊ���/�ɟ5�1s�È�4o��Z<@�ݝ���t�7�>�o>H̾]�}{�-ͪ������4���{֟`ի�./,ݹt��D��N�����"��c�؜��5^�W��i���V"�S>Օ��6Y��Iｹ�����[��y�����{w��n�djx�=��{ڏ������Ǖ�r�e���]�=��X�v�rSf����vn5��Z�a	�ޯ�{|T�2����G�~�&OF4[�D��b;��=�N�!�{����u�q�����a�t�lHMo!Cl��/{7�����c��� 5%�W�ŏ�y��T�4]ǖ��y�g�"+����xUE~�C��w��/��������ލ��>ʔO�k�ZKPs҉�i	�����pԙ΅(ʥ��IA��l3m+a��<7��ɭvμ�a��5�y<ĞeC��� ^Ֆ6%�4�fV)�G�<�Q�6�6VEWGlZ�m�Z]T���Kb���u�/W#��Q���gF��4�X��0��h����_M<��8l4�+u�ˠE��4M!���ٖ+rG"c��A��*��4&�qY��[\$EuZ�n��SB6��/���ɬ�ԭ�,\�]W�Bm�|�����WE��̥�%��^x���^.�b]1������*4�e�*��fؖ�\�P�l6���� \K[���n�-�&�X3i�2����Jˈ������L �Z�F��PZ����l֑L��38Z�hqE�YX�
V��f��d�3mUF� �6�.����:b٭ͭ3n��5��P�jK��ZJ��b����4t�����8�s�Y��i%���QL����XME��ᵖ`e�fy�ض%��3��D[A�Ü��jZ(��m,��.����� O�|�`���\�@Q���5�@ƶl���[�n%���挬b:��c$HC`Й��5��.K\�5tmF�jKۍ`@�c�4��6��I�9(�c��l��.�a���f�@�ט*�cu]i	��V4��0���ڷ�aNa1s�&ԕH�7\�:�E�v �"j���Z��[��S-���i�[�l��!������tt�d�Msq�ƫF$���T,#{-�l0�`�%J论��%��K�v#@�u�2�38��6�F�(�)nH�[t6�1��a#a p���et`���F��=�4�[�ٮ��%Ѕm֌v����H���g�,M��,j�p�#��?ܾ��.�����g�D�8u��fa��{�tAmB���UXc-�Q���i�b�(3qu����[��ئt,Be���f��:4��le�:�o:�j���ƉԊ��[�5����!d�ei�հ�Sl-�6](��E�:Ĵ��3��4Ś&����l-�-���.%��� 5vM���U��I�+32����Ԫv��-U�,uK��,�u����f�m]�al05�.b�L[��l`%�	pK� 0�g�Bm-#[�nH)]�]�)]�R�"��ΚT[Kn[��43��U�V7���V��.%��
�CL+m������:�A�D�Һc�D���h0K��VU�)�t����H�d��G,Ρ-�ae2U�nz�X����r0�q1�Mib\��W$ss��J�-\����Kj�F�$ɺ�)�����0mtH�Uv̸6�aeΰ5�+X�%�/h�v��Taζ [��a� qu�e����N25-f�E�\�:�
�S3;W�K0 )V\�1ȥ(`�ͥ��kR c`j�����Ka�2��$�3�`��#`�\s��YK��)zhl�VcV1�9 gi���@�J�v�iy�.l؇X�&��1���j��%����z�a3�Y2�Bb2�+�($t�ձ ST�uF2�	K��2�h�P�Jʪc�͂��!�(]oTb6ʐF��X[�`���sH��6����:�E����/�';B�v�K�ñZ�����t0@Ii53�Re��Xf��KB�\�fYn[00�,�k�b�Hf��ZG�.�9�M�;!�\�F��ۤ9��J�:h���qYc�0���M�-B��Q�2�XRl�����Ս�p��g3,Z,t����E���K6�͠M��l0Y�ʾ�.q�p1-�[��Zl�V��m	B9���3J9��\�m��62���u�l̰H`�xZ�Yr8�عKY�Ю�,��p���X����Մ��(F��:�b�k��x�y曮l�iL�M���`�U�%\aMh�n����R(�z3C;Lc\�#)1^���%xJñ�7��pv�a-��t�v[6Eу�`Jm��s�N��	�uH��b��.c�+�R�G7%�]h+��a�5m�4��d�K^)���	�Qt�Vj.b۪33���JmE�v2%s���μ䆮��٪�;m3Є�h�nu"t�5���6Fm�f�k�i��ūjD��Mev�d+x��6�>/���itT:��+�pY�Tu�bf\�]�x�9�f����<+֣�t\X�iuԎڪ�-v��J���Q"� ͤ�-���{��3\�e��t|Y�	�:��]]`��!n�n� jjIMK2A�%���f�iY�ՑQ��.�I玽��-�\��)���8��b-u#��,�pʹ�av�I��0�����B�3
a�R�BۥZb̪�79L��]��K-F9��ln�j�V�iq�6-r�Mv+nJ����
ml%lՄ��nJ��%+i��6�"0utfz��&-����J�ۨ9#7k�b�)�+5e��l�����f��F.-��ˊ5�5%\ ��\�q��t�P����X�&ف��F�����ԬW&��c4�--�t�[j<l���Z�KZ5Վ�II��L&��\����2:��M��0��P�$�m\�Ф�l��a�k�!�F]����ZCvC�!�����9�+[Z1�©m*V6�t*�u��U�m&\l�=�Ѝ�hR<lƜJ�5�`M����.�b��R��.���0,γT��Ŕ3�z����!�c�b�X��F��KY���S�z˔\8�X��-X�s�:�v�%`�Tt�S�e��y�鮍.��(`�u
���	��P���+[D��l�m.M* c;"�-�XIv��(�!��t��.jh�0]��1G�lb�X�ض�I�=0��%��6ekIuX	h�`�M6Ց21��M�c@�jkL˖::�&m`]�HR�&���.Z&��Sy�ճ�)�+gl�0�e�U�a��:�%�9�d�#�E�
�q�mNi�;m�X]k�m������l�q�����ųD\�H�`j�L6l]E�+*�fSU��Q���xv&��WE5��6(@3�e�En��/ґҎ��VK���x��f�m��bh���4��G�ʶ�f �Šݥ(�n�%�-��P�NSp��)�3iR⍅�X�E/lcC)Q So<���2�V��#�@8�,���aX-����K�a&	6�n��&w�G���BV��C`�u���6�Q���Y��ck&K��:�JR�k@�k�+�&҈�VMG`-�c0�fu�C��C��84%3j�Ee�+�u]U��+�t%���δx�	�I\�"cE�v�Gdu���%��g*�X��j�)	���
Ŵ�km"@�*au@WK)6��$4ͻYv��KFi��+�Bf�<�^���P�[�3�A`*9[3@��6�ln���b�	[eڰ��Z@�	�k��%+B.�̖��s�4�aC8�z��h��\@�u�ph��XC��[��,�B��Źi�&���	M�Z&�8�BK����f6Y��05�%m���q�@�[ck���Tb�U��vl�E�p�D�(�	�F�xe�s�4��uт�n�P58ⱺt�!tr6����lj�"[��0�a��jˡ��s�u��ʑ�i��[�Q��4����Y�R�����	a��WJl�j�l�5i��i[�C[fRMj956��W1�cE� �%�	NZ71�vZ�L[6S �t �5�����̓vwe�ʦեt^�iYeKZix���gm�3�0 b��^�s��BR��*�l`N��u�-űK�uc��WZL�Iw3b�fj`|��<��ji,������8�K��5�l#���"�@R�B�u��;1��[g��k��6�R�q1�S�����sZ��v(SB�R٭bR]����Ui�kc��Z��n��p�֒�b�]q�J�q�.�.�X�66^+X�Ժ��ŋ��*Un�V9��BV6�2��1e��LlhS�&�Ms	�4�"]���	0�u{&m��5��KR�e]�{G3.��JG.M��e6��rż��˲CX��.�th�-�g%�+�R۬����p\�mΙ+��HͶ `�[�Q�1��Ԛ*�lEڂ�c�r�b��Q�ie7ZK)��%�kf�p]���1���K&��qb(�ҷGV���.���7Z롁�TM�kr��m�T�q�(6�s΋n�1�5�aa����b�[�P6SL۬7]6�蝒X�*F�*YLGV�&4c-�PA.3li�Y���:���iEJ���e�n����\�-��2� �u]e�Һ�pҡ+��e�F��&���&!ū1�4�&���n��+*]9`�ظ֘!�W,��iBf�Ţ��3@�K��m0�F�sqq�&�����H)��R��\č��k<��YH"��d��p�@ǣ�	x��x�Ƙ��J�MFe�B��u���B�fWLX���ޙ<����i�)r��3Lp�a*k�bD�
���v����8 �0�Y���M.u���H���ɶeX�JӳR��s�E�/h�m4�غU�������2�,��E֭��t-���Ŏ���� �(i���Z��F�,a��f4ͅE�[���usu��L�sn�	v������Kl���E�P�5 �(��ݴVxO6��M�5�],��Q�A�mӝ�ٗ13�Cg�gˎ1Xf��&����]nI�<�y�Z-���a�ٳM��pq��ɜ�����8��B�k���8��1�Z9qm���8ʭ�5D�氫Ef�-Y\ˮ�I�#-R�
��W6���°u�71uV6r�����41�Y\��`D+bB$�Q�u�rY��hl��j���Rm6� �B�t͵�8c��#6Q�`
j���5���[s�DF�kC �$͆�ld�~>	,��_<�+g�t�F���!V7kL/T�e,oh&�SB�a	�b���5u)�#&B�i�1�,�2�յ��,b��,��n����tVl�cz*�n$b�q1�ھ�ؤ�����d$���A��?�Ƿ��q�q�����[��� _}�*$�r����H�֊?K��P�HBm���ǎ8�8�5��Mrܨ�+���d�cL�lQPE�r�c��Rb�)����m�5$m�lQL*�Q���F�X�`�X�QFѣ@j5ynb.�E`�X��[��U��\�1X��]��*1�&�Rh�W��(��ͨ�-̚��$�������1I_=��G��Q>���B�fnj�n��v�W3���Ф��k��n�3^�֗9���<�w_}��N��˛]s'\�7;K����i��.��;���\��n5t%,�\8W+���	۹�Z!sr�;�t�S_]^�rbܹ4�$����9�W/�_ϝs��wrh�[���8t��v���]�s�r(Y�c��8����wwz��_͜`�
�Ѳ����v�:R���#e�"�pBL���P��-V�ke��M4��\̂�$�;҉��ڨ9�ݖ,�@�^.��3Q��dA�c��2���e9n�u� ;DJ�<����Z3hlJD˦�(�\��ٕ���6��j��tv�*.,�lP\�׋3b�l Q�2����!*T�佘����%i�ݢ�j���b��)Ʀ��	0��.��l��!<��bl	6t`l�:�����L��W�B�fYU����fq	kqo�sN��5	K���TŷDCLn��G!i�4;b�iQ�]��-%�@��@���`���i�LYs4p����1bԳm�@ա����ZA��˖яLKb�)5��ʠ�m��%vf�v&5�ٴҁk����8��v3�i�e ��T�(��KDtc/[csB9���oe�&(H�,6F�$Զ�4\����톘&�%lqv�kݴ�X�[v�Z�'+��a�%fl��U�BCfc��s�Jl�����h$!�&�p��3UҐ�V*b�7\
r��c	m��2K/i��4��h8&Z;W#%����77]��9`��雬� ѷ��v]<�@���勱ln.���W S�l[c:�m�J&ٍ�V&P����n%��Zֻ�֠��3��JKV9D&t�$ͫ2v�f�p�mu�b,�)pk�[x���8����Yxe�F�Em���&��mm
�m)%Yy�����G	JD�ݠM��v��Z��\�8�X�R"V6��6e�,0�f5���%��8$�)HfڬeV�;Rk�֊�z�u�	� 6@v�`��J9�$ѫ��5��i�ݱ�V�ݰr#r��F(�nf���Ԓ��Х�4Ԯ-1Za���$u��U3-[�����L�il��X����ks-xk�Jph͜Q�r���n�VFfQ��ѕpJu��4�v�5@u��92Z`��M�q;������>�<�������B��h@�`S�0���5���kjT`�TQZRIb��*���ke�b�u�!aDF��9����P�
�dm��X�e��6Մ���ƣ��c�#Q�Y�^�Z�R�J���ai��[%4��a���X%Q�
(��)�e�s!
�0�hSY�"vC5y�%���Q��m����D][h�P���������|3t�};Ǵ��㏻��T�~ɋ�3�+[ۍ�$�$�&�V�l<4[F���o�-T35�R��1�֏l��d��0�� F0�V��5�v�&I]ff*��X�J�|h��g����\���J<�I�U>QO������qǒ^p��u�ٛkY�ɥ[���9��pI�jY��>�R���k�$��I?��l��K6��l��N�F�*�A��e����3v��`�๟�YW����G���1�U͈Z��jѨD���4��L�
w��ۺ�st��^�o7�F\3��]�(��JV�g��>>;n`�$�%^0��q��
�A�I����q^uVN��;w�ta~�̞���|Π��#�\�%=�#�}��+0��S�i~��i�Z��,�Ͻ?-���X�5�;8��,IV��qZ�	vэf�'��K�{Oۺ�O߾�9*����V�ɥ96�vsa$�	2R�_r��Z!E���nO�-�)5�3rDe�=�����sml�����md���┤��M�L����˝r�N�iY���l�ѥf,J�}�o��	7�H<���ȯ=�Oާ���~��D����"R�3Vi�v*WYWQ���$�F,`�	�Ofz�_����8j��퍊�ٰ׍v�Y0E�֑s���_�,�	%$��z��kkM���JہYsu��5�n2�]�a���)l�|���&�z����n��gwVfﱞs�����q~~�;8 �>y�G �>Cf�(yG8��=�A�<{��^�R�:�2r�
>ޗ����D�����l��{!�#��x�a��g�^e�XU��w]�K|�m�wov�S��/�3�ۋhy�VHI��"-f��C��7�����a�.o`CY5 bq��I%>I�Z�N�i��4Do�Uf>f��ɸx�Yw�彺����܆w�� a\�r]�;33���M��!
�265�3�jb�M����=�K3%����~{���I����]�k���y�uS� =�f��#�W^[>Y!�J|�P�X�)�e��,ƭ�U�ݝ��ܶ7�-{햽d���5y��$��]��I@T�8HU+93j��m]m��Sq�e����V��oO��G�(zԈ6�"֛�6�bן�ٽ�Қ}�y�u~��Z��T���խ�����DC�!���u�80kU�ۮ���'<� ��i�+�"�A�OO-�ZW��q�m!��� �L�<ʖ�)8	2L�$T�1�:�F������E>�f�yO�l��o]��]�\?�������'����wlKyc�e�Q��u�v�\Ah�!��0���jg���_nϖf��n��Vf��-qKZv)��ɶa07%ìpo�����	9��$N'�jۼ�qp_F��ʵ3�X�V���Mh�����"���oW�N�y"�b�T������rv��Kj�kǔ��z��_n��8�Kʏ�V}��st��Nۿ�FYئ����[����z'n�a�ˑ2ޫ`�p`�?�Y$eսk5n=��u���ྍ7y�jg@��ŷw��s�;s7�s�$��� i��>�|1>͘�vg�-^��l���D4��d�݂e\�t䧻5�gQ·޸�V}�EY���{'~/�z�_�=#�R����u�m+���+l�J7�Ys��å�^�L5`2�Pɬ�.�6��
��p�mq�&o*��f�a٬����bn���ԃ*�q�9�r�=P��H�X`�)c�cu�����ֺ��Ζ8ÝkH�kՖ��.������4���B��%t��C]��]������[lk�/eeWׯ<,%����b*;�.u�c�����&r]Z9�%�� �ǰ=�P6	W���طn���m�mX����Q�Z�	v��%c��Re��a��x��a�72T�����t2��5EfhY���dd��1���	�7��\�ݨ���->�d�$�%P���f�>kP�8�7'feZ�ѵn52L�t�>��3ᡯ��8�o���Zݣ�M����#[�՘lk[�����J~˙N[���� ��6��tm�{���o|2[j<⩇��V$�b��Q%���``Xݝ�K��X��Y[b%�8�7�[Ƌv��2�<�~��,&LSMjY���d�l̫Q;�LZ6uZ���S���U0Uf��|{ǋ�.��zy��Q���j��!�6����/ދ�yj/�x�s�4���껩���Y� [;`���U ���n�}���v)�c[㸕�Fǜ˄������3u���V5UT�yH�ت��I;�竸Ń/����!lfڪ�*�U
m��,|��r�e����A�����+[�n��Lc�8zl����©���j\[^c	�Xþ
 �w�M��o�+_[��f�_�׮���xk���wb~iR�Km1��0�[q�޶�D�lڼ��*mY�}@(oN�ST��N^i��&n�Bڋ�sJ�3%`mϟY���L�Ray��Y�cr��P�ۘ���bϣS]�b��{i��©�����Ƕ��-�֛Ne��z�ŞOdo��\��C~;��7�.�8����g����qer��l\��#ڤۈ�$�Gxy��z4^�R���Uݣn�f�y[���y5L*�כ7j��1�� >0�o
�1T���:��uxr/}��iD��4�˓�NJ~oۻ�뙦��ﷹo���۸�z��,��MyX�6�{�0I�T�����}2�|�C<8%�	�ib�Q�K��W��F��\.m�	wP��5>y����=zg��S�񛺑ˆW�s�E���`�2r�����=�JѶ��^���*�5Un��֘y��8�A��i�p�y���wm\�����������6�s�����p�26�i-�0Rl�ˑ3�Օ�1T����Ԛ3\V�0��go�_�����I��7sQۆ��9�U�nA�Q���L/ݼat�����7�O��4������g$�yn��^�|���Tn���؋��Kap�U"lk�p�r"��0ޥT}M�_�zZ�/B��1�����وy��8�}��M�X��2c3�!�����5@кY�,e��& ���L����	vM,a��(��fӗ�-9i����x�Ί��׽�׼k��~����)�Ps-�,K*Нzږ�^�����+g3h��Z:/kF�ƪ֘��7�HɪŐ*�
���/u�f1S]��l��ۼUY�e��r��?�z�[]��M�xgG��l����vv��?������I���GB�Lޯ��e�>p�L*��i��a��q@��qU�Gn-�m�(R�6[�L*��ƾ@��P ɒwa�-U ��10�c+h�X��_a��w�n�����������X�ش�M������g�8=�%�։�1���o6s�$PX|�]�����]�2u�ٺ�L5��6ځ�5"fXMQ��J���&&�yκ°�V��%�Ib�לf�]nф�p�!�C.f�	n����+*R!��2��!�f�ِ�M�sLd�s��m�M[M���s�Ya1�`�f]�f6H7��/�`HZ��Bi@��M4t��30PpJuL��n&��YdC��t�UWEx��J
��Ӄ�zv\M��aњ)ěc@`<��⮡4[���m��i6"�\�����0�]�����[��G���;S�;�e��r��Ƌ�{�n���Q�tޫo#��$q�J�0궤�o3e��^dM�9�šC�L��%_�-���b�ͬH�aJ�z�a	j��E�U��[.m�=�Mh��
��S�my��x���m���}:j�����?zwɈ��×��j�Bݩ���Cx]7�S
��ԛۛuK\��S�U[�����S;޳|2O��r�זˍ��oAg2i�'��>���� ���"j�z��tլp����Q�1tD��3&���{��zoWש(�c�BV��+�[6�f���6hs5�Zr�S��{�ߺ_�r�*�°�H��=iS�D�sۻQ����S�z+ �[|9}�r87����^Y�G:8Rs/ĕ
Q�HMj�nɘ{Z�͗��N�;S�;�d�L����)��aT8��{ŏ�g�t�$��aڭr��/.��D�ȼ�K&w֛ӌ*��G�T����L��c!�j���whM�첛������~g+U$P������d����ְMT«��r�nX�0Ź9��tK���l��\�^ž�v��[XMS"f,E���_=�_Q��af̺Xͩ0)srn4B�������m�a.���Zaz$�	]�5����1��J�;����8r�'�cZ�v2 a�u�L����k�N��ۑO���3o��áV�e�R��l0���\�/7�n����|�s��[s-̀P�!�:�7���(R�N���{O���Y�Ui�^)>�ڽ�[\���b����Am���==��y7f{ۈ�ϑ/\�/8�'��������Z���<��#���guԼ_ú���VB`���j.s(]����G�����b�RM/��|b����)י�1ɾӪ�\�w�~ˑQ�?P{�|�y��%�o�g�{���<�X��o��/d��-�莋q��sZ;0r��ߵ.�d����g�tbk�Ŕ&�g�]�Pjczҹ�����_i�\O�^s��0,�w����L�mJ��
k�}�?������)�}��αyg �2�y ��̄�z�{�?#aZ ��jw|�����V>�:43�S*�I��VD!�0�ߴ���U�h<r�Ƿ^�|�'��1�*���j�%Sj��<�9��,��eї��7ym��+�+��F�YqL�Ӳ&��^�L�}&i�ۋ���1Q�n�1���g��p�~���+7Z��y��A�!B�Od���y�}��+ݰ�z�u`=�Ð�x\�(����r������*��U��0�x�w'��D�����=Ŷj���p��	}�7錱����F�觴M���g9�O��ɸ�M3��v���)���5 �]�`}�}�(z�L���:�ʲv^Py�4�w?Mg���}�[�Z�{�lc�a�ٳ��S��L�&{���׹,����,f�R��Y7�N�ds�]�fj�����߻������(�7`ψG5{d�ܺz����sşL+��gl4:����I�[�X�Ge�d6^^	 �bqa�Nz����	U]8*QUMBUI)ܺ����P�:';rwr�W5�E}�ۯw[��$�E�*A�;{{{v��ێ8�?��������WJ,l���u$m{�6L����P� ! G�ǧǷ��nݻv���D�@$y�ߔ\I,�(��y���\�������h�o��"�$�+2�.]���\Ư�v�6�܉
"��v�5=�չE>�5��PV7᭹�6J��-�kp6(-|���F�b-b�X��cQ�H���ͣ�W[r�ܪ7*��t�y]6*���#\�����#k�����M[�����6�Z�j"���sc���W6(�o�r*��%�1�|t��5z�||G�3/rtf�h��Ú=�����b�2�f�fU���ˉ�e�/�WU�������kyzm���w;�`n�8��Q���9��U����x0;��{чv5�ON�}�v�Nƞ�x�?y��Z�d��r�fG�x��}����2���k\>��7��jR�6�xzm��L� �����?�I�ڈ��̦��E�8"�	���ZT%�����$H6�5�W38�2���Δ��@��M$y&uV�t��&�&�w�9����s�Y��{!� ̸��I���8!&pCV�wv��^n!k��N��u������OUy�[��&����/73]�h�5����Jl�����,��7�d9�r缿/{=��*� ԥ�6�w�\�G3��_5����7l��$�8�u[n�k^;��<�A�-��y�JL�U��o�T������� �0r;�q��i�L\mt�zqN�M���]nt��#*§��<[����n�`e4�s~�,�8��W�<�NF��4KHEl��YƐ�К���`��n�������,�̠�L�.���?d��{�sxU�VX����U�v�A6X��2�o���8 �q�Y��՞{�����7�l�iE\Ց����6�v�6Eɒ�e�Uh���QUr�;w���O{��7�^R�p�������b�.���ޛ�w�����;��� �]��\�.'{�̣���$
L�pU��<��=�fg�޽iU�j;��:��Ý����A����ȼ�t�U%y�G�68XH����p��$�ǉI��7_��;R�|�|�?i39
��n1�����C��������&�9�N�"���*⛃֘f��Óxo�!s�U����+'��B��q����t����)�1��N�-`&�{5��H ��{|n�P7m��8-=L";�(���^�W�7x�=����lÏS��3�P �L��&)��zdC�l��Rj�7�����!��ɌB��s~�ڗ��.��C����i���\���Y�vջ��5n��@�vwq8�����*�p�_\�^��y�gv�%�&���UL�Jb�&4]u�\#��X`.�"0�R^H��p��j���s���QR�n�Jb��B,k,�DkZ�)�;�U�Yf�z�Xu�0L5�u�2Ɋf#�P�"u5���3��u�u�-e�q��k)����31Qc]U�%Ņ�DtvM��aF��G���bj�hT��VUw�~���p�OL���B;R&��R	�Oq�5F�Z&^%��l\b�����`�C=M/����4!=�Yk9	;��`��ou;��1q*o8��]6��Ȯ-�a�6�z��2��E�2�bkg|��Fg:��(A��m�#�3N��L��z/�:Yρ�p�������/��s���g�7��$�}>i��u���n)����廕����������������O�	8s�)0��֦i;9� ������p�!2!���^j/Ä�ĩ�������]��e�����EK8�]˞r�=i93E<�Bݥ�&N��M�= ��{���b�R�#G��=�x���r?�[�ͫ;S���?|ﳴ��})�ԅ-�q̣)n �\ķ\�+��79ڑc.�T����;���>w������힫z��o1k���9�z4���u���k�Rj�2�̜�B9��/ł��6l�u_��Rc��	�Q�>�j�_��S��0��-O/�f�^_�#��O�����&������ݙǚ��N�%c"���[���a�6�r���c�(}�:���r��g���#�c*%��'n�
vr���?�M��;�Ӭ}`
!�/7��3�u�� !�x9E��޻p�74�Ɏ `�F�oM�4PUK����xp<d���]����>;͘�|+#�ks�1ܷU��Ưm����g o��p���^N�ŭ=��70B��o"��
���mM��(��n\I�[�,�2d!�8!!��#z���s�W���1Z!�^m�{��XV�p�9�L>4�O����;������n6�����)v��8z�UYm3�ݮ�#V����R˧��~��#�xG���'&�
N^�F�3�UW}��|��[^M�t Zol���e�C�L G�&��L&Q��P��OPX��f���[8 ������mi�^cw�{a�/�n �QŗL( ��X���I�� ���|AI����;p�\�/�b���z��Q6�X���@�����cC�˲�ԲȲ�2r�_]�{m:_�wh -,��q��e�7iv���j�����3y���x]}z��<!�^m�|$��Z��L�Rg�I���ut8^��xh �p��	�L[������M��|�c|��:����;���N�L����G'�A�o)3�'�x8)6�a�U7ϊ�E^ �gz�fuj��1�������8�p.�zRq�¬�������Y����)��Ss@f%/fgB��3B��sI�0/��~��6���n����&�����T���W�;q	�]�3�{���>�Ʊ��
L��&r'��0��c;(�i7��W��p;�y�̎<�H¾�;�|�� ��az�]�N�FM����SI�3��#��&r	I��Y��HFS�NK�_u���wy���{��{�Q�(�Y99.$��&[d���f��Z9=�����K��]�&D8nW���CԎ��;��	�`�'L���ݵp.�L����@�r��HUV�^�VA�~8�ˡ:�����V^:��XnX���_Q��oðx-Z֮�{�*':������SM ��O���73ڰ��.��&e`uë���b���~O[Yq�������k�����������6*ΗG��,y]=��饖e�kZ���x4aj�eV�f"ԁk�V���<�S�������9�g��g�ͽ�͑��������y�+~�ܭ��&0�[;��΂��91w�8U7t��1"$p��-��oA�q�,���4TH�*�qۼ|��y����rMu�dh���g�7��$q���6=��Ψ���\��գ�D��X:��=�þk��'e����pBN�'&���V�ZiTK��oo�޻i ���v��6GV��cw�#��`����[{���W�G�[�l�0V�@�&��6l�>]�	= �jY嗀�KY�>��wW4ECp��y���w�A�|��Rh�����&��*���L|;s��U��`Ÿ�S��c��k��{�\��:���uÈ�{��9���)���R�U<;K%|@���%4Ң�s���:h���,�C���Mm+��c1euئ0�N��r��.�R�q��PF3L� bޢ�u]���MK�.!L)"��jh$ĺ���0p�e�q�PƆ�ƅ*[v06�Zd�h�c#Z2ŦT��a�14��V�u�D�����ܵ����7-��]f`��KFM�Q�Ff��6@�����I74l�B�kR�]4�ѩs*�����ƋO<�����?��~R��]��X99(��ɝ�A�X!�7E���Z����qo���y�)!<�/m%ovYsr�7�/w���4�/M|0����7���U4/޹���o��5���7�:`fWd$�U���YG2��	�x�xP9M�=�z��%f����-a��ĸ�L���o��;���gtl����eZD��Zf�BN�R��pԣ]؎fx6=^h��Y8��%M����o ����H��cv�9�۸g�PT�NS����w`�n���?�!'�Wk�A�R���y���0�]4^w]ʝ����Q������i�9��%���OW6�.��:�1�d�n���;1m��
�\�9ި����F'rH��A�N+9��U@z��K���w��<s�u�K���v�d���@2R�iqB]0Fw�D�,��e����&pR`�J��a�!��ʪ��v�:��cL3�L���8 ��9�N�I��f���i�&4:��ݤ1�|ӗ�0����4�v{O�T�,{�T����з��ɽVҧ�����o��z�g�:�Y3&�8�I%mȺl�®��]yE�~�'�i�� 
��-��| �y��]�OҚh�<��y�:d�׮N0Le��T/c�ps�}X�p�N��j ��������ّJ�nj���&;�	�`10�@E�$�%!��m��O�t��z���)&D;��{��˃����v�A9L���Ûj�g�ڕc�X�8 �L�!��C
L�L��d���Mz�t �8Ok듪���6�&<t�r�!'��C=�;�P���c�&[΃=#Q6�]�ZnL�1�Y��lL�p�a���xa�����h ��r
m>Ra^0
vz�՗�7��ڜC8I�a/;���j��~������Eۇ�y��?��p��}w$�y��48�E˿���.]���hu3W���x�jgQ��ٙ[2�Ɇ�����a�$�`]��FH#=wU�;�αg��;�U��M�/q&)Xh�=�7;�+���ٽ|	7F�����yO�w���</=о���f��y�;�3�����z�ҢF�P ��e�7��\1��x�o��O�ׯ�%/�"�&�l����(=߽�ޱ�2!ͦpA�I�;�������Lpou0pE�Α#Ӭ:\w\8!&�>���IF���=>�6�Cd�����S5y��Dp8��GHsv��&��"�w���s��~�r��j	�vrt�"�BU�հs1[�Y���1a���z�, �`��7�?��@6l��s]�f�]F���5�pg&r;������r�
���&�)3��lG����;��X�=�������۽��-]��9�Ls�D0q�,�Ãf�u�[�7?S� �Nd��4x��p�$���/1��L�+.��E�k��%�i�\��3�Z!L���x�Sy�6�)0	4��v�տt]��yk����e�!'�ws�\Eu�s|���2\�˚�͒�-��-5�~qR=UGBq�_�{y#���b�r��;ǳ݈��c��ʖ�}1%~�D�L*�X���S��F�!F^�xx�%4����C��a�k�-7l���l�ȇ)4Z
{���a�=�������K-����XVp�=��&6�ȣ ��uEX� F.�
$�pzc�s��v�P�
��.sWE� �R��n�M�84�9�fYz��t_��Bu9�Z��-u��+!m�Wݦ�.��j������UypZ���Sᕐ�oʶfU��+5D&eqas�:�n��=޷p�.A�+^�봸��I��6�!ۃ�vX8#}��H�TGK�/�N'��g �?�4�@�0og�#�z|ڙ��cKЙ��l�2�<�&kc��7WWXVh�,Ûܘ9Ӈ
L��9	8*��zf,���C5;x��^�����wn�n���L��c�|v�o�;L��� ���i3��y�M�>���v�8�'VО82p��Wiqܓ��n�_y�;,�f�xf]�̷iT�S���s��_ϙ����%���ᗗ�ٞ�h�ԏ�������y��_/;�;�RG��'��i�o��_����U{��<׫�<>�XE&�����^�u�M�y����A\����O��|χ�u��NAi�GH��,��*�"���i�A��\
hP�5�����_ys㺼�o��i�p��o=����9.�j���Xn����qӕ��g��Ys�����7p���0��������۞/�	C�xv�ʼڼ�I��<d�z�W��{�c��$8�������Y2ж�?j6����#��g�-AF�����E^�|1�|���N�V=yI��P��w�:������03x���|�d�y�^}oz��4�5^��3޴�瞬��}�0B��_bT�[���6������\���y����S=㽒{zO��:��@Ѽf�޳=�=�A7tv��{_-n��1����m�׭���r��*��on:��I}q���9ޞ���ѕ-���%����%o�]�nj�]�Ӽ�� �6��}�KGyN=�%�N��׈SOo�,��qۺuif��^��c���yk��U�%� �qA_Ȼ����!���x:d�Y���C��r��`��<��nEr@0��������e^ӽ�ĞB�F���f�<DZ����ۛ��c<�:5	��U���& �znNպ9q�N����>�����Ցnb�h��^m��ɾٹ>�$kݞ����]!Ԇ�u���/e���g�Oq���%pi�&tDHݱg�]�FT;���H����}��vE�rA��k5֪���*#<)R��B@45��h�,�o���^�󛶞8���ǎݻv�۷���9 �/(�(�h�-��\�ʱ���\*Qj��M=<{{x���nݻv����@��P�D����/#a4���<��o,�nN�Tk��lh���+&�4X�sn��ȷ�|�ە���ۚ/5y���⹰�����鯃W������+�>{Qo�E��+y;�E�&���Ts�r�E�w�n�r��|U�tGJܹ��E͉7j|||T��sE�F�mE�ל���Qs���r�,Z"4{��.�y�5�U�ҷ"}vܟ]���X��h�����h��H4[�μ-�{��*���^﮲���ll%"�[���p��2�7z����7@�u�A��(b�Y�f�:Z�[`ۈ��w-�!C�S���umekL\_KM��]!YUn��X�B9�.* �5� ��Nb]����ex*Z���u�H�+B��
�V���c\.�6aZ�pJ� ��f&���	��J�64�ʉ5�+���֥P�x����<h�g3Z��l�j0��j+L�k�3R#6͚7-�Ǽ�����,&Tp]f�Ie�L�.�v�uuX�I�2��.2M���3��[5���һ��T�Y���Apm�.ٺ2��`5֝fqv�pk.�X���XR2�l�6��f7�e�$y��F��%,��-%I��L�����V��C��)	���k�Pdnè����vbQ�QAn$��:�e6̳��E�5p�;[��"%WU�љHh�m���֦�J1��0�j1��&�ʶ�)r�5�r�ZhP���ȅJܒ6��X�X���q��sΘ���������1F�m(U��Q�m��H�]/[DX� 1��x��SP��\�pgk� 3M4sl�Z%`�rB����؂F�V9�L��:��YEҦ���Q�)v��Chūt�oa�mX ��Qإ���L��x]c%	�B���,��,��<�Ɣ�b�\kuQu������ٸwx��!Q�B՛��ړkY�FXUu�&J��6R�԰��Z��vQH�.� �R,Z&����v��9ۊ�������h붰�����I�,ZF
�5�d䚄���P��.�3f�d�<��Ҙ>%�,5�i�2���Zb�
a�h�wb�kiC �.�G(�!<��w���+t%������$Y����E�KyB#JL�+���Wcn�7dbCQ����[�� �\�6�#4Gh�̖�V��JJmjݤ�p�1��Mrd2��va�)�s�&�E2ܪ죫����s�`�`�`t�魦ٖD%8�f��U����hғ�Γ���q�#M4�����|*��Y��5�u5Z�	��iX6J#Z�Ì��͚� 6lEWfմm��)��Sc�a�XhVbB�#+^Ix{X���v�V��SQex�3��hr�5�hV�P^ZKH�SCq���8	5Т��M�Ħ��ԃ�5�lG��)�VV ͝u����s lȣp�v�5Ζ��z�nZ���y����V��	J�7k�Yw�(�-�"a+���+4v��0�%�m���H�=_Z+�����Fb�-�����|��at2y��nհp[Œp���?�`9�gD
�5��j����p����uٜ!�Bz�W���A;L����|��M,s���9��9�[�)���ՖL�.̲a�D%��V�l��/�2�����vX8 �	K��'����N��5���;A��V3�A�I�U��Y�'�]FYp`|z�	��2��(� �8	K�QE�)8��̎�1U�T�z-Lh�:D?]����-u�*�6ݸ�u3����&r&�2�5�%�;���e���.r��g�Tl%V���1+cbX���ݸM{3Cg-#E��0�u��Q�?��Z�/z���|f�3�L�|Q��yő��k!�Ro8)3�7{0���uL�j������!���,̧��/ط������i��$T-}���ޒN�*�7���|X��]���+`��S��}�_Z�hQ@<�9���g��zκ�R��O(��7y����r;-�6]���Li�2\��p�BpȢ'.����j���&�Vmn��U�+��	�a��4�g>I���3�N<�0�Wl]�˰L4���
N���w;@޴���ϼ�K�����f�zX���|SiRg�7��'�����d���5Mk�_+螵/x�y��A�`����8pR`���kcGL��U�p��X�lb-�[5�]�^. qE��D��G�֖�6i�}0��a�)�����p�nd{.�tCp3u�j�6ݸ��������|ͤO�=���
M�A���i�����j��>}�:�Z�v�ܩD=���x8 �����F]��;��	N{e���gc92>�$�AH�//Q*Mo%w���e��p�]S�jbY^�owf	��w�1�	��SQ�-WO���1��w��,�\C����|$<|fJ!�q�҈�J��}s~<��C�5�p��`O[ �Ӈ!&rI�����u��t�T����O@�7�M�����c�GWU����u3�$��a��5��,'u�U0r�ES�T��[D�t��/c6��w*Qx���tX��r�\?��>p�%&z�O����[���/�C�P�p�8\��%j�i�(k\���.2�՛�����P�r?��?O�[��}�9�L⻻t\gGZ��Oy޴�M�l=[M8pt�pBLR�EZ��cٴ�0���gH�(���`����3��j׀|�i�n�
���}B3_C��^xi��V�r.�ȣ3�q5�[���Nǹ�wV<E�V)h�~��{@���������r�8"�)�aݚ{/i��g�m �&q�y�"󣰽�)����L�������V���h����{��F����Z����T�3�u�Т-�G��Q�u]�g�m���C&x-�Q����:��u���&ߍ �M4(�>Og��C~XfQ�2do2�bo3㮾2e���H�g7�s]{Ĺ�
�E>g'n>��E!�L�|SF��|*i���}޿l%3����6��UK,�n�uQ�4�,�4tͩ�{=}��lЇ��7�(��)8�ux��:�����6�q4b�>�Н��:��#5��A�C��k!�[8 ����y�lgvs��8�S` ��ϛy�"󣰽�,�����L�aiÂ�6�Ewu�q�Zs�O�9.	ӧ�0	'ɑVS��4FnG�ldޔ�Y�0�L�>:��)��&r9�]�x�͐,F�O[��Tv_2�	�p�N �7p^��_<����	�~�o�֧'�_%�Y�ʖ�f�7����:��F���&r	I�D9I�3���x��c��+�;L_lv�̺���S����@,Q���`��r�X��
 �eQ${6j���r�d��1��E��_2y��5�����p�.�~GP�B�.�L��	jd�3n���
C��*��Q��e��ʾ�[7e�Z�SZ��8��qh�pb�K�c�.�1�	t,
.�څ���22��Ԯ.�i�GBf�5إD
��R�,kmr���Z��iI�e���@��kn�uZ�7f�d*7%"���̕6���D�MK�)dm&�i�-4�.B����	t��2�&1�H;b4���P��)A��M0���M�5m�-ծ�=���^�w�v]��}�Z�YG�ec�)z�tΘΰ�Ħ������֓V:�2��tM���2\z��.��E���\�^��< �]3�u;q�7:�ճ�[�F�!�y3��
L�u�����u�"��ѠA���M���7A��u��m��:h�#5�����h�iv���f��0� �dG�i ���uT�F	��Lvޘ���Ɯ̋�Wy�3�N �'
(�'BNoE,:��M��D\���!2#��nS�7��l�{��g �3D�<�����	�g"��8^j�d�r�nP����e�;+^�I���cw�y�x� ���.�ǎ��=��ۦ@��+��"�,A�P�M4"���Q�b�k����t�����\�C�>y����;���"I�A���{���^�1�/!a,�"�����c9�P �8pp�|��!'p���!��{�ٲ�l�rtf���(\��_���ޅ��]�{��ǀ�x�8�
V�ˆ�-�9�0����g�/{n.1�BC�U˺�=��[#�֕F�iDT�׺>0﫶|�����j��zwx�����8��k!�RcÒ�q�H1�+���~"��wX�Â�.A	8����wAx��.^��A�K��m�o���K	���\5�nL����Nu{��Ɋ����%o^ �n��gfi~�޼�Y���#�&��K]�|�ʢ��O��	;��g�	0r��n�5\Ny�fX?�v����pGQ��ΈnwY�ƭ���$�>)1�-���9����w�]ۧ YL�lb,��,1����&�]2A��\�nضn"�j�v��8�{�}=�}�� ��n�:��}���&�Zl=���kH-��k�>Ӯ�	0r�8 ��9&������<v��^9� u�f��z��u�����	���!'�n皽�/9��?��6��Bo8	8	0	0�Ou�b"v� ���uE�0��ˊycv�m.#�!���iϓ-�g�8����}��{;r s��bb+=�@/�������g���ƀR�hǾ����:����fs;|��1���%S9L��?��0mS��eN�'a����ȼg!&j����]9�7Ϝ����Y�6���II����u/��Ÿ.�Ѹ��c9�1��ݳ����ڢ吠gY��޷k�7v+�9Y�}a�<�9	0g �ᴚ����a��>�{.�-��F^�r�,��aT�,���maƤ�f�R`� p��pH�gO���	����>����i�~pj(fb�qβoOwAnxoh+X9�g�8�;�
L�y'gn�{wV���p��M�v�DO]�d���"1�§ Dc�"�r�9h8��������JL��
L�cœy�I�+�j��1�W��v��Sn�(�u�^0w�O�������a���ݖC���g]-��a�Q@��Ȭw���C�����n�j��d���v����7�/�k����&;\X��%���Ժ(Tz�iA(�Ö��N�AGo=��dp�w�{}���Z��<���ĢY�>���B)M4"eu�=��	���'���� ���Sg��kcg�"\Z�9��֮rp�;��.A�nR�>L�� ��4��l �wb��BQ�&:*1ͬ4��n+�ch��Mf,�6�{��o8�����|ɟ����g�|++��S���#��v���&�3�|��Y�Y�l�2�f�U�g�6ɭ��n	"��O��+����Rz	���9Ḃu3�v��Rk�ʻ=��-e � �q�3�A�`���I�H��A�qP�a��=x�љ��0�j�'z��d&�E�����D3��l̶əC�M刬x�����olc��;�� ��?�l��<�ՙ��>��L�VŖ��El툏h�n�?���^o]��-��[�p �����>P� �Ω��/�e4���Lz���������5?���RfÇ�]��zT��X�9c*ԗh�L椼��'p�31����ܖЭ�338����o��*$�����0-[;Q�֊�k_B?i��Us�|��>_��tҤ&,�X�c.��¥�u�u�J�X��C0\m&��b��R���E�f�rXjܵ-J��V�ہ��GP�b�+�&�f@���F��>M#g�W�9p1�
E�����v��2k3C#s�������p�Y�.�u�)f#Y��̕��f��cu^�Fh����F��]�Y�T�ͥ�l��j�0�</F��G����NӀ�
��Ć#st��eDL�*�D/f7)��p�Z��b��h��.��!�(��v�Q���Byot~˹����Nw�P����K���n���$��g"۸iNb5y��n�	Z�6�{6]�4wf8����u0iW�G�vL�:�|=�v�o=~���n�z�9��晜�f~N��Y�eN������Y�����>��Rg ��;y�M ����b�:r�8�wœ�s|�8nn�R���.�''88 Ű,�Z]�K����
7ݖ3���5�V�Bot߮���A��AKHst��]=������l+'��w�'+a탑v�j����mU!j��;�`8vf Cws��a�@0q�S1�F��Y� m	��������1	>��?�o=%����y�Cg47���k-L˹��s��7��$�I��7l+<���9�Ĵ?��h�IIzT1�%��������,��L��{ߊ�_�w~5���.�'�^zn�Vwb���u�|5�^u�G\&�f�m�ҡM4 � 	]Y�7Af|��o�r�o��f;Y8{Ϝ�8�p��|wü��<E���\�A+��D]��ݳ�]������k�u��%�"�2�,���@8�����&BLI���^��3 �p�"���$���1sujc+
�֖�x�3���Ǭ�/7��m��ߕd$��/D7�����\̤<I�r�^2���&�+�h��Id���&�q�`� ո	K��`��ohn��^囀	�܇�!�`x%���:Y�������^e4cm�^۔ôO!��~�����X�r�8 ߚ��u/�=����0�\�n��ZK���#���Ӯ6_��)�Qr.��+M��9��h:���qK����O51��/9��i���ȇ&�~�|����m�_�I���XIÚ(���L'�q�h��/�g�Əu}�p�=�'n��Y_`���v�;������x,���z�����+��}x����Խ��;i[�k�w�.����%����y1u������Q�,nL���Y{|}��f���2FP�j��L����2"��9�ýF?u��<�.b��,��7�&>en����2�#H�C���vy�g�'�4]�}X�6PM[��5o�);��Lc����3�05�}���p�un @6w�������aY�T}��pM��`�jk=h�Y��Q��X��{�g�z/-� �]!zDݾ��ߍ��糟�o/�#^��se.ha�{���%Ru�̤����]�3FBmɂ{'q΁_]�W3��8��n�����՜����>��7�,zձ6.[��k�v��w���q��y�mˬ}�����V#������������[��78���������q�m�y���������?�/x�
~Wg_b;&d5u��fh��n����NWb�|��;�8;�z��e\���4^I�X�g��L�|����bx�>��𛄋����D}�/[�Y��{|��^��W���@��A��?(��:�FVg��ӻ����ŋ=���Nwm�b�7���� ���G�W	�E����S�ۯOk���2j��Ľ�W�s��������֌��� ��㼯�7��)�1Z7���w ����s׮N+u
��@��#yc�gxf����G�O�|�0R��*��ĂY��a��-�#��w��ֺ���5����T�� TD�$�ʹlX�wQ��Q������i��Ƿ���۷nݻ|||<�r	�py*H� TBC���=��c�v��{�}�<v��nݻv���w�r����\�m��������w[�\3�w5E�w[�sh-�o����5{�Ɋ��8����Ѭi�nlb�Է�����F�ݱ�M����(�����<��Ǧ4�6�r�\�Ԩ���p�ѻ����DF�j年j-��F�*�EE�Tr� ��E���"�_����+�sP}+��W�t�K�橜����\��F�DZ"����f���xzA*yGC�[�%������e�U�	H"��i���Զ�zd8�C��pA)5��잾h�e�1^���q0NojÞw���V�����)8�BL��Q� ��(p�e�뎁����J�r:OS�R×�����#���~����g�؟/��O!���៭uWrJbSc��1]�Q7I�Ԯ�ҽf��1�Cg���0���$�BL5�R�\9KOf+�<���p�{�v_/X�ogs�U��|7N,�g�8GqX1Ug����q'�� �m��7%wC.u���|��9M�1�
����hz��
N3�]PpAG�]��y�"-Ҳ/�L��v�ɜr԰�漷;G��sY�̉>�g �8႒���藘&P3ol0b�84t��p�wu_�O/*�����5|��8}�$9�)�#&v�Ftf��� 7���T��y�2jR�R��� cϳ�iyiۏw���7{����0l��M�κ�b��[3�i������oxM4���a�n��{�zfg��	�����bYu?��:��,��][�ݎ�16ps��o7�)��)0pQE�I��DQ��7cV�K˹�Y��`�-1n�IV�m��s�Z�v�XQ%-�3��Q\s������6x��+�/T��	�KU�nt�s��xٝ2�E�=c6F�c�����`��pq3�Ro"�0 ���c���w1���K����+N�&y�s�p�88<�t�=^Ww��-1 ���a��.s�l'yAp�VG2�!�^tX`m`5��lzr.16ps�n�9
NQpA���4Cc�ȭ����A��d���X`#S��S"R�|ݝ2��Օ��P���pF�Z��ݦ�Gx�oYX�^`�;y&��ŋA��IC�'�*��U��;�&T�ca�Vpq$����pI����2	��~��~����w�f4���9vjڼ�ٛVD&��8Ux<M�=�'2|#}�m��2P��b����X�&/W�V&S_�֐)��뮫ڽ�7r^�tT�Hp$�d�Mq.bc���q�ZgqSK*��.�@��9��ZS'�c.1��M���R�«�4�^�-v��5�����9��eb�2�j`e��E�$�;u��K��0���kK.���r��L1�815c��f�剃I�V�k+��k��F�)�`�ݕ�����%��b�����mp���̦��Շ�~�/�~��6%q���йp��ZT�ŔYs�v#Pv���~��� A�g �l>I���W�����x�[�(^4ia����c!&���L�u?5=�&{[�z�qKU�nt�pw�y�R��r��:��RlK}�yټۺ��gUl#7�-�̷2����gy&�����F6s�7jv-�aNV6O^��k�\;�C2�٬�m�[�h��[o�$���]�2m���9�e� �g�Չ{�����1��� �0pF{�w {�������p18pBNR`� �'BO��#"�����7��y�݉���-~#������pE����y�)�p����,��-b׬Jmv!�W\1�ܘd#��k�����B]<��L�����F'�&!'ٕ{�ѭ
z����G�z�j�9yi�B�ˆ��L)̳�k��+P�몲'7�9�kW�4�j�j�#��*���r�[W���`����@�2y4y`;2Gz�V����)���N��j�0��}�����O}�$ߕդJp#��
�Oƀ)�����	��;�2��;ھh�Ȩ��Ѳ�A�`)7�aq}������#D�=��K��c!&�w�vޑ;Ӑј�u]���b����r�Kq�ǟ�&�;8oH�zM@���Dv�Q/���H�8ܓj`�S3�.A�p���ݜ����mg}+\`��v1duM�"�����5���I��a7���Ri�f��`p�V��S8R"��_DS�c��n� �ܰpA���L���GAȆ�[.(1��C3��4]v�Ȭq-Fe��k2��&ˡ��Mlf��|�8 �0r��$��=-B�u�������M��%���؇���T�pn�� ���i�9\�լԶ򝖍�b`��Y����c�����7�	���p�H��ј�sX�ps�I��&p|��a�{�S���W��W���C�ݝ�go��No4n�]�c�N�٘^�!��mK��-3��������������:�	�(SM(/>���x�������\�pE&
L��9�(�[�ʙ��N��Q��p�S{���bۯ��^U^`�{�n��C�]��B&��:�9�gɜ)3��9	G�@)0�x�����#F���wVfS憉��O��)�0�a�q�f�r7\?��h�����Չ3��HK�w{%�l�q�"�t �Х����ր�m\l;c(�h��>����%����8o0`Rg����k�.g������7��N��6����~7׷�Bwݖ��io�%��1�ATS"�MǦnF�"ӿ��[��r����^U^gRnt�:�O�I��$)��Oƣ<����o_0r.�?���0�w3}�C����I������9���+���K�F�)"�r�8 �~|莬��~h#�_4�JL��)�m7<�h�ȡ�N���7���DTYR�Z�g�Ⱥ6oL�w���Xs��{/��H�'^2�Ȫ�gwd���&���DKg������q��7�t��v�ii���τ�d�G�[�3;��(���0J�!}b�3�c�F��&��V.���S����I�M�O�72!�~i����K-)�v{:Z�gn!��mK ��!^�#4��]0-:hK�Ь�M5�c ��}����r��+_ȣ$�>�R�7�!�{+y�㧘G<�nK�)N����7mDv�9E��oQ����I�DIX�r�R�3�N��2ҳ#C���A��s�L_��(Qa�BL�����$�p"&���w�O�g�zlR�l�]^VNg$�}v�҈��?��g"�0���j7���0��4p��qw��*�=u��|��pL.Gf���{�g�[kq1�+�9�d!����5G���~��|v��)���=o	eY������`�R`�(��$�3�ѡ?�w?�?U+Zg^N	7?����S�{��1�V�=�]^����L�?{K	�v��2�[��(�V��f��2�P��e���N���Y+���iV�{�<��j���>�f�i��b4s����R��!��,���[v+�
��h�l\�CM�̷ ��Ux�Фs5e馎Ĳ���B�kq\��pZ9�Cj9����1�Pd�,�[t�"�&�ZM�;kq��(��v���c�D̺f0vfXE��7�Y��봭�5�%-K���*X�.UQ�δqt���܌�(9��
�AH6������nޝ{Gi���ʹ��������#1q����+fm3Y[J�Uӭ�tJ9�,�$�XB9�gV�+q[{c�9��uyY���zc��X��2lnŪ�t��I�>I��&7�*z��d;^�{���|8��r[��Ҥ�w��Ս�l�pH�g��!'<BE��0��Xi����X	��A)7�i ���]�G�2�]�;�U1��%�fF���Y��n��qL'p���[ND�A��w7�9Ñ��R`���nsu���+9&�A ݳ�0��-b���/�p}����nی`ُ�<o�[�<F^��c��X��z��*:����0������]����ʛ���K���� `�X�B�v�fs^�\�n+Y��5��13��Dl'�ǧ���6S�>���I��	�imm��;�YU�H��E�qr��n���ݲϼ�$e8l�����`"�gS�	�d5]�r�M�Y1�3��S�*r���E"ۅ�`<�������,7�B��Oz��5�roN0���kz��4�h�� �v��o��}��viߺ��e^b�M�v�Zޟ��۽M��|z�#q���`�$�`� ]�SK�������Wk�͍�UX�{�]����S�!'��i3�͐�5�ZV��L��o863v3�͌��ͬ��5�^\p�n>�`�!6u�������Ec��� ���A	8pBM⩮o+E�v{������mW^v�],�8�Jn�qn�[q�b`����bW?G�bZ�NЦ$�1Y`� �)��\�.��r Ԉ-aM �m���]>�5�0&1���`�Â�.I��^գ�G�UGV6��
B.�Ŗ1�+��h�檀!K�|�I�&px���oz�50�#<y�� �3�,�6z&��ӫ̉0�0>1,��@I�P�����y��<���XY	�[1�Y~����{����$[s�5��<�lD��g�d)����v�uh���v?5�<O��	I����sH�Ǥp/k�6l֞��@F;P{��y�Q��x����]6Vw��wȼY���M�r�-p`�:�	3�z[��:u� ��o7���N�*�ݦ�UQՍ���Î� �)��q��<<�]�[�a�]B32��G�{נݵ5�덉q2�9x�ڬ��5�*^dp�n�S���.�)8�츧ӻϝ�`"�lY�;�DG�0�]�l7a+��m �Q�hlcGF�Xe�P�=_<�����5���c�"��o���ѕ��1l�p!��7:�3���C���ޓI�����L�`��p��-�������U��n����l=�pN� 0X���D�Կ~;O�%�AI�����
L��[J�8�w�N�OQښͣ�28l7x�e��k�p �c��Fc��C�q�c(=�a�*���
N3���"O�X�FW��1^V�n�巿T�<�}�Rp�O�����(@�k������f��N�����t�."���+q�{�0���Q�=f�z��{x$ /g��hʳ��kz}c�y�~��(�Y3ʰBM���ρ	8��n��M�1���Ԇ�6�UGV6��8'e�z�L?��'�+��=ƹD A	�[e���q^�����֖���*���y\F.�LŻF���x�e����)3��I���e�٭�	����p#*���;=`�v�s���I�����8!oa޼�A��ݞ]��vv����@�⼮I�� ���!k�9J��e;��	ȰJ�^�L�7�k ���LRp���<o��,��jȪ��s����;,�@c�!'�J P�Ȝ��9�T�&rK�V����^VY����=�\p����`v�F�-�AZ;�͗X��BL��
-�NT��I���Ƣv���֠�B��^O$�A9l��t�&{`�폁F��;���fS������Q�o���5>9^��k�3���<��]��G#�O��9��3NpO�1� b�{�|E�63`�}契�����s�,���,�#�i��]~R���q2;N�S�ܻ��^) �Ẽ0���]��T�Ε��ay� . xk�x7�停՛$T����h�M��n����۝�$��L�i��v�� {;H�ޢy�mR�&y�OK�.�ń��V'q��������Y'A�k<�U�r�A^�8������c{�"�0(��6 x��-�������������_��)�L��L�X��G����(�W��/&kq���W�
N>�Sy�OKt�W�Эg8�$T��1b�FY�Ȓ��u��n�|�0�0�Oa^�;�8��v0�gv�d�lvח�\I7�US�Fζ��ak��V��B?~g|���WY�P!�O���Ӛ�)�q���sp�/�B�{D�ٽ����w`{���BH�h?zṷ��;O�??Of��3���\.&��Ƿ�'+�8ѻ�G_�;�7:���>Bc��=c<�e�A#�ε�O������[�����o�w�!���U�yNWЏ&5��j�͚f��<��N��Y�:�cɩ�wqf�������N��8�[��p��oW�z���Ea�9痻j�R���+�ǽ�ЯbλD{Wa�^�ZQ�.ceU$���T(����j�rԶ}gݪg�O��]�����F���n'� �3��z|	�	ߺp�����J1�;+����M^�i�Y� ;�%$	 N���~U��ľ��g�cc��	�\R�"GOoOonݻv��۷{�;��{���Ab�[\؂��nQ �$I!D�<x����n�|v�۷o����G*��Y ����W7�rLQh�*>5�*�o�uA��J��.�Űh(�h67ū�򻺊���ν+���4�cb���ݩ1d��Kk��������]��Q�{ޯ+E\�En�Z�N�m��r���y�,תnm��/<�5\�V�o/-��uo5ylk���U�ͫ�nkr��\�����ï�|��a<r��t-
]�[�a��i6Ua59u��%Gnf�2�6J�9,)�J�6*���U`-v%�:�P���fe0!L�^�R�V��y���
9�.l��".5ml���eԴ#u�k# ��6�!������˶��1v���G��WH�:M�Ɋ�(���6�9���k�!�e��U�j\�E�vѕ����D*���!\��4��L���28Q�f&��&Ֆ�B%��v�`J�W[��хs,�F3U������ݘ����[� ˦��Ze��ze��\��3,8͚�2�v���/�����&��	���	�n�6�l!��GlFi����A�.&��GTR�i�-bڥ��Jm�[�;G���Ŏ%l5����-�H3cl�ø	���ׂ�v�mcmj�����26�F�H˓JZ1���ծ�4Ԧ���z���6�˭H9
X��1�6��Q��ǃ��lڽ��&��Ү�ķ�M�8�q�%�8,M(vYt�ٸm�`�u���j̘I�-#���)�9�Ьs)��5%�J��X��Ύh�=�2�!�A�[P$[l��kG�XiZ���	�7i]�lI�2��u�V;Q���)�py]�_*պi����W�-�R�۲��&�XXf�jf�8Gb��p1����$^���X�v&�� ��E�։�K����F�4G���% �΍kb�,̱���fS�
����im����M(�i��ÖUa�ց��f�]�,;�`�Ѷ-��SB�`��h�Y��3G"�e���4-�-Z�J[�W2��@Inɶ�Eۥ�ceJ���{R�б�E�1���1Ĺq�,fmp�MqH,h��X�9���e�24���e7,ѪmmB�V�Јմ%��t2�
5�t����k�ѩ�]E�"�p�L�[h4�6�WBӛ�LZ���Φ�e +��
�͇2ܪe�-�� s� �0�iK����.޼��_1P���K�����j<�����f�y�}�?3�:�zA&c�3�G	/�.Ѱ����JbZQT����#z�CsZKخ��\iM��nF%�bƚ�����"I�Qfh�:��M��ec�[]eG�-6�!��e+c@���*��Q�l�2� �B�+����b�z�͵k2�ڸ��4v���j4a��&�*�k�#P��]EТ�6C�`	��خ������j�<��'����fe�,Gli���+���(LSF�P e�ՙ�y���fp�8Q�? �0�$Q���v��v��~F��\FCMn�Z�\��a�[�m�VBəV�3y�2���3v�{�3��A�g��m������+���8 ����1Ð�6̚���Y�%�i��^��NR�%&}�c�8��ͼj�.��rM�}1�� �7�� |�����A��͔��5.���8Q�ٸ�-�-\��w�{�#e���������p@"uÁ�>q&s�A�� ����MG0/��4(�|����v��)�*뽳�=,��&�Rp��3�s�Hh-G�:���B�u�`�a-kp#q6CC���!��-�t-kY5f��m�l�9���l����C��e�kPy�k|���M�w���Ke�L�1���&$��L�r6׊�LЪ���0陞!MS�d�Ru+���f3c�|b�eC����w+LS5i�m���̜��Q�ك=n�b�&r<�3���\}�3<D���Y�"~���F��<6g� ǋV?��*������g�+�[mk��$�鷺�Y3*�G�ou���f*~��ɂ��efUJ�l���p�\��8!'q!������o��)�8v;��2"�sn5���˷ʹ��8���^�፥��o��|u3��8 ���$�I�ȓ&��F���ڷ�W��'fa�������"������	?�A���u�5���94��Ⲱ� ̕��Fh:�mm(��4"��Z�M�#�������A3���Ր�I���ĳ�5;��0_use�T�m�n�����K���oe�pv�?���@;� 8=��aJ�X��3A�4cH\�qv�p:�2�u�4���]�u��A8��կ�&��w!轘�BAmoV����y�O�8 ��$�A$�`����z�T`�ѫ�����3mA�+wh����n�s}��.�b���yy�զԹ,w�����w_��;}���(��U��|"�o���`{�������D=un�zξY�TY$�[˶e�LʿYo����-i�խ�;���
L�����|/*W��OS"��v�x��戛V0�I�)0p)8pH�nԠ>d�m����UػP�:���8�M���A�k��L��ɀ��w��ϛ��=}K�~�����ff�l�e��aH�8�a�)+-�S����5����q�ݑ�'R`������{E�<C�U���I���Ͱ{���|AV����2!Ǘ��pA)3���r]ݩ��e��e3�}��U��.9m������SQ�$��61�W<q�MJ����Gs�M��if_l��m�VC�L�)�׹�@�[[�δ�}�¼O���`)3�� �L��0��9;�=���8�lcO�>IÅٔ��+���U���l��Ӥ˳�q8�Ǹ�D��w����74>׼�}�!��:���͑�M�^O�l�ns	���S�t��4L�FX�6E͌�Y��^4&���ުo���Z��A���i�3�>C�i�y����A�I����)4������<S�;�)�g�T[�Wm�����P\��FK�	3��	����ު1f�>��Kc0�m�kN�����ɵ�"򻩬�ش��n&��;�8����|��BN�%&�Y�wF�/���Τ���S��)S@0�s�H�g5�)�f��9��L�-����e�a��F&r
�:�g(ѕ����gx���:����ה��+�)� �ja7�oH)7	�d��`��$�{���r��&+�����`��;\8�l�n�8�R���I�vD��-p�n8
Lb���(8�p�:�q�'9X݃w!�|�A�g��� ^o[;�n�9�BM�.1>^����B�F(�ؼ~N�Ra��,�{)����&��ecÈ�h�^����><�b`��61�uT�U�N�`9ƹ헎䣸��s�t�
�3�Ѻ�������ox�sۃ~7�a(�����϶|=~{�q+WL\D���B]faASce�M�G붴3HD1
�E��P������U@�� 3j�
n�i��%�lq(s��b-f������J ��>���n1���!�V���Cb�u��c����zܭ�=�MH�H��іlf̴і�.i���3��f�҅���M)f�m\�2F�JM-c�Ѣ�^{}��/Z�����,��_Y�e��:hB�v�b�Z�-i��e#l�H�ࡀ�"�Ö�M� ��p}Ƀ���$�*wk"�T�v\<4����n�2���4+M]�B��!̫!2�9\�6�:�{��/��L5�Fc��}Z��s���N\u�³0j�����|a>&�+S��F��р�'�}�������
(�	0��_��u��t<�5Q�Mg���0\S�Q���7��Kd��۾m#�[8 ���{)�٪�yc�4�|ޝ`�Er:Z�[1�I�`�p;n;�]ӂl�pA�p�%�9�e/l>w��y�����aY�I�N��1�%&p&E�g��� ���97����⁕���k*�QL6�-��ى�]J�h��0^5� ��E$�v^��ʔʗJl;�+,�6��%B4VI�du8r7���!���i�ݳ�(^>;�^¿��.����zpZw�㓖��Cظ_�n��f()�To]wp,>�ý���z�7|�۱gyk��ğ�Zi��c�w�-O�b��Ƿ��(��u�5���-����������8nQf]/��c��_�!��ȭ�!9=��2��f[v����u��<a�1W�.�_��fjM�u3�E7�t��n��l9�{�R���9�х�>IÅ{k��U&�]7�;�W��2\����#{��`�F˿���� ����&f�ۗ�}d׷�L�tsqV*toS^Ep�1���@�[Y�A�q��7X�<���@`�0f	{j�֍v�Q �-�c�"�f�;`�a�"�!?=|��sc��NG���G<q��uf̸~�xљ�7�0������1��$�泟$�B)�O��Z/�t�M��dz����w�ꊪ]�;̹���'�Z��BS75�:���?���u���r
dC��t0 ݴ�/�$�%���*Y�N��lP�v�&���H/,r�Mh�3l�nL=(��C�L$^�U�I�-ȯ,z����V��[������T�a�-Sh��j:0���zX838(��$��IÆg,�>�x��
�6�tȇ����ݙq�M�љԛ� �g=��,ɑ��Lj��[iX�B(���G�q:�eSY�y��iÅw;ۛiR�/w�ppA�%���J�Cˋeݽt���}>w��>{�%�K.(���ap���s@�#�JcV�&�WF&̀��|���gΗ�z/K?�?�L�>I�UA�m�
�L���p%�k�f�v�N�D�N��$��BN�}}�[b�6'�D[��C���z���T	��g��L�tC����S:�믛�^jtY�g�vc���AE^`������x��$��w2����w�ppN>z��p�x�fD8)0#�wE�_[{�u7JL���g
�7W�s���`��������彚�R��]�9�|xgxA��(̛�Y��B���~�קy{�:,x��g�so��.mt/�٥�?F��juR�X��^Y�9,�9A��nL��Kg��4W���Ge*��穑3��~#�d�x��C��&JM����|�矇�Z�͍���*�&GM���ʕ��k��K.+Rʚ�F����[��2ܙ�p�jwoz��\ow�[��M��2�y�� �p����ȏ$�A&�pY:�2�r�cY� ���Nsw��EZ�\(��|���X��E�d�������.ym��NK�̲�fSyYȶ�͏�݋���Lf;�ukqg��pE!�L���2v~���&�_D�Md��}��`�!&.���u���8�2�����
��m{�tǲ4z���v�ќ�٭�l̫�̰̮\��s6��m����&^�������	�`���&��q*�T�ي��P���
�'��{j�\����S���L�f�yX@�}�M}�ᅯx��ΣE,^sn��'~ث+f����r~�׬��cy�{�����-����cQ�al��{Z˛�ѵ ���fh�u˦��0�FR6�ZB͈&v�`�#�[Qsn�c�[�Ђ;�e5��fYim��Όѭ�@��D��v�Z��(��]Vխu�9���e)r�6��crT�F\�?��y�<)���Y�ͳ*�j#���e%f�Ԍ+��������מ��US�M�����D��C��A�"��H�eŲ�ce��Q�e#��*�O��������)���˯����|έn"�*��s�^�8�A�ȩ�)0q^`��h�����=ۇjyw.��J�x����2\Z�%�48s���=ս�1�'���N���_�1���%&�c8�b����q}�k��Џ7��+8(���N��%sz���1�8��޺qW8o[Y��ݜ����3�[�A8��D��9��˜�'�ӌ� �ų�NR`'QF�9U����qÅ{7w�x!R��8�=���"����8L�ܕ0��������>������� ���l�ֳ��4�aH�0��B6	rMu33��f~�o�w�.����ɡ��?� ݶ%�o����tY��S�S;�qu����[�(�pAI�J\�.B�);v�a�:����A�*-�ND��W���8Ҽ�E�JTa��Ư����!��RA�o��1s���;��<�r�2
L%v$M{||}��>s��"/��{9��E>5�eZ�A;m��n!�I�9�ۀ�5Ff��T��o��<BMdY�����飚!�ڄ^��M�T]�a�{��ْ�V�	H"�p�'���k뚻������ǀA9��볜��
��w�͟d0��{1�Hܖ��Η����(��$��BW|#x�<���}8�C�b]�������uk{���  ������>)1hM[���!���������6h�K4��Tr^�155�M�䚑�Z�]5Q�Fx�{���ϳ��~u�M��f˃e��?�"��G$Y��{��q�e�u詉�|h�#S�!'ȇ&pG�g��Zp^vz5�x�)��}�ח�m��f[��E����������`6u�Tj���y�����3�!'D'���DPsg;�ӗI��J�����w��:-�}��d�����k}�hÞ
׶�w�g�\F�v܃�h������.
̛�y����Cfڗv{S��xƷ�K���;�=�ը̛^i�H촢��7h{��	���.{��3�Z�M��ɾ�B�\77�����F��^Əx�N����F�p�e�7͏U��h�­x^�$sTT���}�,��pYk�`>��g�o��?J<����}.�A�"�=wQouN����w�����KF����<X��Խ�]�O$&9fOf��V�*J�:�����S�9"��]������&�����zL�WǮ��/B�{u;�+�.\����w��G�_��������)��2w��^>po#��O�q��Xc�d��X���;8�����.e��Gf��z$����&��6*���78�J[���D�r��æۯ㽒Ϸ�d�MũqY��Fi/UR�(�.!WKg�0�e�K�q潕�+�!�����f���>���a3����վ��Jxu���d����Ѐ��]f/L��ٸw�:���Rj�����^ї��?�*&俟v�qxs3�Aa�P����,Q��@��P��[�T~��賵����9�{ozbt}�N������&m�.\_�\���hyܻC�~^>:���ջ���T���~>ʮ�Q=�Ir����>����(�Ɵ(2�@��j�Q Ç
���x�;�0 �'K�)�昐#,�'�����a���>�~�3`c-D�7���#��)�����>�����3~.����R+ٯ4j���qpR;zv����۷o�v������5F������j��ݪ��A��O��<v�ۏ�ݻv����
�9�*6�Qk��5�unb���F�knV��嫚�Ƚey��k�U͠AĉQ%��j7*)Q*-IGE�ͮ�g;w��[����y���h��QF��%��\�s���nF�^Q^[wuy��y�W9���<�:W�y�+t�k��Y���Y�{��a��c�n���y鸇�I��7�AҾ�Q�������|rg��.!'/�/n�B��_�k4\�.�w4J�����m�8oo��n��[Y
Mv�����A�۽���!����F�+�`N��c�\Rp�.C 
�\GE�1�}��^e�#�4��#a	pgL1��7-#Ci���8���%��B{7,�7����U�:��Ύ`��2�3�[�eYݘ���\��[�0���A[9m���u:o��k5wN����E�{��;�s�OZ
6��|�FOx�����lh����o��g���p�>)5 A�0s�v��N�y�=W���NnL�b�^fe܎k��+p�_����	8pk��S༤c.A�p����#�;w�����v�q�C�[�A �����6���*z�d1��Z����޹}�)�J��Ƽ#���{/wxL���^�U�(T����Sp���ԧ	=�> 9Dp9L�V��7`M�>��w��_)S���훜
�8,n�Y�(�pA�ÀE'�̂Y羚�۬�-B�u�`@,ͻ/Yq�rET@DVgn�̳;Jd��5�;��Md�A�C��8 ��y�v�/9�	{���#���f[GN��5�6�W0�Q��!&�aw��.��2�b5�*��>��o�{1�qv�q�����x�g���>��^`�ݘO;�:h��D��\�SYe�ɒ�I�*��a��d��jjx*�P౻տ[$�ԲS);��a�wL+�oWM��q��y����gf
1�t�u�e�n�ٙ�G5��e��������Yް��PY�9�O�9Z,����}v�$ ��YY�d�qR�qs}{9�Ë��ˌ�[�~>k�8��z��o9�l�u�I��Oˎ�C-VCI����`��}�>��� ������)���Voc㈝��,�Sk���W�{.hi����*�\炬QE�6{||@�6߼O�i�~V,J��P��c[ժ4m�k��nמ�X�G:؎��V�)X�&� s�J]#^5��K�3�j"6�H�5��2�zۚ�6K�e�,���GM�\Ѵݞ�����4(l�-�]��� L�3�YH�b;&0�:�)HX&���x*��[j�3A*l��
ԔG���
2[WhE���m�+�R�rU|=yIm7����vk-�P�ZL�q[,�ŋj�(����KBS&�t!��i����`�bp࢏�az����U�֓����Zui����]����)�Rg ����Г��>Q��h ��q�{K7�5��f>Sp�\��rX9
�8(��|l����հ.�pn�����6x�B!��);�"���w�J/^�z�#��`��2�3�[�A<�� �'� v�sv�E8���-���C��'t�pAI���\dn:�x�M�{a��%��Lh}�J;�np��RgRg �ȇ�I����q�.�`����%w�K���[d�5���`�^8pl�r�q��&�uN��d)0��<�nqvc(ȫ��R�4ƙ�U�v��*�T(=~M��nO>bpo"�C.����-��q�խ���02�!K��r�L���`|R`��T�fOjN���D�{znK��n5�x�*�KFN|�n޸
3V���	6�_G�%V�W��}��z�=����-&��0�`�r2�g>=�.u<q8�|��8�f�z�Ñ�(��#.��5���I�C��$�JL�u;S��t^���kyW�r[���	�`�o�Q�BLR��y�󕷯�\�6\C�����q�������X�9ӭ��Sz2Ҿ���Z"�K8#<J��m�_c]����C[�&N�=�ټ��o�����N+��罕:q8����(�}Z��	7�ɑ�պw��<������x:��c�r�b-cm�u�Mn��!.���K6U�GC\��g���_p�??}ٹ�q�m�7l�7um��2��O+���r�����2��4p�'������f�9O��9j60����5��w������*��Νn��3�}M�?��'l~�l��z�4Y�ga�`A�`'� �����$�tP9�Z;�7Ea�z�~�%�{���4gy����5n-�4�;Na(M��������X<��7<ǂ��_�r\��8}�t@�eR瓍/�N�=��&�W���0�Ķ�>�>»�/����%ȭ`�$�"�pRglf��;L��5ݷ���C��n	��1u�e_^4��|������M�۱.��8\�7\9	;��g ��Aq�5�c�#m�� �0~��W���VMc�gN�	�g�?����9I�V�.�$���X�16���9f��QX9wV��n�`E#��N�@�7��\������v�9�\8!&pBLs'!��z����z-�2�2�p��բ9������p� ��|RjЙ��|�����*�S�f��na�3l�I�}ܬ�,�_^4���pNKQ��,���h��r4^]͈�xӢ�9n�pI�����L��<ߙc��l�ev�F�UddgN�|z�� ְq�9��|���E����+�_��`�W3��/͉�l��r�x#ދ����[� �F��:qhhT�E3�6��ޯ����s�����=�h����臇�&2�xT������잚���;�T��3�s��ѸuU���{��X���ז�st\�g ����9I�����s�	X��hb��æ�u3W�l'��w��>�p�"�8 �'�V�Sϛ�
%���Kߌ�#�"�.@lH�qQד�����Rj��Ƥ�p|Fk8 �8pBLL'.��p��3�q}:��7����6�A��&r��5U�ls-�2�!���w����U��wx�$����p���)���#�{��Bg �8	8�pܣ1=��y7���L$�`G����(�6�(jbI
�����ve����;,�{��.��x�ۇ"�Å='I1VK�N�x�?�{|Ř��&wܖ>�3w���:����lu+�d����v�jr��	�ձ̲�3(��\;ʯ@�ӑ$�#�?��p�nO)���#�{�8 �L�\��	;�������<�lA_�0;a���Wi�7����x�s��CjģRM�	*,˷>�f�l�w�r"���(/�Ծo.�J�F�ަW�_bo *�zORf�=~>> |]f���k/|O�,�d����e�%WF)r蚚'V&*@�Wm4֗,1W25lu��L��C5�v�,���4�]��ڇ<��0�Жk�텻fD�4��ٳ(in����fB����ă1.zÌLi�%���XR�)p��3/�6���w:�p�.�pS+������Mli�f��\���P���1���7eeU}���Ʊ������D��H8�"lh;n ��.�f��b�q�̦֚���i�|��7���r�a7l<�ݷ.��]ċ���y;���P��bX�����^ �Â3��p���8 ��ӹ%���l��1�z�h"q���0yW}����7S9�ç��pA:�9I��\�<�P �g<ޜ����^0>��@	7�М(�a�3�=�OtF�Sj$���E����[�C:����&e9��l�g4m6���;�6�� ���W��=��)�̷�ޭ��x�A����&dI�`��pAn��8	6s	��Â3"&����>;���V��Q���|Μn �M����9����W-�����|����s�2��0��[���hm��1U�1*	�K).l�ڀ�#	��{�ݾ�`���Gk�l���?^N缮i,7;���82Y���jz�GShe��������d���k�r7�����c�J���n�S�i��s3gY���yA�ʧ'�x;|�9[]�0�{g��T�gީw����h�w*sQ&��֖�{!Top�����-��kU�����5ٙ07ռ���7n�����A8�K-;��+Μ8/�� 8��4�8�	0^0&*V-[1�E��3�o��[Ʉ\�;�}8�x�u3�Mky&Ɓd�7���o��bs0M���� ����K�}8a���k��(|�����'�&���p����&gRg����I�F���x�խ�.��͸���"{W�K �pI�Rq���63)�>\�G1fgv�]���sa�1�mM���Z�VP��t�kKw}���-�}<����D'�RaJ�QY��"�q�3g��Me;���o[y���5JL�$��&�`�d�b΅L�he�����<`5;����3�ry�!S8 �8r)^��=~�S�N7��<�嵙ρ �g>I���y�I��lgJ��5[w�0���i�ogҿb�� $�{{=����	ȧ��F��2��f%]j��͹5T�U��1%I?s�vp�L����=���xo��;P�k�eS�y7ڸ��޼�$�)8pBL��a��úၩ���Â;�?�&)_m���as���8�&��X�:�;���L,ų�~`����'$���� �s�c39���N��Bh��l�#�����Z ��A��E�>!�I���Z�^������W8cp��(
j��q�aT��
��lJrUtv��}�ն��?�5�)���9��r3�[2�뼈�L2�Rfe{��'8#1�Rpa ����Ƒ��Ǳ��[E Fc��A�`����כ��"��:q����.`��Lӻ�]ƺ���;.	�`'I��|��Ҕc?y��[(�fV��#F����T�Es����I���9�Ywi�E�"	�o��&p�k2���*��Ȁ}����a�'�O��H~!X�3i�xh�k2��KD��D{��'Y�=(�ʗ/��&��3��i�{��Pt��7���}]�η�A��J�>C��d<��2�!	3����!%N���o�g����$�k��<E�Μnu3�Mkqsvޣv|�Ǭ�٭VX�<z��&]����a4����cI��)(�-Y�ΩB�`	fZͤq��Sk��y�0�ÑI���:��L��G��v�� �;u�)�ۻ���A.�O��R`�&����]�,c<�-�x�q�q]��i�l�u�LN�=,�3
L�+y�e�X���'�m��I����?�I�]+c���0�dz!V�V����1yӍ��Q�8>���L� �LRk��bՋ!����g$���R.��[9��d=��u��V^�n�/�d9���P�WP�2�&�Lg����61�m�i�[�l��Y�l�r����pA�`��&�a#�#g4���H?���r�:F�qv�D�<��{Q��1'!>�������Y���"0�'��-'A����M��,���ua�-iJ+L3�i`�D)[�+�m�a����jؼ}8qL{�xp��� qjl�E�
��&���q�"�<��;�q7�q�	�:��|��~��2y����{�7w�ۼ��������V�v�ʷ3_��ׁ��ר�����E�<kq彇VV����Ny�%6�c����Y���Ǹ�y�帇�7s}�c�Gb�}�B+���Ǌy}���e�o��۝ ��˕o��KS��3܂�����s�^�Jp�$�O�Ō�{lj�FT�ɶhRwݣ;��{�.���{�qp�C�҃M5�w�\r����ثQ���@�rg��M���E��{��Gw�=��b��ޏ<�[���������qM����a�W�z�XX}7����ԙ3������~!�akL�y�=꽽wN5F�OG���^��E�HU'7����3D��-��ʞr٩�˷w��� y�ޚ_e��2��S��Ǻg���ӡ@�rgj��C=rcP~���MKیVWI牎!냖��dE2)Z8�>-����W�\D�g�y�;<|�6�݋}}��'���^=�M��ruV!s��@��zt��C��\Lw��F�u)6���ѹ:3�,X�w�{������,��%��Ϛ\`U]gyz?tЈ��{��(�r4zz��\S��~_=ů|1��	]�O�x�wyY�|�����3�@0�N�OG}K�w���4Uj5�AD�5sDW�֋%�U�j�q�����nݻv��۷o������,��j�~�lPHJ��h�o�����<v�۷�v��eRy*HIʩD�n�db�w-�',������+˘�+�.���4P�D7ӐQ�/wE�(|�r�5��J"7��6e+�"4i�r���|\�w����Ov4>:���IQ����h����^Q�\���/uĖMy���������[�I��i��1I��ͣ�vPe$|\+�pY>wV#����F �I1a `e�#�B�t&��pk!RE������}W\ђM��a��d���"��	��~~�z�g�/]R*��ɂ���t��c����ؐcTj����3t93y��T��ݭPBf!v�6WE�l�G�/�4�X�j���K	k��i���ja�(:���,�e��Ŧ\�+y�8���/�r���2�.��8n�3YM4+�k-*��R�x�*5�z]*U��4���|{�[�0S���%��Q2�	�v�Z@͖9���8�`�\m�+ZL(�J�+�͚�-�1c"�6[5�W�
K6�B.s��7S�����T�-�ţK�#`ʍ�����`-���ƙ5k���u)[v��J�R�kȍ��Q�lУH�7i�|�R缁�j�Bf��mʇi�n&�˂aeà�h踛#z��j�(щ��5��kQ �:mD����\�P��)���Y����1s@�ڡ��4�*��5�ԫA���I�I�c8��,�%��Pb65fmB�le���@1`.�V��h����L��g7�2n]�s�1�v�.!�]��sJ;�v���F����(�n�TT��=k���]c��a�P�+��٭&7t��&�+HgV�]�ƹ�Z�fn%͎LV�K�s�`�+�3k��,�)6�55�X�f��p]�����cU��^P���ae]��>D�b5s4���M��Ie�j��&�!N%�l8&е�5#��[�17Z��m�j��1,bb���4+@�mMC�Ը�̋��ݡ�j��Z��W!����[��d	�k���Q�bf� ��	�ZX�I����lͪ1+b�vk*&�:��[֜Q*���@��.	[��+n�Q�jLQ�juq��5LٹEl�ơ]mbKx�!6V5��vi�c��!���e[*��fE�铬f�z��5��k�Wc�],��f��p�֠�(�iA�1�-6!ؖ�A.k�	���mX��� X�6B�!� f�����ֹV��8b��iP��Q���.����)`̜��/T^�t�$?1IF��^���u�UOT/�䙷9&(����2��.��5�6#\����-m]�Q�R�k��.�ܡ4�*�2�d�A�����Ɨ�Ѩl�p94�lִt1�@ͳ��L�8IH�b6�f���nf!P�qC���S:6�JL�TҮ��,un�NuĩjM,Ĭ:��ɕ�k�&���5)@��[Ļ��ʭ4V��֎m�m�$^�;�!6�MzU��K꺢��S�vt�� -K,0��
�	�^���6Қ����}���B���8rp� �l�,��sxf�g�A�-U����&!���oP3����
L��0r�W�x�Oe���|G]����L��y��gܢ���ݐ�Á��ys�9y�ͶܻD�����q����A ���L�y�Ml1�Ų{���[U�����yP;՜���,��,��sEe��2�=�Ki���ֵ��ko�#i�լ�n�8[��/6�;4^���)��]�����x޳�;���9R�`v�Ȼk�ь��4�2qS�T�(���7d5����`�$�r�k�wE��냖O-����@���,%����]�ة�b&��Ⱥ٦��-�n�,���p����n�W�3*�)3�Y9ר�-s�^)p��p��n.V��~Y��p�-g$�o�8$$�i�6����?3<�M1�hP�Vn;�N��ப��f�"_��m��s����~��Q����-�nM��F蝣7]��2�y���i`�y.r{��|���a�E?���+�ks)h�f��7�8�'S8>�½�����h�x3%M�h��p�������p��$�A�Oᯃu��P�Z�h�k�7d5�z E[8)`�����1I���y�!wh�ܦ��9��v�A)5e�Vq���I^Z���y�f3^EB�m�D�y�p�!&I��$��K��k��D��̥����%�:q���
�pA&pA)6��.i�7�_���?~!��faCB���[�^��i�+vo1��z�U�ԓG�S͔Bk�-�fU̙�#n�(����������u��5m|0]��8���p�$��L��&���Zi���g�S �V���n������E���8�����=� ������Ty�R�>�%��AI�a���:��ZiiǮ�)��S
v!�VC��~��Tw���ϻ��?�o��݌�����ë;�W~�5�����^s;���跋pt䌚�"�h�z�vqAN�M�<|��� `��˽�z���_3g��,�g �㉼�I��%.Vv�kj����|:_��E�y�p���Y�(�77�H����r6.���ׁ]�A����o$�RdA�I������i6�j�����7���2��Y�Fs�%����	3�G�0I�ٶ2�`�`#$O�O��tB�ۓ&���$e0%575�l�b�b�T�Mk��i���2�ÿ8Yy�Y	�XfSҙ�����=L׊_3��k�%/�>�;�+�27WL�!�.�L��a���*74����E�A��W�A��Qc�G0�p��	����7ˠAp)�z�_$����Hvr#�k�������)3�-�I��i�/hE�{�'�C�M,�á��rX?�>�p࢏�a ��8��O}�s0�pA�����2!�e�ټKGaOi�1�V7A�g��C������7?p���\�rʷQi�%�ff��2��Z6�E���i�;i���|Fꬬ{�W}n>���n	�:}H�
��y^�Ɗ�ӹ���{��
N�n�Ǹ���'[����ݠױ�\��6�5���0>.� .�i�&��سy9�3�tA����R�R����p���Ņ�Rdзn��e%��U&�/T'oq�n�[Y��I�z몾��ɊY�����0���8�ɫ����"iì{:} f8��
(���;���X/�bw��7㖬�Ĵ.	��ucq��>Ƴ�Q�)Z;�4����W���f�0 �0p�(��I�5;��I���.��a·}��x6\�)@��L��i�!Ҍ���vu+�T�Aoc��\�A&V�U��<>K���x9��9,�?I��Wb�.A�p�$�	E��^`T�E;n��@�ssr/��ڧ/�[�&s�C� �1�8 ��n��[��[�s�Cz-���6^ڳ�kG��&����X�N�{qI��槛�:} ���9�|�=n��ަ�q��f�����	Թ~P˭B�R�c�ݵ�]_&d�/����|1�gy 8 �{*��X�MjS3U�ʐ�T��jS:�1�b�h����Vj\�q����Ri��VP�S�LVLasH7R]f63���n�*�H�2�,�ӝ5�[e�.
.Թ���\���<�Uq5�@�r�B���A�������6h`4fiq�-	K/=i+j"]2R\T��Ĺ;J���lj���F#�U����|��>S�^�n쩹A�ePQ) XFJ��I����d�GGJ����;E�mR�?��z�R���f!��w�FHI��_ew��a��Ƶ�������va.\�IÂw�L����H&����A��s���������{�#%һ�ns�������0r�6��-��LXط鏌�GK���p�y����`��{!�T��\/\4�^�n�mc�F>�i�m�T��)w0���
C��f�oi�>!&�[���הh�x�ql��A2�9Ϩ�ܙ}��es*i\U��FS���>k���gv�BM�)4�K�|V�Gs�M9�9ל�.��-�>79,B��&AI�Vgu�}|�?d��{;�t՛Y��Ȗ$Pͷl�+Q�uDYK02�ہ0e�Rg�	�=�����_�n/� �)?�e�ǅ�{���L���T�6.�>�Y����A���������G�.�@o0��*��P�rC;o�/��7Iy|������$Q*LO�`2��at����7����p6�ž��^w�M��ˢ����ČW�De����p�'�[הh�x�qm��S �8r��Rн�ޠvY϶��	7�� ݳ�M�s.kK���M�#�r�u�2U����vX9���n��p����[����ul;
����ټ��ُ�x�X/{�^g�V���K9�R�<�ֳDU�h�!7��	0	0�Ů��l���k�����Gn8q��{ײh�x�6��a��`W?����	?�]����Z�����<�JC#�
��l�$��Ev��ѥ�Kcq3ui[T	ti^��|�}�C��]!�M'�5,���w�e5sy/��zO�;y�>�0�^,����z�8 ���!'pJ(�d�J�΋���4";�N��������19}z�A���&
M,��P^9��<޴�K{ϮH7r�y�=Q�-۶��Z�@�r�L�q�o��}�uD��)�_�:YW������z�Kc��;����@�"�CHm��*�Z#��1�s�(��^��]�l�=�+7��y�Jg"���� �	��I�$(7��M���sm�������pA)3�S;���t�4��_���9,��J/,m���F��L�8pBN�BL�$��H�NC�1Hè'��g��Gc����."fr����U��:�<`��)gt"h^�o��@!��$�Rxb�qf�U�X���Hl˱7^4�щ�I1��
��Xz��[״[g�Yʷ�)��/���Z#}]�7��nݸ����,07_��
M��Rg!�}���b/ƹ��=������
v�=�o��&����0����Nܞ��ڠ�P`��gaݷ�n\8"1�-3�`����JL:��n�J�m~�X3u���s5������8�a[z�>*��w����#�����C��a���/@g"텧�̓V�������K8%2���O���LJt�����aB����G��lc�z �}A��7P:Dw�Dբ{���>Ń��Ů�S���{��F�]պ�F��I�h<�b��G�C'�lfyNe&��� 
M�{��=Us�G��)���4�lr��2\���������#�ÀQE�����63y}A�CG�͂Pc �,���h�GE�Cdb��Eu�u�1��q������5����ҙ��Y�;B�.jc3��&��޶��A������Rf�	0	0
͘[����?7	J.A��s�0A��I��op �6|��K�v3�r�vN7�)����cy�"�� ��`�rܪ�@��*�C�TV*��s�s�����(�M(��	L/j����ޓE0d�v���!Ū���GxQS�����޹�SY�c�����pq7���� ݰv��m&���A�k���k4�o7��8>"m�Z��I����}����g'���5M�[B�����rjɈ�8��q��K�Zu��(��ꡚ�Pԓd�]1˼l�2�D@��V�}��*n7^��|}�o�䫟��Z�Op���LB� sq]�]M�0.�����tB�J��3���)��el6؂��j�1�E����al4[KEc�B�'2�ηn�q;hw5�m��*�Vgb56�Qw�%�3p�0aۮ����fc�V��2��3v%r���$��nL��6l]k������c%���̥��/Y�ʶ�TKR���G[ŀ�)�m�gk�g�"��e �9'��<B��U�o[���#b-f��]fօ�Y�qU0����Xl�|}�����0�a7xό�v�o3]���+���cތ`�M��d�K�,���tl�M��]3�(�Sn���w�8	3�5�X��o�yg����?�7�K+#����:�����|u0r�w���'w�2���¾�8�ՙt��{;��˞rA�U�A�5�H7��ץ��{�!ߔY���L̢ɬ���&� �n�=�oG��;��<��Rg򉞽/��ԣ2��g8 �pF��g��P��#e���7p࿘]��X^{�W\l�Ǚ���1��ݛ��GG��o/�Z��	�`:�H&pA�I�������,��߅%��%j0��,�k4`s)����mY�e�&�ۂ1ƥ���O������?�F�p�]���ۇ
V�ǖ�<;���6x8V�{_�ɱ��A�'F'�)3�gŊM��EN�u���5�#l^�ڝ�۩*��:�lk�����y�/S�R�x�C2ȬP:��q���Ll�-l3�h�k��,}2C��<�>���<x�ޤ�+o�x__�z:�N]ޜa�e��AnMN�l6ƪ� ;�w�mC����^�p3)�@7l`9�\[���=�p���.fη��3�4�3��g>�oY��?��X�w�aL݆A�p�����=B����g��m��n�@k`��z�޵��&Tz�@�o�7���@)3���$�ʲ�C����L4�����<�9yYD��A�ÔQpBL9�^f���]���x��:��13�����0�q�Jڱ*Ö�{[p��D��},�s���C2���&�r�n]�=�����egF�2s6�a�}�ʭ���=�&eY�e��Oh��I�e	8p��"���]���˼�b1��!��F�x���B]{nDh�+��c�����^+�_!�P�7I��i���Yn�~��R���:�<�a�We����o�=�RD{����g�D���{��,�e�_j~o-ʗF-������ow�6y�ʉ_�a���ՙĹ'�Y���c���7���m>��^�Eɬa�y����������_�����V�&o�_��k��O�W��9���#�DY�vO^H�������������|�r�7�%�dXu��V��M&vU;� Ϫ��,�霪�E�nv)�w
�[����b�^y�9S����5��|&�j���h�ۻ�.L�w������hȰ�T�1\�E�<��zBt�f���}#I�[��4�Q4��z��.��8lz���϶{|vC�gI�`����y鷴�Wa��}����� a}�YG�T��O�%�YW�7h����]������/��_;�X3~���������/���b�87��G�7nhk���ޛ�g����"����8r�l�3d���];����������֎4M�FF��z3���"km���<dܣ�ۚ[�l�!\E���S��O���7�#�-��dY�l<W.ą� �v�bX�yr��zذÞ2�F��0�	�Og!����5�8	>x%������.a�+o���C�t�����l`���(�{�S��]z��,+���`[l�g�N�{�z.�;T��s�,O�?��X�hB�n��˞Ӟ�$OL��^�����l�.�A1�u(��.�rd�^t���.�=�wޤ��3��yq��> ��|�������=A�Q�ԓ���tN�W�(>�%�#>����)�����NY�(��_N�n�g��홲d��]DP��q��۷�ݻv��nݾ>>Itݚ�ȉ��IPD0�˺�~{��Q[�����ǎݻv��۷o���2W�\�?4�R،�nFb)� �I�$�8�v��E��u!)ɜ�yv�8a�d_;\Q?N�������Q2������5�\�T1 �S(L���	���u���MD�h�3�i'���,�%�ӊ0����$�I�+�p��J�PLͤ�&I�6��|�iH�33��>�]2I�޵ۉ��$$�$��C$Th���A�LhA
II.�ȇ�Q���B$(�8�fi�r�Q��LR0>Ed��yY�^s]_��\�W�N[��A������L�t��A���xǙ?�U]>]`ކg9�gF���pE0'k������Dp9�M �S��!&�5�i��t(XA[�}����w����c��88&����p��-��ݍx���)(gg����K��Yc�R�&G���5.��p�����uʶ�(�r�2�i4�ٌ�x~~��̦(Wc�_7cC�K�zi��-�ݰ�ݸXݝ���_rqj��n�og9�[怩�|Q���h݁�.��ݼ��{�v�v��{�����c�_��*]�ޢ1����ְ	/?�O䞟9����"�V��p� �����7��Lz��Xx�l�0���<�M���d{܈�q��#�8��з��U�b�+��7��3�~���āx��� I1s�֪��t�VY��H�8H�����a$F@����!%{��׾�S�w�v�I�K�\U����:�ݷ�3Y[����­�B��Έl۬�뗉������-�-���Gl	-�1.]YC��MHH�F)�41pL�|���(U�dy��5]K�q���76\4��!��&��MC��&[���@�o]�S�� �:����u��b���G6���Pi��{i�k �����թ�v?��x�ۀ���P%�M���C��bAQpf�7��}ֹ���퇵Nd�Ɋ���:�i�
�l0��	7�:�U��G^��=�N8�9c&lt�!��-Ԥy&��4OuE�ⳕ)�&9�;v2$m��e��ڏ?��Ε��zz!C�j!�v�I�ܑ��Sm���n���յ��e�6<Nhq�S��]��9�#C��'ٶ�� ���^��+�i|ݹ5۵��jX<M<��Ǿ�Hy��üfCHf�`�dk�4��ۣ��1�]��m��`y��Ȼ�-�h�U̵�ͬХf�51�]6aJ";hl�BK��e\��V��AW]3l	�%�beq��6-R͒�+(�����[
�К�h]h��bz��Ѝ��<�[�i�S�L�cD���<m[�wd��.�m��B�`iu̬���������})ǆ<�����U1X���6�!�v�-ݲX�����cZ�C�Z��ܿ�2LKU[F��成����yŢ���j�� =WZq��I�I?��x�92��4pMާu��9�������m�׍Ϝ*-d��GcS��q��}>m����m����}`��I19Yg�F�]fPj��m7�s
I�J��4��2�;�W��}��r�l�ܾx�x*��ꦗ��m\��{˧��������.�J�e[�e���u���Fm�׍Ϝ=���0�K�5CS�7�5]�/ĵm�X��P�!�ښib�5�P���`,�ڋE]�ĉ���ˁ�oI�I���[��:o*�n��
���L����Cxmۀ�PV�9޸};h�C�b����D��v\HWX���/r癠�f�	��5�~k�c�y#��UO=K'�kGS��0/���_�0���j?>@�i�0$I�{�-�W�r��a�
�;��N��DTF��\�f�vj�ځ��I%#��eL��`8�IuK+��E���9�:�&$�0�s�BN0�g�bDY˯]���ns�мW��v_�����=�M�zx�;��7��pl�aR�鐢e»�Q��)����s�5^rǻav*�
��c��ߞ�,/���14u�m ��k����[��.-�6h��X�K1w0Av�2+ܞ�6���䓄��q�57�S:�2��ΙǞ�jy[~�a��N7�o�]ߧk���З�w!Ҷ5���^��yv�����m��Y�m!�l�Y���ձ�%Qo���u�t�D�*��o�Y�СAۡ�M�Po����1ck�/V�JU�s1W��@צ�m��8���1ӹ�{:MC��G���<�;��vS]���s�	�X���$��)YǑ��2ٖ�&��v���L�`Ս��6����q���:9��˳����I�M��$��UH��u�ȑ�}S��6�^U��{/����)�[��*G�^�?}ι
L���`�Lܰ�C�6Ƙ����U�4�"� 1b�cH�~��+$$��_j�=�Mv+���M5OyI�r��ԗ��'�LY�:c;7�n�ۍy��
޺ ^��x�������I�s3�fLd�}v�I:M�;5�'��V%Z�rh�U��yg��&�31���&�3H� �2�Q�F7��n<�>m^gvM��5؜��U^׹8E�_XFI���_"�a�����'�S�P�.<6\/xG��������W��t��\��Y6�j�2b�v��`�bms��x��o!ܛ�#v�G�����]���NM��y%���rk���驨��7%������]ǯ�lIo'yN��F��&�r��
Dq�سkCld��m&�i+(
k�M�f%�z�.ï�$�I�Ml����9k,��,��ĭj�
�`O0{N`����Rh����@<0�ޫ̞��ܴ�'�7 9c�$�����O��Z`#ԟ�B$���G5�je�=.�S��ܖ3����Pb[7v��v��4w1�/��!��O���&N�;a��g&r�c��-�3p<0�F(�X�N.ҏ$��&	`�N�E�vjO5���=Z����Yy�U0X�����������
y��Aѓ$E�z}3�񁭻�.�Гϸ�.|;���$&�9�{'y�H�2N��0�i �^��Jo c���B1f���+s��j\&�K��^�J6��R�֎ ���V�n�*���=�L܈�`8n-�f�fi@�Nh�v�vʫ3��B�N��U�e!�Z���k&�c��hx�M5��E��mn �L&
��L��%0�-��F�c�Vkb��k��鱙��`Z�]�Kn��ڮ(\�;�lF���F���B�@��I�a���Z��l���|��?CSmZC&�],u�U�Kh���3h�J�%vm$�+�w�.1믽ؘNL37)��_`v�3��ßWLU�7����d��ڹ�F��R����cow0m/[;a��g&Vb'��l��:I�QL�4t�`���o$�&�1��2�U4�
�$�[�U�-�N��i���M�$�RR읭w�>6ިa�o�nv�R�w�ې�vO<�y5۬��LW��i�x��(`�(�]���v�y�t��fwح����'���`��O䣻�O<��������q>�$̴�j��6fb�v��hMj�WB��frb3<0!�����O����+��r�0݉��E�ZQ������I�'@�w�Ұ���%Y8HpX�ں�%=�wߴ���/�^u$0c}v���]&�~S�ӨF�x�`�٭A4:Ñ3T�$jk�� ��rA�������i(�q����d�x�+V���V��{�;���K.��w֙ⷆ�i�X' ����zs�� ��I�J��X�y�j��=]� ���W��UnC^^hI0w�U<�J���+IJLd��cW c�3;MZ�g�1�\vOQ6� X�]��h��C���￾�v��9t\�\5��˫�[%66L܅oRS$��K�wh��aX�us��������:�������J��][y�La)���{��T�C��u��r݃7wY�)n�
����v����r����Q���$�@H��k���,�;\���<@�{�y�^��(��⼺�O���ˇpD����OZ��gOý�!�ߩ�_��,iѭQ�:h3#4������ ���|@���tn�q�����t����5($��l��6�[v���}����p�&Q�����X�u�e0�\�0�EKȭ}�z��d���N���SQl:�K����̬!��/6�ᴇ���mY $Hnb
s5���/0�,D����ke��kkBmib�[f�*4��s4g��v�,���'I����QǴ>;\t_{e�.�3�궟,P2qޫ�m���-��^��u[1�m����ڦ�D���{s���^�|�3rY�-ޱ6֛�s^����v��wz����w��W�iyy�M7jJG�d��'�-9�e�����pa�x*Fk�v��k���q�������f,�tOLTvTDۉ���[P	wv��y�4��^�=��7<���y<srM�~x�}��-}f�x�8<���ڼ0��O$�p��n�kJ�I�`�p��u�!��4<�h��ܧQ����{r=�M�>{�]�y�Xbit�.u�H�������Q:�0�n���n��SC�6	�8z;V�����h���I�I8�����щ[��a.ئ�Iř��.׮M�I�#�͚H�:�+�`��{�M�8JM5�;C��E��-��d��n�ӊ��=�n8�`�t���WF�t�$u]Z���d󷍀��r�� ��I�a�E�n��m��y%;w��W���yy��U�p_f�ln��$�$��7�Q���7��\�\=7�	��JFh�/q�|ſ�@J<����}�nq_;
5x�`�ƾ���O�2�i�֏���,�7�����:��o55{���<W'�~��4�Y�Ё$<��:��n���~R�m��j��#���uw�<\��
�8</Ī��]uk>�Z�sx��������T8�x�>�oh����.�]O�r(j]v� ����K{ǟ��x�ӽ7��^H��x#G����W:'M�{5�V���'����,�y�c���h�8^�'1ü�������;яo�{�0W����}�7���Γun�Mh�axe�:���&���ٞ��{u���s(�4nnp�i��b&-�|w=�*&����c�W�k��j��X������{���@j�ۛ�g�dOaE�� ����-���},�@�/ϰOu= ��(�#:<�m{Gw�~��'�(����}���³���Җ���زO_	��_i�|��l�:�h�/O r1�o���!(���%����D��=�t�OyÆL��=��Y�A����ٝG��|A����L���-�Kn�̘{�3o�wi�}V���wke�J��Hά�:=�
�駟��t\�F>��͙����um��n�oA���� T��$��[3T���B�մ2m��ڀ������V�![4M��}��Y����-_z-��ms��4�0m�h�}�V�,�Z�y�v��nI]Y`�`��'/e���k��Q��Ҙ������� �pj��Ч�w��1'���t��Q]l2|�x���,���	 HC�a���22�_�!�1�
�fdFIT�����n8�=�}}|i�U�w30�31�ˣ$�% �#!��������q�x����$�&I$@�d`f��fA��XB�dE�"�1�f"��?o�� iI�uuЄf�4J�쌢��5�߯W�Č�H�L1��}�
�0�#6&�d��A%$dd���&��E9ȁ�����LI�)L!{�g�W33fF���H
IIP$�/8���ܙ�%���&nvOu�$�`2�� ��!+�H�{�!��0��!j�p�L�їWo<AI��/�ן��q��f�Y�y����r���Ȟ��ja9,�r���6���c��G�U� \d��r�
�9�h��[M�j���eI����KB<Uq�u�F�38��/Y�+[ĉ�I0V˘4fc5fU��e�Rp�K��������.��K���x��d״����a�����2�*↕j̀L��l��T���(1Z+1�[+�Wc�2��hC7�Dю�ؙ�8%Q�	ei�*�bGWi`)�i�� �� Vֵ��1�X�� J�)
\i���\��LE�UfՑɥ�Zl%�e͔�*�P�֬�漛J��va��掶-q�IiNS��KcqH���\���˴YջX�%h�2��m�]0���Rƫ��5Sj�q�[WS�0.1�KZ��1m�.(��b�l�s������`&U^��sB�E �u�n�^��q0G]�;8ЈMH��eյ��q�2�Jm�P&�&�X�Y��UVhҼ��,���5r�Z�Zح�ғm�Ve�F��.�]x��WC0���/@f��U\腙����j��pT hс�n��i��8uHk"�{n6�0:��2iKq��X��a\FF �������a64�,#�Ae3�csd��1w	�ژ�k�c�
�B�b��������3�4D�1t�%f�̸��Q�c���e�C�k���El.�f[:�È�B������ښ���t���լ�U9���R(��4#6!(Lj�	1�u�:��M]sR��3�f:���[�R(�Ѹ�uX��k)HK&+�GM\\�%	�1�ii�a	�&�m��QS�ZL�
C;-n	kk�Ǐ����S.�a	T53WY��َ4�[�l�v�fZ&WW9��V��Gcd��4���U&n#�޽���J�����k��49�=�M2����K�Iu���2݌]`�hƨ\�Wgj��P.%�6�3n�]��x�0%�X�����]�|N�-���niv^f��8���"k6��5ќ�,Ia3�hmS��E6�.#a�,Q�a���99�Y�4���]-�)im u���%
�l.4A�m5v��؁1 mtuK������LXT���f]A%k1s\.�(Ֆ���:Ķ�U{;:�q����iA�R����%&J�bWg���Ѫ �9cR��]�]���R�YJ�1�.�.�l�L�]H�%#mf[�?�����+m��w��on#�(��ma!SF�eC3D�"l�J^X��b]�c���O_˞$.���w	7�M�j��j�e;x�j�vVSz�Ճ�������s�~���]���5�>���s{�Uz1]�������?���g`_h��lX��d���\��OSM��=*t�A�����m�C.#�pO����?n��t��֏��'�~�O��k����̣o�]�r�9�~���Q`lk�n���:�0�$�F"˸ʖ����nouM�˻-7�����p�%a�W�~��"�ڿ�?5�)7s���%�8�Eܔ#5�PW]�!J.Էi�qK�����~��\y�$��D.)�GpAdG2�!;���?��� $���0I����{�����r{ ~�?@�羐��?���,@Z�ouX}�׷��8]1s���?8?9��*�~7��~2�]���lulΩa�P�������0���+:����m�99����n��g���uSC�y�syָI��y%6���8 1�r��7j��x2�[M���m�ܟ�0	7�������p�\�"�����G���P�S�Y̸y���NU�}$�g�]�w$�n�]�ݣ��X�٩��wsMp���Q�[ynOmpd��\�!(í�_�v���g�	2TؕѴ�#[H�Գ0��r��1�<b�x�`�3���@�Oׯ���̥��7���
���Q�s��hjo �y%p����h��q��W�%{J{Q����o��Ke��Yz��Ǐ^8|o$��뷯����Ai�^Y�v�;��u��f��0q��,���h%Ι��x�C��=�@ݧڏ����Aj�c���> _�4]���2�o-�ݮ1�7�N��ۅ��V��c�v7n{��Y���=Q{��k��
��w[��	�8���ˍRŋa�F6�y$�&���%����L�c�#l�e����iN�<�fm�yո�.������}"v��~{�a��t��]�j�JV�d���.���(�e0G1`�!�;�t�/���Ld�fw��T��9˅EF��� ������}������p}wxOs�30��ݹ�{�ދZ� �o/8
��N|�#�K�N�+m�f�-��`.�)��lA�<O�ٷ�!��fu�m�+�ܸ���#�'S䛺y�͔�s�=�}wYEa���Kq13���-��*cͲ���Y�j�z+�.	����6�;Ea�3W�4ͩ�s�UO>KpA<���.]��߬-��oN�Cf7K�{�z���ü||w�����L�-��E���O1P��]����tZ�qJi���i���:FcȆ��̘!��רr�=|�?`�5�`�ĵ�+-�D�!���9��V!�hc�-A.a�P@�]�;Xm��I����z�v�7:ܵ�sM��t�iǓš���!���S ������+����w_u���wn~��}ݡ�L�Ei�S�
��$�l{��og�f`��b�n�%�N0ŏ��$�Ih`��z�g�7�l���-N	�O7���M�p� �yRph����]��)��wU��۵y�4�g����\<\6�������L�]ۀ��������>6�FRkS�
�ւ{W��9��u`��6 �l����n�/�@��~�����	j�H�s��`���̮�������&�|�Cv��u���mq�D��0�|}S���h��{4pS����s�Jf���:f�Z�B��<D�+���xK(j_#���2TI�[��֚��[�h
V:j�cHQ�&��2�5�p]R]Ÿ�Q�XAa�!H��hqhӬ�1q5��(�Ac���M����
�@cJ���J�eN %t��chX!�qHDطl�J톒����\�T�sM���BL� ���7�
e�2O���,[�4�͘��]n53BJ�[�dˮ+�E7���r�c�o�|�?��]��ws����7䪋����٧{��Ǳ>�x]��M�
Z�s�J�̻����V��a��,3�l�tɭ�`��8���ت�29�lP���_��H�awo�^ ���Lqul��Y�&+�j��J�ڻe���$�I�LU�M�)���2V@I8����~���/;ټ54f�3�'�uR�	'�I�I�VoLE��R�y����ݛ�*5�{����%�oEBcW9l���i����]�[��X��� X�[�k��bU��.���1�d��՞�1Г�둽֢�;����Q����v��$ޟ$�t��i�~m�/�$��U4Ab��4�|����X���FgNxl�ydC�Cd�ٔS�iRr��'��g����W���П:|A�u[���[�T�_�C�)�;���>�������#��]wt���/N�'��Gg��䰝�ɾآ�Y��я|�I�I:LF朚�ٟ����cx[\*=�Z5&W�F�^L�m��s9�>������z���|d�3�v��@��s�xS��ӽ<��C��f^pL;����!�.QB�����Xo�P����aP�[q���@*�-�Wf��@1��n�sKÖ,�Y����Ǳ�O�I�1��M�t�l"�Z��x�*�ʗw�|nh���m䓌����6ғ$���N7����҇r��I��ڻ�-�֒oD���1l��꣢��ęoM���p�PJ��)����C�Gc�
�7e[�ɒ�N3�csk9�)��6(4�o'\���Q�E؛��>�U�6."��Y�f]ڋ��wx� >��������kD=]d�����N� �I�Q�E*�E���HZ�cn[�*��V���ز���1[�woL��Q373޻a��H�I���Bj�yw�Y��okOO�ҙ+�#�w�[�lNQ�S1���Hu���m���J�sA�R��[*�X���5���DPulu���`��3�"�S�M�
)��+�ޞt���b��WYl�C����f8�a�w���T)��H�c�W�-�⻽�ۄ����YU��I��NTg>٠���/���L^z%�nc�0��No%�&�$mrX3�t9#4�o!�j���`�$�$�JKC��̺mx�'�Y��G:[�u���ܛ�j.o)�kjj,e���Z�+�ñ���e���A�R�)>���ny;�U���w��ҁyV�M0��6�.����<|�R-�{ߧ���ff�x���Y^�d���I�Im�ݥ�v�dnR�'�:odZ�f���si���\��Ǎ~���FY����9�RPR�*8̖f�Su�9!]�R8�l��?������k��J�(C8(�:��dv.��M�0�"�j�2�G�`�$�]��s;f�m��o�w���lSE�b�ۆ�N��,E�9��ཱུ����k�	'�I��+����q^3vF��|U�˺1t��$�%]�a�UE>�'a��ژ �P�huӬ��$u_�����o��ltӀ�n��w�����K���csZ 7��z��a^�s.���Y��@�`�{��|��[?hN��a�~��/#��/4�}j��^��{�{s:7����iN�i�#���;������hL�.&��v'�p�`+ll�l�41b噟����S� �}�2L~���ȩK�,���Z2*�Z,Ja7V[���֑��g\�1�M�6�mE�H�LbZ,�@Ɔ2�.�Ʀ&,�5�cN�1�Ս��%�c ake)Q��kq��)��j8$CD�CH@���b�6[��[/�UPv�6���p��j̑(��k�����0�]�IR�)b�f�J�@2�қ6K����������۷�� �n&�
��D���Qs��m�nm�n�7�D3C,�D4!��K�7��IҪ~ˮf����V�*�-V+ߙ��s�o]��$�0>����hv��+�'Xz�SlZ�z��]�P��K{��G�3T��4�L+�b�v����zR�%_�U\�zDv��%�M
���X�uk�ޤ���|��SC���ċ��Q|��v��5���m���q��f��(W-���I�oy$�a�GT�>�,�s�v��pwr���I��o{��I��+�/M������}��>_�1�N��R���A�*�< ��#J��_�m�A����������Q�b��^XFe��F�_����wH	6z��]����A�w�f�%9y��Ӵ7�uw�C�W���M-���}wW��۽Ŀ��*��,&OR�_�s5r�NX5��x��<�ވ��[
�͵�ϭӴ��c��;%�~�qv�N!�jj�O6��$��7�xH�B��^�Y�{����y�'��d��oy$����޻�EEj2�k�_%��X<�P�]�n\�r�K(�,ˁy��fn5�ĵ���=|�f5y�&�LB[sx����L��m��mU�Vc����˛�&�I
C8?�"�'�]�YHl�/8u{9��M��ŰR̊ ��2ۮ�1c�y���"|��G7_%>	IǤsry��3$��4�F޷����jNJ�&qfy���۰6��mM�q�4���^]拌�}ɝ-Z�n�̈���v�ьM䓏% o�������0�R��p��<����G����V�{���4�9!�p��ۯ�s!�����������׋��o�dgzVͽ�߫���y:��O��Mne�!a��s��|n�^�惚Ǔ�G���}�h�>�o�y�>��|E�}�1c[��c|=�>۝�� [�F	Y���/	Ş���"y�w{����@,w��}<*�{�ɂ^h܅��D�x''��y7��L��z֗�r��w�z+P��`燑�Ϥ~yV�޼�4C�a�d��&"��%�&�2k1��&l`���M��㣚:����3��DG��_&�O9��{�y���x�=��=�ޛ�zwO��!���P���i�`{�.��u&S6�c��Φ�ΝH�}�Ѵ"��)��l�{��i�Ex����9LE�=7"��F����}�W�}Aܔ������VCy���Y��HNH��g���d��.�y�m~3�8�=�&��/`x ��}p�h[gw\~��;�r�������\0^�hG�+�U(�]������<��5�'c�X�o^V�6㞲��Ws��{?hڏA���
��"�����E�>��*����r/zԫr��+�Od�+������Z��h4��/�����N��78�;����(���͋Beu����8����P�gL��s�7ޮ�1L�٣���E�k��G6���g
޽#�:��h�^?-�|c��X�
�:�,*��yðw�uGc_���s����Y?N8� @!!!؆2%!�$S�!�B${v������q��<}xy"HHI!#$��T�Ebe���+��b���������q��x���_��]�9�"lP&�?}Ԥ����$����1D��ڂ`�%"`L�b
�w$6d�&d��1	%��(�Rd�u�w\�0@���$DAR�w�]F����X ,�a����X,��d�h�JDD.�p7�\��4d��fD�Pa�E��i4QhfJ,��l`��a��3Q&�
"7�t�PEI�L�Q��bd���}.Q)
IHD�$A��:��^�ל�O��YY���tc�sy&$��2͗�ȷ'�����k �S?R=�Mӌ�3$�\ �m�ȖǤ��jqI%>	2Ph5[]���nG^i�)m���͸aڒ���x<�%kE���	
��ǈu/5ɳΊ�6ʐT�5�ښV6�L���T4ŸХ�?}[�&�췻���z�N��1~Ϊת̇��cXB������ݻ�$�&�lA[t�v7]����ަy���+��e��%��$�����'Q>��� ��I�`P:�U�r���T휂��j�Yy�6��.�z�N8�nGn2e7�����WO�G�\��v9�Ȟ�Uo����,Z)t�C1ɧH(��_(Ơ��[Q�sX+!|-�c
�����YR����I��i���Q]:��yW��������N�֏�B`�L�$�(��WL��e�q����+���w�Xn0I8�][��o��ћ!6ۇ0E��-��Ek1s����+����ձ֑ƍ"��"2�2�^�k�𻷫Sy��	��jˬ���n���H�{� W>�I)&�b��dU���{u�2�������\O�{ǽ��̑!��;�N�Ḧ���[z��$�g\��.����'�bsԸd��IHH��\��7�5��'�P,;������y�K)�՗Y���aWn�u��XL�W�\�J|� `��qO�q�w��nz���=�.��O�6�@	+atj<?6��բ7�fc��>�Wa�a���W{��l�4����{�3sF���}{�/�NQ�>�L���[��&p��ˋ�����u9f����)�JK�{��;������}y��$d�i�2�qD5��tMj`�Ŷ�b�.�)�IGk�XJ����l(ı�F]��6ua��e̳���m���0�	/��A\E�[�a�Ձ�XK]m%�M�$؍�].��2[0r<��b��&t�3�n�Mr�`34�ƌsR1�H4.&��љ�*ˣt��F4��N3`����zۈ�X�6h�z��׿O�^z>��lo�2�A2��f���r9�U��t�ɡ4BZ�AK1c�0�b~�'�M��,�˟g�f��19�Ze`���(e5� ��^��I��NI�T��fu��v���ᖢ�y�K)�5�Y��H ��S��v��`7G8�M��'��֩���+-�2��/�����" $�R;*��e�
�6�۷��$��8��z6k/ �ˆS/G>���{7F<[�|}�w���2U�{B�66X9ip��^utK)�3�Y��,7�����flSlu������粇�k�ȥT��m]�!��c�c�J�X�h��<94��ro��+�[_��$��$�����<+���5���}�nx啰^ ��&��`�T�.�	�-m<��{���y�c���Sê������8k_j�K�C�9v�8�YǗ��s��.���|��w�Ԥ�K8�w���ɯ����Z��5���4����p�h����8�_���֥�v�]�����7K�v$DJ�ؖ��g.�3FK{9?�`���6��ۤ9����V���A�;�fb䳐��
紈˚��ب�'���X�H-�&&�I:Uw��L�&��5�ky�j:k33i����0�)!�>���}�/}��IE7Z�i�p�m*��gW�����,5���r"wc�V�����.`��	.3w���-��������9��^	�cx$�'�M���?#~IZg��N�"����}��4�+�!��Up��sy.�B�ýMu�a����$���k�=��&	y��P#r������a�I��1���J�CYb�pMJ����2u�F�u,�f��v:L�=_g,��yyE��7o�}6�i�+���T5�A���edw����h̷��٫����+���I?�`�����v;�[~�o��[U�k�A��������ٓ
��+}��&�$��&	0	'lF��i6�r�;����rr#�5�b��[]������Fj�������~�o��]l�(M���͘��L�5 +�F�+��f��]K�sL�y���C�7y���w��c�Td�����t���������t�f�	��>	2I)�a!B�ƒ�M5ո֫���/��Y��,;S��QS��%���e�U��I&�J&2DK��$�����w��q��Uï\W=ݸ���a�ݝ.������䨴���ٵ����y;�R/|�2��sW��̋w�N�d���z����o�Ԍ*=<���WǏ���(Do�3hFna=���!,u&�i�I{�̐I>ow�����8�o$�$�y$��ê�C]��wA�����d�7�RM�U�O�ڊ����=O��qa4���S*B�sf���V���]��WB`׌��a�1m�����$�Bm]}{���f8�ɪ�U���i�4z���kx$��0�L������;w��ϓ0�y����Ř1�\Sxn�K�3���t��'6n<�X��r�	%	)c�ڲ9�vg��%&�/��Y����ϩ�K�Xn��Ƈ8-��P��L=0�N�o^�u�-ѻ�5�j��\N6?>�w���xػ�u��0�$�2������Vϵ|���j��ǎ��6�f�I�Jΰ��I�*�d��mc��c��0���#)�ݗC�=.F6ķz��/9����o�G��>����J�&F�#�|>q���c>��H?�%��L5�R0�a�r�ծ��q�.��.][��2�ڭ�%��K�s��gq���%�[����-
\4�Fi�"jV Eq`4^F�n&m����F�رh�V綱V�.�M�B�3B\���bY��Y����KYJ���3ZJ0�ԡ�s5c��:jڬ�����f��e�p��ښj,�,��VT���4�-�]6�v�����vK�M�����~~i��q��s�	�1XV�7Y���w]R����b"�O��)��!&Rq8�u��4�&2�H�w}U[��*u���L�cy$���npM�E��כ��5�+�r�sw�ܡ��~K���${K«{������wn`��¥�G`X�y�`{���:k���5y�I��l��q)@�]Hk��l I?T+�m�;d�Z̽��f��|�=!-��î�]��N�NfD��@�aIy;Gh|�������$���ט��3����ɪ὎=Z�4�&x��z)
��!ó�3Ao8�(�X��Ě[eJ�]e͏Z��)C��0y<���}���&�R[�ak��l���UB��f�[y/"w��%���E��c�����C�g睗ڢ�/fe(�W�zD[�V��iZ��r0mkr��J���T��+����~jG���Y��q�����OFI�G�����~|iV�r����c///n�؅���D�/c� ��U8�``�p@��5b�0��n���������ݓ�`�I��$�ђ5z����{�>^���:x̼#�뫘�[�Uu����s���=\�]޽d�JM��M�`ctX��|'�t�^o?46V1�����?_��ӟn�kj�����q	E���m0]ц� v^���ˋ6:�܄^�t�o�~������2I�I���r��4�F�ӓ~�L:E�w%MW�w@�a�$ޔ��7�m��З�V��ykz��u�z�{I�ǎ�����`���.~�^'*���|�7N�n��Z��0i.�A���Syq�#��X]�IV]64����)�ۧq��]�4X��w�xkcԜqs��x�|�j�,�׊�/���޸aڟ�0�����X�T��:�����$ֵ�;;t�ti��.7ظ=�v���-8�Q́��Z����I�I��>^OYL���n��N��k̈�T+�6�fc��c�:拚�XG�D;3xs���i��[�:�l$�%&�طe�4;l�Me~��������,eIĽm�oF���/w���ƨ����_8��O�I�'�I�����3u�����˳w��t?8��r}޾8C��^���)��G�U�oOp'ȧ	0	H�*�Kt�܌ګa���Z�96�[2�xG7��z��]ב�ڍAi�~^�]y�0��u�����(��Z������X"���z�難��н����n��2�6c=E\<eʘ���i�fXA���l��_<ܺ���o����w��ww����JE&I�IkȌ�vd,a�������ޜ����Z�&	(YL��+WI$�E��b"��f��,�^��*�q��Cm��\��U��ŕ|�I���n\��&�W���)����M�:����JRo��{3$��qd"-�z��漽u�ol���/w���}հbD�a4i�Ezwr�{Sy$�����\�ݮ�f��h+u��x{�V� $�}v�㘭n�t�W�d��%��i�]J�cc��ƨ�q�iL�����&��	2]�}����]6�^n;F����o3�s�e����O�����j��PUQZ��/�������$@DA_�
,�Q��z;�
S1��G,�K-�ͶY��UK5��l��VV�*���eT�U,��+e��f�YU+5Rʩf�YU,��ke��e�Y��*�f�Y��V���el��Y��ke��f�Vm��T�[,��*���f�Y��ke��Y��j��l�j�UK5��Բ�Y[,���Գ[,�K*��l�UA��c�*P�1R �ie�����e�e��ʹ�m,�Jͬ�m,��m��Yf�YVY��j�*�ʹ�m,��m��ifڃ`����o���Q`�`�Q`�`�B���Q`�`�Q`�`�z�hTX0AX1TX1X1X1X1X1X0X0[��� �E�E�E���E��E�F�E����UU� �1X0QX1X1Z�B���lɖ�ٓ-��&m��eUS&[m�)�[l�m��2֪d�UWvݙS-Z�mTɛVY��Z̙�L�*�mK-���^���,��V���gƶ�5Rʩel��Y��in��E�`�E�5�ͪY��UK6����E}}������*������Ӱ���=���|�����/��������_�xO��~I_���������~�TW�?X~������E^��TV�����"�O����>�և�UE�~?�}��^� �w����!7�+�����Q'��Q"�) ��"
� �,��AJ�
Ȁ�"(���� �b��`�`��"(���F
����b(�X�,D�
�*,�
� �T���XSm�R��J�R�����[J��U4�M��fV $E�T ՟�BP����S��Z֭��[Ej��QmV}�W�?w�}�_����������� ������?)�}_���	�:M�����?k���? UQ_�C�'�����pU�Q_��h}���TP��?�����������a��#a���zO�l�>�@hU�Z���'������xm$?Fy����O�5��?�B'�~A�0��TW��~���H
�+���(��
	�_�	g���E��x����L�:UEzN䑉�~��K@�!�n�XV���s���E_�t���}@Q@V�����:��
C�O�����)���w}W�,�8(���1}\                                        ,    t                  �       >�    4��*�* D�BRTH�J U�P�!TH"$(%D��R���)%E��)BQ)(��G���T�UU$�@U�'��� ����B�;� a*����@��v�Uw���)ݎ�PwH�;�n�����    ��� }� �(+��� �()x�� � <��'AB�9 h8� ��Ή�F���-eP��(�稠�c�lw��-��������]    ��>JP�"( RI���o|���yʑRݞ�	R��R���e"Qo%!^��Q�]�O[j��PB�vt�
�{״��("��+���[��@   �Ҿ��*�}�z�J��x=IOw�*s��J�pzj�\�z�wCބ�uGw�‶{��M��޸@9h    |>A*��J�UJ� �;ϐ��ͅ=�� �ww){^MPoUH�z��{t/g#�S{�J����RR�I,�%U�    | �Uﳠ͊�	Qn�����@.m�{r s�w ݺ 9 	�]�     ��  \�*EH)Q
P�*AJ�E^}Pww �5\�]�� �v: �wP��MC�SU�t n܀   �  �}�J	w�F�IT秡[��jR��ҨJ��j
�h�D=��������T/K��=$n��*    ��  �EPE"�EUR%$�
ﾆ�{���R����@wgB��)7(�W@��!J�,���@�9ȅ\�����    �  .�=��P���PF�*����8��
y�N5���=R6w�=+�UKޠ=9;� ��U��;���T�	�*�� hh�顒R� ���ʩ)�J   l� JJF# FOT����M� 43PI�RoD���� ����~��o���_+�'��W��כ������MO�� @��r�/�p$�mV�����Z���j�Z�}uVI ���p�˿����/+�����U�c�B�2Z6��F;"��"t�-��Bd���/!7��z��̙�կ��lJ�+*��T0D�^�-Б�O$�]��f�cn��ۛsK�^�I��[A�Q�M:��Q8�&��&VЕ�1f�X�Tk&�� ��������Q�.��\����&U�{.�8leK;��l�k)�1��qҡ���X���U9R�⼕�E㭊����׸3/
��A��T�g�w,�X�*�W�Eڼ���^����֍=�[�v�o3%Je��9��ڕ��/K����֮de�;�u�NJ��qd%�Z6��+6��fm���T��aU4P`�F-��cRZ%e�JnU�w��guR���]��L�hyy�!9��n��j	�7cŕu���uYT�LH��/[��2^�4�E�{5����I]<�m�AG�VC�8��x�5e�lY2�2�������n��QR�ʼ��e��L�,K�����X.�mԲ�N�^�+V�n�2����Un�,dĨ�q�bElb��[�b�lř�����{6��fúp�j�BQ�"r��YUwջ.����3v�ީ�9��d�Hn"��Mk]��z���Ԡ�H��A�W��\:Ҍ;���1�k0�f�86���1,l�<�N�e*O32���&8Zuy��302�CYҌU�-ͰY"Bl]���Bf��uiY��Nlr�Z�f}Pn|&�[0
պ��Y���OtRxUE�ZX?-W��j��U��omlZ�4��7ov��3a�����Q�fڛO.£S�7Dn�'u��M�����%���T$j..������v���������[B���[�p暺�H˪v5�����n���+���F���؍�wGl3��6Mu�I��2`U������f�kj���Fj���1^$��f�)
�Fەr��˫	�)��bV�Pw[U���[�Kf�x�$��z�*�6��Ri�v0亣��[B���'���m��[ŵ\@�/n%�fe�̐^�ɍ�uP�r
�ɗ���V;YY���ww���l:�#����L�<�����{h�yT�ɵS�I�鱖��&�����Ĳ��,���pho�:ûwzoEe�h^JY�f���ޥ�k%�f��bV���B��\Z�]oqR�	C,�(M^U����1���w���-�mݤ�^�[M@R�ůun�IG-�5R�+E&NCR���$��X0��{Z)ڡXEU��1��,؛NT̻kw4�[�TFA����m�J�w�=f�]��U�i)�-�V��6�V+7���4�R��nV��%,�Uغ��^�	�ɇV�*Ss-�'ʦ�^bGMT��ҫ	X
�XsVeɘ �;�2�Ku��vm"r�GU�wxUaZ~�ڣGm��v)�R;�oj��!,6���m�tj�l�[.���m��iGv��1$��5{�&��"�jx3E����oE	�UnN]��L�m;�;7I2��6�F��[�V+�uy��v1��(ݝ���:���kܽ�e^J���`Y�s6��J�n��Q*��շ���Utd�gs��mEy�(��w�*�gs]=���0�5DQ���7heKw�e˳5ܽ�c)Z$jR�Anث�c,VV=�s��_c�1z�i��S�A�{T"��yx�qL�^�n�6��D4�ٽ�?M������e�&T;��4ڡ�΃�T����Mn\��Y�:p[$�{q�r"��rJ�7�U�M�s-i�JUv�r���4$Y�UR*��L��e�r�$&��vMU��H�9N�;�&�P��W���k"��Ժ�W���˫�q����44E{j��1��Ɯ9�z�;:E12���b̴�X�,�[YA�N�b�B�Ԫ
��F�X�q#�U�M�)A{v��P��S�;��d���B��e�4���8����̬.���q����u��V]-����Z̵�)���X�a�X�J��5����ۦ*͒�֝�Tj��yt{�̼�.\�9N���,����q�eV"�n�1I3�W��e]�z7a;"�`4)�{v���il��u�˭���`�{�r�

�{yEU��,m#cR#�0�܍fC�isf܀ջ)"���Q6#;�_e�M�w����76��{�n�%@/���Te����Ƴ,��8��{�Aۦ��4�d��o�G/
x���v��k+�i�30嵮�O%]6���Ŭ:7`�e��ek�F�G*�-�nܻ�TP�N�j&��IK���֒*����:vM�.�H[{�.���!䭛��B��7jE�7k+pi�5t�Տkd�US-X�	ùT�]�2:;��t�i�jʺ��Ub�aݺwJ���3n�J�\OQI�$R�]e���+hCm�Z+N�5Q�˼��NVQ�:WK${G�%`f��Cn�P3e���9�)a�e���(#+lA/a�XFn]}gu��Y#6�;�E�1���*�aR�:�*��Wzv[���p�Al�Yv�Q��*�ee0�UK^*0aZ5Pv
ٚ�ܚz�r��J������A�͔E���(ՠ��P"������M.��Cv,XF4��6B�}S0��a�T���Q�5Tt�N�QJ)���#wUm��L��Y��T0]նa8�7z$-�6ka)T�K��vd/	y����{#V�i-$�%a9D�Yn���2�`r���%�J,抈em��7�9��42�u�B��*;GXei�{Y���sA�"/No+&�����9��� �ȑ+YA���8�m�-��Ɯ���Ia�\2�EV]@��f���B��F]��]=�Fi�&��̡%��U��j�?���5s)����P+��w���z��r�;i^(�ɑ��z,V��J����ͩ�p1&�7S�$V�Gw%�h=�'ss-B�޹��0l$��oӪ�.޻��"�mKղ������ڣ��;QV�w��5/,ӑ��`�u4]30ͼ�Nc��U�#v��[�kr�&	�,j���\�wS3V�U/a�V͜gj�1E��i�ɗ���A�\*S�4]sS��2�l�f�:*�wQ�X��T���Bn��5��`_ �l[�v�+.b�F��Fl�E��V����c�.�[F�����1&U뵺�ں46h�T�e��f�*e`�>�[�-A�J�K��6qfm�FBܹ� ��3X�@���3s\���&��p]��K$f�0wr����^�+�1ؽ��lƹ-�{e�Q�X�l!�.�]f����u���3h�����F��K�f����4���+$��{+H��l� �D�Yf�X�ѬT��1h���؎�����IsU�	�ph�)&��(Ëok1i��e��`�J��o/L�-S;B���:]��6�%zP�a��u�Ϧؤwk!ȳ&]�Y�&mQ�ۛ����%:ʪO4�Uxd��Z�U�˧e����٪@�ݱ�d{cY�i��`R̅��R<̿���w��RR��a*Z��p�%���Uʡ3\x2�K�RJ.�س�-����*���ݧ�@]L��GswMm,��Hxn�Z!�D����W�-mh����n�Dս�c��(�ʙ7i�۲6�\n�V�8%��Pj�ʦ��X� � ����O�1[��"Pʹ)LҬx�7���ؕ���z4�`����!�ŕ7j�X8՚+n��x%���`�������z;+5�=TΧBӫ{��Ѫ<��ǧL��:9&Es.=YgfV�!f-���V�[�q4���n���92��MZ����P)�yO$��5}*��q��j��A��V��f�h��z���@�*3x�L���3��^Z���{X��ov^���ybUe�^����]�[?c�)V�w�+mLEh���:)�r(��(Ct[�o	�te57iIN��YVp��u>�{F���7.�;T�+#8�噷�nf�CyWl%��	��I��P��M�Ʊ�oSH�jn%�VN���7,мԅ�ڐ��n]2*�6�V�9�j�i�d�m��4��Zp�%e#5Q��i\�*����*�Y�z���P8(Qӗb�Ի+N,2�f顒&��l�P���۷o�or�c�{C&:Leؕ��7lS6�͙.�+��/�DR�A�!��c[n�\(��Çn6�x-��˽�Vw-�{�-�{�*�r�`t�Kv��*�i{t�Pхa�Me�u�z�X�w�n&佩/1��i��Jߖ�7�Ge����5����5�{m�9VB����)��l$�vhKP��qk�5��Aa�����9��T9�L׋D�%И�QmeUTv(�.���h�Xˣ[92ԇ*��b��$��o+p��6+�.�����Ŏ޵���g$�v��v�˭��m^nZ�k$��nb̴r���4+0ؼԝ�K]�S�,֑���@��հe�ɒ=7�j]^�͎�h�V����9f��$�uU�J���Q��C^t&IJm^�+i��f]�F�JX��]*'-�j���RR���aG]Ե�)�ѯwF</JC`F6ȍdad��+����F�֥t�[���F����r�K�wzk́|�[������r�ȱ,5f�8лw�nV���#��V��ZZ*Zz�ט3wf�亱v����&�13�Q�T��
��;�D�b�@�W�,�˚�w[G^�pK�q%YL�;��FL���y)^�bs^+ok53�,�w�9{R���Me[��;�>�vs.�o/C�Xek�Ue�3":�У�V��`ںځ�O*����[��R��j�ok�ٌ���I���l��ݩn�8�6�d��,K[�&Lz$����̸��q��y�HW0
�w:ʭ�J���j(��f��L2�J��D�#KmQ�5�.]��"1�V�ݴv���d^Gy�-�-1a�*���1^�pm諐��ͷH�*��b�:Іiۥ��蓕PE[uSi܄B+a����J���^P�wJ,��Ӌ5A��L{�A�R*�6�0RgY���ù$�+h�$qX�D���(�`�cE�J�&�g4�+J���8䁬� �orE�+NEwSd��L�@�t&,����Uk*��3\N���www��֛�F�ܽ&�KU��΍c.m�W���HŹ���^����[�&<(��0�Y�j��/��D�9������*�ݺЭV����N\bbP=�˲/!ͱL&��v���!+"��=Kb�b����Q�������f�ay,�(e�v-e���]�5Йa+e`�-q X���kYNd�SB-�3a;+j��M����s]Ul�t�nಮa�a�Hָ�
��d�����ኯ1l��k)wW��,�#(��v6�"TK��8E�Ҋ�͒c��
�k�(]YV�����P:J�t�coR�Fd�ywcBT���L��c'>���S^ԁ�
D*{��K&G-�6��S]�̳gr�fٵ��#������/�Nm�nm�y���E�yp�@�ʺ��V�v+�n/��6��Ғ�PN�Kz��ga30L����b�w;4=�8�.軚��JÚM���j�����2&�wt%j��VH�T"�j�3/�Vֈnʕve˩*��nP׶�i�U4r�I6����P۬�qf-@�.�P��˷�]櫻ܪ�Q�ҭ�굷ma����gaW�V˕��뙤lK(�f�%�0��w��X�;̰��wI�Тٔ	��w�Tvi�S��kBaڪ/mf��}� v͙�${�Y�.��J��֤��_Ĝz���^a�o%���T�*�Ҹl�a��M��*E(��n@����ϕ��uاJ�f,�ح4�T.��U�J�,y��b�Z�_��Bk�ջqL{/	n��[�n�[[{���nQ�����I7b���2�k�	v0벍��-%����BL�Sf��˫:k*8776�Ȃ���F��8DP�k#4#߱du��;́^G��/v�N�)J���{4*.K���i���&����i�wx�H��eb+0��q�9ӥ�USr�5�F\�Ugk-���M�[N<����"X�j4.�ur��˭��J�w%#R�J���3"a-˛��}dz%n��`�ŐR�٣U{�[9�ծ�`v����w����n]��(md��б���V�5���9U���8uQ�5x��x�Ղl8�WzQ՛��Bm�� 3&��j����voj�f�)��V�Z���pi�k�.���jƖ�;�]`͸Uk�km���켼��İe�gkF޼ۡb���s6��N�A!�(C	�[
���w��p��yv]Ѣ���̼Z2Ա'#	n��F��&C��;[B����N�>���Y�Apɮ�͸ְf��x�D�b�����7�`��U#_e��Iaڶ������M�:RZf��	V��7zuf�zuԋ�Kzb�^-;��Y��p0ՆTs���x�Z��,�x)�V&X��T]F��
�S�n�c�q�wE۩.����-�c'Ix���/�b�h��aRQ=e��a_ق��C���ʹ�xM�*ɗ)�Ĕv������ڌX�X�#j��=F��u���r|j���7�f��&�!�t*���md)�ǵ�0ɔī�!HU��sH�on���P��ծ�6YI^e��d���`�{�����Wx�ݤV5y�7����uW5�f�
36��ֈڳH���%5L�J��kjT��s(�}�f�]��a���f��;��]-b�r��n�⺥�*�2�ei�I'CތKT��|�:�Gf]��J��8)�dL��ДX�ɨ�P%lӈ�Pˣo5!u�Y���Pm�k*�������n�a��
�;�*��(eʖ�DÕ"�9�kĆ�Cn�[Kr��7������ܣ�t�w��sN4�ee�\²յ,����I�vt��v�B�U�����e�rn��(�UWL雫XX*�յ��^
�75�/�ĽB�)M�&�����T���W����ڷ��u �A@$6�[j(�V5Z*���j���ح�U�mTm��j+k`յEm�j�F5�[�U��b���j�TZ���UQQm�b��Zƪ���lV�-TUZ�b�b��ڋcF�[EZ�ت�ֱ���j-����E���TV�6�F��mU���բ��6�U[%��-V5���mV5��j�TmX��V����jŵ�6�kQ�ڭ�UQ��TkU���ڍ�[h��j��,mF��j�6���F�h���V�V�ՍZ��m�ƪ�m���lUj5��Z�����j BI^?��������K��]��/M�,���ڠr���R����Z�	���d��͵Iݦ���W�8`�n�v��7R����+���]���헹�k
�&т��{u�'V貰5%ЪW�L���4TS�!\(��lR��֣j]�mY��#{[Pi}���SZ�g��5��]�:P�Ԓ
��1%�l���;�9,EdgJ�[3 %m�UL1F�xj���uc���:ҭ��X��h5Em���^���q�w���b��%u|u��z�m�Z�T�j�˶ܗ'J�A�Ŝ����Ҫ��'n�Y7N̷�p{o//i9f�����$nr��q�a���5�k�W��ݛ�
w5���Yj�okK6ff����]J�M��Y�t�^��?ov��U�bT�ǚw8sDU���p=#%�nU�/�<���P[�2�֕ۇ:ӭ#��*��m՜�B�+��dPf�Ud�]�\�\QWt�g3
���_}�]�o
��g�X]�B�Y\e֥�p�VU�x~�ܭ��B��vt���ۨ����H��uN�cj�1�)a}I:�fU�uy����d�T8,zM�[���U�U�(�^��wx�*��ce����w�����m;rѵ��i՚F�y]{�g:e��;�꺮IaU������۝"Bg+�����+�V�9]�X__P��<�ƭ[9�xs63���:�T��W�h�m=�ݸ0%�;4�͘�2�����Ũ�̜i��iK���hS�]U���ݔ�{�˔n�ɒ喸����;:�=[\��W�U|7+A9�r�6�ͽ5���=|Of�]Z�J?�IZ(2S���e��ל��:S�#��f�a?,a��8�l�ڬ�]�Ϋ�U�oT�7�������@��r�hq��Z��P�x��,�V%��b.a]aܹj�Jd+��k��T�+�ڛ���H�ӨN7a��vg=��-:Y雺S�����&�7cK2Cj���G��c�)_Z��nqح�7�TCb�*��0�	�L�خ�8��w��kw�^�O�}AWX�+���{�}�
mD��U�����x��N�D�C{g;д�w�3-ps2��T�'Q����K�<0,�x.�٠��\��4&��Y�֌����w^�U�����p�fuP$cm]m՝o��!���K���^T��zeJ�p�h��0��_4UvMl͊���٭԰:=�]��VtE��<̷�k��r��j�^�.��u�����+)jx�kd�ehU��;F��.�vj�%Q���b��ES��!��m���jW�8��]+珺��J�nfn�mX�A�Lژ	ײ���� FX��Gj����Q��rV�-t��H�i&�[�ݢ�T�y.L���Ǩ%շxu���u;n��	N�&��<ʽ��2E'jLv��&�����Uv�8�T
��|�#.�ܭg2��cu�TKA���wNU�Ig=��(�,�9vF9�S3v�tw�6�押 :g6��Q#�JOqA|v	��j�;�sn���[}�Ŋ�,-=ǻ�`�ۃ)λ��C}�K�L�T���ڗۖdݷ����A�q��5l�w��)uM8+�۾������D�Yۯ;)
�ֈ�T*e�bK��4�
�m��춴��p�pٷ}�x����RRGk�:*!Yً��zU(;˾�t��S�F�%&;;k%u�r�S�
4�����28�>�,pA[F��e�Wq�r��[:13�BR���۷g���|�bYj�P� ��mI}�7eb���8:]��<�R�餦�M.7�yf��˴�k�����0,�/���tC�c�v�7`��G7d��VX.�+s:���^�hA�����r�W��cjn�d�5���u�a�r���ã)îٻ����R��U|˽��:oU�V�A�ww{���ס�����wY[�HP��u,qڝ�'������ڪX�7�ݫ��G*K�S/%�U:9j%K3������ȉ�V,�q"���CJʮ�o��tv�v�J��/^���L1ףr����g�>�(t�X�jb�����P�T����u�}���Ae]G��:wT��֢f��{r���ս�.�{�n���Np��S�¸�{Uw���ް��QhtΡ�2�\�>�����9Ω]NU�Q�a����������y!u��)�K.��V��ф�ޕJ ���%�S�Lmk�?��G`��.�Ws[��Q������o�P����6�S6Ӡ{��]%+��ٵ3��t��4 ���*^���]-�M#��i�'S�}g2��y�+N��T��e��7x�wq����.M���u޽���cYWg�2�pP�b�d�,��ܐ�F����4�ne�V��Ԭ��n��wʾ�V���ڭ��8�ԭ(nSWl��G+�]�S)�춖���Wy��;i^!�A���M���y�4u�D��Kb�uLd�Y@�M:���!n+6�qPLz����vQ�1�H��W�vb�]ǖ��`(U��UA�y�us'$��u_�?��rt�\���OG*v���'��ޝz��쑛d-啝���&�%ivjx�T�D�y%�1#��|�w+zD��Gyn�9�bݙ��n��Z�/7��ZA��zx�m��3O*�����ʲ�t�(�ffX�R����ىi<�Q�s�w�E\.ƪ�[]-#f��`Co+���^VWp������J�2�uw;��hb�7\�gUff���v�6{b�Ëm������B
j�Ue���-��wγ���Y5Y�����^�3-���awO�{�%�w���E�W��4��{��c��,�
���r�V�B�s�e\OuZ��-�����2û2vN�����\��H\�u�]Ժ���<��´����k�޷U�s�u�2dEXb]�E�Wm���ŀ֕i�R�=9��hN;07W�������y��в,�3e�ٛ6��|v�'IlfƟtw� v�a�Nڧt-쵍�5��2��y�bS3���)�'4�wf,X�՚o�ʸ���WnJ��m�Qf�[�J�9��W]#����#����:��ޝ/t�uZ~�o����(+��ε�T�;ںT�ַ�SQ5Յf����s-M��f��4N�l����5��gg�Q�U9���YF�7�e�|�ni��A}zƸq��i�3d8iV��}��]j�,q7y`�ܕQ5��E���g�j�;a��^�%�3t��+]آ���ͪe�Gn���B�,��v��d�.�����N��Y�˒�ᆁӛ[�F�A����6�Ƿ�+/kmXv0;uB+>XB��xQ�Z��N�>á����z2��-����;w�-�}�o����e�m]=��A���b�3�t{[9`)lݾN����;�j��!�e_�S/o3D���WL�Ŗ���uC�ېY솜%�!�Tz���V6����*�� ��Q�,E�L�҂y�_$D�b��2��a*���V�t�t\��Օ��b�hV�um�U�7�f*�6�b2�Vuc/����|ba���uJ�c�j�,�]�W���ڦ�j�ܫO�4�%x�B��u.��|��p�׽2"�6ۻ=���|��7�����E\ⲭ�I`��2͎����|*��	W(�X�����:�=��ERU���EX�5D�n#��닰���@��Ӛ�r��9Km); �t+6��Q`�����\����7�Uf���{��u�0�y&o����CvFO����\O;'۪R�A�w�*웰N�}���r���V�u�B�р�����fLgjQ��,��i�8ڛ���\�+�(�f��Gkp�,,յe��9�MS79ފY�w��NL<u�2�UT낻(���w�!a>�#�c
M}!
��x�X��n�q��r�"�E7Q�M��n�,V$���t,>�ņ�,��q>˽�
�F���6J�h�
��+n�=�������x�R�N������o^O.�)�5U�1P%��[�b[�ѶG9�[��fά�K��3%�-\w�wpt�ed��k独��q{�s��]�@��+{)�S5fh�.!�5�d���$�E�f�;H��a���9U�A��d��њMnnԠ�=T�x�[x���vLQK��M>�i��.,4/dG��X���k"�ݬ��o:�����R��GU��6-�&��[U�ٖyo�h�r�w�9wX����3>�W`��&�t���fU>�Z����λ���j�6�u��S#v�__!}�Npm���1��چ��}g�}�7MuM��s:��k�U�Mi�����a�J�r��ٷ��o
���'oupU����U�YtA�ޡ�<��{챕U��Z��]NkK&�)���C��7�o7)���CkE7�Q��T�뺫�﷯>��y�z��M�֤Ԡ�U�&؂�u;C]��W�j5w�36gYލX���]	u��V���g-�xCΥ�,�UR���9N�ة�jP�!3}�3^���~o���o��T.�ܥB*Ӷ6�d�S7�M��L'��EmQ�K89`���mP#p��5�/���<�*�=��YJ$�4~<־�\��S�˫Y�,:�kl.�7C\���}��;1e��uڴ����$NU��g{bܴ ��d��a�j�\�S����
���3�+w��+�ӱU�h\62��A��[B������Ց\R�졁����\v�s�!(����
�W�V#y�=��/:���o�f���u�S��-���a�6�qr����o��Tv�ە�(����v�"ѓ�V�V��v�Vn���PZ8�Q�V���5����h�O�N[����M�Hww-�FR��_QgQ�+������Vv	׆uTrףeP�o�����e�f���WR=�&���1���ڹB�1�WaJP�˱��R��b��n�#j��J�s;69{Tz��(�.]Ǚ�4�˻����gn����]z�6�`@�ч�]�R�9��@��j�>F�+��hW��Cl�Z*�:�e���KN��N���8�Z����qTĪ��X�u�5n�����7P˨L[�`�Z���5.�Z
�]]Au�s��+M�Qe�z OM�b�R��s��q��"y���me��=o��-���
��j�'�O��R��#J-=38�Fະ�w(^��꯷�?IȊ�y�
���<� ��;L�i����R�'e��ͻ�4�7��+�鵵ܚ��K�m��}����-��sX�h{[��z��S���'�pr�b#���}�Vk�ـ�����A�b�	2];w+������b<�J���R��ֆM_Uf:��b�h�//ph�ٚjqqm���J�7���U�y�/,g]��\k�*}k�y�������T�Æk�@������-ߊim.4�%���es��7�B7�v����+9���9M���\Gst�^іE��8^�p�D9J�aE��r�r���բ�%�z��w��=X��7�i��4�>�:�؜��S����흾NKPU�I��;Zk�f\��}�oq'��E�]��K]fU�p��0f]ޫ<L�G9�[�S�ݎ����[pZ�]�:����#{�R��{5�)��h��1	̡��93J�B�]Rw�ӽ|��G�Y-�hY�v��1m�_J�'5�������֫����.��D����:;,��5}!mLy����yJ���9-��3fͬ�r]&l��gjjBZi�[�u�38�ٵ�F��n�5Y8�C�r*���nh�)�f�(�g�a÷���އ��n.�o]� ��w��C.�d]�[�ܾ�x�u�u]�t8�^'�����l�]4�ҭ�Ų��کu����WV�kw.��iޛx�"H�}�C�]�X핎AXLT]�(0Y�]�KŎ��E���W��� ֶ0e��nv�:š��2�������k��ea�oQU���J�+k4C��t��ׯ���|�_x�a=�4[��~�V�����f�ɶȜ`Bu����T-S��bɗ�[���Us�݀�U����s���]Q\��mn�	[�Y�r�%3m,8�sjls�l����yf>���SW{�MN����#k�xT�r�����v-�8�,��[v�A!J��Q\u��T��WWJ���ݓ���^n�3���*y�uUf�*mr}�%p��Wr�
K2�qc2�\�3$��^����gx�ٛ[ϖZ�ǣ&LY	8+ ��Y�֨z2����у{�:���݌:z{t�[P�D��]	o9Uy\�mfuj�����ڃ�XpUV�;��;P�r��YO.�#��j��c��N�O*���c%q��Pk�
%�|Z�'Eed��wm�2�6���n7 �S�J��E��y��.g̼[�T�.ƕ�K�N.Wc�&u�fl����ƅ��B� 4�
�;y}��AX��c3]oO�U��q��c�o�ڡ%n;�/<J�ņ{)����@i4��ؼ6*��9�y�`d�ݘtܜF�G��t���w�UWz���*�ܲ�.)��b�V+��Gm85�⼭���Z5(9RCl\_!�ZY��1�!�x5h�O�*6���z%]v=�NK��.!Rk���۰�t6�;����PwM���3{+���ӷ�2�8�I��O��N��,qu��c�j�M�Y4n���s+$o��R��\��Kz��)Vj�<�wGY��EΌ�h��͹i�%��G�,�YY�}쳙Xe�9�����(Sz��&�x1��AN��W��k�y�ݻ6�c[\��+`I^�����*�7�"���n�ޛ���v�o��^����^�{��ص�ϩ=�j��Luõ{8ptQΡA_^�//�$�k[}]�T]��7��;A��7�nٚW_gEV��n���m��ۥC�J�P�c/z�v�����N��i� �.ٶ��>�O=E�Yb��1�N� ǩ���dI�pA�� ��M�z2�d����͘qVк�;zk�7K��h�_J���xx�GuWA��{C�Q��uU��&���-e�3qL?�u�
��a��P��n:��cjd��j��b�f�,)�ٿ�� �	&@ ����w�u,�1�̢��j�N>6�^�+�5!��p�fY�ɍ��<����e��q��xv�v�I�\4�s �1�3 �d� ���M��jp,��5���3j<KV����e)�*�51��k.���1��V�-��۳W:����)-n�]�M��f�33��ƐS��&6t늮8V�T�R�a0�[4@����s^!��{`cm��l�i�h�^q�Qo[���1`�h_/<���3����)��9,�`o S���q�]1n�K
kbtb{<^N�n9�$�+p�7	-��l�ͼl��+5��ef�5l	��Er�۱]V�C<<�8l��2 V-�&Q#�����]�m��*P�C�+�k��wl�Un�2&�t���3e�]LAٮR�%v�HA��e-������Ѷr8�����Z���y���<u��S܅�� ۜ3�d�����WM�k���5�KW�ax9�S��[=��ix<%<u�v��8�Z��Er�Gu��z�a���z8\GE�k��k`�{ء�;�զ=����Z��ƍ���%����uL7WNB4�콸��h:�L�[��NLp�ʀAM�U��D֢�4p��͍�v*�f�4CXb!N�"��U+��u�u�����7:Š��7`:�%��֍7�Ζ������0]o1X�j�̚W�4of�c�CJP64�����3	B	�66�mB�=Q�#�c���n��Nn��oa�`uqC��j6X��7��㫮K�ż=��v�8�k	�L�&���Yu���6Э�R܉�*��IQ�ӝ����[(�FS"ͷk��LV�g���"7R8�]���k�^�t��v�vm�� ����{t1�85�om��v�	�L#�[�� ^5bv�f���7C���$U��Zj��FhJ��8�mB^��,�L޵0�j�YBM�b�=���q�/�[��%VX��`!��i����ʄ�K�-6�i��x7`.t:;i댭ل�6�q��If썸%�I�SI�l�\-��;��C�U˹�"5۵j���.�e�*�z�G]�����Q���GE�]�غ��Ȼv�QѶ��>�//OLrv��fݓi�"�,��x�2�/�6���7�-!�ς�6��ù7G��y��v^��u�� �%�Ka�2��X��*޵fΑx��3��T�C����.[qώCc����9����ӭ4س��%�x��il��[	cjRh��Ys0,JU������뫴ڨV�t�]O%a�r���u��n�ԜܴrNڱ�;���n��L�r3s�����3�`�]�.,��`�TZ��f���r��N��U�kNyNۊ�� �}&�ۧ�CĨ�l�m2l
k�уh{q��uկuUarD����^��+S�mϲu�o �=1]����͸��偧%�p����k<��2l����1\�U휤灺w\��f���8!M��m�e]X�6��)�{����C�sWa5n;s2��'LX�,lN{�8P��;.�n�h�f!���-�n<��l�Ѵ�r��<�j�����[vC�X.�bak���n�l�F�9�>f��ҝDn���58��ϳx�԰�{��x��z��t�Q�q؇'�C�D�st\u]f��{h$�{���q]=��s��NW�1ibզs�"���7[��� �u��A���jR�tX�[-/$�f��'rK�h�Z��WV�^+vW< ��h��[����T�l�9̱��tr#�ꗎKZ7�.-�ɌX�[��nuZ����T1l�t)�*��l���i��ٲ�a�okM�� ���6Ls��#�����,�6a�VR�MF4Kt�:n�ݺ���y�nע9���In�o:�Y����<��6�[.��l��J�6�t�2���V�K���m��/Z�j��[t�(���" Ƙ��0�mvqݣ��tw5MMIQ�F]�[���ݩ�f��yb��Y��mK�;X�t��:�UP��wKȉX6]��ͦv�ٹc���-7m;j�/i�Ϩ�x"|\��ui�W9S�C���/6;]Tmv�X��s�g�Pp�ܭΆ��v:6�G��;(��њ4���\B#E���v�̩1+� �Y�T����«A��7�7�Ef炃lrgq����n=EB�z#h՝�V��\k��@���V�(�9��q���h��Mۛ(,t�<�]������i�HKE{Vj��n�;��u���魃��̶],����18]5���ַJ�sp�ݹ^trllZy�^n9�ݴ<��s4k���<��1���Z���\�,��]�D�aA�3��[�!�/�z؆b���vʯN�͚����5�N��=tr�S�*_'�K]�[�[���W������,b�'��݈��;v&�̵ʼ�՞�ȷ3�.KRͦM�В��%bK)�&��u`����]�B��"��`h��)_)5ͧ���;���>֮:]\�z�W��(��p�_		w˜̻�{]s��8C������f��IAvtt�̼��]���N{��.�O9�=g����]&��s��Z!C$.�J]����hʰ2�zF��{'q��+�f�-�	�v�3�9�\�� bj�Y��ԅ�c�[�v�iw��JD���,����Z���ǧv���Q���'/&2	f-^�;g�����u�tn�F<�n���l٥�(�P��˙��Qff��I{F2�%�%�2�Οst� �+���P{
�3s��mIv�������GpvsWC�}�N�v����@��׷$Cd�m�n����u�<*HL"vU���
���Y��!�	�b�m���a�3�k�^2X�*��կm���0g7��ڏ�X#�(K1u��{��t�\�{<[5�`�@�/cGf'D7����LPk��z��/6�[��æ5<�<`KcP����i����c�S�!��J��X�L��7g@���@�V�v�Ŗ�km��B�8��p�H�&B�5Є�Hep<k���[]\��&�A΁��;��s',rOB�XZ��v��ٶ2�E���۠9�kIup�T�X:\���! ���hl���7+��&EIt,`��X�UF;Jlq�9��/8n�ŧ�0ZnkXz���9�d�,���t��r`�gn�n��I��z[^:9�oY�z�S]qM��m]�H��̴�h�`m����u�f6ր���gm�'B����]����0�m�y*_Q3��7`z{<��ۍ%뫌��u�Ò�q��n#4-�ѡ�[V饢�'<��ѝ����B���*���!2��u�����ۣyド�6سԬ�/#��uvt4&�����CF(�ex�USp�m:h1"U�KE��ї�unx�z�'��`�M�5ؙ!Z����1��i���!�<Ywk�Wc�I[�Rb3LKz�Q����uݛT<��ۋnM�2�vh�g�-xz�ۏtct@�(K�h���p�����ol�h�:�U�ĥ�M�P	��h����5��I)y&�F��I�`0�M2l�\]4�vƉf��q��v�OPu/70�t�s��(�MHTe%ba�X�m�������Dc��\�E���c�X�[��[�*�t�6�5���a��K�,� ��$�����[��b�k3)��eYn���e���}�e�m�5,ٌ��Vh2�ͩE-I!�2��e��=��j�H��3�o t;'o^�Ǎ�\�IɽZʺ$��u��5Ö�(%�%6�Y��:�ೀ���zP�f���r��z�t������v�J7c�{�ǣ��:zx7�%�]�\�t\+g�b�qg��[��R@�v�mubx�����t�-�Y�!q�JF�Y����ŘW� �6�n���f��=/t�j�|[����4�n�Zh�4�;��Gb�bd@5��1����bYk*P������ZH��l�k+�s��pWY�u]0& ��ӻa�7"{b��놏nf��U����1���!�m�,��qa��j�Gs�`��n��*۝x�T�4=lFI�@a�����d��n�4��毗����U1v���	��i%p��ؘ�7`�)�#R]k����O��kfa&^� �v���
M��eζ덈�m5�5&�k�r�7�|<�xy@2��33&��\bͬ��y�ǖ9:N#��v�0ǟ
�IF\&��Ja�� ͖�=��5%�E�6�
l8 ݽ��cB�q6Ƅg�K��I����F(8ġ.:������ti	X\�M�u�Z6��&�8�ae�&Xݭp@�:�;=�&СY{TW�)z �\���v�+�=l�k��M�q�ݣ7j�Zd������!�+�lJ3�q�}�]v�q��uwZ�rA��<��Y� z5ӇkGkW,�릉(L�,"e+.,�F q-��J;1�km�ݦ�0d[]���}g����Gls0��6�j��fm��|���xф���?�|�s�b\ ���/q>޷����ܤ�����맳��E�x�W��l�%�6��f�`6ף��|ˎ)��Ġ�v{����]�G�1ض�F^x�R>m^�\\��Rͷ��6c�ƌ��-�����eH���u�\�3��[���t\p/����܆lc�x�<#��t�w��T,��x��(�r6�or�KlG�`�ή.8�lz�1n��f�,4#��(/,ff�'�ON�\�<�Хm�u�2�a�۠�3ك��
$�4!��ǠN���-�=��u���py�c���K8�͝�pj�Q������:��0Q�<ݰ�ץ��v�j�)!��b�G(&z�g��E����A�Ƒs��Yx�t����S�����i�m����ŕ\�of�5�X!I��-Ԅl4f#݇)��5�l�fY��9v�6zN��Y�l�l�LQ��QQlb�5F��%���[cm�Ѩ5���b�Tlm�hڍ�V6�Q�mcZō����BTlh�#[E��*ƲB�DTm�U%h���kIQ��Zţj*�PTb�2����I�5�b��VŌRjؠ�T�ѵ"$� ^_�R��żm-sv��<��t�#�p(���LK�eB���Ô��sC��`��7���D���7����Pu����lh��a6/;��u�n���O#�UO7���1�n��znۀ�5�Y�b�L���+5�2u��i����`A1U��W �*Wa�qCL�*fp��H/n:a���\G.b�\�s�<�P�Y����W�ۧ{��c7q�-q�����mǚ��4T��ba`]��e4�-�l�V�O]�9��Ә㑕�a��k���u�n9��汷nw3��<N��q�E��1��nm�ɞ��6.���n5Y
�\�=�۩�^hN���L8��e����۶�&��G��
�D%��)�l6GV[��݄�1�ڈZ-�q���\��t&#�Wc3��sr�!3���
D�q�.5��b]k�g�s=�^z�]�r`��K*F�!�S0��iQ�\6��s��4�aLy��RuZ�v�f-��ӎ{
"�t����+��CEIR��da5K,ŰR��K,X�f�7�C]م�F�*��]��g�l��U6&��,��&ʅL�X�����C��.����:}]��(�;�u�8��x^9�͵�C���^ǆ1N�O �a�{9��V�-vx���4�3�3H�&�
���.�kq�u!�;��ZD+N0u�ls��1����-��֞�+g���^!�\cY'`x\�W'!3����kd�h;�j�DA3�������G��n[k� i�	��=.B�r�G�Ʉ�RT�Z)���Rb%ti�.%N�s���A�l��V�-�)q-��u��g�a�Tkϫ[��>;���P�Mr%�N7Z�[u�8qn��=��6ch��ͮeR��Z&G@у������j�����a��r��*�+;l��R���U]���-��I���Gj0� �܇i۴�s���_=t�:C�{����
[+T�H��mj�jrr�jж,�xBӭ�Rl�c�X)�-�,IQ�BذlK+Kz�$����ጶP�6�RC�5%�ՊUX��
wT-ᖅ�@��������@�VXP�H��PZq�C�v���;<��T
0#E��C��2�,`R�������_���D��.��.�v�)�,�]��1�rn
5�
��k���������:hF�
�R�l�
�L�0�P&┕��"��b��͠�-� ��(��c��Ku/�%�+�o�*.�z�VnN�#�'��x�t�1G�YH���r�*�!�/���2F�kH�̭�y��q�;�y&����|P ��@�_"�(�@��z���9@hu�"��A��`G�'��y9٨a~3Ծ#Q�����/�#�!_oW��~,��-��tP����=�~_i�����+���}X��dc�@�zP_v���`!��h���=tj�_Ť6�ؗBgj;]ǜ8A��s�Olɠ�	�7J&�DՖ	�P'}H���U�t�ͬ��/o�v�ݝ+r�Em ��^�n�;)|A�Q�źP�{����ET�}�`�?dP'��$R�;�]�9/���*�uIW4�"�|t��)��\AÍ��СAh�a4�k�Xi?vׁPB�}�����j�٨a~�3Ԉ/�@�\}rnC؎^-�n���@�Ŕ���K��t#�{}�/�z���z�bsx�5����_"�|����3v��v{�U��s��u�t���K�9�T^�L�ٻ:V�}㞠�!ShC�|[����A�t�����Cu� �[���S�Ӊ"4�>��a��o_21׾ �=_/� ��?Bn`�a��v^��*�*�iU��mV,�c7�ē�ܥ�l��fk���6���ɛ�l�u���H����u�M�띉����C�z��t=�f/�3�|AmCt� ���k��:��B:�?��O`�^�L�׻��x�z���h [�{�l��G7����vPD2�@�H���!����ԗ��t�s�۵{�������k�*����UWW�y�NX��0ɽ�D����YR�v�GMˉ��y	ͼ�}��mp�\�����x�ބadx��H�2Я�h [�Gm�(�R�(���� ��m3�8{��n򝇐/ h-���Z��=��}�� #҂��T-�ɴ-߈�N�'�]h�u__${�]R/k�gk��r�����m�n�_Y�׎ ��y���$�J��U���������"4��v�4��V[�.Zj6�_Q����A���n�n��T�a�3�;���#��j���෈�~� ��@q���:�E�_K,��k�����AΠ8���u����y�Sx0�͐An�e��u�V^r]n���c�h G!t�?�D2�|[A��ٚ-հע������2�A�k��u����!��F�ozm�P��x��H��h!<�}S{��Չ�l�9��?k>�Y��ë�U|uR5eW*�gj�D���!�Ei�������@�e4�1X��%�X�w�;�t6:�5KGsHٱ��
j�ɜ��Ðx�>U�m[���2̏�#[���4�8t�׶�����7}�2�u;\~n��Ю�J��L��H:`U[B�U#Y��D���r������J`uʭt���U�αp/��i����o�>��U�tK4y~�ڝ�y���2�/�#�=��`�"��",���%����޺;�`ê����H�w;Y�݇;=X�{�E�G���� C,:�ê�u��� ~�� ����/� Y��_���h軝��=Y�ns���uF�!�"��!�������ǵy��?=A��|��G'��<�>ә_x>(����v-C�_"Ϗ����/�.������ho��t8�k|�0�=Xӭ�#�A�R�A�B�-���C9�_�޽U�Ϟ�U譿*��'ՔĽ��t�E���V�n���v�bX9�~��XL��\L�G�����u�iK��ޔUҳuEh��r�ba�Ku��c�iZ�`�CmC�Xc�%ÍL��X����R%҄+`�w��ƈ�b�jͭHOn�r:�u��K�8�GX��d�t:ݔ�����e�:#��p���^�uMt�	vv�qÎl\��DM�0�����6W����g^8�.�Th]�@�"^Ü�0t[�>ݞj�[�C
����f~�^��o}��S���u�Yӭ�붃;iF-Q�P6��)�B�GM�U������(�$A�Y�'���{�<����hM������>*��� [�� ���Z	n���y�[�b�Ha���	Uy�o��w2y�}�2�A�>+�͠�n�=�lcݬv��?s��<�/�!�!�[C<}�^AY���y��k{=N�oqw>�D@�Z���-�"c}�Oz�i�>�҃��ؐA���#t=o���,�9�C��u޴�Âr�
��7�__y�*�H��(`/k:b����/���yk��L��a̯N�-��0�熣U��\�PH�
�<��
=������;m��̝s���#���f�������_��@���2EdIA���8�[�}5�F"�Y�G�,�Z`�3dQ�%!��(� ����L�nNf՜�\���Ht%��f��o����s�����ǣ�E�༮�^�-YQqsG:"�ॡ#-goX�&ӵ����.fbliۏ���3����Zvi,�XyA�C���A��\���.c�G��ӯ�C���7l��Yswp}2�^J�u^�)���ۆfM��<#�9����?k�,)~�o�(@���R�ɽ@o�L�c�� �]�������q��0ﾠ@=�/��q�a]�u_ϬX2W�(����R���]k�0T�	��w!�+q�h�B��Kp�Sd��f>���l����wڮ�m��.늢�Jn\�M��i�KE�5��X�]��a�ݿ�(<�o���i�V?�5yv=��m(�e5Q~������R~xw�;Gf��`�q;���;���}�����yX ��{�ީ��M�^�����Awf�`I	E�-n%�X������b�u�.PD%�J_������	��}��[%�r���՗���<�oL.ɳ��v��}e��]cN�Q�G�.�v�������^�z�وJ����^�pި:�rr�{�m27��{� A/�2Ed"J����=��m�דV�A� �r���%����������[��A;����[e�Y��*�>؟�%�	 ��������!��H��yi�!�C6u�������G��+Ѥ^����Q��)bzt�Ͳ����b��غ���RJ��A�6s��v;�ĝ�l��9��j���u�{���Y~|�A�t(���~zN�Ӑ�j�<�K#q�_�y��ٽ|d+ʇ�?N_ \�$�$����}�	ɗD��;��j������m��7Q������	 ���QJ*��~�w�{�	��H"��,�A|D��2ED�P�𓓽x�׎�1T%�z["����~[ %��J�J,�ýګفI\A��hW�6$�P$1�[i�1�y��2>�͠An��Ҷ�_��C�d�5WY��W/R�uא����b2�ލk�嗸�*�_tݼ�����sv�D��ڼs;j�eƭ�S�o׮��8������|�CH����A�D�7U*��}��y��~���tu�8�Fex����?7,XJ@�d���ð�f7�{�J�Z4���Y?+ �*���!�C,��ͻ(���\�*i���Ͽ����2����2Ed���j��A�v�.�^W� 齯c��{���~ �A|�R���ř)���Q���}�d��,��2PLhm���m]��,?O�Ep$���&H�onnoz��uz`M���H�ܬ�"�($��h,�tO��n����=ӗN��?�A�,Y���d��K�Kށ7����"�A�=����7�3_��h��h �w\�"\Q8-�z�}@hs�Y�� �%� �%
(�Ƕkl�Bd	�a�i�Co9�y V�,�J��|��+ �"�y7�ǹ�}�c�֫��w]VvX�K$������
�>[}.&2�i�[I$�`�SU
�xxF�GN���y�ι���j��^���AR4�:�T,W�m-��N���m��lrd��cf%�B!ie0���׭��xb:z����	M��>�x��[c��.��b�j=Gݫ�9(3$��3�Y.n�F�H�TF6R6��P�Ba3*U�`�`�랷nT�7�3D>7f���Q��N:
�1k�W
��c�.�p=:;k�N�DaX5�f��Y�ǉi6u���_��'���1a��w����K������s�X�Q�f(��0���۾���A�)�A�v@J=����Pӗ�:}y�>��>��B_*�M�fZT�A�\�&J�%�`�%'gbbK�pu��h~{"^jY�7�_��Jz=����A�%<�g�!k�瘇��_O����,+��ٮ����.}�=��e����C��@I�dA% G^���������8��I,z�ǣ��;�r��[�A�PDs�&���H�\�A=��l\��/��#y�;����{�<��:�:P+�����Dn���?�X�/7GEܥ��b��l�A�4�� .�Q��^�Xh�Dtsv#k�l%��ILfT0A�נIjt(�IJ��m�>n�po�/%�8T�w��^I@/j�ߗ�$A% ~�+#���<���)��ުiu�ő�j�E^x.V��t�V��JQ��vݕ2��F.�Q��
ud#3���T^Q�N��KN�UQ�c+�������x�F��}n��y���9H�[����_k�,*�ni���N���-?o3r�7n[����H�:4ȭNU�i�:ϛ4�{Ѡ@;�4/d�|��E(�B�	�[�풳�0~k+�Q`@)@�x��^�ٸ�	o���P���ǱFk������@�)L�YD�<�W���-_�X��� ����;�r�^w�q}%B	���}Ｋ � iP�׬�����,�7R�k���ѱO1V3�Ub�Zw�� ����"��7��'���g�Wqȅ��x�k�Gq0APDq�_��,)A��e��\7ll� �ȟ� �fX���i��H[��������;�@�-P'���D�/��*�H��l�:o�8r�Q�Tqw[y��U�]j}��!V��D@�:��J-u����n�gPy��-���*��.�&͈83l��{v�&C����ēa#�����ee>�l�&��ڜ�j��fk�0�������duB�С��T�F� 6��������A��V�VK�e�c����i�1�.�^Hn�m����A!��`�ܴ�6����b��E���[A��ZM	բ�k�tW�]pϗc��92�HĪ��N�5%̝�o9��Ŭ��𰺲���:Vm^���Yu�l]RrRuyY�yW����v����r��EpD�vu��U[�1��$u��{tk]mSrt�}u���R3����$����k7{%!�);9���^����;\���{ygR��PҲ#͚z'_e2�>�F�K�]�;�5���r*슯��mU���W�Vy�17�LY#B��nK��Jͬ�w�C����Tp=9�V=�s�X��``�Z3��Cz����В�n�S��t�s�z��mAb�ү�Q��j�]lkO�7��-}�:�n��vv)w7��)�$͏���!z���Y�ԥ!+�ڕ{�s�l��Ek9(�v^[r<Z����:rT�5���MܧUV2ha3wT��9��ۧ�[���ꕝ��e"t��"��9EǓ�w�+^1�Wζރ]�%,\�v�L.�+����W�N�aȱg>��HQ�=T;?o<�zӤ*�W[W��������!�F�K�J���!g"jӯ(��F���E_R�7�7�Ù�;7����^[W��0X�m�Z66�j�Ѩ�*-$klQ�h�5��Qm��Z-��X��h���X�جATUQ��Q�Ũ�j-��ƬIDk���lcm�1���k�lTZ�T�#h�Z",�0��EI ������癚~�sy|�1��i�$��_\
H)�n�!�Aa�
@�(���$Je<�\
@Ĥ�Ü凟�>�����f���/�{@P$���!I���RAL@�s�g�$�$�Q~��9W�ݲ�6��C��\
H)>)��}p�ORA@�/�?����;ϯ�䂐R������v�ۇ��`R9E�D
H,��O9wCRAaG9̇���)���>y�s��}�h~H)���(i�x����>�~9�
AaY���Ă����E��B�[|��S)�9ˆ3���
9E�^������9�;�ߔ-��%؃�=�!���m�$�-vFݞ6Y����wj˕y���=�RU������B�s~�c'�) �Q�Y���$�ˁ�tAH4s��o�~��ff|~��=�_;9���Y^w��N}��}<ｓ����RRAaS�܇� �}�-'�
H,�2�W. a�s�>$���Qi
!IN�ʯZ���^��
l@�ݸc<d���D;�0��?
˓�q��+��8�w�qr��RRÿ}pĂ�P<��bAH)�r�~�����f�{�
A���{p� �F }���I��Ok��Ĕ�XQ�s!�Aa�9�-&�R�����W���m�dp��S�vz��H�����|H)
*���i �6��) �0�9p�x�I
C���^r�1�$�{{�x|yW��׺��<�bAH(����X�A~���D�EC���Ă��w��Mp�g1���<@ I� A�_~�������w���Y^~�/��~7\v�e�_s�Ґ�!�*9y�Փ-ͻ�WIk����u��̸��cm^,K]Ss�ǩ#�rŦ�Ǽ*��x�aĂ�����ZLB�%�~���I�9�
B�T9E���\9ˁ�2 Ss�c$</��$�{R�����~7��p�j��ߺ�a`s���0�s�\Bn��A�7v�3���V�����e��L�GM�-��t�{k��x���슜�C�Hhg8ՖU�4��>�E��φJw�h`��
=�r$
@�(���$JO9P-:o~:s�����<���߅ ���a�|H)�?s7/N��������RAk��$��yۆ3��I
�(Ă��^r�#H)*!L9�\1��RA@�~��������1 �0i ����
A��Ͼ�x�^�y��]_����������i ���O�TC%${��x�Xx9�-'��w�9����&2��P- ���z��R*���- ����s�
b0�9p�x��P��9F$q>�wԽ��4�s����o����W��>���IG���{p�O�RA@��Y� �����)��9ˇ��`R9E��Y�{�v������C�) ����!�Aa�7�ZL����~��|�}��i)�GW�<�k��XV~��� ���p��_h�|-���}�W q �P)�}ۆ3�JH(P�9F$RAy��1 ��)�9ˆ2x�H(�Y���I�*�<~�o�<��G������b���T���q��]�{E��$S%>�P-�) ��ypĂ�P9�-'�
H/�A�q�@u�I�S=���+�V,�͠����ˊ�@�KN��U��v��9N���ao�vP{���Z#B�q�=�j�Zv��]�kr��z�|����j�����9�:���BgU+��t���nb�ld��غ�m6���L����x��5��1F�0!*ST� R�+�\�T�iC���v|M�+��a���	�z���:N��˵˃&�'<c��c��=�pz���y^��nI�9�FD�a8�v��G:m v��u�:N���ǭώq׷<\�,�]����-۾��Ͻ���l�Ź�B�ԘrQ[u1�c���K��Pp�ō�%6a��� ��a�Ă�P9��r�RAk�̀�ȁL9�\1�FJH(TC��?w}������7�os�~�$���RAI�~Oٞ���2{I�嘐X�A~��D�EC���Ă�0)���
Af��p0II���x��~ұ���H,4aH��I�RAH/;w@ϵ��os�?y�\��y�
AaY���� �*���R
Asy�H)�0�9p�mw��<��y��~H({E�aI�.��RRÿvጞA��P*嘐X4�^r�J�G��|s��}�X���nE��R�_�/�*�Q����<@ IG��������$���d<H,<�)���`!I��S�]�P2	I�7�� ��Y��ݯ���+�ZA�!I��s )2 S{ۆ3��I�����������S�s<��� ��]��
H))
aϾ�bAH(��n����gy���
AH/ݻ��TAH5P߹p� �
@�(��
H,�Jy˸
$����CĂ����Qi�������� ��n�(�yϏ{�>��m��}��R�e���AHUP�- ����o3 )1�s��c<d���!�Q���o>����z[����?)0k���!����b7s��6J��j@�e�ٗc�e=�${vF�RR�{��<I���H,i ���� ��s��x�_{����k�_��_��8����H)�Q������?�'�wC�%$��!�Aa�0���I�RAd���p�I�9�
A@�(����>��J����������I�9#>A��Us�h`��[�¦~�,�-c�J�i�۽o��׻չ&U���ū��+�U��_���)?���r��d���ߨ����}��8]��Dp^�g|<G����8� ��"���<e$�E�4�^r�~�hO3�V�AH,>�.�_F }��
H,��N�wC%$s��x�Xx0�r�I�
H,�O9w@���]o;�Vcs����[���?
��8���"Tv�H9D) ��̀���s��c<) �Hs�bAa�
H/9wH):s}�wz��CXg��bAH(��Xƒ����C�H���n~#�O�yM���K~�O��<@�Z}
H,���~�����|�ֹϷ���yc����x�Xq� s�ZLB�%2���"RAa�r��� �*�r�H9D) ��� � Ss�c���~������������~����~7�=��<H/��a�aI ������H(��H,��]�¨��h�s��x�_�����{×~���7o���[��u��\]]T n�,&2�:��m���ʲ�k9���N�
H,���߮�) ���r$���Qi �z�y˸
k������Wռ�����H,2�X}
C�w�i8/_M͢��B�^nd �0�;p�x��P�r�H,2) ���`0����)�9ˆ2yI3�_ok�g�H,�����UR����Ă|3�M�P�c�~�M���G ���d�߮�(`��yˆ$���Qi.�����:����CĂ���{w@Ĥ���{pĂ���E���\�3 )1�s��c<JH(R��X|w߾�}�߻����y�� ���s��i�Tke���yW5��P��ӝ��m_N^2�PJ�q]k��=��U6��&��wWd ���e��� >^��,�;�dt�<���$��
AI��S��ጞ���A߬Ă�ƒ�]��TAH4T9�\<H/���r�L@��ϸs�m�j���O���p?JH,(���<H,<��Qi1
H,�O9w@�����������=�
Aaw���Ă�����R
A{o��׷��~~�@R
~@���1�2RA@�(���#
H/9wH)2!L9�\1����P*s�bA`di �����޺���.�\���#�O·g�D|	B�,��;���~�������R>���۸
D��XW��CĂ��� s�ZL���L�����y�=��o���ﯿ����;�<c�\�1\�nm��u�����n����;b�-��M��~�Y�ޟ}fO�_
A@ݢ�Q
H-�2�S
a�r��2RAB���'�\�GNe��+���w2�$�i������?}�}]�s��H)�혐XH.��Q �C���ď��*����/��w��^���n$~-���~���e<�<�ǴW� O��~��Jb�Q�teá�A���y}H�����K�کO1]g�Ӝ��/��p�����CL�� �d��K�§Z�7�u*��� 毐2Ed]�j��4�>��=��A-���,�*�e��	�6��������2����}�d�����[�a�̚S����l�{G:j�r�e�w7�.�/iڹ�5Ү���m'���.�>��j�~�wj[�E�n�R�Y���h�����qMm���y���[��W�d��(f�PO�Y�[������ָ����5���٬���h�m�N&�뚱,�i���)��pDw�^"{�,�J ���W��7�
Z�>��&/.4��٦�dI�%�r�h ��B�:�~ �%�K�J����ή��ŋ����Av��C�ew���sex�ݚ!l	%d�wn�������{V3ݢћ���\Dwhp��/�+�C�F�e��<�"��_n@�AƾFH�%����k��s��/�(u�~2K����{U;�س9��i��>�[-PџPύ�� ����P_d_ d��*�pl���V�PO+5ȟ�;�H�G7i�^�߼=��~;�4D�%`?Is6�M줽~w]Բ��Ɛ׻��T47	��3�ѫi{����:՜�)]״m�[����F��ج5@ʹ^
�ug���}P��Xx�Fٵ�+͙ڌؙ�=7*�&G����\�n\󶞕z.�y���=�(�i�x��!�5�^K����S�uv,�<�$�t<��6��f�R�cLK�hKu�Y����Y��ˠ�x�B �X˙c�l	Cd�d����ʔk��Xٸ1q�2���݈
�d�ݹi� ��D�ҋ!v���6�4�&1m+Մ΅�@Ik�=����e��mip@�2 �f�����Qî�ˍ�v���+*�n�����|��ǭ���d�Ad;��E�1iw�w�Fh� 'n~w� i��٠?%"HE ���w<�	YzV{8X#���X���<��\'��j�Lfdh?x�A�Я�QW䬹��x�9��>(�����}( A�FH�D�9Eeu�g���ft��{��,羠O��� �<�C|bT+�H&��Q퓒l�?/*wa0¾ιHN�<{q����	����*�U'�`�VA�C�@-�`�( �P�����B�}��v���]�ۯA���rX�%#�0�޽Gױ����|8{�%/����l�A�\�n�E�S]��WRQ�BR�n��l�c��5�=}����8����iD�qpzz��x�0#������m�򀌔q���!fJD+�{o]x�%o��OxnD:я|�pQ�Đ4Cu����.u�~�ב��H<��"�K��p��k��{l�����-�d��l����$	$����D�N�g�uB�m>�K�b��f�@��Au�#$^C��&`^}ph� ��	s�����$������1<��v���ú�nt��+�~,��o�Y��("$�,Y���,���A~_#��� �"���������o�^��"͖�4L:���4��?ޱ`�H�%A�_�Q���Xߋ�^]5S�xS�=�&�i�X ��D���+"��ܧs���o�Eڰ��B�V��RҸ�l x�x���o&�n���i�˪N�s�x��Y`��c��*�m�f�K�=�i���HA�^1��T�q��}Ԉ ( D�ł�����{���4��o��A�����E��\�z��i����dI	C��y��'���A�ڶw�X"n��Մ%�^6�����Q�E��N�l��;{��{FT��<���K�����cjP�u�z�[�[73������Y�CļY�ð��M��7�ol����g����J�%Π@;�8���SD_%"�6��ٻjr���X�����k��'��pyu�A��PDy���5z�Y��PM�@2PD"H����F�}9 ���׮��
�.º��w��~�"$��Icr����?{�F�m'톅��n�cmr��z�wg���o:�x���r���/,Eo6�WQ�(���c% A��Ag��W;�5���s~��cm�`u���n�F�@�_ [��?H�IH�d��^>��~[U��������P���f�q[/=x�1~��	́?������k�1ғ+��>(���T!_X�hWZ�R�uר�h�[p>��nc�h#dx�yX!��C���}%h��i��V���]�ٰAmТ� �>�kє������P �$]S�V�m�U���]D{��'Rª5��7`�)U��ְ�^y~t�-Qc�e��>!E��K�o{�U�����c}o��{���5{�$'|��{��{�"!�#$VAD�M��Ͽ`�j�o� �X�]���W�s�}'˯� A��2R �$�~��fj��|���n��}]e�:��ëca9 �e1{ e�ps�LdF�e��ii����iz��F�~}:H��$���s�q��a9{2�!j����/l�1g�h/�g����K�J�AW��z&V���������Y~�A<tϴעq7�s_��W�B���FC!|d��R-�O����#�*����Ȁ�`���X����w�R��<r��N�u��>(���2R �a�E`P�cv��ư7�$FƑ%���)z;Vlg��\N�
����z�T����w;��,��w�`�բ����`�V��y�_}`0�n�t��U��S��K���A����X ����H�T4;극���%�i�Y!�C�v���ܪ1VvЛf�=չU��s��ZhYs�x�bݾ/jjN3��䲥^vO����]�M�w	�k;Aj��WX�}�7e�.vL��r_�M���+{�eम�8�=T���7˱�v�"SNe���7�4y'6@fD�Eˤ������7�%1��"�9��s���A��=O���ըJ�f<]�ؓ�J�]��NuW����I�i���\�펵:t(�U��L����2K�w��L��8�e(+%��v<[�vo���
]I�:�X�}�[l���۹F��IĲ�M��2�.ŮP��V�mu��c���]d��p�l��^�_;��ha��o7%omu�G��o^R<lq7���r��=�p'f��e�Z���� �sjS���A��
��������]Y3T=0����=d�'w%u�ٹ�.0�0Ǫ��添1w7]�Z͗z�6��<�d��X�I��o&u�Sb�}zo0�'*'��!�/e�bo��o-of���e��|G+����UwٗHG�����Uo��+k�%J�o��P��;�;Ƭ\���A�q�W݋v�J��IӰ�۷z2�o����3/�u��'C�+)v�{_u�=�t6�ƶ1�X7P<r��Wt���o�3/���M�u�D?4;��oý����)ަ,��k�re���W�/�ȠkW�^f`��Y�6j���+ɨ���S���3{�6���Px�w,8��Ƶ�U��"]����q.�R�KU󉍼\�Np��Y�B�qˎ��¤+ro*/�	�A[5��!��(��m���cQ��Q�6*h*�V-m�5lm�-�m�lj��-j5�հmQ�*��5�QA�Z����`
 �Ԓ,� ��w0���٦��m�6�5�cs��j�P���\n�;\]�:��śck2�ɳPn�f-b��f�Q��Щ�9q.�����>�&9���ݬ[��0Zp=�,�T�t���L3u�
�U�:�YG��K,p�W�0�p�wNj��� ��������HCE�;�{`�0��یd9��X�䊹�+�]7C���j�{\�WG]s����T�ۯnA�MM�l�S�k��n�B�3q��W9�0�3��l06�k�É-q<wy7�]�	{l�Ǣ�9�s��-cuGz�M]�X|�ښ%%�K܈m"0L�vc��h�VYuX쁤�Y�t�kAP���p���l�\C`�k�엍��4��X'fפOfnk�-.<��"Nx�h$l�@��}d�2ұ�c�(K�l.��n�GV��̇,aYa�m�)��B�a\�*�%���lݞ	�rv�6i�p�`��$�3���uJ�fi')��
�)[��+Im]�.�,�XJl����V]����!s��"�Y���44D�ls�:m�Q���JE��6e��Zƀ5n-�`�����c1�D.l���H9�v8��gs"r,[�\�
�ZB���1���G�M�YFͣL�:��	e����Z�Kp��acc��v��ەu�C���v������B��睡]mN����v�PΤ��Klq����n�e-!�'�etq�թ��ѻOv��DݹT1�0mC��n
`�E�L&x�ٚQ���3x�˖x����uZ��|����ŕ��3�������6Z̘��,�m78	tv��rX@r�vJ��P�m��v�-�����f��6���b܄�8�\D�e���D�cs�)r�fY(J$��fJk,�QŐ��GD�쫑�ڽ��͌d��1�[`D�{p�˦;s�6j��rv�n7�n�XU0�8����gm�[��؎#\Đ�E�&|g��.e�v���0c�����P�/Wf6���?�I:wN��G���эv0ø�s�6'Q����.�b�ζ:�s��H�͕n��Ft���]N��1����6y5�7V��W9H��{kZ���4m����`:�ڎ�/>�O���!�J2��Ua1
�8e���=��y1�7`�nN��:���^S=*D�LuBQ�.A��aE���u�D��!-�ey��ɯm�5�Մ�g��R.�{�?C��`�Ax���x��z.�Mu�C[��x�⨺�c.�_E��C�o}햚�/wp���j�9�{q��s.�F�Vc���Gq+6Xy� �?"��)R� ��n^B��n�è{'�J~�|����j��ۉ�B7��yX ���C'>6!l�=L�����R?3�"Ib���� 潐�ܵ�A����O�V��0G���>����"n�i�W�����~�uT� �� �"z�B9c{=�����v>�e׾ ���5�yO+���Wvj�/�ΐ��$_IC~ ��$C]W#��zOƂ��j�C��o���u�A��d?PP$��/�z�H_D�t��Vj�]�p)x�l6;���Y[(]����J��hZ�2�{{��,����
j��I�O��Sm�;�o%`�p���<��.����6�����d��PQ����$�zۆ�o�W�y�oCT*���U�Sn�f:�����]�q��U��":cҳ#�y���������nZ�u���|6X�] 6�_��}��7E][�$��� N�oU
���X�>��D@��ޠ�|��+ �k.?U�����/,ڼ���.jBE�}����IK���2R ����_��,�> �ݱ`�ğ��"���gt���%��E�{AI�<�;8hά�}t�\?w �!(�� ���X!(���W��ƺJf��7B���N��Wo�+c�Q�� ���) A2PO�osn������~��'WI�jMe��5����L�uų����~4
����l��Ϩ	(���A�ū�y{r��ϯk��̫��7�7���e�'�Yiݫ���ݠݣ�}t�:���}��1��:ϫ�$�����A@q|��Mٙ ���L��!�@��-�d"�($�'�d�󿥝�k�`W���֦��:�fr�S���֮��i���ظ����;��̔C��ib7�~��c�g����<��6�Cmߗ}����
�f��fk�٪��Tq��~ �z���%d$��s^7�}���j�Y�XB>�V�O��fr��{�A�B3�7�@ �꿈�bz�f+���o���x����g���аYZ�����4u�7v*|������@�w`I��))���h�{���J�J���%F��M�L:�b@�-�.�K��c ىZ�&xͪo������YaN�?nȟ�J ��
�wўI��W��lz�4�h׈����N��AТ�I�(�	)R�)��
�5��Z���9��[G�v��v��$VF�K�+ �<���+��=o3���b�z� �q���*R�?%*2/�k�봇u�L��~�^��>� �_#W�DRg.�kێ^�W������ԏ�%B����y \һ��1��,�7�2���R���n���6\�t����ڪU�gq���{Gc��W�޼LϽm�v���A�]t�s���5.e��������~>�Wz؛��M�6�.��k׹�>Y)r'�m��v���KOi1��Cw���l��nTM�Þ��lRSN�v-�$� Q�n�X��	It���f4p�c��*�0���JXA�t-�ޏd���Rt+�I�df���Ӯ��l[?T^����d��wEPd���{�H H�"��A�/���z��àx����X����yibu��Sl]Lh?3�HiH���$^�y�A<l�;złgP_D�BH���p��g*m#�X�������ą�q�~-��`I	D�~IH��O�<�[/+h��ҁd��
6$@)@�o>ݖ7]�\e��~��	�P;{��̄Vߗ���� ��V|AH����������c�s۞�����+c&cH%�-*R� ��{��TR�
ߙ*��L>4}\� έ�c#��"�>�%T�흢�ڲx@��`���s�U����,Y��޴�'��"�CN����G�9�����i�|r��gI���D�u%,��;�tS���Yz�69�g]���Q��h����2����	Q��nM���N�^[lєE.��V��s؟0=z逺��^":�]b��J5�:�K
���ke汃M���۴F��q�.L���<'v��z��[u�j�%ڳ�v���Nk�6�ׯ<��jm�v�j��GQL��_Ap�C�{�!�o�k�U�Sa��T֮�B�<�pgs6��)�m�+m\s��7��y��Gx�FH�%��;���y����"����vGr�������3PDzR?%� �O�(��Gp�8^�����d��{Ըzy��8v���K����� �Ctb�O>Y�+�n�|F�-��( D��Iz��<�o��ח�ll��ݮT�*�����fJJD����.���R� �z�@���"J�a��ٖ�,�F����+vh�c&)�`����P�^��2R �% �CL���vU�ȶ�=�;�'�g�{/������O�A\_#$V"E��uh����KH�G�� �k(�[6st!;H�3)�ۥ���܁��|�{�[���Y��'χ��J�^��75����F�
&>6�TUeL���w�] �nX�:�FJH��d���=���c?9)����ܲ"�O*sWQ	fk*����
�5?��!K;�������a�t�ϒ��3;v�/mM�؞]�}�����[����4����a~F����A:�k�	Ȓ$���P��������F.�����:�"H��%"	���~9�f{���Wu���G<���h�v廻sv�ɻQ4�ѽYv%E����#����U��X��x�&Lo�� qu�ܿ�x���j�w�X���.���-�/<7�L��c�A�z����>��3��_�{����.&�X�wp�i�7{�Yۺ����i%B�ӳTR��j���Z��Uǰ��z-�ۍ�겖��e�QE�lf{�N�����J'��(wXf���,)�C��zD��ݞ��o��в��YDR �"�;�n�K�,Y�:K�������l�����	���{�VU?��Y6�uE�ȬdC�Eu�:i�䜒�m�_c-E�/i5�r���{2��&A��h�G/�������U��
��-�� �nUX�]���^�q��`���}���lz�:c��P~F��������� ��A���
)D�E�y�[�!���]�[����	׺�ފãt#.>5�A�~?b2"���>��W��٢�$%_#$_IC~"J��̪QV�|�fX���ۋӮk��6\Lh �Ι �J��0��4B���R�P��I yV�y,^sp�%����C�3m�Cqr�-���Z:����s����r��ݼGv����z���vC�B;�B���ì�(#9�e|G�K�J�2P�sۘ��m�²$J���_��xh�ŗ�X ����"r����Q�H�_r����"JG�$�7n����I�t��gF7ml���A��Ⱦ���A$�`�f��=�'~��@���/vh~JD��&��}�A�Ϡ���	׳Dc^j�����V?�k͎���7����M��U��wY�q�ѥ�6��4��8:�:��k�ɩu�7<W��4�c�|$��F� ���_�JD��D,�[�D]M�0-w��?����=�gF�Q���ް~>�H�FH���d��VRÁw�2<18��8��G��e�R�����Ka��q���E�3�����F��s���]��J�y�_�:V�λj����S�~�c7��_�"��0{ږ뭉��v����En`2��-�d"�tj�kcw<��z��n�ND��bu��5�}��,�R �a��X�% A��]t6����[���7�/lm�3:�=_]g��OJ�*��+��"F%��@���x�$�3P�g������^����sq��ǽA��n��y�`�[�V(�J ���H�{Vn�X�ٛF����s�;�(�ʝ�of��ݫ�I��s�e��r���&�W�Z�i�[���~�9�j���4��{�h��+fad�۪��Q�ֱ�UfVs�ܪ��.�;����~��X\�к)p�=���@���H��[�f����f��J�a�f��q>���Ns��f;^���\���H'2.�̅7f���30�L�7n�����+�m'�9ی���Z�v�E��%����鍣�s�d6Iv9����{,V��6�mf��N9s���&�Vy�w7qR�H������fE�����6�-ҁ��i�a��~�?+���p��f�f�봁�חlً��(s���p�[��#ͭ��1��\���v�F)@���R/}�6N��Ï�Ӵ��	�W�ޯM�ԽC��1��/�VA�D�IH~))�Fg��e��0o�k���F�B���]��iʹ�z[.*>��AJ�-�Υ�CO�A7%�'�AD��d�� �"_�ʻ������j�7�v�Q��A{�ȝA$�Kd����kv�q�qJ��t������P~�ã�\�Q��P$�b���WUO���j�È"$���"�*�!���T���>�v/�"�y���n'���qQ��A�(�	J��}��dy#b��Ր�A]Ւ�U��6�Hqp�o".��`�m���v�n4���,�=����C�$_\�/�y�5��ջ�X6Ƚ���˟��Nlj_�D?R?I�d�A)@����9;cpo�Z���u��Su1X���r��j�v�g7���Ȣ����L��޺9 ���&^�VR��R���۳|��  
���zR �y������,��'����@�P$D��d�P�w˹u5F�Cv��3k�����D"J_��X�xi�Kw�����IF������o����H'v�C�I[��J$��(��Җ�1��U�������dBg:&��zv�άd^W���@f�sy�{~�/՟�D,�K�J|$�,�ZkT�kc"�!���T/�����[���4NC�����J�$_#$V��MyG���ye�����<���R��ͮ�c�����u-cu����<z��{kJ���uqe������e���J'��
W��l��~o��QQ�4r�UV�
'�P������A2@	)�J 7�=u[�X},|A͑?+܃hn�ɧ����h ��h���%vH�Nk�=�_^Ő@;�$��J�J>�R���͇[�a�j�EF?+]UQ�-���'<��he�3����c(;t�/7l+[JÄ��u�Av*���;u��>��,d���z7*�mGkjcL:�uKT)_f�O.�v,�r*���bA%]�R���+9���6��mmm��4�ۥ����W���ȟV�]�=G+��·���7g+)ӷ)�o1�ً2t�ջ��^���+{��+���݁�7g$]���I(s���|�e�����U4�;}��˞*W �ljx0N��r�&����^����Z�l���\����P��ᩥ�=}��i�6�f�o��J������L�pX멇�p%�V�cS�Xw�]u�,���#�p�Žx��"N�7,��Sw�]qOv�u_8r����G[ǩQ7=�&�gR�.(�paH^]�C�U�f�ڛ%ȑ�T6�^�{�M���[+]��U	gJ����UJ^.B�_9�u����ig�ݞ
�VQ���T�;Y�+N,��[���GP�v;�rK���	�vj��L��]hjp����;;gQ�*�Ĵ�*�L�ر�S;pdQ;�B���&�}/!�oE�.[������c&�u�Ve�F�x���\�;eߞ����:�����Y�;m��k�C׽�v�e����7��/�K1Ȼc�R�SP��R�y���Hs.�[�ǬvS4��1�0�Ά�)�*b�/�2j+�e�o;{/fԬ������z�܇c�y�7׭����������bj�ޖ�TI �lR�Z�g2�,$�
Gl]���o�o��~�=��@���Qm�j�m�ֹ���5����Z�Z�X�mƣm\�r���4I�*�[���������ƬQV��ܱ�n[nQj-���r���͵{�R�y^�7���������� �"H��� D��8B�4�j- �6�H#I��T+뛍�Em�jt���������?o�׊;a�si@.P_�_ICG���S�{q!Y�r��o�h5��O����-��A9J?$���p�����TSD����c��ӫq�H��{u��@��ڀ���C3^;y�2�	 �mТ�O��N��5�WZ��	u_zjB�)�0]�#%�6�g�~_#��`�"%#��_�>#i��QucD��7B����͋�NSw�l�o���A��
Q"fS��y^ePF{�O�� ȾFH�%X�a]�tD(An��t��"��vhNB"JG�"��gx�5	��ݬ�L	��܊8�A�=�fhm�ζ.뿱_��s��~���x�n�t�䎼Y՘�o�Oa�US�Y�6�5Pba'�]�����q헵ؗ��{(�}����Y�;E[�	T���U���������������,Mڰf���v�v��� ����P���Wv�k���&f<A>�C~B��� �%��'|����e�H�O0#n�6��� �6�v�����MT���u[m��t�=z�ϲ��F������D�(�
���;��\l���!��0E*���{Y��9��Y��H��d�( A��uIt<�ĝ���~j��3C}��n��	u_zkh�I@I���A^_��t�A D�� ���dI@IX�	%��|����r�C8�m�ڸL�h^�����d�~��"H����خ�dk��|�J�4YZSўt��"�A��#�Z�za]��ʳ��ڶ=�p�v��� �%�2P�b^�ڍ������w�x��b�X%� �q|��X��YY=�;X�/�W�i��U59bi�D�ؖ9i�OyɚQ�[�.��ް�%��9�@椏�a�龯Q��8�(^�FN��~��|> �O����uvt��*�=v=+m�W\�V1�;�p�m��<�D{%v9��ܾ���g]r�;)��e�>��g�w��6�vQ]���؂�/]/b���)�D��f���fև���ȻRXL츊Ji�ݴ���͖piL�c��8���q�O���<kd*z�s��^'n�pn$�[Yn�_(��{]. 2Wk�,�$�{�����y�Mە���]q��)�V����0Ց<�m��/q�M�|���k��s���v�~IP�~�޽Se��[mBfcH����9��T �{b�2R%D�łd���\z�z�˯��E`���f�nQ�[��&�\}��4��	)l^��#�ϸ�ŃҾ@Π�Ib̔�&J�ع��9]�:�ڬ��p�����W��PDE��$@IX&郰W�,U������~�X�����]�N[mBfcH%�	\�⮚����_ {�"$�XJ�"�|RS7;[_@ϷdHZ�����BPo�z�A�n��$%�$��1�QQ�j�w�qS�q�T�(��)�m�#զ݄����uy�eU�fF9���"#�����p�v���㪝3�5���֊Q��h�N�yE��-�v�n�`��`�ؾ@��։ק��ٺ�r��w�=8F��:{LmY�k3��ò�������׮����qF��`���NN��8��I/����� �8��~�޺�L�k��q��h ��A�"����s���2��݁`�gP
E����Pܽ�¾v:����6��z�4n�~nD��?�
2R#@޳�|4��J�f �>� ~n�9��*��EK��p@�:��vWKc��|��� �R�"��"D�I[���:��R����~���؛�fc~w`H���PP/<cw���=��|�GOg��̶Vg+��)�];b5��3óe���	�Z0���stO��Kz"G��@"�A �_�H;˧�*ume��!z��I�)��f�U��~�A:��H��)	�� ���nv#
��0si�P_{7ʥ�ft����Wb���A|A���2E�������oW�{_/�?/����($��T'���ép��R��N�'�����bN�7un��t��:����6;�zc��YCd'N[�U�Y8c��R���j��U\����]��{��I७�&^3��{��ڸ�wh���0|��V�r�6 H ��~����"�^�M����]��wo�=�"�T�5�{X"�����,)A��I�Uf�+cJU��L	���aӚV�;�C���5�	�PD�_ d�� �����76_�{c��x��[����7S�zs�ڙ��]����(��l2�m�	�YoϿg��d�(��IP�^��5७�&^3�i�T��WG5�ځ?S�sbA� $�X �A�I+�b���٫���l��:��d�f�Y��J{4A�>!&��W��/��ԇ�u|��(�"�J�Atxʮw;���)��N�"���`���h�Z�;�x��\Mv��;�}>��������DC��$�w�G�f�Z�be�1 ��@"N���-i����uҎ�l�*�R�2�%ތ�����t�3����E).�W_7۹�Vxӵ7 vl�����X<�!�w�������p� ���+�J�B(�%4"��uf  {"\텧l�y�Y!٨oc��~n����RT��L�Z���dZN3x�A��]�LW�۷�SԆH�e�7�k2�ʖ�3�*zv����ڴGeӾX�_�Ԟ�a]��<,qN�CgZͩ��W�C  �/�;ܬ�D��$VF2���Ժɲ���m �ް�������L�f#~?k�$�P�R�Y���E��8t��_P	��$VA�D�z3�1n�������y���p���	��`�;�DIH�$B̔�]!�b>�����i�ذd�~�����B��|��k��y�{� DUy�Tq�5Om���j���)~2Ed"%,�煙F��b����pн�ch-Mbe�1o�\	j�� &J-��~�嬸]��t���){�Y��ˡu��g]:�6e��V�/T�ׁ�	%�kv9����M�,�<�f���������v�s�u��%��s���R�؈.�"��`�B���e�\�3"gx,&[�����g�m%���mH3F��LbK..a���C:�R5����ܹ ���8�MJK�l0�V˲B�. �1��"�)�͵�#�)���'N�ݻn�l���ي���1�Ӟ����-�R0s��m�@���!��7nGS�g��u�բF��c��T�B�5�'���|�TŖ����`�[i�W[	�:9ꕞ�3�6�Z�Z�AV0w?X �P_g $�H"D�r���M�t3k�w�_���/=F���A�/��	%�%h �("-��{SP�v����9��2P^��OwE={Z.���<����~���c��|��E`�( D����%����U�u�d�!��s�8b4��� N5B�Q���O�$��z�m=ZoN
M�s���+ ���*pq�ZS�5�?�~7K��8�F� ��X�%/�&J�"d�a��*oj�(:�񭠅���/wW�<��m��u�����_\�{y�._�z~����e����6��崢�6���㋩��'D�X�AftV<�O����r��`�x���Bc��WbՇm�A�F#H�S���:�����j�:�|�"IX?( Ecc��ҳ����l��\�B'�:\���浵��W��ͣ&Rt����B�ԛ�v�<۫�&V��`����l֥S��`�`����=W�P�NK橏t�/����^����`�܀���^����6�o�2Ń%/� ��	"�� �B_��.��x4y�^�Zk{9�e�അ���� A��� ��$����z��c��Β*�E��H�~rX�������_v��(���ث3�\�+�4ȐE��q7w0Gv��ۗݾ���v�)v�F=t/����']�"��*�f׈&w���IH��ǍJu��k�[{��%c�03f���r9
3���u�`�ػ����F9��u���\7��ږQ�4{�{@��ͯE6"���@���n�Amy�[�%֟��Z2 ���2I� 8�]L����N��~V��C~A��#~?ifA[T+�C�J��]ki���b{���y��Z���&�b�+�yK�o0X/���{���}�v�rvU*I^�FQ�^��p[�D�<kK�����Ⱥ�m$}���󨽞.�k'1�T��ٗ�ܜ]�"�w�P&w��:�"��"���;q.���6a俺V�A�w��]����H��X ��KR��p��XD<��F{�X�� ��̆�&����%]_c60�����f�m��zn��W�^�l��nڴG]v�S~�����W�ksW��X4a0������N�w^�Z<n��3��A�G���7D��K|�H�����V"D�kQ�:/l��Х����<��_��u��ػ��D1
��$�fJD?gPfjU����`Π!ヂ��/����Aդfjޠ�g�FH�Ǩ���g���"��K�dA D0���X�5��T�[�F{���M5r�S1��t� �mW�E�AE!%_P�#\l�{S��A��'�f�!J���"����D2���+ ��Tyr���Q� ��S���qސ�W���8�i�ޣ���=�n��z�%�֋�z���ܬ�[1ȡ�wJ��ޫ��"�\�u�)e9�{S���9b̔��)�X�d��5ƫ|U�f ��T�n������z�����	��_P_"��2!�_����Sy�Vj���fͫU묹�9��6���a���k�<%�)�9�u��%A��+!�|$��I`V%Ok��W=������,{��TQ�AmР[� �a_$�,%C�f>��xF1�޵d"�:�N�~�}���Y3�����n��y[�cC�G�0�D�2W��	7�J���v��h�{���i���>�����A ��%�Nj����o��ׁ8��?$�Y�"��1�e��M\ƐA�̂���ؑĹj�D��`�("�B2E��iտ7��l���~�켂呥�
�;��#����,g�ӽ#�.�MmU�'ssړ�9%^քkO�/�I;�����P��C���Qo�ڝ�փ�eg<������sk8��f���a�]�y��i�h�u�E��⏰/����'Z��A�WذQй�-vgč{�,ڬ�Vi�F�����n�gK�W.��2�甑N���غ���]i}b�Ŝ�{�ط���ǤVM�w��l���%T�i���å�̚*��᥌V��T���c��T���)K]aI�ų��u�7t�L�\�K��Gs������!UI�}��)��6�W�K>���(Mzd�*���lt#
�w�r�,1.ʻeU��_o]��[w���F�_J�lRp�emحXR;����e>�T�]{�ۙ�>��R�3Z27:I����M��E�ZgE<�֚�3v�R|�U�ed�;�K�j��5���ٗŶ��u�G˹K�5w��{�Jv�R��Kn�Cx�)*�(�;N�U�0k��vӫ��a�Xkq��p];���h=yO�����ܩ���=Gr�uZ��x��FIr���fM�p�vw_��L��&7��w�6b��H:�&��*�=��w>����}N�ڧ��yƫG2��=�Sh-߮�}�P켣����o����dN�"i��`�׏�%��>i+�2�;i��3��i�޾l�Ź|q�șͮlY��{R��yu֎����������!#�//��;��Ft�顚���T�0:��6��p��gEF4�k��͛v��qwL�W�Św-�����J�:0�h�c��R�Y�����8�Y JBS �M5�-��UsU�Z浹��V��ܫsj5k��RZ5*����cV��͊�X�3�N뚢�-cE���ƹ�E�/O_~��+��:;V�\�$1�1�j:��]�J��� �z:��C�`��N��Zx4�n�ۻ4z�2¾��s�����l@��˺�M�b�y̻�om���ܳ6��P&�A`:�e��$<�\�ع쓱*��'[��`V싼G%t����';��=)`��3ͣ���#�l,1$�cr[9�6:GzRWTm\�6��ƞ��������5�pl/:t�o<q�9�m1�����uX�7X��|u�Z�Z��[���)��چ�(6�R��K
�C��mh��e�i�]6�2�`��vzJC�����vF��i�:�XI��iSx�B��m�f����6#��\Ӵ�v��h`��=gn������n�Jt�&���h0�݅Õ\����s(��X�@8;4�t5�l�1XKs���S���s8�:�dն��w�Z�&T������$���9�7���,�"�ͺ�3֔I�a��p�V�0�lGn�sCX6�v��J�Ll�G��k��犽�qK�8�=
L7Nl��1�ܷhf�"M[X��A�].��p�-��1�8V�-s仈ʄv����!,Q�`̲�xt+�l5V�D���,׉�)�yl.Ddt��{)IS[�au�l:�.��k���d�<�ڍ�ap�
��u��8\:��Xltv�鹫�[;[����lh7R��*C��	�Z����sO������֭��G ��#�cB:���XBy$�E�Lu�]�9K�c�;��U���۰�	���q��aM��I���-+Iq����J\\n�ݚ-�v݊Jq�!��`"G�=к�`a��o�-��s�z��y��cxr3��1iF�X�kB�	˯�T�w!Y��A1�*��E��t��uE���)�r�-�۲�༨p��;-OI[�r:ku�]˷v��ln�]�1ą�<v�i��,�0ݺ��!qd�m>�rKG8y���ٶ�@����\)Ե��A�4Z���ܽvN/N��ݓ��R�ڵ�#U�p���ۭ@6��]�
�^��ˉ6r�&p��9�B�CXQ �hl�怭����٤.����[;.�a۞]`ƶƐ����6ь5��Hic����Ƒfd�m���Kss�mn�窗slR�;k'X6Ԝ�qb4��{�.z�q���p���k狁>[@�1�W7]��~����[��Szv�.:nv��t�v���ir�Kax8�΋�\Jm�~�S���c�R�u�;{=~�-����S"�}b���w��3h,�.r�����b��2E`�q���y�j�GX��[B����e���.��J�A,�!⯒�j�ⷢp��7�v=("�~r-IC�n����uՇ�O'��QM;s��@��VG��C|D�ř)�/GNvt/�?1��/�%|�0�������չ�o��dfo�ޠ���y��[�ܢ9�V>�B��+ Ȃ"�Y���5뷾?h��t[���z�{�������mH�R� ��EZ�xL�g��	����Z{��][s�iMx�*]
kgyc���&HЩwM�]]Q��R���}�L��7�$��$A�y��_�5m�?k��kU��t���������$������4��϶vnɜ�1��k�i:=�9�oO.v0�Ϊ�*�_-��Ѹ:ڥՙ��$��r�=�����_V܋�f[�}�v�]��VСYs��it7�4<]Ă!(��n�콹�nc
��.�E�;�$�q��)�
>�5�$�V)��c;�,{��"��ۅ�wp��{����W���B1��;���ovt�_x�AzX����"J@$_aɷ���b=CH'�Az+ �_n�󭝞N��0��� N���*�UT�㻭ڞd�����]��a��V!�V���J����
���qVQ�~��ws���#o}`�ޠ���2Ed��}���>�,���҃ s����ٸ�1���\�r�2��lL6����ν�������}"A��>?$�P>���bz�.�+祏h�Ƿj��۶,��A0���~	��8]��� 9ڬ���������Av���
�+OPDC9�G�?�e��;ԁx��K�J�	����½�3UVS�px��n�p��v��T��X��ې�Y�䵪�Jz�~T��4e��+�ᡨ��M-���	&�;/J���cG��Ky�cw7�IK����{��q��D�"!�P�	����L�����dG�%_x?{��y���o��4�t�DW�mf�]�{F����a�$�`�("���,�:�S	����&kp��VE�o��=�����J'��I&�~�'��x�$Cd��j��\�=
!�04W&��.���.҈�	)5���C��{I�7B�J'�~J��y�d]��iD������z��g�,3��H���/�����G��+B�d,��$u��� ���G�o�mó�э6���H']�%�2UǦ��]��'�e��Ө A�FH�%s)&:��$�n�Nۅ}�ȳ��|�~��Ȑ��,�ܛ��JV��o��s�"3��Y��a_r��~� �7�\K��C����|AX�
����XIm��Yi�D�ъ��T�Sk΍���k/n������ۖ.�%����6����Q�9���6ڲ'PDC���� Ȃ"6�;����N}�h?����:.��巖�G��ӦA��(�L0����YU[3�A���а���Vw�L!۫	�����\h�7A����\n���Ҽ�-U�^�Nu��$�����7�J4��#��d�S%�/��'�3ʾIH�R�����轡��~Q�a�	��k���������dn�ޠ��2EV����u�A�1P�d��r�$����?%��}y�1Jx]k�� ��:m�Q�A݀$�|�X ��H"Iv3&����WQ�T�1|�>q_�Y�s��.Y���sH��@���de���T��0GU�8��d�AP ���E(����T�Mԧc�3�p�[������df��z�\BH����W��}�Ch�Ir��|nq�To,Ŧ�:���L��˙�<m�t���7��.���w��g��K�k5S��PX�RU�{�]�h�`ݫWh�ܑ�V��z�b�a����S0�J�M1��xm���m����k��d�ә�+�C)X�gWb��P�K��'��W��֔�ؗ �i��.`�t�3�f
68��ݧnl9rk��T�(�5]�rō!��<n���],щ���[RY�θ!��3�[�QҢ����M��IK�qh�kcx��0�"~����v�=�=[�5R'GdK���b-5ݥ��.�&������JN�W��t__D�C�K2�U�Ͻ���������{��
�j]l����dw�qݢ��ܘ.�{nz���G��7U��?8���q<0x=&����G�]����@J�F�Bq�ܕ�����E��X���dwj�]���{��܃�:�Mt6���-"�;����k�m ͂;�{!9�i[�mJ�~���IP��<�u�����:�}�塻]�C�[�W��=A$B�2PD"�$C͛Ue���TU�� �y�ٵ�O��7�4�u�~�����	+>�$�Z��:r�jI%��_D�]��E���d���c3��s� ��J�.�`��A_T��_� A����@IC9y���eF^���뽡r�Iq���A�ؾG����A%#��Xb����������m���J�{�L��V�j��l�W�W�zU�AP�Z�BmTv���J&v܃�YT+a�8�o�s!��D;kj��Ʒ5�ǈ�@/��G����CY���s��Kp$��P�R���w�>�P=����PPE� �yzV�;q>�<:�D�oc����+�%#��J@�c�������L���h�(/z�[��Vs7(��]��%8Ʀj��Qh��ڜ��o��X��q��ȉ�e��^�a��u�~��$��o��������u���������@��tS����?g�6��'�gs�&�͕��&�k��ku23.�V�!�H�t�PF�Q@�X�lv�r�!&_�����ُ]�r��}5%w���,yӪ{��I28�S���Y�=��R�sk5��de�9U��n㔓���{������r!%	"I�ǲ�s�����wgJ��C���K���!Ƃ�PS�ɓ�����T��9�v�B���9���/62��q�{��n����5�t<�{�v�~o�G���)"Y\���]ӝ�������bW�!�V��ڹ[�nʳ��c�اs��9J>�!$RM67��r�[t�ԼחnO[[���)���7�E#����n^�[X0��ta6��5�Sa�ua9��m�[�]��bѧj~��Q�[ҫ��RR+Ǻv����N����bMD`��y��r�"r!%|z�{��;~ϯ|���4�w���B�v�V�����+ݝ;�\Cޠ��$���C�2�����f�����]r����z)"�I_	"4�t��������߇�f�IO��o}���WMu�������ξ��7�ndR�C�o;1��}�&�Y��h�wYxz�:h4j��M�Yk�]ԝ][��iI���N7�=�(�"T��<��uy% %|���[�{�[gUPy�MU��V�r�ڭퟛI{����V����篾y� ��b�Cj��£���^��8얖����M�:���!����|��߿Y��	"��s��xͫ~�U�n�)��OwxR�"w/��$��%T���x)��{���=^9�l��]��������$�ͪx�mWsɲ	"E����������g�*��!.�2�۵Zn���(�I3�w��#{�������;�̞�W�y�n�[X�ƪ�1f��g۸7bH��D$�R���y�~���;�~s�]&����g�8�T�_�T�5_�ײ+d����"N��_]��"�ʽX���۫�Ի�W��-�÷��EK8D������f(��vnUU�&3�l�YT����H�j�jD���ڻW\mf&����QVhR�R^�����c.��(���oG�:j�`�U7��(ީ�h���w8�mE�PiF؞S��m�X�K&)�L��k��8'c��{n]�x.!�V�ȼs�M�
JZ[�����bŖm[f�MhJ	pE	\;f@0�QG��u�z'�,��x�����Y�Q֗�b�ks�-���iw$�+��V�f����cn�#�t�;�A6�KƓ
""�Q���J�J=�r�|��������SϑD�����33�(?D$�JH��Y�Ŵ�_[�����7�}ە���ez3��"����� I-�sJ�i9e�����S�I/ Q�y_���wW���~�l���I�:�+��)�>�-��IC=�w*d�����ic�[�n�e�1�U����{r�g����J�w�$�Ŋ�U����u{�m�ηw�wP�E�T�ݩ�j�w��9�֜�8�U܂�:;���Dn{D�̼lMf�P$�-~k�҄�	"���&��Y�y5y�Ѯ�F֕쏘��/�!�	$�~kƯ:�f��E���W7�6;��J��@�T36�.Q���9Q�{Z���"�^�YW�q�萠_��S"�����F�xzP�o��%�=qY�����M$_���B9Q�vc�w���͟�R�|�Ӻ�֭z/}�<sڽ~��s�O`�t�}�u�}$_	*%/��0՝�7Z~�$�{�n�Us��c�כ�~����[t��Y@�e��s�+	@IJKR�gN�@�[;�/Fn���Q��<>�r�uG�wxvd�V˶�d�ԫ��s���5:��%H�/ic<���
+�J#e�~aȀ���+�$]�k���NzS�3�=�ͻ�si���6 �/����H�E�S�[K'����A��#������UFk77�_�dBG�Ǌғa���x�j��9$��y���W�c��3{���Dw\q��m�窔�7r�fmd!ۥ�:n��r'�t%:EմZ�J�֢OY��q񺣼�����dI����h����Fq,L/.���D��:����ޣ��hz��[��1�|��]�z��&��Z.�UJ�}utw0U�n�����n�d4Nw�4d�*��u[�v�u���U
�zVY���w{�Ӧ^H�{]qP�#�Y*��h\*�Ἣ���:���(<U����-<��"���eޅ�dV.橌�[L�F^vo9P-�Y`74�`��j_H�����E��A��o�&e�a˓��n�5�[�CEP��si�`��]Y��]��sx뾼peB�;�:�`恷:^�륲ힲ�έ|p��RF�Gx���hN������tZz�޽��3�'.(uIg�eE؇b��V	R��y�*��'�̣�g�;�$�T���.�	��L�`����w�+v��0�^ �xeQ�wF�\��]���v{v�F5e)Uz�(��VeL��	�9W=�|G�\���fer7��2��u΁��l�Ni§]�6]E�!�+PD����W� ��S6������i����ᫌ�(��.�=��h0�>�	�6�S�s��Zw���"�TK/����[|��h���]�������K6��c��E� ;��z���$��p�}k��vj�;�@�J���Uq�9!�竎�3r�}f���n��v��٥i�����uV/\�%��(�|�����R�!��"�1@�f!Gb�1K7�˻���xN�S:{�������Y\�|�o�,�@���U�vF�c���nk\�c6�IQI��M����5��6+�
��b��*6�66+����nV2��*1D�%��Kb����Af��d�wE��Bi2D ��D3��%3f��cE� 1MjPlcA�&MIlF�	cQL�ɤ
I�1�A!E��h0�d��M��c b�
D)@��A?a'6�VSMϦ���In��q$C�"�N�V=^k�yV(/�Bz��-��w�n/Z7�;F����½��>R��@��>�90	"�JEB�
|��ջ�@J�ٲ�+�Ot��1��+T�QI_	&#N�K3�B�Ѫ�>)]��G)+Y���t�N3���a�1Hk1+�"u�ug߾��6�}��"���ֱ�/�ܱ\��L�7k�\����a��ފH��$PS��z1̻��ccׯ۬z�F�l�^��}�|��:�e�~���xW%�x��򒤋�#���y�C�َ��ݻ���!���}~����JD�}���-hׇp~s��<���W��5�u����L�m���~�Π� ��q�Ç�[ʸ<j�`pVq��a�d;oMd�d�5��J/6�6�z������w�z��T����.m\���3W�� $���/��J��Z�>#"%��{����Y�8�z�u�r/�ħzD�N��$��J�i}{8�CQ��Hv�zv;kr�O�	�kUj�F^l��8���g��S�I{ܤv{%�y�˽���{�Y���i�� �_I$�$��Ue\����Ṿ��ү�kX]/ޜ�,w��o�����Iy�u��_r�>���IJ>I]n�@�F�׮���f'�e��_��H��"�[�np�~Ѹ���]l��H��mOR���ξ�7��/�}���R�y[ܤ��(	$����fj����9P������~��/_F����>��@I>���̩����gf��Cdw"���!�<%X�i^�uĺM;Ǻ�u�#b{3'�Wy��z���5�u��ͼ�����}�bP[YY�c%H���d�m4L���fe���<1�H'����an��u�RY]J�.�k
:U�F� ����a���nk��)�.�)`�ΰe�\6e ƍ͉����69�,Cg����̋��R�n���:#��63{ lp)rn�Vv}k��UR�u�2�[0�5��G��W�G�&(�y��J$�#�Ua@б��魘��&�6Wec-5H�&^��=� �ﵺQ��B�1����J��j��'F
d���ѲEYi�U�����w)*H�3��k�Yw9��1Yz+�wt��U`�����(� $�����4���Y�7�1�T���volT��ȶD$o}^�~Ў&�ג7c����JR'vV��l��K��[S\�}�y3�q�}���I�H���|��*�ur�r��s�p�{=����׽��)�⑬��6��@(I�8��$��U���JK0s�^�y�gt�)���!����$��^��$OFJ�,!�hp@�7����5�\��e�qb6њ8,�v$#��WB���[��}_	*����]s��Z�e7�OZ��W(�M�w�����}$RP�H�9�[`�P�.�'��b�9Mך�(&D"=�8,>�h�u𺇳0�Uq���,��Y�X�7L��ȳs5Q�����Ҝ��;��v�݅t.���Ԇ孧��7ym�0���q�␒���[Գ6�렳��g/��`J�1�J��v�daV;��ۗ�5�o}�#�@$�H���c�ּ�*~c_���՛~����un˦�8��;77K�����M~�*ts�⒄���}'����8�����[����	�W�\x�W�E�[~��������B{��u��mK0EK,;��=���I퀭�l\��U��KU�̦�_�{��wkwnI16����>�F�֚�Gt���Z��߾�$�����T�c`e�[�,�7c��:׶�z�NcX�}��	�H�{g�p�^���))J IE�u�a����L�1m�^����]G�\֣"�v�;��x&$�����B��O�tf����aj��X-�~��I����:ܬ�Y�Se��kqs��snNS����W��~����o����V�н�lq��Z��I�k|�}ٽz������@�-�;�����/�h>��d���}$&v{s.��|�q;;�μ��&��߶�Cp���^[�&Z�������k�v�]6v;n��<P�lp����55�@�QVo�k��7��+�$]ͭ�]=G�I��i{G�Ԥ�k�����t��!%	"�I̽��թ�ܐWh͊z߽s{1_���k�	<�Ꝼ��ׂ���ߐ��BI$ߤ�;�ZU�^�uw���}��k�O����$@I�/�����0&y�$�{�'맨�ךR���kzr���&�(NF�W�:)TSl�J�G��g�|�r�RF�9��ZXݪ�T���r�����glC3f�k|��͖)m�9�!u%fr��{�_{���/����jG�����B�NS��w���ܿ�_q}%}$��1��x[�@ѣ\J�IZ�z�-�ͻ0Y��f:��b�v�M�Z9�cc���ϟ�|��)"R���w��q�v�E'���¼����_��mJJ~	@IHZO��ƏdUnG׻#^fT-n�z1[J\�N돾N)%���U�!�)+�"�e��u�R=#��s\���;s�<������JD$��D����{kk/�/�<���W�kogxd��nMS�{Z�a�'{���{+�σt�@7v|/26`�F*��&�{������u�����$��v����J`��gr+�.��͔2;��;���A����#ڥЭ0���X��ڐ�a7�.��[h���A7ݝ�O1}-&�uS�F�m?U]E]���5��l�d���R�⺷Mr�GO���^��N
Ր �L+��0�yF �!�l��L�p��ZPy�5/\��;��]�˫��n�z��:���G��8v	��KB���!d��=x�Lnz+�����6�i�;;����Js7�J�#�X���5t��XrX˫L�R�P�v�pp��[/;c{6����'�����ͥs1m׌�G�i�7�i�5��t�+0j�7fQ���?�O6�	�ّ�fLOu�
+�F�r�3�Z�������:���km�n��W[bM"�@+��ls|=�5drl�}�����|�2�*�ǃ����Ͷ��ބ����s��l��7�jI�����ݮ�m����8������_zh�C�_ڥ�ު�~��N�<W�;���)7NX���᭷�7@7_6���?�[^����`iv�o��F����ؾ����Bf���$�͵�l�%ZAn׳a�J�z��J�n�������"�_+���C����7_zm��w�Q���dl1R��VG�܁�C] �Ndӎ���Vz���Fa��R�e8I�(VgQ����_Z��ȞNJ�i���nWB�ۧ�}x�ӚU\�����9���ZC��O>�+��7k�ʖ{x˵�OK�|��z��k��=�FX�+욾�M�m��nx�X�Fz
�y���c�r{�� �m���ZBҮ���y�����M�~;ݞ�M��N�>R��3ܬmYk�݀�A��ޡ������
^n+��?.��yW��P�|��H�/kN�|<��KqU�2�B�^��"�� r�!٫���".� �b�X�4����m|��z��g�g��Iw=ǹgw�']Y{�^PW�������ڃ��Z�r���_��{5�;`��Ҿn�o��qe1�}Bo�t��w@�[���v����˅�UJ��N��gvi��f�9R���Y}�����W�"��g�^d�ϛOk�n묍Co�EC:ٜ��ovT���~ެփt�|�J����gW�;7��^�� ���uS�{;|��ql������m������n���h��y�ٷ�������k�pv��k�t���h��5N�����9���!�����	��GFkHb�1"\��M
�
?R*���H�t��hR��u��M�����߅A��\c������u|m����U��˯m���Ȁ�]�k�nk���cy����t����T��Έ̊�wW���n�z�^��z�%����k�pv��k�+�m n�]^�'�ߌ���eu|hV_7��%������������ܯ(�u~�(��Օ�/w��ܩk���iK��Wƽ�_ao�z�ա˭ѽEo,O��U����|�0����D�֋#�UO;jQB��X��=C�|�_7_|���fwf�ݴc	L=6�i��b��ukGۙ?���m�=����?�B�Ee�*�	S�Iu;l[����ڽ��웱K�fz����fw߳糆� �|��oo��e�]͕��-�}�eW��>�_W�܀n�n�m��E1YengW��>N��������;v�V�9���^6��u~�m����y�vs��w�k=�����w-��}|��A���ߺ��3��	9}����A޻�˛+��[^7����y�zT�x�t� �_7A��U�[Wݹ�\�\�:����n�J�g=��@n��7ﾳZ��Y���Ʋ�N�ń21S��;�ヹ���J��Fvt�V[��9/���+:�)`���앧	�Z��oW*��xV!�q��(��lp<\�k��˧U\�s��i����t�Z�p�3j�P�*��b*���V�?��0s���G�����cw�oo�#�YC�r�c]��6�����1�cs���Mt)��H���a���E�{ݕ��f��v��3f�n좭����[\��J�B���t���C�&��A*�\���u�O+-�Zy��+I��e�A�ꥅm}���]���䭾k3�����b��W1��{mi�U��T�y��4�]�m��xS�����gg:�w	�����SP,r�7꼘o;ȫWW�U��w�72ӛg���B�r��ަ��a�(T������Ęe�:.��{�&���1S��[�^��Cl��;��Q�Ĭ��Y��A{A�q.��w#3I7�ĺ���-�A�+�Q��6��f�8��wX�sU��wma�i��F�1,�=Vpn���}���ƶK���hvS[�]��(��Q�t��])]l'3��ղ7]���[*�������j��u�GٷŌ�e�A�Nt&�K[ض����Mj�Ƕ·���si�+�[���e8��N����R���:�� â7����pf�oY��w�֭Y�z����2�.�7��ӬC|Vva��fiu�w����rGgB:�m�}Z(Q81�U9hfs�řt3�Sw`s�Ikvahl��e�*�G;�o���'�EX����b�DAlc&�mBi0��MF��F5�ɍ��H�RQ!a�	0&�����F���Q&B�h��3$d0E2,IE�6"0$QEbDD"c(AL�2�6B�ThHah4��&��!�&I�SHMJHI��H�J2�!(���b�h�0$D`��(��D�L��1HH�Ra(��ba6A"��bJA4̡1"S#	�02 �211�&�!Q�� �`�Y��E$P�E�c|�uie,p�[�h��/!EٖGK)lbh�،,�D�m<���+��8�mt�z�u��\4�fGACB����D)f��:�%�X	{d�����<q������<"u�����.��ԇ%Ь]�f��&	m���e��X��kln����%����`���j� J��C�,r��M	�Y�l�ni<��'aړ����n�n۔R;1�X�����.g��k���70���d���T�!ݳ-n��'�qqc��f��f[t\Z1�5���XZ��cCE��F���Ep��3.	rB��y� ��S���x��
@��j�n����2��q���w?;�V��tsP���{t����v�\܆��)ю�:Ĝm��9�=�l�u����X�Vm�(n���W[Y�lm�^��<m�BU�������C���CfX(S��]m���΍:��9+gn׋������DCRY��rL,m�i�Ka�\G��w�&�s%�JŶ\�m���`�LsV:��t�S��-�+�����Q�;����F���F9����-�<4޻]0cnq;�;"W��p��@���\F`���Nt���l�/��j�L`)ɳ�-ķO��noE�l�.��lJB%�X,��\�oE ]�3�s�w]i�Űt�Ѻ�ת�5��s=F��{I���!�t�/f���T0Q\==�2i^�
���Kl*h:l�ii���c�q\[�9^Q�0����sZ�%ؖ-���V�f�k`nck\�[���qn3/I�ukS�y#�7Zx�C�ز'k�>�c�s�����%f-��b7�*�������kj�҅���c	�X��Q�.���Ye
T���Y��J`�v��G��j��hG�˶�;�l`L�_
Y���O��5�������鵚ܸA� ��v.;����0"��f�E ��o+0i�]70Ĵ4�b;�h�9ŴM�r�NZ�Sg=/n���k87���c]ۍ��j�2VW8B2���g1�"Y�Xh�Ɣha����D�oO�啁�#y��pE�Ɛ�b��;Ri ��h�c:6
�jmKbk�i���	��'����F�AB����0�X��cNF8�n�+�؞�v�Q���V��8ָ�.mvI1��;<�Z���d�eA4]qbZMn��LV�ᣀ��Y�_��a*r3��ڹ�۞.�I&U��,)��!�6 H�]"f�g�6񺛃���:�j�.[=��ҁz�ӛ�i��m����ߏ�u��j��j���g������,�x�h��v�w���7}�y�z��w������3u���ۀkv���-�����%gC�����n�n�m��b_^ڵ]���݁��{<��M����r�l���Lo'��~�{��}������i�O+�_R�^���=����}�*B�����_�y�u~~޻~~uU�v�R��*�B�S�Ǯ�kg�<�z+�/&��J���Z��=�������~~;�@�ˋ���z�c��)��Ք�1�����-�u�m7K�)�����Wۺ�*s6�|r���U2UVIw��`��S��E_zFtn�P��u��wr�vm�!z�&+F�ϴ���DdY���u.�&��Υ�^3+���F���x��9yv)�YW7��k��_6��ЯG^��=���Nٲ�/��[^s��o n���+X��׻�T���a��nw�u�P��]ا����W��e�J,���6�������מ��_{˲*�3_R����~����r�tuv��+]@�O�n׊��p�9ym��gi��uv�gm'#nQ�9������9��N��� ���xW�:�>�9e:ѡ{�n��Q��J�d�7M���]C����y�S�'y5��k��}R��b������m}�q[�[�=.�c��|� �|�_���j�j�Y���Yͺ��E�7D��򔯌vQ��ׯ�+�2��Y�9r�����>���9^�uy.�o������]�l�֚�L�~��v�$����i�ΧU}r9���KQ�̬O�w`�y�~��Ѡ5���܅*'d���͵�t82mis-�U���
��x�/F�fNdxp���(ɐ������pՒ�F��f�%׮����u�٧1���p
�l�.���Ri�<���|:6�.���t񺙁���.��9�w}~�����x۬~�/.��TV^8�w��'m�V6}�ףZ��6��f�ߴ���7A����0E��N��S���:�yӦ���_cm�n�m���o���>�WG��� �|�<S�=�z��wk��AYP�*e{ĚŵrS�w�+4�D�͐��}_#5��/����]\Y@�·%v����u�*�glN��l��^�.e��yui@jm�}y��t n�m���pV�'�q���V�n�<�I�`w����(6��׏��J�ǡ���b�J��p=Aջu���5��`���hQ V�]�z���_;�ۿ�k}�x'����M=�<O���:>Ɋ:�͵�t"���W�՞��`����{|]�w�*�7��~{:lI%�W�B���������n�sיW�{���>�z��s��3��+�+���n�i���+k3���oӨoW�����˿v�9X��V����J2f�o���K�zׇ��i��ͻ���1�(�u�����w{�R��l����7C��o���W����QL�	�Z����>���s�xuU�GJdn�]�fL��>8���M�oqk����9�Z�r�o�X�G[	{�V�	t�k1Zs,�9�=k��XǱ�q�%�¸�14����uN���Zn �6��΋ʚ!Ȗ��0%a��$1r�͈��#u��c����\�I�c-;m���M�f�	�*e�#�� 5�Z3XU������v�C�Ǒ�i�D9��k���L�A��c�ʕ����hc%n�K	�����"[��bb��h�>u�����B��L��ٚA�r�4sí��*=��%eR	|n�V�<�w�n�w���{��"��2'�׎X���W�˻l��V�@��.�R�Z�������[�GM�w��rwoW����-e��i'�ɋ�(�ۄ��*1oQ����^�����}�t~��{Ý ��i����۷c��n�% ��vy{����3a�1{��ޝ��.�{؀�A�6����aU/ˍ��?,�s2�t�~p�n������U��oůxe[�|���Y㚁�OQ�ȝ�=Oa�����J�ij�@8�;M�UwT�����@wSm|ھ���ד�)ם<��mz���:�<�����}�m�6�Ve�.��kȝ����]��$&������W�K���R�*�y��0p������QB�7A׫��aB���q��}}�ʲ���Cn���W�t��9�?y��N�6b���۫"b�d�A���A�n���`��U�1��oO��$��z���ϛ��C�L���C^� /���7J�y9�����;6Y�1}�
Z�I����{]����������[2o���M��ʽ��_�3�y�75x���������������G��+��䦰�m6N���z�n�N���;H���͍�qo��~����?��������<ƟJ�n\1[,������y��c�[C��|޷��W�y���k�
D>n}�6��:��^hf3�7�5@�ߘ������u��n|zdf���]R��\�Y^9���*����ګ�ܮНȝb:��]Sz�X4�{�q�����Kdb�ۦ�lK��S��y�ל�����8&�/�m��7A����y�I��_��_6�γ5�w��z��T��z��~��&��Sm7_7_=cڽU�2�����Ϋ+o�;�R�/Wޔtm����Nm
�uF�ȩJ��E�����k�l��CY�4�Oa9-]�Щ{\uӛ��3����VW=�	���z���Z2c�{�	<-ɛ�7M�͵���<"��3�y໡�{˄�3"����u���aƯ��oo�T�{��鶃k������1gn�fA�y�����_zW���>n���w�]�)��|�a�@߸yV��7�<>�_P��r�[���q��*\k���+��p8No�5PeJ��=�����OO|v�o0+�<����Ҋ���z���l��
a��b�B�DQ0%�5a����^@́����N�~����/�T�>o�q�_S�z�͵�u�y7����d�T<�۠��u{h�`���q�+h��W>�^Ӵ$d�.��_IC[_ ڰ����x}��:��9�̏eK>�W�(6�q�:�̋XҦ�o���Ťo�ݪ+vj�Ө6�у�z��g�ͧ���k��|��db���2�w�̯g����G���/�w�m|�}�tn�m��.�a����3#��{M�~:Ӵ�`�|=�}�~\�צ��7@7M��Z��]���Ez+�u������ڣuj�@�7M�zG�5���˯uU�u���f!��>�eg;���e�/�l�����e:���6e���]8��̻�I�e_D�ռ�����ҧ�b��/�㫫�����r.����g��ܶFއ�����G�.�Z֬����nXy:}���1�h$}��ݺ1����9� �읃�<GV�ͯZ���T�����'���q�Yy�
*�(r�c3B���euΦ�(�3���c��6��+n�5�!Y.�b.�h� /]d�`��}aX�]��Jj����~����KN���ڷu�˺�ٺ̇ys`�[���h�־_S��D<�7_6���J���ם��ŵ�uUg������n�؍����X.]>��>��Q������U��)����C�_G_��{{	�U��Y�{��o=ه/2_���t�@6ݎ��D���_m��}���a+ȃ�^��v�Y����u�~��{{=�y���OZ�7A��Q���Noff�/@�w[��:�t��b��{��7_|��~^�V=��w����w�.��r!gYagB�Ivj���#��& ��v��B�U�Tos�s�� �|���;PV��˵����o�cME�j�4�P�>�a���<^�z_�Y��=�W*�d<�l�Ths�~���.��J�O�M��Ѣ�l�;��׹�)�!1zǕ�����ҥ�S˧w���M���ٛ�T}�z�z��O6�M�Gf�^*��_7_6����`�Vm��T4�T��?�W���l/ ��9�tm7^�(ǵ}�RhEs_{��z��7��=�×�/�wmvYY{w2�m�s_8���A�m�{��{U�ʻ���৹�+ޘ�wd�/�?P���ؓ�]v�ywR(aϖ�&pb�דt�:�DVۤ���!�[�%�RxuՀmZ�OM�{+�=A����k��V�O=�uH0BÚ��Y�݀��3$f@�Vʅ�o��i�ޭ���>hO{^_a[�����-���഻ҹ�<��n�m���Ez��G��af/-^=ڭHg
�FT���:m�d]��Nץ�bpWQ��/��!/����V���ٕ�]��K٩���jﰛ����,T���]v�.���xrMۺ�����wB���,�	����wQ����V�v��w�����6)���{8��(8��
�32U��G�X4'faf���vFfT"}{7u{U�bT�,��qV`�وY �l+���n�W|�+]xk+o��\uu{��^Z��}�qh\b���:�LI�gE��B��]^�i[z��K�5�˭W�U��wB2���|�OwK��v��̼��|��N�u���S��䝥���/�U3�����%�K����(�Չ�O�e��sy��IgV�|z��7��wԝ��h�_^����붪��d[��ܽ|u��{v���֨�;�E�;2�n�n,���5�t��*Z�zEC�.XGgmu��q#Y�*m�E�[zo�^��R�:����3��pE��uR�3-u&Ͷ;� ��
���Y��j��Y�-R|�w�G.hR'x��{Y@�w(�T��UY����ftZ��5�ؗE��۳���^])���m���`�i�e��ʻ�e��߰int�#�|d�Y)d��X�,��W�h�Yd٥�֛ٝ���T1֨U��#��fda-�Zp��:��f�i�ˁ��w��&�C�G\���kj�ïM�aᓰv�x��Ħ�ysoq��VM�Y��e^k��v�knK�}���)�FP�l��6�Y����y��
�q�\���x�J��!��f:g��׌.Ƀ��ׄ��E2$I�� ��#"DЉ�&,��e&��0��12((h�$cB�bFdB�A�$ �(2b@dJLAAP4�̑�FQ0X��(E���)�!#	"d �3P1BF�QD�F��A1�!��d(3 �$l�HDa��L)$�H�	�X�� � �L�4�&F��(�(��F!���ɖ2l�"�%	�RFah�4�4�I�i���A��!�*B1�D����D4h�H�$ȥ&hAL�D%�b�QTF
ł�~�w}¹��ם�*���m��h��������y�&t�=X����N�+�=����k~zǖ���n�n�m|����<\+N�C��s�˧���S�k�u�6�u������}��;V��+
��h�e�\ź���c�z�^��F�Jm\�,�1����7�}~{���f�S/�=�S���ٞo�GH����ѱ_u*�mذ��J�]|�I�����.*a����7q��.'���L晎 �ד_�>J/��k).~��"����j���@�A�B�Q$��s}*;a�a�'�2��/'��1ٕ\-WP%�H ��� ��W�)J$����;#�H�t��
��Jink���/^S~P�z:A�	u�����T�.5u15�M+j��ƲD�N�|�r�"� y�}}���f�劽G�Q�֫|�R��y�əq{�d�\�1q�:گ
WÀ7�$�IW��(�)H��Ig�G:���Q��S{�"i�ƹ03�պf��q���}�B2R?I~��xL5���+�Teݚ%�O9�!�N�
�n��t�j\HV�`3e��b�@I��:�H!�Т�O���}|魼�ޓ.e�U�8Y���V�ݮ�Î �r$mP��R$�IIM�ǆ����_�q��������NN���7�����K�#�J�J�,�J����O�{�����A	@�BJ��R:0<���슺�ռUg�fb��n�q���=nh���/��E`�~��~�8������.e|�,R�;�u?/u�0�&e�Y=�wbH+7ʵ�ޤ3+�|Gj����H)D�A))�A	H�R��{�^�ȸKt3��}���+��r��7������A�
)D�AJE�S���Ğ�R�Z*��&��Ω��H6�rh֜�K��=Π�u
����~��'j�u�
�s2�@Sڋ�]�q%F�47�J&�aմ�ʠ��F���ܥ*��V���{#v q鎻-��e�4ڀi�b0I����i���㥇��.e�7��:�`x�l<������-fV��[V4f��7��^�ȝ\�"u���ښ�k�5q���7m�l�d���n|��:f�
Kr��J�(� s����M�A׋�#U�<��v�W%\FT�\ӿ{�I~��^zy�O��r&��3��kI�]�턍���v�
\�>ؒ�IP��R�i�Lg{V7B��p#F?e�^�W\�~Ϳ���e�v����M�,Aݢ�&vG�<}3M�<��9uK��/��9r^�����I�H$��QYc�Ͼߧ�_����������H��V���}�WeԠ���j�{�N����_@�ؕ
)D�AJ@IX���y�W�g�eł7`O�f��P$;�<4Lew$�q�p �{�o�\�`�Q�X�ΐ ��+"E��J%�%.p!:�O�R+9�S��/��
���wb~#;�X&��ݳ�{�{�0k⪥d�u��5�E�#�"pn�vI�&�[5a	��2�4þ���0A;�hF�R�RSYl{����/{)ߛ<#�#2���� H���j�Cv�M��ݫ��;�e���?�m���.&���\�������ӕtr�9�ċAe[����+�d�
�O���+��OU��G#V�|~}"^i��w$�~9_�＾�$A d��E����,x,�S��� � JJ�J>����]�G\}��9Y[�A��r_S�
�Ă�A$��Ȃ2R(:7�+�{b��5u\�A�?��JJhe��׷\�짞l��t�_@�Eɘ�<Ȑ�js�ꀃ�D�����H�I3�IK�_V܉��v�3���Q�>������.;�b#��|񝧏ﯿy�ѣ�b��v$���f<k�|	���"�g�_�='Pq:꒥F�~d�������"����Z�7���)����8K2/�骘d܂y������+�2Edd韬�>Y�S�?{��>��vz�L�{s�p���� ��P�R��[7�(z6g���v	����X���K��d�-=�����)~�3��ț�^W\qU������fJGt���Ʊ�kSy��Nn%�j����-U�4��*�OwM0R{�*u_���=�`�$A% A2E`����>���c}03�A4�QJ$JGrQ��aC�k=Je��=�}�;J12��"<�}}�VL�YH�2V[u=�j}�'ދ���g��*�7<"`w��	#�fJ�}"-�s�DV�������Ue#�%��sfb�静-���
K�b��t̸�0�!G���;q �ȒU_%{�zkA����N'��䊇�HCunx�d	���M�~�AJ��w�s��3��4�$�"w�D���5~�R�%<(ؐA�"HI��7���g�H6�~ �{�h@JD���Ģ�omnrRx���eZ��D�H ��?RT(�~"JI�X��U���ړ+��";���P:�wn�@ǲ��gO����f�ot�b�I����˺���B3+�dJ��(b��}��iwc%�r���g�f�(u�y�A��������iӛ�ox��֮^��f�a�K5�ٙ��)Ar/��2P@�"�~��z"���+�"y��Qꚺ4��Y=�^Đ�D����~w!~�>ZW�U;V.�!k]Zۓ��/3���l�B�9�,: ;X��+4\%�ݗ?�y����(�	IM/�3g�?)�)nxL􉎷x)Jڀ�֤P:�@ Ȁ�!��H��C����c`D^�}OdH�ï�K/={��>�]���D��v?�TOI�v�>S��t	�	!%?%XJD�u���;�J�3�v��Uќ��d��j���������v�ǽǅlU��:f�� �H��O����g�}���>� ��= �_@�=O�n��1�^�w"A`I	*��J$���$�����g1���$>�O������t3n8������(��%H�~��,�^Ѡ��g�@�e�ע21����.@��䷗˷t���۰f��^Aw���2��u=����v�ʇ�v�)��U��s[&̭o�z���ׁޗ�t\��a)�����T��nAsnP�Ź�a@���f�؍��M�!(MXJite]�#��3���M�nƁx���Hk��m�aEmqßIԼ����6�0�Z���W�[n�1(p{��pn���;.˸�����-�5�M�b�c�u�;2��Ix_N�{BC׳mp���f���M��fo�3!t(Cin��)���ۢ>;����������m��h���W��s����;^�v-s��������}�DN��dwj��H}������z�g%hY<c�Խ��>Ȳ)��|R�%(�%%4DW}��w��>�M��q$_l����n{c�{Ԇ'&`p;�'�J��{.��c�)sp,�{T<�A�O�$��!)�uC�\::��̬��D��c��q��%���%"AJ$JJh��"�p������F��~ ��
��D�A)ۑ����=�=*�#��I\��A������
�u�T�(�A ���!)�(���;�9�M�2=�>��w�����A'&zA��~iP��J �"ݫ��9G[b��=k�D�!���J������`c`��s�7i���ѕ�.������'"A	*�W�%!�=�[DD]�W�nD|o��`_B�����[����%"A)@+A�A~������۵�u�v���̷�����C�eޙp�yU>��g�7��2�{.��9thѪ�y�2\��{�f��ʌ��G~nGpΗ{�_����:W_n��A�I	.�?lY�z'~9ǽ��?%"JQ'䔫�y�W&�v�^P�}.��~���wwj�wl�7w0��_T����c�d�#�U|��{��DM��W�nDq�������r�ə��|<���+"D���BIb���\�6��9.H�j}��|��E�)OU#��O��1ȟ�IP���{���Y���{�|'����l�6���S��d�):�ܗ�&�.�0,�B���]߾xw��߾���Q'��׎��;�	/d�<&zB�:?�匪Ah/��H[A|ChH'2$�{V��fN�1�{\�C�����n"�&�Vt�r;�A>� �"JQȄE���y���lK�( AK�J>��k3{�uQb�@;�C~�3s:Y�A�fa�ͽ-�:���7��3T�>�#u��XC��^�a���f�õl�uVl[������"I_�D��	�;rjc�)�����6�^�oTRYr�h����,O4s��Ǹ���4r��v˂*�~)G�@�	(;��U��=S���r'��n=ۊ�	���,������CTX��n��{�����j5ʽ�(�Ŏkk�%��ll[�,�ށ��k�BXB�B�[+���g�� �R�$�:(��)H��rquF����7*xZ�$o�1�V�Dq�I:��R'�H �RS�zh𝞙3xc�:>��gO������oV���DW	���Fj�@����n��-��{UP'�$BR'�T+�o���U�Jj���{�'1�r�q�� ��k�ϐFJG�"�MC}��j���*~ܺJ$��N��]Q�z}��	{��>(&����"=�}��E$�{W��j�b�����t���cf����]d�'*��$����ާH�B�%(�����t+��D�R��J~���(��LGO���lh>jo�ͼ��rו?h��?>� �5*�J>��Y��1���ϳ����%!v�n�VLI�q��On����(u
�5��Cv�.��}������6W�$���IH�3�˻}�z��3\n8�;bONov����H;�?JJh��O�@�E����g�f��(q ����'�t�WsFf�^���$��R$�����W ���g��.�@��A3�Y�@�HA�$�_~��c
��G��K���e�o��>����T+�I)IU��G��C��y���9�'�1mW�)�<���^�7���>�q��_M�(mmo�9�S/B����y9�Md��"H��*,��U�u��
�mȗ�rR�;B�y����j����$~�$��������'��"�Y��0�^��83}FkZ`A�O��H�4�uV(z�U���u� Z��Sv�b�����`�ㇰS�QNP�֩멩����J��fU�Q�N��룬�&N^��=K���Tْ��c���mm=����e����PU[�f�	����wK���3��ǻ杮����
����ޏ�Y�:=�C�S]`γ�;w��vT�bo�<�;"ީ/����Zp�2+�?f`�*k֊�۽���ϋ��`�����>�6)(v]v����֚
�̄hV�q�]Y/�݋i;Emسwψ�՝�+{�鱮���Kk$��e�2&/Q�gwvm�-#nv��~J*6���ՕTv�~�2�ԧd�1�&f���sn�/H��.������ףz�is�Ļ̨LU�6�N�rq���:m��6�Y�%���r�iv���&[��j��9��
�8�m;�4L�T���Nȇ"��<G�dT��������$+��2�����k��k�3Fm�Տ��ge-9[��N��)fiO���<j�֔��P�K(3��`eY����!ӡA��RSWir�O��\�g)%K�.�|;o&�W�N���[E�z��7�.�
�K-�{�l:�����fiw��k�R�&]��w&C�yU.ggugv��s4t��rJ�7ՍѼ����
��G���5�0B]�����^�����-�mՑ>��NM]�3�/�Yp��5�n�{��ນ�gws5[�2^v���b��]��+�}��n�EDX��Ȩ"�"��X0e%$1�eI���R �Š�$Id��Q�R1��1((4Q&���h�Q�1D�E�H��"�6!&�Ec���Ĕ��)���D��,h�!2,DjLdƓFKLԘ""�4lE3`�
4j�,Q��Q�f�A���`�cBX1��[���bD*4X�	�ED�A� PlRh�h��`�m�6L`�H�
1DikA��Ib�
ML�B%3T`�hb�F�TF�1E�-,(�4`�FKb��d��i"KEE�h����}����֎X��kli��l.nE� '�λOL�������1�nl`�hT�m���#�Sc�r�\e�E6��;l^r���7=9��S�[����N��nn'n5�\�ulpPtF�h�(I�l�Ԩ5Y���z)^mC�U
��Fe��YDa)z������*�m��\�۬W�)�b��m\��l��n�G8a���u��=�NWPb�̯�V�n�Ů嫇�5)�mF�v��*���s�M�)lb͎-���J����Ğy.�5\u�a*��B�9�*��.Ǚ�vi
�h�n���v������,����`�mY�3����i$vP��#m6A�4V��5f�cd0b#
�&�m^�n���7N���8޸�n�2nT�\z2��Cat�1i�\�e�-��-�!��h�P�4v�����LX�Rkb.��M�s�B�,�v'Y�3���uv����jބV͗����{u���uٱ�Ok��N�A���G�aq4�/;Z��Zp�!�9ꛮ1>9磇��Y�9��E�x��"���ǃ\���<64�����.Nz�%n��m�;�T
���\d�Ջ[��-˹z���zp�q ���6�P�Ɏ�	asLa�#��apS�-�Am��;oQ��ñ�=':�%*�i�l]��%���Y�c�����M�(Ml���t!v]7���n�eWEԩ\����cw�&
��la�w!�wT�G7g�ڦ���WFb�񛜑�,SXPeq�m>&�}�q��������fZ �48�&Z���!�g�Y3��y륛�6;4�u���ǜk�zDթ�9��)�J��P�8SGB�"�k�Ա1���q+�4A2F�4�ԛB%Ih=ԇ�+V�=��؇�9�x�g�*y�<�ju�ol��$@��Q&��Q���!��`<p��7j�ˡ�ȕ�NXus��݌<۠�DKf��sF��M
L8�uYFXL�`7	)�F����[��a�Rm�n89�2�Ɲk^��Ƨ�qCֲn�s��e��pYp�9 �K�Ku&�.1(�72`�L�oK.DZ��:3f���5����� ��E8��P��.��Ç�=�pl�����P���4[�6gv�pg�^92�K���/j�������F���I�\�P��}'�:�e1���z��vV���F�Ͽ����6���X��uI���L��9��I�=6��-�^cfba�}��?Py����M��������������y�p�� �ڈ���B��fu/�2 ��X����	Y��>��\���9�~#S���3�H��e�H��w���A����X�IJ2�o�0z|=^�_B���t���	)
Q􀔏z�d�����9+:��Q�SW���}��h��Zn�L�����J6��u��ρ�$�ĐJJhZ�p���⇭'��} ���g�[eAge��W��D"Iw���H�I&T_n�S=��h��"�|�������p�_\G�^�|A�IJ>���UYΫ��|s��������Sg6���w#n�����V���)���Ŗ��cx8Z�[��^�X���}�+�H�Oݣ�Vm������j���Kz����#}A	l�IO�G�%4C���1�1��s��Ͻ���W^��j����h����vw<+kM2����U�Xz�fq9Y|KE���q��e��*W�VD�^�����5����h�=i��p����H#qP��Z��D8�w��È}��|�$����_%;�L���u~�[�}7�N/�#�?~�VA��J���YP�.���L}B�#=��ز�/��,~=Tco��������I��㏧e��K(W����x�$VA�d�N��5���X���5|����F�C֛��_	����#qP��ڴf�g�y����yӥ���-�@jM]c��퍘4���Ûs��mZўq{�k���@�]ď�+dH!b�����3WI�ٯМ^�G"}���G�6�<� ����	IM���U��{ס��{*����Đ��o:��z�;΃t4l��=��8� �!��3�yeϗ�X/bH ��@���)D�JJo]>��e��k����zH����Lջ��YO%�Z����Xu���B:EU��7�^p0�eV�j����xN��]�������}���Ƕ�AԨP)D�A	H�T(9%[�Z�y��!�E�_
���HW����/y�S�u�q���!
����^7|��$�{\��	 ��QJ)��aA�E�ݑ;����z|#lg��׻���O��I	)��R=w���0Ϡ�Ph�1DT�t��0���La�]�:�9�єM����~m ���~͑ �A%4����vp�	�q|.�	��[����E�/��� �%��K�3򧟕u�ZW�J����fȟgzWtl��{�Ҝ{�� ~�٠ c�%(���6=�mM|E��p$F%B�Q �����F%���Q�[:�1��ƣt8,�}@����"H��"+��
��.pܚ���~j=��%5��W���°'i����Z��g�o��,��h�sZY4��l1^.�e}�=�ѕvFՍ���K��Z�,�w�P�N��r�2�5��c��j�uUv){��y�W�P�#�Q ����﹚p��o���Oڻ����}��)Ǻ�>f�c�'H?$��Z��e�K��Q'LI>����5�cW�]q�ɷ�c1k6����1�5�>��{ I������b;��%�F�h��5�OE{�Td4�A�����IH�R�?$���n�|�)���,Ӊ ��4;w[�t9p��3|.�A/�O�J��-��:b8sS"A��}�)H	)�(���&��E���*ro��>1�O�:�G|A����X�/����d�ȑ ��mG8��?k�D5s����H��^0w��gz���$l���4��W\0����>��� �d��P@�KF�Dh�F~M��R�V�%C���7���_@�P�
Q$%�}�4f|%�fʹ�t��\ѾD�ܫD��=���r��F���W���,9x"��5�o��ԏ�'��Ot��ߑ�d&��۠�q�>F�M�|��F��7.��	<RnîSGwK�XA��c����0Wj�T3��xRjc�uy�Ep���k*<���9�k� Z,\��sn9z�YN�.P5-ђ��aԕї����z�8Uݴ@�L[������iFz�\�F�k�)�]k�ͫ���Mk��&v22����d^ېB�qt�f�*Mg�s��ߪ�\`16�l�q��u��� �m�,M�Z�m	a�h_�������}�$�$�������ܽ���^1�+�?WG}�-y��N���}/�5G�Ǿ �RS@��H �A��j�����S��8��r'�co{�g{�
�~���IT����u�:Ϸ��̉=���辷_+��K��[}���?M���e�KL�
�	}A4��� �������O���
�^�G�jD�-��A)��ܦ���J��8�8|A�f�"��B&�������Q ��m�� ��I�
(�}�(��Oo��!p4�-3Gh�zaP�o�@�����K���� �{(�;�����R�z.7Dnl�c�/����6::/ ���t��o�i�~sD=�%(�A���v��~r5p˵/�
���
��+3{'��Av�
/�A�H!%B�)D�"�vs����?~�tVĠR����-��E�v��e�������&V�wm�c�Uh�l��=�Y1i�����wjn�f@�bJ���[��r��媼?�뿈�"G^�J`�`�
���:�>�����R$���<muA��y=��҈� H?�AIP�R� �!�Óǌ`>��`�*���hy}�wbH#6D�������+���?_�䙪���R �$V;�s}�Foe��q�p8�����s"�pW�_N�竃 �đ�@!%_P �HD�/��Z��f��4?O��!�r�zL�
н�K�TG5�4AjD�d���-��v7��q/�j�	x�f�]��3����"˵.��n��\6p�lzK�[�#�p �ݡ@�)H��f��F'����_P��X�k�<�Ѥn@���O�(�	IM:V͇S��;�F|_D�Jnhv���<��/�"��|���|�d8]�+����%"A�@P?�)H��IP���Hk^�G����m<����g8]��v�VÇWm�#�0�S�>�ãF�Ñ'�]����oeB��ssh�.�Y}Ӝz�B�U58ɕ8^���G�wM@�"JQ$
Jh��ACt��Z��7�@@�w�(�>�����h�f�xK�
F����Ă#���u��u1_r$�H%%4BP$�6�	lX�s�$��v�����ؼF�C�= ��AcT(�H�"�\���j�~&��)Q�q�,<���i�{��g)b�
XB���r^:������Ă
�%u��);ۦ"\��YU��DG֍^�+�QP���"A���RSD%3�P'�w�yw��(���t�xTf�}S�N�P85�N�H �ȟ�In�:������� �D�	��_R�%(�@))���5T:8���YZ��)*/����AԊ��AJD�BJ�(�Z�sn�ڤH^�
���Oۏ^S.r:++<�tDw���;�� �pw�u7|�̆��"`p���AJ�s�Σ�j��w6{����.�:���uӉ�N]�u��i�8��c5pFD���J��mD��b�!)�J�$�X��Oެ�V:Z�:7��z�����pk�(�?r$�����R����[ջnL�Љ"Q�&����`�s�;y�
M���ޒ����
vB��}��� z��:D��A���^����"2褨��=ٯ�,�mT�}B�}%�]����E�.��u�8ܱ=���]1R����.'��� ��?��^~��p5�h�p$���
(�A	H�{���|�<wf>�ipP8c�P'TH ��	)�ґ%(���^��q����*����\I��׽\�;�"��%E��t�w`H"����F���n���A$�X2R Ȃ"I��F�����/�[���v���yZ<�Q��Wæ#�?vt�-�%(��%%>�렺��ȯ`����Cn�t�T1�\��g�qv��5�fn����,�^*�i�T#��y���+W�زp��Tw����,��Uv.��#�٣ݘ�C\f9�"�ʸIz��ST� O��=�D�݌eлZ��ͷk�1$�q��^�蓱�$����la��.) ��nI�U����QV�Z�EV]����CR�ݓH3hs��]�	���۳��q9�]YH��3?ȕ�9z�3���4tx��v\�����Pݣ�ٓ����d�&�������Y��qwWgTƋC�çq��\a"h�͠ǘq�-�j\������`	�
(��?%"{NzcV��p���H��A�OtN&=�����rN���S�Q�A))��f�3o���p�M��{��{�D�BJ��菛��ҡ@�8��۵)�w��78L��"�� A �K���n-���K8���K�b������]4B��J'�	IM��=�!̆s�f��`/�#;��Qd�����3tOY��㐏w¾��Q�$A���X"���}�"JQ'��_%"JQ���܎CA�l����W}�pfr�/���Av iH�R��R�~�nm'�f8?�Z��.5wV�[j�+[+,HV�VPD�I$*�Bn�`��� �P�wЍ�ս�9�F�ۜO���?��cVw>�s̼��X��[7v�&�#�E��{d����dE�詨��VD��1����L�9�z�V�Ġ�+����\����Q��}�6�̙���V�w�kU����j$;�n���J6�� ߄Gr'�
R'��sѓ�#�ю㐏w#����?fȒYܶ.}胼w��H��ğ���IH�R����s��U��zżm+�L��x��G	�~ ��W�E�BH D�ō��Ó/�t㔝z�/��B~"�U|~JD�c�O���/�B|f;����lxv{����TI���W?%H)*�(|=ˢ�t{���q����'p�|}��~!%U�	H����z������m\�M�`���mE1ӸZz�O]%pܘڛ�y��,�ן],�"~)D�@))�����3����X���:�s�ެ�˯e�ψ!俟V�dA��@����1[}o�E�����T�����@��;)J|f8����vD�R���-FpsA�?���dH � ��R��d�?H��m��+�Y�<U��1��ܨeW\��`-^WIk*!���Vw7��G1*��5R2�n��o+4�j�U��;2 �jRc�J���͊�ZEs��*\��P<L������{a9r��x�1����0����Y�TҲS��ڃ���d��޻v]m�x������0[�z��ҳ7*����-j}&+9�b�Μ˼�yZ(���%P�-Dn��֮��L��gWj��6��(�uf�St]4V�&�X��w6�f������^n�C�)�d��GOh����6�K7ul�o2�%��5<�>�:��B�D�f�,�6�����M��We�Lт��kĪ�Z����4B��ڍwFR�ݘ������@����<T��ʼ����U�܎��K����l�͛�;�B�C��0s��Gy�����A>�Y9{7�b�B�2#�������ATAVgUEx��¹w*c�=:�]�1e:ב֭]�n�������5r�+��n��v%���I}I�7�ݙ��*άܭ��x�;ھoEɽ�;�۝|���vt賏oc�D꺚S��x�P����7�<T�yu��"��%��Xʍ�!˙����}2��eW)��;tRyb���]�m���f�zj'%b�6�ʶj�b8��HgV��&ud�Wf�Dpٔ]�=o;h���
�Lt��+���\9��
p��'��9P����Ƨ\�;k�|9��N$.���k)T�t݇"n[�*�m��]S��M�g(�%��G�9l�����/�U�W+��_�$X�`��QF"�Ic	lmE�M�E����X�`�F�clZ�TV6(��5I��Ѵ��h�-2�F*5AFѢ��JѢ�EF�Q��d�4T%i+-%��*ěQh�Z�X�1�h���X�5�b��U���5�TL�Q��5!cQ��lm��cb�c�-Z4�h���5F�F�-�V5�F�h��I�lEF�Z4�HV�Ab���AR�a�)����=�r��.s�����~��|�I.�2 ����~��-t�_��΂���A �����.�����MG	��~/`O���ml�i�})~���%��J@�(	&h[n�nR�߮�!�چ��)1�P��Q������dH)D�A))��$������ךվB���֛02�k֣UIE���A��Kb���E�˯�s�b<��N��b�})H��߲�{����Jx+�y{�7��G�t�ۿ���S�Q� ����� Ý�Ϧ��V���or��ϡ*��p����	���5B�Qaui���#+,�7�̛ʸ#7l�7ݹ��n��O�˩��Y���p�7)UF�E$����t�v~J=��%4JdUgy��X�Dj�yЯ�(�(���]�&<{Db���9��G��R�ϪL�U������4~J=Ө^E��5��S�Wuek��~�6�=�%��fF^U�+mS�An�>ZaݯP���jg�gu
��ԉ)D�JJh�����r��W)bz�uk���X���$^���QJ$���� �s�	OL�DGQw&��u�a8�k��;"!Ŗ�n��ev-��E���b����J���R&���8���"�|}��{�C���s�"�� �\��4 L�_k�yVg�r�����>|.6�{���ĥ<����bH?fȟ�IS��F)L��Ҿ����w��A)
Q��RSY���k�y[���753��5<':A�	�/�+~_$�a�y�VT칗�51^� �n���6��P��Y/���w�����&���I��
ϳcH'qM���I$�W�(��;Kg��/{G�O�ᐭ?h3@��	Gy�obH́ ��W�%"��W=\j*�J�{g�͉�l�n>�KC��19���������N��gnjǹz8_T�zI\؍R��8�Ы�6���nw\���{�����<�׿f6kcb�n\ٝ�u�N��K���X���cn��&5B&�f��66�ǝ�"�Z�U:w���R$��)�;�[+Շ�p�j�X��E�gn�0��T+l��u淬vl!l�i�-�v�A�`��\y�>�sU)�/Via�����Q!�T�f|�t���[�-����w���jj��웅����m��[\�3��[��!��Xd���+��퀨]����p�ݻ\8wWJ�Į�u;���e����Y���G���|��˹.S��5<':Ckٳ�x�nV���A���tX ���!)w���̼�v=<T^�~oW���0��s�+��[�|n8�����r$�YE^?>xw�̔Y2ŨA	*�(��)H��=�����������j����O9��`�}�=햛��n�c�S�������A�$�D�A))���um���ӑ����	��$tT<��J"���q̉ ��"A	)
Q$�H!%�y]��XO�;$jH��[,s��n�ӑ�����D��A�%)nm/{����?���)��m�	\4���H�2+6хhmz���lHWc@�!�����e���e��РR����/NF��u�랒�p��g^V.k=��������A��"�Q$���H�{��
��n�^��Ip�]qj�7�˾�Jɱ/۸�f�{]�
�m��n�o�[0o_�����
�r��Y��ćþ=q$��47WoV�j���6�8g�H?��A�R�_�[G�
B�Q�U��<����)%u�	H�b| ���S��"��k���5��#�?�4#6D�����;�j��DV\@D-S�ذAJD��sn�z�GMa�MO��@�w"A:�S�;���=��+6����V|A���%d����t~X���^���f������]>���ns�{�������A�)8{v���v�DX��Gsc�����[q�b�K��4\�4mĹj���vc����0H��\O�E�n�L��]���:�{����n��,�mNLW��7ϊ�V����,�y�l���ݲ����ܽ�_mł
��k6WW���g�������3`I	-�9����6�݁@���VD��J@�$\�~��r����������i'��(�6��ƌ.Y�r�c'�T��w��5�P�6\�9|�ոBã����Yf-����巼/hǳ����VC͍��$\[�U���Tz�������	�PD9b�2W�H�"Iv0m�oR�;;�����b�_�~�7R�j�=9�}4��<�s��}����W�^woݰ�#�E��ۛ���N�xB/$H����Ww	��mW��`��H~~A$�����C��� �ZL�Y�d8U���Ж����tRfn�)Z�����wN/|�u����{e��X�IN���[���G��b>ў����ٟ~o��{�����dy�\Fn�bn��|���3�'�h����~�1��eS~�珍�|~����H�R��b��f���V��P@��ŀb���Bq^G�c�%۵�n�_�ݢ+����s��	���$�/�"�H�a\wvr�}?oG����z�z�{y�^�Y���	݁ �kqDT�h���we���۽y������y��wK��e��"��'4rjy\lloN�B�;�^$�A�WFՕ�.��J�Ҷn��Q��m/�_�ϛS���&��ɻV"�XBH��TJ�����1�ޜ~~�M>7'��@��D�R����v%;S��K�|ާ����,hF���:]G�있�R���jn$:�F1v!l+�;��M�vo�{{�	�B��(��J����xg���U�+�����u��g������W�@��H?$��}�隹����2|��}� �k����w��*�+�Fx/t�w`H ���`�Y{o�yn(3ւgz��ޯ���S�% �����.��+��.��m�\p �}�4?b� ����/�l1��yP���uiH����7�r��ƫ�W�P'r$*��Uj�����y�����Dwv���[�Y;\��ߣrPe��X��w��/����8���?%���7����ih��ݳj��k��pE�iڏ:a'k�X��*�ו���]mޢ����C�#*D��m�Ϊ[#�.f��/M��w�|�Oc2Z2��r4��靮İYb$�]�h,Mj�d1��,KB��c^+�\�HX����	��@Ѕ��R7Q�Y�Z�F�����iVR%���㧁�<�A�Eǃ;uucKE��<��[KLM��DF�^VŊ�#+v���c�mN7=:���!��Xh�g<L�)p�ňa�պ�����Q�ԉ�8dH���h;WZ��`�&X�����o�n�f�e���㞽�G��:X�Y�e�6�]�7UT���^?빾��#�����D�M{�f'[��e�Mt�qէ|�gye��[7v�7n0wh����k����w�z{�Q�P����ᢻ�AMW�r'�A�$��+{fߣ�Q��
��Q��9�?%�J$JJ}n�Z;����2��Ąp^�� n)
Q����!%T*���{=eY�CSh�"H����!)/��+^�>��:O:r8���3y�~�:�,?�ȓ�.V>"D�J}$�fJ��/C ��'pB*D��=�]���"
j�%}@��A6D�T+┉�ZҾ۫���8��A.6�A����l�t��C��K�R���t:G�"&&EF޸��nh�3dIJ$�
Jk�|�����{�=õ���n�&�rok�#7l7w�`��<>�9���|��B�o�׶2|v�٧�q9��o+-}״[�/�d���YY�M�ڷ���S99t.�Q�K*Z�cR�&���w���7�3�?P�"�obgR�f���'�9A�M|A�?%^.Z�Z�}À5���\�{�		*R� ������e���M�d��w���%|(�$�HĪ�J��H�_NlMGA�1�W(���z<�)���1�����{��� �Gv�ա�q$��	*�JQ��"A���ud�.7�����#=آf��f}~r�͜�1O�G��)��آ׬���f&}B������q�����{V�z��ci�Ul/�[�GT΀'��� ���2�F����hK�#oܔQ����`�� ��W�D�JH�`���s=��e\H �q)�����X)�HO�N�#�X�d���N��a�@L�`��D$A$��C��d������f�q�%^�٣i[��s�X{a����悎1�[8m���o�;�[uY(gp֚ʳ|ňf�����(j���U�][��V{��y���ד�c����"���!�G��S�˔�h �$�g�%���)�/G9����?<��}@��;����}� ����H��@���R\������f���:7���S� ��g��Py�����'>���>m�2�D������LGm3kcg���L蚨vc�85�كvq����z��Y|�e�$��_�����^�qX=����+4��2\m\������2D�{b~ �"�H���9!k;�9|0�~ �E��
#B��cu�/H�>��"HIl�P�;�'Uv���$�@�l���(� �ׯ����STw3�ϧ�)[HW(��A�T(�AJD�T(o�v�ݘ�zj�/�$�P��JE��_V�sK�֓[���z�h�>��w�C�Q�o�YƲ�)�2]��B�sf���f�ܱ^��V��t�
����b��N�*�)l�e%F�z��돤�t�!)�AJ�~IP�R��P#/7�>��u�'賣Y%�gS~����l}����_�K�86�}���x�{r�n�G�jSvzJIC���e���/�UL������	�t� ��H��O��M߯��w�>½m!�]#klWXbt�:n�H ���n,R�V(�}��|}�s{鯩#��?j�#�.���}�Vz=i5޸�A>������~���w\K�=����D{�	p$�U�Qd���#�)g�i���95�+D��w|1_P%lH�IW��	H�R��$�Q�7sD���x��IM�}��=��1zճ��:�IrnLۣ�S�+�;�\M�swj�v�wt����S��1��@�;��6�VW����ƃ��v���S�k_}���  BI������Z����V�m�Uj����V�����km��Z����V�m�mV�m��U�[o�Uj����Z���j�Z�{�V�m�Uj���j�Z�}uV�m�uV�m���V��mU�[o]U�[o��խ��Uj���1AY&SYI-�Tn!_�rY��=�ݐ?���`ϟ �                       ( R���� @�@      �*�R0  �>CmJ
u��P��0�B /}�@�X0@�&�2+�|���0��:�ǐ� ʕ�A_F�5����GH��z=��4���({� �)� �  y
�G�4({z�:�tkTm��z���kx 66�%�����J���7MJkv`���tu�v;����p(  A[ʽ�.���Y;n�C<���l�dV�&ړ\um�jv�e@�}k�۶�0�t�@����h3Ն� 
���  }�M�A� k=H ��K= B���e���(�&�K��     jzhRT�0 `� a���Rh�   ��*�UUS�椀2� 4   3*�)*zH � ��a)�MRT�2h �� i���hT@&��mM�����Q�z�6i)<��W�T����ڞ�63�" ��C�L�
�g�C�DP@��*dO��b2 ����Z�����o���h��v��H��(
�`����*w"e$�%M�=_-���Ͻ`�������r���ϰ^�2,팆@�0���X��o��c��k�`0a!�W����gS5��aڵ�?�O+�����*P��ҏ�w�5
��ha�X��CLft��&v�M��6�)j�S��w!�]ew^�F��r�5B�l���ʧ��4-�1��Z(�K8�bۻZ\�+�0RA]�v	&��N�^KO> �6�uk�j�Hrۿj�8�j���æ�����Uyr�oI��K'���{wO��Z6�����N� ��m)ѹ��Jj΂r}�L��>o`KH�I��vpJ��+�x��Z��'V)��NBl8��#�d�2�Ջ��jL����opL[�^8��+۴����B=��>�{�
u�ȣw�{��q��rg�hZ28�t)�6����g7���dx ��N`�#��i���[³�M�0�?)Ê����vA�;v]�٬��i�q<w�HMB��rb�b\�$:���M�t�	1�o8^}8=�eL��u1ݯN��،ڨv��4�)�Ep)�W���s�l�V�tZ��C}[hZ�!6{z��u�Bڲ�A�0-jc�|e����j�����]B��ın;���ڌ�U3yreu�t$943fS�9k!�X=�w���ߎ0�5}�7[;��\.]��k��GЩ���m��Y����Q�E���3�VY��;qd��Jg*����i���ӹI̽�w5f�����&�m���;�E\x�+��)x�����L�*��[�c��KJ$��r���1�o�N[�
���
Vn��+ln�i�"�nhG�w���:ã6�9��(2���b��J�H9A��&w,�OsKCzu=E�v�4�,hO+���ܒ�<;���K��#">�J�4;�d��8�LkR������+gU��z���	��X9�*U��کN�[��1c���>h �I�-�+�l�0>;�ja9 �
j�bw�͜b�f��>��0B�@GD,՜�(ֲqE���W������v����GaZ�`���1��unɻ�R�8�ZY���n���u卙g�i\�����s�	س����G)�ȵ�s�˥3H��$z��0��J���W׺G�cc����od�b �h��L)4��E���ЗP�w6bX��wͮ5��i��p��Q!8���p�)�ܜ��7��;*��k�s���^�x���4[�����E��b����\�[�>��:[�]��۰n��v�'��r9�ɸ�k��xT�*y����uܡ��X�)wU��<
�cA�%���g!睭�	������0��b�\[{�.<w�>�sah���-B�l�k�+��f,�d,�oBAn �٣��I#��:�U o[��^��w톌j�{�����������u`F6ovu�k����p��v�lJN»l�>��T��{{p.���)�ˬn��S@r� 	GBs�6�"NE�'��v�`�Ocm|�!Y�3^?���h: ㏶�A�5�p5 �5�j�p�}ܰ�w;t0Ü;U�x�}=㴇���zd���ؑ�g]Z�lgNMs����q<��Fvl�@oF�9.�Q��Hn�ZZ�p�;��+S��U9�h��n�=U��Fճ���$�x��y�`�=W�����6uǔ+�{L*xw�fώX�+un���)y�c��Y���D��渽=�4ŗ{�饗n-��ȱ^�;P��3mO
�q}ϴ���cI�mU�ǳ]=y<�Z�_�ݗ�"�Ynpgc��҂v�
�DL�5�]
�ۮTN-��wu��'p�����ӽ�E�Qd�c+Q�:&�L�����-�sG5Ķyo.��Z�
5��+���� ��f�ҕ�jB휰՝������z��"�$��;�@oK������aL��P�ig=�͚8��\r@$U�a�n"`�Z�-k1��׍[���8;�vۧ��6�Հ䳔�6��A;F�Ȳ�}���'�F�oF�%�4ɓ��$��Bf�͙��5��EnsuEX&�
i�[��wz�P<$u�H<�j�Q�.'�^�jp����vs�]�tAaD-���J.L��>����9��&��d��A=7�,M�����Y�e�΂��F�1J2�d��:s�>��ƌ�s�f@����t^탙ם�C�8�E��Uf��6���(Q;8�y��.-��p\�f�(0�q��4"/���b3+7S̕�sI��R}�VP�[��oCt�8ۛ\VYe&���q�G^q�rk"��`�fA(���ۼ4e�4;wg
�:1V�1�M�uk3�d����t7{�̝�p��_v�� ��ގâC�޻q�Ϸ�.�4�����v#t��%՜5�s�����Dbe�m��cuem�[M�١LM<���80K�E7ZW�s't-�7��6!lI�����b,�V�˲�3�������hĳ`�vR�O`E勁{��3C�Y�.	� �o7Tj�.�3���ʒ�yoA0�Q��c!c��e'a���w��;�{׻���.K~G�8�Ͷ���ƽ7Wd֗t+wL���a}��?��?����>��<�vx˃t�r�����9���O^|�^u�2ttz�C��
%   �@ ҈� �-"҈��4)@(�ЈR (�B% � ҡH��(�R�@P	H�B��()H(P"()ЂM
�@+H�P����=G���û^�#o-�b?5 AR�#]3Ƣ**�;s�Q����114@T��i<�>���"c�P��{���N�˫�!x�ިДۃ�;^Yrr|��1-'�33��$δ!T�`ȡ�/��	M/;�>�<�S�P0`�1�2|i�T�]C�Eͫ�-[[��<8�(���a����	���[O��;{ۊ�ig3@�ʼ����§��r�f�i����Sxo�d�e1oտb&N��;�o�`���v�m�\X�LV/U�e�}�ͺ��bY���#ݹm������2`��;WP�|-�%^�l�<���xn*�ve��!�����zb��Oe�ye��<N_R#�n�C�{���[Gu�w��+�9ᷚ�P�f��wf��P������u�8�G��W\��z6���7������N�A}76����Re���T���kݏ�r��P��M}`Ǖ��YsW�)�"#�c���uE�k��_z|3��)��m+�r���'���2`8ø��8=�c�}哽�iA2�$v=sF���kP���7���;�{r�Hbn!�*
z��K�=���&��{���0�g�Y20yS�ڹ��D��y�w)�"�Xx,f�x~aH�`���ކ�C�������He��Kyx�컕\Wq�q�[�\5��\���:�X|��)e���]yT��`����{|.j�p��=��9�o���q��*���Ӟ�w_�r��ݒ�ȪY��8,��ݾ��{<);^��A�7��I�|!����Qjn�n�r�D�t{ˊ�^0�p𹫄�yc��|�xV�#ݿJ{����ݑ����q{p���ћ���=��p��1v�l>ۛd�&}��{��r������"��J:��ށ�uL���T��(pm�y�&g��f��6�N�+v�;��;5`���$���,*[�J���M��!���}�I���"H���X -�6f� h0���ny|=�ӻ�u��{{6 ^�פ�y��&�<w��ǽ1�r��d��V�:���~����J�V�� axoM�+�v����d�쒯&��I�c�t]M�a��� ��6:�c~����ƀ��~���,�a��nw8��z>�$�^��d<�.G<Em�����4\#�ض�a�TW.�Ƹ`Ò�>���z�;\�ۍ�e<�Z�1t�dp���R#�oË���r]���l�Q綯��xyd���p�
�;�,i�ৼ�A7~�=}��߇00-z	��G�.S픬�P�.�<��ۆȤ��\�{��S�	�_Kf��a,�X�X;��F�{���{Z�	Ϸz���t���^;6\D�ݱj�a`�@$�Ѻ�'�}�f���^ʽ���=:>�;�?Y�3't�-����Tۄ^J�l:G\���ͬ��o5�Jwݝ�鞚)}�Ϯ��F��<�G��Ox{�'�,�3�����쩑�9�}�}�����s��U�0�gghrd<j�Q�{���m��x����۩���V���9hgJ�P��]_����|��s��t0٣y���{�,�p���hj����'n4z�	/�D�{:��-��ˁ"���O7�V��#I��C��pA���o�oG�+�t�S�٭rŒ���*�אz{�=q��2�?L� 3^�I��n���4a;|��N�x����ߥ�<�#�gw��v�[�ϤՊ�:r�/a���W#1zI��
D�ʧ�og����*x��J�82�wnQ��Ǘ�@�+;��׵zM���}&ߘ�����qv}���3�O*��nH0�:rܟf��/��������C�8z2����V*������~~�1���vk�Z����9��,ڣGݳs�Ӫ��l?h"�q��}��._M��_�$ޙ�6�'�&��}�=,�X"����F:g�����[>&/��_.�9�ϰ�^{Zϔ^��6@G3��wr�K��Ͻͧw�-+�M
E�G�<^Z��n٘y��p��qS��F�ݠ�m��t�}ٸ��0i�2�:/����m��&q������Y�9C���wmݾ��-�[v=X7rb��� F�ޡu�^]�^:*��ӵ�~���^2��j�d��ު��\A=}r+���� ��1{@p|��ɘ,L��3�c��V,�Q�=M#�cd�~�~��^8.J!)�=ݭsܟ-<~�y8��y�{'�{�x�����,�3B����R���$��p���j����Gy}��Xo�fU�"�t$�~�pxv��W��ޗ=��r�*|��6L���/������N,Y��ߟ���@]�ܪІ��4�lfLE�yUaS�}���3@�]���-Ŏ��.���Fs +�5V"������~�3��O��v�vh�O2����7үL�V��}7�빏���0&u(:�6��b&��Ɏo��a5�`�0���ӐeG��%�9����.#҅Y��(�k�x�f'��ׄ��ΐs镟=*��A��X0�-ҟ������r_R.�*ф�ѣ��na�9�QRQ=e|v�������˘��G�<<2y����2�����gL���X��7��,ŕ��5>��s������ {�"���+D)X�P�s�'izB�0����*�rˆU������(�D&�.AGQ������:4��n���V�ĪB�h&"6�@cA��B,��l��Ź̺Gh�,��@���uT�ؑ��)qG��^Ҷ[��Ջ5ݬ��YH9
�%�h��m�`�g-�y�iNI�%���9n���>U	���n����Chv12��K�qj�T�.��5�ȴ^e5%�(�ک����h��̘z�Y�îՌĥ���m,n� b^��D�H������&ˮJYHa�֙���-s�*Z�e�]�����V��į��Գ-��
bh3ub[A�P�˝\��x�\�#�5�6.����#,Z���QJ��J�uѐRa�:¥α2���8��ea-�z�e ����Y��d��Wm�YiX�9���X�e���l����	N,& hYvA(݈�L�,�*��Y��6[Rl��YWK.�ks��V&��6%��{[��к��Ə^�j�:��̈́ݍ��<D.���շPM1s��s5ƹ�JL��t.��2���]b�Sn�$5��u
k$�%��||#��!|v3wke̬,�,G[�[e�����pB;km���Ku���knj]�Bc!�IK����k�lՄ)u�]������ԁ�]B��Je��1hhն��\[/�Ƒ%k�(<Dv)�eͬ�I���goke����N��\�)��D��*Y+P����`l�i+3X�h-��P��Z�F͔.0F嵲�Wfm7�X�e�.�(۵�]Gk���M��d��,�lY�6ٹ�m�a�Q�)���F���K[e㌸���e�d�%#ʜXJ,�lmf-��0�[�k��,�J�ja�.H��M��V8иƺK-�����M6�+l����"���<��#v��J�4�4lu��fcP[Y��i���ݦZ�B�W��bN��Gq�aYs�����Y�
m5mݔ�.�[B�M��ku;]�����,6"�,�Bń��n6L�-���Se5��]zm�P�K�3n�.]�Љ5��Q6mQ������ se���=��Ⱥ�c-�l�@ճ��#a�eR�0��0�bKLҚ=�n��Ѯ݉��Mc�l�]M�p%&��[��e�t�f���u1!<���g��hI�B�q��J����-��(�f��m7C�X�Yxp�in ���P�@��S&�k��kŬf�7�ЌQ��G�Mhp�	���::]i!Z^�,�M]E��
�%JQJ�I�,����0��X��w iE`]1ak���f�3\:8�mee�M���ڥ3ͯSf�Ys���v��R�᚝�KY��-32F�˙h��Ԇ��6�-�K�=K3hЀ4��0�d�n�&�[1�L�\�3�X7��ӊ(ƻ:�.�LR�l�ji��6��4�qh����7��̬l�5��!f�5��b�62d%������U��uI��z�єͺm�6ʃwK����e!Z�Z�m�m_2�v.���i�./2�$�7K�V�Qѹ��Z%���ly�eL�8-�.�[�I���]ڣ�����]�Z���Dց+���V�n+-G7m��n�6��1m�oY0Z�b�jrrb�`�����6\momT��e6����3i�����<�ʭwb�2̲�v�1^]1�bU�Tk�XA��{l�
][k��cۘ.��Ĩ�W���w!2kc��al�dH�6��m,m@\�*XmM���6X�c����yiY.k:vi�5W<;b5Yæ'6I�           I{v��     	Xl�   0`6�)˛      `�X猚�I�/L�Zy����V	aMv�*�ko<m��ȵuj�
�fJ
��˖\2����m�N��[��п���-�DAWr.$Q(�\Α��$()())JN��ӥUT>cH�`��H�%!��*����PĔ�е��F�[�.թ�* ��
�F��rJ�[KNI�P�6bh"U�(�3���v�����J�q��)M�\�7�0�&�AHm/J��caƿ~�q��6��.�u�1��m��c�mi.��k/X�j�ݬN5
��մ��a1�l�Ii�9�d�]��R ��9�jm4#Kq��ƪ�\�;Yc�2Z�k���㫭�!03DeY�j"�$��������]�[�s�����Ĉ](�nؚX�hə�֫���HKb�oR��\u��K�6��L8u�˅�����&F�����[�`��A���ⶶ����R�2�-��*R�����E�ц�[ -��҅`G�u����mmn�玣t��9�m�����R��̲��՘9����;�6�*[�%��i�L:dfuK�)h�8� 	nL  �` ���:�M���f����^s�)��`iu���.�h��u6����4��mLm�LC]�M�LB�!n5����� P�׿��%������%�Q����'�2�J};��o՗p��J*ɡ4�d��ޮd�����%%
���N���&E�6���)����?a�W.��H��6�ݘ�޽��}�'�mk?4�)k@��&KX�M�ۢ��;_�o�����.|�(��-�_MD��ꈀ�a4t�ȃ�0���i��Ǻ�<h@�%�Q9�o��p�I,�=B�V�U��/K]S�q��
�����m��j��?+��j��\�z�eLE��E��zo?A�/:I�o{��wf=n_(�!r(��J��=��d���;ezѝa��)N<Hy|3~����>p�5+M�B�Ҭ��x�E���V�)d�93��[�t�iv�ر��4>$�Y&�' �Y��*-�o��UҘ�/���Kf6)Vk�{�5�J�\U\E�EV=J絶�1Ɣy�k�tN��<�u�si�UW:�0�A�Q&�{
�b��+D"C��B(��MP�ګ{�<,�J��e��3
 ���Ie�A�e��m�o�F:�#42�F5I3!R�y���2�n*��E#�_PQW�y�xY��J[���AJ���n���ӣ�(���Zۗ����9��L9���J&禵Ee�Z�i�Urjmf���Q�u�`fL�(�{B��L�CjK���M��]�VYP���b�\ї2�C[��&ᔰr5��N��aM�Ϋ�v�� \#���7ߺ����q]��%%�H�][�s�dR��!f�ef@��r��:ٌ��`�IK���qW�ϗ,�B!wE�ܐ��^<s޺�Vt#�a!!ǥ�����O�Q�չ�=�z%#��V�T�%����������ͩ����U�z�p�&�k:�Uq��x{O��T+�OwJ��ΗfQ�S�	$�'N�s��}P�U;GN����}��~Ӣy��)$�׍�mۿ���b��`��T�m�^IJJdI�*
��bft�j#�S����q�q� ��I`�>�1QZ�s5���[9��Dz�(��#AKr�c��	q�����ܐ��z�s�2�=����������̀�u>y���ե���)A>G�gf��O��r�T�L��Q*e`��O/Ech�J���;�{8]�Jj��Z���7o�h����	I�Ţ�:[�k	B0�2�^%�u}��\]>��
f:�M��NC�����l�{�
�"� ����z��ToE'�ř�K���uԅ��w�>��5�8��vLpJ"l�QT@�7�}��J�QQ�B)J+���+�y�(h�TWt	ȋ�Hj�񶳃�(J(���D��ݷ��T2�ϫ��������`~Ը����8�u�ӱ��ĝ�ݵ����l[3
�a&�-GK[��Rݓ]�l�@����n��on�!.9]k����s٦������%q������������k�l\�ͨͦFf2��H����9�0�%(+���o-�OZ��10���EfwwM�����yh�����L3w�y$�����sY��B���(��Q����^s�Yn�����a�����XΛ5��QZ�����A+8-0s���T��!�a��޵��.�뗲��f"����K�z���Vg\�����[߻��srO���~8�ww^�xd���:�\�L)��@�Q((FR�*f&�4�5���N�@�R��Di�A����y���e9ʜ�PqQIPǀg����
�=��R�N?(��Q{�W]>��	�"�{(P{c��˓׸5�H�|�sik����r�Ơ9���i>���x'm���M���
3`��ۛX#�v��ȕ�8�nx��a��}�z�Ӧ��̀�����!��z�)>������^V��L����B�þ�9n�av��x�!��Z�s�XO��o{R�/�������{�˴ѐ0�9n�^���9N�/���$�!�'��ȫq�ឨ����jPd��I&8�=m%������j���eN�PT�U�_����^+�I���l��OpfR��h-*PM?]�T�rh�S�0Fq���!3+C�\�
���h�l�'h\1AKC��Rx4��T�j	��*�J��R�KB"
�R�nD�lԀ(�U14�I��ADU��O�D��S����P����+V�g�|�����3~�$�+���o7���{H�^=������`�eB�mWX4�bQ��ۃ�<���y��]���}e(�&�ˬ�XZ�x��g�Fz�ً��P� P���{��锒2�Ӈᖅ�������y�� o5�vhj�]i���&*6��!`���N�����>}�U��̛�>����#S�F�����S&
�%�&e�J��X�H��*)�}�������6��3Ts��w�����Ϫ��Kf��x2>����}�#�����-Y�����v\�PE%�5�����}��2��]���1d�)E�������h�ڜ+����뽈�)�b�e�.q�BJ���V�Xb�.�ٶ8^гL����ƷXTY��\A���=|��Q&�9]M��r�m�b*���߿���Ś�J!J0D�(( bL����}���P����L%F�.�z�y}��-���.�]_W]��?��2B)��t�������=/��>����QQ�s���|���{�e#�|�2�0�"&"bI�!D�0�3
7M�N�n?����D�Q
�Je!o�N���J坧�PK�D��Ӈ�	�2a19��������Ϸ��cKWq��>��V�_s3�{� =�*�o��zD�R���� ]#g�{�s�K�<p]Г�(��Nd��nC�ꀜ�?[4!��[B��r��>|��&�[�sU��e��rTL����/��%�Y���59�����Q~̅Y�[3�V:�-̣1�~�<H���n/���M5�Kb���Oi�w&�IC��>����6�B��5SҔ0�����ʈH�P%L�3iFܷ��p�82���L�a^��Š&�;�bD��@��m�=w�] m @�"k��ˢ���@4�h�h4�F�1��HV%���|�Ͻ��}�i �4��d�$�8�=j<H��.`�@߽x�z�� ��������G�?Y�ڰ���{.#�1T��Ji��3B�������f@3#�"ibGHt�%$o��w�\���ր1��4V F���?\=���ω��#IrۢCQ�r��� b@9��`:�]��{�h;�5�5�a� �E�!H3"� k�eY�i���@3r$Hq���`t���y�4-h� i(�F���B�4�yڿwZ���ޠ8�=@s ��.�i b �A�M2��� �3 o���}��HH=�q#�N��~6@1 B`�E
4�@b�_~j���3�w���� � oԉ܉�$0H=$ .Q�<j��g2���P��",]EL�|��ى�w���n��S��=�(Ζ�N�}ߚ��m�VSP@�Yn�Ȗ&Sh�0Bm� M�эŖ�ƻ+���(�%x��'n�9&��-x!Y��N�s�cI� �w������ZS"B�b\L��Β6O	H@�@4��gM��;�y
�zs����Qm��V4�$JCI ����ݯ��fA� ߞ�ߞ{羐6��{dK\bGH�6��D��@ā��x��"iH��I]s��u�:����`�D�8��H@��������^-@�G%�$\����}5��羐7�z��@7�vy�a2���� i�D�D���A� ӎvێ�羐5���4P����h�=;㹒ژF��L�d����{�-���q�`@�E�H۽y�z��ԉ�/��4�(h+ �,>�$x �}.�e�b���[�L�ْn�ocN��hXܜ�TI�8�����C�<$z�q2�k�]��|�o H�'R:@c�le�2� k��a:HbA� �N��Nv��~��`�x��"U�@�UhbP�T�sF��@�$\����Z��<�� ���i��:�@ϕ� �Kh�VU]��:�r >}����KXgW�Z�P�-G�����\������	$V�L���y���b A�$	)BNv3j�]�<z�6��Ka�4�z��+2�`ɏb~�y������P�R#.h�])̟��\�Έ0��JQqR���������O}�Ґ�fa��9�������Q��{���5{�N�>Du�{���;����@��M�	-nݺ}��sJ�Ԩ�(�ow��v�X�9Q�q0�E�Q�z�3.�χ�� �>�� =�z��Ȥ��:����'�	U�1�׏���&u���H�1�
��?�jP�[�;��i$i9[Wu��u�d���6�s�}E%\ ��_u���RE�D*\�9��m��D"���������P���_E���}9�Z�ȱ�U�
}�R鷵zh�����=�`�&�_y?g��g&M�0�9�Ar�q���ʴɞ�3��F��s�ǅ�Y_�u�uD﯌��\٬瓇�k��1���܀��NIl��{�������ڛ_zิ��OY跨��^5s�.IN�Ϲ���X>���V�g��3w���<��W������nEiLA�M�P��E�|GO{9y�}W+}��%�)�|�t-���y޻��zw�ؔ�E�����:rju`0*r��S�'ibٶ���?1�Va��1��e��z��q���j���)�Æ���ۼ�")��`"7�b�j �JQj��*+�~jVJ �H�����""7"���@Th������((����F" (��4��%%�JR4CCE*�+C�&*X�bT�Qa1"R�%44��TT<J���X�P��(����*��ZX�"a�PDG�����%� �wvL�-յ(j�5����!���1���0#�LP�R�1Հ��åk�ĻF�I�X��ua.i�D�0��%A#K1�)�-�Y�ˬ��(����YfH�.#p�:��9���ַf�h�i�3��Cٙ�-]jJ \�H�lL ��d��rR0҂͊�8���)C�5��\�-滖m�i��s���tX`�*5���يhճb�6]������1�λK.tݺ�R�-�v͋�� �ɳkTI�X�m���\�0͢�,f��K���mvC�.�a,dڔ�27�KW`qs�6�ن&��u4��P�)n	CE&�X��XZ���-*Vf���n��bfkn�4%ק^XI� ��  �ID�h��ۧN�'��k
�isW�ѣ]k^�f�.�%;���`R��M) ����;��ר�U�H���]n��,rN�:�ɮ�U%�G`\%O>�[�� Fer�K�\�S�L�9��[�{{�=�0�OZ�W�YyWpojs�[W�1�4`�(Tn�.�ή�%B)-����=�i�ޮγ�֥�QVg���m:-@Y�f����ո�q`a���1���y�������pN�	���V��Q�z�L�G���D
�RN�����޳�=����}_�w�j1ɒ$�
����ܻ�\)����F
W�{:{j�D���*��d�]�kO�)�m��B�[�(��y��3�o_w��~�~��ҝ�,�D �o�e�Tw_vt�ʎ}�hԖ)��w��q��9����c<��oE�F�96-�+�������� �=�N<w���ޒ�ʢ���,�׺��=0�F���Ƥ�kj*]�^=s����u--�\A�����q�y�<�����ӈ�QJ5��Z�n�5��J
h�QS�μ��2�Tvзx'�Ns�p������7h�r]�ezC��{�+���B.�_� <{� O���PG�@��s���Sjq/hi�H�(L��a2Q"d$RW�Ӊ8�Oq�@���4�!��U�����xei�v�b#i���Ǎ��MO1aű�x�;r;��yB]$��r���~�%�o��Nm���\�:癩
����������ʊꅙ(���|=��� ~��[\�R��$ƹq�+6��cJ��5&��ڭ�ݜ\�ae�v�&�%.ll�e��mu6֚��[�����(��Ͽ)35�dT�)��2�baN}��_cr��hHr��YGg%E���^�U�λv�W	V����ű%�nUHV�1�r�檒	Bn:ng�[Ξـ���6�O~�Ɋ̮ZYpˊ@���}]QS�X���\c��L��E���]jz��,�:r���_	����{��{˾��������6"f�R�����3gG";7�b������mnEڄ� ����f��P�*-��ݘ�%	�٘��p��_=�=��>���z�Q�O_s�r��6ܾt�"��Mj���̻��Kc�Zfw��G�v}��fN�h���(
z�t��B*�j(EB:��=s�O��QD%���ǻ�Oҡ͆{dLA�kc���a,��L�9׷�5��y�z2���f`N+w���*���	G�WcZ�Wv��$����4@G6��}329��l�Z�#<#��h����cg� �� <���Y�*�ӫ�^K�yӝ�*J�А�A��D�0e"�2���ɘQw�Kk~�{�&�ݽʤt�QFy1U�
�_>���euU�J8�@ܬ��Μ�Q���N�)��}ϡ�v�dQ	BS��q*�<}�KHg4s^a]b=�U�)�eP4�K�k'�UPy*�@��nUߒ�$0�H�ecv�)	�C"��m��1��Pu�n��Il`��Z�L	1f`R�䔫ִk���ek]^��k`���3�ߟ��mK[bv��id�`Q-�qBi���<���nI �o��.���n%��1����&�s�m�n.h��
�����\�:�RB)%a�>uVo��s}��'[�V��S1%@�FD�12�$�#*f&阴FK���q�L�IJ���^���Bks�)�[D۳��KǼW�+�-QG��M{]�t��HC�̊̌P�;y2���އ�)$��ٻ�\-�������{$V8i@Io0���s�H�����V��*�Jm7�SM E2�-�8�>����߃oia�I�z��2.�O����y�Z��U����,�����w�J�;�g��8�N�_�M����Žh�u�;����2�ݒ�y�<��t~���mq�M��ػXW�����-��WU|���߂��f��D!{&0�{܎�;���W�~�x2f�y
vd����/��ԩg{�g��i�����6q�"�����q~�Č=�Q�P�OoPs׳��ׯNTS�Ve;�G<���s�R��h�˪��6 rë,�'�0+a9���U��15u�b�v������qU'�)�v��V�}��}�8s==F{��2n3J�^=����s5�v�n�Η��n��+�V����)9��R�5M
PRQ]����U\`4�j���cJ�D�Y* �(ҋ�7*��	N�J�PPTm�ѩ-�Ҫ�p�cDc9�F5�&��K�w��1� ��6�I�b@�R�q�Ⱥޯ�k������h
xH��wُz���%5*���}���u[svR�R۬�[-�v.h�g&0o�6)f ���V�T=�
�T�s�b켍݈`"�17뵕����0ԮN����E;͵�`�_U���QVH2�l]<��᧨^=Д�	��0�Y���`�r�\�t��{�t��Wg�E(R@ Rgn�͙͞>�?I��o��|fEo����H�D �����y��{�d�D"���8r�UO�:�O�gI���	BZ*f.q�o�������0��ǭ�ZA�`R��^�����ͮ��K�#�u�'����R_{<oq��γb���<sb��)������J��&�"�h *��
ZE(���)F���hh���(B�
����
��J�������xu�"��hg0Q����d�o�+&@j\��6�]qk��Mi�Z�!g ���Qv�֖͋I�G9�k�Ǌ�k�����{���-n��*bBD�BJ&R��-$i����k�M��Q�b�W*g����-8�%�"�_E+G���Li�T(we�B#wu�6̺;�f�K�S�\��o<bHeP߷�mJ�fn؛16����4�P�]\�]7���|Q�V�r:��DX ��i�[[[8@��]��Rд�D%B�QM4�����<q��s�<ݻA��<s}��1�FF�N�ǉ�	E��������}&a"�ށ�����,YJ<��߿~����$4ج�ͨ��nr�.�-t���{(];��Ij&���˽��x��IM�<W�(F2{22(pt��C��"�ьؚ��)�����=���3Q�)d�ET^�k�v�h��PG��oK=���4����'�xZe��@��QM�Kon�龽���V������P�u�u�bKWe��-�A���D�w��d��͛�6�.y���;�>o�/� ���#Lo�E�vʫ�<�|N�����f=��GPq޹����tD�9�$IQ%)�BIB��T%!3)W����o]p�t���(��mL����7��E3��DF�K!o^�w=��P�G*��\�]v��)�0�\V����!(�����U]FY�}�vMU�p�� �)�Z���liB�2�AIP̸��]@�	WTc-�R�Xfe�/1�s
l,��m,*gj.ָ���aim����ˆ���р	��߼a�7��k	��2d���$�+u�;躙AC��!�"�I잷���V�r'c�%�3y������P�V��(�#�W�[��i�4�	T�9�k�W^��,l��)`�Q��S ̨�"2����)F��*�k[����5A�ul�Ui��h��J��p�Ģ����!3�g��O����.ٓ|��(���lqU��g��T%i��]���m���B�����Tu_f�v~����ߩ���J���H&ɵ�2T$��ؖ�7{�sX��A��J��=�:{c|�<K�(��|�Uk\��ik.�Оɛm�;��!@��2f`�m^����^��wu��)gT�˖7��g^�H�����Y;����$��޻ו�M�i��1�Q���� q־��j�f�I>�����y��l���7q�.#{.ܚ�ǽ��$�(�տ�۵z���ߪ��I�oV"�F���랬�B��+L����#��u����(�hI�O>ֳ�%���j>�S2�(�&)�͂�+��M��~~����Qv(�]RTo����xݱ-:�Ј��a��kư�ʢIۋ����|�2�#��,z*Bo��f��p�%��E��b�ꚦf{��{��;�x�-[Ӝz��򾅭�JĸO���b�Q�jb�8:	�vq�X��"Ϸ����ֲ<>4\%2}�Q���q�=.��1C鼷���Ö҅\��p���[�⏱L�P��Q��^�c�wcq�׸-Y� �.k�=.C睜�y%i���<�=xi��n�|�:���wQ Fx�)�ɦ��m��_f�ټ/�c�s>�ա�1go���INO��,'
��Ms�_u
	�?s|��iNf����:�E����y��<��˷����х���8e������}�?��
��'�*.�˰T܆B
Ҋ�Qk2Q��4ޡ��%":�)�E^HrV��%(�!�^��w"4�ol�����R�F�Z޲�RMe�i-�B�3|s�h_/�X�J���2;��2ȑ�ŗ{�7ɷ��+�5/3j#�Mj��W��^������Z*�8�ܷB�bl��gd�6yԓXl�)�ض�зM�ɞ3���Q�bf �=T{]�@���mX��e��K��$�.їg6X�[{UR�����X��f���YE�v����YK)1�J�ᔴ]l3wWY�6�Zm�#+�l���m�,Y�v��5 #һk�9Kv��]�X[ZT.e.&���ۮ��J�V�qq%nP����� %���c��,,v�m�+\�F�\,A��/%���\,���Ӯc�D���JU��3,,�M�IV.+��a �Q��B�k0Ю�oy7�!cv�2U��Qu�!a-�0j�j�k�L)D�VukL���B3�2�=V�ל��  [�@  ���Stg+c�r?�N��w��[m�]�( S@��0!,�t5�p��qɕ�Z�4�	,����R]��(�1��2�q��v�˒�燇0��z�{���lmb�(�-��|��y�+/u��z�؅!uo=�}�3(�Dv��̽ǯ��b�Ԛ>ǳ��ˮ:#dB' ��+g{������o�0�iK)�6w30�s����j�������tc�K��"�����*���{�ٰ+z�P��<����5��l����Ȉ_n�Owc�K�}2}�;����
'0���������/v��D�i�a�A��ƗQFa����ߺ]ȧvn:&)Ul�}��-�mE�/p=[�8�D�=�I:U�ſB<��fJ
#�ھ�zi�I��]�v��7�OF"""�c��}��b&�HP!2J1�����0��y�O[|����G���"����6[�������`�䯶"+�s�d��34"#]�_7=cb��!1up�`�NsβX'�]6�Q�x���H���5�șw��=��ͦ�`�.9cp���b#o�{{�\��>�^w��t������Kޢ �#u��*��m8��E�X�����a�L@�"'+����Z�l���TdE�[���b�o����1b��.k�(�|.�D�ّ�fV[���-ЛF�Yk��R��]K%��`�z�ڨ��\Yv��3/0ZWgi�Z��6I.��q:�B��Ø ��������%R���e�r��	�sm�v�<�LwP���:�;[�Y#S�Ui�.�ƺϽB�gyy��s]��sW��DG�'�)f]���Zy&�|}�Mbb�Im���^\���)	�K2"��^�#�7j`�奣]I����O���&�g,�w͞�]H��Q_g�?�^��&\ē&���U㗜��Y�����sw��Y��1�V�@��̹�珹�5�F��odH^������3�z��V{�KK��}ռ�d�>NO�Q�H�x1tXæ�����}d{�:.��T	'�|��qVdC�J"�7��VR�((u�R�B�v��� ��չ��O����������"�!�k���SX�s׽�0���V�"�mӻ�'-��z$�O��Y6^���u���Ԯ�k O�[��.�F����w'�Z�W`ij�-���wX[�Nk�g���<�^!_n��a��@��.�g��^�}��Qm�hD��fi�jUK�;���]��dL\��)qr`�k;"$H�̛5��'k:f����|��yG�QA>G`GDN����A�I�8��<�U_���bm��r5$�����eC�ZWӾ�=�w�.��mZ[B>��ٟzȷ��n��dzO����Rm���SG<w�v��s�<"��U��{/4�v�\�o~��1�!��fd���GРA���ߠ��U���O��e %+-�؅P�m�U�Sqqݷ����j�g�t�	c���G�o�鸊5.�[4E��+k��
��n�#WMA-�)�;�l��Z�4�J����8�/^֥�2ks�d�br�k�`f��T6t��|���It]נ���S30�G~�G���P }������EY6דM�6�Pɭ}�F��A�׷����Us�{��vvĶ�ӓ�rk��{���Pƭ�QKNo鯵ī��K�79����z��#�ަ�4[V�(
� ����n�5��=�="8_���~Að�l�Y\́��>j5>�R�������>O��[�DP����E>��l�����Ӕ)H���e�&���(P<}�<�c��fO�zi���Dn��߷>����7ϺgҾB[V��sn�5�M�5��Ͻ�k�2��t��*ګD���H͇�ϯ�7�#�a�w��B�bTB�k�ܖքT���Y��K�L����O@U%q|$�����S�Q7}�9���y$m����c��ڍ'��@O����~X��%*��]t���ַD5v�~:=���о)v�1����J�Y<�wP�9e��M+�X��]-�XO�}�,�A����9OG�C�{T;�����M�NM��s�)�M�+���yHSگ�iao.��ܗ�
g���M�u�zڏ�2.�����g����tM2�x���:����v����<��X @}�K�yU��1���#�d��I�Wb�ZP�p�]�5��v�P6�{�_�8-DV|9<����mc�]S2��5�s���S��U���#�d��#��eG���d5 �|�Q�W�
��D����d�$1"s2�%�q�V��V
�%Ȥ�d������n�bZ[ض�-�D9yu2�ADU�5R�m ���r�d�C2��.�-Y��c�A�uv�]�� K{[}�[�x��Mv,��
GO��:��ͭ��lBЉ���e�o�P�&L?y�>��)6�v�F��������A3���ۮ"H�>GȄG,؟P��on7rYR��O���N�����au.�f �A�LL.��|�T���:��m�O"5i� ��7Zt�3�k~��4�P�j��z�SBmZX�V���=�{�o�)���A.J��耈&��@���υ��ǹ�$�+6�&ٹ֮������ H�_{�g��F؊	p����ޢ����Ͼ鿧}�Yz�K�,�Ϧ�e��c ;lhh�7A�����e��׋<�����=��Y��kF#�A�%\ ��;Ͼ�S�>�&]Ok����ֽg�}�"ͱ�/8{w��{��o�_$E�`�� ��\Ll�l�>�!�.y��O��jP>G�@QDA�Gz[���40.}1K�����:9���*���c�z��,�>?��m	�E�(?��4�� Z�E�)l�2iKi��.E�*���ݰ��3�Ji���R�A̻%u������xs 2�g��~�t3krVg3j�2�!�����6�{>�����κ�*8Ĵ��|�)��M^�	��9��w'�u6�sXi�bX�mZo�7�w=��룍y����9̰�i����w�s�g�@��ez�Ǽ���ۆ�Č��o���Ƽ�jU����޹�/�Z�-���up���{��g�ׯ�}|��z�V ��|��� ����7�U���{u����>W�=�`���9�^���*{[z,�����'�Gңހ�+�ϐҖv�:��A �yA ��qjϽg�E��e�h:`�y�$i�յhZA��ʱ����w�4�S��K�o�����&��n&eA���r���е�B�w\���{X���L�����]j�D��-/=f8}'wk��,���u)��A�<��C2TK�� {=A$/���� �7-^U���2$(;�����(�H��!Oe
6E �|T�ߩ�s�h�}��E-#iQ���I����|��}���A�*eWJ�rQ�P(�b�3"�]�xƴ��%[h�7�o�{��r�O�Z��4[Ĩ�uQ=��_:����7c��r�"-�-=9�5��_{�G�jڴ5���jӍ��k����Lk�&�VO�ϻ�^�#�i�#����[|~W�Ϯ����7���L��ko�"}�V��,(/A������#�cȢV���0�iK)ؒ�,��q��Y��%���w_}�<����=4��DY��t�߹���LO����ٷq�0{��E���Uy�σ �(����#�d�!8���G���gJϨ�>��d�רY� �珞�}�qǤ�L��O�2-��"�^�s5T��C7����U���#WQ��F&4%+�ckF��a^���]GA����G �(�� b���WS)�iCY�[F�Q�dE،̮P��"���}�����.�hZL�d/&�]����G�2�bOs��>ｭ5��/�q4툸�\����m�������Ymq��@�O���jCMcV�X��2}�}������'�ch� ���ǹzt�@�#�Gf\�g:�ϱ��{��-�Q�Yr�"9+8�I�s��p�s�$�L�fq��1&$I�����m^�Z�<�d/z��n�͂�[�z ��5L����G����]���|��4/���,��k�e/�j������;~���g�|�c�qBN#�"H3��3W6O[��݀������c�}7N���g�|��+�[��|�{���xi�i�\k��O��[y[��Q�8`�p ��=Gf�3�R]��K�QG	=Y�a��)�;�s[B\�\}JrS��kl�X�c{�{�{����<����{�9�d��DƱ>ّ���ڕ�>��ӞR֯�/z�R�;n������7T}���!0��T�r��p ��z`EN���З���r �=G�Q��I��~�#�o=�}�oۛ͞}����\��B^��%����m��1��C]��ϻ�kMfK����ZC���oYV֓����I��;�N�U�!��DǤ�&ob�!^v��$q� �}'�@DP]7V}D	>��yu���>���:x%}��6��⁾��<�ޱ��"cno.V�5q��[�Yf� �O��ѿPځx�:�愐�� �.X�lWS��ش��&5M1r�j�]�x�t���!b4�{;�{�t�޾�GZ�y�8��D�Aq�}ޖ����"�*o�]Qg�}��R}g�|�0 ��L���wv�BHg���'��#��p�ϰ�"��o=}�4�]����q�]C�3�ϻ��wx�����ϰ�Ϥ�L��Y���7�V졎5�����+�V�*z:xz��gk�(n^����v��R��}ďP�I}h�Fޅޫ;�<+>���t��{�\��.�}4aZuw�v��ÿ<��Nm�ўO����wwO>Ht��ߗE�:��Z�{w���7:�ٝ��Sк=�$�b���Ⱥ(�`��3=�M�����ܙ!���}�r1��b��G��{a��/�+��U+���}�0T�1��{�Ǯ\���f�����tU'r��Nm���{������n�����==���=�Bջ����[�l����7N�$��'�j��D�-�V����/���[J���B�6�1�9�S�T�ȣJ5֢VIH*�H�:���qA)<J��5B("��1UTUX5�eYƢ*+B��-(��E�.�V�Ң�Ljҫ$ER�NB�k����m�H9��E�Ur�;���jYZ�XB�L;vH K#֓B�Z!P*�-Ѝ�p@�[iU�f�m�i���Km��RSKce�,!uن*�f6��kdu"M[�f�R�A�b�F�Z��Y�mh�a����V��R��"嫈�0ޮ�n�SVR�i��.�kCW���[F����K5�a�)l�v��쵋m%�b	1�,�yF�nԅKֶ�u&]�^kiIi�� �J1]n��܏-&r�n��J_-<I���B�=v�Hj	*R�$ږ�5n���%��ŭ�]of�����ٔ.Ұ�vֵ��LR:iH`���s.�]k, �����qt�q�5m��ԊV7R-�Z͠����%f  �\  0EU[��u(��X۪?�C�6�y)uٮ�i#���]Θ���5��f��!�:�K���:R�-�T��.��WȲ��uAРf;����5x�� \E���__<�gi��w�p��C��[��g��,l���}�}�5�u��b<���0qm/�;2�E�(��[�މ!� 2�j�$ID>��x�x*�_.���s�ȼb;��cV����m6��� l�c�m
q�0F��*FDx�zH}i�;�txۭ����鯠�R�`��S��m��(H��)���$)�E�>��";]v74}w�j���̟I���� ����T��6�.�E-���ӳ���ty�s����G(~ e��#�#�^_���(�O���Ǥ�t�ML���8���w���w���5m{![�Ӷ��S��>������!������X�Ʊ,qkO���NNmf>�G�|��}$e٤����ʓ1�e�\ڽ�s����?'����}���t�s����p���@��I�\H@���;v����B񉤎=�Ma�ڶ���JƱ7��^��k�r��oB_ND?gz|T}ۊ�4�w���T��7���	��!13����*`�2�&L4����{�w��յms�2�c&������"�ν�sE�NEG��2{������ᔗB-�������Dz='�F�w]�Ȣ.B���C�d�CN�k�#�4��{���8���N}O����X��%9����n﫷y�}��}&H ɂ$��$�D0D���)�r)�'��m�����#������|�d�rer-��2Yo�\���5m~8�rV*�֌�����������!��'�E�Sq�KU)D�)2���m�npe}Bϔ��t1�M{�޻��4�5��q�!��� �YezϮ�Gun^�r)Ǵ�. �Ϸ�ƴ��k�G�v��j�=����ԉ汬LL���	d>S�o)�sG��"���I���G����������nE8��"ȀD�@��ljꂫ������&�rhR$�a�zy�����8S*�D�I�-���N6XR�8IYI��&�YcX�ku��6�-��>2H�eʱjbs�i�خ�glj���U����s +�������Y�MH���i���^1B8���{������{ؙa�"���>Ff榀��I��[��f�q��Ƿ�,]�6��ƭ����f���"���,�*='�}�R'�}&���5y���j���p� I���&'js6w�"{����0�O�����ߧ���2$lR��Y,�e��~-6�"<���&���_s�a��ھ�y&��B1�k7�w/}^������k��O�|4kV>z���b�>_���G���z,��3�sD���ԕ��,L��G����k�w٧ȏX�kEƲ�|��f�ƶգvi��r,�t�𨾚FD{��>��9� `8E�׭��>�$Iߎ��4E5�#���s >ӤaTzH�Nsq��Ȏ�;wƁ�q����b�n��}�o�w�{�����޲��6֚ķ�8�Yл�s/TM�E��F�/�-׷n�r�Ѥ|��޷�x� ��If.˱x|�}37+k3�� adU�3����Ʊ�LD�X���a�37���о�`�.'�B�KՖ9�B$IY�6@!�0�r���[��%ohd�S���Fл=T@���Q@�#�|@Ѳ�0��w97��O����d<U���N@����#�b{��g��y�t/����|��&�li�8"���xǏ��)�soE��OV
��'�;��(�dWr$EFE��1:Ʌ��_v����L���C3.��ߚ�9�~~kMy��G�^w�뿹���X1�/\���Q�O�����������=��>�;ѰI� #����5oOs^��{���|�kK�DƤ�$�*=$l��g7�yݽT|���q�cYp���DƱ���������sҺ���n��n�'%b�cX�!��z��[�n:D��D��⑛���.���ػ�:���h໊���{�c?�mH�!3�b�C]����K�	Z,]��i�N.maC���f�5��#Bl��c0vڀ˳DQ�V��0l��G ������5���Q�W[�SS)�)u����}�o\��{Z|���cZj�k.�D�q�Nsw�w���zֶ���R���LH��c�����J�ұ��$L@��p�N�j��&^u�v�֟"<b_ə�V!�&$q	���dqD�+}��a�Q�����{Ό�&�iJA��7!��-u�Ԏ!�������ޯ�:�jڴ�������Cg�=�t�N�엤�f��uK����즻"Z�� }È��Q�n���U,�E�I��Q�(��
`��LL�e�.��w���J�P�"cX�>N(�D IEmvkz/��|��߷V��2\bbߞ)y[9������֐�^�#�Gއ��6X��ha��؃b9Ǩ^�d�=麷PD��۝Ǽ�a���~T|�|����115نJ�V��^��{�����߽�og� ���DƦC�x��&}ng��S��>!������t�=9�G�=�2ч��!�cv��;|�=c�`H�V"�m����¶�ַ,ԸX������ؐ� ��E]����Ć�u��@w[�bm�{�7gLh��Yջ�V�6{�5p��U+X��
;��w��I�s}_�m�6$Ϫѹ��A��i�d��}s��J�0�;�ww?{,`���,H�Hu$��6yc�rt_=�k�hu�������+�]����4��dS�7L����{���Xw�=��!���b���:�8���Q��<;�C�1��v�hP^��S��q���R����IU�"Ч�)J���(�J�䪂��E��Bӹ̘""4"U9+WZZF��b<�j��D�QN&� �-+UF󈱃{0RVֶd����s�}��{Zk��i#�G���""��|�˗�y�� �>SՔYq�c8������y����7��5��4��O��xO=���cB������s/���u�r5fC��y���֚�U׌�#r�ո�Y�H��3�(�#n�sq�}g�@Y�}g�|� �zHr��4�w��8�zO����>��!����uD>����tN�b��H☢�}�y�a�~UV����>kH���}7=�," )ܬ�{�}g��A}$!���X$5i\b���O^�x�+���k��~���C'�.��Mm���>q�t �>�eek�4@��!�y��L�ݑ�X��DƱ�LϹ�r�rmwo:C8} I����e5�NB=`����{�6�������B�IO��"H���������4|�"���%j��������a+��ի�ݚ��Z/�X�T�<n"%(M�f[\l�D�F�v��Bm��+Ihm�a������7��=Mt#���Ѷ3:YHW��� �������%��4]�/�����;�� FG��Hz�o��A�oӬ�rS���q�e�5c�z�s��x�!�K�sD� ��='�@��G#ja�0��{yՖA8}������H��i�Ns���������n�K-4�5�؎Jē�j�[a����E�{���zO����#U�đ��bD�BfԘ�z����=�$�H�O2��:��x��F@�f��"H�$A5�;[�:�NIѕ73(���9oj�6'9Vj�1��>����F�{�9�?�Y��Q;��f��>�� ���I1W�ݸ�_G��!�I�D�W��F1G����Y��Yd>~Wu��t�Ď!�c{��Կ�0�g5�}�΅��Y�>�!:���bP���rc�WK.���[��e���u�7�s�}��VE��kN	�$�j�QӤl���G6��� Y�����3�hł�8�`{��w�!���m��ѩNN����=��K�b>���������P�6�:�>Ĝl��:�y{Ya� J�RЦ�faK�o];2�ɩ�ڏ}|�=�����L���j��Cz�ꢍn_c�v`�%Ê��)$��cҦcg{��4�B�uQe$��˘����ْWW~�v��w�u�b��|��2M�ǹ����Ad�݄�Z���H��u�Y����_>i
�A�6��L��X1�Xx�4�wQ�z��{\��TdndBD]��3"�eg=�x��4WL�몥�\j�_;�i��\C�(��F�e�|�5�Z񨤢��ɧoq��h�1]V����f��MT��XU�V2��9��`$g�e|ls-.5�x�i�\[qa���t���t9��.�;�T�$�z^^B�:$E�Э �í���P�Cjں0�u��jOg�{�ypѺٹ�IJ��%"fbg~E�Qkk7]ł<�$���+Ĉ(�w���fP�Ⱦ�À���=4�k��x�EMM�ue>���u�(���v7�v<�����������Dm�ј\G#��
T�J�Ñ����n��T����J��5͍�kY�"�h�˹�hG4춈��&j�vL���=N����=-w5R�ِ)$�mK9�{���ܤ�����}fʺ�{��?S�=F�H�f�@"�^�Pus�m����Wp���ґ��*I���P$D�R3*j�8��^�k�$�R��Q@����9�KwkfF(	:�����jaqB�3ʼ��7�6O�w�����\�T=�a��j�o�/�Q�[�&`b��HmDu@"�^[�玏���i���ġ"&I!�$@�DAJ������gs\,��PE���"ϭ���sLJ��@^��) �]��n�玈��Zwa��۷�����Gt�j��d(�؍�օ=B��1�*�@�oĐL�}�m$�o�=J��>�\�"T,����%DJ ��aĘ+�Qi�)ߧ����ݵ�Cq(ꌇ�j2����=!���$E#�K�226�1�r�\��*
�*�^�v蘏
0BI%�f��5��[Y��T�æ/(�u��w��n�.=V�oMc�����5n����WE�.OT���v����
�K`��n�;�޻�'o�=�[�U�,�]7=��ޛ���I�V�����C<�ۦd�{��aǭk\󸎞�E�g�L��Ԝ���W�d	c���;�(C��g��:�:x�' q �n�vּeݲzf�E��8��2QY.�^YC�%x�0�c��=�bo�o,���G޻�������;��ܴwqFv�兡�����y�Ɍ{�bþ �\�vV���՜3�^�Q�x�O�B���&�&���$�z��9C�{�r/u�C(>� �|
P���Jw�5B�B�*2E�U���iu���Z
R�"�-(I�2��;J����TiQ@���!�F1���`��V�)j�Q��J=����%+�Q-�դ�ZP�m�� FJ��mR�"�%ZR�S%bh�KCXhi�����ӈAV��J�Q��2'eG��^�~�
��mL^�ց�������":ܵY�e��z�G��;m�k��<�v7��M���Eml�-�x6�Dvv�uѰ�m�i�Ya�Sa������b�en��m�au���L�V]�m�*+�քq�U�ֵ��k^��t��6�-,++�՚iA��Ʊ!��F�e�Xo[My��2����*4���˨8�=qq�t��ev�ƶ��Zd��GY�����ap���L(�s5�i�6�hD��i�p�5D��.�ݒ���B��s�XDݱX&4I�9���ԍuV����̬@�Ek�h��,�)JҳK�RV�BlM���Ү�V1,�,��#n�� ��3e�jq��^#UUT �k�   �p[rۙ`GM����C�Jv�[ٔ���Aj�+��ݶw��|��+i�-ŷ:�2m+l�u]�l0#\FY���YwRc%f&c�������3������4�.ŭ�#
$�R%-�4�P����}�o��H��s��E�w��������*��b҈D)�ȯܧ��[��W)�SR�soj�BE�w.��i�)[�L�k*�$��%��J�\��k���N��sNM]X�M�"����f��c���^�Ĥ�,޳�yĩD�H��R�x��d�������E��Q��qs�'.�bjH9��K�@�\�V>sy%�P(��(J.�nm`ҳm�|�䤄D��ϕ�ڹ��PtAU��梅%��:�u�G15i(JL]���#O���7έ�յ�b�V%^벏��R�V��b�t�-�z|F�{�����ͯ�J�Ȫ�>����n��;ɖ��JE�\*���~��+(��f@��WK�ܲ�fљ�7M���W[���s�]�E(p<��5q]��5�N��-�cّ�N�
o>��U�e(V�υ�6B-�nws�0���}u�g�V�l�{��.?n�zAg~�A\���S��$�ܷo��/������� �>��D�!-��l�Fٵ�BT�i�U�Y��=�e:�P�9S
�5]u��\�"JR6�I�Q6���{Γ����в��:��<(�2�P+c�Or�����MMk5)��k�F+rl����$!F��x����duX2���k4&�%u@�Viw[,q�Ŗ�J��n9��5�A֌��"��/��`-��î��JFe�%�UV�gϿ�ɩt�Gc��*T/L(�����;�ǛΘ���E�H����J�ɻ�n{�CO��"��R���uv7�m4�����F�/�kv�n��0�e(J�VáP6�B��m�~�?"���5v��8�������(bQ&B�)ofUk����j�����#]��1��9��ҋF(�Yw+e�`4;� �:G��k�Ե��n��iD"�n$^ggk�� ��']�I�Wy9|���<z�̌J�F�^�y�����o�/�__�K����3P�%��F��313��+��n[�BƸ�6RR奄����+��9���vN��ʥ iI<�R����ӳU�VXc���z7�V�砌���>��_�M%&�ɔE�U�6�9vBv.^@Q�+sUn>��mD;v7^𘘈������H�S0L̘��7�Q坷�q�w�{�	B;au�6g7j�[�,�B>E�IEI��n,{Ϝچ� 웠��y^kǸ�N�蔱�;Kj�ٕU�v�i�5�!��q�5�����[�~����9v|�(\��b�*�fd���!L�L�5i!�t�_9"٘��N�UA^�ǹΘ�Sy�0��p�rs ;�ُ���B]1YbM�#�t��9~�v�/cT"W�W9����:����ʣ�?�K�g�����vz�
c��.kn�̻*P���'�����RH�ʶT��% �8Y\�Ɩ�Y��Ƃ�ڹ�W�2���⊽keq�uhl8Kc�,�hL��D�y�����{�����M-R�.��kEL}��R�ɾ�r��}ʀ�R�_U�e�"�j���J:-mx]���,'Ѯq�n�/���(G+j����N ͟YJ
�W��+�t��	)o�37=���t,��ʸ�p�j��9�n��[�]��Q��[�m��9�A �Μ ��]�j�̕��~�����}4��T��QE�3c���k��[���e�Y���Syۭ�ݻF=�i(	%�\�`Q�ٹ��Y�(���צs�*z�M�L��Xx�4��J
{�����aJD#�= Z��y��Ο��wB��AB�ë�SZh2z#*!��1aZ/^+\©/��qn��W�
�'3 �����w�������[ݰw�1�;���{=���-�.��;�������3g�9���x����I5�{bќu�9�_�������U���v��o�t��潬j�����Ӈn�D�E�w:a��r�\�1޳�p��_+�X��̏m������$>H��%w�_��R�[/
��G-�^���A]õzqN����9�=O�Ns�e�jK<�?%�䑝9�#�#A��dg�ʟL���Ő� ��xN�Fw7���5�O�ZZAF&$�"��`�`�D�Z����PC�b�!3&үp�R+G��J�"�B�;����PiE(�Q��F��P��X14������9"��:�5E�J���q��L�k�(-P�-QlEM��$)h���������O�~�ǜ����A�
Gv��>t��W>7p��(���yΩҀ�c��׿�Y�j$�1���9���EFwU�79Č!�>E,u=h�y[W����%m�/6sca%���x�_s�tQI6LQ5KZ�{�l���9HĞP`��p(g�����ê�7��y�ޚP��<U��Z%LDD��)AB2T�3&&f���+;�cs,�I%vx�t1Fs��9�-B�0��$�QW��2h�`�R�o;cM���e��D�!vk�xܱc{�}�i"�w�G��>�ܼ!�IZ�8(qu�H������דЯ,-&ƞc>.�B@��Va�0`ئ���UɘIk�Ui��m� tH��M���WUٲ�f3���^�"F[���aщu˨���EUU�����c@C)]��leB*>��"����v��LBRIiO5aE���������3>E"����o/���I%�br�n��W�"��Up/�v�7��b�%�;�����p�m)�n������"�r����
<�"1e�C2�URߞ'n �9�^Kx�^�|cx#�ʃ�}c�ɯ�z���XH�=1�t�^��zܻ�Ew&f�H�M��簧�*�(����|-L����(].��UGg\��ģ��,�P�{��y��ռ�,ufL�!F��u2* V9����auh�%xE��.g#
�� �{f���@=}��������wo6����P�̑SB��}��b���B	B������;��jmU<jʋ�Em\V��b�=���ߧ�^�w��a^S�#!(ҧ�7�]Yۍ���^�_����GO=y��j	�@ɉ8��{���R�����p��w����sw:�׿�v��K�� �H{[�m?a�W�dHۺr���J��([s�穬�����͢�������)���sUϱ�"S���g��������sn7��X�(3*���=ݭŻ�A���(�hnX���=�w�% �n�d�vf�t������%��{B������?��� ��F�����R�9�C�%���E��D�f��D�&el�s6�mH���-%��0ۗ��W'��uDs��F�9��]A������Gm�Ӏ��L�C$ɉ��q����{��/�<;1#�Y�Fjys�n�9IQ�P�f�n��)Qۙ�P�̝oq���V�bB!}#h\��{���;�l궗J�lf)eX�eLE5��<}�����(N$�,�Ξ�7x�S�œ�RUX����	���&�\�v^�x�y�t��`�D�Q�ǃ���ؾe�Ƈm3[�������3��.���a����5�ʞ��2�c�@AB2�&W�B����5�����\���$��9!���}���/V���IJN���Y���@���|�zV0�4#>����0d|.�i�s��RP�)z�L.ٶ��<�fH������Z19���v��`�����-���J)R���!V��<�/���@#���٘�]ُ����n�E�l�������CP�&�rq��s��VĨ�]�s��3Wco+Ғ ����E�\��Q�5���8x@e&nD%�AI�)���knhІ/zNo�p�f�JP�P�ڪ"���gkr�Ҧhu�G��s��j���(�S�fFU���{}/�7�h�y�|���u�Y�}1��G�{O�'��*=�1b����, �*f��� �*~x�@P;0��$N��LC��d3��A(�s��~����<'څ�P��� � J�l�e�ֵI�Q(uP~��iD�B�ϠN��6qx�CT�0����Y�P>�����q��o-��N���Cp�9���e��=�e�t0p?�w��l.��V��Ŝ����Y2������􊀩�a:��O?W�y����ފ����]�D?�b%&'�=������{���]����j`��?�2����GP��|�l��S��T����=��!���U2��JdT���\hBn�{�j%ȟ����S禉�|L���g�$�C|x}�,�װF��ȇ�Z�@T�-L=0�[u�46�߆�� �*h�m�ʯ!iT!ƣ�&P�0u!��C_C��sA<͐�����>�O���\�`�!������#�?0MS���㇑�<��I�|Tױ�?������z�����Ϳ�L?��*k�,�eX}�6>Q>�y~�64�A���HaL����c��z{~!�kQ�]A�A�. ��3௣�������>@(
�@{�`��~P�����p��#��:����0N0��"*
�FC�A@T�A���G!j~����'��r~C���^>��OP��9T�6՘��z.KՁ`�ŭ�T0��au��=g�6]@���֗HI�qb���[	�v���BÌ	˸�hp�+��@�&�(
�9���#�;�)�@T��|E�p�`�~^@S�����:�<�c����y��=>������g�d��x?Wa�z���O�G?rz�����������Oi����<�0��1����8K�@T��:���r�~�~�ra��z~=���O>n�	��pA��#����1A���|�_�� ��y< �7=��?���>���)��tf�:|C�`L���{�4�&��bY{�ԓ�>{��C��.�=�`�����lz�5D�:�|{OT���� ���@2�����G��o?Q��E@T�/����C���{���][`��2P�3�M��Jb����
zvx�����]��BC�1VL