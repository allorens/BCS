BZh91AY&SY�3I�;�ߔpy����������  `�|Y�H>�( �R�
$  �@(�w    �      ��}$�TUJ*�z�� }
 �I��T(_��.��\<c�g]�H��t ��{�>��C{�ǧ��t(]��(���v�N;P�  z�[����Zb�.�]��}=:d�V�չ��TR@{�>;�}:�K�k��흵ޜ+���
�8 < �|���6ٽ����{5�:9��;�^�l <��
do>8=#�]������{iV�  (�}n����K�v�pa���Lۧ{�9S^��|j;�l_g�sY*����2(;�'� $w�r��Ӫtg�^�{T�Uӻ�^�K}u�����I�ͻu6�o�����o7n�`�     P     � �S�c�*�&� ��0�&4�`�?%)U=F� 4A�ѓ5?"�T�  � L@ %=$j�T&a4�`0  $@%PF�ъi� �5<SOP�M<P �U*3&�	�F`ѓFFM��7���/�u*���O��@O����(
X( �~""����*��~�	������\6�U��y`���'h�Id�:���̶��� H�H�Y�ɨ��m����U �C�����	?��?�g���z,�����еK�^W�;ԄEJ�R8�>�Z��a�D�>>�� ԛ�>�k���(����<3��0���Q��Bj�;��c5�ca$�}
fԌ���4�T6X�����3��ny/5�ݎg���ܒ\eIu֘�M;�S�;ù�6���2��'�����Z���'|/0G1��NO�fx�2o����@���~Y���F�]�>��O�6^	��UR|��j�kN
h����s��}�U��m
���im�U1���O>�mݮ�o��m艍��q�롼��f��p�|8٨�6����m4qt�R��s��O/S�:A�G���0�K��Ò�R�+՜{��3�զkn�*H����5�nՄ�;��ǲ䬪��6�[n�m�͹eӝ�!Β
���Iڒu�����rk0���ގp��loZz��ɎN���8[��l���a�����8��/��*�Y�Q':����[��8�o��lXе�h#{��qǫ#�Ȼ��[o�}$��ە�7��q[�ց���P�|�&s�e���`�8G��}�q7W�����v:��0s1ݾҸ��xc�m��1ɯ��c}�S1�6��p�[��.�8�hƍp:9c�f7v��]����4o�cz������cf8����'1�w��&��4w���sx�X�V�]i��c��N���r�ݳ2Kܓ�Mp���"�E�URo9!�91�x��kBЛS�ުj6����5�}kF��I&��>�͎���'[¤Ӓv1�d�$��Na�0����-��}�U���;lƍsA��8�c��gk$�7Y�:7K��6�������s���N��R��s��O/la��;��y�f�Q°�ʔ�ez�3�O�i���̒#Sx=rk�����$��9��\��R>cm�]u�̹e¯��K��&�-�WRV$�9A>�ӮMfYz9@��֞�1�c���-��;o
poF��l���F�MZ|�P��_|U��i�R��{
prk�nJyL��1�bƱk@�8F�9��$�S��8k1�e��7�N���
�*��qu��cc���u��I�rL8巃l��o)�Ӊ�6�w�trǘ9���&q�:-�ޘ�[ccLrk���-�x6��p�[�����Nq��SF�����3�r��nXݘ�7��o�-�yNXӈ��>͐�!͐�9�u����Ώx8���4մ��M�pls�9����T�d�l��+�N(�6����(����iІ�4&֦�6����l�s���&�M#�u�;)ʏ�׻Ri���H�H͌$�I0���/y��en������m��b(����x�|}w�SԶĶ�(m���|ȳ�8>.u־)�W��pT^k���O��s����\�N�N���>G�N|ַ��86�����"���J�L�s����\��l��6N�Hts�T�+k�K�Aȋt�c��IX�G&�մ���-`��cLX�|��ې�9H� ��>���iέ�FIڷE�B��qaRq����9�C����6����mҥ��G:����D��#�|4ֶ��O�4�GJ�����Y$�8-.M-�ӫ��\��l��6B}Hj���S��$S�E;�8c����9�0r��M���1�1�cn�ې�9H�!>�i���{"�s�#���FI��'��+�%��irT�@�T��[o���w�M���oP�B���]�:��8u�Qrt�&cbeɝ낼�,�f�f�+�'r9�v����:��	�>ϑ�>{X�>��د���9D�O���a�2�s����\��lU�͐Pqm�Z���$��w'pTwG5ffw��Y�F��3�6�1^�:�(_] ��d��>��Vޠ?P�z|�|�|�|>!��C�qt��߅՝R�϶�X'�`�0LU�{lLZ6�Z}�:�)>(q�O��+�V(�����_���;=ݯmm�qV6�i��n�N�N��&�_i�d;�R&�Aτ?�5�eH�NuC�p낢��-�Ig\�����%��d���Qڐ�\�ӗ!-Ϗ��φ���(���N������s�,$�q�ir��U�s�Du6���&�AϩcT���$Pr(\�1�PI�՘He���Z�m�Ϗ|����O}/�0�+~F�z�㍝�gx��h��J�.�BV,z�1�bb�[Qjx���Ct��ߨL��Չ�`�0LU�w�z&"�{�>��l����[��}���ʾQ�M)<��������y�m���f��sD�~��ބ�+�Ro��p<i��֏�B}�����1��<S�������	�:&*����HO�r�[�\�'�Mʉ�?���N��o񍤷�,�?��->�#=s)��3�`%��B	x�A>|mQ�����I�q��Ho���)��Ө��,�����)ƘsN3�F�:!��9 92ך��F�9Y�).��E�����_O���9���#Z���Tn����)�b�q���[X��fA;u�5KD|��ȢA���<"W2�"mȚh�s�ݒ�0�8SV�+��;P����;sk�}77t��\�.���V=�3u���~� �"�ǖ�⸶����z�*��ۻ����{(_�'ه+��Y\MtN��Ҍ��X0�ykhr�M�{�� �����Hv�"���r�1�L�3�c�K2F&Jǌ���Y��#�l�������k��$���CJ{��:�9^��~��vs��BOsY��t�3���IX7gW\�S�󮇓1�[����ʻ|n׉��a֋����"�{�����}��hynA��Q�[�ҽ٥l�+Ȼ��jM�o[�ߤ��޹�WD_�������ӹ�뾞��dAW�ٴ�v��ǣz�M��O��(�p�&�Cᢑ���b/�e�9���R��2U��-�ㇿl�d��o��{��j�y����מ'���D��w�����5W�Gv��h闈8ot�g�b/��n8"2%2Ma8�N,�cXA�=�[)X8�Y뮼	�5Hw$l���{5�q�)�����jo� �2�dWOv'�I�xl}b\��w��#q�&=��77ِo�7��lzͦ�V'�JL�Δ�*C���S*D]�5�z�n�'�������U#z�������6H��1�9��Z��ۍ���������J�=����i�*e۟�	��(�m�(��st&���m����~0�!����c��0��	�4�nk���݇������KCԋ��$����(5z]��Ռ���~�=��|p���[�Q;2/4I/%&�O	�Nj��G��J;̨]ʣ�Xx�<�@�7���|��ἜE'��r�wsjY��8b۫-��!��<Ұ���W:ņ�Ϛ%�f���}���2���eq�sl����J{m3/�Rr��
O=^�ڱx-9�Oz��<��=�,NY�v`^L���r�e�(�4�d��#�R�c��g���>�7��|x<�ve�҇�M6!2��͗�'t��F��3����$Qr\=3�F�O>ε��ȄXS��s��j̖y1ۤ�i�s(�r��2�F���8���ꛗ{{B��.� �i���������e��*��N=1��f��`g��������m�)�8C��d�#�2nc[��xY�EyMk���G�R[~k�k��0ы��xg1/g��Z��}B0���ٖX`ʆ"5�VM�5K��^�齭��i��v�aJ��>[/%n]>,��'{��6HkS���wqʸ�R�p�fr}������t)�>�wfi)!���n���]��*�������Ri83W�w/����8Z���)ې��Ε�t��;	a�?Tk���(�\�aN�Ma��#���׭r*�)��5�<����1{�L���$umos؁�
��B�:vwR|�wTo:��ˆ�e�@�#���2�ćn������=����$�D�[�+�9�	��=�}��7�Y����k����#Jq��4q��,����n������P���|iOϮ;���I�������7�30ޟ,(�� ��K�2P3Aq�BPޙ�m���I_l���Ka�4��`��)���l�Z#���~=t'L���ܢB���DZnC���fa�<�T��"�)%���Ȅ�Beѩф�ܻ�߷�u��Cs{�&^u�X���X�OĔ̚oBT=�����͍7St���·�5��^�{iUeM".�,5SKq�_���~�$Y��u�1S����6<8r�����i��G���HvG|wh�M|L�ʘ�[ҟb,M�sxsf�=#*���2���{r��Sȁ 6���W�~Y�6�G}��#g�<�<_]�ݹ�î���N{�M:����\�����G�^A8CL���@�;���<����)�	[?Ah�:e/P�\�@����y9���ZW3O~��AL�uܭ�0mߣ�j�q鎦�}㟞`�sV�ɘs�V�4Y��&uE���Ͻ؁�t�5�߫���;�����Z��]<��ӝ�G�jE��hH��%(y�������?��*��kA��0��@TbO�ɂ�W��d����<��|��݄���M��7Z,��u��·�c�I��z�#잻ۓ�����g��u�����k�i9�;��L����KmJϭ��9�6��5��Ԫ���.7�g���Y���%)��"�Ծ�n%Q�Rɳr-zhV����p+[x��dnA�{Gr��f����X��4�7����R�YΞ���n�9<%g/$�ޓAj���P�w���-��Y�W[����������HHW�$/������!�̧�J˓��_�&?PH0���?CG�X�o���.���!�`�$��X"֤r5���"
&ԃmiF¦`���1t,�b!KF*�%���oj{���G�U(,HC��R[���/�j4�/���;!�^�c���^��f�˦�2��lH?���h[�Z���%���47 n"�c��6U�~$4��~?8�����]�'�	bD�i�P�~7ç�8�)v�ⱦ�\M�0i���rQ��J��"d�9I*�c�;lYf�V��]�w{=��*�Е!FHE�[P�-���%i�+��u_�]��CR�D^�n4t��.f���3/xY�Q�h�����({��V����<	�VQ�c9tnĶ�Yn���uڵ5��&�gȾy�ؖ�=��|V��-&ykR���rY>��$e�X�왃 ���w�?*>�M����9�	�e���BM�8:0� ���H �Y0YvOIg2��kB��=��ѡ���thm����0�(F�Q�ԍ�X�\�����D�+u�Ѱ�y�S[d����Ͽ=a��?sd$��rh1����]�:�|R�B����W�$12���X'���Ɯd4ȜQb*��HA��[[��m2�o&�Rv�Û��-Y�Й�|H�q�R|�E|��8~C�y����n��\�(�87cY��,�����Ԭ�~lF�bq%&��w�bn��I��h���7�t5� �,q$O�7�����L�޻��uJHf�y��>J�,�֗�P`@杶g��tt�4��!4!M�N���Z����U�ݗ8J}���1ą�tg��N��������I2����=%4U%�*(F�����`���E��eŷ�]�z������{_B<������~d�dT����Cﶈ>����?��?��0���?�~����d!"���~����9�~o�  �   X X �P@ �� �  t�`� � ��  m�������_!��K���ﾁ}��� �� �`     ���$��  р`p ��
 �� X � X8 m���9���VP��I$L�s��{�L �  � X0     с+� 0@    F �  �8� ��  P� �����Fo/9�s�Q�#��ZG�o}ʪ���� `@ ,  t�`@ 0 �� X      � 
 :!� h���7{��w@4@ v}�%�_4��|��������  �� X ( � �� `����p ,   �  ` �  � 
������ >K�?���) �{��     ��
 ( �@, @(�`  �  ��� �`  ���7ww� @��,A��O�?���$I	����������?'��������v!���Jzzc��	
�BBZ��HB��4!j8Ҹp�j�����vvt�\q��8㶜<qǮ<t�J��B�T�HB�P�kV!P��j�.�X�b�P�P�ӎ�q��8q⸮ݴ�ǎ�:q�N4�Çq\q��cr�{��<�/�-���a���]$�a�B<�z�c�I�$�|��[k(�*jI+� �*���Z�I��JB(���^+�p�Il8 �Q��u!Q��UD	�#k�A�Z�)��g�t�6����Ź&������/��p V���[i["|�U�TN8�'�!&Qq��g�;XgfL���흳�� ��X��%P�ĨX�xtQq��ҽ����N�-��S�m!����iX�Q�f��8a�,`�����g	�>K.dC���v�A�L��e�~xm 4�)�����H�MR	�Ozý�-n�xH�t�����h�V�͕�}���kJfi�0�og���!��&�䩸�4��,�YefL�9AĥL ��"yσ4��1>�CQ.ݒ�+�����ֵ��Y�UNfL����a�ŘQT 9�33{ֵ�seQUC��37�kXw1fUUUS��37�k]��Ś
*�̙���ZϜ�Fh�*!�B~F~F(o�ɭ�)rb��Ŗg)h�庡�V3���k��#cJ��ݙe�'`I��i�4K�d��ܥ.e�\����=�yh(ډoʐ�/�g;�S�yn���L�M$�h��-����sQ��t�8�4Iʩ�)��lM%x�5Z�%B�fH��Q`J�E����9Nw�L&�#�DNuG�b� Cb"a<0`�\sW����0���G��.Wݦ?�q�Z���{6Xҭ�v���`��`r������n!>���y
�I&R�Y��)�ӌHJN���1⪼x��Q��e�Q�$�Dr���a/�5��ce�I�W�i(˖���D������F��S����B+UN��U��t<�1�oơ����og���YEN��d�c*T�~�F& �M���sk����c�Uv��߇W5n�}Ev�ޣ	xҦ�]<��9\�����e��wi%:QR-3��[iIM>t�5�$�UDєh��D<4}cW��E�u)�K�x�uR���F�Xh,��CA��A����)�))�$R�B	��M�[��A�"@L-��*��#j��Ȓ�c�-8agO�2�5�l��a��u���ԡi,�l!�j��F�.���v�+5���,�'d�x�I�Mj)o35x� A�/&����E �q(�i��l�4T�UU;H�6�x�1}$��Y&\$�6B�6&�$d��cG�6��4J`�w.0	l.2,�����nC�iS���Z��a�4���4�!�4\���Y��|R�j����I-/n��*���I�%���)7��7�JL<N�bm��i���M��*�כsq�RQ�%��Ç	�'���ܧ\�UQUEVl�!
��>�a8c1ڪ��!�/�q.�՜��Ь�+�{�Y	�"�ֽT�X#ƀR�H]И�Y��3���kUW�r��!{��6l���`��A�4J;Jm-.�i0L6cUA$��xds���%&�՟"e��@�`����Ye�Y�'ٯ���M��W}϶��##�k�����M�
���h�B�"Fڲ��I	!�{��'�mO���Q��n��]uRHÅ��N�uU*b�Kﵩ	��i�w��i-�͆_IT]�p���,��*t��򵅽{��pzKؘ��'t�虊/��;����T��X���"0�u�3=��iَ��|���{��Y���@#f�4zi�����u�vաud����UDuA�&��p��$^���-+���ۑ5��>r�~L�1 �	M|���/�q�Ӭ�I�N�����WM��F�,��H�(���	  �����22큪�����<Ye�YӏYTfV��՚�|#I�.���0d�['�Yb(e2�Q�9WM��%TddB�\����Z<o�F[e����,�A��S�eQӱ�>u�pM'I�9�R�J6uS(�_�/f|~'��?���D�*5�Q��`��"8(�j�����U~c�g�~Vqq��;�=�ppO���d ࣀ�
;0���0k�k�G�G����j`�c��a�,k�����p~�a�pQ�O�?�;4C���?\���~�Y�c�|aM}$�6N1|^E��`�Lb�!�I'L'Ż2:!����ࣀ�8x�ՇGgI�I'O���,ё�+$�0����������~���Lh�ջ��&�1�upc��Xf<��,^�Jn1�_sAJ$&�r�Y$rAn<4(�dꄐNn9��a$J�J+N�I�B�O��{6�a�.+��ARƶ�Ax���Qc��y���ϑgqH-=��H���XaE��G=%��6 ��/X��#��\�,�F�`�k���n��/?�K�O�M�w�T-���s��z{��j��2�ڹ�����Z�>ɑ��̼��z��G��̼��z��G-rff�7��Xg�8X�X%ծa��Ye�DE�è��(�B�(7YPL$��M�!d?��BPPPZ
₢��� B�>IY�H�1�u����<�I������w�?i�3^h�,��K��TBW�]�G�ʗA�M�+����)�j�2���I@�H5M�?0�n"�A�1� 2y)	Z-O��.̤���^):G,Ħ�-�	uk�Ye�}�?s�����yQh����{�r\��*ؙ0\���"����藬8�M�`����?D6�)�9G"��r�����1nf^�O��0'bs�C�Ӎ�m�H���Ł�R�%��%x�q�Ā�E)B�%�P���1�t��I��\]��m"RW���uab%կ��<Ye�Y9��#����2���Dckf�F&~������&�x��J@�H�|x��2ה���n�Ӽ��߲��K3��TsNk����5<��w� @��O6���Ԕ�QUR�1�o>������Gi�M�x�v�8��7 ���)YORvO%5 �� H��uġ�X6�rw=C�C�c��=X���L�!!CȦ�i�q�D�D<\���O�$�7�Ɠ� \C�$Q��E�P���g�H�z�iaw5��r⺑6�~Ql�*~O�ّ3˓r��)ɥ�LU���oe�Ye��n���)�Y{�#LH��� ��&i�iJv'6��� �% d<��$��#�D��,�.���XD�16�M1��`�R)����Cg�I�]�������Mi�,�4�bF:�"l�R�%���B��L$�=�q��F��D�LI*ZD�>#%)�8O��d�d<Y
 �C��Ye�{�?1B%��Đ����\ԒB�2���"4���)���"��?0~ u�ZG�D�3M{1΍���#�L�����1;�S)t�G4B�����_Yd.�qn7j��m����d�Q�o�����u��:�� �@[D���]_I�P��h��(��WIct{P���[���ST�W����@(��
K����Ye�Xm0�u��� j�	?��$����4��i��'���!ؔ0p�O��_���%m�Kj���%���6�z�	^$$^�FJ��z�7� RD�!�2I�%�@��3�b�'s$�4� q�i ���f�ŏ�F:z�4�i�Lt<a���<�SI3�!��� ��~[{���y��ӯm��%��7�oO)�;׽�J�͍'��
'gm���B׉���B�A����$��c�>q���w�\��xÌV)��i���D�!��� �owדI��1������L�.�[�<��ZeO��"���v����2��)i߳`V����k����B��9p��W37�V+9��g0�VKMz>H�s�չ�Y�q�Ic����LV��C��a�8�!q2�xTV��?�iL>L< //�Q0������F�t��>Hx�ɴэ���`}�ӡ.�d$��]������?Q^K~H��_US*�L�&�N���h�韤��������(i��1�lcu�c�����iY�=F����>����ffc��}c�;��"�r�CG��t	H�Z�� �|$M!e�QAĂi;�I1}JL���98H��ԧI�rH�L5�9���鱺�U*��:��&�g��d,H`Y����Ek�h��}d��W�U)�+��"W�;N>WwG+�CG��������MR\n�b���3fO�	��<1,W���ބ!��(	gg$�L����m��,ބv������1I�[Q���{�T¦Sj|���$��A��ä:t��>V�O��#�H�pQL%#������`�����!��k�d48;��L<���&��B
&`�`��IX'��xQ��į�	��+���	���<LÃ��x8l�ࣂ��X:M�gmp�0{�0�~'�3����	�FN�'��~>��~��ل�����ѐ����hp�X�A��G�pgpM&v2p�Nlf�!�c�G�pp�����;'�d�!H�����+��r�nFBH�����kw]·79�'���މ%)&�3�3*e݁�j���a�ߚ���a�Sp���}=1�%��I��ױk���$r���'��>����B(t[b���Y�SV� ��:���Za�j�h�B�^��^XWaB��0F��#�7#���EvT���܇�� ��Zj��FLǝ�k>�E$N!a]r\���`k7� E&t�`�R���W.V�e)�Pq\O[G.'@CV�f��/fK!��&uV`E���S5*��B���E��Fp�-vPpL9��J�j����_D�LcBJ �TO�_�$���mV2gG�8I��"��م�.���T&&5!�t��k�K�p��r/����v:jao��{;z���b��r"�L��f�b��a˒&�#	�cX�v1�"��{J�f����"�'7��T)4�k�'ҡV���N M�X�1a�l�7e�Bkt��]�t�af���9��Cۥ��xQ�d1%�E_n0��v����7�?�#��6{�����{�r�32��sz�3$�Z�f^f]�{��zC�7�{ޯe��|��I�{ޯe���'�s33Y�s���� a�@K,�0,�Bk짟7K�����\MԷ�;����5ظ�N46����Ь/�ӬH���^���ƺ]�#[ �F3b�i3Yr��Y{e��9;��e�f���33�
c����%�?&yĀkJc_%%m���@g�&h�i���N�*�0m3i����|K*&�-�ܣ�Ѥ��=��+�J��?'���>���Q��%a�n��g?N�X�t\�j�KN�<���1�91#m7�7:�##6�+M1��:z�1�h�5 �����^n���!#�	?>t�rɦ�5�Ӗ��y��<��q+tY�*�7B��?v�	���=BQA����v��-����- �6=������n|���S}�e�hk00��_ZLMGq�"��+�ggF;V���͞!Y�n.���˒p�(�F��� dBk��1p�Ľ8�rC){pR�^�:|%?'�'�w��]Qz���ҝ`3뚅)��]��6s�����/sͭ���&B�x��J��������%��r�})��)��S�6L�+$�a0�`F�m*���A<��	�1�we�u�rj8Ⱝ4�8i�QoI�\�ᬭ�N������Qz;D�5ސ��m�!rSD�vܮE�5fM5:�ڍ�7���~I�������҈Zm3�I{E���J�ڃ"�s@n�R}V��.�&(�/�P�$8O�)ѧ�´�����1�:|��]8�Ҳ����e��s��R��!�������A�Ĉu�a�t�m�,�1�t�N��K�O1�}[�-<���u�r�ƒ�"�7;<���%�8L,#�NO�i�V��md��l�	���O0�I4K,C�m(�&Nos��D��*HU˲7� �@��^|&S�r;�bL�(�u���N]'4�(�������B%�n�OJ�e�=毮]?&�oUT�T6�l��R���{>2i4�ɺ�5��b��1�n&��J4��`� ^�ESU-~944xH	e���!�k�������'��ͦ�@{RH�HBI�Ha�G�I�i퐐$�lN�m0��h�;�զ��0�e�U��a-��3� ��<�F��fY���_d���h�2A�C�T	Ԥ�2��$�t�4R^S�<��װ��W�V$h�Z����@K,�8~>,�q�u|
��:�	��Ҙ�>t�m&��r�n~g�:��-���H�or�ɗ�5a����+Vl0������&�S��PlmK:xt�ff/S��ʪ�66�^�Q8km���T���ڛ�ߓF5�P�[HJ/�]N��'F6�+��V�Q<Y�������+��X�q�{ݸ|Z�QוĤҖk�e&ν5$�B*�6ȍ��������1�G�&�dQ��o&j4����p��wYG�ܝwiI�)���|��#l����f�#�p��ի�Jٰ3�i��ԛJL��	 �`�g�NOƻ��3q�+��2�m���[�!rB�l���T�3A�RP�<�#��!o�IӺ6^Y����.�];���r3B��g�/~�ȶ(��ܐa.B��D��蜣5U����=� f�Ft�inm�ɗcBo��]�h�y-,��G��rܔ���F@��P٠<���LO�Ba��h��;^t��sT_* ��H�5wvY��N�`u+��&a#�k!���	��%�?\x�uw��im�+��<�<��9`i�_$!��m,�6�rM'[{��n��UT�(���Pp��;w�ԏ��[�,�W(�=A`O:��'�m�ԨE�ԩrɃ/�e	����q"wSRr�����p�oi8z�)���'���3R���ѱ�c�6N<O�B�G��օpHB`��(��]�]#�&������	�I�`�&�hK2,!0Q�LpDpk��Ŷ�+�S�g�v����pL:LCÂxp~g�ёQ0Q�M�8(��	�ɣ	�#�z8x�|L=�Ã���y���I���a�`���t��x?�'�ǑG�hplr�CD�L�p�N���~'MK�-d�L�	&��������r��W�ER���t8:r�)>�f'M�����h��Ǩ�����"P����H��9o�F�E�UgP_T�pIҠ�|$g��[�(Rΐ�,\҄�����>;�RA9Xd��b��#���8�c~�l�Z�lt��ps������5��$��-�w�����@n�\Qn�~B�y�(˻����� ��{�컻� ��{�������~�_��z�ܻ��{������{�˻�/y�=~���w�ww��/CA,��0���x̫�m�G�iݪ�A�w�x[��D��zT*��6�KKrk��?_�OΟ"���h��ךc���I��s e6�6�i�?m)>JJN&��1)���Ch�W�+9����	.��~�t��������|�x��I"S�Aa�aX�6����y��bn���,eM�����QUG���q,	\�>�U�:`���3��}�4��g t�INbq��m���ݏ"ŏM���:�h)��Ty<��4R$l���d%��E���ɐ:�H�4�v7?O����aٷ�±Zl�;PG���^���T�"��P���{�?�N��������ȱ��a��Y�JۻDpTb�����kY �X�l��ě��Sf� �*����Nd��M>L�)K~KK �a�%���:r�GI��O'�C�O��⑤�6�'�!$��y$c�q�0���	�˴��@}��++��T����2�c��cL��	��P�ɔ۞�6h�j±Zl�<Uy����"%F�J����q�
t��ѹ"oiȥ��S��Pq���ɤ� �|d{�$$�O4�jRe4�O@2��	6�L5NZ�m-��`a��*g�M$�am����@��	f�,���=����|�5���gp�)7����M�$*Q\΀�.%����EB��M�C��d���#/<Eb��Z���r���E�q��{��H���)-ˢi�Y�d�[ii����Y�\���˃�q,m?5&�XV+��Zz���u��4����[h�!n�7z:r����$�*m�R�O�m�),֑���&�Z>]�v�%��,�E?Qڴ����L�׉I���_�!U��}��|�Lm�i L��]]urȚM&��&���9'��T��%�a�H�}���D$ao9�-:�LOc�4z�XV+��Zt������['n��,�mJ`���N�m��p�X�����Ѹ�I|/�)�.��n,�q0�X��1�rN�z�#u�K��s�c��P�u5���6��$�i�48xgR���ƒ!I���6�M��&�'ҪQ��#8�C��R2a2|�I�%J�"�Pg.�0~ɚ��d�%)@��JA�g,x,�9jL�g�Q3(�Rx�k���	�BY�O��>�J�&%�hB'^�䄄�q6��$�!�0p��9ph����4�S,`p:0�ϮUSTXJ`��>JM�<>�����Zi.�b����C��$0ٺ��(�0W����W(�7Pdjm:���5���g��f�+
�xm�lc��o�����4� p�d���i��u)'>>�9%!��},�8!p�wx��i8�ٳ��q�I	ָ�8�<���^�B-6�\��Y	&���f}�h�q(SeI�ٕ2卟����aX�M��c����5Y����5ɰND�'�֘R��$��x���,h��@ �1tj�T�n�JzZp�P<y<a7�HP6�,���S:�4�-N�2T��D�@x��8�n�J&��/�mL4M�����$W��"xQ�
><AH5�Q?
�fL�a	�l�l`�;\!�c�0L.�d:d[dQlʋ��
8!�	_
?�¯����SƋ/�~���&��;�0�p�W�tȼd|H8(�R�pQ��&&/�K�0��>�����~'ME��88t�|L<L_E����0�>���h�hplr�A���'G�?��x�4O�g���/����M�c��`&�ᄆ���yr%��_�B8����
>
��j
�*��m,	���m����LaI�����&�f�D	R���_`,���-�3�d�H�5�M�KA�#AI��[���i�T��	�u�_{������Խp0s�DV��_�~�Z|{�Н���nv`�#�����8����7�F!i渮HJ���H�D�R�+:E�p�y��$|�8�Z����x��f$d��H6vW�r�;\�$��K��$f�RK1H���e�m��BF�c��V�X􈱁g��I�V=jF�%"d�T��)j��3囬a�̚k��"'
��[�~p�IR�*<ܨ7c[�ٻ�	qƁPܶ�����{�c�0�A�.����X�'k,2\�uR2�z�ϭ�bo&�J,٘N�S��m�*�"�.K	^���W� �R�mV�=sݵ��z=�$�,�kL���1氛�쎀"��P�%f��N�;	��`�*����,ъ��sX/s�v��uN�U���y�Ϳw�wv/y�=~���w�ww��?G������.������������.��b��333{�y�a��u������s�f.v�0� $E�B�]����%lj�L��]tKef���t��A�U��v�.B`ͩ���;\lbf���ǆ�@�A�cc%����=���D)�jَG'�@�{����:�L�룒�6H�I��4͒I'�M'r������}$be�;p�u�%^�p0�N0N�M�:��n8U�o{���U��iD�j���^4��޻��w�jMI{b�*��2��ǔ~�����i��Ξ8>�Iď0�4���`�XV+�z�c�ӫ3X{d��+��Җ�NKKEi7��m����4k��đ�=M�|��{�%_&[MS-���Ӻh�ML`ܣC��>��y�MN�����ӓ�c1.y�ʳs�9f��$�Re0�5��V��S��Z}�BG�?p�(,����d(h� �
��O�M�q�&�����>�O&Si���L-8��q~�d9\�+t�(J��݃e�[֡�*K��5�5���Fʇ�C���e�-4��,�C����1�.��p�L�NPӴȘ�x�A�i��Jq�׎�҃!��
(�B� �Ôq��q�B��	'
�q<v}	�����e�XM$�zz�p��XD��U���y=�y���e0�uĳ#ZS�	oR�I������ oI:�,/�K`�܄�
�7UP�d*D�]1���)����?I&����p1��m0�>į�v������o1�Z~��`�u��gp�B��҄_�S��k������V��ڄ��Gssk/l��m�J�c�=��h��kHbݝ�lC����`��a>BHMӕ�N�1(����v��Ŕ)�'�x��I�:�Ol-0����]��@S���+𻲵�b]bœA��qi\�y�I!$�B�U
����{�G���+j�t�c��Cu���rd<��D&SKrb��NoI��~�`�C����ӧ.%���Ԗ؛Jl>`�.�.{�햄v\�����qa���������B}�J�
�N��AK7�Ŏ��Z����c�GF���hD�!p��#s��`������%&ZJ_�)��t�a��{:I!�)+��G=�}*ꪪ�d [�p�.#����e�s��������Zpn���RC)�<h4�4j2&�-��$���i:� n�$d!����N!���+��v�c������2�+}ݼ!���s����o������N��R�]���#�d�ҨN��x�0H��cY����I����
<�����a>��7UT�g�<%�
G��nz�]˺�|��{�u2�JH�kfm<�&Sa�UN����!���	㨜}�hG��ß��N�FQ��Q�Pa�E[��`�@����,9��x�9Y��,~I'{.��k-��&,�n-"i>7�]�_�8��:~u/몫~$t�闁��S�yòvz}�BxI��4��Z}�	2B0�����×��m�cO��t|f��^���u ��H���3��M�cm��#��96P�+�V>Ut~o���՝ёʉ�	[ �x�y�$�<�4�K+	f�f$p:b^=ac�s�RW��@��$"m4��Yg�a�j#r���7Z�n\���~���3�X_Ē�ZĦ�����\Wj�ҫ�J���5�F�Q����Q�?
'�U�G�Ä0�`��[0�L!�`�pO	��dFpvB`����~>"��#���'������'�=>!�`����`�a�Q�L'F
8(�5�X6a0�p�2>&���0�0tz;>/�#�v.&G	�����0�>0��&��	�0lr�C�����:=4N��	��Ȧ�&��-d0����
8Lp�~r~y�o��h�������a��v��~Do�㞫��{AI�r�n���Sc3ڤ����~E�p�TXF�,�����.ޘC������{s4�|R$�)�%xE:9�=�:0��[���Ѥ
�sw�5�֟��G�d�ˇl�/3<���{�w��o���{����s�îfff����1r��ffo{�y�38�ffo{�y�38�ffo{�y�3``a�A0D���?�E����G�gV��L�-c%���O�><�
p��;O��T�%.��BtB��'{'2�8��z�K1&0K�MݔL�O:m:۶&�>N�BݟH�T��R�I�iV�X����&�6a+>�B�ʢ��Ǔ�Q�Q�Q����t���!��9���إf�f��hj ʫ�#�;Τ�TT�A�R�ݍ���(��5Wf�A��ɫ���ܫ� �$���Q�UQ��l��m08r��JOc���i�S�䰳�C�8��z�q�>볩��5i�O%8px���yaQ�|�7��cګ*�o�MAˏ�[
0�J|���"�,�Md���R	aPDKA�>0��n�`��zZ��b�^�Q{&���q���e�KHK[�I`��T
�-	iUR�'��̞�!��4�������)&��Ty�*�����<���G�:�Ra��ͧ�iO�i�S֘��eQE��Ŕb�E�\�r5���i):H��R�İ� �!���mc�]t�=I	V�G<�a��UH��i�<���i��D����a�Ғ����$��r'
=:�>O�m�Zw"�o[�Y�JԤѥL%���*��(�F&�4Y�҃II^�{a��1�$�T~��A���xD�L:h޷�����3�����t�m8����ݖ��롃k7r]ԫ/	>H�r��u)2����ʒI�U���A�q�ͱeYA׏�O�_����F}27?Nse�^�D���Uc�W�}�ۧ�FUV�d
�miBa@ԣ�H���q��k(�K,-Z�\��F��Z��Pj���r�$+�<
�d�vٛZ���'�H{I�3�M&SC��j�ɻ!$%����ii��A�[I�ϡy07[�d�폤HVU]���uסȳR�LR�W��x�����[�"�H��)	�S(�v91��F�"Wǹ��<�K0�V�uKgzw��e���+�u����S6�y�d��d��h��W[a[Ú7�Ln���'�３t�����Zp�a6�Z9M4���	�?vIN�Iڄ���	�\�8\x}$�P�e0�� w���WX��r��nˢ��[ǩ��L�ك��y�}ʬ���Wjګ*�6.c�}�ܐ�D�{�p��gB]WT��kzM����6�TUJr��	��1��!�1��4Pn�В�!�<�ry��"Dj5���I��5���7��� qɂIG�\:O	�2^��w}y,օ	"ᑖ�BI�>������ɰ�e��(y!��&Ja��X�� �6�e�H�Z9Gd��{	����H}ǩcGq2Z�F�%$M'>M�~Hp��B|"C���qs!��[�^,�*�_�88�!�x��
�����U!�/yk"�`�d7+�M���V�jYJ��7�VX�zt5�Q~�����ģ�u23���Y!��	�%o���8�ƪ�6�K���*�����;��!݈�� h=FU��W�u�Z_���G�
?�O�Q>?F��ׅ
>k�&���
��#�k�#�����66~!��`�=0���8;�Z�����
8*���t���H�Gᯉ�?&�����W����	��xN����E�	���8�����L�&��Eæ����0|�>/�N�����a�`�p�0����*<&��	�0lr�&x<,�&�#�t�]CC�c�10��<0��L��l�D�|��*���6�R�1Jly9N����m�q���[��mV6#P�X�N����h^h�4kFh�g����[��p0e�:+�,�TĲ�������,�cl	�<r�@�񅴊�j�P�dz�����(�f-.al)���Wl��CUG��En��b���%�rØn�k�:i$�XF%I�ڈ�lR1FT�^7^	 㥈C���Ϟ�����!bC+n��N �9P.�"*p5���Y^(&Ǵ��s�Ph�:��
^��S:�3�/u��/n�D����h-��'���]'l�[�^�oK���u
�h��<U�4ya�+�b͐�ޖw��qf���^|����9nF��e%�,�r�w�Ν�E��	^6�!���5���X�_	��,
���XU1���/�Y�o7��b�͈E���Xo;����ǲ2�S�]�6ޮ�9y�}��}�0�.q�������f.q�������f.q���kZ��ž�{��������n���{�UU~�����K���0D��3�_%������An�0���Q;�f�a�l��̌*ӥ����i[o��1�Y�GP|������$���m�]ݰ�Z�.���5����*a�u�3��!��=!9�լ�<��,�8kŶ��#'S���'�;�QI�>}\���	X�N�l[OY�`i����c|tRZy,8�3�,Ӳ��
 &���/K~Ec��7!�v�'�%�/3*�����T�6MQ����u S��䁿���G���h�en���M�Hj۶۹wriA��Q��i,!a}�t�y0Pq)�Zi�Px93�9*��%G6z�q_*�ګn����m�Oǟ}Bh8YI�&��
�%%��}R9C'3!)��3�+/�s׻�;a4�R�Fn�Q{�(�||�0�B3T~�c�Q���r2OY�/C	K�������F�x��ڕ�|��MkP��K�[C��-��5Z����Śa'"j	�K�&]%&��U�Tn��shHHv��O'��#��(����n�a��ު��UWM&Ё���?:JWL������3˷)Kx�Ak�]omG�`ٵ+�>c�1�j��ҕ"���F��+����Ln�� J�Chå�;jk�\P�����R��j65��)�YI�Ұ9cKc3�ߓ��C��S�B�ڗL�H������="D�>$�,��C�fZ{�{�HZW۰��i4�݅K��"s���HHO����NzZ[I>r`�ϳM�H\�B7uP����<���"̎I�gJWJtǬc�*[�kI�2��i<�N��J5�Y�Д�HZo;k�HM-�Bv	�|�-6u4���d��KMh�s�~�O��ܗB۸,*CO(�yHO�i�o2�e�R�M�%�j�����I��mJ�O�|���Y�>��W�9��b,VBF��z�ZCI�4��kE�I�o�0t���W�508���!�_~i����r�q�0y>i>O%'~>�J�*���R�|�7�<�)8A�| ���HBT�oq�DM\�p����3�J;Fí$;��.�7�a�MtH]�X�3&��*쪕��hӤ�Ƥ�uv�`��O��O��صVU�,��,b��1$<�M�R��6�)bw�j�7�I���YV���i��Gd!d؇�aC�]���$�-:��F,i��a� T��k��@G��lyFX��d�gP�]5�ue�7%將j��1�iv�\p�v�;~�s���VR�B������`�'STy:�9�0�-7G~pྒ���b�o_�&�'�zSJ��nYq���ka�n~K����wy{֖���9E��:ل�y�)�����B Cd�p���4D#AdQ�U�Ѫ/h��L���e(��ƒ[�����b����$���q6�.Ϻ�Oo�#U�+�O��v���۬��`f���L�G�t�&@�r��������>O��}>�M:6|q�_�OOOO�0<�ǌ6a�`��~t��q��Ç<;;;;|�+��>x����:^8���W8�q8q�㍸���x�\b�W!�U!j�j�b�.�:h�N1\8p�ºtӧ�q�j�q��Ç�8�Lq�fOdճw��m�W��q&�kg�����h��9�.��{w	ëa���׆Y������FC؄�e�Md_~y�^���t�U[ʑ^�A!}����|[&u��|!�K��=�߶�����9��gx���h��叓���s�~����7^^��ꪪ�y{�ח��z����^�u��{ު������y{��������7^^��ꪪ�yf.��&&a!w�^;�4�8Lx�g06I!i��ͦi�>�|s]�Pqe���L�a���ct����vhTI�P�]��$		<i���2���m��I)a��O��Y�N�N��t��6Q�)�PŨ;M���՜2Q~�j~�����EG�^K\��r5����m��������'R�?&D��ӣg;�Hg��,H��0=�8�ipA�C<@�8!���IJ��j���i���<����ˮN K˦��0��ŷSfͮn�jQ�x�yԡн�#6�Fʒk�R١v	�6�^(G�:����8v\�X��[5l��jE%�fD%$�kR�r�L9CW�Ѻ5�ӕ���q�XM_!0�&�p�L%�Om�d�y8�M��7�ξre(�CM�y��7��%�V~�bk���J���e!��bӽ���J���ظ+`� &�D���9�^v�n]���F���i�v�皕�e����<�Դ��sV��2R`�!1��e$\`��;��	�	f��������zt��5qumش�j�&��i��Vġ�S�=08l���:CB�#c[
��j�h�Q��m�n��i
L�P��m&
٘�����q�b��3,������=���'I$4��gP/&S%�Y��$��N���� tx�ʔ~ pDK '�"x�HB�w���cs9�p�d�8�l��>��{Y4{��>�a�e\��Gq�8�=w~����6`�2�j2�4�N8/�ķ&yI�I�k�T���RH�7��f�U]��>UW�x�0s��X����^�t_
U�\ͷ3H5�����m�ib��\p�2x�zY��76�K �f��k{�Xk��H�\@���f�,��bg��T�̕U[m4�jq4��0�8�.HO&+�%���Q�i4�0���~�g���>��i\�������|-U�E�5��	l�S+��D���tr�6"Y�DN���g����W����I�éI���RKMu��0��FӦ�[O��B±B�OA�wSuI^���&�oe�{w�7�eԶj�Q���U��+�Q�T#G�J��d�a���Љ�!�6CBI�o�#
&�f�YZ��J�X7�B�a8����z��-����hI�A,�����DT�����1x`D:q/�|�Mi'�ɬ=��a9繾z2a5N�q0�쐒+��y_4Qd6B<"&J<QEo`���M�Զ�;bq0��Ƹq�i�Է���QWu��c�UW�Yn��JN7!$�����6�Ő���5!&�;��h���)1���	�0G��B�1x�;���:;><|T�����j�BBB����HB��]Z���p�Ϗ���+�ӳ������_[�o�|�8�]8Ҹp�pB�B���B�,B�Z��\T�!ZՈHZ��Z��X��]\q�8Ҹp�Ê��N�v��4�G�8p�����zߚ�{��@N����+)D
z��$\m�ٝ};���BƦ?DL��I��7Z�v�|�ϔ����n�w۾�t����e��������LB�\���g%��Ͳ��CL]���ǘI�|���HR��&��o���-����:�	�wb�u{(y�JB��0�A�1f�agmפvGf��'���佘d^��Z��o1�ٗ0��J]��kp�\�6n{Y"���{Z�c�}&�. �I�`�E�PC�(ڎ�(h8�Ǩ��,�|WQ�Bt(Ir���:*��;0�_v1Vlp��	�i�,���Mz-�fF�rPj)S�;a��,�)�`�(1tLP�È"�� ��EalA`�%���e{e��N�>F�H�c�YB�-�»W��S}�<t��a�KJw����Ƒk�����z�z݈4�*��j4"��L�ٍ���,��,BI��QV<�#e�������ԓd�Yu8�m����R>3M�P�e8%�c�~?/�%��:�D�j�3��ͪ�����o�^��ꪪ�yf-ᙙ�ֵ���xfff��k;�b����kZ�ᘷ�ffkZֳ�f.�`�!�"a![�Z@g����c-�S�"M�XnXŶ	�m�0^�r����KA-�5�SK̒�vY�M��//m�ǰF�c��"��>��A7~���||�y((�fHB��8��NHe-�}�ڒ��-#��u"Y~$f�)-�Q�$�L��J�c�	�9�Bm�0˺�F�������T�{�;+�a����8�1�[�w֮�j�`%%��I��&]��%%&�h��IM��I�.X��r����%'�ɡ�k,�v��YWx�(p��K���%����a�yE;ɒ�	Z��0��&ā��B��+1i�Y�M�S7��S��c�zH���l��j���|8��jBT�$�����I�BL�<�K^����|�q[L��U'����:�s��?Eב�}�ٳ�c�Uv��(�%ަ0���
�<�<Smpm���M�g�2J%^*ʌ7��6�HD����ؖ�N�g�/�^�:R�]�(�s�0�� o4|p���<"'�8Bu��U��57 k� �ݻ���eI'ĝ(�r$���[��`�;VQ��.g�_�������R����
8,S�׮�����7c�k�N:J�[%j�-Ȭ`�mȱ���Ϛ���i�rJ��Zy>8�K��M/4�}�'�8ID�ϵʒ�
�M�H�r���!��(��������d�7?3�q���G�a��D�!	\���rkZ����
wGa�S��'��Z-:�!�41>O��UѪ>��n��,_����$��)*MK}��`���K=ư�%4�QA5Gh�H�d�p��:B�U�Hյ--(�xlh���]���S,|I!L=?T�WdǒIר�7�7*�[�SFQ��c��R��"FHP����P�����Q9t�M&�U��|����}ω��ʊ(<2�N��i��Fӹp�ChDM��C��^�Ի��^|sROH�%��ї�N&��a��]b$�,�(Klѩe�[0;H����
m�s�-"n߾2o0�����4�y�$���m2��bV��-��ֺo.\�]z�u�~S��6"'HaC=M|mڒ��0�����4��E���`-}i��Vl����Qh�	צ<��{��<'��ʆSdeN�1"�?HLI?�e�ʴ%h�Y�˜���Wy/-<v<O%%���[���Re,�q3���ú2�O6�	Ik���'�&�;����,�Wf$����f0V(�K"��)���-�c�G����w;V0����B��.���>
�4h���*Uv\l�$�G�+��D���9�q(���ȓ�ҏ�'gyx����$!wR���4�U;��$�I�Aߊ�X!Q*4+!�D�R۵Ք�i:�ӜPHT��!��l�d�����|�ã���
zzcӇ������1qP��HZ�(�Ӎ+�8p���������a�ưp�a���'������8ێ6�v��=mƕ�\]B�j�!j�j�-BՋ��:iƜb�p�ۇ۶�����N:iƜc�Ç8�=4��C�H��+K9 y�D>D���8d,v�jB��{Q�L���>��F�n!�ީ��{0S��n܍,��=�Yj�E�6��C�g�nړ����hP��Q����ր��̖��b�+�j.F�Z?�~8}��I;|��������UU��~^�y���j������?{��UW��y{������U{�g���?{��UW��a�4@�aJҮ®$L��;UR�F�8��c&�i�\�N���᭳s�i�f+`m-�O�ïɂ���$�)��}v���d�u'��Lh�3RUJc�'�����1⪾c�1�#!�HQ�{Ld�'�:ϢC���i�D�Ƶ��h����U�6�R]�I��%|q0�HH�H|[�53i�i��v���!��Rd���[$-�T����>���� @��D��B`��#�����{\[�Ѳ�G��bn��׹��r/ZRc�yF�5��]�A��u"�`bK��b��.:�H���٤e"�Ky��x�o'yy<4d9��i�g11�siި��.�b�`���6SE�&���gRFKs��{�dRTx�!Ĵ�}~0�MvI$�i��iy������$���Q��<�#�	.�9�{�qݓP��k¡'����~���#q�5�I�G�a����!v�>/_K�x+�O��"a41v^��&M��9;R����M���H���u�7�6VPc�����%���VF���R���vm8p�$ހ�)JL%�z7$B,��#��x�)�0ƕU��:�b���Q(����Sx�ݟu��Bm6�6��R�=^(�W�,���_�H;���\l���UHJ���$6�)i�0v��D�δ�2���c�:a�+FQ�w���Q��w��N�a�U�0��|��] ����O���3��
��/�<(J�I�܌	\���{ڦ�L��D=�U^���:�/���&�Yʕ	U]#��
N�̢���"e+X0�N���p��d��n�2���#&i�ƞGR�a�"'�8B��7���!�K���x"b%�?��Fq�Ry�J�rS����O7(�oY׬n1�d��[k�u9�
CG	�X4�N6�2��1ؒ�aӳp��i��[>��5ww���vb��Fi$~pӃi��jB��&_Rt��p�'�7P>����RG�7�~��HL�ry��>O�`�%�ˌ�;lj�v;g�����ni����2l��a��U�c����^�ɨ�V5��V��.��E�j�5ƔS�LQՆ���$�[Q٤�L������1�0UV1uUnV1��^&������ƓI�ܞ��I�Ne4e)4�6;�
	bزr5=0�1�UxǬQF�Dq�J�P��H4E�
�t_	l���]9�k���$�a�>�����s]�oZo�*а6�4��v~R3{�~n6��e�6�y�Ө�h6u4�2�qr�UQU*���L&�����f���UW�x�1�mַ%���[��&��e	���V�-i7E�n������F�H�!ZIG�q"2�?n���D�k!�]����*���*���Q�a6�^c5R���e��I4U�N&�:�&�#P��L��k����������A�$�	�~�$�I$��UTJ(���g�����?�O��l�B"(���-@`�������gE��*�Z��G� �XOl�ED�X)�PR)
E!H�B�����T�ARQ*K	RX����Ċ,"�"(�(�b2HQRJ)%AE�T�HQd�I(��5��Ԉ��(�"��(��,��Ȋ,���(���(�%EDQd�E�%	E!E�TE�d
,%0�`�peR�YE�5�#R�Z,Qh�EJ,Qh�a�#%(�,Qh��(�E�RME�eQEQe�T�����(��J(��5F�<mXʳ�d���ꑨ��,Qh�E��QEXeHȢ�,Qe(�X�ЩF)(��(���,����1H�,Qb�YE�,��QR�Z*Z�QeQe(��X��,Qe(��YE�Ib�(��(�E�X��,Qe!R�(QB�Qb�YEYE�X��Qb�(�I(��Qb��YEYE����E�,Qe(��YE�YI,QeX��Qb�(�E���Qe(YEJ,Qe)%�QE�X��,QeQe)%�T��,��,Qe(��)%�Xԣ�X��,T����T��X�eK)R�K*YRʖT��YB�,��(�X�e$��TP�Qe(YI,QeQb�(�E�X��,Q�&RK(�E�T��(�E�,��Ib�X��Qe(�R�K�H1�1 �`�j%�,T�R�(��YK��(�)aK)b�R�R�,Q,��X��*R�,���KK��)e,R��ZX����R�-,R�h��R�R�ZZ,Q,���QKE��*�R�J��QJ��Y)b�(�JT�R�X����R��E��R�K�K%J%�,��J�Y(�R�,�K�K%(����X��%��)d�R��)d��X���Y)b�)QK�R�Y)b�iib�J�X�R�--$�J��,R�,��D�K%JX���)b�JX���,���)b�JX�R��X��U,Qd��X�Q,R��)b�J�VJ�UV*E���V��b��b�U��d�d�*�UX�%X�*�V*��Z��VJ%��Rի*���V*EU��UV*�TR�V*E��U���V*�V*�V*E��U��(��dD�RE"�JE�R)%"��Q%��%�E"�J"�)H��E��$�RE"�JE�����%d��DR,�)$R)"�d%"ȊEBR*�Pb��D�e��k�b��BP�)G���~�(�������HI"�'ԕ�����_�s_�9�������'�O���������?_��_C�?�������e��ؔf�?�	'�ߧ���_�������$?��g?�l�)����? �
/��?��?TO�����}��w�������A@?�<�ɂ*���B�0Y@�����?��x~��!����HġJ_��o�0O�:~���؇���!���8�EU~����?��xI)ZZ�P�Ko�\!C�[��C���Ĥ��"o�8�4�5�5��Ѹ���?������Z�1���?������� ��H6��"�e�B 5j(��
�� ��TTLl��B����%]7���86���_�?����`�ER�UZ*��Г(�$�-R"]����?w�����~/�z����$��x?����b����������I�ZtK_������v��s�?�~�d�/�3��a�=������_����`���S!����$��C�?���u�?���D��g�����'�?�  3����Y�������鳧��#�+���0O�TO��@�_�N����*��a�:O�m4`8|I(��?�Ш�r���h�$���G�[袀)@ӣ��d\�C062���)�?MhN]���������.	ȼ�A�  �+�{��O��Dg��k��EU��i�?�E'��?���t!����������?$�U'������~��	���������?�ܑ��?��������	��*�'�R?����/�п�EU`��!�����������?�柉�0��� ? �����BWBUS��M�)f�m�m4��?���?�i����/��|��r%��I��p�A��}�DUQ4��'��Jj��~g��?���|'�c����G�����Nq"��B���J=d��#�)�O���O�?H� �)�@C��	�������?7も�~a���{��E.��ަ�O�������ȯ�C�)T�i��������w$S�		�4�p