BZh91AY&SY��>ܝ_�rq���"� ����b!�                                        �  ;�o��   D  � ,`�P     
    
         P   PϾ� ��R�$�J
�**���*�T�$�A@ %JI���()� P UQB���(��� T 
 Q_A]�焠�� oXtDb�nP�㠞�:U�p9 �A�n����s���
r�z�BB�U�*�(UQ��ڷ}q�����x��h�y{⨪��{[U���۵���6�7�Wme�ݪf��yG��@ ��)H�t�v@@2�T7Y� �@
}RJ��!(�@T T�*�D�	*� �� ;� 7`���� ��< \ ^�8���A� e�}��w�< -a��hw�
 J��� 	�=<@�>� =+�=����q}N 1�� ={�힀	��Qx -g���v��^� H Q@Τ�@�_ �AE�P��
���݃��A��9 1����/�⪋��1� =�����{�� �w���G�� p   ��B�@>�7����X z��<��� �[�/A���{ ����x �Ǘ��/��`�n��T  �)@H����QUJ�UO ������X  nJ� 2@�>�޷�)�s wx+�C���
  �sґ�W� x�� }ޕRO 	 S�2u�� ��JP��������s  
 �������PW�)T��*�J*������ ���n��t�"��t �� �L� r�P��9 ݁�
 Ax�*)T�� .�� =nE�G 2� �9 wR�N ;w��T7g@� >�     ��50�R��     L"��	)*�   ��  ��UJ�ʩ���4      i�U �*   0�0I�D��U@  �� E&F�)=4d�FF�4)�=L�P�e=C�S����[� 8L�/>i�|)7��z�u�Ȩ��܀��	��E}��QxTS�
���D����
��������g��=�>�v"(����I$��'�QDWى�������*
�?g��z�����ٜ�F }lB0B�T��QF�AP�@J�EJ�
�Q
�
�k � ���Z��Z��Z��Z���+#
��@�U� + 
�B� � +
�+#k 
�Z�� ��Q���+kk��P+
�B�P�+J�B��D+
��c
�R���F�V�F��F���F1� �@+
���PkJ����# 
���T+kkk
�Z���@�+kkk
��@�@+
�B0 �+J���k�P�D�P�P�A��A�D�U� T+�U�DR�@R�F�B� B��R��D���ۀ���u�s��0/��G8����:���b���:,�:9�˃�h�8��t��@�5rc6@�9���3����{�N듡7�]٧Yӂ����r��4 �K�m'^�	���`�_�/^�3�3��&�b�Θ7UwL ���K]���8\�:�M'����S�� :�ՊK_d.�F�:C2b���Y�2'W}'d+�v��F�np���f��]��`�=}8rN�u�.���μ�V䧸dF�V��w)�v�lh���1oN�ݯh�s��D2��o�U@��������A�_3�"��Vɼ����3��!��Z,��;�s�s�1n%n#Iޘ <y6b��AA�؞Ȫ;��ݫ�����w��<89:��]�)�����#��[�m�C�l27GϟC����6w5� L�r��;�wKm�73I�d;ۗw�?L׻:`�rlM��5=M7��8@P�s��0��؃�њ5�ձ�Ӊb1ӻ&��m'��n�lk�p՜��powĸ.��'O�np8K��=�$�2�vu�^ۧ�v¤������gd����J��:UD���ڶ	�hf5�S�˶����m�p�'vu�;	xF���ze:g�fߦX%������5a�ز,��g��G�2�i,"s�>����ݰt�Q�4h��7P�-���{X�q���6Oր�G��%�x�ܽA�ne�VtNh��;��w�\h����^ ��d��L#D�����akv^���-�sA�Bg7�xͬ��
���)��ؔ�'�O`�V]*�l��Lahо�
q�=A���@��Նd���ud�����	yZ�z�����[���n�˖T��YΔ��4�d���N��c����f)5tVx35��Z��q��������S�svG'�Y��X���w2k�y�#D䝓ju�{���P�q�j���V��ި9³�y���崽�"=÷8$lfһ���;�ièvC���uN�:��m�ѻ����ƞW�:��{�͕�p$5m{��	���x�8��NF��������z8�ɵ�ʴ��:`#-���^!�4��8`O�Y�%gN)�%�!ObK�R�7�������]�,.��I���D�N��L}�W2���^d1AT#����� `�1�۬+�VI�%X{i�AU.fɳQnr��Y8Nn��c�X/�2�u���C��f�{��"c"0s��Ț1ø��X�&EV0�FY�c-��6׵ˏp3���Ց������B�Chچ����a�X��kjV�,X� �q�a����9HΪ0�>	;gL`�)��BmR*w�jT�yMa��M.]�Qv��`�y��Ҿ�fMkwm�N��)�P]�Պ�w�B��#Ż�'���2��;�Fܻ��巰[��7m�]�kj�����ת�Q���qt���h�i�r�0�[d�M)-���b�c5��6�^��y�	&`p�Ճ��"���ؤ�w��&L">�����J��ɧO|2]��w3��2r�{�#Nhݐ����^�δ_D*8�Ƶ��/a=x�[����`$]��w:�_b=(�80��;z� 69�VX+����]���;~\onԪn*5�u�%����;I��T�F��R�xt����p|��]�s��������v'�K!4c��hou��H�ӵ pI��s�v�orc�Y�Y+M�c�󧳏9�N�\Ճy�zd0a T!f[�{��]/�����]���ǝ{�j��H����&=�b9�D����0<Q3��ſ!U}�c�ѐ��#ײ)�*�܃��C_g>�س�7�m�h"��Sr�r���Olyehh�{�eٺ���u��>��f�(�3�M�����983�i�uw��<�<�UH���29S��>_K2� �i`9����ۑ��uD;���v�}F�����HA�:��L�������5��V��b}��tY��tG�c�c����R2�ohY)%���gueoLTK)�m㯀��x��b����l�5��0�j�Y���~�r97�K��7��;9�kvG;eX��j��b��s�^cDW�k>%L�l��S�ɫ�uzp-�B�6�L�wԩ��q�
c�J��9��r���Q���9����1
���wY��#%��;�����=�2��bWE��G;S=\���0����h�bڹ�:���9�n�7���xBI��t�ӎ��Q�LΥM�3���۲�ݏ�\JɆ]Z󺑹�8٣���I!�̑ �w��Qp�;:����>�;)��{	= 	+�81�)��9���&����JR�Q:��6X"�ܫ����gRx���-wq��Ǭv��X������7jƲN=u�����4csE�P��R��eO7r3�f���H�6-NQJ��Y�sy����1�廨��Q�km�es�8XUqy:�j��Zӑ�庁��'���Vi]�\1s����P�H��h����e͝>G~��B�on'&��y)��Aր.]�Ɇa*�f�a�&��6C��K����S�K�R9[�P�'
*?MkɈ��y��_gN��|�ѻ��gh�r��aql��p�vt�#T�ܤ�^���8��.���dP�קe�wN�qQ��*]^��e�wi��D����� ����נ��$�Y�p�E��-����Z�f�HQ*�Jtѫ{{� )�;r��S���s��XvӦ�M�i��֞��,����`�Pw�����[�.�u\���` ]��R����DlN��حڇD�B���Ӊrn��9�����7��y�Pk��ģ�i2�v��;6$�B�e�.���8R�sre��4�kZ�>�r6�<��;����/:Zo#�I��EBU�c�Vr��&�|k;����9��.���s�ˢt�W��R N�ئ�׺����yV ��[�ڐcfi��_��M�7�S�f�d�u`�;���E�Z�%M�n���j�U�s�(DȎi�u\��F��nk��G��Gu#ɓ�ғ������C�t��n�:.���w�=���DK�,��2�X�y��kŽٮp�t��y�[�.͇gn�s�Ig)�1�۳�| ��E�+;&��<'~���"��k�Mrd]"�8�Zn�	 ��VUH��n�w�xΘ�˸�+�$^�g�ܛ�Y�Ǭ�к��Ö��ƙ;��]�DMp}�N��ho�����\�Uc�u��}�;�$�d�5��d3��3qk+q��gw�we�۫9��O���� nnmYD�뛎�W&��`ہ�a��k4i�΄��*e�����5����	��qK��(�SGs�dgk�lƐ�a-ͯ[b'�7xUa+e�ذ"��<;���b��X{p�-�9�j{��aKL�w'�i����v❻��E�3���h�n^���Ge����").%c���$Ws�~QT��s�YK�}�ީ�Fw�OY�ʷ��	ٗg'��q��&ժ�M�ΫD,������\2���C����ߥ�wGۺ�T�{9L�\]mR�ڴ�ܵ��#�Z5		�F�R�;�lY�;���la�S���s�p<e/��n@��I$�k��N��"�L}IA��M-�Z�"���k�1��� �;7��)b�%��B�nL�vbK{!{�$p/x�˚ׄ%�\�s�AHtsr�� �E�)غKhh;X3j�p���9�J�w�#.�X%��A�۱/��^lU�m5��jow���+r �^���	ܚ5��'��$c����:��6�]��u`�!ǿ��{��-�k��J`�W9�x!z���z[/i�!N���]�r�Q�r5�ݯ[9��g����2m�7���&���Q-[���][q�;�.8�����<��P3]sP���6�p��/:̖a�&�㹫F�-�ɰ'UY9�dzn�G+�NJ���8�X{�J/u��7L8]g��]Ҧ�Lŷ��r#^�ܺM��4�H����P'O˝�m���v���WL���WwM|�Ϡ��Ͱ�+�Y�Lr��x�@Dö���z�5t5���Y2�۷vw�\xq�볦KS>;7�%����C�F��)Y�ѪQ5�z�T��u�9p�oD7���Uv,�ل����Z�F�'��c����(�%�U9 <zߍHZC,��QѴ��k;���5������NoG�N���VIp�:`�DB�]��h�<�:��
-5cck۽K��z��8�rws0ܦ�ۅ��>V[��Ri�Wiic�Px�ц��V�o�A��킦B!o,�o;Ͱ����͘�B �Zu񳃗F�D��qf�Y�����Aw^�^q�Y�u�v�J(���G�(;p����)4�wik85h�W��;9��]��=0����S�,�����2�)���!�ň3ȗ�q6N�`'�YwGf���A�;��6���ӧ =��j:2����|��^+8��[��OӧAʜEO���Q#��L=�v<1m��ӎҞ�U�RǛ�'. ���bΤ���A��G���Y6#���ӷ.�3p��S,0�/�]w��Χv7�q�ᵓ�������[���vH��: L�o���j�
�c5�	�$4H�W	�Wy� ���y�5�4�}GVlZ�y�*�F�>�T�arj�,lds"�Gf� ��f��p�H�]V6\ -����U��� �#t�i�޸m�gH�6K�)C�1���-˖E�#F$&O�|3�:8�]���x|����;�C�fC�N/Y1���w�c[��NE�:dt�3�q-�9$�f���o��a*u��xr�41,�,�'v�����r�\93x�T���͋ecqӣ���v�y��BO�8�A�ȷ��먒%�̣yb�����9��T[�a \Qi����xa�boR�Vʛes�kq:Mk����Wڣ<1R��G_A�N#�\��7E�A\�SJ>�wbYX,�հV[y��שq�e�3j�i�2v�����Y�P1[�K�]q�H-�a��-�Ԭ=�
}&�C�!u�D����6��oŎY�!{3�S�����d�-\�:��z�y�Xlc�5S�4͏u���M|�7rG*m��i�<aڎ4���x��ga��.�{S`��vڎ��🠯*�sk��2�^8c������Ø^{����r����uޫ6sO#��ac6�7��p�>:��݆��>e2�܇�'Y�mJ��\�� ���(tm����.A�C�uW�؊��(i�pd��5�u.���'���� �=�o(y�l��g��ۛCu��b�����8�@����ќu����u���v�ڞq�ײxYo�"��vJ�\E�4�M�ޣN����̸�<ڴnj��)�cᜓ�z�~�w��j��=tp���1�bΧ��nCR7�Zg��]�2����PZ0�Q8�� ���s�1�VE瀅�^����[M�	��R�&�[yXA��w�weV�����u�� �ɠ <:$M���(�5P���������M��X0�5���sk]뛠����:�`壊�T�n]�7Mp<��T���Z�y��u.K��:n�Ƚ��=�1�{I�T��'��׫Aނ�H���$��@��w�L�Xۘ�s�Km�j`��9��m�n���E#��^Ѱn�z�*&���tH{"�wBh���o+���ގ���f�\�q�m�á�th���4�����=;�D��J��1S�ӶsX�r�.Q�kk���ü8e$�F7x���qטq��ͤa��x���5�#z-��JAsSx�ǖ��;&ӝsZ��aZF!p�Q(A0G`��)1B�L}׼�C@��bg�Y�AOγ�7̺;u�����ۮ�۳�'K�9c+�aYC3R�VO%��z�۲�;9(s���;7'n��&8��d�Ѵg-3�7<6�.�3���}Ŏ� �����r~w[Ů�OPK]�3Y1�<I�g:�lf���v�h����i�`�m�v�e�~��/�f<���B��g5�v��@Q<�h�-Ǥ��Ӌ��(yMH���*�n�x�3g�Q��7Wq|
zSO�U�����KG]ִ^����ߗq"��jº�����*�ܜ��bf�:�P����ws�7���a�'�i�¿]ID�ӳ��S�A��G	��
��r\�R���t��I��]���h���Zr��bN����R(�3rj�gDGM�i��o�:�����Q��X7�H��9ė4�Id��g(we�|f���87�坃Z��2������owor��vt}���Ł��j�����嚙j6�u���j����D9�82M�k��ɥ`] /�ĖJM��]3�>W��R�r!�\�����I���mK��Ԛv�ʻ=C{�`Ɍӣ�{��LM����#�Bg�Bg�u��h#�3d��`����������=�<�ى�ا�ٓH�OZ��f�c�#C��V�̕J�b��و�L����xi\8�e��pm���]#�W�eE���N��|�����m�V�iҔv������,�6�g=���o��t�jY�ɯx/���>_�������}=�|>���<��EU�dE$E$$@	 �b� $�H*�# ���� X
��`�
(X���� �Ȃ���H(� �%�(H�e����H
��(� "�  � "*H�Hb��� +"��X
��"�  ��"�� 	 
�
) H���������� � +bX�H �"�*�� (�2
ȢȢت�*) �6(b�
H�ȨX*!"$�X�� �b�`��� ��X2
X*� 	  $��Ȋ2,�� �	  H��b��Ƞ� ��,�"X"   H�x w{����8ߓ7���/���F)�5�!`ho��xv������6�,��^��Л��_�}����ٲ?F���ы�&�z�w���Q1�~���?n�>{H�h4OnP])�[�fm.�����w|��s�@�$��/������Ȣ� w�v�_1����/���ʀ�/�������={>�������4|���s�\gGZ�f����}ב� 4�0 �Mb��>�vۢubSh}O����u{hI�<�z��W����E���5��!��d��dOY�|�����{��X��g�d��L�Jу|7i�V�m�k�Sx���KЭ�|��.���B����|:���ى�W�^:��
M}�N�����3��<�}_�}�ot�PO�+bs�Ɏ���ޞW�:]-w���ܽI���/a�<�21� ���7W��8�ˉ���ݽ�}��"txNo������Ð����{P��PV����� �Y�M�9�X��Jv������5ɒ�ٻ��]*��|=޻�o��s�Y�7T��q�L�y���ގ�L�q�	����ܿ}ｆ�ϑ���`0�=�!��s8y�x��T�;��#<;���^��K�<{���`������j��?e��_x��9��*P	��]~X���Ɓ������^%�w��Ue����{yƨ ��%w��s#��w�yջG��g����o�wg���U݌\��}3K�n[��GV����7�{}�7:28=��JA��^/���8rN�������s�徜���ٝw`�s�ݑwo�G�/�� %��^<�ɣybKǆ�R��r���0M~���"8{z)sc~s�Iػf����������}~˷//Nݻv�۷n��v�۷n��v�۷nݻv��۶�v�۷n]�v��۷nݼ<<<<;v�۷/[�ɹ��U1-yU����B;��i띁��e.�u�x��߷���e���e�뽹�����k�	�����}{=Ƕ��pZ&��,Yô�;��:=N�;7;j�{=y`�з�H1v@�7��/{~�w=�*񉃦掯үn����'�d8w�8�]�'���orl��2�[ܷ�8`����e��K\rr�j�v�M�%�Gu�S ���G,z1ok�/@c��N�'ۼU�oq���8�\�l��)�!ib��;o{��K+�����9��_�Ӱ��O��W�zu�5���4>Ǫ�ě�,�]Y��.�7�
����׉�����3f�Y&�ʌ�~������Hߞo�G��e�yݝ����g��M�|f	wk�����
�}-~��ب��³��6{7_5�^����=g���oq�,���_�.�°,�r&��Ko�S��X[����KyR�y�<�x���]�<o}����q��E�n����� ��I,��;���\��x+I���9��e�C��Ֆ�}��,���G^pW�
��Z@]=�y����<�c�Yx������q����ټx��n��"�{��PU�E����{	y��š�ʓ�L����E�|T�f����'���t�u}���|_nH>�rN�l=���x���������I�5��OM�-#6w,������M_��˥$�O<�}.�]��.ݻv�۷nݎݻv�۷nݻv�ݻv�۷�n��۷nݻv��v�۷8v;v�ۼk�x�:�Z��Y\�/��ި�໾�?w��^I�ѓ�Wք�����
5��NRn7W)�4e�������^�\�{W�+4�a,�7��!蟕c�B�zX�H�L;��m��޺�z�� <��� ��)2��9|�7P������zC\R���u�\� ���=sr�O�Icc�ۘ�|���yOu� ���{}��	�{ݾ.������<��O����{��:�R� ��d��z�f�ʣQ�/Tc���aL�}�(�%�j�zG�w|׏^�.�CFL0��-F�����os��mۜ(#Ga�
������y�w(d�j'O9�xG:�fT�<z���ū����!�׮����y���!.�c��YX���)+�����5�E��A���kA����:��������Wfvj9�����_�e�H!͓q�"����qV1�	��ʴ>.Hx�����7�*�OÉ�;v��/7w�st��DU��!�E�h��,��x�&���0��gz�n"qo���_n]�&����h��(�h���x��7���u����u���$���m�����}��ۓy��U0��A|w}D�����r������!i d^IP8���0����3NI�� λ��8d�ʉ�8�ܠٹ���c�K��T����k��v�8����g��%\7�i��J��"$M�䏖@1�WE��U��L'�6�[�������FY͝��{jMw�>�x���#�O���z/�p��Cf�"�m�^��O����Ud=�;F{����0)Ī��W�8D��'#�ً{�p�k/��&=Q�$R�q��x�}V��i�sWO�b���Y*\ۣ���.��x�����wo)�tȜ����"���4v����,�$�s�����˽=����\�X�o�r=3�Ȝ0���t`Ū�2<�ߊ���=輦�%��o�����>�%��Eb9}�_v�����s�}sG�;�awM[�-��i�sy<��g����pG�O�9�`���o��TS����}HƇ���ރ��i�py��w�+�pV;ѡ$f,����۹��O�9��;��T �XtOx󧳍V���@�c~�$�rNE��@��-)����Y������!��͈�x���%��uIv����7W��v��5i^Ig����7�|�ok�$_MX{�u���;��%�<�:װt�����;�cǳx���Ӟ�׺O/&��G	��@F:�LS����xa��nw�鼦�9:�h3�W��(�@}��&��^��/z�}���rF��Q���M�#��|�����ۆ��X�u���q���:X��,o��Ɛs{�C~���<�ɹR�5t��Ӎ����|�����9�ܦ����d���[k[����T�ٯ��u>뻞�fCG�Z��'q��f�Q���2_�p!�'��A�]J8<�y��}��|�t���`� �Zڗ�^7����M��d����nkC&]�fK�����P��V�J��C�Oux���e'��������VomO9=^=����l���az�r=��@�tA�ϟ���ξ��;�_zO?o����W��� �t]�0�b��B�	e���*C"*S[ݯ�ۋ�i����{�տex9~�Csdݮ0[R&'�����o[�>� �k�Y>�O�K^d�F����p,���x1�7f�V�A��L[���Xv���_��퐁;�ݐh�!�N��< �Ȏ{-��M疼��I~��֕;�T���������R�<=X$y ���=���e���ׇ��ε���O���]�W�s���¤4�S�ˍ�g���\=�L���������3��~�ǯB�����S�̵a�o�C㍥��%���9z�h/x�_&��-�؞�G7׳s�U�Q��:�;po�6)��������.Ɔ�e�g�����Q-���e�.\`]-oi�z��^�vf�z4��A�v\(h�w��2���+�����nW�#O8���5���qI���7�(�y-����y7'��ޛfI/w��n�n�t�������>;�om~U
e����b�SF�O�͘������Df���sJ˰���cǼюQ���E�h��z���^���rP.0}�k��+�>��`���j��+̝������b,�����'�y<�0��Ւ�q��>>oM��%��Jp���EM{���R�M�)3�rM�ū)��d�go��k@�]u����^����싳�Ɣ���Ӹ����l~:toS���c����:���ˠ�����^�8�U�T���`�����b*�H�\c0�?�{r+�v�g�@�`L��|2l�Q��ǀ̲������1�:���sy�;w���^w�֠��
s���=w���C�X��D�4�x<CH�<��R i��d���*���JrU���n>滘}���GK�չ��=�E�����3���ޯ~ѥ{���z�7�� �{_���ڸ|d�G����&K�c�|����/j�k<�c��Q=<<�X׏k���=�,wh{�~
�����McL����<&��XC|g�>�>�QM����!�g� �+����N�a�����>?{={��E,�qw��Nl�����u��8����z�d�.���p݀��#������2 r�J����8�xر��3}�y��fkIa�a:�L�e�OڒK;��Oz�<�{�n?n��9��=�Ϲ�osTy��Qwk��Ge
V"=V2ɰ��'��&�q�����˹m�{�}��=�{����[��'=�C��th��s!!��N�>���(�g�xp]1x#`�Hu����0q|�F@���c�.s����%�(i���U�$��)���F�_�w���e���p�����/�B̝�c��d�+�O�7����n_ٷɞ�P�6w�S��v1/�7�����������~��n܀��=�/��k�!϶�k��^���gN,�Xc�1�۵��P&^m蒞���d��_�_w��ģO٣��S8������B�A�M��Dz]!�0�X��f��(L���h5��Q�o?�Kq�sH<sݧ��\f1&yra�G��M��ovb����o!�4��ǴV��{���ъ�y|��)����^p���2�Z٢�ݳ��ݳ���t�!�-��vz齃5��~��u�0}�;��n�/�ʻ!���y�3HCY��h��i��<�o`�S���ӽ��=�LEX�U�lO#Ar�ǿ-�����b{f漤.Oޥ�)����s��C}}���� (��`6?�v>����_���'G���g������^s��DS=z0��I��Sk��=̾����G�����q��>���x���;��j掼
7����3�����y�q�(.�V��}��7�w�q���H�����^�s�x�R�\HB���R���܃�m�-z��Ý�p���3�݆�Y�gOEd���������T���}�/g�K������J�"@ø{�=���1cz�+=ݡ��.��/�q���'MoEӽvO���]�N��E�W�׻؆�}ut�u��m�6z&&��n����9]����u>�FOS��l�y�Bǻ�<�d}��YH��O6{�:��1�.���{c�EtC���v��A��y��>�W[-���Erv{�1�7��A�,�n��ỷwD�W,�4t[-�7��ܔ^�z��N���9���xhu�<gY=Gl�}�x�����+�CW��l�^S�Z�-yp�;�<�Oz����o:��K�������^�^�'1���W�����d*A�cM��Z���7�[nh3k��ձ�<XMΜ�p�*�Si.�]GVw���!'��j]�A�� 3I���A��>����i�f�(/����M�a�}�|J��Ή�3l�hc����}�l2p��ٞ����{�m�<b�FQZ�v���o,�SJu�w��ͣ��׳�ۜ�V�{=�F�^"�Q�ļ�vf�y�X}u������,�wc�"��,�Ѭ�]ogc�8�]�Ww
�<s���F3ͮ=�v,'{{?V�k�V�3˲�ݹ=������X�V�/��wae,��6��K��1,৻�A��&�3�e{m���{Mw�.]ḕmz��}����3�*�/j>F��\�<fJ��z/{ը��Y��/=����%��X���c����x��\s����y<��7of����-_H�w{)�+��.r@�� �з���Y�3�'wKL�u �׮j��Ng{�z�w��{x�����^\���������}��מ���>�gٹ�&�|����ܷ�)��|��m��1�4K�fI��{��S��� p|��w��Su��f���R�o:�n�Xxg�
�]��"sw[����pk����{/%��{�Q�	�*�M#�>�f?4E�� zgo��BNŎZyo��8_�;�=u�> o�vf�E)���gv�e呼a"�}�J������x���^N��|�k�߫�6�3�š������>���{�P��3�"#V��>�1f�~>�w�\v�&�o �V�/�qN�/��޳������Xc�ۮo@t��zC�<|�}{��W��Ts��7g�����'1yP��y�*B��;[�9�������7<*���Mt.5C�����Y~GWV��!��E�976+,Ȍ���e߰N@�VA�U��h��wsroo{ÏS�8�ѽ�R�f��^��Wzz���|�b�6r��+HJӌ�ib��M�;ܞ�[�;K=�k-����{s��ܙ��V�V��	��[�s�y����=�ǀ���bo���!�\��{ڼx����w�w��V�n�Ao{�S���#�O{ۜ�#+ݻ�J�x�=�򼈾j.|6�X�0\5��ܲmn5��v/1�y��ҚvP>���=�����ô����{R��f���
N�T> j�we�f����=��o}ן
M�(��jZqa�x����� x��vh�\�³��K��H�$,�Oo_C��5�����Z=w�P�B.���n����Լ��NS}U��	����20���x���U�[�@���=�e.�ݾ^��]ŉqj/��E�v[���Z�������g���= �;���eD2�xt.���P�/�L�׃�tէ��=�U�O<�|��ٷ�Wq6u�>����+�\�g�E؍w׷L���_�����{ݾ���6��H�޼�8�q�����L��+��y����������޽��{6DP�����3}�dm�8�H�����k�z��1��.��͘[Ye��x��g��/�3p&
T?�s�&�K�Dk��7�O�]|�x�r(�bd.����*�<���ԕ����~��|�v��R������>?y��� H���^�}��l� �w�f)�0Ww�[���Y�.A���Y���c��"[���z��;穬JpN߇�~_Ҩ(��1����7����>�=�W�ǿ|>8�����*b�Y��x|y���u�|A�4�MEX�h,�������W+8��2�.� K5�6�����牟6�շ�.�6��ݼGI��\���9�T��Ik�r��k�a�L�K	��Q�(jwZA�����/X��Hs�5����z�v�㭹M��:�N���A�z����w<��;{7�\�����E�b&�PWV�g�y���7�@gm��=G*��J؈�p�ٸ����\�U��n��Σյ������+��S�з���r�����t�]vk��#�s���[�^.i:����yGuMP�γcJs�%Й$�wE$n�;$�n��[Ξ`9Dƺ�6Me�iVm�L�iQ�A��m�ts�`���MjW��Kp�K�Ks ��P�n�Z$ӮhՌ����w[�n4�:���8��8��.��Xʪ�]v�f!2n�Q�ۖuO/Gl���v����=t��_F��Oe��ݐc͛d��+@k4#�,я�3m��H�t��<�cN۷1l=����1]�e�oMnp4qE��{ZW��������ɳ�;�e����)�oR�jqj���1����Q�=�7M�jю�<���cl�f�nGe�KW=\v����^�N眻�;��َ�
.��K���ʻX�JlT˛����8zi(�҃55���^�s +��b��v���խa<n8f\4�����&�5�:7H�cX �ݷ�X✝e�1�[���K�qJsW!v#�D�XTffM�&�t�F6θ����uՒ5#c��͐�Ѯz�Z�x؞�X���W��y�g�g!<n$�rn�����������*����>7On�qh�==�e��QIgh�0.GUve��i��ٶT�=�v66s�U��Gmp>S��QkN��l�q���D"G6�g<�B�G]��ƪYz7m��Gn{����&�$k����έ7X^N���l���s�-�"8��6�������l@�/8�7�j����=�Q�A�YEe\�#�^�h<��u�]���nxRr��c��a��X����8��U�K �"���W��Z��\�^/��Q��c7�ö���p�x�,-�\kp�luc/E�s�6����&���V����.���,2Z�^���W\Ǵ�$�t���]0Pkm�F0v�#������I���u�N��:��k\\u��4��%�e�ka�KcVYhͪ�;Unj�R���z(��q-���@�\ښ�(�'B��!tZ��H\�J�5ru�
�y�Q�2[��]���т��$��1�[\BD���볧�7�]��Ɡ��ݓ����j9���c�#���dR�[�]��.�ىb�C4�^�v�b�DL�U��SS��.�ಮ8�P����i��/$�*���v��+��V�l6��Nn�3v^1и(��5�Q*&ҵ�oFj�,�Ds����Y�G�J�.\�QŚ6;��(�K8�����s�:qm8�;�+��jNia듭�p����Ӹ_b�b�L�
�b�Akһ\�6U���`�t��`�vZr�ܼY�Ml��2�X5����g�cp���װ��<,O<�x����t�[1�E�"�5�1��Jl���j:f,[#E��^�B �{MM�����.ǋ��t��2�H��vQ�	�Iȹ{l;���`���f��j�K���H�s�J�r��u�g�p��L�-��ˢ�X�I���̤�)�����CF����;h"/(����9�irکTuE��t�Yz�Hg���i�\h�{�x���)�2�9���a��k�6ᑡ�Ψ9��Y��!v�tx�����(�y�X���;z�[f��E�+H���n��̝�7]	�Ԕ'q�\2�u���2���P��`���y�/g�qg��/^�0M4�཯�6@�cWh��ږ�J��r�vuhg�]3�
*��6�ci���8�������m�n��V\�uj���YnI�M�Zȴդ*��a�X$�i6Ն\e�66,���ͤ�A���]ي�k3Amu��Sv���� vW<��|K,sm�B]�!��Q���Ln��Ta��!6�1��ԕд%����4�*�L�����Z$YUGsr�赁I/;7ty{Nn�l���7f�rӸ�wA�����2`��˶ᣣ���FӐ'���Oqg�����	M[�rff���l�6��v㮌�+Hg1��q6P��\��6�S���kIcn��F�odsy�A�^G"������:.�{>8{d7eo
yn�Ō����A�nRڔ��6��jn심.�B��ic�!4����U yHwcm/C�Ͳ�)]nLݚ��Ny^�b����E�˚��-؅�4��V�JǶ&��t�-���ҹ��q�j!J����n�v�7)��	�[)/Z2���e�iB�V��.���1n�mdC���f�B&*ḧ́�M�w a�Q�s�3m�c��4p���N8�z�k���@Sk]�v�]���m$q���q�vk�� l瓭�� ^{'mn����k˖M���0G7�L�pjI@�:��L�=�*q�5c3t��8g����M��^�v-�(}w��L�[r�+Sоn��.1� V�@��=L�[PMU�Q�;45׹y�݇��D����t!��Ir\��Ҏ����q$�7A��7vx�[��-p�ֹ���ݫ��np�RZY�WcI��M#^�

��y^2m��%E��ى\�S.Y��������M�"�l�t@�#�)Qܖ������"�kbBɥM1�R2&�OgGiZc#��؜�^��bF5��g��<�'Gq=��Y�:���Fg]����v�!\�qvjϮ���/uC�0���+y:	mtpH�Ώ
m���I���ܖ\�\��v�<�Am���!Y�ŉk��mc�Yn�@�SRT�GR�<�92����ܧd������+�1�Cjn���D��ծ���{l\�ۗe���c��iz^kqtU�VFY*ܚ�Y���I�cMf��������US�栆7�F�l�s��'6rqɣ���%�hKT��T�3&��CC:7G=WZ��!+�U���[���<e9�����\��2,n[��Řu�rYV7P\�+���ŶSL�n�kvi�#�a��ZMM�@3`�ap�Kl�Ϝ<5�6ݍ��.m��3��m�7����6��`(�r�����gY��R(�iը�"�\�ol����%.�G#�v㈠"����ض���*)w �a6f�m*B���αd:�g%X��'Z�{�vb�RX�*]c�CK61.���y�n���p�<ƛdh7����4�n���u�{s�ُI��caZ�[���v�ŠY�����f�T#���9��M����ڰ�5���99L�PV�݊��>��X3	�^�Z�͕ٙ���]��S��D+���,�
;Bj+��H������Y��.��S@`���Q�٭V�l
�w6��OX�ƶ+����	�����XN�"[�=/v,�twEۨ�\q9�=�}�$�z��ܞN��Xݷ�)��!5ݒ76wc��t������X�u�̻��<GyjXK���6+R�B��ґZ��\�v�+c��d&5[�NW�89��vgnx�̓v���WmN�����. ���ek+�B;k�U�m#\\l5n�=sBp���Ҹ�#)hG1.Ȅ7`���z3�yX�	�&N܄΍ڞܑ#�n;hZ{8<��n��&e�]XL��3-F`�65#ʚ)	��� �k�j�5�ΓQy�l��m7\i�ɭ��Vx�t����Tbо[8�V�Մ�@�!ӫqF�J�.w.+A�Y�5lZ�t'e:��Z5���GH�S=۱i�%�㱱�zqGK��l�Kۤ��r�͝d֩�p�'9x�Â�ҵͳk�W��:9;MNѓ<����BY�{u˴�e���r�q5��i0�k���!*/�gl���6�^,�8��$m��P�)�j;hb5�5��=Y�����h��ᱸ��z\�;���A��T�Lq�u��.t���OrTV�Y�Z<�u�^�:R�ާ5����:q����lK��-�|ٽ��Íb�V�s�=�t�n��:�<v5��bXy��rSp�	ö�ʛ��=
��a���i��D-\�N��d�����&�[n@��]R�����]e�Ƀ�����5s��嵋�yi�
'G	j�G�ո�]�P댑gn�h�\S�w��Fn���5؍X\kTSL厨.Bi�z��x��Xqvp����Sm���k-�q`�K8�5c�����J�t���x��㒸��سT��Auto������/3����vU94	<���[�r:��v�`�z�ss���xݞ�U���٬�lm�zk�R7d�V�O��<Jk�:�ӷ\�pg����L�l���^�\[5�E��(w�r��˵��)����hq�Ӎ�[L9����e��4�9��n�@䮱�J�m�W:��l�m��I˝��jL6`lQ�Mz�LF:l�Ӷga7��-Iq�Ō�AGWZ��7`^bv�Zh��wC�@�y��N��W��+��k1	��˵�N��	jq,��j�`�[��=��5sL�r�uvR����V�̀�vܯr�+6��]筰L��n�M���z��>�Ք�[&ckh�f��Z"{X��v1@8�Vmd�t�ۡn����!g[χ����QY1�k�Q�CF�A����%�6Z���l�m�M:�H��73�������3�ܮ�"�C9:�+۴�:�MPBӦgg�u�nv��y&^��7,��0-�W�#�w�/�p��3�{.a�j������eA�V*����X����XVW+���KkRʌTEb���;��ւ�YfM���f���YY��Ң�8Dሤ!!��bDRZ�����  ��,��VB�i�[,�&������J��f[lU#/0�I�@�@"�BT�ǖMX�V(@0� ���y����1���Bڭaⷐ8��0�����;��V/�<q|m���NQT"Ǣ��������Fh�U��ŌF �2�I��J;�QF.�ⰴ�P��AXXb�F1tlL`Rq�U8��FE���Y��ZQQ�j�-1*�ŭm��f%Q��"ZUFDeT*�1+TD|jMh��A-��(����S�LHJDBAR����#kz�AB�J�V�m)Q���fQE��(�UTR���T�� ��*v�1E�4Z�*���X1TPA0ZUZ��V�'2䊠����q!�B ��5*��q���T8�E��Fq>BI44��a�8eu�[.ŵ�g�
���[��YB�56�cE�W+1Ŷdk�����,�{'GN6�
��qƍ�p�LgwF�U"bۓ0�Ʈ��s����y���1��/c�,?�tt��N�庶�m�ٹΎ5m�96��8�0f'�t�����G/Y�'j��:l��s��Ԕ��f^�^�et����qs�wnn���]�;��9s�3j�d�qm]�ݛ�b����0���QQ���:���:"�@���5���۩��$ݺ�.�nj�k��1��e�g���{u;v��ħ�p����w�៝�(��
83�v��֛O%�@uf�g�p��ֵ��<ls�6�|�;���a�K<S�� Oo/�Zɣ��K�v]�f���Ʀ���d��0����[��}�n���Txܡ6^c<�wu��f9�q��ҽ����K���ly�v#��Z|������a�Z�y]��uq�y6�1b�p=��KθIzvٮ���:��}����J���N�����*�r�t��f�t!��K���^�ڬ}��Y�Fg,�&�p�Ӟz��7�y��g���H���jY���D�����=k����f��]k&�p٫���N�d6�a�a1]�>g;X.L�h���Ç�nj�YɊ��!�X�⬏��N� C�[E�������ۚR�^�#�1f��s�A��[��j�Ї6 �s�hD.��Hۊ���d�͖C�����nĝ��ݣ�Z
cutJ/7�۝���ixud7=/����Jq�;v벥��o;н��5e9ԋq+f��<R#�m�ݮh�8��Z۝{���\�GY���W�
)����&��'pi�lT��Kt\OL��ag���푰ư3
�����u�h.��<6㛍ۜw,-�M�a
f�9��x��J�S�;������\�=sU�n2��,cl���x�(�s>�{�����6B�����[ (�%,�+X�E���@��F��(���/ ��bE�@xa�YK+U���N��-�2��4�@���[-�m`�أP^x8{�7".P�q۰�-cZ�����#�hpV�0�mie�F����l(�Ka-,�yKc-�D����<�*���y��獝j6�ieV+~{=��ϭ��͡?���
$_���D�O�цM�۾�c5�.6���I%���V2l8�A�2��T��Z����<���#���������7}��g�j���-vg�W��F�IHB��,j5��D}lA��o��F�����	����Fj�D��䐡D��90��7^Cg=��[B�	��D��������ޛ�:�ۯ�I:.QA�3(D�5<_^�p����n��� ��F�� 3Z�~'|�� s�!Z��Qe��Ҍ>�w��\�g�ْ켉F̵��,��Y�͆�l-^Xkw����O}ڙ�昻��=�7���fP�@$o��(�Ή�ʪb��G�%8�TN�-A �L�!T��}G]׉�J��~6�����M`�l������[��'����T�(��F@��Χ~���!G����ׂ�Y�ഝ.*1p�|F�կ�f�b��T����N�������:�G��D�
eV�|�:A���ʑG�{j�<������|X�_�c㏼����R�1"��󧞀�o��d^��A$Fz�B��׬�s*���>�j�3�&�
%���ĂO��A@�Y�����w��>&j.��x�X ������N<���6\�1LO�1��3cZ�Eh�MNq�YM���&�2!t,Cm��oN��3&fP�[�'�}���$#���Q�e�1�{q�:�\� �y�c���Y�P�B���O��c0>^������+g����+�~$׵@�=�R
��I��I�ޡ�4Ũ!�!�*�N^W��;��A'ڝ��b}��[�+����^���,���to�G^��G��W��о�n��x���͛&�e�8+|-����
��+&���f���/Р	n������j�LDI��S`��{��lnj�y��_�$�[������!��b5i��r�dWĊ�L ��JB&$V����
?V���U�Ya3Y�F~H�n�*�$/Fj�$��|�;���`�X�u�c��1��9t��.��x8'�6��ͩ�6ZK����b�!���`C��#~ =�&�/F���4�P񬝑��o*��X$�̙�B%���A� �-˖�Hy{j���O�󺯉'"�eW��_'������@���C�4j�@_ ���^� ���A��U�w����� 弪�-�_,Z�A�T�P����k׶k������뺑K�N=��$�3�h{1�)NA�;S��V6��}ڽf��KY�ui���V�E>sjY]5��p�:��WO,f��C��nvw+�h*y��\U���H1�t(�ĜB�
�%2�>k] ���EQ��3�(�cjh7�#mP ��{_lf���4}krO}=�-}K#Tlњȑ�@vR�lְk����LJ�Bm�Gf+n��>��/ƴte��ߍ�:����@�H�=��'"�D�/��+�{� f�.�̒. F�Dnl����|G�]苯-ɽ������Fzl�|��|O����z=�t��
 D��4afL̡��h}odP$��!N/n���آDn�
'�w�hS�!Z�r ��I���l�֌d��Q ��H�K�������W�M;������ l���A������;{B�'s=Ua��l7�ă~�ȢA"��
��7w�+0�	(��ؐsQ�G�?z��.�h�ڃ<��۠g�;��6�`s	�0'!�������*k����6�g����#��Kt}�	͈%��k�`�7hI���+l��ё��h3oݓ��<O�xoI�&s�;�q�Gb���j�tfpC"9LŌ��S�S�ֳj���e����;�:��tPOb9�7n�c�L�����u]���D$(��}(�i��k3ˌ�gT�5v
�i�\�;�d.��
�J -Y9���u�G�ls���۱\VU�k]��%�1�
%�����ьv��d q��3�ܶ�r�}`3b�(����ѱ@*�ʡ��e�i�H$���I?Gٻ��2=5(��ݡ@�N��	���苃$!bEYTAٖg���*M=���ߕ� �s��a��P8�j϶�?MՉ{����X�H����pJ�)@�ddϨP ���Q'��f>��ۙ�Ò��f	�y_Wĝ��Q�o	��2fe��}&���1Q^K���7"����P$�{v�꠳���^���~l�f�K �5I���O ��1I��mK�|ߟ��� ~|󓂡�{�Ay��t��*p�/��4�T�ex�C�z�c�K��6�NT�ڳ���e"b����A�� �ۡ@�H�=@Q$#ٵ��+����&�$0 ޯ1����C�t�p�/+�|�������sB�٧dA��LW�[J���d�v2��h{�Kw�>T��k����]���ܽݯ���4�v`���2��]S��ˋs��A#ݞ�@{�< a�|�>?��<����V�5a� �u�
�{f� �@��*�tl�>�z�c۵�%#�lJ��& �lC�7�|�����|�Q$��M��|���*A��M�IݷT@�禐���12�J
�3�"���@�p˜|��� �-������~ �>���r<�9���u;�3�u��l�ާ,�#�v,R;9�͘�?�����f���ׯ_�X\�&&�$��5�$��h�ww�T���zl�#S� ��"`r��|	R��w6��վH"7gH�w�hP$�&$c����Um���A�$%
J
%1��w�D��y"� ��&(:!N��dh*�Td{ʍ2!���	�n[�V[��kr�t��� O/�����-�4�
�:f��`<\����d1�c;R=�{yr+@ ��Κ���{"��Ao�2
1!(��u�绹�|�N��An�2@$��y��.�ω^�"�IH�:&"&TP����~$�搜EL^�3���`w��n��$�������r�V؀T��ᚕ����L��4��5��Y��+� v�u�`ǆޝB
Bd��+@1�.�$�y"�$Nn������[�~�	��=��?���$H*I&~&%�=����_��U�W;,H&��
-fǪ�Z��?�����$�W���)R��_�_�w�6� 3��8�q��^��@$�kg������,TB�%��o�;v��%w'�0�`� Fo� Q{~����e쌝��y����lL��I��ٽ���2{����CG�nk��X��0kJ�XCۺ���^���:�#��_��y^Ę2�X��j�U^̭�(��Iϫ.(P$֥�(�(Ģ`LO��2���1~٣�`�*������%���7�*�M|c"w�ʥGm*��2j">�1k�q�`�.r�j	k�H�q�%dƳ���a:���3�����>�ɛu�[}��Οd	�^z�"6�M~�FVC~г3��>3�������7#��HĆ�sQc_�i�"j6�� ���$s��5O_�N-;*}��c]h�g�[$%(�?#�^��G�LnFR �;1���a��0�G���q��� #~J0������&�Uj5K!_����}_P �����_甬n��W`��[�q��"�Jc��$�VO�顋"��E�ǀI �ۯ��a�I�(�J���������W^�<�#�B%�����I0�� ��ܱ���jˑ�'���xrɁVD]ȫ�([�� �^^�15}�Yr:��3���$>���m~ݭ���ui.ҥGmv���I�&�N�<�]IeF�cv�S�v��-ӳ��F8����=O���ݖ�j���f�\�)����lz��k#�O1s+�	�Z��s��t��Y�9���NЛ3Z��*<󵵻Jg3�*��ďFy@9��7>-�Wu�yy�AT헃���MR$�邻��v\�ΘU�k]��,�1�'N.�;�)��n9뜇T����Y;[�vSz�s�]&&L�0���8�E�	R8�ʠA���D��hQ���u�6�z��5����6����H�{�Z�F쟒�KVsW��7�.js����A~{B�$^7���*��s�"ש/��12�J�c���$��ȠI%��_��t�g}>���|I"/gH�Ny�
&vk�"BR2-�^�ɼ�m*��߂���Dr�Р	#w}R.�e�D�S:h؀�4��D�5����(����Z�m�k�8TH$L�Y�A n��D�Fn��@���yN�fl�	�P	�0&HALc���ű��y(�'j��z�id4jGh��������_�`�IAD�.�@@���E� ��li�>��2�фx�w@]#��Q�@��"�٬�Di���b�1:Ͻ��]qʡ�]�S���<�yyi�Bշ�;�{/K���o���3R�3d�W�j�'L��v�S�j�/R�����`'�״(	9������3t��4���%�TB��bɟP�~$��W�A �=��Eи>�oM|O���wB����
�u���L��B%P1Ƶ�#�UƝ�r	.�Ƞ	~Cٓ4	����:o(U�wM�n��[����X�*����,#5|�fՊ ����B�Q���^��D��ۿUO��4dEDsقlăJ�2)��[@��^`+jv9A��I�20��^u�#���0#��bD�Dz�	��V<o�����u�kV����{��	�_��D_�f�1�HP$�bc���د�q`t%��ZW�gf	��s�p�:h��ldI�:ݰ� �J�t'v��>f��~~g�*(�0�'�?�|H��w���G�H�wE+ɪBpb�f�3i�bz����^ݵ�;���X���~��1&��s
��~��؜�2s��WQ�����ڄ�e�at�yB_s����2�}�HXz\���N!��<�5-��AOt�c���#��{�n�'>�vr�I��׵�tp�<=E�B�Vy�zR�پ�e6���3�E�܁,�r�Z�D׮��w1�ɽ���R:9��:���|K �i��{j���y���4��N�^+<P	��ǳ�<��r��ߍcebe���X�\P&J��He$�<p�}���[a�#=2F�����?j���Ց��3wݝx�z���2���t��/�����X}�x�@��-_.Λ���ۂ�<(;�g9b�9��ݝ;�`���44��v#&>�$bb��� �������9��|�^G�� �ʦx+O�)T��ğ����O�ªLo�z��i���>�x\k�n�kS��n;�vsw�<`����t�w8���A�2��&e��v�FΗ�%���l8��{�&��v��o�`��P.�����'�Y:y���ؔ~��EE�<��]{��/zg>�&f�$<�.�<9�3Io.9���`hi��M�����,�Z6�~>��G|�����=���w�����;�ݾ{���1���-���.-J��N����u��xQ���G��x5վ�@�@��k��w]B�G��C&�(�x3<Y����.���o�������I�B�Ƶ�ß���������UN��J"Bp!V0�
�VV�,V�*�Eln�ƨv��7
��EĪ�Fd����y9Ý�c�������C����HQ�\�1V'��q�TPƆ[�z����H�cMh����X���3�\ZR�L�d���f�ڪPC��{�g1��i�����V$Fb�HCƶʎ�,`�#1,KJ1˴�/���D�_��%$�� ��s^�	�H@��/�H@�`HHQ�Q`D��a�ń	�2Ȁqu�˂ e�� �"Ȕ�K��HB�tͱ��HJ�Ҽ�T�M±D�X#Z�MnZ�J�M��Eff\Cf&`�Ҩ���(�QR,D���������''F��̋ƣh�Ц�d˙�T���q(�2� ������qTQFڪ*-�QV+��*�jV*�,k)NaTYJ�00HŇ(�j+Z� �V�J5�
p@_׎!0�8�+*"LJ �D�hҴZ�m�IJ� U���� @�*�h��9
�J�b5� �DF�*�*���͵v���Lv�F1��Z(�-��Ҹ�������lȞ�,�J�o�����I�	e��=�̍�����Z+�%D)�F#��dX �n���ylYW��5Z �� D���G�v]]@�[��8��6)"�}� ���蟾��*3�r��9�Y x���R�~}�@�u����~�+���n�8�":e���㼦����Kh�oγ�$Nx��}�o�~&
�w~��:�H�X�w���b��`X>u�'�����
���~����H���>��ac�M�jŴm��-QɍO��i��.��Y:�xa�Z9|y���ڋ��$���$���]w�	�&��-`X�o�;ˢ8�H�!`��:֤RD�N��x��qw�^1��M�u��G0Y�P8�y�F�`����
���e�� q;7���: VQ����}����T�w��]@�[�lK�}�����bX��y���D �lCy�9|�7�"cސ���'�ٿ���n/稤����r���$R�'���M0K,��C~sKz���m�[����'�
��7���xE�P�d�~���V������W]nw�Y3�>l3��uߞC��V4`X�w�3�LlB���y�ZԂh�	Yb�-<��x(����z#����S=s�ɏ���3ޮ~�jC�q/�fx����+��}��j�����z�U��|i����߳�Y��{��xE�S��m���ۙ���gHx��w��t@���FJ�u�<:��s�X����o<y�9$�!}����H�����F�����Ϥ4��C�+������K����"�6�ݜ�I��M;F*m�O���%-1��w�E$Ls��)�,Rڥm���� �R	aH��~y�f�X�]������G�g�����H�`R�o�4ñ%a�{����w*f�I�aQ�ޟ�?~���꨸ڏ>��꯼F�(B�k��[�:�jX%�)m<��xF��R	g<�ƺ���;�'�����|"&NM��^��&n8���&<�3���Ho����P)Ĥo�N7ߞq�3�9�;�d���b���:�QI �lRA�ސ!���5� �$��*��s�r�����Ξ��u�"��)h����
ԅJ��O=��0:�� VT�=��C��6s��}�|�?=�8��d�T��{�aԕ����e��
�m�nt�N�*o�ό2u
�H'����|�s��u�.΢!`�^o��	�X��[N���5��(�G�>����J���gx���n?ʚ��ӽ����c�^5��7U"�$K�>�ji��s]F��0=��7��V�b�Or�z�i�r"��|}i?I<_�y�	��m������%�tn��v��lE����]��z����e��&vPkYȄ��n�	6�=3\�q�BF��0��Yt,�����K!f��|s�F��a\օ�K�v5�1"�֚�Z���E�`�����g������C��9��͟��#Î��HJU��C,��tTwf�#�(λ��W*�;1f
�<xU�����c	f� �,-��tc��!tq�|���q�XK�c&���^�?�m�Z\�Cć�9�qg�YP*����牨��bؤ�^9��hdD�{��]���S�&q���d �lB�ß<�;�%4��{1�uۚ��Hu��u_Q��Kr�|f�����r�s'$��I<��3�MZԉ��� 3�Ȁ��"���.���>qaؒ����s��[��iS7��'�K{�sCQ5�h@�8���]���<��+��1s��ȁ�b	e�[O7|�Z�IX%���}��N��R�|կ�&�\n�D2 ��tO�0�����y9� 0���H��몆`h�bR�N9�z��:�`ؖ-#��Y�x˓�y�w�x��5�a #b�ww��`����/�Q�5��o|Hy��}���G�G������E㳷�6gH����	���������t`VAeM���tl
�ᘁ�~s�fD����o~�z#��{/�����Lus35�K�r飝�u�b�1��m6�]�Vݾ���������s>�I�0����l2v!Y����Ȥ�h��y�;�dL�Lk��]s4{^3��R�r�
?|	d|D	��B)сR�9�j~�sn�gHx��M�??����� ��ݶ�"�a����7�����U�}�3��]��o���ϯ��N�3�r�p�U��F�j�E����k�	������C=�{�f�[��)�{�"��+ �����;œ��@���םc����n�"�f���C$.��ϓ�]�n���C�Xo�9�u�Kj��<�=�2j	e ��XkSɹ��q�>yP�)"�>C�ߞk# i�`X�#��s"h�bWs�7���"J_D����C��{w�=��FoǬ���+������1��VJ��:�zԂh�	e�V��/��c�����u���RN��R��Z��h�XS�5k��f�n�ć�9��Y����yf!�w�i�P<9�&����L�޶�D� �u������b�;מk2.�X#b��~_5WD��a͵f";���4|�k�$�.LqZ3�Qû\��d:;-X���
e6����wD,I�e@��#���g���e�[T��u�}�2j	b�)!������~ث��C
� #�!�7C j-�B-�y���dM0lK�n��̟&m-۹�d���P�a�J���י�S5/U��˗_X�? �,B�����֤R�,�J�w�������#Ѿ�������t>�</';�g�?sn�g�?� y�{�,�YA�FJ�}���d� ��#�~����/c�9~�5�y�@�$Q�o_��#�	��L��Xx�X�}�k�]������^�L_A�5�����P�0檪�7ￃ���}}��,D�lu��Z̋��H����W�i�Rӛ����s{���َ�|+���j"ǉ���/����z���lHT�
���>���u�YD��eN���<jB����Kk>�H*C=�yŇbJ��sݹ]��-��'�<Q�O���(ta�J!Y(!bo8ߙ��	������=�l���y�ZԂjX��Ho�ު�a�?X d����~Rv6n��lt�}w�9�4j��	���Yza��Xm�>���Y��n��T-]�z��	��I�ڶx�<���?>��: VT
�d����i�ME$Kĩ�g�4<A�K]�پ�3Ϙ�8ζ���u��2.�cb�=�;d�u!O�xe�j���p��	qל�6ME+j�狼��8�[ݖ^�����MK,��,)�x�UE$t@,y��^y����/|����g^�|�?�}���1��e"�Ɇ�Jv�i$Y�E��S5�U��0�I/vS4I,��D����&0�L�yt�cq�O��+m�蟒A-�O�h$�H��D���v1�f*�YTK�����d�y��_���3�wc6h���}>t{6�r$�{ղ^��y�ǯkk^�ߠɭ�靻^�0�J�6o�wT���$������>	d��Q)�2�����?�+��_�{R�Ɉ����@ ˦[I|Y�M$�����X{koĞ~P! ��f�f~�M@���e�%�&Q��X�u6����ŋ�f�[���fF��f�	}C���|�M �#+v��Ќ|����%�\�{�Nz�n>�L|n��0���NߤʈJ��o���	������nnFLަ�I!u}T�A%�]��D���"��hU�g�5�k�	$�}3�o�U��I�͠�A$��Cs`�g��"QʾtKI��a�ү�З���@��\�J��VV���ƛ��J�w��I$���Xm$_��Ͻ,wUj;FZ�L
V��I	v��tHQ*d��������A.��ӃTil{gʘ��#��}�	��a{݌0�@$���e�ѻ��@���n�#5F.�}�|�M�;Kv���65~{�s��kǮ�Ƀ �[ꮊ镑1I	�͘D�6*S��Ĉ����F�uk3
�]��3\�E�(��Aڽ�OEG���d��]m�?��|��F 땆�mu���Uu�ª��ۓvዳ!k��ț<;[qs%\+�l��!����2�׊�X�M��k��o/ZƋe��F^��N��}��F���W>+OC%�ͣFC$(�*ѕ#PRUy�7.�f�������*���5\���֮����PWhkj6 ˩0�䐚b�FZ�5ոͦ��])nW[�������Fڦ������lJI ��v�`"I��f�Iz���q���	�K�����#[�3 �0
�'��]}>_8d����!��=z�k�R	 C=��%���K,�>�c�����Eoޜ̨��&J��*!(���a��I��Y��K佘���b�˾ذ�	%~�a���$���h���؀�%�#'��7����|7�$��$�H�I%�D@���d��ʍ���,�u�X����O�
,	�V����"p�ݿ���I?����=�u����*���D�P�A$�kƈ>^����p�^�A�S�&�����	��:��z�M8�%n�x��.ڢ9�as\�[\ѻz�Ȍ'��2�L���(ʶi�e����I%���I�;��ٸsӴ(�$��S,4���AA��fTJo崺۔Hߠׂ��
��O�%��\��Kk�.g�*�����h)$x䃱r2D�pu�}x�4�-[�����z�!r[��V��G*�{��`� >�� rw�9�_�n�-���/}����_�������5�f�� �K~K۳��k�����#��H$�JE�������Ci/�Avm3F~O�LF{g�a%ɔ�`�%D%�M]f�b�
�ᳵ���}�U7>�Y�%�K�h��}�C��E�˩w�!$wW�.�n�$���a^��_��-$���5��=>�Y�:-��v�lէ�GЗ��u�I k�T�1W�6h���jR�	�0�8w/���qv��n�&��S8W�]�E��o<mB�3�2�R%tr[^�&�@%����/�_�����A}gB�J1f�ӧCE���i���6A�"bL����˦��W{��K��7���'^�5�$�Cճ�0����@��ޡ��&�ß�jc<m�$Ep�QPfaJ��][؄�H%~��i|�J��a�1�����I�+��:�Iц��$��'6�̈́#�~��K���g��>�K9���׎�WWK��%k^>��������}��cMpH}]I��} ǻ(6�sq�I3������@{�}w�=y�_E������$�瑴�($�ٌ6�+���Ψ�F�����Ift�M$-2� FA�b!(���a�I=�-���{���8��I^O�a$���a��A%���e�cd_�g��(�A=�|.��MH3[	Bi{	3M��2���ʖ�s��c�]-��|�=���5�g����]#��%��A��I��S,�ǼV{�,_�����[S�4�����I��aA�3�8iuz閾K+xd����U�ԒH_�l�(���߻�w��iNN�I},���dL��x�m�%%��L�PK��ƚޮꨨz���Y��h���6i	�h)(S0�`D���E���r����={A��I�|�Q,$���@V�_ݿ���7}�����_�����E�8�4���f6&&/ws|�L���,t��ZJ��ߦ�������}v�x���갡N���p}:�
����{WwT�3(A1�K�]{6�d�;�4OA<�ޥG��uQ<>ڄ��l6A$�2��ZJo��a)�Ю�w�D��=��6.�:�-�4J'����{6�-Ŕ�9�5c�uQ��m��~g��e�)mP6��[z���A,ݖ�M$�K�7�L�Nݞ�yӒ�O�;��X
����7�pHO�Q7O�X���"�y���I%�xz5Dk��~�CZ@$�Hn�2�Ig;���H%]�ׯU{�����w��HvBPF�DI	D�)�M��I$~��s�A0��{QB®c�_$����`4RJs��i/��� ��0&Dʘ��]>��o!ӑ�4N(���}}�$��S�&�K����e��)V�1��*�q��o{�$����m)w�T)�S0"S��:尒%�Uy�(���u��i��g� �D�=�L��A$m�5#�P�����R3�H�k��9~�5��5�l���ɡ�$�U�9r-bʃ��g��檔�^��{��*���7�}�7r$5����Z�G�Т���	��;���m{K|2������+ˎMﭚg��'{=e��y��A�aՉSRz�Ḗx���b����7����(g��zeY����z�U����>� ���{.�}ޣ����<��W��+�t��o�����`�u�|{\�t��P��y��Vf��y\��^�������{���#��}HC���(�ݺ���F���"	q�+�0��DW�#Q7�[^���>�{.������Zfv��1#���_��M�t�a���n��y^4�]��)�/87k�-�T˓l/z���bѵ�����r�V�����}w����r�e�ݸ�7ӱ��'���Sd�Խԙ�-f�R_]�B�X�on���=ӱn�x��a�|���	��w�Ӝ�;e�@���iH+���#ģ�k��p��vy�=��}��=:�����,w�{�{�żY���I�<^�oR�/0�/aP�{ΪO���=�̲=輙�T����M�{����W�������v�>����M@zh�>X�;���v�6��˟e�Yk<A��`�m?� ��=�US�1�wl���M�!�){��.[}�o���t����WO��G�j����Uq�QК�܉���s��A�]����{�{�,�;�{m𺋨�W�0M��p*01f!�Y�!�L��S4ǈ�1i���~�+������u�w�ZL��z�=x0�YG�UE�˕0�,�	R��Hm��b�bG10���9k
�j�'�̛;>L��b3=R��*�#Ѐ���)�rJY�Pj�[b)KB��k�A+L�-g,�\���`��6Y�g'�����>V�]��@�(v%;�1��U��G,8BE{cX��-XĶU��Q�F�yʦm�xr� ^�y�y�x'��W7�3"�%A�mX�mq��X�[-a i�̧u�4��^a��"QYHT��N4(]K�nlgl�4�s1�Tr�M�E6�'30�X$����H�%�⵵��3���Ъ��q��s� �Ђ�$񊘛��R�!��x|�a��ǆ�miٌvBYP�#�W(S���V��F)_$�<���Ԍ��ƚK	^�I�F  tc�=))�ׅpJ������YK�m6�qDE8�J��q�Tb�P�������o9o{���k*.2�W늜�^��*��tșħ$�u��v��<�U"(�tX�R$a	�ZLJS�w��U xu���E�}�@���=�*4+<G6���X�[�B�;C�ĈOjn�huX1��tѲ�i�cf`�`1t�͑�ܶW�'!�(��Ҧ�kn^#R�kP��8�%�yx��5������;@����BS��:'Y�n��lYm��.ޮ0'S#��>�l*��sq\GٱV�wdvh��3���녻\��'��*�깪V=�/lW[�i���F1i�àNgV7Sr5�Wm��F���e���p��q{if5���ww]=8;f�kcC�C��OV��;Y��y���]���=�N�q��z��-p\m5Ν.
�'L��iV�n�+E(P��ไnPb�;x���`��;���fS\F�]�`���;�J���6bh� �F!%l�GJ���6ӳVK����kk��^�IV8LdRwn�1�S==�λzN�$��v�W>V�`C؎G��ѹ��μu��+WIq�[f���+��<G F�f��1W�˲Mb��v7r�ny^��'��z�@BhS39LF�٦ci ������ppt����d�K�z���h�oeH�鋨EY��
��0�nCm�,fܪ��/]�iQf[����Bu���ٱF�Ԛ�������E;���s�\�����[g�<�:w]:Ƥ��<n'
 �͝ǎ[�z؜h(1Q��vv�B �א�=]4W]VىFŸ�_���e�u-9k��k�eс.`)Ϩh�}OA�W���i��&*�Im�i�CQ��O�Ap��)����Y8N�k�5�#d�z�g�����uj�Uܻ��[Q[u��+������ �XمS3s�Qs	��Y���S��k���utOb��n�%�K���	���af'��	�;��iݺ�燞�Q�P��M,ų��ݡc+tLF��L�yn�٬lu� (ĝ�����3�U�rV�S����>��z�,��[M����g��g���l.j�R����������;H���-�-�V��|��:D��ސ�d뭇su{.u��
� ญ�;E������5c�9�(2p�����ɩ7��S�uR�1��K0�0,���<d]pu�ԁ���7�L�׫��3��y�n�+�����0����y�ַld�6�t�H�2ˡ�*�woFz�8��S�=V��]E�Me��1+����p.�s�u�&8#8�&{z坔݌�Úx���k�Q���q�C[CJ@�í�>|���S\��O?�_�|ᒒ�͚$�@$���a���fϽV�M��=j�����2�ICʢh���B�.���g0�A+���"��~��!������I>
����@$ꆭC����E�⣣sŨ�"A�bfI�����-��D�n�m$���f`�}q�����#���e��&�:�&>p3�(#e�W��OG��v�l47Ր�'1��A$B�u�I/�=��հ�D�i!�Ιa)��H<$L	�2�~Q�l0A �]q�Uv�,��f�7�@$��4ZD���Xm��wOy?��R�#�+پ��R���]�UƵѶV�F���
^v��v������ψd�I�cןwТ&bb`)]�on[	 �	U��mJޞ�d��Q��S:3��H�U{�6���r`�J�}�{���b	O=ټ��R�W���>�w�t^��q!tl�]�߿L)��g����+��{��5��M���}�^^���QL�m�Ļ�ｋ���w6���3UeMrK���%�^����{ʉiL�{{7�H�I˿oX���$A��KM_�Xa�':7�i$�M��[��J�V�3hNW��I$n��)$ޞ�`4�|�x�RLA30O��t�[��N���-�[�HH�ͺ	�HuO4�|��ަT�\V	�Q�$�<a���7�( ��e�S���c�I�{f�Jr���T��f�뾯�4�A$�wɆ�Js�h���d���uz�2���[AAxЫ�n�d5�q��{r���f;�*o^�S��u6Ɔ��=~������ ��=b?�$'7���	���[�#Z���a�PI,�X[Hxa"""ff&��ozj��$�OW{'I5��_$��s��H%�4ZI&���J���S��Gf%� G�-�%�{LJJ3:i��D�|9��f����.3�N�mܳ|K�y'IH�@p�<60&����)�/D��<�*<UsͰ�+v�*��o��|�����}�|I$�:��$H-���)$#?~�XI���07�2�"%4¿g0������W���%~�K!$B;:�a$J���>0wA���IO���}��(��/VG��	$�rE
Kp�n��O����	!Y��%��z;4�F���p�a��D���P��%*�8]p��2��i��I�=����{^��u=�Z��*�H����M懲Z	 �jͧ>�"H��)��e�T���E��UC7�P'��O�gE�J`̉2&R�es���Su�7P0��%��OW�k�IB��,$M��Y�XMR�ng��a�0�33J�����IW�A��	����ս��~�v��H�ֺ$�AV�0�i}�W;��0TJ#蛻	>yT�cel���ƻ��$����J~���gs�E����1�{�9���T�Uuo�f��{-���{C��}�?vyh�UD��h����g�j�=�͚L�x���9�:&������'�� � �(Ok��<���x��W�2�|���DǗ�����Ig��,Q�/w��;<�4���!���$���x�umU��޾��x|ch�V��v����Y툁��*��\��.��U�}�~���&Q�pM�$�Owh0�)%���I�����.�;]���$_ v0�C�l����P�������[�K�=�(�U�I�}z�$J��4RS-f��#�\VQ/�g��)�Q&%)��=�w���	 ���
$���"�H�{L$~@���m�G���*xa0b��L)������\�/)$�ݠ�K����a��Hd�U-�z�����զ;]�� '��El�(�#�x����I$���M���.����^�H=�a��I ��D����tJ�����w"=N�Dܸ�^��>���C}q�8_�ŠsUٰ�����d0_~�Iv�kj�M��"jǽnJ�䄲3̻1�iĀ+�߈
1���Ad��	%���\��i[m���K�Yq5�(�^2Mf :՗T�6q/b�3n�n���9��>/$s�Ū[�f����n�]s�*x| vЗZ�a�e�l���m�����9;�)2�����[
�3˝no'i�<�]�ml:�����qhLv�������e�ɺw���z��]���vswC^�p�M ���آ�����9���[�/��h�=kWonr����Z�ƺ��ەaZ����>���~G�DLR��]��(��}��U?�I��;�XIb�Kv<|U6I"�^��6��bb	�2f&Q����y�I(�o1%o��s�Ϋb�|�H$�c�I$�)�r�H��{����}��cb��!�@C>�)%3	��VZHt�u0)$�J�,y��5[	$�]�Xa��Xgz���rLDJ�Je/x(�[�̌��	 ���2���$��g8i$�~�a5d����=BE����}!���!A���H����[n	,$�:��5G��ij�N��
Ч�	z����$�~���J"�Nī�$E�iH�Yfb�y
�*зJV^�6iqJl.���{�7#�B�߿t�bT����%�{B�'!f�@&�u
���ݟv�w9 LR~a�RK��J���}�
��R!LP���s�m ���e������3<�f�����~�Ԏ�'�-A?�ߑ�c;�r��`������y����U�Y��7髿.f+	�>�~`1�1���I P��T��k�[+��4�I?~��\�-����u[Z-���,L�1���>�U���'}�H$�Y5�Z�����h�x$���$J	����!(gD(Hg�L��a�1��.��jR��zK	u�z���	 �z�%���w{��{w�j�xa��@eGk�����	&��Q(ػP��a��/w��b�}}>�Y�I�����N��mP]��KS�~�b��S���Jۦ��� �m�YfXCL	�]��p�B.n�Ѻ���U���?{��e�6��q��v�-�,$�6�i$�I�s����ɽ�]E>�i��I'��Qu���̩��>��K���ů��Y�I.;�.�E�B_�_<�a���H�{�Q,%'n=���O�\2��Z�%?d��h�T��<��۬7�B�
Il��Z�$�e��e��(?��1�����z���s+;�C�{Ɖ�8$�q�'�C������3��a~�0\�Z~������ָ�<�z���'q�=(00UH� Ov6���$����$�ߟPc�}��ؖ�;���"JWM����]���H$���K�K����K�]<��vw�Ft��>��`��s�J���Qg�L��a�c��I/����p���6+vw���%6���I|�Y��a��Hd��O䲨�ꊇ7�d͡�D)���4gD�Zz6���6�3�>=N:M>l������I�0ffR�G�pQ��H$�YohS	 ����J�>�I�׌�d=�^�c�){��ڀ��	�SR�M/���� ���p��}�C�4�D���6A/<}�ě	I���Z�.�9�!X	.�bɓ32$/�s	�]\ZI�s��	�N�CU��3�R��I|��vo��/}	}�z�h���u%�Ǘ��g1�tv�=�"g����I$�Ve2�_�{|�N�^�EtVU���ܷ���K�"���{W>c�������뫸���v����0������Z�
�X��K��ce���s]¿�|M?HC�0�� j���� ���0E����D��F����A$���A��������V��L�_� =Y��I|����6����<|ߝ|}�{�'���f�Q&�����������{P�&iunjh�h�s���gϭmg�,��!~_?K��ך7߻ǘ�Pd{|�a%�o���3S=p�0���@��L�B]�$N�FfeDI>����D�w�'�'Q �dluX�JK�y4ZI$��h��E�G���-�@Q�g��R���0e)-���-��%�u���N���z|v�!吷��BD��M_$�{|�L�Aȑ32$/�['�WI���G�kʳ����� �Wzi��@$OwXo�I.�|��)����56i$�L�^:B �G�!)���g0�i$�K:�~L*%�D���S,$Iw�A��IO�zg�<�'"�*n��e��?�'����o*5���K9\��?XvR��̰$38�{�J��+����va%p��/
op��ܾ�����3�Ng���O�~�0��;��H�]�m7kU�*F�۳���X��$t6Z�c��]���/N�U��mҔ]�Uw�Y���[���6���{mv���xateAa��3:[���:�c�t��)�2��N�CƤ����]vn6t2�غc3�d���:��=D���e�#�V�'n�uQ���y:���{9�<�;��Y��vR��:���D��t��6�t��h�u�L-�1/&�Zh��Ƅ�)f�h���-�n�>ϱ�6���30���:�[I$K��4�H��/�%P�N�qg��ɺ�e��E�u��@�P��� J*&<�
z/�O���_� �	�Ȋ��@$�y��%��ޗɴPK�gr}�C�8��p�:%����|=��%����h$�K�K���uod��?0RH���D��[��0Ҋ:0�%�*D����\�yp���dfXI�<�?�@$�^�|�I$�w����N@�{�IS�a��}�v$L��+���+�C�D$��f�[>��t���Yi,�l2IagK��E%��>1|x={^�}>}��u�h�nP�=���y7<��Ԛmv3�vce8�]m�ۿO�߶��Γ	)�F��/�'v�h,���w����Y��9O|}��
���I/t�*/7bf!D(�3��/���DL�Dmr<J�~>lB;j�j�yv�ԓW��n�s�Q�q\@�Hz\��x���s^]�/P��"zc}�ّ1N�po�ps=
>0Q�EP:�s�Y=��Vt���I"�{���H���w�I��h�Tƴ��
��a��]Q~T~`��Κa$�.H��{�)ؿ�H��r��/B��,��i���FR+urӿ������n��])'0�8�T�`$�ʋ���@=�aҊ��I��m�B~�<0��B$ʑ)A����7)|�.�h?��n=��d�u���$�=i��I!���$�	�c�ǽ��S��z�������iz�����q��`�c@�)��q��!uǞ�Қ������n��%}ϒwP�!e-ڂ�H$�}��aw��4Lb{5�f��WOja��Y+�����Q2"#&
*a��ݬ?�I++<��qr�*�C�����I%�{����).�9xg�:)u�/}[-QkoFbf""I��k�x)��lJA$}�A��K��,wV�DUl���/��.XO{���zN��d6���U������\��G�w����nvkJﳯ�����P�Ls�}J^���%1��'�L��2��k]��u�?]2�۞S�Y�=�W�4�� lR���Őr���e8wWݹ�M�{�M��N�M�/����H[3���}���|���$#!�M}��::���v��o#��s:-~�ȣ�b��ż�|F�T�U���ͯ=�n��=5�vx{=��&�tI�4�4h��=d����h��pV�V�h��G�`P�� �3�LF@�̫7�~bPzg�Ac�����'���ؕ��w�F��v\'777.�q� ;����������{9#���dP}�h!�C��w��}��Liqh��n+�,M<��Xq�w7R/���/���!��h̀}�H@�ƈ}��l�^^>�������uczy�/�LI��
=��w�'�'���vo���ӻz#���>������I)�++�C�C	*��ろ�Wdۺ��׊������gkaY�D� ���7<8�zr���/ݝ��k��&�eL0��;`�#�B�_z�AWǘ�����b�n�+$��g{�7�����|q�J�e�{���'�!�.�;�L�^�\�66 ����[�f��n,�6��������rd���{'�{w�{�s˶�gj��9�>~<�~��l�P��O>�7�V���g��ŕ�g�f��;�|��>#�r�9�.�J�p�6����n}x8^��W���Y1+X�I-B���!L�o˖�|����+���v�X�kٲ͛9?&�m���R��,
�`�GG��TEI<��әX�� ��%C�X��fL�9;7x���H�n&"�����TԽe9j��:ǡ�BS�V*Q,;�͙�����֕�#�b+��-�rO6�,��! ���a�' �#�٘�SȠ�x1�S��t��(�kR�(�:�Y��q�:Z�����6�peq3N��/mLB�*6�b<f���0T*=�Ň9epf5�X��̗**;J��&q���s&#�X���c��SE{f5��0�N�J¼��EEEkR(�5���TX#�Rڈ�I�E�^5�-��3��#DY����a	�IHw�2�e�y+F�n�%2ة�m��UH�V�x��UjQP���֘���Z�e��TDt{�9��E3(�e2�+Xq!���%��^4�lI[Zs(�~�L@H�>c:�춑��g��i�$�}�a�#5B�@�(�LRa.p�=數��m��מI|�Zܧ)|�	W������H$�t�@�9���y ���N]��	6��s�	"�P-;�k��z������zl���h$��÷$A>�a�RH-��R�|��￧����������R��Kmlk*�`�ԗ&�#���h�W�l�T�i���~�!eH���Ok���K���ꯉ,$�HoO4��@��}�5�/���ᄐI|�����{� �H���W�>���Gy�i-���'Ur�%��IQC�y��B>�;����\�*��A>�G�#0�*b�|��g0�A"s��,��=��#eDt��{#BH$�O;�_�%�͆��7�
T(1&f����;�9E�l^��I%�ޠ�I$��V0�a$2cy���q�o�ԅr>�^�6$�^������0�7��n�s�m-ބ�z��ܮ�ĸ.g����`�}uu5��q��87�Mjz�����U}�@z��(�Ұم� J1g�Wg��Z	/�[+?T������ՙZNk�	 �]u�0�I,��p�J����g�uU~����"dB ���s�m�DB��b�x��.�jm0�i�7�^�X3�4�fJ�xx�n�4�D��� �_$�c��/gdp��y�N�ؠ	%�y\��,�����*D��[K��ҏ�G���U��7�)�vU
,�Ϣs��D���p�H��O�ݡ��Ǧƴ���X�9&fd��M�<�Ai"rV�?����-��v�v3n��:�cK%�\	�G�L��!%1I��k
m�5�a$�ͦd��B2;�4�I]��6{d�1�
��	yf�	 ���m.�����PbL�#wk)�6! IWo��s������7o�[2C�I'oe2�I�ʻ��:뻸n�uT�8	��cE�M�!�[-�=���c�xܽ��v�����؞w�2���1�r��pQ�U��1���8�>E~���@�I��8��wsr�5�{=��O]�����i����sȑj^xg���L�<�TCf*�pe����с�y;�v�=���Z� �(�m=��r�H�ϕ2���p�����\K�=�	�q�i��=�Z�һ�j3b�
�볎��X�\��+Ҳ<�X�A]*�k�+u �3R�%�����J�J֭U[p7&�gsc����m���C�&�q�[��-�;�8���r�E����Ͳl
)7h���m�����
��@�f&?"g������J7vh�X	/�{m)���� �(�Mfj��a��D����$埮�9�7@�7-���f0�	c"Mq�i������h$�Q��E��|�����^�D/m���z����'�DT�&dL(���Y�-��D׻hP��In�IY=�`��yw�?%��gu2�%*��i��#HS3$��}�%�}U�c�ra,�TP�Ē^�ɦ�	$�wk��AoW1g�2�J�$�~��K--Ϡ�D�����W��(��Wմ�/ ����_��_M{��XH���XmK�\�j�J��s��_'�����X%v6��]a��v쾲�������3��R6�E��e��^�~��j�faܲ��i$�U��(�K�����Uz�̻�o��$�gc�8t# �(��T?��w����G�N�.5)����l�9�Rxb��H+滪/��&T�S�����X�0>)=��m"���b���8���o�r�%�g��){&�
qr�LUW�]��|�����Q&��k��-
�[j��ѩ4���0�)+���ήq^��:C�׉C��&fJ��<c[�4�It�P�K"�G�]O&fl�	�wk�B��[\�4����Z��*I�
���r��noigexS����	g�A��	 �NH�	$�כ4DK��I�9�������7Ȥ��?%h����I%�4��/�}y�픐���d��_.���B3z�i.8��>=���YK"��i���a���%�Q�Zܤ�
GQ�we�H�h�Zk�OS�����^+����t;��$��i�J	(��d�m��=�N��c�Ʈ��h��Y�m!��
�
D	�3��WO���Mn��[�Є�W�튪i|�	/c��B�B�sz�%�|J�ҷg]0ڍ���4��aK��S+��s��-���ڦI$��1����/p��²V(�p���sߘ�䟔6 �F�����!Gzyy�������TG��rꤌ>[og�M��m�,�7�xy�{�w��77��a�E=0#@Nuߝ��[Kg\���4PIFw�e����x��32b
�������dϏ=�Rvi"z����$����2�i/����u�M(��=F�Iu�0�h���4IRȓ0���v崐	 �^u
#n}��k�+<g|L��
'��ѝ��I|�
�����ϗ���ן��=3�vno.Xn�f��ʎ��6�.1��ʃ��p-n�����Ι�h=���E�e~-�_%�4K�$���6�ԃ{��k��D���ݦXIpR� �Q&$AFa���g0�D؎���wN��A(���H�U��x4PK7g�(|�s�X݀���" L	�G�75�XH$�Uٴi|@%�+��U�1^j�^�J6��$�H[���K�C%L}f�p�]�^]�k�ջ�Ԯ��L$�I �ve
a$H.��7�N}���w>}lU�ԫ���W��ˡ�xn	������&x}d�՝���w�u�\/}��'B;%5���i;:j����뙭rc8�Lu�7Lk��
'�(��wt�*/��>��ʽ>�z}?A���W���~b�I�_��N'��xN��d�sE���#�5ݬQ,$�]\Xk_�7�:���Q�)J'�P�P��/C��ێ�r^]�ћ�L�mF�Q�[��ϙ�=��*A�f�˖�H$��͠�I%�]]<i�Y�{w�S�њWu�2�H�]���S��Ab)%�~J�L��9����s���z�3���	$����6_?�B��ŴPJ�3�6�z�>q�gC��3"d�f+��4�I%Փ���I/m����%휪��$�%��a��_$������`J���t�_�y���1����ĕ�Pm W�gM���"s����Zl����.��K�8�t(�Ӛ�>��"��U��ύ�Q��L%s�}if��5��u��i�G9�,�I}�L����d�;D��p�F�m)�j�()�a�H)b�ۢ����>�x��.ܼ2��<���y{)�]��������-˙5d狳��3�����R������'ww_~|>n�X;f^��]��G	L�3ێ`נ�ny���Ps�uuCu��Y�PW3G���0��[�Ee����v+�
�s;u� ���.V5	��k�px͎� L=]�p4E#�e�e�uݹ��}�7 ��.�9]��r�<Oe���r��&^:7eS�^�tǣ��nvAh���p�̂j۝6�8���֫t rX�N�l�,��4��f}�2n�mq��:z�=m�mt��x� ���לѻ~���T���g1�~�N?0�H$��d�M ��%�L������ns '>����d�a���4IRLȓ��}[�^�	/�'=W�a�~'x����I$�����H$�gu2I5Do����';b�U�S�s&A���c電	:͠-|�1��D���S5=��p�o�f��K��|�P��ZHp�G�И�$#0ѷ�Ao�����ܝ~	$���-|��(�ɢ�ߒ����$'���f�G��A��f`J0DDD	�*R����K`$�H%]�A��}Y�g���ׯ�n��v�g�$�����"PU��Q�������_��nG6̘���;-�f*6��!F(QݫSۤ�5��7\��wϾ�c��%�SW����~�_ J36j�q�%�ޡO���t����Y�����Kkvh��ւ`�D,H��n[�_���'�?��$��9�c��B.FV���p����_�����G�v�������Yޚ"�&ox~��y�x��x�Ż�8�N&u����N�ߞg�5Kio\y��[[f�߬�Z))�J�I�5�b�i	��P,�����"K�mQ-$����RU����\��^���];�E��I�9�HX]xfL�
fG�4.�u�U��[Y�#H�����@I �ٍ��I$�s���S�:�0��\�O��V)ѹS%L���&�۬0�J~�ӛL�ۅ?Nt�Gm��%t�ꆒ	הh������|����{޴X>�1e����
��-�d�u�\�k n:�དྷ1�vƱn������B��T���N��r�A'��$�[]����U�����6�ϣ���H���j���)�" L�P�]��e��7�w�O�%$�I��������m��k�����u�No�4����*!0� '��`4JK��LJK-o�p��W5	È>��o�uR��{&�t��Cޞ�.�c�z���Ӟ�׷����c�|w��˒]\;�k�M�oc�Nnz�[���N��������
�� H�G� :����I$�}�����Au~�i	��,��ʟ�D6��[�����;u	�����H���� �,��P&N��s~h$���HL��̙��
��������Y�įntڷ���A��߻����z�%���]_1D��ɍ� �A�zy�{��xڎ����Cj�łٚ�JFZW7-��7���;BK�YyV����Y*e)� �r��a��I%��L�A,��P�J}��,#�� 係w��$��Wc^n`Q�aDD	�*R�������i&}7;^����qӠ�H��!���$�I��p�A+~;=�..]����g>��D�0fC�.��2�K�WmA��K�釞�,i�]1co�K�|�NB�ϒ_^�iy%)*TB�� ���57"���0q�D�JI|6c9�	 �}�Ba��z���et�"�����[���.Mk��޹������VJ|��r3^���]�C�ɿ�����V��kԣ�<�ϐy�7��,b 8����5��ufE�@�&`J��DS]K�ؔ	$�����Q1����Ny�2Z[+�����"}��(���u�Ɋ�B�`�"aA�6\�جW�.*Ke�0�mkF�Tz�&��ڽ`��W���d(("g_�^�|h��[�� �	/���H��Z���u���V6�nWmC	����2"J�"�YzؠHP�k;{�n�66�eւ�I :c��H��}��v�~ߊF�Th���a�׸"2JQ`J�����Q+�fТ�_%u�UP�{�ÿ�'g�)K]����NT�"R�b��N]�ꕭ"7;���+��LBA$��e
a"P[]�Ohb2�IM\�L$�� L��H��nZW��$'	?_��0\�Ã�~ޭ�B�δ�D�[�����A/���0���-��$�'����5��Fi{/�׳�{6������s|��9��y��8�|�����>}�^l�Xy!6!��͢�`���Xo�\xr[����oo��[��ٸޮʒ��x�ߤ�f���||s�W��u��HVI|E��A�a��i!ѯg������'��k�o_gGNL��_z�z��'L㵒�y�3�b��%�oWji�P��Ѭ�*#�`�/�_���o)��u�_]&�]x�*^��NWVm������{{x�G3gLJmqG`����X���z��ʹ5%[��3H�Q0cїo�k��z�{�eo|�Y�7~��5z{W����<������1�]��{��?�����qn^�����u��{����60/`�Y~T�
�����B1X"�-/+q�HK�C4#%��$�xv�1�g��S��^�M-k|f�?ڼ~�A�&�v�!��e��v��-}��nb�-��{i�K��Gh�=�����B��Bpv�Lv��y"9
�wG��;ǋ����Ak�{��l���}�yY��޻2��R����΄���NG��=tP_��;������X�ɿ �ՃU{�n(s���!�����I����@��O��bz��Bx��v.�-��w��:���2	���A��,�f (�*Z]䤡�������w�b�WTу/z��{/�����n�6�Iz�W�^�پ�@�/��;٠��ϔ9���y!��^~��Ӿr��l�g�(n(��ٯ�B�Y����*V�:un��9�Ww��)�����4U[J��⡍j,�
�AC�mH�:>a<+	�֯������.Yc92l��p�V3r�ʼ@�D�H�G	�����NN��:)*���@���6l����jY��!�(���ř�Ƣ�Y�0:�c"1��
����e;�d��B0Q��N9�`sYx#��4E�H�e�ԗlԨ`�B��E�6
і�
2B����"YQd`,a��f�q:�	c� @̞N��keH� �Ԙ�P��3��#��4S*�c�0�2�]̍`V�*�Ҩ��1ED6�Lb$���b�*�MK��m�����c/KU��kR��Ԩ
1MJTmQ���ф� BH�,�� H
čY	 �) ! ���-KZ����p`��Y�P����g��5%G�p\UN%��Ucŵ�d$zY\@������l��ͺ����e�c���mLS��Q�SԪD��ә��m��9u���BG�[���7AR�����&ۆ׼�	���^������hgeŽ�3��uy�)\�c�72=�mVj��	�p��^�g�躧�z��qg<z�,��	��Du�ݢM�A]zα�T�#���8.��0i�e��u�:�]��,��ۤQ�x#I��0���͑����!�s�֮���vh3��o������n��Q�Vv�93�'��rn�9��βgnz��$.͸���zq����;��Ն�s�pn�N5�9��n�(CmH�
Ӱ�m������,i��Y�,1�n�&� ��a�Nl=&��t�f�^v�zx;=�O6���Z�q�{Avyl�:�O��u�϶\�ͻs�=�V�ᣬrܽ9��O5Au)co�PŚ�i4�6a5C͢��0�Ͷ��9�7��9��u��N�F�ѭ��$�\��6�C�B�h��MF��*��"�	!t�$�a݆������<�'��$�c�vq+�\Y�۪��k�^[r\��:�0dT���y.�:��Җ8��:umtv�e�s�ю黍�c��.�f^^�{g�xɥfDS]I�@��!��W]Q������2F�	�CR��e!��;K��\��&qo<�Z��[,tk�K�M�'9�t���e�0bb��GKVm5&���h�RZ�\E�r˕.�,�(�+�d�l[���g�2��8KIi@��={�v�WS�j����^�m���fÊ^vh��<�K���Z5�ڪ��ASh�3�IpT��U\ͬm��>�����v�<SM��5eΚW���Ҧ��<�7tX�L;���Ƿ4Y c�ݤ;��YmJ��q�u^K�)��=��]�h�%��Ǧ#����ucom2md�e��Yb�Y\e�b^a)���ѹٽ���6V����'PE$��ݮx.i����ݫ��f�<^�덑�j[��nF��d �$�1 ������M�����{���ٷl�@p���33�<Cr�b���OC^t�`HȦ�ife�!m�\9�h2�2F���.4�����W3 	0�1h�ۮ�L�,�Kq��!��Q��e���c=�K�q\C/���ݭ:��t��Q�M)]��G\m�KZ�M����܌m��s��كq=�(^��Gj�ػ-з��M<]����EM�h����c�\۷\�)��h�l���g������Ϳ���|�}��*�IU��m$�K����a!o���Q*���;>;��G�����a����\)R	��3�y&������ݎU��}�#"��H�J����H|����+�O�8�>��K�� ��-��Q%D�b���.��A$�͡M$�H�mwz���_�GވI%Y���ImwLb{���>šn���m�y�m��7ܜ-Yz_%�_�WW�6�1�HGW�wd�xn�$��m��i
��LDHE@�3	�Kr�L�@&7#��	�ڧ��{����K}��a$�[Y�6��%��4�@��V1h��s6��z`@2�bCJ�^�9�&u��P��!�^8y�'�mm��)zQ���JR&T�A��
u��I �n���_$�gO4���v��?)]r7L��
'�H��b��铸`�I��IP��N�9��z`������膢5�7sh���\¶��kvj<#�5C���m6�+��h7wW�fsdO�˰�8�o&x�箞��9ֹ觤 ��@�> ��;�C�i$J]�?}�UgO��/T�΍�u�m�>��b�R	S((2e�$�m
i ��Fӄ),�i�0�L��$�Iz���X����g�`$��߮y,�
C4-����q�n��ۃ�i$�}��k��IM��M$5��́T�"��E���z��0ׯ2!`�3�JM�������I*��D=�!�Zw��J�1��A%9�L���"O����9�Ws����$�EA	K��!��5��nr�˶�ά��A%�K�X��z���&�@�3`�ez���K�sf�i(�����%�B��q��q��ǌgeh��Bo:�i-x,i)H�S����5�a��J�^�������-$�HM�ӯ��BA$��D�{|:�=ܥ�&n�G �MY��L�2��^���$�IV�P`4�H��B�r:������ȷ�7rVDsF�c�1���5�霴��������gN:�6�)Kճ�}��}Wp�8�84��ٓ�]��y���1|w�O=U��#?m2M�$��>�΃(��S
A3J*=�j���!bwJ׮����I%��4��J����$��{���dS>$B��� =�}�}(���c~�	HbZ7��%%���c�]�;�<b|������Ii/�^�KI|���Z�1<H�B�3*A$�P�2�C�C��1�r6K��l5����3+n�����I�1�)�I�,���A"j�h6�I/��6Q�7u��VEB�q�t�H��w�a�7�A3�R&L�p�\���K8lm���;���zi��A*���A%�A���K"�j�g���%s�7�Hv,a0�L����']�P	=�4�"s��RG���S���I|�
����I%�z[S'��TL�fd(@S
w�-��|�8	/�}b�0�I���-��(NwS6k^Ǚ�������p���\��x�)�Y�N��K�\&�w��u���Pt��LU`�бd�?N���e��<�K�Ls1_@��(����׫f��rm��;��&$)Q���Pߒi���_%9�4Nƶ2���$��c�I����iNwM��c��������AK����&fl�Q��C�^ݞ[��v���`8�5&��H٘��������d�fd�1�#��4�H�>�,��Js��i)�x�σ��,�RU�\i��)zt0�_,X���R�Ĥ߾+�-��B^�����(��7!���ÿ4�I$��2INwS$���܉��goT�|���)��
�2f�Վ��B	V�M?�I$����+��I�a�C��J���$�?k�cI1"e(P<�R��t]�q�U3�v�KU��%��IOoS,�H*ܮ=��zm�:�Q�-<�52s>�(IR&ua����I�'�Na/����wg����K��Ci7�4Ia%����b���Edr�,4���(BF}��9WK�;����h9�N�:��:w(^il����^폆�>0���Y�TJ�Jy��FQ�(Ґ`������ � ���!��tL�]�M���ݶ+4��	��v�͕ĶX��t�Ե��+C��,!1���qm�g��r�D�.�<�ŇҚ,K1��;X������b�;D V7\�^�<;q�6�ia�a(F�p ��ѕ�K�S{,DN�k�aЊfږ�*dsV�h����i�E�k��z 8�<�qHV��5u�X�UַF�-�E�1��&\u�[W�wV9���Y6�ێq�A�7�l�k=��t���2�\�Kw�߿��]��YQ�ɥW���\�Q��M$�*�+�iܲ'�=�׾N=އ�E|��n���HV���  H ��30������1�<���H$���Ii/�nW�h��,�C��ꧏ���;��QT����{�]k���"RU�:h���$�oY��;���I$��4I��Ys��${2�
f��L��ᥫ�3�y���H��sM$D׶x�	$����s��[�0��5�S-%É4�$J����s�l4�I%������^�q'wPHL���ZIWw0�)%����Qޞ�?/��;��P�Y�[	w8�L�k���լu��%[�9��r.u3���0�ܴ������>L;��V�Ki��ݠ�A$_twz*{7-�͌�����H$�U��6�Oz�LH�Q���Q�x$�u����V2�D�hB�?������L/]���9�h�Yt��!�J�[��z-��\&�y�Ꞟт,?xX�g��#����3���o�5��eC�c�y���d�*�ߘm$����m��5�=uq��&��j�"A30��M0���Qa"yf��A$�Jˋ�M������G�Q�ޠ������a��w��2�%#0��碫'��=�G9�	 ���4z!"U�u����BBw��׉���W�5;�#U���_VnR%L��T�1�-^x夒S�LB~����&kݬ����a��I$E���A)͎��Ӽ���|���2�@*&@_A��˛�l;�:�aZ��f!�`��֮&�-����$ĉᜧ=�(��A/,���I%��0��6��D�U���`������'�~�!8��M�Pԑ՚��~�sb	�W��:��}z��$�_\_zq����I/	�S���	��?��\�_���o�sQ�/�����Z	9Ѵ�%�H$�9Šn��~�5s���B&��^��=04�&�������f��a���9wh�����Nlzqm������"����� ?� }?x����	$���m����H�2Vz%	��aR���9���w9��?f�I�fz(���t�M"R��b��`_Ά#� �:�(��|�31)�g����[��`BI �v��M,�5]���'~�e8l$�I	��i������z������3�{��}GZS9�MZrj�\9�M�/^��ݦf�lm�j2��5����Қ2$L�l��E�)̍��$�(V�0�]��%s��q^p�E$��u��h�4�$)�C�O{�?�A(�2(���L��h�X�k9�%����8���Ɣ$;G�F��U����&&%D��ڜ�sb� �Uy��$��X���F��d����$�J�g�i J����'�q&%1���P٣��k���}]�S}@�S�A�A W�<��:�"��\ȏ5�P�����"�h�99��y��f芕��*�'Y^w���)�x,�S�<��p���}�	�/;�3m�[�=uu��#��N3�~���+n�$�$�ٷ���?R@�;����L)Pʹ�����L/���t'���'��3��zb�zO��$*eJ�LF�0���
���[���G�\�tt��/�ܴ�lߏ��<�12��g�&��	$���� ��_E U�-���+�3�I��nY���ߩj��ݷ}�^��>�����Wu���$�k/=Lyk�H=`��{��v����R:I��"�1��d����$M�����m�P�랰A5��0����O��l����D�Z���7�>·۠�\;�$�V�(9�Ԫ��ֵLT�9d=ٴ�}5��&%1���Q�|gS�I���!�����1e���m�O��C��L�_1��q d�A�� x�����ª�Y��mV��K#j��hl6��-�����fx�w4g��.�wFK�o2�3�����7'q����[�a$nais?d?bBA�q4J���L̳��8�<����q\�ԡ��aG:�V�]/d�q]�I0�X.���Ӧ�2���xt�cf�2�ib�X�t"k.��E�z�j�kSv�<ن�� ���d��_W/���(�z�E��,=l�я3����&���U롮`��Օf�f5�PZ\���mv)�a\�5�X��ݔ�n;+����6�v���Q|jMlܬ�s�a��rꐍE.%q��t�m���%��~�����*R ̙!-�q���?��Wē����7}���!�w�Mֿ���s�P$;>����fB�&]�mV F�*�|=۷U�k��d��O� A�|��luҜ�����l��f&I2I31t,�����%�x&��1�a��g�'�����?Vu�`����	�@��%L=�꬏Z�ӱ
+��`�]�I?S��� �[��9v:4����j��̓p�̈��&[�|��j����=G0�:��,��W��� ��V�7�����J'j}V'�A�����bBQ%-Zח[6��lLVa�����;qsv8��֮�}|��rcL	��i<�^��'���;̓{�+��E���������ΦO�4n,B��$$�6�� �M��;sF�J���b�"��1G�{my�B��������^әZ#Aء�%��7�*i��qآ.��%R3+'n/76�ĄSG�'��(�3��1C;��5����?[��<(oO�(F�_���x% ę�`@��ݪ	�w��'#���iǸ�?.�$�k��O�֌��&B�f!�ӑj��ofW`�Sv�O��w�`��\�˫>�z��o(�<�~�z*@&&IJA,3ݿ� ��O���7��V�hp*X5�S��@5{�a���O�_i��b%�Ij�(��)0�#pMt��˻=d;v��fM٦�7X5��]n���ƫw����Z�L���&{�g��������	$r��D�xT]����l��5��l�޹����`D�l+_P�bE�.�"��MW�Q���5��l�O���O��4g�d�Qk�:�t3鶷$��J�$%�w���$t��M������[| �(�'��ō�p�=��ކ��z/B ��P:�������)��.�z@��8'7��2��)ڻ�뫧"}5���y{R���{O[nt�c^�]�����)9�Z������{��<��{B/t�ǔ~2	�h��<��\;:*Iz��n�\ًû������������5���z��c��P�z��3�~�{ڊ����[�w�Ui����*��p�̾���q7�M=�gH��X��o��y��q@L9����=��"h���3�6�h=v�^�����Z��f��W��_ˀ�L)�;}}�_���������~����-\��v�75B�}��#���u-���C9��������InDX�g�oȃ�{�^]���=p��<Dii/_j���A���<�˔,H�x�σ <��=VT���`��{�'/?m��K��dDM�=Rɳ����,2`�1��k7�c쏓��?�v_������Lw��м=�U{�5�������^;ݻC�3�qr�5��y������$M}�������s���gT�^<vb"��7twI�Jۋ�.3�T�"A��W�Rx�,�=ML�	������X�ޖ�A����П���t���&`�����'(@�2S���~�������$J���J5S�.<��<�Ƥ�˝[+�|��}���pC2w�	�qzq�'pD}�QܺΏp{<�B��{e���ɉ��^8d��lv��+�{�ol�p8|(\@�}�����P�B����=}I�������x����}�:ſg��|Ls3$\B�㻥�A	JAz�o@$ ���X�A!H������e��9?'8��F�`�9�1�&�`ǩC���T�J���E+r�T�e�Gr3&�NNǁ�:�ee�b�X�n\ʩ�
ʅ����H�D%|��|y��ς��YQ���D�lsjqD�	1*���a�b$�uJD��H	 �!
���L.�-��TLۈ1X��\$2����@�1d	3uG�-�̶AQe`�<�*)�G���.t�" [l�H�R�E��0	<)�8��\�`�UC�G���(w"v,.iu��)��AH��-��	6�Y��N��{�$��B�� [hr� �lk9�+ȉ# ��
"*�JJL$��)���HBXq���Y����Xu^� ��%Z�.&V���Kd-�KI3= r�H�,��'�A���`�I���_���bL�0 M\��_��s҂=g�A��m��4	���z����p�I���{+R��DȘ�10�{��ă���<���5���>�'�'��[�7�5� ��;���{����GZ���@�!?f�&K�J��3m,��vz<xy��n�1���3��@&&IS��eU���I�٢#;��*�{;a�=^�	 ���|	�1!DH�-��w�����=�q5"W�,�Lղ~��MNQ����$�/}�{	mb���&z�e)&L}0"T6�4���LgnS$���y�-���z#��ϳAϊ�:k�I��a�Ԯ䘕J�$$ٷ��dgDo=�\�v���� �yϐ�����uU{f���P�Qŏ�w����:���ٮC�=	��g�w���E(����o��k9�S��h�|����A��{ڮ��O�7u���"F �P��f���t[�8�3T	���Հ�k������Ͱ��:��P'�O�e��%|�����q&���?|������ �":a�٭���	��g�2�mwhH�؂P��Q�ѭ�@=�����pk"baw�WTI1��A�	5�Θ97z�S�����u H�ws��t4��2eLA,3ݰ�^�%	FP�B;�π�A����%�^�z����{�w^r=�pҢd%"DKX�ՂA{ͰA�zɶ��u�$�ͧ����s=w2��&>�*)�5��s�S*�#�����@�H���;�1��Y=�0HU����܃��L}	����6I"{v�ϝ��QY���B#�ֶ?z����+w���|v�N!3�َ�S�6��<Z�O���d�;��+�=�ҋX�r�>w�=�R愿~��ڴn���.��4�����L��H��	�$��g��}���ʘ]��v-���/��5��-s��w�����n�
v:8�Q�^�6n.b�3a�q��d�`d(�;�"���]�܂r��<-mۆ�s��iz�U�;qۮۧ�=���>��k����:lO��WG!zcZ��v�Xmա,j�B]c��Aͦ�]k#*<��6������L<�*��rk1��L�Y���;��Ғ�76�#U��m�s�k�h��5��.�3]���qQ��em���?O蔃2&`B�?���{k��XD�ފ���̆w��uF�O�[��Egsa���bR�@-X�is߾�{��Ψ�����u��~&�y�O��;ʁ �t��2��˩���6͏-Pb�%*	���n�?��o*$�դG��=�<&���`�'�yQ""��eDIJ$D���o_�G�&Bv�3A �s��gcyQ%����7���mu�;5�&{.e)T|���l�-ځ���ߣ{��:��[��y�ª�����$/F�H'�;o�ǟ�_|��eVx��n���n��{Y�ƼP�b&�G*D#�0J�wL	A|���]�"��fWЫ�>�0�3�H�I��u3�~8{�.�����0A3{8h2��a)dL��[�~>�_i���]nR3���nx���K}��z��r�-�����=�s��c�z3�h���L���b}7�\�{羋5�a�S��P	���ͺ�Nti��?�z�~l7>��������ԢfDI�&f`��]"	>���?���!��7�A*r�&++y���V���1)A43�Oo�}��!f�FOG�"A��[͂A?��p*���/�׳Ɖ�aX��J*$).:^ՒH5y�F`z�H#�T�l��4C꽠�?��<�dm��`��x���>��5�i���0���+p@7	�mt�틙�׏'��0FO�X�{���e�͉�k��}|��w�C�+q�ӯ��.��~=Z��
rS���$����d�����u�H���g����R }nX��أd�M�o6I&�;(3s>�NM�3�:+x�'8�����bTD	o��� �$Wn�	��C풉g�2ݨf���Jsqv�w�{�S���ϵK�2�v�>�Lw��U[��H9,�w�y0i��WA��!��&�bR�#>�þ(F*<�<��BO;�~��&}o��k=w���*B�3
�쨸z�ٱ�w�G����m�|A$U��d�OV����MхE^ω[���3�WAJ%LD��f:��������O��¼�D����0OƳ�`���ƌ`��NW"ٹ���}J9c�����.��<�f�W=��oN�z���k��\va%Q%A�{���(�THR"{��{�I����[h���ȭ5�^0dU�d�~5�������JA3 �Pf ��u"���<�L�5{P��{R�oĂ@����$}�nK�V]��lz�y�3:��'��;�_DI�L���V��v�i^�wD༊�4cmNe��� ��c�0@'r����'��3 Ĩ�������;:�b��w�Oz�$��Q��$<�s���`Sp	����)U��<�{�B���!<�;�}��!�w_��f�/9�?���
�s<���y0;�����渀������<�+�.�O�,`)=�ߜ��N�g�^j�cqd)�0����Y�=����uz=&ϰ�^����m�H=�h�	y����3ev�Evz��x+B:%%)�` "d��u=��:�K/cNT�b!��:�ƭ-��׹��2&$�#þ1m�`�v�6�D�KξlN�5~UV�'�LEu���N�����8}�̤�B��}/��	>��}�k��lT]{�~�ʌ4	��o63*�XW��A�nz���zd��eA�lۨ��q��2A'�ǹz��Vu��d�	��@	�se�}dI�"̯�P��s�;�Wp���ѱ�D�u�c�nd�ɍ��I����\ѠOqxO��f	�1Kcr��I �f�M�a�n�ƶ/xw��~'�w[=ۏ�չҒ��hc��S�}W:*��nH�͡��z��U��x���u�����F���͔8��VR�����`�����0�a:�-�n;�˳36�p�]bw:ǣ��>��Ӵ�[0�.`Z@���&���=g��f瑍G5�ak��%�W9��.u����֚�5۷V-S��LT���ym��Ӽ��Ί��{6y�;m�y�0�WR8�u���W����R5ҳYj�
���˱ChK��F�n�0-�h��/���J&�5�mE�F�j�$P�6P:�5�酋���.�luꋧlN��rek��s���_���M&T�0bf~1�}�A=ͯ�����l�9�j��Y�a�t9�@�q��&3L(R���1��c���9o�+:�G��l<�~'���l�L�m�|��ۉ���������$
�>8&J��`L����� ���l��ݸK<��V���H�k�:�$�v�����S�������F�D����z����3���$�nS�O����cj�Nydf��fݶO�%搥L32����w��9�6�^��`��yB�a|��޶ ���s�8���~od�p6��8�E)k����B�6�G.+�u�A������l�i���~�!��Vb��x�$�;�o��Ă~ͩ�=���u�\�K�Gw띿6O��g���}�3&b�*f0zn.�|:��r���m�����#���x���-��i=����O��Y��a�����[�������A�/b�~��󚥂��:��>���|���(�~|��ފ��o��$�O��Uy��d��[���>�k8�(L���|sz�d���{�����u<�H$���|�jx�$M�]��"T)����ϺqG���O^�\�[�� ��sƁ ���9�[<p��2@3�|É���0)�*���F� ���v�3��׶��rs��F�F@y�L�&�?OW/�&��Lb�4�&ji�KĶf
k��ǐ�v�X^^U�w�����A�1(I[��H�U�� �/7�*�Ù27�Q}5m�H��r�_���dJ�%�{�������q��9��_D�g�	��(�H��͒o7f/�+�LUu�:�G�kELɘ��B����]	3�Χ�X�F
�����0�.�t݄ر��12Z�6����}��ຮ���0�/C�׹j)*�[-��o+��a���wYX.>S�q��1#�ַ�^�I	�z�$��׭h�:�(�(L�����ʌ������~�g��&v�(0	��v�[� g{'����%p┉P��3-�����	����focŨr	=�S_D��6HV��f�OB�g�.�<��	0Lē*Z�=s�	�Y�XC�뺐��̝��ؘ!vuk���_>H�?D�0���C��ψ����	������x^��C$۞�@���6O�%��eLD	�BJl}�� ���#2�{��D�f�k{m�~7���l�=�!���lx&D"�B�����ƻ6�A�]��܎��'�Dﳟ�[�o�@���S"&R!D�t_�~g���Wd�ǻ�� �Mve�	#v�^A�o�?�q�Μ�u!<W������hˎ�v!�6�l� �/=�.#P�(nXN�������T�}��@'�Y�<^����s��(�xVB���>����?|~ ��Hϭ�1��
 �&d(E����g�~#�_����څ|���ϧ-�A�r���]4!���8|��T���jj�Gn�����lz�e�1݉�c3[q���m�Ģ�e݅�
��b&S=�^�6A���S��;k�R�+!7��+�$~����?��ˑ*~��`�	^�k��Y�8��������:�O�Y���|�#V������-����DKUq�����J��LJS`}��q���I'm���n+O��W����ks������r��$ȄT�B[��oo}V��ω{�t�7j�P'�~���O<ߒ���Tf�{,��z���`���R!D�l�������f;���n���:���m�~9j�W҆-����	�SJrs�/�G�_*��W~���(�����}�Øg�^��!��X}�f�Z�@������:��������痨�W��g��Z��I����K�=k����-Kw{��9�o����)> n�I�w]�����u:�����h�7�����T��LM�1��I6��9DUQ�I�a��������6�f���w�ĩU�J�R1�^C,xȜ�ȪA�XTm+l(M�0yh<i����}3��#g�N��E�W����q/$�{"R{q$�{��߽ϐܾ{��m��m�!xl��za]۰=���^sA.#է؜�/p��M�_�7�u\[]��z���wX���QP�}븪'�$�ö������oohM\�\@%���4����үjX������aO]�R�w]Zi,'���v0G�;��l��a8��N�������/L���3�&��;2�A����!�/:�uD����e���{���}��9�{}�9%�i6�C~3��j������H�I,.����D[{y��1ڽ�˔�������l�횵Nt{��my�N�&�N�Ǌ��p���7���źNl��=�Y�����{Z�c���m���;c
�w����������}�eA�|�T�;h��}������<��)43�)��3�޸�iY��C�޳����_G���M��=#�S����=ފ�G��dy���Y*���Fk�}���w��|g�S甼��0�i{;���͗G��`ķ�����]�W���Q�m嫭É�÷�Gȝ^�H���6X!�˄N �b��l����R�T����n�(fM�g'��c<����<�0�{+Z��P�Փh�8딉�N�������&��0��f�N�5Y�
��2"pǼT�yT����� Ik����Ʋ���$��E�,% q��Hր�H��K�*�z$����i�+H	 $E$����	^� ;J���$	�ϋx��W�-�g����"��)V"4��4d�)\��Ķڍ��(�EE^%�<��J�xS��T�u�HJ�f�1XC�����$_7X$�KH�&%,�K_$�0���( 0��"')8� pU��Hu�.d�D"�<6�d�]��9b�$!�	`kԨ� `E"<�L����x2��/�@,
u�Am),�F���"��r�D!8�j�g����n>U�%����љ�xܱ�f�Xxu�."�\�w]F���;B�l �-�hB��X��=Yytr���We^l���ɧ`]�7Jō���l���η.ɫ.��}�]h�m��m�Kk��b�T����:���?���|ʽ�q(�8��5a�q�1�.V��6�����*bc�C��]���2�VöH¥�G���4��]E���p��1�.� ,���Щ5H�G4pk���9�c�u�]��O�r+=�Ů������<�p7\�[��84i���,C�.�e��A3	�&`\,؝^���7��x���$�&�=�d�m����r��zl:���8�5�x��e^�/�0Y݇[����)+��%�j���:��j�#[�9\5�p���=ODoR��#l�B�f�V�����n��Հ�p�(����`C��M�ܝ�W��^�a�nq��`�����vmlm�\q�Wa�^C�������p�۶4r����g{]�J^�5�i���M�C��V���k	u���ט�.)6�Ћx�i�p��n&�e#�h5+)aY�e+\:���I�'=������2����t�ܲ���%��{>|�UPIv#Y��A���.��=��Ź�+���gt�{�P�]Z�me���l2��Sk��&�����4��W/�O#��\��',�9c���b�;m Y	�X�Pe��Λ�X�p��!�n�zwN�k^2�<��)�v��Ʒ8�	^���B��'	�<�<�rd%�&�	����F���	�o�����=G�����r�8�t�[)XB��\��"r�����T;n݊N�1�[�Qcq���#WdX���%vݲR��6���!�<h���^R�W���f�m�ogX�oU԰t[������F�f��S���uõF��'QC�Tv���|鵮[��]�l�-ˬ��m句�_�߸�ӽ�C�}흅��<���֒�k��6#�>�ݸډ�9s����n�t�-���$��l[*خ���8#uZ�+��&��VsΗ�YP̶6�1Ɋgs�p۳nu]��uh�t Yh�y����޾*�RMs�o]���}�A�����V�])s Y]2M
��yp]����S�22�����/c�<��Zq�YV�lj8�]�}�X	��\(��M`��im3�f8��@��ƨK�Y�)�]�|����D�3�?���o��_�؞�.�����p�����#ޞ�Uwu�{b�W��X^ߔL�0��l-����/7,�(Q#3�U���>�Z��ggy��͙8��`ǽ���O�]ȕ?D�0f�+T�� ���d�A�U��*���z� �"�P$9���~���*ġ%S�m�v]n��5|�|H���#�5ݯ#I��D��3�Lҿ*;~����3
 M[���I5ٶ�qG�z��S'�	��T?N�sd�Eom�����O�ϵ� �'6v���]�S�HV��!���`6C�,�s�[v�����Uҷc��{�n�O�v�i�OĀMom�[�����s����I N]�pz��"dDL�)�9�l��:���T�P%^qB���|{��a��,k�Y���� A���QԁI2��|;B^�kM�س=W�D���я)SYvo� w� ����'��I�vk`���������^f��C�Edyh3tg�&L(����]/�`j�m��?XqVs�k���P���ȉ�0DLB`Jl�UǺ�'�ft��$��S$	�ζ��3��$E͉]�zHަ�r%ބ%JP%2Sf�z�d��j6�xY���U�$:���'�϶���<��3,ܣbI\�Xx1��<A�n���[�J�ۛ�C�t�s�r��3DDO���Ʉa�'���ka�	:�m�A ��Fbw�&�OoO�^||H9��a��y��B*D(�4�r���.��J+�'J�J�δ�H'�w���FtW*$�wK�����ρ#�>�JDȈ�,<�u{��A�]C�$|:~�m�9g��ôZ�U�9�T�����]n��^�4�FƘ!&�ު�p�{�>����6���i�rg�7:��X�������LX�C^u���C�矮��03���_*3�;�D(��ĳ�]MT�N��Ψ���� �����{jx�&���3�O-���	'�[�ˏ�"$D0%P�1�>@�j����{��|f�ֻt�9�:E H���N�=|�❧������O[6����Kg�낼�i�l�=������I3q]~��=����d�%W��`2FmF�D��'ާ����s�t��n'u�IΩ�@���&�f@���Ͳs䣦�a0n=�ݾ�hd�O޺�?Sv��"�x�Z�7맻�?o�32J�T�Q2[1�h�ko:�$�LzP��J:k<Iݨ�D�O�~�l�؅"d(�($h0z[Ã�_u��߻�p�M{�}�0�l!�*�����(�j�e�T���1Ѣ��Z�S�m�,���C��/o}W2��8�6Zf�D�
�D�:�Y�#���������U�&Nz��!)���G��a���m���to��r�z}��#_�Ɖ�{h0G>۠2rϷ(���lBb7�]�nn0�r��)]L�(i��������x4��]�����mItok3��{���(M^�� ��<�n�1���t�o�������D�'�~����"C�l(ʁ(��5}�a���G�݆�'5s52�!�kۼ�'�]�m����ӳ�{�nz�x±�D�0L���o�3ٶ� ���]��z�<pi�u��=�{����*R!D���z��w޿W���nS �g;.� ���1>Wz8�~����铂+#"d(�($_˪����0�����q~�$�4��$���a�Hͩ�Fs�2�8J>}�%;�5Si>�i��0=YY{Y^�VD��{")G��i�'�6%�Bcj�y�y14�]r^�o<�<�x��]n<[�b�o��b�� >O0�.�5�u�&�tl��ݫs~�+�/�e�n'��N'q��mֹ.�VȰs�F�]a�&���z�$k֗�a�N�s�f�� /[W32gIK�%t�5��\��壡�Z��@�]'a�����;p�!^۲�nZa�8}Wg��ڳ��0d����
�6�@B�I��^4-�6�H�5ׅ]S=������ZY��FQ�r!u�T�M��hjLnn6�ǧ��QmR�.�؈k�K����?�n��n���~y�b�m��Ē7yԚ�F��F
����lA������MvFB��}0%{��E�Ȁg�y~��q�ޮ �#پl�~Ω�Dy1K][��z����A2��)�%[ݿ|���s�2�D]>��r�ދ�� ��� ��4N[|I
I�f�.�n��gfy�W���0� ��S����Ƿ��-��.�i��8~'���ȯw2fd%T�Q2[��\Y�	����?��똎�ްH˫��z�p� �����/v�����3�/~�웑�ݨͣ���'�!�b��%��x��/6��&X�j��L�0%�-�l��F� �{y�H��~�Yb)���^6�?oT�P���H��b&���l�����rn&\Ϫ-��E{��8aԹ�[+��1=ZO��/��n��z����4�{O7�sޚ���P�4�����sS6mK� �� �@��fw٬F�W*$�_����Sq�w����w��EE{��b )
>��{����+���$����3[*;�9�#��Q���G�"�~�A�J0e6�z��OK<r��	-m�J$�����댞�~��3�������	Zv<�FQ&�-�}����;�׃�����?h�ܚ �O���l����?m:S#�Tz��Ԧ�5� �Lut�������^�V!��:�!Wv�7l��wϾ�|�55+v?~���B�w�L	���y��S�8u�)�M c�ۜ�/�Z�L�f�Q����ɫ"������ტ��~�{��A?��6���&��g��Q�OK�vAߒ�3 �D��+['�F*Ο?���{��sa@���Ү��O��`�^�E��fm��N�8�h�&�h�Gk�$r
��B�/�K���,��9���?��߉���bs���Nz��`�A���l��HQ�����o��v6�:��bk٤���H$~���d�]:��r�J}IP�|Nw��p{ LH* Jb�u���FumR��;���+}L�	�׻���Q'5���oF_߽ߞg���y��o�l+�aG\D��D-<���3Չ۶����	��X�[Z�Y�篍�A?@�J�o����x�Ͷ�N�t����#�7��r��W�^�` |w�����3(�FDD)����t(�".�o�D��ֶ�	 �E{��Ig+j~�����F��y{ӖH��IJL�$�E����đ�]"�76��)�޿g�'>I�m�	 �ɠMC�=�%DKamW5#.��J�2��Dvn�$}[4H5�}]Su�u!��H�gǻc������B�#���w���g��Ԇ�6��UM`�w��K��S3�#<�`���^ž��Yb7aI�&KS��k��M|?g�H�?��>{ަo�r�b )
>���箏��W�v�ǳ.�MxY����/�=��r��A������٘�>�Z��f�1�3m�e�K��BZ�I�m0�̈́a&��sip��w�ǿ�441t
cx���g�0�m|$�H�|��f�b�&=�c�z�0~:n�+�r�Tz	D��&�-߻[dXO��K�Fg�]��Iŵ�_	�|��|�y����j;n:�����?���I����O�;��$k/:��X}�h��S���O�WE��\���%��	I��QE/|���!e!���OǏO�� �~����� �v�Ԇ
���Һ�(UY���1"TD���l�H5��7^��y.Ul9Kq@�k�x� ���o�����+;����4��1
�}����v"���l�Zߩ�Y����n�S6{������wۋ7��Y�h�U��o��μ���\�%���>��N��:7E�wu��)��#7�6�Ma���[�,���ny�3Ѧ^-j�M�#��/fhݑ:�d�U�=��y�.w]��Q�8Φ^W[��<>N�,�*��
۱�99���붼
z'�^#F	]���w%���3mtYv���\����ɛ5r�&��5�p$<�����ǜY<���ֺfv`�]U^ָ�:x՜6c�&�U6��KN,�E�e��渼�k�A�R�C�������R}0%w�t��(j�v�$�]��`�7"��ya":����7�A"�o[���dJ$��1B��d�f��e�3�4�. �?U����ow�3�5��vk��7�W�0�&~�&Ͻa;��$�k�|�?W{(�\���\x�H����1�B���ϧ�D1
Q�dDB�/���w�: bk4~;{�A�H��t�$���Z���dG��䒲�'�����2���1�x���� z=���_.���$�o���|�-�>���hW�>�0��J�&� �Y���O=���Gf���)�=��d8X���}}�4#&f$J���sZ���	��7�@����|h=���;�~y^��	���
1��ɘ�G�SgO��Ni=݆�,���;ո�T�\z���W��=��BH������s7�QdOMge(Mϰ]���W|0{�kY����E�]+��R�1���~'����$�~ۚ$���� H�kL>�s����w������R%	�LB���{]�$��Q����'u���	3rE>9���z���L�L(2�g����{�U��,�^VMH��-�|�A{��n�����I�����!HPL��S&��$os���KN�#;�1�U|I ߱�Io;�-��Dj��Ώ:���" V�& �4��!���3hhl�^hcǇ��i�8`�"]��}�ØR�"`J!-y�@���TA�u�*w��+�OO��|Aͷ!K68#&f&J�5aGW6H*�To�P�}t�hܩ�Ğ�sD�O����I�o��s�Ց�1&
����>������`����������IM?s2���c�~�R�V��ʄ�q��>�F^��nyk��#�f|'���mC
����������S��'n�P��2�����r]�û�o��`�-�,��o�{ku�����$,��`��9��s����^p�1��Ü�>F��E�)��ϭ��>���{}�?/�hP郏+`��gW܆�]ٲ��b��&����_s�vOW��s������2\��yg]|4��:o���X����j���c��[ӗQD�ۼ���͊���ոkZ�t}���k��wR�5�g�W<�����?bu�M��^���~�u�^O-G��o�^�i�.�G��/��`�����:�%m�}�k��7]�vw�N��Q{<o���U��mS)~n�zowD���?xb֕{ �����:B(�.���g�b����r��b��<���;��-?1U����[�,�[������3�����fw�=��q]��)C����a+��.4F��|����B��n�uׁi�ɝ|͚���~!���I�=XX�nwW� �;����
a��[�)����y.��/��<�!�����z���u[B��r{���kV��}�H�a�Ed�;b�Œ|���|r�y�����c|��=~�ʹ�c��0��<��Pż=}-��;����7��~����vq^4�Z{{CZ%���Gs�y8��;��@]+��<}�>������O�^��!h��vN�w&��`��m9:�F���Fɻ�4��3)#�3����!�G����?�"�8�=��D�Յ�X�bK#q!	���<� X�f0�� 6�LpW/�%�6rvi1��S �U���i
,8 �XVU�
Ӟ 3��αȀpc���2rrvi^0F�\�psQ�`����U#�,�$�"c�5IY�(�XpW�K^�ԦR�˃�U�31�K�Q-J�J��X�h��H��Qۀ§���Lɐ�Q�l-,%�I��ز�F-1&�AXJKS�a��U���Ĭz�� HZ�j2!����^&Qb��i�v�R$�|x�xA	NC��leHdX1SrR�`�y�P�eihڼ�O�*�,H^��Ea���@��uX��.����j
����*�V�@T�Ӡ@VDB��N�y�X�d���bx����g�q��@��8�[!�ټKǋ�UG�iY�Ѯ$ �z+�3Vc1 pN!c$a-��#^k��C��k��֒����lWd�� ʉ��^���D��v
9{����� �ܷr#��}�Z��P$O]�S	"	%7y����ٷU�s����������QD�I��l�F�]TЕg�,�g�"���cذ�m4l�l,��F�fĚV�	�)3�m j��B�����D�ȅ
$hGՑ�j�6���A�˪46 ��ַ�"�:(ӻ�a|�
C4(�"dJ ���U3"��1f��P���&�2H�Y}��H�v�>Y]���b�oj��.4{�����31)mFV�O���۪ �;��1��ɭ#�ӄ{�64O�y��$���Tc��s1&"!	BS`��v{g�]~���8H;9�A�Oǻ.h�����KcnL���*>��$�s���eı��'5c}�ih��z�M3q�������ts��f0o��8o�W?W��y�Sb�;�  ��������1��2H� ʉ�{�?�:�M����eu'�o�ks�w��~���I�]Ǔw��~$�(/�nlk���	�,���r�&�
Tj)��Lݞ^�ܫ~����N�r#n�ݿ6$����D�Oض�(��N��":�{v�Mn6	$�w��ȿ�����P�G��Y�`9��`J'i=�Z�h$��s�D�|��L�a7�^"�����)ȅ
`Ș ��:�� ��]_A#z7U�c�m�t��ٮ~�}ʾ*��%���R)�]=T�>}�e:�q���|���A#v+��C�_W�h�*�I��U��ɘ���	BS`�uA�y��3�m���#s��WG������;jx�$G=�l�⍩'u>g}��ؙ���(@��jd{.�����W>ݜ.�Ĥ�}������U�tSxVw8��������u��������p������G4�k���<�����u#���+JE-�h���b�	��b��nn#4y�Nvۣu�[��\/I��:-CM*�4΁���tH�df�cl�uj��5�f u�#46����n֬v�,�e��.A�����̥�ܡ���4�B�f���%f�%ں�ٮSKm�$m�ȩ	&�ܯ�i�c뛲Z'[V���.�g���n��Xf��bܶf�&�=p^.ΚS�2�q]��������"`�*&+�}�����+�@$�}|ٟF�DҺ2�����~��_��R���1)��o�!FZ���/Lȸ���$��jt�$���w�Eq�'K��M�����11" �D�'��I���d�J~�Kz�0x�Sf��}|�">٢���B�2&+����Ԃk���N��*�2�D���mcd�OǻY���p��~~�f�'�^7��33
B�-��U͂E|��|��v���HS��E�ύ	��	��s��N�׵�n]��ddZ$�BT�Ą�b�z��	�ƅN\�R�<o�7Ĥ�),5��}{�~��D���&���Q��'�S1�@���T|������N�Cg���W��ה�5#�eJ�d�2�L�g��^�5�[��§��e��9pe�/���n:5�n���f>Լ��ݿI�i?CV�tR��A��a��Ҳ�aH���p�_��eר�����?9�k`�~?�k�@���F��1�vh���|L�0T�7�� _�|z5�/�8�r�1����$g�����	wk������ Ȃ�${ǽ���3�=48MG�I���?�.�#�55�$�w+�=�c}��"y���}��χ}y����N�%a_2�g&>����h�;��h�[��,�H������@�O���h��3�*�4��,AD�ۅ�ٗ��@��7q���nv�1u����Gn�������)S���o�>�u�	 �WMf�3�5|q��� �o�TO+��Q)DD	�*�#}]TA��~�Y�U�I$��uDn{���uV�K�.6lz�yٙ&�
R��#�����s�TI/�Y�y:\�Im�J�����3�����>���]��ئNi�g]����_��j�����j����E��Lnd��>������Nw�U_O���鯁";7����" )�0�}��\ȿyn>�$��+�r{&�$�1��}F���A���f{(
"���2"��B���c��]�P�:s�9b7b�b}���캯�?�s�4I?k����Tsԟ�_��!-B]�JX;[�q0�8�,�K�(&�x
�.�Z۶�}�	����t������>���꾡D����/|s	=f4�lq���~�@����������*b��\� ��2u�W6I?>�I z�u���?�=�Y���=���
d���0%6��P��۴�5�G`��~��d�ۍ��_s�"�Ƿ͛�B��d�)J&|�3��k�<J���u�Z�%��a�;������K�yaY^�P<(�HA��}�NP#'L�({�{�f��)���Иɨ�o���[�f�����I�g��5�;N.�B�WB��{��>'��\���^x����(
`�&��޶� ��.�t*�3�)�.�&�������~��@W��!���x�u�����:P�a 5�D���a��2�ͳ�:PH�83E�ο���|��c�
Gq7�+�w�O�I���u@¥l:X� �wM#Ϸ���9�Fl0�D�W��=깯�MN��ZS���U|kۘ�ĀI��_P ��؊�ev{��@߉U��%&dLə�%��\�$�w:A r�s��6	�^��`�Ov��Od\L)�DJ�0�o��6���ݠH3UΙ$�t(��ut�Ƭ	Dz���Ϩ#�����/��1$��(�l�uD�E�d��e�� ���2~��u_k5��dKgO�;�(�{����0����\)����O\�C��y<�f�9���^�Vj�J2���
�r���=ԇ����,���������#��/���<�w�q���,]\�+�u[�Ɖ��sq�6�f��@l�&���ҵ�fΤ�Yj7��
͆93�k�b�>m�����<X���n��Q�ƨl��Oa��zPYK�K��6.[XӶ���d�R��n�A��{nA�=�x(W�,��j6����XN,S�=<�3�c��n�vd�+;q6���7i�CP�Ƭ+\�;<H��v�a��󶘁���׆{T�v����4��	HP��]�c���?����'6�h�4��|!�F��Y�͒I��B�n�aD��)P�S!�����Js%��.��?�'�@��TI ��Mr@�ǲFyG_�����Ҕ	"$�`뫯��F�t�$:�W��̙�T�f���fzC�b�E}�C��&DLR���*�s�x$gޅ:o>#s6��ud��޾s>�+���t}�5�� �g��O�:&�P�%@�o�Fz���Evn���x
�޽n��g���I=�ɯ�5�}L�����:��o��$n~SaDD�"L�u���e�����f�k3ABMÊ���cm�>|���6�(��{}E�����q�Q �Oo�����f��S�>�
���Y"����10�(
`�*����_���;��o�}d����k���NxO{_k��e��Bo�}��m/-����?;�X�lMy�Iuu��|<�p�w�s�=�R�������oQ?{ՓD}|�Ğ��+��Uﯦ�{q0�TD��(R=�U��s��	')��Z<6��^�)ϧ��PbcIӲ�	&$�g�\lت��b����7�����l����t�����U�]��2Lz�h��.�AG$��2�	���ξa�M޺^f��7�O�:E��l�~=���VDݵ��O�}��ۓA�b��Kv&�Ň��󎻍�N�O�5�Q�F���>}�.�����_��������n�	��k��V+FϤ�7�/�D�O�w�@�t8�(� TP[�������I���/a�o$C}�� ��t(z7j�1޻^�'���beH�*bT����}� �k�G��b�����/ߕK�#�^��l�A�FR��7�3|�,�ւ�3Z|���xC����KJ��s�X;pء_u��������?�t(���Q2�Hl�����8*���Nu���A;��$�t�\���?��~�	�O��($LH&<=�󫯨�F]uTs~�5��1nIW�m���"�$��qش���۽�{�:�B��?F��Yx�7��8��c��i���ӝ���R��f�k�����""LD��(Ow�Z�$��]Q ����3�";��2[���e��`��롏W��Ԋ%f�EbN�p�6>�����ﯶg��	���U_�7����1Y�zk�ۻ�ξRϒ�S
BTLV�g��A'ǫ*O���ݻ�D�c~��v�РA6��(�'u��"e@�*bT��կW�q�L�mQ�-z�+�A8��ǹ��*��z_U�#_8p�T�&����M^�٨xi~��T���9w�&�\�|��<8��kb6��~�ognZ���H�����$�ͪ479��b&B@����c�a�M�ܦW>�D{�V"�eQ ��mdP;�.�c�mV��N���zy�y�;����pMV�UK��r=�vJh:1�6^:���uq�].�������l��Q ���]eQ��p�m}$�#��6��/o��]}�Vc�qx��d��I2"&�B[����ę���4�.�U��]�oĂ@��`Q!ﯛ$΂�Gz#�;�(��f��DL�-�>��@�n� �M�g]��\�Y�[Y�!����W�%��D��l�b,��|ba�v��(����~=�̦Hok��l���ŏ���q@�V�"e(�Ĩ4���|Q��U������K^���ܦ	'㽮�O���u���i�����\�L뾹�:.�/M�����+�u�-k ���f�wd�0�t�,o���D<G�׽���/M��o9<О ��U�� B�^a2y�b���>�{�NM>�X_��ג���k���R��۫�� ��^_��Ƚ��D�g��3�H��E�c�o�Z��>�����O}z��ށ�N��۱N��$ъ���
���J��yL?Z6��м��6i��yY���3�ט�-���\��f�]�}D����5wv�Cf4���Q�;8OK������׌D�l]��od�W��w�C�h�,�/AЬC��zA��˃����o�4���,+ȁT��%Y 2g��dp�9���;�rwT@~ٷ�j����c�h��ӻD�������2����$�W�N��nG����������Y�H�Ǉ������*`
ͼ�x�>Yn{��]���SIOkP���x\�S�]�z{z󷤷����qv����M�{{�SL݃��>�Ű?�qA<��+�_�o�g���^|�$֧,X�b^c��;./�Q���!�)��x�^�H`�l]��z甭F4{[�V��o:;�bP�C"J+�w^���';��]F���o}�_/y�O&�uc�Z�
�<=흞�/pO��p���)��xz{��-�xKz0� o~��D����c�eͿd������C���0N�m�}p���{a�:]�wf+���,]<ƀ߯��C�swg7��V��x��E��M�CM�xġ�k#вjPc��#>�ssB�۱�	(���jI�:q�ެc�4?�rBx>Y-�3ŷh4�&e�Eb��X�����rʣw1FEģ�)6l�&�Oٜ��1�^��*�Ҫnf#[IX[V
*�rىQUUTj,�,�&�����qq�Ƣ� Hp��C�m��H�*0!FC�Ś,�Ml���b-��j �Z'\r
�lW�醳�%8�!W���)�*V JJT��I�c!HU�����TeM�`���C��-%�V@�lEc"$Ī4��XZ%T+X0�θ�� HÑ�-�e*E*YR̴X�)Eb2Ѥ�G�"Hr�0���h�pk�`99�!"�H� "��rRD�6�"8�(��" 	�q@I,P��Mpfk���c�U�#2��2�YKJ�QD�cE-�h��x�'2;i�"�[޲�)) �#ъU⊌z�ҡ�)e���LĢI  $`" ��L$�U�Py�1�D�rfBҨ*���"��c���>}�g�TjM6"�b`�BB盷;/X�{Wb�2꘦6��l�K)Vȭ�b��b�	��n�/oj�Z:����\4�������Ks���=�3�n������%�g5]�v_s'f��<�C�As�lH�`����t�)��ȴ��g����ݎ.W����˼]��:��=�]��a��Q��`%565������$�{M��k0/k7U](�⬶\(�����L��]�����ۃ9����{�kw$ڭ���&�v6�ܬ+%�]��,��9��Ӫum�t�V�F��G��Ò�P�嵮 ;l�)��G�K���I���N�Ғcn/[���'�a4Ϭb��=E��yюJ��t��ņ�Ѯ�<E�}����+�c�G�׳֘WUݵ��e����e�o^�vV�YJ�W-��/����M�a��h3��粬�볋�@۲S���|��D��\ڹ�RA#c��Vb]/Km�2�.�ue�V�5��[S��*�`�H��78��e�V�`��ᬛ���%ݨk��_fX�8.,g�
�ku{�qL�\"-�V��ѣ���D��e�����vY�����)���fu�b�4�i��5^�=h�q���ѷ�y�0h2��&K�sQ����+�VD�:;m\�k�"ěg92�͛�A��UtK4a�C����W$�mt��ɝ.��\��2X���ķ�Ge�B����p���˪ł�g`Un��w]4�w\r뜶�$��/[�y�י	��<:�sg��c[#S���M���]��{p����uA��t��y��,�\���n��<ɢ�Ӻ��n��p��h ݞ�5��dH*	�e6aR�R[������W';We)���f�WZ��6]{31�X�Lٕ��F�rM4��VXG5(�i��n����a���EF5M6n��z���{>3x�9��dݬ]n71�'\7�Z�e�k���&M�ؚ��?>[�|G���M��[�;�m�t��2O\oo8�۱��x�=&.&��F�j�[�r�Z�:MF���+y�M[��o)�um�m�A�5�Ɓ���gM�g�۵�ƛ�ծ������ۈ��<&���m����6r،����l5p��s@�v������G���%km/[C^�CJ�����
x|x��e�U��k]��)�p�T�Zڸ9�kv牥8I^ػkcգd�0�����2�V2��B�kn���ϟU�"dL���,޺�H;~ͦH$����OY�|�s/���n�P$w�)�7��q�#��"B�ŰlߝU�M���/vGϽ�A�A��T	����^ߡ����$*�$LȈ�2�	{Q=VI ���|E��[�U����"�qoĂG�׭�	�{��/�ym�L��P"_�yWfܣ躻�N��Sw5�	��r[�2Wv�������=Tͥ�A�D�L19�6H>�A:g����O�C�~��sO���РInx��ؽ�z�wcm�z��nu(��h��/e��]����qns5���{\��-3DDL��h*2&R�	LJ��+���=��Q#m����u��x�tf���6?v�}5ZoJffd ���=��D��u��5x�����{��z1�?,J��~܏��������\/,X��Kߏ��ێ[�؊��>��Vjn�˄&<�u�)췗\ �@��T	����4	3ף7�g�[�Ǎ��	JB(3���#�"��ײ��h[9�N�ĂA��B� �6�9WǾ��&dD)�	~�|��s��ǈ&|���V:�$�[K�>�~���Tϑ �=�Fe��R���3*K`k:��y]�ϖ���8��+�p��6��&}j��+��љI�+�o�����u�8��ʆ�F.3ar��MfAݝ4�T~2R�
cr�y#�A�d�L��t(����$ޭ�`��&3f����.��F|��lQ3��T(Ɉ�	LJ��fu�	�����0�vMl�vDD.��A#}]͂~5����.y�8�2����333! D��r�Ivc��#ݙy�-�(őxW8����>>X5�Ž�vgX��医��IM^������3�{� {/g��Ѫݣ�QX�c;�'�^ˁ@��>o�\i�#Q�"B�(C�[�Q�V�z�$���A��0�$���&;I�``�O*(��$u�1"!H�(O���?{�*������i����$����$���U]\�D���JwF�3@�����Ef� ה�o>wu)���V}�1t���?�|u��m������]�tʁ���k�?w5�2I=ݒ7-�|r7�]}�+=����{�X�:ԌJ�Cu'���Ov���%_go[��9���I'�����i��qs�#�4�>��D\B�̨/��՟	�r�q>����}�{=�������ZoFT�Ȑ��L�!��=�����Mt�I �ɢ.��=}�h��$�5�VW�w���3=�C�s�f��p��2A�p�'��O��ON�FNm��|�ـ{��o�]0����3�qR��]W��O(8L	�&�3����5t�X:������[������_P ��u�Q�"��44E=���Bz?J%|���n,(jPN/(qs �ǧ��E��\���P�i���=>��tL�oߤV�6;�$�v��A��uۡ��*�"����"�����^�2�)���%��P��&�DXb/S�5y絕��	'�2��L��$�Wc��)��	>��DL�R3
&[�:�� ��ȠI<|2�F~QӾ�	;ݒ(�!u�P&w|
����eAlg=��]��^��Y���%v]
$�=�@�C�|�k^ؽ�l�����5gp4eL̉
	����眒A̷���.qGVnv�%f:��䌝�������t=��gO�1EN�=��j�q�|��uֽ��KY����;��F�7����G���u����v�Sx>����0�.���6��3`��[-&���
�ڸ��lP-�@&�v���:m�����`��h6�Z,�L#^U�5�X���b��:53)���H�lM���\^���$�X��v%5����c��}v��#S\Z'Z���n���G6wB<uzo>ph�Ց�$�)�űXY��c�R�;�ƛǎu��%JGMԭm�ݧ���`��m/as!Ȁ��kCjv7"�q��P.�sn�x�68
�5����w�^ϖϥM4e�����Ǐ�D�۴$�A/��`��~��f:�7�g}�n�P�I�.(�Y2����%�!�sd���yhs��o1@��!+�qD�G��6H%D����{�4(��b�*!L������~�����~�UFE	���p�7�	/u�3wN��"d"��Q3A���2�!��~����}$�7�z�$���N�
��5���w��@�/|
����eA{;����ܪR�n2�hp���� {��lA'���]b��O�v$ X4��������]Ԍ����	b����;��67H��v�t����FT�̒���p�'3�����uF�k�<�U@΋������C�+ iHȐ�	0���V���C��n@��"�־�<F�2MLa��5qE�CD`���tp_�{��m�  ��O�"Uđf��A�a��_���Vwщ�z�Hy~w�B�$�G31���H������_
wo����J��ߵ^ƒ���L))&d�o�V��'��믅���1B=4=U��.�����_Q���b�R� D��7=Ր��"t��q��	���H��РI�!Nt��b���lsOJ""J)*&湢@0z�>���l���L��� ��o6H$��Я�.�������}]�^��߆�n%У��
S;O��	��=x-&#���f�/λ%j��׿�j��5v�Ow�׶�$�w6�_�#;ʾ ��]MO��捉s��$��˯���^����& ����QWC��w>�[���$���cb�P$neć&��}���%���HȐ�	0�j��c�:���};ʃ�"��}UG}�yprc����n=Umｩ�6�U@�Q�����Y�N�s�}|o����w�z�x��~�5U���A����|���Yd��)I3$K�s���oӾ��L��A&5z�=�|��={��}��o��'W�8B
ɘ�L�[�����٭Ȼ��{�{�@����#7ʈ;u|�����{�����c|��W,լN��k���zr�����=hɠ*��-n�����Kp��Lw��$ř_E|P$��l�3�j��	�bnb��>~���TL�x	ό%&Ks���'=�^�����z�>#�S���y?�þ�|GP����u�Y-̻c,0��̉ Ć��+u��� ��u2H^�͗'sn��N�3'O�g��TiK5��@������_i>w��{#�{�$z+9�	��f���A�߰nįZ�ӯ?���^o��v#�g��s!����ѷ��@�D�[S�cGxhWu����]�������6�������3�a��o�$F0fH��'��Ē}ݔ*�m�댚��>��4'2�i�Gă��@Wx����̛�ϒ}�	�:ܶ\����gk���U�-#`n��M�Y�[���k�R�C�~?[~��1��y��0�0�9��L	'������/vҩ���Ӏ�G��[�U{�""J%1WuH��¢g:r�j0�:�[�H=ݕ��;��r�ٺ�s��@��+�(ϊQ&Kmf�d�{7*���V{w|�)�)�h|Iݮ�`�H��vP����RbfD��bC`���5�}���?��S'�$N��g��A�Lw|���\�g���sTx���FD� I�;U�Dc�w��N� ��'��H$�s$P$F���t����ռsq'ӔjO���}M_Ͼ>��X�=�*��Q�����+nO%����+H�fޝtC�Q#|��=wvA�aA�
6Ox+ҸVhn�A�<��"v��d^C�s�8������[7]���.�\̹٭�2��:���'�Y��{5�����/B��l�vcmT��Ѻ�-q�q�
%��{At;�9}t=n΂皼�n�=�+rk��Jvۈ\��0c�Y[aV��c)U��)_]��}���.�����-۝\�C�툹z�z�F�x�ۜ�j���%f��{�X�e��'iE��s8[
�j�������$M������kd�O�r�A?Gd񯊾-��>C'�͂I7ݕ@D��2fL��f�R'[>����ikx��q ��M~���A�sϗ�7��j��wg�ν���D�0�)��]
$Gda�Ny�B]&�[����ݕ@�H���@�������2d���(~W�o��	&/�Ȣ~s������ttt��ߪ��I7�,)13"D�1#����ns:�.��ޙY�eT�&�*�$�ۛ4As�͝�G�9���ϿK�^VL:m�i��� Ρ�sI��v�k�avw���m
d�5����z��y�/D�!�e"I?9����$��c�G�n�H�ɳ@�����S'�lDo��B�U�t��r/
�@������q��⽕m������s�./g��������^�{٣�Q�\Tӟg���Mg
$�};:E��`��s�U�dܽɡyr�0fL���ʍ�$�gm?����Z��g�	'�Sf�����>u�(�
R	*b�vѾ���l��T�	<����I?zs����E�0�V0Y �צ�'��^AF���2d����H=�t*�״)�����Iu�͂~$�o����.��?DG�xeu�!�����Ę�-![p%[u���ݻh�3�2!DDL�X�f"fD	�bGw�_�ТF�f�`���ѧ�`�k3rV�� ��͒iKЌ�@����f�L��k�X����D��ھ���{}B���~=�ཱུ}>%P�c�ID��S���D�Xd_o��o^�k�Q4��*��9��F�z�</��>ōug%ɝ�Y~hzˇP�?'>{��k}8�������)�^"�aܤx	��VÌC{�+��.��'d��+�+җV%-��<����ܓ�{|��^n�,5�y}��Z�C4�|dC,k|��aY���1�ɿ�S�o^\n�ǹ[�Qxm��uڏ�U5�}.�>����C�^Tβ���̃a�])zK=N���6�_��
��m~���ŝ�s9X�F�v��2+��qF����MQ���.��{Ơ��h������_�x=�.!K��V�����%�o�Ď�O!~H˕	�L�c=�r�P6��|����-a6هW��c�=`z)�0�
z$w̹�ξ��\WKp����&-��gH���O{T���ݴ����d����ͫ<���rs�s�U��2�!�{7L�z�̞��F��]uP��O��:����/����[����	�hI�/��8U�|uB��!Y'��`�~L��ܗ}�i%7��.�1MW���^W�>w���y�w����8����m��<��N���r�g����:�'.�ܝꕯ��퉕�sogx�xK�}��3��G���N#��;�/!g�7����>򵊐����16-{�d����\/�R���5f�L���s���<9|�)x�I��9��Xv�{�w��ĕ�>6Ff�|YY���7��!�6�f���]>�%��IXR�R�C��f^�Q���(�p�M�a^i��y��E,��Q��`Pa"e HF#脂��L-�5�KJQ��ZVUd��EL������Ge�2l��gV7�.2�(ъ2��Y�� 1�XF �#O%+�)�D0��(�B�e�6rvp8":ت<ZQYs��&��c�Sj؂���m��e��*Q����AK*N��
6��  	�Qa�U#2�l���
�(ڏKB=E�9qFuQ��X��%�aio�H(F,x�RJ�+6�&�*)�D[VV	M��y8� ��:ȝkkp��lp�b=ֈ08�*ŉ�8,EDX�6Ҷ4J=E^���G� @7�p���4��U�XƱ�EH����! Q�$�lsINP�!(�0�)�(�9$8 Ze��DLe�EDR�U�@�ldH�@� a �pK��U�c�� Tg�*%T-j�Z�+b"�0j9IQE��MM1rգkLD�W�@AXC6������cl�����!r��a� ��	���� �=��l�	 �o��I=��DLʘ
[o������dWm7]L	�����A���D]�z��f��E�6OSv`�
R	*a���
J�퉳��	�9m�Oă��Eok���3g��x�-\���D����m�᭱q�����V'�Y��=��k���w*��~r
0&&|7�l�6	nk��~"��k�yaҎ����.z��A�t(��f4�(�d��{���Q��>��7ܺ�դ�w1�½���+��ٽ~3p���Q�-#�2$!L0�ګ� ��u�(�7CEJ��%��;�Wg$�k����HU�x`�(���-��s�&-ț��;=�DH9u�@Ev�8��S�Ui.�v�
r���"�wG)n�<�	v�8�{���D S����7@���{�R\ Ӝ�d,��L*Uk���H�uoA[��:a7���|*n����	��}��ak�v�9n�y�멢}]4H�]�͘~��V�M��+��$���$���H+�%��e�t�6���f�CB�bC���gϟ?O�#JE	*a�.��A�ʢA�|��=�Y�Y#��	z�k�{��Q�DD�0�m��lI0=�p�|�di �f� �՞���$�@ۿ=Q�^�r��Q��J��&"L�,�I?��Oę���tKk���x�����K���H��u$0�F� I������l{����g�X�� ���lI����,
�4�'����&�\V%"�����C�a�A��*�C�����@�Evw0�'��R/-��Z��hJ�/�ĆE�����ˇ��8Ocj�̼���mz<8Y�j"�b>�Y>Ȩ����wA����%)����.�l��k2\�r�]h{ԓ���FG��63�W���Ӽ�W�Dr�������1��G3uwQ�q��,kC]��Iݼ��5��-\s���}t��؎f��t<:v�H��<���s\���tl:L�\=�m�1b�!X��l�힓<���<\;03rEb��sq��r1a� �n3�<ͨ�ɺ��zѨո��[���k]�nW&����Ҭ5�W��mU�`hBL
��S/����DLĩAO��O?A��[���$Ow]P3w�קS��5�SJ� ���?��xl!)!%L8���w�f��Q�ѣ�ܱ��~���6��_P?~���<%fv�XH��)�����*`7x�ٷTI�쵂��n��4,%�����B������*��0TH��>��Z�bkLv�� �n��z��������A�I}�x;ộm�"5$8�F���=5�D��}B(T�(�������#�>�fu���1w*�=2����yx�: ��83�Y�ۧ9��A ���:�9����pP�&����% T�?GpP��Y ��Mc#�
�>C���37�6	��ݷTDI:<M�DLJ���>���Z^��}�����|����{w(˻t�b��
h �_w����>����>���;�c?Tl營�=L��aL�񃘝ǃ9b�j"ԦR]y���$�חT27�U_��Qb3j~R������@2�T�`��}D�]�� ���v쒳�釗�I�u@�H���D��ݰW�Q�DL�0=��<Y=�L�V۟
��MT�}DcWr�~&^o7��c�Kf*����S�_Q����	D���F}���PA �v�0tz�goDz�wWT	��!�ڢA �=�����
]�b?:�;��Oe�,����s��Һ���@9�-�׮�&*�6�u�-�Vݙ���'��K4lƎ95�D��b�T	�u�f��7_z/�+���}����%�L�
�g����W6H=S�zo�����@��!1ʉ�u�`W��Gs��{��v*>@�,x����()l��E�n����~��^����n�f��=[�#�Q�{����<-�<�\�9�n���_$=�m��>ݍ{������`z풙{#Շ�╄�¿v�I�
=[}L=M��@2�����:�ݪW�{�� G]E�$���l?��E�JS���X_�� �=�Th!L������]
���Wa�o�g�6hH�<�$�s������z�֜�D���~,���kˋ2m(�m]E�{k���.�]�¹�n��m��}�q��l�i������t ��`�����u_<���z��6I/�sd���ȅ˂0�D�xx�j��#���3�r������[$��jc���Al��H̬��o3��$�Q�?E07�Z�$���:���J�ue�F��vGa�@$o������Q�W�D��:��1*PS��GN��<�k���~��d�f9�H&=��}�����JZrz��?������3,Q.��u�)G
^�xq��ޘ}n��Ul�����96�����Γ9b�?y
�ޭ�(�}'����l�7���#D}(!L{����D{�(-�v��+�+���MܼlH>�u�|D{g��D�pn�{̕e����uˍ��Q���j�E��^�<�ث<gDp�baP��u���_DL�0;�ݸ��I��U�$G�x��M�/n�Q�L�K��a�G�=49�(��3"Ɇ�>�΀�������o�r��$�=y�	�=ʉ�܏
ʳQ>�Z��C�V��`)��a���I �+�@$���.��fJ>�B2���{3�@�	��U�}�RT	(dO��z��w����vp�&�f�;�dP'���>��uo;�&=�Fd'��f�
XZ�M���he]��s�Ց=�J�گ� �{6h��m��u鮔Q�r�SG�<��h�y?��۶~4���k)�x���{��c�����bj/c����ḫ�i������5��v���J�?G�0p`���K-C@�jQ���9��ys���[��'����wk:P5�;FE�[��u��̛�^�Z����Ξ��7lm=�s���msǵ͹F$�U�Ҧ��,m9���/l�{eT=�L��sԏ�-��o7d�����v/S㋂:[j�ų`AY��6��l!.�ש���ұ��ICa5�w<ٺ�]
������uS����n��Ζ�+A���@��T`��v*�\���U�*��Q
O|/w�AA���p.���A&}���'�wo��lȾ�:яex.�3U@�D��w�D<�$LLL��{w=�3�0�izz���H'�9s��AGu��`����f.W��Q�cBv��f$�2}9	��纃�����V��y�g�[�TI'�~�`��V�#
D"fg����@$��~����$����WF	��/�>4L���J	�|��_Ē#�{��{a1��y�~S�Ɓ��Xdou�����C���1�f�պ�K	Z	ը�Hf�*�V�t��s5��8)-�Ni[h~}q�ߠ��s:���t�ēy�[����4o=f�=�S��|���H�׍�Hϱ����$�
c�����>[��ꎔ=!��w+�o�����^�}�����o=�6���4,8V� v��C>W<1qY,�s^�;��Z{T��ǲ葞��y>����Uo_tn��ה�"��{���к㛎�����x��Q�	3
T�����${v����w��6�v	�>lOǻ���9�b�"!��1[ҟ�ۨ�*����{޻��ve�A"_GzD�WE����s�
s[`�b�h�Ȉ&a�>=5�D��(O{,f��`�ώQ?z<��g3.E H���_�~����"&J���
)˴�ͬwSQ�Vۙy#�Ig�5�� �t�AR���I`<H���$Gp��kdy�T~$!m�Q��W}�?[��6�������$'B"$��-���	%z��<9��랺�'��uD�!u�
�i-���k���?kn�A
2L�f�ڿ��`����M����{��"b�� |��/-:%O�,ݧЫ�t���y5�^���<i^�� 纃:�{�m��{���0oH^*�Mw=A\��{o�O�.�}�����j�f+<���M���qx�_׀q�$�H�ב_O��|�^�E��$����l�#DLɈ����_P�	sS+Ǎ���i���ѿ%��uW� �^���F{_6kw;rtuZ��"L��"2�{�w=Z*Gr���r�ӳ�Kl���K�:�<���i>����f5����~�I��(I$��3\�+xE�x�A�̑@�^̊�7��{7�t�9��*�A���F��������I��]��$����'�!{�Z��"V�����huDI��"}�`�u$M�n���3X��g:��H���	����x��� �Fa���@�_D��IF�����#����9�RB%�R���^1y�S�eߦ���n����z�B�o��J��ȍ�A,SX*��Q�
Jv3f�������Tr��$�b�$f���$L	�Cs���${v����/�_ܦ�(	�u�OĞ�}n�����������pL��&�$Ke�$�3rW&|Z�X�������gϐ�۲[����y��$���͠�"�HouP�QT��]Z��A#������ ��) L0�魪 ����EI�	��[$����1�"�a���'�	`�&J*�!����	$�uТ	��v�r�şN���E�H �y��w���1 ����1&fP�a|�9+ѹ�$�]��v]P ½�4=������U�'�]\�$���������e	^�͹Y�iݣ�w�2G���B�!+�%�I��g�|������
"��'��TT_����Qg�0`�$Uѫ� �CL@P+# BA0�# ��E21A,H39�p���!���0D0D00@3Ph�  �U�W�X�`��$ ��`����A��*���` `*���g�#1`���Qh�B�$
0`�E�X8��F.(XÊ4Q`�E�PX1Q`��TX0`���E�X0`��TX1A`�E�X�X�T �08UF� ��5���mj������ �Ȉ��1(�&�V�p�����W�������k�g����~�����!����c�7��G������׷��o�^'�"(���W���W�����@~��ADV�����i�� ��"}Q����O�})�~~"���?g����׻��f�?+���%����jl>����W����>II��yT_���U?�UD�PBbD "$XVA  �@ "�`� VEYUsT�*�X "��`����H���3��I��V>ϯ���@E�-@@$F~�~��6?���{�d,_��}�2����ϰ����}�"(��>r��i��?q�/d5����d�9O���g����������p��+���? �$؟^_����~�N����
���DQ�����9��?!�PWG!���2��0wX�O��L'� �p9�K A�@���?�x>h�6{=��L hDQ����aO�O������"���tO{�P=������������w�=���<>)�}��}����{����?pv���DVo��#�|�"����>�����}eC��W`RC�(z�{�����]�"��� cف�!�o��""��^�$�t}D>P����Z��}}��Ưg������~E��
��@���>^!�o�PW�Ǳ�?����|t������|�����)�����e��0(���17�   A@ �)@  

 @ 2 
 �
(�J� P@   �U�� h*� �
 � (+�@
 (
 T )AJ
��E P�I@  ��� QZ� ��                                     
    �  ()�F�U��* �24
� �A��&�!f2�U���� 4��R� �(P��: �r�S��H �(�PEV�:HAM.a��qp 9�*�A��fU!W-R�Ũ��J�9�\�hR� Р�J��(        t 4�R*��IU2iR^��q4(R�r�%R�WN ¤QF#:�$*�T��P���]e\�(U�� sTIf�$J��U�*� �q"� �G#A!�*� @��Jf"1j����`  Z�)��B��$VZ
=� $�   �       �X�PZ�EVF�K6�T�� Ҳh��G�knf�Jq�C�OU�.��[��
�QO   �v�FQr��a٤l� ]�R��s���7WIa.f�ڲk��\�7 �um.f�5U�7S�1���t�����<D �(�  �         z�y9�;SSnvsiW-Jl�ݵJa� �:im�7��������q��wR�fp .��B��Y;�� � �^  9]�j�ծf��\ y޲�y�.�.7+�֗;�]����m�Ln wm�m9�q��m��.M���v-j�(NI@�P<  �         {��[g6�-5���+��.n�[k5nn��1� �kmOy���V���ىs��\m�J�7 �]f\�ښf��r�X PP���H�^�:�i��Gkep 3T�Yt��K����������J�7 ��!�A���"�� 5<���M4  E?!�)U��ɉ�LL�ت��UOԀ  5Oz�h*�   	4�4OT�I�b0'������?ܢ?������ן�b�a��,����!!I���9!!I�@�HH�HH@��$$ I?�	!H��< ���?]�?�~���1���f�-\��ݙn#z�i��U�%AM�Ӳ�U7AՌϮ�w��x����'�Ū�!R�h/k��e��N�[F.��5��zhG3�ND�=v�����a���-/�&-���x��ۗ`kr�&��U���`mf��p��ʁ:;[`�����H�Ů]�5����ٲFv�)�W�g�D�he[��/%Ɍc��Æ���peZ��{0mIhc������A;��i��;v�݃1ԗ��2�X����H5sj=H(^����q��;siԤᱬ���/f���N�� j�fc�6�-I�6	{��.�t�Ij��u����<�NyE� +4�v���"K��\�{d���~�Kʼ��kX�d�DzwI0t�9�0ld�MK:]�_]�XVLkl���ùY�93 ����7m��P5�S�
{f�23����*R����6	ǳp���[��l��=v�+�fm�Ԏ�p,��Lm:6�ɑ��l��
٥触��/[��,A��2}cwV��&���n�Yg2�c�X)MŬ�h!#5��T,b���(-��I�;y����j7��%�������U��f`Ŵ���*�eeɑ`B�6�A݄���(=v�ʎh�{�t*7z��ײ��S�([9�^��˂��CI�]^��������ݝ�a+3/̬���{,խ1��z���
$�nЈȧ"�P(�k-�i�W"!�űb�,��k]�!�ÚR�&��i-�:�ٻw��lʛ����U�8�0Hr���
܂�.��԰o*�Lٱ�قK��#FV�"u+@��զR������ѻ�U2�LCz�ndUbRF7Y��
Wd�ʯl��1)N�nݪ�� )6��6�\;�'��2�{5�,��SV$I����DR�
34�wp����#ۨ�X�T�t6�����`��ЊGu�`&��Iǰ��K�.�#yQIlY,�ѕ��AЃ2��t�S^��16�����,QكqD �Lւ��x�7&�6�+rfк�37]����כ�2�7
�b�س.a�ԙ&4�Zu�`��we�p��z�^Ś>�a�t���K#+j�٦�֣O4S���[�a�,��LX%��Gk�4!����.��k�-zq�1#׷,,u%�a���^42�L�N,a"ī*C �lI�
�N16��*�)��b&�Q0a�T�l�`�fR����M!�ۃ���.�}*�L���6C�t]j�CP�ܻ�L7�Rֽ�u'Smd�Z52T�u���e�H��\X�Wi]�M��̓l�(m�X�e��Y�)���Qː�T��WUsA��x^J�n��J�4�4S�.���VY8�V��T�	-=��a�a36��4p��.��t�F�4����%��dr[ue�k[.JT�ѣ���$���#	S�u�ŶF^n���e��\ͧ����SE���9�V��m0��Y��3Z[���a7�e��ٶF���ޱ�2�`���e�2TY5�싶�^e�cn�d@�T:�"ƚ��y����3st|ȟ�&V���	G[��4~�/@ʹSoq�#V�m����]��b�w�7]�c�{A�f�p��v,����Ź7Zk {�bZl���4`y@dF�[�Mb�ho)ę���V��f�Ԡ��B*�L�MKS�%S>4JN�	"+Hs�Jln�Ҷ]�V˽�r��.�$��]�ܺF�@^a����[��3B)a:kȰ���S1�T��^w�ُ,XTܡ�+a�0�[��$� �J_֍�ՋH��WtcʇЭ���ܹP9(���q�줶�T%M��kt�w��� uղb�2�/���L:)ݝ�E�Y{�hS n�at�	���V0�J���*d�m�ԑ`PE���"@�����Ym�̺957j���2ؘ�S�C}�s"��P�[�K�r,���˽&�#�h��+M�,<�طke�� �D�	*������d�ښ��eY J�%aIU�ԕ*o0��y"�Z�yW��C����Lⶵ�Զ�m̎��Y1���(�F�S���E�`v���1�&�T��O�AO�(fc��	L�&�R�N�%�fb�Fz�	r�Q�� p8(��a���nR�w�!6���W�4���]�n�]`@�h$�{��^:�r�@.���ĭY�Mˑݣ�fڂ�tG)ʟ[;v�e�%3�I��4��N@��U��;�x�Rw(Vlx���g�tV��'��ʻo5Mfl;Z��k��6�ڀ�NP"EdC�!�D;�1r�0�]ՠQj��쵔����.k":�
ʺ��B�-���M*ȉ��#f�-e34LȮ�f�[.�+&�P��`�^�j
�p��zm��e^%�Bb{�HU�(�+vV]z0ME�0�e����K���PdFYw%�h�V���l9[iTq�.J$�l�Jח";�O/d��u��v]�w��l�7@�	T�b�N6Υ�Vض��W��fel�2���|5Mة��МY���5�J�r���)�zF}�F��Q�ۤ����ɖ�6�_�)Z, ��j�m]V]$�-"�IG؎m�uhs.'�����U����Z��se�-;�1'7/^�Z����K�ƫ���K���S��(�k.��!0jO�Sbź�Ć<)�mVS۠��un��S��!B��~�\��ϝI6��i/���*��@��lf婺�G��#��]��n�t�W��h�V��m*+��zn,ڕ�N˂��U��Y1��ؙҲ�b�j�wfڥ��a��(�\�$��T�����*Vh��Ƌt�-Z��M� �r� �k\/U̉�Ӛ��yI��i�wi�=:L,6L�6+���H��+��@��@˖b۲ӵ)c�wm�i+�k1��)��i��tm�CoK͈>md����l�*˗M�h���V�!Y`*6��q�*��ܫ+Dж�{��(��͸Vۢ��=YqƔg[�wv	�Z�LX��yW�X� )�;yn��cn�8tM �w��s\�h��9r�RڌGJ���c
��-��6��5Se"��Q��2�B��"S"�"$�����aТE���0�5�\�d���,k�+.b��U�uV�r�=����G'[�:z�x�۽����Y�vQ���Sĳe���@1�t�B�J��U���;#Oa������(�7JE�0͇�N���U���n)QK�qz���ʖl�H܎��F�Z�N�XGwA����u���d�W6����vB�,S;V2!�j\���c+Y_gE[�����$
@7�R�իpT�@�LB�����-���FD�F�&ֈ&�q;�ZN�~�iE.M��l�	�o[��x��l`������-#���tj��ޛ'�H<�e�/n��[�{.��ɫ�X���{��n�5wZ1T��R�+������3A�p������FTI�Һ`M�pɹCa�8w&�G/,�����bڻW*
J�ݙ��q����r��:�G��6�r�jԲ��Hj�Ll�i���GQQ�S0�Ԑ��W"yj�L���!Yx;�!2�TJ�<��T����e'2E�\n�;�-wl�t �ƨ����XɷJ'y���KF�N��7f���YH%CK��c&hݬP.��"��d2�V��0��eR��F�ݑXܦ\�,�O!z`��]���',��Xe��H��l"�I��B���XS�]�,�n������V�1U��ʱ*nE�q�*���o�H�-ĝl�@[�ʄ�F�YLݻ�t%[�:x�cBó{C*m^" ��Q(��,2�������$̻n�oIJ�R��$)�m��M�CH�޼̦���Sv騬 &�Q�`M����#[$���6���������7�i���ݻ5���6�+ �.�p�F 4\�9��aa������@�3k H�;z&i�2�%:V
��UŴ��ɜ�sV�\(l��t�s	��b0M���;lYs�w0wk~deejdY
{�O%H(mB^��W6��7�u�b֯�V'ڷ&�K+&M
Io>�D��@��LK57�4S�Đ���ni[Z�F��V�+� �Q5Ol���jsb�:�QՕs]���RX����B&�u`�6�:��(�\lRxL�I'.̺�xF�V�j�F��6�K^
�{�Z8���[4~�2��^+�S6�0f�Oh�Fթ�jeٴɛ.є��!l(ƛ^�)�nf���5lfJ��E�ȸ�s�n^���2������wQ+����i+^���f����,��U��e�o-K�J݂����R��˺F�PԮd�2�71W�)�*��
��v�6���7���z,�ll�0�"ai�V^��E;c�`�VJ�5��Y�2��m�a�H�F�%p�,�A�(ԛqm�/�Pf�94-O����������Aj�5q� �H#1�q�r��TN\R�B�oi��d�1Tf�a�`-(y�2D�Ta���7FJ�f� V�X�<�N\"T�f�U��@;H�j�إ�۽�I�2�ۯ�8��D��d|[���TL����7Z����� �*��/-ZVNMim�eZ֍ՙ�L��	������R�����[-�-�Y�􊼬
�cV�̓ub��e3m-����)c�5mj�����o�@L�0�ܼ�j=�S�������!��B����ML˘L�s���{4�p��$�p��jteY�*Zi�
T��E�g$,�ǒ%��mظx�(�6"x���*����	;�u-�T�ͣ��W�h�d���v�]hd�2RBK ����݊T�ܸ���r;3uRy D��j���؀S*��x�5�/�T��J�^���k@p�w�I�c6k�����з����-|��V.!ol\&f���[YVi�Ǣ����W��`��+�S��.fĴ���L܅9S� ��ŭ��n�zj[�av
�&U��Ac�h�)�מ(����^,a�ͳT����P�,rLpb(���`]KwO�7j�@f�Wb���hӡ���R(A8�BRolm��V];ͽ�a�[���9�ckm�7��*�L���b��]�m��ړ!X��+b����+H�"��#��׺��yr�jK.��B8v�=/])G�^gD��(4R���B�̠�a.���];aڷ��+����q���
v� ɻC��P�.)�8�C���W�ښ�b�(�:*BVd�n�t�E�м�c���wL��aD2�+�Q.^	�0NVp�r"���Ɔ
������d`�ƤƊ9P�i�{�l͠ӽo*ޛ�ˠ����Ѭi��RnS��+em��2�V^���B�L:�k����;�1d׆ba�	��v\0G�7fZF���&���/�&'G5��"� �@��+v`"���mU��ݦ�j1�K�B�dڵ��/-e�q�%�yv��St�r��t�^'�^ꆜ߰���"3�Ԁ�0��կE�O�ܭÇڛeմ�F������,*�:̷d%�M1�ّ(�v0"���A�V��dJf�3b� ��b���z%1Z*�A˗P�2����G0��������Z��܂�6b��D,=z �f���dܒ�c��[��,�N���N��Ձ�jK�Н&���Ͷb�v5��)/$	��1�Ԏ��2Z��:P��3~ e�qS&�Q��T�Poq�[N�ion#{o�R���!X7j8�V����ac��EeP�B�:m�3�����Tl���H�i��乆�kt�U��x�/UW����n;�H$�s嫓^�E�+i�ƒ�U{���J���k�xڵ!��8U��,��U��2VU��
�vu^�6y�\�Vb;ch9u�<oq�8j����P�ۚ� W���ݧ��XP̎Kț��
�gp7Cnma	 ���f��\0��6 ����
քn��C�6A�n7a]�1�n�;��:���f*;oB+v����/.-[��w��ҬۏИu1D-��&���W�$��<�D����.7M��
������8�"��w���ř�X�t��f�iĂM��r��f�y��e���[$¤�p�Y�fU��)�`f�e�)���ʽ7�*/&�[&솬�����h^�����IA.��b�F䊝L���TU�.��(����^'���Kb��6��X��]:I��ooMqE��=���-�̹6��z��Uj-����K1�F�T���c|�+�::��8R��`����u�Z�2E�F��`Y���a@v*�:���۴�CٕW�wL��F�\�\ʼ�.|Y���&��4!3!0Fc�(�Ĉ��dDۘ�p�I��!⊓)&�T�B�Hvx^
'-�ԫ�م�pe���X����(�j�D��0.�lP[��Cv��(�Z�6AE�p��YG�=�,Y���u��ԙ�$���t�����m��b��7Eطq�tf�D�nNG��<���B�
g�3b��0�Tو���bZ�H��$䧂����jwcL�Ӂ\R DL�Sȩ��!�HJ�[�i^�V��[t�N�$�������d�+T�b�[��v��ڗ�kCת�:�� P=�m&�Ml�;bT:c���˖��S�,2�,�q�$�#wԫ]Y�)˛J����/5l��
�E�p�r�^��t-�k���Gk��HU�LIlK���R���}*���Q�Ze��Ń�WeR�oQ@�*��n�Ɓ������[e�f31��\����� ����� ��)$� ��*�d�"��R"��)@YP +Hd��	*��"�!$���P�$�T�I!+	
��a		RI
�XHX�$P(@RI�BB�%aI"� (HAd�+T	��+ ��"�,�"��� E ���E() %d���RH�Hd	+ %I	"�(H�Aa$�XB	�	�"�	XV EHE����d�,$��@ "�,E  �H��I��+%@�E���!*�	+RJ�T� �� ) ``�+!
�$�� @$$?�$�	'����������{y����<�
*�-��8Wf䇳�
��C�<nܭ�,KoPu��*�F���{�;)�U"B��x�]�eK�wک[뱹�X�-x�'@n����8��/>�E��5���Ψ�a�������nO���soQ��ɫ�t�"��b=W@�\�{�R��u�v|��f�1+(�C	*"!H{3��eF��>��q�b�Ű�;�����R#0��%���m�6FD�D�C
��+)ºR)�`����*�����{��,]��[�=W�����]����(�FJ'uZU碡jwN	7S�Z�<Ǩć:�T��6�J��B���J����6�IO����w��%�yO��$e�=.lB\xm�jZx��K�tL��-�8��wZ[�����r��`����v0��&�tg7��m\�̼�mr�̳9hoqc�Re��n�fp9�B�jg��{:�K��Y�r�{�8H�X��͹hi�L�6�ob�7:�T]�e�T�S�\Ƀ���^�7\�If�0�q�s��7����k
t)#Ќ���{Z��,�3��ѭ�`�XgKEDȴ"��nU�Ѽ�E�Uf�fc��K&GD�>��������R�d������m�ZGS�/r���h^�c����r_qF���rA�,A�EueYjщ�1Y|9�Ԏ���ѹ2_Q���:Q���$��v�35fϑ�g�(���YՕ:tN��j�5��;�}�(���t�����b�qY��S��+vvY�/.�H�ĲѦۼVؼN�<�����>0�yQF�o`D˚�ux��h�Wa�{zv�D��k�r�EH�my��?-��uܲI�X��g
��'m�5��[�M���<��;Ͼ6����ҷX���֧=��T/u�DwF�M˓4d+K݅t�
<���A��:��JIW���;�J\A�go�Up���=�:�+v�R]�N�g���fn%�f�e`um���q병� Ա`ڗ4i�d�a��]AG^v՗���+T�S��]�1�[����}�@voiz��V����.�A�s~� ��FA��k��%1��Tn!��.�lͥ��_Q�8�{f�#�hlF|_m-o1PY�9�.��c���Q�W�����9)M��-�\GY�Cl'L�&�b���Ɗq{掙��ݍ4�ݼ�������w�V����۬.�B�:��Vr�|��W�Ob�Y�,��5;4���#Ce��qX�B'�y��4�b�BM5�;E�Vn\|W[̱��u�dV� =���H�a�1���QY�����umt]�ݐn��&ѽ�K[�ݗ���2�>��f@�VǫR��;$��m^��@�\Rx^�j�ge=c��E'�*뱔�"�k�P��Zk��!�[L��0e�SX���_X��%��>�U�6�nsV������ԏTIm��z+v�6��V3��\ҳgukvz+�T�m��U���Qm��+mn��u���}u2$�s�	y�0�+���2И�T��c<d�:�������u|�@��k4����tS��)�]u�*�7�(�]�X��w*�۬�Xk���cQ�Ǻ�:k��fPU���U�x���Șktڇ��e��WP��;-_CS���66�2�� W������Bǻ(軇n�T�T�P'Ki�7����Փ@�׼-������3���3UͯT�ۙTSV�HZ������3��s#5�����l�x��ZX&}��{�����ɤ4(ݥ���a`����*6�L�KGDӳ"��;�����ٛ��V�C�����p^��*��"�v+C��.�����_fwj� (U��_:$�Ӽ�^��\7(Be��V;6��g]��)}vɎ�a��@f���nò��n��+l��n��WRc�Y�MNG���X�I�Adt��x��/�o7��c����pW��Q�t&�|k0�'��"� �zP�Ua]�gX[-�x����K�轫4��i��K�j��c�nP��һ��!	�V����� Yj3$h�)�����F�i�v��Z��"A$=n�u����ͽ7c�=y��F�<4ڗoA�O�N��_����7$Wبw3j�X�
��=a�-��U׶_p��x$�r�H]�F�n�B�͚v�$V9�@s�>�]k�*����6�,�5�����Ƣ1�]zy�ј�8�K�E�	E-]St��{��\�˺�U��ut���e���d��Ln�F.׎��1�w�U�J��;B�*ln�Q�ͪ�-�>k���z.��C0[�٨rK��*�F�����h-Ś �r�s���J�Z�gκهB�nD�x�@5�t{Zt��>qH�㮴 ���[;n�L�B�\T��c����u���74,�Vfn����(�3e�\�b�k9�@�c�����fvB� "���G�h����Oe�4�5`ݭ�sI�9cw�{<m	ע�Č�m�ĄЬ"���oIYߕ9�X��w��j^f=@ٳ  У��2Q��ï3�p
��.�L��9���v�����n���G�7/��r��+���o��c^�m���ޟ$u�G�R�'D�іR	�k�����g.Ym�7�Xb!u��t��ř{��T����>鲒:v+��wo�U�rV��U0{_u������~���j��+�d!)�����U֣�{I�4Q�)�!v�+k�b��L��Ϧv��y�pw4���|�q�����[@1:�cQ��M���4����7j�>�UuJvC��/�4.�j�����*����=>r�W<�l��P�9�m]���O"�кmS@������f�y�SV�f
����s���w��F�eM��7_�Ih5deE��&�E�ѨN9)\�&�'K��I�����n�t
���e]:��☽*�����o�fj���V� �ooX��q�d.��ׯ�$�U���j�nJ2��;\����2�Cr��p��ݷi=�� pfdsF��.q�q���Ery-N�2���v6Ԕ�h��+��5��Q ��U���wdp���J�LxI9��x�-�y���r��X<�kk.n��e�ܜDh��^��K��:��$���Y/`�5mF��&��.�,��{�.iǕ�igA�n	@��bB��6b���.⃮��-�F�|��H6�}�y��&��<��6��}����!ݓ�>��f���`i�/u���D�Cn�v�z�hqD���w@�����Ou�|���s)��{��C;\�6]ruv����l�q�!����Hj�1���`>7���9D���{4J�᱅�V����q�mGh�S*�,$�Z����ff�˵ս�V���חeeJy�̳�5j
�W=Db�
]�㕭q�8�&��+nN�t�h%5ޕmث݀����AT��9�:�ؼb36p�9�d缣�<
	殼��%�s��CT��X� ��짳�H�Ֆ�Ay:�w!����u��:�	�y�6��2��s�Qsx2[{���������^�c���VF�e uZ�1��)��[7����I����tn�_[�Y+��K'�p����)Mޣ5$��ٕ��bg�[��z9e�nG�q�B�x�a�	�[���Ml#G���y�mdy�i�-CB+h\=�d'��IɅP�k*�l��7U.S��zՍ�wh�!�9�u��0�{�̓7i�ZFD�5�-L��u��LnNv��vOV�ZAP���p318����{�&퉐F�"��`��jI���]�S.��K3A���Đ�y]�������Օ���N�����7�dD�1������&���r��gi�<���F�۴re�ps��a粩��0w�6]GՔT|��@G��3{gP�m'���Izid�ײ�/�Ӎj{s0T�y��B����%�Z8LѸ�e�w��$��={m(;�b��䎥<d�WV��f�M��g����.ڰ�&R���n˳��U���J�}��]G������ْ�3�c+]�qpĉ�ݕ�U��ϙ0::3F��DM-b.DM6��ƌW4_���i�q�(��U�8곘ϫ#c�˩-�����T����v��ݚ��k;Y�;���{�S���N@��ڄ���b�u\d�Q�c�T�.�,�[j�o��f���8@v�P��e�V�u<�!�ͫw����\{Voo1v�,Q7���5�l�!��e��r��e�̳F��s;�6��kY{`��6@��V�V�Wc�v����-�����/�����΃�[u�M^�n��N��s;D�w��켜�tfd�5��ڋD�q�6��rKK�
�b�A�v��(N�]+��ce����0Qӕ"\{-%;�\Hm8jvFL[��}j�w�̩�:�7,n�V�mMde�|KE�;�]����:�k5���L7��]��w{c�Ci�.��f��ܗ2�V�l�����ͧ���4e�<�h3�Yۻ�gG�xo
���v-R��쭚��7o�f=&v������T��ut�^T�C5$���9F��ټ�.�#�1Mq]e�����|���s��A�,���Z̼��;����^l<Ķ�v����e;a�)F]F���Y���/q�ջ����:f�+�g�n���w����,Zr]�0�gt�ل^�Nu^,�++gE�Z������N����m+f�|D2ü�ش�!a����U�Z;7)NZ�f���6�\{�\��,���ťL)f�e�'E��=*n�aK��ϖ���I�òQgu�a��-�_'r�X�s��ޠ��u=��t�7铳(;O�<��z)<��Fs��nۥ�����5�;s��[ͣ+x���wφ�}X�Lг7m����iΫ��sg�*J����s1074��4�Z5Aow�<�]��+;�mǷ34�]�]^,
��fM�P&��7Z7Eh9Q�E�n�4�r��J�K�XY�R���m�mN��w-9�R�����&�kL�!ɇX�D=0�!c6�);�Ã$7�w�x7nu
g�a�w��Ŧ��-���Osr(��*��yn�ڊΥs��\�v�]#�A[tm�sܦ�����>��N��w! ��X1��k���;C-n��lP���!
�xͺ<�.����m�RV��+;��׸J�'0��3��A��x�L6b7_�����QS�15d�]ƘܨZ�ĹH0ڳ3��)�[��m��U��^��O+.�.���J��u�5.��
��9.;�ESv�4��z.�+m�
�~XUK�YP;�y�0�ʷ�>�`\�mIr�fաD.�V�5; �.�J�ʼXS�4�"�C.�V+��}�8��R��W8�=[5�_2��G�Q����*��a���DpΎ����²���_e���X괆[ғB�6rي':�K�.ٙ�v�<�\�;o.�[�V��r�r/e�Cz�*8�P®�mp��{�e�f��2M�k��k�n&J  �$�R��ݼ9�[�z�r9Z3��0H4\
�(���6�j�u��f�6�w{����={}�	�V%H���J����Ϛ��㫺�WJ�U��*�m�R�6r�L���7�;av��:sy��|2u�[]�8;wR��f�q�vf�:H��v.��ZY�a-���u��s�v�3+�z�����x�&��]��:n�w�΅�4� r�����
b�'3��1�29�.:+����L�Ҷ��w�A%�f0�L�jM<�;�{Y��fR޻���w�{۫	�f4Y�4ՒVvQ�.��=�h�.�SY{��^�nik�P��-���IF;y�X{�;��V�%D����.дsim+WV�v�ZGcZF�Lf�K�Ư��UI�o;#�sX�͸91ctWn�
�;��zs�T6�˼Z����ɹZ� M��oFYB񉡾΄��`�c��۱�i��K0^���a��hZ�63n:0^�z1�BN֜�������T�K��ݡ��|�X�V_&z����avm���Z�bn�:�Vm�eu�CZ��C:��yM����/0�A�-×';�zz���|�7��g.��`[chE��]�tK:��ӷ�֬�z6�����ͽη�6S�5>�<2a����^����a�ar/ms����F�קr�&F5�.��N���"���VzQ]�{�Rt�3���Yq�qk�\�d���H�Bu�8����-�z���Ħ%wV�E�Jn��-�Ɍ���Mv+�ś"9}�j�C�mw�qV񼋑$Z���=[w"/��N��W=$*�1�\[��
a�[@�dܬ5F�6�W[l�z�f�'ݵ��$��֚+M�tGrwF�}��xm����4Y��Y����_v�h���n��hĥ���V�q�`��,���{P��t�޳l�*\`��r�hԲ.U�nTݑ�2��	��iT�.�[U���&�u��!yǢӯ�r��z�\Wwˍ��:t1c7raa��Ȋ��*X�l�i^x>S������r�P�(�颗2��%�O�]i7���%��'NV�L�h�Q�탱|��j�Wk�qn���{8LM�Q���+i���1X�"��0�p����[�@Gq^�n0,�t4c���4!	�(�/�X2��ݳ+i.��M�8�p�9 !����ӹ��S��z����5����ܡͶo��.�,�;`���"s�-ޚ�3�-�1,���Ε2Wh��O����y6o5�7.���U� nm0p���sB�d�52!n�i]�Z��}K1 ��7�N1��P�n�N�����[�ĺ����,�nk�Ϟ���敖m�r�slm\d9���>8�)t�\k@1,��Ni�Z(�oP�X���G1Xͳ#j��+Ybl��.�>��^���l}چ��h3H���4�UL�Jubk|�U���+QWK�0�f��n^����{z򕴷�S�+1(�F2���8�2�r�;�lf���|��z�3|�{����I	OI$�r�?x[k��o#!]Oa�0K/99�"����b�<���5ěa��C�6x�*�y]�[�|����n��i�l�1�s�Lôq:kiz�V��x`�!�ŧ��.x4czOe���a���.S����u]�q����ZԆ�Y��ɵ'L�9Q�[��Ήg]�ۥ��n7l�^ �lez˒4�>�e�Sr�q�ch͋���n���JV8��۵�Ԏ�&0��Q����R�ι���ݵў[q�v�k���s���O`��!��=�nm9N�nun��ny��^�n����b�i���e�8M��8�m�G�w
��\�Ԑ�V����U�o�l<���L��[�u��@I�L�w>��Kt��\�k�N�1\�)m[�:����ދ{9��%����N�^�H�@&8�s�)��LnƗ��<N.V�Þ��u�듖�'ψ�z������\N���5d�v���1���a�od���Wm��f]�����Y�y:�t��O&1��P�۱���\�[���<���ās�]����k��ۣ���]�k3xٻu�s�յ�50��ݸ�vG���׊b�Y�ٷBea���U����iĐnG�c\���Lh��1�;���L��L(��̼��A�g�v{z7s��6��y�Og��������z�����+r��pq=Q�RlpG>��݇�<Gl���6��5�5�<vDݷik�����8v��I�<A��]ɺ��U�9t��盵t�OS��]����5��{j����r�s�n��d7�ۧ[��:�)&����]J���'q�uv �te���B����6��S��s��ؓ��z4�q������;V�H띮�&���{�,Wlj2������Ƿ��0�s���eq΂�Ms�v���9*g�]�������um] v�x�Y]՗OX�粙���K��.��n%�竌�Hq�6ޟZ^]�gnq��n�l�sM۵	$.⼇	9�-�^ڣ�m�<#���N��e�d��qZ��W4ƴl���s9E�}���Mm퓴\k�c�7��ηm;�j�^s��k�8�:�ܝ��.'e�����
n\Is�R�Ur3��n����BG�eu�g���} �ۙ�T��{�[��g�CV�g\ݷ�4��{X��.�s7nu�fw��Z��ՖnL�G���u�u������T�=�[��;�L'�p���D��ú���q��*�����mۡ:r�����<��1r�Ӳ����	.z�7]�a�=<ބ8:{x.3ca����j;7qnԗ<Y��n�v�\��r�7N�vM���)p\n���b4򀮴��K�e��A9��sj�l�v(�<�l�0���.�qcg��k�f;f��;\#���\��u�c[;؃t�oZ�Ҝ��+�`�$zU�1X����eݞ�l�i.=�d�{M��Y'gZä�
d�g���Y��p/<���q=���)���ݷ'���Mk��=vw�#�\�<٬Z��ϫ3gc���<��ֲ���=��w7�y���u�,f\�/k7kQdpt�B��/(퍞ݵ����+��q��:M�Pq�$��[��%�В�K���^�d݅秮�^��{q��;W.z�6�]���8�=A��#��'=�X6�=���q�a7k�r>��ۀ�lo!�qq[��n{DF�:�8�퍍�H�6��\C��le�>p�ɵ���V���n:˞�v�n�����Lλ��|)!Hn�*jxù���wl�w&�vOl�Wb�z��q]����W�&�cn�ŀ�����8s�m�t5���i���ݷnX$ �u,�c��a��g�yݥ���j�-/9�������#�-����ݫr�V�ke�s� �ל�gc{\=�W�Z��s'+쎦�����i�z��!��緇��8�u������V틂c���N'��[�>/67o7K���=Z%�{>�n����[���ю��{Z���L��Y��������1�x6U���'�]�Y��2�9�;F�n6y��곎bD�8�\v������`6x��/Y�+�>��;\D�=z�e���D�5�ŷGN�=m�\�Ӷ�"�m��>˝�g=��<F}��MIZq�ؖ�q狉;lS���׬�{$��۹۴�\�e3�zĶ�x��ԣkm��]����m۵���]n�/uj�ɽ�:�l`v�������ۏ��c>y�ں�ݷ[]�yv���q�v����v�����=�[m��s��ɍЃm�k�P�9ָ�rmu�JHW/3����t�۴x���Sh��О�JN2+�:����m;��n�m�e�wn��ɬ�]�vH{uҞ�n| nɽRs�Ln����&�}@]�N��`x��p�6�xג�qį��ɜ�Et�A�}�^l�:��{6�v��ݺ\�l��Ӹ8sé�g�A��ͯGV%�s��ڵi[��k�H݃���;1�:�v�qn�y6���5�Gx۵[cZ�*
��n�(n��9�8J듶�N]�H�7���Dm���Ճ�u����q�8۰���λ=�ɓ:��݈�v�M�`���+y�v�|Z�l��&8�lm�����GV���d�n�SC�κ;9�+N��,sػv��6���WWlF�1���̅u�Q���e};��˲!,k�[��8|��s��v�錘x.Rb���@;�<��i�͇ֻv9;x��� 2�Ĺ㞵�g�c�ín�Ӌ�<��gC:�	�W��Fxh���D���<�����.����+ta�x���}�Q���u�&Ӯ�6�l/j�u��ڼ������{ucs0N���k�5p�۲��t�;،��x�v����G�ۘ�6ӫQ÷�)�l�C՞�ݰO�m 	�;S:[�݅��
�I�� �)��	����l�:
�!�����[���z�=m/@/�Yҵs�`�:wgfT�=r��뭙�{vl��\&�Go#&I�(#P�M�ͣ�X�N�Y2�3�1m��6��<vݍ��[�$8�ؒ�v�i���;9kū��`1�\v7Pwk�=��	&k�lr����p:�ɏ=NSC����Y�ݽ]S]�\�=G�6�4�svJ�;!��걳�!������^�[7%��;q�:�wM��81UsEJ��pЮ�G�{����!ƃ���vְ1�qݥ�ۮ%���GNq�`��gqU��uvwj=����<���+]�6�go�4�3W#�q�"]����ҽ3���m��یe�U��� �n�7Z�s�]&(�^%�G�a�tp����p<f�����ؓ��i��1��q�kە�9��Z-��-��Ez��m�=�<�ki�m��rX2��=��ʾ)���YC�+v��]�&xӇv��\,���/'��y��GI�m��.i;]z(a���.�T��x8�[(wkAo2�mv���m�ua�tp;c�g[7l����vv)t��lb�����]��
[�S�[�z[�u'��ֺ�f���v�Oq7]��v䲽��Ƕ����Qƛv#��v��u�qv�uPŤ��_)f�v"*랍�5\T+=k���ZE����H۷��g�'s��������t/u]�����۫���:^ݺ���5��K�[f�N�EG���8��R;\�ʒ�W�77lr�6��l��s<�n6w]�m�n6�z��x��1�q�=��[s��u�1�J�S���ێp�sP��mfWKi�/��x�7N��[q��m��e��n�2s̳�;u�\v������.��>�=��v;W��Ӹ�{[;7��,#ۂm��!۝N7]\�v,>9�%��ٖ������q^�q���{�ުt`�۳\qM�^[E�mv^:���KS�p�˟o0c�m��/e�u�.g�=k��노�����r�v��Q��q���j'��%��v�� B4\
ܖXKѹ�dK�D�cn9e��t�h�ٶ+��֎wQ�&Ջ"��][8��8�s����- z��ٺ����/n��a��z�yxva�g�^��q��l'������*\(`s�x�D�f��j�{P!�;r��L�z���1\���sm���u����H^�6rl]vy6�!���4�Ts�ь<��U��waY��J����XPc[Xr�.Rx"�Ʒ]�4[�X�k��`7O�����۰�݇�[6q�k��y䋳ۜb�11�S���������Ofɭ5�m��9pw�7;�ݝCv������^y��%9�n��Yi����{D�i��KĄ(�6N66����3x�SE��d��f,F���A=�euٞ�ܴ8��eگ<�ηdg�;��;a���1�r�Ů��]�Q�Wl:��OXԎ�#�Y�GRW�����}���F̙�{u���93�p�;�y팚�47�9�k�v�t��nAɋ�7�L`���\,�)�5(ݸ5E����E�l^����ld�Q ���ݛϋ�0r��=Y��WWl���b��"aG����>Z�4t��e�Ag=s��Ѧ�R�^3��5�gGl�l�;�8�l�r����7\n�p���q(Vɻ`��v�����-��5`Z�ݭ��8E�n4a��x�۫v�ۍ��4r<S]���ԋӡ��c���m�"�{q=;4a8�K�4�DD^�]mΖ��g�ݣ��r�vǇ�;��\�VT��]t"sՎ㋙{oi�N�v�d->�n�ѫuF�ܼ=�1���ی��e������ѫ2�Gn�(��mў
:�y{ֺ"�[��@�N����i$�y�Q�qsv��:�cK�v�J�۷���.f�l�x����.|[st��u���]�3�e���I�`���:w�.�C�k��Z*��4r\�8�y����Ig�\2�^�_����V(���T�2��ib�U�E�j\���*.+Lh�s
�he� ��@c+C)KJ��.�-���ڲ�n6�n\����֥p�\�)F�c\�Z�
�\�cDTJ�sR�R�9��j�b����Z�
c�Rҥ[J�8Yr�r��mq�Z��"�lFW2�FE1�
�e�Ȃ�)m�3�(Ѡ����̕UVf�c���2�����6�R� ЮW)�ffP��̢K��0�1%UEU�V"V�V�QJR�T�����[F��p�9��9��P��<��Z�UA�Y����W�n+s0DTƵ*"��\���������UU[jU���5���L�1EAh�6(����1Ƶ1R�cc
�kr�L`���e�,PbV��9\�Um���8�q�5����Zʊe�D�(Җ1�%�lUTL�������X��\�`�*��jUs-£���G�1�(��iKL��Sш�j�6�\��Cd�M�7��ul�չJ���=���c�\\�Vv�����n7��H<Pc����\���7�~�����6�d���i�f7mtD]Z�b�;������U�.��f&Ɲ�r\Ƶù�p�ϫ��1]�P�ݳ׮8�c���@�:��=u���y�{>z��l���\���y�u�m�vw;n���Nn��j�E���]���l���s���4��^;A�X/E��'=�\����z!,]���#�3���W{0':����ϡ��kW&�cp#�x�;]�q�W��I��3�RfWF��.S�88�b�<k�\m"F�c�c�j�x�h�Ǳq�fN�ם���my�ٗj����돭���wV�֜��ö�S�����	���G�m��7%���q.�<k�gtJxnve�x;�&�;�3�&��x��<�Uu�ۋɓM�휀6ݽΞD�ֹϮ+�v�v;Ry��r��
��b�#��S��xʇ-mɮ�Ļ����m���J{c�ۍ/E�qv�^ܖ�..��+����;=�3fG\DF�p;�����Wm��1#�85u�X�L�:�:1ӫ��(��lӥ�[��l���;:����x�@t=�y��i�u1�g�[']m`7h�iu�Z��;X��6��msX�8!�ÖֱX�V�gan�I�ϫ�"��d}s[L�{o�l��z'���t��6�Q���ͬtョ�c�N�����cۏ����{V����n�W�\q�snN7I��ZU�qi�7/[y���z�X��n���w�{����Csu��Qi�1���K��/�OHy��c�e�8��=ô=���ź�'>���o7\e���_C����k��ιW��.d8�]�u��j��������K���%9�W%�D��(c��8��t���;G\s�㨜m\6���]�s1��6:�I�F����u���V�l�gV��Z����<�G�ѵՖNچ�]����;�c��)�E|��8瓱簇'gÇv��P�3����!�2��\��LUF�s ̦bdÍ�/(rv�m���8ݸ�;m�9;�</(� �ݼ�۷�r�'�0m���<�g9��7*m�< �s���v�{!�=�0�����y��ͳSUqTn�R�LKL�96϶1�{ ��p{�Á;	����L�d�2��n ���?��
	�� �j����͚�P9����#�3�Z�s���|�oP�H�Yj A��J|d�̆|X��F�Y��+tWOH��T	$=w|MXncY�Wvq1R�!����V�UNI�UĒYq"�\̹��p ��ު�$����8
p��6{/w��E�p�xO�u�"��!�'u�My�{�nw���W}��%�w��CE�!0���t�\�	ʻ����F����͚��9W,n�����؉��u�<:�Db�p[��:إN-N�O��Wmd\�<P�%��PE�؂����o&����]�ܪ�$Yڹ��E��UxS�XH��s��A��q#m��!C0���f���3��v�b�����3R��t��G�EJ�9��Cm���x�%���yr�6��J�ݓu�b��{���Ns-�[���PFmu��z:���;�x  ���������z�ݴ>}}�x<M#�e���0\B��'�d3�|��U`�ŧ��[�0��f�I7�}TH��{�l��ÇUκ�b��f*l��(pM�  ����P;��U0*��r�x�t���`�m$h�`"�z���w��+}5 0�ZH]]U�@'ۙ�Trx(��/�.X3`�D>O,\�n�:�}�g�Oj�������ޛ,��AS�;��Xa&b�<v�@�����
 �'y ׭e�v�ߕ���,��R��]B�\��[,�QpJ};��@�	ѓ��	��������j���oU|D,F2ӊ�tW����9Dl�l�
�������>'��αht2ޑ�Vbx^�9�ih垦���L�iY��2�S��he��XV�[��^8�
֏m%�N���7��j�ID[��s`JU�v��T�h�oU)�-D�%�Q�9�^�DrX��)�cf���� >���B��:^����y<�x�!��}yT MJ͆�C1�DU{\�����9��8���W&�g��$nf�
$�{q��(��Y�8۝�F�i�!.^���v^��Ӫ�М<[��\XkY�c֮�䍗;���h�6Hɭ��I���I�܁�l��D��NUQ �wt�/`�Xa&bW���1��b���|�Q$�ޚ�O��gy5��ח�&��e���j�p�,��`����:YY�`�j��h�x����������T��iZp7�D����I$�On$����]k�Wӛ�؏J#o3Öu�f4Ua��0g-(���<2�9�.�����&�{�m,������w ��5Bk��A�4B��1ؑ��d.�~��D� ��QDCE�f;,2�����a�{P��$9���|p��`����^4�q��EGܪr�:(��I��T.�}'-�ݻFz�9�� ���<��&ݷ��χ��C4a�⹼˪$��!�Hʝ�w+x3�j�\��P �x�����p�E��@�dώ�u�}וA�wq�t�M�(P3�ފo���xT�l5-����p���X`�b�<r�@d�r��h�Ɏ�c�N�>$�yr ��=�D�祳�0Pjsn�����-b��i�x�`�ܲ>ڝ����1�R2�c"� ���>�g����Ce�Uɽ�Q'�/�����ю{sDu���rT(S~�$:����7|��x��v��3T���ٽ���P��.l2��3�E�z��-Y�rRΈ�c��ִ�*�w�$�����Mfu�Գ�;&I���Q���!��Ol��S�Whc�x,t����g���o]����Wr�-�ԓ�`ۢs�1ڎ�ѹO\'�'SE�n�tQ�񰞧��L��gG}\�K��������O4MV�.���+Y�'������[;M���kc�:�Z�9$�4j�����'�{u�D%�c)�L�96R��ӛf�Ղsvxrv��&�q��y�\��:�Sϖ�Zx�kv����w�Oj����?~h^�d�q�K˖=S�"�{�Cz�ԵV����{㦪�0I�{*�>��}8�0��u�AG
��e��&��3�|H�������D_'�:��̱��5�M�N<�h�Kl� �f�Q'�o7�P$��e�[!�;}I�٠H$�ު�9.#B,0S2��T<#s��P�j��{�d�
��A ����A��'m��DЋ�&�W�k��R��l��4�a�ڮ������:��p��MM��4I#�w��><_d��ji�	���=�@�.�c^&�]Su�]��d0��<n\p�z��68�;���/�oͶ���zo$P9{�4	$�O�$X���F�*��� ���%�{M(A!��.$�}���p"X���3�k�[b֩Wn����C�{J\{�RH^��*�����f7�6�-�l�)��V����.���s(0���(�]ܳϑ�$� s�y* �l�ϣ�ն2ɭ��&*�t0�1�n�����99!�F=�	���S��.��:�H�Ӓ�)�-ǡ��D�ɐw/��w7h�$�W\���D�}@M^�k��+��c]�����V`�%�
�5�!�NM_W�;���&�ga���kw�Ex��`���2�dK�s(e���`�����L&PRn�u���b1�i�d�u�������or��~�|Ͱ��$�we�Ux�g�D��FMwP�o\s���bfσ�Ϊ>ï'̍���I�����J��~T��o]�׏�s;7`$G.yAɭ����`�D������@anL%`6SE�����d��젇��k�(�����|�Ϋ�Ǻ�In�wE�����/_D��Յ����h��<�,��+s�-�����Խ��s ������بD��x�fo��u���	5�U�J�Q7	��>��=S6	,��I �����w�ԏB7nE��8G�D)�0���Q-�d�۪$���FmwtNV�� =�� (��%B�ɗa��������j}mt�W�qQ��؆u�ѵ�.�pmn���9pb	�C
 ��$��2���)�鮹�Aɻ�E�oM���=1�5^s��@�����!&a�K�  R�WR��P��� ߻� gJ���)a`��T�B�i��m���.���I���H$r�Z}k ��Cٷ�L
�O�@7�� ¼�J)@`��ν;�:Q�}8�5��� 7=�B��:R�^ߐ�=MݴJ��@^_xw�
�`��zߣ��&ۛ���1�����
���(��3q�\�Rݓ�'9�U��~o��u]TL�,�b"7"���]P �o�<57��꧴b�K��w�$�/rC
3+*8l��l��*!g����4��ۍ-�]h��F{��A���kn}��T��\ϡ�`�[d��̺�'o7�� P�K�������݀�*U儗��KUG�]�%�r�6â2M�.q�5�@E��PgM��Cwmv�gz�H�1�o�E�m!&jGc~H
 1�7P�Eq{��q��K���n�z��O��,����i��h�X�Kg�o]6���y� +vo��<s���@�꽪����#�v�:a(%��-��d0A�ʪ�xwqM����.�O�<^d�'�o���zQ:.qF�U����k�5�w�����iR[�3N��ӆ'�o��m�����uտ�g=o,:=@�(��I7�N]a9z�ΔXB"�-�
Z��Kh���A4��Cc�]v�U�=sz�elk"ip�u�c�9�C�=����Ev�u��WF͎�Y�l�QC�cvad��)8:}�]v���1�["�[p���ٓ�s���
n�i�T�yd��
/\�S�h:i�=�ێ�Z�[s��N�k��۸܌cDK�n���Λ8�fZ�㚧��MW��^��f2��ƀ�<<ٰ ��P�ݨ{$��N�k�)����y�U����GH������k�A�q���˪'����Kɾ��YL�Ge��$�e�O�fq���D�h��ܺNt�U\�P�U�=�ď��
g:^�=5�i�=۳}*3���\�U�f=�*��.���Md�W��A���a�ꮭ� �/rC}�7�(�v�`��&a��k/�.G\�f�E�vH�n�C �:��{{լ8�(�5u,����zޅA�pL�1V�N��By�ھ�)%���p"dē��7�(��ު!5��槃����A;]��]����	�W^�q��h�7<�=;��n^��d�+�̓�w:��P-��x�w�'vo(Q ���P7�"���4&P:k��}�7�+�T�[�؀�Mª����!��4W!n,���|��SB�c��8˘CN�N)��,�HQ��L1:�(٠��̳�e�i�����`�W���E��5=��B�v�$ }��@P��e�/� �P����aНѤ '{P)\��r��y��|��Mx�}��@KE_c���B��]�]��)�i>1�{4H$>��_@3���]ˡ>�mW�^H���4�eBP�jv���M��-tj���Zh
K��� ��y*�f��*3�����'2�m����}�\==�t�W:�(5�:;=\wvŵ�����$ۂQn
%�x�M�W�s�h	$b{����w\��ggU|H���K
����Ki� ɍ��'�8ڶ}��&]�u	���W����@�l,oi7
�#�f�"j��MB�a�p�#z�	�>&����
�%�dݙiC.V+�݌W}�-r����gGܐT^��7�eά-�i2�����.�v�Q.wf�e�؅�e0o�N���/^���	�|�3���4�2�F[��u��p�|Uvܭǧ�ɴ�-��b�d|0�r����ueP��Ò�ͫ�v�b�ԩ��+VRW����r�\�wj7Ƒ�F��Z
&�8a%��(OLE�sv�<g!>���,#.����IQV�.�@*���[Ӯ�i%���D\�qۃh�vM�X�{g��)ـ�V��E��5&�pM��`�;�!d��p��oͅnU�������Mm�
��VQ���D>��Z�&	Z�3��m<c�̗�]_\֘;���#2!Ɣ�8;�8�y�;x�8���% ���F��Y�Qw L��kQ&�l3�`������������vL�.wlY	,��ܥ(�k�g���.��.GH"]85%̃��O!&�ש��g}�]�m*;(�
���H���ƶ[WR�2������j[���k�}ό�&-���gZ�9rP�=2U��kn�+ᳱ��w��f6a�V�h��9-B�%�LѼӶ��x�,7yw���wYβ޻)���u������M��0a޽{��r�o�3�N��G]��5%m�h�P�4���w:���cbo��M��C��#;����nK׵\��������]ֺ���Jf�κ"!fuN"�eּU����ձҲv%�U��Zmj�h��[;�
�$�n�J�j��[��9L��L\�1mJ���9j�mj0QV�-J֪����-rŕ�3FVR�5�IkV�R�QATR��������Y1�R��l+Ze�-�*奣R�Z�ʢ���1ƅej�72#l-,�1�m�1��kKUJ�[K\LX�m\����3+|���q���7v�|�_e�1��U��0�E���Y�R�Q1�G-̶�e�V�2�p�q��ٗ2�,�VŴR��YQp�aZ#U+J*�`f%�U���[�!`��ѱ)m�-��-�J�h�9V�1��ȩEZѭZ�Z-c��"U̸&9�$�[�`)�.V�ʥ����
������Q�C0���)h����r�-�֣Jуj)hՖ5�aQZ5���b�U�Z6�Z���lpg��ʸ��q��*�\��Բ�J%Q��`�%E�U-Ln%-�̩m
�cD���)nbԦZ�ŋ+Kr�J��p�+ZR�e���R��ilF-�U�jYeE1inJ+�Җ8��A*�����|O�󺨐H8^�����- �,�b�0h�sf�z$�����W�P���>��ˍ�ۺ��*�U]~�J��h���zU@�˹`�����5X��{��s�TH$��Ksf���\/1���P�d�m�n�@]���Bط����.�^˒N�NB�����~�|��eBP�k�n�@6^�H$gM�C^�[�_��#����J��d���z��l@M80K�3S�TAe;Ձ��l����4H���D�}�7�^$�
��<�싾��ͨ0 %�8rd�m��P�k����	q#��oީ��܁$���Q3T�Zj2`�J�7��y.G��衫�Ok z�� s�B���{�9b���q{\�fc�&ʬ�c�J%�S�kn��cZz��4�Ұ<k�%%R�=*ռ���Ο}�M�]�:N��!s���eԶf��[,��� �m�Q#ow�����DL"uOt	'öo*��]�̂zq�t�q3�H� ���1��E�P0�#v�ÌN�C�ظ���C����o6��E~�?�~��>zS��۹d��7�G�]�uP/VF���n�C�}7�^$�n�i�q!�����
0B}�v5��z���@H���O�y�T�P�(I@��ݦGc���`&�%�x�NuD����@P)�Fi�׊�������^�x�M�oU ��% ��8a���ڌ�6�qk$���>���}�T�\d�Ϸ�?F��{��x���6��{ ��Sq��J7!���i� >���_ �s�T�)��|�+�͍�	��F����E嚷q�{N��I�l�����g.����(wA}uݧ�����m�n֌o0��}u��9r�=�X����B�$���a�i�dמ npL�q�e��U�gJ����W�|�!'&���z�n����GvMh����3�8�W1�cu��OiBB�@ZL��#�T�\MxCV�u��n�ۓmmTۓ�����銴vc.�jy����\Z�\`��۱�ɮ �X��՟9�vz��.V��Y���h��{uN���i��;�_G��QI�{uƻR�$"î�-U�Q��e�	n����*:a�G3�
pL:�KG��& Cl�v����ϻڇ¡�/D�ep"\2��/���w��6a\� 1��8x�܆:�e(�!��c��Q���<���h���Yr�
�t4�o6ӆ�q�����P'�Y��d�7\�k�ھ�'ǯ�����d���D&�Pq ��.����wA�Y��_�����>R�ߦ���`����"�n� +���$�2a�L�{,��וK5����dUÞ�D�9Y>`�����4l�Ȅ���{K��W�������ǐ��5�]՛�vӅ�r(�i�	����	�P�����sw�AT8E6�U@M��8�k�8���H�}�D�A����)J� [!��.��ѯ��J�]��s�5���<v�7�@:�ڧ��Q"�:�_*U�]��,*�6���K]�GL%%¸|��1f��8�t}�z҃&��,�[�( +�9z ������y~%�1y�� �� 1��#L�g�#&愈$�Z�#zb�Q>:v�X ����%��q	q�����۾����x��
���A��m�{�VJ�<ʠ�n�"x4�jn" !��mss�F�>�}���g7״�-��� �'yU��S0��1���DX�@��n+��	�Ş�2��ug$�ݥ�1�GTG4#n��h�i�u�ק�ނ�$�2`��f��~����>7��4q˄U�DUB�q$l�ܰ@'g/��i_Bj1��&�=��pWqKQ�y�-A�(P�8�T��$�PU�cY�ϡJX,�!Bp̃ݹuD|wszk���eT�۳^0�e	g�=��Ԫ�a� �Tq�b0��1�嶮ոX�TΥt5� �(-�x*$�xō'��_�ٹ�p$�3����y��Q=-|����T��5="E�x�)���z� �n��P$�����ehLW[Pb2VϢ��t�Q����N	�!����`6v�|��"����茛�ogt� �;y 9�ѻK^m
.���1Z�4�>��E��=��^Zu���t7n{]hwk��n���jn" ����Q�#;;��I$��D�^��4����y�T	���P�AP
P,�A�����n��*��y�N��wH�N�����C�MYկ�©9�a�υ�>*�wB/ѕ���8�����AH)�����ɴ($�PIX]����}�ϟ����_w�s�:Ñ�aA�IS��w�8��VJʐ_��~ܞ	�
k<���:d8�!�Dx��vd���ȫ�}�|�ԅ-7���󔅥!Z0+��߷I��R(�~��8�>|��wX<]�;�x�z�M;���`����̒�^c3.`�oڐ��Lb��Xe��nh��+E+wk�V$U��g/��u�h���'�%B����ݜH,8}�-��N..�5�_!������i%#��ܼ�>}�ң��og�z�%@���~��� �����Ct�B�������x���������8�KR�i�T0��y	���#y�lr���n��lOIg��ۧ�Wgll\��~��2Kv\�vk�1��}���e*A}���2m
��RV����0�
�X�>�}�!��O;��g'VJ2�_��rx	��wό.��eu���ׇo�����<��k�/�= ���g���!Z0+gs���O
�Yb{�}���q���%C��~?S�R6����}"��>
�m�����kZ�!�+����x0�K���;��9�JʁA*��o9�ߘ��߼�OP8	XjA{~�ہ��� ����>�6|*j�t"�"
*5�,�z~��E��n��#u	W� g�%e+�����ɴ($�Q%a~��υ����$y�w}"�����ߧ��3��O�Y,ew~�������9��ff��e@�Jÿw�0(ԅ-�߿wg��>98������80+���'�H,>��{�x����D�w�,�dy�W�k�*̛��ȯ���8)�|2�q�KqJݵܧwE�C�]�k}O��SM+{���]f�[8l��Ŝ=������1o���b�~��ć2a(e�	��uc�	��7\�n��ݸ��u�#Pc��\1�!�ûX�1�j����A�x5������^[ZNu�!���s��ZO6]�읶M⣨6�&n3������6̻8wn��^�����ْ�m��\K�f�ptv���%v�+ ��호��ݎ5�u����zq���Y�����,���K=���[��r�a/��m}hӸ^���˧]sǭ����v;E�r[r܈�!�S߻m�t��tf�3?�x��a_ם�a��i%B���}���'P,J�`ϻ��d~! �٭�!}�oa�Q������A����<���Ïn����8�!DA�!׀�(�u_}"Ȳ I�ϧ>�_{�n��������2m
��D�����~�a��aRQ=����ĜB�VVO~��y�f��^O]��@׳�`&ۄ[��%в<	�里�RZ�����H)���_d����o��� ��@�|�_w�Ì��YY*��~����>2�0`0Zn'�O���#+��}=��X�Oa����(�a����gq���Q*�߻� q*AH/��}��*^��㓼<	������Y���7�Z�c���p<N	7���g�ed����~���C^g����|�~&!ĕ�3�s���+T�����N!Y(��Y_oy���M�y��s����}�<KS˖�W�5p�r�Y���"^Wt��֩��{S�qv���nq���oϝ�݋t�f�E�V������jB��~��9HZR�
�s���O
��>~�z�mߠx�bg�s�É�d�T77�Y��>���>E�fExY�O���@D{{�}[U�]8�����o^@�),��6I���0�hy�}���T��0Ҿ����s6K;Sr�c:qiSnn其,���O0�:�7�Hy��~��3���Ĩ~�����8%H)���n^�<	��rs��S;�N����<	�D<�f'B�C�Q��>�dY��VX�_oy��6��
$GÜ��+F���(��L��|4�#�������ݜI�+%eH/���ryH{��E6�"�DA.���𺿺@�}�tʾ>�Dx$�5�H�)JB�`V��s� i<@�A�������sz�5��s$�,d�T=����!�%atg�q�a�]M]k<��x+����x�i ���~�g�N�6hss���a a�}m &k��s����R���?wg����H�rl�G�ĥ�@��˞��R3m�K�1�v��s˔��%�ٚN�9�hE��sR)0�IC'�d|G���#��d��%_>�g��B�*G��^=�ׅ� �#��v6D��QL��:��7Ͻ��$������~��D��(2�!�jA !߳d��$x=7^O	�n s���[HV�+��ϷI ��>��~}g�Dx?���H�����H,:~�+�wN�Uњp��a�¿�?{���
Aa���ݜ��%P(B �Q�FtIN��_*�XbP�×�(��6Q�VWefCS`�R�f�s#8^�5�gEI+��@<�/��ZWW�G�ܴ�=�r��}+��&��m�%"�ԅ,m~ xyF�~��5�F�^����� Ґ������6��8t3	����^u_�<Ou�_ϸx����%w{�vx2mT(���|���C�9T���~��{G]��_��O�d�ed@#������I +��!��q� q+yϿn08ԅ@�����>������� �`V��o� i<� ��|�߷$q��D=���g�'�����{(!��1Q�0��e�..2�����'=����:��ֺ�kjǭ��9��
~i������2�v|#��(�a��~�g�J2�'���P� ���Ә7���7]�|(���n������<�ny�^<���thі����ě������+9�x��}��9�{&�.���6�IP�+'�s�|�paXV�~�݊#��>�>G�PqV=W����m��a��t��D�pMp�
��n�H�&���v<`V����ݞrR��(�Vw��d?v����� G���s߷3���d�X������IXg�s��]3N���80�o;$���b��sÈ��>��a�H(J�a��|8�Xk�_^π��^[��Q�{��5r����QO���fnA�.h����f]�u}��M�j9V{E#���x���k%b�!�9[U�IԒEG}���H����+}��wFn�_f�4:\s.�א*x������'
�'�y_^ȯzHP������x�Xs�����0�(¤��{�{��8!Y++%_׼�rx&�>��Ϯ����{��22F#bM2��!����ň���[<�gT�����6;b�~�~~��Eu����O�:%a�=��0+R�>�����������O*y߷|�����x��s��gJ�2T}�{��8$�,��_sYL.[���g��Ww����a��B��5���{{;އ�<��{�x�ѕ �_����@�J���
���>�$)���*nBp^�O���q� ��7��$�ѣ-����M��}���@��%ed�o��g��B�*$�7�>o��|�w{���aXPT�=�����ND+%ed��׼�rx&�5W�O��MD&��(��o۲T��w������`zԂ��~��g��-��h���~��@�x T��Yb}�}���g���F^�ƣ=�>g�D���dJ�?p��k�th�8fn0�
����m ��Vy����d�����~<�~�@�%@�}��� q+�H/��}�H>�a�������X?;����:�����M�˦�7����*�b�����[6�]����7j ����@X=v�G�Q;��{#O;�:�	*P�E�]���iaN�-����͋�}too�X���^��ev��7$�p�ڻ��O����٭����=�VQ�F��=����/�p����,Kɝe��9� 5��4f)A���c�;��4sEpM�v]p:��D�n�����;��۽H�0*��K�.�7b��hY]JU��"���Ⱥ^|�>�dU�y9�z���K^ˠ�U�gv��Tx/^;�>�����Jj#dky;��j�]��v��I ��Y��U��z޷�gon�t��]�.�Z���rm��ҭ.i��|c��`�����m�c[�Rh������i�&���z�u�,�j�+Τ�6h���s4�S����T�2泊Y	�J[�Ga�����;{�aوuE�I��Ի�c.�t��D���*Cna\Mf��8Nѓ����]���6�C�kx�+%������ɕoS��/1���t���e��Z�`�MY[5�Ω�ٶL�܊�h̜ޡ��$:�*�yp��.v���L��.=�v��6� �v�(ƻכ�Xq�H�C���sA��Q%��R
�H司W+aE���OE�}կu��4���51K�G�[�t
Jgu*7}2Y��VlE��E�U�3����	������Bd;��Tw� .:�԰vK���x�ۉ�l��{�K�p`��;��w�3�՚�Jb)�DI>�j�E�anNC��Z	۩��'=v*3c<���xP�[RեKb���Y���*��Ƹ�Z5rܥ+iJ�h�#h�\�L�)E-mJQ�\���J��fH�32d�.jZ��ڋR��r���T*,���Q-2�*&V�[j88��e���k���m3���P�9v�πˇɻc��v�8�r�XZ�ˈ���%�V�67q�
�������&W����Z-a\�e��.ar-���em�-��=��<�yM������®ص�cr���\�[���Es+�*�TU+mihV�8���,X�&[\��������Q�mh�*����iD�֥�ir�7
ܬ��n-�ƭ��`�Z��m�ڙL�嘢���[j�[�V֥�[EG2QqAKmF�*U���fLl�2�*���K�r��V��h�5l˙1(���j	Z�1�Z-�s
�nS��[��	�m���ɘ�h�r�0�JTj*Z�Q��*R�Z�J%�U��QۘTȶ�Q%mm��b��lQ��W��>��t8϶�ո��tm�S����kr�Y����e��qۄ�8�Y0y�]�T�bDn;&�ڐ�P�ͱ��;��s��>���e��Nۭ7��y1��u[ljZ����G`sn�c��K�.��'U�}Xݧd{��k�v���c]�\q�Ъ+ ��.q��e�t;WQ���-�l���z���ͳ3�ɝ^7g�����ô���=k1��v� _:�j�@̀�#x8��[�����x���N��r�@nzf���I�.���.6�;��˗�����/���.1�F�)�e���l�<�M��.�L�"�]�z�ۀ�k�9x|�ջg=*�h�u��ˮ��l��s,���F]֒Uh���F�S���E���3rS�nG�t�^w�Ch6n�muI����y�^W�n�2����˧�hn��cjv��u<7�T�>���&Bd���s-�v����=�'T����g<����=�7	gu�&�v�d�Y��n<�^��x����A�4'e@[Mq�æ��b�ˆ�iݖv�X���mY��g/<m�9�g���;q=�^R�]˫�i&2;�m�;e�j+sӽ�Q�.S{v۫n��[���
;Fd�6Cu�ݮ�u"����m�F�;,bzxy4�Tng@��h0;�h�Ș��mu��f������wbr[�:�͊����'����Җų]��
�W���^[N�]�9�v�כ�4�Fk��l0p^�L���u��5lk�;���^N�nL򹅊{-�Ľ;����qvr��wW]��p����'>�/�Z2N�t��ql�mn����N�{p�qb����۸x��l;���m��,�Z�d�������^�;���ӆ3�9.��:|l�B�Y��mn�f�]�w��`�NT�uKt��v��4�]��F�������<#�����.8��*ظ�c8����an��he���[��ͬ6]��^v�2Fa��CL!��=K����Tf7'IN.۶Y�<�vK��,��t��ո"7dH싛��7�M�ݵX����.�ힶ�-�^���J����N1A��n�"��:G��Z��y�5�z���^��#B\>�c��ƫ����k/g�cMun��=�:�f�.3�y�Gn]�r3ڗ�S�q�����gm[��V���z{Us��kr�_Y��B\w?[>���@X�&�e��md#tsd�k���]�Ų�^9��]��0f�����C�.9�X���S�{������
�J������<d�IR����C��淼����n�o!�Oɿ����$�B�VT����ہ��{��J�:@�]^�!ǌ
Hs�y��s����~l� ���h����}�$������<f��"<	 �}տ]����@���F/�y���?4�W�#���}!��i* ���}�gĂ�R����n�ug�f{��@B> Q�Pk��>�7H6R�}��{�q����$�a�IC&|dz_}�,�ϼ����5��>H,���~ߛ<d�%H,/�=��C�8¤}����F�_f��|��Dx�P�������I  �� �A��T	�n�d����G�	 ;;��V����˔mX�R����4�R<O��߷3�">@�Ȁ37�Q��>�����W�ϲ���2&7Y��r�MQ��=/&�v��4��{]3=��i�a����v�\ɗ���XW����x�i,B��
��y߶r3��e@�P,�߻� pJ�ֺ~>}��>��\�w���A�!m�v�g����P�s	��Bp]x
�D��{�vq8 VVJǚ]��u�]����~A�P�w&:�T�T��m��,��;�m�����ۍ$��R�9"ȇl�1:3f&�N��֌CE���s�����s����?]w����*Aa~��~�a�°�¤�����dx�Y�>�w�i�����}�/����{�D���`(l��qB��F�?~�p$������vx�yHR���ڑB�k�bn���g}���	��w�Ì�%ed�T=������|�P{n ��M�x3�G�O�`���ާ;�t�˚��T��T�
��������������|8��J��R�����f����H;)B¦�'�̓�^�;�R)�i(d׀��M��g�������l�d�{��q�~�CV�y���aXQ�IS�~�ݜI�
�FVJ2����rx�@����>�vw��˧5�3s������\j�n��Q`�ŉ��w3e^'f�����5q�j���a����Ã�jB��~�ݞp�-)
сZ{�� Ȣ DE|&���QS�f�8�\>�p�%H(T=����ĂÁ����к�油�C��~�66��"<�򌩝���.���������|*�P/���|8�Ĭ
5�Z���|J��g�0�2���+|2b�|,������ఙhD'׀D߹���>@��%ed�����d�	*%`�1�?{��{�\s�y�[߼��(Kq�/#=��R�� ��ݷ6;gf�F��ᘜ5�c����y��߇v�p36�$�Uo���3t��xxyUN��� ��aRX����q'*Ad�����z�� _<�((l��p����O�M}�Nܽ-D�q��>
#����{��JB���}�P6�S��������0k�[�xC# ���w��� ��{|��L̻!�������G�>_fH�{kO�#t��{�7v|�Ԩ�|�@�J����{��j�
A�,=�{��Ă�5����~�/ÿ?������/���6�ܽ��=����Gӷ2/J�ɚq�?>o���V�F��NĞ}������YFJ�2W���G�'�Q%B��/��߼�q�`��������Dy�>�͑dz���2�VW���I�O,�?q�3WkN���������G�!�_ݯ��׎�^w~l��B��
߷߷��@�D
�	��߷3��R
;�ؓ2�����dȲ�|}C��GZ[��g��0���A�T*Aa����8�2Pe@�T��>��{~�v7����q�J�Xk���P<�m!ia��w�Ï�3]��Y��:�8j�"���g�,���o��� i�J�2W��sG���($�T��w��n0�aXV�}��<H���}���{�����
����ɧf+�.W��ii�/��B��
���\��~�K��w*+�[ỡ�w��*Gn�^ve6�R�B�#;Et���&�<��x{��ߌ��ey|�ۓ���������R���Aa������x��R-���}"�!�ϳB��vB����>Q=u��x�R������J�2T�{�@�<�������n��e��D�sF��8Mv:ln�<mֶ��ot�y�׳{zq�XA�`��{@"���O�|>>ʜ����T�B���}���'T
% ���Y Y���u�ٸڟ�8��y����t��ia��}��ǃ �G3�E�p�I@b��`�}S�H�/� �����;�/�D���3���<�����i
�����＇A�IS����8��VJ2�\�w����w�U;��M+{>��� 0~��!�-�ׂ��J����<`PjB����~C�/!���&�sⷩ	���<#P*AeO��~�8�Y��P����vq$�3����a����f��Fynd��u��&bW۾G������߽�<d�ʁD�?}���q�X��w߷[\�?o�i��
��l�υ��#	��I��p��
x$���{���
��YY+��~����@ϻvT����� aG�n~���l+
*J'}��8��VJ2�P�S�πd�4�E	�����WN��y
�C6�F�^b��
y��o�M��8��p�#@������Ʊ4�u8�'�B���F�G�ruN3�����������ʵ�ύr�V�t%��9]����F�y�Nf�c���`7k�T�uuY�d��ͭ=�䦮m�\>���"����7n���c^�X�&`���k���� n;A���'K�t�c��9[�O��{[�F���g�a.',�M���<NѶ�D-���<�i�+�ؽ8��1��<�ٺ�U���\]�4{�1� E�x���},�j�א�[v3��']l�����n �Hb���&�)6�B? ?�����<`Q���w�<�!m!Z�������4�>�=�������bk�{�É �w���<C�J�����(�\��Ӛ�H-����d{<@DzV����.{@���dԍ���y2�T����|8��*AH/�}�~��<
C�a�.��v��Ѿ7n|4�>5k:.!�NAb��~#����8�Y�J�_�}��M�bJ�V��{�͟^�o�ϡ��T�������g'T��w߷'�m�g�x�5�P$@�|;~͐3�{���֧���`XԂ���9ݞp�-�+X���}�'� ���}�ۇ�cϼ�|�r���ACB�����9W�Fm�\S��#^G�?-�� ȟT�
���߷9���g���=�@�T?w~�È�
�k��n�t�JB�����ۇ0+����߼f����@*�И�-�����M8�uJu՚}���r�n88~�?��.��9���v�ԝ�����
��YY+��~��&Щ*%a��߷q�a�{�?o�~�
����Ă��+%_��ܞ&��f"~!C��@B>W�O�`�<)�dZ�߻Vn�b����d��+D���v<�1c�F�5�LW-�B-�� (��#oNر ��|����?�$�y����vy�)i
�oپ��$������ۇ,�"��=s3_+m�w��Α�$�,�~s�0�jkN��4��˾��$������������_g��y���
A`z��������K�'�|,���MZ΄��b�X�d �\�!׾��?s���9�	>GҲ�%~��ݞFM�RT(����}�xÌ+
¤�=�����No����s��c+%���[�rx�@�g�L��Y�7�H,?}�{��x��H[@���H���8�x2<	u�W�d�@�P+,No���q�+(�PD��Y��>*���T�*QZ�=��ƹ�۶�\3���D�:����N�Jcr�E��]}�S.)�N��
#��]|�u��PB�o���x��T
!�����d`�|o�������JAw~绁�AH4�����Ï#�O�����6��E��ϤY�ϼ��e(ܷA�;F��qVd�ޒIP�%ag7�~�a��aR"3;��dx�X���.{�>���Z��������%�e)�<@�%a�?{�aǌ
ԅ���{��R ������|
�U�nŨ^���I��5��Ŋ��`�+Z�i����M�[!�2�c��W�����R7��55�_q�H@�~����4���+��~�<g*AB�{����C�J��P|b���a��g�F��)���澦xa�#��f\���,e@�P/}��|8��+���Q�?l�������_�<
C�//��&x0+My���.��ˬ�f� q8	5��ݜN VVJ�2W��϶y6������7��*	+
w�9�!ĂÑ�IS�w�8��
�YY++��nJ"H����b���#P`$�(�����׎h⎷U�M۷���#[�o������4�X]f���ؕ��|�<`V�)h��������+c��׵�xFWݓ;9�p��[�w3�����P��߻������7f�Y��+��8�_����$��߹�Ƽ�}Xy�9�g�KP(��}����AH,5���n��
x!��fx}��|,�����Xp�Q�a��� ��E� |���Y+��>��d�%B���7�I��ѿd����O�G���H�=`�Y,ed������@���y�u�.jB(Y Y�]}� dW��䶺�����}���<�!RFo��߼����Y��;߷3��s����]9�E�v�Xc\�FM;{��j��sz\:�;��}��zн*�2,D��3T�b*ιA�nk?{��~��?�*�}�<C�%ag���3ژW53F��4��¹{�퇌6��RT����"Ϭ��Nv�Y=*�|H�.s�;�Ă��R��߷�t�aH�k�|,�>�V����d��B"��/i��b8ٺ-�]��*
�{l�^J��zD���� �&!8P=�,�#\�'P+(�YY+����<d�AH,)���^|,�#����d;��=de�wgpB�J2�����iˣ��llְ�֋�x���ﻇ�RO��l�U�| ���"�!��C�|i�w߼����@��>��p�8�R
s���>��o����~V�_��q�u�]Z�y0�a^�s�����T*Aa����g+*�g���������i a��Q���;��x�R�����q�����u��iCa��U�	�_g�,���c_��y���%H/.���M�D�
$�,�����q �� }����y���ϭ�.���VL���eyw�7'�6�C�?<�ʺD��aL��Aa����������ݞr��?�Gu�f�߾!�����$��Xs~��p� ����b}�{���u���W׳� ׿V�SW�}&�Wb��vy�zy������sXG��u5V�嶏R�T6�l�óf%�
\��r�����������dt#P�B�����)�qV��<uu����;��ۓ��ר3�.�����̸t�t�=;�����	s�[r�T�b�%΋pk���֋����I��zS�
���c`=v3���;l�q&�.月̱���n{c��Fb+�M�k�cJ �j7]�����꺜�t���nB�q���Ƽ�����n�v�v���5͸h|�Ofr�aխ��3vQ�03�Eۮ`��Z���e.��������\�L+���Z�!����l?���T*J�a���p�*� !��� ����i����C>���k���p<7H4�-�߿��8ߏ�EM^��3(q5�,�y����'++%f����w���Z��i�J�IX^o��y0�aR
�}��<I�
�c+'��y�����{8��n�=����Md�fkFx)���������?}���� ��
��MQo�<��#�@�>��}�q�+(�P�}�{���'_שBpP�4�ExY��<��@�';�/���{IȅID+�}�6q�d��*?~�����k�϶|���?n�������K�f���͟ �'�6[�؄��> �@�}]�l�q��� �_{���h}�o����z$�/����a��aA�Ib~����$�B�Q��������<�I �d݌��v�3HA�������@tbM����c�do=sܱ�M�����틵����r����XR���Xs�}�Ã�jB��}߿wg��-)
�}��πdW���[S5]��8���/߿}�q�+(�P?w��g�pIXP�F�s���53F��4����y��$� @D{UQF/KA��S���'aNe����m<T��mɒO:�s��b��P���u�R,���>�e�j���k�?[���䐀���9���d��*�������+X��>��%��Ps�('r���}>t�T��t@L�
Dx"������ȁYFJ�_�߾��d�	*$���7���段��}�=H,>T߾�vx��
�YR���n�+��A<�!�	 P!ϯ$��_�R�=�|G� ��Q��I��߾����+(���p����}a��s�����I��x���C�J��>��a��\�\�!�a^�9�p4��*J!X}�{���'�������w�ᮞ�Ă�s��� r%`V��߾�7H)�7��n<��;���ϠQ��
pRL�8h�%��9��V���uڜOgTl�;6׳�^޻�������&�0����su��$����M?�ʤ)�7��>/ɪ@|8?M�v���A�D� �K��O!����O^�N��A����>gz%�k��m�Ԧ��["	F���AG6��A�ٓ^��Wޝ��,��v��
-�\=���c��/v�!v^6�n���&t�ü�޵�n�ZC�w�����A�ѻ�}#].��^�8��,eK���:0��1Z���}˸��n�U�b	�2��(�la�ݭ*��n��Y�j�/�oh�p���,Tވ��L8wf�C�p�y�t�"�7_1`X��9D]u՗�;��Nh�],iĚ�.��3��6�V$���r$��
�ĄE[���D�@VJ��mct��:�%]ڷ���K��t�LU�\ی*V�j�X�_a�X5����wq(J����b!�55{��"q�Ktf��{;�r�T���z�{MF[�6#$;�91*3k� 5E��_�WWI�͔oj�_!sV_of\���tV	/�Ѕ�e�����*�%48l>(�t�%ƚ*T&��gMBJgvYVn\@À˨�u�p��e�g��l��O9��;I�o2�^�b7N�|a�ٻa,Gpv)�.�I4yf�n�����,s�y�-�"a�IR6��X�4ޚn�^Wh8�5�+�L����V���.���ߢB{�5T�T��W��ɩJP�,&��B|F�g"w�Nk�sFڎ��"��;��X�+]A�/;"Vi�uo�=޾ٷD��ŐK�w�`��3k7�9Lһƴ:BT�4&5��y��;�םVb�2�����־�R`9�x�M�D=ʔ	���|غeQ�U.�[ �a���*�d�R�
���]�Mâ��=W��!�*�����l��V&�t.'1�E�Әc�8�t�zOT\��zw]q��SD[m�)a���iJ��6֨���.[n*d�bb�k1Ŷ���Jb�C)m��VѫiF2ѡ���k12��c\-m��%E�f�m1�L-\fe1kh�em��û ��ʽ�����<o`�!�_
n�����;���U�8�v�x�nA�w�w��K�b�V#�̮S�*`�\�T\�-�Km�X�`�KSc`���g���n��)�퓅���`�8�ۜ'.9���p�s���۶8;`�	R�kZ�4E��Kie�3� cxɷ�ɹ���n8����`�7(��B�[E�֖�,�K����"[��[k-mDAƙll�E��h���UIF��asr�ƮU��.9h̴�Y�-JUF�+�q\�Rҵ��L�q1ŴՈ��(�j�j��mQ�PiFڂ�A�Q�����*Dd�T�6ܸ&-��m��b֕Km�e����Z��b�E�[D�Y�R��*�F��֭L�pZR*��4��KcQ��5�S�H���s��>7�!�M>�*�k#bjP�@a�yweP�˸��l
9�,��ݕ@�>��yG�K�l��y�̺�� ��L�X����D6�r����A��飹��]E�t� B��I _Ne
;w��#&§�W9h���EB�Lv�;xѝ��C�6V�u�-Y1�֊�k'R�n8^��(À�@P��\� �'.{*���;w�OA�7E��	[S���*�!Dn8-�T��	��ު ������W+���{r��*�gD�
�۽TI&�n�8Iy����<a�>m���3;��gv�� ��j��[-�N�I$f>ʠI���t#R�7�N�MX��t�tnJ���2�6h�H���|E����lvu�G�pX���@{�݀���ݧ�8䃭��y��f��}A���2�� _7w�8�]N*
A��&�z7k���{��^'ٵ_U O�k#�jM�A�T��ʢ|O�����;��uqai�s$�u�B��oO�7[!��;U�_��:�=��ba��D�Y�<6���4X�C�\�����י���|��ԉ��D6����D��MI6n�$\dצ`�v��N��U|6a
�:g.@d���ԩ�o*�N�Ov�Ux��f�e��K{E.�$��;(�z�P�S�:��$���e�I<�f;r
Sn�3Ă}���D�f�e��3��-MF�U]�S
Tt�s�̿�޹O��u� 
�肞�]�	��z�U �$7�X�b
B���AG'�@$�T&t�쁁i����j�H#�����Mx�n��[Z�B���Ɠ�kԕ�2��cŗLf�V1fa�N�خ]�6 ����1[�C����Q�:1�b�#A)����_|; 4���V�n�Ǎg�W)�`mρ��\Y�r/g�ǆ�0��D]6�h^�,�Fڗ
ݏfF�[���k��1ϭ���jp�y9З`�u���</l��h�^˂�pc���:=��m�����55�������
�cԵ���Cٮ�ѲN�H:ɕ�)ɹ���=�yz�M!��(ŝ�m�\�r�Ńy��g�v�\�����u�i�\g�mn6���t�p۬�����8��ֺ���Ύ�M(hÈA�_x,�ʢI��7�$/_eW��q�����1홮�'���ؒ�.!��'�{+(Q/�7��Ȉ}���	�7�$|�*��On˧�\��s��67���,��"{X>�y�B��so����kڻ�ڢI:f�=7ϲ��(���lAN��w�o�p�ǂ�IozC�47۽N�ܙ��i �ײȶ6p�@��B����H7ݽ4޷�H@�޸�H�=�r�I���n��ӱU�m�Ä�������_��Y����s���q�����'���vn��������HC�0�p(��d���*�$�^��P#Vt�HG]x���7eP���؄҆�80XuAwNU�(!+�C�y5��_�w<$0g]Z��6����nb1Ts�ڼ�q�٧n<�V�YFN�.�[�".aA��{����#���$���Ux�n�4O�6m�!.�0�y�X�b�(16�����yDwwzkĀI�.C��V�z�<A�y�({�䀮�l&��6l围�p���N�=s�~�� '��P@Pc_[�J͸TuLW�v�M�͈-��Cb
p��� A����~��8
��J��*N�$�c__)��w��w=/|�n����u�s=b҄Z���G�=������qκ�2��ٝ`Y$1T;8�@��@��5U}^� ����$l��O�ـ�z�u9�Yww6I#sw��L�� ؄����q%�,�Qc��h�)��$�ޡ^$3{,B�G��M�M��fk#�J0��a�ϲ���%�|b�nT9L#� �M6N4��Zf`�h˛��!��O��N�_��4+@y-]iwhss����L�[<��ົ������ ��sj:���_Ox��s�Hξ��M�{!��CjI������;C�� ����O�'�����=�
����H\b�I�
/�@s����M�C�Ok(Ps=��u�j�J��y|�1�nP��=5|4���Ƭ�K�;����*��B`7fv�c���h�C����RA�E�\��lpc��ߟ��|j�Z�w��yE��A�נ��z%��p�acw��5�U	���X��l�C��������^�jj�7�
�*r$A>�}�+�a�1�B�]�WC��A�(�͆�|Qy��$�<�|I��荼���|	8]���H�}�^'�5q�	�p`��wet�V=$_���|O�n���.�z�b9#��G,k�E��N*�㍱@�9�������S��:�Z6V��:ʻ2�M;�JԽO���m���]e�~ ��]�̈���|=����t�ԆA|V�aD(A��I�2�D��ߤ\l7Q{W=mש��x�* ���T+y;�����Q2��B�E1��Bl���E�d��^
\����n�8�qci��~���QeEzE�����I�w�(�O����rC�o�WROa��= ��y"��9���8b8BF��P���R;K�D�=���SHP���T����o�{RbFl:�p.s� �[$��3S�TI7]�4O��:9w��鼚� �gu
��PRF�Đ��p���Rv���^/?�C�w�� �Sz^,G�+�H��Ā���}SW5�&!&W�>��AY�$˴v���'6��P?E�~�9��rP!ֵ��kf� ���r	Yh�XrVu+�bȮ�{QعX��ŕ��eɎ��!��X��Lm:�� 	��~��mv�����h��VG1<��)v8��:���P��ncA��\s����MTa����hݓ:�c��Ŕ�f���ج�.�Δ8uD
pjܯ�j+�љ�ouÇ�<�mڻ7+��H�.�v�����ntu������<�rv��b����5�<�h�-=q�ns��ֹW���um�l�Ar\�����B>ێ��.=u�Xn,��sۤ �.w����r^K�n����ƫ"<u��	�n܎�|������'1Hc��vfW�{���� ���'�ʮ&�^��;o�h�-�8Si��F!�N��ڷ �K���fn.������$���2	��f��UKs��J�����Q�N�WU	[��H�.�Q�;n���N��P�	#+q�@��$\l���Ns�1�_D�N�|O����� �I��~�v��Dt�b�(to�띪�c���P�Fe�����dO���sz��e�����#�]vH��7�@�2̜�$�!I0�L(��~.\7�rVy��v�\���]���'6C����M~����rµ	�	�\̛��>'�mfL�A;�}J�G��J��r��׋v�-�@
�d��Y`�(Bn�n��o+N\�mzm-��n�~zx!0���Pv:}��(/+F�7��㉤{�z�;*�l�X�j��'��}�Vt���n�;���	�3�>��$����4H0���Σs9��p�e�Ci9��w I��;��}S�Wj���lIW���}T	Q���A��P��=��r��Px8��Io�I�����@9�r��>���]���)�y"�!��0(9y���ܑ��nM�=�A��rH��}T>'���TnI���W�����_;}܏<tlԼ7��B�'F�CK�z�[OK�Q��uv�������������f�]O�ݾ$�yB�$���R��{�{LH&��US�!�	�&
L:�����^T�S�N��u� �=� *w��D=<"T�]y�:P���#�Ua��-��ݗ�7{�h��bC<p�tC�C�۸�Q-C���s���:-ج0o����
%\����������rLs�V�G����ۊ�M���ɯ�����ۯ��w�TI#>�����'�Y*��N���]ΩR��C�;��B� ����^$�E�ꑮ��Ϻ��&.�ꉈ�Aci�ᖔ8BF�\� P���z��|��<���\�(�}ݵ@�@"�v}&͹���B֠�@~�:��6�nP<FKs-��o=s�+�Z��-�]S�($���o7�$��$�����	�{� 
o{7��@��o�~���{ݵ@���E(I#2�nA'fI�nNo �M��X(�H��ڠ	�E���A={���s�}5�j�D���a����I�<����ۜ�$&�gI;b�i#��j� �.�g�A�h`�(PCm�ܫ����ךZŸ�����Q?B=���s�E���ËXo�6�e]�~�R`������9|���kQ��Z)݌�;���2�V8����8N���eh7�x�,l�\�&s��2�Nm�uD}YlO���*P��qI������5��@|�:ĀH�}�@]��r��:bm�qZ�ٻk�c��;�h���;�q8&\�FϪӻG�@>c���A2�P�u]TH$Tk�hP��=__��IJ.�5���  #��@����J	�$��j{k�H���5*毫�g��뜂A=o��ă8�����Oe�}��q��	$a�XmψY="I'��M�X��DVP��]3����A$u�ʯ���a�N^	��G{|����-m�뒫[�@>$f��v�LΫx�O7�!�i2H���#S�0T(PCm'�{/(
>$�Κ3u]��ٕ#����s�A"��S�Qۜ�
7(���q걄�d�C���Χ��To+������2Ew.�v��`�n��N�v��RclY�����m �	x�=a��b7Dj=�Ȼ�ٰn��{@�jl�TB��tIҵ�)�&��yl����{2�$�p]�n���F���y�z�E�N�4	_%�{8J���vG��.�ݼXc/`"_[�4*�a�r��a��꘷j(����3�����P�a�g�we�]Fj���k8�[��V<�ʴ![�I��H���j9|�8�w�d�Y�;F���
%��h��ٔ㧲d�U��gt�/uΉ3(m�ԟr�x��kLFF�fj���ʥkVЃ1�C����׉���e����p�&��/BڕG
����%�F���>}�u$��Un��S����de 1٣�݌LV�12���C ��sZr`���׀�K�i)�Vϗ'�}����=r��]�e�w^�7S�Ne�B3z"���|���S ���}Qt��t���7g��̻x�wt����![�-�M��۱zo��|#sb����w��场V�B��K����������[�8�őf��WK��f�����xY�U�5���+�G;tGy7��O�
��d��i��>�`n���3j+�:�2v�K@�ycit���[S6Чe�/ >Rѝ�6��� f��Đ��F#a�q�8�g5���8�#ӟ<��+o�2��-�[Z��=QBv�
P��9gy+�^��q�:��.�J��V7���ze���boU����wR��J��hЭ��)Jը��Um���j��eZڭQ�҅�-��KV�Q���#J�֥Q-�(�DkB�l���e�ҌV���6�Z�%E��2�XR���"�i%UB��Q�IUQB�D����PYm���ffb����V�)kb�"�J[b5�Ķŋ�D�m��m,�F6�
����F��JU��---
�F�W+\cJ�6U�����mR�R�۫.���Z%+*����V�QU�YPZ�R��1!Zª*6�)e���e�֔Z4��4��Z��X6�DZ�UƬb�ƍ*VյQV��(��+QEYY\̊䭵q̦���EV6�m� ���h�kBҫJ-�fU(�m�6أJTmR���(�V��ee�6����X�(�h�d`��VփV����iZ%A�h�EF��m�֕P��b%��Z66���Z�[K[YieŴ�.�MR����
،DjUmm[h([e{�k���Y�:pW�l��1�x9����⮞^.w6;�H{p��*m�7&�4ⵎ�s�8@�^.�{4���덷;��4Q�	��ڝ�6�Rl��un�']\;�g��1�cm�,����n�Mǳ��6ݟN�W�wa<���r�v꺔9�sՋ��v�F���=X�@ʋ�N%|�nC��ŝU�n�h�z�븺K�p�5�+��M֞�k�����n�
�U7+���2"�˴���7$�qx�F���\��i�q��\���8w�W��W>�����fϭ���1�b�:[Zw=D9Pb��gګ��q���H�x8��c�c��	ݗ��1���D�c䭥C��^v'��fx�ͬqBu�az�����:뜺�:�;�ĜgvÎ������c�)ǫ-���>o��}G�>��8@����P.˦��]�rC۳`�0���`Svx�n�b�v���^d�.�;SX� �9U��tgF6b�#L����m��i1��C���F�͛;�n�
�70㳍��fpc��A��н�y�۶������@ئn�zN���r�U�p��k'�g��V�WCv-m����ή�`'��x�3��O1X�<�q{s�Q8�ȠrX��J�{�k�N[En��gq�ti4dw͞Q�l��[%�aó�e��kE>��3�亽`G�8�n�I��뾮�ی}cR���9m5��tv��[�Z�݂qܧ�JSt���a#���z#�c%�܍�-u�z�u=q�Ƕڻku�K̳��mg�
�mɰ%+z�n�V�γs��m!�M�v�p��=>�<�4��\��%5c�;%�K�s����\�<����
�ZE��#����O��(kq��,��v.�T�i|޴]̪5*��->����B�݁�m;�m�6��%�gb����"�l�.(5�y�����c�<�'8炻g���w<sF��ֶ�Kmt�U吪���ﮎ��Η�f�<�2��h燥��Xl�n�7m!d=gQ�ۘG��GYz�>I!eˤ̵�f4M�\.�,�nW�p��[(v<�O���ؖ)m�v�.]=����J[++tq���+˺���^t�gb�1�s[�d9�+j���9��D�k0���c�-��/I`�nՋ����>������Y軩���%=s1X���7W�xR�u�sQ=,l��0ro]v�m=^�y�;1���xE[�������7�5=pmn��@��.A4=��7�&8�n�n��u��uz���ճ�]k��n��s���|����d��p�9�컑$oe
 �O�vyV��л��r_ۙ�hP�$�jF5�(4�P�	��m�x�Yq�o�]�bI$�>��o�:����q&r]���$���R�C0�0*�f����|o7:h+���5�EU���$���U�@7��4Vr��0�6��'���Jڠ����'��UA#ss�| �|���Pt��{�R[���%&�)@tv_H�Hm^L�S�۷��Y��� 
}��U >i��{��{����>�?��m��l�r3�.x4n��箵rD�[�8��#+Z�W*�;7��Ϙ��b�H?Nm\�/og�A]^�_8���p�n�(Q;��Tc��L�Ba��9��[�6��y��Zw�dʹ�ڽ^��V������0���cu4ng������;��C�� h����41e�^1���Fvw�=��Mx��M������v�A�Y~'�i�� �iC�$l�]W����e�	��ۋ�\v�8ǶI=��T	�5{!�ӰAJ	�$������T�Dl��>.�zkĂI��'Ē7_eLY�x��M���O�w��@�bڈIl�r
/:Y��177|�N��P�S�D��� H�>ʣpz隮Q��m�Xk���SR���|����m�0U���b�n�s�1�� |�2�G�;��)�Rl��\��U��9z ��V���^�{{y >}\���DG�,�`�e�
 �{����5Q��ٻ�� �S��;=�|Iސ��k�vp�����&7W�S~��$�D� 'K�7j�n��b��K֥/Kn�R:����׽u������1_�N���m=�T�K(������D`���m=���N�v�*3g�\����<<_Vw��H:k�0I�ϧ�^u-e�A�Z�Н��U,_r.$��J���	���U|���l�ΎSh �Sk���	�K0�0*�T��oszh�Bz��:s��@�_z�j�^� 9;ھG�-V��At�@��(d&�H	���ǆ��]ͻ]k�N5��Gs���׬�����߿;�7�p������9�E�wMY�1{�<k2X>$]��Q36�L"�d��:�����񛈝9���A"�o��O{P#F�2�Grx!�K��xn�-�$���^���@��uc��ٌ'��E�oM}��[1	��u^<gr��x#&��L�d�o��W�ٽB�ӷ�l7
KUӽd��m(,.��+��V�[��t��%��]��3��To{ë(�n�\"��J�Y�G�����f���j��P9}�xx`��;wU�C�W2�!���'�;��xH8v�|��8^�T(l�ori ��$ 8s��c+zR^��·���ߟB��O�LX�9&�뎸[�-�dx殮��P^7.!�&��!��{���Y�������H �{U�Wr�!�z!�&m�(Gt�� �v��QZr��*�M���g�P��Gl�MW��E�wM|Iӷ��̲/ǍȊ���e�F8L"�0IPPZ��x��I\���KE�ͷ��	'י�T	�'��O�Ih`�Q�������m����:�� /y��@1˭�
���W2��M�EϤ��$s���C�Ba�3��ͬ ��J7�d�l4o��D�*��T	 �=yNV�M�9���x9��O��z�4�7^�Tk
�R�����75̻��Z��U�=�n+V��eP�Ķ:��ۍ�*����������s�b:�)r��5�[MfL���oV���/ k[�cۧ-^�s����[s]���K�,-��1�<�]G�����n�f$oKN{ݮSh]Y��k�kʬ	[��#m��>S�q�l�u8g�r{9l������S�=¬�x9Yv�0���ɤm��ٵ�;q������8�89��������Bɸ�_t6�W=rq����\4.M�Bv1ٻ���/]G=�D���Fwj��F��CI� �
b2�q\�pD6��#�9�eP$�=y	'�]}Bjf,��^y=�Dx��.V�
P	fQ��������0�fl�|x��I �u��$�����O<��a�-���P�&���u�Q�l^�C�T��v��3�A7[[Tw���C�
���n��ūzW�d�7> X�ۂ��/5�D�/7z�=
���8����i+q��pă�{�(�|w;zh胒E�Z�7�H�ց��^H��=�H*8�*�KI�z���#	.��R.�t��!jB�W>��9��ϡ��rV�]����f���?��ÀBa�3~:z�$e�P�<H$^n�Q̜�ō73��&d"��K�u�(81�k!��q��}�B��ދ郑��v�D_<�e�^L_�^����u�u{u�sD\�n�
�0uNw�{c���tmi�w��z���w<�1,�̗�J�����x 9��2I>�.��$/>ߪ� �hՙW��0��f�l�$� �`2`U���$^����R2��w��7�va~�\�(�k� ��� Ì[JI6C
����V�^��A�w�D���F�z�u���8�ۚ$L��8L#
b�	��z��9��pyd�fj��#goj��>���I�=��IEi�һ#�`0RK�L9��v��C�����l��Y�(v}x�Rx������`�m�~�p;��B�۽4$��^��ͩ~m*�(	�w��L���ppS�S��㵒FUާ����H=��B��K��f�P��5�ww7���z.m��:�A��X(���}��ҧSgۓp[{��xs40��DF�,L{7�jr��xno+�����^'v�6��p�0����Y[�G����3.����uP$�!�d�d� �L
�SY��
!,}ot]S�DH��"@$)��+���Q�@�	���/O1M(E$��s��ݟ2'^U69��B�OtQ*��Q>$99>`�|*v���S"��B�܂	Tb)��Oŷ��o��Xϝ�"�z&�����H�ϟ���3�]�!i�� 	�s���~Tu��F�z���'NHdZ�G��Ӈ��'�UHP���'`�0D��  3헢��?/��}ЯY��2؇"�4̵Wpʊ�<������� ��!�7qJ�GM���|Μ� �����&���YpCl�P�M �������;[ˮ���4=o��c���,#��\vӿA��d�������u�*j���f+�[������7Z~�`��Oqt�@��z�^+>��T�/9��H��C>v��{�g�<!�t��c���B.��W�j�h?�?~��6�~B%���'t��L���۸��#c{��]7UW]na���J�1��Z�%��R:�\�9��끍��{΢,%�� �hǮ�Y��	����� O��M�]��Z����χ���C���u7H���n��\Z-��d��⃼�T�de��>ꭥ=]T���h 67�������zo��Ҡ�뤽�r��m���^]��wiy$�{�� �#�#}�}Rguw�|\�m�6:w�jV�]"��*4�m�Ω�Qv�u�n��]os�a�Da��bWw���Y�ݲ�`�-�ݪ&�3v.m�
Q�ƫ�� ]�V	��{o�޻˻H >:7����+��i�/�/}T���
4˿��].�1�ƍ�%�F�㞝d֑�A��������0��jC�e���{�]GN��	]h�^������[��{{����*�l���4�^8�'g�v�Ӕ'�ֳ��;vh�;���oG@g/��N��*vٶ�7e��os�r=�J�݌���t�>4���Ca3�ȶ3�c��(��\t�v�<�u�M{u���.��(���Mssˆ�f��Se�Gjⱔ���C�[�'��]/G��΍�mj�*-(��e޷�V�n����L�X�y�t���u�y��N8n����4�r�ƶg�j����ۊ�)�Lц۲b3|�w���ӎ{k]1�0�t�.��� �#��� �Ww�Oਊ�Ӿ:WE�ݯ:���twsiPM�M��A3!��x���އ����g[Ĭ @i��_� +�� dԮn��߼׉5��ʰ/&{�F�F�n� n��n�|����;�؎@|dosj����E�:-��?'U-�ͳ��!���������.�0=�w���Hʐa��',�U�2�4�Ů�)�2M�[{m6 d�k��Y�~�X�m<��ݷ	$��sU"v�ZW7=}���f��
ɂ�"ˆ���,����tE�չ��q�T��\��uu��M�����1��6˅$�W+���H$2�j�H 2{���*ʧ���������m�URFC�
���4�ʦ�nŒK�>t�xL�B�]ѽ�h+�糒O�zs�����0�;�����ة��w��_S����nG���J�w�0}܀ja�7��{�Vw)Ƀ�	$�]��$�X��&�;�N�����^v��q�q0G�L�D�:ix�� >��n/�+�w�Q�|�"}[�� ��MX���UB�F	m�bS�
5W;Ι�k���L����U�d�kn� w��C�=�/Sp9<�$lY������8b�vvmش�A.ս0t�D�ꎪ�GK��H��{�wi��ި6F����0 �B���ix��u���<��u��+�F7W-�/agql'=/������
cȕ>򨅮�l .s��� ��~anМs�����|+�m���k�ۻ	(8�,�!��CqF�5�T���g��ۨ��l ��n��DF��ST@��Uܮ���������8(G�o�J���ۢI8w:zR%��m��I���wZ��Li"I�n�j��~�M�Y���a���N-P�be�ĝ_x�I�Y��p���R:E�$��ch���qer�w%
�[�h	���&oi�Թ��s(��D�ս���(\�Q��/�����n�vK�J����\�Wx�`�ɶ9mκ����5K�lMd=ls��fT/�Ѽ�*��Y��p�ە�ӖU�T�cz�_r��]�YT�'X��v��}|,���2�Gg��n�԰3:��Պ��F�k�\���M �r�0d�!@5Rfvc��8�i4dÃ`t2����[��+�~&��ov�^�\P��'�&j���7�u���� [m�[yq���=�w�"���/�g3cQ?����#;hk�d���u�P��5cZ;/*M��os�u�u�w:�Av�q#�`� ՗��=f���/��P�u��݂q�;R]�z*����͌�EFJ1�yA_r���Ef���o%�J�ګ��*�<d�o&dz���)Ui�u3t	w�LQ��1u�)�)�M���V�TC�Y�%c��dT�/V�T9��]c*wfww�<��]x5k�Vb.�h�mH��X;h,`�Lh�GI����/��졛�I��8l�eC[^���5tI�d;R
N�u�}w����q_={��wfۂ��u����3D�يfLxs7;�o: 9-�햺�xq͠[�f�Vhh;��F%���B���WBr�M���^V������tܬ6���X��c�'f���n�K���
ҭL�n��K�g���/s{��g5�F�"�,DeT�j�m�
4h�+TQg�G)J�-�5�V�Ҵ��mKiZ[Km�UP��KB�ZRT�h5���(�`(�����Qm��[J��XQ��-*T�pmDJ6�Z�lU��Z���kh�b"�V�iU�J�[[(�ekX*[bV�
0GU��F-Kih���
U��A�meJ����
ҕ*6!ch4V�D��ж�Z�6���R�[ic"��h�*Z5�+-�V�Z麲��h�R�3\e(4�
8�D2�J����
�U��V*ѕEQX�m�T�b#U̸
cQ�"*���J[K+h��Ub&Z�UiJ��ZZ-��ZYQGVc�"�%ʵ�0PF#1��[JE2�����(�(��R�֭j�m�հr�E����*Q�R�km��
��ģ(�-�mX�1R�%�\e�TKh�-��R�R�ԭQ"���[EB�Q-�R�Q`�Xk4�+����҅)m����jG-�̰P�U���Z5:�34
�E��a��kE�������ͬ��� ��>���I�w�J0��0l����HT�Au�����k{^� fk�`�R�DB��%���s�W�A�n�ߒC��b���4.�
F�o���&��IE/��{����W{�w ���� B��UK��o��0�䴁ZH)Yq��qk�x:7LvYy�0/CG�k��R�q���;7�������M��\1}役�v�Iq��f�I �+�������*��NFh�ݷd�Ia��)lZ���pSP*���i��S
`�g{�͌��}`���s�B���L���mr�⫽���ha�mCi�n(��窼%�����>  ��}�;�Ns��������c�m0Q�=��/}O��EMg6�A�ħ@�s�� F<�LI�λ��|fۆ�W!�:���Dn#цvmB�<E�2N[�Cx��G�f΢��N�.0kԶ�:���xڑWl�n�xxxL����\Ԃ^�鸘#�&TLJ0N�[b@|��'L�N�/srЬ`m�tX��H�Y�� @evuݠp�{�|���x.���+��2�o�i�燮���Z���n��A.��ɸ��[h��(79U�@D.y�6  ����ꨉ������nb\�`]��L�^�(����7{6�Dr��GMW*�1�:` ���� ���0Q���]�2�]�б��7I^튒?I{'�"n�0�(�,�Ƹ��N$F����	!���d�a�rn�!��7h./�/m�*��u�в#�R���Y[�w~Iy#�w�up݃���eL�[�$�B��U%����pU5�w�B 27z��y���]�^ۮ �3s�4��n�����<�q�^�L�"�g5&n9W��w��i9��v�Ε��&aǏ�l?\���ɖsjӉT��MYZ�ǳQoY��.���D鹶v]�p�ʝ��,����ђ�Kg)�R�<b�F�xT����.�v�d�u�s�w'��E��Ӳ.gqغ�⸷M;(7^������8X-Խ��X��(��nQ.u�i��s�d�܆�nʙ�ey6�dK<s;�͢Ν�n����:I{u�k��R�%�t3��Ş��G�.��t:���b-���1�v�63�C��ܯa ����X�!���-=��q���q�^v4@Ztc�ݺW.2�g��ʈ@��{x�����'����m� ���]�`� Y��~={�}&ɾIh�l�H:��`�9�TO����W6���nю5F����b@|Y��E��i�ܐ �M�w��Z661Z����-X��Np�%6��ݻV  �7��s�8Ǥ��<����M�g7n�$���b�E�n�$j�!�yzc;z3�S�ն�+""�o?0
�c�!���Aѣ�)s�wi/@qڛ�����>p��smH ,}�7+�W�{��W{Ve =��wa#x�nH>k�$M����  (vv��6o�9v(uE�ٛf�k�n��=�mu�z=By=�m��v��w���X"<a��e�mu�Ig-�@ "�c���!���;�m}=ٗv�#��mHz�&�`� ��LJ0K}۠�<��˱�1[�XO��mk��w8A�1���:�^�oe>�W�w�]��E��seq�{2D%�>�W�DHn@]�ZJ��������gu{�� ���??�@|+}��@�V�s
j��I
�c!�" �����	$�����I(&,owN��L���N��[�A��^B벤��CC	8a�8cGOH�1ϕ/H ��D�4����OĚz- 7�ͫ�{iz����'�3��SK��[0��6I-�PHn�W��l�&�r��Y�OZ$��~j�I?��h�������G){�D�[���c�TM�d�c�#�dz\��n�YO]���;h��<�`�
b,ow(p"!�E��v��!�D,}���]�݅+X�^+�����M$�]�&�؋G�8A2h����� �3�������x ���$����tO�x�4����v���kc��Hy���!�B�n�b@�n�V#��ކ,ά=Y0-�ű%͕{G2�ỳL<���g;��WK:w�d�8���I!��tpJU�ີy5�ۛ����Q�_�_�\~  @�{*�H�����m��%Yrrbp�p���f�'N8�;�{7R$Cު�䗒C�{nɰAgtuq�%�f�������Bvj���CC	6ˆp��]��w`�;��DFzW-�녞������� �����#;���9�G�#s���T�$Ȏ_�G�q �� �a���q)kmk5<�:����s���f���Y����DL��o^6���wd@Y�<��έ����V�o�@������w(pF"�Q<�t��Hn��[m� ���� ����s"n�i�np]E]z��o`�Dx�0�!�˒�$�z���� �:;��kA-��3����
�ٸRA�K4�����������NbK�뻷v�gw���
�1��没�f�
���1��@�vE�l�5=;��������J��wv�1;n�n�vw?u����;i[��ۛ�Yr�	{1�ߤ�aLFLgFŚ�����'�J�϶��N������ \���}T!H��m�ݹ��UU,ԃ�����A��!����̪�Z�u�(=`�(�T� Q��{;��燓�[��y��u㱛�ݶ�z�pa&�p�.�[{�֐Iy.� $�ux�G[b�y�׷:�	$����	t�1�G� ��$73`l��F��F��k���Dv��*	����I$���T,�=}`Û�	/@��P�aP�F���$�	����	�.����yz���ߒ+�$.o*M [=�X"<a�.
��;�����u�$�=�f�$��Z 	��7}��	�*Ėω�٪�;��C�<�aD�O�O+���|�{^���<���R����܏PD�~5�rH��=����.�T�;�w۵�13�)�7�)*2�i
K���һ(�K��h#����=�vhJ-oXb��e���&	�d
u�qF�}�<��(���˛��1���v��Jx���Kѵvc����z�ֻ2t�ݶg6�:�S&�Fa��n�C��N܃���t�G9�'��R�&�����ɞ�k�����C�bM����u�������Z�d�nյaZ�Z:����;���V�E�����p3����q;�����v���:����y�c\�A�[۫v��Q��]�����ӷ7a�l^�%�y��Ϛ;O;�����yƉ{Gg���$8%�w��؂����^S�h�[o*���{ww7yU�>�țۖ� ��[L�5�PL�O�"'Ҝoncߕ��b�٩���u�2i��{T�H/��� EFVϕG���[�u� :-W5��d(��w>H�I�d�rA� t�=A��{rp$�C]�W����ۻ	(;�&XF�`P_/,Q�*�p�_R��MIM����wh ���\��Gϖo{Y&<��]U$g�$@&(�4iU=ۻ"�goM4��O'�]n� S�t�@}�]�w� #;z[F�Q#�AN�N;1�( �M�ٲ��);�ۛ��ǋ��U]=��Ź�Ǟ�ߛ����yRf"%mw����4��w`�@,��p�=��������S5Ͳ ����Y+b
�� \��|� I�JFY`�Ӽ;�-Z�b�˳v��NvÃ����gEZ �D�2|vD,V��ŏ#�[�A4-�L�[XȢiv��W�#�;����w�n��>#?7���d�^����u���?�e�R�����b�-�ݺ7���s^I$I�j�Z̯d�
�[�ڿ�\�m݀�3;�ג[�s�z$Ê�����z"��K/�m�[q` ;7��@���2l�tI$�	)��5��3(��*���ܶ�@��7�>���bF�w�I���m��?O�{�H��B�eU.f�1��ei��"m�NO4q�gl�k!�q��z�oS8=���(R��㋅��ׄ
��a�QZ�h?�$ɽ4�� ���O���Ϳq��ǘ�m�I������puwg0��9�ai��E��Sz� @.��p��s��!�>������^�"�5��U�clAP[��ԕ�I'C^ez� %V�c��9��Ҏ��KE,ɏ[�x�*������6��v�nz��!�;���sd;�{��=[�yZ��觕уc���3����%��?����@�W=���{*	�ϢJm��m7�z�]�  �ni���"�1�H�+�[&����$iX�6���sIb�b:pc���	W���4L��M�7yx�κ]��~���p��\�6� *����#���Uz$Lv�|���Yp����� ���Ռ�V�[O���^K�ƭ>�Z��lz����ߟ��Z�(��TG��߀ Y;�6 *���YUm�W{���!l�Sb���4H�Cd���J�;.Ť�XW2�|�=U��E�c� e_svv�w���R�"�=�`��P[�{s�q��{�Շ� ��|B�n�@|�s*�e_uݠs��2/�@�M��E���8t$�A�eS@ ھ�����0�y���TmRb�F��5fu9�VfV���VZ�nc�|F�"���4�����U�2:
���Ի����'M��B��o�Y}*'҃��Jlݼ� ���׏b���#���t�
*_:������#3���w.P{��_�y�߲�;�fX�L�Ze���J�)��^ң��f�e�Dst/��������
=#���U��V g������S���z+Ѝ����W���1ܡ6�D�4JTOr���I)xwkƼFJ�ު� ensv��s��]r��ۓ=bn�3ԗ�3� �L�	NC�ܻV �;����J-�u�?�u��v� 3�Ґ��-��DC����>�6��Yp�wR� �OV�a�D��~k� B�e.'!��Iع$�N��eAn.U^P��A��Hk̯Uo(m�;y��&Ow$�$��� ��E�~j���,�1儼��J^��ؗ[%��(pC���I�J5�gm\��3$��ѹU�.`F6��SE�>s�4Q�Рѩv��5&%�Tl�q�'eh�i����L�Qf���vZu xr��y]$ᚆ��c{�Uo}�B/o��o5����������`��s�	Ӳ��s9��1�dH��X��N��8oxN��&#����)��v��)�2���}�qN���
SDǽ�C߯omJ\V�]���~c�_dɷș�R��	�׳H���F�rwPT�Yչ�� uq�2I�U��EIuj��gV!�ḟd�Ʈ��H1F�N�&S s�<:p�ɗz�3B��n�.&�Al�=n��3�{��=�l��D�'F#��`���\Z��k��gu(n���[h��2������-���*��e�Pb��O��^��n_f�ȎM�jw-��`[O���qS�&��QcU���o�v�V�!���װ^��}�r%=��ݞ͐Pu���u��ꡉF�aD����;�ƛz'R�v�R��WV�1o]|�F{�Xws��w�]#2����Bu=[PΧ�J��J��K�SU(s+���{Z����L�nd�}a���_<7�>�ox�wjK�=��wR9��F*�[�+y�z݈��lvE�&�}�;���v6!j�U,f�cT0�h9�RAZ�R[�ӡ׳��7L*i��"]��8����t�`����[@U��:���(�R�����Щe-U�iDƙB�"i��+cYU*5�b�մ���Db���b�jQ�Ա��0��N&-�����%h",�b��b
��[j�X,U�֢h���ҩEj("ZTZ����%�b�Z�[R�i�Z2�[��bY��"�F�T��T���mm�1�t��64m�km\��Q[T��E*Tb%�q
"���[*RŪ"���m\�2��V��Q�)r����cR�Fыn0�.2�*�5�����CBU�B�Y+P]8�R���*2�VQW��fX�R�*%*�T���B�J��ZV,�6�]9���ڰ����� �!JҌb�(�U-(VTb*�$�4m.Z(�e)m�Tl(�U�1T`�V�Qݎ��7`v��cH�;ݵ)l���V�ҵiV���ԬX,�ږajƋ
�l�m���J��2�QF�Z*���U�1G�+R��L�f2��+*Rڋic�`�DA����Ϛ�%\�b�9Dztd���n�˴���Z�q�C�D�G-]q>�r��v�� �x����9ܾ�px��ۮ]�n�Mi����!��m����]� O6ђ�r
C<LmlOe�5��Y5
5�)=nc�����n r^��5�;�lb^�Ul�͌ݔy�u�㷵^ܦSN��:ۮ�����шK�ގn�u��n���j�#������k�0a�nێ��A���~��� ��g��/@9ܜg��������䵤nmGs��#�A�&a�����vOi���l݌����[���	I����6�#<cb���Six�ǶKu��ՂwC��c�1�M�a�%��g��n��n�=�W����8���X��
���gH�{�t`��ۊyͻF8$;z5F{7��۞��9g�_[}v}��[�\\��	�㇎n2ୗ�q��ɓl����8�pg �dMۄ,a�����c��b#2�O%۠(�i�ތ&�V�F��}}^�R����pi��ۮ����I�nOn:�R�sn��[���dA$����;��/��۱�4qq�r<����}gt}Fw�U�ru����\��Ǳ�g:���	�g]Z���}Yq���N��R���p%��d'l��!mk�N჎�wh�v�Â}m�r�`N	:�i��ݟ�3�;͓�'�ݰ������9��]��c���y���ʜ��ض�>�z�rƹݺ�m	w%��6��15[��{��nr#�*�5�B1����W;q2hNZv��!l����W��Qg���J�y��M���������G���G='����W���]�m�y��;<7[�=i�.�lo=x�u��h씾%�E��lѽ��{v���wk����Y|MWP=n��v�w��a��1#]�ڌ<���n�sg*�"��v�y�:�iL�v���Bs�eM�uǶ�q�ګy�u��.�._	��x��&�y���OWT���ζl���݁���=���spt���nΗR]Gm���v�������0L�^t��w��n��ܷp��-�łp�7�.�#q�mN�M�Ml��[�cl=�����eo6sٱ�v�u�v�-��[��W���n�cMx^#uۣ���G��cu�<��ٷPR�Z=��2�n�]9ܻkr<n�q��ݧ)K�Ի�y�n;d͕鍀ֶ8v�x�U ц۬s��kv�0&)���kK�L�\'\E<,�R:��Vwu�\�.�v�v��~~�?���p$s��nۈ�����H ����L����nOTaI{q��E�n��>�Yk��(Aaڪ!�y^�'�D��*J�V�� �=����
��DC�y�9&F�Q�݉!c�B��&=�"�wU�H �d�4�@Z��fl����u���ù���+�ɪH��@�-�	�4�z��-���M��4�]z9���,��o�9~v�9H2G��V��"�"�����.�����ʩ#� v��?�f�Q��{�{��:�Dk�s~h�B��m�V��^./�ߨ�۵Ġ��	�{����(��:ݱ�&ӹ�q�Bm���]Z ��G���Z����8�P�ePh���T��]�wHg�k��\�e�jH^CeU#v�I`�a(MDCAm�Ԓa]�&b��`��l	�Z����]���XU$nq�i�꒥m��h"Ҧ�f�\�g�o��wL�ų����̻���
��w�|gr�����rK�I6�]���l��Nۻ>����P�|��x�b�m?�`�A��\.ճ]K�e��Ne6A�Y��$�b H1T�[�YJ���5Q� Y7uLݵO�>"�v�<��L��A���R@��Y%��d�b��ݜ�I ��GM4�{E�=-�7�4I�rZ���rL .����Ӟ��N��yW*&Q��]���x�l-��n�v�ឃ����i9pr��mz�B�`��=��	D&	���
y�*����� ]��"7k����B�{\�-����¦E0z$�O����O{��|�Ӯ���R̥T����>������mx��8�Tf�_c��HDUoz�)^��p�FP�� ޻m������ _.���f|UE+[���vDܭ6�;����삟\dHDo�Z���8^���
��WNť��Ӕr�*�Pp��B%B�U��r���nMF7�N��T�Dv�6����	����\B(C�T����d�\���αM�
��`|��z�*���ʛ����	@yb�1T�udU#I$/gcm�ٸ�/d�{�M6�� A^\uP�W�A�ʡJ���<��~�{tŝ٫a���/]%�e�LA[x����v��!� ��ob�,��"��j��a�o}�ׁ z�0�;�u�ˊ�;�F��<���٨B�CD8Q҈�i��m�}]�lm�͂�w-�wS��D�u����d���N5�u��6�*MU���� [9�6F��ͭ������ ����4��c�e�{*'ҁG��)�w]������h�"*7.�� t�:�`-���%䐚p/GL�hs�u�xu2�������ǖ���y������]*7�]]<�����ʆqu���(A���#�������.��p!h�RCs2���3��=����΃#�Iݎb"!_�V&A�	vv��,�Ug�9o���\����=�����FSnh �ٞ�s�֎6��� ����������=����?��|�T Yu�6 �>��m���������(��s�&���0фY�U� ��r���v.ζ���c��]eS�ݝ���+�v6�[7���©�(�#���˝�`;�)� |��i�|�:e�̘$�4�xR$��ʪ�J�qSi��2�~�6z:���c5r����� ]�I� 37`|����ܿL��t���XI �v�RJ�V�Pࠠ4Xo�z�$�����G��:�˴���n� �7[` �����P[W���.�oS�ζb�ו#kr��w7�:n^(�����A��b�����ب`�Z��|]m"���Φ�KC2����f��Et\A{��
5z��0vD֪D��S����bx��Of�ʾz�&�yn�غ�!�-͵:��)d�����K\��jW�ʜ{p3����k����c�k��g�k[�Xu�p/#�[���;�\���Z�wZ3�pV̲�O����4��l��[��pW;��T��z��3��
�3��nX�a*�� �s���<�n���O�u�ö	�<�������_Qpr�H������[d�#��g�ɧ��su��$��툎�a��8�Co��R��3�� N�r�7	���?O�
���� 7u�ޘ�ZL
Q�I
�t<m�DD֙_��]U� ��|xy�*� ����½޽�sţb�;��#Ā�!zS�S�m0���j��{-f_��qo)�DE�n��I���R�%l��Da5���F������ %�S`�}f^�` w|��W�L��oy��L�!���*����^Hm��J���Ct��Ğ�4�D���*� ��f{z�_тvɂ ������v^3�KƱ�\�ޫ��	�9��N�v���%�lVj�%��4J�XbN]T�"PKN��	K���������Tm;��ˣ;UTA$���3[.�Gpj��6oq�ؐ}�O���ܡ����"�+&�ܾ#@_��*��m��]��`8[\2]J�7{���y�b[����w$��&�qx{)�H=5�{�}S�ɀ Y��Z�w|� �3ӑoz�)(g`re0�H�T��[�`|.�� >�.r���ܳ�����| F�7�]�i���u��,�'H#�y\�V���|�q��Ҡ@ >���Q����;��D���Kɝ���9�6��#�T�� ��:����};w�Oas��]Դ� Ww�� ;s�a\�Q�dq��T���AF7�
D�����cwX������i�{+������^t�}���?�)�zbE>�8"��c��x�b��sl1�\��j����m� A
���{(�D�#�%Jm��a�_K�W%���S�H e�:` ;s�Q6���M��lkw��٤�OqٹW���d^]%�5ϢH�h�'�"I�V��gb뱾$2�Ee̻�w-�ؗjv��8隞�aȮ�3�"��B��=����O�F�E�eM��/���Vuފ&�d�纅)�� �k��H�D��Ϳ�=+OJ"&f C:+-������ooD+筰W٭�>�co�d_��x�]Y��n(!T�Sa�ނH�0
�ᢞsl##o��t���C��כ�>6��0�:��<�Zv��J�z�S��Z+�!A&�L����������ڡ������.�bx��������b�?J���ymr��� ٴ� co�_��Sy�E���!z�[L�y�U^I
�Ȧ�h(e������UH|��q�ԇ��6����*� g+����F�:� ��`-�(�)���0����j�������S��۬�@ۚ� "�o��l��!�0�Q
$v���4�[�P��>����`� ���,"!c��������`ٖޯ�Wu��7Sw���*�^�D{��Λ�O;g�J�U�[��MJΉ����#�Bꎣ�J�f�I��9B	��

G�Ym�|����S}2޺uQ��hc/[T@ ��I�����b�+!�b��(B�6�$҂Lx�!,�!Ob,�v����!�{J�z{<���?�FK[)�|u8� `���TI$����<�df���H���mP(�X�OҡDC�A��Ӵ*�Jv[�m�KQ5��Z�y�lD�r�H��x�
-����:������{����P�A�3I����$v^UR	�[N��Y޻Ɛ�/�T@ ��*� Z�pXa@,1Tu]n�,[�"*': _^UD4nss�=�[���|�����۠ʛ��P��L�8H���U �K3:j�m�lKw�dhm� B�ny >�[d���W8��c�3�b�S�&m^`�.�Q�b���3�P5�9bɻ2�v�DC��23�VoaDd(�:�CeƊ�J���gԱ�K��	e	]rk�$��z��n%�Z����P�����`7Ĳ�a�5��M�V]%ɣ+��t4l]�Ѯ�o	=���8��vܓ�s���)��n]�:ӗx�؍.��[E�b���{uf�Z�Ǩku�V0�<��κ2l�v#(u��-�j�t)h�:���w��\\}:�Glc/l����+��[<�QV��-��A�*J�g��n����Ž��hvk/mک�4v��PPc��P�`�ᒁ��=t�46�$ �Ͱb���ͷ��ݪ�RK�n^T�7nh�d�E��a�.���E�_Cۭ�� �<��I$�O$�����U�����L�	Hc���!DC�A��$+�j�y 7�i� _��]���zm���� ��x�dDf�6�W���(�G�%�Q����8����J��]�T���73�hE�g>ʿv';��D��B��m&��"}�Q*Sh�v���ӣ��B�񫭷�ގ�,�ꦀ@,�޻� F�����t6��	&�!	a[�
mg�cR�4���+��:�:�B��|�����B���'���4� nn�"�堇+S��6D�n�#c�[T@��w��Ҧ�i��IDC��Ym�A�oC�K��I1vi6p�c�s�������f���{�1B6k�S@�n�q�u/��E������v�����Ft�eH���[��L]��{R�D�y��v�@x� �eI�S:�軹�)�)�0X�AMv���B�̧@ ?.��[���oOF�w$�I��K�&�A)�`�f��밵��������^-���Q�9R� .:�׵vԮ����ۼ���nv��D�=1"�zc���r x�7�s]�v��U��m�� 8�K?Q$���{C����H �di�D��c��t�b����S�yW[#�d�c�s7	�]�����c���&PW-ɻ�6^F�{^��Aqו/��x�]�)�ܻ�%yv�ڠ�
8C�h�A-5�Ө�yV��Ӝ���D -�n�D0=yU(�=9�$R��w�D�lr�������$DFC�n��__#Ǉq�6*�"�E)�f����]��q���GVޱuP�&a^���t��;�T��J|�uҷ� �RA�L}gy^��p����/ s���E�v�9Wۦ3�%��,6�m^9\�r�p��е���x�H,���u�8]�p1t�46�ц�`�4ko3gRq@�n���t��-'n�t�SV�Y�y�=�;�9�ˤ��kj	օ\%�%��wJ��;NSxonn����L>��mk2�ح���g3��3Î��[k33N�w(m��5i>���Z�� ���R�eZ�T�����d���c:uCNӢ��e!�;���]u��D�x���6��(��̥΂���=�f��̚^p[K&�p��M���cѱ� �l�BT̩V�޹�Uf�s�#|�t��`�y��_:���d�p
V��g_|Fյ|�0֡�0g2!bF}2r ��3^�lh�D�w_]&�p�,n���Q���ЁB)L����9�:�{QA�؝r�P���9=z��R�b�<S̚�^;=*c���G�i�z8f��#te�wv�Tt.�����iB�v�����Ѵ:�T����p����}y������\
΋iд���o,�{�����vfGv���_/�8yf!�r��Y�8$D7����D�r��+h���>�k�[/4��w�6��N��b7�(����ج�ۋ��7.��Y����<����X�͡�yu�y�S��TvRͱ�w%Z����R7r���۳u9�m�ǳ��H@�EZR��2)�F&Q�jEX:������F[UTX6�[)��cX�X���JԔQ*V�T������Q�h��ӂ�h�X�մm)j����IPDVXe*��V��JZ6�Z؊���KKek�fJ6�ڋ-ZQj��D��("Ԫ�ʊ�(�Vګ,k[J��U��2�0tF%�J�-J�lKeJ�f`�b��ն�-�Jҵ*(�T���ckbk.B�F��R�Q��h�ˍ��R�$r���m*�Z�J�
3�i�����T-���e��Z
��pR�V��e)J#�b��K��Xѭl�-��-�ж�\jV��P�*�����
�fem�Pֵ�F+(�+QT�Z.Ze�TF��.Z��IQqӎa���\\
�\�䥡UQLj�k����-��JWu��j��E��[rAD�H�	l��U�"P��Y�MR�]�^���ʂ�0���4�o��;w�f��Օ錨��5���R  �1� y��wʜΠ���-F�jR��p_�(�b*�	Q{��R[���+�*6�z��J��Z��g?4 0) �?9�y�D�����Y�ޛ�����p�+۫q�W%����n:�fN��Ha�wh.`,[�A����ϋsnGMs���M��R �y��Q�+�&zhS�Ը����K� �&����P��CĞ%J<�T��m�A���p�p�ۯI$
�X����6�A-è���>��F�^)n�Gp}�ޒ'��tk�I��{��Ղݏ�g�߳��[S` >:ct@��{��$�LpP��SP�D�s���u���d{6q ���: -���O�NPG���mߎ�zqZ��mv>\M��;,;چ3�m_N�Y'i�uL�qE�1��Bs�rXͭf��E���jCĚ6'4���B$��ɀX�g���֒I-=�4%R��ϝT��o��>.���f�%g�U=��s��%��lu�6�F����mwj�)���B�������|�_6�N"~��zg�����[������$��r�u]�]Oz1F_��������v��v��B�ZT=͵DF�k��=}T�u�Ώ����@|tvkj�Z۝���+�C���>���'�R�(�)�{�y��F���� �:�u��wE��ڜA������[��fn=�D�x���Sh6/rv���W3���G wz��Xvk���\]���o�(�%M�
$��]Q(D��0C�'�K�H7�KAZ/���a&�y���T|:r� TXo��R��<ٖ 	�~V�������b��x#�2�Ni���v;�Z�ʗw8L4w���z��1�)JsG��#gk�����D���w�����ߏ붒6��8c�a/km�����E��N��l&#�\�9�i�h�-��n�p:0�Yq�Y�(录+u�sm�N���^{�ʬoZs!� v��3��wk�-���۵�|]��[]�]`��r�0m��mvEL������;��N�ƌ�V창�\�x�{3�F��#6Ӯ��6�՞�'�<����g�Z乳l�ýB��Fv�ƞ��ك]��Y�y�I뇃e�f����la5��SB��7��|eҵ�����j���d@�S }R��a�Oݠ�$�k{ww����n�I�e�?D(m84����"pMH�9���7�.�@?~��� ��/��6��}R�+�9�uդ�:�v!��P�e�+͢����ü��sȜ�k_��$FF涕 p�T���aa� �������O��גH*'z�� �w�b�沎���̯$��Lշf#b!�J�a���:��7��gGg���Q�G*�t=�- ��)�D +�qx፲;hwk'���D�B �0�o�:�6��V��]��&z�O4v���~�����>%z"��GC|�C� '���[�7��4�� :>
D��}Y�e��a*+�y�@ۓyU�!�����{�x���E�V\�`��*ȃ�����+���-U�ͬTv��vQ���7|ʨp�'�Gnﴟ�X��>�7�� 徕'N�s������~p��Q3A*/��W� ������+[��kپ�ٴ	�tJ��INw���yY���0fL������o��[��"}}�Q��t| >��@ ��z�w:�U�$ 8������zc���{�zT6���V  ���iQ��[��&�Q��/�$��wy�Q"I�%1&��x�ݿ�����>��x\�6��dFdeݭ���:�Q�JW��7A�������_�.Y��.��w�^T� =��v	A�f9|~����X�F�(.j�4�_wUt�0��.&�-5[U)$]'hX��n'��� �޻�	��!���W!�����!nPi�Z0Y(4h��'��?��7 
�U�&���`+���'����d=���f/9�e^��SDe����^�.��uhg��!�����η�aܼ��s����������ݯb�k'� ,�޻���ؔ�V�/�a�
*k�Q}��\DM�!�LE�޼�X ��w\�F���#5�#t�6iE�ۢ{}����Q3�E1�smP >��Ӭ����Wk�DE��̻�� ���舀��K`*��^�/� �*��d���7p^#������z��qA��:�{�w}|�����Q
"��\��o�i�ٯJ^H�c��Em�]N��������� ,;�Lױ�1B0�(�;W�T��T��Y�.�y����� ��mQ 9��^	��=yw�
��W��LA='�6��T $�� ^�̗[�s>��܈���n��Ai��f�.��e ��E�D�m�{�h�Sھ�=�d�'G9�H�X]*Z�fw]��y]��w�ԺWt^*�ɹ"�kn&���_��0�DΈ�	��I��K��epG�aХ��U�\k^�+��f�[Ɂ�� جm�@�}l��	��$��ܪ%%���G�ⶴ�p��̷1 ��6�$�;Ϳ������:�h;+�F���/׎8�0�Շ��Ʒc̎-v�t�WM��1#������q�]Vj�Â�8)�6�zR  Z�`�o7h:�ڣj{���g$�sfzQA%�6�*�I*�����,]�9X���h2b}]�-���]{B�쮠 �4���DGb�蝑�OK�77l����`LD1��b��rq#D�ӻɲ�����`{&:�ˊ�d� HZ����f�]����b%m��h��U�޵:�e���X��0>��޻� 2;uڣ�r$�%UD���;=4% !vPn0A��D��۽�q �S'���q80��9� ��]�	 dv�Zgu:��3/C�a3J�Դi���*��-���lrg,����//��F���y��f���:����X�^�]
�����w�$�p��-2Æ�{kR�[c����=��5�H{D:��;	���#N�3�=;���wj�Z���N������d�j�}g�4��I�m��:Ɍ<�1��<n4��s��
ݷp���:�ɑ홹�8�6�^�\�c������i#D{,&6����맞��o9B��x�U��{O����	�)]�[��ֻ�ޜ%��yWlh�iua��5��5�n:u1� �R{fu�gK�\y����>|����x�� q9���3�yڰ@ ���*�>��/{����R�'��_i��wo]�K.5ba�D����2{�pJA̋{�K$ȸ�֝ v�]� "tդ�����x���g�=$��@.b!&PQ�Yv-N�ܚ�Hӫa��C3��L7\�j@vv��E���ەR���1B%�X��\v������>#s� K�v�> {��TI$�`^��Z�u�J� ?vV�ߒLt�P�*m�\n��&�&薂�^r랼�'�NI�~$p �0/D�O\�Z��]���_��H��Ɨ�����ڰ��:����|b7�����|Pbe��RP�"µ˪�n�� A�۔� �}�XF��y�{�D+j=1��5�ݠ ����dd�l�bf���e�[�b�+M�I�w����~����v�#�܄�4�3:�zD`�%�k2TYpjn���&��n�;=Ws'Z��y���8��o���n㖀@"��7D��_��`��ۢ{-��ل�l���M;��"1�� k���O�����$�<=�V� azj�$�/��e�0�R�컫���}��3S�CI�@<WE� �w{��dS�H�(��Hkvb4'�H�b�%�o(T��n�s�d��s�����r�H�"ZA$�S��6�~�� ���ρ7���D��
]�i��Z#�fۛe��Ղ��xѴ�;��0�E�X����u�R�H2c������v�μp�j	&V����;""*Fh���R'�]���obVþ1�4%/$J��$�ok|�@]��`W5=A����N���K�2��:`�s�΀;���y*O�FM{r&qݙ�Rs�UU"Cc]��4eڦXn^x�]�k�t�Ŝ̴k]�E�^sn����[�[�e�x��AID9xkLݠd�.qĹd��KM^UJ(�w���H�wd�E�Zj
���F��)f�k��¼��5�����y�H�̻����:JĢIqx۠�a��I�*\��J� tf�:>�jb�g[c�C�r�@-�����F��ָͦO�Ry���7����8��kU;u#����HR����:F
����8��@����̪� �n�s���63���ɽ�""�b_6���>���{��#҄za��OY8=)y*(b=;1�6r�EI����	��!�C��N��ڋuK�����d��8H��P=�<�2 '����@}�12&nﻦ"!�n��:3��A�o�ˈ��31��@�+�nJ7����f;��0ͷ/��qo����)=���y�v�h��n�.L���f$v4n6�hf�x۸���x`;: e�ǂ=��J�n��+1�1����U���˻k�ۉ��*T�>�;�`D�x5-���ﯛ�I�In��m� �\[�������-uJ��?����K���x��8��Dm��k+�Ð��v9K���J�3�������Y	�����{wv"63n� 
�|�����=箞��v�� ��L�{܉��@�J%6�R�Z�����-sܛ����>�ܩ �.-�5DDd�[l�=�~J4�7	6P�i��2�C���@E�T�
�q��"Uun�	�27q�D	\;�tLN�33�	�M*���:�+]���e6�%��G^S� p��03w�ޙ���]��}:�m�y/O�A�����B 37���ew�����Z���s� \�D4���w$�-�OyI�S��D����A����ъQZ�p:܃�1�R�nM�f�Y"`9�0[��^1eܗ2�뽵ɹ�Q�nV\M�*q3��;9�yTyOwv+�0<��B�u"�{b�9S�e��T�c,Z���c5��q��!�;4���:��Jia��3,�y�,S6��.u�>�F�-;{��o6�ǚh;U}��FwM�
^hm�Bs0�`5*���&ۭ��w6�m����.�O_]�N�e�u�v^Ύ�U���P07u%�gWVҾ8���OثjE�tˤ�C�z�s��J����U�<�ٝ�Y��}�� �ӺI��YjpivWD�<v��n�vmJ�:��$�Om޲�t���ȵ��u��R�T��1	�/2j�7B�R�'mKb�7�ƨ\��!1�yB�P:w��	�� �t��^��%�����zܵ�^_,]�N;�ܗ��J���(�\r�R��� 	ݍ��G+fp��޴����Vn�mcN���}�UX�ն������n�y�Cw��	l��	њ���{C�;-+�3-�Yz(�[�y}��;�e�vs9 F���[�L=q��h䮷���*D��+D�y���4g72�n2��{�a����6��6�������0��9M֋"���5[^��r����	�Ύ�9b�����yǪoT.���A:�-������Dc\4���`�ё��t�'�-�ݧUY��W[˳���������u�F7!hf���s�3Ə��Y涝�ij��q۱y�5׸N]
.���Ǹ�xo��5����
�������=O��E��Ķ��q�mۊV֨�
��k�*�h�˙�Jb�ƭj�(�b���5un*�S2����b` �E�t�F9n�r,��\Ũ+�UMT�j�s�P��l����-�Q�iQb�-�eL����2�"+��������,Zآ�Z"�n��IKK4�U]4cZ�J�S2��K-�RٙE2������Yl���Qq��YKb� �[Q[V��5�1jX��Ŋ��օ���#K*:,�[F��knZZ��TG�J�KEE�DQJ�e�T[s[r��1�(�b��X)���h+�5L�Ԣ���)KU�[u��(j�Uf6TV�EU2�S��DHcV"ƶb���YM5i�1���5�Qf�J�\J(ZQ�E1*53,j�J�-l��8�ʸ�waM�8�0�fPĨ��lU�Ve������-�[nPŲ�X������~������N�Ak'@]rA��ʻb�o����S�����U�T8���J')�8�<y�b��k�ݳm�m�c�lh�c8$ԐK�F�g�WG\�#:�ukG�J��	ť���]�ţby�e�#�O ��v�Z�l���ٹ1�)5�[�^mSp��\�;g��v��b�M�����խ�e�kK����vn�m���n}vG\�:�硋�zf���n��^�=���!�Iv١��ʲ5����qn�m��q���ӽg��a�s���,��0Y��c�X�,�v��w=Y���6:���pv��o<gOdŶl�mf�9&6���̈́��ۃ���n�9�Ð��e��ۃ�.:�6��8[�գg��1��c��ܝt[��r��Ei7QmY�op7]�p7��H����۵�yF�r=�j����Y�ٺrtORv"�F��ON�k�pc��8��m�[m�k��qO6L�h��x͙^�`��Gv�v�{7ZC�7c�v3�:rQw�;�;ǚ�Ώ>ǣ�͆��^�A�n����Ɏ��r�����e��{ca�	�,�;s����]�A9maS�Q�M�v��]�<�*vW���۷Et�qd�[[��K�ɻ.��vD61+nĳуK� �q�H����]��l��q�7rrk���s�xMk۱��g����{�m7A�qsV؃{<v:x�q��c�-�tk̡nb����[�!͎�t�|Q��ۮ
Tæ��}Q��5�n���t�s�͛��:�pv�����t�b�g��՜����[��3bl>8Ju�8���s��7e&�ׇ���/�j��v{0�G���ܧgt��X�z�[�Um3cGX�t�n���%�*@����s���3���A��%m���%z�.����g���'U�ZF��i�{e�6�d;�^J���@����'g�n�ɮ��kL�އ�۶m��S�x��=�c����8.�ɹ�AМt9hg�]��nk��tu�����c�M�g�9k�p�r���1zm�+�u�Q���Nz����=�9�U��z���=siҸ�u��]�u��`Q��]Uy9�y�zۯ9�E�l����y�uҖ�k9n�k"��`��Nܨ��<nŪ1ۗ���Ot�f�E�y�v޹�ݧ�n�..o]Wk��sg�l=�+.쩬��m�{`��r�B�Z궇t�=8N��{ZU4/\���r]�WXw�6.�䧃s�l��&�І�ݣ����߿5rx�*H���/j��k�m� go]�R.p��tt��d��"��j���Dpe�

P���6�Ť�}jZ�qF75�X� @(�|�!��7��$�L����˙v���뛂L�.�x��x�%6�1�$ n��`����^��=ՙ9�����@Hff�݄��	0����iq��*c���Ms��}G WyͰwN�`:$��F�0���y�ƍ$U���I�z�l�TCp�*����~���c�i�o�-�'�*͊E;�L���7�� > ����Q��v�����L�����k�磁��i��y;1��"�%�Om��i4|�G��/xZѢ ��VO$�޴؀A�����۵,k��\�esk#�ԓ�@WI�m�k���P"<�a�
�Q	D�.�u��]���	��uо;7֪V�<#Ѽw;kB~�kL����X�ݑ��wd.�E��&q]�;{f,��]��1�\�|��7�� ��ݧD �t\��a:�K�h��aAJa�7�v�^K���4�	zzn1�B���q-�|�� ����������y��pMBb�	1U�m�����)�,�[�_D��w����`| �z-3X��` ��I��[�dˇ��n�x��Ny!��B�ACv{l=qcj7�7<�@2O���� Q�^�U"�vB}(s�ۿ�6E���w�<͘5��cS:S���N��5�	����h���1��ɶ�"�	-�e��ݤIlv�5@�(���B�D:(q�������o.��6;v��q�^JgҠ�AT�絤؃��vo��Ul�s��  ����>@$-}��@�n�>�}B؈��a$���Ɉ`��*;����cM� �H���]߂���޽B��=�c��V��c;�u��16"��6YyL�0pf�v���mAhhM�Z�w��1�^�BrUyS{��� ���P�����x*i��W�z����[�@|*���y�����u)LUv'�1�7;5�K�ݘ�	�pap���n�?�`�w7)­j.�j7����Z@ ��7� A�����5ً����[}�鰄kP� ��2T%�����i50-fw[�k6��4Wͬ������,��S3�Dz���o�T��4�$�6�qm�!k��,��X�䴃D�<kr�T��a��Cp�%1Ko{nŤ�w����V]r�A`�� ��w~H����/on�M�	O�Z,@�Pz �hN�N����v� e���8v+�ɜI$сtX$�=��K�����FOtȥ�/25!Gm�B ����� ���jcw:�r��)��%�����-U�s��Xc�k9V�HI���ԗ]>憦�sѻ]�[5q����5��s�'tlv!�q� ���n��썉=$�{���b�~'�wj����2e
QU����� ngsv��S�;�M]� � ^�1��DG�I@J�cr�ͭ=��h���g��4�E*�C7����_�!��S���6:�B@ ���jȈ��Xn]�Omy\�>H���� /��m���<�Đ)S3�Dy�������mm��˽�M�t �[��w �B�ݦ�FQWս�&g�-����)zf�l?��iTR��۱h�F��6�3||�_guݠ;u�{55)L�T�*� p�]�r�q�ԉ�꺿Z%��ݩ&����{*���l3ш������md���"}���؟su 1��y]���"w�ݰ{y�v ��[��|�������o�c�r�'(ӈ;�Q}z ��� ���qm3+6R�v���ie��m�����ch�6��c�&>�Hĉ�p@����<�J7<NԬ�v}�+u�λ>��l>�8#�j�Ti�-ؓ��d�׶�r��g�����Ǯ�n�����4W������z4�Ɖ�v�㎯�u���f��k]�}qKw��K!>�4m�8�[�s�v���+�>�Vv�ǘ��{�q�۲�]�3�٥���ω���E�u��]���l��h1\<��Ż"�j3�]��t�I��^`ܜh��3�<^l*[`^�X�vݳ�D�0o���2b!(��s���˨�>��O� 0}�Zí��{ ���9wv�	$7�*M�j#�jXl�$O�9�~�>�(N~�ǯ"^d�of:h"##�*b����?c�ճ.��� ���P�(0ۈ&(�Cm�`$yR��q��<t�s��Z��I��$�$�<��j�m�� ?!�Ҩ�;{�EQ�ٽ�U$�$u�DCH��9�aۻ��Ϩ(�ݳ]�Q���ד^���a��0T�i6�����v��:���H��h�f��H ��s����}U)��̬�NJ9���5KL]e�:�d��T�h�s�wgd�ۭ����<j�������M�N�{�$'��`��62�Q�����l;��uOy���l��xڢG��N1�BL9+�n�֒Q��-�>�Yƻ�>��c
�YO������m�<�8vA�0&ruH�Iڻ��*���}q�%�x^*�b�eV�9��+Lꥻ�U��6:� Y۽wa�]0�&C�n��QP�(A�����˩�����+����Ս�)��-��� >26� �w��=�;jE8�T��Co.���Z]��9� �u�:����� fި-��ag���4HA��W�M^ۗ�a�TDCe�Pzkz��D��ْ��b:+TfK߀��s�^n�v Y���MLt3��7t]� @"%��0�TQu��g��&l�[�ݗ<g{I9��x�v������R���=mr\�t|��w��~$�'>Z���Χ�}~����H?����ud��G�	R�{����%�l
�����ۯT��I^��ً Y��� 3 `��.�nˎ�{�Q��..!(��sAF�eѰ�	�ɡ�D����9��Y�ʍ���)g�Y�~HZ��k�pF���r���hL�WSC������ծGF���I�\<u��ܮ+����f�~u2� }��v�@!f�6����RO����I$�'��|�MFC8#Ԓ]3[V- ��KǷr��	 ���(z]���;�\t$���wv����A� �&��z�L�ٍ:�Yޚ��'�]}�v ��[d���s���]."���rz:ֈ�"@�L'7cs�a,�������T��cu��,ݟ9������OF���3"/ܑ�y�v Y۴� ������EӿnF�{��Ā Yۭ�RZ�E�JI��43�KA���C]�V���m_[ϬD���A�S�wj>��TC�o>�;�"=J�A��b}ʹ�������9s�}��K�'���� !wnSa%,7�U�)��R..(I0꼣���d(����<&�h��?jD�D���7I��y/e����Z#m\�ᙻ��k�Jn��-�^&�`�\��../����E�w��Ĕ�ؘ�A��&K����1��c
�Hl&�ו�0�R�ɿ$����qE(�ӈA
}$���o5: ��v���Z�@Oۗ�"PZn��J$�����������ݷ3�jG�Ľ[���P{v����v'�f�0'/n��w�����뎺eب��[\�2.��G�|����B֤Y63.<���2I:j�Y�q��	������Ew����'z�]�]��l{j�P|iw�Z ;{���J(�+�vN	Rto���a(%L�I�V��@n�;�� ~\����#��8� ��� ����}n|)�DB��u�dfv�Q��oR��i�@��� :/������m�p�p�	/,7[T���Ԛr�f<x�T��}�X�t^�5C�!�*碷���u7�۽�v� 8?4�NUR�Xo�{�}W��R6��Î@)lyg��=�2٨e6���2�5܎�,0���W
e��H��
�&��U�Ք�LHa�����U�Eà���u�u�1vGvk��qv�$�q����GWVv�v�ݞ�s�����ٞM�l����8��;�!�{<��=�n�n�Yt�qrP๡9z�y��ѧ�r:����}��]s;Vê8�t��9{s���{m��t3��C���Y��v��V�R�6�a8�-�����d1�3r�r��g�V�<:�l)�a�/V��������uohn^ܼfs�֖Mԯn-����p۶�`��g�o5F��e�"e�'M]�'����, q|ܿ��=fc����þmQ 	.�޻���cj�,0�A*�yq��Ң#*�{Y�]3�����,�޻� �nb"%�:�j
�6�����)D(I����*����I,/�V�H<�ȫ@%���q���Sӽw~H�����)J����� EM%G+��U���n�)��p�AU���� q|ܰ FE�~��x�ҝ���
�8ۢK��X�l�9G*���(w�ZI$��Z��t�:���i��m�"A��!�d[���RR�p��:�<�Sl�]=��HC�En+���ÜO>)�fO��`�@����`$L�T�.�� "�Ғ @+ר��Q���[���ӓlH���׌߫	82��,U��exT��I7�Q�*_>���+l��u�rK�>�z��v�YpkS�A�17Q����!xs��\�Ф*�t#��X�،��ru�4��^+�@(��u�2-�t@��+[
h6�򨫭�BFͤXa2\8�T�9�L�I�S��$�Ui�9;���&�4j?4� �y`[��w��nȳ��tU�����7���y� ���`��yR� ���{ya�̈%��!��*���2L�}�($�]���ʅy�������@��U�{�y'�E�Bj�3�����9v���]��.���l5��k�U�煼#��BQ. �Y��݃A0�����G2ۢ A�<i� w7��c�����u^�\]cj� E���$�,�m4[)B)�4:��J���d"�?^�ޡoi$�~��V�$���N�n�^H1[/3p�/�Q2w{�	K!�G|L�{�f%7��1������9�M�{�]	p�W��ͭ>èC�((�6X�6U���s�G9�e]l*�]8�^*䔻��]ٗ1u��I�VV��(�s�ua¯ws��s).oo��{�3C8��T�_o�-�.���:sT�OR�&�d*�R��|6���m>m�C�)�J�$�ѽ�\���fv䶢V�A�z󹊗w���00�\�>��i#��je�[���Kg}�`9$�J��,bÒ��z����RYiu�_%ܾm�Pc� ٘�1�ޗƢ*�r�
�u}�IX ��ը����c�1]hz��-��&�.�]>'�:�$D?J[�)���dI��>����yX�o/X΋GwH�C�CI)z:$��,�)�PwrN�Z}��+���k'X�[��s�z��kE�<�LT�+��mLy���ѭ���|�Q���)�c�g�V�XLկ:t=��W��oֵ��aN��`&D!01]C�,����]�Ry]�od�D���ײV�uwݖ�����i���I��˽S���A�YB�8��РDwr����d��Ҭ�N�Sy]]�oN8m6��[D$Z)����ں���������;B�� ˌ��H[2n�5N݅iĮ2pk�=��jL>ψ�����4��^�v�$�5Ut��\�y�����V_ܣ�X:�S�,�Ө�ͽ��CekYy	�-�U�ǍǷ8�V�dLdD�����a�V��"���b.%�Th�p��V�'�0���P�2�ȹ��z�c���B�9Z�tlpjjh,�.�n�6����R�K�HK�)J�Ж��(V��K�Wܹ��Tq[��P�hUmV�5��&)r�L�SX�ۍʆ[1�c�e���q�.1��V�\*��B�fA[3*��[3�mq+QLn	B�s�*-���ZZ�[V�hˈR�*,�\F���Uq��e��v�<x�<���p̥-T1��+*8���-X�2ڶ��ˎDA�U\�̮F��)c��j��ZU+UұTn\��L�32`�����Z1���ƶ�AG��m[Dk�.fV�J�5X� ��2\��X�J�[K�l�r���[,�c`S;��vCgq��r���rr�.�xG8q��=���p�U@X$G(\q+�8�ihW-�Eb��es�1�6ѕ��6��ɍikKYR�mU�\Jb\Jb"�2��W��n%k�±�b��r�#e�r�Fcq���m��K���<��B����<�_ m���H�7sz��@�{eL�@*���%������d��t6Ә��vw]�t_[i�D��)�Ayq�|e���}N;"p����
����h�JK��H>�Utu�����ٯ� /sz��D�>�*�l��S��CR�Y.�LKk�=�r3٬rvz���:���
�8���lLD�ZߍS���@�]�;+_�D��v� /��@U�o�v�Ҭ��Ey%���v����bDKo[t���=�����z� ���tH�y�� z�ю����~ŕ�$�3�	R���y`�Aћt�6|vԅ�OFO���F|ݙ�whH!�]UI����m8�0�Ա�\�I���� [�F@ ����I'�� ��ʅ�?*�^m�fiJz[V�{)�=��tV8��`ep�n�����3�ó
�2\��z�L��NY�:�j�\�MZ��l�QJw �R�Q>�T�ci�Y�/��D�G繨�O6�H�R �#;�U����:����wc,_�U�5���ub��l��'a��t;v<\؎xɷ]����QN��8,�ͻ����C2��  Y~�~a�1�Ln���eT�e�� ����|��g�S���@��+	�r ~9z��}���5צ��f��� ����L���+�R@Os���ƅ����%C6j��bDU!Z�� |ec�� X��B�:}.�"fW6Ȉ2���j\�Й"W��%Kg��^�N7>��.`� '��R Lw�V�$���{�����69�:�&��������6��a����r*Z�_Oy ���y罙�I�p���C�"�[TA�n�sv.3|b�P��/ww<�uN&��wwqY���ϝo98_�Ԩ���ؾ{oh]�e���CgT�FB<��IU.|��d=��w[��	.)��pD8�I���FT��I�N{#����kv3�$jv�f��:��uuvC��n0�s-��ee\v8���z�q�t�nL��"�oO7��y�P��G��G�Ք�P'v[���`�\X�Ok]ø�m�)2����݌u�vG��V�r�P9��,���1�ܶ�t=v5.y���Ōg�nׅ�`v+�c�Y�f����Kv3S7���a�۴�훮v�b%��`cqj��U��_�7ϙ���TO��G$.��� \�۝��G�i�v�V���l�d\�P�����I�pE �w���	uW�f����ö]s�W�s����H���,t���G(�ϔ��:heuK@ ���vD7�F��}�=��� Xڢnw]�1��B�$�bDN�[]U΢��K@���jZ���޻�� ]uͽ�[�8��	�I��͉H:b�&�b)�L:��ﮉ$������y��@��@P���0>��븋�u�6�;!��G�z�۪4<�����Q��(Am�[��.Q��P[\O+u��Sn���6o�ߟ������Zo��I&�;�ŤI z�U�^<Uև6lwE��'�o]�Ix̝��S�LD�ys��R,���(v�a�����*�z��-���I��`���(�1m���̇k9�fa��fO��;�����g:q��Ă3k	0krY=䯳���^	�=5H�%#�t�[<{�:R����l�!��>C�C����/�4�|A���G�v�z�� _n��� �����s��gɆ�aT�Trx��v
����n",|�0���}v��<���H��wa$,gM%��2X��[γ����[�|v(je���yw �H]z�D0qo��skMrP�D+��B��c�/0g�s�9���v+,b��;�������߿��m>����N�+ -�t�$ Yo�����s��u��݄A����ە Æ�11T�y���ڙ��W���  #/��� ���`�H�P���������H'��l�Ğ�J��Bڼu ȷ�:>@|ܗIQܕ'a����5�{jB���Dy�Ƿ������v`���PT��Wb���������v�D��绊bV��%F!U\��r[|�����}��h8n��[��h�zK�	$��mT0l[ʘ����v����y��Wky��.�m��q��c�T��Q(M��
��w��71[G���E_7L�.-�LC����v�" �=��w���0v���C�Z�^v������)6��Q�u��;s̾յ��������;�u ���4�A%���v��]�N{}K�
w��� @�%�f�$�%�	�4��eش��X.)��Oo���6 ��9��{��wh;T�)ݓ}T"��� �ڎÆ�1Jm��4��w;J�Fߝ^/L����8��%Z@���F�.^�R�Rz}*]W���߈��9?��}��� u��wl�2��H��)�Bnj`�X�ћ[3�^Cs��Ѽ{{�͗�N��ջ[�����Y]�!7@��Vڣ��Gr����;n�ٮƸ��H�YSM!.3"-a �{}�+���M�7���A�b��3,�f?0����@ ��%H��ny�
��YuwY$`�6M^&��E�Y4c����=]1�.8�G��]D;���~~�o��c�T�%\�Ɯ� ���_� �J:�Da/W��=���I�4�c�h���w]�Ic:q(���X�
��g�>wT����m�Q:�r|@,��_c��s�o<wT�H_g4����h�Ɇa0��ח~�� ]{��|�O�o��a��r ;wy�� ��`��=��31���0�Բ�1��Sn�I,�˫��PA}���c�g���n@NU�ݤ�a���!�Q#����� �4�Hܟy����@.�˻�]{��"2���$��Z��j�^z��!vfZ�`�;LO��JK�W(�蜛��7q�]AA�ݢ�Pܬ'�psG��q&�LP,�ۂu�YD�y!��GV��K�Cm�p��닱��n�n��������c����7fݮݷ�J���]�gm�����k��۹{g���u�۞o��]�M�	����pw6����N�ks���=���ѳ�dO]������ԇc�p��Qh��^���gkcx���/4�l�q�#��=�냋��mv���p]=�t;�a�g�<�%�zm�Ss�F��%�A��[ŵ�d�L��+k׍v�u&��/�����Ce�I���q�ۣi/$2�&�$	�������3"�D��U�(��
�nd���z��0�,*�9s�D� WV8&��hA�}�~�H��r	�$]r�_P��xsn3~�^H*g�7wb�`���I$�ue
 �P؜���h7nNzgy��
��ݡA�^�@R��4Xp��pj�G]���;8(�`�GuK�A=][T>��J�[��ѰH#6�|$\R��Cp�11'k�(P&�w�O���|];|�X3Y�A$�uu{ws��g��r2��J�����N^Nu3��![O`޻@.�у[��.Yr�ۮ�n�߹øCE��8`��F�s�Iʺ��|On�P���U9<"T��W_M@��Ȇ�D�NP��ު'�7���Vv�H����E�
d=��E���4m��s���0ne^�Z��r��L�jC�\���Ep#��B*��A�7�ݧ,�A>'�Wy^�ۻ�@�cTĖwZWס[�~����0�L?&P3�;TI=��4I&d�!a�[wv�N��I]{B��n�U�eDD�DDI�S��~SY9��� �۠(�A;ݽT��s�
�sO��eME9��pXp��pj�:�;.��[�Mi�i���Jݾ�� �f��
�'��Ϛ��=���E$��^�@1�D�Wm��/4I���=�8�-�/D��W����~y�b ����WfUM��MH<��$��va�\U>���;;z��1Z!�Â�0T�39���3s��E��}6�*�$��ޡ@���hN�d����$J���M	8��%3սTH$�۹b��ZG�|�Z���N=�
�����1[����3��$ѷ��C�6Z�Cq��V�t��*ZΏ�ُ���
�{�Ǌ�&�q���]YovxP���$�۹g�N0���~L)�z���� ����I<��$	U�\�y�`�b8��T�$P��*"�b"^��> r^�w�:υ7z�_�l��	'�U�T	x�n���<���A/�ԉ�8��*q���=�F��@q
r�>×�*t�ApRu�3a�చ.!���ݤ>�� .�@�W�{|ƾۙ��u�TH'��]ϙ�Ȣ����!�29OD�װ���M"~��P W�n����H+n��^��Dr��=Vh��8N*G��2FU_M`T�v]�mU��8�gn���wM@��6�C�0�	N�oS��<�5� ��N�d���$3�z��GT[�ѕ�o(NbD���F��\�]�e��vذ��ݹ�|���bt���@g����X���A��ŭ��C����x,�dV��f0ɃTg�
�v��W�����۶6��r��H	��J�b��a��/+��3�
�KF0��gBi����k<�,���G=B����[o����LD@��DB\�ɖ	ڭ٢A>��T���qQV0�o�I;Y{B�d�Ci�E6b�;��3�X��M���d�:�6�I��^�����������;�
p�� ��$��ޚ�IТ�0�#��Ő}�Y�@�H�����h��C�Ⴈq��=�1D��H7��^�A۽B�H<z��R�:g�Q��,l�P�*;Se�L5��R'kz�ĂA��r��Q��s<DA";�d�}w��+���۹��I	FHH@��H@��$$ I(B����$����$��B����$��H@��	!I�P$�	'�$ I?$ I(B��	!I��IO�H@��B����$����$��B��IO�����)��Mч��(��9,����������1�A@�� P �P�� � ( (�B�  (
H� � A@�AFJ�� �AI
�(P � �T�@ R�
� 


JE@@(
  P���@%JU+�hQTUPHP��T�di������H���(ki�m"��mRB��
*D��*!� �GgP��"�H�!%!���� ����  � $�0!���,���� Oxz
p�=����Ξ����� ��L@2+��@�P��� �� ��B���yҤ�������>����;� :�H

 O�  >��(��
�%*U��`�@���d ף���ܤ��z����cҽ�p��'@��PN ��`��� �@ �   �g� @���(Cy�� �����{ �{ �� ݃y� v���C|Ѷ�u��9�����@]�� G�  � ���*��*D�P�E����op��`� n��*�lF�o<�ڣϠ�f�m�n����gTH�ʩM�ZUx�g�u�*H$U�  G���z�J��J�n�*�b�PN�qRF@�E��ݺ���D��DwgUD � �  <(�eAIi�H�B��
�=+v9P�@�F�(b�\�
nDNZT�]�t��\�*�vꀧ8��&%��P((�  n��Ί��ª����r� ��uJ�"%wp:���ħ��3��lB)ݎ����J���� x  i�P
J�f(�����^ ���cwrJ�vuQ)���Qn��)��襛TDd1R�"��A.mR�tBJ( Px  �;6�X�s �o����u�A��9P� h݁�T���O<�a�������à|      Sѡ���M�#C4��Њ~LBR�P0 �#4����Ѫ�jT���ɑ� �0B'�U(e)�@       ��RT�D        HH�)H�4hѤ������<!�'�������~����o&?pFÕl7Z����f[>Ԅ ,$�����!� %����  �� �	�6���� ,��>d�U�O���O������R?�����`( �"h:$v!$��4�Hh	��0А�����ۓ���������_�	 [��9�H����W����d��G�/Ϻ��$C��?wQt!�o����~i�Ceq.��k��z�e�38�����Ɲ�so^�emGZ��Q��x|��v�K�Ȇ\a���3�4�+[3wC�:��4����=x̘,���٘���s5��6MG�9#TY[��˫������7��݂�mbձbs3\ki�����'�f\ڨ��"���۪{p�R��Xڔ�b��s�ٹ4�3�(�DK�3`v]j�ӄ�*�݇M�#$)��\��Q���T��U$TC늖d�7#wG+c۔w\k1�D�4 u���<�jvZڈc��-���kl�h܍�d�N��r�\�W�{��Bh�e�DA�i�--2�7u�̏-;�s����VN2�.�ML�����5T�������N��Xw��Mc(�,Zw03�f�Ww�����BK�kD �%y�e��0�e�lj.�9 %nA�[�fi��QV�� �ф�b���!�Q���ˡ�2�p"�����b��I�N��D3��ؘz֜18兙	�9)b���p��NO������%yX��a��1�hISn^�bE�lA{n��T����[ӕ�-2�hj�3o�9uى	�4��X�c�}�g�b�>�s�$]��Ƿy&kjD����\ǎ���Ů:�"٠�J*�e�/P�÷�3SN�;I�U=��pb����Ԩ�ݭ���9��+&充%M�['��QSMJ��m㻻��2�m���M� �X5�"��^}�A��Ŧ��ׂ��f��p��۟˳w�L�U�(��٦��&&�ţ;��Y����n����Mڄ�k���c��w^TJjT&�Ǯ܊Ү��*Z��P�m����\ʇl��շ%�*Y�2aGY�Y��ZT�i-��j�$��uy)��i����0�b�Ņ6&}b��)5�:�7h�3j5���P��O��Z���:U	;�c8�oYVL:��&{�2Q�ܱ�#di�̽�0�)x.lV@{��L�t��*zʕ����nk�R��,f̄�I�_�m^[�y���
uf������n�PRe^Pl�XF��`�@o--�;a�e�n���L�[���u(�%p+�jjv�[�"&�b�ɯ4�!PT	��G1\yP+T�wZ�J�j^|�M��e^=9�0�h��$\�vE�˴��װ�Lt�R;I��Rj�v^��J!d$��E���ŗ2����W{r)�/a�T�����s2���3.�4kc6KZ���2��2�B(;��(S���-K��YL�k\�����2��P�i�mXv��.��+*QKVh	�R�7@ʉfR�!�ܶ*�xB7�A�1k�[�Uk���-�4΄vd���û�LWO&U����w��m f����Qt��6i0�R� q��t�s��#���z&l�]l�2�t�$��	P��y@���x�wYz�ʄ�W�X�e2ł�ŵ�U)�N����P�m4�^hjdYn�E�J��mͼ�R�/Em��g�\�CBdᄋ%M�rM�d�(1Ӽ%=�h �z���6�e�U�D��2]L߰Y��qO����� �זU�q��pܔt�u*}�{��I�Ŵԋ�PS��iT<�XԳ�,�t�/j��yw�t�� Xf�6��Ȯ��i�e�&�1i8�ni�7!�+u�r�B� ��&��^\B��諊%k.�$���N��jk��I��)mjX�(��Kh�);y4;%�)���� h�����,0a��sn�L�Vǩ^K0-5{�2�Eh��{��ӏ(̭���
Vr\VodOS�ܽf�m��!��y��4ښ�ұ7VX��,ОF	�%�[�[8A�(Ix����t�*Vs74���Φ�ڼ��_�L&J��DE��jVj�D�&�}d�X�k&c*7�D��0�V09Y���b&V9�N�%`5���Uкv��^j�D��f�"ݭzjV�S�j�Z���6Q�f���Y��%`ғ�)%D�eX�Xw��Cia��*z�N&x�;Y�I�5��FX�c��>��9R��q��̥�-��jX�.VT�1�m�y�ٍ��+(�
a���;��V?�����~K�YY	0�ۦ��z(&y]�-�V.�����Gk-K�C��,kDWt`���j̷yunDBfe�{�)c����5��XfT�Le��/&�ж���vJ%���P��r<[?��%wk��]%�:�j�� 8��)���V
9�.�Kյ�4�1D�;opl�ܻo&EW�A�YӔ�8�M7+En���%�i:��d�3#$�"(��e�X�WN�Ǣ4�ڵ�f�3z���-�6���V�ff-�,Hij�hִ
Q�u��ЙA��l#��A�P@6��7+-�T��ǈ��j����T�I2�@ĽX蛸��뫴��qR�hކ�RY2�����"�!�7�yO)��F�!�y	�cW/oL�x)�'6�Cj��k70 6�y�Ƣ�Zu�!��oEL�����,гtX9��^2m!ʏ�w��i�K	��7t�]�2L�3n�bѕuke�P�;�H�{�b�1Q�{R`��ddL�[M݃E�wy����ݳ#�w.�08b$' �Է��#u��uu{��{8�a�Go�S7}TpT�ӢA�2�T��m�#����7���V���ؒR���<j��T�8���Ku�H�"���rٜ�����뽥fv�7P�N��!YN�gsH�F��{v��d]uzV �V�N���`m�[��-��dy��6r����數앆�[�P�F޽9�*�ǔ��m�%��j�ӛX\����j4��St��nnط2e��۴L�8r�n��K!�kZf!n�������^!��V�y��c�j
��͕GJ�X�t�C��%��6���^DnV<̡�A�T�c&��4��l黵��fR��J6�`�-V�J[FGx�K#>�:Ұ�9��P�H��P�bxT�b�H���D�-�ȧ��b�c��^�7rӊV��uq9��*��ב��P�?n7%YJ�
o2J�յm�bٱ��gD4��⫨�: wk&#bH���yG%ػ��ڙ�²�ܐYN�j�Kh*��HB�t��b�h���E�ɑbӚ�ܙ��#2�nyOj�����2N���&��qމW��b삤��p��9X�P�5� �b��ͨ��(0����Sl+��,je�h��͈�6�Qn��)�em��B�E��TR��	����ۓP���N�8)�J�o�wP�����uڦB����e�dD�J�Β2"�� 7jАc�#,b��A��2)���:�A��`1�(���vU��%���,fg�#C)E�[*�s-"5k����{$��d*sU���KK,�VL���t	��WO9.͎���g4Y�,J�O�X�Z �rs`�Ow BY 1)e �B�ђ̆��6m�6t0�4�t ���rv1�����ʰr��O+ld��VB�31�u��]j���!��Cfn�6�ݺ�GΪ����S���y#T4i`b��;Tj;D���*f�o6�Mˋr�ݺi�W�+Rٗ�#ga9����_O�[�:� X!��Z��)���Lm��r��VG�Q�jà�5�6�ˡICX���5V�d��8��.\WH
y�F)/H����K�)�Vf�գs]�m,y���S&\�+�b���Y� ��U�1��8�J��%��-X4Ed9��ŅX#���h͠�ޖe�b̙���VQF�̆6擫�MB2%ܦ���`������o0(r*/cp<b��*�Y�-81]�V4�G�e�s[�5�IZ�[�fV����5���f��ˠT͐�g^���f�{j�d��pP2�˩�n%V�kW�L˰��wY{������pS6�f�:2�u����(��bn�8` ����RHt��(@�F��bXΪ�M$RKl���Y.ܬ�,;�t
�YA�$�~ܲ2�J-�f�m�����Mz��1wOvfLռlͧ�C�n��{�y�%���3 ��u(�6��r�2�)�i�4�r�n���g@�P2J0V4o$-�9\cܥ*h�s��u*�\�v�b�����5l��,^�gY����:�^?��ot���K�V[B�#cCD���5u�w��PG��`�����]=�g�M�eJ����od�e��[!֡ne�0;+C?	2���hE�����)me�w�<����U�.`ʵ��6��u��k;�YO�����t�P8������T�IWX� ��F^%�]�2�������BƯ�Nu������D�/&k�sfO�T�)�.B��v3���¶��n,c�5��4��X\���,*�'�57��)�^��jZ�#��NIX��Y�b�ӆ�8���XvI��lV��r�=Wo�[RK�2�1�D*1�*)�7skfV;C#�UxӬ����J������;���َ��=Ե����t�
\am�yr�g[�&fهGea�aP͛��ɴ�%�`�ܥ��34���:wcĴ�4Ę�n�~P�I��V!s�N��K�[I�;I��#L���� ܹ����j�	Qܸ��j`�p�{%J�w��r}�lCYW3c˸UB���[�`"3�B�jݩ�u�~�2)̊�@)�T���djq���4�m�ؗ[���v*n�����^
li2n�Q�/��ܣe���0m˺9��ۆ���A[�n�U�Q�L�a�N=�@�P�Aŉ���f�l�X�]�v8�����˭�	�N�OZƆ�8H_E[�`����kUe����S\�jZ�Q�wA�8�n�j�$E�%]���r�ɚ^�e�}�:8k4� ��҆\i�z&L�6���ou�:��Sr�cK�5�f�,%j�ګ���V�zT���N9�f����rn���j�I�]m���n���X� �}8�T�x�FK�tg����1�l�1���sn�]-�o7��TSJ��h6/t���,�x��gh:8�b��R��NO͕w���vV^���1����&m��k͓E�+L���5��Rd	�����ҽO��R-�e�Qn��L�㸅���b�fJ�k+��X� ���[��iOmHR;�H��"I'���D�kkZ%͕b]������x�Ve\�v�W0�B1���ӛ�b�#m��eV�H�&�6�t$��������@���gV
_2�pSP�x@�D�0�԰�a�u)i8*�p�ԻF>���x��&^��@���OPɥ`���c�U�T&�;�
��mٙq��@{(ٵ4��Xw��f�70k^���TrL��8��-TwG�u�b�t�B�P{O�ޓMҒ���R~36!��l�N��$5�i���ZΓy�b��c7j܃4\�r�V��K�J��\�k�6�Y��ʸ�UM.�q`Ni���3o@P�X�X3❯�J�Y�W3��`C0��,i��1�w��($	���m��D`��p�!����r�X�Fnv&N7	�fI����8T�2�5vиM!U��ɪ+&��*�Q��;N�S(��
��ZzlP��Q�(Dl���=�&VWz�V�?K����u�r��u���LVX��(�M;YA�È1KjD˛;�A��e��dO��9go���p��m*�2fS��c�0d92�����Ԧ�5c%I�o��2��
�3C�G�:n��6Fǚ��X�"\���4�	ZΆ���iq�%'B=����c߭�]�;tw��hh8�׀)�d��j���ù�b��a2��n<�i�nQ��6��Ɖ_��(��m��&�Y��̺j�4���nU�E-i��J]w�f�U����Â��lU,���*B�h��M儠�3��MZ��)Yx���ۢiZ�]^��QRT[��^�sn�+�yeA��=ҏќ	���B�GF)uw���Ha�J)*6�F�]��еJh�{B_�-���ݺ̗wl^e��Nl��1��$�4C!2��S`yX.��ȱ�!S#q���DJ�u�X�crb'uv���K@��jm�kL`�A  �	&�b�"�&p��k�'����JE��U�+[>ɚN��X���I���mF@Vj�
��j^ �f�L��܌"4\���r��(�����.�-�#�aֽ����\����ek�b�A���e���=mFge��͛IX�L L&��\����x�F4��eEB���-��cYB�b�t0'��*�4����;�������a(\ݿ���'m�=+91���?��h�R���ay��[�����/�ç��U󭦔�U�/����t顓��$��m$��$/�Ēl�#I&�m	�` M�$�I ��N�@9@9@xF�I�$&І�B�	(�"4$F$i!&Āl�6�B� ^8�'�:C�'��HI6CbHM�mH�/q<q!�
���q��]ܠ<q=�/p� ؁���6$���!���$�I	�@�Hl�I� l ؒb@���I��4���J0I$�@#H�I �Alm$$�Ill@�m!$�h mhHI�%���4�#H@�@؀Blؒ�h��@(ЛH1����~ϩ��>��O����������� J|C/5̀� �/�$%�߾�BF�p,$� �9�Ƹg�^}��>�1+�3*�:����X{�B���!���8�&�M�2۫N+Dk��qǄ�#*Ң���w>��<�!"�%R$T0w]���©�z���'�{T(��{��Ү��p�Xi�u���з<9'�9���Z�9�Vas �9���BW�JԮ��s7�ঽ�JZ�*s�X����գD�}���חY�)��j��kәr3�Q�{U�1�L^�iz0c��8���Cn�.Z�av'S��Vbլ��n��Mg+Ӑ�F4��y�������| �&���w��Ϯ�tN�/�_d��y�T��e�{��3���Թ��VE����330���S���f�Z��H�n�3zmd�u]�h^-�7M=�_5�h�NRo]��r�z�b�M�}w��y#�`��zvhY&n�t�VM�2�/�c���j�Õ����="�z��G	Bi��W��jvҺChe� ms�3�҂ͲVa����w�ȴ\�2>x�oiC1��ͽ�@V}{��mAY{|A
J��k6��q�N6l@�7J*����2���{��^͏+��E�XZ��U�����Q��R[���[�nd$d�!6L`Ɉ��X�:6s@�2�}�C,mK�0'Gt�^m�!���O����W�Ln}��ҠBw�uf�76� ��u�l��/$9��b*�7��.��f-��+9XZgq̚��j�󑐪+Bou�����&D�-�7,�fK0�iE�_[be�̬�qwT��_b�Y�#�����Ӿl�v9/Z�6�U�-f��)��8or��"mGr�\Äc��pՈ�&��\�]�3NVe��)2�4��a�2)mN�"&E���M��+R�b׻��u��uN����Mv�n�rf	-�B\b�yC:g
ʌW�;��<�ʧ��\5�-�-�����vtT�����#mb�.F��Z��2��7SiT��m\��y|�tM�{2>���A���)���=�.9JJ}H�R���̤�WWTd��ź{"�j�1ZA�Y`룠��f��8��c�T��2Vn�:�n�Z���{i�������/fF�[36�۰td�r��	�DMT$�����/D0�n� �"Ʊm��2�)���A�Q�Qm�4֝�V]%���&M��͐��*Fe�o��J�s��bn���[G��3�4R6NB���rƗI���a+	�f�%��7���0:�J˸.���{�ҫ9;vKtfV[�zQѸ ����Y�^��\��������>��h�Qn"sX:�c�p2�a3lKNAx�S ����t)��r��:���wXYP9�P�q��)��f�d��;5���BN�o30��W�r�sJG���o6��;���lg8vgr�%��z�n�I���l�J�X��zgtޤt�g�k��z�{b�L��� ��������V374v̨8S��YS���b���;[���nQAʃ�D�	q	����T���S4N�f��M��������F[�P�|�i��Z�mH��� ���^
�h;V��T�ΦdǏ�p�4,����73:��`�h�����+ �Y�cnn�)@m�!�TT_gN4�+&��X�]�^��u0�i���^�5u���P�\%��3!DǮ�T�.�Ɖ�y�	��.�69R����B��Ժfn��45�f\�7����OGe��\k_f��U�u�#����:�v��`f�w�a���D`���ś��	 Gxs�4��k��z�l����k7�{zn�nEc�.���F(3:X�������vZ4�����j�Lu�nuՉI�&9���l ��f��3ya�DaxqL�-���.�VXfKX]};�����)�N`�/��ڒ�.�i��[���Frl���J�et�����P��_}x�]�JQ��y}J�Z��e���-�Ww�����-մ���9�|z�n^뫹��&���2���rKY�,��L��0J���;�H�u�Df�|�B�� �)3mS&�;�{Ȧf<��*�)�^G�=�n�s.��R��nR���"L@��WZ���eЭ���(݋n,I�|�;# �a�+�TFJE��?�ۍސ�kY��.�+th�)M���
"���ha9��D���P�z�=bld�I��e�J܂Q����EAM� �]�x�Ջ-
ݺ�S���Y�f��Z2�	n^�w�7r릯�����b9w��&�=���8WfU��M��;MZ�9�jn�2���v�s�f��d��*u���e��`���[�MB���Ky�Vf0�5UEk�S��NC*`a�/,�߻z�ykd���"0˝�ŉP�^�k�3�����V�<>{��Br�Mk�ӭ�p��0�)�U������>�˺�|���Fq�}�Љ9S#��f�Css��찺�ŷ�b��-W|Oe�������A�M��ѣ�t�Ϋ�uG^��צ���A�30��Ӈ�����ɑgg�l�i����v��V��=riVw(;�T�ݕb�^:ܱN�Xf��[��Lڄu"��8��KNI��7�����˴��4����@MG�Y�Ff1��sVX��8u���.K��wT����i�"��]�X��������E�ԃB��2f['d�?=�F��Ħ5o�`�l��Ӥ&�U���U�1����zj��������Gu=�s�Oq��qա�.�p���ܯ��قsK��*���S_|3k���CRs4+��of�������zu]܊9��
��;s"Ru�-6t�J�-ݥfe�Iv�����}Zp�/j�b��[�u��l��j��׸րĤz3X�^�9��<T�G)�/z����Ja7�1m��d�d.��7��<Z���E}o�hHz���#$�Y�Qg"j�t�FK[�N&�d]6���c�
�}}j�݊��d�=�o�<��[ZzR\Mj�{���N�c�v8V�4���۷U!k�XY��4�
��JU��q�����3��6(w��T�gi��Z��b��x���]�^�,����"BM[^�*#�ޫ��C���%����ۦ Vf���7��$e��Jx�姗ǳ:	[8���%�ˣ��:���e���c&%R�ʭe�%�d�ؤ˾b��=Xs>(��9[�:5�t�^�s���.d�f�g9�{���e���!k�2��o[\Vq�������Vn��ĩ��ʱ��aH1��r��E<D��λ���$��3(�@̇w:e	�޲�C�3�Z6밾��73.��{���7$J�.����N��eͣ����<�t�/�J8���.ZY�(����f�p��i�8�T('f�b7����ooa���v�ۅS���z6�8x6��Pa<�X�,�uW8���Y`��0=�I(�xG)]`�)��T5)�:��uY�xa.kYVa���}A$1j]}��R�O�*����b.�蠠��Q��B�Vh7z5���l����EZu�e�}�󰙫�-����;2�!��i�Y�mnc7-�}Ov%����{5vc<.��j���W2wA����N�9]n-}�$���Է ͜&X���)-�{������E1������­��Y-gPvL+��g>��Y77c#6]h��^�C9T�Q^*�]��F���OA�F�8�X�B�1a�%%S-=���J����Cu��/$��R�Ї�d������5j��g���ץwָ�X;�ǝ���tJ�Y�w��˥�.�Ù/i�x�ୡ�̻�w�{9�Y�p>l�X���,��'%*�#�I�������N��WJ4������h��IO-�t>!ږ��3�`��ᨪ�՛��6Cl�r܂V4z�U���RY�jŒ�k�w�K��հ[�~��U��^��9\<��L�՝��E��wF�J�V)q�'���L�4yv�=��+��A��}o&�ղU�JM4	nrV�k.&�4B[[I�&��݆ڝ���Z���e5��;*��r_s{f�Ռu�8xV-�7 ��������{������|�l���ܵ9뺛N�p,k1�yյ��r����\�:e+x��{Fͫw��{��],��p)�#"��v�db{�m^��e�1�z�Ö�Ԫ��6�]Z�*wSP�����o�kkO4�J}���a�a�ؙ��
���-�n��E��q�[��2uL�/����/3��f�I�7�6�"����U�y��H�^T��<��skC72T���M͝��U�jXu����;8o��]��F5�zzXܑ��ya2d��하a��Wi�[�	.�͹���ޕ60d@�
�za]��i�@��]�M2��4ʈ�F���X��R��Q�lp�Z�X�k��w�\b��X2#TaBcD��n�CKvg(kv��q�o+)����:k˧�s^�}]y��T7�Եc�.v³�Ё�e����7К�eE���7��q�Z�>�\��r���˧B�j5fq&P���3&�RB�w�+ŷ�h͆�;s�ޢ�"�;�c��@�4*��L�Y��W�r�`�{���]�C܄��W���æ�nV�k:����f7�K;iح�J�'�ɑP]Ks����b���u�7��/k7U��Y��ˁ��9�X@��P��v �;�j5՛���9��b�^®�QR0]17����tY��LV�"^=�hL��[}YGD��VW�@[{3��\ȐΜ��{xC`d9v#�.�̽�n��`�]�{̺Vu4�P�fQл#��񶞇)*�
8ǈ����H )��@��J��+`�m��7]�٪�g�⛚�强�����N��<�o�E�S��TݧAVV]��k�sW@��h�<��b��9�.�w�!�e���Ǆ��K��u'��w�09@��s���]'`�`����nu<����բ�)n�����,�AGd̶�;ު�F�,	y��P��і{9R�3%�L�n+�f��a��͚{V5m3P��e!oro3hl�^o�\՜j�Z컔>��q��w������Λ1=5�D�k9f�N�NU�}��2��p��G-�AG�X�K�����f�dͱ*�jQ$=6�D��� �t���߆2�.��QğCP�}w�Ok�ƍZ��-��7GXz-�;E���7��7�PmF�(���f���*�ȥ�T�z��|7�fni9�&���kc(�5&�7�)��(��N޻��V��3)K�eZ��5#i��1�b�J����IXX8�-����o(b��N���,�ɀ1.1ִ@�?>6@��J�΋��٧WSo�uJ�սceLm�z��	�q�*�c���[��`[�.��!�������K/3��f��dN��aR2��܉ybo۬ý��>}On�H5�ME��5���se1۹���H�̼����7�o��5qޒ�f���D�-]�DWe��0��n�\��6h�]}�.I���m�B����t����ݬ�����i��3���0v�[�{$;�a_-)倗Vr����e��pM=̕��5�1.�6z�U:�/���X�����f]���_#�W$|��c�^D#�;��:J��G�z��Z��kr�*�j�)Aw/��/Mg��Evgã����$3vjHp��h�mV��:���X���ұk���݊Q� �:s�j-��}���S]�}ײ�N^3��V�aA8nӝ��#)�Ûv@ԡ��j�
��5bq��V�K�������d��� ����|���'�m�΢�-��q*�I4�\����/
���*�]a� ��f޷�/��Л��a*�Z��Ey�F�t�����]����Yr	fwU���}%��Koz�S#G'qr��+��������;���x&Sg8o���aE!�m�R�
��޷4rz�rM�x�u���L�ʫ�`9۫�xx�+�^�ә��F�+a|;a�u�+k-
�7`?`Vi*@��lY����[����ve�юv��aG�5�(¤l(�5[XN��b!ұ8��]J�gv`U��E��)�_#[��uݰ,����P�7��ΰ��Z ]�<�	�i�xx�Z2�-�CH�D��4D��Iř[d�F"��=d>�u�����_q�!��΍۷���ﶁ�fr���F�kS�%`������_\32W%�k�6\�V���KS��[d��U������&v9P�f��9l�H��Q��h��r�j8�=��o]b�fY�g��=�/�����yۼ��)-S��"��x!�D�9����fN�Ujrr��HQp�y�����CINFXS5ck/�
����&}��c��OK�N�M�:������qRt��3n���_K�xf�Y��A��qGB����K���S�JK�`�|�3��MWYxU����gq^\�3Ne�\���I�\���8_Wd�ôz(U�8�ܞ���s�1��x5Z��oྈ �1���A�$�[��� ���H>|>�a$	��[䵣�[��W�k�RH��8z�Q���[8��)n��X�b��^1Ό�e��]l�MLң�Z!�c�On�Ѹ
uy��=<�>{:�͞E/Nn��y�oF��=@�檍n"nΦ�;T
;u4�ٸV����<x\��Yrt�gl��ڥ�Ħ�,�f�W�0�ɮ����ݝ�:���������۰[��6(�B^[��]l�k��k�En3�6N�@�C�DOTU�)���!;��#sbJf�$��`�-C� ��1n��u�klgQ�Fl*��(�(�R�;Te�f#\ر[R��P4�c!N���uWk.W������_ttmy|��&�y���uȴu� �N=#�d�'+���66�Trle�ɷ6�V�b[G	����e��	6K�Ɩ�Ơ^ʋ@���SQ����'/bu<�un�)*ݮ�V��,�-%���Y���fލÂ�m��
ݭ#ب�^����c)�,�M��i�#ۦr܏ARq��xcn�	�S��֎�h��1�6QJ�,GJK;�
6��p�b�m�-��7�Wo
�B���ld��z���kAtp��RR�J�X{0��9�&�tׅ賏Nr{�t���J'6M����O������h�z%��4�.�c�U�#ch;5ȧ�Ӈ��I�*3Up�4�lfk��C�[]��qɦL�§�7,�{LWc��;�l��vHE禖��E��1ۅhZ�c.$�"8�ѓJq��jK���՚ʽ� %�b�!L�g6E��:�;� ����N���n�i+<��e&�1�jy�8�5a��9c[[�"TI@�6-���.7<�r��:�	��,�.����\Ꝼu���	<\\���Ӯ!aS�ۖ.d��C�N�R�֎ݰ'F�Us���8�-���,ZLJ�Q���u��2��W\��<�m�R&&�)��E&&�3@z�29��'S�TM��sea5�ƥ�CBPau��X�k�g��g��!�u��f��6����t��Yph�A�{vXva�Nv�Q;1�>s�|���I\�sC�m����n��<�Cή�����s�L'b�X�E�l��,�`�R�B�pu�1��5���u���m�<5����gY䦢��r����k��c����hY<�6����`\�Ό��Ј�n��]H���y�7V1��N�G�Z�>9�:;�6��.�Y�-�p���v���i�א\���n�Ǵ�/��r��$5�>2�^��I�Vd�������Ү+��,���b��E��m��M�,�\UBYQ�"lR�ɐ$f۳ˀ˧n���n1WjX���l
�u��hK��z�\a_e��+�c��=�A��.3T��Ki�@ۓk��Z��㶸ٖl+�1��Kv�E`8��E��nmv�����V�d�\z�����-�n�-1Kkhv9�1��A�����>���*�r�6���,�fRԳ�촄	e"F�*`�s�	�Z/>=E4E��Z;\j�dr6clVީ��&q��%��x�ygY�{c$c�Έ���= 6��3m;�3�<:�x���xy<��\b�u�
^�f��۵� �$,f��-��b.ƕgMi0u��0�6�t�����a;�}��+����M3�i	�d,��3m��	��ј�\����&��(K���jX����t�^.�]���kS�	����o�kI��y���10�A�WW��pn�a��7m�t�]&4YH�$ؘ�ӷg�Ğ���c�=��f����٦r�+(>Æ@�n��%�а.�Ve1���x�=�S��9���S��a���H�x�9\6�tҎ�̚,b��F��+�׳.�8ٶ6��mNqj��F�.��'.�5�B�E���k$fjg�M�9,��&e�t��a��<�-��%i�y���JF˶���4a�Iħ�0�eU��[�x�w�n��H�|�q��c��]�,��8���ɩ1�	e,�,C<����s�q�f�i;rT	k6�ͥv����D��ج70h�LU-��U��ћ�ņt���r�h�&ρ�zPY�b�n4͹Q�����K.2)G:63<j��M2�b�����KS�DZ�����p�V�̪ilȖ������a�#�Xl/]����I����D� �[�lB�C����3��)��9�מ�JbϷ�%�W�K�����d�f;>s�4�2]������f7KfIO��GY��fJęWheB��b]�pp>N��H<ܸ�'���=��),	W��d��qv�dō	�D��a{G-۳�C����٭��IYL����X).�	�N�3Ż<�Z*L� N�;s.�um�N��2Pg��q͞����ù4���r��`�ٱ�oR^&�C��doE���y��9ǡ6{[�E������gP�On�g*��o>�'�9���6.F�˰���`=�gcɗ'��<m��n�'�q�ٹ��i�Ɔ-�@�7�q�'Y��!˸�<4n��`�1�ێ5�;�{Fk�����]�^��U��v�t���W�7KGt�m�]�4���mwY�dƸȚ �`���".޷�u����'2�p�s�l�kr�b�D�К9ת������<D�Eһn��T6�pK���&�W:^�ԭ�"��;9��\��\o�<�xg��X^4�wgX�n�Jb;����dS�̈́�R�i��hZ�Z28C��9����nvpώ�\�;��,��-t���NyNx$4[�� ��ID�Egn���u��0Ԏ+��l�!�A��Vt�v�x���j�.�P�s˻m�uh��CX�a`�
��%(QKǜ�I����f|a5�����dZ�n�Hf�ͩ�����5F6���&��M;^y����ZM��u�h@�)�񺂭�S���8��٩��R�y�Is7�[K���\��"���7���P��Cc��6䶍ᮧNz�T���åy0Kt�f��Y��aJ7m
gC���{�W��n��q˭$-֑rh��H��f�3ִ�ġG��Q�눼M��]��ۣ�j���I���O��(F��a%���v�=+�7klұ
-�U@f����0C"�v�V-@���oOi���;�v�F����S��m.���L��b�I�9�,�OPu��4U�`���"gF����{%�n�=u�(��cBcM�F�I��[��wC��s��=�]��<�9� �8� ��)��0rM�.��c���5-7���,�v�qq���3��0���z���M4����7[���"A�vm=�x��{Z��Լ�Qt�-���n���7O	�sz�z�gt�о�>�2��)v.5Qd���ұ�p@��Z1uM5�G��iP���JT��A،ӄ�vtI=Aݵ���ú�W���4�g���v쎔��v�-ov2�a-���m�G/n-�Gm�nI���
��xn���M���%��3C�ha��Sh�8-iG$Ԫd�Z��@ـkmV��`B$]+j˂2Ļh$�Uz��8ל@�����r�c�[c�]s�QwAWH�����������\w20�jGEv�	X�I��ZV���ك�R�j=�u��Ρ��'�K ]%m�⌙�;	�j��`%�P^E�����v{AR��������tĩ�[�m��M�5j��+��zz�F�u��7zc��w;������œ.��-��-F�58)6�/[u���Y������X���lc�٤M
��rt)dX�
8�޹om��K�����l�g�l0�Y�j��*܃+�ٳ7c�$u9�q5s��M���3�z�[cq�;XQ��Un�g�͊�����қL�����E�p���R�v�Y����q<���=�q��E1�vȜnC�Ӑ�k�\\ݰ�M#˥p��G����	˭��e��G����n��9��2[Fƚ�!A��&�q��6������)�.�K�nz�z�`]�Gtp�����hv��9��k��6B��Q�#��pQ�<s�t].KE�T��=����v�hRrݴ�RZ�U����b�ve�[V���Ys���ASv�q=ne�㦖����#X���J۔��Ay�O���k���s�x��ll9�����ȬZ]
�a�2ka��w,a�r�d�ݮ�^�<	8�S�L�@]e�V%�X7����t.ys׋���GM����ܖ����5�u�c� Nɮ�x+�ێ)����`�r�YPMXL���Z�[S�^mك�6M�ق<܎�t����T����vR�%(j��j*����5�rjg��j�B#��bЖ;puq��xȇ[�tp�a��� 6����!S��t0��CHM�T��#�-���(�8*FQ����Mfr����8��u,3(а���l`�J�s�tм^�#��nۄ�� �S�%�gu����Uwܕ�ؓ�&S�z5�n��n;Ñ��]TGq�ݲ�4�l3�D��j��J�4r���(�OI0)3��2A!"��+��%�+R*d�=
�<f�B�$(�/���Q�eY��^I���}�aPPB!z����Q��QT��Ud�3����ʼ����J$�P!K�&��CZ5rm��"BCʤ������yJ��$S��˞̮�z�xхA,++���g�l�e^E��z7�䒩�$j{[ji��&L�T\l��>ӊLCr�y6��݄�it��h!hv	n&��t�z=�����WX���$���z�2x����h��r��h��T���5�x�wֳ�毵ھ��d�{�Z�p`���O��lv����r��:xT�Mt��T�n������4B藲Os䅯��(��͞�!��#q��F�Ħ�S�Io2~X����n���R\`[��W<v%ׇn �5�Hi�v �3�l��W+Σ�2W����m��cu�N$���yf]W�3�6�E���0n��Tt������t��B����.^L��$E\���\�	R�iu�FH�ޫ��D��G]p�Va/n���n_y�#��+q�F����F�xtkگb�Du�l���-夬��;5����� u�-�?��G��1��{f���;�(f�2x��S�7s�뗮L����b�B��u�8qlW=[e16�-X^%�[��v�2��,�9���属$�#z0[oxxg�*�t������'�"���z=O^�;;������j�j�P�ð=��Ϧ˳n��ge  ���,[]�����h���O9�%�R��#-�G�z�u�X�,@�S]�i�[/��E;K:�7���:l�%ۇWF��A��%�ly�oa䅳mF���^��]+%3P����C1gmj�삔Av��b ���\c�����:�DWn�k�[��Jٚ-�h諨�n�2��`��Ę%t���n�o6�-�1nx7G)�PF핹�DI�Hb$,�`�ģ�uV"�;�m�p�q����̺���79��d۶���2C5�I7e! Ք�=nr!��H&ϭf����2e���:K+�`��bX�]�B�3Y�U�fD7x��� C����Ĳ�c7d�f�;Bvz�AF��ma�-M]e	H���K�.u�*����ha�^�O��V���I�����sX��� �6c	4�%x&��B�AДS��76N�r�L���us:y.�Gp�}�O1SL�Tʍv�`�E�V8'(��M�y���S��s��ooh���{{�0��n�H˗�;Q��am��l���W]�S��gB��2j�fíFڦ�gQ��쎰�6ι�֩CdԹ���GEՋD�ָ��̌a�-�gr���&m��h)�9b�ͭ6d�Fõf!��.6ƍgN"�Ɨm�;��Ӵ�#�M�fq���wm�Ե��Gjv֜�����~���r}���*��G�s��.�$m��c2BI��Uh���ߟ���XL��!�r��r��֮�����^��~'�+���dk��pLz"��6I6{B"<J���o��{Ƕ9P����jһ�(T�O��JPD��T�D�����r�^{��$�}~�4I�Ok��$�$(�������w~�|go�5D��b�H�Γ$}����vT��{��$C/:\��|+޲��,Z�f)�X��}ێC���}|��Q&����]�E$�y1�$$�9���\�*����s�z��{��*Ms���7!0ZF7`�e�+F۶�&��	��"�V�V����|���c��l��`Bk��6@?��n����Z:���֞�U$��t�>�OZ@�&R�=�t�#�#�ݣ���ɾqTQx9�h�7\ToŮ���)M�غ�ݣ#��*vڊ���^�5����ז����x�W	&��T79�d�;=�UB�E#��3�r�)A^��YAQ�(IF�<���$�3=���&��ސ��H��@#�Γ��D����P�H#C�V�V�
������YX�]d �Mvr�L�I&�=�BI&���=�؄�{�&�m�d� �!D�(��Q;��\s�����Q&��t�I4w�d�����q���o�s����]f�:f�YB���Wcjp�\/�s`�:�1��4v~|�~զI��|5~�H:$v�B$�/q�����Ǯ��[n��$w{c��W�!dU��R�g�-�A7G	�Oq��{:d�h�Y��!$�v��rI�6��z�r�����D�b�&#% b}1)M؍��>� 8��ܢI8<����ݰ��6�"E2su[�ɇu+�l��)©���n���<�|p������bu��s��^�4� |nU�3A��;����H��lI����b\t�l�7p����R�����Dk���Mh����J$��:Y~��v)�$���*IJ��%ihP�>'��[��ksU!�^GΔ
���}'I>$����� �3ΐ�;��_L�X}�;f63Y�[�E�=����>��v���]d�t�ڥvmt��HM�0^k�&�OoJP ���׶o���W�{d��	��uʨH^�ehUڤ�R�_c�ɢem�y��ub�&6��5D�Mz�rh�����$��7����9�lO��V�B�!R�&���$��6I&��� �38�f%�q'�כ�P�I�t�~�$�D��RW%~���\�����w'�I�Q��P� W�ʓ$Tw���l9R�޳8�u��)h�p9��u����nŪ���k^՝F�)�X��	�g��=��}���Qy��3ω5FZ��B~�+D���
�B��k�Ο�ɢO��\�����=��ē]kr�$�5���$�~9��!��R���^�� �>��C5Z�c�UjZŖ��t��Xl����O���RH�B�g��3�$�ksU  ;�$'޿%�ɟ5��L��\�lMfj��4 0���@�*��:1	{��|go(h�MfyRd�M�l��TO\9<��,Ǜ^͛s��h�j�RF)F���d�~'���B&�}W�v�>� �&�5RtI�Fw��Lj�]d*T��gٓ��)�mg��Հ�&���$�N{���&�}��d��7:W����&�j��~�Y8�Q7����G��%T$�O�E pj~�t�Ā;=�T �I;~�\�U�qV����K�v�fTk$�ﶍ�Ǫ�7�trnVTL�5f�u3E���	�����b��{t� o�{�R�����m4�Y�v.K'�똹��b,l'U�$���غ�������Q�\�� ��E�Q5E
�h����P�l�1�{���5�ۭ�%�uݞ�s�]�Qۢ1�[x,�at����XU��7WY�+�2��5��	s�X]LZ�4�M��zy�ɠ��3`�'��a�tfs�5j�E���^ҝ��@�d�e(kj���l,�\����Z<���?~��uF\����h�Nv�bQ ��u�N��&5��I'}�$%�)WV��EZ*J'���BL7]�)J슳�d�k�w}��	'o��B�L���۷è��
 4�R@�Q@�>7��*D�t�(�e�?q�+q����I����U$����bPU��]�j�RF)��t���^9>הI&s�Ģ@5��됐+3ʐ�|#0���4 >���1����*�T�B+�(j�?Q5��M���m���~�$�g�I��LI�t�3��������M��[VهRX�C��*��9à�KUx�1�sV��Wv�����j������{fI�G��)�Hfy�d�4%xe�u@�4s}$�A$�=��T'��>�mXH�k�k�4�������!�r�냖�ā2%���/^Ȭ���zȻ�0*� �p^^ʙ�Y&U��;�f-��"r�^x�Z�� x�s��BI$fy�d���/�qf�o�}�	��]\���6(T {ӹ�H���2I$�d����J
�k�����oĒMQ9��B	$fy��P��v��(�c�/t�5gޕ�`{�C]%8~$�Gf�N�$�>�lT�َ��$�^�}*����5v�A�j�?�?h�v�Cd��*�A6�$���!$�;9�d�O��'���e6�ob�G��H$|B�����2��� �U�H�׫���#����G+��|��Rj1����28I����h�g�ITJ�Ƶ]��!�4'k��|�#J�D����s�a?��U���i�D�hN�I�H���B U	�Ľ�zQ9�_d��ڰ��k�᧾t�D�3��Q:�p��I�/?
ǜ��<&L'��i���Z�-tW	]·�T�-ή������y���`8zJq�G|o�f���и�L��$�u��6�·*V��b�@zrr݋��C��Ě&��S��� �d��$�'{ڙ�sjF�a�C7Γ��A��ڱD����р%3}�� ;dW.�n&��Rd�$��l��D������#l����������k�3�4�+kaq	\h�ukxH�c.X��b��]X�g�������6Q>>Yy��&�$�n�%h�G��R&��wyl	{��֠��&#�]߮"��pP&�( �. �캲We�H��p�Α��Hq �wd���w�HA%L��n�}��t,�) J��J�>�BI$�{�8h�MK}�#��w���Ā~=��>� I���	���Jʥd_+}{;�����R����I��v�	$���K~�4���ļI�)<�X�3�ٜ�V�����6t�	����l��L�(���f�{&	�n:q�57Q���B���2	� �TL�S�=��N$�Mf���>/bw(�$��ޒ|H���!�H���4H���+]]7D��LI)�JI^�h���<O���g�fܜ��/4uf�ѫ�������TK���۞�D�$f�S 	Cێ�&�t]�OOgw�Ztw�с(��>��J���z��WH]���]?�$�^�dw���[����BI4I��ݪJ$=��:$��>�=��E��O�4�غ��Y
�(e�8�k݊�̚$
8����*m��zvI���?Q5��I�'��:�B�ͥrQ�fCd�se�h}~�$��������HI�=������B�y ��Ĭ�JVU+ ��I��c�ɢ@��r�m-ŀy��/٩�(�3�� �����'i�����2k����了;��*+*����מ�xI�ƙ�+�z�E���]�۲���ed#gv4yc�t'e�9G���|�s2V�Z4��#.�	�xa��%�xx��K����^��v:���v�.�8�vm�w m�zƵ����lsAɇ�8u��N�ؕ�t�����6bű����K�Q�����C�Og#=��w^.��{]sD����*�9�b�&�9���g>��vz�,릥Q�/[����
��u=�/l���Y�U��3���q���8���XN�\�D�g��@��dn�7��o�������+|H�Ύ h���H2I'��um�w���OyJ��43u�и ��V ( b��j�4M]J���}?h��j��I=��!�h2����b�	���W����O�\�O�@$��[ J'V��a�8x��&�	$�����?�la?��Hп��U�=x8R[f�� >�(��)"����	"���w�V�5D݂�a��׌/�4�� �WGCA�����{�#�?=���u,�Uq�'/Q$7��$Fwl�B $��S��oo���(";SK�h]�d�vМ�F���TK����q��f��>�|�O�Վ����|�:2&gk�B$����	�e?{r�z�� $���P����R�
�!#��)�L��W�zc�xT��mWgV����]�]�=�;��>�bp��WYg�@{����1b��n\,���
Q뜚�X�J�xD@����O�4I'=�S�A����vgs)�d� >��`�)F.�*D�F�|��8��Y�[F�أ�ZI$љ���DDgsTD�8lB�H�KD	�u���)� �x��}��%�fyҠ����n|H���	s�[HՑVB�JH��8I�<�OX��-h{�CI;�d�I���=��!�?�:L��_~���)X��A*Ƚ����k��fs��|8���BԲ�ш����~��?
��ݤ`͑��$�H��c��D��g� ,S.�V:>�����'�ڧО��a^Q%x��*"#rs�i��K��$�Noj��D���I� nRnx_�eX��2����+�V¤$w���nHo[���u��<���FNzo����i����x�+�"���sӨ���P�zoxe>ȏr���/9�-
i�[[�e.ݫtF]Q�gq�Λ����B롗�A�I�;F,){�2nF%7�c�3o"���ޮ�I^��9�"4
u�^�ԝ���]b�ޠ.�eo�ӽè�1��\���,nq�y��v�ԯ-�g�^*.�3��ؤ��y��i);�7*�:�f�ssE���+.����Y������\gj�N�񾓞�bۻ�ATw-��ߏj؞g=awf	C
۬��ru+;rt�[;�-�%� ][3Hޞ���ܲ/�W �攮妖�b�u����5s�Q��z�<Q����e��:�0�
�j�rr�;�)fa <��T�q�R����O���� o�\\-56�n�7��V��;�w��L����*�
�5v�̶`��s)��`����ώ
0m�X�Ku��l���.��ᥝ���s���%ʞ��J���^]3�������+���K0 �2
Klϟ�Q3뙝���Q��0Vl���XU����"w�3�5<�]����e���Y�T�����P���F��80B8���F��;>3K,>@5a�,u�'��l�_PΙy1m�z7��,���)B�͂����/;U�ݭ��rT���,�(q}�>��q\�I��h NZ��]|��'�t��P��%/&4��~x�7�	�?��ű~.ދȺ�t��y/k�/w��#�=]9]"V�FÝ(ZL���r�rj�2g���1SOؗ{d����ױҮ9�%� Iu�1NC<<�{ގ�%w��ǟ�#>1!�3�#ZeR$FN�.��������*�d�l]��B�{�xO�׹�*d�bbyyX���>��$<�L�X��N�ʭg[P�{3�ď�
����]+��fC#�n�Y�B(a��{������@Ds��L& D�K��팓s��]r�z�`P���O9��X{�H��G��_W<�9$���
pް�C\U$�4HOt��=��#ʽ�ǒ����.���(����r<�5<j^N������ɝ�4�^�'����|�Oz���Ҋ�ۓ*�R�c��
,<��>%(�:�20�E(��yyA�3b�ͼbO=/��S<\��a�Sɫ=�IT���{Ǳ9�ɽ/���Y8'��B�j�"�I�ɐ�y�0�{��*���)-�����2,2�u!��T���kM���~o'�[gϞ1����C"_i�{�ޭ�Fk�<P ����$��*N�]�1��ncJ�،���I�MQ�^��]!v�C�c��$�D����M�_�lzw�4s}�BI$d�HD���{���|��螏�4�5�ԣk1�)),�RUM\�0,q0L�1�n�*�??��#f�-iR� W"~$�]9Sd���l��m��:�;_{F<&�|� �$zs�ɺ��4$�H����J�HzD��k'�&I$�}��*��i��w��P�c�|���ʣ]9��&{\�OĚ%�{/C,R��dY�h�C��'�'�I���P�K���+�V ޝW��8�BMQ4�T�4I����wqN�5�.�7���P|#bZ�چ�xr���.��!D��6F��ݝع������+�۷gHW+�`0R���H�6����
1?l�43�:L�Pz�*��1O�^�*�$���U��`xN1�	Q���
�$��ؤ+�t!�R���($n���y�䪫��f�Gk�>�ڶ�,[��k6f�ϯ���hՋI��c��$�;��*� ���(����<�1��uD��4}��!5 �]HՑa]�J�L��D�}^Y}<�S;�D�S��E�@39��$�I����W\��%ݚ�jR�Mה�� �_]݉zl�Bj�4H��g�$���=3��n�yǞR�$�Owl��D������C9���Ȑm|5�Χ1p�]E�L�N/G*	&���rUI42yҳZ��ٔ��h�fF"^:�஭X?
��g[��[5S�vko(��}���$�G�{nUB	5�ʐG�Vׁ�2��Ǜ`���`��F��[a��g��	��3�\U�s�2��������V�Ѩ�i�/�άf� ި#U�l��rPD"Dt$�cU*h�2ƭ��wYf[��¸��[�㣎qv��p�qۭ�m2��y���n�6\��:��G]�5-�����z�ޡ9	��p�M�51�K4�tw8A�Q����]�� �f
�2�%�h�BlC(�J��X,4t[�`U��ӑzjȷk���{>��Z�J�[Vl�a���sB�s�I�n/R*mw'��t,l����.�q��� y���h u~���P�Iý��~$��t�6ׯr/�����3���	#{nBj��^��I"�B��YL�}�υZ+�0�nT&�4I����$2y�Q&�{j8<B�܄ʃV�j�XDZ�&�$�&�ySd� /h�=�=ޮY��=2�4I={�rh���I�M�|��!}wi�2`43�C�3���BSɀ���I�>�l����4���H{�T����$�_	(ן:uL�I3=���������J$
��I�I$��{d�k�^��❀9z�J�|/p玑�+T�������3$ar���\O��(ի�Y�Fnz8I�5R :$�=�BElNi����B 5Cs]&I���@��h b�/t��Y���ў�19y��iX;�:� p\;WVo'�K�j�x-��\��!�tw%�s�)����%�KOq��ԡ�I&��&I$�g�I��5�s�/^,�)p��mI"�\j�6@?Q>��>�N�u��̋+�ӫfw�q5ݪ����#��lJ�.@�شA�J	�w���C;��А)�T�$��3wd 	G/��t1�\��P�GI�J�|N�����i(�ْB~$�=���P��|5�D�����Gsw!�I��m�yo;�'x��e g�Q��M,��F�b�z���;�[�x�%⼹��?���＀�I6�V�T�&gc��Mk/�ے�%R�w�n���y��D�$�v�b��Q�V��{��T[3�P�{�'*�Mh�f�r� ���m�A���B�uڻ�:��򰑷@��i1O�^�*D�'O�g�$�/)��MX�'�y.̣r���jGm���M��n9�ՁsY쫾��_
�6U�΅9�-[�w�%2�|��/~瓠��<u/.�A|;��7�`~$w~�*I~�b��\-X$�B(`\�-C���/�I�O6'�I5���%I?W�뫂�����$,m�$��I�&�A��F��M�P�OG�J�4O�j�����Wp�~�����I^̒h�Ѻ���0=�n���v����;af�+�%��&��i:�L���ym��U{�I��j�׫�<}iE}f�<&��	$�O��b��I&�w]X鞬�d���{�J�O���ەP�J�2*�"I���Ú�D�H�A��-��<lmv�Q'��n��Q\?D`�]]��!	j	V�x�t�h���$�M_j,���5<$r��rj�5���E�
4t�Ťh�(���H�6�b��IGْ� �Ẫ�I�c�����G�1�tưUM�r�.'oK��!_6]z�����9m��Y$f�u�r�|N��^���v+��Ϲ��H�w��UBC�V	$P�Q�s���M����W��~o/��$���I'ǵղ@���F�BB�$�p.L$ eI��)Q��� �V:	f맬��0�+�W���~��Hj�g2E 4N�j�_"�$�g�ID��~�ޮ��E^�ܨ@k���=w�j��f�2Uvd��j�{�����I�;��� =����D�6<Ֆ�'j,�i����pdU�
D�k�'�ã�����>��I�'y�k��k&�V��0v��I�Mg�J��T<]rA�`�*J'��+���oIB�c��IR[�pdĈ�Iy�]ڒI��wF�7����C$�9ղH��<�a$(�(��Q:}���s'P���|:*�H罒BN_{nT==O�缯�~`瑡Y"e,`_9�Co���^�����QD�
uk3�ݮ�J`e�CN��#d����{^��g��d'�O.��\�y�:̢/�\���+ г[��cYIms�@WU��g��-�cv�r�c��R�4��qp�®ى�5��qiثB�8�6��gp�6F<�#��.k;��LB;Yv"T�7�Ʈa��T�/�hU��֝xS�.�u�mr��풣�f�Ů��Qu�tm�F].A��mL���q4��U�sXݴr8Y'�6�&����HJ�l,BJ�̷�TV��ً�~�~'��3�j|�_ac�H�I=ۍ�D�~��m�H�~u��+��u��IێBeA��F��M�Pʢl�%�z��!�Y�������&v�BI��mϡ�F��ϳ�]��U�&�:Tz�ڣY���$�<}�)BHk�'�^���r�?7�� N_{nBi��g(�$�_	�GCS~�<X͍f�$�%��BI4I��m�I���	:c���r�C'c˻�x��5j��T���:('�H���=QN��	��Y�$�I�Oǯ��Z��$���Vd;�v�;ҦU�u*�Ǎll4��l�˾�/i�v�#�hP�js6z�Vl�j���G�+�B�Pw9��I'N�e(I$��V��X��|�v�������_vܨi`�,����ԣ�N�$����׾#ۛ��A�'�b��p�[��9p�g��fM���Y�v���^�u�2�=�}�p��s=
td{�_̻~��T&��D����rQ$��uU�@j�חo�O'�L�9^ѱwj��FM��U(h�D�v����&�@����q ={�� �}���	tr��Q_Y����̔pO<!��Ǵ0�O�v�	&�>��D�h�=��^���Xߨ�F�ӭ�u`�,I6�{Ū�~$�3=�}��4I���ܔI$�]I����{d��_�Uܶ�Β��7l�sO������wJq j�f���C�P%	�@}��a\��CpЪ�h�D��g�HN3��Rų/�됃D��=z�H�υX	Z��~���>n,�qi��v|o:�Q&�>��E���{d�I"�fV�{�jAp�8Y@+I%b Y�YVOğ��n�P�$�V�Ⱥ�&�j������a]B������M�}^^��g��b���{@��j#Xu�[#	w.����[��:�?}�9��o䐒>V�F�$'��we�]A��F�ݪ&�@%y�Szh���/�M�b�VM��$�MN_{oa�o����>$�z迉?7AQ��B���2|{�#�D��m��v{v�vt]}�΋�MN{�%}$�����rEc�zz�s"j
?���tR!Q6�����.p���ا[�8r��3"�>y������-������X�Q$��͉D�$����R^�Z�����:�D��?��bU�9�ʒj��j�ӭ���C��Ò�"k�I'��$$�0����7�:�W��ʼ�kV���A/��Z�F!$�;�>$T���=^��QU�'�D�s`J�F�܄�Z<8Ք�I$"�j�:��Q�Ɋ_Ě'ۺ�$�߻nO�4I�t��]�}�NC=ۘ���waE�vm��U\qMEp��W�q�v�3�e�;a�����j��SՃw���jC�wX�Q�s��3�I%�|�.AYn�^�uv�&�a6g�EĚ&����&���$�tI�HI$��{nB ���L����%��}�;�`�F���^r����mXWx1��;[(���֑�p�|�K���kI�[���̌	��lP�I?��O�O?N������O� ={�%;TA�U�I��o�����ؽ��IrG�=~��$�z��rI43��2I9�u��QĄN%�}P���G*HU���>'���@���t�$�K{��	����\�3�M_v�hg��d��8��A/� ����ՙ3�0��I>3�P�&�#}���I$�=���q�f�g�v�D�;o�؟���VP
�$��Q|�)�D�}ۮC��wMo�/i��I�L��H>�y1��滻���<{۹W�?����p��g3X�nK���1��́ӹ�6���ڗ��<�0fTSic�UOa�;2����$��������T�\5z�n��<��y�<`��ًNF�=�ς�N<�#	��A2���c.\�V[E�b��7R��E=�3",Nҕ��s�U��zF�3��ʺ��S	"����y��Wu��P�S���ݲ^N�+�u��;�*͜pܕz�D�r�|%:U���l���ۊ����(׽�f���>��=��i��IPh5ك.���ѴF��a�2������k\��#U$�,�cLܡ�W�7DH&a���T*�wJ��X�ƶ�L����6�aj��[K�v�b+>̍P���%��;�X�퇸)�΃�E�z�`=X�-�l4��{�����V��s�v���TnE�����R��9`������B�9���پ.�횵k���kr��tS�q���Bth�H�h]�[�D��j&��˽�7�\�ݝMl�Ұ n�uαgs+)X��o4�͜K���6�o1g\cf��dv���4뀨���:��.���B��oh{m�L"L}ӣ��w^7��U�e3ƕ`�%ww�u��7z����گ+�:������7pH���W�zgÓ���N�Ρu�E�l	��$e���@&Pޘ��� �ɣ,˒Ax�R	E�kh���
�4�R^5M%��hm8o[N��YF�Ň�-���ӳ��ն�bڈNc`T#�l��|~=��G�o�����w�ʓ����g�֣^�Ċ����d'�^�A*��k�D��)+��w�U���6.���U��ʫ�<���X�g�Y4aL�J��Bm0ZǙϓ*�˶�U���a�**g�2z�:zY���hW4��.��3<浺��y�:�+���<��'���')��O�EGĭ�)�<�mp�U��+Ǚ���m�Oz����z@S6�9g��y{���ǽ�O�􏶴�z�����kc�yzb�y��z^���OD�(/(��n\��mxx3�^�xL(�d�r�������B

:�B{�y|�!��S�b�я@^�aG��U��)ޡ�^�{B!�D_!�>�JP���P(
r��fs�;ϱ���/ Ԋ���\d��2���%�n���Үx�&S7#�ϙA̦}�2Om��疳�N^TW��M����������	ԁ��䰺�D�#��￶�?+V���Y�g5Ιf�*&��m�a͕���O�GQb�6�};�e"kX�vX�"����܆��n���v��"d7n�s3D������pg0�n����b.�����_Q�ü����醢k;e�ʙ��f�3�.u�¬0qq��oGE��������{-Nn����0�y���+�������.2-�uY�K��S�s�����)��B�����,Z�@�(knf�i�a��.�y���t�]���wF��獶��Q[�x�z��l×�����-�3�l��6ag�GG�s�I{
xG��= �������A�=�{p66MܾA��0�E��1����f$�����b�]Eʻ���b��S:�u5���2:�6ŉXYT]((mm��xs���[���N��P��;iyð�lrKŃ��j�xT�ɘ�ol�Ԅ�妖YΤ)\�K��9
�ֆ�H�h�ڈCjLjx�������T�ͣ�ǉ5�Yf����S�̖k�0�n,�c{=�/NF�'�0�U��4���Gc�7+ɱF#��ַ6^z�{r��PQC�W�>6L]Dͬp��9��粼( A��i��h�*�:Sk3u�0���Թ!ab���к��n{k+C^�<���.�ܚq@���^�`�F���܁i�k^C��+�en�lŸ�I4���ˈ�.1��3��7����m�i{��X��=�m+�{U�ĒO�چ��X�����W9-Ìc$oav ��ӎd��{e={Og9x�z�&���#l�qH�X��A��:0�`�b2�Ku�6���Å�i� =[�Ԯ�=�XK4�gE*�Zl٧
P�l�"�,�Y�#�+����[B�5�ب��X�J��i)�n��٬n�z�yz�ƞ���6@w=�^Wlt�;��t�����jV�í��6g[Bg �([lHE����{K;"��d9:.�6���ֵ�:�m�[����,[�o[�J�+X�!O����~kv1��˗jZ��y�h��r�ۉ��	d��٣�°R+,])W��5ȻC�N��=��݆\�j�[2FX0b����[������hFdtXe�� ����|�ǎ�%���� 5�ndfq����-=�m�ֻMqXo��_��\��%V���^f~�$�9�3=C*�Hw��ݒ{�f�}s�Uݙ�5�k�ˎ)#�u�d���*˾���.�#!��J�3P��4��{���nA0^�
���'��n� T=�;<fI���!eFi
��J_{�ӦM�됒@{8�W��: ���I�$�T}��*M�#PH�Bc�.�F����[;�nfp�@�kf*tɢOğw�ID��Mj��ev�����?P��@1�~QAK�U��T&�4Nm�%\���޺L�I;��!�'ڽ�C^�$^o߿�l�+6���Q�)���&�&��lO'��]�ҵ�3Ggￇ��5�vUOO�f�t�$�N��I ��a����{/R�-c�����&���%Bg��꺻JɻT!��~��}Q�9<jgy��(�lu¥���5y�_m�,b�.��aH�/�����*g �wY�|k}=��3�hOl�u�m�����`��?�$�?���I�I�j�a�B	2���(�yu/Q)кۼ���.�"�>�~���ܹ��%1=�����Xǘ�"xDA�쒡 =��d&��MN��*$��׺?���渢M��*	'5{�I�kۊ�y�W�ܺ0�c�V礨K@/�I
HY��޹��f�ɣ�����.�@:�=$�����T �^�T��ǌw��ø�C ՚����6U��[�]�Lx���tҥ����f8�����!i/�W��шI'v�'�p�h�T=��?���^=p9�6O�{��W����i!�|�$��o�W	�X�P�$����H��&�qZ;�5�[��&����H�v�BW�.$�^�T�I�g�Xvϕ$G:�c�*q�W>Nͱ	̭�W�Y�w=���|;�-��8��]-��C5&j�%�j)��NJ��� ;���(�TI�����B	$g�]&I��9w}E+$]�FC���l��jc�I8q�W ���BI������v6�t��<:�5�2�&����@]�����H�$	؛;W�&����d��ې��'�d�I��c4*�rW�.��Ҟػu�b��uL���Ź���ږ0���98rPI.�ƴ�B�~5��'碆�5D��T�$��>��u-a���s��Z� ����I��@�F�������$�D�����g�$�x�][��D�=��! @��.-�ͽ>��}	��8q�j�+V�*ʤOĚ'���&�4M�������=D�>�V�$��n�P�'�Uj�*�@%y�V=h}�u��I4ו6@��n~$���_�,�ݏ�6Q��u>��5}m#iS���؏j�:�J�M�C��*,���.�d�AfR���1Vt!H���6�uSM���	��"~���d����7��"��2Q�=�Bh�D���)E�@�.�W��W㫉4�GV� ��l`BF{.}����a"���"�H`�nu$�&�G�\g[���P1�m��Jۊ��V����q�A*�R�1SZ�|�$�;uʄ�~$����%�<>�����F7V�D�3vHM;�_*K䅟�@8�u�'��t&/�b $�{vHH��*Iwm����o��v���B-�I<B(�_\P�>��$�t����<���ƺ��V�$�Nol`J$a�eϡ!g�q�j�+V�*�����ʫ/�@Y��@ ����$����{q�'��x�qϡ5(���Tm"Mڡ�v�D��U:gO�
���MOg����'��m�'� �:
�+��rvT��
g^dƊ�9�ɳe�0y��b�? =,�D�֙��F.ww��"5	+Av�˦�7��BCf��7#)D-E]�?���4	��A�e����wJ=J[;=������,��(�i�H������B��$��e�4�wo�v��m� a ��A�˯.�!���1+�{J���4e�7��/A��F�{�t��u<���sN{tݱ�� v�ĵ�c�to78��b�n����I�!uqj���{\�\�50�tƱE�L,bJ�up�0.�]]�1F,Ji�r�X��ъݕݭ��n��@�wi���! vϔ4I�M��N�'���*���l�f�P��v���?;D���"������RTO����}����lx��<}�lMg�Rd�s��dӻ�s��d_�x��?|Og[��kwU:d�'�$uM�m�y��jI$���uaq�C]�eI��$�:�F���Z�@O�5�\�uh�+vR��$����I�$�G��7��u�3֣�2uʄ�A��q�j�+V�J�W9���I�}ۭ�� �A�^���$�F�L�I=��>�\�Jz'�O%�2Ǵn�Bʮ�m�e[�7u Qp�į1m�
��һK�oQDZD�j�>��9$�BI'õU��$��g�@Wss�e�#e��\��uU���7G�	v�y��̺6D�s����~S���b�R.2�T��q�^"�П�c1ms�E�p������:�X� �1��i��ݚ�&��=Y���I�M{U���'��U�I'�����U4N������"5�y	V�4%�Wb�����ê$	��!?I�ҧ��v�̝�ĒO��պ$�#��r�/����?��3�莝^�tI�|'�4@$��� Q��m�Q�$�}έ�$j�'�v�F��Ⅿt��j������+8k��b6Px���$����A$a���#Q�������~Ͳ;Fc]GLݯ4g��f-��SUR��`�[�����XS7Lտ7�¯|�$�ݺ��B�O�}��.��䖣���tI9۲C(ݢ���*�eg�E �3/��͚����"1����D����4I#��tP�/�ː������7C�(.�"��wْT&�?�}�BH�/�!J��Z�Ur�g9A6-=���NأJ�6e����,��Q�Z�W4�^��9�he�8ƶ����
�$$�����0�~ەP��4%�Wb��p��u�� ��nx�e��ğ�ő�MQ x�� L>�WD����Kr+ 5�B~V���Tօ��HO�I:7U:D�y�u�,��$��I(��{nB �#�	��0�i�gy��f#��@�����>on�.EפP�2��͞�՛8�}��ׁ�%f���~��z1	O�mω$�>�V�(��G�a��v��l@�ǁ�6U"�$"�lNt����3�Z�_��I�x�m�H�պ��<���8yz�o��P�{l -"J�A�_g�E	&���Ua�&��	Ү�����%{�I�I��mʄ k�պ$���4��"��0{�ga�@����(I4I�a�MD�u,�]����vNM�{u�r���zLP��8�n�2(e����6�&W/w�qxCKlq���v_y0�Y� 	V_T�K��w11$��uwwhPp�z:h�h���ʨ}C2�������RUh��V$�g�1�x��)�����ǥ��%DP�m����r	��	؝Ґ�N�N#0�8��������Ǟ���6w'	Fꦉ$�}�� ��^מ�s7���=���j�VU��0��K�h�[TX��}ҁ#"$��ٵN@5\{][�@?��BY��Ƹ��*��mO�!��6U"�$"��4I {;\�I$�K����L� �O�w][��I>�쐙]gq
UiU��=m�0z��}���j���S�I�&okr� �b���ٞ�x겼��i���a���n�#%Od��I��N:�'[9�s��*��$w7c|I'��Lc�.f�]��nϔ*���ÓD1X���s��D�.R��ɹ�7�ǔ�샣kU{,�;����b�Nk��4lD �Y�Tf3�z� ]7}�r��uO
m��J��d6��:^�1U&�4�C%D�2�V��۩"��Ѽ�a�G!���vvڎNϫ�xQN�O'=pd��
Mɴ=<��5�<�h8�]cƏxiD@7>;kp����[�����2����Z��h���ȗF����h�<�j��1����9]"��kXt�i��U�q�iq�F4�lyZ=j�f�C']-�NK2eKfp9�~��m���7fѡ߫�1ӫ gn�P�I#��NQ5�����/��E�$�w{d����Q�����ID����s����y�;KT��$�I���$���I=��>�$��.�rox�(�<U���$,%��>/��	�I#��>pDխ[�r�G<Vz/Q f�$�M��R�"xo�6U"RHGG�wnZ��6I%f�P�h����)*��qQu���)�Dx�޺7c�"$JQ��$yI)�I�'|qS�Qb�������:y�HI�@���s�D������_����|�1�`�g�����vR^烃���G�\T՘s\+�^|�lyb�[�[�λ;$��I�dpNx��%�O�Ů^9������4I'{�1+�h�D��tl]����Dm��s�i��4W�ػi���ɥР�y�u	[�����k8�yj� P��������z잤MdЕ�L�J��xx(|�?ЀI'�{�I'?T_�I�M�\��H�[�#u�� ��>�GOt�p�$�Ӫ�tI�KU�W��>YX��zj�$�� ��GI5Ⲭ�aX�K�^\�ve�V�����m�I�8����uo�M;۬&�XuH6��d�=�)P���n��T�V�nQ�9��I�}��T>�a�A~°�~���RU��tH�=�}
5t��0�C�����p���>��f�2�n��ć;O^���4R!#�s��B�D)@�~�O��O2�N��J�*iUEM��r;Qe�MF�j4�;�sҶi�J�|�M��q��ͯi��iSQ�W�ek��SQ��MSG�y���2�)�e]玩�1C�U�Z)�4�=�k�j������UN��=��M5mi�5MSE&ST�K��]��1X�b��TҪ���cM-��R���=���v�,����e�f�T�+9nG5[��:�Qq��i:h���#e����
�STTJ��������*j�M�2 ���sڏ��㙜;鹢�a
���"oe-A�wp1�x���Yu��u$8oB9�f��.�F�jΫQn�Z��6ov��-�����c��u�7�L\��nr�0J��I��[�[����,�ɰ��� wnG��j ��j���l��������]K8���9+��� �0�hMLg��J�b�8�^r�'#h�[�~�+\EiL��l�u�vs�Ɗ���F�lIi2�ʋs��|�3J˺ȓy�54+�^]�q��ܻd�+8nVG��n欢�N�"u�ڇ����!ZK�ׁ���W���ee?�}L�>{u��o"�Jй����-��|�v���7�����h�4^�w3;��Zi|2nI�]��'��zF�﫷N`F]�ާΧ��m�����5Ðl��f��Ý�sV.�X��^nXq���P���{ݬ�� )u�q-��Eȯ2H(vU����k��6'FkV�\�L�春��a��U�<h��' p_[KiZ�}T�8�9݊Y��ٲ��][\7@q�՝+e&�s�7������l�N����(]ѕ'�^�[Xeb;Wv�d]�����o�I���)�R�r���6��J��tpJ�c�pnX;#����2^�� �o��}*��B�_X��v�y�ul��/���r��6�N��o"�lu�S�!�3b#�sz��]�U4�)��{dRe�ӮՆ3/3:m��\޸�{�Y�-�>4�6�l��|
S���ULޚ	؇�	<y��y!$�m�`3Ů{�@ǽ�*>��y�t���2ϴ�y�g�jS���H�Њ�P:	$'=�Dxuj��C��N^�*wJ���/H��H>�ه#AU\L<��jr7ɚ�Q\�����-"�� ��<��a^Ex��Zo.��rfG{oQ!(ffL!�%����M2�W�%��IQl��v���W��%�ɄU�^2��n�;6]H���i��O�8Z���T��mvu�\�9�T*hŷD�K3�6Չ�s���9�7+V��mri՛�i�}��O����cFl$�/[C��&rC��)�k;�ɍ��ٗ���BR�ɓ"���d�릒����Pv�96��2\���/1��	����ϛ��Z�>�E5M(�h�=��ma��STҍF5L�o�1���4g=+��x����4�Q����3��;�w�n���Me��.�Tщ��#k(�e4��Ҍ�s�ΚZj4�4�4��*�{�FZ���]μ����f�԰�zLT�4\��#k�4ST�\����x�V0��Me�)��wkC5MS
j�Q���w�4����ޮw�3�mq��C)�h�u��Xb�t�1S���EC��1���4�SJ��V��ej��G�'?�;%��6C%ZD�����ک�}�ï�����8g=h�\7=M���_���Rb���i[Q���9<�MUD��U�s��-�b�T�1ST�)�d�}��Q����I��9���jTP��#�>���me��(�a֩�߹�4i3MS�z7d�F!J�I�'�D/�)j�ZU4���Sݑ�������4=^��Em*t�iS�e4���9�i[Q��(�d�}��-wQ*j:b�����=V5a������i4STʻ�j��F(r���E5�hh�w��4֘i�j��0��j�;�s(�V�MST�I��4gX�Of��խ�me������5M**�9�4�j*iJ"��:L�V��ezf�T�+9nG&�ԅUcƖ��M���l�u˾o�ZV��%MF�f���zLZj�&*j�CE5L�\��h�Zf��j�Q��&M������z�U��7���3��s�����b��Ύ4�	�=��*����)9�nZ�z���eK��9�]�/]�ީ��,���fL�BIym����5L)�g��cMf���/���x�ÕJX���5L����4�4�Q�EEM��r;��T�N����~��U��]{e4���z�t��Q��tҦ��^�w�e��SQ��MS��u�^F�m�3x������}��U��u�n؛8Śh�#�z퓴�(�A#s�Z���
L�������K����Q�����m+j5��0��5L��w�e�iF�F�STѹ�g#k(�b�g��I:���Ң���1���EM)J*iS�e2���(��4Ҧ;��eUJ�1$�1Y���N�15���o-*j�D��_��g��/iq�ǻ�i[Q��(�f����kM(�kI�5M��r6��Ʃ�aMST�̎C��dW��g޳�>�Os$ �1
p;4�4�Q��w�e�il**iF�G'����4���iS�SJ��kP��2���v���Y��J�I�J���s��Q����LT�:�r�6��M�2��}��ʪ�2�j٦�g���M]��W��a��טSTҍFLw[ɡ�kL(j���e5M��.���:j���TҥP���i��k��2�U=(Ҟ��T�~���D�O�v&޽�~O�ٶR�KL�飳�����Ҧ��T��k��-�b�T�/���f���y�3ɢ��U㷫F�4�MST����r�6��Ʃ�aMSTT���ƚV�~B��3���QX$T�&"��m���5P��@}z���PxSv�wS�&�ڜ�s.�:�]Wj}Z5N�S� ��:��5%J�0����QSe <;nΎ��3���N�!��j�ͳ�v�a�v��ia���z�mˎ�)bQ㍰<
]�e'��=���g���s��=<�fɩ
��	�c�Z�Ѯ7kQ ]B�-���Z��뮖��s�ԒS�=��\�X�ޛ�\]p\�V�u!�'ݶX�</c8�i�aî.�˳Q�07%GsZO#����6j񁕍�]jeti�I�5��9
�
�<��]�`Q�e_�ؾ�����s��ZiF�J�*h��3��ZT�ҧC)�L���3����(�i���~�iSQ���F֢T�t���tÕ�^F�cE5L����9O�c	�4�Y���~��Mi����aMS���7��g#���9W�d�YkL)�j�(e5Mr�˱���j1[���EC��1���SQSJ���y�{k�D>{^�Ͻd_�"d� �Lb�zi[4�]���4�V�%MQQ*g��b�V�z��e&�j��c�������~�7|ֻ�#y��m�5MS9\��ma��-�j�ST���ƚ4�5GM�c1R�0�>��!��w�ϙ�����jc��m/TTҪ��._�����v�iS��ҦW9�gM-3N�T�N�T�*���s(�])�z�Yj=�T�~��{����I������:l�E5m(�{Zŵ��MST0�����s��0հ���kJ��J5:z�뱵��j4�Q�eC��1���������T�f���Q���iS/:�f�����z��1H�U��:e�G
�[��ơ�/�g/��G�����~��<�6�?����:}���l���5U��J3[�1oC��LT�2�E5L�x��h�ZiF�\��x�G�9��Zj�v�����J5Zj���3|�1���T�K8����a�J�V6�š�T�ֽ܆���Ҫ��^� 3�����Y�J"�-������i�b�Q�� �k�R��'&7�3{f�Ug�����������a9��y��:�*NV�}Hw��E�w9�,���2�T�iFW>|�t��4:iS)�J����|���j%MGLT�7[ݾz8�O�+��k���-���V�=*6r�)���i��CE2���M+j4�Q��综�ZaI�j�Q��˾ފ��=}Xb��b��iUC}�1�������*iSQ����[�4ҦQ/ϝ�cV2�Ͽ�w�|�c�~y��I&����n1��/��e��6!���Yc1��Ww�S���;�ך�(�a���ε�4h����V�B8SW0�>��$1؏�ϏOg{9h**iQQSG'����4�������u���^j4�.��M-3C��2�M*j��;��j�Q��1ST�a��/�N�u'����'�n�OJ�̒�ٖ��`hۂ9*��f1�z�
�uѴ��+|�~����{9UX�QMu���mxa����)�j��{x4֚�
j���j4R�{�ckV�b�=��CfY��il*���4����)EM*t�S7����f�Tʬ����J���-3C��Oj�6�ҍYQ*kַ=�g�Im�߽�|b�T�1ST�M�3����j�Q�ҍF��o9Xa��j�Rj���g������:��U�h��5M|͎��V#uJ�5�-:j��{�=5��TTҢ��9���"1����^e������f]���ǵ+FX��{��V��wO<n�ݍ��'��X����B�^>���lS.�7oUG�  xxNv� 8��m����ZiF�0�5��m�6Tl�X�b��Qmh�ϳ���2�z��v[�y�CҍF���r�4���6��˱�4q�;�� Q�8�[�fr.�� ���yܣ��3��IT�c��+Yc{]���0#ڀҌ���1[	�{Z���qO�m#D5[�h����09�s9Jڍ(�iA�����������I�g')�N�B7h�sA�ԗ"�Y챝�\���	�8:�+����v{����:��ƚ4T޵���"�@=��9ݍb!�s��l�`�zi�`F��V.�5m(�1F��g#h���1f9U�Q���b�M���X�a\�l��m9�d��ZPj0 207��9An4q��C��0X��78�z]w}���\
��r�1��r܏Q�������41w=��l���J1��9�2�أD#G1y��^w��Y�޽�yh�4F(�1@g{�^FҶ�J&�J&�;�s�[>���PĬSuJ�6��h�s!��W'�o8�w�1�� ƹ�����h#'��de�#�5;�ejr��ssΧ��:]�g7򺝯9NM\㇙tj���M{��D�B��ح��+��"7����j�Fs�bLVw[�� $y*a�0�|�o#h��4C��Fυb���v�4i�3>�p�[L#JF�O��K�K%f�~{�KlC`k>��A`�؈H{�� ��PDh����a�$Fcaʚλ������Də
<�����P	���`Ҍ�`�5�Zf��
������8m�+,	��r6!��l޹����Dh���V�4[Db��k��s~��&��X�g/Z���m+MF�G�F�� � ��_��&P�IBπ��EOkYyb! ��ܼｗ��z���~�#���k��c20#Q��z�1��Q�e��{��Ĺk@���|>>|"�':�HH����6s9�l-�0�(�h�߯(��20*�=�>�z�]��8�G��s]�\؆�W}yF��w9nMvU`�x��Lw7����<Wo�l������!��f��`��(�6�M��4X���1Fw~��m-�o���_w�LCiiFgڼ���X�j�0:�V6��=u�d,xb$�"�o��GpDsٞ�"�Z�����2s~��6X��A��9yE5i�F(�=�r�6�h#��f���5nm�x��~s�rD:�&�i���s�8ōL�?r��=��n�gU��N$����z�b�fG����I'I�}�۩e-�����,�U���vf����`�\E�\7�;H]��������m)�L9����G6t�=vz��.{{���1����l$8���Z�5��<7�q&�ϵ�l� �7H�f8a����2͋z����6��z,Y�r���Rn;1��v���ݗPD��ݴ��닡��5s�cR��.x���W'r�h������4�A�@�K���]Y�������x�a?��ٞ�8�b�#�9���ұ��6=�r�lCh=��m����}f��6g�� ��Dq�w�^QNƂ2L�N�OcX�w960#ڣ�}�n�?H�ě7��1[1F��.��E4[Db��b���yJڍ(��-g�罯�E��Y@c���I�&D���Ӎ�ֲ�b.A�{��GpDb�c��w��jg9����`FA��ױ��)�iF1F���^@��)�����h,6���bt	�����-�-ʯ�
#�@��@>��m䱬4�5������b	_��3��n�^�&5��o�=�k�E;�{9n{x`�<Uc��h����l�j!��(�_��2���\�1�������G#D��h��#a�f��^FҶ�J5Q�ο�_�� ���v�VSylDI��=h]�7B���:�aݮ4�'k���R���~>��������^�5���b<H"H��g#��Cb'����`FL�w��L��Ez�ܢ��J0��0�5�r�6�h��s���ǌb��i�M��^�[����kv�x�L'^����gƌ�(�N\u�U�m�Z�Mk�ٷ����*�Qii�9�γ3s]�`��ˮ�6�}�c���!�4o՟d�5��MF7Ϝ�An4�!���˂PDnTw���ރ���QO��FBgo}��u�xĬ<Xe�^=���c1�4�={�b��4A�4L�v��f��+�w��!�q�b�������mF�MF!���`V�`K1��p�)�	"la�`�Oә@�r�=���� � �5����b"����l�6�5�z�kP�絚9/Ia�l׵���m�]��x�ꪱYE4m�3ٿ`,alQ�bG7^���L絹y�؆�����An1���w e�wF�v�yE;h#+???}��o�!M�L���(����Q5�=��kz�4J6g�W�ϡ��f8vY�$������lCbVҌ���-��A�4F��{�E4X���On�3�g<b��ޮ�6���҈j3���V�`Og>�3S����6�f�̢���{7�`�x�5�;x��~�#�Aɻ�r��mZ��הS�X�8���w=��7x�6��F�{9��~c�1	I�4Ѧ���ocb�#J59��䱬4�Q�l�o�~�c���K�rx_gIٰ�Acu����dTێ�	�Y1��-f�v������_V`��+7�s^�Ģ9��]ʦ�b�N��?��� :{>��8�6n���!ڂ#F�W��)�l�7~g(���Xx�0��{���S|ֽ7����iF�Ҍ��x,-�4D�!���h��M�&�3��/#i{��V=�ûVҍF�MFc�
�l	f=���:�S�vi�Ӎ�ֲ��BA��s��؆��z���\��e�8��FC�2�����s�����a(�&�yEå:{�ϟ�����}%�z�V�ݣ�G
m)C`b�h[n&��DĻ�1:f�������vZ�WQLCf���<�آF���v�Zk(�`A��y�]�����������b.B��`������mׄ��H��&9�e%L�,���z���m[J5��ΜuU���o�a�(�#D�˴Sح�`{��r6��Pj4���s��Ζ��g�,��?U<:���*���G��̅�D�D$[�3���84����jo�����с���W/(��4�1F�y�^F�`�=��t3�����h�4F^�x痡�]����끶!���h�ג���d`k|�r6��h#�D����g����;��,�g@���a�v���8�z���%�ۚs�;���o�/�;���GF���9R�M,��	�ʯ������0�1�e�4�'���`�b�lW�v�6!�cJ1�7�ొ�{U�t��\��#Dֱ��)��#�!��9yJڍ(�iD�g}�`�3|���|/ʃ��W���U`�HX��y$:�h]<�rC{n��v�2#e�5E�>~�����P��h<8�[�k!oDR��s��r; ��AMd�́lCeG�j�B�������k�J0�`{~�r6�M��U;(�`uUX���-�3�}�[b�#J�Ru�w�����̛��������؆�6"ԇ}���!�">{[֊����5�y^�QNƀ�!��R*J��l�`#����$�bQ4�5�o�V�6��#B���ȱj~�������$�څ+j1�l���
�����G�+UX¬���9u�d���,�jt�o��؏Hu���!�Mq���9��Z`FFh׫��)�y�]���:��Saj���i�4M���x�!);F�4�}�0�ؠ�4�Q���k%����W[���	���[Ac�q������.r�&�=����gC<e�>�cy�gS��S��kj^$J��;�ޓ�0ָJdCBE�'!�����v�L�ɗgD�o	��,mBI�W��l��[��Y�Y�K��:�v�.��"�'$��`'+��^	��Vu��K�p���6urڲ�����M*�b��#{B����vx�+(r��� �ک�G2+Se��MVͭ�M6{3W!�:�ɀ,Ϩ�N���@��P�Q"v�N��E�gs;��8�'W��e;��Q�5�Tp��Mf�_K�����-�2�]fe�����z�>��Yf�&{n�7JC��_#ՠ�֮Aұ`�궓W��i�L�Aپ{�V�Net�@_X�]י���ms��`E��7��,r͈ވ5j[��nr�\5������w�����3�k���N�Op�F��lhٯ��'l�M��Ӷ��y��wȐ3s��䰞r��҅m-γ�@P������ێi��j�;rn�S:G�V����c<���We��]Ҧ�{�\M���YST[�꿷M�8;�q�I��X���r�
ͥ:���s�K��N]e�\��9Xl1�754�2��غ9�ssp�s��͋�rz6Y� ��m�]/��ojR�ÈXzH�0��*</�)�������ZsK��{|V�S�M�:.�K���wgV�_M��s8�9�ɮٳ3��kW[�h�v���2��r��Jyݦ�of�J�omG�o�!�bQ�f���u�'�?�����?{=�	�sJ�+��gv�\I��Ѝ~��G؉�1=i(DȽ<N{x�OϏo<�"�L���N��LԮ�C�U�5�$/<U*)�W��<Zl=����T��l��-I	;V�욖d*��x�OmQNz�2(œ��ކ���1*j�uw#�ex\���Qmp����$�+��hV�%efM�v�2�l�0�9,,7�Ss֌��A�8��	�.�iVg���&Q'�d��)'ՙJ�2mv�	<�FT�Fɱ9ꚉ���J��ֺtJ"�0�58�VInxP��H�員�"�]S�9�6"N�'���$*�H�HO+�؉�_F�0���)jI�� L}�O�?�*]k4��QYFZ���SBTܘ���T۞4�ݢ������K�DR���K��c�^ݞ����[��N���6g3��a�e�����;<
�g��T��T�]c�j�[�w�+f0ƣ���q�*f)%��le\C��41-hBĮ՚R\X)5�Xe6�3o<����%\�N����k�X�ڸC�;�FU�(k���P�e�XG����ϕ3�|�>6��yLs���2R]�� ��Y�&1�nW�+Gm�d��9Ћ�s�U��3ʦv�0L�բG[J��n�0�[nA[v|!ڜu���iH����loH��l�x�Slk��^"fX�N��l�5Q͜5���5�����'3��[^����q���FcB��$�jk���2��]Z�Ɋ�۶�ǒ{)_���Ư��1»���!�3b�X�����ha�xw����<;��d.F�ٕױ,JF#�3KM��;	C0tz2��Fa�bQ��\pv�S�qB�;=x�ؓ�!�����0]s��i�>H8����2X���7�]i�3n��#�j�ͱ�)	�M3LH�;dX�ʝ'�g���v��iN�:�����Pd
YC�E�vEޜ���;s�����.+gs�2]Z��'V�@x4\�K�:מ.-q�3��:�ꓩ�n!��0LQ��*[�װ����m�H��oR�9мZ�n�IN�xG�:Y��� ��7�,xh���8���e��G�2�ع &�X�k-�,#ȡ��#+�8�tpq��s�Z�8�u69�s�nBK����n�^��lc��q1Cv������4���-sԚ�΂f��M���eM��Ŗ2r�arb�.���7�DnY,췍N�V��j�a��zݜ��)��+���L։�eDͳMBhJ��_������}��kW-6���2:+F��%gFR͢�L-���[�pY�@]�������؝W]����h�X�Y
����� γ��x�yT{S���zb6v��*���8j�kOe�õ].;bM!!�8c\�]�vVC�ژsћ�b�T�lc;��y�a�MeG(��#ٌ],���"ꥃp��q�����7\��7V���d1,<�v9�[�p��7��������gcXx��j��,Ck�iF�J3���XZb�Ch��q�Z)��#��ͽ=X�f��ඕ�Q�҂j3� (�.�8s�)L!3)A��x�U�CoD$]��\���1Z����G�s��e�##5k����j��F(���_9,=�sZ8�%�5U71��U�h��h���XL-�0�(���{Y-�4�5d`s����1���g7�؆�6#r�w�.���7�=����gs�zZ
&�3(���G���,������k<��iF�J3��`�1[�"h���uh�!�[�w~�il�1��g}�d�W\MF�MFr���-��(�UUa��,m��˯s!iሒ� ߹�7G�{��x�pZ=��2oW܁l��h﫚�)�iF1Fa���-�ƈѺa���R��ɀlp�(��*TDđ	�y�mp��&[�唱;3����e����О�]ǑƏ���cb��1���k%����C`k����A�z<��Ɵ7�!�:ưX��7��u�k(ö�2'5}g(��c�1�0���P� A�z�؄q��wuIP䴵W�K��i3��j���{�l��rTD�Qa0�@O�<���}n��Ȯ�8IF�Q�7����&��{� ��i|���lCbD=_=�F,h�Pa��`�JڌCig���o$�u6c������xx�L+�f�8�S��B�X� � �9�6A�n4��}�s|����/^3��X��Ch��5�a�l-1Fa�{�-�m��#d�J%!fT_����;�� m���4�Q����F���F��`�AiƂ8�I����w9�{OS{�|؆�7\β�;��-���V�%bd`w��g��Q��Q��7��+a07��^Em�!u�jц�h�Q�`{~���j1��=�o����jK���8�ҽ�'��-����[8�����z��nkA�l��eq��ʧ���7XS�bE��F�����2�7mq����sy؆�kx�*����g�6�Os�F��Ɋ0�=�s�����P�7�b��i�M���`�أҙ�>�5Ŧ�˾��YiF�#﹒�q�lDR�7�.�� ��gC5���1=�sٞw|�Q�!�S<g�T32��ԑ'��o���Op�S���Ҍ����l �#Dh�]�c�z��.�s�?5���S4��F��W�Y+yR{W�މ}f��
�v+~ �9E���`���t�G��s���l{������s�)�����;��0[�V5Pj3�9���^���*`uX��h48�^�k!�{�Q��z��w\�� � �^���GA���6X���{YE57w���<K�<��sZ-�4@���ea�`���-�m�׵����F�����[Yiz��\�!�/UN+`hd`CW�d�!�8�E!��x�pPDpa�ﵔa��Fk7�x��߳J�����+7H��,s֍�"��o\�cy��g��6����1� �7�'�Bw�^�[,�ҍF�f��ొ�F(�6�j��Z0�m�u�����G�b�X��~߰[J�Q��JFk}�i������<J��x6��6/�G����8�s�u�%�ĭ \�x3��&�8��s��@�!��j3U�k(��[a���u2;Oo84F�{>,��o�:NѦ�4F_����(#J&�G'����H�$A )��'S�ϑ��}ab��SAc�N1C|�����a���^��FE�t�2e	J%B�"����l�{<��l��r�k�(�6V/x,b�b�Ch�ߵ�a��Dbg��`��﮵'1�����F:��x[?
K�'O�8�h9i�C�5]I��g77�]�ɂ
�6���$�� Tg|{��6ʎ�����W�	 ��K��iF�5���X2�/����0:�c�4N4T��ebr����//x� ���3��X��L���o(�VҌCa�w�`� :z�ٟ��Ͼ�g���ڐ٭�%@`��#������J�ٲف�юn������7�Ae6؞E4xh�֯�[aQ��پ�K����;�s%��A�,㝣���b;!�g�,C�"8�v��ׂ6|�D���D��M ,�#�u�E�A��ͥ�߬�>Y���o��	'�]O�ۜ�H3gj�r�\���%D̢R���s���4(��B۷c�'+ĀNC��$��u^$r�BA�*���P����G0�ݤ$c�TH���T��T"��ɡ�͚�9�(L�BR�P��{j� ���t� _Z��g���!k.���tI>;�z1v4eҗ9pbfnr���Xu ��c��;ƛ���3o9]���T�)6릐��3K��E�'*�#�`�|�r�_�6���Q�#n�U�Jp��t��u�]���㍏��]�Y^�8��kCY�=s���f�i�.J۝�l���ܕx\ ���r��U͵q� \u��R�e�69�/m�}����k�Բ/��x�MPW�уb����hM�Gm�#�5�;8��H�fyn�c���6�6�/Z���g7=���әtʜm)Xܸ��aY{/TSQ�6h����mXBk�1i�3Hԕ�[�._����At fRF�7U�%�j�$�5u���\��� ���	B�)��3(�������҂�	y� Y�����(�x��d5�wԦ�-"vq!&eM�ں�A&��P>=�oASD���u��H$7�A ��ׅm$K�
&e��Qgm�k���cAWmQ$�=ʯH�޹̭uNŪј�'�ǭ��ë p
ѡ	��Fz?��
���j1��P$�<�@����;�ֳ���oz^�@�B! �P�2�+�$��"V��K��.��#�4B�ݘ�_�|���Z���*��kt
��n������~�����Pۏ�>����j�*�R�ߌ�(.sZM��4d��(=��nA���N��2-P]!�B��o-<r�4��Sco���7���v�ˎ�/��$�Z�ox���s��Sm����F�����d�մ*��)(���^= �� -������(P��P$�w\�h!��!2�EJ���W[â�k��eHTH��B�$���h�;9�$j�Lol�n H;tꏺ�\�2����;M�^sT
ׯr���v��۪#���H��T���X�m�Pb4K�q���H���,{x��}�e/�<%����y��{\�IP�c<$��*T�_��.�DYΖ���{[�h<U�N��w:a�@�p��Bdʒ�ʅ5S�TD����Yj�GĞ-܊;��H�L�����䶩zxRQ3*Q�u�D��� ��%�C�|w(��SԖT�ޑ������IX�u��Ȯ��}����Gr�j�k1��v��Ǹz8�X�ݞei��$$��k��_9u����󗌓V8��EݢX��3��<�
�oē��
� �<�ۑt�P�v2��'(!�8P��E%7}�u@�|�<���u����kē��uD�s��K�<��_<�-��"�gR��thĵ��_:�Wn��M3��Z�k��vf�Ͽ|��F�W��,�u�|H�Z�A=�(@��1I��{qWC�4	'{�
��$��D�x��?-1T.��!�O��K����k�I;�(P>*���k��9�ӆU9�wTlZ���j�����{;���캱���Ov��A �<� R8rxRQ3*Q�J��ˇ�<s��$�ƨ�O���^����'��I��"&1�o3��-shZDj�lI��C	aํWn'�,Uؒn�a�G��&��4oE�n(��6�*���K'���6M��&�Ə�"e32���,�%���SWm@=;�:�Т3:�P$���;_G������9�YAZ�h�t6�*\�aŮ��l�%�Ga�V7*�{�g�~�U���׾ 
�?����-��h�v�D�y�P>��T:�vB�I+�Qg���$����Nw����ڢ|H�޹y�sǄ�.�����Հ:��t����P%��H�=�7���7=�	�ފ��ޖ��g�*��VV��O˟M-��j���>�;���8�"�F��;����C_��Av�>>�
���0%f\|����`C�� =��(h���)�"C���C�/U�@����y^��\�8��	�H����ǀ#B�+u��oxB�1��y�������w�O�c^8�b�F���
.��2�;o2�싰�q��m�5�φ,�z=�a�[�6@����N��;/3�4̺&�3��F*�H�
�݋��kF8�P�޺���\�zTǰR����R�"�\Y��44�ik5���3μw-����3�tP���������2�#q0y�=/e{JN������U��tc3q{qi����a�@p��5�ې_6xQ0H����s���?_��T4K�m��|��$`
�� ��lj5ڞt����h�ڠ@&�6�r6f�*I%Y�ۺ�%�n�W"*�%;Iu�H��TN���a���ʄ	�
RH$�E=n��&�|I��W�=�j�H'#:��� O,�B�R
�5ɵ�Vɜ��p�wn$7�"�=�� (�n0�����.�m�P�A�2��%5S�T	�ٹ^��M6�=���=��A��
���M��߮�u�#ҥv�d;l�n)kn�Ұex�L�",�1��U����y�`��O�B��{�K�РA�yU�r�|�Nl��;ā��Q>T&0l ��bfE׷B�+����H4;k3ә�ܵ�/p޺hÑv���<���XKՕ���bx��{u�
��u �V7��v�\9�����hn��������'��νG�x���М��È��g	�B�B�I$����lSۍ� z��I�����[y,�ݭQ �w�W����:�����AY�i݌���Ŋ�>7<�x �;;*��o\���]y��9�Q6�W�F% W�٭MP$s�����be�hpG'eU
$��Q"���P7SG��~���~�m�J"��h��F����N3�Cτ�s��k.f��=��~iq���=o~z�I ��$Yc�e�T	�=U�H%���CyX*� �h:��_��	t�ܘ�@V{��Cޖ�d^Ⱂu�����Lh�A	�Q��D�Y�t&�~��E=c�'�s��u���&��=�q�P����ɚ.�o]�(EO��p�"�=�˽�Pa�ml�wH�:7��)؝^�|����)�ǵ@J�OW,2��+�`Di6�6�3v�9(���2v��؉�g^Y{Z��qC�դ���`��y�`C����t������R�^7�*&vG�4�h!pkog�4��t�\�������k���TMoU������i)�N�-�\K�>��Qʺ��5�dVPrά�C�Ds�V�WK�����^骄 ��d���S��d��*Æ�3E���	�J����C'U�d�ժja�+6B�7�Žvd�$��r��6�FE�ڷے�픅��+[��0h����R��SK����X����/�Ҿ���P�֨�����D�[��]�լ�nI�^�s)I�_@�{�����N�w�"����&�*�6DIyοA{vǒ}���Z�֪؜��6�E��7�r�����X��� �r�j��G���[��Yy��!��b	�J"���	��q$��	$HۡX���nd'gI�|����B�e��N�i�,�Nl2�͜�����wڵb� �G�H�j�NW3���u|����oM㕗G3Q8��v�t�ޥZx�l8彺��#�\��
�+4}5����޾$�{�0]h�9���K:�ث�ҳwd�C6M��BS�b��yN��1~~�b���Y�FdTM��ľ�1�2��>�0�/M-=L�g��y)�UdR��]��C�6�b�n�e[]���T��v���$�
4°���L����1+ ��E�K��4.ֈ�Q3&q��u�+��Ƞ�\�r�8�3,�qU-ǜ���Y�K�ԗea쒵d�]*�r��)-U�=+̑3��Tʍ[9�2�J��D$�쓙����%^{%����0Ɋ����F�)h�L��9�y�$8��W3ë��A���OȂ<���<�)*�(�IRHB����2��R�H���#];F�PժHy�V'�5{%�AJ��֍�p\2O�] �+Ur��	hȋ1WHA��,g2	W6��T�ru��Y�?��<�~s���>$�weP>&�����F��II���DΖ /�`P�}-�W����SR�|rok�V$I�0��(�(=n�@�y�W���/�͍xY�t���h�N�:���$�T��K�Y�@��l��i�k'7���\'4/L){eh
X)2�=�#	!Ņr�Q$u܊=�Љ:"�p�Z�x�S�(�;�&��eHJBJj��� c#�e�؍������ۚ�{9Рn�RP��70�O%�&*%(֘;�^D{[U�IZݫ8^T:�YL��ځ@���uD�P�ca'�&!DP=u�\�S�%q�vEezA �ۡD��{���ȮT��!}����a���<�zm�;ۧݖ,�U�0�^:ǻ�r^>�qrC֥Wuu�;X}�� �᲻Y��߰b���T�
I%%{�6 	�kw�}Ӓ�C�]O8�I�mW�'���u�
r<���>|����:�^�mڔ��kk7:a.����>c��`�rAQr�����gk6HO!����>$�j��uGݻ91\���Pk��%�j�#�
�ф���vs��x7ݽݮ��	;5�A��U���#�����+^Dr����l�A)	)Q���{/hP'�p�=���Ix�P$u����Z�("%$l2f/$��E{���
� ݜ�@��z����9,P�7�TJ�1á'�&!DKr��uT�]i	rm�#j�����hP$��3� v���z�Z�4������6�3aZ©���-t��wo0Q��x���k��֥��u�YkKw��9�;�4���{��#�e��k%�o3��6T~.��דY�rM&��v�B�s��Z㇁��N�;t�r�=��ًۮ%�K\���-cIeip��ѫ����m��<�����/�r��A���O'm+��玎��e��[��Q��b��0^����\ɮv�n�t��a�r�G�t�����E�{JN��*��m��j�\'�nX��f�K�v�ra^ص����N�'V�IQ��p��J(��W���	��TA����N�b{�lz]UW����V���
f� ��s�&����;�-R�Nn5D�}=Q@��+q?6�v���	�$FB�ٮ�B��uRA �UIrWj��0I'�m
����Ӆ�D]�A+����U�b��Xt�^� �������o�Иq����(\�H�=~�j��m$�>9���_6��3���$���3��
�"��W��Yؼ.d�\�[6�\���*�-
[��vr��jx��]��^ �v6�+�ݝ�����8�V#d�|$z�>�����kt/3.���s�����}�+&$Ι�BI+�:��٘�%�Qh��κ��"gQN,xʬ'o�47a���Z�r���^D�լw����k+BaL(W���݈��X+��)��������	��� Pɗ�+�'n̊��r�&C�eE��BA9�@�m3�c(�:k�6�(�o��_T �a$!x՚����Z�鸛�g0�gj�@P��u�
�l�����|"I��PRv�'ǳ]
[��>�cZ��@�O6����mU��#���4��R\�X�]k��-�m�̗�a6C=��Imab�v�Wχ�a��Sߜ_���X;9� �F�j��ODF�؆�<��q=���k��^��TU
F�D���� �GTMiȘ�A��|H=�רf{D�V��P͉�*��"�H$��[u@�|o��D{�w���;Y��nL �.�Һ�}^��-=��3(7�@ȥKgt��7LCbQm�zNi����(��ʣK�{�W,��H'��B�>=�t(��A(�(�+��s��q*�w�ʉe��y�A>����w�is$w`'���ī� FB���s��(o��V� �管��O� g�[��=~��<؏8}����z���������*4�O�ݜ$�	eqK�፸���b�����$̙)(	)�n�x�K�uGē{=p ��n�����K�t(�#6e�D]i!%����G����R� 
��l '_� &��q�y������aU�6J%����+�}��<���"4E�����s[�P ��\P$j��$Y�)�Ro�e֩�mk�x=��R�H57T|M��Ǩ�u�7����iJ6�܈�t0��(ș��`Ju#��*Ǝv���W	-�����k�έv�᷼�	qVkWg�5��VC����$��^%D�Q0&QW���O�3�)��ɶ��O���I!�+"��Π��Ne���٘�((,��x�Â��ze���ܺ�j�̓ƛ�/՛8?�y���~FB���.�D�6h�E�u�4����o�'HP;�l� ��fI��B))���@�U�{�'76� ��VE���Aтd��)�F����˄���F��_MЂO��5D���{;b�hJkI�j�({3��T'5R*F�D׺;�u��y��\�� ;3S�{;�qn���@��D�Rڃ1 _H$�����P�L�:��o�s|�ͪ��D��3D�{qРO��eTD�̄.�E���5�XRZ����]L_wja��vT�9-��˘�X��B�����]K�wjK�F+�զ������� 6����ATL��Q���Þ̾�{<�)vݱ��v��+G(½���9���T�N{� B�8ЕOn���c`�9(2h�� 7��ʭ슝l����M�R�	c���fL�+�c�uaa.���u�J;/k�l��7c��;��.�ֺ�({]tÜ�v�u!����b�����Ī��2etvi`��ޛnM&���ӓˤãۑ�e06w#��-���}����e}I�}�$���D��gb97u�PW�O�f�$E��FB�٩�^�G3yǢv�D���T �|H}�T	#���{�^��(�L��f�!v� ]XT�����n� >���	�Ӧ/�;q�'s��^��p�2"%$l���T����%�N�'KP$�g*�GcʠO���.�t�WA� 
�q��):��J��PV
%�{#`V�NTt��� �@7o�x��r�x�{�13�J��_]P�Ί�P��E)���O�C�U�̕�X2uЪ�B���X��>�|�LXg����λ�$���Q���Xh�����@P����#B���f��W���Q�c6�ĕ��6��+��O���S�0�d�O���W_!�����Q��9�9�dd-���̦..\MU�݂������^�	�ܡ^7�ӄPb������2ف �a$!x:Gھ�e��� ]F7���.��c~"��$�� ������OmD��;Q�I�
3�@�{9�bS�}4�I��I�wB��s��H��6��A#��G�..'�����D�C�Xh@$ns�)u�9�A��^�	L�%2O\)��,	�݄͵\�e�g�۞�H�������O"���H�q�У�;6r�@$ns� �Y�N�y��4��+�vj�D��E��|����^�����i�ظ �Xh�w9�x�_	B#8�8�����j�KF`L���e�y�P>ۏF��qbhY�5���yw�cgbn7�.Uˬ�ꄿ W�c����%Z���^��vO�7�x�vj��� ���9?}_�o�>Xh	��С3|`@-I^7~5<�k�����cx>�Q�;y�A �vxოJ����	\�� ���dJ��SU;�@�;^%4��e�5�^'��n�gb�����?~����6+nq��ԅ�VZۣ�,�H6W ��"ʤU�)������TM���8s�ڠI �_!��o�m��e��\Q ��*��Ȕ)Q�^D�8-��ɨ����$��РI쾯P'O��#5�My�VH�ϐ�����@|o/�
 �&��)�fP������j���_U�j3eEQ�;��e%���Ă|H׵D��Gd]AY8�//{�>؇=]J����P��ڤjj��������B�;�B��ʑ=#M^
;X����"��f���y�| �M=���	���T�%x�Q�:$�����.��ʈ�2֝�ֶ��@=��@����#賂I�Q+���^.����_\����X��[,�3�Y�4\����Ɂ2%S))�S}U�I>/�ТH&�{"�ȧ�:�Cݏt�U�A �_P�{5�Q6����(]�n<��m���I$��G����Q���1q�x����7�ȵJ�@�X�x����0��.\�]*�����d�o;*���-�Ms"��u�!v������1k�	V���I.3�Eٜ���ONR<�W�n���35�2�"�x�:יʈ�ޙ��A"5�y��	�gU�!6�f�s �I�z�,_���]��8v�I6�L�xh��ʖ���H�3[ϵ��vWh��'�{x��ӤW^,ӝ��NS!@�f%fAJ��xy�^��H0X�jkl�ֽٸ�¡O0�{�e+��v�r��h���nf�Õ�`6:���8>]fv�Wt�AwZ�f���Ւoۈ;$�W�r�j�c1Rt�is:Eb�Bh�&���ou�wO�SnY�}0j�Y��&��K�-�0,3툼�n!��=l��:���{y��9J&0.�5��h�㋫�L;��:���}��G��}�us�n�ҝ�IڽT���7j�Qfŗv���4�y����+�V6Q��X�q��O��o���b��ȢΏ�h��@^_ty����ԥrwou�w��dw�6
ؤٕtY����B���ӽ�/��8l�gK�u�ͱ[��n�tC�0�')<″wt2�q1�{ƯE�Hb�4���WS3��c~�R9��jn�[���;8������)�r��:K���ta�}YWAk�qĻ�R�8�K�'�:��t7��� 6�b������a��h�� 8����+2��B�Cƚ���)9j&�+u�w;�D:�ؓm�+Gk�+�-n���jU��a� \�]�Ӫ>,u����Wg`�ь��V�=6�����@�B.���s۷VV����-tM�4$7�ZW}��[߯Ϫ�UJ�	�\/(��r�#-"����]Y�MN�؍\�g�HEAWQk�Dy��H(OI(��fB\��ad�%g��Y��ʢ$�����%T�G.ug�jIm�g���"�{��T��˕3�a���B��s�yм/Z1]��s=�r�����m��E�	QA{� I� ��=[
���d�t���0��0�-����9eVFk�Qs�Ē뗵�1G"�"��TP�4v\�T��,K�OJ0������R�A@Z�UAB��L�g�nk��e(��eL���ѵDs�""0C���^]R5�(�3L"r���H/49�(��rТ�-5Η�9��L������ߛs�9����/�W|�gm�9����"��k�n���x��T��;�	vwqu�uU7'���r���tX=��9��ϔr%y��ޣX���ñ���\�s��6�����/��ݧ��$����8]8DB��nڶ�H�V�94��r�0���۴����.�q�o-�r�K�r0���m���L���ݍ0x��[�4���n^箉�bT�|�:��_V�dqY�I�y�T�%��om�L{yųB^��Krc�f�v0"S�a�`�8N�p-�n�<����1i����3�6�PX뙯]1H���X�p�!���SgOg
]<Z�z�}hX���ųQ�m�,�� ,�};4�k>����/P���w�m��p�|�.v�2��g݄�łX���׮5�y�qŦ�d��p��'e����;��m���ՃJe}i�Cר�œe@�ۃ�c��7!��gI�̮a��B�n�׵Ź��$ބ���Z:1�M��H ��J��g[G,��"[�-�OU��n��G��9�f�\G���8��.}�Q���8�0y`�tY�W��>��kstv�q�]����
����e��")ecr�	�����5�#n���y��k����k��6�4XG�T�c�Cŗz�$�-=nn�q=Q�F�)�l�ԙ�8BW��mSCK���e�[It{"�k��nT�M��\��;M�v���������Ƴu��(��G��b�P��Ζ��v��v:�s�pFn�,.X� ��KtѮ)�J�\#1՚R!.��Q �	�T�ꢓP9'�,OgW�S���W+�ƹJWun�\��f��c�U�nd�im���a�z��ť"Z�=+a�v+dd�V�t�tP�5UR� �����ݡ��l ���V<mi��m��T�!�=z��Ԯ\A�l �3��g[����״��Lȕ	�K���
V6b��-�\�8�½�'�*2u��Ş�pͺ� �����nyK���F�����*J�W�����[�]�FZ��m�'���Gfۄ��t8er�]��=�EO�Kl�e�a�y��Zr�ӝ����&�*֝��U��%O=����u��B䎙aQ-�#v�=����If�)n��8~@ ��H���@��(�Ag^W��ٜ��h�"f�OU
��kĕ̱ ���S))P�g���K�Vgwq���Zx���h	���i�j�$@�U7ԫۼ�H�"%$j�0{2� ��j�O���W��v+~{�h�{3��}f�]���K쎥_�/���	� f�P�I���S-�P�n��;�4M.�L	)+����Ă@=��^�i#Ľ�����n����I=��݈���9	���$�Fb�����d��Z��|���H�v����D__�~�[Q�(�8٧������ �sTz�[�/Nu��Hy���D�������Z��ɳ�Fʯ-*��7$`�f��ێ��ϣ�Gu�5!�H{�����z�wZONY�Y*حڗr��21hAus)�4�_��̟�%��@����,
��5�;�.PAw��fʠ��V��{T>${�b�$��POo*k7�p�3q�	�;���~�ԊD�)#`��C<�u�Q�I��TI$��ۿf�&v{d�iE�b-�j�?��Fo�A �A���I��<'�j~���(N樃���lX%��:��5�}<�����f�Nm�� ݧ�{F��8w�2����cV�d��U�މ��t"&RWx� ���,����&��q2囯G_Uy��`����@Ф��A�����g�Yc�ڢ/{v��o�h�lnK�0�����-)	^4�r�Y ���R �x� ����w,M��Olj��
��`�Z��^c9	%󗪐�@٭�8��BR�{����8�<]�N�2R�1�����w9��˯�>?}��v,��!�^ѵt,�T�J�{�lC����AI� �>'���vy�������$}���>V4�))��I�`�d���~7SҸ�Գp+p�����./�hٜ���v&��}S}�$��13	�5D;�8�/�%>�M��y�	�c���tb�Wl����7�H��AL�~��	�� vg��3�O�e��o�Ұ��a�7t9��N{�7_@��4��6r�� +��]0=���m�Y<�<��e�\n��5��(�+�Ms����+Ĝ���{l<���~�[s�'��gUDM��A��%x��֮к��=n:���^4S����cT	#u�9o'zX�A�^�Ld��Z}q�E�(c {�ד:�Qz�U�{��'�#P��5���Tl9�r�ʚ�`���%eX�u?�ߦ�ON�fa����_�D~{�ﺭ�7���"7rhN��I=����$�g���Y�ѩ�p
�U������ciW0^�F�%e��v�_�g��2.T��O>|��'{�I �n�we<��53�&���,��L�� o��ER*�%�_d�PkAgM#���|I��TA=��8yk��ާ��;��7x
���Nw�7@
�|�Y�g03��E��쑾'�:��O�k�b���ɘ#B̢��afzՇ�H;-�$��u����NFE`�f�U˅�]U}c`gB����k�m��$鷒#���&Xx*f��h�٢�%��M�F�Y�B-CR�a���á��ǵ�Zsz��I&��G)e�Ǽ0�q���O��b��u��ø�����iiɃA%)C���uK�^]�����of�ۻ��w ��@�tr�X���eG����uh9-��v��뛐؇���'k�Mn .�	�y�+���drc����8�'�Ή���5�ήn�r]�'dB�Yds����ݮ��>x�쭍ئk{p:�R,�^z��ճ�뗔�1Xy;:G28�T��V�.�m���Y��!�㩖xg�c��Y�%���.�H�z��ǧ�fT����C��$�[z�Y���=.����s*Y�	&�7B��w���r�{��@*�V�#�=��h+M�E�s�S�VO�>Ǽ��'��8���}:�BV�e=9w1�R��
�������레�o�c�����`=���t(
�=-��?������i)+���dz�m��� ���� P�-���U�0��y淀^>�@���dVҤ.�P:k�yI��U�ƣ,J���T����.�O�ؾ��M�rs��$��DĦ3C6�X�"T��7�t���������N�]74^3�l�YY����2�_�4�u�$�6�F�����EOYІo��^�% Gj�!F��fT�����S�bWY�;�x�t]ca��FR��fi#��gkF��M�Sӛ,:Ƿ�<��I�2{�v��|,p�fn��Pt]���7tM]rŷ��#�����������9�P��0(	��� �ϱ��>��p�))�1)+��B�� �ƨ�|vl�Jo��'Υ :lO�S���q�*��+T,z�H�|�!����*��I�:�	�������Z[�D` I�T��f�.��m$�����{�J}ۖ���$J���[�B� ��틬����}}}����e�r��%�p9l#512�d&63p:��I�3��[�^}�cRy�$$������D��;{v�1���DE��T	$n��`���
eD��[��!�;�L�H�ǔ	#^:�I ����*�5{~�(!�R�wj��i]���>��j��V��͇sqn^��<�J�t=mZ�;���
*�ͰJ;�-IueM"���Y�p�f휱��b����W[YS����_�s�>%�mP�����Ϧ��% W�J�`�����R��F��	�ovŒ���kG"��OjoX�z��q%VR�j�'(z�GR�	��f��T���VH��^���в\_\׉�?'�E���������W��0i�v�T�"4�$��=ˉ�s؊m2MX��?}����y��_�> O{�} �����Av���}R���� T��J�wbȮ�H]�B�����O�z6��u�$�s�m߉���O��&��sy]�����#D�Д��Y}�� ��l�(�Q��R���y�P �۷`��}r((�X@�ʒeJS4"�U�B�����>7y�b�F����o��ޒii��17r˴}���f]�|�Ҍ�n\��\�5�%�!Ofm�6+CS2�S�k��0�gS�K%�����P�K$�鏽�#�_�8��JJ"V�|�ƅ 7�ja�1������>轹�<os��]\`��u��2�W�.taQ,e�S cm�7'WY�M����^�-5}�����P�R�Q�˻ ��s)H��o�Z8�[~��'e�y�îg�J$�<ɠMWW�bt�3�)+�Օ@�{}"=������i�e�������&sWq�YY]152dA�J3(�(=n�'�39Q$��lB�U��3r�C���&�I��T	��GI��$�W����+f����d��� ���@�u����h����v`�o�hɼ, fe	�)���{^�y��E�R��מ�r٢A׍W�$�}�yW�S�U{3������7#��Բ4lffy�d7U�;����i���$7f	��c��\��Ƣ�+�5�+v+�#��Q����O��.���ט�X�WV���ά%�������B=�*��6�����]N	}n��k�*[��ԊQ�q��f�����^�qSf�e44� eKXш�mQ�k���V�`�c��1ŎM8���CGb�lЬ�*G�v�u îJ�F�:{>n���vwL�"'gHf�{C�6c=���ɨ*�(U9��#2M�t#��Q�ݵmѓ�*�Sg�����¶�ns�Wy|�5@�A>��n��{��-8��Of:�H�T��T)@��ѷX�62����dgg*>��n��4��c����������(����񿀡S���ӗ�޽��8�wZ	sj�A<�m\������(�(��q=m�[W$�I ��T	�;��߉����}���q�S��%��xJJex՚��~�H:]��2�+����+^*$Ay��_�}x��y��W9ݽ��h4��j��]��Y�,m��,�XL�<��(HJW<gBfP�*R��S�T	$�]>�U�:Ŋ�V)K�	#��eAJV�Q$�V�d��k�ϥ�
��nfK6r�V��I*
�#fD�`�جݒ�\є
KsnMF���%k��*�S��1{��)�_x��s����!�x��v��\���yˬ��Õ(+�U��=}�@
�L?��Zt�ۍ�I�����@�U�$��� �J�U�zK[e�a9pp�r�w`�;�D�����v/�]!�	��{6�ő34fA��%D� ���|I��Tɻ����B��>'�z�Q ������6��#�t<AE����	@Q�A�hx�q��ۮ\�]l2oZ���}~>�;�n�楼_X�n��5�PI'ݙ�D�P2Qق0!��W`�Cw����X@��%ZWm���(�M�ܵ�l����<H;���ٝB�(����'��v@W�|���""�v��^�$� ~�d�h���Ҁ5X��.���LEd�w4�����r%��.pNqg��	�V�ӣ`M��9����aw"1�-�{E����e9���Z��X˰������Wfo'øXLG����WN�0Z|��NRal���²+�����a�c���˸E��p�ԗu�7�<͡�����%�u�
����l�ۮ�sD��p��ɺ�g� �rl���[�לFC\/X�*��K;�%IM��w�.���;gZ�5��nf�d�/�bU�rv0��t��؀-��8&��.�l�c*��;;OuD�:~�Za��ٙegeG�1CoL�C 4��xfY����c�S���r<����i\�w:��P�}��r��h3!Z�d9�J�LZ!ɝ��v�5�׆ ��s�g`T��*���B��@���0�5�Xo{2aF��5�^�f�Y�����-GsXQqT���$%�g�x�{��bC-Q9 U��]\9e�)A']��90^=G5���5�k���n:�I���3����ؖ�8�5,yz�Kh�]�-�{K1�x��V�g=ʻ��K�������tGlKDuXŷ��6�4O�VT��M؃v���b�=��Jw0��Fۜ!�霵L��a��oF�ȩu��aȑT�DP��h��v+3���t���#!����CAl�����{�|�vy�����u<�=�H����%u�g���G�������̼�*�(��)�86�y+�Teۊԗ{��K��PU�ew�0��vLV��
�Su]]EP�1��ݜ+<Դ*<Ե5vڃg�a�J���$׶�
KQd�W<��q�:�%Bb��z�Z�����PS�%L4Ǵ��[3"0�O3�!LJ�2�Ҋ�+fʑ,rܒ�$/5���]RL3u,��-)=�-O-q �tr"�C3]*�,�M���H�Ҧ��&�:.��I��Fa�I$z�N��*��AUAT^UT�!B�G�i����4�$��5�ȵ���]��C3Уմ:���Q�cd%E�d������E^AVL�3#]]������f:�U�_3�y-��E��0�#�B5�I����l~���f~n���^Z�
�j�K���JD���:V*�x�I��|ۍǅO<	���+>��4�
o���*	Q�)+�=��z�߭m�Ö|FN��םT	$�΢2o"J��_�G8����@C��x�ԡa��GC��u�����x�̃=D� �Y��A&�5Q$�{;
4fVr+�.�JڢK��@��O��U����@�{�Ҁ�����r��Ez�r�I��߲LL�(��j��tH12�IR�f�KڢA'��`�"f��S20�%ds�T���~����)DA%+R
2vqF�f��:ɖ� }�T ޽u`�����}�1���7�H`��r]�>�N��YvSNWuN����$�m͹�@�],3P����]�����/�Ū�J��eB2�J�
����]Y���Ub��v'+�T�μ���hW���w��/�=��fZ��S��95��u��>.�-C�Çq�`0�we�Xպ��
S�=����B�O�g<1=��  |7ى�>��S�wW'��W����&f�I12t(�D@��uDy2DD�
NR�I<�mX$�w��Uܖ�]�ah����IL��kWu�>#^eG�#�:��5h�]�	9���O��b�(_�m�ʢ,�Ju�<�L�"�%�B��I �muY���(��Ꝉ�T3���M��f�QH�	)Z�Q�����4%�!h��А5�U��H=���$U�����)��w'2�߼�螣�%L�i3Z�s8�B��@U�j�P�gQ�b�|l�t[���N�0*F��ՑQW�c]��W�{��jɓ&yH�h��4�-G)��Q6;[`�6�"j��m�6P.�W��pK���l[3n�(vt�����8���v7\�
�b�i�x�8-t����=��J��ɧQ�퉕��-v:���L�[B��y;zǦs�ҵ�t�Gn`ۣ,M���%�mX���.��`��.2�o�G�����.�n^�`���e�.ɑ�ѹ��g��hY,`�;s=����4$��}�}"R�R�JD~��~�H#w2�I>�ު�Gsۋ#�fh����5\_��QJ�II{�n�2��׸�w�� ����/c���%���d���'���AݷB�$��/P<ԫ��b��כ��K����}�^'Ю{��IL����R�@�n��HԲ��΅x�k퉹��a�1���\�AV�I�L�Fu�	���۶�ݤ���F,$��$:��A'u�ݧG9�=�����tǠJ(�L)v"�y��t��h�%̶�؎��-E3�j��}�kKjR���̪�j�$��j�{e�*'�u�͐�y2I�r�E-ڑ*fT�R�"_���$����`�-�\�
�d�tHaj�a��Ԟ�1Q8o�G�[��N�C;%��B����ʼ 12�'i��EL��'2�kT�������Q�@�ߪ��k�lX'�7������Ӫ�	�Ө"yI��)+��^f��ݐO�]∸}�fs��K�گGk�]���v6��B�W/k7����}���P �o���	�;}h�zos6I���	��g�I)��ao.� �6��,�3�&A�{�/ĝ��)�'(;[����^0X��!#0Q�j��*:el$J�l����� ���[�+����}���2�]���Cov���Ty=��'*k�ct(��2���DR����u�J�LG3~�z�mP$Ff��t�L
�#�Y4�{@5��\ʔ����[U��6���@$�zu�ї�#��*bȖ��c�v�����`���Ke>���ݷ�k� ��O/af�)�-S:��0�*�cǅ��A��5��ݪ��$o}�ذ|O��֨魨"uI��)+��+1.��1B�� f�.��r�����y��/4o�r�eL�Q"fN�(�(�Z�/93Z;ETv6<H���� ���(�w�B�u�C���@�K�HP ǌ��T�jLo������M�aƌ��sE�9�e�Ͽ�{��5r�����_�T P��:���t�m�^*��f���v��@+Y��"L�Fu�	1��WA� ޸�U��H=}j�Oy�~�s۞���>��@R�>&0�g�0>�Yev����A�N��N�:t�s��wj�V�魵=y��B�:�*�$�c�@��݈/x���TK���S���6J �+1LAaN$I��AYШ;�@j4�j������
�����ӻ���w����I؝j��AJ�I?yE[B�{�F�ıC���qv*���ڠA ���}1��V��78��&�Z�.��B�t�'�nϠ��/�b9�!tm��B.em����~��~��Eֺ�	35
�v��T�;]��o�J�W_*�%��F&���C�	J^5~5�[b�;��x���A}�*��>}�B� ���	��^8/����
D�R�%�A'��vHQ���'��Ĺq ���B���wd	���! 	)Z������Đ�}��V��Gn�$�]��W�-�/���H��n�NavU�V����[� t�t����R&w��w;��Q��Z2ս�C��pL����ݍ��R�q�06JAھU|�Q��w��:3��]e-N���e{���%{�ؖ8m��7h����F��]1�!M�5������q�cBZaF	�v޲m�ί�\��u!�CZ�����$X��a,�����0��n8�-�B�,�FP�\��w�Q�v��
�ԭ-j�&��`��4�	�ZҲ&@�\v/<a�]�r�B��[�ܼ�]�հ�B��Rv3�jĪ������U�ٽI�\��&'����:�W��ˎ��=������e2�nfF�0��e%�ծ�H7ݮ����@�9��fU��yT'�V�5	Цe@������$�[�دĒO�w���%�Z����+^`n��WZ)]�BO���Hp�-���7iq��k�x�;w��$���Mx���?)eB0�
����:r�DacH}��`NE��$��F�t덊��2E+GyQ����:�� {�UbOЕ$Z7��=m�
�n[ �3͋h��z��;>�T��D�HlZ�Z��nF�C�pOi:�ٳ��^�G�������eʔ�J ���ՂOܤA>$ngU�^�Q�A�=��`��4H�Q�#f$`I_j�� ���<��ň�(���T����~[�V��\�i&�Y�m�E���_\r���n��Aj�,��]!�����Z��(`����fr�J]jg[���ȓQ ��
fQP,�:�$^g* ��twL�\-���)���	�>��F��A+�� ֮��&�A�T(�Hy�T �w_1K��E��z2�H�L,�@�g��!!B�@���` =�������)� {r�	�Ϊ ���ػ�{Ϟ|7�Gݹc�r�8�`��f�.�qf��Jr�c!n�I"�+6�Ճ�Q����O��z���x�A;��ߎ�2�>���TH;}(BmL������P;.�şd�AO;I&�:�k�v���h�!dA'��O���8j���@�I)+y� ���R�����O��]D��c�w]{y�qP�+P|`�A�8>gbΣ��v�u�p���x[���j�ɓWq���#La�Ymp$��W�$�wg�"MD�t)�D@��{s� �ɶ��,��ά|�ś��t��T�Lp��P5�ݡB@�{����UFÄ���+�sĉ]UD��|�߯Ļ�Tr��O�3ގ���I���ʐ�;U�c�F9뇃ԁ˵�	�g�:�fh�����5��Hf�
�ʢHo�՟;�Tu
F��r"	����^�v,�c�&BD�BR�ȍ̯P��w��.z��A ���b�w�N��N����;��y@U'Y�Z�
RJTh;w~�O���^CK��|b1u��M�f݂	.�Dҍ�;"a# ���ެ�<ӭ��q%ev]������� :��>�'_Cw7��o�ԺLƅh��21-�VFwhK�خfU��f��Y�1\��L�|g����'<esj0�+�{����whP�k��I��TEM>��]f��>���X$��'@P��u�|��[PR�n���K��ۣ�����t=�p��9*���WY���N%[��Ffe_�������> �/��؄˚4 u���ă��Q
�l�$$(Z(��6)�}Aס=����N[�^ ���)$�qo����Y���"f0����̠(�@;|ר���`��U��ϼI!ż�� ��^!��jՂRAZ �����{o�7�^���2� ��z�vk��W���GDӑ^�P�K�0��RJ��&H'��_<�:'�� %�_ϧs`P���O���0%����Ua��f[2+ ��8!3��ɪee�Q��V���5�q���L�yF�z�͡�oU�o@p儱��n�N�ԫ����H �p۠�n�3��=��q3F��x��J\��qҮ���֙�����Ӄ��⁗>f���[A:ѱ1�D�"��lf�pVj�wsue��{ֲYj���\'�n:(,ۺy���nN�.oe�����J�Y!9��!WD9�*�s���ۍ�����n����7�7%�᳍�Pgm�����<W�OB�cu��(���[��o'	bck!��ϲ�J۶Q��n���ATy}�n��x��K��>��{>AU��W\wu>jdzmn��(^��1$]Y�9V-�#��
�{י��"+-�5!��7�.�l��
��oM:Qj������*#��`���]�X�h��j���d�j[c|�s6n������Qf�8q��e�鵖E橹C_j����Y�NԒ����aP�7�L�][�ó�P���W�i������r��ogm֑h֞�V۳g�]�+V yԱ�J���պ[�#�}�>���η;-J֕�Sͧ�N*HN���4:��_n�����w9פ�sح�,�s�ͷ3�r�{�ǯ���9�K1����գ�yw�MǼqm�(XTj6�n>U���r'8��~�O�ﯟj��Mu=�玝x���ƕ4�m�ON=ʒ^�F]��zB��s2jܼw��)�PQCx󓁔l����  D`�W<�1$���m��1	������j-svF"�y�m�Z�!TEQZ�6�����ɱd�e'�e^��Mv�2%��MF�\��E4)=�U$4�3L����fn�z!W��`Q�DE4�3wBBԼ%v���DD�[2�{����Kʞz��
:��\��/3�z6�$�����g��O<I��\l�M���Z�S���'S7"�"WUL�(�rv��Bb����������G�zaA��mH��=�nTA-[aG�ʢ��Lܣ(�*�JOTT�](�uLH���B�%"T��Д�򨲢˙2H�L7*�#�]�w���W�eþ�+%Xt ��gϞW�,q�L��V���f�q1�l��. F],�m�4�\����	�(��Dь�#�2Ú�m�lq�[��/���\xI��r#ᶚ�m���ͪ�c��)��c�+.6b!��N�\�q�v]5�c��phĐ�n��@�KW"�h��!���=�e!,�ۍ[l�8��m��`�6fq&�k0R�:�lۭ�q�s�ۤ�\xJ�&�s�&�l`�jkV�yʄn��'eaJ��>��𭧨w�&���u'�����JI�<P�ŗ�$�80r+֤���礗ۮ9:�I�)�[u#��-XxRr���N P��Md\W=����=DsXv�Hy�xx ��`څ�K�)*����O\�*x�9}�c����D����+h��y�:��M�L�Xݘ2�L�q���3sK1��Y�d9څle��y���1�bv�n;P�l٥.�45�F	3\�X!�ձ�%�+��y�V8ծ�K4+RR�f���p{*wGb����Tgz�3g]Dݢ0�w�w���b]\���C[.%J\ט�-�viu�KnЌ՘z�P^$7m(#��L[�m6�􍗇�\����^��ݧ�]۶:��%��qń��1�˴���C0{C��c<YՎR�뎻�V%i�ID�����l=��(Y��9,7�gNn�{k�	z#u�:���\�,fT�i9�+�D}�!�'�ͷ3;۱h����ĝ� �tY=f�9"\'F�v#n�u�jE��R��eD��}v�{kb�"�������M饶�^N;6�U�f�.�/*ip��)���Ekl�KWkH�m�>mq�+�X�p�utz�X@���(Flln��\X�5p�Ԅ�<g��\�-�m�R�j�fz9�[+�q�g��#^s�vh(]\�Z��LA�����h!C�v��a�dೈ����,lu���]�j�ǃJ�YnoL���햹K�-V�ՖcD�ݬ�s�v9�Pyѭ��f���;���!c���z��pB1�͵4���.A���N��M�WFvo;Z�('D���ƪ�hk��k���Z[k-�bd�]�8�ukbN*�B24pd�mP�2�5���0l���$�7n��CN��PH$��l��"�eG��>��#/Z	�_U�H�9$��
M�O��r�D��2 �h�̢�5;�vK�ڱ*��`�ˊ3I�>.�B�=��łf�L���sS�,��"
DP�'k�w6�}��k�R��N�"��(A���V�B"T�A��]�;�O\�kp� ��B� ��ͱ`��잊���{w���|�fҕ&! ��Hc��J�
��;�z�N��67@�O=λ�lWd׎�b��Oc�p��	�a��c<uK�%�r��M��fйs���R-�)<�/�V�A$��;�@L�z�g���lWd׌pЅ�����os�>���bd��&Ffe}�s~D�s���3.���1�/@�=�|k0]�s�^R_7"�y�_
Kw��91�:��Ι뫉V���N�P�~�!���q����F>�v#b�&��2�M(��k�](Ùdb33(�At��I:m�"��6�V���	�'3u�	�}���s"
D)D%��C=LoJܦvHŗ�`�C�ܟW^u9&�Oj���H��XU{�1*�BR��̠�׭Q�|ĄA$-�wd�8�}]y�^9���̹P7t���̩(H��]c��g�\�'1A�s�/U���%o���}��pZ�@�f��(��
��l�3|�G���&:�C�ةմA�M�������2T�)�n�籼��I1�|O^uP>��$����]s�s3n�S2EĘ�S(�>u}�(��w�*$^��e:�6T�w��n[���]A�kJ�@==����N�"���{�A^oL4��%T���>�4�K:v.���C��we�NJ�n�g�$��
'�:��
�L�233(�vv�k�����`�Ui ��ʢ	'-�Q�����ׇp���+�_GAfD��y��{�'�·i�����i� d�n��>��B�� m� ����v\;r��ݎ���	���Kx��CQ��Vy� a(3	J��\C�j�$���8
̿w����g&[7���n���6��D �s���U�_��)LA=z��s�~ۈ�#so,\H
�-�
T@)%nv���n>�� ��N>=�ײ)@^���+;}�]�P�&��(P�T+�6���a���U�H7��v �x�*��������F�а��M*��^_�/�PΠK`ú<�h~�ge��C�v�C�&�S��R-n:8��ꉅ��D��fen�v�m� �5���s�U��w(%K�O�wnW��x����Y �:H�#``�v��Tv�>��*	5��Q�Kkf;D��=����&JQ�S�@ǻ�g��Ok�@���n4X��˼ڢI?v�H�7������Ъ愳fR�X�uY8��	��ܱ~'�^MP���BN��}��ESĂFիh�8F�e� �<�GĀJV	�Et^P���
 g��*P�ܶ6�5�(�D�I)<��Χt�dx\rT�<;r�<��:`+ޑ��o��P]�bu	�0�"�Y�s�YɃV��=r��>����I��y"�=Y����R�s���U���|k6X]ܨ�)��TK�Y5X��f�q�2mf���u^^��cu��:0��k9
����Y�_>��={�j:�\@���[lS�=$1���"�Mp��M�[�Q�.�՚l]as��݂��^��r6����J��v�B�X��Z���*��c4�clL�b�"��9��y�s��7��G.�pC�nܗk\�����۬��ms�����=�D6�j���3����c֊#��Ԗ��8�uhx�P�W.�Uڷ��8��ݙ_[�zWb���)t��.f�C9����o&�$>O������ :��z���k��m}��`�<�E8sH0J�R�Tb�H�O\���rR��H��&�����U�@3qx����b&�e��XU���"JV��A}����jt /tNˮw���^O�ugU45�)D�*)$0}�����)��#@ +�yӠ(g��l�dY� �ՃD�l6�5�U�h$������ vo�L�m]�V)�b��OF��$����|s_eو�M�����O�K�ɶ	�D�e�iZꝛ��X��g�<��I��\�۟��Y��v�i�C���|� M�j�A9ϲ�B��ʎ̚u��!Xّ&D虙D�v�m�%\)��{��L>�zN<e%�йؓ�A̳�۷p��V�ӌc)_�{v��jRQ�VE���Y��i�d�r]��ۉ��tu��r$�u�UI9��ߏ�Gk�����|�l�%izA�W���BQ������ �\;����S���O��N�xs�;B�c��$!	B�Gf�Y�{�d3�*�x]er�x�z���㝗r �,[ 
�~l
N�Z	�*)$ю�˲H<s��]�y�.\ېH�YB���|��	=�43q�9��������~�_Z�\����Jj�ҹ8�p�CF^������v�)���˳���l��Ui_�����H7ϝ���ܑ0�OJ��e�{:���bȉ����"�5Α�z�1ٴj�,�k���>$���݂A'�q
6���ɱ�v�"'Dl�0'��� ݚ��bω ���|O����jzf��Y=Pra1b6��"%�#iM��N^F�T����j�i�;��d����&L<2�J�/S�*͍������ez�V�AXpq0
�R�T+Uu-��};tiw�.�'�+qQ$�Y��0Љ*�������Cם��>s��*
A a(W�ٵ�#���atyah���H�{v$��W�=��@�U�c�5�a���b���A iw`��
գ�ѥ�M���κ9_�'�?#��\��U�d��e
$�w+���ef-�>�J�h;~�>��a�I��E �	$�� �����4uC��mn`�Om�I#�<��տ��<����6I�E�(U6�ׅI��T$��v�aʛ��v�$��z��uQ16"8ɉ,LL���2��f��G��B�|�Uvw���ۙz��J��6�m]Lg��.����o�A*�v_q�Δ7,[T�w�2)�Vh�ô0��������c{���ꆺ�~2�A��d� ��T��P=���{uƦ�����^�y�TA=���^��ȓ5jT��T�=Be��b�՗`���i3�f�qZM[t��D�s%j��v��s��TE a(Y�FfP�	w ������g�m�oj�ҢI�fmQ>T�Q&B�RI�ӵ�b�A
���{��z�$���	 ���݂g�{���~N���5�(ڥ�I)*��7@��R�Wt3�9���T�P;9S���k�F��6I�(�(P�+��C5�Y�$��@�	��w`���Q{&Y�X�7���Q5�&Ǫ��$��ŒAo(Q ��&��=��(����Y%�b�Ǜ]%��J��7���;a��\7a�Y�wz�������u��|䗕���1�
�Y�;DA,����������t�v���<#Km6pK�zs,��v�cs���`�t=�mf��������Ѡ$sF�i�����`�t[
�b�Դj8�X�m]�Y3��VX:��s�w����<�a��ۣP��m�V��0ڗ0
h]����B�O���ĹvC2Tv��K�q#z�]RZ��$�n�N�x��zy�B��GG��!:�/S�����s��ss���3،�4uf��s���?yM!E��T�P�	��V ��T�]�sO�����w6P���'�aU��h)dF�*�;^9�+�oM�,�{�]z�yب_R�|��oT��	@�ч��`�s��DfO��[��H;ۮł	�/;I��D��JUc���)<S!*��ܼ���
�=���S�l��P�}� �7f�E�@YB�?�s��bfy?�dvw��y�O<�,���
�gP��C`��	U�8!-���n��ݫ�:@�[��\��W�V�P�8o�`&�>�M���[>٘�
�́ƌ��YT�B|h�����A'1�P'��H%?���~��f��!Do]�LO �+�*;6��m)���/V�q��J��S:#��jmg^�e���n�Y&Vdj��ܾ��H!�b	�ΪS��7s�׶U=�P�R
%vDm�xQ'ǷH:7p˻ڳ0�U��c�@�H�Ϊ�A�J�0�L Mx�m��q����H���P$��uD�^�x �	Z�E$b�&P^*R���+ă����1ѐEz�j���:�C������0�r�c��xJS䀘BA�e'�� �c�k��Iݎ-�����b��}��e��#5HO	u����T	$����]���?'@�����5�����(I��]�d���Q�6N�3�D�y�U	�z�аc-�E`��^�N�t�&
Qj^�Aۮ�o���q��8��.QR���H8��PY�x��� �cܹL3پMgS�˦ػʆ�Kơ�R�ʼ������`�!���
.�4mؑY�r�Q'kYt�V&�cW�֜���tyW�v.�[�%�r��)����7�)�x\]i*ԧ9[RЭ,N�}�,���v�ٮ���P�f*l�3$fnWs˽v���%��o���N�r[�1�c[���FND8����9��R;�ۼ=w]�ts�G�A��H�ؽ!�i��x��NY���Ť��V¼��U�{�j;���y[]K�5Gt�;��;�b6�	Цf�wx�@�$�ڔ7"GN�[��C5�ӂ��il��Y]si��daq��nw��R���ƻYK*�����Ni�г'�P��zP���d��lŏݷ��(��ٕ�������I�^���֤�kyy�LL��ޔ�Dv	�U�*+�����٫�fj�V�f�������x��sC>��v�!
0����t�L��ClNt�7��^�ύT�˟m<n{Q��z�i��TlLVmEp�Х�/z"�6�PS'A^:���eC�M6�촲���gN��ۋ˦w	��=������ɓ���!������sH᭫��ڷ3&m��*fJ1*��y�^#V��;�[}��q�x�ظE
�g)�y}��8�L��pU��x�«ܠn`��0P �Q-@�%�;��F���~�g�*UQ<kұ1~\�%W��^�լ)#�D�%O*k��*�}m4��Z�	�5�\��<UH��L�P�\B
"�r2K�L�a'�F���y��3ȍ"�2�8|��f��t|����&�"���Wm���꡹��Q�\��J+�2�RI�y����e4
�1r�%#ف�]-��s�ī�Qd^�^�f�&zz{iL�#q������+-r<#$�Q��*�BW/#%S�|�g��$��nP���D���ԣ ��@$��$�˵��I��EAW���SB�|�SR����*������f�a	RVjEy{��	�C����8�恡��^�TPo����!E����Nj.���y��9�y�8�t2�J4Z�e�$�Z)�k������-� �K�<����=����έP��J�AD���Dm�_g`�)qyW!��	 v�;��|^v)��tR�b�B��R2`!!AB/j��$nvP��CsqV�N/f�A#g:�A47��% �0�� �@_7��b&��,X\[
f�b�-u�X��
R�Q�X�h�YPQ��p��&P^3)W{]eP$��\�n{��H��zO7@
�o��P�&N�&g���TJ^w��7<�{:�H'��b�o.K�ٗЍU�ܮ9�T�UU�;���w��m�sO*�.j�nx∋���~$��������Ta>"�
(����jcfi�H������P f{���#����I,�*�~�Sh
�zދ����ϛ�ӗ� �H�1�i�����X�D���i�}"�rO�#
�d��-w��2D�W�«H�Wh'������.:O�+��A>9�D��sLuZ�qx�F��g*(Y�E.�� BX�X�3�6`�s�1)�\k�mZeڷg������Ġ��0���`�7[�W��:f�U}[�[����`�kj�"���0%�2���&@fY8�V\�:i+���|O��j��s�z�s�SK��'�Y��b��d�BaE�{T|I��	�*�u��k���'ė��nv'�fl���3�bfQ����nf�=�",����-��x���wp@ښ�3��P$�#I�)!@��O�w�l o�eIY�f��\��I#�r�Ēy����C8Rw����+�|���ֱ�n'��� ifJ̝�6��; �\M��Y�Uȁ�]��yugS���������I���Io��xFk�&��7(�C�d���\�v5n6������=��f�6�,Uv�f�37Q#-3`��!� J�-gjFk�[�q1��=zѽ`Ku�+����
�s�t�����	���\�s�q�g3^6����؄ɜ�&���e�\�pj�-˻e.z*3d�Hł�i��t��='πgS�t�@�v��îc`�b�m�	S��Kx����E�HS+�%	J3(�|GM�Q$�x�ĒHy���9��z��h�ʀ ��$*���Q"BI��,Y-�Qք��d�۱G����ڠO�y�����ٗҲv�ɺ�������"P^3)[�i��|��$D����ՠ�;�j�$����L$�ЄB �-�n��ws�t�$��T	$�΄��b���q>����t�� ����7v�	��J�
;q.+1G�K7�}ϲ�I��w`�A�ب��6j������y�C��.v��q�iyr$E�+��byv��NpY�M�t4]��s��y|�R�_'���	��A�ب��Bkh��N��HǺ��qd�)D�2�ՀF��
��R�I�Ɂ8��v��S�����ŗ�6�j��E���n���ٶ��*�ɐ-}�@ڇ�C&s>��.�%%	���y�k�nv���ؼtm�*ftC���U�AE@"BI�cz�����I3����# �qn�"��O	�&�ذH�؅��ӳ"P^3)]��R�#'f(EU�ܦ��3;Ofvkb����j�ڔ��)��`�b�\�y������KosDTE�_]�A ���>'�:�K�A�j����L�i���h�H-i4�s����z˱X�a�I��#���)*Vs0`p�S3(��I��d�q�
 ����'9Ӷ3v�;������*�9$$�(�P�a �nu�C�	���A'�qP �gP��MuLM��׻d���(JQ(L�7�k�Тu�z�Z���y<}�p �8]ZY��q[W�x�i)lP�媓0���'54
�gv�wpج��Z76�8O�gb����:q���� ]*Ub���M�o�u�*�9	���Q;3�P$�|�aެ��7�UZ�M$n$���^3)_j��H$�>v-��ˮ��PC�@��j�>|�]��2�M��I�#bL�m��p�:����h(؞l�����M�fV1ň�D�B!Gu�Q���O�>wf���5[a�}��O���T	���jb&en�;K���0�&T�F�� ��:�	�s����f��]�;2wĕ�����!J0�T��$A������r��/��vxE�u
� ��wdW_��RR�Re�N��K������H�iQ$�gs����9���8��\UcQYN�ت/�;�ɜ�s��"h������T8Fk3NN�:e˻���-*Żˉ	���*�gJ�¯����P��J
!$���H#s�U���'9/UUI/;���5@�uB�7#LV�j+�%L� �-�������X����Uwf:nfc�������±��Kxc��@�o��^sTf�Ȝ�)Qj�"s���'_k�fg�`�#QB!E��B�!S��E�&H ���b�y�P$�3��+�f`Z�kx��L�12�5gf�o�	����)f�T��c� ��H���~�A%�4�
 0�RD*�)��>�tG/���I��wd��D��Ό��w@�)�4��O���������Q鎩����mQ�<�"��B|Lbۻ��5^'�=���X�7j�w�8�ܖ��R#F�
|�T1�w-d��R�^"Z���;{�nm��;��T�2A�/�U�b��W��?�^/�#� m��Ί֧q���Ś�|=��h<]l��m6F�9�4��ж��(��y��#�\Fj��r��	��a�,��n1Ĺ���f�CJWVLA+��݄6��w3�G�;���Y]�ܖ9�h�n��,!f�&�\�[sǤ�9|2�:\��H����Y;���%��fڱ�5j��{%���S��$B�v��	Vj���c��7d�����G+��x�&� ����˲�f��N�:�l��nW&K��h�tٴ*y|
�B�]�^vd��$��,��8��H�y�tI$����P�O�|.�����0���%�`��% el�Z�D����r�$�%������_�߉��T�d�=���݂�Ԯ��Т)���힙��D�"�xD'�
�'=�����o�M���Tc�^ 8�RT
�-���I�w��.u{�i윸p���I�I$����P�DC��7q9\s������ �S(J�[�CK�g�lmwn,v�i4i�e����?}��jդR��N1FE^d�h�����t��ܢ{�.�kź�t�ĒM��>������ȣt�R�Ug�%(~&Om�:4��r���b��G��8��%Qpϼwq�c5�#'�5�����ov����s����or�9�h+�7��S]h�ي�ɢI;���I&�߽�*h��L�%�7K^To��"��"ƾ���@��p�D���3��<T�d���I'o�˟Bi/��Q��Z$�[<�kSފ�����r� ]}�	?Fg�%B	���MD���!-R$�qI+��(T�O��J� $��l�ܭ�w�E庢MznI	4I���ː�I�s:�';6�nơ}�FA�b�*$I�����\��<���W�b�1�h�͙���@𿢀5v���3��N��*�$���I�^����+9��T �h���&����U�WiYD�_c�L�q��Z����寡4H�{.O�5D��t�ĒE�w!��[�P�S��U��R�&Ϧ[�����*2I$�~[�|���tlwv�N�t���ʖ��ve96�>��Q���+�$ɏ!Y��g<^��Ot��,��n����x�s]ӽD��?�� �g�&Ik���H��H�Gݙt<�z�x�<Ov�P�I$��t����b�5�dV�9�^�`F[ݹ	K�Ŝ �T-
Q���I����*k���s��Gs��(�C3]'D���}��>�&`b�-��ݯb<���N"щ[	�Ykl*����ڸ :� �a��`��$�r����(V��p�衢I5���$�TI�g�HN����U��ɶ��hfy�d�
 +�X ��9F/t�	&y�o�s0�q��$�&�g�'_h������ 4;0ff��b�ߪ���eU�7j�%�F��ӦMI�n�% H��Ef9�;{�&���T����I	�Ϸ�VE�J� ����{D�i�T� ?v�$|I���9^�-��(3��Z�څY�:j;�I��1
0�H�znoq������۾�e�)c��]z׭	׋G9�gA�I��uD�����ڤB�]�d��̒�$�>����egK�&�EI�I����H������<�Y�>��TꝜcR���kL�E:b���w&Kq��ӎ�uWI"�>�^6|AQ�(w�<�ɢ@��r	'o��'���ǣ�сhn�f:N� On9P��@���J�СR���@>wrA[ګY$�j{���D��6.�R	�}�#h�сX�j����B~$;�I58��:��>�K� ��� =쾄�?����Dڰ��WD��m���Q$����׽�!&�#ٮ���A��]�_h�{�B~s��� �*T��e�O�$�k�ʛ+��ޓ��P�O�)g���޷���rH>kaI���~c� �����q��blm�$H!  J�?*��	 _�����/"_�11��DX
��)V�ń�,;��b���l�Fu�dJ����1Y�K,2�(�b�H BHQi��@�3L�o����Z��FQ���z��M@ ����=1.?��w�������1pPl^�� �Qied>�@��0����oKP��;
	�j4Xs��-}Q�P{��5�,�$� %�0]�q��*���O�M%��H �0ii ����6�6������/�������rC��Po�!H������@�bI��	 [��d��_�����i���*#��B�����#J�E���葐O����*�
�"O֪�L3����>Կ3��P~�Z���b�"�&�}�T]LY�J2�?��FB�s�HBB_��!$%��	$ 8-��r���-4��?��������@}� ����?j�/�B���J/������g�>�}����$e���O����Z>��$g�}��E�������� �����������g�Q	  K?��uP��?�#�V�_����g�Qf�g�����"�������_��A���ꌡ�?H}�A����%���~��@����@ ����i0|�����?��ȶ��3� @=�Q�l�bH I�T�@ ���������2F���pGܨp�� |�K��(��dA��Y��@V�Lm�����)P�ؒa����� PM,�,���>�?������J ����	v�0T��P?jC1H�@g&�췀�B@ �!����G�]}�z�'��~��� }��| �ɋ����/��ÿP���r?�`���~��>�,A?�?;P������w��J�r>Ԍ���c��"�/�~K럴�������!����#h�@ �K��/��G����@�}C������E����
�������Z,�4�aHg�����HT�D־��������|aa��$ta����������h\]>�~�_�}-@ �~�/�������>��Z�ѱ��A}���}P��6���~>��?���q�V	�$ 	�I0��`P��� �;�k�����?���I _�_��B���``>����+�;��4�~�A�j�ZG��0bG�Ѐ/���!{괿�rE8P�/�p