BZh91AY&SY`���J_�@q���"� ����bF��              ���6��!k�D*%RT�D
R�P$!"k*� 4ҕ**�B@�)P�
@h$   �j���J�WF�bT��H��(�L�G]%֕P���&�i��
빊���M�T�-0]� ��UB0h�W�G �);h� Z�ђ '�MhVE*�R�
��B�&�
��DE�T6h�)*JK\��Ux{YJR��$%%HH�)�JP {��N��4MXzn`�>p����=G���kw��2�6뎬/n t�7s{z�W���(P��6�(;�}��A���);2)( w;�=iK��=Ow��ƕJ+Jg/MR٩/-�uW��Jz^�T"�D/oopzU�\;��iB��׻�S֕{�������m{vy�P��Cy��I)=,V*�6��IP 8�\�����%w���JQ����j݁M9��ҕ�4[׶�x<��(��^{�*QB��Sǃ�J�2=��^��J���.x+���yޕ@=�R���0���$D���R���;�T�LGyo=��T��ۼ�J�t��<���S��x���+y^{�J�){�ͼ=*U�lr�c�Uz�j�y�P�Wiwz�mn�KuE*"[+B��RK��T��y���T*���zyR�Z���t,�H[����U^�(q�{�C��^������uZ�M�7�4*�o<�^U	z�/l�JlkOM���UJ�iysM�()Sj�U[-�5��JP ���UPu����%S�Ӝ+l��c׻���%J����U(Jv�{�W�F�t�wnt �ƀ��p(���@މ"���a�)7Ϣ�P ���{�� }K�t�+w�
��0 n۳` �8����� �ޓ�4 zX43�{� 7"�OFUQ���QG�%)  ܾ��o����Jw  �V�@��ݞ��9��\@�=j{�P�=Ǡ��/
f����B���Wϔ�� 92�� �����y� � 9���  �  �w�4�=��y� Ge� ��I/`ٌt�F��%$� 8� |�� ޲���l7�u�  �O�=�����)� �� <� (<����  U@�   50��Q���CL�P���D�i�IQPF  A�	� O&AIRP      OMMJ��h   �	2��*��   �� �	QISL�!�ɣLA�=O(b~������7�?g�����^e~���ȗ0^����䮷ˑ����� �
��  *�?H���Q xX$?����,�'���_��gʟ�?� h?Τ�I�Q ��yA�D�\NTE�����?���?ɀc�`�0q��clb� ��\`�8�1��c��1q��\cc�Č�.0q��`����0q�l�1q��\b����&1q��e�1�LL`����11��db�8��11��L`���`c�8��1q��b�8�����&11��Lb�1���11��L`����.0�1i�c �0q��bc-��Jb�8��1q��\`�#���0q��Lbc���&1�b��!�`����0�0�8��%�q��`�8���4��&11��L`��0bFc���.11��8��4�1m��\b����0�1i��\b�8��.0�&0i��b�8��1q��#���.0q��Sh`�8��.0q�c����.1q��8��6��L�4�1�c �-8�Ŷ�\`��&1#�)���1�c�����.0q�����1�b��1q��\`�`��8�1�c���%1�0m��b�8��1-���.0q��`�8��Č\`�8��11��`�8��1�0q��b����&1q��`�����0q��bc���&10`�8��c0q��Lbc���0q�1�&0m��`����&1-��)�0q��`c���&21q�c �.0L`����bS �&0q��Lb�8����\`����&11���`�8��&0b���`� �%�q��bc���[���11��\`�����`����&11��LaL`� �&01��\`c8��cƘc6��&11��`���A�
`�8��&0q��b�8�`c���&11��bc���S�0bc���&1q�L�0-��Lbc����[a�R�&0q��`�8��c1q�����.0`�`�&1q�c��1��f0i������b�1���1q�c�	�H��)�&1q��[-��ض���b�38���0m��LC0q�����%�1�S�.1q�c �F.1q�c �.1b�`��1b� ��X���1�c0`[%0b�1q��
a�������`�.1q�c0aLLb� �.0`��0���1����1��q�L\b�1�0�J`�1��\b����-1q�c��1�c)��6�1�c�10q�c �0�@c�.1q�c�1q�c��1���1q�[�0b��0Lb��1�cb�!��0Lb�1\`8�1�c�	���l@1�0A��c �`#�Uq��1A� ��(�W	l@q�LA`�cC���� ��*4���\`#�q�.11�.0Q� 0@1�.0q�b��Eq��0�"��G��\b
c��-��0)�!�Tq�0���G�\`#�U#�*����b�A`�c`��q��0� ���\b��Pq�1E���G�C���cb���cKb��Uq��0D�8���Lb+�Tq���\`�� m��0A� 8�S �b��U1��0�18��.0q��\`c��`�8��0b���01��`����0q��\bcbF.1q�c8��&0`�0�.1q��`�8��1q���1q�c0q������`���8���#�1q�c�)�C0`�8���b�����bSb��0`���\`�1�����`�1�c1`���C6�1�c1q���1`�1���0b�`F.0q��b����1q���&1m��\`�8��%0�&1m��b��9�R��}*a�?���Uy(/�"�����H�s]�Uޚ�kb��l�Cq���a��Fu(�T�ux�D�!e�^�r�-@XBX�7x7n
.k�s.n���CL�i���֩m���=����J^,�i�HT��FAL�(��aD�]�7s�)�u4���eneXpm�RYO$; Q�G1o��BDi�ۻ��A6쭛�����0u�Ȑ��C�ǂ��/���Î��J�t������tڭ��
�U�2��ކs�h$3V��X
�#�TA�.K, �-�#&��P����s/0:*�X���L��D�`m�֨���Sn��ӹ޽�&���On㘆*Ȍ�Q������,0�t�a+�J�+QLL���4H���D��B�K,;�`�%�7����L�eRl^G���YH�ו�i÷emj���"(ŔflGN[�#kը�C(j�QCمb��!X+K�ӹSjI�6����kh]�mЈ'�	r�^Y�4$@ä2�lE�<9)�@홣&B��Q>�L�DLӛd�4�4Һڡ��6iQ�6��5��X���õ�lfEV�Uņ�;�X�M+\2����Tɶi
	�V�%�x�Rc�4���,'I��e
B�Sn�D��R�R�`>�e��ER�Њ9b͍F�J��P�(��2RUl�k&�1ǵ(5y	�re��r9�^,��,��[�ScA��' �kp�u]��K��7��*�[eL��GV㥑,r�]]�룤��4�b�����93.�8Lf�;U�Y7�WD�5Y��9%5u,�!�ݦiU��M�x���Y.\����
�[A驛�	(X%[��Jȉ�%�r�aZDq�"�:��5÷��cɧ4Ԡ�kkHaܱ{�V��h6�����P�t,2��ӑ�#���QL�/ʉ�U�lFH���u�=�B�ζ�:"��D3�"-�˺�t��3KFTNL"�	T��j�Z�R��j��[s6����A�) n�+c%����E���
�<��Į�U��7d�uz!t��9���NT4���x���e��4�jU�McW���T!4��RZ(!��^��Y.�j��̛�ӌ��;�������;��V�!��j�eih��)*{YP�m�lf��K�yW��TF%R�&S�fR��&J1���ĥ�Hp�Y���M�A��j��r�p'~ӺȪj'��X�mR�Qצ&e��R�qZ��!�û"eTVh%�NR܅K�W��MlaW�bC1Ci�
G��(U�z���1�֬Y*��FEz���&�lm"��������[�j(_�ط*��Z�u�5���@�i������c����o%*MF�p�͍c2��m��hEٓ��dt��GȄ�`�Sq�Z&�f'Q��t)�9�e�k%�yj�a�m�Y�
��ӬZ��q���M�2���xˢn�-^�ugi`�5Q��4e6.V���"!�
1P��bJ���Fz�&䥪��S2J�˕uVrΨ�Yoj��UiF�$p�Z��@�l���8��`Ղ�$(*)b(l�m-)�KB�6�vC�.������/%X��$�/qBS�yQc�bȱ*���xj�b'.�x���M1t5֙u�d:lVRĘn�!b�n9x�RPՠa���1v��ke��*4�ԯO�V��z�����=H����:�@�N�{���S�'��ׯU"�vR�x�q�j�;D�Uw���2�L+^�4�LÁ��wV��G)�M+n��C�Z�(�m�+�qd[EE�),+Jq�5fY�Ț�����lEV��3v6Ð�	eِU����YwbfК�)�F�5R��֥x2#��$Gvb`J7F��L��m���L�n�m��"&Y��m{f1�r�$ԙ3"�{u�:,�����2�;��;�)طF�T��S���8]U���^+eM*I�Na�e]:9z��ʗR���([��)�c�ҰG͕{��C�Z�ɫS�nޛ��U
���U�&��!�,Éh�2j*�9DP;��Td��wy��ʰ2�i3\Uw���u1�SYO!D� ��#��]Aq�aB<ea�,�j(+iˢ��4X����[ܱ�pf���I�/pՅ�S0Mf�j�Mmm�+"�m�:P�;�\f=˶wp��P�8��rR+v�먋��D���j')#xE�33�6�)jW�؅���V�������:/3*lMؘ�@������[�-����6��zl�m�no���h����h�)��A$�XÍ��a�p��Sʺ����ZDql�6�V<٤�лZY��ܺͫ�T��e�"-t�YW�[�[������ޘ��0n҆l:��q���̨5�Y�(�F^k�:�CP�I�f4J����㬚37�̲�Õ��*fŔvI.��ڬU��'���j�y5Mթ
�o��%�HE�1T��b�4����+�wM��r�<r\���Lԍa��L\U"/Pi�'k,ʑ���"��fH��.�� z���*�s������K -�����pù�.L��D�����f0^�t�U�!`�����0�jީv��9d��w���@����!��,��)��,�4hLM��V�ɤ��b2
Ƶ*���y�anV#�X�	��F��j����ζDŘ$�����QJ�0�K�bt�`C����^o�)H�k�smM��-6C�j�IE���X�(���T����͚
ຳ5���L�j�k��`�\k��e*%��1�e'M@�U01l���G#�Tp��6����<�&Un,t^ڔ�w�=x�������ݚZp��J`����KR��r�]���w4tֺ�C���Kr
�4���7B$"�"X��sa���ѫ5k=2[��6Ș�c��윒�7�z�&�e6do��ފ����W�ŧL�p����ed�ٮ�1Pɴ�"�o6��V��((,w �),x���t��Wy�/�ŕE /n'P	Hhb�ܗ���c�T3*@d574�3X�,��6��0�Q&�7~��nRqd����.��d�n��V�1��w��j`��eษ��80������Z��w����m;�a+�0A/Xj"�=K4�k*Yy.����bgcw��D��E8qDFI�Їj
���H��.��C6�+���d�ܬ8"�R�5`MS����t��ƔథZnDr�Z�d��`�yu�:+i�S��"��۳x#�Ƅ�nA�Pɰ2�� ��i����Nͬ��D�2���tj�v�*���L����V�X�Un���K�p`�v��Q�JZ��uD)yq+��	"��z�u4��/ș5SUb����ll#swUƴ�e��^A����6����Umeݐ޼J@6��1��RS�k
�0��n���RU�Y��R�הnf�;���׬�Q��B2�`����0h[0�iZ%a�܌�-:�r��A��g)[�(�V �DoK�NV��:;�h7�����(b�$h���(by��3jo�-�,�wNm�aH�u��
Um��f�"�ĵ
�t�unP���&�0ͱnM:Ն۠yjf:rl��7`,Ycm�6�蹶!�4���
c.��ҧ(�z��.^L����=�4Ѵ��{�a�\^���q�";i��� a�Z��w7f���àm%%̠����k�gC[�2�,23B�x�U��[�����E0M���7��Ț��F14FS��Ul�0R�*L;�J�լ��x+73o%�
R�;�������w��6����ј��4�V�LӗW�mñƲM$��rfhFQ�%�Fh�����<���*
�t�jCF�wN�KtR7R�l̩v<�5m��2��w�A�QS��9��R��y��'T�i�Ö�v��2���Y�u�o-�CxΕ�qamŊa�&�ۭ7�(�Iq)x.��n�㎷Z�nTa�$f��+oU�h��F/h��fee��n8�D�,^'�Тi3Vf
�#fG1b�o%�H�"�k�N�*�ÖZin]ie�RކF�J�*^ᚣ("F���m�Ӣ�#kZ���Ej��L�%�yFű�4��'"�f��r���$�J�S���l���Y�TN�PK=sd���\�rU������,e�d-��86.T�E�0 v�ȵ� �n �^���-���-ڲڭ�ӬW�������E�"��GR
�n�[y���q�Ե�p����8nU��j;y{�á���nȓ0��w�̬/�ZPr�8L�Z6�Y
�4m&���1'2�Df�:R�x궬,GS؝ͬU`��mMա��a��՛Qc��{���RZ��
I��VZ�c�VN���3��`[��y՝�(ڽWf ێX9x��
ڍY�P*����xk6��t#��2�y3ZCq��"���u����`���Y�Sԭ��Ğ�w��D�e[�< "R�ʍՑl]ֆ��uڰ5� �t=�݅s	�)T��S��K(U�o�q(���qŔ a��S�����vEG�J�yPT0˼�1J��yQ6�Z�d�U �$�ll�܋Q���LK���z��;j� ė��l۫kH(��V&�U�i����Y��9�z�0�U�n%M:�st��ڦoN�kL#vܸN�Q6�l^�)e�f�H��G$����C��*Vl#�O�Vm��V0�!���VX��6�Ȼ���kZ�V����;d���V�fK��h��#������WXAM'��m�N���N�e'�Z�ZX��U]̪��jf��F�v(4�\� 8n���hY�Vf1h^�DɄSw�-��c�k'R���Fv�0كqz��Ъ�g�uu&2���j3h^�JR�I�x2��Xvg����-S6�XdF,�x�ӋQ���猐i�41p%�[�������������m"������FV�9�i�ɳ[���d����[��f�i)w�N�5�C5/�ÑI �x�����n�b����aP�y0����.T��xuI��fRdmn����X���a�Q��+�g�]<RL�e$�V�{-̵C�Ĳ�ݰD�݈�O`���]�"��n�Vh���-�Q�"��4���O����? ��b������W�_�����ݺS�Q���;�u���R����c`�.M�f�o/LF��'aV$�-�[ef�%͹Pd�72��Ѫ²���푒R8�f���wN��IT(h��ne^+�F��#k�^K�e]�2�%�Si�܍�b\�U�&�a�-̭���XхZ��nI�ר]��!�pUӈnY�m�-D�*�n� ��rB����N[b���3y��ԑƜ�Up�f�ƈEԽ���=��s$�)��ǄWOe�*߁��y�r�̠ұElN$Hl�bc�9L [w��Zv�Y6������8�j�����<hn�e�BwyA��J��ކUH�Y�L)���6�S_�z�*�qP��MU�i��b�w*�2.�i���MK��<�Uj�mP*�Z�)����J�D`��E����'��x�*��z���if�Iڦ�(�I�M6�+�p�%�B���ug-IĚ��N$�ҪO���KTjR�-]���U\��q$�I#k5RN�5���Ě�8�5���{��ى&�����b6�j�]��wP��f��z��%"I*I$����X����Ĺe���|��T��U�RQn�H���I-���OT��T�(��`�LWIr��D�"�R"Ӵ��2��k�<N��)4��K"�D�i�t����]W��ȩ*JR�J-�T�����j�F��8�/��}�g�?�b��Y�usWJ�V����R-�4�GU5��$�����\�'ԢmsW�s�uiZI5�I@���ڳV��G�i�1&�Vj��N�Z[Ԡ'k-bS���|���bēI#���(�N)��jMN��|�[�Z��J��Dj�cJ�>-�k)i:d�]���NPek�lV	i��"냴���4�u��3wfj�I�'`�|���]��m_�.�j��S_D|]H��%��ZW��?.弓KVmp�*��|��#�m7Z[�%mW����$Z���x�%K��T�q6�+K����_������q0JX��mg�T��Z�F�JjT���-�SZ�]�mX4Ղ�bR#���>J���W����m6��ŀ��%6'��"��>K\ĺ��Qk1kW�r��%��Ӵ]2����8���bخ�+�1�6�.��J��X%��IJB�,i�4�o[�4R8�&���Y�t��K�h*�#��#���EI\Yk�mkX�Q4�(�Z6����F��TM�J�rS��ڶ#�Z�W�ڧzb���I|����T��V����T�+�|�8ޤ�N�55,OEQv����bIZN.�wԔX��IZV�#�]�\�-����F'�D�\��kmKWI5�;Q�Ҥ�W��R��yo-��]���$	JR�G�)\T	ā`�SVb�J,IҺF.�NS�R�������o�(�.�.��w#b�J+jbm�֋]iDq]��Z��*�4л��k�}:�4�UK�N��]�ĵ)�S&�I$���\[��dUiE�>O�Z�X����-�Jޱx�d��r�_]�*e�z���MrU�V���n2��r�Wj�Y�AMg.���UnŪ�.rx�����)ID�<��*}�y�s�V#N���J���TX;m��M�U����*�9^���f�W�j��Wj֝��%M;I.IZ�%��MT�j楣���U��Q"rT�Uڤ�-ib��o�(�,K�U$��"�-J�Vuʉb8�Yխm���m`��qU1p�qH�Y�V�'��E$Z-$�U��J�I�V�I*�5*N�Ŕ�M�j��:OhҫV�t�(��]��ՠ�TմuV�I⸩$�
莬���OQH�NM�IZiZJX�q+Yi�1�U�RJ�i������r��~�@?��!�{�
�`��]ן~�$�I$�I$�N�����ky��y�WV��;��MOٱG����r)�G#��s}o��..��S/�PҖ�G+�Q)�����ת������whPV��i�"�ym�-ʗi<�:����aT�͵�XV�5j���G5}rd.�e�x����*�B���Xnp��.��;Bc���mye�!�����вp�-��gs
N�o���d�UՑ����T���)V��eQ�Ġ�W�":�R6d�YlNr��ӭK�lF��]�Mƒ�3��F���좸R�9��y�H#�ܤ����.3"�������/���u�as'l��I��H���O(4{��T6�g>�2S�C��ʹ����"H��1e��<�F�Z�����k�QP��P%�ӕ8�)�pnD�.X��Y����/�v���U�̰
- Ms�t��8�rw�M��p�-dt�wdeL]{�C���>�u���R��AY�j�M:�l5ʈ�L�;���v#�k3�}h�;�� ×���p������3��M��pë"��5˾��Z�f���uZ�r��/�tޠ���HՉ�f*oOݯ�W/45�0�2���m���u�i��uj�
�mm]!��e�Ŗ�:�E{3�;J�{�&���`��WO!}���ǜ:?m⧝�G|5펇�����esl���zP��]�[�w  ��.�0k�ɽ&��j�:��-���7�Zv�zc������,�6d�s�f�#E���0Ĺ]Ĳj�Ō�A�X8�5Դp陗�������Oc���6�4�z�#��[M��,s�Jm���\��uH)�-
�:��b�\�(�*���CsQ�(��/ʴ�^G��Y����&+��Dn=
�q׬��-{!J�=�8j�a�B�,y���� 攩�z�h���̷ut��>��aW���$�Ն�Wq����pV�"�ת��7z��Rq���o_!���7�P��*�ً1Vǈs1���v��9�*>�����!.�BvY�Ŝ*��beu*��l�g��T��E�*u���1��c���^�D��.��5��]c�KY�!��h�1.ZhQ�]:�*̼��u���M]�Hc�pI&����� ��4yMI͹��,�*�<Ͷ=��޺�D���,�ͥ}���FZ�M욕G2�!�9cy>�Tv��8�=�>�����\��QUcf��u%<:���] ��2=�1�0g�"���z��#�Y/�]���O.�>��:�,����a= r�s�\�V��!�p<���r�	w[YӾ�*�<{����k�e�[]��1��f���@ɂh����8�QWO����n�d�.F���-�f�,�5ۦdw�8m]̛�WkhaI��҄��y�D�}��4�B�q=sVkV�/��)�W��5T�6īP�uкĶ�4�X�8b��Q�}ǜ�Qw��%NmmL^niG:�Ҩ]1�R�o%-�c���&����7�+V!G�z�V�0f��QcC�W�����lq��������|��/6��v�o�ˉ�p=Ouf��|�ۡ�o�fZ��[�D�먺!���5�FBw8��,�hC�Ũ�뮾��v��wM�ǷbwF�e!ٜ�� ٰ�G�z��<0�������ud�6�(s�p\-e3c$���s� �ҁ�S�]�I��� {��}ۙ�>�p]Ilv�����p�lh�X+�K��q)j��Xw���c퉅G6vk�H�5�Fk�#5�ձ�;����T�O
\�������j��L`�1���]WJ�^�]v������㝯��0*��ƛ�;Q��q��9
9��V�E���h�b�u뜺e	�y��P�{�e��
tє�sx�B�ʪ��Vx���3h�c �I�x/Vj�ֳ�v��hc�P�r���1Ta��dUݙ(ݓqH��V�X�6.ޑ2ap�������N���*�mǝû�l�y6{FL�=�4�l�Tq]�[���Y�����bċ0�]���7F���^l=j��a��s�[�'��bG�jcWn=@��,��ɑ��v�s�5�,�G�;3&2!+���ƫ
� �r����-YԺmZ��V[�zΞ��\w��ҩfLc2�
�nTP�w�Y0"��Ʒ�tT8�Zp�̼�{���b�]!8�8vKKq]����7x:��m��-蕦�t��%iX���x1b�V��B��e�_NG����n�ǯ�nJ�հ�,ٷ@�����杽�Gf��]��I<��F�mnn��4^X[���A>�f��0ժ���z�a�unLQe�`ɫ��n����d� 6��u��*\�኱�lc(����Ly�dcۑ�G�:r��~S8k��3�n�P�vc�u��I/�4�:%�S��P,����]����3z�#��	�Q����2P��aa���VT.�6�38g,pr��Ғ�M����Y쥗GcAq��Z����R��i�����ɱ���Z�܍:*�E�

љ���4p�))���a�9�n@����I�4>����������f����&C�v����7��V�;���Ӓ:r�Ε��VdΫ(�����|�
K���|3��Հ�I�vWm��/��1���jzl�jK��_<97�=O�b������*�J��STCy:�W`��ŷM�
����U��j�7�s_K��Mu�Ts�K��Km�.;�ɫ�0X� ��k䙹å�C��3}�轪�N��+*�L!�7Iݻ��`�o��Ԇ�p����#c�9.�5V곪�j28I��ܭ'����:��{u���R͚�i��)c��ȝgM��v:��ѱjv���t�仂�g]��.�{���#��v�mpX9���V �o0�j�s�l�Vc�+��:�ު��j�/'�(6�I(�I�V7㷮��ҔmJ��o=:�t�se��'_W�)�C@���h ݿ���;	��Z�	Z�85�/IE�#j(e��P����	{N���J��%gJu���1��Ҩ!�p�)K��;7�y��FXް�Ȩ��\�����t������TaS#��=��:�ޫ�(��������QlD���(�{yɦ,0p�x��}Ƨ�X�E�ɺP��AN��ڂl��LS=�sy���4���T�^�m�jv�ѝ{ۥ��T�˞m0�y>�f�rb�N�-������X{�u��E*�/7��l�.�c�]]+���E�q����y��.Лv�n�L�#���K�^�rAB۽T�N8��Cc7Z�T`Q�[�s:�����y�۶6{=|��ΖɇC�LW&K3e���&h�CY�_����撚�����x��J�ژ;�~9/J�Ƥ�wj�*�ޖ-��u��}�@˫|�b饰t�s��Z�P�cb��<���\ޮκε����BZJjg�9L��]�Q��r�Z�T0�pw��.�}y�w�Gt���5I7����9F�:��˙�eWK���-���뜏1i��[�p$��w+���ǵ�-ސ�q�]�';��`��of�T��E�F�k[�Z�{�v\ڝ��)��Q���0b+_m�bݼ,��c���Ue+ʲ�c:&�r.�+�Y�y))u���D/�<��r*� l`D�2G*���[x�'�NX��E��&Ï��s+��p��܆s '�U��7�4�c��/��о �`�Rv=�	���^XQ=�}W}zz�^Qs�P�b��2�h�+��3	����.��Mjt�x�%.�:�D��qw{�����9�g�dx��<�WI�8��A��Y�D��,���-�Е�7�WZ��j*U�ڮ�U8P�ȉ]ʔ����w�ܮ�$�u=(��ᛔ��ֶ�BXqr�a�I87�²m��T����l�>�js�[f�/�/#��q��[�c��f��g銘�m�&�dC�@��,Đ�n�E2V�����u.zOi�ɫL���]��1��Z򪑊4^=�`�ܰ�8��^�VK��[7�٢�`��8�eP�$�k���,ZgNR���ݪ���56�8�ۜhnZ�Mv!r�4ޞq,��q��&C�Wfܜ�!q�S˅&��� �O����&txiC'v��z2�yE:z^ݚȖe:̈́��)u���[�1���ᙛ����7�V0G��Q��dV���NG:�q��^.�n��ƭ��Q���͎�L7)�"p��_Ѱ1�B�"_j����̏0s�Ҕ��\{Ĵ;v�̖����q�r1�)E��P���.�r�3y��v�g1P9��f�ζ�d�t�.�"�Yzf���y/��ۏ`�%�yXù�p
r햏d*h�ܘ�B��j�dH��6�`{d 3keA�%�[�`Y@N��g�v�����q��m�9�GJPw
�#U��Iw� �q�P�3o.��av�ɵ%��o3��FԱ�3a���u�P��Y$Aϯj�dRl��nhK�J7�Ř@��U:�U������unū'vG�̃4rK&.mT�rgRj�K�\�v����sWu��en�ĉy[�����3�ZY�-؏�.qE*е+n9-��1���k,��ͤ�;�;�� uw�B+�w������T�]�vn=�]��R	y]{�����&
qm�uUĞ�^p���o=
�%U5�,;�����`�,��apn���������7��8uL7+���O�U��Cl�����;Z�ԉ�����|0"edN�N��(b��{n�b��t`3��l�30N�h�o�\�_3فNt��3�+.���v��ס�A��y���5|kEN�S�(_ɱ-Y��5��X�ή��?�߯*h-i��xl��[�e\����w�:*Z+;oigE(��،Pwk�*�2�.uf^��q7������7z�]�x�Ӭ!�j��26��� �M��d�;-�Hx�B����T9�K�Wj��Vq�Aʴ�����m�i�V���qJS��]"����Sע��)�{ma�=�"�/�[���39ѫ��&�Ԧ�c��\q*W\z�uvAyq*'��r���}\1+��+p]��4�xx��.R>�����X2
sH�:��aQ��DYɣzX�Wsc�XN��M;��{Wj����&�z,rġ}�e`���;/�
�ۨ{Q����c���M��-��6�Xڻ�rf<�|q^KIL���.\���+a�!2n��9
¢��̷�,��b�Lr���J�)�P��_\�>yPz�8T+(�[p:��'#Z�co/FLp�|�Xk��HV�v�m�s��.�Q�<
�l2 ��j�r�.dC����2m�+���,��/ Ɯg����4�Ѹ��I����up�4gf|f�Lvz�9}0Q�0��5ۨ��].ѨA��9X�[���h��w�[}�[��u>�{fƲ��Hur��3��+��m���ksN>��N����JR7�;��Z�5���;�HEr��,�(���h�%��E��=x{�����Μso�cy������2�]Mo��HS{���w^��I���R>���o�vL|�b��s8�;���ኪ�/u!;!���wU���v�՚�'I$�I$��-�3Ɂ�^wH{��@b7=�<����r&@U�"�y^�/PFy^�K�Ʋ E[� �FCj�6!����y$Q��y˫W����w.
N�V��uJ>�Z�$��(��)�P�;�M���s�W=�{��O2��l[�H��}�紉2�@t{zݲ���9�^B��ny\���9:��Έ��ҁ� O+����hG�"uԩ�"ug��� T���i����RT��ya��6P�!�G N�@. 
��yة�Q��&�Z뺱y�h��Q�) �p"* �?�����A D�������?������b��~���������/��.�NJ��k?����u�0�L��P>9U�C���p]}��Sʿ<M�`����Wf�(�����Y��/�3K.���M䜷��r� �KƎU�Kb�ך�Yrť�*-}|�������V��1�W���rW�f�����3&��)p%h�՘����;�.7�cŴ�k����T�8:԰�;؟��+fLWc���(T�ν��K	P���.>�=��	�x ��u�n�a����mu�K�`����uT�G�cm-���ؚ���k�ǔn�;�n%b��k�h�t��2^�VM��:�q�Qu��Y�AF,��i�]N��ݒܜ�}�vF ҏ���g]\�V�R��h���|������Rc9�t�JnV��د
s:�`F�t�n�os��'4�% -j�P���{JocyI�J�_It�e��n�a̜�9;���R���YHb�&��,�EWK��v<=��:��`��XU��a��L�D,.a�ܖwy:�9[� �yfa6Z�k*��1O��r6|�UK��ܖ�x���̹or�S������'ɉS�2���`_:�_T��!asVWU�
WP��/��.�j�)��pGt�^^�[ܭ�G�\|z{q�]|u�u�]u�]tu�]u�]u��:뮺뮺��u�]uק]u�]u�\u�]u㮱�]u�]u��X뮺뮺�뮴뮺뮽��u�]u�_u�:뮺뮾1�]u�]u���]u�]zu�[u�]m�]u�^�u�]u㮺뎺�]u�]u��Zu�1�]u�]u�]u��]u�]u�]u֝u�]u׷]u�]u�]u��X뮺뮺��뮽��{���w��^��dÙ`E8��Kd�M
�O9_F�b�����f����[Ƴ�
8;�1��}qo�S�W(&��eJ��d�8������[��@��\�SM�5��^�k�7�����nd�����y�hvחR�M��6��Uuj����2un*ܽ�����i�hʚz5���]��::����]�Fn��
�d�q�V�X���n4��p�ՙ8�b�S�J�\��k\�x�F��1�p����Wvh�N��ZIK���k�\p椕fd��ٛ��GY7�m7ԟEbj=qۮ��ŦVP�l#���0 ڿA�/���zR�kre0�u�U99g�3'!�T��]����Wّ�.��t�F�\Xh�m��ٔe��ӫyu�zF�F�ǹ�3I�a��i`'�s7��sjؕ����m)pZ�A��B�%��g��.��({�x��X��(Qӛ}2���JP�6�P�@�w-���V�W�sVg4�������H)u�E��%�S�]H�:{���	����N�S9�7w�PhX#rU�2D�	�=�hT�-��-��T��[Yv�)rs2هj�)p�����>~^^/oo�����u�]u�]|u�:뮺뮾::�:뮺��G]u�]u�_c��뮼u�]q�]u�]u�]zu�]u�]u�^:뮺㮺�u�[u�]uק]u�]u�]u��]u�]u�]zu�:뮺�Ӯ��u�]q�]u׎��뮺�n�Ӯ��n�뮺��u�u�]c��뮺�㮺�n�뮺�뮺뎺뮼u�]u�]u�^:뮶뮺�N��N�뮺��vH93o,�GN�|��쉝�I%�*�ˋ`�����U�ksu)�M��U�l�&P8k5�ؼ{:�f��M��;�h��c���ڔ����H��),F1��n�,.�˘ݕS�[[
��
�����E]*Y&o%�{ ��Ap�]�,�U�s���-ռ0xz���]�%�U��W#դo80L�o�yKP]�aά|'y�ԅ�."-q���wE,!�s�ZyQ�:�I�5����w��b\��oL�c�`R�P�*��1�p {W^��c	q	�w1]�f��뎝�k��D�����k\���F45�]+��J�뱣q�\�t�FGMi��f�����Y����[8�W��U5���;')Gv�u�^0��gC�^4�hj9ۃ��
�䆵c
��n���w��z��}�&�jY�L����PMۼ�����(�Y���Ԛ9DF敆DM�M�q&]uR��m'�F��u�����ΦFK'�����`��]�����=�,�)A�4���f�B�\���'N�����A�����+�<�U���iм��n|���~�>^�]u㮺�n�뮺�뮺ۮ�뮽:뮶뮺�N��N�뮺�ۣ���뮶�ۮ�뮺�u�\u�]u�^�u��u�]uק]u�]u�]x뮺㮺뮼u�]q�]u�^:뮸뮺ۮ�뮽::뮺�N��n��N�뮎���u�]q�]u׎���:뮺�:뮺��]u�]zu�[u�]u�]{u֝u�]uק]u�]u�]u��]m�]u�^:뮇�y���X�H3U�CT�'oJ�|�ɯhn��Tj�K6��犺�v�*��K'-N��8�p<�yo!ݮ�\͚}�gM��'�r�S�{�Vu5]�,��r���g�>`n� ܒx�x^�y�JS�M�s�����j��|}�yi���7+����)U�����yX�k�SQK8�1S�f�nX��U;կ��&����b�Yn� V���;�Er�y��j�z�����'z��
|�)6G,��.���)�rdXfr����ݪ��p�p_<���뮌���%�������̠����� x�Y��uO��ܣ
R�vt[c���A����K_J�x�9O��촢���9D��G0��)�z�tj]�{&ժ�m�/J��UP:�Q�������;M�Ă�:��NR�'n@xT}��أ'[��*8ê�e��UwN	�L�ٵ�^�h�C�R�+�qaí��h�n���*�:o,NL��-+)�j�Ʊt>��]{����#�f.@���Գ:��m�6&:�r��[7>��Wi�ڽ8VU��7R��QS�X�N��]aG:�8���ۯo�N��n�뮺�Ӯ�ۮ�뮼u�]q�]u�^:뮸뮺뎺뮼u�Zu�]u�^�u�]u�^�u�]u�]u��u��]zu�]u��:뮺뮽��N�뮺뮾:�]u�]u׷]i�]u�^:뮸�u�]u�_u�]u��u�]u���]u�]zu�[u�:��N�뮺뮺��:뮺뮺룮�뮺뮺:뮺뮺룮�뮺믎��]u�]u��_	]򼫬���fVy���[ٸ���[�[!a�Y�h�e�u�;P6��&Q�D��M��U���;�(�N�f�U�#|�Xq�7σ��u%�i�V���8���6� ���z����n��r��r���8��Ѱ$6r�R��g��.hU��̭T����^�}�L��kp*���5�^��5KzXR��u�=�N�t{X��{��k�k��K����V'�E�E�hw����u\�������W���f���s1�^I���.�&BХKR:��5쭶-I�umɯ��b�"��u�I��^�ho;[����@�a)��a�e��7���J�����PD����ٔ+7���Lh�z�Uv]���n/a*`Gi0^�X*c�b�v7;������|<Dx
�H��V�����U��x�{"�����d 4�9b���O�2My�x{�A*F��Wӳ�ݥ�f*�aU�O��R����{oATB��R]�<��̋#� Ȳį\1�����k�`�����:�	%33N��!������{8�`��ϽU��u���7���ƘkH��W��{�ѨM�1�t��Uê�$���!B�̐F�,�R��i��<o�����Dްu[���}� ��#�v�ų��=���͎��M�f� �ˣ+�۱I��hr�x%\<=z+,9;"����rUGk_�b�!��K"�P2eP�Yj��eI��圪����
;�@ܮ���{�p5/�C�$�w|�NW��2ު���b��l'|�W����M��<<�  5o4�zͺ�u��V��R���!�N�_ew!�*�;�ݷ{e�-�՜��d���:�.���z��˨�'l^P�.��fR���L�ؓ;1wb�R�	ն&s��ʷ۬�k����/ �i#a�a�q��U�@d� �,{�nbi����}�S�Y�R��72�O��k;b�M���Ց�����ʪ����}i�ה,��<b��G''U�j:'�3ͦ*���{�=��lL�[Y�ʸ�ܶs�M�Q�|{��m��=���6�r��v��HK-V��K�,T{Tn!H�;���.~��E��Ȭ�k�w9*����w޾:��SB4��	t��zqꏞ%�ٞ�x]��yEu�*s!ZCl��y��[�k����V[rڠ$/@�7e��f�3�Y�9�����K���Y�p���46�:D�vQ�rd�)U��{^��iɦ�[��Lk��%#�k� �g�n�.��Z1+8�����M.q�mF�%3Hƻ2�������.߬E3(u���P���=����|�Uл�iu�kc6�&�y�^�#6C�mN��A�{�c2�h�%��J�
`��Vs���s�n��|�z����kX:�f��%�tq�9�=�5wZzN����9�g2��4��9�����F�
������E��_ =�!��[�ٴ7�ݎ�]4lU��+�Ş��%���H�����ǖi���o)B�Z�~�{09v�-����CW���r�QO����<�c�uz�����k��f�<<W'�Mkt8%��:�ts�mj$,}���)��Y�E%&��uL�V�t^pt�Aj��@WDvo�{lw
�ܸ�u��l!��[kܩ�Eھf .�b�̓���@{�Bf�]}1�IQl�a�U���K�g�FGdhrU13n�*V��|u�z���N�Ś�]d�Ԭ+�2s�E�̜�u��P�k��h��h��<1�X蠯UE\���0%�ʥ�-dU��VG ��w@^��#�dt)����v�R�*7��[�V� x����y#y]�S�Y��r�LP=�V�����̝8�p�w��AP�N�Ǎ�o��(9����3��.�8�y8G��WM��zWi�f�<7g�_t�n�����d��y�Guث� a^��ܧoqi��_����%�#Dj������1r7���r����ڒ
���Č~�W{qS�o9�T�.7y���*�M���!d��ɕ�5b��R讴u�˖sv��� ]; y=I���X���&�9G:�!5���)T�Ǡg_�|$j�Cު�|�y�=;4���3MܗBu<Ҋ̣��Z��F����4�YY�!���k��{#�����.K�ܗ�D�s����>�U>܃[�� �.=lk}�4�rJ:�\�ߖ��(0�X{{��;��z��T�����lR���r��A��vle�bA�nq�l����sr�6�R�pyzmfd7ϰ.Շ�CtV�p���5h,�x6���v�L�碄E=�v�z��>[�\�h��Vr9���i�\.�u��yWv)b�p`���;�G�#���l�L*�U׳��)Տz��"D>�ђ��h]���6!ڎC�*ѭ�r���/d��`v'�ڪ�e��Z�y�TQ�ZS�{tg<cR��Ń@���Ma=[]3�He8��f�zD�hӷ�D�B�vP[ێcA�S/d��X�s�ܹwV����!�Yþ �-gP���XdƦ�=���#���3�7SC5h=q��u��c�dܡo./gNn_�G����S�Sr��z�UqyY����y���ݨ�Ѻ���AF�Fj
���Z��I[���vJIڬ}إf�V SrK̷����f��ȅB�3�wv����^�e�Ȑ�yl*[���wt�l T�8�J���p��V�.��ٝde�O*�2��ڦ�k���b�N�f<���73��pP�3r#c�P��F�vH�[�R�V8PF�9}U��p\亼B'-�8%UT�%7BYS��P)��B�λ�>�uU|�H,�80����OړCǊ��U8��f���J��N��ԇ����a�g�[X���cS��h&̏�a\7+k+S�JDv]�\��;{�'Nfvk��,�W�&̝9d��]6U>���3[��*]�'���~*=�}L)��(�,�}0��T�5�}�:6h]��{��\�HJ�-;{�M]�Lǎ$0�ke�C#ٽT����lw�G/r`z2a��ה�]�I2�X3^T'�GZ��W2רg��[@��VVfW�0/�,wS�v]L�	�lΒ\����B���Xx��b-ӛ�A��"�GNKٳ"��^Nͬ��6�o
�2����r��[R�	�>�V�7k�1�e]�i��S���|�Z�ݾz�����[G4G^\�ht.���8�B6Y����݆�9����z�46�L\7;V����H>\�+�w\�}˒��֕��C�x%cz���`ч���[���ӹ˩3+9����l�M�㵒�X�[�BZ�
�H+�hv��s��,�Iͫ����7V���k��l��U�������#��(_�W!Q�o��զR�w�Cn�PE�~�T�a��4�u&j�a��UҭZO]6m��}�fQ[k�"i]Y ���%P�c"��w���w���av勋��'w;�y$őZ3F���>܌�r��j��ے�i�Y�h�ܾ�g�%H�kCC�X�9��5z�Z��EV�[c�`Z�mR�����zm�%=b'��ӜkqV<�.�*��a&�ܫ�z(%�*��lv�����+K�7"˹η�ih����s;C��꺑�~{7��2�ޮ��v)�qC,Gj��
���j�6�^��:���a���dW�r�k��2`W27j�ZslM�jyz�����]�ڮ������8m�\�����ި *�������������_�������CXT�¯��xd̪�e���u�����G�����P�Z���%F�hHn�%�$␒bN9	�$�������l"���!� |ED��7
(@I���&�'��d�IpI�Bm4�m6R-��
E��$��S�S*E@�m�c-H���A�������-DD�I���8\�#|B9��!�����=qዹ!����'��y b#�H�, cM�����@��������=�y�r����ҐI��A1��邍���A`�	
P��hTI�"cH�"Q)8�0�rq����M�HQDL)��J(�FJ��p�dH�Li��QbB"1��#�<Ͻ�.�/���=zsʽ��Q2)	,�R���M��<l�_���v��Yr���5�1�x����'�D��J��ٍ�n��̳!.��+e����L;.F*�jg�����j���s��W���UqW��W��[�H;�ы�a\:���9�G��ygl;0m�
�v�b�o�����=��3P�آ�I���{�T�R!���wL2�6.�S���N;��ԗ8B��ܶ�u�U��`ӷt��h%�6�9���}6r��yC���׉S!��-n�0��1%�i4�u8(-�A�.��I��lxI�lx{��[@�����8^�����3s"�]^ɦ��jaf�
��F�Y#o�QJ�wc�o�X��E��8�����Lb�g:(�-I�rV�0J�m��qQJ��v̶G�_m� |Ž�݀N�4N5����4�h�-l%���:��;�51k���X��X����_R[XOe%���l�ru���q���3�������M�l�ڑ9�Wu�p����-��}eWt�b���\V�]C����JI/�C6p5�ȩ�jaɤ�l�k1�c��NG]tݝ`�#*��֘*�^-g��.�33�wP\+s<!(���1�c��0�H�,�>���s�㻸�+���y��z��G,�s�8���/,AEم$I��p�T�����
$�i$[��Lb&�I��软w�o7�E���{�Y{�ݽr��n��);��n��($D�EF[bD�A1��)B�)RA,��!q��A���T���#.A\-�፨C�����D1���BZ���!%�r$_$]�tz�����<�G���<�Ͻ����r9�s��t���HH�I(K.ّ�ʍ��jpЧ{��S��-��z�1�d������tG��/���ǆq�Lc6��&Ȓ@�(�d�Q���M���A��q)p��z=���^O3���=r��Q�D��!%�l�G�<���z��^'=����8�s�����>_>��q{�qG(B1�"j	9���)Dd�8�A(b�6J��!�b��eY9@�["2ȍ�H��Q�9E@S��i�&1R&�	����;̧�]����M��,>�<ǟ����s�-����M�p��"&�f�-lA$��iH�H�F�r6���i�p"�Q�D�[I"��'گ>��y���U�����"%7!8�Q��������dI�À(4�di�`��؍�Hh!"(BCM��l��H�$G����'q��=�G�w�����,�c����kO���������p��!I$#ErD�M�,��R�a�l����?SJ���	�K����������"AE�"����===�:뮎�뮺��Ǐ;��҂+[:(p��QR�EQTo�*2��\y�ߦ�m��Ӯ�뮎�뮺��Ǐ:��P�g}+d��w9L��?t�r"�E	1P3�U@v�q���]u�G]u�]x��Ǐ�������f,}�Yr���S��d��	��n���{z}}}u�G]u�]x��Ǐ��}ﺐ]d��/aT�������B�w6w��Ǿ8�|�2|�����	EUCe�#����s$5�ay�=�>���F7w���Yj��Ң>d�S2o< R��!�ʒJ`�e�7!�
$�P�Qlnd�jN��5�G�q��'JV�e�Y(������l6�J�iAt�^�������R�fj�QST��`Ϋ�n���ӱ�L�#������rx�1s�����+�I�!@>!I�����;n�����Ԫ�j�.uiR�!��{U�+~G�����ԧ�d M!��p��BH�hc��|��N!'�Ǉ�&��N��	�X�QJ���&������;���	_>p����|��<��stX��$�;��kl�=y���jK�=�>8�=��q>���z�u��S˖��$�I$��&HL�I��-�N�|���`�6��n���yˮ����f���]mr����Hq�r�����f���s����keL�,��d �q��4\Rq�a����y��ۏEǸ<L.|�Z�$�6� ����NH�wQ�1��j��y}^�$�w�
A$p�
o�� +����������Ww-��:�/�\q���/q�^=�s����{9�s��x/����	��a�̍�B.�ޭi+,օ�{��"�R�[��,�ͣ�KC̏/#`�����%JǒU=�,^J�ּ1/T�^��eY/�]��H¼e�Dh���PM�;wQ.&y�ǥ3e��&��O�zA����*��dfA%�	Q����'V��J���XĲ��H��!Nh������w�a�A��ZT�ݹ1�ݕ�6tL��1��um�a�;���L���e�§>2O�n|~}r��ʠ�]��� ��\WF�bc2�ɬMn�D���R�>��m��-/��n6@�g�
��-}�ⶥ��H�t�`��z�L���-����4�/+�$����)Ejӊ58pf�i�8Qsfb6�3I2U]3�w�*n���#��|�q���N.�ӳ>5
q�/|3n�^'����\/�Ujb��7ߟf�k혷r�#J�����E��*��3�:�l�=TĻ�{EW��`�Ey����N��&_&ح����y�::��ǫ��]���F2�X)Z=%��b[Ċ�{��7���<<<<<+�lN'Ϣ�{��V3K'�8�],�u<~T%�׭Ϻ_�F��8r��'I^��6�N��������&ǅG}s��bYni|v������3��^��#t-#hE���1�>��Ƚ�ï��RIGe-ǵ�4�\}Pe���h�7�I*�<��Ul�b��\¼�J������bs�%� i�J��@�Ł��X�@1��u���u佢1��Cgk����])����y�~�Z��]�'2񯎧�m�m}�{N�h���V�R�x�lקcUadI�hi2��[v�2�j�]9��7�/f��r=M\���E��55��di��HJ<���Ժ��R-�u�.�<�q�6�'U�Ck`N�Q(�m i	,���2��8�2ET�f�QWYf����e2�A���U&$@�"M�+kZqV웙5�8U��Jl��mB�]Y��}�&'j�%}o
#��G�x�Fz<M��{$��գ��qb����0��]�r���p��!v�+7�ux�ytLrJ�7�)wU�1�c���\��겯�l��W�a�Q��=�ݛg��!=�瞙;KPGĭ�(>)L��k�b�R�)�]�1�N��2�R25'l��&�@���HKv�A��{;�+I�5���V3�/٤˯F����V�Ƈ���%ғ5�)nJ�TsvV�1u�����k��eф�[7�ӥ0�;�qD�Z�Ń�le�4�V̨�^�fG�m��N��-�3��8�U����0!m�*ֆͽT�H�ɜ�Y$��� �g�g5��cݲ���J��AĈ����a�m5��T��wA�j���ej��yϻ�7�l?/�QOɧ����e���:�d�#ڃ���9y��t���mi�	q@�kV������Q&����W�F{r�{�R�S6�zS����Ogr�Ai���w��j�U�z��)���n��h?���R��K>�pV�TqAm^������D����U�j:Ȟ�\�K�"�_�ry����00�n�\��{��ڝ�6N�\vަ�rĺ�n����ؾg�
'�i����%Vq��/hK��7f�U���aA��1�Tά��������"}�f
aV�ij}"���*�B6�},�aI�g��^����ײ%��gdZ��V%)�n��<�QE�5M�_���Y������l��e���u��7�,z���t�ԝ$3{*����ɇ.���û��m�d�r"��*q˥�5m�>��0����mj�8n�٫���|�A\:�}	�6=Q�wei�/;x��C&1ݞjt�Gu(�&u#��l5��"?hƸC�s�Yy��e	ؖ1�z����p���;$��3�4 ��e��c����ͨ���k���a��M���n޴^TsT)�5�6=^�5KÒ���Lw��oM�W�rL�;�x�b�Kb�����"h� @ݬ���0"w/�T<�ѹK1��#�L
�\6�RY��sLa;�P��|��w�v:U�1=�`|70H62������51��ʥ.f�2��w�TP}f��E#�m������"N�ڈ]���eu�w"��
�뻧J�2�\~�f�N��\V���ˉgi����U/F0#1��N��]��:<6ʪ!y{�C\��3�G�ǂ�މ�0:��坙i�`Y�Bٻ��3�P)�����W��J�ѱ���<��m�Ǩ�Ľ=�x���>Uӯ�d��ᅿ�;i��}�u��DV���J������܋��͉�ˢtGV���eþاj,��u��}Z�Ic���{J�E��N�Y�^k6 �7�(9�����x��<_��!G�&c��T���੬G �(w���i�����5�D/c������)��\�FV��{�;F���>]��^![��A�Uёv��;��d��	�$��W(�ūӆ��e��nB�l��Ri�F@̟I6
)�a�3���R���^�F ���eL�)�Q��9���G^�mږD��nouW��`�� �-�RR>@��5��������;�,.�Z�#L�\ZN�Q��N���ò	�즗�	�E9tC�ͫsf�{T
���g5�}�^4�H�j�����M�/�,YW��w)�YޘZБ��V,��?x#�;u��ehU�n2�aɚZ{Ս�Y�UXrX��+��co�����S����{OaOy��,+�������7��;{l[��������۽��+S�s�����h�q�����F�aC/]ܐd��!�h�y	f�W�d
Z���ET�>\�p�K(DN��K��q5虊L�X�F�pЈPnjI2B�lɩk�v�ùX��d�UU^���.�ǌ���TNɐ7�1���	�}$�8���j��2������5�c�w����e�LL�w�1X_����#���)9������W�߉%�0}�l�K�>���j����L�Ze$L��;����+ʥ�07o	������ƚj��d�.�"�y�)5;B�L葹01IE��22)��br��O��_4����(�,U��b
JsD�@͠	�w >�����|���I��Q.7�}���=��@[�^QV�␝�=	z�8#vo�b�_���/{5�ۗ�xY�U}�p:eY�TZ�1gKB���[���g9W��ʃ�r-���g`���Q�
�5W^Q��˜�	�Q�
�捎��EƖZ����ӏnnv�d��D��&;��>l�U���c1���~u�|�����{�^���-ڸ'�������~��&˵7vG�<�^t#�L�[�M� S@|�޵��oL�u%�N`���JcT!L#!��ǫGgK#^�H�l6F��$L��{r��|�f�uR�a���#n�Z���2�Fd�[�h��$��q`��5=]*[k0^�4;��F�
^��}�Z���o�	�F�l,/��9M��iY��TU�bM`��2H��& �ɫ����6\=�l�+v%Zӛ�Ī�pu�>]���Q�i�őހy�tv��Gu�.�o'��9�Lǐ5W������ Fl��E��ɍ�S��MgV�g^c݁ozhiٓk�z����[��(�j�R"�~�\��4�yd�[%�gO�'�3�2�N��}k�NVE�R��C.�vƽ���Q	Ո�y�UuW���{��[�+F�犫kr�и�DY�#�.o������-��>#]a�th�]��UA{���k=2��fl�I˦�vK]*�Y�|���x��1�H��6�κ����[�x7T!i��&dl��`��F��`�{����5rN�Y�؁���R^��l�ܑ�yMw��ޔ)Q���7�osr��&�@�����i��NO����x��٢����-���$ <;�p��Y������?�)�����;Dȓ�����}R*�s�:M�����|i���w�4�5Kٮiq$�Yzh�m��({�02�ilsƨ� �<�k��;lN��:�J|!�Bg�y�d�A% 	�-�a!t-� �0�]�2��=%� ?�<q�@�'7�+S*�l�
K��$ͺ�H���ʦfl��*Z��-�7s�F'�b�V+׉��M�e��Vd�V]k���Y���Qw@߫��ŁBS����纪���T,M�>N%��Qsɽ�pnd�][e@��?F�c|�]R;j�WԆACL�ب�n�m\�n�E�DG�(��_����w��.����Ƹ�˅c�8�K:�ڐ
ά�S	[��ۏz0��h�!�W�V�zo]�ԏ���c�'|��S:�@�3<�s��\�Ƶۓz�ΜOb�Y�;*��9��v�b�����Jt�Gϻ`�S�\�!{s�|�ˢ�$�S�隳K&a��5�,���b�U�VNnz5	ڊ�ճGsڦ����^����2�QնA�2/�  1�W�#=;K�LQ��7q-H����fm���Z��%0�2� N�;�ao�7�A���6��W��l�|�Q�A��($V�ǹɣ"�Q%�2.�<;�`���փ½ʰp2d��W�����YS�͸�º|�Zhϛ�y�@�6Y@�e��0�Ю��Vj����T�}�UzN�`��f��(@��1o/�,0Cb�zI�S�3*��4���n5{�|������P�8��b�W��ܯ`.�eh+e�dK��i{{�n��x5���x)��݆[�"_]�5�U�*6V,rM�^�]����}��/EP��~�����5��u�D�=�6!`78jٸ{c7,�R�2;���\��V��d�-��!�-Bx݇�������SWqP?� �����3�4gv7F�.Y)�<
�N��u�0�]6N3J���y�˸��8z�¨xU� [��=�˹�qA��d��ݾ�6a���x���h�=
�|��G���I���rLgu�B;�>삾\#w�W��"����CsV�ŽQ�wq"�i�i6F��-	$6v��N��B��T�>��FP�N�1�kegK���^�VvN��l�ω�,0L ��w��w(�CM�ZN	A����>�b�en�o�:}�����CF"i\�V��o�z-���/u�Y3Z�$�tݕw����R��ߧ�sf��yo٥] Vp�� ��9��{N�^�3/�_�yY���Y�k۶e�x�[�/�^vFG�H�- ��k���F �T�*-Efef�dj:t���'`�����}�E4���z���)5�����8�^��p��0�r�|y���	åG�>�y�Vd���b7j~�pF�\<�K�fE�@�j����k�E�P�Iv��	�.�:�Ff
��Y|�Ax:�>�ᓍj���]w�F�pt��u�yzX �sf0N����J
yػ�l7v�b�4�I��-b�N,����s������&�JbVAWh���L�s	��N�n�ζm:��8�ε41X�w�Fa��$ȣ
���z������!g�P@_%au��� ���.���Z�k�с��l5�¸V�'N5�l����,�#�/�m|�x����+�����˰d��3��w3��	N���N�o3(� 96]l(2^�),5g[��k�>z;f��e�mǴ��:�A.ts����T�]ۗ/
!�I�릡���M�g"H�/w���l�q<�70�jWew�"���s�)e��9�Wy|сNf�n��;2�Y��n�RS�AFՆ/}�K����ges�:��!�7�<t��ф[9ٵ�:8Pu��\��ev��E9��=rN��-$>��T:���.������ם��5�'�󰢼�M^A��盇G>�Л��7f�v!�G��K1���s�'�;��èEB���JPp;���vl�YNV�6�J���0ă���v��R.j�DLTAĉ$8[e5TI��*h�BJ�;�&�/��w��8H'���q��ų̌�q�2���Klg1j����'$X�g�As�U��H~|��̻%>o�Z�,�y륚�I�ٱ����Q�w�S{�-J؉�}��k��(M��e�^�\��t��M������\��zm�rNWq�V�`\�7�&h�{�'��t)k}��K�7G�R�@�A���4ȇw �'�:��W[ܷ�gsά�:.$�f+����B�43�Tcj��"f�I�}p����=.xp��p��ʬ0	�&�+���S�]�6��l�z���v�˒�J��1W�׸u!Rޛ�>;;��C(��)I#����&Ĵ�8M`��:RT�U�������w��И���=�wz�U�F�(���<�vZ���!���w�f�)X��McB�<p*�Qw��/Sڪ�Ӎ�����hZ��q�I�{�u�ۣw`�WK���l�uus��2������+�9�:�G����wV��g(q�^Zշq��8�<���]q�ݝ�gs5�Y���_3:N��AF��
z���y����O��u��8
���w7��(� ټ71�à����Ρ�lZ ��G�Z] {�ӷI��B���S#^P$�v �y�&UNI:$�N�DhЪ�"/�T�	+$�[��7�==�:��룮��8�:����yʿ�$.ǝ �N|�nw�q
*���sG!������=>�������뮺�8����H���.G��X�i�^���K痡@Sul����o^���������믣��뮸�8���G۱�%�)�r"g#��7�`@�E���\�c�|x��x�ۯ����������8�>����w��h�C�^����UQ� �SJ����K����$�g.9���(J+�rNR*E
�\���Q̐�q��7��UW�^��q�7 �XYP]�s�쨞b����{��eЍ
}W"��P/�;
NS�G2Q�u�Cȏ��g�C�E���]�c!Ȼ�iY��E�=s;��2y����:�$N�t����4��A{�	�F�C�c��Ў�Є�Wxq�$���a�U�(C��jJ�.{�v��OQظ���ۗ��/�xyxz�i��Ji��6���}�=�U@��j�~���ͼ������d#c�}պ�iR�[��c����%�VcmSSy���������6)����%������|�)�?�~����Oo̟
�T��r���� 5�Om�M� 7�g�>����s��a�<����pT�^}N4^�"��<�o	�V"µ���Z�q��<9ry��-=Ƨg	@0�{�)'΅�e�X^���9S������#g�h@�Rل%O�{Q�9�,��>z����c|'��J,u)����|>ug�|��~b���27��Y�z��w>>���D$"@���H�I	���ֲ��{ɱ��|�|t�i�=��z���<����XkPW��+I����_!tm`�$=<��y��p����p9S�_��%�>צ���t�n�q����"�����Z�$�BT��{��H��L��\]#��z���~��&)1��}}�l/��O���	�"�a�z����b���DҘ�����,8hP=�;�������t�n[��INs��� �eW%�&���5���x�οJ"����������<�G�W+��lg���txK9��*|*�����*���\�� ���Ȫ��;��V�؈a�YMe�Ṅ���$�.�i�Z���k�����@=Պ"��y:!{�ծ��[�Z�� Ǉ�j㸓}����Bz�bͳ��+����(s��M4�M4�SM����=��ȵ����/����i<�
��>M'�VQ}��ց��[�F�d�����m�͙ mBu�D��-��L��Nۋ7�4��/�~�1���1s<��c�]ً������sX{�����<+�GK����+�s.
�V�:{֞�o��O�j~喼�z5��A�|

��6���ݻ8������-������K�|�}#��G��h��0�-h������&�L"�8���Cs5�y��G�����=�{C�:Q}a����h|}��	�VE�Ce��a�4���t�R���-����xy`p��c�>�;��y�8����8��Pj��y�c�V�଀}����F�_MgL�_7�<��~� �t�0况WT��.t	����
 ң�S�\J��Ԋ�������{��֟�����\����\�y0i�m��x[:S@T�>|���r����>�d\�)@����"��{��a���e����|��_E���K�R�g�Л��nb����>�à_����^��Cγ��.� ����O��?8o����81��e
Pf��S{dr-�^���?_T�3'�g<�/{m��T
l%Vq�X�q��LM��%�w-�Y��M]�랭�U�É�͡� i�ʕ����`��k*9��T8%�b�N"�[�G	V�H��M��z&��謱:�,.]{��J~�����yy ���ۺ�w���\�4w�ԩ��ٱk��;�e*ŢL��xXf��4����V��V��p�qE#��8��� V��-�n���o�8�=
����P�"�@��~`7^��Juk�xuGO/t���o&n����*{o����z��~��x�@X�{�F��Xzup_������{��UG.�{�%,0�P �m7��^�,��r��O�������_s���@#^z}�[��h�4��K���ɌGW���� ��[w?�7ax���f�� �WU��\@��zQ������,v��خO�x{�[�vc��0��<�i񽌙]?��=����H����}Ʊ���6�kb'S>*�St���p &�/�� l��y�(�>�`m-��^�5����괸xzA����ͧ����{���)��oР��0�gՓy�ws�p�3�q������'�����nu���tszR�ڜ�G���8��>��'���g�|�D��৤|g/ޜӱ)��
�Z���*�fQS�Q{��!�K��BR�|:}��5Q�>��+�	Ӂ����	�<������	��O�<=�	��Utݖ|D����@�^�P!ly��ʁ�l��\	w�ą��|��+"��d}6��K�)XH��hO�a�,��<���?7+�����΋�5}����ϭ��ُs؄��	�q��6�W�d�_:�>#A�H�TQ��	���m�cu:7zӓ���8;3{K��̌c�|d�e���s�����Û��u&*��M4�M/���ƶбXJ+��faml��>�@oE���� `���'I��1����%��k�f1�=�/3�d�p#����3���Lج`i��i���oV�S�zK��ķ^骦��Y����/:�)�x=�hGw+���~��d�Zc}7���P��A5
�=
�{�X�u�E3�Az|1�yx�\�������>-H;�p���x?��oƒ��Ū���rs8 ˃���T-P�f
VQ��Y����|	H����=dF����j�dܞ5�,��Jr��RXsW�����F�c׵�)J�p!e� =�ʌx�+��Fw�C�xݿeNh3��+�V3���>��p:�l7�������`8��o
u�Q�a� ʱIN��GM������*��\̝���8����ų�K�E��.Lb��x	����MN��;�ݢn,�k���x!����7�2�D�<�L->�Ж�s�ЙPW�����e���������tI�:��?�����hD�0�_�	���/���OP]c�t���%��Wä�ߜ�y����}i�k9�8XF]�6�0�W�efn����M�n�9�me�k�S��P�$�����)�ٕ���u����T"u�;�ʬ7����ש��ڳ�k��Gۜ����w��M4�SM4�@�y�w�H[�P�0��5�;�<�L�-�vF�}շ��c������[^��.z����]�i��`�θ� 
k�"���_�ߒ'�-�r���AZNk^,��:u��?��}.�)�t���mȐY�0̤�h�;z���X��W���Q�I�a�����,ӝ�,;y�u�v]�H� կ���ݡ��CM�m��I�-#���l��������)%-]��ʟj��
;��g.�D��S1��4.��BX/��ӏ�j������"��iyVK��+�:'3��׏�Uj�c'�$���F䀘N�HCL?��<6e��;m��곾�ݲ<>��^��f !N��{�x�����#��)@<��!u��!����j2��YE�OL-������y��W�6E1и,�xH~���	��y�H����檗d��I^�=���{���|S@��\B����tާ����X9z���p �n��C��E��\�^nm���kOs3��%�'à���q'`	d���4�b{�Sz���Z�ɭ��E=���Xt����׍����竣Ȯ��W~[b�����eۗ#�*��C�R�y�65g���Ͼ�Y�\�6R�2*^oc��e;N�,c*\�]�T 7:����7vC��WU���#%�YwK����d�fo){��\ް�%�M4�M4�M5G��g:�z�ʼ�.#� �\O������u�}�+��H^��wus[9��d��2�Θ�t�ٓ]�w�<�{���[0��b�g�7\M����p4�#X�k��ú� ^f�ɘ�]�k:�U��3>m����ʟ��Ǉ��;ί\����@��+���rܟR���oU")���}xWE���Cu�yA��n���>>?A}\��k���{�=�M>�����=�Be.�����(ox�@|:���X�B��/���Ԉ��vc��yl��k�<�
���MU�y��U,ph��uϣ��N2�[��1ټ��s�K�t��ا�ٓj�w�ɿYI6��T��0�.���>��x2��I�0=* mk��k4;��
���.�-.�6V=����b*�q��g��R��$�>�2|���.���|5f�H�/�:.�����s������令�����}lxi���&S�} #��)7�����YřN	��w�ɛ-[���}=��0��\a�N�ƜTV���!b�������~uy u3����%��t.�zM�ؓL5yP*��u�=4,�<>.tߗ++(�쩚�7�B=�ۖ+��G���s!�+�3�R�C{K��ۜ�J�%nNK�s��v�t�J�2�;������:�7�N�ʮ��Zi���i�qǃ��D�{>r����=d]��}W�%��v��H��=���/Bd�ݜ�BGs�x:|/���|�E�B���tٟ/�R��*���X���om��2x�\zl��� ��4�J��[w��?��[^�V�������Xkֱe}��
J�
a�^�w����܈�W3����0�硍�\��� Q��A�\C&�)N3҃n/=1R�,�I���z�1�k(��@x�q$<c������=�K�l�tq�'���<��h�
�]\�����Hރ��+9J��v�M4ӾJ��|5t�����[^�~oe�".5�m�����t���#�o"W,�ϋ�Mh�<��pz:@��sf� W�_43��~mi�B�����\�|y��oY�<�8Mw�e>��Iz��(9�/A���'2�C{ۘ}�O����̹ۛv���~����<���s�ǽ��M���X^r2��=D�x.,yW4.���"��'(�"��!�zuuA�k�]��5=\�y�P����X��7�y����:Y����9��p�]��A���YX�5.�0~�ݎK�u �Ƨ�zK
[�~�W�@k	=��iw�s�<nZ�\ʭ�y�э�Q��t��S'y�f��䕫�Mգba��A�s�v�CU������"d��^�]�Vj�)X�^옸�C�P�T�Ӹ�)���)���2Aw�:��zvwrv���M4�M4�I{����ߗ��� �ߕ�⇀�]:����o�k�w�a;^�;�;�ҵ���t_��zۺ��V^k��<�@�om�� 8AǙ��*@�� � �]��~�ҹ�>Kڭ�{=MUWu��]��x�ʞ&�&f�2$�	���2�k��{C�0}��)�ܛ��.|fl��ێ�ܲ�v���.�ԕG�\���������v��� Z )���^�訿Gq�!�p$C�{aO|�ۏ�4;v�7l�3p8�z���B�L]�������%�{8M�{^)�xh��め(�,�}���j�ρή<~��إqQ�-Y��33��m��0��dy�����j3s�{ʡ�����g`̽:���T��2 ,hV��5�{��W���c���}�;��a+�w*��\��w�yc��O�j����c�s�6>^(��ӊ��u1��>%� ���9)U��d�~'��Wk�����oc[M<5Ӂl�ث�B�n�o��>�kԧs�H�w��T�bS��)L|��=]^o�1P경\g�Xx�>Z����o�س���/��Xt+����.�=ۄ<�kl�����r��wujM���f���c���ҫ���۷�M�cc�c��"p�?���U�P-լ<pΪ��A�-��ݷ9bWB���B�����z�wԻ`�����~zi)���h)��L�M������	��}��oA�E͆ؖ-�����_����K]��w�up1������5�y�����7�[ų���s
F�X� ���v���s�
{`(;�/n�.��T7*z�t��<g�&<�8�#Û�Q��)>IE��p$8�C�z�]�����\vMwo�sH�ҘW���>�'.���=������a-�-�,�noM�e�6�,;:���tlb�DK4��)���=k�|�L@ROq��ӓ��y������`C�o��[ɧ��z�Jx<h������xa[�*=��txB���:��v�A_k�`|��=^049i�,B�uKR�Ĕ�r˄ oԼ��S�gӮ��@mnD���03��A�`"P�Na�/�o;�Ϸs�D�<�Z5��G��@�˧�@gF'�gz�H��\�W ���;��"�yp��C�_O>����ڴD"���h]�pN9�}Mqa���@�:�!̯{�Pw
1���Mr��Fnz�zTU�MZ���<i����Mw�0xG�]>��j}��H���H�;<�A5>A���#��E�x�fn�9+�=6C�;%JT{t�.�k�wR�Oc@�^k���������ۑ��H�T�WVX��t���������d�g�f��K�2���^k���﮷�\�>gq�ou襹g�j<�gX5��y�������W��j�m�r�۸BI!	 ��ל����;�w�gP���3���0,?o h1��a[�u�/,�/s8Tڱ��4��p�� �^X7��P}��g9񩝼�b�v��Q�����~�u���������Q��O���W^N�MB�Jz�Q��0���x�F=vn��G�X������3#me��2�	���\k9�׆���J��=���*���j���+<G��T�����7�gJ�C�gO�Ls���E@�Θǌ ��]j��ޠ�}�͞���8��vf�r��',pS>�2_8�1��O݂5����+���A���yy6QLP0���N3]54���(i&�::P=�'��]^X��]��x7���c��9cϼ3�{�4z-|}��f�خ3&5^��w�N'��R-Ov�#p�r��p���x,>?9�[L����ߟ_�)��7o+�x"�8>��pt�y(%�c?�gw�{`�������p9�G����:����Þc�YH���[���aK��EX�i��]�T��'�ȑh�9�V~�r��_�k�5������_W<�S/���W�y��ފECA��S�J$�#���8�]ZԎ���v��ed*�f�5��G���RV�N=�&��������SJ��u��f�̹uwx�\��"�}p�ۼ�Ċ�t�Qd�/0(R3sks�ԔG[����gD�[����bs�~Q ��w*��� mV�P����z+�Q��9o*�';8"G)�:��a����Y��:�g�*�*,���v+^�L��S1�xtpż�A�0���&�]nv7\s��G�r�f�6�i��=z����X��\�7HY�wY$]����ݗ��xq5��s��z&5�5�y�G�*<�Q��cJ+Qw�6��!]�:�N�Kj遚���DFu�edO�-�%�9ڍ������ށp*.��n��W��T�&gm|�����ʒ�=c3��r|j�lS��b����vfB�����f҇���KM&���8��aw+ayf"�Փ��S�p��0n�7w,^V���<.flyf%�A��B�D{�2N�j�	NKOPPr%�H����]��Ka.��C�+���:�zX�҄�l"U�����k&� �����v��rD�.�,P��U�"�&<��j�|y�2�%�Ɉ%h�Bl�E��>5B��(�dאH"Q�Z����TqJ2�s�A��(떙D
�{��rZ/-�G�P���RU�@�_�!ܛ+u����S��'�P�Mi%D�1T�v�0BW�Df�ۙ���zC����{͉9)c4eOrb`�{�����/�e�K�XE���1�1:��'��N��	.�A�e�Ե�]t7��X��`#�G�wv�a<t��]Z�ç��9�(y�{û��Qeof��i�N�d���K��R��(K���:˗�]b�ۄ%t��Z��U��[U٨�=��E��a|��6v�]�<Yy�Ѓ�J��Y�V�#e-��y2�)��*Xl�v�vԾ�"���J8t4��:��;��ԭr��m��.J�gr�#j�VRQ�I�I�dx]�\[�MMU*��7�ű���ݮ)#��iŦ^L�� K���P�%R���a�O_�t������ɖ@�T��\��5�ñ��u}i�²�oS�՝lr�|��H�t����u�8>���d���_
����u�H8ƨ][�d��є+�S�E�͑A��V���Q��b�]��+��{��)�e8����.��m�L��Yl̣�������0Z�;����(���¹q�̽�̴��̈́Kս�h��}}�C-�K#�:�)\y�w*p�/;VN̝���r	�s3�C���w�����7��˗�	�AeZ"BTӔ$~��I�� �{y�L�u�6��Ӯ�����>������8���� ��%B'�S{��]��]�۞T˕���m�:�㮽��____^�q�w���T	g.�g]ZDMΜ�#\�C$����z�G�'��m��zzu�]{u�:믯�O<q�����t�l�D*J�HH��2�����B��F*SU�Ɯiǧ]u�^�u��믯O?7������}��T&�������/F9�qa@�D�b�ܪ�{�:���9\��e*�-
���#%(�M�;�g�9��(�-�9¬�0(��#9�XBO��U�xӦ��݄t��u
j�� (sV]	9vQ�d����ܔZw;s���q3��f��Q��J�AH���&*ӥ9J���	��E�O|�����;�I����.g����s��ק�.���#�6�E$Jb%$!�*6dj9I@Z��F�D	d�d��#"�VԆa�x�\��-C�9Nǂ�Ӽ�`��K4�,�,�k=%�+��7Y���.+�{�c�rrH�2)B8�2�Yo<���^����-�{�Ğ�ǻ��g�={�z���g�y����ܳ^��#�뻄��ב��w�:��{���N��y�Ce\I3��2Gi�.2$��j��N��aa���|<{�'$JF�2iR�$pBԄ�E��]�G�G���m���m�-��[A� �����[��u&\�߼��U��q�Wn��k��2N멵�'r��+6��օ��Ҥ��p��j��:����.3��M�$�U�����4��^���l�H�Ϭ3���=��]3�m���q���;���pJ�+6��0n�!�=��L��$�̗�w&|2n;�m%l,��{^J�9.ĲZE�=[SK
朽�����y�ύ��~�P���}(��P����،���c�@)<ۯ%��Cx��Eq�}5�|/�OH�$1��y:耽2����[�<:��Z��XW���r`|�s�{�����}##;�09�H���~�!�w�Ȉj�~U�-=��&�k>R�&�������]���l�ڪ�n���'�����޺�rqWP�	�  �2�)�{�gNZ]��
/͑5�2K��4�a�y���}��N"�v�S����0[ ���Ni�S��U�	N����ɼ��h���@��מ����|lb�9��H_*�랔s��B`{|���F� 9RB�+2���r�+��;��?�̌b�CE!g}�=�=O���d#�3x�k�)��%q�nc5�tYff7�B������`��> =���g�a���C�"1 �߯���u�Rs.:E���_R3�τa��k
�B��דxT����s��LK3D�}`��P
>���.�:����t��k�2�"�VvgG�;b��������Fs�;fvUv������0 O���1����m����m�	 9���}����߃�L�0/�ѽ��N��
1=;��Gq+'��k����@�w��F���V��Ʉ����nc�׉�n.�5�ݩ�y5?�g�D�f�	cVD�G�Ǩ�$]��ˀ������p������~e�W�z�5y�}u���.{��L���xw<;��2l T�Q�>%5t��+�`�>qM�`�����T��3q�����FKt�H�S�k[�e��w32�쿀�@�^� z�`�s�Ln`c������ŧ��#?7�k���{i����_V��Q:h� <����Wm�xb���Ewg	�|/���	�e�0����5�D���ݣ9��B��fxV�俄g{M�_���}�����&:���Z퉆d��uSskm��n\x&f[�m�۱)���y�I@Z�Y�Hft��-�k�ڜ��j؛�wx�:PM��G���ݼ��)B��cuW|���7�/�����:� ��&��c]/��G/��m���{��>�'�����2՚��@Qbe���҇��o���]kI����c<�.�il3%�9�n�Y�r��+�O�т^�3�	=�	μ߯b�uع$���n��G;��	�Y�"ǬxB��� ��b��3�9�|��e�����p��z�:���ez�z��g"R�0�gG=��멽8��ޟ���m�-���m�P`<�< qJ��WMr�0S)�yg��!�/|�v�f�W{N
/�b��@�`��]5}�Ofp��޶
���]0-��]��\|e���c\_�ۺ����C���쮮�=3�� |����`�V�s�	.�3,����^>!�+�r}�6�4>�+�֡P����ɱ�� �N�=Ù ���v�3uNY~U`+I�����'{g\�a�y��i�zP�����6�:L�v������㿎����)�7����}�C���i%�$�	�_�>n�|�/u�̜�FCpa�#�-�1�!�vǁ�w$�hO���S�� �)��j��[�����LcC���F{x(�O��O��a$Dxkd�dJ���}j �����VS�#�7<���AB-4��7������H|��D�����37�[�xBөg����򾇖�/��U�e��7T>8�T�6{s�k�lO5P!�-���~���K�l��*��+ҫH�(y�~���gouLO����l�i���L_e%�����͔���I�y�FŰ���`��H��ߐѾS���̖�n�/o
4(J��jً���=:���+�c�R*�����Z���n�5��*US�ݺ���s��냤8u�ofp1�%���N���V��q5��2���.ڝ�fn��ŵ��v0�����~�����lB�m�m���=���<�f{���S S*�2@׌�M�)8fi�������,tk�L�U�I�0y��ў��惘��V�.�rC6M��K?��C�dB|�a������Rw���{2F��!@+����{�{�F�<�s��|n�>�sL�ِ��1�`��g�]�+)��2��h�H&���Nz<Z���$���A�l�?y�:\�_o`�􈓓��8�_uZ�S!]g]�N��J?{�k�	k��'���(�z����qoq|�`K�ȧ���`�ڔ:��d�<�ǇF��ԑ��>8���e}86
<E�B���p����{�1]����������H�pp���|�����xDu^ %�%�OV��~�R|�:[o�� ����O��,��^c#Z-�0�Hݒ�޶��OZK���W,��X@�VW�wN�D���2iegQ�<��^"��]�&��&������@.��]/.�M������;�������W�:�\?7�Y��҇��;�� �Eޡ�s�ڏ@\w�
�;ڝZ�+
��xk���+-�8��ݺ�а`[Oa>ݮz��ƔLc����o8�L�T weHD �%�w]�!��w�<<6��睦0���,�����ރ%u��������
��{YA��:���|�eY�"p�x�؁q#m� [m��\�m��A$�q�~3�+9��M�7��)�dU֒�i�f��o���<1+Oe-�v���5Y���+2!�Y��k�#��3�c͹�ʶ�9@��|�<�a�@� ��6`��M5����'�.��k���mf��-����?�v7H-=��my�� 2�l860΃bݮ����2!3k�BƲ���w�M� uGc����K��ff��<��� ��
��?bd 4���G�Ͻ������<�'�ȞsBc�Y>G5z��v�?�a��Hu�W�]φ�����k0f3����'�"�K�����}���I�x=��h�gɐ:s ��Շ>�����]'��c��y.���2#�m��=���ri��{J������p���(�������A�~�Ӱ��D�TlA뫞��xq宛�>�:`�FTd��`|�Kֶ��wP���R�e��%iʉ�g���x�k�PͭI�� ���Ϲ��B�k�s�ޝqߕ��~]��w��P���<��S2���+���!�>G=)ޒ���oC;�<�,�X
�%����;h���L&���k��9�^�K��⨽_�*�}e���z��z��005$��6��<-�<���(�Æ���Bm����C�۾�.�(}+��N�.�Nd�D�˂Vt��tr���6�66���\�	���>���Ă�ٳ��N:|>;k��_Y#]�c<��{�M%X�2gSQ��1�9��{�Ԙ'��7;jUw��{�����Km��m��."F�m .*����^��~��nC�= {��F�B?�w�`Q�5|h�-upiK�_��:sN�}�[}��
�X�����G���>\4���7�T"1�����_�>6��D���GS�B|���{��ή��n�F�����vԤ��=��<c��.��Vx4D(����y}��/5P��G��Ҝ����g��OOypZ�6���<|�9�<��Dg�i��23v�6\�Kݖ�Nyg�S� �sl܁�<��Y����j���"����$}:i���*�y~�0L^��=�{8`;��*���s���`8��1��ڞ�3E�f��!ᒂV�"ϵ\�VTxnU������,��]��>_P�W\~�!x�kX�˞��2��v�㠎Mo!�U.������_��@� �[ɨK�~� �ϧS��OV��³�N�7�E�r�E�o�����N��ɭ���𧤬���d��p���_�xk��i�'���<��Ω�OYq���Z[ˎ���g����uQ���G/�"H=`i�Y�'�*i�|~{&r����ν>�%��~I���~[[�}X̲qr��j��ve�W��k��Lj��z��1�F˿��xg�M��@��ӪQ�-F9��w�>˅lY{؅�\��#�f���X⾨{Bv{y�:��%�� �G_��. 1�� Km���m�T." �F
��,�'^��7�o>���=�d�j������(߻��4��<�>�����#�O�*@�r�m�2!�7	9��_��噏
���ؒ�2����h����t�Hח~�Fv��\.zs ��<�]��z ��{aB*-���!r�+-�j�ߘ������$�K'�Ὅ 2����s�}5WW��_50�<�'�>bJ�k�L�P���^� �Y	�oT�!�<hD��ө�&�u��߯�r^��I>N���qq��K+�Xh�����y�r��L��8(��C1h62�Z��~]ٸ����P��������'>�3���R�X�1e���8�~��S���Ə3XM�e���A�w�X�z_t🕿��'�Y���>�F�VQ~�
e�]�Kw���綟����/�y7�n�kFo��iv%g�.�og䠤���{�+�r���Y��>��k�US��u��=߼7�����a���ޘ�P4M@��{�'9�1-���Su{��`��\5�C{�n)4DM���6k�0\S\:ol�!�q�*	p$)�2~aHԢ�� Suv�M0C�mU�����үU[��d�Tsn�f�Ԫ�&�p�e��u,46��n�uH�ʭ�}0"�^G�$Q򧽹1�|�iӋ�����f�A�sB�MR칷u�n�����)��4ⷈ����H��jm��[m���m���$QS��y���}�_�{��?*�yWT�|wm��o�<��-��D��o&�|N�Q|嚘'v�qYʒ�]o�j�};�J=_� ��w��p�Ad!�=�h�Q^<R��:m����nٔ�Uդ���d���JW�2�`�"�~�����O;��ùJ�D{^�S��z5��H!�\�Ķv+���O�.��^�rK��f��� �᧥s�t$�]=�@�L��@�k��:0`5?D��#B�O9P�����y3k�w�ם�=z�M��R2cbr=��TϘ ����W�	
}*1�i�к�t�ⵉp����z�v-e�K�8n	����'�P>,����t��C�<h^���ɱg��^�~�P�$�r5:3�üX}o��Lg�V'�}n�>ۚ`�v9=Do?+���69rΌ7�9��	�]��̗��)�a�������EV��8dM�����P]Jry6F�\�:a�#Sႆ��q7�~U�Z����'|�ta�0V����O������i��A���6���<���,$w�#CW<�M�o��\>���{eٳ���E��@[/���ھ�
��!s���ƅq�ژ�!RM.qڞ��0�^��"b�ʢkr�[Lm
��Ȭ���8O3�U{�{�!\��#o�n�F��q��1�]XA3�̝tTȶG�֐�z1����{u����f^����� �o�j%�6�`�pR6�b�m�� �T�@�Z����zT�<�
���zz����v���h������d�;y+yjS����)����V%,������(�~�������C��w=L�z�Jr�ɭ�� ^=[ռ'ٚ��rw��:��n^���x�7����[�dkF�F�Y'�.SM�=>�^�8�͝�w�.p뮓z���[;zۼ_]�'�xN����fj����^>�/O�%��t�Ssy�S۷65K��h�t��Y"N@רk����\���W"ѩ�֓���o&t����U��)���{r�Y��;8gwgfgvp����	<
���Oi۽�8�:썱��>��A� �G�`K��_�{V�Ÿ[�������"����Xy��C��J��7ϔ{�����9�aS�N�CnG��]TҬ]ŀ|^����)���V� z*����;�A��O���u��ν�N���|����1����1�-�#$����p��X��s�
�FVŻ�v1�Ё������:� ���M�����|y��]sЗ��Q�j��ķ�H׌nOi��ۓ�fUe�ʪ�ؽ� ߗ�sܪv�"�H�k�TG�/�3�y���Db$�LvFֺ:�r����7�v�ʂ�]Ƅ��u�Hq�l�T�K�Y{���G8���ȍ���C�%��2<��>���D//��*Sx;�������
��A/:�uٺ���h��J��vؓ�:�9�������QK}~lm��Km���1��U����=����f�pe��֙�O��P!�`@iG���:��z<wR)�P
�۹�<w�xxw]r����}�H�J��K��n ү}�c�� /(k�Gri8/Q�v�Ul<;?;V�O���0Kd
�o��3|��fyXꖀ�M��F�;k6v����ȑ����>F7s��zf��ށι��A|�����$d4�3l�lgN�|vۜ�N�;�䞗~�c����P�H{i����
3��A��޿X��]լ�L��.[�N�d��Y�z������J����0)��T���|h��1�iT��Srw|�8�x�.'��ozz�
jœ���Z��M��?���Lw<�pDz�[F���L �{OS~s����"�t�8���a nE�q���ۛ�ò��B�=��7��;���������aN���l�[��Ҕ�1eٮ�X́co�5���)c�8��tI�i������e����)蘦����$���������ݨ�:�y�<��f�|�כ� �m�vмô1�J7]��U�δ֊�}����&c�V𮍑�_��Wd�L���8��0�/���\+��ugr!D�1'�)�12��ǹ;��`3��i�釫u[v7�[�7���"
�T�',w|k�6�r�m�`��\˱��䧞C�\
�{,�p����:��Q���&���V�����<47K��:r5��$��5��5|�h�35�]:4�R�fn�u��F�n6�2;S��k�����ܙNf������E=�z�t�6�Z�����E(z;w٭І�ʉ��-�z:��ubI��g1}Y.v-[���b��XƱc�S�7+�M)R�5w�}��M��"
نq�&��1�[ӆn�9L�u=�&i<��d�w��Fu9zb�b{�7��`��m��.�r�v�S8q�驽3cF��U�L˓���kR'���I�T��>�t:�#��B=b-��B�[T�i�;-���7�����G:f㻭UkG�@�=����Ys�ne���sV&3�Qf+�u[J�<[�9�9�7ֵ�oT,[���7�C��ԧ��])UR�ͧ���k-�<-�zy4�~ƺ�ea�r�M��I�A��|���0q���2��j����O�"���ƻ#���^A:L�h�G��*��H�_����|������*"H��Fs˷vkH�Ek����f��2�N��o"GMc@.��i��I���K�צ��714@�����,3��l��sާ�~H�ﴓێ�!�V�P���IwѽD����W��"�����F�R,���9u��5(��3�c���+�*���кi#=%�e������s�`�hWd��f=�.���X}�T��ն{"y��r�q��Q]ՈMƹ]�N��3�UL0_Vls��b�4��U"��B��ӻ�.q�6��L˻�0#���p9�U��x���'`����u'|.�̭{ų�e����YF�����5�f�auֱ�u��;���;��a�f`��w���Z��*��U��!�/���ea���+88Vb=p����u\��,���<�-u�5{.�p���w�7NV�aw3�������/D����p,��U&�O��v�Ė�F�:宅�X��OCa�b>��d�r>z��۠�P}Y����l�X����G׻�U)��j�CY�H1-�/�ug�<����Z޹��P\Wu��`��vV]�1��bu�ɚB-u@΅�`�0tus5	l���r�lB0ѻ��)|��5ћW=}�X�-�5�����G�qO,��iI}����._�h|�U�D���G3hj-Ïm�>>�:�ۮ��]u���Ǐ_^��%,*����T%B�NTw���!ΑU�6I���q�u��]u��X뮺���Ǐ������2�)��#}�<B��(*�q:J�����n�5�u�]u��X뮺���Ǐ_^��ڹs1��N%�e���$!
#��fS��m��Ƿ]uק]u�]u���Ǐ__<�HT��PQy(�q/D���u։>�>�ȸދm�����Yr�5��2"Ι�,��%�L��\����DD"R_�T+�2�EP�����ˢ��	>�۟��~G��J}�p*�%ba��DN��B&�"��!Ȼ�"�.QTH<<$�(Qd��'�sw.�q쾗��Z�᧒b��\la���CC�i�Z���D�k�;}�:��7�c������?H	N?�����h%Ő��ڂ[m����ENW������ʠ}��t�����^=�{ϨS��[kN��û��5sq��aUl��5H�~�Cܔը��4�s_yJ���	\T6�F�Xz�
�d�Nq�W�FGV�ɨ噶w(�u�����zw��3�>g���!2��ڙ��^��]�}��*���F��)���$��V�_S�w�����W�=}�h|��>`�������Zo�K�5���p�7�����N�i���	'��n����_>�t	/�� �k����4����ٕ	�DsbX��hWɣ�7v�;�.xL3w<�ݚ�Q��u��2̋׭@���`S:y��j�:�d���m�S�ΝlvpǇ�79Yu�WQ8�/�ڞ�w�r�{�A ���Y��--N;2�J�S�w��6�
3�	�|�DG�{��Wj�Z��}��X�0>�r��_���� �=������	 ~��GX���i��N�S=�H��Or���SGt
n��&���Oٹ�۶�����g�m��E0ۘ�s[��h���c߰tkL8���mɸ=%T\\'c{�`����[���6~��W����A[�s~bAc�s������zn��&gK�'ݰW�UB��ٝ��(�eM�o���\*7���),v˰l핱_a������D��Z��Pα��/-���M����`��H�m�%��j*  ��f���o���E�2�ç���>[>�|�.�;Yj�3)YM[O8��� b��;r��x)�4��Fh�i݉.�B�8�S��-�.�5�)�V�)��gY_Y:��3kuC���A�����⪏y8�oP������y�xc�Q�n���70�1e�U���ۖ�]}��znj�;^A1�\��1���p��~hO�9�]`c�[M�#M(Q����������t���u�yI�T��q�"0�,��rqYQ��ju�Bu��d�ݳR|n��C8�C���$�������!��*��(���?��~<8t&v�]D�0v�Gfmt�}�s��~�Yޫ�g+��i�Ĺ������o�U�u�u��ޞ���A���k�=�}Г�����U3~f}�a��3�`ON;���ow�#9ێ����!ٖ<���5
FH׌�E@^i�2����\
[(X#T���9:��h��Q��TG喂�W|��PO������o�ibT��4��I"s��~<i���V��]��*L�����R�f֖I!��>},5����ԩ�}]0l��웻��`٭�p(�9of�фɲ��f�(Q��i1nݣ�^��ڌ��[�� �W��x�m��7X�m����j���y:}���?���	3h��͙��i��c�ϖgpK:��^M�:�)��z��0޳�b��Ru��j�
o�a#��m~D<d���\u�z�>�f�9!��{��J[�@XʱЩ��{TI$�o�h��zHa�p��ؖL|$��ƾ>�Z�����]��y�Wox�`xO��N���T3����5LLΨR���C��{������񾦞C�#,��A9���'��ql��X�ug��-�2F�=�,���X�����<mT�����n�H?�}�{��m��`��OУ�^�j� >q�@�ܒ�Y�OE)�k31��q�׻u���y�_�k�o���7�!"-*�ެ�ǥƴc�a��u�},���B�n�R���߫����1Y�eyQ��A�? �]^�|���vƉN����Q�z���+Oӣ�ޘț�RkN�֬;%��E��� �z���o������,5����W��%�>W7He���5�N���h�����%ldWwJ`X���?��ضã�=��L�C���s.[�c�`����w���N��9����S�ձ,	0�[���=�\�,�uw;�3��L��M�;��\7iˤv�2ve���9���<S�lۥ�I����\�]�wm�Unق=�!^������FV_��O
����.;if�ꮂ�[��.���ں�ǻE��t�y�������^�l��m@-��m��l���,�����?u�s|�>��������^�ߌ�׆D�B�T�G7K�tP�}В\kNA�]w����*LÝy��`��W���ʀ���L	m��-[���pV<�c�G��td=����0�d��k}�R3�M19������<y��:�G��L��A^��Ft�nO�pk�<w��CtWYΫ���ʜ�����b � ��_)y���9�b�'B��;m�vm���ө0���u)�j��u|~{��q
�)�����K�,{����M�A�H�e�M�jZx2~rD�M;��ɒv`��$�k�9��.�:��ѐX�	�ˌ�ĥj�QƓ�?<H�Y�|O�.ܾW�+Ѿn��b}>{��['��ˬR3�)��\��v��_90�<?y:\�y` s�q"��0�o\��Y�c2�I:���7Ni3�xt���p�K����W��폶�Y|��c�`������<�ؾz���G3�o����6���9/���#�|�а�P�4��<��g�]������p���g�J^���d8���D�f��厱��=���J|k�ѯo�Vj,Ÿ�u������5���z�Ū�훓������F�""��`�]�8z��K3mt\�y0�����=����Έ> W��Ǩ 7�m��m�6�m�\}� ��4���b��GеP���#����Uꋗ�o��0Ba��R.�1��-�7F�͘��q�sU�����|d^�bs�)bѼ�I�aGb�:��z����p�m��]��
p�r��@n�j�7GG6�>��ˀe"����?��uV�J�23U����{�M]�u�ČV�S[����p�Q��`���D�7X�4�ڞF�^�y��-��n}7���)�7�ג��F���=+������pM�s�H2��i�ys9�<�0ݪSM�4%1]٧�&�o��
xw~Ա_2��#��X'�t��}�oS��OQ`O=���ܳ�d�#'q�g�;$���,r�V A�Wդ��ZD8Q�hH1����e1�5s+ݣ��:3���ݲ�w�S���'���,%�j���j�=|%|:��/�<��B��Q��}-�B�U�����);�	�gt�I��=��'i*�+��M^Oc��^P�NZQߦ�r����";Xs�_=Йȏ~P�s_���s��Le�o����8���GE�RJ)�w�\,�}�^����P7���`���W��L�Ƭ�W�}k��/jͣ\���iKD�����E�<uL{ޫ
9���k���o�c�UZ_@�r��:�Y�1GV�g\��+)��10�;��Էྋ>����SoO��m�B�m��m�਒($��>߳�~�߻�����A��/�ȷ�.a_2)�'�ciw�|u3]���و��V�4hv����_dgk+ �o�`��Q�j˩����/!1��sTt����zҴ�w]�ݞ�|=�u򥽵��㽏�P�0=!�N�%<0s��So��&�7f!<Fe�e������5'̭)Z��j�8�nb�����Yo�1�oH>p��~��Ʊ�Dԫ�+;��]���p�3�!1�dЮW>�(}��-�)3������y��9Y+�0�v�m�uS1���.�pgkj����.�Û���]��cֽ����s+�2箚1�r��4����0am�ކ��`s@��b��J9>�xm�H�����5���p�}�[�Zl��pڽs0�	�:;�gbO�^�I�y�,("J.�lb*. -�=z�Ei�֮����|h$S�J���)hc#c���'hB���
����!��wJ�Zs�~��~��o�2��^�j�Z�}�>�4��h]7Ɵ��~ٲ��$�7Y���4s��y��fY�I�nbMG3���ƛ���L�D�|M�ŰԬ���ʅ�+����T�۪�oC�ݽKU Q-�tU��8:éx�1��yC���;�wr�-s�=̚��"v�<�y�[2~ 6��ؖE#m�"[m�"�m���W>�����:���J�Q�w^TŢQ����7��m��J�跋���nuvh;��]XV�c!�Ϲ0��rR*�i�/���~��ޠK�8�MN��`<��K�]P6�_9�uc�Nr#�{��c�"[�F�7���=�~J2�+��~j
jE��4ɥ��!NOf��U�x|9�]�G����y�(���2F�g:�aU�/B��35�9"�-��ݱ1s�hۍ�'\3p�c��(�sUD|�r�&�:�n�S���1�]'6c�T��Hnw/
�V�GSe/��}Y��/���D�� ��� s��_"��PY�r�G/���ͥۙ<�2��N�<��3�'놠�<w��(p��c�oLy�����x�0�by����;��ݙ;��'z�~ȏ17�K��FTM�����	��wi��ݲ�Ly�(��������^��b�&���,>lb{j /���v[zy�.�e���%�h�%A�5'�߃�o�R�N�#~�ֽ���t V�Ũ�'@�8��w����g:(cK���$³�^�vgX�:F`o<0�p��8�.1�c���N�jO`.SM��o�������~w�)<y;�ۅiRTa�����L��n�-�����͚9[��q�I=+*ƺe&#\P�ӱl���u!>�Yו��z�e�d�p�;ŭ�s:�9z${YÜ�i�.�ls��=�<��ﭣ��~"8��67H�m���m���m��g�yכ������7�~@}j=��ȥ��y�xT���Lsx@���}S鶞tļQ���Nҹn�k_A��zE7.���[����=5�$|����GA����kK�ESv	O���fm�"���Js���&H��ꆯ6�/��}�<���x���W��Q�'���	�[=o̓�	E� ��O#h#4�I��}��]i��s�v]Fj�GCq1���L�ar'�����oF�ϗ�{��h>}$��}zO.�k��C�ś$�3��*��Q:j����x���{ y4�.���qB���s����`Ys��Y�����Ӝ��Z�I��_�erZXH��\E�iz�d��[2Ԋ�p#Xf��rv����K��01>+7^>s�����&7�.�;D��z>�:��'�+�-�M�P��eY&=�\ox��S6�� {o駣��>Tx�"O���Q��G���_��H�L%	<�-ü�P?�{���܉�t��G`\�P�x�J88�j'u&�����nH���DeeU,2,�71@���F3�E���40�lwd
�OM���7�t�;���@����ҝzۤ=[C�=�a_"jVκ��� ���g�#�#Y(�a{�.%��<�8��(�'�,�kw��룣��!�#�����`���j6�m���Qd$ ��w������:�(���<��<����O�pw'��q��;2����c�֞��9��՞�|	�����Q7�dPX�ۮE����E4���a�z�oRF�l4��v��#rU��e����^��5�\�!��z`���Y�������at�%��Է��k���6x&��c=+��q�S^�1�|<�Շ>S8�s[���-a����u�TcD��7��ዂ�������W��W\���֫'�E��l��{�@�~�&�Θ���:!�ɓ���1n�"�^9�{��=�-�-���Glo��hO�km���n�n<{!����)�y�5��GL1A�n@ߤW?u�Z�=z-�2�5�U�r�7��Z�,S�M�7w�d ��\ђ�s��1M��A�V�@ �G6x-�2�̦s��=��=w�H�8�����O�w��>Y��8QӛW<D����9s��.4���tt�e�����y.��i;�b��� �|��uTS��H3q��~�(�����*�Zۗ�������k��#;Dm�Y�nR�1 {]�j&5���m� B �C_���p�.����`���y:����jT�g$2���8o���]��f�wx���^n�5�b�?ダ>W?q� ���Q-��E-��UF�����rg�t�&�-�n�t����ZJ�V A^�a��@�����n���\��f�e�W
�e��S:�gw�%?z�{kPX#Q�Z�������G���a5)v�Y�K����L	.��/ж߽��"�g�5��X�O��b	P-+`&���a�x�fD�5�S]_Z�t󻙦����l�[���;��vk�R�n�K�f�-�J"!y��8���k�2����
��>P����Y��t�����,Y�/=@���a�Ծ��U,���yD����}>����W�^X�Mc�$�y�A_�*^��Z�\�e��S,Z5�����c�[�#lȉpΙ�U��S�ݷ�^45�)���,���>�
�}x*�nW[܂�H�?~��R�ʅ�o����t�}��j����R�k�?��	��f!���YT�̄��-j��1���Y�|���i�ǫ@U�`�e��H�s���ﷹ[�4J�,!�B�fi+�>A�S���k	Z����e0���`F�c������/{~�0��1<�AUםK�3j����k	��;�C�GNӻgF��EX6�K]2�F���7&,Z;{�#k4�.R!Ǳ {%��]V5�<H>����=f���������9z��٫���8�)S�;^��GJ7]�F�ޖ�;�K�D\�ƣ��X�օ�ppa��Tt�`�ie�W�A��l-~�z�b�sv��0*�21�����Q�&��[6�R���H7o����dD��/��jne>e3MKQM͎�o@=�Cz�uɝy'p���:�K9��ż��t7D�k�V��O<���q�}1_9�vq��R\�M�:;Ĺj{_L�Y[7�뙆��w=�.�n=���q�sb����G���.�+owMvgk)�w�4EL��bVN��3i�Ә-�N�������ɽ�ݽ,Z���G���A�X�[����"�ѲWg(j�3���]2�3��lm�i�WϹ��j�3����:��,�L7{ D�<��D,뀒���w��J_T�7	{"��i%	���E�V�;_]d�NU%v;K�dpYVd��e���Z:j��m�yn�ts5O`�o��y,"�9Ic���y{rndj��i�D�iv�*ҶSq�l1h�(�_
"�)q�/$���|�~���A!ܾ۶�F��"��潦M/��J�e��Mr�A�|����VK"8Za����Q�Ob�d�)Q3%�/6�z5ۢ�N���r���}��-k%\��B��.̎�_>�ɹK��˯m��&�X�f�����^�N���v����wR�nV�34�2u��v��B7͜z�Q��)�_�;yT�R���Ɣ���/g�8uS�����-��SF>A��^q���6_*{��Y�7�\���C9.���ّ@g,6���c�����J���ݽ�`��UV�*���Z�s�fʫS:Ηj#�x�\��bw
������X�ӵX�,��^^��a#0�����b�^_�s����ȸj���V(\8�/�[�2��9������E�D����4���%�Y-��r��X�=M.|��A�4s�5�2*��R���:��Fg"DU!�G ��8Y"�9c{���;V,4;�B��-e]I���Z���w��un��^8QUp�й�wz��ծ���54���n��V�T����ұ����&vV��az�m�b����m뭒��de�u]|,qK{J{�'J�.	�� A�o:PU��f��5/�k��������NG
���	>W�QH�H�D~$+��8Z�,ҫS{��j!$TG)q�n8�����]zu�Zu�^<<~o�����p��E߆g
���,�Ȱ�*���(�~�v}m��m�]u�^�u֝u׏^<x���亨�� `������kkߟ��A�gNbp�����8�ۮ���]i�]x���Ǐ����~$��EK+H�2T�ٕ��\�U��(�R+�-��q�u�]x뮴뮼x��|�7��ߟn�\�t��EhEY�!J�̹���I�����5�����(�IY��RD���+ �������U����ӨGJ��!�o�,z��DmYZ�*�sC$�U)�W��R�T(�U����:RHD(�QED�$���;� M<��}��(*<�*w)ep��ԏ�[�(T�N��eY�D��PI�ֳ���>��w>[@D�2 ��I�K	 ����8B� �āHRB$�@�p�|�q�8��zo,��GrGyjH�<L��hKq�8cP�0���|>u�;y.�#`4{ؑ�c�T3�����8�D ��t��F�M�bR��U�*woOFj"Ze�K	���|D���@�@Fc$��$dB�3�&gl��)W��S�އ��y.���,q#��:��_>���j�=������U���{�/x�Qu^��Tx�O*ur�1 �%7#�@KE��i��2��D)I
%��#	��ʄ0�nY�H�L4D�9FQ��9�r��� [m�+m�؍��h�U�|��Wi�ב[/�󵵽��k��Rv+t)�}!�.,������;i�i�Q��Q�'�d_��i>@������LE�^f�����k�r�S�؟a��<�|�Y�F�gKu�)��9���5���|�s���F>�����/R)�5O	q�7Fr��eʖ��1�����$SJ����Zć�,{`������e���c�N�)Z�����8	��2\g��P��54����G��cg��k,��d��++5c;7s�cXcH�R)�.VF�M�������4��Ѭ6;�V*���/v���^���%s"YLl��4����~�oUB���F��`cgv���F.[���8~�0�/|�h�<�(��YV��O�d��i�t޿}>��\�%�R��݀{����?#>4xKHa����8y���[���d�	�{���	��\[��˜ͮ��G{v��g���-���3O�����Ͼ=�Fx�4������?|���|��~��Hl\�MM�����d���3����Cϝ~�X�@�-��>x<��J?bJ�G�=�f):~i[�Y2�[�G�o`�a�6WU�9<RK��*�G��e����9��{D�l�����"��H��Wj�G�;�p\�(�kU;���V����*��R��e=���H�d3�N����$�{9��|ݫ;�gD�Q;i�mR�m�m�İ���m����"��wޞ�����`ݖ����HQ��f{�AR��̵Rʼ��� "8�t�wYf���4�E�k{N�=�~M<�D��g�1bG(={6q=c� �諝W��[R�}�w�E^�#m���^#�G��v� �����+���RݪZ�f%=�Y��|�iݧ��ثgv�e�2���D�|��,8E�=�Ǳ�O\c@�!��,��LHf,�u���R�����ƅPKҵ��[=�S��ȉ:�s�*�~!��:%;*�Ӷ�~���%����GO[vׂ�˻���sp3}�̊V�>0��+�yÑh5t�}�|=ʲ/5����g����Y0�z{��� ��w�/����j���x^�a<:=B����[����i�����r�=%�V7L1go�^aT�W����X㙒�qS}G:Χa����A�r�^�ĶځQ���n�#��$��k8�՚%�W=��o�������F�K֎~^;� d��A��hj���B�_���Rq
�����n��:_b��:똮��0:�e�tq=Z�Qո�i<m��qjQ"��d\�u86i��hg�f��x���W��[ܯ�i�+�q��̔0wM��C��=��vgT�o�	Z=r�Z�j�QY�3�V��������h6�m��m��\@<�<=����[��q�Y߃y���u�v�� ���O�sB�O��Yr�
�}��
mI1hOvMMdl"t�eo�+�����/Ö���(k��o���xǈ���%z�u�����oPŦA�s�7���( -���Z�rɕ=�zh����p/@�Bh=9���o[.a�e�2Cc��R$nė%ٓhJ���w�^J�i\�}��?��ռ��긴2�e��}��`q?�͛9�������EϾu�x|�$Ky,s=��w������3-A�{�^'���Aq�-�=ŲU�TG�j/���t�����P��d�iv����ö�u��7��^j��/��X>��Oy�}���c�Z�kw0h����׵% �\c�U����B\t���	^b�'������|<q��}#��_��ix�lߑ�}�$�ehȔ}*�
j���z���xx�L<��;��ޡТFgw8Z������[���i��p�
�H���%ؽ�r�����qo�l6ޚ8���d���uEߡ�;]�*�]���Ѻ���?t,��?�V�i��e�8�\�*�;ǈ�_�k�>}�מ���<����s��
ݕ�`n�=��&^-��u�:m;�O��Z`�t���i�t�7��mU�7;�ݺ7zL��C��|�����l�m�m���'��[�D#�s|^�ą,#|��S�Pj��O���i�����~��a6S<ז��^V��ڻ���2��[���d��1��Ƃ�\}+f�.=�����3GfM�uŔ5B���>�K�r"o��@�&�ŴHC��9�H�K���=�$й�"���Z�	ǣ��Ԟ�ݾ�<��e�ou;	��#r]z�5��SmxĴ��P0v�눇��c[��J�q<36��Z2[��]k	S�����A��>�"�狯��,�p�ɣ�vJ9��N�����;�JFO=��I�_�O����C��V�g�
/�=���R%أ2wڵw|�J%w�i�q"O�u:F���[bS�]�k���\sp�SQ�11�V����ܭ�|	��a1aq��~��#��ʱ�������n����$��^K�u�� P�z��������$3�f����Y����2�
ypn�f����W���=߶�à�|�}���bt�Ռ�ѬH<��И��B*�F��,��^�ʚMzϱ��4���w���q�X���vkrz���˒˚�V��V�v`���_*�
�7.1}[b%�<	�cƫ���[�;C�Zu�Y�c���/&�	4h�j���x�ޚ7`�ڞV�y�l���O�|~n�,�m�Ķ��x�G� �Ġ(V
בu��7��1�S���v������8QJQ�������/�ʟlۥ��ඇ�U��;3����P���FȨ�v�wc�|o�`�t����m�cG�zk�	�����!�"i�k�E�P�;۰�Ci�"�2��-�]�ڑ�L�p��l2�tv�S�c�Rn7���Y~Rǥ���i$g&�q�"�������&}�#��2%<#r�ۡoV���̸�=Xv�;����
9�l0j>s:Tz��h(F��ħK�0�^��|=�!�2����G�\�ktA*[���ӥ�Q*"�_|���]5x�~��>���Z5QL��qj���eV�'����I��C����,1�rk�Cmt����h�esR%U�\r:y��&�1��"[�ex�78]�����<zh�����<2D@M�Z��5kD
֎���������J2��z��'�tܜ�[
[���oX]��X!j<)e��n?_{zn�,����ޘ0�3�="�D35{�c�-����P���u�gʒ��a ���F1g���|��y���������:�X`��n�����BdL���r{���{����S#-3y�]w�(�U
�s�T�����Z5c���D�vd�;{y��5.f,+n�I����y�k]'���ްO���	 ��� �K��)����k���ݢkuk:\�]�ڬ�Ou���k�W��j��xJ<
���Z�S;H�}�2��!����-���m�-��D^y��4�7��|`0g`pn�v���R�ۏ"�S*���N��Ȩ�cĝ�z���]Crp�Ň8�xQ��u����
��{�`�ͩᛟw�y�-��'#�gBfl�U��Iz�32��w�$�}��8}І��#e%���B?�]Yς_[8��Т�ߵ�D�[��wgHE�=�I����o��z��yC-�>�@��[��3n0r���F��t��kV�_����{�T���L'�ީmO����m�n��KQ]��d�r_*�M��1�`|��cОEO��{�o�[@P=BVv!_�#W)�������z}�։�6��=��Z�)� ����1����p����|srt7���"�(�g�u}��a���/}���}�x�V|<�m���>�=k
���avƘێ��"�Y[�F���A'�����!_�EiPc��h ��ݘ�\!�,��2�G�Okb*�cu�2�����u�]"�(wus[9��c�p�@Ǔ1-T��0G���=�^��]����[w%Љ��������k9��FR�]�v��J�od�$��ך!8/"y3l�������p�"���-�Ia!���rNlw��z09������}WSjk�33B�����s����� ||�� ��mm��C�����}���7��Qe�GGO�k�LPP'��/�Y�Q���w�}k�zCP�Qj���"ךC����^E#�f�-��z��_�[5@�����Rkz��]8����:������!���+Mp���M?c������yz�t�:����ʲ�Ƹ���p��{mh���Z�t�Tȝ~����2KV�r�Y{�iR{��D��Zj���\���]U�	[�uϣ��e� �_O@"|A[�G؈/Z��rZ�P��02�(q����i�ac��1��W���C�mimv�;�դ�b4��-���]�f�N�n�f�c��gX{��x-����il�a�v$���-��@�1(����[���Yp���V��[A%�������1���ޜ���N�Iz&L�۸s�kK9��C��jy8�t��Y�0�\n�y�g����Ã�h�4�)�C�_:������Q���@!��34�i��#G�敛K�i��<��곪�8bIGfٖ�ԐJ|_�t��Z}�؜��9N�_|��}Z>�}�
�^Zz4��蚽X�q�M\��B��9W]jD:+T�%����Ԛ�P'&�B��{1o�����$�ex��5@5
�+�dr��,Y�{�F��Ɂ�N��Uoo7������D��tͩd�m����Ϲ��>>>>�m���b�}�w���o[n}�?7ް2�,�v��m��L}�����"�{aB.��g�܁�� ؤ���z��c�MhqJm�Tn$E���ֿ�7!T�i�U�~��	R�^{�C�2!0㝝�=�{]�8���J��[Ç9���_Rw�q�sC��]��U}1�c���6<�s�����34
t�>��À�έr�Tt�Tx�������;7,�ukpѮ=�=��'�6K�hj�t��rA�zm��;�Pl�\f?Z�}=�]wok숞�d{��xy����h/�-^u�M��X7]j����,�SW�t�i��2f^b'�6���@��ϧT	��w���!���7K��/)n9��22���i�n�S�Z{��P��t&\za���6@��|y�a���tm��zO��WZ�#�ۍѳ��-��c��R]I���+�u�-\dy��F���&�4>���R<��=�;&wI���1�s��B���N�s�:OL�uI`�F�jbA�÷n�+zfx�݅2	��B.�-�P�ʱP��33sY�V�S��r�U�n���	���̫M�3�sH1`���؅+��ۘ�z����fh�u��쬘^�!��ٕa�{�q��f�T��dj���Ko�lo�vH���'�����W��m�-��R�m���ξ���¬#�Vs�w�¨aȎ���rWX�K�9�U��%&�xlO-��C9�}�@c7�ۍ��n���hR��=�ٙ7��y�5gt�A9�/`����\&x�C�uq˚͝�+G �2�E���膛췑�+����p�ҘO��/D�y�k�Vo?U\����ͽ��������j�Q�>�#�O��Q�j�NϾ��2)8��S�(j�I����r�����l�N�;\�	C�ǆ���!?y3-Bh������=�{�ز����HG�9�ԘB疯]�4�oT�+Q�`����_�#��YUa��1�^��=�he�߱�z�|�xD�w�, �b��}M�3�ӹ� �j��-ԥ�m8�қ��+��oM��f)�S�t8���lUn��i&��L����y�y�ф�7=uH�l4ɣ��a^������u�G�z��0߸Nwӟ�a�&s�=;�֮�Ù��d�Dz��V[ܼ�b"��~���}�e~P�VB��{���Lj��.������U��n]�6�,��og�ۗt�׭r�w���)��:����G� ��	\`.��=װ]�v(���ʐUL�Q	����.�u.q�ّl��;ޔ�ud�n��R���onl�g���	�~����#];٨�N��	����Y�:����U�[en�0��1��0���)���sXA�0�� ���@����b[m���b�y�y���y�{���f�/8�W<��ybG�UJ:f`�����ǡȁ�i�/5�U��i���H�^�`��������b���wB�=��5���!�P]�_>��� i��勶�$Y�wvv���v��<3�T&9�i>-�Bɏs\�Xލn��K׺��P	�����wB:r�͂e/,/��0����_P�g)���>]xE����W��I��4�0�9�b�q�s�MOL3ìW�XC�o����D��u���c�A�k�s��gf�ڪ�s{� /]/s:�g�pA��`�:�+�XL��mt�,���V�0�8:v�����}4��3F8�n<x��;5*��@Ӱ$l���i`^� s��RǷ�ߓ%b����mJ.���3 �$8�*Y��	�>ʩKg��_��z���M��F{D$�
"�[�>7sԽXF�H�O�uܞ#���>�"Z�/��� ���;յ�e���S;�	榑�@����~���zh���P}�F��	�7!��Qz��/l���?V�p�xi8D�Ꜥέ����;H�$!b�W��v��Ͳ�v8#:N���Q8&��3}�u�*�;zm�QWYl�%��N�@����vś�Lu�)q��1��1��epy� �#���b%w����e���Z���in*g@]�0t��E����n�9�ki��+,>u��s�SE�C�ђ��g�ɠ�Tn�e�]�|o����0ņ6�A�FV���
�v�cN�˱�8Ei�^��q�^�,_A�,�ة��e����l�/����MbJؒ�d.��s�,aY.f)>��ғ��>�x��޳F�����H��ti�ܟEU�αb7ܓ�ڝR��&K���z�Wq�WT�z����0�A8L�@ku+���� ɫ��Y�%k�\ҦmC���ݖ�ؼԴo\4e�G�@[���D�Gb���+x*L�@�ۜM�au���"VhK�[&~/R��*EөT����D�xn��]�r�L����ͤ��13��u:`)�DU�T\�t.��5�٫
����F^U�Y��/ ���xs��:�P�g7F��E�w�)�]�д5y���R����Ϡf֥��!,�k �"]p[�B��e�՛ٹ��7n�)�VG�!.UZ�OlqU����%�������'ȋ�L�Z���
���&5J��,�7D�����# ݺ���!MZ��Un_�>�Wm��k$=nA��vU����Ԯ�X�����3����S����'����o�c����B��>���8�O�/oqAT�I�G�>�o�z�~����/���;�w��^�k��_U̅\t�L�-p�+z��j٦e���:�Sd��:���)+��H?Z�{h:��&��/tB�n�Y=;�L�cxǹ�9�:f�kB�� !u�5�ѳM1v������˧mՍG��3�l��__����O�O��
Qგ[sjj���\���_X�S=e���on\ќ/�R��'�q�9��o8�Z$��e���Ŷ�il�oF-屛Q�L�F�	������gd���h(����0]"w(��%�̹7e2l���fc�7��E�{}x�wוދ:����b�nƬ�k����y�j-��N��!��ufVIJ^�ٝ�*t�Lw]k-�!;7{sNQn��J�#rZ����'���*�P��C^특��q���N��5>x��e���h���d�������DRx:�^A~��h;��.�p������;q혩(�*���޻bV�N�E�]ꑚ�:��v�oD&����.�*�6���"��W{f#y#`��q�ZNVU7���]ה��#�F��?_���7V����O�u�P�e�Aë3>��D~���!2�֕��^�@/_}vZL�{�|���7�����^:�:�8������g�AU�j"[5*De�z�TG3*3��3�@�W���}q�]u׎�뭺�Ǐ^<�����T�VjU)Y�Ћ���eu�ޜ������u�]u㮺�n����׏_w��U��ih�QQ\�0��H��U5H#D+R�o�6��u�]x뮺ۮ�x��������~S�r�ATUA�dr ��C	��ͳ��1��"!I!ov�W|�r �E�&Tb%[B=s�!��O*��^�����-
�#~'r�G
��Be�YT�dQW
���N詭9R�/:x~���Y�P�P��R�]D �U%%���hYVF�Z�2T�˲(�)�i*k*6(HF���N�NhF��gH.�}�$�,Y`PT&f*QQ5L�!UME-A6~����w�~~~}�{*F���ΗoarGL�,6����ڰ�q�Ks �����{9�y����:��l���v�m�m�m��5}}�����N��,�)�P�՜+��v
I�B˺$?|����O�^A�XA�w![��Cݞl{n����Z�9�Wϛ/���x�*�O���"�c�Pc���W�P��޸���3����P!�۲Y'���n�X��C��������4�q!������X�u��i[iNs#��К��Ӓ�bK�]"�y�������A87��5���0�n�(؋��������M�����^��q�Ϊ��Q�ӨX�c����Xk 1:��y㞨䜤uz"�4⽵��;�.=Ё��r|��-5�$���^[��=���7cz�a����V��ZÀ���/�<�q�'O���'! v��D�Gc�$st���������e�=��C�%+(�=��gH!t�|o��οC�m���'�����S74�J�t`��ݙjpk!��7��UC5z.��z}a>��vO��cѭ���
%�k��Si�w��C�o[�˳��^��wL�&4��^6}���C�3��ţ��!���ӄc4*_���uJzJ5��w�X3�"�K���T����i*�u�gn�/��=_·��	��yn�Ĳ� �G�"jDx��S�o5�W8�ۗ��Q\����Ĵ#��	r���q����s��w>|�͝�s���[��]Km���m��m������y���ѯ���& �j�i|��'٦Y�f�E�'�'���v��g8���sUf���L�E8gsNz`sY!���H�ؒ�L3&I������;z��B�1�|���7��.�a�7~k�~Uƨߗ׏�y5C���d���8/�82�in�sV�-t��y�f�ߛ-�j�V<�wМA����'��d����9ָ|�Ǘ�꾅�����`K���sxy�g�]ㆾP|�X1���u��+"���k��O�!�xf�
d����c�SV/A����P~�����.:g���X|I�y���C=TVE��tFQ��&CfּD�KL�	��|d�n��CSN�zK�T+!Ja,�ݝ�|���լ9�in�v1�*����}��|W
��=\��O%9hhtŗk��z}�N�r�<�:{�]��0g�jM]ԟ[�qi��%��zڧ�q�C�G��8���$��Ӡ���g�`���Xc"��bL"��DB�᧍��΢�۹\x�#;�xO o����O�(�i0y��<�i��X͐��f�~�z6v ��]�Y��Cn%��d�]�!�N3�b�%rW�<���X;�J�2�Vι���v�Y�fv��GIm���%}�鋘����b���scGS�Jv�A�{��z��d�o�q����x�6�m���v�m�w���>��f�W��GU��ܧ�ѭ�X"�3��'nЛr�ʍ�#a����y�gn����&S�*�~:��o~��m�l�Wā�����������=o�� y�N2��Zy0�|�-H�e??s�Hq��#O�c]�d�ͬ�6]bQ,���M�$�Y��@4�|`WՌ(Q  5��2;�XJ{l<� W����$��9�5�O=5[����h��qp�(K�e^�
�<�q>'g���'��~�gcCs�0k�Yc���N�o���%|��Yϕ���|h�uS�<`�5�}<��Q>f�	Uy��6���Y��k4�^��&Mw��0���B@���\�����m�W��A޸@��#b�3�ӓk��5��߹���zn{D�3Tb�,^�Ƨ��:�H�TF���d�L����qx������=���7k���ߙ/z.)�)3�%��֠�^�޺缊�w}��[i)�bL�j�b��L�����υ,��v;jb����+��vY����/�#�� ���+��*
 �|��1���7u���T���-Yp�z%���5��5�\���F�:ζ��Nt �֗r��b]�Ki$Ood;}�$�/;,���`����ڱ�ג���v	�/nK�a�&�+zQ`���>Y7�h5j�'9�[�#E�&�����{+�|��s!���M4�m�ݶ�k^������o޴��4��ǥ��T}�.q�!t�a��������kQ�%�$���kᾯ�s�O��V϶�`����5i����j�c�Cq���焓B����N���*wOS��Ɩ^�y:1g�7[W�������)^=VW'��	/
@���{5�C�9}cDu8��--��D�d��}�OY}�ps4�=��fjۺ�y��_;"}w�u������n����uV�j�.Ng�
8O:�#��9����,t�����4��ȴ��W�p!\"|��r �4�\�qx�>��Z�t�
[Bq-���l{c��۳�~��w�߳U)��3��|�����t��w���cq��P���K��P��>��eٹ����[0�7�q� >�#����G\��X!���v}�ͻ�1������9��q[w��������H���>��3���F���hc�[\�t}A��P��_})gwF���y5����kH9r��A�ְN�y���T">Y��{�O��4I_�N)aN�Ո7,��n��6�%�2���"Zjҫ�p��d;؇[y����{���7�v�=�����U؍��h铈��Vƺo6I���s�̮\�O÷��4�v�m4�`w�<�Ow�ם�T៼߁A�����i: vQ5��������8�ܷb��f���_���~^� Y�<y�������Ǒ80��I��_S=� �u_��}�<!�跥����-���EM�������3M�������6�]�;��;^�.>�
�����,+w�y��,{�,²m/,v�5��i	�l�v��F��vn�)g���v�
4W�}$Ņ��K=7�|`�}s~l�O��_5�F�h�xzV���B��w�$����e�)I��������P�Gڬz��F��8e����]ecw��0��\�ȉJ��結^�Z=��z^��pP#���G��$/fD�|�k_;?���"�zm��X�b🷺}��<���$nE���|oʘ[��nd�}����$�H%ĉ������Y�!��|C<g�m�nD2+�t���b˘��4q���FNj���`|C�"��1���sX*�y���w]�na�3�x�{;S��v�G�9��C+64<���">�:��b�;mJ��n�@��;Qe�#S%� Ѣ9^G�u�;a� O�>U��3O��e�m�Vѕ��;���	��E��P�v䆉�e�Wk��0'o3��ם�'}������M7m�ݶ�`}�,ҙq����|����	.`4S��<7��{����K�U�	?f��x�!��ve����������y�cYt����9���E�˃�H~�U�tЙ���6������<^=���m��k�
I�s-�g?>�~>�m{B�~�� Ļ���]OZ����e�'e"�FT�t��I95
v�N�{g|��kjؽsj��$�0�A�z�� vW?��Kk[ 敲�������FAp{.ov�{/ǂ�z�r+��W�����u�r�3���<�L[yu��c�i�C����6�G�`�����5ʀ�6���8��k7u��2��80��u��zA���'{��ʺ��/L�Yd[u�|���	�����+)N�x�g�\��}"b�ji������$�9e�kQ:�҉����Iڊ�s��P�n����PN��czöz��S��m��C�����B�n_�q`�l�UV��}_�d�Y�_u��hb��<cdt:MJ�]
��2E�em�u�:��K��>�([�U�p�K	�؝kj��u�ڍ������G����$K��d�*U�U�M��Q%ф��w>���n�w�޺r6����V��J�v�ќa�tbA,5m�٥ԫ����f�+�s������Vy^�s��9^lGmf��6�`ލ�M˓H8�z�&���z{��r���jW�E�~�S����5�'��$K+U��U� ��Ci�+��;A�ڇ����{�}�&����H���j^��}>�â<���G :䷋�l�d�l�n�\MYقV�ч��:c`�A���ڵ7����G�.����<��m��6�k"Y�;�]��>&;��+S��g�u�\4�����p&!�6\�������ds磋±G�F�{�U����޽�c�ʭ��s�W�|�*���䪣���"��`���I]ӝ���.µG빼T�0������(���p��@�S�1Q��b�`�oO��s9&wI�7��+{W�r��CͣMy��`.�Q��"��"?ď쏲��c�dK��gؖ|l}S!�wN�������)Y�6�윺F�К��R�\&�hȝ��z���n(Fv��r��VNZ*lFor���8Ɂ$Ss�XR�.�'�)��*�]�eJ�5Ң2.�&��~�=���{3������G�ʣ���/�+���>�6��'����GD<u*���8������b�'x���猼9��*O����<0��Tz�} ώ��R�.%��G�U�q�W���Nt�S�<LD�����ּ���$�j�/�YJv)�!��#a�C6)�̾X!\�eC���q��6M��הw&���X���l+:�0�g��P�qU�X��"����oi���)�DL�����Z�f��F.EM=u��<�n].�t��#|���;�{���ըZ�kxkJeD�d>�ws�ꚇ�^�y������<H��W0�u�"D=��t�5�U	�_x��E�/���zzRK�ͯK&�h� Ϝd�n��'R����_bŵl0��7�D��4bo���� ����e�f�o���s�=��U[�j�ꂑ�E�|�G��(���|��_?X�0;S�&�B��s'���ܓ�Ve���4<3<ݘ�)�L�M�6��
ѵm$��dY��_�؄I��%6�I���u�{��
T�!��\Ħ���u�����C�v����g	�YN�SO�$�>uQ��Kk�%m���}:?.{�������?����)vWX,�o�������fi��R�G��'�g�Еj����ŸބN9���(Ѯ閏E�^�iw�w�N�t�a��#�vQ'6�T��G7f7!հ������ �q�ta�v�/��g:w�;h[�����L�}�%v�J�=�,��aF��Nc�]Ni;|���ywEb��?���#l,�N��C[6�x>���y�W6дI��J��y��T�c��B���`�Kj׬���D�Y��g�l�0%Cl��)\����F}��{P�-y����æ�gb���X�O
lk~ j�����G�G��ނ=�4k�Ŷ"����H�b0��5>jͽ�c�Y��f8
#�[�0��Nk�52�3;8��-�5�g�M��\TK��ë=^�e�Äz�Z'2��N�<��o�P�K���� YNO��b]���׎�f٪�]�16��X�|eKC���}�� a�>�,���w�0A�waIY�����C5�0��/P��]EՖ���*<�ݣ9o^�/�y)m��7t�M˗��|�����m���m�d ����w�f��Z~p�7ɏZ!�#� �M3��5EO��wO5�#oJR��޺��%�9P=�'���R�h���z���GF\i=�a�x**��~�������x0�}��f��qθ�a�69��#^��ۍ�eUWUN���W6��p����D�d�x�i��$��i�M�uv�w4����܎>� \�-��l:�cdWMR}z��柌j�zsy.�ߨg&R�q��y�8=�}�.n\_Ti�K)��f"n.%�"d;D���rW3��}hz:o�dl�ߘ%�mzF׎t9�9/�۹Rv���
�ԖΟn�I$)�o�%�@T�/'���Y�[�kȉ�~]!��������184�����,��M^�5R�N�{���4k@���ko�;݃.{cr贗���j�tέ�K=��%�P��*�5��m�+J��1s�_���ν��8�O0���SqU��������խ=9(��QǗau�Ѯ�Pٺjv�i�f ��th�mZuսI"u���^-�t18��G�/�bW��c���O"��i�
�,Es	;]�^E�ǝȪKh�@gV�0DmN�v���J���W�3NKg�ɕ+t��E��8_��|�8m����h�	*9{Z\ii�v��#K1moj�9R��[ePqE�� �d�(��-u�{�n�����yܜ{q$����f��r��-Wǳt��4�ѱre��TC�ofF\�h��qt�bj�lfZ��ۥ%bJ�^��}G�Ly��n�(^�t�ٜ���oSs�6���l�&H�X9��@�T�U����*;�x��S�Zʊ�4��Ɓ��V�%���oer�G�L��9y��.���F\���\.a��z�"��f��Q3Rt����i;�E���V��R��
�v�z�f�Ǜ0��j�#؅b�����1��x6���,K�i=1�y�y]���Qû�#�o��d��K�6󨨵?uy좳���B8gQK�:<�55`�lr���[vv� ��g#h�Y��ދ�VءWU�k��G�WE�P�ZX4�]�6�����Rww[K��\h��������	��	5UW/�v��5���3��ȷ�a�̚}���`=cS�mV�I��2��R��Ԟ0�Vr�0�6�သ�����: ��ݗ��sW�x�9іj.K�s2����KH���^
}��G�jV���֠�Z�7o��B_��$5��³&��&ԕ�4��弼�	��v���Y�������� ̰1���*\,�P�Ql3&�^:�8^K�k��� 2TP��Z]v{�=�^�e�	���*wۿ,�0s=���ý��˛#�:+T���3�����{��V�T���ĺ�^���72�
�5F�ǸR��b��JCu�_Wgd�:�VP��!��,Y�']{t�9Q��{�K��M�t�v(��|t[B���[C5uq�.����K�����/1�Q,����R�����5���t8K�:��
&U�R�:6�9�N���#�����3;ɚ��BٴM��u������n�`��V]��^���m�wu��,��T�����{�]0�.Xls��w��lꛛ���=��;�qҩc+�:���1��'��Dck��=t(ӷ\�Y�rm��ﺵ�y{��V(�R}�HF�<��"��V��&��w(�d���aDEʤ�}�X�)&<m��>:�:뮶�<q�K|���}����2�	R�5QIe��_\J#������I�SR�����[�<}x�뮸뮺ۮ�x��׏����?�.�hH=QR���L��Z�� �UW��}@����m�ק���:뮶�<q����߉<�@�%J��d��+�UT�ps�VJ�ӑQQ�+��]o�����<u�]q�]u�x���׏��gs�$�;�	\�ߗz
�W"8�߷}�3�AA���F��[9�u�G�Q��(��"+���/!�?L����N�\ ʳ��˨��K.�dEqd�eUʞ1�\s'��+��EEPI������0��%Y\��E�8UHl�Q��҃YEATHt��Ϋ�l��G=�\����9DU�3�)R入�(*�D*�ߎ��]�T���D(���\=D霿��~���V|wz���	� �2XH@ g�9 -CP��a�`�)�d��P2re�h��-�D��H\G�0Js��f������5/�N�,���|�l�M�!P��p>�;����H���pH8�A���A��-+ M"�jU#�YiT�������&�\�pd*D	e�"q�Tpq#e�H-��q� Q��H$$�`�rI I�#0���d�Ym ̒6 ��`R��l� M��=t^9_r=]�t�o��U�[�oxd�����{�"�������m���l-��$	|������i!|�5��/}��-�ij􉳺"X�
�{�N�+a�äY��&о2���G��?�]_=�r*�������pV�'G{K>�V4���ɘ)�@����M;5��ӏ�[�Gcj+N�`՞B6����BR���U��;���v� V4�ʮ�j�#�C�zA���"���~8�&�D���n�OX���[�N�c3wv,�׀0�]�`���4Dn5�&���Voo(��3��O��Rp��q�l�fO��NG��vyu��dnUH݄�W.�Mo�7!�ҁ++w#Z����n�H��ߢ��$���k�4y�n�VnW��*AIKml��u#�����H�� ut�ܽ����nV��%Ą�!EJ{��~T$�6�{��|��9r���O.�q�5�ȝ����*Icb�4|�E�g��u-�(�{���B����麟,����5j���*�D��X��po�r�.uϖ%i!�j�ŧc�����!ɮQ�Fg�:g����ݯ���S�벧y�p]2�=��؉�ʕyA8:��T��Y���r����|��\��<��bS�M4��m4�}�|߯oߑ�`�?_W�!)��}�@W�Ӵ-o<���{�[�ilx�v���=�6	�Q\ü���9�/}=!�cs���]c�� ���Vd�dyM{?��97z�p�S��0�������y�����W����"�#��ɧoSc�f�u�����`�Zz����d4q��㾘ܙ����^�sՆȻ�F��8��f�f��C�&ƿ�l�ӏ��*���ļuZ�L��\F$�淳v�Z�x��}��:x���01�}"��4_��z�V&��P]ٝ񠗉>��aHx�:P�|�Z�`f1�ol�w5�'4�i�z��:�:ԛYk	���\����ޕH?��y0���i_�%q������i�"��.�9�6��M�De�c�]DBױvr'��I�sRn��4�4�*�dz�U��ߍ��h
�&�⚬̯�w�]SQ��ŧoqZ����̘6L���o�s�b�F0�$��ޱ�f�%{��|��,��Z�,i�3������]e�0���\�\�:}��3\77+���W]��8g��M4�M4�3���7Ͼ���d�1��t�-�V����>x=^�"T sfn�E�|�{�dg�i�O�q�^g��,Nw�O�V���*;RK�9�r�z�p�!�;-�����'��w?W�Fo����˧�1�=�dlϙ4�V5wܧC�oM-�mkX�m��'��C�bx�g��k���ǻS��M33�9�V�{�I��rM���?0i��f��A��k�w{bh�s��5����KsNn��6q���7k�8��|�{��&��Gs�H�1�V�Ҵ�3R��^7����]
;錠��r{%���N&��D���5�M{OJ[�9Z�#t����O�B�L4�y�8ѝҕii�7����R*��w�eL�5��k��KfJ^��� � 鲽^�§s��yq0��ѷd��Pe'�>=@@��^��"�$�A�uj����j=	&��C~����0<��
��_����� ��'�9��6�tI���+.!�Rmen��.1��Cq�>��.>��R}[��[�V��;�A�����A]��h���eA���;,F*Pjjږڂƃ~/G�<�?����?�(֙�g�7}����0;�
P�T��*�����Ϊ�0��W
6{ݑO7��tA���Tl@�q�(gg���ky��0����x��V��U�l�&�G�Y�~�	�f��&z�LBzY���0<=�%+m�p�U���V�M�i�Y�UA�ê(KF�f�BLo_W>�A@x)t«��:�8{�P\��G &V����	�o����v���3�C�t�@^�Wʯ"s����T��;�2w#�D֍��Q��2��؇xv��|B���һ��x�U��~���.O����񚦻�k�\�G3���]��s�{��F]:��Q=�s��ť�'�+�Rdݦ&�s���=�P�#$������nB�+F���+Iu�ų�m�]^�'8��g��>X^��W�L�d��Y�0���CT�4L�V��6r~�D��ڻ����ڈ�d��F+��&����򖪽���8kQ<� Y�3V9�V�����I�,ڒ�k<��\�S0L�}�,���������mH����h����?�������}�ə;<�Ϊ쭆�����U��Jo{��X�+s]�w]��cW+�� �s������r�Wb�$�:%3;�#R�%�w�J��v�饻�蠪���ٞ����*�oH�����DbaF���2 ɐ�����2�7&�	Z񓊮ڝ��j�΅�C|����\�T
�>��3�ҶR^H���PL�<��n�&Mb#�`d>���p,\��s��Xƻ��S�KU>f�w��x��S�*ppv��<f1�F����Mr��l��^�;�P��ܡZ&��۽�4�W��Agյ:�>�^��8�M&��.����]���m�[�5|�qhޯR	H�VR�V��{hx#/�p�`L�ԑZ�9���&�����]f�I4��TK�����ڨ�W9����������w���6��o�}�Mq��쒺
����=��I������
�%פ0����9�i��푻	vu�̓i�&��3U�uJ��n�Ý��F�]v7���q$w/:u֔��zg�\�5-�6��3�t`��L�o}�n��ܴ3d��:�P��3:��3�k�|tvT�-�f��X�� ����{<�?�������|։����j����>�W���fH��e�P��%�Kb�þ���+KV�m䑎�wA��Z��P��@}�!t�T�v[*)BaLY�r�597��m%�t�ų�l�1�=<�?\�[�q�8��j���n���+�/܊�#�k��Վ�/�yo�����}��t��䍿OE�yۋ�e��&��>����w)w��n������f`��C��B�]+��ߛj����i,��B8a�a�(�����Cၹ��&���y3����v}MɿG[�+�[��0��-�ڲW�|}�=�K�q��Vy����}hǞ�Y�<k�i:{�_$�%�{U��G-���̎0�{1^eړO��v�\0�O���f@�k�%�Ǵ�Ż8�\`�͕~؃�cOm$o'����Ⱥl��k��������<Qv�O�,i\v=�DR՟R�`7���)�ޱ�+@Fͻwѓ��wR���6��:V��7s��][_"wWΔO�|�];}�8���5����V�+K|�<7{b�N��^[������8y�ey�)��M4�M4�����ӎ"���e���&�z��)ra���5ed�l��x�ucV�W��Ʒ�!�`�����v�@*���(�3`�z�����i��I��!�:��ee��3�`���ub�)���흋���mVf*�U�E+Ѝ�D����:�����ΰ�!�Of��A�y�rX;�0vvv�xUƚ�G���;n�[��L�,%�)��'�V:q]��Z���OW�5��3���� �`B�)�A�6��*��]�Yt]4�}�`L4����ל�d�>��[��Kf4M��3�{�"����<��<��0�0.���<������u+v���v�aU��&D�_��\����-s�����v��@�#\u�t�3ۄɷ�'k�� Wb�u�H��v���J$і����@�s���4�vF�r&���zK�{��s�8h��'sZw��He˫�:�MK�;����A$�T(� H�|w����%�����׽����cμ�a�s�e,�p�'��;#���'y����}>2���B}ն�M4�M���kw�}�����;�T�,��=AL\�z�|��G�?��*Ѷ~If������,����i^��a>�3
�C3Z����Z�v������ԅ��G�u���[���[&J��M�!�մz��j <����մ��3�`��I��#G���p
V�=�	��8��&�0�R��h�膞��8A��+@�>��\���h����y�!;�bJ;f���z�!����B���xE����~��b�B6U<Syig��ڂ��DE׶�^v�,���P�j���z"���Oo��L%�gU0��%ڶ}=ZNO�d�*%ԍ8us<���MֈI���H�d��My����sHՒ�÷r5[�(e9�3ʬ5�<m�f{���V��Ӄ��]V�wwwM�oR�P��QT�͸�P�ssq��.�^:�����G���oçn�ˁ��W�T�-D�����v�y'
[��}+�җl�_���LN�te��� ��|ff3�Y殔���B����ՙ�gd�:�'�'����);��~�>��_���������?[�[�G�s��؇����}�L�f�m��ܕ��(�M1R`p<����5�S�������/���:��r>㚺�ީ"M�O������8�&�ָ1���0�}�5Z���f�MGw�(U�r_�a�t��h}׏f8C.��{���eBx�֧���iXqI�:{Lf�'�.8_0��F��|F�e���3��ޘ�e��H�r$�}��{����ȴ'�a3����~��g���)��k�Ź7�^G��`u�[� ��+:���=4���Ү�U윍�}K������9oV��gp@�/7:�F(қ V7w���?��j�x�f��8i2g�+��32�W?���wPuL�����lOtQ�e����q?!�˷��%ϛ|�Nz�Bu�}��H��=��[�]b���O��k.휝�b��R�]#��,m����^���u��T���Up��$Aa�3+6��tϫ+������}��W�k�U*����{3�,ᾊX�"vN�������Gk�u5ӌ$0hV�����U%��C�F�6�Wcå���F�Bޛ�$#n:�0��I��l�#r	�3�5,nIf�uc]݋��v�[�����%�㯭4�M4�O���uߞ�}��=�����Z�koJ�Y*ƫ}vO�9�{�ə����y
0�S���Q>垩L[�D��))[J��(����τ7��F�A�!�63�y�!������<��ע#,���bP����6�Әv��Ԯgx�3^Mz�1�t��q4� G���z�3�X/�����j7M!�T�IU������q��O>��@�йV�E����M���*l����Ows{*6�Z��q�+n�՛V*��{L�wC!�""|�ǧ�G;^�ӍK�V���뫊���s��6�z�ި҈��m�`	���� Q�$�u{��Z�������U|wd��>���+{��O�ߺg���;��-h�;�U�`waU���W���2��>/����r��Yۛ��G�1�S�kK�]@�̬RZ!�}����B�v�i�W�w]s�7Ǥ+f�a�'�8FeKۂ�����������ܻg��$��޾6���e��Z����x3��<&V�Dw^eYp��S�6<��\�8�u�y��l]��{��-��ːc�u(8�-�c3i�6s����W�@7*�ې��FnB����8Ej�r�d�{��E�'LѸ���K,��ٮX��-��-��Q�L��j�.�{�؃��Ͷ�#�K곰.z�pZ���7�!H��]���t����-���;�R��s�m�z�e���Xr��#�9۽s伾�%we�<wnz��q͛-3�7XE�v�`S(�Zn�[�k�_v^,6��ע�T������8j+97���+V;3D�TP�6׭X�L�׉a���m!�f%[E��ƞa����7��n��qJ眅��ŎX�M���k��UV�gEJ.Zުի̶�t���]ddIHnp7�1
dB����a�ˬ�+��$CA�}��$�0m�5�d��-ױuΧZ8(�B�ÚZ�O 9�=d�F��,��g��R�U�������V\&�
T`E��N�4�1�ͷzW��{����Jujw�|p���+wM�:U6�b��~s�ICEUc%����H4h֟6a'�M�G�9�m��B�io��L
�\%eʵ����	]\����P!P�j��b&�%a	g�^��>��)ً35ܝ�	z����j��{����-��.[�okp��C=�&�4�WKl��ViK��$����xD�6�wR����V�3���$5u��<�����u��D�}��`ـ楎�cX����L�5QS�e_+�ځU��KL��O_�VY)mN�j���:�m����]X����"�c{�e��+#Yn�1�v�
i0�{:R��1�t|����7�H��C9%��ݥ.i����L���,G_��.[�Ӯ\.���7Yڼ��Jzd��T�[����e֞ã.���F���K��;��Z8<`�n�e:��oB�{���*�V]�}����p�a�j��f�Nu��<��*�3�=:�����ኝN�O��8z"����=*�+��bT=��{[�%��Q&�����u6��\h�.�#y�2��tJ2�2/^C��N�ET{h��	�:�1Pr���B,�V��Wu*0L��M�̙���JRu���n�]V�&T��Y���/��Y
@ֿ��Z}r�����C;�n����S��*$:U��D.U͔n��_>��w>��cz�D"��v��i�@��$�x��mp��^BȹPUTW8Rd��I���n��>>�ۮ��:��ǎ>�����(�T����De�"R���NAU�r.W'h���\��o�����������뭺뮺�<x������$d"��?w���$��;S�'�EE��UEQG���6�������[u�]u�^<x��������UQ�G����q������_$�H�H�Zm��׷^�u�]u�\u�Ǐ}}}|焒�"�
�I��#V?#O*NR�D���I:�C��Z�r���_��&W�0�,ZA����Ar��ʪ"���
�D
�T��#B��sP���]]�TF��.
.��*�.US*���E\��ˆh�0�QUbE�r�E'eʫ����T%��W-\�'�\�7�B?t�kY���Mʂ'�E`��5oԅUQ�*'�W�afe�IV�j������>�����_����3�$t��Co�4V�k%t�iuۺ�N�S�tkN��ʓ!���ܡ���yyyyyyyyyxwL��}{���s��S�D��������= ��<��Q'|{���:����]�mc�O�SL��x	7�^>��"$����/g��0X�R�ԔF��Q:Jþ��˂��u>���ݨ��������K�9އ�V��-�[{:s�R!���mu_mX��}�5%��1�/����\=6�^N^��|�zSl��|y���}#�>�3��gJ0���#�R����V�5�j�E;��;���a8j�5bw����_��0�L�z�;x։�4���y}>�e���	���c��ǋs:�O�22l.Ѻq�;�Y�7�=	+@]T�CM:�C��뛗E��?]����\J|j�/���2p9	W���^Wm�h���q�t�??G^��gs"������^(H�a����Հ��$��^ʆ��r��c��b����D�<�{��t�᭮1�Y�[\�j6�t��+����Y|p���r)��:6� �� ʰ�M<w������h��� v�9S\z/��,���ܨah2nos�z�������;�7���M4���Қi��>������T;x y�W�,G��V���E@﫻�YF��H��Sfs1U%f�W��s360�d-���`���G�k��v�cg_fWo(���0����ᾇ5�;u�¤-�8��uϞ�;��Ro�ߔu�>Ӻp�JQ!-�
�}*��Y�����ӱ݌$����y�M1��҃��p��0����+���1r6�yl!�_�Y<�+��Zd����	�f=�CJ��ۀ�ߤ�3[%�6^^Wf~�{�{$�KR��w��	_���Cn����ɿV�;Gp��(�{b^y�wr7�o��/�x2c�9Ӱ�i����35ԥ�Ȑ}�u������8R�Vt(��.N�hs���4W_}��+�]ǩ������<n�0q3���*���y}���bf
��Ur�6�N_��\ڨ��f-�l�"�7�tC�Ϡ�o�����	��d���08�;�T�.׋�T�����(l)��¹8����{�L	����f�&.���;;fv��q-�Z�U�+\��8���������������g5Y�mɕ�w~�7��h���6���}��$����p���\��/�*��m:v$���WSDSë�C��3�!��P��_��l�T��Y(�dށ��6�2��L�"��O�q�Q�c�wW
��;�.���T�74苷)�_m�Wm��ա�C�{��w=\�w��_#�ް�wԡ(�n��q�}JI�2r��C[v���4��=hy�_#�cݞ�;��O�4�i �5:�y�ju��䁽^�!�.�r-y��>�q��|���=��⑳p���Rcި�R���8�u���*��ѐ9�fk�����܍���.�+U���/�oޞpF������fj<8�3}u�u����>������Ĝ��?�*��d�G����0�V���~vguT�F�	/";kX�]4�z(*�Y{,�TW�X��͂��)�9�qR#:)OH}��w�R;�v���--��T^���i�{ui:3��$O/]�9���2��:�,�95	s2��y��M����Cr��MfqB\��;&9���_5$�ݻ���
U;�G��I�-Oj3�4z���Sc;Wf�|̤�Q�[�F������G�������ܣ�r~FM}U���xw��A�Q@�t�O=8�Ŋ��WvN�INµ�3UW�[����p�FVl�a�掽���,Y�x=P�hz�YE�_�Y뼻�>ɚ\>~��t�#���[ؙ�Ȫ�Ƒg*C�.Ԭ�=������k'yxg�,�>[g�cg�8'lz��fiC��m�Z�k�މ��U?��g;��$_�9�y� }�PN�zs=i�T�ju&�lg��x�I>TX��`u=��?*za1ƢkD�:0-�����8L�J��&f""7}��E�F�8�U�a����Wm�tr���L�S<�q�ݧ�t���-�j��<MAmt�jC�D�b����;�7Q��x	PIt�J���Fǩ�����F;?:%*��0p��!ݵ�a�o͟ U#==�
,��߈�ti��:�mI������FK5m�{U� v��SN��wz����U���$=��i��0����<�=T۹���K~�zv6�t�;�]�9M|U�����>��j7������@~�����������ŋԟ�L�x���t�蔹���-��ކ�퀵w��k�����Κ���3����Ds��`�._���+�QÞ�}���ej~u��ꋌ���9�Ԫ&� Q-Az�q���.s��4n����Z�sT�Y*�z��Z��l�K6��?�V}/W���L��3"�;�����#�>����I��5ܸ�2 @xkF�Wt�g6�0k:#̕�;�7�u�gv��g�i��;˸׶|^
�S��e�GU�3���]�nC�^P��ث�D��w���7�w=Z��VK�n��f�˧ ;�齊�$�=��9����a�-�K]��V��B:-�3��f������+�1u�XWol��$j8[p��K�k����E���9���s�д[J;���pZ���l�;�N�;�x�X����C��&y`�0&\w#����鐚��jE��&�Z8LVY1�w���[�ǂ��g��Qf�W�V�Q�Vv��a�J��&o9�|x8J;���g�o���s�v��3�m�f]a�=|�*��r#۪ܬ+m0S��k�G7�s	n>��M4�M4�����������;my]R�vY��9 �=:��g*)L�g���z���е~����sSN�W@@뛊0�!�����2uRV1�33�g���4( |�r�~��۸�n���v��u��ڕ:�v�]�r=������F�����J���	i�fj�:{��N6�u��h8�v���*ʶ5�u�Gnd8�^�-$��Z���p�X~g�,���d�0(�|�ja�0fbMnR�P�Y٦�[���J)�6�X�NW H�px]�hs���8��	Y#��L��k��uu�'���L-�W��(e�fv�#x����醉�ᔅ��FU_V�k�D��w�λļ�2�C+�<�v��OK�H��ˈ�$e�����\R���ҦB[>��dS����t�5����Wݛ��R�\ʊ�B��4���1�1mV�$����/���H�>���ȫ���%����G#�
�V��@�-��M�w���	�	w�]�����f���f\i5X�ty�2x��.q������~yyyyyyyyx9�h��)y��{M�z�����ve����tn�=�ܹp�]���[�j5��4ۊ���5E/��+J�@WJ���5�7Dx��5&�[�\��Vd��(�oV "|�4`!���.�~�7�������b؆��\�Ni2(כ$��#�9M�S�tG�!�t��
�Wo�Ckhk�6f���ֺ�]>����\��Ϩd��s�X�cG�5^�x�R�oĩy�װ���q6�]�^�N��Qhfp	8H���Ə�I��}�i�⧲��[��fF:dm�V���� �����n�>��AYy��K���h?W���:*�ю7p��k33k=f,�7��R���on�z����FpO�uR#�=Q�S�%�})��a;y����+��[Q'^%����&�x9�7N�O�	=����������8��+2�yik�A��^��eJG�����2񙙣������ް��d�k��큦a��m}I��^�N�m�R�N��"C��<�����Ewq
;x�sut)LyB�T�WhW�k���W��#���f	���N�]�m�/�Y�3jU��u=�s�WN���Du@��G�N�ND�ܛ[�����fN����i��ii����6^�_�M��Wq��4�Y�����4M�\�ȶ��q��t���ɢ���%^�䗉���ڷ/ϔ�����b���`����}U�"e�ح3 �t���*�U�x�L�756ņ��9D���<���P�r�����f_��-OO�1H��T��Z2����=��W�}[k��Y�y�30w	C���r�*��c{Q9X�uC�N�=�s�Hǖ(Oo����$�W~�{\8��g}��{Y�*��
��l=��,��xl��;���~�O��co>~�z�����1�r�}�_�n��m�~^�;��ڐ�Y�YR7b�'4p���d[٨ɫ��^v`i'��DML�����qhޚ�	7�M�yi3|c2]��:Ŷ�U�3/�a���0�Rk��R������[�2�~��_b��6�"�WMr���*���>��fإ���ੌ \��D�A�R�0��ɶ�!X¿x2<o�1�wz���^V��v�2;;�IC�X�[\ez�c�gdt\̑g���:t�g��M��2Q/��^^^^^^^^\����0'�5Ӕ�*�}78�y��Ǭ%�\�]���"��;��Z�˭�j	�/rX� ��vb]�SM�?��C�a������qd�q�u��=f׫�I�*�WtHu~J�l�M���n;����x4�Y�z������l�MH�OrR<�[-T��������sUfrR���Zx�c�)͵��vx����<���)��gkf�k�=+t�Q�C#���@��S{��U��$�:��U����ET��P�%����n[�Tal���K3���Mn�?�&��b~��|gjzA�W^ft��X5��-q|f���8�n���O��|�dȃ�6���*�3��]kj�4DC�FZ�»���p-�����0���3��^ݻ��9�H�>#����*�d���7�S�AA5�g<��FK���US�����}��f�q��Ju�	�����bD�l[���3��t�Y�p�ʽ�M
�$J�����m��,�}3�^Y�8�M��r���/�y��en%����L�7�Yȣ�'%R���v��M4�M4�O�O�μ���}�~�{_z�)Ğ3�ٍ�nI�hL��Jy��8�ٜ��~#g�k?Vڜ�O�y��{�J �\.gD�P�R6C=�u{+��x��J�0����4%�H��%ў��4���#�ݖم��^cI(ٛ�79���P݀�0�w
�8wӛF1���_o�/I�Rp1�<N�H�f�l����vv��U溛]&+3L$�#-����Hܭ���p�"'Ǻ��1�y��p�]}�/�Nn��~һ��q)#�o�ξ�ܿU�-xl���{���;n��6۝��gUE����o+�
��)��x�������]��!��P�ѝX���v��2\�g
�u��v)n�GwPI�J��6��U>s�uu�uEiܕgR4G3{F�_�C[{/]Oo� �vBr�W=��H��6��N�*i{sb��b��6]�Ӕ*ѝ�O�G܏a{��5�q<���WKk^����HtG	w�b���jŬU����egB/+t]l&-���	��ZŸ(��,����l�Ɨr���
'�z�]B;&��x����Gi�ŭ��Y�t��x�c��t1Д������7�dm=V:³"�����J�����m��.�.�K��Z�V�S�:V)[��8#D��M��A�����C+.'��JN'�CL\9㌘��Y.)�G��ͳ#L= �k�UA%���ڗi�D\z�h�є����7ݒg$�3�a��G=��v*JM�+[*��C�9,nI[��f�,���Y�):���پ؞cIV��h!��n��.���b� c1����rg:�w�[B�ޕݰ��xf�e� 'r�gO��>�4#sgi�۴ij]�v�;�J+Tg7v�����EsQ�XLn�i���e�J�.��	�ܪ�p�۷}�^a���ڗ6���ܲ[<�:��O|WB2n���h!����qE�vo�h$�vԪ	��k:��Q�=:o0vX���2�,�5z�L�U��_�����Si��w���v����ʻ�GQ��9���7���Y��v�;Aǰ�U��j=���V�IP�F��b'���$/��,�7���PC�w�աH�i��Ytl��a3��56�]K~$�M��C.&����&�@�q��E����f݄D�MUԩ��ė�IV�"�'�O��C2SqN^��K`�����ɗvM����J䩟oE}#��ܛ���"{���6�C�P}��"�A�Ð� �3��Uԅ>�-�݀��>�N��zVL�W�c̝c1EӁ���l��eξ���䆳��qd\��/\J��r֊���QS����
�nh����+�=m Lc�}s.�����ky\�d��X�Wz��1�S�B�^�����xڭA��p�po,jC��D��R���!�xҨ7yK�Uq��s�9��^�i�H�CCS`Qc��k�ִ�����q�c'2~���9O��i���k8�$�r���7�9�m>�b��[C��fv�X�U�Q޶��jPw]XRb���k5���t����_5������z�V@o(���W�9��
�xN�.>��8�\�AM�h@�C�h.�vI'5ᜇ^'�� Ʌ_1�*�m��*e�E��B�vX�R��\V)�$X����J�#4��l�N�����e�p`@�����^�[g;��d��v���Ty(ok����c���G*��t_l�j�2�Yu���X�T�4��[�����=��y�QƭIuΈK4n�X}@��ϴ,����O��h qD���M?�*�\�9�:Nt�΄ˑ����C���Wy�I%�2���!)��q���^�]i�]u�x���O��I<�A�!	?z�Ӵ��}ɐjH�$�=��Tg^�q�����ۮ�뮺뎼x�㎾��p�D�i>ج_�$Qv]��%QY"l(���HAwD��U*�}zqǏO�����N�뮸�Ǐ8���S��IEPȲwIW+"J��q�+P�
N�y\��F�_^6�ǧ��׷]i�]u�^<x���_^ö2�"wE2m��,,".(�����\"��I2���\��%ˏĞI�;�L��B�r���w����>TE�f����ˇ*��s�9
�g*��#G�||"!�[J���HUAW(���P�?�K�_��������y$ʢ�'2y�Չ\y*���+G�aҊ��W�p��F�Iwp���8Ty����y/��p��R��.A�b��*�(���}7RxMsnI�C�r t�Oap�D�\y#�Q���.{KqkŔ^��z��x��U>E�|%����.��&��㷏 L�E���rH�[2I�3��8H|r�T��G(f�.m�.���9¥���(r�U1��2��s+��s][pW^v��7��o��̠���
�DA,��F�p�'� Ȏ(� �D��$*!H&S^��5���o{�y�y��ʾ����!��l�<���|�Z�
�aq1�,3e�H[�xa18[�2X�����D��q�F�i)�Z��e�[�Hч���I-������������U��B��L��Ϩf��>�^�x�N�K6��z��,7ˆ*bl!�Z���Q�ޭw�U��_���ǉ�O���,q��([�̹mM���v���$�lw��ă}��V:���z'�2�K��)���$���}�o�dGzT�p;����S��1u���{9��q��i�V��`�X������}|�iS8��������͘=+#�1�@�p�!�|�~���3�,~�_�{g�Զd��/�m��E�[�o@p�̀��C��
�z:Ո��u&<��٪C�(jl�E��'4ćc�h\7��kw�;D��B��]ݵ�,hGt�U�ծޯp�BndS�00��#���z��oz�Ɲ��t�,�.�3SX��e����he%��R�[�)���/�ei�:8����L��U��N�yK}`�-������30�0�5`�W�7��(�u����r�[2�v!;5,��;h_�f���(j�5��,���͕y��£�T��4��J���Ifc��K�I���ז�'�_G�:�\�ौh������N7������o7���h�P�޹�U4#�Q��n/F��o�0�;��:��Q�z�fn�*7{��-~��9�H�QY�.���D�*�����6}���JS�4�x��p���{OwN�ۍ�~�0+��>����)5Mϑ�Y�.�.|=��Q(6��M%<�6e�Ϣ}��p��a���̦���ӌ12��D��+�K�|�vzH��=��9ݸd���ڂx��:�ϷJ O^���L�#�2�,������y�ϨTZ[%�矰ۆP`wG��BI}���޽s>��ޙ�=I�0mޢsek��M�3�.�_I�K��M{��cڃ���ΏR�lW����)<̞��;U7{+5Q��oD�{v�gll���}�=Ɯ�K��r��b��orY[���Z��D�f6����F�X��`��"�]�גּ����e��5�T����T5��;I]�b~'��A��_V��ש�ŰM�δr�u��L�Օ9UA�v��6@ڤ��|Z[ԺYY��q�����.�g�L�7k���5j�%�d^N����E����Ε;A'�{��_����� Z[��9�v"�G��<ad)��6��.�p;�.��kj��;ƔFc=�b���H��:��[VN4��'0�6;DNڈ�<����opzޘ���S��[B�`oJ�(�����ࢳ��uY��o��=~��9C�J�A�<��y���s+ܽ�(��n�Ѻk�������Z@�P*%���x-ŋLǥ{�q��d1����:;N#>�5�)Ζ�F��<J��O�d�.��s��痪��9�!ݯ�����W˧Β�ʏvm�@��~��Xk�Tk%��e��v�o�$+Ӯ:�6#�`D��kֿ�U:��PgH��dw��y� ��m��EV��x�vl�8]Ê;������=���UH٫�Rި��_��@�u<���A5���;��*��Y,�3/�Pp�z�ړ��s a��ev4�/,R�KE�FuWJK���̻S�W�D2�n��V��������6���C���X-&�}���ڜ]]��(`��Q���t�
�ˏY�}g	�����d\d�rD���a��o7����y���r��WzK�
X� ��g��mol�uμ�wF��x�n�w������8{��y�pA�^��ޗ��x��aO�Ñ�9��� j��'Z��m����"a�0��`D�H����:O�-򷐨���U�4���11�f�J4I�)���b�/��=�; �d,����ۙ�5�������Z�`P����n��5`����'��{m����i��Q�z�Y��<���I��y�.���RR8q���Ը�,(�ϳGH|_L�E�mc+��z׽rv�9~H��tma$�/� �|��.�z�Ӛ��ءxuet��D��qCv��S��>	�Bn��w�f�>k,GMUtU���2N[^Q˦1�?xS����� M��(K9���^�#,GE�����UM�j F�̻:��sm<n8`�I�m�î��v\�K���`��K0�WH�|x�d�&0�J��ف1z\*�XgcV��_^� �+�ŻL��N�>�K��y�P�Y��@�^R��kF�p��xk��Y�M�Y��T��n�]`�Ӥ���0S����U�yS|��7�*?a��c��糷����ՙ{��b��g�f��%ֈBX�X0�[tНz�L��m���퍿�y��G{��=����nɨO�l���ݼݥ�3��x����+����H�`���Z�1�%�*V�ԍ��u}���y�lC3L�h�ڣӻ t.�v��V�:��{���m\�LP�d� i����~�;|���?nw�䑖 ���W-��,";�Y*�#Kz��v�j3�^{�����;��&�17�)i�}^��7�7�w�3�����W�r��5Æ/3��*7_c�#�-d��w6����])�C��f{�CnLl����l���(G���0di�<�wFT��u����j:�R��1�.Wk�2$���1��^��<��8���+�S��ܶ˙�[�OU{�]�H�Xz�#w��vt'����Ϊ�л����#9�63ّJfcgDfOV����.4�(v曋���]{8��O��E�t���.�w=��u�{��(����wa��mΣ�c�qjd��x���&̵|�Ռ�VEG2,5ǥf�}Y ��|`닭[�({}������� zr+cդl�3j^���q`��#e�\6��+`>�:�g��;ȕ��;Oe�k��/9���5��WVŹ�`�2~�K�T���	gw�h����M*���5O��oFs��`H�2�S)�.� �TԺ���q��cl�`��=]Wg)�����zH:0´��8t�眝~��ꫣ(߶�LW������ff ��qߚ���}z�I�w��жd������J��	����O+�SG�>'�l�j��}	%��D;�7�"q6�o�������O�-ԛ@���w��@�l��Cxz�L�j.�r����zTA4u�<�#���5���pV�Wp����:���t�y����ve3��U7�.���'g��ՏY���=[��j[yE+Z�)#�η�c�R{��'+��w�rk9�t�s�\��,�����w��4Mȯld�`G��e�����-�}�7?hsjڼ޿1�>�#ā��>�Q߻\��w�tŽG�RmM��e�᳹Ҙ�f�ʉ�3��)g[����Ζ�[�zt�߼<8xxxy����ͯ����"�)"
��_����>0׾�^��[Xb��.���ko��#�u�F[��|źmn�t���	ko0�� ��q���M*����m1l��쎎GN�Zw��K���� e�y�-��{󎶽�$ռ m�&�$N��N�OW��H�X��X�i�Y�w%2�Wٗ[_տ`3t��`��s���Ow�z�шW\n@
w|9%g���ݒ�����f��:;�9M�W�U�⥜�oռ�����s�c����8���5R��u*/U!�ހ�LML�q9u�z�z%�6�+N���S��G�˶��?���Uz9EN�zP��[���zw[mCU�wr<��fm��S�@��xw���9��!��哚��Ü6��p�1t�tٟK���;%��ݞ��_�[X[]V���gM�?��U��H�����0cQ�;(⥷�0�����v�V����s�N���!Ӯ)7��e�W0�aQ�%�w�e�����@�%"7N{�%[ؖU���W���*��ܰ7����\D[���ι�}�W�����`F1��#1-�]m������O�.]>��|�;e;ř��f�rJ����D�op�-t�y���붛;ܛ�^D
��rRjE���������~jQ��G*��0��7��B�_F���z���Nק��K��\^{����:3x��5��?�qm�xC�Ȍ�Y����@���\2�k<R|�&�mA�k
R�?O�k�36�I��0�dtq��=��w�2;Fc���'KU�f��U��;�e^�2ϖ���u������������Is�yGzz�qzZ��"g�R��f`ի�do��F���J������ϑ��3V�pj$�k#_;�z��#�� U��1� ��M�2��yu��,��/h�z����=)瑝ـ7A�_g1��y��*�(ѡ�z� �gA`%�J��W��H��(m�׆��>�<�2���s2�G��GX���3ͥ�,ɢk�i��|t�&��o}|k�V�����8:�d�넒D�Oa�ڠ��+��=����Ғ���U���wk��+"N�!��sn&R��PwI}�ά��'���а�wߞ��	�{���N�«��0#���`�d�;��)m	�˗O.�sN�}Շ�RL파,ӝ�U��k7�9':�M6��Ͷ�8�|����b��_YȏD`]�_��o#�2��Z&cw'�e�g_0��a�u�&��� C��v<�o��w��L!2�˺S#,������.��3w�� ��G�лc�k�{���"����"�Da�?Gzϰ�Z�r����$����J� ӹۣa��o-���j���9޾�U���|���ˣzNw\�k���S���u2�%�~K=�<�؏N�#�djv���L�y^-�Zu�����T�]cz=�G��7�H�Q��=��!�-��a�r���� ��1���7$ٖL�?xp"�>,�;u�ۅ�R�k��k�)�ݠ'_��Ӧz[�%�k�R��:���.����Q�N>d�M��u���S�1���:}���d`Rϖ���	�Fǐ����lD��q��L��N�?}}�n	�6BJ�|W|q��R�._��7�����*ڽk�f���n�t��-P����V��,,�9B_l�ɤTү���Է5�xns��u�]����f��y����1�c.on��\��������"3�/Ҥ>nx�>�0��u�d�K<��c��r�h���|������p��\�Z� ǾU�*zL3�Wn�,��0"d4Du���q�ϸ��W�v�q�T��]��ǩV=�j{�̜�P�Iҗ7$�NAλ?k0�	��ԕ�����e.V�<�Q:uٙ���8{		��%���3�\�h�궬h����{g�Q���n��1�k�=�O��3����W^�A�*ޙ�W�'Xn���q&hbj�ڎ��)Tފ�z��e-Coh��Ɯ�M�gh�*α[,�9�qn���Y�}V�z[����f�s{���a�,m��f���v5fa��5��#C�Tz�!ю����E��u]rǋ�\E�=�]�e:S���N�y��f:��X,�@���'�w�J;έ�T�q�� �##"��{��v�ft��{�eN�=̧�_��ju���#�$��3�8��U�O!NYY��{�4�;(���شV�m:�9�K�4#��[�۶��%&�������aVh6�иȳ�8�\���ԩhi^��u���� \C��ܙ���:����T�	ofn���P�ȼCF��Q�%I-��Rv�0��9e)\&�����ɜ&M%0E&�ukP`�J$�ݗ�1���M3Gb�l��sn�T����7[Rf.�����%8c�����!{�_-)�]��-<���/�U\z�e��)���UI�CO�U�%Q��A����ӥ
ڼfz�r���&�Xx�� o+2%�:�<1[ :����%����si�,�;��%ή���D�t	��+��t�-+�*�i�q���a��նM��ݖ������T��M:^
��_һ�7o��4�Wl�DՇ��&�?^J)��k����ד#������UH7��Gh��N�C��ha��6Ԕ��d��v3(gV̝/V�M�~�L���P�;�����:+��sԝt�S�{�gb�:Vb�a����to���hՉ��[E�qC��Q����Ù�y������V� �N�HP;�m�B�o:)5T��A������T�J*1��@�("*�M�B����?Y��3pT�#�Iت���������,���W�+����q��_��a�ܔsl]�Q������VԺT§KG 9����2�[M�"]�S�q�� �[[,��%�.��5u(�@�(cH���dk��f��I���p���.�-��K���))�g!x%���CZ���TD(r��u�T�zk��tma���@fgd��֩��6��~��4�YXo7=��%XwjX�r�<b�����p:y��)k���֖8�l�������\d�����7�Oud;1�U�����Gc�V���)q8���_g�,�)��a�+�qP9�9���VW?k���^��q�oL�U��[��=�;OL�4���J��M�W�Pw�n�U��*y�k�0s�(N'����;Wz�\�̮\�e���o�3:+�k8�C2�"��F�9���im��h����-$E���~�����hs����K.�0���6��*n���L�i�{T��X�+��Jt{����"hag�ȵi'2ѯ�H��Z��9��V���囋V�l�^R:���w�"�P�ޢgf���6J�N؍KD�pV�{�;]fq��V�������e��)�&e�Dt�R ƃ<	$K\��'{;
?���G(O��\.G(/�*�hlSZ���ǏOo��>�:�]u�]x��Ǐz�䧨ܻ�����\��I$QE9�4s�ȣ�E�X�Av[��O2��8�r����׷�===�����:�]u�]x����o��{��Z�\���B�+����e�dD>'�uP���HT�*@�>���x��������u�]u�Ǐ<u��H�
������m2g}�q��~zz� �~:Ew�����4d*l�'(���;}z{q��������u�]u׏<x�ץ�$��n��.%r�t� ΄Up�=\:Dr&\���Ap�/���YAG���Q��ȎE�DEd��;�

tR�>���As8_�Z�w��Թ� ���$�����l����*�a�.*�����(��e7�GT���wn�gYQ}���7�$�_�Bc��r�Ys���T>7�)�<�i^�E��*"�E���w��K"���4�TA�u��ΰ�! �G��wEEη�QEUx (x+�0������@�}���2KiNO�^�7��.�,��E��&>�X������r�قU�������� oFն��r�<;��fa��R���{���o�'-�F��O��QB�48�A�I&�����7��āM����	_�(���������[ml�j�r%]Fq"�YBSΫ=�tb��g��;3�6�3�M�z��Z�~c��vN��hՃ:d ��]���g����j�­��p�c�u�h�(�m���8�۝M��p�ݦ�:�Z����zaW��D��wc��5������^ɦq�`����a�rY��]~�U��be~V�Lj[kNw^��q�MP�;9coײ5��}q��;��tL���}�N����K5�;4����H��
GF�6�.d�0��桹�*/K��LLMRg���q��l�U�~��d%!'���sybiH�i٫�7	v�j4���
�㌼�+�,�d���[k�.d�*W�Wj��i��c�y�\�XOٙe]��8���˺L¥��k��#=W��P��u��&�}Q˽�}J�w]�Č���u�s�q�z���gA�cMp�䣝�f�=%��8w�y��o7���:��U-�*��z|�3� G
P�<G�^hs��Ŷ��yo��'pN�l̈́4�y�^�'��ϟ\.���r�4��J�&�X���afp�z��Fd��������W~vw��8�_
P���`y�樈Ƕ�ݰq%�roZ�w<+�z��#w>3Oi�p[C3��=w5�&��h8���-ͨ�s"cҽ��SV�s>^�~f���v��w�^%n���4N���;�o,�M���]�q0W���U���0]ٯ- ��c�	d:��!�?;�9����a���F��ە3�┪j��b��ޮ����ֆ��(�}C`=�q�J�ꉉل�z�2����Y:u��+M-����9�{80jХ�R�fM�ͧ*�:+�k�a�6�2E�p���Y��W�G��{�� �-�f�W�?@`U�MeXo��~��(:Ӊ5y4b�	�N^5AR̗�j�}s,p����P�����?_����}J�g�,(���( �=���={}	͙�j�����ڙB�Y[ʞ�}�m�R7����Xy�p�g��j�woVl�4bY���P�~���� ��.��)�!ߎ�`�7껯��7�S1Y:�H0m�a�а���4�Ы��ܩ
}�o��w˛B�ͣ�����D����)��cۋ��D�t��N���=�u���k�7w7�i��2���=�q+:E︚w�o]�Q����U8b-��\�7nn����$T�� ��31�ׁ�B�0�쁺KQ�Χ�j�Y{�8���ꉷg�x��a�=��bޥ�_X"a��Q멟���0�f��w�c�47������|�Qm��ȫ�wŬ76��ŤV�vk�##1E�s�鷥>ا�i��uoPg��I�g*��ӧӳ�C�	����^#4�	#M����-���u��^4��tBV@~�ZdP��&7#֌I9U��!�gn�w�}o�mqrP��lΪ��Acw���[Ǒ����F�܄��y��Rzw�K�Y��K{�7"����|����awd����;@r'œ<��	���b�emQ�i`�w�M�%�A_�Tkn�-Ƒg3��	��Y7~��.w#[��Yv���7�c��!��Yv�h\�� �����D�g�R�z�Q},ê�-e�u�L0s�|��
�UW��y��o0���v�+KZ��������$�\��+�}"��.�=��j'�&^�l�{�����Lg���l���xxh��ԄW�]�{�Իi�Nxs��خH�����ǽ�ϳ�	���k��k��3}Q�H�8���%�Vz�n����
��S�����M��9�LۣY	�t��S��O��o����H����e��&�Aq���:&M�����=0+˪��W"̦��^��h+}ղ�[����]���48S��3��VBU# f��}�|�>����\R�jZ���)��4kp���k����	�:@G��{vp8���[k��S��dk�V�à6�z��'		����� XK �[���uv��:���{"�O�`#7|���oUz�c�2����^pm�Z�*L��
LE�Y�'rkl8���(4,=�;�N���-$��+����q΋~Q��A�h>Y���C>�1Q�s+���m^ۻ�AK���f���볡D�׆������B+,�tu�d���!5ػ[٧ټ�A�m�:��<<=^������:��Ps���DX.�ժ�tLO�Q6DgI�#�a7M6�	w-�J�ez���
AsL���<��wD��cճT���[��'Go�����nߝ}�y.2�.��H������b28�'�H�I��TM>�4��	��?,�ٗa�*��g'��Kv��׳s99⻧���kh	~�/����4��a&�:��R+_���^�m���k�7�w��7*�;N�_3s�k�����FR�GW����u�+U�9�퇱�ZB˒��xx�Xj��Y�/����܆�~�cgº 0������`��4�wp�g^�RG/^^(���x������bh�gן9yx�jB7����k�o`����wv��ɞ{3�t�ݳ�g�*�i��_f��#��Z9��tݙbp��Xlu���N�s7>U��}����}m���k\to4y��1)|����Vs�ܜA8/��l��w	%�QS���^7}���0K��I�$�mu�c�-��x��7��b`�'k�u.�=�U1�b]|s�g{�o����������&Tb;Y���m�`�n�۲�5muڍ���$��8�J�QG�E����l����
0C�v3�񸨛uZp�lw�ݗ���y��~�#�ϓ��nA�В@X8	���Wk��z3�so<�!��{�=i��J��.I�p������^N����ضqfQ�]�N�Y��3��{��S�ݮ��c���c���댒��0��S�o@�@z�4�L�X�ſ/t��s;��A?]�%Xb24�5n��£�C�I�:*c'��f�%cn��z�C�gk���PHw�����NQo'i�Bޙ��m��~�'C绞:1�!�4��d�J�.��*���걩���{��YRp�R9���`L ��7���~�gR��O��3ϯ&eZ�9;�wZ��IZ�Ase�ոG�)]�鎛%ǷtN����ǐp���i��ln�C,S�9{�{������:�����}|����w8<��o���-�<I6��SZ�e�Yܾ�6�w��r�����;���1�c��:d���]+���ݖkN
���B�3	;��c'�� YӊevJ�@!Ѕ����Ϸ:�X�[�o)��wrm$��n���:�RH�]�0�=�P�}�\;�`Du�`����v���4n�R�d����8#�C!��'�aCo^[��Y�eryi=՜d#K�w�?o�q��/�ɘg<Ӄ�����zk�m,��c�H0`f���k@�������4�3��?i)xO��Mη�����I��7���������O���ܕ+�[Ckz}�l���΄|��90�F3T	:���r�P�8I�}r��NU�Hɮ>��k���dY�M�Y��(S�6=ȓ���*�����*k{�6���7o�ㆾ0�Ԫ/�ؼ���
��f՞����>�CJR0�/�Pk�9�ǂ_������`�{�EnH��q�O;��Ԇ;�^&q�a�X8�tÚjP�*�e<�E��{��qǏ�ܛ3�G&��{�;��vnfe����|@e�ؼ�Ηme	&�m�Dԭ��'���3GS��Y.�=����&��f����6�m�c��ZM�w���� �o0$���*��D���#tʐ��H��⡛�t��r'�A�Zq�0��2����\���6V�l��]:�(eR�ͺ3���Z 3�b���o78nn\���[����]*�aʀ�|Ӥ�沔t�{��l�۽�75O�W":p���+��i}6�8��@n ��k�Ґ�\�L����{�g
��~����`�^�l�tk�%���nF�=H�����M��jGw�ػ[&2.�e�b1��0)�S��餣�f��&�z����!�����X��v��E,>��vF�pH�b���7�	n�a|���mJ��[[f�=���yK~ZdDj�W�e���\�=8ƚ5橵�����[�����x�=�0���� �����[�����^K*
_G躝�K��i<Yگ<úRq�N�h]vOF���@�+�f=L�Eo�2B$d��#$p�|��&�t�Z+�Sښ�VZ�=�;'#�o�7�t�R�f˰�o�x��tJ�g��):N9A��xxxxxxmf�0`����`L�p�{�<ϒ�9Q�35�b8��Xʖ��2�Z;W�����L�٬���t�3���C������Ή���oN�s'T%�.�z�#���m�9��2[b�m���}�/R��n�NC��^�˩��U��5�-�3Pۅ��޵�����:�a��{�bGj��F�xL�#7�=��@]n�`FQ���w�	n��im��s�3�X簶�wUؕ7��uErkfm{�֧g{E�$H�cI5��n*%֊:}R�yс��aGNƉ�qti�v����(ʨEz���I�x�wn	��&�{�:��[�M����8��É��X1�a������{r�cI�Z�N\]H3q�q��A� �>���dQ|u�fx���j6O�2��򛽬�^��
�C����2t�w���M21�K��{*u8"�W��Vq]E�0�V,�1�·,�Ps��l2g1�5��3-���=!7�GN�}zf+;1)��n�62��׼$��t�ӽ`�ޞ>> ��=]%J��O�ڧ}1��m_z:ENǨ��J�q��~�x� ��7�F�5��k�g��F��8Z#k����q]'�XC���q�im�����nG��d�I�;O�m�=���]�_�l��6�4m�e�����70��2��/��ү`L���Of�	�0�5Zi��1���������;%�Y�*�&��t�߳6�6<����M͓��=u�e�>qpFg?R`��K�gc(�Y�Kz�4O6v�KZ��s���H��\���^+=׷S�_���,sG��I��ǌ��]6K�4hj-P.���w�T�Ro���g�>�9ͱ9.����wN��u�vT�z~�A|�J�'��� {+�o˚���[��o`�r���3��<��%T�����Oz��?� U���
�?���i�H"�������YQ����`FS? �g.�2cgdˑ�`)�0�L���v�!��r�ː�!�!#H�#H�20 d9r���ș� �H�2Ec���R � �H�RX�!H�21�B0D��D@��B2*d �0�3��2hA�`���a(�F��dB ��FD ) b!�@b���bD 	���@`����@b	���2ld�8��1��B H 0P�� 1��  0��HD 0��BA 1�0�� 1��B 1��B �HD 1D��B 0��BN��p�B 0P��D 0��BH H 0��BH 1D��B 9TT 0��Q 1��BD 0�1�� 1��B HP 0@�� �HD 1��B 1��B 0P��D 1@��B  1��B 0�� 1 �1��BD 0P��BD 0P��B �B1EB���4hp d6 C&06  0@ 0@ 1 @.��@ 1@ 0D@ 0�  0P@ 1D��@ 0D@ 0D@ 0Q 0P��R!#T.���e2c	��p#�0�vH2T 0D��!�cB����3�1D� �Bm�S"p ���0�Lb�pa��H`�1��X2@`�1E����Xb0U�`��B��T#" 0U�H�V2!H21V1D�I�������� 	E H�FF������g���@������!��L?���?��/���(x��������~~u�'��� _�������*����@W����?q�C�X1��S�b���?c�P�@W����'��-��__����?��'����Q'� �� 	(@�A�� "!`	 �V
��*P�$H�DX(E �* �$b	`!(�F" )"!A�@��@"!AH
HF
X�H(A�@�"!����
�	"����H����� ,"�" ���
*�QBDBEDBABP�A$"E@�A#	�"`q�0��9b("	�A"!���@�@H DH(@H�D EH�@H�DX E�B"V""V �F"�Q�$@ �������V~��� �"�
 �H (�����/������	�������w��@Z�A�?����"��O��C����8��I��'� ����R���� ~T ��A���~�����DP^~���DPW@�R~��%�qx6����W�Έ�.>�p��, U�����c���?ۘ *�����r�?�g��������?xf��?��D����C���@WO!�HC�?h ���g�y��K��(��J���?�����9���N��� ��!���)��;�a���}_�����1PE�����q���
C����PVI��N6���@-�` �������O�/�+�5,�#Mb��)B�&�h-,ȕPk��P�[&� ��(*Z�MeZ6�"l�-QM�[b��ѶȠ��)�IB�U����ūi��v���vm+nշu�-�lr`[%U��;�kj;+1��r��i��M�Y�+X���d�RGf��Jō��vc��m���t5�B�)4�m����K!%d�͚]�Wm�����Wn�ȶ$͵c�L�6�a�a6��J�rui*V��m�mm�Ħ�eM�%Rv����(�m��v�hԬ�j�  u�>��j���X���]ۘ��[k��v��{�����v�^�^�ۻsRN�9��̴=��;�Uw��7rW��yG,���]�k{4=^�󧽺�N�Qwk�]��2�j��JZmkn�  wn$|�H�clHU[5�}^�(P�FE���D��e�}�o��+�O�f�p5�{n�M��{4��mݻ7W�׻<��m�g.z{��@vŮ���vފ���g��zշ=�ײڝ�٥�������2|   7�_l��n�疵m�U+p�v��{λ��Nb����۸��۶������-L����ݧY�K�w��Ol8���ڕ�k���Z��K��cgl�i����n(�;�ۮ�   ^��SZ����z�մQ�����Z�̯e2�����[�OR���{�w���D��W�J�v����k�[Ca�vsx��We\����W��z���ke����&�#fU��   ��o�������U�{�v���o��۫��.v�{ު��b�=�����Y�{�ݱ�Z��Ow���Vu�]�{�ު�yoez��[Gw���KiKA��ԧWnWw�  �}վ�uk7V�UDw:j�OUUz+˼Ƨ�����vw{�jk���<^���  0��m���p�#��� ��.�S-3f���f�LYU�   �| � �\ �;�nt= 3� q:��  ]���  <�8 ;�A{�^ � jz��� ww��l ��vڭL����v�6��v�w�  /y���zX��  Y,P��0 �o{O<  ���  Gu�  ���@ �z{�  {��:�
n�QD�ӴY�B��i֥ۜ��  ��  kiӀ  �j�
P����x  8q�� mt�  iiˀ ���h 4�wڅ]�x� Z�m�ڵ�Ķ���$˧:�ڷ�  3_)� }�{��x �'�� ��{ۻ�� ���@����@P󼻠  �4��޷� π"��M��* @S�0��� �)��b�IB`d4O��T ` ����T�@ 	2��FUP� h3R���������Dڟ���M�Bܽ3N��֤��J�4�ֆ;�A��e%sj1�����|��ק���1����m��?��61��y�lcm��1�����61�O�  <�LHW�MD���HJ�+��`��VL'q锈8(^�S&5$��Ӵ+��F�pi�}�1�pCr"]��w�B��Z��)j�����]c.|�퀪i`U���m�$��6�m�sl|���6���$�fO�7QK[�2�"1u�G���[�n���wKE�.R�:ݲ*�Փ7Q����K�����o�Mk�.Ou�/t�x�a���45��1�b����#�ن�&Gz�,�X�f¦��`��[n�K�f��7w���i"4�*�5cf��&%$	gLx)��孹���7L ��tY��Z-��5��V٢��w��f���n��{�)�i�3*�&�(R��(�q��P��K���{��z�}���!Q0F��Ѕ�*�&�Jn"�(<92`o���Č�!��)�d��qű�3��:	��q��.�Ȳ`�$�`R՝��f�����iK��CEij��Z��
�P� "[GV���2��cv���L�n���V�̦�B!���x��
�<&�\V�.���4g>������)=��K8��k�E/[ѧZU���
��J+�mb|�ǡV]��r�H*V�ӫy��/�����f
M/�8r�%#JQ�!��ûDJ
ѩZ�9q��t��X�Y��Y�[��8EH��v�-k�*��aS+M�ڊ�R0ft��j(f�e������-|�d5��W{�4֖ԻVl�a�wxZM�#��C�U\8)ACm�	]d��*r�4������&Bz[pf^0�aO2+gU�Q
�|rӷ�a�x�W�����i�n���v��%��8y���x�qMq��ё����I�����&�F��R����n�\�h�U�BQeI����حa�y�5��2�2D�z�;�f˴�DX�V"��:�PN3������p�v]��$7e�h3�Vs-:��m r<�Etp7Wh���c��ۭ�)�Y�
a]�_n����@Z"���I�Xf5D�#Z�FX�nֽ3E�ϖ7�C�3Zf4�(�Xm�S�W�ش�+	�{�]��3V�+3GV�!O�u��F��i\N*��E[o-���^n�ChA3]6$�N�PM��$�CJ��^�;{m��sV4�S�Z��Ho7�����0$5V��fimQ���U�����bl-�)Q[k-�L��d
�X.�ȶ�A�����,5(L-�s4$�.�U*ӓe֩r< гo�ً`�ùn�@!�o>AͥJEP�R��U�f��8�OD��E��P�u�j��9�JEлʛ�+C�k�{(<M��{�Һ�u$��n�
o�2d�f��3�\ �H��N"+H�kQz�٦,B�-���6���{���ٰ��ƭ���`䆦�L7Mˈ�4�B���@�{(�X���;n
:�in[��b�9h�Zn�I��[2e)�SpM@q�d-��)=�}Q)e+�L�ؕ!�Ih�J�`<)-���%���w'��m��ppj�X��Y���*�m2rQ2���4��X�6�U��2cɦ�R��[p�N	�ךh�9z��b��)�CKF1Wzo-��1\ڨ�P�0]�pJ)��mMh<j�;kV����B<�W���-��E=Heb�5f꺛����бq����Y��@�4�fXV/�42@ь뎞*%�r�R3�Z�^�f�m�d�x�Wa�W�K��ӽ֕-t�ml��h���b͒U���)���֯��Ҕ��f������0�5�SywA"]�	�+bu����Um6Hl�(:�|�bd�W�_�n� 8��WYj&�<#Tȭ��(�K#�T��;����h�cSx�}�B������Ð"����<@���z��@T*Xܰ.��;�ӥ�V �Ȩ&��7r�Ma&����NR�T��D���b���[+�V��E*�,U�ø� ���SU��rP�4��`7�X��e
��4��H�I��t��e�8���NQ*3���&��u��9y�}�ъ-V���\4+yD|i�ݝ��Q��i],t�-�X�cK�@ݒ�c�"�#�wR�]�/b��91S�R�uq̫u�����j��P�����z�xr����u��w�k%��T�@��Ď�bG-���nV��]�V���c�R,��1#��b٦�<�ŲLס����R�by{���g³]�*�u�ƤѬfe��fČR��p��$�EJÊ�*Jl���+C�v+�[{�m�*H��gMj�+!g����p��CCkS
F��c)�Y���Z)ѻe�X���r�7�@ mDotN�Ʊ�{6F� ;Y[vm;y�mJ2��iۂ�
������k@��b:%=W7z��8"ّ[ni`�۔� �Q��wR6�ř�n^�1Y���
�Yb��*���A1�R�4�Ov442�Yj�[�y�ӂjg�O"<�%糃�ϵF\Ĉ��X(�͍�X�n�% Fi-��D!�7KH�B�� Rnf+Bl�T�k���j�c5���Xjն��C��fjwA�)j��NC���e���:���֚a��A��hl���GX�d�eh7`�����E�Z�J��UZ�nH>r�����ݼ[m!���ٵ�)�� c�
�c��FTgM�*L�s2�����`=0�����E[nk�y4(Wۃ�q*������WbEm�P�ܚ�,V�4J�q�wc+0bV�:�K2`��3*6v�H��ó� �)c� Y�dU�b���(^�Y��Wj�ani'��
��ѷ>WXU()��lS�SaY�I�`�WC�zڍ!!#�E�IB^�[�1�r��TNk���iV�c��H-eh��
b�x��X�^�4�1�u��Q-���3x�.�Wf��":ފ2ۥM����P^�İ	�5��T�sE-GD���"��!����
b�BU�ɲ��,ދ�ZPY&KR��~�h�S:���b�>�\[:���f48���A[n��F3{yT�,YZ�Ts/A�~�DD�����7]�Vb.SlPcp���x����8�/���h��=ǜ����%��a�
�5�*��3
ߨ��&飡\U�p�i�#M!�퀡G-�ЬH��͢�h8FD��ǆ%Opf�iIi��v������s��V�4jځ7B�.�e�n���R�((���t�a����W�4�!��X�4��y��I��i�5`f�kse�Ԇ�w$.S3(e++@$ԑ_�^Ya��6f��`z	��"a�V��P��[O/Pv��ަ� ���VR�y�J���h�Ff�{�m�[�s��	���H�f@i�/r�����.���N7��i��J��и ܹ�/C�+V�hf!I|��L�4Q�n��6����b�v�+���V�mf�ԙ���e�G��T]���K]����RQ��˧)�,�B����)��fXא�	�[���N��"��dS�����~�B��wZ%)�ɷ&i�R�1�D��B������QiW�S�jPN��Pv��w*G,۫��i��PN�ډn��a�Y[�-VӨ�����	fY�m�kK�p^����8�րm�ƱìnGj��J���-Ch�M|N�`Y�q���B��v��~��j�o0�gBD*<�^]ȖZ��tK��i*�w�+�Z�m�޷�0n�6�x.�[��@u�R�'���Q����C�lW[�L��Z%
h"���.�@8���3%�dͽ�A�,4�vd ]
ݷr�N�B�Z���r=�BTդ��Y n|d�L��@��4��F���,iMejY*g�j�eJ�&5�b�b��1�Ն����]��jL-�\��Ga��Ps��>>��⳦a�6�'a	ZZ2�W�:�A���\�B����km@h�� ܬ?];�v��5Ga����&нz@�D�I[z!�Z�Ka�QXfa@t�mͽ�m�Qt�蛦i�6�qf/SM�N��;���U���r�<b��$L�r���X���-mG]K�pғy�;j�f�=�rY�7	͇8[v��e���J|����V�lls�L��uY�w{
���x�	�u��qٕk�M@#�+qV���A��̺�W�]�Q;��B�T(�T����]Ѱ��m�ˤ��JTԬoQ�Xs);2E�M
̋��Ж[Dy��d�$���ff�<�(5�h�����ՠ�F�Y0֗@X�HY�FƁ�i}wjݤ-��J�lM�N̹*,�W��n2*]-��oIO��ꭶ轩��nJ�s������PGc�l�S�A�")�2R��ը���.��:��gb�X�e�"�5QA�%PV\"�T+"��	f�ʌk��<Xh檥Za���piS�n�35�Kq!��,"F�Xo/.�Z%%��֍�&�f�쫩7�i �o)=�Ejo]^aϴ�n��m(���zi��Vvi[v�6U��`V���b��Щa^Kk�6U�b��֍*B^4�M�����e#�]cL�Q^�t�9��)����?zy��s�� ��g�;�Y�ב��QU�=x$n帷 �	�p�˩���V�4�;��<V-$n	�r�����i����
PlkM۴a5V���Mv^�V-5��la�`n�^���*���o	a����%�� �S.��������ªZ��fG0S�0M�,ڬz手��"������֙���3tmb�ݨ��-�ب�d�@����L7��̛v��U�a7 �V�)��:���аP����;b8�ͩ#�F�R�9���BA�v�� �A�Z�C#�`���I�k�+J2�B�Qz�5T�����Ւ�擂�e�'.��w�n�8��#�t#Y!:��V4j]m�{3M���Xw�Й.,-���St:Hi ��a[�f��A��{NMPnm�i�F��^��P&WŅ[T�Q�$m�؀�\�V�,��1V���&j�+1$���It��t�w4��������q�h'
����R�W+{M\%?������t�Ę;s�O`�ϷI�.,Ǉt	n�q;6 �E3f�5dL����mG�)��$@�T�STQ<y�VU4�݀�pB�x��]�D]0�f����PU�)E �l;h]�Ň%v&�ɩ�֊I��ȵY�%b�k�C���5�Q)�L�3G��F΃��?=��m�a6���� ����h\a���j����Y����L�m��93r6��%�40��6��ʱN "�ދ�ch�m�֖�m��CMG��*�%K�-
ɉ,��S-���i�e��r��,I���g3@���{Z&k�7�m�B� �ܵA�"ݷ��Ol��[[�IGv�1+Y��:�V[H���\o5
v�֕�լA+��JslO_�ӧg�`�E�@�ܚy�Ղ�[��0%7i�)V�%8���|(�8&�[PV%��)R#T�]f䎕`�s\�Lz� 2��xn���V�k��T�	'BޓW�Ws*iʰF�G�;��������5����f�HM�jM�D��%A20�d��6RlUư�7xM4`��<I�heh�[�i�q�����X�썁��2h0�RT�v(�Υ<˽��8�iܺmWs@��9M����`��+�4�	�e]7z H�����`7��s�1�=�Eqnƒ�!2-:�2��`®��*����jV ���e!旁�F�Wm-M)X���&л�BT!$67Qn&�iV�h�+Ck��]�eHeX�.���W��ԋph��� d��y����;���2ku��d8h6�	<��`X��
0[�Z�Mت��0h���YGwS�(�cu'��*[w���Ӭ��CJ��Z2�̑�����X��m0ުPikP�>����J��!zh����j�!T-�a����J��e�,�V���
�s(V&s �RX�Ye�4@?�@�뱬�Yz��KV��
	�gj���R�1�9�f�X�����Vo`�6E�ň���p$i0ڤ��Ė�������
�n��E�n�hZq������7%`X�2���R��X���iMt�">3������/��O��,�n�x���N����M�vk��=(JŒ�5z��h�M:���<��Ò���r�F4
��I��Л��o4ef���1�(l��z�mh���o�-�jC�#�	��LF3����$�œ1�`�ׅd�pk��p
g��I'�ԇ��,L-�9��(��:��H����";��ڶ4�3Y���fl��&Űv^=��`�v��+ښ}f���*zd��A��L� ��*'gAw�m[��RF�Q�[6k�O(�w�F��Gz���8�E��C(8�T�b�ӌD�J6��7@1b�.��
n#�}anÅ����0*�f���Z����	7x�U��m�^�)��Z��w2�,�j�Tz߁�p�J۬D'"&�e�v�7�`7k��v�^�F��%�Z�wF��т�I��
m�Ў'W���܊����Z�RʬBѨ���v5���*��M6N�9�ɇ.�i��ʋ��KD{�O�5�r@-L��7J�] ��6�j�\���SdH�u){��	\� ^�t��V%�F�k��*^��z,ݕ�)]5���H؍����1j��y�h]�m	Z1����Pn�4�SѻB��4\w-�Q�;OtBbV�S�:���t�0�T5�B+�!-_`$��MA� �B6�� �	�&ˣnT�:u�,�;A����{�����eY���SR��Xڹ�0^�4�AP��h-��&��?$�����u��Kg&�=d����_kAL�w����1�wEb��:����I�DY�ҷ�d��9��}Dx<<s�������V��O
�/�m�ؖF�ٛ��ˡ�
|󂿗���xnt�n��X=c����[�Ŋv�R0C!��ه�B3��L>��b7=[Nōi\6���ppsR;Zx.��k)	}���[��b�z�{��g��\��ً��u�|3���.{#=�X@?zdZ�t|��;@.ī������Qޑat�{Y��s+#�.uL�"�.guq)A�؊���m�.M)t,��5m��8P��j�Ҡ�0�a5<�/z/$�ϼ�l�"��������Apw9@G ��0-�d�T��NZy��G����M("-�#���麻b��~$�������ڋ������h�ܦ�Ⱦ亳q�|�)nbC���j�2�Į�����j
�<y:�hj�c\��2�r|9�(%2@�VB�aM����жf1���+��K��S�0�W�{$gۖ���m}�r�������P��ޤ���)�]�y�n呃�]5��%����7~c��jTf����T�<�����D�=ןh���V����U���_ךp+;[5�B�M�spu��L�W
�	���x��Gm���zel�s�l�u�5��V-�Tj��5 p����7�-Qq6V�mA�hWNW�Ag_
"��ӳ��g��gdeg\�i|!��#U�|#���oǱ���}T�x�8sL9��.��HulUС�D�e���hI�8j���jn�<�W�nҺ,[��J-��}��u�&�S��E��VY�R�Z�Z�����op�tL�D�z=i��`��r�Ä�}�֌��k���e���(N��R3oo��	/����.�s���x�<6X(��1:�1�挘�����g�J��f�Kt
7�O͇Jd����p���$0�1�M�)�>L���[�v]�k�y|/�0���89���}VG)�F[l��t/�岹����7ˉ�/��P����Q^�CJ$! ��6����)�V���;Eh[�e��c,���hU�\�����u��N�����89���bu����8�������8�僶��7�1��0���N֢��.�`604�
UL(.<B��{݄��8�.s$�vRg�!����wUm��'�e�l#�3�%1��B}\�ڤo-q4ttor��[�sgTV�B��c �e�lR (����e���6�:��x��g�`�Jv��qN��e�nVr��uXQ96�4m���ʩ@�N`�dn�x��{|�r�Q4�+{�ʶ�U���!Yb��T��>�����"}��<X��@й�$�R�,C��������f5�}�yڛB��(:�]��v�k����	r=pn��h˗rA��U�9����R���NgR��tWs��˻{5��m�O���S���z!]�9g�їIh�kQ�y�v�8�9G^3eX�@ӧ�.��Tf��4�wLjT��ٺ�VK��zH�/e�}�ڝ��ov��82p�'�]
x7q��l���}�
ǃKe�Nd(�&����e.8��}��V����a��������:'m�$��aH;�Fs�U�M��CV6<�Y~Y/���`�p�Ŵ����B�[�% �]�^�:�n�XW_a�2P�0�s@L�D��	��:O�ӖG�Uh�pVg`E�(�B%�=��ul�<l��2��`�7I,sp��2�t���jE�}8���W�Եi���j��hP�jevi2+MA(ZtXt�8�H���&Z����!�z�,�G�s����݃�J'�ZU�w�a(@*|�P�e�&�&��v���0�V���3�p�[�U	ۡ�I������V��:����k�/r���C�f�A��ciE��;#� =�u�E�x��t<~��{L .8��O�v����T�a%gi�+o��t�
f�*��=������[4vK1�`��&�ljNA6hc�0�·qq�	Yل+U��2G�̧>-�ׅ!5;7\7��q-�.*���j0�Ӊ}u6�+�o����	l�x|-�#�a�m	Ϯ�Ab�)���ѫ�f�5,��0�08�ʸ�Rp5*�Ϋ�*Wt�o��E-����h������?B��a�@xOy��6��^�ْ��}�b�e���
�ͱ��̭��Id���&,&�C�R�5��ns�.��� o�E vz�����'/f�I�}X0��*;�s�.H�v/$�GF*��x����k��:�\��{jh�mvC��܈˧ٹ�����­�b�p
*5�C�A_^1ȽNƖ��U�l2�e�3"��ؑ6E����}���i[|7Ϙ}��vj�G12�g5���o�ͽ���ƟY��W2��tD[r���s�΅Ħ\�I��+����☼�dY(�۴���!��ca*+&r�P
<vy�����nq]��f� �]�s@J��{s�G����ô+aB���w�ȉtm�5���<b��5��y{Հ��b��B�k�[�pΛ���0���3d�&!��:�:��d�b�=���8�n�ιl�7Aq�je�N�� �Lº�S��u����P�c:<3�Ҕ���l4+�rmlMMg �x� �5@o��y�1e��j�/{l'`)�IQ�{��Ȅ��K��!�&���\�Y;���Z@�U53u�H"�\!�׆2	���&�|���Ma
!�e�R2 m5�4&Pݮ�*%#\'Y��Fh��VjV ���]G�)d�$VsVB�R���|7a��Y>��p����z�l��={ƹ�.��Ȓs�\�����Rdj�+��ە����ߜ�-A�J�����C
��X�3��3֪�&��I��ݺUFu]6�jL�(j8�Y�e���2POq��k6>��<�<��YerT���F݆:i�p��{�{F�h�-��L�V� c�׆	����]����{���ҩ*ɩ��)�e��Nϛ�\�i9�O�sh"�tiϷ�Z[1�kC<u�ĺ��Č]x�*#;�\�A�uip��XN��6�,�f�.��Ii
��e(Nv����i���f��ES�V�1c��������e�|������Cvu�t�-�ZNB���1g�9��V��e�l&��l�7ӥ��v��~���P�=;��U6��3f��P�,D�QvP8;EQ�C�[�3�(��5�����S�K�	�e`}\��<� ��mLV��T5~��'U�����9������*��7~.]<��mw�mw�[���&�P>�� z�=pN{I���g/hR�څa$�bK"Qݥ��|��KNwO�#%�
�����O����ä�T�`�8�6�����<4̽~�wk�y/�8��I�3��Efeg)M�9L�D�#Aq�����r�߰CF��QQh3�Wv&hcb�wH����d拁��=�غ��ǡ����g�� �f�.o8�hg|v�Ay]���{%&�3�'��y
V$�`��Ү��ΓݠҾ��_8Z���8lpxť��2.�)pg�e���:�.�9Gv��x����n�ty��K�&e.��V�z��B)p���nZ��,�TF�u'��Wo!�f�ڰn��7��S�=@V�3��i�
�<"�>?E��}bŇδľj̮P��:�o�K�OZ��e�|�}] �\��_��<SM�Gt��;��a����:e��S�c��u�)��s-��QWi�k5�S��omZ�
�w�D���W�=~ ���F���*j��������o;�H��Pޱ��%xE���yZ��|m;���7N�U��uMuIj�c�ɲ8M��V͐�r�$4lٻ�t�[v�NU�]�NX_u����9c-��9{wӵb)�iJ6��G��'+���#6��9Ñ��f��=�����=k�Pǎ��y�]D��2�сK���/�lDf��	w��s^B�fl��ꥍW=�x`y��V�7��0M�u�T�b�,ua/z����XU������f�˶b�"6x�*�Mb��9�[�F�����=L�Ԧ1"W�Xf��+��g	pY�5�bqmɫ�e���������vM�O'Lx~��4n�V��3/m)��n�Èi�o��$�J�Nj���o] ��¾�n��˴�Ρ�h�_ip;듯����Au�=2�6���>}�צ!연��у�Gg�_�i�RN�o�uvf*���PF[+h#v���m�x`�������N��k���p��2��0m!��Ӿ�[�]����<�<�il�Γ�O��v��Aj��&$���2����U�Xm_R|4��f���H0Wbg�ޯ��/|�w�-�+0a�qf�޴#��v�/�-�VP��kn癸�w˪Pv��"�R`�3�-�������ʾ��z��U<2�箝�vao'-�u=��{�K؎<��*l�LK֎} �̛Zk�C�}��k'jg�cM_wQN��X,�]�iyԛv�$�'��8ΰQ�iU���-�s��	W.��K��i.�Db�"fu�"�u+;ڂu{|��tm�2��x�(��}Uz/Sx�=�x�l=/F$��2͛��v�/��㝳�e5/������o&�Nx�l뼮O�ǲ��J乺�I�d������o�{h���T��.vRx�o�5J%��<�.��8����z;��={7$ͬg'���x=�q��\՘��ҽI��5����PH+�������D��*;�.��TQ9�� [�Uz���%����,��X<��N㣵z.��)��Y�Sk�9Րh/P�Ҿ·�4�n�H�a�Gt���<s�U�q�c�{.+�\�o��S���E���=�i�.��Ծ���|����0
��6��|���}��=PI����&�ia�%�z3V�,» K��`�������

�A5w%a�J�s5��[o�`�3}g1N�+I��%��G3i�R�}�U#�N��UǇ�w]�K�	�{TK�݂��Nq;T�T;�M4����𨃡��M7���K�Pl�B�N�A����j��]�E��ep��7�hkX���$�"��2k�xc�	�$�L�m�K7٭"��޻�,��wת��FZ;2�
uf�G��[���x���M�����n�Zh��Ke;|! ��C��AJ�q�w+C[�<Z�!2��Vj�	d�d]�_Wה7Mj���:�k�ޚ�� ꮤ���]��}���u3�Gz�(��}X�dQ(C��f��s��� �[�"vnV�86_���kkC ֊�;�xk�v{WYkh�2��-�����xpnR�s[�Ǜ�X��u�W��)�{c6�m��ZU�h55����`�ò�+f>���I�GQ��6�/�����t:�(r�>�-�"k2�f^B�fI|YO�o+k4�X�w#��3T�շ8-4��4��W��z4��B�i�]��K��ʝ�i��;7��lY�w#l��}����w�2w�z��]b�
;�WB#L���a,�yF���[�79�c��@q
t�ݤf
��S��!]79��7	v(���f\AU��@J��u�ú�s;��{[�(x��l^�/4}���B-�^�N���w������Ӫ]��[ej�T�44��FS��侘{�L>�����7�-)�&_F{�S�w,�MDr˖��[^�z��'��f����J#�m��{j5��Y�"̽&��ܓ>˲�t��d�~d˽�Y�h�Z���:�ap�s�z�O!\�Wa�=@@k�u��dg�����$��b��j�����C�Ի��\J͛��T��̲�������9�߆��.�=�[@�h�N�ˠD1{���j�obi*`� .��i/&�]~,<1�!�Y
�5���L�coF�pd��e�& �q��S�G-���_�� �فY�"R�����J���n޹3\\V�+����������@A�U=����G��ٝu�u��	����L��'��K�r���jUÙ%�'J� �1}���H�v�2{��:o�L&�ѽ��m4#\�� `p��Z�c+n�qݨ 6��N%Wv �_*�X`ag9Z��9�+.��Ҋ��Mwǩ�Ya+ؓb�I8oEZ���1Sz�R"�R3,'m6��:��9x�׬$Fܼ
�����j��zj]�\��̰�r�����u^f2d��
ҥ\�m��hHn��ka��l*{nٳ<��Q������;p������^6,_���O_��'fK�Q}(�oJp� �QAu�}=��U��,��bU�t�_�y2L3H����X(�ֱ쯀��+X��xn1����̪���@�F�sF++:���MAtZ�w|�ZB�Y��o����h$�9Us���4C�!7�N�6�Eo`��t�����AUn��n��O�2x��Z�R�0�.�ј�.�J���$�Ж��0�Z��/�^Wru�}U��7��� |ω-�)�g}���t��.(�ɜ������zz�<��=q\$\�v����&A\z�d���D��[b��*�*Mcn�T�dK�.WG�'���-\�%9tڇ�|ܬ��u+l�*oo��Ij�o'W\�I�<r������0Z�����S���]�k�M��a�������b0��CݴL����-�AI�{`ܴ�޹n�r���Hy����{{�^uިk���d��oɼ��-j}�P����X�d�
v延�y�6s�dʂ��&7Xf窞'q@��x7'Z|��Օ�Hv�*gBouû�ߎ�ص9�^޶�� =�x ��������;dS��}S
4�݋������.�}}t 0�s+Q�B���m\�Zݥ{����3�)7r�oDJ��+
�>˜�a��պrl�mrق��D��p�`�Z8���7�&�ڟQ�&p7�g�Y�a�lKZ�Jͼ�*�F���!�b�-X��_��"��{<Iŭ��^�i��fo�����^ǫ��Z��,Y��xs[7�O��iA�--�++��E�1�:n��#f�����w�E������Z)d���K L�#[Y�B�&�o�"�-���x���̋���Ӡt�(��Y�hvn��Md5��<i��WL@���Q枝�2�h���T�5W�c����D&j�s����X��K��2�2�6��Z�*�����Y���uje;�Y��y����`����,�Ys���c���),!g3�G�h
H�z]�����T��Je�'�Aa{*��5;�o��h�-�^&��Ԯ���S�o�eĨPe��0x���d-Fѳ���ԋ�
e�.��k�wL�
����bYprK]IS���h�@Y��y�+����ӉǵnL
�ָO������X@��o�oM,�u].q��-�&^�`Ze^¡nf�n|N����2�S�VL�����]�d�z:|i�EYRao�P*����̶�eR�re��&n�T2ms��=H]�����9c��
�2�O�Y���P��)o���s*���^({r�=.x� ,N�3���w9Ǎ�C�Ӡ�k8�H��o6^�ɖ�c�wwx`p�v�'�bEu����Z��V�؃-r����U��t��_�,�v'��[W�#P�*�Q\�="&ޝ9��`�l7�D��B�m��^%�9²��kܮP�A8?t�m3���wf�8�7ٮm`��(�e���L鞽o,^(ܺS�^A��%��3�)⤣�����6��w
/ħ�ô�\��Q���s�����>i�\C��!'bmA�l1YKGtĦ�Q>��Sgd�G�\Xk��S>�+�[�{.�9�ㄬ�#7&�X}�R9����@���pi�rT�!i�����ރ����i�܉��P@�4D ��#��i��;ӡѴ{]�l���woOS��soG#6��ݱ0KH0%�-�j�]< ���}��4�pZ"K��
Ϧ�!rj�dsH/�S�
�k9Xz.G[*S��.��f�x��j�cC����T���Sx]ic9T�j�uT�_٠�e�T�Qj$$D�}gv�]�#*��L�3h���H���&��,��}���[w�/v)����N���dx*k̲�D�fH��iL��@�#2j���ОT�|�,���B�Uf��]�̐q��䝜�%�ܞn6 A	�^��[}�2��u��7���6TJ
ҵ[`V�<6�bKk��nK�2Ь�e��,�ȠN���F))�4]c�c����K��|^@�t]ଫT���_]J��#�Z�\�J��Y�nC�����[K�NÃ(�r�q���F�W>�LT4 ��6���t�����6�s��;�,&)3��<ʰ�
����{ ������6�K�TFv�?L�H5q���z8or�t�#:�p�-�sg>�ur'�iR�Ԣ�;ޚ�0�����֎�9ch1�n넮7-�Ul]���%�\���<ңw�x�ш��}Yɷ����J����"
�Nm7��c(�R�t�R���[�\����z���hy�FU�fH�6I�Ѱ*�^��J�Y����2^��fȄ+��������Nb�rz+s^��BucK�a)��s�\.���S_
tYS�+-:��^Pks��ĭb.�M1`��SF�0;r(��J[\�ÃS���u!�ʴ�ivgv���E's��Ζ:�w�m�[�1�F,,����5�����Ce>^'Vz�򢂖qӖ�c:��}�c9�!1�n1j�CKZ��[q*hT{	��ľ���[�d~�Ѻ=�ٛB�bY�	��C�����^�u��j���%��G#�y�im�n#�0�Tƀ�}������R�P�ݨΐ�r��Q8sx�.�@ɉ��3f������p�)[�B�LS�)#�,�f��1�)���`zUgt�eY�K(�@�c٧f��/E�E��_�y!i�t���[�.T��݈{��֎��������+���]�@��i���"�ઙ.���n��T�uB�F�)\�bH����ӵ��x.�c��VY�pLV-����Bk�NqXj����N�M]�1;�0�9ݖ�� ۮ�� �.f�2m^�G��(,��%7���|��:�X��k���ɯv�nk��rZ��p�������݀%��2�''����. �.�^U���� �x.�����@xp.�eQ�AC�����dt��6�a�:ʘ�D�KN�S�K�e\�DV�ʴ��
#��)>��w;U@����XC�L!~j��^��^ť�Ѯ�P:��!�̺K-"x�&%jر{D�;��np�匬�bu�v0.:�����h��&�,l�uӲ�&8TR��,Q͚�����u���Ɖ}]��#H`�o���VoS��CwfV���pY�drKղy�E�;����!�7kӁ�7���,^���h'� �ǹGEa ��dt\d����{�3�wGN�]a(��]�쫔ƊkQT��Y*�|�S��Д�����5���sD#������u��b���u87�:���P�1�Yv��[�K�JN�Ւ�;I�qwX�*���厠�����9z��u����$�;I�ɑ�ֆ�.��&���B�0/.������T�'΋��q��\���+��݌JIŜ�6����:��q3�۵
��R�Ć��N��i���=o��xrHW��&�i�8^p�^�n��j��[/5J�M��s�}r�4Zum��e����I�d��Ǣ.JB��X��z�3兌�y%�U"G��>HdZpz���㌍��{�cr�Ko�el�^7��8'�����軺�Wq[5&0h�W�����,m�`Av�;�A�7�A�!v�E�`q���h��'gv�h��;T-e�<}���L�\.�	!�B9�9���ˉZ*"�| ��w�.Yvɀ�M��
F`ҷ.��8����U��YH�}�a4�JM1x-P3/�b8�we���n�|E�R��n���g��y�@e�6%v(��V�:sQ�����3�h�GIą��e㕦=�*B��]&��i�._tҜ
��sme`�i�)^������-|$��8�'9{&�AѢ{��Ao).5o(�/;^�if���` �V�:�{����UK�{Â�ѫ��X89�&�X����%�^%�������H�*.�dxvH4������[���϶}�\B��թV*7�������t2ʦ:r�{B�8��=�k{'."�y� �&:�Y�;��̢m]@je�+o���U��2�t�=�}�>��Q��
WޒS�fW¿��*��J.ق�l_;���66B���l	H��+�!eq�FmNW����H��.%�7��7���@�����������8�[UPY��(."T�a8,Q��j�C�2u�Xd���@� b�w �_2���1�C��M��2�����R��Tͥ���/E��gm�t�m���>a;�ytZ��vC��<eA�ׇ*��Wү
-�\3Z
(��W��Ŕ�]I���Rˣ��:K������N
^5���f�}V��������B¨� Y���sY���_Z�i�ǔξ��&V�N*�Yڃ����c�o]
v�hؒ$f�a˧P*v���m�� �0�����f�v�N�YI����ч��3� �kN�/�bCX=8���n�����z2�B�5�	��b�Ҿ��a+���c��-�e�y���S-����f�����#�9�����W�`���{wɱ��(�8���u�K��-)��
�iB�U|��Mb�nIU�w�k�>��S���^s���6�¨w��ﯳd�J)_�-ݴ*�y�g�� ���lƴx���Kx�ѺJ<��GVT�׻�q-��m����>ù�ݧ_���os�Z��֦	��`2�9�a���tx���n���&��#Cs��pp�]�}���� d�oy*/�z����˛�'g�;�hy���$�N)�ܶ��'�@6�E.�&]�ڈXh�� =m[��ݾǷ٦�Aa���Z{W�Ť"�j]h���܎Z�-�Sgf�2 �u��LB}<o�Y�F彘�h�JU� 3��[�3;V�|�{��Q�O��Nu��F��t�������W��}G4y�Õ��c����o,M��P?N�F]��VS����Ns���Y�CD��>T,8�z�_6�c��g���S����7��d��7E=#m4��$' �.nvU�J�v��`ނ����*��:�om��Zߜ�.��LƄq�m�����]�7D�M=V9Ф��
�g7��Ź��.W �E��@�[{ڞs<2^���pGR����Z�ty�-v��K����Xy�/���R���M|�q%D�ΐ�@�T �ۛf����{X����}���[�B���0����N��:�f2
�Yj��I<H����}�N�g9���$�ф�ܘ�"����xv�.����b�����{��oZU�`�Ό�i�\t�.�N��n�N�@f���lG{��,��	�C^�7$�W�>)E���y\�����������۷�X}[��}����׌ف�+V��^��{)�� ��}���^�01��/�(:T��[׊
,\4�V��wK@���"�{$�x��=x����,C��KZ}��*Ӡ�d�]�.;ƍ�V�#���,���*}����ٛ��V ��_��9�B�F��Q��<E��`��/&mw8ǁY|x0�rw<GiJ����G�<�P��gur�j�7���򛔉��{]���Gl�
�7Z}�A��:�Eۄ*9PԦ����g��+9]+�V�w
+y�h�q��Pc�t2P=���M2Crp���r�Y�Z4�S��	�/��:�LJ�_f�ͫ�f衰f� ���٣D6&'x*�{���k��/O(�]�b�tA�/��X�4��B�T�6 ��ܚ�Zx�/�N;j���z�6R�7 �@F`��㍞�uS���6F��|��~��=���U��~C=���W�<뾗���;�#/���f��P�5|˼}�:�[�:�ɻ�U*yƱgXCg���*f��c� ��*I�����V�Յ2�=���%�s�q{�`�l�m�mK��E\+oT	t��l�)�W
�]��S+�
FK�P���,A�{����d�����m�B��V�oHI-I�4Ll�<0M��x�Y`Q�nY�BŅ�]Z�D�9�A1vu�P�=c���P�Lt��.��Kf�����Qᄎ���8}���n��(6N@��P�*��|����/W�*�|�<�C��n�w��n�9J8\�Y����}��F��bd;����|��BiY���a޻�hT6f-� i���)Y;�;�-��;��"b���؉�"�+�#Վ���G���fM'�q=�$8V6�7C��ٲ�kEةc���vT��w-Q�T+oxw&�|��3x5H��Xi,�V�«D��I��msw7Es����m�`�l��z8��vqj�i�F3��J�\��]�V)��j��*�oIp�]���އ�ͱ�.������:����<2Z�~��qX���?-4vv`
�دL[t�|`�m8m9� ��w����{��س�j�=�9��]�E>̐*m��2͍+QyȎ˻��㤩N��Y��2��E���������4�Y!��jt[��Ie١'-г��
gp�NA��ں��0RB���6*�&�Ά�������e��-<G�-�8Ǵ�H5��6? �n�.�[�Ă��U�dT���u���b��j&�`�t�P�C9]�t���͸/��G��rQVgF�8Gi*�r��t����f����ʗ���	]�=̤�����{�5稒Xa�u��v�����a�:���tw%=��-,El];�����I�WZ��(:���YZ�u:�}g�*��6�d����n{[��W�{�j;Z>�gB�qd��0e����Yb��L=Y�/s�^�ewZm�+w���-r�P����Ե��XA��r�걇��������DR<�k���{!'m�]��k8���:�$n֬��V~�Oq��*�y}׸�r�����ٓ>l��g�2�+��dz齼�C��Wp_���p[Hٵ�[Lu�y��zq6�m�<dSbZ�ق�b
�3Q�.�U�W_^��=ϩu7�g�c�J/��ѣR�mT�b�9�$�3��A(���0���cNP1��!Ʉ7\��ñr��W۽ľ�W��m�B�.4��ØS�t�i�w�9��Yq'�k�)bX�1�;|��= %��kK4���z�b�Ը�UU�©n��ĝ��m���Ec����7��Ӫ�7tN�r�s��U��.������ig\6�ǶLY4^U!��ؾ��]�%3] �Z's�B78�(U���@���J��$(����VV��bl�n���r�-n�W{���c���:�9`v*M�[R�*62�W]Y��Q���KS��-�]�q5q<��M�W؋�yC��v$S�l�hn.�i���a�f�����Ȋ�аv	��z;��T �F	���ټ�Q�^��	�Nθ!��E��$���y����#�t{Bh�����Sy����
s7���pD�G�;���vJ�D�]��10������-\M]�x~ZN+���xx{����{Ι(�>�1)�pOR����� 7e�r�V!ZK�o����\���j��en����'1*��+�8�J�	��5�f���Z*���(t��\���8N�+�.�5�$7�M" �
K��p�w�h�����u�K�e���wOTge:� f����"_sS4K��Ր �\���p�;��t�t�3�@f�oW.���e� 1��-V�ɹF_��ޔ`�<; �:��nA�RFTw��YD?{��۽r�����'d��9�F�r��Z;7�g�T�Q��E��18ܫۃw1���|��I!|�bg�N���4MT2r?nt@��u
t�^�/�*밇�Z�{:Igd�]t�V��Y�m"f��ʑ�{َm�²P���;BYw �����vwU�{7�2&;0����XӸ�}�]t�Ȏ��� 6�=6���(��|j*z���,�&�@rW��4�Z�60vU�o^�<��C�:L�6�bR�&�����u�n+cOҲ�hv焚�ժt�ݐ�^6춎��n|�p����1,���\y�J�͉Bt6k�ьە��4v���bՂ�C��gc�B�����˞-�u�f�O#��ƽ�������z��CT��.����nkF`t�.��zXB�
-�ɋMʺ=�(�*�o�mjGZ��Cԍи��&���r�]!:�d:�� �C��/}�T���T<��pYPO#��y��NUET��*���̩�\��^
�UAY�QO-.A�AVdvr��+�p���쏔9��I$� E�aռ�r5�w(���^"Q(�V�ݵ�(�����U��ɋx�t(�"L��TshY!��%y�2]J�"��".I��)$x��#/�ЎTr�����p�EZ���S��t�'k�t��!"*5�iQ[�ꨕGq
y����&�6WU�
+��N��̰ČJ�$�elΚ%4C�yŕU^aE�\�ʳHrt:H�QUPQ�*�QS�r3"�H�su�\�R��w]��J��^I,���fʒL��"Ҥ���'Q�rCwvr#���V�T������������̾\��'GՏ��(M'w��F��i�9}���D�v����L�8���t��ݦ��wJ����>��^�.0@a�l�k�����J�:��C8�k���y�W/��Tju<�p_�m�\)��Ïإ�G�#-g�<]*��,ũ!���ն��4����Y������k���,�N�e����S1�<�����Z�\k��.����싰�fv�j{&�͠��bpվ�0��"H�f�{�B���n,��b=c9	/�GK�K���}�ǈVK�]3B͟V�Nr���^ue�9wJ�ts$8��֝Χl9�s'{AA#�i�5j��qFE�&9���`ߡȾU��ذ7�pչ���Zʹ����S	)����ȡ�!9~�O���`�pOm�$��Ƿ\�(�	s܃�~&�_9�kn�{�F������;"n多�Tԅ>�C�O�`�N8� �n������-{�,�݈
���Ѻ�{,�ӣ�WT2�u��7�	�:D�����&<�q7Y��]k޼]K.�c��jዂ�y�2���A������5�x[��W��'�8<���UM�����V:)eطў�z7y$�<���U��3�f�s�+�Qj�I�j����W���;�d^z/���5�Y�o1l=)�u�D�R�@`I�u��V�����<�'��b�b}(�D��p�9���gN��B�%�w�򽹕��>����y����'^����G�j,� �u�`p�e����2]	�[}��	�$�X�YO��WEh9{^��������2������/���>6�y^J[������w�逻$���T���Ԃt�vΝ�N�E�Jӭ�J��ݙ�{ܠ���E\�HB�)�~j�GTyvL���&��q�(;�9%�ȭ��=�S��j2��k�ݢ��)åhY1��)8���PC�O��/'�Mnz��ǫ�ԕ��	�H%�Ӯ��fd�[O����I޳ӄ����懑�c>?`B�\��ǍbJ_-����s�z!�3ã�HɩY�UU��%=����s�9�"p� �{�H��ʥ<�QN;3��^7T|�Z�[C13r.f�5���~��J3]���'s��"���^�����^/u��#�&��v��L�3eU�\��FLF�U���9���H�`�ZY���Ηx�?/��Jv�$]�A����j��Z�$�vO�!��GM�"��L���a�'|c�tL�8�o	���Sފ,��O	�+�J"݊��,�V:8|{�NO-F��wEjWj�i���g��y�-��W��n���zY�ׯ�SYJ��:������Ƭ���]]e�9��fW�/L���7�<4�����wLP�J�'h�z���o����5�Ni�u�bes׺��^�j�`��X���0r�.��޷$��59Ȯ�#�=(U�t4��9M�y)�C��r�%��Kک��g�J]�����f��<1;>��c�W(2�K��z��GZ�}���|{E�?7{Żh��tr��Ǣ���w/}
��Ω��q�@�·m���!����X-�r�nI�t~:%4�����בucQ��\���ч�Y�c�مR�F	�
{��_0r�gxj�Z�Z�ސ�h1��I�.��zbjf���N�Ž����w�⑩SI���&/��>���Ėb|;�WE�I,�>҂w4]������n�cCǥ�s/ӛ�k,��τ&r��M�p�&a&du+�H��zZ�8��l�t��=է�v����އȲcD0��2V|�x
���rꠊ���{F$�um�9��G�����8�`��v���R/!!n)�'u�.V: �.E���&y��&���*+,�aD��l@
��t�O�Q�˥�����n�2й���H苛��mw��V>�${Jmz���^�LkQ��5�p�a���!M�伖��^Q%���s� �¢T+ݲ�7[�H�x�7�Ra���\� �F����1n[r�*���#� Q���A��_O�������wGz��Y(=�+TE��瑊�͒6��Wu��;�-��T�]��<+�+�|,0�����7G�=�ኚ[G=����/���X����:��?���[+�XZe�\�z�h�t�\�k^�¼��l�������j��DN�!��T��w^��"���z8�2rp+�ʯ���Z�-�~���m��w< p=#Q��7ʻ�xVߵ��jCV'�Ç�(b�����)�!����V�G�]�Jc��د����BΜh��+������V�E�m)�9��+Vu�U,�m�:d��$.G�ณێA8�7��C�}���j��w����quEDuk����Z�+���Ҋ��SK�W+��!�o�ub���16�H=r���-g��/u�;竽s��J��>t���\��7M/�q.볜!<����ͷ:b��5]��ڔ7��(�Tf�;q�^���e�N��B�`��x��Ti��?n�{m��I���V��&��x��lf�4Qj����'�42���]��[�EL��ãi���.��>�b��)��C������\��Ԗo4xzU��U�M'��c8;�16�MP*��{�*�3�,�3��\#J8�IWn��wx�';q>���na��!�m��uh�f|�� �i���b�	$8{gF��>&k7y���E^D�Ş��m^Gb���
��U�Mz�j��H��z-�yӏ}�����(?��&�6�8>[��hߔ�e�c%�_C���_85)�'��Qe`�=�}ʌ�<�Q�B+����:s��7Ӥ�fX�	F+{���7�6�}�����Z��L��e����Lׅ�V�/��������^*�J�8Q�ƺ�ncxu���.$�.���G%4�|=�Pz<y�S=��ϰՏ^�����o9�����rl��wj�X��OB�k�#D�Jw�ZCL��S������b۞KUf�b�Ǜ�Qq6}Z{���uWa��R��\�!��ub	]��#���^;ɼw�����w�;�GE�t.8���z͟n�_'���	ν�_Y��Y���`�Q��z��g(�N>���J�V����&b�xS� g�*�����o�^��z@3܍R�\9��:�v\fT5����u-��U{��dq�r�w=���k�hg���Y���SS�᭳�U������ޥ����#��Lg���n	�vZv��L[�w<���Q�d�h��:��Q���o,�,�v�����Ӵ���.��JN�z�ԧC�6 �{%y?�?��\ͅ��@{g�� �|���(��L�M�q�{��ݝ�g
�c�jک�~߼����o 8�
6} B�H`�V���n-+��#:b�����tY<�T��#Z!��K�h���Q�^��'�Z��SHh��cÞ&��є�ow��L��F�N�4ޘ�ү����q�'˯;
��b�	v3�3 ��䟁�{�l�\
��& 6�J��r�5�y���p�;Z}Y��8��b�\��/sA�,�ț�#{u� ��C&<P�Lyd6��+Z+��.ϴ5|��tf%��Bt��~�q�^���d���s�Fz`is���>�0�X��t�Y���_v=��H���z�~���m3�ݷ�,iiv��&�iؚ AfG8��$iĄ���㰾�R®b�ߥ�k]dS�e!iw��Һ�)��E�g�~�7��AQ>���]��<Ӫ�2��wz����K��,Ƿ�9��2o�������jh9'jK?X@���l³�����5q^`��8*�VG��ܰ|__fW3[Tyŵ��V���.�o�DV�哮	�&��<k9�],p����צ+����8� CF��-릉cS,��-�a
b�r���Ƞ����9+���J͟^��R��hU�g�_�c�����>����ެ�U�Y�m=;^.x�it{����Vs�7��*�2v�F�j͌�wOG��n���m��CmY�./���e��gv;(h��J2+�qY]�'�f��4_-�q�����_�G����T��U���ڧś*��93fgb�jM��m����i��OV�.z�WK��O����K3GD�h�G��F�;�t� /���^��ܽ˯d;�Gn�6�E �1O)�׵���#Sya82��a�QZ�S��U�:�ۤ�^�zkG[��瘁�TI]�w��x�4<zP���ix��i��%4(8�*��SY��?Ezck
�t�r�gR'OZvE��+��}/���hB��tAe��Q\M;�B��|���}3��h~�*q`�mv�P��*��i���ygs��\^�]_B�R]IȽ�'6��#RN�i ަa �z"4kȺ���+�0[BZ1o�Y�����'�y1천�R����^_@�x+��J��h�>]�4�Vڭz�VrTT�>�ʞ���-,K���H�>��\H9������ŋ�әU+eO[�W�%��5s��{e/>A+쾱���y�����s0�]Y������r|x��
�$���TH4Oeu漒_�G��m�h<��;���6�N7R���a�J��j�t!�)wpzJ�s�q��M��wD.��n	%��W�w ��|��
��59���*���ڻ�虯p���+#�`td�T����4DJffyԮqa"B/��R���N]6�t���b��)�#׆R[mLh���Jϙ�P�c4.]Tۘ���>~DՉCMHY{=����0Y�'Z�]�}y�qL!#u�.V: �.E��eɡw�"����k�|��+`(R��V%//Yb�K�?�ٻ"�G�����Y���c�7�1B���N{u��d>��R��<�G�]��
�O���g����s]�{���}���}!���G��a�X���}��i-�*��c����
b�X�K�~��O��h�k])�ƒ��@�����9�'��x6�.��D4��W�Վ����?����k>��M<z�"ҵd���bq�lB�|���<F��<D�ls�X��I�J�L���V5�����j_{�W�ԗ3�|��=��}:q�lF�|��7��-�,�Wʜd���z]�H@�h�/o^��vH�V��Z�7`�V�ǝ�\�^3]Om=�iK����^��yNLz�~���R��T��J�H�}�3�o}���Ga���/&Zk�zg�\��3$�Z; *--�Z1�2:�Y�AE��O���m=;r�@{z�Q�MND�>����}��/��k��|��{��19�M��Hu�ڕ��v�f!��0�� ��/N�
6Y���R� +��i*��nquറ\���tTn��^o[�;^z�:�K��&��I�
<5�8)�s�Z��dq�r^�`�YjNTt��w9���d&�מJ/�,��e{�آ�t$�p��@�>�ŵLӓU�s}������3ogc,D=�8�������
�0]M>�"�z9Ǯ��X�S�=) 5�lܿzeH�}lI�eN�a]W�I����M8���.�Bʼ��`w@�$Wt���U�MC�Mh>�ܼ�uV�P�w�HD����Wj�Α�+�3�����V�6�.V
7�H�^TI.��w0D�j�k�~\���#�� 4"p��B'���y(�>՜�-��\%3/6�N���ζ��q� ��}�KT��%�o婓�7�k@�X�U3^���W�U�	�/F6�=��~�oo��>�,�������.$�yp�s��O�ǏjX�vs�{�/����
�=._�ˮ���l��:V�q�v�i�&!Ŷg.��x��v��6�K�`�{����ō��}1O���j�$�O-9�0�A��m���{�h��zvK}k�l՛Q���qsobՙ[G��\��*i��3�7�tPl��G.oa��.�jN7B���-�O�s�&�z�:��h���a1���0�5��h�Q����)<o��&�ZX��zc1,T16�&�ۨu����9��t�y�wH�F�a$(�s� ��Kܗq��-x���YWb�m�V������M��g9�>�ޜ�y�<��:f�gu���Ƨr�}����Ֆ�7|�h�����������g�S�{zPؕQ��I0/"�j&��f_���������#�ݜ5�����i<��>�!-!�Vr�˿CO}wt�]�AGX�76ͪ���]��9<�w��g,s��Ǖ]CI4�SR�g��C�Ij��Wry<˱w}Y�َK��$���>nF�({,�yZh{��+êI:��E����3��˗���ǜ�Q���t(�^w�ֺ�]��z��p�F�{�`<e_s ��iP��VVjm؏޽��	��ʐ
��T�j��x��}+K�p댝e'P�<{�.ۻ�-�S��s��0A:�(d�,�+#yEx�	�(�A��������;�z5���)-̕v���o��򂗳�χS�X�R�XU@��$�Yʢ������gQ<�R:ޮ�ٽ<ŧ�i���ۍ���Ƭ��aQo��G8��(���=�No�R��]x�ݵw��ϙ����k8*�9�3��qz[��,�(OS*��#���<2b�;\r{��ë+���&��ˢw�e�����\൤AN\�AB��7M]�jn����AdL�AM<�戜{�`v:z�P�t|�ʲU�$&+�Zf�%���O��r��*:Y�^p>�]mfߝJ��G��yv4r�5�C���Q����Hµg�h��\�+�LV֜hֶ+f)�E��h��Wܬ�M���rDr��,ALla�md|"�%N�WI��[j�S77/Z�Lċ̉�8ׯZ�J�0+/x�W��	�:��>�������uE�Z�1�E}�F˧���Ò�Tn��Lg���м4�w��������/c�]�{ Y=��y�Ԡ$�c�1y����O6�����x1�Eay �F,�^�� �j�m�{nv;1�3:�$V����n9�;P��FWçǜ���ʓIY�J֖`2}�-y����<��}ڈ�ݡb�aS�4���/���W�B;��ec�.�;����d�*�����2n`F�� �����w����6*3�K� S�U�y�b�� h�u����&I��-�+�s���֢O%:+�h��*�v��f�a��mձ��:�ѽ�S�
��Pt�Ga����g��~@K�7�&�)p�^ԫɛ��rfG�*�I�k.��&�o�9��A�A�C��T`��Rx�)���I�$]
׬���J�(9���`8�)*�D������H�زO�`�s�}wk����}:�f �gv�ێ�cAR.��	��mN+�ۍY���$y�rR��P����m5VHo��-�	?z�����!�Ig�9���o���l��U��sA+�rݔc���PCF]�����Yr��\�%�TE�{�掙S^+�SͫZ�F_�]�ӹ"Է������AJ<8��3��.�6��%M�}6r���ܻk� j#	[��q%�m�}�W�`�o�[(o��5/A�m�q��]��S�ħl��.*��F兲����c�OOo9�������~"�"��V/|}6{.Y�3vpY�p/��L��]�`Л�����9��'�jQu�Ÿ(S\��βx�E_-@Y�Iva��_"��-�.j��AT�p�{
��k\y�v��
h�Yzw挷�mQN�ƨ��D�.�g 7�Q��&0	�1k#k�r�M�#7Y��р��z�V^'��v)jJ�P�çC#����SHU�ZE����D//C�I}.�����ϯG�hTj����L�l�k��B����ɷ� @�Z*\�;]#u�
�ic�.ά:,��Nn՝��no��+Zܙv8�.o]�`��iɻ�n�"�4BI ��ī�**j��Vl�!e)��(�b�AQ�䓒DI$TQU%g*.�T*n�%��V�kOv�"`�S��r
�ReTh$�iQDfV�XTdE�*�IЪ��D�JáW Ņ!fȹQA�%��DR�FXYQj�rEV�\0���	�H� �6U�����f��P���P�Y�ZI"e%t"�����$�R.h��
H.�Z�QR��S�5D+�鑥'U�Y2�+���K��FYh��R���p��K�.��+�[J��] �:q#��Ċ��(&M	D(�Բ,(�̴����"�3,ˤ�Pܝ��U%%�\�S2T$�(�"ԴKCXGI*����W��ӥ[:\͒,SֱE�vX��Ȍ�"vS���کb�A��.���2��`��}*����[�`���9�
b��okbf�d��q�O�"?<j<(�i�aT���"���޾Aղ��_�> I;:|���m�I	?��O�i7I��?�w�]y!;���3g��ȁ�u�sʸ���(����S�D�>����Kďa�nN����F=;�ڭ��=?S�0��wXz�~$����*ɾ�����V���x�q�ēz�?��|O�D��X�4#� �G�s���8c��^f��[����""�}�ݺ���>�F޾������[�og��H�;���|�M�	'|������C�[��M���0�yv��Wo��Ν�p/���Q�<� $9���烢���q��k3z>�}
 Q~�/�@��>�q���<	'�^�G����mGF��'>;s�������N$�~��� {I	߿�vWՂM;Ͽ;�������.\Y�����@>%ڸ���_OѯM�޷_	>G�}�}�+H���>�O�70<Ͼ4G���z�{�}�{L
ڏYF|q�����?�ra=��͔P���;�߽��m�N��?�8?=$��#������D���~ۨ&�}��E����+�	"��f���c�ǽG���i�z�?����n�z��x�v���~��|B�O~���������;����]������y$ݝ1 ��GӦ/=q>���r�լ'br���$x^L�t#O���=�ϼ���'�9?P���~'&w�Es�Ǵ90���Q�e���܇���N��u���ݽ |I�]��;�
=�Aq��<�9�v�ퟶ*�+�3�uD�UN�n�/�0�#�p� |>p$�Ӵ������r��~����{Ohx����<w��C���xzL.�=��]�?S�aWz�G�&���אw�o�rs����N'~������r����|����� ��'*G����I��;�i��w�~o�|�ݽ;���F�x3�>��#�l{�^��A'ް��~��M���{>�������~9�Dx�>�RE
>� ��th;�b����싪���]{ۮ{ |I�~��~�.����x���}�zw��n@�{ϝ�7�%O��~�D#��}}��|ϼ��]��Q}�<��k��~���v����7���>���.�#�~�{�I����R�ԩ�w�Po�}���'����3��y�W��C���0�L��an�U�݌>�U�+�:R��`��<zA��A`�s�����qb�`ֻ�b
�\O�nһDW{#�e����\�]f����D�kM
�%��g7���l��Sߨ���OQ��ߩ�a�?�����'z����z�����k��ϞN���<I����x���'�|=}������_-?�?���}��|�L��]�m��ߟ�����ӽ?����~�=���~8��zO��ǧ.���B��O��Lǀ�=��� ��{f�}��s�2=�zO��@��Y��{�@�:-d�բF	u����O��iF�����o�$=�8�|��rs�í��N']Ƿ�ې>$���x���q�^!�ɯ�뷽����;�����~;N���'�m�;�}鵞/6$�+�E���^�b�#}#|y7��|��bw&������=&}������s�'&���
���޺�0�[.�~>�x�$�������;~z�O|Bw�����h�AwG!e�+�������� >���������~�|y߮>}�9'۷�w���<M!>����Ǥ�F'x�G߼�[s�<@��9ӵ[Oğ���?����I�����'���������rU8x�j�]B"�>����������
��Ͼ����v���v��	2�O���}��?Sӽ�]>�]� rN�O���c��bM�z�'���������oIɾ�;N��q�Ϗ>�	Eȣ�}����_�H���;�2�q����?�^�e`�!��C��raw�?O�?�ߎ���s���;���I��'�}���o�rs�=��ǤԜI���ޓ��ې=%�y������	ߦ������G'~ww'u��P��"5��C�c�zv��ǫ��;�i]���m��w�vܛ㾼����x<�����;�������㏩���9g�8� (���_����a�l���녳�ּ��ӑ��$��>!�DD}�����N��ۜ~o>v���r����ɼBL?�x�v�]��;ߖ>'��������a@��������
o�O��Ͻd\�������/{�$I��ݱ#i��C���u����>�K�F��}G�������<L4>X�};���;o�;�z@��>8�y��o������>�{C�~��	2�O���z@B>��*c�}� !W1��:��^���^ g�d�Ӊ�[-���C�k���%�f{H",Mʸ[�ĸ�.(���K�vV�����ͣ.�⬽���SR��X����1Hge5N��c%b�db��R�zE������Z�y��|:�S0���×Jsf��RG�=��\�D#�q� /�;�i>������`�x�+��Az�
���<}��<O�q�}���bw�;��t~�����?���ޝ���s���ܮ=�&���׾�߿�Ϸ��Y��*���?�=$#�mC>�q��y�$��v���x��_�翾������O{�~;N�w��x����:w�Ͽ8��u��r�����3�'�G�}[��>�ka<Eќ�]]�ξ��>|ȃ�>����9�;�9??`9]�P���x�~[w�v��߉�K���w��ܟ~��<M�	S�?��v=&�B@�C�(��I�y}� �$�>�>�E�餳;�]�z+�yC6�h��DAE������������;�b=G�o+o��x���nw�j��ߝ��aT��x����h�<��?���\s���HHG�F��z�d{H�<��&�~��#~QN~�Jfs_0~��#���}���$����X��'~8R�;r�`R}餏�'�+�@���ȓ�@����z���>�P*F]�NN�fny�5^pP/��cV��.|�:����8�\�!�e�����-�E�8�8������c�K/lzz�ڨC����ZMHt����T6���Z�����d�m����ޫ�#�dѡ�	�tJ/y��:��ݸ��t RF���~O[Z�>S8n���I<2��F �TNK�CxD;�z��bDgWu#t:��|U�FSu=�D�'�Is�N�u�vI\i� �k��Ɗ���� ���V;�a�]�WUW)=B��Ғ�=�òLY��u���]uf���]Q�3c�o���UY���c^�j��������ʜ�N�i��/����q}&�	{_����*���K�	ʲ:���AA�6�gH/^cVzl����t���s*��#�nbE��,t�Z��Oy�Ui���\Y��fR������u����l|�]hѰ��,�#$���#<�nY��g������S���1kd{� 4���٤����x��<~��@\�̫�J�rɶ���W��L}E7�e-L�i�-h�ϙ�N�p��ድ�SsF{� �/Oao��]ݧAl�0������0�d�ҧ��l<7���lt�0v��;Ϋ�Jaz��zs��(E���g�ߎ{z��7� �T/n�5�}���~�����Fd���C}�'���l��9���'���+��|����'��,�Hm��32ܭ��1� �pR��L[^�C�J������9�>��O:'����cӒ���Β]��{Ī6FUDJ�5�3��>�xk�ٟ>^?�����~���/3�j��+���V���ϼ�,k��^�j�F�y]�2�U��2���'�!Dч*-��u6�rd�W8�X����M9~���cʃ��ZI��MHQ��;Pf}��RV!�k�-	5�ڶD���j��؛e�lӬ�7C�<�=���P�=R+5�G%'�#�ҙ]]��w�u���������7���9u��V�uۍ�5�d�{NKu�0����J��n��.8y�y�;sώ�9	e�ʇo#l��Q��u�`�]qv�t��Sp5��F�~����7;WT2�ii0��d���srm�9Ⱥ�w�x	�<D�Z{����:��{��U��rGs�Ƽ�_.�b�)������npM����V"�$��� ��S7�k�,�\����K%�����z�b3� ��W��9D]������W�2`,��'Y�Q�f�
W���:=�X��̚׊.��޽u�wLL��!���Z�� `�%�K`aRPۨ�5]o�v��dZ�N+u���<:2w���a���N^鮱5��h�hH�.ɂt��u+�-�t�;�}��y��FOV��JNt�f�"���`�6�caAUx%�̣ ��}�cGN�������%����b0���Ǣ�L���{�����j����#S%�C��K�ۦ�oO0rV!��і��E�p��t��ԫ���u�/P9=ьu7b�h��X��څW��Z�(#�fԇ�`ar�ڳ>��W�3w%���c;�v-{n�5:���Ur#��2��W�[҅g��V�,�*w�ƭ��ɩ�4m�Έ״m�/����E������`W�����d���DM�N�e�� �Y;7Q��G�u�}�w����Q�	s�0lV�b�֊N�,�(wk�#�:��a��ְ~וg��B��T��ݠ�L�%�*�cީ�Cu�Ŝ{�k&�������=�{6�@~�Ϟ��$���lE^͠��߷+߰O=遺W��U��s�I<6zp�9�ɠ��|����7f�ּ~��mW�[�M�A��� _i���Qe)�(>�O�i��8���Ӽ���h�*�d<s���rz8UF�2vlɲC${_wPR��B�L�1qN@�Q���P4�Y���ka��;ɛ�k(V�*5�{g���B��x�<��+��Z�Jm{y_�A7���q���u�[��z�
�>�8�F�!k���?\x�b��Iw�Z��D������pog���i��|qሪ'Ͻ��^�<�T�j{��u�W)�׆�
�	ܓ+��+�
���-g�'��/;��5ԱJ�ܯi�F��Nh!4�Qsx��Y��('r�]���tߢ<��y����Ի� ѼUu�Ӻ�8�#��tc�g��B6}���OsGܞ*��A^<p�G�����X�uQg�c<�3^/T�7!�~����C�)n����h�� ��r��=M��J��C�nXP�8�E'w�8�ݓw��϶,�6:�r�{P�{K{bJ�
�ǩդR(�X��zp�T���[��9vM����Q�Eë���b|�OK��r�kЕ[�f�z�^~Km��f41qg+>f�sl�$<���(y�v�N�Ԛ�t�'��m� �,�6�)��\�n)�'ۯ�r��:b���p'g%��Ȋx��#;�H�[�b�ȭ��K;X��z˔k�������r���N��Swm�A���E��u�]��dg
�ds��R9ܣ�t����xW�c�b�=��u�تͩ���nM&y��o��=��LS��u�V���-0�:�k�i_v�[�݋�sw�h��UxB��V�!��T��C�n�����s'Mv�֜�m]ߊr{9�������*�%�]�z6'&����Wt��f��3f0[��g�U��Zi]8��gvt�����?��؟?!�S �;�>��U��{�V�Zb�THf;{�X�a��"�%�k\:X��rv}i�l�:P�|~twL[��=�+-K���+��y]˽O]��*�P���;�K���
6Y��Vz\���ȧ� $����7�I�ٽ?@(]i�g*T��d�ܦ��^� g&dmws�:����70�Yp��xAG�h�{����ZV���o�����h�p���J�Q���`��o�Z66]�5j�1u�ͫ�!���γ:�*[��sS|�ù�|��}m%^�ō��<�bmz�{�N�z�C���+I��u��֠��y�yX��R���΋�٥ZC�s�}�p<�к��E�y��8�u�-'^L 7��t����8�^7&����6���H���Q�ה���7��`v�+]Ozr���^+�n��U���u�(�Έ%����y������kƲ:��@�#��FA��g�]�W�tke��%l�=2�k����S�c�1@�ς���Zt�qΗ#�!NҹL��#*�o8;����(�K�7��'��Mq=
�l�-�N��XQ�m��U�,�ah@��ݵ�]��'�*�[���?7L}PUS��O���3��+�!��k�_$������zdw��p׷�j\x�=�����q'+˅ y��^=�mI陪��wm�rz�if���)�r���گ;�I��7�FY���y�s�͛�sLh���awB�����o6���<<��ظװ�87��_mV�a��~ٞ�������B�C�v���0�kǄ��@�R��6x�t�)�0�E�9+��J�ݎ��-��a��O�� �� zr���>��#��74`�k۝�א�:�: i�A6s���H����P
�8y���=��(���e�{�b�wT��F����Y�_z:��TE>|���?�	!S� ��n,���8���0/��Y��W��Ok�;�]�@�j'������Yf�]�R�@��P�z��	��ʧ���g�����6^}vљ޸�§wʿV=�x}��T��gӡ�BM$�=�>�uaY�S.	�*n�tߢ�ny�ݐ8ې'��k3�J�0���g9��|;T�r�M#-Z��R#��ɽ�uT��H�\�{�\F���I�eXnF��g6V�n2ީ@��Ƕ��h� ��+���jj@a܋�1H�BgZ��/:��{��U��q��#��ˇ��jw�.̵
���Z�n�Et��J�ہ	�W�Ϝ���{�u6��keG�r'*tӾȅ]����öt��P��lA:���(Y& Y�(�hW),�r��Ė�u���Wk����0�����W��'�>;�O���f�߄��`�0U��kmZ˨Lg�P�}�7�y�$g�3��;�X�0�Rt�4:k�JAls�O4I�z�Ͷ�z3D�*��n����s�
�][�4�ڭ�Ya;�b�aQ�^��?d�(�����x[�(/+:�l��nٲ�IPԾ�-�#��h�6��V\�Ս��Nْ��µ��$� �7r�:�����7�)�.��E����R��E�v(��ë�z�� ɷ,l�n�W?�����ݐҖ�t��S��,�%�����@E�dO=���k���i������)L7��������>N=!L�;	�^@u�+g���\�-XZ���u5-��d: ����4>_g���A�;\\�8(����m{��ܛ�����KI=�o4g�����4B�AV:5�l:|�Ʀi1�u{%77ƽg�3��2�0��_x�Wb��v�k�8���w
ߒ���v-,���7l���|*�Mr!�߭�nA�Q\5�oE�z$���d{$w]��{ ��(�{�!^����7�Z��;�z&)-�I@Wd�ِɠ�k��^��AJzj���ׂ�N�����7��x?�|V�})�� 8M�(�m0vS$�n��#b�GBW��hu��������.z�|-e�yGM{�J�����SKuT��E��ܫ�Bce̄��uE<��sie�w|�F�&랰Nb��d-N\"����PC3��!v���;�#m�\g��Z�2���@��2s�X��]�(�wz-b��W�x�w5NpԺ���+:��V�D�o���(�됣=�kȄGT�{��;ܑ��IE� 5��D�zk.np�ޤFQ��H�07���r[+^�1�,h:U�8z�Ӆ7�פ�ll�"���K�yT�w�M�J�k;Nt�ű���6�h�1�7���_�)��$w�����%�7Z��(�}�p&U6)eu�[���q�͑��Ayι˺)�2M�cg'��ݼb���Z㦤��1���g�ʱM:��h6�Ё�V{�:�x����ٛ��r�&ö�'V��1k9.��D"����|n`ڛW/c��"�u��VV|����R�Cg�	-=&IR��i%^y�@�=���Oo��~��G^�y��e۳�_�W��o��wJz���$JV��`]�/2����+��;�>�7�[��"S���}��Q����[�M�/���w���-gy�ٿ@��[]l��t�Lȶ�
�\R�R=Z�hf� Tʋ�v4*��T��(�gt$�+ L���V�q�� 
�l�� ��dt}f�h��Ӑԃ���l�*��Gy���gn�b�h�j�yݨ����8�䇔ǁfe^h-��r��\�9�w(4�v�e��|$ua���72�!n>�E�m�Dj:���Qd�[Ӗ�[w�Ld��U�d.�i�Wٷk�B�}����G�烹]>�v�X��v2�y���bn��n�3�{��b���K��U�-u��H\.���Mʉv��v6M�YZ�gA���ʅ� ����~���bP��e.�MήŨuN�2�4v�� �'rꮻ���WF�VY3Uf���:VJ[W0�{R��:t$(�]����[$gs+z�bLx��W���vhg8�d���{��x�o��,�nv���v7j"i��|�r ��u�n�z���u�*`8[���"�5�Ö�D�f�n=��9+��6��^G��8pX�;����&2A��q�m�b��wZ�_wD�2��ԇ�e�7���lY��,��t����iV��y6t���]�}:v����pǯ��A�G.Sl}�k�潴�`� p�W�R ��[1�k�n�ގ�@nH�;�]G緦�����x�c�oYM�}�Lf�����pn�.C̛ꔧPK�%A`�M!]{���Aʕ,���S�J�=A)��Y�X�0��zO��N�����c�p����u�ٽrI���I������d(�m�}�����/rg2��K���I�f��:�V���n��Em`6Z��I��b�U�����4/(�;���Wڲ�p���u>����&vuɏ���&q�F,�_+ƻ��7 ���ҹ7|o�f����h?J����O�>[��Ȳ�!Ï??={�����,���s"��TEВ"�:��³TXjF(W �EYTHt�QU�֡B��Ľ�M"(���%AQ*�:nVҴ��U�ar�am0�dJbD���r�:�UD��af��iB%����l�C4�6��
��eq:�*�QI�%Q!RA-N�#6T�f��a"i�+Z�j)EVar4�J�T���eK*�*�نF{��\���m(DB
����ĭK�&Rh���Tˑ��Q"�C�,
��J2�L�MP��H���%%�'"(�TeDQD�����U*D�rB�)S��t�XJӗ%KX��V���r�E�y����T%D0�T��+�t���"D���YΔui&�ZtS��s]��B)1����RT�ΙV[D�J5�eIE��BĢU6H����P�IB��DB��iy畑DF-)D6A��S��YJғ*�D˒aK8TI(JI�u珷T�7Ϛw�`�O����;ׁ���d74{5��\�|_�zM��y]��j�;Y��g����9�����<[v����0O�7���ƽ��gt4�PQ��z���9w�$�B4�U\`�&l�z�Z����~���-^�*�����i�MQ����h%�K�q˯o�M2�Ƴ �w���
�#z��ܽ9�7Dy��Nh!4�Qq@[�IfA��u�Z|��\�8���z��g�h����t�#毣&���B6W�����O���W˽�4_[�&�VG$H^9���dq��]�E��U	m�Y1�Ng+>f��΍��8������{��X�-n�c�#t(890tvв�`��Y�Q_�_R��a�yD�D�3�4���h|H�>ޓH��:C�Dh(��E��R�n���ً�x8��]���:-��n�	���f��S, �)�y��
�����Z/ܯ!�u�A�o{�K���!�f���^�*Q�c���&)��?���[<U��Q�ugC�Vm�H��w�rƓV�˾�rÌ)��R����b��T��~����GD<��A�Y��K��&|~=gJRB�*<�у���*����ע��Ж�H���Ľ�t��}(�ώ�=��4��2��{ ������RM%�s�<�����E�^�^������G^ʱ�l�(m؂ٟ!��ݬ,�m)L���Ûw�Բ�N�_�Ux`��=��DJ��賑q�қK@!]���:!q�]�Fh�Gn����2�ދ�j���oCLg��iFlJ|��`�2���s�8�U��x��y�u�Əg��v_�~3��V�hYׇDٰV�1jM�,��4����܂o�u�� �	~�a��'���g���H�yQ����ӥQZ�Ji{L����c�_��ޓ�)�Z���۞�Mׯ<�ϫ|~�C���+I���N�x#Z�5�8q�=G׿ؽ~ms5������\�_/*�a�Lrc�Q�T;6x��uQi:�H 5Nl��{�{m�U�t����O���S�P�r����)kmW����=�#m�"�M#�2���{�R�?4
��Έ'`�H2P�^�F���g�9t�U�v+(�ې��f:7]��d����|��]Qfۉ|
'`�A��q�3��g�w�N�M�jFg�c9Z�vk�{���o����9�����Z��@��2��a�*.�U1�D�Wq�G�J�}��3b��rE2Y��Җ1\Vu�������i����"�|z��EdU�[�a�*����`���Nl��PY$�w1�&!�~��bd�Q��WAQ=lmt{��b��(s:�rk���� vM�4T�Ջ�9��[��e��ơj��xx{�{��{ơ?�9zGwN����� ܱ�T��D��/NA�����-i��0��t[�$��F�5��\)_G�f��<<~��}t91�p�{��I5����aC�׊��S��ؖ�j�2��']�APB�K���`r3��
�[͎�Y�(n��^� D�g[�'����E���c�~�����	ON��ey�?)����wלƞ{䶣�Bc+�u���Vl�-�B�8�qe¾^�贮�'/��5u_ݓ��q�N�G��P�3���K'�.��$�'D!W��q;3�ɂ+�(��A$��QN�?V^[Ԭb9�א��w����~�Vܣ�,Y=��'���:+����s�.��[�����y{X�����N9w]k3����F�s��c����ZI�5�������n���ov7�W)#�R.#���$���)���#��v#��׹�#L���V;��M�d�{���"0<o�mLA�$B�QSy�E�Dr���f彠�"⣅f��!�n����S�5�ҁ�ߥ�Ҭ��q�p��
Ps�t��Lez��30�5ކ������eU�[j�%JҪ��B�J��N���^(�.��J]ǆ��#�u��m8ѡ���ovN��KV�,M�L?���"nW�B�锜����������-޶�[�?}�|��j� JҬ���L@�U�^�.Y�f��Sih.�`���W{��զ���>��uW+�b	�S&�⅒c�#y@:��nl 
�����Q����C3���9^���g-��W�Aj�f\zGt�}N<���:a<�d�0�oDNp����\��vܵ�{Wn�?C-v=��)�J_t�5�]bhz Afy�'�$�tVu��yo��n��Ƈ�-Î��B�&n�2ju��'j1�Jwl�Y�p�t�d�����9�`���K��Y�VJ�O������O����8��&j��f���`�������n`�gˣ<jP���ye���;}k�����.x�Wg� �f9��~��y�u��b�[��'9¤H�A�:�{B{P�Vf\_!X�܋��͈�R0I�Y���s2��nl�
�VWu	�C��Y�y1(%K�%]��L���m1�M�����c޽Fd�f|\8���oOb��ۡ�Ϟ��,���� ��(�7�{�w�wZ����_%o�t�_t�i"�0��w��B8�ȍ�f���L���#�}ห�=v�ϽiV�̏ۿH���7t:�<���>9��;����.V���;�w�6�Y��l�H�qv%�n^�����u����W�}�W������9�Oޅ�� �6+�x�l�d�,�-��[�*y���ׂ��7��>^���ΎFo`8��ozrg;VZ`��(ޝ�S�#� ��7�;�3���/���y��@�#��59+Z2�e���)Ea�6�T	�@�"�'I��wD��OTt�����̧�6j�p�^2�9�z�
��-z%6����B����JA1�쏫����Ob:\�d'�@:�C�C�Ӝk�+!���]��P7����pi-엑�}W���=Yo��P�.6��ф��!术�������s�c".��_1���b�n/Rޓ�'�	3������5�z5^���Wq�2�@��?k�\�
H�^Uɹ��������&�����k9�YfC�9 t�@h\d_,��˕nJY���;.KtF��^tP=�V\n�m��3�,����S��UM�� =Ϋ�B�� -��F2<Ή�=��[�=�8�5� Wb?z]��4�����u�N��7n�.��/;�V�mKWk��rW��p3��nQ��U��5Bӭ�{��w�s��uf����o}�<w��Z��.q�t�;XC��V�O�pm�I��eӹw��;�J�E�/.�7� ��s�ڝ�׏�6�X1�B��H�ιJ�=�e��u�6�"6���=N�WQ:|�D�������ʧÖ�pΠ\^p��R�Ώh��i8a^3$�����?N��>���ۮr��']<�����Om%��T�pc��5�sng��.39>�{�Y�9Z�:~����uǝ�c�v�����l۾�ڟ��t-1�\��~��}�ys-(V#xݱb�Ռ���ٮ/�rg)m���0�7��Řz�w��g��o�-����~]G������rI<�
ҧp%3�����&��|�k���^Ķ�OoزnutC�.���w�K۽�V�ef��Cu~�[OTK��VmCk�U Y��
�"i͜޾����qt�Gk��2��9���7Nn!�=�����f��+.{�.V���bk�"��]tûm����]τ,n��r�R�<�=}X�/x�
���uMa�y[���8�i�b��Z�YyV㽭x�#j`[<���?�P��f�⤷{� cT��1��j��_&ѺIT�d��Cp�9��^)Yg��+�l�{yL:�|�'���ܭ�	b2�0�݄�F���pXΖ���ǺTog �=�䎘Ƹ_���g��Юڊq-�`|}� [5��:��j�Kr��Z�_��j��t�7Y{n;����ڻ4rw��^.�x��oO���ΐ����du�-y����)�����z�kW�f\O��矹�#P.�U��P�U,wIo�y,�u�)��oR�8�V�l��&�i�AR�A�/hx�E‹�ɹ�b�m>����;o\�q�2u�I�w��!�c
�k�؟,m�IМ�U����[jg}.����&�C�L��X߽�S�ů�k>j��K[#r�
��;J����åS��@�q�w���r�]���zn��Kq��s��+����I�W0ߧ���Sس{jL�*z��8�H�����:�s��^��'�DF��0�"+�c�܋aWc+�wvT8����$;������6�S�O��ކo�@�{e{�� o\�*.a��t�B;y}F�M*�xڞ]����u�,u˘y���������$�w��kKRL۱aV����DEM���B�sΝ���^�8�R�.>��J۞��˓�����
�r�-U���%�K6C��#�^!G�^M�0�yŵTOl���H�i�=�6Alwﾯ��������O����V�E�ucn�{u�S���Vy�e�|����lS{v�_f�����x��_^��-�7^�C������ǋi�%鉞������UJ뻚��B�\7�ֻd[m�Ԇ���s�^�S{\q��F>�Ң:��
���'�� kz}vb;]+\���8��{5��r�2��>�8�F�k;�W��_Z��i�z�Dk�/����>��p��f7S{��7�]����V+= S��B.�s��l�JT{"�����V�觺�j��Bױ��[c�ꔶC��������7x)��xJ�zښ�Ư*�m�c�j��,� >�:'�|����4�OL�U�$�����.5@
��P-��.=����OW�+������;b:�\ވ��M�ˌoXʹm��1�^8��-���ٹ*w_!����H��o=Z���}����k�������삡8�9!xgh�p��,�ȇ��7Qcs�-�@{a���Sd>��sf�w��n#Ֆ}Ws�x��~u��~2fIN��2�T`��TE�c��t��;�	[�������d�"w;d�Aܱo=��}T��x����	�Z�l��r`���ċw����^�������/��4���1w^���27ݴ�9=�gH���w�����6w�ؘ��֒���;��#�j�3��y�˷�NS6v�f*��\�7]W�兝=���]��q���ry{�?g�?y���@��;lײ�Я�*T��O}:ܕo�n)q.]Kcj1ſ5Bc����>q}�̐��� ���ؗo�g��
U99R��}�6qA�u����r�-ꊂu�ʬ�.6),z�7�9�{M�J�Ķ�;X=7:�j�EԢE����T��Uv��.��II9��w<]��z�:���Dv�;�:��|3KO��������,Oa�~{^�yד�u���d���ֹ���j-9ȨǸ�֎]�n)=���V�s=����~w���i�o�����ɵLT��eX�"�^�a����4&$1��]OR�>Ѥ��){��{nRU��y�{�/n�Ossr���1��!�9Ix�G3��fVK��A���	��y��:%���9�]ǹ�o�G@S�Ƹ]q�e�l��I]׫D�Ĭ7a-�Ҁ1VHfݩN�[n �����v�l��s��eW�/?\U%J��}��ͫlc�S�7!�b+i�%�F��n�x�,#{�,A�jN��WN|6;u��o�Y��s��7]-+����d�_wi;1�-��෠�^/�:nU�����]��;��3<*�m����r�:�HN9H`�/���E�u��o�'������#e���v���gQv >#�r��m?�˔�u�0�\)ܜ�juC�z�KU���"��]�/����p��R�'�b��S�����ЧI�X��I*�'�7Č��OkS������w��{���耎t��x{��~h�C� �_��<�=�+��1���F�;�,��������2�~e��3�{��	���߻.g֗�z*-o�az�Ռb޾E��Χ�T�MD���e���H3^��QϭN����l��B� ��F�쫰���nfg�����.�2[����l�5�s�Ƌ�j�v�t
˱EYNDǭ�y�9�y�#`�v�齉���m�.�,4�	౷�c�t�y(=���S+�v)#w�ܽ��k�!���X�i�K�v`ؚw���K���T��<Eg��n�O�X�:ݜ;u)��<ΔN�I�:�=��:�����)��YFޯVW��������mNL���v�P��fbH����w��˹��[�gd���j:����b�xgiܖB�LowS�]�
���Ҧ�t��a�����]���[^�珉_].�7�l@�l�}v�����e�^˱1LĭH�n{���3F��YU�i�����{�x���-}7W_���:���l>�<�&�Ç����:q�FdjY�)Oi�Y������A�DNCJCD�Ot�7��^�w@�f�l׃{<p5sӈʥ�O:Ay��Q�~��Z�����Z$��R���
�^m
��0D���&��NWS��v�V3T�ذ�\0EJW/ný�����ԊF)�Q	�_^Y}M!e��	�3�`��w�S�����e��.��n+n��ź!Y8��q�g��X�4rі:S���TLq�h�G\$����Fm�f���3��Ǧ��}j�CA[b�}�M�֠�;4$~�Ռg�����+Ԓ��C���d��q����8X�w���>��=��+;p"�溡��up)A�I�����nV�&�	4D�{F*�������7��ٗ u�Z��P���F�"���r��PJ�}՗l8�Q�x��^�te0�ܗ1k�}��;R,�e��C�H��Ǔ�w3���}X\ܳmm[\Jہ�%$V�%�����	�k%�e:c.4Z�V�ËWT�)��J8���L�n�}��J��Gصv�����vWs����nw{\Vh�� F�����l�h�o�������s�9���dܝN�j��1]�P�/��*_g$�4�O�a�ӣ��x;VR{�	�F���M��*�75�;�<k�k~�7 Vs������!��¹ɷ���m;J����on�ظy�O��WR�3]9g�!;��F7j�f�IHY��ei���k|5^��Sx��f�� �j[�ؚukz��-wV ���n��!L�-v�Y*�/����Ɋ���`�J[�Nջ�E39��V��<^�/7�YيH,N����.vͭۜ��hF��dF�ļKn_����b�0Ċ�M��̝��	��u(����
"s:جlq�Zx$4*%������d���m�c2�8p�X�RɅv�!��=04p�jYw���_^��V,r̐M����A|�f�)����	Za�H�Ĝ�4���L��Hl�0F\�4kd!�8���E�
a��ad\-.:�]>��haB=�My5�=|U�C[׹@�J����ek� ��2(�j,�Ӝ"ґ9F	��[L�H��"i�"��DC�Q�$a�2N���D'"E�$�̪�i2��%�!d�EĮDYbb!�Q�G]�,�Z�$��0J$��Bʺ�H��I*���'���f[ �eer�0�r�e�RI�­ES-�aVYe�*��&j2�TYQ��I-E,-��h��1J5��ʽ-J�:�,�H�\�*+�N��jT����9��Q% �B"D����$CC*Z�-̊�Y��9�!G	JB��,ZJK"�S��Y'��"�E�9S(����$j�e��(���9&�եHr-Je)�	��jH�s/WTгI�$�f��#Ne�936jTs��Uh����C�u1hY����Y��Pf��b!�J!AV�Z��!�+P�:QJTʌ8�+���QhQ&bD����dhY�E�b����{������o����@ޞ��J^���z�����K�v����	mXV���m�x%M{��.�p�]��UW�U�9�ך�����Y�?��ɮ�[^|�5N��^�z�\l�`.�8�f1`g;n/��۫};��Y)��]��+5��t:d�S�
ו3i8�yőSwf.�s���� Z{6�m�ѣ��ף�m �롊˞�K��xf��I�T�m�v�wR^�Iz�����k̵����~.��(�g��z�\�c`�������6nD-}S:�9{t�s��7��C���5�o�L�|��6�f)�|{���j؃��@:�{<����y\���5�C3f꽮��s����HM{����Q�:��V��w��)f4懟�歗��8�|��T9�5KR�/h�E��8Dk����Om��^�U7\��a�Q�'~Ϝ|7���|=O�,�n����;!�5��*�6��{z�m?��MDN��Ǔ�W�ݣW��یz\\�
�5�r��+��Q�2TX#ֶ�w��������@_r����]G�sz�#F[B��V/cPx4΋�}�<Տ�د��֪(h�U�s��Mk�]��Q(�|��yٕ۝* IB���e�8̀���s���^��<[��c;�{�oi��}_UW�V����ƣ7���S�ʗ�kNM*�~�T��ڣ�U�~�j��c����lru��)���-��s���#n���ހ/7�Vf�Lw����d�I���y<����Dע#칕V�mV=��`��1Bo�u�� ^9�u��Ě���Y�g��~??g���<�׼�^�9juM�Y�=�a@b��%��nM?-rlndS��Y��yk��7��v<[N���T�=�C��70�]�_{��w�t]Q�cu�,�ϝ�:�(s� v<[�-o��+H�F{��&�S�w����+v@��"�6�m�m5-����=���W<��EKN�[I�m���!���\��xֹ���k�J�"�`m��.�S�h���U������K|޼�.��4\�%��#Z`�r!n�zgY�h��=Bn�|�l�rq8~���z3jތ�N�4¿�t�U���4�y�9彦�m�O7���&����C}����ՅQ�<�)I����IK�9�P�.2��n�W�������G��|�}ߧ�0��l���2�ˉ.%���k�88� q�>=���%��c����ul���f�쏡T�����~g�VS9���ߪ�磌��&`ft����;J^��8���Ŷ=N�M7!����F��}�����^)��
�U�!S�*���v�G<�3���T9�4T��Ư;�Y��m��l�����	�\P/������I�v�0��r%�QO�*Ŕ�(�s�|��<��HN�Yg��Dv�M����s��`fa���w�p#�-S�z������Cs����ra<��!��������_'��<��[�Ou��ܥr�����#�Џ�J �G��s:}wR��V�����߮��^<z�4�)^��P�[�}p�����{��w bᏐW�v��Ͻ�ߋG�Ź�j��kh��̞~4���S�y O��v�̋D�b�Y��:�=�\VLT\�gd[���1Ak���]�`s�EOD8O�\�M�?w��;�V�>�ݶhD���"�c�E��ln����>�{vÎXMI�8�N��AL ���+mxۼ���`fPR7r�v�{�y�_���9��K���R������_R��xa��h�R�f*9 ���]��fEҥ>���J��Uo����>[Ձ�k����}+���w4�N��7y,˳M���<�z��si�	YW���\��ض�U���.䭩�.��ٸ�ߗQ��~��-Z�8�L�� hg��GWm'{=�W��.@S�Z�BݟFzu^���>�w���D��7���症�(v�ϲ�w���eϻ�=!h@ֿ}����]�9LEs����)�CM�cVo�~V�c��q_����]�t�/y����c�B}�&y˗�M_nw��w�:e�=�o����Y�9��;�~ݐ��z�x��5���^�~k!�`�D����TbaKi��or�G�S�.B�J�+������_n���D�<G��v��tټ�0�r�=^j��谜r:��2y�"�j�/d{J*�}=W؋��Ot�f���J���ˆu�G�	ιH[��dU�K�c�k�����%�v����>\v@��S�[Ô�����/�%�G��Q��w���m�2��|�*��c@B�_&��/��ޅ�*iC#�~�nh�/ �S�{n���͋ېЈ%�M9�9�R��[�+caL���a=��0qw������^ @�q�"z�s���g�=t�
ˬ{�B(�J�\�r�ounNt���W�_Wǽ��Js~�\��_�$3�I�g�=L�[�|��D4.�� e1t�J���հ�"o֗n[Y�Ҟ!t�L�5#�;�,�xj��]{R%J�Z���a�L�r6Fb�����xf(��x����x�n�nw��Dd��y�8��f���wa�<&��H���C�lb�^�;���Yyy~Ԭ ������]�Oq�Z�ue�`�*[��}w��<	äpCOu������X����n%4�K���Y����H���&��|�mO���z�M��߰��:�E9�~On%���Y��p$3+�fo8�81��&��O��^�܈OU��K�יk���^$����a?6dP��|�ʾ�+94��tQ�#�G_?��UB��iy��C�w!���������_q�Y������@9��y"��sʇ��fiF�;4Q���ބ�u.V��7P��s��-��Vl�WQ�#�BoV8�^1*Qvjf�u����j����O�:�w�;N��e=+[X�w���:!��;ۏ��T�Iw��V�:7��������s����=��;��o�I\����
��>�uNB!d5�_m��O���B��ļ��+�W/,dǓݿ���lz~�e�|T�4���S.0Σn'���1��h��̃�C�Zh��߽�e'��̸�q��1ES9.�~;�c�S���t�2��\�욝Y8�#���R+_���Aqj��b��<Z摊m�$h��\���9-eՈw�6��3I�YS���l�Fs3ws�ZXy�P��\3S>{il��s���s�vnE�E|�{�}���'Tg�,�����1{��5���~�7wYp��F��4�G��g�M{4�Vd�SoӐ�U=����Ԝ�_��zk��&��m�^��;=^�Saugrc�|�S�[�UcW�]G��~}G�;���u���x���b��֪�(o�^\�Xr��,�9;R��}�6qA�S��w�ܫ<S�.�4vNzI�阱���y�*).sVU�(�u��f��h�5w�t���Y[�|y���,�*<��;*��4���h~&>�,9Z�VӔ�h�o?~ov{��r���w��J�t�$*���嫶�!|c�w���E���7�>�e^��so� <�;ϴ(��|�V��'�m�ȅ�0ƹ�g���i���ۭ��E�t�ݾ�����g^���{���L�tP��N�/W����ZmKx�R8wk���U��jQ�ð�H�e'}�h�xKah@��Gw��ZVq��a�d��^빪ɵn�[�=��e'M�x�uk�r��g\)iъ�Uݯ���j/@���/)[�[���­��2����X#1��8�]��;=���.3ޫj�_eY{}��W��,���gD�!A�ȁ�f�N�[ϵ���-�l�Pחw�f�z��?<�KBF�����:�~m�+�*�5d=���j^�\R��8�mZ��g�!�#یߓ�ldï0�X� {�r��{h���w�E�Dn.�d>A��H-.����Mi�4ہ��=�ɖ�=��ܳ����m4�g����=��dd�N1��H�׆�U�u�_��+1�5c�Ӎa�Ũ�%��Ǉc8��-���@�er��n���xv=���v�Z�ch�C����{p֋ەu������9�3ם�УkF>׉��<���Gj]W5˸��p�#�u�=���^��[Q���]Ǯ%��槫è�|��}��D���2���~��5/<�Z�/D�_bs>UBg+2y��g�?y��{�䇳�5v�j�(����>�V��S,�7!=p��WgX�-w��]��[�G�K�t�[Z��O;l�%�'n[Y�躡Q��\# ee����	�Tu6o1Z�I=�sחὮGgb���rVԁ��T-��zE��1y����6�CugMDki�D�{pVmCk����
���:�N��v�wG�fݗ��|��Y5�GgT�nqNo���_6����~8h�k�a�t�X��|�"]�a����hL�/���y@vνU�wOub����q��&��:!��O�r~��7�Bו3�|���Wۖ;���q�r9�U�\�:ר��6����/ �����!�����6Vqr���%��W���Af��O1����<t���Z�a��҈���gX�������٢E��[��/]?m��]��UȮ6@����\��S�]Y���#�,�@�S�т.]���K k\y�踖��nvwb�n2lڊ�Nu.m7������uU���gᯎHe�h��'��4�s�W�����
5ޒ�)��<f޴	�Ѿ	��0�Ȕ��|T�Gd-���k�[�O��m7�㓏 �Z�K����;����vBq0�3�vG��eښr��#5�Qg��&�~��o��ܸ�{q�u�3vT��9O��gPj.s���BCv;*�yt�.�'k�Pѓ�Ϸ[Y���#:I�f��xmo���j�r&�ò���ff�&�O3	U�6v�.�>C��Jy�L�2z���U������sU�Yt���na���n���s2���s訹�o��[Wc譆�=�q�n�js��-�w�����H^�y�f��Ҟ_aŹ��vv5�G�w������<`'��-o�.���>۞�kkά�x�����GK�^L�&ܣ�s���"��[�����|��uv�w��gw���&���*��4`��,HVa$>���˫-����wX��l��#[�inH�O��A�k^��%���-��S�m��:I3�}�m�4�WA���`
Gd]�������"k}�Mƻ(���w�mpr�ͻ�:|S�q�ꪪ�����	��q��UR,Ɇ5��g��m>��}��{�P�;�
�J؞�w���n�e�=!hF��h����r���<��/ޗ��ͭ�N�FޠV�L!I8l�\�VzE?k��ZG7b��&u�{Z��:P}��[1g+%I�Ω�KP��_�[�Vz����9����wʓ�\��:��D��i�U�ů�g<���C�}���s�9j�K�������[mlY��H�������s�v���8��{)�?'Tyx���ۏ�@V����LU���nB�z�*�sT���f�&�O?r�@��<t���NZ���kz�j-C���,��j�ǵɠ����z��Z:�N�f/8�͎N�/�m{�x���uo}��-�^�\��4����茋��cvbx;�sb�%����52=�io��t�w"����z\��1v@�G2��Y�v�X2�IЕW���d����G�;z#��/�Gtg���A�U��\ҝ/3Q��h�|��H�͠��I[���IzE,I�Y뀢�;j(�ܫ�����ڌ5��nw_e�Ze�����Gb޻��
l��`d<kqzo�C�D�ė!��sgv���6.�����z֊{=��Nܤ�+����93,~)�g�%����7jxx]u��چ��-���tQ�#y�4~�����P���#�<�����,@>8�ѱ���ZG:޾�e�P�N������w�2��j٤#�%:�!� >��c�:u����w���m	8�k_JbdI��(�՛G����n;�IO���5�+Uh��k�ѵ��hR]�d+���A�}J��As+��%��Ff�.�c�	i�V��**��(;o�)O�m`�X(5�)�w�{zO�˙GqK��Xg\%+��ɐKͭ�*	uw�K�:���i �̤�nҢnK�CS�����	Ic�X��q�pi�qnuW,�<�֟M�W���҂��:я8ݢr�ȺgÂ�#����ͅ!ºV�.�.w���@��$ѷ-�v�(\�:��FP��<|wjd�䱽;�w�MS[\�]�8��=����߃�'���EVz��_^8�BL
�V����à�ū����[�y�r�8制����^N��aT�<�@�}�6��4tb=U�T���)����@e�uQ>͐vt���(�9����ܦv�E��F9���菴��D�K@5:�c���7Sf�Z�{TM/�V���e��<NZO�[�\qMt��a���ܰ�|=@o׵�3�pe��s��#ÝV��� fR�':��SV��K�ʢ��C�����lNĖ.w|v�e7h03�{qZI��5H���:�;�]t��ԑ�{f-�&���mwrw�$>D��
\��u�]���;��j`�*�u�>88>�o`^*��Q���ƴ�=v!�#&>��#�r�z9�ˡc����.����х �cT��D�k)��n�q��_�>���٩��q��tmMo�u�ۯ��ͦ�іYf��B��B��<�
�'��X�2��o�����g�6�;WT����}��)���	���.s	�x�K�{E@�6f��dQ��&�˸� 辰ǳ��pX[�1��xf�EcG-������0�7�|#��&�ݫӼ�۬%W 1�z2t ؁(�u�.�蛼
NN������"Ռ��0��;N��ŝ�
��C��)YEt�^���w��d����t�;(z�,�pAS�����c7r�i�XiK,O�-S��0R�%�N��S�o*�3M�aF�^�r��s5��%�2��!%�޹:��)�A�L����v��;����ϱ��P�F��$�šeZ��da���U���.=uU��2���$�q(���*�aj�NW�Fi��)��ZT��	�����ʫ:WR�IkJK��8���eUs�F ���*��D��2ZVQ���g",�������J��E+C�ueL�J2�H���\"�D4���eU�sÖd���aQr�R�Q�Y%E��0�ĂM�IZJa)R��D�1hW*��D��(���d'J�9Q&�EG8��
���7Ej�Ff��-�a��w*
,�Y*BDg9Pr

���@�t�B^��vUPU�K����* �д�$5
jH"J��ʫ�T�����̍YQ!�Y�*Ω��Nf���
�Dr�u��s�&��榑t��s�����D���iEUX��M��*�a(fm	�����G9N�҂(��5�2�LdDQZ�]%R*�+�EPgEi�L
U*U�;�zr�(��TB�H��=.�98"oF�J�ɶ�t��&�Ѷ�H�w�� yu+ϫ�L�\wu�If�.V���;n�MTY����)���cVھ��������)���mP�����N<������̻{��׺��s�����CfM��}3ӏzYJ�|�D�V~����<��3̑��v��u���R���K˗5�6��X�B:������kܨ~^:�g��������:��3�SS�,����kl�uI��w����2���g�Ԯ���z���x����N�+��c]�������7u��G[��'w��u��Kю���s��"��#�ԭp�������q�[��Wݨ>�}�����Pw݆��OIr���<�v�W[Y��/�'/N�D�u=��#������(�Z��{���)�\��`�vG%<P5��/9��]ړ��N��v�WۗݸdWq�2�}���n$]��,\�+�n�}��bNv)<����k;��e�`�}�w��X��!�հ��˧����}�����h�G;7�:������K�XR.'\*�M&�L'X��a�f�U��[�5��ާ����'�	���/�݌������;�_��'k����T
�x��c�EDNK:.�㵎En�}���t���r/�����-���r[�5��^\P�}����䞇��yUrZ��ʄ��|�����b3��N�J�/B��|#��m�z����u(y�'M�n�u�@�-b@ןpίb3��s����ywB\]���7ΔY��c�5mS�h3��6�z��z*3�L�Շ��73Oo�[����{���dQ��)f��Ҟ�>�k�Ǿ⏡ �s��a��ܵ8��:P�=��@z?����.�,}�&r�'��<�vW�cKM�4xL2�%����c����Øћ7}"*.}�g�®Ε1��9{�$Z~�=��s(]^{dYȟo�S�l��2�3��G�߬N�8�W�>��Wե��,y�|��u �orf�88�]��P��v��J��@ڸ���t߆y}�0}�S|�C丿O7���C��R<�>���]n狫é��̱8YQ筞V1P��fJRU	�I2ɶ\3%�s�vL���1о�[+����~��/G[�h�21A���ʛA�j^� :�yX=�N7%��ɻw����q�ׂe�.aiN�0&3��f)���[4�r�cȸř���}_U}T\�q^(��͛�fߤ-�*��E9~5����,/6�vY���^F4������R�;�䗪�UB���y�<�y�)�o�錼��b77T��y�;����h^=b7"N�\U5J���8�����(�ȶ���i�sNlE��.}O��Ĝ|�����3��/�����̛u�pگ[g�)�=N��!5!���:��@�(�O,�N�B�w��N���u˴6-���D������;!m�'м��T�{��_��^�&ߞ��;y=k�wj����[��1ˆu�@|$s�W�{xU�����"=�3iB}U��5yb��
u�Zط����-�k�rgh�rn�R�y3n����-�<��K7��=��k�j-�>�~�mV������5�Z�y��L�֖�+l����;7"����<��O��<��<�::�[�+��I8�9׭M$��лm^o1�$>��AǊ��[���#Ϊ[�.Q�s��g&��h�]�u�fWf��`�	�n��uT^�y��Y��!��ntG{�ښL|2�z����޵^�Q�F��nM�d�jῼ<<�:�ʮ��}p�Z����;�w[7|�̮��3M�TN�ʌQ�{��4RKJ�=�̿6�)g'�,w����qz�i}�m���jx��Gg���ۜ6�goE��
�0����N����=��gUX�_9�z���A���_2�K̄��Q��ya�f(��Z��i��]��+6�mx���0纟���K^�g������;���v�&�l\;��<�Nb@|��7�ϓ�\(`����̮�g'[%�Ѝk�Mϡt�ι�߹�{�硘�ëվ>�Ң��+-�o^��4[��|���>���kvsEȍ�޷�]��Ǥ�nn�wi���7=2�Vzi�\��~���ʇeJ6R���;c�4\�������S���&�kbm�8�5�=k����:�*{݅�^T~�����~E�v�0���sEK7��e��y�G-a��K8Q�>�8�P���7  �m_NZD�o�yƸI�^و>Se�s���j���H�0��h,�)�������#jW$n�@��1��g>��N5���ʸ��Q�n���l9WΓX5��QTTZ��?���{���g���l���b��e�
}����R�=CܸgPj�/5c�j�����峊}��]F}q"�����&Fw�E�y=���g����������s�(C��	�������'��=q-s���Y�%�gʘ��fW��n�7��]S�'j��������3�Q�=�FE�5^�G6ƌ�Rb��.+��?s�۸k�#]�*���R(ۙt!��>�^�-�-�cV�Jy�Й����S�y��fך@�y�b��2u�����:�"�y�Qs��;|,S�sϩ����x��S�'�;����պϷ& ��=�a��*�3���:�5z�.�'O�w��K�M�y�� ��Ɉ{��U}ٛ/-�L�*vX�]�!�r�)�_�ʐ��ڕ=��iJ�oW>��׳���멒��}Z�BݟDv��r���͏�zg�5�\�U_^�Vo$X�R�5�ds:��ah�)��{(�{�TatO^�!��m�N{�=�6�Gw8�؈V1�K2�4$X��u���`�-�����t�z����-װ�ᐦ�̒���{�W�xO�D�"����ƣ��J��~����Ҟ�1����2�"�v��6���n�p+Z؃�E��N��1��Aak��̶�#9�m��'J��k�k�~ط�*����~׋b�=��8��]}��1�������B����͆�­��uJF�b��fc���ܔ�����8]�}�z�x��秧��C��ʼ�*��\d���6���L�ݫ����9��*�*�i�	Ϳ(;�X廞j���e�E|�A~�q9&{����WIu�B�/h� vy?�B������pz �]����C&k�h��*[|gϸgQv!�딭c�efej��R����M�n��L���{^��Qz��g��Ǣ�>j�j�ײ�Mф��)�'*=�<!;Ye�j'3�*��)�Y]ђ9܄t�;hc+&���wV0��&�iv���Ι�Bg��O?/�"�v�D�Z:�F h'�nK��'��ǉs��1��-�S���oFxb�Z��@��/��Vp�/��eAc�n|�J�K,��vG'���q�>]�3H��Y�U�]�[N��h~}8A*t�8M�[K�G���d�Q�nHǟ� E�3��{ĕ�ā�D�˔�*Ëk'�P����o�Q��g��X�;@��&�>�(3�v��x�������iup�}{[��w+�����iP�����i�O=��<�j�����V&|���Vd����u���s��pw�MdK���Jo��vK�����i}�F��؞�>�M�"�����c��S�����On
�^^{E�!!쪆s��}��D���ʉ)W�^�Ա;p�k���~�y���iLk=tX�]]̓�vd�
~ޕ��M���ﻳ��^�{�k�G%��/i�S���e�o��s.Gu��)�\���&���ʷh����m��ݠiͼ��l�s�5x�]��t�D�8.@�9��]��X�n��I�ɣPu���yѷi���\�5�=3�TCy��q�:�mg��dh^D��n	㑭ьB!zlj���aLO��֮پӻ��/�ˬ���������ބbw���&YA��.�y�f>��`\��"�у���1+:�|j��~Cd���LEˋ"�Vw<@T⺃ >g�K5���\SdQV�VA�jR��۟��E�Kq#=�̏?}Y��9���Mp��|z�.���s�S�S���ml���n[�8v]�k��W}NFnʚ�f�Mǝ�3s:\�y���Ց7�$L�R��:v�b������C�8���ux����F'�q���V����o�#}k�6������ҞŜ}gj�;��mV�bm3���Ǖ�9gvz;����eGHف�&�*w�:����YH�mB��������EF궑Y�����6�#�Q���b�#��w���K��>����[
�,�b�������[��k\�x��bm�[�*�T�Q��l�v�\mD�{�}����o�M5����Y�[���Ŏ���*���z���޿ �l�
�%�1�6mvϯ�m>�϶Zͧ�w�>ܙ֔�NjhV���a�@!�T�`p�sj?����5C<��=8mP�{��[��HZ�(�+����3L*�W�[��ao8�[�l�F���K�P�"������n���Cb	&7�c�j�LV:�zm���=E�������ث�{9��Mm�Pk݂�]՚��循�j���,]������G�sN�i��g:��Bz�p^7X��cY����<�;�j�S���gI����ST�X��5�FmE��N��g�S����]��brӐ����2�^���z���a�#f�5�G~^	׷FU{�����a{dȶz�Xך�.9��M����u��>n�b�M�)�9�'׻���]�]ϵ���˂߲��[ʱ/���T��{�/���������M���=jv{�W���t|���c����w�u]���ǆ�m�^Ͳ�
�LO��C:�y���9�-l��&<��Dot.=��V��v�	�1q$��;B�UMڴ���m��\��'i�{p=�_N��k�v����U]K'v����A�q�)��ݗ��p�ܳ����w�op�`o��扸��d�xǹ>�y�����yZ^��`�����^�C�y��Ju����YR�3',�+��Z�mݱ͖�p�֍����n�uJ���ٔ�on�I�u�����.�<}i3w}����^����U>��_N<H�@a�����uo����&6�ڱc�ɆtR��L�YNJb9yY�|�Z�J��������z��3�X��U�EB�����B��;����uvk)ؑ����TJ��t궵�����O�N��z��(T����	/'�z{�q#=; ���e^W���;Z�n�; �s�D0��>l+K�Z�*U�Q{�5��u����m=-�J�T7�*�v�Tt��Q'w]d�n�{�[��Y9t�j���̦|'Ey��;�at�֨���\���.�0ւ{�;�W��|"[Xq��ݝ�馽?�4�Bt߅�R)V�qk[mp؎z����?]����5��s��Ѫ����[�s�.��9V<����=������G�ۉ����S�{������o��,��$�GNSԧ���%Ą���4Y��o���_ԡ�Z.��}���R�X�;gt9X}=`��!l�e��#)0��A9!�.Q���dU�ҵl(�����,mR��l����������ݚ-Ea�ǃ��n�Iq�Ȋ� #X�5�p2��F��3�Ó{@�K�T����tl-8�V�+*d��4��ޣ2�8o,嵓g�����_�}m:fW�[���}��+o	,DEKѡ���Y�F�0u��Pd�f�nRiF9%r��0�0v:��Pۨ��6{qܹ��9+E�Y�3].�ar\�\xn�Wh�,�OXv9p"�u��#x�ԡQ�t�U�~~f��"�=���sV��������{�݊/vE݁�"���$�6%IF�X�r,U{88d�B��y��a�e�k4���+�I�a�5��Zw9H��c5ݘ��s{��
^ah���-�nojXsz�}�|u^Tn��r�8�Ä��
�f�Ŧ�Q���W�ɱ:gWh�q�"{q�����⟽ure���l���,!C,�������sUn���P; �6���V�\������9<�\#w�:�t��0c�O/Kt� �_c��9�_nDǚ�z��TH���w��=��|�N��v��7lk���7Xo���	�d���OkX9ιYabn�P���͝f�N��cC�)�`@+�EH]_(��a�������|��Ut�Jނ(�u�T[�d��O����F����&2r:�锉]YrjV��^]�����e��^� ��ඩ�t���Q����W.��GU�)�@�
��0��ٜ
 �A���tw�t�2����W'�*Hk�Z5�ɮnֹ��B�n����dJ�sh���	��e��Uy4!ڄ����6Rw)�����s���������m�JQt ޳��7��Wx��p�n#��7�f����D�x��o�1x����4P�|[�׼肋?�,9���K-��[���T�d�:�m��x֭�|����o�R�v|�7,A�;�6�_]��@@�/VpYJ Q's2��ḭ:���R�s���ԙ�r�5�ļ-�������ef����Nm�@�Z�J}B���JĽ{Ս���Oz=4痭��QW:���1�$�ɞ��r�2�磹�Z�ң�U��Z��������*7����u� �K���F'o�I�Vo�4�,]�X�6a�>����˳A�z��,Ȫ����}w���)��B��W[Z�%��������|�T>c/�^R�|3�)�64���\V�ᐷDFkp\?;�$�s���V�E�4����5�/�p�"�٠�¶a�.���j�m;��gE'�����}�ڭR�B�>�웜VƚM��iۈ�yu�A�J�4*�����p�Y����<Ϋ3B�(9�_�D�lؼ�c7��ȧ�;�="��&iXӈc���q�B�ܒ�J�k)�z�����=y.rL��M:�ZQD�DEp�Q2��PUDYQ�Q�"�����(�,X[eI��T�UUZЍF�E���I�r���T�+�
&�
�8D��DS*��KP$�������W#�iHT�Ts�%r""+��Dr��R�X�DT�0ҹ��AdPNE�Ar�J��Jk"�jGw]�D�"�T��A��3�kYL%�nd\���IAQ�
�\�+�l��
�y�iE2#D�!!�I�N)�Yp�(�f�$�D�Ȥ�TTGu�Y2��
:�1jv�+� �TEsԹ2�LP���L��D�uH�Ye,��Zr�Z�3�P��A$!G%Y��TE\��8r9�QI��s�> �	x�H���7Y�`fT0�O0�gK{�<n؏B�V��w;ǉ�MN��f(^��xe��R���ٺɼ�;G�>ˌe)ro}��y3�����ʞ�����5��M�="a8��딅��|rUa���bg,2:��vU&ڙ���w�5�mS��Qz��mǚ7�E��+���5�Q'��՛<�ӕǙgNr�4�!�M�̩���>�k��~�Vx+�ڦ@�����2wC9�wΑ�P�gj��R�4L�5'���eY}�l��է�ΦPg�w7��K��K�R��R�:���zZ{Y���{�pf�p�n�}ٵ���4�����l�EȆ;GBv2���b�-�����퐽�q���;.�{!��x�����f��t@#v��x��MN��rxEr.7g��q1P�MdK��^�!��P�@ճ0�KKv�&�I"���Z��f_Իy՝�X�wNm���On
�Wx �2N{����0����8w�[&棺��s���^�y�v�I������R$R�N��<;��BV����2�
�*l���774�ՖiL���J�@��(��A�X�١×t�`�)�l$������w_�Y:>����� ����ۤ���*֖dڌ'����[�g�q�W�2V!�Cʽ�[�DDε�H�׬��+���ڶ�kݻBoDs��ӱz$�ތ�f/{3}/�4���[ћV��uJ���{^�5x�q��r��p�����g+1�5V�>j��s��`�M�S�sQAs�c��5x�]���A���!�T�c��m�S���F�j_�Ƭ9�y��^�p�0��|������-�=˚�[�v��k��f���d�bS���3��i����Nl;���u��3m��k�A�,�Y)�}NFnʟV�)�w䍪s�7(d9�סD�v�7���]�{e~9r�_�_HWO�<�<S2S�N�v�97a��`�=���wb����耞���K��_g+[�)�wb���;��ǭX��^jq��G�?w�����eG칕ie��H�P���%I����׾������$��{<��3k�!��+H�Tk|�#���ږ��9|5N����;���Y4m���H�f��#Kvov���t�.�#tVo�e_�Ū�zL �!��0�r˻_�;H�]�qP^�	�c�Χ�x
�/lV��5vū;+����h+����|dEE��{�+��ȀU)��^r������G7
��L���t�����x�Q�9x���*�E��GJ��R �N��z��<qu�)�q�;o�筅����{��<S_�;&GSݥN�'��e��I�
v
Əm��6�f�Cm���%���������%�Nz�����d[�N��d�}Z��]��kNǎ�e���̟z.�z��w�ם���ϲ�w݆��zK:(֑͕"SU������Z�mz{5������ܽϫ��Ȯ�r�{�b��O��-�v1l^�룷��M�0�@��Z����q��3��'�\H�»D,�6�Xx6of���'�}�؃��^EYq��ݠ��9e����>��8��d�^wi;0����A/���s	��S�f�z�[Tr���ކ��]f��g;���L�\�Y�;e�vy5����~�����۲�Z��ܱmi��{I;x����W9��]�ǆAᰪ%g�3r�<�i�-.��jnv���J�c�5ӭK�������<���:�sm�.�{��[M�z������U;�݆h&/7'+T�t�N:J�0Jo�n��:��CɊ�[c�F�gr�9�2����ʗ�3��� v�.['��L'��w�<��{o;��������'����w�O�k�wp9<��ݦ��K�}�늘�����$�k�K=�ֻ�o�Y��g��=^}�׽�}�B����Cnۍ�Y9{��'L�6���yZ���X�hL�g�<�j���2�Y����(���,��=����ѻo�����ͥ�|����s�������������|g��A���-�����m��k�E�Ȇ;m��[���(�F�깷��+��.��o5㵮h�P8�`����-W?S̶D�iiג�~��O|�<E���{����Vkk�v�U�}bp�/Ȝ1�'�t��E;�f����[_b��E9����6���[�Sh_�=d��Rۧ�-?*�^ԗ��R���׭�?S�8��b���<n@����s.�=���F[�>�e�:Xz,l�>=Ӌ��SOU��:���n�\���R�*� �廣4?��(0"V[䟦�^a����;�m��=O���CSM�%U�dKù14MfZo�j�F2��7ɷsz76�t�1����y��v\����~]᣷���n�_9n�U�V_���n�fL���]�Z���1՗.޾����u3�����}���]�)^M]9���Vm*���O0ʱ��f��n�
i�9�8T��ߺ}u�'?a��n�D��Zqylɯfy����g��^�l�
ᜉ����8�u���E>W7+D�_L�ͳ5��'j87��ù�
����ˆux�	9�#����%�J+70��uf����.$ryf�,^>r`tgW�׽�~7�s�h=��M���.-k���Uro8��Dx�O�,���R{Y�=^���;b�`�O�. �b��~=kw��u芭.���+TFk���;/%�D�x4�{BOk��"��
��<�e�č^봷��7��q��οV3�����%�[���Յ.O�_żwܿo�;�6����н�J+5T�2��h����/"��8f<��m5G|���ږ�gx�I-�+6	 W2v_�w����X�Kԕ�2��'�©�A�q�z|��yk�	p�Fk�����4H�/{V���e�s	��GP8���e¶����~��{�P{���_��
�0����=M�>ǋh:��t]��^�;�-�ػm�Dp�0=�z���m��>���w����	s������w�����H ��F{z䔏��@O�B}�b���Ƴ�����"�`�n�/}��m��u <�f���М�K��0�I�Pn*g�g.ep��{%��֢dxEgY��܍7��g!l��|ۦ7#��ô%�c�srPA�-�}FQ|r.����IU��]L�ux���x��õ����2�lW��cOJHT;�������|B洣�X֪��a��U֑�sk�TwJ�o;��Uq���n#�H�H
}����Vv���3��^=j{<dt�#P[��:�K��G����q���:��s]%�z-Kי����.��^�[�O~� p��R*O{&�����[�"��D�G�7�;��9����:k}>��y�]�w/dܹ�Z"Ldomz����q��^�5)�;�'\᩾Y*��y�+<p��w�}]'۠��dYD����N�0<P�i�2��
ݟV���g*�\�1���r�*�*:�/�����G��'��K�������,03�*�N�&Ԭў�n�AQ���$�_i�iV�@0{��F�'�m<!]���=������X�k�8���Gæ��F\
��Ι������P~�^a���pzͦ��Ht�w��u�G�R��e^�BOW�=T��������G�(��9\�t���_��T�JMG�U_{+M�{��=꺎�枘�q>���Up��?]��o���?9''/�Q
<|T��_��}���33���(ul��_�1�n��T��r��;�x�Tr�\v��8{����z3������{�3kV�pg��'��<��\���Q;��J����pv����xx�?S��V�4���M@9�g��>%n)����UG]z��������Q�@L$�q��\�>�ѹN2���UY[܅��vп�^܅��%���6�;0�(�#Qp>'���/m�=��ч�4]�M�J|zl�B�B[9MS%�и�U�^vS�s(	�b�wS)LL��z���w\
�7[5��ߵ[���x;zg���;d�ێ�qۅ׸�i���TA`�0d�v�"�n逶�ѕ���=^َ��r��a��y�ß����)>*��W����di�7�@N�=n�O�LQ�z	����8�B�%��g��mR��� �A��Ǜ�v��]9����/��Nݥ�K���,�-g^��2:"��D����ݽ��z�L�g��{.�Í�=���@��g$����8�d���K�����䫱�.�gM������#پ���DZob��ck?��d
9:��|ws���s�7�w��uD���QSժzb����^��-P}Ǝa� !0{� ���Y��Bܩr}��q�&��A"D ��~���~Ԡ�wU�E\�Qsp��<�|{jEJ��Ցa��u	m��Uv�z�]r��ʱ��MoX7�k�A�' ���|ĺ����r�X�_k����q�X}�N�j������E$� �ϸ�y������&K�=�:��oP�+�`�7���f�K������јvgn��ޖ�X����5������rb�~��&�����t=|����YS&���͡;>���͜���j��y��a�T���ҟ3��Ǫ#�V����##˨t��t�����yV<�y�Qu�:��Qך��L��6�t0ץ;~�)�`91�~�	K����%]�9oM�+Q��R��]eI�~V�|����w�"�f�B���;og�ұ� ��k�"���9&g���7!i����w�֪="�_�_��jݟ�E��c۟~�lX�:�{����ߋ��Qs2�*'�Y��\H�M�6����b�����1�IWP�H�<��T~��i(�=�T�)ݏ��Ef�aƽ�Qե��ն�Q�#J+n�щ��4���j5��ۨ������| �dw�H��p�y��h4g���dɒ��;���og��[j^ʉ,�׼ Η��u6����zj3�����Ȟ���C{�_�]l�2>y�,����N��3�c�_`y�h^�O���:%���p�OF�Ү=�a{�x�o���]���#�_��]��.��]y0��.U[�묽Kܰ��T�p��]ӟY����,R�.�Vv��Σ��.��<�O��yhv�	O�31z)����:I;�e�1 �S=��P]�]XL�}X69��w>��n;Ԅ���Q���Qqyi����>���~�u��P&�Q��u2��*'+��z)j��������`�e��[�>�����OFq��o��Z��*���M�sq$#0_�@�|f�A��eC��eu�����ťe�ũ{�{�3�/��v�������E̒�����8H
Cډ��Og�8�f,p��>��kw���`��B�'�<_L��yƼ>��B�]WI��UD5�	������yv�ؕӒޝٞ�6������9�:շra'�x����G��}B��<��J�YI\�{D����j�2�Ȏ��_�����zX�G��p�J�E�t:f��zD��}Q�Y6��:V������!Sӣ�ͮMM�q nT(<��9��Χpp �s��X�\��W݂��k+���Ӽ����*̖�ɯ�7u�z�����Ր�4S��9�=�e���\�p<r����.����︇��D��-�X'$ŝ�30�q��"�6�  G^�fM���7�ٙs'U�l	�0�������۲���%�z|�G�����{��������7�=;/�G�;��I_��K��.2�c�Jv�a�ϰ�8�m1�rc�-�쾻���Mf��^=U�r=�\%gm������9���뎪(���;���+���{�.��꾎���k�`r����� l�^��U�W��w��g�9�;�,dx��fQ��awD��G(η�3R���;���~,	�ۃQ;׬�ϥ;|rz뇷��/�^ܢ��-��]3r��ʾ˳����t@3���M#WH��C��@��"e�>�=6�u�c.�&�w�{���^�(���X1Zz�b�y� '~�+�uX����Ƴ����V���3���=h� ��z�y}G��K$��0�LU��-���	�����x-D��(tпm��׽Yw��jw��WG*!��*czr�r�3���@��#��-��2���*r'�{P�3��=b�o��=��^������\�_�ul��>�8!H�?T�!����XU�rN`5+>��TX�_�:�N��6^���t��-�9v6��4[isdY�Y]�L�VA|�Eܵ��3TFj���t@Y7x��Y�s�l�v"3a��i�,�½-�8z�랸��F�ۻ�V,o+��0�.��4���_�nTb$ct�x��f��&
����t����d��K�=7��X.c���W�Ԩ�{=���y�e�}�aOuy�N7<��E1��s�n�#,����R�s}e�0�(�j��.u�e�4�Im�B����W�nb�U�j�*)2�� �D*���`ŏ����H�tR���ڎ0���ktg�8���D.&��t�DCCw�e�eu�ek��V���5��z9��N벉<\Q�'[���):�U�5z:��Д��n]��2�.���H�٨r{����aGqz^��C�g}�q��f������zb�ϲ�ܴ"��F�F8��Eu�Ym��Р�Qa\���vic�B,�Ń��*IN,��j�c�|U�1���[� �t�
�3JYMj+���Q#!G��=��-�{ܔ��w�>ã.��b�<M�L�p`��i	��`m�Lb�V�ކR��7�v)�qfw`^-�A-}�*,���h.
�������;��5,]P�SJB�]�(�Sx�[�k�P�����#>Ɓ�����ܬd;m�� B� ��B�X�8������q�O�l��w����w�>�����g
�0�܎w����h��b�	��j�#�J��ԟRs6��t���V�U�x�7H}e�7���0U͓����0�e⼡�8��f��I仧@�i:Q8�
7"�ɓZ0Ϛ_#�A���gx����]�+�7v:|�]��h��wYI��o���Fq��]��Ӊ����,���6�����H�	�ܧ8�b���r��51���G�^b��3��y�CI��'�˹�m��{��6��,� �(j�V̷u9<������E�"gm���{����'�X&
�o��I�j�l��>pޝ�^޾�z}�!-�FM����?/g<ۮllp1��$����w8��z���wX����Q)-r�	�2�����q�.��ɩ�Av�k�Q���V҇�7n�b�7ײ�����s�ۊ9E�~�o�f8��j�0h���k;A�-��#;�-ɗ�f�jI*4��[��#:�g�����i�aGV�+���;\Z��C�X���+���H��$��%�hu�-ЁM��'ֶ� �7�e��.��ǜˎ��J�wt��)�}w��:bXn,9��;<��iBX��/o{�$����nP��:FB�6ۮ����6����0g:i[-�yb��fE��&��Ί2ʀY\h�]�[�� �Qa:-7�;�ï�9v,Y��t��G�e8��*��L�b�e� ��|	 ����uAQh�"��uK]ܜ���Et��YТ��Tk�T�)6UQ�L��9�J�\΅µ"�l�4S�y!y,�*/R
qB�aA�PQUep�=H��9ʊs�i�VADG"���B��PG("+R������4H����QQAEª�W* ����͗(*�e�Z���jQ5*����^��vr�(���e���¢.\����"9¹r�(",�iDEG,ʯP���*�Dz@���R�P�\9F�TEΘC��TDG(�wn�(�PQW*3.Q\��(��Ey�!S�(��E\���fQ�TDR�2�J�28DI%JJ(�����h���
�ZH\�D�ʪ**.�6��TPL�
Jа��*�:�ԎQU$]u��(�5��*df|�y�\�	x"AB����%����+հ�آ�=����7�5č�������齹���^�]3��g��Cs�*����ֽ{����0f��������=�q�ps�IQ}��{�����o���K<���(��1
CA�u���J�� �2*s�٨��]h!�yY�����q�/�:�v'O�mZo�C���3��=�D7����sYX�l�Ǣ5o\��Q<��<�X��{�y����Ҝ��Ϳ6�th
����$�$�t�诋������T?u��J�I���\NЪx=3��*ǳ�T��2���hz�z2�Ts�雪^Pܮ���z�
����>Ú�+��'����ۺ����p��ޜ�>�:M�gu v�]_ܨỎU�2��ӕ�����J�=����q���=���n��d��Z5꺇iM=1�]�s�uW	Y��C~��c�$���7��2D~̚��O,�[���Ox���>��<�m�*��
]^������ܯ��\�{�eL�o�ҫ؟o��{���5* O�bpϏ��<
��=��Q;��D�~��6;�>4���ɽB�go���?\�ȇ��^�MG�AS��n������t�N����B��Y�B�k+�;�h�jPr�н��,�L<ӄE���9H��x�xl��/,@���Ǧ&�L�Z�{��vc�A���^�j���?��̝��2�.����e]G�^.�n{K����F��h��<W,�v2W[&ޕd�h�WXp�+����G��?���Em���ަGkې��$���5v���n�������lBn��gW�1bJ��|�*Q���*��K��~j�K��	.�e01T;��J`�[{�u����nn�����f|vֻ�Cީ������;��hs�{��,�ƨ��@)����|�ntӼM^�s&:�u��6�v�s޶��I�W�r�>��|c�4��������>�;�P����+�ٛ3��u`b�tա�}ֆ�;�i=fG]x�z�������٢��9� !%������6/^Q{{���}[ǭWpQ����=��C�X�5E���wV�n��U˪.o��<���mH�R���L>5�wQQ�F뢶�o��OzOC�p�&k�W��|�K��*d�:M���9�_��91�����9*���e���Ч7T�G����iOq2m�P�׀��G9��}���f�-�ᬇ��~k#�겹���:�ׅ\z_�z�����rb���7�= ����z�Q�}�*d��H���b���Pr�sݫ�L��jM��8Y1�x-~T-����n`A���`��/I�f��w[�LT���k�
g2����j9�o6ǡ�V���E��uc�	H���]��4a�ڛB�ۣ�"�������9^t�m�7w���nl�F�9�Rw�>�,z�Ua�J�r3�.��7�7�w;�+K���ORqؙ�Z�7���7rbW�\�tc1�M��T�a>�S+�V�*����ҬW�z/:k�{%{ٵ�}~������86�����I��0l�ɇ�YU�qEq*����<<�_τ�e��Wڨ��-HQ��J���WiK��.ܯI�N����^񿌪�)�xe3���Tc6�U���!�s��^��ny��0B�{�.#"]p|rz�3��!C�[%y%��pd���+ݒ�I��)H������j�~�Lo1�P%y��p�S�]���#}����$�IT�Wq�]�������8p]N։�ӝ�2�TP��.�Vv��Σ����0�ytL�5�3��1'k��y�{��D�
 E�%��AvEՄ˧Ճy��w;h�ձm���G�-�]��ޙ6���%��j�4����0�3
���=-���A�Ȼ�T�nh����sx���vb�}]~+���o��=qwlU�uQ�r Nn$�g��T���O���.�PN�b�}�ئ��7�����ݗ�a�����e�(�}#����zi��ԓe;�=�5R�{z��4S��8<[��#�&�ӨМ"��e��A��c���׹uO�MǇ�.�F��h݉�DQ��s��#;N�u�^�Ur�=��_��6��"��<��tg������g�ӵ�m�Yqu|j�]Q,_��9�$0�Nk�靦�cw!����O�o#يlWѬ�ꄶ�,�D�}3�%�q�O�8�.g��UQw{ދ�S����=�r�S�j���*<V���z{�{d�Z��LZO���z�@u��(��4u��;z)I��UIcQ��I>�#��hD��_�WOx��X�D{��R��x�����7���VUg.'g�S���2k|�Ѻm���.d����>�c����!���i�
�û�x{�sA�Wd�:�n{�>W�1���ceW��'�x�������u����*���}����;�ݰ��<��{�ƺ>��O����+��{�+$�) �Ύ�(��ʯڨQ����V�o9Tx7�������x�M�gY~���9�U�W�j�����Ȏ{GN�K�2���{f��W�ڛ���*J��}[!���Ł�jN��02%;|rz뇷��(�{r�p���T�.�r�a��JC�*�6k��
(NGb��U�hr�c޸�N���Eu`�:9���T�������}b(d��X��V�=�ژ$��;��zee!2�M�$��W�^޼ٽL]�in��Q`!��0�����{DwI{��W`�p�ρtR�U��e Z��M�Z�1��u2�ota��$��b U����u���Q�����@������Ivf-2����y� '�!�4/3O�to�6\�q#|i���������"�����R4��7��,P���F[7S<4J@��1�����;s�Y��s����?*czr�r�8K��@��JF*�C��5ܶ=�yL�*%^��u��=w>
����nw�Gܤ�����#��V��3�x�c��@U>�Ȩ(2��fvPݼ�Jo:@=�LM��f���N�1���}��wJ�n#;��]��+��dzܹ���K���`G9�@R�dTN�o�¼��.�g�/�}��wu����1]_�T����{��EtJ��%̐��D����욾�:��C��E�ԉ��;�LC�>���{��h���]o ܼ��r���p�诋���������rž��Sy��hj��[��%b����4�3#=�p+�gLܹ�yN�q�m{�C��5�!GKnn|�C��7z���WQ�K��瓠:M�u u�H�}ʎ��^�(�NW�gGG8̡;Q�J�`r7�i�k�!Ak���]���8������������ۢ�v�(d]
{7,[�h�����Wj�,�ZS��LU�Ŷ��o1�dQ�*�a=e���+od�Q�����6���=�s�u��n�B.�s��%�l�{�_�~�[����=�N׻�~b�ytV��uW	Y�]������?9''.:�����5�g�J���O=���tm9�>��Ks�ዕO�>K�x�����}iB�?#Ohx5������i��жt��sPr��x\VMx�<
��01΂���;/:D�r4�gvUS��{�3�~���76z9*��{r�<����aL5�n������� e}~�$��S@��.ٻ�Jl�ឯW2߫�������~�	<�If��4gjўFC��^}�*fn�ً�ڽ�A,�9�e)�^����yHo����;)�K��@H�P��=]02���r����$��{s������g��x.�OG#�O��w��q���������j� �1Z�ߡ]%�-r8��.�Zs�l'n�p�Ȏ{���ܤ����p}p��t���|p���Y"q�S�[�y�=�D����`� i\g���ά_��C>s�7�w�ԓ�v,oE�)����dޯ$��=w늸�,�c������@Q�zf������C{� ~����pUT'/�{��+�����
�l���U%��Ieb�$��E]o�4�|w2��e]�h+k�f��!n��������JR[׃X��w���T�e�b�vw4��|λ�6w)�M���K2y�IʫS��'��Agn��h��[f}�����8���z9�h�U�E\K�.o��<�A!�2.%K��ϠL>5��oq���<�0�W��M��Ѿ��7�ԁ��^c5�*;���f=*��9M���Uc�%���k��<�U���K7G�~5�&F���iK�d��7�:��BȨ�X:M¹<V�|ϝ.����3s+���;+��>���W�~5��w޻��WI��yԌ�r��<7����G�z�GPoq(���ܨ�:����<}���ǽ3A����##˨t���7�v�_@��:No���y��8z{�y���&d法�������9�>��Lpx��E��?U��02����v��&�#�V~c.d�\�^���^�`7�z�_Օ^7�6�P��}���ue��J�t;�ʭ�2'������]�{���'߶�#���ͯ��W:���xWp�I������{wYy�z4�~�>K�q���=u��h(n|��K,��3}R�?r�F꽕�K'g3Z�u�3�1V�joƙW�P%y��p�S�]�� ��7�/L�{^��n.�Mq������<7XW>o�X�l��ݱ����Gv�b�𔫮��ܵOY	����P�A����[*7$~K���7�C9�o��W�U�>��(%st����7��&]�\�q�ZE��I�*��_��R�?tP{)´#T�p�&̨y,������g�T����"̄��2�tv����;|l�S����\⋏Eu��n���Q�p��O_�P12�[2J���f�v��29��v]3��ȕ�5o3}�����n������f�Qfߤ�N�?����n�Pzj�'�Ǽr��}���u��II9�;�>�g}���9�$gUS���M�9 '7����~�6_�G�k���fV��Ե�8��ӷ�[#�kj��{�'4�.:v�������^�TK�;��s�@M`px��O�h^e�Jk��3�҅d����Ko��3Ȟ93�%���>��B��U�o�y���W[����ԠO��&�T�f��]+Ƽ_�l��mT�I�{���G�}W�c�2��g�MJ��Y������7.���M���_���k��V�T�NGL���.��A��윷~n7��q^7�e@��˙5�(�Yv�u�׼n���ͦ<*>�]0�^�DP���i�Y��hQ��自�3y�c�g>�q�z��zfU������	�~�3�q��׫5����w���;ۈ�{WY���12{Q昣gLd���n�&]8j��Ώy���m�W��1!J��}�g6��B�p����p&:���;�֮$�VM����ͦv��IC��<�}���,�dZM���\����g��罺����R��x|��7�G��������������Dt�G�����*���Y��Ǘ�ڿv��w���x��=�w���d���9�U�W��L<�ɟ�t��i��-u�U��8	�<����G)��=���N��03��߂��w���~<�~4z~.��5���D�����@ߔ?�����'�'��?�����C+}49_�w J�]�9N���+��q�YR��}���9$+�=�;^�ߪQQ%�X1H�LI<���	ߪB
��cۖVƅb쮴:oJ�ɽԧ��3K҂ފ�c�ϥ��y��Y�,�јP$�wF[7S</���!���U|�M�AU����X��n���-O��M��7�+�(�8K�t NH@`�Pa���.���{��y�x�ܠ��^-�qz\r��;�r=}ul��3�x�8����z��2UVN�v_ck8	�P*�sp��c�Ӵ�dC�m��}�+I��;���w|h_DN�Rz9��s���=�D���#�D��Y�,*�=D:K�3�<��Ϻg�L�����+�����kX���6ȫ}��W��^l�RT�tV!�����+zki�q�3��0+�}[�P�h߶[1�` �*S�����i1:6/u1y[r�gΗ�e����ݣ*3�{r��_x�<�{  �W�	���{�,�une��SX"t����s��~�W����5=4��2G-�H$����울�c��C�[�!8�_q��\}xk,<�u;�M��5�q�)��A�y}&�M���^ר���釆�SY�����ʿ]��Ɣ׹�ݚ�э�7��i������w�)K�����T��^a���$�^C�����~���1�ON��]W�ǗP';��}t=qʎ��U�2���ps�%t�+G����g��l>������p��3_G���S]�2<�+x�{��J��롷��g��q͏x��U鬫�)g�O���!TO�]N3�Y�9���3���}*��%׼r7���PI����_m����^|=����4b̩��!t�;�f��'����zX�u�����_���F��t���G��_���MW��k۔rO�{�5�*��W�����N�]���/$����ٷr�jTyZ��WW3��׃�y���/T�p�%��h�ڇ �%?��k~���KKu�G�3��@/t�3���Ȋj�E�!�g�[��`��&P>F;ҋ����֞v�B�3)e)J�ĤŨ پ��f��vmust"]��ڏe�p��(���*�M|qq;P��"���p=V�K|:�eƠ:�X�lb�{E컜V�^Sh&'L==�+KjJ��x�}�;c���޻�!N�\���oo+d��HV��m���u����ǣ����^��/;$���ׅ�Nœ߳)���h�Bk���,#Otxr��Ҩ�E��i��l]��3�w�<%��B�[�Ɗ;[�p���7s�	V.��`-b�{�<T�p+���u�V۾�*�N�j�K�y�{	x]`��@�u�50�CɩS1��]6�A�Etlk�S:�|�gو�S�ZO��w��<l°��Y�����>|NR9@��\�v<��H�x��9/O\3�R�6#�c6�(��ih�նk�z*
΅�q���guQt�s 
����ܘ_�a����p�嘇}�*F[)�w� 殴�E�@�"�Nqy��������jot���ũ�L�cO#)��yx� ቛ�6��۔�8pC>r�%Z�r���(��E�"Ln�U}���*k�VUE�9\{J��¤OQ��*w!x+Nl��m��j�ekۀ���Ι��;:�O�§a�S������U{�p��GXn;��2}�)������%Ky�߈�n�V��9�m�,��"��|�=��N���]fE�t��n�h�' �O)��켍ig�3����'��co�t{�y!�k��=��f�Z�v�u�$����a�T��(qmTxf���x��uЂ�*���"����#L�N�*"	����^!CVg��̈́�.��^�W8N�9#D�;��w�͚�h�T,N0S�a�ð��]�.�u"QN�w�hv�-��F�D֥�Ӱ,+b���M:��&,�L�yI �NAj��CC���xS�V�.�������)�_-�+��R^�� N�E2�C	h����U�6ie��M��ػ��l�/xf��nf����=��]�bsY\'�ǭ��&L8���sy{@�wqm�)g y�!�gO%�{�}�3%�kh[I�e�.����w:��+iТ��,���,,"��5��mY�wGZw��E����V{�K�x*��0�p��y�����T/u�u�����ʲ��� �_��d�Uʎ_{I��y��|ӈ�
y��o(���p|�ӱo��C�ނ��f���2Wu��1pK.�x��/VE;�wy4�}5�|�Z��©��6����ۋ��>a���
w�̥f۸ju�M�u/�� Kɂ�2v��v��@:����B�{°~հ��o+z@s[��Z%��Y�9wѣ�JaCs��s3��#f���Gr���m�mU���5��4�ⷛ�a�{}�ՠ�{�^��ve���{�*p��7,|E���G���eC��H;�x8��A�0Gn5�_c�\��:��7)3��6���A>��$��A>
��j���\���ra�DW,���rdzH갈��8,��K�U\;��!DE^��EE�Ȃ�)̊���B���G"*U�(�:�Ȋ���.h&t���� �P�"9TUE��	\��tU��s�$\I*Т�\*
�Va����#Ie�"���Ur"
dD<�ܮC9�����AUp���˺%U̔�ʊ�H�r".TU�(�R)�H��L
�D��Y^����QAQ�QAʠ�*�Qr*�(*�DL�R�r�$�( �r�*(��t�UZ%Q[��L��0�")͔DE�� ���Ԋ�A99W"�][ǐ�g�Ȼ��!9�Tr���DUO"�=+���+�A>$����(� I����=0��
§-�7���z��'e�$w�ln�X�y�u�Iz����ߔ鯻G���g�y��񠊄��b����j��п}S9��U*�9fQwz�\=�.�Dv��Σ�����3�Y�(�愧�
�1��'=�� �|e�x�cb*e.���a;�o8xg=�h�'�����9dL���Y�s������jH�1���(�8���_�eq�	���)[Z9�Z9�Oc:�]�\uݭ�z3�'S���w�q�G��99������4�J��%�8��zto��~��h�c�����|0��>�;��uE�3D� +��R*%K�����7ђ^�;S�{��ã���]���}H�88_3^����n"]_L�Ī�ԁ#|���V{�(ɞ���-%�?K�ۑ���}b��t'����0}��^��Y��I̛���+�(�<6���J�ӝ��ON��K��[�~5꺇q޻���t����9�wj m�{]~u�M�jPD�̩�Q�*y���zz3�68�DI�~n~��GL�$>٨⟽�.�/��{�3������^��>���D��>�9<��OF�O�F��d}8�Q2�{�Cs���BZ�Hmң��ǝ�T9�����l/��6��u?g����c|Fi=�oB,�������T��a'w;��&���V��Tꩩ;�����f�<��3�[��3f廰�wM���o��O���Ak��>]J	��}7s�YU�ԍ�};�=�4:T�l���ˑ~�ZN�t�5����Ux�ħ��8����Z�Y��&��Я�E˪�FD�c�r#�+��.W�qە�;��i:7:��6eT<��*:�m�[���y��Q�����^��\FD����O]F{!��/箶J�K,�#��^+�63 �V+��Z��+�L����R������Ƹ���猋������בE��5,z��g���v��>2�B�D�3aW��<.�RU<��	\G����.�R��|Ͻ�WD�]Wu�]��kz9�i�7��=fP"��L�o�AvEՄͻ}~ֹ��}>��`���σ��%wz�����O���L����/� ����2��"�R�\k��7�O�1�R�{k;ΟW#�}Dy��=}wlWt���� ��f�@�cN����>��Q�-�k�L���=�ʎSԑNg�y�Dt�x}�F�u���]Q,\s�<��ĽH�Μ3譬}櫀��n�j&s�X��a����r�"x�tϸ��k�Wϫ8����`F;�Wx}�R���*l�9O�c�w���}@ػ�6[0�J��~<�d=:�9=�n���A36�����^ʃ{���f�̾�Ҷ)��*���n���{gh�D��5gŤUW�'�����-�p\ӯ�{�q��74 ��]�[�u�:u-�I�ڢ�Ch9�h]9^5~�ƣ�$:շra'�x��g�o�Z����7�*�t�:69� WvR�T�h��=V����c֛���Y��N\���,�VZ��_O�����%Rxl�Gzty�W��FTwS'9��������qE����LxQ~��i���z��b�_1�4���P�7�V:v{��o1��93+~�8%���r{
���eK���5���=,�=��^��
�xR��{�U�Vv����7�tA���QG�/��ɷ��}kܷ9���2;����1�P�>dN�w��ѽx*;�y3�]/�ץ�qڏ��rz���%~<|u?P���m�H�7���{pjw�Y����9=u��cзoT׫��zz����N�j��F;�׷<]�%�5��e^�F��!�~���;�%y�ȗ!Fu�v{�W�9wۨ�-�譬	a��1��R�y,��Ţ
�2�yd�=R^�*-��d�ۑ�omm�7�s�e3K҃ޮ�9�~�i�n;��]�f�a�-���ێ�5���ˋa@*I��tz��y<Y^�*�k���o���c|g�Q�7�n�\2�H:���
ek:ɜ���\�K��!�-��
�� �(^[�<ѹ��LlV�<������s.�>�N ���m�M�k���!�9An�5'f��C��w�?g�L�k�E��*cr{�ò4ωw��	��@T���k�מ9J�r�_A�
}�Q�<�]��۵�����I�]��ul��3�x�/=Z���O�K�^�@G	;� 9�@�717�)�����c�o����ZM�u�����;������qFbp2q��r�C��TQ�������ds�i@,*�Q��As����g��;6�r;j�v����Zu��j��2��J�!� h��"�J�M_���W��c��ا�}=G/xfۺZ�':G}Ι=��x�u�_d�O�T�<��kC>׌�}��׾�<<�����&�aN-R���̭�Uɸ�]\�Gu�{�ދ��Y�7.lS�vlv���g��.����{?v�?�9��i�0�;#��zs��&�3��;o����7qʽ&Q�y���?E�Oe�z�(;�/�t�wJ�='�Nx�5꺆���]�=��+#�롽��@e�����~��w�\ͥ�@�2ǼI��uD*�u9�E�9�>��Ks�ዕO�!.��dK�M��~���8 X�O_c��EI�_j����S7��<���l]�tkѣ�ٸ���78����2���%�ZC���v�K0��ᶲ��G�]���ͪ� �X���A$ARբ+ j�O4����X>ۆ͹s��9.�Z�V�Z�i<�W������L.u?��ܿߣg_�dE�6�ڼ|�3��s���0'�u���;����h�7��4}}���S��j�.U�}�nQϡ����5��ʨw^�F�)���HB��<���Ǳk7<�oHt,�'���2���+���=�.;^܅�)�Y�6�ڇ���Qz+�]�˫\�Wm��9��zey���Y��������/օ���/;)�K����#S���[�y~Ėt���FI:�=T�3�fQv�����x�9�'��:��s�Y���=u����.�y(���l�P:|2P4nbIK�c�6t��{���N�(�_/}�2o��L�A]�ю���,�c�0P� i\g��v�:�1p�B}qO��.g�}QS����Q���]ʖ�}=T�+�wM7�Dw@B`�P��zf���Ϥ{��55Y"�3�#�����/�Ώo���ȫ�T\�s�'��$#'��n�X��٠9{*��
�wY��r����g��T%���7ԁ�5���3^��/���W�1r��S1��q��y�hw߱ �Vkoɋ�)��x\��5��]�I�Q��b�BHT��.��I˱�;��wzܵF�<�d���ywN��=ѕ�ķGc�W9V4j����X��ku�p��]��,,��<�����N�=���������՝,�ʭ�i�]?�����+�Q��x�{�í[w&җ�ɸ}���x��B5��L���q���v���J1��=�GJȁ�b�N��Ot୏K�WP���rb�8��q�= �j�3OS��{ΰ����P��:8@�}�2[��[kG_�+��������UXbҮ܎r#�F��5��]�����Ǧ{�6��u���v�̜�9Q*�a�er7����LpR�!z���c�>�9����t���|�v��;*;g�w��39֓���MA�Qިw�^*z��4E{3#��v�s���� Lgmp��Uk#>�L{�wev����/�ܯI܈N���uW�g.��'Y�ڎ�oM�Zݞ���3qG`4o��^r];�9u��ϧ��=�����[%�[t�٩O���[���5H�(�L��%�S)L\E9M��\Uǝ@�^w<d_��>+�]���A!356h��W{�qq^���v��[/L��<tAw�
�E���RU<��	_���/2�8��Qݨ�i_�M�W��O_6���#4��7�,��e �>��_4�w��r��&�*����i��n���_�X��l0ţkI�R��vp �Q�&nuЀ�x��7�\&9��覝Gu�A��%_�۸}�5X�o:x'�p�T4�7�֟��SZ���k/�\ç�Y%�]�mn��B K��s����
�/�m�����|��F����a�{;�޿��%q��<|��HO������O��?I��0�a~����s;;wc_���H�~z��a苹�P�4#���>�<��wQ���*���M�9 '7B9MM�j~�j�jSy�8t���ӹ�돕u�Y9�����StG����\K�%�������u��$��z=��@c7��@r7j&�Wl�y�	�P��#�9�D�Ι��xݢ9�*�FP�`8��9Y�vg�J�#w���;ƅӕ�W������V�ɋI��*:�[D�/[���j������r��ê=���)���K�#�XLV�q��~_���������:�/�����*|��L�!L���7�;��ދ��2yܑ���(��x�Q~=���)';�ϵ��E���|D��Uׅ�]W����/:�t��t�ێc�|��2����o�>�C��Tl��z�G%w��ݬ��>>��m1r���.�=����+��{{�~��䃇3v�Ϥ|j����q�O=��eW������p&3���|�z{�GuW[�bc�`s����Q��e�K�t����#�a�/�tv�N��	��;���%,��p�T[���&�y��b��rѽ9��KȰG��C�.�ͭ���D���F����:�)������;=Ҫ���S�V���Mݪ�uɻ��gQ����t�����6�s����ON�S��}(u�NQ�r9M��'�{pj'z��=��m*����/�=ɨw��#�[��0�Gk۔]�%�5��Q�>2���ex�厠���=X̚e�7|��>����sr�]X98�os۔rK٘�ARē��9=��%]'ï�y.�=�ݢ�ܚ�5�k>�9OS�K� �4��=ŒX1�U�Ѿ>Bl�W^�^�{#+7w���d�O\�o]�zKS��B�oʘ܉�_�p�n@�.��)O^5�k5-r|T:��g���v�[>���R|U���z���y
��mïq�5�4�o��Or�P;A��"�d����&{;�t��t�#��x������zI�q�ܶd����A�|��ꈤ�@�p$�{
�x���9��
�8���^?J�Zgpg��5��g��}��.덁}Y�q.k��2CP@����TI^ɫ��9S�Vj=C ���>�I��-B�w���q�H��3�oC��W\��Mĩ�y5:*������q6r��<y��اv�w$��s��m�����V�w���@Y%G
�E��"7>q�:o�`��ޕ}ﮇ�C��MY��c(8��8��Pul���8����{�,`g�o}��[!��ҧ�<������ȩ=�v3^�����u�"`����x��1�S�޻�Ԫ��s���O`sC�ї��gL�K�����{����y����F,��y�_~����c�1�7�k���������������G�g���� w8�M�n�Q\�Ϗl�hX6t;�^���|o�q��]C�Jk��G�Eo��Up���5�f"o+w���}>��_�p_��Vi��no�H������Y�qDzX��_ҩ� �;���8�B�o�%.Y6�ֻ'�v�3����v��8s�t��3�|��|}Nx~�������g&z�*��Z������2z��=��{e.U�}�nQvp�펚�xٕP���R=v}=�U����6�
"{wچp����H	u.3�N��~���xns�b���Y�%��6�%�dG�<�Էjr�-��]g8���|O��@L/:�fẄ�r��DK��q�d���+��:�s�j.�j�@vN��P���&zS/�2�{�a��x�=�x��;���#������Z{Z�����H�9�g�鸌j�=fP%@�sS)t��l'n�p�����][ڙ�[+�~��O�?fB]A�}��7����WS�j����4s4,�T�x&c#r��Os�
�{uQ]�cLQ���\z�ui�8+����E�q��2��Z[�{�����y��u�#�dۜr���J��42/ik�x8�鸵��L%�}ɞ���/ٽ6�
J�n4�缼�qe�n���W���Q�c�0P�/��q��ی���J$c�'HS�o�����9�9϶��>���w��t�G]�����<q��G��tu{J7yx�?�x�w?H^�ꮌ���dxTk�h3��y�&��V�q�}�Wꋛ���<������~�NEg��Jg�GK������R[}&ᾤdq���k�w]p%�t�Wy���2�n������2{�hu@�*KG(�<_��~�[w%"��/����׀�O�~R�DM�.@pD~��j'���t�-Â߿<V/a=;^5N~']������N�._��wdݻ�����:�z���D5�2y��-�����x�\S�q܍�=_z��-�]���g�z)e���6�Ύ�����5�}�����X�2q}�*%A��=���n��4��ň�]oE����dH�L\�w�q*{ӑ�C�Oi�����Fw������zY�F!�t���R�Eg%~z��a/% ;;k�S:�ؕL{�wev��+������N��_D!Nh�H��,h����na�g�M�qgсu:I+�|�zz����_;�\s ��Cbf-�*�	O7���-Z�\%� �7K,S|uŃ��+���Xw�8��
h�x%����O��#�/'N������/���Fƍ�H�o=�����#<y,ԭٜ�h�o��ih����ff�V}�#�b��l�qC���M��b��{����7ݺ85��|�<���{�殳Ϥ�Z�CR��!�&�8�P~��yoB�޻�s�
8���wՋ���s+��ںK
w��7�����_݀^�4B�Z��`����[v0�tTn����jﳃt�@E	�_zH�q�TD���o�:Y4v�q�뤸�;�v],S\�eZ��fG������ԄU�3%�A�&�H"�IDk����]K�g{ 8.��_6������Qu��I�[;�z��y�4�!��[Q,z�s=%h:�OK%rF����x+��^^��l>�	��^��-�믤���H=�{H��Z~���K�6�k�ʻ;gF)�R�CN�_);��� �o�-ҵ�!�n�P�}��{r���5N��돹q4^�^�i�!��b*{p�9�W���Sƨ�b�Q�zJr1�L^]�y�H��R�~�B:wcx�1P�:;�c��w8B�a��ٞ�N� �`S9���5��� ��3�sZ�P�;���S/*���B�=X��U�a�C�{�C3���J�A�I�K9v"�נ�@Zz�-����B*��2���	_(>�r�*nSMV�񥣵����u�"�,�Uh��N&�F�wIǋ瓫f�x�q��]L�F\5�rw�$\�|**�8.�d��M�_0ƅ�-��Gq�xb����L�J���r�X>�W�	/���WeO2y����h!ֶ��Q4��
����B+��ۯ�w��gu��0��!BX�V{\#�s�¤�s�y�5肯9;jnM
��"�C[�����w�
ɋ/8�@D�Z.D�Ѧw`���:��B7!2j=~�/AΫ4����F���]i��|�\;O-{�x;�|��:��5���e.��u��Q��w-�5U��g�yX�P�p��B���_r�9�۞��6c3��ߨ�yf�zi��} $��5�J���k,�7�\��΃oj��
�/AA��]ݪW�к8�q�B�]a�E��;E�`g'�&՘ާ�B},�����yY���M/V��Q}s0�wp�%9����%pl�+&��h�D}�������~\	���Xʰз���g}��� M�� N�7���m3���Zwo�)�G{�~��6�^m�`�I��n�ෛrû�Nb�aF�ŭ3-	������0m�:uJ2!Jɯ7�\��4v�Йe������VRj��>�x{3_rwx�#���u���4F�]3|�7\����{;-[H��MJ$0���mW90�c��
v:�n>�)<�y}զB:���*��� !�Q�)flrH���vP\��.U"����rn�!ʢ�U��P]�r��EQU�!:�.Q�"*#�E �2�2(x�A�8S(�Aw�#̈�9�p�*���.W"�$*���ue"eE�|HQ�婑�WL�(��L�(T(��h��r�D�4J�w)��p*��HPr�W<*�#�N��j���H��U��9Ȣ�wE�u
��8Gļ;H.;��TG"���_*FhUr�W�*w�z��PUȈ��\+2/u��`TE\��,��.QQPE�|��)�Px�R��j�T|Br(y[�i�����8E2�eJdG��$����"8\.QuO��/$��8��Ӳ*��HE�s��<���ES�4�����L�B(���r*(*'���^w�R!�1���&z������3�R,�9Q�,��ΗSu"&��L߅���� B��Z�I�9�Ûw��>)�r���aJK`~TA��W^���F���U�@O�u.#"]p|rz�3��О��S��9۷��^���i@=�6;�g����&pe	��yL]9M���0=���"ᾧ�^<�����6OQ�{�U9�!E�ރ��7�^������6@2�*�����,�J��2�G�59�3	�W���6���3�+���;p��v�u�a��,�wK$��@H8�S-���Au��lx\�.����G�-�;�g����#�O3��G���	�����d�y�L�� �PJ�E���=�k�F���g����|=�"�aҥ�����>�<��wQ��b��ON�r3O�.�c���P�ƽ��I�}P#��w���eC�U֑�3�<ϣ�k��>�#z���Mt򪔥��޺v薓��M���n@GzbIO�¸F��	�Im�8�y�>�q-�9i���w��7�I�|���&��TG,�46�9�4."���|v=��=�Ɏ���z�\��2�5��靁�>��_>�d
��WI�UDr�5u�=w���O=o�xΟ�o����vl�����[�fs�ݣUބ(E�%���6�툽��x�`�Z���т	D�D5��'��ش]F�=ec�:�4{��tF����\d\)�bv�K{X��)��a�ʉ��*�0�IO��ĺ��N���X��jơx�e���fy)���|�����t��{ ;�񿷣*G<��_s�#�����;s��:�{�<Ү|��S7�
���]!q	:�9]C��gU����s��S�2�8�	Gy����ޞ�!E�s���Yk���������f�մ�S=��u�s�uW	Y�x6���9��{^qD���u��<��Kﶨ�Q��+*�l.'ư��a�%Mk Ӝ{�X���p�W0:ZP�Ǫ`�Sy3�#{h�܉tG��9G�✎Sq������;լ��X�F�]~���kz��ʖ3ܝ���{r�C��-�tׇ�xNFY��^Mec�u��mES������VkJ�@ך�'+��K�u`�ב���W�%�X1H�L_�3���f��/�'3}�F��4��	��0/��V){�Ʋ;i�S��iR�H<�>���K$���(�۞/Ez�T�3R�������t6r�Po]XײZ�=����LnDOz�vi��yz���abwb�J���	�擄'�Pa��2��r�t�a�nw�Gܤ����#�}�!q��ꊌ�7n䢡���5�ƶr'�ISR�7\���C��r���^�a�t�8���һ�rg�V�t�ֵz�,p���8�m�޹�������Ǎ�Osk)�D�^{y�3�ww!v��]�v�u��,�h�W�"�2��¼oT
�Iha�F��(���B=s )��P* ]10�،�����c�o�㌭�<w���R���ۺ�g&JN���ݳB��TY��;��~2*']oρaTg���jC��+�mZ�Z�%�XEm{��Gw\l��늹s]&��UD5�dl���9�|j[Mt��͉x��1YrF�]��\7ԉ��<�q�*!��A.���SD�8jt{y�|��������'������ڌ>9���W'�Wu�{ 9��ތ�γ�\o3�(3��������M@���������?h,y���k����������@��Cѳ�J\�9�������(����e���W�gG]*��Կ�~+�z���%5�c#ˢ���F�u��k%�{�^��(��	���Co������no����ߍn/�/<	��]��z��M<���Vy"���T��=���u^���\u{�W���޹Ñ�:N�}�Pr�O�b�&�e�,�H��;]7�EZ����k�@ږ�k^@ȕO�9Ӄ�J����9'Ľ����*a�ݱ�r@b� �����؁�X�NE_�Q�4��.r��]���nz��j�G���ؼ<���;���'�nP�Iv+�+4Э���к�0N��W��۷ƭ=�k��Jvr���iCF���{�r�웃�7!p�>����%E\Zo�`LN��I����:��信ի.ߋ޻
��	I��9N��~���s�b���X�%���^r=/E�n�j���M#ʈ.b���n�@\o�<ǝ0��Y����Og"��K��\�K��.٭�sϰ���P��۔�'�e�:IJc~��L�E�޼zg�����m_�Q��}H��ź�oCcg4��3�x�cTAwP��@�<����]9l&��4�M���יKe`��l�뼏G)>*�9\[�1٧�x�8��� i\g�
g{��u�b�"�u����|���N:C���ho��i77�n⻌�;�99�/��ê���9�o�e�(���k�L���}ydp����g'x��:<M���/��"�]Qsq�l�el���wy�'w��[w��ƫ��>U"���g՟	��}��-��m� {���y3^����[q�F�
�ș�dnO.����ڢ܁#}�1WS������j#�&}�n��R��7��ޥ��������U�陭���C�E}��r2�F|zƨ/-Â߿<V/au�:�o�ѣy�����t+GV��Sr�tft|o[L�����LgBn��ZH4-_Vhv��i���orq�rg؜�+�)^�7,������5�N8����z��ӏ�{�p,�Tr��<�y�vB�g3��ED�	�^߫1���9�u݅�(�q��ut��e)�[u5��ڪLv�����Ԍ�&��T��s�֎��^>ϸ�ce�y����][���J꧙��C�X�[]���:f����u�i���G/T���ʉP}�~��F}<�|j~�w�}T��T��s�k���
�X�*����ҧ;g�w{�#3�i;�5&zaVxm�>���Z�[��tWUq�=ī�W ';k�ʪ�FD�c�s��җm`_v��t�"Yp���?g佄���7�e�W��n(�F��py��]K�.x>.z�3���D���$QP��ط�{�t$�d����Y6/·qS<�.�����*���;�2+ܮ%�;�O�s�}��<�}�n\%�����<Wc��3a@(�%JU<��Y�� |_�P�\�]�r���Gf�|+!�;w;�������=ŒyA����qS-�f�Q��Y�Y�EĮŮk�3:�Ǵ���O3��G��w�	��9E��`&����1<��w{�.�kUy�w�ϼn*gGiϮ�*[���|���o;��_�wlU�U���f�Ȯ���R���X��ۙ؇v&Gt�?��b~v<X����q=��%�H+�3���)�����Hp��V�pb�(^�
�<:�����nUެy��Hg:�Ƈ��Z���]W�l_�������ݓ�S����3G%Q�Q�Ňf�y��wN��j��#��@�
y����ys*�H�|�}����;^�u���D��z`V���@l��r�]*��.�-� /|�MD�{<+>���imr*�"x��2�!��א�k5�_k'{�x
�z��.��ܪ��46�9�4."���|w�$3^���5�/;��ց=�c�����Ϻg�odQ�}B��Mʪ#���}~�a���-6g���7>طk]����GF'C�o�x��+�z.`{�\ɨ�G,�c�+�;k�Iͺ�_���w��+�n�6=W\�]#��uX���2=�Ǯ.�W�e[�}�C���T�j����<���ިS����'�����U]㐗P�"=�\%gm��]�4k�쥐fm��s��#v�>>s%�meW���_Fc9T;�SZ�+��F��_z��{ګ.�����kUc��y3���|}�����C�qhw���S��^���m�gR�o�z��U�Қ=�0;��[g'��{_V���(���-�Mxz�G��zi�r[u���?a����'�N�Ȥ�rF�9���>����	���5��kΘQ�g�ڬ�r��L�m��6���O'+ �yA�,�x�7�V�r!�Փ��MS�6�ڽ���|��%@�^{���Uj/?d�2~�a~�M���G��.��Y�N�M99�������k�')�>�讬���1}�nQϞK$�b�K���U_�ko�'/�U]�z�@��Ha\yՊ^f��;_���"^J�$��;��ZM)�ܕ+����ĖtL��.(�#qS<9s(;��IjqC�!�~Tƞ�����s�4O������9�h���P;I]���	�Ĕ�U�9l�Q�_��A��ݯ��x�}�O�A��"
�9���M�P)��uz^q�����d!��@���=��c�Ӵ��܅TKxˌ�\��v�ܥi7��n:��йuE��q s� )�_����[Ƴ�X_Z��Q�\�Mܑ4�5��#z7�|���g�tϸ����θ��s]$��� h�/jE��BUl��N�ú�ꞵs]��H��ծ�\C}H�ϣ����x
���A������4O#�8�����FkM�e��z�u�2�}��vS��W&�:�g��P���]@�L��>�eW\N׷�k&zvlR4�{S[����ߐoN׋���S�m����� �~�^�f����5�X����2��jxOۋ!I-��q�4H�k8y����Y�ҹ�Ƿ��w�%�ڋ��5p٨�;c^�v�H�X�V�H� ���: {:�֧��	�}|���[�l�������Gv:|��	��&����p���v!K���G�7�c���NI�w�s����t���װ�3~/u�Uܟ�5�;!!��޶.���j�<�$�^�ڤ%g�~�Y�Z����~���V�߰/�.o����ܞ[���{����2����(���>��g��r�v�T��t�;�5*�%;O��j�&i~o��jy��G���:#:�Q:����O�9Ӄ�O�*�׷(���/sx�hMһ|��jo�-�q]N����_��}�@$�q�s��讼��ؾ׷!7�dg��;=k�qy+7�#�I�E#�eT+�2����&o���~t���Y����j�Q=��P��Y5qQqY|�@���-u�V<�	.�e01T;��R�����}fQv��ޙ��������������P�Y|ڸz:s�(�>����(	�d�j��/詔�r"̈́�Bsۦ���P�5I�m��N�W'���W��9I�W�r�>��]��>���Ā�(;+��Ƌ���Ȱ����o��=W�a�+C���wR�n;�q:z��W��h�r s� !�'�\�zK�pz3+���ԝ ��t�%�{=��.WU������m-&��w[W���)wn]��V��,4��nY\�MU�ݮ7��9��xئ��?X�ΓQ�7��y�4`�fgE[��=�T�BT什�	�WZ��
&�d�;���8�SY�#޼�Jo?��Ҽf?z���Qܭ�>�����>��/��"��.j�W-s7�ϣ����$q���x\��|_��脶�M�ԁ��^18��<>�~w�*ǜz=9�j��ҜԨ�#ܴ�5���)��q���]}��W�=�����0w��.�'zkVp���ky��_.�d76:O�]+͍�daڭ��w�yON׽��~����QC3��Yܪ�.BOT�Y�*OD>��v��t=|���eL���gGI�8S�q��2:0T�2��w3�/-w�O}����{���t��:o��w\V�w�c�,�]���W����_��,��<Z<������>��0�G�i��N�D%]�;�GN��}��H�s�}�E��FD���w���=O|{*6ⲫ����*�L����J��FJ�=�;��J��~���{���:��Ϛ%<�ڞ�e�v�`a�ՕXo�*�@��@N��ȗP��͟�1�hz�m��û�Y��wn����C/$���2�·$���=��{s΅�+��ߞ	�3�_�{�e��u�����h��!�@�qn+�ՙ��D�x�{cyˈ����u�w�����[j�{����;w~��$���-��)J鸈}l����γ�|��흗�͌�j�1;p�90�4�g����E��σ�ũ<s^K��{��>�7z��?�̏��M�﫲�|]y��zg�v: ��ͅ ��T�Bd�rf��>?��A��[�՗~�Y�-{*(w��=|+;h���Q�sL/����d����&�X�{uw�6��̿-�g���g,���÷����;�v���B|o���ȍ9E�~�?Q��v��dM/n>^�q����o�c��IvL���}�̌�+�~hd�$�mr��3�lNO<������S��H) #�{����0zv3�P��]i�s>���:v�wD��d�]��w�'��j�7�]_��z��-����A )j&�S��Y �9�a���\L�y�L,�ɟX�{zi�e��%�5�*Vq�\�I*d��dy;ƅ�S��W�|k�5=:/���M_y��>�۹1m���:g�og�G��}B��<��r���Ddk�_�Z�-��%�ua�L�{��yٮrǫΰ!F�w"�u����7�����ʁ\��Ms�#�����b�v���毳L)S�z��{��ǅz�����NG�P�7�uX����q�z����irEg��#=�x�X�Dx���1xw~Ė2�L`��MzJk�T#��`'
�̾����ҭ%)��)�H�I��s��f�(;v��T]�Y�4�!�P/�Ny>�(s����(Kl���I�rp�u��{���Xc��\10�ȫ���@ݒ9���ȶ9gI2��5m�o��T�+�+�	k�5,��NM��aW=z�6wv����u&�Ut�b����t�$�W�;#�4+���NIz<}�l�qȮ��7},+#`8v1`�W�O�;jU�wT9ǆ�Z*� �3ػQ��1.߯Mծ�X#"d���[#t�]���uf�52뒔-Vmң��h���۷�$�䂫�e����wzw����wQ�r Q��,V�Rt��ξ��</� ����/�T�M#G-q��r���uB�J�R�B�<��%��J���]b�ʃ���
v�K�� <�D�	c��~M|~�Zڒn�V�i[1��`��<ۍ�0��7p��������5�e�O��9�W;:L����*��{ڍ�+L<�&��F���vٖxI��ѻVl�ᡃ�ћ��m����e+CD]��g.�д^v��~����k�� �
������5)	�l�'�3VHp���j�5b�e��	��4Yҭl�&��uaD<B��:>���kU	��|�W�}���1���g�nT��Dn^�'�y,�|��7^Te ;^�	�s��ON�.��m�A�pu�I-���&��	(s�Y�,�͎��Q��d՝�ť6�ǆ|؉� �Co&׎S��n:�[�[Q����N�ت�*;N�u3s{Q�C9[���su)F�����)a�/6ԧ�1ѷb��4iҮ��){� ޥW����V�Y����`;�4�'� !b�r��'g1���|ѣ���Ҭ=rh���� �\-�t�i�vpl�Y��tw	C�$��ry ��M�t�M��Z�\�d��A��{�d�VZ������my���&-�z���]�A����kb{���V[�o��֎��h�83_ͺ͙}�ھ!�}����5���xo�L��cjۭ7�K9�u1�X(a֣e�z/����\���'�۲����ǜ5�z���J��;�ɡ�-~v;�8��s��k�(v^i��-��6'z�}�
�/�i��,��?	Zn'�>Hr�,�}%%:��c��ã��+L�`e��V��T3ot���π~��ri9�W�bz�n�Ʀ��t��9�+��Le�V��r�p}זd�W��;ђR7!v˫�PjR�W{м+��3q�;�ۛ1�f26mq��o�9�H��p�n��%33���8j�"��=tt�u-0v�y�� n�Q�L�V�Y8Aٔ;��aq�N]��ش޵b|h���E���s](٬>h�]*E첔!N�ܧ�+�!]�h^l<�L��䙅�TTDNdUȜR.��U��_�*�ם�we
�E�u��'���Er
dUDG"Ԣ5
�g�i�κ���A**+�*���"��r�x�sWP�6r�a$QA
�)�J �����D**��q
�dTr��*�(*x�*#�/X�����g*�A_�$��ʣ��R�*�A]:U���E�ܮQQwS�a�$�3�EQL��9�G�.Qs��Zr̨�,�9��O(��:�w�ۢ\���!9Q�� ����G(�EE�.UkB�w�Y���neADr8Q�%Nar(�rr�����D���Ph'�������#����C�j��sP��(���up���J�� ��N��F�;��N�=:f��R���  ���ᢲ�q�%JʳZ��8��\>�,>s�|���������X�v��wVL��b��C{^̗��_��Ƣ=[L\���ϒ�x��xN���M�=�+��ם������.�)^�����2Z;�c�&3���J��@�R,QH����K{'��z��ݵLj���Qޛɟ�t�0-�1p�j��>~C�)��Kw�ZO�\�3�c��{yykZ��	��3���������^1q��r�<��}�^���x\W��ͬ�;�Y�Y����Y���3�tl��{� ^���N���WVY�u�c����Y%٘�t�
eu!7�Q�����-%�m��s�Ґ;�$ ��V)y�|k�X�q]lr9/ԃђY�Y����'���N;ou�I΃0�IΨۊ2ْx&v�Pw����8��M�*cm�P11�h�����vv��;q� �o�(	�ql�(�/�Eܠ�:Xv!��-�{����&v�����qe�7�G�M2���7�B.�d��]17�)��gN��(�²g����t��@����s���V�y�pv�:��йuE��q s����� Od�5R�Q[���Q~��P�V${���A��T\B��3 !�Xb�˶^I7$4LG��Zz3C.�/a:f�Y�%�ǒ��a}��0���c}��r���h��8��Ftr���p�L�4Z�RM:���E\��;��	<,��](��od����P�
�n�x+��G�_Zd9�g�}�>�o��6�Vu�\D���J�!�� hP� x��T:�/�S;�:N�M3�o���Q�z�_��"{"8���ǀ�������L߲�K�sۮ,�+k|�$�%��=��7E3��C�vS�\�Nx]��i�hx�k��:쩶<����khށו�2Y�Z��A������~=F���ת��z�O��:H�1�'�=:�s������v����׃8~1~��~\�^5�'�~/�qז�+.
%��I��^5�y=^1�؟#���+#�롷��g��99q���C���*s��t���p^Su��s�w�f�ɯq�m�1r�� ��;�9�\ur��8��߲"�ٴ����o�{iޝ9��(����x�����=~�t�#'{^@ȕO�9�8;T����^ܢ��/�C��+}w6b��hҥaSI@�TAs�^�F�W���:a'K��S�g����xnG=�u\�L�l�o������"��ZI�I�h��;�3��Qp>'�� n9�e�P�Ϫ0��ezv�W_��][�)7Fuqi�(1G2�/�k�`�9��Dmi�Q@l��q����*���:w����	�jE�ޫa��f���l�_��7nZ=�-T�:W���3bsQBE��l��ɜÛ^\��wœ��^���-{� >5�-i������jB��Gr�w������%�L�& b�rJS���3�e=���xo�G���N��~IN�4}E��>��� ��ϴρf� ���0�lnb����E���j/�6g�X��	̼��]�߳��w����)>*��W���vi�7�$� �b~ 9��ldg:�mv�g��z��U����V�C�u����ZO{�'�c���w<m���
6}W�����m�ג�GD��O��;��^YV�+C!ϫx��8Ώp��@����]o=S�/P<�j��5=��l��A!���TJ��Ղa��	�_%��m��g�kÁ�n|�@d�q�����h��~|�9�T���)ω���
�����èշrL�,�'��~�����,ny���&O}��^|x
ޡdTs�&�]+ lب�;����*�/��W�����6��)<v��+v�o1���t>I]ɋ�}�n;���R3�� .YS&��G,�mh���x�����klȤ3n���-��,gG��1iS܌��3q�|gs����^��������2.�W	���y�����>�Փ\	;e��,�9�)� Tbx�$�#O�̕��.w_f7Wl����uĎ��wl�� zԤicsV��f-������y��C:��F����
)V*�ŵ�.��W,�X�� �)��9m1:��';_�f��e�?}�c�G�i��N�BU�ӛ�C�NGl�����FV����ʪΪ�-�r��-
��fHu73��)�������\��ddD�c�{�{�l]8�J�	� �^f���ز�'�ui:7�s���u������x�
�΀�K�q[͝���{���+z��O��=��q�}%��Ydؼ�L�w3�b��!��⧾����O��U�̷�X�ח(ȵ�O�����]yx�� �l*�e/�Hs�{&Š����Y��\��W���
Q�G�����9�a����7�,��P^�w�=�r֛y���ã�*g�7S:˫	�v��29��w#����R�w_\vF���LX[������V����8@��0�B̒d-��^��{T���6d�[���o��T�0��p�����q����_��TT�9 /�rB3�~�e����P��]iNi�n���ԭ��]�׾���'�Fں�j�]Q,s�<�A )�=���Og�d��g���/�S/c��k��/v���Ll}�#+\9�����N�[G��Lt},��+�pP1Bۺ�𼼌�A�g;̻�昇�Y{��
"�&%��'y�<�3Wi���(.D�h�IyX�w	�8�5l�gi�N�uv]�Y��)����n��7G���`���h�<Nq-q�O�8�.g��%U�	����q�xҎ�#�4}�"��=���<��{$�]�RcЗu�9�=z�C�@Q�+�ܪ�9d	�to!�H�����e��L���DR���҇��:���+���雎��7��N蹀��\��B�3[iũ�[t��78OY�;>��/Ƿ#i�
�]1%�zr<��Κ>������G�W���͛���6��@��'&es3�Q���P�'���/���x�5��b�UWx�������� t�Zy�_���y?~�\?�"�]��QX����,=bngU	O�a�s��P��::=�|*j�Q��Ԑ��d�|���>��z�(��7�>�'��.���A�*r���9��U�s3J㋩����g�^�B��5-^�"S��"z뇷��׌\v�\���|Ky5��Q���EN��T�=�uu�,��3da]頕ǝ���dNS�}/�WVY�u�b��{r�<�I~X���-^>�Ws��SШ�S;�Y<���P��>5�,v��c��~��E�.���.x��^�>�葬Z�Dzg9Hw(H��v��o�"��l�Vl5ytZ	��s�-^�JH�"�I9c�pq=Y@-���/�BS�a��7!l�[���8��0؀��z����j�I2��[�޸u̔ug�\�<<�Vq9:V� MV�J�����O\�N*����fI��߮eo]�{%��C�!�o��O&�B�F�d�¤^{u��a����L���� ��������̂��y������YG���x�x�b]��v|�G)>*�����V��3�x�F8��$���T��&�=�z����2+8?x�"r�s]c:6����]⣺V�y�pv���TY��;��Ƚ΄�(�׊����;]��Vjvz���.��s��'8��덁q՝qW�MĪ����O�����}m�U�H��R+�:�j�e���ڷ�C}(��X|ǀ%_{�=~����duμJ=��zvh�G ��g�}�����ÝrJ�M�'\�w_��ϗ�f�V���R���.�F\
�}X�n\���a��f�h������x���W�3C�;�pjdmѮyUY�nd����� ��wC�ʎ�9&Qޜ�"Ύ�U�늗�|n<W��PWX�~��V^fsj��_=��1�}�s�U�V}����������I�ˏ�D*���w9�蝕��3����k�*�k�|�T��sk{P�rݽ�5���jb߱K:1b�P���9�5
<ғ�Re���2�Us��d�#�k�]�X3.GLs�����D����l�v������	=.xzwE$���Jn��v�rN��=���q^���I�u����{ϸ~�/�t�c�J�샟B]{�#zk��r�v�T��t�;��Pqn���)��ټԵ�晸�(z��A�� gҩ�����l��r���G˶�wτJ��{��g�Jh�f�.��z����ǫ�
�΀I��;N��~���ᵏ�k�?0r��~9J6V,���	=��vS$�q&Ѩ3�A�d8	���x+�:y̳*&��CxK��o�=��[�@�&�|���Z�d���`��D2`r:�!�&~���C]���X�]��9�~��W����g��l�;��;� ��ϴρg�QP��|712��1�4F����4��=���]|0o=�h���y�������>��QP�J�b��K����;Y��/<@��w��ю�1p�C����+�����Ez;���:�9�W�޵N�h���Ob~	f<�$����f����!
��V�9;ǜq�&�uh
�ʮ�R�p�z�����TT�'6Kg ���*^�V|&�	���Iߛ�@��.��Y��杷�����+;�/��`��7���D��R�P�CJ���:}��W����aŊ�l`0����PPN�+s)�8L ��O�w�1{O�-�{�:�$�j�)�{l�!k������B�>=��v��eH�����۠��C���q�5����;�k�s�`�%���_˛>�Ʊ�����8̬>���U�	��>��{3��[ց=rz��d��7�:��,�sc��U��͊�;��O�£_/m�9wO�)Ŭ�w�Oz��ں�Llbq]&������r�dG,����9l��V׸��@���~�J���ԧ��F���UXa)�\lyu��Λ�;����z�rə8�8��u�Vc����,{�P^ެ����9��1½[L.����ѽ4:T�ݳ�e
�9�t�<3ؤL�Ԕސ�֓��������u�^2����v��UV�
�3�HK�P���~�z�z�[��n��_�m�I݄�Iѹ�^�2��W��n���ߋ���:�u�{����ug�)���:'���z�/=�!=u�Pw�Yj&pe@���S��!�������{c�6��{����?w���>+��q� ��7�t�3�;X4�8��^�O�4�{c'7)�u��o��d5�QC�̻�]�x�w;��.��<��,����=����D����^跳�	���}���;ڱM�	f���0���{�=�xP����Z��M��z�M��F�e��2��:��;�?�����\�,�"��M�{�C,xRv�Y�WX����P�C�v42���Uܷ\I�)���@	ڻ���MR��R�{.�$���pI<���7ua3n�_�}�O3��G��z������d�J�wu1pvz�[�j����;3
��Pz[2JN�w0�R�ъ}M}$f��}�B��8��Vg�M�9 +�k��
�����9�!��T��Ͼ�W�#�?Si��jC"}�~��U�$iݝ��;^���#z��ע%���<�	L�J{<+~�q�Y �;kz|oj��s&�1oM�Ѿ��x�D�q�>�^G��8и�U�nUQd	���4�]4�+�~��Vi���BյRcГ�<r#�z�@u��(���+��Ҫ��c��Oh]��sr�+�~ܬJ{Ư����/R������<�q^7�P/�2{Ez�᳃�^�S�`���s�א���f��?1�)LxTz���K���yu3q�V:vv��d���'&������\]���̫�g�Q�u�����9���=~s��5�Ek��JkU�{/��Oxz;j���V=�u�m�: �����O��ʭ7W%��p;�37�Y����~�����&V��G�si^:dP��`4����"{����B@�rt��^M�Z�ـܶ���i_o��t����S�Y0�[γn�۱���|�ސ�[A�S��KM8Wj��96�\��S��b��e���R��W}>���"'���>���o^�������.@�@���ꜣፚ� ��.��T���ӠLgm���]�0
t��������^1v�\��'ķ�tׇ��da��R�T�.[ʍ�s\n�C*�4���vD�:����j���1q�����O^�*�I=��/�{|�w�7�b٣=H]L�o��;��!~갼̾5ޔ;z"���s������$�|'�ѱN�Hv��G�t�',��� Z�r
\�L�\��z��Z��k�<) }��tuѦ��P�!��6�=�Ö��.��9!��-��2��w(>^�8V�eQ�;���=ޟ#��#��y�dz���y�q���Ą]̀���P j鉫�a�ꚋ��ˑs��Ś��u��=���z�0�s����gu�ު�4=����8 sP$�P���8�oM��r�Ԕ�x��U�j
�H��]h �*<\tϸ����6�g\U˚�?}ۊ;ԯ����[%�<d�L�D��vL�.&��:�����>��]|���r,����m�f1����L�����1���c������pcco���6��61���lcm�������1�������6�cch�61��0cco����m��lcm��1�������6��61��vlcm�61����
�2���5�� ���9�>�GP ((Q@} �P�����  ( � 
  � 
AU@�� T��	  HR�
�H

����R* 
�
UQ%EQ�JTI*RU�IB��kR�$DQ��D���RUB$QB��*$��r�
*U)AQ(����@��J��T�)R�)H��
���%"���B��"��P�(IBUR�HT��TE"�5�  ���ܦ9���s���
������t�֥.��'$��+�ks�q�mQ�����Bʰ:ԋ�j��	R�* 
JI�  r�(�V)��ź�^�� Z�Q@Q�EX����(��(��:(�(��-����(��(��B�  X�n(�(��(�b�&�u�wR�UJ�ARJ�QB�m�   �xh�U����v�� nVV��]��]�vT�7-��5-n�m�n��Z�ճWM�p�Wp6Q[��a�n�uR�P�� P����UEx   ���9ۑ�06k[��#���T��\#����Wv�t�9�і:�e��N���l�㫪��I�Nӧn��]��S6�US�ê5v�Z�TUJ���$�R(�
x   O^��zmw\K8ӹk��wt�B�V��:-N��Ӭ��[v�jq�t�
��\u����ہ���ٮ����n۵wk���u�����ݑq%R�**U!(T.��Wx  �޺�,��p�S�u+�n����۱��u��)ۮvۢ�d�못n貺t��:�K����tîݪ��Zs�U�k��`�wV�v�`�:�T4��
�H��  Ysڦ���5sV���Gu�qŮ56gl��Ww]���m�1t˺�u��ۻ�6��JU�b����u���,WJmT�+m»��u�����Rl9JJ	R
TP��R�  ��:g]]�v��"�֔����n�m��w�N�n��v����F�Ui�P�&�23]��i۳�u���J]����r檻�2�-�j���
�AR��"���"K�  '�7���g'rt�J�.�]GW\����5�uݗYm��J�Ukv�U��m�]���v�lC@�M��X5��ں���s����mT�p���R��J�
��   6^<�]��n�E�J�V�k���mvfQҷ:+W`��Q����mmhn�9р��VÓ��[f����S��)P  E=�	)Q@����a4��M0O�J���Q��5Oɤƪ�4� 	4��LUT�R���f���������?��̝�0�Ǹ�s����}�_}�{���	!I��	!I�@$$?hB���IO܄��$d! ����������|�3����+i�^��u�$N�`��Z�W�*��TX+	*"���m"��S^-V�ue��'u���y�l��v{S�oU֬�8��U���H���=
˼���|0T��b������͒�K��m�"4����r�4+�6ҥX����t��u[�c%F�ဧylк�Yi�?�޻]5V+���m'�R�U���.e�f��:d���,J�j��RekY�V�m[��q�A�c8^����DHR���e[9�ʑ<!�ݡ���h���Ô�U��Z$
j����Ù�p1z0����J�]�ڳ��Ð�@�Ւc�.�r,��պ�ڰ&�Z��xٱg"8��BQ'夊l�T
���[$5/t��qGT��5zi�kTo�̓����v溺 �L������􊺓U��7���J�UQwG-\tu<�Z�:���L�;W8uI-�;W�%��\�N�f`�[E^U��;���@ڻw�r"f�i��x��f�[�YB���ݤCC`b�wZ%f`���W㱛l��+ٗ��WZ٫�jV�t����`ٰ[�X�Fмv���q$�[;��1�3^�T�F��M;�Y��v��q���	f��L��Ev=�i ��ާ�<�0bM\7m�vV�;O���^<v�)[ǆc��+�!�r˫9�.������S��&����Z�D��M���ߔg��ռL&e�z�v �W���Ŭ�)N����vh�)bܸ����v��JB���芼A���ז�v6�%d�d]
Q���w�r��R�Y@m�J�K����:��R8��͋^����4�D�/ ���l���@m-hp�v.��k0�t�E�-1
�wJ����6b�MR�Ԗ1�U�C�7Zv\(��ʲie��&�8�hc��azwoᕍ]ckV`d�Q�&��Z�QB��l)m�uP��� F1�D����C��T̫�e�bi���8qi�nKW#���=�W��X�$�{(�֜$�;��2���k[���vD��1�}�mQZҒ@��
$�/ٛ�ʺ���jtUD�,�bjŊ��-fzm�8�:�ufR�x(E@,�MkHX�iNP�*i��@��
ˀ7A6Ř�0�ejy�;�.�"�#`���N̎��&���HjfU�'u�mѼ��qHZ�A���
br����uuB��^V�ܔr�Waa�J��n�qs
f��.Ű-$�j�T�՛&��`F��є��S5�oh�2Z�֬�8��1��Z���G^k7X�v^Q�Q����x?2�8��4�V�$Е�ծl����칷)�-]�r�Խ��䫍�m���5t�7[�Z����Ҥ��X�g
X� x�S��(ɻ��@��/1��F��&7�]M�ۚQû��cm*�[4n�DD�>Xn����[�D賖-C����z)m�C+Uk��dwf�O��R����?�s-f���6-.���z��fS�Ee�w���;�ś�,f�A�ui.��e��a��āVt��������נ��F�
�6���<T�Oq�E�M����
��*�Lb��a����c%�;o1nV�c	D�Y��1�*�2`�4hZ4U�e�CU��0�KIdɢ�|Ee�Yw	b��N-B>�*dkP<��0��^^m+��4���n�#W��Jn�kE���/%����!{Zd�
k�o�ۢ�Hc\�t���}zU��3�u���t�F��PLV�m�p��j98"[W�7]Ct�DT�H'E,�Yr�j�nhZa��&F�6���SX���m\��)饏&�T��ay�<�U��+L���iN'j�����I�k]շ�QK(SxF�t�(a�_Z�˺�I����8l�h�U�u>�����.A��w%nâ�@���2��S^���"��M���{�'K�%^˻&��a${�Sh�s*�Ԋ�%U��/`i��HY���`ֲ�%m\��mk�ZE�w����X�!���;Ӎ�dJ���$M
B���׫o|1�v�+8á~w���S&�UnJI�Pe��U'���#�6Q�/i%���LWe�Ce������Bku�&����N�;ya+XwJ���v�i�:�Р�Mt�Ӕ%����Q�&@�M!]H�P��˺ˉ&����ѷ����b��bX[,	�P��C^��i^���-�{�VR�9p�ڻ���v��wh\���8���v��g׺ۡ�
��)bݍ���b��q	�̛���Om
U�J�Ik"�8j�1+S�B��cZ�-�/�l6à�0����`i�F�,�rT�J�,AR��e����sr�֞*��E�7D� v�oBq�J����"y�a���I#@3�������
Ve�6ܹ�I�-�X-Tś���t+a��*^�/p��z��������;fitέU���d?&t00ekY�4.�9Tb�N�Sl=��sK4��w��l)VH��c��%�wV*�5Ԏ��m�RR�j�˭O^�{Q��&Kwg(�6b{�5�����]:E#�l�jrx�:�$:<V��|�u!2�Y���յ.Z1\Y�n9���(tHnQu�tM�Jd�M��t+k(�9k �q��-n�d��Hlp���n�5�$p�&��c]�b����0����k�4�`HXwkme;n���J�C�ѱ���Z%ϱ��c����C���`�P��B`�6�=e^�j[)^݂�;%�g�B�a�t�������#[l�%�]wrR��eU����. �y�n旹�$$�5�VfdL�V1��f�3(IV�7`��seq?@]���+{�N��>�L�Սc� �n���G�ed
B�ʼA n��� Ņ��Y��h�*���2�Q��uy�%\y���F����������P������zZ˙��{YFΐ�4!�;k��i�cv��FҦ�:Wu�k�{t�rP4��i���sn���Y.^%��J���{wz�l��F��:Jk�²�\ú�c�QA[wP;�	O�˙MPm]c$r�whX�ɒ��ɡe��77X�B����vqM� ;vvx�:����2÷5��f�2��VVnb&ab���"0d����H��P�T�MՙZi��>�k0�6��)d��N�m,˫��!ఉ��� ]j0���R{�Z[=��a����o��_�Y��fJwE�2���k�Qa:�ཻ�8\ d:.�*�e6�]ʌҤ�%��r��&�KM]Ŷ���%ZW ���L�,�KX��K�`3�%m�m�@��S�}z��KX1����p�]<`c6�d�n�t�Y�"�FJ/Q�U�6�(k6��w�fn�EhYt#ݼp�-�u���hLJV�q�,Ɂ�K �м�R�'v�&�pZyw*ދA'D�ُ���َ�X�)�#v����%KtE�ٕs �Z(P��6-��5�K^�V��\{��H҄��/3@!k4�ۂ�-D*9�=T4*���a,Ŷ&�����f��6���B��e]`��H'H�N�B[�2ȗPGCa��`�{ @@����&G�l��B��b�V�Ii5��$�D��'~,JpMI����1��;�z��
j�)[z�lt�2�B��Fì%�0F�T߱Vl�R��$D�q�o�!��f�d3,b˷�7��Oio�K��&Z�q�N�SKP@r�����/)V��,ÖoK jx�n�I����k��N�m,k�c3QP�li����
3m��`���l%�sS��[�CEr���(q�9��zk���Λ:�t�V��C�ZgFS2�ø�{S��s���F[S#:0BB�h�u����z.,$��0lR��	�r�on���l���w�]���;yt�XLXt�
2��.��\�+����f�uR��f-�hJ��%j�9��TFf��xK;�T4oN�x�h��oKk!NGH�H�7"����H#h���ܭ4!"�ߖ�u-��Ȗa`����6�#QaeZw����m<ܕ�
��'kJ��*X!b�l)�[�K���M�Ӵv؅b1<o8�жw����]dë b*I�VX˳B��2��!QWx���w`��lLVRKWR����u��m7����Ӧ��XX̇E'�Oh�g+'��c6��.�n8�ܬ�X�E�Y�`A�	]�^��Ǻ�P=��Y@���U��4�77m��de�YYQ7����b۱-}�	m9��v��a����MK @jtY[LPǷae�Ŧtz�j@�#{8�yz�w+ t����㰚=����U=F��]0�3�Go�zҖ���S5��1�cӁ�7���=*���V��n槮�yӭ�!��̠�5d�xpK�k�PeF���"ݡ��ް���Э��Â)uwu5Hт��[��ņr�8��	
X	���6��T��׀�˕*ؖw���]<��|Z�8�\I�R��`;/7n�T�
}1�-Vie���4w�u�]4z�YA�/�6/���s���9{���C����CM$r^5[&��R�\�f�ZV]��l�6�k~�ψ"��� Ѭ�rE�f*W�bΰk�*:�+Z���/\���OM�����t��5�̴�����P�8a����]C�;�d�,F���ov-�F̋�:��I��Ժ�Q����e, �9r�%�2a��SH
@֔���e�CUf��7�͙��&��{�����9v�;��vv޴���oJƅ��t���T��"g-����i�T�xS.�{��ihX����Ѫ��j4�.ɶ�'ymL��F�(h�U�X��3���/�H�54�'��/%0��X�R�H�X�`x��D+#ƫgqe"�ۼ]���w#�5AY��e[�3�ݕPm=7z�^H��N<8��t�� Z/+�s);��3]f���QN��$.��V,3Y"d�4�Ƿ����+���z��8��ף7t�{@w��%=YY��J��Il���¯yY[ZY��C�+NR�j�b�^��`�m%E�?h�dM�)+ ����̷�f�35�jf��VQ��)1ڠ��^F��1趝̻��+�3^7t�&��%M"�Ӽ���Q,�r�������w�F���E������I�qC�6��9fA��u.�t����JA2�������F�©�ٴ~��f�s��v�� ,�T�v3�N�t��e�S(M��ۨ�7 �ݛ@�ۃ$�i-��)F�:ud�q:O�M�P��Va�
ܲVV#�f�Ż��x�6]���G�-��7������֝�/��f��pn���W+h�%i�5>�\ā˲�
{�*Ӵ3+R��-&��H'���JL	V]�C&�Ye��b�Lɖ3�݌@S-]s�Ōw�4����҆��[�$_҃��Թu��,|򮊭��6沂K^v�wO�S���Jd�J�6�.7X3F�!m"k~{M;���'�]m�4��ſ,��\�Q(�	Ӂ�4c%�ͼi�Ut��Qb,��bX�*�zU���x,]�Ȗ��8A�b�GY,�ŧ"�
�͆*�JS��+��]Mo ج,�p����5dۭ�X;.���1��75��#r%cwqeYh�61h�Z�J� ��8�;N˷����f�\{�#�=���[y`[�M��E���8,V1��W`Ыť|�;Ӊ��N������t��Ru�ׄ�5� v�=���җF��Y	yj���oHU4�9���3�,��{&Q�;�i�.f�c���`9��۳y��FC�=���$�5;�b�^�k�he]�\�
d/Z9[ۮ�]�|A��K��K�{H�p�O+��5XUJj�5-U�Ȁ0+-,Ai�E���vKw�J^ժuq��<��&�4E#kIɿa�{�(!�3��k؜W��G2�4lJ���Z%��Xӛt�-uu
Y�w�%ج���4[�.^�;�X�1��K�f�r�!bĦ�+��=A]cM�{v��	>f��j�nf1*���J��7^�lD�ǖ�D�Ѡ�e��&�d�D2�jܚ�2�^F>o*�EP'�^0�a���ut��fP��d�7�ѢݙV��V��!m��o Wv�H�*".�U�r�y�t�n�'YNҬ�c�b�� ��[Z�i�5�wK©c�ß��;c-�3ǘj�|�:�f�j��nK�ki���Ev�^^�GkKR�X�J4(3V�z��t-�t�W�m�0�7��q���5he�����v���A��e��m]�Ks�i���0��	�6��&�l*øn���jm���c17�[��mv�-Х1A�Zr�e]��1�Kʐ[6�l@1F�v��۫��Z�k��/@Lژ��_	��Al*M�w:;t�U��Ad;R�:q�tnh��c(�^wk3l�&�kr��v�[53	5n�����M��gR��5���#��K�H��;��*ܺ*�=� �܀�c�Ko��][{��(�"3Y��e�U��0� �5-�H{G-V��[CUl�m���9�p��D�.$��w� ���)�ޭ���Y|��x�T�%ˈLt��Je�%�W����&[4ڏ��וt�5[%ND
�!�V�5�5ܺ���̼eTW��*��v*^�D�ӣ	5�n�r�X
���]��vmlXM�P�6*N�d
�p�֨��*���|���W!�L��ˀ�3+0-I�ĩ��훼z
��u��Դ ��޷M��M묢�웷VDC1LVεo>)7��+e�xU�6�א�̏V��[����vo,-xҳ�$QX��A�o���HC����5��2�ЛB���u����q�*�\�(6�Ƿ/��*$Tr�dʸ�9�gT�-���Yy�d�����^t���Hs�F{���1w6�Ԇ�ĊoB�R�96��o��m�08�I�����	2��}�t��eК��g��d�&�l�c_[
!�q5��0ԭ�xoXΊ���|e��t)�۶�T��Q���Z5�r�[�Z��ᄈ�/z*����Ӡi������4�މ:�P����/Z�v��������eY�)^�o�T	u3"����c}\��1<ē�νf��o�q̽�C4�Rs���)>zͺ��%X�0���r�"�f=�V�L߈B�Ǯ��+�m�����MЃ�Ҕ�!7h�tk��Y{�f��j�_N��/�)� #���#�v'N���\�.��/��f^��gu��$zʄ�%�9ʓ<��J���2��� z���T�1lO�gp��Y�D_Z���p�Bu��y����r�u�.;����Fqr�aԕC��볚�j$��#�׹�L��O��V Yꔋ�^s{R���K�97�[�30 8���������d���օ3��v�aL���[o;���1���ZŽ9Z�Rk�ba7�p�y[��p����,�Xѕ˾&�\��@!�.J�\���W��G']27�(�;FRӛ�˭J<2:ޙN[]�t.ڍP�V�W�q��2b�T��IzPeSśY2�u���يz,�ؼ��)��/9yV���	zɁ������4��\�U��ǆ��W�:��A�����˽t�0�y\+3��aC���t�NgW!����YW�W��ֈ������#C:�[Z�����)���̡�պH5�%�0jX�y;�`���[�ⱽ.;���xK��)%i�B���FlM֜sN�N��m��:R'wԁS��&�������b�[Z�N�ާ3U&�iz�i<��]]���X��*l���1�Wc�9U�p��eX��_��-��ZC��wPw��"�E������u�(�]�6O`yB$�A����{d���Or�Tn���+TB���l�Q��&
f�w����Z�<x�R�#��g4��rR�����\[�N<�d��V�R�x����.�a��L��E�ָQ���� g��K��zBy�u4;����ZG
��"�7�k�m��]0f��`
�e��[[)o��.|��P����-�X���fe�%���,d^c��B ���M��m���Jv�b�n������k�8�G�֎���e��8t)V�S�7D��btz�鬼ۗQ���Fe67�Z�W����=7B��^U��?%�X��|.����I�X:�-�`�H蠠Sw4�f
��.�Gv�W]���Vpձ�ͼ.�j�BV�V[�_*=B�T�r�-�\�]	{G����M�K��c�Є�P���it.�r���Y;�=���pp��r[0W'�KPDJ�{�����|��L�v�H�50��ct����Q��Z=���h��kgwg��b1�	u@��e��ա��a9��(��ݡ����q������*�a�]�v�t�OGq&���42�:Ѧ��ģFѫ*Y�n�8����h-a;6��_:k��
�y(��/,�@D/q���4
�e����/:�8Od�"�Y�ʋN*���pH������~β���.�
>�wW��W�>K�ٵ�2i�U�ӻV(���\s�:��/��6M�U��I��d�TY�*��Q�q= �$��YS�^4���Y���Co)c���]�¶�n��>S��q�"�����Kp%4_F��Ɏ�"�zY�1uh�aT6��-͘�PV!yK6O��K�����
��Yy/d���{��=��W� ������c	�׵����}/��cL��n��&�4��N9]2gY��nA.��]/�1�Nؑg��8(�.�*6���s���q�67��	Y՚�CIlsQ�z�z�D��*���U�b��s�z�M�}���oHƞ�z�R�R�w:u���g%Sټ\�Q`�pv�8Cj��̘j����*�%vD��kW*���Į���C����n�Xyi�iW��wɢQ�b������V���y�p��c.���	�Ʀ����L�seMG��(�V�5p��a�Aѷ����M�[�-�L2�׭�V��Ι>�Y+��S��ϻi�]C���6�f��>.��PU� �z,d��
��v5ݗ���XiY�yfp�fW\8�o�*�ƞ1tuRB��0�|��x�K]�m���^�]�'
M+�� �ˬ]}�v�s�"���7u�*��;#��F�o��ݧ՝�u��kU�ļ�KP�6�;��˹1�V�}��)GINiM`wY��:�CXMI[�j�ʬͦ4[I��[��8q9��;�͕v�@{g-@�t֍j�wy�p$�
��;��Y�k}:����=\p��,�*G�K��k�3p��TŊ9�U�E�6��t�j����)M��O�G���n��32�W�ښ5ؙ݁wݷ4;Y�����W�S��޴2"Yi�X�Kmq��\;���y;i������
Qvj󹭋�a��6s����K��n�"�Y�3��p.��/��0�x� �d
�/~ŗ�iKs���p��RyN�}gw���ݫ^kIYDft�ՑT���B(l���*ڒ��ڮ7��"{�`zvPd�Ϗ��G�-������ǰɊ��*��e:�ÿ/�p��_'�ޕ����DQ��L�L��޺��d4H�/+�~��I�T&�bި�Ǻw y.1���P��Y[��q��Y[D�����SLM�O�+�3�CmgsT�ڇh�����ǆ����i���gsE^�Zե����Yx��ְݚ:��1��2��N�@��A9��]y�$�S�9�?���B
R��I���d�ib�%���%�uHS�m=�=Y��YV�A�����<�3��0��H�̪��'B�u����Id������!}V��Z�`q8��zò�9y���ٙՑ��kU`�9d�e�Tf /��������e�N�N���JͬK�+�풤[�]ܪٺ��Xg6��w���IPsXrqYɸT����U�n��6�r���u]�c��H����`����sl\�c��݁����]m����*{$�%�����՚s$��Κt.n�oĺ��Q{�V�J?���A`]t��,��Pv��7巈���6����o 6�� 4�+0Z��ҌRŚ�
|���K��.�D�y�n��Lt�^�O��a3fMt���u�Nq�Ww��.�|�pE�z3�u�$�Q�8ѴH�Xf�1*�l�e���X�䌥�Wl/W�D�B�6x,�$�y�.�L|����;Nn�&�wrQrG�E���U���Poonp�+x���N8uf맵�!�n��X��*��FZ��R�Y��\,���I*�o�"ε�V��G`Wu���`���Pkl����H��e����8����bU�H�n�'zC�.���e�A�1��7#��-�⻣N�^��Wv&�G-p!��c��vWWQS$������RAwWQ �[z$v�]j�������a�	N��I��H^|�0#IN"Z�CX�kn�΋3��\.���Zl�n��vxk�uq�"|*�k;�e����Bb6��=�lR�uB�>�����C�&3��n��֣����C$��)��Y�0+�����۩����v�r�X�~�]hDo��g��]J��)9�-�<VQ�(�f��U���Ȑ��e%�e�Zk�����X:^<�����|�C]�f*\!lBE����eȕ������[g�6X�����GA�rA��V8�~6�V���UfU\���M]�������jq���҇Y��b���]��f�زZ����ktC!I�F��7�:�T��7Z��ܧ|�oS(RJG`9�/�]���|VoH���;�k$��k�S�M�ú-�Ct��V�M�¸�e�7R�MZ�,8w��W�1��t����@��w,��o�ǳ�V,x���j�U��d�;��n�
��g7�F�,�l��\�X_[}RU<�˺Ҷ*>��đjx�#3~Y�.���@
�������vr�	w��P�v�li�2ra4Kܻ֮��x��-�]wL�Q�ݔ����&���S�Qۄc��un��7�]E�R��m�Z�Yd#�4���Ah�w!�4X�b�p�1�m�ఞ�8�ҭ�
�&�_it[�C}ҙ<5��v'*\��9F�;�Mz٭��N�1��3���'=8$J�JћG:>�db�.��ΐ&Ewd�TF�G��yM�R$�@.?8mͤ/:-�u- �rCp�n��<�9-�-^gB%�h�o4�o�%�7�S�qO����d�r�W��f�R�ݮbݹ&,Aj7I3��P>%YP���EJ�����7"d��x>7���5�t�"�[�r
�%�r��Y�Ԯmƫ�)3�K��T��)\��u�a�Fd]9m!�:�gɰ�wV��7��k#��-���X΁��j'3usk����Wb?D��t�ɓӘ���S��R��M����#t�N[��ye�C(rB�O��R�%;������8*�Ʒ�4�|�$�,?GڬL�s3�ḓk� �	�WQ5�ֵ]�$jFZ:&M=[AsϸvZF�3�t��K��WL�ɬŋ��0��ʜ��Oz�(�v����غ��i�T�Ϋ�W ���6��lX��b��޷�R�;\�F�N�ǅ4��Ʌ�I-�7��[�c9Rz(:�C���oPA����U:��MP���"�Nʙ��f��6Y��X�3P"����Z�;������d�e�:4�1|��ם6Po��F`�x_s������,n���A��:>V3+��P�ݎ�ǧw-��|0�&&� k3{���*ɔv����vgmj-bf�{�)]r�Z]��ۊ�)�m�K]CE�V�g"��o]oR�k�7E�-��#���9K���B�ns{S�*���L5ֵ;�^e���,l&�u/�Aj�nŕzm�RȬ��L�+���$�""�O}�V]2p�B�m+: ��j��sr�����c-L�*�]�UͻIV�#���գ���=Nu.�#ɑN�:Nc�}XیK�E�N�3��m!��l��;{�tOUE�i�LG8.S�2����2]l����ڙu�\�}vR�>�u��+.R#�=�c}����:|�@ax_i/0 ��� ݣ��|��SU{:j޴�^.w�4�a�]���*,j>Ne=}�&õ��L8�G�>�v���`�պY(b�mS2�nħ�t��u�u3�QI�;��ӎ�m:9Jڊ(^`Ӕ��_
ݗ���>{r�P��3{�gH2�ub��S�����0��
a^��\�:8t����1N�r6�t�q��oi��Lb�2e���2ґ�f���k2
L��o(�Mqq)����+7)^��5�ӄ��`�вőD'nY�N�.��P��.�YU���{*��� i� ��� �*+�X�)�׷�[��v�`�6d��9���܀��]��3R��kV�_M���4�zWj������v������Ă@B���;��U5�'1u��h�3uZ�"|�E�jn�E��K8e���;cDTohK��zv���W@�d��橂3p��I�d�:�4pw�U��_(v��uvmDztX��$��Ob��e��}�w^8L���ڃ�R�/��ٶ�C��ػ
Z_=t���K-��X\��9y]��h-]�J��S�ދv�w�F,ǰ�@�����%�q;-^�}m�P>t�V-[U�Ikݡw�ַ�n�M�ppsy=�ԙ6où.����C+��Y�3����޾JZdt��`E��u�޲-�����<� �U�Nm�T#�Y
%U7���䘳0R� vV��i��efE �޼�/���˩܌��|��f��tS���8Q�G�6��4ڰb��2�o%��LB��YR��HQ�v�L�Vu�щ���qLf����KJ`�ٳ2��C]L�<�0"d-v%����83�SjԳ���촩	����I|&"�{nq�`����l�/�v�F�����S��H���颐|�ڎj���7�4Hk�E:��w�!8u��` ���k���Y��.�{B�Y��*��<.�>�g��/�۸�T[�b��:��V��i��\e��[�u,�H��s2}2����z(�YN+fb�v����w[QJ�X�����f����^i�8g�R��2���.r:��9j�uϩ9�T�������LP����Ɖ<�Vj�Np��o{����t.+^��"ChNa9�8�F[_t�Y��d�R����t��p]s���(ȫ$U�)�;y��V^������#��iZ��lȮ�v5�e�3�'��ǜ!�v��?>bN#s���$���Y�f>^��JD^��L�*u� /���<u|Mu(�rr������@��H��du���\���Ө���Ұ�v�WW���-�p��R)ۥ�b���[mR�nu�l�4���k	�����$Q7d,�LjV	6�>U�^���&�r�:���j�������Է��>f{�y��G^L��ӝ����1 vN�0-Ƈv���@Z�J�y�l�"gym���a%%1��CK��lމ��H��Bu�B5f����T�4�.���a֡��A���xk9�\-�_s�k܇��4�ǰE'G(���a�5:���2�ޝ����tF���&��\����˥e>!���*�H�
Ӿ��Z`���&.	]�Y��ޤR��r7{��ʣRIr�0=���	!I���~���-�-�/>T�-k��0�8��6VU9n쿦��7D��f�&��7f���if�,>�k�ܥ�M�ݻm�E��[�2��c��ݽ"�R`�� ^�n����t9�+�W]�2u`��43k)�C�W*�9�m@�<��"=��9�>W�t"��c�`�sC��͗���
Ysp[�w��Gv<'�K�ViV+9��`3���9�|�B��m��T��&���
�ӷ��C��moMR���6,Y��Śn��S]M���'m�]wɍ�Y�U�P<˩��5��z�<Ef��du0+UeaZ. Fհ��:=�u�A�Xj�K��	���Q=�s��������E�ն��Vq��ٛQ���t���E:�d�݇[e-#6���R��;&���K�pn�<�u�����r��y�!��������p�yY2�.� .ݖ����#�\��<��^�ǋ���smO���Ӈ���%��2и�+1�wJ�r� ;K�OFA����U�nج=o
I=��Mԓ
uyZ����Ӻ��؝�u��r�6�FT�yE���K��*�$H����ٝ�ڬ���	��9�3�f��
����-��z�J�jBv0��/8���z��v��d:�\��R��X��i
ׇh��mgX�5SZ����'*mP����:/6�=��[�^���C�GY��m�}��\\RX�o#ѻ(\�^��m�.VO���@�Zf*X���
�7�����qjMҺ���՛�Z�ͮʋG:|Ti���TZvB&'�jnV������ۚ�A�(1�m/�f�w;9a1A��ʼŵ�Ê�<�:�ƷF9 gpŤ�(�o���ʴ�)}��v�
aܵp!e�a.5����r�@������N܆�&�Ꙡ���x/Ƥ�(9}{a�v��k!�z���V�D�IX*9�Wv�	g�]�Tx�����q�t���v�����x�Ӭ�7AM��o��X����QK��hӋh�;�Ô�.A��(OH�˺�`�o��!$Aש�Vz�/��@���,�gi�.ZQ�I�7��G�b8' ���#7G�6�S�-k��2�C��ȴ
3+L�t�lQ66+�Vtݐ�l�V�2�r���5f��x-J�E�MXiRf�F4Ӭ̮����+�hG�w�rA����m-��7V7Y��]yDag>O�2�`���#մp�}�7����jժ&��,�:a��t8�*-K��X������F�s��mMx�pA(��kx0h������+���W�ef��P1��w�ϗt.��9��z:��eҺ�����GFM{���)��-ae��ZM��9:yI�Փo�
-�4.��=��{2��5��kC�Y)�R� Tn���`�[+8w�f!��_P�;Pn�ݸ� ƶ��9F�.�SP訇$p�b�^�xze5�֖��/�1j˶�u7�$ѺE��m\]>��3:^�-a� q���+o��ʓ�A�]ǳ�v];ZKs�(�kƹ+Yr��_�Κ�5�ۈގ9Ǫ���u��F���W����>	1x�I��*�!0�s\!佅� _Gd�p;oN�����'v���Q2Vwo4�n�D�
��dܗc��t�]Ϗ&Om�ywr�W�nd��hA]���l���+5�/V��ah�Z=��4�5b"��'r�Cz���T4�V1�N=�0^�a;\u�+xؙX�u�/�WV���Y9>W�i�N�����z�ݥw%pt��g!��㡢��Q�Z�Zءo�F�3��E����e=�O�.��
���#�ۮH����F���@
\c�MK;�C%#��ʤ:�5��Q��ɨ���<�%Ѹ]�+^h��g`�,4�v�ɴ�Xx��73���ɑlT�]��8�O�|��A�|vl�%��ӱa�����S�!��/v.��v��&Uӵ���L��`T�|��ls4�;�9��P�J�i�ۺXZ�"�lD+�eq�畇y�ty\&�iM1X]锫Il0�F�X�-�']�ک���u,j��bŭi=֕G*h�`�����si�����nd��*B���5�����k���H������{r�ы'P��.�L�Sa�3iu�h�u� �����lƷ�\����:V�ή����ɣ�'����w��3����g�N�r�fL�{�v���ԥ�N���/mY�H�̒�����&�Z���K��[���u>|�ם���v�ƺ㾵��!�y|����Ԩ�.嶉�F��� rQY�u�KW�X�c��J�X3[b�.W0�x���6�:3�G3c��t<�A�Y�w����o�0��W*{ɇ��5K���PU������Kytw-0��˙8��'.��ְhhRܻØ��慜�p��)��R�J�Zw4�^����e�G���ctu�'`5����V�8;i�����sH;�V��>g�v�J�ƹ���J��Mى� ��Pv�J��V�D��$F��K�8�y�ԙ�$�t���u�J��dc�����[�-�酼.�d}XM���73�ȱ�nL��c��F�R��Z�ɩ� u����U��Eڻ�ԉ�7{Xae�j(XA}0fd�Nv��e6��H�7�ZUS�Z���ۙ�)��Q-�gYk�W+���wّ��m^ Vܒ7&�ÔR�7ϰV=�8�]��y��!�t�qa[p�{و�U�$5n�{+wJ��i�	�e�$Z��A�qT�eU��_d�@��9������/��Xڌ��>w��]S9�Q�Y���4Qr���taN9�ى��ƺ��\ùSo�oP�On��Īq�DkW_sC�4]j�x$�\kV˺���Y�78vH�v��l%u���FN6]\̼Y�Q�.'�KB��c|N��2��l٩F|z�cvOd�:�r��{.o�u�}Ӣ��ѻI뼣cȔ�8͎ �;����P��[�9 ,�MIXsOm�f�"�BÛ͛�|�h�7;Q�;r���� �����h�Nb���[�B��/�`96s���y����nY#��6uʓ��E��{���g&�<>܏��.�q;�٠�� b�w;]��������q�;2v-YJ��ru�;R����N\T��g\6�H*���� ���k]@l�p:�΢�],��0����6dW��>.j�=�A4>�ע�M�$W3|owl`��ݳ���ٺ���REt�s���C���m�H���E[\6�� �t.��
M������b��u)c��'Yk0��h�B��c�\���tqeZ�IT����C.�ڏ@�I:�� r%]����`*���-G�*iP�Tp7�=����7�� �h\�(�ZZ�+_o>�/��S�����)��mY���s{e��<SC���_>p�#���"oq⚬br�)e㛆�j����]�P��h��>��/E�j�������MoI�Nn��nF�`%�R.���������Zv
��w��t[���*�[�����ra4%��b�~zi[�
��bn�ʳ/-͂��/�ݻ�TO��I�w��*�3n���C���	�}R����ԡ�N��0#q��+*�WKf��U����e��|+gc#�%k�m˜4���ݫ���S(�Dr]s��+Pn���F#�r�h�9N$6��*v`T`Z</��%=����r(68~z��%>ΎZK���;6���q�����S���t�'�������)؏��7���$��1Sn#b�WԗX����3���rv��2m��i�YN�"��l��[���"L��T�)J�kl�$�뿻A8�;J�$�Œ�8��	S�VTf,.����UՆ��lF*զ3�%��4R�]�������s�*K��Yc��2X���t�[�q�ST�����+��1n9eޝR[9�7	G�	����]�:��5�\���M�.�9� ���^��w����<��+2�8i��f�Mc���R�
Y{�A8�����-���r_�WF��k�b�a�w��YN��e�}�ݝ�A
Ӌ�"u��"7�wa�Q�6�8�����#2ܙ�5Nc��`�\�-�3��g10oKG���9�vH��Q�!�q�����P��y5�>B�c�Me�ʰ��Ʒ6����uq_VRj�܎��ĨréMF�Is3i�,�ˢ�r�VVȢ#
�z��{�q�sj:5�sǆ���1+�}�kB"��Bֽ�
Z��Wlٮ�nn_.j0�\�y����'ۮ������R<h���ܥV�ׯ6����2�v�A|tw��qQէT@Wa�)�m�B�j��"4�:��oB���'�<�Ɔ�?9i`$�ҫk�%áe(s�n�DVb�gi�o��RέM8�Z-3/��/�+9v�p9�Y�ΔsCP��+؀�(��G�K�f�!�VА���Qu�s�*a�QZvL��-�+��J:����J�4	<��W_�p�Cަ�T�v;]!�Vq��L,E���et��͠���7:��CC�v�U�{���qG�d;�A㶙B��pK��ֆ�gz�nK��u�����J��М4�&�S���[ʰy���1P��}��|Ȣq�u����Μܗ�@[4H��I���*�[��\�X�"V�L3���`Qh�K��Tki\+�9�+X����bf_@�R����dé|�rX�%�H�2�^�'T�oa:j�b��� ����W��a��Q�ea��x*�1Vn��{�e�����+��Y�]����v�tzϹn�`�Y[��l%���;%��1q��D�ֳA1g�� �����> �nL�����Q�����b�$}Hd����1Q�f�:�5CM����ؕ��%_,O��]��kQd�4�Ò�=�aq�}B
�u�H�q>�܏P�S+[S��,�O*nd�>�L]�5k�v�|��ʕ���9�l}�W��6�be�s�4;wf��b�]��S���f�f+M/�[Ě�)nʄ�쮐�|U����tk�͜�[��5]M��e
de�m�������c��;�t�AX�w<Ŏ��	�<,�vY;.'t��h���|�^�Le1�U��Q�{g����芓(t�m/(�U�a��H���z�V�i<Fn٫TlT=�NT;���Rշ,����u75��^R'f��>i�s{�WCLr_�B6�@y?��8c��<:��;V�yvn|�[�Eєx.J7��`�D�j�RҒ���5���^���ᾄ�A)T]X�KG�.�<���p��vZ}rJ�����$��ǻ�DR�VgV��"�Y	L�"�6�B-�^��\�*iYd���#RT�t?X����s���+u�1ٓ��Έ�U7/�b���m��	���h;|���M(`�:V6'E�7�h���Ex�Ȭ��g�̅��z��T��i�]<(L���u��R���#d� �ڮi���5�įYN�r�H�M�H�o%�G �����
�p�=y�k;����ES��'>�������,}w�uVq�$<������D�3��׈V��R�] � ��O��km�[xSu��16vԭ�6x��l���MΧ��c��|:�n,�l�з��`N�RC��oj`��dv�nܧ�fGl\qoj�z�/�$[J�V�*��V��m�++ak��.T�6J�[��
�͇x�|��o#��Vj�(��&��R��yB������L���j�g$������fP;�]%Hi��mT嫛���;}����1���1<bU���6p�
צ��P��f��Y]��mp�th����ֲԳ�2�nl����!b��1)؉�Y�J ���8o)[P�noQ��R����H)���)��:����f�c:�A���=q��Të-ݮX���HKS���Z�rj��0�GB����oN��c�$l×�S +4�pw]8[�8>چ�oML��c���:���`�g1��Z�Y���.7nIYvf��2![�$����ae�E<?XO�l=���Y��	W+f�r������D��,�AD�(�9�@ܷ�n��¯lSd��n��*�4f�ut�Kg�w�("փ���Ιr�"���r]�gv��1�wlVjq�r��1'��9`��j�Z���f�S9��'�WZ\�����X0�:��#�oH�UvN��z���ޫ��8�m�]Yvw����"]�m
��f>leRS���[t`B\��^Mj�ѥ�Ӛ��2d��Tw"�e���o O��B�݆���!��̼׆�8���[͡V4 F�e��0�)��������̭ 
ꝗWI�1F��9�Ѹm1d��4����>ݡM����6��\�i����|w*ʲˬ��}�AE@S�G�.� 2�9�eNc��B�K3;&`P2.���Ǧ>jR��$ZT��e��VqZ�$p�S����F�vME:}R�v���^�X"�K��_vS�%4p͒�:��B&����м:���+T�F��]{/�a!'w--T[��W]̢�<��w�E;ԥ�-��Zi��r^���:ɽp���ʜ��;cx��B�e^wdM�gG��jbƺK��t�@q��u���4l�eNJu�K4�ӥ��p�.J�ܢ��e�=F����,��(�#lܥ�Ь�Kje�J����Y�a��p��

��V*!jgDv>�%��.U����c^;)����N�y���*6�S4�z�N�tϥ�y����'Y���4�uk�=b��s�5�>M�y2�������Y2tI����C������=�O�d\�r�۵c�wMS.�Df�N���d��Si�ɲ��^�6��q�q��Zͬf�.nR��Q�M֌$۔���� V�N]���s֍y;�m$��a� N�~��p`��؊9f}��u�}+"��Wq4��&�D5����P՘� �y��C��D[;��kܔ�����5m�v�V革�54U�A5�䒖_^$���s�9��r�sa��mN��x˒P����M�w�5�*�T
����E|���U�]t�A`��H*O��E��Gh��W�|��c{2�k���3���{*L�u�:�%��r�<��@]+�A�%;ٰHHUb��\��{�Z�+���oq�'0,R�k�!�W�f��//a��e鮺�	�J�b����#q�2)N���R�iD@�َ�,�b
���Pm���N�q��l�U,%Ӫk&,͕���i�U�<�v���lD����2y�e����MW,����)�]P��;�P�9(�����V�Mꎭ'��]����J�8�0�mA�l���Ѭ =��f�y�P7��)-��I��F��׍nn��<�U����Q#k)��{��n*z��0�T.R��	5K��,�CKT�iIՍsnd�*Ջ���[�ٔ�^��V�+��Q�(G���e��F8�,q�LRI봶1׵(�Ͳ�o����ݷ?oN}ޡ�GMAk(m�j��j���څJ�QKJ"ĵ��[X����PQ�0ʠ��-KZ  ��L	l���b�mQ��%�1p5ZҥYZ����j����ĭ��5�X�cQp�0��`���VVR�cR�Xˆ�[h��#�e���Ċ���F�UR��6�0�[T*����e�Vڵ( ���UZ�D��T�.1pңKjX��kV�[Z�,Å�[J%�P���J���4P�j�cZҲ�*U[J�-X�L
E-mj����
[h���Ҕh"%ū���ҭ��llU)lmJXV���Ye�Z��8K-��D�Vն�,��TQ�5Ad�`��mJ�-
�F�R�h�*�b��	h��m
�K[�
��b���-��ḸĪ��Q�QB���\-G0����}L�N2)�����ufЦ*�{��^H�Ou�h=���p�zz9� y���y$Un��e�$6\7�s�+�s��W&��Ǖ���9񚫏7.�\�J��J�mQ�ȭ�z�L�Պp>���(��n��ޠS���h�-�r*&'Q��ɉؽ����g[�Yv�H�R�)���#�1�:ϑ�x3�'�:����5�1��n=�Y����/,B��n�^��"{[����l�c���^�sݺ��n�lf��u�/Ҝ�b�y���ɋ��9ն��c)n��Z��Tk	^鴎=���8��W^B��K�d���ٞ�������٩Z��E�ݭ69�p�/w��m�Wz�к������޾��#2���(e��fse�r^���N��A���{U�m��������څ;�+g��c�r<��.oo�S�|۞K��z�ݡe��0O�s2l-b��+|h8²pw�������z{7�?�^�2=j�V����3r����@�ķn�ʋV
���|%S�9�B�j�:m=^d���h���k���*׸��%!#Ve�j֚,.;]͢o�9�z`r�(�ջ��V��&����ndr�5Ȣ�̩!�p��)����Ế��f�+z�bkd�@�boI׫;�Ҷ�x�-|;:�P����Zr|Ɲg�r��x�������h���޻��P�Ң��ח:3����#4[g;�D�'-�f��5����u��ί7eה2��O,��..�#�*�Vj��i4�r`�wc�+ޚ����|�ƽ=C2C�M����t����M�+`�Q�������&�)���s[X�=,���=
��1w"z�nV�X���w�����V��8t��
�M������95w4k���76���d�C���S���R+�N,�c��#/��Z�Bݵ�
5BٍF#<ɛ�7)���U�gdZȃCv�
�S�\ɭ���C�Z(�7R�d��][ys�j�'<y3�-�<7�`��Y�X��cל���6V����͵��euX�#WmvJ�-�7�4�b�����JI�H�jw!Qh����R��]ʺ��Gt�_:	c��-%|s^�+C�ĺ�p,��3�71��'�9�$Dڡ�sSj۫����n�zm�(%Nv�m���$S�%a�/�l�]B�ىZ�4����Z��l��ђD;ޓ���o�0f�3^n֛���^KM�����eq��o��z+�k�5����!���ޤ[�[�}�5��T\'�)�b���M�_f��5��t��ƅg#�j�6v�Nr�V�0��y�95�R��	���z�E�/ӭ
�L�+YW��1wO��-[�	�f���M>��~UyMۍ�f�Ї�i��4m��n^�k^TC�\uqo���g���u����V*QJ��:N���ǎ����v�(_,,[k/�o]������>9�ݖ�(C�1�:͊�L�)�Wy�<��|O��N�q�k�b]�{�R���yv�<�3�kc9���^�����tUO�uC��G�����:�}���� ��:u�:��GK�z��r<J���W��^���X�W�|sVx�2���1^QRx=��10G�����m˺�HhP��뒖pǐ޶
���fy�1��O�';/}aߚ�U�8aLg�^cͮ��k��w4�w	; �/����$��F�=-��j�o��o*h����j^�jF�C�%���1Ǻ�Wk�Wa�c.s�,=��}Y�n�C���&��5
,�_l�Aj�βxf^��'�SJ�s���)��7\!��C��&@�������M��!3a�Ro���kw���j.��v�B���cCehM�úaQ/O�(��e��8d\�A�R�J����ސ.�м�X��n;���a~�1��f�S�Q�ёۍ�Pf�A�C���sꦨ^e<xw57͊��C�36�^O57z����zŏ4Voϕ�7�]ziBU����J�#5�z9�	wU���Ye6�0?wVi�e+��9��S9�Ĵ/��&���B������­���z�|p�t����F���yF_gD���#�$�>;�s%J�j��i�[���s��W~���z�n;{��W���l;V�A�A8�u:�N��{�lOk|��g�r�Bya�-��I�`s�q�WWb��IZ5�O�r`3���b���cK�8[}`л[����͛� 8�u�6��|���`�|�*�9�[������;#�����)-��wB�"��ˋWwL&m�<9 R�{� ���T��-�%�����T�^���yt��]�Ǵ���2/�5i$��P�=.�n}i+�N�پ|�6wf�5�^�]���.z���{�]�c��]��<k�:o��'���s<������E�TU�������9Sk$p�v<v�|�&��V��'�Tߓ�w�J����)#�]x s��Do,w}t�k���I2�թn��.����/[�Ø��)�:Om�l����Y�y��۾��Fs�"��r��W��g%8!+p�&�	3�&s�UN2��{�s�Ě,F,�{���9�b�u����^$c��򪾜��iZ�Ɩ�1L哭�e�O	]7X�ׅ�Ȍ�n+�S��]^�Eorr�X����d̆��Ӳ�ۿt!u��r*�^\�ɻ�/2�:�x)њ�U�W.D�9��z����Z�o@</hז%\��h�ɍd� ��`4���w0jۛ7x}���xŜM���ض�^(���&"; �z̞������7t���$M�>iޭr�f=oZ؜Ru���%�]B��qKIe�oT��,=l,ћ�����4z{7?i�J���*c5=*z%IYY<�a�j}��ϯ�-���y��E3~�f�������禙Ŏ����9�)�خ~{?��}6�sf�[����vߟgD��s�v9%ņg*kgNj��lz�Lٝ[E{ԧ1;I����O�^fť�be�Sҽ�b�������!~�hW��43���J�6]���R&�~WVUj�L�o[�ՏI��s2�w����>+K#�Vt.���:{�6�ׇ��Pٔ&)m-9Z��v^ �l&��u��P�ۅ9B#�K��N:��Ɋb��C�fI�=ېL�%̦�%�ǳ�>9���
^]x"9Xɚ�֫7�����VG�gj縟�vqrh	OzS�Hzz�:"[e��q�٧z�4S}�C�P���/��ھ��ޔ�)�z�VS��"IB�[��*�S�ܐ�!��(Ї�P�
�r��;�9C�=����~>co<X[�'8�/ ��)�{����Ba�ki��^�| ����]u�K�7�s�E��M#�4���6(ڜ�Fv�n���&�ތ���Lq�	�qk�.���MzT��|B]p�:&�}{g#f.�.���wq�\�7�kT�Y���O�	���k�u�������g<>�͖�r^3<�=|���(���9�ν�Wz�`i=�tRM��=��S�9[���j�V�Q2Jzj%gk_a����.n��P1!�H}_InXY,p��[yby�kq+o�ڰ�]�y��ܯ)�&�~�lSei�s>n�h5��yl��^���M�ҳ�x箳UT>��9���U�X���o��op�{�/��F�}pz0��w>���a�r1��ٯ<���1]c�`(���9�L�WD�j4�o�ԝe�d� VJxЯg)�u~+�j���1E�Iy�ǻo�m�o�f��������t^�	օz�2�yK����l�M�ġ�Ca�V_��m>�v�T��n�����_������&
���.=k�J,5�ׯ��-C���ro3��J�&;��)��(�CBW��zd��>��kҒ��:����=���n�6�>/V����ȾiT�ag��*���)�bzb�~�T���5W�ۤ�Ҝ�1V�8�W�.l�{c�g'c�3�}Um%Y"L��7��B!B�LskyL%���f��&��I�V����e�R�w�+����Φ촳���#0�L�X��q�6t?���z\�B�"�<��HW�4 ���3˱F�ع�X��x��lV�L�El��=�tk��2���v���R���E]G�wSNf��n�����rY��"�<o�����O0f�w9�JX�kY�d�*L��u�\��T!����s<h����~�3{�o���>K{Ґ�y��X/9y���r�W��tU>|���;�)+?<�+-=mN�t����d:]��D�M���ohC�v
�Z�z�)���g:K8�s�ig��nt�X�^c�b& �n;��l�41���L�1o?�/E���9�>�l�~�w��r�*�
��^e;ǧ5�͉�"V)Zך��\��Q~h佽�	a�~(^�/�.U�K[��B���a���V��0+�K���8.���f,or���������Oe�H�l]�����H-��/��"��2���:]��7�.�Gc:�3rv�//�:�v2��)��\�i��ѻZ��@���NWgJr�����ZE�TW/iuM��
�˾�6(4)�����ߓݠ�:h-͉�43h&�oj[6�f?N9C�i��Ho�{�Ϲ��͚��Rݦ���J���aж�-�O�r�\��+/�Acl�\xg)�r��M퇩��v�lW���0�J�vD�d�.'v�Қ~�t���=;�P��Dr��;����z������\1�&{�(s=:�?|���A�߀�BX����ZR|�(|����5<i݈v��^�Un��z��:P��=/.fp_\���-9fZ��%EvJxT1[���\�����>=6�p����N�2h�5��C�&�я���=4r@���˽�J�s~O�߆�*��K�V��[B���"����3���I8Q��2�:�lt�M������U�*��g����Utʽ�iw51��n����7{�+:�{I��r�!܄"�1W��g�f�ZV ���H�nCx*J��Ď6t}��F�n�V���%�f�g���F��
褩V�U�V��"��;\�&]&D}�ѓu����cÝΈ;����TJM(Β��-�𜔵x!ȫ��!�M�Y �⯊����K���&�J��YGOZ���"��ohB��oM3�������#:���r�.��|��K5�..���&W2��!��	]7X�������n*��Qt����=2��v�%F�1��n��Vmߏ��ח�N}U����w,荤�����9��P$�x���7kL�x&[�;��΋�m�sY3��m1�D�ud4�F&XW(P���2/�-�V��o~�S7�j�o���$���>��N*&��V?ND���b���s����~[䟺M�r�yhQ�Ƈ����)#�Q�����G�zPڬ��fuo�y��Rr����z�bqp��PZ�&�uos��Ifv��1�gk��Ȥ#ӭ��g3�V��\�P��Qjk���R���������iS��i���s�c�[���\r�%�,v���[�==fL��5��,�M��(Em�S���K�~c���٣84Fg�0�%\���G���e��ӪP����ߋn�i1]z�H����2��+W(l5��}����w]��&�v�\7:��`
:�cH�ni�|+�p<� W!�Y"�/���d�(̚��L	)lg�q(��u^���WEd���F;7T�7(E�������ܪ�h�=a��L�#{��3���\�be�����v� Τ��;���)u!c���]��f�.�C�����r��v��`�C,eU�Es�3]s�	&���$��]oov�q]ܦN4#�M��X.b�bf,���];��՚�nZ}�	2�Ma����VgT�e1�vgP�+�T�v#��}�1�s���Zi�Sa��D�L����e�� G�j��;��ȯ��*�7F�f!,o*�goӨ���'��Wl�6�-�%�swN�Tu���Q��<���l����s�:�E��p�,`wl�V�n��q�a��#��.��aS�pTk��mKm�Rdg�R7X� �&�M�p���Ӣ'�Q#��c{�s�Q��I��7*��3i
J�CY[]������e��w�K�b;���ŵ�<\��
̂�Z�w��N�ɷ�q�Z�d�ma�+N��[w�a��1�6k9ڎ;� �솵
�݅�B��m�J.5��|w�c���v(پ�����x�Nɺ��\�*X�΂��;X�]�s.�}�u�x�8�Te�:ϋ���S:�8�}��ѰG2�)]^�'�q ��ݹ4�Wqʜ4���+���Z�:=sgPC�ّRR�c!��K:a��pIvX�����L��{c 4ɗsN&��y@����Z'��u�ٳ�D}���ߦ����t�:�t�I�if�R�g=DU���Ӻ�q�Lt�{�ۥ\��5�`�zf�°��8^�*�a�,�rXn�(���l��% ��Qk�}��z�
ȯ{�c�8���X�n�M71L�uJw�ݜ�C������4�\���s��w����̗ySe[�P����׸���axGe�T3LwV&5ȩ:%��=�!=��ˬɼnU��kÖ���i�g�!��C���Ri����l�n��k�{B��{	¶�����*�d����d���M�6h��B�$W�W-��r=� 4��+E���K9�j��X�i�uj������↻q��w�&�hje��e�\a�H�1F�6e(Dޭ	�*ܱ��κ��r]%��g3IJ=��S�O��r����PE���p]>�t���]��2uh�8�@k�]�'��v���E���2�T��Z�eC�wr]��]9�����X���ǥ�c�[뎊��9[ǥh2�F[��oU�V��m�=�Zů;6�I�
�`����d�u�s�;v�� �ڲ���ƮF4n�imn���K�
s0턆er1Pˋ��/!�@|$ h���eŬqL`�pb�0�R��[�U��+m�Ĭ����5�h�Zj�,H��*�ID%�Z��ڶ"���QH�J�,`�j╖Ջm(Ŷ�U
[
0�R��Ub4eaQV�cQ�DQ�((ơmZ(�Q�����J���b�,X+U�kUcR�-YJ����U��VV�m���j�*5��H�[[(����U��5FȢ�e�0�L(�Vڡk`�,UY�-�Ŭ�J%J�Qlh��4��iR�(��-���V%�����X1�H¶+�bʒ�-)[R�e��h6��kKm����Ŷ�R�Z�j� ���*��)kjU��Qk��a(�j�e�X�����U��TF�Z���T���)K-�AV��P�1*�7V(���"�$FQ�[UT+*)Z¬���Җ�Z�Fڕ+*�n�u�7t{8��;�%e�g�GEw�VVn�Է8ؖ���%�]��9Ʈ[��������.F���.p����8�\r�r؎+o��V�Z{�ǳ���t2�x��:fz���y+��ګS7zE��캝�"�{��)��*Ǉ^:";���X��;����*�X#]�+�lt�M����}K�dO5�znk#b��Qp)��4��W^@N}\T�V�P)��+�P�6!ix����em���TΩb^nɮg������eO��HŘ��to��=[uP�OT�;=fsHΆ�h�:*�|�Y{�Һ}u���{���c#\C��>Sz"@���K+Ey����WW<�ͼ>�j3�h�Ss5��ջ$G���u���@��b�+Mc����1���Q�J9݁ʬ�z��ɮ�bU�g:��V��sE�f�n֖��o=C���c�'=`��f��=�"�q�VSV=�(V[�1�͜�ܵ=��Z�r͸��w0k���n��\��I^�2�X��g�p�Q�U-������3���G ��*R{Ĺ���][S��CivM����6���S%Z�m�ްE��M4����K�D�\p^�5���qD�Y��ʯ�Ί���ܸ�kpMI�7�ճ5{��7ܦo�c7��]xZ�U��)�zVtWd|�\��,��נ�t��9'��y,��eCI�a��'R�ά�1�M��Ѷ���O��--�|����Uy^n�m�����U�\g:��M]	�v�,+XX�5|�9j��凥gZov���n�z@n{20��S{���6���E���f%�ް�$��a��V����.jL�s��'e����_����'��T����{�BS��WSC�#�՚n*�Pk����!�xP�T탕C�_FM.���幕�V��r�o5g�awl�����ؤ��t���@@�>�*k^D(b�2.������X��MN��ٷSe����RƱ%�A�:Z��:S\�5��]���R����X9�����Y����n�Cw��:�TL�����z3pK��rK79�����]Hu���K����"�j嘭*{z�}LS����e�f�qk�4�V�����{��5,͕f���ٹI��S�y���iw!)�ҡ,��2 bz;3v�K.���n.	�8�T����K�f4n���#�<W��I�\^S�8������K�R�b�G�W'��9���]�~[��{�8Z%�tu���Ssu��ݢ{�m��b��Zn�LS��@���k_;K7�.��������R�C���sꦨ^e<xw5�\�ܝ��e��ݮj�Xa+�68��q�8��Q{W�Q�8���΢&#���=���7�����W�y��ZS��g<9��'�O��Ri����H8�H�P<��g�W�Yb���Y���s{zx�2q���|��:��T��:��oS,�L�[��N��;�d�&ߒh�0�$�{�6�|��޼<���Q�}�@D3�.��_��[���gxƯo��[�^��OS�,6�L'�~�x��L��4�:�4�m�}1�L�OY�N�a=;�2u�o�5;�$��>�>�	�o�N���<�]߻��\�[�ݾ^��N!�Y6�2|̘�l&Щ�l:��y��u^�m'8�2j�m�X]ӏ̓�7i�N�a:w�d�O��g�s�wy�s���w�7����M0<Iǧs�u!��!��'i�,���'��.'�u3�XM���N��<��i8�ĩ��!�N0�)�l��.|{0���u��8�\|����l�L���	پ�m&��=;�I��q����C�ÉY6�Ò�Ci4���m&u0�6�bÉ6���{C��d�o�&s��ߞk6�X�_n������pC���')�U�4jI��;1n�%b��K۝y:���x��� �����٨�yZ뵹S��ǁ�c1K���kvq.����b��&s3kH[r�o��͐�n�0�wo�T�m�]8�b�"�ԉ�]���\TNn� ��� ��nG�'���:�oNwx����'�w�T�l����+2���h,>��P�&���l8����m����q�G;�{���o�G�>�q�@g����(z��ht�>v�xɓ�`�'�P�'�� m'��ϻ���'�|ĕ	����Aa�@�M�i<;�gþˊ�}5=�|237W){ޣ����d�N��l�Ր͡�M�����~bC���!>@��pm�S�M��h︄�2�!���Y'��}�J���۽4Sng�P�}s������#�}	*�6��w��'��k$�k6$��Vq�4���~bC~����󸓩�M ����'�F}�N{�����Ʒ����Y&P���*T���IRm��8��&�4��ya8��y�5���ԕ�!�՜`i'Xfox�&�Za��=@�=��?T_`��ض����w3xA��Dw��N��&f;��N��^{�*I�ޤ������d�'ώO(N06�Ohe�	�hi%z�z��L�����ߒ�������?N��J��p�OwO>A`}�
��4�Ν�T�d�w��e�u���J�w�x�d߶LRq�i=t��P�`u<��C̏m�1�Ґ��>��w�1�v��|%8��~d���O�Y%N�x8��N��N$��{��4��߽��	�&{�y%t�;��)=~`d-��#�t������뫻0~'"�3Fww�HVӽ��'Rg���h.Oi'�u5�Ad�<=�2u*=�'�8��T=7�@���L��^m$� ��C�t�z����f�E�f�7?9���_dRz��a���|�C�ChLSL�:��vO��.uI=C�svu<d��Z��u*=�'�:�������}�}�v�_	Â{D���Go�P)�[/�[ZV�+9�;hS_Z֞���k�Qؐ8�����}ģ�yBr����Ǫ�,�2��t�"ε��%hι��6wZ�0\���C�E'@�ӝ��������z�n%z�a��3��xu���u�#��3�>߶������bE&�03-�d=CI�g�I�&]��N �h�ɤ:��3T&�q1�N&Y'����u���'��OH�����Gw^�9Y���4��}��'a��̟$�����O�;�|&�!>g�����O�8���L��Ad��}��'Y3�&�q'YSHM����}|��Euw«�c��������}�d�ӝ��N���&��$��>}9�|$�|���H}�!�x��f�'�u3� �O>��N�`;��݂FOӿik��w&��=�y��}};d4��s�:�$�y�N��],$��&�;�:����μ��C<����a����2i3�a�m'�뢧�8Hݬχъ{� �,�}�i��C��%`y=��N�sT=Y2q������	�N�Τ����qi4퓻����m6w��%IԆy�N�Y8�O��J��}1=x��������}�̜N�a:��������C��r�j��&�;�ud8�����$��Ri�	��0�e�\�!Y'��|��E�ӻ��]��z��ޟr��,3hI��ff
I��O3a���*2u�!�C��I�����Xw�oO1�i��O1��3��ջ�U��7�y�|=�E{�-� �&�λ(L��!Y6���P8�i4̘,':�f�mI8�3a�M:d2�`u'��{7�q��7�}����b�"�U�������Q s��>��i��s��dɎg�Y'P�{�T�'�w��+&Ҳd��6ɯ)���&���XN!�����W���:>�?N�5��yb>��l�|>���!�7����N�����>Ag{d:��>��|��L�g�*T����+&� {�'Y6����ya8ɶv�M�p�y��	��#]9��ɎRH?zX.`}f��ov�_Ń�( ���>q`F�y��OY�I�g�^0���-e�����1E��i��H��,mpu�D)�I5�շY����-��Fk9E�Q����+�vF1�z�^[�d[��t�p�.�Μ���?|�$�Cl8��d;=�Hi�<��:ì�|l�N��;�
��4���T�I�;�|�I:��q%J�u����}�p�/� �ƺza�Nt}��*?zVM$ˤ���l�6e�I�=a�=gY�z�*V��Ad���:��)�¡�M%a����I<�}�Y��y_�)����?nrB���h�L��ĊN��V`m&_SG�'X�SI��>����z���
�Z���J�Ow���J�g��zÌ�]��A�d�{�5~�f����@���&;���2O>縒���&�s)4���hu����L$8�e53M&Y:��=��|���AΰI�a�7��,&��q�;�8`��z^�������OR�;��>d��&��6ɶL���d�2g�k�|�$�39�H���!l�C�L&u�Mf�g�8� ������� �ձ�v��bDM<s����|�v�3)'�zk�8�Ĭ�{�d�&ߒy�L�I����	>@��m�I�|sX�C�m��ٖI���lx2#޸���
R�����o����'P;�'�|�Ԭɪi:��7���	���d���@�O�$�}ĝ`|��g��5;�|�O�����Q������������ה>���.��0�B��q$��d�VR|Ì�JΞЛI�.���I�x8��L'���$Ӵ�퓬$Ӹs:�<ϼ5��W�]�cv��q̿��:��L2i'��C�x��g�I�f�	��d�V����q���d����d�a�N���I��� >#�x�}_Z���(^�kw霻_r��z�i;>߾IXu��1��*N ��i!�M&qL0�I����ēnLXq�iX{C��d�=Ր�'s�����`u�L]m|�a�'�퍨̼���Y�>��z��M\�u#vy��\��;)G�*Lw2�n���塧K��9V�CW�̎��b�Tcj�b�ڸ#Gzć�Z�xg]u,#�	vdX4çI[n$����U�	c��77]�xz1j�z�1Fs4N�[N~��G�Y]�Y�w|s�,�3�{��x #>d�,I�~{��%ABy��q
�h)3-��6ɤ�$�N'�m�a8��Y6���hqi>}C������J[��������P��Y�|>��E��x�>o�:�a<}�q	�e�=a6�C\ϒT&wgP��J��b��d�g�m'S��n�'�v�}��ok�UgsT�kw�����2��'�|�!���`i�y�m�h�C��O�e�;�u�d�}��hfw��%ABy3�u%d�VL��q��4������X���P~���V�򟇽��D|���:�!�I]2�l$�����:���˃,�a�ӝ�:̤�=�	�4ɜw>�u#�0J��j��u�,N<?|3oWvs����zȃ�T�d�'����	�O��he�I�3=�ԕ�	��Ha�C<� �$�N\2u!�s�m'�,�(N��y����F�w��;�ǙN+����Q��i;u�'�{�M��g�@�&�3�!�S���I8�Ol4���L��Jʆ&}����L���|@$xF��J�I�V�{[�s3��(�ԕ��H,4��{�Y'<�$��N��E�o�ŇI����q��xf�^�8�>�i&Y:��W�'� ����i��E���j��#ބ��0q��)��'�Xzw�!Xi��߽��I�&{�y%Ւu��Rz��Ͱ�i=t��RHz�3M&Y:|���Yw1���o��y�2=�/N�OP�s�XM3&���N��;�M$�'�Xz� ���L�޼�$�<�^�	'��R)=~`|[�H}�}�DlWOcǓ�ݜ��XN�M�����d�Hu&�\�ROP�n�O'�ѭ�u'YY�X8��M�$�y�>@�'{�6�i�����#${�D����:���u.��3%�R����}�O<>�%�W�����m���3)����Z��y�
\\��l(�m��cyj� �&b�T$�=\u�֦V���j�U�_6:�:��-��4蝶9jJ�R�����p�`T�N��W[2 gC��
����;��ֿ$P�|��-��2���a��;�x��L��4�:�35a6Ì<1�L�OY�N�a=���{��#�{G�>���q㊸�+���3=n��������|&�!>C�Y>O>fqgM�Sɛ ��>�u��(��i8�ĩ�l:��t�6��M�w�	�h���ѳ����u��������}�#�p�߽}>���"=��d��$>�3�8�d���b�|�|���|�S3� ��|͇u�����i8�ĩ�l�8����:���~���1�2o�o~�4�|á�`�N�a=�بI��OC�Ĝ`|��=�N�>�1%d��C�m&�Z�6�S����maěe`{�{�u���7py���ݝ
��M�ggl��C��o�'���:��l'>���M�vwx%I6�'�ϒVd3�`��h,3i��M%&�q�׼��X��k�7�۫�s\���6�>z��'�����:���=5`u��<�>v�xɓ�`�'�P�';`m&Y8}߼%a8�C]ϒT'��!Y6������Z�//w�����o��=	>d�t�d�a�e��8�͇̝ՐP�&�e�����0:�{�x������OY6�)���M�)3���Y'�{����̸�+�8w�������PP������*N��u&�4�0XN2|�3C�d�O�|��d<՜@�M?0�,0=C|l�H�q'S,� �����x{���7��WZ~�_m�	�$�� �M!ӝ��*T�;�IRm���N�m�O�|��@�<����m���ԕ�!�8�������6��h��f'�[3ko�s��,�����!P��g��N��&q��e�u����%J�ww�+'=�>1I�M�|��P�`m<��˦� i����ܕps�M��?B(���Y�YZ`)��{W���;-�b�b�V8Wv`V�)8twS��bQ�mĸt��k*i�.����aBŚ�-�;p������z�l驠F����
l�6�s�����S��Ӵ;�p�H����Q����
��aSU-F\_������G�=C���$I��g�F	����N��2w��C�� �=�T�d�w��e�u�����+�$��"ɿl�Rq�i=t�Bq��ߺ��=�b"hڹ����ˡ���=�>>L�uM^2Jʇ��PY%Ow�d�=�ԜI�*�!Rz��~��,'��縒��N��)=~`y���y�<���&�[X��?x" �=�O��Ï�)�4�>Bq'��:���I�C[�PY%M�:�	���z��>eC�}��>d���ͤ� s_{���{4w�~��twY��>^��0�'O{��z�̶`i�������0��I��>C�N �ROP�sx�L�M3[�Y:�	��ԝd��GfMvγ_�}�o}��Gޣ�|����>����6��2sX�I���2�z��ϔ:��Oݡ�'Y3�Hu��.MP�I�<��8�d�����k=Rt�����*?
>�>j>�>��'C=��>I������03;�|&�!>g��"�����,�$�*e �L}C��Adߴ�IĝeL��Fn�C���{\u�d����'H|��I�����L��a�N2q������'R|�]�u�<�8$���|���0��2&4�b�d�!��Ad����8��?78�.{��G�dA�}�I�N��}�d��]��a��1:���Ou�8�O̞󸓬��w�q	ԇ-2�m�����OS~�����'p��ݗz�[S�g�� 2>Xm<d�9��:����&�q���8��{���'�3;�N�������ӶON�����g���*N�"���|Dџ��Y�q)?y �ȀO���C��L��N$�a���mC��r�l�8ɶN�C�Y2q�=�;I<d��`�O��<}9�@�'����ߙ_��[*�iU�����S�Xd�;�ݜY�^=�cB��3������o�m2[}������y�+W�z��a\ʼ�?'9��BwJ���x�ԧ_@����]��s��Bӓ�-a��2�ޠ,�p2c���a������\]�j7oS���}�q����z'��'P��A`�u&�z�`��I��f�i�	�T>d�CP�8ɴ��!��� u�N�x�xɮ��}���6ػ�M���3�;����8�H���`�i�N�8�m��|%ABgvu
ɴ���q&�i���O3a���g�͇�4�S��������|tm�uݽ�R�ǅD�>&�;�`�fY>a��hN!�'��|�u���$�XO;���iY*m��)��	�O��l:��}�m����?��6�6f9���G�� ��Z�)�3�jft6�}��U!�=��^ہf��|�����{��{y����/"'�>F���ټ�0�����ם���%D��?>f�z��gM�Ȥ��ɁV��lo�+Ms�NWN���U6�'
�y���VXۨ}yr�@�j�[�>��L�ն�l�Vnu0��o$'j�h䇷�Iaɡ�m��*����5Jy~�*L��sY~�rz �IYkw�j�w�sbh�m���UjΣ�fƿ-IJ
�O<���e��Z��학�����c7�a���ՔV��<k| ���E]m�����P����˓�w\tt��=��W�o8����{�l��w�\��y\l�N�v�Q��0���o�i[���;)�'5�(��P��j�f'Nf�\9WW���/r�Y���7L��4�cR��ZM�z�Yc��,��j�Z�Kޭ1w�{+�%��@|���/ټr=r�DS�{_o'0ƃU-�
\�����+���,�\��OL�D��c�}����h�T�qˊ��(.�2���wیV�:WerZ)�Z���Q�E����S�L�n=�+�����c��� �-���uc���̰�0�n	��6�՝��L���Α�1=F�I�Vծˎ�[�`9
��ׂ|��\�̠
����JA3W�����up�NS�<�ݾ��np²�bd][0V�y�oL�{fY��73��Z��0��n�i�h�S��:�W*}�v������$tӔ�����(L��n�Jq�3t�6%��A�Ą��J܃���b�����h����AoR[�"�H���� �R<ڥ��Me���WR���Ga������	�]:�����7��朗��ۘn�سܲa�]c���lQ3�7�E�<�j��d\h-yJ�Tq�[A�N��:�P�4@�Y�r[�6m�k3Z�{۰V�$K�p+�;2��*/��*��PW������j7�>$nW�,����266�JVo>�c_[E�b�[iMIm��gpi8Z \�x۲�fZ%�Vݺ[����]�ӸR�J��%����w<M�K*]ά��r��Yx����hz�����e�)�Nixieh��l�e
�f8��2k�kƌӒ�Q#h���]�v���x�Ś�Y��v��ꁔm�s"u��D�5^Џ���̕�LEffU�bi�qB'V:�۝R��{�rw��u�r�o�g�r��R��I]�w�����-k�n$sQR�
��fvq�;өcR���j9x��J��]e�*쬵�ab�-�Z���!�u�c�(F�����%�EK�q��}�-9E�b��R��*u�d4N�����`ұ�{�	�R���ۻ�Ҭe�Q/��8(�-r�2����hմw����t��#�I��RW�	��@o��ygN��^]p�Jz(n�I����W�g$��c�o!Ի6�ν�Q�X7��e��,���ƫ�����ùÈ MP��_p�ةB��fJ�銺�r�oXE�;�����H8q#9kU����v���z�0�b.3�ql@��f�s!CK�yH��T)N[
W��r�M�no#׺+ 6���[�}9i\$:A�����ΧܶV�:�+Ubp4�qu.=ً��gj�q�VF�b�|����Ay��y�+2�t&f*��t�pҸ� �`Lt��m��V��L�ٕ�c�n;��Z=��h�
���m����<����趇g	M�s�Z�ޯuk(�(V�YX��`�6�V-��-ZթZ!R��ō�%-km��*H�Z�b����E"����[E�Z�[J�֥%j֊�4�e��R�cF��k%��Q*TkjZ"�mEm(Ո�+DP�Q���`��K�B�X�TKKmX�m
�l(ŕ��H�U��RЫ��6��T�D��D`�)YQE�"�ѩXT�D�EB���Z�Tm��Z5�DA�EU�-l�DEIiQ�J-�X�ֶ��U���K-��Ҳ�UA��XT�
����QPZP�[J���b*�+�)F��4D�(�ckKl�b#X�THڵEkb(�mcXT ��Rִ��[)*��+Em��j[j��0�*��*#���UE*X����e���Dm�F��(�E��d��0X�1kD�AH�V�X��+EQD�Fъ"Km�%2[B�TH�IZ�ň�j�+R)R�#mZ֔�lhM�[{��Tz��N�W���]C��
|���J�z:�x�$��[w�[��xp�5�\�4j�ŭn�eU����x{���c7�W4����`�x���Rr�{����ov�^Pۍ��\VWzr�[u]i���b��3|��g{9O-�Y����N�� Mf\�Z��{�G=���Ϗ-�t�\�s����ĕ�|>Zx`�K�n�[�\�]=ӝI�h����(Dr���偉HW�Ii֊���ky�].Z}`&w���q�_I�C3|�����ܼTN6��yE��Q��X|���Е�̀몼��1Q���]���3�:���A%����01��w��%ϡ�x� RƱ%�OaӀ�%7;i�y�:��i�.S���\r}���Kΰ���q迪O5�+���\�i�x��N��,Ѕ�5+ns�����ܢX�${F)�3�zdT2gmCt�R�r�u�]����+npO9X�^c����[qh�Kwy�w�iw�u�2չS�I(�t������~^�\�`�����p�N�`��oU\���RN;T��7��+DR�z���]�we��j{gm���a��ˤz�M�2b��e��	R#�zg����V�S�j��������ʞ��M�5c�3�hr!��`�6�t!u�W5M^\�{Ա�K�n���wh�$�ōz����ݭ6G$=��k;(^׋�˕q�:�d,��MV��6�1*��b��k��L��Zl'���w�sbh9Y�qD)=r��;�'��T�J~�LW���7�͚x�nRݦ󵕷zis��8ؽ�\��ı�5Ѭ21��t�^���Dr��M��>��/��X�ފ�=M�5���ꭌ~6t�9H@�lU�F�����#�'(��sN<��hd�ioe7ڦ֨�p�ڈ�R�Rg�F�k���W�1�И}�WA�As}j+KͿ>Z�α҄P��*#�K����9�j1�K�J����KLqJձ�J�٤�+|y+�|zm�T���&��}v7�lr�̓�VϦ�5�l�˰1�
���O�޽*��D1�Ӯ�w�d
��C*� W�H���9��f��gƃ����ym8M\����d#{kk��E�^$d" ���)�i��-~��{��6�o)v̭d�|���GҔNc�y�mn��m����"���]wj�<���ۚ�vc�}D�8?{����Z�x�cjM����9`�*k^Q]{c�:�]b_;��}X����3Q�{����3��dM6xסv�)�"��yC�+6���je���vV+�um�9�EQ�I`'�ptgbjj����\��U�%�Xo��y�n��N��|��i���VK�U��=+�qI�����Y��$�IO�z"}��)*a��4m7t�fݞt!u�Q�����ɮW��Ԟaֻ˝ш�����A�Zl4q�L�f�=;usL���N������+˕r+�]�N��޾L�n֛�=ެB�Z�V��T�o#r��ÓA1�E�mʏNKv;e
�R:��sd�r��Z3wcw��X�>[��-�^E	jEt�B�C9g�9܍ھ�Zͦ��a6��}��1�ݧ�ѷ�;P�ϩ��C8v]���D`�z��rDv�T���5�T5�xT����{�������EG����EA��7)��
z=8w�!kv���z5]���3�ۤ��&�v�nҊJ 2p^� Ǣ﷠��0�a;�<xɝ�f�{��\��B��Y��(��Y+�`O����§ö�
Z~|�n��'�O{��~
�'o�<wo�c��)�cS���Ja>������-�k֜��������Ƽ�y��:�w�g�{�_]��y���~��o��Ĥ+{4|�>=�~|s���n���՞.gl4��X``�0�������s�K�W�5)�JV6��G)e=�t��nj��1]W�y�%�P�_e��]*�]׊���Jdh��/��9v�;�h��z���/��SbWUy�������O'�'��i��%�����n�9��1*Q���=��l�S��:n�T�Ã3�:�5:]���>�[���4{Q�1�wB�࢞�ftPm�rRN���5:��Ӌ,>�C#]�jɾ�<�q��ͬ����X�b�eh��Hۃ���Px�E�q^��wD��,�����Ub��u���@��a���.\*nÐb�۽�2e�l�*9��qk��j&b�Z��;@��ǒ��B^�-�`�����ۈ-PMN���L�P��&Dѓ]����������q��wu�h8��X9%�����H�=�͡�F��77N��ݣ:����xxxu;�)ku�"2�g�Xq[�!VV5B�]xdg0o*^n���8j:a���7K�SRj��J�M��O��������yyr�k)�͔�\���9�P��J��c^����yku=�k:^���C6��ȡ-c�������1�Y�ӭ�jPku��s��.~���F�y�}��6|�ç������s��ٳUѝ�
�����{z�[�^�ym�ہ�ݿ*�Q34�����˹\ɛɫ] ݬkt����#��R%y(��[a`��Fy�)�s�#dn�1��:��S
��6�Ɯ)��LH�2�㶥Db�^d���Y�g/���@\��i}���ҽ,s2��<���k�H�q@�&
��"�O��Z���.3�Ԍ]���V�܃��Gwu�Ϩf��o,�D鞖Y,�KQeC��4k�ty���Y��u�����I}Ȟ��Pd�_������EX���r`|/e�A��0�|&�����K�f.er�������q1�ELI�w�[J�����1�͍�,\�T�eY��w�j{!�/%��w�MG�q�{Res�Ҙg�U*�.��"�+n�o:�ThbR.N��\����.3v����lم��p��[ֈ�8�8��4�ۚ���QQ���&��쯗5�?y�!נs�%��R���t�<�E�w/��\��vVM>2Apb�)��U�d�<1���犀���pT��������kA��B/9ݪ��K�𩹼R.��A����/(5��ۊ�������\U�ΡO�csǺo2��sN�[�����PX�Y�Q�!��Y,K:+|��]�Ws�^8oٳ�V)w�𔲪йr'��K�:�5ؕ���r������,��u��V�����ǳ���{���,��R�j�Ho�lFo	�9[˸Ga���C��n0�.�*MƂ�^H���f�����CkrUVS�Wz^��@�Ю��eQ���<~^���o�كz�����j�S-rz*���,�Y�Zk��XdG��csdz��B����@�>�ӹ���o��vߋ�R��=1�&f�idyz�^��x���q��f����]��x��M��o�{�%g�,�ȫ�*w^�1[�{������N�`�ΔTX�E����f���������<پ�y���}Ε&�Ch"���@s>$'��J=̀�uOe����f½{��Eĭ�@�#��E��W�j-�w��=�)�ݙ�ݧ��x���{x�ZV5����}�Wq�'h�yN�@[ �x+����{�5X*�im�1u~r�a���,�q���C��Ĳ�JT4�򔫝Q���s�4�G�z�I8-���(��Q~R�>1���Q������T=�%�"�K;Qos�k7;��Y你�]ÂC�'['�C~�B,>2:���P�L&��G*c�|�e߲o3�yO�.1���HkC�.���S�{�*T�9��Y�s�		u@2y6��U�ϙ����� lC�v�$J.�TC�s�a�S��(��<�q�S������ؓ=���ٽ\��[��E|��X�ڲ�
��%��?���ff���൹��٘qs��6Y���6�qsdÂ+$���kJC�q�7S���B��N��6��$����L[���ѾXFAs��4΋�q��wf|�Ţ�w��J�V��z���5�xQ��4�������~�UO�ڄ&;��7%.Z,	8Dixg�c8}��aT�F눩2��~�ҲN�`g=Mh�w�R�Żk�7Ȓ��	�� ,IW���G�m�^�(�J˕�����X��o
Ja^d�0����>�۹MF���d׹���}�K2��}��R���ϸ棖w���o>�m)a��Ӱ�c|D�j��%whΕ�޺�x�E[q�U� ����A�<����������d�:���*�E�g�J=62�����9�{��PJ/�Dx�����xZx� ���^,�NɊ2H�S��k���V�M�3��9�9��5��6�_U�7�僅�0*��Ǵ�+�`���,ir�f�f�����ӳ�l���0�Xj�ŬQB����&�fΉ���\ܡ�x�����-kJ���*�uIr��T�E�([T�1xS�;�����kX�eu�C�e�A*��NJ�:���yY�Fd XP�\��L�G=���g�"��g�ʮ���\��l��Jz�ݧZ�u��t�q�Q�qp�ZgcˢqMBq��Z2
㚼dXa��]�jd�lz\/G�s�q��@L�����Ȯ�~lK��	슦�ac�a�|�>1ٳ\�c������2��Z�<'_U��yL��	+�4LOb�T#r�dX�(������o�޸3�GZ�L����j�!L)�o^��5��"GL�z(P�[ָ�mO+R��^��ʇ����ɒ��g�����\.�qz��t���>��K#������/+�C%�lx�P5�@�&U�7;�F���Tv�NAI݌���N�~��ی�ް/x�{n,�����u���ʳW@��ݴ5O���N����t�W{}$��:���=��W�L��H��,G3�c-���.=�h�X�a���@�s%Yɥ��9�_�_}U_W��n$�'�V��Ӌ�:V8����q�N�gG��"2��{ԬUq���Ǡ~��mK��ݔ<v	�e1�Nd��1�c�JM`�#U�RÄ�I/{�����;&vU$[R���J�L��Qe��������JD`2%hwOa�m:��sح��R����ڂ��חܦ�2�f�DW��,�n	X3�:�CΉ�1A�[�v�3&$�Ʃ')���Td�(Od_��9�O���P;6Ϭ�`- !囲=��P�Z��`�jJ�ڋ+b-��%��6���MIΞ!��ɦF^�UVX�I՛�U-�V�eڍ������>�Pn�'������D3�|M�ٓ����*���Bt��YOZ��Z��>8F����˱��I�s�u`��e��{�� ��oNh�����*��v�����`*|���Z< u���O*���y��v�<uǞ;�չ����.u���H�ӳ�C?g�Xڹ@�t�o�y(��h-�D��1�w^���.��4<#o�s4`>����Ǉ-t��J�ZL)�c��(�K�e��=�a�zϵ�u-/�ݓC�V�K�a����u�.�qN�Wcn�Ŵk�j�C�h��IR��K���D�ب���;��6C�wh�q�R�
�ˡ]��&�{�� =�[�ó���n���ݷy��
mE�8B��05�`�jTER��i��`�]�d�x���<rXpQ�ܧh�������αR�0�:����<�H��Í�]Z���on�`�ݥ�8��#��޶l(f�����c'����frZ��P qX����N�\�V��ܙ��)Wk�	d[��P���f������~�����ߏ{G "S�]��{3�N�/�}򣢕SЪ?�o�2|;5esH�\�L��r(��P�����Ƚ�v0l�觑z�wM�Z<������W�A*jz#�͛�Y����p=���Ë�z�zR��98'q9���R��$��a|��*Wv�:Ǫ�q���Ҫ��}xu_��ה�c�Z���̧h�6�F�q�����X��]�ќu���^��P*:��
�׋&�p(%�b�|��\�����~V��^��v" �Ŭ����J�^x�泾�!��{�}���*�^o����Z�sG�e�gD^#�X=Fֿ��z�����R�"�d�l���.��lWt�ra���\T�cL���40�[�z�.��h�Y������n\��#]�-���Y��hQߊU$^-5�=�����K6܋����N�ۉ�Y:dtjrg+�J�6�.gt�C���nk�QY㏑
8���]�KZ�{�H,ŝ�y�|�ͫ1w{5���+w�)6��x!�.{��_pr�Cl>x��2��O�l�m�*!/�!�洛������{s"��J2��i�M	�N/���#���2ཨ{d�j�V@"�A�Ѝ�b�&��!�W)���1F����jTttk �G+x��o\�Y�:�V�TU�A�W��I��@���jm�"�T��c(����ĳn��%,dk2r�r�l|�喷��B�Uu�f;�\���N\eG�ϟkZ,��ux�[��E�`#k�mL~=#�1]#�8ag�h[)�b��>7f��ڂ�f�RYI��7d��� K����!�zNӸ2�Z��F�v��6�N�w[8K��t� 
�d�p�3s��ܫ��0�j�R�x)2.���a����=�R�x���\��`�Y!���ю��s�t�J�I���>��=,'ϥ�Z+6�l�3D8_[čm�>����#i"�쒦��TXfϸN�R��ֻ4onU�,�F�x���;w)��[b�ed=6�*KT�:�{�YIڮK�Z��
 ��}t3	������h����ĸ	���J=�O�M��veZ0ȷ��e����9���v�4�L�]La�wV�6Ѻ�G�:�њВ�R*�΀={���-���\���L��*RfN�ܘv�VN���"|�ep��t�c&a�R�I�Oh^�^�7�݋[�h+>J��LV���B�`kR�[X�ӥʃH���9�������'Z1�;n�t���qa=�k�	��u)�n��[� 7��V��k���
4�����G�N�{&�e�>��F(�y�d{-�k��X*U�Lr�����j�j����t�zH�%��pS��&U�h�ɻ��1� � �����Xq���v�K�8˩QD�l޴r�_I�8B���N�l$ܲ� �u9�Z�S&�����nIX-4.	���G��'f�&�s��2���Fѽڠ'ya���5U����xk�2[)I(j��5��î�?,��kr麙��J�am.�u�;��#��k[�\��Ot�V%�T��b�g;�9l��\�l=j�U*T��_i���E��Jѫ+�|k�$�n�g淼V��v�sp,,�PҔ���*ܘ͠�/�Y
�O{��t���\�vf�(Y\;]���Z]f���>� ��:�k�j����Z��6u�]�
b�6�Л=�7�gk�R���)1^�q�����e�W%�Z�t��݇&,�k�����6��Z�jkg�YI���@y���y���;��Ρ�s���Ň�+bR�ҭ�*X�؅B��AZ�E%���`�l��Q[E�"��Bڊ�"�1��Y+
���#l����XѶ��J��*���B֨��e��%)TPX���*�QZ�dA���KV�֌����Qb�-Q�V��QV��5�"-e��2������Kl*m`��J����QPUkX԰m(��R�%j�mX����m
V�Tl�j��PR�Da[mm�YcZ���jJ�TQciX�eX#�AE���V�l���bĥ�R �e���)�DUU�Z�T��R�mJ��+�e��V��"�5iT�VV�k*
Z�j�`�m�A�ն�*��P�ե�*������E�2�(T��Ub+-i[[m(�ԫ+A�(��H�6�DE���T�j�iPTIT��2,�Z�Yee��j�"�)+
�%�-eE�j��QF"�`�-j��-K
�E*�UQ[ZTU�Yw�}�?m�;�z@an�Q�{͚o
�<H<���;fj�Z��$�[�A!˗lbQ�un��Ne���c;g�� ��𝆈����b\+?��C�^쾏�U���@Ƿ9ĺedZ��Xp�7�l�}~�s:���D���^M��e'P���^��yO���2#`ex��D_���U>��8.���jX��Cnu�N��>�3V���ȱsiAL1XUc���L@oٲ�F�.�7z�Z�$rY�/;w{#v�J�t�y,�c���:�;�v�W�H老:�yҊ�$Ȑ��˹EWob�̼5*<�O��xؙ��n\p��K�lJ��ʭklR��?�����i�mL^x�,-�x/���C����4S�f�R�c�>Ϳ>�uFy��7�ψ�|&���x�UA��|=ssd�_	�i
��%�Яx�7�C2sc�q�,�x�/ό��n�yhm�n�Wo��in5'������Jd���P��Nʐ�`��]�h�,��0�����B�Ks����R�E^�g��R�ؑ(��\��0�)���H�s� =�n��٧�����Wga�R�b/9�F!�X��-��ZcQ(oV�_^f�����߈E��{�9ƵR5�wN���U,�!���֯!�z'w^#Ze Mf�KpV	\����\;��)ۼ��m�j�Μ���wo�,գ:Snv$�͢1;^u�Ҡ���C�h*u��^�m�x��M�ؓ=��F�#tŜ���-��ꪡ��W�Q��k�'h�|=�H�VŊs�.��n+$������S��ǡ�-n�f���y�ʥ�6k��5�P��M�^3��\a�R�Cau��0����;����]y����3;��l匰=X�?�(eU1�P�;��ȗ,#G2�C.�F[�~�W�["���«�z�4�%��W~�G�����,�씒�쁄��b��WJ�Q�qw߂I����9�ݿU�o�v�iJ�݊n��M���/�t�S�8I5�ST����G^��HV�Y��t��}��2�&l�����Jr�o6�0o��jZ{�=����Ԙ]�˨X��6�(n�'<y�W�}�*��sb.Flߦ�"@��X���Hx��+�
�9��K�q�s�S�L�[��ޛ/�xmys �e=�v2D�(���sy\�0?=��׮�O�D�w���˧��g��3���6��6,�)�W��}Ӻ������@��@pxo��5/�~Ӿ�j��+�hy	���9�[TU��S��~�X�$}����tܝ��˺0��1����h_d��ƴcv���8~���rx��f���?�o�a��Y��Gk�����˨�Q7;/y��A�Ŭ�=|`�|Xr̝tvgA\N��h�\��Hd�4�BT�_U}��}d����}=x)Y�2аﳲ��Qq�����/��"곞�5W��{�1�G�����顝)�$N��r�Eh�k��k��PU�('V�\
*
��m��p��4�G-��;y.�!��	8]�(P�b�5�Ĺy�Z��.%�T�py���@�7�t�:o[7�.�|nԴ4���d���&��T	��{��h�J�s��)ŎV��E���_��9��4ΛnF�����r�ٱ]a�#(y�kR��.�BP͂��;X�G(�0�E�� Tld�zV�gB��ϺS8/�����	�꼼�x.־l���B�!��Y�S�ML��N˗#C������`ؒ�	p׻�'/.����у}wc|g�J�u��iĸ�4����+" ����G�����v/�^-�sђ��$�"o�I�b�y�!ָK�spU3���F��<�4�3k�*�6=ؽ�ٜ	ҦG������g�+���أa�;bړ�7��ɦFg��D�8��mV�]�n�V��UЛ:�f�@���S<�t�7YP7�1d+ח����˂������6�P1�K�E�R�L;�y��%�'�����\k��'r���Ϥ�G)q�뺶q�GB!�G�I�hr��O�6�2�d�[c`��F�+�]�y?  <u����1(Q�8��\�QŃf�K�Or��t�>�2V�Ԛ�5Gzj]�#!��3�N���x��h�JP�:+��T���f)e�Px��襳���8{�G��:6�s^p�����Ī}�g%�+$�����N�I�dqU<���S������ӳ��P���xN-F�(����7�!hF�1^}����w
0w)������]�J�Q�{f���jwSW�!�s��q���"-M��������p��j$�C�%�շ�Qt�bcZ�A�2�T��"��͗�l���$x8�r��c$T�V��1��;j��ם�z�(��g���2t'#z-3<����vhW�Q���=���䧰Z�ܛ(pg�$"�W"����Y�<�te��4'C��2�㢯�����{~d�vѾt{��9L�Q<&��F
O��+}k>&��G����Ӟy"���ۆ�èY��]���z��7�!�s7ցb�h�V*WJ�r	R*v#�͛ꑛ`t;g�[�M��ưڑ�GM�b�{
�N����\u��k8��Q�ܽ��4��[���uڝ%MQ]��$*E�VE��J4�e�]���v(��V��&��lṬ�M���Vڤ�^�Ra�6.�M�lF��{�UR���Y� =� �g>V�4(vAi��T��Kd�u��p��yA����D�40���YͥV�I[GhnkS��Č;-S�/��[���P��"̚&��+�ڱ�o�>yP��ռ{WOV��Ō�|%y�숉�]�7�`.C]��Q8��e�muBGn�P�V\�Jnn�27q6G��5���W��627nE�R	�BD`�v����
��[���n��'�����Fu����;d/Xw��r�C�����Ya]'�ʇ��{������y�������=��+�g�4�~MJ�,��S�Ƭ2#y^1�͑���
vr4�'x�毞�=ա��qx�ޏf�t*�.����<l7���Y�3��E.�B��^���qԤ,���}ӡ��	�6w�:ld�@6  Dzq�By]$�ެ~��f�?zl�0ia�B]2́��YO�dj�L���y�_��v��3֊�=s���_��ձr��3�n"O(�c+�4
},ڗH��>��'h����3n]C����Bj�P37��u�(�ۍ��xW�;�䙲�l�ܬ���Sˍ˥
�[2� ��,�j�en�wGǛ��l*TԌ��	�`D�q�\���l�G����b2F���;��Iu�\����v1簑n˛М/$º�˻*ڳ VY� <���f�;[�GT}�38U��#��+��vӵ���m�:-�0�?w��x\�AZ9�ׂ=�ɢ�G�M7T�����3]񋽋�j���5�6S8s,�Tn+�_h��f�F���5J�͚�P��f(4у�j:�¬:1u�Ϲ�=���O��c��t�ly�i,�{ಕ���9<#"6V��L�u��a�$Ұ������=��?9�8��)�!����(�ʻ%��6 �O��t��M��4s���e�8�zY�I�lK|~�u�&u�<7|�9����"����%Q�9���{9�7�4 iV�%F��T�P����r���2��T#;��ܔ�h�#G���z8�P��ș�����W��
�(�����^��.���׽*d���
�w1`I\q ��;�i��C�"�p�z�D횫�j�]���L�n�Y㹓N/�]NɈ�pұYn֩�ԛ�Ha+���t����TdQ���R�C	q�.���gF`��u1[��^ٽ�Sl+k��G�gj�V�+&E8�RH�R�{αW�fH#p�˨�P���-��k��^)�+�2U���݌����k��0.���:·����Hnu�ޖ+|�W�P�|�2*䢼��6���ap����s����7��H�a������G����{��	�p�v�ђ����\r��bsǭ�Y����7'�\�ٹ�����W[vz1.{y{[�#�dfCXfV�k��b��s�{Ϟ��$צ�X�Ň�yJ����x8�ft��Q�B�8<b��9,����|8A�����vێ��
��=��o3&�j�A���GOe�M�	6t�cÇa���?i��(7�5�����Ղv��J\��Q�k���V���+i��W	oΣ��Hu�T�x`��{��������ת�Ϋ��-l�9���h�ĄvD,uQ:-��Xv�F����r���t��W{�7;��a5l�o���#{+�Lh��@�"�p/��zD��ڎ%����x���Ԓ5)C�J�.�|�*��f��5�KCK�x�]�h����������+k�u�=\�P��2_Sر
Y������)è�~�hٹV)�ـlR��h��\kC�$���Z�$����*��Mb�1�d�s�gB��Δ�������g�V��ax�d'狈|�d�e�u��9"M�v�&6jڸ�"F�ʻ�+�^���6'��H��ƶ�)���7t����Zp�B�>�S�<QժS����8��]8݉:bZ����:��q�+C��
�!4��7��U�x���ۅ�Z�f U��m�%�BG���I��,`�V�uS�8\�����`��(Ĭw�ݿϙsH?58h}�ݏ��eDG��!+"Ĺ��E ӵ�ϼ�c�H��ױ=ʧщ8���'(A���r2�5�rNSyV,y���BVE�r�nz��4.+�<ӑ>u���w���c�V/T�X���ؕ��_L����Ö.umZPL�9Jռ�/}Gm�ݘd�X�碌�����������|w�8i�钶���q�[������s�).]����@Kf�JQ��ڦ�idqs��ʋ�Ŀ���w5h֙�t�a�'��/6���J�y�Zm]aO��+��;�,����SAN��RN�1('���
�i	;QYñ���/M�����חV��A���B��T�_�\B��d����t��ܬ��n�K��Vvaĵ�1������
���Xӄ#��K��������gu���L�iq�G�s��N��l)}h�0�T��V�^�G��(]c$T;R�|��0���5�[�v@�C͋}��SV�}���ؐ�:�M�b��%�e�,l4;E����Z�Q��ɷ*h:[��|i*r�k�996wme*��Y����lu��E�+]�u+����ԅ�:��ݘk��u�G%�B���B�����z/�bV��������6����kB{��u�1K/s�L��L�9�i���IF��:c؈�Z�1)�˼�r(�.�f��ۂwZ߳�'���s_��cmI�Z|��x��*��_���k>̥���H#�Mhd�1��1֙av��Ql���p��2�������w�α�~IVӿ'� ׽i�b\���z�r	R*v���'�nR{p��kǻ�Þnr����փo��a�'[I6�(��o����N�h\��l7Kk{tJ�:����5)�{#�W�M83��R�%Q��Y,?���+��j�m��E��Cٵ=}�[��.x���jDD��mě�S0$5ض"}�������,���Ż�p��wgG籶����'Jw}l�F�ȿc�L��(E�l�w�_��:_\�w����n\��뇪7#H�.|Q��o՟4-�8g��@{��d1���$��RѬ�ī�o��z|瀗���;r,���(o�ؘx��yN+ՆDl�����ej�w�`��WWV���8H��.�e�l��[�s�ݓ�O�]��F�玉�F�ُ�T)��5�)6�4��h�&�����v���Q��n��QrWY�ȥۡŔ�^���p���ۃ�0�|fm
e�8��u��]�Ф�n] �+/�m�ᵕK��{� Lm�r��[Tv����������/rvb��FH��j0^�6��9oN�#o�ԡ}�-��\��9��-��Kݔ�F�4ٗ�����P4��+{ۛwh]��WVO_Ri�@�����EЕL�{Q�6:k�Z�C����tq8sEV�������iHe�����J�����$Tj��\Q��K6��/Lz�Bv���;�f�D�B�a��Ƥ�F�!��~Ip��]�NЯ�����,O����E�0�T�\�]��21�Wp����ȟ	�Q����k�]�X>�ښ��\w�
���%'^��6����������Ԩ��J;bD����֑e����pR�+��Ei���{��Pz�=�Q���o8�ۥqn,�� �J�`�!B_�x\6���9ɸ�E-�ЪEdz�����FY�Ÿ���(��ɇVI�5�#��wi����hR1f�,��)��6e荌Q�w����ɹ��l4΋�8��v!���G��Ɨb��>:Ẃ��n晷�vԃ����q��2�)������v�܋SB4KR��P[ޛ�GZǕ�.�wY�)>M�T*��:y����X@�3���{�;'b֥;5�Фx�3�
��-�p���7������{�(�D�lI�]l�9��j|���<{G��erY<��g ��r�$c�]% *8/M��("���B���4@"��e��0-h��������%�j�:ͱ`Ӻ�N�+���Nh�/��K5��T�^h�2�R��h:�m��-�Y�b�Բ�
۝t�u��p�Z]7�7���.�ŎZ�B����t�*�5w�����V�����6\6tP�㽱����XN�|sp����ˡ�:�-����K�;#mm��5vp����fU��ݩI���αֆ�w��7��;��F�Lo��݂�x��n��շ���2r�7k�_������Z�q�Z�4C5љ�*ɭooE>�9w]�[�G��#]�Z,*Xo���d��LEuH4�O*w0cm��v���������s���� ��[u-r��F���,cƲ��}�4��ݶ$�ӭWQ��a�y`�������[z&;k�&�Ux�̖q���U��S^i�f��+x��&���h�l��C�l1�EdHtS��"\�]|H��eN��PzfP֐�h��uQ}�����hz§[b�{���P�}fH,�m9�yj-k>�3 ]\C���tA�NjtC)u0���>����f�E����Y��ÎW&�N�ʄJ�^��,�ٙ�zL{e�%}���7'N�)�|�T�3X��c��`8����;
]�F��N-ȩ���εqe�n�=F�k��>I��8ݝ6��bV��϶��}A��P����:�m����S8s'�8�J���D��oٍ���[�Kϕ,�:��#M!�u]���v�g�E���Z-r�F���.oj��t���>�I/�{\:�y��¥]S��gzΊɢ��q���tD�X�&�t#�����n�bڵ�-�0��_��kK����7���0a��ef6+!Ȼ�*��Ι(w[qd5�cj�Ѿ�tE��f������
IGu^��й�5�h��@w'�C�K2��A��]Gnt�f\;n�fs��j�m,�u)�U j���t��(b�z�(��x��`_��%�X��B�L�9r=��-C7{�l:0^��s�Mvʤ�����y&�Yi]q��]��g�|��zK���]��,��^�� )z�Q�|O,[t��h��u1#�}�P�+��4�=�o=Ffe��x"�t�]]�͘����ڋ���A7�:�C7BE�BQ��ɦ�ՃR�D��k�%X�b���Є�#*�w<�襤����v�EΩ�7[�Y��6�whޱy�J�9�^K��Jr�Պ�"ŐPF
L�iA���k`���DX����U*�EPPh �E��A����"�EQb��U�«KDH�DQV�Q��eVQbAQQm�����ʩJ"�b��QV1+X��#Z!QA��F*���D*����ҨV�UT�� ���
������(�V��ETm�-���lmQ�KXJ�1",X���F[UkZ�EAV(�X��b,�����[VeP�1E�U��P+X��"��A�X�*����"�
V�Pb�Z�*���EQEQaQ��6����[E�T��X�����,QE�V����)DU�1�QAF*�"*V*�AE��"��Dcl
���D+��E�+�F1Q�E �ied(ʅ�*"(T�`Ҷ�V)
���dDX��-��ķ}��;���!�Y�6�tS.�!Or�gM\�W�8�uk�R�T�	�lYw(M}Uo�� uV),���lLH;�P����Z�������*��#�kV�j�yu/�P�1�C*��ڄ0;��ȗ,��4p����ݗ7�e�@M�Z#|<���l����]�>�P�JIP�@�c���=�Wݘw�;'A���a��J}�G���GZV��O����v������U��Z*��4�;�9�:l�]�}��Hcz�aS��ͽ���2�&l�>��Rp��FH�����=�0����}�Т�p�5���ۑ�����Z���:,U�G\؋��6�{wP�Ӕ����"��S6x�Q��N�SԮ0��յL��U�v3��qj�P����8v�d[���c9�Μ��{1\j����d��\h�j���]�͗Oc�Y�RϮ!\��u�N!>��f),w'��Z^��˔O�ڄ�-i�*ǔ5˱0v���R�W~�5	�o�e�=Ք��P���j[啴�_ԫL�c�ֽ	�*�o�GVf.1�~cgE�-�&�XL��ƌ�V��f��=A�Oi��ڦ����{t9����ʚ�l�7��n9&C��Ϲ�kr�!q�Ô`}�ʷ)ׯx����h�S���=�-S���1�˜.�Ң�ɱB-!\�jߔ��w��͉%���p���:��zu�L��{�B�k6AWE��e⌮��R��(_A"r�t�*����D�={���������i�yΖ�k���`��r�{Pv�]�D0� K�B�n�w)��C�)I��p��͇/ɕ�֠[P���}&��nd�_�q�
Z}�h�}F{E݄Ϧ�:K;6gP�>�T��4/z(q��C]㘌P��|d�0�ҥ�r�v��ÿ
]��Rں
��՝%Y����n��E�*W��3�����T�j�cJq'��꜏�W�{��_��9b��;���爚Je�g�Uma�����tw�
�e�|�f^�2߁�l�Fܬ��m�'��R�o���o䠥�.�3�;V��!�o#[臤���||�w8Y�!�$�DܗLM�V���w����p��}Oۆ��{sv��Z�wq���]k��GE�zX��ĮsDT��ZÔ45':oWb�ë:�r2ev��ޞ͉�-�۰���,P��8k�ʜE��H�gN�}:d�y�2jH�N2s�דx��絜�H�z�ʅ���8t�8d�es�����Fpmf½��J�ag=�r<*����7oN�nb���-ɺ��nWjX�er��P��.�e/���98�`u�jc���d�ΰ��{)U������t��jm>�V�SR@G���<�y*)�3j�0���*`��T='w�.�پ���޺�X�'k��m��8hv�ī�G�׊߲1A�H��I�-<��UaJ|�L�>�D����vf��.Wl0QJ;c�\{��6Y�91p�i�W�3�Wg�NuN��w��w�G%D�Z��D��C͔�3ڪ���V0��}B�Ko��2�>jU�ܼ\^ܝ�������.�Yt�,�R�����ޜH��*�D"0Vdu�+
��4��iJ!�ꡖ�(��(����4�T��oGy3<�����Yc\H5ᕽ=������wQı
��y����+-Z[�y{�ꅉ��f���c�h:�Q��u�p��p��ح��t��#\���W��S�C��5�6�pmOp���J-6��n6=���2���-=�f�2������~��D&הt��Y�":M�{5[ғ��t�-k7n�_,J��v��@T���Eaζ�l/���Wvl�{'J%4�%�!>��3�� �sմ�P�yTBw�F�P�£dC)`:u��H�q�F1�L�q�i�2[O�����O����n�f��&�5�c���W,�6h���h�o��p���rQ<���n�Ň��˓J<1�]݂.}��e�+����ܽ�kWK���V#Rpe�F�jL\4vuξYʺ�`�Q�+w(�����*~�ګ#q��mN�����i��>���}����5جl�q�VY���6�g��dK(�#"�˝�ܛ�q�#]�q�.���t,zP&�����!�#��\&�oIXt<�y�����,�>�dY�k3��e{慿s�nV5�^"��0��s�J-G�]��Jj9]�ջ$�9�'�������d'(�aJ�,�u��S�Ƭ2#y^3��9%'6>�\þ��o���G!B���E��{Xf���:; ����O��c�3}����X�J��}�rN�>��ả|�<���O�]������w�:/֨CBt���@捲:Zu��}�{A<U�߱�*/i@J�Y���YO�dj�β��'n-��K׶je`]�5(�G��R�ܕ��/�f�+�4S�f�	�7�}{i�:�^M���f)�Z���o�F|l�&�IA�i
��X����q}��b���s]�6MZ�ܕ��FAc�V�U�z��~Q���P�+��1|��Cm�e�����[�.6�[LO9��;6`?�^����yq��R������I��zs%W���{8�`�iG�t��-�Rހy�G�kZU�����7>W+wi�#S#�i��z��,���l�Z�Ipj�k�ӭ��]2��C(G؂�o���/}3:�)<��� ��W	�O����:MM�W:�����R�8�*Pyڃ��
�z��U{W�.(-�-�q(��Ҙs�=[�7��+W�9�P��EbN���Э3��K��t������4�̕������8}��:lȞ+W��a��E�|�8����S�u��v�蘿z���?a�o�ŀd�!�ڄm�ɹ��l	�����7^��J,�q!���nzJ9l_R���r�X)n���q��U�'9|����G��\7�7��r�Vw8�yt͒����Z�+��_[!`���,����־~�R~��e��w(e��:g�צ^�2ǁ�z��]���e�Ba8}@h��Ҩ-<�x�dӇ���n����;��}d���$9-��������w&Z�͞6(C�"���pz�"U��N�t.iq
�5 ���ꇘ[�����3�fBq�x5�=o���[tu�ۭꉬ3+:Nlte&��x:��"}S(Z�7'OP�Z�<�p�y���^k�����R�읮�=�1f�p�%-�Cը\g��P6t���C7HQt0]d�B�`�"����m��O��.�s���a��6�-XG�eM����i�ۼO��u^��*�����c=62M�v�#�VR�譽oL��@]M��
X8�9B��ir�}�U|D�g�ͅ�^�s�R���
��Ů1:���޻�e���8E���:������¥��F&���x�O`��]&8�rNz�Y&�q�#2�`$4n������f��9!������an4�U5���{I�oȮ�~u�BC���E�R{��BI�JQ��g��E�闽8FF�4C:�TB�њ��.��0�ky|��ɕwco������#/�(�6�ѺO�I岵�A��%�8�	=���W&�[}��A�:�o���.�غ��9]��٬��wxױY�y���C1U����'�dYVW�H]/��W��.���Y���C��\���-'^��bXjd�f�f�H]��Q0#Z���FLy�f��������N��	�z$��6ݛy����6̓�l ׾��LJ1P�R�I��#�:��S�ㆎ�q�7칫�2���^����.D��|j���"0$���]؃��P�G��^\5�7+/	�s5{RVA�!>U6�%��ګ���ǌao&��뫕6�g��Y��߮d��ԭcy#��stbi��,�����XUZ����޼{2�1W�+���(�U���s�/[+/���M4���,l�&�bc2+��Ӡ�Q_./3�K�s&~��Rw����EdA����3~�4���D��n�Ҳ� <	Y�G5Ì�֥���k!.cs���Ż��K<C��_��,�Y�J�j����(�Ӷ�p��Ӯ�R�qzt.�˵p�fˤ^�z� �u��5����X���R��ĸ�xi��;' ��ΰ���13��������1}�Y��`������v7a�����Xr�YNW=n{�Wm�7�;���٪���S�3����)�����8����K#��ێ����O.j��IR�v�#��..(�5�n];(=�l�a=�5��N��E�ԍ��OP�]�� C{agD��1��v�3�j��|�a�e,t�du5�F+��œ^�Bl/��Dc�\vS-�Y�/��l���q7YP��={�2�dK�����X�D�]�#���P���e�[Sʺ��C�]��G�������c^���o�%�´�h!��[HM����O���)�o=2]`���f$1\�~n�r�5�k{����Gq�-�X=��X��g�eY�5�Œݭ� E�`�6K3�e��3��ݫ����Q �On^�v�6����as~�N.o�л٨�,���T�{�C	��<��k�ww2:��g8��Tow��� �M��Ws���{�M#z�]�k�����_����d�З�Y�A蒚1�^���+=�I��X�?$�E��蠯^\i��\������T_5���}ٸ"�&5W_y���{��!�*�Ox��pƃ�ʄ0�t��C>���WR���:�Ex�Z�Z���=È~�h/�1��������!��.��lB�hW�3Kb:��\��kGGR�J�FF�ޞ/�^8o�e"(_PJ���Q��3l��<�A͚,�]�^(�/����j�Β����{���Y�0y�w��~Y�B�($�_�0��v\�2�S:�����cfUؾ�}3x�F�z�gM�g�=&�lg�gB9^�w��v���������s�}�[����C�X��*���ע�l�z�
�����S�xuiqn<�0�=A�.���9;Bd��TFXήF��}ѩ�Q`���bn=�́�+e��^s����tfMD�=����䑫��at�~�E�uF�Ý�,=T���i��'�8���7H[ܢ�r�)��P���J)��Ni��T3)��T���7}VUq�tbv���+0;;X���iP�F&ͣ���I)��;���V�Eӄ3Gd2T������4M�����MuG�5� �K���,��RSs:��6��<3�a5��.�g�yd�Q���7��i�ϣxT~B@��@�Δ\^�.�*��8:]6���������U2�����;3�}sv4l�N���Up��K�P�2�(��Y�
},��dp|g�ݩ���,��^����ix�^8lyy�ϒ�zm%��B��8B��a������YEC�ۧL)x˛���v(�Zp�M����tp*�b�A�i*�4�1w�j�	��Bw�$��]�a�傮��)��y\��$����IQ.Ԯ8��0]sP��d���m��S5��⬄_��\,
��n{����=��\}j����@�<�z��ܭ�3Q>ϒ�k�Y�Oeb���x��p��/�o��:ᣇ�^���f6L=�G-|2��zX�~��ي�2��;���w ^�:w�F�+��m�g34xX�Y��i�oV�ݍ�i�B�f,��z���J�V�cז;�.��I9�º�o�;"*fw?���7�y�ri�9���n���i)w2����ܗ�%�������� �ur�q]��,���D�Ǩͭ�Z'](�i��5�+Uc��O�����8{�+R���+X��7�)��᎝��$�I��<dÆ�r�5[޾%f��I���Zc�'8�[M�*�V���ѩx�o.�QO��b��6�I��b��r��}���o.���"pheJ��v	�h:��;u�=P]�"��˥PZ���(f<,��y��Q��IXS�;����C��aS��{{B�{q�D oca�>9A�����]:�Ý�N���WC�٣�?P��	�Y���#259��֬l>ދ]Fh����xxZ�'��+=�9Raͩu�%�#!Y<UOS�Þ<��P����+�[c�e�fك3���y�^��:��.^�O��:,ϒ����*T�T���8���}�&y]��e���N���E#��v�V�$'M���g�n��n���/U�R��q��BO�����[�^�eJ�K�'�����֊}s
P����sU��(Lӟ(��k�Y�$,{�彛C���DbL<'�v��������E��^��`bAՐ�$�2��8��+�K��'��v�0�T8f��Aq��夺�^��	3_:�>X3��<�o�����wp�ᐁ���Lp�K�^cI\�BbD���]Ṕ.VAp�_ ��� �ї���N����$p�}��o�B��=�+L+��JoqsE3n�:b96#a:�ά�Fv�o�}Htͼ�eT=�[b�*�-����.fy�j�8�l�v��[���G�%4;�0�t�gXh�;`�%�X\��J2а:>��5M4M]�`�&u1�6�˭ggL�Y��R�Q�(���p�Nˤ�nb.�d��ڸ��*�@z$�F�w>�;�~*�f��c~�ח�p�z��b��(8�%�P��ެ�VJ�N$����;g��H>����1Z��f�lŨ��n������s�C�HQZ6�i+f6o�n�׭��R2;+���.ճy��&nf����q���u7���mҀ�7*m����"�CE���)ffK��{�^�l�`N.��+���\�: ��ԫ�+k @v�3b�R�l�g���	�/園�u��\(�T�o0t4+�}v�Ɔ�{:�Lٻ�P�˂s�6�5z~�wjp펹ڃ*��>7du���Y�BOG�Z��y��C�\J\=.�+�0�gV�Jͬ��:U�j,��:+wv]�;��@�;�gsr+���nQ`R�w�&���b�U��Vr*��B��ᇲ�'��*�gfk+!X�\Xفl��f����YccH��,�DV"xujv���w)��7L���Ws֑ˏ�� '��̓p�]&)�Y\8ə&��C]D^g,U����泘�����-��)��2Sx��R�s��ɋ;����Y����o;�kAwH���-�n�4ͻP�v�]K�5��FP���ބ��~���8����x��}+=٦rAӚ�1'�Vr��LٷW+,��D�\�%˺T#����;zD@[S�ZсRoa���2�=��Øe��כ���SpՂ
yڮA51�k�&���#��Ad�w��ɔ7��P��6�}�ڹ2���N�¸�gL���0e�6���u���D�biQ��D1YbU�q^���-ɕ�;JI�قve�W����Z��j�ݡI�(e*��m��l�
�8�����)�8�yK�b��D�(��Ŭ.�وR�tS�崷E�)�C�e��:�w2��z�]�bc��Ί�����Tճ��m�t�D�:A�u����J�X�;W����I&5֪m���$��f�ij��mc�5.�J�l��x���i��Y)�2(v���<'@Ok4+*�f��u�H@� ���Gzv�h��B�vw0enF��T����e/�#�_S�iLD�8��y��2�S�N�]��*�1��P���Qͺ�0Z{/���/dW���΄�.8B��7�/A�&�Ȼ ��t�h9L��زwko�',533FT[�PGY �O&b�]i�Wr�P�&� G[�n&E�X�Kw6E���	���SU����0��a�:���].n���<k���;&-�����<ZB���ܠ�T��B��nR[*�k))_b�	� ���}yb��+R��,��eJ6�UPR#Q#Z��A-��l����jư���J�"-m�b�@QQ+R#Z�YR�QjQV%)Q�J��VZPh��եKmh��E-(��k(�+DD�Ե�ATIU
ZQR*"�,X(
��+*����"��X��F��X)m�(��նP[eJQ�V���X�U��+Q-T��E���EAU(�ȣ��)�����*"��()(�1m
+�$m���Q��b*
��AV1�""��Em(��E-�m*��DFШ�**���(*��F#��*�ih�F��PX�*���Dl-*�EU�DU#Q�J���+ATb,-(�����Ec�l���Y`��`֊����HƵ��aD�*�}�I `��+ra(���Sr�M��a�S2!��^���29�+uu%��]�r�T{x�;�Ֆ-��ԃ�J;��US׃p�<e�s��B��?������P؝����W���ʡ��6�q�.]�Ԃ"�gMh��[��ҳ���Գ)����3��PV"�R;"٠��gJ/:yS��˜�+���I��s^a���,&��C��\��ƶ
[I3�#�1R��Uq�g�_�Qe�	�ˋ	Wya�����i�3�N؉��%"0$���]؞=撖hug s�-���M�'u���ͧ��q����^F��^:fOpJ�D�pM�sA�VTd�(J�}Y��Ln��1M�%�:/}M����Aa����`+����푓�Eg�+�"�^Xe�w�����s�3'^��G��� z�1��,^݄o#*��1���Ü��p{��l$Nx�`z��/���r��ܴ �smr1����YN׃�o�.�4�+�"�.uC8u��#'tc��V�>J	���5��a���Zy�\l+�)�����oՆ]��ZڍEx_{V��t��S�ϱ@p�[�\�9��׆�Vt�7�e�\��u�甬_���-x��)fs*��t�<1�_lX�&U��A�oHze�������m(��p��Eh/J�=lWo*͂��iv�6w��oI�e�֑5��/��7�QΙ�fbPt:�v��(d�]G3-5�M�u*�N+6����� 6�'����U(%tj��l�$G-��tJ{#*|�n1��]��ӵt�3�M�b8���L����ԫ	:����q��e�#�*��/zZ�u�5�����U7�����u>�`J��H��۪~�]C��=��4�uѴ�r����_��üy�t�̜���}�e�eD�W$���CT���T��r�����ˬ�[�Ow�3����^�ζ����a�$���*��o�2`��$�	��V�&o����,�ma�>����kZߤ��_�=h�H�[R����j{�Q�Y�?l�����{�I]d��s���A���_��P�h7�j0�X�֒��]J���mOU�(�{�fΣ�d���@{kԥ�w����X� �1.��J�d<��u4p�_"�v��پք�>����1��$V�A*}r*7��`.C]��}�fq��C<d��s�6o��EC~ˋ`�fJ/�w���n܋�9"�
C����H{�q⃗��|�6e��v+烓3�>�٦�VM�\ L?EZ�v��s۪/�U�:�1Yio/Lqm���b�m�3�J�;6�98�כk�2V_d�R�Vj���M�Ke;s5�d��E&;у"��;ۭ�lj�q�gP��EiOo��j���zܜk-A:�������<`�Z�q�<Z:֗�����TºM}�e^�r�(,��W��j�!���Zs�:#i���m�}��'bP�b��gθ��qI�q���\*��eC�P�vT�[�.��#,�l����4')@UӅ�N�Qඖ�a���Q�ǽs��=���t6飠�l���.�;���t����L~Y.E�j���1ݯ���"��7niZ|��
GE	��`�t����.��w�.�MS����ewr:�޺�0槯��U.^\`r�eBY�Q+;˖���zmCat}���fh��Ƕ�^�U}t�m�P�%�r���K�鿒Py+��P��pHy����m�����gs�yz���9M+O��&�ėj+\��`�{���-�g�в��v[�׼�`�'5��:}�7{�*�J�)���W7�IC%�E�t)\r�W���7�v�����ͅ;N}U����Y�����(��I�7�Z��;ҁx=��,&gn��Ւ�o�j��
�`̙w�A%���9M˃U��������u(9�ܛ�EY[��LLW�j�K�`�#���)Fb�3��ب������S��Ĝ��\���roa��A��Ľ����l�nt&E�c����� E�������;��Y��9��)_^j�7��'�2'�����n���V�3��B|N�.�x!R�Վ�c�1�j/�bc%aéCg�E������<c��C"d@����=�8#f���'I�i}��V)C����x�Z�+}(eU>ڄhFl��j�����e�5�΢���-Z.F����w�JY�$Y`9k��L`]县�Y��y+�G��>�8���;8IA��X�_�R�lG�Km�=传�'n4	S�ː����M��N��$��e�ާ����d���{�$�$��W�R���m�bL���<�b܅�q�����t-)��p�����g���S^�@G8'g7pl=����k��~�Un �D�19:�1+T�]�.FlĆF
ʤ��p��*���a�v(�����18�[��n�wy���I5���V���W�U�;���R�Y�|m}О������K�[��o����hd��0�{p<�}�j��n��Z^�+�w4��%���T+T�Vߡ�tΝB�mWm�c�C�E�RUF¡Oo�^�g��[Ě��J��
���+8����-�IYwllf9��2�Cv����I��L�����G^f,���f��z��%�wżL�.�9��휺��=ӻq�>U��N�3��rRyLA�>�N��k��^���-�蛈�&7�\=o�	��>o�F���_R�rt�=�U0����4`>R�y����AՐʈQ�RWEC�冡�ob����iN�=�Q�K��u�PV]V(#��������D�m^Lh팗h|�Ҭ��Vʉz�X�*:F�Ǣ��"BT.���+"�Q�]L�<�tn��f��5�R��8����H����+I`�,�s�$�8�6'���^�������DM#1�'$��wmf�.�a��p1���������o䠬E��*�c�j��\fm7��ir��:ӓV���v[5��N�vx�K}���,8l)m$�Ď���+«�4ώ�c	�B5b�#d��D�)�����v�&�7%"0%LVK�u�J����<v��Z`��[��v�ˠ�g��>��"�>�u�V���bC\I{$���<+*2̶,��ڷ�W`�d��y�����x?��e�a��sT�Fl�M���%bsD?�Jy�F�A���9тy�d���7�l��l�t=���v�A�fB�t^+���+;N9���@�	D�:ܒ�]w��г���%E�3��]O�qs5�����lQ|���h*]��ط���i�d�������M��"��,N��%��X+2)�7�%�1ﳴm��C9�/4M22���F�FT!~��K�g*qQK�.�M{-�Ǻwy!]�n�t�|x!�sm�r����;^�z�à!�)GXn���j���"�R�ia�1'��8wV_k�`E�XnmJ��uq.0�{]3V����־��cV��z��D���j�fjv�3�Jq��\b��.�x�Nʠ�1�,o��D+'�v�+`=��M��/e"9m����C�/z]�g���DR�QcM{֗{9�����y�M�2��:�{W��ը#��q��t�3U����Y�JWӏ1�:�jЙ�~�	t�#"󍎱\�/r�{q�ݶ��������lqy�x7��	��=�ޫ���/�K.��KQeC����`-�5�{�iv���	e��%��l�^I��saNPR�u��V�٠���a��j���U�bL�ⳬHnݻK��6�ph�]A���Sz��[.�;.�Չ01��OZ�F�%u+�X�P˕�dgA-aY^WW�q56|��!�c(��͓T+>�驝9 ��ʽ�9 lغѨ����qe�Gi��1k�}��F��s��}
�&m���8%���\3���f�s���!�`�ט�>�-+�vjL��a�Pr���vMf�ʱ�7wy0J�*%���{+iC����J�ܨC
0�Im$3��_$���Ji�E��ӻ��8U:�]d�(X"��J�)`mw�������yr����`�k3�(}�f6�rB��_q����J:�©�k/i��l�-W�S�"�c�0!��g��O|+�7W�wҊ!{�V�tbjX�;u��E���o��"�Ȉ��
g�V�k%��:�/M����]���ÐҸ:i�N��WJ�j�Y����ַ��U�9چ55Zu������8F+!� }�~�j�z(v�G��5^ʤ��b��μ���(��o5�����V�}�4���B��zS.=���WӦ�mt���:GK�%>����{$Ⴣ^���BP�3�MPyҞ��c��s���էw��a�ep�wG-�*c���E�|�zοW���	�� !
�������r�:�<T�9Ea�1Am���T^M���`t�W�*���T4��9D���+�ό,�څ)yR^e��k'!���Z�v���4�4��v�#�����A�M�>F��z�ל�"\��ɓQÖ1J����[w��3���(L	���f^n)G�]�����?����I�����d�֢��܇�2�J�[	6�3]G��*�)�7���j�7��������q�^��p�%�F�^M�����sJp.�w����Q]��e^���UR�vKdH��M5�H|b�syp�P_�+#}3(��TS"�;��x�Jc�u�w7��W�NJ��T�{�Ex�����#�c��XTK��+�T�M�WNܥ��˱��#(�Nef�9��Zy@�Ù'����\V���=u����.���M�����%-�(c\�</k1_�Wח�����'�2'�ظ��BmWAЬ2o�����aK�ٟVIu~Fq֕N;�x/q.��F�'���+sPc5�o�I��ᙗ۰����:�d�y�G�(F�](wQ�=l���<��p��B���-������M�;�r��H���2�Caw�'���X�5�Ƹy���F�R)}�"�ė�gd>uՆN��{80�s���bW��8���l���A��Z�������8���P��rv.7s4bjA<��"��Mtc�1�jvLb�I����ck�CZ~��m�Q�CՌQfb���,mh��;�<Zc7x-%��Dj��R��Ʒ-Vr�O��}\޾G�p�m���N�F�����[l� ǈ|�������tR�l<r��maȜP��H\&<Nmi�Rn����ո�U�����3�T��$8"��3f�+*ӥ�s2��I�Ք<u��UPk���xb�0��ǶKF�y����uEd�=e|�k���!s�UE�oE����"�f�HDg�*�6F5����r׏���P�ܹ{]=��7���Dc��;���q��E�{'�ڕ�I�Q�ƥ�9����oڒ��,EF!X�{p�Vo��r��c�Y�ǖ϶�;��OK����-+�w/T$�>�C�I�Ç���͓��=�O�葘�m��s}J���#UÊ\�a�&:�\<Ry<&>u㼻�Jxq�H�g�Y2KX`��!a��+��4B-L�������[��]ʥl'1,��0��\������Y�Ə
O�����ɍ�.�wb���?T�� D%�����qQu�R��\?p�޶l9��x#=����fv�*��ZGK�zYd��h���hP؝����1Z�����$��b�ѽ�9md��M�;���,��t�v'L�eA�kR�U�z� �9p��,�q:>~�n�N�tr��_��m�9q����Ms<�ŧ�v�X2VTU� �Fо�{yk1s��dԛ�Ā�/g8�\��u�G��Ⱥ�WL!z��*�yܦ�)�h9˪^��rwm�y:���Hh�ffVtXQ��\{�IW�Җ!ZR�`:��8�o�-h�LW�K
[I�KJ�&��;��l�����컥����6zuE�=WV��o�p#��1X�kʯ��=w�8��>��*�g9�̜Î|ޑ_O��P��+��pխ."d+�86Q>bO;�����}j,�i
���l%�\�G7S8h]�F�.��p�f�{9�%�+"'���2��n'�
��y�!���oڴ텀�9�q��i���A�FT!c$c���P����Rʽvc�6�w�A�&m���8p�6��`v{.�������9�^r�z����H@���	�RVf�vF����}��e$vcu��\!>ȼ7K���^Ն��CR��gWWXS#�njf��r콸��ۖ������hdqu<��f�o�����Ӽ��f��pF�mV��%G���Y'Uc|�6Q�]<�������"Dr�D��1��v�3ڪ�;��cy�E�w˽!�$��B��]LX��U�BԸ�PˎL���͏)}h�|e���T2��r�5�;y�	Tc^Ss<�,��C{g%�-[(�뭣;y�n��l�6B�[ux��} ��q�\�b�U(P��w�����d���ִņhy�i9~C%@u:<�/6����JV�]&������5aa�6�9sb�Ԅf�m��/��� Mɼ�*[j}د�k�%I�2�:�����u�7�A43�LҒӔ�ۭ�x�SHt+t�w9>p2]�0iaV���
��ʻ_Af�T�޴�k)�I,6��o7���ң	��*?�b�Y�u"XQ2�Ք0쇧\�hta�� �i�[V�u�5<�z�o�۽� +��2\��Qa��tQ�K���';����p�;V�j�s^����$�s��[X�{�2 6hc�"]r��b5�t�O$\R��= �Ņ��-�3�+ye>L��C��\˒�*�k;;Z.G x��Gv�l��F◗��uKr���[���M�si	��z_1����|�o0_����%��V��������I���r���n���Yǝ��2J�On��c��S�&.y�yz�+\%���v�"xLFJ�E��Ҳ*v�˦��5�C�CNU����:�e�Q�ט��0�{WG:ڌ*Z��Z�O��/.���S�XU7GV��i�:�>x�sXW.����w]$�fU���E9���|��y�{��ĥY4+���)4ZK�mi���e'���yV{Dڈ^������[��㔧qy�ޖz��X:8T|�~8s8�j�+t(͡�6V������Mm��k��<;t��{y�VjG��7��Y馕K���){�U�>��&rF�Ԉ.m��Y�W!���˴gr�^ɑ�ɑŘN���N��]���ޥfm�(-A�9���<�Wh��LW�p��l�w���d̲�i4��):��򱼙�G������VHrԒ��= w�K��љ�Pk��k	f�ːMR����"W4�φ�,�41ZBQg�.�r��KI��V�ܩW��D`=�%�g�+�c�(�6�Fn�W�&f��a K��)D�]�)��TYn^�h�si��3�U�9鹒�f��x^WR��W���Y�9�~�κ�>�z��ц�B��<��i�ޚT�6�B\�|V�߳�!$�2�f�ظ�;�nC�rtsTSF�`A	�����5[O8��JU�G	`�5U�}eCCStC���q�;H�=�?=�
�R��{�klR�(�W�6'�VN���Rݡ��Eb�m�X��g�i�N^5q,��Mg@�"S��
���&�5mok]��:,ފ�-�ö�8`]�\�%��T��uz��C��%��eE{ ���:��%b ܺ�2�Cc��y%^譶�/d�ϝ�z�F�ˢ��g.B��� ���F���oY���zMc��^��&Q>�k����kkqI�&L\�d�g�+_`��!��k��#|����d��8�P�|k�I���
��(�"*�bFF
1FZ�PUF"j*�EF1X*�1F
�Ecb�P@Q�K����b�UDA`�Q%h�#��l*�B��UQEDTA"�"1E+,T�ŭB��+mb�"�Db�Q�Kb���������U��1��X,b�R1K`UElTT-Y,V"�DAEȃ��1AF��DDX�V[*���V1E_�ha,Te����SXX��U��*�R�"����YU+��-iR��)Æ�X�*Um�pV3�)�b�Rʪ�Ƴ�,b""��Z��1f-�\%J���EDŬm
��ťlE"*8�PÄ
�)�E�"�����,Q����}�X��/�+Pjѓ#��(�R{�n��ne��vD��dt�9�VJy!�w� �$�����n���v)w����6�!���FoC����"P��`� V¼�wzUtER�ݖYw�TV[��@�N9��=X󹜠�3<����k�f��ȰT:H#OHn�{�iv��燼����6�]��o����d�l[��R�\%�ɥ���r5ȃyg����w�w{vA8s�z��I8S�{�|3"ʎ���զÕ���k[�����@���䮥q���O�=���뙻�30��:#x�Y�}R��(w���C��j(F(�bOZK�ki�%���guFg�)�e��h�w�6�0=f��_.X��ׇt)���|E�^[2��5�k��6��`^�Xy!}�宪8=x��$C�f�w.EF�&`'=�6}o}Ǟ�Ǝ6�����U�x�˲ȯT<q<����Y���9E{DL��k��2��k���&Ĉz��o�\#�a�����Q�8�0���m�
�x�u���U�Ꞓ�8��`���8�����])+(C��;��� _rÅ�&�m������`
W�a3ݖ_�n�Ѷ]�n���TCS�=��ϧK�R��l���y��޷��J���U��C�a<J���ǓZ�~�P��=���mީ�6��Q뭊�h�И���^�iuI3��S87�Gw)�pڷۤ�6 ��! �6������zf��ќ�rig>��NS���#�fA9�=~�!Beǘ��w|f;5��`�(�6ն;g��؏�9�{�@YӴ�{���<�H���.����&!3�fT��2_��c�{��I׽*��	|V��֩��U(Q�Z�c:Qq~�EԪw��t0��܌n�ή�ӿL!��Չ��3}r/Ūv{��x;R�z�EW
)J��Ļ=7YH��u�Cf2��5,g6��N�!��\g���u�y��7���8�,��̨<���S��:=�I/0A��ݽ�@�zױGl?8�U�)�(��x������Ņ.��VF��E۽�鼾B��թ	H�p*:Z��B*U��;|��2!�u�=.�2(��0f7�	�G�ܟ�+�w%���߶�kR���,�ն��[�"�B�ON���+�h�g�"o���]����p!�f�])�,P�1�rP�{Y�����9�࢙��ȨYڎ����p]�j����K�\�t؊�"��֕t�V;���B�by+ڨ|t+��"P��Rd�|�s�fj�/����Q�wj�.���^���A3E��ō��6��&��[����8B�|�nJq�����4��S�
GI���|U���4kV����ᕈ.��Vɢ����y`��ֵ��]�ˣ�:�%��z�ͽ��a�w�cE��Q�a��-�P��F�q痷R�x�u�il�`����{e�S/���Cs
8'$��]ԳbTD1�H����u<^�L��$鷜Z֚����ˡ�Kޜ:�";٬P��0tIK�%ceO�=v͞�^Pj'-Q�Hf������M�Z{}x�#��N�wٓQX��)�K%1�p���a^�u,O�����ݙc/���Ŧ�f�jV@��Xϡ��īՃ���w�d[ܡ�	��!,��al��6�o8��0��F��z,Srs��\�ى��Hz.��
�-x�r�@��:�pv�fu�f�%���=��1I��m�a�Qͫ���6��+`��D.	��B:�k��LM[��H�r��t�[�Y��<�~��ߌ���X��qW(�%<�����n���.�gi�d�"㐫��PV�Z*{�#��Nߕ�EDʘXuD�g���F{���۽"����;\�b��/!^X��`>R,=2���k$�^����q���en���e`]�ya��G��*NV�P�}�Y5����Z�j��`�w��ˢtЦ���f�∬���ݵek�g[�/��|�9Fw�sG���{Ϛri�x��1����5f&0�[mᓌ�NX��ʽ�[ڻ���, ��*��F�ة\���z��ER;4lR|�`pO.��7dM
y�8�j�l�~��GllЮWP�]r$r��v\����]l���WDӗ:3�-FKW%'�vs�������t���|�h���a
��1z�+
Wl6%�7ݵ���Ϩ�4^�C�.�q��-�7�x) �0L�}�x�`�G(T��NM���-�o׶mll�ji�R�Η�N��.Ɣ�k������m$�ؑԘ�ZB�;;�����p�,xk��Ug�C-C�97�%"0��1X.�OZ ���]�Sz��$�̅{ϙ�Z=�A�(+>���c0�<����=~
��~D��5Ė6Q>��I~q�w6{_�x�]~;�`�Y%�9��p�܄j�r���tā�H5�ݓ+"�[�֗j']�{Y��:j�UK��RÔPod�z�%l^݄ldeB2F8�̕�:��}�9$A�c�#���q��*�����	��ތo+�|7�c���7~���,����gԔ���h(�2�2��Bn��go,�qu�-�sp�t����wK���%eXu^��Jٱ1�G��c<'<��;4�M��p�v��YwH�O.�� ���<q��ӭ:��q�N�=l��Ü6��
�wfLE���Չ�\̮P܃d�|����K��ʆ$�ú�ea߾�ڰ���?����a]aB�q^aDL[we���`�{S�0������o�<t����=�^^��<F�3�¸�j�.OJփ%�QΫ͙�o���<��!�)�|���Ӱ��si�T-X�糙�ף�׾xb������T2[p7�%��P��st8�~
_Z!ӵv�y!�n��du��¬��(�Q0V?�#TP�T:�F����,����%ܽ�h�ٲׯ��(NV&��[�����ˆ��
�K!���C_��7���W���a&�G$"^���f��ї��O���|i�naA���P��ѳ�Z*~�9IY�$+�b#J͜R��|��Ӟy"���[jO
�m��4y&�۽�
�͞�}��ޛ�xO|�A�4ƴ�x�پ�G{ P�`rG.����+X��-�,}����d��#��s��\\s��:��b\]�|��^�,my�)���|F��iu��Õ�#�P�M.��q��y�c��?){�]tỠ1q����Flt�zX�1^2��y��yn,txs�*nfilh s�[�ц}�X��^V�6�'����D���hX8�'v�NMĤi;S�_WR&��k0n�*�d�.&�3�Cx���Y����X}����S��n>x�/	��_�P���ְ*�'�om��Y�f�Y��sG"f�>���ڸ��`��__�Ϭ��Ϲ>�^:^�k~!��{8�Ɂ��޸�e�8�u��m��6E��h����;�5�:Y^�z�*�}��GsI�F�d��^"�����%"��-��o�ٺ���w^UY�2'�u��&b+�Ӌ+ٽ��_Y�py�p̋����z6+.�u6`=�[���QegN�����7F����l4�i3p�!�l���^��(���_Jwg0s�����t��=35��y�[+(\�5΢��m�6v�V�8�0���p!
�����ᴋ�T�s�fg�OJ������ڐ��e��-��[�{����i���5�j(i���Q&-o.G���� �ݺ�w5%Y���<n���ǯx'p�^���(�(k�%�GTFثE�L�'մ�^�M@|+��7Xd.g�ٳ�o+Mi�.i��'�E}Q��c��o�W�6x�%�(=FU~��Qzˑ���a��w*p͢�z!~���Y�L�ta*:
9ծ�[��j�$�jI����ܜ��m��;͛����Gn��\���]�U��#��p�b�m���z���t�+���ޑB�����%J�P�<�p���lMJ��4p���\;���0-��u	�z��U��{���=�`0.�r��P��ZC>um�ڔ[��X���z-ҸY��J����b����s��N+R�ص�a�צc`�gŚ��j*Ᾱ|R_[����������9zứvL0�H��֕b�j�6;W�Pྥ�����o	��#����l9��v}��!Tpo�q��]����E��+��ua�z�]�sL���쉜q�M���-���7j�&�7%.Z:Q>9���I)�h�dqƯ~�'��荷�7�ԓ�4���Hg�R��Ϥ���x�;P�*�m:�q���9�zw�~�7�k]C.�G�}�WYՒ�d�𞕅1�,���8IK}�NK�&!����З��;��T�\��d�	x��b�����,/�`�k�7���j��{Ĝ5�����ݹ�z�^`��7RB�Ed?s�=mj�F�oX��n�tߢ�gM������/�Y�)��wv%�D��b�������w��;��,��9��H��s�LE�y�a^?�3�u9ײ���N5d4��8sZ��2�=�\P���Ҋ6Gm��ks-�R�'bk�Mf��G��������7A��5� �ФT��.�Քq.�ov:�\�E�+a��#��'���+r�x7NS}\m�Qb��h��3�b([$WH@���Q6��ʎzm�C�Fßc�����l�{�{p<�}�]�7���l�7���e�x��B���zz�d�@���6Yh�ds��[R�8k����s��S}K�lN��e�{��K�n�iqO���*%�5tb��/!K`y�`>R-闽9挍]�OLSny{��톑3*�(����V�n�HܹQ�w�m�b�備��Z�̴77:�T]R󶠫���!��/�D�Uu���d\9G��g���1���뺜���\��ޢ�6�qz�H�~�,���h��#���C|�\���X�-%h��e�����y�[��5#OK�y{�͛^
F̲����J�W�_qȳ9ڻ�Z�+,';86���4lK.6ka��8��՞j�a�ҥ�11X�a�c���ؑ؊�:��̸�����V.g��p�.�eE�(e�sMTIH��S�R��+�t̰	5Z�m�
��3�~�����2��}�wՁ��5B;�6_���N)�r���3kg��Łw���8�>1ܷr��N��Sj�C=�H����{�HCmɵ�����γ;��u��[ʑ{��ܵx#Q���G�;7E�ŀ�n�f�).�g_a�kz��ufK�T8I�6�Y�(�k�������>���__��V�����&�Y�f{VR'6+�$o�^��'6���3��P��^Pf��cj�T�����xf�懱��]5�eݔ2�N����/�,��%0F���F�Zv��':o��ܚde۰��^"�u�y�~�H:=z��ɇр��a�R=,h��<ڛ�h;�cyὫ��ٗ=T�wk���I�@��Hc S�Θ��bO��pצ�^Ն���r˃�X����W,� ��N�v����w���G�$����V����!㼳�/l���.�Z�Zo������p�xG��eֽ)���"&�H�\D�-��âS��S�8�$�Nz��a��mx�a�I�)^w����xw��e�Z�C��%��n�iR�t渤��4��r;J��1ٲ�R�<��G���r��0V2El+�Wb��u�x�\�T��՗�����Q���tlICy\�[�|62x��e�%��!��[Hh�&监{v*ù�~�C���;D#P�b�-+�f���	;C��w<������l6�!P�mw�F�	��q�Ҏ;�J��g<j��'��.��j�v�6e�ڱ5��$|]�z�k���c}q|M���̙�C܎;k�r>�������Jb�^�P�=�lۚ􊾏Oyd�\W��@6��0�؎˭�bbmtW�N.�B�}�I,���T��C�<n���p;��o�����ܩV����w�)im��n�1=(�g�\�T��F�7�G{<���!�p6)�>�7O6�E�R�M���!A�g�$���n��ļ:�}f����u�*qx�����#��72�w�>m:�8�6D6��a�����S����x������6�̉Io\�xGa/j�ލټN�U����k���ș���+ƮeŇ\O��{�>�\Sv_ ��Il;�ź��$���&7z�6e�8�u�����6^#�Y�6��+�'�g3ok�Wy�m�%�s����}�]���-b�=�0��q+�����۽��C�k��ƳB�[��a����oI�U,���չ/5����{�e�2uQ�k��2��[��ܳ�{�~+��>[כ
^�0zc�L��afϩ��Q^��(�l�aҝ���=��͘�]�7 �L��]@Dh�Dȳpu�ǩ�C��
�����W��1�\�r�8�Y%֜gc�y�{8��E���gt��0;���Y1	�� 0ZF�mY��z�<c����z�pZ�m�Xj����Qm�z��!���"%9�v�Bt}��_0i�Z�kؖ�f�vb�yW�g�����6�meW+5�%-�hj�X�:�-	���T>�p{��m�����s�;D(u��ǆm��[��)��n�u����&$�<VG�^���Շ���:\9(3��P�m��]�Xf�Q�gM(�Z;\�B��'�\��L�1�F-�(�[��{q�R�G5����z*�n1͋�C$ce��
.ˊ�>����V4<$V�W����t�5�Z�Ԉb�c��>�rv��}�	�{h����R�>��9��f�w3��@h������l������Z�k��l������ţ%���5�Up^쭰�;B�(�S�2��u��;�23{;B���D�5�1�E	Vnԋk�a��Ym|��.�U��Y��Ԯ�=ӻN��!W(��%
��&nF�u��扦��Rv��!Pv:�{�.��=����MVR׬�N�/���E����,��VkLU�+[��I�J+�Ԇ�ж�^�;]o��q� �3v��[
�����!O�Z���|r���_.5��Q-�5yoI���� �Ew#�Cf64O5<ѫz�Dz��qpIr�%ε^�v낭,c^K��ʼ��S2^��伝�T��ngH��­�Cީ���@��t..��qF�:H3Բ0JpW-ٹ�A�;���{Rm�V!��9�;TWM#c��$CKq�۝K�9Z[P��*̽��t7#�ޚsvJ����	�bl�ƶ�����*�{�n��`�9�����nܕ��M$HSv��)NHG�&kc���q�-C�n*�y·ld���Tv�f��=�V�·���uqR�>�
7��M�����!糖K�]E�b\��kfѤ&�H6PYx\\=��;#�SE��hr��a?rE�V�pN���Է��\�qI�@�C�<RWg��*63���`ğ;טi�s&v���1v���);6��ewZ̩^-���o�AX�g��@��N��g[#j��P��ܬ�s�d�c��:NQU��..zf�A��"�B��u�gy4vJ�t�I������c�M�f�NGQ/`gY,u�5�Mv���� ب�z)��.��$D���V�d��%㣵�����m��+�H	��Vj���)��v;*S;]����ƻ::Taw;�k��r�m� �i�.�k����{� �G;/
P�*X��®5��-�s����Co;���jX����P��Ζ��|)wa�԰ۀL��*a\@�/&�oJ*�vTfP���a��xr��-N�Ԭd@���o]�B�{ ����#�aZ�0ű0�L8D��E҂2F0QE0�T`�b�DE[Lc���J(��ZamQb1D����e�E�J�U�V��F��k0�L*�*�b�1l�X��E",X���Q��i\!�-���� ���Qh��,�%G��QU�(����-T����TEQqj���Ì`������� ��K��������qB�\[��-�E��,�E\5�.-űFZ�Z��*"�X���Q	(�,EX\%E��(���X�D�b�Y@P�TE���-h�"*�(�0�"��*#��,U�Db�m�1L!�A�����b��"��m�,���*�b6�V+hc#0�00Q\5���ҴjU��Jʡl�+1J-k�.�X�URA�H"�~�����h]MC��!��Z*�l��(�O��9��i�Y��ʆՙ�����x��|�\���5��&��nXi�ֵ9�X�+?Q�.Eފ���1Y�Y�����WQ���j�|c�f�B�K����p�Xb�8�R,�T�;m�=β�S�_����0��(�Df\��N��O�;Mg-R<0�6�=+|��M}���Ƚ/6%F�ԡ�,��3iJ��E�ڼM��v_kB��s/LP!�Y2�X���N9E�3�H�>3�����"=^qMz�Q/��/$����]�]T]����O<�! +��V)S�4p�����#�
z��QP�!8�旱��oT���Ġ6�qˡ\c\԰*��'���5�2�o!E��I�6���gD}��Nk�n�'<M��WS~��"��z�=��(Wk��>���jW׷\�����!��]�k�$����/{P����ad�籭*�.Վ�lN.��x?�#�z��[J2�*]����68���=�.�F&f��YڗvL'��}#|��;��5�^7A��qz�bl�m��dr�}x9�q�X�l������ܔ�h���/�-�6�4O�� *ǇoK�QF�����cY̖3�7��t�2�A�_����6��sj�PB���J�$7�꣛�����;kI�u��;�BZM�
��#j���<x(�t� �,�k[���hj�nÜ���j܈��D�)];�F	�u�nN��1��5���ybyg�Yܔ��d&;�������9�ئ��MQ�6Ґ�i��^�hT%IϏQ3�E�P�ߪ8=�q_�aO��d�=�C�Io��W����oؔ�BH�{6����Xv7��&l�>��
5�@ʆ��l�B��B9�8s��pr���m=�-Ƥ���e��w�֬m��X�n�����:&�"~��?z.	x�ckznnT��ԩYq�%
"�J#'��d0�Wb�a�bX4�W�U��B�|�&�vnߛ�Ƒ��v\��H���/!�(�+�}�ʮ�ߛ�r{��국h���u�ʁ�~��՞Ҥ���I.֖�_�9�	���ʞƱ�@j0�
�A���B1%��	���th�G4�P�1��I<��Q�HY��X��@�|�Xze�K}��S�殤�#�[��Wo}�C�n�*D�2��xD|�c�2�J*�;4o7�'2Z�>;�����?('�M�{Pzƻ�Pp��XK�z�
�[ָ���+���̆ߍ��3-E}g4[���*5���[l��(�\����`�$�J���8�urg���`�7W��%�.2s�j�d�&���L��*V�:@�xɘ�ᆸ_L�q�ڴ�	����J�eL�^0�.�`;��Fe���kD�t���.�ۘ��9�"vtX����aG���)��s[0>�p�	o���y#����R$�w�
�C�ii�!e��3]�j�C��)�t�j�����o'�*X�8�Q4�5�]W�[�'��9;up����Fa�A׮z6k�V�ͯq��[9ҥ�q���Xp�R�J��۶8�|؛}��ي�-)Y\E?��ƙ��,�Ǻ��X;��䔈�dS���r=�}���gZ{�
U�u��<��|��kJ
Ϭ�0VY�߲R*�5�iquC&�J������&�����̘�K���7�aaYQ��/(3r���l�x�ϰ�h9f�Ad�Λ��龄+�G�d�L+'4Dǌ3�a�r7��%{<8B���k�-�\v�Ǵ'=�{�9h�	C�1�A�cs�J�c��T8p��xɥ��&���$����8ݓĩ{�2���Y]�B�<�p��p�� \��{*������zn/j�`M��Tcx�����2�vp�I�����KҎ��Ӄy:Y&�8�ʬf�Oa�)�i��h��+ 5����x<3(8�pѯ)�8�+�y+��:�=f��<�vyN>��aƋ�&<��L���;=�yef�~2��<#�;�l�U�캙p��s{#�W��mՄ��$�\]�������yi�"�4�c'J���	Sn"��s���˧g�5�\��\�Ԉ��R%eq{\a<��s�齺�{gu�'2�%�p��1jmE�>،ى�U xе."��,���X��y�kS�56��ࣥ�)�8��ޜK<�	��,�R��/�`� VÏ����������9���B��H�\Y��uѴ�r�|g�o�2x�K.��KQ>A=Zv�<(�R��/��&e�߄�[�q�dfJ��o[6פWJ�ֻ&���[@ܓ
�H �&�iU��.�$�~�B�^I(����-��<o��H��x� ׼�k�=�Ig�{e�^�;M�1I%Yf��y�	�^Pm�^��5�k��=0�w���4�����3{-��\Nu�n�P��� 
�={	�����9�b�`�C}�b>��^���2�����z�逻66���v��Y43+#����S(���OЌ�n�wo���N�O>��>~�F}0$5؍�h�����p���0Q�ɒ����S;8���z</;�L�+����S<�9~��^���&�Ț�*�qf���K؜�Q�tf����RS���r���i����3�h�5)��Y���z! ݮ�:W}�z��'DN��)�����X6%G�����X�w�ڻ�x�8��;'N6���dTIUyv8�k�+�,M��0�f2�bp�~���6.�:W���X�
�|֟;Ϳ�V5�dx{ a1{��)x@Wn�ݶ���~�s�5ʅ��K�N}������uƞS�x�.#`l�u檈��فa�;�w]�W��zϺ9��P�V�ǃn*
�׶mcnr`^�<������ѳo��Ԟ	ә鮭��n�ƨ�݀�T�N�sǹ=�����8N̍�#"\��k�J���b��Z��
���z�<5)��i�t�m�Oc�[�{�;�m<qx;i.g��\)�J��T<�V9�֔�ʺ[Ϧ�Cp�X�e��K%9셥}y:\9~�tJ�E�C^Jg�z cq��۩�W�:�#k�:�P#�,��BP��Q��>1�zbεu
]J�
6:ra�ܷ��� �/b�e�b�b\�eQ����$y�N8��1�å���~�H��nxwOω{S�����o�J?�F}t�
��]gr��=����e��޾�+m䘙(�gdA�T�����6z�w�D5��n�h��u_�\ݝJ�9quq�A�M%�;�Aue�}J�Xy���,��j=p�e5�>�s�F]�Q�n�rO�-�+\��ђ�{�T˳+�����dF��y�cq���q�{����HUvvb�+�q`�^�@�&���3�ڥ�֡>�n�>_^�omL�`�h_��M�C����lqa����鿁�'b��v>��&Y$x��*�.Վ�v���}w}%�s(p�	����a6К�=�:lt�8{]>��Q��C:�d�.�ц��R�r�c���x��5%.P�F-ML���X��[O҆US����Ĕ�h�ѓ�GU��4�W*^V�	pk�{��=��0��^�뎱w�:ǫ2W�D��d&s��#�T�����Wϥ���/^o@M�+,�=��������T�F�&�X�:cS�cqS$��o�쎹ǳf��vT�K��}&Z�̓���J��G�"�N[�xb�2�&ɏ�ܮ����E$�Rj	��%pl-���9��Ղ���\��E�͛�ҧ��q^Q���LQP���I8�.��wsǜ8�������d7��y�Qb���7g"61�Sr����(>}��!�{#��Q��'��86]=��Y�ǖ϶«�-۩:�T���D5Ím���$r;p�$��qj�w��3U��Ђ�hu�[�������h5f�����J�XhDm�Q=3��UԲ���S�LM=�3��v�\e�����*h�7�>��=Z�+�Z�ұ���Nh��4�a�e���t���)u]Ŭ�E�Ӻ��������I�q�#29�L-��)y�J:�q�c��m��w3��uʝ�|����i�}�j�&8�������z2�w
�>����D��I�U���\�_��
�vD<�%��ؼ����5���{��}Mt��z��\��¾4]4�	�ӯ&v��2�@��/�H�^��o��dd����}�k��`M%]-��j�>a�+�b��e�\^�䎗��}{$�8�B��s�6T�Q�8m�kC�C�'���z��v/�����j�����נ<�lة��ٖQ4Ƶ-�����Y6ؙ�ʭx�Gd�1�)ޚW=5��ޕ.F&j����N�؇BYY����s�r�zJ�d��G�R��&��>:���(e�s�&�2$G���x�5s|>O��z=�"ME��h���S�.������Dy��K4FÌb�z���F���ZI�RNSyV VTd�	Y.Q��
p����,_�֢p] ⻕�k ���-O��=6�A�`ʘ���ڹkv.�|��ncWl��u��L6�O��K>ӑ����Gg���j���蟬���;p���%+=D���u7��:������A����p��M��]�+{�R)Vp�ڰQ��,�Y�%:�&^Xf�a�
��$��6i���8��w\�@.;���;���̋�Ac�=ɌPȼO{u��>^4?r�������F7����J;��Ly��ڤ�K�p��
�f@^F��d�QAs��,���Yݎ��؋ڰ�	]KvK�O,ofM���T�qCj�
�P��8����KZy��~�i�)�lm�8��v'{�#��9M�/��I~�<Y�<lR�
�J��֩7��C�DLr�ϦLHH�є�V�����!�7O���g�¼�E���l�R�J�Ko����D���!���SW �9Bc�ڃ4e���)}h��/zp5,��5���}��jL8���������˓|^%ú�&�k��U�o�������%�тv��w��[�����c�_jJB��"=U�ܯ�T�ȡ���fÚ����k�H��u �d�v��ݓt;���Ldc�ع��\d*5��:�x�nu��N�g}��+mx�"k���6�0��U�ۼ{�4��{u�VITv�)�n��Gէu��i	Ĩ>Ül�t����^��,i��
���lX��5 i?^g��.����׫G_�*>��Tr�q�w��d�N��[����/&u���H�Ӑ9Q�Am��Y�V��R���Ϙ�y�J��fc{.�n�����GnD��r	R*v#E����Q�����.3�؋Գ��Ŝ�����Ez$HI:����k�wT߇<ZL�+"�}���ea�
�-��\��H���kcxr4��>�Q�!���aͅ�/R���p�c׎��v~�U�F@��U�ݚ%A#L���$�%��l��6�A�sw��#�ȯ���u��T�<Q�g����)�w`=^,�������`nˀ��)���2/��/�����a���a�S��B�XW��6����jc��d+�q-W��*��ۯ5���{ ҸO=�9� ������	@{R��<�4S�r�^��t̺%�u�!ڻX���k�����u����Ct&r�~�|���ZF�L�Q��Ec6[�{(�b��=�q�֊��i5F��=��K�nx�`O�q����c �H�
FE	��8i#�����F1[�P�Ga��R��3����~mS����w�4�OZ��&�kT���e�_!�{��g+��A�����С�wIqP;�Ɗ8��]J!���ҷ['���ɖs�"M{P �]b�3�rnڢus}m7`��/%����Xe��þ���Q�Z+F��!��a�2r���V��s���i[���8�+���/r��B�\b��HX��8؊�n^R,�>�l)t�1�f�N���i�]C��;i���q�V��[ʥ�bfp���	��=���%叮���X|g��}/��^�.�<xd�5��O^�\��X0M6���T�b\�a���B��X��O��'���L���{z���މ�W�H���=˒�`R���k�z%¬?�]gr��=8��<��"�/=�.nsX{`Ib�K4�ڥqałg�
����g�J?�B|��'1�t�kNNu�T�^T��xS<l��\|n�Ɇ�H{)iYK�c��q��_T��j���D�ᰜ>�N�6:e<�K�����~�;R��f�Y�,�:�"��dV���Md�-;�՚�{S'O02�ü�8�l���du�nbJ\�X4p�-�8�[��U���]-UdĲ��k�V9�9k����X�,��>�%��Lw1r`���Fl����cw&�R��ss���̻b��p˪��'��x�x� �*-��<�d�>	>�z3�+oh��(��,yܨX��	V�enc��Hڥ�qr@�(�@����L��*v\�aȸ.��[����_!G����Մ���@>�Z/U��gC-@E��Y�A�ʊλ��5a��V��%bR���a܋ffCB�\����k�F��B&6b�k`lU����Ol�Y��M��m��!���꓎T�|����:I���I��������}W�V�X6�j����%�`��e��Re�w��ޚ�$�T��k'���Q��
R��%�,w�p��S@�h��%Yo��pO�ũ��ʐ�Q�Inc\�r9$��t2d�sN��͗�q2c��&B�^�~+�K"�)�(M��H��bv��eZ��JG8Ժ��f�iľ�i�N���;U26�{�DP:H�y����<�ժ
m�4��,�.����t�t
}x�L�v~��2/{���Eۊ6x�ԬSv�r]�fP�NXr����Ub�e�vf��V��Y�W�pf%0�g���k�e��n]粰����u�����\H�Ӟବ�P0�K�7+n���1c��H:6�L3&L�Y�����l����Yx��S��s�J�|��W�1���l�hG��M֥sG'(Q�gb���VՃyN�K�BB�`Yx�)ӏ���}m�*��,:��$M� ڏ���X��ɀ3�����v�SU(;�EsCk�J��.��.�N9��2d�ٙ� ,�m���E�EG15�5]�9b�|!vY�t�
�&a�w�Z�	�':r�i�B��,����*�Q�b�11�! _���Ō������}�X�\M�!.�髢�NYצ,	Ph�9��K��ہ�<����W!,�@�>��*A�2�*��`m�1뼽�*��VR�O��8�َ� �Es.��Ud1G���������K2�¦蕆�2��q>�[�����͟f<�c�dP
6(���\��zm���^�ⳁT��蔏+HV�n;����K����D�ϕ��B �\��m.;�y�ve�	仒�_Q�𸆖�Q�b{u��,]�#������$���-B;{��E�b�zF��9���dIes�8,�=,��2�� �ˢ���b�r��(�P�M�v7P�$��{\͸v�/T�їIF��`��n��6e9قQ:-�T�CܷZf2-��t��X`٧u7N��f�\��1g���t�:g�P/q�A�(r�>�N;:縰c�t1��uc�n�챈�Ŭ�}��f�/W�e�*��{��en��E7�(�⭚"��Z���(f)��n:w9M$�<R0w\ᙠ�����X0�V��y�Ƅ�v���ַo%Ea��s��ţR)box�>��;
�**D��b��[�ܗ���V�{H�,�8ʇ��j��[�7�����b�c���@B'��d�,�FF���}�4�tx��X�7nԳ����̻1�X�`r�U���`�(���+�q�8q�1kD-%b���Ķ�"�)hV*F(�����m����iQ��51[p�(������"���Db�`�J���0�,DEb��1�����б�Q�S��
�QAqh���
�
�U�1Q�-��QaZ�.D0���������YX"-mh�T�T+Q&��	Q����,b0UUQQUb����m%#���ږ�Qm�U`���V��-B��T-�A0�UX��**��T��8�DEUm(��*�UTQEEPTb�a��ūTn
4Ū(�����8k�[K�
�XҨ�e�UTF*�AT���"�����QX�Z��,�(�kEV#Z�0�0����TF���*1���m�����>�q�m��>]E�|w��1�n/�3�u�P�隷�Ir���K��:xN<t�`�x	��O{�_��ՠ�\���)7d��W[����>αM�FE(���`�D(�3�o��ĭ�|v�w���j4O
�\��.A8hgr�/nFd'u ֬m��X���O��x����BE�����U����,���r׏�آN�8Fy���^�^���ÿkt���u��]�S��K�8�wN"�'өR���Ug!�?t:�]��[.��(����t�Yvb�i�t#��{0��wB����������VxH���H�jWE�>�R�a�U��W@�+zN=��Bz���uq�iD�]"�yy7�^��YL7�	3�u�J�(��)ͥ|R�.OR��Ԟb�l�9���h�ă�!��QWFl���0j�򂰍�"T��g�W�5�m�f��|�2O-��j_�����R��8�U���`�7��B��s뙧��jR�t������UG����z�g�H��%��� }ޟ�J/q"uhw8�s�B�fC�-Sظr�vyM3��j����:�<�lܼ��e9���|��8>��xL����(�YQ �ŷ}��Js2�i���3��;�`"��F�%��`������f�hiutޟg%�fr�;UWY����7���&�u#���㘥{]�E��H>؆S��X��ٙ}�cΚ@nV��]���J�d�RPV"�xl�4�F��"��K��8�S�Q�\���sʱ��`���)f,��frGRb�i�Wa3�]E�=�*P�P�QT����mlE�a���=���.`�T<���s�%d\��~�DM�C��CָԢ��.��s;�ho��r&�L��A5��$��n����(Jȿ	r�nz��7P��+���^J�)�mr�i«��X���lEg�+��0ϧa�r7��%
ͨH�ml�sR�̎j���Wa���h����1@|^�8����W�8f�4{��E�XŖ��Ԗ@�wϷ{q�b#J]9�F��S�F��xd�QK���,���Yݎ�����cN!w^3�6�q�C�<ή7���SN�'K$ײ8�ʬfN�F-ۮw�sc�z��Ֆ�j��./]��p�7౬]ZVu��jDM�uH��q��]s�Ɛ���6��p��Z��S�:.=��",)�4�1���K�����G`�p*�޼����u-&�������{Y�;�Op�A�c* -[u����rINb�uJ6����1+����ά��=��������o��x��A��:�;19W+;n�;*�ٜ�G'.D6����1�����@ņ�4�u�;��$��Ч
�'C�*R)�9楞�'��P�����"�u6���}j2+X�N{	��*�"��,����4�uѰ��Qa�Q�9�(��f�Dt֤^���t��^��.j�X�u!<+��Z]�y{%B緭�k�*�G�dg��w���QFC@��IVJ\�Ơ`�ֹ*ā�<��C'����x��_�N�f��<����vZ��M'�a�f�OZ�3y=h�H�ZJ�J��;T_5��t �j�`��qtyַ_%kf�7,?E\̡n/
gΝI-��^��+�\q�ncՉqv��߉��7�'=钶D^Ѿ��? OQ�!�Tl�O2hxM��/
S��;c�ov��*��Η�q˞-9�'���T�ܹ���v#bsG�e�f��9��&�{���) ������#oR9�p{��ʉ+꼔��p2�W:�����GL{��Iܫ;9g�ah�.|z��;~�q��1z�F/C�	�{��+�jY뙾h�rfY��] �jO1����m��<ƽ�<�}��|9��)3�$������wׯٻt).8Z�]�R�n_v�%�nTa�9e=��G��>�=6\�΄.��T��fz����Ԇd��Ǘ�����ȴpi&]d�ST��#׊M���9G8	ym�~��7�Qb�
}�׬TS:����x�9�=��r�ҩ�f��|we��W�ܡ�w�����g����6�
�ŌM�C|P�75{�a�%�ʺ�ŕ=������=Y�M��k��5/�W���>�����62Ԃ�dd����*ݸ��0Yz����i#3H構���E���3�.�mS��r����O^�L�G��Y}�я�{�5v�"W
b�1kb�~|a�S�f�����y�f�vθu�̾耘^��jt��Έ�<L�%�]5$uL�1@�p�/�	E ���	�(O��w[ts.�U<���̚�<O9�/2�޵��0_�Cج
��,>l�C\�)瓄"�^�
�jӮcf���܍e��,�����#�c��h7.!)\r�W��5,
�"�][k�Z9���![-�۞آa�WCH77���Z���т{Ƶ${���Z�N*�3݄��mR��m�	A��k4�v(�x��r*��KҮ�fË$�cZU�]����_h5v0�4[c�6�sz�p�n^�f��=+���*�{ڂqյ*A�'5tF��È���Ζ��wU�2[�������[x�k3��qˀ݌\�}���&�8���t{��4�3�����!�Juɣ�ˮ�Үx����槰��At#������fQ�}1�^�:t�L���E�����:-C:�d�y�G�;�¤�'Ԧ��[}�e����/���G�j,ׯ�עU]��97�%.Z,}#G������s�[��R�f,�Im��too���nK��K5�c~�k�� g�����ts��2�M~����x�Mh
C��'l�|�C��!�g����|���~�8�Ұ�>���I��S�6�a}�A�&�H�+������>αV��lQ�P9�\a��a#&�)���T�[��qN,+�^L#�����p���hؙ�3E�6vw�6&�Č�M��͕G���^c��vVW>E!�U���z-�V���V|v(���8Fy��݌�q��+��ΰ�l7�n��� �� m��2��
�Z��}8edWh�9y�Gq]#��Ypƺ�P��=���i>0{�.��eiz�\V��{P ���=���������cۚ�O��#l��w��;~wAST��w�h��~`GV�	슦���å�!3w~rǙҮ�Z����y�C�k�年5�7�5G
p3���u��~�b[��\ƚ{-cY��G���Ye�BK��Էo��#�ݢճ��j!��7/9�нr9pb��^��;�
-VZ�9����!ɼ�[��ig�^.�b�/��$��Wx��,=2��FF�ud3AL����Ѷ)�#�`�^P��=l��uOH���j@�#Xs����G�'���z��.�"G�v�X�Cx��Ec��;�c;�S�6�L�*VyP���g��{�F�j�k<�<�<hVh��0I�z���iO^%�X�����(�CX�s�\}��p�'1����ym���l�b��c]�w�^��a��oJ���a7�^���T~
�U�:��/zp*t53T0q���8��gG�*��q{�aR����G��6瀸�.��p���ּuS�"��c��v  �]<.g�R�Om%F��c��{��6��u�'�J2����k��Ue�z�.j�d:�\[����)���M(&�l�$׹�9^o*�²� <	Y.Q��*�Ð�{/�+�yMVm�O���%�s��y�GLNm0`���6��bV'4E	���;X������W�D9Kmh�O��|{5�i{T�sZP��8���c���&伷@R͹C��Y
�)o<�Xrby�V�ϟ/}��,�Hxo���}l�T�g;�� �p7;b�P�]����{��Y����۷��j�����&���`�����]�D�7ϒ� [J>��ӯvU��ɼ�jl��lL�w�v�r]����*�a�C�;x��繜�iC��MC���|p�;$Z����,���{�7(OJyKbBh���d�k�sN��UħS�ĵ�{#��S�߫$�姖�1aHvy-H����7}����>�A!�9^�>�K����
�t11h=jPO�pN(n!��i��Ja��|�9*'Hb;�D��3ϕ>SD3��^b"�n�eP�GZ*��ܡ�=ze�9�^n����6e/rS�:��c����0ڗ֎�^��jY�k"4�H��Dc���+7n��R���#�8�嗸6�e���7#�X���#Ǉ��
i�:61��;=�GR�A�Ă4�iR�ׂ]�y{%B��޶l9�H����)6�s�U��o3��rϵ���Fʇ� x�=49��OQ<v�msPz�>��̭a8D�~{3g���8�5���/�#�(��
�.�=N�/�^Tq��C�=<��Oo>f�z2����E2��m$%�/��R������=��"J4�7��kgN�����憯]��N���_�^�g�l;p��Iy�T�Ys�j9iW\�ڽ�P6rB�4�&D�t��S��2J�w�rJV�.�Q{X �wWoK��f>�D�&�5ßk6�Jxv
�w=Տ>ȆA�Km.QPĎt�}�\�X���N/�OQ��!�Q�!<ɪ��x9�)C�Vd��,�����n���tϥ��c�H��^5[�������$5؍��r��	�Z0�x-35���z}#�[os�X%�y��҉g�~A�Ȱ1Ȉ��$F{��˸Gb�j��M���X"y�S����
�_�Y`�=�8B9W���چ��"sX�]_K�#�D�O������S{V��jҟrÅ���7ۍbw��=��+ڳθ�yN)ﺴ���������-�G*�~��Ө�"����{�E�k�Vn-E��8+����9WɉB�os*aW�=�q2�s�ץ���Hy=T�M8ӻ�O�q]�}�v�!t�v��R�^����潠��V�x�(��Nជ"�6��v��{��`�i��ӭ�N��نa*����}���
T0�Z(P9�$ŭ�������ʇ=���'ٶ���1oG`S7Q]���b���#x=�3�����J[HW4��Wx�7Xd.g�ر<z��wm��ߎ��W�n�+�H�a76�S���f4p-��6n����;Z�rg;1��g8ĸX���!���8�u���ޮ@&l�JvM��p��5��G��_.�,����ى�Ć�˾�w:TL�E��wn�]������"uan0vwWksgh��n��w���"���0X*Ē�1�g�꡶����J�g[4ء�����gK3�����#�k�2Q#_��E�uJ�.3mF|O
c���@ r1,�K��ߥ�-��-�(e���j�+�,��Ac�Dㆌ,�ѫ�p�'bW���v����J��Y����No�'�"�'�\|n�Ɇ�VI�5�y���X!�tG����'�a�*�}Y�@��X�JÆ����b���:-C(�,Þ��KD�-���H\���8��t��!n^�K�^<�Ƶ%4�Vʅ���p홈WpZY2J��ˎ��Z�h�n�a��Ip�Hdq�W�֘��¼��8pk���r"��Uū�+W�rs,x�K%cz�&$��7��%�,�w"�O�,HF�Ք�7�ɧ<.:9/D}�Z�$�m������U/��b��遍���U�BJ�AUώ�B �}V�Sj�z���z���=Q�$��p��	�Y���#259���M�L]W�x�;�y��R&Y*/�#G�ՅK�[]��5r�2��,�N;Ӕ��F%��Y>Έ��ʞ�JӨ&v*�y�e�9};�s�sh�F9�p�s!r�8x���4��=�i�Y)��ye@C}�^Z�C�+XeI}Q
�Z���:�ZV��{WFI����N�ּ�`�O�.�d>���u�Z��;I��p��Ϟ�&V|W'�./�۞)��f��x83Y�^�K���R���R�����R��K������8E�ژ'WN+h.��{��������e��V����\S5�ڄ�g���a���Qp�Ď����r�Os��Y�!(��a�R8���L-;򉎴W/ &��$:Ȫa�ܚ�6"�H��&9'<��,5��`>R/����5�Ɋ�����3��xMi�#�RofLMvr�K��D6�H��J)f�=�I���8'�M�ڃ���W�25�ї3ʔg]��'+������'���,OKȱQ��g���t�[5��#w"��9���2�U��R3�<K�$�8��E�!P���p���SL��7/��u�-�:fX�QB�����\��|���,� '�3��%b.�A��e�:��=��*t5g�]�2z�����[g�[е���O|�O��1(�C�[I0v$u'�J�H�7(�����ȵy�C;=�әb����!l�T>KE�Nnp�2͜�^ơYCX��:�ݹ�[��G{�!c2��ǚ�2v1��Y���@��(��#>����Kjt�7yc�3zDʾ:�]`yO��{8�:x��XJ�M�d*3m��jw'J�=]����Ѽ���h��8��4������6�3N���=N�m��$&Q-��gi�^�+	��^1��;&e�e$�c�!ޅw�����{񝪩V�HQ���T�8&"��fT��X��Z�/�1��d8q}��j�g@:�5�-�v8� ��gc�:�7"��m��Q�x;v��c76�L�ۖ��`���9���64�1�N��pUՄH��T;7w�͟GnX\��0IT�)�8n-����ڶO�9��85����9����J;�.��u��KI��Iծ�WN�m�z�=�ĭݻ�T)[����lz~'ؕs������3'c�]x/0���\�h/%M58V��:�����j3;l�LZ��Dζ�r�L��cm2�|��ʰM�M�j��(Z���s+�G��O�rO�Ӽ���5oH����[��0!Z��ˉ]ǲ�����V�e�01�.p'6� �@�No!f�j����r�#�Ƥ±��Z��@HG�ȡ6�YB��G�^���0q��p�O]��	�v#��uEq�x������"�)�k� ��sY���dz��:H���sQ��J)��7��%�)'�]�ƙ����Z#�}�-��2�շ8��gdզ�U��^�6��W��G�d����řمt/B����;%H�T�7k]:���]�mA+a��3�!�͚��W	�o��=������v��Q���5R���P�rs*�;��MK���`d��J��S�J�z�.C+�g��'�)J:Lf�2�S���C��͂#������	=u��ؔ�\�^j)���;���;hVR���"+Y��0�`.g8�DzRw`�)���@���2p��4��*kf5�(�˕�2��47��=g�{�<\^�ˑ4'���:\�4��چ�U7����tw9[��q�2�N�zAݮ8��Jb�M�8w��% �ڱʨܼ7��� _c�90��yZ���E�|5Vwe
EZRh��u��vj��?hQt_u`��c�KM�F�И���d�3�s���%�s��Gb\䎶%�^T�%;ň�+T������>�'e�n���C%CHAշ���o2�R9`�ytA�M�Igd�|��D�.���)7�n]s��E�"��|s�j�z_a�:�Dpj轔g@]+��1V4ڠ�o��$ד�V'n��p����7u��CE�O��q��֏���@�5ng^;����������( #4�m-��OtX����	.e����S��Q)���,�l����u�h�����]H���M*�y+����z�~������TEETG-b��-��
(
��Tp��ZWPqJ(������	UXT,QPT�Z�k*�m���F��T�*Q�µPKj�Zتb��,T(��`*Ŷ֪��J���Qb�DbTj��(,(�(�2�q�PQb[
 ڲUR�Kj�Db�7mf(�b�.0X�kqT��3a���-�b��aD�F��QŋV��cm[KT�+�f(TU�QVEE0�Q�lPUF*���DX"#F�DQ����#-��\XQ�(�Ռ�UEEB�"�Kh�TT��J-�ـŔm1�P�Q@m+RQZ��*�F�m��)�����1B��մ��m[�U��,P���X�Fb��iDbThU��p�m\8��b�TTY�%�UE�-ŘX��b�[ETh�a�0E��*(�UT( MZ���tÇ.��[x��%;�j�9���yIzyJ�����$���/F��UU-�Z^��Y�����5�G�fD�rAӠ���M�7��"0�J������=撄�]kJӎ��(Z~\G��ߢ��>A���6U��n�CIq�)~�`Z\D�̢M{�����{ⲣ 0�+�\��}�R�0�33��)�<Xw!�����.8U{��FN��į��S/,3mi�K����N]�s�s�ӛ$���&���^݆o#*�2F8�l0p׻U8�v���K:tʲ;&vD+]K>��^��A��A�C5x��X�x^�`�F��d�QAs��,��#*6h���7��uj�Ǩ�l��vk�*�c`�6���p�>ţ����X�X�|/STo�c�}��0<uǰy^^�h�l�͕\b�P3���0�#F��X�M�y8�x�텝���ʟ)ۀ�m�^b"��N�����O�ƾ��3����=��V�ҵ&=*�����0��S��l��u15��R� V�*C��w�w���v�<���$U��7P���R��L�A��m����(Y�
��;�lg_�A���z�+�&#��z�d�=�	uo'��p�[�w�s\3M�jɆ�'.q��l���\�܌�ke.,��r7F�n��M�Λ�ƭ̈��5��U�o�u5lĻ���A;;@]}�fC3�q�[1m��b��.�݉]ʕ��л�^�~0�(�i��COHj���%�#\2�r�7O���Ι�#��oC����3͉c;kن�ϲ[@��F�*ر"��^Mz!͜R�hv@��Ȓ�]����=�e�r�H���.Lu���X��J��\q��'�Ȍ.:���zs����<C
U-���vse�QB�C�I�I{�H�o���TwFo,6�ҙ���¸�XPČs����p$f��!��K�!��d�|̬�T�B�'�o��s8���ޞ,z��~�DW���T��Ȩ�&`2�G ���%YfIz��þ7��z�bH\�L%��{2����ˆǖe��A%������	���D+�~m(=���iO��Ar_n]ѱфaVI��Y�ɒ���/��0o�D��(C.Y@։�vμX��Owe�@z��A U�۽�P��bv%�MJ���4�S�uiqs�@]�	��|ա2e�uDft�0�w��	+�X=�6�{I����6q?��9��37���j�uLA��ck������ �k/��ް�����++��	��@�۶����n�n�W7p9#�n՝]�L���N��h�Z��<Y�����L�X�*އ'3(���3��Z��6:u)�vp�Wد�%�9��@�C�S�x�ԋ�)ݜƨ=��K�q�w����_D��9T-8v����f��G7�j�AA"wiyҋ��EץS�gK����o���}r{I�fZ�h��;�ia���է��
�kQCHP!�9D��.Z<���g��Kc5��i���̩S�S��t]���lk��S�pؕ�R������H�\c��\o���X��ѱ�p�e
��,�2���9�9�O^Kw^��$����џ{�%�s��_�Cm��䕓`1.���zzfu.]�a�催=}�L�w�w�(����dQ-���mR���g�x��$$��z�}��Y�r�b�e�s������t�/�łt"}\�tE�atmn�!Zkצ�[�ɲ�Y�*%՘�/�`�|}����M���\|n�u�0��!up[��)�=���f�M)��u�u�/ ^��{�E�^;*���9<-Cf��z�I�kw[����R�0z�Xd>0Wa����jك�e�Լ^<���Z�s��u�ߨ*�S.����>]���x�����O1�32�N�ʒ�ֵX�i*�v�Fk�9� /c�خ�y{�c�T��2ԯY��ͼ9Y�PMي\�dg�r�@��<�դ	t�(isb�-�aܩr�����ud=w�+r�rŉ���n��n9m9�n�;f^n�M1'4p�e���y����H�@��u<]]�c'u�`�J��I��jq�v�����w"��1����r��W)�
5�sW��P�@z�Q�v�Z�/���&[��|�ǵ��aɯ43k�����ٟE1���y��Ui����²��.�e{9�O-n�}���vmy�3f����O��ߩcKg�EEV7Oud!VнG\�\ٯ<O�-݈p�D�*�c�
g^l)t׊��5�f� 'Zx��[�in��*EӮU�|��y��V7���̸��8�~^�4�ςg�����g9��-�L�ROM����~�u��oʱR�P�!NЈ�@K>������m����;���7�j�a�v���O���x>9���B(P+��D���xgkc�M�{R����E�Yx����)�&yj��c�$I	������=�'��a�sF������Fu�'[αˍ�,���T� �ot��|��6����w�{��r�T������1�F�\38���NG�9x�YFEҭ'5�s�w���]�g���P�hm�mL�1PݩԶ�W:�"n��S����N}[.����������<�%�A	٬��^��y�՝�- �ҍ}�s�+�^Q}{c�e%Ϯ_;�l�nW�\�W"�o+��9�xN��$
�x�.ɡ+f�R+�N'�c��R��'j�u��}[3yK[ɻ�9��	ވt���<K��n��[:�x�966�P�j�6�u��+͕�9�
[�>=d������?�g�v:���
�){���.9|��mb& �n(wS���z��,���F�gS�+&e���N�-��ޱ=u:��)�ã5|��7kM��=���v-D±Kf����7;��3L-�/�.]�e5c2P��9�e�׾K��]9�g�[�oT6��<���m�JB�;�sJEd�W�
�K���~���F�E�9fn�J��[�����y���'��ʁ�21���(^&Fq5�*�2���6q��R|���K���H�j��j����̫n���F�YE���񬡮ބ�*�6��sK+���+#y�@t����̓���՚Bc]���N���ӭ�B�7��V�[�vT���.N*�ޑb�嫲�u���{9tr��i��M��>�v�mU�7}�c
�(TWQ�����[��n�$jPmk5��G-V:�{�{)��
�P
)B܍�48V��A���;ٵF���jRNP٭fE�F��)>v>OK���j�X]<�"�*8���Z�4p"�	��S�!q�Me�W�;�+|y"4����v�m�����l�93���:��oW�kXSlvǟ/w2��h�z��9H�n�rRu���ϕ޽*��)#]�s�\Uk�+��]->g�iMY�N���=JN�:x�kd���dP{��|�vS��=�mX�Xzzf��c�����nwB����<e�ɧ��jo�����j��{�� ���~�c���f�Y�{jG�üHΊ	=�C�vU�W�[d�"�ezo���̵��9��y�U��}�4w8��lӖ]X:�+��7�)n�d[��7YT<����f�\�ٙ._q;���z��d��>�߆�Ӓ�Pz��7�c��.��/��Ily�W\�řx�Pꋛ��gH��v�N��(!�I��J��HɃ�p�#�'9����	ڽT�Ej�o�]�3$��Fp�9�>�f�5~�w�У�����9~��~�k���RH���G��3;TZG%���Xq�</h���W"�ڼ�B��u��YUjUG[�(6�49Z�c����An�� ����b�xD���[�fnZ�Ɏ}�۝n��4���[��q>ΉX-	���)�,�tJ�JVS|�ƶp^.3��*����������i��o[ އ6S�*��m���s_�q�;�U��e-�׋��N���33���m�{Z���v{a��_\W�+Y����#^����5��8��EHT�U�M�e�=Օ�|ߟj����Gb�GK˝�U_ze�I�?L���@x^'U;Gu��._�MX|{9���P����	o:�֦�h+�ɷu�Z�r�=$kR^��ϝ�MJ{ҟ*@k��1�e
/��V��n�l(5m,\/�ˋE#Qsq���{;3-5��(#�+(����&m��n�
$GW^�����3F	��֚[���ʶRб֣5�ש96�8�`��!��Z�vw�SǜD����+�,w �䶬J]8X�-oH�r���k���.	�
�t�K�B�WQ��b����F�\<�:�o�:�����U7ac�3���4�*�s��;x�%q��n�������Y֡�nrtSTT��%d݋��/�f��䐸%�7�4!�L-�W
�1f;/:���ߓ3��gb��|�6)���Ћ�R4t���{,C횕�.�P�vmdD����Ѧ4b�]sz�icz=��z��=q֤r[�w⬗G�]B����Uy���[�P	��(ܾ�Hk̍\�K���{�Pl�-�7u4�c��[WҮ]�m$l�x�Z�����6똼���|�����G$=���Xrh43D�TN��\us%�����n��r�l�z�-�\�W��4�[��uy��Y��;�8B�ܵTO���)z���=�՝ZSB�r���.l�Os�$nfQ�$��|�o5��L�m����~4�*���޽�S�N���[]ti4��K!r�;��r�F���t��D�n��Z��Q}�����᠀c������EqqII]�(țw[��RH��ӊe6�흖\�1��Y=���c:��d����oV��K:vN"�m\�M���X钝��is���r?f�0�����;����2�>�X׽�ѯ6~�)�q��;P��'S5�|��o�M�F����mQ�b=����0��7�~U����vx.�idT"f8v�tY���{���"�c��%*ް�$������)�E
+���t�I����:{��RsӴ#Q�k�b]�{�R����.��W����U3S�������q�Tt�e��)��B] Wm���^�Е����W5]�ԑq�E¸H�=j.<TD��<j��6S��O0f�^�y��h�����HU�J�y��˭�.��ݑ W3Ƅ.ɯJٶUq���S��e�C��ʍZ��Try��ݴ�p�o��'��-�=o��*��Г�{bC���v`�z���cwmkQ,Seh��Їt쫻�ܨv�5����[�W��V۞�;y�~�~���{�􇰱�z���;*ͽ����aɠ����R�:v�������t>z����9��{�# ��� �l�h�b���ы3ʵ-<&�KЍ�wv\G-�*�=�ڭj�\�n;��\��ݲ^Չ"�c�_.Fd����skg;t⽴%e�+.�N+�= ѕm�긴T�_%��l��yr�ERt=y���@��w=񓏗<�ܽTڕ�j��V���b*]�VX�����]d�wv[�f��ڙ��)�ݮ�ww[B�h��v�gJ�؝���J�Y(W���[JH=w۶��3�R�j�m���J�A���:&���N�WJ��_���u�'��F��
���"��M퇩�㷻j�+��F߰l�\k
�~�'6͹����9�h`k��<Ϋ������)��V*�P��؃"��˹u�n��{���F�t��|���z�P�[��oϖ�ĺ#���9S=���9���eDk�K��B�i�щHW�)>OX̘Z�W��I{�&��h�������#¼_ez)���}u�݌j�霄����|»�wJ��g�JS�+���VL=X���D��t j�Zz}Z������I��$�	'��$�	'�@�$���$�@�$��	!I��$�	'���$�$$�	'��$ I?�	!I��$��$ I,	!I�$ I?rB��BH@�~�$�	'�BH@�~�IO���$�	!I��PVI��yJ�@�	�` �������ׯ��� k!!T���&�*�`J�f��@�&c@Z�	T�V�Z
U�
(�h�UP ��
���6Ւ�Z�Vj5*kf3Z�2�նٽ���������Mi4�9	l�'���eD���)���U�������ơ(���i]�r{��і�-�m�j�*m���UE�*��JkZcm���bb٫lhm�%��-M�4*B�f�Ѫ��%�J��YQ�l�,��F�,i����  ;�ނ�U[ln۫-hm�֓�e)A����l
)+L ֪�s���[B�R��R��kl����N��`j��m���T$2Z��e
&ݷ2[�  p�+ARZ�5Z�kM��MVZ���(j��km����J��ƖZ���w[] ��V�mwmJeZ�����
(P�EQ=[2�d�E����k\   s{�
(
(X=�P�E
(hhL��Р:(t4,��
(P�B���(P�B�
A���
C�Р m��xR:�i����m4Zj�֕JXw�u�K"��bsj*V�ʼ   ^�4[U-����ldm$����Vuݶ�ʍQ�%2����(Յ���JV�P�����	ܮ�l-��\��S[7E��J�P*�V�ڂo   wW�m�٥R�ڀZ�D�P�Ղ�l�m��Tm���uCl��cZ2��0(R�֫@lх�XRu�e[Z�k6�R��S��0EI[*�f��   ۼ�N�w+r�n�;�w\ӋUZP܍]+M(J��-�R�Y�p46�5�]�C@�4�3B�K+�ݴ�P��nڭ	3
�e���mQ�)EJV[V׀  �=��5V�k�f��K��U��u 
6��θ�*�W.Pj��
SvEQ�Ө
cpѩL�5�3m��kFmP�  ڼU(���A�T���P;WED����J��PkS]9�Qv��QV�ۥu ���@w4�Jٴ�m��"�S5�e�  7�R���w:ݵC0�@	]%��A]�����ҪTn�Tj���b�ٝ�ӊ�U�UR�lT��ջ�fl�k�  c�5�	�� zW]V�3up붠\:jյ*��s�]�u@Ωܥ-[M5gWuv�[lr�EtRU��ۃV�R�Lh2��   ��
RU	� ��a�`L4d�)� ��j4 4�T�I�R��4 `I���*�5)��O�o����~���w�2���|���%�&]֔a���]@��1��������vG�x$�	&�! ����	!I��B����$�$ ����������_�X�GY��˃X�mĶ]JsY�԰2��m5��摱7p��V������	U�s5E ��q�7p��D<�s4��&l(^��j��O{��^�ZSN�x��J�J�8�څji�.��SFj��r� 4�'^�{�ŲnC��[6�x*�'j��fPwb��F�Qж��9�[���(_i����w*l��5�L>	������U���fj�SdT[J�6 ä���f�y�˼��Ӑ�c
�L�?D�	��.H�3r�:�w���I�5%��GBM�5�Id�G��9r&�s�#�[��e���1Yy����m��w�M�Pv�V����e�=��[T�j�Z�i�f3�o%k�J��W:Eލ	��ۃo_[e��Q�p��fع���V/XWf�e��2�2(GB���Yi^�ܹhYia Xͭ{�v��S�e0k1P�KD�����0"��T��GJ�:���[u9w�i�w/]Yk6>M���0��.��dRM[�����
N�!�@#e����$-ެ�1��͛��eaE��������gA3Y�N�s3e�f ҡ�wіZxZ6��m���;�hE�7;_`��t'�x�'Y��n��09�h�bh���_{ע��6H�tm��E��.�L����EU�`�˾�Yt�3c#}�d¦d�>{-�{O�Պ��M�i�w��0F,J,1�Z�S��4�(d�Pn�M�j��������n
W�ΐ9\�+W\�b�cd��	�ȉDn���#E��x#O��:֊�/h��{����O��!R��D4웬�G���Q�*��f^ͺ8ʶ誽�6}�Ue�cջ�Y�.�n[CM�
�[���&D��MYy2�`��f��K߰fd�t�r��d*�I��av�E-^���Vzh��WW�֘���z+Yc(�ኵ�V
4!z]�w��-�n�,P�yZVm��4�\t�^�ܘu��^�(�T;)����Q
�a|!Q9�ݷ�*�Y5K�WY�V�I#|]CY�O�A��D2\ܐQTp5��e��Z�QYwv�4�����r�7,�v�F�`�T�����qp/uD0�;��Ĺ�y��"ed��n Ζ,�ݚ���[Q���D9Y�6ʭѩXV@��J��~����^ŶC�ܺJ�]���� �Nq���y��F�d^;��YN��TXh`��4�R���Y��1Cڧ���y_b8�B�XZh�/Z�Fx���f��6/Cu���֮�ٷ��Y[�-�6�S�)P@M�E�ǧ*�mnl����*"Y���d�XR�����Z�J]�n]]kv��	���h�
��+��� ����W�yJ���R�0��n\�Xh�>\�^�����-��$�j�WoÁӬ�z�u^��g{b`VU�%|��g^�z��	�QÏ����.]l�b�2�"kc{��.��)��`Z�I�RzV"M���٠Q��t��m^XU�(�ow`Q^��t�Y�w�2�t��Wwf��ʅ�+�c.�k8��78B�ڕe���hrhQf��&�lڬ�H��˰4h��-�$m�9pe��Ŏ�m�,���E	�-�M��xo�GVZyE^�L=��m�GV0�"p;�{k6ʔK���R����۶1�v�")౨��������.D+e,�4Hd��1KQ�{�4��lle�)��W��ڭ��X9�B���Ռ��!�#�ȶ�����4���{?<�w�O�# c�<lҌSC]�KO,���/>�Ct3Cp��@����j��V=*�9
y��OY�+"Վ]���Qd�V,�Nk[��zs�1�K�;���$i�7�ۚR���ե��b���p� ��@1fq�[��2��o\*��A������˥BXeZ@�ֵ�5a��.&_��U*ƴe��0�#%�H�SI��^B���ϼt���G��#<��k�Z+;u����1��ahR�C��pfp��A550;D)�y���:SoLf;��(�I��23�WKo^k	#���qlF�������U�gR�b\�i7&�����Մ�%!a�I�w��sw~ɯ.��wC��GZ�2.��6�b����i$拑����3�F�_</��[ 7�pp�ݺ62��@�a�9v��i'��5x�PT�qjж�n�U�1��q���ueۦ�3����L�[Ϭp�Pyo�4�q�B�m��h[ Z�m�e����pX����4��j�*�4��MO�W��pk�.��qZ֞�����ޗ�nͺVN0v�����hs�骮CX����e`\
8�<�V�!���Y�}cJ��M[�k�3v �Kg�+5)1�����R�R�śNP��,F��vu�z@.������Ֆ�۶u�=��}<�M1w��N�O��6Nh|R�Y��ZI������ʚ9���R�b9t]L�ߙ�[B��6��9j��5ya"@�)�f],OnC4쓤�c;ȶb�;4t�lO{���7�n��b�s4n�E�i@m2y��g�+�m��ɮ��6uSõ�Ϲ��=��4rda���T�1�a��<ۖ��6�I{�+0HkFP���z��!�@��t
u��6Iu�<)˼�`Wz�:,����k S����f�'gTU7YB�4���Dm�i�4t��W-g��_�t�a"�S��N4/rƫ��1m^ԃ�Mne����c�t����3�IM3{w��6����A��T0�Kܽ�.۹�a��������Hn��Q�����ɔ3('3�S�5*��d�`1�k�����&U��G��T�z+-�5���8��/���N�1&L�5�k>��ۀ������5�6p��c|�`�݉�R)d^ƃ̕{{�)��mʁ�b;1�ܽB�a��*4�&TtI��i��-�M�0����5W*�ػ��f]�wk<��Vd.��O^��.�6�N�'���9>9+S�[�hsDa���<i�Oxg�n2����m?87����%�wF��u��Z�˽!Z:�aL5��s��W�"m!]�S���u�:�X�H�J�0���7���נ�}n�a&��l�X�<M��\iB��vR�,�oᆋ$S8��ܫ����N��g47>��a5[X�H:^�ܑ콰@-�ٕjfS,+��s���Aof-�z�͖CJ*!Y���<5ڗ�,<���~��a�m֝�� �ͽ���*���n�F�1h�&Ȭ<2h��������QXH�or��� �[��v�|u��v�mi���Z��w���G�Oa��!9�M�v9/�5�n��<XN��e���`�kߒ���"��̠�ݬ�Y�a>�K�!%7~��f����:���A�)PJ�B�n��C �fu--5E��*ỡl[s10�7�����1��@�l�"�k b��µ�մ�^���h���$,�Y��f�V�^m���x�-��e�����7̻w#V�#nc;�Ywku�&�3.G7cu	�l�#�*TW�	̌�
�v��c{yysWk3i��5��8A��<N��d�<I�0Ѻ�,�/o:�7�p����9I=2b�79}F�
y��X��^-�I
,]2��vsI�He���d�M��4��t��Cf�	��(=�(�N�ͩ��j외���GJh����rPK
�T��:v�d�]�S51�^��&)�r�ژo� X�)�@C�ں.�M�`n�&�d�3`�ޣl�c{kVlvo2� V�"��P�r����&Zۚa.�<�iV-E;��5��4�ne:.��n�ݜ����Ysl�A'n�4��쥹��m�-3m��S�a���ՠ�Yvw3G]tؽӰ]�"����hڻ�zN�bfQJ̗�ee�7�F�<6�tX9���Ӽƛ�*�t���(���d�+yX7)3Z0]�g�c�"!f��4�zTU6�h�aZŧP�'��wC�k7f�%A5-�k���%m��G��ka����Fj�/FѨ4���M:Ŷ'�az��]Z�}��:0^�M��m_!���wYy���k�[b�=_h`��W-�rR���%���������爊igg-�N��g�d�y�(R�w���t%���7oP�T����ج�3/�.Ώ�^:�b�!�Q�A�|�5��~�[v;�*�9s�A��fV��g�M��[BX��&�n�aX�ʘ%���s.�[�p��"0�=ٷkd�R��v�f�:TYm�*kZ�ћqֈ⺛���P:D���n�*4t��J��i�Ȉ�Ċ���6�^���oHWN�7W%n�4m5׺�<�s���ũ�3^���-m10S6ML9�����aX�=�\3G�E �����ޝ������OBKZ ����!]We���g���2+��*K�Q�"ֱ�R[ �ǧ}���nt��\臊�`pUû4��t�1J����2I9E�o��#ܯ�Z�ݽw�ع�'P�*�0=t��5�u���P���Vi^}��̺��e�f&�칀�n&���T��nod�I$T��D��Ax)���]���-6Ĭ�b�X^3vC��7V�3#-e�y����v�k
�|�umV�.��[j�4��wU�LM�rKV[�Ǭ�(�!#���W��y�F�9N���+[��ݏ����(�]��R��I��5c.�[�3q��*�솅�b�D
i�-u�Q��Ǧ��z�D6���;p�	!C2�f�pI]��YCwr�'�,���9z��Bol��W@7B���]i�u��zb�F'��{&�hA�(3ZN��/�Z������S��t+u�W{j���?Z�e�O�r��j�4���I���5�۲���`��[��^�x�Q�S*�V<�kvFoY,/Y�*:%|
,�:�[���9�6۳�[Wf��5Q�j�vC��?9�����#�Dx�A�|	�'Gyu��槗��.�Ҟml�����ƍu��k�z�t�����{k�(��x k�t��Z�\�fe����	r载�_M��nYכH,��af &�Sـ�Ɏ�E���U�b�ӡ���[��އ��a�C�6�a/sv�堋1��fn�ۦ~@�ֱf��7�F:��K'Q�˴H����H�b�9�(�a�8����I�)����M��J9�����]�m�m�M#�ic8�ִ��lűf�$��vH�˗v�m�����w��Ր!.�i-۽��*"o�X�x����ĝvq��`��e�x���K��k@gw�A�RQPe�s!��4�6�@���Op.�W �Y����Ç9B��7��R�[�c��$8��[S0�FS;��
Z��t�E����cr�;b�����<��E�h̶�C�E�[w)�-���5-4�< %�VUи�S^H2V-y[qJ�F6��Ĭ�b��YV����-�N�U/X\Ӷo��s��5ec��-�6h�V$��o����m`�wx�ǁ}YaXV/%���*%Z�陔2�Ѩާ8n���F���;��w*�Q̦� ��,��`��y���ID�Z��V����N<<yp���óxv�ø6�%��Ua�N9��:�w(`��cG˦�$���(�K@T+� ����wA�n*�P#��R�[��b�·��6wti�;z���hȜ�lZUm����XO�v��]m�:�1������~�"kA��vG�t )�0qC��Q���{o2�z-�Q ��:�Mn��\�I:͛2��N�͡2�Ф��壎�Yh���;�TWlE��׊�	� gM�9{��l����[��t�öX�P�bVY�sX�r[P�F�ۢ�a���Y`:e|^*�����1X�<t�OE����\�Y�g~���9�a=*�Uk�e���������;,r�iM�����ͫeeû˰�ا] )*���[`�OCie
����g������%2/cԝ
`u
�"�[�")7d�Y��S�{v��9�0Y�pd`��v��-WH2�[�����O
y��q=��v>|��oX�� ��K�6V,��PhF�cǆ��ͨ��?<�E'{W#�+ ֔9�`d�C	�SXʒ���G�O��4�P�Ӷ0���{��h��`�1����ӹ��LG���]l@ �1���ee�9R�j�t��U��Z�-�H���z�Z����Q��A�(-Xt�8f�Ɯ7He�i��q������C�Ĩ*�.�:�������X4+��G�K�N��fb�zb�F����*��ss7i]MX�+6��4KYR���A��X^	��BZ�V*}k�-Tq �1�x���P�۫��̼۫�n��k
��С��t�V�$����I�[�E�LЕj��{�d7�]n��Rӣ�"Pૉ��f���+�F���*��5�KjVe�2�J���dŤم���������'����9�/݀�L��"��Q.&#y�=����Z�����Z����	
��H����R^e�6�@Fڹ���0U=��ڒ�"kWQ]��d`��Q��]`{xk�l�F'-�a���8a��[�*�b�x��\���"��]�MA�WwG�aR�E��L����_R�֎��ҽ������(�$q�1m(� (�L�3��,�B���nlh�[r��4.��m`��WѼ��*��[4ګ����E]�q��	��Zw7c��At35��VE��f�/Zz̇,��M�䍌�s]ͫq�c2S�r��H�Y���j�Y�e�KFh�2eB�̥^��F�A�9$���f�Tuee:q������9�EA�w�Z�@p�z�F��gk�RWS��+��)u	��ʂ�qed��	<�I:����	 ���B{��$�}(�>sB�0�P�Պ�B�L�������8F�]J��yA�+��{�;��Dru
٫a���:��{�?D�Rd땯S2=�3�z�����dIW�A]��Bt����]�WZ
Ӗ8�`e�Fo
Vnsr�n��e�[�0IZ�Ys�(D�iE�j]�[N�ݺ�.ƺk�Գ[玷�+�
(��y.y>8(ېm��}�%h�M�OX���f
S�y�Z�1+�t���ڃ&°����#��7/ ��v���|"�ޗZ���O;��F���L�*a��MLԁ���CO�d�_s��Z��x7x�}�������������3OE�,y(V]�9�vN�g6��be��N]�M��k�{�e1��nR�X�N�Lw��7ʖ?�w\n��u��FNϒ/u^#F�er��m���ZR�sM8�
��kY�{k��kr�52��pU��)���`�k�:�*�j�ַw\�h�r�`�z���:���FSJh�G�t���R�[Δ���3��NK�^v�C;�u�V)��C�-�z_2�uS�茁r�3,|�N��q���U�h%���	�);�(����,�ڸ�ju��L4�����kJs�y�Y�<�]�fuZ�k������M�a웹yB�DtP���u�r��i��IS��tL�%��ql���_<�Cw<���@���p�/���؞����re��ܥ��Z��Se��fP��]����
wA����6��Z�-_{)�~��m�u+Y��y��*��C�^2pb����jmFhs�"�w�����6�O��y��D]+A[O]�v8�c+|]��z���n[.��C�;�e��|y�"���Onp��]>,`*�3�[�N^��f�5�dJ�t���8�U��,���E�t%uhP��Ѹ�Y��N�F:���9
�0T62v�R�=��
R�Q<�\�q�\������ٶN��Xt)�&���
�2]��@�޽��P�B��KM���j�I����s�ꡦ^@�X�<r��=la7F! ĠatkRA_C��$�7Ey�,8�5ãrl��x78x�x�E�}��2���<�mX���%.ŝ�8�.��",��s�q�y��+u%o�;�q�2�}{9�̙2LT�Q�J8��=�x�N�ohJQ=4p�8���m�Q���cU���ϰv���;6yU������x(�N�|5{��Ⴣ��ufYU�����c�K8��,��ok����F�����(��x��w]��pxumԭ�V�����\R�ְ0�z삓<Yɇ"�.�E8XӥsVV�g��]O� ��n�n�h��w�r�~�3<���"/W��O=+P7/U��u;W$�8#b]�섃�3�xʯ	���(�x�e�����3�Q��
��Z��m��-�j�0�0����o� ��^P)�G��F�,ŅG��X�v�%��/G�c0.��<��@}�ĺ<���wu��.%㺸et�z0t����vd��ہ�h�������Lv��]@��5[�P�OS���ù';�J���l�b_6�Px��j]���o� ��R�X�(��xuf�9��	�H��{��Ӹ�u0�{s#5>QZ��&R`F�°�B�6���8�[�<ۂ`ц�	 f�^�D������ʽ�Ƕu�g�al���򚑢�5��|�e
}��V���y޲�ɳ�L���C�f�Tqm\�ѭ�V������@wsÍ����Z����7�����q�O��G"�Q��et��|M@b�*��:�K���r6a�~K��Q�39�	�;����%�a�F]���S��e���ܥE�M����5��p�	-�p��o�n�5����}"�-x��n���߸ h�(�z:�Zٷ�M� ���fE�Dl��:ܑ�L��� ��Xgo2���Q.��a�yJ�z9>˨r�� o`T�nw�i��(Ը��n�A�C6�R�7��]��t�KZc.Dh��Tt��m�I�d�tA	����⦸:g�S]��鹜6^��V�k�3U�3/gW�����塱�D���/݌����4�>��<6J����٦�f���O����\�A�[F��{�Z�� ���ٚLf3Z�n!o�6ِ��t����mT�'M��8Ϻ��%_H�	7�o�)v�����LW
=u�	O��������އx4V���^�гo��<�u������8�KܔsDp..v�v�=/��MbeWhêJzoVc��r!1��$�Wn�v�hUl �I���J�}���������Z���i��wi|��}�eH�7�waJ��U����p^U4M�ٷ�p[#���xL���+Ժ��G�9l��,��J�\��.��Z3Rs�s)�9V&()�vF�y\�F�S�l�H���MX��/_n�����HPw�o���=b��x`�9|D/���'s�9$�8�l�띺א��Ti�.���i ��m�$��P;t"](���w�ZnR��f����|�5�eSݎs�x!�)���TxZϗa9{�d���u�ĄNBnm��n�p;��Gf9L򺖦*������>_s�'�h��]��������Y]g�֪�ֳFa��n����.���L;o.I9F�܄�l���]b���I-��א�n����I��uЭ�G7�O}Ĉ�{�u'\*�Q#0_&�-�{Q_p��F�Z��_)	mh6����蜂�+'^!ϳ��iև	VΨ����Vݔr�$����,*Y"�ɐ�e��u����ʈ�R̷��=u��'{:��T2kqV�2NU�(S����d�-��$jh͍����[fs���dou�`�iޔ'2���Q�X�)R*~}�F���D3�r��c�f��U��ki>f�8d�+�%Y9ɤ�̎%������
)'����+�WN�h���Q��f�������].��i�&��CER�%�o�eF�e�f42�X�� ���#�n�b8�v�6�EXʣB��؋��� ��m�^m�F;����m���|T\���f7�:]]*7��pf
9�MJM���%�J�k��T������%6�f_�dmvk�o{ea�*����2�d���_����բ
�l��	��.9���P�P�)�X��z�����{|/�V���%���8�b���k�J�X0GW�u��T��n��-�%�Q�;qm��k���f�p��A5P4�w��c'4��Mդ��]�b�%�,����"��n�.��.T�c{iɭ(��]��4��uz��B�&NXU�W��/��]�q,r�%]#��*���Y�m�#Q>�v��f
ܬ�D͞��4%��N�+�9J�>�k��퉴�v��d"��u���\a@�|o2�]N^��9�3;tn�(�nTN
k*f�IPu��7��t��Wр���S1����Z��$*S�"�w��i!o���8������u�T^�lUV�����u$o�I1�NҠz�J�
���ԣ�f��69��MT'�뭲��s�l]�FZ�M�;�v$9}۶xJJ���s1	�ȁ5>V��M�h�}��uV�wz���m�U�|�剅`��Qn�&��h����5�������J�Q�;0�s��
�֋vW�u6��qw�s*�f��a�����ue��F<�`��=e�ޛ��z�s��#V�Hخ
�b�l�خa����ن�)�e]�ǳsh}VQ�Lhx�!��R:l=���懽�Y�|�v�N]������-�z�0�&������1]w"3��lhj8vJ�f�ݪ�[ɡ�6�;R�\w��%����p�ӛ����Y@��'+�Yg}Hn,�IM�\;�L�ӡ��Ǉ.v�1��+�m�K��MvK#`�2�e�f����4E\%�H�TϤ��}�;���f_L�v�<��(�eq�����/��I����Q�h��sut��u��&o���l�x��r��YKJ���
�0�7.�Q�r%l��� �Z�7�� �d���ܬ�*X�̰���e��`4_s�G���яc�t四��Ӄ.s�씱ښмik*�zn���HFv�J8A���v��:��b<�DKUn�\4oek�M9:S=�sJ�A�ݴțG��km�3t�ڣ�������.�*}�Men�V���G���*����B�1b�Q�j��m���١fv�p{E��"����%e�SW�+^��{}��G�`�9��y�r�<��E����-#5I������F��ŒF0���c��qm�`³�����P��|��A�	ޕ���5�L����(�.�sѬP�E��w.v��:�ԁ��z�an�w��;�\@�vp����v�b���T����3{���/�pꔗh��4��������I�o_ƏG���]�M�ƙ�"}�V�5�M����)g��<h�_OfI��n�� ݎa���L;���_њ^sή��N�$U7MbOA�(�8��������7����Ţ$�y(�or��(���b��y�����}<~P�	TlH��ϱ!�m�j&&��
��w_)����z���u�I����e4�s1>g�O�0�����wu%�n�3Cjorg �r�Nk.�1�s�k�cw��dt	���8!��6+�l�3��V4n�u�a幸e\8�M��̹�ٝ�6I��>Y}�Mr��@�eJ��$Ż�˹ӭx��O�:k�<{���D:��;S�ѱ���홛��v�3/�Ο
���
��\�.�mX�)6b�;�ͦ	wk�5���p�vp)BJV��O躛\tgZ:�]ij�ۨ�Բ`��w��%5��97�ԡ�we*o����2���y��<bbM��n�U����/�����e���pi*�ֈ#I�5�L��5}4xD�Q��׏D3���7çL��"{q{��M�xs&8��Ɯ���'��B���e�����ƍ'fp�)i��Y�Y�F�9Y�����.U�r]̒}8�b#�M����3����[x� �7`ں�n�Wwǝjm݈�d��I�z�Nҟ,��h-�O��~�Q���ć�Q{=紤:՝J����]2L�d"�ͻrm+$#��log��r´�5蒵���87��D��]]B'�"��WZo���8�l��U��;]w�me�)%n���r	Q-��g'X��X�U*:ԟX������&bZ,�Y�~��t��
��c�b(N5Y��*�W�f�I�	��l�YN��\�T���<;�̶1�C���qǼ:#1S<,O�ѭC���8���J|��z:�R�:.|�=]XP��,�0��+��^C��Fʮ�#2�}����o[�V�8���9��M��!����ԋ7�U�l��j�1�6����7 ��i��g7���]5���F�h#�'H\�Ʈ���=�M怹묮F��v�#�3�@EƷh�E�W���
��f�jҸ��K�[g#&��;hڝ̒y�J��]�Ϛ�z�vq5����{��e�,,L�z�ɔ���!w`e�y�~[�4�ԻX�H�&�v��12�{������+;���;9�S_>IU�s];��&�,�o+�l{��D��*B����@^�[���:�`��ɀ�ç*bi>D����"\�ܻ�<Nm�m���l2�x��g+(��2�K��ۃ
�v9�rN�ƨ`�pA�c�k{���X�y�}tۗ�t��_#��v<N�,�-�����E�{���jJXa�8�;�ބ֭�H*������YH�����YrM��s���9K%�0fh��f�]�w
�\�R��&�i��A �m��k��M`�i"�w=��c`��,Yz�D�v�0�w|����Kщ;T�[��XU�%�5�s�����h[OT�3w#G51�{�X�v��o�gNE���>F`1�ݵ���j��ɳ�M���6�����г��鼱*�]<�!h�ˌU�2Wq<��t�^Z��(�Q�k��}���5�C�S�C�(^+F��v-�"�9�����ygoq��A�T m[Tέ��T�bQv�@7'5Y��DU����l�	c]��WԐ1F��S9�[�@|�ܡ��K��i����-S�q�z�Thj�m�v�|>�4�N�_"�'A�ۼ.�N�Xf�4#����L}�`T����R-mYz �X��[Cc}R�� ��"�m5��9�uѾ}�Q���L)_S�_e���D��V }p�Ӣ�s�ou�;"R P@��{&��RK�����ΘO�����ռ��aeg�)&]���$�Ӣ�ղ�Y4F®�^��4�G��B�#ˎHr�y�z��3��']�'>j�v��T�jH����(��,�b�D�q�v!��W�RY�/��\o��M��.b6��� �+&�ß `"�j�G˴�Y��7(�[��vz��^��x��C ���ok��Хҁt��6�b�#ݤ�3�]YG����|
knv���T��XZ7F��pbQ�I�;P�h��n�.f�=�:s1�`�Cu��+�Q�-E���(�NQs�8n#֡�X�j�y:�(e�:�D'N�e��c/\ɪJ;��;�7�u�#:r��'c�ol���<vٝ"�Gs�u:>�F�m�{2#��)&�:�r��J�J8�oE'Cq�Y�I��f��v�/1�X�뱊�Z�.�N����#��x��@ $HIO���������V��.��y��WA����X��u�-l��%�݃�{Z�-��'O-��/�4P���"꒦e+ܶ��E���2�6�G�uA��\fbˡ�/2A���&"�k6���R�5Ž�9����k*���xv�Pd%�*s�#�n���:q9Yt-4~�Vi�SM=�
��S�:��-`�]�_P] 	�(\Է'l�o�]sz�n+Y��"���b���P��{
?.�}l�$`u���ylO�����Z�d��[��n�pgS�wK�����V���d{[*u���C��і��w�O@��&I��m�׊+n��F�35]����9/:�Y]����h�MЀu��0ĕѾ�� 䒽�]��wg]m��ˉ�Fޤ���o�������{�cbㇺ�n+�1�;a�����)J��m^9�%�՘.�C�Z�lx�v�[Lq�e����Q�t�|�x1�O��ŧXJq�m_r]�nYr���1u�!�p��
	�2�gkE�Z0I��vc =����x�r�ґ[1�ek�F��Q�QR�Ws�T�rj�)軫�V�(/m����M��u�M�64[�gF��/�w��1E�=����1��ĩ��oQa�dNI�шaG%��s�ӳR�i�ޙGjn#�7ڹ� �Z�e_L:uolYU�3v]D�u�"X�0����4sL����<��;�ݬ��9�'s::O��:��aw��Hk{P,չL�&��^�%��Ǎr�k&�ԬB���ӗ�F�Z���1�A�_I�kuW=`��s#�Q%�2SX�%N��,���;-���7lD-�1\b���3	�h���۫�(��]آ�j
��S%�]k�q�f�{T�rM̢>F>�E�i�R�O�ٜe;x�;��H�����s/B���F�N��'E�Oj(��z{;S!F���B�Q�5�bZKV%V�o�fE]Rv�k�Ǆ�3
��3�8���@�ռ=U�Ϣ�m
S�K�:b�7ҭ�ޜ����AY!�h'���7�� ���l8�hhq��k�.�vpЫ�v�D���Q�:kh�iTYgx����M����u�.W�ݭХ��Ƨۤk����o�K�Z�je1:��]�`^2�N��>+��S5��5��Ӎ�3Y�]%��������S��y��ᤩ�sce�e�B�|/r���֩YǬ��i���)�2�2��%��k[|]��8�r����e&��+q�ǹݡ��{@Μj�ӘwoS��EW��Ӷ���v"J�Y�1ښ:�V������Z_'ZI�1�v_bA,��ư�5���Ԏ��	V8�j�L�U+w�� �p
F(���F�5w�+,�=��*Ǟ�Ө�û�$2�F���9����ڨ&�������Ľ9�K*1�Y|�X[�r�h��t7�U�:,�$��}�HB��� ���]�&���d��!{L�7)�x�f�$ޞ�d5۹5��ɽ4�pl�O�ǫxq'�v��g&U�bv��`�Qj�]≪1ͻ���E���^�	��L�-a@�ǉ껳�bH�4�u(��x�>�\'8z���f�6�rZwӪ���CV+Φ�4]��ؘQ�r����%�"�%����xD�A���b�Y�䊼x�l��	졙ե����mi�7V>���QH/J����/D�R=�e!�S%��wj����l����439�H���=w^M�����h�=3N�� $����Rڡ~����m�\�{,���p�$V
�FJ����X�&M<;z��g-��|�wchV5�^6�b������n�
�i�]�T�5s��L�X���)C�C7�v��b�I�[�w-싯�,4�U��E0�CF�99A�Sxb����'K]1�N�|+i4�l�[ܾc��.7z��d�h���v�w"5z��%�g�7s{�6{�of��o	ă�V[i;.m��8��%��RN�QI��A�\�f#���o���{��AWm��ky����Ƀ2��^Qc#����M�h]=쇮��p�1n�kY�Gp�ɼȦPu�q�r�[��}\���\��������Dh�,T�z��@���i�[���b��j����݅�c��-:��lH��m��	4��͗(\�8&ܾɵ��L���W�����N�=�B>�Ƿ�gJ��*7�e��O]Y�2�,��j>'��ޫW�>N��ٗ
kQ���'jUb}��_m�&���a�Fs�h_I��/9Y��MM�ka�C��۹�����6e��Eώ���|;,5j�v!�M�w��0wY$�϶��|�a:Bq���9v��,�me�=$W�r�K�r����ӷի`�����}�\�(t��%����f���FJ�����{Im�7ᖾ�>=�9�n����^y�+���mA<�$��b�aE�d�N�v�b4�=uخ�o_d�3l�r�O���9�Xy�[D}:��Rc�÷y��ie&����Q�Y&��+N�y�U��;6��7��A��E��5�h�e	�1�0�����������b9#�m�3So�!%�c�.��̎�i��Q���j��W	Gt�lvtݒ ����m�˒҆�矔���"/MB]�;��/ul�V��e���m����ᮌ�r�C�X4��d0�g��n��j��Ӥ�Wϳ̗����U��Q*��	\�v��\���>G�Wj�`�ی��+�#p�o+�%�+����᫫;�d#�fA	�<�{S~D�g�f��
��7�-�i�
����[t��}�mVE���XlWin�:�J�hv�P�\X{8��¯�/f^fuj�OtӀ,��Bҏtvn�X*ŝ��c[�7B�F�פI��c=L�0��0�=�Fx�Uy	s��W�;
��;����.8��џwC�e^���֏��6����t`�V;U��Q��і�b�#N-@�Y�C�LZy`d恰8���f���Cӕ��5W�[���3�E��Wvi�,�gvv�L0�w1�j��>�#��8a��R�`^t݈3��
���+G�s[�-�N�`�������ɬ����}}�Hm��
�:b�� �Q5*Wn��@�`���ʚ��X.�(\�׃��f�6C�r�ܛ�8�a����H��c�FB�6��)��aQ͎uo4W^X���"ҵbY�e���J���zy{*���f[��V=y�
���cUΖ.���M�@[�\8ԺG�lrv��ft׳�4����p�i�qei���	��@7�h�
��5�����t%�,h����kkG.`Ҷ�L����F�Of*��3='���5�w��
��M��3����c���t�7��	�  ڎ �׉��{8bJkE�d���g*.VX�&ZT�j��B��R��:���[z�=T��Y�ۂÛ�5�F)����`ڴ�/1y�K�#}_�>����Gz�f%�Ō�s1s"��sF�&�WB\�=�ne�(��x]�LH���Kc�\��h���m�@hv=e�x2^������o+
��!14�Pn�5�s��h#ؑ�B��h����?���;��H#c�Ǯ���b�#�÷kD+N^}k��J���J�
��&]A>P��2'&70_n|�>e���Lc{�|�k�/�k���/OU�e0��̆�"s�<FH�XO�͌z�w_>�0��I��3k*�4�Jd=:���F���-h�ոk���L<�V6��v.ɉ�^�;�:.����&���J�V�f�]8�#��%-²�e�D�W�����Ĭ��iPY�#H�nݽ�yH��.��� hӨ7�4��4o�f�]�¡f�t�������ݘ�s�h�w�p�pp�a����.�������"I����'�!,r���
�Ys�ۥʵ%�
����9�Xou�v=ww��k���^�:�Y0������-����e�(μB~�zw���|ʢh҈�ٽ%�_p�{8��X{����f�����qs�)��ӫ[Q;�������ʻ	!8�ʽ�cE�<�e����1���88#�wZ�TÖce�wm\w���\k+z�>�|�R�\���5�n�U
��&�7�?���;����W�A�g��w򆰓T��C!ƍ:�qZ�ļ-͜���Ʒ���-≶��ny�����ҰH�YGc?I�qօ�W!2����ݨ-BN*Â����SNۖ�k;*&���;t�!բ��[!�ܯ��M�l�eF�^]b�ic��5�eXNoq�n�ciZI����Ww՗��0o.��gP4PYD,���ܾඋ�S-5���x�v�D��ȉ���O�ڝ�T��	Љ�7fhS�*���+i�Dقj[�l8���X��;�uw `���2�~�)�/li6e�\:X��<��~h�WL�q�#͌�|��Ň�gY�>ڐ+�Oj��*��o3�IXB6g.�]�B��җ��	e�k�;.���U�2Kw�_��h_A%�hCm�b=w�c7�=:��o�!2��a���j���֔̄��©AyB������&�(��q��M�mI��K2�K�4�êqp�$Yy��׌#Gv��PC���˶�cc�qP����g��:/<�_=�xC�UY\C��'6,*����<�*x�8Իް1�$�yy�\(L	>e;]X��B�+�:��̕`��\���v��<õo+\ƞ]�ͮE|(���$�v%��2e�`E���aS����2@��B�E$�G��+Ȧ��T��-<��=+��Y[�n�~��G��i[[SɄ�pv)gq8�Y6��p5�l�j��h-�4���Nˬ�Q�^���M
h@ӱ��z���rc�2�Ơ��j���ـWT�9&�wWpdejJ�K֮v�j����]{���T�ef,�튫�����6𝣮���l%�Q �]҆)e��һ �l�2R�M����i0��{Ŵ(x#<_�5�ˎL�o�/��}�(#��.W��zTM5(��T�O!B�$m��6JTn�`"�K]KW"%a���HWZ&�.˺��d��%=���P�������VU����n��!���C[R�I�N�t���]�!�ϻi�[o;������@��煢��E�4��3����g��g+<�<���L�x�ZwS��QЩ���h���5Ԏ����]�B���j�y��no+hB���i���5��Z^�"�H�|7F^���}[v�"��1��E�V���U��x�r2��%a�s�+ 7��PeH�1n�KK��o<���Zu�mNQMSn�F�ķ�]��W%��3�c�r���\������
������]v�p��}�DS��uMy{�r8b�l�҄�����|[Tvg<�%�^I)�)��T�f}ԐW�\Nw+Kk���J�Wf�Ĳ��t�ܡ8c�����.���T�%/��:�+x�ME�v� �T�,���h�yr�����!Ί���AK�k8�ѼrBpVvZ,���S<��Yr;KN�2į��w����y
?{_��0{�eh�۸=�iq�⯬7"`-��QB��o��(���0I2�+cے����;3Mj��*j�a�kWR��318F�b��p�y���[iv�K��9�Guq�����B�T�|�bL�YIw�J�li��P�z�T5�N4N�b�}v�Y�c��Fl���u�i����bmi���g\]ϖo#^J�7o�\E�{E���z��T6�,6�\0n���T"0�Q��D7[QG�'��])�n��-�z���rm��dT{��7rk��8��r��l����Wwtƥ��a���#+zJrf��O�ʸ��%X�;/S�й�.Ԕ�m4�KUcV��/v?aѮ�hq��b�o�y�wxbXՆN;M�Z�;��)�^�`���n	`���V^�2�b��J<kf]���u����"�ӄX�)M�>�YX�K�q��7�Hbd���#zFn����,�p�]��U�>�-[�{Φ��8���~�p��5lծ�8-H����qVT��KֶJ��E��j�˂�N�W4�a���T6�vm#N`�	j{d�m!�@�rJ,���8����%l_Yy�����Nw���Kiݦ���I���|�~�̋������hr�f�X���j�a�V�9�9���[�X�1��:-fU�j��(�!\��ήM*9��z����A��lh�Y0j� ��qE����3�4��kT�t��[ ��f��+�s��-�.��|N�#�kF���z�w^s	qk� ��-5����}��۾{���7+wk��o�Qx�D�����jk4�b�JD"-v�b� ���˽b��_u�e�c�v��pȪ�^��(������M�@���Vv��	�R:6�n!���._nU���+R�l5�V٫��l�ܦyp�eJ=��.$o�eڢ9�%\��n!�ـ�Z��;�,�#�8p�=��Rr��Pabi���.��]�f�����5n���$n�����n�&Fܮ��g*��.�ݡ�=���!�ɍ�_Wc�i��2*���S��=Ǧ�IV�ᑺ�1��1���AuhW^�,��h�[ǅ�tɬժ'��2�A�tW��'%��[Bk!<�5yϘ��f[�U$gyA���+����m��[�W���92B�\�:��&�l+��N���U�^�(�̊*Xr�e�k� �%ǧkH�ެ��k3�ģ�;.m�Dv����h;�{����XFB"��"���{�����kv�o���Uu��e��P"����x�W
������ٶ�P̃���Ғg%B�����{;_���?	�ߛ>>f�����RBH��|G_$�@�:��9HKw����nT�sI�.E���4r3��0��K�HӸ6a�C��+��ݢ͡�ro,Y�;/��%�G*�dGeBGJ�ؑ�L�X9���V�����۝b��V�s�Zƌ�i��"Vu�&f+�M�ñ�X���cViW��$�*mqȦR�&Q�˄[F��K��>-h'�ڶS�Q��f�J'U�=�{�nKJ���_"�U�x�IzA;��|}���F�!�H���k���5i��Q�����L�{�3]3n�+1P��[�6��b��\���p5k:�Mv��(q�|�bA�ݵo�6n�L�৆�7�d��n��359.�'�i��/�a�
յ��8&�e&H�B�7"�}:�ʙc	�ހ���pѕӗ8�0q"+i�b�ҝY�t�b?�m��7|6^S������eͫ�9���j��hv�(]9͑COe3�ӄK3�jO�su_3{�o���r���px��!ZR�z����բ��'�s�/^�o���/����m����i�:���\��x����3 �1 �[�y���2��ZLW޹�dّ�+�*r�������UP
Hm��?k+��ƶ,���dQ��6ҴQ1b��lX��XS(Z،w�"�*QQ��b��:�*,WT�++Xڍj�QbbQc���Fڪ(2��"9EA��Ŷ�����EH���J����(�E��(ZTr�n���aF�4тbږ҉����Xm����
1UQn�+�(�TZԺk���k�����Q����R��ь�*"�1�(�U�ܥը�e�����R��FT�D�%eV �[E��Tәb1KB����J1q��uh��W)E�B���j�Tf�Q�*:J#mT"��Z�T�LV��*���� �A�TX*Ѫ�,AjQXR�U�kiYm�3H�2�Q��Z�E�)`�FY�-j�eX�Җ�b6�ikP��R1D[Jʣej���Q�Aeˊ�]4��<(5�@��]�d��1��W����C{��:���t����,n�C�P���杉�S��+��������t����q�?��1��t�z�����V��L���ӱ굤Lg�Iܫ�H��\�G}wx��S���ߏ��X�j�q�T\X;
2�]#c\��Grت�Y{<�w�F�)4E���}*�������Є�NA"�H�D]à�����uU�I��m�x�:w5@�~���Yy��z$^K��T�A����CM��dqU1|��0�[̼Ɵ9�8���c�1���z�}P��pê��3�*�8�Fʋ��!L�,j�r�&شftl�m
;F=aHP��Re��w0HL�q�D`j(eз�ӱ�=]�L�c��1Yj�[��{s�����/��66��F�L�"\��T5�3؇�{�ڋ$�Z��QI�/�,v\L�}�pDllc�}�^�G"��˾-�X���&e���&�d�
7I^�7�E��o���'c&Lp�U��Hا�U�'?�D�㗊��R:��y�ŀJg�X<J|�e�T{P��9�`ߚ92ZG\��"�B���&:<9�� ix��C33Y�}��^R�89�(JY/��4lN��m(�meRU��Z��EMq3�,�lIl���s�#�9��6F��WH��`�ݾ�g>�<t���Ɲ�
B��wV`I����۸�tujY�.q��ލ',�[��$���$*�ܵP�N��~V�b�|F�F>��4}l�W!Bߦ���x�#��(�"�����K�E�����ϋ�Cru�cci�]~��^�C�H������q��śtVeJ>�php��S�y��G��k[��ǈs�8�W@�}q��*�E���Mg�f켿#K�絬���wv�r�nBr�J��Q\��A�ba�����Ʒ��V@~R;$u�)��$�..�����OH[|�E���Vy�U�@:!����W'9`��bs�a1ʫӋ��t
��		�j�!ɥ_^�>S3�ڻ�9��
v� �����G��(���L[�qL�ʱ.:��F�Kg��b��}�V:SOK���;Uu�=瘺R�X��.8$�8.vVU�;�w'��9Sp���J*$1+�9�D�CnG]wn���9~���jڗur�cFс��C�뛤��`�Nnh^T}�i�u�3x��F���{z�����«m�������+h��+9�`N��e�C���8Ë0��0�o��@ׄ�~h5��>��%�۔2�w^g.B������m"��6l�J�Ϛ-;�
w�:l�ǎ�7z�:�4Br���z�U@�e�tT�Z9�.��:�b�-�Ɗ�D����v�%P�
���ǀ�^,�My����9C��G����o8sg�8dY�AW�"뺗�u�Eٮ�%�C�?/�'�ʫ^�ҫU ��Vf�Çu]�R�4!�r=1�^8�:�\Հј5$4!Su�S�O�U���(2���Eͤi�����|��Z�)p�Fm]���~��	u�
"���o�u=E�9�
 �MYC�m.�[��R�lY+�c"��V]_#�B��Q���"b��Fy�$c����TM�rѴ0���}�2�j������\� ^c(A��Q���y:F�\�)�dMX࡝L�H�y�U�O��~�e�h��!�k��.�:�@aH9W�z-Nztu�{�z9��q.��]����gzj���V,�[aL1BzSz�}:��O�}�u��-˕4�f�ÑOt;ܔ�f��Fp�<��~n�d�!@��A앆�`�����t\$�[�ov��e��J�q/r��p��i��X�[/&c�)U���lW�U{�;DE�R�fI�P�n
I�7��9˯P��)��	��V�aN��#tZ��ڗ��B>
� ��)yz�ش*M��s�sN��9\x��� ��+)t�3!� _;�>)�WNz��u�^z��KB��E�6�W֍ב�-�55L��4�^$�.[�63���d�2��ڭ�l_��g>���i_f��w��2�5s�]��ߐ	G-�-������V͗���Pl�
��o�vu�*,c�7�TL���OTYѥ��~&o=������3U�^���Q�ֹ^�R5�x.��^ �4-&���Y�����鹽v�(0t�"�ש�
cr���@�r�x�{*�8�����u��b�C�v��y�Uk�U�cH�z��M�
� �����n����	���`]�Ǳ�����s�ܹe�����7P��s[ 4Ί�
q&�<��N�@���-�T���)s���kn �%a����G@�m�1M2�;f8E�Ezh�qr�l8�Q�`��E����w���!��Y�b��'h8uM�oi�By���P��Uk���
����j����3�g$�^�iֱ��k��0��>�EgU�cG���R���k&��$���R�]e쵝�o�\�/�}��p��># ����f�6�o��#E��9�v���1{�|8w˵Q�rjYB�O�Fߝx����XO�uѣ!��8�3���<��ϛ�2r�4�焠4r��@AS�*�^�կ�{�K��x�F��7�@&f/QxgH�����2cm���
���4J�u��������ǸE9{��|�zc�
K�b8nĮyk��y}�if^��j�N�U[���3.F��S:�>=��s�B�y>Y]3J�{.2�ۛ=F��^[M�9[8g�=�o��V��B;�$��g Xe�P음�ꕁ�Q1aH�U>�;B�
��
����5�_%��w`�b���.ĩ���i�p�R�r�E���j$���Q9��Yӑq]���h���"G0*�z#a�p���[��M�W�ӊ����<霊s#:c�����M��u�C�1���BtGL臞�Q�<ʋ[=.���?�76�{��$WM��AQ܉��A�vg=�G��z�����#ꡜe�3���$=�`M+^�W���%}�~�Ĩ8���P9 ڥD7.gF?S���NA��զu
�T�Uv����Ȍte���Es���O/#��z$X.2<iR�ծ��ݷ��*�.e�l@�M�xA��[�S�*Jo& R���*ˋ���<"�	U*��8��I׷k�[L��Y�qlQ�|�Vz��x���3�L��N�
t�y���j(e?Q����������w,��H(Œ]d;n�rI;>k�d�{)�� ]O]׸�xy�T���ӪfM/��nk��i�P_^+�,�X�>�s���� R���q�A��|����Xf�.�+o$Zf�/pf6x-	�"��g��
{Xm_�)Z��]���/2������oL�CR"\��5wJ�awx{���Ɗ���V�sS��~�U��_Xo�~���]G3��_ݾ܇����~�u�^X���
����Ѷ�d��=U���>��]��>"ꛝ�u�Jl�����Y��B�臁��_PY&��sd��4Ng��n�n�f�,V��d��g�VF*Ԛm�m�+S�ŚB=##`4�s�hڷ紳4{U�r��zu��.�k��Au�y����ķ��ת��H��g����0��3��܂gX���襞}~��X����ySz����Q�а�~�G�OC��laA�
�}�n�v��9ΜSq���;�+yU���6�[����Wd�4c��B�.����X����m�w\���i��z�ck����!Z�2�T�(OE���;Q�F�k	���a�O���Ve��u˼�[���]uZ�1�\kE*��W>��8���r�IXql���{��0[��1���V8k1�i>�L.��F��g'�ݾ�+�ܥ��<�*��3R��c;TX���S���Z���f��;P�3Z��t�C'��g�r��\�L��)-���q9��r1�u�$������F��r�mHQ[;�}�3�*�|6'rj�}�/����+�Ӂ�O8����s��I�w
�2NKs���R=������r�����⊉&�{�t��6���w�5,x}p�jׯ+��C�r/Fрrq�vDu͊O-�:�'6�C܂��tqθI��]����md�>MT(�x�<|u-���V���<��F�Fsv�-���vJ�TF�~�ӂ,r�؊��J�H�9!X���"��RnY�}���'-7�f��X���R 3�\մfIhEC`�&k&�灜�@]���2/7Ne�S�E>m���-F��1�9�FaP�t��A�6}�-D�7�C�R�s�sr�ƶq�f���b7�Y,\� Y<�c=Ee�p�*��)e�=�&(�}��Ů��ݐ��{�}������Ql�l�ns��U�2��Q�ۏ&U�΀�^ȢU@�=ۓ�α���> .jH���xk`��#�۠0������8yTm���R�oƐe�SA�Vk.Kf��7�{�ѺT�^���h懷0>Y�iN+���m�`�����7�����:�۲�o̓���SB�;�����[�,h�=9�֤F^�&oؘ��.Ռ��3��4.oH6k�O�ӆ\��*�6tW�
��Hs�������{5ν�9X��ؓ�����⣚�J�\k~����	f�^�����qL�\9�'K�/D�7[ͺ�k���(Q�UME�ʐᛚ裲Ј)��ƚ0�%V�wI�ќ'��V�c%l�����Jg�u�}�^��b��syJ/-�/�.k[S�{�C�T�)�9�nA��]��ȷ;�y�;R��1�41x�����q�a�KrG�\D�	שR�>ŹUt2r[�����ʎ�>9Sc���Q3:��r������(p_w�:K�GÃ[
4��(z�n,C\�	�@K2p�tܬΝ��ǒRόJ ��jp��Ӿ{�/"�@�����uto��tiu����R]m�޵�[9ȉ�'��H�mSɡS3}H�%g��ʉ�)�,-��4P��O��������}srۧg��r \�K �N$�@��I���ΜddZ�v��kZ�B��;4}��nG@�m�1M2�8�����@����p9Vᥑ�@��o�(�%�_+�hF������1R�=k
�M<�Ӛ�u���C�ɞ���z�ݩ�#�ӳ�a�-ח�+��q��٥�˻C�h�w7IC��z�:+�"Dr^�빃�u\��v�P2�+&�h��6��/��Ԭ �r��{�V���+6X3�Nezh�%���7`�t�����붪Ø��j����x�R˯Rk��jY훍�3��Y���PΫr�$z_�W+� <g��xe�}��o;-B�[��8�#b�
�R2
�r�aq�~-���F������M59�ĞZ�B��fM��E;(mz�B_�V�'�̓�XO�(�z,a�#kj�-P����K�@AS%Z�~���
�O8�����+L����# �ڛsg�®����:[��W8�ߙt�+�P�뛫�̲�̉���F��6���H�,�v��׻5�^.<�^�b�j�nk��֪��J{P�_'a�uJ-�y����j&�h�r�_�U�ڰ�7�:�����F���Dlp�p�A��s�6�_PN+s#��\��ғ���>-2ige5Osx��V0��+��BtG�ȪQ�<ʋ���x.����a�"0�Y[�����R����%���W���!}}��hz�ZV���	�88:�^��<���+;�ͫaߔ�/����\�j��HlumbOۚ���3[{e��6�Q��}s�'Y�~���enf�M���V���"P[Q���׹��\8����=Wr���8#�;�2�'����u���	�.��p�޼��$�\8��m��l2G@�Wo�����U<ѯ��R�H������a	���*Et�V".�rz�7N��\٤�(T;�9���U��t2)��v6oD���T�Al�uQӎPBA�ڎpf)^��CJ��l�����9�d�
R|0K���eƇD���i�Vh8&8*Ԣț;o'�����A<�;���T�c��V:��i����b<|��oV��>�������/V�MX<�g��\a�\T_AѴ\�����6U���P����d����vq����z���U퀚o�u:�c�o��9؟c����t�a���71�o��y���G�mL"���-�;4x7c&H��{K�F�>�J�x)9�/":���p���ٝ��5QIo^%6��!�(CN�o�WYw�,����{��l��),���Z.��]����{sD�ô�vk�2\1
!r��	���}Cfh�=����n�#�pָ?ql3�t�I�*�6+\*��|=CC�C��|�m�nG �:��6�E-�fL���l���{��k��0�����atVΎ��=�Ĩ:3���)�čxT�i~�Z��$��⾨�+��ry�b�,ˡFJ�����5��eG*Фs�Q���:�/�܁c�Fl�]�K]�w](x^`SA���4Q7ܡ�K�pR�������l�
*��[�����]u2�ł5,k�-�iG��n����˶( �Jl�����`仒`�����8ъ��S�7bk{]�w�7Ü��S�@�_�Ѻī,��6Yv�JYC&c��Ę:,F����VWӎ������&�i��!�˳��5��(Ы�oC���`��X0`��h2r�f���/�b����ԾR2ȅhG8�N�.JM
�=]�n��%er�eKUƺ�d��:�)���:,�n��1���}�c��\j5�\�7�N��ػ�EǛWa9�ʳ�-�'-�wq�K�+7�%�r��ֲr��*U.1�1��S�d����ݣˆ-<�	V]���)�t��[y�D�WJL�b�jn���v���egX��i��AʺG�eOۃ�C�Ѫ2�$IC)!�9S�V�#\���bA�ha�K,�푽Çj	4nكL��	Z�(`'���fK�w�g�}n�Yw}6Wl�A	��!f���E��a}˄���Mc�H0�.A��Ivv��{��k�=y�Z|<�Q	W�7fs�h��Slչ��:��a�S8���c��;9�TT�a���7*4�,Ϋ��fM��f�����N�X�Eb��gfc� I�� T�@ᣉ �Ŷ�4P�hl�p���XMo�T��� ��콸Z�����[)B��S8����'w2ju|,k����P�.�	_\��{3����ǇsxP0<�NxD�	��ݭ�~���M#���Y�V�43�f|j"����� �+�R�Y��WX5������n��.�+q����p��aف�f�ut�p �:��[J�-��	ά�B�w��%��-����U�x����!��!O�+�a�F��;�g,ag(�waӮ�Ѡ#x��+�3���[��w\6�̌�<�w�u?������S�)W�kcٗVj2=��d������C A�Zzv,'����L�B�ù]c�:�����h蕗A ��m4y�Q�m���䫏);n�rdR��'�,S������BS��`�.L��UxZݸ�IW�oi�
��r����:�F�<3�����:]T�l���AU�d��'�np��E�������>���)cG#r�B��YäujFQ&N�P��6��VȭI®x6�^�Y�e-�S��P7e���ܵQ�`ab!&3��!�^�c�s��o�q��{� �Va�T��9�4�W	�y�
r�����4Pg��@I�;�X�2�O�k��e=B�칰���-Z!�I�;B�Q-�gU6��wW���,
i�|��ev�ovP�T�3J#J���311�Њ�̕��*�KDE�UA�����Z�J�m�B����(�H���V�Z���KX�h6֍��5j�孥�+iPTYm�����mTZ�r˖Vb��6V��1�Q
%[[j���1���mF���&�Z�\�m���`��bDEPUˍnT�V ��CY�cjbQ�+T-)[mG-t���J�,U�-[XT���X,T�\WZ�[��,e)Vj�#�R���*�ֈ��ZX�W)��liJ���keQ��ee���YLU�u�j��pDFZ"QEQDh��J��эk1�#��p�b�4���"��Z�3*i�堙F�.���Mզ��iebֲ��q���E�-�pUq)K+
�DZŒ�s20��K!x���+l�V�x��o��j���oW��z�"lIWB�ַ�y9`�Ŝ��t3z�j����ҘX��;���|�X�a��k�5�6��PeB�*^1@�����+.Kͥ��gM%��R�[�P'��Q0�*��Kl����KPs˃��ǰ�;z�+d˼���D�;J����P2��*{� 8r4:e���P�+�9D���̨��wjr�q�J��](L׻���tu�s1�쪰�8��`)�CR�U��w��4Nb?z�ND�ɈRC(�7�RX;[�~�<�ٕ8��5G���^/������6էϯy�z����`�RE&E؅] 䜖���*�W��S;��l���NLPvpe�
sa��Z�_�$m�B�{nQ����(�眎Fрrq�vQs~���J��pg�-����r�>��� *]Y8O�U
�,\ڗ��>�:�j��r�S��F$]����X�M�kei�t'�,^�/�=C<Z.�tJ{���>/�3I�+4&G��x�ٚ�M��\$�S�@fp��h��@��= ��M��9K�%��%���L��|rf���uʳ�`r�W)�ܓ1DL�h�w�s�(bĴ%��+9�p�yG+c�vt�]�u�M5?�o�.ȼ���͆���Biҙ����4%��z#������ev�r+m��bmR��ظӌ�$QIX���އ��Q�oV��1P�u�zu���UԾ1Y��=Sc�B,��Ӯ�����6+��]C��%����f��7�!@�49e�1D.>�d�]�Ս�{ó�aꬶ4��bɪ��M��>�@�t�l^ʈv��x�ʼ١ܷ��)���qSYZ֫���}���8
�ۗ��*��#�۠3%+��z-`|��q���{I�c=K�D�ݣ��'&�׶�!��lU�ة��aXɭ�B\*��+\�$�jݗv�^E����8��X� U]�P/�����
땦�`�R0W����e�������=�C�}&G{P�21�P�R�hL�FR�
��K`��U�^ĥ-n���<��%�]|�p��`\K�S�\��WG_�2:M�H�L��^���n�����Cߺ����إJ$��aU�**�Dt09�̨��u=p���e��6^gT�{��GD�����P�ド�a���X8L�{�#�c���i
�^�{^Ҧ�*1u�U�e��dQعV�F��jx�����o�}����%z� @{ז�h�f�Ӫۻ�pF&��.�����vN�d����M�ML�~�`1���f ��Q�v�ls��nWԗBr�[k��j*ga�8f�3�	��t.om��d�����Q��^��è�����񇲣c��cőF���K�v�t�j����b�r�st,AR�hB�)���KE]|H�:7C�C����%m3�~[�M�č,���db��r�ɗuH@g�k`�:*l�N$��ة;9���%�P�C�	;g=\�V�������t
��7s�P�s1�.j+�@5]��w��gdw,�>��1Om߷�b��ٻ�N�C�Da-��i�C��h!�j�x-
�1��E�9/��} B��"�Y�a��a�j�]�y|��A�gU�a*�qKVf®f0��y�����o,�8(�{��W�yֽ�*FAV	�g0�ؼ(�6�{g6�8�E��BS�nS�)�*��x��"�j�2غ��3¶�-g��E�v4w_?pBx�A$*��}V�}�T�F��_B��ΚS�dt�b��6��̗**��Ze8��b_|��[���ɯ<#�+�����,2ˇ2:�#y#�+�f՝R����`i�qp�z�0��G�)6�K��y^=��������Ec�-Io���(��Xս�
�[ ��Ud"M���J�Uޕ�53��K�x<�녋l�����Ms�]�^�2�o�4���6�Av.q]E�䲟I8}�e�iGI�99nm�G�U(1Y�\+D�<+p�;�J���8W�J�r�E�������oevc8�TK��8HF�c�C�
:�-�AR�@�C����LAt0���Q�-�|0��r+���P�c�EН�:!窔z�y�>�z�����O���}R��Uz����j���ʅ��0Z�sME8����	�
g";�������V��x�.FN%�J~��t��z:����E\��@�7Nd�~�U�F����H=[>� {d�i嶱i�_�������J�����9�8$vK��T�A�zY���]f���$����3�Y�S@Z�#)����JH�.�9_��ܸ�:'[L������+����ז��׫;l�V������/�oMǈ��&[L���U�E�z��2�~S�L����O��F�x4k!��~^=|�o����ԧ�;6,ĺl'�zƗ1	�b�P@I٫��|bdU�a�/ѿ�)9ؗ���D�e=������	�Ȁ�?�5S4F�����k����<7�wa,˝|q�=㬿q��G���`wn���}vzv}n�����*�q#���Ӛ,�Ј�΍�E��8�����+E�S����H*@Ю����(��f��΅���y,���%Iq�	��?|�W�7/���ق_����P�C��Ohاҕd8����̡:�E(����՜=����R���1��0�=��o��l�7�L�40��< �Y�8OA���De����m�kA�8=Q�P���P6�]�Px�ϩ[�����ޡ�W�βU�uI��vj�b{1����Z��ȹ����ъ���^�̆�Y���B�LY��ܞ�*	��z1�UшpJި�JZ�ш��u���P�E)g��ᙛ���ʚ�=��՛��G��)�8W@�l��v:���]��j,eV�mҋ����kK6ӫ�M�\���J7���D��J��y���	D��lu8t'���"�DN��G�-�tsStg�\����U>[:=�WGX��c��]Sr�Ԇ�t
��		�LL��J��E�w3ۙ��Z�>����o6�(�������L�ʹq�5��n�MX��l]3����F���7�&�"�qW-�; �G�������9SU�D�gv�d��{^=�}��X,6��u���ƂK,tr��}�-�*.a��f���9d�ٮ�~䫟���mߡ��74�엝�.M�NL��^XǕ��ކ[�?Z�;+{��Ӓ�x�H,�]]6;.�b	?���\b��:!�/���+T��k�{�X�[CJ��H<�ƧՕ�`dc����7V�7������UZ��p�n�w����p���8Uz�>9~~���	+�'���Q����f�Ɏ�y�% Cq�b44 ��z����-f��,W�~���8��N$�6����e,�s��LJS0�&@dC�5m�RCB(�= ��M�*R%@��lN�Z\"�̳�{�E��r2&���1�P�t��6��̵jq�-vK���ι�!ݭ��2�6�$|��Df�P�UĽ�b��2�8c�d>�,��D�<9�M��Y�b����M����Y)����cJ�'�O?��]B����	����<>���������0��\�+�9ZƘ�f2||�Q�"���ᭂ��$tt���U�N�c�Xu.KV��욎�pR�@U�{�ٮu��ŝ�lU�أHO%���>um;����N�c�s�$F�Q�s��qb':�N*���t�B��"d�4cv6ܡ{���4(!�[Z�{��kl��]8Ӭ���l�I�J�s �{�X�wu�=��3/�)�ܽ���/��y��ݳ���}bR2��,zlb�[Y)���[9��G�<'s��T�̇�A$�ݟg}�z͎.5���4�@�*=L�V��_��6����)[��cV�c%l�����VWD�+ݖ�삨��i�(�����#b'�Dg��p��:�͹��v*s!㮋S�t�Ժº����\�\&�;;!D���U@���R�7ŹUt�2r[����ڳ%⽷�+��BW!�D�8w=Uة���/��C�|,v�%����֜��{���o�FXk����_��J����M�Lj�ʛ�*1!��C~�		��W]�q�u^Y-a�{�j��O�5�c�yJ:����Ȥ�����<�~*�"��36�Ĉr�dK���{O�o*[��U%6#��u�;���2�=s[ �:*l�8� z s������A���o��p�`�"4��t��S�c�Jv:Ci������1�pZ���vx$ȿF�����
{D����n�o>66o$�n�4Y
%���F�J�:	����gyds�y�g��r�Ҁ��H�^�,�9g�MX˵P]Oy����
����_E��Y�V���-9����b\D$r�:I{����9�	��e�e�5}�k��Ο��i<O����'z+�\�n��ܪg��^�����&uٻM2P3V鲆ٖ�2hp��cà�{��ًv\�8�c2K:�;]~��]
oybs�*ϗ�T�e,E�P>JǤ\,m�:U.�''�����%�������I�$ʋ[���&��B�H�#\��ᾃ���৏���Cs	q�5`�Xܕd�d-��w��S�qW���6g��f�gx�
5k�Ʃ#�l����G�5���n���n�����\XuCrv04�T�Ԣy�	�K���{��o�@ְ�O��#ڥ��
T9�2k����E�	�p]WE�p_T��{.��4$ĩx=U��l�n��5�,"pu3�Ã����wS���RCz�ٓ%���0neOT]B`UW�+ўh�J��:g!̨���T|]t=� �[p��cv8�ߑw�z�:q�ԇ������i�$Db���X�ڬ�g�YP'n#��yԭ��ŭ3W]��w!l����]�g������J�l���|�V�`ٖ`;ۣ3C�Ot�\�f'%�L��#�(��n{dlt��Η�X�y;5�w˗�]��`x)��{��'��ˮ�rN��!�#�̫�y^{���g+�o �Ƴ��EɛW��l"��h���v����È�N{g������+F��8�AU�j�h��_=��˽�S�b�/�>!Ey��{��rpN�m,8zu^�⧜z�fv��_9����U<�!�s`d�
R@�p]����P�\_���j���p��H�*�`��Y"�����J����V��G���ES��������-�Ef�����WG^�����(f� W��@V�j��T�}���>�E��D��mf*k1m�y}���U�������H[F2hp�����M׺�x:by/��s������c;*�6��-Er�����Y
=iT�!�u�[tvk�d\Ɏ�hV���-M+��M�\�5
x�{!�\|E�s�ͣF�Ӈ�L�>��N�9�`�h�>�5�-�Sdӎ_v���۠Ez�vkD�m�T7Ɨ�/P��P��@��O^	=�mX��9�t[���y��g��m���!.�k�v1r��"�r"憙p�SV�>)PnCw�5mf�3�&`Q�j)��7���x�y�j���SB�Ŋ�96*z\�b��Y�H�.$f��#�d�^(K��axf����Jҵ}��è�+i,��
˫\���*���I���g-h�]�:�S�\#:�+Kpt��/�v�����W�Nq�.�$x�*�\��l 4;�=������']��E�]1�.�����&�"~��G����7�5|4����p�AyiS��~�m;��swI�g92�Fo�����z�&a,J�S�*��bTD'#����쐭M�-�A�: D\!8Y���z��2x��L�7~�H%��R��糾�+��Ҝ�v:�n�mH�)�+��Md:gx��{����bgb�WW��57�P�g!�	߸�3�*���m���sĩ�5�m{�5�p^����UR
qS� ��<ayO�4�l�1�v�4�������E!�3��1�P�m���V,�q��0<H):���g�l������N�4w��b��W�<6� T���1��]QC{�l8¡�;ۦ�+:�S�i_̞&'f�4���Y4y�Mr��<a��O��=T����Qa�{a��'\`�M���K�;��Vv]Y촸e,�Lt2 ��d>��i���Ci�z�*O'{��d��1/)Ru
Ɍ���`�~�Ì*MRcO-�f̠�(�Y2�6�@�4�M��I�}�*�����rb����V���
{�G��ϲi��_̜�xw��8�D�w�ͤ�y;�۰�P��`~k+1�{���)+yE�O�uI�j�n���8����
���Fo�>2��ͦkZ��G�P � }��N���o��g̞gr�k�f�;���`f2T�9�4��S�ى��q��|w��!Xm�LgyE�$i=��E6��TP?g��&��BϺiwg��]d�:ǁ�T�:���l��<�a�����f�d��1�N����Xz��m���)�C��d���I7���_Y116w���!���g����Oq��nV}]u���Dyԏ	��ע�>B�6fd���=J�1���>q��� �@�y�6ý�Ă�-�����Ϭ1N��QO�si?!Y:��:�����l*���ם韕�O��`�8+Ѻ�P`��2�j<o��`:��hͧΓZ]:��rb��Kp���:jW�U�\�ܲ���'F����`��j��E1/1q�����mm��]�������'P�F�LS��'V�O ��Tj���N�d,�:���R��0}��Jj&L�6Jg:^c���Z��WX�[7�F�e�fX�ّ�o���6�!�݁�k�7��T�-9Z�3h�����nGA�l8uW\�c����ϑ�h�ou,݇*�X�%�q��v�"�t��]�!q|��]h^�e
(<vf���0,;FYlI�ʑT$�;QKw���	]hټ�k��*�&�SV
*�S���f���K�X�� ��%t���PI�_-�N���A�ή���@<Z��i5G�iZo*���X���HZT������Z�ёi��::K��'[���Y��MS�M�;M���Q��[]�{��J"�k�Џ�VIx�f�]+-!��^L��&���~��7�[ͮa9�HST���9X��V0��w@'D;�����i}IM��u���b�i=���u��o,e�hQܧ�W*Z0��Su��}Cwl8�$����Vj�Vj;���* ��\%�1��ǜ�@M�|t����z�]�\��V�ЖVa�i������:O6�;�JgJ�܅�;un=	j�a�ak�Mu�����G�^��w�ʕ�E]�*���4�m"�����38�J�*ޓ�n�ԌF��5y���ggp��݊��4�#����ʍ����>��uj��f��^�\�qأĽ�t�v��򠙥R܇Fؔ�s5�����tD���۠Gg&���3f�ǩ�1P%v�89������}.+�����!�.��Ruh���D��b���`�
��rg� t�lkؖ�ܮk Q�hꗍb�������]�J��)��vRp\JՀ�ry%[�7��6�r��q�0n�N<7�7)�͛��1�en�[�h�y��"��7�X��+�:�#O48�fǓ�̷���{�����y���cLmZ��w�he�b�p4s��c������C�dz�1�X�BI�э���w'x�4��z�o���f�1�*�^I^vB�9E2e���ÞmΞ���/���$$s�#�x�3����6<�pg��y����y�o;Ȋ�/%�	�U0���3NU�wf���eAX�9�i�"M�l8��`x�3{�*h��[�IWk�3nܣY�>]�[7�kVP��	GR뺓.it��5s�Ϩ�a�f��ׯmWW6wh�&9��������A;(����t��_[�u	���R�3V�Z\`�sd�����lC�ci�e�2o�ry+��EU6]He�h��ن�,�'ƴZr+L_;.�$s	�^p���b󶓫:���8pDv*DmG�!�0Mh���Z����w>��}��w[(��բ�j
R��V6�QJ�4��\���QP����Zʂ�E��Y�JR�F�bb���m�Ym�JYQJ��:qL-���m��[iQiZ�YmP���fTin���J����bҖ�Z+m��,��)TV�+EV���ڵ�JV(�hڂ�����R��4��U(��c-ڊ�R��U��U��9R֥l���h�-���DT���h���Q�0�e��mX��`�̔mR���h�b��Kc)R����Z�m�j�,eıb�UZ��[m[T(��QEF�+B�MSFKB����T1��[(�b��F�E-[V�*���fZQ��--QU-�+
�+j��j�-��KQ�F���降V��*!lSN �E-�b�-E��jեQ�����[JT��J�E��[V��AkQ�b	[l�mm&Y����m��(�iF�cj[X�R�F�R�"��9�c��p��v�3=������[���#�o����4N5�!�`_R|�^u
(�80�&��5pw�=�+qK̥w�n�l�w�{���m�����[���f}O�}�h
)X}�I�'�=����5HTެ��O�Oy�g���'��
AO=�h�qYR�z��XqP�?K�`q���k�o�/λL��������iw�>���#��6Ϙx���C�}�G��1i�}��AB��n��d���)1ӤC�1��o9�}7f�~aY�M���ϙ*ny�&�R
z�����cc���^�mw���_xl DyEG�3���R���a��Ă��;��x��*)=�p4�0��CI�{������y��0�ACg{����l��ɪb,4§��y�����6©��d}����x�ެi\��V�<2<T;�p�x���O�iE�'S�� T��ܧwa�k��a�纇ڤ�
����i�$�ĚJ�{�1>d��s� �I���M���`s�۝*}v���~�\S1x~� T	�dD	^�Ɉ�q�>M��M$��d���5l�'ua�=�� �>��ʲb�u��|N T�}��m8�����0���Lg﹒i�2W����ߵ�y����k�;����(����5�$����٫��<T+1��8�Vk�4ϘTX���g�1:������Xu�"��V�P��9f��2b���`� �ٜ*&5m�Ϻ����k����&�܅���+1�y�� �����%UH)�)�:�k�r��1�}M0�
�_ǔ��h~B���16ì�:��p��}遛��oH������&ީ�G�La��?d?!�y�&!�(b,4¦r���ɴ�B��73�m
Ì*k�Rc��Y������{J�@�4����'�^R�~��;�O�&���r�����J���gjy{y��~f$�Ğ%�ti �Y>q�hc� �߻��x��XbO=��6���;ˤJʞ�邓I:�C|�f[?2{�'���AHa�u��K �3���<f3S��]J����㉤
óʡ��N9���i��+�'��i��+���d;���!���lI겠ny�5�Cܰҡ_7́�k+��`��|¢��RǶ<*�<�c��;9�zl_��n��]K,��7�T�4�zW�+��v����h��,��!</�W����眡��[��:�Ws,���	�i�5����F�X�	&J���r�G*�XutkS8m�.X{n�f`�2r�?�Y�y�=6�5(l���͠����W�� ��v���̿�@����
���d�
�P��a4��d�O-QCԕ�����&!Y�O3�{9�l:³��ֲ��ΰ�s'�U ��4ui��q�o�,5�B�������/�����ο�@q�c�`�H�i�Ɉx�E�Ձ�Xq���N����&�ŚN0��ۉ:�f�d��/�J�0����s�b��|�M�a�L���Y��Х���P��/�v�\}�( D��>^�Si�I�xk��?2�����a��=B��Y1�$�Ğv��ALd�}Ͱ^!R���M0�l1߾�iiY�g�s%@Qd�{��{��k��aϳU}p2@���&ݵ���6~d֬<��H,�߲:�*��aY=q:�Y�V~CI����va�
�d��i ��J��rN�AM;��������Ϸ�[ݮ�YG~|p��~�C�������A`q���ϐ�6¢����i6��14���'��C��,�*AN���SL��QCi+��>7f�z�gY7=�v<&<:<&=>9;N �:��{���+����Y�z�'UT��a����,돿s�7�B��y�3���*OfͰ�1!^��AM��bzw�)�H?�w,X�I�1�A�Tl1�s�Rb���|�����_�(��N���i?!X{���a�?��:��`_����H
/���m=@�>���d������l=a�Ri
��d��c�}�)��`]��}Z6�᝟}��;;���*</�+_h���1;� i+?;<�&�Y4o�4�E%I�u�|�l�'uO���6�Xo��wvu��y�kB��=q? _N�D�O�4��ʼ�"�9�j+�rN��_�}��Wvg�)R=a���Y>�)�/�	<VT7iԇrÏ��$���egP�|¢�Oh�g�1:����,:��OgXL�Ζ�⬓d-2��'�K�xɌ�sY"��+��xs�q
�a����a
Ì+��'�H,��d�O�*�J�O�8���Xq��!_���q6ì*�&3l>�P�H�Ս�2V���r�(��"zN��8��p`��'-0����y��7ۀ��S*�rk��7=����'0c�����4�U �=���a3á�A��|��:Ye����PK��Q���lx{#�� Wʬa!>9�-&������ע��}U_W�^Q{�8����R
q������&!����rb��1�r�m
����H,+��/�$�
�j��E��z�i�+�M�g*Au7�I��8 Lx�B�.�?�t��TK�D9d�����x����r� ��8���u
�S�w��>|`��d�{�]�x��]��36�P*T׼�Ri ���Y��)*O���L���:�����كҶ�t�������� xn��8�ז2zϐRz�Ǐ�|�O�?3s�$�6Ol?2x�kd�$��G9�q!P��1V�{����˯5�h����~��~o�����3�N�k)�q�&�s�m �a�~�iq�@�*��S����!�~I]�s�J��+:Ϧ����
��{��x��) .�*�>�����U=��}| �~��ߵ���6�@��=>�Qv�����aY�cXT٪2��1�	���a�ܚC��1!����f��1=@�:�f�O��d<H,6��0�d�*��'b�5Lw��[�w��,����a�P+:}��m�+��βT�cY?&'+�6���z����i�aܤן`i �k~��u
�S~�N�`�B��~�k(�����~��Y9�nH��N^^���~�\��S��w��IR7�`~eOIXnw�P�'���0��0|��
�[l�βVz�bz���<����!S�M��7�B��
���i�1/2�V��S��[�շ���C�{�:y�&�(��Nr� �!ܧ���⡴��g{��l��f���H)�cw�h�b�wf����gXV�
�����6�P�>�4����l_���74B�rrA��wU_�z�g}�I���+���i��`~?s4�Y*u���9�4��S����L����'�{�l<gɌ4���ͤx�e�%H)�k��f���AQ�N�l��(F�:�7㚢9�~��zc�<OXwE ���ojM�<�CI��1'��~��m���w��Xm��Sӝ�6ϙ*M�������&�<������,�e�;��x�2�/���8���M�V��h���Љ�^q�h���<�[�^̕ 'ug�]�n\e �(9vg@⹗;3���c�V�_�K�ڗ�͈���R��G��/���g��Rs�����@��'��)Z�\�\[!��b;,��V������NodJ�0�O�� ��?�y�ԟ%E!�������!S�P3��l�A�a�qRT7�d�eN"��g�����[gY��0;���w$3�za��?\mps�_٫+[���{�S�Lq4���&�|�M!�X��>C�y�k'��6e��O̞�<�&'�I�~fM$Ԇ���R
k�'2��c8�~�M��Sq��oL巘c~�=��꼴X� 1 �?k�Ì<E��Vz}̓H~I\O��`x���C\���~B��'���*M_�i�d�)<�g̕:���1H)����g]�<%�Wυf�IK�~6�c�<�c�|�&�<a�y��P�����P�����1����k�%b�O��{��%B���M (����Xi?{@ğzoL6��E�a��A�L}���t�
�վ�J��q�yǽ(m
��OS�:~�I<C�d�<�e��a��o��q�|���I�TY>�dS�O\`�C�f�A���������i�̱Lg�IP��>S�'K+z��;�F/�ǽQ遐"	^���d�-�s���Ì*O=����$��t���d���b���!S估�HV'��&ߙ=L`y���J�d�QO'3 S�
0�w�*tS?D�o����G�舏ds�}����R�����C���R
Vy���P����,:�gWL
��+���;�<@QC��hi��$�>3�Y�'��![ߵ�϶w��4>��q_%��~G�G�{Ƥ���d��?eUR
q�氨,��^SH�L�1�����Af�n_�����6fa�bN����&~�V,�q�|�� ��{����:^Ի�3;����eg*cc�s�T "Gß�6�i�����P�auE��l8¡�;ۦ�+:�S��Q2x��M�I*e�G���)
��s	� ��j��I:�~�w3j���r^����M.G����#`}��A���g��P�$xw���ꤩ<;�4�'�����g0�:�d�[tk�,����
���ć��2��(�Y<��6�@�4�L�{��>P���Y��Iw#���=m�JvTʎG9i�j��yf��͘Y�t.0��]k�tl���	���}�]�AnW�.�zn{�{\RPk;�PRo��WE��,Sb腓�OO{E�r³�umPw�銎�qR�YZK��j��G���� ����sq+��8������2m1�s�d�1��d�S���D�fw�ͤ�x̇��z�T������3���,4�AJ�9�§�:�$�j�n��
�� B����>�߹^�|f}0<=I^��?2b���&��@ě|=�L�'�܁���aXVi��M�9�i��S��;�j�:�r�&��x�0�5p�a�i1���HDz�Us��K���o�=��z t `�14��b'�c���X��<Ì6�R=�Y��b�<��L*w�}a�a��S��,+
�Y���6����M��mE��P&b�E�)�nOnw|o�\0@�!�����YHVO���'�T��̟�~q'�Qg����2u��3�T��~o��l1 ��bVqRVkϲE����S���I�
�ԪN����9o�wٕ��Q�2}��#>½�� i!m���a6����Qt��R~C�k
��5�>5g�2x���Ն3�J���� ����	�eH>ٿl�݇
�����ֹ~�0t.����ӏ3x�ǀQ1�t�u����f��'�~C���>X~a��N���
����S�L@QM��
M;t��l�?!�~d�9�zn�0�³l��wz ��J����69�U[��/�U����� �ǆ'Y����߰�ԅa�:���!��Y����6��TRw�16��bO��� �d�]�<a���{Ef��bLJ�aS}�y���'��7��uV�|�y��}�@�¡���4�Y�<?Y���M��� T��ܧ��!�o��`�rj��*﹆��O�I���w�!���f��/��O�h�wz���;���k�{��
m��Xc�� i+<T�ެ��'̩�<��������ճ��Շ��� �>���bɤ�6s�|N T�{�4�d���3"�xLl{�G���S;5S5i쿯��vO�J��{�����l�D�+*A���XmP��Փk+4o�g�*,�\M3��C�c��<��E7����AC�6{̛z�Ɉ
�|�������uy��}�'�����S`|�t��F����	f}�$�C3��~lo�pn��q�����\x_r[Ѽ΍� �v�ո���)��^x�)(�;Z�^��1Yg�¿���H�g[���_"�L1�~�z�<K����&�6��^y3~rmY��z������ ���<q5��� (�����`u��&��L̅a�
�CG���Y�M�XT�U ��dS�u���!Xc?}��u�H/��&���E���16ì�>���ς@��γ��S���> xFϽ0;繦|������7�&!����,6¦r�ù�i:�a�^�h�VaS�QI��gf�4���ɠ��S�&�ܿkR~e�!Y�
���+>�S��11��G�0=��ğ8��o�4�S�'\|�p4��H<����x�0�V��y���f+���Jʚ��I��B���,�g�Oua��ݚH)�����s�������{����ٶJ���/rN8�@�6{T1=d띠y�4������7p��̕�g,;�)>C�w�z��<��!�XiP����4��eu;�6ϘTRk>���߼��s���w3�r�`Lz� lq�m��15�d�
�Pѿp�z�d�EQCԕǈ�~�D�+:��wy�l:³��ֲ��ΰ��a������掠m? �N3�.h���/�j��I���]�Q�}YV��;Wf�~aP6e1�a�b!Q|��J��1o�q�Y6y��6�a�Z��Vk�LO��	Qa�;�<�r$�+�;f�E���￾��c���\�������{�>�zb��L{�z�@QqO�ȦӨ'��`������|&�m�ۤ�
�5d�x��y�b)1���6�x�H:��ɴ������HJ�+/7��]:���{��qu���L "G�pɁȤ�4�NϾ�|��?2kV��H,��~���d�
h�5��z�u��Y�'�O�v��va�
�d�=��z�_;d���O��o~w�������8$���:���)r��g��3i�ֻ��g�i�0���{��m��bi�w�<H>�b�QeaR
y��)4�M2c��Cĕ��Mٴ��Y�M����f�sz�����޼��>���+�+<Փ�R=ga����*���'�:�θ�}���)
�yvΦ�z¤�~��a�bB��3I<a���h��i ��ܱb�&0�L�����8y�ٽC��t�T��y��2�WruZ�K����	����*��5�Y�y�:�Mp5:|���d�5���e�
K_5��:�jՠ��-4��jću�M���îF��v��|}�T�^Y��h�i=�!�~��w�����wڹ~���J+�t�c0��@�@�27�E��Tѿ�h���a����
��<�M!ԕ��~�S�M�(�Njé����s�h9��^P;�i��?e&��=̀��Lq��߳���鷛�����D�<"��.�/�VB���y��'��������Mv�N"���*}�g��/�#����22�!3��^���i:Y��9��M��Q&l@��c�Ѳ�k�bGx��=�Mt����b^�>s�
$�eu�n�ݣs��P�H�j�=���K�
.�8�v͇s���]w��"^���PH�jdst�uW���(4c�E�BtGU�Ϫ�x�Ό�	�nw:3}��P�.��Z��Ȅ��\{����n��<RDE^�p������GTQ�gw���j�j�^�j���^�°g����O�;���R�"�3����Jo]:6�Nc����&2nH�&�a�Q�'!����UҎ�i��v6od4U����v�n�O ��7��c�Ք�A�@�z$4�"4�k�Ǘ�lG�ݽ>t����xl~e�������Ն���5�WG����PvSC�MT]���ʸz�A��5��/b��ң7.���VX�[|&"-'�
�d��qC��W�y�����V�GrJ�g����̔@$�X���+e�*�{w�V�|=��o�G,F�Wv���}dɀ�s��3D�k�*�����6{���`�{v�[�L�����]N����}�W���m�;y��J��H��,G���bj+"(���	���eʰj��\TV���t�)z��Tj�V�S�} �T�`�D�)�A�h�M_�G�Z12*��!���u����e�zDnfj�h�O���X�\E����q�J���z7�Vd\��=K�e�齩x<�ŭ����S0`V1^�%׌�s�6�p��=>��N:��r#'M�6kqH�&[���3�����V�*&Y�	T���{Ɨ�.�N����w��*�����_,�3�������VJ��,�u;=�CL��4E�����*�_�V=��c`��#�g}���% �α��������WPgc<з�-N�GG�`ͭV��3l�S���=i+s�JV��\yE��K
��OXn�C�����=��`�v�}F97����d~��2���T2���c.�>ƈ����#�B�)��$6�&/�)5��\��� ?	�� �R�"�ڋ��Dmy�B�:���g�m�p�+��+9/�Nf|H����o
�:��t�9n1��}~���%tǕ���w�k�_=�nK��G-d�;fMb�i�7�����Kף`��:K)����c\c�)�86n��)���*�n�ң8��U�0#����!�ڻ.,.絥�*� �շ�Ʌ��^%�x*����֔ry��@����0L�C�uz(�jldې���7i߸��,��U�o|�"�՜��	�%:ؚ��n��T�v|�&G�\�*�}��xb����v�ե��BV����}i�6!91@���>l�8 }�����T��A墜��+سl<#��p���,��l�J����8"�t2$*LD��D�����<"6����)ͧ�0�������:����_�)�P8K@�aΜ`5[2[�J�6��O�U���{��rDi�*Єs��Rs)ܫB"���L2���\Ն���[�Q��eo|��k5P��e��L��x�]I��Ʈ�C�9��!�P�u秢�\t��G6n��Ř��n^v�>�
"�i�{��0�WH�.T6Kr/�0�P���9)��|b"�oS���%E��)e[1��}+�S#=�iC)b�b6<������Y�!�)W;�vh����%:!�FFD#����t��$W�Ey�>/E���{��ה�O&��~b��Z霯aҿ)%��;��qPnrE�˥��M^�_XV��K)�����Y��!�,Ք���{�=�EϤ㲋}I��oQʉ�A3/�d���}�|�!ih�ٛ(�F���2�������+מ��M�n.]���� ��k֛��X�FG������t�Z�\��@��ٮ�3rv]]���t��H���1|��0�&��±����j1�?/�oU����(T��ZH�1 v��c��U����*�A����*GC����	�Ρ�^�+�4T$�[.�]KLIܼ��U��
���[ܧ� ,��9A��'碝B�����N��V!�+�q��ԓ�#��%̆�ũ�3�/�tM@�� ��*Q&���k�u�Q��W�w3C.B���8#�lȷ�ju�%Xr\I���
WQ��/�Q���\ٷ�6���/�u�| ��9���Vx��۞�у�CG�ߩ�Bcr�7!���`����Eo�p:T��ޕ�}]sa�����{ή��r��Aq A�� ]��|���;\�V�x��y*n�r��2%nu�;��L���R��s[ fa����b/fwp���:s�+�MX��-�����D�~���ǂ��m�������vj��G�K��R��s��j�4s��m�N�ge�dWɜ�o+��-��a_4�`NX�W8^���err�	)Lf��k�x
�m��J(FoN��[aɗ�h��Y�z�U�j�īa��γKTD\�~L���pX�F����u�u�FS��b16�����{�@S���%���=4ҿ����;����E)3@�ݜ7;(t�x��	�cr�yk}�KՖBX�|�6��VrK�p��k.�9�,B\�(=�_u�݉�o.�4�e���M���C9a����)�B��B��(M���Z�ӿ"��^� A<��.�ڃ�_"� 0k��M��f]����7�D�N�|C�� �(	ӷs��՗��о���(ǣX��ɢ�E]����Cm�����ʗfSqm�|�v15[!�P��H�n������Ľ�R��h=Pb�\�1��]}** ��qR�i�D`���<璇;Tu.j��ZhN�Zs�,$�Ė��vu:hV`�ھ���Y�sB;���/&ı�PFU�p��Ab4n���>�
�����v �znű����o�H��*��WC��ٗ���R{�ͻ��	b�D
�A�V�FrU�H��;ʑ�}���<`��˼���V�I.�[:�9Ȍ<�u�VJ�(GPRY��Q���0G�-��z]Kyn�/k�V�K�d�E�e^��3�mB�E���~A&�?l#{#Fm5���I'�����W���ju�z��[T�o�l���B.���
L���:;�B����U-뉶6$�\ƨ.�b�)����oq��hΧ�i_8��u�Y�*����ȶ��ǈL7��#���H��(��B���y<+Y���O�5$�F�����\X�V��I���M/^��{�Ő���A�=��4s��P�xx �uo̟}$ђs�;���v"]̋]��u�G4\)˛�i�K�7 dy��u������f�D���؏�#Lb����wVmI�Z��u�4��9k��!��ܠ{z��8�+�p�a����fǦ�0C�,���Fe;ov�\��$
������s]y�^�{����cAq&�`K��j��+Uh��C��r����*+�\{B�k��])��S,}����ɪ=NVgcYll�K]�y��	��.��MH�7χ1;:�J���V�F_Y�}u�(��Xu�r��m^�/��=w�a����6��K�b��N7�qh�o�m^��@�ѭxrv�"c��������ao�g�z�ctK���/9�Z\!�^^s��<g���C��3Ѿ�j֣r�������5�i,�l�T��ۚ����tft����2��[��w��A@eؕ�) ��b
�e�x�f]cj��W��H�û��0���h��h�z�]-a�yj�+o[>�@�s	�A� I8s�ڍh�Yl��d��-�FՔ�E�R�V�Z4�j����*.J�b�������ե�u�)��i���Q�KT��Ŵ�[D�Q�QR�q,�T+q3kR�ʕj��V��ږ4aQ��D��,�V��hk)���m�"��E�Z#*��UKj��V�F��R���h�(��QQ�-�U��J���e+J��T��h�d�Qr���T�l�%J�V��TF"�(�K�]j�\��嶔U�R�[M9�T�%b5*�VңJ�̰�Ȣ�V�V�PDn��mj�mX��U���(��*�b��[DF�R�RZ��cj�Q��#b�ե�+D��[a[ThV��DZ�B���Vk\���[L*�,��(�klT�*�kUd����QZ�J�,AE4���mmKe`���XVQ���
�Q�Z
���`���F#QV*Q�i�QPPcܵr�*Ҫ(�(�h�"�VL��R�[�l]a���h�uuuk�v��Q�K$��YL��9��bc=��P�w�!�/�������N��^=�B͔ h�|�_F�Ҹ�Y� =�x;8�2�νS8#�zf2 ��u��'˩����C�O/���
#	ni�E�s�k�;m�(�W���p��s��!�1�V�z@|*`SU.,V���>�#!{�	O�r
�B�8Wf�)�Kx��chp��},%A���0tvhߚ��Y�@������\8�F�@<g��E�b�>�:Z���q�˫��&T[V�c�95H39�����5`L�|�![����*vUzb�3�c1`m8pw8�Z.�N�����w�3ޡ��#3�ZDַ�
Ű�̾�^Ep# �Snj&\רHF�WD7V9���L���4gD���uMv�C��7��J��D��y!�ᆝ�Vx��>C�EK+O�j�)��`�7��S4�/|P�}7]��nѼ��V�K�T(�E�����	���D��ݽd�v��*3�:��	�����db�29��:��W�}1Ң�����/eףx@ܙܼ�O��\�2��)?[= ����&Jo�?G�1�n��<Rz&���.�U:ŕf9ʓ��wam;4�^�jLRxW׹Q��,�7k������	��:q�������;:���x�8��*Fr�d��9�j��Zy�f�w�Dkj5�Κ{.�T>ܝ�/o��xd�Z<��M�K�+��N�H5���l^]���߽�� r�Jg�ؙ���
�L`��PnC�V��r�����}��2��u�k�hQ5�!)�M�X3'�F�`�4��yS�5�jڱ��kV)GC"�^G63���R�r��O�K��Ц�{�:���������#L��1|��� Q�k�zu��\3��7n^����G��0t:'�[��爈�xR��a�>Nݎ��*���c������H��4Ӟ���b���6ʂ���|ꇰ��`
��<"�xQ�G���=|�j�^qI�T07{~W,FF�T�`�D�>M��-ɨQ�j�d�!�nu�m��,���M��v�ɨ��`g#8Ӄ�E��9=�T�/��O
�����h
�� ���Z{��8��}��"��)T�8��s
�#�����&z�$�=B����Nj�7�q%�`��-���xG@���
&2�79Y� d8B7'aD4�S��08�>)iQ)ܧk7�FՖ��f�<ޥ�{��SZ��خp����%�^�,���<j0ޮ���y��v
���/���f�0��#R����㦸���2N�P����[L��7V���9�[�9b°�ƬI���eZ.�����q* %d˛C{���J��s)n��'Y��sL�
�C���N1r>��Øy�yw���:�}�W�<嶫���Ԯ:o�f�~d7 �Ε����-�l�tA��Tx"����0^�V���$��_k�s�q_�,#��H�,�j�<�q��:qN*��=a��#�>>T+�S��t�(�J�,嶵��^�!����~ʮ��ܫڵ=
")��V2�`XGd�aM�j�n#�4��˟=H�#}Bka�Bp@�3���Q[V�*F��>�5
�����bk⽚��퇴k{���)���#�+Dq�؇'ԫ�@�nr
������;�7��0�w�MJ���7��!7�!Bo&�o��/�_Wq���G��DXS�7�%ι�G7t�6F	�{�$so5t�=VTk�������Brb�|��S���44�k�}u�һI�rY缍I�Ǒ�aJ����!�Du���������dH2���JTe	-��xxz^��N0��&�����o�o��U�UL;�N��D�v���芛��<ɥw�j�V[ĭI��@��Ƚ5��@XC�~_;O���J�B"���b����?zE��C�͊LC�c[��O�/N埴�,T����t���%q+�ykL���>9 �1���;ξ��3cf^��u�U퉠�Ss��u8Ǧ��ٰz�E����������%7yk��7�pD�yKZ�E��[ut�d�w������Co�;yӈ�v�U?Ժ�� �~(AW'4+�q�G6��	�ڻ��}��gڟL������u}Yu����WR}�
�-
�;H�)e�C­���!��'΀����%�F �R������
�,��D���P|Ɨ�:jmm��ga���z:���2�]�O���GثD6!o���J�p'U�r�}��/�!n��t>�gvojNj�z�l����x����q���*!=W�0>�ٮ�Ϻ+r�4������9�<9�Qa�#HM��cl���1
�W�>�j1�.�(��͜�%5 �P`u=[wl�X��X�ze􍁧�A�٨�R"=s]֪��FA��^dOxz�:����D/[Վ%97�ٖ���R�{��^�V�}[J"�( ͙�aX&T<7�O�d��}�(��qp�Q���G)�*[�v���tN!�-Q teJ��_�EՅ�}8�K��okJ��]	(��׍�Py���X��*l?*`�W�] 8.�@s�K�:s(,6�E�=�,�f�y�[��N���֌>��)V��uu�B{j�R��D���a�QMP趖%>��ANZ���5��Z�����o��.�d���Y��8^�N�ү��J���~ū��5�v�m��=�x{�R��ܽV��.+��8���)1�.)�ݖ���;�M�����>�h�D�H̠��֏]厉�Lс
\z�\�]����V�����hl�mSɡ%�N}����ܻ�/��. {�|)�0�F�iP�aѵ�����W��C��?	)R���Jy�U��K&����ν(� ���)��^��{ą�
��G���#t
�	pT؎�Pۉw8J�7ro1���91oׅ�1�15�4�)u<=w�	�*��/p�Y���Lϲ�9oz?{c���
�mײ_�ڞ(EA�|cj�9�����2\NNd�hڑ��ֳ�]	�NH357}��8E{:����pck� [tvhߚ��C>��z'j_t��B���y��\��lL^0NB9��c)�7�Q�eɄ�u�ڷ{s�d^�Aj����iǛF��j1g[�;8�*���%W�+����Ϣ��HF߆�sw8�Z.��v;�׋�K�ؖ��o(9��h�#�k�
������ mM��r�+5�.���Q��޺<��
�4m�ޛ#V���Y�kI���@ˊ<��]n�_L���{�p��J��[��Xޮ�FY�5"�v7ݳW��jj�~������;�-J�j���T2=�Z�m��q쩻��tf����bG:�Tq���re�����3QF>ɦ�C�� {���r��-�{������H�J�>*$͋��܌\��� ��\��	��J����B.��|f>�L�)�3A�݇��R�FD�7j%�
:(vPW�F=S;�P�n�^��Z���aB�,��z
���,�����ȷ6qȥ�O��0��Нܙ�Fs&Y� ��E��bg���Y߯��̟��;����|D�r��aI蘕8��Ƀ\�C'�'���yy�'3U��.&.6%!#c\�룹>���\���I�T��l+��$�'u�~��ٝF}�u�F��K�u%U�յc�7P��-߲����vD&��sxu�T|1*�|��\:��������)��}2�L:�9T����\]��ؓ:ouFtf�>���*�Ni�T�J��Qtp�,��_"+��-�l�GsyLU�VTy�T6uI���ڋ�e���lp0~�4k�l�}v=�9[1�1eؐ3!�TT%t$u�P|�o���X7��F��5"%�hS�}QsHJ�Tך����Iݡ��/ݰ��F�i�32�3K'7�Kɭ�cC3�Fn
葦�:�,1YCu�%]���k{/n�t|/F�X���o;2��M�Tġ�c�O�z��g��h��ƹ��w\@�q�c@�d�[m�Ѳfd��pSͼd�ppͻ�3X:�J/���ﾵ��2w{��1�w�}�B�����uc�l\y)�o'NE�6o��V����h�X]��no��l�.�>�J%�e<D��]�.U�>���7h�}����L�kL嚨O��m{�9:�/�x�o;%�]���vk���x�T4����=#�AM����^�o[z�u���Ռ�U��<�'�S����D���j��Yf��s����5��%p�T05�t���|]��C��X=�,��ς��8%{��;�Y�w=��;n�Lr޶��~���O}�R�u����ǜgM��W@���`��G�3&�d$���QX��O2[G���-=�i��Ih�'�C]����\�H����m��t8g5���ޚ��~��9e�U��n�芎Х�6:�����0��V6��N�]~��c��%JR�j�$��խ����u�t�S���#�V/PHN��[�U�Ź�*B��Cm���4�Vs��۽z��Y[�	�Qᰠ�w8�x����U�V:4���u ��{�;�X��{D����Lշ�n��n����c�t�l�814����엝��ٚ��.��R��l�xn�ǳ�z��u���:=����:�e�	b��r=�����00�E担e[^�-����]Ъ�vx� �����q8�tʞ���@*ʽ�~L�Ϭk'*lNLP%C`�8"=�(�Q�ѫ�1Q:Z�݅&�R�X���96\;��G\ߩ<���`��C"A���P�ڈ�5�{6�,i3�r��b@Rx���t���x��U0�m:
4(=s�Xi����0}U���)F❽險���]�H�5ābǸ��v�r̭�-�S1L�u�YE���;���ۚ��\��`ԑ�2.�����x��إ�I�
�\j��񕛎���˔���:\5w�����_Bo�E�i�{��Gt�H�,\�E�ܘ�V�c���.�ʽvn�}[z�h��28_�;áK(Ž�D'��F{Pҁ�o��8=֕����l#��i���T��G�#��qy[���͗ ����Il�O��F�E��b+&�mcMl�b�ꬔ���m�
/�e �^��8 ��Bz��`}W�]���F][�ob%�w�^\n	9,T��ꮊ��&���B�my25��~�~��^��ܚ�O�j��!�K�S�~8�O�ZEeot���A08��bX����]kɘVYtSy�t�@VG��G�r'UMզ/���/h�Y�DE"��`���D*f��%|��������%����7В�|��k�vuü���Ou�� I57�(���� =�:��֜�޵�P�Ä��5µ�b���"�;!]UR��`tB��T�*"��:��ԙ�{��ф��[+�tem_*Q/{�ʽ�5��Nʈ�e@ \Җ丑0e�,�Is%�_*ΐ�����Qnp:gj^L�D��:��H��R��,U@��6�1u�Ό�b6���ʁ`�S�������u<tKQN'@�!E!��������Ku˖���ĨPGOB���<�.{�ŗC�S��/ w�׵�o�sN&�;y3[i�7�j�0z���4�:>�=���7���WGZ�#������"*,���j�m*��osz�:hC�:��6
�fcfݒ#��r����ߣ���0�Zt���g�ն�3�{��Y}����P�yH�Լ�u=�xlQ��y�u9�F���;�Zwlj/X^��	Q];o�n`��B��\���ך�� vMuZ� �l��u���a����"�wkSkU��V�n��F�z(EC}Qiex��/m"){���,�������t-4��	yP�ԩ�f-}G����k��g��t��ϵ�ޒ�aY�D���,�+�_Su��{�X�8�Q����}x��]���|��e�ÕjT��ǽ�kۊ�0N,7�{e�6��v����힮�ڊ46Hٻ �����������Rb5��Q�j���:Ϩ�"�u[�1#0���V@nk&���Q��}w���� KҒ���I���b�l�������an�t�{}�W9����ᩅ���ř��sY���^�e��a
��ff� ����[=0���� ��>V�����+s}[���!&��25-{Ӌ��+	U�K�{iՆ+�1�c���P�z��t�g��[Kpp��G·u�ӥ�J�����=u�|��e�1��A��u
��7=����7�����鐥@`)�*ƠE�	�p�+�ԩ��;���_�����]c㘰�����ɛvjݻw��<����|�>
du�ȷ6�E,R}�)p��C:�����.Dk�ST�ǝ(�Ul7��z�%6:~�v>"a�fiXu����
�	�cy�vvr��������Ȇe\�(�et��r���G'�C�$MB�!j���}%��E܆S�"��2F?R����5"�H�~�����~�uҽ�_R
��Eh�i3מc�ɵ��}(20��L�7w�u��i�q<���)us�K]Vq<ᡭ��xb���X�p�S9�ꢞ��m��&"-C��azN^��p:|$H��Y�w��`PqG�oz���k45,��j;�+M7��o�c�I$��Z�e�q���}����� Z`��B��>�;ӷww�h�6hՄ�+���ֳa�D��� v]mL�Z���ַf�L1+��<BU����Pr�s4]�]zJ�.�z�w���\�6��G݉����"�l��}����L�[�ۥ`��I�tn�t�F#���Sa���ůp�W�f�iܻw9���&R��E}ZZ�M�Uj�(��'�lJYK��'�q�d���f�x���@�9�v�=�2��׳��c�$���ʀ�����Րɠs�j���_.i�eh�q��
Ԉf���BEyh���1�3C�
��s��`�m�+\T����f'��{���rmo&�i̷�G��_B�T��Z�[�+�4N	3�%�A��Xo�y�_&�ԡk,DV�`�Oo�)Qe�K�jB�&�b宬�hLK"{X���3Mv��t��R|V�����P��:�D٫S��%���h�Υ����oxwda����z\YN�pa��ˬ��<ҧ�mW���v��P#�ha��;��qYH(/i�Ѧ ��K'y�an����.F�(m.�H`�K��E�6�n�4n;�G-���VX�Ce�j�ũyv\wO�L�`���ʖZ��J�'ZT�efX���31/9��%4`�AOC'�t�ŀAOR8����Rŕ���n��{�>�1�r�Z��n�ӽ�Oi�^��J����jSN����#��f�8p�z^�^���7K�rBd+�z���=Ww�䮰]�}�>Z]��+V�u�P�7	��b�,mj�nVf���V� VԦ�A��t��ui�� ⌺"��ׂ2GN��Xzu�#;[\Qٱwt����Wm�{EQ� �5u����N�q�e;������i�v��n蓑�d��w���*��acי
A�'�g�ç�2�����N�Y7�^v�f��.��tj���k˻�'=X�Sh.{���d�Y����>xkd��S��jY�z��ńb���Yk�����
���	�=7E7��7��=��?6o;�S.М5ف��ۏWi�[���et��5�:�V4*�Jap�v4m� ]d���x��\��JM����m�l
�MΥVRC:����AE�ub�ʾo.*SBP�fi�F;p�ɍhiҝ?moVG��*@+i�H�U�M�-��&��%Y�Ȍ7�{��Tŀ7>+/�]&5��z��j��6w5C�+����op��IY����oM�;X��˭�&��.b��[=�%�u�}���'�0WM	�0f|r�Q�m����%�֨�jʑEF�P��U��U�S�eZ�4�Xі--U[eI�*�e����f��-���TTp�jIU2�F ��`�ֹ��s("�b!h[R�X�L��,�R�kZ%j �AlV�QDҲ,����*���k
�U�Tq�m�.R���)DQb"��h���(#+Qb]Y�C-ZZ��1�j��"���#4�Z+�f-U�V�Ue�J���E���J�F��j�+TUb[FѠ�"�[R�L�c�PYʵ����mun��F�"��DQb%(Ң������AER�ET+QQ�����L�Q��6�Y������Ke�ؗ4�J����EUEuL�F(#+Dr�UR(,b"�
�Ė"�ԭh��V7M1Zږ%�PV)iDE
�,�-�!Qm�eF��RPj���U�T`���:�Zy�8/���iV﹮k�z����=�E��uX�vn�΁�x)Ygp���kO.Z�JѪ]�3^�(}_}U�V�<��-�r10xU��x7�C!�G�J�	���4�9�#����ǖx����d;����˜���Q�ONAO֯��T;>�J���D���0�*��+ϋSF����;�E&lL�·�C�/�h�3�j[�'j.��X�{6 �����<#X<3ֳ 6mJ�w�x}�ۣ�Pm��C*�Δ�ؽ<�Eu0���4���c&�J�T�����C�ϯN��Z����7c �'��pJ�G�����7�N�G��l�4�!-ַ�G�OQ�������n��ߚjO�rWB��]��nsFф ��-�w44t���ks�qe\?��o9��Bs�AV���4R&��-�Ⱥ� Y53if�,+�+_;w���F�w;�+y�a;##cPٚ6��6��b%Mj�j#b��z�7�(�<7�7N�V����sj:_mz�y܃�{+�Յ�^��]���<��;�5)85����Pl�VuTtT;�lPT,)K>֬cd�� �:qJ�����"¾G[/��0���NCWx��i�J�շ�G��мU.ܮ͒6�K�7&f�7E7��2�G]P��1��\s���5i�������xʉ'�Vz�KѮ�Vf>����*��|����rX�X}�s��4pl�[�W��ϔ���|��t<q��.�=�� �˷[̧��+}�'ns�4c�V�9��P}r�{V��DE9э+	�9V^T^���V��	H��s'͎z�VM���Z�=Ӆ�X;q}�9Վ�<�z�kF�\;�f�\�\��2�*G)���V��ꭈriW��{؎	�/�el�>H�Ql5�x�J�(Ś}�s;2�\u�A��U�uN$�x%06L,4zH���y-�l�
�{��0V#J%Js�; �Ga�	����Y9S~���QQ-��p\�r3^ue�]ފ���~*�]��)6\;���:��'�э����D��q13�c�̚�&�$q��7��	�@G+���#iVt�3-:
��W�kE_-�o�Y4i/%��m�9ˋ$���)|���f�$���������|2<����׽�}F6š����N�S�s�]p���`Ԑ�d]�����f�)9�ꇃ�N���˽�OSa⟄Ny���v�Զ��O�+���K�u�C�R�Gt਌�
����<{���Otv�0G�^WA�NkT,��!��]lc]�j�� �#���Wv�A��(Z�r�@:�.+�]��J��@^n�A%X#����q��ڂr���o��v_EY�תL�o�[�R/��ʟ;��|tU��Yz�e��q��^�&�����x =�j��i�J[ĥ&?z*8Ef��b�Ga��,��Z>�¦7<��;�Z���w��w��^���ɳ�h�� f:b6.�D;�ǋ�6w�E�/Đٌ�@��8���L�[�����Y]r�v(�GB�@a�A�ݮ��A{@��_@�>�ٮqZù�wQ����ޣ~�?h�Vʏ��0�i	�ކ:\����B�my25ڌs��qt26q�[2$��9��S��s�{&mז<�^ʗM�:{f,L]+Ø:�[���h���5�j��	�/xv��O��%���a�DV�������_m
���(:X�E�P��"�R���՚�B�\mJR�ͩP������(�.]eKBf:&���UD����<DA7��H%֖�dK�����Z=̗:���Q�vg����T�"�_).$ˈ���4�Ns��;��I}�G���p{��C�X�m7����@��N�eKz�]��}�^l��{�z�|�Qk�4�*6�|ǰ�wF�}>գg+��d
y~�ޱ���q&L��UZ��kW.��6�h>���VŲ�z^�Ra�W�foܬ�/�fD�l�uI�g�籑c.q;z��L�{��L��<���#: ]�jΘ��;5�f_>�B�L��ׅ�]�pX`�ٷА��'!D�e]�k�+5�� 72�Md���t�ݕ�4"��f!��S�L��z|�+�x0ͯx�X=�𽰁D�����\�r�x���=���0�L該�8�)�lT���b��������4g=^%y�1�	��}� Ljm��N��f#��W������G�)�͔��ʦ9tkl�M:���G@���:7��1r�μ�B*���O�^�DR�r|t��Wn�%s�G�M���#���+�_,�]AUgU�a*�p�]Y���:Ռ�ܝ+�9U�����qL��ߨ�׹�Y���م�Ō-���1�up�����}�<̕z�pY8�j��L�d�?-�s)����f�]dZ����xi���nb�!��w*�xn_�ݺ��idnr;�9�Fo�$l�!>�Ԫ���1�����뫿mq��[�l��%�j���A[�Sf˙���6�ꕏ��3b�i�\���#��GG:ɐTY�5]��ɦg��v���R�X"�d8su�})U��ʉ�k��������%0��(o��2X/�K��S���/ՙ��h`ĵ-�,u_,Tj��c�ow�k,��^�E�#�Htb:�b����~�;�1��Ǽ�:��/3d�n�<�	��GL�;i�v�~6�f
�ng���{�oz�y�]vV�C��3���J9����(��3��{�3�����l���)u ^2�Gpl�sn��R�}F�@��ϟI��b�SU�xyQ��,�U(��J4~�z]_��%7�q���`���M�;}���iS�G����N�D
��gҊ��.v\��	�]ٳ+:�y9��<�m�[�r�( ��̑�Ԡ�&:r��-�8=AFT�70<�J��7�g{�I���V�d���h�UZt��i��k��S��
A����tqq���b9̞�����P�\C��:ʘ^4
�6T_���Ft,��ɝs��rz��-���e2(�#F�q�3R�'j.]1�f���"���1]R�N�gԭ����u˩1����#�#vY��3"\��./�ь��(�19Y�U��a����ۀ�ov�paѿ�)�	�<�S������ܿl`s�\�����JrĢ��7�V�u#�zZ�;S�
�a������^&:��
-n��C�T�Լ���DD!�pWf-v\��'Syq�A��"����icte�U�*��.��[�qbUl<��D�:�Qk()Ss��'pf��_p�����1o����َ�qٛJ��8�o��Pq���#���.�P�����u�?����cM��y����c�G����M�g4��{����h�*�&��	H�,{���Rf�� �#�%]yg����n�߂��	�dd�YЫ�]Pj�𮮹N�V�u��3�W'To��߮ha��2��+��K�!�:α��ޏ�k�oF!�����D{$�>�<Y�&�'&�i��A��lg��Y"���X����Yx&9�P�k�`z��.v#���a��4���+�VF0����A��NU�Z��*"��+
�1�[�k';��ku���6�kSC�Hl#��K�luKW �{�	V�`�X������.z����t.�����G:�{g�S������y
�3�eO�A�ܡ��b�GJ���|ѓ�vʐ��]�>Hs;2�K���>��Ҭ�ğmx*Uf�Y����Gd�Y�U��%-u�[��:pIS�p\��{�=���NTߡ91@�TIl��{!��{�R=g/�r��C�R����r,N;���:��'�с�:"��7�f�]yb�ܬ��/��2Q�@:��j�m�����������ZE���w�c7��]�� �9�ʐ�ͷ�(E��^��c��J��f���.�-I�iz]�K��Y45.�*y]�&9X�E�"������:���	��S�8�P ���8G�_}_Zn�&/]�TlLG�#mŊ.�:A¢��ӎ��UcUL;�N��e�C�0�F��-Z�^u�R�CQ芛(W��t��]) ,W�~VW���@/ygRc<�����,_�s�Y�P=U�jڅOs!����P��� �~:͊_I�<��/<U+��ј�٫�d�\2}y����@y{6 ���&��E�¦	hsc�=Ӱ&OKt+eG:.�q��v�(Œ�L\Tp��u_�;ȕtcC�"b�h�+��3_騂]�uT{�.�)R�a�W����s�� a�P�"�TC���x��^l�r/dS�1;�-�ɑ�S������>cۂ�.���Q��{ҸKj���x����N7����OU�k�ŕ˛��Fcjj��5o���+�06*�l
�Qn�=�����b�kɟk���X6ՌXr�Jɼo5�Z3���Y��WM@^k�HB��ȃ�7��1�,
��\�A����>�ӑ�n+�+��L��� ü�!�n2V��L�FV��@x��^��c�R��{|6�A��Ov��������(u�����]����YY{{AC��z�3Kn]��U4rψ銑B�Ǉ��`�R��4ؘO.spEo��ٔ���ҷn`�r ������ռ�Mx��V�o+��+�w\�U�V&ݴ�Ƥ[����zY���g���:�`��B�n*s#�t�ܹu�-	���XV*� �/;*7e�v�*�f��_�R�>�{�^[=�d�מ�vu�=1�ʛn��v��3��6��|��{v���=@P��V�3U�B\8#�aFZ�\�K�.�t�N��^��]t�ml�*�O"�r^�DW�z����+��Q뇲�����z퉤e;�ŉ��'('d ue��'����o��ЊJ�!�]zf0�J��iUP�a�^�>��EM(����)sgN檈�~�=2���h�4Ί��B�I� yL�l�	�sX�V���ƷS�9�XFX�*́����'\!�3s|�W��@���É��SB��1{�[���
̳���zh�%���_�G��P|�ګ�sP)�E8e)����o*�mfo3'u���~�ӭc=��|L��x�J�-OU�2<Z�W�U���߆�:fY̽�����>��,�X�F�=�7p��*6,an�`�1�up��N�/�sn�ޛA@Y���C��AS�[2�-j��{C��B�6��kQ�Y5m
۳��'P�`�۴��Y��;o��4��G:#{�iT���dA%,�#h��m�zrc�[��c+V如PVY8)®��\��z0Tq�Z�í��a��}_A~�ó�M��)�C�V�K�պ�U��%(�N�o�-���HF�M�F�N����5ۼ֪�S<�^��+��U������5��i|��̗8Q�`d׶��.��E��FlΖ�[�V��B9�S�n��7�eŇT;'cG�S�Q+�b�o*�>��Dj
ʓϖ���GWv��sY�GK�~٥/X�Zd(Su�},*��=mډ/P��Dݸΰ���dfn`r�/es:�n�*�P����uGG��{��{M
vʙ����E.�]f��omNN�nBo+s�����qt'Dq�V��R�P<ʋ��������ɂ�?G�&�� �� ��������e���g��sg|~���9��Xg�C����J׳�Д�M[��B^H�d�q*6_�TXw�:�T�H��9��Ԡ�&:r�Et�l��AEp��Z|��]�ĭ�ъ;e܍��ԣ��O/#��{T2T{iR���s1�jQ�R��5�-��s�0��o�l�n�b'}c�A�ub�r�U�i�T���@J��Q�ֺ���� �y/�;(c�3���ɫ݄�I��U�r��.�k^>�]'>�7j��`O�{j<�6�x�)�(ݞ��Z�u�7=��=�M��nn�$2]���{�����t	*<ω���M���f��un��=f�]�v�ЃR?ꯪ�G#���#����v�M�E����6��3�L��Pe��a���(������h�'>�}y���<�X�E[=5ߗ2�Δ��N��%B\�M�TVI�S��:vv���^v!^�c�Vl�~�u�D\��dP�G#���[��[з��fR��d���t�^X��+���g�Dkh|g��"E�]t�'?�>�/�\v�{<��^���*�A�S,���C�$߱��0m��%�8��d�K?n��/=���C0LV�f��FOG>��qy�263Ϩl�gb�`�u��]W���	�ݪ��RًýY!��}sCc����0�/v�a܂�:����Wc��q��&w��Pgz�d�,�%MZ��0}s��A�$R�u��ݸ��<'�?1c��{ޚaˬr��)�ީ��g�BQ8=��Z\ ����㲏 �n�<�*]��6S��>S3�ON�X��vHV����=Bx@��� ��Qڵ�46���s�j�0h�fk2�ꦻ��e�QH�6��I��U��X�Ӹ�<`	�sd���i�����[Ҧ��u�]�D�)c�:=�bCz�0��ͽ�$z���Wj��X�-Ũ����ڕ��f��լV����M`�A�]u�fm��p�i*��!�{�z��V��H��t�0�Cm���-,��/��R*O!�Z-�puζ��w�M��  `J*;J9�D���Or;L��Ky�(v�lHە�pvU�h�U���)u�;��1(�X���7rE��ރ'#�̈́�˔Oj|�ja�gGZjQ��Fh�k�_X�����1��1��=�M�����fE�t�u}]��M��r���6�T2ӥ�V�r'����P�dt�2ޅΚ�14�����ސdj���2���7:Ԛ������<]ok\���{U�U�q������3u�hd��s��`6@F�!�Y(V�}_vB�lP�LMo*[��n-�	�:�8umM��vpc���{�6���-��W|���k����K䅙|FkL,�z���U��32�(�4�tR��I�BvX`�C�=o�DWS��|��<Y���,z��s0��E��u �k����.k�0`�ıVZJe���ȆU�;%G{W�{��w7�V�
Vy�Ȧ,��%�<.4��Ī�7�Y}�:�S�]i�u�r�ԉ<n�lZ�a�W:?z����rݍ�Q<5ڭ�Q��#q;��#/Eњ�ӹj�.z��WV���FMȊ�0^��,%�R�A1b�8]�\�"d��;L�Řm��[�frȦ���am��{MLY{�V,ٛW��RfEj���<�9��@U*�ˎvC�#�	�s�:��vح���ԝ���.n���I���3��ה��b�><�z���ݸ�2��㕄�s��!C%��4ڠ�v^�f����Y��ab��j�	E��QH$��� *ܛO�С G�al���Ʊp��R«�&JΝh����b��^mw\U +h�
���n�LT���T
��GL Wz��h�{:��tB�S�&��Yr�$Tї�(N�of-{h�������1�m�N�TNn驗}r�+��R@Z2Q��e��n΁�W:�V�g%�h�s���l��a���Q��aX��D��(��Z��@�z�eb
�<{�Ģԯi�6�>�QrQ��5�s�ή�ƇP'�ś��<���>'ݺ.YF�l���;<#�U�;�'n��C�K�Y��>0An�o����(uθ
�i+�\.�3��j����}�����s����Y45���tC�n�`��ޭ���������}�G�Y�=G�9�SX�l;��(��݉k�ۙtベ˺Q�,(��Ÿ�R&K��$РT|:����Sw���(<�*�����+W��.��C�!GR��m�c7y�-)WX�f� Hxev������>.!\��GE
�*�;]�z�����,�h�P |�-��"�+fe��EC)*",Tj��.e`��imI���U��֥UT\ITAX�Z"�J������j�,E���J�ZUE̸QEc-�F#�"9h*��6j�b�*�U1EA�4��UX�!F��"�#*T-uJ��Pm�T���1��M%E4��4��,ET���1QUTEPQA��iF1EU�"!YX�QPTTTAX�[l�XŊ��]8�Qb��UU&�f
��,QB�U�֢"�T�
�QS���F0QAb1T���EQUm(�����"��#$U���c`�#E",�����b��"�k`�ut�V ��AX�G-,AUb,F(�dF$b#��U2�X*�A����Ub�ZVڢղ�m(�Vڶ�c+A�PU����UQ�̪%aZ���D[b
��ҍ��QPEF
�����v���;t��PJS��bgLmށ��
g�sn�^�X/��[�N�׷���;Y�o���hL�~��72�\�y��=�?�8�nf:�m� �mH�#�P���
�j�!��z�.if���x�$j�QW7�t?Y瓿#��ʇf�m#t�<�I^	L��p$�숽T�J�ū�kS�W93�@����K�s�\���ɞ������Brb�(����R8(-���^��9��<>�y�C��Z�+�x��VS�vwd;(���I��cvtAu�|��j��C4g��6J�k���md�>TjB��p��7����Uꩇsa:
�͛p4Vm�%��#G\eX�93��OԾ
�P�T��]���;O��+�t�M d]R8�C㙫GwS�0HH��:�sVј5$�"�= �f��]��	�| J�x+)w������U�R٨��pT"�q�z�p5u%�Z��Ot� ��u�U׏�j7�Y,\�"��&,�b(gPpŤv���=4&+|>�¦6&�f�s�y��'��n�(��b�����Gه�r�yጡ.�D;�ǈ}���e��������>��Y[���Q����y�g���زm�.�7h�$z��׮gU���}���Pz�����ۖ2��g)v{n��M4�?��'�e|��;|s���b�j�rj=���.I��E�;w�`���q�m�Q㈪"��N��o�DF�7����]<�1X�O\O�a���(ԑ[[r��$[v^��r�n��R)���Hf���9�v��ĺ�y�X����*;��S�Bz7���peO{��ϧ�VP4� 15�8�{��!v簸�M�`��'@�"��.���(J�xs�V��F!B�|�J�Vwn�ʴ��J��0B��Mۅ�d���H�k�������_/��sX�
Zt�j���q>S�{:�!�E@ \Җ�6mH�&�w؋��Qnp:gj^	��C�WZ�z�"\�z��\z� bG4+�D�SR,���Ns�=>8��i��*�l>[��>������Ո'�ÃPՃ���n��>�i���u.��}��c�D�N�z�f����~�De��Fd����PF	�.���֩���'����r�r"`��~v� �T�hE%Sخ�%�H���Pb2[���$)�A�q�����J���(�5u)utT�C�4`L�"�������E�R�"�ڻC�<H��{��`�ŚΧMf���qn`��T��7��T��Nv���Y~�k��f����4�7�ƙ�a�{����r]5��҉2�m�����c��C��2��KY�������*��Y��YVz��P�;}��L�N������o�6�-�W�W�@��`�������w0S�!��u�CQ>��\]���~�&��L+�MC=�xi��F{��8��@�%���aQ�p���T�"`v�&NnKË^�ۗv�Hف꬈a�,��j�?��V	~����uW�x������b�b�Sg-˅g��������
~ܕe��{)b.���9�M��Q�eɄ�Ӂ�{�g���u�A�RA�1]q͵�3;φ���fnr
�O�+��z/�iۼ��h��}��CVH�8<*dYw�W}-{�}CG:h��$l�{��i��h��3����Ë_�D�i� ��y��B�tBuc�7ӧdm�B����_�2���A��R��"�i^��q�b���j�E�lZ�r�v�)v5�-�C���b�
�lOXn�LL<	�ށeųo}���V���[j�|�#;�P��SS�6�_P�<�u�E�62M����{Ժ���Z���>�l#Dv��s*=g�Q`~�z����	Lz��3�3##"�Y#s���;�`�4�ML�\~��fN��6�������f�t�Z����]��9I�Vv���ѩV�n���D���d:2Nb\�s� �]t霺���e��ҳ\���L���WBF�'�O+JJ]�@|suﾯ{������ly~v���*�sO Rz&5z|�`�3q޻˃�����ꖨ��B	����G�x\u��a�27֩@��d߾<:����--{Φh��)��]�s�Ѥ�(T��R�F�V)GC>����ٽ��<E*Q ���v*��8��C\|�a���}^�8a���Z��b)>̧�Z��P�\\�pE��-������@�8\�p����QӐ��)�|������h�
uI��;QwL�"͈�V�>������K����SA���z5ߗ�/�X66��#z��.]�흙͇v��Ӗ�M���8�MGG�q���KA׃X�����s�>�G�ϱ?yǍ��@{u8t�z��w���ty���+k�b�}5a�"�G���$T��P�qWh�s��D錶����%�x���0�n]'1ɞ����g6L��%�
��v��_Q7f�T�+�&�Z]�zN���bNh��v��5�)�Y��g �[̈́����l�[���������e�u
f�'��^J���OD�ә��m�]}���M�^q���!6����k���6:rzYWG8�6�fh�.�O�Yň��j#'SV�5�wi$��Ƹ6(*�n��.P�N��6�w_\�ZA��Q�}�[��z�&U��~�N��+p�;��\1���i�V� :α���خ�:v��sj����Ϸ�61o�[A�ݨ�O��~V�?`O�ϡg�R�u����ǰ\tn㜍��ӊ�Κ纊R�[�P'�=|U
�=m1tNx�֗+�z������ ND��3wp�x����S2�3���D��&r�]J �j�n"���E	�4��j��]h(O+�I��]bS��8�b���ԋ
G@����5��x�ֈ�+&�gW�g^d�z�4��mHQ~&�L�.gfT8�5i���x���:LsK��|�춅y�s)P8!W@9%ι�s�
��aߓ=����r��	Ɋ/�3����]W����z������6��g���]����ݐ�P�(Ry}�"6P���\wj��vj���"�C��b+Ԇڋ$\"$r�TX�eŁ�x��3��̮���V^�B-�*�P �t��5�#�Ծ�g��������|�>$R#Hꉄ�b�ݜ�Y]�z����ٗ�%zY�~�Qg�����M���0�l�/��e5\sp�d)�����{ޘN�X��;J��8�U���zi����j�M�EYK�ƾH��66ץꀻ��9�a`�u�,L�gټ�3���M�Ï�}_v��?7=]{�t��e��W��L��u�正0jHh2.�0z���s�r���#b��g:���V�b;U�FMF����7g��Oz�)����QWRC�S�99N�D�j�Gm�6!��Y�9�ړs�2ꛓa�A���v֘�^��^���]|�v�K�+x�Y�z�l�=�5V�۬ ��9��E�B��z.�D;�ǋ�6g�wS�Z�ydv��)�D$c'��REmm��[�v^�Aʱ�z-O{�>�[����"�����ϰm{��+�MhX����;h�z��'%Dm�*��@mk���K�=^�<t�>��+31�.,D�Vl��IM@�=��p�A웭�"�R-Q�6&�L�m&�9Kq���>��F=X�y��Z����^zf:2��J��<�U{�1�ti��ya�4�Y�b�đՔ�/���-�6��Q��Ndst���v�������}�0��F񞝙����j���
���.�}|Z�yh���Zd(C�l�E��;����>���{�w��ٰ��yiRU�s|V���YY������{r��C��5BA��v�r��+F�U��ٛ��\�Qv��u�2an�J�nT��3����K�ʍ�rL9���s;o´�e�|3�T��7���d�T��M[�$=�ܺ"��k��ķ����w�����Q?	QPCj!L��9
�<�.{��9�A5zqS�
�v��O2$;��gm��� w8]�g������Z����{*�N9k:��Q{�A�J��_3��ULu�0.B�+�[#j�M�R3C`�L�ͻ��\�0U��wR�y(flɝ��'}�u��/;`k>�\��C�4`gEM��N$�@�;9��ZI�u[��lZ3*2_��"��*O�K���t
��3�L��c�bj+�^h��Eg���z��\T�ޱ�QG��>�^� ���7�a�u��P[�Us\�k��eۺB�.��9/իR�nJ�����g�|2�Y�nXJ�$";�	xUԿY����|����N
9���,yUmL�ȥ��23
��v;���ӻ�k���ٷ��VB,L�h��=�&�T%��u�?"K0>��AS���0���&��kz�ʴ��^��;�|�{�+�Z9�Fo$l�!>���V#<rt�z5�6�u5M��=�m�!En1�^���o۝j�����[�=����&����+<�h���SK�[x.�>��]\�Ч��?-jR1�� \fNbvw�)�^�)�b���xv��mdޛ̕��Y�a���w�h9�7T'a׭7?WՃ�D��~��WWq>�W��W����7�eÙs��m�O�D�M���\n�e$���<Y���qT��i���Cǅ`<}��nӰ��Xz1J����TsgJ���b8�K����P젬яT��K�
.�5=�jU���r:��MC���Ee�F���Q�XU�"���n�KJ�P��Y�	��{��~�z=qO�Eq��m��u�~�ڞR⡭�3�w��+�L7N� ��L������"���띅l��M�"t�+�$d�]t���߅�����hu�"�(!�s;�Ԡ�!1ӐjEt�p&�����st��J[k��a���.F�R��˳q��{T/�%��R�����&2^�ś&�$z�^��)~3k����:�M��)Nd�/�_�T;�,�a�v�&j*���T������/��V
�hY𔝻�hiSyҘ�>��h(#:��x����X��������f<}��ȖȬ���\Lh����ȱs���:S�����DWR�Gk}!�H�h��t좶�[\��q	]�T�B�׼�Ӫ�er�ᳯ�5���ң(1�� ��j���\!�{V����fP�q\�Vh���S�71����&�k�{�yV�x��s#�c1XZ��D�:ߞ��b�]��(�R�D��m���,�w��7��	��׌�\Ŕ8|O��io��x:���侰�(0�t�	+đkl�;�����	���9<�U0���ؼl�M_��.���S�x��F�>��<r�Eٹ$�=��\�^��K<��.�٨�wM�r�����7��Ƀa��$4"�<#�Mn�b�O'��>�m�kG��X�6">�Y�A'aD;V�b�vFF�x>��4g��W���X.�e�^���T�K�U�a�����χP�ꯐ�����Cr��UX�q�U����Xn9�sY�1�S��>
�1	^�G�-N����϶
�.E)gZ��A��}��cY����1��qNU�'�7}�G�*�+����ʥ\��z3��E���ZZ���J7���D��+w�/��쐭M�>l#�`P�+�9D���K�vxW�#��o����W(xhl+���:�tu�s1���b��q�!@��^��B�Gf�<rj飲Y�u���و�b�z(��ldې��r�����	�|6N�+��x���e�
������z�������-F%	����m�塴vh�2Ґ������nw$�ҹ�N�:�.�$�ȫ��X�6>]X��%���Vؖ�e�c�*��%��\;����.�j��A3��Nj��r�3�;��Ě��K�#;��^\+uw�zW�7���x/�5&����M�w�U��K�s�; �*��sY�^�;�5��q���-��/��)�p*�;~������?�UK\$�HѲ�p�ݐ��띇��v+pMM	�A��#�bn�54tW������@�&"�Hm��BE�"@s�EA��zì}4��>��+��ܢ�-��[r�m �R;Μa�z"��诏P��.�t� ,*������n\�!վf�6�6�+*䱴�z��")����S 3�\մfIh2.�����s�Wb�tT��4)]�}efa��q�1�\����F������LE&Ϭ��
"���k=�&f��d�tͷ��s+3n���oN
�H�0xT�߼X�EgPpń�ð�R�1ol���i��Ƥ�қ�V}m�0��:j����23�� a�D]ʈv9[�!����{�L���r��<����7Cf2||�Q�5��+l-�
/���c&��׵*I�Wڵm�od�vK������{5�Ϻ+r-�S�Bz|ކ:YX=��}�n���b�4�1�e����A����om�ñ�!6D���Q돎��9�����k��:N�!ɽ�[�ʳ��U)�(&3P�mE)Xvë��νv�T�Zcr�]֫�2b���M�Y)�2p{����ʹA:s/^�Y/h���@G�oNkUƑ�P���֪��}��-�8s��3'�Rs���J=���򖝶/���j����.'�'���μ�k,;r�|���o!=쩏����/�Ї����SfaԍD"�Q[,e c�cxH��ϡ݋[�.��yt�!&�Om�+s������1�Ǹ_p�l$:���KFɤz���8%�OⳜ���u!���Xgg�z�:\_IB�qhs[ �2ܷ�EK$����i����^���H���
N�d������Ċ�a��V-�9�;yB��'�<;����<xn�ڥc�3�h<�:ˊ
鬉����>��ٞ��t{a�y,?nuZ|�� �p��.��Q`�wf�[Z�_rz�Z��Sә�^j"���s���b�Xa["��8��J���jHz�Ι�Tzd#~�2�b�P�e���o ���>�y�D�X��T�T�^�qY�7��,��\�G�[����'o�`����C��.��ZA�ڑ����Qu�}��wt�8�ʜi]�q�Y��LUX��q�b<��q]3�zwZDu.��c�X�(���w,�@��	W��j�c�i����y�������z���z�m��c�q��4��S3Gu)����=Iu&b�N����n	W3�#S��<2��u���Ϸ�[�5�S<2����.�(d�6��B����V �b)�����S�l��M�W�,r���bʻV�%��\IՅ�q+���u���h]I}[xuY�(N ���[�ܬ���R��\~������4�����5;��r��[�%�w�͉e_F��.�Z�M��rh 4�O���vLiuoۃ+��vcM�ť`�w�����X�}z4f,u��ࠛ�n<�e_Ww
3�)aҠ5���Ms��}��Тr��[���]��62WG�5V�癔Ɂ�u)L=�<̶����Z7�h�&��>�����+�ocXbZ��[T�J���f+�
Ј{]�B�]�m���e\8���7Ȟ����򶅧v����A�2'|����I�LmX�8޼��8C�8^q=�D�"hɑE�ؐ]2�{k*�#Zc!�>� ��CFɳ��r٤!$�P�B�xK�J����gy8��=�O<���T�=�Wi&��D�ǝM���M)cP�y��}���BO�D~��X����z7u}��(�rq��Pwʥ��ϓ��`Һ�����]� K��'����mjȉ(����!R�0�Չ�ro;;]�M�F��'���I+DT�.�k��RWӻ�j��(@~lb��*�e��������ATb+Z�TZ�DG�9��T4��*,aR�*�[��mV����EGV�U��MR���Zk!X���"
�EDb�V(����2�("V�Y"�h�E�� �`��(�XňȤ�DY�*�c�U�QE5KH�*(����@\�QTX(���*(���" �i
�0b�b�DE����-1�b$�Tik"�2���eF"0�**�TQEED�4Q2(�Yp�2�AV*��U�`#U�"%eUm,��PP�)4¬Ƒb�5�H5�b�2��QF2)Qckb
����+��*""���,UF#�\j��Ae��Ȣ�2�Tb�D�UC�EV�qUƫ�M5X�QAcTEUCV�b��*�~��>�<�`c�� ��y��h�z��qƑt���mf�4��|���!w4��{wd�n}�ڨ�[y�����C᩷˛�V���;�U��vˋ':�g*Jj��r(��3�QbE�!�q~�穗J�^+�s�S޺w�O��ݸY��[/&c�+k���x��BuѢ!�ɖ�q�;��9�6 ���A�.��)nsfԃ�Q��Nds�����-�k��qf�2��o��6�6�_��Xwꨀ:�`sT�D�|Z�~�G�X2\��'aA�:ٞ���0������v6۵�%9ø�V�'{/.]ջ��@q?l>�p�<��ú|2�d�ږeĒf:��t�x�7^S�n#'�a���?S�"6�h4`FJ�ʍ���F*�y�mD��N\�i�06�<�st,AR�hB)�-���ٷg��4;��
��9��SӢ0�׷�T�ߣ���̾T�̳!��4`�:*l)Ě@��U]��z�.M(��g*^��t|4R��B�ev&c�bj+��Od1��檖0�X0�i�7�ߗ�<u��[��ފ0��J�:	�"��{5@Q3U�m�9v�����
��Rܱ��������?z�E`^b�{�Htm�gd�D�c�A>X���>�_�>�pLɌ$�x�g{�ft|n�Xɖ�\�<Y֯>@����|S[Na�9�˔p�\�y��ȷ����G{u��hs�W�|����*,����d)f�"��>b�>Fʻ�X%�>���fu[�;%"ի���^���י��:�S8��¬��t�>_ D�R�]#VJnǮ�{ΰ5bpɜ�9Ku���Z���j���L��ջۜ�50��ܪ��պ�^_2R���o�#��T7G?uiy�����+���ZY&]���A;�\��N/7�Q�Y�9
������zel�(3U��h��3},�
�ɯW�S�2�Cu|ٸ�Yqn�vN��ꕞ|TM
}Q�cwW"P�}B�kZb��J�b�R�'c��*�f����;�tZ��eF��ܾN�w�l.�C�T(�E�
�"��ZD]&�i\@�1[͠`m�@�L˞��&3�T�{^�O#GT�'��~���c�Z��&g��gȗ�z������q��\��_yOEb򠆅S�ԥ1i����k����6j�R/�V� �`���>��'��2q���^^�UNd5�:v����ǳ�2J�>�^����˦34���Z3���EvRF�p���Y�fT������c����/��ك{�I���&���\O�V4��'�;��k�w2y�WǏ$��!̮je[́\9V+/�W[�!�A	�v��tM{w3W/�ޔurۜ����H��|0�vwJ���y}a��}i���F�/�����`��p{X}YHN����z��@�e�\O��n�:��*u8��vrY�c���iw����� ��Q�47�entSw�іBF8��na��VJ�TG1���Ĵ`�5�Me�yBۚ�:U����L�p��5ֹƣ���;�T��C�rZ���M���鬷'3��`h>�ٖ�:�7&yj)VN�m�Иk�����/��}�K,���i;����J;���f�{�ƌ�l_-������5qA�Z�ֶ�Oi/p�O���Ɯ�ԙ��'_�(�c4+/Pv�ҙY��׳Q:�;Y��W+1�X�ΐy���	�.�YH�s�Zq��U��[坆�0s�ϼs���dp��,c�'�^��8D�[�]H����J����٫������B�K�	�lU�93BZ�+�(`Lc���&S��c+L.�֚���G+$՝�+Q�kǽ�l���h�����P��g��BӻM���";�iV�j�:�d��˸�흕�͠�*��K���h�R���-����6H��G����I�0�0)ힰ�E �.!P�WUb��d\�d�~q���~eWy���r�Ӝ��8�V�c�9�~
z�F��8��[b���[nmm��r�;ذ2� ]-W�/��;���>�a��v����v�'9�s���� k�
���Z���M"9�#��M�e\ތ�� ���Ӝ��̇��@/m�ꮩh��D/]n�����"��Pn��ue�}�7U���� ��Ey�:CmC�*�z������ʔ��f��§W�ZHe<�R\ڷi���
NJ��e��A�4��XV7Q���O�J���]�iv�&Z��<��W������t3�F�z��"C������1�}��3�;�Mߛ���g�x]���A�(k4v7#�̥ݻ/J��7�t�,�tr�#{
�OxK}s�A���#&꣍��g=��|8��sF|�-Y�/�ǌԏM�y�Ն�"�8r����P�3���q��^:��b�{�c�{�Jb���]��i��ۗVu�9hng�9�))�j��6���B�]s�r�x��fA��^Ն;�9�,�ﾪx������"7�7H��v*��\�W(pζń�����ɔ�&I�7* `�z�����*,��:ҫ>��a=�m ���8��(2��8��ٽ��#����'VU��{7;�f������f��ҧ&��(__w[.���skKw����㛮�zBz������xC`�8��R��3̫��Q�,N���C}���-��jۦ�^�/r]*��P���\%	�Q.rn��<�^�u#s��m.:�d&ڷK�=���m⛮\6��f�;�f���PѤ	��,���Mߴ�:��18�ڶ��h�u�v��*{���m�Ң��r���Ӂק�j�j�K�~M%y�2��ެ\ur��/T�.�2��̵4���W��;V�az�Dl�W�����n������0q�OqX�rH����[������|�����R���YQ�Ϳu�7�;GH�%��?h�R���Ѽ�@0d�EA׊M�Fﳲ��މ��[t���	-�M��z.e�(R-Ԭ��딷{ّi>�����&#����<e,&�;��m�[1�r��R�� M��m`���a&wt�\�^_[g�r6��M�g�6ܬ�7���IE��e�yc>��$F��`�G��}ˉ��nÚ�Zz&S��{m�eV�.�5��&�p�()��4p���Ήo��������U��;�3�|�5$�����t�x�G���V{)�7��)C�iu�8���.�X�qǚ�İ��w�����hk��ro@�{}�㲕�J
��=�O<H��o���Q���a-�����D5q@>T���'��O����&��G��R���D�"��P˾�mykXlc��-\W�����+*�n�0�2�)�o�ڣ}v��"�le�\/Jz�������A:����g���֣���N>��5S��vnp�2��7�S�[>s��������}OR�:�8"��c�����8D�X3���W���)��&osOY�ן��e4=1V��UN����]�շ�!^�Gʗ���� +fw$x�j�w�n�18�>��r�'X�6�W�\zP�,�
�d�yAWs\w����zζ�Aqϗ��wir��bh�ބ���>��a��!�Ek[�����^����S�a��Ժ�C�L�~�B�_��vVǶ�eٍ�j�w���X1x����c��r	��8r�-���k���SM�p+���N��_�iUn�<��>߾�8���2�OE���c0&�M�;YV�$�j����V�;���O#���6�H�ۊ��WF�^���b�l���E�*�zS$Gj#7gt�+�<=�l�i��R��*�(�-oq���ja�jGY�L=x2V��]���N������5�݇�j��אWV���E�eW�S�UWV�����¯(q!���dʛ������M��;l1Ag�!`��򖧼W�* V���8��u�19�^��=]{ˋ���R��}��Q3�����e�y��9���L�h��Gv�*�b��#+���a(t�Q��j��M�=���4ƅ�6��+(��S���ޭ'�VVޒ���A�}�e�ż��D����2Mov1{r�����Z�92����Ѯ�@���Gx�D��<i7l��n
����[�6�Z�]��P���"�HՓ)�8�n�.V6��4u ��Z��CQ���w=L��h�0F��-�l�7��Z�x�j�WmUօ�Z���q�L-R ���@Na۬���B���;E��L��ʐy���6\Yxޔ��+�`j�H�>jwK�YH��h��4}��Q��9}y17�r�^�Ӿ�c�p,c���Aw��q�Z=�"�bޕ�i�DhVot8����d���εl��:� ��z����*��U����Y5!�(�\�)n#̷��Ҹ�P,�J�,v��V�6l��∓k8�Z���^"7�+����i�j�S���s���tD�{QOzaB��&��f��O}�h٨2K��*���&�=�����po�9�zSA[��_-��6�K��/*^�S�BZ&;Q�ׇ%�t^ѱ�3�����oB暶���d
J)�:m��qU�z�oH)��O�䊵�!�+pm��ЕΎFf&�zL��a���0]lf���pE�7�#��(]>o"�PX��!��}�܃
2oIY��MF�XI����s:�v	K$M2d�Cc�e9�z�D:�/�ǉ����Q�,��
���NGX��:����d��<:�6�gM��π;�9��-<�}I��(j22��'ͺy������=�ݭnb�%k�*db�]���d9�<��qR��5������'W���eT$��V��˦�o�'ݷA4xY�Q�A�ʊ�Z�U�'��d��	؝:����e�K{��	C����o�jnG> �����e����U�J��38�!�h�N��	����"�?!�<�dl�I�/t��#��MNaW�X�]��B���T#����s�So��f�����qY��w�Ocb���;�X���LY����V��=�C�I�2��O��^������^�[ޅ`� �8gj�TD�;c�9;{��G��a�a�鯏������|�;7���ފ�臾�2�ܺs	���]:����;$?N�\vW�����jå��\�u��0++$٢пWV3+r�޻��Z)i1f<�"��v̤��<`㞞*�j�W;9��2���C�ȯt�L�)�&�Jn�٢���Ʈ������;6r�E�Oz����e����b�/pr� ��Ȼ�h\*�v �J�_<N��>�6_�07T�};b5
iu�n��q���N8��aa�Z�K��_�J;�L��+��DH��8O*<�V��sqCXM>xd[�t�=��Vf�狮Kl˰��~T���-��D��;z2M�ƙ���&
�v�Omv��}i6��ח���WW�P�5&y�f����i��i��#wJ���M�֞H��65�f�r.Z+]�4�Y�u#_�"1����9{ˌ&^�5a��^,�N������X|�~Σ���;O>�&�FH�E7a8��aR�]��z��ݤ�=g��ԑ�/�2efkmI���Ҩ���ފB��<(D������Qu��7�k��IEK�mfwq�^]���o��4��g٭#���U���^{]��gf�����)���'0��~f���]�X������pˌ�ƨ������|<��9�2�+S��jG������Xw4�3|����=�RM����g�A�#����u�5��o�������q��뻶��|���v�Rr�R��o��D|Q>�ό5�Ԫ�w⚸hĳ	�f���}x,�0��zi�eZ��*��|4������-�]���
�2���X2��*6�푽���o[�+ƫ�F0sK�Q.z��^]�q�XE�X���t������])�],�"���{+�8^�Rr&�[����&�����7KFY�� 9�
Nfa{�V�ɔt��.���R�{���DV#�k[���|�1#�Z7�YQ.+{�>¹�R����-f�B"�D����콵��*��4*�A�:W\�����FF4�\2�Ǒit�w���5p�/��[|��k^Gz�<��^vDc��p�=�d΂��<������o��zG�"�vU˲r:�!�Q�m�w��B[<	۷�.~|&���`�q+[SM>;�1yNp���5��'j��B��ӸL�:A^6i����u�u����� @Qn�i�[y�F6��vE�����kk�e����^SW�_t�`�V���Y1��ѓ�^�WW��Ϲ-)�H}���C4�ߛDG��׳��:���ʸ���K �z�-��3:XXO0�l�/.s�S�5�������%y,��`�^uu�dE�x\j�'���ШX溱��nJ��zkoz��؞�A}~�ϣhzF%��͐`0e�����؞ e�#h�kn�2�������ih��o��&��7�n5�J�8{���ąiL2v���)��C�8v���i�u��4�N�эؤ�DyQ�q]r��t������M�M�����*�e����N��7o������Oxob]��Y�N��x�����pu� :�=\��rG�!�ӻ�k�}�H�8�Cw&�tiZ�7��f'�W+�
��uw,R{��0�b�M�޵���w���fQ�N*���6ձQR2h�vC�Խ�,s_У��Ǳ���Lx��TJ�X���b���ԻN -gi2��;��w]E�J�H�]�1k�Si�\�;n��[?�jCݼ��W���t�T7H�Űe����4�yL���{��準+����J*+^:U������{�!�h�oz���v�J��$`��+���e�<�����s�]skj�Zٖ�����z��;�˳q6�
�`��Q##�(H�R��%�zuB�˰ڠxe��L3	_��I�����V��,�p��dv�\�������R5����P��+���ۣJ7�y�痡k���m�[���l�=|����u���� �o[���9���k-ҝ�+p�MX��e��V\8�Ml\x�h�f�f����~�s��}�Ԛ"���1EAVE��
��*�-T�UT�*�**�`����dr�D�A�"���"��UUQX����"��1G�*��5*�ETA�X*��*��X�F�(�MYE���!iX����@UQA��E���F,TbF	ZQ+F*��UT]!X�#A`���1��(������VE�q�TX�EU`*�TETAcUQ����%��Z��E�0T@`���EU�ը�1X�� �*̴i����(��V"T�TUEU"���DDUV
�DV"�V���
�աDV�DUU�mh�EEZ1X��QPPX�eAU,�&��UUE�Ȍ��-*$F-�
��A�*9lDP`��3�Ͼϰ���U=|��6�4�|)���b������v���r�X���v�O���H1���W�_zN[}$���
q���E��9���۳�r��5kXlc��!������d%p�Q�§���f��YT{���0�lP�ԭ�=[�^�{#K����0�Ε����R5Ǳ�cN��b�-8�g��w�[.s�N��q�y[�N�ק:L���('+AŢ��P�@V=�����P{x��W�7�{<�g���XmE;��جUX�:��]'�ѵ.c�s��l��"B��X�(�V�9씣�Ca2$h�b���1����R\����R�OW��>�;�����m�v�V/*��̱�[�8ṇ�����ۮ��Z~��5kk����#\�-#!��U��d�Gm���f����SN��Օ���*�W2%��us��Ro:S���M�o]�+
��Ҥv��'���0e,�O�⧍Cs��k̡<,Q�w��OE�uc5%p��j�6�U��>�:�n�r.�~�
ǧ{O��UڅM�V�6�V!�ҭ��a���5eĚ�0M�20_8a(_S-魱9����o3�N�`�a�F�C�?{��=���x�Μ3u�D�{�v���2��%8�CTN���uMl�Km�4QwR����3�;y��;��5)����4�qBP��e^m{�3&�e�[����*	���|7��J���|.Hj*k��Mfk-���l��ֻ֝�]<ʺݷ�z]����,XJy�u�l���>J��^y���M=�f�{�t����]�7M��!^˶����ְ��{T#c*v�N
�������͋t72��z���-��>ƅe����u"��il����0�3S>l,ިU�Auy�e��=YH��h�bν��"/�rX��L�>��uL,���y;�(.�z���x+�s����UkpH:�r�V����KR/�-��;yOl�}�aq�؆褳�W��w6���'�Q�e��JM^��j�1��:X��d���(j*�+��~PP�����Q��[��7��.jվ+2\Ƿ����.����Ռ�O S����]aVF	Cl�hK PIY���t7��|��j�����m�y/�Y8�5}�U�1��k��ט�|4#����2���gE�ys*:Msw$��U��9[�Ux�W+VS��ݩ�p�֬9y. :2hڲ����5!�����:��J(n�j�q�4�簱�1]S�j����\���_���c�^՞����Gj�/]�үF����\����Yy������v��)F���m�`�&�Q�ѷgbv���
�;��`Z��ĉN������Rp*P�de�/��-��4���lE�{5��T�~�?��h7CO�J�U�\죌�����묳6X��9��Q�V�K|�Uy4���y�[��LI��tu�ޡz���km�^Uښ�De6F�/�C����ЕYL���or�IWƎ6��nj�2�̃;�&�C\n��W�.�.���0g[b�s��]n��d��7Rǐ~�v�Nj��^�ukj����=i����6Q1Դ0/
�������J�F�"��ef��̽l�܂�z�ڕ�gg��n�RJ��}�2��S��ˀ�x���z]:���R�z�`y0����IY&;�v�Eh����7�w~˞�����x������a*"z�}{�I	~�a�~�������Ü������'�>+75��<���Ay�壱�iۋ���G����<1`��e.���N�倫L���}��j
�����F�z�i;�d�)���;7��ԏ�v�c�'�ջ�\�f�r<����ӛ� �xߐ{Z���g�m�'S��A���CP,��W�K�͸���L��|�^�ZS}����v�zu
-".�w�+��vv��d����{��N\	������9�1ޙN]*v+��誇E��ں���,��c��꾽~�h����}r[f]�K���A
�9�-�q�pIy�u�Uf�*E�\��~/������I��ۋ~i{m^�ȹ�X3w�Z��1�S#yo�cd�*�W2%�����ӹ)(N2��������7�N0$m��
|s��cd`�G�G.'�S��H��S��b�\���%ܟjC�P�W�vz{���:M����/�Q.$��(��j�j�s]�J�yR�+&�U��P��.�������'��}�nW���My&���Ѝ��{�w��f���:��I��]ך���Nu���	W�ub��:!\�9�K���������"Pg\�Rс�9�M�N(�)�����{����mM�z�;��F�d�`�5���uyV��:U��[�J�d!�3˸��(ח��;����	�7�%����*���gw���Vv��Xs{����-E*{\3O0�6�an�kZ���*�ѳ^�T�9<&��&A+%�z���x>��~Ao�~ J�E�x���|�-����^ܙ�6!L���ս�f++_�(����}���IS�ռ|��B!R�����㒞�'��%i[gH<��p�ջ��E��hq�#Z.�oЮ"rƄ���3��5K�*\��]*��S�zG r6H�:��h^�R��#w�w�(LfW�n ��2�js�g���XmE �.*�b�Ub��@���5��m�a�r�8�{��K����-B���V��d�
z+̈́̍S�K�Ah�
+�=|^,"�+
�ẺŞշ�wv
;Z��aTF2Z�k�0��^>���lV�Ve�-��
Neι��UϬ3l���6���@4*��@7:�_9��3���^^ ��g�U���������e�;tD��׹�ZL��`�&l�������v	�O!�u����m�v����&U�4nw��� 6�9�u=�0�(�ڍ���[^�����FE�g����B/�bo*�;i�0���]B[&;Qq���*�>���N��9�yu�J��Y.�u]}�d��+=C��&�*����[�;69���y�]<�RX�Wä��O$RqBP���eW)�}�,e2�a~z��c�����W;�e��=�|�^h8�5��Z�W�yX�f�JOZ5��^� ��s�>ފ`��M9梦�B*�C\��m�P4�+#���Z���957�U�]�"��9M�XX�%��S}��s��K���]��vq���XQ�~��U��.��i
˶��r��ְ�.��ia�yzJl���D/~��o�<�'��VU����
�^���F��JI�%e���Mv�:�VgY¶��v<�Vu��F_;��|q���&�u�=�݄JrP��+x�W�$ Ѡ��E����)K�W��I��Y&Mc�U���|�����ɭ�p�r	�Uj���w��gv�ݒ���އ� ����#}�G�G�����W�{�y�f�;��e".v�h`�s\��#I܈Wy����ԇ/4�e��;7��{��]L��A��V�)�X���o�Ŏ�;�qn+�	��֭�e��b���z��vhT;��e�Y4�.)�0Cqq��<ڱ�q�8�V,v�J���/`�X4�{�H�#}Bu�#T�'���7KU�|F��F�}��hO�L��u���=��}61yPCGW��p�_��Ȳ�X�w�ғٷ�b�IkE@���α�C89���^���~��Bs�KD�Gj az��0]���g6�Tq�q��+���iԉJo΂'m<�8\^��y�]�YSf��o����~+�������y �Rp*P�de�o&TD9o8�3N�`�3�K:4����>s��z$�V��}���R���x)��f��)�^�^h���3|�$Yn�owP"��Dգ�
��;g�N���:��q;X��qN�8����gG�]�o�Wrמ�J�[F�٩�6�Ό(y�_�F��)� ��z��sH�qV�zu^,�14����kCމEM>e�3Yb�{鮷t2ANNR��2������ɠ�r��#��5ޏ�<|� `���i�c�Ț�wW�jpU���P���S���)G���}�5�	��-d��3��gӻ��W�v��t���F����fd[oy���5�;Q]K�ɭj��t�k	�>��<1ʽ�W�}�@Q�h��B���|'�����j����A��e\:�3��5���S]To��]���:�Ԭ"���{���{�q��d!�ې��?{�/��hc^�;@�8��25�n��9ٸ%Ҹ�8�ziVT�����/�b��Ώ�/��O!���:���{������<������zc8�I/|*9#��;b�P�ҹM����j3�!�%���s�j+9XV��B!5mù}�=�r24t`v'��dK���j�r�l��^c������q�6j��W�c>��t�\4m��++}P��U����<��Vǎ��ևw��rd�w�n	=҇C�j�m����WsD����+]0���ډK�R�I�g`F�c�x{F!��\��w�X�2��6�m��Ÿ���so����z�ͥ�c�閕JaK��䆅�s�.Ό{Ol=�A
Ci�5��K�ϸ�=�z�I��|ۊ��留ȳp۽�U�Z�D���-:�R�>ڈ����*��D�����m<�V���I��}\�q�ƣ�UH�����8�c}�)��L�3Qb�w��l��Ҥ�;;D���CQ��Rx�8Q"3�����6���8z�3��`�@��54�d���ں��m��T>��o�2�0F�=A8��^�錄l�������|"�45�N�98U�Z^����P���f�����[E�z�In��a�����>TѲc�{�) gx@f{=L��}Z`�%��W�0���|�W���a0��n�/#�\JF��k�xv�*�|}t�cc@�Ԭ#��g^�
6K+Z�7��p^z����55���,�)��h)w�w�����6޸����/Z�&L�d��E�W�N�fH+���nB��n_i �]n�ì�1O�$�r������^�7�J[�+�ޤs�f⫔j�h�e�-���K��o7�(�jJ�U��sr����-8�gZ/9��0�M	&m�p���yh�=�Y��t�z)ؽ>�ڰgZ����1q���m<����ݖ^�$�b�!��s�`S�=a��.!P�S$_�P���sb*�##S׉����y��ޕڅ=ƣ�jݹ�aOCa=����cI��\d��n���KF/̮��������r�k�;��2��z꺾V�g����&��N@Kq^=����~;�ߋ�)�,���}B��f��~I>o)a�����5]Ո�Da��Ҭ�s�2D�����yʍge\�_3 �I@�ä6��Up���Y��Pn��gr�'���{�:�w�y[��y �N*P�f���ruO�O][����Ǜ��sx��~��HΊn�D�Z�{`���4�qkɬ�#��LHS��_t����Q��W�:6[�E�9���ݐ��ls��O�T8'�X�����v%������P�vf��Lft��邍Fg��]��<zP�yh1���:�y�� ��4��彧�A�/t���P���JB�g�R��ч���41�Ӯ�}]E��|_����>��3���ܮԂk�Z��L!��P.�߯?tȢ,�c%���<a�T���lW�h[�yw+.�'�I5E�5<����c����Wo6k-p�-�!Dz��y��}����W����v�xtЫ͕;�&��b�8nݰy$���u'q�3��]��rhu%#zsL�h"���,��t<���w%ߎ+!/���c�^�;����	�����c5�R.��DC���We�06����걛�2�#�p�{O���E؁?|�Ϧ�c@�Xj,ٷ�pu	����@u���b��/)��kC㕘4���2���ފ����0��lk���4��`�P��vR=�+ޓS�e�I��D����� �YY�>]��fP~����E墺�By\ѥ��:�'HM�Db�y42�]��pEK�ۮgJ�''���3PT���g"C���u$$�7enht3r�CL��T�c�����8���O�������"qd��X��,E*V��X����EL���.Z:�<V���j3��2]����U̍�peZ��F��I�MeM��j(��r�H�|ھ���Z�ѝ�����f���rY<c�I|�WA/�����+>�ČCbo+f�qladnㅵ��Z����CX]�D�%VVD�;yi�ƍܑU˅�Uc��diō%��r��MZ{:�H�Co���95���l�݋]7��P5,G�5�� �A�������ilg%�Ivв5�&�')�a۹i�иT�Ș���q!o/�-'���G��q�p�n�v[���r�$h���)Q�4�Ȍ��7x�ch�PTD�-q�t�7��������;]�.����x�q�Cn*��9����j}��hJ�ھ�\�WX�J.;/�>�u�E`_��}�ʀ=���U|oZ��7�V�O�+�LKTh�z�]إH����/�,��P���K�r���{]gO�&i�g�r�����[��g1���vs>�3Ge��C��?��´�_<�ezC��^!����xgjJ�+d�N����r�M��ܗ�ӹD%]:n	lޑ��Ō8��v��f 4����a<�΃vvg��6�
ϭ���d���JŅ�3��
U��ۜH����ˠN���3��PU�[����e��[��Н����[�z����e�Cj�%5a�2��g�҆��e�Gs;I6ɖ]�kwCӎ�}Dn�������x��s� +��/d�y��VV�]p&1�B�vq[D��\F\����x���U�yZk��l�}�vB��U���ރ��g�1��"��~˘�Ї��[���XސU�� ��m�F�>Vy*A*T3;MJ�ͫ�������Q3�*5���EUb*��2��U������Z1-����DD��T���T�QUDX�������UV-eQYX��,QQ�娋��M5aATTP`��b�j���*5(骈e��Z1b*(�F"��PF5��D�"ZҢĭD��\¢���1AEm+[Eee[j��Eb
��(b�LJ*�**��2�1�M�#aiDUQ���TX��1��"�UX�]\�(��V*"�s%VV"���2��X��T�+`�4�Dt[�[UTb�5U����UUQ�R���1Uf��R����G-��AUDƌ��*�(�l�UQY�Q��E(�)�J�Q-�%X�Z�SV*�T�("��EX�+�Q&4H"��I�U��t�$��u�"�fp\�ͦ�,��W1�h��*^DSq��S��c��1��$��oh*�e�����-�++r~J�����J ������l��w�ֶd��	�5��*��^z�tr�>Յ�	C����}�gw`A��r���l� ��!W�RÄ����{��-��=�/g�>�T��N���QAn�a�����¬VQn��Hf4�< cۣǗ{�<���:CY��t(�y���}�P^u�h�i��uc8c"x��{*�V�1�w�-S|�;5���^N�
���شx�H��:��>=��uv�g;���v4��ջe���X��z�}�.�ܡ��3��Տ��;�'zd�:����V4�#P,�i+t��ld�VT�3@x�=����H��8�	�(��V���P�#S�G���?��O#�/[���P1���-_���4u	��JQ@�wKWx�okqs*f잹^�z��w���tRSD�I�B,lWbJ&���<�dy�����c/������Gm��Hѧ ����n�����{�E�G�t׳"�l���m�y9�7d����n�{M
��a�K�j٭��"څ�+�)�=����4*���ע��DҒ��	>ߺ�c���=g�C>R�����=r��iG�o�n^�c�ǫ��:/O!��d�fA�W��CJ�P�U�*3�7u��J[k�bx1�̦��@��6pZw#}I��J�ս�.�u���=g,E��<�ǎ5�ent2�U��e��k�T�V��>�9�<�(:���t��¨�(�E7~n*����Oz\jh��XRMMfWz����u�Kׅ�T�8��ϓ�^�ͷ��''!�̒���Y�C��KPe�����@���������1��;����S<����p���Ҭ� 5q@>�����=i�ؐ��;��Ȯ�{�s�o�R�t�\(e����|Vn��\��b��FΈ��n�%�iwP�F��9�b���M��]��#u��XE�OV�׳����R1���:*wb�QS@��eA�aKϒ칧B�@7Z�^��hv�`:�2�O�;O�Cpm]�4��fh篬u� �����b9��.|�4-*yԫ��Y������  ��܂|�I��]}�gY�ee^��bz&ػ��g�9(��]ҠOh�GI�����-�8�֋��g�q�����Ϲs_KRI�Pro4��T�#��X3�\vV6�@�����Zt��ϼB�Jvt��`�c8�9/£�C�"v�j<ZD]&��],�7���%�_,�b�>ģ�E����~S�^�9H��8rͥʜ�2� ��mћ�E'e��ߓK��p��%�eڗ��
0����3Ou��Jo*�";���X;����W���U#Cn'���2X��ڧv�&�1��{>�DU*��!����e$
�7V5a�ꓑ��G)��]s�޻�V8��dm��>8���\��O�T(��,���i��B��ѩ��^u%f9~�%)xz�g/f�ǧ|k�h�2��Jrc5���ձ��6)$�#���h2eg54��g5�y���Vy,ez���b��fk�ۻmO�ݺ�׋6�I
<+�����-f�X6���}�A������=�Zj}�;�Eb���C��C�2
�1M��~Se����9Z{�/�<=� ����������﹭�Y�nR�nN��Ȝ�SuZT�����S%��^�|2HEf���ץ/wؑ�gj��L�SEJ��&m�݆���c3���>{]��ɭ\P�ޘ��?-�Ud8�s�z�5���\��Wo�{`m!�P{�h-k㽪�'��S���{���F���jo�ʠ[�t�lV^�a�+h���&���v�R�c����hB���[��F�k��8�A�Ʌ��DRL��w��#�gY���Q����'{�A9Zb�]�ӆ!���{jr��=A$#`*H�@��q{|���XmE �.>T;��{`����jֽA�ogh`�)5�J�F5Cjݹ씣���&���XL;����{ѩ�;b��~�G���|���q_��c��2��ծ	�#��Y��>��U,׮KU�AOW�������m�\Y�����x�V�Y�RB~L����H��+iy5g2�:�u���)���K���SC�n`)��o�&_Lkj�����V���'@�z�m9_ժ�=O]��@��b!7F�ہ�N�V�b2����T0����}6��r�+Zޑ�85�NC���=g�C>Bv��l���7[��;��=z�9���Kj݄�I��i(��F�Ub��h�Z�E[L�w�s�5��5�x��e�Vw#|)8�	CQYj���Y��q����QOrV�,2�K���}���4H��>��Qbh��CY�	ֽ[�<��	�/¯���ҫ=�H��M}��j*n��7�c����·��F���YnN`�Xm�G�M�cR�A�uOXW1$D���a�ZƛޔTY��o�S����������!KP��l.�b����N&�;��Yo/;�v��4c�O�MNaS�������N�e����]��%���
�/Jef��٧���3�򲓝qt�)³���uf+�ZFh�F�������{�c�v࠺����*_s���IR���:K��1�aj��ّD���1�'
�n�1ayX�٤=�3*୊9�ه�3�YHѼۃ���i���$���ȭ��(��m'ѱ�;��R��^�˜(��J�]!s�Ȟ��:j���=�g�G-�-���`��2d��Ž+�M�2�s����7����v�Wz#Hx�A�j��e�EZ~5C����G�W{�>���������;aɉ�[��)��l.���q
�B�i\�\�ϩJm�9�e��T�6��ü�m�}7m(w/��b��!��NBR��貵j���L��Y��^"T c����;�iN[�A{TgCU379V�`1u7�{��X+D�r~;�_��S�V5��-3 �����6����׽�}�]k��H+�1�I����Ϸt�]P��8����j�'�Db;ۼ-q�"q�#m�U�;㍑�igC�ɣ�Ί}�igp뺷��߹qd����c�p��O�rr�`�Q�M��qP݉����k��s��S?P�C�����CY[n�W�.��,�9MӘ�(��{���ᡐ����g�^����`v�k[z��b�l��u��w��v�K����&��⏎�^�wG`&�:4Z�9�=�H���ʉx�M-3�C+4d��Q�^L�:R�V�J�3GeK�B�/�m0�Dr;B��pc6 ��כ�Pf��g>���C3��É׉�Wx�ܒL�Kx�Lmp�<ƥ�����ӳD5qMխ�:yd�|z�nG���ֻ�}�nv���u���C.�w�����k��>yqA�{ڹ�r�� ��Z��B�{��ޞ�YT>"�>�^��E�OV�㓼�d'p��
U�[hN-S��Ţ�3�nzV�\�lv�L�V�2���]���^r<s��������'{_;�T;�X�knz�PiX�\ ���I��o^�XNo`X��N�,v�N�%���*i'P�ZZzzܕW�n뷼�+IZI�<�
����m[�/%���C����Ӂ��p獉��{9Y������
H�+US�ɤy�v>2۩O�\P�� ��öz�e3׶ '��^���v������pOq_���iTl7�q��S9+
�ҭL����]:�ˬj���ќ�#v�lڼ�1�oH⯍�v�$�̻��D�y�^���܁�Ή�|e8m:�k��I{��W]Ć��W��&�D�1$��E(+�Kc��ͥè���K}�Bf�o�3CtR�_��>L/m����O��81�7t�+�<�^�υnD�������{�Y����ls"F�>��_�#R#�,7Ѽ���`<��U�\��w�G�=)�	CQ��WA�:�
Mʣ�	�Yo�Sշ�{�ۊ��n8����d�C\N��yz*ݘ�5���Ky��X�e��Q�V���	C�&��o�Ij*i�����]חc����Ǝwj��S�f�ժ�y}N�e!�[����-�Mhj�	j����=�,��R#������:�v��������A߹m-kv�;:m���{��(�&Q���!rW/p��M�S���7Ha��ԆB���*�<Úu�K{u�����f���h�{<��|;V�Ք�Ζ�;v����LIK+�[��8��O̶|�;7<])�G;�V��-Ջ���Y��s�iM����^��5�}]�����kL/���W�2����!���CW��E��$��W櫜���[��z�Q��E��-����'S�p\��;R�j�j;٩n݉!�%��Ցw�լ^G���d��S�8�d�,���dL�Tʾb�E#9:6�-�qn+�XZ��I��Sl��ģ�w�j)�\UįJu8�9e�-l�1x`�'=�6�n��1tq�M_�W���c��049���[�=�mc�*q
�Ty��|���C��_��cᘖm�g?Xy	z�ē��z�K+���%(=�E����n���fcf���̣o����2��2qo��}U��H��}�=W/v�i�V�c�|�����H�Y}a��m3"R���Hm��q���S|�Z�#RqqZ�L�3����JvÒ3�<�}�N*P��H����a��l=��\��gF�Ήo�Mh=�=�Z��C����8�!��n��%�O�8[��y��;�JK�N���;��%A�(ǂDuQ"�T�w4v�\t��"���YYn�W�v��*єޫ�4%��B�N��U�'����ntx7�K��\R��o��9�����npb� Q�R6 |��2w-�(�r���Ϛ=�� �d�m�"(��e���d���^2u�ph���u�Dg�,L#�`�S���i�X�b�Oy�*�D�l��eHY�������ܿm�"Eا��q{�+S[�hq����^8!)�j�>��<+�,���_�Z?y���z
ӻ��:C�-t+4h�zYV�u#
�+B��^�vz@L���f�lkb���	�/X�	���߾�揄���.r��s���R�[!�vn{���PPC9z��(w�E8��bdN�ھ���ΖZM�Z����O,~��v!���d�{��5ߩ�K��3,UX��ȹ�&�J�@ƒ"�N�7�y��e��{KS�=aOCav����B�ZF�j�/�YYj��jz���X.߅�B#Z�/%�S�X�%*f�׷$�~���nض���~�8�B���w��簻\�iV����j|����y[VVi��&�鞌C�20�v�*��S�Z��}i��g���}�y���)���P�Z�����s�a�-�x�
�#Q�6rt�[���e^�W`��ʍ�+�矫y_3t8/:ղ�J�RZ�,��D�h�h>9Q8����]bp�K�Vk�zn���_VY�+����cM�/��`�j���*э�¶�1��&lv'uJʊ�0Q��Le���c5{���:�ݝ2����H��v��h=`�Q�C�K�S�\o^���
���+�lV	y��T����+{���Hu����ky-}\�X�o;x��T��Q�L����#n��]���f�.Z�1����apӬ��3h����^ZA/<$=�E���zDcfHR�ނ.��!��c��\��V�Ԡ��$��vmU�pHP����lx��3<��"CG�An�nÌ�Zo�ף�rp�`(��C�(l�\x�а�ڲ^]6�I4�z�t�f�]_��^KzG(~��[{[�m� ���eN�0�O,�5�]}�@�U���^׆�=�S'h����DvGC���&啧�V�]J��ݭ�TN�{���\%]��իL�N�<ւ�P*�3�F�]έ>B�r�]�I;��W�]� iOU��w�u(9��=ml.
��fZ��=vsX�dɣ�hk���3vD)N�PlX���ɛ��R���Y��Ÿ�M�����J�I��^�2Ĝ���l�3Pȹ��>ͻ�8c���#�ǝZm2�X�	R%�:��*�p�t�8�T��&�t��"F���F��b���Z�l��%a��V>��XD�"t)-����� ��S)ү���CU���w��+���WQ�`��^R9 -
�f]�~Y�e�~U��%u�W}��c�F��د�,�2���槴��B��<��t���m4H�\f/xa]\u.X�TP|�����{�k-��ew]�t����˖�\��Wg��)��U�i�ƅ+H�:�u$����' 9x�l��a�,�c ��q��C��VJ(���j�H :M��e�n���ۙ�Y��|m����Z�Kj�u:�b6�KZ��$-���9��'J�a�"�֪Ç�kIB_|��=�w�H�$�՜1�r��[xu��n�B�X����n����y�=����������ƈ�_9,�N���N}�Q�۝Z���'xD&�^⨴�fc�6�tF��f���oO3.�����έ���u��A�
��˜�ޅ�2�N�D���J�ޓfm��Z�1�N�n�l>������#w��L�&���o��
ߛ�y�y9)����uw����Nu|��A6�
���ؤ��\�2�������ҧz  ���!�ajb��V%�̬S# U���=pQ�2~��.�=�M혹�f!J-�q��n\5���F8���
#x����N���s{���Ѭ�}ӹ��}3�l�t�Cv��y�Z�X��U*;s7v9$�����~�F �z�F0D�ł�*�,U�C�bcX,T�,PX �R*�����*����\ajUĬH����b*")�Q���X���#���PH��lX��X�QDV"����:j�TH�WQF �f5b��(�-��F#�Y@U���1b����@T���0b�j��Db�
�i�GT�Gm�,UE�ڌ��%�A�����b�(��F"�1U��UQV��X�,DEETc�TQ�,v�"(�������
0UDFn�AUݦ�A�n��DDQ��"+QECIQU "*(��dLeTt�bcA��"*�E��3&A,SM1*1U�1DTX[,X���(���l*�Wm�7�#�EQѲ�(���QQ��ԕ(������EU2ګ4�X.�`��]3�YC�U[�z0�}�����ݱ4��&3�pY�ͣ�J��įT�ۏj�,Ҭ�������_Yf�uo�sN:OSjNc��*~���i�`���~+���}`6pZw"��׳�r�D�2��/U׳�z�����0�z4m#��eߓD�h3��_CFf`��k�핝zT���%���(k3Yj�����ׁ¨�(�E7%E�iQ��>�{�!�r1l�zxY�Q�ML����襩8�.FZ9(���7�{VL���(oxN�%��|"_q�s��W��W>������cZ1W��KY��Xm�٦�c��t��dLl��~�2S<0i�=C}G�>��	^y��U/���I<^7��φ�b�5L=R6��K�z�eQo��C �e�V/Jz��{�T�o��sϔ^j��-wB�s<�8D�[��D��c�Ğ�Y�yu��V�w�Sy��њ{�jH�'~�L�b�]�Өc��^�c��G�ƽW�u.u�P�b�T�Aͤ��P^�.��|�t�<�.h����y:X��,k@u�Gy#
5�D��N�����l6-[��gw*�[zR��m�d��}͂Uh�%�f��dl����ԧX�i��d�s��W${{r��:�+2�h�ܴH�N�L�w
�`6ڷK�읱�E;���F������^fP���hΓ����)GH��j݀����##Gp8,��/3u뤌^�*+��/US��4�=�#\�ٗp��w���U�0�:���1Q��d`t'	l�ո^��m�S�V5����쓧�o9���osz��?v��b�^Ҳ���qVo�t�+��g<��4&�5����TNvU���:Jc���dP�1��I��}�f�&�:w5�7�畷F4�I�T��'
�N����&J|��Lĭ[i�tSv���d9��ɦ�$JȚ�]�/ �ͭd��h1��V0t��茦�ފ@��:�hM�d������&��t����n�6d�f�{,h:<=��;+K�
���Z�{�s}y뷵�-u��x���I�k����ƔI�������dd�6F��=�6�r�!�`�ùĝ^��y׋b���8����wZ�/�b�lf��j�/����<3ٷ=��ֲ-T��Ov��9�45o]�.*(;7#�n�� V��n���r��V��A++r	$��~�
�J�Ç�Վ�^����B�]��]�E.^p?C�\Jo'�(-���{�Aw��f/)M������p�bW]����}'���S<׏D�:�7��m9A:�m;tqOO��u/X΍�Rn�ѷw4�[Y*�V���H�M����k�[ފ�����"�2B�5���3x�����.r���&|5�ϓl��Ŋ{g�Q�vV ����Kp��+��\���2Dg{���]��g�-�v�R��Q�E��menu�}c��Bq��U��|_:��G!ݯ��0��ˈRs�
���꾹c���碆/*�	��JQ@���/U���bE��8��[���{�ĨI���1u���ۍ��{mL��l��^�.y���ƔN,]��+�+������L�4�
l:m�C�#	���I=���D�-I�V���z�Ef��P�u���b�g5��+�+��3SCk��N ��|I�T����<��x�ުTnR��́J��]6e,<��"�7�s��sv�i���Iif�Lτ�x�wY�|�Jͣ�e�"?K����{#��E�}�"��,4�	#�)f2�&S��ӹ
���Rj7�v�W���{٭�G���
@<TTxˋ�	��T�sa:
4(7V#��؊�<7+=��y��M�3U_�*|��]� 5>�v��yN��Bt%S�@b��i;b�	�O,h�����]�۝�7^�=�%Y�(AW';x>4��sz��1�G)w2������Vr�h���[��'�G�D��{��/�s)rnT"�nv <� �h���V���=Y��p�v�G�#|�5�b����>�|Ɛ��MA���Y�;����]]�ؒwG;�i����������v��2�6t9�(��bO�1��
57)84�[�މ��Kf/��Oƶ��:�@a��Aʿn��S����:�7W�\��q�ٛZn����Ow�^t0������*��[օ8[>O�ڌs��q`D�V)s@�YGj�I������{���`�x�ϩ�tlf��cR3s]�):X:�AP�8���\�l�ZE{4��:�EW|f���/?v����_n_�Z:�-F�D7��*���:�h%Mf��@C��C��}�p��#s�p�T�ۋ$}-���{��Y�AK��NcY:M�c*5v).;\�P�)뺶x2��E��8������=��%ݻ����%�^�
��"�؃]J"�(l�3I�J�.���K	����/8��\�8�Թu�."6%^!� �H��J�L�9�pj�`\�Ue�n��b�W!��,��ovu�*,c�8�TJ�专. B�Ӱ�'s��[f��N����ZXѡxj��VO=�q�&;�P�)��\5��N'F(qG���ܑ>��zF��|ߒ�P�G`�+��C�PpN9}=]/\��)�v�h����m�cQȩ� �%������S�N�g%CŎe;^����{��N�X*I8���Y=��D`B�U<�<�e>��].��1��J�E�ȫ�JkS�S+�X��H؝x��㙫`tw?f��)!ؙ�pCQ^��~.���'��n��7gペ0�.�s��Z���{����p�J�:zx{�q/ ���"�{���,��w�5�s/:V[lF�x�1���Q�E�V�H�8*���vh�V2H�?��	��
��*
�]��ǝ-�dr�$>�,d����c�:W�ے�9�/��;�l�mowIk!�鸨O�!l�'�&��FQᶏ��	���p���yͼ��8�qH��.H������/Z���9�B�]�1Iz��>��]��\�s�RdUT���v�9s��X#l���W9�reCE����/f����	��i�8��m/e�T��QV�W̔�`��O�+ųѕ(Fd�2���"�b;*��t�����ќ�)��k����̭���b���ْ�j&�@�b:�jOo��{���ߋ	yB8�tK�Q۷<*B3�ŷf��&�:|)���� ��\��s]v^���EŪ]��ʴ��)P�R�ځ�'a¿2Tc��dN�*'�x
�P�!L� �Iw�Zȉ�\��f�۷~;���L���:F+s#�6E�r��'�@b1Ҡ7�:��*�ׯ�o.ײ���Khs��=@�*)�\.�μN�r�c�����g̯\^1(�كݳ�wXۼ�F?���(B��%�3�� =�ޑ��]�=~O���3S��r�*�k����"�C��H��9�������"�Mb"�#!�푰R��*��ȓ����G9�,
�y Hމ.=��(�@l�b�:q�D);>�2���(�+���xԹ��d��]�s0^�$�Hg��]�y5I1�!pT��gu�N��$6�W��1h�E�~;zss|4������oUJpE*� y+��!ޣE�zd:�]�l�c��xt/�e
;�@tÜ�͔o��Ɯ6��%E�w0���
NL��r��
�}���������^M�	���
5^�!��V��0祬��d��*�u�sK{n
v�ǎ���T�o<�����F��Q�T��#X<�I�9۾=��FI`���\T�v�m#zfDK����Q�P��&J��q��z�ۅw���5�)U�P���)��*���~���6�F��q��U0�{]{
�]����y>����j۫�9�\�����&�>�*��'/��^��(u��}Cؐ�)so��h���/�:,�3�E�Y�ϫ���u���b�,�-����W^r��z��x��������U\�H��������l�gb����&*�KS�Qޜ0v���d��6��un+�p��t1�P��3��2�|�:���襀>�Ex;1s�~�,�eq�[����"�{�KMg�qܾ�϶(�ʅT�X"��;q��jyUt	�ډ��5��hl2���Y}B�ϕ-��M1tN�s˄�=�X������ͻ���I�ط�2�����T�+���S�һ�ٶ}����}�9�~y�������F:��cÕ���!{�2���`2@,�l9ʤ:�I!��=mޞ�n�)�{{jJ[��.嫵ZU�Y�y ��8�C�[�Ǥ���o>�-#����EĈ�"ሞ������C�ߍ{�/z���,O64^f1Bk�{�����Zw*�ܫ躑jG@�^�����b�\�Vq�3Ƹkw�|7���wfk+�3ЄJ�%��|�fGY�c6�I�Ӊ>��T@ٸW�G���"�-��'�Q�8�j�H�i@~�*S����*��}L�O��r��'&(R���G���#��q�V�$8�W�1��S��\�X6���C����[���pE��dH2���[f�Zr"ug&�x�`��b��r������\p��\5T�s~N��
C�8"C*�u+�;	os8�MnR�/�����\K+�?k���>g۪�]E�"=�������K�=�-��]p����5%�	���*��f�*���<vP���;�;��M�]:U�g���ЈT�=�_Y9U�
"��H��9�
���t2]�
����^Ș�0]e��C���#�|�5�b��"b�G��Tƾ��f�+fn���S2����r�Y�S{���!j��I}a%WLP���8u]�u�kPF5�z��o����/ �2�=���M�=�t�4�l��(��;������k�4QK�,��]����
	\z�:m�ڜ`�
_5�s7NG@�Jn
��&����䶨�fF;G�r8@�t���Wn<S*�gC�{"�xv%���B]b��r�����:�X���U;��$t[�0� �X�=�St9�u����\���{����Xb���1C����B�*EE�'�¿��"Ч
�ד:�F9���.��k�;�Ѧ��E*W*g�j�u�%�P8�d�4cR;��42Ol4�];K�n�+r����v������%l�����V��$��>��B��r���\��P��!��
�gݹ��˪ԥ/�6�B�;U9�����3�/&c�hb�	L@�09�/(.��u��V��D�h�#
���NKi��x�:=~�h�@���π��NI�ꭆs����g��a:�:T(#�aFZ��鸥#\�	�@V5��M�f��dB��	
�ŝ���]�_�/���|����a����}�F�+�k`�);�b��b؉,��d;��t}��ʡ���z)�,�J��Ô���G:�ˑ�K1:���Wސ�Q^�[�R?t^�i���[�XgZ��|^L�`�����zi�jh-�m��d��v`�ϓ��1�5+�mKU���.g-�wgGs��[��s+F�W�&ﵾXcꖒa�F��*8n3��7�'���C�.l�������;R1�%X��ݱ��WM֕���^�<�c�^�-�!Y���E� �E�Tғ�`��;Y9����u�B�2�l
�v��	��#D��+�ЧP��(��5��Q�z�|��3+�_3�V#��#�QN���7d�������v�8���T�jce�pM�^��(���~u��3�i��M�a�,��B��nXďC�ԫ X{\�xW���y��G
�9�,{��S>���\���F�?%cr���-�:�����Vk�9ɕջޙM���x(��{����C�j]B�HHan�fhV�Ŭ���g�!��B����U;�^��i�O�Q:�,����kG:iNz6:f��^��# �Snk��\O�����Q5X.g�y�%���+���9�,���d�`I2�R�SaH�U>�;U(1Y��b�J 3�v���������S�2'�^�E��v+�%F9�T2'y�WGBC�����eN�׸9Y�s{�8�{�kiU08���0n������g�h����Ͽ9��$��BH@���$ I?���$�$�	'�!$ I?�	!I�$�	'�!$ I?�H@��	!I��$�	'��$ I8BH@�RB��H@�XB����$����$��$�	'��$ I?�	!I�	!I��e5�Md��ou�!�?���}��������袊
T(�B��H���AE �J��IB����  R�TP�I$��D���ʉ%�R���D�TPŤJ�T�
�	U
$D������PI H��*�*�RIR��z�(p �V�P�,RQ�R����cIDS0b�̥	�	1������N wD��PmT�Y	�A��)i��A)(@ء�!!@)U@�u�1�m�6�Ul�I��H��� 4��w   @  e�  ���B%U�۲�.�@"��	���J�E�E2٩!hJ�5DF�*	�� ptk
F��D
���UY1%6�)ScT%5A"�AN  YC�"%-X���Fl 1�AkJ�B�kf� �l�U� �  �
S4�1�F��l�ٲ3e)���6�6
Ф�R�Km4["iM4��R�+c( �`(�*�2V��l
ՠh�QC	Ji�c0
-F�f��i iUD*�(p �hbP�BU��)�c j�ٕ%�f�fkZ�4h�K �P$��EI. �65#&�CRJSF�M[T��Y�ik2,- �Va�@L���(  &4i�)"�4  �   �x`�*�� h�224� C#&�挘� ���F	� ���T�# ɐ i��E Ba	�dOS&��{Q�z�=F	�iA&�C"�@�`#y5 ��4�f����I�r�i;��W��J�][�ZZ��0�(�*2=J
a��������@�� ��	���$|F����X���� ��QT�$����%
*�8�����V�m�Ö��D[R�S��~�Ɇ�lJ�9K���dH�#�8������z��T�".�]6�u*^�(h��ݐӫN�ի+�ԪDM`�V�����'�6�YB��7�𱉭��N'Z�����p��mެQ��۪KD��eS�uZ��a��G�4��:��q=��q�=I!��e�Ͱ����u�7�s(Ls���c��e^�B�IW�6�4��M�^*�u$����b�y�Nj�Z�H������ض,,��ؙ�NXx^��VӺr��-�@�^�fj��F0l�5����9eImMvѲԬ�ܧa��w�R�WGP�q^Q�/~�`�+^����FY�r��KA7��"/��*�7ڎjw�^������#xNq辫ǆ�QŒ"��ˠ�ՙ�ъ��)kC��'&�U������ӠN��;5:'q��Aa�{�BeQ�Dۈ�`ʹ[Qʲ���عs͂�#W���Շ-V�k(�9L��W��3SL�Ͷ3��`
���ݧ+EN�ki#���z�*�nhYy���ol�(ӳb�t��
8�YA$N��,�]n�\�����{)<tJ��м���G�$b�J�z���%T���2 [U�3x��h#�hYl����� <x{�P��$i����<,sN����Ѡ�.���C~{����1fn����bA�F��\-QXr�Û`��rm��,��٭������4�*�uJ|֥��m��[�vN��!��5`rimv��B�Vpa(��J��{:��sJ+�*Q�ĻZ̗gM,u�j�h(v�%���s\�r�:��g^.��d[ZhI4�Ju{Z5��R v2����#X���1��m�WL��jI�n��%��if�n��V��/u��+�ƓYz�֯(��M�y�4�V+�37V�jkJƨ��g\Yz�LȠ��"3u����C����P��Z�&���i��'�g���T]��sic:b���V��e�G*���Ej���kZՖ�4\7E*�u��طkR��e5�a�jC�{wN�V��$��H�S�V�I�9�f^Չ�Wݚ��0�D%��Q�G-'R�8�e�rA��\�	'�F��۹���Kה[8�WZfL�[PQ٢<W��mT3k4��([��͓kS85�������T*dPܥ�3fK��0^_h�Xz��X��I��3�M&�=u-�����.T���y�%�����P�c��ގ%�CC��=���ޜ��f�Zib8�̺F2� ���4�KH�PO!K�:�۾�rD�/���,N��:�l�N�\���d�ܼ�IH�ݻ:L�*���M5(KU�^�
��m�@�G3m���������Z43%�4ѕN�����q	w�Cc��-��ch�x)����ܷF�̈�Y�5̈^�k~�B�Ff��t�;�B!�)]���#n�{���������޲G6�X4���iDV�R���"x�����QT�x�Y����1`=;�X��6��� 5��t��%��h�ԫUt5���V���U�&Ui]Kn�%���r�&PW{�2bu��%�E�m6�Ұ�����n�Q��1���h�ͤ@����L�e�b�ǎ�C_enr�F�Zu��=�1��n��iA�6�)1.핺�ʊ@�P�O5�x��U��v��k��պ8)�2Ke=�0n�Dl�\͓hn��UA�&�e��v�i6S� >�]]�����m�RK1*�d�p�屢y�2\N|kA���
n���)�a������ �7W�$�W�uT���ݱ�n�	7��NGv����O)�n���ie�Q��+3,9v"Z�%��xC��۬m}=��r��F����6M���C0#cv�0�m�e�f�V�kyq'���zP�ƹ����i�m�[�|-+I��#%�\����%�����1��oFު�T��'���o*�QwOl�]�2��0��$/I�ArSۢ��K֢P�ڵ��,=�^�Q�e���o����b�
�9t�MS����4�k����F��x����w�,�V���5���5���jg̕)��`ؘU[t��vZ�ed]���+&&����s��йׯ0.�f2%�\���h�����a��;��R�ؘ��r�Bwx�k�T�Z,ST�G������L���3�ܠ�Yn�j4!̥�2�]�ܕ�V\x�M-���?��R*�������rl��>�n�d�b,�c��Z�(l��;�u��ͽ�1:Q���&��Kf���ַo�����q�\��:
��(��l�gnwnf�0�j�6�W������L$J@��ثi�I�8r!z��lP�Ut�Cb5�xh���"�ްm��.����` �{>6�yr�s�7T�O���)劔�}�@�ނ������c(YӴBܨ�9�	�2�a�6�gk���f�wP�oq먓[,�w�hY*�b�C���l���b�&�1�a�Z�F;Eû�8�6*Vl����9H:�okK�Vܬ8�k<�/6��C���>+,ͭ�/Q�X�mԆ�-���f�*[	4�Xl��C��k/�ͫVUE�f���U�(�櫨\L�Z�m��pN�go+uA�<��ZY�޻z����������r�$]��RL_Q��]f`0�kS�uwJi�*�6��ѕ_Ȥ-�{R?��p&�]��%�uRՇQ�UL)5+�n�b�f�Ƹ7���<
|��W�)fb��nR|�����9���y�7Þk� �M�c/5����J�B�d�W)AHL+	���M�+�n(3(ňP����?��_X�x�>�I�M"*֋4�o�Ӥ�������WHs�1��V�tΨ����?\6�(*1J6��o=Ig-�UyZ�e$���H��X`��&��zE3��)V�v���d�H��H9�\�'2cN�1��ט�f��n�#�E�H��eeA�Ox�
߮+"^QӁ%[�+Q��,�P(+K	���A�x�=e6���e޴��G>��,̽��wQ^0ʼң�{r�iֺͫ�uf��I�j$h�w����.�C����NeMld�QouU*X�L2j+[�wY�IFe�H��e�ћ7U٬���t6�)��I�\�f���£Ǎ�9�z��6��-��
�8�HCl`l?��'ƖC�f��i�KT�;[gF6+��-;E��T��Ռ�*�Ϲ�-q��.$૥zt���ZŚ1�e��B�\uj���+.Xd:�2�N�z���(f���2��r��z-㿴mjږ�`��Z+0�����hi��Q��]t,��8z��p%������/�+,����t0Z��eɔ�訝%����,��̙��R�M�;3~�U.�V]�7r9j���v�R6Ҡ��� �9�oOvn�e�e�Eb:��~�d�1�ݍ���`+v�)��g���XN��QQ+ڒѷG���e���#e��$��²<Ya�MI,�2m�՛�3�Ė�Hsv�,�G�7YL�W�j�q����ì�T�ٲ`KRݵWWT	oP�G/+t�Av�f6��,m�z��m��	|k��]����ux8�j���Sb�m$��4R��Dڤܗ%Cf&���51��2�[��Z�q�
as����?��n�+	���Q@�Lu�u�:����'��A𣯺���fΡ���V�Z$�t�b[��[T����i�K��>&���_wcg�����&����^�u_=!� i����+��[B�v�	UN��7��]�a��t�0VȪ�Wj`lS�rUV�'-16�]�X���"�5�7Z7,=�L�������R"[�K��o�ЪuL����Z&\��#w��a5�E�_E�
&f�%�1:����ֶ��s4Z܍�hG@�;u�ާG-cL�~����#�A;�|L��H�����ءCt�������P�[�vmZW4M���0�5�r��	�)P2[���M.�ȥ�;8s� �A���E��<�p�e�.Nos�u,��t�b����eo�S ��:[[���6wp�Zz����0������I���ddUxB���\K��Fa�#�Rrot�����g{��&�s�>t1�1L]��fwM8r6����ro8x�|�T��Yif���!�+sUଊ}wl���`[7.��R$�r}Z��b�7¢!�#R�pu�e�09^PG�����@"wF��yo�[�xm��sv5w���u�9t�_'���Y3-Xu�f���(n��:�/�v�M�-�I� �)�p��f����K��!\�7���m޵xyĳ�-Vjv���/EG�tP���#'�9'6��������5�7ݭF��u�uJ��dtU��h�$��u�`"�����O;ZlX�/v��*�ɓXb�:g�U���M*��s\��Aa�;@���� �:�cf��0}��7T�;oNo C�h�h�˭�:���A�_<&�q�qYzV'�QG���w[�L���}�a��1ϰ���{�`��K�����Kݽ C��f�C��>k	��-QθM�񿱄ʷ�����mZj�\(Wv\�ٴ0e�v�(��Y�h���!p��U��<�D$7٣�!=�R�an۫C���|W{DV��y�w�����m㫫PK"�S�t�����L�[R�AS�c��h]m�q�.� ��Α����n�����2Q�{$�ut�)(Lig���q�Ne�\_��<Y�����+B�U��4k�l��[�ڷuE��}J<u���"��U+�|�F�'tzn���^�n�|A���53(��	3�)������U�m�vst�
u���,z(\fd�fQ��;��o7���*�I��ܽ҃䣪���<�5p_%�\���IJM������ �:�]�ՋN�V7����v�&�<��i��b�Ba�D7�;�����/Q�.Ѿ��5�A;Y;En-�WL�I��֐39�AykkX:`}d͊s��a��Uٚ��끡���	�Ζ�xCv�nm�X�'�]�����(��MmCR�QU�3
]Fh<]6q�ʳ�z[}xʔM.�%�'���]`.����0�ٽ|�t�'1,��u���Na�;H�"�r�ohvX9ϭ��ԁ=]y��!v��Gf�M�'҆۫�fX��I1M�����J윶M���J�l�$�aZ"��W�w��{}ٗ���N<����@�aRN�̭$ܳ}��'y�A�%��VdO"��9���V̴��ѨJr�u�[!5�M������W&��T�vN��5�˲�y@:݂�� �gWeQc��xM��jC2��pL̰���rv��n��]ueF�5�l".���YnJ%E��|�R��PŖ��+���S�G��-�r��\�ۡ�J��q*�Г�x2�D�
F+v�G��&X�y��EuJ�Z�g1"{ˮ7I	bN�0;X���(<W�0���@��,_*ޜ��5�6�ZKS�ۈ�0]jXj�tv>���v쉜&��ށ���U��.-��N�e����L��1�Z�,�)fr���;Me_V��o�;U��#�UʙP�A��z��R�`�w}�)�p�\r�
��˾Z��|�=|Q��[��Ӯ�Fbw�'\ѕ-7���KJXSyu�+HTNM˙ءu�"�P��2ƣeE�� ���u���[�'t��v;�I�l�e`�w�r�η,9��P̳�5gc-`��w����2�1
�u��D-�t9�+�2�r�h+d�[���?�Y�i����s7!{m�EgRݧ�-��j��ó�	J����:�:�BA��c��Y�1���̢�f��/p��ՠ4�ɥ�l���i�����~\��ڄ�-�t��ത��{���P�j_jT�pڃ��C�*p;��'�u�c�FoOyJ�.�e){�cE�������^N30Q�CF���>A�5P�.�{�o�dS���ۻ��;#^��ֶ=zeҖ���{��w��pX9v�m��x�;�O�;��D�S�l��j�0v��K�O�#��*�.7�Wl�Nv�vE��o2��:�W#S����%��gy�p�{��*�n�9|�r���"W�-�uŖiX�wrp��<���X
�)��/U�ӴfL��^Ң�,ٚ)A�F/���U;��f�h[�q5V�t;��N܆�5U���T�`�w@�/��u"��ѫ��:.��1�y��ѱF����K�G+e�7
a�c�Mɪ���r�Pphǫ6�R-�k���[�gv��x�+7p�&L4fl}�+H�"
"�v�(��n��(upb�Wc��2�}�}�Ν�C8�f�w�uȍ�׺�q����'���AJ�-S��
Һ7�M��q��֞��7aA��'��x�X&�Z*=�D�42�J[3�<�P�a�%���<܏_9���dX�6'm���z��fgZ����|a��}U���$*��y���	��U3ܦ]���Nk1i�WL����U�'HE1�5����N�_v�¾��RZ,�5�/��^�8;���c���ncܳb�p�U�1�{�)���4
4j.f}��;��>���ϵ�w �1Q��ef`H��o��Q���u��,!���ss����\W춳c��=��l0f��F�"!z��Vd,K4��n�]��[G]�ee����]�:�h����)UL\Hڪ�,KQ����޷�:{�7Q�>���]��d�I�.���i��;�V�Dm��Y@
����E(t����%r�v^���&��\9�Z�f7�в2�8��B��򲋱0WN7C�c%�b�uL�ctS#�J���uPUwr+�q4j�x0xB�NFmd6�"�\���㓛w����c]�j�=/��	��)���"P�C-���P����!MK:!������2`ү%eV�W�2�����oi�6-�Ɩ*:c�����Zˬ*��C�Tz�QC�I���d����w��0Ń0uj�6f��L�=g��籛��{ÁV�I�JR�`Ƿ�vl^�>x"|�H/���6��p=gT�w��p�\Mاj�itЋ�t��O�D-O�ݘ���+��®����_cV^�1v����G�	��R��(ѻg�ٛ4Vc��szru��8�Nط�)b�u��"fY��Rqm:�#���z����Bq2���x�
S�0H�G^!ս4K���C�L�|�̈ri��WLo�w$���Qk�FB�����i�&�@�n��gQ[bI2V.�a�g:뛈�F��`(_v��㬹�x�� ���ъ���E��RI�tf'�9��Mʧײ�wnH;Re�u��ܒ5���&��8�w������c�3�x�<�O1��јHUڔ%��ʛٰ���Y�a��0��b}�r�@"��	��j�[�+[��9�5=d�`�X�r�F�c����V|1��)� 7�H�AK[�ybsrrܜ�w9j�m\(tFlv��[RI�I$rI'pI�m�M�����H�YgUͼ����Q�rf$�Qbt�w]sD6�x�˝l�+�U:]�j񋼷4�	��R�Df��4c��×IѽvsNqj�dS�X��k�@E�8��:�
�;��J�����E7�!-�ڛ�@��K&��� u��;|Vf�ዯfmințu�Q�4��U˫�Ba[��;�؊[�$��*�ve��=dY�K7�*���uj�޼�t�{�2A��8�8{ �Rwv�2���LA�k����{y=��%�c,�k�T6K�����sx�a}0���[R��|�S;�s�X��<���{�=I��V�3�T�p�w�b��\]�z�e}4�eV�����E׎~���,�p�Yu)ӄI2VM�.�<�fS����x�8l��L�p��[�;)}�6�]f��.�R��O�����oW0�N�v2_h����1�����eD�az��[���J��Oö��e�f@��r�c�/����s4q�\Y(ۥ|�Qg��8W,V:u�`�1X�oe�� �ox���Q�+���P�,mH���o�G/a���\xv�*�WN��k,g�,n�%�]"[#�*���t�
.���l���Z~�P���/t��vVρ�3�"A������ؕ7o ��-	6s�wm�e<��~�+����h2/���{�ǁn��\ŉ�غv�i΃�� �]�8f��V���% rm
�CӸI���03��]Q�r��W��W��OX�F�fa��I�7n���]�Gޱ���d�O>ƍ�y8��r�F���Y�6=����J�2ۉ����z�Ȕyˎ��kY�e-��K$:�tu%"X�`�kyEߔ���ɘ��1���l�6�����wP�X��A����6�^ۆ�Pv���V�0��Pk�mu��U��$����m;�t;-M�L6��v��pۙҖ#�Ӆ�(�O��WG+�9P��5v�2\F�OT
�)IGpEԖi9�Lf'Zr�gh����\�f���2���]�`�ʜ��s����(�Ćm]pȆ��&�Ҳ�J'}�`P`�Kt�/��8���W�K:2^wV1�Ҋ��f��-�#x�l��#tٽukN%\�ق��xM��Ԥ�;b�\>��mL�y�Wu���ޚ�9�X�F�3��à8�� hE����}4� s.�+0��]���{���� ��˼����ơ�!�<8Z��u��q����U��
�|4Gn��Y��(�Gh0��-Vm�߭��G�<	�'A6<�r�����ֺ����h�ŉu�W��Z�}�-��e-�vԔ�>(��0�09sk��;��� �ژ�u����U��c��4�n�^(+��*i|��1ui����n�b[�-�;�������J-ɷZb�5�/;F����<Fm�6��Z�q��A�T�xX�(!�18�q<#h%]�8F�]�fp�{g%�T�N�Ӛk9��3�a�0dλ�b�+t(��p��E�ǹז2��-�4��	`�vPp�\4��#@*�O��Ŏc/t.뫮fɹ%1�LS1�U����U�u>�k�v�_�]�-�[�d��a趥[��[��-ʇ��Bڡo�0�b84JMKw�^�y�n���J�I!-����;����BJ6��Hҗ��ڄ�B�v��c��Hu�h�̚��S�w2T۴����%�����yYmoD�RT�C!T
k�N��Ⱥy��S���g���%��7���k:���7�˨�o�gn�;�_,���7�mh����(^�}n�3Xj��|�q��Y��2���K��Y��a��r���T��x����V����\Ah�C��R=�ѷ��xS�7^���dӞ�5�C�%M �l�zkn����Ԭ�w�_R��NҼ���dV"�]`�up-[�n���X�nP�'�Y�+�Ȣ�-�EQ������s���P����[��d�Ϭ=�E�{|�`���Vc�6٭6�Jc��A`湷>�U�c�1�ܭ�zV�����k��ZA�Z�TY��X�X��,��3�M#DHS}�O.����l��ؙ�`���-iNu�<b��3,l�X3�8�5d�:�#{�Y��i�N$�Ԝ9&��˺����O��+�
��Ik�[,^�ct�g�3�s�tAD��>�r����=����g�va��2�Ŗ�u"ſ��݆� �M6��&��:�V���0��Ӻ�pw�W����N����[MT��bd�ruT���0ChڽР �ݨ�͡eu:�Mn!��y�Ey-f#�h�K��s]��� ��;6����%��iV뛼	R�$��>gY�n�]3��&nU���X�wdv$����yit�l���P(蠺`$��e�Ic]�)ثk�1�.֩�����y�.,��]z���)$�z���{��.ۺCi�%�!�MK�щ��V���3�X�[8YZ�e�����Qk�t%��k�f>_f��	�w`�5$9K�m�!�*�)�mPYw�]�#ʱ(�)YM�&q/�hE��G)���/HLs�]��ʭn��K�R�����N�s��UyF@��?�#�b����Nf��nv�r٫T�5no^𙯡�7+������WA*�����@۬�M�[,�Y�tUٹ��W_q5k��ė5Iwp9�V�7��wuo}���u",�՘h$�px�Z��qoK����p#qu\3*��U��GS��hL\[Ա-�Q�\Z�\�F�@�a\�+�˫�6/�W�ǒ}.�xo>�}ܷlHØR�n����@�4rGD! cFS�
��W���\�rT/(��R�Bӝ��)�ۓYD���6P��n�;Rż*��}�ۥi�5�
��A�{/E��}֎��g[�f�^dI4�n�5��8Q,Ʈ�{u-���Hٖ�`��R4�J6����{V��S��P'5b�Ķ�ۣ��p蕡�t��Y��3X�g���Ty��8[�H&I|�K噋J�3�5��n�x)ɣ��%wlh��Us�qU.�vI�}UH�w}5n�R3z�s7�WE�I�_mi�Ꜽ�RuG`�CΪ��GmNCEgK�Mo���ړ[S�"������K]��z�`�&3'l��>���PK��\y�Qa-Q]��^���uΑɆn�Wk2��K�ܫ�gȵ���`�4�u�&�*^�O5p�;iw3cOR��b���Y#�'f�v���p�<���2�{�N�h�/A��}���4�O�p��=`=����e]��{�խC�e�Z��a[㢄��r�f"!f]��ϋ��hJV����u�N�N��I/ �wx���ԇa���p�X��\��\��┣9�+1����l�����7���Ý2�w%��@�n�]�u�@n�:�t	f�����2���p����:\�WD��h.e���'��*���K�ciE�b����;(�ҹ�Ԭ�n�[�ni}�P���y����QF�0�+���0���3|-'p�Y��휄����	9�]m��A�p��tޭR���8槌�W7�$Ō�;1��G��t^0l;�r�[��CXA���1D0k�f�������	bNı𽼗�V�ݺՎ<�T��o�zOs��2�%�p��1��8nV��vp��bj,���� ����(��,��ŷ����t���(��f���6����o�=J��;���C�S
�f��"5�R��|�'}�u1wQ����Ȭ��sl7b٥�mJ*��	�u`�D�4���d\�s�����X���s,�pT�r�U�l�ߞ&�����֚�Z��G��"���}���h�&�;����>��ɕֶl��'�Zd�����a��k7�j���A�SjAmmM��%��FPزᳵ|6�lV��h�$�3�f��Ft�2땨�7R-���3L�҃#����C�zF�1<��|��Nt�l^p��4PxݦѻtAН�I�����;v����W-�6`3�]
uo���1#�cOC��ը5�6͛���v���mdX��*�j�QL��Z����P�D{O�ƍ��k�
�#���VZ�Q6�:�+5�cr�`�paZ��vu�Ң�m�b����כ��ҟ �b˴.�k��fUu���	���^�4�$!�Zy��Uԋ<h�ݹ%X��HR!�e[��8^�6Cu{s��痽��e:��o}��7Ӵ���@ *E4�H{{�}倉����}���yߦ��>
vʎ�YBua��ef�k@Sk[]�����˷2̤�-N�c�Ǖ��ۮ�n�w��ލ#i�b9�F�r������[3m�9U�ytrԐ�2:��L�BҘ���SG��GJ�wR$����b�\����A�E\�c*����4�Lwo%cb�Is�n�<�t�Ir񪼬ĺ2"�f���W,Pl@�ǚ���.�lW�h;�3��T����;w�N�l�:Gg����(J�1��݅'5QA,Kr��+V�VV�ط!�r�ܣ܊�Y���%bL-��vVʫ�{�'2���JSb�"Gm��ذaΈ�ɥ^ٕ�+ޕðX�5{��kb�XD��I�й������	9s6&�L��;�O3)	k_d��dG�e�;
Ѯ-k_,�N��A�+kIۂո����̢(��n0�[�����)����X�wnV)V�f�ckִ�D����DՋ���SLE2ى�Ŷ�jL\����[��d��D�hc�m1:u�]!K�PS���#-��H��0C�]9m�J�k*"6��.U�mJ��z�&.�*#���m�m-��R�fDq�mEffb�auu�bى���2��Z\���Z���0�2DC�l��-0j8�bT��Ln�i`�j���NC���F��s�]��8sLɸ�ybDŸ�Ï�ޅA&��̄�H�nmU'�����?����s��^2� .\G���3�޷�v�܀\j�ON�~�w�yg�P��C��`$l�n_�z�P[K��K��r��g5m��՗��A]' ׈����!=��-��ۅ/�CF(�jkWN��zZ
���&��9�!��sUg*�w��Ο�q�>D��G��	K|�Qz�S�*�ô5�����M�o��M!�� �a��̷_�����~��2���B9�u�4�k95���=< �Ӟ�E�t����W@�l�=���ܥ�pF�G�A!2v�§��tw�u�{={�w�t�v>IJ9���8��fnޜ�}�5(�4�F`P�Vl�2yfb��*����v`gr�HL�٧gˢp�	��!����哼󪱾��;}\(DkU;��][�xWvk�mq�����Mw��:D�'�&�����j\����9[R���۩�8��ooI�}pM-@��f-�[&%
.��� ������F�e5db�Yt3{Q��}�;C5�C�Q��
���}� �<�V� ���'w
(�uV_���{�3�Cs^f�{��Ī�v��Q+��`�N�<�zkFr�]hp_-ݲ�y��j�e�i*���FEf��[��7��Wn�x!ڪ�#������@��Ӗ��d�G%�!���~���n4Ў���u��DJ����E��}�\3Q�."GO-F%ToEC��n�EĦ~xXP�k9鴏<��o�W���T�ՏN��qm�%D�m^��Ѧs���bw^�j��'UF�ck�Ѧ��L/�޺�������}�W^���\����)��5�g�ּ����gZ��#x ��\���B9+�O��<}pȲ�A~�C٣�<�fQg�n��<
,�;}]O��g_��s�����p��zU�C��C����a�Z<��¯lN&�ТMP�D?StS���S�5���ִ��er�MCA�cc�Ъ�:�+��y�I�cmʎr��ϙU����1P:��A�1��˘뷉�X�+�Z�2{F�u��b��ݬ�m����YZ�]\���8�����Mm�k3r�M��� �B�$�f�H��t��w���4���ͻ��������{�6߶���z3u��2x\��+}gs�z�.9߁��Sb��Le,�zh���\�xk6`ح.�;7�L�aol���wꋸ�.QY�x&W�e����4p��Z}`C�����]9ڡ{mccw��b;$��2[�_1bwF˫Ӽ7�963u���C��äӼ��]qU����qD��$I��n�zW�B�1�f��z&i��<',<sN�x��[ʰ��3g5~o�u>z�}�K��AӁiq������]�G(le�
b�N(~8 	s͵���/��H ��bõ�I��s;�h���;x�+��7Q�j��p|��S'��+��~%�qEne���|ߒ�J�K9�*�$F:b�Q�'+�Q�\�� �k�V�l�Ǥ��i����5|�#��8S5��s�1p1�:�ͯU���{tk|ɡ1j9�!C�t�&�l�|�$f���LJ[ʚ`�ܧ;ݝ�NlG�s�Y���R���
1ǮG�7�𬘚ڏQ����v��^qlj�N m\jDD�W��"���fg��|��?mzmw������0^ֲ�i��%�=�W�tz�lK���׶�y�3W�VUVkz�5��`Y�����C�������o�K�|��w<�aVYzk�E���.͆�(���-�il��Id��嵔�e�<��ب��i�����SJ-J/8���%+k��v��^��O���=ub�|ћ��&���wH̺�z�]hu�t�/֬Jvy)o(<3���XӲ*���������n͚Tp��A8J��p��Y\�w��Pd��%w
�����}��-3��Gx����(&S�������G��6n(�[��e,%�±k����OX;|j2bʔ&G'f�3
V߶��6�ob/kϪ�B��=�n\?e�2����T-=��sZxcݜ���Aj�q����b�}g<VÈ����D�mK�HK�y3k� �z,\�msˬ8�f���54MC�;�F��57�өz���ݖ&�X[u����gF�V�sU�Xvm�g8]V��B���7G��%O���C�L�?�~�1�'[L��>ⓆDS��r&Y�G�D��/^PY��'k����H[/���;��>�n�z8���r(͂����2mf�u��&��}Y�W��[����LI�[�,X��/4J��:,�<.��8��z��C$��;�R�홸3\�lh���Y�]��b�B2�nb�Ϳg���c��&�c��hVӡX�p¾�*r��xUsѽ��r���P���iUC�\�4��muߵ�i�դ�~܅�r���]��#�F�F�Ql��̀x.�����8^���
�O���%A�țs�ߺ�f⇁Ռ,�s ��G�Yb
e�-&��s�놿Iib�?yZKѐ�r�3`�}a��v�z�9߁��['�c�0���)�����z;r�p��hE�^S�yS0��Vq`�"��k8vLN�pr#�'���3Ǖ���Z��p�p��վ�ؚ��-S]�l��ō��{���߹A�a�\��6��eG�X1OyF����^m�k��yɾ���9���P=M1��*��ۦ5w�ަ�PR+wM��.����|��qo٣y�BVU=vn��n۫�!83�t:�W����0�¢�_7s�<Zy�wv��X����~^�9$X��U��2Fn�4u	���d�/3Z��h+5�ݏ�����]$���{�ժ���,o��S[�eȄcK�O-����|N'u�,H���<VJ��>f�}fo�uE�v#Lָ��Wm��a��^��;�ɹ���+�Y�C��CPܸw��S���Y��L�*����ET5�x�^�4o��P��g���[�n�L&z���5�μ���i�ո~����Fw׋�6��ʍ$��w�O�ϊ�8�]m�ާ���kr�;G�ٽf_*�G;����?t~�گ�}��J��V�ۗyw9LR
��kT[ Bh?��ybdK��K�6���SOU��g3%��iݔ�fGL�xݔJVzʤA��u �1��ic�k69Ew.mL�\2�V���&e�&�;� �Z��Ktؠ���c<j�h�-Ю�k�ܩ�Rzr�
��{*U��G���������@���˹h�c
���HU���o1׬��8y�E�T�4��6w��M޵vfZ�R�r\X�-�Z�][�����,ޘ���A{�w���q�@`�*��f����mV۫_-��Dmjq4gU^=����C�,�:��3��4�Wpхe�xR7!�k���_u����0��ܳ"Quɝo'vr|��6M���y��)|qۼ�d*=tc�ݫ�`=�hȶj����v�jk�*2�gX��䡔�l]q�Q����U�d6�s����S�c&~k�ZfgTz���%pt�D�j�|^��B˖�����dk�����1K�5�ʩa��A�c�w��]�Z;8����l���݄錶x��ѽeÒ��"VF�w(�2Z�V�9��1�Y�>޵�J��U�混�ԯ+��S8�Eҡ�Փ>�:�tf��h]�:��tk�S�!r�ھ*YQ����EZ�k�\S�����'J���޳�f�ֵ;���u�f	Z쁷�0u��zx+a4ާ�W-n���h^v�&Ӿ7��t"vF�Ğ��l�V�՝��*+�$��r�O�n��T�)vT|lQ|v]���|��NǬ9��|9�sU���q�Oj�epX@2"�.8X�TQ���x�� [�vuouV(��OX9��\�%<X�.��S;����_���� �H�S.�0.Ys	s0�V-�bţ�q���b���A)L���b�*(���Z1pU�˃���P[�b�
� ��b��TQF(���*���X�ƱT��+V[UAUk�Qb**��QDQ��b�����j�8�"�ت��:h��b�TV"� ��ic������o�/s>�����2# J�Ml���l�0f���&�5��K��$�^�s����-��4ν뽒�Q�5Kq���U���fZ��7�e7���R���ruJ�<���{����,��Fn������!��nnߺ�7�\[%n�ť637[��,�!Z�����hє�
OWb�ei�eX��Dj�.gZSV�OCs�9�ξT㝱���t�^�-��P����A=~x�-̇tq�	�!����n����Ѱ0ؾb����A�G.gT-�Y�W�X��c7��5P
�bVU���Pm��:PY�8S�8�*�B�ޯY��߫��/��F�&�:X9�!S1��3l�0��\���r@�3�Ŝ��������:f7�_�nXƠ�7���IXf�oj��bz�����q&�����o6�_jGu�|ٚ��Q��Ӷ�72*c,�	��i%�������N	Q�6�� �%Ȭa.����wή�'Ⱦ�V�7�ܰ�q���N瀞�uy���F��O�^�/:�&�D�2/��8���%֊'��N��B�K2P�t�{R�^��:UAyoZ�������Z�����W^����C��J����_f����W4�oG�j����d���Em{·A��Ի��تn�df��.0�q3q���2~���
���>�8+�7��wFh�E/q�����(��R�y~׷�6�0J���w[��e��V	w��Ol��Vc)���:��<�t6
�,��}}��m����z�㝂z�
58�3W^Ɯ��f穢�#WI���Ð4���ة����?^�[�8�z��=
3?������������0=a��S�	�ۺ��6&�V�"��dj��bFHl؞�ƷaD�[1a�ً�ɛm߻ICT��,���镽��/��vG�GA�'��S�V��P��Bo8t�����@�"Rxz�A�m���V����[BHg�~u���{��{G��7���PD��^ �m5{��z4`�7��^6��2������]��W��u�Cs�*��
��ìx�VC�j2�-��h�p�e����}C2�
�='�=��ז�ױ��
�8b�/3^T1^1X��Ԗ]Yƛ�ɒ���հɸ��Ψp�N�\Re�m�q���!uY�x�"�n�<\�{���d�{R"z*~ϟa���t�Z������۲�;����p��nŗt�o�k��h𭠬�9���O�\�Q�;w���;vI!Sƪ[���+�:ă5��E�%��S���c�k˔u�E�9��|P,���:ef��_xyT��x�7�=�	g|=W�0V�V��rU�v�egJ�T����GOh��}�P~"6W��o�;�mVga}�{1��5��x����=�\.D5drW'��97�f�вz�^gdb���B�V+��w�e�SBe`��}��g���4�/&�-0�Cq[Y�b��$tU���u���G:�7���L�#W��.��
s;=���6�T?9�v������XR�;j���;�<�˼g�y�Ũ�w���S�+'A�U����Sz��n^�H�q��rG�ʶ����\s��ب͡O�18-)Ula]a��67���sYI�s;�O�"�@x=�{{%����F� ��as�N�R�fj�]C�z��o:^���S�c"�v�߬��;����o��4w���䱎z>=�l9,��C�QC�d�=-�B;W(#� �kgL��(��H}B^}�YA;Գ�Q�=�(�<J�]X�[v�1�#z��s�1Qz�c:�M;�4:�ϗA�.T��e��<�4���_j:v$NpktR�j�Xd���r�b�G-y|N�Ȗ�*��ub6�:�.�>����%�ݑ���<��Sɲ߻�F|PL��;�K��o��A�������\v���(�3ظ��Ӳ`�^����>�x����v+1�T#��j��g�)���;�<�r����~i��p���*�sȋ�^H�����$�>��~t>�y�]��v{J�ӵ���#����U�3��`����u����wv�"�n�Q�7��t�.�`���&_^_k(�-8��$nz*(#R�w�<�9}CQ�{ճx����Dkuz��V�	Y��ս�}�(LHC���h�0`.���wΖr�A�̑�"�"�̹����oy������jڻ��?w���OR:�2��	�u����Q�S���	�y����1n��=1!��n�Y̜�x��4�J�݆�W�cur:U�H��<��O�/ǧo��>��Q	��d�*{��羈ܗ�;�8I��:��̺#��]M��XosZ��d�)`X���M\Mo���T��S��>d������}@a;�����޺>�Y\�1\�2|M���8��_���ZȎ��tMv�7���'����kω�2���Vn�����a,:#�Յ.�=+��!�&U���*r����w���n"�}R��V�Qɭ��~�/�W!;�*����!����-�9��8�m��6�ٸ ��u�O��8���_�����2Η<)�U�I%�~�8�H���T�sЅ������61���e��oc;8K��
Kl�#{K�6�]Ε�v���"lcq.��=���L\(��|��݉ۢ3�\��L�<��nom_�����&m��c_���Y���)z�5�I��;:`�⼄D������9�n��y��#��v���@hzY����B�N�/��x&*t7�7jG���D5�\!����[���{�E�=�En�֤�Ha;/"�9ꠡ���p�Zr������+��Z�	�������ڊ�S���w��k�!�����t�|��n��S_�,��zͼ����<֢�r��] m{�A�x��%�op%lv�y�����~�J�"��v���sg�Sx��d;�����dnu���tv���e�T8S%߶��|�EE���X����-�د^V��ш!�y�i�%�c����o�r��5������ε;�����[�V:(�{�o�m�D��}1���ڌ�ȥp�õ�ζ��'˫.rvj-U#���-�n��o�i=���0R�2�ɟRD�BmEÍ.
E��ۃKV2�v*�\ʽf�æ- 0BE�:v#b��}m�r�Քj�9+��\�vk��Vhܺ�"�� ��k��Dvg��x�n��H=?j�(.a=�S㽧�:�b��#�B���ծ����.z�a7^S��b��hʘ-����Y�VR�J�i��|�F�&��#C�6v��CTn���ԅ�� �Β�x39r�$O�4^{�F�}ҴF�
���k�ۢ��H,����$BiV�ó65����	��
�*��(�GP�ac5�����*�~pɛu/JM4�q��XR��uc}]@�s��D�V�Y`M*�	�i�yyK�	Fds��g7
��6o�wVr�0��
�c�?Zu�.9��@�fOI�����5���s�4�ɒ��`V'\���1p�_n�6�u/��*G��6��2�WL��A��p��y�гq=��V__s�v��cպy�2L�L�B�ת���N4�t�����,�.��7�ږ~��D��w�n��v�L�#!�>��޼��(rr�*i���N�[����$����AC�3Y�.e}�� �WܫJ�z���UZ��Q�t%,�[���W�����Ѝ��<ET�r���W���lcú�2����pȦ�N��@hl��@���r�O���#�ü�5��^I)]{H��rb��n7Jfd�t��kW�]n�O��9� �+!8�p7 btW#/6�a�@�Jb";e���XnS������PY�||��<���G�AmUUdT���*UjX�J�҉V�X�"��"֢T�J���6ʫ-
�)*5*T���DJՕ�*���k(�F"�b��D��1��EDDdTUDPEc��1��T`����Q��TP�X�Ĭ�3F
*�(1X�1TE�����E���&"*,b�b�-J������ߚދ�E��~y��½�VoWa��(��8Hu9c�EȤIg.Z�d|�3��x�T*G��U��1��|�I�<Or��	yQ�N�cؚ(��)��<��3]����I����;�`H89z����W��XU��Mp�C�z����1AUs�ux��T��!�/�^�~�Q�z�Ph��^������+�z�,M�#���gmm1���v0%ai*Qn�䶟�H������]`ݣ��uc�%O�����<���yy���0m�:�i��Պ�3h��/�8Sˮ�w�����=���Y����7\^@z���F��\5$%;:����o\�*.H��=��ܬƜܚ�a�dq��wf�r��$���'y���yX���'���j��L.1t�>f�e��v���w˭��1��_j�;�f�L�}gs� U8SYk.�i�#r-�Iz7=�BR�Ws��I}m����/��s��ӄ���g�s�1�E㌰��/({<�(�{v'�<�L��O�W��Y��6�i�[K���Kn���]����P�ʚF�o/o��zn=�jx�:�x}�X�����b�pBQsu��[�;.W�h٪h��Nt8����יwWљ��&�bf寡�9{��ml*�\)�b-�����id��\n�@���[Fz�G�:��뀎V�iU�&�"֤�4�J�y��T�#
��pH)��8����Z$*��N�-�`^f�׵I:�_��ó�p�[���[�5ei� �7�f��9�&ׄ(������:$�a�t[8�cs��(���Q�ͨ�v�;ʆ:�%�^jx#9_����~�YFQ�Á�zy�PtV�M��qѭmcgʃ�<���^;��-��Y� B�q��(�ޘ����k�����z��ͣ�μ*o	ۢD�n��Q�'�ӕ�H,���.iԩs:��Gf��㼥�e��m/;]#7���g��7��XA�
u3,�7F>j��ݓp�"B�*�t�Xu��R���Eq�$��<��JD����@ʙIqk�<����D5��S�!��ʘ�[D)3�{����F��[ˠ�oz��V��s�c��`yo���Vj�F���ō���y�~�¬�d&:#����u5<�=��G�ӗ/.���#n�m�I�~�A�E�¡^���c;���
l�
��u�PF�U���Vf_����{�FM�lK��k��te��8��ԫxB"g8�՘�6
y��z�̋�
(����Yl*ȴb�9Š�)N�|�u�1�]��ݻqԟ�zv��)�S5A,m���+��xR���b2-*�rƧOu�ң��i����3���'���c��X�����O1�1h��7❞�^��Hu(H˯P��糪��[|�K]I�Q��������1�U�k{�T �'M�F9���^��L�����YMT�Șbhi��p�t�PLue���S��}���� ֹ�">�����s������,o_��owHYN�(��%q�<�2B`�j���x\��I�A���B�O:�>��{�z吏:��mf�/5�f�kU�//�|VxZ���zW�Ocsā�9e�ǫ�N��oe製D�5Ҳ3BX���Ю�{M%AuVx�n���p�h�ӽP��ө.��G��|�ݏ�c����O'��J�7q3�;[��-�<��$A��]��N�jCD�/���ܼk�rVY�N�e��i|�|�f(,���Oh\�.$aSu�wB数x�m��G�ё]QG.*�tƂ�'$7�/s�������T��#=�cExɚ�ON�2z���[N�XC�zn�e���D�˺bx��m���KH��`�i�C&Wq�ㄊ�"��w{�An����	E<��wm��ڈ�o:V������������b��q�a�&]��7.W�4ޑ��
RUta�Lf���g[��1�2�yp���h��&�Y0-�*î���k���I%#����z"%��kc�'㈲=Zt
�[S�7s%�G�=������s<��	�q�2$Hm:��m��o\��=�Ϸ�$�Ʃ�HM}N2,&P=@��5����'T�� ��o�I&!�@�z�:�r���9�s�8��ā�ug���4n��w`z��&�l��m�l%H}톓hM�9�:I*O���O:����zH,8���6�i	ċf���OO�|�y� ��M�!:Hk~䞲����owϾ�>ߝ�C�x��wa'�����E���@��8�:�|�$�$��l6���4��Ntv�}���}�O�C�3�C�XN���M0�w��C��2��C'T��8ä�w�6��,��^:�EYk{[z!O�L	����������d� �X0�^sO�q�t��Y��z��;Hm Ϡ�ͭ�Yl����)���}`ϣڀm��I<Cϩ!Ω��8���'��H�i<`:I�%�y���/�{�{�N�>d>� z�j���t���=d���:��q�2h��:�8��m�2xȠv�x�k��}�z��O��.,����̠��n�xQ��b��l9�l9qܕ���>mԙ�ձ-Z�a��
�L��V��#��_��DEo=m��=1�=B~2�m����bC�*x�I�z�i��M2c6�<awd����l��[뻂���o~k�xȰ=:�<@��CԁXt�X��:a�m�20�O���'l���G��::�����@�$���P�M�|��Bql��+
�L6��5H0�VE$���!����8�����9��ξ��y��'�Xi>�Y"��O���`jr�0��	�2|�]Y&���d��ݽ��<������ąH{�0�$���E��Մ)��Hz�ݓԞ�5l&�q�bC��2@�2������ok�Ha��2M��������X|���d�$�=�T��q ����'��Y!�����s�{����!�Cā���ROXx��V$�� t��H��@8�{��@��0 ��8¦������>���סM$:a8>��@��m��=Y�3� m򘁦]XI�&��q�N2A�~��:���]�}c׾}ߜ��i�	��l�0>N�%f�Đ����fRz��'l��;����v��:d����F�F��u�{��VM�����p�@8�i�`w�;H3l��Jä��0:g��!�"�Lğf���G���o헼;���<��@uM���Ժ���U�&�����ݻ�
�'�L��и��񫃡��`�r���R�o�'r��K�]��s_����{�o�~4�t�����<a��$?�m2!ēL�� ��OY'l;@�!�Xm"��>淪��>��>�����;I=I��� �08�i�M��|�4�s�;C�\�m�L^!��!��}���/3���ކ q!P�I�R@�I!�񇏌&=�=d�'�v�6ύ��C�N���l6�}���ֺ�;��^c"�I��$ |�l1 vùי$�'��&�O:��g̚>��@����O|�5������� 0��7�I�E1�;@�&�L�;d=`Vtf��h���|�t�@4�w���Ϲ�;�}z@���6�{��� k�')!ӦI;C�-�Cl<N���$(uO��0g�������7�m���=�ϐ�K�x�@�ԓi8�!6��r!&�m�	���'�yv>�̺���o�{"�6��=a�$>gal��=d� �'~���E�q �'�I�=B&��I���]��s���������>B}�I�z���(��$+!�0�I�I�&�E$�'���F�=d����M�.���;�s��}��L8��'�!��X@�HCi�8���LP*O�H�v�w̒��G��u�D�'�Of��e_z������/ ��/�7�V��x���d4�J�D�,�V�D��;;3��އ�	>}W�Q�uH"
�政#��SMq���l�D*C�'��2�
�hM$���!�	�a�V0�ϐ�wf�(1�1�R��u
>�%���LD<ܒ2x¼`w��d�u���$��HZu݄��jwHC>�4����s׮{�����q$��8���!�Xc$�ѻ'x��� P�g,�I0*N0����>a�ƽ��zַ߾��CI'{�1|���N�;>�d�	Xr�I�����G�� t���`yεr�y�o$>@�:Bv�a�VH_��'l&�� m$�%Hzä�oxHf�Bi�4��Y'L:N��9�l��}�w�2OX|�)l>H�|�N��'��i;9OP��0۶M��C�Noܐ�	���>@0��}�r�}��w�_x��W�'L>gG�!�"��B��4���q�7�6�l�����O4}Bg;9��?>:��u�v�!�'�Rx��&������!�vyI���E ,�2m�z��Ψ2g����K{:}�믾�Z�λ�z�N�ğ�x�>��Oz��&�ԓ�u�$�E�$�0�N2�m�&��bC�s�����Ͼ׽��C�HLO��C�>:�0ϻ���d� �jɴ�n�,!�bd� t�>}־�1�{�pW�,�3p��;��Z,�Sa�b�na6�0jtX�+uG�S��
R�G�Oc�2+�������(�&������;Ų3����2�M��*:�U�d�v�4�9���n:�,����z�K��í�[��o89ӣ\��e�����.!b�|x�S`+���5�8ӫ�2��uS�
���c��w]��r�Vt�Z�����K�l'�fRErV���SN�����V9䭀���|(Y5bN�DSyI�KW�j,�F�6*)���9��Z�2�Q��J�-1�&�\�yk;q�sr��[?s���`�鋫K���m/u���.Ŕ�2���&�1p��-4�WB��1����/rP�a� J�hh�v�P�h2]}B7��>��L]N�������^La{F����&bf�ʗN��<qv8��3�S�x����{�}����{�%V�o%��w\�G((!�;���Nl�P�D�]�����\ne��qf�:���so�դE�ΪmdeN���wW	MvNn9���7/�(�F���V�ӭGD���grX:��@-�r�Fe��o�*�33D���+*mr̿�C�v �\7^	�ml�L��n�\\�Q���-�(�ٰ�5��J��=�rV5zH���z�od�_eL�n\�e�fr2�\V.�{��(�W`ұy�X�W�u����*2�.;�%��C��B��S㔕�vV �s�k���Jo�V�pc�*鍔�k4>�̩����va����96[�Y��/GaG��[�0�M@�Y76��x��Ju)�kZ�z��κ�j� "6�۹j����>�ٓ��d���CKTX�Ac�b�����DUY�
�#
�������PX���TPA�"�UX����Z��TbجU�j*�,V#�r�TAQAae�(��6�1�V�,�G(�e�U�AcR�DT���[U��jZ6���EZ�ej-���qYe���V�(�YV(��R��	�{�f���e	v�4��A��t�Ծ�H�7.J;�h��(yjէ��=�yZ|�+�"|����r��C��m;>���<��<�j6Y��sw⼝Et���xm_*PjDOx�vvr�p��F���"��؆,�%��G:��v,K���t�è��:��u��`�B���iAu���<f�ɻ�ӏ���Ou��g�S��{Pln(�[�M�2����J�-��}�z7�����v�X[Uؙ���2�N�D��Rn�N���!Z�z�_�Ʋ��%7Q���ݺ��-�#�u��{==}��o<�(���C��s�#l#0f�)ʒ���ζԻ�B���5�x'i�&����Wu�yp�(���[<�܅.��҃�E>n���mR�_��G��Y��B���i�PP6�������� �ƻK�剏 ��ן}(ϭ�#��s4H��3�����ܔq��v��,�ʵ�&�g1��O���Z|꛱T͛s�1���y�1oK;�E��!�[��硐�[.��7�1�CZoύ͜����֥�B�{ݓ�C4�c�8�q۰��b�q7v78=,0��u�bRE-��88�V�t�ZJz�n�g�R�go)��l���������a�бevRH}�j���� �B���n�.�\�d��o�K��"
5y����)k5���Gw�������e���7O%��興�1���c7a+�p�
�����:9��;NX��=T'�p�vF�F�����w�\3k��wk�{7:ο� ��V�[%%�{ޏs�õ�Q�~���.�7�4C�w3ՙ�>g�p��U��G�^;Գ5�룼�xR����D�1���q�wr-u&���H�f��&�5��pXdSǗ�cyz�C#�bmyCm��<6�0��ݒ��ߑ��7YN����m�n���%�z�X�ʎʁ3q����F�Suu:� &{3m=f	P#����h�ś%E9b9{y�ch�U�W�5},��Ok��ndg�!��{��� fFn��[�^2�r$㟾���﫛m���ӹ�p��m�=c���g�sf����R�i��0;�.�����4X���W�6�)�$j��s��';��sٽ^$���d�&�ݣb^t��(��!��^rhL�5�\�T�#!<17�̛�P�P6�=%_j�F�5�A�B|0�g���p�6I��3U�継tS��o����3��W�D���08;�kƫxi^���J��1i%�:E�^y,��p�`�jY����:��t��P�P�l���:P�-��϶�^���e�=y�ЦZ��qj����X�$q�Eդڣ�l�:����W�8k��Qf�$��E���*�<M��(QJ�v 0����ވ��-}³�u���eY�ɕ���Yf����5���ܽ�g���W���Wْ� �by�iԔ�f��QS����B����Õ^��Sk��5�6weӬ� nL\'�Rfh��ߎ���G�ݵ�$��{�:a�7�/L��7-�T�c4<}�f�"�z�J�.l��}��g�����%�^�в/ا��)���5E8���#��W��Eѳ����e2�竧�_W��~��P��p��ԗ��C^�,?Q� kxl�>�Ꙭ��QA��c��Ӛ�V��`܆����kp�%w �t5c�ܩ�FKO.侈���!=|�or��-ݎ��Y�u�I��ث@O�&ۗ�O�qZ�{Z$�Vf��>���ܴp��QJ�Ł��O[��m��y=g���9�2c.]�X��Cx�c�W6��m�ҳd֧�S���1{zt�2|R��E�.w��R�qG�\�*�1�p�8C�F�+ӳ8I��q��!YV��g;8�yk��i4����^ɳU�nݟ?h�g�7��8$���+ε;�w���B�}���:�h{Q�Znߪ�����������ۺ��a|��8�&._f�ż�t*Kz���/=�7��KB�s�i�˴�K�ޏG��	�Sc����z�w,S~L^���Eq�Y�@�q��Nv;�x���f�ƥ3����c��-���Jt�S6�$���0�GT�ܧ��ʡ��3��nsˮ'|�s���e�)r.�﷼�y����x'��tmX��=9ߜ�WԼ��B;�p�z�Z�_^��U�����}A��gV�_=��,P��I���s:x��jP�$o��Ny>z+�dV\��-ў�����d�o����'��4��^�116@6��d�@����C�X��jo|&\䷄��:�v�,����o�S��u�Vb�\��-_wr�;���=���Ye󭿰F��7�,/�����.n�nx��|�P�6�i�6�f�\AJ��rCsx�*�p;��QX��Q�5�l�c{��=G�fzM��Ά���ۤFm���N>��~�����<��5f����F��T��X��
��={Ԩ��EG*�y���N]�Eg$obf9�X6㮵�Ɩ`s�q���j��sO��Y$�ގ���^�N�j�2+
�"�O2��9���]/Ӥn��T9U�׸��⏺�?v~�@[�*P8c����Ԯ���e���h�⸁~�ٞ�
��n���<�6�{�U,�v�;�n�v%V�9��l;�w%�����|���f�~�+���%���\�/�/��0�|���ǳ�����4��K�=#^��1EٜK����*\9ͨ��g_k*4�(�&���:B�|7_=R��,��X&��!�F� xu�&��S½�����x�M W}��2��AOM���=�C���y�����~5�&Ė�V�8��ե����Y���[�w���N�ޢ.w�N#��e:N�52"f����/8a �� �z�d�-���wc��U�X;��7C�7�N�Ԩ/���*�	�k��S��`ggT�-���n�sC�ټ�&9ׄW%�:����<�����UUQ-=�k&�G��Xf�b��y%
�*/s	F�/k����vP���[�)��*���.�"�3Oi�x�`��ݍQO�=�W�uPn_Sw�@S�Ϗ�d>@3�������ۼ�(����i;!Y�1�������h>�fڑ2J"���N�ʃ�I��5�lX�t��x��s�I�mv ��s�&2�P�9�s�{�6����Z�޴
�mP2���~�r��D��LmA��ן/���h�����St�0Z7Fa�.j��"6�8ŗ:�P�+nT�nQ�x�0�U�\+w00��VWcKbWw�����}�w�Z'O���M6(Z�	�]!�Lu�^O�74!���<�	�\��2���.����q�ѵ8̔(�2�@�qL�$�R�d(mȭ]��먯��Yq����;�y"����]sJ!hB�J�4�cpٶ,��gX˨hե��Q<�vfU�LD��8�|X�{7-j�����l=H�*ӜnV�oFۉ,�I;=Ƨc˭$��"���
m褰]kS!,<Twl��>�\�/qY�dm,Ut;& ͛r<��O4f%�ܷ� $ئe�Y%͉���	Du�(A�j�+f�i�śB��J���sV:�W��$f��Ff�M+e��O�V��*7�6sq�&_�G�=�.��Y��.I(;��7�;8m�&Ŏ����¤I���+���Y��$�oa;˫����Wtd��͋-Ezɽ7�i���nh�@��Q\+���d0'�,'�c�����-���\�7�ѕ7L���)���$%|{�2@�S[e�f���`��zI�sp�֏��y�+]!�w}O��@��z�وi�xJ�yaP��j�������Գ-�z�ٴY�+凚n����f��^z{�7�NܘU�G*���x���.��u�T%;"A7��9��{[���&�A��\�Ib����ܧC6�r9�]�M�Mp�G$|o�.�����R�;���1T�ܤ���%�ʆ��I xX�{]�8�`�:�1���2�5 q�gEzM�MN����u(�V�I��؀�H\'>2�:0id�ӪH�F�3v�-�UV�U,h����5|s�X5T�aFҥ�,Yj1km�D`�AFۙpb.*Q��\�P��ZZ��ecJ�F�+Q�+�TPL��h�e1V����Ub1m��hт�iZ�Ѷ�-*�e�cb�UB������e[IZ�-Kh[
���+\�WZ�)P���a�j�9�4㋫X������5����UEJ�ui�D�n.3Yn�m4�,�D��ʨ�j���X�-.d�摶]YZ"e�f�G��E�-m������m���*38(O��H�Y	c��|��w�7�'�0`���
�Q��9�fϵ�!�%��~�ޏG�Ikm:�D�v��$�R�;_l�d���BΨQA�V�-��ݜc1�S (;~G(�j���\���keGlU�+��l���Vw��h	[,h��&��B�{�U��[h�Ŝ��&�<�.1>Ǿ���c������j���Z���9bl5k���H��z��Wl.�`���w.�o�KQu�����=�2J��f{���f^�*�(���L�����Sټ��ֶ�=�S�~>�Xs_�i�y4^|��đ�9K+#�[�z&w )���WӪ��rඋ����o�U󻳤rjz�� W ��\��о�q�ºui�I������+���G�'�M��?f/�%f�(-9{.x*�]�!Fn���:�Z������ۮ��u8c�o��=Oġ��Ě�|����d��ᅶO�3=X&�>n��*��ǯ&	�})�)�����P��SF����]^����D��w������L�x6��;�\��U��)];�<��lnO�<�Ic&�sc4n[�f��|��:/`�}V7�P��~���z�\��z�q�%HɎ�G͒�\��*�z�bt��wi�We=�����N��.|Ft�,���L/�=J�����5+���m��/�N-�vSC	ۼ���o�,�SJn�	�=4����k�z#�/V>B����`D���َ��#��D%�!>M����U�$ u��0�5��Y�ًOgn
�G�T�@g�d����v�}s2m_m�Ta�ak�K������yD/R�׸�:�/�oS;�����E���e�<sC7�A�~Y�_A{�E2c���+��ƶNt�8%�V�9���-wk�������L,��.�C�-k��_^;܅�;=`���2'�����ܗ����=d�WmU	F�t��s7{9�f�ּ���r�er�hD��z�5��Vxx@��X�Սc����:� ��� �")�'��r���$�U�DRM�H?}��a�Vw3�tk��Mƀ;��,�����ƕp:��r�1�O?
Wb�buO�Ї����G<���3��)�7Vl}�{����os�A�`2dH0Y��;}��}��u9إǇ����"�]��!hюx��ݓ��S��7�4�r^}x�����z�yѤ��#�U�e�W3s��I�{wD7[�=8<r��!ų~è/g�[����vhB��G������ݞڣPw��e�5&GY�F�w�Bga�f�ۼ���j�Ͳ���,�Ι���Ӿ:���Ʒ�6-I,��/{D}q�9n(+�ʊm�z�-���z���+W��{ވ���rk8���L}eXب�K�����9SX�����/����/��9�1��]ʑy3�s��`����ilԲ�}4��R`�if{%tv�@qQ�tB4{-�i����`r��oO����� �����y�&ʃK��՗�x���v:�1��k��S�Ш������|"�LM����{
�S賹¦;C9c�b�Z-�6܇�}^.��x�ѽA]��k�ᣞ8�>��V������+��
*�4
S�-�h"��?�o9�w�'���7v�����]���R_n-:���L[���X�w�;b�Xï�lz�M)'�����H6�}cr2H�[���J����W>}�q*�z,��k��Fus�;�F�,�,L�~tV�L=r5�	��G��c=cy��+β����Nb�!�>4�B�����7�~����.ԧL��S¬�r�m���<:h�<9��Sj�ؽ�1��;SȠ��'q�0�o����$�{ �]�Z�q�t���	 .��)��V�=br��°Y&���.�S�XOk�w���ZY��(@�P���w��J�°�?q�ݕ��]
в}�vɖg��2�����0�;sn�i��[ʇ�>R�^��Gz&�:"���]�}�T��0\�)'ﾯ����/?M/�������O�V�bx#��Ս���3����*,�$�u���ag���g͙�}W$���������$�.�(�HA�X��N���R��Wܸ$�(���Ubuh�p5�l�TN��;�4���Q�m�ri�Y��}y��y�H��޺�\�7-4pi`ܚ�Sn��=x�R1)�J��K�+
7���S�Է�]�[ʰ����}��w8j��o*)���ÛU^L����עya�ݧ���b����հ�4,����@%G���^G�ӹ�������;j�5W�l����si6dN�n͇�p�$��U��Un/�?���|����k;��{ ���O��������ժ�K�wX�I���o��k��b���EA�f��˖��I�̄Cל�Xalߟk:��݅vշmҤ��	3��n2x�A�f���mGJ��Ɓ�ٳk2nx�R��w��R��v�}�lk�klD�㾔�i��\���ː\�K�?N3a�����g��f�9rK%���� E�a@"�N]v��*�����w�yu�%��Cג��"F��@z�}��kq�m�ZN�`t�w&�i����Է���!\l�S�e7�����%��5���>X��v`$�Ԏ�_{��B@��Y��b~�'�6O=L�{ڲq�|�u�-:���i�k;c��wMk�ٶ2�$NX���an��ؚ�'�y���w�dJ3�{b�����Vh>�/�r�<\���O=56�˧WZ�o�1�k!����!>��j�uA7۔�yԨ�+�<�KL����4���@�)���o���}��B;�*����>~�:B���~ò�G��#����zDC@'ƽ�<�`����~�����ٙY��7��V��t�"�����2��e⨺���(i��W���'�d�(�Ѐ^����c���	|��ȱH��h;�~{��U�Zk��7a��7Y��5/g���d�jp~���&�u��L	��Q��x�憎NE6�T"==U���[a�������WGӕ0����t	�bs[ުMݍ�P�2`��U��*yOj���V`��E�Q�\���GV�ۗ�_7�b_��/v��U�v&0֍�Ww�Ԓ\^t0����+�����p�/���c�I9��]�#�5c�T6�l
����R�����1�@������tG�U�[�l�?�Z��g^Q�&�Z��n�w-�ĺV[C����lD�Ǻ�=dVcm�m�]�q����E#4]-�].t����;IYW '@t�����#�cP�Z���T�m���/�^��gR��������t�z��c��=Q��@��q�8�#-�&��#�(��y�e�Ρ���x�lл�˥a���Jo�`���C�^򒕭��T&t��:�����^��n,[Fj�ޓ 86�n�Y��qj���k�>�D�Q��Wa<��ۊ�����0��F� Z��{�� �C+SD�첮��>s�+͛K���M��+����M��̺R��en��mБ��i�X˫���qq�pd�qر����i�Ө��'kyB��������fS��!��.�8��@p�����,�yr�4�+��XޘH�n&KH� �Q�2�q�ގL{�j͝��Ř��\����5B��!]��p���M��:q�K�4�W:��L�w[�'jg%"�&�K�*��ܣ��"��nEK�3�[�)�em�Ϙmk��j��:;/ͧ����ZUl�!��H�f�mĬ^Y�ꒂm�*�wT+�q��	k�<]6�G)Fi���/,��2R�OY�~Ƶ�����6��⑜o�%K�tb�k���5��X+��v�M�9;� qͧZ������rlC�3��8G��z����#���ze���&�}z��
��d�������k67�Қد��6�����Bd*���y�j�Y�v~̝�� b�Ws�\�՚�6q��l�ݵE%%Xd�����8R���T��J���'��a��v��s�⶙s*6��L-Ƙ��.��-\aF��[u�1T2�+u��u�b�4敤�fj
cZ¥U��b[X�U%��h[E�5�-b��*��!�Ym�TkQ�Q��Y�@�J���`�
�L��F0D��u�(��-���J�D[lGT�ŉ�TƋ���E5eA,U+Um(�5t��b�2�,�cV���1�D�3
%ˌ�]Z(�J�2�3�e���U���֖�TQ�+1�Z ŊcE˔�U5n$����e՘j鍹�e��%��r�Mh�i�U�\�M:�.��kn6 ��m�m�j�CT��Me�Q�EKh�-pKmkJ�������~��7�����ݧr<��epbt�+5b�XF(f��
�p�I�x�D{Z�w1)XP4}ۧg�1�[���^��O}�ܠ�k^ta*��[D�R��K�M�2.5b2Qɋ$լo:53�q�ƺ��j��}��i0'�|k���V�׍��	[���X=`��ɳ�RN���r�V�y��[Vn��]�4Puz��b�Ľ=���]Tg�9�^j��G�C��8�ǭ�N0��9q�=ԇ{>�׋��ԫ' Jb�X�OY��+X��hk��x�Y.c���I��ㅂ *�r�9�������\_k�`d.�ՅdKyR|���+<��ʿ[�];�ǻwQupcqF���O&�zn��"õ�1����$�#ފ��g�Q�֧�s��w.�^��:wsy����\��MWt�|VE�p��]�nk.��sW���ʮ��=�yL�G�6�y�,�SLЅ���Y�
g�A��r)�G��;i�� kMF6��^�=�]k�O��d0̃~ί�o4L^O��r��^^x&��f���׽
����>C��?4���ළ��u)}��W2A�4s����m�V����=~Hm��x�v���0�a�n�khJ�ɸ����,W�����=y+8��bܾ�;���(�ը��=s��vz��Jll*f>�/q(�,����=�'?}UU~�|�o�)����]Υ�aέ'�{�*����,������Z J֢B�q�9h�@H��jg�E��=a��|�0�nGr����}[gU5�(ě�s����xX�УI��O+ɭ�����0�]�%���6�i�hgW)�-P[��K2\��,������Od1[��>Koay���(AG^�7���	��/�� rt����O@���7�[��$��l.el>�o
X��u�,}s�;,�$�r稾�ڣ�����%�z_�zGe<X8��8���ֈFY�����d�9�N�o+Z���ͫ�T�8�G����{އ��|��������M��r���=|L��1�wwj�P�u�4V=�ve���͆l�Qo����?o����Ў�֗Oi׸<��V��ɫ�S1�g"(t������uǪo\Z��i��w���e���u����ټ����lU�,6�,�YUvO�o+�%��wy�ʉ[���6�L?3�yWP�vt3�P�c�t$ ��Gx^v*�A`��-��E��{�$'F���~�ˁ�n��=ε��q@�"cpE��zAVF{ϫ�^�n#O���i}�x*{U{J!F�B���^l\i:�7�CޏwR�٦t�FS�(�v�S��M�]ZJ��z=�Y��of/~��{���;�.�k�D���|��|���}"7�Ϡ��{HWdu5;
E��ۏ�)��@�σVhrV�z֙%�A�k�[o2˂�Z00�y�5����Pl�5ouυxq��%z�s�����>�i��VPy�GB�Jw d�17�l]�-��3"
��ݘ�O��#|B��{��|�֨��kݛ)w���/�3S~�����t6�n�[Οb���I�p�H�<��A}\�Uj�����Ff7w���a�K��-ꚪ�
���-B�NO�]S̽��sE��]a��ⳣ�l;z���P���MnH��P��Zw�%�{��ͮwZ�vvU�/T+̽w`r���Q����9P�4{�I}�[�_n��s��==Ub�X����7-�=����Nt�rzp,3
;v!8�ӝ�K
�����o[ʘ��z�T�Nme��J����5�Ώ n�4�&�\�� ��N�è�Up_TѴ']˼zsFB�0:[�w�d�j�x��7�r�Y��Av:J/�X�S)d�MQvo��]�c.9�rz���Y���skZ�}�jԅ�
jj܎�lwJ�7�p�j����3Y9�*�^vk��ʕ�WY�PхWM⦺�$	�6	;�q���{��M�� ����$.��|�^��g;���~�t{6z,0mxM��W��e�!~#�cY�~)��a���o�0֕����~�˪������\��P�"(o���CYʇ�hw��O;�w�s���%�ˊ�P_;���p�gWeseicmHw��e�s�M��!�X��p��۩�ō*lu:�ou�����S��w���}k�>B�:4���;Q�?r�o^O��3�J��@��<��o4�j��$X�������,�v�Psu��U�(�Kmv=���gT۩s��K��v=�9���W�%�}�u�&d���/��KX�$&~͚��'�Dk	�UM�C�y�OfEG9ލ�p��z4�3X@���f��u�����M�j�?�YGN6[��)�K���Z��P�:�4<���n��[��7�N��V��#HӇP��=X�5Nx:����D�U7�q���J���pI��qJ<����Mj��8J��c6��{�4�B�����ڟ���<�g�m�ɳ9��P�8����<�`h�_|�����|)���|���;k��Et�2n�eU,�o�N
k�	:���FJ2�u��3
�:f�2\��B�`o�4����ڒ���叛N���~DA���0\T�œ���a`k�Ǩ1hv�֏V�ұM���ٗ�f,kl,�V��[茺���/uo9.',j��,�e�Q�4V�M�M�#��鉑X�w���J�\O�{+Ω��]��W�e�TޮwϷ�=����+�j�rKg�N-f��<�����/p�;T�4K�u��x6a�w��6��0���7�/�O{G�O��r�Pxѯ:k���;po{��`l�7���wwf��mR�2�R�la��"ڂ���*�kJܩ�wv�^XjW<��Z4�N�	Z܅F�ꮑF[w�L}����}9(�*�nr��e�i[��O�����w�W���b�Ϲp��j��i�Ao4u�^�{�	����p�]N��t��s���i\r�(]���M!�¥�&an0���f]ed� ��{�|���C)�i�Q���m�߸g	j�e�白�}�Y���]��K ��������Ø\����=�B��ľ󣴝�o+ؚ�X3.oa�/9Ȣ��,1:zp���q|�4�Ontyo�b��Np��������6����&�wk�Zd)�:�u�I��k2����E��3�&M�j�����U:|{�N�$6�r� ��H��ʴ��ݢ��a:;���8[�z%�۳/EP����s|�)���Y���tU��u����7_˞��3�ی�gv�;�qV+H�����+,bZ:bU����U^4���j�N�o�b�7�\�E]����U��iZw�Q�S��Kc��PgF̱�e�V����5�dk]�E�s���	>Iw@3:�R� �;4]�1�F�yw�$fw^�E�yAc���e=ұ����ċ�oo�,	����ý���]j� ����gYQL���Q�%��={�"�۪�[1
4�rs�<Ҥlvbz��XY!��uD��(�H��������[�y�i�����2N��s�����)������ʖ�f���4��G;UԤR��gIb�6�mWY�C�VG[m� �rqvob촯3P��݅��9���eg�b4�#���5�:��
�i�͓z&���Ǚ��/��8lCHYj���~�1,�����_&�_�)�"-k[�y����#gb���b�JV^���1��y��t%���(�^��l��ڙ{i�#C{���Z��拓�lL��L5x�I��:�T�u!�+��Y�z�ռb[�]t�3���`=��pB��YI�{� ��ce�iu���o�a����ji�$fB\/dx�YXԗw�2�I��d�Z�wV�Y���1�fMW�),W\2]=эvb�t����A]��SJȲ	���V�R��ػC�G)*T.��.5I�1R�k�j�UbȰL�D��
*T�H.%KiQQӆ5j��fe� �1%E̪+�ime�b��UTDXT�WT��Ѵ�")��q�u����5��J��(ֱm�V�̒�cˎ1@PUUUD�Mj����eM$�V����sVeѐ�Ց�����b�Q4�\�-c�*:ek�SJ˖P�&�2±ʫFcSIh�&����UEb��r�q��J�s�����.R��
ʒ�c�nR��DTQ%�3�����8�i�N93,��B�Ab�A�W��S\�LѪ�ˮ�ד$�4�^��38mjuy;��C/�1�#U@��ԛ�"ӟ��>�k�gx~�b~��xi��U���N$�C�1m�7#qC�QTW;���;8x4S��]��۹f� ��} �,�ب��7؄��ħ�`�7Y�:�	dʌ�B^��yI�5��ܪ��8���tg�c@�׺�j�x��97�;:�u@�DLͳYs�0��+�D��Gݼ�x޼�Y�ɞ�^��8���6��/��Y�{��Bg7����):��7��E&��=q��l�5��=hR�p��&(��5�M�֛�f�׋Yu�K*��W�R\N�y����;V����)����	�{{�\5C����JC)�\J.H$��_&�H�}~��Ԉ����F��C��5R����xp�[N��8���.{���{��[�er��`�s�Ŵ�)&Vb�nksٕ�-�i��j�g�����2i�9�{E��'FQ0�.��ݭ'&<wB�ދCb��Q������2��h�r��U
D���0��Y�ݙ�\�X,B���k܄���ݔt�0��N�ݯW?9~��(�^d�Sb�Ɔ�s�`݁�,"[;Iev׺���M�O��\��HgHɌ6�ߐ̥�^�V�k����GyB�s�εd.�(Q	�q���@XcU���6�Ț��[}QŹ�3�#GGS�d��ę�&���i�m��Q�}G�����Ɖ���=�8`���꣫c���_y��
:_��+�����r��8Q��4]Izh���'���VW���V_[��١���kE����Sl4;;�~��Z��,b����Z��c�4��k%���9��S��_o�>>!�:���&�b��t��w����v^.M�>�ϼ�+��#�#'����a_Y�Je��',�&'iLΚ��pvĈ�dB3�S��SF�x�R�w~�ݔ������j�"F��L#�+�B�:�r����z��TS��M�5�	ӧ��yt��Y�@3D-r�+�E�Ck~�|X�����b��@���j��ctiV$2��U��B���a�`G���*b�ˮg�+>��v�*�g��p�n1_eΉAG��0J��,���H���t��ܗ�}��m����"w#��
���8D<h��+��9�����ޱ��9��׈'�Kz���n;6x��Ԁ��WX�Hv�{��8��}kj,[� ��'l ����lSx�6p�i�Ιs3vd/9��{6
��	�w0�aGA��9��5
��w�^�[�����:"�6e-?o��џ5�䷨O���.��cm*�^R^�p,E�d���.���~����Qj=ۯg���D�ٞyN�;����O+�;\��a#��q���"y%�(�G�_A��+T7�l9�f���`��;�/zL�M�d�䬨��'k�)H�4�])��-,$[��T�9/��?;���P�vԁ}�#����z3�<K~���[�i�ӈ����Q�k[�yGK���z�I���N|��7���|�e)��&NfT�Z���R��������&��3�D�QҪ��T��9�U�5��H�#g��n��-w2�=W�,����0-<��_v0�L�[vA;"�9cF�]Cݼ���S{H�������^�Ǜ��wZ3aD����!6{V���AN���$gش����pw��Շ{�`����f���;kORw��)x������"������h&<�T�	^P��w�b�Λ��V�<Wֆknxs�x�K��˩]�ц��<,5�v��^��)U����ִ�ɟ��7��r��~~,�g2׼2ez�o��[I�h��m�c}pU�t]t��F��#�<��4wCE��������GhL��b
����1GƏ����a����F�-R;;^	2s
��Xv����j[ʝ�s���c��l��w]�a�ܮ�P�-�:�l-����٥G"[�����y�R��<���F$�쁱G�|��TqL�����n[Vş����\w�p�(����<Vc�O���>��7�!~�,�[���8��Yz�R;'5��9u=ݬ#��b_���EH�j�}�����T��fgܰ�����}�؆Ri(|� /��Ŭ���9�kJW�l�Nb�S=p#C�S5�b��q'�p!�"�:{z�����sc�h�ܷ�����=vQv���e�3�_�����C�/-=�3�R��y<BD����w+.��՝�нLi~��%@�T���,�3��Ӿ��u=��]՟e�_�\~OC��cՎj"A9��Oo��3�����憯k|:���tƜ8�Tt������������2彺=r�,c�^Q�4��㫗���ޗŶ��'��U���3���F��Z��������OIW����Vg��̀���!v�6s��!O2q�8��r�Y��S��w;�覨���r��C�B�Z���v�nđ߶�}��L�<5B��Vk����p�𮘸�n��o[�����-h[������9f��cO�
�P'ǭi�E_�в��f���<W���̮x.E��ZK
5�_��j�;!+`�C��f�F.�l�x��v��ɖ���x���śVƝ!�,�B��4���rj���^��TF�(�>�zBE��t>���Խ���wD춉]
/�<����K9i�ߩ���E��W�Y㢟����i�J�;V0�n^S�ܺ�5�z������'�`���:���p.2[̇Fه��E9�νIY�
2�H�"���+������|y�z=�DKL�kzM9��6�euDd���0��L��*�-֤FҾ8y�+)L۹�|��k��#x �]0��1��9�ј�=�K!Mc���ě<x�lj��q�Q\n2��k��mr�0����~r�aҷ�z_s�|V���_��_^��Guq%�b���8D���~[�uECV:�S݁/�:[̌��qM�dL:W��}kIb;,Z���@eJ�{��F�}�������'��LI��+@��̘˃*ce�3|!���Kڹy���;=V�<C�_w1g
:�C�ⰄM�D��FGTKv����w�'eͥ���?1�F
��r�/o��Ըѣ���	�u<_x筍��*=p��}�ͮ��"[Z�%rv�U�����*�</|	������d����ikL��d�.�GXqo����c��W^
�m�85֮���y/�DD{{1�ټ�s�GڨD.�í}�JZG�
OM�%m�j���j���z�PB�_i���;CQy�k��}t�ue�O�^�ۗ@�����0������-~7Y�=��/���}o�0���Y�,;)��1m���DH�ͿctK������P�9�q�7��5��^#s�l)K�U֭���|�":�z4~�\G�`Z|���_���MNN`yխ�?�fOΣ�9�~?Dl�~�h�Ԏhפ>�J����o{h�2��>5��O��~@*��c���
&���h�&��n����
�nY����|uߎS�^�����	Ƒ��z^�����SP%j�8���XG�GgHC�ۻ�^r����AXk��e�-��\����[t�+�n%������<{�]�:t����8�&�So�;Wm�"�^��rqRO�_W�V�<܀�~W?�~1�
2�����ʍ�O
>7�nb~�r�}hX=H/[�z����]��r6��ͺsB���N�=�^��2�Qb����b㺶/����<��~�b���w7UN5ྡྷN|a}5�������U~7.MUm��;;/��Q��zhĂQ���O��+�2���giw�ә~�׏�_�n�<x�1���3��Q��m
��� ���)I���Q�~��eq�_ �jkt��������/{��6�_gL�㫏�Y���+^�Vk'd+�6+��q���u�[kn�]L�CΠ�)�,%3P������?���pj���ݐ>A/��b�T��!Gyq�&&���?i���|�� {tH��X���%Y\їEԷo{���&�U���Xi��Izj½c4���WȞ3X�j�������:�^���ߒ tN6s�n��ջ������.!7jwq�ek�����T�"�`��)����pm>�c]����ڊͲ��%��k�F����{�A�р�q�r��r�h�|�R�0н����V�r�����TPRQH�w,z��\���g5�*�n���s*����Yy8���o�����;�Cb����+�>R�B�#��
��u������W{�����1�ʇ#g�7��]%&�rD)���4�\̭�$*l�u��Ǔ+Z�L������ߏls2jw)|�/ufd�����{H �A�ɘ���gnh�"�i���b9m`�I�a�]�a���X��.&��49M���_Si$m�L� ����r�g'� \n��<���C��:1M�3[i5l������v
b���k#*��J|��wi#�w��Gf���6�N��H��s�"D*��+�����ε�I��ԗ��UU���w��?�#W3r�a� ��woM;���+wR�Esi�S����l#�c~�z�N�,���2�ט�=���c�U�V�:�9W��T&��y�؅NɃ��]Zs�M�|n��m�,;KP��Θ�ۓu�w�]��]��zY1t޼��N.ޡ�:K�*��8ɘ4f�v('S�4@��&�0"�*�sOjga�"%tfZ�RK��ѽ<��0�*��mȤa���x����.�z�6�ٶ�s�Oz��j�뤦 nx���Xp�'ޜζ�w�눤�
���Lq1�%E��C-�B��!�鵵
���-�J%�Tm�U��9��10a��B�k)��iiB��ɘ����2�Ar�
�%d��Y-��3I�Ajk,P�k��20ؠ�$D�JȲV�����kr��nG,��ز��2�IL̬Rb��E
��#�WV�f5U"�˔PR�1X��I����ո����V�*Ue���V������2eZ&�L�[E�X̤S�E4��㬹Y1&2�&1J�R�t���]2�re
�H�m���L�a\jL�V��5��#%�P��Ӭ�q4~�����e��U�O��{W4��YpE�8y��>���4֮ų���fD}W&Y��rl_Kڄy�E���A�Kw��+ݶ<%�Fx,!X}�3�0��d6���w��PgQ}�~��J��s�{�˒`�r��>�!�C<�zT��z�z��D����0�X8�c���dV��.�lٗ����/��l{
-q�s�	�������=m��є��Wג�:k���*4q�w�)���
D��xd�n�ҍdŷl�DE�M�Lu!��B�b�P�gdS�;�Fh�xyB������aZ����t����õ���tۄotg[sQU_TdL/U9Co��9�ОvX���o8�Wj��">�|ívz���!��Vå����:��+����sl�J� m��!RڜE�����0�;���Q�\WX�)v޶��uH���1��d涮�@�p�
s��U6y��{���qs2Q�!Ʃ��_C�1i��6�Ӡ�i�oA^yͭ��f]5����<C=j�e��24�E�vߢ^�y��a�<a�N��_��a<���L&������ �@Y�sӑTYj���;���g���u�}�~�?'�^6���ee�~���T�u�oGv;���R�:�\��T���n�UG!7:2�f9�ؘ�m��eH�,س�yq'��<A:tߓ9��k`�[����FG�Z�S�Ś8åZ�ځ��F�%	F���&C�2��ʛ���E���㼴����u�s713�P��l-�(�ž~0Z�b�g��]K"�x|f�x����\Nj�a�
M�p�\d�wmMx�5ʎkf�}.�nr{'2d�,�7����s�����R�6�1�~�$!r��Q��}��9�3�la�tA�c��K��<%�h�y��g��>����R��^�1C���:�փ��r��e_mP������o�c�|��6|_,5-���1��n^O9yn���y��[�~�����J�O����{����sV�}O�4B
?jd\���p�D*,=�e|k:�f�C�j��a4���Frg`xG���������i�yȐX=��������ԸE��e�	�-}�x�j-8`��q\4~�3����z�E�*ô���"�L�ء^�+w�ʄ��q�B�{��i'�/�!�sFf����-%mS��1b*��>��&�$;����C׊�j�����ù��m�=�wQ�x�:���/�y[Cqkk���;w�R���f��D�f�6գ�ќ���cV;wE��-��0^4\`$乢E1u��^���{N���4j׊/�4#5#����9�6��8]xn��9��X���z�X�DV��5�T^v>>��|V�l_�Um8�g��=�����4�&P��^��m�ji�~��h'�mi�d3��dyw	���L�ޕ�[a�c���^&ofAdV.4a���9}��%�j��ct������L��n���ƹQ�ψ�M�pȽ�/k������t���3����=՝��*�C��D����kx�R��H�G���;5�sY�qO!�_�3�2�l�=�>9�H�Ǧ�H �� lQ��nd�eu�5ʿo5�e���9��.;���?�\TVQG�!]1 ���:��L�]���FF�F�h�v���,�J�5�>�s-F!#`��p^T�fq��F���39�V0X�r�����6��z�r�����Lqcm���8��Y�2��%�F�-�Nʒ�!���ən�'�5�fD_1���!�bӋ��.�_w���4w�ܘh�R�b��L8�@w+<��&UN����}�C�%\c�_��^�(�K��2�+s�����݄�Y�6��&r-���]���vQ��m���uf��H��ƈ��W��	�����+���V��`.��$���y�כֿ>�B�r_#���!�����*�n�o�ݻ�ͼ�����y��q�b��z��@�`ʬ�{��ٻ����(/��Chba��Fs�
({�ګ���{�z*�\��y��[(y��QX,B�ve�� ���\"�b]K����FH�5zn��}�+
����Af�՗��I�:�=g�BukW�J���]��*�Շn�"���JU��[}M�����%-�}t�ߞ��ڛ��@��pSHe6�v�wuN�G���2��,",�������j'iiWLf�Ʃ�$4D��U���xF�{p��Pg��ؘNTs��#D�ʾe-�x�,K~�^>"�����r��|!w_�W7]��骊����u
j��(F|aӘ�Ä�� �J򽘨28���ڡ�y��Z�jo`�xyqŕY�}>5H�x�d2<��ӡ����5�S�t4�T���,&'i�xg�� �r�ŧҙ:���+��p�~�*vg�ޙ�W�#<U�uiԷT�+-��0�������v���\�c������HC�cڽ�H���71�Z����^*�x�B��أ�䲠�g��){8�w���8�cb�}(�)��3NбBp.��ha�Ngr�:���_=�6\RH�pD�]x���ۤ>����W>$�\x�`��&sq���s��o���þ�1��G�YT�:aR�kV;ͥ���j���J�����a�w���|Y���c�?i�����67U�m��k�i}l-�a��?���k�ٹu�'���6C+�A��O��=9���S|B�	񻧄�:{neJ��ѧԇ��Ŧz�;?.̓3�&�@4�F�v���n�D��2:���0^?���Y�l���K|~5���jJ���p0��0Z�VCպ����e/R�V��s=v:�0��m���=vǞb�L���'�jKH~�3����$�K�ZjWI�33|g�v<�՗>���>���9Ξ�{�mM�O_f��Z��]�l�u&1��g�w[����`0�.��� �B�Kz���S��)ޫ�}R��V�Q�}�o$6��F3na:R�����9"cj+��_�pOTw`-p&D�7�t� ��4;>8v!���v�ws�ig�{ݨw��d�aYa���cX�zb\|���`�"D<�+����'�M��\H�/�C���`��Rz���}�k��Q�L�n��y�ӣDm�苵��l��Y�}���
F���ޞ�	�,4t���2��
�4EK�P�Y�ꈣ��?���(=O��f�b&v{o��ێ�������0��mҕ`��9J�p�$XQ�G�U���ؿzl�!|��<��&ofAdV/0֠o�����s<�(�y�,R������pU)��\�Y1�r]P��6�'9�/1:\�~�#�+���h��-Bx���3��ιy����+��S�[�w�젢�@�D`���V9򠡼��p�[r��)��{:�u�b�|���Qd���|T�m������!�G(�l��0�������C���ImŚ���$˓�z���NH�TW�_�TfW�[�ɮW.w����9.;o��R])�P�׮T�X��Y�[$�e����L� �Jʅ;쾩�f�(�yJ,��>q'
�.�÷ޔ~as��S��*��X�D���>B_����Q��թz-#b�G����j��T��W<�'����� �q�Ez�"z����q������#e�z����D <��:���g�-qaǧևf�(�xю�n��~����"}�h�@�������9��	����}Eݹ�3Z̎O�#�/V�	���^�X�7�6"V�s"����:����ҕ�s��e����Q�p8�(
r��E�܎�>��ʏ.�eA�N�CN�����j׽^�%�پ\o��j�+�p��N?*�������q1j��u^�`� �j��	lf.\�j������U!ەc[��ݝ��u+��Xl�!�FŬ�'.7���K����ԅ�3ʹx���F����*	��t�<ǉ���hJn�|��	��5q�_�L�T�{+�(�m����G�y�Fݻ���Y�C����4���E]�U���y3��0Ze�{�����Q�c|ív{��9
���^�nS�ҍr�V\�J:G��o�
At�����8y��K$��hZ
jD^*��<x�l�sX��r��1]�Y�D%+�t+	_tZ2Y����YY���]��$7r�	$����'�3O;2���}B̎;�
z��u���u7��Y�a�J��L|;�QdM�E�[����{2��AZ�󎷰�MPqP��n� Z�uW�P����k]��X��-ע�D+��:�Fub���$�� =r�{,h7�y\
Q�� �kz�C*�ʄ#�[��u�f-p�_K�R��od2&j�[��Ql��`)g�鋍m�qc�/�q=��A�3��n�;q.��.�r;��oUWK�2��� +��05�NA�ze��mʊ���QJ�v�_#mR�pu
{��]���9�ɪ�p�x�_qHtړ_lO�ʝ[��l�ȇ�m�����!ϳ�i8q�7�ٚ]�v���<vQz\�k95�`�8���Wr�C����<ot�	|59Y�4�#d���5wά9v&���5b^N7}�����+#S1�kF���j�Q�6�,֠�C3���o��5f��o�s��߉�)<Oo@�fʶ���S%�6�;�
�ۃ�eNAU�X��@��g=4�P��V��-�ٔP6B�J�Y����9ԇ�c�+�V5��ymk<b�n �t.����a�ٚx��qs��G�G�/,��ֲ�ͻ�Ƕ�Y��i�
��c�͔���Q�}�{�B�D��f�y}��
�:�˪��w�j����Em�)�Y)�p�78\�ç$t�gu��Ʈnȡ��N��gO.̴�'���.X,
6�q70k�Mz������rn�%΍>����S0-�^�����y���y�;��Y�2fUS��&����f]jU0Q�\K���0ʶˌ�In`-h�m�QH(�b9a�QrѹLj,r�WM4ܲ��f$*E��ˋUI\Q�r�Wk�S3I�F(,�WL�.\r�m�T�C�UP�̦ ��,@�,��t�!U��1C�� �i�6Y�+UĈ��J32���kZ�R��Q�*1�2�KQ�)���m
ʊ:��"�.ci����-.Y�(�10,jZ�U�Z�c-(�h��J��j>��:��\�}0��a���E��c�B���z�xv��2p�jL�
NRp���@�c��b,!�(�n�yw�.���.�;f�W�<�"��"��ӖEE����߷G�����s��g��dv'dE�L�-��V[��ӓ�A��Fb�F�<����C�3�3��5��$7��8Wf��w-�dz �dW�����Ě���5i���5OݛV��}�A{��Q�T*��Y���ť<z~-v�{;Y�iYT��N�v|p���Z�C,�D:h��:�w�w�����L��8�����a��?:M�ٳ[��']�K�f�ݬ�v�&�{ ����bb�!ixܜ��u�{��z͓�c�B�֛(�+?X�l���U~u^�V|4�\�J�9]�H>J���es�[��/���HdO/b޵im^�o1��fA}6)
`�KY����!NE���fGA��B�c��@���Ѱx��,��L�z��^�y��%g��eYmx��r����S�����ll�Ad�&K}��7�!��V�� ��W�Y���WLWeFM+S	5�B4��RU2��C	HQ��g&v<���q����{�[c֡��w��E��K�qk�� ��r�l63+V�Ǌ��.DQ�&\��jCK�Ь��ó�cu|���U�of�j���="��(p;xƞKI<o��|�)vN������7��!�����X�<X���6;���+ �S���}��5�Ŝ��t`�5�荟h��~�ՙ�pu[G<��KO��p���g��t|@�U=-D�4J�O��-U�v�U�s��'=|^6�@�%hܛ)'.���s�I�����,A��{��þ_F|�D�ܙ����������u�S�����{%���t�+{��Di���<����{>GZ	��SP'L!�>����T��5�����Y�l;��A�a���&/a��O7=������\v��a�F�a�R�w��np��|+N��Rez`H�j@��t���2tb㺶/�w�����u���B~tp�	6m�,�\�,����x�[���:ֽhs�X�G�Nj�2�w�Q���WX�GY ��w����w##iu9��PS�t���Qpo�)J���e��J�9wW>+1�<x�Z}��6����Z���Q����b�C�3��'�N�G��T�Uk�>z�����m�~���f����݃	�����X༎��S��x���-`��ao�q���������1���Y
�PAսY4����|:�vlb��Y�B�jD���71E�$��.�O�Q]D��I���ʙ����� ���7唉C��K|���n뻷���PB�Di��ua�L��B�x����C�^��u��u(�/�pa=��H�,;�3�0����������N3���d�!�C�w�y*3���9g��.�x�w��,�k�m�#�35�>�P��v��z�8`S����	��J�x���e-:gs�53��`0������gf�\t��=��F�������b�ϖZ={<�!��-%�~�S�g*�<�z�STA�M�c���^yN�t�����P��2�(vn��a�g܄�h��j&��(�/�e'.�����X�ش����&E[�}��]GF1��K���h��Qp�(�u�hi*��v4e��g��)l�<���x�d�)%�"��.�p�qʱ��ޯe,�,�!��T�i��-���w�<��(=�Xk�N���y�>>Ѕ/|���W?�F��e��ޱF�|�yl���D3��ú��B��nI�|5a'���f�мS�(z|�<��e�u�ꞝ~��p�lx�>/�ɇ�lBAmӮC�Au)��C��s�݇���a�zD\v��8A2,�"������tﯻ��O�c�����}hodRצ%��?Y�L�6��r�2n�!��DoO�|�M^|g.'Q"{�z~�&9v>'Mm0�t Hp��1�Qr$Lm��n^l��r��٠� Y/��^X��:Ѕ��],<ZR�p���g��~��<����E��ø��g7i*.41����\(������Dwȴ�0�&_-� 6��VZ*�zxI�KI8�i9Q�22�e_�گq�Tw�K��(�YL���]՛��t�yX��bV:�T��_�T�vm��$oI�@�o�_[���ÕH��7 �胼|B[���	�z�|����%�_!e�Xl���������^�8]���[�ζn���mB�
�R��NI7K��;.BYTv��l��+�l9KO��#QG�9ʈx���R���{��7�.��*6z\���&rBQ]c˵K�[N��ކ�lz��9�!�z������wmR�sKc7=��P��-��v�e(�1��'r�6tѣ���U����v�F�q_/�C�<��7Wn�$,�C�VW�S��%ư�M�)��0[�y���^Z��J"Kj�bN˧+�b�`c:�L�K5-��@�_�k�u�#Ĥ���0�%@E{/��c���$M@�t����*,���a�`��]�{�"�Pham#��g���t�1\^%�M��h]/�å�<�҆��TB��znnz���ѹ��~oOiC1a�����.5J��V��y��_������]/�+�;%�f�2��wY��4�b�n<o86��m^�N�Fq��z�S�Yy�e-�7-fP/~�V�-�#&0Ҝ�q�&۷�'&%�-M�9�l`/�A{���O�>5{�y��~��w�5�a��g̹��?�����tnZY���W��L�v|�;�Vy�u�g�� ������̓� �7'��k}���Ǒ�t�vL���|��Ŗ��p�:�L;�(�Z�+�ڐ�o��78�՗4�&�����]�7�S��2\�)"�"Q���:fz镴/�.Yx���]"r*�Ex�|).I6.�e�:iNK��K�%C�Pk٫rh�3s�SJ�4V�����O�����_3��+V�}	��g�tj� KǮ�Q��tb[�5��d��W}��(�v1���MV��>��6�-(p]	�s��j�C� �v�r��ۙ�]~��0�VS"�)�"z�2��9[מ�Z������C��-xt��m��E�����d������yh.�5��n�LV����}y�% 76`q$�>^�#�>�ȕ�z����a�˒d98�p�kF]/-�3:2�*ن��*'F.?&1�j}�;�O�|���{�X3+�9{AG;��Y�Ң�.��a�v��q�Ωa��S�hs,Y�WNZ��t]I�0�ǑY�:.Q�܊}�ٗ�֭��>_Bȉ{��]!���������}'��Y����&zVR;�Τ��Y�/k��z��e��z)�Q�^��<g+��~)�!-d�SA��f%��WM�{�g�rθ���C1�bg?��?m�U�W���M#�x��	T���b���c�j��i^��&�}��({���Ao(К�VFӗ1�Ӽ�3�e6����0��|�P�>�!Ҍ�1�31��<f��DwW�r���xȨ�ㄜ�0��Ԉ�^,�|���B�=�'Ѿ�y�5��1^F�nv|f� ప5N�-�����v'D?,՞Bמ�x ,�7�e���n�:ʴo��H�o%������hO�mda�e��F�nT�|ǚ�+$B�پ�d�z�e�$z+�c=��ͦ^U��'0�8�O��9�X����Z��vD�k�N���w��p�/13Ǻ�O���`�D���j\��뙆�u�B�r�s�ghSqgԾ��d2+�cmx��Ė-q^�~f�:���}~��A>�g��h��*B�yTB��4p}(�ݽ��7�"�����+W���g�%�V?����Z{W��dxѢ����=��f�T�r�ͥ}r�g�b�=���n�;���/���� ���U�LI��O�9Z������y�4����v��L�S��f�5B�b����+R-aG��Cŉ�O�c���o���/�s��W콈�ыƼ��z��>8n�r���z�h��KW�C�n�^�������!���dN���sЕ��<���
���ͭ��:�!-tY@U���\��`����BT��cn��V��NY�C�ksy�{#L��f�����(�!u��`���R
�� ^k�mB^\�a��9��A��P�.�1��;�p�n�T,�m��fp��$�ӻ����1���_a�αv�{u�c�j�^% ��$q1�Gjq��;V�a�k2vKH�,Jй}7��_v�3BԖ�"t�߄��-[Z�F=n���V�ݱe��������Ԁ������&^�����X�rvO6�>ł�t%8�.缛؆�
�Iǒ \�g-�%�Y���K����d[i�M�(A�㼫2��&��S�$Է�wE�!՗��>�4����u��^m��P�0<�p19���PZāi�h�[��<Eԣ2#%���r��x��ۧ�h��ua>.u���B��s��o6����:��3t~�wG;w�h�:���9 VWU��:�,��������y	8�-;�7�&�l��5|�䣮:x���Z�^Hħ\.t�l\�������5Ҝ�	<M�x(\�Bg"7ݣE�p]ݾAp*u7f�][w��e�����`Ǹ5g�̃�����%
'���7+/�Ʋ��Z��j��}4e�7�v����зL���=(sw����n���2�E��U�kq^�)b�e(�>?S�,�Bc��]�������:�Ti���R7�%YO
79��$	�#��6�7dijK�óNlͅ��b����.�+Y�uIo����֨o�x�\�s��/�"iNZ1��--j)R���ҢȪe��,EEFED��

�E��1.4-���ab9�ELʤ1ƍ��LC��JX[k3-G`(\����LP�]PYs3!��q1%h$�RٍƘ\W*�,U��bYZ+h(�J�E�\���)l+-,d��[��]a�%���8���V��m�\j-�a�X�J�*��d���MU4ж�KJ��`�11�%T��Ub8���W~��ʞz�p�0�� ���MZ�W8,`S��nKE�()�c�j#��6��*9���	��B0(�S"�0�؛sٺ�56G��zh桂���f��*�f�2\�T�[{�φ	.���������0�)YJ&�Fʝ�ٶs;ZI�Q1*Q�c�S�)Z�*F�S>�'Zo����I���{%��E�W�#�)C���!��a�t]���gQ�5k�y|�)I���E�/��x�^�os��
�
lg���⌺j�"�����u�'�{�b׺yet���x�}����KOn&1�����ƶ�7�6���$��E�ۥ5>"��4_�W�q(�dk|]\�'��S���C��f����H,[jƠK�g3������OV�;���=�%�c�y��1ɮ�N��ȥ����a�U�J�tR��t�W�k�� �k�nR������.�&�=7b�)9 �sy�#ܬ��XG�;:f6/W��a��^�PZT=r{�{ciC=�
��ۃ~ʊj�F��sR�1�O�CĻ$�ו8�yx�@�ѣ�b��P1,�����fi�T_{����<���-}I#e����zM��i/U�ۜ�v�]�ا��B�}�G��V���MF�f�4����?c���T�D�l�JrNW���t��B�x�G�|��]t���"-�z\�],T)��R!W�f�@�&n�`�
c��l�`���\蓾@#u���3H�f��ﬡ�)��CMŧ'��5����^#lSI�;GݗY�� ���}�I�H�s��1�^Sߗ]�m�:�]��qM����pp�y���muʡW)N��w�c����\��m�\�X͂�#}�6%gJ��15��"٭r񖋐�$�rA���[kƂ\p�H�kN������qk��v׫�w�-��3��g�堻,ֈ�����PN�3�������Wy	8k���d��<űǼP�\����^�M8�����)��=��W2X�����PG�d�}S}}�lV���L�P�#�X~�v�f&�4F�^��ҋ)�eɚ�^u)r��J�&�����E`�F)�/^n�]�ַ�\nn�:Go�r��F5����m{�4�y��Xླྀs�=�M	}���C����g?��l���y��w��Z���\D?�<@��T���(����5RM�K�{�Z�
�.|P'��ӆ�8'=�_\}��|��XkQr�o��3/��p��vi@� 6�=o���q^��B��b+�N��H3!�}�����S+6�	W
��L�h�\K�܋�&���	9V�)�c�~��R�(�����<G��)��<2��ܼ�Ywެ6t�k�G	9��kZSSh^!
��d@
l�m�;f��6åq���j&���!���{�+�^�H/���Q�/yg���E���wV���5ڭ�\׽��Mrg�z�8���M�y����t1뻶���B��/��|����C"�*|�SF�q��ı����ǟ%�J=�o���{�� ��0�qC"����y�$��Ʈ�{o���ԁ>6`��{�7�ȇ<����/�m)R��QY�ziҗ�M����*x�ٸtf�ȔkΎeҙ«jv�N�Gǹ^������:�[�Q��զ����ts|&^]*���dXS+��Y+s-�S�\X��ސ�z�*����Ƨ\w.�F��/��T�#e'��1H�����أNc],����7���<�֒5W��B�	ӽO�t�<��8l��"�}L��ZK���I���絲&-ӆ�,��dq|�繂���_l/�"�@ґ|��Rdͺ3��j}~u'$Eғ#h�P:���Ykv���O��R�-���(��p�iY�
=�Q[��V4�1�J�!�-�yJb������R�B
Zr �����H:\;W쭕���ڹU�<ڸ�&�*9�s��H�.���{RW]Y^�u��Xn�?�
~4b��}��A��i|�hvO@bS=�ݗgԆr��m� _y�H��%(pI���K�r�d�U���:>CX�����?�A����C�[l{U%w����Y//���F�5KQ�]�qHnjz0�q�V	HR���F���L��oa��v�U���גÄ��<)G2'���7��S>�/S5\��P�6L�R��6��W�х��Cܑ�ZG����1�����\1m�gQӜ-�~@*�����{��n���d�<Zf�Wg��<�5��2��Ǜ���>}��u��m�돻5�K0�l�k<�����ą��g1����'Y��s���^X�*��Fj
xXk��0H.�f�i��BȜ8�o;�7<����*�s�.��O�#��iu�eg�v�}�F���s��ZC;|��/���t�UkaS����{�/�Z�(A�4�8�	5�-�x��5���Fg�w�ᚇ��^�~�wu�d��=\�g�����)�Wɲa��״�͌q�E���.�����P��YKL$�ʮ�#�mn��k�Lb�vsU8;GӇQ����k����p�[��E�[^[�W`*/Q���x���S^��zEW��S����`9�b��2��%g.�Q��N�a���T�,����eY���d��q����5��OR�C]1F�_�/{��g�����:�;���e��y� V��:wA�oS,Lˀ�/΋�9\^9�B��LZ��L��n!���Q9f{�.>���7>󲋵���"f�FŤx���/W��Rg�6xՄ8,I��T�s�{P�!9��7����*K�g���"�D3U�&{��N?.y�P�渕����M�٥nbMl��>*�ל��&k���eխ�=��e�ڑL�y֮>>>�����Ѱ����;+Z�õ��w^�����S$�⾼y�,���Ḱ$orZ�G/[VJ���e[�ʕ��͹s�Yк��tǮ��C����r6�����Z��,�<x���3P�G��~Bj�T��d�Xt��S3!�m���7j/�Gwu���!���!3<�y�	CUy/3n����.�����C�n!�63���1���7�j���c��1p	��Zp�g-Ղ�@�8v��C��uW��C��g����0R��U�@��d�^CƠ2[/�Ww��kւ0����)a'5�,�H����kƲf����zZ�VD>,�!��#Nj&��󾾺 ޅ��Reg��t�_Q��cǼ�g�k�H<w5��Y/�{ow�C�x�"��L�t�E��
���<��z�{N�<֝��*���m\��\�b��#-x���יy`��L�M2�W���;vH�EF����ʢ�ީ��U�T;��N�mhy�;S����r]��xVj���Mm��D�G�&��e,��x ���w�E��|V'�j��mgf�D�}K�'OL�㶂�b�"R�*�eR�{G�]�o�͞�����K�0^�+W���g�^"W)V����{�q��\��N:�Pj{����[g@R�}�oJ�}۸�+�XLVj��_�Q�/g7��r���k��(M�h��2���lڰsm�7�^���"5<��{��w��e~�8�Z}�^9�ܓc�5���_v�g�������E��������[�ʿ{:Z�O����Co:J�g�&��4B
=ԗB��T��ee^gD3���Y�C�h�09�C�ȲH�읩x\N�����jt��i[%�gz%SSe�+H%p|h�¹-��ǳ;N��ef�G1hss��2 Ti��εx��E�/y�rs݉.U�?LsS���W �䉎n��'jDe(�PF���Ij��(ʜ� �v���)�ux��7O�UO�������i�gz�����J��׈��&$�9��AwW6�z#%�3&qW�^CX�R�"#Vb��h��z����$=��53S.}�B��A��=yS�ޘ
��ҋ#A�3R;c^���=���G�X���U�מ>��(|@���x�������D���b�����
��v&U�Y���{^��ួY/���or�� xF�'%�J�C��^��<�6����Nc|:���MU^���i�l:Y�vQۣ�v9�ow��O�~������ڟ�j��4�(�9H��(������@>��ȽϿ!�Գ0���S:����]���`��<d$�@
� ��hXz	'���o�I�Բ^P�"~z�  u�I"2��0���K�g\~��63��YX+]�"f冐�1����ڷ�{2�c`�1C �QV��R�D�u{���/�Ae� � |� �N�bK3����N�`~kU��~��o��w��U݋�!#U��2�M����Fwx��D���k"���������Zp����K�vXm�h���a��eNsj�%́��$�  E� )|���UAE�O��M r:U	ΉL/_��%���6�-A��Q1l��%��4���m)��Fi�lI7?(vd&���S���<?���c�!�(��Ɇ����&V��7��T����bM� $��]� �.}��z�ג�-����7�j"��b���!���K�j�2<��B�*� M�E�{_4`���t�2]�`�	e@�p/*̪��b*��C�lȀ��/�� AZ�j\B�N��Q��	��PI��XB���mi��%$�Z_ �}�D	�oa�Ղ�S�D@@����
F�=�����vd����4�3��c�$����Wv<�xǊx�u5��r/��,�  n:�A�N�iܢ  o_Jx�q3��OC1=���3x�u�Z�j,L���0�i8�. z��7���=��|ˤY� ��2��D@@�l4�~�̓�[�Y/��̠�Z�RA�W}e�aP�� ��p$ (V�fh�<O,�mݐ���v�2�Ll��!�Z�fKy[�'��TȂ!���$���B��rE8P�겋e