BZh91AY&SYN��@��߀`q���"� ����b*                                            � HX �}���Ly�     �  ,      U         P           ��z�$��"�T(�P%(J*��J)%*)H)���$*JJ���D�H�(�� U>yH 5T� )Q
�����bԀ9��*���*�[��{�4^z �ΩAws�$���B=nl��w�D%��N^�(<���   7���64h ��o8:�|���*��{c��%L�_mJ�q)m�'�`>=�� tS� ܩ�������b g��� <  � ,���@� ^!I(UU""%R֢U l>}��gB{���}��` ||��
x 	/F��v��ϰ� ��|^ 	������   9��@ �Ի�� ���H�|} 7`�w� w`=y� s�>� <o�b�< $�=� ����� <�s�X �    w$� :�Q(�T���۪> ;��S��9��`/G ��jJG����{Ͼ��� }�=� <o���x Zǟ`y��   |�H  `^`9�=�sȥ< d�70��݀9�rt��x �cv�N��b   My�P 8�QQJ�*U)*J���l}P@�CBC� ���J��#Ҁ;�8�ݺR�w����w�* { ���  � ������8 C���x� ǐv 2 �w`ǽ�K��x�2@�!�   9{����$����Q*��/��� ���0C� ;��� g 4v :1 �ꂜ [� e � P/��>��|@# ��$��<@���Cv c�p �r r�n��� |      �  } 4�&�( FL@� �~	������ �4� =�M1*T 4    ��R&����#  щ�14 �H���S@44 F�h Ԥ�~�6���COQ������}��g����ߧ��~��k���O�-_\��{�}|y���C��^�1��T/�U"�Թ~�R!�ȿ����+���_��_��K�/��D5ӛm�����T�~���_V��������������_ɩɥ`�`�iGC���D�"q��j�f$�R�hhN4S�Jq�N0�)Ʃ8�Uƥ8Ś)��)8�`8�R��i'S���Ʈ1�q��b�'���'�fq����.58��8Ì�a�3K�8��aƪ�Uq���q��8�Y�\j8Ҹ�\j�2�0������+�Uƕƪ�*�J�ƕ�U�q�5WWWWWW����j�0�Uq��ÍaƎ4q���N4q�q�8Ía�l�Ǝ0�'8ʸ�Ǝ4q���3G8Ì�j�2q���d��Ǝ2q��N2q���jq���k1q���jq��N58��N58�q�jq��N2q��j�0�S�3.4���8�\aƎ1q��N1f�G�0�G���S�d̸��b�'�Ì����N5\e�8��d�'q���h�3K�8��N3�Y��d�'8�3*�Uq��8Íh�G\i�q��UƎ4�0�4fq�q�q�q����N4q�f��d�'q��ʸʸ�ƫ5\h�G8�Ǝ58�Ǝ58��'�l��S��a�U�.58��N58��'�efq��.4q��N58�Ƨ�jq��NMN2q��N58���d�J�K�Y�q��N1q��N2q���k2q��.58��8��8�Ƨ�k���Ƨ���N1q��\b�K���1q��\jq�Ɨ\iq�Ɨ��b�S�.58��N5Wq��.5\fb�S��e\iq���Ǝ58�1�N2\a�N58��S��ef��ƪ�'8ʸÍ+�8٪�Ì8ʸ�q��W���S�WW��U�r������+�+�+�UƜif��K�WWWW��2�4�2�5WWW�UƳ��4�2\i\iq��.2�2�5WW����Y��Uƪ�*�J�*�4fq�q�q�q��*�0�q��ʸҸҸ�q�q��q���\i\e\j�0�Fn5W��8Ҹ�q��3G.1\d���*�\j�h��\aq���q��EfD�Dq�UƩWR��GC�IƖd�1GG*��Uq���Hq�8�`��
�a+�U\j&sW������3^�O�}}o�Þ���k�.^��d��2�����v|ć��kk��Wd�8Ű�U��PN"�F��"�q���:�h��Ie�^��6��g+��c�Z�,�#;S�I8+'�P�{�;f�o��L��pI���!�zG� ߺN���Ţ�v+���:o'��Sfo��� "��f���ͭ6��&��p �=xb�k:��	\�ZH¤ś�9蚖��'$'7�3,`�F]��:X'G��-E����om:�׽��NH�� ��;i�̂.�˺���4 &4�w4=���B�c6�T2��ԳQ���w�]E�p�z�ՁwG�L�9>٢GJє�]���p�:�j_}���1�ŋQ��
2����&k�vP�݃�-�rӕ6owkoY9�6W�KqNX��#q/�=k��ɢ�8@�.���7ɻ�t:AF�����ݺ���,a;�I�B¹L�y�x;w�{�u}Zۚ����j�ˆ�V���ѿ�6�3_����Ț��_�8��gc"�Je����R�,Q�m6^{��Gy*��bb�x���"h�" ͚������6�Ʃ���Áϣ
�7bۏ�7����Ou�H��ܒ�ܺ��s��{]��зa�� !�Af7�'�xN��1C��q�N�e���Pv�V�t.O�N��386��w�7�bi%���H�4vtMi*�Sʾ]K��[��l�`kYc�7�`������wQp���l�ž5.�sE��uP��9�z$)ݻ;Ts���K�F;p֝���Ȝ9���G�|/�*۩H���5�u8+�ls�{ւz�(�"L�L$��@:�F��ww4Ֆ��1�F��5�����+|3P<�u�q��W;�s����4�t��hsR/5��o`�v�`�q��'�t&]�����w	^y�Atqty��vv&N���{��WWq��i��u����
��sHp���V^��4ؙ;���z>9��v��p��"�{�7ϾZ�;��&�]�	��YSD��wxoN�����aܒN�c�����\�ѽ���6ѧ��#����zǳ9��T4�������b����H��󱠉۸0��é��o|�P��{����v�ݸsSƻ���A�u���g`�75Ǔo��,;�ON1�y%rĹn\޽�Qr�.gC����nG���C�;p!���c睭!f��gO�S;R�եtk���V�����^}�"d��RZ�^t�F�Sygi=�Oa�4��D\tf�Œ9WN4;�浄G�l%Pn��$�ڮ�j����Be���}A���޹ېME�2��k��/a�F�0������s�haD��o.�qR�!��f̌�a|���2�Z��E��j{��[���f�g�j��{����4\�Hfe��Awx�g�훲iu��3�g�r���(L�S	yl���O4;�3��ч�ve�Ʀ��;n���9;�ya�wܯ$��p#�p�'�z,�]���OuG�l�9f��3@ă5c:G���c��{b�Ǽ����I��U�d��G�v�w2f�:������굄3Wp�z2o[�<d`�ڷ~�b�M�RqD�b�#��6�e�\�U6���Cк��{vӂ^C%���qnm��\���2�f�KJ�� t�&�v�x���S�5�W�2��|V�i3��\.��]�{���x����E��{�gc������v ����V��`4�t�W�Y�ѣ!�Ð�U�F��&n��,�7��4wT*]wWCN�w6�F -�q�M�a��S�b���A3�){����{�ɡD�>ʊ�/K��4�>x�ef�gGUE=��2N[��@8�&��z���ӎ�����y��ON���˥d��V�s�em���V���t>�חG`�ʣ�̿�¸1퍷F���D� �^�b�1���8�M�,����[o��U�&�k�c��^��[s��v ��#y�3n�
���w�ۅkq��Sz�r��t��ɣk:8a�NѢ>���y򷘝7�S3;,�8<m0Ob;��;�!�L�G��C(�Y�kз����; �#;/NwN��9 ��&"ν>{�2��B��a7"��l��O��������{q�+���𝷡T�Kp�8Y�yv!�"��0������!d��b���f�G ��v�y���Ëx�֘.��4�[mP�@ ��~g�G0��(`�w�i2*%���u�n,�d,e	giMÜA�c�f��'&5T�16�v�z�9�����F�]��o�ʠz�����!!6.�c��=l��	�NH�!��y԰沰*�5A�U2U�j�c�2%U���ڴG�n<޻��l�׈x��O�u�Hޓ��p嵵,���Z���'�Bx�*T�8yr1d��gv^|�SZ2���Ў�o;n]�M���'f	���1Qq�˚�����%��5g9����5΅��[��/�5N�uV�-�u�B���a��	9�`}������nm��p^ /�;2bj���eO�簐�=�p�n`bh����@r-�Yu�;էIP�ۜF�&�M$�͗�k2Y�ǭ�c���[^!����:�sP-N��Q��-8�}��Y��*�Q�s�|M�0�/����[]����/��X�wf�P��\ؗ咍:���5=;Z�� �7�� ٹ�K��8p}�LG��)�Ӥ"��hH�Z���׻���Qn.��p�	\���d;��_:�GʽѶ��He���ܹ:7��k�uC���*�<�����y�>��4K�p��u��X�i���샰��b�xn��תnZ�����)�ݪ�.�,�ű��z��8 &��ė�ަ2r,'�5vqӣ�4ݜ�3rO��\L'`F� ��j}9�ky�]j�}�ߎ�ى��Mg%��\<����c��n��q~%P�i�9a559�kJ�۹U@�8R,	2p��g^;5(!���������B����m)8nZ!��l�KV>h��ck���G$�5�,��ݵ�f��6
��5����D#��<k�����A��Z�� ��iU���\�	�ޣM룔����hro©����Z1�Ҙ���1����k�
��^�*�q�]2�µ���0%�m1W;r]���g�}.����λ����6�t��~}����ҷf�@��c�k|��+6���n��i���]ïoJ7���?n�l��y�S	��9�s��_��]����l�ָW�Zv�N�ډ��d�<cVϊЀ!��wA[��Qw�����0��	�+9!��������"�~\�^�3���q��}&G�v�������.ɏ�Y��0���JX���p|B��ro*����Q��t��Wn�s��zM�2��c�w�:���{5�kfN�B5n�����_@iµ靿"s��­�c�CI2@�vUc\��g��r��!�*���H������s`mo^�Wn�f��R�F���;X{w:G:G���c��VuLnB����\8F@�rަNv,�#���B�*�}4ռ��57T�c?�yn�Yk�N��7T2�۽��h�{��@�ø2�-�N꽝����� ���Or���Y.�ݛ�S.5?.ӛ��P�N�q�E��SpC�y�!�W����l<9��Q��3 �3N?����r0!Ap�>�>M�u�ؖ�.���,"z��`7��ɍE�����wA��&	fۓ��J6�ڀ�:�f$́��Q�jo#.�z:\��A�`i�]�j|"��;X�μ��Ɗ)�<8�=�S�N 1>k4�����P�y��ƾN�\�.���!�lh͗`�`�f�I�oek��H/�}���Е�;�R�a}�X��l
�K5�qt��#��e�<�d˃)�э���h�5y�����V��2n�Gbu'��K�P�h��\��m 92�h���H܇����-�m;��s������X�uK���J�zwp��Z�ͧ4��#`�����hsvޣ\W��8� F'v����Ro9�ٚ��G�p�Y�K�,#��.C���t���|�8����t^|����] `o�H�'��,I�O%�j����q;�d���sٝ`|K:���c����y�N����E{���ڳ�Hbа:`�K{�PgV\��~�X�W=�o�lnDswq��)ú�S����0C`c�j$`��V8S�grDc��&��K��L�qr��5:��jS7D��q���I�+l��(o�N:{z�+˹ӫ��b�o#|5�һ5��r3���ql�90fX�.��U�F��"z޽*Y;��-x�N��]�rC��R�6V0��o=;6f��L�Wf��s�%�АFM�!�Ǐю(M7����t�T��K#����52������S�־������xE"$�{�z*`],v��t�ư�	��Gbm�Wk�_��Gp�]�5��p��� ����D�ƗMe� ��d$'�3��o
�T���X7TɤR2c��+��ىtы�h��E��x��Z�����zrOpN��s9��}�ol:ƓwU�)���J�.�n��;G%�q+��,'�y�����8����sv��whE^|��Y��c��v�kSv��.N��v��Ҁ�5��[���xl�����sy�BI�%��g5�K��ȵ�� ��{ ���}+�$�b��c;�ܔ%ps !''&ΧnS&l���縎�I=�5�[��we���e�r��3�Y�u����sLX{&ֳ�AwD�@ �"�Թ��gW��g:ݗS'@��	�@�۱��\{5
7�%��������_ET}F( )n��yg6�xu�N�7:�q���6f�Q4�XiT�a(�p=�{4٪ryv��V��;'hO
z�Vy�-#X�#:���h�'�T4RD�JȈ֧uN���p9��x�E��H[6*)IQ��X�<w���!uɯ��0���v��/f!sw-N<��I=��6�4�쯭<H[W�3x�^�9�2f���� �u�4��q�,���5T.�˜���7�a#9DMS�4��k�s_�f増�W���)>L�x 0�欛�5S�z���Ӗ�<r�s\�������S�6��5=ך���S��ۃzz�;4GV-��E9Τf�u;���(wo-�4��b�Hޕaç�n��fr�Mʁ������١n���"�*�v��=n^�6»�q��)�n����ڒ#9{��l������o7V�2�=��S�stT���3� Y���;N��r:�;l�1nov��52�Q��F �nR�Z�5�։
�f�1�ޠpQ����od}&�]ݛ��7o$�XĮo=CKc�Ɔ	�5�lK�*����=�݊v��fE�HދOt���z֒OZɫ~Q��M��ӼF\]�]�	��j͸�����j<�8�X4��9��v�PQ�N��9�C:a8p���0���#�l[����H�l=0�q�y:.<�	�9-A�{υ�v�s�}���EDw�����[�p���T:8��5�H+hө��݈�47r!��u�˅RJ��q�q���@dM>+fE��v7�8m�pthDYױ.��W�wh�wd����͕�Ë+傳�5W��:��\�i��T�U���M)5>��#xAQ�U�VozE@�_	��͢�subw���x& z�#4��Dm�̏�7+����j�KwK�Vq�ブE����,މ'�T�ڱg��El����&�Hw�n%��d�I+��ꬹ0�Nު�k�;c��w\ݸ�kS��{�ݞ�݁f�����fC�q��}zv^ǲ��篁�ݜq:&�}�lc�����k�C��`����^Ĭ\1v�)�ŵY��Bv���!���<5��ƹ��Ǹ�ra�����c|��9ҹiu�����u�w)�M<��y�;;Ȓ�|"���X��ssv�̛�;@��3[xY���$�c@	~��f⯎���ι��~�nH�7���y�;<~�&W�f���i� ����_�5������ߧ�e.��a9A��>,$b��(=��,{vA�A�����(ѥmsR>����pT7,���Gx���Z��7�\Jy.�i@���7F�4���>���T�q} �v~'}�O%_���'n7�QJ��/t������1+ ۣ^S����i'e��c�x�VC!�~w[�X����}�H��}<J������v���(��&��2��*�0!��Cko��NA38���MD�{����W�+۸B�UԖ�V��1�K�H��|�t��i�N�k�i�l{�3f7�vf���N�i�c�<���~'sɆ��o�X�{I�&�+H���|�	��ɚ	�/8�����.iH�>��ʹ��?����T;�1��ޤ�ݒ���upiGv̀�o�E�\ѼL#"�+N
��y�z��	��� j��D$����{�z5.8�"�D]��Ű���ol�e��d�w5Ѧްn�	P_��Hnoo��|w.c�rv!2�9N�v0��J�^1^l��w��1��m8�MsFK�N~ۧk.�N�����{�o/�����`�U��W�*�n�ׯ#*�]��y'U��t�����{0��ר[��gv@��w��'�)�n=n�'��lg,Ny�kNn6�G�}�<'�h��HGsݘ!zȾ���t�hCE����� �P��������=�|[���� ��h���D~��bX ~�<�ԫi%�s1U̪橵R��̐��sJ�Em���j+�ĥ��+���l6ٲ"檮d��B��lJ�H�$���`�̥�G4����*V�VʶA�mRsT���-��eS����Kj2�撜Үh��Nh���aK�9�+jV�m&��Rؕl6���Vț*��m�W2�sJsIUU�Ske`�)[6I�M�l���V�V�Nd���9�mP櫚\Ҫm梮bU�@RB~�K�3��)�.�����<�������0b808�a��I�g�NiZu��O � �tx���h9�xd�+�P��q��8ߢ���#�N�]AHb�D4�LPȓ`p��8��� e��,eO#�LC`�HLeDغi��Zo^�߄��3T�BZ�g�5���<)�D���Y%9��#8��G�W�%y�e���D�:�141��c^�JI#K�̚p��M��x�sr�y�A�w�;���պ����)$�Ťb��\p��g�	��q4�����D�G�pa@�Q	5��2@�QS����6@>_*I��mM�f%&�)�����Y��������6W ��.t��Z�SL@&����K������ޑ�<^	0�刲Ƃ�|�̃+E#7<��b�u�MP�RI�^��u:�)�g� ���=��P�K+9���x׫�ʥB~�����*W�������4����"'�����?����o_����޸������e_�&��#ʐ�����`�(�W=!�g����s���c�k:���~��+>�`���C���{��xn�9OI�|}�7�Q�"�oor�mD�������=N�J�,�ugv�'��vEga<�����r�C~8�l�5"�z]�D��+��{����0t䖞���O)��[f����tM��`߫;���
���1Ȧ�d���&��p-��h�	�+�<Əg�\ꇥ���\�e(y�`Ŗr��{ҏ��5Wq�xyK{��v���Spc_MՒ�%wZ�&C(��V[�FP;��rQ�o��w�t�������u���d�Kg��s����������"s|;�׋��X��|��G�bK��FO�� ��av���f��	�����}����-�~���6-/�����;��v�74j���6{������m�Q�|[GT��{�u���+wx�q1�� �l�bs�J�^W7�ѐd�����xl�t�^wsü;��W�'G�Յ�q�uF��r�"0��_`���;�|�#w>�Qϳح?}컞��@2��`��y��Jd����L;���O��|�,%�<�aE���t�׬�9������*�OE��ϬW0�tŪ�����{/Vv�s��Fۅv�^���4_fz	ծ]�
w,�h������_�,=����C\�v'[�l.�oP�G�x�t�_|��}����}�믗]u�]|:뮽:뮺���]u��]u㮺뮾]u�u�]u�Ӯ���뮺���Y�]u�]u��뮺뮺�κ뮺뮾�g]u�_N����\u�]u�î��Ӯ���]u�]|�뮺���]u��]u�_��N�뮽:뮺�u�]u��]u�î��N�뮾u�u�]u����]u׎����u��뮺뮾]u׎�뎺뮺믶u�g]u�u�]u�~���_��8nOv�S�� 3�O|�$7��\^*dЮM~�x�gp��uz�8I��}�
��'����a���K&y���Ź��=� X�z����H�q�ք�|��}�k�{���S�<���\�Z�+�����]�罗ޙ������U���/ٞa{å��}O����<=4*:z�,u1���`wJ9�;� �g��&y�>�7��m'�{y��SR��㙞����ȓ_�Q:o.W_����/�n//dh���Y�/`�T>۰p�q}�X��&ŏP�ueP�E\�Ȣ����+3����Y���=�x� ͧ�%�6��w�1}�D�.[���׉{3l�c��<���\�iv}V̜�i�б��î7���}�%��:L��mf,Ա%bO�cᾨ`��'	�'x/I.��@6��P=~&�OP|���7������sϯ>��zd�}u.P�=�₳<6�p���Q�O%�F"������}����y�O��ߙ��:�4�ɜ���~�7R�;OP-�zV6�[��/�V��б��w4/�ﳜz��=%��@�o�מ�wx.�T{v7�򕩼ϻa��f�;ҳ���Ln�{uV���U��<��/��w�wr������s-�s���w&=뫖�����l|*���eaI��^輻R����;����}���z���>x�1�E�C������[ccccc`ln�뮺뮻:뮺뮺볮�뮺믷Y�]u�]u��:뮺믗]u㮺뮺�u�^:뮺���]u��]uק]u�_��u�]u��뮺뮺�vu�]u�]u��:뮺뮺볮�뮺뮻:볮�뮺�뮺뮺�κ뮺뮾�g]u�^�u�]|;:뮺믗]u㮺��]u�]|�:뮺���]u���Y��:��������ll�bX<�q~������!{[� #��_�k�`��q���Cˊ񙝼���Τ�O5Ž[�=�R��7� �W ;�ؾ�����#w�}�2dH�[:��x��=f����{��cF�����W�����'�I-�2M�?ٹ��^,I���{EE�e�|;V��z��̾�����_��77���x6ݜ�����A���W���߹IO��q�����2��s]�k�?z�wwe��.��0��bk�X���Ǚ�X�H��C�s�{�9����W�1��}�y�F�޼�p�ބ�&w���+�� Yd��x�N�)gz1�m~x����%昷!# ����q��Y�Po;����k�=ğc�Ʒ�K<;���oK�^o���-��6��=���1`2-������+U8��E�}'��q����>���l����
�,�x�Ƕ����o+�3�{��rύ��� ZP��<s��A�9�Z���;nk��V�yЅAP?v*��f��u_T ���+�mV�|/<�x�<9�wt��wMB�sO=<�Ҍ�e����z�����{V��>�wʿG��J�ؽݓә��'��0s�@��ً���t�PY}���TT_U�]�Ǐ�y�.͓����a���]L����EJ�=�R4j��3���������n�D�T61(�֪��Err�D����Fɾ~�Y�3�<8�_W����˛�7ytܨ{c�J� r��<P��zb��+@�ǵg�Jd�{9��)]��^�^��@&�����-7ں�M�����Uqz�s�/Ҝg؟{�@Ϥ'7U#����{ΖN������{������n +�����G���&�jXơ���S�&i<�=H�܉��K��;�vk>�����r��鏟���⨋�/`���=������p�d;�Q{���&M�j&��'�����P���Ѵ�{5�s����N�����Ouv���γ+9��+�b�3�{zOP ޴��� ��:�og���}���4�����}s��~ªSt϶��`�5��ڢؖ8����������ӯۿӼ~���J��V�#�|+���ϰ˚G�������ܺ���5F���vi���4]�%�[={�*�G��A ����(]�~��A*�ϨZ|.�A�j��7E��z,�&����o~�]ۯ�L�8��{���Gǆ��Ӧ��o!&���_��hE��p9��m3��<�h^�ehw�V��;�D� ٻ|�Q���v��։bl���鼹�zl zW�_�eE��R�����>��|yE��{G�q��>�n=�i�.{�s'�p�w�'�wC/+1N1��D�/[1����g�}��B2g�K��2��jz�F��O�D>,�n8����"L����O8�j�$�u�}v�F��>��uG˺�Z�8w�f�(g#��,j?�&������y�[b�g=�W9X��̽��v�]�nq��D��}��ַq���}�=�#�;1k��!�����z$E���a���8�E�y�]3{}�9�>Aq���x{ڶ��s�7�f��|J��	��Q�����D�lڻC)�����^M
�'ύdg�����#�2/v���@�X��h���y<)ܻݏ7�;��˾W�C�x`�;�?,ѓ���r��X��\��x
R5�s��t�]����%ܭؓH�DSP����=n�*��7/6R�{ �c���N���=/x����������a@fS�sP�:��ܲ�p>��זw�&�ɡ�8��@�L�EǲN+ӊ��Nwz{������9�u^�=��F�_v�1�K�N��ɛ��&�/^´z߻ï�70�wҞ(�g������Λ�K�{,�|��gǎY\Ϩ���C�~��\�^9��ٴe���+���hq��OtGs�I�;/��!m`�������}�E�@b�GV,�&��� �=_�|D���3;u��+��>���^L�M�l��r�vx�4�yxL�9�/+��iB�:M�}_99���x*�&KI�"�N�w�g�Ou_ty�p�'�{=��{�K�U�G]�,+ȓB�ފž�m8�|��u������5�s�4PQ�{����~:�6:���C+=����'^�1��_jsl��{�<T̾�xY�Z����%��t`�4�@N=7��C�0>[�,�M��_��y��4��9�|N��)��S'��c�xnz�������,I<�5�9�jo:'s1-ޑzD���S��Ü��5���:���g��4���G��$�_����*V���A�{��k�яԡ �����lh<�/�s���+��\)��{9���9g�{��P�h�}�r߼�o֬��[�g��w�ح Wݩa��Ә��f�ݽ����t�ά��كg /Qu��؉ �zG���k{�ݪp�]�Y�gڲ��f�s}�d�}��h����E������fO\��ݥ���y���1Wﮨi�q��F�M8���U���^��Սn����ߢϖN����ɕzn��iߧm��u��`j}��%�b�}��舷}����;;#���6ǭ�Y;��{��՚�����ƅ���Sm��d�boSs����^x2�|D��ojω�N�6_bK7�(�泜w���n-��y�=7���݈�����xd�"O��<�۾���T1�I�=���[��^�F�0<s���sR����Oð����<��=�����Oq??Q�ܬ�Ozq:�z�wb�{�?u����(�0���on�}���/^����u�����U�Pǽ7�qZ�9��Y�Z><=����9��O/wK���zL�vL���w���A��D�k�/m^쏼I�f�n�[7����o�<׶t�{|;Z�}4��p����ͺ˼�{�,3��BRU�k߬ެ�w������V�#r�l,�to�S�����p��U����^M\c����n��|~��ojo~JK}�=�ս��b,b�vu����ќ��w��.�;ݣ�TerzK��G��,Rr�A� �˕�0�����oF�f�P�[�ֽ�[�d��>�wf۳z�6{�"AK�b^'~�bS��{�"�3;��s��%�r��B��3�;���Ff ���#3!E���a{t���=���z��Y��:g�L�p�7����_�v,���%�Ǆy�;U��o��u�8c{����l �x�.�m>%j�Z�o�/N��o����仔k�3�҃��]r��l���Po@y�v�М��u�" .���X��g���\��>/�I��|ǱM��wސ��r��f˝���/��� ��H�5S�M�O����u	Kǧ��������<�(�#m�]�i�O� '<�����V9#�O�k��S���K���)��E�M	����#���+\c��V.'I�^h��"�vkX| �����A��~�v8=��C�{�����{�wsש����/u�*a��p��'g����\������9��xD���Jq����*o�غ���K��r�>,{p��^)Ƿ�`����ٕ{�״�$��#�P��1�Q�8�Za�=�������2��^��{�p��3�+f�|�իԟ����7��p6�Q�q�%���̽�8��1r�~�s�>�$ͺUk��G��`H���(6�7ܸ�7�n5���8��A��~=۷A��������r`ժ���xEk�<���z�D��%_�r/0��k��3�'����J��IJ��%�~�t��C�a�.��I=����Rϟaq��#9Ύ�S�[�aA�U�� �l�{�N��z@����8�f8۝ �;#�l��I��w3��ԓ�zz��@K��.��{�]}����}3Г�s�� ��}y$�{=ޅ.�*������rL�#9N~��c+� ����Iv<ݣk�K7=G���վ��g�-�>Kw=�{n{�-���g h��j���^35�Ʋ�ٍ�儮g�fjz�����X6�����G&Mzj�D����rC<�t�ޞ��ɾh���B�x}�z�{ܭ�{Z�GH#�ڻ�;�=�?�]{�2�of�D��
j��_%����v���N��s$þV�1$�N�,^��{\�м>ӻ�����Wu�?_O�ꌧ��UL���nc{nZ�`!��0a������=#�����$#�yа��b�}P��{ogaw{N����Ĕ@<��v_]���B���2�g��\�a��:�\��ly�ӆB.�����7tikV-Dd!z ��JXR�x���� |�D�y��O!��Q$������O���q�i�ؾ�{�*�g��>�>+���N��O=��o�w�p�z1����}���`�[���V��q��'��ڥ� ��Ò�ζ����g,d˯�	5są0�z��U�ՠ��:�ϥ靾GU:c������a�y�|�>��漧p������װeݩ�{�^ޅd�L�zn��������F�i/d����	}��{���9����ץ���]���_^!�b���b�+W�n7H�X���g}���$��3�ycx�t��1Ŏ��p��/Ϧi��2�>��9���a�wq��>�kxf��\7bZ)Ѽ��ɘ�f�{l��{G��z�����!�7�{�<|Mk���O[�þ�"]'�Ek������Zucr��Q/l�{�<�8��}�C���'�`��C�H�U��R�oy��Y�W��GT���7�"�91��G�ҧ��#_	<�Mٗzᛨ�#��!��֦��T�t�anz�hk�/�����/��G��|��Y�^C��t�AJ�=�6�/{����`0�7��1�r�fgZr�k���xyE�ZhԯT��KS3�BA}�����w�;�ϳ���sx����}u���;�wݱ�wOxM{'��J�b�\n�}p�f3�:�ӱ�
�3r�}���w���#�eHB�\�7_[�z5�7T}��P�nh��y�����(���_�����������>!��{�4<w.���\�+�\�Ok�V�9���$��s���6i�=�O�l2d�v���[<��f�<�'ӫ*��f��9�Q܆��[B�ΐq��.N��x����������]l�����ma������n��[��?aIm�,��2�,±ո�P��A��6d��ˣ�y!��U��[�����CK�{>ř?�����35��W��w��g�������H�o�ח��_�����x����2e�o.���ч�� ���*d1��Ċ'�>պ����-YGQ̭�aaj2fʑ�]��i�.x���K����/�6����*M�nf!�	��3L�Z��g:����b�\�pM3,5����c�t�]t��f�(��m+f

Yc�$f&�M��-�̱�!8e���k+F2��-�U�¬�1t]D�ΉH�
���I-��F��i�6��؀,��%��C�l�@Ѝ�ѣ��Ƌja/k)0]���\�j�� �,+�Ds^!��9v͔U����se�����֤E��!FJ(e�^\�afm���L�`%�`У�1.�����2Y�b�������EFۡ�H�]��t��˒]z���*Mnݢ�iD�M���Xa�G)c��R���Q8X�D�kI�cYK��1]*��j���k��h��h(WA�ƺl�*[!iB5)Jĸ�ۣ�f�a[JFŗQ*i5����D�s�f��K���2��p�Z�����1��E���e�+m������+��,�c �֩H0q�doin�m6�-	pZ�,e��V�[��H6Uۓ1����m.4ҭty&%Md�e!��u+^���PtX.��\ꌰvu��W%�F�\JV+�V�\�i�"�Ͱ��m���6/,2����3���Q�1
K�@{6kp͗(��]��P�m�-��0��tv�0���ݜ��U͉�V�)�9�k���It4-,&�lrL�[�R�v�p�c[4a��uE ��X��,*�
6[^*jWe�����X���U��)Ymt9���M
���IJ����
 ��U���*\c��+eF�;Z�8�cs�yIE��Mk��3M21��7JK)�-"�A������f3���+4c���l�uf]�e s��7qrss�F� �v3\�p9�(͵c��!ĥ�Yt��T�(캂&&�lq&&�s�n[�΅��ѬtrQ�2g;�Cl��#��� c��6�I��(i�VY�`"mE)dH��n��붧	���dUȥ*�+1%(@���d݌sA��{K��k�Hd����v�S5���Ym�U��˔�l�.��z#B]�SVeD*@�G�輨v�U��X	1K�J�.Y��CY�EIkfL��C]�lH�q�)au��6�08��a v%�^,5������j��=@�.fj��ւĈ6�ژ�{j�	6q2%1�s)��D��[���(�gv��L;+��fjL�9���2]*eU�ڹ��3"�؋�m�Y��"�m��l�s"��z��3N�(QٖH��P�CL4������x�9���(C�Kf{F�v#�\8��$�T�W���]g�"�Z,m���jcA��!+YIt%;B��5��Ԕ�[��0U�V̅n�8�h�C� ��(\%j]�Κh�J(4��H[�l�Mc��Z�b����4f�MI�)b7D���[�Mn�L����h�pԷ�&�����q.-Q�Mvn��{)�ݓmqH�[F��tn�mĽC���PѤ�1h(��\�F�Ɩ`sI�t#c��fѪ�s�,�iڅ*�X���i4H����7nb4Mr�uLK��y�l�0��V2��6���76c�&��ֹ���[Pѱ:��u�0��LM*��[XČ��4�0�hl�^���0B�5�d���WJ�f5�5\d���Cs�ͻ+�F�Ռ�ыEմ���ι�L�g���Ƙ{T��Ԭ*J�mHi4�3.�H�.8t���#m�iָM�A��.�t��kL�Źe�8(@�-�GW֦�ư ���A��q3�uУU2���묡0lQ��L�[6iC;2��D�{p����p�%IT�A-�q-��0����ɻCh.#ĵ��+�`�n�UMY�'�-�9��]]���rL'4u�����T�DH�a����t�pba�.3tX8�ɦc6kz��L�9�.c��%�	�����ٗC[���M�!6�uX�� bb�s�K�Y�^�i�&K c��+�,�Q�7��4%�4��H�j�W\,i(`P^%v���eQd�,1�oi�$�5�T.����X9J;�4�Ψ%� :��&�	�cd� E�����M\"\�XD�R\r@-5��M��m�6D�2�@�ً���&YX���Z�7]ְT�e�vr�M��m��F�ݑ�F��eu4e0,([l1�ݘ鶊��v��[�8��C40���E�L�Dh�2����LѕYv`�����`Bֳ:L����զ��u*KK��Ҥͱ�5�F&2d��It	t�2�)������LE�x�)-Β�YMtJr�� ˅��M�X.�fSX)���Xl����R9MQ.�ݢJu�U	��.���f� {6�ٱnQ!jЎ�����eu����[nɄ޻GL�an����j^ɶ���-{6� *�&`6�:��mFnř�6�2�Yu��m.+á`s�P�4��t6p�si��.��S�\�P5��GXe�\BRf;G%#,v��vV\��2�Ck[2��ŮӃ)�镳G\��c��c�"�U �]6He��鐙�am�Ε�
��]�9�j�-�e&lu���N!-��"��A-��Lb��-�5.#
q�`���\h�3X�՗J*\4��ٺ����u���,��lJKÉ[�U^�`Z�f<+ ���ئ�a
�cf������V:�B]n%ZY�@�!���R�H�*��0����l�R�Yt&���Lķ8�U�V��k3�^��Q�VPXM��L��5��&��W�),n�Ќ�⣭5��^FB����\k�aꄍ��Ŏ�t%\�Ґ
b$.WL�Ml(��њ����@�F�us��YST���l]�b��9�ĺ�bQ�ݜх�+M�Z��U�ŗkv��ZJnl�m�b0لA��If�*YJSkZ�	�HN�❩B)�f$1�X����E�e[-�8�P�f��LLLal!����c!����W[���.��(�chZi��z�v�B�P0�\�Z5��.u�k��(�����&h�����[]͡A�W�̣il�hGmSr��x�3C��)�V,:�ق�^Ca��2[hL\���GX�s�!��mlm����7MR�I�um��e��6&�+[B�Y�q�ĳ��&E�EM��$���as�[i��ui],h�]f��de5e�A�
��Ri��¤��]rI���M���K�+�m�͘(KdJ:M���ƭ]�6�l;:3X7jF5��!�q�W5e��i���SMY���0K�V�;-���m�t��qf��Ik�V���v��k��ub����4)(��5�Ux���J�mW�g���x�a,0]nYcN�d+r���.����ԁ�Z[�ʂ��etX	��n�D�"�hL��F���͂�^k4a�`G.�͸�uI�]#�h���x\�.�;D����i�M�aq�],fR�҂�7%MV�Ɇ�����e��6nĵ��8u9�@Ι*&��θ;m2��B�[�P�%b�KqK)�F8ã0�8^��r�kr�m��0������H����8�9� (��Ic[��k�밂-�ƅ)�n�F[p� ���
ݲA%�ؚX���ė���b�����8�kT�	�k5��u��֊
6J�$:�-��4z�X�]m֜�5���-�5���;R��1��$\�jئ�4(��nڡ��L�y٣�#]E5fns��{]��TfH�5�h��- .h���aD� ˴�5����s�0Wj+R�X:�M�l����G\M.�	�l�4�[fX�.9��m�C@R�Ů"$��R��9�:ʖ����3sF*s�`mQq#Qʶk.5vwZ+v��
�],E�U�u:��amR�����ؙ(�L9�I���Ʊ�229fibb塹3M��x�yP��M#4s��ɖf�f���"�b���B�51[�,rcs)� Ƃ�Ř�umEa�kb�bR<S�f��ƍ4!!�Mc�5
]](1X77h�d�4���)���K��IR�mm�1R��-Z�pck-#s͗@�CX�Ȉ����R�BR�6�@3F�`n�&�[���Vʚ�h�ʖkM�� �bTѭ`�X�ܛ$��rRi�$׀�����	f �Ɣ�F�Ch��+�^�8ܮNV�L�D�3M3�3�������8���(���+k*�K(��`�������%�\�)���v��"/�U6��suMs���6V�`2�09�F\�c4�a�b���)w]ڱ� m�"�kR�^��RQ`�ՠ켐�Y��@њUnlԫl��ѵ�`]�ޖW�pkV��h�[ st04u�VV�f��&p"�nQ$��m���",�X3i
A�f*�J܆e���MWj�h8eʪ���X�l�2���s6[-��7D�3*��c�#�[��ڳ*��L�K���Rݫ�`�UvUUUUUUUUUX�����֐M�Sy�'��&�wC71��1m�f%�q��m��y�7��(� �\3�w{pD��㸰�`V�ZLJ���1*�³2�*��`ns��.\���nc[�sǧ�}?����_n�뮺�κ뮺�|V�77͜�9��.&e��m��\�����9s��\Ͷ��χ����u��ۮ�뮺볮�뮾>u�gίXP分["�1�
��b��-s.0�+F��.R)Z�)*�`��ƈ��ċ�70���r��ąAf$+1*���"�E,�Uyn428���0YRQ��IX[`�\�X��R
�`��P�Z�ŭ[e*��l\AVEm�̅m�0#������T��T�R��
|�q���QU`�UJ�(R��v�.UrԂ�
�ܥ\AE���²�Ҋ)�-��f��8�m���^�ω"Ig6'��)f��d2�%eH�\ۦ�v�
��Yz�^a�^�NHw�G�F�kN&��J���9��]:w�a�~��0���6��&-��al.�e�C^�4�ue6N�L:5�К�ДCB�e��j4׆��"WƱ��԰�a�F[y�b0n�.�\;ƅLm�\�64ie��ԺP{]��m,�CRP��1�� &��Y��F��輳3�-�m �:���e�宫�ijM��ʌ�s�����Y��k��T��Tn����F�- :Y�6l�j�]��	v�����c����"�ճ�r�*i��G[�d4�=q���K0�Z$�,���z�1�U�j����Z�ۓ'Wul�i*�r�˷�Ci�Q�˱�A��HikN�-��)�&Kn�F�aRk�Z�t�,].!(WB���x$g��n���$��
ƶ(j�L���q4ՙ���9K0�j5+�@�6�0�F\P�k�hƹ�bEsԚ��jZ�i]�Y����,6�ɛ�B�A4�n5t�Z��W:
R��^�vI����)��b�&��/e�6�8ݔ�L�@�)�p�$��(�Y�C�Z�ly��@e�L�k��E,,`�AP�v�F���-i�QtM�kV�� T�h�P{�DT�hZv��s%�L,m������ܳe.�
e��2�"ԥ��Lێk����v�i��ե�m1.�1D��Uff�X�9�]-斸��P���g��!�%�\�(���6&\K\[V0��������l]�s�J�-��Z%	�J�Z��
n�����P�ĳ0�d�̽M(�#㈊0Wm��r]jƵ�)1�(l3"�J��J�v�3]i��oX\�U+��2��nWF,����H�#Y���Y�͕��D$E$cT�1��I���a�k�s�sf�3����P{Bm(��]���46˫�ʪ��R���7T��1�l!&�M��*ۖ�X�*RѨ�K[X(����F2�V[R�Zƨ����D�	V�T�RƔI`�j��u%j�yZ(�!�*�Nl-V��h�c!ר-YT�0���x��)K�#D`u��%%ZVR��P����j�H����6��6��֒�T�EZ�%�*�j��c-�,9�eX�m����}���2�~I�E�Ă��`���N�� ����}�����(�/YW����>?�A@�z�]��4�1�٦��H�ڜc@`�^֯4Q��r߀����I�x�AzY�`��� �~����͘g+b�[� �;�����������^�ι�)�c#��!ުZl�N�촒�6�\<�5�-��h	8�&$�%'�B����v%� � ��x ܬ;�Dx�%��fI.�\nАK{� �;�h���}C,A�ˌIB���ٍ`�,��c\���stu�
���]F���5���ew�篞��3��nm�d�g!�Q$�A��Te���7��  W�&	0����1�����_�����k(��0�,Zf�P��o����,I�Ԁ��>F?�D�g�`��N��4ĥ�O�S�����|-�� �Ή,	�网,	$�x$i�<K�{Jfԋ���>5�
N�(xnz�  HU��,K&U����ٳ6#�햒A����P+Vit��"]@�l����{��^�^�L�k�ɨ�@�d���HFň��"T
%ij�p$����
�њ�<���6�g�sw�ZC\cs$H�w-�Ę���g���O����Xe�}O�)��$%4�6Ͱ�.���WDE���5Ֆܙ_�����r����ĒK{o �I/��m���<�*V���h{.jD�A��MQĄ2� �o���[��& '$�7⺸� 
b�������y7�J�֯)��m��X}����B�m<q�1�����A�}��;/��9�TK��h��l�<�3.Ç<W��VIl�W�wc遗�m�Nu[b��%!W�7�7�v"�<�����,Y�b���	�	$�^ϲ�]�aXJ8���n~��3��j�\�%��.e�2Gg6Y>�e�T�ۜ*���v7|8� "��]�`#ѹU���
_#=Y�h/��H$β`�����<� �/��`�HK3e��E�\�W�ꀃ��U۶�rhK�9�4U���;�h�s��"m�H�(�e4�$�r%�Ü�.%W�S���n�H��'�zY��lLx��x��d�/b�N�8E�P�|H&2.dr��كA�bD��]˜w��}%�j��!���ҧ���yr0�]��@��䡝���,N�Ƒ-2C���������g/.��~�0Uzd�s[�H's_0K��{�J!�f�֭�]z�>�W��r�{���Y3���9 =.�玾�W�hK`2p}��"�����DK�ŕ9�S��b[QM��W��)Ѕ �25�K�˗$�v�����˴��l�PE��%���%�n�b������G�W�-�Mx12�.�<\�uҍ���{B���$ȭ�;k>��.	� �@�Y�b@>����F�$�Q�S�3r��݁,H�j��'0
�b��Lf��ݵ
0;��>��I�I�e����;��C��)�m���Yyu[ri�G���B!DAynK�����u(�G��'׌bM�m	bN�1-STI��0�b�"��eY������~�rH2�g���3j�j}�׷�S-,�3Ide�^D;�n�	o2L]��c^_�/W!�>��g5�� �o����y~t](/���td(=H�}/�~�=r��_|�����A{]<�h�sW��f����{�٧���m�罾��B��*D�9� +5,^`��&����#�n�B�I���&]��<6%Š��c��̹ˍ�n���f�ʎn�V5�g$�W�]����.�d!7a��L7��0�M�q��jĭe�4��l��bU�%�.�-VٲY��� �����Ҏ&8�K�IXV�8�k,pTMs����e�]���y�ƵI	�J�Mh�\��b'e���&Кm�MGL^Z�2���Yl��p�[Zi��jL�����v�iF�*��g Vm��٢�V�[�#�2Ł��"Cou0�Ep8��!� ��p ��Y{�	/�ǔjI:�L��>�r���K��1�ڟK)�\;��.�?�*�@$Y��!K{�r4*�p�o���9F��;���`��r�>k�x�A��IM��ԯ�^z��`H$����gci�[����u�å�3�	���r�h�7��	��U��h���^�����UK��� �CL�k�ر$�̗��jR�2�< �	v� ���,q��)^W�2r����lXu��>˥�bĎ�\��Av�F�v��f�ef+�*E3I�����?M�3`=�g��́,_.�I�Ad<j��}r�k}����q=W�M���.
0`@/������?�K~ЕG�⮝���x��$#�0pә4|w�DV"6!P�Ř	�;��J3�c�/�7�޺�����g�p����]�ѥ��dŋ�/n�2�|��1$�w��bM�x��^�ckTB�0T(PǍ���\�Q��&ߑ���e1%�n!��p��K�'l
��aҀ�Fk^�wR�c�x9ɹ� z��b}/��	c���=�}|�c��޹��w� ��D(�/!�:�R	nۉQ�Pݪ�j�M�l�$d�C�!栈9��r��2���`?��-�Io7���\�l<�
,�EX�ͱ5�K��J��i�)c�[Uc�;�� ��Ȯ�&@�N:�Rƙ2,f�f�\/��2	#���I� [��W�h�dbL��w��Lo��{ʵ �*X[R�Hd�c�bv�	ݷ��Hk緰q{����hs���V�6 LO`�ǬX0g_Ɍu^����sVپ���Q9�}qY�s�C�]ڵh�p|񯼆�j�h�3a>u(�nj�����8�Ã~���uo��^� � �;��!��g��'q I���Q5�R$���l�x �X�n4��e��}��� ��fk	�x��&�O�����?�����[��$��^�i�Q��%�-m���J���}����M�S�Z�
FgG4\6�,��Z�m��¥I��<N��/!�&����j��e��31��$�}���P��el)֫�B�gM����m��6�?~�@e˾���C~<��0�K-�a fs5�h��;S�(������ph����4O��(��r��2�P�w�(��;$ĕ�r$�F��/���.͸��%�m��7"\�#Շ��� ��}�;����ٙEF���}����@���؉�͙�X�-�d`�or�p�m�|9�~�v����ܲ;���۴&r��}
���p{������E���$�tt3�[�Q�ߏ�c'�_s�h,9�}�/�&��v�n�w�fd �����.۴�}~ o����l� ٱ��h�P����ߜ����f��مڍXR+�lI��̚��7S,������m��{3�,M6����qǘ�U�i���e˼K��y
Lf�1$>��INc�� � ������$�O>UA��{�O���` �l��M��	)�Pާ�k��r�+<[T2�'��&u�Cnv$�Z�<�>������o���8_�2	5��$�-��@���'�$�n}���[Ηݜac^)�A�ٖi�&΁����	$�u�q�nM�E<� �T����ө�xqIx5�k/�$��B�\N�a�.�4x���m�H�,��NȐAc�����/1d�X�u����ω��s�2<�zp�����$O�^���Pn2�H����g��Nt�k�[��N��;�g1_���N�g�=�<���1m-�$\{�:�����Z��V��l*U���X�X�י��.��͚3XcL��R�+^fr��Z�+�ֳ=sјq-��Z�IYm���x
����ړ���t{%tݒX�iNmbs�����SR�Ձ,�]Y�ю����-c1nev��kW)X�Z��kB�R��Ʊ�3M[�][K*��	����A�&LV#��d��s1VaISS��Y�ن#�pm���d-Ֆ*h]�6.������їy����A�6�X����Ғ4�����Z����H$x8��x��w�k]��#7{�ln_rک�����Ic�׆$�Q+��oL^F�8�H&�d�L�j��׆��}��Ӏ����j�d�b�9�P�b�4]F���- ��x&�i��g�%5���o^��j�v�$�X�o���K�ȕY��׶8S3�xr�|�=۹3J�m9~�6*���}qxg/F^?�q3�%��nZA&�^,|�!�-.�ѵrb���Z�@-Kl�꧳@�у]�bb]�16�;�3M�&�f;h&F�^��(^��亂�	x5��=�3��� ��`��c򏖃l�L�wq�oD-���BP�q@�ϢK	�O~�'Hp��ﲝx���[� �)���ͯ����g��mI�}�z1 ����m�i�pHn�r!0�Υ�G��,X��W�S4��}x�%�nZ|�����y� �:x��%��@��w����5�Y���o=����&�m�R�}���0_r� ^����?|�O B"��3���zI�nE���fy��!	�.� ��["b�E<�ﲱ�O��X�	��6��� ��T�̻ �:��(G���ڮg^�[1�-���H��!��"L�r�.��,NK'/�ڮU�S6֩�
�r�aF�9خ#-e�l�ͨ+��������Ւ�	=��|��9�$�v��&����=Y��	/�s.�(]��P�� ����|0?͇X��/@�A!��e� _wdH���o������=��{�K�q�S)r���9�-�����
0��O��=��h鐸���<c����f�7� �v�Cu��G*m���������������/݋�ݱ�>�WH���2��fz�;Z+vk��wiĶ0�_4�J��%ʼ�rq�`l닩P�����1oC:�)�O3s�h�nv��{�Gy�6��������m�cp�_9��$�/���_pλ�;6���? �ݜ�+��x]���湱���V�3F��C��،���<����Y��!����X�ls�Fi���-uļ_u�|���#���J8M�n�,���b�=*�6���b3��f���$�����e� }��bF1��<����f�>�	�t�g�=��G��n{X�s�6�/���X��\�e�=n��i�{��!;�����N���I�sx�G�nq�F-��.�#7��u��Fow!}ē�����U��zn���ܤ��(�Ì��R�<&V�u���V{f	�y�;ǔ#{f�=wfӷw��K�th�6���lA��o$	�߆��9���3{�_P����p�'���x�;�o�b�����B�^�����F��<��~1����A��yf��{p����$��u�s�Z�)2"'v���2Q|sW��n���Z.<Y�g�z�<�2��W� ��5̀{��:n�ۘ<!e�oB+�Nb�8|��$��k:��[�.}�����9���A�}˅V�0m��q�K�ǥ�Z�ⷖ<<��d�)�Bt5�����N �f7�q0���R���q-D��/O�]{u��oooooooon��o���;�n����� D�����S0�H��0

 �_&Zp[��&�tk^hY�[.��t�yz7�:�Z��Jt���������gۮ�뮽���=����͛8>���J�4I��*!��{�e	�&*�bKK+ZbB�eF�-d�,��R�`+�u��^�n��a�R߳�X�ZLk>����:���pQ�
�	q�h����`��h�y�W7"��e#��GR���28�[L�����f��ئ�T�h��)mŭ\�`���N����	x,� \b����¹dR�=���׈T��T,�����:ҵWSb�����0.U�LKJ��wuPf
Rĉ](�*�U�-�!����������m��h��
�%LkZVX��C#+Ɖ0I�D�9.X����e(�Jśj�j�@�^45���,��X��r�3)��Cp�5�2�3l̠���gv����1��+QE��P�)��GiQbj�lA���q̻�1���1��(�m��N<pc�����WQ��=fٳ%�X���s|�!�5����-7��C��H.$+����N��R��O�n��s(0� ^��Yw����8M�>���~s񋚹c�����O�[>ur�̹$�,��w�Rw,1&
Ԉ�����'x~�����u��(�>s���7��4���vw������r�%�Ad)i��n��
���/~g�\{�������R�����:��@�y��>>&���5r�4����׬�4��[�O�el�*���Y���!������ͺ�b���\G��&�e�ΰB�.m���Q��5�a]��{�������n�?��>G|��a��T+%�3����A`v��C.}��Hq��w�{�����O�&�O��{�;�A��,3���8E:0*Sy��}�3&l��xy�����5\�v������3󏼽z���{�P�Oc�2$�7�>�Ru�Id�!a3��Dj " LY��Y����Q�����t >"�T>�c��sE�{�C��=���9�Y
[;*A����ؐ�(����緿^p�����wHz�,��YS=��xE�P�%B�/￷Xr$�����󽿿M�WM�L�H��aS�{�"���^v�i�Y��`���4�,���zd1=+���?F��n�:5!ZY�d�w� @g����r����4�̏�rt��#'�~`����~�.]t3{=o�{݀����i����?z�S9>x|{p��,�2b�E��{�!�XB��#4�:����Sі0��8�P�%M���'A��!?|��}����cY���8$'}��jB0dϟ���Oy����<d̷g)�)9��w�A�TճG�f�2�^��7� ;ZƗs6�rA�
h��>O�~qfh�3o�H~k߻���!Kd,�3}��5�B���Xh��{���
"�`h��Y�=�b[ #s��(2T+%B�>���a�IXS��ɟ[����='�<aS?y�@��T+'GFwC����D�h�L�Qg,!
����=��ć��+!m7���U&`J!�4��;f?��u��dG�`T�����������@��}�8�D
�(T�M���!�:���a lnW�L�ln}����m�"V%V~��8� �+!FV����@�u�c�{����r����Y�,=�K�qf?�f3�%�f!���׌%l(��w�|��c��Ę�~�����~ҿi��t�5�P�����0�l`��>�o�ɶ�i���)<aS�{���Y� "��#����-���Mm���v�jv�1��w�ύ/��-����]�;H|�r$+D7��w���	S�eV���U������DQ�8���d��4�٘���]hbQQ�F��ej�^�X7��ɫ�M�m�W�L �雗�ͤ��a��rvOnj)��3w%m���ݽJs�Ĺq�y��Sh~�����|<�՞��h��d��:��M7!�Z`�-e����4j�,Jl�`�i�5fJ�v�Z�ZS$-�G6�ڠ[i�=�������muh�0f���`��	st�!E�g�&,��vlԖԙ�� 
��驦+���mځ)�\@�T´�]�3,+c
��.������,sԣ��le��u���K�ާx�ӠŲ�޲�4�˜3hjڈ[k�7e�6*--чM�>��o2�{��? VQ�Y*o����'Y�IXS>~����9���{��w �0�͌Y]tAf�@D ����S|�@�HS|7�#L�)�
��X.��a`�f��Mm"�����V���~$+R�R��~p�S�+��rם�����Ǧ�h����_}��� �۱�ȰUU��]��* ���'�*g}�u�S�a�c%B����j,�@�@dB!��@�����6�wu"x0�`�!m7|��8�/|��0߿w�	S�%K�</���1��L"��u�S��{͝=�z$�Q�FJ�����'Y��+
��~�+�
����2���u��s7�<Q��������YY3���$:SQz}���ʫ���<H|�=���I([!m ����1���k�_�x� VAO�w��!�Agc�3�y���q��LCJ�D���	!�a�ӷ>�4{�����,JY�v���k&�m�p�l�2�1*`�=n���x����&�V~��~}"Q�mf�'��������Y|���W2������2(��R�����AH_�7�����J�|-<����ZN�C|���%N�
�=���.��xC�� ^y�u;�c*Ct��/������_��({��B��U�.�Q����#s2c|NFVN��-�\<
����s�±4��j/G�U^��~�)'"&ۛ̚�?�&&|����d�d�,IXS?}��¦FLa�� ������ �Ȱ�^��#�j}�#jj 'R~���5L�w;�������z8�R�JZA����ąh$+ �����d])�����COw@aŘbs=����ǿ����c��Zs߿۬8	+{�\��.�='�<C�t0z��S���:�	!9p��� �z�a�w�N�)�<Bh%dajr�aE�� �)޸2�w��*}�Ci9�8`� ]\�DQT�':x_��a��so��/Ͼ��E�����gFN����v2��w��;�%�0�A��q��T�I���B��J
c��
\/׽���>�����~�_"F�N��[}�]7ER5X�]66-lh��
kF�,X\�翟p�ZIx�9��Ϸ�uN�Hgf-3^�c$�)ުT��9^YS=\a���ˏS��umm	,�y�nE�-`��׀$�O�)�A%@���*=AC[7���Q&�K��e[:&w�Xzi��:њB�K��<WJĸ@��
P�@�uB��s�J%%�4	%M��{�'���.�n_�Y��uxz��b���ч���1�k^+�^�q�x�_#��/ۋs�Gryݾ2be��K�gw|���1�l���y,�ğ;�>r��$��Ǒ(J
;����(�	�C�9��������M��pbI���o��
Hy��%1�B�$�|~��Ɨk�S1�J]�I�k�';^D��pD�pB� ��vu�y����BP�v�8�t������
Y��
}�B��$�ouE �J�:o�\.\$
�l��f�3CY�f�t����Y�큲�]�6,m#��0-�w
&�d���y��$�۲X�$�I�{z��mU��'$Z���r9�52+z�D��$o��
F�^����
s5�f��R	w�{���x5�/BRI ���Ъd���>�z<�(�g���룑�U���~�V4�
)é^H}�R���d�JI ��'F����g�s�As;����
�PI3���ɩk+8���!B�c��_:���˚���K36h�I2H?>� ��H��>���Օ��sرV9h1��=SwD7�����H=�O_9~ss>����AN`V�%MV��1*�bʪ�O'V�^�؅�N�B��Q	���&LY�"�oH���$�k��Px%�|l�Q��̒s ����$.�<�~k���I�u]
���D-�zH�ȭ�y��{��}�pMQ�mT<&�%�m�v�h����E��%e���D����5E�V}�����
 ���=gM i2I'ջ4#��Z�=�B^��7eb�k�wB�k:t����G�&rExpǨNL</k�� $��������>���2lI&I����I0I%���,����A����d�T���
��%����YuB���es��A ��{-�V��9������S�S;�Oo<�\�0��P ANx�%WS%�t�OQl��m�$�
y]M�Ky�e"N�t�\��ٻ�V���<�����"�H)@/ �ϒ�D�s��5ъ�0>ye�P��h���>�94I��יD������w�VX��l?e�Vn�/��~��@�9��>�v��X�oR
a`.&��׫>����s~��p���~x�Bϔa��X�WeX�2���;�^����~]�	��b`�(�����-�6�XEŗcZ݂]����J94�#�8�v��U�(�ґ�:���[)������ke&���kl��\�z��i�� ��a�F2�*�fj�hM��D�BgM�Q�ێ c-�%�t��藿ØyB��-��l--�F0c	�6b�7Z��2��6c1��LJc��#�����^xx��U]ck����intm�f�m��ev4�<�]��#2Fp��@.��BҝV�Ѐ%���%�t�P�	v��'���k4���{ٚ�	$�{�	���?�H-��v;�M �ʽ�>��k5W)�s�e��P��C%��"�"�>�"�J�u5�{	Mx���a�I'��r�E zs$M$�&���F;�yS��.�_�y�ä���D��{�U%"�
�rIx�9���M|���yg�=��1��t$�Fv^D�I&�͡TA$�w�#f����J1��I.�x ���#���d��恤�I��M	V��{�y�6�(�ϞeV��V�
�ŉA$v�E �X]�~���%$W9�s%F!ܼL:V�[KqLٮH����j:3VS�;,2���g���`�b�pJ}�RIzs���%:���q��y�ƶk&b�9L��ΑB�#͵��Y(D1wFC݅fꄤ	��ߗ2q?t��5�y&���$�L[e:�6�;����75��{�#Լ2��X�Z}����{}��gF������) Y�;�;�s#�<�������@k;��(QL��']�U���KΣU�X7����IDNg�)k�O}��3����	9�٩I$�Vv�Ou��s8$�@&]=�(Rv�w.w�b��-��t���$��?�5'������d�f�$�A ��ೕJ�j($�I2^�q�xi~�{��ʨZ�N�Ow��MH����I* AN}�2��ʹ^	$�g<4�>Q�(��f�Id�Тi$��*	&�[��s���=J��l5�13!���<L+����c����
V��[+���,{sfw��w�A<A8u����������⭚P�'�������P#�Xi'2zF�"J�Χ&�L��\�%����b���\bqW�Uжk�WM�i$	y�GF���HT��B3L�!�G�n�K=�bXI��1Pa��0�<.ڡ	*g֌�=0��d�l�J`��ӡ����sv�=B��yYr��2�1�D�r�W����Hy)��&��j3�{^�g�����;9r��"@��L�7��g�]t$�Ht>�=�Iv��)M{�����>��z헾ӱ��)�������.h$� �יI����s#�mt,�fy���l��mǼ��Y*�#r��RC£A-�y��w&{v|i�'z�����dg�n^�I������#]������:B�p����dq{��,.Os��ᯎ��4�R�acjl���30+Wl�t�ɭn���`������mU�q;�v/eT"RG/� 2H%�"h$�k}�I^=��5�v����I$��w�R���t �
'��	{��I ��3��?t[c4�qS��@$���f�ݒA�y��
E �׉��A�Gl��L��]A%�:�L+�G���H%��%L��K��{B���U1�$�ٯ�)4wl
��Fxx�;����]{ǳ�����7��u��wt�{dI$��'&�s��:�uH��ߺA����㯄"ޙ�+�]=��n��.��% �.{�o��t�������٥-���?�g���dɓ �d������ʾ�A��R�% ^��c;ǻ��3�H�3�5+�#�W�g)��RH*���(�Q�t(R$�e�Ow��L����Qh_S���^11�U��+�B�ntv��1T2�;Ks�Y�k�ü9���FX�{�
AxZy+�y��%�4i$J���9�9"rs��{����)&H�fȦ�����;������ڹ֔M��c�uA��M�>6S�I)��@4�Q�QA$��� ]��j��f�>4�W)Ca�P�8u#��$��4�	d+��M	$������[��,7���$��]Ц�RK����%�V&�qt��wN�.�6Q�s�+������̭$�zrD��C����x��Iv��K��[5I2~�B���J�D'ta��X���I�${q����8��N�x�gc:Cj��CS;�ȭʌ��A�.gw]�%8�p��B��1���zE)&HSEQ���PVm��9�f������(�=�BZO�՞�=���rI��w�:b�pJp轊�ۭi��bOY�A��'n���õ���ۋv_Iv1+�`�>rK7u�k�ϊ�m�=|ym��o�$��t�{e�����ݬ�n�
Z7s�u[ޘ�zק��M�]:%�ٯ�Ph{=�M�{���z{wW.=���y"�q?�����o��;��p�r�gQ�%=Ms�˚��c��C���J֏�a����%0!8X�+���9n��5(U�=˃�^�{�[��pg�#��j���ȧ�_f������}l\��o��3��=�' @��Ս����?�G�g|g��-x ��l<���\I�o�W����V�M-A�ۏ���M��:�ƇSd�$ݳT�@TK����\��A^�����gz`\�Dѫ�w�$�����Xz9��.�*�YK&�L�c��3��ܟsxO��w�t�n��3�>�y����~�+'zш����1D<�/M��/�����������'�>�k6B^��n�@���ױ��g���т_A�<;�~o_~Î�^�h��_a��6��}:�O0~n[���MSm�Q�B|���D�����.t�yb�z�:��?&bQܠX���pq�:���|77����'r�I�L���ǳ��7�{��H�n���.. ,~����qc�`����W�y�@8�H��	Ⅼ��nnT</Ŭs"��� ln��/u�����.�å3�b��6�we�����&(?	ǕT��"<�>ZP��a�����$��JIK�"�@����~F]/�,�R�"݉�����[�h�V1j]-X����B�Q@�?D��^cD!��~���Ω7�h���d��׬! ���#hW�+6�te��#Z���e�Z[m31�ٳ���v}��o�u�]u�Ӯ��oooo��|���X��h�:�QB�1b���5�.$�5̢���X�/-�z�6Vۜ�Z�>�O����]q�]u�]}:�:뮽�g�=�s�斥�([�S/r�E)J��e��[B���S�TS*s
�"��ơ�UYm��mw%qiNZ(���EkUJ�X�8�U��Z5{fe��a�XDI�Ũ)Ʊ�q�ض�l� $�
W̴9׿8�-��⒣m��l��mV(,X���(q�u�"pKERm�d��2ڈ�rʭJ���jh����3r�i=lUdf���ڤU�1��cV9h�(��

A30.U�5Qb9j�(�Z�U�Ԩ��hQU�(n�AQ��Y0H���19w Uq��"�沢#.Xf�*��X��d����+"��+e`��m֘��cTV4jEDSS���&%I����pϏ������͞&C,��8[�t��U��壮�"]�S�iUX-4)dq�XM�6��0�s���5H�I���ҩeq,D�q��2�9қv �F���F��X���)̴��]6D�gYf*�]]k�`���]G�v�#1E��mv��JY��I�p.���T%f�Κюtz9�m���K{j�skb�����i�8���`��Dd�F�]	���La�,fj�Énr�f��Ōz2��3K#tkf&���mVW��ڃc�0�+#�M),M,�݂Xf�i���R��F�r�挨��%Xն��s��l�4��@+�E�&�%��1m�R[+q�Q�iz��EIDe���J�1�C���۬tf�K�������2Ԫf�����rY{VLU���7�6�0��e�ܲY�r5�i���`꼌i�����A�mRT��h5�  ��B��Z6�R���I��"!fc��Tvژqfu6�A�mJ��]Q��hή��4m#��!�����my7&�X����0�CS��B��VZ.�;GfT�,u�i�T���Rƻ��hM�v"�u�D���	��kT�6i�%�q4��.AbVj�\���\�BL���a0F�ܷY�W������0��:Y��.�R�C���%�c)�	K��!)����M-X�@�]����lŅ�-
-Մܮ��B����,V�Z6ᎎ�tZb���mk2]a	���,*���C����E�V��"c\m���VR5�D�i5���]�6Z2ZGr۳�`�1�MÀ����aFYeE�ijJ�e �Ŗ���3�%�h���{A��v�q�)���m� .��e֔�IF.F��[�QV������)��r�Õ
f5�B���0b-+�Z�lf���k)l3���(�\�\�f\��+�U`����OG�k�zy��wr�8k��x���#?O� 2dɅzN�?|>���V6�ͣWQ�fժmP��5��)���1�Е���̰�].�t���QEc]Bn�A�%s�e�.8��4��[���&��i�&���u�H����e���Yt�ԃ��m��ɺ��fҌ5Z�qm��k�?J�#�F`���R��+,�1k�����0KU],�9�1�V��������:�y��P+6vn�J��6��H1�(�k[H�6���iZ��=�����P�??O]�$��%�/�N�I$w��@I{��5]m��l���M%y/���T��*����]�yN@/ڶ7�x���ǈ�h�MM�T�&If�m*	!��J�yRA-��1qu3���_�ERA�|��' �2.�.�{�@��H�c�槖J��wŽa���֎ ���e**gwIws��Sj�A���;Ѥ��s*'���8q�:m$�\��K�"�)u�̭gp�C9����Dn��PI
틤M\�:Pa�˼�*6�gY�� 93��M�^ίs���#qH�g%W�H�i+�y����
7���9MV{��>u��/{oA.�2��D'�n҃q�,���6^�ț3Leql� ̅4r￧���*����u�l�U ��H�s�59.��(�"a8��.���5���$�LU޼ʘ����D�1��O]�&T��}�I��U�7b��חoS������qv�Xx˿;��?�c_���w�w�oW}G^������faH�����.�/	�Ǐ��?=���ߟ��6��-}�M$�Q��	<���^92�2����Ug�[����؏�,@i�)[�y�I%�ǚcI$���3���H���^Z@E0I �{(P��A ���Kz�
�S��R�o�Y��.:��b}-��`k$�	�y��p�d�ɜ�c%l��z�rʞ}Z�}X�x�>�<��O(B��Jp�F��UȒ~�|��	�uY^F�5���ē���I�	�ۦ
Q��Ut��=X�C��Ot=��w��a��b�&�p� �2J{X�R��֦y����h����Ϻ�Q�3���le��3�:IE��H$�I[=QL���N��>f�iD�̢�I������=�H-�I"4!��OB~3��v�_��i��4釃��Lv\��I$�WOT���1Ɲv=�_��Ҕ4���9E����'�٣K�����H	Xw��1��fV�����߉��Ws��^\��j҄��?�䁫�*뽪`�뻋h�.���e�N�G�vu���/�g;��߿��J���yJ��Ǌ��ώ�y��	;�H�N�˫�k�#C�N����1����7j��V�pgwK&�hA$^Y=QL�d���@��>�N{���I��2���|s\�$�UQ񫩶��$7�!gP����K�y�K$���@�H���TS$J�w�sԩ����w}Gۢ>��~��gl�&M�������M�Q�ۛ���#v4J�Y?=�~��;6�I9���i����BRH�%��2�VF[n���Ca=��H�E�'j)+Y���;�O�y)�zj�A"�4gNv	��m��΃I�A.;=1I �f����M%/^�F^���*;�$�'��J 'wH�Hz �У�`�eΏo<�HgrsKX���	���� ^�$�?u94�$��᥊P�5�J<�LAvdb�g�E����{Y�Iv�Tմ���K#^d�H6�3��P���c:]?��"��'�ë�	�)[��,�+Z`�(`<��)�U�Fz������n�o�3���w���\C���L��!x��Ķ�ry���9���Ͽ�6��7�by��:�K�bE����D�I�2h��簦a��-�Z��U��R��	{���J�)NN�=�� Z�l�Kŧ�[Y�L��t ����TзM2ָؕʚ�j��S	<Ef%��0�A�嚲�$�&	 sq�	H$�'�ن2H�ox���l��˧$�K7��l��GxxO8w�-�W��h';�����Jٞ�Eτ$�+�ܦP	$}�%2��.��^"z��N\Խ�I��Mg;��x,��,�I=��1��H��WOY{W^���̗��(,|�2���IGuP�I�<$�1:tLB�
!wRȬ~�~��	0������A(ٹj�xgE�z��u�4�e��y�.�	Hh>�B:�$�AEݲG��ڕ%��;���4!��}|��TN��O4�r�e�@'��ԉ)�n�ޗ�HH�@�ٛ/���ɯI�ʾ�X۾�tG�v�Kض�y�k�KOӌ�sN9��U}v>��$�MƛS��7�w%cݎ�CQ��8�ĆA��������&��! dɓE�`BE� ����]3q��؆m�飙Vű�6W]����۬��!\
�5����¸�e���%]E�`m&�LiH�B�Բܲ7Z��@���"�yv�Wf6m������ۦ�魛�d
e1J�6���SX��1����l"Wf�YV��7(ݔ���[P�6XF�M]m6�!eu�6���Յr�&��M��,���'�I慆Ь�:�f� ��^c�s��a
�`��I��'߃9���.9�_.b�A"c�f��H�����RVK��\A��g-`~�-(��>�СI2� �ڏl$ü1��j˧6��;��h������P|��@?uЪI�t��󚾙{h8�q���w�A�*N��!��<�ލ��sF�E�W�hBA$�:��^S�4�r�t$_��U,d���:��NIjh�lW����BwE<�9�Y��g�9�u�ٕ��2H%캚4JIt>m=�I�ܒ�"s4�f�:uO�
Hz��xx�Q\�&!]��^��wt�\�T�T�{�����ō:I�~��^-�A$����M.~��B�d���I�Ӑ�wL��[�9��a(����&1�j�l`�R�2�֙md
;T[U������C�p{~'���I$��ݚ��Έ��rM2��c�y3�02:�}4j��8t���S�IM�*Ө ����'�bQ �>�B	�٤����r)dC�\��r+Z��՜�Z��7������I��B�=���޸�ok�z{7h�
z�t�Q͗~���y��eZ߀3577��2dɄ	 2fy��K�/���r��gj�I���)�PH�߳��2̘�
HUx,�0A�P �{�y���I,]�ZRH�
��iڋw��˽�'BI"�b;i�'�xI)�߽���1��M$�J�����}��gz���p1�pI%��C�K�D��q����T� �m�!��u�5�wXq$)��/l���M^�w0���,]�}� JI��4ꗺ�qճ�{���f�	=/T�$�$�b�e"��"����S���fS�E�1�0��Cv�0���4r��r�	M5.�R4u�c=�.�DFe�{��:(]��h�ۚ�gwI.[�D�H$��"i%���M�f�x|�zd�@$�r�"}>D���;������f���������j�Ss�	4��/��Ry�:d�d�=�H��x�|srE���l�{R�I�I�J�t8<&.!�l�빞�;;�J;vh�42hhI"�=�F)�k��>��L�j��M�FhzN��X1K���u-��޻�qn���P������fO���{w�N�yM�9>�� dɓ$���s��$@'��(��~�hU.o{��uA��^,��G�C��+���	Z�P�K��B�$���Q5��Q��\v�gn�H,|��B���x�D't�2]�ȚI�5�Q~�<��q\�	:��Je"R|�$�@$�J�Rv���a�#��Ǘ4TJ��1�k\f�V`]�JUZ��\/30 3\�`d�z��(wHC�S��\��D�q�4$����c�RE�ݿ]�z��v���k'����$}�(R]ttQ�P�9tLD�񈎉��K��W��UXbM�>H���vP�h������=DYш�淫�b����+Y���M��m�
.�MQ4����H$��͉&�$w����bg�L�����H$���'k�M�Rh$��Z�	�F)Pd�|�������CC&r�쫚%�,d���*$�Z��K��6�\@�b�̰�^T�z�SQALN�r ��%ե�v�ݾ�P�����C<�+�_,S���Ӕ�~����eqkT�v����_�/N�/"[ǏD+dfxd�����T(R�����]�1G�i�ϕA�ä9<��n'y>�x�l%�7�B���=J�I#�9KJz��:��;�'C%Z�È"� ��X�K��%`Ź�	k]\�f��h�K�ٝ�=�=���D't�I�wI�+�i2D�d�m#�2��QIU��A��7����+Y�3�uկ�T��7\a�!QO���z��Rq��K���fW�S�i�(qϲ��IϜ��������_v܉6)��
>e� b�F?R Rk;�(�5�A�@H��]���m�~�8��IE�u*I2D,�2��z�"��@)<9�k�u龗��X/�� ��M��M%�/�@:I �׾S!  �����c����q�ȝIʎ�3���#�x< �(F<�׬PI |��Wb]뢙��3��RMA�2I[���� �zx��v�C�'o�O��s�{���c�:y`��8B�����屓J��:w^���=0��U��bQ���ˡ�~��t����1��1�^V�b��h����os��̙o32�-~������$�ɓ& �g|{k�K�����ؐ��F��cLf�kإ�g���@���J,ɦ�٭��љ�sIjB�ԋb���q�!-.��z��#X9HM	M)��4�v��R2��f��i�YI�e�^�`D�,�A��	��2�i`�a�K�
�M+�p�+H�Miq�$KK�,j�0a�Ѵ�1t]��1�l찲��S�3_1GL�SmUrm�Z35.n]����,ѕ���_{����.� ��;��θ�#,���x�|���Il��EP���}�)k4]C�V��As�)��lFv�	�:��]�J�\=䞷iӴ��Q���^f���vH���SH���tq�JY"��p�J�_j������	��$�.�ݭ��m���D�te*%2\Ap��.ɟG�$�8���BD����&[�xM"!�@�*��?Vl�
>�ɊGJD��R59 ��=̼M��!�WGR�qo�;��X�;�)�<.�E���Ux%���TZX�J;_f�nF�Gp�噉(z�2A$E�jD��:�T����.+~�Z��~��<�.���T�P�M�Zf�h9D6`�<��j�&Vm����~��8���s+z�2�I,���H$�$ϝH�u�������,����J("�GE������N����7v��*��	"�'���Õ)7���-�ɨs���߆sy4/y�`{����7yQ-~�w���w�(z��z�BQ�I�S���+/AJ��T��%�����`����<[!x���+i����������9l���~�y��ak������ʒA%��ʫ��>��*4.�(%D't�M�]Mʤ�/|�4��|omk�q3T�u"���$�O�H��]b��0�!'�b픿yq��]��^�e-~�p�$�ȯ
g>	�7b�PIȥ�ܼ����d�^��@Q��<'Ȉxb1
�'�{��T��r�S*��%>�-��$����� �$��J�I$?r�*��oE���k�Fem�G���m�akպ�\[��]fi�A� �3C0��Z���`���(*I$}�٠��w���S!'��o���ܢ}u�cK;�D�� ��*T���𜢡�R��\�� Yh^�>��ק2���*�Ν���X�a�"�~�"S�p����ew-��aw2��'����>Zu��.� ����W.q�@%��L��L�3��Z�yD���IO�z�IHBxF5N����-y��B �݁��I���T�=���DMɀx��S��^V���r���\�'\�Go����k��kM��W��t�͋Ӱ��Պ����{I���O����X�o��C�н�|:ڦ��M緼�G�sޯ��߹��>��M[��⯌�W����>v��`���,{��r�纮w9���^n�FiPR�s�u�����"�=���e��,�ׅA��<
h9�c�ٻ�����/�4]�Ē���w��Ň�z���o����)��{y�s�}�����+1�tp���a���p�]9�c��_C���<�Ko-��.�79���ܶ]�}������	�,z/t�~ٚ��呲�T�o����<�������_��$��k�%h�AO�g�����{����[C�_��}�����DqND�����'�����H����Hb�/���������Π�(V'�樬g}�{|��b�_�͝�b���;wpgk}raUU5���w�ˊ?2�nL��h�O�{ǌf]��Gof�\�\��v�����]���;ѳu矼�����.�n�9{]=�)JaJ퓘�X��\�U��[ßʿ{[���@��,���y�a��Y���݆�6h ���<��3Kѩm� ���_#���v<���'_7�����+��0��=��>ɳ��8�(|}ek�w��{��8�=���(q��
��wo;�s���W$n����Q�^��̑��7�H!gw�򘆉D*Q�Qk@^����C+T�*,��h�iӀf(���R*Z�"e+���9^=��N���u�]u�]u��뮺�{j��z��ˍ�m�[9��QPX�*�(����l��B�4b2ҥ�UTB#>Z�rq��{}=���u�]u�뮸뮾'�ΦrܵAEX�(���1*J�+E��ܣ��i�Q��KQ�F��DA�J!�r����(�bPĪ�-�b��R�m��J�X�DR&�8�,-�X6���[��m�핁���EE*J���QfZ"�EQ���ʊ�*��PE�
(�����+G�Q�֕F[51�6�ı��X���t�SS0*�Zc�Xj��D0��Ĳ)��UfZ�"��"!�0�R�����V��A*TE�EE���Y���EKm�eF
+��+7.,�T�Xq��Qkg7�ūL��ͬ�m���Z*�PX��Mpx�A�U*TE\�Tm-UKj*�0UEQA-�-|)�h�QQ`���Er�2����%>�A�T|J��֫��[ssnm�ʪ�����KǏ*��KiDڒ��}|��9�ǎ�>?�NM$����3������wN�Kx�ʋ穥��8�=����I�T��,Ȅ�Z��e�D�������|'��Τ�cש���A`��9E<
��ԉH$����U�G�#Y;���1����I���PL��7OL�������^�Ѓoۍ�䵘.q�(�f�u(m���V��5\��R٣�j~����H� �D�h�SJ��BK�ʷ�S) )�:x��w��׌���w�^|{�zI;;���(2L���N� �F"�^%s�T�ȧ.��Y��\��P�Ml����i���d��t��i�	V�{�>���q�B�ntD'(�s��=r�E��'�#<ʐ@$����y��S��䓁s���RK��=\|ԀBv�:І�c�=�o��.���v���O�1L��Y�KC����T	$������^3��=��H/�=���m����`x�W҅Q���H��>�ï�������`���9.�!)Di����`�G��K���
^<x�ֆҍ�!a 綽��xr��y�Ը4�?xy<`�x.�֝	e�]*A"���:hB�b'^)�s�(�RITzx�-d�w����{����b0q��l-Ա�!0˂\9�х�]�eݗG6���S.���h%�`I-��r�B&�����*Y�&I%qѴ�/3�u�q=�wjw���W����k�)("��\�Rޣ�|H��@�"��w��U	 �z�c��|��Z�`���K������Ke��$����F�{z�!���D(DB��K�qԩ2I(n��M@x$�A.�����jiG,��Gё�I���OH���-sb!9EC��<�U=	Y�=ȍ-0�(g�����PIC�ӒL2j�g�[E�&ź/��(�3��8i����S���av,��I$�.� d�v��z�=�������$�v��A$��T4�d�
�у�J�k�8۫�����v�V{��4�<����yni{���ٍo�#v{�>������g���w6��������wv`��������|q�1�s��+j)ky�s�9~D�^���O<yT6R��'�����)r1�iFTV� �ĭ�f��]B������P���0i+����a��nZ�v�QU�4���bn�,e�� ��dFP�`m�t��*�1��,. `ʰJ[���ZiD�V7`����]�Ql����Yg�vW��l"����.Rۡ]4ЖK dЖP4����Z!��v�ܹ9"m�����i�mZ�R�*��S`v+�۬����n�a�Bt>ρ�9��1!ӯ��K��� �������@$�?j�K/��FGn�S�M$�$vl� ��;�+� �gm=	�V��q�Zw��O���$��_K�I$ \��CJ)'����T�/�m��Q�L�pbR�]�P� ��Ϝ����n����G��=�h����H$�C���JB\�*e 5����Bn�-`��ƈ�����x�n�)'�Χ4�w�sd$�s;��t��ך����-$�׷;����k������R�	es̤I?de2�aP�u�D��R]�R��	$�q�Q$��i�K�ϲn%�b�]���B��}6�	�m.2�/f�ЛqpX\�%r�vh���O�؝`r
t��4Y�qTAy���yiI$��:j��=W$p.|�����'*�$�$�H��t�/�X<`��Ԋ^��NPT�NeY�V�O�=��`�L�y�X�I{� �;ϟw�5�/��g�{�z�����a{�A/-郇b�~��76{y
�s���y"A���6sp1D�$�>V��v�y�e��}4��D؆A慛S��:Z_l��wwO����ǏB�&Е�@�K3ʚ^���I$H�kąl���O}>2M��|�����3�~�r�B&�����7���h�H�_�.�Qd�w�=���Rhr.���S�RW��(��O�:hR�/�AB�e��^���6����$$�3��
 �/\�%&lֈ���H�I��[�T�z&$����$M��	SO^���x�vJ����+gvu;Is�UǼ�>�x��A$��l�+d�Σ{�M�ivb*�Qg��˵Jt��($�fڬm����J���%Ml�ldVfRWL6��~��O��	�*j�m�JI$|��
�H%L�GoW�%�jvѻxO���ucȔPH��l�R��.�9%;�3��o[�M�PI��Y���S�{��a$H�5Acw��;��RR�y�]Ow<��Q!:�O�c�K8wIE�D�	���z��R�)�{��=B���/v��xq4<vw�����^�Ȏ�T**��_"-6X�YX=����>�{�Ͼ�������r�7�������KǏT[![[�_��>+�緞x���t�"�H��Mh���.P��(�º֕E��-ޒ��>�s��$�x��*�@'%s�4i$��î�s��׭K, :K7'�
K(�x� ����#nf�$�	�x1�3�9^�N<ǈ��p���o�4i"Ȥ�ws��^ty��t��Jw(�aB��C�{��lh�����.V������+��l�j����;��Y�?o�'�GR��;��4As;�K��<�!-�y]HH����ዚ�4I5�94i$ݠ�Qc�ֈ�%b�>�=�)$Z�T�١��Z�'�њR
��:[�F�%;}�z�l���]=�5��mI�A��Z���3�� ���:A$��Ǒ(���l�oX�?Z랃�I!잚4�D����R���U���C��ߦ.=��{+t�z��vw�gD�H$����e�$�Ә� ���N{i��H�w�%��nk.��皔������BA;�Ѩ?����/.�i���X�>%Ú[�B��R��ξ���?��6vL�
ɓ& �`  �`G�ﾉ$П�-���s�"�&z����O�GR���rN��?{�J�.$�I���!>��^g�I��f��|��N	r�!(��XͲ�e\�p����M�Թ�q�隴Ξ���$!I.B�Y3�V�wIy����̤�Oݰ$w���x}˜����$
�t���;��Y�<�z"Z�/=��z��kkf�e��$���{dH$�EO��ݾ �%�y�h�A�P�(,��6ŕ2ӑ@�I�}�@�V���ډ�B�g:�%{�D� �$��u��A҆x0�k��[Ư�_�G���o%{�l�{܁$wP�j�iUw�KsEX+�O!�{���ĒH+��h���U�@!���O���Eܴ�!wwUc�߸�8�}��Շo`�no��T9!�Pm��\��?p�>�v/y�s��ɛ���g���e�@��w��wn�g��\����)���H[�j�a��z��~a���O"��ǐ���6����Zҗ�������^.��i՚�B��fhFEi+�0:gZʚd3���)l�1lՎ�ʍlI� �v]�(�3t5�;���ԕ�`@y-�gc&K0�q�z�&��s\웄#�:��]�+\P��,e�-���H�U`8x�c�ƙ&%z����
�]�7@��]���k1Mp�Y���!�4Ա"m���vc���̭��ƁX��n�[.I��f����W~���%�P�!<GP"�� | �Ή$�&E󺪍gG���^ݲ��dK+�j�@�K�4�T(��̥�m'��_�D�@$wGuL]�TM�8.��_O�LX�wwG`�iړ�tI �k.�ٟ&(ڛ�}y:q�����"��Ike��3D�n��*�;�%c�����yt��	>���X�WGoU%{���?g�6��Z��,$�Vu�Z�$(g�^a�~ʠA+;!�+�m�ȼO�(WG�H,1�l�d��ouJ��F���h��)	$���@���J�4)*�麬*����,2˪F���J��ٝ�I[qNS�xw\3#�8m�h	���a��z�~��d��]�4	~�"�M2�OspY��c����w���~^z��� �)A��\�fV84|�?k�z���C%�s����%z����Q�:��c<��������J�-��x�<y-h� *��$�y��O�e�����z���	�}��Gq�a�d��(@�L^�u@S$WgD�$f`�j>�lW/h�1���n�A �̆�2�J�K�
dR&�����ޚ��0x�U\�pL�LP-;�֡M��GL�=�K�b}�)�L�π'�769ߜ� �(sl_��$�
�Ȑv��'�{q�`��۠R�:�u�oH�Vr4�1᥸Z�eq�߷�4H\��E���V��r���b��4�nw �T	�٠��r���{���T��d�'�)��p�c��Z��Y߄�^�x��I{�D����8�S����>��>�k=�D�%ߺ@�Iw�K	OV�\N�u��i�I���:w9�~�p`w��/N����`�O�����Շ����e�O��x���A�����7�u�;���o��%򁻕�p�4�N�|&͞>�<�<�Օ�ʫ2 ��������>�����������$-�9V!0Ǽ����i�(�R	c$	W�I ������&q�H�ڙ.��+\�\�Px�}�^��I0ő~��Udi���瀅6Y9YsLh�^@�X���:�z�����,UP�.4��hi�j���2ґe�AX9�Ùp;�5�Ɗ7��S]X۠�?>ϛ{�&��dp�3���nĒ	��w���Mf�u"��ƻ|� L�
 �t��Y4�p/n�"�C<d���^� H�G/���᮷��	;���H�2%�!Xd��5�(��<#'�*�NٱW�$@&��Ҝ��H-�d@��H$��MA'���˙�]H��$�_7�h���9�˒�s �x�g�wWy�y�٪G�3o�l܉c�ى`@'̑��eD���G�@���_|^����0z�Ϣ�}7=����-�/n�=��ǧ:��ˀV5�k������x=���)w����;�xwιpG�	?�2d�ɐ�L�0��
��Z��,���םߤH&�]`�c<x��g ��ΐ&w:F;���w�H���I]�_w��~~{��i��z��ޑ����i�Q�\<e���4B�bS4L!4�u`��g����K4A�U�H �_�6|������>�����͌�k��H C編P�����IC����%�/fU��D�S���CY!����2dX��CIq3��=R�e���j���� �C<�꾪Y"X�vL�K�ɬ���[��c@�Lu�MI+{�^m%��9O��U }�Q�DN��΢Đf�i�$���B���k�^Oru-)�Ų]��NŞpM�wF�N�M��E�
��U��W�5�����X�Vv;CIw�Kb*�{.q�~'i�r���ӯ.ͭzyOh���5��읝�b�F�?^�Y�YV6a�w�f��~����2d�=����7�>K4x�(��<���
�n�3x����t�=h�c��q۩m�k�G��<B�H�x���[˗���=��������}����{��L@������|�:��f]��w]��=����{#�-ǯ���f��.�k���w�ys���:D��y௕�W����9���t���Gy�͸<7y���_�ڕ!ݐv�Ob@��墔���49yѧW�����P�����&��ĉ�q�O�.w[��ޝ����jb�!u��];:�<��� Y�:ހo���G��y����Ǯ�oB�G�����S�1�B:9�[���X���q���$(ŕӓ��q��!��
緍ݸ�k���W��ن����^�w֨�f�4_stw�=h��_�!�������Ih��&O+�Q����������ر ��z.�߽�zy��$3~�d����y�=p]�iE�z�{/#��&o�2p�D���/g���ˢo@��_yo/
�2��W�k)�B˓��q#�nK���bi���B�1���١>Ǟ�{ۍ�lǷ���c��qk����,�x:;5��ɾ��������,�X.%��/��d�< )��6g:q
zԏz������4ȼP��s2���d�MF�tgo{k��,�����i��i��gT8���L�4�ζޏ��hԃ�%C�}��	]�ݛ���*v�zhdY m��pU��F�	ژ"b$%�F4},p�h��.o�7��9�1ٹ��0�G�9%�<k5-���M��ʇ
Zo�x,Y�����Mu�]M4L#EU��n�]��|�9�/j*�UVE��Rv�e��(�����!�����m��UQUF[b��z��[m�x���|���{{{{x뮺믗]u�]u����o5Ŷ�8�'-TJ�
��F�ETQPrʤ�T�QeJ� �����[�嬼�ּ�+�Oo������������]u�î�㮺��U���IDQ�V
�cm�������Q�S"塍U������ˉ��E)h�k,Db�nҬVڛiQLR�5�bQ��̶(V���和Q��)[Q6��Z1����TiKj���0����[a�c�ՋUm�kUE-�m�im����Z�Z+�11,DQAq,q����X`�*1͡QM�&Lۀ�TAM��i^A.Z�YTX��E���D6�Db&%E��
�E*���m��mQq�ʙ���4�jQ�Y�X����b#�e����Ѯ6�A���Qb��EUݰ�\���U-���b%�ES31�Tc_��*����h�8�v�"��������E�b�F��/��xmar�.�#�kmX�6s٥�دl�΁̹ԫJ�G94uI���Υ�ZO�ض+t��0�u��!K����#� b�����r�҈L�:b�����!�
�#N�n�J���LkD��T�95�-n�e4��n�,�fW���x����")�Lm�v����M�� ��Чk �.3��,�����+�\[�«�-���֔3G!`]h�T�唵�c!sr5Y�-u��s�fvԢg*�l��`�r�v@�3�aYs�D�����f\�,��`�E�**k3�9 L7n�5J�V[H�K�S7Fat-b�1�aj얙����&��eh�Ż��e�V�6�Mur��v�6a**��tvWG%�P�B:�K�D ]��4��+K\���4qmH4��t���Ҫ��������h;��F$�[Vjf��)�r�i��qݢ�k]�m��,]4�$���n�ԡk.�&���X�i�g�u�����e�ƶŶ�0��"(�R55f��u�,�F��R�ѕ�*�32��c����L������l�ڒ�D�r�38�є&�\CXHu�ք!l��䁵��L�&@.��[�!-%�&�0�np\��9F[�,j8V��i���G�����F��a��[<�T���B^�h�ieƚYhCݫ
kj��Fr:�aJ[��%4��-J��i���5�Q���GK��LP��B�c0iu;U��,a�����-�o��)����8���i��F��b<�s��d"�0M;҇389� �cve��.��tY���*\���n�-s.�R�-�8ֲ�(Zi��GC-�B�U���f�N�92�cJ����6�.5*,����x�<�s�jk
���ݙ�M�*4�]���ːBXU_<�$���U�B�nW*��%pnks�ܷ�r�a�x�Ox���V	 �%ӗ�:e�v�0ڌ�m�R6V.�-�bj�˹4af̤��)
��Z������c�T��c�da��̦:�f0	VS�a��[x�5�X�֑$05�JK�;+L��3kj��u�xm&sD���:�MV����&彥e��Evu�m����l[1nM�u�T���[ ж1^�f�l6�VԎ�ʔ��U�#	JGuiYCg[��h��6��hŵH̺[��э&L�?��������x�&@	'Y>�T�
���cJf�4V�.>�ˎ�s�U@�{�-��U�~wB
}�*��&X�/N��>;ٿvMR@�H{͙`A`�zD��e{�r;�'����y�A��(F*�~��!vdI �x]S��yc��oIߺK�A��[���'��'(�8��߶/+�f��p/�D���b9{b��Y��h'��ɩR��9tr��n׺9����9O��V}7I �o׳LH���|�LyZ�]2)&%ߺD�d�9�4���������';L�4G�;��6������]5;Bk�A��{ k���d1�)�X�!����}n��x�c�9s$&H}��'�����N�gӏ�&s�@�@%�^Hi��ᕠ0��I;q+?�p{���܏���AUذ�4��>�t��U�7�ZנyޫP��D5�.Ǜ��jOd�N+�q�y~纯�-���͹�H�=�Tvv��.C�=]����^ޞ<U�Ǐ	�d�@Y"D�"
�9���y���ٓ��T�W�{ĝ]~#�.�͙�9������(<A�+�� �|�bu�������dj|�~�A ���	%��z��'h��/�D ��1"�������ε
H�Vlx+�� i���(�d�{��;������d��l���L�4>�wt�(g��V]P$_;`�2��em��������P�nmW$���`�}��������G�k].&���+�1f&�!WGG`����{iB�]K��C	���O��\���@���D���"�%��i��TO�p��TLY�@$��ʠxd���;ķ��m$�{v�ϯ���"	  /3����F�KK�v2���,���LM"�SbJ�;��O��@�@"�:fX�v�4��(��.VqH�	���d�}|��ljV��D�s��~>�Nm��?�g��	E��vY���9��}��́�ɓ X(̙2b�Hȁ|���Q��������v4�'�m�}rj�]罼ܛ�F�����IW���$�H�Ι�e�+�_�6�Sq�Y2�=Tpz���!��$
�1��$K,���p���ܮ��W���cofAbB�2|����p����PZ|�Zif1��ݗ=f�5��b��1��\�4ܾ�>����Z=��l��RjE�&3vD��H[(�~4���hU��.�t��@P%�1�gP�4g�V�S��^�x�Kܯ2^jm���8���Z����� H����A6��� )�[�]qOz.ޯ3̐�%��N�L�}bI�I�S!�S91/5���Ϸ���	3���J�}2ĳй�^�q	�U;�utd]D�z��lD�z�@����IbZ�!oTa���r��٫�{3B?�hߞ�G�����˜���i�ݩ ��vl���V�J3�^f�5��Oߤ�dU뿴��V��>�o3��;;;8g#21E�A��X���9�L�'�+��� ��G����$����4kǕ�cL�;2	'�㌂H7�����ʝ�`qAa��ҥ�k-4^#r8y�1w0m����m��)��7}����]fP.��Q��!���؉Du�hi]o��иK�9��L�!�dk���@�{4>��9IC8��מʡ,�1=�O��_��� � s�a�Je����@���φ�L���~C���T�^�Lr��Q!�=�m�l	��r�n�A����O>oM	d���Y~E���Rx��tg�	�����׻@H$S�mS	)�{w�/�������H�d�����3�N� S��Uٳ<�h�7�%�q�A,x��l˱�A]�"i���~Qs3�.��<N�TdTbY�z�^n2$w߹N�T������^���9���2�GM�"c��Jg���p�}��C�Kt���Ð�t&d/�o��0�:S���(�I��}�:n�&�
$I<��k���j�@��;�\��-͆!��^͗bl�e!���CM�]pl�� DV�:� 0��܅�B�B��e��P-i�x[�l,H�Ί�fܗVj��L�\�YSZ�YF�)6�lix�H��5c�+2)S+eR;1b^����6kA-4��E�i�ˢe�Mqn#���:�j�]h
y�0��ȍ�thb])6e�&�(bd�萱"�e��ͪ���?���c� ����4��d����D�%��E��}�+$9}�fO2�E�UZb�+P�����[�:t�Ƕ7+��,�cOy��wl0�]]���y��#��Γ���B �n�ܦ���"@ �L�O���Avi�s�̂A76SFPKJ��ú�0�{�|�����UOW
/1ޑC$\<�T�%wF�JK�l���(KN����������}72@%��>�{DɧC0��<O]窘����L�K�F�ˢ�%���<� �OBxH��u)�(��g-�Q��6��%�]��mZ���s8=q��u�<�$od���q4Ƙ���iְ����-+�g}K����)�1@���I`I��e��
<9�g�t"|�ro!�n�}s���WK2+��>���WO���=�\�zX��k����)���D9N���?v+���ջ���x�݄��]�Y���Z<U!��g�<��<���Z�i��{*�� �SL�d��,���O�LRO����@�A�\�Bx.�� �Wc�ң��ykfc���vKKJލ2	��r4AwN�3����W�he�z �%�OzX`N�~2Ao���A�+�|deG�I\t����<
��<�]C�x�{���}�"��^�����H%�tY I+w���_�կ����}~~�)���"8��#x^�2��f\�XE��k75�%퍝�]�}~O^���S�P<�\� ����	 ����z��W�h�\��P���8�5����xI<Ho]S��Iϼ��{� �d���̂H.��A�|�E�_2石���g!��1�z���$]��CKS'�� p�<y�G����+����[�Ӥ��3�]\S����Wl�5�w����w�k�xbK�-^W}������o�����F3�نH�fL��5lV�2���~>/�m��׽�=�?��6�ܛ�rxB0#��Yo��a�X7hv�J �W�v��wW^�����6� ���g<�ƶ�w.���{�[�E�/���6{�v:��&䖋��$���DI}��B����_�|ѽ�ڂ�1Җd�"4ueps5�m6nͱ����!ǽ��!�(����;�!2���D���5'�3��;�����g��2!gwP֋.����x��{�$Ǩ)yu�s����?R �3j�2F� ��T$Wf�n�Ϲx�7�r����p�C�MչQ�x�� �(�X��H5��#tp񦢳1�� �\��%�c��2F5zN��p�ϼWy�����_6|&�����(L�$dwL�A]����t��˂��J���uG��ux?En�����Б?ۯ�"�׊ث5��}�vۻ�۾z�~����n|��_������Ǖ�Զ�����[������~o�]��W�|K�B�&fqY�USϟd-����F�]W¯�z��m�c�2˹��ȯU����>Q���t�9%PvK�4�&����K���G�ژ-���iZ����PS�{$C��P�Gu�fU	6�3�d�d��D�M�y�����oFz�;$W���2�i�����Rw7�n-��B伅P������� ���H%oG&R-#^��{�]"xw��W��"f�S�%�(���z���p	X�+��@Z�q��;��x	/����"]�M�9Q^x�~��G�Hٹ��""磻�y�$�-���;�y��1&:�%�.N�xpaϼ
�>�%�>vȨ�Sb��fp=�E��Hw��&�h�OUP��IYʆ���}�Ng�����,/���M?�~���a圷���cF_����/�xw�� �o��<��o��}|z�����?��x�'$�@�l]f[��: w���ɓ`D$X�Ǻ�[��in�\l���bU�k f�z��.T��)��!�@�3��K�SR(�4�(��˙�o�&"lQt���]M�HF �P��)
�ż�X�If��ƺ��"�����Ͱftc������h���)fh�Ke�l��6��M5�g8l�)
���4��z�b��WKi�0̖mQk��ͺd���j��9���soW
,�E�1��-�i��b�@l6n����gt��"���]K{� �?oK�n:��_��[ �u&�$�h��L���r� �wr�����*�$+��v���o���L�,��I�)�ѳ�M�� Up�n�u����Lq �xƂ�BIѶ���.�*d���=QX���W����LK�̉$���@ǆK���C�wuގ��3A�L�A{ [$u�+��1��ݪb�"���ޮ�pӜ'��D�k���T@D(�Tcz�=]���ɗ��&�(�H%woP $�qi��Cwr/68m�I1(�<�	k�V�A����:���¡��� KZq����5,�������<�~����% ~�٠
d����M���{⧖d^��T�%�'��5��Ƃ!È Q~��&�Nx����gU����@��į ���L�8�xo���HO�t/:v�q�zs�69�J�p����	�����ק���Ǐ+�V͛-Y���� C��v��$�8��:ZAb�����������'t]C!^ʾ�`Đ)�|��$�Y=�ʿxTq�N�b<���f=݂J�A���BP�N���{��{�[DWL䑥�rH-�Smo<�$;'�\
z��~�=#|� �oٴ*�po�wQ��nz�IY�
e�~�44p�����E^{�@�B��i �H~��,|�x!��oU�#���u�R���ř�i5άN2��``c�6�&���R1�ɕ��|��q�a_��߯>��^g
 ݙ �%���Kq�s�6������!�:X��A���"�PL9�+�q$N���^��w������WoCI��2ǩj29We�EqK� ?�@|����H��D�P�Kux����䦻<qgyՁ�پ:��q`RU�zo�axaM�����'wg����O���QF�a��}��g�=j�7DX�!����$�ydta�㛰��A<�u&�^|������=A���dq�*�/�����I.��1���������L�����w'�o�Ґn��ޚ?v\�-+ǆ��G����z��	��;��΁�X3$��Mm���[pG�o&"+c�;�o�P���i�>GUOL;ni�����h�t.�ŷ�2�j������&JVuϸ�{��ys��M��T���MDk��&�� <w�{���O���Bzm�gi��o�k^Uh+Ż*��5�����ŏx�B����Ԫ�����}���g��ٯ_��i��{N�C��]ѓ|&����ˮ��k;�]�vn��`�<�>Y��n�xe�}�ug�o#=iȰL����Mr��E���#C��r�|����[O��ؾ�=����3���|2�~#zz�3��s��������8{��<9x�A�׸q����M�{�:ʸ�ө~�*��5��P=V����h�{���#�C,o���9͛.�Ж��7|}��X�NΎ)���.�CWZ��;����3p�񹦥�o���a��x�9�o�~�z�u��Z�����D���Q��}o!]s�]�r��]lW�F!��E&{�^�p��U�;�欽�-�}���R6�y��P"���u�����Tׇ,^���8�z����D��]�V�}������;��W�	�0瞑NNVk+ߠ�;6��6�UQ�p>�rX�X�.A	�wi���VU��)kJ��j���r�"���ő�g'gg����������]u�î�㮺��_��\�kEX��h*�ڊ�V�)X��������Z�s���z|=�^�������ޞ�u�_��u���j�ֳm�XV%e���*�F��i���[(1�mE�AT���r�PDE@UT���8��(���#�[Z��pjEUQ2�+!j1EdQ]b��DD��"�1*��(�b
����j�m%1�Qjc�b�/0�Q�kj1��EQUu�"��E(�6�DP��ʻlR�kZ(��������-����X���ۙ,E"�[m���8(�֪"��e�մ�)�X%kj�*�U�T+YQEX�ƣh�l�Xe�(�P��+U�����*%�v���:��G-%-U�Հ�+�J���Ŷ�
� ����5*��A����'��l�ɓ&`�	 ��0-7��?	}�����J��:М�����鸞�FV^�l�1W�@'�H/��������	w:���ߪ�K�\"��y��dKĂ�ݓ@-�:4@\��*�}2	 ���D�X����Fv�+0@��y���Q����q]�m�0�歖�Z.�2Xи��&��lT�	�3I��t����Y�\�è�N\M2@�nD�K���.\)|Ɉ�>��gl�bgA�3�ʈr� r�wL)�m)�?Dߧ{�=�%�9��z;�%�����Z��ͨ���̰a%��G�xNR�a̓]���;G3��d�Q��·��Z(��9��nK	�v7�����)kA��9���\6=�g#��4}��%�����	+{��<h ��5��Qy��'�x޿��Y����/Z��߬�t�[���V�7�u�m���)�����{���)o��=�L��%1��V9�~�9��j<����M��7C���o�	b��uADy�7�4��D�@=�T>�H�U'և�WN��.��y�h2��YI���6�
�q������u݌�փ�T+�7g5��~�w�sc�O��~|�$�@���$K�tH'�ɮ�b^c:D�a-����.�b�!��:���<<9���I9ј�w�f��`$�I�{���,H/��$��O#z��>�^��&7�y�@*(S�6	��"A �GN{��}\<H%\{s�b����}DXw��C�}�W{b�C*u�v*�/}�4Đcw&A,@�O��&�{��V�����h>I[A��9�zz4���$�^�𵌰	0��M,Q�Φ���!�DlD���<�OR�S0��W�wA��n������z�D�V���+��ؼt7��5D����aV.�V1T�G�ܟ�<A���>���0PҞ^�wל7���̟fL��1�
��w��n[��r��v���f[��ۇb��|/����/"\z��7Ui�ET\$E�L�� ٬0MH]ne��M�LI�R�a��s�Y�Yk�\�du�CED��R�Kr�Z�7E�I�(�7i�̮v��]q�kG�6fK��A�`��eW�;h�wc2��,΍&3
��i���%�Tw7�Vf�J&���Y�Zh���*��˶z�ؙQ�A[vq�eʺ)��6�������+l���pc�͛��i��n���C�t�O51~��1_��ı�ٗ�'tN�C��
>���@%2����(M�c;_2|$�Dn�����H.�Y�=U]��s4�Gs�j�1<8x��O\	u�I �L����|���O�;6�7�"A �ݲ$�a ��+%D9e
��ʏFPz��f���)�/����z���|��H�$���-�E�s�80怠
�lK ~͑�u�P���$_G�L��{"A$����'�3�r"�(�"J߯�xg��YM
htF&�;0�xt�����5l�Y��������W4�8� o1]W2HW��	$����R�����r�ٶ^��A$/lY�Cϱ�D"�xU�q���c��w�b�ω#Ę��{���=`�Ľ�gNY��sp�,d+U���9�y-*C��Tǯ��5UXm�Ԫp�$?�{2a�&K�@` ���?�$��C����fA �}j;v:z�_6jb'	�q!�R*����"	/z$X�5$���z��z�a����d	bIn�t�"Y�1R�<�Q��7=~���=S	���������I%�L��b^e�:�dw6d���s�����F_S���$�uӂ���Aj���a�+��O7������
��̛�硐�HM�yT	";�d��u�����g��O�����c����J/�����M1yF[����6ƺ(AWh�v3Y�jU����;WAŷ��y�� �ؐKc{�WFW	���z8� ]y,��=�����#@��X�,��J.|�q�62� E�l�&%�s0� J�=�y�1�Yɳ�֦�_�,�1%����fd ���HB�a���>1� ����^�mG�m����7s�9��Û�+�W���eOl�u�ˬ�H����X�r ~XzP�eʓ���v\�|� �2fW/j�)G_l��	c�̻*iz�{@��A�t���<G��:o&O��7���$��wH�����ј����O\T�#^x����nm"K�ΐ��ޥj*���/Q�$ngqY�$���ԛ�<��z�P)9d�:t:���'F%��f��b�6�n4E˲�r����g���>|�m΂"x�$cse�(_�H>uX(�+h�NvTǈ,cs#'�����9B9��7_K�
�i�b�lx�9�� ���	�ِ���О���U8o,q>��}��l�c`�5�� �����b)��2��d�=}�qU=s�̩����� �~�g��7�<"�C��}��3��&c&-�#,�D=�Ngtp�i͞���!����3T.e��!���]繤x�t��K݀�̈́c�{�^����l�l�W]_sN{��q�19n&C���e���!�%�����;@��Au	x[�yX$߾�y�����g�5�pq7�
��Rq�-�2k��y��5�A����c;K��Κ�-�l�-���vK�@�j�&-��o��"�1����I+�%���d�(r�#��.1̿d�Yy���{P61��Ovo��� _�H��U���W{-�IV��X �9��gs�,�ˇ�ѻ�ob2I&{G���!ρ�W��wwbY2«��zY&/�ܵ����2z	¼Vq0�%��>��ݯ�=+\�S�3m���[��U�L��A	��l��x�Ik��RM4{�pD"9x�L{����H1��3��<9�0������� �Y�2�a�K{�L���n��*��x�a���T���hU��{7�-����_���0�xy��U���ƎW�q�=1���;�=u��~��[��=Ĩp�c)��P�x���2�n��fJ覍\����YH2xo�-�1˨�M3*�r5�6�X[f:��u��3�`�%k
�b��dYc�՛Kq���e��k�5�����Is1+,aR[T�bK��u��ł	��� X�Qd�T�nVX:hQҕ�+v6J�CF���e��m������@��UY��FiL5V��HŲ�T��H&�m���J�B\̽uچ.{%cl�ch"XG5�{h�,U�3C1�H�˖���mfn�Y^z�4K2�>~���썺-v�����_�y�_�c��KGwL���O�T��|��C;H̽�$�7���"D(�@����{\W��r[�������K�}2I,c��W1Ly��O���]B�Z�g3-ɇ�B;�ؖ�.�$I�Α(s$%�D��O�cbz.R�2Đ7ۑ H1�����P��l���J^�����9���$���$�g�0���u�g�	d��fA���[��*w�dz�w��$Wc䀹�5�g\��9<3��ƺzLgd�`J�~2}=\��j�Q�x��VH�+	)���^&F"Y��� ��j��:�.�tI��mWTtя߿�=���k��c���2I}�<�hފ4��}�\U=oSH��yѫ���Ch���]{����SSa��.��t�O=N	� �]酀o��2��5(����g��F]?�.�/��CR	��\�7�و�{�$����;v^�='��(gY���҈�o6�dɐfy��f$�%�.d���[����{X�� �5�R�;���1,��o5��1�!9vp�M��}Պ�Nerld*�$H$��d�zܧ&xt��t�[ۏ��(A����C�W�4��oNv^��v6��6|ӖՁ�P���ο��o�`F���˿������L�A!n�$�X���'nqA��(r�!�"��qE�pq��c�`���k����)n�m�8�ѭaf+*�g����I���� U�C��d	�@���M�Dk��ё# �b��J�2Mq$��Q�N^ a��2]��yF�b=$�B��2@�&E�s�dq�,��mL�+�D��$�ctI�]Yk
���id��gD�	�ŌO�o�yE͈�̜�Z1�oӚ�]�T�E���;��J��D�K�ݚ����b~��3�XT��E=i_�̀L�
v"��\qԖw�,M�$��!�Ø�n=����yo K�=H�:ɼ�	�fIbLv�|��mw.r�G�v{��7�;ߪ��4a$��o���|���]Z���U=�ѳf�@�GgFlk��2Ĉd�[�3�>�U��HRz�p1;�b��qZ��Jq�h��8��XK����(�a�mT�m��ҁ{��|�"��@ �ѻ��G�{��O^>�22��u�U,s�����=�$�]#y{��>�c�H��jJ`��b����{^����D��������T��r�I1w�$��gV��4��td��� ���M�=�@�w/
sB�_ŧv��=t�ո	cwy�9 	��A/�q��%����L?�V���A��o���Q�,i�v�1���u���P����a��ӿ�=?��f�';�z�d�-�ɧ|#/� ��L�2d>!���~��-�8�Į�IX�(�b1��6I ����B�$ٌ�F�L�[Y85ݰ$��E��f�&"V~X��x|!c����+n�i��Ѧ�܎ەP�k\����]RS&W���{r]e����l� �@NgT�	w��)�֪~1���Gg���X�� I�=mX�ҁ}�L�s��"�ꣵ�^~w���WF�"�)�����Y,�����h:�"\zV��&-��KçxsT�ut� �Wc�A��>/�^kJoW�5� ǳL�	����@����!	����,�Ecʷ�(�c{�@��w2ɦzr��HI�@u�F��{MM3�O�ޙyf��t�@��OfI��$C*���Y�E��NV2[�d� ����D�0ɫ���"3�l��
����\�G�O�-����s[�g�E� Я�ӟ);}���6��]�����Ō�'�=���޽�fL���,����Χ_v����\]߇y#������{��=��-l���x�P��sޯY����"H�Y�8��{tGN�1ə޾��<=����>ӳw���r�Ş5	��TǞ8"ǔ�.�����v���T��>���K�縭��ͷ��%o����x������WDP�n�ܮ��	�g��{OS�A��4s����G��u�Tzugi>��K�f�/<�<\�� �������ە�9�yw�D����:)��@<��:�.-��x�(+��6u���B�;~��0��������xX��� �|�	��%����p�5��M��^%��[2���!oC�r�.�jg�����'nǹ��Rb��f����O�MM$�{$k�7"4��m�O�}i��W=ݾ�A��N����p��Z��J��P�i��*s������N�v�s��䆲���R�{z�R˓y�;N�<f�pR���aн5lk�\�F1�1!�BA���Gh�"�=�N�1�1`=]��Ý�=��m�9N�Ѻbx=�ç����v�PԎq�q��S�:uW��碜r55��=��#OyOhp{v�����Y|_?+�d}�C �r/M]�J��>E6��Zxկ\��7z6�G������_���(���&����~e�^o6>uh��$�M%�	"�d\�/QDX��
Cj�T��&��D4��런?L�H"�p�Ɗʢ`@�1���N �NK�V���i��L��)���QY5$3ā ��s�O�!�W��ζ1�@KET��6(��U9e^�L,KJ�V�����͞>߇�ۯon�����u�^�u�^:��=s[��f�ͳ�fZ(҅V%�C-����E���
V""�b�S&�Oo����������î��Ӯ���]r�Qb�?�Qƈ���iF"��mjvX\o,��b���mAF"X��DLimKch����J�A�,�("�W��"�1����C+VQX�UAUE��� �%Ee%���b����U�-�Qm
é�3�F ���'Am
1UJ�EڰS-*UTm�.am(�DCR��(j�1��C���F/��[h�
хeEX(�8ڕ2Ո�Ĭ��ٹV ���R�6�E��	a�,-�29^j���ml�����m�eb�`���̥H�hɬ*l����sZլ��ͷ5lֶ��b����s-��i�յ�������[+Z�
�M^څ�fb:
��l1i�/���R*T�v�a2i�����[�@♠�kR�/�0�[yΌ5B<&�
[(J���@v�&аn��JՅi.X[�wPCJ	,�!����t��i0^�36�m�+��3j@`Dj�5)�$��a��[\5ԘpYf]����ڱG9^,f�c(6[^E�˓2�����6Ťݲ��q��Δ�-���:V��k����")eXBdV7���%��2���b�#6`��Җ����b������HC ky�UL�-��&p��Pl�9�VȎ0�i(��͔e�Лj�dj��+Z	.)M�Cb�v"�Š�ͱ�I��6���U�tV��-��e�j쵫vqmiMT����=K�c8���փ�aV� 2�$���=h�0��+
�ʡ�d�j�45�a���Z�k���a�p�3%�ҹ�2e���رL�[-WjZ6��8��"���cU�!�v��fȣq.R�cn Rj���@�t�5a)H���7a�ԋa�
�ͫ����ź�SHsq�UG�1̍m�pi�wh�,Z6����4�f\]b)�t7��`*�.!�K]��b�����2�t�hR��-�t�]u�eva�(�pZ��r��J$!B�ц2M���QmRƉdwu�!3\�ͫ�S��K1qJ��Hv�3D���l(��sSiN�A��64�2XQ���[llΖ��Z�-k+0��0�s10�cQ6�s�8����4�L�Ⱥ�[m0slɵ�mK+�m2��Ӂqq�RY�/+�s5��{8����em3�5��±F�B�D���5m��gGl'g[���֮���T1�A����i���!�5�lQ�;4���B�Kbܺ7�����1\d7��7�ج���R��UXa٥�4.ʹ\��T����E։^�����$��S��=[kv��&)L�u��)f�<�a��H�^�e�V��X4�5�Z�sd.��ݜ�k6�"�%������MV��Uu�6�q��u,�(V�Mh��̯V�-D-Ĺ�3e�hkL�#`☆�m��	3�՗13�(�P�eLXn�"�\nv�e�T�n�)m=�W��h��(M.+���ջ������h��\Ц����I���ˋb�,�I�H\����G�6.�߾�~O�m\̿{�~�����	$n�H�1���Ʊ�D?�r�
q
@I�hoz�I�~��.��P��p,�o�� d�oL�Lh�����-��#���JP](����,I���V���^X7/������D�#{�e��jg�F��E������S3�����ؖ%� d�3��I%Wm
�����d���%�MՓp��x�\��t` ���g�z-�vV����`=���-,���F��N]�/��BS�/tn�H��ϣ֮ 8Y���2���LJӭ�`9�-SP.�[���vxr����:�]�Јp=�q$��Ap�ё �A+�d	/��d��� 컁�Iͽ�%������x� m�s�o�j7ￗ��;��c�5A�Ǯ���9��L��Y����sn�K_�p?:N��cFȃ�<�0rQ���Ȼ^��jgd2o�f����$s�d%���%ةeZ�ճ���m���çObx���w2$�w�CL1F_f�OA�m�����_{e��v4낈�^A�2��*������uD�	��h��j�>�.�����[ }�$SxA�y�B.��7�_��1�9q&j�"��ʋw�fX�!wv5S�D�H��������o!"�~l^+.r��,k��v�iW
��l,�9��v�*�w��(hA<@Hq���	W�"H$�������T���N�v�{��I��i����<�]�ЈG�~�&�Y�gz6)���ɒI�����Xǈ�w������j�/����x�o?zĐH*��H�L����b�|�O޿��"nUz�����R�g$��_��Cxm��׼�1���ѱ��bw�5L>������MS75�B
]��d͸A�{ֈ�%shdɓ 6��	 �˙LP+7�I-���	�@x	�<�W\�C\��)��bX���4�
����%nׇB���!�"s���w�)�B0��=�$�K&po��Au����bZ�2	%Wt��s�������=P�I�ܸ(��,�
�J"4ez�n�0���\�Q�ҍ厙�͊p?'�����ֻÝ�+�ᤖ!e�I���2V;ZĖ�F5�}WX�@vl��	��'�CB	�BE�n���8�%���s|��/}�<�1/��%�0�`m�z�3\���#o�����~��)#��a�����_��� �ݍ¹�_ݞ�Vx���vd�5��$�� ߴ[��0��x�Eߵ�����x	u�؋x�� ��d�`X��6���Q��]|�B�t�=�4��ſW=ٽP�N��<���|Df��s<�z�{�f��%�i����.����Y�̅�y>{��W^�̛[�ggd�|W��@W�O��S�U;�̒H+��j��#�D�	>� I_v̂�@@�����ӋeVw���@���ͷ�<��[�W�5�3ל6�.��VĚ�����2�Ԫ���>�#uq�����P �3�|�{�X7�3py��"@'ם#��}DB�]�̃�ѥ�o��� ���A�Ď�ِH$�� ��=5�J���x�8.4 � $$W��� X,�'�P�O�O��^6wt�$���-*�"_���|0n�	'DDB�w��]c��Fu5��ENĶ�V��	�
�?s�W"���_d�W��\I=�]�%�@x��8�\4�V�d?�������/ ���dA^���B��Rj�S8}-�u�^:e�f�S�w�kn��ٽ��׹u��i�O
yy2-�v���k��G��;�w����KgO����2,㊟�a%��3qH�s7��+zfhᆘSyq�9�{9,���=o=�K�7u�] r�H��l��S�܆�m4pV4!yxLWL�;A�t�ls)6؃e5c���h�Q���]0@M�ņ�9�c[I��馑�f ��ƒ�D�g�k�E��I]��l4&�4aN����M��M5�n�[�*��H�5^{1�9�!4)e�ɝ3�p���X�a�)�����S2�v�f��f�JC<̑ѻ\B�L����v[*���Bx���PK��.��p	ܹ	nl�$h	3��� �>�#1�4',UêJd�Wy"q��F/�)�׊��Ri��Ѩ�ϵ�8������#Y��) bcרӐo(������pSÙҲz%�r���	�7DV��.ؐH+���Ē�r�R��=�L;()�B����Fi�w'��d�.�H�I��1K�{���i��q�A|�H�5I��D$�!��XM�d��$esQ��f�$	����$���1��ck����*YC}.�<��eu���R܂�t�3�k��be�b�#E��b#�,�|F	xP#[Ϟ�&�'��,�	.�Rs���зY�^�֠)��HG��CHD\u����˺x����e�����~^y����	I~��-+�J�����y]�����{�7�Fm�1|��|��<cƉ��vJ���
�'�݌'3��U1�$m����_{L��g���	Dmo2dɐeW�H�%�㔒�� �#�N��ק�|���v��5x$`�N��B�� �Ogl�K�3��3.�� �I�A��H�މb| ���0�Úv�����d���U)��p� ���A���h��OH�@���� �h��8ò�� $=��0E��t�l�˩�O�ڽ��z߼��ݝA���w::��^%�Ew��J����:R�#ՖΌewe�
��1[2h�`�2M����6���>ӈBI���^^�.�Ő7ױ l�";�D��5�S��@�z�I�[@��.S��x5�{$�
�0��U�i�Z��I5�� �C�t� ���(f�wD-c�>]@Bx��<C���b��;:�i��q�>
�Ñ�Ԟ�����5H
��V���S������XQ��=�<�qw؍�v@=��xu��������(�(ߐw�ͬ�&M󀼦���fl���t�\E�	"�AB�ͯ����f�}9���s%�U@���ס�S�jÈ�b��r8=K���p]��K��&YM�s�K�=�}�ۥ=���LKgḺ ��2���C�th��v�g�rt
X�
�P���(!f�,��&:�P\q�k��S-�nї���?>O����������l���TX��:�H�U�ؿ�@0 ￦A��tw�?IDc�HȰ,�Y,��eW��]����T�4�$�sj�I>b,ﺠ4������F�,���$wl�g`��y�t�C�=7�=bH$�]��A>e�����z�{��cd�9s3���G<�Z[���ư�)&�̛��kΌ�:~nv!�dI�I�/�yH$�oC�b��3BL k�~������C���=Ս��H�����O�:��]���{�������3?�e:0��簺�~QG�6��e��Q>�K��MFz�������%�y�鞵�Є�q=��f���v~���Yg�ɡި�a�s�gZ�H�aC��u�̴�.X�?n�I��z�M�b}�s �ZV3�ɤ�ɂ��y[��[ h���c�A�15���ڱ+�\�l�utat-��[ti��'������&p]���Y="I%j̐� fwD���yt��5=��^�$f*P�D���F11�n͕�4���Jd
��I��p回:E1��a���9�>�%�����N	���Sb�M �}3@ H$3��~�������^vQ�9
��֚ ��{l~D:t!��;;���l�+����ַ����_l�K�퀪W����y�/<���uDeaC�DК͑$�����M[�����f]{�X��2X�-<����jQ6VN�=��������ܫX�]f����d)N���r������5?^qzzDR"���>��Gv]{+~����r+|�{�����<`�3ږ<:u�f���%.�y?F|�Ye7�Z����@i�i��Q���B�Ě��Xe�����U&��e����,@Kkne(�I��2�IisH�z�*L����z�Y�3��ԩ�m��b��v�l�%�Q�vkJ�hcI��u��� P��6�Up0�5e6jR.��cX�� Ѱ�T)HWc�V��0��(�T��J���s�BP-�&��le�!-�KŌ-+�&���I��2�ۚԚ6V�g���|�#��՛��7���$n�D�I�����b�?��z��+W�Y$��n@��T��O͕��$��l�z�]��VI�fD�A,g{�Ac��n�Ɵ�Tw���Z$w(AP�D���Ă���-$�U�ϗ�ʉ��ɑiMwt�
`��N	����x��M�=�DY�s����̐9��dX�	�fL�*~�ٰ��93��J���V��_�}Dr!�űb�d�U��g�q�*�>���g��$�����;�!��o�T
N���`!�yn�8�b���MZ,U�D����-L�dL�_;��D:"�B���d0�"s:$H\��AL� ��b�an7��&Y��K=a�C�hwP���a��[>�٧\T��(#���b�P�*��L�^��u�����T�3w ̸{E;�I�2@=��CK�8����������ջ�W��cl=w1F~��2d��ߚK	�.e����ɌRW���E9$�.տD;���2.�؈lE��RO)]F�]��Y�� �v\�b˟�I"$o� �J"	B����0���G8�l�9����Ia(�BǽRy�:=��r+��R*���E8&"6.ץi&�6/	[qx��#��o��&��$�,�$�E�ޙ1#���^�IJ��3K�ђ� t�\�:��!˨�˥�:�(#�D:���� �hw����&�@ ��gHIbo{�Mo��í�X���=2|0�]� �W��!��e������1�}��9G.3�2$RA��H�wL��AN�"陋��w0`�s���u�W��]��c��Đ��nb��S���1�l����?z����2�}p�{<<����zK�Q��v,��ޛ�;�1���yo�Wg���D]M�����P�v��>.ޓ<D��s�w�-�#��6~�[�1q�}��gw?b�;�0��i�j/�}|�˕��4��|����޻3p�fR�j��O��7g�e��W觴�	�T���64��G���>Z�P�W�*��y�j���`�z�F�~����ۢ�)�{R��X��e�SgAf�>[�+�<=�%��'�}'i����|j�Wk� n�p��r��I=�דg����4<����y�ޑ/4;K@��^��#�o�E���N3e��'�زc�.;����k��^^U��R�y���ýnL�Nb9.�1��Q�F�-$�3~���ϝ�Z/�^^��@��g����q�l�=<��`�����Zb�ݏ ��D�"��|r�/��`I�(�~\�����h�Gȁ��<4�l=��`�/R��8�_����`w���<�6^ S\�;p�Wy�3GY��g�,ީӚu������	�Y��]��r�*��~�u������$K�����r�.�ս���
x��s�;7*̧�w��:���a��ED�1��ރ=�Ǫ�#Aa`�Û�~����x�W�s{P^�yg�\����o��K�/*������	�a�C�x�Q�;r��V�ZU�8��Vhfx��3Ϗ����&����2�(W�x����#��M(� ���-?y5�Z��<~8���B���̧Ug@��� �N��s��}��z�5?{���<>m�w^R��"�PX���֭}�s��mm[5����T��pyK1�Db1����y�u������ۯooooo�]u㮺�>M�'%'Y{j�[55�� )�7v��E+(��c]����\^j����|=�������������\u�]u����m|i|��^�r�.TQ�Q����IE�����Um���P+*T�VĩYRѡYUX���"�\���ְ�'�ܰ�R�U*�֨T�KJ)��J�T*	B��B���O�b��mE�V6�UdRu�֦��[ki���նi�ln�o4������R��KE��C��z�J�b2EPF�6�A�Q`��`��Lq%g�,PYP*V�*��G���e�b�V*�RT���ω�J��5�q�yl!b��Y�,�����2&������'ᬋ �w{�I��I�1H�tS���Ʉ���Tv߱D����0�&����,� �!�ޢ�&7�b/czܬi�֤fE��B
�� �(��\�D�\����=��4���/�����\t�C&�����z�.Z`�!oP%��kse��0�\nq�hG�ni,���r��fT�7g1=��C�itm>�`z�Ԁ�d�gD�I$F�́���l�v�U�ה�@2�ٳF�(�~D�E��˦����&�T��8�y{2��2� ��w�P��}m4 �v�<���p���^m��d�d���%������~R��Z�d	/ݲ$����Aȇu����(��� � �ې$�H�˙	�C]�������~��V�(�/-\��������y�o11x���f����|Qݔ��%6+�PۥyN���2e��L�2o��&=~� ��^�xA�Aw�4��$γ$<م7�T�(��$�t�"R ��]�Mع�6tW��ʘ#�@��a)+<bpk�T�CJl1��t9�ڹ�q�6�-�lb���
��B��B
�� �;�>�d��ܸ	�ܤ�D�L蛓J��ޙbIk�d�U`<�䈈H�[�[���)��ڙ�1z��ӻ�/Gб�ܙ��A&k6$�H�����Tz�u��J�^�t��� ��w�BP ����G���A��� �
��p����^��,g=��	<�D��*!�9Q�U]��B۰H�nZH$~{3�/7�ە���dX��H�#8Y;�9�?��c�������yW�Wy�z.�I�{ H�ޙc��-����uzJ�z�6(�S���E�����q˞C��왽����G��G1o��?�g�ayy��m���s�X��f���)��9s�J�4�>K,�����i�|�)�PGC��ix���Et���;����t JA(W]	��ݷ\-�%hYY��~��m|�\ ^�v�ԅ;-�,�UV��=�fʫ�ݳ	e̫"���.�3�\3=U�f)�Y�1��P��ؤm @��A��e%�S ]-r%�Fݵ�f�c�j�&��16T��Mh�ٹ����Zbds6�ΔIJ��j6 ���4�z�Ł�r�]�"jks5�˰CcV�։�ͩ���S�����D�;��*;$H&�2i� a�L�w�AU^9�I�:b�b�u���	��KL��(AP�D�j�"���nS��?]`��Hd.g�H$�vD�&@���������֒9���P�tDD=�w.�IEftI�oI��v��^�� �\^H�1Yݓ$-��%�Q	@��#��dzn�/��Lk��Y3ĂA=�ِZw�W��{l=��	�����C����M]��-L��|�}>��*�b�g����ɖ&�#[����$J"_C��"% �D@��nq�3 	s�,�^[j=�݅ٙ�]a����f#[}�3��X�{7bG2@�)�fO>*3Gu��:D�X��D��=�GbB;��&O=�$��
{늅�j6U��mq=:��K�	������ϧ�ӞCظw0ǏP^OG���e���'a��ǔ{�8"�j�I94}����������ـuy��$�'ۿL�3���,o�	�K��ɉÅJ
��P���L��˖�&=}{�H�3��?9��Ăi�9�A,2U�0ZX�$̟h:�'t�D.���w�OwN�5C���K)׊�7�e���D�0���H^ݙ�]�"s!�Ʀ�f'�}2b��V洞`���}�r�*�A;���ѽ)��y�A$E{&A�I�Zo���4q.{C��Ke�#�븩 ����:���Ȍt�Qҙ�a�6�2!�Q��=�,I��b(��l���3��)��$2G\ŵ[M�&|a'"(�c1�[Õw�BP�5=t�lDf�P%���H�ZYfȷ�@��4c��4l�9B!�U1x�ly�"�L�*pZ���]��T�W6;˱;1��XCZq4�9�rLAI���o��6��gާ9"K�%�t>%�U�O�G�ԑ�2<0��sCC8���0����Ŏ�~�̐Q�"X��dm�(B�	�C�]ޝx�y�S� �����.-������..��{��c��fNp<�;�B"
A2ۺ��mo�K�}g���A�lq/99>�ӕ%�|���	�ޙ;^��P�-*�.\����2�`˵E%.�R]E&hK�͵�.��#���
,�\�N�"+����"��9����[�ĒA�ޝj	;ߡxx\#S�'��&آ[�s"A KmΟl'�x��"�W�D�/;�}X�߼3��I$)��K,�wtz���?����콗ф�)ȅ
����̕�LI ����9�O'�/xķ�.���D���"r����q�"�w;Y���]�%�\�K ��ɐ?v���8�|��{ț�3}���fL>�&�b�KY�g-�.In~7"9��k�p��x�����:~W�{u�0]M���=X���N��$�����8vvvp���$��H�L���������$Hd����O�yV^������-$���d�b�Ț�1��{Q{�\�c]kc�h0
�6���W�T.%ъY��1.�Y��gDH�C^�yBw�C�:[������U��,H[�"��Țǟt�� ��t�%����]���<G��Sc�У�K�{}W[ ��ν�d��$O1G:wv�����a�l�A
xO��շ"I_l�҃�Pʑ������d�vgcUH/}��i��I�IȄb��Ǻ2jUb�+˒� ه ����
θ�d��#;�^�k����b@��bFB� ��E��$�y�"O_���(O{�m\tɆ(�g@�8��$yH��6���(`���y����{9-R��q��/e�^w�u�ޕ��5ӹ9$=��,B�_e�9G(�@Mx���Jg�i�Z!g�syw4�w-�����e�d��:+�g�����5�f���L5��IZLѭ��ZA��s�A�V��8%b6ah0����׬%v���F�۱�%!�u����v���e�X1��Ь�$�lF�6������@�d�6MP�Tx���u�K��-�VZfj8�J�u
�Φb��8�)sYV�d\�CWm��-����X����D.��f���h5GR-@��+�����78�/ �~��$B�	��C�ϡ�+��A$���0�@2�^܈��^�7��z@9�,7{�8P��s�	ed�Kk����X�`>�"[;j���H+���YQ鞁�hQ]	��&kr@';���xPK�xy���j#f$I7���ܼMx�b��CZ�t=Ʊ�S�r66pS�x��^��ʭ���/i�x����"D���4��b��u���H4z�鳑��e}�/c�ڄ���P�>�I$�w����i�_�Nf\��_H�e�v[��&{�����7���~|g��]k��*���V�b�k����9�:���X��<13*��}�}����pE�$��� �4֟��Fc��F3�&ǣ���(��"M4��8H����k/WN`5yx_;�LK�ہ`צ�;N/��^럐~|��5��������;�{Q��o�	�.�R�������?~^����=xq���^�x�o�hgggggg��,H�I�2D��>�d�t��]	�W�_�Hv�9�yBN	x�P���1��I0�nx�QZ�5c ,�H�CM��T	ȭ	=�	�����G�7����Έ����a��4��w$���e���ui�����Y8$���D�#�9#��C��!�]����X�}�q�"���� �=qZ[��$���f�=Wp��)�D�	��^<L3V��ӊ���F�׫-Eغ�8�H�s���'�<Od$\�F �^q�B �osbY�"X���:���lV���4�����D�iD�������'%?d�$����E��Z�m��^����4	/�2��wgT���[Wq�kX��^H����R��iv\I,c���ղ��{��f�m�rp��.��FE�y����g��^:�M����ܒZ���@~�Q�g��94}9w���dɓ|��r���n̂O�'�7�uBN	w���<�i�;�vl�`s襺��騒I+6�I �����IY�7�R��y	H���O��xx%�,Y�M�c%Zΐ�E��w�����1��e�'��b���R�rf|G�s�=%��1�I�����Gi�x�srS�nI����6��RU�&W�����M�.o߳��nd1E�:E5!��I���I�w���Gt���mo�U$�u̐!��^�EȄ`@��R��9�ܪ�����F1)�K��A0�;�r�'�����7X��3^�C@�	��T��e�b��%��A@��9��֒X�jiD��H�Y2Ac�"�	h��,��B��R����n]-rH*nfH �Z�=���1�j-fl���*Yq�{����qygHԏ��r�?o���{�����Cr~�>����v'%�+ۓ�5Kք�f]7�7�,�2gݵ�ʙ-�U�Q�	ܒ�	!��7M@G~ىv�pF�������'ǹRK��2	�V�,��%������V�hA�l��8D�Arj���(ghB!�7O�Qw�E�8sɸ�J��,������e~��\<yN�e�
o�2��Kd��g��x�ދbI��N<|�w���h��TH$5wt� �m���"�?m��ə$������ ]��f˂��fı!2F:o���U�F�XE��|�K$H������C6 i�h;��b�=�o ��K�4�;�%��Fպ�!㔱/��5��T;��@B�O���핰�n�{�5��$>=b%��Ι$
޹�h������ɋ��U�şGxnY�w�{;l�xu+=@~ӧ۶l-{F��.��]���<����*ۉ�{�<kN�ülg{)����;����\8h���Á��\4_9����=��ܤ��Bsc�� <4�����v��$��l��|����<7@�Y��,.��|ߓ���w���s}�'��� ��o���G� �=a��+�Oy�#f�W�����&-�;�R�vt�y�>���\��@>���Aܲ�o��%ɝ�ڗ7�X�[���*���Q�u�o�[9+�d�K�h��\�lż�����?{�=��}7&篰x�_���O[D&��P�j�Wx{Ӱ�#����/�ت�\�^&��g�˭��F�#�߹���zk��kQ�?e��^�:�v~>\=��:�`������]��깮�w2vI<�~z�:
$tNx~�轾үoW�y���^��5r�׳vk����n��-�y��o!�R`'�����Fm�`n��u>���oo��},9�۵هM�[�@�^ۅ��/SI�PA ����Qv �ey��a/����^]�9R�8�ݏn*5�����т�����o���A�J �G{���8��Z�d����5�$^��>���7��>:{��M�[L�3"�,�	 Χu�9�&�>[r�-vF{���{����\�Q��W�e�/T��=dR>4�}6[Fw��DÃ���128�����L�\��%�g�ڤ�^jC�R�<r�lq�S��'�w~+k{u=ސ5,�-a�� ��i$�7ӭ��<�l�0�pZ�f
d��2�f38�p8����C]��L&�4�"�A��E���Й64��?��*�� �ج�H�*	��m��m��lm\Vs[9���j������u��u��������:뮺���_W,[[V��U��˛kfʶ��K�<�m����u����׷�����Ӯ�뮺믇Ü��H�C��c̥ܰUTWmE�����UTkUPFE�����*��>9�
����D����UbQD�%u
��*")!G��&5,b-h�V�K�& ���^3���6���aQb�
��dX�V��r��b�Ƀ^%Dm���q��A\w(��u�e��G)b�XnVޙ�';.�;��Ʉ��C�Hb,*�HUk�^$�E�V���e,1�PԈ����P�T�"�ME��'X"�H�(A`]�YX"�cgr�M`��
��*�CM�����������ʽr�FՄإ�rm�Ҽ��u��͆�؋��v�N��a�ґ[tn���0S@���n���\l�����l%�h��Aך=]˙��2XcM�q��n;��4��"�\b�B��hk���o5vv�GZ�-մ��,K�cS����98X��iFh�M���\ �k]��Y	�����8d��셍�ҕŬ��B!,U��	�c-��\�m�s�AڻPݢ�KʐR���+\X�Q�V�����%�Y*��9���`�Yf^
��n-x��U��S5e�G�
0uf�hk��(M4�K5,���\&SСk�U��6��� Z�Iw1j]�].-��ԅ�,U*U�.̭+ŵ���]
��u-LҢ֣r�����\ṆƬQC��)N#h��Ƶ`�"m����\X�R�v���jc�@�U�ն�d�+`Y�x�k��[���nR�]���l�3eX��n�̹˝�+.�Ջ��*��\�[����3,N���ke��MYu���44��bj̽��
A4�JT��Y�6ڲ�KP���ݫͲ��b�5]�n�b�`V\5��l\�m�p���`X���[-�׮m\�0W`-**��m��X�y��t#�A�]1���k��	��	����8%Sqq�]\�c!f��,]t��)��l��+4IW�]�d� �`]cV����-�����W[	E�+�4ѻ�cv\dЙ�Z�7�$������5��Ћp�Dt�[�(L���諙f���U�2�P�%Y�e��Y��mL�F��V�^&�"l����%^��YWa���)f��%� -�͘[�B�K4AK������MĴ̲�4�ˣ��ط�B����i��0�j�n�1It-��UukKtl\�ar�+�Wu)��9w��o)�f^����e�~�z�=k<�R9����L[�B�m�7��R�1[5�Bf&ly`K�R�[�:�MW\ۥ��n	od	[qKQ��<�kI�[��y40��U��Қ[�ɪX�9i�ۗM�jVm�PMn�.����A�i.�n�����`�*u+�$�� ��L��g%���,v�Wl&tj��B���k��`�g5���uab��2���Ku+��F:b��g4c��tyP�\�Г�J�		~�Y.I��$-�%�{�A[�[r�1��BY����V~��xP"F1���vG�A�=1WKk�Mwl	���9A���O,Y֤�󌝂u

�U��"A%_t�$�:��7�ގ��(׳"A ��wt�;$�>��A��J�
3�z�P���=	%�e]�,��g��J����Q-�2�����$���Uf��@�-�g��'}���; ��2K�6�J��R�z�ٓ�xx��S^�̩Z����VY�fԩ`���:2̋�m6N��o0��J�p��c�KK$�\��['w�Az<N�����.�R{�P�&�k���@HV7���)5�;�;ۿ�/�;�ݬ����!boMUIW챴��}����-���0gZ�'rI�� 
&G�������5s�Ӻ��nhdɿL�ƂA$���	�-�BN��7�ៀ��Hٮ>�AD(B��ng�C�ާ ����S5[ǳp�B���$�}�<�FA��@���=z�\s�2İ93�����Lc���}�+u�Ut�L�y͖�V5a ���`@��b�nK�X]�D���:�rΥ>z�l-���e���Ϻ�	�vO��χ����$	O�L.��05)�d�����CA�����mZM�tka��e߿g�~��y@��3��� ��fK88�tt�3"�ݯx��T�<���R
h�:,��P���z_�d�}ܻa`�>'ܛ=%�$��H���f�s�ƌߪ�Bj�󞄝�HMk+՞� �k�"A �g-f�M�[3�t�=樕N�ؠ�{PQ!���rwe)_o� �p��h.n�<6��=��y�F���k��ϫ3£�1oP��rKx�N��ɓ&�;+�@Ʀw�y�$���&IMuX
}���P#��}�d%��Z�d����L�{�$d/�y�B7�q�y��d�cD��u
��{}s$�$��n���k��lv;j�`$��	!wt�3��3�F�ؙA JG
�D��O����*K,؈�����g"bh�fpf]�u6L������#Ȅ^	�*S���'םH,��d��z�־o�ߖ�?[�b���2	˃u����}�Uu̖�S��Ow����$�r�bI$K��@Kt��N9Lx&-����D�
P�x��G�����i���4�$��[�3�%�+˴�W�2A ��%5Us��� �C�c�W��x/z�//3��� �B��l����Ӱ�s���h�G��(%��Q���Vޙ`��v�]�7C��/M�TN��n{��e��*�~B����4��W��مG���,�/�"��}T�qN���P""|��VU̐B��/4廬��ي�H*vL�,I]}2�rk���*bI �e��Iý���R��A�,��YeE%]���u�p	s[�n��1�6�HpS�T	�{y2F�|��#̑!���4��O�x���q�A%vd�ē87���E��zÊ����x���o]�(�IU� y�1#a���dfM������~�$sꝇ��x�TUo@q�F��D��ۓ�]�&Pw;Ga
�2A�c��HTH=�v#�����.$f3�d�OM���)9�v S%�8� K\\Je!�kK{�NZ���4~疒)�<y��d�<)�.=�"�J�r$Ǫ�o=M�v�.�e�$v�q�H�ttɭ���b�P�����)�m�b�A����r`K�B0{	�R�����!��}����0�p4���={ �>80�1a��к��0��h��Y� �;w���O�~�K��u�8��rf����%�fc{�j���XB��ai��P�F�xBP�6V2���Ĥh,�w�
[�R�{�Z7s���Q��\�Ң��.a��6�k�2��`�j�(A�!k5SP���)�;]��J�J �\�R��c5-H�̩\�U���0b�u.Mr�m�C+�lG�����M��˛v���bUS��6�R7n�j��:��nv�n�V}������.k�����w���Ke��@���V�׼�QQ�ؘ��sh�A"�#I2�ug�pS�To{��2ċe��y�n�-�p񾋽�ēލ�,H$wwL�A7��\ע�1���:QȄ^	��Ttw�H#,��(�n�k�6�9��I#��d��_�g�K�A�Wnq�}Zin����tQ,	 ��o52~�@��w����%񥡫�t(s<xp*����z�� �A]�-9=׻�a�I}ޑ Fe��[�"o/�;�8��|h⼝,H���3L:�f��]XG���em��38u�m2���G�_\� �!�y��sD�l��v$�I!Wl�2�{�z,�Y�l�����H�̙$�`�|���2[O}�����]?����_Q�L����x{�/w��h`z�{�XO�����d�Q�{{�ɫup9��{�s�������B�zR��~�Zŋ�e;	=�l	�W�t��(�6�����ۚ��O��>n�<�pS�T	}^��H_���&���
��}>��É$oṽ�}��RU��r��	�#�W�"3�[/S���L��T	$��ğ3�s�G!�t	��DOmL�q��Ѓ�������d����I����s����1�k�ɖ�o�$>�H�[��A���iwd���[y���a�v�H��@��ً1��ҍ��Ґ��=e��%Q��G��ܙ�X�H��$������ˇrk���Br!�S �I]}4��x��.�;�HU��z4���\��SG�r��� ��r,�|�' �soxV򉫟X/�%����"��<z��V�ȒK��%� ���-���+�<簥Y�$=�̓5&=X(�U�W)rV㷝�O��۳un��=�=����+ly�P��yပ�@�ŋ��j'�H$�ϤH0�?���3���!�N�AP=]^�}�b�!`�6�{�dI��$���;�V��gs��ȱ��� A�=�S�u;�>��62��f�?*��rG2Uqr$ӝ�[w�d�@E��u�#|� �WQB�g�6��n��Ɨ:65�*���቙X��݈!���O���4�>fD�IY��2O4f":�_������"y��]�l|%��Zl`J�	D�,�����I�ͬ�Dd��KvH�$�����	�g��<�hYĩ,��mQ���n^ܻ �!���k�Ϲ	%���=���G�x�U�%1$7��H����D@xJ!�Cǚ�>�}Jx�����$�\KX�[��e�,
��X��SO	�í`������8������"T���I[R-��^�-q��_�9��k2���ۇ�%�{�U[ä
��,Y>�O�D������r�V�z-�!{�1~�*��b���ZA9۳#Y K��bW?{r^����m��,\�	��+%�4�:j�֜һ�qcB�]F��fԌ�?>�^�b��f�g�Sϑ��A�݁ �)wt�8 >�p}���J���**d��bX�x����C��j���m9�؟T�����,Kz����@���- �땚����u�����\Db��d���X�^��?�clpђ����X��� �WwL�UG\��vA�B�����7s����l>S���=ĂI[�6Ɖ~E�dA���K���c�/�o/ʹ,�����ߣ���$������N�J،�[/�X�ߣM_;�Yo\	cA��N�3�=�}�PI{q�3=�����z�����=�8�>��-���{��W��yON�瑾n�u�;M�����֔5��#?{��DU��[�W7��J|�M����|�q�w���S�R�]J�#6��Z3$�sDF�jKz�0�%���7P�5����F�)��´`�+.�@sM���4[��0\J]����+�.BjF^(Բ̓m�,�9�x+ihWf���a"e*�"ԅ,k�	�Mu���u�hK^�� �aL*FL��dBYV#n�%	f�m���vqf�Yg��g���2���5f0Aiѱ]���v^�c��۬
��l�5�&Vh|�>ߝ�5T�3=r�B ��Ι$�B��Q�%���דu�KVz�	"<&�.��]D���t{,˞����zb� �'�lP ���Q�H3P+-�Ǻ�h�7� �<��j�/���.��d	�����\k�I��ndWk�bGh���."
��ӴvF�>'5D�븐	�V��|�A�����ʁ�%�����1��h��G��9vA�B�����ȃ�=�������}��ì�ޭ�`H+1��$��.�C
��}����z^�Μ�S�zk3�Q�4-�hub�+5�	n!::j��P1
kCs��i��H��	`_����rc0`=�a�@"K�ٓJ��{�z�'�ib�24�2����.!ʁmv!�ݕ@�7�^����������3��d|o������qY�������$t�7�f��Q^(@����no�lg��}�*#~>"P��Y^���H��,Y���И�+��d�%���X���/�ټ�{v"q����Rx�*@��S�r$�gD��&+/z�ћ��j��o	e�F�,	��c瞸S<���*���x�ョƥ���v�OR<���ft�$�M�{>��(��B@���t:�����&H%vdF���j�=���oL�A{�9��{;}�r�R.
\��(L2=�����k4bW+���J�3�嵊\Q��2�a�/��� :%���o<�,IbA,J��+ُ�պ�1�Ҥ�1���@��}��������=�Jx�m�+P�	�C"Ko_Ic �WwL���۹����A��k�Ä(
� ���$wL�H��ymוw-���B�^�rZ�?t���.'|����z���N���{:�JbѺa3N�Z8�:C��0<fXTL�� @���xn���,����7z�;;޾���h�1��ڽ�ܣ?	<;<�=��}�n�3Ь���ǖ�P&m���w"��3��į{ݣ|X�a��;��=n�4�|��Ƃ�ˤW���Oz)&W�r̠	4��^z.>¸���ue�R�=��m�Ou҃/����5�9./!�f��.��R~�岸�|s�ubƙ�8�ˑ��C=�ǂ:���WG$��~2��&�������7�������uV�ӽ�դ����Φo��o����X�+��+<_��3|_����k�u������Zy�������]S|N V�F��{��ݏۼ��$i�c�Y��������~ʆ{�OG����B�?�珎��~�v���}����-z���*�5d�ך�;�Sa�&�R��=I�}��!w���<N��<���_jy�&��_x����z׏;p��bS�����Mb{�j@wgg2�O��vݓX7�z`�����K{��d��"SI��|�KGO_L
�̺�	�H������u7q�{�zU�Z�QT]����F�h��'N��Zr�d�E��t����Oz�}w�ٶ�s�n��^3�+ж�yz���L�{�wޓ�絼����=�&��f�w�<�����`�G���@��/���M�Y]�}�3rw7;d��|p��{,nO��H��Jz�g$�	��b��[յ�oZ��+;�ּ�Ύk�9y�>�o���׷�^�������n���뮾>9�k����<ֱ�lٴ�mz��V��sV�����W����|�.��������������u�]u�����9W9�m�5EP:����X,6�J�TPU"�nP��B����!�!QTF&0�Q�si��*q��B(�2��%�q�A1����`T̰���Z�E�IEdX�+hVh���^��l�աJB����!Ԃ�k"�B�P���U}��QY*V��5*8�VOY�E%DE�ʥ�7Y*L�R���VE�)�c"Vk1�Eh"����	�������+1��
)-���`�\�,XbJ�
�r� �,�8 45��L�>��7^d�]�H�dޠI�x�s;�������`�y1������D1�N2@GfH����ŕ4n;��_�$�Ēvs�
h��	�x����I �-�]��c���~�d=s,H!w�n�1������'���^��{�~K��X��޻Mr�%Un[���\��Ρ�.��3`7uk[��V�_?g���.�Aq w2������@����~� �e�P�|�Ƨ��$���]�U���!9�r��������&S�:}�\|Z�TY,	���	�$ K&m~�&Y/=���}�$�)�_BP�B��TW1�x&"��)$��n=�~�S!77M �B��R���ykx�{�z�ү�ih�����(��bvHح�$�,��T�goH�gmuz���u���6U��h]^�ɮz,C޼ۭ�Y�7�Y҄n�K�4�z�|�@+����-�_K��1�=X��x�C�*個��$|����uN�"3�2Ē��T�Jl���/y�X�+O�Zg."}�������aY�P@jJ˅����7]�\׵�ka� (���$DA����ZA+丆(v�H��,� �&��q6���fA��ؤJYt)z�q�0���1�ϝuLI������o��X�W=�d�-��얻�V@�Y^�|���Uy:~wD'& T�M�;v_D�(2@E�^�w�p��{T�I��$��,�*�P�
��o)�׃=nI�QR�Y�={�$�X��Mzjj��ޡ�,�j&�d���:���{���/��T����L��:�R	%���!��gg��'�3�<Tqz�N)��aDx���ߔ�s�0g�W�·��h���zu��j�)}��Lı�A����:=Ĕ*{���eЮ"8`�fk#9��T��1̷��c{�zu������,�k��[�����R�j썆6�K?�
�cf��bЋls��U�4���.Z`v	���R�^V���1���99%�� ��Yo,@��i���Г%Vݥ��LB$Ũ	��`ܘ�-���n)`�f,�i$W,Kp�QsKr�G+�[z�P��̎k)h济1�L�����\cme����_<�O|v	F�m���5t����75j��5%�&Q��2�?���?�,eL���������y�ɒ$���k�x�y�|l����K1"�:dV׷u$DA����$�Ŋ�y��u]J}�,H&�:dC�t	.��ê2�:��x2
�q�4�}"e#�2A ��j�ʿ_�Q$��Ι:����wHE�r��N!@B��zjͿic��H33� c$	2�%� .�q}|��ǖed�rdtpH���	B	<�Ɲɸ�I^� ��=a�w�~8�	��bI/��<���N��a[7�	$�w� ��C�H��+Kj�f�����fL;�ͭ��-�7Y��z�>w�Xh�P;�^ɐI ��fI ����E񨇏{��Y�"�[Bg=#��&=2[�3y䆳�
��kZޞɦ$�Vh��yrg�l����g�"v���x����x����\;^�٧��-`J^-l�w����'­�#o���2^_�2}y~�&��[�2d����H$���2 ��I���_҂�����;t솶易$�!���x]s&;8\��$�]�L�'v'� ��P �G�x�*��=I���C��/�
�w��S�Y�w�O��8>1�L�c�s"�jDz7�I$��Ɋ�^�S3��N�L��!�x㗗tBq�
���Hz�bx�E\~��H���4�[czy��wdę�uV���q6������ร�p)��F�.�ln�iV`�ʂX�(Ki�vP�Gl��X2
���J9���I�΁ �ds�%����F����9=�K[���Y�OcP(���T��t�b|f{#��U�a�&����%��Ζ�d���D�9{'��S~����[<@�a<
���b׽�$s$}��fs�ꑾ�qN"�~I�7��絸�#q�3��oi~3�x��VU��ɞ!�_gg�z��KFy�&�*=�3�o1b��OĞ�ImϾ�"�j�	�!��
�����T��E�![�ؖ$O_t�X���R�����P&��-#�I>��ø��������2��;=fT��I{z��~�H%��AvH��٘�H��y�R�@=
_񵤷(�M��:d��٪��r:�G8e��I�;���NC��wq�o&�X�;ٱ,A1ݮ�"o6�N���y"A ss$M6G��ä�sge�7}�z%�e^��7�ؐA����Ơ��Os�K���z�H>��&���E@�߽� �#�fA�G��V��l�dh�A"�vd�I�떒*n]gx0�'�T�<���zOcǫ=K�F;��d�=�O�w��Lix�zt�U\Jr��21ň��=�]~�^G���R�c�quI��#�q#|��<�n?<�	�������9f�}J2�C���"I<�ŋ|�>��e�irAۯa������W{�e�������
%ڙ{s:dH3�d[��L��9�}%�T������N�-�{IO[Z!�5�`G#��������GF�U�D� Á^��;�	Ɉ;�߽"H�܆��`��·͝��زc$H�H�i%��Ot(I�wxN�*�G=�"r��}��������$f�b[X�V�ɐM2��3=��`�ty`�D;�&P���$�ۯ&X� ����:n�����s��R%�7�-,v�$�$sH��l �P=-F�;�4qC����pKO\H$gD�$����NzW�m�UFk�;ng�)��Q
5���DM��I���gI���C���$�{bL�"�[��z�%��xM�]Tq�Az��jj&o�~�@���~�s��pݾk���}����䟊=�/�!;��5���t�iב�����>�((y�71�r-�{�w�����Mm���&�6�R�ʠĩ[��9��XbؠgT��╌�s�e�-�b�L�1�1.�����[a#֩k�u��ı[,j�)��3�cX;vI���f���k�mi�b:����r�u�-��w!J��T���D��8�P�%�7�nb�h��
����w��ؤ�Y��	�V�k���H��F�ɵ$�EW��k6V��&�YGQb��"��#�>�ߌ Iq;�LR��jE�'�y2H%�7�4�\lBww\tl�X1Si����B��2L8�`ü���T�{�,K��O�n�vc���B��,���$���/#"�g�2����Q�	9�	�Ǽ�K䀁>n�٦)�1p�f���� ����XfdI�@'�ze2X��8B�˓(P7v���K�x�h�ca�Qc��-ד>,)�������{u�O+�7 �j��a@�����%��9��=� ��l��oy�D�9��@��� �ٝ	$�"]��,��.�P"�~�����2�w1�L�RFg�8�5�l���è"�V�:��(Q����� H&;�e�@��}Y�=C�wY�2"dH$���2��%� Iq;�LUvĕ��kAJ'g�'�ˤ�xT��4�k�{�[C;�wـ�l�lt��[����{�!�s}���k7���5f&c���j��9�2�bžU3q�I%����y��ƾ�`I�(�ܷ�����8=��Ɉ=�ݹ�A&;vd�K䍣#���{��A�̙�d��dr$�F���˼(w<=�=��Yɢ�ׄm�$y�����āގ�[׳����*�p��$f�%��%��)`�(C×x{b��4ɑge�~�4,�g�����~��,H1�qm�3�������lz��R�AB!�.�T4r�6M��$�^�J�2i�n�d�3r���*Os�e����T;����d6�B� �R�M	 ���� �R�"u_��T	d�̑84=�V����B�2c�Ȓ@%��`�(��$�Ik��hj�Ig��	��^��~��d���$�hN�y��ܡ$�ϻH0ɖ��8�2�>������Z���Fz�ys�a���*�t6,�l;WJ���V|��)�}�(�^E:��]z}���z��Ȳ �ibž�y#�A�{�i���$����x�NK���Phux辮�"��E2LHȋ�i�,��|��Rq۝܂O�je���"
wB'�n�$�N�:t�xZ��^=Q�����-��$\\Ȗ0�����y���s���A����6�����(F^��.&��.GF��C���s؛?_G8l�.T���̊ɰ!�>|����u�xx�;������c'���J�z��S�J�V��2I��>َ${�#�$�O�"AL�0�2����9���O+����;�!���1j�0��$yؚ��n��ũ�x����=�%�{� ��s�`�$�Bt k]�GH|&��(�!��d���D�A��̳e.6;m������yc�ħ�|�j�[�	Hۡ�9/NF�Oj{X�`��00-��Zf$K�*�p�<Jo��!�z|�z�|21����5�ŋ|���^��(��|�b.K��Y_K7љm(y�\׵c��Ϻᝥ�flI$�����C���y�O�z�JĈ4=\�k+Un�-�����6�Z�]Pk�sE�Z8!�&�������4�P!8�׷R4����e�nd�z6dC#�W�>������s̚���Pw���T�m\�����<@�Ȩ��
	ǌ� ���	�����J��q'��c���I�'�9���y�d�"�3��X���vݭ�~�ĝ��K�;�Zj��Jw�Q��4tt^�͌�ށ�Q�=I�ԲY�1 �$A,��e��%���g�{��+&�I��ۉ�E��߉�C��"QU�2�윉b�3��~���@�5]!4���q���M��=?������y�\�~������O���m����%��R�'�r�yb�����y�EƒfD�L#M�������Di�i�jaj��#M�������(jajF��MP�Di�4�4�jF����i�4�4�4�`�Ѧ�0�L4Ѧh�SL4Ѧ��V�50�F�i�L4Ѧ��i���SF�4�Ma�-0�F�i���MM4i�M+LZa����h���1i��4Ѧ��i��50�F�4��F�i���0�����zk4�i��4��F��a���b�F�b�4i���54�Ma��Mji�L4�MM1�Ɇ�i�Ŧh�F�V�i���0�F����i�L4�LZa�U�h���F�i��i���4i��50�F�i�L4��F�i�M�i���Ҵ�L4Ѧa��0�i�4Uf̒�p����V�J�IV�%i�Vl�V��i����i�+ׯ�fQZh+5����%��,ْ�c5T�ʋ6b��+�R��N�`�l�T�f�Y�4�f�Ze�1J�JW�yO)+32�i�+L�Zj*�U+5�i�V��ZoZ*��8.1S�9b�4��F�#MP�Di�4�4����T4�4�aah�5CM���)�jF�F�F�F�#ML#LQ������5|}j��o�d�,ȕ
�M���~�����������?�����?���?��������`< ?�;���I�����쾿���ꂈeg��Z"#��֊D?����W��ʾ/�_��_������(���������x���|��������_~������5�7-�k@�5���[*�hԤ�fRMb���e�+M)Xʕ��j�Jե+,�ZX*ʰU�Ы*�U�hU�hU�ҕ��VV���IX�*�jJ��+Ud���+I�V��+TЫU`�B�������e*�%Z�EYYJ���cIVī,J��U�[TR��b#�/�Zܟ�����/�%P�%EmJ��U�T��~��?�������j�O�T�_����QW����z��u�Կ����W���_���|_���ꂈ{�ܯ濏���_x���D?�_����ο_��W������_�y��H�j�q��r�����V}L
?���i�M+>�(��a$Q����Oد��}z��~��.��yʾ����}�y_���J�������~k/��5�5�9��
!���\��?��uz��W�ﾕ�[.�z��U�_K�9_�O�v�������/����_;6���~��_νU�>�y_��_g���g�D~��W+����������?��k������e5��AV�W-� ?�s2}p"5�\(N���N��@�u��@ h��P(ȶ��24�  j�R��[4R�CZV���u���� �R�Pt�iTԶ��fR��l�jm$ V��
�R�"�[R�YP���(���4��F�Zm��!@)J[k�                                               �^� ��Q��J��t=�xƊ�` F�fӳ(W6��5�E!VZ�  �Z�5�Bta�[b�  ��W&����AX �r9����*�nU�P�K�p�, QG�� ᢾ��}� U�����|���s>�B����ٶ�2�    �        � VX�{� ���}��`����W��y� �] 4{���Ɗ����y`}��`��O}�  x{��Ъ�`�m[x   sG�j�]w �>���U,��0�76�hS3�p��s��;��g�*���\�k�UK�X|�(*�Z            =�c[��>��yuؙ���r���-�+P���P����m�cK�w{����5յ�9��\� ��B�r�\)W7vV��T��  =/�J��3]5,n ��Q�#������m���n5��˘v38 �v��]N��r�sme�݅M���)T�B�UU���   �         �ޱ�[���K��m+m��驈�k��Ln weV�˻_]Ҷ����͊sn�V6\�*�� w*�mr��l�s��(Q{����>� >���[�m�V�jUv�\ J�f�m�+��q���u]�4��Tٷ eն���V�cns�f���J��;�j�->���O�  �        �zҭ�3uY����Z�;�ҳ2�n)G�< j�d��4��9h�R͢�L �UVf�J��E_Xa@��   ;�_-QQ,ڡP` m*��5%Ue�(��@�5r�R\ ���݆��j����BV�/m| �?L�J@  O�bJUM4�&CL�iTj$�4 FAت�f�� 2 T��i2�* �M$�*�  �����~_�(��������m��ʕ�Kt?T$�	'�L���IMHB!!��B�� IO�H@�2����~?�������7���h��owuS	��9{���R���iLIe��L�u���Jj����*�y�[�^V��Çj��cn��Omפ��-���0ŖN<c�m9��^`l��h�BRXR{.�kXъ��yB��T�\���qnJ�� ��)W�Pn�N]�i��n���8Ѣ��~����[x�۽����h�),�J��͙��v��{CK����-�kSf��v$�l��Um͔n���@v����Mނ��3��wfe�c�,�#LvQ4����"fP�3ꗠ6�[�����),+ ӗم��;�B�	J���	B
�W��*�WzJ"�-��&\F�e&]�M��x�وv�rP6���g
Ͷ�LS���J�-;;�ܬv��"�j;V*D����]L�*�7�";wv)�&3uHϓɂ���e�ה�s�-��d	
�6U�����!J�+F�p�d-B9%e�eȬ�ÿ:JȎY��j܂޲�IK,L.���*�3����d魚�����Y4�	l�bnn8K����mk,EW�N��z6���1��BCNе���eH�+���^eZ4Ϋgt�ӱM��O�����<Pнf�i�-�q�+p\`T6�Q�\$^l.8�,�tRj���¯N=(��r�f�x���3n:�r��ƃU�͍�[�kV�+�U�V�0MJc���Q��Tsށf5�k)����%B�f�Y�u��}��²�הF���$�%��㡱�Y��2��Ǧ�/!KEme�
m �Ȕ�ī'(ق�R@�4���.��,+*�a]ĳp��gK�i]�{V�6v-�{�,���O!j�j���($���j��k�]^:�a�̲��H��f73&]Ƿ���>n�@撮��}6�(�q�y��qcsk-^�*ȼ�{��w�<i�#٣Aw��"��zM�-�(\i�x�L��\wQ]m�Ӣ�	m5�Xȍ����^�m�u	���3�1�IA1�N�Ox`sq҆h�xsK��uJ�7��iL^��˒,�b�(D�N��u�f���O�Vb�b+���i���d����e�"�p]��۲���]2�^DSۚS���l�x.��+��K����^�v�H-�Ҩ򠩀�Ү��g�V�J�E�i�3n���=
[�fh9NԢ���BY�"Z�|���#�؍��4�&�`N�]ڽZs#ֳ���Bf%���!*��v�=k$zp
����]�`�d(b�@���r�,��*n=D��b�^,~N]�
g��ےB�vۗU ��=�îRa4w<ѥRM[��n�����`���-!W�T�խ�bnJU�6q���r�Ԑ���D8h6�on^�tj]a�{��V^4�⁋w��'h��=EB��:yebI7�Y���\yx�+f��Rbfԭe-؂M�t�?m�;�=w�P�%�AT���]4bݙ�,2����c�ۙ�M�W��wq��&�əV���j�R�9fbn��[yl�4�zP�G!�lN���yL�.\�X�<���R/	`�nU\f��"��:�4��0�e4�C݋���<Y�!e3�+VSUr�h�f����U{��j;����ʿ�?�Ea��v")K�XC7u<����"�
��@LN�Y�
G	u���q����D�G�p<���;T�6�Xn����V��gJY����� p+��A,�F����(-���b!4��6U�hvf�z&�{�HV�Z�r�+�获&+N��34ֲ�}�Qc��V;�F�)M.���D4"���.O��+6��$�����b��k��T�fM�s\If]�hD�GR�CVѢHNQ]�H�g�����.�I(\�Q9�^V<oE�F\ ���qVz�{Y�j��+N�m�Vv̭b2�%�n-��8�#B��)s+0ٙnnc�Gڼ 
v��O7O��:���`�%^e;@e��nl�R�80LVp��Y�$2����������W�A�kp(f�Ѹ���y�P�̔�a�y�yh��Y��lS2�Jϳr���-иRfM�JN����˼��WB�
 �-�ɬn셴��ѽj��xұD-r�ڶ��Ӑ�wV�˻w4�g0���xX0�M��x[zݚLM�oYC~�&^�h��Qn�������v�gQXmCv&��Tp�)�bBs\���Jm4�����I]Kj�w�m��7�0�L9�_��������*y�p��Xp�dьZ����d��e���(����4�7[�2Gq[���νÎVN�3�H:Xh��Jm��vحZ.;�V=+	6v\U�x,���f�̒��I���fјE�<��)8��5�͉s7#a��F�Ud;	�Nk��ɷ�֘�Q�Vy�VnTsv�Ʃ#�ʂ������-�Ei�n���i*�п���3��u�B��%%S%֊��-���ڕw��S�Ц0��A���n�%�W-֛Dk)]P�y6��-����C�f�`K�@���2���*��ݺ�Pnmc�,���L°n�-����v���ꥲh���`-ض���b�Щ I�ݰ�/h:��	̽�'3Y#2�L��[��7I���e�c��z�`�Q�p(�Z���J��'���� d�7v����%��]ǖ��]�VR*(m��nJ���,'���0����(���Ok*�#�QX�t���f�y��ʹ��EG���)"�V�&��[�x�2����m�IL���!m��6��A��[��.Cv�#3Mv">�,M�r^慘(�M�z�ܷ@�V\��aWWx��(3,G��>I��B�+������~�+E��/J���a���$��n,
�ڄb������
�aۡh4oN]����,E&(�L�
�Ǣ�Ѣ�b6�P��6v�R �K
���NH�j��F�6��v�� 9nX��/I��Se2#yB��P��.]I:��U5o��!�lѧa�ٍ�Ȕ���w�ClaD[,r 3vY�b�vV�ͥZ�Iɞ����������7����(���nV�-b��CS1T{�j�6�R��i�#�z3(�W�$�Wu���:�Ȯa$�8���9���EGs�N�m�2��^�7#�An�H5�]J��[xt]��I[l��4��Z��,��sh�R��5	�f(+kh���eK ��ƔZiOh�b�eÅVK�̀d;�PaY��un�w5nm���`ɥU��0��*J�43��A0=QP�[+ �˔f�.�p%�Ic-�
ش��jJ̒�`B�)8��.�]9�����7Wo�A�����1��z������l-5�Fm�ˊn�Y�X�q�X~�<W)A��C���-�AE�������wAz!��dnS���J�n���F���J�hn;�-,\w�?6B��ҕHK�˽�{���Af���ד)L8�F�[E�{���:���nf�@�7� S0�
	[{�D�i-)��/,����֓�Ī.,��F�2�XB�֕���J�[�,���Z�;J\�qYͺ�1��l�{f��1(�ש��sr�z��r�ø��!h�>soe^�����P�pQQ*"U��Z�R�nju`��ҷ���S�f���ôCyb:���#�k�{-���̆�bX�(^^x����ʎ	��X���#l]ߋ��d�C�cv���GqDt!m���[gЦ�s�6p0c����mˎ�E���W:��r�5�p�f���*S*��,�JPdI�� eak�Ch�T,I�����%��	�r��6=XHq
	�8����������A��6��f��7�1��ԕ��T���j�9��d�)�Pb�ٵ�b����{A�"�C�-^T�,A�d�E�H�t)k��*�Zd��.�Tʋm)��̭t6���K�j����a�R��n��=��x��4ڄ��0�R,� �73`5��p�hJ��d@�PW�P{N���3+lR��.�Eh�bw1�5Q��Y�v�a�֐�T(c�ܛ�4�̸w�&�]�ҫ$�p+�;�_kFh����D�P#_�LV�wm䱖n�;� �F;�t����m�N:�Pk�蛭ܙ-�Z��&
�Ykl*С��e^c��*�S�֛xD4�ZڅU��V����b�Ƽ� �l�rY�^�#��0{"�V�%�دH0×���fՓe��v�(��j��$�Q��`������U�d��͋5�"�+lԕKan���&G��+��275�n��FR)i
��?k��w1�c!<8�βYOo)9�Q8C{rٌ��m��&*�|���R+�d��[ǈ+W�����(�-�!Yd�6��ʸ˕�n9��2HVƍ՛�������&���ou4�=)�1�̻���9f�۲ݛt������dۘ2h��.�������*�Ae��5�`*����e^fMf1��&�P��/4����j-^����Cj݋�n���U�/JQк��h7�3(��Â���D�,!,o&�[���Nb�5��%֧{x�����7���d`+��a$ZI�ncY6V`����8��(�4�#f��2��p��T�;�X1��-�Na�,G�@��
r�:F��"Ѧ����c	ڙ�ɍ2�<rؕ�t�ƨ�n�,�U��ׯ/�l*�\��CvZ�#6���+qT1Ê�O5*Ts(�1!�\Jaj�����z����d��J�~��%F4����1�ٕ2m��e�rT����f�{b��p[�y�P����J�N#�MV+��Cc  ���G+K�ە�u�30V�:H��&�@F�cʋSP�6<Y�QSHje���`��݊��V�@m����&U2��vV�v�e�h�$�7M���x��U3t����$)�e���kZwy����dk�Ow_�j�VD�Oƍo5�w}7+�J�K
����{f�q���J&�!oU�5�դnʍ�;��WWoc�uoh2
.�P���gM5$�oC�e^F.K]g�?O\��0�=DZ�ɦA)��d)G��U9��yb�M�¥�O�<��f� �,w�WۍF--U��̂3O��m���-�J�1ɦ�8g����b��p��=��v)f?:�N����i
����	+I�[�`��^��#2�[R�$��M�a�V�F�5�8���ʺ��D#>��4~-�!AU�˻�JO.��ko	�F<��D��9�^��31�v�<����T�I����s.b�Z	W�Y~�屋��%�N�ZBn����X���Iʘ��l�9[��䦜��J6k<�4�e��X��Le�j�h0eX�rI�h^(/h�2��3C�孧Q
o��Cӻ��dE;�G�V�[��ئ:V��AL'��M�Soq5C��uY�
�O���Srm��*�5[2�׈�ߍ�K!��UvQ�c�3���V�*:��"�a2��x�Kj���b�ٰD:$n]�Am��n�XBw�&�0�r����[E�+ũ:�Xr-�S,��S�w\wV���m��s-A�8� ,��4U�d��� ��mbӲ����I�Pd܃w'o5j�"+Lͺ[3p[HkU5��T��f�غ�NR�$�%�v<ϲ��L�3�ƚT��L�n�F9h���i6h�HG�n�{�P�f��@&%oR��4���&bK\�B*ߞ�/X��D� +��;��騨U�-�ۺ�1��f�5�ffmZ`�7ij���(ȣ-���-`�p�
>Y�neթ͂�knXP�0���Mx��Noq�Xڬ�)Hdw�p:�;zi7/&�8�1����32�V7�d�����XSBSE��.��Yb��µ��/+r�ܳy�����	U�ܶۖt��K0e(�,���//Ҳ2��Yu�Z{@!V�nX�yaBd�n�)�{�ZpJ�5�葘v�	��bxfѣzbq΋8+_k���7���n�i�X��	^��[���L�������9=����nn�w�Su)؛�0CeQi��c��G�*��s�V�޶*ո1�N���>�wr��E<dz��D�c���9U�z���Teʲ���Z�c�AhZki�F��p`�̭�"��SFɲp�(؁`�3.��Vز�*P�EVE�yYb���D��wo+Y&���Ĕ�8��CWRZ��E(�x�L�L�E��X��Ȳ�k�.��M���X80!{�ose��`fQ�Zn�5krPRHҼTȆ��ն"��6b��^���[��xHm�4cv�ś��]j���B9	t:Y��ۄ@q4��&�Nc�e�چ�^!L����F��-;�"�Y�եf#���.WP
z�RGo@�)�,�sT��j�yY������u��ѫ�N��	�R�%R�n���s���N[*��W��H��Tڛ,d(�:vyT��:�]V7qV�cE,�s]��%�N��5���K�
�<�[{$�l�Ǻ�S��cb`l�
u3��ϋrϳ��R��g*��V,j�A*e�sv���B�FI��
��5WR�[���ݖ�6u�]12�h5�Vj��������
������Nŭm�G�b�ƘSn���ooF��ù+v'Q��I4�b5e-!r;�av��˔VX/mjL�4yGV��F���yz�%O�Ā�Ylrl��SU*/=I �+�j�Q&�kMއ�a���n�K��tjJHf�x�b�*� .�/��i:K��9ܼ���|���=a���B�$��X V�A@ I���@ XBJ���HI*$�$���HAHIP�P��$�d$� ���� H)$"��(AB, P	$���BHA@$ (I*��$�B��`Ada��,$$X@��H�	���B,$, �*BT��B�$R �@`� �B�$��I�� ) ��$�!
�!Y +�R@�,��XH�����$�� VIB�,� �"�"�@��!�(HdaJ�$P�+��+ 
�AH@�	$X@�  �H�	?�!��?��������_u��C:�텬���4�wn	��V�ns��U�G�gc�P��ɚ�C&w'�Չ]Y@� ��W�W&7"���`ݻ�0�m�d�O�jek������:*F�%v�g`�������ݤxK�Uwz�Q��}���z�Hw#�1����S���kאYT�f�����G���B�����'8f�RR,�:WK�3�rYQ���I�e��|61o��@k�<mKW]�3/8��u܌��Ĳ�z!z9j�;�<O%v�yZ�Y2ёd�Ⱥ=L9^ݎ˗����f�v�Ӛs��@��1�\�pn�Hn�Ty�����˲3]L�f��sn�M�}a�s,å�Ƈ�oY�i��G�α���6kU�7++
z����og)���ѹ)ecA5e�.^j����a��T=Flwj�U��z��9],Y�b�W�q���0��&�A,֥^JÌ�B$�S�ƹ���f��xZ���w	��5{V1�R����;�L�c�6���	���V�ZY��M�����w���\E^��ݝ]������r�>������J{|������8d�-9�`'�s�b�Y�o5�|�u=2�^h01F!%,X�fӷ���m���hP��f�o�5�J��:�t;[y+�詟	[�Km�zlbP�R$^�N����p�����R��3��t^�KP��륬��F���^<!y�M*Qp��\ֺ
]*��ef)	[y�� �����o�p���gv�WZн����S��V��:Ks:�8�\���ŝ�6��K�޷{�j�1-�˛�[�Jc��s�!:QI�5�Z��g&��iN�)]� �w$���z�(��qBuAj��npQ˨)uZ����T�Y;��q�N+1L��̎��ƣ��?_1�6(7w4�%�!VVf���5M
���:��|���l��\�;a9:�׸��16�(��m\���3Bf��iزF�]ɪ{W���ck-���;��=X)�dGnhe���̛ǣ;@�`3��q��3+=n2UK��%ך�5G
���%<9�Z��ע�{��S���b}T��D�!6�Ar���% v��3���!n�'5�����n��t�/2���+}�=W1#�/�S0�ދ{}���;�rx�}����ȕp+T���wȡ+-��J��n��o�%����-�ӂ2:�em1��f�&o���������睧���r]WaN�ji~T��~8f�h;Uj�D�ؕ��wK������]��Qz�ӁA[�Pj�l�//b+�!fOt����y"�P�n=����?!���$�E_kh����|z�p�hf���L�]����J�����Ǥ8�	>N��S"B���<�ѣ��v]v��у��vb5H'�J�jM
f�Kz{NR9�z��e��)�˝����.����˧4�j����� �lc��Wb��F�c�*mY\w�bcH���*��yQ���4n�ת�뷭͚yX��k��������u �6a#�LpS�㻖1Q��
رy��>eA�r�h×�eaGA��&�
��L��6�L4�}/���Kg�#�QlU�i8$�!\�t���r�
h��GKe��S�Lq>ՀQZ+��<�W{�dF�^�h�C�ׇ{��������Kbkb�=Cb	d����5��CF��B;��&��hgs���v�ō�-َ뛧��Ww�s���ъ��;�����y��Q�@�Sӵt�\v�E������t�ޙ�2�*����b��s�qZ���������� ���ʘ3()L��
;�5�e�����1w�����<4�IU��ۥ4��ao�:'�hL�m��
(��6������4��`��f�f�js���N��zm���о�E�Z�I�z�)V�P�Q����� 5��.���7
&�����kkC�f)�y��!w�hmم��K��;�sQ�Q��z��nLܣͯ��=8�)mnG�k��ӎ�Cu:�c���*<��ͽ�U��g��n�d�ø�M��*�j�s���۱mk`εg.�U� �n�Y��@D���Hv��Q����;q+	/��L�������x�,�$5-���[���ajYq�����:oH}n���>B�wB�N��VvF8D�PǬ�䊮U��� ��~;X�M�k].;rr����Ѣ2i��5���G���b�����g����yy��w���V��x2�y0�!B��Q��4<|8r'i���r�D��k�C_�A�:�d�n�.X��̫�lZ�i������E_��G�Jcny �?\DM�5�+$zb�]�͠�O�:��k�-whgd��`�s�G 2���l�o_���];c|�:�-�a�Q��b��X�<�E���jޯJQ��,���t�f�	h�,�u*�י���Y�$��<g@�:^9�b��["J�4�p�c��a�m1�W�y%LAͫ���M���NWGݭ�b�sn��R�����J�&�T�óA"�J8gP�ǖP�����VN�J�_O����u�R�\�I��Ձ;�]
�z"G���^ntI�m]�Y�vk��#ζ2�l"�޼�2Z?g�.KX��oM�Z��9\��1۝�uC��9��ֹ�WsR#E�����i����P���ʨ
�j���{��*T|ďw��G�Y|,� ��^5S8����q)����2�ejnu4��5ñ��C�Ӄc�F�&t�Tq�Ps;+[�ղ:�yg��z���Vj�W�N�w��b��u�-��#�&:ؾ�k��Eδ�a㻊Ԇ���Z��5yf%M9���}�@�8�r[K�i��THn:%�fQ�S�
����\z�ٳF�9N��'fmM��5_3@@M���������ih�o���υ�=L���ʵ�A`��v%@�"`Jv4Su���<
q��s������gN���*���	��c�@�{�eG��-�os�����`K�*Xu2�X�ŗ��-�%mfCG3�������V����g'����3���|��+��	���2�� ���L�m�p݊U�(X9����J��$��D�����]֑���f|�7m/�S�Cs�;�s�j�]�Zӗ�\�ebPS]���&V���y�����������-o�Mx��K1��9��ҭ84?��f�퇹���5���&.M6��82�:p�h�i��כ�gun�(��֍s�!Îeq*m����f�A
�x�-���r*!P�)unN�AY��t��[��ioXa �以�:}���b�e�v��C4�����4����[�zU���q[�WЋ����hS��������d�����@&+0؝�bf	Y����&K �%{�2�d�{%;S��#�ǖpwe��qo���Z���C�6���0e����m�S"���`�q�ջ��V4k�s.��x�%��X]�f���Y��#�Vl� ]�uV�})ȏ�o�ܞ9A�_M7x�#��=XØ�t�"I�ğlGT��Ah.�F��Z�m��S:���8���̭0*��	UaUzO�I�̤�č�m�n�W�\��bP֭��M�f�Q�����.Pk᷑T�'�V��X��V���y�x�^i�c�j)��e�3L�ݬv�[�(��z��G>��>P��T����<�wZ_eԧƐ�;Z�ς���ћD��N����i�V�ڹk�6��ט�/{7:���<���e�J��V�ȹ@H��HV�/d9�_ݼrS	r<U);W+=7�z�i*Ό�{��}tt�r!W���rE�j��Q�LcKcԌ���*-I�2=�.��NPY���i�N����P��w٫V�0�t����9 �x��B�7��i��Q�*_6!���Ӫ<����W��n�r��ې����m�����3"e��ei�@��-+��	G3C��:�ͪsGd�.J�po�&���ة�iyљ^ԪK�66��ݑ	f�觋f�v�//�t�LK����Vm�L���m�9��c��� ����ښ���f��x��U�n������6�.ՖLF�e��gΎ$xO��M��q�P��[���w��cX�D
2�J�#�KJ�U)}˺���"�m����nl&I1�-`^��n[��rf��S����u���+��
Y���r�݈���R� ��+�e-�a}ult�@�\ەֲ&ZT�<;S/h��8����r�62n��Kn��U��M�<EZ�E'�(�i�lL��p�s�Wv�G� �jR��\o�Qn���+s-ttٳ	���+9Arf�,�j�OW�(��č������cYN�wӯ:*�ۃz��Vժ��4RN�^ɲ����4&�zl�vB�M.���`�u"6I<2�⮔ܰsH�8f�T⚈]��KM#\`yKDW-��.v͊6��驝�,l�YI�K�D#����Z9�����˻�6��}]�6�Zi����EK��W�u)���@o6�ujG����
p�HZ���X9ל�q�{p��0观�UG��<�;n V���Yfs͛�}v��1�s7�m8��)��3P���T�ow-����v1�d&U��L��A�8�:��X;�;�tlɔ����uZKp�[�	�g^4�}i����_6������3BU:���֌������S�Q�V6�Zm��m9�֏>�:�����F�f��F�ɽ���X%�|�O{�,�����>���Z�b�e)�(%^\�=�7DB��h޴�
{E[v�կے��c��|V�ٝ�v��z:b���̧���]���tٵ^-#>Z�S���[�It��scx�g��Z�jcw��ɾ�_�m
�Y����ݟwdn���|�вߓw�5&�f�Y)U�ߠ��o<�oI�\��A�A�O�7��lS^MV�,b�mZ壛X��%eIX��]�����Vж!�oa����B��k`��U���.��;Qx�cZDŒ���"�$�4YkN쿺�\%P/�kor�y���²O e�<��@�Ŋ*�Xఢ3WK�af�;��D����޼aq��u�1i����x�cZ3�b!��]}F���
�giv�ҤN���6����ٛ9C)�UL�c�j��!w:��A�C��Ǆ��\K:ŗ����ۧ3/"�e+9�W�M]��:*k��������vgs��b�&��R��;2�s��΋�������	y���Ö��=�S����z�5������˗��P�Ӟ�L7���k\)�e)=��^���:��D��9��l�mv3���#F}}v��G �(ąuڮ4q�4�v�!.���zvQ�&[k�S]�/�Io��k�pJ�a�RN}
(�F�5󿙲�����бg(��{^"M7^LG�����r�;���R-f��R�V��+�BZ�K��s2�"�|/���ꖕɖ@;ʹs�4iwpF�*�^�׬Z�%$���+:�\�b=��u\�}T�.��u�;��Jq�M��m�{��j�
���Yr�_a�3o"�����if����U]�q�7�*hYt⼷S)�<,	m��T۳���~4j�1^���ع{B�ydǨ�����0A���cl�rweջ|)^J��v�
.�f\�v͊ÔA�4Q�>v*+�M��g�"U��� ��6w�Em���Oq����ȴa4}�󘚪�t3�[���iV;5�ʗ���K}rU�j�lw��0F93iNb�w�N�G����U~z�8�Qфm��{��kd�锤]�Xr�Vi3��4�:�$��1��j��K[�N�$)u�R����c��"!��v����/T��r���K2m��U*�42�<jz���@��s����=�kn=\������)*�)ѾIpEMٔ-�ø6�Cgm��䦺$*�1��'3�"��3(��棭s\@�So6�/��v��R��bd/ۥ�I��!��#��us�1*�Kz4�֩F�x"��齙�Q����9[�����y��s�1�B'���Q �w(Rͪ=���^MNvLО7)[����{��#4sP[X���v�IZ�+zEx��I�50x(Q�o�4��9�1��!�KiCZ�Ӑ=��o��}�r�uNwJfVtX�N�̭ɩ��	N����Č���sN�Y�Eض�:9h@���6@Z��GV�ԛ�U�Z�υƒ�[Ʒ�u0Q��2b\�c[X�e���8��G���="�|.�[�R�}�!e3��X�4�&���Z9|�Y�Gښ�iG�o�ag�uZ���_�Z�@���b�l�e��6VV�u�e^�1��(�'v��oA��'���r�x]9"�w��o�=0��N��U��q��i�O�eN�m�r	<:��n��r��f�V{s�2��ِ�W��6� ��pN�b������jL�yH�GUc����	4��5jU�����)��;��]�+:Kou�ҷ��=9��< �/,�ͺRl���2c��g$SYZQ�(�o��g�	[�2�ܙ�H�p*�6h��o9�=�8J���E]>�Z�b�˺�6u[��}ή"{~�0ma�[��;@W�^j�6�iu���h�Ύ�Zgkw���	��T�t�qS�n�8�an�\�Z�n��U�Ć��eRz��g��1An�]ۮ��(�+F��һ�S��^�!r6�3E�է4Ƿ*�K�Cz� �+��M�j���j7:}|��J%���5gq�^Ү��G��a�ܺ�tXX�WP�UG8m(�\�<�N�N�)0#l����5a���E+
��G�7�c�@�*��c��P��ZGCUىF�����d����n����]���'��T}R���77uc	N��c��5=���d��eї�����	!I�$�^o<E�kLv��l�An�&ch�ya�hH�z0�v��6��]��W�k��6y�gn�e7Yre�q���\�ք�.��c^mtP��Bs�&#m�M��ŝ���[8�3��ųc>��+Jqv�g�c��G'�9��V}��9S�3��P8ܻj�y8n7wo2�3�x���瞰-�>�K���a-����k��{�#��rt�g�וcq��r���v���v�y�Vի�7#��=u��ѭ5��h6.۰k���ڞ�\Y��ۖS^MV^7$�6_�yy6�j�;�켓�ݜ��'����-=�����nHx�*��c3�0p���L'6��ŋ�X��_n�y��l�]=�w����IN٬��<���A��ڽk#en9���a��N�Is�VIs<n�Y����fV+f���ku�$#� d�=Cnh���/F;�ٸ}�1=�q�;.�v������cl<ޛ��sk��|=�N�(]��]Ǎ��
��f��ͮ��̧�R��`�6.2�<$��ݢ�$���z:��:uҀ�rc���'�K��m�q�s���O2X;���}v]��s���t�nrI�|�#��]B�ND��K�g��ᴜ<����+��<v��.��r�ɷe����[�h��9wb���kR���Š��E2�G#���Uo��wn/<m��\��!n��f7m�+��=+Z�u]�s���$˨�u�͗��솎�l�v�mX�G��!��[7���בgEgn۝��dl��b��\Վ!��Г��{�lD�l�Q�ۻ�&ㄮ�2���]lۡ����t!�Þ��#s�I��Nܕ\�
��q�g7@�����A���ܛ��X����E�3�IvM�����E���v�;v2����-nW�M �Ԝ��{v��;t��n���;z}��r�/��s�눴az;91�8���f^�3Ĵs��-k����;m�]�7��Xn�:����\��p�q���>��Lʳ��H�csݢwcs�#�ݻN"�G\s�v�:"�[:��9��=u�6�Ձ9�sdy����s�/��Pu�Gv-��:Sf�/iqۭl�l�l��X�iF�';�홳�� J�+t���snK:Y�t;�.�6�������t�;4���L\�W<�nr�&��Nb�y�����n8�s�a;X�zwj::��������W[+�f�-�t���Cv�k�m������T�qύ[��˓�u���c�[Dn�%��eS�=���0�{	�&$ܘg;)y@۶�g�N��}��0��L�L�vݮ�<s�W�@gvNܙ�ս���pܺxWlG���d��ld�q�ᥩ�,�]�-�f�<��ݛ�6*PMk�K�m�tez���<s����ݡ#�-v���M�l��>�\�-/=�k��x�9ݝm��n�ulr�i���d���\�ٺ����Nփ�=�z���w7k���x[�2\�rk��7]��A��8��>��1m��v9ۢ��\q�r�m��8S�r�F�+f��G˭���Gk;y����a֯+;=���m���}٠v�uc�Z�b�����)�bݣ�"��<�� ێ�s�ЏM9f79.ɮ'�p���m����:��ڌ��m�t��ݎͶm	���!&��F�A����!]�;h�-n{[� �ݟNJ��guʼ�G[w]�nw=n��"66�'Q�6�׍�۹���Ǎ��nM��vՓ��3�nM�c��nk��m����%�׌�Q]q-m�j�ϖ�Z���1��bSn�%��q��m$�+q����E�<V;nڭ�{����q�,��}�m��BU�r�g���xv�9^�-ʰ�r�c¸��P�x�	mM-˱^��Wc!����n�2�V��e��l����d��U�Fz�z���m�{	�dJ��ݨ�Wm��K�V�׮�ۮ��,ۮ�Z맬3�s�l��	�N��g���=��Y�wa:{[lU�u!���0��էl7V鬦y�{CƱ��Oa홮x+��/dlk�6��F��N� A;��Z;m[��5F�J�\v7n�p\�!Ψ�n�n�'h�:��cr+�ñl{;Mm�o���f�n��7h��P�f�]�Jp�ݛY6Nx���nB�'��ٵ%�M=�=cW`��]��N����[l�pQ�\�n�g�#&�1E��uI�d��.���h|�s��n�\���uQ�j�)!Q5�Q�e8�^�8�,ݎ�N���<FXV��Di�c�sGlX.��\��ۖ���g`�����;,d��y�<*l�0h�S�M��3��>�]�vov�5�{k��:�O)����nq�m.�8�W�x��c��n�$�Lh�v.n(������y.|����[r�۝���4s�
�v�;[s5DKC�`x+�b�,�Ɠ����q�ۭ��:��y��>�Nh2.�l7�a���Ge$�����i�|�ۡ�dtrd��<$�7�n�&���97:3E��m�O�<��b5r��V�����q]s�1vQ^;GWi��ޮ'�����w7I�=��0�x���xuF�jq�'��VxS�֕�''��\8���v9�<�.nlp�\�ɶn-�R��ۍf�@�
3NEknݸܽr��>�:�zv�VN��&���'gc�÷\������ iUU�^�M�ӺN�e7n�Idˍ��\x�'�v��qݏ�u������<�jW��E��;��\c�q2�.�:M0 ,��7�ͮ-���`�nK��<��zx�M���om�	װۅN�I��ky��^�������[���O�vz�C${zܧ,���Om�
=�Kƻ�Gu�ں��D��m���	k�F:��������r=�Җ�gm�z��6�rv�
G8讷�q�8�8S�s1��������p]j�xt�oO�g�G��ի�0�̻ �����o4q�p-se�;�،u�z9m������W714��m^b�n����6�/X^j��Zm��(�g=4�l�hQ^�!�޺�ӻv�ڧ�Ӯ�I�r ���bnNl�7bD�`;j�B��9��(�ݺ�xi.�c��V���v��v��[�t]<V���=Չ\y�����k��[��zCS�5�U�m��wk��v��|��t��z�k��$�@��ȡ�o`�����p�=�ؽ]q{vbɸ�����[ƁY:�mg���N��,^:��s���iՃF�z�wn.�d���`ݮ2is�n���l�����H�͹��v]ٻ�d4�]��n��` ȭp9ܲ�X;1ܮ�;,cյ�.1�m��ۛ���a�<�1��s�����MO[����P�J�<�ϲ��pa�>��y�;�f�]m��F�]� �S:��鱭F�mh�^W�
�����i�5��q`�DY�Zc8^9��m�K��6�f�Fک=kE��0��s���۷g�s���q�zۥ99������ţt����ŧ��lh4�;m�n/we�1�2�Gk��/����j㮯bck���f�5���n���u���uաȃ�����*��1�dlv�q��˃��)���;	�=qn��/=m�y�ر�u��m��N�4��Ԏ��;T���<Ul�b�v�]�+3l��Ŷ������+d��ik[��n�4�#k/��G�#w#�,��6e]�uLn��tv��g��V�D����8��;�aN�v.��z0v8ۮĶ��ǯN��ݸ��۷��Nn��n�H�K5�.jK�;��׷�Σq6.�, ����٫O��L�m&��h��>�	�3��m����sѸ�^�l���S۳�b���ܤ&'m��"�-ۧgB���qk�8wo���m9�����Dn����wl�[<����ݻ���b��o]�&����p��3Λ���Du�]�sq���{=����q�CD��m��{z:,�m/g$�3���<v�x_^��woT�3z���nٗ�쑘���kfƐld���FHn�L�sɽ ��lG�S�@v;l<�U���t���<�������a��m����e��#k�l׋<��l��mۀ�lڇ�ƵˬZ��۬g�L1v�۪���c��6�-Ŕ2]�r����^ݍ�%���ve�HV8�u'O�nu@�p��(�kn*����x65������,��8`ݮ|�=��x��mͺ���=k��;���*vt��򙹋qe���b��Q�goX�ձ/N��ˮ�MJ���{�3N�ٴ���z�#k�Ӹ���:_C�ya�\6nt4Nu��9B�����X�&q���v�n).�&��.�n|Cw=۰��u�b��>���kP���z�mq=��.���u��\���ۛc�G���g'%��Wl�W v�Ws{�h�,Snܺ�<�x�F�^�HCӶ��';��^1�5fά�<�n8���wn�ŶB��`'u�q�r�q��<��в�[Su۶:�tŝ�q=�[/N�:7��s�u�n��8�wo+��W��#�!b�ُ`7T�C��;�q��;�b�s��(%�፻\#{;n˭�nƹ���v�:��D:��7�����&�. ݓ=/M���t�(�����ny�j��}O���U3ʮ����/Aӻ@D��6,�6˲�צ��-V,���I�mm�ظ��n�u����r�v魻��Dq�u�'�G��m�7���^x�%�7Hh!�M+�����p�]�۔�ls�sŋ���k��nK/vuݎ��f�Fj��Qn���bw�Z3�p��:+<�G6�ض�]�U�ô�ks�hK�ݚ��A�k0���O��ओ�ݭix��4M�[s@�\�j�T�V�[\�.j��]·:*�"��(g]s��ӜTc�ՠ�Ţ3+]t��׮�5-�WZ�r'�bnZF�卻0GVN��R��rܹ�ҙ��̌�n���GxPx{zz��^��k����;���GV�0�PXը�KR�m2���h�%��3�q�Ų̵�� �Ŷ�\�#�(�K9��Z�p��ḻ�X��"8ʑ��Z�j��"��[�h��s%�R���\�1���Pq
���r�+B�,P[J���R��,V֩Q�E�\���Z�R�&
嘆�n��J*�X ����Vh��8�1�c�l���։fZ��q,TX���*�	iq�V0U��˙h�a�Qf�X�E�\m����ڌ�(�)QEEL�r���YiEP�,b�J�6�m���(̮f5*��S�Z�2
c-ˆ �R�2����T�AD����YET-̬k2�ԣ���9����L�V"��وPq��Z�R�Tm--q�X�+�VbTV��h��Q���
�*����T4ɌMR��!�̹[U%�QE--EY����EZe1��,Y*V(�H���k������
��3c�L)��u�a{k3M�5_
b�u�̻W�t��m�Q���ۮ�����ת�����n�u�-N��:/�b���W���u��ŷl�8^J��8(`�'�&�I�rյ���^۞�\�j���[���p�\�X8ѫf��̂2�r���u�;km��s����-���y�J��l�r�QՓtuF���n�h7.��{p.�������ΰ��\�t�{uqt���Ɲ�ݷ����]t8ۮ�A,�Vwj�; ��o9�A�|����e0��/i���[3���]ZϬ�_=^�q�":Jp1˞;0�v���r-��]�ٍ��qZ���6g����������d0sw��/c���7Ud]�6Mz�]p��M�e�n��k�<�C���y�nN���:>]nz��k1j�Y�;[<{�q\���<8�.�ڛƅ���b��^0u���p�;w\;a�qӽ�l�;zۓ7>���s��;�zیg@;����b��֐��m�����zwK�=PMvz@.�)n2g�l�Tj:��]�wm�n����(�����T�sġRO\Í�.����|]��^����C�s���<�Mv��1�����(�v���$��ΏI����v�
ۭ۷�՜]�'h�y�-��aP��ۮ%-�m�@�g�C'�6�v�4��nَ�b��@Q�ZC��ԯne �����F�umO<�[�8������\���vN6ۭ�u�{^p�W���6�5�2�Q��1�V\�7 (s\W��Uv�s��1dw���f:L�3�]���*�̽u��]���s��z7���s��9g����7mnD����碷a����s�;����:=����X�nڷ[�u�E�-mƫX�dӻ��l[���Ӽ�c�C�z��>��YNa��5��f�u"u��1��������P��Y�k�q��`շ{�����2�;.ò���=�"c@��*��n8�
f(��X�ᙆ`9V�#,�{ e�ySv��ܘ�6\v��|����ls�qD.
܍�32YQs2���3��*�WTƙ�˙w��vr�0��q��]�9^p�}�n��ɜ�v�<���*	��/m�a{��
�e��9�(�
#.a��֔������]�Q����6���('��܏Ϊ�)nNc=B��0�L
�'���[��%�o?r@�x,a.���/'J'⺣��L;��_{����s�����(����z�������I�i&m2e؏k��?
��D�ֵ�[˥�i
����~U���yhF�A$z��J���܉�Ϳ]Y?HU�P�I#=[�[#�
�v�����VH����R2QJ@��9]R� ��[���s̯H�[�H���`O�V{7�(7�K��'X��l^Қ����͠�>x��p�X���X��܋��q]f���tdJ|��!��iq�$(�]��{.� >gf��9��_�+�/����	���AVz
��Q8"q���5wC�~�B�7���=d�˜�] ~�y�te�T10}U{�t��H��a�OT[����F�9���Oo��q���W��H�� .�av�s}T �vvց�o��
�Iǽ=��[�V�$P3�ty�(	8��ł��U�/-�w,z���IUޔA'�~� �缒|�M�L�w�[�9�Fnu	/�O���{��?��wY���N���%䯉��&�P�cJ.{��7;hT�yx}�\t	=�+�I���,=����L�=o���o��jn	��'Du��r�nx\v�k�z,ۡ�[<X6G	C}��?�H�A)���=+�A ����3��ve/.��w;h����J@��۲R�i=D�$(�U��iU
{����M�p -�$ ����;� ޝ�b�������k���%a����u_ę�ޫ �~<���M͖r�l�395~���չ�z�f�::wP�o.�����V<{D�v���H��5d÷�����]��*����4����n�$��L�Y�`D�Ў�y����L ���䀬o�W�P���b�0��l�u�%��)�-4\m0e��u�!W�m��8.���G��
�>�_O�Wt���w�	�wH��.&ف2��2�rz��H����[uqЍ\4詒��.��M�c`�`1�' \컲	nnՒH%Wu}�t�#_e݂L�����I��F�H�9S�'½���W��l�7�H�����y�7�Z�c9�
�OQ$I
8�f����%u��r��aq���g��go��� �҉z�a��]����\�ܲ�������.��AY}H��z���i��.���n]�Yá��f/l�1-�	�j�in��љ�.#��W�4�Ղ=Û�l���wK���[T��<��<�q���%=�](J0 bhGE����N�ܗ�\7��>��5��֐�)�B� �{�}@�v 0�E�O���q�&z;1�,݅�霽�u��n�8�As�<i̛	8:<�u������eٔ{_�ygz�	��_J �H&߷�����3��e^]��݀I%m��V�	�ā(d���v~?q�C� �Fo�ՄW^�V��{�U
c�-�{�Y$}���O�)H R��6
��7�Y���f��m�=���Uf���� ߧuY)]4��H�Tq������E�T	�eh��ݨ��OleBֲ��/�Q���8#q���5C���4�=���
H *���� s=� W��CQ��=*'�UO24)]0,�[T(K����>�wR�L��(����PG����2(�^񘯴g%A�NTP���ݸ<,�Tj3A ĉkf���\����W�w�Y��ܧ!�m��ѥ��*��S�r���yw�А�)�,9)���k\y�;ץ[�-�u�c^ݼd��x�V�#��A������kv}#�]r�n�i�����-�(��w'g(�ۛ�gq��m\��y5������GZݹ�\�웑`Si[�G"��\ͱ���899k�� ����[��yx���:��tf.Wl��u�l��H2�6V:[+�����눢�&�|��D�͛�g�A5��]�"n�\=�r�4d+�R� ��W�$d�� [%F�]�7��=V���K��p���  ���+g�������O3wK%a�0��,H�I@�V݋����]��A��U�� ����'�k��>��_�m T�J�r�K�&���'�����&���B��<���q��?J����	[`ٔf` ��~�iP@P;����l�Sw�+��� 7�<��|(｛���){)�?�Ͼ�-iB�V�x��nwF�,�sm��j���=�z,H��0��=�����B��ǳϒ@�=��
���[AOK��[���}/+��'���݀Ho4'N"����ꂏ�e�~;��,���J�M;P�F$�U�:oE%7�Zͻh�j�&�fQ�\��ʽ�3	C(�m�1mY���^{�/fI+��k\��c���OĊ��ݟ�wJ �k��}\%]u�G�am�%�\m�eksz�� ��J�(W�G�$wM�ץ�
�y > ]҉NC���b@�2J�W{eg�E{���U�I��7����gG��m���H��%���i�
]�r��$�wguT3٫6a���*�Q�6���:�m
��%B�ʻYl��ee���2�J	m����?W�̃�0��ƞOm��6T�:���������	�����|ߣT�Q�vm  
gy sZ�]j��wï��_���U�(|6���p�R��z/���x=��ڀ��vւ	�߷�X)��Emg1�]W����Tq��`��,�0AǾ�Hvz���y��,�<�y�_��i#թ�S�wq9�~��{9�9-:}|�˫�ٺt�#��m��,<9е���cq������y;�\%Vt����O��ž���q�ɗm���g���㨐WvO��~���	�=��=�y����	\}"�	��I(=[W� ���T=\S��]��;kh +�'�* 	��]���1��B���Y�]�q�s���Ճ�]9f.J���8��%�n�ZwnلC���_ߣ��
�)_���(|H<�z��+'��B���D��k�$����m�F�΂D����P��e���]�@���$Q��A���O��w��J�#:b��逑���I�^�{��N��B�P�*e%&N��O����3�����B��!0�J1X�m�ul����CK����OӶrT�P;���s٣���
���
�&�_����t�l������r�T�!��i;��en^EN�{��w�@��>s[�כ[�[�7,|M��J�{U��hp�Z[�
L'l�v�޻$AU����{�uC�۱ (d�ھ�(�ހ��a{���H�Sq�?A��y�s�`��r�>���.ol��m������ߠ2r����� ��mYoUh�ԇ�*�*������Y����i�
]�r���E��k+�����M-�䪀�Q��m�׍I�.����~�ɗ����O?H J9��.��U{�|I��Ki��jQ��+��K��ݓ�%W�Q?xt�pH`�!j��glnRb�zc�@$7�V$��B�$~��rjyl�JU�~�$=�۰K}�8�L1
�IE��D�Fuvط|깼9U�y�`��:Q�����w~�2T��e�I�.�BB��KS2���VP[���r��CJ�<6�T�l�s�Q�4�P�L�Z
̶jՋ+��L���<<�&DXq�TN@�QF'
L<mwm�N8��nϓ��'86;�Mgy��0n*원�8Ӓ�n�0pI��ĸw��ƅ@�mÍλW=�������_;�mry�YL�k����W�O78�ϴ�W��9du���܎a���i]\�����v���7�����4�e�M>;v�V�q;i̻�.�9.ܐLpg�ѩ���@�^#�5�a�n���l��g�zu��c�˵!ps�-�ͼ=�����c�'H�~�������L���λ �~*�eI ���Y��^��'�0�UB�
�ҁ,k��&C@�@�u`�{���༴^d�˯uX$�Y�(���H����^���ްL��W���T�K�sn�I�^�X'��f���w��~+oe������i��	G"���ZS#�Ok����Q ��ޫ�	^�u�>�0UW�P:=4�0�Z���{��~&t��G۸|=�n%LV� Sk�K������+d�b��Z�Q�cMI��R�urL��pY4�x�a:-=\����-gm��8�L?��IŽ�G���U�H%OO%T2�heǔ��~Q:��Р�׻v	˃��&�̻��b��h��|�h'ʷ%���Tg��b޻�L�C��)q�u{w�}GQɼ�{�i��c���F*˱*e�A/�l��- �r��M�P������ ��ܩ g���_�]����Qe�~c^��� ��nd
ޝ��U�~�b���kq���;UP����f���ʀ��
U���=r���+s��Ww��IS�'w��j�r㜴�
��#_v��O�]���r��tiP@P9=�A�P*má��/�m�$���X���0�[~�������n�+
=�;v�m��;^�S	���-=��ۑ
bDq6����@Y�E^�r��T� �Oj�> ��яM�֋�Z N�˲�����g�A���(��w:WĀr��x�Z.xy=��A+�� �AS�>�8I�]�R��:e{&`$s�s	0�D̻�ɽvOĕ;ҨP�5Ӷj:��uj�ŮÞ��� � j��m�l�]��kx�����ԃ':�j�!�o;�o	��،hIx�wWU�K�;����v��As���,�]gf�z]���:עV��1^�u�~���)/7lz��w�Y�YZ�x��ZWHZ��{XoA�N�ѷ����R����4�">D5Ko��=�+W:�μ��).�9�qKOL�;eCjx^��]�n���e�i��ctx��������[��tZ&y����H����^ދ���;���PVU<�9Y��H�:(ʴ�]�.�;|�#u3��COe�C����))�w7yRz[`}����C�Ӌ���pI�.����C���pQ⍝�9nK��®u�:v�������]�2J�{t=��GF����8��+J�Jz1m�PP���+���2�}�v)[-9���d�2��Z����T�ʄV����	Bi�r����\���l^c�{�{s�9gN�l�u�(�m�_�,
�fݥ��ug�<7E]�k{�37kE���ѽoE�0WwW�>�Uݙ���5U�;r&�Zi��)	��ۆ�Hy��T���j�����;�J���-+��7S4ð��p��ꬌ ��]�䆙as�,�]z�[h�F{8�N�0��P��mu\W�gjy\87씊ܡ[S�5�z{ko�G�|�)k��ѳ/V:sҩ;�!S���z��k�s�ˁ���Uy¯w��X�@I�ܺ�Y�L���̺1������&�BΪ�pC��,�@PMP��W�����e�4�AnkZV���Q�Y����k
�[��U+Ke��i���E�1��9��Z��\L`
�F)�db�Z��Eaij�,KiP��aDZ�i�Ŷ��ն,��FҨ��2�+��*i����E�MD���Z�Y*�+m�h�RUq.R4����ZZ+D--l��Z*�����U��8cF֔R�m�eE)h9��Vc,ʥcR�+ZDiKm�kQ�-���Ȗ�ڥkVWXh�J$SVԨ��)jҌPbȳ-���A�AR�(��X����C��Gp��<������n1D�b����a��QH�Y+0���J��L2��*�b�EQKF��2b��b5+Z�hU��Q2ɖŘU��F,�UX��ie���m*#�*"����L�F�jT3
,1�TI����l�؈���|���߼�	*{�C�a�ĐI��}U�MK��j����;j�$�T�Т��y,���s�)ce��9y��Ӡ~~i@AR,d�>��Wu�}{��{N�(�<�� tͪ����F�,\9L ౟;�#����[��q��,@���l�5�Mv�f5�7G|����~�N�%"��{.�!Ol�A$�Wu�lv�,k�����_e�$��z
4�+6R�ܾB��r��~�<VH��P���(A���H>
m����%��zv[�A���(��w:WĀIίu"M��j�=����H*gJE�w]�J�~k�I��j4e�mu�`������R��	&����vo\h����n�}㷃�qHK�Ff-毠�>:Fz��[YbJ��U�^4knJ��yԯ���ˊm7[<zV�����gi �wҀ$0��|YI�H�Um�$.��<�0��>&��Hίm� �~ڢ�Lei�ƫ��,0͒v�q�oD㴝��n��f�<u�Wgv5Y�f�1u��Pg�P\���N������.��S���W�Q�ޔA����R�e��QH�_ge�v��a�F���@UB{�j����y* %(����)�?X��rDPpH�j��ݿ��[��d���5�y̬Ѡ�N���� ���H�d>�S�p�f�-g��ѴI����(o�{~N����t7WY���	����~\o�k	��q�e�sk��$�ҏIe۩�d^��V���;lX$��Y�w�1������K���⧪�-nj�@t�r��&�fؤ#�C�aHF�q��5[��է�H=ì>�;!^]k�	�1�_�)�HqD���q=�sA��Żw]�t�z�h��;ø1��g��k[��;n�in8�O!�v��۲ĺњ�l��:3��mv�@�DB���s�{��D"v�t��sۈඍ���ˮ1�P���E�so<c��Rv����D�u�]	�<�X�}Y�ܯ/+��=fqƄ���c<�i�M�i"���ca��%v����s'5��:����t��wOlg�ŝ{`�Y��g������L�$��#�w+�Y �~ݯ���_�!u}�R�u�cN!��_D*��g�P�PK��M���ޮۙ��4�L����IW��	<�DrsM��s��V	�)`����%���v]� ���$����J�/9��h'�]��� �SΔ	�ç�Y
A�"-����ذ�s:�`4+ϣ�B���mm >���ӓ2�ؤ�;ޙ�.�j��_�ă)��Q	(s�	9��.y h7����wB~�_9��Vlίa~=�����(D̐2҉�Y���rh����(u�=�=����܋u�����Oׅ��8�����`�J}�D���ʳf�׶��ļiTʰH!=��~-��!�$.�Һ��,b*��g���Z����4�������V��`N����֡:��<7��D�n�%甗ˣ:���X�y�2n�A)�Fä�d���A?��
$���dX���i���Ρ��uEe)�9:�|I?���dA��b�T�<���^������ �}䅌TCz���EW}�n�u����8�wH��[�d�����&J��8��P�vBqᯰt�S8p8�f�Ow��d�W��&WE�i��,�@{���d �D
�����ì�++%B�����@�>G���W��%پ��x���iuX�N�8�l{y��D���g��նI<1��U��-��3âA���(�����~�T�@q�$�T��?y�}��u����w�~�Ԃ����g>�^>�Þ��y�H/߿k��xH)�{Ͻ�:�^��sZ��l�㑓/�0�#���a� VX�Y��~}ޞ�����O����
�Rg���y��aR
K]��u'P�������:���k��|޷�8d �g1�ɐْ�v! Y�'���:��Z�������9�B�B�0���Z����7��^�=<D���V������i��l�;u��㗫�m�>��jð��E�Ao7���V�����ʫï�k+��"4!|@����{���td����|��C�+{��8�u�\m֍na�¿����[��_����k=�#�H��n����JʁbT
k�y��v%`Q�� 
.�~��r~�W	�5^��|��������ף�3}3�ff��f����;߽���؁YY*As~k�1O�����?s�u���ĕ���{�!�aXPaRT�}��H,�Y(����ۓ�1��kX{�����fh-g���{9907��p�=�����9���������߁a�!��-������y��z���]�߶s���![�E����� ��)��G�{���\�x����%H(�{��u%a�i�V��2j��6Ì+����1%�7|�s��.}��7���:βQ��@���è�iu��|�>!�]�U������߾�{�
�_=��r��nk5�]rS�&��>�ԂΌ����������IR����ּ��o�|��C�>V�IS]��vu'D*AH.o�}���{���!L�b�B?	��e����׍���
CV�����9�H[)
�i���9N T��?}�~�0�z��ȡBqO�.��i��0E�:�W�ܦl����e�Eߣ�ú�8������������9�`\�d!X�(3�ug�]��:+]��w߽�����o߶u�+o��e=��.6�F�0�¿��7��
��Rs߶v3����^~�u�ּܺ�ؕ���vq�X�
�>��KH6�����W~���$�o�&��::˺N)
6]w�N:�����7u�;mc^9un��3g�������e�Z�O� �����ޡ��H,��Ϲ��C�*%ag��܇RϽr��_>���!�N'���:��
�R����N%@�|���?	�3U�xu ��~~�a�=`V�=�������s���߽�ϥ!iHV�+s���@S� �����p�:2VX�Pٽ��O��w�}��|$�7��?j��MWN���º��oa��IP�(�a������N�� �}��5��]����Ă�����?op8ZA��+���=`V�<zy�[�1����`#�:�P����u�۝����*A{翷��%B�*	+
w�{�!��T�3���ԝ�������x�x2�X���>���%@ #7����Nf;�,�~n�P�+RZy��vs���<�S]�f�ח���o|�9N T�ʝ��}�u�d���P��~���:�D���?�r7�7��+�K!g�z��D�Nx���a{�r��fA�ήޗ�(��-k1
�c�xV*��6*X`���R�Pc�����zw�-��b"v8^���<n����m���W7lTv9��I�	�����:;�˲"{w:x��m�pj��5�n�;��|��^7.��=�5��׸�2q��7�ۃ��];�y�x��{�:ƻs�4K����u��q�B�����k���n_t:��׳��yl����z�w8�B��Qѻ#��<��q.:���|����qu��	94q#���3·=���]�@�����m��rZͫCQr6���7cn��n
�	�r�S���(��U�n�g�8��a_u����0ĔB�~��nd�eH(?~��@�J���k��}��q��{���z�wp8j�iH[a����ïa�b�>��\�䯀d����������������v�'_3>�gFM!RT,IXS�y�܇XtaR
J����l�N�Y(�ɫ�=�}��ν�گ��D �9����q͌ "���y�ïXjB�����9�Bү���D{����¶�s_�DW�j�@��J VT���}�u�d����b���u ��ޏ6���5]:�6Ñ�u�o͇5�~��m'
��V�{��:�c*�Y�>��@�J��Xk�g���������_ν�X~�<�p�A|5����ܹ�sZֱu�N�ַ��:���d����3�n!�N���������"�$�,�}��C�:°�
���=��I�
�R�g}ܜM l��}�_y�"{s���b��G#�c��[�m�n��)YAu����ovd0�7	pD�q�{�d'���𕆾�?l:=H)-=��vs����
��]��18�S��8~ӭk^ߞ~�b{�;��ԂβT,C<�϶uĕ��=_�Q�Z���Ӝ�Xta_�޾�pbJ!Rk��/��������K�����YH`/E�yO�
�X�"x!��pwٚ ��ml�{M&�*0?n�T������I�KL�0��s��>R
y���bVk��g��5H)��?_?:>��~���u������F�.�rW��ĝ��?l�t@��d���\�}���B��T��}���y��g��Ͽ�߰����T�L��=�ԝ�����������z{ܶ��3Fj����ϼ�^gwS���m �2�3�}�gi
�i���9�(�Ybw�����oͯ�ny�?2��
!����:�RV֏v���rj�u�m ��=���$�%�V�V����?}�����Wx?w�@�@+�����`XԂ�3�ہ�R
Aa�����Y���������ƴ� ��k�۠���K.�a�gX�7t�ܽO`�[v��k8ŋ��p-6�rDL��@��#�@��%ed������&��*IXY�y�܇R�s��y����:�����ݝI�+%Y(������]�?LĹ�4f:�@�J�_s�l;�"˯�,3�i���/V�i�_ �_"��\׿r'*Ae�߹�ۇY�J�2T.����t<�ݞ!ԕ������yu�\���:ã
����4��T������gY(ʐP;�����y�n�7W��U�(���3oQ�%��o�p��oa��\�2��9ܖ���M�V�\5�q������>�$�X5�3�w�T�iK�s��ïFi��G�WYq�F:�k�19w߻�Χ�k㏟����3l�����=�gM!H���s���°�*J�k��ԝ��{��y��&FVK\�>���M _�s-��Lњ�cèJ��y���`PjB�����8_(/��ߍ��ea�N?(�"yY�'
������w��%H(�ߺ��0���e��ۥh�u��U��� �y���#�Z(� [s8�m]\���e7!d�x�2�@�����:�7�a���Q
��X~��}���%R
<��{è�8滯?z}���?5���w�� ���9ﻇ^�+C������s5�U� u��g���J�k������|���g���ɤ*J�IXS����C� ��y���gR'FVL9��;���}���o����A|��d'���G����U���jA@�_{��$��H/��^a_ߖ��~�H)����}��ĂΌ�
����vu��)�����7Z��4�!�W���l5<Ǿ�����ND*J!Xs_s����d�*�Y�u�#�O�aG�FgO��=��Ͳ�U?�*� ��y�>O��G.s7��d����7������[�K��2��)z���.�O���[��bfW6���N\y������B�þ~��p�r;�(�M#1� ���_�Y<��d�������
��y����纾k���x��q ���yϹ��°�*}����N�VJ2�VW\�_nN& vQW�4g�H�`�HI.	LW��bnݽ=��v\���@Y�h��������c4f���~@�+�w�v�����{��9�B�HT��s���9-
���:���� uxr���2�������?}�8�D����ݾ:�4̚3W\��pa]~޾�
��T������ɇ��<�^��q����@�?}�:��+�`V���p8H4
|�ݑ19����+z�t�E �9�~p�sY����D����Τtd����>׻8ɈPIR5����o=�k�u�f��y�:0�(¤�3߽�gRu
�Y++�{��'1���M\.�v! Y�%W���~�4����~�^z��jB�����9�B��+C\�rNA�@��w}���}���}�������=��}'̣%B�����Ρؒ��?/�/�ִ�m�9�q�c
��5��� ��y���L��]��ݟ�
���6q ���y����AH,;�~�p��Y'>�l�J?�1��.J�\GQb��.��[iT\�@�:�d����K�B�U��U��:��ݽ5n�:{�]��tAg��O78��B��%jL*�Z z��sohp%=��߳�%�����Ӧa���蹉Ai����]�3a�]/C[wX���[K+٬Nc��ܩc�+��*�T�s4��yv�OU�;-{���c��m��݇��J�F`ȴ�
�v{���m��mьa������ab\��0�)�#����唖1���ƴ}oR &T��M��ĸ��t���rKهVЮ�8��P��Q+k/0k�b�q��v��1uV��^7
��US�
�/Z��YO/i����!���]���Ak������UR9�Ǩ�OUA]N�(i�G_ �J��6�P�b��n`�m��(Y��2�;�U��n�����QY���yb�o]N⻜�yҡ��	�@z{d�VU���B<��oN�Gxrͼg��FMlS=��땍C����C�d���j�nQ�@|*v�*-�!��a�ʠ�v��W,د҉ͺ�c�k��V��E����V{�lk��bB�n����֞-���V_U�S^�J��*X��t7�j�=�c�w�Tkr�.1ˢ[k��qCF�o���J܏p�P�Wy;l�Q�6e2pRw��z��a*7��5
oil��%?u��&X{u�9��Q�:d=�!Iem�W����][Z1��݂s�3^�W�:㕞*1��;���l���ق
�t��g`�*�;�K�߻�Ǧ��*�h"(���R�)��Kl�lKmZU|f+�Z5*�F�+��[mU��0�*�D���
�E�T��k[t�j�hե�m�T�lZ���D���-QU�ܹ1�)�̵q-�ң[T˃��1Rť�3�Ū���V���
�be.%D���Z���K���J��p0J�j��mlX�[E-�K��V��T�A�fXd�)TW.*����WZ4
��h�s(�bZY��"���m
*�EiE-+s�E��Z�iul�[[U��*�uK1�,��Q*�"�eeb��FکU*�s
�X�[�Ƹ0��&%*�D�ҊK1�LVL�QV��9f&-�b�+m��%����ꬨ���K�-R�Qm��kkd�b)��ڕ�kq3"�F��]2V(��Ѷ���JՅimeK�\��sT��H��Kh���Em�FTEKmWVѪ�e��(�QT+(ԣ-�3.QV�0-�`��j��h�Z�rխA[D�#�I]i�PQ�rʮR�T��+q�r��C)��6�h��q��V�/uu�����Y�&�n]��V|n�qv�-��1G��m�kv�v�q�C��eR�X܎����֏g8����cm��ݛ݂8.�C���[�O��v�e10 �;��#����m��v�zH�n�ձϮ��g�`�YwFh�s���=!�/m�n������N��ӌ��'8�س�]����d�ljx�W ��@]W$�ˀ����=s�i�]�y�M�z��p�cc\�-۱^sV�N�΁��b�%��8gv�qW<qۺ)�j��qם�y�vi��Y�,��AV��+��qk��(�s�.c�X�n۲�	l{lY��8C��ʦ:���j�<mX�5,���ny�fy�\%�������ڽ0	��y�K�t�1oB��2��5���.K��� :�Q�O^;v w;����ލ��\3�C��-=�"���Ln�.���[p�Y.3������{q�S�)������.�8��7a�i���gl�sJ�[�X�b#�.V��pgs�i˹�Ϸ	�x����+u�TG��㇞'�� S���d{;k�Ħr�-S�dyl�V,s�mn�l��x7Z����K\��y���ɷ!��� �.��*'@"��73�9�9�9��`D��M�la�Gr��j�vN�t��ׂ�U�v��݈�]�Ӽ��]3��f�=6�<Q���{a]֎N�+klۺʂ$+m=����vϲ�=���:#���ۗ۱f�����޵�uԭkn�#m3!ˏ;�v��랠K��J��׉^��Cs�����yS�N=�j�Kx[69^sm�g��i������8���{t\݇�n���:ׁ\s�n���ǎضG���8��E��ۧ<;��}ԵIu&�v���h�ٰm���p䮶�wGkl��̝����[wcBh��gd77�{i�,��U\ۻd��LX�p����7\�D�ݹu�uكv��v].��v.t���Lt�ǰS9��)���fdծ��\���.�����r��>~s��]����ѝ��;C6.�s\=�(�gs<�ȪBF8��ݣ��<#�*�7Ny�ڻ=����Wf/^��k�<:��m�y��ak�7��2�����rW��^�cx�<��\]���Op�9kuf�6���k��v7[v��V\��Sn�n��w[sAwl���c�����\~�ui��#g�gv3v������svlq�: �<�k�l���#q���;���9��u�pD;{���*2��'��G�#�߷7gS�����W^g}�C�J�V�}�u�A�a����=>?g��a������l�N�Y++%eu�w���B ]Õ��"ٱ��#����0#�H�>�#W�ғ��z ���ЈT���������S�eN���:��J��P�\���YoG���y��8��J��7�5Li�isW\��q�u���Ða��B��B����}��:�`ʁR�?��_Ͼ�������T���u�w��ă�H[a�}�ۇ^�
�����f9���y�Z��O��������q����|�Yc%{�y��2i
$�Q%aOy��a� ���}��:�z�߼~�^k�I�) ����4�B�����Q�f�����8%a���v�X�h����������q�~�]�����Eǝ_���+(���>�:��J��P =���a#��{�ͩV��|��8uh�ΎP7,����<�v�\�'��+�����F"Oهȿ�)$��~�¾y���bAI�
��}��:βVT�P�>��@�V�ߏ~��7\�?{�o�� ��>��wT�il?s�~�:p�*��<�*2�'%�"�g~ɴ�1UD|G����:_�?G�້}����XC$W������7��U�I��[��J�٠��u�N�e��k�UF�%R����Z_�{��=�O9v��LB�*%a��}��q�XVaRQ3���ԝ��ed�o��_��3��.~��D����S�C� [60�,>�����z�R��߽���BҐ��
�����ߝ￠T���+(����:βVQ��P�>�ݝC�J��{�j�k�j\��!�#
�_���9�zc�߽���i'�*K�>�Ͼ��u���*��}��tJ��R�{�����|����w��HZXy����u��o�~�-r�f�W2�.���8��������׻82b�+��4������M��$�/{�y�aRT��}�Τ�!Y(ʐ]{�~���d����&�B����p%u��q�s6���O]t������x�1�p��9=�0���>E�K��� �#����X5!Ih�����*Al߽�ہR
~���k��xw�,�;��wp�:�YY*{�����+�x��}�֍���:ã
��u���%���w��y�<a���:Τ
��}��tJ�R�{���H)ʎ�K�n}A�����t>� ��2���\ֹ�;�>�����������p*IRI��y��}�����S�aM�DggI��q���~]�"�m�{8(o$�����R�Ty�c�GV�!R�����U�.�I�xY�WNQbB�=�V+燇��S>�xmx|aXQ�IA3���ԝB�X��A�߽�ԜN }��7:&k5G1���÷?u�����s�_,��$|*�?}�{���-�+X���� ���{�ۇX�>���럾���z���D�y�9�82	tw��9nfe͐�L�����)��y�ݜH~�~�=���������^��Ԃ���k�{��p� Ґ�;�~�p��w�=�q�>�C�>wm���C�<`!��F�(	�omsK�62u��1�D��d������E�m���׿����2VVJ�������
$�)����!Ԃ��]�����������O9�l�N�Y++%eu�}��:7�yr��E�Y�H�V���a׬
5!�{�w���G@�}���ii
�i�{��q8�R�VX����ngY+,d�{|������Ӟ��og�u%afs��}��h�n�C�;W���m ������ۇ:2�Q*�oI��� v	Xk�u�>��)
�����ÏFuw��R��䯀d�����c�W���N�i ������Ă�XY�{�܇Xv0�)T�L����?f��.�a��T���G<-\6�S�<=6�sq�o����g3�d�>�����VXާ��wVJ�
�e�8��ΖվG5�u�8�7d}/��� >����׽c+���w'"b�����5�����R�����`v5!K@����8�ɿ�����C����"�ʮ��DY ��?}�}�:βVQ��g|��A��?�M�����	�Zq��r$�4���M���t��R��Z�x��󬹎����w��SZ�Y]dֵ��a�a\�ﷰ�
��*J!Xw���Ό�%P*T�{�� #�8g����~�{��,�Z���- �B�?w��ß��0i��Z�fe�'bL��wgS��d�ϻ���-;��&�?~��C�*AaC����C�:°�*J&w�~�ԝB�VVG���{����O>�ܞĨ]���\�\�h��8i ��7�v��!m;�l�JB��sž���ٻ��uͿ� H�4��|Fo}�p�:2VPd�X�w�~��:$�3~����u�F[��70�a_�w��{�K�Է��s5u������1'�T��=�߶tgY(ʁR�g{�� v%`V�^s��:{�?s�R�y����ף�k7��)�.:3W5�@��������v VVJ��]yϷ��d�_���~��߻��Ͼ'�v$�/7�?ra�0�,aRT����:��VJ2�X����U��2��l��=��i\�oڦ����N4R%�p�/|��o/z�D��Uࡩu�?����O����}s�:x�ݙk�e�u��{�ox�'��onVwI�C���i��|�I�鹼�s��ˌ�gY훝�봺��_7\t<r���ݮx��\^�Kv��c�g@���˷u��'�4�Ok��Ta��ړ�ܰ�\Ȧ���{g�����Ksx�EŁq��kX;��k^N���W�p�ݴ��=�v�㲆{��GgPu��4�Wo/fx9�;s�o*�2s�]��7f���tO\&ќ��5n��ۀ,���ݭ����벃ڰtW^�Ma��\�L�j�c�~@�J��}�Ǭ
Ԃ����s�����(}6�]�"� "7�H���Bve<�Y�'��nH,�d���{��u%|1�;�Wt��H�Cª��l	^BT*Mw����w=���Ă��%@��}��R����}���Rgo��?r�[�p�Ai�|�0hᆵ��˸OD��>�ΧP++%H.������D�
���z�:�o�g���y�8�XtT�L�{������eu�>���J�n�~��b��h�5�4�ȕ���>�{}u���� �s����vR�B�`W_���N*e�������p����>5��'���Ȁ+3�P�>�2��#щ�$َ�Ԃ��������RPB���~�g`β~���y����<�u�Ty��l�R�+X��s^n2�m!XO�����c�y�޷�C�E�����eY��7v�<�&�<y�Q8��ק��ݬk�,k\uۙ���h��{�Љp`q9?|#�#�_��'P*AH.������J�X_�w���aX~���k���<I����͝I�B�Q� ����p*=��o�.��r��R���}�ïXj}K���솗����tO׎h��O7������ܛa,��iL��}n�<�\\�yӬw/8�V-e�u�8���1R�u�^�����H��;�~��␶��`V�����
�
�@������ngc%e*�����_�����z�_��u9o�
*��~~������$�%�;�|�gY�JʁD��g<�ٟ�y������*AH.���
�R�s�>�lß��0P,1�5�`#���(a��{��g��?FJ�_y湳�&!D� ��{�}�:ñ�H(�=�gg^�ޥ�c'FT���ۓ���n�w�9�9��0�ᤂ�>���~�,jB����϶s����׏ޟ�~v���_o��S�(�YS�w�w�������7�P�>�6�V������~|�Hzv۪��c`��+�JuE;,vۃv6�j8�h�2)	�D7qk=�����|,�?�G߻�l81%B���߻��:3��e@�P.w�~�Ԃ��v���}�~�������כ�R
A�a���ïc����U�:3W5��������l�u��Vk�~��<��u���Z�gLH(X���}߽�:ã
°�*o~��|	~������o`�;����>H��x\�u�˗�P:�����v�XjB�wϾ����>�~�{����x�u=�(j���w��꒞�I�iW�𗂎������Z�����V�+e�.fS�������G�Zө_V<����=�7����*eO}�����v2T��@�{�CG����-�#!E	�_pa\������1�������H)?!Xs~~�gFu���PJ�fwϽ���Xk���n�|�ܿ���~��������wp�AzaϾ�0h�:�Z���@���l�x�d��������ɴ5�ߞ��t��蒰���:ã
*w�~�ĝB�����1u���� ���x/s�o��?JKk��shیDۅ�&܀f�:f����[m���ogs�ډ(#O�wti��@�_� �&�������Z���3����t�-�+X��y� i8�Q��w���5�u�������ì�%ed�X�w�~�Ԃó�m����չ��ff����+���l8�i*#�w�}��>��=a�߿sp�A@�T
g}��H,� �s�$��|���ɵ��[c�5�ʯ�}�z�`V�9��W.���u�� bpI���vu:�YY*Au|��82m
$�X���绹n߿kˮw�}�=a�
°�*g|�ݝI�+%ed�+��>ܜM�X}���:&]i2����a��݇��s�4�����8�XF�,���wg:R��
���wIȁQ? ��������������n���>�r��C\\tů[W�Xgy�����[t)ф���˱��􇮉E}�,��o?��ί}���l=��w9t:w�$���'�FJ�C{���:�Xt���~���5�ӭf���0�]~��$�%B����>�ѝd�5Oݦ���)�@�*7�~�èJ��X���7I ���=��ïF_�rF�:�߸��i��ሴ`p8���d�͘��B�V�^�y�&�m�j^�g��������sWWWY���3�>�ΧP*Aed����g#&ТJ�IXS����C�;V	��\�^s�y
��7���gRtB�VVJ2������6�K��yu�`�ц��q+o�}����Z�)�E�Dd��8��/}��K������B��i���I��@���~����u���%C����n�}��;��힤oOq�Y��hsY���8��¿�>�Ã��%�=���ѝd�*J�����Ny�������~@���F�W~}���R����nz
�g:��ˢ�Mf���w���C����{��u���$|	���p?M�D�
������y�aP3�{��$�k߷�6����&�VJ2���w'"m�>-��5�9�%�vq�X}�~�p��R�3�}��$�q���˞R����r��(�Xw��p�;+,d�T3�{�Ρ�IO����B�݌�8��M�.��U�Q�����P��T�[�#���gm1�+�����C�]$I�3I�p�{�ظ����E�|���{�Sn��ꀰJ����rd�6JW%�niv��ln4Y��W\�$���=���:��1i��v��Y��	-cl[�k+gE=s� �v��I���Nw9n��O5:׍Y���U۬�5�%��m��͔颬8pE�v˝�Ss��3m��h6Y-��N�xq=����r��ܠ����G�r�m�Sgg�v���9�;�0�*�;svd�Kt�a5�űk�uY�e���/JF�Ӷ��u�k���Y�������6[S�w������o������B�����p�'c*�Y��߸u �/����ۯs��_1����o��ɺA���o���z0+��}�ū���uu����I�����AH,�w���;�;�>;����l�2m
$�T������C�:0�+
����߶u'b��VO>1�{�y����g_/�wryh]q���f#�n�5xm ��y�w0?5!m;�l�iB���k���������
Agk��|0��� ��߬_�P�?�b'Q��������/V��oJ$�e]�?���I%Ž��E�(�?v]z�]Y<���hG"�w׷d��P��p�]:Y�)��ݡd���O�ŽA�[��t-&�����C J9��vk�A��H�p����7l=Q���Ͽ��߼Om��%p9�� �U����Aq�*r�����|�{��'⯷����E�D\)đH'����;�JQ�{�u.~�[��䛂ޛxq_�Vz�U-�H�l��r��/��eT�
��!\1�ݫ��W�o��,�Uݗ2��g��<#��� ���}Â��|�x1ַ�|��	���d��ǚ!ȉ����mu݂A&E�A�A��ח��ѼS��A*��v	'�"ޠ.��FLP'ӗ_;�W�'�"uVU�A���$���y��l k��ﺅ�C�R�F�j4�bڠ�'�vguU�*�u�Y��I�=�`�dY�(�N�8_n!~)��-V01�&Dl��b �i&�I��[Wc0m�>ۘe�h�$.2�%����:�*�hG"]�H2/m�'wP�|R���G<+P��� 3{l.�&�R�d!�����o�$L~˝o��Bmή�A�g�|H$d��	�TQ��{.�/�S3<H��{苅 ؒ)$� rw��gգ��u��n=�4�̼�,݂��ׇ/��GL�f Ϊ��n�?f%O\��[mP/�d	�$7w���#d���Kk�_!���s�u�+|	�J:�f�z��Í����=qp*p��o���Q��O���_)�O��ޟUg�,�"E�c4j|�vi�ft��i�sy��H�{�Z�FX�o2;e�=`"s��u|]@�ok�3��h�V���>�ɋ3gU�8�k��.��ū׶V�ݨ�f��9ylͣ��aCS[�}�K��h�jl,�us2���D�;���m�IUm�0�Ȑő�Y�<�=@�띌ϕ�X�	W��w6�V.�����a>Y����l�f��mm�C����:'l��嶣����5t�+k2��<ʻ���`���Km����+�k���:7��y҂�V�B&� �{���qۻ�1i���w(��^eus�W�C��)���A��wN]�WQ�:b|�v���<�E�*^��]:i�zxiG\.U]y*�;�X.��8�����z�E�4t��nj&2𥳐J�;��Ro�i����y�"�/�7]��o��%�o��V	Zf�붝�39v���s�K�i�U�&;L��{��T��+�EjD\�{�v�Y��2�C:[�h�DPvY\��.=��g�׷꿃�2��T}���M�q\	:G{2�������@�m����e`:��擼��Bu���U����o*b�!ow��r���m�����V .�W[�إ,��U��~��5ާ�W���*մ����X�bX��Ld�)KVQB��i�̹�-�\(ҵ��-�8�4�D��*����Dt�1Dt�T5SU�bV�V6�6ږ(���̤\�q����[V,1���r*�ETH�ibڥ���J�R�kt�J�pF�Y�b�
,DL�E�iɖ\��̸":�Q�*(���k���JZUJ�-�[h�X�ih�-�cB�mU�h(ܦ*"+��(�KY�-+��ܣh*&V�"��2PQ�F�U*T��ك�[J6�ZX��J�J��!Q`��EaR��URM7
���f���c
ڔYJZ�5
*#Ae��QVKj��ґb-��m����Kj2�A(�Z�*�P�TQR�h��1m���(��کi*�U�X�,X�U��QPb��fXƖ�V
�aj6���Q�F%��j���Z-�#T`�ֱ�f,kc�QU�"��e��5� %�ޱ��_R����h<͐�d@�2]���m$׫�˾�|H5�� h�9  ����ۯ����
�m\8�mJ�\��,�AW���^��	{�?��ǁ ��uY+����N��W�u�_�mIq��1@Z(��Ǟv'�+��4X�Ev���Ê�=��������*��{ΩH;;�`Y �����c����}�pɠ㷴�&�j��ʲO�*�iE$����ł��q�$ߵOL�WƷz��{���=mw��u1�|�o�U���!Ev{�l �W����B��s�1*v�N�T�&{�R㹽v	zk0��E�"�A��ܮ/=�(о�j�c��TP���~Ǹ#۞��C�8�ƅ�AV%�fjʘ�n杺-��x2�\���ܶY;Orc`A���yܮ���'Nts�h2�˾w|7����������y�L����!����
o� �MNzj�1�qb��du�z�W���~55�#$4�n�e�M(b ����)!m��z�y�W^[��ݞzl�ˬ�=i9����߇�p�n��侱d@+s�W� EM�G>��O���׷�>�g�U�{P5�ߍQ������Ωݺ�b�~�U��M�g�
�ݻ�H2k���uQft�Q��`�*�<!��c*)%ή��&O?i���|Z�[�{K�����r_ As_PG�{�����iGvwݛ��T�����Iޝt,�\ɦ�97���o��ٱ�N�ݒ*l�m��,E�
�����Y��gq�:�p�U�@c��Is��@��M������7]�ظ�gb���\{h������d��=����hFU�&�{�/����+�������}.�F��tY7VwL}���o��|M�k�
�XSY���2����ֺ�R��9�bL�n����Rztx�X!N��4v�r��;[[������܅��[pݶ�,�z|��Д�����5��ph�O1tdސz�v���9'���{]���ؒ���4vs��Ӻ���#i��ٶ'�us\���U��9=�ɷ;���u�U�d���62�˶NӞ�nqv ���*�m�����͠�۫�$���(����ۣj{k���֝���F��\����wFBDqI����݂I�{C�I$��vs��7��}��C���tu?|�n �)E��@�į��Uu7~w�\H$��ƈ97�Ř.\p�����}Bc�	�	�W`�th���۰A�;Y�^��ҝT�s�$�5��Y7���L�h�2č�d�.���upn���X	���� ��7��$�����ߡݝS�����h"/uC_4 �
��w�5�?w[P���Bήf�����>�fp���y=�| *w�O�pgy�i�>���1�P��l����������%�n꽰���8[g�����i�H�iE'�>�A3�`Y �J�o]�=N���~+1� A���;c!	!M���Q��H ����]�g�Y�]o&p��<�^M�yQq��Ն+Ū�۰�w^`�����܈�J�G!�q̭x���5ktYS�!���׿���x�����~���HW��vI�V<����r�'�&�0��P.N�J��{U �e
�����>wϫ�$+���'(L|�jFR��d]+��r؇�Dy�B<ݭ
T�$������]���^�Oה,�Dp�2č�d�.�{v	'���S�GCu�
׾j�|
��T(��ڹ ź�S��u�rشX�:đ��������c�����Ѕ�B�b1�ty�M|Ј�c�=ۛb�$��uY$�{ʾ&�Z	��o����f��_��X��i�h���X�P���^{L��w|=}�C�y�VH$�	�����²/]h$6<;�!	 m�ӻ�mu݂~�m1� g�V��|$���pE;Q�v�{1vC���=~Y��2��a�Q�/���7.�ں|4�pY}&���A�b�)vf�������c��� >+�y_ď� ���2N+Ѕf�1J2N��I�냫������A!�ڨ�/;���^*�@O�nu��hE��4��������2	/{�F�v���'�,�%� P�.�o��Cu���@J������~G�kl����糗�<z��Ξ���ʨt���	���,	�h������r���y}w� �\^�d���GC�ٳ(�;���A �����Z�Y�;�so��K���w4���)�ՂA��T$��{�X$l�������	��06�QI@��iK��]�Oǥ�5ƪ�{'^�H�9���wU��c=,�-�v}'Q�ī"� ��iOĽ�m�%W����;����
̿�QQ�����q�=s��wPZ�+�����R��9$����S���בm�Y�&�Q���_c��| �����50�(�0��P2mu�$���V�]���T�8����*P��T���K�K�5W<������}�m�V��mٖ�Ąٺt���rn�{� mTR�A2�w����S��qW㴺��
�?y  �]�D��2!O#Tr�u��T�of��c<L06$Q��E�[J���Z=kp�X����!�_��0'6y�;�j=z���boj)븗Ǣ��"hE1ܵ�����	͞��D5�3�(�}|����t"=}��  ������W�&b�!E� ¸a�X-��n�#+�^}� 
s��D?�&�憻v1ů�_K���I}PxS��QF�&n������M�:�{�N��c|���k�fDg�|NwSh @"h�n�Dz�S�-{xm`�QH�m^�~�鶝�p,�{����sF��a{��wv:�^W�����/�w�Ä~��?�&�~���F��=u�-O�|> ������pœs�ny{j���x�k�����;g�ՅAڟn�n���ǜ5��;��=w]I�ַl/���t�m��n�գ��pKgqnnŷD`.8b�Fb�9�I���sΚ3�g��/��b��wYk�7�d�d01�	��W��ΚXt��l;�ݯ\�ι�Y�Ϯ2�pq��ų�t!p�k;��q��ފy@��x��[�#�61^���7l�U�{9�7
@])�w���cMR��=�R���p$�O;j� 5;�X����j��k��� I���
�A�������$�[g6��.�F���s]�Nvۆ Ѽ��@����72���A�X��bGUk3r]��K�^륀��ͩ0�O��)���h�F��&�E�ަl�Z�C.0�;���ہH�M�^�F��K��7;�Z���mZ�l[��Uftɇ Vd�C��6Q�Q!S���t �/��a5}q�"whα��> �2+ ����d����cIg��=`������<�<+�hֹ5u��c=n˷\ه�����������Ŕ�m�"L�'1��Ff�N�>��o)�}�Ml9��e�K��jHټ�������l��٘Y�T�ex�;dr��^�:���|��Q�[� a[]���8�Z�������r�6uq�Ҟ]#��SM>gj�7����Sp�v�duH��f÷� ��{'��~h�_:�[ ��vf >
�=5>J���=;��_
�V.4܉��n��]^�H���y�@�j��잹9\�����4���&�3 Ib�g��Ċ1#���~�2^�E g��,�ݘ� Ѿ��<H祪c'n.ਐ�ժ�K��po��P���w�q/�_%;�}qp}7<�� ��, �}��g�|N����M��K�wۇ�L�)E98�q���!(m����x{��cvy%�77;]�ȔY7��}	M��F�����2o䳞�� >w�n"7����Uz_om�D�Xv7D�_��0�����h�$D��	��d��!<+uy�N8�V��g$�@|_of`w�M� ؛��U,um����g��u�FHXj$��m"��f` O{j�� �f_]���y;v��=s��"���K�<��t֘������$n]ع����I�l_���y4n�Hgz��X�3}#n���O�� �O['�[]߮�"K�t�n�
�!���4��ݥ���hub�p#�p���� ���0 �loyL�V"��Og�m�&��c��fE��ܹ^I$�I��XU�g�y3<I����`H���*�E�f���"Z�ZNVD���2�j6#RԸ��ohg��;9�&`��W85ɞ����s���>��%��	Bc��=��gI'��V�	j���/����rj*�䪝�m�@/���%3l:d��M#R�ruO)g{�z���}��'��p� b����n'��ױ=�}W�@].W+d	�3�*&������Ӱ 7v���Cٕ����=��@�D��6��|�jh"�R�)���}���8y�u�>��[A|��t��+��m�uF���Y.64����M�W��m�#�1r;;*�X�=,��m`��~!Ƚ4����YIdž'[�Φo���]�-��@��Z�Y���¸E��F2�M1#�	a�ꄓ�ߺ��U�$����+��Ri.���h1}�Y]��݇�W��W��	��%	 `��q�lc\��7<f�y����^�$	�8A"��n�Y�a�3�F��{�M�1~֝�@���2!6�0�Wc���\���6"b���a�z�7��,(L�,-�v�bIr���nnC��W� 
K�:i �e�va8�xs������\�v{lTh��QE;a1�����n0 �����Ƴ�ޒu$5�p�I�����A�Z�����CE=�H�S�,���؈���]p���� |N���V[�&��_^� �%U��[�V^^d!(R˛]~�($��(���_�ǧ;���Z�D4�{�3�D�U��^%=��+z.��ÙR�������A�.��*QٶQm���Щq�	)^<EZ��`�ݧ��/L5��FY1)��,g]W6���MCr�tw�����۹9�r[UrV��4�oφ]c�؉Z��l}�BqV8�!י� gU�t�G\�����ܘ
O5,@j[��g,��m"ћ�~Y�=D��ű�2�[�E-ׅ�T�,�ʇLT=f]e`�LX���V���]m��]W�$D*ġj�ʷJ�a���N�bg_]�û3��d�7(��]g�F�)ř��[�^�*p��L�U�c,�0�98�@g0�xwhC��f]�G3_�2��sF�^Wi�捼��d���),؛�\Ff�n�����D[X	M����C^,�̆P����}
�(g]h�)�6qD3�GÝ��qu�8�w��4�`s+�^�qI{cr�j�k07���a��tm�ܡ�2cy�-�k[u���y3,^�)/=L�Nm<E3�aW�
i��������w�5w��g���N��/_2��);��w�]����*6=�ϪdI�Ž��!|��8,~�� ��ݼ1oj箌p���+م�q�:a5MX��T�y��׶0&���M�ܲ�d�N��f��wU%`j�]Tr�ų�|�t|u�B���kHW_�9�/9�u�]�uƭm�[+#��5Q�}�mp������e�J�&PY��{}^��{��N�r%VGݓZ�na�������z�b�%)X�R�����[@�-�h�K[*�Qd�VѪ��VE�D-��-�h�V�lEc�Q�J����*V��E�R�����H���әj-Umme�kQ%��Fڪ�A*1�Ub��(6�mKeb,DR����V""�KXŌڙt�A���V����QB�)F��9�X�e,j�GIV�ҖՈ(��QF��m��Z,V���-��%�P�єD�*(ղ�[cD�Qmj���U��[�UVۗ1�h��j�F+kh��5��eʱLUR�Jڴ�X����T[�b8�[�-
�T����R�Y��U�T�j��Z��TiD*X��U�V��-uL�,�Դ��el*�YS-Je1��J�Z������S��F���+*V�����+�8-kZ�*ZY[ZQ[R��1���In6�<̎�-ҚM:+��v*M���by<� �k�v󌝺9��.ņ�ku�f��M�tO[x��s�q�#���Ӯ�K[�y7EW�ʽz��\���	�t��o��kqʽ�0��Pz�,�k�����9���直��[v{�TL���@r/�l&�0ї�2���y�t����)�����Ζ����ͮ��O'jWEm)]m�;Ogc{m��8�#2�9B��Z;Q�ݠ�����v칂ֳF����;^�p��3ڌV�Q�e�=(�]�y�m`5�ë/v9��筛v{p��mݜŸ�Qr�򘲠ȸ���k8�m\��\��7nd猌�t`gj0��dd!^�[��ۮi��z8��<��<����҇e�x��=�1�g��� )XN���#4�\O4ܦjKܝ�Zxqa��]�K�����v֞�y[��m���@e`i�n!�=��c��]F�!�u���;<u�2�ms��S���mse�n���mtn���ҝ�7pr!ۣI�Ãiɮ�eގ�mۻ{&n瀥6�kV���݁�t��ud�dѸ6d���v$�R�+76���s���۶�:��ヮD����=���m�f��yy�۶y���.{�[�����Җ���e�8`O/V�|�q��lv��ۮ]��ɗk6��N,��'g�O9�7ˏ�5���vw	ڡ5�زu��s���|�Y/E�nP��%Hۇ����]en7�se��[�g#nx���F�msp�kX�'�q�n
\�z��xܗGv����v������+O=�N^���;��Z�M�n��z�����ѝF�v5�ۮ�t�\ݓxc�7:oC�z�:�0�TD�t�4�yl�{N�t�ڻp\���psF��R�Y�q�sa�{Nޭ�l��Ύ��N^9��>5��m����z�nz7<�U�c���=�<�0Wn�7�p�B\�Ǡ�ל��zS��� �^���@���>:C�չ������S��W�Z �j�7Yw	�՞�P�J�P湌VɌ������s�#��m*s"^�n�s�˭8��v�Q�x��C�{[�����GJ������3�{��*�����8�t� 5���z�\r2Z�pWs�ٷn��Nԭ)ű*ׄ���:�?ϖ����b5��8�g<c�@wf�"��f��g ;E�;�K�m�5�{;{\�E�.\�v��g�h�_'�ϝ�q�C��9xfm��y�7c�iaPh9�N½\�������sGh�nȯ=���?xr�?�e��b7�ᬯ� �w<X�N����?NҊ�������!���٘�^O
�DI�F�gy��I#ƾ��C�>3�SR>_����	�O7$8�ۇ��=״^�ϩ _���D��	���_z��&���~�V@��P\�1���n:$�;}�� �'}<܂�֮��d�B*(�o�}�ȼ���π�7oy���w��0&/z��Lɓ�]~�ջ�$��٘J�Da
F�b%js_7!�1}���_��o����9�˲6���g��	&���%���F��_|���;}B�gy��6��m:�l1b�k���<�y�nT�9Ӷ���߿zJƭ�v�}�W�� :{m��1{�M /�.���+с�RH�tI�MQ��bU�&څ��n���]���A�N������]���Ua���̭RJ�W2X֯A6�&o\��M�c�ȱ�vf�P�F]v�)l�Ai7.��b͍�뗢3�|�������{uWvz��1"b���C@&�ɲ;��iˮ��K4d��b7ts�]xDJI��*���.�p�mN��h��`/�A3[����c"@�r��gn]�\Ew+���n'�>A�c�@ 
K��`|�����2��;~�ٜ�w����(���)��&2��`Y���[P`���}m7d��֭|H���a$&ovf���uVB{�/��4�n���kY%[;��H�h�����W���q��.9K�=���H�LD��'z�"P	L_kv �{�"i��>�H�����Y��X�n��!fB��*�[��$�dr��.�q��6V	&���Q �߻�"0/n��)�]q�s�~Ϩ�Rb�TIQ2J��h2��@ ��� WV�^[��K���m���2��Ӎh���Q�8O۶��E}��2�TW�^��^�{���^r$e�{׾�6�~�S�����>�|>�[��'��k�U�D�?W�vf|�V�#%�#f�Ǳ��w�3�Uf�.7�����0 :>s�2{6�j3��ؤ�G���^y��D�� �����8�"t}n��I55�+&5�~��:h{��|�N��� ]��EasZ3ԃ�eĄČ�H�L����s&^�ڻ��}�ݗ:��v�?�Ͽ{� f@�����eo;�o���| ���5G��*�c���0d[4��{�ۢM�+l��UI$�
�ɯO2���&�����I�n�;> �{ّ'ry�$ ��Z��������F��!rd!(R�ʮ���O��_��~���kݧ���5���0 �ܞ�+T�r0D�i�#u��Z���v��3�o̢q ��� @)ܭc��3�_�)��[&Q���-zk�J�n��˭�S1�sH�m�4Oz!��i������9�����	����#���ٿ-��|�O����~��)���1+6��@��UR�����N2����ߢ�O�t��%Ě$��|���ޗ�X��VS�W>�"�(�ơ-����dV1�[n�v8㎝pB��V�s�������}��A&NU���I$�U��A#{o������?t�ni�m�$�M�N��>��VP� �QN�N��{}�{��W6S�y��@}>��4��K:�$�n�{�N?�yݿ$�F����U$��*����r  �7[��˜�Bڎo�� '�<ڒ��N�u؉+����Y���QK������N+jw�b9��� �7>��I&�<����ۥf�=d��Urb������S-�3[N���7��H���w�߃$�I5D�I�3�����E�6�Ul������o}�U,�L�tw�k7c.Ift�Z�D�{���&N�/����0epSL�1���zm0�URD�k6{s�ӄ��M��u���v��t�3�c���{�S��iƑlm�A۝n;E�0�W���]��d����v.E��r面8�v�!\�v���bB�\�X�\k�mpn#��v����]1��nσ�a-���h�Q���î��݋��ed�9wU��ْ���l����.8��/'=�b����	�i�gx[qǛfa�9��;;aJ��������סQ7L��.��l�B�ZI��]��,�oh�e��D��/u� ���1 �y��fR=��qЗ��λ�-3QO	qb	*Z��nb��:S�y�8�x��v�� ����h���0ȹ.�}�W-3��{���EQB���N�:�<��,��c�8���'z=�D���$�ݪԓ�(�����؍Cv���/��ω$�_*X~$�I���� �'}�k���?o���	���Q��o�u���!@��jJ��H�����s�E��=���=����u�fb "w�Vî>(����7b���y��B��Oi�5�D���ۏb��n8�;��	$�~����`���,F��[k��!�s�y��@|��[��F�7F��*���Ud ���d�n� �t�e�H��S �<�B�[J�v�e�FH0lD�F2�߾�~���o���g��MuXT�����ҕ4ˋ���ъ��* P��^������$��9��9> ;����`��Sa n1���柨�g�YP�b	*Z����d�D����� O-�Mzs���z���{_vf �H��S`}[�Y@"���QN���t>�EW9d�����w����@|���4�����~��Ĝ�����s� �Фh�#U����m �m\�=���~�{��G��s3 $N�����/�]�n`#=^�� �D�Y�&A18�E�j�S������^��U��3ۛ�$�C���ϼE�6PR(��U_{3����հ @+����E/{��}1��쿷{{3{�M��8�(�D�$Ī�l/K��D�	���M�~�6� N���C@#a�� �SK �/.�O���~ ��In��Y��d�H%^]B�	+��n����xؤ^E������;����Y��#4���7<�}��u�P"`���^�b�jڞ�Չ�K-��.a�G|����gٶ+;�����$�EO{�� '���> ���CT�VF�B�K���r�k�ŗ~��86�j�@$�Qh"���f�n�ԕ^���M�Y�Y@"��P��q�z�@ �gsİ��w����זhh��f4���̀�G�Y����I	�Kb#������v�up�[�ɢ[�{s�hc����=����N}�fLT��D�u8��Ϳ�b������u���U�b���U���#Y�4��x(��8Ap(��RWvYĩN��NB����_�@|��z� �s�m� �X�J.�d�b�$��u0&b�S*�m2舰��k�A�����~�  ���	�%���tNb8�\&G$��g{%���,�:Z��O��"7N�����v{s0�{��a�vʯ[�譈��C7j.�����"��-nf����^M�W_h�gf���kzn^�,�"�eXsz�Q>�mZ�b0�|�s?�H�Ji�j6�f!A%��o���bHwߪ�t�{�q+��e{�//��"-�o7����l2�.r��;�wG��ݼ؝��hz��c�3Ҽ�q�c7;Dc��RM�p�
@�Q����P��A,�w^D���t�H,S'�ďx봤���g�3>@%5�Oڈ�$�j)�J��$�2����}7{O5s =����|��u6��g�������4n�J��S��U�Wݙ� DOzv�R �5����m���� ��ݙ� ;��!��"�tI&�h6"wa-�A��u����k���g<X"=��0 <θ��ycD@؈]{��l��ѐ
�f^fV]���"G۷3e��AN��o��D��$�.K�  �G�B�f$+֟_.A:S�D�uW��o۶��hr�s�Y��N�xU�x�ƻ��+�H�s}ۓ��.���J�EP���}�{��{����ܒ[j�]��v�x��l��c���c��άw`�G:�x���On��\���Q�t��ƭҽCv�J�R���rFӸ�{7A�Ѻـ�bݭ��Wns��RЛK���nݺ�Y��8�C�c���V%�gr+�����f��a^N�������i�S.��%��<ciݍJ/l�ϵ�l��q��X�rh��x^�Ǜf.J,�̵�+���۷��^;9�dܜq�:,qr�i�6\�~���qtu�=*���3�w3 ���� c���>�*�}�m��C��Ͳ@&�/�UY����A�Q������M�B��7;n8 'ޭc@|��",4�8{�J�K�����L�)	MH��D��7$@�Y���Aޜ��9�:��� �'�;mI F3��󠪘�&�D�(�ʮ}�ji��o�0k�/.}mH  �=e� Y������ĩtdƾI*�~����3��lƃc�O#��h�;�rS1�G�r����N�s�ۿ���3{ݙ����{v�!�uu���1���Զ�.4��-ݽ�g�m���թ�|f�����{ﳄ�ܐ�U�-�yv��$��m
d��w��tM��}ۍ��6'%���w䬃�K��[TK��]�T b	.��.d�/�N֌�>�=�[��3�T�=;ӫ�S��p$���-ƍ��T}(f]zi�ë��6�;��B2��F=�u�I%�����#� ?9�e�~����"�W�]D�;+�o\�� �<Օ��TӶ��a��� |�S^�������o����ڠ�I!����Uz4Π���܊�kg�����Ϻ���D��r| {��oD���x���жz߰؈�mw�G/�����Ap(����1 �I�N�RY&�݉\u�lF���,�����ϒ_��}H����u?�<8Y�������Zx��cnK\&f�:�M�T��.N�bU���] 1R)�D� �]�r �9:d�&�?_<� X�����~�~]T�I!��na5H.�p��7~��8��*��*	���v��� ���3 �ܞnH�/�ѝ������9�q���AIp��z�bA#�=o� _�ڣ��J�����
�w[��y�F�c��5�|Of��� ��R�;�M��������xo�&Ƙ����[#0mv��xN��
 �Y�=Z�ƥ��y�RL˼��I�S�C�u���x]��섬�Hl��^��'UȚ�X�Xe��G�Xw�wz���0ra�ouW���jӮ�����f��p��z�:i]}�K����6�b��`��=*��\�]ټq�-`��X������(Nկ�sҤe\���ݫ��:>�дk�̋Z ��r��*4��g�gm.#ݠw9�v�	y�W���-j���N��Jm�9�G�������]��P�I�2�����R���an�S�x?dw��N����Lvgu�R�K��s9��[��[�/�%q�=����)%��a��4�vP�ݽͲ�R���^�jL�g���v�L���h!���ջ˻@Lս��{�2�'P�f�ĥ����)�h1�//zv�ܾ�r�v�gM����A`��z���U�.�gg�����g�A���(�;N��ԫn���gX�{u%-��,�@O�7�4���V�r��\�o�V���6��/1�a�z�1�k�C�>暇����D���*9F��dJ:�j�m�������F(8�`uɳ2i�ЗB$ӕ�񢽙n��+޽�����ّ.��=����u��ȯ��oOea�'�|͕��.����o��r��u4.cxU;ͽ�c��z�1L�R�'��Ŷ��c��,�Ӂ�Nѽ��)��A�p��D�[B�P�(��VT�F4[
��x���a�qUA[lXѢ�TZ
�*Q1+l��[kE*�eT��0+X�.�0*Ѭ���*"��DLq̨ʱA̸�+*�+�nU
����TīmQB�`�V�E�E9J�"���+b*#R��q��&�Y�j�EUF4���
,�\��*�����A�����TAD�c[J���kTUb�����i�\�Z�E2�-�ږ�h"����PAE+(-�cGL�WN1������4n\Qb�TEF	�J�]\G*3V�jԢ�-%��2�QTE�J-EE�卅���	kV"�+*%h��
*��TbT��AT�������FJ�U�rՙV�X-h���[UQQ�"�5j,V"�K�`�V0D���3�%��TZ��r �´Q-�`�"8�12 �V,j�QEQD�Q\J6��D�(�_�	5�{������ٽ�� N��o�
�5e
�U3
����VBv����+� ��  ����� <ε����^�uU:���/���f��:�z�*�nE�s_6��f��*��~�����{t��31A�=���$ |y�w��:�{����|W���!�9P@�����sr����a�$�hN�t��9��~~���-�7�n�������!� y�E�R�-}Q�.5�=��0��$����/�I�GD?T�*�m2迀ER�^���u͸�w'lh 3�ԑ��u�\����	] �0�1�$)�Z�������s�˦���Ā�H'���6>����0� b
�M"�ݸ��
�,m�Q� �>�� ��Yh�[����D�0�C�_p�>ӲϦN��������n�*�)��D��%��)��xՕH�B���O��J-xVJ{t3%FK��K��� >?~���=�� TR����v�
��܈�7�a�;�<�7�̈{�U�M�@�fݩ ���ݘH�^�5�����A'#q��i��%���sۋ�.l!�8݃1f��ݺ���)s�Ͽ�r��b��QQ�N�Y���r o����'tٖ���܏�<��@��u�e�LP� FK��K���H�ޞ��!�{�;d`�z� ��ݙ�h���gE��wm�9._��d��d@fI2���s.��@s��=��C�r������5��R@{;�0$�L.	p�ے�坏,���J��d f�� �=٘�A$���%���N�'�d�_z�6\ b	.��^�A"^�꿚�{�h��r���� {���`�<ȕ�O$[�=��ׂ��Crǉ}�]z*��F_���������R�D��^�fv3s4�5®��)��b�ڡ�jjݻ�W2������>Q#i����@;����ٺFǰb]-�s��v�����=m=�;u�9��@A��u���݋�7/P]��xw��Oh��I��q��[l;z.v����i:ݲ;��k�u���[�(����㧲�lsւ�k�L�*$�C��I�N0p60�{D�s��.���ͻY�q��q�i7c��<�6�0om�;v��nQ��l��u�n#���`������(�$6��u�+=�q�:��p3,<�\�B)q	=_�S˨S%%��� �r���Ζ��ǭ�ȱV����[��w�$�QoZ@a-�	����"�++gG��^�o�Oē|�� �%Wy�������5��Kk�&	Q�A�#%�[.�3@ �ͫ@�v^�z٨ ;_�3>I�{�,��&b<Jm�lD��_�8��P]n���	��y��u� �E����;��VF��fg�3 ���)
�����%�Fne6 ;��ΗN��g+�:�� k}���O�i�� �{<ܝ������?������e��!W3Vs�:�3�	\���c���ѡN�wNx���O~���칺�랺�+�/�w1`D�u[�"�^�Y�W��o2xRMm{���1 �'ٵo��Z��EJf�Uv�o��r P��Ɏ~ֻ�Z<S#j���7�Ȇê@��N�ge�]��ɫ�`�;2��v���Q����Ϫ�>��.���{��ﲯ���������p�^��Ԑs�F���ͭ�X�{����'[	Aiș�'7��a$�_=�l�8}����{������fհ�#o_R''�&	Q�A�#%:��x���"ɥ�w�o���V��>?/y�X.�z�y�4Ho�j����cƊ��lE.�JV���������^�{�^4��N-Z��@?9|�Y (��d�}�Ok{�b���D�BBK �c��Lݺ��hU�״�St��n
�`�<K�h�ϸ��1�ے���ܮI|�Ks_]��@Q{ͺ'϶�����t�[��lĨ�J3_]���� b	.XU���X	~��j�^�����U��@gN����vdF ���S��ܣ2�� �mP�"����UN�v����y� u:�*�9�����ki�j�}郶x���{[ԟ�+�a7ꃲ���6Kq��}�闦��V,�E��Vi6��v��L߽�m0'��i�65 �:y� ����3�'=pN̠�R���a��i�א���$�Eİ�H�/y�D�Oc� ���8f��ď#X���͒Tq}�w�[.�3�I!Vm[V�ɽ���=�����sn�$����:� �"`�w{Y��['=px��s��xZ��1���n�97�&͹��[x��c����hB�J��R뻉$O%ܟ̚$�Od�h^Z�"4;��K��={D k{٘�X\�DT�L�UA.�;ٔ��|���^�OW��oI��� ���`k�N"�6T����Z^*�Ϣ_��0HX��$u~�=X^� �fUL�f"{~�ܖ�M=S̀��٨��k�����K�	{VuWq�%M��B@^���� '��p� ����ʽ��j�:��}&�x[=�%!�l2�ќ��k3uS�,��P�̱rť�\e�&cxb�b�U�(�d��Gs.���һ���3�$�~�ۘN:�I�a(#MQ0�&��6��ö�P�N�M4��fb��}�� ��:��9�����#P�q2�A�`�1f�"K,�n���=����mq��Ui���7I8������y؈�R���&��1` O{j�� ����9�G�S�����=�������S`\�dGD2*��TSh.�m��*��,��Żُo���N�j� /��* @�]��<c�g��]U�X8#��A5U$������> =ۺD<�=��Y�vz��r O{����/��^�(���JU*���ONe(��2,+��D��[=��$�D�����'ӳ�������tY�Z�W�i����ALR��Ut��ӡF���an:��րUז�!��gm�D�}���CE��FVs�����{����w�G�7��o2)B��XhT퐫8�>ႛ�س�VR�fb�ZOٷ���|�x��{�k����� _�SZR9m5I!$%ġ�&�6�.ܫ۵�r;��c��I��q�u�ջ; tps۪�o�[Q�t� �F�kst�Xi�v�^<	�g�r�oqڛ��������� 8ۍr�Ƣ�'��8���}�����������]�}C�7j؇����'ewQ�Z��gl�ڻd+�q�l<���l]�8!/7��E�Nv�I8Q$y�;�q�ڱ��f���_X�&T�[���N9Ƞv�:�g���D5غ�:�RN�D⩳j{�����G�tt�QR?�&���#�s�z�ݙ�2���]���|��t���o[T ��P把/���.�u[٘�ZzAQ�]�Vc̫`|\�\� ���3_%@�f�I�0�
��'IQ�!m�)��5�� ���O~�����>��BI&�]|�
�?M��`6PG��	�r$�gfK������m�2��lM�qR�D�~����7��}~rDR�ɍ������>�#�*���J�{��d�V�Jߒ�=a�W�e�."�OY� 6������m�������{��U� Ò�lF`E�seM=v��FqbXr��k�1u��V\����߿��nE�9��.�{v�D�o��bA"I���@
�kb�vסY{�I��vf$�����bj ӆ5e��^	$����%�	m2��X�mHf�oy5�r-��I��b�Q��F�}Q�l����ĸ5"n�魚�ḵڙ+�VS�ಲ20s��L{��_�)�/�߷��o�I$�O؀
��H{$IC���U��^���d��>��ESd��f, >�m[��z"s&�e�x�/�ّ���Si ��D���R�%:��|�-��E��x� �~x��k�W���O_T�C��ҏm���`D��m�Y@�S̩&�%�o��� �w���;�.-\{%�\��+��O=��@m{���7ϭ�1��a[��}M���H܁(�X�Ϸ[����'g��dݐ�@�D���HyQ�����$�.�d��n`Ē'g�Q7�D���c	>�ޚ�V�s2# 6���	{mQ R�TU*t�^�X�f�s�'��a�U��� u{�� ��O2!��y�-�u�5 ���1D�)%UL��ޫ�D���	���o;��!3q#-=����c��i��bvd	���ݧK�e�����432ԵB�"�~��Ӡ��^�M�������.�
(��	��'U�������<,�.���(�3@D�d�ȢMQ&���v����G�Af���	%zH�����Q��[r k�kq��LP�h�}��<��Fo��R@�Ͻ��\fe[��<h�i1 ���$��%�v�Nl2V9n�� 3tl�թ]v}�tw����~ۆ���&n���M��O7 Dy���L����W-k��� ��+i|f�n�*B�,A%�o�ۖp|�.��fWc1rܷ���  ����<���| v�[�u�����_V�u�@��J�4�y��k�s� zo��su;�G���3�:ڒ"��va9��QO\07i��RoK��V�lߢ,/��� @}�}ٙ� |l�K�XG]�>��}Fxdʅ��I�򻮁��xCj׮k��&�#.��R��7�N�^p�w�❛Ar�x�T�g~��{���U�G{��jC������0��&K���ك+�{e�媏x��M�oU��k��c�vf�Gd�j'�f�����	�uj��:����@����&��u���Dv���P����61����Gq(ȅ&c��L�wm|���� �[^�p�TB�M��vF�gג@�y�����pGz(D�SA2��t�Dw{���zEJxOT�r ���vf|�^�l A�9\{0Y�����ӎ�%HS%�$�wݞ���A�i ~�j^o�w��Uy�� ��ۙ�"��u6�m@8"�K��[z�����e_�{e�<N��ns�" :��� 3}<�r��=�&�i�$�{{3O�R�!�8����[*��� ���s�����ko�W�Ϸ������a #4�9��trQ{V�u������W<!��h��%�tb�]a"Z�v�63�Oh��<��0��I檳��v����٪E^�Ρx5�Д���
R�,��}�O��!K��Џ8ͅ�;x�ատVee�����ݫ��N9j����;ONPK90��E;���V�[������� ƆVm8%�x��~Ic��Ҫbj������,!N!�����'	;�J�+z�=8�9�8E��;Mc�"����Dh�v����-�Ǐ)���\�V%��v�vHړ_4n�m>���Z��g���yu�3E�*-���D�h�.�	��-�ʒ��)Sr����q�������/b�oE�0ҫ)�¶H����sz�J�u��"�aIi
���T��z�t�j�m���c�ż���6��׳�z����qLy��/��[o_�d�u�!X[����ɱ]�Ӱp^mWV������p�E�Zޠ��(���%G�=I�^O��l�������`�N��E���I��q��\{,퇙C��"�C��}睊y��v�{y��g�ä�>�víq�*5G%�,wm{,l�T���EA�ʽS�]���Yo�wnҥ����:c�2~V%٦o(R��3i7�7
�!)��~c�y�֜�!���Z	��zf�Ld�pU��]�Q��Ti�Q�$1�51U�Z�GZ��5q�:����+n�G�W���켩.�2�b��ķ~ͽK�f�]���>�7�T;��h�:�db�
d�U�MhQ]ą�7�ޖ¿����`�$�}j�����+,X��k,T���PU(Ņ-��lL���j�"��W-�������Ш�*$R,��3�����ҵ������؍�+"����PDm���Z�fe)F�*�c+R��b&�UQ�J�A�A����G�AmRŴm�UV*��T�Ѷ�V��lP��*��1(�[e�b*�Q�Р�lEQ"�#�dFADkUt�-+�`�r��VX�UVڶ���J�E�%m�XȂ*��1\���[(��D�UX�iA��(�Z�l�������TD�TBШ�-�8��i"��e�(���T��TXԬX㉅�D�T�l(*J�U-�kb ��*.fd�t�*�jQX&5�-u�Ђ��-u����A`��X��QDU�U���F��b�5��`�����jdEAW#���,�mX���ʠ��-̙m��m��L{�T���=�[��y���:�G�;;�׷�`�t�oI�r�덭��V懎�nN^��)��u�4]h[��v:v�k��N^L�V7�� ���kug�Ȭ�E���Ѐ/>8��cK�:��px�<��6;�!��1�W����$��.͝�=˱f���x8�gU�7+�\���}�ܻ�l�Gh�;�xWqX����Or��c���<���.ۗ���q����>�OcPvP��u>�wn�����ٶ��^�ۇ��t�h�Sٹ����s<s��GKĽ�Vm�>��i���.6�ݻ�;�X������c�爺|۵�vxu��n9`D���������h-ݞ���[�=�r2�';E�30]Kڧ�d��Rsq̼�e,�ݸ�e��vu�&�Y�Q�lͽ�xA�����=wl-�	ccv��X8�hz5v��W���=N۶ƭ�c�k^�s��e�b$6ܺ	���=��ѩ+�q�x�n"��z+sv���q٨�RNrVE.��9�@��h�<֎;W�rk�c�v��k�'��������ga	ݮi��v<&[�\�Z3y{�cs�s|.מ�G�s���`^�J�x�sf�r���e�����Ŭv��`����zֶ�7�=h6:�,8佹�=�"��1۷�|�n�s���D�q�Z�ccv�эn.]��^.�;=.O[qvK�����ݹ��n��6�6;7�]t�A �=�Q�f.�;�v��3��u���T�c��.צ����V�=�&�]�ts�rgT=��aܽ�;	I�)�1��[�i�#͜�;-����YR�l�8.E�n`���eb|u=ō���ٷP��Cs}t��0�\���֙��ݸ���y�Í�?��n��a�` ��:읎-�ͮ��������}��k�hY�u�v���8.��6����]3�Ln+r��'7�v�����e��踭nL���/f#��u����]]0Z,���Wj������16ƈ��|�剮��.z�c�v�'��;cە���t׍�rZ ��l�Y1�ݵ��/gMm��d�5�}��l�gj�4�Ƕ��'�u�8͗�c�-�C��ϷX� li�մW���^����Ϸ=�͑ǫɮC�7l5�N�ֱ�5]s�;�����mr�vr�'�q�a��ۛnR�/7��qF� ���v2��f�[L�3�u����V��2��s�t�HYlv�ct�n.]d-���F�9�������b5Jb��Q7y�� �m[@|���/�r���+l�cމڑ6�Q 2l�o�~$gJ���9w�P���t�<@��f�>��{|�S $ܝ�"@(����� �mG�¾3L��g$��7"�MQ4.�5�_�����O_���o�}�A�ڶ$��λ�3NY�!L� �具�ܚ�(M{"5�um �@x��MI1�y���n�۶.h�NĨ��h �4���;��]4����2Y}�޼��jk���xG� TI�;�0%޾S��	�w��V�>p�I��	��`�.P�s��9�ދ�خ�շ��Y2㔹����n�!p�LHޔ�%p	/�Ia�ڍ ��o߷��=Z�)gSt�� �}��aS��t�JB�U)�����3��+�*�nx_�A6?M�c�d�N"�Y�;m�q=��������8-���!���Ɋ�w:���L�����Q��k��_$���Q���fb �"�:TA�^'~U�Fq��(c�K3�.��$�/�����ߙӾ�.�K��8��$9����}ّ���B&����wG:�W�>��.t�RI'e���n>��@�;��D�(Ȫ�I ����9fD\�2X�J��~��X ﺭ���.��z���ު��w��}�~�� N����_�k
���m�hAE!IFXr$A!K�,%��Ɏ��Y��e��lz��^�������������T���3�u���x� D��p�g5���I7��x�1��$c������Z�D�-�#wi��v�K/�^�a�ْ�k��m� }=�"{mӝ9��}�Y���ߨ*w�\р��3%�	��f�|��'��W�~$��c�s5f�\�;�rªf�Wm��jC��DwM�+��q^^���X�������Pwōr�G��������������ͲMM��.�I|�I���"��]�)u�'�ӣ����=���<� ��{�n"�#�\��#�)V?���tI�ӣn� b��a�' RHӺ��uܲI'kϷ�>����WS\����3�:��l @�<ڑ��ޥ���SSTI ��a�΍b��Bc�[[)��[�b��\���#}�E��X�L�_n� 6��l" ��1�y�jc�Wo��a8;=Ҭ$��:X)F\H%գ���X)y��5}�f/5�OĀ}�ڍ��_-�}v�$m����ν<��x%��$J"�m��RoK��),�{nD M{
�=��u?#1���I�����<C��%�"a���۾Ⱦ˿D�c;��
Y����:�@|���h��?>�ȥ7U��U�:�v(����6��4y4knQgY�Gm,ILe�؜Q2D���ϻ��%�*H0c:��w�,~���gĒ�v�i5�f��W�$5m_�mȀ���wPj<�V�oz�?��ٳͩ '�ݙ�m=�����E�cWg{l��n\�bxt���ؐp���=cv,F�Pğf�}� \�I#Ok�z�]���nzy��>~}٘s��z�o+\�Aw���6�ٯm55`��]�k+1b��=��$�DrN���q���#@Aٳ�4�@�������gՃG�9�NЖ�P*�Q��2A*��q�� ={� ~��˚Q���� 3g[�"��vf �^W�UADU"ڑ�-�J��|.�_)�A,�}w'�>}�� Y��L�ŭ2�ޏ-ti$�k�F��!�f�0�wke��� �ڶ�ܹC+�E��|��1����Db#k:�AV�����q`�0*�5��zA��^��(��^�Kԕ��i��R5,��1�޸Rn;꾊(��8z�4�΅�婑��e�&z�GV?��۸\��V�Na�KTn;/f:q�s�6�1ۓW�b�cm��=�Z������:y,�ے�dݲ�3��H�+u�<�'��ѭA�'���7N��_$�6���q��.:�c������n��k�u��Y�t��[��ᣏ]���خ��sf<{'F�3mǅغy⽋���z���q<���M�Rc�rz31wl�p��x����Kq�Tc*]����Ͱzd�T��]�7���۷f���E7W8:ۍm�J�-��G�W�$5�}.���@4Oc�hD�@��I؎�b��r�v�I+���	�TQ���"wV���`Mlz3:�� ��sx 	Y��DDv�w,�ï�J��9�R��֜�Im�\�w�s ĀI�u[@|	�Yw�'w'�π@??vf$�@-��ɱ�t
�TmHL�K��=k�uٷڳ�� ��<XD�?j
� �y��-b번�Z���ޮ�a;��rD�2ۑ����*$ ���p��O2+f�9sp�rq"I<�eo�_����[�>��C�O+��׬8N����l�۵���q��]tcs�]Wd�
QF�J��!�f�10�y�.����Vm[��\�gU`�G�-���uD�>��K�Q���e�C
�_�Us�D�u�f�rWM�k02�\��/y�p�Jǳ���q���*���Ap����H�H/��8�"��hK[�J
냖�Nߌ�0ȹu�)��/������ :���/u��b�Sh��6�r������{(MR���)�;��` 率��������M:7�=�@ugSa���4�ϔ�6�H�%KU��ͮjs�_��r�׵qO:����7B��gn{�s���K�X�Rn���$��Kۏ��i$�m�]�g��չ�/*�����ۆ��"󧬈UD�ؽ��+�&�� ~�5uӉ"�����)�Nq���c�h�;�v�yn��G���Z��F�v�$J# M��	��v�  ��֜�	~}٘��6�q�ϲ4�<����ζ��Nz��
F&��z]�`Ēn9*F�UWfʿ��D�~��� /�;�� xG��WS�V\�IS=�q��a(c�iUk�D��z�^}��H-+��C׵�Eed�+:��՞	e�c w)o���/rvҨ�Rc�q�k�'�B��>�R0HI�j�$[���*�׾�B~�|+���t {��� ���٘.2���UU5QNٜ�9��ݹ��u��Nb ���1��Χ����l�ؐ{;v�߱����F	.�w�@ľI|��m���g^^^f�����1��W��3 Hw:��)W�����yR����߽�77Z���s��=1�u��'v�k��<e�Ld��RO�|K��(�]w����ND�׼� �w:�"<����'F�n" b��$̕�y�M4%T�d��6�J��<�.Y�p�4��6�A�q��%�[Q��w�����������1ݯS}�� A=�V�"'�ˆ�<�.^�>������� 's���o���@��Y2s���9	&��oآ '���� F���v�ݟqup8���w�\|��Jl̬TzΑ}�w9{x�e����;nn�؇��6��y�5���Sz�ؘ�ƶ�9egx��B�eL�߀�}~9�K߿f�`I}j����\�(b�v�F~�M�@�O�׽u��9՗�@%W����@"{6��>5��	�<�������6�8d�0�l���e��l��d��8���+%O
???~�7bT����"�ݹ�D�u[@ ��c�ymz��D���S�4�31 I�t�Iz�.�NF�%�.�%����ϱ{=>�T���sŀ�'�����o� )w�}��m�?p^�H�MB�27v�ޗ$�K����9�p����=U���@����[z���y�)>j�v�]��a͚.d�s4I�Mr��UQ&�$���������n���(��H%����%+]ض�&��n�8'N&��r���e�h���� */y����|h�<��\�v�ps.
Ն�5�q�Nk����N	�K����ڌ�8���������w�P	�g(�� z-Gk�wɦ��W�fl�l�mjL�5�ד#���3I���=Xۑ���o�{h񹍽���8���ФR�:{c�����OI�t��W����TPŎEK=���ƧT7]������Ϊ�VV3�؝b�u��힃a�8s��p
�o6�nα.�]��O<��c����Ϊ����v#m��Y�bn.��P��/v9e��w�q����������;;�l���mή�(���5���۰�ʹ�4E�d��?��~&��C!�_Žn�C��=c �vf��b�(�Ǟ�6 �{<�q7�B*j �����z��I&����G��ھ�~���A��>��@ ��®����{BH�B]����K�]_�w�<Ә���{�>��ME�V�}��PD秛R@�}ّ����PQ'���)Q��b���nd�oF��@jKi�@���s3�Dﺮ}��_mH^�.�I^ו�!�T�H�c�
�^h?��/ӳU��Oz��nq&gc�a"Pۿnf$�Gg�Q"�˙�k�~���� ��m/F'jy�`Cm�v琍Z[����bdM4p��I���t�X�1���v?�5�׋���u�h#�mG�7o�z�[iI���Ⱦ&1U&��C!�V��r�$�[�}�ik�2v��N؍��9ؼ0YDQ�β��o��V޹F��u돒Y�Ձ��U4�:�F�GC�ؾ�:({'�TX����e�G�����[���@ ��~�a����ݩY��n����
��(E*�m~���m{��� �+�=�Yq���h	 �7ݙ�$�g�]���B]����JR-TL�~<�w7�gzZh�D���tȀ�m�`|���Ż>^��U'0t$��������Z�D�-��W`)7��H��紞�����<�rHc��� d�hQ&��"7ɬΘi׾U���������'��\j.}����u�1�iˮζ*�������s�7��t�9��8πA���h��s�Q3��gL�_�=�� �m6��5�Fq�D08c�a*�wv�>�G��z�y���p=^�h �g�R��o%�$.9u�.���b�&pH��5�]X[�d�I|��]�I߾1ߞ�V����J�Pwy2R�P^�[��NPDkY3C�ȗ���? X����1��%]�����K}�U��'0͙p1�]�=\�}�5���Y�[�eiy�AoI5G�5E]ڋ���p^v�I����-[���-T�y�Ht�R�G{X���#��"�X2)�U�P��q���ßP	����u�3��C�t�U{��Ud��vAvi�h�d�N?+�'�Of<u��;O;N<��w��Y��
e"�V݅���6���^�)9]l�N�6��o$�F���J�v��< �\�t���v��Doum�fA�,o�Guԗ�����*+y�s����i���ə�����`�ѡR=r��u+r��6�+�/�ڳI0��T� -(��\��~���J�ێ��Vϱγ�k�ͭ�L��%��:;0�ޞytʏ޵)����A�ϯ��n��'O^�,Rĳo��L�48�G�9q��^K�{{ծ�#�5[��vI8��3to#�p���7���
�^on���K�>s��z tw�V.ن���m��S�1&��U\��KY����8�a8�����޷�+w�¡���^	Ci�)���5W���ǿ+i�ѻw٣�1��4���ܛ;����!ִ�4�ߨ39�z�3�6K���r ��yܸV��GT|�M8%vT�:䣚�K
�kor��f�Zm;�-�퇠���1}�e�T����y{�o,�fb:, �cq0V�[c�Z
��+;��^_�xL�����}yo�4Fbpҳ8䰆����u���:��������wX�c���T`�V��1S(XŴ�DTb��%X��(�e��*�����b0c4�mq�**Ԫ�k,L�+(���"*"Ĉ1WN�Uj�UƘ[D��`��s3�Q-�kX��J�NeХ(�-�X�QKB�,Qb*��X�e\ʷ<cm�v�'���Ƹ����+iJ"���kh�(�lu@�[�1`��Um��"��,n&����i�T6ҥ4�b���W2�1�)�]4DPSFҔZX�U-����&!b�kV�M&��e���.j��
+4�(*�Z�-c�)Q4Ԏ-Y�TJ�s+ejc*���XfhQc��\�ֳ�R�5��KZV�T���P-�3,enR��.*MZ,q�e�ITkF�.�Xe�ܦ�E4ʊ�%bRň���ڪe.�+����b�5�+��ҵ
¢��
c(�*֨�.�`�JT�PE�EV�
&Z�B���}�D��M� �<ڐR=��N4�($����۞������*�=`7�l ޭcH����{�ʲɵSr]���T%�1��e$�`���V~$��&�MWd��z�4�ݝdCA�����Α��Z����>o�Y���<Y ��t������q�n�����-��=pu�㔹��������F�&�Uަ�A�l` �{��ɟ�{��]�{q�l+��@H]�ڪ��<���I��c�O�ٙ����%G�:=���x �zƀ���{����9Y��vI9�׺g$���gK�H�54�]� 5�sİ>��H9��|Ī$�h��� 7{�K�fÉ�#p�eW�w-^����w��~�| _��� 1�sx���[�#��}�f�P�iz�U�:�2{-��wuŨ1��^v�i��V���N�7\=�{����z�i�0�M�)5�$@��a�z z����UY6S��R2�($���߽���I%7�(�3X�e��wR���@}��s1�7�*������w�lC�Ē$T�����	<g�*=sbNz��[��n�t���~f����Tp$S������-��K�}��>[��s�/\�r@��]����6�Fۅ'j������%�G?z�t�va7�o�����H���f [�� �D{f�z]vP���[���Y�>�}$
&��'�ٙ�$�W{j�"/%3ܮ�3y��L�"e�s1"R��L� ��r����2s�������ן` �ӵI$r���ή�@4k�;�'A%��Sg���8eՅ�w.�I�~�iˈ�r=M�AY���+}��� ��nL�LoS��|�'9�Y��9熊#\(��z�P�����c�d��q_N��3��iW<^�3q�9�:��˨���N�rQ2�[�$Q�=Q�M�w:-9��nhy�ԧE�<��^��cYxP	i)e{t�͞�c�V�N���]t�ê��}u��IЅq��ݦ]�V���g��1�<�R��n��틈��0��\�Q��7V�s�收��mzM�:��vͧ�h�r띱�;�W��;>z��{�u��.ɖضC�����m�]l[��	U� ������n�^�yd�E���cZ�n�9�S-��(]��QS^����n�AUQ*P�UY|�}���H ��U�> �k��
�=A�]��n#@���Sh��u.����M:���9�3*��2t�ɍ�7��`|
�u\D45��jHe3.�u�֌�z�x$��rF�m£�%v�����Zs 3�\p�ͩ�u�1$I��iAm�뿚���!@�a���{}��ص���ͬ$�I��  ���^ǽ����5�.�zoK&x��Ĕb��W�R�݇"���x���9�_O�9p��က��n�D��n#���f����1����)�T���)0An#É����q��ۖvy�z.�v,��h�����y�Y�mm��7M�g��� ���dG�����/�-�ӈ��9������(&�a�]X
����I*4���^���&��j>���.�<_K�y�6fE�^�����`����;U�Ɍ+�m�̀	��/Xλׇqnl~X��Աe� 9��� '�{3:5�_�������ɜ���%܉��E�����<�X%E�'� ��	��6N񭻏7=����=ͪ <{٘���ێ3n�+-�J����=��"+��t$'��3 }�n}j�W�C>I ����$~k�hI��c�Oo�0bIջ*�J�$���F���w\�>n=��@ ���w�U���k��_��VAqF�%�T%B�:΂r�5����>������^���v��C��~��߁�!����J]t��ܿm�ؗ� �m�h=�1q}���d>7oʈ]�ۘH���2&��� �^:�]�)Sh�M�1;Ew�� Ǽ�|�7�.�)!�武���vC���@�U��)M;i~��` ��{���$�w�V�֘C��Q�N*7�m�Ǉ{�,��U����՝C��ioY0>v�E	�g ��Pme�K �۝����A��q�c�Es��ɀ�~��H���a/z�.�M6�)'6�<$���h�^b�HS|N�N�4�u\0�a�>@W\A�3��I}ݝ���w�֤�D�1�"VSޔ ��{�-��.w�Y��:�;��o� '��o��l=�՛�f��w۵��߿��]���àr@d�dRMŷ\<N6��<&�U�e��$�>�x�~�u\CΧ ۼ|���m[ z�#ܮt����+;�٘���m ��S��#�r�䡮�I,噪����=�{<�Dy �}����mYBW^@�U���g�^��#��"R&��E4����n�  �~릀H2�^�X�Y�[�I	 ѹ;�A��G���R@��H��,4J�˫�m��(�Z��*��ؘY�y}V�@��`h�׼�݇J<���Yc��؃m�e^�`.<���M�Rt����i�
��:�W��h����.��,�"����dP�WE6�F0��-���$��T-�2����`p����	1��t��폻*%�y$�{�A|H��*� >���ϒ�8�qޔ��������p����vۚܤ���u�1�;Qv��W�~��Ҫ��UU�"k:� ��[� �$ƽ������޷��qTz�1I�� #���eG�(�(�T�M��|���ɠ�~�ݝW�  ��:` �>�ȌH1��$��uc V�&p!��8[�%mغA$[�����}�Du8�~��q� �����_u����(�.6�pGl�n�DO_tV�Pݙ�j�k�#c/�]/�I/e���D���T��*���$~��>���.�
%9�r��^S��MI�=����o7,Z�N�����ۙ�@N�����ڎ��5���P����Zk6���y/��c>�NE��:�v�^S:��a{$q�С�S�9�v��^Zu�j3����M�=�݆�v�=��v�{n��n�]�9�{��=4���)ݎ��=�����"&���q7v�݄ٔ쉷]�e���2)n���Av�۲�y���.wl�����W���ɸlCڸd+p�ic���Of�������۲�[��t�ʧgs��W�ç(v����ɍ;��y�[ɏ#�]D��asl[����I�d���+�f��[<۞�β�v��-��k�tj��1���D��-HY;����Ґ����%�ӕ- �1��2I$���� s�S����}F�o�� ���v��s3i�!�%vszY7�S���Ԟ�kieDu�ۡ ��n#ﺛ� =v<��V�b�y��Q�J$���2['[�q�=� �@�����:���9�Z�@1�s`2O��{��[�S�	�r�quD�<�w("h_���b����0>׳�Q���M��L����$r��,�����њ�7��^�Y��^)Mb���u�cx�DDﺮ"�y��{�+��e�=l��2}��m��HH'n��݇cn��6��axn��婠�?�����`k\�������İ A>�U�@ ��y�ĠyT�N�y��$��;�=똒e�RP�����r}����5�
�cy����9�g��ak�����t�[:�=cB�
ɂ�̸v���/��O\޼r�S�H�qv���h�w���Jk��o5�$�o��@ 4k����ꍎ�VqO7��TMMTR�pN�_� �N��@|O���9��P �N�  v��z��h��� 10�wi��`�+�k+O[*2����� ����"c����)�Ŋ{-��@|>���B���	�*�f�
��Ӑ"7kİ6��v�&O<Ш�	j_"�O���`	o^�{3_�L�Ͻ�=��dH���=����:�s3<N�n=���]s����훣�?�b�EL�E*��o7M��9��r ����Ă~��w�_�ܮ���ҷ&�$�i�D/��@v,tosLO��թ�u�^��3f����{\�{vfD�횮W��Õ�F�̛�$;�m�1�E9n�]�>�d��$ ��|Dv֞�X�ޯu�^�����ǝ6�h��؍���|�'ފ����;�Oyz�{t����A�ｬ�=�xa�sCŔ��$㜬�\r k��""��f`K��U-9*)�J͵�b�������9 }��s0 >'}��.�":N�^ͻ�� >*�[jAT��)�T��m��b� A=�a�����M$��c ��3 @��l*�u��WrH�ME#��5{� �{`����j�@�t�8J"0�)����"O<I��P1&h�����*�]��n>�� )�u��;/Ӽ3��a|����5�6ɧV�6"�Fڊ	R�λ�i$���Ou�_���7�'� c�����U�"�J4���Gw�[���ZHw�܅����uk�۹�b% ���U��	/�wTx,N}�����  D�]���L����B��a-��X�Z�M޼�k��>X	 S��p�D���H��]��*�F�"j�X·V��;��_m�љ�, ���-x�����*�2�..:��<�����
�����I������?c�ͲO�{�0&���)H6���o� �<�u��WM��N�w�����1 > ��ľ$O�.�%VsC���Z�iQ���HJL�u��ٻ�[��VZ�%�5�iU�î�7c\�ae�2�yqF �&��'Y}�� 'wj�	��X�&�/&"������&�݉|LC���ha6��*�R�݋h%*��&V=�^m��'{j� <�y�"!߷*q=���H���.j(%C}*W$I;z��1n���Ow=@ O�i���%�[�͂���ې���.��gn5��f�_>�`  �=�Z ��nȡ)�x+���0�s%��e\R��UU�A�=�-�z���a�;՗~f�a���[ޫ�� #Y���A����ͺ�}��O�K�yZC,t��T��<5��6�g�ң^� k�p]1[�d5ǥ�>����8�N�� �v�A	a�)�dT�u�=�fl��4m���9ѧ�Zں�r��������f;ys1k�|�+���z�p��Qk��p藸��k��R3�	�D��usc�nĺ�J@	�c�L�;r�,�!C���U��h���1��C\�|�b���W���ba��v��}|��Ac禣}����,5l�wH�QO�7���^���8�c;k�kN�B)nӛ�]t%�Q۾Kx���n�0To9@T�fԚ�#	=�.�;ؚ��x�&����;��c�b���l̸���W
qPhQ�����26�#����2���:;7�5d�@�p_-�������{i�Ne�ud��!���]�븵p]��5�+����/S1��3yth�Pq�
ó��v�nS��,r��d42U�ͳZ;n���A�~®-�Фzv�2�}:��K��'r*�2Ƚ���b����Թ�$e����ٖ���r���b�j�b���ŝN�屃`�Gf�a-T�2�v5٘7sҕ�ZnDqFm�y[�4FL��2����{R�ݪ���i��Mo:����Yф�W8j�)puĶ[�NK.cZ���çM�|�͜��<��v�Z��ͼ�ek
PԜ���.OqT�2�j��1�}�x�����xC��CIK�OԸ]��)8n]
X4"UK��3;*C��������}ĀH6n��#��Z��Klm��e�#�.`��R�2�9TTQA��b (��m�PUԵ�m
5Y�X��lh�U��J#1��b"�B� ��-ieecmҨ���XưY\�0�Ŋ�.5��Q��H��۬�DPE�J+m��XU�l��.
�)����PUX�-��3&R�����D[n!Ub2e��\D�iP�[E�Z4�b����,TulDQ�W)R���D�ڢ��D�҅bUiKK���Z1�`V�%D�-B��EX���5!Qb���m
#-mb(i�AcV��n�U��Qq�YT@�"��� ���B�ۂ+b�m*2�J���QUV���ic��9iiYm"\B�q���K�73/$'$�v���hJ��`����7P���Y+�E�<<�oe:s�W�l��u�Żn/��c�n�V˼�^��6�b�,��&�p��c��Vn�V7m��q�3mvP�ۜVrS
�vꇥx ������pc[���cu���D�dѮ8��yss�Z:�:	�� �;��z�*��ڷ<��]���k�x{O�s��£��;<��ru�؎��s�ޭ�CE�����de�p݃���5�ɷ8�;p��L<���my�t��x���X�M�o<'ͺ6V����NWv�ۄ�r�<���;;cq�cn1n]���X�l<m;-�[xi��Ѩ7N�v.,ΨU���ڣ����\=�p9뵵�Z��yx��kG�v�{p�&}n3�=�'��^#!��gm�/]��p�mp�ln[���uq��ٌ[x-�d��beNv�1b�st�|g��l�ZMi��q��)/n�ї�7� n�c�װpL�=�օ��������n7����݌����,��m��˜�cM���s�s�r�:{e
��&��ܸ�v�;8R]���s�cpv��];�z׮1�uj�=�uJ.�#Ѩ��ף���.S3�6nr�����]��������c=t޹��3�m^i�KnN�۶�<1˝ڶ�^N�]�vֽ�m��[�q���m���2v'H۱�g�j��#ֵ.�u��蔭��[��������Nx�D�e���秠�fmX��kX�W6q͝��z���f��#=,������
6۵Ӓ
�pE�r��n�l��s=�8��q�̷6�Y=�M{�<PV��u�ێgOn!w��.+�ݵ&��.�$A-�g'69ۓ�ݷ`���9	G��4U�Q5tl�q����}�;��.P�$ۍOom���1ݧ��(��������&W�����\�㣗���n:�竳�s��n΀kL��[�:\���nhu\Z�Uł�����Ga�RqSӆ;u�7h����s���x��s�֮�M�l��ډ:����k�v����Y6��	�Bt�#�۞/]g���i�⋞C��8�n�.�9��[�`����hݴ�j�Og��G���g�&�������\�*�ag8��;�Cq��u�<����t\\�]�@˱��n�pW�S���̜qXsqԵ�贙����v�ݵ��-�7tb=��>9����m�P2v�B'C�'������� gkt@�_{�0&��*��>�M�D�{����#�R���n��K�{���=�<1�s*U��� @ 5�s��_{�3�~��)4���.��%�u*�H�&HT��Y�� A��kq������==������;�T@�}��π��|�	�%Ȍ�agU�k��#,L�a�v�@��f` ����9����_$��λ ]�$r P��j==9��?sݚ����m�k�P�P�1�@����ς D�m6�:jw�/U�M��/I-��	D�6� ���tA�(�}1�n.ϲ3ۢ���Xz�
~���w�]�R����3�=c@�}�>� A;�WJ��ϔ�͘����$ }��������N$���t�I%��-��u]ǳ�S����X.������%�=.]�B�}h?�ѳY���rn�0vk��v��q�F��/P4�U聗T���?u��D���vf�H'���A�sUU�os���ɗ�%!��8
&�	DT�����	�ڶ��V��Ǫ�{�'v^ZV�'��$�w��;����f*�
��Wy�$�L�2��R$ĒM_{�D�L���M��;�A�5Io�`:v_��%H��,�d�H%���}�ޙ(���S��x D��\D0����\��l��uz﷧$��B�M�W�D���m�@!;���P:U�$���L;O^�����ڐm��EBә\wn�bI$��Ҙ 7g9�w1�~X�*����ς"'{�l�y��)QE**���{��*q�DvϟlF�m���@N��� ��9��������{����j��߄��5��H�&��������B�=��˃���Rֲ�?*��s9���û�}ym3n�ui�6�>V���j��1�fk��˄�ׂ���z����:WaW���ɻy��$�{�V�7L�����A(�(%�[.�<^�y�u�+x!D��i H��l�%G�7�a9-�s ͯ�A;�K���/F�Q7��d�UX�@��y���x�~��\zm ���h"c٭�@7���@�"&�l�����|M���ݒ�Y���[8�ѵ�<+m��hX�L<���}����[k���D�"@�?n �)�6����{���2�]�I@-;�p���kA�#P%	7�Q����$�G=t�R��jO4D�/��o�٘����wwQYy���K&��J4�ERS��q�u� ~�x� 
[3W��W@��k؈i z�v@�;�sx��݄&�\0HcWi�t��[u�z4|�$�.9�N�	�{s3�@���5�ސ����;Z�J})&N��*�A[R�N�i�V\`T�eާ睛Sn�N�:*b��DB��^r	�G�H�}�t��ˊ1#�0EM�k�٘ �{V�����_�=��j�=��:h��������Qv���w������0��P �q�1�f�Z;e�u�㽶�%p�K����q)S@��9���~��rG��fm~D�����Ē S���A=q����]���m�d?{[ρ^'3�D҉�&���g7M� ]8s�q���*���ۙ�I'���7�]�$��J��RF����u1H*i�1��f 'Ϫ�D;_C=���d��{�� '_K���}D�n#PE%;KO�����ڇU�}(����@ ��m�� �H�=�Sf�\D�m� �^y�@K݄8��"j)UACh��S` ���Zw���S����l�T�Q�I�M�ؕ ���{ͫ-��=-:����\ָ�L�f��������ȪPi�s��T�&�"���7fM��B�c��滳�r�=����Q0�N�F&��6;;2g���<3 iG��:UɎy���np5p��7\h��	��tg@�N\�����z���a^,�_�����Ý�;>V��;v��Y���%3�t�n3=c9�2�f�h\�O����\\��۷6N�|��X�5����:�O[rV��W$mZ��YZ���6�\L�q��Ex!ے;qX�un�v�5��[]���FS�X�� mӶ�����OYL���su��ߧ��㪚�Q9����q�"'�մ  x{Ο�^��|��uO�nf�f �G��[;G��C
AI$�Iv�5�wI"�Ֆ�����>��>��� =�ݐ!.N��/9�{BH�i�Q8%8E:f��l�݀ ���S�s-�_�#P�>���H�f�j�=h6�f�Iˣ���s;k�"���_���ݻ ��u���t՜���vwJ��Q,ۊ%IW�����oU��tAڗ>�H��$��;�Ν�	���k���)!���n����0x�Um���mwb��R�hs������{����q�f*($-(���(�sٻvHw��x��Fc�ι@�FvoX���DP�ƘC7�;7�P3��%�eL�`Hu���;�z��V�d����Us�w��Mwq0�/
�ԁ�W�+�夔����r�hmm5����y����@b4�L�I?���O����7`�́��k۳����d0��H$�zug���v��IFI���Z��u���;n�����w�#jŧ�D�,�"R�ޕ;<��ᩌ�ӫ�,�� \��� ����u�07Y�=�=u�b��Ki�	B��j�wD�;�͡�&���{[O=�* ��uX ��r���(�ܔg�>`�UóklwJzy9�c9^�q�lj���90s��g���P�3�y�G�B�����`����H%o]}�D���mZ4-c��wd��lZ��
�p�����	w��\��m��y�Ԟ�� yf��fl�˭�3���H���60Z�F�F]�6W]�	+�eA ��,m24&s�{�Cus���r8��Fݼ�s�X�V��<�B��Q�g�>�t��Mf�a��!��X�9��W�W��$�n�$���Q#|.�nHؒP.w\���=h�O�d�� �W��h U=����T6.�SΡ�5�_��H�*'@��`��J$׷��S���W�#��#�g�� �WW�|A ����59�R��obx�m� ��̜��
Y�c�H(�<x�B�&��4�(�����?Pi��S��Vw��$���Q ��/}�H�z0;���$�oP |�٠w�"�H�Q�T�7՝Zph�����y}CI'���s�z�p�:�[J�5V���qA!iEE��DЧ��HC�E��&z�� �ϴ�.��y��6���Q��l��3"���-�z�{n�b@PsfmP Qwj*�OyH����\�g�1*V:}^�X��q��Rق�m7Y��ѽ=C��&����#���J�5�������vdy����A]�����dM�%շB�w��`����vYd��Z���V�����+�uزJc	��r=�c������6��pxŸ"����l��� �u�rzTN�R%({d�� {׾�T-O{PY�+�%Ӿ��>yw*@t��p@�9(��]��c�c��j�Zr
�3/���Iw��:�x��ٛ���� ��*F�F��).�;^���P�;ھ �cz+Z�ͅg�� g_��K�wX���!P,C$�T]�`�O5D��3���� 
����])]p�8�zHO7�s��a��2��eu�ĒWV������m�Ǵ����þ��A^��W�2��Z��[m���ov�6�os-���X��.�P;s���3Xgp['�*���I�"��.�=b�]��Ilc��|K����iyn��:���ͺ������;^�H\�3�cv�jW���î�GV;v;#;W�{e5���Ӯ&�	�u���Q�``���#n]�xw=c�����;y�ۛ�"����8�˶u<Tk�y�3ͽ�E!�euc�˲�g�3�(������qkڮ��ڛ�-Y֓E����ص�++
�㣛n\��۷L]j�M��cz�3^�v�N⹅��x��7iy��	8Lb$��x�D�&ē��iR�-w�U� Q���b، ���z?v]�A��۰	�k���H"R��3  ��[6ծ;,�'g�/�ػܐ$���t�	�B�E���rH��a ۋPh'
0S���޻�Ҿ �\7��QN�ܨ 1OyR�(����
G$����6_�*^>쪽tH/+�VO�PG���}�����|�z�v
�q
�2@`�E@��(���|������v�IP@P=�>ڠ����}�Y�^����DK�	 P4`L�n�W���ksvi��0�V&n�jp�tc�f� �ެY��  3o � ��n��ou;�٭O�Mi (��h�K8�M�alI(���������G�mia	Sih����WfpU{+�9����NB��2xX����HaK���f �0[�Od�8���-�0K黾�A$���(�@���M
��;�o��ǵ�l�h$me����	�J]��r��ӟ�!�G��OP~�����`$���Q���u���	�
�䫭�X-�f_�]���wo�%{v
�P�9�T�V��+����Y�����Gݪ���9!�ʳ�~�	5y�W��-k���P�
O;~��G����vg#�e���A���W�cbN|ThMج���b�`��(��Ď\%�;%��F:�q�����!hh�$��\{��$��ٷd	��u�=4��u=��� e��M�gU��c�r�$I�e\�]vў�\�{��
��ڀ���Hx绸��U�QI��	�4\8�6�3$���HP����� P&�Y�>Z�V����bj�^܈�awZ�Z�ۇ9hW:��2�]|S}�.��]ۮ��9���ݨ���ܲ���^XX�%{��M�S9yLt4�D��5������X�Y�Ы�W���=����f�LUA�o��=��0�"����C���X��nR�*�e�,�rA;-e^��Y�������Բ�Y�;�-������/t��v�WG�$��B���� ��̇�F�T��� \ƻ����.��@ĉx���͟9�Ζ1*�ݽ��ށY۫�ض}Ɏ�ڹwG{��Ĳ:`j�ڃ��v�Clv$5#���}\Lj-�	�Q�¹{�=R�X��c4�/Qm�ټ�-Tʨ������n�� Јf��T�Yʇ<�]��4�j��EIo֣j.���._pwbO\]����rM%�!�w:WJz��Y��z���&c���e�p̦����ZGU�w�r4�N����88�ڢqn����S��o^Ws6���w�����c�0��j�5VRYb;y��׈���7sX�F�p���y�����N��v3�����U��s�B�}��˔�*��cC:�.�h��5n,�����FYr1`Y��ir��!#cr��(�VR�`\kibܗD�֮��g ��lm��]����3��+���x�[���6+;��{���9�I8:��<*so�6<w7~Se泻%a�f=�� ���4�M�Ƀ�7yͻp�^*B�Q��xF ���S�c'n�\)�IE\�U��ꕞ���M�Ѹ��Q��<�����k���U5k5+��ZÚ�����]��(�q��c��5-Q��cY�b`�ƣ[QkQD̳J�(Զҵk+ZTC��F2������Q����\��q��1Aj%�wj�B�FkW-upb&��U��ު:����5p�J�USHQ#6�V;ى�V":�EM&���򉪵MT1�1cZ"�T�Qf���Q`���u��e(&4Dr�T*�Tv���PFҰb�D\���j1Q�Y7n�]%�Q����*�h�����
c�Smej�m�EE4�EUe��J���Re�c1ޮ�EQF(�u�E5�m�
�VՊ�QEdSQ)��R#��4�T�l��)�kX�`�j�c������
�EA�Z���T�pȪ#E�5������lm�+1+EV*e
5*"啎�UTL�]QiR�R����kZUm��V�R����*".%�UY��Qq�b��UX��R�R�ŕ�\.8T�QEr����o���z,W#����Ura��y����K�U �.G�/m:΂AO+�� �k����/�:j�rF0�����Hn-@�S���NL��A ���rTn�v� Z��T(}���| ��h]�(d�;V�'�1	d�N���i�oM�{<۳�=�v�g^�c���a�8(Q���6�Tr79�2��`�k3z��H%z�~ˑV����io�� �߼��
04a�J*���|Et;��s§l�� 
�>���h=��YX���;˯G��1�2Ԍ���b=�� ��+�`�E�w�ڃ�O�,+s��J���H��B6��d�^��7+��՞�>�Pz�����mh (����EA		�T�"��y�ѻ
��U�I�FX�j��z���ẵ40��X��Jj���kr�=�`Qj��V_iy\�q���n7�fm%Ċ��w�'ׇ�Ȓ	8����UJ�7oz��uf�w�.N� �l��iE�J�ylgx�*Y�ǟ�D���C1�Or1v�V� �����(�:�e뜙�/��vv�A�S���nN�{��B���>)E�$3���D�7x�sH�u��;D�Q��p@�X;�αd��uk�6D�oW��}@�� 
Q{�A��|0P�uw�hO�B�H(���l�I���$�t��γ������'�	����~ _�z��Ք���FFSH˱ޱ��>���y��m  sS�6zy1�Of?�)���T��-�qӐ"��Q{]wV����X~��V������[� t]�Tl��9��~���hq#w,`���Dܩ���W[�H��Y���ܩ0y�T�R�Kf����*{ϣa7,#��E^���+���%7tP/��ϩ���w�~Oh�9�v�1��m��/j���H"$C��C��v�vKJ��9Nxg&�9n^!^75�S�v��ڌq�vz�����&+����<�܊��fz�l����@��{p�7�ά�v����ힻm�yUv��&f�/8����\�$�ƚ�h����n\Y.:�t\��;�&�N8�ZX���l1��]�{m0t>&p�k<�Ω�Q�x��s{Z��5^V5�:Xqn(�$�3�=,�A'��z�U  �]�HPg��U��C1N�媅ק~$^���ĕtu2�N�-�3z�I�%,����Z/NGe�]�E[=<��\�F�r5~��i����M����
X����,�I��uX �1Ё������n:�����g���
/7�A��DbQWż�xsZs�B~4�j� 5�y!B�^�^�����y�4.o]�H�R��h��iv#�� (�vh߻��~8z��@}쑥@}@	��`���W����.��NӸ�j���M�n%�k@vnA�N��7|��(�vqպ��x�v�F/��"� EC$���v~�fﶬ�I+o�P5�#H��u���$�&o����I�eȒ	8��:�WĀ���ۻ�5�U��	���"{t_OA�߁��R�-�s�W۝}O*�ݨh��V�U�)�ɼ�b�%W
��5}�?��pN���j�^B�
�~��$���Q�[��xtq���owĀU�Z�	8!Q6���]��?�҈ �CD��w�� gI䪀�(^��
���M����݃��r^<z�(l�~l�ھ
-{kh
l���C���h��%<�2T�AiE@������c	�3*h
��ʕ@���B��wU�&�fb�YFY�p�Q�2Z�F���h�@���c��t�[����i�I�z:�]m����v.�F{��뿉$װQ$��w�ϙI�G�N�5���J��^ͣ�e��c��P.o]�d�X����|��( (�6�����T ����W�]̌�l����	4Na�Ϊ� �n��'�:��{�8�mM��µ�~���Z*��|���fz�ac[���6-=��I�<�3g�&>��w�Y��m�ɚ�-���)�)72��I����Q"���`���z�	IQ6����C�����z� �o�~$��� d���z�.ȼr��Lś@/�m�$	8�n����Y$��U�kio��N�S6��Tڭ���*@T�O$-����T4��P��-�T0�a��o6�'^k���wv�r�<<�ؘ�a�������f{\҈%�8����n�X'�G�]�$��E�7�P��\��(��䀬�e_��i��mv�޻$���!7����>O�+@�oJ�	k���#+��dA�^���?L'��1d�����'�X,���mX�nq��p���Y�$�o�샕��H�Ę�܉ ��˰s�@�=|�*>�c�PA���  �<�@��@3|=��V�·�9�s�eu]/C�0��~�[.m�V��(5�����D����2ŉ(Uri����H�b����{�~�[�r���1���˿�J�0CRDM�(�g��*�镶a�h�p9�Ɩ|�(��6���V�����w.`p���_1
:�f�ܛύ��=���x��qu�|X�2���V�z�"Z�<;���IR6�����>���T(P��߃��s�$?�����=�����&9"�T}��$�G��w�u�I��uY ���_L��x��{��Oq'�0�1��2�I�h��}�6� xnkK7=� )崙�?��+��1d������.oY���&�%��yj� (�6� )l�"I�)[���M��d�Aw�J	H���˔	$�޻��72�#w7���[���u��e��7�S���n��8f����.�k�K���]��c�j��kgn1�����A����m�r Sw/Xw:�ZYՙ}Gc �US����P1a�0���83�-��y��1�ݗ\8�œ�a|a�׃��Fqr/<���ջ{V�p\,�grݖ�f:ݪ�.s�W�����7+�젝��I�;���y�q�\]ۮt�1�<���&�G>wm��h�#�7��u��k�u8���Y9��;e���)����>����.wC#�{qm۪
y2�ڻm0�Lu9+�m�*����o'p:���{q��Y�+�u�<���h����}{mD�i�%^�P�	+��_~&뷮��t��I������ �$͠%w ��e�]��觕 $귓����{�k� OP�I���L���n���%<�B�c� `iE@��(A �wm_��41>�]��t�@�L�h
[��c�>��ٍ�ѕ&���'�V�%^�	��˔Ak{�� ���t�1�9����G=e��}!f�W�����3Ӷ���6��U�?F�+���y/���ҴT3���1�6J��nl�Ǉu���VԳ:m���q�b��݈+�:�ݱtC�9&8�"H% R��.Q$u{zŐI?d�u�4{�ے�4}�/eI���O�]������rOgfW� ��W����QY�],����M�z���z�T3#�ҵ:�V��Σ+�g�z4��쓕�{����R���֧�Z^*��3����=���guX'�rgu� ��ʮ��<�:�,��&�R0T���w�;~��?Lޫ�m���Z��]���>��r_@<~�@Qu��`�$@�Ҋ�o�Urﮉ'j>J����C�ޘ���V`��?gr�{�7ń�Q�є_�W ~]��ow��u��A�n]_Ă�7j� ����4�졺�~zJ���LF��A$i'�ݹv���sKٻ����2�F�EB
p�I�x��a`. On�Y����B�+{(W�5n�L��T;s�.�]��f��>����܉ ��K�s����_������.�u|(U�<�� y� �`t�[!��7IJ��
�H
)�����]�Oĕ<�h��ۇ}�Eef�Gw�o9//g
��C��S֭5�����[��<r�9�]�.vK�=����؂z�uf�7��#B����6��KkO�Yc�$���B��D���b'JF�w`�ܕ�4nmuX'�
�eV� �w��EѨ��3U��� {xL�Q��`$�om�V��H�|N�� (��
{;ʵ���-�8�0B"E��=�kaa"��Ϡxg%�hx(5ӺF�����/��<NSKj��	[{(	9^ޠ���.�=��$V^� ����D�8�I@7��f��W����ۧ:�������� �w�/�^A�_�����i'���$��)vs���'kw�X ��>w��`݋�Ow�|yL�@q{ʗĭ�� ���r<��q��w�� H.��~ WE=���?y:�s�ۘ}�i86��w���gI���\�⸞� t��u�W^�w:�Ń+~���eu;k��5�urw���~[�n��5Pڴ�/�xW��S�
��ub'JF�v:�ݢ���^���4���[�H�mm {��*�(��K��o����l]�PyE��HCF5$*0bQ�$��]��E����Nd燵&�� �0`B�	�'}�H�r$����(����u��`�~��벇	�l�(��䀭�	7�M��-�.���������v��x�}�{b���=��/����E:�<��*��~�fC1p�(�wB����,����"<I�ﳧ������
���J��	��jPT�n2��Z�l_���uǯ�AޮʲA"vo]�IU2������֕Y0`?fef^��� ��t��L�ED��[�s���H{y���7}�[��$���$ I?�@�$���$ I,	!I�`IO��$ I?�H@��B���$�	'� IO���$���B��B� IN�$�	'��$ I?�B��$ I?���$�0$�	'�@�$��$ I?�b��L��9�6�͈� � ���fO� �G>t*� ���
 �*�  ��E � �  E
�R��PR�� �P
PP
�  ;��3Y��EU�IPH� �#��eEEQ���Q(��D*R$��#B�Z)��U"�J%6� �UD�DU:m���                                     @   �      %)}�A˺J�rE��:����j�j�A��}�v��oJ g1�.�z혗�;޷E�����Z^c{۪�y�J�R�Ѷb���   t��|���ꗘG �]G��ۼ�*�bۑЫ�� :]��� ��49��frҮ��y��^�{ԝm���IA�&��  �        �/m[qvŰ�k���r�6��񻷑�/xw���*�s��U*9j�Ś�v�9�����J�� ������P��PX�E.ę5��   J� Х��8�����
 �(�R��3�P��S�(U�T�S�73B�JN *���)�Х-RS�g@^Z�)W6N}��)C}�5$�)SY�  �        �
��������P���*�T)ze9� �. hm@U�8�hr	Y�,  ��cUq���i�_   ;��ҩ���h*���j�o0aQ��/fs�T� �N��bNwu*�r�R�r 9ɡ1�*z�M�  |         w�Lڋ�J�h��9i���Q^ۀh�aR�&��/z�	�W��#� �-�������M���5)o�  E��,��*� ��*�D��B�s.���W֯m� F�d�V	���{������1��@!+KiK�           :��=��c�u£���on<�R��p `���;S�O/N��[��z�qǐW� �&�W1Ԁ�v<�v�v2��  h��Ͻwy�N�6� n���.w�u���� n`�׎�v�+z� �'m��j��ܱNͪ\�v�z�y�uπO&���A�� O�bJUM4�&CO��J��� D�*��P��  �=�&
�H��	4�I���@z�b�7��?��� ���������������$ I5~ֿ�H@�l@$$?�B�� �$��H@�0! ���?�_��3��4:���k9�{�f�W�dd��z\$��p\��o���\�œz�P��%F3�Rl=�N����/g�����5���LX�F ��e�#&-�RY�j�q4ܷ���l�9�>�1�v6
y]A
�[�9���˴T�D�,��R�p���-H�r�{��1��8gUr,�sFs�f�Y,����SQX���2��CU���)�ifo����;�l;l��uv�X�ܽ�ٚ�̀f��Ѐ
��&��\|�L�s�$��n�^(ڒt آ���GnC���Eŭv���JY�Y��02�� '#��ݷ-b��v�
�u-�[Ó���d�{����,�H)�8LԺ� K�x����+��'�8�����-�"6�J��"W*}���è�&7���T5�s�s#�&LGk�.�;�E
���AB��j�xuZ�U�p��S3�r�Q������d7m�nF�č�ޔ��R�Z5�@�($�8��3��Cp5�X��ޘ�ݏ㽋u�/sz�3���h��
:��[�E'>��k��gp)��;Gt�ZJ�iі����#Z@t�n�.���3�)ܟo�zR�^�>s.�-W���E�* C��E@�iN���Н�pwz9��i8ߑ�y�×f� B��8���{���'�ї G�n3�d�LӗM��5���wF�=��_�w�9�R^j�-�V>�(�R���"���]�ћذіH0��T���}\�CM�-��q�E`<E�����E"X�3���!_\k��,K��X;��k/�hS��U������m���[�Ŵd}�<Zu��{k<_t�gQ������U�Y�i�w�<�M|;[������br`�Q���*���D�sl&����q�g)�}��ǸI��)���vN���H���"1!�)(b$��E�ͺ��1��.�4�Vh�]����l=�z9ԸJb#tQ9���_k��{��n��+"(�o�ɣ�pKm:�Hhp3].k�3�f��a����b}wW�$��1�t4���J#���e�.�H��ʒ���n���#6S��46�Ʀ�M��,�2A�����۔�w��ڱ��D@��2�iJc��Z�8�㎽|�f�9��nA����N�Rt���k���l��d�'�{�5��Ξ���.��e�gF�͌;�ѡ�SQJ}݌��qK�*��z��OJ�q�r��,�Xk6�2�9E&���!t�M�汥��aˬv��������ݳ��rn��9�.���t=5��+�$:��9pܝ���.�Tu���>G�`���o�+5c�˻�7t�S�ᯙ�0d�/Jĥ���3q�ݺ�]��Ԉ˧7es4�nEn̴p{m�΂�	9��5����K��뙨��䶅,Cx�uj3))������-ޕ��J��qhdH��)7bU���.��L��{��Gcp�iv˰�o��,36��K�4t�5(�U�c�B�X#]�:�Yr�$�v�;"�2$b�s"Q�=\�;��/>D�Z�G%�D���l�l�fDS(�N���J�����k͊De�Lg*���fΝӚy��Z�=��h s�����������:�k�D�f��4��5�Ej�ɈҗkI:��2�5���1[Y�S���k@t�r���R�C�j�6k!n��Lx]AyjTuOki�y۫���q �]���T=w�u��x�fA��\���́�i̭!��ٙ�ZOj�*�Xu)���qIXŽC�A�>o:��m7%�i|-Bol$�)��^�m��,:)藹�Α�*�ɺ����GR0Ґ��&|7q�w�(��)F;g�-݄��
��P�T0�i�{7�ԋu��Rg��5����_K�\���iM+F鰆C5+��6DU�� ��uV�QK#4�G�6����K�B�m�&�ZsR�Uw���r^	[J��[67�I:Q�lf���p��Y��ZŚ�k賡E���*5팕�u����ĵu�e����=5����`��+��17pC��9K|�x�PV��`����#ʓ�wr�؈��7�D��0!�K�S|zdk��7K#��3X�gk2sǄ���2X�q�.Y5-���жÂ"xnv0��Γ�4�����hm���3�#�JB)pY׷&�{�Sq�Kwp��ӷSd�����U`#l{�gṼxZw��n7p�k�0b�9v�������\nH��r���k��;���J0r���h���
�c�v[n8�&hg` F87�!�-�>*Gʢ�X����{4��m}A̎��b�{^Ų�w��X�����zʗ�����-�R+�ŉ7���ޛ4<�)��X��+��R����{*��gFJ�;l�#޷� qu��IqI�[aՋ	���y5�.�ʹf<�2��1�
�j,�]���a������C{���>�I�&A\I��L�w�a��!�@���s�R�1�:=͹�@�Wٻ���M�ql���ج�]<J+fdQ���.�HN�����˦q�U6��t�7��ᛥ��OL�L2<N�7T�@t=4[-U�*c��u�.�2e2��J�y��m��y����u'�a�߭��t��{rp�Gr���R��C8�R=�2g��<6��x�f�A2P����r�O.� 9�w\GB�-�`��:nq�!w!ή�.�t�9FE2q>��Ň� N.=��GN]�%ε;au\#.D-(ݛ��`�g ���淀���W-�gC��VӜ�����Ph6-�rJ���Aa!�T���of���qnq5���8P� ��\��78澙�MuȹR�\(}��a�3u�e5F(:#a�
�2�t�u��{�@=xM���S=9,Ӻ��c�$4�[t���&��U�;&ڇt��ځI�������:�뭢���B�G���r����9��ֺA����4���Z荺8�.F����٥}��3���=��{#{�s�W�w9���/��b8��ī"'K�$41�Q6�͙Z���KOd呴�7���+][���,�7�+`���Z�۸�Ud�CMe0�c� 79X�XI��w(��O\���n/���o ���<��E�qr#q�q�ݷR��c
�[hZ�yhX���` ���w_#`��]��&q=�J��� s��4pZ�䛒���#^G�=m�s��0���Y���R|�1�8����)��Ϟ#0Kx�'n�@w�L:~	3����F�Q���-K(�-\+N��[2�7x�LI�˫��w\Od�{�k�n�QYq��ӻo�7k�,�hy�&��;���ٍ�b�h<-��+/+�ݹ��}��XEE�&o��8��.�� X�t;�P��ݸ^���J��Րg$� �6I��N�t�
%��o�;�ke�P]6W�>	W�T�]���k�/d���(,�0+!�J�֌I�#�,`���{1��1	���\
tf���ճ3rރ��.�WG{V Eӝ�}��g�a-�Y���k֦�79Fk��`�0`�H"���=�d�YY�D���+&��]q�2��r�Ct��xvP�T�i}n0�B�n��\��cY�=�c��ֆj�^�T�Ŏ�#GX�Wt��bHt3{�M1.��`���X*��gsf�%�;�ȵK9�ҚC]�����/�R��r(f؇UVp�T؊C�ax.q��6�3T�TE�"�8���}�s�wvoP�اs�*p�uُ�{\�|�6������Yŭ-|��9��o>�y�0�:[.be����%����jk"�S�����|"�Z)B(d@ƈ��V��2��{Ԭ�M��� ݙZޔ��:pn��\�]��N���EMH�5��7�e��854I�
�Wd��2N��7Q��\��Vn�u]�h���������JD���P:�']R��*Q��/mn�ht�@X��V=ttlQ>�"(2�t�v�;:��9ј\W���3�u��;'Z ї�31�6޶P�G����@���7���ӥ�����r=�2:$r
�f�k)�M�F�#��fP�۲ƃ؀W�����ەf��hң���4�{[&�m�����ciZ���;̓���i8��-���rV�m҉9fC��b*�k0�>8`��5q����4�M��F4��y6�3U-�x.�(�_r�;%{�8zuV�-��7�sd���c)l�	&QbB��ɿ9�9|i=3�3���͉`����K�GvP ��{��[I_YxKhXt�!-�z�G��%nju��Jgw;ec@@wA�6��V��H�p!�v�N���%�Ճ���L�7B68��(�
R<q&s-I�kV(g�\�B�^n����jS�uŹ���6R[Q��I
�9{OBgKQy�.����1��vv�/4��iSX��.nn%.�wQݍ5z��x�^��݊l �)��77V�Q#�P��o!���Bf��u����s��.� �n��{ZJ�B��$92@����æ�l�J�U���.�4e(�����P�g\v^x[��0���{y$����I�<\�ŝ܆�ZzϞ�v�)��s�iY"b�-�����IF�Lˁ�7-˨�éؔ�����Zu�n�w,c��v%�V�Oq`o2�I�)Q.KW�fLbb���<�$�.��j��g(WI6�9�	Pn�k�D�G�	4�[�,��k/7������܏O\-�)[� �.Po�q��$�X�ᙼ�V�����Y��Q�ju��'َս��y�54��nL����{^�ʕ�SS)��w��}�\��vGq[��GKRka�MZ�(�K�x"ς�4��FU�L����A�z-�v�ov#ܺ-	���%k�:���0g6�w]��MgHn�.�"��ٲ}�r�]�!��&K��.XQ/vݝ�q1D�ж��K����ɟ+��{>�0��.�4Ь�9f���8�L0�J4Q6�ސ���Ե������g7j�(�<W��PB.�5\J�J��aw��׌�1�u�F4h����*��7���Еԟ];�� ww9x>Z���R"=Gۛ���w�on�*�=���D�vA�ZX�Hq���ܔ=�8	���L��]Y.Uj�(�;^9��o^�G8ofǶ0z1\ku?��JZ�K{�r=�]�.5���]��)�"�i��&�6��2ޱ���S8��i�k�IH���tv�����zͷ������V޳�1�����rU�*γ\K���o��T�%�KKi�gX�j�!2���2��A_1]�^/\r�H�+�U޴���[Xp�s&Q���}*U˵q���c3��)m�*E��1|��z�ӝ
|i�gq0�+����Q�����#%����b�Zdn*0ne./�	v|��$�z�uɛq�w�AnH济^2s�ۥ��tC��iV`��\�ঃd�����2��2����5Ε;�yd6N��-�:�r`�cHI7A�J��X�nn�iMLJц��LZ���M0nk�F@�lt�ƹq9��x )��s���9�r�*�k-��^L!�r��v w{jŢ�uq����^��hy��$ ��9(�u�l�� ��M�N۫�T�Rt�=�滭����w1����4�A0L��-ˤ�+@P��T�)N��pm�ۼ�Θ&S� 'N�]�Y�Z�%센�6F�l��<�xv�NL�P��֠�6)Ǥr�j�lj�N�^�0��)R�{��l�ےS�mˤ�y�[p�7Ḑ�ŌK�B�rf���i�ޱ)0��J��"B0�no]g\��u�ˢ	A��|ݐ����B����{��5ډ�(e!0�mt���O5���R���Vl��Y� �)>���>����}�F!������ �2��l���\��!79+׀�YOV�,����sM�.�'��@��*���a�r�L��l�j<�r��X\��X�!�-�Ր��f�v���i��u�NO.�j�\�v��k�һlk���x<7t��j�8ɗ���4��7�q��΋�k�����YM��]��I�z��5l���@�r{���p�ەLܟu��cy{�m�2��n�~�s��iF|�:ه�W	�:�)��b����kq]0ȫY2�( *J��ܹHr��U˜&��M�i#�����sWL��v��i���[���:0�wc��؊β��$u�Ğ:zk�sD�n14ۯ��� �	inM���ǯ���*��K8^f���+���MH�dŊq,�jh�"���]Lk��m{�����`�>�齃�+=�1r�m`�6�vjy�!'A�v���b�8���*g;�n�_@���\�\<^n]��:�[�����Ǿ�m��نE�[8f��b��9�GodÔdV��]6����y��ͷ��34��ݵ�v��'"]��)�;sT�P=�7�k�ׇ; � �:]3��]��Bn묫���d�F�Х�U�Ŕ�wk�����&�7]°���
2��ܔL;�{a��t��j�ݝ;���|i�~wf�/{�􄄞�E! P��	�X@R+ �$ H�@�@$+$ *@RP$� ��$X
�d�P!��I+%d+	"�T�P�))E$�"�`$ R E	+ %I$����(HE�H�I���R, P"��
 �B
I$RI�!P ��H,E��,	��J�(HBBII,�, ,��B(I$	����+$��� ��B�Ad!� , E��@P"��`H���Y ��@�A`@�**B
���BBE$!� IR@�"�	$�
@�@�*B�BV 
*I(��@$$?�xx{ʎ�����ߝ�
add����U���A�qq:ܬ6�� !�fL��*]x��@Hf��6Ǽ'ڤ&�3Gc��id�'>���>�w�4�h`����q&�˞��H­����AV�'5��5�_	w��?�&�for�ڧP�3��oJl�ם�v\�|`��d�r�}�aE�0��ˋY,}�k3�<��Ω�*�󎭥r��v�f5�o
��=է�T�d���k/�]Ρ��}��#Os�fn��wl{}� >U��0�Vj
,ܡ��F��EwR+̼�8�,&�I��訆��Ѻ�K�'��5�q����c!]'��=�<�K�|���W-r��#�z�/l�>���v�]b���S��*�9���s(��n�P�UZ�0�@]�T��$��c!�L�0I2��u;���b�#.r�l�Y�%�+Uoqܷ(k|nŢ#�Ӟ�"�qwg�aD7ը�&��x-���i�� .�n:�nɗ�E�E�����f�T��=����m��d��ˈփ��%Ԯ��;���Qv��jx8A��CE���ո��M�	�g+gp&7Zmi��n��w){�.{�w\�n]^�#���~]F���k>2?�v ��߉��mZ���Qg�W��{������P��O���Ef�@D���\��ԩ�8�WS�VTV-g���(*��ю%�W@�z��)p���o{GK��̩�/��&-��+ֽys��3�qN�'7x't�T�OK�{�uv� [��f��P������6�ypxz�s|��,v��s���F���L�'�7�����8��pg��rA�-0Oa��},u����յ����L��)׹��ݹ�Wk�Ɏ_P΅�P��y�R�]=��mU�_)���i}ۨ͆b|'L{/ ��:J�Tew6Ļ5���0����p�1�2��6as���&�(>��mv�ݱ�R>���9���3�J��	m��G�潸�k���{��,vct��*P�x�Yi�:S���i�G(5�u��/�V>�ّ�'�Dd�v��x���92�I�����#ҏF����GGt��"��W��5(5�U�<4�'z�j�%u�W�_6��e(f��m,��g��*D>F.=�>�y�fn�ZHW�����G��� �GJ[è�e4�陶mpzOd��Eu�Cj�+���yݨl�Nh��&�*����ˆw����OD=��ѡ���ڂG�YZEe��}H�5Lx�_�등u�Q�����;cWOr {���j]@�� E]�Wn��P9{�:��l0���H]!���7_<��n��l���ugB��F�� ќ%���W'k�5�n�w���G.]78
����-���@�'��n.���uqR���d��r�ꆺ����Kb�e�ޝ2�J���+�{{g�6��Ԋ�ȩ���v0i崆=��e<��I�XK��1��N���nv�D��F��`�^9�5��Ҭ��tj5K�6����Lt���c�EmGƉ�y	9�;^�"j�ʺ+� �F�t��).�u�;�u�M����8��q��=��xh��%�1@E�)����c�k��]���;(sYq���WV���v<B��$��.4'T�I��4:�q�^kͤ?���2�t�/EWf�N�����+��O��H��WT��uh`�Xr�������>B9�h1mE�R
�^�r�cz�s|�׌�yB��]�yڕ@n�;�ϻVN猓�y��XS�/�d�/]���|ɑ�����I�%Q��]��͒yU���eܳ���vs�'��پLi�x�@�0�]4��/=�z��9�}xĦ���i0�fg����u9}k+�E�����Sk�ugL����2�:D��:���u_S����.���9$;�OGh�{w�t]h�wfXU7d^�D2DT�q���,B��t�>"��k��{j^�*���r�0vŢf�rBL�׏/]�6'hmz�!�X���ow�>�7R&��3&�`Y��o'{y�*٭�a�YBY)4�^Pr\��ڲiM=�NYg+��4xvp3�r{}��t]�G�;*������>��:O//��|��/>>���g~:|���Q�`�0_d>��9�!ҖÞ��n;0���!r&��x-���1�m�m���n�cnG�Ʊ�+�L���w0Y�ŝ/�e�N�����ڹX���(�9���ʵ�c��wC�]2�ߎx���jX�k��l������v�:�{���H7Kj�+�z�8FuL a���&�{���s\�C��h���(�������IE�>2�*-pwQ�bNc=��(ӑ��u��M��"�g�`B�R�x��8���f���(�L8Ѥ�m��!��L��ׁ�J�3A_T�v�|�i�=����]�oQbd](J���{롖��R�>\n��d�UyF.s%{<����YW���ɗ-^��1$��}y���-;�0����bӯ�s�s�����K��9*�!��u2�%���E]�5�O�V���ұ��5:5�-��CK��wx��y��z,���I��Nԣ�$�np�k����4E�}h>�H��-�~��^��ż��9��L>I�[����� �Ď���W��K9��E��Mk�8w=)wk�I�yj.h�(��������9�e�:��˳�u��3U:;)�j�Z[�"���4'��W�����,�*-j毎�D`�͉�d�P��KXCF�XX�E��Iè�f������f�.�<֊���f��(����p*ۇ9ԃ�M��c��u��Xz�c�u;�q�k�)�%�H�V/f�=�q<��h���ep
�J�<��{X�էg�6g?����z:2�y�� 4�����Q��na�0��Թ��%N����P[6�i���-_F.Xu���B�U�ӏZB�񼶗;��yړ����AA:����g�wm������r&8�Uw�����NX�#�b�ccm�q�H���&��kXîڹuq�q)S���9���aJgD�x&+.�K�k*K����G��q2)�/�B-N�jP�,Ĭp>'��؆e.��]]W���}տ<0U���#��;b�d�p�o.�w4��7E�}}���bɦI�,��V�}!��.�.�'I��������i��x�sjc=�S�TJQ�M�@�; ���K��r��GFU��̍㕗D��S�<�c��VM>C.���X���L{���Z��Ʋ:�B%��|�}+ҳ�����Oc��«=��iNx,�{$��Н��40��Z����O`)(=mr���{$lS�b3ϼ�O���[#���_�=��(����]k�r�� �t;��pm�u�I���yEn|xN�i[=������M^<}<����e�{�JKL�k�k-��b���}lL;՜ȸ�(�,���*��f��9�]gb�=�2I���=�2�,&|�^���u�{�Zr#{c5�>xP/�^dX�16���V���N�)TW���^*��ow`�B��y�ܱ(�>)�](r. ��ù�� �U|V��mK݋<�f�T+��0�^'���/|�D+�
��
@���2���׍�^��I�&'wǹ�ה-�K9�ϯ]H��*a�E(r�Ae���xn�|X].�����S��ĵ�j������"c�.�W�+����2�l�/�y]����ܨ���;.��h��B�q漴��҈���V��ys��0�묾��]ݔ���ÕH���s�09���{g����=�,>z�=�C��yk@�1�x&R�9��ْeԇ�]۶/�������n �
��`�xf��Jo"�9�	úEУ��#�$����Ɖ��m��'����Gwy�i�m�+�t�PۭBiv�[����u�ݵj��K�{�P9�>�g�vR9���gK�U!Q�+΃&���rO{�����t���C�z3�~�ל�^5�3(CHݠ5ڧr�9We8lN�̰zS��"�!+�\c�7��S����vPF���Vp�ZT�@�n���q�L=�o|�wX�Y�w�}\DLY!�SY�⮻R��4�#Ӂ�=2�'��A��\��Ҳy�u=��úmB]��>��bZ�|57�I�?+�� �eΙ��G���M�矖��7�d���o�w�­�y���Lxseep��W�z�`�P�tL�b�ީ+��[�	űaO��j�.�\��Z�"���̪].���J��B{miLG[�G=}����}�g��T:Ռ]V�OS��Q����1��ؗEHgH���kZ��������H���`���ڪr��l�1�x[�,�a7+�T85`���=���R�Q�-�_y�~��f@Z ��e3�f�d�Z>D��;��.ɝp�]W���0�sUdz7x��3��#噐k��R�Tw�׷Hwu�?��DzfM=k6�w}�{z���"�#hlYN�')�TC���R6'�Lb��(����֐�t��f؎�m��|���^^μ�D�k��^������B��C$%���4F��Vt���SX���n�|���v����u��2�G������J��ƌ�1�D;�ʬ�K�ÇR��Yv����W۬4���Ƥ9m���Io:���e�2(�ݳ*t*��E�/-���Jb��B���pΜ{����&ߋ��ˬ�p�Y�M���vS���q6\�h�;��[�+d�;�5��=ޏ��/��X�����i���
q�]Am_<��gdŚR_|=|��x�׌pz�\gڱe�f<��b9�IBǋls斶�-}FM��.:핶x�����Hv���2�\���(�".�`�N4'B�f$VM�j����z��(�5g�9c�!�s�U1�� �(��v>���9�{@Ǎ>���T.+�u&ov<�k6�9��7͢�z��hΛ=6�>�*q��n^�N�k��R�ZRˊ���yO����_�t��Ip��q��u���]������?��� ӝ��9 ��}0ٚ#ܰ��.����e\�vfKRe�&���F��g`����&�}�x5�3�����\&���|�6-�م���|�^�7">�sr�h����#xs��Y�<t���YȜv�f�롬H�!����x���v�d�����nvR��z�>)t��U�i�v�����E5x_T�<��G8T;�)�-����hU�P�PX}�}�7�9�C��x�ȯT9�q��\pѼ˄��0��j�h���AHbg$l�#��&�n7v�f�c�x[T-����(�F�Kڶj��N��t�FQOk�!��L�x�=7|0T=~bU�4��yb��`o"�����i��^�}��T��=�������5������I�w�=d��<�*�K�f����S67�{�;L����� ������^�cp�l�ӊo��̛�O�
u�.�.Y�ב�YhW	U���n��M��>��7�WLΙ[�FM\�:���ʦ�{��_(1���G����ew!�{�G�Q8v�.b�R�iu�U��O[Nd�.�0��5�0��MF��1�ŷb�lƂN��eL �㾁[ō�;s�[��˱�n�-�F��qu`��(46k�bJ\��:�J�VZt5�靼Fbhn�&�?3D^3�����;��t`_[�t�K^�RI�ӣW�a��U�w��W�������.Y��I�E#�||�)�J&�l룦�x�~��y��6bW�u��T~"��=I�б3�=:ݼ��97��v�xu��̎�:�#�G�5q�C��p�����w9�ȗ%9Hd�Ss��I�I�ua�x7�I�(ll+a�_$8��<7n���!5�����S� ������6�3�[�>�c����|��خ
]�s��P3c��ut�[�A��]\�.�W�t�D.'���7R�p@��J��0"u��NkAo��x����D5��xJ�mL��Q��W��\FM�Յw�V*��)��c����d�����@P�]�u�K��X�Yٯ�?Y��V����t���Yof��IJ�@�ٚ㫕�{����8'�Id^�w;}��l_�C���^k�p�Y,�T���*����/j�:<fcq��8�<Y��ZqT75r��7)[��Ǹ��
�J�Ȼm.�^�K����4���j��g:���V������Mv8�o,�P�Z���x�r�`���쪅��C�(p@���Fϴl����S�f���	5mr����A,�ӴFX���Aن���ظo&Աڰ�$Т~T����\Haj���˗�>59�u��
2KѼ�=�;�Xz�_y'h�z���F�yh�_G,�ٛ�g_c�nB��V�"��y�f�Y�j��⮢jd#��c�[�Fw$b��g_ν�E;�fZf9gf6�󧖎3��D�zeM��t�W��h�h���ʧ+����Uc��hff.��)���<QP��t�f����m�'�Pnmj/o��r�t$�if����Z���t���w|^S�c�c�c�q^<V��H�E幟]������e�תIz<��RՊ�T��g�������-`D9W2ۧ���1�̈́T��%�����^�����n@�r��[�[~��ay�}3)�z��ڡ���5�eG��u�<��ݗ���9�[Y"N�R����2�u����{7j���9%~�=*n��3q���-Fz��e;;j�*\��aͼ9,�M��1�Vb�D�+Tv��O�	k��C��V��2�6�s�+�
]�]n�E;6Fr^�}0�nVռ�U)F_�UW�|@�p�I���9��t:u�]Zږްj�]D��Snxy��kn͌X�̈́�Vy׌a3��lݺ��cnz����c�Pkn�2���7pu�2\�ڳ�N�l�c���I����&�+,i��v�#v�w���-��$[�74q�}OY�)�4�Y늷iq��Vۇ�o*�oG�`;q��	�@��y�6ٺ�t�(
oV-�n.�y�.�7e�^��v蓱pU�����yD��g>`�`��#��q����U{��t�8h�;z뮶�n�#�ۭ�̰9跮���XU�`$C�mfMy[��l�E��i�sյ��Z�6����m�n�`��I�.W�:�R��v�䱛�:�ڵ�\�����8룮 �^:[+���v�ۥ����n5teSc���x��x�6ǳ)�����
��V��ۻ7F[�n����N�8��N��"�gs��y؜]\r��ܵ�{g���e;�\�c<9l.n�k�������j�p��/��^/=��g��=��r�=o<�%�vcT�Ony�rnz���Y{b瑝�=^uvs�v��s��An��K�%��{\����!B�:75�k9���^x��nݶ�S�p��n����Σ�3�ΰ;�ړ��������Zމ�t�uP��]��6Ȩx��9�{ �e��;������������\yL]���E���Ť��'��b�[��O8	�XŹ�q%�;s��m�ڣ玉����'�Ѷ�P�״WŃ����&
{i_G\��s�m�u�=��M�����k��cz'��!����[��#j��S�uqF���q��Z ���gp�p��rΝ�й4k4n����=�X�q�@���t�&�v�ӎ��A��\�8�"�pL]��#;RAs�u¯9�HYxz�w%�� ��s=;aRY�ևm�ɹ�����-#�]��k��VvI���wY���M{b]⃱�N	��^;TS�j穹wv14��V�X�gj�y�]�J�Z��\@�y#��qE�"띬�vx�K^�;��LUծ�sg�5�7oe�[r�F�^�#����qB�a�%���٠|+�piۧ<u�s�����m����[^�ǱҝJ���;e<򝺶�p�%Yy{=a�Ŏ��ܲ�Δ�9���	��m�OV�	�.�ָ����Ys����W���kF�m�|m[�0a=�ׯ��Y�M!��VS��(�.�l����k��:�+<�k�2��t/���L����n{f�p�C��4ú���˻l���#�"{��D�lt�Ut�]'L3�Ϲ�� ��g�êxޱ,����Q��Mس����cv;<c+�NՍ�o8d6蹝=��:��:�>��`|�z����`9Քzw=��'g��v����vqs�������Uk6�u�eɭ������y��2��`��v�1��`k3��]�v:�k��l��eݷk��s��8���3�{�;rtk��s�l��ּEӦb�(ǲݹ����:Ӷ��t�V6s�d�\����l\NOo=������,��ӭ3�.��y�=��9�����3G5�qҋ%����IcscX��7�y�+Уu
��W�痡��ynwP8x����]���g1� ��]g��v�zn�z㎰����͖��;���Nm�ב�y3�y�싶g�:���A�Z�BN�8��z-��8����9z8K�����:α���ks�ѭ��K�ь�p5[�\񸷧`n�Nj��VGs۰�Z5�Dۮ�)'�sz����q��dW6�6�qʮ�����n9F�`�Zy+nC���6�l0�ٙ:������"׵�ѽvc9���Ic�8�klv����:^�q����M��j�|��E�]<�Y�r��s��%�N8���l�x�&���7p1\Z��o([D�[w�F^OEm��pz�Ӵ��'�t�Ikf�J�r��[`�H�vw9�e	U�M;�W=��!�܋Y�m�mp�M��b��������[��a<�^Ľ̺9�N��w�Z2���L�3ދ�%��!�];�ɍ�nm�։�ns��\mt<����dn��=���5rZ��jË��kG.�;=v.�mӵ�.^s�uv�t�[�)Ӌlٳ�.���ۡ��Z0�ce	]�w:t;{�v�WnU8�s�*�;�y_u� ��ݵ���-���f��\ݷ&���jT)d-�;��ǲ�m�lO&���^0�۸��,"����GY�3�u�;qwU�leu��m\s�۲���{8�i<��h��@�˶p�4���clx��v�r��YѯL�	S�x[$��.B�&��8�q��m�n���XH����v��6q�U��N�T�����{Z+nk�vt�R�ݒz��>5Wn#ca�z{��ۮ��-��6v�OGf�lϬ\��V
3�p��$�jٶ�q�y���[���0�윘���ީ���.��.�M2�����$��TH��ۀc$�;0CCSRoT�3جx^sϞ���ָoZg�m�����[�ROG`�h�l�tn���nr�l���_7nO\pu��7FN����LK��ͷ>�v=ڤ���G\�!ɍ۳���e�5[���NLtFls��1�Z=�rY�����^�Cşn�+{g���/=�byK�X��Nȼ�Rܶd{Z��ED��g`��ܧWn�ȯj'i�ز�:5^{$�ml�^]� �s�<z6��qb�n��a9�G.M�r�����i�s����kq�m��:��=[�rϞ�Q�mh�ڶ�m5�g�.����Q��up�vrK�0JCw3u�w]9kN�Bv�n�<��c��;$�&�n�vݷeâ�ts�Y엦�q�wg<��m��q����j�.��}"A��G�3����Z��r�,�*�Ɇ�N,�C�Ft���Q��y��е�[+l�޻oWbz�ll�ٌfR����x^8p���I���!�w���uhܢ�ɶ
��۞ݵ���<�q�^:�t�l<��S�7O6��3��6���n1�h��츟� sc�����]�=n�7a�]�҈S�g�c���yK
<�l%���ݢB�����.Kƭ��m�Av'�ɗC� g=�C�z��N����ƛ9�Ϸf��AK�r��	]b,E���ع� ;s�v���x��t�W��-'k9,&�{�M����&�r5r�p.���nu�!��콎7U��s˯m�յ�/Q&�q�{le�q�[g��y��5ܩ�y��m��3�1/�2���]�5j�kev�����x�.����;1x�XL�[����u�n�`�'�n��1�u*�=��ӉMͺ���u��M��w#�Z�z�n���E�x��\p�����{;�.ۉѝ���1�4�� #��9x4�r1��֭��rpv-['n���T8�dٛ&�v��pp���ᮜp�WQ�����ˋ<rw�9��@X���۝��[=��y������glV�����C��ɣ�:�Ck�n-����M��l���c��������]�/h`�;��\ku�vh���Q�M�;��0b��ݦ8��I3=m
���sK��;�������b�\����wd�����펃���� ظ�w[v�]h��R���]>Y���-��<c�ݱX�8�JJ<�n<���@�-���<I�n�i3�Y�B�{v��q�9�Wz��z��=�����=��z�cpt.Wf��_lO]8�v�nr�l]D�,'�V�{+���^	�*M�ט�a�hv�P�:\�+ѧݺ� ��/;;n۴�F�Ԡx�v�ƺ�xd^ǰ�̼zx&�M�w�;��G[�»9wV��Go����\��=rl�&˞�b�;N:�u� vǐ��ݻ���lX)D{zն냝��u�15��*�]�`g���i.�avo��}m��őΓm��`��g\�����ۃku�w��Y\igv�۝����AĜWV�޵*[r����{v���ݸ�"���)7<��¢���GrlVK2<N6\l=�8|�#�y��\K����gN�]��έ�)����&��˶�c���ݺ��F�ݵ��Aqn�n:��������)�������n08뱝�{g�}���s�1�2�{n�k��woop��8K]���ے-r���FGm0�M�aA��������x�ۭ����=U�ͺ6��{��닭�G`n8�/W�����9���7��[�iՇ��;q�
���\���+5���f���ڳ���v勭ccqH<�0�q�=z$�;pmh�oc�S����dI��o)�۳��ڸ'�\[WYX�R}`r϶��mq�5�����z�v.w;�g�wmb9;l�'�.ɰځ���CQh�v+����M�;%�c��#��rmj�M���N�&���Qvܣ��0�l��O����u��퍺�l�k�ۍ���v�vo�����ò��v%�x���"���D;0K��U�㇁5�Ҿj���T�t���F����[�ɱ�p��.���笼M�D��4�Ef�^�u7�q��^x�&v
�g�K��r6��ֶ���׃ɫ���-�nL�v�P�a�G [�����!bL	�l^��Lv�cV���ksi�q�:�
V�ܱ������%�웗�c���C:5�3�X�yS��F�5^|�y�Q��.�����tm҅�r95I�8�{vٰ)׌޵7Sm���-��g)�v���;����A;[�tk8���:�{y9ր9�glǞw8���(���;l�ڷd�4��x�n��rۗ��W`.�`�yzT�ʹ]�����#x�4ν���٘饭���Es�k\QE�ţs*u��k�nLV��=;nguƸ��\��Vvu!��M��=r���j�9�~waTG�f5�)Z���4�������IV�JQ ��UHZ�-��R���c2�R�ʭY*RѶ����AL����j�\b����[1�q�-�A*-���V�Tm�J�DiJ���V�`�TiW0��+Z�*"��DX����Ѫ����Kl�5F։H��T�֌R�c�\U�-�"T��kmY*�V����ڠ�3-L������U��-KQ��m�����DQLI�%�R�Eh+J�chUUb�m��"ڶ��)��a[j2�-ƖэF�QQ�R�֥kQR��R�(��-�-�KRع�ceZ%e���*IYTJ#��b�6QR�kbڦ$�2�U�[[F�m��%B��EJ�cQ)iab,Z�R����W0�pY��*���ZZ�e�,j"�`��*�D�1��m(,���m�ҙ�1f#)cZD��jV���؋���-�E��KVT�-Z�*[cEnU�Z�k�f[��*��$�;�o�V[�qզ�]f�Q
��n�6���ݺ�;��?;O��v/n�8!�q�#�%�������r� 7�%��\=���v8�u]<�Y�^�����[ccU�.N��ڭ���F�kmR�pq��Px��vmu��^p�����{wO݃�7/]n{[v�+!�a���-��#���+�KóӇ��6�GF�.�!���c�v$��l����Z�v�����֒艗�s��1�dM�ǋ6S���*X�Ϻ4��'c���&�2�|�'B17�.�ہ룎J�����w	�u9�m��\���វ����l�#����5�l¢nNnǺT���oA�v��m��˓�C���ۗb��w:���ݭ��)a:{X��\x�	��e��]sW����X�1�Wd�p��I�����o���|�.�=<u�ӌ�`���U�q����Qs�tm<P�a��=n-
�,\�<&�Z�x����g��Jh�Fϧ����K�� 瘺}�.���s�>7|�6�G>g�ʦ��oCmT��vy57av8��-ɉ5\��1��e9��x��F�9�9���mq���lg�à���P�l�o[��=;m��t�;y��]b[r�N��6y�i�v0]��r��t�����@n�[Y��7���9���<|�����m=�Xq�SkV��gA�n�h�윏k2���Zf����ܦ+h��<Kۉ9���$��s��O����I4g-��)��X��'i��m8����\�*����jDԑ�W�Ȧ���S���r�덻Y��͍X�秷kq�h9�sq��.y7�f7n9�p�@�9	)8)w���6��|qv!��%����c�(b�9�\���p���v��cے�[p�3��7d���l`�B�m��+&8����n�b@5on��n�ǡ��ʔb�v/cF��v���^������am�z�v}W#n���M��g��H�W\�)�0�W.Z���%�-�j5�ŵ��1Ÿ�Xd}���v�d3�a��'��R���UT�m�Lr�ZXa��eK��%��s�\��P��9���^�݁�|us˘��.!�n��ہE-Q���2cF�3�Q[��/
a�.ώ_+�ʠ<�^˰>��\��c����.}�)��.G�AT�=�B �V}���pK`�e���'.��,>]�� Sz�-��튓���R�~�4 ��'Z�����x)��`:����CD���,�s9����n���X �~��@[w��x%34�6ػ�@�l\�ZBٙO�� ˓����IM ���o=�u;k�t�ޞ� �:�� V��q�"(�pS�1' Z��*���i��˪��	*�>��[� ����Cw鳷����ߢ���#N\I*%9���z�Z@|���j�F�J�%pfLJ��:����߂"/7���f��~��dۏB�bnF2[q?;�U�����YL�I�z��nq�Kۃ��ʑ������L���e�4��r�M ��~� 	s�Ͳ|��^�s������@��r�k����L!�����컱i ���|�]ƦL��V=�S���d0��d�w6?�-��{u���y�`6�z�E����������'��<��d4gº�De[)V�˷D�oW�h� ��� 
��V<�LN++ڦs;�)/M�Pa��1������ A���v ���9���Og;��c~ ���V�ft��"jyE�{.f]�]tش\�"�|�����w` ���Tɐ�6�㲤�I{c�B��>�Á Jd9r���w]E�ov�u9_G{l����d 4�N��d�?��R$���@�EF�ę8�ɂq,�F�5�ˋ�nv�'3�4u��5s�\$�Sߟ��ߺr�Ĩ��29r����Y۵j� �-����,��AzLZ�-�y��=�D�n��`����f�$m�(=�[I������r�� {�ۢ@߸��z���7�<����']�6�T���%���˻�@ �}�� }��Zת�Ӯ�z7�Y��H�s���v�W.o:䥽]����r�Xæ��u"��)�d-���˚�ǡ���qo����}D���ۨ� ˞ҕ�o�p�����0W�GFF��K<M7��A�I����X�n=���}8̇w�z���V�m zk:�-T��B��n�_êA��i:0׏�æ�P��^��,�뻿�"7iT@�V�q�Aӻ��w�>y���X}9�DdOQq���zj���6B���Z�{V������k=!8�����޻� �7�: +}8ȉu��Y��".���Y�#2wJ�\D�7��Q)�TQ�/_� WP{�r���y�E &w���%߲YI���޿wu�a��:�S0�\6��b�M�X�2&BNwCo��g)�ݰ�Ҩ�}8ȏz��Zr��� ���=��gggt����z@e=�N��K�N3����s�.����5��RU-=&�C��{�D�O����n�.�S�vo�/L�G�U�?O��P]���v�n�_k��x�^n<��MΪ�4:�AA�m�A��]�!��o{jՍ���t��qc�~�eMQT�H�{���_ Vwmڲ'���}>�������9�Gg.�3��qx�ZKF֮�7���3���뎽9R�>�>���m�.�g�����i�@�0ܟ)  ��ۻ�*�o�͗z�"�j�T@�1�K������5,%��ʨ������´�:���j]�
�<{^��f����wu���w��E�Ni ԧ1 �ɤ�=pI&��+E�D�K�&=9�ϸ 7�߂ Ef���a��8��b�*�JT���_u��łB"9���"����1�k��;��x�#@�{����6�R�	�	p��uX� /����]*�Eǚ��$�ov��dc�����𥳐Bts�cč��~�9�<{R��sS���p�a���R�J�����W�^;��8�5�^�ʑ��1�U���Y�vep�2[���������PLW�v�˷�d�+��S��Gn5ˏs� �n::{s�}��}�ls�a��l�Jp�m�n�:z��É�������y��9��>6�Ό1��[W�끇��^Nl���]��Q��k����]{o��e2���"}Mom��\�5t:5\��mln�x�C��ط>:����6��W���n�ڰ+x �.@���	�\qv��Lx�\�p��&gu=N�r�2u�f���߿~�:�H������� 6���X$�}��]R=�ԫ3{�\�m�cz;sv�.�Ƕ"!4?�r�R3���-�����[�t�r ���v�J�U��oi���}<� )���5,&bk˜�]I�;��H$��]���þ�7n��}�o�A$і�֑?x��,��4Y	�.���(Y����� ov�Z��+�����o���'����$�ʪۣ;�"��bn�j�~�>��&�ۜ�P���^<�N�l_<Wu�A%��v�Y�X�����z�ZaDP����e�A�Ƕ1�FF'��熸�nz;RЉ�˴�������.��܄�Y��v]ڰ@��_ ��'_����]�:��� @|c����z�m�4�?� ��t}�+yTeس���8����\��bqz|�./8L�x�]��؅S>�M١��f]mjT�V��esݬ�� �>�]��"o�����:^�X�yyW�����*tD��EW��vҚ A������"v*�ܸ���X��#J�uD����)ݖ�	3�6(ׂ�=�uC��I���bs�A������<+����-�n::`��~�t�,��$�Թa2�+�:�y ��j���[��7���i��������v��tFҳ�9�b�!� �CL��8�K���{R���k��si��1]�H��1������L�Cp�XE�=YSQ����!��7���@�=10l�V���}���������J�$Cr�U#��w+ ͽ���W��7q����� �����n�-����[���N��^�ޱ�S̶ӈ���� �m�mX�JK��Y����d�!Dd��"�5ϻr*�����������n�i��m����lW>,��>�8d���;��\��HQ����+�Q �v�ޠ ���ۿ����P�4509��Qod�^t4NWE����fv��_�#]��[��ʞU��\R[��&E���8A2`D6(���M���}�[������y��� ��۵d k��J�z"��d������<L�a.u6���ٳ��dns�qs7'`M;�m�J��q�ot`Ԧ��%���S:�� �*{�6I$�]o�i6M��1���"lϱ����AۻV���^L)x1!��E7�a��$�>�(���a��@ fn��_�|�u��>	Z�5��Ol�}.��JJ{��Æ��!.D�]V}` i]�4 eMY�����kFǷ-��:�?��h ����Pa��� �4�.:4m�k//d�,@$W�W`�+��� [��fgMq�{
k{�t�3#9�*Dd|���>��3������h{;����q��K�B<���,�v�!S�^�.���K��β�
o�����$�d��Ob�	���5�njSQ-��cv�LS�s�� >�ʻ� ��o^�����li1;/���E�.��;z<�E�n*��Y��l��k�;���������������Nd��lI��s�ۻK�$�����K��|�sF�J�^_��V]�$��UIpOuBM���hQ��|�:�{���i詽��D�v��T�/�ǀAK;#��OO�,g2��OY��ʯ�*I$���J$� c닥���^��t  ��=T��'�[�!	9/�+��L�SM#�>۪"���r}��9x�v�Y�@ B��`�H�[��쨅9k��[�iUKf�?dm8��$k���7s��6b����̓f�	LϨ� n��<�{�u��yU���
�p�v�Sl��/'.cħ֪DPڑ�b51��݇؋��=�^u�p��S �;��� ĩ<>Y�@�74Z]��un�7o�"~-�`(	�2aR�F��Y�;]=�ssg'mi ��du�����n0��{k��<q3�gGn6o>�n܂�����g^$`}\qI��Q&���k^V��9�x0�����$���f=�����(�9Ӡ���T��,n-�Czɶ��ێ���s]\��s���!���Ν�N݋/Y.7V��	{0�Nj#4���v��	F�s����8�A3b{���a�n�W>x��q��q+;ȱ�.�v�[w������ۓW9f5�k�� 0ܗ�D
��n���yc�ݯlG�9� �li'-�I�Ʉ[b�ڞ�K�W�����/Ǯ)V� �.d��~)��� E{�-tp��w�ԛ����m�٨��:z�� ��ڻ '苟w�r���>�ӌ��Wݷj�v�&LOYL��~���� ij(� ���ګ ���=���$�B&@��6�a�F8qU)�˻�|�6�t<��W����^��@%����"�:��Y�y�*��A�6�`uܬ�Ȉ�(����^m���%���^̡��s�e�e�l;�_l{U�����w����\�r06�H {�U� YӚUJ��Kv�V�cwm�@��ݷQj�ǵB�L�Z&� �}����W��^�V��bCQJ�ʵ��h=�vy��R�R��(��q�Oy�����B\�0
ٞ7���Ws�T�!�z`�;�
{fEM�n�/%�v]�Uq�i 3;n�Dg<ҕ�T��ՙw�Ih}�؄Y,��8h�=�b��u��t ���X��o�����ۻD���M
K�zv
l6˃F�2��n*��.]�{YU�����P ����t*o�	�芽����{�''/ǚ8��4�k��D�����ھ��s�V�]�� ��إDa�߃bf�t�����xߝIF�;OZ<�i���g79c�*�����(��G'x{��2M4�P���X �����������tI�vni\ ���Z($sq�R^u�n ��̲MQ��~�_娟V=덭Mum^��r� �=�T�+o�� Xo7�P���,�Y�Y5�ir�Aa�̢j�P `n?) yVw��W�}�'�	�3p:n�"�s-n�u�����G&�NΏ8ܕ`��[:����y��Zڶ�\boU�ۚ��ځ���!�)��i�Uк��!=3M�u�}��%��ڞ�姖)[Ҝܷguܛ�]��owۄ��&�}�8Nk\�W�>�/��8.c�Ft��T[��)դ4�[���ܠ���|�v�����������Ʃ��� �l�`}�����XE4Y�cx���A�YF�
�2�6�. y�{j�Wz�dYW��֖]�O�\V�)�u��^�:��H��i�9c�_3^o��76��Ҽ���o4"|\\6&jA��܆��At��|��Ogts�l�"����S��]o�z0�I�&Z O������H��v�ގ����X���.�ޔ�%;���p�xu�w̭N���,Z������S��Ǯ,��o�.��zl���.��F/�X��q��K����b�;V��W���bk1�7D�[�� ﻾EZ�I�+|iL{i�ۂ�p��&gV'+�,����N�PA��;YF57dg��|��)�E�3;�˜ 8b�V���BZ�WV���)���T��w�,Ft�?6Όx��֎e^�tf�{�Q������w9:�:�N�{{�xW���N-�:�:�j-s��X�Y�;�ϱYם�W7N7z�i���v��)���|f�W�̳�J97@˃}\��ݭ����R�{�nnN�f�qB�;�*g��<=�x>Cr��e^�A�lҽ�A&o�M�F���r+�x�ދJؕ����#~߄�0YK*�e����UX"E���K�kT��ֵ�Z�ʣ)khX��*"�Z�h�)Uk+Эcspb�m�YAkZ�-UQF��iZff)jV5,�ѵ*�,��X�)m
ڭ6�%FѫH�(��6�J"�Jն�qƍ��E)IQ���AAekUĹeTm�ˆQmh�إF��TF�aB��h����V�-�F�(�ER��j�iV%���m���B�eF �AV�4)KR�،(1iQm�[J��6������5"��m�����F�*ƔRҵj5%Tj�hZ*(���*R�me��+Q��lm��JX�lR��(��*��e+-TZ��)P�*[m��e�%j����*��R�D�(UV�Q��VUJ�2�mmeU"5���5%J��UeF�h�J��-h6����m�ղ��QT���#JR�҉mD���4��J��E-��E����D��,A���-E�)R�Ij�Q)hTmZգJ��j+jZ[m�TE�ն�{�7�e�R3s�D }m�7��9�2�$�26�im�u�H�*;�ya$�>wAQ(�������{o3�es������|����"z9ĹCQ32�TQ�V��U��T{�v6����H皪� ��7��{�w���wuUIY�����}���)���ݺn�.��o[�<K�魮�'��s����ȓ�>��e�a"6�>�z�i�@ ��~R |^���n���K�;x���?q����o������.Hc�-��#��wj�7�]Pͻ�[�WΏ�Ho1�  E_vݫ A�����y/8ߨ��[NI�e9q
&�#�� �A���X �^D����)GztȎ@ky��� *���Z^�*tA�Â!��PKz;^�ڽ^�����xo� ��i�A ^����g�quW���>������S��x({�����^��,�P]T�ҋ�gI9�oc�Vkܰ�1�W�{z��]ַl�%d��Kb:�%%�s�)�8�ۑTW�_��Հ �y��ZUU����AS%  *�������|���J	p�AG����,s��)OWF:�ۛtkb�tŞkug���0�-vI��͇��73$��rG�<~`�
��H:$�I��րw�ݺI�r�+y[��x"�}ݷiY�/\�5. d�@Ҩ�)r�G�_���* ��n̺~a�]۷w�D>�t������"�~��e���R�7$1˗
���7L�$�<}:�K���~��	���"N���I�ّ'}bn4�؇��GFG�d��L�p���K���š ��u@+o���몛ܽٿJ {�wv>=�(jT�NeT��Υ4|��臘�+�V��N$�ޮ븋Hc��J�����D���5x���v+���aC�,ڋ��"�m	�Ğ:��%�٪�6�����!��%���=CW'}�ǣ/�^�mlŸbw��N{�{��3u�qg��mn8�i��4Nw�Z6�����{U��v�۬�)�;\x�ce�巷=�Mi{`�8# ݭ����k]{HG��u]���.���S�qqh��B��c���tn�-��7:�29�g	�jm��lt�+/8���C�^4m�>v��-�5�2wo=�h��lX��wiwb��4�&j���X.�t��v��.�|-�s��.��zwu��4��vy�NN�k[=�q����F��ߝ�����l�)��/��Q ��wjh@ ��o�'�7�>Z�&'����˿��n��Pq�ىr�j\�ۨ���V�)�gz�d�����o~�έ�H"ϳ]DP�cq�z��n`C����\�SR���*(=N��� ��~��Ց�s�N۾��A#6sJT@����o�}�J�ܐ�3-�T{;.�<�OZn�sޯ�7�ߒ�E_v��f0�p�a�C��)P)�^����%9��Tc;� 6���5�i�ZإRDJ}>�)m�7� ��۴�X�^��]\c��6'�."E����]�`h(U\�k�����>�y���?����h��p�e9���=H ��~�@i?{�xG�%[{F\4}��T�47�ߒ.S�����$U�=���&�
G�y�x+5���{w�7vKש�8��$I�IX��c�]��z~��Y6g(�!�x����"�`��yk|��Ǹ��Z���O��%z��~N���~� *����$c�G,t=���[Ij,g6�F�,uy���DEgnUF����m�gU��� +o1� Wݷj��Ӥ����ġQA�u�UU~���g�R�� �*�{n�&��y��ى0P�\ M���rO$�E6�Yi��wv  �y��Y����Q&\D�۽$�HO��d�D��:3ȏin��~�R�Pv�YKF8{\K�Qa��Qh���-Gb�*!@b ��[>���a�!�Aw�k7� o{jՇ�s�=K�^\e޾�^�h�3wv��.|o�(`�0�6��Z���$��	�Sӗ�=`N�� @e��ݤ��}��� �$&�a\��g/s72 ���e��A���)y�y�d�'�a���D��G�r{Vg ���5���;�P��u�%E���x�����FX���=� `�8/i��3�w(s��hd�&�^՚�Be,��{���tE{�$�߻��P|��k�:"V��̶��c�RG�Z�TY�n�ӵ�u�A��uQ`-}����mU�F��<<�����75ϓp`&IP�R&T��t�'���<�dHw��{^m�'�$q���E ��߃7wiHW��zDd6���۞:��]ɻnH�K������;a��(�Z���yۭ�i���2Kk9��v�#�ͩ�@�����lV"�o)C�y�z��V�����5�k�@�mzۉ��LD2Itq*��$(��ebK��V,�%ϯ]R n��|�I삥�^�/2y�իs�iB��19�MPq۴���龜�g�&v}n�"�mXm��Em�7����f�D/6�Ah-���2ɽ�H3W�v|�AgU�R�[�o�+���t�e�諉�w�B�w7�D�:�4]��v]n�g�ܷ�,z��j;n��ջ��u3�����BG�du�
�z)k �$O���IlV}I�z:b\�$I#��N� �+����*Lt}6���܇=�/�	UwZU�|߀@��wfU[��틙�m9���9��!�ƺ��2��i��Au�t�����E�p�����ˆ����J�Ue%4F�q���w`S����q�9׹Ң",/��޲fnHc�%�T��˺���3�7<z{T��n"#�vvݫ @�O�{��nm�T
v׭��.��DD�pV���7s��"-k�S*�1M���s��>��b	����ڱjܬ�A��f��rN��(��������@�{v�� �}��DDU(���F Лo��y-�d!���C�n������-�X���ŕ�HI�w=w�H����ꬁ�]/����t��W����bI��"jߚ�ƥ��;d3�Q�<1{�{zOs�@����˛[�\�+�!����MT�QZ�y��/!����(��E�㷩��ɱ�h;l�V�@.j�t�y+t�2x�R����;qc�NwF�67Y�:�Jvv�g\y(:����=�[pjm�P�ն�u����s���3�nƍ5�H�y�u�!םV�Q��v�\��l�B�똷`�����ÍK����&�aݟ]�|u˝�<�]w=aő�h�v��6�����hθ�,���!��{9���S��ӴR�R�V��uŧu��Y��'��k<��u�	���q�� ��0���'�'̈���ڵ`�;5��wF���;�R����"���J���&"
a��i4�뎀�s�b�嗈�3T` {�w`�]Q����\/nf�v����L�M���%�T�;�wiX Nͥ4�J�똟3ʧk.[��".�Y �ٮ��S��D�p�P%�yd+��y�9�-��S7{V���>�u@$ͽ���]]r�W����]�as�B��19�MW��v�R�����|©��o�n� �F>�t���-�����L-�gq��~|���w���y�;G��X����a��b�I��v��mvH6��r���k���&�n �G㮷n� כI: �n��$�o��V���9�>�� @|v�i_PG)�$�#D�QQH�m�}$Fx\>����ӓ�v-+���'k+=j��Y��t�{�����9y��o���s�
O�nĻ�h����`����_%��߫�����@����O�N���n��3�"
�D�s-��@�N�� �� zjUeN�$��7;����U >�����3�,��r�mU"s��+��[{�;��|�@�ۆ���	O��GY�yڂ_NZ0$���T)'�&�%@`�T���!$[{�V-v3l���ɩ	'���H���� ���^Mk�ȹ�o&���z#$A.%nܷ��M����al�8�6��]���ncd�-�Jۿ�ߧ��܆LNe\϶�uAz8��*����[�Fb6��Nj����-�`LS3-¨����]� �z���k���t���΄�z? +s���Y�eHfo�j��]�H54ඤp�����yH ��wj��n��HʖR�.�U5����L�no��R�oTU��r���AZٵg��a�o!������E�y�0�k˩j��2#b��<�3��|��K�|? _����{�zfX�E�dEN���9�w^��H"��� e�mU�@#zoN���kͩ�S�HG����Č,!�%��H�ܻ���7��:؉^�V�vOJ���<? �ݵQ��ޔ������Y���1�y��^o5�����n��R�]��I>ܙ�Q7��l��Dm^��\8,��^r�Ǥ��� �����n+#g��#�Ay�W���>2�&9LNeU�o=�t X�{}7�x�!�}��v�w��"-^:���wn�-[�uҢ�N���
�pH�At�uڰ 3]�'Q���j{\oFOP� >}�wdD	�zWʃ��;�KA0����a{K��恓-���l�|;WV�s�=H����u�<�q�bu�����y���!ր���>�b�'�=˜�K�h^:KWV`�������r:{f��x/8t�Eq�wߪ����Q&���4y<��D"��D
@�O�I�w��������n�<U�]�H${��W�U��PMH��ӂP����!8.d�		��&
��Zںa��c]Oi�t�����w���lH�r��[U������o;���'�O���%��Q?_K��qw�d #�oJ�uڶD�q0J��Q��6���nwnu���6�&�$��>)Q m�� Xz{k�3�>`�|m(pCnT53*&�;��:�^��C��G��:L{�{h�3f��i$-E�c�kn��`�9�}�q��U|��*��'G�$�` OD��,Vz�8<`?hǏ�E:�ԛ�M4 �d���m�i���ڢ�lW�&C�9�|z��8w�� ���ۻS�
�R\I
g�*d�fb��}�H�f��Ie(�3.p��N��t�y�Q���A�S�_��W޼�}��5��%V���zi�?;�@t���Zjʹؠ���PA`ʑb$`���+�TF�o����t���{!��n��qutK���m;�\�8MK���+-�8�Fa��uTKjwr�5��ˣ:��S�k�w�*-j�*{�����Q���QJ"=�N�$z5��q٨��KA��Yet~���a��}Ʌ��G�C�c6gA�@t�r+z�J�S[�����I��Vpu��X!�.N�������7ەڒh�m^\+�o��uhH��=�+N�z�%�����<�V��u+�#�Jm�Q_�{2"NeI\�*�['������9�mBU缒�����s�n��Դ=S��n�>=��-�%�_`i���#�^��/KqdN�r�RMWTi�Q��7d��[�uY}��˲r�S�h�f:�erƀ��.���|�<7�w��$��^�'��Vڽ[E���o���D��йOY�����G�u�[�F�eN��f���<��ogu�#�e�e��+^������c\(�����|Z��<�|��|=rdzйco"��e�vk���{&l�g�fnP��c��y�ɚr���M�
$w��y�[s�'�5s�?o�J͙���K$�
�xG�5�f�;���u�}�d��;��Щ�@t2غT�^�bn'|�Ւ�3I��O���&�d�c�0Y�׌���u�p��YI��3Yu0 Q�A(
Z6��m�[m�1�
�lJ#b5�[j���iVը���������"#,��5Tb6�ҥJ֥-�-(TQBցm�D���T���h[F�[Qem�iQm���m�--��T���JŶ�-(ڵR�mV�*��,��6�)Q��2ʫZT��6�m`�%T�[Z�R���[+Z2��mYF��*�T�ڵ�c+b�*�D-��U*�-T)h�Ĵ�Q!Q��[�J��KJ�(��cZ�m��+RҖ�im�h([-dm���Kl6Km�-(�id�QmieE"�U��0Ud��mk�J�Q+"5X�E+Qb���m*�YDR��PVҴ�*�!Z2+mB*R��J�X�U!U-eE��b��A���X�VB�X�[RRءRڵ��YYZ5����j"��"�DTZԈ�dF(֕
�*�4mim-��V���FR�]�by��Y̹:��8�Q�ce1�;����x{t�i�tL��r{r
{���ȝ�z�>,�y�ϣ��V4�ͮ_tŸ룷C��'6x���6;W@�bWn�;hIxH��cV�齝��p;l�\%�nl[H�p��p��wc�F��|����Q�t�O ٮ�Zt�`�m3���^��0۱��mX�y\���	9b�y��i���V[�[(q�q����w���\�ms�9�u�&/U�-��4�m:]Š��9�����D��n[/�'tg;m��N��x�v�;<��6(؛.j�<����m����NRz{v;c[���&��ܽZ;K�t웂�Y����l�n���ʗ`�&��ٹu��1Y73���i�ާ�v�1<z��sd�a앗Mn��u�W3����5]&��ݦ��o.����Y�c�60��:��<�98�ڷ�؇�8�gh6T�z�p\xnq���ۤ�g&����TN*�٤�7�u�m����ni<2��W�%���ʹ�n����э��y{�xs-���ʖv��V.E:u��`��ی���q��� rݕ���9�B�;�'���Fw��rY	�aW nmx�gn����WDu�Nm�/^Ī�<B�6\���-�;yv�.w^ñO�r���v˵'uq�y��g��x �����e�#��C�n���;�y��})�oe�n���^x�1ݢ�շcjMv�1Ӈ�b���k�sv�76����·��5�8� �6^]Ggp�v�R`�^Z�m��S�)�j^غއ�V,v\c�n{;t$i�n8,�s����p���\�7���8�l����79:(��ͫ����������&^S���GUL��#��r���Q�r�nwm=Y��`w���c�/M�뷇m��vdO ]�ڈ��&ۍ�ۮ�m�ݎ�Gny��hK�ݎ���ⶌ�p=���m�uj�S]^�/A0+�pl\LDrst7s���������o��!ۧ�L�G��;'u��Z�u�<V��N�ۉ�<\���������q�0'�����3<�v���+<d��V][vJ��6�<���)�>P�/Yȼu���Aʼ����Gq�N3��z���z�v��Ӯܽ�<=���`���]��O�Mnpk��;7d��r��k[Q��wl��z��IPTk8��q'b�A�E+��.��ѭ)�unn�7t.G��n��x�x�j�����=�xĉ�|�c	[�ߜ���s��� �u���� ��U`\'��n�vg`5�9�+n�I4���D�%釶Z`9�Y-����˻VDz�^˱Z��r���� p��+s��� ASڑ4�X0���~��,\"��e(�-q��I�{�d� a8fy/^-3Pþ��;n��ό�p����%���z3�ݰ�K
�S� ��v��D�ޕ��tb��jMj��-*yD�$�n0�"�`�4�?y��4I&u�V���^dJ��{tB��������vA�ޛҨ*1o�ߋ�7���k�tsW�=l�m�k�ѫm;�h�8;]�tk ������~���#��E�,���ݫJ� �ޛҨ'3w-eT_ww:�A6= ���VW<�d��dEN�� ����������ؕ��ܞ��컚�MLu�z,�r��Ϧꬺ�q��`f��+���GH��*����x��((�T�����5��� <=�+)A�$����� M�T@ϻ�|�N����M���0�q-��s���@�=H���/Y��+x| }�w��J[��W� �ظEÂ�P�%�ya�������XN��M��$�;� X����R��[���r�3=[w���񔡂mʆ�eD� �{��@|��&�Z�7�C�&@�s���;���������ߛ�D�p��j�<���M�go	sqp�6��׵E��=�Δ+utv �h��m�a#0�M�f�ZA%��w��A+���ɇ�X���Wr�����I�s�M4��&�a�"�	'����q���x�WX ��c� ;��D;U��{w.K�L�\L�Zڸ�-�	�*�L�	UT�|�ǀ�����)�3ƱW?��r��-��@�Ӵ_N@���&\�םgB�x�[�n�swk�9�p��`���G`���Ȣ�f4¥��> x��+���	�ޚ�*ۿ�� N�jf	�#j��˽�b�79lƆ �j� ����|$��ۏx(�/2	�E��#���7��44��-���H ����%D�;�J���R�kw�� >+�����7U���"�
&cDN�c��1�5�����˺��GN]x˙m������-ن�.y,�{AQ(%�^�H�]��v��V��cC��E%D sw���9��`�Fa�(�ھ�i�ouv�D��R�z��9߀���xߒ���Osl�D��~��(k�gp9��H�9���a��H ���ڻ4-�}=\�Pn� [��Z^��[(�
l��y*�z����Wc�1���wv��E�7���3<��t����6���wƽLn2��.�{ty͐6�w\��
�_g,7�l(U�,8{y��r�g�x�wm_x{�'��lt)I)-DD��a�����2I4O~yʊ�"@���}�wo�1��<� �W��Q�s��N�/����}��),O��C�. �WF;=��DqD1�G:�#v���*�:F{^�����0�*$�8�\sI"ws��։':ޙ��T�@y�R�L7p�%䗖fv�ܭ�a(1`�����2N�c��b`���z�� Y��v�@$g_�=H>��-k�
�����꽖�
�SD��uh��H%�oiPu�WkYe���D_�y�WdK�:�MRG��.�Xf!6MSN5B�q��9}�%�K�^]�X�I+��;_�_L�k��c�]W�<8����ѹ�_�&0�X)�M��JI���v���!�\�K�/$��� �l�D��0���8>=�N�C��\1�g�����Ųr�x-���B�x�kefڈ�*��rR����Ȉ8��]E�EL�����NtE ��m��m��{���n�\ҙ5v�֯'IoAˮ��m��y��dR�{�m;��]���V؝�rP��gu��kg�����x�e۲�;da�Uc�0\�[���t���J��ӌc��=�'*��!�;=u���ݻz�v�s[o >a�����t�뷳��\c����;v&�Xl��&��ԸKe����#�����/<V&��玮����Ǧ4�0̞Þg�����t=X�����n\5*I�����we�� ���h��$���H�I���uto�H~3��Ob��jLB��':�8�	Gv�x�����wAw_�*����d�	 �9~����ZBܩ�`��,��]P	wk�
��A,�lϒA"n���ή�n�߽�� �7o�D }}�$ϒ@G�n0`�,0E�]���v� {�7H��^g��+s��NT���@���	�|j� ����MbQ�5�̤JJ�wj�h��Z�`m/{PJ�$�&�D�[��v<�j����<
6xW�2�C�k7�69۫@���b�e/c]s㴞��%��R��$��of�pD@d�2`\���h$h�� �$�ĕ��ۢy�#�&2ũs��p�$׷rd�K|��ә�mz�=�wvD=��>��>��XG�NI�ݨ�uhѵ���#\�0�����m�m��Hȶ�K�����)�Ǵ7��1�{�m%�{�����pT� ���h�I+��4'��s/��av��]���0��UR��fR ��H:$�3�{&��jo�v�� ���4�I��{�e最X���L�4�ג���ۧ��N�$K�l�D�h����:${�x=����� =��I�$��fKp��$Q:뺶�I�m�yP�{�=0��KϮd�d$���ۢm#�oMz���k10B ��4;-i#��9�]F��i]���5e�SF垀�Ǣ'hf�p�&�1	�0�fRI����N� �y�>����TKk�OV��2�Ix-�ݺ6:��� �tw{XF�������W�a�Y阴���n��_����T��
ݯc��	�r�L�n��$���DD"�M��R{�wF�D�^Ț�I.�۝5�պH;���s�K�-ǽ2�P�-���b��MO֞�Zz�ż ���w�����Y.�ʺד�b�k���$Zܕ".5���<2+�$��A^}�wd #^ҥ@�fղG(��Q��1�o���l@|}[V� }�qR ߷@$:h��_~$[�����=�nE`���H7�=Q@2�� M�_������iNN?7g$�;�|�Q 
�{�x=Һ�akT�hS�~1���#A�i�1��1u���X����$_��rIa�ѻ�4�(	�H��}��b����� ���"eM͚Jw;y�.�s7�b�%yv�P�I'\2�E���K[N-$��f�5dn_f�UG v��P [�� xqn%��aw?{zü�\�p��b�"=�o�E��~@ ި����~�ڰ Gue*� >�}�@�,��*\�Ķ������@u)�T|�s��(���x"u��ϴ�s펟]lz�3Ke���ÏC�v����/)���f�l�66i�c����h\}t�S�8�@Vh�Z��xx{�؏���I��ظMC	��3
Q���~@ �7�mTn���U�)�H�i$E�����5ݻV-/M�&�?:ͷ]�>WL ��T6�#GSǎ�X�+'n8Nٽ���+[mH�]+n���~}�ܴLI1\ݾ���^�� {�ͲXr�R$jF��V��$���6�S�'\�~�3
��7ݝv��]�ު�
��^�ӛ�QQ ]�y U��v-hM���/5tu��[i�*`d�^�E=�~@ Wf�Z�""=��a�A޵��A��� 
�ݻ�����Ɉd�4�*�ټ��L�^z��ܗ�H��ۻ� ���v�ʟ@�����ā�=�8�v�1��\@��y{wv�D����x�{��z����q� ��ۻ	'g�ERy}p�g�+�Y�O��9g^A��Q�����̡G�q��Jg��v>l{nrUy^f�$J����A�@�������}�ۀ\���7v�i3�C�]NԹ�'��Ϛ�ڹ����6�w;y�9�whLp�X1q3c8%����!Y<kb.��m�.�#��:M�-�0`�܁�Nw6��n��Z�lM��;s��N�ѻv���ݞrq[i�פ�'���v�m�y��듻=��ܱ�c�|�$��p��:����r�Y'��}/K�E��G+��i<�&kqx��o�3k<��{cv_��[�"�=[�����*�=�xW����}d�PJnf<�k����>��@�[=�$���1���8�fL�I$on��^�N �2�AuInvM �o��wVM)��q�/�H ;3�����J��+�gz����"k`ߒ^>���C�5���$�9gD�%�Y��z�:�RK�gf���� ��`w�]>�}�"�w�lB,2�0�Y���>s!����ꂻ�����=ރ���"�߳}d�+%eOc1>���p��v0�A�A��>��%l��n��{��P�1��3���w�"x�a���=֭�0��ht^f2VT�9�w
�2S�}��>��t�ރ�˩�ٜ��Ϗ4�Ld�ɿ{�����q�Y+0�}�y��Y��&2���<�>��2��| ���r�p�h�XG�	8,�a)KZ9��&�$��-�7
ۇ��U��2ඹ�N��*�uj0bi�l���'�G������<��C���=���gFc:�YXbc1�O5���T��3~�=��Lvy��t�?e?}���'��c%ed�$�]t�#`�>��G!5$�6�5�N�\a�^}��N2c2e�����|�U���}�7ԃ�va������d�)X�"&� �����\6�����D�˸����8�^���qF�&�,N�����x{���������Α�>�J��YS'�w���N��c2!��`�k��l�*��b3�~ۿ7�ٷ��p;ć�mO���FA�<Hnf�T�Y�ͳ���>����+8��Y��e���y��k��Ɏ&2c�����y�WV�p��y���G���0}�>G�G�e>���p��;d�Wc1�<ןsf�Y+*p�|~��rW0sB��YS����8}���sݠ#�>�>D>��'~�~l��gP�c1����u��Vy"=@��z!}�t�����ô�`��d����=���p��%Oa}7����mѦ�ѣ�d�����7�I��Lfe��Y1;��}�_"O����}n8N���a���{�w
�'Xc1�!��`�kϹ�L�pf3���C �"���p�`#��|t�`��}&c+|��7o�X��Z9��oH�1۵W+��+�d:�>�xr!w������a����w�'Ì��{�vgY++&f0��{���1��Lq1�����'S��&'��_��s���3!�מ�gN�1�Ę�qu�٦T����sd%�D6ˈ�}dY��'��>��Vx�3�w�߿z�_'��3��vx3�1��a�c1�kϹ�L�88�I�32e;����<��d�,�L~��}��^����B���x�>�s(�"��3F��`�L�N��?kϷ�L������Y1=���o��<f8$�b`��!�\�L@�/y���siW����V�Ԯ
^��J��B�WG[�[_f҇bF���ȸw}_U�p���Cd�|����O�y3����>9q�R�G�B��p�C\�t�m��ܵ�;��fv�^I�(
��Z/+c��N�ܮ�s#�	 ز�99�ś2�)�r�Y�O�P��s�^�xak;���g	�6�\�G�`�I>�NI���8����>�J ��p�ݓ�5�ojJ3;vt%��-`,�z�a{��ݗ���V�>�;�է��G4��9�V�q'�8T/���D��z�n$��8a����I
��u�gn��ʙP&��'
�E��լ��㩠^��5N�nʚ��Z%u�g�� v�%8y�D����7�m�S��5�}�+�m��H5��F�2���;{��q&n�4�}2.=[1t��G��܎,�(��J���X\��
�h��f�{�lrS�����b�/n�Y�5�������ݘ�곲ݽǂ�A��N��Ǹڶ������}��s3��Ǜ�V}�a6Q�����rn�N�:Պ*�z�H0	ި�v�Hد�q�0�*��[�H����kh�no?�Q��b�|q��~�#�=�J�5�y�˟w���Wa�($�����坖�V����Wv�]����r��o%����bp����Pfu8nor���t^'+k9h�;]n�or�N���5=wɧ�7�f����O�[p���VL�r���[K7E�\O�"�W�.�9F��sf�m��Q�Qk[k--YJ��m+*T-������))D��m����6��EB�X�Q��B�J�m%QR(6��`����ʊJ1T��Qj�[h�EE)KJ�0�V���4����XʢV�U���ڊ�KDh�U`�2���F,���h�bD�ZZ�J��kEPE�e*U�Q[T
ֈ��cZ�RX�F
(�TU[j+iJ�+k,Z��h�F,U�DV����m+e�Q���mZ�X���[h6��1���1Yic�lQ[V��)M%Af$�KF�TQAm�+1%�J�ke�
�kef2�T�mR�����-KX6�AJ�Ѷ��mkA�1�Ȋ�Z6�qY�[LQ������.&T�#mDIm��X�*"�km�&6�S.*b2��JZE�X �
"�5P\B��U[eb�Q��J�ETUT�2E`�Y+YieE�m�e1 ��Q*6�XcTe+j�kj�3)s1X���  �������0�c0C�ȟ��٦T8�f!���Cbw������1�Ny��ƚsf Г�#���G}Ӳ󑰖����]~�:�YY?e��y��ٮK1�Ld�VJ�~����'YY*yd�fQ�Ut�#��ׯ��g��G��:�٦T�a���y��պ�\��9��Xb{Ͼ�~3�!�1�����b~���gFc:��������}_����c����Rq�c%ed�����}d�+%��d����s�½��LL�s�+W��S�D�p�$@�� ���q�B1�sZт�s��f3qe��<\[��}��T��.�x�S����7���LfY1��LN��������c%eLc12��{�Vu:������~���y�}��ʇ��f!��c%O߿~�}a��3g��y���֭��tf'{�����&e�ɯ9����������of2�W��Lq1�����O��LL1�2���{�Vt;d�W��}�y������~ٌ���K����Bl5؄���Q�=���޳+%eC���O~���јβVVJ�×9�7�5b���s���Y+*O\f2T���{��y��r�d������½��LL7�|��h�ѭkX<�'Y_��Ȃ>�_.���􏶲{O���>�>��bo߻�}d�+�����2~������%egD1���5��c*�w�Z�7
�����b������E_˭���9O��|��6߫b�Yt��r������[�ҢR���K�)�Ǐu�����HBO����b�O>������|"����C!��}ԝ�3��w�p��'r�d̳~�^�b(/A���Z�9��h��Y�>�"��ٶN��8ɉ���ʞ����Vt�\�1��y���S�1������s�_��>���?��WeG=��Y ���`�<V%����h��n����.??{����x"���+%O7��w�|���b�d�����ݝf3����&3g�o�p�W�Gȏvm��0���S:O��Ȍ�{�̞yf2VVJ�b}�y��^�Y1���ۂ��L14}�E�>ӓ"�`�c0�&3�45�zܕ7���}	<f8$�b`�����缅gY++:!��by����eC��b3�n��+W�uv�i�=6|4�>���FG��n��k��ĝ�3����+8�YY:e�����{3�c&8	����S������u���}��u���q��LeO��~��;d�Wc1ȇ�o�l�VJʜ�o�2�˭��ї\�ΧXb'��'��B�u1����>�A���>�vtf3�`3�11��'�o�p�T�q��#��L�}��w�'����~��_S�����d�1=��<�+�Y����vQ�E60�8�������b~d�fY1�d��߾�}|x�98k�~�9<='̌>}EfWW�>��f31��O�o�l�VJʇc1����}��a�x�`�.���?g~O�l���@X`GD0���a��\��
�t��'v��0	�m~������@S�t���oI�V�D���.���=�	$$�ם��H�f�f*/�9�u�zT��#���UcV���Y�Զܜ��wn{mb���h�p\��/)�3'�Yy^+F�}�[Z��-sѬ1�5S�4�Eˇ]CӼ��/X�rq{.�����q��%��5훳r���s���'[j�Y����ԿOb���^y���Y��s6s��lk��mln[[]g\<��{-�Z-�Nܺ�70�6D��|����ۻ9�x"�Z�9�M�[h�e��8���������f���Y��6�$��b{���a��:�YY2e�����{3�c&8&2c�1���ﺰ��Fނ:3�셻7�#�3�2���<�+;�&2���~���S�1���|z����Vned���Ϧϻ����}�|��r>kuK��4�߷ݟ1�Cc1�D�c<��ٌ�8�1&8�ḑ}��w�'��c%ed��s�����~?
}�{�¿��&&	�ߋ�8,�L1V}�E���rdAd�fY1���~�������c�&>� �A��f}xf>�:���:�ڟ��'�1��C�����͘��YP�1��Fbw߾�~0�'��s˿�f���$(Y����"����/��G���L�Yf2VV޻����d�VJ��ɉ��{������Led���>߳��������o����#�}�v�C+%eK�y�[�u�W3Z2�pY��&�y���!�1�"�Cc1=���bϠ��'�����o��O��|"�w�1�'�0q�əN�����O,�K�c&8����{�W��d������~��:40�(���b�C�)䋭͢�j�aѲ�L+�=������o��a������S��|޽ٌ�J�e��d��߾�}d�+����f&{Ϲ�!Y��f3{>�����z}���>g �o{��f!�c1f3��O�}��񓬬<9���&K0�'�}�|���v|�{�/A�����������dh�6"��'�;+ՠ�J�����g+r��9,6��׉��3���D:#�' \��0�J��\�f�.S%�sO����zs�~a��כ3��L��c&8&2ba��߿��'���&2�VT���gC�L|�����������ǠT�\�>�>�3%��V��0�U��YS�Oy����x���Jʆ�b~߾��γ�df3`��`��Ǘ5�>�|�xc*O�3++&e=���o�O'�c%�f3�|�����Q����G8l��ʄ�g�G��W;�A�`?}G��F�}K� �4[<���؁R�
���{�$x�>�>D]�/����_v�k��m�!���C�����a��3`~���5�[���j�p�1'\f'y�tzβfY���c�k���Y����9����y�W�c&&��o��O�Led�����P�;�&2�$�c�y����eNf'w���g�o��m�0���-�۞:��s��7c8�\'	�x�yQ����;,�"]{�DCa���'����"~��~3���1��3����P�8�Y��J��<��ጬ��'����i7�u���翷�O�Y��1����ׅ�H��xq���� �ȰG�5�혜++%c����u�8�޿}����Q%ac
�����aRX�I`���f$���}�u��m��of;�������zȲ ^���(3�f�8m���?y��<HP������g)
�k�y�������~�f�ۜ�]��i�3���C���h�9Tǩ�c��	���}�����՞�eO:�t|�q�-��̔4;ȡ��&�!$����~H)�+���n ��%B�����Ì+3�=Z) ��xY������"���덫�
Aa������@��׿p���R���~�`{{�����y���a���w
�`T������kYs4殴�N$��{��N�d���"���@@��;A�g���#��}=P�80��s�vc'T��S���#�E�ͥ8x�Z%��jAB�[ps�V��l#�'�c6�m�ӸF�ҦuH����7��q�*!�����|.���R���h���ى�`V�!z����E�"��M��}2�g�O߼�w
��
	*��lĂÂ��!B��Q��	�|��� �=~ #�N��{��F������}�>D�^��f���
Zw߿}��<
C��˸�
����|����#��"�8XPڇÀhd_��љ��$���=���l�N�aXk�w�w�y�s�*AI�
��s�}�L�VJ��YS����'bu��~s4�2Y�`E	>�Q�����b.�~kʐ�i
��矶k��H-�
�~�����bJ�YS���ۅg����]����ׇ�]ʴ'e�o����ATnM���<�w���:t�`�߄S��,�|�J��"����V���n�� !?���*g��i�V[���h����u �����a�RT+%X~ߺ���1�^�x���<�~�7�bA@��;�L#X�
Z{���;H6���o��R
r~޹�H������00CI6��m�ˬ6�Ϣq��qh��i�Ӗ�c�V3�y%<������w�ԋ�kK�
|����٤�H,�%N���蓨Q%aF���_�
�Q㇧cf}�&��Z����3�X>FJ2�Q�;���:'P/�;��֮f�nc��:����u�À�B�C����s˶��{��$�h��O=�����
������
�FJ��#ȁ��I|�&r�8�>�$2<	�y��2��hu��� ��
���wa���VJ���}��8�d�*J�mP��wNZ��~����G�"��I�}�`q ���C�}�ۅx0*S�;��p�8�E�=���E-���H����m�� �oϼ�ԝB�+
0�,�Ϸ���80�%��~�Ͻ�9."�t[9�>�#� |�{߾�:'P,�w�1��ˡ��8g������8�����v��vk�HW_���~47y���R��{�:�S�e�}�ۅg*AB�;���|(�#��a�S?}����T	��Y(<��e��-��
���\��B*~�!��́N`-�tm���n ­Or����G� <<<��⟂dP�=�wj����s�$InS���� ��{�l7)�.��ӎ����y܎�8h�q֢�8��]��]h�����^�����;��ֺ�k�=�E��k��׎�9u��Ct�j�ov�0��Ӷٓ���	���β�B;���.����
�$e,��͹�ng�vΙN.q�=�<l;h���7nºm�\h�����n]q��T�v�.��N��T��Δ��u�*����8��g���(%��O������8݆a������O���$���+��_�
�P8%@���~��3�ә�/��x��-?o�;�;�A�x"�_Nς4|!��Ap�d� ����2<	�yb��K����^���>I�*J+
y����VT�
��w;��4�������G;h���zȻ��G�d ����������:����u�ÑĂ��@W�Hdx^>�D/�9��}��|��@��S����~��¤8��P�w�i�V�^�es5���`��TϾ���s�{��w�� �~����d���@����`p�<	���� �&cV����b+G�hx"�j~�k��"�xp���1���bO����q����d��w� 
 8�� ��i�����?T+0�%�{����2r2�Q��@�}�t�Y@�S��`�p�E�����L�g��;�Y:�0e���u�N]%��Z�tl�j!����J�f|$��(�߾כ$)i��=٤��0+X/~����؁S�|��|�鍯��8�Nk��G�}�G�  @����V{�����㫅��Xu�Oy��l;�JVM��}�g��k�n������椀/j�w^�z]�b��u�u�:�i�o�N�{�M��l�9w]Å�dx46��I�v���[+��IO��y��͟��J2��}��4��k� �~������A��74l|HN6�꼹�G||!;��֌��WW�)�I�����AH,�%N����N�aX}������yׇ�w�s�B��0�(�ID��y��$N2�VT�{��������i��� ��|�|*��{;i[�6M��܉�HR���vo��k�`T����N�K+*~����Vo~w�}��Y}:�����@�@޾b��|[�y��sZ��� ����6x�d��?}�~�+'�~?^y����P<��ݜH,5!Bӿ�}���v��E�S����$<�����n���8�uQ����v���t�ܺ�b�#]��;���S۱p�j�__n��6ˇ���O{��8�@� �����:$�AaO�>o�;^�W��#�:���u�wc?�X�׿�q �q��������'DY NeJ0P�(�,D�>�>���(����b��)�E��5����H/�
�;���N�,@��?}���+9*$�f��^���6��S�To�q�|��RH�
Pd�8�S����D:��Y++��_�q��YP(��~��e�g��_w]ʅY��dUڒء30ڗo絝v�x&�Y�GU}�
�A�7����P׺ݜĚW6�]�RX\@����n����w�����?�@��w�����k�H)���{�;�A�!Z!�����W��R�3KP�P�i�&��z��b�1{Ͽ^��Z~������T�{�vu'P�J
����+0�*%�y��2s�o?s�����Ȳu�������'bu�o�/Ɯ�Ѫ��������ą��-��>Ѿ�o<Φ���������'>���N�(�X~��~�+8�P���D;���>�>c�ӟ2a�|C�I�����Q=�.�>A�[$���$��Ԝ:��L���'��o۠�P�*!�0��'��|��vt��2���5�p�� +���G�P(��w���1��򧟾���i�B�C����¼f��Pچ�p�PȰG�3�(�����9�]k3��LO�sg�N�RT�~��r�T�B��w�����ed�+&�5�o�������~��߿��8���+��˚��tg���]�~q �)h����)
�Z�"+1d]��Ro[�� B �����³��
��`�{��8Ì+~��+fZ�70�aS�}��Etԯ�T(cΣ@�<	�����}�<���*A@��}�l5�Z������ u�ם3���Za�ّ{)]�؇<Μ�� �����[X�5��B�p���R�V�;��J���+��ve�v��M�ww���HI����+���w
��7��l"�i�&��#տ��"� "<	����,�Y}�����)�����9
Ñ�H(���6������VT�{����>?x~����q�>w�6��ss��sm�:�|��͋Saw+����Ԑ���Q�!�%b���7)��u>=`|��5�À�B��P?w��7�����~�݁Ă���v]a���?�}�sp��2T(��b��(�Q�G�O�m���	 ����a�IP��|�����b����vtf2XʁR�_;��`q�
G�	ﻤ~�<	����9�˩�V��p�GM��0���وb$��O�y��'++%H)�{�Ή:�XV���Ƿ�������u�*AI�%N��q�����*AN����
 �ʥ��CD6�||;�y!Ώ������
C���s�7��
�}��v�H,�����L
��^�t�=�����  @ux�0�)�s߇+fN�V��XtaS�}��P�Ad��?{�~�����������P:����l��X��i��{���i��a����¼��U�z��~��'���#m��E�֔�#�ޒ�쳌q�P�?v���෡����a�z�uZmhZ3]::#+."�AG�{��c*���b]g�����\aWt�Wz��u_���'���V{���G�^��0�������5�j�70k91�)k�'�e^
���Q�㯟.���ܯe�csw�������ɽܥ�@�q)+qmI�;e�6��Q*�#ք��������p��y����x�bp�">����W���<qFY��{��\%��C� ͦog+�a>��S��&�lK�^M���(��.�7���6�fn^�xO$����-�fJnžo}���}�����i`m=��A6�����]�)��d��x�	n���Ou�{ L���i�NS��/�}�Qy�'e��'l9�ӷurŖ	�G��t[v8;fsh[}u{6�T=c�-����EK[Z��[�8���C�sӛj,���^p�7���{���{=q�`�3)����|��c^�(b���9��Bt�5w�`�`������06{��Q��k��+�=�ٷ�c�����B��Q7n]q{�S�\�yɳoh���kH���D��Z�9������}�@R��.��0
�.W]`:�|ͤ9�p����}9�G�V�p�v�����=xj��93^3��Ip�[�7*�=��N�)���Wf�W��[��(|�0e�;�����M���]ͽ�K(Ozd�*^-� ��j>�sǴ�tҮfeeTQY�,�)K*%���$m
"�Q�����H�R�X�jPP��(aiF���*V��Z�Z�Ub�Ŵ��lF9AB�*��+�V.-��eAFZUij��DjUR����W��LJܸ�Z��*c�U)\b�1�m��eE[J9h���\�1!Y��V*JѩV�TE�J��AƎZ��PF�cĬ�#8�(�T����D���*T�UQLJ��a�(�\�U2�m�f\b�-���YQB�����#��J�m�j�J�1�5��-*hU�T�k��V�$�Y
0Td�bfZт���iZcq�\j+2�Qb�0jV�j�+�c��U�32U�5���4��&8�c�6��R�f2W�C2�q�����F�@� �J"�h9V��X�ʱ
���ۘR�*��
�KJ��%j��+3-�c�T�[�[�1��F��
�Q-#����B��e��?y����m��l��1��::]���9�iw��y���G��u��W�^�r�����j�&Ƕ��A\�Pn�A2�s��s���f=6-�nZ����l�	��v�7d�YTv���\�O�,P,k`#��=s��<v۴W�LS˸�������=��gk&8s<����]��Y�����ŧ$�n.۶�ٷ��R�ޠ2�VM�z�;o\�Z.���&�j%����[[m1Y c�h�،�[�s�L8��;m:�nA�c]��U+;��8�,��[R�Gq���x
�������c�����b����ᵺ��\Aѭ������L]�kGaYu�#z�m�
���m�C��8.�.'�zC��؎��6r������������ ��ڱ�S�lX�N�6�s���qζy{[E�Zθ��/#����r\���-�����2�ٷn�:;;l�\;qX�vv��,v��qv�%{q�t��)��nL���m:�g:._h�5ڡ�<T��`����N�/�q�;�ݒ���Œ������zs��]�>y�nm\k�S�q�{g�rr>�ÞM�`+��ݛ�;`ܜ�
�&����e^�Ǝ�A��N�y�-;��\u��n�d�pW�b<��zvJ�v�y�+�>x*����n�������@{V��u��m�R�l����<=v�v��#gtUձ��aςx�l��WZ�'j��۶ͮ-W[�;=;6�+s�v�f�)�۶���}�����;H;��6㰅�v���.���S��@s��ǚ(LX����W�x��`s�	v�ll� �,�Z��ö�Z<�48ev�)�]��%89kW
/N�����K���,��el���ۏ65Wmu�]=��I�����)�(9����U���Œͳ�܃���p;`�Nø����;����ۍq��m7=wh�xr����皸&�M��<a�qzi3u�|��;F�è���X�sױ_��������}ۭKk{�&-�5�Xǵ\vZ1�73p[#��S��'X�q���gjń��^�g3s�Qj�u�u�jXͅ���'��N=q�,\u�r��+����dʓecI1ÈO��ǚy�6�F��:�n+�qwh��xM=�[��h���9��zx�i�|�=�5�Vݳ�m�c��;u�W]�6F��g���'�ڬ�qX:�t�\+����Z�kټ����Wn��8q���ٚ��t�����̺k�Z����?�Ny��8�@�����߽�gRu
	+
0�)����B��
�����Ο߷��9i�g��&�oﻣ��ed������}��������tesR��e
�} Q�<Hxe�F���Ql�����ލ�R��Z0*S�~����R�V��~�*AC�*����~�e��|�59��M���f���aS9���:!ԕ
�X{�5�g��YP(��w��o�1�����ޟ0?5�F����{�8�zR����n�0*S���)�浐�1E ,�#���ES��� �td��%L���l!ԕ������°�
��RX��ϴq�7����������d�+%eL�}�d�'P)ϼ�.WV�f�֍�lA�=��y�T��� /s�&���;_}x��t/���Sg�����a���p��2T*J��}��80�?�{�ϸ�^��}�_�l��ɖ���.e�<���)7e^�ՇD�k�iڵs�F�q�������󎮮V�C�>aS������N�Y(������²q��@�~��`q�}�w�7F�?�[�A2<%!7r ����?{���*ANf|y��]5ѭWY^ �"No��8�@�������1�����u�	�D�Sm�И���\w��7�t(�����wL�ʉȴU��=������v�ב㹯�H�O���ݟ�:��+
°��k��R
AI�;���d���c+$Wgވ�"!�H�=��N!0��N`u�9�k݇#� �~���7��+X��=�oo�g�߼��=+*{�7�p�	*!�|�GpV^k��h�3Z�u��Ã
�Ͻ�Þ�w��ONk՟��N!Y++��_�pf2Q��@���g��@�<H_�wH#�nu7����@��r|��d�a(n!�Th���I�<�G������ﻤX#�@�g�1_u\jg�{O��|>�5�°�aRQ
�����2ped����>D_}� 
 Q�\8�]�/�툴���/A�`�݌��j��1��Ʉ��m���]����C9yܡ�C`���'�|
>��^l8�AH(��to��� $+ﻨdxvz#� I���O��2T����>��aXS�9��U�f:.�p�:�S߹���=�����w=�V��sg#1���T��}�����
Zw��`w��i
j7�B0��u�b�h�wO�6|!D|}��]5ѭ]\^ ������Ag���T�{�Τ�%H,9�=��}��W*���w=����d@��)A;�j�#m\�5�����nl�����^ߝo ��f�j:>pk�Mk�?�_P�w��B���*J�ID���������S�{���ƽ���e�b~�G�qG®�H6�V�Ō�HxP;�h�)
сZ���{���t B ��}Og�/��VSϩ�o��?	*;�4q�#
��k�WZ�nf���9��L��wa؇R
A>�=�@������{�{|�|B �����H)O���݁ă�R�}S����$p�2~���u��I}J=��6#��n���X��Uԭ7K�+!���-m��L14����1�M����d|��;�'"ed�=��}�C��G�>�=�|(�"=��T?��G٠ZN'��8��������<��}�:� 9�Jh�l0T$�
�^H�x$���Am�03�L�ހ/��6�R���g|��xS���lρ#��(�@�M>��_T���{��>�=��k3X�rH)���퇨u ��������c*J�ϟ��Ξk�3����g��Z���i翽�`w��e!Z��s�7�`�G�b(��j	� 	ߩ�'�v_Ƚ�����J��S>���!�%aXV����Aa��H)*w�|�{�����Yn">1q"yNf�KX�=��k�A�T�p�}�p��n%M�\]iK���~�`�{o�*}Ep�suWr�&� ɓ:� �q��R
y��~�@�񿼿Ʊ���:�:�Xo��{��RIh���F�Od|�θ��)��l�B������N��'���7�*%@�}�F�paX9�/�r����b^��t�[u�W[+ۻ.�c�XÞwm�{[n.:����u��0]{�L��a8�����DEw\��C�(�d�+w����*A@�*{��6�X����3���w��C�i����`vv�l�+P���sp^0*y�}�a��l4�R �=�_H�/�$i��}n����љ"A �*��I�k ��}7u*,(l�XLm�1�'ƫ�ρ>'������2��]x�v;�V��"��
!�������"v�&Ӟ9�>$�n�&|A���k�:�<����JZ/A�L��i�$H�ڙ$W��+=�]i��3}��+�� .��S�"����٪��M1�4a�/FZ;��x	cENI+w4�y��:w.����x��j���'j�ŕ)�@e�o;��zwTb7H����������`A�`�l�\v����\�<Wm�x�6�ƹ��;�����׭����Bw&���pL�1�M�H;-�8�F?�Y.�+���e ۹���=�F^0]�m؎��uvs��ݲ9�ù��6�`{u�#�����s��D]�sI��p�8x,d(�q�me���ɖ96�������vٷ;[O=[��@�Z��GPN=���s[ry�q#ͻ�3�;��9���mF��D6�g����~��4ܝ�� ˬs�AY�H �vuW�
ŶT��b� ��ɐD�Y��lDD78T��
>9�7����έ���I�i�� 
ޞ_*���_&���~n��;~a�[a(mU{��d@;��B��<�,�<��Ø�g��U�	"so(Q�B���	���r�W��j� �SV�Ē	���I�x�L�L�k ��b{��nwz!80�^==�B�$�rv Km�	숒u�ȒNgf�x�y�2C�t]��=2��Ư獳��X�b6�Yc�{bkuv�k�;]bB׃![n%y	�B���������f]����}� ��'j w���Wfox[�}b�N@���7��[f��C�~D7ϫ+'�H� ���ܔ�1վ���a���Ƶ��uY�&��W��Y���*�p��P�W9�,26�ҍ�T� f����A#�s����xg��[�c������Ϊ���؃�F IYU�D�w�d�	��Mk��<�������^��{y� ���D�P�&ښ������W[78$M�$�� �s[�����y.�|}Py��/���$�g:�6@L 싐�w�"�� �t��*}�i*T��@Q�y!ٳ��K�b�4P8���
\Ò���m&mwYs�iz�:���D�Zc<Ab����4�����u���(b ����m
 �l�O�$��ު/^d�4flV�q϶�'z^>]��ڄ�7�#kk���wS�'�y���g�A��3�I�]�U@4-&�ɝ�x1݉�ۄ� _�����Dk/�h�F��Ω��b
��c*xF]����LR<Δ���ۑ��M��щ��.{��ݚ��z�nj�Y;��v|eA���<����3e�A9w�U|e�b
��1J�����]�J˝\���@ S�ܕI��ьt�Ȏ$��D<zg���� �Zl���\�$��v�$J�kT��'��"A#��$��ݯQ��K �
��M`��8��T�lLr�un%�	��p%*�
Vۣ��\�{�����:6h��/����H5��4H�&��f�{	��2�<���A ��t��Mi`���DTw�:�b�j�6�ۑ�$�؇�G��G]�Ux�H��j�wv��\����vp��wA�M�
!�D��]TH$�_mQ$��`�&�7��#�u�'n����<�h��!4EU»����`�sU �|����
������ ��ք��b��ۼ�o�-=���X�Ř/8s���~�gS�h^+Ϋ��SU��݊�v�y��2��`"��(ٸ7��xH�¾�ʯb���6eD4@�9�U|u��o��0����� S�ݴ����:I}W�11[2F
��e���p�w�lč�q�M��lF-�����[NT����~�uha
!����$��}�Dx�H��@)0r�
Y	<�� �@9׻B�.Z�& 8%�mu�Z���O�]Z��QY6O�>��ڠI#\v)!u��:��=�z&��P�p!C����@�0�5�]�r�eٔ��;�Ν <�rT	���RJ�7��M��Cp�vz[�o�-�R� ��A$��$�+/��:���	u� ���Dp|{!��h��*�e�ـN]��W��(S�>%�Q ({�E
Q�ʟ��R��
���;>'�]��O#��Da��H�lSz�����&,�׻mK�;����G��ܔ�4���l�B^�|n+w �5��󗪘 [���̉$����M�:9=��B�q�q
s��j�S�m�$��q��/���D[�-ҙ�k�ܙ�g�OTf�1Z��$9�����rsθ<�>rt���ۻ3��lv,[��e���L���Z�����m��a�6)��\,�h�k�m�󻵜ۋ���G���Gjz�q���ԧc�����|���5Z���ǫD�a�� �;S���V+�v"O7lq)�"�S��5����=]u�����>8�b�I��Tw1X�9z�(	�1I0�o�Ce��(�*�U�U�MI�s��6�$�]�@$�ު�$�Le=��(����nee$�
 8%��Ղ	>;w�"�$A<:�T�a��:FGLv)$��t�ȝ��B��PL�f���E&I)l� �2ﺨx�n��N�l^U�`��J�J�;����q�@�[]U��ݪS��1vшC{y�bA"TUĀI"��j�"�{j�];w������i�!d���ܼ�u� �m.6\%v������q�����;��}�Ɨ	�43��"��f�>$]�mQ��ݵ���Ñ��"A ��F.�4�2Sd|Vu�z�Yr�a`������I<��{����w3
�'��rh��>1���l�V�y�Dy��nq�wn��i�&y�/�V�����r��1�8f���$���M���(7�:/��zQcr���<����bCBv�*�I'o{hQ ��e7��Bd��Uts� )��*B��"�\2�5����c��TM7r�h�	���R�+��Y7���	�+��$���(Cp�C	�T�wM|p��ں\P]�j {��q�K���kt��o�FS'V�����K�͹8��낳��k�݅v�z��a��ߟ���~�iZ�����Ox�n�vkĀN��#�h���UT/\zi�P�z��x>;p�p�8"t]l��6��u�7��S����n�A:��$���A{��U��a�a�6ALIY�SD��{ H7ԇ���8���	��D�ż�һ���,���{��kGj$�$R6�ܩ���U��>�Ǘ�蘎�t'G���eu�F34��fr,)�*��́{�V�*�W3m��^�>5{ ��-�oc�~V���k\�={Qfb�_hD�{�iS�l|�F�}ܦEa��G9�`^��X$�e��Z��v�7��yx7ƗތK�t�����{�s�ԇ+ދ�|e���$*�{�ٗ����5�������n-z�A��"}��O{��՛����,5����-����.��q\M��I��=�[^2��	� {���ν���9���g�	�8h��[Mw�aL�ZA)R�s[�p��ׇx�wq�=ڊ�d>\��gK˵W��N7N*�#pws���ƹJ;�НF���*�q<�Yuhs�:.�|&���mvpT�n�f6�8��7�]�7�2ϖ�ύ|է�����5��M�f���h+�O�CelT2��w�r.T��.�����gf�U�������VCԴrv;q	�nmݦ6ԉv�J�,��9]y2߫��mc�X���p�A��v�T܆.�w���K:�n�WS�_m����.�E���ߞ�8o��v��kq�| �wN����8�q�����1��a���S�;�zv̈́��P�,F���O�d�O��e ���ԺG�rWT0,uoc�3z@�0�}���³�p�d��^C<L��������f��oyǝ�o���c�9l�E0J��H�-�m��F�EEEUbe�j�V�QiX�DUed�5���2��A��+%es
��U�AAqG-�aEj(��mEQF&2�̶,mQ�����!��(�[B��)�b�F*�f"m-(�+�KaQ���T����$U�\f2#QS30QQPKj��B�b �4*�-��m�j�ţQ��1A�*�lZ��d�2k��J��EE��+j�*6������E���(�Tr�US1˙L�TBңiQAq�G���LFb���YQKV��PDP�+h�Z5(�,FcF�"�11Z����B�b6��-aKs*�V�X�X6��m��Tm�s(��30jQ�lm�ŋ�QEUV҉T�k�%A����X�R�i�r߈M�����BO۟m
�꯲$�v�Yi��J!�ȼ�C����g|vD�@
��@P�yy+��~�]���"�)"�*B,i����ޚ.Q�Hc�;ϒ�x�/h�j{��ļ�ֳ�_8�����v��*N�4뮌gJ0�뮹����ʈ��m�7��X(Cp�6S&�K��}���>�~�UB{��O��sj��;Q|�Ĉ�p(�i'�F��N���RG'�ד^�:��H�H�����>���L�ԇ�A���m$`�Ux���A���l��L	��@��c�S�����

>�T��1�a�)6A�$����f.��	>:�� �+ov� O�V������qj����£ ����=�ý���7��]�p���}���hӣ���+leK����A���+"�5՜:�(<O��+p��Lr�6j>���0~��+��~,4�P!D14:��D��o�@Th���]�P$��ݪ�A�������ӽվ<�,�<�V���s�0���tsas��4�>:7��ڭn��~�?>��llR=p8v�_��zh#+{j���S����]đ�}�F�kK�C0f�ڮ�/kk��@7�h��y�	��T��@�7gs��o8�	���Q�M&!�&wk����v�W�x�]7J�z7+�"Az�hP$��>'��4�i#8"�x���8E�ΙhH�a���O�9]�TI#T�F�ǻ0E�Q=y�zjo*�>�}��[0-�a�+:�kă��5�w6=9�q�	鞉@.�oˋ�R�'��V���7^[B�F���gL����5����X�=sg���`d�lk�W�ӆ؉˶Z�����G�p�&T���/j���u�s�X!8��d>���h�ú�Wei��7c7�n'h:��r�+8͓�a�]pj���	�.�&�ȕ�qg�5�k�!N�d�ֻ=n����c����0j������(�ZL�aM@��7:�:b�{L)M�)>(�6�и�n�;\�n�g���[u����O���vlGm���.�s[m��U�x
~ϛ�N��V#�Hn:�����\V���xS9���7\ƣ���w߾�Cʈb�U�TA;[�B� �]�{'���/G�XұD��9w�Rq擙@�p6�4��3�w6҉"[ڕ�0�n�v��F�ˁ&ۛc���r*u0P�pT0[
�L�N�,�\�O��K���s�����^>і��E��D6Ri1 ��K��;\ue� �w��(�o3�Jt�����t�s��\T�C�nH�N��ژ$���l����t���@}N?5H
��Ί�O*�g�%�ѐϬБ]�m��, �d�
wgWd�������O]����g�;[q�9盏��Jm<�C�&8���
>�՗0I&�s��.yl��/C��7�ĨN\f��r�i��BP�����>3�dNul�畨��~N;�x��fIXp���v��D�a��ӭC-X�͓�4"4�J�JÒ���h�*�,>*X�/������x�<�A$�츒Mf�M
��W]��v:ܤ�(À�8(9�ó� [��-EvOz:΃˗� �G{@JzyW��s��B!�P�l*�v��Ȏ���L6�����` OO%@P"���*wye�iD)'��;�Cs L��$N��P'�]n�
��wo�3�)l��
	�����T�����&��a�n|�|�H�pX�+e����9��۫A�4x\ú��0S�/�f���H9}�"�#+3��Z�"��ڻf�3oz��]��l8��O�5ՁD�5�Q%ʣն�'č��D��Ϊ�U�&�kw�.W�L�\A�NK˝$.�HUAAM{ۣ�8ߧ5���]��7���ی3k8�l���fDS�{����ݮȴ8����FK���=��$M�Rd̿U
#�J�ܤ�[��%p�>:_fN��P��@[�j�@]<�_q~w=|�ݩ��*�H�u��B!�P�l*��[�Gđ{�3�1EQ��#L�T�e�]P$r�:���&�Ľw7�l��~D���љ�mq֫4v�i�pa%�0t؟kn��^4&H1�x�#�I��0�^��I-t�H
�m	� d{�Uv�@P>7��^���C���)�蝛@b]y�z�O?s�P P�y/���zG$e8�統�Jqט`�bm��@B�?.�V(��F�c�I����n��#�3��	'{1�/���	���!��پ�'����62�����H;�j�x���>'��vuw'{�@�`%h�l��=��n,M9�`S��!��$>�n'C��:�&��O�D������fX$�ך���D�����jf6�r�"q�"+'���۔�%BpC$�<vvY s��<��3с��H ��@�OO$&���z{J`
���6-�9B�ι9={v!^����j�����f�V��j���ž|�������B!�P�lD����Q�w.C$���^4{C)sE�u�	�.$�z�4��������u^#&��TMW!���X:s.����D���oB�G�tG]�.~�ڃL��Xn/Y� ���^$dL�m[�0	�u��-f\Ifwm
��i�ÁApD1%��鍳]�'��G���{��H��b�S�ur8E*��k�8�pf�Ϛ�@}<��Gϼ�{������}�TH$��uP���k��M6,Jo�zג�<���Jn��ʹ���Nj�Q۽��N���qo(�؝	E^�2w��;�F-�l�@�ɭ�l���Y�+=�m�V��-,�Ӗq����	۝�ϣ��tn4��m̀2o]��Q�(���cq���@\mQ(�s
v�]�� u<��uwa6x6;��̣��7!$g)n�PŻn7E]z�8.'ig��H7Z8����c�h�uj\;����
�P�|u��D���˷t�d��,s�Lui[Ś�wV���%�����ɇ���"�H���^�.���pa�Tô��;=t��z�wRl�	�q	�_��`I��ٯAy�U�-�{�@j��|H'/{j�5�8�(D8)�a��;U�B�6�Nq����U�I�T���C��U��ɱ�uˉ��y��E��0������>$��m
$���r^'�c�mQ>$wn�W�$��u
<2�d��.J�b;�����Ƿwj��V=Si@s��H?�A��S�}�o�j�Y��m�C0�1 ���':�NYh�I�	����w�������5�1���T����F��m���JiaA�	��-a�e-h��n�Mg�g���n�u�*�����맮�]�p�����@={�^�I>��@3���n,U��+ʞ��Ɨ� ��R<ԛ%pi0\�r�(�,�b�l�]V^_���iS�
�ӷY���i�Y�"J���ޝ͢%F��蔖�5m��ם�K�/LVX:�w��9Γf�KJ�#�[��>99!O}pmP�
��͕�6	��	�78���[�@�s���%��}$9ז	 ����(�����z�ƛli���5�V�.����| W��@��d@Pt���~�:��N�g��4�)Sk��`�	l���F�$m�t��p�&�H��#	�<xD��Κ,4vm���K?�m��3<��byqSTU�8������$�<g9����xXX��*�o� L��"�OO%Ac�z���7�T	<��#D�����. ��T�%@P6w�3`d������� '3���wz�5@���'�����$�(À�I����DI���I��x�G�M��qփ�r�;/Y�{YƓ�"�e�gqɜQz�7v��j��Wi�Nݨ�L��^�f�����R�j��[�'Ďz��>'ٛ�T	��؄T80��(l�qG5�v�B\&���7� ��y (
���L�|�*Y��a��s�vgĎ�ִ�`�8!�9���Aw�B���{N�8.�^���}Y��D��n�z{��A����-�<A?�o]\�۲�9M����q�x�V۵6��������AC7l$�a&�l���F�$���m*�>m��W=V�u ��<�������M�)��$!�3��G"���\��o�6h�.�z�m��C�l8���;~b 0K�(�Oz�D�7�T�0k���Ww��������I��ꢶ٤�H7'�co���j��#���@P��Z���
��� L�ʝg9,�7՚@O�>��y��l=
�{�Q1$��y$�ccX`�Y�nk���~��#��=�T��'�E��k{o�#n���k�n
*0��$t�v�"��HS3�:��7e�c�v	���@������ ف��R؞��ozt�̂ш�D6`�|�(�Y.�nܗ���S�8�\��Mhx.�x�������)�-t�p�ڢ������"M�yZ��O\���{�G��܄�, �������n"�l�A�٩�H$F]�U@$c�I2.��랷5'Z���3'>{p��PD2D?<���F������ld.5{�|I˾�A#<2H���"���4���k�6��X�W[>#^�UA#v^�}��Ն��d�"��H����xQ-�M��lÃ�슔I����dH8��S�rqX<H��j�H$n��$����^:'n�9S���^�Yvk�Y�ee�KdŶEG�5i�NoV��[gL~ʦ�/)�B8nO\4Kv١���ʆ �;�&S�E)?ywݍ^*��D'���㾀^�K�U
w|�Sd}p)�h�9n���f4z���{�\��k��\e�[�]�E0ݪ��o��T(R:�ɢnY VJZ�])˖�,�h�f}t�f�F����6��ZVpX�v:. 7�N�Y� �{�P��B�����r�L %��2��I9Y��ݽb\;���ә�m�)����,���
JWd^$Ѥ�0��{�?A�yz5�?_(\>�q>'4͇�YE���숅JI�.�SU�����}��=�����֧r��o���L�6�M��2�+6�����ܶ瓱�E.=q�̓=��L}�M֎�_J�E��h��3Y��( B5k�ϐ�lO����,h#�7���{-V�˹��~���ͽ�B&��k�a}���Z�>΢�{"O��NoJȺU���މwp�S���o��9vބ/�_7(m�MX��$'>�G�.��=�e<Ո�)e���;3�ӻou�����<�{~�/v��Y�s-X���*ݬ���S�3���N~�H,~#fays��������;U�k��:ڝ�n��>1kK��>u��ܗS-��c�K�����䬂��q(6���'e�U��'ѻ�1�3*3�;b�CS���+8s�0&y�}��������ya/mSe����c�u�m�{���L����π   ��,�Y9h��UT�U\h�hV��L��B�31b(���("��"�69@�#b�LA�E������J�
9jQ�f\pm�+���JV"�UJ����s)1��1��q�V!��A�J�")�P1T[B�[T�-����r��V儬�,DJ�1F��%���*[q��Y�rª6��L�D"�R,��
(�b������Ķ��T�*�VѰQK�R��-Q�[V��¨�ڂ�DDXˎW!�UUmGkH�r㔘�lL�(,�Q@YU�HҋUEAG,�c.Qb���0�5��T��m��2�cZ�$�U3,1!�LF�*8�JR�r�E����Tkw����{���זZڰoZ�� �w���8��2<�����#q+f�|O�ݴ��n�[[<l�ӎ�î�= �>.83mv�l���hm����ss�[�u�n�S�.��
��nV8��5���x�͕N�9KZ׎��=�>�n��/+j�պޜ�.ˉ��-�j^�|�	��mΎ�<k�k�Ö��C\\�p��mpQ�x��aܜq�����q��+��6ݶϬsN�90��h�=�r�۝yǳp��1���^��;�g�cesv�KƵr�q�7f� fˮ8�6��u��t̞����5y���Xӭ��؋r�x{'5W]!xyC�9���wI��a\���-�%���8�=�8�>���z��!qkv�ݮ�d�{sW=�p�Xu���q��l�����C�.��.�Pn�ӓ��O[���\����6�rv!7N;�x�W[vA���Y]�E��(ܾۜ���MO���ݫ�8z0/`���ۂ,lv���W���cpR�ι wn�aћM;�q;��x��Z����dl��Wl���s���W=�{�w;n��蓧m�W!�NƄ�cc<�6�ۑ����������!��M��n��<��4��kFB���Z�x�Ƹ�7.�wn�1�]��@xy6��'�.�����nŽJm+��]�8<[���0�0�ݗ�3�m4X��>|����=h����푇���`�ݺ�Y�n��l�m�Kwn��u�ϲj�m���\��h�O)��� ��{v�Gb�b�QG�۱�l^<玤92�G����-6�l�g��۵��ݍq�l�Ng);\c9��h\n#���v�ص֜or�I�h���=c����]]�-������=��;��ɸ�gz��n3f_l`<��.:���<��M���#�j�6��Ƈk�9�#����K��띄gla{pۍy�����{��G�m���������v���&n.���6���O&����+�Ս�p�JV��V���|�v�4+����9ҏ��euļO];y�װv��b�N_������h��h�u�1���/nnPfܘ�#��v�Onz׎�c��#���n 	-V�������y�sي�Qm����ڗ��7x��s���9 ��y��ݷ�Ѽ�{G�f��Ӻ뵐!��@�e�D����-A����w[��7�\�wó���#�Db�h��N�nV�Ev�e�A�;M���G3V�i���n�,H��q�ЯO�&����S�1�q/��=�^��
 >W4�C�=<�}�v�d��Yt$^��$����7�Èa	ٞ�I챘�tI�N� �Aܧ�I���$ӋLk!gc��Q6�d$Xa�)���cd�on�	5DH��C���I#:�$�ol�%�fCpeA�ę͛��Md��qv� ���D�u��&DN��Wپ��g�t.��(�
h�uneQ>$���mS��\<�fX��5��NJ��MI�T��\���5gW��3b�����۵ngێ����Vp��/nCS��v���[�������p�11��.�I5۝4 �ԞH+���A��/�5�G��@:������78���[�(�g��u����\��[��A��-��c�R�n+���l��2�˭6�D'rݼ��:��+W�Y���9��W��V-\8�P{+�$��Ρ@���F�� �Y�w�~��̲����œ���$>k�� w����{��_�5~�F��U]gl�ݡq����3<�r�zi�r�	(龚�|)�ܩP糧~l��s��z��7bIY�ۀ[J�H��StIL�Es���X��>���@ �����CR����e�@}�)-[H1҂�C9�:���=v-3q��g
��y�m��5����￟}p�ĸ��5�j�*�#k{f�A��$���yl�Kѥ@
k��\v4��g*���1'M�K@ۛh�e7�{��ȲN�v�|t�dH#+\B�Y��FN֙������)�M�]�D�3�>d����ӳ��Ɣ����{̊i���mg�VQ-;��*�����}%��o�ۏ<�-��x�]�j�rY��9j.���� ��ݪ�5OdH5�4�aD6� O��uvt0���ЃYݵ� u�I
 ��K��)G�Z��63&ȹ��`ͱ��X������$���Ư��-͢|�ʢ|N��� �Y}�@�&�QK8�؉D��V��]m���h�8��]��.�Qʼ�<v�wH��»��ne�!2D1�wn�� ���((�ʺd�r�:ܼ=�,^K�C�&�b�Lpڿ0�2C�)�T2����k�Y5/c�/4P ���H���|V�gkz@�^�T;��dp�M�r����kozE2]���2�֒	ɍ�$�V_uW��b�C�8��v��7���٫Թ�־���5�}9�J�'��{z H�K���3������TJ�v�MP&o;,@f[��� ΅�5���;�{Qք0�RTb� _M<�vܢو�"i�!���R�H��i�ц�@��k��u۴,������bږ��}�Dr���K�;�ۇ�\$ ���^j""!�<����Y㫞���b1ژ��7M��=�ߟ�{�Mv�^�~}��b:߻P Qw�/���(��H@X2b�I>&������X�C�����f��.�k9j�s<��3/�h�.��}pk$n�
�x��1�*��f �Fk�U�T	 ���ejY�u.w�����^�)�@�ܐ��i����1 �ڊ�d�fb=79�����\�'ē�ݪ� ���G�\�ܵ�7[4<O��E�H�C�0��K�T�����W�2�qs�^�*�A����x���R�Lwm�rC;1�k��CuxB
��%�2�}}D�#m���3���m�	>��:gu�m���;x
��sZ!o���'�+(�c�&<�#�lt�6��{[\�y��d],6-պ��`�8���٣�l�K���ׄ��vݪW�p��:���Q�#�u\���TP=4�nƁp��Q�֓��o�BB�η;����۝=F볗L�sj���}w �ң���k�őЗz8	+!���JN�)���r�(P�ĻQl�K�nw �GX�ٷA�DXg��
�#�1մu��u����ThR�H�u��y�ŜH1u����F�\1�z��A��H m���T&l���=�k�w��(���	@a&�l�.vXV�L+�vF�U�x�M��Р��%�zd>\���Э�C�����jo��3�!�N�㛝r�;.S��H���� j�ȒDhڿ1Y,�h�NWe.��Y�$�ݽt(�|M��$��t�)��V�r���X9o���L6�2\0����H�v�zF�)�����O^����%� #~����i�Kb��m�r���͌�rz��^c�g�u����$Mi�6�P'􈒦\���!�1 È��z��h�fw H$e�uW�z��(���������"��D���4ڄ�%�$l�uP$����#���A/Ɨ�kU+b,�ej�z��1��(�R�A�1F�u�t���<�Sε-���]B���
^Go\��shؔw��!@|q�.�����P�kH|}K���9wb���f�0�"�U@�s��A ���K�>t�'3���
�o��P��"I�.���>�ƭ�Âh�b@3�u�]�s=��D�zvC �|.�v��>���f�/+8T�2��^��i����PaCF���{U�A'w;kկ�y
��J�F��� 
�s� �ܒ5��t�q��oM�a!��(eBTe����y��^��:w�6N�2k�[{����R�A8HC8�Ωd�}�@E�vȭ��%��yE.wA��گE��#�C�b��!ڽ�Iɮ��n���[y�@�oo���IwW.y���M�q��m7����$M��ׅOx惓�w�vR�x���d������Sf�xN���&��Xj�g�t0]7�	��J���-�TQ�sPy/qo]�й�܍�:���U���W�{}�G�ïM4Z,"�UFK���D�JӮ�� �;�I$�_mQ>�U��cW8Ќ���1n�l�&�F�=�t(��$:JO?8	S9�V�^J��#�m*y��iԞV��c�T�m8��I��2`r48��۸6�M����sl�{@��M8�H��*Sl+��)��%�o ���~H���H >r���~��h��gzt�H;��B�P�)7�N��9�iH,Kv�hہ�3Q]0�wĂI��T	$b�L��K�l��+
o4�Bo,���P�=�(�sU��#%)<�S�u:	#�7hW�΋�$��&[h2\1_uJ�C�n{�BG�h G��k�w-���κ0�B��q�m8]�Λ��!άY���m�y$ۡ���������{��N��x+$�f���6*]��P���Jښ ��l�EfgMx��.u�yo��^S�K�>�<�h $��_
�y�dt�T�C�?4��pXm��!Pb-��i���b��â��uE�h-�������m8A�8;�tO�u��3;9/�_�Hm�sq}J��w�A�g�sA���pl�{UӀ�nX��ϡ�\�۞��>'��yo�I��T}���#K���y�Z(��s���%�!�sv(�;}�4A��K����b;�Z�����xd	��T	ݲ��DҚ;5�ҕ���c�2'3"��A{�B��3��vw;��B�vFlG8h��Ɇ���uD��f�O�B���>%�;2	�;��T$�{��ɜ���}��|kW��yk��"^_jg.E:nv˖0f��6v����Q�#/�v���q)�b�6ƒ��'��ƾHg����Ĺ���B�H�X8��3�F�qk�v��z�]���Q����+�0��D�ۮ�#Vv������>�����v	8��v���s���Y:�B�q��m�sC�M���c[�݃���s��d�������[���l�]"��v[����=����$�:�!]�o��8ls�y�Q��gF�w�l��8�ٶ�]��kv�8��snD�#W!P�m/n9C�����σ��	�w��ߟ���j�0[kxs(fgH�A���K��t��7�.�������f-��`�>ɭ�s�>�ӇZ&f�#�3��I ��uxP>!�w����e���:bpu�b ��M�5=w�D��w3:|z�a*s�p�@���O�7��T@T-�P�P1�`ă��C34��Yd�Q=�@ ��͡@��xu��nmT����e��P���^.�v2�J�j�$(�DzmX:<߷n�h$tf�
�>7��@P$�Gb]�t_
�2�x��� ���A[(X*z��ٜ�\;cc9k$�gp��V����Ͽ����zŶ w���Q �os6��A;QؤX{�?{�K��`Uq>K�@>��{����6���6��`��D p��]�v��#i^�V�/�We�;��]��n����S<NN�}))j�0Ï���;�o���f�m��S�g@�Jn gz�,\F� ��3��H'j;�5��\�����A+5�fi�K��;�uD��A$5Nc�]�҉q]�'�3hP$�Gb��n�l�����[xz��3Y=WT	=Qط�+�*G�Hh��\��� �Ѫ@��)C��@��9�j}���Ml���V͓#)Q�g<O�9Qؤ����E��z��z����J��ndcj��K�zZ��9�z�N.z��=��6�2k+���C��<W����.�95�^��0�����H��|kԃ�z���=羡�Jo�*���x�E����67�pH��(@�y�=ޢF�̉�$��ު� Mc�^��m�dޙ�8nB���2bv$[y�@�IC�[o��-$˂9m2=�T��E�=cJ]���Ԩ^x��ٛ&���yT%�JB���=�̛��R@�>c��ry����� ����K���$�,�"�zBk�:�Z�w ��2�3��k�
��K�
��M�������|Rg�xc���yK��P�:���A��D�I�\/P_E\�&���halk��Տ�M��̌���E��V��A�p�F�j�|A�u�F��p��+���2�Ax�{s�극Fk]"[S��2o�.��eW�G)�����1Iw����C�D�-C���m����<1�3{seΨ��Xк�!-�u-�ȹu*vpb�Gtg��s�n�,��k&�gcB�Fw�cf6ݗ$H:j��+����������wOP�gEv�c<��|�#B�-3�Wi��F�SX�P��D�������7o�Qz�U�Y[���7p8���}�]Hs��$̺,����X���z�B�9ѹ��λ��-dKE�%YX�jѻ��H'��|����I����U+c�_#7:-��9�x�G9�����l5v|��Pt��A��]�䮩3`3�5���O���e��""�L�<����uV&�\��jȫ����gW5yy�K3(����.�A�{ė���F�Ѷ��w�]����{�N&�#�]6wucuݯ'f�kC��s�KxB�h%r�a��5#�3��e,����k��e�
-.�R�w-���gE���22�P��n�f�?y��~x���^�F2�(����,�TT�hѱ���#�Ge��e�VUbFZ�CR���V҆R�*H��,*�
�2����QD-	TED����"�"�"�,���Lq�+2�,ik���m�iYRYiZ��.3%�X*����J�YZ%���Ym*VڍB��`Tr��TA�QX6�1�\�Z�-�[l�ٌ��Q�UƵ��Kb��fULn&��#1�%b�ڢ\a�j*�ܶ
�Z2ڭ�)����)YE�b8\m��
50�bT­*L�Ua�jZ�ʗ[hTZ�W-���Uť����.�d���C.fe�µ���6�%,���bR����b�!ijRԩem+�*��l���-�e�����VԶ�ZcrKKF��r¸���Fҍ--���5��k
#ZQ��2�jإ���"�כ�AF*܉�3/z��6��P.u�=��Ƴp�OW^����� )��� �gl�*�����n�I�cm�"N $�5�0�w3:�FN�nK�a�F��Z��Fm�U|H}'�&;�lp���~�n��l�[�����`6��/��ی"v���콸�l��]���;{a@��0 �����'Ǯ���  >}'����̥�ֳS;����>�z	 ��ު$P{����B���vkz�w�締q����fv��oovhM�gW�r�u�˚��7���'�%� N��}��(��R{9��)a�u��$/�z�/s:�Dv��8�Q�8�L=�B�zw�b�
��h	'z�hP�U��"	0�>�s�>T��������pj�8�(�@z�:_��[&e�=T�k�`�<d�)<��бy��? ��U�B�g�Qj�H��ТO�鵃n�m�E������ *s��P����	�ɩ��6M�U{��pX�C�n->˧F����Z�ێ9�%�3�U���˂�z7�b ��pX��٫گI��ʀ�/@�����^��J4�D��Π(��J	����Ω�Q�P�ݽ��[�:	��y�@�H���#���1J�T���m�@��������j��oP��O�ܖH���ʛ���O�:�k��5� �FC,Bpߠ6��]F��ZE^>�$w[B�"���Iu�N>�iS's!�|����GL�z����p�T�2[�gĝoݵ��[�/�
����>%��S��H{s�KW�s���t}·��)�h���MB*#٨%�}��8��HXܨ2��5g�ѺR�����zͥ�Mǋ����Fk�.�
�H��6�N�ii������r��xݷE���wf��7h�:�M6qu�U��W]�@;�����U5�8�{��q�y��%����\�q��;Ҝ��5����Ǜ�gR��u�lf1�õ��P��ҕ��n� a�.�Qf�6�-��p�u#�9:�i��ǜ��m�Nܙ�7���%�m��g:����[;�ۭu�*���ӌ^�]k���`�s������mGojݜX�z{{ v�@0½�<�a� � ��/6��N��k( ��$2��[�߹#�ۙ�}�g��7ܠ���mi��_�o�P�뗅k���^���ӈ q]/A��I�|�]1�U�ɚ�u�(��J	���9�,[{�@		�NA����>�r� )��J��`�H�N5�x��.�[�U��|0{&� ���
�N9��m�O��"6^�x�Q�+-�=� O�v�����{y�K6$I�=��Ξ�K1m� ���N9�K�v����~�^��{��H�i�]�/�PB��6�*\�����hذu1��Mè�������
�7k��m�pU ~�@ �y*�����R�j"=JnbA ��ݡ@E�vڀKP�fbA{�r(<y�u�Z����tw�2�m���⥇�+�u&.����'��3�yw<3��tS�]�.��P�kGr�E��V  �}ʐ�<�t����筜��$L�a��8��P}[�+Āw3:��v��|�lfÉ/��
�s�K� ��T��3lц�	�:{j������$����s�6�᫯"����u���A��}C�H�l�j	��w�Av�_͹��P�d2&����O�m�Ux��� L�P�����#+M5��T����g�:d��[���F՗hyMs������P�Ǡ8fz3���$���
 r��)?۞��uy�)c�淥
��ݡG��`��f	IC�&�*mEIW0�[��Ξ��;ovh�5u�H'��owo�Kޗ\H���KP�fbK�Dt��A%oݕPg^Yu6U�|�W)bPN�S���]��ڲ��ɣ�4�s�{W����%<����/�F
�bY������|��KR��F��+5k�K�� =�~���H��6�fn1�VMvW\��'EI��\��xڤ(
�r�Qw��2�v#u�fz�+�|"�l�F(&�x�Բ	���܈�
�_SH��^� R���96�,�M��X�9�㭇9���!·1Y�:+���� �/j��ݵ�1%8�Q��=�X0�&`��Ǧ�j�����`��Y}�^*gq�ͭX;�6�=@��o"I[o 6�2�ЋqDn�R�>^��y�C�<��r�h(��@;�dD�us�E�.�&����4a�H˾��+FN1sY�g���ȟEe�U��q��� ��S�&]!� �n��s�P Pq�ڌz��g5�s{X��Gb�pL��w�V�����0 �6f�Iy�.��I@���ͫIԵ0kdMS���X,�����g?��O�5�a�,$���j�P |:?r�J��D���@>��`O�̽ڠ	$��
�	�����������:[���tH�`Ծ�<;�۫��X^�Nxё��w}�w������/�5m! ���� �E����R����@R�� 6�d��,�� %@��uz���3S+�der�� �H׻T�8�ʕ
�5_] �:�E=�J�����L��&� �g�a ���Q���Ozv�nr�2��}�}@| q�m.�/&L� 1U�g�c���]�Pԗ�P�8�%@P���W�)�Dl�U|"�<i����Bѻ5b���	Y	�܀,�$� w��J���xg�9#n�d���&����B�+�R�]�:^$v�C����~�Oړ�@Fn�<�$	Ɂc�,�[�.�@��;�r�I9��&K>ߦ�l�㣙n�lZ6�nݱ�3�8�7���r�'n�y{�0��v���i�[=��n�x5�h�s�������q�u՛[�9k����̜����\�-��&���{A�c\��3����{v���z�����=gpӏ@���Sd��cc��w�����vJ�d�&�;��)����9�ln�g0�x\���$��g<���	�5��;�;RB��d�{���e��W2�!0����d����c1���$�{/:���N��2n2s��U��^'���^u
TL$a`Aa9;�kH�-�^
Gܦ�( ;��@P�xD����g����29���-�!�Ms��I ��d�H'�wu�:���$�{�:�	޷�I���0Ȅӄ�����q��a�M�� ��mQ���xg��ޫ{����Wя� {;z{5U�!7��2\�N3B$��}�F3�\��_���T	���>$y}�!N}.�O��A���C��\"��v�����Y��M�=�vŝkSs��w������=��A�.溈$�q��$��ު1�F�Z�X̐d�H�H�H���&�E'��鿺� ,�^Н>c��xE�L���������W(�飠�{�q�+Ā�-u�y>��b���4�m��擷�+׹]*l�K�]�h��� ;�em�E�g�D*�	M@*aD��lT�I5��4|��3փ�tu��s�0�$�y}�FF3��&""D���W^�b�|rv&@D�H��T	$��w<##�uU��Lc|d��-iq�Bi��Ԫ���rF���Q�m�W�V�f� 
�s�����m��w�#���W
+�4n����Û�g+���]�vɠ��Y��c��	����	� ���ƥ��D�r�h�A����յ����%��:A�ސ��h�p�A��rQ��a��_�gn��#�A U�uW��{y�Ssr�uR+�G'��E��0!�f"2����}@P:9�H *X[��ޚ$c{ok��h&�j�E����q4��{;�i���-�W��ͨ�.7*���n���iօ�L�j��AG7Ԕ(��Ϊ��O<�#P8R��9��f�F�b�OY ��W���͡D��xs�m>���؇d���Р$[���a�b!�MW���UV�HX7��-��b��S萠s�*ܽ�h|u�u$��􉈅-4
I� �i۵+��Wn��bs�j�ODk��x������}ҥ��a�p��ڢA&��dQ;\�Ɏ�&��,ͥ���M*(>s�W���E��SZ,/��0U2>�9��ƈnjp�Aμ�r�b��{	�������9�|�Ƒi1�2�Gi_!>;B&Nʦ���d�f�uP ��L�h�6Y��*��^T،��x����
���>$/7:�&`���8��d�)�%I&v��v	c�%y�M[���G����b֕�x��o��B{�od* ������]J����{2E[8�)@=@�<�B�s�&�0�A�S� ���M i��s�nV5�Gg_UH��'����Ԡ��[��]/�JF�r9Ci���b�]e�y�����8���͸๼���Tzx���ѽ� �a�b!�p&���A')^�����+/�1d�Q���9ە^#�/��#c'a�d�i�$k��d���=�n�܋ޤ �[�@'�U|wU���]m����^!6`�2bD���Mof�x������zDU��:��I>'3s����f�"�~�iɐc�����bM� I�[��+w:�ng-����{q@`j|H���`���1�S޼�����f�Q�n'ۑ<��{{�@�H9��B�|�߼Z�^�o�z�ñ��u,�W��݉�\�&��ـ��У������אd�Q���J��<����"�t<c�+4I��])��u����|���:��W3|���\\A+3^v�P�#�Mr{����+�������>�|5�L~� ����M�++�|˫  �V�f�
η8h˸�Jz�<$�����x9W���cf�,L��]F�5����ߝ����~7;�@�y���d��x�z˼�@������*Q���%�:�241ڳx/�R�Cm��[[iӼӽ�ڈ�3����%��_+"�v����g3��t�MD��˕jq�+�5
��9g]plx�wKD��B���:J�\��~/�{��9Fu���d9�<=d~�?N�J�}6 ��ۚ�����mc't�`����ʲ`�&�
��8���㇔a
��t�R旘��������1,�̻�p5�/\B'_׼w���uᎥ��S7ݛu�2��������
����)�7�����)�l�����H�;���4����i�[��2�+�]�Z���75Q�FG����;�	�Bi�LO�n��f�V���(U޽=my.r��n�7�l�;�b��t9�����L�EyQ��j�-`dh��\�t��,rtz�{�/���v9�-����T%���Lo �[���|;��U��8N��Qc-r3��Um�>�d҈�B�7�6�y��d��w���oLW񡵅^=��4��ë����J��K-kFZYF�P��խ�m^32%���Ʃh��iV#mDP���(�b[iKB��\�rؖ5�J���%�s&Z`3"� Ѩ��b"F�diJ��-�J�Ye�-R�b"����R�TlZ�J2�-��J�1�b�KV��ک\�*�"ѥ*��G0�b֪.eƢ�ֱiVV�%�-(5���H�Z(�b����X��5m�EFKj����Z�m-Z�+UD�5\���RҢ�mJZ�SDīR��X�P�Q��ڨ�%\k(��Q�c-�JUh�ih�j�J¨��Q�E"�Z5�L�Q�5����FUAKJ%Fڊ(���8��)����V��ţlKETBҪ�2��q�։iX4��*���Z*�j,(��7�1lQe`��j)YYl��D�RPh��cl���T�1*���ym���ܩ���y���� pn3�&�؞w��ϥ��]����N�!�Z�v:�$Y-��7�jݱ��pe�q�ql�a����u�1��0t�Y�;L�,u.knx�4`��G<�������s�[p6�p��M̂[Wn�ۂƔ��h���.�1u"���f��N��:�n� �gn�u���ùn;ko@E�����a6�O�� V�z��8"�ۇHq� z�}pח��E�e�]�+�6|�[vw���i�i,�a���nۣ=@�.]�>��@���,\�9N(V��kn���x^Y�3{y�]�/.^��LmO����Y�v�c�D`�6�^��:j콍�:��;9n:L�lxγ��dKcv4�&��s��۞9�+����hW��MSY�:4z����u�=���4��#nn�>�G�nqWO�]�6%h�����u�BvV�ceeEŷ��\`��gC1��ȇ8���;X���ގ�m�&���b��5���H`89����c�)t��%�+���襃�K��C�;�hY;^s�u<(b��v�+�r�g>�9��'�I�t\qKľ�ݹ�a����VZ�r��+6�˹"h�}��ێ�vq�띸{Z;�S��m�z�:�#nm�q�����2�uǐˮ�]n�V�6�;/gyj첕��=��pg�,��2qv�.F;譬��ێ\7�-�����v���9v���z��$�uθ9"���;r6���y��ѤA][���s����n��4u�ۄ`��m�φ��ek�n��Nq v�v�s���)�r�1�����c�3a��Sݳ�]���t���� #0��[�Ѻ��p�N!g��sl<��x��5�ov��zM�	�^v����L�N�kW�)�mf
x��k�ud6���q�6���q���!Ρ�Bn,p��p8#��9`�ٸS������[:�5�.���^���͒�;r�]��v���]�G[�*g����!5̧;�ǭ��[�ݰWJ��[u����%����Tr��������n�����5���Wt&^:���v[���n}{v�8NY��������\-���mmڇ<�w`���{r�t��p�dƫ�.6���t�?s����;1�<��6q��n�5ڠ�s�=���Zq�r�ab2��ō#���n�'��,�Z�]K��<�m�'v:D���ٍ�0��ڃ��;nqg��	������g���q�=0A'�s��>$��t�=ý�;S��p�H$}���@�3�I0Zn����>4�k��Ei޾��G��HoӒ�>��<�P�r�^M�%��~�A�a�
hOL�UI�3j�"���`��n����2����
'I����x�À�P�s@ԭ���������^ ��͚'�)_!U]=�Fn���u�my�-?(i �ں�	;J�@�V��W�v!S�S��A����Hʋ�&Ww(�96���(��t�\�z���&2�b�W���9I6��z�tм��0b��pv�H;��TI$��@��-���OnP���ꢨk��!�PY*'�qOH�@���Q|��H��Q��u�8���8H��\�a�w��{�7�q�CJ'=J�Y�b��w]�I�w��B�k�*m��Z
��e�yݾ�> 
�s�x�2��O��9�4��/�W�ٙ�I0Km"Q٭�H9J�	v�T��7��	�$�^uz�)_)'��&9sbɑyN�z�d�ت��ʡW&Ĩ�+|t��=<�����ʽ��$��N�Wo,�D8.AC%�R�P��ٲ9�M
�Qo�h�UU^ �E��y��@ա�c1��s��`L��u�������,��;=1v1ȝ�h���o`���e���=�-���pͫ�@��{"	 �y��@�����ٺ� ���R>�z-�`�6�C[=yT&k�|�=�M����E�A���U�}9���͒z�Ϯ�T�|ؙ r�Q �)��I���9��ڝ�R�n����[���A�s�W��:� sk�E~�;����,9Ϝ�zђn.f�d"��mwv��lF�=�
��k��k�z{L�u�V��@��Ϊ�38��m�A�f��g62{�(+�V(
�;iBs��;�&��BfB$u��l-�&[&&����^�}y�F�l]I'�<�O�{��H9��B�S�O�<T��6��{z_kX�x����bb�<nz4��ϭ�i2�H�!�$0^p4�L��ݔ T�<�P�~�(���wx�yۇh�{��G'��@��L��ڹ��ϴD�
I0��|O��v��6�V��W�*�t�t:��ٯ�V<L��U7�%@|�yU!@�N�;�Kg:Xڙj� �{���6�i�P��J@�O��������b/����y�J���������0J��S���'�.�y�q\�Xy��*�\{Y<�z��W0k�U?.x�6�qkEF6��|n�ʯl� ��+�U���N8�}�T�s��a�^SGf���#)^Ȇ��-�$Fwmz�e�P�Q|��)��Q������Lr��1�� ��7Zx��6��ٖ�<^����u�6:�J"�����[E����x���$�|�*B��~;C+_��*��}= N��P��Y��b��l�4i���P��ǚ���A �g^m
�7Q|���Wu,��Ӻ����rI0[�S#~ܚC�(D_��U =��X�=:�^������Oe�P�|n�����C@bj�}w#H!�DC68� ���P/�E;ܩo�&ǴP���_;�p�$qbc	L�*�?D>�{�P�l�<�Ҫ�7��
s��:�{^蚱�¶d�n�#��hӳ<?E}�j����_L�v��=��[y�z;qꄫ��X.zb�KZ���ew�LpEP�X��l��L�Gs�N�7�x�X���I�Т�{I��]�ҏ&�i��a�z3�UMn��=�<�3����V���Y�G� ��^{n|��3t�kχY�Ǎ[��ŻX{���6�꽴s�u��n�0V���/�{��{�n�c�x8]>*#��J�������v#�XFD�9.�;��8g����A'N���"�˵÷YX��9�:�r�;;��k7[Kj�S6x���0� ْ��-�U÷�E0�a�)�Ǧ��Q��+ك�A"�j��H�r�5��QӔ(	Qz����xh��0TC"c_uQ �fov�ܛ��@�FT_)$x�yݵ@�qԶ��I�;�6.��k���vL8�Sd�����'�AQy��έt���`ڋ�$��$d�9 ��-�)�>1�w�}�Mx��	�q�>��n�� ��s��G3|��ɢ�$ԻN�h���&�b�8�.~�6�2�+ >/:���'պDJ����~ ������ؼ���0T�Nr��f"�Ջl=�&�ԛf=l@Vv6����[�[���7[S?ȁ�XN>REn��E���9� �����{ݞ|�DD{�r���9R�D�!�I�U|V��Fuxf�HP�h���u�ԷYN���6ʙ����Dꑕ�5�o�~�l�@Ҝ�����̱�C�G��������{:�%$@�v��DY�3�Q l�%�d��c����8�7��$6*)�w]� �ͥ4|	)��ּ{s��C� �f����9���\B
 [�LЃ�B�T��j�� y��""�w�,�Q	��	%[w�c֖�3�"�n	LҠ�[wN��K�iW�|�`��<NC���'��w`|�;]}D ,���]u����}(�43K��C!H���ݏS��u�-��nx�\ҧGk=�֍t������^���t�s�wǷ�.��#����|?|�o�fF����Xhŭ�L�I�2���?l�`���&D֍g����5&��3�����~ <�u@ 1���$��4�;<ef3�5y~���L�Ɉ����4��SG��z�� A�ՙ����%��z�
�-�������1�8oRT-�<-�B����z>�5�m�lo�\{��=�AZ֊��	�m�<I>��k�A$˷�7<�IA�7	"a�F�[3�yQ՝�/,�q��h���F^�\�{Ú�T���}�ѱ��aġ2T6�r��al��4�K�Vvm]��[$[PS7 .~�u_ ��~� �F?O4˔�m(��_EVr���W��)��p^'<�s ��n���Ĩ�k��\{u�����Sm��J�b�	2������ �^�]�A7�}���+|�� ���Js�� �OZg~���~{}=��G[!���h�-n���|2�:�+ A�{��P}5�)�jg��:�s=�Ǿ ��ꨰ���Wo��^�����@ 1���=�^�]�3�&!D8k�Uy-Uݗ�0LU�n�DF�Y�	��#�ofmݠ3�f��m���k��z��W���n�Y��J��_FA%/IV,$2i��$����'�-�T�}�6�Ӣ��F��ﶰ�]��8��p�TdR�}��H�ꈟ$��;)�
6����o]� 3v��7�TM�R�[�7�^��D_�$k��Tx�.�ӕ��Q�
k��
0d�-KPI)�&TOY� �n�+G"�R��Cc����߿�����c��f$��y���> ��ڵ`Z���دV9[茰|��Ff���f�8��a�%A1�	6�C+|*�ۥ �"��j����3��e�����"c��1�z�����f!����'�{z���|3�����j'�tj�q~�t�H""�3�Ҳ���~�S��	���sWƳ���뼣����
���� @}��]DP�o�K�x����C����p�%D���PK��j��m�;_+۰w�uV��]Q [w��^E��eЬ���F�B��pF�k�c���t#o۝��y�n_&ǆ���{�Յ�}K���e{��a��(:�37EffQ=�v�r:'LCq�y�p[vwnv�]����WAnV��l�w'��m�V�<[n��z�<SF�C�g	�����a���iy��և��8�����T��n���W��'y1���K�s������v�պ��.ݬ�[���v�m�qû9Ϡ�#����zM��WU�I���6^Nڳ[�B r[�����'FK���O�x�oH����=:�;i��8ܼ�q�kqŭ�h��ӽ���\�h�y�a�<A3����5ؒV���ZA"q^�)��m�7�r���S��u`�z�nҲ5�k�7^L9P�f+0 0��u�	�-�֡7w:��$ ���H�/���?��6�E�^}Qk=��l$�IPLQͪ���`_7@ ���"��L{�^^�X;튤RH���&}�<Ɉ/��O�^Q?G��1��ᛤ�aOר��'�o�� Y�����^���~؆�9�[�� ���%�pI�-�;I�%[��vJ�yU���}W��[��5����	��c��6rrN�6n�(s)������@�<��\�Ip��
]ms
��L9^�P���ڂ��$��XV?) V�{�
��'�.�$#_��7�N����7�^KC�$m1N]h��}��THm�{��Xv +m���twb6�F�;��l�ʞ��ж箝�_���y�T�J3*�6�w�
rز��8��
ú�t8j�s��U��]Wu�f�2G}�G� ��o�|�_v��A55/�����?F}��ɇ(���s�2u�A ���j����#��~�ϯ�uo� cy�� �2����+�16�I����!�UC�ߠ��w>��mǾ@ ��ۻH�;]�7�r�ꊈ�^n�ޒi%�#���ق�|���'��~>�W����X߱�$�#3�n�- c��J���D���b�QE���<�����t�M
�6��뭲��.k��|�wt�z�e�iA0�.)<8��ph�z���X <�u_r�ʛ��\�'/�y���� F��ݫs'��C�9��*�J�~������g���N����YݵV <�t� ��y�d�*����F;W�hr�)��#\�.d !�׫�@U^o<����d��*�.���I(�������D���3������5ĵ']oT�f���r5wO,�7w+�0��"m���T��[9{&���<��=�L�*mt�+kŹ9���Er�f���˚x�wي-��c�6氏{iJ$���G�a��i��56��W����cÛ�B�P��rf�z{���vl�V�ډ�[�/�p�}DS��o{v��fp}T�y7�f1�|�����L�}�E�x3�=]�)��"ns�yu��\��Gm�_v�3�f�vk]V	閞F�
��ކ��0���mI��~��mc�U�B�k>K�3��&���<F�˼}+M��q���8�ɘq�N�`���ҏXl
��א��=,�Z(�WS�UV���u1�3h�2AP/wEK��ŗ}�n�k��M㞺WIT���::��8ϻq0+�zj9�������3ս+(ukV�m餄�B�u���#�Y��}Ԗ76!�8���w}4�pE̳��y��V���й�_��͇\�{�o̝����zÂ̾�l��{ƴ�j��}�1�{��X�V�2�'���υ�m���=��;�Z���@U�󳹾����ڶ7w��TB�4��V>kI�Y�y��Z���V��7T�p��ac;�����G�I����;�.��Iڽ�O+sBo���~��vo�Q��AJ-B��sݽ:�-'���`_M���V}���v��e�8�L9�a�ǧ���|�:{]��)�=i[���y�N�(׵.7JOqؐ�'˭Lf_ܗs\	W����Vx[�HG�e��j��,j���bP�=J&Z��
%��J�(���ki��TYEZ���3Z
P�����j��b��m���1UUm����Kh�P��XԲ�eb�Ѷ���hV�h�PZ��kj��bX�E��̸e�UYP��ɌiJ��W-�9�U���j�eDJ%ڣ���h��+UA*�U��ŕR�[J2�V�Th�E�lZ֔�pp+jҖTB�5��F�*,T�Ѣ65�[mm�KILnU��e��*R��Z�Z؍mh�m���VV�R���"2��A*�YJ����Kf\�[[�"��E���E�jQP�Ԫ6����̵m��mmm�R�����-W1�ն��Y[j�Z���ij�V�3-UŔ*�PD*ܹ�+/�">!cyM��׻�Y <�t�8�y0��9Nb��<��z��m����j��H���H�n��Ź�������ͻ���c�`I*	�) �j�hA�|�%Wr�ɹ�a�H"�f�DDR����;p�;�*��T`m�-"�4�)����r��ۢv��VQ`ء8�ݬ���w�����*!��R���\�n�]� L�~� �۾n!r��_�=�ywd �9��3j�C�$ja�Q�<�H ��N�WQT�e�=�Y ��uH �|ߐ�Nn�g�Ú��=�Bl���c�TG��B 0/_�����=�/�Yv�@|c��J����o�N��49	���U�����w�Ӥx���x�3���>�޷�>�'{���=&y��3�.�A�a"C�u�gl�v�*�<������]���n�k����7|�>��jX4wS|
��b�L��;��r�f7�����IK�U��ys	�8�e<LP>i 7��ڨ�>��b��A�v?R@|����� 2{��:����Zy�Fgm�b���t�K�Wn����7b�Ӽ�ʺ1Ó����jM�6�a�l�;wcS�`D�	�8$ں�h@�q��3;���=
�T�{0מ�_* @}��7�V�Q3��8/�^S��wi%�:+#�}ԥκ ����fomڲ�{�]�n�b�S�6f�H8�0H԰����lB@��r@D�L˻�������, >��� 37���\�X�&�l��>������y��]ߏ��APe�Hwn�� $k�毷�rք\p>������C��m��eTQ���v fm)�������@*�~@ �YݷQ�g?E�=�Fb�H�;94���8��9����E�/6ym��k�����S/qZ~L���'/]6((��n��TN�hCo³�Z�^؊=�[o�N10��N�y9��k�Pn��8-����
O5BN4�c�y�i-x5�+�n��y����\<��t&ֽ&����	���|�;��wJ[�<q�<Rp�'��1 ��7 ��Y��/m�6:�ͬlN���5�;Wn�{oG/f#�#�\O\�L�>�Vp��;/Qt#vwx�����,�뵱�	ġ�ЯOb��ӫӼTg#\�zv�`�q{ [uue	�-�t���5s�Fa�O~�~�C�!3	�b��Rc%H�U��To�@�'�Q+&i��O!.i��zI��f��ѿl�8D�I��4���W�D�d��0�'g#`��� Y��w`|5�s� A�R��o��wF�<� )4J9�^8Xϒ;ϣ2�x��SB $�
�T�v�Vr��8�@|m��ݐi�ξ��dͪ�n	n[�a5H�W>���c^ 	�H <�uH >V��p^�׫�_]�s%sP�!�	��]W���T�@��	�t=ؾC�� ��M��~$��:*�A%q���"��b3�)m��h�2���6�<�M۞Ҩņu��ն��3�3`&�fbI����i�̌���@���]�uQ�e��ݐv<��K�;��0��1QH�7��>�O��[B_1������͛��)�ǧZ�g�7ޞ�|g��è��|�9|��u1�zN�+8F~"��N̛���Ƒ7u�Q�d�I���~L�l.qO��X��b�ĀL���H']]'@D`_?}  {[����߯	 ���+�" ��o�eu%)�a��.�ה��^��QgD���"/�]|��7x�G����fʹ>�WR�X���t'x�a9`�dD�|�es����vl�>�Oڇ���S>ҩ�[w�� ����뿬��{���ʤ�lY,�6��^;⛏-��qZ^����0G� ��}!B��*����&c�~��w��� ��DD��w`VdhB��7us�R� 7z܄���2�0� �iki%�9��#6�n�Z�q�wΏ�@|����H���m�~$n�R{*�P����h����IL�d�S����3|�x ��䃢@�W{��l�Y|����h���]�'���Vz�m�.��#:무gH70g�Ͷ�Ơ�[�{7|���cZ��5�Ͻto��i�kw�� �Ff�]�'��#��	�R	�W�93�ί.PDp]�H �u�uݤ ��?:��wo����9����PQ3�&H��Wǲ�n��@|�:�<Sj�f���6ɍ��ksN	&@[ݝtI'n/����<��v���[����gf�ʦM���]�N�Jw���H=+Ӯ�淓��1�`�
����	D�Z	q9Ʋ��H �o���"�n<�ԃ`�w}�c��,o�����u��5�!�1�uH6��:��^�g�W��7��H��f�u�E�7'8�D ���rj��ȍ	!�se��a@A�(����Q �6� |�#��\��0Ψ��;A$of�ڲ �9�}A������)�b�`^����|&N	(7���� ۓ�TE�|:�͙�ʬ"����{P����'Y�[}{����#���t.OF�u��yۗK�=���O>�7��u1�c �]���O6�;ɉ2���eѰ��8��)C���u՞� dǤU�wۼLIf &�]w` �ǚU�|? +�f~pe�_�X���8<{`�Khuc��v�n.��'��&�>>��d�F�}�{{2�� ��3�h@ ,w����+7#=�$� �#���H�y��)��88.�\��g43ӳw��Xz�v�5 �^g:� ��|? )��_QGF�����y�le��DB-������4���@ �/G@ �R���O^TF�i�Ψ��X��/fK��ClQ�-s�}*�5����_��tDF�y_M��~H"fom��cD8��N��"]W:�����#P�0�1�,�j����ڰ-t�f������O�[�۪c����r@����(�q�+O�u�8S�ٝ��\�P�z��by�u�^ϫ���۰Ϋ��V;X	L���k����j�{��1D6l2O����y�T&�F�G�N�7��F��+w�������n<�q<�3�$�&K��nN���{z4�n�Tݛ]���7ik���{`2=�܊����q��E�vu�s�dյI����wof���.�kq�n�f�囌���F7n]�;�u�>$��['OaEՏ�OojtV�뮺��QVz:99/%��z5zt��k<�a�r����//N���vj�aTu��KV�;u���ߟ���P8��L��4| d�����v�g#�Лڂ��O$�p~@etYNf$9	q?U#���@����]�iV;��[�X�h�C{� '�ͲĤ����z�oq>�s���9��
%�2&�p����X _���������8��Afnuѱr\�$D#
l�ERZ�z1�?X�7��R�3d���'e��D73���<�w1�r���"8q��$�<�a�a�Ip�
:w�Š ��,RX.z��,zr��gnY�$�Hwvuڲ��]Q�{�����j<*�;���l����\'�69�s�u�҅tv:����(��0�㹡��-��3��S�#� ��ڿ�	��]R��檺D�ԳEŽ�L��^���Z^��\�@��)�v�H��*��qO���h��I�]����M�V:�X���=�-g6	�� ʿv�bm$)�)T���"y-�/��ڍ�-4Ǐ�|�.�ͻ��Ҡ V�����7��U�˿|I����y0�!�K�����˿� /����D5N+
��t_���� �^g]��#�������C�R9M��$k;���N�ҫ@ �˺��#K�~���&]�]��#�0;����h5�4pl��1�ꃋ� ��~JL�dDهf��Y{W�	���� 9��D$2#� �d�/jsqd��.P� �o;Z|�Ş�M���\C[�=���s;�ΰ��n��[�ÀÃ
pĞ
:sn��N+ݧ@D`v7�{8K�*�a,F�V��di{����2�$i�����Ef��)"��Y=���;�:��_k�$$�D_DO�&e���|�^k��{3�������` &a�(��M��4 h_7@$^����:�t�)��z�m�a׹�a=�n���.�+4���d��깋��m�m�7'bU����4N,�M�t/��7N+�z����TDA��7�V��E�"�#>J�^q�/�ϓ`uy�r��@�]Jh ��x߀@|Vt�~���m3O� ��O�_��H�SU؇0�r�!��G2��H ��UQ��<FLdR�G�
�޺��o�}D���<�4������ҹ Y�FX4�"d͉������{k�ŷ]�F�d�3�魝g"܋��	�M�&c���SQ d�� ����AQ/:2Z����N}��>��~�^���jQ.�r�({���$��)�����ɬ@ e���D�*t�@:'q�����rK� ���pZ`��Ц�A��9}�Wh +=���~w�3ί�>[w��xF����N���m��M�PeRMm����g���� Xm�I%�ٷv 	l_l03�o��L��8`��S�y�h�yw�W�M��ٴ.���
GT���=���@^� ����V�^�eه�u��4�kx������K%K�6��*��&��Z/�zv��Z%%��bb/qO�Ꙉ��X0�n#� ��λV@���Ryq;T���u�B� �hB�lD?c�ĮS8:�cq�F�"b%��s�;��O�?��
G)���Y|��� ��� i}��	�J�޴NTq�F�Xݠ Ev�ݥa^�ydG�nK�����Jh��-���-�/]��y��qk��T@*�Mo5�SZ����n˸jS%��TR{z���ͥ4|
/57En^L�u�����- k��TF^č9q$����F��y�T��햙'�gl�@D���Ω �X��gn��ז���= ����i;��m �i�4����I"u+� �����d=����ۻ	R�o{�7��m9������B�� IO��IO���$�	!I�$�	'���$����$��$�	'��IO��$ I?��$ I?���$�	!I@�$��IO��$ I?���$��B��`IO��$ I?�B��$�	'��(+$�k3q砕�+0
 ��d��D��� �@
B�i� (�P� � �@   � R (( Q@(�P�� � �sփ�4$�@)"B��WZ��RRT�T���(H
�T�hԑT�P
�P���T��B�R��w�           }                                  !C��r�*�
N�rn0w�o< j���WM��u!С���� ��kѢ�h��ҕv`�g�� � >���� n� � ��6z�h�`y {���Q� �����{�����Wk�x��� �	D���  |         |��|�C�CW3@PɠS���P��}�T�j����>ǐI` @�w�� x�F���   /4����Py{��fz��\ϝy�p{���������� �Fܻ���oXW{��ͺ2y���j�K��*��*6π           =}
s�>Xͽ5zgM�u�U�s��_/m(�]o /a��r�W�*�*�3TJ�\��4�����R���T����}�|Q%R���:�)*\�T��l�P���p  ��y�)J�唹��٪)I� �JR�E�R�nR��<����Ҋ��T��唹`�	UU��� MQ{*��s�咥%+�)}��-�x��]L�uѓ�I��4�v�|  �        �_M����^��r{�i�m8 ꂻ��kh&��n��t�{���{z�� pt)����@w�:�����|   �^��]��y��3�p�S#=����n�͕́Wm���(K�� v��C�޴���j�j]�p����Jj��6HE   �        ��\N�^�;�R�l=V�gy�W� ҅Y��P.��08�����`�׀�'�ޫ�<ڪ�T��]�-d��  �����ۥj��� 9������5��=���u�ǈ�� pҋ3{�&�Vz�� ���6(> 5=2���  S�`�)P   �O�I��P  ت�f�	������*R�  $�HCR�4 ���w���#����*�3��<|#K�K#P��~n|����B��	�����$������$����$�P$�	#$�������_������0��fn���	���:]$�lm,�Α��*
�e4ۚw�9t/��z�m.�����<��x���v@G�e�1���]l�+��9f�Y�r���}��'�u�:���jV ���mYSF={y5�����_Xx�ba=ݏ��rY�u�u<m�{�d��Wv[Әpg��9�8n��4�84�On�d��ggN�S�q3"�	���9�{,�f;����
�s!�Fkǫ5�Y6ޘ^N9�~0ڣ��cEO�p���,QPX��M��R�ĕ��U9 \oA�>ڻVlnf��ʙEӑ��aý��9�f.p�<����Cϫ�9����"	�f�5뼻u?���T/���b�3��8͹�5�f�i=���F*/,J�]�ڟe�(\0�g(�Wd���1U��3��7����������7�\��ǁ�#"�[g�b�V�qT�j�������K����s�E���߻��p��6�q��������Vk;3F�h��q여eu�5 ��q��NGJ!-�;�H0j�3~�CX��-��r@�OG[D��GW4����_�cjûKZ0|k�H�M<�T���a�\v>���u��N�˲ٳT��j�u��dt#�ϑV$pʳ^�L����!gvX�f��NH�eɫn�?%K�dќ���4H��+�ٚub
���.�#��{�����21욺=���Wo��rHػ���Y�����8�t`�W�5ӣ �ߤ�圥�ô�ͱ�/JɗLd�ޔ��^����lu����wa������S��,٤b{u���v��X�^��+�lP�U�3�T46_)�_]k�}ں��n:o.�o�N�a��{6SڍNJ �}ѵc�R,�޹5q�x7��p/N�0�^�7�oC�u�@��0nu��퐰ER�ޣoE�s#m�[̋;�� ��j����.n�]ÕL7Ȳ �O(:��tyc��E��	ph�W���OA+F��Ƨ+��mf��v���	;����νB�	Q�վ�о�ud�ǳ5m���r��5����a�̗6o>��l������5�z]�8��oIr&��Zۺ4�H�:&5����f�Y���N��f�Z��$[E����=�;dFC�$�i��Jٓ�'���VBYj���-�����5���fW֝L]	�2i�&��&3!ub��p�r#43��{&� ���,�ǵ��f6�&�C1��ml��0D��ʚ���dW� o>�;��4�x~W{S�\��6B�f�3��ݦ�U�P<E�È��լ&��BX���h+D�`h����/mp��sou�Wgj��8��U��a�%�H>�hD#��@�k��0&����B��\�ov0����廫,����[�CSg{�R=��o!G�8�	�>)�Y�{���Z�u��5M;�ȴ�Wh�Y�]��8�y=��d;Ű7�+�KU��Omν,ծ}�k;�yq ŴLx�.n��E=����t��% �QP|�R������Ew3�]�g�_���_��	8�)�k�7|giŢD�>�n�v��d�>Yz��tRr�Ҍfe��� a���[�$0��ʴ^��j�ʈ)��_����x=�����\�`$���vP�g�X�H�+z.%�5�� ��$�aK"ՉM��F��.�w�8(���`�O|�9�q+�\p���c����ȋ���K�1�j������
5Śz�Z�{]�[ױ�Yh��8���V.ܯ��L��[�]v�?����k���oi틠X����U��4F,f���|.Q�iK��uGa6��˗��w8�?��&ꯌ;��PE{��^�l�G�%�V�5%§:��|Bѧ��*�ΟE�I��8�Ni��uh/(`ݵM����u���U��כľ��2��%���nrwZ�.4���x�	:l8ƺ��hܙ,�S�`�I��;{&�Df,�K�����۠��RK��%n~A��H�<TrPb.�8JL����:1�Ёw��(���95��{	T北4֬C�sK��M{�:,�x�nv�5n��3����U�� d<�NgIl=���n����'�Sn�n��K���-��{���ڂ�x,�E��m[6�n�����M^�e���ǥ����b����IP��ڵ�ɬ�c8�q�ۼ)�!���$���K��������L֙���6��2�2�A�C@�1��5��Fc�?#�
�մb�ܗ�:��ةG���cwL�OD�,O��� u��VGE�w��7���n43{$��u�jIwm}��x���By>))c^�g�����8h��}�ѷ��+��_w\����VM�B���PO�[u�T��ymc��z�GU�v�v��Eߢ�x�X0�E@+��)�A(uV�v5m���$�����K�y2(��Ӝ 쪍�����ovM���w~gGQ���r,w8Loh�qK� �S��i�*�8z05l����C�46"j�*
���������$�F�a�Պ��Nr�ռ��֮RC�C�Ƞ�{rS���wp,ɻ�_Uu���4V��H8��;�/`��0�Ͷ�� �릇�D}��Ҳ�d���y��K�!%��79�v�3k�Őc@qީ��}{7�����*�k9�r��
����[6E�K���S��V�{O3�bi�C6Ǒju�钼	����t��lihc���X�P�co6Ő���5H��/ru�)����E���E��,e�&Cz9c���p�-Æ�͒���߷���ż���v\Ġ���_��]tS����K�Y	k|�7w��Β	��eq�̘n����`�+E�Pi#V����ݚ�Ν�f׮RwN�x��o>�~y&pk�8y�d�'x�q�U��gsm�{��=�ѯ{�Ӛ1�)�d��#vo�$��<�C$X�`3��;��-!�eGO��H4���Ӿ+�n�!�$�o'#��M�9�y�^��4����V�ہ[/��In0+m
K4$�Ĩ����N�c�&���u_%G�C0,�8$ݘ,8r����<	Ty�p�A�=�;��u��s�֋{�u�������\4� Iĵ]�e��wnͧZޢ<��_h+tG^t�^�q�t	˴����r����:��'!����.bX���ۮ 1;WWa�y��S�m3ߐ�̯�����_%I60��7W �����FŹ%�n�;�W�eO]�-�en�P�T�T;p���}e��v�:���+�r�е2��}U�����]�� ����	Y�1	Xt�t��-9�5|D��1�����~�U�)6-�R���NAF2���(3yV�����{u�(�#�1 KD�֍Wh��&����[R`C=��z�Ǝ�-��U]�����L:BX0=Govv0���=�˷�����#+��-����l�K��5̩ c��Ǻ���!by"����<�c{�`��1wݷ@ ^�ĸU���-pd����(=4��=;�l������0P��.�e�"���d#Xڰ�ĵ�a[Ёr�*�����o��Kk:���0�`�y��0w�!ٹw���[N[F�v]-�ef�ADw{�-���[�� w��9��uǷr�7��l���f�����=�;�ZcW�~���>�`���|zD�x�^�6��"�S�]���,v��;H����ԁ���;O�(�����<�0ґ��W��+�QTޤۯ�.og>�0����=�SІ[�� @���hޥK\�px�F�d1���z7��?��:(��P�v=u�N�u��ۧD&��{�7���`�g��Y�D�C�Ӈ�y��7FZ3a����צY`����46$�m��]�5�9!Xӛ�TҔx��Qv�^�SrX������� ����&�ĔJqf�Qm8Q2�^�ksf����{P�"gs���Z|h��6���Dm�,��ˏ�l�3펾%�s���.y����ob��P��+�*��7v�Td,2�K�im�5��*���Psp)��a�t��b��<��I�Ӹv�������Wٚi��;�v�e�VU�یn1�푠��>���7�h�W�,U���W�^��q�"*
��nW�K��׆pX�C�%�����v薜9���t��5 5֤ �{��3w-$�.1������oXǞ��<�Bon����6N���.R����K�V���7���=�\VF�R������4!�T�k��oiV�E-�qe}ݽ&��fN�K����r��7x��s�ɽ�����cZul���=3^�n����\VB�BV/��0G�}�^!�۽`�I掼�#���e�F���o�B������)t�$Aw\|�j_u�)nv��8��U��u)�t��s����tÆ����:�b=P��qB֜�GOgi�z���i^]���lؔ ��~���i�H�����;3��w63�����V�����*z��I�z<��Г�h��~�hHcb#�H:wUk-��f��\@��w��=t4�9�K�٫&v ���y���,S{Ỵ�U�{~u	�S�& f"�A�E�8lõ��g��<k-ME��6�]��Uc᝽���e)����]�̶���:��y��%��ɭD\9yL��u�9L�k@�ut��r<���y5����)N�W���4h�S>%�6s��P���)�t��ͮ��lB�i���A�'l�!JH �[�K��>�f�ƟeoV���s��t�j�w[�oD/	�f%28���F5�(��Nz�ϲ��A����A�����EȝTȞ�'7n'�z}��s"�f�,�P�2�[�_�����b*����n��3f�L���iq�
�Cg9���8.��dlCRd熼@x�k��\)�}�d�wk(���i`�!��7NZa	�p�;�$+�ї-ʘ�o��V������θ��/t�K��X07�C�1A��Ӭ�J���W�و����2إ�*��xz�s���݁��V��Y`f�ːq[V��-�~ڇ��;.P�X�$}+.Rmo����ڭ��q���/��̝#=̄1勚@�2xFo�t]c�u�N��ɸ����a�w�A�N�>��[혠Ib��-᫊	uܚݚE+ ����+<A�c\����Z�K��C��F���c�+�K��x���뚻�$�H;a�-�x��=������<��ձ|���si��]��{�w!��9)d��m6���3���x�P�S������H�n�$ݼfM���9�3����wW�'��6w���f�ׄ�-��&�	?	�m�阹��S�B�Vr���^�t �p�&qw��pi MT���6s�/���vB�]{�]�sY�d��j^Q-Y�+3:}�,���cݫu���&�MӚ��}%ءB	�#�;�D!v�:1e8��C%!;{T��Է�ޠ�V\�ڢ`�;�5�&�:���\�fm_&t1X�x��.Ŋ��Z�܌]�nL�{�I�f�2��1.K��s��q�e��/n�8K�k���X�Wwr���q��4l:(Sb��˃dGq)U&ȧu#0q��:Ae�����ot�V���WP<5�����[)QN�3�G���;gt�&���ȲTr��i&/N[�][:5s�F�Fu�T�ځ
�>��k�v�v��_F۾(%}F��o2�>g '�E�;7���{,����^���eǋ��p��x��wv�s�v�<v17�:k�	�VF���׺1z�C�dW�4A���M��{�LxU*�y7YtO�6��^�L�(�+t�r^��/A U��o]�Uyv&P��<M�l����[�����;Z�c��� �,$�FuW4}(wU2-v�nθn���\3 ��#��u׶��iu�I���e���<�<������C���7 4� Xv��`�Wk�[���Ƣ	ױ��O�3�D5�ͩ��JFͽlـn	KQ݈2�-�B]ʑ� �8wW`�u�x2�c���{��X�$R����p&մNP���n�5G3j��ٰk4n�f�C^�w���!��P"P߹�]`��T��j��`���@����*hY�S'�z��"��0�<b����JEf�f��eP"3
��RZ|�+�z`�Dp���,��3�X�I�=PhaX��\d�������c�kVL`ۚM
O�g ǃ�N�a�P��I��ί��v)#���@��.�wU�Z�x��ΠJ���H}k�ھ�1rf��۹�hDn�n�LDaO����a�.k׶.4�r���k&�Ѯ4�{/�K�/�.�ULu�d{'�n�,���1����#`�e.=�&U�;�u��+�y���"~a�2�u�v�QÊ�Vi(Ѻ�ν�X%9׭��w{D������Ĭ���9O>�G	�V��qGA��*ブ��H7{���u�f�硎h3�N��68�����z�*��J����h�{�����18Q�|;���� �B����P$XB� * H�E  @� E!$�H 
�,$��E� ,%d*H(I+$$ J�B, XE� � ! � �BHY �I	H�"��!(� RB(�P���"� ��,����BIXH�HT��RH�V 
��@��`I�Y����
B@���I
�RII 
BH� ��,�����H�H�! (Ad P!�� $�	%d�@P ����
� �Aa$� ,YH�$*I"�"� �BAd+$�HBE,(H
HIm �,� � �$���B! ��{��{�5�����E���̱�n+6b�$�C�+�2���r�ܮ�Ñ�z�>U{/`Aבe�`�O�pR�#st���v�yy�'�gq�-�59����ڒ���#b�h�=��G�؇I4�w�f�U�x��_������+�І5I�n���&|��e��=7��\�5��L�7�����ǀ����&F�����l����NUc��%��z����=C<=�y NPNYY̺�B�\�`�^'�rW5��cs�d�-dF�7ӽ/�a��b�nv�`��f�<1ǎ`E�-t��ބ{�h��jК�B���A2�S�Qgs��7Nn���;�c���1�����oB	76:U-ы}�^��H%�-@wҔNzo{�ė�}�>9Ũ�zc��z'y+��o9r�G��V��7|��ݯ��g��g�g�i��O�3� 8�6��������+�V�GU�>R0WJO�X˦��Lk�ږj��T�C������O�P���\N{���^��� �U��^'�/�т��K����}H�N;�6�{;W����	橲<��3΂iY"�Mۼ��V��w�&U��i'o#�7;�n��N���(tǮ��Rj�].��f7�Ǔ�ZzvEוelp��.v�0�688��q^P���/-�?aB;<�a{�uZ�{+��l5yg�f�((�?4���N����KQ9��Wm�������?-�a�.�&���,��]��O�)/��8:�vm]��}�R�s�h7%Z75������9�H!G-�gM�.�3#٨?\揚�#S����O_(};�O��x�3��>�k�":����ZK��R]��dbl\`xz����d�v?����X<"���9��{�c'���'5��z�A�dԞ������)	)��_#�lݽ�:�O�z��w%�X�]z0v���tY���Q���|��;2{�}=@C�'�w7[�qP��x�}��Rc�7���↥݉5�I����W=�Ax�n�;^>\}�kx! ��2��c������o������T=�+2{w~>���;�-E*9g��\���0��}��x�����Q�y��w��h�ӬƟ�r8�D�9=�_��<Ǖ֯mGs�H��l��.�4s��F-cu�������i�͗C��yה:(�,Eź
��h�=��e�����9����A�����۱L�����>�}[>V%�~$F��/��w/�L[=k�<����Z�{�Z�s�{p\��u){�������n��2ǰד��\��	�'�w'⮒V�9?ko�"���}�x=�)�c�,������^�{����g��qr�r�m�s3�����5��<pI�6�^M�M=�7 }9.l��?/Og�2��"�ۼ�΃�ʎo��B�������M'R��G�>�^n�>�
���C^�"�^�۾������PrL�1C䧫����&��{��C��J�|����37���tv7�7�x�_.�dy 
]��/��/�T�1������_I��t{C����JM�-�/G�.hU�3~�F�t�qN�8.�r��;��F�����L��GU�L��}Q�����ٹ��Ⴃ�s�5��H7��pzM���>�^�n{�m]�Q���{�ԏ�9V��׀�`����#�ز#'{^�ê^������g'�I0�����I��<��;B����ԧ㏂�5͝Gdع�Ӎ���g\�h��|��͞�ޒ(>�4kMtӶ��X>��K��@{ޢ)�������`}f�I��Y~������E�����{4��;uWP�rg-�@����}�=xc#�/��+�]=y�r�e����Bl/�^��V1�u�0�^U�j�� =�2������fѶ��*F$o��#+c���l��ˈ�t��j�~=��}���!��KE2���}���a[�}���y�Ǟ��R�K�R�3����B��19�d��W'���K#�P܉�y�]�!��v��F^����W�hx�nu*��c/����/��/u�^og�wwT���w��Յy��s� v?i{�J�f�����w{�Ԟd��O�[H����U�'����E���� *��{�a����s�r�S�{�[icF�U�G����o�*1��{A�=F
񉁳�u�_B��,�w�g1��=4�ݓ�{�Z�=��N\�e�-�L���@�Z;p^{spy��3ܤ�u�ލՒ/NW�
��ob[��q��Q�#��a@�`~��vԮ��>�罱�~ފ/\<}�D�i�r>�w��~E`�ȱ���>�piӆ�ݽ=�y���sBEbD�'7�6�@�Ƽ#�x3�0n٫j�D�1��r?(�J[܆f�����?�܊A�!��?>�L���n;����w
q�;1 �2��VL����e3øa��O�ݤ!�U�دN>������WQ���5� 2�wמJ�y_+��};�;Y�~�ъ������{�s5zۧu�����F��{�^�U�^��]~Er"�r9ۄ���9�k�f��<y9���T+�;7��1�N��N{b����]���u��Z����}}F�ܗ��=�E|�uwI*��G��f�#��kÂ[��D�;���|C�*�Gh[�<f��A;0v_{�ԇ@4Ww�ޜ��.��<��d�.l]5���N����<��gS�qp2���_QɅ}2I�]��.ᛲ��}��6ݠNMg�;��D2��ӑ]����եr���fԎD�@�����P�Oo��i��.{�)�1��#��I�kzpK�im�:����#۽�g��_u�y�Pũ��1��O,�׃�={5d�4�״�'��+�=���!���f��(�gA�6xM�{�zlFc�Q�͌�1�{�Jf5�C�k�8����훯2�7{ͷ��y�9�<�ѝ2�C�l�]��=�S�\��|��9:���fR���?r��_QY�un{�K�l�;�n\�r�8����=q_A�i}��<9��wyᚽ$C�����J�������*����k�f�Ou�y���B����kp�iq��:���y�]���,�F��bs�����P9��8�������>����`ѣ�\R.ꣻ{;�d���������vz�,�?�K;���ǧ�M���Ű7�!�Q������y����z��>���Ș��<��??{�zzg��
k�ەf<eI����8,c��?qc^v�xaO�z{i��3�a�%Y��p�,Qe)9�9=�u���"n�O��]�8��;�Tg:�^~#�V���y�HZ+'�$*���=�V�1��gz���D���:����-�y�rb~ @:��H"9�Y�u�����C�l�U�UF���yvy-�</�;�K�N)ɦ�L1�G��o�`��B�d��!臚�o}��7�:��ܽ�ƽ�Q�-��;9.��}�-�x/w�.�ݞbV�V���Y�¤p��p��ۚڙ��2�տ:�;�y�'p���k����»f�|My{�ۣ���@B�!{a�3%P�vh���s_l�UsnI�a��N�:�V�E]�5��Sl{�����rmɗ��Hܕv��]�n�Ƚ��"Z]�o��$h�Luu��u���k��,k�����;�wj�y�g37�k�����Y�{�J|�9���i��;T�X��;��wo�R�3ܲ,���^��M�ك۷�ܼ(��.�4y:8La��u<4��f=�|Z�u<�Oi�$$��oaܳ2��&O�XU�g/s�ov�,E���WzU�>�"X�n�E��83w�!OrK8����D�z��,���;z�Xʎz��T��^"/3yy&��`�g�U����D��=�i��c�1��{n����ah{=�;}�\��0���C���{z�f�$w�S��Z�=�ˢ�Ҏ��XfM|1��3�^c��7�)96�G�jΕ�e�����g~�@���ka/{���WҜˑ��KJ�<�rr�f���5L���&�I�0�o��Л�B����=��Fcwr����m4`����f��^�+r���2
����^�K���Ͻ���Q��N<G��](bn���s�.��=�f���h�p��_h�Wn�'�6��&��c]ɟv����)�������5�\�ϯ����sF˒� =y6�w��,��[�l���I��#����Q�Y��qR﷜�:������/,|�&k���z@z��t幥v�V,�qa0{������.Xsf#'nox B�b�&����w�}]�w�f�"g{X1�F�=�;�|�0�x5yI�3ާ����>QU���0W�_�0sZ|[��|u���A��*�^s9�/��ؤ!W���v�]��{�2^���.��$��k��rQ�����zZ��s��������=j��"��sD(�/I�{|��|Y��87yN��mݩ�Y5.���L/�2q.u�;7��_�m��Fn�ߺ
���p����Wu���]�k���:=�ܹW�}}�2��3����O�j_\>O��Av}p|�	_,�t��~�SЄѱ�? h�7xb�J����w<�ް{'Nv�F�Ųr��{�W���b����yu8^��Wq�"j��}�'����� � �v����/����|wKn�������ƥd��g'���Zw�x6;FKқ˽n������Ћփ�}zA婪���>OZ�����}3(Db�~I�u��Ǉ�{��ع�Nݬ�{8Qp6pܵ��_q����қ7:l`k��h��CL��>Hd�)��Y8���a�-S�'����v�R1��/����h��~|���F7:��QNT.O>=ϲ��L�f�-}���o�El�[��0sb���]�	���W߸Y�i:�V�C�e[巄�Gϫ�V?������RyJ^�����@z�帴)94��<|�qހw �v�x�p��+~�o��@��U���͑���Fg'�>�#��^�������{I<D�$�H�O��=�v�pqۅ$����T�h�VZ�v\'ݻ��à^�i1��]<����Ōx=�u��Щ�*��մ��We��A��gk�q�5���=����y�h�!�u��'���G�31g{|�rEמ<Ϟ�q�3�o�8�F_\�i���y��O%S��]���9�l0�m:pe|1�G�ߣ�݃�R�^�ޝ��������,��o�7��zb�-�Ě��J��qHt�.��*�n�2�8�,��S��6�cMk}8�� �MS�u_?X����w�R<)y6Š`����vm���}������޶���d�˸��P�o��>;������Ƶ��.��/=w4��^G������rs���=�7yov�=��ȔXb�m�ޮ�_���zC�N/�]��
�e�xu%�#���B��e���率�QG={�{�{/��'��k�<ރAM h����gop���ό�f�L����q�#<�\s��i�ƍ�|Ꮦ��J{ �G�FT��7��^�^�ӣf�0#�ጼLCg�_d���>~b���Ϥ�a����ck<��.x�]L�MP��������"#|u�=�s���u��S!��%���W]�w�޵qž���K	��Y���x��r�Fd�o�w="��k�r\��jwcdxx��`��z��MB���w�uv�<ߏ`i��r
�yS�L�z�V��ʎv��Wq��[!y��7�'���^4<����k�//�X�*��뇺���K�Tf���O�ʜ[��!��o��o'�|�)Fz9�J��x=�7t'�;�v>���o
G�z}Rڰrb��<8[��%�O;{��g��vg{�����)p�ǵ o\������|�l8���`��d��>sO����e-x0.Y����j���ٙc^K&!��}mjd@ӳ:k�	��6��O��i~�;;\�ɾ����w��Gx޲kkx_1�����ݎHL
A���c����Ia���|qԃ>����� �[�)���˹�����!�2|O�#�#F�U�N���0z�Q�at��T��p�{�lpm+��mG=ay�c�ź3�ޛx�qj
Fv�����E��xmѽ̓����9e��y�{rӓ�Ii/;U��(��l�܏��n�r�nP��V�!�G������ݕu��A��$�!�?TC�գ��=_������{��P�{ص��r���K(d94�gg3�o��i�~|D�f��&�{�鉏d�ى\WUO���݇��{\
��s�A8���9����C�y2�h�V+�J&�XO6'	�w�D�z�c8�>�,���x7p��'-{z79�:w(ܷ��"��I/�D�p��!���)]����(-�nx�7���%��:>����yH����S�./>�!��Ր~K'�g�`}��֤'yG�[D����4C�N{���H�!�W�Ν*����uVz종qk��:��b��@��y{/����Wܫ;�B�;Z}�mc#t���e�K5�{�Ηtc��y����tS���$�3r?]"�/!@׏{��ٱ�ݞI���&����]�2���D����<���u�	��0��o�e���\pØ�Y����{9�{ى&�t�IK���T(&�M �Ř��G���@���x-�W���w���Uӣ����^ǔ?1���سkq�fq��c~�Os�.�%_��?���1�7b���p��F�l��4`
f��om��	��Ј3�d_8 �@�:�_K��2�d:�$3��D�cQ�@�<���>���{�^�9:�N0�=����|�����/.j�응�jVP���=�g{�����X��li%Ƹqɩt�IWN��e:��m����,v&�$ش��my���l��
�:86�6y���)&�C�ˁ�q�ۣ�v,b�L\�rc�r�Np\k��G�q��ix���kLrq��ୁ	�Bն'D5���]��n��-d���Cp�]�ܙ��-M�89+-r���^�q��,r�S���^^n�]I���k-0�w��HƱ1��WLtxm�َ5�kq�����TG�F:�p��x�uft�ڬ�į7��<e�{�U��n���7v�f���仐s	Mb��@q	s�w,9���]V�d��t��X��n	�Ҡz ޲qG��σ������/\;���Z�<v����dZ��� okaa�Y�xs7u��=O�ۜ]p��`^�5���Q��v9ۡ�]��v��c;��a���4���v8�t�8�mu��N�釄���j��j��A�\۹�y���e��A���ۋ�^2���kUz��y�7��dk9��,S��rt؋7ZK�v^o÷m�wt�^V�jŝ3��˲wG	���7;s�mm�=�s;uUt�m����ky�sL�e7m�
��m��#�):DP̈́p��:�G=d��oNy	d�0�FTv�����Y��{qv��Er3h��ק�̓۷kLLf�U��Hn�Kj)��O	�ڈ�"�	���ފ�k���vWm�8/;�Q���q��c�k�lj*b��n��q�OeP��`<�<��=s<�Cb��r]M��6����K����ͅ,9LF�� i/G;�^�Ӵ{g6�٬x�'3�/Qly�n�q�@hT�Sb�`�ez��7a:Gk�n��t]�v�z���n�x�3o<�sX���_ΫN���e�4[9!$���b�o��ζ�ݙ�Й�sJd��S[��vǮ2�b0��wi:�Yݸ��2N)0onմ�;)	��&F�ػuvޫ^(�j➻zx���6ݝ5���X���ս�+��Ƃ�ۈ-�ӹ��[qq��y}n��lqq���nN�꛶9}���>�������l�.y�]�v�xl����69�8�\�q�{6d�ٯ=�b��v��ܪ��]�"6�U7L�{k����3vPh��6^�3�F9�cY�R�'v��(����hm����!l���l<`0[cAg�0��G=��u�V��-��Y}nE��v-ܣP�=�:���6�&�ʕ`��<�v�@|���q�������[��y�Z�՝-�T��[�	�/i6+���l�wk�â��Mr�@p��:Qݵ��r{m�%��%��p�m�t�<Hau�j�\��6�;N���k�h��(A�g۱۶G
���r�<Ŷb/"��k�;=��-�Ip�m�3mے��<\�F��*���$@��cs ���s�t�)in�o-�Wu��X��Xy���}n<�3Ś��	��=�ur�k�����C�D=���� ����ݻ��[��¸���cO^m�9h
��+t�yOk�;r.��k;=�s��0�}2j�V�jC�<�a���	��s�J�x맜N��6�㵜=�:�^rq�/���⥢7�N �.n.��8:�X�iL���v㱂z���!�ό���"f��ʆ{hX��]��u;9m3�t�u\��!v�ۡ�/^I�rm���V4���f���c1�����F���^B�nݼf6��0�/m��e��z�y/Y{miSܝ.7zݹ#\p�<��V�]y3t�x����1�gnunh����u��xF�[�lw+Ϟ������RT����u�nbݰ-��]��;k[��� �D�8y�a���n��r`x�v�.�k��n�n��'�C/�c�h�<8���t�x����ը�h1��]�v]�ݮ�y��ܖ�.u�Ϯ��˝�c�[�`N,N�Y�=�ˍ��t�5m׻@�]C����vƱX����qnu��^!���Kv��7e}\(C�W\��m��s͸L���C�����'6���;tJzwn���ַ&����s�����kΒڨJL��Y��@����Y�V;���@6���uƽ��z�Ӱ�9�J�d�%nYσ��/<�ݱ�ۂ���.�e��g��ڻF���#g���َ&�c�7؞x�/�GEvy�7����q���uݼ�m�.v�N��\��ݎ���)�Y'��\[�6;Q��g�E{��qՕ�G��1�E���S�[u�,�{C�֫���k�۠�+�/�kv���8ۍ�.�5�i]=����qX]w5�f��a����Da�qt].1\.���M������{,;��.F�=��m��;Q�����J��+����Ƽ@�^���oQm�=�9ANNñ�C��.E�@�=�h!ubŪ.��A��qX�RO=�Onv��n'u71���so3��d�<3�M��=��͎;t4n3�01�ûsv�����wo:���ݍ+��N���櫭v�:M�n	��
�^��^��7!�u�)�y�Z8v�:��t.vM�u���{l��^��X5<�c�[h������u���§v�r�O{�N�x2v��y�%��Q���ez۫���`8��J��5���Ggd�omRd�x�N��ݶ}���������n��n���ڮ�6,�s�<N}v�w>�$`G4@�m\��le��C����:�zN�>ź������A�+��G&��=K��-��1�C4��2�B�����͞|���m���Ĝ�Ǩ8�{^�F�;6}�C�.�p�����t�
��l��:�w%�k7���բz����]�Y�ӂ�ۧjѹ�м㱡� N�z���{(�OGZ��v�諢^5�qрF8�bw�Ѽ�z���u�,�|
N8��s��-����K�=�+��]k���y�y\�څ��k��gn�#�Z6���H� k1&���ٵ�n{v�$�j�V����{c�ݸ7�{/2�Ŷ,=qWy�/j�t��oY��Ǝ�S\!ں�7n�%S�e�\N��c�mu���n��v��Y�=���tcJ>�[\:N�K������S�sH�8#��c��l�.Nnw5���bt7���σ<@��䱣Zx��^{J�l�>�U)ne��V��v	�&���Ɍ��rp>�k��O90D$�5��]\]����!����I�vu�[��v������t���
l��v�wb�"؎��:w��:�ۮ��q\p	.bⵌ���;w����sۄ�p����<�rs/)�����֖�C9[Lzoܰ�c�foO/A����b�:Ԉ��,�����]�ݗ�=���� �&ݭ�vsa��J�n8ݸ�S1k�V	�ԏ.oU�֍�<�0���P���殽�v�˻r�x�;��F蝼]l�\�.�q�gz���lCĮP8ζ�\b�2�l��Zy�<��G�6^7;�B��v�s�v�cԹ f7���鞃��ޓ&��y�������=cp�k�nz9�]���hCvz�vH�:�$(��է�c'nՖkBç]Nvv��OKs�����i��r�n��{v���	ü�����c<뤐M.�nܱqr<��v'=t�@�����y�l�f��u5�g>*��i=�s�v�O8�kƙ�!���� ;�`��q��<vی�p{�/t1��N�e��\�6��x8J�9v��OM7V��ݑ7fz�p LٹyJ�ಌG��\�vۃS��g�S<uĸ9D�qsض�g�{Z덻s�-n�]uz�n�8s����^wt/�u.���:�&����/19�vZm�yMp�u�E�N��<�cs��s��7]�9��G���p�4y7c^��׮����n�O���z�t�Dr�9�Mt]s�^^�	g��[l6��ݺ.�����k����n��u��9��Si�c^�ܵ�ь$�Ŭ���l�"���۶Z�\���]�'��u�v�cG�z�u!v�4�'H]��F��EX�WA%�a�J��5�m;�C՞�N�U���z�����RN�M�sv����ܗ8��z�[�M:^��e�����7o)�N��tݲ.l��&�x8��ln�ݎ��;�$�vG�NL��v8{��e ����ې�1�%�$��gv���k�+[�ƭ�=�y��L	�`���s�*3 t6��n2�h��������Oc��mێ����c��i�e�VN,h�f����\�Q�8�i-�ι��n�a[�ۋ������s/��g
���m�g'n��ڸ���Ff�`�����<�sDC�(�^u����IԞ]�v�n�����qn�n�K�������xp`��hzܻ\l�3���r���+����Bؓ'g��[Bq������n�᫅�+�z��Q�D�klvqƹMd3cj.�cw;����Z��ڷ�G���pp���SV�gHX|ns<S����ø�^�[�{A�Z��ū���%z-���[�޷!vb5���������@Y�]//m�lX�����5^��؁w��)���݆t��f�ɍs��t�U��S��qϵv�N�NHOc[d�//&�.���i��K������#��Vܹ�N+�=��z�Y16W�o9v�uP�y�C<��kl�v�01�M%Z'���M���r�7\N��ˣ�1�m��G�⪥�����+���W.����ѻA�˝Ϟս�����Q��h9��L�ˮ�j�L�N��x�&y��A�t��{�2��ƶ�aM��q�m�:�5nu�pJ]��k��:��6!.��׍�Sn�6%��
ɳv�x5m���n�I�U�ᬫs̴Ug������N���3���l��C=�n����0[:/�"��n�\Z���]�Dn�q�1I�zwgI<݋�����Zns�.�����+Y+*��V+cJ�ed㟴��+��Z2����Ekj�Pk+-�Iyv,*aS��m*�ŅJ5�c�h�[Q]��ъ��T(�R�,�
�kX�QQ��������DSk[m�K�*��jԭ��V,�l�cK
�1b����%-�-(���Z��R�k*d�sjQ��
�v�Ъ�sX�J"-��mD��n��W�,S��Ķ�"!VҲ*�R.r.�UZ�Ԓ����-��mZ��jE-)`ԅmv5�Υ3llJ��E\�,Z�V"YiZ�iQc�ҭ9J��AUJ�婊�q�s`�Z�ʙ)�Z���Fҵ2S-YR��Rղ�ԅRq2GPTchV�J�֤mJ��ڢ��Kk2�ʵ1k�U��-��uYW5T��b,�-�b��I�s�����1y�mԒ�j��������u�F���t��YhNv�V
�l\V�5�v�cdCs��n��n�-����&�݇��gu�u��u���Ż��)��|Q�cw%��.��-�a�nSuݘ�j1��׫�\�ܛZ�ӛW��)p!�n�V�ƚ��]�aq烁�d���04�8��AZ7��1��x��W�� O�b���Z�3�xN��C�ۇ�(q�[n��뮢������F�e���׍��J�3�s�;e#����������C� �<��ܛ�v�b��K��vz�@���A�wm��<'��ɓ��Wl��������v�� m��zKjv��=U܇b��dJ'�]�{Pn����t\p�g��n�{wǍ�\۟���n8�K�� hM�t��VA'O:�wb=]��nӀ�<���5����F(��F�{��==�G�l=me��\�^�'�pӢ�W	�^�䷮N��u�KñOb��탟%��'��s�s½p�f�1�1���9{> μ����׭��7'��kqb릸�w'�k��nEY;m�[Ec����7W&�ݷE�Dp�uǇ�<m���u��]���,C��F�n������+[�=Wΰ8�Nf�����Ѯ��M���~��F�ݵ��q�o;^ڡ�t��ipgl��i�[v�՞��pu�s��]���j�=�9����u��y���cۄ�{A�m��Y�&�i�n�kM��@=b�S���:x����}��8�=���n�MF�
q0�.��f��t�[�o�] �6�c�N;v��f""v�s����$�9�g�i��۱�s��z�l n֭���v�ꋲg Eq� �5˝;=(vđ����N�F�Qe㚸.�zN!ݬ����'<�/;p�u����؝��V���K�i�؏����7M���o�;l鈺��/\��k����s�J��5��xI$ḙy�V�vJ�9�mV����tmT[2�����n�kZܥ��1s��^<�<��������ci�s��N^Cc/l���ݸ7l<����۟�61�xU��C(x��v|`���Ll�[T�"�\R��<� �8�98��� v����^2�9�<;������.�ɜ=�3�.��q��ȝ�����߿}��#9��H���zT�y�� =5{P�[kN�l��ɚ��I<���B�f6�D0R�I`�~T���l�w��a'����A>=q=!x���X�=U��V�6��H���
^}��$���#S��b�*U[�><����|v�t�٣��	�	h��=��g+T2*W�	ee9'ē{/�	�v^�Q��<B��@9�t����dE.%$t�تDk���J}6��I�xĂA�� O}����zW��Т�)_��F���:��9���.��/nsZ{N�k���W���������Rw�I��A'6��H'û/h#jU�=kR	� ��فK���E��NK�T@>ު5S�����e\�V�^ݦ'���9�#8Cʜh\��+�]m�����i�;fi�yS�g2�9"��c;�o�Z�3t���J�>$�콪$۫�������J�Ǒ�"E3��*g\�	�ohQ�b¼�1b�KB�'�y�콚 ��/-�N)%@d������j�s�3�.I$Y��+��-����6��¾����`K<�f&	��.������R	;&�rb�N�{z��	iI
w��:��:�
&!p�v��{[+s�n��[t�8Z�8v�z�;v�\>�L����S.18�����H$�Q$�t,�&�ɼ��L�@�r�w��F������t7�|H,j���a��{���z߽<��z�L��r{��l�W�A8���ʈ0���:���g])� �v�f�����j�����Q�+%غIVVʺ5W]��,���zT�_n�Ժ�}�_V,�������O+��i%��pG8Ǜᢡy�.fOx�@����R��t�x�!"0ۊ�T��z���Y:�>9UWB�:q�G_+�RE#���:fz�싎�S-L0[bB��S�=��b:T��e�����#�ꪼA�F�R	$�W"����8F������' 6�r�0���n�s����)l�$�27>bS��^h
���DgBJ/�k;��UU���|O�yٟ*�ɼ�5{��}T	��NI3�kQE#(8����_f���������EH�t�A��s �9���z�M��S���9�l��b%?�L��l��v�\��yڕ}���Y��(�{9$��W0|i����D�rz^�FŘ%o^`�Hdܹ'��v�ِI#�3k;L�r{�'k��m`4Di�l��fe#3�x���)���s_��灖�Wnj6`�	w�Ì#�w���k%��߱�̋��,�$P����"�Ь������U/U$�ͪw�����s�4	�{���I��f~>5���Լ��;��m��v�i�M���<�a�z��gCō�9��le݊7@��?>�X�҅C���$���Vd�	�3j�ojLU���'7�k�\��A��r6hDNBJD�j��UTA��˙�N��@+1��s��$����^�Ř�y�i�ft�L4�`'�R{�l��^�W��2����%�R�?֢� K���p`ٚ���ZF%T)D�_	\qX����6�t�>'Ƴ3�P$�M��;TC�� ����|a���N|_=�A ��LB���l��r}]��4��N|R9�ݱ@���u쥅�0�����Us�84oy,��l��[�sA��'�ή���:j�!�������yI���-(�R�.6�r6C�ca@�E����.Ŏݎ�)�3��G2���%Y��ch�۔᲏.�k]�L�CQ�b��i� Y�8M�X��<�]���Z��m������]v�m[}t��;:��\N8�8ݏ�c�-ksk���xH+Z@���`Wͼ��W�;��t�`;bݷ���Ls���9K��OaFT�I����N@m�9���t�$m�n�g�v^'��2�����y=	��Ѕ�������ߦQD�J�/UH�F�f�H=���{�v8��ݺt��ֲ`�ٳ@�����*ciI/�����j�F��Y	}�B�I�v�S��SR��/�j>���iF�����뙃#�vđݶ�Oh����2L�@���H=�ܓ�8N�i��A8�ړ�+o�)���i���#5ېI&����Wm�*����W�����}ۅ�?Cu�!���W""6%fU��޺�1�[TH'#���W1(�nοavR@����rc��l���,���h��Ӷ����Ӥ9:}��b�u��q���D�|Z��H6uڟI Ws�>,��y��75�T	��v���g�.@��J�|�`���a˙q�f��O����)I�ֳڪo1��
��ޯ5|��$�ס�7��)S��6���v]93�7�vM��ͬ��;����c�>�&��s<��$�]� ��W"1�N����5��j'�r�� e(�-3&�I�%G])$������m^7.�j�iywĂ|�y�O�A������"�L�M�P=�U��Ffd�>��<��=)������V,9&�b��*�i��A8�ړ�+g�	���J��t�ݣ�F�Y�I>9��D�f�VϷ~��e�\t�2�*0Y(�"���9�;���Fp�@�WPD���zk?����~Ќ�?Cu�	�9|�Dx��ͪܑfzR�Mw+��F�p�A��nK]�^��jQ�V�l���I$��vd�f�Mvd�wq�Ky�]��x�7�H��iM|�`��ۙ��> {�d����up�D�GDL�s�O�Q�=���0f|�Nn,h<�t��{�ND6�Ed{�F0�8�ldRJW�^+� �H��ڢg��-2�q�ܐV�����SY����$���B$^�t�$F;P,]d��wQ�(�yvH71{(�TN*- a��%���5S@��]�5ے�+	��Yq ����(��v�����s����!�j��Wb1���ɖ������{s�8�`tGS˜�4�p�A8��P�GăY����юԃI�6�GB�<rb�P$��u
��Ҁ������H$���F��v��Wo� �H���>��h\M������m�۩�w,���T�	��}�U�:�	�
cC��zRmt'33��$�c�>'���qZPIi4���ꮓm����b�I��ڢA�׊A �tu��3QF�����v�F渺Wak����Dwo���a��n��ݼ�
����7sPee8s��A�U��v�9�$8�}�B�Q�-3&�I�$(ۥ$teϕڼ'��vɞyu^'��R	$�G\�'��b�;F�U��壪zƫ�{F��vG�t=��g��I\=oL#q�sOL2�.C>�'��
 �&:3e����^)�O���$�IdR!�=�ӄ�@���I�=K�(�%$w�ߕ��{`c0��̉����I�{�A$�k���>ͫ���yASOk��{\4C~��JZ��\uJ$��'N���Ԯ��utH$d<�$tuD��#|��b��n|a��T�E��	ٙ���3�A$�Erځ#Ċ�ͦw3�`�9\��ٳ�� ���iM.:�A��ٕ�b�c�"�+��� I���ü���u!�������pT
�Y)�OBRf�7��ZY_��}%����B,(�f�7T^A���R�9T�͹�l����'��X@��AI��I3�\�x�]RV-���;�^&��#γ��ɋ�$�t�v���Ng<�3L���]�ȧk���ӣ��>�EzK�΋�'�����9ᎍZ{�d�݌:�/�vo���.!�n37m��x��o[��\��u��7�u1{2���: �������tWlt�n�]�c�Z�f머�h{
�����`���<�^m֚۟�땍�[g��U���>;o�pY�x�::�sh�������a4a'|����GteD�	����qK�k��5e�����}��^��e�p�	�M��9�U^�^�G����EsZO��.��H5��4H$�';&�������"���RGO|��̂�Ϊ �T��:���������R>5��4O�=�4Y,~��Z��InFGC'�3g���ww6h�GB�J��]:��L�`�E�i���d�@l�
���O����&wD���#y-��	�of�x�yf93bɺ3@�X=�AR[yZM�d ㍃@�:.����̜v�|ݾw���r���FاM��ߟ��A�=���zQS Fvf�<����
�#��5í^5��T	�F��e��)HV�����t������n�֨dv��2&���$�^���{kOR��-��
��gy��EG�qڇ�y�l��F{���Ff�U���A&�wL�x��\'!>9S�Nh���t�UI�܂A��F��E��)2H=y�4A��R��*H�a8ԑ�w�v���>���N��U�YnI�k��u����V�'��P��(�D�P�~-���I ��\��6/*�w]T	����Aϗޡ�${��9�pT���L�,kc;��N�QUӣ��V�6=鍢�1�{@�k������&
��}��f�H�vĂA��f@<r�o�.{���'.���b}ӋZ�j&�"7�6|�X~g���3�3tA�� �I��dI[>�%�*w(�'�����,BE��u˰';Ϡ�Nxk9�2�nx���r�b��O{�٧�.��Ek�Ot�:�x|sz0�E}l}�f��>��{ݥn�v[�l�2-t���ݻ�9��?p(��	c�К�~���_hj<^����GS�As�ttC8�Is�"��58���rɨw�:F��m��⢄��ݜ7<kk��-�!_���>�l�V�N��Uh�9cetm�ű��<����w|�
Ȩ�/��ʙ���co}��=��J��%�\��R�W���{��d*'�yF�t��;�<ѣV.����"[��U&GJz-��n�?���U���������w�X+C[gxY2Ī���g�z���c��^�mǉPW��y!��}���h~}^)������{�"^����xm��9R�&q�,g4��D��0�=����c�ۈ�jQt͜w{�cf��-�J�:�^�oMB�;6Z��6�"Vr���H&��0�7�0{tP�+f.�������oI����X�u�aɛʺ�,�T�_.�r�U���x�;&��t.Yq��~,�x��ܢ��1��q[�	��������7��~�%=F�*��ޛ���o�� ��^Ω�Z����*Hs/,/�SfD�yak&��x�:�\��ɚF�!��,0::���/E�oa=���n����'g�xyg#����'+ޟz�j6O;1��Й��v�ݱ��=���I��e�B����i	������F�ܕ���<��A?W��.���ٜ0��J�|������u�)�m�������
E"Qլ�Ѳ�mm���j�4ͪʌID+T�+J��%�*�SR��j���B�VVd�8b���Līj���恒��[Vԯ�-�qb�ƕ;q�C8��W�n���3�*�aYm�Z�b�E�B�ڢVV1��eJ�nlL�cmb�.J���j�,����9���q�PP�H(�YD�-Uu�S �R��%QY��al�%m-k��*��"$�NR�,�Dc҅KeTjX�miU*5��ţҪ�[+�(+*Ȳ�R���)iJ+X�m����"9�� ԭh��s�mR��-��%8т(�,WjdL��[(�hQLͪ)Z{N��=�ؒMo+�{D� ����l�go��� Z����[�̒	�����{V:_*�N,��@�0ۆЅJ�l��A���@R��f�Z>�v�s9Y	�_fЫ��ĂsX����N=�.�x������뮸����L����b�H"�n��T8D�P�~-�O�I9z�DI��ڢ6M�_^غ�O�wc�I'����5��BI����Q��(�[6N�;�1��A5��ω'�}�TF=�(��WZS�>��b�jP���Q����Onf�
U1J{c	5ܮc��}�TH�����H�)O�ۦ*��#|��R ��5�0�|�3�4߆52�xO.��܌�:����OnvXD��!�ٓέ�ř��m��< ��|��t3�͟��){�����M��W��%gf�8K�3>{^���}M	�%Ss�[n#�5�!�P�P��+ �j���O��6��$�R��]SC�1�%'�B?��D'\#���eE^
��k��#[�n�cl�V������HC������A �Κ$c� ��.eނ����@�R��{{:h-N�N,�"�u^<�9'ǷyӲgEut��p�i�A9��U�I=�܂M]��.�2Ug�dS]�eN��䵻�D�z��$�gwY{2Et�����}ٳ@�H=�܂}ә[P҄Hm4��2�P�;w��wDV�UQ����'Ě�WSq�j���>%+ʚ&�ˍh�P�\1>+n���A��rT���&�z��,�d��mP�	u۟	5ܮb˃���؉�})�Ңoڻ��]�o�a��\�%'΄�{�՞���}���ȼ��fmAn��ý	"횜���r�F�<1_WD�D�&���\��v5��ip�@fh[�� viI�>we�mv�r��WkWl�8o<I���]Y&��-�7�]#��#����Ș�ytvz�n{n��i�0m{�����s�)�,Pό�n�Ɛ�^94���ݛ��O[�s��7f{q<ݸz�#Ƹv8�[=�yse����卌�|�w@VN����l��3s�F�hy�N�c�wN���Cub�i�G[��>.z�땹���H�) �i�(J)ML$�U���m�H�v�I��dp�P�r�ʾκ�ߦJH�=Le�QE#t�W� ��;Ur���&�nn��t�Ēky\��N+�����S���O�WE6�,�"�uG[�$�A��S����ގuUq�m��$�k)�$w*25�֠Bp_�l�>-v�!.$D�
��kx�$��td�O_f��jhQz�x��lO=:��(D��J���S�ۙ��9Qb
U��>.�\�e����ڣL����ۻ����r�0�Fǖ���9��x4G���͖���;�G]�lѹ�c������e����|	��kʈ��͚��;(\K(���� ��U1�X��L&Q�-M�5TY]y5w>�����E��./����_/y��to�g�ey�H$��|��weƏ����Bt��{��\��Ѷ�Ӂ.�_I�Um�l׈��&�Uk==����:�h�ڂˆ��f2��bff�|nYѽ�{v��I��S ��ٲ*��Sp�d��[���t���pV��}KdA�o76hG,��#zu�3�����Kf
���DB,?�nK]� \m12.w����9 �f|I5��B�<�ܚ�zrnN��=���Lpa��p����$1?9��b��e�R��cRk�N��ۏk������߯}�S�S*�X��w�6�(	<���ғ�w$ve)U���U"$_vuQ>�/[	�-����d��w�|������\w`�M�f�	<����ͽ��<����MwAU�)��eۂ�P:���D�G-�>$S���r����`�̺&G�C�DKݯv5ѓZ����S,r%��60��r�="ą����r�jr��%/2��j���<O��{T	$��rD�/C	&�,�m!��dB�L-q٬�%)��$�I�Ă:�VV�{�>�κ�F��T�b!��C�Ǆ�Yʦ*�nwtժ��$^m�
$��s�|O��*1W�S�*�X���@� #�p�:���94�@���5�vxv��r�n��B!��o;����)��ʆ��}�(�E��$�G_:2x��DYٱ=3`�@9�LONV[P�ͦ�QSʌ����8����yR����ɧ$�A��s ��W�tLAf�^�v���)��E�
ܧ${q\��x7���iSu^$�ɷ$�A��s�U�)�8D6�C����k�&�6�7đ�T�{yY�	o�'��U&�k��*k�S�������uƹ�F%����~��e'<pb��1g=�f��W>�>��T>���(��`��̅|	�%�a%"ʆ��nA$�we
�b����i�'Āku\� �ܪb�»�d��m!%�4`��A7�m�Hו�N���Ntv͘�G�(�\�vzk?���������������$�r�\�	�7j��zޥ�.��$�s1Y�����)���Mϊ��^A�N�qD�#z��'Ăoq�N�nУm�Y����q{��OV[P�ͦ��M�	 �ݪ ��}.�w����u�I>=��} ��f��#��z�A7
.��)ܭ��u�{\H�)2A��ڢ�ɥ����_L�r�t�ɮP���D����S�� ?'��k鸺�1����g�vv��>$tdғ�h,T���4��<^�5����H��_�ޢ��6�w�cw���|�;�g�rV�����4�v�\�=�~�����-?ߟC��x�{��l�.�l������ܬ�{r�%�;���]�<s����p��X����ȡ��Z����0�Q�/�q`5���2'4�^+svcfܖ�Y�ڲN�Ҍ�olg��*bWr�ե�z�����lv�d6�v�ex甎먇n�O< p��4�s���mʙ'�T�
c'E��ծquo,���\\�Z\��Y����YG�n���[H\!�옭��5���v��<[��8� 惪�ѫ�����p�x��_�ܬ�Ʒ{hQ$�tdҐo6nB�6�ܭ5ں`Ef��}n��e��`��UЧ�|�i���n��k7vh�}ѓK�m���6�����#�Œے��M�gf����E��H��t�&��f� �:2iI=8r�mCD �M��|�q�:��#m�n6i	'Ʒ�a���L�U�x��A�a�0\1*;)O�$�b���Os3�}ٝ�@�=4����W�z�������ѩG�BD$�Em�г{Y���{4ic9u���s����i�%������_�a��8-H�n{�A ;4�	�s�>)��qC��/�dn��P$n2���"�q�R7Nϟ��}��t��9#X���>�1Z��闫�[Yy�˜z���Ưf���C�.�n��䋷]vh�8��fJ)s�N6������� �Sw?A#��iI$��ȀH���o��ښ���*2�`�X-��{�N)�خ@��IvcV@��gdÕ40:2iI �kyYU�Dj(����[y������R���{ă��ԒI>|�� �wf�90�p���(��$���a��6��������z��~Q�"�.&�I�VD�H��ڣW�nz3rJ��|�	hYf�ƭ�ǁݍ�B�n�����|�Cvl4tt5(�ћ����6(�F�>Q�JI�$��|	$of�
ŝe�5��Tf�A ��>ڜIQ0�0CNT9k�Azz� �>�d�5��	'�������D��*k;�ǆ����f'��H
���#w��Ϫ#��}�`5'�{޻W��ɦ����r�b���`^��{O���
�K�e��OFI�q�ځ;vU'���<��B/��)<�L��'��;}*�<١��D�U?���9��O����\� ����P6��RPJ��׺��\�9[����UO�����$�te��T3a���}������.(� �[r
[�T|I��hmj��ct�GΈ�FӲ$��ݪ �Ri���λ8��W����g��͊֎�aL��C���v����|�۔Z$�h����|�j!2m_��ʩ�I����<rm����;x��Ȁ|H��ڠ	�]ÎlC�F�$�q�H==7d6ߏd���I$}��TI#�&ԂA�#,��5|!]'�FM����0!F<��s�ǯ��J2\����g>&��*� �:2mH$ȟ�%
P������>U�ﵻu܎[���I���@����R	$�W�"ϖ����k�R߃*~t罞�X��~�j����5�3�b����;��,�6����o�|8_G��{��D��o�Ο�?:>E;��w��8u�����-��}
qI �~�V}z+h �h���N�M��>����b+Mw�������Ļ-=���z�qڝK���Ic�y����Z8����`R������������}�)v�Q$��'��vgƜM�鼮��=�7*� ���R͜�!(a8~pۢ}�'�����7"Ȼ��}��I4�	��ȏ8�Ov��GE�Un�kbF0\1�W���$��g��^i���5;M֑gf���H5ܼh���F��1��뙛ݸ~��nEА�p��>>"�]��;�v�F�����T���$��k��f!�-Ґq�ـMv��N��]�TI��1}�H&���>'{7j� ��kpD���i<��В��>������E^�e�������|w7n�6m�\�cƷ)�{_Ct���/���'�'�Y]�(e���H���}75����p�[�Gv�MiWwڕ��]�#�={dl��Q�yo-���ȝOz�L�O9O2��3�tE�Q>�@����`�{��f��e�]4���^�Ll������nu���/	���\Z�ۢDAu�mjS�Z4��+D�2'�ߍU6e�I=�A�����֝�n����x,���4��� SU�T�ך��^�ŗ���/.z;r���wtf���q3�	��_j��\$��nU<߰������Aǘ�=}f�6���X&{�{a�M�\m�6�C���v����	�����������'{:gQ�jه5�ٳLȼ�3�zY�'�GF�����{�I��	F#�_]��g����.�����_r�~שط"p��!�ʫ��/.�z���7j�T��5�צ)�6���E���D��`�ʄ�y#���f�����M:�t����ok��W1���zV؆��q8�����h���q��7��{o8OB�&���#�/�@RˣO�i��˸zw�nW/{���s�*�JR���90�3ovx=�}#�M[&���*�vy�g�/��J��OU�.˪0p�akK��{��k�8���-�K�`c8�c%��>�ν
x�qۼ�>���&1�b�#Ju0��d�D���=2{X��.<N�g�ݣ�߽�]6>5TbkF�Kkh6YmVҵ*�ѵQ6�ԭUٳ�R��)�E�����`�d��E��Me-�1Uk���Q��Ȫ	�Em�lX)FV�[o	��(�F[PU-h-+E������j�#Z,KZZ%[m�*9��[cRƥԣu-��Vڭh��[
��2.��Um�
1Qc��-(�ˑԶ����ntjU�D-(�eQ����YZ�cJ[[l^%��j��j�+dQ�YF��K"��h�*�Y�u�iZز�փq��%Pm�(�kN[�R��L���6�����U�`�R�V�Q��R����lcmXZS������,l��5���j,��U֢�[j��v��.-�+m+�[��YZ�UTSn�cq�������L]�]�g��v�g��'k��<d8�a�WO9��m�e��\O����ǌn��6xS�0�#�@�d�%l�o^t��7����8��q�Mluu�y ���Z^q��%�g��c���뭼99'qm��z�ѱ\��1W]�)����Dn�^�m�r�|�=rm�9eu�W����o!��Ԑq\�q�mg�ɑܖ݇�㧝�zس�hXNx���0#�aʑ1�c�S-��Kv�,�^:��;LQ��mڝ�>�9Wn��xm�tY��pW.zG��|�z4�U�T�����F��%Ɋ����r�7;�Z�-�g�n����aZs]�v��Y�zn^k����yR���d��4oc��0S֮3v�g=<le�v�y�[�h�N��v� �>���n�u۝��Q�-ui�e�lq#��f.x�.�8�)0v�����.��s� ����<��퍅�U[/;��\��'t� ����Gnn�d^���t��E���:���
�R[��x�Է<)���v�zc.{���J�k7Y�p��ݸ�=�s�,<$U�z�k8��ō��+A���.��n:�;^�!���f�IcˎqoK�{�]ɳ�u���J�r
u������ű/	Ҏs�����I*6�ZԖ5�t�(�M�f�n�q��wg�^[O'i�C��1���`��Ԟy���F�=����n{f���v��s<�#��-�d�t�����a����˳N�ݵ�j���&�q�Ziݹ��ς[s�\��h����m�gG]'�[H�W��v����f|���@������<hq���G='���B��@��0�z�v��'�h��&�t�nۏ6����niէ�)��
sۗ-���r���l���q�q�[v��]7J�k����a��&w=n3h��RW�q������ֆ��h!`�r`y��]�^�Zσ=��N/5ݧ�T���lve�c�]0��u��=][�s�C\3����VD���V�JF����0�������d����Ӭ��za9�1��M�]�=������m���� �n��ƙC�<�Ϝ]��a㭤��cx��ou�y�mnK��u�=K�qvZ���`-���v�t-�ib�x�T�vp{�p�<�=d7�gӵ����#cC�=��/7Qss�ܘ������\v7�B�j^��Ŷf<��#�b�`Xv"�2�͜V*V����r%�'/GV�tV�Wv��f��9)ڰ�a3	y#7�F��P
�h�z�N)$n+���ݟl�{�6��=0H=ج�u���,�Yd�[b9we�ؙ��/Nf���/9ِH$wf�P$�K�5�j,]��č�9l$�	���W����A$�ݪ ��<iv�b��� �r�\�'{7f�릣�
Te���=���y�.e���|	.�L�$���D�)�:HN�E-Ҧ��`E��#a�u�I?r��9�M��ԇCTkē���(�v)��x���>���2!Q(�BAQ?D��V�EŶ�a�0ۄ8����k�ݭ��]��Y���}kC�hAh��oVϠYݵ@��q �������'�w�o�O{�d"�cwf�8-��Wq|+�/h��Mn��W��(qʧQ���[0.M�\�vcȚX�dq�4v��T�p�=��A�U���!���v�����{=�v"���5qy:�%�[C�����Mj��On�� A�ئ��j�M3ٹ5*z�ge��%��ݞ�O��MĐA�55��Q���ӄ���ݪ$�D�I>ٳ�m�6�>�3�w]�T�����j�.hA#�MĂ|I��q7 ��vumP'�v�cBF0\1+�TI�v+�C;U��^�@%UUU I"�MĂA �r��.����/���M�N-�]g���uk5�g�h��Z������<u�Nh
�ߟ�����z6%�����7O�&���#2Z5�E<����sT�	9P��S�hAh����Jك�t"*�t�T�v\�Q� �� �A��s �C�3/4�{;\�'���
@��03�'u�A �~��K [�Φ��]��*�.`����-K�:g��iOz��.w��z�~��y��x�i$ko��+[�y�'��N\䂁@���-@�ɻ_x{�x�U�ٴ$���r �K�����������dUR���g,��M��RI$�s�>$:�v�hP�2�$tu�&ե �h����V"'���z�lQ��XL���� �ҧ��O��+"�O{����룹��tA!��CTvEݧ�;y��:9�l�S��;�-��]�k�*��
�!�c�^Ґ	$�W0Ao�j�w�A��9��
��T�A��Q�m�8b"T�ǘ�n`�r��4��A�,�ž'ă��̂��v�.g*,�{y�ւA����nBE�����A&��k1�f�y|o�*$�����ݪ$[;F %�\:�Ч*����,S0|	��ݪ�$�ѓiG#�L���������Yܨ���t�bN�E���_������sᎎ�������A�x��S;�|P,d�Z,ѽ��y�������O�*�^-�S%�m��Kﺨ��gfԃ
p��ڙ�����{-�I��ڠA�FM�Fr��B����B�G��e�ۯ�K��n\c�s׌<M�pu�Ogu�]{\�HO2�5�H6[��6�7�z	 �ݡD�	6�X��좇1ST#���]P$�w}�0��D#hF�P�Z�c���6�H�ո �H��f�#ǋ�S�@=��U��dَW0E�����-U}54H��R	!�Nfۛב��d��=}�TI>�yHH3�ֶ�a�CE���X����DC�4ev$O�9��$����I5ܫJ�����˞p@$fOfa#��	�d�DS0r�]$��GO��2Fܓ7��^'��=�>$�]ʦ$<�1kT�'��nZ���S���݌>�g��޹|�C�}{���<��O��,sǫ)X���+p�W�2�>�U�� ���ʺ��<=�{����{g����.d�i7	�Q�9q˦�ex���eg[�퇕'l<-�r�n�vs���ѐqi�<Y�dz�v%�n�s�]�a�]w=�������Û�N�I��)���;g�o��\���"�ip�.j�M��s�n�u�;plfC=��věhn�������&x'���q�֧���s����ӣ�9��V���
���tnG�S�(���y� .����˓�[(�KΞ���������Լ[6�*�eQ�/iI$�]Ό���2�)}��I>S���ð$̆DaRLr�(��+��շW7@�FC�R	"��H�UMN'9���Hj����b@Q}J|	$�TD�r���N&���,��)�|k�T�#FU�D�e���ǃ����;U��H Qs��� ��tg��w�v���zL�&�"�=BA��v�e��Z-%'vVH�H5��U$`��"�=
iH$����	>��گx�u�c5ŮW3D�����@�fQvm�ٶ��q��:x��N���
"�<�������?D@P�Ah��lK�� ��	$�f�Q͛}kz����P��$��I&�L���)���m�\���1�e�]g�J~^��0��5̞���پi�n�b�o<�f��I�x7��@������>wE�y���Շrs~q��:�51z�^�� �����A7��ω ��f�Q �:��>�,�nF}y4V
-�ft�7z�v��|L���O��M���M��p(���@$�f�Q?����([b6��
�b��b���^$ڥr �M���x�O���8F{Pf|�B�|��X7<1�0$�%���z� �[yy�e�]� �;�v��zR����c*����ͫ+�k�Ƅ�=-������m����wH(�U�.}���P�^-��ܬ2	5��4	�<�&�Ɠ�{���i��'ӻ�ٟ����HH�.2"y�+5�	�HG�ĜRZ��砐E�v�	)
x��������Oy�r2�q��2K���kă��)'Ė�=������H��]��u���|^�bak�����2l�[�`�;oz��|�	���{Nˋ�RgT�}�$�EG�x <'�����mQ})	�+��-�fu@���yǴ��kFmA���@�.R�O���M������,۪'�j��hA��U�A��S���F#gA"�o*�I>�}JG���T�=�h�2��)Ï%	�-?2KF�h���=1�����is֨W�x#�<�Z��~���"BQ���Ǯܣ�v:	�s��h?Uʸ���O�3	?��$uun4��f6�߫� ���c��*�ꚿQ�/iO��]ʤ@>&�>�[:���ۜO�;t4$m�<�Ö<RI|�DE������Z�`�m����FB��-5�p�`���}��!K�O����$�|H���ٻ<*����ծ˽Ӊ=ی���h��̛���m��>�U홨u�J~c�gd��Q�v�\��;�V&�ӂ�G3���󜯞� }S���w�g߽v�F��n0۪3?*2E}����0������Ci�H$g*�G��vh��#U��!W]���
W@l���D�%Մ}���\T?���b�V���sh�����&�v�c�+]Q �Gv*� �G_n�w"-��%��Y$nr��V*	��!��� ^t�Qb�͝,�p��luĒ"�� �u��W� ޷5��A�=qN4�d�\��L/�IH=Ҳcݹ�TI�.�Yb�󭘢|I��S ��۵D�'g�Yq	� ��Ԟ�fb:�"���� �u׵On�fHM�U�h��cǽ?_�����c�($L�����T|O�ǫ�7c�ڪ��*�ْI���y�� �����Uy|쬍Y��;ܻL����G~�}D�#S����؂��ӳ9�������O�	���Z�$B	M9ʤ��-����<=��|��wG�n/R:1����n7g\��>�.70i�ftj�n	��>�l�]s�ۜ��gw�\��㍷ƀ8{*�z�3�|�=�!a���Mۓ������4�{��`�GU��6q��m��f���{n����v�Cg��$��O&��l�8��3�l��׹v�t[�0i�8�ƚ*Ǝ�ǔ뎺�ٴ�vy�,烯N�瑭v����
�8v��R����l��]ۗ.R���@���s����|��RD�p�O����P�n0ۿ��کI/�j�$�ǆA�eJ��D���L	ݻB��6+I�p!�2�]*�f{'�[���� �[۴(�ņA>4�0��X�櫹n:'�R&! Ceê=�5TI<�a	�LD�w��i<��"A on�{�+8D����I�AL4���J�zc)]�w;�Q|���&��`�"�E��;Fx��U̞�eB$)�/3�N4�ă����;A��L�}�3�(��+yT�6:��؜	况�DH����l����i��K�^pt��qb筌�`suu?�~�tZ��m�1�v�DA���	 �]Ό�U)X�#���Ӥ�1��'nh�&&��6恙�S�������z�t�̈YW����Eލ�[��YI��uS�f�|?gx����<���m}��l�4?:71A��r��w�5��$u��zv������w﻾�~�UT���Lw��G+�0���q$W���|s�T��^��>��gj{so�g����G�߷}J�㯞�k�N�`o�<��%��؋�OُH��Gv�2G_n����;7!e2�i�$��!CiA��C��� �۝�QP���/det�$'N��U��6�v��o&��ܹ�iA�&��CH�[�Ut�R.���3YX�t@]�Byqu~~����źP�[�M�H#/P`}�ە^2�'}ݜ�k
1OJ���㹉�"s��p�@m��m���j��n��Y04ݦhV�ĂGWnU\D92r ������TW	&��6ꁙ��$Nv�Q$�P��v-Guu)F�k���h	���B� .~�^�ug\x{Rtyeo�4O�O��X�Һ���օ�V2e�}�����Ǹ{�����Y�?6V�/<2�p5�>Zd��R{Z�j�{���lm�ۼ��������A����"k)�H��:	��#n1{&�֝��NH�^=��<��E�C���cK��Ҋ89�U�p�g��N��.|�+�7|����N�w���z�!���$������w��/=�	��͓��(-���VhD��}�{�[�wT�N��<;_�rnC�&kv��~wm�y�m�Wn���QL�����5��o7���ɳ��ـf,��>�ɷ%�Rߔ�)�lFb��9]�_C�>s=��Jf��l�h]��f��Q��1Q���.!tQ�$���է�}���|*Z�Gw�θVw��FhBVNh�M)=y����^�|��ND壺�ͱ�0�K�q!')�ƫo��n�-�\��"n)��J^s
��q]��n Lk�^9F{|�H�u��7��-{n�u	Ӽ%�x<
263�$7�Z�Q���ل������V�5 �gL[�˂�{|{�g�Y��b��#+;0K��E�H�D��_Tn�W>>��ރ�E��Oz��!ͪx7�b�t�[oi�e�Տ<���v�{w���e�|5�n�L�c�Ǜ����Tj�CJ����;��|����פu_?w��ֹ3�a�!k�R\�����Mƀ�]��~�+X�r��κ�(b�m�?�E����mJJ��eh���X
(�PQ���TQKJő�i�P�-�Vf�h�E�-�R�¹+""�v1�QW-k���VK�Qcb�0�%e�DZ��-)F�D��Qژ��UiguЩQ-Dke�h[kQ�X�
�m"�VZ���B�9a�%AZQAF���Ѵ�m��Im��Ŗ�U[[TDEb5
�J�Q[i�,(�fB�4J�����(��0����"�QcX�UEF*�эZU[lm��,QV��Tj0X��,�5�6,R"
k9��U��ʭj�[j*�ҋ�QY��"�Ȩ��e�b 4B�u
��"*<��Ҕ��]iJ���[F���kEX1b"T�T���
(�� �j�"��(䪬D��UV�0g$QGYU�d����8ɄSjoa!}���V'߷�>��ϝ�)��L1���aH��];j��W��. �m�8$�ܪ �K�n4�Mq�"�,�k�B.	�ˇAn����J�>.	"�LG�W�A��ɢI�FM�ߟ��������?�� ׍x�K�Væ��Z�ɺ�{��v��2��t�~~���ء6�ԿM�K�OVnUH�t�2���A�[w/7b���Z*!O��ٕ@����PטpچJ����A �[�`����A$�n�
�K� �Mn,쪻�f�ڌ��(��-��v�H=��ω� ��T�Æ����I��ʯ��4��/�I�M�$���Jqjӫı�)�\���џ�+c�\��I;Z�t<
�D��U{4���7��5e�vn{�$q ��dgy<=z{�/12��,��8�3��5��w��g��	$Ǫ|���;;?^�.1���M�N"G�$��1���RnR��;sr� o�Q�O�5���!�������O�'��G��7O:�h���=V��[D�&�u��Y�2�(��!���!�e���w�S@��*���j�wc��.wlVM�Q?�#���I���
�4I�H�~U�=rfle����w�$�td�kc�)�[��N��cr�5�6�����8H$��8 ��2,j|T>��H'�f	$�񟂾��Fܑ�nA��rUG]�ꁛ�M�Xd�A>�ZC ��̬�U��1Ll��@�ݙ&���&!6a�D��fc���ܯUŜ��C6:�I>S���A��q���̪񎻄���R�::^�f��d�T�Z� �ٯ�w'�����˴D�y��<�n9�a>� ���89�����S炴J�T��[�NNf^-�~�$�+�)�ѼԹ�.׃�7ދtOFԇ�`%�6㳷\P&����V�#V�7��p�G'em�ܽ�|lvݺǍ�Ӭ�{��V�i�Y7V��\���Y�n�;�����"�8��,`Z)��&���v��kt��ݡIWs�_;w<n۱��[�n�����ݎjm�i�m�O1���8ܳۘ�eT�
Lv�\;+6c�8�h,nl��u��h��ܪ�yu��v����Z쯄\?%&�n�8BD�m�؄�>W����Ntc�Ou�Ux�Z3�e\f�Y.̒ގb���&\:�̉p�)��s6��� .�H'�יT	37yr���=��y�p��m)�;�,@'�7+�I�����!e3��n�d��̡^���&��p��&*���ZRn�ZUU$��G8 ��ەD�w�ё� �.��������d2҄�I�۟ovE�Tg���<�ٚ�J�t�+���̪$��td�q��py���
p������pQ��N�ۍ��gDl�[[x	]��8lv��.�oϿ���6�t��L�nMN��"
#2��T<����5���';�(WEP�`m�o՟�, �*���Z�۝��k��G�s7������Si�Ʃ���L���X������a�݀�ݔ�Lz�<4HGqws����*4�W��{y��˃F�C�dK������.Q��Af�U H$w��ω�u��ƍ��fGP�!�ߘa�N�a��3;�xh�{��Y�V��:��$'s��x�J��81�a���DϷ�َ}{7w�\I�w"H$d�2	�[�Us|�����+}y��`�,1�I���I�LUj��H$���66f�b��vMn0fr�h'2]� �Mts��y���]<:��7}{��#B�J��m��m��dT&,���<69�����s�v���|�}��bs6��Ɠ��*̓�I�\Ys�D�\.oT�wR;��nC�*#�u*6� �"�$��:�� �u��>���nv ✖$@��$�,�oI&��~6��	r�@S��L���\]L�Yi�X���_5�ц(<=1\U�����ѱ�+]J��~�ȇl[�U��$}���I��;_��ws�������GM�0]\c�+3~ B_;��e�K���oSUi{�}�|�3QQ*��\�v۝��Z�Rp 4W�� �VY@݋&�I�J*�o`��No�	�z�EE*�*T$�a�;��>����|�6S���}o �T�K� �4۸�H;��[�]$?nŷ(��/<Z2 !JB.(�CV�OF��sc���g���:�I�(���vzk?{��?i|\�%<:���D��_Z�I!�mӘ�=<Y�V�[���PI�ˎ�
#ʻJ�ʆm&n�6��DD�Ij��a[$̸7+l� ���l _8tͨ��^�����H*D�"�$��52�VK`HQVR���z`�Nds������D�EQ��0&�l$�*����≬Jo	��qW�����y-�=�9����.Ȯ��.��+:mė�qWgs��J��d�e�|��u�oV�?v��82�HCTıP�tF9�O�����x��q�t�Q�㰉A�Beã5���2d�S��&ʛ���Lg� �w^���o%�	��9�����jv?�!�7c��:g5���ˋ]r�I��m�ùB��@1�WN�_�������:�o��qt�w�d�a�Ԝ����9W��g]�$���ƑD(q�S�O�4֐H�TS�������S$@g�dۀ> ���@�Nm@�R
Q�>QsJ�4Xm�L��Tu�쿘�aNn�fc���r:�:oǀ�>�e乖�w	��{�D�
8L�d��+��2��-ߵ�����9.  zu���EO��x4������	!�Rl�e�˅��UϨ �8ˈ�ŽU<o�F�o��`@n���D��m|��_�_�U�aj���/��K�H2��r;p�:�L^8f;|�����.��8ً�Jb����6��8����D���~�J�VNR��Bn���~w�����m����)�,�W�ܷ��v�fe��v7n;5Qm[���s;�dڼ���U˶�d�mV�n����۞O)F;g�2�q��;�]���p໮n-�c&R����{kCs�X<�U�:O<����l���Ks��{ c]��G[=��c�o�t�$�:�ڹ��A;�z�9�m=�.I`{0MtCӣn��%���&��Y�≠���j�ԙ�%���&�n-��%��v�)�,�kO9,ֿ{�����y�JP��rܿ��qNn"� �s��~>���K&{�&�m�sH�;�������T����0��q�w���K�,i\�C ��NK �u�$�F;�Y}�Gv9�jg��T���$���d��O�� @oA'du��ܵ���������O�E�8[y
}0�-2Zry��l;9 b�����+�q@ C=�V'v^K���6$0��ww���Pwz螀�EM)I7r���� �VM�Ϗ�A��f��	/��Q5#��D`Dwc�4"-ͷu)u�[��4R,����x�C6X�xǅ�����wǵ��N���b����4Z-�)��FB���=�� �켖�1��a��"
B����$�}��/�Ή���1JK�U�0��Gc�3��g5��j�J�ӑ�+W/n �Dn�yt�_<��Q"G!3���������X�zv�{���ɪ���H,��k�ڷ�~ x��p�� f�X�bɹ�/x�结�L7�K���8Z�˓&�=�����&��L�3Y"GU{�?�d���]L�@�y-��3��"�E$INN+'x�����	��ۈ�D@ G��%� �Nx���+ب��گc����Nzb<�l*�0�l��i�GLΚ�`=�9�;�9�)󙾃z@"ǼӀ 6�dۀ>�9�"�=�O*�o�s�/T��	�&А�p�"�r��7E� �����o�
&5�TPG7w�����jU/~��݀@z�d� �NK��$[5�C=�{�&d���%����3��*�J�������^��	�y�پ�ۆ� =x�m��q0��������m�O����xE�=�0\T)��W.η7/���)��| -���4���t��$�U�Y��x�`��ٖa]��ڄa\�u^�ӷh��з`�U��2`3x��v.���T��[�r?{����Z�����"6y�j"w���Q ���L$
M�L3�m��Vj*�z�-� �zK�� zg92�4�:�h�\��ۗ2Ι�t��U%RD���!l�3a�7��G��U��W�F'{-��o�tL����m���ԽsE�!I
�pc<��Y�QAn�+��:�PP��9"$��s����o�u-�0�l��i��3��* @|�$���t�g�v�ۛ����v�p�pڧ�i�
�c�E�$�[7��x]-;WF�W=�>#���� �sqH8{�M8��N�#.��UR�H)KLZ'7����j�D�,��khƘ�j��hDG���
	1������L�'2�U��ǥ����g�.�ɺ&@=ڵ�� �y,�6�j�n�=�����m�j�[˝��٢��1��C�5�a\9�.j�;���N�cm؜�:k��N��JS!T6������E�t}߽J�EAT�i+L;��� ��Kcs���� SI�����[�O��w���Δ.旴p��|w���ѽQ�c��wE�׫L�hF��\M��Q�8�#9�.���}���$��b���*ʸ�  3�\� D��[�у_�-|���,x���_�@.�{U��J�0�-2ZuB9��N��$����N��WX� ;����Y�Į�R�2p�m�p�)I6��â �����X���w�ʞ���'����$���ӏ�#���eR��H)KNG:�<���� �su2�s��� "��^���)2�9���]���0�N_��ۗ> 87�S^W��j�]s�G�� wZl`D��%�� ���R����=��w�`�%D�S#]�h4Ti��o��Ŧy9-����v�ۃ��g��b�Ƿy�q��x��Sw(^�����Y5:6T�"��:Yv��0���.�Xb#�㲳싛˙D�R2�UQ}ӓ��Ba(C9���EB������$w�������X�h�8k�z��{��j�钾���K̉�T�8zgU�<"�乯�u��h��o�u�9s��^��x�W�v���W��[����������MnyۏNIZ�*��x���-="ϗs���0<�Ys�<�;�J���Ӱ����q�P�/������f�a^����9��FОz��?{����ak���{&�Z�Q.Z=�����P�%��W3߆_{J�I*��G�}*�Sd�^m���L�����{�g:�YY�,��Z9 �<<ps�`�:���Ux�2��a�#�"`�,���=Gw��]x�u%9sM�C�<+�e�;�3t�mZ���l9G���8X��{1)Z�j����n�����8��a�6֢�^C������ws�Ƞ_��a��Im���E����9�B����"�_����_��n{zw�`�mO�)/�C޻�-C�P!ǽ]��:NVd�)��Z��pgc�`����W1�v��.�s��xhy��˔w�*ڛ�W**fli�j��1�UӺC��Ň-]���=��{.��f{���V<z B��?A���NՅ��K������3-�]�~�w�j}�yo�5�r�I�l��J��A�VB���J��J ��ʊ�V
E`���"��Z�E��3j*��V3QaEX6�U_,��q�)yl�֊�PU�,E�5�#����l�F)¦���(,E���1����R��ڶ�U���dPY�DDC!R-M��T+P������QX�Q���-��9�
���VBů�`�S6#m`�eB�Vd�/0��<��M�"*�� ��Efk+ �MaD�U�J�"�[Pբ�l)��j�%��m%b%���m�,�Q���ֈ�ն�DT���
��V�(��e"�6)F��]e�L+ �����`���Eym���
���%AAdT�F(�dQF3��.P�(�%B�V-eQ�b�h�+b��N&L���*�E�B�Tvj��24���o7d�����8��r/bR���8C�'��{;v��v+��c�h�s��:�Sێp1˒mf�놻�]��<����Z��8`m�>��q{v��fP����S������=��{\���{m���5q!��0�n62v�LXy;{D���t���ˀ�x���c���l ��n݋���:�����Z�v�
�t��/�m����>Ę3�y��9K�E�n=u�:i�z� ��c����p�۩ס����[�S|Κѻ6#kuw�q|�u���ց$�9˭��ܖ��i���<��a���GWnN�;�7��s�ƞ�g�;n��m����۞2v���k[��I����lggi�21u�nx՚�d����ڎz3��i�7<���@���Ӗ����6�-]�v�Y)�=v�iq�z��ک]��^������W�U�e�.4gn�%�u����Dn�B;j�}C�o9�F3��7��Â�=��^L�<<3��ŕ�Z�-㧮��YM���ڹ�ݻq��^2�����k��t�ng:�۳�F���b��Ss�g�;^�kR����Su��R{v��;u��}�<)Φζ�8$8�tO��n���[�D��ea�:�%��v�޹s�5l�#���n�|:γ�O�5���i%<ݝfy���3�6�vh�t1K=���3���������a����N���;��6��X�Kl�w
<�kn7��w'@��5�z1��*x������#��8�!Sڍv���3�^�����In��v۳GSx��P��E�ط�C�6Oovz8�Y�孕q+�n�,�8�z�wn�>˄���9s��-�*�A�nq#c�>7cs�l�gH���=\M�8�.�]f���;r��m���g���Ψ��u��[�ٸN�:��{|ƾ|�m�z㝞�đqٛq5<\�m�Dmqv�Y'�Wk/;�V�����Y�(Ż�:D\L�U�������mʄo�;���s�jۓc|��y���Kf��܌aQ�㎚���v9K��nՎѦ�M�����^��m�n�Ti��z�Z(�R��n��%���n��8�6ny�xG��l(�ݝ�ld��a����e޹�۪�v3�7t.�۶{�t�۠�����ܻ��Ȝ��mv����K�<[v�>��Z���U��j��[g����������qMnɝ�Ƹ�Վ��T-^�rZڄz+����뎻v�-j|�5���}���:煪i+_�˦��3�ץ�d�6��UD�G7��}ή�� �w�o�#�n8�Q4[�����D�%���U56VvM<�W��O���_�� ���$L���6)����j*�Ψ�z��a%*�ʥo�U�M����ު�� �=�]9�ۗ���2Gw����QޫA��.w�IIB�SI9��\`������/�Ug��fn̮��t6�wB��;3������Za'4����F�� vmm����?=�1;�s3/�(�U�$��̮�j��$����Ix���*�m�LsB�e��l��i��a�	C#,�R^=�}��)��/�ܶ�po��|����E�M�����s��r����p�e��)�v"9��L��@Y���i�y2�����6�#}�L�F��G\�bM�d�:���k�1��bKH�O�Ì�ݛ1�������DDU��f������ g}��-�3�z&������TOcH��Q%%RSBʴL�ӹ�Dg����c��~�� 6�up� �õ��w�%BSJRS*��:��g���}>㢲 �,��3�f�?��9�s]�_�d.��m\ ˌ.{䒒�4��s7�{" �z��t{ů6����U]꩛ xw6�>x�����f���ՐL~&ۋ��q���7�N��)�ø-�<m�y����%&�n��9��	2�Bf�CQ�� ���p�3��p
}�z���ހ%���E$��˻ϡ�!�%�P��9���q�.���Oу�S㼚&H;+uӀ �yn\�
��<������t@"�JU��	&�n��q=^��S��fs��z��j=Y����������sU!E_^qyϦKQ��u�A�E�>�8b���#�c����[ScSple��� ���ö�Z�""�˦��L}Y4h���TH�L&ъl8X��s��ج��y: ��uc�D@ k�r� @q�g�^220H��3I/�_f4�٥�&	�As�w��>9��9��*:�ݭ>�]dˀ7�n[�" ;��r�/+(M���p�KREd���&���㱻<xy�9���T�n�83g�mr�<���}>��Ue,)����+��;��` O�W�Tm�<T��~-]kqD���r���4��.pف(���9���yg��Z���=�Nm���y_ȒTvw>�S�G�;gT�����{�q$?.��O��o����su���͸�� 8�+A1{�S��Pm�\�	��Ě>ݞ��	f;�����U`@vv�w�^َRJ.��7U���k&T��>䒱��jk��.�'҂�(t�������cZ1G�r܇@x�q���%�z=�ԇ�k4g/Q���}�� 1��/VtI45���U)L��IM�-W �{�����>���{C:��p��S6A�ϳ���=A�~�޻ع4J��m�S=���'bUuF��Wc�q�L�])ܽ;N�yŵ~�w��-��a���[s�B��M�۟0���������i�c��3���6@L�W>���s�HJi
EBN���O����'���W�P�|��=a�|��Y��&B����2c{�~vt��T���&B������hd�@���@U��oe�g�ϳe0�|��D��%q_��ȅ�(���t�IP��2���~��g�q�� A�ϲGۋz �|�]f��DXz�2J�I�M�{󣤜B��T�
���~���T��~�Ӝs�!Ȣ=|B>��(�����{Nj�#��I�Ƥ�y����t�!�&C$�W{������T�
�d30����d<g����j�s���d2&L�t� W��>U�%~L �h��:a�9��~��x��IP�1�f���6}dy�t��'&���y�!2m�<���N!RT*J������y�2%B��߽y�YT+d��Q��>��L%j�^�kSxʋr�	��C�~�r��2�-�:�u��o�bo��w�![�;�j��[��Ph�nuy�#������ㆺ\l7����ېr��W��s��wY7n$��K�Ә��iֹ֬V��k8���:��
�<����/���/'Phe��u�S�G6�v�6τ�r��I�m�0d��o]����V�z�gg���p��q�[�O\W&�[[;g�"��M�u�:���J�v㋱��A���+��]���]���=i��扭��.���oNcD��c�th���Y���.K�u��E�W!���{~����p���C�x��d߷_�:N�!��2�3!�=�޺<g�d�
��Xo~��^!��a�����|�C�O����{��'gT2J�d��3��}�YDy���VK%��l0�	#�AX{ξ�}d*J�yW����^�r����^�:���Rt�ԙ����߻�!RT*J�g�{��9�3�Ȁ��>D@�'~�W5:ދ��$=S�R��?�9a��p(�Q����J�{��t_�*&&��}����g�3��d�d�'8�
_������ӈ%`X����޺�ܶԅ���C��o���r�)8� Ȣ=��E���_,t0 Y��d34fC>w�޺<����P�d3���u�0�r�r&���~tt��������W�����%B��|�}�L�YDy�NI�"`�MD>�T�3�}�3���3I��Sȏ���� C|�}��~��s��@�&���κ�hT�
�d3�|��<��d�
������;N��w�T~���S9���s�%A!a��Tp��=���y5�Ƿ��9�����,�h���~�a"�e7�$�|
 #�_L�Qy�d��3y�;C���fI�!�B����2�>���1�q�vH�B������hxjL��&Ck���,��DW��$�a�i*�d"T�n~��}���Y�~u��|���!��"#2�q��4�wm��uC.\���P�k��,����cM��w�kn�D��V�ll�b��z�A��#�������o������x�CD�d0��u��<a��*&�����:8���IP�+���׹��}~�x�S'�
w�+%��l6j���"�!����Y��L��!�&O�{��N��|���y�_5q�3sf��Щ��L�C3'��ߝT<g���3!��2~���G�N�ςPȣ�P�*��Ԑ,�YDo�z+���9{�q%B��V����W��g�2d�2c�9��gq;$�T�
����u��<�|l�өwM���>�RT+|��ު���!���Ď������QH�@DK_\�G���d303!�~���G��!��}��[���W 2������ʂ�9�C$Ƨ�����NΨd�
��3?������x&I�u;��8����M�0�ASi�8%�0�%��8�[N-)ֻ(.�m�����k�ߟ������:[�N�T�Lÿ����#�L��jL����G;���L�IP�������d"����B>Wo0R��p@���=��U�̆f��d2d�����DI��B�$�I��� I���Ͻw�������R>;޷��>��;a�:��g�3��dɒd��9���$�%gnI��>���]C�*J� y��YI'�GxD�����j� �a�ӄ���(����~��N!RT+;fC>~�޺<��@@�@DB #���re�:";�#���5q���M7b��W��U��}���w<��m\���Y����K!ݯ�e��)y��{��￞n�y�@�~���C��!�g!�cS����GvuC$�T��Ͽ�u�E���!Vvd�Xm��P�=dZf��z��y���o;Rx�IP�Rd��~ts�N�ړ!�0�g��u�;B��d2a�f߿;󪇌���\�S�=|��!�S�'�;�������W���<�{��:�<��d�
��a��μ�3ę�{:�{�u<��Rd�L�&�s����N!RT*J�����z�!�2%B�~��Ϊ>F���T���������"'z��5�Q�W]���m�
�V��4��;7][�T͵�������#r�����=C'\�������*�fC?������%B����߿&�|,�>�����v �0�}�ﾎ$�%{fI������]C��2L������9�[�my��J�	�w��(�Dz�G�'��Q?uVvNm���?m�Ύy):C$�W�p}���}��*x�C&C!����_<�!����@G��@D	�ڎޣY�Ȕ����� #�Eq�~��I��� I���g�]��A��&5��X{��<�>�&B���$�������{��n�������8���fg$����߿u�<C�Rd*J�Ň�z��Y�@��~0�bp��2~��S��P���8�I� #Y����<C!�d2&C0߽���<a�9�9���{�~y��2S?l����\i�3o2��HF�8
ߦ�W�DE*vS�R��/./�a�����c����!|��m�7�y�ϛ�������� �q%~�$ΌϿo�"�Dy������K��a�$�<0�����g��L�9&C�Db_�C#́\�:�یs����z�_�ϟ<�x�O2%B�	�޾|�!�J�g��d0�=���G�D��2�gmw�򾸌�ش�E�SbM�C�$hr#��n_;P��k��tAS�a�Y)	S�:�>���W���!���3߽��v�I桒T+����Y�$��dD"<��/�C#̊"<��f�_m�?���zώy���u�Rd.����+&l�"(}W(#�$�U��:O��7�tq'������t��vCվ$_��F�� 2!d3�~u�l<�C$�T�S�_d�G�`G���G�����͓�Gꗳ��a�"8V�S1
)Ȣ=�3�~��U�Gę�rL�ISݿ|��e'HmI�΃�z��U��O�p����]��y���O�IP�?~��Ϊ��Vx̆C	��7�:8�h�>
a�~��D(l���|,�?O;�k�U�#ڠG�����L�̓&L�&?s����N'bGȢ<�~�O�7�Fwê��:>���L��~��U�x?�+afp�x2�`5=!�B!����љ���=��!�>��#��O�,������s��Y�x9�G!�cS�7�:8���d���2���=���ę<��mh�D�z��Wn���F�oV�{��ǭ_7�[�y���{XĈ]k���<q5�o�4�5��_�gP��p����ВQba�
I�z�c���͑i|f��Y�e���Z֧��i�ֳ{sz�<���o[m�^۷;�*t�����2ܦEI����b����m�'�m�I�BӮ@� .�q&6;v�X�-�x��c��k���Z�lnm�`���o3�>�7L;pq[��m¿���ٷc=,��<��[t�#G:����p��ۇQp�W�y扠�gP��݁wg9��ut���u]�\u˓�3��a�^K��������뾂�a�d��I�nvQ��l�#4�!�&O�{󣝔�!�I��a�Ͽ>�ޡ�<C!�s�k}�量/�����{�����fC3�b!�vHd
"H�!��]$�E6w7}!�!����]���I����߻G�°��?w�C��
��RT�o�tq'�d�
��G>���]AdP<��y+��99���D<|�nG"�bI���b:���FI�+;d2J�~���]C�*D�d4L�a�_���u���~>�f�"� #�� "<�����'gT2J�d��Ϟ�����x&I�C�&8I���)в=Y�WOd�|��z[�>��{��}g�I��*~��ލ�'HlRd3�d3�翺��RT#�@��#��D>-J�c~�ħN��g��a2uy�Ό��V�wᯜNB��n��'��Q����
��Ry�f��zό�&~s�=��׷��'�T�4�s�{2N'bd��9&f�}��]C�<��!u&C0��<�(�Fς #|����}">�7F� �V��ݵfs<��nn���Ú��[�4�!�N���{����
	mCI}��G����FOP����*���z��3�22��{��>���r��z|�����>$�5=���FI��I\̓9�����uș&Lu������%�G��!�k�X6G��(�"͏��Y�_����L�Yt�cۼ���I�Zb/uTE���v,�By����7��@����;R��/@����hr�b͌���T]���=�����{I�������{�!SȆC&�d30��z��Y�̆f��o>����c{>'/����8�a��g�w���m����<a��:�޺#�%B���3���޲��T�
��ێ|����z:��޿'��30䙙��}��P�5&B�I���߽y����*���:��k��RI����!���"3��o��s4C�>��fh̆}��:��!�����Xo�z��yx9�C�#�_d�G�������	#�d��Q�7��υ�~!�F�c�RL�I����J�	�w�_�u����!RT*H#�]�d�z��QrQ�i�d3������<�d�
�'�y���������d0�?^{�(� #�YFlw���J"�-ۚG�\Ou�}Z�j�z����N}d�ݣu>N�*G�xk�NB��o� I���9�s0�
��C$�V��zσ<I��*h�&M�sߝ�'�2L�����_Ǿv���>u�;C��\Rd6�齔@�g�C�qV �@��[w!�y���_�2N!Y���M|���&>��e{�@��ٓ"Ϭ���
��Xo����uy�a��I�Oמ���;�d�
��}��?:�[�|4�"<�Ck�b�XM���:I�x���w��<fa�2jL�.��F6��d�
�O=���*�zۿ�Ѣ&f�i�(a�Т/�+J����aPi�\��:y�N���_�[:���%G	��+�7��+��UI6����#vM�w�n��ŻZ�)G����<���*`�v[���%�6���#��gR���\jA�r^���>}�O���	������8����DR@�^k����{ݨ˽ynK20�:g������&G�yjCn!��d�p>������M��k��Ͽ��
������$tiX$�3��4��غ�뿚%��YB��Q,�.��Ύ��x~'���@�M���Z���%{ll�W�.�'��v�� �®��¬�+.�O��TS[�恂u��aG�y+�~��Q�W>�g� q]���E��}���ey\ĩol��f�����֯Lb�"�	~����-���i�����d�w��^�9���il�~��gK�c�EC��xȽ1c�c��yf���o��j+<������td��fB�7\;I'{���}�|4��t
�68�
z��xl��q��	�o����v�����Rt�7=�A;*�N�]��w���s���H�6����Q����#d��)�$��9���E���U�O��}�imW]��F���X�Y��oa���.�=0�7И{�<�&u��k4�m���X��������z��-����x���9���!ǆ/)�6Aհ�<��G��60�`���ʶ�[�i&�yH���'0YCx�n8�C�����]|����ϒ#�J�v�)��(FJ5���Q�g���lDF(���P����]o)U4�J(��[B�E��2�b���ZŬ���VNZ�RZQTQ�#��Y�
�Ĩ:�M@��PV<B���Zł��ֈ���
�ň�$�X���q%H)�4�[j��""���B�\���b�2B�u�m�)X�0�Z���V����[ET̪&��+
�*��m���1�"��RQ�*U��J�����Pm
�,�e������"J��T�)+S��VE������µj��5��5���Znl�
֤��@����u�0X�QdmP�P�ADQEW6
�*T��-��@��AJ����W"�����R���O�>y�x�O�2%B�	�����P�%B��T<L��|��v�!�c�ϔ��K�m����<>
 "羙w'Nr�2>���@��r��cP�9�ν��&p̓&��d����;2N'i�fa�2����Q�G�����>��@K���k���@mq��I&�ǈt�!����td�B��d332���"������_9�3_q��D �2�>y�{�x��Xx9��˽�ђw���fI������u�"<�׽p:��Fx��j!�p�&�e��srq/c4;��n����.��玵r�_��-�]w..���ԕ=��w���uY���39&CjL����F����J>���}3�D"����T���rz�����y��z�x�d2J�C	���~td�B���yn����;���:a��3��|���d�
�U�ZG7�L�I��~�� Q��>D�2d�4�s��̓��$��I��>|��]C�<��!u&C|ݟ~��>k��<� q���s��
C9��C��C'�οtd����Y�����޺<g�d�
�L�|=����?Z�A�� �p(��mO���td��P�+�2L�gϟ���,�G�g`�pY,&�2Z�$z���=��uY�������}�I�ړ'˽�wI����_�~��P�
�d2d2��~u���l��w����5��]>k����ŢV!���D�7�ܽܠ�B�S���&Y��V�Z��3��)�u57x�����n��}� 3�����y�Ӥ3?�=�����-����<a�r��u�;B��j%B����[0l���2m\k��^��#�"��vd�N��&f�I������x���!u&Cia�ߝ����a�Gf�;�gkjM� �&F���u�l�[G]Slۉ�⍵��0e]��6*�7������m��>!�z�N�>�ѓ��Hffd332����ty����Xo~���uy�a�:��?3�':�_���T�w�td�N�d��2L����z�'��dǧ�:��w7m����T�3�~��U�>$��I�'�s�:ot{Hp�$,���� �T+��>��p�
�d2J�fO~��f}gȀ��� "���7?V��nNg�����2��3N18�MHw9�ht��_y����|C$��d�
���:��|g�3��dɒd~~}�4}[��G� B#����>E��f!RT/����>����o��y�U�0PP�m)�d
"��S�8�=쿻�������v��2�������g�d2d2&C0��?w����<�a�!�cS�7�tq%￙��mu�?|�7��G�^>G�zg���&I�߿�ǅ��^n��v�a�����g��&frL���'ͽ󣝔zH����u	|��{x@Ez���<�d��f�������3!��d2&Oy��w��l&\�~�䋳_�\[��N���ȳ�e�ö6Ҧ&�j18.�u��i^s�w��.%��r����{��(�O'Qs�O� #6F!qOl�y3����'Uu��-�;�4��H����f�]����`�uGV�񃚲�rm�`�:}<�
�(�e爳)07m�h73�۸{tu�d��w���D�ny|u��xɐ�j.�i6�ņ���e �ٛ�.sˮ=�ԛV��M�;a��3�E��\�;�2V8^�nŵ�:�-ƺv�in�SmW��I�[�׃1qg��f��2�+/��:����A�a�Z�c��3�]�T�sy��;�k��A:��7�lD@IC_��g��� '�y�A��&5�j��=��U��&B���$�����ĜN�$̻�~s�>��$��]��]C�<5&B��]a�ξ��!���!�=�疸�px]���!�x�N����!��">O�s[��>���>-�L��>�$�T0��~���x��!�a�d�?m�I�T2J�I_�Ӈ���=Mo��L�iDy��*b4Bk�6���g�*x	�wϾ����&B��cRd�o�ts�N�ړ!�0�ͻ�~�z�WњΝ{��� � "L!��>�>��;g�2������ߝC��!�b�<;��ܼ�Cj� 3�~(���}2�d���[�Wǯ߻C�J�I٨fo�y�x�8fI��*|�ߝI��2L���(���υ��4������y��@��2K��~u�<|a�Λ����.	��^�d_��jzC"�@�>�2������tx��_��}��Ϸ�����C�2��μ��񇃐�4r&5=���Gw����&A�~��,��"����[:Aǎc�}��}���;�6�:i��ݶ�ȯ6���83��\\\.�^�0��`(d�{gGAe�M���=�虇�u�޸�i*%C�Rd���I�*J�{�2���z��S�����#>�+��i�"9�\���fC3Fd22}���v'Hf���)�a��^n�C�G!���3�D#��G���ϝuU}e䧢S~��߳��Bxf�f"9X���}}<°�;2R��A�/�P��������Vgu.2�d�{�����VV��$��d�d�7�9��8���fa�30���u�<Cɩ2Q�@O �Ew����,��z~�75q���m��<C��9���q>!��fC3�g��u�;B��T�����ekY��T}��}V�d>Q0Ð�*}��Ύ$��I\̓ �}�L�QB#ȏ�c�FL�Rl�"��`��>ܖ}�rd|�Tg�����~gq�2Rd���2J�p�!���������C&C!�>[[,�G�4�F����WޒI� "�:��ގ!�t�a�<�~��8�y�y��C�<�{�t>!�i�d���a���޸�i+Oz�\�˿y2N��&Ov����8���30䙚8�wL�Y�"(D�=��@�`�"4����0+{L"� ��h�
��\O�����3M��#u���^�܇g��������#&�6���d}�#���Ƞ@�332�3!��=����%B� B #���ki�,�YD|#v�$��{������ԝ�s|���8�I^�2L�����޺���d�0|����x�׋���Oș����q�Gę�qD�}�'goӣ�F$�C��IP�d3����}��*y�d������q�T+<fC!����` ~{=z8���D��@�����p�i����<�C<��z�<�6��T+��z��<I��d�dyD�l�����k�l�lM:n^J¡�t��Υ�����m]�����B���T"ů�:��َ�FX)��t�֑�I�}�9`�����(�����y�t����&f$�������u�jL��&Cb���{����C=zx����X��j|(�$z���Gh�gs����������RT+ߞ��G�x�C&C!�!�`��{���@��(���P/�D���1��a��%{fI��{߽u��2i���W�n�/5��w;<IS��;�~u�;IY��
���~���r��6���~7�������s�́fO� "�m�W�� �B%B�Ȟ��z�$�Vx̆IG/�D��@���7�^��fE7���^/��l9��ױ�l�Wu�q�qpLGWF������م�o� 2=/��@���2Lj%B��~��\|g�3�d�4L�&��=���N'bd��|޿�x|�y���|g�y߿:�!�ԙ�&A]Y,�Fς #r�B��Ciu!�x!�{����w���Y�,��r1?/��>34�G� 2!d4!�}�{��퇃��4r&���~tt���%tfI�����~ݡ���ͬw>E���!{'N���O��y�:I�x&a�:��\g���39&C�%�����t�!�Rd2J�l�~~�����!���S�!�����{���3!����`L���Ύ�q
þ�?)���M���<a�(���O��WU#O]�G��O���y�}���%|�d�2L���?|��'��&frL�|����h�����t�����&3L�Ӑ�����t�=��z�_��d��D��>��,e�vuWX���^�{�F�#3.h˨4�Y�����I�#�xc����%B��;�]�x<6��u��>�2n���'ht�IP���gϿߘ�� Yg��R�&jc"�s4" $�f�{��y!�T*Ljo�ߝ$�%{�g3?�{�����E;���DE�C{>L�C�E��m�ڶ�[3�:������Gn��Z�V����=a�}���tD'ZP�)�,�A�ݒ������2_w�::6��gF�ߞ��!�xD2��o{��<Oy��q�̆fd22ow�::C�N���w�nj�ח���8��!������hjv4;荑�dtGO��}�̓�#��2L�2L���Ύ�q;$�T������<C��
��d��߽�/]�����'z�Y�| �Di�:��yͻ�vT�y�Ї,eH,?}���c;@�T
%`~����_�w>u��:��?qRT+���1���tt��T��3$�f}���C��ę02x혆��mC.	#�E����t�����}��q�� /(DC[�&�N��Rd3��w�~��<C����� �>s�,�g�l��\���ϲ���d22o7�z:C���	̈e4	����H|,@G鯘<|CĘ�2L�a�u��\|�L��&�O����#:�G��&f�I��>}��C�<<��\SȀ����K Y����Dl+�$o�#dJ깘��
Z�F��w�m��΋ͳɞŐ��D��
���뒩��-n�ct��ҾD-5���l\5�	׏��0Q�xgS\;4y�wÖ��n�h7&�g]�v��������W)D=]������y�n��1���۝�o�	>/��wn	�H���B�\�s�|���ڳ��T/v�9�m��$�׻�Xݧn8|��gg�'�h{��@�Ѷ��,:<���m	�y۰�tvYq��*6��]�^{\���]�Nzz8�:3���qh#[�^�fn��.[kuZ[���d��z���~V~�*��ݧa�ʉ������v�6�l�o������'`�Hffd332��u�;B��T<L�|�s�L�g��D|;��V�sZM�����8����GI;�P�*%p�~�zg��G���[���AIBa�B�T�Lî|��3�ę
��|�n��g�~���v���}$��&C$�WO>{����<�d�d30��:�>�|���@D	��̞+>���OxiGޢ���4!3y�R�QI߈q����_�y�A��&5��X{���>3ę��2d�2y~}��~�����Ӥ�B����33�����P�&��T��=�_~u�<|d3�� ��!��ү@�,��_)�GG�~|��{��:gl�d�
�߼���3�8����a2��y׿;�$�>
 "<���$z�$�~�ϰ�;��$�`̓8f~u�u�8�"6x�i�	��R$�QB>;��v���rL�ԙ/��vRt��3�]ܝ`���@Eml�xYhd2J�f�u�θ���fC$� �A��$
"H�9*3p|���\���~�
�*�=.Ƌu��M��۪ލ׌��Iv�vrE���S�RO�mG� i��C?;��G�8�MC$ơ�_�~��L�fI�	�d������<ȠB#��&����gF_�G���o�Ρ�)2�����t�i*6+��qpK	"�� 2,
W�"H����|"��g]O%י!���G���19����^��<�=}�+�n<���חn�G1���:�����;�,�����?�=�ȁe�=���Cd2!�m�����<r��I�M�����'gT2J��G��������|(�!��BE���&`$�0ӡdz��S��'�fa�2%K���G]�t��&@E����GI�f$��_}�>��'�22�����t�l��3!�T���tt�bt�`���׏7!(pṢ>Q���BmR����!Ę�2Lj������x�!RT�L�&��=󳤜N�$�T���_O������|=D�D�x+�>��_dDu��!��7p�'�7���'b!������� #�s�E�Y�4R�	�sJ���Ѥ q����˩ Y�	�r%K���GI;�I\̓!O}���C#ȉ�����$��D|�g<�7/qR�SdvӶ�=�6n�nYn���k�����i��w����M���H����G�w���x��39&CjL���Ύ�q
��^�d3�����p��d2~���~{�t�L���������d�
����y���Hf���O���my��x�3�}�ރ��8��Sֻ���!`|!\���YE�&�2`���;:I��2L�9&f#�}���C�2J��Rd4�ί��?g��WL�8��DW���|� ��w7p�'����Ύ��:C33!���Ϟ���#<C�a2�|^�N���͞�6rm����6�gű����l֪��tŸ��N�s�QDU�D�`�y%����el�Ke��P��bn�7q�����$�� �C$ڛ���GI;�P�+�2L���k��#�E��.����&t,�A��S��'�g4lU�y�t�Y���jL������):CiI��d3���_���d�C!�D2������EU���~� #�>DG�������@g�"gkCM�������z��<�<�M�d�PG��;r͟Y��鸠��;�2��G����Zɗ GR�S�z���n�7￧��]�u�[��v�üi�z���� ��B�v�� m8[������c����EK�����p��w+���>�g���s���b�N���V� ���7峎EJd���)��N��~�f�;���w��K���d��sL�Y~�� �9N�r1z3�9H�^�	�GL��q�j9�]+�2P	yu��D���+ދ��-�p!�խ� q����0�$ m�<F��҄�y��r�ыh���8t|�~�p$�����֡�0�<�ۯ��E��;�\�@݊7*�s�5tw`��3G<��w�.i(�{`�퇽��ⶤ-��4�k��*u]���� �Q�" �������&`$�0ӓ�C_e��D��}U5H�}�r����ֱ���~�gN�G�֤��MLϣg�'�q��Gr�6�6��7N�皻>�k�N}d��)�'Mg�~�{:��"�?|���S'��W��  �k����FN�����L���2e��_�p�$Ə�R%#n��}4DO*�����>3�l�;��33�}ނ'��gU��6���&e8p��Jp�Й��p�]����檷��߀>�W�̰��|�.f)T*Ng�WD�jU����]�z ^�i��)k�GRA#��}z'h��}�}����sBxdD��H@�.<x֭�έ�T�7���V޾�2�1�D�Aݕ��B�·�K�Q��:�
�HI�Nx��VL�ž5�oE��H��N
	���67ѹǽ��#L(�:=����^^�&�������.��C�g�{���~�~�5R=9ӻ	�'��7}ĉ7\e�#��$�ǂ%���[�5���{�Ě��c�&G�E8����ڣDF���:��W�
�����ɹ�v#mw�j6�'	�n�ڨ���hۑ�z̦��Y+Z�Z��vj�F$�ܠ�S}�u��:n�=ur� ��|'tv��K������j��_o*��<�]����?V�l�`�#=�nh�l<#��.���+rj����R1\��n¶ح��Z��]�Z{c'Y��p�Q|T�D9}�*��q^�[�bd�7V=��a=}Q�o�u���b=�=;;�@*8�;w-|��Fnŏ����%��z�cP���hs�������i}��s���53��]Ǐ�~�~����F�;�Pc?v�G��u�÷$�oV@�&O�B�V�s"�ԣo���-�d��#��5}oD=���}�m�M;�l���7��n$كڇ��}�K�yu��6`P���+|x{n��]r\g���h���(��]Z�c �7��(�[1��D�|w=�?$�F�͟j�Yf��Kh��t�=�/o=s�'��=��n"WX��׸�zE�A���y�f�]�iO�3���rD�����	���S;G^w�X�p�SY�e�&�|����7�jy���t���*�����m�p�>'�3�O*���{�����>}e^�`���h�KN["�����5[rd�[T�Ue[`�B�IPY���8<B�Ͳ�Z���m��8̚�PZ�5
�h�V���)*�F�T�1�8�,U��EU�esP0YiQ`�-I^*C kb�Z� a���Ҍ��3%rB�XJ�*R�ԕ�X"�r�(6Ŷ��V�33(ȭ��MJ�RjJ�
�YZ��TQaR��PQ-����KB�����V��,dX��Q�mU����v(B��"^Y��T�
�XT���DXJ�AH*ŋ"°�+)+MrAUUԬR��Ƴ�4���V��g/4�k��Mh6�DBT��U�F0Xq��������դP栰���(�P2T��]��7`�Z9��,X�D���|�s��q�O6ϸ�9ӌ��v�t�#�ݺ�+pp%��5���5�s�u��kf�f׌����n�z,pG^�m�"[�݌��ݮn�k���S�o,`9y�tōү%c��٧�����ۜ6�v�IO��9�ܘCaUGM���ֻq��X��ޡ�=mӶɱc{z4�������n�<��]7=��'e���<��o.ܓe���e�S���g���>靧r�6���u�u���<>77�v�v�N��ˌd�]wN:+�A�=�ώ9�Ͻlc�lOdck	�7�F펼��/<���N������ݹ��ļv��6��m����˃�\�<6�Ac����d|zMGW�9uk�o7\�qh�Սm��n�n*[�6�<h��XM쥵s����2F8K\m���]^���_|�2Z�nq�q;�����#������,i=n1H�K�n\���3�%��>r�.���ֺŔ������.N�.n].kG�NՔ�u�n�<�q�:�%92a�y����!��G��sd�'\��.{v�x{8�#�)��ǃk�íq��t��#ĉ"�jw�������V���{]��cY.{#,��
K��ct�m��2���81sDm�;�^��v��J=�{=ѻ�=�G[b+m���mv��˦�7.��*��.��]�Dzs�7[-u���q�ۧ��i�{8����ZNPf�;h<�[���f���"��$�n�mۋ��]sr��ֺɩn�bk<�NC���,�\��-�GA�pk�c��ڬ�+�E�^[����*0��y-�=���3ƣ�^��v�M�Gf#U�N]�nC	75��۱��^K����I�ܓ��/���]�5��q΁��N��0Wg)���Z�:Г�sϵ�h6Gv��*^��;��v�g�!tnึ4f�k���	bXנ^�.��籃��try��I��'=p%e�n��k���:��FClF[o<�wb6��ݾ�|�d�Ы�r-�vy{%��γ�u��h�rWF]�Zʇ=�n}c��ۛ��m�n%�� �N��m#�{uV��g�CYϘţ�귭��އ�1͞7]����v�2�8n�ɀVnDN���o��z���k�j�x�#�uOg�ޞ�a�rn�v�[�W=#����3��.ص��E�+e�Š:r�S�c�ֵ���)-���T���m5n8��������{\�6�jmnz��6�������� ��F���g_�� '�j��� �Ŭ��[*�]VO�:����p$@q�Z�;����5�d����g�h$�O(ȳ����s�� �V�V #{�($�^�tD�W�5y�d��	�O��H���*���mu�3<x}��ܟmZ�L��ƭ@wencHzuZ���%��~�j��g{�����E��D ��p��>3�s%�tW��WV�r�:��0\�!��3���&î�: *�6e�]��ǟ��W��l��f��>�K�@b�]aW^�~�~�o����7\m��n�sOS-6t��0e]��l2U��M�۱�W3�vO�@/�ۦ$rX�3�+WG����w��S6��u�@�$UQJ'.�� 6��(�c�����,��ُb�t�wv}��d��9�+c
>��-�*�G����݆Y��
�2ر��n�M�C7#۪rQ��;2����GT�ܿ � ��V��}�,c�;�G�zFΏ��LU�T�U%I��O��7�D@�r�	���i�^��=�e��;��I%�l7Ę�
) J�����������+9@�7ͩ��%�o�>�9��ɪY��l�זϾ	�3��.��)(��(�H���^ 㚴+����[�Q�9k�Ӏ" �9-c`@sW�q��p|��/��><�|$��Rd��k9�R5�n��p���`H��r�<����;��v�(J|Kۦ�U�l" 㫚� ��sTNo�6u��� �1�"�dD���l���	E�J"_����8u���\�iG{b �k� H%�쌚㷃#���Vy�B��Rp&��P�\����$�\ �6n�����i]��IC��q���{Ϻ��I�*�#�0�b��r�L�:z�o��lt<k�.8Uq��zk�]r�����>������1̿�?df��kM6�(��&%�]���>�{�z=�2�ɓ� �ƪ�� �3\ξ��3{=�:S�F��� �k�DJ���US�� ��j��}ݻ�.!��7 |���h���5�E>��{.^�[����	\����:n�gv�zŋ31��*\�p��b��L���6%%R�	R�[�y���� �բfd��Nh/���9���^cp 9����l˙�D �6��Ӵ�3mZ��uVq��<kUp q��$��e��,��>��vj�J�c	��l��%��߄I%�u�G�|:�ʽ��z�|\΁�5h���o�uϪ�h�AT�R���k/br���垭x֪l�|n�0 9V2�`���yyJ��C̩��t�
����_��������Ҙ�����o9���p��0ýq7��sE�Ԯ���Q�#A�Y�x;�DDC3���}W��UUU$�D��?�o�7��c��E����e|@�ت� 3:��,K��],�1�p���G=f��m/3~(��Ch�C���N�9|R�ٴ�-Ө�;Hsr���Ͽ�>����J���U� mu� U�����=�����D�Ƿ�����-��4�(QJ�I����0�P��1_6vx^U<@ع�� 䱍� �ם����������&�	���T��WWg΀ʷ���$[��E�p�ٓ+K�W���Z��HI�Y�%��2��Y��\x�F��N�J�*3�L�ec�G�@bYῂd��9����X���`A���K��\UR�	��
���W3!���yl��v�{}p���t�G��2fe�Y�""r������9�H�B��x�r�E�-�;�����xoh��&�]�{7u���k$�M���ow3��n�����+�U��ZTn�_{�m��I��j!��Nv��.����;�Fco�L��]�5���S�����)���j�8���k�l����Q�;J�G6� g�l���E��)2�,�x�u֭q��\۷+!�]�^Ck�#��od]m������ۦϰ��O��	��ܠ���Y��6��+��ծg^�[�2V���k5e�sm�����Z%�����Š�x��9�c���r^S\�n|�,1s�!�-��,�YW���qZ9����~*���H�RX�^�_�� r���a2mW:����|]�kqD�%�XO,%u$C�#n�_55��$��As��sr�âgo����؊In���y�k�<�z}�	8��%s�KL����Z&@�w=ы�|>�ޞ��Ի���>6�up�t�ٙd�"�T��)w/eJ袷�\�rf�U�\�� �uV >�O6p^^�6/�
=��:������j�q����(%����[p��y�^Ǩ�#x6Qԧ�	1���#�$���<y�M2�i���Pܗg�ٝm�7h���7)8�=j�'�h���ME(T�z�<8���� L��W,;��zc��������_$J\�c� C����r8�2&�_5r�99�Y�{|���eQE��]˻3tDƳ�b�\Q�!�pi�-�s��K�\�צ�+�U���/���̔��d/��\}PI01.���>��S��ֽ��q^R�Q�9w�K��]��b2B�m�䞶IԾ���a Q..3:kOz�Xn �u�� o�S`G�� �)JI6sW�����U�g~�p��� u���"�Y-�ٻ��|@�����:�f��D*V�5sO�@e��1��wG� ꧕V =�M�2GZ�f��+�l]V׮?�;����tqVh�i���N�v�Vtݶ���~V��v[\�����}���FK�̺�*9ՠ	������g���e��ImeA�s������@��a��pG0��ط9���U�V}��=t�'�}��. �����Ԙ�9�L����asURT�%$Ӏ]z�0 :�<\�>
��/�ћEeɧl��D�XY������ �̑q�e�0T�3J�}�؎�wf����^�v��_�X8��VT�㡚={�T��B��Q�b0����k���w+p@�-���צL��S4�%UM�F]T5^�"������� 3=�����[�����a�Q�@��r�u�@%R(Q*��kWU8�	y+�#}�}���R�t�Xc�r�=k�� E�Z�=�!ܞiׄ��D�P�_�$JEN��ٻ�@s����}���|�ut_����۾�2�/~���W. �˭e�ˀ#����5�>��X�n���@>�k�_9j'�)L���Q���dߟ�<~B���b�m� ����P��$���}������Won"�D#̢Ɋ�JU+�,[��&@ཫ� �1ܿG�z���\�2������'bZ�M��h�2��3�Ւ�6/�W32��c`��^�\@ {{]��`�"�����Ѭ3�۸V�j/���J�禳P}Z�ʻ�1T��az�v�w�!�L�jaC���l?��G�s��G�{����\�$IP�U7�2�� 7߹6=�o��{~ȝ��+"@w������3>��n"+��}��A��
)�,��(�Yfx��;�۫���r��t�ܱ�j�������(��B�T��i��`�ྫA ��r��y�T��IY���l� ��������B.$[iG.���0 G�*Z�r3�����z@ F�|U��nv��$��=V��SW�7kI��/)��.:�(]�@� �ٚ�0� 	ɗx�ή��x/*�'�=������S��S%L�*��f�����R���IG����:�${;mˀ>#��rdz��q��Է���'���E�Q&BuϦ������������T�L��7�x Aۺ����:��n 1G ���s�gH���z�NZƓN�-̼�˼�0J��‏��uM%m;�k�DM���};���v��/����QjFwOk+�^HĪ�ev|�u��Q$Qf B���Y#�"����gu�!]uۃ��.�n���X���7n엷m�a�;8��˶۰���v˰�R㫶y�e6��Z���c�y�1���9p���ֽq�s�.�ӮCF�����ۃ�qxC�\��Ӝ�Xݝb������|�i�:y�<�޻7�A\���k\<�3�9�L�7m�Y4m����0���9�`n��z����nA�:݉&�!��Ԝ��8㫣���M���a���ol����$U$�%UY�=5�\ � w'���:��l4�W��8��WMg�D��fjo��Zz���5I[:��?�3N����m���Ĥ�:32Dn�ۖ$u=t�@�NY�闄��<6�e��P���Q��)�d�`@`��a�ޚ+��jw��*�^�  ��M�2u=t�s���J�)@TҧLSW����|�V� ��ˀ S�Ne��_[��;/"���	%��Lė������2���Y ����9q7����Ǜ���ܷ/��#)��	о��d�OFγ��"<CpYG�\2Di��Q�:��۱��βkkq�==d����������JJ��R��\̰#j��� *h�jf6+��8�b���a$����:�2k�B���IUSgP�� #"s#}x�U)����U�b�6�ѥG=�$����xLn���kBt*ĵvރ�{��e��w|V�
��9���V��ZR���B����>�#�?Λ�>�?Q��L��t��rcH甙ry�����;�S��Ԅ��s�YX�:� Em�����y1�~빙`F��M� �ή(�l8)Q1U4!7 ���U��f6d���L�2fg�U��gjp��/^.]=�q; z��7�藓)R�SJ�M�T���5?�Z�t$�sW�~�y2��m� �k�D��j��&vA	�D�wOĲ�	�:�f�ZH�n����Gm��]ͮY��.z��6�ߟ����j�R��OD
��N�pk��&�m��{n;�;�����ю�~6�Ȩ)
��IZ�]�0�#E]�>��ˡz��0�&H�uVv�nO�ϝUG�EG���	!�Ǔ��P��r6��MtD�>�Nﾾs<5mL��U�e���7=ѩ��9o�:;��ׄͽ̡;٘j]�~��m}���K<�)�l�6v�x�c�v>��@A�uRE����7�<c��]�eQ	ܒ,�|���ш�G
e���v���ɒ�!�]R}����ភ��C��~R�Ѽ���zl����M�#���Ş�2�:���v���ӏ�A���;���}}�Sy���~�m�A��{��%�~��O+lg�~���yk�N���\`t�}��o��i��;��Qmð^�Z{5�fNGW�աy��
a���"r���]f�[a�W�l��62D��j���J�N�V�FՒ,��f��^�Zڳ�b�	�6�[Z.f���o��T{5LF�f��B����{�{q������j*���tlQ�:L^<��^���8ac�[���=�1ft��&]ۼ*���37V�^~���!�Rc{^ޫ���87��n�r����!�W�U�^\�����o?B��.Ma�X���g;�v/h>�dxy�0���ݛpz`0�|�!A����W��0>�]���
/×M���� yC�[�����On���-ႤyeXE��8%�x���c�.w�CȚ��V�q�7=�F�L�\�3y`��_�m+�}��	����zu?5�y���g��0@d�����n�j�a�P�<~��x���1dޖ�Á�\�7f{N�з(��$)�Ft��85����^c����/( �jRo�R�Z [�3˽�ga�t`π�R��eN�dPQ-PZ����>j����DH��ڦ��s\��$���`,�P�+�����2�)m��98���/-m*T��X*ɒ��k*�*�V-C2h�j��&fUPx�����%E���*�"(��F��IFE�M�*���YP�]J(�V+P�`��J��6.�Y8�*(�1T��6��)8��J���&������R<������%A�������T9jq1EV)3QU�DF[bJ�a��<�+PW����V,�X#"���u��V�E�++m*d�P�quх��z��z��-h�IQd�(����(���UQ�v��H(1��4(�V���E����j0���,W���VBݬm+mb+���d^5�
�X�`�G���DPYR
�3�V@R���m��U�UE+*�+�QAAx�/q�o<�y�� 2�uh�����_�N���)�-�JM��3�`��w�۪	����H� {3��ˀ#���|A�M{���k��\_�ku��߉"�!�-E. [�6 az��6%CQ�ٓG#ij�몷Up �jl$���������ʏO\�[ch�@6�IPDC)�f�m����]���Ř�����u�ɞ��d����ߟ��(�@"�z��Q��! L��S` W���'�wٔ{������P�!3=�����T!	',U��6;�YL�`�b�d��u� GU�� ���N��;+!�L6�JB�(N�]�p� ����d�	��v�~����� '��[�� ��*���Tii4�J���%�kz��� ���  ���M��_5�2����BC�L�;r��I�8���T%ytLBw�������)�'LD�oa���F��Rv%�݇ ��_���A~
�]�� ���m����wͷ!I	-�qs�^D���:�G�w�z	��̯�^��`@���`��s��Z�����u���{���x�3��,�\rj�/Ʒ8Bt��Φ7W��)�7��,$�A<�|I!���"��D=�u>��s��&N��U3��S��dnWq;pw>M�HGR�Neƺ'#�)E
�ӁQΪn�f�OS�����.` ���`@�ί�I=��V��>i[��5DdR!ER�RI���u��g�]\ ��U�N�ukv�l� ��Ne��s�A1��T�IU*P$���i�+��������N!�3'���Xݚ���\g�侬�I7��K_���&6n7�Bʸ� @>�M���z��ݹ��>��e7 |�c��H٩��Br.��J�Q����l�fI�N�S���׶��iک�������4!.�C���'�RA��H\>�]���9w c��]��7�q)0&��@�d밺��v��,�n�:��.j��zr�\	�:�u�<]�p��Smg.��"l����mϒʾ��uД[�L�pn����{]0�F68�ǌCd��Kp��,.�40�ms�uv,i�68�b��ݳ����v�#Û#�X��]8y#;ƍqxu�l��d��]�^�ˣA��#�.��j�<��0������Od�:9�({fI�n:�G���c�T�f�<��bیu���{�NB�[��)<�'众c�( ��r��Wve{#���`@O:�\i3
��*P��ɰ��z����Yq�wuy����X ٩�	��;Z�z���z� �~@�	F��Z][$�%���K�&K�G��3��Y2���]T���f�Ԑ��B Q�0�Q����]�;˺��^�"�}U7� {۶�e� u,t�;��3����|�h"c���Jr7
I���Y��I/��t������2�dڮʫ ��o&�&d�X�̙�9������ԃ�0	A�9�kS��ۤ�#�GJR-��>6�fq�=5�����S�ʈR�UCmZ� }��_�2}Ա�@m����͎�ʩ��������B������$��U�S��̒�>7��Qp=���F�[�����t��a��{3w|W�I���]C�#;��Od�����9磭��݉ ����+la3��V�&k���֟�S^��|R#�?�&b��]u��l &b�-d���Ϋ~ ٵ��$[9ѐz*��T�CQԯ	��quC7��,-���u7�� �R�M� G:�#ϼ���饤�_v��s��#C��A**I9@��� ��s�g����#;W��d�,t����s�Ez�_f_x�f ��Da�P.5
(�f�����x�d�v7`�����Z�q��n��k|���}��d�UI([}�z���S3<,t�a |�s��u|���7�:WustL�s��~Is��Y�
7��?$��	X�펖-Pݷ��0" r{J�<��|��̚��8�=�yU]�/�!�mA"bHInL��ۮ�	��T����ɧ{霝3KG}�EvC�m�C��&b��<U��8iyM�����L�����6�B�،{}���)q���*��d�oQ����Mޞ_$J�\� ��W>}���p(U�AR��뮡*㽑�"<�| �i� <� � ��֯�ܽ�2׽��鿂��`xgEz
�B�O�*�up� �mku=u�ả��̼�yM���1բfg}նI}��y/��������y��c��3<Uԝ������.{u�$��r�N �,B�S��49�D�#�S�nz�� &x5ՠ����-c�9�\cE78����m6��V�b����$ˉ}��1��L�.�_�E����+� &H�W:���>�h� >IW�g�"�7��[�]ė��jj\*	T*�T6u*�@ �k�ė�s��01��W�I:�ղy$�-�5l:�MZE�JM�GK��h�^�=�Օ�:*�  ���2���n,Ӌ�̭?f��� ��kq��5��y��2��/vb���˸�2�W�}����אz/
~��=�U������~�����:�A��<HC�@�*��Rnu�8t�����luC�����]U� A���D�I}&��_�w�^�(?>��f��Ւ�E������+���/��h�-��[^\�j)v��W|R�P��Qέ'������� K�H�e]5=�c��TDP	�>�����"ą���k2�{�j�6e%�;*fxo-d��K0l�ꊉY0!}��^X"8L�)%��|�]�$���Ā �/�Ȟ�XW� >��խ�3'%�6�^���j@SH�J��:ia���S�>�+�������5-�̿�6k�N＠�����Pn�t�N3n&�N<��^X1$��_b�%�-����y����%=g��$����vNeO�۫�0�%��(�mO�U���8����7�V��XY�;�>^	C���zl�dt�N���Px����ip٭ ���e�t��}�����>)&�M�܆�|�/&�����<j�ػS۹����c��7Xx���v�[����>g�ri3۶���t�ӞЍ����v�Hm�ܜs�[�����uǝ[n��m�ʈ���k�	d�F��hD����CgN�Y�[�9;7�-�Ғ"$\�ծ2�幋�vD�Ųm����r0�X�MW-ڰb坱s΅�Og�.{.
Av�����j��d�ٰqɟU�;7p�Sr�k������˃�;���}����|]<J����:  �[��` q\ө�G�:��W�̊��~��I/�'�6q/b��JPUBi�5̿�'<�{�>��t��� ĳ� F���yKs�J����(ٴ�5O�BSIUˁyw��&H�Yp��+oأ��R��XL��`��2@\_ب�S>`"8L�)%��%��C~�2���ܮ�r� ⱕ3p ��^釫W?Bu�+Ks�:$�����I�SR����f��	��C��'�����݋�� ���"O���V�e�I��]Ǻ��!QB�e-tSv�9���uC�>u�d�Eh���s=�R����ݳJH��)S�m^�D�9������0��K�YWs�[[� ���_�>�o�
AU�7]u���}3�Ee%Q����m��mH��/ڈ+8�"L�w:,���x2�ղ�[�v���,�}��)�N�C�5~���n���8�_bA$C��U�/���Q ;�\[����*9�'������ �D4�t�B+n% g�����ȣ��9Oإ�G��L��Ͼ}p5��h.�c�\�n_���������.2@geu�� ��s\ک�L�E��e=V�L�v#���[���������e�Kb�vLʝl� ��|+� %�VۢO��W�̜��|�ܽ�}�~R~���h�m]���@�v7��[��H���Y���d�@����zi���-]�1 �������9�����Z����PDRH/o��8ɥ�M�[.Υ��`��}��7�P��Ǵ� ��;�sL�v+��\���T{����|�L@��PE"H�p����ڿ@+���%���u��j�'c��U�Xصz36��Qe����yz�X���~���y�m�}7�w�YVy���mq���X5�w�u��K�&O��d��e&\�tlVL��J:�%I����o�� &R�y��� #5_�2����w5L��I8"�UU�Md��	�F��ˊ𨈂z#m"y�su[���s�@Wue�  >���[ 5���$/ǘ���#�jE	$����Z��V[Y����e�Ҽ���qOGY:k?�w��4�m�m��C�U1^�'�]�0� �j��W M�7��y����=ޮn�>=�~���}�DDԤ)����-�@2F�����F����� F.�Kp3�Ϊf�
ٚXd�z��|_�R��yDs:S��4�I�<�Ӂ����Z >��M��^%n��� غ�-�A�s�A�=#(�P�*�I�W]��,�Q�e�޵��FUk�� '�շ���{�O�*e�_��=��s���%U��B0:��{�BJ��f�����F&'���E�h�G�oL�93(a��Y�N\�kw��n�z��R�2*J����5��� �yնx��ś�M�s�@F��Ka2@q�T���_-�Q{�.f���:D��q��A�WI�ܝu�F#z;]���k9u����U;Ӟ�r��7����`pe��,&�t٪�c��i�	�;ܵ�1퍺v�<Jv9��̰ KW�/�"�'X"8L�&LJo����J����2�_m^����+��dD�[4�����
����M�L^�;�Q�I	4R���b�@nW?�L�����n|$_� ���� :�mA�b�J~l8��)5U.vT�s+���Q�6ffx�Z� �#ً��:�z��u^�s����ڸ@�w�ƛ�l(�b]+�1���;�ᔎ򋼛�V7���w�L�w��04PI|���%��:��t�E����L=�Z�h��d�֍�E�ä��`�z�yIr��`>1�����(�| �Ut�y!WJQx��g�)y5ʭ�be�3I]X��ךrb�.��8���q�j�p�/=w}l7�~۫�T||�MgJ?>��{�ޒ��觹�Mssv�>~X#�On)7��N�i�q�%�{=�uDMY`-���{����C�ዮ�F�'���=�/���ț;���������Վ���G/j7�%/_l����i���m���"yY*M.����[��qr�xs������-�g�����ە�E�YCe���r�x蘝BW�`��>�����}��\Z&��P{Ǎ���)nQ{�M�����k�v$������G�N���=��f�E8;���u��!;��6���Ⱥ&8����5h���l/�}��d�5u���k[���3�����e�B���Y�}�����|�TWB�=�f��S��G9�!9 �{Ɲ0�FL�������`	�U�4���
|�����;̷���C�<�����}����z�A���$�cCnc��}�C��\=[��.�`V
�7�ߺ���o�z]�.�^���ڂ]8֯�j�$oM x��w}��rd������W�"���'��W�n2/�{e����?s(��&:�p����b��'}��I�=�U=�q�Mw]ڤ�<d���x�v��OI�t7�gz��r�'r��Hyqt�yc�(��x���a|^H�J�[�Tn��"��{Dd�tQ��\��D�	QV("[jK�aV,��E"���Q��
&�3�yN&TK�FZUI�ʤ�k#Ӟ<�/V�W�*t���X�V�`TQH�J<�yB���DXVd��P̨#\ª"��IR,N���T�΅X���лe5�IPS[]i3U���jJ�rN�38����dW4�!�W�ul�E� d+j������EX�UEX������%Z���T
���J���
,�:b�u��� �8���GZ�X��(�ޯHqxʒ��X�V*0F�b����0�0X�d��21�
ADdV"�d(��E�Q�`V

dڒ��^2��+�V�C���x���(�ZÈ01�6�d�Y��5��
dY�"0Rkb"��mm)S�FT��� �DX����d�VA�j�+%`,��uh,塭��� ��ԬY
ʋ:j���,���2Ѷ*�Ve�kEk ���n���'����4�X��Σ-��x��qS�9��</��cLx�6<۲���FxqW ��K�{e��NË���{v;�Ŭf����܌c��q�������Ҧ���p.�f 9kgq�;VҜ%��܎�\�V�V��{v�n��y�ő8�C�
6�㌷�
u�q���<t�� r®�0�� ��'���]��e�s�l�W�&�nFܾ�<�ݧ�����V=�z��d��B���8�p��p[����k��ng�fN8E��;=�̞�W�����:g�n1�̍�1���0����p�4�8�]���s��v�kc] n�����=9�Bv�vN7�ݗ<�����=
����[�7m����n��<��o)�P�u��
�GFwn�4k�����x3�'��m�����O79k0�6F{�b����p�iM�q���wA/8�U���m��ƻ�����Z�<��`�N�c��KF�!9:.���Y-<']W6��jqɝrZ��۲Wc�(8g���Їcq��cY�ѐ�8%�m�\�R�ȪW^�Vt;]rqq��(R�����hNS�@���H.W	t\n�:̳F:J�\<oS\��v6Ӟd�(���H��X���;5�u�������Btp�qW���W��eNe�z;��Y;=�n�:��������ݗ�+)�.4W��P�����b-�ݭ�-��I�re8.�nk�t�8�[n�5���溺wH���OkA�;u��6��[	�:�׫���د�z�D� v6� �X�qݸz3E��=����v��ב���%vw�9��{1
^�������a��I8�@�Fz#{gݲ���jU�����f����vv�j��*[��ۂ���9yǵ��J�yHn:m\p���a��D��nN�)�{5��t<i��7l�Yꑬv2I�X�N[vu�������)`�Ù�a�!�v��b��ܽ�sc/T�Μ�7�����r�u�̇k�O>�/���7c�1vG�����u�h춃��xwlh9ƺˡ��S���m�e9�pϔ��p{���ۮ��X�^Q��f+=���kmŤ��5�V�h���w.��uj�]C�[�g��b'g����I�GW:j��pM��n�E�r-��[M���r��m�]�����K���`�-٬�^d�9��Z�7G�[
��l�������щR3$�:�w�ᄨ�jz���"P�yխ��V_����]��h0~WW����G>��0��e��⏷���+�k/�Y~R�~�L�ݸ����:��M� �E(�Fɂ�_t� ����"8L�&L)�bp� ��/�s2�r&6�ʾ�W D�٩��@:��M���
"e��H����p�t�nuE�٪����� ���S@ @i�Ol��5칚�y^n�W�+�(%UD�%Ga=RI$�u=�7E͞�	�42�k&Xi����w��>��_s�����ߟ\ik���ˎ�g����n%�����F��$-�����v�n�o���Ǿ�x�9^&}�u�0�í�d� A��U@WCIR:+;{~ރ�)��@a���v�,^��0��L�k�"zs#��8qx�zv�P��͞��MͬY�X�����Y�F��i�=��;�jX�<�6�[oާ4��ޞy�Z$��� ն�̸ 4�*����"*�T_�av��ӫ�I��F�$u�&ST���7d0 '��A |\����K�K~j� G��۫q ��n|��F CL��-�u�ګe&<����L-��&@>6��� '{+n^f罏H~���d�M�9��3j&*��/>+� w�����=V;��u^:l&H5���c�4�Ã�����_��D� Q?ͩӍ��嵷fW\7XoEք�<�\݇��[q���?|� �	���]��^~�I#��,"fd��Z�T�ϧ��]�O�M���� ���i�UH�UP*M�]�7@AsW��.K���}�h�ed2d��j�  �����Hym+��dK�S���ݞ`�o i�{J/w�̨@�:���9��_�T�z=4�W�������-P`æi��{�w)�d9�<oT����`�fmy�:�23٪��/)-�gM�'�٩�#�:6�R"JJj�NX-�/<��ۤe�� h�W�&fN��r�d���i��Kw^���; �*F@!�Jl��:�Cާ@TI얛=�Uy�Y ������������i�W~̸v8�"zd� �D�M��ܷ�i��ݥ��+��ݞ��u����ݞ����#���()��r4I'k5�� ���l.�Y1��s8-^D��u[��z/�)Lʪ�)�r�N@_%Uܕ�¨�[�B�S�"ټ�\���m9��=e���U�#|�8C���	O�Ҝ	w�LĢ 
�ZJz��<|�` �nr��G�.��Ic<P�Sr52��m.K"x�Rt�Q ��l> =�N|H$�GX�YZaR�������Fm]�z���.Ε3 ��xr�NΝ�Y6����3�=�݌��N\+ ���6iw��u-�,�e8y���{��T��-�0ۄ�! �NI�':6�+�w��V�O�����FlӟH5�ެ�P9�1yqi�q�K���v���m��ؘ���ݨny�q��`��}�Ͻ��`��M�o�� �ɧ>$�+W\O����e�l�Q�s�U�|O�lӐO��Ʌ��L��\���NT����?w�0�O�\t�A�_y
��sޜ��Ok��m�-�Ɨ䋀��:�О!>"�:��R��x��qb9�p�F�M) �]q#���a�HCNJ�����ޠx�&�T��A>�Yq �Gvn҈���r�!�y�g_Q�����5BSr53�vVA ���2�g�m��oP�޲O�'�I����{�vhL�/[����oޞtzv�pN��qR�ު������e�m��&��I���2&��z^�J�?����vW�+�����ɿ�;t�`��
�^�E���u����ݪ�k�ܛ��{g��8�C�"x9;n^�eV��ĺ�m�[u���,����<=�=���kf��z�۶ֱ�-��۰�7[��u%ym���@���s�t�G�u$�Mh��s�7Nc\�Wk�;lnc�nm>/6�֦lu�y�� Ʃ3�nu��Y��<��.����u�n�9{Z��)���n�V<�;VX��.���q� \�x�l%�#����������~�N�v��� �J�	:6�"F�f�Tdg���L5g:H��Ppt�$Gr���3��+�=Qs5k�	��$�	kn$Ovf�:�r�6�]�H��ҕ�zO�w�_���`�~S�?�={�^�	�S�����W�}T���n�.@@��7�6��i�ia�-4�	�X����r�Ld=� Qs>@�}��@�:1�˕	�O,���Ďz���(�l(��;��N�����`�����d��gD�nf�H��JL�5�j�{� y�c20L��#m!p��}v�;E�q���ξsl�\<��Nz�����Oߩ$uE��ʎ�Gă[ٴ(OF:^���â�@~��
~����o�"d`�M� �ʿv{��eoO;��vc�=�V�A�aY�e���	ֺv����$����OhSo��Go`�s��ʻZ��v�(��� �{6��x�t-�A��a}wA��Җj�>�0�6Jn��v�UO���A|3.�f���H���8��$��Q�d�@�q>=����>ɰk$L����UOԤ�A뎬����8W;�WU�Q<�Z7��z!:���)>����t�T�ˌ�ۼ�;;���rR�I��P���+��ڄt��`��A��֚6ݸP�T���h0�"��Q��a*�ۼ~%���A�!�����4I¶���I�Z�9U�����}�iHs*�҈@�q�p����?q���su�O�a�zR�Aq�>@�����uؕl�ʭ���K�І�e2Ĩ��$�{cj�I"�;�k�����EP}�[5��5__z�p6��vO^K۲ې����I��w�+�G���OfV�7tN0�8[f�{ ����*o;Ē��RO�=q�)���,�L6JnkǝmC�,mT<�nk.	<_b�H'�����{�6w���em�'Ĩ��$��Q���@�p;�f|I���H�޹��R��A������f�pn��Bq������?��,n؊�Y�n�:U��sv���ɺ�u<`mV����כ��G��Ͽ��	���#��ڠEŶ�+5�X��M�uO�+l�-���H���=B�*��0:��k�` ��g-��Ouf�A�ˬn:��k�̝�m��!%:�bc�|�$���z� �쾼p��E���k3�X��v�jP>��7��0�25����
耰d�X�����I���� �Y/�L��������H�;)M����~��Rnl�G����?LO�׷���ԿH�Ҳ���O<��
���i��WP������U�t�V�L�1��7�Ɇ�M����W���&�C��|f�jTTĀI7��U�I�Y*A���G.���)'��Kq ��o���$�r���h����1��, S	�a2`�w��8�Ɂ6"�;p�B �koz��t,�%��Q�L�¥&�蝁 �]��D�Oq�%�R�P�o�����<o"o|�'Č�ͪ��e!%X�wB�Wʃ�����[f!��H�ƥ�����BH�;
�[���-GL�i�{�TI>�YHH�
V�M"RI0ꌨ��B���uD�y[TA �@'ƶ:����⻻*�>;F��	�,&2Ć��� ���˲���'��o}�cf�����K�}�7�ދRn��!�rQ�|:����/v�]�tR�e ج�u��a��jB�d�\�T�
�z����=t/I玆=�{��W']�L�|��:�� p@��:�.����hk��;�˽�����m�*Fn�[p9'�z��7-��۶M�ی��m�˓��ݭF�^��D�<������ږ��ƴ���	Ӱ���D�Nv\V��xã�^�+ ��H��ی�^&zB��L�Cx�ǁ�Ev#V΋L�!7!s�ݶT�e�z�n�x�����3�u���u���v�-k��q�-�p��)n��R�L�Z�_ÒR(���%���f��YJ|A �V������k'k�:ӿ�&��*D�a)~Sk?�˽j������ٯW��]JA>$��	�{	ٗy�_o�fv�$.��I.0�DBu@l7�H$�S��'ċ��p��UY�$ю���H4w�Y*�i-��	2Ӑy���6�Q�|t�j��|MF��$�flخ��GC3Y�o��'�O�{+E��)$�tF̈́I�sgLٶm2q�z'qH$Oteϐ ��ͪ<O6�a�wl,�T�%8�cg���U��;�uXկ[jL��cT]Қ͔m<�:��P�
(Aʕ�>݊,�}�w�^5�L]�#K1RY�{T&�ؾ� �����ħ!T�M	[�ykn�;�xb�<�1�Vb]�i����L��|�� ����.?$��!�wˤ�!L�n�D�0�2���hr���s�a-l�?-
=�w�l��̸H�wk��I�[q �O��6����t���5������*��HKa);�u�}����\��ccU��-{N�e��HٛP�-�R% I)7���:�n�켹��H1��|�$����(�t�=}w_�&���2{��
N8dq9A|���$:�O�+��%ڛȞާ��WQ �E�f��1ҟo���G�V�=��p+��c�ZԯMcֻ<����8�oDz]ț�$��{>�_"�e��pO|k[��$��l�$�tc� ��|�z/�����X$�~������08�
�nԂ�k{ۚb��fא$��m
�Lb����%��J[�b�Y�r�I8��l�7T>��D�x�$�,Y��m���P�����X)\��qΩ���[�E�ܡ&���Je��7,�5f#�����C�e�Jx����B���D�皨ж{��Y}/z������y�a
�ؼR������EGm�6v��T�[�0w,��t����]х�l���u��8��'v(��H���e�!#���\֓e�x�U7�ޙ>ɝ�TwI�#��/��������1
�[e�)ɻ1I�P׼��]+��t��DY��]U�7�� ͺp�=�2���=6l��v��S�G��<~��p/-���k;<�Ô�<�0����� J���*���K��S�{T���������xg�6�nBz"Ԕ����z)n��:v�~B���$��ɭ�^H\�7�jyx�!T��z��&�3u��{�j��R8߶53�{+){;n7�;���˄�Dh�e��������������Q��ৎT�zݾPl�K�����۾����W�u��Io��ݮ ^^^]�,�C�V|Y"x{r)r�N�"��5g���+D��9-�������,���Ս��u�vRu�n᠆�#��R8sӇ������p�#�=�:Pת��F�˘��>#�7�7��O,vb���g�q睅�LԞ�9]�n!���gr(4R�V���Xe+�ǫcw��x�ۃl��yZ7��<���_�qiDV넀��G�TڱP��C��rq��z=����'�t�5/�"Z%P.y��v�����X�C⸭��TqimP+�XT%b�F�dQb�ʗ��]n���b��H�T�3F*��d��.ےcQE�3�:�Ȳ"��AH�eC$桙:J���b�jZ�P�m8�t�ń�%gNul�"�V9ՖE��(�L9��/)�RfVDdPQ�Z�\0Qf�YĔAb!uԲ/6aDAAm,Xs%AMJ�����P��ڡP�-�d�2����QV�D(��V�IP�g5*���,*�EQ)Zªd�,3�U+9i��Jń�T��QQ�XX��"�6�C-�[aX��o5�J��ȠT+�x˛�f�S%IV��,-lګKe��J�B�E��X�Z�T�.UA�[hTX�E�[T塘�(��Ū�P�.�r�6"��AF!V�Q2�*:�9uKY+�1R��Щ�jFұJ<r)�V�J��]���	ۛTH'�/=��e�RŜ�{O;)����=� �VU
 �N�:S�|H5����DeeżU{(@;�W5�b�[�n	h(�����I$��G\�Av���y�}SDi�JAƶ:�7HM�T_p��S�B��)��6y�ٞ�ӳ��\uu��.����v�n�o������V
zm�O�g^l��:B|I����p��헫z���=��H<qҐO�l�6L&Q	�A�tŜ�]"�v��s�5���N���MtuO�>+l.g)�l����'��AP�
b|��ԂH΍����7Z�tYq;׻�NB�W32��u�%���@�	[�Zݓ�A��ԂA�eD�	ٛ[r��g7�*9umkUuM�1a�mI��;;w}Ä��6��KQ�/N��!����>��z���Gg����GjX�;7��vlӣ���Ԙ�O���f)H(n,����۝B�{j۝��l�b�HQ�ݙ�@ݩ"�7t�g����5+�8�
9.�����7�ݛ�gp���{8� �U3 J���y|�&E4	oG��RH$9��Ovf�!f��Η����	�ݔ@�$)��r4�y�UͰ:l�E�Vw�w�$�F�m)���͡^;9\/
��NT��5��|J���I�3k������	�}�����#E�3��p �[R$�fks<xu�ЊS4��*/����>�@�*-H�w��ڟ/�Ϊ�GB�]��n�!G��a�u�%��U)T	 ���U� �+iI{p�ۻ��:�A �ۙ�D�H�YJA��Ը�P��׆��凳|K:���l�OzX0�}��Z��[<� �".�S�����^x���N��˪��p^����n�^vy�[��d��q���	 �6Ū�Z�>�Ue\:|��r���WdN��`���˶�3��l�QvN ��� 'v���&w���A6ݶ��vp^^�x3Ʈ�t'G[
��(uc;\�m���i����}v;&���v���ɽ�b��E��b�`�2���^Ѳ�����%�պd.M�v�6��C�D�Bp��n�x�Ռ>�ٱu�n���+��W��ޔᘴYW�5������L�p��Eg���~s�&��H(n8�{(����A �в��7�-ݼ��R&P4����ͪ%zs�DJ����3�&�	�c|��#V֓7'cs�#�I���A�YJI&���®�;#6|�����BM�P��ν����HU\�s01��J��CI�۽�$���t�Z<R��I0ꁕ]7)�d�X�&���GB�S�@'ƺ:����LgH�v��hn.)d%�S�%Eu���Fԫ�<�G�UUP�.R&�:�.�ݟ��Y~�"�L)�RE8�����]�\�u]m��:֘�lH���t]�TG5��?�����
f�!��o����+iI$�Ej���=��Y��j�/����[���X���\H��)���l/
�y����z7۾����u��B!d[�	%�t�y��Q�rͨ9U�i�ն�������0_r>�=�@�/��q���ݪv稑eu)$�kc�P ��5�Ù�����:s�"5�,eDD��$���S��$���$�g��i$��Ԥ�kc�|���Jl��	6�0�op�e�9���l�� �|O�jʉ�'{3e�@�0̈ٮ�A�u�|H� 	AJ�~��}�����Ś�2���H#.6�x�fmP���#;����u�o�E[�5\Lс��*�Kpm�@���ڒ�'.�Q��1}��O��f�v\1�V��IgF܄I$wfmP�|t�#ʨ$�|��g�)ԛ�DdII�
�D�)�4�qy�>$V,��ݙ�@�rN����W^8�&�#.!l��A ���]�LGy�[BbL\�Ib�;6)=-�ߠ��G�	��iȪ{�{��]�I���!�W�S�f��؎��<L�n�ˣn����됁'�3j�1oV�dÐ$�������׾7阔�˩��ٝ4	$v'Q3�mȃ��EԄAUÉM��a&�' ��B� �èsƪ���EQ����ȐH'wsj� �v'Q �O��=�K�!��!0�n`�-�_[��;.���B���ξ:3��˱gҚ���������0Ba�q?yH;}�^�|H�N�|x;КW�mHǷ_Ogf�3�q�좢�%8bV���6��Ь��,�P�h$���D�Gbu�A���i_c廐���<�]΅R��	7<���g��D�I�[]w!�U-��r7ē���^�����M�̺�0HdH�ߔ��� �]U��|n���#5:�����:���!��S7��b�i؊��zFk��fS�Tw�rv��?���K�ߧs�p�L�M��Nt����ʰ�<�w/�{9������1���d�1`�U��<��qdo,"�����M�S��I&�:��Ӆ�7�퟿�����=`r۶J�q��3�ڻqI�`�ɻ\������wWE�����Yj�Xr�~� �è�I�]p$7E��OUP$�u_\F�d� 5	�5�Q&�慷F�^Պ���D�I=q�!
�%�[YS�n�}�QZZE��
m�غ�����ې�>�xe�آ�fV�
��t��z�Q"]�R2�	7]��~�)�ҽ*� �H�]p'�{/gw�z��5c�w����iJ
�Æ�}��2�'�o�5{ں�=܎�$�mj���El�m�����,��ߔ���>�V3>�7E���sʁx�7Y�J��n��Ϊ���2<D�s�m��{��=�	vx/"b���f��<'n�O*׿)D��X"Bm��ۣq\��;]n3pl�A_d���\����2��ݹ��mԷ9��k;��3E�Y@�
���/���}v�=��Yv�p]s��m�{ۣ��tl��1n;u�V�^]�;U��\���gq�j��v�[n9ꭲ�Δ��{�/d�Wm�t�x���]�6MV���^n;k��t��ꃳmk����n0�ny�u��������ڗ��	��͂L�lq��b� sJĸ�f����\C�C��0[���OT�E�WO�$6����U,�O\���'p��A$�Ȯ�����hm�m�ڄ�D�g���c'Bk�Hث�|H$m��P$����!��o�w�>��)�l�1;!@5�{T|H1�t��R����MdVJĎ����<f2�H��	����K���@�*+�3��H��{T	#���[�6Ep�ؔ렋ؽ����	8�K.u@�ꪢ�]�� ��c<	�Jځ>'�7�k�{]��OhIf_]��>�
��L�@�h6Kl���iMa1&��M��-��m�#�u<�]_�������M��[S�Iw/��$�k� �<��q�f�v��X5ѓ>@��^m�W�s� �(�H�%�~s�'�����۲.+����}��c�q�ೝ���p:v�[J̤f�n�5g���g�T��|eU�WVv;	Ζ�K�}�ަC���K]3w�:��<�ۏV����ﾩ�H���I>=�����6#�Q]1�>Dk}���i���' �<�I���	 �웇�[� �	���H��2RD���HQ�"���$v��/�a��Q ��LO��+�E��s�%ԉ�>wU�(l\m��l�!���m˲|�����!	��ʯI�t�A���5�4�Ӓ���ʰ��mխ�q']��c6��nC4�^"���0��ۚzy��l�����	
s�:����t����v�$��0�u��a�;^�w钂M��$aA1H���b���=ٯ��m�`�	�����|z�=F��Z�X�o���˦�"	
����[�J;���8`�H���y1�T���_�WL��A��Ky�}��G��}a�-~�a�Rr�wt��ˠ�=��S��p���oO9N[��F6��N�C��7�W��G:R	#�:�i�4D���W�����"n�ͫ�v�}36[�$�	qmĒH��ڈ�	jpaSa�J\nH���(`�]��UfJǴ���kc.��콪�.4��Raƛf�������^�n���YӃ]pt�5�P��m��}??zm[���We1 �w�.|��'�/h>�J�Q�ǀ�����&�:�#�F%dB	�Hh��Gl��fZ�s�#�ޒA�n�����D�����Bl�D�[�I�6����7��Ƕ'e|z��k������v{t	^�\	�#�/j�H�z���mB*��<�5���r�TF��M�_UI �:x#{��S��k��~u�V��Ģ<z:^M�0w$�1b4��A̡���j�,��{[}ڏ�	qx8�N#o�q��:��6o��$L$d.Pz����H�La�黫2�+8̉�}]��@��ӓޜ=��ш��ߢ˛4b�P�`�j6�m��tG6`�G<"K�g���s��>�b�5���J\nH��.�ed}���	���Ϗr[+���x�D�	'�{{U�@��2�d���ۖ/�^Z
9br\�B��I���A �LH�d��]�輽03�W�0�`�ɓ0�ڪ�$v�rI'��M]h�Yh�v-q�'��e�z�c�$M�L68,�Ԁ{btӭ�U�7�\��f�h��o]1>#n:�x;���FTn�Ul�Ux�}Ca�z���� �Ys�i⥝/x,�sκD{�w΅P~yw��	!I��$�	'� $�	'�@�$�	!I�BB@ Ő� '�$ I?���$� IO�$ I?���$��B����$��$ I(B��	!I��IO���$�P$�	'�$ I?�B�� �$�I	O�����)��w:����o�9,����������0��0    � � �        P �      �       p  #@ �%@���V�EP�(
�P U
 i�j�$�EV�)@  T���� +��              @                  ҠR`     @�_m�]jumT�Ԯ3U��3-/]8�7� =�+]uڙIٺ�T��U:����f� ��������'P DP/}
��}sm����km�t�S�� �j)ֻUnv�5tk�i������ �GN���K��Ыn@c��gEDU �A�6kE�       �@��=�GOmA��Eq� ]@ZΫT]`�� �s�F�� ; �Z���+����Q6<}�iH�E|k�w|�{W  �g/�w�^��O6����@� �Z��N@�/N� xP���肒��        ���M�:h� ��>���� , =ހ��t(�`�v�(n�� :{��`�@��� ��z� v�r�-c��`��=��s� ����z��z7Ͼ�����Ŏ�Δ�����P �D;�"��   }  R�.{�[%*�;�Ϲ��kc�����Γk���-|���*[�� ��f�F���3sKm�������U�wu�����]��{X��� {Ҋ����wO|��U��oz�g�B��r��v���$��,���l��O  _}� t����n� ` ��N��hr@�F@�P ��**�         �X����� ��r)$� ��M��XÛ:�)u�v(�:�5F� �v��܆�:9v��@ x�$�=_>�3WN�j�[��֕r�c��
0t�e[��Ur�V�bk�]������f]jU8\�*���     ���RU$       OɄ��J0 ��	��B'�R�5!@      S���EF  L �` L��
y*�4 �     �JLM����������6PmF�<)��>O��~��s���$6�^����>�^�˓7O�	Bu$9���
~A��C��) 萁!h!$&�"��D�@�$�y���?��O����bĄ3! B0�r�В@��!�0��t�P
��B$�Hm!�����X�$b���������	!;�BsF�5p�@��Ώ�m&'����~T���,��E����}�T�j�UZ�����\��(-�A±����zt�����(C�)͸�ޑ���Y��5L�i�܂#�@�3��N�Y��K78��V��Ib�R��)m��{)�Q�^����M��S���8�����r��(��bs�s�|E ���v�g
ԡ�FCΦj�jw��Uu��0fQ��:Q��(��|�:�c+���de}b�k4|�k��Y����s\��wq�;����J����J�ѥ�Y5D0������dؒ���#p�7Dsw�˳�v�:�I�0��ך��|V��A�c�̽u�;��@��v�c}�[�yf��������D��9t�8s��UAݣzP1J
\47MYz#�� ��3DM� �Ý�P�#�,�!׋n�#G1�*P=�rb^{���"Cv*�֋����m�[��ѓ��r�q|��y������>�1ș�Q�t���qF]7^v���(���ɖ�P8�:#%��Ýs 0&q�si�����Ep��h���Y��_ڀ�;&�1��������Qٺ����Ý1f�k��|2�\��ͺ�-�V�C���'�t-ܰ�X�ڶ�C��r��/v8���f��oQ۽��&Ӥ�o�5v2ǃN�
i�I4RY����;E5�<�A�P7S�JH{�K ���g^KQGv��Un��\�@��݈a�-���]�2d���g^Ws��^��INB]%����;όo&������v�w��0e�;	K/�˗��t�vUf5��Q�9�#p���4��/n�f�;#2�.�o&u����.��(� ��:�s�U�1�"��X�:���1��Nҹ ���nh8�^Ǡ�;tl�u^bj3���ۼX�h�.�Z�֞��<.PC",��v�	=sNSrv��s�avqP�n�!���b�E�2��CvkѸ���u�V3��\�q��ט�{�CZ�N3���VR��j�guqUƚ5�}rj��2�9��[Q��7̓��DLsVcΘ�|{���=�՛��.��O3bc9Ӵ*�i}�V������@��V�:VH7š7�e'�p�w7z��Dw7��sq��������+�H4};q�m�`��5"�Xw�5I�Z3p��ւx��vP5�a<��6�87�܏K��OF��1��Q^7;;�Y��ݺ�|�v�ҧO��9-���ʔ]��Z�UZ3X����u����q^�lm7��o�Ft1��H�q� ܕv[�s�^'�>�����o�sj��*Í���=��|�gv�k���y�z��S���� z.����`o7�)�WFc��q�)vFМG'�ۺgF�YȋZst�N��/�q:�=���;�Fu)��vC�fޝX9n)fe���~��̨b��
��8����ųyi�pLK�XwT�0 w7�xvf�'C�E�]�ܚ����k,vޙ�+��0APU̒��3X�7������p�9qu���n�S5�<O�㚀}�|��ݯ����VM<� v=i�ƹ�Y�̝��"�X��/�i	� �w8+T�/i/'������1�s�.<	<���%9t㤼syÜ�C"�	�1i*g`���2NPɆ�� �a���3a��1cĲ�a��峂]�Mg�Z)K"(��{�j�"V�[F�nu�`�L�����_U�Q��g��wZ`?�hX2���1��S���L(E�4&�t��gR��w9�w�ݛ^&0�k�l���b�_ۯ�e8��&�L=^��"�osW�����YÝ��9���ЮQp|��}�.s�Vᜎ',��0�b�9f����.9j܄���经1J�}uS�].t\�V1�s^	��/�'��u��s��77 .����ƣ �(z�c�W��%�1��1**��t,��db�����c�U�&�Ȏe,׶GII�u>�܏��y2VH9.u{mk �1؛�+����u�LAY1ig
xg]��ڹ��Cf1p����ON�������n��)�Dy=$ށ��ƹX�ܧ4,s�ƒ���sX'�7��c����,ѹ��13��g]��˔(.������]�4����U��G>o-p�q�5ۅ��J�����;�Hr���)'�frT�>Ў����<[7�9z�ܰ-��*F�&�U���V�Ap��\��r����������a�h��`g$9^������Wݨת��9s��S��Vj�'�,�px^I��@1�<Zxsg5���Q�\�y9!�i,�oH��`3��r�9wz��3�^���ꎽ3�Ƴv�M=LgC�t=s����l�m�7-���P��oS�7�=�z�K(� Nv���.H��ܣŔt����J���7�p�Ơ�RhX�!��A�Y�F�5���Z�Ww`iqA˄o,뷖5ۂ��}W�s�p���'+�?pm1`�KN8nޏnܻ��;x������0��f� i������Eq��3��f,Ҏܛ�Y�ʳq(�]�=��JǡΖ��rK�#ʄ6��[�p�ޗt7I��.!T�a��n���7{o�i��o�q�C4�NK��t��H0m�N��ǛF凡
_����=�G�5s{<�&U<�j���b�9"���D,%汕��Rv�MM��-�ɛ#ka1D;��v��j�
F{W�h�J5��Gw�f�|�m;ټ�������i��VsN��M�'�o{2�P==z�!�]
mݸ��zP��Ď�7��'C�oj$�[c��.�P�7�@͉�a���g���gr�oru=�Ǻw,ߪ{1�GО��H%0�\g*����y��Cb��L�����u����ͩ�:on���I��`�]�G!/3�#Q�;pĜCu��{���%%� ��K�vR����ǃ�"=�V��P:;z���m�>��ّ[Ǧ����>`)��n)(��Aw���I����2X0Bh6�o�R�%ϗk��7���q��©�p���˯S���5L�#�X�^���$ύ�\��v�qn�W$3��Mol�$@�a�����v$x�t��I����@�!:n�ӛJJ�b崠L�[�^Ō��}�gf�1m�Gc�������N��ud�(y��yI״H ��T49UH���_���p+6|��fhż)�q�Η;�9aص�@����w\�Ha�!�vk�6m���Pr:{����R�������8��:7�{G]L1����Ӕ��8�l�n	U�Jk�M�?&^-H��XY�櫧e��yB	��8�
c�LԸ���������zP(���<Mu���X�􃵾�W
lѻ\�]t	�ۯ�㪃T˛hǅ���--�T���b��nNb{��u$�=�^��[8�=y��H6���'~/<	#�;�ד�9_�\����}:&Gd�ږ�n'�\Ĺ<Xh�of�&H+�\�t�Q�o���p5�5|�E�QF��s���+��p�O��:<��H� �/t�:�Jɱ���G3�p�Uv���fmZ���:�o>:���B��i��[Wn]�9x�5eWt�t�ں�>xK�
�Nt�;�3T3�چ1�g�?�reێ5y`��ۍ˚�[I�vVB��u�
w��װ����yd��uj�q�J`�WL��7�LkD!�7R;z�F�w���s��/��^���5�q�"뼤�\���7�J��BC�|�ц���(�k�r*�n��M�`�ᇊp�y�Y�I�M,wviC��d�-\YX�t�{`	@ڦ\ �4e'I:��u��_�e�B�f��Rb÷Ot��7;����oXn��fS�wb���M��1��������݁���L�69��᭍8��� 8�h�^��Ts��]`d؄�&�^<ꙅ�4eo��h�-h#MdO�N��j�qX�QeK��V�7�Tu�>��G=����po
;18L�����̣h@�B᜺<����kq�3�7����xM���n�]�����8�m��D;�0X%m�O��QK.}�p�ґj؈wu�.]�13ӎ� �L�
�&wC���ܑ�2�x�4�`m��w)ں�;�Ð��=���:�����y�������p��;gMoqe�e����{"��7��ג �������h�G�V0���dA����ik���WI��1�YRӑ��t���{p�u��n����a%�!'��I�Et�w+ݼZWsj�Ѐw�!����Ǽ��fB�
g$�!!�o�6]]�����ŀHᱬ�z`�v."툡V�Ӡ�9EՕ�O��=i�=��!�;aۍf�{��P����~��w{����x��j	a�ï��p3T��0�r<w���W�D��P�cS���"����!p�e���խS{��m�,�t5�ʍ0�{�Vn�Q�8U)�����`=��oh�Wm�g\d�F\�6��_7a�fcs`2�6��b��ă98qF��k�����t���<��Z'�ZPΠ�FH�z&t�">���v̧�����"s�j��j3�$�x�z�F�{={�=t��(����M�9��h�;FQ9c�M�r�e��{��h�ps�:��3���?w>\�:�T�mЈ9�y��-aj��U]��L<��Eڝ���y�]������݁���J��wm�{�����Hd�'I�|���Jp\�&9�wg.��^ODJ}G;�ssP��R�:���i`K1���=R$&�׼�Jn,wq������w�vrӮ>�ꛛ`<VQ��]�/�jr�\ݤ`�c�u*r��L��m�3d������x�b��{Zr.[��*��:�꣎�S�R�����ы�:�ʹ��H���O݄LV�_j�"99 �\{F.��`�4Tٍw\�5m�}%Ig:c(��t�J1�܃Jj�'��kN�)�sGO�Q���ǒGoM��M��8���]���n�a�mڈްt�{�ch�Kxɥ�N����cw�mL��`�9@3��r��"�]'H����;͕՞����l8������1P�\�Hxh����L�ي'��`78�fG�;G@{�X����r�F��L�㤭	*a��'[6��)�.��Q�^$s0�!�(�<E��G��7�I�gk�"�\���Teڑ�/k�NJA)C��Y�R"�Z$�/6G��M�6�1-O��Ӯ�:N#������6���^ʇc�0�zfq�pM5��h.9����&Td��/Ȭ&��%�	�k��cJf�R�)�a��.�4��f�^\�ð�V�}����WrŝK0r�N�i���/��B�{�Sp�ѝwV�|\0s0��� �ۄ�n'�g�.wq���ӏݽ���#�vkw�f��VܸZ�!ss�q:��S�j9z�E.�L��g�_|݊�5���
����p����n�R8�R�{'zͩ�2�ꭶn�b#Own+��Ü��h����ج�w:�����n�b��,ĳl-7�;"{��kq@˛��n��F����썕�\]��6J�����]�w{��d��j��M��u;�P�����C�{�Ǔ{q�ړM!��^& a���+���w�"�����X�h��B�Q��ϓc3w��t����t��8�����r�$��bF����.靑`��a��'y�n�����bA�S!\��̈́��n�Fq����w��с��`	 1i�9��4������孇62��Û�K���ɻ�g��D�s��8]�6^qR��惖L�Qh�t��g.h���c�{�h�2w�^w.n;�RC����<�َc L�7�S�7sV.=s��`CT�����	T�;���ZV$w�vM�+Eɜw*o&�:�ʢ�	܍"�Sl|��8�cs��㛃����s��1�ѷ� ���=���gb�uoZ�����?]���>OݽL��Fb}�|�~XǾ��7l>t���}w�>��xw�C�B R! , RC�$!	R��%`,$� HH	$@ P� )$( ,���	d( ��)$�) P�XAd�� $���  @H� AT�		 
ń��H�+$��$���+!"�H�RHE!$�B�@! �a��+R ��	�$�$�@� �	 $�RJ�d�%a ���
�$�@H�$� *I$X@�	[HI*EE! ���
�B��� �$RB� Y����HV�+)	?��~g�������>3_>�H��B>�3�9�$$��-�@�t��*���$�@���g�ۿS�+:?�/��S7��P-����^���so>�(
#�xS�=�!�����{��%VǇ���9�K�s�c�;�Z*E�ӷ!Ƈ����@�3�w�R���ޗ�ɲxQ�t��/f�;P�Xu��/�p���$>�B=ۥ�h��wO���O7/[=4�wT��ko�gξdJv�hk���5oi�MÚ5��P����xv��W�Oo\U]�ӿu�7qy����t �Z���:u�χt��I0֍3ďzP�x;�;'=K;��븳��u�j;�TD�@t��x#�n��@آ񹰑1\�{^�h�k
�d\xY3���W4y-~�dLJ�y�ۗ�p�wt�݆y+9�r�뫇'$J-�5W��I�o6�� m���>���g��Bs A�7wZ���40����^��s���Rk�L�_�_�9�d�G�u6-h�����f��H������Lz�� �IݨrŎW���roG6�G�$�Pׅ��2�ݼ�����Vݭ��d,�|��V�f6.�^�����vjŸ�����wNi�Y�K��(�3ޫyof-C�e;��0;y.pN����x��H@���<���EӬ<�Ds[��u�k����N���e+�"s�����%J�Ba;L�xbk5�[fl{��k�=짯5�y}#�4*��mYgϡ(�VQВ��#[jhw�Ny�K���M���i��f<����t�g�{��+yf�s�
�&v��#�n1us�;A�{-���pD�3J�Jnܽ	����hPpl��ov�{��ԝ����+ժ/z�/}xQ6h�T�aj�%�f�����k��6<@�V��� �L�Ϗ��	7G�|�Xg�C������yZ��Aٝ��GwyJ��t$���2[Q�UA���ZdD��(j�kC�o{8N�^����U�軬�y�#4#r �bꕷ��maW��$���^&n��:�h���N��h~�&��ґ��@C���u�P���y�ry&MɾZ�|g�A��Ǿ�ԫee���Et���/t�_%�>~��_�� =�}��;{C0r���q_{��7��,��]��:�}T�?5����P������!{a�Rcj�M�����O=�Ļر�a�r5���Ws��FRk�.��Z��34[�����9�7~>����W��$��`Z�4n{ɯpk}}���ʭN��x�^v�z�����2�2��"3bv�Vn�����[���*�/d[�5��S�W'���he��9��~���p4�Fg	�7���1{sm��z�Rb���؍��v�*i+��襟i�ͨ�|�u��S���iɽ;֧f/�� ��{B�@���}^t�OZ�m�O|�=��|��{��}�Q~������Ybn9�jw]EG.꜂��KX��ns�<}���.�Ic>�w�4O��(�Π"yyX���+1r���w��Cȸyb�|�o� F*ɏ�;�Kجz���Ӳ��ǥo�]���M��j�rg^y��ү�EM��g�^SS���N�*eTlձ' n�P���^�{x���c~T�mk�9�,�(�D��p��ՆO`�z�4���Nj� 55u���\9e\�-K1��{`����tD�����ZM�޹���o}wڋ�Aj��Z��M:�{%�^�t������S�1�G�k�ώy=c�S{u��TA�կ7\���{���\1��ъtmtgk0��=�g���/7U��z�s�p}�-��v���������t��/n���s�sJ��d�����f��J��|_�d�|qÉׇ^�$���{���h��m�{;��x�`NnpCP����u�����s��C��4���Glһ���{�_H�g��x���=O��@�`aqFYt�(Q��3,ԧ@��)^�xz���\������ Trx�E;�}����Ǘܶ?e���y��������]8����u��7�w��}����
0�t��cp⚘��w�9�|v�7;7���7ü���K��:j�V9�w�g�cB-D�l�F�3H�Qx���P��*|��n�wf��Szy�=�t���1�=a]O�]'����铋�j����dId�p�� �<'�E<�����ו�����5�G�������}�|x�8�Ľ4���l�O�^��X�x�[��3���w����>�*<�x�Źs���t*{������)�ٹi��9��Ӻ����w�NA�>��'�w7@�x�+U�E`��7�:�3tB��g&�8$!��5>	���u�]�i���/����G:-�Ofx���\���No��:p���������h�l�ͻ��Q�0`��+���� ���ǣ�(�M��sz���׷8�>�`�v]��y^\�GfRNKk͖w�.ha
�9�O��o-�y=���m��B_.!��W���}i��:��L;�x��*Z}����s�-\�ǰk�6�X���+f���Ѳ��0.sP��{v��Q��sy��Ub�/tb��.��J�w%ؗ��.{s��[�91E3������6�0a\��^91!�y�:�_�b�S�O��
B���f�����X&���ϸ�_i�{����|S��2_�b��B������鷧��.����mgM���1(�J��`��QumHQdQQ�W��'�۠�G'�^�d���(�[�KW�)�̶��Y��t9�; ���U�_u�3�/ySs�>���]r�nJO�����+G+����q���Gc������瑢���e]�`֒@�~���Fs��c��u�{�!�.0�ά3S^]�j����o�m|�^�Ծʋ�+�8��wf>�+�)�䒓�l�5'|��׍�؈MM�Fгb^�	S�P�L^�"�YY�7jz��/
̋�\�Ѝ��U��s�ǫ�àԸ�aC�`S��M��vh��R;-�8ʙP���ܝ�?a�{9T�������ݧy��ѐ�]d���Q�8��฻�{6��>@�3{��`S�g��g>�i^���������L�� d^;�@9��wF=��k��f��eb�Y�6�^w�3��5
<z�<�>����:0��^��K�߲�����z���y��f�>D���^��}@�I�|嬋�#�N I���y�7np���~�]?m���E�$%�.00�9�8�u��z���������n��NLCC���C����w���I]H�ـ�"��	T��A`��wG<jce^ݎv�v��'��^(3�=��m�s��s�FnE|�P���.z�r���X�<F̛�(�A��w�Fny.Y�n��'��o�qLys�퇕%Yԁ��3*4�KP7bn30�gZ�z*�X6o:��O��� �<��_�8�פ������g���a���=]�=�kFZOBvtW�;��̆t�s���^���r0��UA����k����-�������,�����V�W��r�w8�i�������p<���;|�v��{�1=���X�HCy"ʣ��J���\^ߊ��N�ͅ;�/�y��I�.Y���bR�r�w��I�ǫ�`#P�Uߗw6�J����i>�6u��0f�	����y��dz��N!�\����V��ٵ�D�r��Og"1����q��׆#�Y���v�Σ���Ǯ/ Շ/��Of�i�*^�-���o����ޭyz':�=V�yȖ<�Up�o�@��Ut�- ��G�tE'���k��Q���}�������^�Y�o�W]�C�W�Y	6������d�S6����m�x��4����9r�	b�qhzQ����d�y��b���/��M���H����ۑLb7k���6��a�W�gڭ�*�Qv�7}��j���sN��Gk�$��Q0�G��K�ܷrC�%�_d�\�L򷴍��2��U���p��Xq�x]=�u-�����>�kl̽C!�Xݼ��s�#I�ѻ�grv�1z��Cp,��v�2d�m�NY��av��7j���n�(��_S�/w{r�k��&�(We�JjPv��I*�fߌkk�qbs�t��$D�Z��^Y��24���;"�CYb��eF({�Ү��v�.A�C���"=j�xw���e�mx�;�w74�%N�=Մa�V�ћn�����D��1[��0-9��h�5�%��̺�l۳�H��yxm�{Ø����ܻ���ڛ��=c�ѣ�)�a��]Th���r)3�[���I[|�sP��U���:�+W�����X���,�t����̉�=��>6�h�t����jPju�������TL8�^2�D�̮N��{L� ���KS���jw��>5�e��%�܍IŮ��Өn�'ԧ�	x��M�cV�b��MRΤx��C�YCU5��^�s�r�t��\�s�������k��2�'b�BqZ��,���wb	��hp�z�ԩ�LT�}�����V��+D���մ�c��g5�`J�{*~^�ְ�0�X6�!�(�*�&����v�v��{���o>��"{G���ݭ��ĉ�[ݮ���WD�=�Q�L欧�R�yP5���Ǣ��Gw?5e}tvl5��b��F���&is�s�ü�ѐ��:V��O^W]�Cszf�{i��n����ő�1g�Nӏ�ŞQU������ݣ
����g�����ҽ� .�^E�t۫�Z��:�,׉Ԣ�\�K����z2�l�e�{x�=��/��vy���8�V����=g3hc�1	�B�a��?9
{���J�CyGU6�i��ߍ�X��iZ�1�g��>�n���/<o�w<cs�&3�x��e�����~��5��b'6�r��D�B��3�*����`5_o�'��@ǺX���bl8(=�ݵ]�h/���p�[�!�ކ��AGג�%<M[�0��OwN��ez^>��¡Leq�]'�3G'�D��ȝ�;v��]_1�<8���[vg_���I݀����C���������r{�W���9Spш�8�Y3O����������ޣ�{6l8й���ٚ(Y#��k�pÇͷ�{�����dM)^k��S7�m�_�L�7g�	��-���i�{�j��M���L�u�|6�.�/Bb���;��A�>KQ���O�ɂK�����yN2Y:^}ď|�=�,��˶el��N��؋������
3s�,��Mꣲ2P<_��B.ܬ��!E��9Ea�($Jl��?����VҒ��ܴrc�!���;��o/h=�y�yPU�b�HN��j�`kH8RF�b
E�
u�L�.�b���|�{�=����0�9�UF��B^(�v�%��v$V�-�7"�O����	����|���F+�4�Eȸ�3o�j6�w��d=���w����ǽ��&�n>�s`3���ؑ�A��wr�3���D�Q4�nέ��pol	٠��q���g���8�������C�ٰ͎�|'m\��ATL��#��92q�^��!3�#c1��k��V��̹�f�{�=�﷈ul���̑i)�+c(�2D���Bw#0�͝1I-#Z��c�㻍�3K+�3�-���\sp��y{`N��I{�\�OzL�=�����y]��o��XGS�j7�qj5��%T�nM�%{*oF볹�)z��w=Aa����5�2<�z��ft�bu�g?x�X&�EX.�=�Ox����Zx)����������ox�{s��պ��]6���;M>�+�|4M�S�Ż�x��<�7�`)¼�o0|bTܒh�}�a$�82D�Ӻ�E���Tb�q�&��_]��񾹷<;��n�����I�z3|6�f�Ep�$xg���|Vo�kB��e���z���|.��Q�wc͐����7��F�+:r`1&f�C�.Df�{����(�`���
���-�}��4|־bg�����Xj3=��]2�!���0�'�h�������=�Zw�m>9sc.��y{ǲˢ?*+��#r�l�61�ؽ'FkX����#$�0{O����r=��߰x�t�4	
.����w|�6���.��}�;�i9sL:<޴�j��-�=�[�z}�Oggc:E����r�3���dx��yN�5��MW�6�����ϑ.n�K��;ݮX{Y��'vT�-����OpB��I�d�`<���&Bм�(W�u�F)9���n�:�Z������>��.�kns�Z�'�B@$�A"��I4�h ���9��ʃUr�k�y���ѵv,S��3З\�n��]n��0��ik/l�k��%��醼�'oC�u��y�;��YgZ�Иq{�%k��ɚ�z��N��q�˲�Z���.��vw7����n�M��v�ܜ=*��O]qna���ֺ$������^�=k�֋�����O��`�ݐ1:+����k=�����mH=����l4�d�nZ��^�¶,j�3��`��v�E�'g�y��!q�GiӎM��^��T#9	���m��l8U]�q=��6뚝��b�μ��xv9�4��v��qb��.�ЊF��M�*���1���������FG����צ����˶�r��1�ݦ6�^�a��^#gۣ7r�#�'s��>���a���hd�n}�n-���!��mۮ��ܝq�m(���rp��vс�y�J�'dE;c��Wt�����'/ku�]�x����ӂ*7mBNq�/��}��s˫�^܁��[��P�9�=f��8�Ԅ����<��9��l�Af���u�wN�6D�_j61�X�[�Oc��$�+J�'�� qz�9�r	<.�ؽY��������5s;=m͵:���s���LvE���6���И��V݃��Î�a�=k���O[f��=a�:�*�ek��촺�mq�i-�-�u������e��.ޏa��]{,��]<��M�Lӎwx���Hu���������m�����Y�����h��r=��wzn��9lv%2vۏ;�[��x6����&I�9���6Mr�k�RZt��u\.N]t78�tuk��:��V�x��[k�<����N[���M�1�9��Cu�ղm�F8�b7����-�8�n�>ݻ��8lS���r������n����[!˗/I�=s����,��q�q�9ۨ�f(�FN�5y�N�tvێd�F1���S�R���wN펅�������y_U�sGkv�u�jݶv�Ś�����<�a�Y���^�a��b�A��jV���)pn���u�[�������y�s֧t�q�n3�j���]YG�=�6��8���p��j���]��nͻs��Z�<kE-�]������=rp]�u�3��;jΗF݉-�e�z;���.�Qqɺ��nu�Խ�5�KRY��۱C���k� �/Qh�#g��n���y�]F�ƩH0��Q�B���N��;������������=�'���kN�h׳� K<=����e�V:^�����<n���ՁSb;=�l-�p�{'"s� p�k��������l`�z� 3n��l�:7%���Hn4F��0��.��wh�(s���y룬H����㓞��r�3g����]�����)�]D��z����KuÙ�t���E��6����=��[�����a㰀�I�����X#\nڮ1uˍIӴ�&\<���ݐ���e�Gq]�g>.�m���69k��lY��d%�v��u�0J�Ep��7s����c�U靷b��f�Y�KۓIHl���u�7@��$���0V��kn�1ٶ�#�6�&ڌ�k��7���I�F�j"N�on����u�a@�\���]��^4[�soo/m�+h�]��bSh'��mz�ոB�nGvr�N+����a�@�k@ᮮ�E�%ў( �k���w#ϲ.�n$�9��W.�)�6��d�A睺�3u�/��.������y3�w�i���f5j��7>'�֭h�9�.�궸:�5�s���d�7,�p�ln��n�nɍ�y�P�tezjzmp=������`��֭������Bjx�n�[/�m��b���Y�`�觝rf���A���F�y���v�G[̀�[z��b�Ս&����α��=���u�d�5"�v�]e�T[���C���8���>d��|*����Pt�{m��������<�V��Wb��f^N�Y{qf���.1D�@kP�M�5����=w^���ӇE��\F�wh;�u/=����Oj�$8��l����1�z��[8rp�K����W5���s�`0	垭r�<�Y��nB�)z��緰�66�����umV�K�i�ˉyS��]ێ6�š5�{v��6M����k^����#�촫��B��9���0�iju�yKn�q�7/;S�r�|��أ�B��G��k��fTwr뱨�ݷ��<Ƥ���$�nլ�m��{b=�U]�]vܠv6�����g\r�'�(r��r笸8w*����j�l�z�ڋ7���X��rw`�ݫ�=m㵶�Ìa^1��s���mƗ�:ь�z=�8�ݜxڬX�۲u�Rs�c7�{VM�yQ�&G�o`�.8��\�f�ܜ���ŽoW<�l��U��@�ڳ�1�;s�9��nj��h:7OX�/��u��c���n�F�ۏ;�(��o6�M<��lXR3��G�ە��װ.��69�f9zzz�ȓ��Zq��pƱ����f��)�c<t�sG�GWe�sR����y{3X�r砧o[t����I��Ӹ-�۷88����Aݻ���!�;i:���t��Gu<��
�g�s��-7�䫋%ݹ:�c���>0ٽ��p�qz����պ�N���Pݘϸ���1ٹ�8��e�[�F��h�j'9��]eHu[��x�]>��v�`;[e�ܸb��6����Ar�q�oWU2l�K^����/9Ǵn5j�{X[n�:a�q�&��@����ǋ�=�-n����L�k=v�N�e�\v��v��n:�,���WIkz<�E퍉|p��p힇����'\l���앹�it�]n7iB�:�pnx��΍Dj�����[9�:�FK��^�LM��n�v��=1/jB�'C�q�tKq��ŜFϳ�&WH!�ۓ�[�KH�;qr=�l��n�
b,e����h�hLc8���霛�N2-��]M�^�ks<�h�ձ���|�n�{n��ۛ�OJX�9�ٸ�nx�v�;�(�Hn{=n��%Λ�ɮv�dθ1ώ��r�f���&'z�$u�Q���n�]]]��.�8:���Ɲ<.��=�n۳��h�u��)u�c���(²�-/;��q�ִ�d�8��)��˳�����u������qs�8޶.;v2�����!ݶV�������c]��J�1]+�]t�OloI��n"6u�L�]�W�\6��b�m݌<{�;��v�ε�L\�I3\�cֵ�^�A��T{k%#��F��K'\v��%�&]�nh|�V����\����YݒW�ʜZm�Y�91q�8�ݜݮ���r޻lu�np�n˂N�� x�l��}S�c��EA8:�H�8�ء�y�p�c��փ��HU&�<=n`�^���ԫ�N���\E�h�)���x:ދ\��us�����{v{rl#6�������O\;[�����]���'&v	S��ܺq�e�����C�Zvmǚ��z������}m	�iwe^���0��Sl;��Oj]:͞y�wc&[���ʥ�=Q1��˙^ŋ0^ܾX�Qwnَ�Ȏ�9ٵV8�B�u[��\�(�mj�kn\�ɧ;r�m9��+3��m�͖);�n+s�4��8.{')���q���kɞ��w��8�]lq�(zڼ�p��v6��u�������(��&5��
���G�M�v��{z[n�U�p`��f2]3�y����v�ݮ�v�g�+�ۮ��ˠ�N��
v�NM�1v�����9�:�v�֝΅e�{:�i.Ł֣r�^�5�u+��ۣ	����G����s�ɞst���J��#������ʍc�:(*D!�(�s��Q� ������w0��mj�[Έ"�D��]��f�Ϊ��,�O�^���=�h-�nX|7L�mt V]�ź(tu�s�݌5�V.*�6m��\f�����I�6W�&m�Шۗۃ�Ta�궕��yI1���ˤtn��Y�1��r�9Ɗ�T#��������O���o��G6�(��t���G]�,\�ۤCO\�<[0�R����V�6v(3=��m;��t�ۮc�z���Zٽ��\�Rjܘ�����Ǜ%:0(���Ky�&�R-U5N�Zj��,��$�UJ�UU6gf���њ��gj�B%���هRÙ,]u�-vô�:�Is��C�"xS����NlEy���n�ĳ�71���l�>�s{�`ꎹ�����t��H���۳���l���I<��"PP���p/d�A�p�*�*`7�����t�7���f�ɉ륱��0'EHt�;���z��/BfΈۢ��{d5��ɻVf�P�n;qn�/P�F1����)]8�;O\���Պ�=���76^:�X�;�Y-���ۮ��tm�`�;N�{f�^ݴ��[s��o:y�D�1]Iec�#�ְöxv���)A�	�g��o����q�ǸG�g�ÄqlQU%U�+DB(�Җ��cTJQ��DciFE"�"���E��Z�#�a����*�@��[e�Q�J�c��Z��2Хp�bF"%���ZʚH"fYcJ��#L�-�ȑ���ȒB�Q�ZE��[u"Ҋ��w*R5��ݪ��
�R�Z$������AK�(� �ҍ(� �.䔤U���A�-�V�%"%Z�V���\���hPX�,DUF�jK�JV��T���AV/Ib�J��iX���m�����X+P�Xa��
 5*ł�ڊa�a�,m*ԕ��T+#1J5V�
Z��.�%����r�J�L\c�Eb��Ʋ���AC	*���b0�k&*(�E��6�,-�[vL�j#�#@�q:QU\�?��w���!f.2I�]gE�N�o<<�s�lFű�5��a��H���]w�����,�\C�;2J�Y� �}nN�Wꍲ�S�˭��ղF�n�X�\�<������d�DǮF�u��6��̙����1�=�x�,��͗��\���u��S'[#����e����#����/�jv9��^0u���&ϖ�2lHp�B8��e��z�A�rk=�3�ݰ�.���j��p�c�-�j������^�N�q�n��mZ��c�W�L����]�^u��9Lc=�sv�P��
ȝF\��eD��&���N��.q���d�=9�c�ʝusq�׵��}�]��o;u|����	��h���sl�t�Gj��퍼R��puv�P�!m�2�;m��O9������n�5��yu�o*��'v¨�*�x�^[���n	�8c������\vul�z��g�G��d��Kg��tG`��_�N�w��Vz�Z�۲n�<��
r]m.vL��5�u��H��4��R��v{f�8gY�.=��m���G:/<����W'���@=�	����3�`���p�f-�{R�1�-Bu�f��7�:�볧���.��,i����Mٗ��	b��,g�n��8rvv���㎑U��^�T��˸磎�nC)���+�o9V�g��4N��=���iŢn��q��v��ڏ.��.�����]v��˷N��q�v�<�ˠx�l��<��\��R�՝2�ٓ����t�a�Ŏ���M�V�J9�s��^�E�9�p!'00GM�;s�&����|��t�(��ܺce���G8�Pn��nݓ���2�S��)Sm.��=�:6��݋i�;����z�Y�������	��yv�n�qɑ�ySa9܏lq�x�y��7��y8���
`y� ��Z�F2���Z7,Q��۱�����G/�Twl�v��Ǳ������=��˹�6���9U�g�s���ϰv\���{)�|���ܮ T3�˷.㟔uĜnN\�<;�eɢ��G�c H��~���O�R2��5lĿ��������v�Q y�(xe�i�.���}��p��_�d��쩈�����-��A�h�ޅ�v�����ǖ�^	!Y<j�A$]uI5����4����zA�?P�@ܚ�&�H/�� y��rb{=;��|�	��$�@�u$�D�pf)'����܁�gM+������I$�6�$�H멤�H-����k�k/;���m��r���gX��r�F����U
I$���v�{y�vL\q�	$�=�SI����$Z�ʇt���Y�ò0��\mP�7	#TR��f+Sa�5vN�{udR��quGK(C~�� �v�ɠ�+;{n�%VUm�(�5ҹgo�,�~����}���H�K�E�o���	}uߗH?t�I��~}xR<�m�dSY�z����r7zⶮ;��a�yil~��<���?��⽛��Y؜�u�oj/�Hι�	$����i�Ǭ���30y���7��@*ҵ#��m�� ߽��{ ���y܋�Yp�Gc��$�Iywweش��dF��u;d&�Aܛ���~���ڀ�B��
H������$�9Qĺ�� 8�ɑ�$��e��O۔R:��9�)׻w�D���uU�'�ӳ���6�I%���v��G*8�Y��k�휄��m��81��nG,��$b�0Wu��sGn�q�m��{r5-D�}��)�\��Q�]�, �{�ݤ^Izrx�y!�=E�Rb�G-�|�����G5�U�eA0�8�TN�Dy�;yvpNL�I$���˻	g#�z�&z"k��fV��Ђ���#-*��n���{{��6�� ���!-1�;b�];0�5���*+� /���Ƨ�s��7/{�%�O�z���G
_��<6/]��m.Ɉ)v��rW���Ů��&I$�^�Z�0����<v����=�gw3��7��A�w�֞� }}|�  �S	���.�#SݮŤh��bT[!5��0�^�c�����qrN�-If>��I#=d�I�SI:�]vN�S��߼i�5cO�e��A�s�V����݈�]�Shd�፤.����̅ۃyM낞�ۻI"kc�Q+�$z�M%�[[��9�>�3;υ��Ak�5IDb��?-	-9�C��43���2~ݛm���؃��w ���. U�qo���|d��u��#���Jڶ�����w� \��`| ]{|�չ�嫫�t>=�ט6���.��/
FKc+Ve�7�qs��+�[o��D��ކd�	/��$�Y��nX��j;taA�<�gt��#o
i��}��+���w��z�[�w#�.s��O>�l3���ǽ�"N���L�9�Q�Ԗh�[��F |�����:v� �dz���
I$��n;�T�jk���]�Ʃ$^7�SI$��n�[=WK��L[KF���R�e�	_��kn[O�-P������Q�b����gyQ�*���q8���d&��;�xcb{�A���~�i=���f���{X������ޕ?nQH�r�����w`���^��n��f�a� �����v�]�+�^ƞ�q��T��9qB���[�YUH��n�;��I#��k����Ix�����=������QJ�v�C4��My뗋�4鹡I$�����$�Gq����.�v���\�O�%��[q���׷�I ���
��+rK5�SI/$������A$���r�-��;.G8T�T�s�}�Y;'�4���4%3�xn��`z/+v{�b�/M{u�}�e;�osfb?�F7�Y�c��!x��;�^��׍<xFK�v��=��ݭvxy ������SC�'��^�M��n:�м�����ίnp|�̅��9�1��e��t��ge���w74�p�wZ�2Zp�z 鄩18]��5��s�s���c�M=n�1�zĳ]/n���9�7H��j��U�=j��O+�6(���(l;
�<�7����/k��wGk�x�G>t��������#��!^eU%�J�w$ߒC�H_"�;dbO.(����H�wc�iy��`--ӱ�'�hO	��cK_�y��$���˻	q��"�J3��;b�+�ɤ�F՘3`�1>0�o={h�u���H:�P%l���햑)]�����׊Æئ}c�ȣ͋�����7�f������O` ��L� 	��L�װ�um0�Uw�l���#��$C���a�d��s��܊8m����[p�I�ퟋd G�Zd���l}8,�=��] Gc�֝�*m�Vq�s�F�b�]q9��:�:�*ܮ��=�+d��n��g5�mO'�"�A%��u4�{V��8<��݌ ��L�K��s��tv��F�{�� o���[\}^���kӿ�o �i�n��Kv6�d��b3V�d�׋N�n���z^}� �+;��]7֐I �'�i$w3A"vNc��k����f�{$�0ɑ
faC��7�L �n��c|�/�ٮ��� �k�}���\@zwf���*Q>0ڞ�ۃ����z�&<��M=�������ﹹ3�����ۤ��Ob���-�G���� �{�ծ��U��!�N/�RH$����H$��v]�QS�[���Nђj@*O��'T�kR�g��Z���C��**��7UUs^�^�֪�Ws��L�����6 3�r읹ق�peu.�"�@�]M$����(�t��T��m�@C��j�u�8��E$�Ix۩&�9���֊�SS�e�f�}�� ���=�S�RI���qݤI,�=�q/z�
p��H3."�����TomI���_6��r��g
۟���r���{��'7�)^;:�ɤ�����X\e����H�[O�@���^��?h��4�[��&�t^E:�.�=&BA�Mz�H���.��K#��5�"R�8鷒I~w*k�%齚�ڜ���4�3��V�=�SfE<]uj3�� c2��I$f�]��$9=�	�����s��GF��ӳ�p�[=mdi麢n0Gc>:4�~���є�Ŏ�(���w+m���޻� �<�s\�޼zfԓA$�ܻ��1���R�5���+}�]�;1{g��Ƌܝ�H����v$�檑A.y���eSxo��}{��+,u�.��so=i$���t"�H���(��"2v��I$^�[$�Y�RC���+
(�0Ë��4m�勤@{�\�͛	$�kSA$���D圥[}Sb�`��X�m��t�SC�zK�%T��3b�ؑd�Ν3�;��Z��S^�fD1����ZH.�޻��p0K���ə�� ����aşj��:I��Ov�M�ykU�D���u4���O���
�����X*����:d���m�oWMc�8���A_�"����=��9Q/�w����l�{X�  ^��ϐN�����Z(�w�E$�ƵT��+(C�1*-�:��RIE���v:��{�э���\@ ��;��w��zn{��~Ϸ��R�3�0�K���ws t�cb}���]@ �l�����^��q��K��ڟ�;�({N�v�@�B� z�H�gc�����y%呖�R^��+�����ex� 7������{��%�mQ4@���Iy$nv[<�jo���4�2u�2��VZ�!b�qYt@M��^���������rg�ꡃ����o0��ϙ��󅝾���|s��������ypc�}deo3�'��x��x��IN�PR*�V�2���{v^;�s�I�u̐"��{72*��q�.�[7+�؎�J���l�A�w57AuK��yM`��]�v�pr��v��'tN�[�{Rc:� crlGQ�����pi�3ќ��P�Kg,�g�,��i{sqsU�е�꫏,D,v�PR�6�z�p������ɛ:U�ά�5�S���ψ5q��}}p������x6oY1����  ��{���Е�"oz�]��tq<��^H^���ޛ/�2HQ>0�
{on�$���u*�b�H�rI$����֊Jӎ���u[;�f�1j�X�"���'�{��$��'�A�&��a"Gf�o> �y�okc�}��AE X��ږ��WY��dm��H^lש�^��˴�I=��?����F�dp {m�IWw�,k(��z����{ t���&lbpH��M$I���b�%ydu�Km7.�{���C:�+n�2��b���<\S�cx���qq�^6�Kh�ڝ���u82��4��/6�8H߽�� ;R���W�Gd̴�	$�7.Ť�	r�*&Rt��mM����;n��Xt:�y�k]�ˍK����ܚ���b���Un�D)��.��O��l৉�.�����ڧ�XK�{L.���)-��o-��o��7���혖H6�ڶ�<��O&�"bI�
'��ׯF� ���� �i��~��7��jv� ���ol`'�W�p��	L0o�ueRۼ��͍ʤ�]�1�� �ᘀ@|��������76.�<�kz��Ϲ�ke��a�d��s�����I�-�'3z,�s�.�����RM �빚I��S�'����ӚP�j+�u2��j�YZ��5�#,%R`INq��\bR�V�{��`�v�
K���k�ލ�N��)y$G��i'��y���49y���7�� ���^��:�F��	����Iu��q�Q���cg<���3 ����s�9����۬��f�S�EE��`j��Y���$;.hRA$����������\����fT�ͱ~�{iV�y�f����� ]'Ba��N��B@;�f���;�&$���{m����T6A��b���I�s�(�Q�~قj��H�h�/��;h[w�r>���{6 ��3A�ߣ��z�|����ׅW���������#&��%($P��/qS|ʘ�x."�{���MWea�s�в�~��t����L�;Z�]ئ�4�T�]]�߇��C�6�7�����Mj�	11�_Q���s}�wwX�:�Ƒxe�Oxu��9�������X�J�N^�y������e�{8[4�3� &����W��9�����Xs�7�u�Ƽ�; ҽ�:s��I����L���z$ə��G�}%����Wh+{s7�xȜ�>̈2S��ؘ̺��qqU���F�,o�f�W��/U��Dy{���P����0�<��|�?y�-��S����OҾ��Wox�{6��F{VyToM���T�@���`�O�&vk�/�`9��,dx�HƳT$�x�Ҹ��iZ�.�٘P�s��׹���D=�R��]G�aS�K�-$O�|/�����P�U;��参ս��>g{�j�ޞ�v�>��5����Q�o��w_w�n1�����=�`5��i�[�F+�f��zT"�-�H
���C"έE޻��E|?�t�:>>��xؗ���%�ԀȌ�E$���*C �6�LYE�،acQnU�,���l��ԒR�lTj��F�#Vڗ*��[.KV��*$#QhUU%I!r*2A�%�#,�I ��%ԻL0��n-ŶڥQ��@m�������(���J���0�H�T�մ�(*-�c	m,V6�G���#K�h�BD,d�G%�	#Bȅ˵D�����#H���S;�����W�q�lnw(��Z���[URR�B	��F����V�IA�5Z�l
��b(�2�Z����n챤XF�V��`�lDrF�,�K�H��$b�2F����F���q�#�l���5��R1V�-ȅ�b5$�&�Ȓ�HA��mM]˻�v��QTY
�DA������4;	�dr�Mi.iI�V����w�ig�=m��c嫷�<91�{����û�8��6�n�� �cCh@P�
���"ԓW���FFIm�8�P�|}�;�&;��B�A�@��pLm�0"��7�έ�^I�>�T��H��I��6_��1!D��aNu��,w��G:��0�ɀ ��۟~�$?s߻�����#���_�^b�h
��wa��4^K�߱ص3N�D�fU`@�5�3�/wv�� ������d��޶�n(����⺟Ѹ䃔b�6�ai��5�\��X��`S�VE*�w�yZ0�R��0�K��ι�D��_v]�8�p�YT���$�$u�<$��\>�9�C�?['�W�[-�R�d�}Zd��8_ߺ�Z$�7*cv�k���Y�K�nJ�a�Z�hЯs3� o|�y����ſ��豥*�N�I/۩�$�Ae�e���g�:!XW�j�b���mo��M]�(��`  ^�;��h����--��)J��Qu�Lhٌ���]�
�K�Zɑ]C�xûw�L9�v��̽vf2��-��2�e�oѧ��5n��Y�~3(ą���m$������nb�o$�ى	/$����E�ݙ���<�7�ڜ~�2��ӑ:B��V �t�۫�Wm��;Z�b�
6��Is{:����X��!o9��bA�w����˓�*����Q�z�D�a�ښ	 �����f�9�s��"6���a�b�|����nq��Ł�6}�w��� >�0G�uv/w�{�sռ�����R� ���Mv]��I%�r��^I$:��V��k��v� {����0pŀ���tEO�ɈM0��U*�3�<y΁�PI��6m$���UI �=wR/;���5#�~���q�ٺ!XW�%��	�;.kԲ�p>X���z�UO6��A$�}�� �9�ԙ7�^�z��ܑ!{�N�6M�tt�wNUs��xv^,{t��&��K;CY�hs�?A����G?��;�Ϗe�:�9ɯ���(�2�$I�����s�9�9��xɶ�ZT]L8q��`{���n���L��:qu�H��	��Nr8"����x2�:湻oX�SntF�ۓp̽����y�3�壤{=c5��<����E���e�G�:x���ywNw,�%"p���۫5�Il�6�#t�v������gSX9���Πn�}-�rӰ�v���\�ͤq<^��z���t"��4)�U�|_���V�O�Q��޴��KWeE�@��M ��q�Kt�o���I ��R�YA��K8C�r@������~���@8N��$�I�SI=�F�	̩��d��}R��,pΆ�qk��ŀ������]D:���I[��H��뛉�ww��ad).���kW���G��s}H��Sl{���o�����ዕ�{���Y����k���UT) ��W���֨�,\N�qT�d�3 >wyq �9�{��[��Cs��w���Vȅ�UB֜�
���=p��	�y�+�E$��Q9*=�yH�Qߋlf��ښ	/.hRI ���ۻ�]�JkU�d��q��1��n =ڵ�ӵZ�_�
����'�nGVn"��&���\�]�2�=d��wE�sa���5�Ak+�l��j�Y��س�j��	�ʶ��˖��׹����	#�u4$�g��Z$����ueҔՔ�%Ubh^�f,��w�֞�w��۞Į�גIw2I'�:�;���2��c���=;��ܲ=���6�Y�]���(_n��7䗖t�U������[w��pw����M�3���	�AT���糏BĐy��D�ߺ�A$w��?���F_��N1�~?)m���nM˞��QN��]Ս�.��wT'<A��|E!V{�g�����!��W���>"o�	';�B�=F'{��~�5A$�{�-� ��@jQ�)������:T��:-@��ͮ�]L��$�]ݹw~I�Y�f�"��Gis(4����D#X�)|6B�z��I߶�,�9�9�u`��!���.�b�嶀��$݌��"`��{btO��֟i��v����6�-?����L�٦��n����$�v��wh��Y�ٓBc�ɒ�%[C�+�[[ն�*L�*��wi$�K۳f���]��W"�Ԣ�<����b���tH($K3H3Ӯ��wqa�h��ݭQ�$����Nl3��I#�u$����ٮ��8�S�����#�_�F�Ȩ�k�#m�C��^}s��dqRnWL׺�Ӱ��m�3�׾� �x��`�@'��.��K�����s{�c��3����_�����flR^H�!���k���˫�޴�^Gl� ?oyp ����{]�z{vn���RZP�]���8N~�h�I����򑮚���\ �z�����ـ/v��iڭe�9�=�w\i�z1��@��M��$�������e�:7�6&�9Uӕ�mֱ��#���eNf��gn{�Pﶌ���^�);�C�\���L:�N���n!^���x�fb�?g�ڝ2a�*N�*�C͟�s3� �w�5��^�N�Eu�>����;��� s��7���=�3����l=�q����rPƸn����>5�
�e��Œ�s9�W�� ڗ���|��0����*  ��{���n�s���z�>g��� �s��^�O�VsNB�R]=$w5��k`�g9&��.�x` x��b �ﹽ�b��c����gjxd�ݹK0�bTBi�;UR�I+��wi�Kr;:z�Onk��� �oy1 �����������&fQNI���49���ݠ�I���h$��v]�K�%�8o8����6��oyڱD�V;/��9�s]��цn�N��B�$�mE$J���˻E�ta����o��8� l�!�>D��=Z�>喽x��3Oq3�o���+r'&ael){C3oi�rw$Yl1��g��Zz��F]9��9)�h�1��߫Y�Mq�#7;qu؝���g����=<2]2k��6g��2vri���n��j칐,�h��=n�k����LJ.{\l83c��r6K�Zf� ��r�%s���J�νk-�}�6v�g{2�:8n�����t���|�Ϝ�67;G���=On��������!]*v��=lم�cZ���mes�v�@3g�<��kkf9H��8[��g� ���m=j*�#���VU��ߏ�n���?�ǝ�T>Kw{�I Yӆ�!x�F���b�K� ��s{[s>���mK4L�v*$@T��I��|b��$���7` s׏A�i�p��׳S&�[���v�R]7۞ִ����`���FF�n�.����K7�.Ţ�Ags}��n�P�/�RCF���s38������)�'w�k{�H{���C�y^sQ� %�szk3�-Z�-v�V&H�U�x��2v��=���������x��b�/)��c��۶�§N�ƥ�ݺ]q�W^75�X�;����4�W�)V����e��s}�5�� w~�� �oy08����ۙ�c�Go���	#�卓��q� �+ ����@�m�'?O�L���u���(��`�a=�͝����["�#:k(ʸ�r�l�W��bT�{�k�"&Zݺ����Ǚ���iy"P���PI$�Wu�	f����T�������� ��8kA�����������os��#��s[�I$��P�D�9]�RKj�a%H�0�D���}wlh[�^�N@���� ��& m�}�5M�1g���5u����C�q�)!�E}��)�	^��k-�췹�n,E3)!5�*�A.9s�	 �;���Ι������Gs�=��e��D!*+F2G��t'=��qh{��4m���|�e��~ꃞ�b�Q��ؘd�O��4Np����m$xy�����z��Ń����滋J'j��~$�W~����2I���T#|�^��,\JI]u�H.��M�#�0T͝���6hm�*�ǭ#�9�� ����v�I�gi:F�ޜ�*bl9��A+��vo"j��7T��I�'Xs��g6��DhT^��p�֛���R�,龏���,��^շQA$����wc�|�Ѫ���8f�g�{��_7��|�;�R�A$77r���	%�����1w�׼�[.�g���]i�U#����~�
H>箷��y)w���U��RIwn�H'Z�M�]S�5�T#!k��]�N�l]xdݷ��\/g��j���k����K�0&���z�
"���$�-u�(��Bq[몢	��m����a�Sb%��u054��'Й�ޛ$����H'ֺ���!�ʠK���&dLJ��E�x� ��`�,B�9g&!U�W@�H/7[`��k�	Ŝd�%)�M�c��ظc�]S�H*�2���8���V<�թ acߒ�՟�n7��r�v�9��螱�.���ܣq<�.����u�T{��Χ�y���?� ޷��m{��1�%�}�U�O�<�b�箚M�,���'�fOR��sFV�Y�
��$�J0'�v�t�`ۮBMKV*�*i���F�j*R��?������RDA�"'?x�<�`���A ��u@�1m)�C�T�WWlE��7j��#�����~K�� �r���;l��{]���E��$�sD���������oD#�&"QM�7Rz���$-����.���뚻�0��$�w;�Ӱ 5����=��-wԬT�o�S� �d�� ���D������( N�i�c�`�%)�T���	=������t��3I��25��I ��t������H�)
3��r���Q�Q�S�slʶ��[��ݹ����q�9��v/�}��@���N��w������^���8W�Hy�\}c��Wiԯ��s��˴*��U#��-��u���Y�x�2�Uaz�Ҋ']��`d��6��1hl��jS�3V�y���#b�HZ�ޥwCv.���w�>�[��k�9F��[��p�o�$�[-�
�\i��c�9�~L��ӓ�W�@-�(��/G}�/k�=���n�3�3v�i^�q�E�-�)�]�]��: l�v_7�����܈O-�ԋ��c!ɇ$�/W�M֌S޲.��y�{L���!+���{qw�G�|���n�`�n�(g�(� sXq��1.�gI\��QVɗ���f��_b|�^�#~{���b���q���=�P��f�8rz9�;�cRة��w��g�O�\��=�3��A�^���/l�O{<;u˚}�6p��iL�y8�C.'vq\��*����PN�3�^"��in��k\�U#E��"�
�r tV(�����zw��&n�/;��gktx���^u~�G����=�dEw"�s~=�B����I�@�5�{��Xp׺�)uڀ]�1����=��������S�e7P��L�;���+8N۽�{��x�p�p�RW�6�w֭9�tJʎ�۸�x����(Qb�,��E"Ƽս�����5As���&��tB�F�C58��ك.�&E9����:?�=����Da"C`����.�w���H��ab����W��T�)j����Q�ݢ$$�*�l�ۖ�eZ�V�`�XF
�FLn�F*2ThD�1D�[����H%�,�$�H���Z-��L�BH%H�P�������m�xG�=����KՖܬ�Td"��Z��M�������{p�S����eQۀM�ɎĮ��T6TJ�+znj#Z���܈�z����-D�QjA�P#�.�V��Y��R� nU����x�<����:@�)�(IeڵqFڶ�#�*֕�*�eVֵ-��`Ÿ�!��*5iE��[d�e�����)�"��DH�2Ei���
�HR���l�J�ch��LZ��ċ!얂E�EQ��iX�%�FH���ar�d����A��%�V,���b\XL�D�c����w+��r�A.�`����7��$˶�ض�m(�Db+iiKeȫ1%�JQH��"��$�Kpnk
Ҍ�&�i�!�!�⏝�]�����Gr{Y�uڡ8��,�f�\���e�v���0���p�֫Q�)�gz4h�ڠ��N��G.k�맷hMƫ��4O85g2�`*��L����X��a����$gi7�v1j�ݮ�����{�uϗlN���!�x����ӳgp�����!ȋ<��]q�n���܏m���j!�"x�$s��v�����M���3ԯ,�s�Q�5��kOq�M�q�b�y�t�ORq���FVm��nq��Pv����ռs��v�=����k��{kO���V����f{:��+�B��%�Z�o%��Y��#��[�;�g��ݝ�÷n����=��úus��yV����^;F�w2������n���!���p�T�lu����;n8[��v;n�Y��v��KK���<�g0q��5���uY��S�L�{v'lnl@!��`zM���i�kqB��xB�L�p��n��qIs�t9�ΉĘ�rq�p�2�t�]d!�aݎ�.y�6I�� �y�zS'�g^�����6�Bg���U籵�:�2���6`0����s�έ/�3��$E�+�9d�l�+=�{Wm�e1r\�a�)���s��ڷFƗ�G9]��.ی�ۖ�l�}ǥ:;��3�����=���jy�]�H���h�\Z:���%�5���gu3��&v��6���y:�(q���E��VDw/�vE�ey�n�ݟ[���@�a �@1�K ��.��٣[;p��um���ۗl�M�����e7Z9�mpK�n�:�sGPm�,�=��\��A�n���ř�lr������5m�x\�q�n��%ٚg9��j:sz�q��8�j��jj����M��G=jL�l�"㫋l�1�=��\m��%6�<�]mC��Kn
Nǜ^���.=��I���#8���ޛI^kw=h5=���/u�;d����Ѯ�[kq�m�ũ�7g�N�Й�*�tnܥ��t�b�x�#�E�S�`����ɛk�gg��W g��k��<��7�	^���G�x�oOl�)< ����x���ts����>]����N&��Hs�ힹ�ɩ�k���j��y��<Q��(|����w��q��9�-Qn�k��֭�TB!�"�w�{��d�$���!��7Mx��	{��ߎo	܍n��3�-���'�sc*T��
��Ռ�=/���G3
�U�x�ĂK���ǎ	ҷq-q��,���[��(S��1hl��H��m�E%��i��FEܬ���W�%���!�Bb%ߎ���yP'v����$���^b�b�U�97��t_U��ę�Q>�����>8{$F%��˺��Q$��o:��A��Li����Y�ҡ�H�cN��#�	$�4ڌQ+j��mY@)D%"*>mKT��Ϗ�i���6s�M�Y���o6��� ������yu�Q ���L�d)P�10aP2{g�L��2�	.�+�=ELq���M܂w	,�dG���#�Cz38c�ï�*.� mdN2)��t&Z�������ݟ}?������ ��jI/�Iׯ�7��ISF�:59�?~�� � /]X���C���0O��k�ɵ֤�8K���^靧���P�Au��d�p��$�s�A�\�so[f��0 C��J)�.n	 �<��VQ�v��v7���$�����7$n�66L%ݳ��< t��YW��]�T!\m���VS�S%O���&'���Oi����s@:=�_q��}6�Ft��sr$Dqg_���HD���x�v�6D��{��I��	���&��wD]���`�O2�~I��7���&w��O�o�� ��Cz7,��3fT�����i��dR�>��6��B�#+4n�ֈ~�|j�vXO��Z^p��~�����1s��jX���p'��������aD@�c����r��(��Aq�W�$��2 |�\��o�0O���6����� Ur�f|�i�}ʢ�=�۽�J�uM�Uē�y��Q��t��Y]���n��ɺ�&dL�fA�Y�knN�'���Y ��:�j�C�IC�rTw{�b�yQLD����A�$Q%��c�īz�䩴���������pvZ����ՙ�Arͺ����xV�O�%�ʢH}����MZd������G��D��B%6#1�O���l����7�dHE��I���A%�sa��T�S
�D�����iOzh�Ύ���g:��2������R9ݛt@��^�0��srͨ3�LB.���9}����n	��p�����f�r�)U���z�.��^��641��D-���t�n��[��!;�j����^f��d�/PWCh�A��0��˹����&��n�z�xMrz�y�o����������(�@�ʠI �n��_\�Ң���(���$���S���(J
b`��F�D�t��3����ɻ�A����$�'��Bι�w9�è��]�pk����3����*m>vby�W��A���m�&��!��x�)L�J��輩Y9I݊��ζ�$�yq>#�����<큠�M��2Ϗ{�	�bj��V�O~�n73s���c>���� �\I$�;�#e��Z���,��ݿ���?$ѐIn�R��m�c>^�gpF+�����z����'�F��w�2e�(
�g�ԟ��j�nl��~K�G��b�i��>�9�^ޝ���G;n�ew}�P��kN�:�x�g;���6��]�c4���v.���n�w��.�i-�wY�7�6��\�d��걹�^�ϳ�u��L��|��f��Xy�b�6��Q����d���lv�����<ݹ��o5��Be�sv�+I�M`( j2݌�N+�Ih�^�b�z���M��p�E{v.,@� �
�;_yί'a
��+6������Gm̐H���.Fs[��x�V��O�ܿ>�Q�:XH�,�d��bm>%��4N�;q�[�`_\H$�r(�T�訍��Ek�R�JR�d���R${H�A�t�ۂk�?Iݸ�7��{0D#3#�O<��}�����'Ʊ����j5�Y�	 �q ��s�R���2�<O��y�5vv�J.��`]Q>$�W<�$�_w6�[�^}��FѨ,��uIY�]Q��jr/<�i��p�ݡ�*�h�7juo����D7hC�]\H$޽�'ė�΄�E��̗&�"AS{TN\��TR&" L6k_6���>�w^��~j_���>b˫�lmLFn�܇�7j�𹪮vnx�Ἱ$_�k�[�����	5{^���k�9_����	;o�A/��A��������󞽜o��U�P�#��E�z�+Ēgkl�f��+�v��} �>��ͽ{��g3�$s
KY�w.R]�4멠H$��� �o�r苮W���\�U|��L������yL��c��k,"G]�P��so��~��/�y��sضpsjρ��vB�;-�km���V�nq=f�i*pu��e����=�U��eW���A��m�O��D��v�����I��t.=��� "fR��"s�e�wG(�n�&������$]�H$��2'Pw�8�tޖ2J����%6k_6�#odI!�a;N�޼�[rʹ�t�ٯ�y\]	�yo�e�K��wý��ٝ��e�s@�8CK�����M�b��v�����\;A���`���_wU�P�#��E�O^燿CZ�i���'ƶ��$]�I'���\��*���|��;z�D(bR�%6�s$�o�MY6����h��i��2�$7��>�s�Ｓ\�o��XV�U ���l�g$ݍٞ��Jtg`��%�m8J��uMA��Y�s��>�ɒO��wTT��SW�9��zz���A�� ix�D��B%7����fs�����ӕYt�}��>$�s^'ǗN�yu���=���!s	�J����N�x�K����k���|{���u^�M��
�%D	LWWWu�T�.�N0I�"H'ā�uT	����fCз��ұ)�Փ�a��<��1�r{�QĬqo���h�!f��s�.5_�J��q�lOgAqeo;�������I񿾉&�d�JR�D��"�L� ��n�EvQ�YzO��@�Of�
����s"�G**=��OB4���oF��m������pbx�6���à����ݳ^�I��\���x���{�2�M����c��WF=R��W�I�ڪ����BY��$�~s�@�߃�֮Ӻ����'w���H={�^�Gd�U��*;Ӱ̒�9�	2R��،��W�v��2	w!�ޙ���s�y�M	��oKK|ρn�n�A{�������D��׉$���OVH)A-u��Ct�E>� "J��3�ͲH+bH���S�x՝B�I���d	s��S&�X΋�5ֲ����n�\nIg?$y��h�<������,��gہM㊣��(m�X2
,wP�搑�Oю.�����{��Uc`���a���v  ��8�.F�m`v�]8ݗ��և��n�5�j�m{f�G��Ƹˍ�o�s�Em��]\۳�ݣ�7j��g���[m�t�M"�Ln۴�L�חvb�6'r�<����2ۤB"��gq�'�7g[wc�c���p��yx11�p�Qe�,���e2��ֳ�Mjk ��gRt��7N��+ms{y�٭�]��m�1� �p����vQ��]*.�οJ%��"�9ڪ�>���t�=Y"A\2gZ����{TH$�����	DC���)�jv'����=W�]���f��#�$H$�DˈE�V���MY=W!2L#2"#�##k1�O�V���td,}�Euw�$����'�Y"I8��I���D��v:=[{O�lp�d��O)�H��;�u}�[/wW��w�C�s�[�E�!�?sR��i���n�x�`cFt�ՂA��I;�t0f��y�^������s�_㑷[�ɖ��#�!s�j�5�'װ�q�?�������W�����;��v�'�+bA>$�M��:uH�5�/��kI���U7�Z�(P��d���
.����6+'�H���Ӿ��N�VP�zwV��
�cX��sc���n����P$!�{�4n1t���.����E�s���Ն���/�����s��� �OWH�I�}7TH*���{nu�V,߻���!����ǗҶ�o~���>���|�{�m�T���d��;��O��Bd�FdDG�h�yb�Esf5��S� !��
$��ZfC�ž$t�&E��$)L�Jk2��㛼�Jogh>3.c�M����vs`;9{g�}<}F�Q��+�p�	Ǯ�S�q�San��v�� I�E*߷ߘ�d�7hC�~ԯۓ�L�	�9�TR��3#˶@�9��~9��h�L�f�uՁ��a��moF�H���~ ���A����[��{c䥄-�d��{Y��h�v�$���ﶍ\w[�r#�w_B{ƽ�3�ٻ�vx��U.o;���-=;|=�F9��qA���c�C6{�Z��
�ȑ��l`�P��LҲq�Ze�L$�zk�w�|��垃=�W�J4�^�7�B{���{7q���w�2�N�$�O�[��ĕ<�P��v�9���{[��RK(`����6����@���)��*=��J��
����N�r-��Zz�#k}�%���z��|Fyjev�v.��6[2��~�EL�]��y3Z]w�'n�Yһ�u���h�_�g6�"3o�^�Ԛ�Ws"����!�=X�o�e�����]�L�.�t�}+����1�MVw�*�SWGF�O�=��+�0��6�~�s�9_�og�\����7����{w��yf�{�[G�26����ې�KSS7�
�>��v{����#���B�V�1�	�슨��.�){�-�H8���9a'��;�Ý=��7\�v��:�XQ���t�õ����wcI�31/�O�qw����Vo�������G�x�~���RK��x�b׷ش��]DWeg�;��n�=�e�����[ܲ��2� ���v%�y��ri�y��2-�1�B�}�{���q��H�����䷄8�pQܻ`[�;��6w_wv;L����p���P"v��ךE��y��V=���Ś��|�{�0��ת����bp�<Ի��R1V�#	%WX��[��w�\��2�E�F�S2�I����)�ik��-�-�,���E..�/ �^NL��1�|ݣ���!.UT�[z�cE��F�]�d	r�J��j ��Ķ��R�S�`�.(�
�*6$�$jS%nm&�QrB-ܶEQ$�ն0�EV�����Z#QX"�k
�$�H���)inTK�kCJ����1�iE[`��J�*�W,
���kDDL3�����\5UV
+
�rʂ���-��1F�I1��I@���BFAQ%�UT�QX��*�L���4"+IQ�.��w-"�*�Á�1��ТkƅE��r5jIiU0�a%i��I.F,�h�KRҡ[������V�ZTU�kh"ň�6(���E�ĭ�EDA�M1�qЫ��mF�kE1T��!V�[�HI�������LA>=�'m.&!8"`D�L)���S-h�������I#�ͰH$	�G֜)��9$U��U�M�k�]�fh}���Ѷ��o�����'ӹ�� �v7�~���N<Ś,�n�1w��9�_�e-��l�8���ON��\Q*5^���L.���2ff�^=a�67��@��p�]�l��O�6	$�v�9���(0eIP��E���]���mU���L�@��m�ͷ�7럻͊W=���e������a�D���	(��8,etu�;oxI��o�	����L��������BsՊ℀z���I�"I�;���qD�7�g^��{b�Oj^�&� ��G;ˈm�7�U^�4��ʼ��]bU�N�Qb]�V���HӠ���Q�������".�XgӖ����2�~1_@�	?fWS1:˂|�y��I��H�I=ۍ�������&�RJ	�qِ<�n�GZ&�'�Wc����)󩒧�o��N7j��L�=8�� �lH �7�f]�V��A�����	�����B%7��[lM�L��y�I����ݸߎ��{�"f{��]�����ZthE���$o�]?NA���������&w�H$�n:d�갶	���2��#+�m;�
�NmĒA��`l�4�X��y�� ��N����KHKV�GV�Y$uv�i�4	�>�H}���v���ٷ2S��q/�ҚPD�Wl���$��r+&`^����=��5�h�W��7l����Bē��F��o�a�]�b1W����}�f �o��{z6�[ni�sə�����3^{c�굮S\�����]�p��g��^�DE����ۊ���� ���l�]�Ⲏ���E�L�:��^ۏ;�y�\ݨ�Bݨ�on�֮�/t]B����h�`\f��;u�iʽc����Q�[fN�ˋ�Y�����5���t�c���gn�Qmф�ۮq��� ��^c;�r�z���rC������9� ����2I�޶*��T�S��Lu@�;;?}��	�1����̃���[���D�$�}Ϳ	;[��t��lv�=bɁ|�_��bB%66u�d�A�޷�|H5W�����(	{ͲI=[�L�W�0���%B�o�ofݡ',���{��A>�޶�"{$<t�#X�Ӻ�>ͫ`�
I�el�>��lI�pTk�u�	���o�Od��ދ��{����bqY $�����6n�퍛���;���ϛ�­�~-��)`�{�kZM�v�m�I"{$I5�qه|2�<�lE�����j���<^�%2������ͯߋ�;m���H�My|�X����<�C|�ř����E���Y2*vb9F��u��#�I��y���Ş��7�*��}E��8�k�-�%�&$�G�h�x�&{`I�QY����n�m�I��H�`s[d�%��M�s�~����Y�>��ω&r= ���GF�2l\|{;u��P���*z�A ��u���̨��x���l��ݟH$omca���u��snG�#��-,J��u�w8��#�n���&X�P�+ ���pt��]�Ƕ�$΀'{k=px���Lյ���b�?r����%q�=�����g�D�
�y�l��9�$�����Au�J�w��J����ǲ`#��Z��(���lI$�	 �s���3`������i3̻���;_��A�e;}_cU��쏹�|�)�>�炃޻�%я��%��|�޾*���K��|
��p���>��<`������$p���U(a��O� ���[�6��U�"5������joxe-Y���D�^�k�]h$v��l��\��ر�r$�^V����o���p����r-�"f
1��r�����v�𣖴��S{��#�{y
�￿���{�nLe�S�n�U�滭�Ҟ�y�q܈�� t+N�	���t�KA0&a)IK`�>��ό7�;�Uq����	�X�'ăռ�3�&���~�v̝S0L�L@ɩ���t�>"6^O9��"�W6	$�o6�킹
bLIS��g���S�uL��3i�0I�������6l�|�uy��K�K�u��x��Zru'*�FE�j[-�N=R�߳A���dW��qy�V��*"�`DԼ���ԩ�P M
_���`�k���6eܬ�?O�gă9�H3�%�x��ZE^6I]����7�$��X,´���k	��ۢ�ݤ�z�]E5vٗ�ݎ�Y�Cvq���5���H2J�J��Ͷ� ���ߘ ��y+����]mTד�m���l1�1�n��2���6�3��p��rk}XH�FVsl�7�$o��ju[�;��Z�3	JJk���l;�>'ăϳ�s�n��a]����� �ʜ%$;�A[��5�޹Ho�g���ސ��6D�������.5~������j.̉��`�8�H$�s�f\Ts�U���s��$�d�������v��V��8c���S�PS������^梷T���ʘZ��Mfm^�ꁢ�X!�J%u���҇���< �;~1v[�b}��j��+����um�֬��Q}�uq�9g;�������#�dM�^FWS��Nv�X80�x1��4�5�}ck�����Ov�r��C�/fC�m��3�����ˊ�A�wz���ٸ����n�3h�#�l������:ŋ�h��qr�֦��PDf�颔��M=9].��7V���j��Z:�Nqь�3Y E*���_�hDVC�'��sZM;���$��x�Fi}{{��9x��6�3}IsYd�$�����֓㦯33K�++�w� �͑ ���x�=v�s�w=��d�%��A������;-�0I ��$a��	����H"s$I$�s��t�+D0�SL��]��s���Ǳ$k��~$���^�p��,M��URo=��mn�U
E��g�~$�v����Iv} O���d�g�������2wuʣvGQ�Zab������N)�툎�p�4���Q�y?@���`�}�	7���$'w�?�՚A�ys�&������\x�T/L��Y^z���یBy\^�;�(�Ʒ�����FH�Ȫ�c�q]v*6:�C��Z鶧 e�R��E����K�3�> {�S�� �w�͒O���6>;j�z!�Q5&�@���&S&	M�;v�'ę�������XL�>CM.	��V��	sy��9>���P��@P�uB��n���ac�u5����$Wd�缷�;��9���>��%p�f�*[8�[`�͉�up���l����0�H3���	"�$I׻�hP���(��ն�^<��4��dP�8������ۃ�3������٩L�2�H�*:u�2L�ka�+������m`{/[u��'��?V�����!�'/eM����3j���o���:��I��5,]97�iq.<Q�*�h�����vĂ	4�輻�dHY嚚<�e��=˶��������|��W�?��<��3���B��]���0Lɛ:╜t���������g>��&��b��I�TɂU8�z��;��"iEV?2	�5yI���uuHU_V�e�]N��~gǧ�J�
��I$��L�Ʃ�dP�����5y>�����2�وf�l �X=�������9�n!��]�fְ�=1�DU�����͵}�B�AP&�*s�u��d�͉}���&��V8J;v_vs`��W���8�L�*$2�W���� ��9�୷�����>�t�Owc�Gdp��8"qՆEs���S2`ʄߌN���}��2;#����K��g)��kr}'{��$MF�Q��^�z���T������fh�nbI'��9�d��o^�	�7��9�ơ)پ���������fOq��(�{�	��u��[=3����+0�;`��MU� ��X"�,å�{�E>�}�Rߟϸ�q�����{���#7�~m�ЯEvȐH'�ۭ�O����AJa���Z�伦IH)���v�vJ��vu�0�R�c�j �$�T$uo}���T�PQ��P$����|H1��L�̈́�d�Ȉ��ݜ��>ͱ�h��J��T���ОF�� �gTjs0�	'����O������V��g'\�{fmDL�1�P+��I>3�������齮ׁ�I��m��D�v6kX��J�
T&�Ná���ܞ��h����>����꾐Di쪩/�����g ��B%B���x�$�΁�nf�����[�'�k�~/:D�,�e>�~��=�٧�_k����M���g/h�4)��Avo�wK#<=�Kce�>е�݅�vǜ'�4g��yL&c��!r���[}w������{'�j�gn��Wu�.I� ��.�9�9�ܸ(w��;�v�����S<;D��&L��;AK�k���n�hk�������C���a���}/�6֗Ϸ�\�~��ce�������q��Tx;T�φk�6V�+W<Gm����z�b��b�'���A��
���ٰ,3�L��g-�i�[�����O���Oݷ<P>%���;
pLW���q�U�ڃ.��^�,K�`��r�j]�Mo�{�7|���'�=;�B�z�A����7N"=��+NG���;�m�e�<�J��mAdsW���<潱���Ǖ�rpx|d�_'���KPW'<{�4zc�݀[���a@�'gz�y����e����|�����=��|:�NtŻۦ��K�����+���<��o�Z^�L��[���R6�) �`����=R"�x�!��<u��#���ݏ����S�u�J!]�CY��׮t"�toz��@�רc��Zqы���y��]���x��cճ�fQ�К�so[!�N��]����a�N���a�8wS/"q�{�S�+z�jut]{~�����v�/}w�f�������5�F��{�%�Ջ>�ޖ+�4�r[h�X��b��NBD��:�1͡�)�)�(�eA�����[aFE�T�1qF�Q+Rڠ�@R����*��TPU-�&2]�#lUZH��D�JU��@�C�*�-B�"�l- ����D\�m�4��LHҩQ���ƣH�%�*"���AUb$FU�e�X��HJF�V2ڃi�.ֱ���C��]�V�Hҍ[Pi����Ū
�D�ڕ�ʧV�eA1eX5�J���b�R%d����������hU@�X����-UR,IPU�1b᪂1��E`�X( ��"�,X[Vm�X�(ł�E�QE�q��V�Ŗ5����6ʂ�d��"���m*Vwpw��]�g/�l�L�^���G\lq�n�ڑ�뫝��ۙ��Ynʹ�\<e�ԧV����}O>m�p6c��y�9wW�`x�Y�z;��6�g���:\��0r�nK5�[agn�1�����n|�La2]:�C�����r���=��;���G/m�q��{[���l�n�lqg��f��uӸ���<����L�E�p=��h����Y�v���؍�jtg�;�x;G�n6a�c*L����+�|����6�g\lVr��6�kVqϝ�xt�ݕ���D��j�)n6--�W��y��3�N��cIT�r;ɣ�u[���� �rX�s{�8������۲i�q�����d۷c�7�Ώ������f:2�;qtA����Pi�.��tr�ܻ��үo� .�g�ێ�]����k7�sc�
����7�f��8��n�Ջ�pҽ���v���g��٫�E	�������nz������nV��v3���ЩWX;]t{g���4c/=�p�qnܚ���;7g]�zlY���ɓn��]uKGN{�@���<qV`�a�筒�\�+���vW!^M�{6��R��ul��xH�q��.dZ���c��xz4�vn8ؽ��g�4b�āl':����F�o.EOm�Y�ʛ)�v$�˷��G���&�q���n�e��A���݂ R۞��������sc��xi����5c]�9�{#�.'���[v�m�<n�W���&>q��̋4=�ǣ+�:v.�2ۮ�m�+O-p��ǷB�q��Smun��ƺ�{.θ�(��ש�n�[��+�_7i�\򘰙�ڧk����ƪ�Vj���z�8{���-���u{�Ѹ�ή�v��&�0��:��yBW��P�3��٨�;;v���jw���Y�û�����|O�Ӛ�#�Mu��^oG*�a��<p��֭l���]Fݕ�Ktؠ�X�kA���cmv2�7d�a.���,m�>z�Nx��3�L�k�7S{��7I۴s�c[NŰ;�!�t�<��˷=;t�����M�"M�MXzD����w/]�ɛe�6��W5�".t�jk�❮ٞ�Bm���Fm��4mk�+���m��z�V� �� ���B��J���������P
�����$eocgĒt���T�A�әX�#k;&,�
�3	PQ���$��(�3o��wV	�vs��t	$H�W�6�n����^���i:�I`*b��t'�o�Wz��}e����NOnW�Α �ڜQ$��T��n�tM��4A&%�6I%�H�N��e��G+���~rL�-���)f�F�	�w[���D9�n�����O�N_6H%�ȟ|N��l��2�d�{9ekS��  (�L��r�����m�u��n1i!\�X!O�L�=o~��QR[��}��_<�@'Ď����3.��64F��������NL(��S��UQ���0HQ��`S5d,+q����P����^�.�gH�b=��z���f���;�6�K����3X.���u5��������/����$�H�{��ٹ��{p2��nu�-ϝ�����*�oǦ�i�H�T��^tFoJ��	�D�ӷ��ua+D%T̂�����>�i�Di�W  I��a���������>�#W�˲K[+�GJ��^޴�n��t�r�"oz��ݽ�b"��]��`�Mgu������4;�&dHJL(�ǭGS�v8z�\�д�q[��� 8'-��A��?__�'�\	�TD����`�s{)���O5gA��>��
���zf�w<l�N�v1��E,�'�����{L�D��P`ν�6�92�V�
J�T��#�hi>w{����f1L��sI\��yw%�����i{���G|`8U�7n�;f�K���0�*o�ō�����%�*����� u��	f��?o�L�3yL$eADY�g,�E����h2����O�����P7��m�V�k~$VnAZ!(��d%-����$I혣U^̭�0��l�H3{٭&�|�SSjf(��yr;F�,��d^Ӹ��j��n�:�Wv�����u�S;x(d�}���ՠ��#��ն&wwd�I��r����ד�\D�u����ܦ'_�ʙ
T&Ȏ���o/z�-}}t8�v7�A'+�O�@ḫ�����=2��\,�r�4�u��6Т~�a��:f�fЌw�7ę��`?��%W,0�(��TF�U-��px��N0���ߙ��� �y��LNZ�kj�V5,�E�s�gjӮ�j'��Xv�"wv�E]�20�[o3д�����e��	�Aaϊ����{���ٞO~n�ȹ-��/�	���f�f"�fd���[��W�X3���G��wv��q�"Jչ��U��:�/4#������
�Y �
��{܎u@�*&BSb�[�� ���$�O��c`�̽��'�����i��.w'd��G/Һ;[�eD��Pe�uyB�&�@$���d�rƹ4�L�R�z�8�҄9���I�L���>$��e0I@��Q'��	g�A����R��!�3F'{,�FA�m��I��$��b:%���3�5�B�J�ED�)���l���ox_Gd��v �	����$���Q�_J�Ϋ�51l��7B��E#���ll6���^��-(���&,N1�j���c��%N9�y,M�%���N�]*�����f�m��U��ϝ��U�& ��ˑͷm�}��:{����M���'>y�j�̗��9ۍb4�s��۠U��s�N��\��sӺ0y�˝���km��Ϲ�Ј$��v�[^���n��v9�n���S�KcQv��9�x1'�=l%�,�l3�lŸF�WX6
��'��+���d�5�m!� z��r��0q\��Fy���qr�l�8ŧ���'�p����`�ߎ�|�I�r[�K�0��{���)��م���S1$��l�]�"7	:�԰� �?Y ��i[f�$z��0	���l��U��N7��+"&	PbDI�]��~$c�q�A ����Rb�:�M7#<Dvm�8��.ff&RaS�T���)^Q �v�'Ę��A�q6;ʪ�8J�&�[$GT���B� ̅�YXH#9ȓ�][��[*%��%y�A&7{~ �8�D��6.D��
�WB�Q-M�-,3\�S�n�<���y�qn�Z�o����J&k���֓M��	�&��3�9;�n�gzsd�@1���0��RI�.ˑS��R���Ȍ=!��5w��RUV����7[ą�g�~{�m��ƷqS���	b���sfniДO�x{�y����I }����P�m����^��j��(��d%-������2	i9
"Ν�`���l;H��DŃH��Cq��['~S6�0�+����Os� �k޷����1�5����J�bf!&`��$w�t���9�Ȓ�}O$c�����5��5�/3�k�`���U�',ePR�,zꡭ�5�V��'=;	�KH�q�J���ε��ж��0|�s�$�=�l39��zk4��Y�?x�H�Ұ��&DJ%7���Ac0X{���=`�|s\H �޶� ��+���zWD�A��0Ǌ�(��90	�ͺ��j����^����#����uoLqB2���S�vɺ�����e�7Z1l�gN�*�j��z����(�v>��jAs߭�}]��h&"LD�J[i���{��';Ėc�����~~3��P�#Ouɖ,ӥ$��
ă(ĉ(@�uU`�	3۸Ø¹WL�^��
](H&���A���篲�����~��~q�r��܅�q���<u�^��tm끞9���S��\������Q�m�|�� ���e3˄��:�b^��$O4AǚwB#I���:d5�yIz,ʃm
�>��߁>$��c�iD�Pc�Bx�]\X@�%�9�߉'���c�fɡ�fb��P�ۻm�O���S=��x� �@F���gB嗲�77�0	3y�LO,��D4�pJ~����A �0&)�������Yu�g�Ƣ�t�.$�P�YuB٣gGL���߽� � �}��"��F>�L(�	CU��	ö���$d��}�7ę�ܠ�喤�E2�w�wOcp��q���
��������v֬�6�3ɍ�p�ڣ�WJ���U:�Ub�����i��{�)�	�Z�����M�*�m�&wwdV�(C��2 �0�2v��B��"���[i�U�ANf�`�ye� �S�U�=��ɮ��=R�""�I���$�;s]q9ʎ�eKʎ�x&o7`�GdY�Tyaa�J�N�=v���eL���2H'����u.�Tec�	5�x� ǯ��$���i�;q�3��3{�uf&�#6��$�� �z��6�8���& ���ŉ���aq�饫�J�t�w��GQ��������iݤk	-Ȼr�Fvg%��[{�����x{ӛ�����a���z�=s�ۮmg+;;hU��򭸿u���GP�y6�O\��:��r\q��<���w������!ۓY�k�'c��W�v���l���	������w=�\����y��G����܏7>�κ-�y�dpm��E k���U�۱�r�k���pk�v�6������5�v�g���u��n\�]p�i�Ǳ�9�ⅲ�0s�ݮ�6Q���]���v7rJ�!no#x�L��
#?o[�3U����͂Jڒ�%l����g��ڐc�!)�"�n����ɳ9.:�2I;�dI:��`�:�"#)�v���.�S%����������o�&
�z2�t����Hދ2	�޶�J(P��F}&f�g<9\��3�9�eI#/:� �7��Qp9���I+�@�D��{hi&w{�˞�"���.����k{��A>3}�ؼ�;}��׮�=�R�,-��n�'���rbx��ꇰ����IwP�.�7��`���:���{6�I"o��,jю%Q�]�]2���~rJK&�s=��M��m���U}�3��_���fE��n]�u$�N�Y��t}��gvy�<�}�zg�\�7�oSv�!��K����wȂA�3n� ������!:�m\m��H��$�2J��+ù������ʉ#3`�B����t�'ķ}m�Io���k�8��"	�	�:�'�\���$ܧL�L��S ��Q�6�'!mV6	qH�B D	����獃�ڜ�ں՘�זM]�6A;w{!���M-��^�=x�/Ŏ��L��U�8�P�|"�j��� �>pl��!_�-R�.m��j)F��K�����Gbd��ldt7�m�	37�=��x�$� ��Xl�Y��jw3��h �ۍ��{!���N(��`Vn#�A��Q2C`�>l2O�jr ���HQ���ξ��~Z�]���^���
� ��/��^8��R������]�V͛����eg����MO{_���8��rsp�N�W!�6v��|�!����Ay�y6�����[��@aS�ZS���x�sD���j��;sgo9S�:���|��4���XV��ĺ½�o���2'j
IG��N:��X���w�0P����plӋ�Nm���f�vj6ʋ{���w�V�6+1��w�x([��y?z]i�!u���\��E�qG[���px%b�<���U�ޝ�i8z5�׏_zף�gjt�u"q�$}�Q�����=�ड़�R�]+����W]Yui�3u����mAg��A����[E�j>�=�ޙ���<O�ś�{�K��h����3D[I^:���#<�۪I���hC{�G��<��JdS���v���"^����l��{�pn�������}+�Ա�;y{���Sї.��5Q�M�Fma�J�Iz�BB��Œ���{��lv�{�g�yޘgy�C�*���n�A���U�U��>�	yo���¡��������=�xu�6��CTy�kOQ�&��+:��	7$�{��z�h�8|��am�;���ys幺#3rg22��	�B
�P���U�p�Jh:s���sY�t�[�<Y�{������R�/H9��ŧ��Ƿ|��+f��{<p�+�DǛN�t��ιw�/}�㳱��eTP*֠�Q�aP��%Q�V�
�6ƶB�����k
&�+"���-[j����Q`�J�"��+$������6�L+&�0^���A��,U"�(VTX"E���U���V�Z�HT�L3	0��%I�JDX���b��!X,�Յd
�I*�-(VJ��eHTR���m��eXT¡X)&��+
��kQ��Db�騌"���PX((VV[J�VT�X4Vä��-��T!P[[ ��B6���������ϔF8���޴+��Ns21J�d�I(v�7�L��ŕ��$��a�A�l3$�|���CJЕ���s���<�&$Ȃd�l<�Q'��S3��S@��WM�E�f�Fbf�����i9�}��G��� 5i��pvn��\���H&T�������o�T���\���;̀H�9�y��ʎʯoY�Ҁ2��x��4+�4Q@�D����H�oUeYh��f�� �x�� ϟ7�M5y���iD� �{�!!$� ���A'�^�~$��mEdz��J�vfE�'č|��+��$�)Q0CU�b���t*�n�`5l��o��>$}�b�d��J�[N.�ٍy�l6��{�BX������/�}�����E�9��D���eF���`�ϣw[���7Yf�.�~�Gč��>7� �HP$����$���q��L,Z�6f���� �[��U�cbF.�]�]���W-B)$�>j�Z:�rk���n�c��z^�q�8,$�j��Gs��'I,*���0�7z�� ��{&->ꚩ������ݷ����H�B (3�1!gVc��z�v���{L[�Uk����`�IW��	#,�j����(�ĢSb'�[�$��{ �]t�E�D
"3��S��<H&�^0�^�0ɏf�$$��r��c��K'�:�)�I[��?�qu�Y����m�W�	!J������`���B������=T�V�B��o�vE�76`Ou��g���Fz�RU-VV�w��1�� \+²����pּ�;�6.��/=��m�ӓ�טH]Ws��dO��Ix�Ÿ�i��փp���eF��c:թN�(\���;�|����u�yn�NyMx��b���j2W��y2����6�q�OF�ϝ�v8]��.*�.{uݭ��%�5ֹ��ORo�b��}�:�s]�y8W�`��%�F[��m�[n�V��6��̅���t7;������;jv�SK0v���M8Q,u�n��y�.i	�2�&z}]E\ݝ��W�C��QG@�7k�>�G�Q"B�$��*�`�@+7q�A�dc�Q�F�m?lK̛��lI]����9MXU�����S�n��c���WH$����vE��*(�����߫��o�i�i���9L��v�6.'��^�6'�,�>�\q���J%7���Qx�vT9�{�A��d�1m� �|��*s{5�&z�dt!��$� �3��$��{O�۳�1gf�1���� �|��h��9�Dy��N�]�*�H,`}���qٻB[��N,�_8�HV6Z����*��%���y���'\�������G3�5�2mFW�M�0�yu��`d��"B�H�o��lT��0� ��*�tI�NN��K-���X����e}�Ώ���u�n{6�V] 0�f̼����L5��o��ne~����]v��$��S�9��L���L�����߭�L��V�+4a1f�A��d�l�۶�'�fቍo����q �u�[6)hD}&&���ʱ^�F:�'*g����'ę��9t�n� ��	+�4Q��D��;k�gw��ݺz����~�ĂA/�-�	������/vd�A�xa��َ�>z����N2is\�ó��Goo<W~xq�_,qr�&󙊏�����i�we0s�7�^�/c��@%��o��a�Q1���o�d��+�v)VI"���	3{�� ���EF*����{ff	"��sm�I3�����]!��#�횪�79ֲ/�����l�:]�Uφ8�4���Cv�6ݐ���[�[fFa�����e�d�{�Ml|O�����H���3Z�(s%H�d�l;Qsi��1;�OĐf���A&����Ճrc��B��O�u���O���c��d�3�2�[r�=�yWZO�o�+����K�.��T�F�8�b&+>�m�ЅW�NUSW;4�Ǳ(<�7g.��IIS �vwRDB%���\I��LI7�V����b�6I���00�JI�A";fG\��y�Vx�L�v6H"��|H;s���:��}��j��	I�II��g[�� �F�Ȑ@3	�.4�eP[׼O�����$�3�2d/H�"D]���z�ؔY ���`_\I ��{y��Nݑ�g���8��a�w�@��j��we�f�Ƹ"E��Xsļ�S�e�6v!8���4\���x�r����PZ�2���Q �w�e?�-�gT���[$���G�����hU�+��a<�n�Α�sI�+��X�6Kz�G^��.���vR��nD@B'�T��g<lF=� ��{f,�
ڣ��Ӗ_:�>"�������$`��Q)����AGr*�h���ʲ:�=>׽��O{��_i)(݉y�l����p��/���w���-�峼��kli&�D���{�i��1��
����B̝�k\�>�q$��l��v+�e�췯���I��s!zD2 ����>$��a��wU9��yq^$>�oĂL��7ә��D��r#.8��mE���xi������,�Jz��xMz�G-�<�\;*���79j�.��,�κ��g?}���6�N�h��^z7nڭ����Zgi��F�e����/:��[m���;�욋��v���]��ywm���ոmx���Nہ}z�|&���<�G1B�;3sϡ�@���8�r�a:;d��R����ʇ��pU%&ʈ�n���j���ۍs�UYzv���f��9�Cƺp�ݥ�5�x��x�l�����0�s������#Oq��μ��h����ҧ���-m�ᚑn�r�'ē���o��)*H��s=0QOs�����t��%�X�W�o<a�0��r�Τj2�fc`�I����Wyq
]E����Z�P��Bn'{[�A����"��R��� HQ�ф��ٍ����S00�JI�A,�
�������'v���$�'w��I��8�t�����5zr4"��)I�mW<d��dK��F��'�v��&�	 ��y�:.�o�yr;up�URE��E�k8R�d�mmrk=r��!GS�U�U7��Nʏ��:�</[m�|H3ݸ��[����H���	w7�������I�)��nT�rY���jN�ag��b�7�n'R��*�K'�,;����������h��֕!��	k� �;�H�^�lRn��B
���(� �ʾ��$�g���H��I$��=�^}v��`Ј
�LM�`���A5X���f�nV�NQ�Q�{��lEy�^.��������#~;��A�%�2	�_?2I�	'�����+E�t�$�s�LN��$� ���_��7)�AD\	q���}q �O=�l9�wy�m����@V�,_�"��2*+%��U,.�7Hכ�����]�<�����_��1���ܿ�S���mN�����{(�.�;7;�b��	��A3�"2$/H�D@v������p�7G$ˮ��d�M�Ē=��v]D�yo���[bBb&T��ꨒA�����q�\4,�8�����)��w;� j)^d����W�TM�y���i��>�7QZ��;��=[����Ǫ��tA�c�������sn$�y��A��&��Ϥ��1��r֓�Lx�l�� ��d���d���sK*aP~ ��yK��:xB�m�����}��Qi����k��ߚ|:�6�X8�ޡ�� ��k�s�6ɱ����Q�3ߞ� ��S����?U������mTP,��x�����]�ѰO4jn�*�,A�|*:�ߺ���.\'�h>49߰5N��HQ$�y�2ke!Z���
�=��4�h&�������ֺ���(ƴ5Q
$�T7�~�&�n0�)�x�x-e�2˗�8���'�Ͽh�U�{{ߜ�þN�=��J2�X%@���4��k�H[L���7H6RU^�}O��~��S�&πD/S��IgF&:0�
�I���m �q���T��̛m
$�,aXo~���>�����cG���"?~�tm(Z�5�5?{��'!�p��9���R��<	�=U r'(n}����Vs��R�5�;�M$��0*^���N D�j$����d�{�^�n�L���;U�d�ҁ����yT���w*���LFV��zL&��\c݊5�������2��@����q�4I��p�vKr��Ѧ��D�{�d6!���X<��1�d����q�Y�w�r�q*��w�l�`V�-�\��d��
A`��}C�,
��s|?^�O�]G �r��l�UU�9I.ݷ3	��I�����1WA
��j�us���dr��䗐/?w�6� D�jTL����P�q�4I��ڣ5T����z���f}|r'\�\ɶM���ed�*u��Eq8��t��d�˄��hs�`i�Q$(s���ϥ�	�9���D�k��{��M�
� VX��{�J4%D?g&��^ۜ�?9���m�#D�|��X�2d.^��G"w������J2�|󾌳,�e@" d�!����~�||(�Hg�{���P�Q�����4k��}�%aux[�"lJ���4q;���K�z��3c%e*u�sy6$�AH,-����e�ID*���d�%4���6g[�d�eH)�{�̓q6�M����e�W&M�h8Ƈ���IAy!��@Ͼ���D�K}�X��	�A��{`q(S�j$��e�Y*IP�C���2m���	�|��;?����Ob�l�3�]�
�`Ww���P�4����ov��z���髞�>�psCWx[��	󏧻�F�i���ܣ���dm�xbm!�j{���qҼ����4�Kw1��๧��ly�잕<I�x�!�ë�p�P�N٘Yn�Zwg�a��h���
@h~��޻��۞��o����Z^~y���~g\iѺ=��d��C�^^��]�3��A\.q!x�k|t�2��c�f/r�=�.ԉ�ڋ7��[���Ӏ��#7�`�=Һu%��U��w������̪=��������9#(>;�)�|�����:���}��<��jj��DW������ݶ�->#��N�X�V��l�s�����=ǵ���C�G��y������/t֯� uC7�tuyp���4յt@�k���֟1'k}�x�����-M
إ����8����#�)�����i�Ғ���'��}��ޯ]���a�f��+�{A����\�q�:�6��J���ϵJ�1���u�����Hײq�H���Ƕ{"$`0;1uբ���osmL&���1ռ�u�7}�!y��9qxMC�hۖN�-�=޳����oo�>�;��O�7�S|Ƅ��vqx5���W,O�]���ױ�P�SV��=p���1��)��Zݠ2�>�}�W'B����n�����sz�d�n`�y��ĩ:�J�7955Є��HW�k&l"�Ntfr���!��ZʫAE�D8����b�
��"� VAdYX)b�-eIX�DdDI+TV���L!+2�ZXT��!R�T@R
T�VT���"G.��-
e)S%TTQJ���)m�Y"�j������TPXt�8TY�R.��+
ԣ"�E"�i1�En����[L�@�kIYKeTm�(�Ҫ�Rڍ)iQ�EX�e���R�K�E�F���F�U�-�m�)��a ��S�kQH�E%e�F��FڅYD,UA`)*2g�A`�K�+$T�b�JJ�K�LZ�
��aP:Jȡ�J�Q�*Q��ֵ�UY�U�(
a
��"�TY"�j$��J�n�6s2f8���<�y4�Ŷ�h�{3ksKٻ9[�2ՍN-���'�q&��c9��t���oFy��.5���׾|~Xx�
�p�3�틵��ϛW��5���s���z{Xܜ��܎�5n'��Ϸ[n	�t/f�ʲ����r��x�(����h�H���s��ǎ�n��hqӷ����y0�k9�nu��kdp�v5�9���9���2���l���&k�Q�3�۴D����67[���c���;�@�9V�!\8������K��[�������2���w=���s���F��=\�vM���x�n0����#���۱cv�[ܷk�7�ژN�gf6�81b�`(�]�Vpexi�-s��d�A��|s�!8tvz�\�ev����(�����F�vzۢri ��x�:��Uol{�[��/�g^z�۠n�{]r��wϟ#7����;����;�fv��3���8G��]�ޝ��E�ۇ]�F�8�t�nqrD��s�i����ɂ�4B\�P��e2�M)xwz6C&6zz�X��\�8n{O�\��޷8M^q�bv*˶��7O:�볻ֺLpW��C�n���mȣS�q�����hn!\�(4UpuHm��jc��v�-Œ<璷:�L�C��\���[m��v�h3vf8��m������Z���Q�0�N�d{'�:��;�k����:-�Sq�1���sγn3�b�]�-v8���� �+�SO;;�`�&6ڲkO�.M�Ӊ]pv�.z� �m����ۣ��C��vZ�l�5��I��3��˝�ױd��<쎸ښ<�n{KVw.c����/`�^�����ڴ<�md��ܜn(5Q�ٖ�U�W3�l�n�j�6�8��s�<kpq�웈�>3Gv㪽���B6�ܖ��.$��
��cu��Z�_⑔�1�*P��k�Z�R�0Ӷ.�4����;&�#�
�2(�EEh���&)%pT@�v�ם�D�ۇ��0?��s�'�H��7=�v.�:Ȗ:{A�Ĥhv�9��ʖ�}%��p']�ý�ٮ<�Ƚ�ٻpV�l�v�i��m���U�v�G��n]ڥ��6W�,�jÁ�뗙v+��U��Ǎ�sĞ8����U���Pm�R*lJ�S�[%O�����z�8�C,>L*uߛ�!�!���YX<�����%eH(�߼Ѷ�|-���結G��6w��C��!���=�c��$ߝzCm���,�#����Y@�yC{��_]��N��{�}�'�M�RV0�,���æaRT*J�{߼ɶM��Q���cX�k�َ�a�� �h�t$��p�#A�49߰4:J$�@>�̚H.�H)�����|\����8� T�ʗ��ť�
$���y�m���
�ޓ�F�&B��%
w{����S��aiB�v����5L�A@�*�=��6��Ԃ���w�w@k���y�I}�O_o��De!>��SA���xJ���`D�O|���i�
�YFJ�s�9�pI�&�'>�)�O�u�ƈ��|�ƍ4D�����2i�q�����=�@�%���z�	����e��IjI���<Z΍�:]�8�$�t����Όu�0_�����[������4>��4�(��
����5�HV���R�w��H)�1�Ks_�2��F���~�1�5Q���=ﻣ���	�mv�	nV7�4ѱ�&w�wA�%D#U��{���>���}?E;��wΗM�D�9��4�<;|9�=e��5/=��CMQݔ����J��W�Ud 9�����M^����a��k�c2�FT
����Ѷ���R-:�ߎd����MoѪ�6u��I��~,3�e��^��q+5�{G�j5Q��ȉ��hY�#ȏ|:��~|�	x�<�I ��<��y�i ��}�Ey8����#��	�4�4������#1������A�!Z��`T��}��AM�VR}��'�aq�;�s޲<���;�h�+}�|y[�9ir�F҅9�{��"IA
�c+�;�2:�f���R�S���6�R
CrӮs�d��)
�߽���I�q�o������[+��	�7O@5����E�uS����O�D����ʦ��)�T}T�U�*7�k&����VVJ�s�9�i6�IXV���{�:a�#r�}|���X�	#�Du��,�}�>Dx+7����@�ߟ����\�/g1����H�$xt��'� o���'��T��>��4�p@�D
�%�����U������>3�t;���6���4Bk�f�a/&J�Ѧ���>���n!��
�c+��ј̲VT��W�n�H�c�Je��2��u2�X�N��:����+�tnÞ͋QO�v�*�����A��������PC�|Io����ԅ-3�>9�6n�R����NFJk�F��q�^������C�����%\��Lu��&ěH)�/=�0�c
�RQ=ߞ�&�.{�:y�w��;�,��;߾���'!0��^��˄����{N��I ���tm<	�:}r�g��M� �_em�� �b^��t̲T*J�C���2,�Y�G�O �F-8�}�s�$�Fa�:�5ֹ6n�Sn�K#�j��N�)>q:��N�~���ܱ�K��h�h��s��q*!R�;��2�YP*T����6���������z��!�N��9�4�y
#���Qn��]�E����k "���"�#�#�o非�q�N���ɴ�H,+
����a�F%�*y�=�M�led�����i��'c�����o� 2 ���b,�2�!��J�����q(�!D���h2<	��E ������V��q���<���@�@O_�e֚������{���G��*k�ͬ�^L���G��D�״��4�eJ�8�0@��ea��C���%@���y�g�YG�"��$Vw�@
ͨħ�̛��`>��7`���^������{}>@5aз�ӽ�����|V�§�����v`�1H��FB��jl�H��g����>1�u$�|�t����Si������M�n2VQ��w~�G��N�$�O��|<H�'}�0�Ri
���~�̛d�+%Y�������d �8�߫���W
���Aߍc�����vp�R��X<�j׵�=������z�aߎ/U�\�O��|ƌ������=�s&��h��s߾� Y����.�j�N 0�q�L0��J��*���d�Aa������ܱ�K��8�ƈ��>��������}}����?R�&{�cU� {��M07��Ԃ���y�7�AJy���{:|j���e�)�}���+��݁i]�|�%
P�ƪ&�����W�Th�Dh�����{�K�k;w���y$��T{���L���B�)����h7�?7|f332�q��Ə�����|rw��s�G$(P3�o�7�Q�FSAk�����
�������w����{�y��C�J�C���h�G��&�4mr�y�*�FXi�N��|�m��VJ�×��23�O}����.s��R�S�����A`p�)����r2F!���Qm �썍�ݳ�˷�W�ȹ��,nIL�N~�
��=Y<
�~.�緹��*�k
V^a���U���;���|V�M>�':pʮ��[��x`�aG~���i�vxL�`�t31���K+�ɵ��ub�{9�n��.��4m�z	�.�7��� ��u�.�C���zg��:�W����gl��%���ݎ�t�zwn�cf�m�r�Þ6�o����/�Y���s�M���Vk���/7�z��+`��l���P�H�:�sY���㶗]���U1fÎ�V�0:�3�;8��k$�(�|Fӭ����_����1��1���M'��R
AL��ɴ�B��,aX^c��0�
�]��9��N�����M�n2�Q��������h�?/U�\�M������2G�Hx=&��O�O u�P�aHT�сR��s@m6�R*s��0̲T*J����x�{��{�掴F���F���{��h���＆��AH,=�wё�2VT���x��/��M�s����ĢHk�}܁��A��a��}CA�R��̘��G�D D0G��W�zfT�2�VQ��:��2�ؒ���ay�;�0�#
��RT�~w�M�s��7߽�L2i�����w���7����a�2�2�q(Z=5��%
P�~�Ϩ;C�����d�?{<>��Ͻ���*T
���}C��R
�ݙ�>�>O��W󋆒��V�n[pɚ�Ѷ�٪"�u/Y)�S2�K㝞n�}�[2���i�戙��w@m+����9|�#:d��J�O|�>b��'�h��w�4�H]��@�
P�C���QiB��sp�C�1Lh��'^k���Af�J�m�y�;��
>��^�B��S,Z��3n��i�W�V�0p|7����� ��[�M�Z�P��6�zy�@��+��$�>>^+|ӿ��'Iߚ�y>"M�D��aX_�{�a�%B����}�d�&�Y(�z����_h�7�#�=���@����.DJ��{�D�
! ~��h�!DJ4=�!���k3�vӴ
�����:��J��C�~���%G5�I�4�c��/tq(S����N޾����ϯ�|
U�FKXwy����JʐP)����`,G�#���ﶀ��Tq���ʅ�}�(�MHk�ڷ��U�W�SI=Ϻ�M��
�YFJ���G���6����[=�x�bb�!�XT�
��;�̚d���YY(�C߾��,�)ݣ�.5OﾸώJJ��.���Y5���C�����{���2s↭����mߘf^Z&gǚ��٭�iĢ��w�w�Mn��`V�*]s�y�6G�#�7y�������}������22T,IP����l6°���̹&c�7F�6�=ϻ��!ġk��м��<χ'28�O����>�sh�A`ljB�������HW�[N��+fX�:������7�M|Jݙ�^���]�F��jSU�J���y�i6�V0�Ns�}z|��}u�8���fY9�j>��[�nmu�[�sSn��t�d5���dC��2�N����~;���_�;��J�-{ݟ��a�¤�Oy�~��&�Y(2�Xʚ��@����ym:^�	�44g~����n����=ġJ3hw���[��k��R����h��H,�s~�c�>��Ng]����{��4q�4C]~��N6=a1q�m��<߽���H,�����эW;�M��޷Q�$@�߽���`��H[Ms�y�4�Rd���$o�+���ֻ�Y�@�s�Q��Ì�Q�,	�(sk�Y�N\m��q��W[���~�ׄ�.�~'�W�{|������d��y�2m&Щ+V���(�G���=]	:�� Vͺ����FVKS^s�d�M�k>>���c-�L�h81��n�C��4W~uQs�́�^��M�
Ad=�膡c� |<28�=�+ ���B�����.31Ě��/�����6��*Aa���1�d�*�yGA�Y�}�Yʟ�~|�|(����s l� �HV�߸�R
fk�����1K�NRV{}�G�����>���혌�����ּɴ�B�*Aag{�e�F%B�{�}��L����(�V�}`�8�>�1�/qd��wdŮ��*xq�1�V���+�1�����x�w��j��'���O���YS�w��I����}�N��R��/>:Ǥ��P>;��d��B��;������̖���O���h�"A���7Ρ�d*$�X��w�г�~>�]��/���"�hR�"���ηj�Y��]OmuX8j�$n��D����7*��_~I�k2���u�戞�=��TB5PXyw�P�&YP,J�|�y�i��.���;���Isw@p9

#G�>�-��D�~�{xJ��1�@TГ�����m�����n�{�i���́�;��aXY�7�a�aR
�w�2i�l��2�g{�\9ga��k����\N C{���ave�D��ƃ�=5�%B�H�w���Q�F43���_���y�~���z��>N�H��'o��-(R�R{���Ǝ�Osq6e�-�A?	#�����7���YDp�Q
�FV��P�&c*J�gw�k|�|(�C߾� LvU������k���(���Qn���=�n�cf7fb��8�J����ġk�Tj5Q7�}�J��v}�8���+64F�k��a ��%�s�s�6ɱ���VJ2����6�@ɼj��l�ߺ7��o+�ɺ9�';[��TE�KgL�z�"&3������H��/X����VQ�w�qK��p���UȜ4eG\n�pXz�YGa�&�p:�ͬ�5�>78�7��^�nD��ݞ�pcX��q{V�t�:���:�m��T����L�(�#�n��@�!�;1���Ͷn�vw�5p������v��6��l3P� b۞ݎ�뜧\�-���� 2pj:z�f:�"���Z��^�ᶪZ�{<\�c��-#��ƺ����=�\��#j��W����te.����,1r�>#A�2{�E���-���4�]�H)�{�2��G>�:���?4ng2�J4��}��wG84F��>��&7$�e�$�Z�Y!��
����y��Ó�aֱ(P"D}߾��4�@bQ$7߾��!C!D_���{��k�w|�C|޲�x4&�����e�b^�SI<ϻ�M�m��מ�̛I� � 4F�_�����ϝk�[GZ"K*J'���d�&�2�VVJʛ���7�?7̶̘E/6q(Z<���6���뭒<C����Aߩ
�Z��My��M�T�����| ���!9�RΔ{�@`�" ϻ��6�ƈ�*~�$6e�-˄�ѺaS�=�I6�d�+]��0��wZ�p�G1��bTy߽��cR
AMy�9�77H6��;���a����{�/v��j��9�ŵ"�$��:���k��N�㶶�G<E�;��G`��v�Øg��������)���O��j�Q���{�d�M�A%H,/x߹�
L��^o���}�|���J�5�{�8�)B�pj&�ﻢ�'�vu�\�M�ߊ>����<	����/����R͛Ș}x�=��w�z�BD�aW��D��㔤RySN�Jus�z-�eDOj�f8�r�ys��| �mG� �
���y�4�@��'x��^}@�ȏ@�����/k �&��#�џ>�~	��2�z�m4D�9�4�6�R.���Ι,e@�T�%4���əѧ�iG�"��I�v��(����ϲ�t�D��oo"�]f%�6%}�s�8���ϼ\�?�3+,*u��M�M�aXB{��Ѧ��)PO{���ƫ�_=��ט����d���c*s��ܓi�k���afL���6�p����j�%
<� go�A���﷢]us�;�8����k�l'�-y��(P��ﻣ�h������}�}�V��z֐AH�Zr"����6���5`$�k�bL�t��������,�n\'�bP�7���4��B�7�FY��������bπ�Q�K�!���sQ1i޳�d$����<)�{�d%�ݙ�^��q+=����B����zη�w&�����!�%aXV��s�e�Ib%�;��6ɱ����z�M"G}9~�:i�  `S�l�\�M�����ID�
$�}����F4(S�=�zn����6j_��w���LCL�l�Y���W��h�P�{2L��y2k�n&�9p9@ȷ'ݫ���Pe��>���y����Z�y혗�>��O+�-<�zj�=\H1����~��E�ya;����X�������z�������+�6ټ_YG��d�|���ܘ�p��%��V�[�[i��q���h���\��G������_�^�/���12ӗ�<�^^��{oOI���x�Q
�	n��oM��ۡI�ks���]��{�S5�˂�G�I�R鸻W�cV�
��L���{����g]Kp�ܱƃ�쇼��V��Bcqr��]�P�����Ϲ���Gw��W�bѰ_N���5���%��}x5�����<�U�3��haQ����:�;K�rVN��?.��K�]Ň=��Q��M�n�@�`(�LS�B��/�_�����7�Zr�.޷K�����V�W��	�iH�I�mo�F}����'��uᰓp��Y�s\��R���}}����қءYB�������Q��[�Sh�-�%���kxq�^��|,�Gg"�Ae����v�I��>�ؘ��OwP��D�޳m�:-
ݺ1b�Ew�8%^��{��V��k�tj�/I�Ŝ�����w�#�z���b��?���9�ٽ����~T4�TA[f�
��.Qa�*�IX6�ak`�j��
t�h-���� ITc%eE*,�P�0��Ő���
�$jTB��K )EIh\bZD����5�2��A�@��T`�R�RVB�R�eE�d���0�RF8[kN�Œ-db**+AeF[VT�h�,b
�
�D�*,�j �'L�&�R(�`�V�j
Kl�������F��V����*�1Fʑ%��t-�V�DAm%$Yҭ�I��AQ�؊�$鸡mZ�Q��J�Ԃ�,(��V�Z�,Z�
���R�Z��PX��ĭX��0�L5����>$ w�{י���*e�~7�P�*%B���ɶ�4F���v��Dn�G9M=w�P��_�Y��	�#�����3P(��9�d�m`V�!!���t��=�3������hg>�1�����ڶ_E,��m�6��{���� F�5Q(S~���Į!����^{}�;H,�z�L20�(�ID׾�̛H,�Y+*k�{̓i���?{���7!X�D%��AE*"�b���WrK �.%1��K�Q��z�\�TT�M��m��X>g]G)ih���ɭ��
���Ms�y�6�*y�]�y�2�]����P陃%B�*C�￴q���Wל��d�-��&�ġLy�����Ad�1�=�9�`����I �s�|��`m� ����J�;И�o���~��(ǔ�D�;�|�C2]��^��r�����8�,��YFJ���y�4��T�ÇZ�=Ϸμ�^��t�#
��RQ;߽��l���P�
o�}��L��푑�˄��hs�`}���~����R�֐��u�{�[�+Fl`T�\���N D�h{ϲ�k��Y���g�l�b��k)��6L5�S=n(�ѥP�&C؝cw[��Y;`mF�(ҳu�*�'�BH������< ���>T��y�L6°�<��L�./UcP�AO5���8!��B�Q�����G�}ꭑ�xg��@�g�Y�Q��J!!�{��9
P�0Bw�e頉x��.�[j�{�̋� �V�욡���p;m&�3U/$!�+�7?����E���1��"s�ލ��J��D�9�2��J
����0�¤ٜ�s��v _7�ri�c+%����7�~��qן���̘Ao6q�_�>�rDx</#��a�NG�{��|�&�)
сZ0*]w��M�T��YR�^���J��*��}#� ���|,�#�n"K��MQ�"f��t�P�C�{іe��T����_^�W�׼6�����i�}�st�e!X!;���uMI�}�8�2]��^��m'^k���=�}����;����Yc%L{�o&�&ТJ���/��a��*J!RX�y�~��&3�q�uN�*AM�߻�6&�)s��0Vץ�G�~��}{Bl����C�>�oXd��bH��~=�s&ˊ��_Z=���7w�h�XS롧S���'�➫3� ���_;K�b�V�.�V�hn�B�̫��~����������mzm8۲�\���"�G+�v�A�g��Yٸ������ٸ�����;f��9S�����
p��`��)�]ɱ�g���@������糹٫�C=���/Tv��k�G�q�Cj؝:�6�}v� �V���W<�8]�뎴Oq�M�x_$���������6���۞�.n{Kc��&�,���r)��5��r��u�+�-���݄�3���|��R�1���~d��ȐN��S�7��nF+�q�k����}�D��0#�&	�Ӵ�$����j�[5���$�o`I��`�a>�c�n�z7����.`�0	"%�F�H��/r��>}+��B��\K���}|wn����@�d(�EEל6��Vc$E:��$���l�Iǽ�7:�OFH`�}�>&�i�(L�d��Vs~$�u�eT�cۺM��$q���I�=�l�q�cb�U!�0b�mJf�SF��3��f�n9�ps�5L���qA��P�������W5ƽ�#����̬Es��
������*�x"
�$�
��+�I�ܽl��9�|��H*����	FĽVp��s�b�@�c}���3�Jn]�����Uw�J�he�I~��oYI��������<��5Q��^7�vo������@$�|� ���%E�{0Y�T�k�l�L�`G�L#Y=M��A�ی2Dv�z���Qu��A>&��[$�{)��BR	���#�����V�Ti'"v�I�q�O����������7�Ip��,R:�`ɏ�]���������ӭ4cP3B|H��� ��7`����5՝���U�)H��T�k�8�f�ts]��W)7i� ���A7o�����L&R2HO��5�H�݌3�H���g�r�	��$�u����e�E(� ��$��Uaq����A��2�$M��}Q�l��evM0
s]w��V^�﷭~Q=��b(�۳��O9�,.s\��7�^�]�T�0<!c��VB�*,e�=��z����I�7�#5a���S�[la�S��gKρ>$�������I�ك�(#="a�N�k�1��0��S���$��I$���wbG8!@��7�CJA3>>��驒&�/���幯ȋ���6A�9y>ݻ��3�!F�����x	8�쮊�ꥐ��f�٩�]����q�M��2Nm��E)Vs��^R:�P"���x���>'����������ݾ�z����0��HD�!6#k��gs".����dO��D�Gm�P`��U�9,fU:����PB8��I����`�H9Y�yNj*�����48Ay�$���	ڽ['�A1 ���[��aA�/�����	�f[d�q�g/�?�y�/]~�0��a�K�*wĴOY���D��x�~���ݞ�!��ǂ��윳���v��S6�v��T��.��jymv}#�|O�&3��)="a�����u����C�]�x��A ����$����*�Y��=._u膤�� �M���\��NЯc�U��t[n絉�cS�l-��ފt��o��y���L��m��$���D�IT[��~7]Ewm�'�0�@��AQ��;/��w�2j}�X$�}]{m��H8���p�;�*�8򬤌�PfIO�պ�$u�c�Gr��*��`F�p콶�$�{�O�p���0� �}��Q�evϺ���'*�)��=�l�Iw��qRk<ok�0Hھ]'�A�(���[��F�ȗs��<�p	w��$u��@.�uo.kPw��.
��.���UO�Ԗ�e���{4��'p�8�*�V�e���.�sa`[�+\e�߱S&.��;��ow쿽��v�@n3�0�Zy�ۤ6\e��n��Wp�eۚ[�g�{h7Fy�k�LWlu��82ѻl��ޭ�s��[M���;HvW&k��=��5m�uה�9�3ٝľ�\�`�GCul�l�U���N0p��6�;���5�#t2q��.��/;Y܃�"��,qVڪ��Z��I��7g��S�F;����qa�*v5"E]��M���a��dJ�݃�)="a�u��I���>.�'����q[1{���o��s��50I���K`�ڙ&��	��3��:I8�q�H$}H>��tv���zOL8P((�TD���;/r�'�<�I9s��S%�n$����w� O��IE��\�|�z��A��y�Dc�l�/v$Gm���=��ӭ�i��7�I�5��#�4<Mr�RO^����8+�	��>�n�$^tH$���l�U"2�ز�Q�T��J���YKkF��T.�nf�^�WA	���nT���.���S�*0N[��Đ�g�|Av���*�.�v2��<���	��ك�(#$�0�F�U�_���8����/q�R�������9����txy���gX�����Ȣ�̀�<#-�����m�UH���|$��D�H�o�l���OU>�N/q�C΁Lf|}��>�H7��L�/�q�㺲�$��AݿoZm/]X��ʜ���ٞ�_=��rw|H#{fH �f[`�q�e-�-;s�$��$��*"�2HM�6�[ ���q9"Ыs��7�I���`�s�������{�e�Pf ��%DLDc X�<<�u,\Riz6ڞ'Yr��Mߏ����y��)�9 I$�{L�Fm�S|>��3ƹ���m�U졙�%Ux�kt�M�z�Q���7j��A�;x߈ �_e�����޸�Df��A>3�t�z�w/�����Kk�m�L%3�4u����ל� �Q�K�	*�r@���|2j|==�z���M�ć�����NnEz�s�ۙ���D�4;�Y �71�Āso��{�!��LϏ�k˦����;*��fa{?O����$��O-�4mK���uFd��2������36d��um�I �^�Iy�z:N$�f�)>�u���b�64v-n�Z�R�����;�;V�ׇ=V���1dȉ�Y�2N��6H%�D�5��`wBf�3v�$��{��Vp���fF�=➍CB���L�I>����$��I�� ����v�uV9�̓�H�TP��\���g�|I2�"62��}�����w"Ġ�I�)�k�i����1�V���]`�=[����$���a^���*��cp/r���HԒ#{��K����J<��ruZ6��7�ù���U��
]m�ݩ�~�&��6e�@��@3>>�l��I �g�O�2�n�:���Sw�'���	'î��J�R�g*1�����#������#�@鍝���
t�WI<k��X�ă3%v�A�)H���|��I#/�I ���3z��Zz���o`H����#&`ȟC`FWk�t@�,��u�{���{������S5�/��-��a��D�30B>Y�'Ğ�ܯ2%e�U�"8�/f�-�|H$������a��7d�30��%C`��t��Z
��B��$�Y���I���nX�������3�1�&3"|��ӭ�I's��ݻF-sP�	�I�ȐH%�f6	#;� E�q�7)��ڥ��Y��Ehw���,����5�PL:�������U�Иʏ'kvmDR�ȳ�K��5���5Q]��6��b�Y4,QY�ǟr���������������難��!��v�/k��Os�i�ݞ>�ޚX�W����3�x%Q����w+��-��M9�޼r��L�;�r�c~=Ĳ�~�۵,�����|0$E��1uj4M�	���%�Gl�א�n;����������r��v��Y腈�O{ 揇��f�r��p:�a��~y�d���uX�B��i��ҡ�jy�W٭6�<����'�3�9���PU��1�K�Ϣ�h�Y�ӥ>�vݦ�c�O�-~�B]��~�`͜���{� �M���T����H2��5�o�QH��v���oU<�h�|��V��9������0�^����7�e�f�2��9J��v��~���c�3���9q'F����O
��	����{wHl�g��u�W6'���/�r��`��O����W��\�u��������0����9�Z��$���N��u�����\���C��� z˞���i�v������m��|�{#E����,���l�k�������ad���v޺����1��%�ka��t�f�u�OH6{�x�͍<Ӻ0�
�KS��f*�s7�˜MY�Ӎ��pm��u���6A�&X���
�1�g{�Wy���e����X�TQ5L8)R[Aam�6��KB��[j��X�%����R��lX0aQDV�@+Z1kU�l���@��UZ�b��T)YPKd�(1�PE��QEԵӆa�J��
�
ŋ"�
���P��iFR�
���"�#K$���h��+�1�������J��a*���������*V4*�Ir"$H��e��H�"�B�*X6�H��h��jYVޮ0��U���(�0"(�-�4l��%�0��$j1Pī���%��m��Ս��ь�a��)0�EW%cV��R&@��k."�	�V���+E�X�&-im�(1�6׫)`� ݵ����߫�\jѳ�ђ�Rg&�n�x� ���^fٴq�Oks��e�N����K�&MŮ�!��I^��� r�s��1oF̳v���%Iu�۠�F�c�c� �^f�ɼ��=y��Z�L�\��;k3\{%�hX��Tփ�N�����BB��v�7kl;ȕ�k���mݭ��n�AnU��"�z�k��筬�th��eϷ\S��ۍ��["��A���$�:��1x�(��n݋l���ۃ�q��s�˓�y<X��5��rg��/N1��m�tk���5�n�@�h�����N����x���ll(���;��;l�nmu���zE����)�lT$<��r E�����e���Wpv2���9��p��ve����+;��Nw#uL)��Q�t]sv8���d��s�۬N8zx�ŭ��{��<ei��&tn��e�Ȏ��a�N4VZ��E����۷a�u��t�.�T6Y�½��˨�볷�Ch-��tV���3���I{Vlruu�����YtGf�vG�-�^�v��[��<��k��x��U�V�S�!����q.7l�[�f�瞷�1lK�A�S� 9x�ݙ��;�K1���sڸu�2	�h�9&녞M4�ƃ���;k\s��˧�yθ����$�{L�ۄ��n�)Suv�Z{�۷X��s��'���O<��/7[�7b�s�
N�vw�z�����9��x98��0O����I>)v�vKt�:�!���:@�]�Mڧ�j��n.w��j��E��W=uB����z�D���;�z�.��<c��y8GnyY-m���u��v�T/l�"�3Iuy vkl�lѩ�j�x��>�=��^NƓ�e��Z;v݄ج�ͻS[tku�U8��X��י�K���[����YN�����/j��\m���6�[FW�r�';/�Z��(��Ǖ�.�ݞC��ɋ�vF;n�ݞ�rxj�����<�OS�b�pp����M��n�m��=v���r��)��q\�mnM�u	5��R�scn��b����<#�����֋x�%�#��s��S��.�E�S�R��m{P�.'EmN���V��.ݚ�j�6�%0q�ۢ�6�!kz	�2o�`G)Ϗ�_�l��_ge?I���ɫՙ�w�x��	�o��")FB�R�Q��)������tm8�I =���$��luڅ[[%L���3N�k��3D�����H#{�$�R&yV;��_�n�S�NwfP�8j�AFfG��Wn��o���$�ה�H$}ٍ�I}���z�����ln�b`��LC`�w[�$����&���-U�l	;�(?��E�gv����l(:�b�H�F[f:2�7�m.�H���N�Vڮ�7I`k~��,C�_��2m��I��L�I��F�ȉ��ђ�������7Oz5"���M0F�L���(NB�l�O	���Cn6aJ��P෌e���ؼ�HvJ��Z�z����b�9�'-�^�kBiY����:귶���̯3w�#���Kuݕ��z�<�*,(��u��6���Um��2�p�s���9ݘ��IΥVL#&bQ�Cb2�ZX���T��y|�$m�O���c��gE��09��"k��f�fFfG�6���׻�˙��H�f����j�ݚ߁$��� �O]�7���(�u�%��ؔ�"�LH�����v����;=d���MVے6"�+J��]�j��fI1��v�dG^�|Aw��ͩ�)tx��/��&�[ڀ�z��p�2a	�5ӭ� �/����b�w��N�D��vﱰ	�3ת�M�O;��+��-ㅎe5y�'�Xes����Ъ���P����A:�#����$�g.7Z��v1�Z"y��#$3ސ0�:r�h��e�V�ބ$��*�d��Md�T߄A�;x-/��~�ֺoX,�s2d1Gz�U��&�����*r$�ۻ��}�ى��z�Wm��|w6$5��%)BfR�C~����>w�o,k|n ɠ	��O�n6A9���>��Ж�֯�\~(�W�*$d�����f�o�q��������Vs����;cC�jouV������wf6ͱ�,�x��f�0��ݓ&�3$���Wu�I�ً]��Yn'�w)�I7���d]��=��8��&�2a	P+�:�~'ă���0L���A�}�i��O�5��L��ٔ�ވQ�f|}��"o%QCs/S� �����̊a$<�7}S�K�������A"RшiP���ZII�X�&)�7�L�c����>�]���7�h�k]�\�3��˴8s�ς�sP6��i�p Յ"�j�gLP��_�{e��LD����I$��wl�����Y9��ɋ	!�: D�Yg.H#���t�'Wu�[g�)U�$qP���[���}�]�������ݤ�	j�Ȧ�(�����WH��Uj�S�w�E����a�c�ݪ������^{1` 9�����9s\��� ��ɭ|�����������}��ޗ�]q�ݭ��T���@$�{5Iy$qI;���9���74�0��q w�N�)]&���kT��kJ�[0������(���$Z����]���&I��*�,y�d �&g��Ya������[�^O�/r�n�X�Rk� .�� �﻽���wEҴ�̱�0��'�^�F��=S1al�4يь�^�WS1�/��Y�G9��]���y�n�;���^�Dh�X;_Uz���+�r��Bgh�	���!<:��pZ�I$wd�b��m	��/km ���l9x �x��/:���t/:�u�m��{p%f���wn�vs�n�
2YLc��W���[�����m�����t�V��&��]��Llk�ݾ2����v�
�:z�Z����Z]��quTp�g�����Zk������5���6�.ש{n�t����|�E ����ɹ��D�C��t޲`�v�� ��w{��w��[[��-����/X0��py�y�uڝ�3Z/=��lo��x�.L �z�@ {}�w���/n���W�ë �~sUPc�4=5/fN$�����m"Gnd�,��,}�r� w}�w��x�:����b4�wm5J{��@��A"D��
�{����>��L*�����>���kx�^�zQH[AY4�n{Z��$�\�+�]vf�G�F���I$�{v�$�[��)���,��.�v1(A�;��vb�t��S��v��ME\�bQKRƧ��e�;ނ�D�?���˙��|�{��� ��b�Dw;�3� �Y��v-!�wS��UHj�=�����%r�{��c	q�*Y���ܕ�l(����Yw�D����������{ݾ���:CI�:-ڗ�k���a�nl��1��;s��I-�컰�)oN�PJ&��忚�k��H���HA,	|�{��������`�A��f���}�{&�=�ϐ �}��l`���=�1�c�4<��W~�×^ر�i� �}m�	$�Μ5I$�o�_c�}�̭&��*��Z7Xcd�3 ȐT*a*��
�$kٓ��̾��	e7m�I%�8d��H�����{w�k'gu�`�s��ͣ�}�qF4��1��<�z�M·v�]3~ꇫ�;(Փm��u�%�@ 팠�$�^-�M���:�GA;DQO7_E$�l�C\rCd(R���Y~CSo[l�*�{OH8�O�o��T�I ��Ցt\k뽴���0���Y\5t�k�X`������A=
� I��%�|S�3CsT��h���!צ�E�ǧF杈73n�Q1��T�Ky'rx��V��ut,)������$�Y�f�"J ���H��Ђ�2ϊf;^�57�ޮ�-��$L8�
�D�]u4@$���ˍ�֎�{� <����&�Rƣօ��g�Kw�9Ѹ��uF,1W).�f�$��3@$JY��l�-�w�"i�l�~1�.��am$��H��D��jv����n6<����)��v'UL�?��. Y���$�Hgv�ݥ�d���I�K��� >y�e���nr��Zڲi��뻻H�uW�k�iؚ�%y$����H-�ݻ�1|,sy��[w�6�5<u@��|]=!v�W� �o��u��8I&�K����`�V�d�s��2�G{�]���U�
pf%D�N�G��.��ь���Hnt�$��Y{�ݤI;�:�D��g���ܕ�7�vg�mq�v�ʵ*+�:.��Vp��i�ǉ��V$�!���Ĝʑ�/X�Q7ǂB/�I�ƨ`AJ�g�7�8�m�l$w�	��IvE(�*�B*�I���7m�� wژ��qv��'z���S�g�,d6v�.v�f�E�V�-QYX|2|�eR��o�O:��G�Nn��|�{�{cb�kS'�u�ˁH���"\I��~��[�K�x�kU؝U2�y����/i�q]����$��Kw{n�"R[�(R+�h�P/������E0���7�"R�,.뻶I���t&�IT�L���3krAB�l��(,�ݻ�RD�8�K\r\j�+���H]����/����M�s�H$�Ku�RI$[Ꜫ��8����N�� �{��O��<��J����K�$����s���WI���2��$�	g8�)Qo�i& :�
��7օƔ]X�1[��
2�*�����)�V3/ấ��ң͋��c��2��3i�^T7)�J�7��5�Wc��\�^���j�/�E��	H� �j^w	�o�.�@Ϭ����'����b�֬k�����+�+��M�#��9����t��9�P.8���A�N���v����K.�)��Ik�u/���Wy��U�v�Ӯ9�@5;]�Z�v�˭�=�;0r�6����]�i.���|�X���_�H������v��5���Ij��궴p]O��p�hó��LnYݷ�#�����YNm���E-Nߙ������D���u餒H7�$���h����v�?$O��I6l�3)2�E����T�Uw��b�3l}Z�֒I%����/$�o�i$�tb�Z�s�u�<��S���N��i y�� ��ϰl@-��]���Oo� ��������qKHD�%�C�����?]�bI{A$E�����=ݺ�xm~�x� �T�ɓ�h#PAza�骡Iy%��u����=a��o}�� �}���@�s��w��%�ݜ�75�Gxձ��C�'A��sڍ��s�\b�j�	�rp_�������������֪R��v׀ع��Z���o0A�dϰb>k�s�>8�D�-Nߙ�;v��	]��C�߉�o�a���Fj��>W��;���}�H��ia�h,�|�.��ӵ��6[|_�LZ5 뽣��V�+w��I$1���G;�]�)-�Da�	ط������T�� ���T�k�wwk�I$�o��=�'�uY1֒I�ji$=���ѽ�;Z��GS!�@��B��"��J��!�T�H$��v�ߒA%䷜6���7�,�<$��C�J% 1-�~��H	�}�W�k��2��i��'�2� �﻽������XwuM��w}�W�7��V�VҎ6J�-��:��p],��[�(�U\�|uFJ�c��30 A�����  �=�3�׬�;�eπ����`��* NU+��y:RL�[��u\�H$�B�7n�"R�椚Ks�s���S��^V�<�Y-N_��/;�w`��}0@Iy�c�L�&q1u����L���3�k ��@��oKZ7
Bcd;Zu{��Ɲ���'��6��yt��i�.A�ؽ�'oz{9�-�cw����<�Ȯ�mk�a6�]_���~$#&?��G_����<���k�Q<g�yѮ��ܲ�>C����}����~���/ ��'�i
����|������0{�{{<;Ny����i��K*���Oh1�+k.F�&��ͽڂfBzV7&����'�[Qb�l�ݹպ�A��
	��A:���d���ި6&�k��w�{�9_O�~���y3������}xb.vs���`S&���՚�!Pӥ�
m(zh@u�����i��0uq#�z�Kf�~�)����op���wop�t�Dz�XwD��5Zk��L�ܞ_g�ι��yG�����U$���pSw��"i��x-�qw�*;	U2�j�~ۚux����!�d�}�&|���C�R��T�}�^���i��q��z�l��{K��M�A��v���ðz`���f��n���|9��pS��5�o�>nZ�9�gw�2n<�-�G<�s�u�V��q�Gg3�'
���1戾��b�0G��Q�����Hf����� Gjh��S�������Ҏx�:�ն^��ZY�y7��<����ad\'��}����9�s��=��������qL�#2ڊ"��l�"m�6�PiD��LH��mC$�D1"D�J�RʹKim��ň��*1T��B6�)H��*��Tr��+C�ck+iV��QEE�R��-�rG,��y"HC����e+Ul2DZ�%e��$ɈZR�R��q�"
��""&$UQ2Qw��B1Ŭ�$YU��h�Db����cJ*Ҍed�lAUQX�%IH��V⌨�[h)p
�m���A�������P\2��LR��@[m`��m(�mAQ�mFۄFڅ�+Q%)yv-(�жƑPDzJUQ�-�8��E� ��P�*�,E�Ub������-h",v˟�A%坟m�I���U$ٲ��!)�� ���W^j�����$L��6m"P�樚$}R�3%|�ʭ�Z{F��;_���&CZA���L ����m;��OxOW�vI6�9�X1ֽn2���Ѭ݅[T��6v5<Zq@b{if�nf�MOX;�ܩ���??g��e� 1-��u��@?����p�IuM%��o6�AOk�d�I��I��9.2 ��J!���U
D�6�2����I�sSI�o�h$H��沽�ss��4��E#L�WL� �b�J	}4=Iy$�m����鋎9�}m���ј1 ��e�<�,��'�6��v�n��#Ob��8n[N4��QK� ^8���I/,�ݾ�w�r!�JX	d��-Q�@ػ�[+�����./$�V���ޠ�Hh��)eF�q��k�~
�P�I���xȋ��G��d�Q�B��f 7�{�֘�X�-mEx���Է��pY��=�w��[;�8	��.�@**�|ȩ��^w��d����y���9Q7`ج
�)V��)����D�m�o�Ja� �����l�}��m�[n6h��i��
�RC^��H
̑�AAiHK`�~��I&�dnE�?O}��� �s. {�w{���~���n-��y��:�"�:CF�ۙ^ o~�u��;혫�k��B��Y2M$�ov݋\ځRa*�p��_n�z<����x
���^Iy�v��K�ޑ�U�mdNDa�s~ˀ#�3��%���5��}��iN��4�cc�錈%�u4I$�n�3�"L5����*�Y��aou�0�粷3�=�owg?c֛��i�:v�}�Ӗ�;�/��{G6y����
����+0��H.�FZ�2o�����K��԰����JDZ��>5��%̍����[���KF�X'���9ٮת��ck����v��F�v��O8Vh�	�n�O;P�:���^��pF�8�Dn��6��Xǳ�*E�m���u�X��n��i疒��7�^�gF��g+���O6ƜoPL�-�q����Mvn5Q�xnZ�/ct��/�e��\��� `3m�AQ�8Ky�ٮ|(ږ�K�y��4Y(�{��X �����=� ^�`(��v_Gڷ`�ښ�I#�ێŤ�0F���IJ CZA�z�xj�ʎ�37U׭|$�f���$^S�B�"�Y�/+0��[^���N)�~@jԊ��[>�m�\$�9�F�H%/f�{�*�B֭�$�=����� _{,���2+�4hSj�t���s;�X�]�I$��D�I�>�
�_VOiʼ�K�y��Z^��TPzE�Wf�����mM���76%Y��K�u�wa"L�H�Ey$>ˈ:f��iJ���F�@p@�}T/½tq�,�4�v%���\G�����}~O����s<7�<��s��� ޸����{+{��pfY�|��Y7{wv��H)ΡT���4Y(�z��٘q�n��������[�+?+�����D��^�/�쉑:����T�혼�X�`�;o^�DRDݭ̍Q3v���K�Nl���@�]M$I���;��v=f�sjz4;+�A7�j��)����������A�K7�u ��f�o.�#�p�«���{Z׺u��QQ�[[�� M�U�9�e� ���]�Y�Kn�Iy^u	5�V�2T	�	��ڪK� ��u���:R�K!C���&�HKɒh$�ou�;z6`��xk��;ln�\>�Ua,l%���y�]IԌ=��!]�N�BK��"�~��#"�R� ����'�q{��I'��~��J{v޹@�ykpEg��P�R)$�����6јQ0O��]�m$��O�ԫp��h��2M��Ey(r;��сV�p7�6�F���*b%�!|�H�{{�ݤA)��Ի���+'<}T���F{w�f7�S[�5����efc;�wy�B*U�[�ב:e�]�v��6�f�3�(�_�����I �����[�b�$ʀ�&�KN_#9<�5�h���� ��w{�{@�����Y�����e�'=_��K*�K4�w^������Ǟ�Ω���8��p �s�����{�U��9ͅ�������\���1��������j�]��vL�4D��M5>t�Y=����T��܏����W����Z{����\A�y����:�d��O	8I�o�[i9?i�#��5�A}�� �TՔ��Mm�sD[��C�/y$:�n�I)ޡ%���٫������K��i�gk�ZA$��h����Ŏ��ѓ��KI.�۶M���q�AFj�*b%���S�gqX��Iy(���&�Jrt�y"D�̭W]����+o,�b���\c�Θ��hPrx�����3�.sx_�`�	��^���RjKٻ�،1"
�e�o�'7*f�p��`��#��`������j��Bzo�Y�RBsf� c^�́2;7���o��$�A}z� ﷕��Zgu��ݓm���ڶ�ۍ��s��s!m��a R�%S�%A\HU9]3{��p)mw�f��wZ׾� ��F  ����v�����rgw����� ��`.�~;F�[�dz4�/s0i�Ü�qkfz�u݂����� g����Kzq=Y�kjz����dD$�NP5���l��_r�X�q�s�Y���{� ^�<� W۷K�����b|Sjy����͜�a$ʎ3A$��ʚ�D���v�k���yI�w�yq׈�k��Q�%�Z��UI�]���ZYζ!�ÑuI3m�w�ˈ�{���y�c����������Y�T�8�����ӻ8�d<��p$���Ώ{�ay"��л}����.��Nۮ�>;��k�?��/I�DtF����Q&z�	2TI���x6�RGU�]'��g��c)jq����cv�=��q�ּ�k{vm�l��7;���X�;v���"��s��u�=��]�\nC�䛲m���jwm��y,q����o7U�=��gCɳ��5<duڻyj�F%�v�MPAg[����9��9�a�mTF�KfХA �ҫ^fD<Y���+.n�ƫ�!��Pn:��;*NPc�n���=�?8*�IB��KSʊI$��̚I����I�y&�y��[h��0���\N�WH��ĶO��I�E���8�wY$@$��� �����`sX�o��z'�`%��ghЋ~��F����$�W��ٴ�E�`���A\��		{2My$�{�ٷ�ȈI82LDC����}km@/;א�I���J	/>�g|mmR�٭^^�H�}��x�|��!S��1�{]�R�| a�b����*�I"���$�O���m��8\���v����]G܃E�)�gk�R��s��l����XZ���q���*�f��<��J5x]�0 ;��z���>���"�Sl�b�5`��M$I�ζ̀���ӥ��!�x��.�O{��v�fjW���}����1�ۋ�Yb�d����w[����F�^1P1��9�����p�T�8�]�~��Tf��O����e���7��{� 2w�o Y�yww�d�j�߲�ݾ���<�--�V���m� ��d���]���{ o��7���|b��G�bv�$D��������n<�	]��I$<���UI�e�N�"�xWgt��S�nR~��f�"hX5n��	G�kA$]5J��l��Y�5�	:�׭�a��+xY�q�e���:�|�;�Z�J�=��n�1]5�ێ�n�+n�9�������N_��{��{[ o�>�|@=g��@��D�}��lb9�$a�X�(�-�7�T��|����g6m"in�&�@��	 �=�}CU���y�i.� leLJ��&���&  ]��� ��\�ٗ8������d�YŚ)�j�}A���/�5�2=Hc�����6��$\d^�H��M�����IyTn�&�H�4�h�4�H�KX��O���?@V��< Sx\��{. =�w}�������Na�{#�ځұZhl�U"PJ��]��G��G��Q~I8檒%��&�����~��D����Z׷���*�d#X�rT��P�CX48Ĕ����v���O�nʎ{o�7c��$��|��$�s�&��In�m�1�;�GW�=&�d�LK ���q��7ץa
��l=׷~�Lel��&�j��"�H�ճ4�I.��RP}m�7���y`)8/
n5,�j=i
����b�	/%%�l��:5.XI63�[��������4��j�)PCL�GGz�g5��%��M
H$����۲l$��g�U�F�6f;˔��������6�\T�z���x|��#����hmVp������ڗ���S�Q�q�$�$���h)�����m��~%��2��.u�'��9��H�v�h��l�J�	����e�?Oݵ�;A�F��Lݪ���pMr2�ێlt��(�U^k�=*b-�jG�\��I^��I"kc���5��2@;=RMy"�]�I����3��Jz.�T�K��jzI��D9��D��f���H�lq�H��누�gw�`=�:��|�v���^�}ޞ����a�H$gn�p��&f�f�I<��wnŢ�go�ab�U�%�4+�f��{��/%�$�yn�$�	WF���H�ꕌȸ��9גK��-�1�R��փ�����Ņ\��1l���N��컿$�4�̢J5��dX(��'���S�kUO���	!Z~_�@$��?�'H��ά?�`�����R�`��@��������Zٞ�ԅZ���L�p�j�E��� M��$ HI!'I�	�Gi�H~��,���R�*@�d,���>�0�H����~N�j�_�~�_V}��>ɀ�zO�Q&L�ӡO�c��Πl?�֓�7��Ǧ�)4�w&�a@r`=��s�߀	!?���?���������D�rO� @���&�!HO��,,�?}?����(}����'��3)�����i�Lϸ>S�>��@$��?�C���b}��{���	HC'���%5���H ���Ɇ��렷��ԑ�����C��X1���������L/�$��J@$�Nϫ%�F�^uz4��[0�s! B0a'#Ҭ���2<d�#�j`��̟/I��G��	 B|I��%>ɠ�d�����>�~A>��S����?��,�2XZI�Ϥ��I?���?#�RJ/������*|}�e�H�����3� |���>F���	>����4t�i��t�<�Y����}߉���Ͼ.a�2���}]�����~S_�~��&Ϭ�d$HO�O�dc���~� ���|f����'�@����
2�|�IHF&'�	 B�?��� '������i��:���P�蓿�'fB���'�I��@�A�>�"xLL�I�C�|��HBX2d��6}��5&I���H��Z������	�O bI�K?t�aiM����E����H����}�~��C��HH��@�Q��h�D>��>�'�C����<��?Ğ���O�����'��#�!�����y��~�Ň��1�����~ψv��! B}��>y�ϛ�A�K$�����w��H��O���s�������������^C��>`L"��ߐ7�;�ܑ�������bC�C�>BL���$��ϟh6~R���>�������8x|�����2$&�︓�I�C?�c��#��_��P�Oݰ�}A����}^��aF|�ݫ�vd�RJ��?_��� �$'�B$����	�>p;@���'���w���  I	���~���D�>A�}Ԛ��u)'q������d��"����XC���!=�����ܑN$��Z�