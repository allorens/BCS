BZh91AY&SY*�����_�`q���"� ����bG��                ]��I �B*�$�J��UR
�*PA%�H%B �* ����UQ"Z4�I T)�(    8dT�U(���PI):h
֠JR�5)!QT�����b�RI$Hւ*��
��z}����v��*U�UEUND��3�lZ��H���9h����ʪ�\�U(��r�j��*�kRU)**5��I"�*��V���KuPt5T� )@z����WK��阫S��nmt:w[a��m�{פ��#6UJ;u�����*�5;5u��pp�խ����Fm�v)	BD�%�AT(�})B��;>%^���_}ު�G�����Wm%EUO�U��=�{�P�CkG����
��roT�U�*{��λ���G9wP	J��Ο{ރJ�>��=5zb�T�"Ga��^>��) P�{pR�Ԫ�GOvܟ}�҇�H�Z����{L�*^��_{�*��{������o{��}Wm)*W���tUM�t��{��ĕ{4Ӷ�ڏ�M
�����σ臬��*��b���P��ҒR�����UW���}o�|�R�*��{���"��������^���o��((W����^է��`�>����D}�O��*�j�G�ꪯa��2�Uz��R:jU��h�`BU�}(�( ��Ы�U
"�z_w�U^��jw�C����{ʪ
���O���a��8�b�^q��j]�<��(�T��z��U�k�w� 0�^zE���U*�JJ"�|})E(���*�z������ލ�O UV�ǯ��=��>��'�:t2��x H�1��W@��wt� Ҁ*)Ush�*�*�ϨRR���K�  V����  sw ��{��<���� lw �t��l�O��7�4��T�v����EER�}%J��s� >i�F���W7���=��EP6��: ׽�x� ]��u����]@ �V t������ճQBo|�J � >  �����ˀ���[�M1�� G�� H����s�� 1��^ 
]���RHU��w ]j��} U�| o�@ۏu���-���7Wp q�t@�s׀=������
 sv��� >    �     z j`)RP      O�F$�*�  � L	��)*�� 0�  �� 1%%S�h�4z@ F� I�R&�J��0	��&	�0FT�z��*jB�%=��G�2@4ښ=��~���	?�?��J�9f��`���:�mL���襞?ʾ��삈*����@AW@T�Ȣ���QD�|�O�������AV���|QD|`����E���������7�g����lc�1����c�q�c�1�{y��lg�1�c��c8�1���1��ct�3��c�:q�|li�g�1���3�c�3�cLc�3�c�1���61�|g�1�c���1�g�q��g�c�g�1�n��c�1���4�1�8�1�c8�7�1�g��q�c�;q��1�c�1�`��c�1�n��>1���64��3�c�1��qǎ1�c=�1�c�=�1�1�c8�1��cM���61���1�c��g��q�c�1�61�c�lc8��1ӏ��1��c8�1����q�c�g�1��q�g�q�c��q�g�q�63����{c�c�1�c�g�1�c�1��c�c�c�1�c�q�c�1��c�1���g�q�lc�1���q�c�1�g1�lg��1�c�3��?c8�1�8�3�N<Lg�1�g���0c8�l�7�q�1��T�{d�S�D�D�P�f�P��Q�T�����.2����)�	�
c �*c �=022'��T�D�T��T�P�&P�T��T�D��P�P��T��\`L`�	����!�����!�3 c"cc �*c"c �*c(ccc c(cL��)�����#��c
c(�\aLeLdLeN�SS�T�D�D�����Șʘ��8�8�02&2�2&0&2&2�2�00�0t�Ș��CSS���laaO�������������c"c ��@�P�D�P�1�1�1�1�:d�E�P�������ȘȘ����Ș�8�8����ȘȘ���cc"|`LeLaLeLd`LaeL`o���	�	���c �
cc"c v��!����D�@�T�P��P��@�S����!��������+��3�#������	�)������ �A�Q��q�1�1�>3�������
c"c"cL��������L!���	�!�������)���q�1�1�1�;aLaL`Leq�1�1�1�daeaLdeL`ed`~0��8�22&2&0&0'N<��Ș�8�8��Ș�*c"c
c
cc"c"c*cq��1�1�1�;eLd� � �?S��(�q�q�q�q�e�S�*�&0/��	��c �� ���0)�"8��0	��
�aq�Ld@�:dLd&P1�q�1�1�q�q��V`a`aGS<�T�A��A�q�q�q����(����8¸ʘ�8�=8�G�
��0.20=�8�<dedd\ad`\```~0�¸¸�L�c(��"|ae\a;`eC�P>0�/\eC �A�q�q�Ș���8Ș�=��0��� ʘʘ�8��ȸ�8�?�zg�q�n��1���8�3�c���c�q�gd�1�g�1���g�g�q����q�g�x��q�c�c�1�7M��?�1�g�q���c�q�g1��1�g�q�bc�q�`�1��q�c�1�g�`�q���gǧ�3��g1�g��g�c8�1��=������8�3ۏ3�N<1��q�i�`�q�g�q�g��c8�3�8�3���8�1�g1���&q�g�q�c�q�c�c���3��8�0c��q�g�1�g�q�`��c1�g�1�q���3�c8��q�`��8�1����v�3��1�i�`�{c��8�1�cl��2|q��0c�1�ݱ���1�g�q�1��8�3�����q�c��1�g�q�1�g�c��`�1�1�cg1�1�c��8�Ɍ8Í�`�q��bc1�q����<Rc�1�c��&1�c�1�g�1�c�8��1�c��1�c8�1�c����1�c�1�c�1��c�1���1���1�c8����1�cLc�1�����1�c�3��ǆ1���lc�1�����q�c�1�cc�1�g�1�g�[�`#�R��z�ٟU�yI�^��i�M�Tr��J	�m"r�GB'�#�1�SK3��u��r��xU����l�ɢh^TG�\�9f*JV""Zӱ��MK&�Ԇ�1�)!�.��j���
7@jVҴ�J��'�VG�0�oکلÛ3i�б4.̤��Ni��#;w;:��e����YcH�e�H[ ���{��j�9$��j��'	�E��@�n^���-ڗP`��a�a6��h�)��Q�7f�a����@��s,eXRlM�F�5�t��,؉�P��i��7Qw<Ù���T�P����tm�V�^]eҐ��i��8>r퍲��ב|�bV�.�J��G���j2Sܻ�b⊅fR˒���n�"*!���swFoN�jj�qb7���<1L0+���=�glT4�=�A�=B̤���r���^�&,������9ALsZ�h� m�h����E����)Rcd�[�X-Խu��n�f�h)w�J��ش

%.���f�5�A�^[k]���I�*�n �i��d(���2�
W����7�黔n��=��մ���fc(\:�"�i�V�"�sAn������*VP2�b-����S2�R*�*S̤2ʳ�ĳWt��Y2ΛR��� {�`�K�Ҏ�Mѓ%fV\�ݲ��Vt�N�i�e��t�jB!7�@�EG�>i�(�ih����+.����㑗��7n�gSŲ��:��d �%��M��S,if�!x`6�ÔUͰ(�q/��૊>Q�^��&��&�˦�T e
R���C�̢3�n�6�{����Eyh͛���&�ƅ�1V�(I�[QU��qܖ.�ƥ�[�!�5L�'Nȹt��r�AC3Nk�3h�iM7b�YyQ]�ɖՔ��w��ά�w�4^P�Tt�V�&%�wbmFܥ��U;m�"�׀8�t@ν"�^��Zt��(�w�£���	^�D2=�4ѓĕm
y�%w�ޤȆ�R�Y�X��D�j6�|�i�R�Ϊ{�
���9C[��®�dA�F���<��b������`���������6�����(t$u;��F��O2�m����
��5����@Zێ]^]��m��&f�P�I|��*A\��L�X�� �$������w��4�ư�Z��iMu������	���`@�N�bt0��/�-��h�4�4�a��st�f)Z^5�b�*���n�e���㊵�F�h��e���T&Mz���\D�ɋ���VT��Thc��P�"��Ҋ�3w3Vb��=2���Tf�:*ڦd�ֆL���M���KŻ�qA�V�PI���F�c��ذu+�Ɇ1��٦su�6�FI3vd����Sf[��NQ�J�NV�GB�Z��Y���[�u�X>"|S�j{����9R�m�.�1PD��Sk*f�kn�*l�����t�PEE,E�8�B��WB!��1�����	j�D�R,��o�Z�`8�q�J��3[&J
��twa���d�kZl[��\�����b�%"'Qj銽���,�%�u���M�2�x�G��ĳsp�;��I��z�үke*��r�Y�+lL�w� �WS+h�k0)%�����"��ug�NvƝ�5�P�@B�mІR�Jx6�L�l�h�NX��;d��$�	F�л��/D�o^�x�1(�4��;��U���ʽ�톔up`��r��� ��n@�ɭI�f�G$0on�h��M�ɲ�e̶Z҅��GH�o(�`��P��Z�4|���Ɲ��6�M"�XKCH�K�았��N�v��y�,��\IWv��S2�Q�6-�kopZə.�����N�Q�x&�Mx��ٔ����ˌ�"�w>�.4�w(b�2��۽�(L�sqQ�|��P.�T��s4�6R$�vm-��f�ƫN�-�m̲����ةVSmK�߉�\�)*Э�;n�0�b�9���	�m�9M˒K�DD屭U�&M�v^�Y��Vũ
�b틩��T�ᢶ�a4ʴ3t��N�יH;Ti���Kl��#z�1�Jb��c8��Z���j^1R;u�v�r��*���Q�CR��S�&��ᄲ<<�x�!n���m;È�n��ʸ�����B��-F�7�mX���F�m-�v����E^!'ҋ��0+1;.M�1SC,䛊�a7��c�m����SqW*�mZ�0��j���*ݬ�\��X��)�f�f�jDV���d5N��'3Me�x'�w<vV�26=�n	*�kՇ/.]�ӳWX�-;�t'��v�J@��y#ERt�����3�v鲞������Mk8��E2J���"�GF���f���&P��x漤b1��zK56U#��&����#�{Vf�v7v�*UumT)i,_�V���m:�� -�#��#$�;��r
�PLj�j��H��r���<����;P�yilŀE�6�f��))�Q�Q����f���Q�d��̛F�n��ǣt6aā�Y�^�%�gek9�7���4�Lئ ����K�N8a�4۹.��tQ����\ú��m���)��&U�(���Eeb�mՠ�ke���R
�2�F�-���t��M�Q�{�VX��!�K)9W5(n��n�r�G7J�aD;)Fߢn\��%����2�2�P�t�zM9$˧v�jw���5���(�ӎ��EY�Er]b���	�[{�aJ2<�ঙ���Q]��H#���YzPu�ВƜ1]/��.\��F��2	{{YR��9&IR�B��Jތ0)Fؗ���ˬ�l����ʺ�{�*��f�M�SR�MYr�r+�1	���*e\�7I� �M��[L�ѧH��%	%�Β��������hV��[�L7�mz�5��jdqSh�����2�5��(�[r����$0`>�ز��^T,ֵ������)��*�����hJ�z�Ɉ]�1=�{`�h�Dװmչw3k5�b�����]�ӥ�:�ь�6��!����na����d�脩d/�RZ�ne�3j�^.\f�fR�Y�+d�ӆ�7sX5�*m1Q:>d��Q,�:�h�TG�C��N&�l͎֝�yZ��䙒ն��/ɔe��4�j5�����t�����jB���ߐ�B��)��) ���x���ͭ&AB�vĻgfˤYon�j�[E�M�����:[�Y�^[�%czN���Ӛ�bpͺTYz��r�dt*������N�lE뫺���윌f܌Z�䒀��F�-FC�v%��2RY�Sǂ񕦖ր�ݙT���b�+���21j٩u����I�.��d�n�������Rk�m;�U��my/.�C��b�R�v��j�ԫp�Wr[�Q+l�Y��.��r�Mq�h��{�*��b8�
.&���8��:�2�döDS3Z�#�CA��y9����aꬩ���i/P֪ٔq�5C�x������0^�ĉ�qAjJLN](��(<ao�H]�D&��ͺ���ndÌ�	�h�-\�y��Y[E\��]��y=k��ɐiŖ|��v�ǂ��5�E��є��2�nG���n'2�w�m��# IK��]-	Ze�yt�j[X�F�`�e9�O�$we�y�9+Z.|���84��V4�cMe�,��t6�ʻ:�6�]�qZe7 �=Y�&Z�mcxh�b�@x2�N8(�k/XIx��-
²�WJH��Ҳ�_\%P��#W��a*�:�&"�9SV�O��Cf�
�	�+T�Rr�K�F�?��[g
E70�us���rt:ir�� �F�N�1��ˬ��;̱��h3t��A@��^�m+��x��&�i�ٻT�9SH�R�*Q����/69�b�5+���\�=T��5ZX����r�IA���N�����ݸe��L�%C��e�Y)[6�j��ne<�s�J��G����L��Vk�jGt4�Ɇ,h\7����9�i�{���(8��I�q���0���Ъ@�7��d_Ɋ�)fn��<��@��dʤ��R�m1^�@�R�B̑�ǌ �ڢe��9em�M�����)nЅ���v��Tf�m����`(�q�a�t�=��i[uwB�پ���@%��X�"��p�����֖۠F���f����bْ�S���z�^B��3�GM\��0��PvE]�2.U��0��r�{hf*�2[�5�5f��5o��HV����CM��\[Mn؋I�M���2��U�#E�f�.�e��d+73jf��0��̨��mQd�ܠ����Pfh[��3]���)�e��F�@M�G�F�U�-����z�j�6TV��ǹ�*0U��l�
�X§�yW�����t"4Y1AZ�1Nȫ���7v-!�Bcak��p�p'�%�7�;F�ʼզ��I�F�G^cy����`�-�6�H���J�g���An�H�v,U���2����є�uwr%Pؚq9��Ƶ��`����ɺB�����������)�;0�b�
��4Z͡�8Q`��Y����b��N�L��%ֹR��
��<��hSͲ�r+(EY���Ӻ�z�J*�kp���Ŵ��,P�֨k���1�cߔ�1*uz�����q�d+�ٙ�͊3A-�	PR�qX��1�,P�o1�����q����6Jʊ��mjVN]{F�EF�P�p],کK�m�d�Kć����1�3BE�f"�n�=���p�&��.��n��a�a���:>e㸲�YnE�xU��눺D8)��tӝ���	5ӮнDX��=�b�y�򕊍�ŁU�j���v`�R\�Đ��:��#!f�a�WeܰT)��v��˷a�Gj���N=d���ǫF<��Dƕ�vB@]���~*��m�<��ҬbPI �����z���P��U�"`��`E�la�5��F�)H���#E^����<m���"��u�^R�bI�bOu�g5�LxW�̅l�\-�	ÓS.e�C�E� �ڰ�uB�5��-l�䱤��������[YN`��$�a�D]H���F�톬ռ�["#$(��N�zN*m0���Ɏ}�KB9B�5�+�V��6�Z-�:u���<Z��wYXi�ԞX�b��(��,eUȑd��-�2��j�i��1�(�˳����9H������Ǝ>�4�ݸl^7���T�>w�rv�a%��3+&�D�z�o
�v;��P8K*�Üy�≴g	��M�ހ��d��w��,�+N��|��l���x�g0��C��&���]�$��8OC/o$F"XT=�i4/	��W���x��	L;����P6c)ӼB8^�0��똌Fq�3Lަ�����wY݋���N>㌸R(�r��l�sx���8���;���K{i��еP�q�".�^�f"������]�7���=��t��u6X:���&�e���t�x)���#y��������{�w��G�h�cy�AR��^�G��#�%���]�y|f7hZ䜷��.���ٕ*䓚䝺�A��i���K�����}{���7���6��7$���I��+��l��ԨI�G@q�ϥ��Ő�2e�eoӥ�+��Nk��K�p�59�p9Tb��,=��V����ӳ��":�9ː8>m`
�{��/�+u>���V�\��͜}��Zt�(�wnKt�L-�Y�LӫR�:�Yt������b2}!S������Qy�>��.[O���;4����7d��������S�SH�N�K.E���p�&��v,���oe��4�ڃ/��3�l{;;��x�$���ol��8�r�f�J킬��rv)gVŚyN[;�NF��Ɗ%�kN��d<�od����
�\:I��]J�q�L7��-Cxa;�wD��)h��7�Ф<��9��7�t@J�e�A����ƫ8�B��^Ǚ�ػt2�Vh[e�(6Ƞa:u��|�����0��MJt*����ޝ'4�����-�D��"��P2%a<N��3�s�',�9CQ�Z��`�r'(Y2%Y�"*���6q�C5J��R8S*�u.
��&�˛'s)�>��d�1�z�8z��1���(-���1dq�o�P�)Ґ�7���uX���}Vn��[��,�$2���q�W��hf�B*�>ہ�϶^�Szv�g($aW"$��]ox�;�i�8���tKlP��L3w�pB��wq�c7��*�%i�nͲ��s�ǘ-���o/���Y��wA���%�(]K��v~�1e�BdL��ӕ)�_yٜ�^[����@<��Т_?}�aA/J�l�8��?�tH��,�6�C��Fɸq�e���4�=���YZO#6nMDB�Du�eжm�@#��Q*�Dq��;��n��+'�a�!��!,�Y$�CI�:ΩX�(�G3)� Hc��9eC��/��˝g�P���+	��U�f^�wd��S1�H;�2c��&IXR;g�Nμ�%�C�E�&q����	�z��a�A�=�a��ͧȻ9٩��C�#���]�g4�+��/OPp�V���e��FBY�r���͜z��W{$�}M���ޖsI��]��Id�P��C��)�Pt2�))}�P��x�I2A�4w��@�"����=A���2��
�Ì�8����"$��f�՘��p�B'�tNa�{�;�h$�s��#M��:q�2�c+����a�E��:.U��ð�#8s��[k.����d��"�����K=�������x�$�ʡd�N"Q��^��O�ih�GN�ܭ��r��Zݜ���r�di�x��Ȼ_\_��6Igt�ws��9CI�E����L��]I�(u�����p"h'-Ҵ�Ww�C�2����$�(i#
[��g4�9�0�|�}s�.�O4���2?/�a�"{� ��8�{o�[:�~W���{y����0K��9x`�]��-���o�iTs�L��+�9Y�8�P4���wY�_�Z*Q�jd;:R��x;{��	]v�o�CA�%B
����Ù�GZ������cܒ�Q��Vj�tn��+��#�� '��Σ;-\<�q��$�DsV�w�������z绷��F�̑�82&��]jd͂�q��^��3�j0��#]��b��1h�8������UE���*!i�������l�l]t�&>yZx<��	IX��N��3,)��5���5ݷ� �EfKZ=h���R�i�w�	z*p=���X.H�O�d��=�f�|6E�8��v��4龾��d���T�Z��f�[㫳�qŖ�wݶ�+IRst!ӹp�ҴXg7�@�%����L�kwd=|n�d�<n����� �8���l�ʥ9J�Aq�Uޗj���3F�aw���s�=���<�JaEH-+R+9�[�>���p����9�5�j�VTH�x6�)/�_q�1^}�˹���VX��]k,]\��ՠ՞���2��OmE�q�+t��S��5��>HХ�bU�pu����t�Z���p	/=43��Q0*v2e�b�ѵ��Ȯw��h�O9��#"�*R5�n<�t��9.�B�%Cr���7��{v����݉��{�:,���R�-�
G(̶�M�[�L�w6�۩d���Rًp�E�b�A��jl��2���OX'���ɮ�Ϊ�o$=��QB���I�4J���3T�I���>ޠm;CL9t��<�7���NN���t��D��!ݵrWb��d�.�VM�q�.Z���/q�7�ۼ��f�&Q��G,ۙ,d��Ӻ��k+�%��</!ٔ�c)	)&�0���6ź���	��6$MV�vʚ����l��H�nw�^��*��f�;��;e�wyjv�Q=�+��GG	%�:&Ma�l�Ɲn����U���}�=��'`X���ȥQ����0�Btk��f�}��:{uw��4T4���ev�[��M��G�j ���.��t-�w�ݣ=��B�gq�~�$����n?�n�ntr_LF�]�U����M�4�:��ڜ�����1�ڗ©T�ᅉ9l�<5J�1v��X,t&�j="�8���G~��Ԗ��fm��Q��Wq���[U۝s��	�����{A��@eb���u��ڝ+gY/�"�&���&���	��ʹ�>
�ө�P�u��6�=}�v�fWL`���=�G��̭���ڮg+(��L�\��]n��Hu*��Y�N���_�33��K�˻�3[<�=vG�f	2�u����эV=��;#�[�o5_�n�T��5N�ٰ������u�L�	�[9|�ά��M�����os� �>�Ofw=|��[YO.-�Wp��읾��*"]�"t�8J�m�u5�)��w�cy�X���:�����.����6�\��x��=g��RŚ��CG���b��]��R�gj�˖b��i*��.�B���?J}Av�0�]ٚ��[RU��I�OM��vv�ԥf�K���44� E��&��'e�7��1�e΀�^�Kwzm�/:��:�4��=0R@�Ś2�`�M�:�nۈ6�[e1eݔ�K�)>t���\.�o�ב"�bKR�vP��a֫DpT��;�Eܽܕ#]}���8]X��>Bc�I\�Q*N-��v�oQ� �up����r�
�<�e����۝����\}Ӳ����#r{olw�%3n��*�9a��V۬�4�p�{���n��b�R5Z�{@�B�8��P�j�e�.i���ٛr�y�m������f�=Լz%d]n��s���v�X�G��0"�]sK0�s�i35br��m7�u���hc�,�������v�Xq`p�tU�,�m챣�0�ྀQ�K�
�ɷ}���U���wH�ǖҾم�D�M(j�)oU
֥��P��]|�.L)��f���Ulf�_\:C�(<�F>�vF5� �Tj1P�f�3X����&n��%���& q���$=\�Fd��ޙ��2�_p�c��غ�z9.��X��9_d�7&�����ܜ#��)�st��J���,� ��:E}N�:��p'Y����d�L
���RWgmn]�2���v;����"M�8���T��V�|�<wuKi��w\r�5W�;/N�R;�m	s�/p�U�D���ڲ[�7�lMwAl�XEI�#%kP⭮�������@��%�J��:��ҜM��u&��n���i����	c�7y�ݎa�(s�aë)�R�H��ͺ g]��K�c��8_u@�gz9��M���+t�al1Y�_�25ښ��(V9�e[��+a���8tp��--� |6M�+&��|V�!�7b�������h;�f';��(̖�r���U����ff���x�Vm.v_�sV�fTjSN	磊��[����P'XR�nH6��7v܁%�+2�ʱ�V�NںƦɂ�R�ڋ^���iҀp&�I+�ہ��)czP��i�Ž�.�XvA��̛ƻK�g�����{��aGl��-Z��D���w}Ɏ�yWOM
"lʵ���+��<�k��Wu[�I�:9f�zq˫�_bX�W�+$U�����L=#��ϵfc�a�/'iU�+�ڒ�+��<��Ǜ�H��q��Ju�rU��8c-f`�}�=�b(O)tj|�U��4���qKS�)R�6��w:'�����fE��:ڜ�A�`,�dv�S�Wj���\�{x�%��t;Wl��ep;�Q��>��P��ʹ0nuqѲ�:H�|	�m��dgo��ȏ�8���z/��50��}�wp�]@j�=��Y)��;�ͣOL�F�-Xx�4e�9�ei4�ͳ��m%V&G�hm��������t��)*#VWW��[ht�� �6��s��.ޫg]൭Yml*t7A�:D	N�sDG����d��)�a�bXip��`o�oV� Mf��!Z��^�`A�)f�$�讹٬e�6mg&�+f��y��;�Z;Q{o��Z�Oc`ꌌ��R��Z���H;3vԗ��_ t���(�GB��\��F����w7ڞ:;K���gpi'����Y
��iv��Ok/�t���Z��]��Ϻm�&�Q%�6Nn
L�|+Owf�1�̷�N
P���Z�Tغ�{kU�Y�Z���	Nn9`��L��7�ά�PR�ˑ����*�m
��L��S<fl��\���F�]����f�d�tU���Ɏ�R�Z��Ã.m<9���b�wm�OO&���O���6g:�����A��/+>&^.�9��#V�]�]E������er�i��o��t�;�;5u�g`]ՙAZkA�X���.p�d����B1:<4L�V���b]v�v�I�p�+����O"����4�T�3g�ەF��/�]YoDi7�K5�/�t�;�k>�˳��I>��;�R���XҚ���}w	��W�-�q6�v��nWSi6nu��q榤&w+[�t��VN�t��\=��S�y��k<-u��Pr�s9ӫhX�.���v+e��3zh��y��$[kE�*�W��$��M-7���p����{�\.��c��q�/����(�d���]{�J�\j'��'MŽ������iV��&�6��n>u�O"J�c����v�C�̛�qeɧ3{yk�)0o:����r���ؑ�_ m�2]ՠjZ��j��{���7��'u�WX�P�\:eF�-���t�A��*�*����72^k�w��g��=ľ�b�J�zr�y��|�f��!���W�1�a�#哐�[�-ڳ;��.ƙb(�P�r�C�%���]��bL4F�'0��+8���4��:��҆�:��,e5|�m���4r@c��,��$�]jB�k�s0�˴w.�9ܸ���-����]Rj4�f;H���+;%h����4�W\�m�	�+�yF�ObV�f=����V_Y�G������J(�Q�"�����w�(�R���w�gW6�v3INe�Dx�4g	6�5�tp�-aL�kV�E�r�rIN󹑭X���N���̏�̨8��&qLi�7x�ÝөO/z�L�˪ �Zs���+D�Oz�M��X:)��Sp�[�H@^��\��2�Us�\��4 [��P��#ҍۡ�N�!Cf��q��M��o��^,ftWƹ �6��6��5�3��]�$�:,]�𭩪J��6�`9�0�j�93��	���71	h�𠮖�kEm���rZ�7qbo]K�ҭ�J�k�����<�2D�\s�{�7�ϝ���[��װ���)G�`8����"b
�@�r.�x��K�S��������1w,���������V��z����a��E���_jd�o;y5ك&�.��z�˕��Xi���d����<Pc{�C��;nz��%����.*�Z�ڊ��D�!���*$�>����l@�v����9{���3��i<X8�(h���ҳt����8(�{�bwvX;�"Dl$JJfYT`�ݎ���$�1 س5��"�6�ݜ�mZ�4 ���-�sV�z�!B��{9.z�8v*�l�WK o_(hγ:�x�ͥ�U�W>yg)�7�oQ�0���Z��\�75oһ�����	
;��كav�����Vo]�U�#IW(�l��R�ʽ�#Y7�މ@��Wз�ܜ�{�[.Dm�S{�2�<�{���b���r�;z��]K�rj΀�	Ι�7V�7����ܛ�Q�1���u�p7\T���['<��S첕7u���e�s�����P%�4n���3���9���Zo;8�=�
�[���a&��'|�o<�m���{Jĵ(zvb�5K��S7�ͥJ�̲P�m��ú�Bӛ}�RF�zo���:�>8���o[��L4'qނ�`�h��]�{��t_�bٜ�-\s�:�n>�^[�D<��������|�Ȼ8ugp�>t��gu6e��^��K̝zD���i�kF����;hò���>�z�S���fC3�B�ޜyԸb㝇]��.L�r�Y��t���̡�KcJ�W]+�*��r��qp�c���;i^������R�ɴ�na],�ϵ�������g^e�O��3��德ݎ�s����S������/аx&�C�ޡf�͐
�:;�#D�޵�Ψ|	�ˡ�pJ>=�I��WN׬uC��ޜi�^��seK���I���C�f�(�cM��ӹ>�T#����r.][mۅ�P��ܜ���X�\5��t�w�8��
βgu����8��� ��"H  ˰חn��¦"j,풩!�H���
Wn;�� ƥ�.�>611.X���`ڠ��CT�D)Zd�,�e�2c�@�KLMhBD�Ku@��>0"NJ4�H�T���
s0����H�h����8g#���dN��_,�u���ܘ :SD�@�Wz���,�.�BJ Y�2l���Z�V�I�ϟ_7��d?������:�N����x�������� l����c�>P�ȿ��/I��Y~{�?��I+W9#��@Z2 Ä�{dx�(K��9�~@��|�ړ �y)�._o9��p{� �y	��r� ��g�r<���|�� ��$>'�}����?�N��,��;��D)T��!���D@�^M�� Y�> 4�&}hDD�ʆ�H��%>��K�& �o͝Ǧܾ��"q�R�u;fd�D��&L\ެ��,���$�]��ܠR�H� 0��{��,F{h���I�m�UW3��l��:5���Y�½^�SH4%7C��mT��!ҫaG��)R��#'۷�Xj
�pz�Z:�Nѳs� �I@���)2\@&�I���ߞo	�/�{�u�yJ��	 k�҈�uf
f�@�� 
A	d��)O<�T3+:�?�$HI����?�B��)�������X)������������w����#�:H���?c�܉��٨:�p�F�wKy�o%�\�F+]���r_�0�.����r�=���r��u�x�{�;[�u�\M�KOf�"}F��S%#�6&���.��
tL�p��/����wKS�{ɢ���aP����|�TGk(H�
X*&zX�U{F��,�֯f�ּ���D���MX�Y:�ī��{�kz �~�Ua���3�lgk5����]Ɯ��6�֒暗�qØ�+|o��2Uq��h����=ʹJ�*^b��MM;X��ܭ���pS�c�j���t�8�����uh�<YUZ�u�yx-`
ё��r�p��Wo�0����1s��1�������.W_.��[�i�9B+��c�k/NO�}{gf6�ܜz[��b��L�2ۤz��O�T(fd���q8�t.���֣�]���lP��B��� }��J+oK�p2��y-]]�T�Б�qZ��*u���u+�8��;ej����r�+�NYaN�K�kSP5ZroLכ��E�!�ݕ�uJ�Lf�nr�s&v-�8kom�6f: m� �L�{/ιi���JN�&:o5w����r�W"�]�s��{���zy����]{u�u�]u�]|tu�]u�]u�G]u�]u�뮼u�]u�\u�_����뮺�뮺�Ӯ��n���]u�]u�뮼u�]u�_���뮺��\u���Ӯ�뮺��κ��]u�]q��]u�]u��u�]z||||z||||u��]u׷]g]u�]~�������ۯ�㮾:�w�����{���pk���1�W*':�ҭ43e;����{Wơ�Q�k*/W�U��og���g���ki%�����ǻW�g8���#9�Jǵ�I`J�K��oq�h��:s	��]���!�];�z�Bo����dR$S�5�����u�sv����	��i�;����d� T�XJ�eJ�����rQe�ޡ�Y�Fx*{�h��A%!{�%j���}�kR��X7p�w�u��_YT��^;&��C��wV��D3e*���[Y[��~�6�;�*��u�L-ݓ��L�w+�х�*��Fos�3T�g�\X��%,�<�[V�$�e#uU�ν����Rf��{��k���ccq*��A��ҋ:^�W[��j<"��邥��y�0(p���P��?j9���{�\��6��t���Rؼ�]��Z+�.v��үz��r�Z6$'3�bW�Wؙ��FE��" a�!͚<���f����0�:����.e�&�6ڠ3N�^5���3�0�L�ʌ}�'>��!V�z���s
���l���r�ת�@|��������/�)�@�����\s3%� Y��>��A�5��7��b��R̍q ��@UUT�L:�X��o�ڠ�fې�J>�>O&h���e
b���x�>#n�����9"� �֪+lpV��&��0&ҹ�<��K�� �87:�|uǷ��㮽����]u�]q�Y�]u�]u���]u�]u�]u�]u�]|u�u�u�㮺뮽�뮽:뮺�뮺�ۮ����]u�\u�u�]u�]u�u�^:뮺믏��<u�]zu�]u��]x뮺뮺�κ뮾>8��������^�u�^�u�u�]u��^���ޝu�κ뮺뎺���ε�ub#���L�}l��(��0i>���Ã��W]�A�]����Ҳ�QBH�	����O2c���m�v�/��\=� �1��<��+-��8Y]A���3�	�����4Q�^K��gz�� E+��Ҋ���`�o��[}_>Ǘ.+��-�.����h�FC��!�v˕=^��@n�HU*���,b�U{|�{FE����#^�D3�a�d��Wt�|��ځno{��tj��6e��Q���6}��-����S8�Շz� #�s�dU�+7�Ƒ`ՠu&j���߾���)"c���Q����oF]��m/��y��O'r}k)��a݊Pk�w��u�pگ�_�����(��1L��f�@m�#VI��|�1�dbJ��|�UU@�c��B ǮL�˹ỮX Цj��l�\�������{�w\��]/��~��#!�(�eۛ��Uy�hmZ��wwb6`o�P��{Զf�*��+/�:�{'�R���`F1 ��w�װb�U@Qz�-�v�5A���U2�de�75r�Vh�B��Jo ��n�Uvp�P:�r���$�[�����!�o`��e��SkJ�u��yշ����3�;����'��:��mL�M�¥պ����'�n-RW:ݹBp��*�Pἠ�Õ˟s�⏅�S\�v<]�yVF�����䫺�]lї���C���=9;n�4�z��ΫƬ�#�r���$�[wݗ}���{���8���]u�^�u�]{tu�_��뮺㮺��]u�]~��:뮺뮾:::뮺��:뮺뮿]u㮺뮽�뮽:뮺�뮺�ۮ����]u�]~������]u�\u�]u��]u�u�]~:뮺뎎�뮾>>>>�����뎺���]x뮺믎�����>8�뮺뮺�u��:��y�]��:��~���n�ob�b��{���u��9e��c�����[ť܈��>�,�}�%q�"U�)IS�Y��@��`�z����;�̈́J(�xmf�};�J2���ۈȸn�U�mzVsrN�Omǽ�u/�L�+7��u�}u��js���.����i���L_](w�bb��+��uy{�è>���~�s�^��j���9�E9�s�R�S-�0�g��	dv�����6�7"�g��D[�G5gGƠ�Kq���E]*QZ$���9��N�A�=�*�K�9V\��r��T��W��{G�Ȗű�nfw��W\ز=W}��N�bkC�9�C���w_.�+9���fN�MGF��T�J�Np:���ҹz�^jw)+U�ng=$�/Riz�Q�}��A$QO;'hB��+���[]Ĳ�U�9������I�-��l�E!��b�.�E�.�m-���&(U����ٙ:��ur��c|t�֗۰�IW{�Y�qj�jt[���n�X%�+��ݝJ���ǃ�v�KdWtcAA
�����ָ��[��� 7]�UW�ͅծK�=ޞ�_����{��u�]u�u�㮺�N�뮽�뮿u�뮼q�]x뮺뮿]u�]u�G]u�]u�_g]u�]u�뮼u�]u׷]uק]u�^�u�]u�u�]u��]uױ��]u�]u��u�_��뮺�x뮺��|~�>3��㮺�㮼u�]u��]u�׷����u�u�]�{���o����c;i�:��m��7�&����m�5�W��w�\c��F�
`թ���ͬ鮶�J흲�cք�����w9G���y\�Mh���@�d�\�s�N�ܽ���F��k�z�F��;��r4'H����v�+�QP�`��`E	��s4K(t�.$6捝h�D2>����l�P�Z�4(�A���]$��V�fȴH	.�*���)uh��t�a��s���v[���<��ut��	]�� 2Li�,�y��D�j��vtҝ��ohfn�����Y{$�>ɝ&VK��	�Ŋ���]����b�u��tCv�WkS�C�1C�t �yv��A�HH��G�zR��5�]���yMT���I$d�+[;�v�`x�t��-)�a���\�Ѩm\4Rį'N��T@n��R�v���v�c�o<9_����C=��-�YVZ\^�kl����b�B׬N�`�k�ܣv�=|��Ɍ��s��YY��s�i�rs��v��\��{8�)u�{0���s^�v�Sn�<8^ӻ�37���}a�lg��������>:�뮺뮺�u׎�뮺뎺���]uק]u�^�u�]zu�]{tu�]u�]u�u�]u�_���뮸뮾:κ뮺��]x뮺�n��N��뮺�뮺�:�:뮺뮺�:뮺�ۮ��Ӯ���]|||q�����㮺:믌뮺�Ӯ�������ۯ�u׎�뮺���i!��L�y3.���h�]�{B�p�v�1��2�v�����;N@��`bX������\�=ށ��W3�TǨ�8p\�Wn�U�]
�W:Ӿ5� �oqp��"N� p����-ɿ�`�r�'FY��.Xk�B���$���a�|{%�s.6F�y���F��
5}
�*Ӯ�a�w.z���nfg<M�TCqGI�݂�L���h;�-�9��n��E���N\����WG*�ʛW7yۮSP�����:ؾ哣�t�y����vk3a��*�
]aE,Y�rI��w$��-���9�v�R=(uZ�!D����{l����k��2��
�OxGM�f���hQ�\�&t�n'��I����u]����`KG�n �}P}�U�l�Ϙ_��;��S\���+3�Y�U�\/���:"3{��ժ��Y,˂��'
����с8dR�ӏ�Fʕ�#�q�k��Q��f�j|g��ϲG�J�s>�j�U�ˤ�+��=Q:��t�F�{�mpt�5�9�qƖ��ݗZj���^][y�����=��}|u�룮�뮺믎���뮺���^:뮺�:��]u�]{u�]zt~:뮺뎺��]u�]u��뮺뮺��뮺�뮺�뮾:�:��G]u�]u�뮼u׎�뮺����]u�]q�]~:뮿u����������뮺뎎�뮺�κ������ۯק]{����{���w�ݽV�a\�^q�̑����1G����9�E����p��#��;7m�$5|�ї�[C]5���c+]5v,)݇�t�zχ�r^e�T:�U�0�Y��Z��eM��Շwk��Yt�ٹn�e\��V�w�}���G�};��kfu�EpR*�f�A[��x��E�V�ee�r':�z�jv�y���v�.tr�a�/)S;K�#��Гɦr����9���&Uc�(��}nC:�8�@r�d�\.a��ofV˴�tU�!G\fp�����6��y�-���r��]�E1	�i�� �^&o&Q4:���F����J'��d>�&L�&���4mN#����+�ڥYЀ�`�+��m�ͦ⹗b��ei�ٕ��-y�=���l̢N�M�)�v�O���� Cq9�wq�v��7U�0��Is.�l�t�6ߝh3�v_R}��Ҫ�ۛ����ƺ�k7}h q���(����-FK�+y�Ճ�R��f�[wȡ�M�� m(lr�D��v��\u������ �m��'$�B�,���+�|�]���.�R��������]N1�]Tymono�݇�&��;%���m4�n|u�q���\��,�[ʍY��j��Ό4�M=��ݛ��h[���f�CeG��؇��[�M�Y�<x�.�s2��/)�E���u��ut���C5|���-Z�Иz�z�4�=�6���D��e�l�̪��y��[�&wq�"xU{�Uxڗ'cvZ)65�u[�Q�B��"���Ok��V�&����=
ا��&k�%,׼��P2��֨b�7`=�s-�^q��l��D���y]�3˖�n*T�1e�2P{�;y�A�_������ܻ{���ܧD�b���J��w���B�:�R�%[Gw9�{�lF��X��e�y��{�O��f���鸞����.�ӎd�^��d<;�d���1#{�lgVs�ڭ"�ֱ��5�z�����u��o4pP�����:��s1T�,7�t�6�.�m�f��y�o�>=����^e���=$3:u�r��*���9�e�4-����m`�{E��_%�Qeh��h�Tk��n��,96N��ٔ*M:\yj���O#cxwi���t�Ǚ\���%��-���K�q��ׅ��*ժZ�3�b������;���=u���β��ͪ�L^�Ր��z�(9;q�l��b��܍�vT����d`�����8�)�+}˩B._8�)+F�V%ؑ�����S�S��r|����v������a]��|9n��VU�K1=x���\WAc)ƕ�c��өj��������b��X���Ƅ�{Nmd��#y&�.�{I:-#�Y�sB��l�OFz�)�slIK3K����>;2K�����Oz���I��;\t��{ë�Qi�Ю�<M�N�Y9��v��d9+8�{=�v�no:�#��@�K-��C�>���h�;�U�
�z�gv�GP�ք�k�2��{ka�:�Z�����t�*B��96����7ft̺�Q `��UN�X呼�9)f�����Y�wV���-T�ZFM�VesR]Ήe����$V��uN��)�
�J�^��q��@V�OM���,A����#dG��+1P���-t��'�g��8umVPk�٩^�Η�[V��M�N��i�\̼w�O�;�;��N��f#�W�V�&��Nd��.����Gbb-�6v�����9LT�3�iVsc�|��&�`crĿ�"c ���a����\|���\���N�$/�v��ydͬ
��,���߈Ʌ ���svg6�h��Wz���L�&��*���U����0ϸք��}�I}4�?\	�@X��}�� ��]h��k��f4r�]�n�G��ܥ�Ŵ�~]��#x��%u���aފ�>������Me��b�A����.�������&��:��7���9[+-^�F��k���bnd��p�r� dT7��O/jK�ʋgSo�7���i�����]h.ѽ%�G	S����W�ݭ�sy'+�2���'p,89��k��2��̄��YM�F�gz��O]�P
X���Y6�4��9r�e����xfj� ��ڧRc�/���5�32������"�oJ�m\��%���v�ev_b�Į��U9����Y\�_fWu�&�*9gb��3��cT�-�pWV�r\�ݷ:L��0��Z ����mU�i_]Go;�&ST�X�
�HJ�6�K���*��]�%S�`VL�}�KtSɭ����z�?����""#�����?��?����  �#��?�H�?�?��LL�7�����wy���7�f纝�we��v�x��ܴ;V��S=L��\�!�e̦�
\�ܶ�j���p�6s��/^ֵ\rH�e$W�����WP��7|o�q�v��qz�T�6�^R����˫���u֘�p�?�ݹW>n���k��c�����y/\���eR�ڳ��wc	�W�ź�7]����n���+���KL���铵����Zs��{���Gw���.�{�5�c����T��s�i�n�W7\<��n�k��6�z��C����V��6��-+e�Z&�ޫ�sopڸ{�ۄɚ�l]Vs����FT�D���l�	L�*eH�P&�+�z�̭�nS�nM�p$���l�=j�vF�u��][+�(��fو*�+��iq��/��!<=�5c�����2&�NHc�214:Iг�[ct��%�s��2bu3�a�i���Y���b�3��"�4N�I���Eӝ$��s��+�u%�@UY3A��m���#(;�5ʷ@UnD��q���Z�Bg�8�Y��u�@��s��@�D�ﻑ�G�G�jn�m��-hb̫���Kv���fH�e�),��}Ћ�gwL�%tͱwY��E�nQ�y����1�gZ9C<h�餻oh��R����x�W:h�.�|��j<����"��g��֞y��y�P;\է�7p�����S�N��1й�pg]�؜���}�k� �[)��us��[��T��q����uc�4�3��R]Sf�s�������1�q�7*hm��y�r��%�F4�� 9*M���ևgH���!�t�e� ����/�9%�����4g���s�t�+�M���ٖ�z_;�ۛ�Uj�/��\9�����^�Q����#����d��H�"CRd(e��6�9rE�̖�s{P�j/�/q�JdS$󙚒�L�.D��[L�-����\���弪�6�앸;������j4�ni�L�~�q���m(�g[z㇇d{�K���ʜ�v��j�^�KT��{����~v�+N��t�^r�h�qy�iݫ˺�W���׊׭{�.��=���5�R��f����h��p��sKUtݬnG��v�wwu��W�^Ì�/\��A4�-�S �a'-I�$Ԫ����[��7;���vM�׌��.�C��U��y\�u9���No��9^�η��vi4T����*H)S� ���3%�|��nw�\�;Gt�tܷ�^��Ҽb����W�P�җ��v����r[N���m�z�㏉�A%D��E�L�AL�����װ����/������۹�/c����os�/]���p�zw�f���.{7�^�5���9�Z�^]�]�3ws��e�$�FB2��HE����8���my�i���x�J�{��T��E�m@�A�L��Pr���D� ���%�L�i����mF�����$��jR�I)���"�v�3���U�&ێ��ť5nV��<�����; Ժ��q�q�ww�g���-8�y���{Qm�w�l�T��zf)y��6�;�ν�R��NA���4_����V(VT���|�����f�y���O���ӧN���>:�� ������I�R+���9?����
���2[@Dd�eci+T*��H"�
�
�`�FBz��"�VJ��AJ���AC�]C�B U� ��r@��x����������|g��g����T@�;� ����)R��P(K�~@�
,u�0��̄QE"&@(�z�g;XdEH��3"��J����1�
��j�H̅J��%غ�Kj"jД�D��lY`%��&��,����t�ӧO��3��c1?����%h	iTOid�Ɣ���Z��j&.VV4�D��DB�f��%K֢�&j
b��3N��gN�:t�����c)>��_i��z�N�fch�E���mY���䢋휙ơ�S�|���������������ϧ=�{_x�g�/y����9�Ԩ�5��x�#�
��|�IJ#"��(d(���ۏoOON=����<{go�?
�Ne���L�)�s���)�&`��2#T���"�ϭE�5�C�W�a�ƕ$5�m�P�lz��?2����l�߻
(x���h��ږ�
�"�����H�kɜn��J�C*UC�(ņ%�ꔨ���M�F}�����i�@�\�:�^��q��wqu�����Mܥ1�����c��Թ�A������Ӷ��sK��.��W��Y{�Ca!6�� ��%�K����g�i[n��e�!�2�ów��NY):��&{�U �!ə!�@��=�㞷s0�S���^9�[^^�n���<����=R�:�\n�7�y/R�c����������vcz׭�j����*��j�;v����%.nK�z�n����{��ȧq�g�ܵ���b��
#�����ط�c���܊q���|"�# �;�渨�\W6�57��~�����̦�݌�ˢ�4fhᘣe�p���T *p���u���^�!Ix�g�PӺt��Ae��M��"�ʍW�-���/�U+�J:)��eu\[Bw�#t���\�7��^#�O�����x�Wh;K�Q�%\�k)'�wB�0�UG�j�I��o`c��L��Q�- �1r��4�"wM$p��Sy%or,[��d�+99^�Z%EH>#�F%`ll�c���6�ф��S~T����R)�
��Q ����d���VP�ݣ:d
}���
�D&���0\J�u��s�g�z{��ޫ�}��'-�"���{L{
d�}�� �;��J]��cdR��:n哀�b���.��2+O�@��EYRsӗ6�jN;�#�y���N
�N��Xg��B��ɕ.��_S�2�T���/H�w�Y�����}�`�|�Q�I�n��z�r���ڢ�����%c�b�}��[#�aΝ�n�u�^O:��kZ��e�V�h�[��.d���Y�e�d��N.�E���d���=|w�Ѐ������|;[��נ)��>X�'�'��@|�@��FvmCc̉S����ǛC��� �/*a�_d�3�Ӷ+��o��כĽ���!��Yo7��K���A��|���[�C��l��B��Pl�z=��c�z�$����ezV���	j��t�U��yw�1��Y��8��3
�Z�.���}K/$�@f��!�_�X�ͧ5W�̴R�h�E]`7�@g�{�Ϣ�W_O���89��&8�s�Y�����>P;)�!���ț�Լ:Md���L�SR�3��X�[����e�ͱ�d�/�*˕�����Oꈝ��5(,�=�[��iHr1�|�m����*5 �3[ l�wTY>��L{���f��s��Xi��0�Ib�x!S����>O���y#ude63��������"��DE��$�p �����rv��O4�������bE��kM���u�s)N��+V�7���c��s�K��NK�#��@SB8S��t��wD��C5�}lu��w���m�R��JΝ�{�Z+�W��xTA��ӢMb��+ӎ��F�Ҍ�Y�F}Zř��9�sm�2�ؾ�~v�C�3W���2	�z{$
�x[�򿽇���^�y��d���S�y�}���l��S��>�M?��T^���VA�Y�E�߷�V
|~>��X"�7��b=�UG�gN����j��y1"��']��E��:�
�{�ٚ�0q��6,H;��HS _��R��XKM-f�F�`���-�w����u�^����Gßyz��+��k��!�Cj�Ux�Ҫ���U��-�����k����K4��r{�I�x���E`���7ޙjWi�B������
��.E���D�{Xx[����\�������4�Z�X�eL1hw�+�^�/&��n��{��eUYdN,4+��H�ngF�x��v6�S�L�5T�.kK*K}_}�7�Wʇ-t��T������jVEI�8�x>��@�.$V��ˋ�#�E�fހ+1:���״Q$��$�'�F�,��=g�}-5��ꥼ�$H�+&\�z�'N�*R8쎾�&�`�ԧWT
�& 3��#�Uso'	�o⃓�ﳈ[�|I49�l����3��Ҷ�["%�9ѥ�ײt3��7jv��\��V͟}UW�V�����x_��5����HI���B�*z��~�s�a��~��LRQ�U0i[ն �W��)I�1���/):�w�b��R��>�qR͢)�v7*�)R��b�9�K&-�[L5Hx�	O�㋣�ՃafH4קKջ���|�������(|.�k���r�0/fy��k��IQu�j��r��\S5S��L�y�KV�-���NC�r�fE}q%��~�o��=��۞߮>x��~uf���룷^}���[St�wW�Jz͙�˛g}��L�H�Ƭ��_ۂ��;�+פ�����&�0`�ݼ�7�����Qr	�j*8�^Vy�h���C�8.xC���ѝ-6�����u�Xs�1�n=K��y �]k�����WޗvM^��C��Vj���`��;s{).��禷]/������F�z�Y���&��&*��f�Fa��2�����ԏ���'�O��.����f����=΀ Q'[m��d�ؽ]�����)�h֌[|�_�w�
A�p��w5<}QvW�Fi�>ܲ}��0�_o�������Vjd�Q�����8��;�6��׊rjx�&R��V�l#�P���۞"��F�QW%l�'ڗW*}�b������t](���|����Q�5 5rRf}��#�e�s:6�[�I]�H��#Sv�,��g�G�*��˭ѕǳ��e���~m�TcT9�[�㹺���i�Q~ڟUTx9M�C5��p�]�i���p���4�R��g�h~
͠���h���k�� JTy`�n60(�d���ft�T�vZ�g4��|V! *ͺv�֓MKV��|c��ܺҠRgf&CDO��JU��ӫ�*�)��d�_��g��S�%Ww1t|w#ovW{8?�oZ��)3�[��rW��IB�j����*�+�9:���Y������/t��EF0&;����^X�g%B_c�.*i�ڈ�b�gv��e-��M��N�)z�*�%>�E�%�.�D��x"����5����t��kS�mL���/eE��4l�7�F��R�ڛ}T釙����
"pU�wD֣��L�7�Ҕ���T|:��B��g��YRq�U��9Y������8�0d�c0�>;pJFY�Bѧ�s}[;�_�O�������4;_�x9S��[L��N�wf>b#/�Y*��䴭Lo4��c-�Bu����߻s'���x��z��J4[�'fҭ�ViY>ݬȭj�JǷ�<��I\m�*<�m� �څR�v�ܪ«gH)q�"6=6F�8bD=��
�gqӂ�O�~"��( �@�)8B�1}^�Z��5�rf��m�Ut���N���{x'y+�g�Ogʐ�(4Wbt:׾P�w�3�B�2i<�\�=t��<_<Q5o�٠Ӧ��O�j�Bwъİf���³eVC�`�<����ߚ�~�_��p�:���|j��L"
�W���&Om,%g����ӳn+K,�Ë)ޚ�m�Wګ�j�t'b�F���liaM�l��C����Z�zrf�Kl��}�[�İ���ou+Q�3K�άC 9�^v�I�����0�!�:�ì���צf�l��$#�
��L�Rb�\���M�pI��o%���:����O�XՒ�T�-S��a���3�׉	�U���B�� b
ǜ*��5I���4���|�e�}CM[&�Vm�`'	cUxC�Tm�i)�D���-���8���T�4<(�x�YW����${���a�_�}]�T��Y���+1&���Ӱ��!$+G���Y{�=�7G������$�R�� ,Y:*����8��*�$�zE;k_?�9늴��ݷ.2�"�ԵV����e ޟn���%
��*��%B�����gymd᥾uv�o�g�a91�-�����j=i��s;�-��~m���P_�=����^y�ޏ�+ʏ=`��*� ��M�szc<K��#����^��ua3�K��TQ���N'�<b��o3h�Yo�:���s-y�K�w<C��6���fN�Պ�.��l��z~�Y�C�B����t���Ӽ�*�X�E��f���=����3S�;Q�^.+_NŮG�HO�M����W��a�յXv.̚�<�VL&S��z;R�m�����0]=}���d�+�5��"+/�#Tt��&�6��)!�M58�rΧX�=�L���;�6Y���(шӋ����`69������T����t�\U�//0��a��"$׾�w��Mɹ~��yC�,X�	��%�d�h��ёO��-
0XAcݫR>�gm��0.�d^o��~T�V�%YiC��{��yE����$0�]��u���V�U� To9���;;��T+�L�da��R|x�4/I�6J��ݶ�w��ܘY^�͎T�y���L���M��9���VNW�-�4�Lԇ�g��|��1�n�#m�^���z�����o���[ټ�����b?x��&OI�{y_;;"�PF��4(?P�ϼ�>����GHR�],úOIv5	9��7yP!yqȫ6`AW=��-grN��$�ԪC#ޙO��c�����/pr+}�μ�]�c�v��*-V/z��3�aIپ���d��S�JZ�����=�D���4hK� P$Az]�r-9�!���{ٳ8��nD��2�)!�s3%�%&`�N"�*�:k2<f}�������^L,���ZV���6�.�w��==���a-텘6���؁�KW��nz��P$3�d�.�uT�F��w贲�i�����T���5`4i���e�V_V�X}a6��a-[bb����y����Y�5��ju��O��i$@��9
��y�$�`��,5Pq��R�ήقf���@��p0�B(�bn�����(N?���H�qy��e���(��J��"����D��!f�d�!kk$lO�xGE����T_xХ��E���5+�F-L�^ZS'.|ш�s>�f~���	��\[�2�wΧ��A�C%Ô���δQD�MW����Y)�҆�u^W]E,sm�R�-�ݜ�Ev*�O��`]��몜50�=5O�B�H��|�;Ӽu���-L<~	a���hL�"�'�RӾa�B��g�1=Im���WJ��}��8N��;��^�U�ʢ(��gc�K���n��J�KK�3��9��w�+�p�8�����;��4����zKI�r���7����g(Y�.s)�z�� �C>l�}����vY�72�g_�^�=�0�[됶�}�q�l��yRj�3L,�����^(1q�)t�Y��N��0nNM!R�X�E�е�5$�MID��+ٌOvϼ����z��MS�-5$���7�)��em+��vMH����gL�3VS^�F�ީ��V����af;�Y��^�;��x�Z���t�S�{�ψ�)���1�[���Ϲw�J{�n,[c;����oG�Ʊ��F0���Ѝ��x�{7e�6%{6�*�췚3*]�f��{�*��mʹ0�D����z�5RA���ʷ3*�[;3L����������Dy;�S���g��В������Ѱ���ʋn��.}@j�f�f�f�[���Ɓ���<��#�!�y��f^Ggj�cI��ր����Tb]�փ6�vѮ�t�B�=�)n�wA`��}�1y8�6l�x蕖��r�9to\��\n"[�'IO�$&���ZZn1��W١ʱ�6�^<(tq��5��7#�[�t�X:'��s��ޫ��Sk���ԃ�=W�6Q{sx�3���<�ٛ�V���wa����S�Sƚ`�枮hN�՛w�e�rY���,��Y��#�̼�)84�|h�F{���xNR���v3*R�t[Ui��fG��2ۍ����V;+vWn��Ɯ�.�)1C�2:ѕ��VgGq2�A�.�_]έ�W3�'�Q�Hnf���S��y�)ڰ4�*����0l�d�6�0+n�o�� �!@5*�ˮ�<*�Eu<]1����O^���f�_�ٻ�V@W��>�O���y�nvP� 9BUŇev�,��9y��X�/_=��bG�Y{N�.�����:w_H�yG�]1 �Ĵ�y�^`h�[Y�.��W�����յ�z섩Q2�,�@O�a�1�W�mlёzΒ�ʆpS%A�n�!�:�+tl�=��O�G}1���W�����e�Ku$�RA$J�ʔ��t��2�B��ISa��@����/q��=��yL��s^���T��`�{���7D6���e���emļ	y��
�
t��@_jh���7=�5��(r���:>��Sw5���̝m#� R<@W�N��b���O/k^9o�qf�>�w�,�������/{6e�i�xr�#ss.)Zu���T�c�(^��#��ݓI���t8ᷪ����ɡ-c[7\3$T���ƛ� �d��ڴ�e��MBp� --9BnF��&]�ąC��W��{J�jt)^��tr=�Pj2:[G�F����������6[�GiZrU��1:���k�L؋��9W��$@� {��H��8��gpڔ�:T�c*��D�Iy2���8���ߤ�'�c%a6�BE� \2+�� �*S�3�t��$�M�e��jU�w�^�+�<y�9�:;��p���[�!���ٝ&*Ej����7�rQea�Zm���zvs��eM�֦[�+�>��=�y-�q=��x�\�Բw[�V���u_H�Z���t�0v��,�&�Ֆ�[�]�sv�M#�;������z.�{�iM�
�̃T�����|U��y�ʰ�T����%���]5��vQ�gٕP<@�S�a�eb�EWS'2�<�" Q��2i3���}{zzzzq�>:����5���3�r��
u�"������������E�ȧ�DXug����������Y�_Y�=3������&b�VLb�)5X�,[q�-��H�����i���������|}}f~?�d��s�E���j�]jT*y�fR����j[eA�e�{=�N�:t��g����4g�Bz��AH�g���IX��z�T֓[V���~?_^ޞ���G__Y����>i^�AO\��ɝ����,.��\�x߸��˩V�T*\[j³<~=���===8?__Y�>����C�(�E�Q�.��h�ȍ�m?'��/���խ*��=��,>��C�y�BM�s4Q���[J�4���+@�)QEF.��8ehΥV�X�]k�g�g�yo�j����v�)UUz�5Z�Y+m��C9�U���vʳ�a>�uʌ�3�]���j(x�.�0Z
�+'�s�쾧�Y��YR4�s=Y���θ�\�]8�����|������۳�Cv���ۀ}���3���0���0}7�\���bO;��cb�i� a$	�7��)Z@�nA��X����ח���Wv��:���kz�; ���0M���S�C��V�<�	�����xN�H^ A�Ȋ~�+�i����:YБ�1�^gɐ$|�y ��x@��0�l]��=���*K�o�zb��M�<��w�s�s 0�Ԝ
��p(˶|�M1bE*>>�2���]���b��v37����=��@��y��+�>W�7����DV�yTDP2��
J���,�~�~�\��V�>��|%��џ�v~�M,x��CkPo�Ǽ����Pd�F(g�g��8��"@Â� !�'cC��㻗������x&�wD�n��L޼�`3�.�G��o$: �p.�N�Lxv�vy���G��χ�>I�].�d�0��.$\� �g�oѭ�^R��6�^���5��{%�����5�����{�7�&NRo��C��;W��yS���Ӭ�-�Nq`��z��H�� |�L�̗�̔���pމv�Ȥ��U�<���}��Ņ i�`q����9�-��&\����|���H�����D���%j�[��Z������̗��,�ހ��J2��{�ט��H���H��T��T�߆�W�o4{ؓêi�𮣦�%�۝�W؟B�s7�a�|Xs���7�oK6:�Q������o�]w��Ϭ�#Yc+,H�81Z�	 <�1�W<�{'�a�1�v�$�с��[��>L K@zao|�Af��h΁L��ů�E?e�V���0�l0:��p����^�����P�f��ff�������2�&�ݥ�2s������| <
鹠X4)�l����#�ϜiB�@���=�� V�ncjЉ�!�$���`�H��k�h�����x@j�o$���-ѽ-���_�쀹�5�5�$����,5�t@���h�����j/�I�xf`3�9/�8 9����c���[^��b�|0�7��cx,�7�-ᑎ&�m��S�"�.�>��atHF4�/8L�-W�A`|}�r���1PDo�4+ʥ�S�m���!�x��ak�7��Tk9$5��#�Rp4�� }LKY�@58@���W�H�����u[E`�W���9[�� ��;s3!�0f���R7��ܠ����@e5�^?|�fE��1��~���S6َ{��X���P�b�|��)����1�y�P.=,��� ���S�T��&]��{����T��D|+��;g�H;��x}�΃��|�vI���f!��ض��J�&Mm�F��w��f�����J��>g<x�ɖ�T�l�dҶ�u��%�=B��Y`q�$��>���� 7qj��xqӑoN�ΓY�n�ծ�9M�uӴ�.̨������{:��
OC�h����Y�����޳7��9/���g��~2�fX����>r|�n��^]ץ�a�|��=���m�J�2�JNxm��c������ݺ��Z����?u�<%��z���0{Tcx+Q"�Ú���)�3�o)t�����Y�Y�R�5/{:��OJq����p���N�D06����_�Ò�9�2 �nO�:�\l��?2��;��%��1�0>��*f1�p����?#��^A˹|��#�H:�'��9�p*��d��ů)�_����������e@ڟM�5�Ґ�E�+�4Á����G��nY�jvi,=Q�Y��o	3�\.7vǽ����༲5I�_ݿLhR� �!@���^��$� �j��A�����>���7�9Oᦣ��wo��������
5W-0�
� �avI񐇲R���PvOgSS{1ݼ9�����큋�u�]��N*��˜ۮ)��A`�� �z��h�:rrS����a|�u�.$lȄ\|y!�1�@I�]��������7Е�n ����{h"���k����&=���h�	@tg�nJͬ���*|[`a!���ʈ�� ?���t��v��Hƴ���y��sy�*�Zy�)�ң�:�}b�vG���2#� �zȟqEJ>��1=�
�G�f�ˍwȏ}3�R�&q��Y;ji*|���5�7�@��Mδiwԫ1	�Y����:���'ֹ�׭�O�.�Ґ��^#��TA걮�n�����Du�a�ڧ���e�ЎӻԮ<޽�k�=����[���pV=�ڙ}�(}��j���I������Ώ<�׽{�N���	@�Si��`x�P��2H��)8��֚���1S�|�ª�S�tjUU�v�E�Fy�k�8�w`([�>5B^P�4��,1}���Λ/˚Z�m�٠���aVxx7w��,�q�g���g���M��c�� ���/�>>�<�v��3ɶA)�t��L��|}{0�wk����.x�A�Q��Ϟ��s�����E5��!���7��چL�J���K^��{�����fܶ��*J̥f���F�jc�w�\��)��3v�u9�:��c����+���\�,ַ�]Ȝ�Sjm�)���R�1�+�����2��{��pw.Y!C(��!��<���qY6رL�s�<�oq�ް��Ɇ�3q��5<�b�k��y=���H�msw-����:�5�<�0���vҫn�����+���
h�{h��Z��]��l�7�aa�ە�D�P1�]�C��L�¼�
t�Ϭ{�Ab�>�'zT���u=f�E6�d}��0?����a�ώ����5�[�g�=��<{]u�R�m�W\]��eI�Cm㭍̇lԥf+�.fƺ��{����� �>�n��t6����q����qѕ�ut���2u-�K-��3���\N��=v��%X�3�Z�|Eh�}y�k�zg'�3�'�3<O�|�q��^�q[�X��8���HN}>���z� L@we��+�M�#���C�E_Tpo�t�,����]##��LQ���ThR1̉�M�\���*N�i���m,z��V�r�{������e	�X�l�y�ZPY���E�I�|���-�)����bu<���o��6�������:`$>G'���ߞ��9$�茋WD񨰉Z����'����z��;�5��J �Q�j߉>|�)���3Ӱ\�(ٔ��w���S3\])����<�,b���������<,� ���~��J=��#P�uˇ1��JCo|@�G�zd�u}�?;��U�?���M��|;�`SL�p�YY�e�|ST}�����Վ��D?�/U�\���Z�]��е��n:�'�R�uC3���VAxx��kT�c��EUO9O��$;��50�Y��W<^�3�Afh�~���;���My^6�SV@a{�LPfm�\���J{R˭�̝�;��]>�g�!�����K*�Y\�߅�ڜ���0�6���_͋�-�O=���^gr�����#FPU�����t�i�B��o[���\6�����v��c%H;�=?�d�9�����k�>����_���>�6>�鏻M)��]��Z����^��. �}.�qݺ��\�����jvc}b-�8m��ñrڃ����
��`�"!<j�� (t��gP�*Ho�q�<�T-H�U�Ә�atKyj���k���j�������v�kz��3��m�ikaV�f�Y�N�%q�/���k9Yb:5Y1R
�ݎ���
48�!����5)LH��}R��9��x��>D�zM �|�N��}�A=s��=L̂#¸����q�7{Q��۞�dw!]��O�ƪRD��"�O���ql���a�Z犹m�Qۗy�Ԕ>s�,�a5�7�(�;1�A�c��|n�cS�,��)��)@��z�'b��m�gv�V�1��~��H�{c�d{�T��x�a��d{ˋ�*����瘟n����s=xS��EPޒ�-�p���FX��#���2f

�S���<7�����5ũK��pgڸM~�������雑;���͘Ł�Pƺ��R�ZJ�>t��s�!��,��7�=��>��
�$d/�zC�*�NG��u݈������^�-$@�v�`+zOM�s
��H�ə�����<t�eӽ@0h��bFI ����2F�pE\�~�<��ե{u�Dѷ��I�W��F3��u>��7��EbA�N��4��:��ۙR�0�cf�x�6�����k��:�ι�Y:MѺ�xt.P��M]/��8������W6�Z�V���CH
��%�%���>������q�s^V�.1�g{=�;�w%��	�(E�8]Mj�����Oe<��/uE	���S�J>�4�zdy�>5U��:�XY�ϧ10�l����M���Lu:�f��q�.��5��Y��+���tk�����N�P�s�Y�T�7���r��qm��z�@v�c���H�A�br�l�J{�m	-g��j4��c���r�����M���!�.?���i���P��fmp(��\�uЮ��V��5bɈs0���CS(ܖ���t6����q��Ns�r~O�S�'��
��I�49x�k()�������XY��oh�"o>�
p�ڨʇ'�B�_aʲc�l�b���;��R$vZ歊m�}�=��+���VL�D?� R��M��%�b�0LLw�@Q�����0� !�݋m�e�|�������%���տ��zO,��Ҙfnz��{��[����l�z,u?b����ӆ~�?a�_���:�"��q��QҠe�N|O��HS���e�ao :��^�N�P�v�c�.���جv``��Z�����m�<5z s����z�);x�'���U�!�6��>!�:8{�-ĸK��F*��36ߚ I����v�<o���9h�V_N��ȱ�x�	����CV��КR[�_Jr�0��T�x�gW"U
�����̓��#�E-��/��x��`����c��������?D@D8�D<WgK�-���hb!���~�T{`
�W^|�8��\�_·ܤ��|�:�Տβ�f������\u��f��L1�>J@_>�L�/�d�?Hu��#���7��v��I	�>N�cU5��I�r�(Β��vg��H�,"���F>!�M{�3����ԧ[���m�h�U�w�ϻ)��~j���)�J�Tg�m�%�7��:���Hz�J#�'�i�-�ׯٷ��A�}�� r$Q�Pɏ0_��zLr��ڻ'#<�ZS/^'	�H��Ǯ�K�(�9��G{��M"�g�^CI�l�8��K���`hC�ߧ�t�ǝ�ј}|�QBN����˸�a���%)�Ɓr�(���������I�!��>��Ӿ�x��w �ex��9g�<�2�n�ך�;)�a�(�㼔B�^TGy�fS	�&���<�C���S�Ȕ*�������`����@\��̆ҍR�NF��#�Lp�����#=s3/�SvR!Y�K�8@F��1_�;ٓ�GDK^�E�2���]�N��x"i�`����fX�옇�ݸ��{��ݭ��T�s���HA��ީ��#wu����I2�'�.+u9�`oH*�j�֌�R�:H�KY�[6zyvA�%�]u�z޷�ъ�F
B��+�	G5a����g9�������啘��:A��.�lf�5ͅ4ֵ/F����w�"�@	H�3�i�Ά(to����G��7e���TO�E�sq�@a1�}u�O�w�b��6�r��H��#s7	�݅܁X�� Xcl�t/�n���^��9�l�bTKt����8�I�&�Ovvk��㜈K3nVqc�/���M@M��tq}b����\g����	�s;G��B��5'��MjND*'9�����0�5!|�E4S�<�<zz��u�I�e�u�����kwO9-���-ev��S��BC��U)��je�"�0~��ߝ��V>GɅLd����$ɀ�|v�ԩZ��f��-Q#��v�Δ���y�p����9�����J���AGhKBa-	���S��}�aN��4S�g��a�;��b�~��ӽ�ǣ[*�u��i�zt�w�2Lr ��%��.tz���*x�0S����OK[^���|p��Y��ְ֯@���ޞ}<���D�׍]�j��'p�P��S�-zX���eVL<>��}B�c%YA.����p�|>$�7 �+g4�ɑ�+����Μ��t������Bk�}�Q��3ْ���2q��ᆱ�J௦�n��W����׆�%�[�i�)3�Wo�֎2���f��G �OtJ:l�v��������B(�`�Rw�-���gKR�pc�e.����z#Q��-�v��7	M��T�t,��}�w�����:��?�2o�0�.x{�����.���q��"�f�<��2�9 �<� � �(.��q�c�]������تkq.��!�'�3�q���h�8����r��[qo���B�rb�@Ɩ1EZ�p2&�9�Fp��3!�r��)�����j'Ae��&�O��e�9�6���0�c���6�H��9���U�79�q���ҏ�I��E�{�=�yU��CJ�o2]����m�a\�:g��U2���<�p��zKzBp�a�ｑ�Vsf��e\\҈� ��>p�ԅ�7��R���qk���`���|ak�i�.�/k�s^�uhb�]�7f�g�S���G�pp�u�g�B���+zL�O|��qj�xy����_=$�'\��W��M�l��o��ᙃ[�(��� ���8�=%��8��ӭ���.D��6��5����m3��{�T��m�4 �a�vD��k��~l�[
4�KY��?�&�kr��r�?�$��WT(��sS8��}�D�CRma)+h�k��̢��Ϸ�N��<5��S7�M��|ڶ q=Z@����Cv?3�����
�v ����������si�G�և�R�d�]jN�����p[��QG��r�Jo�f���g�j���p�����0���)����x��i:����T8�oU���ư��<޾O,�>	�%P/�%��ʘ�g�[[�t��%�4̕�m8mz�Yp6�5ni[��X���$hj���cn�u�yN���&(d��.��iDw\��5�6����ibd�m�Bh/	�[�A���yO]n�er`X������vz���4/m��=�<�g1G�̩��%�{�|]e��0�B��n�(�x��Joda*ƅ�Y�����^��b��+5C^��˜�Ͳe��ģ0A"�8�	.jƼ�nhmN���W�]��8,���痼��b��Y�mw,�>]]�tr�|��¯���}��e1Z���ę7��[�,#��B���.L�8�	��1��u�7�,!\�"����<D���1OT Wr#�0����
n�wn2v���i ��׸�g���-{�aٔqJn�/kp��L,7x� �E�\�Abܬ�Z�%{�N��}[O�R����f��"u=�e�F� *��6�Q���A�:�#¶�j���t���{]Rۭ���AV˖,-w5����i�=V��Ǡ>�nفM;v�ވh�5���-%���c�����J�C��IJ�H��U�^z�裡o[��lĎ9yI+,��KUa�;mr���Kn�#����W\�����1<��X��e��"]9�C��oR	@�ޔ����р�WP����U��gr�κ��ν��j��淋:��s�'�=�`��Ρ(�N�^k9w��F�Ju� �br��x�fNR�P}�d&a�;�i�㹽7O��=lIR���}:v_��`������x@��6��pJk2�5�/�>�{3��o��c���{(���]�{3w檙]�eO��.�dV�8l>-p��|sݓ�������j���L;R�+����Z�ۯ�6g݋����L�ҖyR:��]���(P�8�y�;����#��&Q\,Uʓ���� &U��*qg:�K�l��Ưl��H�[">=N�K�->��';%Zc@��W��ul�n�*C�VQbȲ.�l"Ŗɔ�/8�r��记�v��o+*�P���9Asݻwm!p������<����zh˖^*l�]��o�Tb�o[��+��t�=[�ތ'7xc	h�ޝ/x����'[����ѻ��,R�����1��Y,+����4�3�WAtgFP��(벞s4��Ĩ��oB��CTU��[�eӭ�G{�1$���=�\2���3 D>�@q�f.1���vv7v�秓�ʺš;��R��Δ�C��oQk�����5�K+���&��\z�+堪Q9F�D��m�ن�b�(����%>��)J*ל�����đ�ݪ"�Z���3:39uS֧�Q�V��,g��?O����ӧ���^3�ѝ�*d���z��D��m��r�?�յkYV<���(��Y�Vٜ	Y�i����������]}x�Y�c���>P��ѡ�\ʖآ*fV_Nh�+Z�DD��L��ٞ�+��τ�x��{}~����ӣ㯯�����S���^"ş-�`��E���+����Qk-��ں��g�ǧ��q����|}}x�gO�(z2��[S���i����J��J��AGT�Ҷ����r�3Ǐ����{{zt}}}�2�џ ==����**R��
���Ǭ��j�DR�fǭ��"�1���	�<z{}|qǷ�������<u�4�
#�9'9=�ڕ�9�%U4��c�=C�3�Z�D�Z"0P��Gm֩��4�b���L z�4
Ȫ����������W���Tdu�>u��E�N�8dm*TWY�3���|�P���#I@SI��e�hj���X]T�,+6�������j�ݑq{u���J^ۋ�bٯJV�{�ܜu��qw3��w9[\�5��{��מ��Shh�.AnK�ɑ22�{2��Qs��y���U�]֑l�M�M�gX�s��
������:����l�m�.����e�)���3$�R���a�Ln�U�xN�u{=ש�8����q�7qQݚu���=8T�w;rc�Tn绵9�rZ�n�ۨ��J�s��׻"�iy��{;[��F���D�.L�&d�H�bAs���jL�q��qn��n�q��@��aH�FT)?�$�>�/�~���u	��NXi���|�;���$ʆ�"�S�Z�݅�s۲^�*�^gqSH�[e��)�G�a�5~Y���!��7��Trbbg�8F4E!܄�C�ǟC�y�V�\���Vn?2�#M��)A�{�|P��ίz^��H}�$n�����[<VH*�'��S���ek���fFe�##���;�_�޹��L2t^�� kmuq�Hϫ�	�(TjU��-\Y�VU52j�y��:ny�Ƙ���(M|��Kx�0JZ��H�w��󋆟<[���>�β��ܴtǠk�Y^����H���JGǍ����$���dˋ�J"�ۣ�*��}+�e�s�5�拕�i݀�1���s�1cAU�ޛkk��Tņ}0*�[nfb�,.���?y(�
{��N3�-���J>��l�>~��J{�"ږ���a�3})�+�'�/��f���B�~���%�۠d��] d��:3k�AT�çGL{����P~u��%m��C^nwϙ�L�A�d�`|�|:����,eWz*A/�G�E�&�ym��+�C*�����x/5�x]�E�Q����D�y����c�K��C�""-B�l�w���>FU�ⱀ�܄�x�� !�˫���K����#a۞��C9���Px�i�]|�&��eE ���[{;��3>Ѣ�׍�|PtQ�/�q�&�Ų�p� �lX2a�]BQJ��ޕ�;Z���cn��ڋϦ|����7����w����$2�'*C�b 	3$�`��Ĝ��g��n�m:�}s��:����ׯ��+�ɘ��lZąD[D�}8Q��{IϚCUUYפ�x�jM<|��q�׀�)�� ����?�yk.m)�W+�mp'ә.��a�m+ �+�Q�}Ç����*+4ȣ�2\ ���N��՛ʎ`va6�2��}ܢ�:����c�C�S�0#b�/�װ;_.�������n1��x3(��Ӕ�֤=�)�x�a�֠:;��z�\aR~U�׃?���L�� 2�X�*��5��[���V`m�5��)��5㾎c>0�ce���:�y����Ez)�c\Srvc�0�����ʄ���*��\|�f_'>��D�֟����t�e��_݃�r$.T�D���>�nb���J-��� �K�b�������[��=ytRA�j���!le�������9���&��c�^�^�&;�̎}�&�3"R�-F���}8^��a���x]o|n3ЛNJ���f��i�����:���`�嘇������Ɗ�UW�D��L�?'7�-�����Gº���q k�yIbdծp�2#�ɥ���L�D�� �&�i%UR�_�o���<�ԏ������vd#I���Y���%�����h��on��ʛuB: P�$x�ܷ�믇�FM}R�ϸ�܉���5j�=6T�$X��W]f��s���޶�rP<�;m_R�V�]�x��M4:Q��ߟ~�����?��e^�
��N�C/��}�}���Y�<@/�̔vDzd���y��vcد)�GlIqez�I��|
���qޤש�j�ߡ���O�"@��+}pz�z�Dn�+�h�+Ɗ��&G g����4o�d2'���@T�*�3O�X;.^=_q\:�r��/�TL(��ĩ, S<�v/Q�k�#c"w��Kt��[1Lv`Y-�M`H]]�������~�.�����D4yM��[���5%(�����o��c-��"�$U�?Ddxd��E
wLa��X��(���vV/8?7slb��.��5 B����{*����wz cc[g�X���0|b��?0���*�Kln��m�T����r��ou[^1c���õ�ji�}!�D6?���χt�qED��r���7ѬM^o)Ur���a�{�O��c���*�"�&��p�*QQ�AD�c�??UzKz��ʄ��:�=3�SPp�6�X�?���`}��xxז�s��i` qG�\'�ƺeO���|� ���.d?�����^�ҕX�4  �� {�+��<�
>4~������!����τ��<���G�EtL!,0Uq���1���>���7sc`)'N�6�s�E�Y����4��+Ss�/A��3v��ϗ#�\&"�������;z뫫P���\;����S�B�E��ޱz�.�n�Ë���J�R�e����>��:���~+!�'�f����0�#$a&`<�����/�{���}���i�-�6[x�w�.b|��3�nd�9v�KBZ8P\���$�sǆ:��*���Z�)����@x�X���S�3����i�f֢��jpr�Y�|��y�RɉrJ!2F I�2�˧�@���b���61a��cpb��yV!���g�3�����%]-<2�z�ݷx<��E����������i�Ө�3�kʟ0�l;8L�9�K�Vm�y�Z/� C/d�ט�޼��2��hϜ�/��A�g�91���m��=�?Q�6)����=}�)N������صz$��~�x���1:��FGNL��ؚ�S�f|��I̞��~^����N+:/�7<�ly�M"�q��yz����R�,538g��<�]{�{v�f��:Ӯ�f��
�	`���P��tTL{�=O$�.�r۶��4k_8���ծ�E��Z���|�}bvI+���,ey��3>8��Ş�����׋i�9c�\�|�H��t�=����vw`��k8k��	ז��v�EC���+�@�p�Z�h�/����˽ȍ�6J��q/�6�Kq�}}��n�ڽT��P�J��PC�`n�Z�Syr�NF��O�/�2#Qo�:��t�ͧ-�=Y5n�e�k�m�zG�b�n]e(Vk=�+�Χ��N.d%�Lf��V��茹��Xh�~�E�D	���S�Ȅ2�#�P:�Zޜ��I��z��b�kg~��m��/3S�Y�m�cs�]y��J�;���T�*����9*#w�|<���ih}�,���`ɉݑ9�$/2�"�˳��k@�ӫ���ֻ�t:�ںw����o�|�'�Z�17�hm�|�-���^�z�-"��ϞN[x��w�8BV/����v�y{h=S�쿹t-Y�{�m�$s(��E�fb�܍�x��1�B��1��M��2'�V0���b���8v�<����,��,�~���kC�&pg��þ��x��ZD?s�Sߪ=�T	�`ީa9q�y�dz��Ռ����;�d=�jZ	 W��$����>>.P߼�.
���@����l�{X[?� $ז�����v�� �)?f:�yx�F�f�W�T���;������C�s�_��]9!��ܼ@f �����p>�C�4����=Aѿ"V�8n��E�w��H_t/�9��FK����3"����9?U|x{�(�Z��2_�ʔ�"�˖
�dY�(*�H������r|k��H�X:C���6��*�M40����v&�����;ǜM��qrn	Ϝ�br&F����:$�=}馽]��O�f�7��px�,���j��p�37+0WT�����f+\�E1ս����9�],��QE|�⿗��(�k[<m۞��( mB!�F%�m8$�E <�;�w�}�r�,Z}]�4⏾�Zyk���ˎ,�T��m��-Sq�s���_+�t����Xd�Ta�DTռ���"=����Zn���B��\b���,fC}^鶀S�qSܴ��Fc�^`��=�۷���#�w�����	]HĊt�#�0(���
2�`�+�+E�����&sN�
�Gᚰ	�S��EҲ�y��@�&��~�+��(�ˢItC��t��謐T����c�nB&.�S{��a��ߵ5j�Ȝ5*|��c�#��\8s-��j��{��n����qM��>Q}�ڼܖU
��_�w�fx^s�W)SS�{X��fq܉��	��̫�}���'㸡���0��N9�:����@q/���O�뀟,q�%NFE/.��Dhvӵ�>7_NQ�<2�,�Yf��-?C_�|���NAu�������.����h�]o���3�5h�U�Z;_�in/��c��be+R����ϥ�����0���YN7ם%���z���y@1w����׹,"����w��Ǧ���$E��_�0`�ɟ�>~�!�to�T�8*QqW����[L�Nk{4��'���o�ע��A����{�|�x{�����ة{�F%}/'L,�K�=�؋r�
��*��4|CR\݇5 ���>[�r�l�.���_�l�cZB�n\�t4|�zMT����=8L{��k��ڇ7p<5��Oiel�mD�L�9e3]�7�C��e��u�Y[�#�~(��{(��a�Xax���ʡ�O7���y���O{cTϘ��	�ثp�T�b��2�v�~�4ڿHW��"���$o�/�j�fӾR�J�ޖ��t�����	L��F�2OBTx�a���NY�۳$6����n���N? ��~�m~a"��l�S����rT��p��~���$�)*�f�[9=5�E��ͨ��\5��ԈoH���
�s�y�5iZ��h���i,/C�#ڤO�^p�.^xS]2�:��&]��$4���}-ڐ�:-}ж���b��f<2{C�څ�@A�?n��~����4�11@US���ip ��.Wz`E�G��ƏL[;Lc����YP�<�����w��h��}�>m��΍�1�B����w�#8 �<:G��X��[�2'=rڑʌ#f]�9鶨q-S�~b���_TU�Q��\0��q����i���%X��}XFX���������	]�	Q���-�GY���Ɲ�g4Kn���4
�
F�@��e�<:e�=Z���we`][��zg�춌��LU��Un���a]p/�G�{�E�V�8��%�
�M���ute����c���Ї�.�ZX;���-�r0V[��y����H��iꛈ�89��z�9������=�{�Ƴ;۞U��i�ݙ�l�称r���q��I���3]��{�%)qK��p<o	*��2>k���Ϝ��U�D�"p`Se�C*r 82 r���AJ� ���~�{��Tq���Y��.w��5c�o_tqq@�*�	��[gl�W����,x~�)B�M��;LH�H�G�KgJ�O�O������lR"�@O�yB6@f�M�B�R��6�F�(�S>�|~��5:���������vwA8!��ͥ���5���نi�x2�^d��v� ,���^�F���ր��~�`?1�2{��T�r&cdH-c��$�y^��������ՁdK��eoR#�g�a������z�1�:x��|e��^Mr�����r0���t�	'xѫ����p� û���=��>=����%Ha���+�qE�Qe���`��I�e�o�ٴa��C3u;G�%�	��`W�taz��s遲�dah�]��51��s�٣+�1=7dD�?����;"��_��u�~, �Uߍ>YM!�&�U
�Hu���5�J�!��N�8�̘�cT���p��8'�����zr���k�7��1G�[q:��Y����Z<���5�@����P�J�1ȟF��JT2tZ�Hި]KV>���Q1B����bzDy�U��2Su6��>=݊�G��C��1�~��O��� #$Q�G6���TE�R�,� b^fᛜF�V�K�k����E|����܊uxe_n*��Z�ͮl�҈��}<\�K9�Bj�π�bDt�%#���R	��^B#$�	)$IR@'��}��o�r�`L�$�#2�I(���3�~�3��99�^����ʬ����e9% ���L�$���R��I�(B�g ��x�TMq���M��p��c;Բ�+m� )+�D��څ�4]�ѳ��d
�,6��]Ԇ�=鱷�^��y�����wmSw,�;�9=>G����/߷���Bn��F���m�ޞq�X�u�)���?4�-��1��	��1�[ыO]�y6���90�/>���=����y�$Z�z&��(���חm�2�J���:�.��xkˁ+�հ��sr� J��c����6H�a0]��l���d4��}�d���4�MM�\bs�<���#��#��.�I��-�+oD)� �*/�X#o>t-u\�5�����aݐ��Ɏ�lt��J���v��T7�mE���T�)�Cq�Zr.B�ׇe�r8���t>���������0�p4���s/�c�Ϡ,�l��w�����&%��ۃi$�Hn�����U)���Ek~Q����>��)ޒ�i�=��go�ӽ�$��k�Z�w�,̻���q�W�/�7�a�H�,�D���(�ւ����lu+������r�Uj���1�*F�/n.����-i�]}��R4�"�8��73�'!\�VY���X�kcl�U�[����R�X	 P��A�s�󽯇$�\��^cǐ�S%<ɩ�x7�����v;�\1�ӏ!�U��Y]R ����о~��a�XeQ�Ea��J*������{��	�a^'��M�j��t�0�c�2|�Eݟ��$@~o[m\y_@��b��t�\��:���FG�w�7��>n�5>� ƿ^�mTj�Lty��y5�������l뾭|�Z�K3k�7�&��$3ז�߹�nH����(a?sd��"�L�U�oN=��{��|o�˞���v�N���5��Bf=����� 3�k�_sgV�e�c�|�w=�=�X�G�ܮ.��Ю}`�#�&Iӧ����^�p�4�5��H���3�3</}��{��SC떹m7��OED�Ϝ
�STҢ>�<
9��˾��z��ق��޺'������@��"��xP���}XbFm��JG,���'�(��g���88�%�s�NS������>��L��1a:���q�+�Ӌ��۸�,D.>�<"���-�G|�|�Qz��s?���~�����s}^�������B����|�霗�|pSH� �Ӎ�Q�u��[��s4à �Ʈ�� 4Q^���ˏk��C�~he�yG�=��C($kv�!����������V��m�=IG*Oߴ�6�ٔ����d�#o���)'tT�Z+6S�ʱ��y��|�YNB��������4�I�|#��W:}��;�XN�kar�λ�z�T#�aP��:	�s�]�.8."��[������ĝt|�WwG�s�j�1�.��t`P��T���S� 3%jh���ՙwS�����h=�V�sq��Uc=x#T�O쩸�;f�^�rv-�����WK�����J��ԛ  j\y���1�79K�@�:�ޭꝳ�n��U��>��o^d������m��K^��j=�a.�����YL���=7�����G��Fv�Tu��x�/��ڶe]�aq7+��+���ٽ`�����HZ�]M�\���c�_Wgm �+S:��w%s�I��sщ2��ķ�`��̼��m�[�ru�bSh���bL�����n�YI�#�s����)7޷^���Ovyc�{ ��:1]'V:牍9�e�ַ����fm9�\zv�.g�����[ƛe�n�R�m���9ݙ�V���З��&���,ᇸ&V�q�!�ub�MmV��c$�����HpU�d��H��T����LIS���t�ٙ���[���8�`$�<bU�7��rVC�_�'~�9�җ�JĪE�N��@$�j�g��E�I�e.�z������*�1�#L�n�
Z�	��ęE�&�p}����H���VHP�܈,�`S'��iSF����6�	Ѿ�Z�����n���������o$|(_r��'-]�m�+;��\a��d��o�h�QE6S���[�jw)H\|�楾­o���`��Mb*�,��"$��qy�4���*�p��I�^�ښ�䛲4�Rd�R�ؗ�U���0�n�����;A6nW#(x�[6yT������\O������N�AS�����7e�鬞��@�n�֞<�.�Mӎ�f��Jl�0̬��ۥK�V��B�������#��"v��h}Kqlꎌ��4� ��b��ۛ�R�Rl�O�<����k���_<z��{뭥z�"�TO1,���a,��}�q�:�5dN�>c(=�F��6�5��듚�n�n�49�v���vCm\�n���[6*���,�����SH+g>�f͔8�d�r�X=������i�)��aW�j��d�s6>(���aPӪ3�w��*�=��+�u�t�{8�&>@��ha����3�K8
�t�ي]�����D�'y���31� a�Z;��V���r�8�2ܛQ~`�|@ �(�F�j(2*)���ԟ���jlYu*�F
���I|���O��8����>:��:Ͼ�F�p9���s��L\�(�emh;i�֭Z���S{ረ�!;W�q������8���}x�g�����O$8�E���E�6�f�ֈF��h�*J���_p���S�=?����q���>���:Ξ^��"�Å}��ӾO�
��e�]���0l���1vR#Tm�3U�Q��M=�Mq��ߣ���Ǐg�o^�s��U1��V���G��_nL�ո*�*��ej[+���z}{~������������u=�<��*X�0�Kn`�U�V)�䥵��Zd�X�4ϯ�o�{{}__^<x�ξ^ܩ�8�m����e��U2ݡ][��<����䋘��eVkW�.h�kJ���d���S���i�Db��+ѹ\�U���QTm:�d5,�,�Z��;�F
�KK3�U�X���E-R�c�f*�V���*e�E�҅y�Zĳ�a�) ��`��O)���<:�z�2�j�]v�6��Z�9	zyڮ�]Ϻ��@m�U1t���]݇^nf��ξ���*���Pa�T!�R T B��f�e%�G�+͍���75c��ݟ�o��6�/�ܺ��Qb�=<\P�ߘb7.�69�V�v�O�x�K����9�;���ʳ<�_��k	/m��3�}g+ti�=�|i�f=�kZ�m��1+���$�Z��˧0�����Rd�rg1�
��;+�2���+���X�1�z�f�qb�������o=	/��h�����%��u9�X8T�[����R8��FPݕ�l:p/P�=�g��:�d0��s������Õ�r���[+�����1-M�23|��a��^�Lk�|�9�47�8��f5���s����y; �{���|�咏|C�0ᜋ�p�$(�+�� ʙ-&&Y�ֶ0�mi=49A]�,�RQ����Z�&YA˰�%ժ�>^�lu4U�q��>��Mʇ��O�!4��RW��=V��9�ǐ���0�yZj���K����m�|C�w�f����(V���'��ۦ��*�߽[�Q�
{{"��u���A�>� 3DX���|6�����Vx`˝�'��)P�(�հ��+x0��ԑ����uV+��$7Kb������:����f����߶���]���_^�:��Q����fj���~����mI��71���f��x����<���`�@HeT!�XaD~H��C�>���>���e�cu~��*�m�򤬓&�	G�Th4$�L���p��}<;6 �9�v�;6�Y)V0��B�_eD<�]��˽ۣ��x\ϱ$�uQ@x�<��@��o���h[k�J��1����f)�.>���6��"۽��fi��&c�f(���.�c�� �>�s"E94����ה����:iԏ�ۛ�e���8�$Ogow�T�lY���d�7�|\Z��H�<h�ي��]O�Zc���m�`L<*�q��)����?Ff��Y~c#<���<��"���bS�H��_O��S:e<��#X����LG'���\C��^]��-H�e�o�I��Y;��L�B��6��L9�;[V��+:K[��_��Ǡ"I��2���	X�2�N.E	(fu��:�W��.����"'����h�R5f�g\��nʹ`%8ͥ�ԋ�`�i��do$.�n�l[k�X??��D�;�C|�����,�qFm9&��$<����]ϐ����a��>�L�y2�2&�{;q&s�4q9��1D*
L�6e�p:m�L�e�mg�qA�a�z
�)|j��eٛMHէ�����I�݆ޓɞ�[��Oo�E�[SC����Մ�B�!��2kz�7���n�zL�ڂ�r����@�a�@!�BT�z�Hd�!�"O����r�u���0dϼ�����Z�!.Q��%H��32B@2ȖB�$����b���� > P!�w�A�F�:�?�D�b�)��|��B���>������EL�nv×G�����z2KH���M�&M�<�CS5ea�|�.Z7����g�k���Ng�#ٌ,�V`����W�N��\1���o���-���#d�xU�fD���TI��=����˥�]��z��=�-$�34���%�6��6��S"�b��j��:��ءo�6��F�P�o��&��"�m�Π8���I��}�c}������SKbT �x6>6=��k� ���i��E�UGy�\͵y�a�y�W�r�������1���H�}��}���ց�ңC�c��!t"&�8A#�m���z�����{��O+��t��k��3v��Md��T@���h��eY��3=f�W�f���O�����8�dL��E�f]ڳ�����_���;ꞕ]�*AVFw�.�)
��)P���co�����f�='`-�oW���\w<��ϙiP�W#tJ�=���`lL[�k` �*�?�1%�e�o������K^�I�:��n�XB�Z��d֚\�����n�D���������u�����]FmJZ�ˮ����7n33�2�ݝ��Y��:�z�\�(_򪾣�d�"�!�^�Dx2�C(rG�*n|�~{��ߝ��|\?����6c�`ǌO�w?�w�n{<,K�w�C�k�/-ꃳ�}�Ʉ�cƴ��BmWR%<�G����~nc��O3����mۘ�N��A����{�>vw��lE���j~0!IÂ����:$W�^M>� ��J"ݵ�M`��ǉ��=��;3�d��H+��ԩ��-ap/\��!cm�(�O�n5�li� ��P%���
�i����_|G��EG�s+�H�2㈘k��\yuV�ɱ]��GH�8;�Ņ�.�g�y�*���7�N�9Ҙ8�~�C�^�+�}�Sc�2$�.�Yq�#$�L���a&��9��O�of&,b��-�a�c�q�>29�(��I����[��2�Q��f����'��;�Gƃ�O8�BU��U���H�Y�H�	��oD���L�8�a-j�u*�U������>0y|��}�`؟��U��J�>����h��ɏ�P�>��ْf���yu'�w�^�Ã ;㜈�7�:�2�w�	]J����P$��������Ճ[������ݶ99K��iw4>H`׌ݨ8�f��N���4:Rq����B�{�E� ���$+b  ��%�h�E�Ո�}�t���AD�@ E\�R��y]�k.>�}�mZ����v�}������;3;��y(�lM.�%,�ѝ��'�����_
��e���� �0 C"D�@�#�|���{����<k��.�{���3��f��D��3ی�����������e��TU6沰�y���0�_��H��Ә��}�H����� T#-ɐ��9Zݯ�q��v�ƋK�,7����	>X��X���<��P���v�nؿ.ٍz��q,�4�Ί���sՊL�U����7Cz�8�4wAנ6`���,��ҟt�]J.�r�%�fu�� �?s��&�&���* 8��4�?k�!����a^�	�{��m���ۖ� &�;ur�T9;�qѐ�v+�+����ÛS�q�6c��=���w)K_\6gc����>O0�1m�E��!�p��9��!×�sb��W�-sv�DT�V�����ˆ7.��%�%�F`�^pΡ~��c�Kw5�����Bf7��]�aeJ��5b��g�-Q�|<cWEz�OHJ����AvcH�zF4��a2�$V�eމ�[���}�˷6����(�.Kj���O��a�"̆`oy��~��Q�u����ɘ�_�E1Pi��3K ��;�Ջs@d���
���<�P�8�W�w�����������;���}OT/]^��%;��7�j!mG����P�s�;,XN乌C���Q��&noY�?���}��HdV!�N�N �>��s��x9����>�T)��ʥ,"܂�����J�E1��hK���`0�^��������W�@�Oܨ�^��H��-���o��SB�>�mqup,��liwMt.C��V�Ώ�;�|,m"��!ȡ�Tǰ����޸��X*�p������+��\��r��TԊJ�ޫ�hm?��}����qS�)�3ɍ��`��xoAJ�i�H����6넴4p=>�=y�<l��-���m�jk���M}����Ug�M����[�.�cA	]Y������y�a�hפ�(��G˶�P�ʃp?Ztz���/FM`w�S~��a�)���,^1�58�Ǫ��;���qݡ���0uO����J���]`P�{3hw�T�.��?���,Y"�-m�Q��V��L;|鎍�O�����uY�:�t��)���� �ϘL��`�m����B�<S��dя��OD�['�������o#��ұ�� ��+hJD5�������M~���Sm�I�tJF\���O:�h޾F���3��j��d���\�mP��>�3�"�	{��c�[{$Yŧ6U�	$�7�to7O>����.{�2p����Lc}�Ǟ�oG�����������
?�0��d���paVS���*�@^r	X�f[�2�12
�R�׽��\el�	IKa3"\���
H\d⛇�vD���Dr�(�	�W�fe�H'�;�
c:sUr�]O�@��g���}w|pi��/��]J�C&�[Q�v��P�kl<��?V�*�xд=$�~u�w��|��Xj`f�͍�l�)�B
ͽ��ӵ˽��5�r�!O���.+rh�ϟ�*�{�`?�4N16HJ��N��}��mpw��Y�
�,�����*�g�7C�K�1����Ey��$T�}T��gZ�t�_ݘ����@���ï�Hk>BX��+>>�5�H���o0�3�8��������͙���;kt����ϛ�c@$߰&Z�8v~�ֆ�n�|���`�"R=]�N:]��>�x3�h�p�-��lL�*�,2����̉�����'�ӕ-�������`��rY�
	�/Q0<~�=�2��r'}0��Z���<F��yW�9���DQV�3)�a4	$���9�|����j�ݘ�G�5|W��M[����p�p���C��/�*��_g6R���𻶲w��}"��s�����X�!�S��A7T�	��4�YŘe�N��u߰\<�+6���#���es�i�Y�F6I�uՌβ�S��~+DI�+�#Q����D{�wv�.o-�#Y�aWh�;F�?gs�ف��o@�YPfd���h|n��l}߽�����n���U��pdR�!���(��x{�KxCwQ�s��k�~������J�H?}"R�_A�l|]!�brr*�%��P�[)���U.1���r�5��Oz�@�İ�W���Z�Fn�k�U?}"�������h�\f��'��f�l
��݋g��_��B����z����#�,��0��]��F�>N��3��5'%�iػ���(���p��'�|�	P�+��VT0�����5	ɬ$�qo����{����l�	�8��65r�v"�Y�	��^������ۣ���B�����C�f�=~	cߜ��?LH弶_����-|�=��y�v��5���wBi0@���p.��}���O�|���9a�Ly�3�go<�z�L��������d�m_�Q�>d *G�}��.3�i��y�Ev��	T��ov����~N(���pT�Z�
�d��Aj��j!��H@�kB���b��t�e?[0l�7�V=��0T�Zt�p}0���B��錑)|+�y����m���ؠm��O���W��Τ����'�'��R�<����H�A�_�p�>i���E��}p������+���#ڽ��ڤ�xwع��`�v��[���aqGd���^�.nʼ���-ȗC����b�}�D������Á�#�dXd������8�{�c �����%��z��c�Al��_ډ�[�La�vWyH�8=ό�,1��,�m���6�Ve3Zn#I���jC��~"Z�ܫ0��!�c�9��d�[�A_62��N��\�5��ތb��nZ���&B�|�V�l���v��v���Ѽ�T�	����q_�s�)��׭����m��u����}�<S���w?�]G:�Mw�	��Y�����HI�~��ﮅ|w�'���4��DF�l[���Oƪ|J����{������ �Y�61a�O��K�lu��u�e�ۆ���Mަ���F��{��i���
�Kq�5�'ɧ"�l��>=W"y�����{`0�2F^#*�}�jy�gU�F|+m�N��4E0�APi����;b���Ň�|ß�|3�ݱܨ=�l�u��F/�&0���J˕�Є�_�G��]�+��~"F�m/F��صj���1*�tݝ�����q^�������R)�k�L+��*�H�1���7�7筁[�4EvP��E��*��[��R���t��u�X0�����F�{�� �O�ٕ�B�^V��B!�^E9=ݥ0o��.1�.��V���y�#xa�G����1v2s8o"���֑�A�00$0�00� ���+{�Op�Q,-�bl�-�������?��;���\��G���.'�:5l��H_S��}���{X]��5w�Z䰇�:�Q>d5�;�糸1�1����eh����"�6�\�e&_A0o���'�EOT���8�^w���@�C��F2�`�`[?]{����m��q�D��bW��gB��!zA�
ٌm�Ⱥ��Ez�Q���o-q���G�A#�H�?y�=���aj�DZ43�Z]�g������;�f��{{�{"�p��z��D�1^zh��v��B�#h�.|���]�A����5��즒�U���?;``G^O�ئ�zـ"Q�k~�6%zP��� R�����"ƞ$�J�����L��_E9�Vϵ�4^��)�9��:�����ke݌jC� =�v��ЌKO�x�?��+�c��&	���m�2��u�t\g1�Μ�&4��7xF���ΰ�ۗ�s�/[;0NY"�yH]t*��ne�z���K/9���`�+"㷻;�i�����x�2�\�P�B�,��=��S)E6�[��9��m��N�h���h����̱Hz렮e;��%�y���E�rmf��x�{I�Ur͞��n�ev���`��g+$�S��9NB�4tnB��n��Wl^bڼ�X�8o�L҉��s$��Wy��Ue���$�YW+��m[�@Vp��wM|�&�R��jo�X��aB��� ����l|koBKR��6��Ԧ-^k�}[J�0��+�P#5u��ԓ���֧n��4�
��i�����ܗu�9�]��@��Y�ݺ��A^QRGY�'+L��4�M�Z;���N���O�!���8K�X�Z�nT�������FsQ��r���\�P�J�6���L"��u�u��u�u��ƴ��Xp�]�Ծ+�E}1��bL]�V��}pf$m�m�M���U��SS�ž�էw_f��0t�\<.��qm�:�9g2]'t�	��T=,P;�h�v#D�sqvN���R�2!��Sc}�Xã/���@,�Ǖ�3*m�$��3ij����:��Y�KzlT�x�V�(;n��N�A[�I0��(
l �a�o*�f��c�(t�B�\�&X�'f
�G�!���[�g��n�q���׆�4��ݬ�<��(K��AU�i�(_T-�ù�i����_.�`���)	 q��H6�B�TT)��?08cn���\;�dZ%��X�Wz�<5َ>��ۼ�tڽp�yWE���36.K6�f�8�{ܔ�tn
t��.�Z�/+�8=����Dp�h�nj�_H�w������q��;�p�ms�(��Q޼�H�c�$7�u:��]]s��v����:t�!"npЌ��f>�V\f�jW�����x��l��/A�&�L˹�!�Rx�!b!��ٌ��Y�L�b��Ps9�g#L.��HŪF��Ht"���n�mM6��3hό�2_[���`}�v����z��qK��R��˨��٩��f#�1�1�Ү�S]��26��R�m�׊`Y�`�NbJ���3wlS�dO_q�N�eK0)r���5.Zi�M��=#ƪAsJ�[��m��`��4��/�+��Nv�g9�pg_C�I6�)FMݮ�LY�\��i96(��z�:����Z��t�k�V�1����-��41�
X2�.�יMZ=�2��f��H����5ٖ��v:�`֞I� kO3z�
{�ol�&�<�ѐz�� &�.Z~������m��r^0e'5��%���7*hU��!㬪9eg ��%!4��&���vZ�e�o��¬kXV/�s����KD�\�s���������qǷ����׏%�ў��?��J�`���o��Fҕi̬�-S&I��j�����;�g�������=������Ye�џ�?�`��7��e����ؑDJ��
�� �*�~�$Ek�.��4�t�y?O�{|]}x���:zET���F��6�̩�PF��V�2Vfl6�!AԱQ{hSQZ�4�������=����������Ɩ���g��\�b*V��D�a�i�KmO6�ZU�s_�8|��?��^�qǷ����^3����T?Z����[F�r�(;i���D��J{a�����Me���ڈ3������y=�'���O��3�c>�~���6��i��sV�E

S_zv�i�b0Y�e.���h(��l�m�B��Qh�,V%s
���9u*��QD)�8�
j�U�'Z��]fλR�v��Q�q���U�Z5(�Qm�p����b�R��±�9'�X�4z��T�h"1TUE�fX�--������+����8�N�ku�^V����+s�{�;um���nuD�[�h�H1��]��"�>I�Y��jT9#���������WpRئ���m����3R��9��[�_����%p�Y��9od� �H�>7l^�D��n+[��7g��ݸV�׮���ͧuu��)vע���[������q����E;���S���S<�VC	"��R��)�UL2Ke4�̷^�7;mkm6�����w�ml��;g��v��;g�#� �@2JD�H����%"�H�2�@��>����g.o8L�-�fXm��*���nL�M)l��0���G���v9�c�� �E���@�q�_���BTA>�<� �W�46���rӟD6��1L��/�u�)�v�����{���}��5m{]%ƪ�n�X���=r$R���0�Ly���Ґ�����g����gj
P/N�A�H��3��>��/2i�/�!�����3�(j�,��JV�Wp��<���Zn����O�i�>f
/����k����;̄�?j�Z¶�:2�ݍ=��%�W[~V"��A-�~a�:�lׯwF �|��(�dG>���$�oH��ܞ����۩O�[!@��]�Z���_w���{H�q��	��e�ȣ h8����`d�x�rz������8g�[�j΍l�q�z�ϯ�RL�m�ЙA����^:�S������_Hv���/�[!#���U��y��Wz⎿�^���s//�T��)6�D7Q�=_OT0����dJ$܃��g�Hc�����Hޭ\� ��fpDl��W�~�>\��7 ���M�Q(ܲ�>5�ϙs��mNO+�]7��q���]�=�з�GS�̝c+��ކ�C[�Dr���d��n`�LZ�_B�x����oʐ�O_;ݝ�Gz��{�5��wlC!�Ǘ�P�Y�L�ۚ��n���N�`���ğ���"�%	�+�$y�yǘxy�� [G����
�m?w�z�jX(|\�>�A������ԧ���>w���]K�l7mR|�w���� ���k��d�@H�h׹�7~~-,G��S���f��fS�R�0䘿-*�f?0���x��X������@b�_~$�p �$gշ�^�>���{��l��������w�n8���p��~�Mip��N�Q���U(}�B�^s�2h�U�Yq�ݼI�F�}�v��3����X<���G��\�T>b�P�8���(��?U}U���˜��/���꾟r]7o����v�Wݴ���
)��ЮG1��N�5.8ː?=��	Ne�-�r5$�*�j/-�~�!�ժ�}X�=QR�G�|�l0�7�)j1��a{T�c����f�P1�������>e�\Y��;^,�k.E��pn�߸�����Λ�3��[�m���a�t�{fQ��俻�k�g�.��*�91�}HK�C���z	T
������_k��~���r�3�c� ssQa���!���C˜Wv��[Ϩ��¦5�����9����-�k�{Ҷ�@����h�au.�ov�.��`��]�Tv^&W��Anvq�8,�J&�5�.���};:Xr�p��7l�!�݂�T˂�=J�L�57\��t�)�1�! 0Xey!��!�Bg���|�g�����r)�&��]�4;�?�@f��_9h��*bzH1���c�n��E��L��ry���`'א���vn�1����u�����y�y�92����vv�5k�+�oGk��)��N�,���+?�D�@���[�D	~�P�_2<�H��g����t^�Ɨ��5��|`���H�Bu��3�^6ߡ���O�	>����P������jXl��
$�џ\���B��� ��|���)50i�!gA�>�Fy�!Ԏ�~���t{���K�*x��>�"hK���NJ��`�>d;3M?���<��Lg��L�����3�8O-.+%�_��֋ٚ��}!yo�c7hY���zh��Sfi	!�ի�<y��u?�.��w*.5/�����z�����H�ڍQ���tB~c�_ﶆ ��8}����+��Hkk��B��3��J���OXӵ���Or¸mD�j�na�S�nA+�1��mm�
���m�1C�z��ؼ�l��F��տ��*g����^�x�Qx�걿YѸ��/�@):�)�m�,�˪�5���A��  	������V.�zc�Z��S� Ě�����t$��z�R̛E�n+=P�o:P\���9��Xg[�E�ܟ�	�'$�� �
�H����ߞ�I�WG[;-q����Ռ"��O������b��C�ܧ��Pe�u-f��j���j���;�n஋k��CE?�ts��Ԕ�9����������nG]�k*��Cow�ݴ�.:��QGo	��ND�����S�7!��6~$Ɔ�MI�0Ȏ����������ȹ8^�M���1�2�Zxe��7X���ז��M Ae�I	���!��Ϩ$Y�;C�3�uB+#�z�����x#�߂��'|���`j-8�<	7%�=�Q�S{)�5u�a�$�n	����&zou���40o��U}��O�?������@k.�K�)�T(�K)�ʊ��3:X[����<З�2d��r�M�}�=�L%CT�)���G'MS��6NwI�1�v�v�a!���-������v�+C��_\��3n<b��e{�jG£P$i4�k����L���՞��ƗqMr���u�p�)�ξ��8�&̔b�|�c<�o�B���*�qwq!�d��+>+�d�Ǟ��}1��ց?�/�����@�<7Ƶ�N��ޝ�m��:֨,D�Ω�Z�M�E���Gs�
�>E�V���juꕗ���=(��z;���-�￿~�]�w�]�s�Xd!�$H$O Oؔ�?����M�~��IrT�a��$˝���^��x��CJ���1���{�睫z��w[���nS�2$CrL�֦��C
d8���'������Vk��[-b%�oH�����	��蘆��2�+;�*��=���t�思��w�X[*9M�`Y�o�%�Y���d������n��Œ܌�$�O꧆����{�Ny�_��W"j��	�v�����xk�Ԧ�����WJ�_���1s�퉣B���YJ�U��AvP�=��5���V~�f%�T�!��H��<NT�L���2ų���eZ�hܢNrlⲱ�s�C*��]%�w��$>#i��ur'��c��U�u=�M&�c^V�Xk�1,z��u�V�Ӧ�g��zy����p9���	��'΃|ou]\F��zw\�����Ag����[��;BQ�F�;�������;�?F�'pՊ�Q����I�&�Q(�'蕧�^�1z�|��~e��F�{a�>���.��j�gjՌ�x��|E������͆��l��D�v�c����u��A�X�#*�qj�5��t��Ȩ��Ƕ�u3N4'�}D��p(m-�-�<C+Ɲ���狳u'@
f获T��p;�i.��ۆ���';@�wb�ӎ�Bԩϟ6�R�R�q�:3.���ޫ���`!�N��+�>�y�wkC7��C���>z^S�T�ok��;�]=�������n:�dZ���\��Cvc\����Fx3�� �;���Ckr{i�^���c�}��xP9��v�xE��;pێ��U� ��T�hC7���酈|��33��|nl�ΆS^�Z��Ny��(���G��.|jzf�-|Q?FYL"߮t�2H�Y?q���Ǿ������O�H�ۉ�2`�A���]K����5�z�B<]2}��:2��w鸺ޛ��ힵ֞ۤ�i1mېU4X�7����t�8��1�X�6��H3F�A1=��՟}C�!�X�pJ�%����LO���W1?j�V�S�2{�z:g����nY]�|�B:�r������^D}���t/��,�t5�2Ж��5=]Ǉs�P���8�����)uv�$�=^hm�y�L�%�*�)�x`'���JI�L$�
��������Jnh��e���wjco��Rux��y�*��ӥ��5�����D�c��g|�n�b=��
�.�2�jR��o�j�o��Ω����^�7T'+:c�R������j�W��� ��G;�훺t�|Q�^p2u���e*�|c�uAޘ������q�t�����Z���[.q�fD���4�O� ��2�$0w>OnJA���{r�\������nG�p�*q�B��m��4Ɍzc�,�� �ݩU��^�]G�3�f���;C�����j���y���H�"�eW�Fh8傘��:˷�����l��p���z4���m��4�p�.sܤ����6��oT�/%��������VG��9�O��f�]�܈�0RS٨���<�[����>�IknU�t� �J+�}������3|��F��l�H��R[��):k�	�}̌Pu�T��)�a�c����zU?�OD�G����`��@�55	p��ij31z_:����^�Q��lw8ð%���y*���=��a�.@g���P�^��fceG����NG���<���z�VԎv`�+�ghV�����2'Z��6ʜ�".��r�I��i��_?�@P����C9啎0ɺg��8��HA�fEe��mv���71��N;pǷ}4��ˠEU���>�QT���C�x���fr~�)�<M���ԮS��Ĉ�wm`���F�ܤs$,����M	7iıU+ y��pG�yZ|D� �QY+oD�_a��/F_V,꒘�S�G5�t�q,y2���)Jnx+*��g,�mUt���[�v���^پ��y�{�����0�>G<g��<�����:u������{!H�7�ǛP,�)HU�%���fm
4F�J;#��ȵ���������_ڲ;銇�L&5��#��C��1��	q�vĩ�O��]�D�`M�j�&JH	�v`���8q�[;P�-�0!XΤޑ��!��;`kky��9_E*3��j�&��`%�l��-4��#]s�u30k�ҿ{$�J�I�*� N-*%�p��������C���S��ش����� �<�S5s�q��sL����uB�}�z~�Zy!$�0a���Ѧ�rm����Li���[޼�qk�<�[�c:��zΛ�/͈��0�֏1��|h_X@wA��'֮b�Ȍ��h�n�G�k�Wɢ߽��0��+��î����{��'�b�"�[���믅	�5���m��}�Wx�l��J�q�|c���	���
��ǒ�l��~"׽��{�ԗgμ;m����u^ׅ}./��9l��{�����c�^g�m7d�j���kq���o`;{���T�O�or/_
��7����)'�f�o��u��OK�$c�/��b�b��y��^��C9�2���r����a�$��z^=�t���Er��E5��r�����g���m���8���C�2N��!���@��a�
RjL�L����+�gZ��4�M����v��jj��i����M�Pm��PK�?�� (L��(��6#$��b�^���l�J�����25���� ��qٶ�5�-������Mi�̚>2W��J�8���qbا׵qt���5�Ru�n��us���Iƅ!�K�nQ�Y-��N5z�5���;���؜��c�Z?���o�R�#�׃������}����RZ(Ć�&M���m�8~�5Է�����|�J��IB#�|���R�h�z�ܦ:��o]�~�̑,<6���`p�l�p��N�6x���H���T\Ѿ��B�Mz�<�ʥD�r}7���lF�Ag�kkW�k�&�>*=-��h�Jی]);ڷ}n�9֚oCO?���כк)��5ְ��Z���v\ɺ�\rg8�����eNL�"HS"W6�`��
�{6�S��_|�/C�U	Y%֫�� �mɀg����Ƨ4fS@��~�}3����C.�WI�ѐ�E[FsЇ��@�VД⨳t9b�E���l]�W�[H}֝��m̷5JȚ�[`��Ҩ!�R��PY�Ec0Tf(w!����yj�=�u{��=�َշ��s����L�>�ֳ��N�
����R,��|K:�<<�g������̈́���7S��a��
s�?[�ܻ��S�E�a�;�ߔ�t����mr��?��{h����*&�����O��XC0=��᫝��Iֽs�Wt��+��g��;@J/�f�G��g0���mR͝�4ڶ-Ӕ�i��A?1�_No��1t�=�M�:e̠n������]���0E�"6OF��c�xXm`�2h�;�f�Cnz�D����[����zO��������f�V�0���x(ɏ�C_�<�
��S�E?6˄�X�
jc�(\c���2��nĔzFpٳ�#8܍$��a$l����#QS��*��BU��k�쿕�rN	Aa�P�2d�J[h"�>�^�c�.u������Ƹ"p�R�~"ZϐC�|��+o��~�5�ۻ����3�1��
[b�ӎS��/�3������+�	�,��Nh�v��6����n"���K�窸f� Z�b���4pD��튘.P&m�[RL֙)5�7N�	��sO2Hfc��Z����4\z�]��6�0-�w1�b @:�^J�|߯v7�N6�I������J}���8�Ѻ�.:�t]������tpC�pN���]��z}�gn�z�v�-t$�S�̥�>�0.Y�̈́�:��#�qU���dFٹ�k͖ظ�r��w@	�����/q��s��I��@b�;�SJ��O9�v���R��x!���n����Ϲq�ϥ��ξ<e�*��2L��,d���mf���%Jo�2����H��ٺ�)<Bu1��O�!�#�Ɖ+M�zV��
9V-��RG[�8G�5��̧��vVά� �!�b�tv�4���� u���f��xy(��԰��,h���l(t@e�VY�(�W:uk�D![����ef�`�4�y�d��2|����0�h��p�S���H�`{� ׎�$ú�}D��;�/��ݓ,����#��M�wsx�Z�պ����R�[�.�7 <�wv�����R�����t䬬۳�(��ۭ
 KL�,���֒;7:s�3c���5�[��U)����|�h�5�e�w7iE$�&��e���Z��"�cQ�kV�:uG��XO�<��2lq��u_��>������vq�U�|T��9l*��=c�Q�ኙ����߲N��В�n��:j��v���-��7b��&�.���*X�H�?H�	t��bU0+r]�����ƊH��D�*\=s�Yzn�@��'��C���\�2��S)�Ȳ4�(��2���t�8��@�vz��B���Q6T�e�;��J��$'�ȕQL�ژں溷�1�P&�̄�0vFBy(a�u:ȣ�����g,ͷ��� ���5�r,�Ǣ�Q�GQ�45�m�]�d����V�<�^�D���ӷy1_S�,7�Y�k%t���:N��������}*TB+96Q�T��
�Q����Oq7�����&���L8&��)*QrK�֓��cЕ@��[��gg -����G[�S	87mFKΤ�E�#�!V\����C�Z�N�u-��+]qn���N�ifP\Pf�:v�V���}}�bz�{ۙ��J,�ޡ��o�kO5�ky/��[�v��[D��:<��\�-��wgk�4�������#,X!�Q怍�"�;��n�ڡ���6s6�����,��1fm���-�Łq�����g�:܁�A8�'�3]bѣ���xG
H���&1���R]<:��% �s��*j��(:�|�t�����Yo��T�Wk�Z����܆Wnn��)���]�LηS�T����\��˥�]D%ö�+-fo�w��/��"(�'��h�S�j"&��h���1JkFT��g%Q�3�Ѱe�:t�<�O�|�����>�g�;�SG����IU�,kU��j,Q�����[UNj*��:i����y?�8��_Y��?Y�=�ٮ4SY¢fEV*�Ov��b-��vu��d��"��X�	�"�g��ק����{}Y��ϱ��}}5�?dl3�TH���EAEDFsDS�ȫ�*�U
�D*Qi�����y?O�㏣����~��Pk'	(�9��"�QAEP��'�TC%bx�]�S �u0��Eb���wo:g���׷���q�>:ϲϲ�OUTQ?{j+DM��U~�F*��,<����{�L~��|g:&�[!f�O����v�>���>�ϠzK^��6�ET[����_�|1�j7�\UQ+(+5��n�sF#B���s*1Eam���*���[
���)cJ�QRu��M���*���X�K(�Bm-�E�oz���#ıE9-�X�j�>i���`�b?)X�����m�����I�d�r�Os-�bނ�w����6\��]��I۾�{�7O�u�s�?C0������"�_ކ�����uE9����to�"E����
��SN*i�g>���gE?�*|\��z#�3��mR���M�`$���]���Qr)�����	�Z��4����g!� 2�S-��(Vr^�����3���^���1�;���u�U���b�.�Kh�n��y�� �@��L���o՘��6�4�g}hzl����e�w��p�7Rĉa s~|�i�5�0G|�����Z��ggN7�:������Q9��c���a&/���Z��77_�9�*3ͬo�K����ˁ<�R��<nF&Y�0��;{ʹ�>�)���{aSэ"	�h݇g�p@��/��o$��ِܚ]�m���v��>�~Im������|`��+k�6��>S8b�ym����C2���������7`ǘǰ,�l��p��Y=�U|��)p�����ZY������H�i�=Yh���ը���b�f:���~^:��cҝo�Jz=L�V���3!{$!��	��?`S{J&w��f�w_ln��}.��e��w(�OR��\�{���*��̴�=]F��7�F�����Jy�D�Y*Д��V�3��d'u��_��6G��~���W��� ���wOt�G���;�@��Z�p6E�z\ �֒��2f,k�����w�{�K�fƞ��z�݀f�㎀�n��Ԡ[k��5�<�|�8Pc���&8����ǋ����w��J a�H<Ϳ�`�QQ?+� H^?z0C'.;�����>g��i���/�{������Y�`;"%����;�{�$c6�^���"a�@�8~�xU$dR�AU�ﾛ�)6n�7K�h�7LT?a�6�w�B��0���36��@Q����S�L�3�&�m3w�靣m�jA�7����6ПK��7���5B]���C��Ln�L{R��o�L8����<6�5yR'�}^1#=rڑ<F �	%R]3�eV���S���Q��pw��T6�0W�Z��]�<��,�n2�%�K�f�;
]c�����}̞�h�Q�ݿAza���h�>��>���p�/a���=V�W>d"[�l���GV�s�n�Q������`YG��LLo=���xǙ}���9|�}�����>��r�c �Nu��fO��J��蝗X'
��z��	�ܾ�����ܾEg*5m��V>J�WtK�|������_vT#�^,�/9�:v�����+WB8fs��".�k#��ܺ��4;������%�R���@B2$bFV��"Hw��U�����hL�-����5k�,4�|p��㻷7N����b�ە���{��(���H��)w�w�>����"s���O)j̟����$,49x���_a��+�"�/qb��vy0���)�]GG���K��:��@vĽMe�;�5�<��X(\�k_��]7�<!"�_���H�������ܨ6�.���rͮ���ϭ�4��=uXΞ���B,�g:��O�-H^��)���\�	O�f4M�X�f���ޓ+)��w`��>`3_��8U@=	yn>WJ彫�|՞3)=��)JF5��k*�5P�Ms��:�'`�㘲׾�a��:k�揌��ᐱ�8��'�c��ٚZ�����x��D��s��|
IHU/��@��O=�MϬ$���7�����mvGd^1'���q�({��c�>��#\�3ʊ���`N}
l����l�J�[��=�jNڧ��m���gqZ�[MJ�O�~��x���K�`Q��Nku���*�5����u�7��$e�[bx�W
&3�"E�2��˳i��n��f�X��k�~U�Ա<�b�˺W��ˁ���l)tU�E*o�rd,Yr���f܉��m�RٖN
|t3UWhX2�#��@�'�s��
ɧsL�;�t�Eݲܧ:f��=]/�" ��\��R��[�|������s��~}���C.OR!��E'}�y�y��뾿/<l;~��&Q�OTS�]6=>����`�;#�� a�i�o�U�w�l���� 5D��WQ�HVg�La�5J�u�#u޽7�kr"FP	�i��lu�ɽ�N�7���ΩƆ�{���_��c�d��˭�U�!8��9��4����2wj�5sD/b��+�rݔ����[����y�빙ݓv]f,�g��sRs����q�#ڻH���=�]���6��� ���A��>�}���<���fR ���TĈ�N��ٳ�{	����םv-�� ʩͭ�S�d2{�)�W\����C��Y+�|_ٜ��F����כ���[N�w��0g|z 3��~z�p�w\ӊ�3�ת-̶68m�r�g7!�et?�hf^�������>�.ܦ�Tr�C�Ҭu�j��˶����=�����_�>t�)l�t�H-A��G-E�{�K��v�M[6���i���N��s���s�<	܁�l3u�Yu�q��dͩ���F�y[��]r��p�����ã{�O���|��{ ~���)P
B���R0+7y����(\��ᜰ��'�szcH�2�bQ|�O���-�빿��H�Sw�Ͻ>]����o�+ש���/�yƠl���+��T���ɜ�V�L�|���b�3�8kQ�a۾ח*�����K�#cy\������f�xɞ�f=SQ88���zK^M	���}�}��7e��>��2��-GO{�~��]:>���55��&�j��=Ӌ<�v3��'X��'6�M�kL.������OR_T�p�wZ�Ώ3z/)2�����A�j05$��E�wSU�@�1��7��cO�wkO�~F�K�VMe
����QIuT��x�[v�XBCX6�_��5&���:=�DM��^�]\��њ�W��{;;2�)��/;5�߭�������LO�.��_���=Z�g��S
~���z>i	�<x�.FRy��6���2��-�����5��E]�:<0s���[���ed�{6{X̃�Q�Mz�%D{�`H���Ӱ��P�����T;�T�5k6]�8�\1�v��⮵х��ѭ�]e��[۷b��%��U�~�~0���Ǝ�2�!��OcA�W�ԣ�յ��{���}	?����?^�Q�ϣuF�X`��y���H�m���sd��i����w�Q�_��͝6�HN���`�C���b��4�}�!eO�}a��8��'���[���U�3:͍�1�D�*d��&*�oI��9�`P*O��Jʡ�k�g�?->��uZ�q�.KU+�T�oMV����N^.�y@��OW�2����=�����/���UP}#��9�^V'S{n��\m%f�B��aŹ�|���
5\@�S'�7�rgu�(wޡ��s�!��YL��	w�V"�W����Ӊ-�S�k��Õ*;�U�;�x ���@u���ǲZ�K��5�u��ioy�o�%��Kf�$_� �xe��VKp��߈�~Ƨ��YėjT_C1������e�=uz�*{��&b�zvQ�E��φ�5okΉ9̺�SL>�V�oow�Ś{����res@�W�L�����]�����8<��F��"��o�}N������G�F$H� ��P��(B�q�2&SR[RBS2����h߹��)E�٘�FPm��J-�][q��ۻu�\T�@Kd��73��z}T0'�X1��b(	v�a��2�����ռ��Mdf��h2=/|���x�L��(X�>]wM".2�-֫�G&�ეxc��|\��`N�j+��x����fbDOf6d���(���k� 3�fk5�e�q��뽳xQ�s'[ML<�L�ލ��Rc{�8�uufy+�I��ސ�)ὢ��8|�+G\g����A����u��Vn�]ˉ���G4{rO�v�]�"�>�M�f�Ɩ=}}�މ���w}@v����2<����\&�8l����e�~5w�f��lef��j*����{��-��u��� � ���A5����u�p��ɛ�2詒m#3?E�p�(߸HoT�t=�#;�wM@O\�^ճ�8gV,�����c�cs��X.��K%C���-Z�/e�_��<�V�=pd=^!��ʝ��v!M�x�Ǭ)W�V�J��ٙoFȲ����Vȼ
�S#H:B�}W6]������˖�B�q���)���[1��חc��hs�ݞ8�T�+u���1�O��ә����[���F�-�\޾*f�#z��.}�@|�0:�n�>��mMgT �f��J�Mӣ0�h��v��ˊ���/���( |v���(1�,3��O�N+�ν����^:��G��ͥ�rP�Av�9���Ƚ���׫�w��]�`g�.�8�\E@��`N�m�s;��q"��;��h�g��+�����}�S�!�v(����O�k.�>�R�g�T��2MH����v���`n1�����rws1��7���2�����E���~����߳,�����cP��t���<�j�	�����-n�5�OQ�'��u�Vv�����UA�ٹf������>4�{�3�)G-�J�k�$o[܂�R��d�������7�,�M��X<m��3Dv�I>�x�����z�Nr��<�W�	*����
h�*��0E6��i��iGc 4�b�(��@E�s�]������L���[�����2�M+H4
*����n�'ˑ����n��חZǔ
���9��=y]��A�D����P0+�d�k�x̀��� <����<��O:Y(��7O�N�|:�&��������=��VrZ���˪�M����Lɛ"CQ��ٳѴ�ݛ'���Ϡ��3��7Ov[7�^m���n}����"!r���}Zo}a���p�"f�oNT��,3�d���f?��S��+{pJfϽ����ϖA ~�?$�D�(�A�;��-�?��a�i����0�4ɑg՞�����4��1"�Ke�n*~S(8Ħ�-4叿�T@<	�f�.��ˡ\�n��&�h�H��츽�iH��� 6��/y됨��"���ɓo���k���*9y�3@_H�]��z��UR���v�oL<�<��ø�v���O�S�G���sW�K��QdFO��+�f���S��ʻ���X�'�7�Qn��ϟa�K��i�7�<k�hLxݞdHư�ʧMͬ5�Q���W�������AHn��k�ۥ�6V���D0���M�G�j����dl8n�/�Yi�uv.�Ӫ^�\�W��wW,�{z���4�\�͵��ģ��� y�y� a��^l��!;�p=Q�W�|��*�3�gk�o��� �X��e�uWx���g:�r󜺔�2&-�%*�]J��<=�A��:&�@և��3F��oi�O��(蘈���p���mY�Q�=ְ��w	U��1��� Z�׼��]_�����\���%�_�V�v��=&;2�Ӱ����5���їt�m��W�h� r���ِ���{���lӭ2�]��n��D��wl������xe�}
���
Q��ߵ�l�����Wv��3� �X�`�T�7�c?�ҹ�fsC^lQW�;݊a���zUf�-����^*|N�ƭ���p2M��9����qӄ0����c�}�<���/�/f���ZuZ^�'����o{&q�Nw6{���[��Fj�@Yۭ�10��׽��<7����U�����c�y����~]Rۨ�]K՜��p���n��U[:����L��k{0�jܡ�KtX��ڙZ޷|+���ƈ���NL���޽��7ƴֵ&$+jW]�=Uttz�lwČ����.偱v�=��^���5��@}/����1��4�� �,��ܰ^mdj�R:%['O�1׷�����X�nS�죇R�1M��1�#��LfJ(ܹ���_εIDt�������o;7\����S�@9zZ�g^���8�>����h\`�#�.v1u-Ɠ��u�i��L��zw=ԁu��]�:���dؙ}�hŘ� o6N��wY��㰻=��C�E�>5%�a��OE�pn<�4�]�J1�֋����ѹuu�u��j)����r ����Y�6��]*ˮe���^�p�b�1����s�u�ۨ�!�l��̓iKP>Ѣ�Q��N���1N���i�_����Y]�gt2�\zd�l_B��V;MC�X���]�BR����d�e���)�7t')Z�7n�Aܒ��Ǉs��;��6��3(v���A��gR�N�L��ܫR'�3&u\U�۩�ua�n�m0}���A4-��t� '��r�U˖�n����j피E�Äc<�_4��Ij�]���8X]��S�'����s��4J0W;�v�qۮ�56��;��n:�и<�I�*����+��k�㎺;xu��ᾦ*S;�lQ�˕}�v�l	���Z-Ek[�֬|鬴�j�)�j}���Q�Ӵ�vs��LPЛ��˼3��P��
�J��b�7��Ơy����6�2���=�uf�:���|��`�1Ndm�AΥZMe-�̺����W�<Ol�
b�7CI�a�-TŰ��d���L���e>��m�Տs)��E.$��l�R�Ti���W�/<��%*Aȅq4��Iz[�9�|v�ٕ�nj��(P�F��٦Q�&���ո_\*�qqtN��F��� ׽��W+�\D��Q�j�;W6�5�����ts9j�K�\#��JT�J��;�	���J�7��˨�������sM� x�&n��K�f��;��O�\�ɫ{L��_���k��r�e�$�N�K{w�U��ty\�S��:�0�2�qn]9�Y[Ɲn�m�nK���%M�W2�92s���o^/I�k50ѭ��R5�^_v��X��t�E�c���bD*�r�o-����c�v�zM����z���!ca^���`)�[�a`��A���	]u�mY�4JT���}>��������ϔ+6�-�ZQYmk(�mAUV}I���r�ǧ�Ƿ��������3둟��>���U��jE����(��(�,�U�G"�"*����G �?\{{{{|q�������~�Q0DEE�UQBĂ,�U��PGR��k\��(�8����oooo�8�>����:l{As�c���3DDE+����EK�)mj�������k_:�J��:i��ӧO�o����>��n�z�z��r�ϟ"6��e�U���Z(���U�QSP�ΞΝ:t����_Y�\g}
�>|���4�ڙ
d%�kQU�Rڹ*֎k���:*�gO'N�:t�{}~���Ϯ3���8�EU4"��**�XҔ�Qb����eUU�Y!m_�QTl��
)�I�iETU��J,QE��i�UT��eF�*�o��-4II4�1p#�T�"���%b�� �'�AQ�"[b�m���#F�QU��PDQ�^~e�ҝ�T�\�ݩ���rk׬�㝶��׋�{���Q��添m�*PH"�e"K3*T��2�&e3����&Q��ҕ�80oj�j�����I*����M�a�vD��+L�nq��X<M(k��W�g���[Kӧ%�������\��9�u�K�l��ۆ݋�r�[��{�m�\�a�{Sn��z���b�^:�崽�����ښ�]�+u9�Ki�:���i{r�Ƽ�qR�ۯNޓԁ�'c��[�D۳��m�!�,L��̞���GZp����\�^���i���qcy���a�kg����g��x�o��%fZ��rR~��͌�Z��|�^�\E
��� à<�NEm�d�2���u�8���霦�!���C�,0�#8.n^b������ᄷ+��xh#yV}�^L�C>�R�>�l\^���Dվ�c�}��=�,��&y��,.��4����s�[�U+��~��i1��v�^��S�>�A�F���}>M>�bS2��j2� 1%��0��*�l1���Ǧx�C�X@K<����ȸ�髸�t	�Ū�s/����0�Y���V���VdP����Nڽ�/y�T�oDܭڮEܵˠ0a�>q�گ���O�dx2v����Lz�Y�ٝ���|=���:U?����0%�Ǘ����.bm�}\����h5�k�������~�"���הbPl�k�kw��9LD4hԠͣD �6��˲]-�7j1�n�;���\��.�{����̛�[���I3�T�ަ{�	g2�q&u����O��yP^�y�C��IZ;3�+׋�Vh�].�us[v��DD�N)��:cS	�V_�%.��l�*';��N4jgL��Ȥw_�ggQ�jǎ��lZ�Fv����3�#�q�'�Us��ke,��*Q�17�;��ͦ�9��W0�1��W
w`��7۸q�Q������7�ٕͥ�q��2ʇ�}�ɪ�4���NN��+�0\a�w�����e��c��F�P#��nut국۸o/o�M��s�X+(�Y��kSܶ�_���U��f����v3�k����f��?�%�J/��Ů�e,��Gz���EF���  >�},~�&O���M���P)+�A�a�7�ڏ�ϐy[��Xұ�όՉB��`�<`藢�W��uZ�iN����l��~���v���`�{*�˶����U�����TU�t�K"
��w&~�^�rƗr{��f�����㤣�٠k:�m��뫅v�Z�_����_�,Px���)O�Q B��}�B�i�=�1pl��_>�%mWMͳ5��Q����r}�6�ʵ*Pܺ��lL�n�����C� z�x���.��:��R]^ۼ����?�����R;�S�:���FŠ�n�]s�ѹ�4�u�חcշn ͊k)��������\�A܋�or��i.�m{6���ٻ>ԯ���M�T;�5J'���h�zB�v����=S��i�@���r���մّ����S���e��x�[}�Ʋ����h�Q9�<���'�	�,�I��͙��7�퓕���X�4eߜ=��y�6z;�E�G�����X&�z_M���g(�w���:um+�[�3�-3���ö/�j.`���7H
P�OS� 1.'�CKd�8��m1��˶	���<a-w�Nz�9�v�z�bsL�9d�rvvwacXط��xi�Y���ϪR����SVT�N��<T�j�i�"�n@��e^cP��v���÷ y�4����7�V�T�JZƺy��7�V�=6*�ʼ�����B�)��}��moI:A}�]�xl}x�,TiY0s\�'�J��P�.�+Y�'ٳ�b���d�a�f�X7�Kܢ�T|����d�-��\5�܀-�3C�>"�����	��n�y�!~�t��v����T�^�٠!%������}WTK�Z���Ihga����9vj�AK\Y���k����(޻�ɑU�]Tғ�M�Ŏ��ཋ�*��Q}����0m�fk�����e��r6y� c%!vN�� T� �
�9r,s�1�S�y���7���3\��j N̿^�mR�L�<��gdW><Dߎ�t+����=����:���&��O,֭@7 �MG����	��Vg��vWjyx��2��\"vo
8��=���F7�n���L�ؽ����;+C����=��s=;�5�a|�����/�2Mf7�>5���;����(���;$������%�V�����ur�yv���f���oj�&>���+��+t�ǵ&����vج�Ι�iրB����ҙ�j2���ޭ����:��{�7�֚P�yr��;;r#��~���\)*\:������iof�E�9nAJ�i�sƋ�D��"	���@�`ʔ���2���u�M�V�{$����NK(mcQ��q��rqNnhv���A��{~U0*�N�t��4ڠ,��'�$3�V�	�]�ҷ_z�t�����C�Jg8��՞/���<x�(Y���'oͭc��������-v[ަ����o�V6�)�����|���W������f���+�>�ڼS��Ɲ��7���*v�k"�9��}�W�`8��/\.�T^�����+�6�}�Duf�23m6yh��n��k2�� 2O4�DY앱*��<*�9�&;������̊��@ϙ��Q���m�ϐ��ɇ��̃C*t�OG^/��q�kM�����T�v٨B�6)��7����8P	�A�D�W�6H�������j��3���rb��T�۴>yJ��#1y�%�� m���%U{0m�)+㾺�C���e��&fI����!��^�}�]�s0kAyzl�yǪ�=��~o�k����D�"�Ъ�f��U��f����[��ecʳ́CT1h�/:N0�7Љsk8L�I}sM���7GrK|��eU�D� " �z��U<�f����nY���47K��Ϩ����?��X��D�ÿAf�d���]�ޯ<�g39�v�����̉�[�,؍ߪ;"�SÈ<�vE(���E�Otu��.���%���^%Ujb�k�;�y��*��NPod.T�!n`��S��U�q���ԍZd�wv��|��{-��&6s�}e%d�o�ʼt�� @��v{9�<C�d��}���9�Vc�:x1�U�'�]�O��}����.������s+1ev�L/TKS�gC���F.�������F���7�;��Dg�z\�2j��0V�@��IQgn[�!���2��g��SMn����֍��P3�0�఩��`-���5�t�|�S7�棖�[���t�R2�}ǻ�\(�y��9 (�K!19Ew���3�f�<bA��
jl�r����kr�̵J^��W���ZK����yyH3=�U�:NK�C����+���z���
9�ފ`���܏^,��5��Äɢ�ٗ}�+���z�dݜ�5Y�[0�{4gt���o�<k(ԝ4�8>nߪR�/���U�eX����>5�ͷ3]og�������+�l�`��F���=y5[��2R��G]GKS�]��G�*�էWR�j��K�Y`d��)�}��G����˳_z".;g��Q4���e@�X.�6Z�U=+�"�r8�]�4��	ݛ�����p)��`9�Z!���&������ը{�y��n�Sפ���\��I&ܽ�w�����Z�ޏ�sѪEl���|��o���ˍn�˺���w+i⛭�6:f�-��Kn�A2��䪠�ч��ץE�+cL���KG���f^�Q޿s{piJT�mwo����3�n�35hՆP���;l}�=��?��	:@�����o 8��������n�T�H<�"z�5�g�G�Wy��a��=��U���n��@��]���T�󊂯�2i�\�����2{ݼ�}�H�C�	��!v�:j}���0�B��3�R�{��o^˰\�l�y�W,���z��:��4�ꘕ��+�u ��jʵwøH�����<> F�"B�^v䢯 �Z�ݻ���S��`�y����i���#�	�]�9!�n:�D�c�)O(jS G�吥�^���'4���!f�D?1Ƽ6��x�ܘ�?�z���)��-I��-Bi�A0oV�S�,��Fb�;96L�N6AT��0*�6�����]�}!cα���~��0W'��s[�*�o7�wB< ��O�Rk~�@�a��p��n�{�X>Ʈ�T�څ���]cQ��j�^����Z�C�fQD^���kY���ߤ#�:w���<o#P�Gg��i��"1����=��D�����@��ê��Z���A�<wʵ[m�X�6d��.�=/��%vb&�'7��+�uD��߉�4{&�;ߵ ڛu�_��WE�'��Zq�fbeQ�|�Sq�/q�$��	H���~K;���>��m��ىl�Zz�c =Y���!��;h2�����ھ�԰�tH���JT��Z�2��Kem��[��?j�o1�]��VЬ��L�QI\�ӥ7��m�C��j��kP�b����gPQ-��r��u�O�lǎ=�5�v������>d@��2(,OA�!4%Ē)L�
Tڝ�]�k��-�e��)2� ���)�-Z�����#�ڦ7m�����o=��m��{�^��F��f�R��h:0Đa��lcoIX���o�w[ܜ�$_z�E��l�4��ƬoYMg0 ͜l�=<��L��L8���=�i�6����3��_3uS��馉��6T��2���!���-{�Α�݃���������j~|g��Ժ*e�ũ��dE�j��*�:k�ϡtm���5YY>'}� 3�����o���b_�譧ܤc�^8kY�;]н��H��n���Ƭ%q��t-��޺���ۊ����s��{03����"-jQY�/�=��~��8��uw; �8�ek�O�<ݗB��e�j稞S�������^n�;Ct�ՔI'�[.L�J����~������x[x�t��+�$��ْ	O���86���&�/Lep`���̂z��"��pV��{��?evC�.;N�
�ѣ �mf�D@x��;�a��V6�̺-�l���e�s��K�^��v�����ڝ[��`���u�Ӊ|���X��Jw%��Y\6{�
�@�Ƕ)&�X-��o���w}����ӎ����\�]p�5�8R�-����	���o����O	}˷�[�z�BT�^\���Gcwr����r���!~�� ?>D�aEu�gd0f��5�OpoPZ �_�{�}�����0(������ݬ�>Es	��6�"+��u�wJ1�](��P-fN7>���f^����Vܮ�o�^�d�]'W�hF�vv���z���[o��d^6Na��C�ɢ�U�G���K h8wfq�_:���ve�@u��u=u�w�	�?������3�9��7���ݞ�u��B�wf�z�rR8��+���V58�N#f�a�������v{:��6�e`f9�M��nܜ���m�7�54�kO�ݎ�A����5ː��1��\CL۰1z���w����}F�_w��:�3�7iԵ��Η��б؇v����Ą&I��;��1J�E��S1闅�*!|MnU��E�˴��!�l`���E�Vf�0.� ��IqԧK�W�gei��N�;�a	���djc��rxy���g��[�����9��5�X�x4�2dT	��(��;�*�%5�J�G��l���������Fj:P�*Ӝ#�LT�d�y�_h��ʼԁ�6�Z��i�)���㙍r�3����2�N�-�g8�B�7G�S&lv�X�.��B��<�ܮ�1;D.:��:r����{$���٫���g 7/pv�RW#䁣�'Sk33��KQ(�v�,��c<CG_,Vb�f�ؒ�1�z��#gq�(n�������T�sXz��Ծ�^�;��k�U�Y�f��A��۾T+/Edz�S we��rnﰢ��o�h����`�*ֺ�3p�Ǽ��1K�ܥ�wgu\�Z�dN�b���s6d$����s:/VF�fnGs�@��"�L��Ք^i����2eu7���B��c#�-`Ⱥ��;��9�;��*�*�>Q��� m(h8��:�o�݂R�s��8VCĹ���k}0�{�n��W.�(�P��B��Q$�
�]e$M^����usSI�}MWu뵺,���哨�G�R_ ��vݚ��8.��!2��GY�lsgQ�B�3O���n��fV���S@���jMD�Y}�患��z�I�۹���յ��P�.�1�%�O1N��&����U�9ˎ;�=�4紷]��Nޙ����(w#*��)��t��|�s�8��g>Օ�^��:w��Yz��[cv�ԆӠ!��4Y8^uS�N���N�nᙷ��]N�[Ot]��l�w�k�K��O;����RK�fڭ� ��U�:�[-��o �
��V}�)M0D��T� =ޗ#xwA�޽�����X=
�Bz���Mԙ��,��c����X�n�4��\�m١k���]�9>�ז�u�437��N+���\�z\C�#��[��ˏv��6�k����8�r�\i�����«mP��.��;YL�7���](��g��D�YOv���N�:u���¯���K�lb@Mz�u�����)�ML�Ѣ�n͹����]�(��q�"i�f).�q{g	�j�u?5 ��#ܬ�����a�wʖc��u�d�g��Ra��7ï�"M��\-�$�����8p璪b�Ա�*>ɡ_Nk��(9���f��j�U(1��Q���	$逭N	ٷY�,WQ���d2��*���3'6{Z�?XI0DUE�[��"��[F
�'5���J�TQ�========��G_Y�^���(Q�X��)�Z�m�F
��mW��T5�����3�������ӯ�������N���TQUL���q������k�+U`��$e���====?__���3��>�%E#W�V������Q,_-5[l��g��N�:}��I���gl��Ow
�����K�ɽ�j�S�h���V	�(��~>��====?__G_Y�^���y�UTTV'��J�ұ-�>2�
���U�� "��Qj�Dm���*$�� �<�g��===>>���>������\�\�d��b[�+�J�E檞P��{(��E���+V(�E����+)EQX�3��Ub�fq��>���byW�U�[�V1_��:�^��L��
��V/5��Ȫ(��2_�	-EY�C*b�kV�"�,���D�EATO&�g�^�wb=�g��8u#|d��ז�p{�<�P�НM���X�ޫC��wn֓~H�	H�s�9(���쉿eh���jȍ�v��xI�+Xd��0�oN9�5��h	3 ���Sr}�޹m-e���ph�<�uVT���Q�Da���}C�~[bQN-�,s1#a@l��F�x�eq2�]7{�*��`�h:�҄�����F��;�-9W�뿯*ӏ���9 �H'�y���T-R,_z�b�,9Ƅ1'�z�*�+��0�V�U4�ݵ �@b�d,鉯]�����8�P:}�J(��7��vm���v�4�#Ft��7KQ�6`OO��l&y~�rry����n�}�����*��H	�}�T��H�^��i�*�����9G{Pp��Q��vM�;���v;����z�F\d�=�w�kXK�M���=W�����}V+[Ҥ�{�-u�^�ڈN��/ٛ����	�ɤǷ��ܷ9s�g[�;����K�]\�.���c��ʚ��;�k�RC��'����r�s����رd�1�U�u���Ô�Z�3i�k����O�.ј:/e���Ė�y�v�>����������Aæ�/p�����Z*��f:Ĩtᔫ���C�k��&�#FM��a���@d.'V��nx�g��FƧg��X����.��a�."�����CJ�gݙ�o��:ș;�ly�?�&�O��`�a�m�=La�e��b������j{!�35�ۮ���֦�pU�z����f�l;�NW��,�1eH-3���T�W�!'��{�e�p�P�-������٢𪸿���MO���D ՛�\�;��������ٹ0��Fa��>�Xf@�.3�BWz6�����>�9��5@�c�8U^7i@Χͣ/_�� �F���DeTq���������!Pi� �r��1/}��`=_>�v��쪵,}��/$��E_A7v=�/���X�}z3�z����Mu���ͽ���~�k�.��.��W���s�8h.9W��y�I���f��"�+�-�::�vV����8T���	]���͏x����3;���F��nwn�h�l�H!��}X��L�s������;Y����D�Q{&��zM�2RD�g�!�D D C��4�9,�be�2̄��}����q�-���F�D��m�$��:�&�էӪW��mn��52�2E�)�U��c;C��;��P���)5�v�h;[@)��[lԫ��k�T�jg�,���d�5��K�Huߛ���4w�?=�ջ��ߪ�;}c�M���ԓ�'}���>���o6_ykV0�oh��3�{�c"����<G�m��Jh���o�}�W��`�gz$^1"�%�v���Vù������f�s4e��ۍ;�ժ���F$�T�5�^����DI�ճ��@�A�.�����U�g�ve2O�ny�d�_��6�K��\��d�S�.�O""�7{���� �=Ӝ\O��.���dV�R��/w5�;u������H�I���������~��N�q��o�k$�!1-SP�U4-g1n�	�	;v�3��2�÷����ʟ��+��Y���q��)QL��Z0���J�0�m�5� �j،���9,'qa�,IӬ�}�1
�.K��N�������Ig�g-$iõק��w9(�+���I$�9�W��3eu
����%9x�Eˬ��3��?D#�0�^h�v��и4u{E�\�=����k�oWn*�������7��=��R�B�@'40lV=�p��|��qVp]���zNt�[�FNjUHk�s���p=�_A�J�E V�Ǿ�z(;y���Q�1\�M��)�X]���M멐6��`EϖE�=�'�������В��op�=5,.j@F�'��W���pRƚ�(�S}����$�}���]�.�<q���j�>8���m��k�l&+RL�l�	h��c"����H_`����A����t���s�mC�YtH���y>�������v#��O���V��;�熚���wT2��zK��{9q�Ӽ����+��@���U�6���D���:A�+���0a����LrU]��q��E�(��_(	�L�yJ���;^k'1f���î��/8&H�{T�k9X-������]2��K���U`W
��ԛ�xdb��T�+�$��Kn	���;;tWA|���r�mə�5�r�P#sY{���������0fwo�f"��������� /��kb�J�v�a]>����8�[M���M-���uGa��'���v����x -u�gP
{��tX}�q\`�O%�W>"Z
�efK2�_z�nb"Y�&�]Ǧ��X6{:��[���U�a{��Wٴr1��7҆�����|ޏ0����=giA����ggv�B�n��h��(��`��R#uo���}��<��`6����j�\o@���ZS1���4\Ɯ��������}� aV����8�SCj�B�E�F�z��S�c��)����r��b�W�K����ޚ��M�*��(d�]��a~t�����@k��,���o��S\F㸵x3�3_%�~0��6d�}�.���f��vM1K��6歱�o���� 3�55�4z$��aqT����0<�3��������\�;��r^ͰI�xN҂T�J��U�m�l�nԗ�zb��[#~q������|=?�/͜��3D��(|> UT "�E����K�2>��x�����R��ϵp�G��e�����}ӿ�j�B2�@�m���쥈#:�;Fm��7��y���4��@�E@�=�5j����}k(3�(��l��U;���{�p(���MR�Ѽ���6tR�_V��Yh��Ҡe�(��ff}@.|SZ(f�ĸ��d�N�c�%>nT�m�6��z���;]].�#�c�7�>ţ},�5���o�}�j��mT�O�ϴ�i�I�j��MS�����ۓ�|�syw��;��&��ء~f�N�Ĕvt�UBW�uW��u6��8���v{t���k��2V����=��$�9��'m���s!�?@�ff�_���F�w�5�l��Y�1(�pd�]�����c��u��N]�@;q��'.sc�T�~gk��,��U�C�;®�v�.��|���P:�b�{'U�{6UE{{�r��rkz|@�����)�m������f���d��e˳�(��ܼ�t�=�E�ݛY��(U��g�{UqqT���]çR�o�"�"AiQ(&t�cѱv�8�EԵD��榧5}�nձ�e��;�	��YL+����F�f*Ֆj��v,}w���/�hxՐ��(��?$Rv��U�{[ԥ���^��}��}�6�	���h��)��,��u�La���w���mv.�3!���{�>�er��FOl�E�a�ۛ��0rW.c%I�&�u�W��!�氌�z�c$}�bE��$�W���N��w��N���cqU�"�{��:k�,c~y׳�C�
�٪�6"�VuV˜��ӏ���L7�H(�yt�kR����s<�K�-���[��ͩ1ݜ��C�>���J��d2��z
��P�%����˻֏zUO��ΐqeB��J��kMh�d!�X��jPc�!�OH�1Y���V3F牘5&�d�[�LFo@-:�5�#Ĥ��Юc^�94�=�QǠVc<Iۙ��K�+l�5"oKXk
fRD"_��z���ض����5m0����EY�S�k7,�Ky�ԌJV�*^�5���'2��={\(��T������I���"�__I��vT]�deʷ.s�BI�{�v�t�;A�_]�ꕻ�� ㊓}�R(Rg�U
o:���[ŷ61�9�N��Z�Ӯ��Ʀj�u��N��9EW-IK��Œ��`�N�>��}� ���:���z��wO��̯O��z����6�x��V�+a4��T�w�����,h	v?f�i�#��v+�)�>M�I]O]T�!VC?i
P��sg\���h���o[��]�p�k3����������5��;i�Bv���;x�Vx�M�6E�����ն7�j�$�����%����7(�?6�{[�]�!�mKS��7�r�ATd� ⫬� ǚU�:��K��3徝�/�4��"���bPI"��H��}s��c}0�7�K�m�c�1���yL�So	�u�;��(�&�����r6�z�_�a]�x?�,ct�[֙ޙg��;�ܓ�Bt������g���8yFt�]�w��]������m�ϣ|u��H��t/��1_p��R������R�Ҝ��n��;ۤ\o`~|���h�������{ԋ�u�h��vbț�V\U���k���~��QW�o�7|���v�A@:�Ω��c��r�����ˎ��N�<u^{;e�ofgw,��d�x�z[*�%Un�WNlw�<�2�G�����(�;�+_\�w_��"�-��f����W�Z� g���_�n8�m�'�\v�컢�K-gC:�JR��ˮ��q���p�YVڨ
)����N�y��j=8̬f�ZM.��\�����Vz���l�|�����a<��j�Q����X<8w��_7C�Ol��]��Ļ��7r��9��<:b1��i��l��/��[kژ?��Gi�{�vgMԴ;5K��(���;ьζ2Y8��|��Q1�Z�)������j�ێ���^xkw]��Q��h���A=�(��z8����o%�_B�<�;+:o��%{uG��Z84�{F��v�L+�WUN!Zrc��R�K�t�o7�7H��R��+nN
�R����g륬����̏fC�p��i��_X�˱��sTM6�9��*#�����'�wx��� �A�F%�qB�ٕ����g�=���N����6q�:<��oE�ΫA�òI�<�Һ���a��^�#;�������0� ���y�͹�r��%P�7�nv��9 +g=k��:Z2X�..1�*<�xV�'�Jm�|JD��KFc��o\����1�^j
mٯZ"+3_��7ǘA�E�hJ�%�ؘ�(����½����uc.=VO��A�UN<����Y�0ә�l�{���� ݚ�Q���L��.r'-tANHaǊ��]�6�Ό01������h4xǙ�����Su�xei���׭��Z�����>��@�c����N�;}���*�TL�^�RT���.�F�c����PB���(6��E�4��M��*IqV��4�G�{������8�ԥ��u
Ӭn���ѐ�U�2��->nU��M�v�0��nfk>ŭ�Q�e풬�d\\Y������!��/mz�kk��{������U��g��� ˹�*@�Z�Q���rj9�V2��୉f�Sɯ9��r��e��V�'[o�Փ��y!�Lx�D����]�j[]��\�t�ϯ1�{�ܫ� �,\S��67��M<�E������ϭ�tT�r� ���6�VP|	8�W�7qVk�	�.�3=��ێ݉��*(4�E�(��KJ�M<�Pd�Kh���6�	�+#�(+w$7s����]K��u��$�IX��쏧���H����;c����H�о��%�h��ԓThi�w�⎞&�iҳq�Ly�ɉn����M�/,'����+���g.�M�S�B����.mr��U'r�c�oy�
��%
��=jMu(�лi^vp�B�^SG9�W��SR&��j�Xz�T�Y���KHU�jL���8�� ݂�#u�t�q�6�uѦ��9M���z�� ���sK������\Ո�	#�EG5'P�����LU֦y��Z��8+�����]
F��7E���p�-n�v{H���:'ق�Y���b;S6]��$����c)�$S�Dt���h�ߠ[�b����zs|��J�������	�� �A����xou�u�E-K����B�	��]������m;����Q,���k�'��K�Lw�σ�}g��ei�?��AK��ru��&��l���*gv�_���xJ���H'V��3hY�+�p\�eո iA��6�m^;�Ԇ,�VbO�e�+�|wΦ��;��R��a���>���+�5� ���F[aR��&�M�
S]�V�L�1��շ�XmD��.������6���{"�r�\��9l�kUv���]�fT��|fs�ѓ/-%�5Iw���*t`�P����,
D���#�il���<*�^�K�7�����f��sS~���U��uyd5Wڴ7ݔD<F:wxwR��k 4��Ɍ�0l4&�y�+&�Iutw<��7*!��TjR�m�F�p����B��t̕����I�N��h�G�Y�6��L�2������p5ܐ1�}י���958	�7�`0�x��'s_h �����t�j�[Y���+&/����G�ThR����w�S!)�X!�M�p��Q+�SPv��_y��|���rv��e�#�V��2�H��ȫC��y�v�?�0W���%3�=䭽o���d�׊d����]R������U]�XU%Ncg�����Q§-�CsBW�)=
��������3��M܎��һӘ��3�)��4�.�*�>o��<��U�R��C��n�N���V�[�E��%t��1d�I���7b��A�^��ћi/w� �>��E���KH�$i)B
�TD�,�,���E�G.A@M@O}zzzzzg_�3��:���Ϟ�9r��Q;�̧4m"�)R*�WP��ʞI�'��ק����\|Y�^�z+�-�\�=Nԋ"�b"��l�m�kF�B[j2�'?^�����}}_Y�^�����|B�;�I�"�D<�j<�D�*�z����:i�����������O�����j,*#R�J�A�J�_���i�+f�N�:t��{='��1�='�DE԰��`��ަ�R�A��4a\궫YϯOOOOO�>���=>����.qં"�#m������khV�ڣ�gԺ�KlA>943fC��Dg�('�J�X�|k�E�kb(��0�""*)͝b��E�Vڨ ��Xq�aH�$�F*�Z#��,�k����ŕ���;t�����֝��v�r;��\��*�K��|�Ţ���u�=w^�ڷ�G�k�#nJg<9^�{��c�Y�M�S�*�ݡ�%���՝`M
�κ��n�J�v�'t*��t�:� �<x�
=YN8*��Bņ7r��ק93عn�/	�|�6�\�v�݁Mh�u׷'u�[��y��5+�x旹݇�:λ�"]�v֫nݬۮ��sv�oc��ky��wv��z�5+Jl\9W\v7%��{%���>�q�	������8C9��n�OIR2A )�O'�V�bڕ�k���_?�}���P�����VZV���t�����Y[33;0��)�t�z�-�ɭ��K�bk)�;#��6KD��;N�Rb�;�{Z<{	��n�+��w�������g��ܽ�t��/>�;�Y�wU�s����^�aV=	9�|�q,32ØՕ�������"������էy�¼�U�yf�z�ӊ�^�dí���RNii��{"��ι�dѺVw�e�V�b��a��Lo.�fz�Cfr�ka�ڠ'.Lmʻ�!�z�QKr��&|{ׂݵc�[��Y����,�J���n��E^�a6��`>�x/���y8���?��_9P�B]��d�"�96���8��P�0yu>�kM����,��U�r^�-yE�i`C53�f��Zޟ@�g���4��i�RF(���p�9W7�j��kdD�g��/ƺ�F��k�%��tU:-h����/�h�ۃ���3NWu�ㇸ-���C.󲤻����fVӶ��YA��A�^�6�'�}?v�\F�ww@}��;��#��H�Tm$s�(�k�Ų:-[��
a;�q�����8��9���{X�a���'T��������7�U
f ug���;&��W��`~&�5���N�E�k>���9�,[���/l��9�@H���۾�fŞӓy�簾����WuAt�fK����	��:U��3�A��iؠ����f��sF��yW����Ҿ�Wpcٔ!��eTv�B��������2�%�o��+gN,�= ק��@t���Gc�0�ꕏĸ�L�s�jz��wx�aZ�\k�#'��ww�o����u��B`��nc����9B$�i-e0S/���i~��'�;Vz�_H�>����Q�$XA,l���3H�\0}��7�ªgp�'�d�K׏�gJ�Y�34Yқ�����q�'F�{i�';�q��a8�٤����jxa�,�5>))oX*����o�ɣ�9��Gq��KZKF��=�ͬ���k%،֬7�<m�{N+�>�K
XI�O�6t�쇺x�
�7B2�h� � "4A{s�7_wE�++[��1�[!�7.$��M�+�Ө{h�sNt�{M�g
s�f�&�N�qH�*��*�oZY�}� �F^�����"�y陙��s���ac�3��=4ojg�.��{����إ�Wt�g�v��2�U���z۪��m�x�����#WLZ�*�i��3&�1�6�9]cn�^�U��$�˧L�͡��:<�s��������x��R_x��mu��,B��T%v}g��ܠI�}K �m|9���7
{寄ߩ���<.��S�q�M�7�\�Y=aS�2�;�aF��Sйw���j����3�ywt�iuTݬ~��Z(ʺ9q���U��oHݽN��U���}]~���r^�T���z�*��Uq�x�NDآ`�I� � I�Ͻ�W����Ȑ��*�����z}������w��x�f��u��e�(��YR*Dw7�΅�Jv�fc:���yo�{���և�q��EZk�=�ۚ\�V7��坣�ͤ[[����Ԛe�Χ43;����B:>L�ľ�ѽݐ�TZ��}f 0�������L�8�ǝ;��
�8����'��,RQ���X�D � D�w���S���\!3���`���r�U����g��'f2]7jy��~|:�[e����o�����ȏ�W��f�e=[뺸S5���BXR���HS����Em�W���;�K��Ucg��<��46:Z������D���WV�o�2:qoe��R����T^�18�}Qo8�~g�N�wd+���ʀ�q�o���/j=eD���f�KAi�WuP��g_��C��`ڛ��u���9a�j[N`y]�_u�	���:��H� d�v��^ �L"ݯ�:_��$����z�♁ڌ�����Q�~Ш6��Ct�3�|���=n^)E�[KeTKyn'�,�۩��C��>�E��]�;x��-W|9b����%�0��RY,�����ɼ�J���T���i�"'�;�V4�:k��s^	�o����&	EG�����#�MAޗ��˜pj�uN�/,�3Z��2F�87�\�zJ"���Z���8i׎���'S6�#)�y�#�31���6�9˜�c��J�e�� ��7�����n�`�-ѩ���T Ig����ʊ��8n�?u��o��|���)��Q�jv�MMr����b4M�un�sJu}߿�Q�V���W�Iwa��].�3B�0��gj�Vc�'`��1ڞ���{t'wf>��7=�G\ld��@ս���f�[o�N<Vc���8���V���y��J���Ȟd�ΛkLb^�nw������U���]G(E�+�l�����˝�X)�$�ַ�\�wv�U��[.������C'0M�FmV>qm�9�u��x��c�
�b�9M`]8խ����I4.����*6=G}2)���}�0�t��\� M�Zڈ�e�e�S���ᥲ��Ta��o&�;=�/]C�p}=CcC�M*�W[�J�V-!4�A��C��>�^���R#�C)=�3W���D�9���v+�P��;<}�G"�3�;���"����	�oT,��`'�3u�y\��]��- 8�YĆ�������G�n�c3F<�=jG�U���)e���"e]X&�s&�_V�6F�wGX�Ef�wkʇ)0n�t��2��9^�D-��<�zͼ���P*��<���f�>m��+D�[�G�v��˦��8����qa3ۍ]L��]SM�]�Rd^�'�W!��!�1�r�̾8k׺M}N�g�ϒ��4"����W�TԊ#�W�]o�&]�����"gG���_74�f �ͨ؉�����{S8�4����&��iǖ��>������ת�K7�,1�N���0��7g�@ff�CQcy�������+V�7w%���jӵ'�G��o�~�0�t�����<_�u��
�E#H� ��~� N)�	��u�U�i�{�m\9Q�kv�c���'-�tL�y�x�ovvV�I������ӳs�n0�{ YQ�kCtd�s6Л��Ur��}+'�z�������fA����l���t��P�;�UIY�bC�X��h�=#�kWt�;��`���N5�c�)�W57F�����4B��F�o[gs�mKY.�1?�M�Ont�J��|��f*��,�Y��)���H3:�f��Z��W0f��ʋ�;:)�n6������^��:�{C�׈m
*~�^�y�y�]9���)~��g�G>7mUr�GL���ܫg�M.,�3l���4������5�k©�q����Uǀ��[���<:�!~���@e�Hv5d� �6�S:}q˔K)�D�Ku��ZM���&�=-*c��n���?K_���"L�ǟg c�6M�8g�����ݮ
�ۘ[5vlw��}	ʀk{��2���̵�4�a��t*3�8g��'�Ֆ�3�9j�x��;KARD�B�w�xTՋ:Vw���|��x�����,�6-�蛞N�3����;_�'�Lk�k�YUk���&�_�q�(�W���qu���~��n�}��B��%Z���Ṯ�e��_"@��{Ums��x����c�k_Qmm6�Gǻ쬂p�E=ٿw��A�i`�8Ī?�uNΡ�{.�~�$}F���x��F����x�+ǈZ|j��r��E���_��t��Y~S=+U����X(�I�1� y�-L�#glEM\��nesD�k8}F�u���z=�,b��`98j��V3`�M�Q�E� �  �������☞��{7�<��.���������C����'+':�k��M�zԪ��3�e��rz���s}la(��JZ˳�L�	�	���Wg��"+��Hu��]v���}{eOE�P:�lfj�a��(u�3�~��ATק����C����L�s]C�ctKv����ټ�-��P��rffG,<�d����W<Y�wU2يb|>iݥ��h��}@%��c�����~}��ڟf�Ǜ���'>b�W}d&KFKD1�/t�֘O�Ë{}'R���9�Ԓƌѹ�\��D�@:ݙ2�"&���l�����jDF����׹ɺ���[�'��vT@�b��7��)���F�b������vN�]�����嬍Vj��2Lu���Nsp"ݑlF�v�d��D��9:���>�3ږ�α8��Q���C}G\6f����b��aqձތ8�k#����mh��T��ca���n�-8B4a�M�;Ovwu]��ɜv�ѡ�z����ڹ6�Θ��F�H,*�����ǘ�-�c�J�S��늂��W��{�� &��,"Ae�As"L�#jF��1�v�M�`�R�%�{Qqz�ܧ^�vp�Z����L�s)�pd�vbh�*�T�R&Q�IM�:�O���̲�.�n�����G�jӕՃcm� �4x�����e��C^�2$�G���u��D�M�3k����U+��������`����}ѣy�!��6kw���XG%vuGL{)�[0fi<�a�"��U��e�B��n������.��J�E_�������=Lg׉b�!P~�fe�$j��U��Մ`5T���s{��,��tj=��7��kI�kM�w[�h�n2����/�x
�A댹�����	��^*�7S+�Į*; ����̚
��=q�E��{�֢2(7���7'�m\���Q�i���ٿ������K�5���1�jwMm�S^�c�c����P��h�07�K�k0m�5%�\CTw�����y���e�������Ico隒k��B�0�%X�TE���=���Q��`�(,�]-=��vgF��D	9ׯW@����(t2�n
D�惑�{{r[U:������!Z��:�j�\����ؠ?}U�U�ǜ��;���״66�z K�4{�̛������B�W����]�|�+Y��@W��Ɋ��:��3��X/z�
�*:�볡e��[�TI[��M+m�@�g��\�Fq�s�׬�ݑ��};P�tӏ�N4�{�=�9�����Ȍ�:ȑW���,����Bͻf-����T���@�;��w��4��摡�V�+�Cf�ܻ:c���D��}z��V1X���`k��k9���8^��Try���� ��&A4H ����_b����H6��&C�<U�Q��޵�V,�����fX$���n>�g'�����a�y�HYWF�T�7n��N�7;o����E���G�^��}Q���"�nW��hr�#�JcӈmA�Ú3]��� �UL�<�f}Ǣ���@C����e�"g:EY�fp�̃���y��s��l"����(C�3�*�9&*oP�YiYi��=��4T�>2f�}����4�>�7L��Y%�=���h��j���T�X�wsR�*V�c�^4Fۭ1ُì�h]Ǎ�NJ+]'�\�
�a`�Fd:��SZ#+(���M�F�ʸ}�;�[�`�D�nZ�9f�o�{��`���1�ֳ�h��]�7��J���t�T�c�kWsE�ѹ��cyl�,�v!io�9w+j�J�Cv����6�w8QYG�ھ�EC{�����f�ʻ�b${�0 -�]�uo��j��پ+]�T4��$���vN�~{u4�k@�|��<�<&��HX�7����i���U*�]nM��ܙ�)�fzI9e�ž�&�a`�������N���`;6�j4|��x���V	�F�kmp4^'x�UP�M	9u��f�9���Ke��4=��z��:�D�-��3�X=�a|�0�����H�R�g�*^�;P�lQ_@�Z�]�|.=����Nrl�ș��
tN�d���nּ��;G������E�t��~��5"��Ʃd�)�6N�إ�A���Y���P�������60��ćJ�|n�4��0f���@q��5*"�KQ"�^��ܽqF;m�MV���?�{������h���QO��8Z����F�[��'2�6Ң�2[-����G�7K:�_��6}A�wQY��k�>�rs�Z7;���z݉�gW	 �uݯ���5Z���1�b��?y�lp����N�v�pez��t�5ҡ[[M	6��t$(�b�2]ȷu�V\1��. �,�=Q+��#��h�AKd}�Vh���tҎi�]�2I
Ѵ�1ź
!z�2��\�O��	�����i,�>ө�Nv��f6ت�x,2�3&��w*xf�/o���\���q�����K���j��Z��|�,�[��U�3\�'��[����l��h���y����⎢�85f���'�eho��*����@�z����6�a}h6\Ekԙ����PtTUM�g#{j�.=���g������j�jȻ���<'u��En��9���f�竁�Z嗌�b�J�Q��V37�5ÊX��y�)�6g�AW���Y\y$tT��ٔ��
��D�d�[��m�g\H��uӫ��&J��@~��S�ok͵�2q�X��َ�Mĥ�˦�s�Ԁn�ӛI�U����dX�-�;:��Wpr��K�2��n��h� \��}�8�O*�҈�֏�Q8h���kE�Y��3$�q�����������|z}��m��ے�,?Ac�˔m���*x�ݧ��U%�M,���t�ӧOg�챟�����}��*L��!אQ~�����+O,�5ں2�=�'N�:t�?���~'����U#�F���>�>5R#�i�3�����:{=�:t���{?���OgOg���_m��v��&�NIEX���l^���Y?yN#:y>��====?__3��ӯ��|��@�/2��U��h�O��N`i����������������:>�>L�����9�rjd2E\\�ğ�9�K��w!P��kmE�
,bK�1��>o�Ug�T_M���}aؤ9�1AX�'�p�+*���EX�rT��ԊO-P���*��AE-��X�R
m�DEv�{���|wy	:�g1��r��p���?ud�E��P����.d]��ės�J�{�l+����
"C�F��TW���WR�]��y��d�� :�@�]vSU�R�DF�1�/�ۏeRj��F{ ���P��Nd��sRcõ��Va�4��9���G�u�G0�7�j=��W�v���>��j�kc�Jb����\_NU���ֱ���wZ�>�:k�xt���E���$�u���\���KL�f��
��_|�
��-|��c��⳧ �@Cd�ڜg#6q��ش��I�@���lנ..��Ǡ�\��.o,W>��/[�۬/O9� ��O�5̍퍏l;�]�F:�#T��=O[Js����0��v�n?x�V,	W�J�~W�����T_�$3��jJ�XY3�o�-��f�T�R�l�	:
ƈ��}���*!(�IP�h4p������� Z|��ªu_���w�3� ��.��u��U�O��g���bH���@��d�]p㗛A�eY����	R�;W Z�{2��'�=,����/��-�2��9�J���`n����ڱ��㴺�);��w�{�%I�Y�!g��m2��ˏ�g�&#غ�[��qZ�Rǲ�D���9,X4hW�X{��ig�������4j��a��l�<4�F�3�73F����'�z�:�!�|��Ly��1���W}-�H<~���8��#��)\�c"2x�������IH�`;����q�Ǯ�Wd0;�k�K��d����x�?����]�U����Mհ�
���cu��ڸԭ�wf�[3�%�W^3��=இi����N:"c����j^�&���3&cu��i��2������f^���Y���A�CdʙU�tr:�+�f������q	<�wc��nԾ$&���p v��]�oz)e%'�׍���V�W6���Շؚ�È{c���Uy��%�(E1�������p]���vNO�W��H*�C������`.����;HT�&�ت�h��˭%^���ηWCE�>�GTR��I�IpS�E�;6B'sf�0��JӶ+^����|�R84���u+pw)��q�pǑvk��g��u���m�\g�m����c�g�q(ZK�����J�/����q��:L7��?+Sw�~�·���Aѽ��^�j���ٷ.�7��j3(532��iʚ$[�O���y���:]@���	���$�6���t�Zku���1G���k�3]�Y7ݷ�R��ϱ��4
�܅�Q��h�ld�3	�W�;=�P�c������>��'���a׽��{ۆM�v��s:i�<�;5���6ӍBS
���k�\�Ss~F���w�}��Wnc+�X<��Zju�e�w���J�k�埊���d�$"HG���vl��%��h��p����`��^#���m?M��g�{���y��/y�O2S�\U5r�\���GX��O�N0��s�L�!���'�lY���["8ﮅ׮��=�g�TbMS���R��窶�;==�Q~`Q$P$�<�I%����Ϗz�S����^�\W0�M$/B��\��#�_cr(�z�q�DUPcP��'�X�I�}n�gt� }k������ݛ}+dԇ��53r6f�o(�u�\���y���#Km�����H�]D�4f�5N��<���!L�h��/�$R����̂o�x�}��{�s�YxxF��ql��j��2L�����)�1���hn�����S����f�l�,ӭ:��z��+����[k�
E3x�Eט8�:a�l���U�����v�}}W٧knp0�x���c��8�LY\..M��OG
�� ���f{����,�Z�,�����b���П1YZ���n[4�+�{	���2J�Zۡ;r�:*Y,�'96��yo=���`���ٮ��ܣ�sB�s5���z�זR6�޾Pγ�=ݓ�+߫;�ۚxk=�FA��Y�IߌHGp	Yd��������̌�@���^nG�B@=Ss��f[T+޸�}GzFA�{����6����6G��2Fb�u�'�;2�_n�f���R_��ƛ�T����pp8�"����&N�����7'#z�磷�\r�g���h���?�MǴQ/~�o��}Sz)�wn�̗Y#2��,-���C�:�'f!3g�`S��G�\�Y��|" U�%Gó�W�P�=�)���x�#��N�n����ϫ@�'����:C��=��x�w��t��a���(�$F���XU�,N�[�Ez̮��M�K�!F��,YA�=9���ќU^9C�~���-e\MT�e{�F.9Wά;D�X�&���Pw�g��:���?Rvfg��s谭��2������iȷM�޶�b9�X��:�1����d1�K�j�2}v/��b0vu��D*�Kp�~�����<Ւ���-2���"�C�S^=���%�R��y�e�tN��	w����<�2k�X͠7��%M���^��4z����fsxr�z���QJ��f�b��S>Ӫ�9�e�Y����Y8 �ݙ���O�/�y^�O��;rQD�DUg�xm�f�O�^�J�7=��=��Ou{Q�$�ݪ����xqnK�l6M���|�<�_����kSs�;��[��Z�u-�Vn��8S�l�1� �p5q���m����2�	'�ۋ�����D���kf�6��i��>{uG��|[G;�xN��Jƺ�8Й��c'�V�kڗ��	^}Ǯ��V�w�>kr���/FN�1�|��[��/�;s}���$��ѭ��Ԡ��F�  D ���U���4���9�9�`� ����[�������q�u�,���(���Z��ؗaݭ��3A%>��2}���?t׀���Rݝ���5a�J�s��g��F��S�`��֘���nh��l�l���cw�áBݯ�?^��^f7\r�'�}&@�:�
n����cf�Si�eš��9M��C]�Q";:F���y��L}^��9��1��M��o[�3�A��!��fӭ��h�z�[����o�&��Z3���Ro��sw�^��
ƥ�����;����P�ɔ3kw�Wlϊ:-�z%�A)�Cg���}��TƘ�pV��{��7�vk~��6�m�]�pq�Ԟ��K
�aQ�g�XR]�k;���3+-�tŮ�b�`N&�a������8թWv����\e��9���A�l�|��5�^����x��<����oh�4e�yD<ݵn<�,[d[0T�nǗ�g.l�d���y	;6��T�y�-�����L�j��/�i`��ɪ�N3����tBv�.�8.�O���!���h4ɶ�SJP�"fT��Y������vCM�L���bCneɛ��q�z�p�?��r����Ċ%I��sG��HϽr�����}�삎t��U�[tԴ�f=��)5d�G�#%��C�/����ϏW��)����el��T������u��c���s-���'�ķ7F����3�56u�12�n{�-�!�`
���e��6^�ʓsW/2�w�g��jPm�W=�+��}-���wr���y�E�m��Y���v/sE�s���$0k�V��V���Hg�E��N�t�{���sS��\��W��̃�p���[]�9�e���w��m�O@��n������R�r��8��7f=}�͎1��8��<�֎��m�$"�����99�u�a��\w-�?�Y�K�̹��zћ��n{]��!;	�H�����e�l_�3!��6��]>k�qmʖ�2_�2�b���:��f��6���]��s3*N����S�ԦfrG[��TgQH@�PW5����wuWN!�dr��Y�A��)��Yo��t���y�C���+���X;Q�P[���L�
5�'�8�oy�ǜ�Y�0��|�=t�]���{��Gr�/G^�=������\Gkk������s�m����?�R�S{IX6Cy]t�v��c���[zEC?&��3�}y����ۮ��/4F�w�r��f���A��UU�ګ�w\��>�4�tgn�aO��\�u�u.�U�����d4D�װIn����nE���w�kM��n� =û m.��l�W�.�7��x����Z�R!��k�}�٢d��逊3 	����+��Q��~x���@Ʊξv��7ۤ�n
��n-��#;�^�~�=�=g�6S0nԵ{3������,rt�$��m�ԣ��H�(�P}�43�/��Zx�r��G;�m��Z��p�T`�l�h(@��2=��l+�m��ꤩ|P���~~���� �<�W3��eHwl�z���vV˳u�p�pR��Q�3�ԯ7�����r-�k�q(R
�C�d5HW����է�m�s)wg,N��]��)X�l�n���6���qkA>钍�g�}o$�Bxy�S�v��o1�RO��1�;"��#��݂5��`Β	g�|e��0M����Z���"]�i��|�����ʉ������i�'�*���u�M{z��y��j��EWp=ј�~���33o�L�/#���0��*^��Nq���y�;y�k�2��-=�Z0���g-��.N_|�����
 $�'覾���x��[Ş�&.���vx������L��*m��8s:��1猀���="7՗B���ϹN��|�c�^�[��M�a9�s_�o0֤>{#̺�=͸�u,1w[.��$�ټ��@҃�*�j���v�-���?7��`Ju:�0�5w9\E5�β�}��W�C���Z��.Ǌq�~��c^��m�x�`vz�;�&���{��� �"j��-����Ut�S����TӋ���^�ô�<�ؿtk}�&��ǿ��!G��Q�N�o[��_U�9���ɝE묓tP��3�K��$�P�ۇ��o��/�M=�y���э��1+���H�=a�Gk[�N�Ǩ�����������%�J�H��;y�����}���is��q���3!�&={'˵g�����ʡ���)R�g�ͺ&(�8���*2�9z�3�� ƿ�O�(�u�+Em��t�=�?q�|���D�2�jCOc�}�Dw�d����)}㙹u�xW#�.-E�g�yN��FzFW�Lj̏�ދSU콦j�	`��\xI���1�Ҋܳ�R������=&���8Փ�����ҘG_ӄ��2Tx�|[�V.���>m�U�Ϩ .�x,ݗ�]ш�g���m����Z�&�ؙ�ژem�wfY���4�\ײ�#[��l���r�5�٩޴:љ������H�(Q�팫��ۑ��6!�G�2�pn�ʰBˋ~���5����ļ�3zE�U1 0�ڎj-FV�V�n�S�������`�	�b�� ���ĺ�Ϗ���?��W�_�?��K����
 ����AEO�>?�ǈ��PQN��|!��>Ns� ��� �J�H��@�"�������� !*����XBEa	@!	 ! a H�E�2�D���*���B"!(@�(�*�>`�*�@�(	/P��$H� `B�@$ �z�q!D�E B�	%DH�T BPP�PB$T P� B@@�Q A�P B@�$T� �P BU@�	X��X��Q�!"0!*0!�!(�u�>
0! �!�!0!*0!(�!*0!*0!"�!<�p�	Q��	Q�	Q�Q�`�BA`BT~|����X����H�HB� �A0! @ @��!H�@�,@ �q�l���_�� &B�AH���^���������������?����?���?���~��?��_�?������DAW���������D_��QX�������2�������A�?���_��?w�?���������C���	�@s���P~��s�<EUPeU�UP� h 
P�Uh@DJ)�i)DJDH X�ZZ�`�bX�`�i Y�Y�Y�X V��E�%V Z��%F Y  ��BQa�h�eA` ZU�XF�
� X�d!X�Y�hF@
E��bE��YX$Y�d � (D�hV�`	V`X�dYV%�`�e	 ��A�fE�V`XE�V%XQ�`�b�V	A�d�`%Y�	 �`�`�bE��e �V`YXIP�d�` X�b !XV`X$FT Y�a�` X�%X`YdY	F ��`Y X �Q�$YVBU�Ve�eB� �V%` %�d�`eD�
Q�V�h`YU�E�XaZ�% �i�iV$%XR���V�b� ZE�Y�i �hVAbUDI�IE��D�"Q�D�
Di$�� ��_����F�E
Qh@) V�T�����������O�AE((@hTT�P����?�������@��}���AD~��/���g�����������<c�_����Dt?�؟����O�* ���_�C�0���(����C�EDp?����}!��~�C�`����3����8	o�������Q_�R����C�?�������� ~�O�0��<ADs����p
 ����C���+��'������q�۠�����w`(��i�ԟ~��8���?�>�����7���D_�=0p?�Ay��˿����Pq������)�ѡ��KF��0(���1|�J��*��%	UBT������HF�)�i��`�P�D�Q�)*(J���b���PEI*�*�n�R*�UEQ֣,�U����*��3V�Z͊fY��V���h�k@�5U��b�-���M��Zv�d�-
�j��l���Z�-�ɚ�f��Q`ӳ���d���Tƌ���ZVړ1�"ZȤ���cK[I�eeb5[kYk3k(�4ԣKiMR��m��b�SjZ̓f�ճf�-e���M��fiU�M��;� �
y��� [�u��[Zjq���Z髶\�
�%(5����R����MMn]f�mvݵ��gUE!�U���)���Uvݭ�Sa����յ
���M3$յ��Z�x  .�CB�
v���Z���"�
(P����B�MD�ySU�����v2�Wke��ֶ��Ml]��SKV���R�B�F�ie-YT�;�٩kmj��Ҷ�k*f�66�II05�x  6�U[c�P͎n]S4j�Isp���a%)T� �j����*�(���֔���R��宋U�#����7m�e	[-�Y���ՙ�  YꁣԹ�Ԯ�%In�\�N���v�ꮖ훚J�C�ݮ��@uv+l�YŎ�ۧS]v�T��c��Uթs����V�ٲV��Z�Yem�^  �z�H굩t�h�SR3f�V���S�h�.pj)Щ�'B����)JU]���UZԷ\��v�U[�F�q�[%aY���m�X��  n�jʔ�N�M
��TiT���p  9˜  �` �g+� ��� P5a@ �� : .q2l�l����R�̭Ҵ���  w^ hoN  u� ��U� [��  7u8R��ۀ�
v�N  e0  ;W7  ۛClHٴ�RҪ�,�X�  f�  ��P(B�0  �  (nvp  I���M� @l�� *�-.� ��Z�4  �j�6��i��Xɭ� e�  =�[@� C� 7[�  3�U�  �L  ��  ��`�7  4g\� ��*��l��*���3M�Z�U�  ��  vv�  �m�  �*`� ݷ  � @3�n� �9��&�� 
9���+�<�iJT � Oh�JJ�3P ��U?�=BRf�4��@O��I4��S�b�U*��  IP&UQ� ���oۋ�Q���+9�#Z�e*��4�D=�è&�`�0Xn�����=���f���o{�7�;�h
���@?�Q�r�+�XAO���?��U�tɜ\#�U���ͪ�w�&�2*��:4r��ڒTi��`��t7��w+T��Y0����6���ʒ� 5�z���YT@���n�Mbb�ҦʬX)GPY�]bf�f��Q+�7�l�a$ic*��׀��e
@'��Y���.fS�E��.i�ɟګj�K�]YȲL�� v4�w����gY7��o4@2
F8+q��$m)ZظNۦ���H%a�J�Ki���S�4���Q�3�w�9kFr�ED���6d��x�t
X���ڷ�C,P8�t^�r#F+qR��6���.��eN��x��f��n�q9�����g�1�����
��f��Hb�$���2=�00�M�b���1m���hѵ�f[FY��V�d�h�7b���52�j+]�A�1P׭�����`��p֢m���X�T��/"�&��׋~��ނQnAaV�	R����C�=b��V�#��tĆ�K灪�Y��KC ��ov��2�:� �(�U����ER��d1�x��{`;ڹ��Bǡ���T0n��������T��EAb�Q�[�TvͼŧuR��fU�X�SlU:�4����`��q�&S�+Z�t�mo֛7l��ط�]���9M�`�W���%59����&�抗�K75&��J|]�ѥ�5v�-=�c� `e�̅:Ua�
�<��2wn���G)�@�\���]B�k.mGn��G V*��h$�9�iѥ2�����v�̧F
Z�v>{��QїtO�Ē������R�7g,��R��ѡ�5�,�DN��6�P�Ll��@ĥ��lVӛ�̯�J̻��ߥ*9OjD�~�
[��ye���f�+e���<!$%�R���ӷR�@��^�B���Ux��jHb��V��)���Ӧ�1v��E*��Y��R��p��y��pjÙW��V���p�YB�9� y��G@��2�v��ƅ+��ð�zE$�n��`����r�'/�9�#(^�
�S�#*��w3 {ne+`�w,�gS5p���toiL�h��2�ix��R��m@sq<"��6�<�p8b5uf�Q+\!e	x�W��+i1t���i�0D!��n���ǁ U�Km���5�A����u��iJ�d����7��Pꭴ�$i��n���
X�p;m������N6�:�bHiE��c�;���k��#�gdz�4��oSiC������
u�϶�-ݡE�c.�B������f �"�<� Z3kU�9 ݺ;n�*�C+%LD��/%*.:�Y�ۧ4z {yb&�fln=C��IN�{ʘ ܂��[���
�"'�MӇ2'-�A�f��Q���VV�Q���M9�VQ�Ziؓt⥔�w�ᆵb;������>B�nbGn*Q��s3�T��0ުzh@�N��,���Ŋ��A�t���sS��d5>�.����N�4��Q9bQ�1j���:J���ڵF�CF����wN1�^I�wH��T�-�Ea��t[Ĳ�سq�LU�N���ڱF-���A$ٛN��(@�ȇhK�س2b�gi��Un��I��P��L���yz��-��мXR�~gV�_^�Ñ��HXڇSF�G,տ�)[OE�����3e�lf�~%��k�Q�V +9�YJjp�n�v%Su�����X�	ٲN��F�V�E9nn�0���t��ֻ��"n=��X���G���e
��
�N��t)��+g�s���4�~|�r�i4�+��*_[vr�6
v���V��p7[���ɸ0��)3�屎���F���Sd��0Ӽan����Eg�r�)�n�X�*&�]dP'���:b�	d�W�%]P�D;�n��P�6�::�� &
Amd���k.༠�H�k@��?��Л V���&V��Sif��,	8TCbrB�5D4	��f�%�bU�����*Zt�Y�u��z(�ť��2��[� �(�bwB�[J�h:����KcCsV���.XJ�C���GZEթ��B΅hյ6; �̘n*Y�m��0%H���Qf�Q��tv�%-�H�8�b��4�d��ӔyfM2�/$*��������z�"Y�C@٭j�e^^���x`��Ňkiag�)5x��Z���"Kw,^��Ow�W��܌�hm/h�]�1n�p� �Y�\R�t"�gz<��;2r&�p��j,�b��%8��+���%.�z�9����_c؝bfa�S�I-2�Ej�0�32��/.c�;��W�N���bEp�f�G[@�5jY��p�Ǹ*DU�m�
 �BI�Ď�n^�V�nc��oE`��
��J���u��HnPO*m�m�N�Q�9WQd�����o6M�M)�S�h����E��<��Kʁ'X.5BU�y�[u2%�(�Z�����--��(����f��i�rF2�h�����$Am�Vn��\�aaY6�#�IY0n�DXGo�;h�kPv��b�t�*�hG/BL;؈:/�r3SCl�%�>�������{���o啱bj�0��ik!�5?��w2��*%tsV�% �,��۫�qV�E�N��LT��K���ӥ/ֺf��A���cB�'YZ0����I�WZ�e�O^fR����§�V�� �=��Sq��&�^��u�
r��<2�L2+y��0�eZ1Vd.�e�ʟ��d�U2&,;���ە��݀����y/Kz��)�B�T�r�\*��%���re��{�D��$d�����/c-[����^]&�-̻��H�\��uO+A���`y`]Ip�[9�-��X��ڱ��4�.�
ƣX*"x r�7� �E�$l�EݲIv��A�*)�3D@��u*�f^Qu�,�ݽ� u*ȩKL� J��jr�����&����omJ���{~���k�L��~EDp�]��2�ܴ@m@���!�����̫/!�tm��fe@�
<�1����(��7m�M0ļW��S�
Ǎ�s+ �OQ���-dM����P�b�D,�D�b�+�n�:\,�sU=�%]+�*7X���t�(�[��f6�t��1�T�G{+L��~�7����v�%d3c�F9���b�n��̵�e<;E�;���h]X&[
-��E�3q�cMY�7X�&��i���wun�&Ɣ��-ӛ�ږh|ۣk*;av4*���X葌h�*�P��vM�,E+$��7H�Q�S�.enl���ڱ4S3��(�M[����l�b��Q�p�:���e-j�,H(����7rȪb��7n㼌�A��J�l��"rY��V��MJ�C�d��g.����t������H������	E��g#�H�2b���Y5�4`l^�z-�)^IZ�+t�L;5��:l#l@��eei���ӷu�V�~.RygX5�-Zz�62�e�	��Bw*�*x��j,��.v!;�`�+S���k3b�
e֥R��/\�Q i�ӎj�� B����Eޗt��d��!I�-�ᢓ��T�֢;1k6���S�@f��p�W�f�KV���Wć���-��2if������¼���	i���͍����aָAy�b(��&����ᤨ�n��>�-�v*��MĆJ0S�g/-Ӥ)�0����J�ܸA�m��y����1a�gw[�Uv��y�jG��rou$�K1�#�p�Ɂ�EZ�H7��U��P�iʼb�3�v�P�$��PB����"�����7*k�ؕ�AK m���
�[�f���x�i�ӻ��x�?KmRօ�W��ݧq�� H��*�]�Yh��	�B╣m¢�kl����-^�Ԕ�[��m��30kM���� ,�[b\t��b�H�,�W8�����7DE �Hf�3x5����Ծk�I���V�!'�@ݴ�_�A� ���I2��	�Z˩��`�7P��lS��RhA��L�owYHj�Zc2�sP�k]%��!%��n��wESH\�o1�4�8������^�k���ɺ~�[�H+X",R�;������i&����];9Ks^�I�,@uT�B3�k5��j�׶����j�c+m:	!Enm���ށR�#B���Å�wԖ�Z�{E�ۢ�7
Id{��,�הfY����:�ۘ�4ͫj7Y�.�X�Rt2�)zYZ���[Vo	˼�!�a`�70��n���,F錼*�@ٶ#-ꚋ��nJ�#���8q�z$-W���d���H�,��a��S���=�۸�m�p���vBX��ڹ�K,�K	֞	�Z�C�N� u�2������e&�+.-ӱ�_c�xd�OlnԘ6��[{�͈JEsQ�7w��m٧UC�e�3�mn	�B�KM��I�`�6�M��S։�G�iV.�3h!u5Q<��G���VR)� m�m��ں��-3h��5IX�ΙwF�&���TA����P��.,���{!획ɨ�U�{��wXJ�y����]�b�m8�X���N��$/V[�vd�A2���f��V��:��8��
�A������;�H�L��u��ҭ4�D�S� ܕb^ӗ�N�]���F�C�L������(�b�7lQ,�j�a��^�G$ѱ�&2���vj��=�_@$��2̭�h��&%�@°V�Y�e���g �#ѰQ��+��7k&P!m��gA��X�����8ڦ�Fj}���x���E�w��a�ȴU�8S>+��ao��l���!^"4=�-T֣o�F+��rΫ����c�Vb�Ј<3j�_J��2�b�	�śgaI�¬݄�\T��K+'Z��؍���e9�l��ѕ�B�N�QX^�d֦M��"� ��Q-����kl�"��eSB���bCOk�z|���T%e�̦�#�nJƢ�ѺVV��<���ƨ:@�U-<�9ӻz�Hǉ!�c�S7B�.�O/otl�٣X�91�iǗ�է����Bhy��b���^�O,C���i	S������ �'�d��Z��::me#��
 ��1��⣓�l�!l�*h�v��/)ͩn���s^�.�Et��rV��Y �H�̽nΊo�HF���٫E�\R��p��d�|�w4��4�o�!aeM')�x����įC��X��l�7+b�{���(�x�iSu�f������,�Sk@V�2T@k���T�z� T�T�, JK�Ӗ[�!�v/#9J�����f���-=��h���c�E�0X����X�p!z��Р�&�*Vht��EA�s"��@m�w*�ң�3)m@7v��kF�Sk	F��U�]��W�V�Zm�J��y��PP[�@4.�X$����|2��S�:�IN�& H����>نe�a�Dn�!F�Ԫ܄�̢>�nm�1�ǈ�.�����K�Q�m��w��S`��Z�p%Eq42PU.��w@k(f�Vڔ���]!�J��f���J�N#*7G~�p�H�y{J�N؄��Y��Rm�`僷f���lV��v�(�^+���k,ӽZ5�7�e��*ڈ���V1�SQʐ�W>A����V�mn�C6?�V��լ�P b������S(�ZAh�"�,�T��U�4è�hS�"ɺ��.`����Q-�nܠ�ԏ��V��Eͨt���&D���X�ZWD"iɷ4�yCST�Zf��'L��Դ�5�j�6#5Q^IM^07^��zڒ淟8�e��]X�N�ӣ,m%�b�w�b�L/1�ƶ���mO����7r��q�nP�ֶ��6l$kUX�ܴ��Y*J��R��%=.9���"��7�����T[$Al�$����ڠjl��oN���B-8�֕��@2.`�Q]@�qӣg*����U�b����4Q�gi�ZF��h^������$fǆ����OH�B�r�[dX[H�,*8l�6�{N�Fƨ����-������E,�zs	*���Q+��*�jKu橍�`�5}j���T��*3{$��@Z���r�r�1kwϵ`6q䭧Q���b��1����&..8�A������b�5!m��r�V�K�0$PqXO9VP��9J�F޲-{�lL�6N)����T*d،N�NXI�\�������c4��YY�c�C�u�^��]�]%i���n�OopZ4�'
���Kp����g�ob��5�����RQ��њaPe��ڱ�@fXC����!���L'��!�n`��!y�X�f�)K��fk�͗X�#�K�f
��Y��=n�<��\,٤9/X8(&�d����xD�`��u��������+6�B]:ZE GPz��d���/��B�̉L7��fՔ�.�A�b1S�R��Y�׀MA�g/Q2#�G�N<ӹ$�2���4#����\�6�ic�4:&ګ� �v�m�PN-Ղ	%n'Jd��s6�E�ڦsS'Y��^m�Y�2-#E�?castQ���8ʶpiT�gd�Ⱥѧni�NָKe�^+xqn� ���ƭOq7p��e
OZ���lK�Ky�b ������ڀ���%op֫40hY-�w��U��X�
�c�SkV)S#kr�,R�B�(v��j�c̗�y�`.�gʎ�n͇4�)z*X%<A�����I��+v��[�)/�;@$"U�i�<'q㺰�P�j�EB�^պwDP��Sub7��՘��3���ͫ�R�!23���tb�)U�Z�5�m�?��(�-*q�W�P5�7�P�r�2wQ�Pn�{:��=�R����R��,�Iז``��q��m�gq��6�t([��/<Hkz���5_��>ԥ�F����{�,���Z�kQ��`0cUv�|����t��ml��訋��q�y|������ܯyd��2�2�4��X��]�>�K����ܕv��ً:W,E���n��%E�8�"�I|B�1"n��y{4ҙI����I�k8qo?F������M�Sv�.��^�dn������:�}1��~8�q����	�U-�ScLCsO,�6�^�k�7z��F�&3���W܆�2�v��e�Ġ)ΒA�����K�\m���������O��t�z̼L5/�#�nof���G�3�1��21L�Yo!��ŕ��uB�=F�R�n� "��RL���R���N��_9�I�&RYi7Yy+���E�Q�[dm�A^�Gd��勁�Es�{p�ͦ�-o>���ݬo+t���5��d����P��}YY�wll��nZ��qu(�L�}�<ڀ��N��Ι��|���}AN!x�[=a�d(T���T�U���;#_e�
j�.����u�G�Z
AŁY�=������㆒i�WR���>�-5�-3oS�YxW>̓ Ve@;$�'�$q���J���
���yA]*�E�h,�w�)}��N�l7q��s�>�̾���^���e�Ap�;�h�6�pE��L3��*��q*;�>�Bg+v�_f.补�Z/9$�
�b�&���|�u]���ܾ�DL��H��:�J@)d�+������Y��1t��ӑr8lTTa�9m������V^;av����F��Ϯ��<;s�qgF�$�Ԇ��=�-���em��x4���Ƭ8��ņ����X���������9婈Z��o�v�w1��H-p��ŏ��@���ۮ3g���m�m5zևAD;�
�@��f��e\�i	H�)�.�Pu��k�MmW��j���d�e V���|/����8[l��0խB�Zb�ǺzX��޿`��Ed�ޓ����o*z���e�����+�C+�ҴV�i��Ρ�E[�w&�k��J��S����km>���_��PN��n�h.h�:�Nt�p��"2��rm�w�y'0��7����)�:+�)�����/k�d���Չi��>�����siB�9Z�ed���p>H�Xv�	>��O�Jn�&�-E%��\��n]o��I���h��-\��X�
yբ'��A(�ޢ�l���]p]�0_�V�y�19rt|�5�mGJe���&���U�Is�7��|Wf"yU�7ܭ��qs�͊�T�J_Q�gx_'l��^��[��<�{��q�I-n��/Vælp���A��r"�����X ƺ�iV���r��qr;4G��4����MM�T�����z� ��lDv���#z�Ү<�Ί���ݛ��X���!R���n���v��z=��i�c<��}1{����~�孉(��2�:��c]�!�E�r�)g�}/�s���[oB5��}����{Q��\ow�z*ʊΔiH��:):����b�sQ�J�֠���]2�L�zYu�����Y��{i�^�=�|����p��wmٴ��{�/J7ªWp6�9zzl�Z��aWg�S$�o��x�66+p:�3;2�_��O"� =�[-�v�X��۬9�]����O7�=d�L�Sٳ4�:lP6,�¬.�����>�}لlr��Jc[�&'u=�Y���m�����Lq����a�y�*�n?<<��ݔ8�{}u1Z>0ei R�vE.N�\v/n��q���H�u�gLy�a\"�<�c��][|���b�BOl^L����G��>	���ɻ��CGU�p�O ��H[�j�/���گ��rF�b*JE
�?L�<�g��v��!�\{��T�]r�Kq�X+�����}���W�C��(G3�C����gw.}P %��|r��rum9VjD僼Lu;1��p<r-����"O�òy�r����展�]=8=�&x����r`�_pP��gB��8�'��au6�+[�+*e�#:�x�:)�����:غ���ۣ�J�fAf1ea�{4U��L���7-���۝�Sr��p��R���?+�-,��U�>��J�<��J�zX�\(|���#�}{%,pX�y�#`]ac�k��kE�׳D���]�b���Δ�_���ڥY���fT��yƺe�˸�e�UX����)Ko�mIF�m�[`�
��@ֽ6f� C�S]dnec�ҝ�S���Jb�tc]���V�Jַ���si�j��� ��K�c�_�"$Ǿ�C30������c	��`e?\oh+�CwⰎ�9�����d��NlV+K`�יt�̙�l� �uן�Ȍ9�+�9�d�!���x�`����^7�G�f;��1����.T�����kZ��P��*z�;Wogs�D�xWMY�ð(Y�Y�ږhk%��9����G�f���t��<^�7�O�~�ޢq�Z�u��o���j��a]���XGN�j]-���nf����yJG-,�-y�7��ا.u���G�8;\]�~����[+��<�L�ʎч��r�c��_.ǈ ��J��-lU`���';�Ҷ��K�h�*ި��FVۊG�Ҍ�Ά�YA�~ջW/w�0��F��.\G0a���Pܻ�Q{�3���(J
	1�>Nv�gLYq��u�O�����7Pʻ�9�F�Lҝ�rK�nf���N;ԁ53\e(���oSM�/�
R�GǗvQvn�IWqB��I����`ȝ�k��a7�@�9���V����	�1;�0��Ƴ�r�\toujp�\3��5��!]��J�q�R���w�hݿ`�@��PS��K/@=�����:ѡ=��r���)uT�U��c�5�����������S��n���B��^X{{�X�6I�%_=靲�kK�iu�8Ǵ��Y�i�kr��<-k`���@A���{0���Er�PY�˸H6�T����`.�ͷj���M�L��K�SWa������b"���=W�����9R�7�*�����1�����c�{<{ �4֊�"4�\�ѕ��v�tT��'��ݽ�X�w7�9���e�~z��2����c.��qb|�P�8Q��\w.1*;L�G���9�Z�Ic�GX�eY�Pd�����3)<0cc0�îѦ0��-�k��7$3v����>�q �x��!Z��ˬ�YJ��A�bM��{HwM;e���WoR��Ӯ��Pe����R�e�e��=��0ݽ��&tSL��sk�sq�M�wN\��{��W��A��3��a��7�tG����$���M*�e}3��WZk�l�Ⱥ=XU��%Yi���aj��.��a���*6�Z����f*$�7��tS��-*�t]G��-�X�c[��E5.Y�35L:�n�g��:��B�7W�8��2;��y��S� /9s�Nz�i����R��������J^�m��^Ň�,ܾR��|[����ٚ������{@�gC96�d.��+,�۹WQ��Ȝ�'k=wr��!_̹�����z�{��Sw��mf�N�B�1��5�J�,�O+6�\����1ݣsjl$�hh)��U�q���l�c:b��kcu
˥�3gR�Mu$�C}��,<�x*�qv��v�f��\�q��{E��<�]���+�y7�ʱΗ�$�;,�)�Q���j��S�;9��O�m��e��ǲF��{����n�\$ȫߣ�;ר��{��܋%bv���l�\��hU��H�s�
~�e=����-���n��'�ͱ�:ٻ�t�ֲ���}[Ӈ��=�tH��Î/�њ���́�����ض���ޚ+{v�ʊ��3Y꒭c�kJ]]Rʉ�ۘ�����Gj�y�0��K~!�M�S��S�N*�u�`��H�gݬӽo,0+x��)nD򕼠z�WdY�L��3%�\��z�����D�E�}e���{LMy�2
̼�K[���۠�Gk&�C&7�uu���b�q������U�W��r˨��Q^r}{7�㤩���O�ITp�	ohn�O�f���O��L����RC�2���Xp&��m�N�}��yč&�s���v1�*�� �k޴-zK��j�n�R�6_\�Se�;�,'Ք���w%졾���E�ZT�ߦ,w��X.1����F�;Uνun�mܺ�.�[kl�3����m�<��Q��C7N��1�ȸ�T�gl��_��U�1o��Q��4o�����dv&����+5������%I%��5�[v1ï&,+3[ٔ���T���+
�ɤ*g' d�K�_�ա����֌�uXX�օ�h-�vk��	�}�]��3;�+CZZ���a*4�z��<D��D��^���"��Z��j6�N��p]�*[���ĳ{�0�$`t��aӛ8�9�)�;m
(��;u0�]�����.�s��s��#'L�1�]n�U��g�7�r�j*��:t�tU�;�֣�����qJ+y��*E��=�ef�4���q�)pP� �Z&��PK#J\z4emFwZ��[E�N+��c�69���u��:[����:�mp2O3�\�}�_�� ����Ê>cE0�wi#R��4`�3���6��]�uaϱ�efF�i���1c�A۶�u�hBm��dy����� �:�Fd3,��ٷ���<a��o@oi^�yj$u.øe_d6�k�a-���W;0ˆx	�맴�nx�DqmG���*�]V�{%�͛i3�,/:�Y�Z���m�ӆY!ӎ�:99s��PeH�c	�6�e���e�b)�[�[4�9��oj�AnV�]�[kR/�<�RҀ���_�J�L�vC����ӘGcn+����[O��%R�=�e�Y|�'�Bny��[�g�a���Ý�]��(�]uZ���DBY;v޵��՜{u���Fև
�ɔCsR�� �Q�fمnyoQQtz��w"��o!�C�$��
,���#8̽�6����84�x�a�s(XH�u_��αXn��/E��Ɗ�d�ͷH�қ���E����G�:x:ji�2�o^}��O�F�"�M��ۦ#|�oa��C��|��5R�.{��x��&n�J
��$u�ǻy�Y[������Ŷ�L5��e9�}�g�&|�:�|�E7:t%���6�ˈ�Y� �1`�N�v`������|`C�4��>�t�E�y��;����������+�ÒX��RHy#m���^#g��K:�٤�Ƌ�kr��t4�qu:����f�9����U.��;���$r-��sn@j�5�B�+��:gN�O��a����~q����y���v<���"��'e�r%\�t���nµa���|Sô�F���5ăgiA�jج���T��L
���t�z`�'����x�E�>	� ��m Tz!�����ep��8<.o�a���t��N����\w)q�t:�&K�6�M��<Լ�`���{Q&{$�;;�� ��2��2\3v'�iq{�'��p4��wE퓝��Ȕ��f ��WR;���c(;[k���b�!*h�@XxhȒ������Z�+ ��;���oK���]6.;�@I{o�5�$aw%շ��������5K�JW��y0L��%laj��S����L���=(�n��^E-�9�ݤG��&��B���ި�ȦU�1]�^fB̍3�x�xsPnv__o�6X׍0��˔�ަ��\�r]�E�Z�����*���l.km\}5��c k\OOt]��9����чA#� G[k��gFe�(��U�+Wg�`���..p9˝`R�c7���})�А4o�GV��f���b����\O��i�K�h�앶R����(��ݮ��ݖ
F 4-rl�kݗ|�yN�����A�;5X
]�(�;!��)�eۺ7ک"�l��u��_���v�q]�ğ���;΍b��Դ�:�!I�7fe�(���ŉ;��v	"�+�@Z��ڂ��y�`�׺qU�Yu�4q�z���;W�܋�����m��4�����#/8Ѻ ^n,�N\.'���W�_���о/���"����t��`�YS��̃\U�����\�Z3N ������o�go�
7n�%��K�#:�� f��1@3��D��ή�� ��:��c���V��fmf�YM�xZ���Z�7Q��8�7Wsf���.��˧v�#�,�u8)A_8�����#<��m:³$,	�˕"��.b�v��*0�e��eC�N]�4d����#���MJn��A��\[M�r��(<�ާ�a�[3 �m��b�W���H��F��u�2�c45�oD��xt�@�������Ҩ��z!ʜ����o>�Y�K��1@c�6��+6(�(S�ͫP�5A��3ӍK[Ve�a]p������o,���6�*��bin��v��9�V���j�,���tevĉ:_A))��A�+�z!��]�Wv�{��Թ��m�r��1�D'�T{��u�I��Qf��=��y!�dK޸c�J�����__z��?K��w߯�*����,W�%w���u,�z��:�;h�{�:�2�uŚU��lv�M�����iO���uh�1<���蓷�N��Kb��GBK���r�צ����@-��x�E}#�[VJ�/�������B�oz<�i�>a��˭�d���f}�ff}������y�����n�u<
~d� �2���]G)�k�����y�ʎ������i��J�9s���c�����O\���4kZ��^�wU�2���4�]'$c�[e��W}���r��Օ�ߗX�n��mm���k�X;\;i#������9��)�j�W���M=���W2����]-W�orm���}Ѹ�d�뢇1�U�*Z���(I�lcI�@�w]����T����y:���Z��V�sW�BFAzh�#�;6e��-��h�WFD�Hl�')��^Lvw���z��3�̾���+t��� \ �\�sh�;B�ZNމx�l�9����4L���N;Q��;�_�J1��(�vJ���Zι�{��`{�]���y��*�*��q�t5P���t*��6��\[�B���Z���l}ݪ�^��ф��Ӷ��BZϽ�����n^�v�����n!9:���x-�o�Z++/FR�`Us[%ݸ�
fu>Xv�ʛ�X�h<�5��t1P�`d/�p��eXv-�fB87���*˃�� ��}(�p�*�9�7����K����\�踉���<.�`]�0�˗Q��f���瘫�⻨��(K�x��]g������Vq�z��n��������y��t�	C�0�$\��j`�ZZ&�k��q�=y�]�q1���ԋ	"�����rw���0��2����G��{d�1`�xM[Z�ywd��i� ����	^3�xT,]��D�ÖV��1H�d/���r�6c���tQ�Ƃ
��D�]=lQ�*��彬[LU��;s`A�x����)��t�/���%�@&D˛��Yf�n���=%q�Y�/jJѴ�Q{��#i�_
ã��1�A]��kP���n�ީ���o�q�c���6/��,O�i�}-��^${�����M�s��>��\�+��MY�lȍ` ꧲:��Gi#^><J��ۜnu����5m'PS��\L���X�n;"��;$�l!۫o���1�6�Q�^�65X�磫.u3�-�?:���`�����*GҮO{'˅�p��Ő=ڤ=��p�Ζ�.��&{>%��@�f�|���(<��/���U.9�s���.�-�y��ȁ�+����f�CY�:N�j�7*���Y8&*`!����y�<��f�{�}>��<b����}�Ԭ!9������3��Юﮡ�GÉ˝f����,�e��B�]Nˆ]�ܲ7��`�X�����X;�*bT��E}u��p�]���N�l�b�����X�	:�Ls,Q[��I��{hHq��c�����{j���K2֚۠�VUN��aq�r�UsXr�'�z��ΞmC��1�(�{4�r��5e��^��N��Na|�+cv� ԝu;Z�'��=PXÛ��[���+�[n䩜k���h�.co�F�Z�Q~�e۩���O%k����s;X��K��л����J�ko��ϛ�xa�sE�{��EcT��XV�*zn�o.����7ږ��L�wt�n�K' ;��P��h��m{��)h7���>�x��1+��&�;"�	ܫ.͐C|x+&��6���ǷVnRMGj�*̏l");��Ӗ�VJy�b�C�����6[B��[+;nX��e�����.a�{�n�7A��ٔCMa'������O1]!�s��]n����[��mВ�U�[n��n�kV�9X8����!d���6��J�u��9cA��o���W�$�=�}���S�3��c;���ٸ�xd9ͦ��^�.�C(�gst��.�`X�j��x�Q��\�Le-�5Y@&�s���ue ́��xԤ3&9u�v�jp4�;m�g"��@�|�,�q�VYWb�������ܨ�rp+�b�z��3�<�([��p�o7p�B,��W2e(��vcWIۅԔa��gh��dL�.�����GU�v	w�3V��v0c�c�ըi]3�i��\�y[m��ѯ����E��gv��ٴ��̈́���j�>�����̌��r�a�}�P�y)�,p��pj���	3�6Ҙ;��m]pBt�6�Vq7��g1 �1G���%�$uq׎_Ӧ5Y}�7i^�T�bM�(m:#:KR�z7,r�^�V�nmXż���,T�v�l�1�,h`iH�j��h��
zȺ/�_n&(ٷ��-s�'�ᙩoHr��>�qA�Xz�:�,p[s+9ݷ������Sp��U�$�p���P^Y�1{;�܂�z���<opk��o�{nԤ������<��j�6�����j�vn�����CӪi���	԰�-Ǫ&��aD£l���4WQ0�Tn��+5>r���,�S�Iv���,ŷ�6��N�[����p��pmc]��^[�B�A+Jb��ՅwNg&�����1(o-�踪�=-��ͧ��J���|���H��1�9�3[ݲm��gm�#2��PX!��E�R���Ev*�`��>ӷ+�f����̙y#��T6H�_Y���`a��E��܀](on^��i�/I6���0�:���`���7�c��I��(ތTs�7�#I�M�*�U���I�;�qt�ŧx�ܞ�>5�B�ݽ��q�,
d�mGNJu�r���Y��]%�I�_u4G��ܿ��af�澒�8�K4΢�Y��
�/YE��b2=��L^�I�/�Y�"�i����΋_[��"��{�6�7X�(n����>�I˝}h^U+�U��ff��=P	w����+�޶��Uh��	t��9���U���W�6��Kb}��O%](w�k���o6�[#�D2�xU���nP�gK@V]��n�νNm�x��U�,=s�-���:u��S��Z��:���8�F��sm��ᴡ��ַj��(M�9%+8���7���{Ɖ���r�PTp���FB���>=37p��9�c���'Bê4)��g����w�:_b�j���L�r)��3-	�a���h|wo��͆�O
���5��2���k��������T�m�9��6����oj�A� n��o�H��9,@�ݶ��;��z���;�I����9�������ˮ���ё]�X�}�Y}v�ץ��G��F��73t+�b.���E6�a�,����9l���4���2�ǵqjK+��7wsir�g2�������E�˝��J[ݹ��4�K4���0�R5Ů'F��J��;�����bWX�jە,I��� ��[���k ����*׾:�ym�'+����i��Xªu���[}�(�s_s�{KK���>����ܸR�.e�ްy>�3�@��1��Df��i;�zZ�-*\�#+%��2j���$.�.��y�{ڀ
�uZ���Srs@.�C�6�2�=+K�6�,��&͆i}w׊c<ߤ�U�i�nT�av�A��8�ᑓ�u?u���٦ⳳ��c��F���T/&.�c[%�+��4�� $`��@�}�����Ob��,S�WUf�c��m�9i�������ݔ��|�$�ˑ1[V��*b�r���zYD����g�z�p�䦦�hV�{�u�|�,��mY�ov��d�1����v����Ж�$�\�n��|H9C��t��j���Ed�l�aK��u>w��o�w�Xu]�<��T� �{��Q��+��WJn<�m�)U�V�
 Ʀ�I窘N3��==��u���4���֢ͬgC.Uu:l�[�.�d��X)������R^n�Xː����M�a�����Y�0���Fͻ�?d����� )E̘��V(�5���h���Q�H.O7��L�r�Z��o��M�)d�1��НaR�Ў#!���S13��39P��/r\,��vi(��$�V5m�v��eq$�e	,�ޯ�P���fpUo�f3�L�zt�M4����l���gu���0<�h���;t��_;���n�n �N��
o�Va֫C:����b�^�� �nFN�8n=[�4��μν�P"���p�4�\Ҟ����k)�&"�<�v��-0��.�_v<�E�hյw�a�_^�#*S��vt�x�bթi�����K����=e�kt�}���o5L����'p'87��(`�e̲�d�Z�yfҧN
��vy.d��`=��2պv����Iq"�����5�W<�Uw�:§.+��Z!� D�uZ�����Н[�6�������򄱪}�1h>����ZD�N���B0uZ�ѐ��
�	�H��EU�M�c��a����!�S�.�eM	���ɛ�T�㞓�,�Gz���7TH8��%_����X���.+ ��+5��>P�$���ND3������$�#5́C��L1��;=e�6��!�kR�۾A�(�!�غ*9jB�U����v��E���7D��6e�3S����g�T��е���̃�h�ŗ]��(K#�؛������/"|��w%)6�g�0t<c�� �j��^�>(g; {Lg8�u�1*�p]��ɧ�NX8N�3m�32�.,t	%f���˧�QKo5��=���ld�s�Y�)R��0-�>y�9/��f��j���
8Z]ׂ�@�gK�f4��t������[j�LSo��Q?I)�D��0^BsTqU��o#�?\m8QD��+U�o��7xMpaƂ#nn����7�7W�x�'���v�љ�z�#�_V��WX��i���e��Y!G;�L����N��G�EN�&*on�YB����AgG�^f�L�\E��	KmD��95x%o�()�r��pǮ��SϹ8�;R�N-�8�;L������l!���C�w4k��-��:Պ��f[���z�v��� t#&��;$Ü�'���78��j-�<��w��6���N�Ss
�s�5�5$s9�v[�'=+oyX��{ZVHغ��]:�q��Y��+h�t,B<����{����x�@͵d�{n׈��#��{��a5g.�Y]il}x�/a���9)O�B�K�Фz�:��0ګ�"�X��j���$�m��$�R�>4,1I"�C����#ۥhw*�����f�\�[v���{5³yD3���H]1�Z�6M[R��X�mV6󆱂˻i�T�X�D�6>
��ґ�y���4v�cUm(�Ť�3p�B	#����:B-k��P�.,e�}cM�г�R�W�1v���`Z�n�(ԥ� =�̺ާ�]��E��E��1EO!ǭٔ%���U�^ v���@m��ޏj��m�z�c��U���nz[ݻ��-](�Nj�N�<�-Y��=�pW��_�{q���T�%�� ���]ѓ�m���b�n���u��Qz,�L-Ҥڵ# R�:�(R�lS֏n��yx�7Ϻz��x�[�u�f,�������BZ�v��p1{���19�`y����W�W(��j�w���
�ս�®�������Dw.��i4���7{x�A8����{�����2Jth>��"��n�����5�x�fK\���Um��OKtʬ��٦��Ԧ�<����|t\�R��4�Y�N�ZU�d�T��x^����������}�p2
ur�F�;P�[���vTwA�R����Zw$o=��T9���˚���[u��+��M>���[+{�:WYJ�K)����h?%]2�^7K�+!kTĖ���Yk���k�ώ�ɽ[n�h?�yX&p`fJt ��ʻ�Q�ɪ�Tghɝy���A�ԏ!t��Kgi�E��k�{;�_U���0�
E�#��pɁU��0D�>�t�W>�X��F>��o�mA;]1]uʷ��^e����8y��nWs�<ܡVn�/ҭͼv��,��R��hڴ�,�T�B�+�k;�:@�R�SuZ�a�8�t����LkS�8��yz�}GB;��!�]5j��;�<&v,mi�կӳˇ�8E���ٗιIؘ5���>�"�j��;�1Q��愄�x��*���mer2�����۝�����a�{E���4 �j�ƪ�2���So[x��;�0��tBXG��J�u�$Kȯv
7qTWe|��TN��%,!��,۔��g;,�a�2�]�B�B;8 ���û �\t>�g�q�4�5m���H-8]�/�	�Q���n��Fcwy�*jL��{*�8���Xπ��n6�nz!�����h�Un�d�R�Ѫ��Ķ��U���}1�9��M �z�2���6hN7]��;9{�t�w��]�A�(��E�|�=�u�]\��0=�s�g#�̔�ѣ��O�NH1��n�ڼ�m�9�Y7�SǵiE���P��E5V�,����t�ސ�KuQ���]���l"%���uc{X��y�,��J�h��>F�U��T�ʝ�M�Gˮ�b�:{pDNb����2q�G�����D>� ˇjU�e�.��l����ӡ���H���)[����ڱW�/���\�J��@� �.Ӻo*��#�}�l=G5��aF�|��N}u�Vz��)���XÜw+%E�Vb�0���z+���SO����a�0)ז��Q��.��Q7�(��W���nJũ��\�T�4��{�箂��9�������	�	���5[�Z�jkj�a�X':r�ki�0&�r���]�L��K����쥌�ta�z��]5�U�,ɑ��khX�R�sN��KLT�q\�R֋�y�tx`���Zbk��$����(�[H?p���`�H�>
� u��JY���!�njH�b����Xx>��̜�S:��ya�[)���>�S�镛o�-m��L�1c��V;�tC�0Z ��c�%��U��W���O�7���u&Z��wx�������Y5x+]� �U]�޼C]�S%Y}�,�+6NS��/���H��"�n5r�:8;/�-Y���v�EV���ӵ�ܥ���Χ�E�CGG5^%2L� t��M���Cbd��04*,x�v<�hVu&K��M��@n�Tv@��'*`��ƶ�Ge��j۔*ɡI���<+Q��w��
�aUB;g��F�^�P�Ϋ��Z��|��3d�XqV&|�P
�uR]�m�Vr|�����3�V�Mx�7�sN=��AG�ͼ{��,��[�>�*«��^_R"�1fӽיce��f�f
a#��}B��T�r�B��j	�E*Z��#���	ܾ��P*ի4�_P�3�1����td^r��e7u[^�Ys��l>i�^Wp*'1�z�ڽ-
r�˛B��Q��&�V�2�\���wV��	B�,�9m���ޜ��f����_b����.U�W^��t��C���PD���`����0��ǵ�}��81�Pw�RJ���5b�b�t��[���x)V<i���@�[���·�{T`}�s1^���
�䩶�1a�Ly]�n6�tv�'5�W�_G(8�8�wݗ.��9]8���'�g�HǏ��J���u�s5��b���G��3CH�Z���P7cD�RQКJP�hC��	�T�5M%)BR�]�II�颀(�ZSK�֗lv�Ji��%S@�P�Et!�)�F������T��Ĵ-]e�!���:B�֚�t8�:�C��Q�CE��zN��:t���[cl�Š:4�փ�7`�롢�:^��Mz�=��t=�N컱@t�v]��K;!l�R4���A�Q7C�-i5�JշFb�"�[�Rh]��v��t���:Ď���Z���ERX�M�b)zh`�ѡ�ׅ���WK�f͹�6>$��֍�`+F^n[m jT���(��h��GN�Χ�J�F�U˩+Z�Ua7��S{�rEm���?⫦��?<˾`�K(�������T�Mp�6���w�P��Ї|S����&F��P�C;�F }������������-!��گIki���QKoHm�b��77K�ʜE:p��ٱL(/>�������Gş�ibc7�lft��![�Ƕ2�:�3el�ab�S2c!�1J^W O�����w�C)ݪ�ݴm�9wz�S��I^��՗���^�\
v��Ҽ%W ���k��w���.�O��K�h��,G<ߥ�����o=�mu�5�~��Rtǭ�/�	�U(
͆G�O�Ck��]����J�%��)�ִ�4��>ɳ��\傽*��e _�V? )Vro)�s����fs��.ƌ�+�]Mj��=!�k�gӎ���&/)r.E����#��0@ЅCZ�6�=Z����Ue����o�{���;^�z8s�h��.�������KL�AnȆ��Q�h�OqM��0��w�Y��ʼ骮}]�G�e{����Q����as��n� ��	�zu$O
,��!����#ة�t�������1L�},���32E��x�)7�j���H���'��������k�|��׼�eU�����Yw]J�����B��.Ҹ݅�&;4�I��9ň��=��:���.����:�7_o.0{�V�J�_{���AI'�:��NUk�[� ؘ�9� f��펡���W~�/��}a˻�'�^i֖��i�܏^���;Z�K!��?��l�&�rn!S}䲇��}�*�����V��/�n�pk�0�� ,�Z[I՜�(���{u��]������dLxԡU���&6Uc�݀'r����w���I��5���Q@(�|;�E81͙$phf�q\됵�:2ݲ�٠����6U�鍆 X��z_�.�bo5�&c.�#��h�4���ԥÞn�h����@�Mp�~�<� �h���*�mdV(��:��!�
}v؎�!�(���l汁�#�㡦&ym�#�����q5�U���R-vP�.N��
Q[)��*���Z�1���T��cF�2��#�@�잭�~D+HW�,�ci�;�\</KD�!���y�^�!Sj1�'�
r�ΒDG��8�>e,��Fj��8�>  �|V�^ Xy��>���I9o�����"oz���{������Eji�\YI��j�����+�HHs�TG�G+3���^ڼ겥Nݲ�*�M�{M��#����s�gb�ty(,u�妣�%��3}L�K|4���,�������y�X9�c/��r����u��v���3|�͒u�s�f��:�'k{ ���A3���u�U����ԣ��5��-�3y|����R��c��K�@$ͱ^��۞���U�
jg��_��x�V;�vz�±�}戎���M�l�)(h1�T�U5W�cFL���a�c�N�}�k�j��Z�|:CfZ�X��-�~�x�t��y+ |���=�g��K���ԅc����p<|x{|��u������F�Wo���M��M�c7��=�e-<����:�B�}iW��p�^8;��M0�����˼g���xqLW��Y�=>�K+%\��l^�1Ӗn�Z*�*�O\]��>��V����:�Kŝ���R��)C}��ʻ.Aв,>��{����@�O�x5������+��ܟe��8��?z�fwSo�	n��ي3b�n�{���:p�>�Ht�(���r?6)��O�T�r�C�Gҷ�<Kr�)���L�����wR��^;}{�<υ�5ࢥc��n�@�X^��[9,�d�r���=���֌�*,�5�XD�㵝tq�mS0�W�լ.���Y��{��y��[ٗ���_Q��}���7:r9�a���]�kV�Ӝ��e���.;��q��u�J�����M��O�fbo�egƟt���O��M�z50�c�3����.���w����o�@�kc�ru�wk<�]g#���
�\Ȱ�OZ�8�]��PYA���XڀS�@c�Sϛh�d�%2k`6&�Va�SU}�`\�j���������
����CU�@o�Mz7p�w������ݖ���l��W��!��{'�+����^�EZ��u�>����Nճ�`�a�!�}ǁm��ό�!���mW�ҔpzZ��}U��◔=�jާ;�ٺ��/���U�ɴMqW�	]�k�aB�w�c�i#Pmx����U�E�U�Im$TNܴ-ԝm���8�y�a@>�3=�)�e��}�B�kzOY��2˯thWv�'�ް3Wo(��n��W	��x]f*a� /��h{&ƀ��A�J���E^�b�},�'S�+S��vj��5g��n�����~@W?�!��Ɍ���k����1��U7�S;�-���d�A����#^R0i�T�>��n��7��xo��\)�&�B������`^^oP}٬�5�|�xJ�/ݍ
�~d>�����f�NuWU�PQ�Z+�xWaʿlumT�,�k� WofvVEL�P'�r�)L���O���t�b�z�"���5lX6w�wd᢮Z���Y����z�r�Տpd�a�y�R6��my��{M�/W����R{��u���0r��W�bw/ҩ��/��ግƙ�m���W��a������C5Re!�PA�����܂5��z!�ќ��yK7����[�9̩�x
v�&Ҭ�����g0���,-a�^�A�֛~G����\���ҽ۹�u��O�l�����ٜA�PS~s�B���ŕ��Og[M�Ll�F�N[Y5���ދI��4�uI*��0=����;�+�X�|b�5w@����G	���]6l�6��WS��Rs�yx�d�3:�^i�X���p�[ukĲr�*�J�<������_f�t���-��۷��1^�d ճ W�iK�>w����ϧ�Z�[�m���!�z@Q���p���j*�t5�^��|�8A����1� 4a��0���@G�ĸ�4��Ȃ�n�yG[�(
��%ݶ��
�2662y�,���Q�؄7���D�gXZY����ۗ���%x��	�k4T�}u���Y��gʐ�z�h�tS�2.6�T�ke�Ld�'�M�X,���Y^ڸc=춉�y���
���xQ��]j|@y�~v�#�����3UuGm��7[�L]����ɪ�]N��μ*-&�>r�͟?f!i|�<8����8,Y
�<��<��"fE�!;����|��˧��G�-H��Z4\zk�}�_Q�&�6:.���(^���,)�ɑ���K�tM6���FA�a��.�'��%�ŷ��xz�{p!�0��傽mk88~c��rs��T�W����6��.�d��y��Alϯ�W{���^oW��#��/�CW����(�u暻���a��#n�b͛贂��B��j}'֮�f28O�+����S괰��̫Y�1\-�v3����Sq�D��+]�e8�#[�*���}0ϻ� ���֫��V�\��b|�2/�ؘ���e`So��f��"$�,�*κ��O��mr�B�U(�ǵ��]ѭ�%]c���:`��@�o����8X��_h�>��{-����zȫ��d�낲�#Q��l�D&���������0$5��E��*�`�זa�o-�Ж�v��bw�^]r�����c�f݄��VP�O�5[أ�b�?]غ�o�c�����sX�a�hf�v��X�,��A�C���ND�P��hmE���e�azcbv�)�Z�R�����{��l���1�m j:�]8��\��`�@v��x���Fw�H C_-��,��"�Ou��gm��.s�+=^DbA�Q�����z�$e�Yo��fE�ҹS���
��1��j<aa#�r���6kF_>�*�iv����G[I˲��f
�qu{\"���7�y�0�8o^{�
��5jp��:q���[�.�ܩ�r��5�ْVU��O.�ɛ�69��[SoYF:�v؍�2a0T����N@��4��vi�c�Q�T��`�7g=R��O�`�jE�<V�O#ʯ�� ��j�E%*�FT��~�7Vy�>�bC]z��W*��KI�+]�)�청�c,���c�Z�N��@m̞��ؕ�p����>C*9绹�Ii5|���ETuLM��Z��E�{��w*��n=ƹ��x�[�{�Q˸���^��b�0�c�*����9[b'."H�;����e^{�{w���"}��h�Sb��vu@z3�lG��:��EQD�{�_{G�z����϶��jXa�N��)��j��K~�"F=�B�?^���w~� "�;']�������:��3�K���!W�{7C�l'N�e�%�p��S��ۻ�o�I�ޑ��iR�AF��7k�y�V�puQ.���i��>�W���̩$�"9Ԡ{��7�`l����s/�����E]^����oV�
�i�z��T���:��5��g�yc��Rm.�G�^S�9�����Y��Y��[�f���7���,���`���-��qW�͵��e�#}�c���֗j�ً�c�	ջX�����m%�:%Փ�5ٍ^}�AՑ�GHo�E�c}��Oy�*zB�p��+��9G��f7�1��8�98����m����.<��)	_m�ǀ�o��8�Z��������w'G��]��o�VZ͊��$���2Ҥʧ%
>�Hu�q������b�b�sX)34�R�������Z�'�Vd2�=��+�`���F�u���*U��U6!aMt$5%iI���6�	L�ϠCU��-��Z�o/[^5\�$��r~D ���*����vz�nq"^r���|��aЛj�N^�t|>��/�"1;���­AR�퐴M]��{7*�ޅP���n��>^��ћF��
����7Ƙ&�����+�^�,�z�S��-@؝���*|g��m�t��PcE�[�1�	�6�ڷ/Z�u��^%wWRc���>��i������q�h�D;p�y�
k��������j�����z����*�Ky+�@� Wg����7��{��Y����k��֠�}��=O"k�;Nc���xX��רg)��.n�a�򡹜��<��h+}�v��rX{��;A���X���SB�n��Ûa�����Z\����@��3rgWv�����ڬ�I��|��0b�ƅ�),���RF�>��A��/_�֠����U<�z,�h�>�äI称�y�M��o��]���K�Sy[z��k���dh��B�Q�kJlbi�}t���Rw+m�j2�NI�Ɇj���-DQ���С	�� +�bC�ʬ���?���7H]ou��y	-��ݸB�����V����|e ����)�%(H�6��z炙�t>�`�w:^K���w��5��s���=���z� ���y! �N�N��ygKO�/6B�]N�4�!9Ѭ�V{�*x�<����'{=u�zzxK�����aז�;�,����׆�>��k鐰=X�ǅ:�x�4Ǽ�6sf�;�Ӂ�C4�A�aNtc�u;�*Lێû�r���o��-��U�؂�o�h�D���
�{�k����\����gd�kȹ!ӂ���f*Z;o쑌�X�Q����:[ݝ�n���ob5^����]`����#�ח`_��t����U�=�j&��rϩѬ_I�n��&PUg��|�"��[-����Q�a��`�f ���@D���}�8�~���H��=��Y�-U��s���S���rn#s�Dw;=���"����#�z����W]��+k��>I��[z��9��1����,(;Up-J]��F*Wt�]�����:;2���k�L[m�P�k��5��S г ;��z]�rPj>:��Iqs��jԾ��^��v����S���WS&���69�h�{����"��o�':�� W��,���� 43i�v�	�ϡl�}�饯~���c��A��^jj���2v���k�E��
6{Z[S9F�!L�0�h������6����;��OS��̜H]gٔ�f�+�~�c5o ��R�N�vj�tS�z/�bG���6<1�{��2w(��f��Է%p�ZS�ЁY�>r�p
�> :�[���
wT����@,������G���E	J�MӜѳ��?@�
�������? )g )j����xe�6-��7�ۻЌ�M�Q��m`_y��{���n�bb��b���%��a�S�A���/N��vil���u ,,�^���0M�1�]91�ޅ��l��h�+Uֲ��T63m�p��s��[o^Y��ݟ:4{yk;S�x1�U\���^��z.������Ǽ7�{V?W�*��;[��є���Ƿe�@{)'�7�Y*2=UL+�t����ϣ}��ck_58�@fz�L�ۨ r-�S�]ƝBǸ�nG��]a�d���-l�l�b���#�gY��l��;���jrDc9FvW;���M�������av}��';s8���V3H�]P���:rcG���ޠ�m���W���8y	o:�}�"�t��M� ��\���Vo����B�st�Ǫ��e)}>��:�7����rɔ.aw&�=��o�1j����vr����,\�V��ʓv[(̫�	t�J��A"kix7�!4E�y!\�/Z��E��T�G�3�'����y��h��i"3����Kdg2uBT��
ow��s���\�n�FçO�ϭ��O�^& p�\[�0v����Z��!��5矘Ə]�[��6��^�ո���q�J�Ҽ���7��QU��������f�KWi�(�3�R������Y��8֭�p7N�6$�AڝXn͑Mb�h<��J�����V�}�h��W��1B�u0����;���p�&ۧY�D{w4��z�)=�D|5��3�S�{;�d�[�cc��r����em��uͅqW�w�OB���n���ڄYYޔ�dl����܊*:�J�<¥w^�3���J�r�m�Wy{�!ƈ��kiM�v-�[o����$�0^�������.���L\��7�	G,��h,8{��)vrvg��a�Ϗ�J+�l�#��i�V���uns7zFY!�f���\��v�����O+�C'�cU�P�".�k�X�1�n��z}��A�fe�L�]���EX�4%�غJh��2���0^R�<]>�l�U��T��u�e]Ez��nHWRv��ɩ��c��6j��1	�X��V]8��P��y�y�s;u����Yu� &4�{�SƳ�x���~����'�rZ�������O%��9��z,4T{y��"�]̝����Y��x�]Ij�ˏ��/<70�r�^��n�5��ʴ��:.�eu����2�Tm�wr����H/4���D6��ݻ�3�]�H���$�%NΎ�ۺ
1��wN�:��1�U�N��b���0V_
�H8P/����I�.b]y�kwhPG����m�N+܆��2���|�pFB-�f� �T��a�l����ʀ�]��_
ɡ�Y|�<��ʍHzk�AZN���.�|�b��p�0�� �W<�V�C����qx\��䆲U-�T7,��]��;l�n@C�j\E�"��ӢOVeN��3�{q�P�o�.�'��ٵ5��J�Ք�{y}np�gt���bM&1�
qC�	u��@�Y��2��s���z^�]�Ȱ�ʥt��Z�f^���-��>�����>�ԝ
�e-y�#�og�ˢP�O�#�;ӂ�a6�^9[�]oo1]�u��V���OmtW�������|�,RglW��"�͐m�{�z��f����ɵ��I�/����!·�J9za���w���4�zt���A�1K�$z-�����wJy�)|1y���n��(��#}P�y�:%SwWҙ�]�롱;���ך�տ-��{��@=:5ٵc�ݸ-���wں� �I�I�M`��DLI�Ļ��t�(h�i���#A�ݸJ�j���8�:�]!Ht(�i����QAZ:�:v0tih����+C��3m��gI�F���ӱ�k�4%u�ꍱ�{�����;[Vڡ֝3RF*QV��)�Jf4�"h"i�P�2h
����hӢ���Tb�F'[b"�N�4�1.�:�
�[h�F�Ql�"�ڍ�M-%�h֍V�X��:�uj�Y�ݢ�Z&�؋Z�Z��Ѧ���#EU���#�5IX�m�0AA�1�*v�E4Q�ն#X�kA�*n��"��PVګLcTN��U�S�n����]d�
�[���Kj
��>�+�(�D
�����pV�lð�������{�w\YA�P�a�ʇu��]���6�ɼc����9{���xo�7�h�Pg��c�CHd�<��.!�}���`�����|<�q��i��y��������=����C�C��Ѿ���׽��:�h�|���|���/A�����1�k���\׌�G3hg��3����4��~�|Hy������	��z���|�:4?n��}�R�'��/G�܇�̆�ǯ�{������;{��>ψ>A��x��Ӥ�)������Zُ��㙱� ��}.�������x����z_/o��ph��>�����O�u^S��^ ��4�wrkA����>`�~���o_<xi|AA�7���HS�=��w隬����5	����`ԣ��w��C��'��?c�u��O�}�>~|��h�	T�c�t?�i�}�~����N�>���2����y���4��=S��t���4:�%��~�ޥ��7p�zk�ydޯMK��zI�Wy�z]'����4z���!y��������e�>ïpy�ϝ�0����;�_��	_�B!��OO������Z���{�`4i'��~<����f!�n� s���q��S�v�<sx�A�M�w ����{�o��}T��@~�G�����/E��{�~��2t?�׹��n��>ÿ���'_�0�����C�������R0<���Y�nz�vz7r!�/-��fF����	Z��>����<�z��v��?O�=���<z�P�C����q������S��^������4u�/��cI�M���C�f!������g��t=�j-�*;%��6��N��� �A��8��w���{̺
���{�'������z0��'��x<κO��?#������%?��u�2{�q�������4>}��쟠�>^ ���`>ƗN�������'	қޮ���ᙤ1����� z�xïG߼�����/x�O��������>@�ܺO_}��<ǉ~]R�;����:}��u���C��׸��rz�5���>�>�5OO�A����nj�q��4����L'/�Gh���{q���:����/�?���K�c������5�����~�P}�G���Py������~T��K��� �u�=���|����6�_�������7�k�t�A�ֶٓ�E��Ͳe�볓g��%��n{�ׯsȬlm�X3~��e ���<'�(V��t� A����2��aĖC�W;��Swo�Rq��a�3��M@E�ኇC�
Y��+G���}x�zzqP)V�E�7o_(e���\�SqN^�w@9厷��:��VC�HUAU��6@�~�BW��>��4?.���/BW�=�����	Z����A�<@x�|��Ǆ/��������z���|����t����+�
_��|����E�g�S�Od�FRo@fl� 75K�Ɨ���<��d�����}n�������Ҿ�{����O�?�8z}��CG�x�l��7�B�y�]QUi^B��m��ws��4��b��ƽK�:~ǈ�s��it����~���1�ܝ=�t����~����'��<�������)�=�=A�{@d=��׹f�!]�G��=�t�38ohf"ǽ��%����E�������0��^��(�/��t>O��x0���=��%{�����A�F���'���O�:_wGC�'����oHf����Mݷn���/^w�ϟ}�}���:O��~G�>C���Oo��=@}��;׏�����i�����������4�>�o�?eѡ�u_܇�J�>~x��z���'���C!������$�GF�*���_>�B^3����p��0�g����?��}���4���߾p:Ph�����_PcO������:C�<���i5��C�4:�}��͞�zG�{�3 ʳ������n̮>x�������C�m^��~�kǬ�O��׈?�x����	O�=x���?��:C��t���A������GA����'���}����~�a����=�=���y��Y ���8gF�P|��|����璃C����Q@S�]z;��c�_wO�����'��>G�䆟���_%������>���^�ǈ=���?o�}���3�~�;Z��-�����s=����ѣ�}�˯�?��=�|:<�}�'���t�ow���<T��O�Y>ǈ?C���):�h=A�~�hA���/�;�C�Ӟ�#ͣ����=�ݴs���gܺ4>���޼P�%x��ׄ�#�%i����0~��:_G��<�_����?z��x����z��|A�<A�y����h+�����y��po&�H#ހ��1��^ޣzζ?	u�v��q��ͱ���q�]DJ�Zs�|���!}~BN�eW'x�}og\�Av��,��i��+�M,���i5�k��YKNY*�4mv
v�̂����D:�wm��9\s���� ������5]�����4���/}��A��?G_���:]���7a5I�����������y����'��|���|�P���������,��=�Cy�4�{��6N�u�y�^?���O�t~>}���OPѤ�=>����]:��;������A�����</�=C���?b�@S�O���M?���.��|����5�z�-٬5f!��8,��.)4�^c]f�&j=�%�y��K�h��>���>GCt�K� K2·�6\Ph�����K"
�	MU��+4Ӗ�Q���=�ۣHg�V��P;2���)Pu�v�V|�y{*��:{��xE)5�^�<�'藖cnp�w4{ۂ�q�m[�|.�1|@��X��M| �����9�*�+�q&��w;��S�﫽��jP����r��<9�.�%~7�v�$8\�3��!�.&���&|�md�+�|f�p�m����F,m,a�PB;)z}K��%)D����xo�R�fQZ*�7ږ��EbɌ��E��-J64!>QY6+�lǲZ�-��נ� �e�F���\����.��*۔����u��L�^�}a�ý�'�Ӆ�q9�DR��f�W���kq�A�����Z/�@��m4IZrK@J6sf�;�a�?�(e>�P�蓐�Dbl�rlB�H�%ܓi=]�:r�d�{5��τ�h�Ƴ&֗�����o)��
V!�ǽuk�c�����'IZ��ע�K}h79Q=��9�ԏ|�������:���.Ö�:��pJBBH.k�춀gɊ�s+s�����)�O��lt~����u'Y������=�O~�+�K�L�[�~Χ�'TM�'��'ܟQ�X����J��Q���Z;��c�a��i�C��x��?c�]x������]))�������:{2�P�5O܇�O�e���v)4��A^���u��K���F��N]!N���(1��@�iW �~h^o���x���#=32�4�����k���]��bi� S��֯�̲���|g?0)���̩OX��h��5�ڟ62����n��g���ٱ�WP��>�.�8u���>�Ʀ���^ڀ���h����R�v�����Ƶq�uh�%Wg��cVy`)��1yׅ�
�T���+��Ľ.Ğ{:���B���8��w��f�yu-mg��	UiL<)��|�(���*������yy�Ǽ�k�>$E)�L���/d�����N�/pב0��A=���k����0�9��6IQ�n�S�T`���(��X�ϻ�U{u��.��Z��"��l������.�_�~w����gqt��l�FO{m�܋Y�E��'I�7w=!$h���fg#�z�)f��+��jn�}Vq-��s�x�Y!"����V�Úl�xNQ-��ݦr�}�}6�z��3���ʸ���7o���q-㡰�<���9�ϲ]��窄��Fu��_o*�F�'M�S��j���fI(�K2Jn�{�㹯b���KG��0�?��-?8k��+
җ�=����r�T:j������0&�s���t��!�蹷��;��
>��݀��-^�	jwl
m��q�D5��gKg��	�v�6���ի+%\��ؼ�FɖW �ϛ�V�Z ��ϭwp��3{c�z���|�H�4`�e�eƺ�`%j�L�
=��n�N��[�8�m�� O��V����X832�1��x5{���!�ܻ��vl`Id8�,������
j�V��������g�M�,r��&[ѩhO�Keh���be����<�y��
�iܫ��Ǐ	X�W�U05Y�WwZ]ޢyd��ӆ��XS��`r��~cO�G\߶�ڮ\Jwb6=]�Ⱦ�����k}(��g[��n��~u;�]P<-ְ�W�U����)��F�ݭe��5���Qx۳B�cڍ�� 'L��ªhR��Ɗ<>�2x=Cλ�q���}��-;䋸�#ӥ�
������u���wC#�/�����5(E����:I��xF,���+8T�4`e�g�Y#ݽ�7���<:�Wb�����ɮ�%��R��ݏ�d��7s�P����oY���3+n�2�{yRC{wh>�?>��nPД����-�nO�Uf�}j���,5\<U��S��ZS�{J+�	oE��`x�e׃���e��~�VJ��^�r���v�EF� 7X�����ԟn� ���u�W�u���y���yT���S�컈�{��y��ͫ�fD\8�a�uw+�{���ƪ�����3�x�O��h�Jb�b�V��b��bT-ܮ뺷��S	q2��-{�{LVc�Q~qe�yM�0���N��)׿j��J˃�(�z��%;j�H���xj�W�TP;u���L ɜr�/i�ԅc�����\k��ȚN���3w�q�9_����WS�x|���
�v��]��#m�U�ĸo��i���t�z�V=V-DL,aKN�\�e����W����;̾\�W^R�WAzz����xV��R�BڀQ)Q:/Y��h�c{eߔh��[Es�HZ��PZ���E]޲��פ�f��Sz�:o`."���T{�8�t2�,�=fW:p����,�;�
��Q�W���,�w �"�Y#b����%�;��15�5S4��wv��%��u�s���,/�^�Ev�B��Lt�vvo�~RՄws�X�0lgeb|�G-a�H���|jK#y墳���y��k���u1)��b&>�:�u.��X�N�kc-�X������v8+�\��B�	�]�W����a��ʴp�i_�y�/ڪeIBڜ\��|f�n�6���ټ�V�U�BǶ�/ӟ�_�s�5]㵘�zU%�UJ<�uO�ʫ�vƲ�ͥ��ng��qR��y� ?���eyR�Y>�l���T���3.��b�+��m=&�L���	+Ukf�=�C`���u��^}�*�U���Q�~�Z68W����jR���a�ָm8�Uv%�@b�8	Kc��04@-th}p�O����ǚٮM�)ݷHy�݌��kGn�V��h:Zl���'Θ �>��3i�����޸Gh��C�a��@85�-S�R/i�7ܳ���b�|�ν�� go�������i��{��յ.w��<���s�x��M���P;7�/�kO ���%��B�V�y�P���ӂ�t���K'	rۤ���FEgZ�}�s�Y�2�}1��� ���~;����|��|�̯$'�X��w�[��E�>F� ��J���ѳÙB����ʿ +���0�x��^ՎEC6Sn���ݫ��^n @wJn�1�z�}�G�%�ҧ�Hc�IJ����C�ڝ`�ʻ��.�˙�e_7|(�g�.�����g�p+r�U>�F%x���9�2TU;+*�cyk�
����������vI��5;��*#u�X��bLg3�^������5�>cι���{�ˋ�m�PB;)z}JwIJ7�����L|,�����o}�����S�L:�-�X�p��;ف߹�[~D.Ϲ=�[5`w@��]FUؽ��W�e�B�ag+��8�����w��W8����M[y`&J\;�������5��>�`:XQV�
���Ѧ=糯t��`ի�}�������nVLmW>��t�Z8=��[�1s��!/�6,�?��/q�x���a��������`L�R�#}�8-_dʯ{��+���j�R��o#'��	Tb�5w�<<�����Cm�>�|���I���m����s�6<���G�K�fH���N�bǦh��qU�j
��^Su���k�(d���Q�g���Od�� [6��<ӪH��ѐ��Ѻ��-5�U��;mW�R4���K�Zu������Ŷ�C����b2�P�-�vJaAyf�����s�1�y����d��#��I���?q�+Z����ι���5;ԏ����~^n�s�!�5���������tűww���=x��3`]�9�G��T˅s�"1�1S�i=�C��;��^���YFJe������]�P�Jc��kS[�P�]6�X.Ա`��;k���]c�69�e1q�Y��eNw��<1�mk�����?���&k��s!m9b�L�&�E"F�S�A��>���W��^mU,�~>M�]��0$^44�oy_�Lm���J�׹��U�Z-��J�iL<,@����Gu���pR��6n�����`{uп.ψ
���T�xd���cҮT>A� ���ֲt��6vV�� *p�/"�z�XZ-(�pj�?�5)8#��hL;��^|8���\����-Z0f).ϥ2)��h�kP�h1�
�>��0O�\>򻃥��b8�ǎ�ޝ�Ǻ�����0��Wsj�}ia���PW�˖�u���j�u�Ư��V�ɍr��K�&��{ �����`^���Uj��iV�M��m�@��|�Z�a�������\N��W�3ѾN�ֳ�7���z6l�h 6w�oֻ�8X��������F��X�B��؃{��R��L���̤��P�Ϟ�4j���փ�Qxv�.���mV�-z�U��6	��L�k�BY[�A��T'��k.4�z�6m���k�
��b�����{�h���]C��[\��3���@��8��sś1 7�/bU�ge���i)s̯~��z�4��o�?F޿�t�mo���S|�]�{┯ڝ�t.F%GL�(I��tn����ñe�L��^����G���zN���}UG�Kq�%�����Z�2�;���n�d�<�a�jx
�p���D46��il�6��@�I���e[4&[r�SI=ٲUkY�4�!��uί 7k��<�<���l��B���8�]�=]�_
X�["Y��=�a�F ;n���l�LZk�����z#ӸI�V}*�M�5�S�e+v�+��1C��X|-֦O!;C��:�P]&�سq���O��K�=U�d�{��-�����vk�׬�r�S�\<��\�f��v�n���@Mn戬vD�2w�k�yd�p��lLg�y��ߝRX��>�����~����6ͺ�ƀ�B[��
E�yT}a�4<@�yZBysyܶw۲l��$|�p��G������~c�j�`�B��A�Z0$=��k����ȼ���}���V�q.�b[�=�e�[�\���U3�a�U��-�yҀ��A�N��y���Ë	\U=�~vW��s=��� ���(z�!��u螴�+��\5�v�����*�J�@'��y�N�No6tK�k�|����u���Ϲ��#��AY����]�0R\l?Ns)�BD�90�z�+��PP��^�;��N�ܴwZ
^E�R4`s�m#{��n49�˕�IvFd��]n���%�q�5������Yz�i�i�>w#Y`�@�����֥E-��r"m�]�ԍkN��;�q�=���+U �<����>ywN����/xv�����8b�:�L��6R3���1��s�q�o4������k6����&5���K��l�Wa�^�n*�v���<��O�Y��������TZեY�r��ܳ��=��/c��7�wGw�:���2��K�dѡ�l�7��>�{; ,���aea)��K����	�*�V��5�t�e�+{Eq8���l��.刻x�Ijn�}tJ��x�)5Sf]�w]1Dγն���--��,�F�L�a3�x���L�Mi�'�Q��t�k��G
S-nT�&䫮���OG1>�4�j�Қ�[��H�h�L���2�g��f'Q��M�Z����j��.����e4����:b40%	� n��d�75LLZM殠��� �Ul7�\��u�X
7���[k)�bVJްa����em$�ug8q��b`���:��J:�oT�r����WP���4`B�����p����H��n-��v\f���7���2��晾��<n=����khY�^�c[�ڝ�����@+�S��`4o��8x��A���e��X��'W�ZA��>r�I��u����zv��y烵+e�W!��]�p���݂x3uً&G�����<�*���9����U��\g�D [6h;���+b&t��
�f�>Y�нΫ]�m����˜���r�{�uQ�$�����d
���P7M�r���i�/E=묻pK�ib��fh�̣=�L���N��C.08�b��
�ܭ��}�����zR�3��P>X��tř�����������}����R�P���Վ=i�toi�gZ[&��jE�=>U16c
�0�^�G�v���� �&��9SE���>Du����1�AC-�:']��#x_�Fv�ih����s�u�v^�om'w�����s8��A�ÙCI�o���� ����b偌���5��x��}� �� 3',-��<>�fԦ��ZI�o����4��̲g�eV��n�z'��}��w�[�6ws~���H{���8Ӗ،�͝�<nLx�j[����"=!m��8g����<����ܾ�$ �W��'l����f@r�V�����sXZ���
*���[�Э��ӊ�w�7�}1u�F}�&���#����)�݈ӕ�D��΄_$���8L��J�������<Z~)d��'-z,�}�U�!j��ޫ+��v�&mY�C���ܒqME����*�'Z�14�P�%�5�b(�.�T�3���1�Z
7mt�-�ul�Ӡ�u�6tth� �*-ֳUQ&����]�V�حj�� ш5l�DkE�v��[��8+m[
I��)�7X�Z�4E]�D]b��&�-bӫch��v�GmѦ�c1PT�4mZ$��X�����Q���8���X7c�
�#��J	��:��lX��b�$֓�QA��i���v���AIT�]�M�lU[h�&��sc�j�Qj�c�)�AE�b����6ttfn��DIV��:�-�k`��mA%;un��K��n�h�7ml��Mt⌧4RDWWc�㙺�b	�{�ͩ̔!�O�������ُ{S.a��%�[g�J������[x�y��Qݡ��{���k�R��:�Vln?��k\�ܾ��{)W\jq���ֺ2Ү�\1S\H�1[!Sn�	��2��,[MAy�zo�!��K�`�`��Y+�e��Wd��j`�R�@�9��d�}X��s�R+;�[�Wy�3�hy��r���"����t"��ݷ�~b���9�rB�B�ӯyx�jK��ϩ�-z��Qxo����V�O=~�R�P���p� ��w�{��7�7�(v�͊r�J�S�����K�u�c���q�����_��=χ�o����&A$�Gm��*U���KGbT��OO��s�5]~�4ȿ�ɕ�v�vY^>k%�9ڇRm������ӇO�eT�GSA�@ϫ�.�<�xVO��,1:� ����r���u�Ch�����}	��J�v�TF������:ZǵD�����G���O
���q�ِ�{����y���f�a�7εt��� Q��dS�#�]"��j*��p~����ۉ�Y���z)�6��ܦ��1vjvH�C�M�� �>��6����0ܠqVDDG.��[�r��S�q;E�V7w�Rc��뤬[xJ9e9e�O�� ��l�ܮW�lT�6�� ��]��r�1�f`; �"�s�h��l��v=�嚫�d>��P��L+-!�z��)���:ۇ7��Ç�Z�\^'��oC���9r�N�5���w�U}�UzInF���'��٧��5����,��C)�K�i��Q(�8�5\Ђ�j������Z<���E�k���୿Tx/�ŏ�ʷ��KP;7�_����䪞O*�Q�Oe[z��V�*]�>�=K��H��DU�t^�0�_ي�w�Z�Or���z���� ��''ޒA{u��z����qN#��]y�%`�u7�nІN�q$�2���a������e�/��٭��#)�&���g�TU2ܟ`�k��o�k���vR���N�)U�,5�z��rJw�y;��p�=z�1����IM�`�Wk��>ǵ��ʭ�E�,���'����e�W�2�5[D�7C�~�r���oi
�����aB��NMSՁ��RT�__5b��/�^!�~�=�mo�~������CzN��b�͌��ٹ0���xi�.�� �v�8�V
���|O^�#H/�}���F��]E�;o>�+�;�u�n��j��SR��	�q0Gz�|�����mY��2�R��t�1�}栂Q���������������cWf!�6F1�\﹄�et��S}�j�9kF���9#%�l��u��lf+�)�� ���C�6�E�W}�Y���Whx8����s9��bw>������Dx)�*=��
ˡ������"��'���������d��q#f��緰��P�rT2�U��"K�fZB�Ƨ�#,�4�r�]۽�	�s�V+��Zo.��X�A�$�2��:�1���ڪZ=;J\	fw�i�����[x�o�Tf��]~1vщUb��s�9�b��A�������{<�����=�9��z$�U#�r�V@��Nڙ;^�La�6EM(h��'rL^N�ǧ��b�� �嬲��ꡌ��T������^cޗ}]�s:�G�뢗b���&�Nދz�\[C����i�;T{�k��&�3v��j���z�iѪ~]��P���ک�5^ˏk��}�ґ�u>��1���	R�9�)���g�T�x�y�↯ �ܭ��*��.��9�(/^9��.��i,}{\��<w�K�*���ޞ?{�������M����Y�ܧ�� �=S}�r�4��Dzq�������;~���-eʳu�Or^�zֈ��k3RWu����V�c3S��M�E&�2�M��_�S��W6���RJl��5T"��N��;]�d��;5Xd5����a�J5��;�8�S�YWo��E���9�A�����Ϊo�o:��p�w�pVئ���9��y��Z}�M{�Qk&s2�c�a�j�;���t�d���3�o�j�>�2�-����Wz>����-�Ve1�ƫ<x��L����Z
TΛ�h~�����s�9��5^i�JR�hnȡ���1>��h��Q^��m���ݣz��ӵ-̖�[��F�{=��eO���/CI(��V��ݛ�v��9����/�Z�л�V���k*��u�k-��QQt`e�^ơ�w8�}�ț,�s�y�Bɵo�}ꎸx�Z�K�s�Cx�"���~�<�Ǟ�"�W�/d%P�"�v]�U��A�6��	�?E��j�����􊺻Ʋ���+hJ��1�Y��od|���aW�:�"rU�rp�����4׶ײS��mJ �e.ǥ�y�^���.K�A��^��<c�����/a	�i��N����;�l�oɄ�zA��I��)���V�;���1秭Xޗ��J�����F��P�T��4�t�����`��.�׊]��o�ܫ�F���yͽ��*ȫ���Eg
L�)�.3!���x{a�4��n[���ѥ�/)KW3��
�̥I5ښ��@�/����ٟ�-�X�\��е�y����n�Q��t�Dk��z�Z�S�3������a*�l�7S㩶�0�ь0cL�ՏL�pT(��ړ3�+=z�٬Z�&�fm��4a]�.�M��o��#z�aS�c}�M��{,��z��h��Իj����;�������⎼�T��w�;TS��+�毥���v�ȡ͢���;��Cy��p���WZ�����L�=���9Fk�Ć��;k��߶����m����<>O��ˌ|5�Giv����E���{��H�o��^v�غ�Kھ^�b.�2�����s.����*��mm�j��[pT�#(�6+���������o�ѡ�Q+i�x�^}��ٟ?7�>���uy�"4���xk78�<-�\N�6�_^���a;���P��O+���-�@YxD�]��-�,֓y%�jӐ̋-�-{r�T�T�g�J��M�>�l��`
�ņ�\�l��]��f�f!�)���q\�y���&��wo�alU�-���j1���i�ٳs"O�y�x�0�Si�n����r��f���u�&�}��u^oɾSs�8(V ��]JVc
nL�h�m_I���L���o{��7���iшj�?e��fUE������حe�6���5|_�{)U-�t��U�<|�&6��جz�-�{��V���J�O*tv�x�뿗��p����׼�,L�҇�y0�K���w�.c��}��aJ��?��$�,�%�wϔ�)�lj�غ��*�jT֧���OZ�(Ҕ6�v_I�TK��R�8�\4MM�',�|���%�O-�ޱ�����O�����CC��)�%Ke��Q��t��o������G���ꃪ}Mz�;F%z��FԱ�"��V�M��F�N_,��蒭�{Բq5�;������ƿ<���[���7��g��}����os��O�C}����%s�g����R��,׈Q��"��^m73ӆd�O*���*�ٮ��ʹn�>���B�ձ�]Z�Ã�b~�4{���y��m>ܞ�gw����#��	�DdJ�eGH&���u}��<�M$�\��ye#�[��O&iY�M^��:|��#%n��8K<%��Ṛ��b��:c}t;������S=��z��f�"9��][�~��i׽��ץhYRY�$2��j�%˾{�<�Ԥ�^�'�(�f������3y�S��Um����<kI��;ڲM�7)�Ѫ�X7��x�{2Q�ӽ��h��wp�j�\��$ϩ�4vx?�tӾ�q�S�x���*������g,��j�_��T=�5l��&V<
y��@������]��_B:�i���e������MF�'���m��N�ܫ���އ2�G{ګ���e@�{ӄ������
��j��-����j-u$c��s �qX�H����o��n�tL�a�fF�%^�|����&�S[h�;^�J�Z��;�]�G���孑�=U3$�j��������M�2�g�3C.�3@&wSM+kY�
5��1M���U����U#�.���w��Чɺ�/.X�e^�!^զ����Lk,�wYfvZ�\5��J�Jh�R�}ڪu�K��)f�F;��b�8�=���kh���Z��9X<���1�Q�*2�����yέk�����P�9��.�I[��nk�x�ug8���B۬��ޤ#��}(���ո�q���Nz%�:t�l��J�;<UcgjNM��7)��31re6:���TD��}�p}�u��>ɗ���ϑpW逕�Y@��{��{�k�;*w4*ڶ�ק��M���]�v��h�m�!��}�ɯ���u��n��'qI�L��+Zj�bu;����Ax��ܭ�3m��P�I�t�3���y(��4�ȭd���=Zט������@�%n�s�*C��=��?U{�k�yq�B���N,v|������u�N�,d�&v�"�,���>BI���3��j���L�}=)�v�>����z�/�G*�g���ۘd��B9?z�l�g�gS���8��w5���w��5�]��� ��9��C*��}<{���KW����1'!�_:��ջtQ+k6�Te�jJmW�{~�w͵��ژ�f�I��oJB�?t?/�]��;g}�g����3�f�A�;ʜ���^�X�]^�^���-Gn���K�ZO��4z.9�'�+_��O̭���Ț��7=�/?m�j��;�B'�M��E{�&�-������[���w=�n!��;�q�Z�;�2/dW�ڠ���9o `ɝ�n\�u�f���+B�2�w Up�+�ڼٷ}AW��ܭ'b��|�q�f�Ր��	 �}��˖�ǤE�;�U|�ff��N��EΫ�-�Xm#r����z�N��ӽ�>�����K���2�v�R�r���ת.��F�������:���wK��Qٝ~Y�gXZ�!cl��m�W�V���DݲXJI��:���^�@g��◞�za�WI3���@�ګ�R'^��K��5wD�$�H�/�GUk��DQ�w���[)g��q�)�=KAzL}n�{�Cm�����:�������xf�u�\&�O{���S�b��^�}Puk^^�O��x�Z�0���A�F�)cϻ���L�^ʯ-~4��]K����'o��x��q�g]�$�.��[Q�{�3^Į���.���JSf���L��Q%V���[6����N+Kv�����c���!�Z�v��۩����9]�y�/��s&o��s�O�*ztj����S�t����+�ȩ$�i�=����̫zr���$[������w����oA%Jǯ���e��z	�Ȯ�����fQn�;ï�N�r�h�k�@�����og5c��9P���)�@���/��<4��l�^���6�L�,]5�^,[�iv:�����e5�x�rV�B0�d�Ͼϳ�>������/ji��#���v��ފN�q;IO���eI��y�u�����ƙ�[7�W}�=�vC[D�=�N�S��(��v����fx�[���4�t�>Ջ��\�\���Lv��mt��m7���50����S��d���'fvv{ވQ���Il�"QW�'r�����(ؼ�Smsr^V����RmU&��*{��vk}��o�x;�uk�?R��ɻ��
�U�f�N-��S�y��1��5K�[<����{U/Al�D^`EDP��{9���n�l&lq�h;�lP�閈ioq���=��Y�=]�q'�K1���L��f�˳R�^�?�ƿ��񩂏iJ4�X��q��]bWP�+k�8y�s.�w�b�U�W\Z�_լmҏa�H��*��k8x?�"ߧt7�ɤz������.-��������Wy���*gT��λ�w�Ĉ���2�˫X�<y`�L����]�fÎ���sh�Ƭ���b43y���Gi�Jr�BqI��$&7ol�(�Y�tMh݇�yP�!d�lu�g��ޏs�Xh�ef��a찃��M��ݚ~�F���:��,B�R&�{u����j޼=y|cx)��$8@l%Gu<�{\�Þ�Kd-ۑ��Wd����p���/қy�Ļd���8��V2�0�W|�Z�+�P���m-;��gq���oj�v�x'�uگ-�]�asx���Ê�	$�z��@KEz��,,��f�=o3��� �'a<��T��A&t�G.�ͯ*�5s&"uo��ť\{�$� >���=�2��f�x-f�*�{e1ʳ��}Hդ@y��xQf���n؁��٠.���`�������b[DծD����""j�X�ŷR%A:����Y�[�Q%��u���ݫ��k���6�+�U7�C��}��7LЮ�`�)�J�V6C�vt,��/Nr�w?��`��=�d�Ww�&?[4w��ɜM]�|�gU�bj�n��ͮ	��s'Z�\���z�dzڡ�G!�έ_DПq��೯h�d����(�pwx }Α�Y3/�W9б!����Q�/�d���L�%�0D�2)�e'Z�s+��w
H���[7�U6�6����`#q�<c{X�"�!sB���s+w���/�0���A5OS�9{���k�=���%�$uf�n��^=xm
�g&V8�v��LMU/Od�
�FkV9�e�itB"Xx�6�e�yMI� X�y��%6���R94Z6�@Ey���Ӈ#x�պ�O���s��q�������#!��N���}�K dY0rO-C��~����Ot6a�A;��C���j6B����RѮ���������qq�-/�sYӣk�$.6�ĳ 4e4�'�����\�!��l���3G�﩮my���gx�=:�b�ovm�� u��V|��'J��t����ϲ����Z��K+"�V]�}W�9��i��=Ś׉����|���:����$D�ޖ�bj�s&<0��Ĳ�W�W�]��7f�sA��/��`��CS���Ng,�"'{ߑ��̅�	��a~l�*֞a��,*GF&�Tʼ=n��9��]m$��fe0��G�g1�=c����"�~����w��+Q�
jا\�{���:C�����6Ƚ�G)mLd�T�u9��(=k�X�sk������|�Q����[�UzU��u�͔���s�ݏr���=i�����g�b����������8t�,U�k�jJݗ}�M���t ��a<��-�a��y�Y�\o{r�m�N_X*�2\��hΠu�3�/8Sssn����;�-7=�]�E�ݧ��ۼ0}��Uu����M.���v����i�tU֭�ؠ���Z� �Z����'����ܒvU[�vLEն��DU7c,m�j�Q=�Pc&(�h� **��Dkw��c�2CPL���g���U4wn�5���6��b)�豊6�AA$DWlΪ�u�Z��F"�
툊bj
.ͱF&*�"��=b�i���V�B�M�I�UAT�4]ې��PF�SѢ#�QCm�+��EQM��%�RTD��:�l��kZJh��*(��@Fκ*٦�Z�*��4��"��M8�V��MT�ŋ�����ֈ�*h���`���Vfъ�tP�gͣUvٿ��oۘ��ֿL�<FW��^ݽ8I�}2�&�4��ם�K�\�4!*�#��W+'#v*i�ڐC�>�]-�C(]��Mc2��33{�f�&$Y��T�W�P{iNL�-��K�����}�"��
uo%�
|�n)�sV�[��S������(m/ ��[~�u��^H��5�?;���t�g'��8����s~c��P�8mgyq���_���y+�=�\ɛK��M�7�qz_�5�r#HP�OJc�_�*/N�_o{;5�U�CӀ�^�M����;���f�^��?g�v~Ua�)O�Y�g��3����5-��X���>�ޜ�K�f��M�������EX�;<Ǻo�}�SzA<3�~%c�^~�������m�vw�}ƅ���^}KU�])��]Ov���-=Ds���*�g�K��Q�ӕ�}㽛�yyt�]��od��x|�d�Ṣ���V`2�L]eN]ڥ��_�|7�6Wp��-5�
����P���Ge�^�:+Y�<��{��ٱ�eL�%3!K��4�5i��M��T]�]A���T�b�}0����=�c����=�R�o:-�}��SqI�.�����#��m�}�U`M-S-уn��$��+��B�<��pԡ}�ˎ���X�3z�z���D��oa��m$u�(��4eK�e�DXu�飒:�.�'HEyW����T�������������������5�;dØ�y�U|r�_;Ni�b|}L"'B�@}�9�����~����Ю���<�{[�I��\�����_eA~��^�{����.��|�~��U�w{�њ��#�Iq�K�_;�����_���R�I�)��p�u��FcY�����_���4���8��O�-�9�w����U/I�͏}�B�����(�{W�]�g��_�ˋk����:��f-���Ż��X���6K�V5m���kP���d���]�$�d;s�X3\!�8�xȷ�(�rךB��&������m�q{U��#o�C�n�ѡhi�Ɵ�!���bW{mer��2=8���r�N�(4YH�X{�e�+kmm��[k������z��w�n�ҥ'�A�I���ڥ쵊�{��C�x������p���*��Ңgv��i�/Mv����W
�H������{K�os	��ݹ^���L��0�l�r�譙�B�G��m��#�e��+ �a��T��%LͺΧWc8G�$a����]���]3��õ�s�;��[[���*�r��K9*��n ���k�e�3cG$��ns33{�j)f��m[5[̣6/s/VR��*R��;n�6lm�||��Jj�a@V�3jqs�rNE��Ǽ4��K=��.~���Ư����U��y�f@f<���.O[�����p���=�yZ�й�?z_K�壄��C-V����T�����=�2�1E{}	��UL5=ݨ��a�Z^]"����������3��}���/�ׅO3X�g���=���*z�5�zv����'��1�K��f���Xn_�S�݄L���r��(�V�xY�Ie������/�r��b����Ÿb��}e��ZN�+rm�ݟ��̊kKj�e�;�L�IW�!F�����h���I-e��K`li,�(Dn���!L���J��5-٫X��PُZ�j�Rz0ڪJ���%Q���m���}��rژ��O�,[��^�}B�u?o�.^uS����#UX���=3���^�~Rݺ��S�V�M�R��9V��VSa�����wӷ%�+�3������N9�f���ǅ��y������t���FD����EV�'X1���}���y��2ӫj�ɣ�ب�6�s�q5����_�$�ulym'��r�v���O��z�y�q�Ʀ�-��W�Į�mgܸ���T��V��?%R�����7�sܮ���w����/�Hk�K�r�6/]/��!U�pi��z��R$���w�ǜ;����,�x��J���ߏ^M���sjN[���Dľ��M{��_��{ݴ�]��{�Gx��9��/)ޥ*�[kݽ8u9�68T�i3�h�M;�T�-��4��t���*�X�s��/6V��^9��Ϩ�]{��&��t}�h����E��B��f%��������1���qB���9�X��g�6z%]4��M����n�S���c56�2'\t�����P���2��S��(�Nqy>R�b�t�dVlM�.�F���#�V�f�M����fS��ܿ#�`��v��b��8���y�>�ƻx���jg!�,�4� [rv9]X���#R8�H��r�c�o����,��]�<�d���y���Q��`}u�+6 ��7��\q�ڣԦB�̬�5�M
�Y4���r�vf`��8d�H�)�z�׾����w_��J�5?{��o3j�9S�i&["9�|T�F˶8��Z�I���q�jR���P[��G3_ �~�v!~�ߑa��c>�N��_̈́'mL���sHR���t��E��d����)�ã�v�;�X��u]{�󱔺����_V\�6�ˊ�.�P�>�Fz���x{�ڑ��h�C�Ӎ񪗨�Vc׭��|��9Ɔ��b�ʕ�*����^({�U{��}�V�0v������3��n+n� ��EFZQMz�[S�1���lSF=J�ƥc2�jFC(�4��������-�nfz�]�R�9ߊ��:p��.5�}S���w��8�$���ô�4�}�O�ί;�A҇�c�i�qO�k��$$WGk��^�C�E���3��d�b]�V*���҈�����*=��%-@xm�jv��m������@��z��r�슙�TL�u;�/u׺�ǌ5���Ҩz*s1�#Qexc�5�q8�`
U�7J�#�ʴ ��	�����B˭5����川2�_��C�Su�⃸���39:�ij��Yu���/�:F��"��BԪ��]z�m���}�}���b���q]��VWynE+a�wZ��x�{%-V�Jrv���g��;�Wמ���5b£n�ٴ�X���hmH�5��B�3Y�WvT�$_��m�^W��3�&u	�O5��{ilB�͚ǕIG.4��^�|����S��z5-��ܞ�h�m�S,7&[b��Z�n��K�]6G�Qy�vFQ�X�ZN�'BxW�u?mxl�_c���3h��5|r�_?	^��e��Jn�;ymG�3���p5�T�쭡+�	{گ:�S�/��O�NՐ5Ͱ�բmcX|rr��B�ҽ�L64���	6��Y.��j�e����3�;$a������ks"�έ��f�5�PW��O��mW� g���~-b]LP(j�\�	���>O;���>�=���|�����񰑯e�qڣz[�e��g�b+4$צ.��W{g�o˩y�:�Oo��˥S�CiyӼ΋8O�*�]�ĭ��O���7�+�����kIb�9��v��A�L�S<���$icG�<��Q��n�Q��;�G�������)k�iR�{;i�;X;l�kk�����{��>�p�v����	�B�g=T�g��������T�q���m�4�W��N�;��}_}�w����9���<��䣟r׆ן˩v�[M�gO�oz{L�8��r��At��k��z���yu��b�u�N��c����+t ���tP�zH����Z������~��г?�U�	J|�>aL5mƻmo�e�=]l��^�[#������U����$\��������&�X�~�oT�����Ʃ�={��-^�1R�����F
(��F/j�'4����kj�~�J��mOI����xw;�oM�.��6�<Vl�Iz��?p���5g��<�)�5�	X�m��tL+�C�e�R^6�*�p���4)�+ig��5g�J��M�ZI��&e�.T�1���J��7)aW|<k܇��w��1I֓����(m�]!v�9�6w/vr�Y/L�+�M�ک�ﲕ	^���,�߉A�����EL)��T�f�@�t0R�zZg	����}V>�&u�k8�ͨ���}t�]�W$\���b�^��������_Y*إ�Oix���9����(4Y�I��Y���kX5g!���y��{�ѐ���꽘�~eT���}M�	KD�jT�Ʋ�b]X��<E�c��f�f)��z��SdF���I��w���^�I��ٽ�ҙ�H75�w]�<���}�����j�X��)罵7'[PP�� =P �t�`���;��P9RRb��S&r��G�X�>��Ԧ��:6i� �o"�m{���P�Q��m�e�ݶs�_�$�~]K��<�Q��b��I��==9E^�gH߲O>^��-�J�>Į�Yˎ^'��4\E���=T��v���k\ܩӆ�gyx��k����K�r�6R�нgx)F�t��:��Tl?#]V+�{�7.�uAԹ��}
��y>}3��Z��~�����)y�UxR���Y�i���e�������{۵��[�su;:8����g�ë���yƷ�g�����q��a����n���cW��1�<��U�S�A�����{޹�b�lm���Jht�x�63��ܚw�;[M]lhP�nc+Z�G&g��W�S��٭/sd����#9:�9�>3n�~����Z���������*pQ����i]LVc���������f��F�%�~�>�t������vJ^V���A;K��$�mOt����!|Sg��f�'��y��P�f������f��h6m2��oڬl���D?��fI{�.��[�M�d��l�glAly�����]�.���(�2�ّ5�ɝ���Õh+�w�զ5�l3,m�N���v�����tN`�j���P�<Z����>�#*r�����h;�&Ņ2��-8pe��Fbg}L���A+ϭ����jj���h�_y^�΃��P����D7PQ�[Yysp�n�{Zi��\�$ݷ.��>5T����X3���J�(�ب�|C/T��eL{�<ẁ����<��,/�8�y���j~�����v*ʎ/Q~^ڥ�L���{�j�+~�`�����늃����R���%�W��dz���K6l#���O5y�ܭ�U�J�h�������N�sxy٦OB�>=��Z
Y�t��	��\y�!ة��g�/�~"�h���]kł�Z�Q}/h�h�3�o����k%��U�0i��եG�����c3��b*P>Yo�6���G)��"��y���Lk�����Jݦ/"���H�s~o7��%�wt)Ҡ��w�E���oV�+
j�5f�9��-ۊ�<����Yc
Ngy�G9e����w��T+}�m�H���v�?nT�醫{��+۞9����i���Ω3z��ӝ��P�Ώ?*q�)�?,����wyYW�UZ���ݘ�u�S���~>��锷iVN���;�%Ȍ��b�[��>�A?Us|��O;Y��x��;���s���JZ����*��G/�Ɑ���p����=]�ž�<�������xf��i�n�-�Yų;�n�j�aS�,>r�G���Z���ϵ�н�~V�4-�R]�_Ki;����&�d����k�5�ȬZ�뒇�IC��g����{��7a��iw�g-w;��Y2T��.���򱊤�I��d���}�r�-Ž��Z��>��Y]�Y��k�z����zy41�Y%�j��ښ�5����/y:����9:n$���^�>���1-�u�}˦j��U=�Fԫ����6H��l$7~��e��⼾��V_bO*n��Y�V,�4���I�����+�'�18Wkq�Y�z}�Ӿ���p��΄���ӷ|.�{�e��ϊC+5������ӽF�bI����ꦐ/�<�xii?b��B�^{�\���_��mTr�6ѻ�й�`V-�1������������������ �|�W�+�LS��V��t�u��ʾ��m6傖d�FJp��`Yb��윫���/q��sq�=�f[���U�ᛃ�?x�կr��#I�O�V�!*�
i��=
2�tZ�	�e���*��� w�s��,�X��Y�yݞ��0v�����/+c��M��K��+vt��ܞ\k��!{[�݁Rh4�.W�뽴��7�r2GVyY>;3�ŝ~�{=ˎe�y%1m=|y��$�E,�XO�vk��h�Q���3�^���5�xW�q���y&Ox�qa�9�e�ǅ��$���FC�^��P3i(���f�V
���u]qW8k�v̸8�54G��Oo65H�{��i��G�`�o�D\���an��ٓ��Q���=�7��9&��6n��B
���	��K�tYC��W��/��⧝>K6gk0'xq��8a�t8-�NѱKw>��u윴�v�ՙ{4���xoS�;C�_pZ)�����3�J�@S�O�����}7���Ib��.������ ����@��KI�=��$����
`�dr�D�eɈ�Q��|:��+��8�%W���Sk#(�T��y�{3��]�PQ�#7
c����f\5�O:`��{�WrK�p_nl�[��=Y36���F��<��'|���"p��M8�U��3sG�1p��g՝/,�	�)iS+P������M�x�n=���tr���s�=�q��~��d��-ŭ�J(y\w�E��V}�tޮ����aL�i���ν�m��d�}h<��\�ʍc@�x����i����m�t��C�4h[*8��䜎�T�즴a5*״zY�+Z�^����˺��HrZ��%x�z�*�w�U36�u�J��ӜIK.!-0�@Wl׹�Cf��P��ڧ0ݮ<�X0Xq9�L-R�i;���s����{�>�y��o���MW���Ь��n�ے!j���Q�QMX@|����@���f�f�%�}�A�T��3��]z`��z���<�F��B��G����y�T�f��4���U-�(�%�­�ط;K��}#i�;!�ʼ}�>�Ҵmgov8���du*x��v{�N����L仱�Φ�#i��k���_��VJ��p�;-�Sp�&��1��>���6"�O��A[�k"G%��[���Iu3��C�=�,��7B�TI�z�z�.uEj�����X�qe�av�c^��r֢��R�Uݕ �����)|D�s_���y˩�<���#�1Wc4�T�6آfў�"��Zw[�X)���6Ɩ*�"����U�Tlj:��U������'F�]tk5APh�
���ikZ�;�Vخ�n�DVź�-����$���PDUI;:��.�%�TU՝m��[j�b��17mힸ����j��ڪ������[�1[5���Dv�WgTUl���
(����h�,l�q�V7A�F"�g�Ttb�wnb���Ls[j��E[�Z�nMl�"����LRE1A�3T5OmEIES��k����Zݎ�8��&5��UE%DM�M:ŶհSUk�5;ijh�&�����%����jfb(�j&"��,m�� U
*�PV�o�^Z]Lq���ٛ��1NjE�(9��#6��&�2@�˞�oݶ��\h�傟Vl�饢鬢ș��}�W��2�<����?�D���-�R�i�u�Iu���7Ȅ�K����Ǟ5�C�O�2E;`��v���kW�PZ��f�Q��+n�~S�}k�2���M��ّ�#혊�2�v�Zc��a���*+Y�U��}�{��R}}#��s���寍%�~^��ԣ�^�VWw�~(vvb��L�T�-5ڙ�9�������tӴ���4�խ[aM5�f�8�TV�7l����-/�w(
�w�n!<M���J���Ϲq�k�������,z.�^2������D�������܇�go)�g�Ү�i�;�o�W��<-�e�Koܯ8�1�����n>�;���{L����W-��Kn��()�Ǚ��#�a^ڢ'G�๾��g�^�	�ߠ7�j�f��ԳY�I��dh(b2��%^kZ�dſvC[TOx�{���\�Ƽ�x������%��w\�ou����o���ct��L�kj���l�39ȭ5h���"pa*���1�<A�y�^���io��Thԣ�B�M��{��ұ���BgJ=��`��+Z�X�Yx�R���^��J�K��'��ao�<xz�
r�ŁE�ʀM�諭�+j'�Ȭj��ԅNg��-��I�=�y��,k��U��xE��V2�[QR�O��ݼ%V"�)YmE�nj����U^���8|!��W���f�)���3AG�&�eTcJ-X�rlVhM3L�;���ˮtI�>T�D�z3�=�;�T縛k�ĩ��LY��k���N���X�7u��NS-g��v�3a�M�릵O�q��>��x��[�g�Y���@[������̜I��(�K��.�M�ٸ=��L2:�ڞ�	��O52��X%�qm��z���>vQ�o˽au�������#��=Jqͭ#|�l����&���#��a�C�-�c�_�X��R���L�~h�y�W�ߡ���$,��ݪd��5`�d���񙬝�.ʢ�/�]�o�O6�2���}i�<�/rǌתM���>3�my�{�%q�bWm����;�*u���P���7���_�e�/�{'Zh_,�Vj,��#�����n�R�޹����&iї�м�~卩x)j�hg�xq�AR���=�2�Åb�qz;�|�I|���V����u7��+�k���P�=;���QM��ŕ�F�tgf���/6�UY;p�h^�7��I�4���^E��OM��a�R�O����sm���Hj��<�Ŋy�e��^�p�h�u����9����ۓӣU��߇�F���KɐJ�t#���#19۷���5�U�Ɨ���;�Z�v/rb�eΥh���uFk��)��?z������_���r�ɓi�߉���w��®��}���U��.�6����)ٖ�R2���P݆���,���n�=��L�xe���9�ۘ��y��cw�׋Ϫ��)�}E>�Qe�KfӬ+��P�l��R�W�Oc�Qp��u]چ4��q��M��TvN�V �=E��4r�#��$#��|��:��vD�<��E5���W��1�	�|��ŧg���;S[Z�c34�N�m1�f�mJ��8�TlM�1�(sP�$25���`��܀��S�`�ft� ����K����*���ZG���}i�i;W��,��0�V7/s��y�3n��%2�)�/���S��CA/-o;�ɢ�*�oƖ�Tp��!�;���c*�ۈi������|%�tҢz{��M�|�^OQ�Z���V�t�̌��gdD^�̼�u�wﾯ��:=��Y,ۆ�5�K#L���1�M�s�{�2���=j�z�jHN4]�1��B��@ip��d��S|�Kǝw��y�D��\Z<�����8���MJ=;��o���jc4��n�L��5�M��*SF<�;U�VѪ�e�������Z�^���w����.ߟ�b}Y���ک�����^A�w+ma�zU]��>Y{{�ՙQn�D���Qok!�6lzʨ�ųg����})��N�]��o��N#������<i|{�6���i����ܟkg�t$�.���L��y�}W���Ͱ�� 6�O�*��R�B��<{�Me�c˻#��s��5��W�����_Wxy�=]���*�ҟ�o�����s�R�qAw��_ooHk�ח��g{7�4w�޹^��LN�t�3V��vV�=ٯ����9�k�Ǽ7��M-���{��[,�S�Lkǵ:}��۲�R%b�����.׼��2�߃���zse��um,´�˝��:�N�H��5�9A��9�Û����Ɋ^���xV�5�������^�өx7�A6�=�I��KǜN�nP��1�v�./ym�����g\W�wT��!sTf3�w�r�v_w�y��dþRZ�ql�8g�]Lȕ��Z���a�-�V2u��0�Ț�pl-c�4Q�ט�$��}kR���3ȷR�YdE��b��!��7;�L�n�%�o10�luY-+UҋQ���l�8��3{�K�/�����6mIB�ni��4׳�e�q)��e��q�UY��Qar�u}j��`�[�L��y�\���������w�R��3��bש�ᣟ��>{Ҝ~�������"6��(�ڋT��{2�vI��ޘ��Y�En��������ȼ~G�s��3�ߠ>���{~^(o��Ui��}�=Ys���-������W[�Xc���K���}Ju��տwy��m����4+.4Zg����T��]�w"��=Z�k�����u.w��@|�{~�Zݗ<��s^�Vs^?Ni��&��_t���%�_D�u���[\���%�ԩځ��f�u�kߋW}\"���eCtv���b y��o�����P�$���2��6ȫNY�Ӹ���۵
�£�o��[�%E�o�8��ej�ؗK��ۮ�#����8����s��W����G��JZ�
C1]���ʵ3�����b�Z�*���~��#h����5γ��<��P���d8�k����'��]��z��녱{�r��uG��S����P}ӭ�.�Ϻ��ǀu�S��MG�^�{�G�<�G�k�F}�߷�@�P9Y4��՞�����)w���b�q��{�~=�i&��J<�s�~��<�;`J��Z�b/"��Gb�-��׷.���fZ6�+R����p侑M�=w��S~��8�����__%[E�nZ���J����I_x
�Ϧa�}K�m3t�=��z��Z횛UI��t[ܴ[�=����z��<]xv��f/$�{L}�.�k�)�lQ�t����e;e���k���V�g{K���o�����)M��jb�%�d"Z��	;q���<^^Zx�k�YYޠ1�<��\1r����#a��'f�LT6���1ª�2��5E
�z v�[&�ڑ��r�<�u�&�-�g-SZN�͠�#����;��¬ �qt��h*(����#����l�b��d�]�����8�6����e��v(�k�p�W���:�#vw�� ��ݧ���7W��着���D���3�]�W�{���=ū�ֱkt�1�Y(ƈZ��N�S�n�b�M{����<Y���������k�����Ԗ-]K�T���/7���.]�gr5*�d�i�-^ډ2���H��^�<����8�cy���pGW����}I�g��)�{��4��L�|���\5�+o!><Tn�qY�@��j�a״ڝlT8�?nT��s��k��~bC^u�[�[���ߚ��y6w<���U�C�DN�#ئ��^����|I�Q���ٞ�SOޫ��P��؟^?W-�++Ǖm;H��{ݵO�]�_���uhݬny�YT^R�R�d�W���������h�����Q�i��z���!'z���3/n��,�YLֲ�J�1�F׃f����,�y̚��;\wd��xf���(3v�S1۸lV26�vS���5���3k��*�9��z��{ڔ����/����L����(�n �4E�,JJ��ge�����u�t�=�񽋠i��?����iz����t�J��	V2����:k�s7�U��h�u�FR�v��G�6��w���r��ϋ�|{�tm4���U�<u;ֽ٧���	�U^��m�-�
��f�MS:4�{3�ҥ޻]uㄓ8LS���5�[�>XO�<����~�E}�S=S�k{Iz�y*��;Fkb��vպ��M$����v��}�י=S�x�X~��	��5���K��mM�Y�T��2�f%�r�k~4�K��ނ�ކ�i��V����ۺ�UZ�A[L5�V�e�;ɻn|�|��������%��͸�g����;m��6C�ڂ�j}1��eo	Aۓ~��:��a�i��'��꙽��ol��t��R�����4a��["���ʞ,�fXӶ�8�Ay �sԌ�f�jQ�MN׬[6��W��ܬ6Sb�~ȓ��~���&ߦ�Ϲk͢�T�Lym?T��gyp�����u�3�Y@�I�
�|��k�HݖתT�n��5�=�����y�������Ze#,id����F���i��B�q�Eٗ���E�D����ܔ"��*c�1J����u�t�)��2�N܆7;݉�K�%sggu!w��e冠��7��e�f�<�f@�ྩ��TX���vE�`�
��YnuA9;����]�ޒ�{�l�̏�Uwj�W����=�ty�S�)N!g�f��gE���N~o�V�����Gjy���g��_�W�g"�g�#��.i7����-����NYL��u����.U���X�;�Cwei�y�cEhe+��u3��KLZ7;�Ugs̮ݛ���l�5�t�1��(��Dlz�5��Vw��{%.W�8�Vz,4�٭���ڿ+{:�����#)4M]���e�� �Yl���fz���O��I������cܖ��B��k|�$;�mPy)�]6n
�E���dvy��o	噧��vײ_fU�<fG���&݌t�gf�)�c,�%�j����"�����g&��mO>:�=^UV�S���^[�(�m�2��\�§�T&x��>�a��'WS���������R��
��gi��*��j!�Q$�vT9���ul3 �/�S��[��9��k �ý,>��q������1I�>J��}�Q�Ss3�`�;*�����k��^�3��'9Ӱ�N��Ou�$/+V�x�Ϋ����]c��3WZ\�q�%I����:(���,���;E,��D
��wy��mǇ�{��X��|�X��ū�������G����U.�b���.��aW&��?[��[�Ǫ{����yo��ז�"
�]K���T�=����'G���:�ճ�n�zS6��}�(j�=�ܭ���ʆ��s�����R�c�5GБ�g�u��h���6A���^ⶔ��~F����a\�q�ٞwZ-�W9���T��v�3���%��.��^[���o)G�X����k�v�unE��؟���p^߈����v��>}������w˼�K#��~l��_9l�>�'�>�i3�Gt/}ϤƽYr�l(JV�I�vt]2I*�R�:�#�_]>��W3Y1m<�G{��饞�ř[kd��d�[�:���}s�U�ud���]���(�+��e<�O�z��S;Q9��eg7�a>~�݇��߼��<��㝓�^�Nk(��"l�K*����!�OT���տV2�n�[�3�X�+���M�.P�YL<� ��I��)EUflJhޤ\�CR�n������J�L=%����bu���w7*GX��Ǹmg\�V�I��0�B����b�*b����i�m;8�1^Uۤ��A
.vV����;WO;T����*���燪�3�7 �����9fX�E��f�e ��M�m�N;������]��Eh{#t/��,�����"��*��{�^C�j+YwI�"� k�V�5:$�C���;��h��c�#vs���Hf�����ie�B���3sk��؃-]�`s*t���|�`����}ȗ�b�b�4�:�;�����)#����ulǯgQg[ǜ�O��P�(w��W/9�{s�� �~Vx�.�!`AW
�}�W�_7�`�1����Ų���������N >Ka��[z�
��5���ٮ�g6�bn���e�ؖ:*y��c;"fKB܏p ��q��Ά>���p���Q�W�/�I!��lw�gR ��;��K��|�Rc3���:��[�#8���,���1�A"$|Kx�Wu�{��[�y�d��)��d������:a"�5�g��!S�r=眞>�ttloR���n��q����Z��	�c��O(���7�Q�������N��V ���^�-]vVP�؏d\a�Ļ��XE6�́W0�<;B���p=�ټ+i�0�!���J��j�EiB����z��xл���/���,��}c�K44�M�pX��pC���+0��v��״i �?"}t���j��ڝ���rYdB�^(��o� ����#{
­<�4�{}F�*/ulS��3p��G9<���(��lu3F��)�:���Yؐ�Z�B[�B}4v8uG[{�f��&��z�7��Z해�3����J��Av*9�/S�+u^5�)��B +x�jndFh�^��sH�իUx�Γ{���� ,os�V�#�=��pE:)�7������g�ku��u��sܵl`��|�Սգ���Qm�
���SAT���=&�q���l�,�a*n�6=�V�1�{��t�K��u�P�t��#E���1VA�l^b�����֢@�Y�W�6j��y���rl�:�+�g.͊�xR1My��m�iSㆷ$�x2yc�����ȫ���De��3�gB	����h
��k��ϣLk�Q�1!Hi�tVwG��;��f�p��*;���횒�-��
�NS�8����C̓!�Jhq��8&CW�_m�O �d�۔vmkIU�ufSU��?������\a=$����K�T�GN�^��ٮ!b�W�a�����X���kS��Q��=_fޮf��^ֹ���6���8->�ƪ'W8��h-����u�V
@v���ltYf�6���7e�wo�W=+����@�����=۴�M��T�4�EAQݵWc���n�h��e��T�V�TT�QEGcZpEte��X�"����DUMtb��j��h��ݷTl��h�*�h((�������*�.�)���ݲSb�#m��&�]�
��f
�1QQ=�m���m�5��TTE!A]��CD�;nٶ1ATQkD5a�j���"J	�����6�ETU:%Q66����D�6�(�*�(�����h���&(��4n�Pu� �RP�CQWF���;j4i(�������(J��cd�Q�L�DHDMAA]�Iт

����V�i((h���i�����|�~|���{��Ͼ�����)�s��藪�7����(�/���Ԟh�.� ��(�l�o��+��1j&�僽��类PP��F�F~nj�cO��5��M���<j����
�[�A�*t:��[ް�Fz��'gi9�r^�9S��U~���]�J�O*tv���:'�����X匒�*5��|}��%D9	�G������}'�7�b%�=s�D��lmm�,�ݗ�S�J	}�f9U�T��m�Z�"7 Tʹ�xH�?	�OK�rZ��zv������fJ�.�Ym�j�ƪ����+X��Y�o���A�����%�9��UG��v�5��,4hz���?"��@�����-c�`��\��������"�!53m,�~(m/ }��u첡�Z��� T�>�퀕v�<�׮�>#2{�Jk����g����S�o�j��%q��%s؆aθb�Lm�N�y���#�D)�z������t�+<���S��z�ּV�m_��<=�Mi��u$�5�nx����w�)��N�V�xzv�/'��VzB�b@�:�}8N������7���o��v�n*Sw@��^;�Ə1��`��lh[��ܸ�:!4t�-ޗ��Ksh>�I�1v����#���=�ژ���ث�5%S6�>j�I�5��`Q���)5����������4��Vi|�HfEh}�|m�SUg�*߉��������֘_+O��e�o;��0�ϝ��GC��w��b��aJ~
����5��KX�r]���<�w��w��U���BW3���n閚��{�D���K��-�C��ت����;�:�U>GJ�Ie�v��B��C�~;�N��H�^�Mk�]����T�����z�|��9�Xrz�ߊ�z�/�A��-9t�ω�	��F��?_�ǹ��;}\��wm:�)��]E�^j�ۍYLb�,��ă��{	�d��9y����|i��ڍ�:�`�O����kt���}�Dǟdx���fQv�a��c*�y`�M0K��V�a��w+��/m��-_�8{��7�&�:K��(�.w�Eot��ǺRŰ�g�EF���a�Q6�̜eAV�E� ��b���)��<c}�~�-�K�g���P�5��%;��F��s��׵�e^�6b��[�A��ʢ��řD�@�y��Mnv:K�d(��۱j�F��;0W+A�.�s��^�;��tDهV'5Xs�S=�$n�;��̼W�}��nw�}USĝy����V���8��sԦug�Қ^�:��yd?��9p�blB7@f5�)�/ds�8��#7iz����>�S��{���;�e'�i�.[i�w��� ��m�'�*?���$ҭl�
w֘���[�"�r��>����H�ܠ+�W�^J�f�n�uCL�F������H+�¬��!}{Z��]���������b5�C���Y�7�:ȫ+ǍmQ3��
n�e9J��l�9�J1E�?�y�S��l�u2����ʹ\�$���Xn����t����<�5��6��M��c72�VZ�7��a���7tʊ�r�������J����ϳ�oݐ��OA�}�K}���9��M�����N��Fm��q�D���ڵc��w��w��)���LM-{��e�s!���#'����j���gu�z�/����W�P�]R�S�r98�zݟQʋ�.=��b���5F�Ī1���!Җ��.]�CAP��r�p�%��ֳ��|{���)� o�-v�:o�e�$�XG���ʦٳa����B%G������®���{��ֱ�1��O&@L��D����Ds��E�ۓ@��4��Q����3�>"�n���H��>Ͼ|�,uο���O�J���b� *n����D�bZx���h�#"�M��-I�-5��Z[��C`��1w��s�t�Z��S�a�o=�?0R�j x��s�!����;�XV�g��;�n��k;��Mț��My�������-������㡡�8�y�x��nXRK������t���.��j�����*�;e���a�6s�/n�٘�;���k~��̺ _Oq#:ƃcg�.jk���NV�����`��]���Vj��[���,͕� 5��&�z�'r~;���-���w|�c���cok[���	Pw�X���O��o�r����ߚ����S��R��m^WB�̡n��]�mn1��"��j<�.�_T>T�]����GH
�p�|ힴ���t4���WF��M�4�󸶄�i�e�egd��eod�y��Ι"�£#���暞�a0M�������s�aU��d�#��m����9G�VKj�:[5[Di�2�u�;uu5�5��SF���X�T`I7��N�oc�H�'�]���'C�?T��u��n�[�k�8��Ձm�rQƀiu��?Z�`�F���.�Ma�x�U~�����+\v���n�ʧ����4��j�*]<�L^=�gww��&�ԏM�N���8�kؚE4ϳ֙�&��B[�l4wd����Jz.&i����}��o�dÐ�����>fmȪ���x��;��t>�^gR����@���e����%�)h�;��s4Bݦ�X��j.hD`��ڵ5=X���3"�S0!s�s����4k��l�T�j�qyjvK^}YP�[z7I��ȱ�suΗ�L.`knk+�TbOg��*P��SYp3�v}G)���B�@�:Z�ay
0u�����w����n�2�>F#,���N�DqQ�5SY;�%�a���b���L����b��0<^zr[��km���7�S�v"����������]�<q�ڟ�S�t�(�9�`:�<��;��u�}*��}U/Kr��ܮb���0�:x�	�m�L�?@�zP���,��/,&-����{Soٗ����>D�,�fx�[��b��Y�=���f��6�1������2׳����T�x��
0��@?7v����9xF�n�z�9�5�d��.;�k6��4���홈�a��&���m��uDX�G"F�;������ᆮ(*4���+�se��47E�:��+M�4@���tg��W\Жθ.r�7@}=<.��K5=����Є��f��{����Z��N�:�ݿÖ�s�}Θٷ�{���Y'�m��svftN�<S%˥��R.�f�Řxts9�o9s���'GÇ��\�sz7�(��6e��:V����r�M��X\儙���R���1��i� ��o~f�4���8ӫg����@|��zy�_�!g=6uC��|--��'t�9�7��d��-�΃�.V��F�쎈:6���p-Kd8뜄 v�1��Tv[�C%�.NWA��� 3��{��r�	asy��b�o�I���a^���w�g���l�^s���Fy�~���J)����xG�����nI���#^|�8��@_�,��f����S��Xb����૫�R��	���A�Nv���ٱKr�_A�< =l��ԪX]=jy�Eq�6K��fR���W=����wys�öV�6vS�9p�gb"�׹�ص�.���%Z��df�ROF�)̸nw�R�B��e^<��ϘZ+n;n9��:�k�	��H��^GL�a���S��ӽ<����Ꞻ:9�(�����f�0)o;���u�̭��R�-�G<��Ǒ��b��l�����Tn�n�����Q�4(�����F>aB[c#��#ڧ�S�t�1��{Ng{z�����m����^�b�ߘn������=z,;<ʩ�4J�wL���7�(�~_�u� �`(k��~Y����t"��|�cd�;��ټ��((c�F*�s��י�%�kzK��<�$��w+�)�n�M�Cϴd��u��)=�塃/�c�P!/Ӹ�k,cp��n���}��~�2��n8o�'���\xeվ�!6�c����֡��N���w���^a#3��v��=�^u�+�\�
�� �������9mtUT����g�����v[V�M�S-pբ�����R�;N�� .df �/�^�:%��1踱�j��]Ը�����뎈����Etj�O;V�9��8uy�������|���=���T|�Mt�t_k]odt�����@c�7�*,����x�!�����-���ш�Q��͛��bJe]�x�(U�ř�����@^�"gTpې����P�3�qC::_Lp�n�,����j�l��C�7���&�g%���Zp/�� ���!���r=��-�`�k:�@n�R�zy�;2P��s��4Yׯt�
�)�h��j;��.s�	����tc�2�=�+fmdv�~�(�|uZ�����NBH�
���ٖ~�{N�N����v�[��'9��d���fY#m��7%qOӲ�����̀#N���O>�����m���,=*��*��_�Mf�~��`r��BDz���Z�a�:��Tͦ��K�t�S��� ���g:�]�M�pV�4n"�����;sM�,_̱���w6
}n�O6j���1�γ��J�����zkr$/6ײ�����^��fmM1�$�W�֏�zZm9������kg@_\|��)w����=m�`����7� ��S�kq�|ou�wˌ�x��yL8�T��}ʑ���U��n�Q}T��?#�`r9�cD�n��vٳ�FOGKp�x���x#aYl	���n��9��'Ïl��X�l��Z�֗�~gՓ�	~|�-��r��"�{B��'.Zb8R�����F�^M��m�k.9<�[��ߋ������׸��\a�2K�r8��a��SPZ@yi��o^pc�m8����,JwNDt)t	Ɗ�2:�lU3�j�x�F�;��W}�w�r�4w��Nq�2�: �]r��Ds�;B�-�w�	��}�F�f�ܕ����n{��bV"��6�?F�I��-��øK����{I.�rцYKap���T�=����g�MY�����я�.J�㡗����;���9Q0�	�}�euӲ/�ӡ	�3��mט�U��k�Xg؟{t8[l�p�m��DK'�z<� .6�[���u*���b2����n�D7wK��ϐ�FZ�.Y\�Ѡ��۠m����\F=�k���.�d���NN�zsݷ7�;�g�l��q.�3~T���Ǫ��jU�5��6�-��KM���~��s�a?��c�g_<D��w��X������U�}��P�o�8츋���hxX�a%AuE�{�5 ��M�"�
w#72��B�;��|&e���� �a�7v��G>l��m�^��Wl�nWfn��/_�	�+��N���Y�¬!5��M6�=O�}�'�.2�إ���o;���i�˲�:���4N�M�q`�~����)y�B�ū�׿���X�mjw�=��y��F�t!F�>}��l�Y���cD#
��#�ɐڨ�޵��:0�n��:�ڝ�����HH�'�m��M�J��Y�F���z��iu�H�Y�[��y�wA�~r�W��-l!���	�S�3N�-4͒���-��nD^u f���WY��,'��ᦜ�Z�\$�J[�F���T�w�vK^Z�.Yd�hab��x�;�L�Mb�`�s�m���~�4��T��
S5�#>�g�r�: \�B�@�:{'7�
���Y��\Q���q�e��'J�x�n��S�:3����[��YW2�֣[����A�����/5�'�!Ɣu�����ӱ0�6���'�Xݲ��<s�'`:F�̈������~��a�=�`�uPꮹ�3���AШm~'�y��4�q����w�\���~gaA3��]�lܽN�G�����t�8F-���mu�ٜ;2�[�Z�M�ą�f� ������p��9 ��w0.m�,X�Z�kX%�����r�WWB��d�'�2i���ޗ1�򙮡d��o�+xj��o��(�ռ0ޒ8)g�/�DɁ����C�0	��=wh��`�dy�3B��z�{��N���L9��%ݳ�ߧ�T���k*�D�!b��mƠǭt � z9����e���J8i���=�K���kή�]�9������e�fa���.��癹��[�6�@��Q:���f?'U�����w6[�[͔8����� ��d��)㕤�W�Ôd6N�������}}�8"��D.W.�0�ۡr�<.��+�-����@ǉ�&���B��8�y��lt�����a-�9�:�����!G���U~�>�~Վx�O���\�R��+���t�Wo�m+��:�����x={Tv��y��'=4u�f]`�h�ǻ�i��݋`�u�n��4z���{�\@�nB���D6��Zu�\{k���4��m"����:����l��	�=;O��+UM�$��+͎�)�)?5���P��c�dҼa���2�ӪH�=w����\��w�D�@+y�}���	jz���\%��L����v�ɭ���)�;�'(�Y�;���?a�u]<(�ã��Re�� ��6`^:�>������s��p�ᱍӉHs՘�gF�,R)�Hk\WL5k^���v=��C�\.ު���T��vy{m���dކ�W����K��P,#y�'O�r5��L�_��h�:�r
nq����Ym�G����;!��r�	 ���H����t�{�]X1��۹7j[3�ѻ�o;M3���n��/y��`���N��-�)\�|�ټ�N�̡)4�(�B�	�Ý4���CA.��NK�|�V��Ky�=�'@�Pܤݥ�Q��n�[a�&<1�^[��7G�6�*�፬�V`�+���9���'gw2�j]1[d������[`�x������HK����;�|s�K�ÚT<4qw�]J�G��Vq��ị2n�����w&wR|��p��)f9�n���s���$�/�8�P��c��c��foGڭ�M��׀�	��OJ���S^�Ŏ�f�j]�����܍�J�³��Q�Yټ���{�>����nzj�=���3��J���oJ�&%X3R�{�ٰ�x�a�5�x�^"�)0h�����*�[���=��A���� �����R+�H�TF��KÅ���\�e���ćcI.ܙ����I��u��Iŗ]ĖSm�p�����G�U<6����y����=i�-?]r��g�rʥW@��0P��In�!A�^$��)�Y%��31�#"JBlS��w�z�Ifh��C�	�k�����f!��C������˷����t��B�=���jSܜԂ�Ƅ}ٽ(\7�8��i�h����d�a���2�cÑ�/r�N���xc���p$�e��zuP��dP�}1��+h1ۧ�I�ᑻ�)!J�c/{���#9wF��I�=͉��oM�I�Ŋ��H��n��=rt3t`�f�E�b��+AxpR��;yY�]��r����U�7�ֹ�$Q.��šx�'(³�C���L��L�TK_���q�;��Ȕ��)�����T�ͷ��8��fzʷo84֕%�٘p��ܼ��,~Ԓ��Yx']�uz1 �_8sZ_r$6{G3	1���p����f�f��E&�0^I��:r��|M!�9v\�"�׎̛�|DWB���i��m�5읰w�4ɀ�y}�Q�d�V�J(�]AW��XWV�=x�:O�G�=����������oډ�����x��S�r�Hy��4L���Ǽ�J���Ǔo�6�1yi�K6����I{�M(ʋʡ:�p#k�7�7F�^qu�%ܐ�Ӫ���}��Y�)7����i�Qo�	���n�r�0����
�`ɚ��QrR����*Al'���fӐ��4�N�A}�ݞ݁io]N tY���d��8�}��O�1��0�гػt�P�/�Ѡ�F]���l=Ӧu�>����~�ILg�go�������s���=c8z����▾Ќ��2��.XCB�����{��Wt�1�ՔμY�rF����f0/��W�Ŏ���?j���Z0t7nH��x�����׋T�@UP(
��
(��1Q$A�QQD�)U�1;m��bm�C@A4QTD��,�T[& "h���������Ri""J���)(���	!���h(��ъ���F�(��

J�&$Ҙ�#F ��"��)��F�@�����Q�
Z(��ij�JB�b&��4��
i�A��B���D� +@�!Ѧ���������*J*����hB �(J
�(+l�AEPP�j��m!C��QABP�t�PPDDR��EACEU	PS�AhPED��S@Ut�MI$�U,BQQ-$MU5�5CCAATRWU����u�(�����K��mq��}�e�g�7�%��gn(Ү;@5k{�nj]�v�ީ��������-O!Flf�^�,4�͘e���L6.zJX�b�����g�=�#���[�/qP��ƀ�~��H�d`D���:V�t3uJ��,ˣ�YTĵuQ��ɥ�!K��	Y��է�ݟe4\��-ЪhW�:�wl�������#����S�!էaWk��;�r6��C�2�� 3��(;dU+���U��l��#m�O�n`�4��μ
?k� �+�!�WL,��/#x���ꪗs�Y�4J��a��7Ӆ��agRUv9�����M��i���G`�Q�T|���RM�~x�~�Y�%w�Ez�W�O*5��Uf��ݞCK�7�]�v\��Q9
p-���q?s?��Dd�\�.~_�p>���Sd�eF����6=��9π�5� �-�HN��Gyf]�#"��d4v�1�RM��Y,v9�N�Yy�h��~R��ⰡWOe�?y�@;mĢI�/�p����([�ō�/z6���b��(ڼ�����Y�f�ѹ��g�]��6L�p/��8q� v����)����;���S]R�a(I]�l��'z���J�s�%oh�c��N�/X��`h�	`�{t����8��z�U���w���vvS��=�:<ٖ�vwɑ�c�
$M>�9R�j�r�}��t�<��Kn��TNS�fT2S�������W �a��1�<�����؞�y��Vx�Jy���|ˢ�����'�����B��t��r�&��l���;�Ś���V͘c�*�V��N��C�h�.��3��N�]�	W�ŋj:l�%T�D�vzi���랈�ĥ��_���S�dCi�O�jS�3���̺O���QQ�=l̀FN�1j&6�zih��/c*��H�4P�V�ǐ��L�B[֔m��Y9��i�(���&壆=��x�=�pV�J��_B�Tm&����:Ge��G#:�4N'�9M��yt���5�(��M�<͵�F^OL��ldN'��tò�0,Kd*�%��֗�S�[,�s�P�9���X�i��)T��f���3Yf�mVq:�vlR}0�>��k�[�	c�~l���LM-{�v\u�s!�Z�:�u���%_c�����ތ<Ǟ��n�#���q��<�qBZݟQ��\q@���Z2ь�|~�a3�ۻUϧo]���A��s�t����] ��F�c8��Ap���[�=L)Π��f�k�OT�Y�O6��Xy���y���l?0��P6�GAY�Y�OC��t��ɜPd쾊���xs�ٮ�����Wy>Ɲ)~S�7Ov�ilC��o�T=��\�b�K����[����u{��2�5MqH��)S�:Niό�ִ��s�v[��
+)R{��;!�[<dJElL���h��*��c���:'#��k�(G��CE�����_�K.{� �3Q��e����ˎ���r�y��X��,����'�^�홎IDZ��<��`��1y��'j�@�{��D�u�p����td�Y����W.�m��8���@����κj�m���G�^vgm�r����Qne�^Dou��9n��e*z�)��==����cWi�<�D@z��;X������v��,�p�k:���_Y���������u��ᄚs!��E����z96�Vl���nn��>��\�t�}u��&���e�M���:�z���l���.��Egt�<f`U�'������{�>�u����,��V:�F�/����z»w�پ�ï����B�]���y����E}P����}FY���l�	lO"�!i�N�V�c������xT�������e9�}���]RI�s��Ӑx-lQ�UTat��Q�L+#9���w��t,s���M�pQU�.ynw@,zhׁs���M=.w�5;%����~>i?�k�K�h��ܜUv!:h9���p���xqd)�A������!)�����=X�ɐ�03�.�ɹ��j�3�W�
��c8<"N�}�.��c�MO8U�����K����k��8>����Q>��[�,g5.����ؕ�b�����3��-'F����L�����̿6���6����y�c� :�����#|��kC���S�����0y���SU�ǞM��N��M�2�=��ð�;�nx���ʢX�4X�W���""28T�}�c��T�"��f�
�f�:3#K;�k����;�8��k�O���N�5OM��ޕ�:��;>��rE�j���4���t*n9�H�7�{!������vME�S��F��Gnns<ܰ�g��,�֬�[��j��6��l�,k��6�3�LM�ڗ׉"["�������7=�̕t�yhP8쳗��kϷr����zʲ^�~��uIj�"�/Fh��|�y�;TC� R9��:���H��۔+�?�=��Uoqo+(_n��tm��+�aw�S�2�gH�����E��e�4')��Y���.z2xY�\�ѕ����3b�`�{^�Y�"���7nU0�~�v��:�K�ɾ�z--��fy�w��2D�׋���M����<�X��z����!�\� ���;
�oE��Ps9��i���\��_L��+{!E3���E���λ��˨����fes�Q�!�ǰ�6�v���;ϴ� ˹���;ޥ�/��6 �D��^ػ��Bo��V��X���η���I>B��/�fU���n�X��5��Ǐ����K%;�K�_�E~��w��~�l���af��N��Z��ՎBy�"ml��FG^P�S���s6�=�k�+}=m�v�:z��j��h��4��x�c�j.�QZƢJ�dlY��[=c������*P�>譛��p��_A�t��װ#�U0�S֧S2�Y<5?B��M��{ݭ�!�:�ع�1V٠��]��ן���K6�J;L��Px뀖4l��ݱkD�H���6���s]@s'�<i�;-O!Cf�ai��XVGOKuxm�AB�l:EUa��'��>LFо����W4)�s��hSQ���;�Y��a�����8�wUu4�����5-�n�v���3b$���v��^,x,����[��hSu���:��P���e�=��c�e��%C�舸�r�U�\��CJ�e�&~GZ���Ǧ��T�bM���׃���ï{�T<�=m7�⪹�w5F��Q�=3s� �� ��DL���x��w��w4�U�¢��l␠�t�e]e�ޝ<��G�0���2� t�P�r�&e�6��5~�����a��c���s�qD�Ժg��c�����g=�[6�����8�7�&��#{g�侲�Z��u���kz�)C8C7!�³%�PG6�"�&���F.�F\:+9���V��(F��)��%]���e.��e��RVU�HV�r�c��o�~�>�.��xtln�mw<����S<:����E���s��i�l�s�@��Lظ����9
B~}���h+9��۠+�-�}�0�QǞW<Yym��b���{WS����h�ڈ�����C^i��t�f|֟�>:��!��8	m�Ny���KM�C%�޶)��盺�Y���@�$��X��~0ד[�? +��[� [��y����E������_�r3V��ng��c�WWDX���H�fW9MM��L1���t�H*'�d��`�ۀ׻���H��Ega�t�%��'��,����n����y�D�<�{�M�%?C�7;�OX\%�-����5�N�ʊ�k]P�s{ FTT �h�aF6��6����_Zd��ﾋ�(�$���!)l�$C5%f�T2�a���(�T4�5�j�[j3l��<�� fT)�!��Qj�x��:Gg�qC��-}i�S,�.Z{� ���K�S?�v6VR�j��9̤뵻cQ+_����c�8�y
�	j�Z^Z��٨�(9���z�9YQQ+?�1�G�.�"�kN�z�����W�v���v4U��ƶ�GY����iy,��/o=z26ߨ����)�\9�ף:�T���C�ڎ��)g����g	���/ڜ��"��m�=''�1�/j��'//:Dͨ"�7T������p��[������:��x�Z��\gQ��2h��FgE\F�p����9x�9m�#��q~����(P�v}G*.���Y[!B�Wπq�;���"�̖C){��>%qNeG@,���4��r5܅�9�7�B:5u�)���""�*�뵖p�ݲ���=f�B�nL�u���@<󇂎3 F�GAv��}v�<MT����Cu���e߶g0�[��0�|�:'#��6�����˜o<�����}Q	�fq���ҡ�����n��;^��e���U�Uw��_.�¼۱�>f��m��S�OSom��7��M�x%寫�༯v��^aS��u巆Vu����;a*� ~u)�r��/:F4F[��z���ϗ\Pޠ� �2�!�u�Kv��żCoZh�]���R�9B.��h�����ی��Jx.:��/vNi�NFY�cCu� ���p���I{!�~|�{F�����g�^�I���,]o;���i�˲�:���4N�y믺�"��apkv�1�i��U���c4ný���~�w�����j�����E�~����o'lJ!G�^;��{������mD��=�{�N�@�IA��}G�[���j�ݕ��[�`:�x0& ���,r���z7���ed� jq���njK���y���x�o�8��K1���U6;����D6��A�Q�:U�ڪ��2viьw&OlI�Բ����f�M3�����:*�fӾ�4��dHH�'�]���g�N?.3p)��E���~�І�
�p�FYC�S>�[��d�;�wAi����ܺݐv��r��1{�n�ۮ�=�[;o:x`�]5�`����Ӡ5>�qp�)��=.w��ӻ�M����Y���n]�3r��>���4݁�CuJ�&���K5�#-nψ�4t@����ܘכ�	�m\^�-���t��O�c�7p�,���'L�Yǚ��"S��0��s��O�^��rf_3�ݢ����$q���v
�����]��?y���O��Y��_kFł�pfbڮ� r��ǋoPE�W1i?��t+O���4Ϗ8�sv����w�*�q^*{ˮ����ya,���a��e�������Zʳю�m��QQp�R�v���;.�>nj.y�����Ɠ�����(v\��O�rʚ�9�zʲ^�o��NZ�i�.����#1��1'���ޗ�G�fI�"�S7�:�}+v���Ue*<��:�mm8��7����n�k���r��u�	����'�7/�
�"^:�����q�9M7h6+K����@�9����i��u��Zj�r�boI;������'f!��.pe�r�"۴A��	Xi���d�����YݷM/-�*f�r�|4��Y@c�7V��@Y��v�"��.��9OϏc�{v�8�*����2㭯��J�=���/OU��h�簀��R�1���K>���-/=��Z�m`ݺ�2��b9#�Jn�4mV̑P��p�|�-i��9:�! �Lpyf��S_UD���:鞄7!��۷��w\�Y]�9�P�d�z���L@��{�5��f�p��gD���:O`����k�nc�@ueS��CGU����	�=v���ej��h��>�~��s�]!�t��"��^�W`\ܲhK#�v�J%El��tr��}^O�M�R�a��޽ee)����/���~l�d���k+��\��|�x�toA
L�:�N�fJ�̊eحD�X�3�+�#f��S֔�#�O!-|�¶�Y��(���d�N��D4cX�fj�������H��� 즅0.Y�#�УJ4=Gu�#'���6q��;E��!�-�z���9h���^q�D�7�[o�fQ���>]�P�|�Þ�Fݺ;Y���>5
�*`�t��{������KPod*P�+��l����ڔ�������l�.��	�w���5�;�a�Y7�\`P��U��p��xq����wW����e�l���w�So5�~Fm��,�h��bY�:�����`t:1�
���E���۷%�H흧+��5:7!���FXO�`w<۸���=T���1+��eE���q�1��//�]�C�s2��2q�sμpeu���`	f}�����r� ��UT��Ւ�ݬ�x�xn��vUaH�7F+dCl��kހ��t�ƠfV���Рq�>w��n!uc�<���MeTD�f`��R+��ǭ�Yw�(v�vU�睡s9��8u#p~K�.gu��R1��ɩ�6��t��D)C)����z��a�g>�p�dt�	݂����|e�25�i��T\ ��櫭*������ɝ�L�ܳ�KuռV+�Om����"t��ݩWcK�g'%�OSt��z�n|�g�w�B��6}qB}�f2�t9�r�2Y��z�rYU�l���_NG -�#�n_z	ǃ}}���^c��u�v���o{t)'.��g]A�j�%�I�|~&�n������a(�;�̀ڟQy�(�h�.�:&�:��r�O,���{ѮF�\����ў��Z��%�`6V�ĕ `4�����"�6�ŭRT2쬚-V)tuN�V	+F�uԋOd�� ���]R�`��	%0�|��������9ڹǼ|���>��{�M3Z��X@�6�v��7�M��WQ����n�|N(�by�t��cC7IM���R[ھ���9�Z[R�82G�p��^�hE�����wX ֫���"�8��`7/^�u������)e��WD,̕���&o1a\"��C�C��/��e��_p��"Q#��Ź֝�S�����K�X�&q�o^+.f2�1,�gEq#�.���S��v�L�޾;�*�8�t��W���I����a��2`�w��UO�-m�1�Zt��n��
u��|�m��Mife�	SO�O7A:�R�[\�3��j��/2�G
W|έY��to77�_\]�Ø�6%�O�8��Pܯ$��!��yo'�����kЫgX��	{�}l8���,f����6�N��/�i�fV������v��b2Vr�/�L9�����֕�逸�ӹk�^��u�g��gҾ�M�U�@� ���~^��J�m�N�=��7}6��r������_ҷ���$J��ُ�m��}��� ���k��U���XW	K��~�����yC���cU��Ddv�"�p�q���\.��]9��.�B1�YW�]�Ƭ�y�Xv:�1#���j��mD�0�q&�W]O_�i,�*��qJ\���f�T�n�����# �Ex�*X����%:�)�#Q]@y��S-to2�@G�ƾ�e��齓3�X��	c��YՌ�x����sh͏m���	�a���\��&�f�+g���0/�>����_"� W�0��^�^Wj�V�d��m���ʙx��W�o��m�jڦ��ӥ��3���'UNd��w�*-<��,`�� �uи�ZB��]��J�C14�+���h����#���x v���JcZ>��
pn�a�_�Q��F{��kFA����J'F����U�;5��&���}�<W&�1	����U9M[�̺��'M6���0qP ��'ՠN��i��)�`y��S��=���K�b[F��3��L���t2�v�f1�EN�Y���Ҧ0��.���)<�X���R������fri�����,} �+F(��2VW��Y¬�^���^��l���]����ɘUf��ᔲ:�|up�ڤL�� �ƕ�c�Y������Z��i�ݮ�4J4��p�}�<7&��wm�1�t]�N�M6/�a��R� A�O�qn�ʵ�|A�;�CX}�,Ev�����5���Ս X�0b\h���y;��X�����Yd���V_{;h�\��m���r��Iue>��[B��Vw�:��<xw�X�S��b�m��r,�,�}z��**JH��Op��()J��Jh
)�i)"
t��hh���	*����
����(���A�Hh&�4Z"(hHi�Hj"�
b�i���!*�"�)(���JiJ
)������b���U-D�F��!�1-4hCLA@�8��i*d���(�*h

���Z������RUD�R��S�DAH� �5�B������h�(
���B�$hZ�$
"
�����*$�(�"B�� ��P�,T�HSL�IT$IE)J[J�ihZ������뺶��a���{;�Z��R[��&n��dMV�����Yt�1��u7T �g�u_;�ib�O��%U��$N�>�	pv���՟�̟��,���X\%9�"=��>��N�<e�Z���<s{2@�*6����ʏ(c�U��*��k���
�Y�z��Z�֞�y	K6B!�(�5���a��^���;���76�uyK)��e��B��8
�f��ʅD	j��/>�H����e�lh�O�r.��_X�bn8�O�D��t�7/EK/�s�&���:��T�K�5?��Q�P�����&��Ddf��_T��|	SvI!��L	]�ʚ˄�}n�jǨ�r�UB��Z�ǫGe,�z���{����1Gk]�ӭ!�ڤ��a��J�H��#���ǧ#7;���'9�7��4��x�bz����bU�v�N�wĮ)�~p7\����D�lAJ���uT���n1�Oy���捂2*�n	�.�L
�Cc�k����9�v �Qu�:����K-�A ����:��9X:���9���:1�V�%�������:��C^�g�4FP��o�N�i�`!�*&Crq��O-�Ln*�*���>����#fc�b`7ʷ��US�[1ɕ��+AdF�E�d�ק��6�}�Ү�x;�Dr��љj�ݳ�:3ձ��b&tٍlǺv��I�ַ��*f�۴�#{޲z-�	0���=b�Bb�Q���}�X����ӆ5���O[osp�PP�6�m�r..��!�����1�K,S#8�./ݺa��s���2[�'���Xw�����
 ���<�ͭ�}Z �R��(�eq���_T[��u�	m��l�S۸�뜦��b��+r�q�Z��^��^��L.7�m�"Y(��K�|k��-����M����m��d�Ce\vY�{�n��'��p����]�Ӌ���0��[���<��kʧ�s�:��:���>��w㍾����X{����S$_[�0.��jw�+	
��$j�A�F�]є�z�DZ�y�~m��Ŷ|���ZS׺f��U
�	�}F}N�oVD��䨡�������f���Wq��D��Х�cG	ok�RʙtO,��)�Z�G���	j��f��Z^���wBF3Ɇ�{̣S$�z�m��(e�d��|�]<+^ࢪ˄���xj�Ɍ��(y��^_�F8�6�'#-�n�����C-n}�(�=�W��g�:s�E�Ze�ݝ#�Q��/����Z�����L'Ƨ�1黆�g�Xg�a:e��⥺�\*wPt\����S���
@���ʤ�x�F��Q_״Wb�������_�B�=��K@E����Iˣw���<d�h�oQ�7�������y����Q���,smf�����ͼ�ԇy��L�z�v5��19�8����^�Q�ጵ�k�$��9�D��+����_�E�n�6(Q�f��=��;]�!��8�#�U5gA=UU5\bp��r���ۮb�n w����g��M$X�j�sgԟ�e3B��</m�I���\�]eT�(�|k����~�P����U\��Y�k�;�6+�~�r�R���=�,w&G��:��9a-�j��U���N`�΀���9��r��p���	�:M3:��WO�gh����]�8z�g��O�v���D�t5�6L�	mw(���缺"�R7'��8xnP8�4�2Qi�V�Ю���(IU��ؘ����,Ϭ���Y��#��}��%�wDX�nؐ�T;���,�%Sӗ�{��g_E���R��5�^^��g�|����P���6?W;	m�Y�Y�n!Q<�k�����j����nm���C�7��$Tu���^�|�-i��-��[! 5C�x��8�UGS�3Vҧw->�]3C+�M�k�v�7)���v�7�j�ӽ��T�8B��?;&�� �㷙Փ�;qF�F�Y�W`���6��ʇ�������L�]�q��LLlU'S��}0f+�]:!{��^I���h[5旣�[�k0���=먖9�����.�0b�X.�*|����ϭ����	oJ7<�{���Ι�������W^+�����ח8P���e�������\&����'��h���l<!��͘9�Y��y�i�w�؞�>��m*P�-�[6"��
;>��"U3���5��U��KTJƶ��{��2�\\sU�Y����M����Nћ+����e�t�;p��,���<�\O50Ζǽ8��<r�3x��q\�6h
3���S�vZ�B�͌����ݕ���������nɾ��ax�~�g�٬�."S�|j~Ge��0"{�|:�T�e*(����OV�Q˧��KwByea�#��gб�P����$����c��<mgJq��v�^tq�+������m*�ܠry�p7��õǪ��Q�%q���m���F�����t�r0��ˣ?��x��u�+��u�9�^Fq��#�2^��,�A�;�ͥV��pZ;g��0�ۣ:���lt�K��_���l:+�o���=X�����σ���/ʞ83~���C��2�؇�inc\a�Dp�dn %�g�^�6j��wӑ���;?>�w��|r�#'������>�>�|���HN��?:�[5��.��B���$n���}O���j{%R2��N�hGm�V�н���|5\��AAAޫ�.��n&`�v.C5`��zA�4N>�'�'���h��o�+��rX�.ww9W����y2{9��7閼3|�5ǡ=)XVu�gwy̜�<\���n�^t�~]uA��Ɍ���4zặ��XP�]<Y�kO�{q(���(_��3B��Z�w���+��m��u�	ޣf�ѹfQ��FZ�rYS]FɛN�gg�K��'��KV��v�; ͷ >���J;
�ފ�o��	J���n��g^��\��+���R�n{WoSHegI�~��3L�м���j/Y1�]J8,Nt�u(!*�x�`��75��97�T�n�����]S<�;޻M:��^��)�tȆ�ڟ`ץ:�*+e��u����i޷[��K�fc�ʼO��1�l�dM=iB�Z{[BS�(PH������mC�aOSP敷�u�n�s<w)�-ɏ9�'�'ؠ/*&����5:Ge��G#:�4\,:�nӬ���K)η+��|���)�n�aK*anR~%0��فcL2V��~z���yl{���O{=Y�Uu�C���)�r^���uWT(�t�p�� %�-�7�d�0;fr\����U���m�w���c�c=�#,y��mRG-�R�TBr%�@�۳�9za���k��7פbOMK��\*=�R�[�ˢk��ә�h�{#�ȡ�i�ƒN[
��zo�ޜ�6N��cgso��5�*鴸\8�I��r&�k���'�gM���ki��/yv��Ė4ʍ���b������cɉ=��=�-�G��뗸u1 ��{���s�zۗ�O{�f�W��Ti��0����qf��晝t �ܠ�h]2\�lMK^q�gU�f���M��M��:s,J�/�v�Yu�*��?F�#y�Ͱ�ÍZK�.�1V=�əwї`Uֺ;��F����ϝ�,+�����oCŧ�я­���㡎Mv�وhb��m\��_���j�����K �K��]��<�uɨ�,����'�^.�6�u������8�еm]gH�w6D3m�9K��q��;h���������n�d�dJ�q��|���~��֭���_@���[]눖܄�����ϙu�	��3p�G<�!�8��s��Ơ��$ט�$|�s�O��u�Lh�0�N�<�̔p�k:���T>T�]�Ņ�ڌo(\��Lf9��t��o�9�ʴ��O��g��+�ɾt7w�Zye��V�Z���uZ�|����ܞ�Zk�rpmB�\*0(�G)ߴ��p������T��[qgS���wv���]�y�l��,�������P�zh�!�B���r��ެ�	�;{`��� ��v����N �Xk:����
ҥ,�7^V/�?(� ]���_i����N���Y���ٚ���{ژ���ߥVY��x'�3��
��f�x�p��Wm�m]����X�RGw�,.��Q8��!<�=��n�n��ї��ghV������4p�������'NP
�ϲ����@��}D�vT2"X��s]7*6�e8�0��o2}�i�fR����p�m��k.y�}c�F�j�զ�V^NM�k��ϩ�v��VT2�oF閲��4݁�uB�1�\t`���j����A݈�Í��ە��Q��H�`i-N����l�FOi��N�T��+�pg��m:%�O*�ېs1<�\�ϼg���W�䋎��)�(�7l
̌-�{�v���8M����)t���q���
�e�L�Ҟ9�Ͱi�v}��rE�j�sf����Cm�9�GzT�8�ڥ":��j�o>f9P��N���T�B��Πw(�u����5����8=��f��P{�VIn׊ܬ���5�C�9���׈ƙ=���Dϡ@��u}��O��H*��l�挜U���Gx����1�1�wb��g@ƻ�,:ׁm�F<3r��a.��̓��
^�wGL�B��nl*k{�{�s�P�-ӥ�%����;�u�-�� ظ�ז��Eۺ����3R�7���g7༴��
�2�Ͱ7g��i��y1�E�l\�3Z%f����n�j�,Ǔ�z�\ﯱf#M�#�ǌ��W����fc�kn������c�,\������̩ʊ�W��ų2B^<��|"��Vc}3.f;�1�H�?�0�2s��uq����E�f���尠�eS	c���3rR��=r�v-L�����)�qYhW���#���_x�k=0~��B5��9X��a���d��F��nfaR��Fa���P�n˓����F��{e�K*��jw�3��T���x�m=�ͳ[��0G6�H�m���~����Hp���;2k��Ge�[@�+UM�5��V�z(��&Y;���wCx�c�8�D3o>��r��B۶��ھ�!K'��xv)�N��r.���d�����'�j.��L�.�O�Nџf:��7k�u��|v*a�2j�>X���~<�.8���|?}�&ݸ�w-C5��Z���z)֧��63O�r@-}��O��K������~q�(��y��z������0;-�1�.��_IZr͍�uf��q��*��m�^����qʡKX���2��h�5���00KtuM
4�M�;;`z�k�~��m+5�EgǼ3�`䶩����G�B2�y@��H��@�g���Q�_�qG�/��T�7}[�r�	�ZU����Ax�f��LV�w��7ʈ���Dw�r�W���sԅ�o+ܰ�
[��V���7�y`�<H���y���Y:�'bw�կR�9��w �Kl�-�w_nH��_y��o��f�Mټ|���n��:e��1O�>���.�%u�p'\#���#x�Ԁ�Օ�Mg�hˈ��z�m�9�)w0�z�a�%Q���3����x���̍@����@��={R���:N��s1�r�f8AC��#�ݶ�N�X_�.�eq�������'��G9���*������[r�/�~n��D��AG)�>>z���oc�2�π���#��i	�ֲ*�q�;9l��J�������x~�x��2��1�g�Λ�~�n�/8P�/GZ��ǜ��Qqj���̵z@]���O9U�"�����1�k���l5�_�5�MoEQ��}���$�r_��1wF�/5���.����ފ�o��	J���w�G_:\���&`J;I�jbqOM��B���|�u����΀�S�/>�-uثE��i����/�sԕ%r��ן�<�?S���]��;�v�{S�atT�󦄰�O�fS�y�j��	@�0��g��Oj.���te�*O�K�#Z���-N�Oa���d!")(�=�����V�B�m�ȗj�d��.jm]l]���f;�@Tr�]o�eK��KiheY���m���=�pG�|�v�@OsC�3��^������E^W�����Qɒ�#��屠
%v�[y�r�v�Wy:��E�8M���ý�v�^��h�6��Ӛ��}�y��e��r�^w4t�S��#f���T@���/4�����6��E瑐�����^gTs�c��[s�O���d+��6[�[��[���gь�~��^��o^�{��rB���-���Ƅ;Ο0ϵ>]�En�S .��˄�m�X���������W���[��fy�4��-�x�2k�t�|Py7L	�9��A���w�x%�W	�p�B�.tت���%Q���n6�ؕ�9� l��qx�#s���x9Ӡ�vœ<���(�3���o�FA�Sp`KR~Ô��Q�2�X���py�rm�m5�S�^f�۵L6��#mӐ1�6��[�]��"��Z{�.5��1�ǣsc�v�[�63�A��V��ʇ����`#�!�����x�n�o4Yg���'�_u�7'e��ib���;�c���~��˺dc�eo!�!$L�=i�|��8�r���A�d驷��z�ƺ�q��6�� �ltp�g��t�k�s,���X��t���vf��]X��eU��1��4�z�ΝÎ��3b^�|c��"�:U���*'1f7R_�wsuh#��`�ߴ������5��{g��y�T[�(#˸�"��󥄫\Q<����U��K�Fr��Thnc*$4^��[˱7��Gd}����NE���Y>�;�}�.|9!�&��u��V���pdI�2�4kK�[;x� ZG`zĨL����6�ess�	�^�2gH��{N�&w���F��d�ol�#`�D�O����s.���@�.���k��Ԣ��F��kG �p{n��*���L^���!J{���T��ܾ���9�t�oL�ۺ－͜��:Gt��2�5�����׸�;�h�Q�`��Xr�NP���޷_�1&��*����(f:�#o���Dc˰����"uU���7}L��Uj�i��:(n��jPv�4R�Ŏ�.�t��ͧD+�����y~���*�#�zV<�S2�oq 3�mfh�][���K>x�͡����s���7�a�=�ϭ�T�f���T͡�SG������@�;����:Բ�0�5-�&����E�$��B�/E��Đ��>@ L��s.��;�]�vYQop��B����T�蚼�e��t���|��{t� uI�n�F�Q&�P6���ۑ��vp���D�`�"���Y���Bݚ�W:��!Q��&m���z���Qͣs��|�A�	h�)1/�Z���b����,x���x�`��i��b��R����;���hR�XҘ8L���+����DH�2�Ln�E�Eqod���T��)X�G��N�u=~� ¡^�^v�q���Q^h�+��g��sq�}X�2�Un���$
D<�=��\�*��_f�K��G��Si�c�0h������ jݮ$d�qj�z�Z�q��7%��n%��cF�t�Y���+"Y�\�+�D�1n�
�bw;Xmd�ZWM+읏'�BJ��ܐ�]��h�;�m�1��ᘥŉ�,j�p�=1+��R��Z/�sx��{N��X9����;�0��{�C���*�6�fV�Ͷ%�j�:�f������T�/{t_%��T;3p�p�NY]O�����(���yP�1�;�±X�l7�2���u0�9u���J�bN�ƻ��AM�o׳Nb��+�>��Rqo����4ad��E�[����HǚJdeӼ��1��B��#9[5ˇt5�zQ�@ւR���6w=�-��Pv)R�2v,��"�IeK+�G�+n��@vu��m��kL)O�:˺&�i�,�Æ<��j�6v!WM���S{Y��7�`ءc������)�wNW��;k�T����T�T�AML�UJ�IJ4L$m�"F�"�(Z
Ѩ��8�R ����&����������!b��b�")Jh	�(R�(��)���)5��(�(b�h)ր))��6�P���!BД$ES��I@�SAQ%@��Eh4�44TCTDR%�:B (�����B"���(������B���cj��] j�h)(�P)Z
���M:����MPvJC��K�HҔ�P��+l�Z
hu����& B��t,T&�[�)��(�UWP���Iї��>�P����:b-� 5֗��x7��������,�կ���w�<��{��^0��v9|	�H���Z<���>��]�����S�-�0�� ;6�Eq��qY.�O�vS�*�i�v7ek�fݻ���W�{�LX�~��P��p�|�H�N���f�,]o;�hO֞�b(�B���+� 	�ۛ7�|�mã���JG���ވ"�\*0&��jw�*����dp���<I�l)���΀��*_��^�b�:Z��cL�sH����:��N��Ӻ�xu��x�{���]Z�m�:��^�eo"+r;NG:���G
װ���tO* ���Z�ut��,�.Iۧ�'�n�6�V]k�e��;��k%�,O�m|ݒ�	o?WO
؋��`}nz������x�1�JbS�[Ҋ�;�so�V���z�w�S�Z�YP�y�N�Xy�hc7T�B�\t�)��""b�i}��'4���v|�
 \�GM
a(�|�Xbn�Y��a��N�V�x@��w��kCt��te�s����7L4r4Ŏ��$gWE	Ɣm��P�̌.���rg��P������.^�mX�0������3�/�@����;>�ʋ�,ER��2ԟ�eB���5��t�U;wCZ��b��*�y�X�ƞ��C��[���j>Xo�K����~Pڞ��|V�ME�}��1�CzƁ����?j���k7O�%&�5N/|�=��x�uڸe��37J�_H��D�f��%���9�q�F���u�����C��y�v�l\�4v)n����2�K���	9�*`!�W<��}������������[QoN9���wVc���ӱ��b�{ >��s8ӯ;�4�[r��0�q�`���Q��×g���"�9���ŕd�y�q؇B�]�W��Y�;X[�����MŪ�E�ׇ��r736�����
�{��������0-7�-��y_����ۮ�^$�������C�g@�w\;��^���'��\E��f��m\�� ��6?W;��p Ѣ�:}MxfdTSl�����~]P��{t�[��9���"m��'��rӁk��ś#Xk��i��b�ΰ6fT�}=e_<�]�'K+�����d�4)aeZ��t�|v�L�T!MKj�[sW�\p��0\�fĈհ��(�=\�P�5���6{ Bt�F�=@{b�QFa�[1���[Y�F��q{��<7�����SB}��k�Z�8K��	�v�:*��u��y0Z�=��b�W�;�����y�*�����E�\�͒�(�9eq�4˟��='�.}ی�t�K�ؑ,ne��9�X�f�]��EAZ�@��d�B�]��$�}Y�'��ޱ����cb7e��Z-o�7�t���������x�n�W;1>J�C_��G��|�V��sn+9�v�uX7���j��{֓o9�a������J���[%ϺC�;^�^���lS���NF���P�hفr͐�����<}N����PS��Z�ܬ5Դ{J�z��1��٬�q�<(ʌ��a��xI��L���SGL�dB�B�iF�?,��Ɣ�~5���`�r�'�s�##��O>�r;��]�ʬ��2���T\�������m��d��L��;�V�̲B}���g����O ����=N��xjw�^�����p�LƵ�D�V���}���<�J�w^ʎp</m�HG�|׎ j�.Ut�����YÚ����W�{ ����:P�U.�4�=��Tc`;(f΃s��=��ty�=H{M��f�v��k�ˎ����1H%	c�n�rpu�����Yw�(tle�y�3�<�z؞�u;-ƈ�9��[zB��p2��������r�#'��g����e��xk��GKp�X5�g�ٞ�6�Yۂy�6nN�=2�p� 5�VL�%���[�aB�t�f��o([�O�+vBߤ�F��9�Ő#۵��s�}-̲����*��~ɵ�:_�5�_�34;�G�iꥯ�����}z�g~�6�J^�,��om�g�흜vް�v�k	m*�rb�[f
��i��p��^�X#;:[�]�w��O�w��.i��8��M�Ms	3V:\�3J�&�j��l�P�rp/g! .=� ;jy��?YZϽ4-�6���eA�\��0{�_���D�ru��e�_��g�ۖ�jw�y��olw�s� ?�>��У��K�N���}6Ǝ0ڎ�TeZ}��w׎�_����Ń���`C5r�g�w��-N�������"4���4ҝqؚ�����uj�2�a2�(�ݐ%�=>��:uB�&���>�u��BS����zv]��WS�fA���,������l��NQk�g�<�� ��f��6T* O��x��:GZ�NY�8�k��ήq�U������>Y�.���Z���nRy�=�a�q,Cd,�3�oRS6�"���s{�x�����b�j�������ʻ$�P����n�kwV=���G����b��̎&�^���vY��gǞ���T�S\ňiQ	Ⱥ�|��h�s"#� tfs�	89������.�M��������n�w�✧�1�qЈq�O'����y|�wtY"=�-2���/�dz�M��-I�0Bo`C(���k衪��l��ׂu48����o��t��w���4<�^K�pt�u�l�7�p5mے�F���wʘV0��{K�a~��^=��6b��*pp�3��p�[����{�{�@�W�_H��1�.jPc���6r��]'(���u��t cɚ{�kD8q��m�$��.�I�]=hnf��S��?�nL�7�#UGAY���˼Fw9����1ͣc�28]�2Ո��-i��Qkj�	��w��Gs����7�%�W'���2�t�⬲������D���R��ڪ�͝H�豢&c��D+~s˝�q��'��8xnP��td�Y�{�iSǎ<žt�e�LG5�6�E�k)yl� V�G&8��@��}�=�%�z�>��m%F����j��Z|�3M����s���==��/�p�����y�%(��uE��Y��9�������W�5��zGw\�׺н��"��a��;�;O�8���\��[�㝲z͸*a�xT)��v�����r�Y�t�u:%#]�t����h�S�iU�w:��<�R��H�M謽�ޡ��`y��\���[+�$�m�gtS�Ӯ�6�R`];�*���s��M&�{΍����<ⷼ�3��J���M�ڔ8�B=�=-��<(}*�쵰ʆ�}�E�c^���6����T��i���_��b��8���vB%��xi�(���'�P�4�9.��U�I�W~�V{���JG��Og�#��R�Z�xS[�V�>ܨP�π䠛oD�cU�O��M1�kM.��4��~��!��rG��Hdt�<��{����tU�l���[M#�3�g3��չ��}y��{�~P.YF�0�z\�-N�k�eC)m��"��Ȧ�4����Uy������kO�����ts�ƼX�7>����D�4���ݯ7n�3�v��6��=&�e[ڻ����F�r��Q
�f�g�e���,��"ẺlP�J6��(t6d`��m����e]w=A��Kw�c�c�����[��vh]\�:�#�4v�DbedDjO�2��lޙk)�.ۍ�^%Y;�7M��u�#,y���6��,ˮ�9U��_�`v���5�=庐��GLR��uB���P���6���-���6�t!�y�e������<i��[���;�����S�qƧ�$�\�SN���Z��xۖ�k��0�z�x�e�fa	�s�_8�tE��dn$e��J���ODM�[��uF�r�?.���ע2�g��Moqo-e.쀟^t�KizD��ƣU�v���wc�fc��Q#���]��g��|�*���o��E�kN/�[
�aKc��)��AW�x�&#8ىKpgn۰�����.���맢�ܬFa�&Mn2�"��0��5��D
Iy̵�L�E��J�;�`��dk��y���A3A���T��˭�5���f��o(�fSΛ.�TM���4�ݨ3%��L��� ��zP�|�ˊ;>k�b��G6��t	�.�vMv\��u&�[n��Z����Wѽ7t=�b]gR��򰘰(v�bQ*�Bs�E����؞��ͩ�����fΊ)�r���Wb�{�V�5Y�j�DU�n�.��\s����0�)/ѧ�8��!s�#V�>�g��J3����nƈFT=v���wRd����ۮj���(Ӟ�t7����#�Ϩ�[N�#��Vŉ��tu<�\�	��D�K�DZ݋��QF_2x�3�9��R�aFu<��木d�FɏQ\s��.�	��igF4�+�j��7�'����#��7>�*6`\�)�(Ξ�N�٧��:�t�)�=��Tz	����z�{���{y͘nS��Zn9��H��[�8�l�ThSQ���;324�K��S�yE]����P�8u�9�6s��jk,���:�\����v�Dk�y���{ꬮ'�
]��;a�����{%�O ���D�FXO�4r2�n�oc��I�[�3Qё[7��c�y���(��j�;u��&��c�8;�dpc���].���v4������|���,��"�����3����5��h�F`;(l�0c���lt͛���.�'wF[�xۗ�0����� ����Ok����g-�����q��Z}�:�'wG]�Iy-�?S���us�*v�}M��x>W�#���t���p[�B�Ϣ����ռKyhs�ٷ��ߟ#'���w��n�rpu[���B˼5�9����_�N�^3��ׇ���nWe~Y����Dp~�}�M�3��;�|/<�g��oc�2�π�\ )6s�U��|�cu4^��VsH�qp�=���̹��5]��tsf�U�ppf��5��y�.K�x��X��]�����Y��F?2��\N�%����ܔ�:(^n���^��=>�=��������̬bxn���Fk�6d���p-c��8��ϒ�©�����_Y�	S�7����G�v�4n/ܤqj輯�ɠZ���mӖ�r�P�U�~+0g�x�k��,�b���`�,�����qui�tn��G+/b�َ���g��{N�N��鰸J[:dC6���Ŷ`�V��R�l��sM�9ۇ�+e��ܺ;��::��ͳ4uB�'���	jwZz��%�=�zR�[2�=]��[�,w-J�Nr~�>~�n��Ŗ�3��'� jw�-�aa���Rj�e���id��m�粹��b2�lh�{M�dp˧��M6�(d�JO����فc��H����=J��;�n�A������=�w`�n��ϔ]�-�0����x�O>ݚ��w�)s�z��yy����2�q"O<��>��od��[���Pvigj�M��aL�U��4�*2mCqM7lh��I�x\�vn��#���j��%�yv<}'9���S�/-Oö�0��Ϙgڟ*�vӌ��=8+��a�Ap��W#��j�N�� ��
��Y�n��Bx*:��\i�q���e>{�FY�=�����aƨS��'*w��S���>�Oc���4�[��9^��.���W��׻ )8����qd.)η]�����U�fOI�uˈ��%ȝp�n���:��L��0)�l�p��Q�i���=���T���ӎN���Ơ�~��=��{
���2-�i����	f)h�R�1u۵�3��	�㡣ڜo<�<�dnX9����wtn}��)�(���\P&���y�dZ�u߲7�_�x���6f8i%l�9�.w�=ĉn�0��8:�/Db�б��uػ�U먋3�<�<�d �c�����w!����v����۷mh���SS]��~\g�J�����A����6�X�<r��
�̀�!'j�e�\��	�5�c�y*��+��W\�i�нw�*�,�z��8���^(`�4=B�]��1�\��qW���)'wA��� a���]�I��Z�����9��;����أ��2��請A[�Y
�\K����f>Yr�gi������ё��mN3�S=�C���I�����-��PQY��ܮЛ�fJG�\ѻ� ,j�Ӣs�̿�����ѧ?M�y�#^n��z �T�Ljw�f��J�uu�0�틎�h�ܕ#�{8(n��
;y���[)vI��M���(zE=z:lN��+p=\f�ޮ��4��d�w����oVD�G�~��Zr����:8W��)l�\"�e�Y����=́��b�/�+�ja�� �8�����ʎ
�>�[��~Q��3����Nt�.d��K�Z���Y�:��s����/L��z\�4얼�eC)m��2�VF��=�5��TL@�n��1�b/"�D��s�6\Fm����r�
hUH�yj~�z�v[���CVjS�T��O1ͅ�������~.L�n���n�!���E{���ϭ��,�h�"㫦�
4�l��:ߴfMT�ƨ���Zn��w��i8�q�ڟ�.��YS��D	\��_�.��B0:��F�8���6�$�4�dVlO`K��Et"P�/�t�>����R�G�_a飴�;�6�X1OLHQQ%�n�`���n��r��ʎseY蜄,F�t7�r����^ wd� G*�p��H��ƺg���SB�:���z����%⭚[w`�mP��WJ6��t�ͥw23�Rh�R�"��N�Xj�:ݼo�������x��{i!nͧ6�G9aܲ%;�9��5����D�4
맼�"Z��{��*�Ufc;u�ݓ�X4~��>h=��22�:��
���:���2+�*�����vl�&#��6_/���іz�[��� �FJ�-��>��u��|�(�Wf%;'�.C���~�朶.Jj�YS��ȳVCSK�2Ck���g��WA���r��|�WB>��a�`M�������ռ�Τ�X�υvj�:��79<�m����;���K���^�t1뼝�,�."b��b�q�dr�2>��$�nǄ'#�6'��d�zs(��116ú]�{wn��<i��1C��h�_a���>n�)`V��YT��1wB�^�3�L����t=-��1�)\�`��ݭ�LG�Yoz�l�<��d�(�PEK;��<ǳ�^_a!������r���5�^Ü4�����绒p���e���N���-i���o���P���=wR��k��W
4�wq̘pN�3���H�ܹ�<�*3z�S+����v�j/�Q����7{�E�W\�]YQr�l���r�f�#�8t(ޢ��e+kG	�ul��\Ch�t^m�X�g.o�	���g+&έ���
��i�x�h�7��e�^����)�ߡsp�M'R�57mV�̣Bʉ����@Fh8-N��盖���?a�E,��B��[˒f���6-K�3n8��+��Rt^��h9{�*d�^��V�>&�ķ�i��YG2j8��=��/l�����S���֭��FQi������;�qw&�T���9�=�΅f�u�A_b��η��۲+��ղ�s�Et�.�w��}y������R_8�}Ը�.���c8N	n��9Y����;0/T�K�c>\�Lu�MI���
vt�f��o���:��D����ȯ8�7�$r��w�p��r�X����fm�5����\D8���ȫA��P�beo�^�u�a�����c�����}�tPN��*T����v�Q��4�7[��Y�g����؀;�2��s��(b�kݕ���u%�i|s�Q���gH���:�:N]��ER��2�'�wd���y$��iӼ���%��b�mR&�6�t���<]
��{�=؎yZ� tܠX�+A���\�8n?�-�;�z�ݎ
�M�j�7���k`j��n��4�c�ո_[u=ƴ^�ˋ8�|`�V�}�P���edĝ>}{�c�h�d�_���'�厜�y�������ű#��wb����f�-�n-��h�����t�n��Оl%�F.wm<�òʵ��E֚q�ۚ�]0hcfU�o)���KMP5#ݴr�^gLX1+VZ)�M�-�
���YRi3�gA�.�h����x]�!��^�e��x>i����!���&JE�R%<}��y�b�e����o<˹������t\���M	l�Jh
�쁢 ���E)���z��)�h��QP�5Z�

�)��C��4�%:֊�������E=i(B��Z
bJ�ZZM�[�UM]�RФ�5@QN�����K��äJ5�i((H����(Jj�JkB)
@����C��Ƃ����:]�((,d:M4�!JS%t�"b�&�R�we���
R����JP�C��S�t'@P�t�b���1/@ꢤ�h�4�����"����Ht��EH$UC�*B��ѥ:F��:((J�M�]���^��4���)w���;ر��V2v�L6�^�R(Jo����mJ�Uw{C������ߧ(�����p�-�n�,�1-Η�]���&wr�_�E|�-�/5�N�שׂ%�������݈~2�|�_e�3���K��Yf�Np�U�ֈ"0�*�D\p���PSOQ�-e.�e ��-��L�ʃ��C��܈�sr7�.9���tE��ۚ�p�c�����u눼=^��m\��P��{pYC:�$�n��l�ZaͱV�+Tv��K��e���YH9G=�a�q*:�p�|�s�U<��טjb�z'���2�! zc��j�·�E^v�-*�B�M��d�z:XY�ڴRavڮ.�O�-{���c�rw�3I�ޜ�\�D�հ��d��=}�<4bE�2D��4iy�[���+���\�s>�p{2�mE�jw�k�X��>��
�+fƲ����f�	Ln�fdV�9��A����X���R�amOZ��	s�d�%-�v����p�T�f������3����_Tzx�x��Pc����܊�l�8�=i��R;����� y��Q1S���*A�����U�ۙv9��:���s�+�äl뀯#�㺓"�(��ݖ�������e�]4n��է���Iw��dA�y���j���X%��ǯ�����gP���Х��/��i�r`u��Y����B=�>�b�8ṅ�F�
:땬�g���b]30�u�9%�}�3h��ŜD����SO�1���%k�'rV[�?�~�7��?f,8'y��ʷ#��U40��a�ܻG"`W�j�����Q:󢪯����/&a�/n&ycN�ݱ�ۏ�P�{~Dq�s=�x�R�.T#,98��Y׍S26B���7�eS�pv��먣LN�ʎp<-��4�:�	����˔�
sy�a�\��r4���fw�gP0��<H�9�t5Vӹ�*�a�U��3���m�x�F�l7��y\%��jr�y�j �j��/1�8�x�F�.,v��`x�B˼YC��2����ko4��q��\��wm�'O+ٔ:�-�v�s�����a��=F��w9��<�tZ��Ƕ���ݍ�XgN�h�5���?<�x���=�Ldn�:n|���t��XP�n�֏;Og1D�{���ݨ���,t1���@��w!9龊�Y�\P�뷜�m�4q���T2Sq��i�Yr��ڣ��yt첹}�������(ٷW���KgEs7�c�W�+n�3+��/��y�"ŝz�r-\d�];�=��Q�w�r���}E�GE<��@-��+^��G5�r*A��2�=�f�P�kU��U�H)t1veܽH�"����
�Q�-��ީ='�+q�t�l�w}'N�Y�Dd����w{��%�|nڑ�,e�3z��Wg%�'-���/C����Z�W�Wn�Xp=��`�R��pK�d��u��d:3�w%^O,�n��!�+�yjw��-N������U	��Z��l=�sH���Gm�I��=���2ϻS�r�U{� �J�A>6���VE҆S��Є	j}���Z' r�"�^��ޝ�k���?V�u{M�E���:L�P�ؠ-��Q��ñ{�z��ڻ����VY~f��*Z�(r4��O�otp����Q���>i�y�_M�,ue=,���J���ۮ�C�HT�����-�������9SvI!��L	e��,�a��9>�\��Nfl������ǯBx,�
��K^♮q�ĭZ��zڞ\p]�Y�w'ށ���&�ڸE�n��͜�4�xcS��;M\utت�^����_d7K=�i�|��횷$�re��د8��=쎀*�*#��w!i��m4d��Jn	�.�^
l����Vb��ݬ����^�ݥ���<ã��� J�� CtsC��[�M�ַ��`�VSf\���~���Z.�m��`Q�.1���p���8�}r��`!�Q-��~�M�_����^��]Z���c�?�Ԑe���}M�↊h���oQ��{��}���%���2&A��P̙Ϩ��k7$	dhů#�r��%�y\�o�����r��B�*͈'���b�J��n	���%�X�B���vs33r�(�Wt�����Pj�'N��I���k��R�Q��}<���!�fc��k�DE��s����ϖ��f\�ˇ�	j�BM0��O����!K+4�qw,��Ql.6�� ���u޸��A��KӞYܠ]B�l��}yU};��ܬC����td8��\�7Wر╇�g�>����]�O�6�녉����&�9�Q��Sb9\^�T��]",%q*<�'Q7��֜Zyl.:�U�2�Hָy��[��z�k�v�+w�R|]�-���/�Y[�)踰v��H�W
�	�S���:������$���f�q�>��"{a����ίe�i��im��n��5�5�<���@�Zl�֘�]����FVmGd�����S��Ȑ��by��M�C���tp�װ����'<�����5�a��U�}�m��������T��}N�-4�/�N(�3��߲���xJh��8צ;�u�^VԿ9�\o?t�ւ��S	�����얼�T2�}ӭea�c�@�T�u�#>�̞Q>����S��ˀ��[��8��*�!M
�iG�_Z�!��=�����z�kX��Q	��M:7����[��h����^4R��H�J�
��(d��k�h��t�p�g�d��o�v���F=��&ҁ�n\�޳�^�;:�$а���������ו�JȠ�w��Z�wP�sSX]ZY�e�c��9���s���?���<��U�X�*�PtS7;?#6��SE���BE�Q�nd-΄%�<�=Lf�5�㧒�#��m��
~8��O�)n��v�Qā֙�g���P�L����-�U�5����3��~��Шm~'�m�i�q�����,eU�,%�k�\g'<���W�U�@ډ�k��?N9e5Qnl+=�����t#۽'��]�q�m{�6��
��i�ݩg��̸ݗ�p��Kx��*�]�9�*�xk�\c�3Kk������*nǷ�ˌ��jw22�����ĉnVa��(Vh��OQAKUDa�(qw�Y@?�'�����i�-�1�y|����}T@�̃�}n�.[����;��]�\�d�w�=��"̵��w
�鎐�D]��K �(�a�\�%dvs�gT5���������5�4oTA}q8xuC�*�c��:3P�͒�V�+;!¼~ [m��^��SwE�͓���V�Xi��֬��]:�L&'/���`ڮa'��]L	�{�-I�ޖ�p��<m[<�u��p��~�z�{�7d���Q�l,k�t�ӱ\�O+�^@j�S��q��&��5��.�l�]�x,�54A[�_ڲhܻӷ��z_��t{�[���r����`7���c�+5VwWRf�ંo{�V*6E��"���N#"��bLJj�<�*�}f�omR�o-�jG��̼מo����u-`Cu���j/��;��4͎�)l�4%��;qjP�PY���hJz1�h�|͍�V��#�c4�68�<h	=F��Ԫ�T�� ����]���;F5����
� \�m�+oyA�<��	S���:9^Y)2�� Y^��-������<Z�#������kxw˻������פ��{�q��'�߸�.̧�����NxK�HDY07ԙ�B�E�6��:m^�FZ&:��2~¥�#'���6��וnGuB��k��YXc��[��Y,����}��m�h���$q��ow��|����0d��R�?�zx�SN��_=�����W����]�f]3�m
yD�Z�߃�`��p~�oe�~	������ځ��h���//�K���sq2��pˮH��8�����9mg]Ի�
�Y�bU�le�wkv<]7t�� ���OH
��?9x�R	�,a��t������x�VK���;��F��&�9��R#2���d�v�bp�wAs27 w�����8��{����oc�9���ܙrP5s�^	�%��)N_���:�_��ѻ�Ε.V밙!�2�VR��i`^��a
����U��C���G��>t*������)�����ȱ��+ל��;�:�X �,f�n*�];^�~~��[4��������M�a�����no�~����e~�0�W���[�����	��L�3����o+�?]7^ۭ��ok�N~����C�i�̵󡏏�it@��w!9�k�neu�	޻y�9э,�����εV���R�FZ�䲹}���p/��8x�
m���?aR��A9[�������Ӿ�k����¤%Nt�yt�)�P���h�w�y���Q�w�y��}E��pf�ri�im�S�6��U�]�tb�}:�w��P;��%t�4�i�Z��Q�.{���`�l�9�ջ+6��~����2���e�/�i� D�t�l�P��f��(C=56��bx���twN����f���΄i���7���_�e�k^-���%p�f��,d�H���~��s�oq��U�DT����;F#�lO�r� �]-�5�)eL-�O�ʗ���E��V�+��N/ޫ�;r���� KU:����Ϫ3
쎍҆]PEU;0�cC>�j�
���s#TS�gqp��5[�G<�duU
bik�U�.3��?"8�6d�܇�Q;����m�=J�Cv'5و���� %.�w��aQeD)Π%�5`���S�I䧬��DA�޻o��0'��\h���gx=ݓ�:ȇ	w��H׀���h������Z��0� ;�J��Ȑ�.���7��{���d�^�S���DP�f]R�S�r98�5�>��nE[utت�5��f�Tb�7`쓚�� �s>DqՇ+gws�}��e�\����"<�㿔}��U=dk��Le�jO�r�خ~h�q�d5���˝���P�:��,y��϶�t��z9�X��gx�
�:ss�R��ݔ�-�e�f��b��	��AG{#��rxSn��ij��Qq�m�,�%�O'���(:2�w�R��ؽ̜I�^_�kb�S{�g9���C��?
f�r��q�ys��9^Ǧ��+���e>�N}-��
�Z����ˠ{�m��Vi���[��"��\q��:8_��"3rP~1q�ŕ�QD�:!�oc���~�=�"�l��u m�e*[�r���qf��尦�
���=
Zf��ng]ۑ�8�*��Pp�r�#0�t�{M�$Ty���&��S�[�q���N��u�6؎`�{�R�����q������%ٔ�m�J�~'����vzd��p���z�a,�g�r�2p�t�{����p��#��Z�>4(��L��[+�$�m�gtuC�)��07���@|�8�{�5	�GRu1���e��� �oT�Wbt����C�ݦ��(���p�}o+A��@��q�����x��/��g{BN�á<���գr��3�Ý±Wd������Z�Ǡ�����h}�.�t��sKv\�]w����X���ixwVD���by�|ai�lP�}3ͯ�z��A��A�
�?Cl�r�ܫ�����)�v��� KU>�-N�-4�/�N(�8��n�C�A�Q��L���v�e��'����Yq���[�5�\�B�a5P���;%�5��z7M��}lvڮy�4r���V.1��:8i��)�H`���聸�$K	GC�5?v�Ԭ�~�2�z�q�sR�Y�cr�5s>F#,�{	�>V犖�q
�����۳�YQrEǛ���m���sYe�J�Z�e�����̌
Y��]��~8��=wL��X,;�x������_�[���\���m�BX� �s��xTk�<6��F��~eu����|�7^T��k!��a������M׷1zk���T[�����9X���6�0˜���@�9Cft#"f#����8z��K �}P	��03����YS]�9������\v!Эw<r.q@h�<`�3oc[;6�P�DX��q"Vه�����+�QAM=F=�Ĺ���{2����oZ���e��w�	�c���(e� ��_:��}�!�*߈^���'lե~.���s{;�G%��}.o�;R�IA���h���}o��-f����|(Q�&�M��ٓX ���7��XN�N�j���CY�o��n��L�B�i�Rt3�o�c��gO�<k��<yv�	�w9f�����t�8:�ބY��[�Q�
�'ǍƝ����������q���n:�}ΨkynˣE�ܬFa�t9�{Jd�h�dC��P����;#���pk��*� }S}�;
�ltм���-*�B�p���:`����}�(=m�uw/o f�?W�#�if?���l�\�tЕ���B����Y(h̶�n/_����Mz�ݨ�=#{�kϺ�;O��+UM�_D3J~ƛ�S�Q"y�������U��)���n�v�	�"�-�tv�}BE�
����T�}OZ�h�+�NT2Q�/�v7$��p�w�OE�vwy����c�9��(;Π��0.Y��OZx=ct���@h�7����\̞Fw(�-j߬��ُ.�����Jl:FZ� ���v�%]�,s������,��~�󣣘ҎG����K��to)�S�O��-��9�5�~�d,�2r�\��0��Z_��v��yi����ۼ�c�Ήr����l�L3��������{���TE��*"��@TEr�+�@_�@TE򀨊��DW��
���_��*"�ꀨ��@TEr�+� TE��+�P_�������+�P_� TE}�*"��1AY&SYQg� a8_�rY��=�ݐ?���`b�����JJ�j=����(km��{�h5�Qh4 ��uL&�kmU�
e��h9���3:�ՃJZ�֗��ච�2)��۸���s����RE9�;k5V�b�,p�kZ�m�5�����m����i�e����[B�M�l��6�T���eB��mV�͢mB����n�i65��fZ� n9ܲ���ɐ�*��
� ���ҕ$�F A�i�& Њ~CR�Q� L #  ��&MLL`���~%J���a40��0�bb���0�D�LF��e0M&	�G��&�M��A&�R�ښ�ɑ�4�   j��v�{�沔���*��KB��f|�RA!		?iI d��!	 LX�_���1�=�>6���D �T<	�z I ~0�A�RB�*��ƺ�(X�Ӈ?=��B�?��?��d��?�a�,����?M�����!M�9u�ΐn�]S�{��ô���Xn��;��Ie%��b��l�-�B��t1ڭ��fh��d��h�h�j�A��U*�	�j�^�n���T]4����5׬�j�wMX�Q� ���*��$���ݚnb����[��)M�l�b����Ck(�����`v���.^��n�*X1>�R�Yw����k^!��p8�v��e��T���-L(�f�T��3&խ4���T�j4���N:f��ѱ��L�Ğ+ʹn�1+��QR��X�������b���e��=�inc��
��ژv��٭�Ml��;��n�4;��SF�T���f���[��]<ySt���0Jn�dL����lL�h����U�� �C�Ֆ�&�����t���Z��s*���%4$Z.��۷�&�Paנ_�I��T!Y��\2}��ڋ]��OE5�B6�s#5.�b��6P�����tVm�S�B85��q�Y��Z�ˈ2� �B���3��ޚeX7���]h���s��|���L�4�6�S-a���P��������Z, H55�w2Aܥ�dJDls(E�~��o�O�u�g,����f����[���d=[���� V� j[�olMI����T�F��0���r����d���٬9m���B�O�&n6��a��!�;�Ď����[��4]E2�_(傢0���V��\5[W�a�3-��v�\P� ����p�tR�U�+l��U���,���&���b�
�7�54;��ejh���H��!��Өnd�y���iɬҴ�زI:����;;Jӭe�36�W҂B��_8ӻ4�ӛG .�6��EǠn�Mݚ�[�Y��'�QXL;�#�&����;�e+�Vn�X�T�"�m]a�L�Sly��&%�K\ATd���w@���cײ[�09���)6K��eY�{2�?��%n�X��u��u�b�EY��m"t2QE��2�t�).�?#t����q����-�7�m�TO,n� �azһd&����J�7Ct�������W�P�m��^֍��Yd)�M\���]���w��ֿ??�?����d��x�%?�#�O��l�۽�����������b����x��f���Y�����h����Ǖr�G�E%wW>fh���p�� �����Vx����O/;bk|�Z�.���ݖE�q.^a��յ6��tB��zek�M�p\�u_՛eރ [�j�I��F�9�m?M��E+m�����T.������4��2�s\K�x��z��n�SlV>������
��ۂ�P�EKy/kT�Ŋ%�����*����ċf�,3Q�e�^<��ȴ?����2*99��]Y}�f�nV��[�j�%ʛۜrh^����p�&�j��"�n"�sV�.�>�P=���;��Pk,�M>/�B\ׂ� b+mlR�a��(��[l�,�h�佳7�]qW����9�2X�����*�<* 5�l��!��/7��ph�'�NRlJ�S�m.�K0vN�sm+��9�4닇5/��bq��9�����w.T�.uj7�;1d�,ݑV�3��*1/nUs�S�GtU��:Ő��{~��=0Ix������ڻ7Z�x�^<�\5w>���Ld-����,��Qgka�%���o>W��*��:�,��wW�\��r���x���:�s긱X�{ڞ\Mf:hOr�����&.�m6��ivQ�J�H�J�aM�9��B<<�^���G�Gz�+���(��ݫ�}�ٲ��˜��7��Tʧ���W݆:�sg��
�e
2�4�.�ڋ��VfT�U��t�=����x���-ǂ��5�0hƋTj���\�,����/&%Ԇu ��V�s<[
S�{{w�u�����v�y�\������X���ӭ�h�6�ZZ����Җ�ۭ;�2������ �Jܬ���'�wY��F��%?fud휺Ns�S'C���Wj�c�7�b�Y�[O*�P���Y��u�4��p���f��(�8��b|���)Ǡ��F�%H@Un�D��>F�K�ty^�hjn�t�����p"�(�O��ƯL��TC<��ErO�c"k�}g�ClV���L���S-Q�@p���uR_(]�ñU�a�6�q2�<Ij�úz�k5�w�xN�p;�Nt�/�����?����31�8����	���E�h��-9Mc�Cq��i�a��-3��B��F�;#��f���"Ŕ�R�qd�3��;�>0�]o)_:[p���@�o;!���T�qft�=�ò��M�1��3J��#u�B(�����u)E���/ge[Ȣ�!x��
t׌�5���/�Ws�,�aG��>&n'\�b���ޤ3,;ԅ���JB�p����|�?nM��[%�^n�F�h��)��]o��ڵMOj��gR��u.��Ӗ��Q��wd-��\��i��*�SӰŎ��3��� ��1o:go< �x.��2�0��"r6c�}��<���L5g�Ve�b��n6�.Ƥw�F�Ng�L�]uϮ5�p���x*�ݘ�Q��s����`D��j�m�X�<�T��R�l�x� czS" ���I΅X��^�:��ү����}�MQ�>��:n��\�:>:¤i��4��:n�1s�mR���9����*���tU(�EW�s�EI+�G�v�l�G���N�d�m�2�Y��n��n�KfՂ>�oz*����oY�j���`甯c [�x�T�(gb�v��q�P�\Z�)�-yb�v9����u<4n��M%���t��:jý�u� �$��z�R���5�s:t��]�M�Y�����	$+@/
"ǃ���S	�'"K�L��7�/r�+��m�Q���kޫ���5%g��4�ŏ������L
%tV�I��074mL�[��x�~R);a�*���-�c&um\(`�P X&�&����ŢLQ
7��jn�ѥ��������%9V���5��fU�*���tKs0Is�ɔ�\A�FLKr0(|�"�z��o4B�Բu��[�	T]-�4���`��Z]ٮRt�]�;V1R��aj^����M�W�A�Gy*y�j�Y�ҫ��-�ۥ�N�LZ,r��ٮ�sZ/D���y��M\�%�oXt�w�[u�%�	[ N���hJ3�1���[]�7HbF-�R�͇E�f�7�P�֨�\e�D�$Ӈ��a/��#C�n����;l�*��I�����	�vQɍ}5p����p���g�-�] ��l5�0��S[$�;RxՐm��ݫu�[�SӘa�&��	�! IX/��d2A�����T~�o���:�^m?�(�d�E�]<`�nk���]�w�L=X���HL�{�*��T�Թ#�lYaf	���x[N[�_9�T
����b�b]�A]�������;�S���/f�����sװ�ӖY����6)�v��e���;�l��X1���0E�J+ذYm���h\�DTUTʲ,+�H�V%,�#
�+�����7����l����dqUe���s�t?�m���ЍJD~��Uy��3�\���ɕ^wx͂������z����d�'��� =��4�~����ټ�Ǫ���𲕹�ϰf;m����
���6>����mMy�G�t�wϷl=V��feN:!^����m�cg+��>m��ռ�r�;� 宱ZŦ�ZNC�W�1�����Ļq��:�0uf����1u3�!b�ڄ����W��ke^RQ��u犝�Z�~ܺGʼ�|��D��yM��!�6.V{��	X�4�7����_��t�v¶a���OW��1���(���zo��.I�S������Ȃ҂NR1��Y�Yx��T�wV����1�ز�']�I��{�[X�;�z���U����g���^Ȝ����Q"L^v�}�օ@���Vо[ul����d�{SfxAՕf[��nk�[��|1x^��@�u��[=�s}�LɁxXS��9��q�9[�ݙ����x��nÓ��Q���??)��)�r,$Fe߫f![VtR��Ϩ,/�=~���_j_T�I�9���%t����>������u��%��u_��B��}��QP��x�-��V����=�	នT�J��ת-��L��՜��
~�
����I�Œ��}�,YK�F`����We=�i���>v�C��<x�ƫ�b�b�m1c(v�(ŗ՛ݵ�3)<x_B�(Ў�>򞼰_y�w��s��v�����}o�I���M��G�Yd_���ً� �=�;����oVa\�`
�3N׌O���}��{;#��)2�>*��+Rʺ��λ�ȥ9���t}����Os��j�A�^�Ln��y_����99��MVV|5K+��S��t��r5F�H	p���~|�>������g�Md��(��^���o6�l=ڗix�0���m��p"�Kp��i�&����W3������/�rCk,�#���q�"H��d\��'t���)+D�=��=A,ǂmL���Ȍxy�p�N�m;���>�c��W:���Z!��	n��R�%D���DʗJ�ʸ,�9wd���j ��$_�c��������#�WD䄩u( 0E.8�c6�F�wrK ��`f1M&��+M̒�\�61���N���������FB��P-�aY(����*QZ��@ @�O� �z�_=Sy��VgW��Cf5]�m޻��F��^[70��XuZ0Y�=�l��!�l��-b��3���7Ƚ��F��O��%������l���|I��ޓ(�-	�����%���|g**Hb��O���*һ�X��4���N���_�s����צ�a}ETzqjh֬W�s+��/۾�.e��MPO;R����;��Ugk;w[�Y�.�:�;��nR_z={ބ�VM$��bBu��^w�n���d�$�.�!� �$�$�I;�������N$	�$6��	��d�$7��{�	@'�O�������&��ԐX V@����~7�C��X�'�I6���5�@��0'�C�ChO}��d��C��ϵ�`~0�{�HC�Hk�I1$��ޟ=�}�����01����5��N9M�D�JW#�����*I>a&��ya!�$4��齐I�+$�d4�
�X�m��P i��$�$��	�>�T{Ѳ}�D���s�!���pH��4�T8Ha�T�{Z�[s���ۣ�Fx�P]\�4���D��XM^����������s�����Ԥ����}�ݫ��a�و�ɉi�-�P5��n6I���&N�-����&_�_�ܢf
詎�O�c�}��?iY�X�+n��)�|�1�7w<�9)�TcUԑ:ggU��a825���g���VI��3�ڽ� �Wv˝�'N׎��('1*�1xy�x=K��촨-���k�e���B�%�ۙ˟c�f��u�"�K�_�{�!���=����^�~�>p��x m���L�U1�|+�k��4�o��7���y$��H��((�5ѹ}�(M����F�SE�O\f)�i�[�t��,�0�U��Q�>&�"&x, �a�!��u�1r��iuT���-����9f��,�j*u�:�K��8����yː��#���Y�VJ���s�bq\�6.r9�\uf9�*����%�~�)�ʔ�3�+�O�����?�Rov��~w`qq[�vP ��GOUtk��T0�]��~,�:�Z�՝���nߙX��U�,$��ə���#Y+�|�� ^N����r��r����N�NIAj�_#�r��$��r6��'/3�n.��`j�3�_]������z�n�ι���9�r_j<�F�:�rg
x��*R�[b�)F��^��h�L̷��L8���]Ɓ��?�YF<�AһL*�)�;����]4�H�(e]�.�����9vm(���S��������efP1��dǎc�Vn\k27���XۡYg)�2�v�,e�u�7��կǼ�a+E�-�,-�,X	majZ����X�R�Ȣ�� �J����~�u����w̡ܹ?~�=����q����b��䈯?q�,o��
˵z��`�bTJn��Y��I"�q�׋Dz>�Y^	���=~��w[c���sٶ���ce	��Bɲ*�����]xP��0��� ���E�"k�O=|����À]�7��椔��WP�Z��+�h�-c[�Y�%��{m�{z��^��-�-�FL���
�J�3YB��~/t���|�&�����yt�S�mjɏ��w�v��?3Of���/u|51����I��z}�غNyz�33��i�Ʉ�̧����g�]:��q�~5�b�b�*N�+�L+�����Y(u��{{p�{���|>b1�v�q6#��y�\���8Ԟ0F)W�=B���H"$T�}��Vn��T��\k6��oy̟'�݊T2���旎=eLC��Cl��z�3��'c�i�u7�����=fݳH_)����'KqSo̺��s�߷�&'ɦ~eLB��y��7Nk��p5am�V�%4�.��szw�>�ߪ������>�����}�!�13���&e�9f���?76��UM�㧎���{�����1<f3���>>!�*�1�o7No�<m
ͳ|9e�9�;���,�Mj�>d�m�+�4�)�x�fݱ����+�m4�Xk��b ��a�|aY�ٍ�r�ap��9��]��n�f��r��=�G���m�D]>�����(sT?O������6u�>8�ea��Sė)�i��L������S�n����n3�b�u�BǰG��D� ��0�+<n���%Lj(�t�}C��eM�^��C������[�׉6��/n������!U��ˮ򏰳biⷚ��w�M�ވ��@�"!���l����n�b{��m�Ͱ�N�Z��κO͋_ԅV3�U�PT+����&�
����i��|�x)�i��jC�ǉ��k�,���T�a]�k�~���'P��+�7e�+���k�� �C��$"PYʼI�f��y�8|�DH�4|Y�>B�
�/.t�OԻ*�ײ�v^�-�;����"v�h=�<���[����:�ى�+>��j�ǉ��fS>��i{�7�QN!��=��5�P��i���OC��g,�̘�$�+����w���
���}���<�������$�k.����f����>�0�B��ӷBf��^]!�/{�v=q�Ǩ{�m=M�wY���$��{Wy�5V����#7�y~Y����m�CN�߼�8�M��|͸�T������g^���]�W��ow.k8�7E�o�c���ꚥ&|~H��
�iW�X�c�*��T�W�*�^�~�Ξ!P�e�������N}߾��i+6�1=f�yۭx��u�E1(���^h~�N���B���G��f@�1�]��e�R��Į��M�z��[�DG����3���`��|}�=B:��gZ��P����4��q��C�Xq�*bq���;��n�P��2�}�z�C��u���a��7�:�;O��x�l�i4�ex�{�3t{L��8�x���[��B�a���16�����R���1�x�:�=�;������%�1�Oh��I�9$f���Su�X����xW1SjC�yU8�mU՝=�:�.��-�kJ۳B.vi�v�Ե�ؗs1R����	�ݙ �J�Qh�W[csMC�9l ��	��ݙ�iv�]�ٻ8-xEo�x��ʼ���n9aRj���Ñ&�DP��1�Z��g�YIE[�1H�:iZ��eFّ���r�v1��@�伬�f�#ku����OS���TU ��\IRVE�XVV
��-�ڠV�
���"T�R���*Ȉ�K�F**F��BШ��Ŷ���KeX�2(��>5�>���{�o�����g}>O�2꟢hc*g��<��s�3��hT��u�����8�=�����)�3r�N���4u>x�Cl������:��;N���u���La_��`ӟӐ-���<G������F3�N	�Q���M;Wz���<M'���1�=��x"˔�wT�C�o���E���d�cf�ZKq��)��⭑����G� X��c�D��D��M:=������LM�����/ܖ��>��"$y�T�c5�8b,F�2���}��h�6�λxʛB������ۦV���o���8�Lm���x�fһ��a׈b{�7|z����tE�LCc�Y���L�(�#H"��S�i�0�j$�_DDDC�G��(~�J��9�i�h�z��_3	�L��2��m�.��;˷i��"kܩ���"E��F�A���1���뙘b�P��u�b$Dh�곿Y���;�y����&�|e݆���}����i�ěg�;����SIY�O��w�h�gX?S7J���+"��¡F�O�S|�1ѭ�\1N�䐄�|� ~%a��x��5����S�T����u+�ӏ Z�~g�w��ĩ���m�d�I�k	�������M*�p!�h�xE�����<��$K|r�l���(q����͗�����Eը�$�9�l��q�D}��!���r���Ga+E1O���.Jz��P�FT�Re����ϘJ�Kz�\lB�/S���[Q'ja�H��!S�T8�r�Լ���5G��&��"|Z]��+l5d���n�#�������˶|�mxz��섡��JB�W��Ho�ٱnL$E���+�X�r�������?G��xo�bG�9�@�c>�nf���M�k���{m�&ۮ嫗���h0�	�VItU��B��Q�����YZ�ıbCj�,�9���ou��M��G�_�\������H	ɝ������<X]�i2��K��b�6�%py�P�F���Y��� ���V(�
�wc�T��̶Jq�S����nq}�{��{>��P�#���;& �uH~	?>�k,#h�3�P
�;�v8G����i<�[=3��m����5��uA��G.)���\���d��ck\f�x��������ʔ��ynʻ�8��q9�V�� �,'6�����=��wܵ�L��@��+��A����1���m�TW��ۍw�)�,�~�]���5orL즯��uҋ�*ȅՑ�N;-��uu�W�cܜ%p��IF.i�&	��{������2�_��9���v_TՓ�uv鵴�fvY7
��j�������U�I���6���牆N���
6Z�i�f�C���;���5f�m~��L1K��vY����b�RH�(*���ޥ�xR7k��˜�D]�����*M�ǽ�q���.N�{��'E��c0` �B�0Q^ұF1T�
*�#PEPj[edX���P����"���Q�Ң�T*�R(�**��F
��XV6�PAEdF
�De��TJʈ��b[h�X�Q�U�"��[r�3,�
&YD�w7��һy�^[Ż�DDDM�i���S�_j��omFhRԴ�b+ӈ߼�H�b�s�~)�wPiJ��yJ�ѵ�.Su༞��T
j��nxaÊ��"������-��1;���DE�W�a�?]�\�]���	�<�.]w�������*R��u9c��
�?t�|Eh6>�։cۜĎ�y)yGka𜦥�J��`��ǝ����j{��軶��R���%�I}���v�ze�a��~�3͈�{���A��k���WE�l����pJ�锴�ɱ$i#q�u�u�x�O.��^o>ő��������C0�Y�ikF��r.����l0��1��:����m� �]Z��g&�i��y�gY�Я7�({�5����1@Q����U{���o~��g+��C���zc��h-L���;����a��]����[L��M���آ��<�K�<���M�2P�5,'S�툫ج�����C���;����wr���}Tdב� C	��m |	 ���m���5�Q�mI˳;'åv�q�~�b;�v;땾|���'� �r��&jQv����Ѧj��sm��@Rr����DG�\�4=B�VxI���	}o��v�e��$�:��=~J<U䴣Z�K�0�]�Q�x�2:��wZ��<��	wI���%9wv����}���I����^m�E��H|���洑o�
�DSaV`���l�8�r����f�9�B/,��T��3!�Yٞ���yM�pm�� }O�똞����i}Hf ��s߆�O*~���p1�3��Ѯ�!���Uߩ�b��7j���X�~�ygVG��gd�����c]>y/���:��Ȫ׍�v�7^E���ވG�f�	�Ͽ=Œ0)٠R��s	T�U�Z��<��S�_e�p5�y������mTx*����6�WmK;�IBa�qqa7ZZ���9k�p,Հ@�g.�p�]�4�:K���2k_)N�ݕ���[�u`����������uܷz �4B��j����~�'�����d1�U��Sfh�lc�(�S)\���	]ϟnS�U�Uu�b��is��ǹ��W8m��������&n؆��R��+�4�ro�ݬXbUl�̻ʌ�]��cel�X����rq�.N���̉fEJ��E��p��ع�<�u���DL5"��|�3D_,*��V���yb���%U��2�EeKh[kkD`�-�Z1`,�SR�fF���,(�B�XQ1�YC*��IL�ɉ�R�H�0" ��Y�w�urǚ�ן��"��(�r)�D�t���dd���8�����D��p��2j�v��%j�1���G���wq���R�B2�`���͛|%@i]UV�swz�M8�·����""2�G�y����Ȃ�w�ӠT���6�K����ګF�_kKq�L�d�fR��)rr�/Z"$s!b�A׎B��	��~H�ܱ�]�i�yu%S��5cgcz/�G�*�M��#�S0�$V#�'��9��]U,���F>ʔ#�ߛ�,.���x��I4�z{ь9l�IE"��W�_}�r���F`q��E��c2���; j�5u��ʣ�z�0���[$\}^���V���%f�$z�v���
0(|���ƞ�����r?��=�{老�ڦ�feg�.f-<��Z��u���+�n�UՏ%��}����>���?c��RW�
nz��Ѵ�7�f��M���zI�����ވ�Z��q�I�SJ:��(� \����Z���G8`�z��@5�`�����lж`�����T!��+���5�y&�˯e�(�_R�f��(���ýL���D��� p�6O�S?g5|0X�|+3_)}�zFv#���g�OKڛ�;a;s]ӽ��Y*���폇3!vއC���0�gc���7ڦJڬM�fa�G�wV�B�ZĻ��{1n����G ��8ϻ��Y�1PDݺ)�C��:8�vȹ}91����L�x���"���ws[����=b���
�ޢ��u�5�ք�z��ޑ��ٹ��M�+�}��}�*�:�$���N�D��1�&�5����(�G�NT�S6s�^���b�rY��+^�9K� ���lOe3��ʸxH7"��Aڼ&N5��<�x����;7':j-�|;����l���c�]{��ͫ��N�.w<)N�Wu�c*��{L��z�t!<ͷyP�c"OU�"�8kB\+n�sH��R+�W]�2f��w�\8őЛ��ggh��GJ��T�Gw�]��@��z�o,��2��W
���$�h��<V��c!��xN;(�JEJ�؆�xB��K!PZ(��e�Yl�J��`�]�Đ�F�7KSL&�^Z�0H�T��r�U�oIVaÌ�&f��]�7޾E<��b,�6����G,���-�%\s+\j����,�m"�V�ڊ��m
5�[FѥZ�G��	��4s�gZ��H�ܜ�׽Y���ҧ/Wk�N���%u�	��{��#XmzKo�cɬ�J:_�پ1�d��0xڮj:(3t�����[�]��gC[�B�7=�,sƈ���mE�ݒ;�,n�G4���7{�\��3P��n�4z����+����QfP��1���ԮO�����x2���6-��J�l�K̦�*�x�'��.��r���T�	��V`�z�E���p\'4�E��4�u5�=1%]���L\\��W�jf8T���1��x�Q��z��S�;"&��}it���guY~L%�V�^�0�i۶�ɭ�Ib�{�ox�͜�S؆��b^�EM�EB���p��Շq�n�����e��s(?[A�sTY�};i�0Y��6�m0������O�bnfb�eKUQ�wg_���0L���s�xh*��21�Ą�
�^RwF�#�9��Ҽ�r��.�{2t�Ֆ+?QƎ[��9�e%�� q/)f8��>ԛ'���K�G��h���-��w=~�F��֏Z��O�=����efR������s�8�X_x"�7�m�-�b򕠷o��ܷ]�P\�o��{9�eS	���^��`�Ȗ݊3p<E����ҝ/Yn�P�g}ު�]ᯱK�1��}�gtм���!�ɯfc�Wƀ^���z��GWש�|�;j�Q�+S&:��� é��%��u!�� �ya�S��f�;w�X�����2�bט��+�xo��^2�DĒv����^?<�::
l�C#�%WG��,i�G�s���[Q�=Ҡ���e`���/ثZ۵�z3}�h��j"�'�W�K9�e$z���R����g)��W���p�e�����$���՗���;ۛ��Rc�f����j&���6d�Z�lc���]�V!5�t��E�k�����*Sr\�eB/�Gj�5t���e-��eaT���@/jՕ(*���P��q�V^qΥ�On�@��7.� ����c�˰cZ�t��N����HhN�un &A�<�;�Hŏ �I��B�.ʲNKV�R�li:$�b���Ti�p`f�JMջ4���F�<i��z���^n�Ǎ�՜nڤ� ��w��7��n�����dme��
E*+)b�TR��J-�mJ�V+H�Q�
�hڱ��q�#}�wM�3����-�m��%ye���t��뼡�sVd B�����ćp�	���������	�+,R����r�W�uk��JZpeӻ��{kZ�X�ό�6`�lR	�3^u�� �	��XtX�lm�H��sQ.?^�j��.] ��[�� �����rjmʡRn��e�6�����N&ʛ���[�^��Y:^v���8���g�߂
���ew��_�0{1X�tA't��fb�sT�H x'Y�[^'�@��/�/%�Z�B��JD;1淚ݵ+���~�22%��kQ�b6��Y��<�'so�}�A�V�]f��u�
�*ϑ�iH �րw���F�1dj�;�;���F[��:<6����IQc8Y�q�]������p�6�iL�yV>ǧ۷e�+��k�׮:�N�+h#���b]{Dt�5p�(���5k�I�L�S��t��,e��kՇ^55S�L��-f<�f"�f�v��\(=r����]�9P���{b���x	#K����YN�)$��\� �4$��Z��7����d|պ�޾�v���^������ ��<�^W��x����W��L�.�t���	K��g���b��_/Xư�0yՏ\�\V������Z�r�r}��rK����U�3�.N)i�����g�r�������`�����49�~7�f���׮�d�2���U��q��*[sU]B�I�a�K���&x�o���6߰w�9l���
��z����7Y�[�DS�e�E��4
1ah�n{{����˽K1E�].љ�U�{qU֣��WPUb)�w�0���2����*<F�ʬy_�iDо�O����R�6'��&;�^�j�$�����+���k���af�tS�0��W���:y,���\��y$��i���d�o�6q�S36uu�!��Ԕ�Ya�@-�WO.�o[3z2��μ��\�pP,2p���4#�KPܘ��L^m=�P�S��}}U��jF��MmZƢ�zDR���yh<"Ց,�v}.ѳ*輲��PMܻ� ���,�f�P@ �Vn�˺�\2Ey�鼱�^,ס=f�L[��9���7�<څ�YZU�����J�ZZԭ�-QT�Klm�DJ�Ҋ���2ҭa�O�5N��͞C5�О�f�8JH}B �Vh��շJ���ل�}�,���������H.9�[(/H�i��}f�C��^�}
QˢCP��ůoec���I�]�{N1���,����Ξ�%S�1��7���P���]�3`T�wC��5��8@$L��� ����9x�Q�'�v��y�V�*�^��l�{��9m;�d��t,%�ٶ�n՟*aZ��,<'U	hBlw*�Mu�Y�U�ZD�*r��b�����`H0=W��resǆh��?J�qk{�Y��mn��R�骺A"D|K㈸D�'嵷�fȄ��{�j��᡺
���+�&��F�g�8���}���g��w���N��3ϫ�I �>��0/f�;���/]�����c�Ŋ�N��J�ǑD��۳!=;��å��3 8�4c�8_5y�S�s��`���=��*YE�sNc¢���>6�b!�7(�P��Wb�׋�=vF����J�or�'b�Wl�̖ꦌ�N	E��е^|��w3��8�f�����LuD�䍢n�'��gM��*��I\�+'�uh�Z�V��V䳙��IIE��E��l���'rd2�)ق�	~��ǯK�Vc����:��X�VLau�Q�ju[b�R|k��7HFr�_����5��U�YyY���%�ب=���f�txE�Ҙ���Q����-���쉻��II�;vM�a^���-��˰=�����O~w͡�0��sܰGF绦+|����U��P�RF�6�û��N(�q9R]�Y�!Tҁ��%�1=�e�4ma=��;�:Yw��:��8�5�۽�t��t]We�Qn^;�PjT�+vq����~��nN�*���8�Q�Bz�G���F���,��t%�)\��u�T��£:koi0�T,fT�����T���Gf��(i���D[���D������Sk~Y�^Jޕ$���iQ���[�s��&b�Bc2��m���cav'Փx�nj����Q,��r�#p3�(����5�9C)r7�WECy\�s�3c��P&�A��J��r\�����-�;qrwwK�QYG-bO^cy����8s�m��Ħ.��k��{��4��im��*
��V-KiV�Dj��eA�TX���DQ�����$�5���S�vz79Rye� �{�^��&:|3��2ŝ Ӿ�͡�
�z��S�f\�x��x`C·-[�5�F⚌�.�N3�b�@uXb������k�m�((Zv�(GDy�if�c��K��1����j��ᛡP��3�D��밸�&���2����٨9�/�Z�h�7��<�ړ>�,��wu�>zs��Nl[�ywA&D�<=�͞�{�@9��N��X47zпD��x�'ƤB��0&�'"��W	��FvVGފV�Z����>����7%FGg{ʽ��J���Z<}�A����B����o��m�d�_E�� u4�`3;~5X#�ͪ����亂VR1�ݰ_���ЛQє�����y��Yw3\V���J�<����SpZL���\Mc;]�������"�$8v��M��n�lH��gMĽv*q��˸�HR��uc]K�,�D�ox��s��3����y$�}�/#��Ý�i��A�2<r�^�_�w���b��̮��Ǳ>,:�3������X0�.��Z�0�+��~+����w������yJ��'s����7:4_M���:��t��P!|n_4��w,�f�S�NɅb�Z��/��J]��.xt���ҡ���]#��d�����]���$�:N��=��_�׶���|����$uu��w����a��N�5���Z��v����0�|pT��\bp��|��q�/\f�v֌㙽P�Q�8��W䮲��#�P+;1�{�щ����h�����T�������E��fӣ��4��44�/˗I�M�6���e�?�+�v�"����j�6�h��~��H;F�b�G��٨��K���8��ۯӯ٪�_���J���������1��I$	 w�ag��$��5O���9le�e��<)�?��h��7�_!�`|Y I� I����o�dtPJi0?@v����ݳ�f���	�ܲ_����	H�/�!��W�Zﮚ����v�^��u
Se�Lذ��7X���9�C���L9�����;0?>7;��w�PT?4��:��ͻ�� @Z;�P��UP��bK3���rM�����PzSƄ��3��0��r(���7�
��w��}��p�"
���0Jof@U�ds��~�n����K��h-��o����!ٟ&"���3z*�YO����LT���^��t6pG���$��t@�:U�}D�S)[)���B��Q2�<,0:EAPŨ��¼�6��e��g�A��rXy�0�̳W��Y��=c#���8����F;�
��NvN�15�<ɕw��o�?i�,��Ms�� $���\�q+���"(�� �<7^S�E|�;3i��
��q]��h�>�4K�h�2 �RF��I�@��O�$�$���:���J�?	���6!�l��p�FBHI���b�ğ��0Z�����	$d�I��I�O�d���Ͼ�̭K�G�ϡ�9�l�-��7�^`P�)�$	��s�:��֛AP�;� x0$iz4�����>����h5��sI�q�1�Lw�`����n�"�;D:�I>�x����i$PT9�Nt�g��v$�I^=^��#Ȋ
��Ɓ^v.f}|SĿ<C�ˡ4�.`��:z�%h���Y���V &����;�N�+��z���;z�%�-o��˝ʈ��p�l(�vlH�R�aT���Б�ܳC��d[���q@�Y�(/>��T>��0jA�ϓ��۳vJ�nf�Ԑ1�m�!�J1VKqR���s�TȂ �y!z0�3m�w$S�	�j0�