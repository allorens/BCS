BZh91AY&SY����L߀`qg���#�*����b�H��IDUUT�S�                                   �((���  <                                    ��DJ��*�P�U	�)UT(�
*@�
 )EER�U�HAHU@ )"J�QJH�  ܩ�H�UR�P�I@S�}H��E7n�Ewc�Tn�*�)S:���
��PR���Gv(q�M;IV��,�`   ���  <}��q [���p w0� ���q:�c���z3x�I����9t��Z-�� q�w�    �@ {�B��UH(��s�+�= ��0{�� ��: 4�w��m�����y�A�l�������ǡ=8 7a�f�޳�   }� ��`v>����P��4@� ;��c��z
��)G���� dɠ��`�   ��B���DQR���P�%A>�}� G`�� -��� ���@������vzzRk<��,��ǰ��    ^��n����!����'m���� ;�p�w`����(m���d�� �Q�=���   �R � �B(T�P);��+m� 2p�vtDfIU���I8:GNA��wp{;��c�����v� [:��/{�    >}$  8�>�}��zLu n�td
m��ݎ���
"�)I`�9 ݺ@1��   �� �  �@PJ���� �֥U�� �q(7`��' Y�.��Wvp�9@�ä%٠Ϊ�g� 2    x�$ A�|��*����]��q�v@�#!���BK  ݇W ��Gπ (H$� � L��J��#  M4�� O�IJ��& &�F1&@ѡ�ʥ%?R@      �d��EDрM�� CFC	=RQ*� �     "DM=H�4�'�L����ڃCjlQ�_���>ϥV����>�Am�S}'{*o���_]{EUEp�� 
������ U�?��
����H������S�������=���j*���$�y�4����_�P{�A��"�������)�`��)�SŦ)LR�%0J`��)�S�٫�̮�]�]��-vZ��k��f�vj��k�k���1
`��)�P�i���	LR�%0J`4�)�S���S�)LR�%1`4�)�S1�	L��1Jb��vZ���k��ɖ�6�-vZ�����ٵ�k�n�)�S�	L�%1J`��#M	L�%1
b��)�S���ٮ�2�e��]��-vmvmvZ�ل۳k�k�V�0b��)�L�i�S�L��1J`4�i���)���	LR��1J`���+��j��k��en�]�ݕ�6�6�-vj��0Jb��)�S�)L��-��ݖ�&j�ٵ�k�k��en�]�]��5٦j쒘0b��i�S�)LB2��1J`��)�S�)L��e]��]��-vZ���k�Wf�f��L��٫�We�ʻ5vj��٫��,�]�e���Wf��]��5vZ�٫�k�rje�f�e��]�vZ��k�n�2�e��]��-vZ�ٵ�[��T�i�S�	LR�%1Jb�Čb��i�S�L��f�eBnͮ�n�n�ݕ�5�+vmvfUٵ�[��ejb4�i�S�$b��#L��0b��i�S�)�R��[�۳[��en��en�ݕ�5�+vV��[�n�1`4�)���#LR�3n#3+vmv[vV����[��f�Jf�e�enͮ�n�ݕ�6�*�mvV��L��0Z`��)��1b��J`��i�LR0F� ��LT`���"�q*�em3Un&�k�շ` �V����Q�*1�Kj�Jڻ5�-�vkV��
4�T� �1PjB1i��LAJb����LPb���*��T�
��A�(0)�)R#)�)LJb
SR���!R�"��D��0E)��LJ` �����f��m�ĭ�Ķ��D������0E)����[�Uĵi��vm�v 1Pi��LP`�� �ڶ�֪��[�����Lb�F�
4�E��ĵ��Z۲���n&�i�LZb��
S�)L�21J`4�i��������ٵ�[������)�S�)L�1J`���+vmvk��mvmvV��LR��1Jb��)���)�S�)LR��1
`��)��5	�k��f�e��]�����	L�$i�)�S�L���ң�]~#�nu���?M������ƒ�zB���,�m�7p5�tol��aK$��T��f�ZeQ�in�Y�!��Q���N�1��"�M�d�^㛣t����F��T�w�X�kͽU�|ۛclRvm账���72��(iԉ^ҍ�7BǢ��fћ�#yZV)��Ў���$�^,ɴ�+jY��yd��鸞h
%�@&G[��Z u1�Kvv�pR�@ۻ�.�A�݅5
l�1�2�Gn�IVV� h�!u5�4��o3�)L�/sj׶��[��"��,�Uə�U`F��K��v,�ph���X�D�!��G}y�ժى�h����v��TJ��a�����N^�a�)e�1���7��A�QKٚp��XLT��Xj��i�Y�%*W��.��:JCbf1J�̢��дk��~��(�=�Z�3t<7x�л�y�{(�f9j�ԠM`��<t6�3X�FܫW�V�F[��$�.���#t��0ƃw�R�o���)K&0k)�;���
5r�;�j�P�8��	�C�HR�[[�m�n�`�u�������R�ӣ����9���ͱ���Ed���'��F�*1l���n5X�a��6J�ڀ�n�d��º�(���;oBv.��@�k��z�Xf[�6xjX5�w=%f��Ƒ��!{,Sͷ,-�km̺��K6��{V�R�)W�25�w�x������ԥb�ơ��f� U��j�s,�1�X��h��Ȃc7okv�J��$�m�p���q���۽�j����捔6�� ܫ�*
�eJz.[�T-h�kF�Fi��\�BB>���*�Pe鎷-���ؓZ����2��f���)٧l�y�1�;�H*�mVSF"7t���&����T��qB�E<{����i�c.V�X3i��7��]]��N9�f��i��;$Ӵ2+�c[�mo0�nl/o��Բ�$:tBnf$Ҝ�j,��G��B�Ĳ�HՍ7�r��@൲�\��`)�R�&6�q��n�s()"���V"t�F�]��T$�:xcئZ�2�-]���݅;6���²�JLZU/R�l�{�4�`Ӈj�ۈ�%,�;�s
���p�g�IB�b��٦I�
Q�VD�ս5���AR��0۔�]��gt-�6Z�wyr��a��P�j���%^�Wr�����C/s2�I�eG�n�ı,��^�a�[��o5��{:�o[�X��4�2L�X�������ЖC��LYt �1�ر���ǃpo�(�ȭ5/%�ljV�^�+hA��{���+w|^��e<-�ՉN��'\�W��1�=����$)74�n
�ٺƥ(�Kn�!ћhG��ce�G{��Fjs��V�/�5=��2��=3t�&�q�;b��!ܸ#��H�2�6����Ė�E�]Jq&	��6x��!bB�ab�5YAm'{�5n<�4ި(d�Tb� ̬���{e�!yJZ����Bĳ���M-�[[ur��r�r;{�5P��`�� �{�uI���S+-l=ɷ(�+�����Oq��Gx��˭����&��e��N�`�w�x�7�Zݽ�����f��#vd��P�lᔱ��RF�"�u�kѕ{sfxE<����o-���V�9p0%J�ov�Dfe8S70Y�3�!�W�{�TэA��V��@mYӋ4` �6�ڸ2�*�(��;ͬ�V��0��w�6�%o�n���T�;�\�)b�6,dM������ -7x���!�.��Ė;��+]��5�^�K�G��k%<:r�^��g%���T6],��-d-�vO]R���@�F��`�Ӗ�;����[%�(6[� B��h��d�5D;r��Pw�ǚ�ۺ{��`ˢ\Ҏ"RZ��[�j�R"艅Էz�y�Q�sFb5 �ooo70�n�6����e�6�k��Ǝ\�Kچ$��J�*,��(�<0�~�8���C�zsp^ޜIʵY� ��%��^��f��;�E鼤N�J�fVeM�{DCu0��F�)'�6�
%I�WQ;x0�n�%gk-����2�5�v���z4d�I�+cp�1mb�5��n< m=���&�hw�(`��)=�֮<����K*�Z�9n�DU�ͺt��A��;��*�[Ȭ��Ǻp��i(Y[*L�T�t+��T�+���˂��#��uݢ��y��r�n�n��.����Ai��4��R�Qe
{gY��.���b]��%�Ҟd��V)n�]�C`\��e����tq��`�w�e�7�=tn�G`�vи&���.V��x���=.;MX�BG��V뼛�IBm�Knh�u��H�eD�mY�5&���n�ۥtv��[j�V�x��č=L3�"�b��"ɬ:�*�9n��,P9�KB�F˭1VaͶ�t6f���NiI+#Feٔ�dJn=�%eB�7.���$T�U��+F�p�jQ)z.��Ǻ`��^�C�i��/h�sP�Ұ�Snx��
��nj�Ѷi�ղ�I))�ӱ(�d�Ŷ^lD�,�L�H�֭��ˋu�U͇2�Y�a�Yd�	:����aZe^�0�b���f[��V��Ô��j�4c�I�����m�nmշ
�ܦ���U�6�!&���x��5j��ť��.�b���m�2n�-���X��x���`z�Ç��T��)~�בe書$;[�1*���K�f)��ūl��bΔD�b٠Y��/
�mPi���@�Bmf�We���|T�ΛO�IW+.�S�嘅<�3jZ�.��LN��-K!�tXŘk���	��=$^,�g! ֍�<h�M�v�n�����$ѫ\TC���ۙ���˞�Q�m���������cJAK�D��́�h��X��km��[-]k]n�\�-��L�x�mnkR��3+.���H�I"���V'6nm��! U��%�9u�	d�8I��a��Ź<�f�ʔ����f�y!��WP��Uh.�`�S̭'q:�ѵ�ۍ�Q̣	7z0��R9�F��m��������q��n#g4e\�4}�n���o��+S4�D����G�\Z*�^��,ݻ/bz����N�X��޵����Њ�����e]�8^�1�K�W�᭩��6��ڸo\�r��@�����S\7
��7�a�+F-n7"Vn�&�<�n�����ۆѳX-�R�̭�̅J٭���CБ\��KwzQ]Y��ŀ,���Up�j�itA�T��L��Z8SӔ�̆�Z�f��w,պN��h��F��oƐ;�yV��\j!�+K��ܩ�尲)�S����w�(Bƈ�J������J��ӬsM�EŐ�� \f��Z��@�	ړ����&�R�����c-�Z� ��n��f��3n3�I��a��F�������X�Z� Y�=��S�)h�
��z0���c%l���9��36�5[VM<Y�(*-M�n�
eO�xH�2��W���y[�]m=�
�0L�YYj��
ʩ53f�X�i`n/,˱����A���Y�V�T��r*��U�{�[Ķ6��v�eZj��z�˽aݼ�Q�f��S]�b����z[7l"�	x�^Ȳ��d�C���������-N�e��x2�����ڴM����e��c�2(Kv�-J{{��$����EZ����.����iq�������wf��J{�]N��>\��Q���8R�<�B�;�6�+/���ax�jT:�l���/F)[����[���J�\��V�7����J��k��1�"CF�-�̨�G�e
Ĭ���b-HVQ��o0�2w��iЫ9��d귗#g���иu^M���ټ�s�tv�2%*�J�kF�jku۔�3d�*�x�:̽N��Q�,քn�R/E�����i3���ݭ7Jx�1`�{Xe���m<��wZ,H�.fڡ6q��� 3�ū()��M~j��s�e�*���V�:��t+@-�gE��t�f`BS�Z	��A�ek///gXO,)�5���{X�3�qJ�Vn�nHʬ�޸��07���n��2�\ˌ�=ܐ]jh��70{��(bɤG@i�rTSr^Ƈ�s׷RDh!�Gp���9�� S�W"�S�i��,��l֍�-!v2�j�SH��b%+Cy��[�M$�%�l��V��`�е<e�nJ��v��{��4����e�iH���2:&+����329��`yG�ùv��G� [6�+R�H�̫�2]]��T��T7F��Cl��+P�ғy�V]���^�{u��]�K �
h�[t�#��i����ފ�ܧE���m�c����" hbA^Ia�mlƍ]9G4m����	�( 3p�{�El�a"��T&a�+F� K�,� 5�0��k�p�l��Z��	CVci�O
�̬`k�L��L�h��C�oZY�f+J�f򡻤�[u)*��*Ɇ��f-F�j�T��%�x�d���nف�MƀW�(��n��gNi��Ԓ�Ze�MX�y�J�y{Kv�3]z�:���b��+V�ÇƜܭÐ����� ��^�,ޙ@+���9J͜$kQTB�b���t��:۵yg�PB;x����O\W��@�b�tց�v�D�Ps.n=T����"s��v3a�wKX�vh���i�O��EWl%�P�4�����	����H%�ˆ+�]nݱ��{L]a���lVJ�JTcQ9��
�Z0�w������7dԋtEF^�V����\,������c��nXg�۫j���ne��[5�pT�d�I2(��X�(n� ъ�#"���& �T۽�C`�NT� �#Ic,��Vַ���Y)�6X*�Ƕ� �CwI��j�c[b�0�b�e�d^�P��ͭ�ͻ݃�8,dz8�x��f�d�dh���'C��r��/m��Vp�K�[M�����`,�2��]�$X�������Y��^�� hWJ���w�kv�e�ҭ�v�O	[�!#fj�,�+p��i�aё2qᱵhօ0�J��H�!@b��n��B��4��^Ûi-Tv�R4L�6�a�ڊ+�B�Å�
�b:Rf�z\�lx���}yu|���[��������4���m(j^D�@�ʳB�ܓ2F9��۶����t��#pk�	��͓��ݘ���X�u��&[-Ȃl^md�V��B�ѹ6�GV���B�rI���K��f�*
97p�P�o6���PR��n�����ֳu�r�<�f�'I�h'(v�ݨ�r�l�c��0[Qa>�U�R�36�"
>��
8(&c�2�֊�:�5����^�`ugȮ��=�N�JCB�K%���[3t[���̾&�k�^[\�G�3x}�E�4<ӰI@�]h���yU��
�f���J�y�5�.���v޸�mi��KS�3C 6�EX�`�4={�ف�I8̽u��F�d�)^8�h���Q�ZD�zĦ�c2������#K��6�sw��t�������(��ņ��J��jy�
7Vh�Pj:�t�t��\����. Z��4^,��0@���,������pI)ŭ$\�YyH�C�q�il�j��s,��v.�S�QT˫$1���*��c�Xڻ�/����zJ��v�7��E�Dͱy�����bs]�5�l=7��幃.�nc6�T����%���������&����Z�i�RPyY��RTYLE�At�9j�ǂ�Lv0��u��)�X:v�񫡶�0'�*C�RTV�f��+u���!Q�oJ7D�#(^_�6��U�'Y�F�+r��73��N'v�̃
C�n���$n�^a��kL�w���"u��0�h5�%c�a�4�D58�,%J�$Xy�{`6�%��Ԥ�сkMڸ�<��YY[kL��]�C#��4��[a_�U�x졙p��!Q�8.�+�.:Bi�$�#�2=ByN��2��4�J����{C���˭��RƷ#�Z�:�:�n���l☴i�������V�i��fjyz��e]-8�[xN`!��EP���Y�w�/m�J� :jI�XASoF��Ϋ:2�s7/ssh�)M�� ׯ+(Y���M�BmH�ŇLe�1����5�v��t*fҴ��J��6˚<]F��@45Y��׬^V�,��-��If�V��ͥ6[��tVeK�v�ڱ�ѷl`wrX ��^���0�3f�ٹy{��\�c;�i����yVKu�6��YOJ�{$v�RO�(q4&�����l�'	�)@PK%�5r�6]��������|/	Zl�d�:N��r�%��:ز�p�d�$�.���7���]���8N�K�Y�%���&c�wrbD��JaN�9��L'�D�hf�v]�iճP����Ǹ�'S��#
�a49������m���c7gQ0�7Yc���a(� ���4.�0�J���^Bx�d���d���$����IDL�yd�t�9���~�>M������-Z�c{>c���	n�D%�{(T��k���MxT6�d�k.�,��d�:J �|^s?e�a&�4'��J<���LX$�:J*��-(o�I6L$���p�'	D�z+�W)�a$�{�B�&�3y�x�J�6͒(
ɠ8�&C�e^a0��-����0�)e�`�>_��<O��y��J�U�Fَ9�ss% IDB�(�#J�h
1��J&�Ý�,YT$�	�	�u�F�CeYݐH$��gM�~;��K�,�aMea?�ݬ�h�]N�mf�x���p�*�$���<��}�-M���Ѓ-� x Kp�o	�ٶ��|{I'��t�'�d-�80�d�G�^B0�I6���%����ZM�#ǍM��0�Qd�F_@� ���K0�<<�� �wb��h��1�.��=�ַ@i,�&���+�D��sG4�7@�n=�{��� |0�=��~�bR�%$���OJ)����C���w��~A���������֔G�Pd@��lV��Fڢ�X�X���j�kZ6ڨ�ѭX�Q���V�V�գm�ű�����Z�jƭQ����Q�Q�kmQm��-����֫kXլUF�Q��X�KkE��Ʊ[h��*�b�UF�m����XգV�Z�Q�cm�V*��UUj5m�j�ŵE��m�j��Z���6��ֱ��F�h�-�X��m���Q�5Z-�X��Q����j-��E�bբ�Ջ[H�""��(���9O�q�=ǝR�*���֨w��s�9[/V�@���+�-V行L僓���"%BAy]j �n)�)����|���
��uh��t����B�D���@wqC}��{����u�ܗC��j�.dFj����ʭE;�\�L�؝��	+
���$@모�ý݋W�b]�搻���D"�Q����"�����?���|~P���'�?���,�AG���������3�����>l��ϧ��U+�����znw2�Yk*����xs��n`����Z����6`�V�09@����xKR���t�\�s��u^escb�T�[�W��A)1h����U��vz�U��ʯ4bem�`��i��T��w��mc�<�Lם��1�Y�hZP���5}v��[hWս�z89W��ʮ#n�"_��ڽ���ֺ�^j�958���շ��Lh�L�Ώmm��2��P�zx�p�z��/�y�O_^���"�:�B��n�r���mݡ�W{�����8Lq��^������F�څhY�Ͷ�Z6��9��Gn���t��/b,� )5�EרN���l�J����I#�Go^ݔ�z�� �ie����Ŝ�}��ے�y�v��f]�4:[��S��՘�qf���������u��P�*���������g����m
D�m���hӺ�fZL�*�(9�B�@�T,���W���K��(�p�[��/K�<�N��V��S�7lc��%��U�{t���ܭ�d�)B����;X�L�*VGn4ê��x�aݫښ,.=�U��z�\��l\2�v��3n��2�v�M�^�l�����(enr�}f�9`����k뺊ҲL��UT��`�OwX�ǄS�{�ufWR�)�z�t�b�Z��&d����n�zx��qӎ8㎜q�v�8ێ8�=8�8�8�pq�qǎ8��q�q�8�N8�8�8��8�8�یq�q�x�8�8�<qƜq�qǧq�q�8�8��i�q�x��8�8�8ێ8�;q�t�4�m��8�N8�8��q��q�q��q���:q�q�n8㎜q�t�8�q�v�8߻���{���w������+�[��<5�jݙ�Ո�h���2��:�ĳ	V޶n�k+�v�ϣn���ܭ���bGt�5��t���T��Z��
F���{Zʅ.����E#�P�����^�jm�c��ޯ3wetR�+d��8�E[�����������;��Y�5)R������^U�wN�ҧ�@髭�:�<+{�0q��mӻ�48&<��Ӛɶ���c8�8���d��?`�b�\��R��큮�!�0�����x��_<�O��V�	��ס�z�6�u͵�Z����8�M�g.�G4k�YO�o�`�`�h�4k��'1�=�ʕ�TWf�*Et�)��";5w*���U�,�GLh$�v�W&��	ЮR�Ԓ��Oʱ�S_,��}�D��;W�<���$�2F�To,!�i:Uv{��:A��r�>��#g�1�t5����N�:�pٛ:�m��ʑU��e��U}���	n�YT�u���wr���U�u��in�
�jFs�tL�o�K����ky4�V�.�	��X֍݄�i1Q"�ѤU���M+.���\�pJ�6Ԡ��s3yW/����b4��e\�Vr�{WpcZA�[��
�b�,"e�-��2`��09�z�Ч�������S+Y�o�۴m���oX��,��tRy3�ƽ<����w��pq�q�q��8�8�<qƜq�qǧq�q�v�8��q�q�zq�m�q��q�q�qǧq�q�q�84�8�<q�8�8�=�8�8�8��q�qǧq�q��q�q���8�8���8�m��q�q�qǎ8ӎ8�8�88�8�8ノ8�8�88�8�8ノ8�8�88�8�{̬쳹W��yM�4P�����nrǉxY;ڲ���y���Zw�t�}r�J��a�����#����4m L��sз���x�:�嬼 k&'��JV6��� iu�S *!�!������;(;A�gh�.lJ��۞�'u��L	,VB��MWv�ΜT-#��y��ޯl��{�5�dݺ���w�Wx��q�������k�����Ĩp�szi��t�n���ɝ6�T^b�q��- ��n�c���;�Y�u�ݕ��[�s9�[0!,5�_V�2*4�����4�x��k0�۽�@�#�z��|�	��3�\\���8������El�.��\Uە�����iX\[7����s`���]�wU�u]�,LQ���ͩ�)t��$�m��Uf�ԩ*��h�-S��-5�pǵ������<� �rεG�u�`��b�M#����UA�h�y�-����tފ��E,�S��d���(Y�ϒ��(wv�9:�U(����������&W87��J0�Z�XEJ�wsYoC�4.���Vv�VR찜z^�,Y�!
1���;f������+�9����5)�i ����6R�] �\��q�#�j��ub2�ÙZ	D����Wv���z�	{�Q��s4tP��mz|�ry9�J� ��6�{�CY|6��pqB��G�q`�m>#2�&Cx,�0��F����n��f��c|s�RŘ�9i����G�V��Nه��\��u�3k���]fl����y��4�uB�t���s(V�˺�0N��A]1wK�ѝH���"�1�'�'���+Z7�3�op!u5%'ۂI�)�wW<�t\�Zch�j��`���Y�HۡU��9vI(����`sW��޹]�Qɯk3j��&{$w�2�r�j���N��a�ӝGi��I�!��;1�Јm�m�n�5n�uc\��Sp�|+�
!\ δ�u�yr�ڼ�qh�2K�]ɉ�^�u�ݰ�Ha����/{v��E�q���]�j��s<7�JfcG:�YJ�zFk���V2�l��s	t��`Af�쭽�ZY4���Z:ṚhQ�Yi���6���v�4���V�/\t��%���xE���`7�����3o3���#�i�e[�
U����/c��D̬������\�3��.\�-b!�Y������,߷#b�U((�b��8�MЩ�9�ޮ��dK�mMٖM�(^,O���wϦ��;%N��T�[ĄN��l(�sHg#�����ٸ��Zk�i���[��B[�^֥r��=�"��d�:�lm�i�R1�}���b<Ҭ.Ej�K��zFR^$������
�����:�_c��"+U�X�a�|��oGB�y[
��vu�v��Us1��g��.���@�MCe֫ۡC9�z�Y��wI�l���<d�[b��}����XqlLt�ۙZS͙�OZ}�/|;m�/�_R��y<cd}�tZ�+��-�f���J㘡�+�����&TV�pW��c7E��ٱ�֊��9]�Qn��]�ib����<X{_�fq�8n+�;���v.���1�1�>b�r0��[rJ6r�m��P
˔�yACmy�镕y��{�s�7�c1f���ϏV�� ����Ojty)MX2�;��N����ݓ��p�i3���/k��/oM�����aWY��r�],j��m�=hq�D���k@�e���tS��v�I�`�a�Ge��uSrmY��E����+��ݪ}�(���N�(jp\��yƬM��+��S˔g�*��G���f����Ш������*O5��f���dü���L���Ωq.ކ�b�+���cMY=wyW�ŷ�R�٦��U�*Z��7�З�Fֺ����RV����4��ّE۲k�n���=�z�����ޜ7&�C1u��¥�%�WD�y��]�eog!wܖ��� �D�9x��f���lgLz�t���f[�7af�=��"!�{����!�������nSqY��U���5��/<���S�pf�1�*b@Ƒ��9�я6�2�W<&���f��wu�Zǫ��J�;����V�yE�V䩨�L|�T낻(vo]�Y�.���q)��</�7X�ŭѧ֓�=�BY�Ar+�] }G�Y���n�#�|��x4��'X-z!;�ٷ�ʚ��7��YЋ{*�8M�T���u4�r�K����h˷�Z�W�m�3��׆���E7� ��+/fK��atO��lv�sU��8WU���7�ZݽXXܷ��杉�Z�_`�!�N�uha�d�#�&Yk�h�u�K紳{S`j��Tw�y���U�OE�������|#[ʺ��N�j�Z	�0v\�rƘY���o���5�9OW�L����9�/b{�;.\{[V�������ܸB��8�9�GFծ;��y�����m�LW�zFٚ����cO8���7+=�������J�U�r
�i���0���w�;��kE>:0� ���Q&���[��Wm�z76��=݂x��75E[�բ;]��Y�۶:��u�8�%����x�ʲ)Y=��Q�.��]�O�z�,u
��c������2���ף7d�V�)���M�rT�˫TMc{'mǽFV�=N;��+wP�m
�l�t����(fF�P4a#R�3�ӂ�X��N�O)e!�`�`����+�r��g��V_�|�SO�VЮ�4v�o]�컬���WmX�'wf�l��yv�hn^���0��)�\U'w�g9�^=�>��}-��uף+x� f2��ږ��6�V��:��EYv���<�f���y`r�`�w\Ϋ��:���\���kШV�u��zб8E�S�0H��5�L`��zZ)�۩f��_	g]�G=�s�����y:��*ƞ�;|5��t�Nq�I��0�R�9vU卵ZhP�&��������fqd��o[q�O�H�a�z���h�]�p:�a�*��"��9)��w�ݕ����P�Xx�<��Q��4��<W9�-ǡ;��V�ͽӮn�)�Yn�Xytw�t6�����y�̒�U�t�����m��]�Y�)���+6�fs�Z�yJ�̥�[�s�tj�ջ-����,�:����R�K<���2L*�Aw��<�i̚X��SpcW�\f{+���,լ��=��\��Y�{ޜY��ԇ�EOY��d��g9mOo;v��b aН�g5;��m�n�.­���␑��s+��ɔ��FC�tV��-ٲ��2�%EV��|��ع�hw �r�s'�@�]��I�ݥd����ڗ\��30�}��TN7Yn���'a��uHwkC��f��X��B0�}������s�<�9W�!��Wh�ɺ򠹧LV�.���M��_1c)ƈ��Ӓ�g�/Ӥ�rz��x���*"SoC��%�S���·x��VMc]�{���.����خD�[�:z��>]�K/ h��GPu���+��r�.5�T���vZ��a[GF�Br��s;]�fVe]���r�:\�t/��7�mtrh3Tj�5�fHq���0;P��� fQ �ն�CI��{�=[������T��=�(*�c�+@̫�ɋvA���죁Jl�9�����:�{�����oo4�?'���5W���C��N��V����d�{�s�$��b�L �ŋ��\��6�u�{�³�W�����s�]b�uOE������Z��ѓ��{v^:}pb켰����Y���T5���;+��\,�	�[�W;iNyaԾ��D�]��A�����7L����R��O�v����k��Y��
'��VF�l�+h��ܮ�]OJ/�Mה�w:f]}LvX�XĎ�|}[��Y�\yʷ�T\l�;�"��!J��zԤ^�~B7��y�^���koM�u���s@+]��fx�F���)��98�b=���;�C�og�J�sH��\9%/��e�MMu����Kܞ̼����xU�]f��!��ڒ��������A�p#c�x&A9n K�i�X*���\��G�h�Y:X΍e��b��F�7oT�����`s�t����b���6�	���w�sjѴ]���~a���IX���lG��Q��*�\��Aõ�|gw+���<R�s#�X������;g_�Jbv:�Pl�����Ւ�v�搾+�4oD�����V7h��'�3�Zg�z�K�;�>R�}g��ʋk�����[U>���`�*����{,��E����t��ԴM�.���W4��wu�g4���x��=w~�h2m
,����݂N��;���w���3a��Mi��yJ�ՕrX|� z��<�ԝ|�൒o1V�ˁ^�	�|n�ye^����ǶҲ!��益�hWM��"#w�<�ם�]�f�t;xV˼��VA6���Y\�j��԰�:ϫёAةD�R��g�'|�H��3VY׉Պ�rV�ڥi�s�p\@�E����Ȓ�w��/B��2��)fw<���e�\��z.X֊t�7�+��9��2�"���r�����`zl0��sMl�]:MbQS�wsj�W
fT���]�n��Va<l��cZ��S,(v�r�xh�=Zwķ�ך��+j�����k�������f��V*ڸb�ݪ���q/�mu�Xi\�8r��=��Q�'�1@��i��x�^gCI+�충�<��{�^z�e���ٙ���2u`�8ĩ�VQ��4,��ܢ��^ms��ү0p�+�u�zJ���l^t�egq$�٣���3c�S�3���}��`�!��[06UP�ާsX5wU���k2���ۨ�9ӝC��շ����`i�J����ҭmh��}����y��*.�R�ȯU���
�m�}�p���{Lll��B0H)-'�1Ǫ�x�:��ͼ�-۪�gc�v�U��K�sqR̲ x�9���v+�p��I{��.[�t�Y�x�����iX�޻����ޮs�e�X2������j�\L�˃��e�ԢC�.N�q5s��N}b��=T��b)�3w�K-\�<C`���!^;�|sU��!ͦsn«�5o�;�nޮ�����V�W��]G��΢�t����ǔ�a���bۧ�<�i��e� �v��J�{���|�u^��\�;�r,�9�F��z���W�;imL��QӜ7PC<{�xH�ָL�����O{���ɞ��b��@V\*�b�ꄞ^�O�EU�����~ϯ����_�����_��W��n���"v�'侧�B.��V��)a���|+#(P�`�T�tM��.�y,&t<�&��r\ùPȋ�xC6���|}��N��˃2���˓J>ڔ5�΅�а����îYn�����k�	�lB��b=���X�n�JS�_<��U�� �B1�[�*����osm�֫��`�xŮ�+�+!b���V��ýA�Kaףv��K���c�����8�ݽ���tN�a�w�O��j����]�ݤ9��,�l�q����Џ��on�^�p≣kr�O5	5��x����p$��=n�,i�h)%���")�]F5LkI���kGe�`n1�����r��Ǜ�6�1�
P;%���4�ݣ���A��)��.7k�8��x<�&#J�iHquq)11,n(���X,q��e
�(^�bw/0Vf���]q�����D֓m� k��n�e�c�U�^�!*ѹ��nvy\\떳ԗ%�c���k��gM�,��}v�M����F-m�V����[-�JX�5����`����9-�����o1\vY�:ɹ;d�v�����.]S�8r�l2�-wb���YT�X6�ه[���b�0oD-Yvy��T:�#�[4�ש�m-���On��mۜpcSF1vNPrC��.5��i�qP0)tl�M�!�kj�IHh�����b�idfՋ1�0��ɗo
����^ .�+��]�:{�����l`�li+�0 �����Tq�m�u�F	���ݮ6�î޶w.�n��]uŎ�VW:ـS��=��p�s&�z��h�ݴ
{n��t�t^�zzv9�i�㑜���㮺�+��uAqta�ָ6;T�k g^�^��5#z���'�	T�%�u����%�s���*C]���8L��uz��YFA��1��	ap�'�8���,5#���Ua�0�1�a�Bѓi�q���I�8V[.�H�6�LJ%�r9���F\�\H���N9�x�����~��"x����@�5��z툻1�N��y�B�u6�uE�n�UT�q7�f颎�7'eͮ��*�Ffm,c4��bu�فZŁ.��@Vx7lo&Ɣ�tkbq[�\&���۟<6���9�*�a1�Q� jI��N$p%��ѻl�&�)f��۪܊Tc��u���~l}ƶy6����-����v'5U�/�ɃC�6��ȕ���݋��6〗N����0��7gpR�����u� ���+j�\�Кl�%�ִXm��v.&)�h�`Kc,�x,��\�U��:7��oh��۷��=1�x��;�8�u�n7]�Uɶm���1 ����[���SN��*�Sۈ�sv�v��Y�+���S��N����:W�D�Met��qd�se�r.����ל��r�gY�)�n����v���h�d����K��q��N�͸�N��:�Ҟ�ćT9���]��5{-R��`�[��Ym9 �V��n�1l�Zg���lt�l7]firK*�@q��LFŘ�%�\�e�)��@]���u��竞��܀r��y�o|�@&��,,�k��))��y�<�͞JY��T��%�]a�Գaږ�^��H�K��X�w�V��X{]�/;:��r-i)�&�sX;�)�=��M���g����g�[�!��P4�,��f0�޸�յ٭�{��qs�S���r�ј�I���ㅏ^xƺ:ǬÎ}�B;u��X��2rgz�>�K�m6F&S���zާ%�rk�C����;��s��kf�*������;s��/�j��;y��R��cp۞e�]�a0�hJ���W�]���v9k���
[,[��f�"�s��� �M�E;McaHY]uNԵ��n'�|'�N�eL	������n��6�l��i1l�p��Y;�H�"�^ܧm�b�ݬd�8\5���X,X����-�ڶ�x�ni�7"	u��^��nx��Gq�v�f�	��]�V`����,���,���66�����ll�V���3guOA�s�7����2���Zc�q.�X�FgL�1���&����t=����3^�&�{Bv��N4[o9�B����d���ݢ�Ņ����G��|����-)нZ�s���t�I���ͺ�#�����w�ﯵ���;�D�^&2d��������b ��m&�y8-K��n�G�5��4�yW⪊a]@͠�5�v����1<�¸>��#�^ێ�.3:%5]`��W������N��:��.�o4�]3�ϋ�ѻR2�v��1�����s��f���m�%p]1T�̚5���q`�:,<c�5�ȹܽu��ps�eO :y�;,:��]�E��e�5��,4MLDt�:f��鮊��GV�BZ1��³5����<�&�qY�7%ōt*J�ޘk��30-�K���"�G�����3m),�+0	i���0�5��5�i�5��<p��ˢ����679n����+�SB�Fc��*��Ua-k4�e��g#����۝5y�؁㰆��g�6�,\.bK0@���,
Zi�V.ׇW�n�X��%\65�����S]�FN�G$㳪vx
IC-ušh��ց��{$č�s��5���k'��0�x�n.4Ȯ�]��y��r������P�%���BW\�����c=��Ct[�BS�vs=��]f\�tc�R���[Lc)�8J����7g��kN^����Ѻa�p58qqɱY`f�J�H+6�Yv��Xʚf���n��^Ӎ�1 �llg@�8fV`�3X��t��0��Nv��n��Cn�5�׮���p��6�q\g4��G�Mâ��d�^�����쳫1�!]�l��K	��� �κ��l�q�`ǲ���8]6ɵK/lHBT-٬j�@�hl�]��N�U9�-x8���q�Ók�vc����vÈ��m��r=�Z��˼�����j�b��6��ܨ�k���f��׍n`��a[�e�,R�IL�b��U���� �L�3^ĻXQ�l�ւ��.�R��lx��3��M++	��)!n��h�LCi^}\Ü��.�5�l���B�2¶�@Y�����GLF��<�ʼa���lk���A�������r�v�Fx�9S���k'\un7Ǝ��Q6<��؜/<��#�pv��VƸ�{��롍��:�l���1B������'��lMI\�]1kX2�-W�G�m9/Z��EB��f�֭���	��|Bdk��j�Q����I�A��R8�u�����i2C
Glkq�AKL<lFٮ�����Z�a2l��v)�lhw]t����q;�\l�8�^ĸ7=�I���H�H�^�T�3Q�6[lL�KF��Ӵ\C�pc�`�#[�̱��l��I�撩�붘�W:��'	���'7Of���� q'9�Y�M狮����a}^�;As&|-�92+��un�	r�=Fѐi�������#�{�ۢ��Jl�c2ʴc���	�mu����ƕ��r��â���`6��O
�'Y�`�,uM���۲$�aF4I��u�q��GB�:F-�i&r�Z��SS�n&��FS,6�,���zS������a���-r�c=P;�Ơf[l 2�m ؖ����L܊v��n�|�u���c��=a,���[���vy5�W���M�ě]��c�#c^��Pg�.K�v] J�GG�e�]q/��v����`݇`��W����{��gQك�֭�^1Ơڭ͛!�u'=�5e�������O�h/3q�q��63�/�9
�[t��/l�Ƃ���vK���V�ԗ�:���p6��kZ�'d����7�Ks�4�%���88�I�3�HͲ��׃���w���.<�xۮ��mH���0��1p�[�b�i�H�t��[���@�v#��#�+�y���^`�{}|�n�K���<l��v�gR糶BB�#�VmY�sI��pg�&4t�tK6ô���
l�:&t)�^�lv���U�6OGol�:9�6�c���d�7foc�so-�Aŧ���4s�����^�����y�Sp�ch�%�^6�y�k�:��T���FblP�:�uյ�iep����9'�B<��{�j���q#�*��K-l�0:n�K6�,mm���n�y���vw�ZL콙�эF�� �`�Bx�(�j�
q
J��證A`b�b6�<�K)LۅxB�/6�ڎ�d�Ů:��m&:�<����7��]�g�E�C���}���0.��kYL�f	M-�&�kˬ!-�T���e���<hWh};;�}�}ٮ�u��n�����@h�&i$�� �����t�&pY�lչMp������J��(HOE�x.{�$nz�KT;�F�
ܗ�˵˶�N���t�v�X3螹�B;3
�.����4T�VɵѰ�1�i
�e��ջs���u�d����mt4�*��i�Yu��jjB��ڮn6�Bn�(��c�cjn*mr*5lt1��V�4`GM��ں�6v�q�x�:�pOV㞩�dͮϊ0t�����ްݳNnngi��Y�j��p�UF�kf����9�s\f�=vj���j����Z����훲���ܴ�UU{'d��ޛGm�}���n���k�'����9��Vx�ٴ�9%BK�]_ۈ���ˍYu:��-������.�c���E,�5�C-����˟��Ԃ�k)���.`�J�*5B��њ�f9uI1�u��؟98;LlD&֬�֙��a�Pi�O;�ҔI �ttx�Q�g���qIIe�uYRDq��N5�{,��v���$�-��4��b��������A�!����͊�t���\�7����w�x���.�.vPL�=q�Q�m����j�6��i}z%B@�S�s��8��m eX3K�E��-�X�1��}��o��J(2=�޾�QJf&����BH��H0 �1��<~��8ノ8�;v�۷n8���KR1��B��b7�]E�&#~ҺF�����P3=�
ZV杻zzq�pq�q�nݻv�����}s`�������B14�m$��(�D�>v��ݮL��ݹ�D�{�%I]6wZ�,b�0�݈�k�21��u�E!_�,�/wb��uE���d�cEF�L�e��/��D�\5��B�4_U�F���W�)5��ެ�,0�5����m͙_�����ӝ�޺�9Tl,c��m_��!��#�p���r�r4��w1�_�t�7e{��t�9�����ݷo��/:�ss��纍e����o�%wp���k���d��f�b�5�A����ߟ;�:�gv�˫��]wn��r�����R��a(Ci��mN��W-����^B���'6��ws��7,�v��ws������l��Փ����G���L�
�&�n�v��UQ�!�w��{U��Ok3���bسtC0�4�@�w�u�P
��mp�=K����Y��Q�Q�Q�5(͊�]�],%t3��km#��Bƶ[8��B*%����n3�p���nY�=�s�e���F<DݍvWgmD1��3�и����t{^u٘�p:Wh�P�Kf�	��:�b�3o0�u�Vx�8-�i�E.&2k���F�v��s�$]\��\q�e�V��*���Ң�k.�Y��d�ƃ���,H���n}N��c^�����+��Jӈ�^�-c��- ]��4v�َ�!��ff�7�h׳��t�ݗ�����x�גݬj)ūM۵Mn�X�@��&!F�/1��W�cdxJ�N�8ֺ-����`u���O���{��M� �v�����.܋�Ah�Ր�^��D�%�,�v��l�Ɖ��լ$Fi�Q�z���7M���g��m)0iX �8��ifn�b8�����:��eڝ:Ŝ<�4$���Yl%�1[��
.�R5�g�[�=����^�A���{P�;V+n�Tr˃ՀV̤nZ�4P@]c�v�����7��T�㶢�Ga�*L��Vˋ���vݤ�s�k�nGɖi4ؙ6�7:h*� X�`͵�G��Y���BX��8���nTd��{[v�:�`�f�b'Ld-̗\#v	�.a���n]϶� M���؞��Z5��B[=���Jv��r�WrֻUQ��v�+.v�A�Q�ep7ذof�h��`X��`�n$����lR�F�d��#�8���^�� nU���θ��=������m� p��N\є��ItFb�P�5էƈ-�8�d���J�&���Z�[5SL�R��A�$cvK1f��GSYLZ�9bZ��B�D!,FJths���5��GY�Sa��]��Yk'�{��;��^�{m�_�=�=�e�+���E��P[z�P��h
�¥�-�D���j[R�HԂ�B���+�+e����qeiఔK)^�ZD�J����,���V�G�a������8��l
!!X6b-��t�o)eHW�Ж[jZ25%mX�T��+F�E0�9t$Q�U�d�:�F�nf�8s3��T.X��n]ˮi+���?����׭(xSf����np�[%��\�,�K�:�}>^�k��6|��U����t��M��M���Ɖ���˥�M&��*�����gg٦���l��|�m�߻o\N���&��܇��Z�}
�f&ScU<���5��ŀ���l��P/w[��jsE
������0T>�̔����|�����U$�@��һ������Tƌ�}N��M��iخ}+�;&2M`4B�9wl;W�9�Q�Z��4"G���-�L��y�߿aw��a8�[^UUP�н��ñ����J����z/�V��@L�2�˷����&Ѯ����D�݆�KGV�sQڻ9�.�n9pi���l҈|�d��of#�k1�T�k�	/�4�*_}K���,X��� ���}�=^���ڜ��Қ����ƃ�]}���W�T��>���x�fЌمa V�/��Qz"�޲�ư�Lŷ\�Be[CU@��ţΟ�;7�[Ul&-2�M`w��Ό��E��>�����E̔t�f�4٦��z�a�Iy����DZW�C�6<~ۼ�~���ڜ��R�� V*��M�Kj˓�w�����jҰ��[X�Ѹ8rt�G;��u	'7:t���m�+��8�SUS�Q�L���Z��/��=����Y��J�T�m���o�6���z�5Z9nӹ��7V>�x�v||}�����)����xt>l�f����/sL��a|'?���J{%�ʽ1uE|�]*b��T��Bj�G&L��S���[}t���T��pUA8��Ƚ�@����b�T
)���_}�z���~����N>l�&�5�����ۡ��^�[5�L��}J�l�ꩦ���V~�t>����6���'����\U>�)�^/�#t�laOW���WB٣��sqo={þI���_>���KͲ��v��q3B:��qx�f�f�2v��q �Ｐ�4�~T٠��څ�M?Wb]ݿY�����ﳻ}`PCi�y(<i�M���j�U�#�n_13�u��(L��O�5�q5W�kU��{q���R`�M��2����0|�>��Ԧ���}xS��0��2��V�N�/�ݨ��0��}�P�͡�=uq�|�3/D�����m���9*]���8�/��̱�1�m�'P;0 �H�*<�+�Q>�rŦ�G#ė�ו��A�j��^���;�b��������e33d���ߧ�捧A�Ϯr�4=%U�T���HU &|�jܟJb]`A=&0�x��l�OX"���'mڃv,0k��l���&)XO>������2�#�����{e�}'�|��a�����k�YW]���`�y�p�b�fN?�ѸC�]�z^!3�/;~����٨L�2��D��KѶ��_�Lr���&t�-ϻM6j�n�>��)�d�ۂ�5	�2�\`���[3�,;���ȿ�a��C^�[5M痙4�����w��v)�O���s7�.�[�{�
���ES��uL�����6�M�b׵g�Uy�λnΞ�\2��&fp�o��c�;Y��W�d'�5]��F�F=8�4ral^���
��Ur������ŋ^`Ufܙ��@�aӕ���U�׷�CQ��0b4��f�T���{M�-v�kt/gtۆ�.jL;f$�[�T�[q��mt/n��Q��s���O5����"�[9OD�����`���u�1�Wi`L-I�m�{Z�o4�X�.Z���G��yܩ���o7]u�͡l�&�e�c*��,R�n�.��n"ͪ���;��;����}��������A��b������%0.t�g�T8)�ӸP}�s���Θ��T �(�^����Pe]T2���j�.<�V����/ן�	f��#�f�eo�_��n�t�jq;ʻ��@\���9y�7#���_�ں�wG��u����f�sY{��c��q}��4٦ו6v�/>"�x��/͚ŤE�r߾��g=�@�����w���_Y���>���-�����_���0?���s���{�꧆�ж|�uY��}{L�r�E�Jѳh��Jm��[p̫`�%Fа\.�3fT��ÿ���ǽ}��wz�oh^T��\^�9�.���T,����yKYM�M�T᪐#S,�B�I�E�����h����uvL7�os�2���+��"7fU��8�lVd�=����	�*
,�&S�U���㶟@A���r|1��.+���(\�̋���^̟n��o��h�F���X�^6�f����0��}�
.�ϗ�\Θ9(w~����-���3)��a @8��}��3%ot�w�>���>�닱ǻ�y�gծ�K�5^�jC^�6�y4ۈ����i)����L^���D���t�ՠ\,�M��&L��Q+��3	�D�eQVc�=u4z�v��tu���\nn]0�q�B�Ґ0F����k5\���o��<�`��1O�Ѩ���t�A �[L�b L�UxUU@}��gЉ��9x�N>��u�Ӎ۹�X̻�X��A�BgD>E�˳��(V�����m�l]�}��3p��A��XQK`���� �*#R�kN�Yӗ�_v-�ܵkNuM�s��Co�t�Qy�V{[��-j���`(�9�K�Oj�2}톪�۾S='�[���fr�)6�6�� =+X��3]ݻ��٨/�WV��	�8W0N|�����ka�˿����^o/xBW��wz����ww��� O3(
U�X��h
ɊE)��-��=�m�{qǓ� ��Q��
�kt\���'խQ�8;3(e��\k�B�z��mع	�a��a�ʐw.en��v�.2��F���a�p7�f&�b�wֶvj�C�kD!��D��n�l�x��Y�F�ggv�y���b-��b͐)��O~Ac���vw�gަ�6o)+�7sZ`�e��
�.N��/|�вޮ�u��v���������%2�N򺼬��r�H\��U�/���r�D��Ӟ��H:0�����x�H�e��w�Z�.���R�dB+,'G��Ŝ���	�2�ꪑk��gm��xU�'f���z�h���0�#�*�6qJCb��bE!s z�6�oe3�=�^v��/l�.��˒:gM3���}��� L�|B`=(L��ʼ&��9��}�u؆�ShM�(Khy�n���]Tn��\0�7뽽����]�h�A1jl)�f+��q���zп&����٦����g^<(|<MK���}��B1�����f��^M�S�٬i�D��9�o̪Z}M�����gS���z���^q��u���g�$�H���z,�l�%�Iyݺ���Q�WhUn��e�T�d}�E_e���딳7zzvA_6����G�0���I�y����姺;;뭟1_V� ����h�/O� ����]������RL!pb��߼.ㅋ��<��#��o����"�ۣC��%��v鰤��&�	�@F��Bk���i��$���P��-�j��,%(b�`A��2��u������^�n�v}�ۍ�z�=cqD\pm�]�� <��1���
K�ʚ��⣞&B���mM�1*�X@�4�X��e��+���ۊv��m\m�����&���7�6�wK%%Fee'�����X|�d[]��6���ƚ��9Y�l�1��愕�0�^<a3i��a2��V����#3�\��v��-v�w��8i�٪^n���J���5�f'c���kۃV	�>7��'ɳ/yuR){cqfP;���30h1�O=��������D���<��4M�>�}]����M����`��H�%�4�ǱKv�d���)�s�0��\�Wq�ϩ�^>n�y�֩��\x]�Q�vX��&�3Z؊���.�����=��}���J�-��X�T�n��w���Z���kT�	Q��oY�?����-����ߎ������w��S�3��]��M��@Uk�j�5_c�=�p��[5�8:�G8�0V��^.�����K,�ϡ�ޯ���LN�f+�Cg"cwWJ��[��tW�1��bŋVdh(�"�~c�Ys�[���#���~ש���M��W�R3]���]����6��;DM�f��&��v�UI�.�Ɉ:J��&뇶����}M��>o4}����{a0��MTr϶�כ5Wt �t�;/=׽W��w�O��Ζ��0�e�T�L��S��
�sj�!�wO����)]
�4��.���sa��Vm�ڃ��'�g�o�F 'P�A�̡r�ά��D���%_+}���Nu�ݯ
o�ohw�W}��=#
v�>o4}Z&�`����i��sw�^���7z���Qa����R���`�0o������ |�jG҃ż�Z^�oj��s��$�W�-`.�iڽ��H۫��.�x]Զ��ʴ+v�u�t�g[ �Ǚ�i�}�ެ;���܋#��ܙ�mW2��-I��V��g.�MS��HBO�_gw���ɍ%-�%����2���2]�;C���rL,�"z�uк����3��:�`�L�U�;W��>f��v�]��뗼��DⷋM��gB"��vJ[��Sz�̨��a,�˓+
*�o^YX���z�����y�r�T�5��{�uȺ�������󷆝[�U�͹`��Ԛp^ͧ��wԸ�͐ɽ��ԫΗ�r�ōQxq2��U��E`��]Դ��c���
�*�{��G�Q������V�[ˡƷz�����*Y#W9�/������]AC�8�N��Tbp�s�����k�s��ѿ2��՝�j�Iݾ�I<���3ϼ0��n���jZ'�_�y;ls+pO��m��Ϯ���߯���wA�:�j�AQ�5��n;^�*l�y]���.���KE2�R�����VM9K"��d<�i� ���Loa����+�'1y��j
�R-�> #3Q�U �^�ۉ�OL����fT������+�b�+5ߝ+=��W���7GU�D�n�M躖�_[/l��ݔt��X�
�N��T���]`wM�,�C�0�'�٠��ijO���DXH;�p3�(
܋�D���,f
 H�"`枌 �}��z߬P�S6̥c����BD tAʼX�z�7W�#w6�_p������Ä�$)Z	�ѻ�q�b�s��ݺ~{��g[�.n�M����ӢQ�*\�?�K�4���]��HKKB����1��P�m��㷧�o��>���8�ӧN�qƞ�'�����!�QcB�ӄU�lW7wnm��Q�wv���.T;�s�ƣL(�C�1�O���o���>>1����ۧN�>>>=�L�T�U##Lnd���m�f��wr�ƍ��\wj]�_źP�����+��DcEs]5��b/*���F$(�]������W��bh���s|oM���c����P|r�E��7��yPk�*�b�c!�{����mdT_V�`#\9i�sTlb��5�nb�$U��PY���v�h��u��]*���su�͢�ۉ|\#�U�*-����h+W�������r�M�b,W��������;]�z��~�nݻ-�3�3gӾ�yUPu�#��������ÑT��3��S�C���n>:#��gB��p�
TE�qd�٬�&�wX̧,=3^l��<����;���A[��4��H8 �j.��9:��Z��{����
�8NM��z}G����M�L�,�-� ,.�Y�6���z��'y>~��K�ke��Lcf{�q�@�'6��)l"6�B	�sM��XU���lRS�A��9��Ǹlo�;yJ������[�w�7�y!,GJƎ��Nj��0Ʃ �����6;3�x4� �E1oy6����KkWz��zH��ݸ���' �'u5H	��C
Yl�1k��8��
�A7 ����q�ef�Hj}E�zr�z�}G��Ce�8$f&v�vERg�7]�l��#�l�T)[�kCy��5���j��p��y��)�7kp�ˠ���� =�/�j~��Q8>����z�-���A7m��e�v�̬����˯�Ϟ��8����Ύ�VW����������3��)��!8%���&M��7Є�/��b��b�P��2h.�;*��!�7��l�@����T��<g�d��<t� �e9 F�����������.�,��2jqq��uR�,�,�nA�Z�Ε&1m���=w��,����^��2ʤ��*���W=��3�<�w|/�zsn㣢FF ��L:��� � �Rr=�My�=�hu�f� �,�d;������V�ʩ��Ӝ���B
b�\8"��$WT=37���� �����U8p����XƬ���f���~���d<�ɗ�F�F���M�wd�A�Rp@��+�}W������,�X��U�e�O�G5��6_8$f �&����@<&�n��=2�/I�(A�K3}����4l� &*��v�%�ռ�W8]�4�a�i�������^A[�Q����3�\ ���5�����s`ڻǩlP��s%��r������]��㕶��>��	M���jF@�HX�ƼJ79���2i�w_���B7�?��ƴö�Jg;V�3��Տb��k��yڎ�e�#�e�����'���Z:q�뗱�6�c�� �S��IPe,���9�;���:;x��5F����qul�W��Zp1%��l�z�3�	Վ�:�vZ��z��!a9VKd|�m��Z� �}�W][[�$�j;t��X�e���au�l���7KX�.�]e�Ij���2Py�q��+	i����)YVi��qj����%���u<v� �9H9a��;U�pES�5RmQ̸yݓ/�n. �$��'{��8̹�S_&�2�@Ak���#*����~kR�a)؍�`���ޟT�n�Vs8$e�d&܆�ER�^F�+�0�*�p{�9�A��/1JA� 4#�\#�T��e)SwY���##Z�1(�g�v� ^T��
�p��3������ ��:-�������L��;f�eD��~o71p S�Jc�h��7�l݈h>�f�^-T�U!�*�1�*��������4.p�*���g��&���e��A�n8�)y؉�*s�Ѳ��#?P�Ѻ&�"�).��j��䤶��́�v��	qr�����7Y��D@�$�A��Q�N���s�V��z��C�^��#�;�×��ȱ��vi�� �T�6Ņ�jb"�8!�z\��^7���_Ģ�YP��AR2y�6C�AX`�=��򻎾�*�ڒ����;�hx#rd��׃��hSky�&LCbC��H=���{�͕��F�1R����Bݢ��ETn�F�	3��M��kT�U/1e�0��#�����v�}Q�л�l�pH�NXCn8��wbRT�:2�<2�QܫR5�59�Pr�pU,]nw�:��S��׼ᦓ6����v�ex��4"KS�q���aE�r�p������p�?�4E:�cz��T.o71q��hucv��T���޴m�����A�ː]�
�4�M�3]\��Hj�s��%��֛5K�y�}}�|�F^�]�E�v ��`�E�V�t���W|8ޖvq�^�} �,X�,�Zhcv�]�	�NEn��<eų:@ܝ�'�;zý��މOT9�y�>��z��5��\�XF�X ��W����S(n�Z!���b-Y�ȫ��=}h�j4uQB�R���˨_�aW�>�W�Z;�=���WU��x�'Cu�aְ(�0�md����!���)	����&L���̃KM�X^/*_�𣙹��A1H#N��3�$*�Av]�F򧙶���������$.p�M��]�{�sk�=ޮqhU�P,&�G�3��*����CC=� B�O#�W<�\ t��$r�oq����$@�'��k��:�)��
;�4�q�M��e�ۋ�Y*T}����������m��6�:�.�B�ek"���bMXa0H ��s�d�O?�$�~�?q�E���5"f��EfJ��l��L����k��c4�X )� է�Lm;uxС!�+��>�Ü������:ipAn`�ͻ�u{�Zw������d ����U]U�ݻg=G:���xe|�D2�,�[���dSB�NA�V�)�²,��t9�6�B)9$'���S��H�N� X̠��/\9�D3�8r*��7y#O�)zm�ZV`X{�8"��v4��kɭ���j#�͙�f.>�)x�L'�CH�9_~�V�s
�kAz���������h���=<ޗ�g��K>���|�4���-�%+�հ
��z��ם�z��D��I���=�m���m�%&C�}U�������H8�Â*_�xV��H��A���w���84j������Eۻj��e.�Qt�$y�/��A+W5ac�s乌i���n�k��Xٍ�.�w�*ZA|����q��A7i��N�p���Ps���8	�Vw�u,�m���u8v#�8 �T��aT���B�A�s^Q~���6��a ��v'ma��ȿz�tLOI}m�����=j�
�n���Mx�u����[�Zo�8'�
U"��9B�$>��^&.���ok�@G�^�dvױ��WZל�-9n8^p��!�nԑ�'4b�}辠 �iH5�t���N ��Xws�Tp������޺��_^5��}�1:�l:�r�pU-h-wgN�����N0m�(E�]��=:*g����p ��A���j�K@T�g����M�b�˃�u<`��;_	I`e�X�X���S@Rڵ��ەts��c�����wG����q��ءm�؀�fy�L�wf��%1��x��v��vz,j�3v;�z-��d�"벯.x��z7i��E����5t1cMc�-FSt��D�4),���v�;n15�-��ST�
�ut�1O�ڌ9�*����5�'m�b�49aLR�.����-taKf5��H9�aIq�^��tvC-^v�ݗ���$t�
�D����Q~���XVg����S��H0�$`T<�Bı��`�KaXR�v`őkƘ2fʻsGS�e]���e��+cAmw`�
�yö
����F��6b�޺̿=�� �X6��aE&v5H9�R�Rv#*z�\[�f�C� � ݧa�\s���p����׼����w8"�V{.������;|Ֆ�ѕad�z�"C��6Q�Yl�H8�&_Ͻ��H�ʎ!ʍ��T�OQ{��q�' �������NZ��-A�[F{Ϗ���R��P T���l�&:�؃ѫ�x�pX���X��F��v���KX�:郰0Ū�My\��n�1i���R�#��R�ĩ�\2�[�A�l��C�7\9i�`n�n�]r	B^�a��"��M �&`m�c�Wmt�5�%�6��Lm��li]���Y�}� �����@)��h7i����_W�h����k��qi��լ�t�a���>b��@E �HSc;FfW��4f�=�-�-�4¯��>����d�BTt����Q��G
u��}�]�ǯ�����Cb���ү��CɑV]o�O������[m��D
��+���e�|o画���]ke�pAa���7;TZnT?z��M��'(ח�����P��p������u�;����M��}%�� ��NS� ��g��&��{�(�f	�<�m��� U �3�~��mמz���š��ńP�y��Ȋf�BRg1lc�Ð � ������>g�#������3�v����g+�/�� 6\w8,*�b)Q�=u1�N%�F�5���k)t�+M���Qi� Z2v@�ц6M֤���A�R�)kK-�cyi��k��^;��������9����_����+��Q� o-�d�s���$���g����[w��CAN�	#V�3�^��mמz��ܥ��L3��Hj���ѩ���������>p�v�pA�p�h�gj�aqZ2yV��H^�f�+//ʷ{Q"�;`���}A�]�f#�u�y�z��}bu ��$x)zie���#qb�V�^)� ���A��mA�۾땝k��}�^��ke��,6[q3]۵#Xݩ,<��/���ɧ[Ϥ@�Ln׶�o�wus��K��y�fS"�6M7N����fM��B9�r쓓�ȓ�R�Rp����qfo���0R����o�����)qy����`�8-T���c���f���\D'I�.��I!��KGm�Vmч��f��m�%���]����_;�~>=-��
b�k�ERalb���j��v���Ʋ���Ƶ���r��+���aR�u� An���h ���nPm5��
�k�pkS��b�U�׽ޮE���8Q���b��p0�bz������� �"u�8,X]�"*���̸bn�1���^$k�Tx�U�M{^m��7)q���A�R��'ɮ�����U;��1�a0�Gbl��偪p��w���ޜc��Ah�Ń�ս}��O�����vA��R촆o,,�n���W�\e�rd驀�m��Y\U�fA�K5�te�o�:����Pëz��V�{D�Ӷ�@��l@U����2��Zm{�,��Yr���Qd�}�Z�Oy���א�WOq����2�<9�y�5H9`{�
��S����}�:��=��l-��B\lS%��޵xܖ�Kw����s hA��|�і����ǥ��c���Ue��lº��M��Ek�s>f�U�5�	�Z��&�9i�-��a �[U{�b�m!�\��LV�����Vt��7�����`FZ���Qy~9���6��L�'b3S��(��y?&ݯNf�-��-�	9X�#:縗��9���e ���"� ��4�؊Ba!I;R��(�q6�8r6�g5H8靪���y��"�vR�7���26���|�p�mX,�W��R`���R!�#0[��+��m�!ö��r=����o+�/�2�Ł�p���v,j��S/ ~��wx���E��ZrIf�hnD�]��.�dƁ��)�յ�ff�4�h5�b��9�����co[`��M�̩{i�R���G��� �����֍v���Yʳl@6�\������r	�x�&pČ��A�EK�X��s�BI�3��8��������u�#�]n�e�Yd�ʷ�����+E´�]zc���>Z]���Sv �ϭ t�im;���ގ��_ٷ����)��YH��.�T�6A3�Du.l��W^�/bcS��[���ɸ���YvΫ��*:��ol�`��s%ٛ|tv�l�b��嚎vN5%��@8�b��V�+jWuK̎�S�՗o�h�eM0�nȝ˚ɹ��������Gb֭[�尥��wR�tn�d�*_+C��& �T���}�
�����:�d�ڧ֘�B�[��}���a��v2��=؃�t{/2�������1R[-f�M�y�(&�;L�㓸ۥ[g��lk�.g��UۥVs6��c�$��oZK����^�pfJ5���v�݃gl�b��e8��×]T;�3�����ٌ�-Aǯi�SpT�}��`ܱ�t�����ڵJoq|O���Kgr���gWn oU�C��uh`<����U}o�j[`�t1f�w(��#�p�Z�9-}�2�A�*�˄H��2��R\7&��^�C��\�����c����Y�2��j#�D5�na��Avx�WKZ�o��.���B�G�~�ʟ��V���l��ID���Ƙ���E_����]Q�Y\6	�J�rT�M4㷷�oo�q�8���ӷn�>>><�P%E	��J�(����@�i���qǎ8�q�ǧnݻ|������_W)��Z�yҠ�c��d5�w�sV"��܂-�]БR�6`�dưFH�F����j"��\���Qb��U���I��.���[na(�m�E?Z�ۥ��J *M`6�j�QF���(œE�E�}۵rh�cb�[r4cF2Xڢ6/�%���X�}6�[�36�y���*/-vWƹ�rۄe��8�O?�^�Z�'X����SR�zwn��|u�}�2��f8��N1�r����69z���f�%md����pX��ѣ�����6aˍ��3K����y�PL�im����bBU���V9#�iP�,ͺ-m��x�0I�4ʉ]a�G�V��l�I/l��e�[�H,�Q�,Lİ��oZ���Y�LS���z�f��u�ݳ!cTp��#�v��viG{a�͈��\��L"C�iu�nŭ] �ѸrkA��B���h�'`�b#q���x9�s�98ظ�t�1����l�*,, �%�gD̻�v0��nƒ�6�M\\�tKOIS�����'>������=�(A�S��xsD�)�L-BͶ@їH����әK,�Ҷ�-�s�]&[c���n��H�;s�˛[���v%j:�,b4�km5��X��m���Ta�5��RO$�]�f�N��p��Ʋ��g�TM�sP�v݋��2�M�I�I�C�4���G�����M�`ڮ=�x/#Ѧu]�����3��a�Ҙ��� ��v6�x����C`��:�m�k���*\�v�h�.�yN��&0�ڛC"V�.5�������<�` �x����4��.23Z
�2�Uѵee�8"�b1ѻ&���K���nl.癹�lp��0�Mu�Wm��!�ܕ�c%��ԈkkP�|n8��;I�<�v�����1q����+[E��SGOs�t
�p�3e�\�5t�z��h�^��^^/6�q��j)s���Z%5��j$D����|Vft�Q㇞����:{4a{<wnӑq$��#�k�qLn���ϭ� 7g�����/^Q��{a�8�mMrl�T��`��f�t
K��C4.[J�ٺ"%��<<�m#��Fn�lk �1�{5���8�n�͌7N;��m�&��U5Uq%�Ik�h��iL�~d���w4f��C�7�:�W+xm1{L��(ҩ�I�n͇�Ć<��r��֊�j�∱��bm6��  �*Վ��w�*�	F
81��MR�3�B�8�7n^����u��3�("�Čԇ���"T�2�pY-�D�@�����kF�E&m��n���I���bcv�5��c0D�la0\.$f��2�e�����/m@������af�ZVh^�bc��2�",k�-k]�
���'g��-֡�lf�PĳiLm���{����>y3%x�y��W�����Ճ��6n���M:�t�n�w��u��5e0�6$��z���2Yz��l����ǈ��;>���������LW���sf�8��ԲV�z�h �s�#�;�ñN��j�eW��FZ�{)�H"]Æ')ɜ�ݝW1���v��-���'ucT��5�,?< s�(-�򞼣q#�Yd9ʲ$y���W�Bӝ7>S�ϧ�ݛ�p���Aa��	i؃����w� �',2�
]2g�;TA�[(A�@;���qw�U�����D��nl�pA�L�ًΘ�5�����@"y9� !��Z�AȪNX�p���G���[t���uVt��-�;>g� ���8c��۴^�:4'��ٴTL�mrd"N�{�$���Z�G�&�m�# %.�6sf�m��;g;(;j	��`Ah4���1��8}�yZ�|����E:�w�����*B�R��yC��!B��58fv���%~�K�|�8�����B�ebׇRY*�3�K��7.����Q�Ig�89�c�Bx�Y�]���.���$�<����K����WWd;���G�UƟm�m��*�A�y�=��*�B{����_׵��|}k�����s�b.�Z��n"�ك�]�\V�v ���5P�My0�u��4��=�~�6���B�l�n;)�'u0sT��H
��2�b�6�;����S���Q���|>�y\�|�Zv,/|ilTe�����y��p�A�A��9�Rs�@ݠ�k;���|bf@�X�O]����|=54��9�m�CM�A��L�i�ZΛ�y��s�~��u��G�R��5@S�Z�t#�\���s�D<A (ocNr�H�A�A�A�gv�gm��ӈZ�)p#��X��ĭf.����L���J�̙T��`�Gf��g,��a0�ǐ�+��6Ы�ڏf�������/��m�<�UU����v��T����������RpA`j�3�=�ޅ��hW����nGt�/sa�z�\�:e;�����f
9��=�IL���z�`��NF��s�������mm��U`��/o�xg�ji�����M>@|6�8"�z�1�^c�R����%��>���R2gv�gm�8���/Pn%Qg�%L�mH6 �R��p���&P�������,l8��θ���_��V�F_zb2�n�<In�MR�s~�ؓ����ڋ��p`C%\D�Ɗn�F�=�ru�wPã�/d����y������������!j�� U%T;g7z�����V��7�����N=6k�,�Y��X ��`�FrpER�0�JZc3E���l�<E�g,L�`�3�׻V��8���z�Ac�����T��7A���fzM8��S�"� �An+��f�a�{��nls�^���@] 9�6۱�[1c`�L�]��z��f�"}�����咃T/�IU��]�y7�{}j�Ì�"r�j<=�%�*��ٹCE[����a�̮�  {�gnv��,�3��7�;w:��������u��nR�=�FA驻�����>�ؠ�m�

A�U�=��(}e �w��N�>j�`Z[����s�R���A�+3:�%GN!k8���rS�Ac������A���Ї��9�06��9�	��&�A: ��s��Mz��䎌rfb2ȇ��IɄ�D�w��Hi�L�7�8"�8>b�����k����^�͕�z�^��-F�)�w�>,;ɼX���1xMRpXePJ���I��J���j��[�8z�yC7�fz�oO��P�y�\�ERg}κ��A��"��r#u �"�Â*�ؚ�/cD�zРŧ#��+��{=�Z�id�a�C��X�{����=2:v�Mv��y#mL����������S�:��/w��b�̮�X�pAi�/��+�a�~�uT��8ʕ�y��	9�c�cf��?�)���x��ߨfо�|�_��sN��į1k�vh�lEږ3o�����6��n��<���2�qW��ߟw��a �;��8�M� X�����X7/ȿ�φ|���&Nu�=�=ݞ*�6�mm��QD'F��+�����}ٽ�MJ�X�i�h�S5�-�]���tQ�z�$[T��ظ2�����R;mN��Q9u�\(a���h��ɺ�%��=���v�����lbon���s�^GM��-
���z�@wZgì�7>��90�윮�+w)I�A�"�MY[��c7EY�4�P��ruƓ�v���Z����A�@ٻ�wn�U�gT�K�HZ������e�ck�,Y����+c��/���� �'1��XUh�6�o�k���ye��,���ê�{'r���؅�ܵ�(�r9��J'�v��<�K@Z靁�@U&��㷩�q��h@>8\�\�Ugt=���^�͵Ŝ#�˂7SUJ����l"�2�A��jr�-T��]拋�2:C'�:f���=~�Q�N���=i�T�4���C\�9͖�Y�Y��닶�&�C}Yd9�c9\��fz�tV��F8����K&�PXw�ݗ/���;O&���p>���58"�:`MCHP�R����~���3}�~VUg�R��؁��Z����8l�v�T��F��xq��z��N�%=%�st՜ȶㇵ[����nF���ÞjK�'�މߤ�}G,-T�XK&T��h��ow>d_��p���x������f<�����d4���H}HA��X!!�}� ��/.����Q�0�$s���r
�Q�"�gM6�1]duv�v�e�����;��7�Z	���H�};S&R�#�ẻ�[)zyA�iJ(vh����2�|�h��J��`���2���|ã9�w�[�~�]>>�Qm��QdUX;��e�'�Y����
ٯ�1Ŭ��A%9t��`�P��uћ�������8�zY��N��.	���{޲r�J$��u��#�.ty��3�!�uÑT��F�pRa,hG	����1�s7r��d;��CU'g��;��./�j8I�M>A�2a���>����B����k�,*�Ѣ��p�V%��vN�zٱ��RD���Ίɾx��k�(3���*��j�"�Ll�vp4Q'APIw���4A��=��]t@��ё�6Q.�Un����`�;h҃�Ǳ�E���Cvg'���~���pF�
�T��L�Xa�J΀E���&v��D8�
��k��!T���=����bָ��9x�;Ȯ}��zȿI��Gy�O�v �r�8.���\�}�y���i){k�P,�N���h�r��'���������68r�!Ds�'b޹��0ZkW��7�p��u��bZ�3�,_Su{�y�Y=����mU��l���=;}<*��x��@�_7)�^�� ��&�9�fݠ87u�;(i�׵�a
x��o
��0�f;Un������:���1��=7�R�����[N�nԂ	�PҘzՐ���W^�i��bH1�ü�׽�笋�Ҏt8�Ƀ��1�.AN=�Z;9�/tw�����Y��/簣���6��l�m	���.m�VF �5��)�f��'Ƌ;�N=�g�������|�-f�.b.���+$�3_&s$�sS��Rv"�:� ���4}������lh�8t�jX�9��w�g�n�[i�|��UU��L� ��� Ƨ �;Iو"���' �T�t��<J~��j@��"�'w^�/�j5�y��@8�p������NY0���<(��/�ُ@L��#ɞ���U �&�6�l�>yžub�-���N���o��Y,e]�����S��xrV�f����&�<�=5ө,Y� *���L0�F+�Z�0��D�]e�N�]�{D4�l-��@���rs�(���V��� ���&Th�8�ݞ�}a�l�q�r�V�ށ��W<�\��n��"�ݨ��7^\��Y�ua�蛵�@��DC��JOl��w�i�dK�V�x�[��b1<�_G���z7���c^N&�;��̎��Y�(�-=���vj3P�Aj��.A�p�U;��E�1)�L�yϬ6����㦪�:��o�%žvZncr��#V��^ۇ~�>�  Y�NG��ݩbԓQ���N1�g|���G��3�x���Nzz���Z�#u"�ñ���T���<w#��b�f���MΈs����N�U�oq츸�QɌ���{�8�G?d�-K�^P�Ё��]Ɛ��P�AN������$�v�`��e��MS�vJ��k��' �ZC����S%n����x��,P?J'���o��[n�w��S4����P�vui匤zc�U,G���M�O<�f�:�U��3;�W/v�T{|}6��m��;O��s�n�2QP�"�'P�w�d��-��6P^h����cL�,������6��5٦�Q�������v�ݝIf�nu�%�	�n��F��c��M�MkJ�b��6�c h1�ic�Mca
�K6�V�S�Zg�s��-B˳��Wt7��tc���j�p�F�#h�7X�w\E=�줹�7w	�����ƃ8Km�W��ؖ>ے9�G9�^�n�)9N���UQ��<������<�0[i� �;Q��A�qTsz����/A��m���zȚxW@i�@����`�E*!�R��'b��|:��E���kRUegwq�Ȩ�Q�4����AǙ��hȹ�[�>
�İ�p3�pm�j���D[�TF](�ݨ��s�r��wpA>y��~�{���B�vZ�A7��A��hT�S��Mv�/H���^�Wz�G�Ã4��dۇ�s�gV�@�o|�i���#Z��J�7�z٣mڵ3�����j��j�����*�v]�^�&);�jW�û1�}P�N'n|�9�9ÃT��*��|�����/�p���5tn�
	 �+��A�L뉒�0�LGM	�	x�d�)�!9x��e7�C@B�W�ک7Md�d�ɵ�hS��c޽��l�Bl�g�R�x��R�) on�[�[��G{��U>�"���έ�K�"��?)Aer}����8��k3/�wF�lһ�x>�c0�%t]���l���*ܦ*Zߙ�VC`����Jt�m��lTSZ�:��a\��
Ͼ��v�}m�o��Z1C5��s��T��eL�@�vwe��w�<���2+�r#�yh�;/L~�9��s�-��sO�,�t5���PV�؊�<u��څ�v\9��ES���Uǳ�M�]�O�X��yq�`�[����Uh����N�N�T�� ��7h!�7kز)`������9���[��#W8'-f�- !N�Ʃ���O�f��_�u�lԙ4˅����#�s��K����E���˃�}w�_��/�{�ǘj�K��J߆��c߽0�N.��]�v$�� ���4�0T�Uy�T���<Q|Z�6�
ؗ�zE�\�����WV�>p��k��A���O36�KSd�jd-'oT��� �T��5A��8W��x��������v�4we	G/��}j��V��cu��Tok%n��ǊY���W�[qU!,��M[ө�ЁB�*�6�5��4�T}H,���!
xC��/"m�ZoM��tWS�w�k6r��}��۽����h���6�ɋ0s ��N���RhK�D��jn
>W4_RR�ţWvs�a�Q)4��[G٫���*
��G�ɢ����*���kJb����K�z��:S����b��S��Rx����ӊ�jYVo�]�X���Fg,��Ρ��r
��+�]�0�����B�cj�,Q:Y=�������4�9o�u��WQo3Lk`�u�^oRӕ�*�
�Xe��j]3���x��лzQ2�̒�M����5]����+S��f�]���5�J�Zw\
f���]�ϔ�i��{k=�=�����7�kF*�E�����[.u��Uu����<��X�L3&�B��{6�J�\�K�}z�[�I=AQML X��Z��7�T٪���f��LTҀʝq;���ue5�!�⬺9-N��:��jsTH핋�5{�����I5����]�6.�E-�u�Ik�ʥ�u�`ō��c�޻��{I�1V�"c�w(sI�՜Y��5}�n˲�W����/FH:���We�mu؞����(���n֕��fty81��m=�E��+;9�hݸ��u刎=���k�����W��cTإI��גi�6k��	hx�\��tDw�w�"ٗ��o+�j�$ A � �d��c��+y[��j�C��v����������i�v���۷����UͪK1%]ݣFۅE�Ӎ��ǎ8��4�;|zv������$$	�
�#R�X�gwe��n&߯���s��va�����o6ߝ�4X�~v�Fэ���m{��jI��}[�k�R�5R����
��Uw���F1��j@�[�\G�W-��v���a(�5�ߊ�S4���ZH�1��ڂ��;֋�W-����b��Ph�[�S�YD������m�D���N{u�\�_6���-#5"���NɌRm���q������ m�`E1���k��oofT{����SB���`�O{�@?k��l��� ݠ��V�؊���qS8wvv���nj���TVt�ncr��7]��A�&�O���9}�iX�
�@1R�٣G2�J�J�	G,s��HkM�v�î��O�χ}?��O8��p�ߐv �8v�ם@�+Wͷ�&�=;��G@ؔr�8#-݈N�Rp)�LU ���WV�ǢM3�2�5i����b�{1�ޘ\&�1�y1C9Ú�*H��̹ç��-�)&B*��SC B�ERgN�^���"#�~N�8H>�O�W*z��)gN.-r����j�&p���5JA�E�}4�se@�9�9LnІ�כ@��\��6�8'-"h�X6�����4tI�(��YX�&�YвWl�ٶ�%��ʚ��%�u���w��]]�^'�n��8�J��f�3|�^��>�P-��Dfe�y7õ�̮�X�r�p*�ȩ�ȿ`p})��ߣ~��W�	��A1��5��0�v��ۋ�K6�^]S�[$��rv^&��r�Ԁ�.�]a[`�ѸD@P��Vs�8 �:b��]��v��#�W�ô���%gN.i@�K�{�s�a����' �T�T��� v{X�9��h��u#��7�@��\�_6���h9�@�E��.�����+_���) �֜nݜ�媕{(�rg|-^��
�Y�7'ojj;_��xC��A�4h�) ���ё�x�}��B�mR�/C*�X�vw���"Vy��A�9;#m*bmEvYv��Z�9i� � ������<���8�5�~�Nѭ�	�5�<2������FbrS�U��A�Bx�~�s�DKy�rɬ�A�e�YC�Q~h�O�q�B|�wy�0w��c���]}F�ϰ�Wu�l���r�s��Ĺ���[*��㏶�m��AdQC�;�d���O=S����%akI�)p�f����Ϻ�q�l�\�hF��p��=͡q�Ñ�����4���Gn�NC�D���eB�<]��P��0j�G��Tu�\�s[�x6���=�[��l��2��#�[n�6]A׶Y�*��ֈݶܼ٫��lٝ�z�����۞�O�ycŝ����ss7&�B=&z��\�=,�Wv6f�41��PU��#(8.6������y���͇q�q�6-=w;͎qC�sŎG���:��K�A7��@�z���K�Nl�f������a���ǣO:G��Р�@M�*�r*��X�"�8!��Ub�ӀE��o�{�;W����w�坔�A�NA5Ko*��P�x����'A=���p��A����^hd*����]g���VU�z���/�o��#-3��qR//
BB��=�ċ�0{>K�_}	�X�����Rv~�Zc��U=�?4�8 ��;�O�ݻ=��zJ��L��[!w�<Fbrl.���k���cәGCW ��:����}~�o,���r٩���,j������������W���v[�a���t\uզhv+�=��AxF�X�Hc���@�p�T��*�>���r��HK�_6�8�MRucg}����]cSU؍�ذ9����,j�� 7v�w���PxuQ;��~&�1W&�Lh�{���W|;�<�f1���|��K�x&�2�ky�=4k(��1�*t<�0hh+޿g��T;;;8f2� [����q�~�v�����ܨ�����y ���U*F}�<�K�끙���:�pAj�ERg����8ؿE˛n�3�ۤ{������\r�w]��Rp �&�^ ����~�^筝�Y��"*�8ɳyp^�F�[*�ڈ�:F�r���j602��n�h��p ݮb.�j��^�zŗ��O�kUwI��Q�)sA��s�N��C�Z�����<Vϳͼ��m�hh�nb�n��$R(p��T���ϋ7m��Ad�)�[|	�@8�p�U;��v�^��J:�\я�+��Q��_���4w��1��x���I� ��Aȥ�Ef�r�[���V�v���p^�I\�/���C@LkQ��Fg�����l�X�?��*��/���B�FP��p�I��������n�ѵۺ���`�YwS]�ӡB�ZK����wk��vq!n�f�Aҳ2�v�&P8�+ޫing����� +m`��=�8�J8e "�T��U8r*��׼��Oq(��L�T�6�GWEs>8���,�@PG�ݺ�����!g���MT�К�bֹ� ݡ�֔�P��_��c�Ë�˂��B<�/�mcV���/h]��MK�{#��SZo�_���ͩ&�f
l�y��\X��{b�筲\��w��;�aT����6��NZv ����.���N�>գo�wx��(ᔸ���Bz����BA����HQH;�����T�O>T ����-ۨm���S��s>>��w���]��Q��h����A�SI��䜂r�07nݠ�v㺢����$�O�]����s����V��A�p*�y������&�A]�ĩڪ��Z���sz��`A�O{�6���㑔����1�A�v1����Q�3���q�eN���D��ʔ��+OM)��[uX�hPs(w�˽Ze���1qV����C������}���y:�=6�mKm��J}�G	��1�BH�;�.H8"��}��A\�oX�y�9OEs>?FJ���NӤ;�媕�`׾>�<���C"L��KXB���T��v�[�¸�gfv5j����Ar�9�E� ��ݷ�n^�(��m��+ڨ��b>4A�p�n&qJ�5ڒ	�9Ǻ���㍞S8\t���}��������w���3�cF���b���>4mE[BFX���k��	���MU "j���"o+�tz��[���5J.'Y��%q��' Я�����
�PE�A��8]pa��#���8\f�w^i�5��_��f��ƍ�b!�-���2r��x��F�:��ܧ �v��VC��UӅ��ǡ�x���q7;�������� X�P6�84h��S��(�^<����TM��hj��f[߫s:�� q_U�t�v_4��̌L^|�5TM8Vm� kи����n��y����>֞�m���h��[��Û^>�x�t���R��R�^�8��MS�t�&���tu��;�7G�w`��sh�73p�eN-�p����ph���1�2��3�v�^]�2�����ռ�G,���U͉�Hg;r�:��5��c1�%@�M۷%�ĳ��n�M� �rv��ϲ�cb����Z�vwE��������݉�1�)2��X����I6�	�ħyv�b�GR�[`4�śM5/=F��6a��i�<��;I1�1�q�3�ڲ-�
�^����y^[l%�ul	[��뷅 ���pr�����4�cT���]yی�f�b&�v;�^7��z�3�m���3^��
�ge�ק��b$ZC���N�gjz"Rr	�����Z��h��$�*�p���yfz�p�\�c@8�p�4\��N�]�8����|sH-�p����iQ���ߎw������'|��T{%e>o�o���U� ��MF���4�8T�����~I���X�C[k��_�z�r�O�����M
�b�\�;Y�=o�ͮ�{=�_}��`̻3]��Lh]=t��;m���7�Yf�Fݱ1=z���|�����@[��
�@-^Nۙ:��{�y�+�%�m���=�>�^D���� �c� ՠ��*�8"�3H8#��K��俽�םtn.��΃z�<��rRq�G�<�+�I�W����u荷�.A�n
]f�{�Vfs��o�ж�mE�����F[�4�㦴��YY�����W1l�r7S;��ɅjIZ,X/IȬNAcV�8 �� ՠ�|�]����٫8�|�~��^�E�9���v�|�D���>BB�K�-�ڗ_� �D���d��v ��x��27�ܻ�sc���Z<��(=����h[��*�9Nj�pANT�9�ND�	 Y$�m6ŅSޕ�h����A�NA�p*�� �T���yv���z�`�:�v��*�����Q1.�hp7�b����K�S�����Hy�5N�;DP�gp���9�z ]�i�����5�;���v�L���Av�&'Ӟܱ^���)ܼ�X}�{#�y��r8N�-���́ ݡ���ߝw��8r.���"iU;;T���k�؇�����W�,ε�6��Q�Ŝ;*.�J<����V�H�V�a"gV���f��`�ŗ����̻��?�D��K�G�s[|������H:�W���|WQ^��`Lbrk�����%K�ERc�	�*Z��[iÝ�,a�-N��f戱}��#3��7�	�A���V�R���m`�FS�:���'j�� �j��r��bYyg�T������Y����D������<h�~_I������b�������h�qt��X]-�ԥ!�J����Zu1I�;UCC�'���Q^��m.b;7}W�vf��=�L�=��zU
B�JNŲ��K��:�/�1�`�A�-���4E���BFg6�;[f8����	�\����jisA�����p��N�f���sfdY��|R�r��u;�Ӡ��7\;���,�'3�!^�j�C��n�X�&�.�XYv<'�{��E���<���Y���|��!=A|�Y
 I��<jd�^}*S�{���ܤi����9�1�t�@V�����Y9���bg8)�v>r^o\��=:~���j��ߚ}�]U��5R�� ���]��n���y[��|���>����'��ŋ��BFg6�;e���݁�Fe;�̆��u��@�?z�`��blM]�GD�ׄ(v�ڜӹ�w-F�d�
�X&y9m�9�L���Cg8vA�2����uq��n�����9�2�\9�A�*�8�B�Ы�;[�6ͺ�L\�ჱ�vq�A{){k��
��@p �Y�r���Uww��	�N��T����A�����Z�
��$�E�r��󾇇�TE�_�bE�e8�����h�w\
�b*����R�xb�|}�����3���8j��Pܭ�w���~�:�����x��u�����P�T�*D�
�P�z�U���v���lY'!�
н�+V����v��Ac��x55�媒G'�*�Qh�01oc�L�Jy�c��u�GK봧w�ƻ�����wf�䣃$�X��Ͳ�_(�Joc;lwi�9����V�%��� �*v;�;Ȁ�o$�t��1�ɺ#u� Kl�{�{&v��������;f�f=c�5nEOv�m��]L:e�Wd��t���K0`n��+��r#����}ۅ�d]����,=��gM���!�t�M�eٺj����6gY����eC�����h�tyK�3;k��])w��q�(�N;��ǵ���8��U�m�
��V�T)Nj����vR����sS����#��3����t�H�K����4��@��a��ɛHf��kn�-��X͵i@�� �G0���p�Y:�vlb���[<ei1޻��^�w�����йs��R_iut�Ρ��u��/��f���Y�f�u�u
#7B��]��.�r;EC�w�)-6g</Sw �g��SF�9�z�1ȴ��R�'r�om�&	N��)�����C�����}{�V��<�ͅ�h�6L�e&�|�n>{M	��ɯ;oM��V�F���zzK�:�lH���7�gP��k{kQ�fWSD ��٨��Q��wn��m#Q*��N��ee�[wu:�JI�u���n�ût�m>^IW>`⬧�5:L�N�K��c�X&�<�p>ۅ�cP����Eh0�r�U��r)�.��5ca�f�W֝�.Y���qd�Ʋ��?p�i��3`B�4~>}��~��3Q&ɨ-"Z
��!�V���:��iǎ��<q�n8�N8�o�ݻ|||q��b*,lT?F���Pd	�*�q<co��;q�v�8ێ;v�������I��o-��nU�����y�^`_ί<ԗ����s#��\ƿ��y�h�\ƻ�s�?4�>��,m���5ӪT�@7t��rB7T���=λͧ]�h���_�w��F��o+�����\�4����ݱ�_�����_��eo���U�+r�5p��.77+�u��w���Պ�"ܮQ�6���߄ۚ��]��Ł�1�&���WDj�2s�s��r�½}�}��6s�9�`ٌ�g��H+۔�F�8�+e��'I�&(�m��Ę%���:�i�&��j�Rk��X���/`%%�T�8yC�r��=�.m]-����I��_��44�����V�=ڒ���'%rӴ�X��ے[J��\���-ی�J0M00����2�:; X���lv��]Y��|�9�6���٘ʛ��c
�Ƙ��3l�[e4R�F�4k�H��c�D5`���t��%� @�!��]�=	��t�NF*k�u44����Y��;(���6펇n�΋\�7g��3qô�M�<���y��v��#ԂV�Z�+g&�՜qj����}�E���;q�[v�9΋5Z1"5!�Mn���G+���g���� �Ӌ�]��.�\U���Nָ��Bxxf�ks��M[w��u�ۂ����n��jt[LD���=tsJ�k����+��p]���tw-@��P����LK�]8=!�/CX.�7.��w�����p8��ɽ3�63kN�]�;���&陣Z���:u�sl1�Z��!�evc<f��L�����$�E���+��(%BE&z�ʔY8.^T�����!ڔ�y�)�w/	q�� %��`�ٷq�S>�3q6ǲ�Pݫ�=��찁�i���!f���]sZѶ�j��)˚��
�2�p�MQ쌎43\��Ql�7�z����S蛵�Æ���뭄����s����vm��	�E�=��%(���P��9,�f,f2�:k����8K��WK��nrrμ��Pk*!s�2�sפzC��.{Q�5��tl�����5�z����q��/8x��e��Z�UPjLa^xཥ�2�OX����q=�r�f�Q��t��p0��e���V�1�ª��-��g�}��s#���������k��3�CC��E�Na�9��lh���8���<%��m�.h;`��քs�%�V
9�k�{:����f�$ݺ�%!v��v��O�t��.� �v��ގ5���h��G�%��2v��ToQ����77��kmY)���[��y�z6����#�Pn.w����iѸ^�<p
P�,]]��YWv���&t������o����Ŗ�A�B�Z�Ale�#M:rF�6{9R��" �x/�|��أ.��F�T�ANgv����Fg6�8��Ϟ��F���75��C@]�x��Aէ!�B�y{�Ԇ1�M&i=팮�ttⓞ����>C�t�5��������zp2|��lwn�8"�݉�BtV;����X �	�G�v>?�<��&�N 榪^-T���<�6qX�>X�|�m1M8��U �wۯ/{��8��m�g-8!�hd��3	���X���r5I��S#K�����I^��kg�^��}gq�v9�,D�a�|��C���A�q�8�W�w�tl�Aw@��`��ղ�f8:���#�cku� Uwi�w�,5��#��P]n��L��i�6�Eb�~@y��M����
{`{ֱH �҃���T��5ܻ]���A�S��!�����e�|����/RT�`�f���kzS�7��
9v�OE���6L4��4V�٤���&pf7/��D�I*�z|}�m�&�g��Z����kōϺ�C����C�2��LP�p������mƀJ������5J��,]�c^Q��LF����N7j��f9�9�N{Zu`g�;F�"�Y��)�80����꣊�\�]9�)9U8r7]ؚ�q+�U�9��a<�n�\'%9(�H>�B��v-���R#^�1�e��[@�c鵳�������]V�E�����yͷ�#-8,n�r*��[�A�z�#�G40g�v��%ظ��sa4���NN&ܨ)�ڲYy��t�1�85I��'��k��tM�����i������]�����T�
��YJp�R�)���{Ec�����F�s�O/�K��9)؂� ��ى�����h�5)�L��C�s]�b.ӀA�p�{��*r3��Sk6J����Imv�}���ݥ���oc���[M��3nt&�$oN!��%�� e������C��X�4�2dɾnic՗�v��!�^sm��He�b�T�؃T��T��ڄef�޶	�MZ��5Kr�u�bƉ�s�Ӽ�1� & i��=Nؒ2S�S�nd.��"�3���"�ï6o<6Ogb=([vЗ��Ӝ������ų���A�T�� �I��߮"�3%!HJn��V�P �H%oH� x��vR+4v�I �& �.K�0�$%��>��/�9I�H=^�^��q��|�6X����'��o��.m.��ؚ��' ����.�����wS�z�y��6M��;��f3��m�ER��:��󼫦;��؏k� ����*�9N�A�Cm�;K�����n9|��5��!=?���'<��jk�� ���-U.;�ޑ����#�(` �xFjgN+���l_uxC����C�i��e�}��!b��<s��2�8J�j�u0�VDl�#+���WN�E��.����ee��W=b��o�-��2o�sKW��o��AǙU(0��8jd�$�BRț@��%V(�'h�mg���k��~i�8���5ı�N
R*�Hg�1fc[�~��d+.�D&�\����ثULD
����)t�؁]r���������t�=Ӈ"��ؚ���wS�0�?,���;-p"'�;K�F�Oy+^���8,j�r���Wp�^��v{�Xu�q]��}�;�D8��l�p2ӀA�p���>ێ��s� ��M��A7��1F�5���T����Ս�$g�71�7�o�Ns�y0pAo6�b"��U8^qo�9�T��"[u�1��՘�6E�sIb�~Xa�t��	�'"��_xR<wKa��>g�A8鹍ܳ�n�s�sj�eP�.���NM��.��w�;g�:y͗�br�4�r*�ؚ�<H�R�Ѿ��33��s���-�wu 8^�o��c���)vw�r��(���}��M*�������l�<	�9��U=�œ&��F�}�T��.t�q�]úN��u!���X�h���ј�Xmv9�d�8��V�m�C�y���vg��x�KAS�GPCָ��`�W8����7�cW���ի��*`�x�T`x�$1��c��ݰ�#�
��<�h����{2�!AΖ4�X��-+�5v��gGG;e:	��}����{�.�tݘxƁ�f�p�߾O�o�}i�Sl�$'������/��֍5�p=�Qؓ��N�/�i5�˹�ʼ��)�' �3 ��_�L������N,j���Ύ�f��q��9�p5�T^k��fM��4s���©Â*���
�R߭���U��|o���X��吞����'bۨ85K��o�g��[e�2�h��#����t��ȪNAaT�?��xZ|�]��A&=�/�k�!Њ�j-�L����`c�pD��T��̦�6�1,�=q�mx�[����T�ٙ�ލ�әx�$�K�!;(�"��&����Q�`�pAm���RU!H�/s/ۜ�ZG[�+P�]��~ǇR�8Yp4���A�vpnӲd5H	XM;���]ֈ{ �H�A�6�!ݎ3�{1�S&'u�9)A]��;R]\�Â���c�v#�� �S������R����9�|�&�
���� u8r7S8�q,`ӧj�L�3�0tezy�֖��l�p���@

����O��A�O��˾��n�sx���/#7���=3A���C���߂����{����q;6��g��}W�'�R!#u5RCѵ����~K�B�H��g�xT��G~��ή�~����< ��Y�U9w+E���Dr(P���BB�!��~���^��AB���@1�8"�a��������z�[/��bЅ�V�r�85������
��Bd�U'b*�9�]���7�,9�N6�k;f=��/1�I2W Z<��w]��!�(T���b*k����� �(${#G([����[8M����Ҧ��t*�e"i���w:�Y�1@�k�9��Mv�9�z�f@͋�0�vR��P��yсwT�U5�*"�3��L��s;M[����v#����{������k�G{7v3�l�Bo9���-2��'`A}�"vo+gX�;���N]�h@�q,@�N��RΞ��}��D~ڻ�{��90mb���X�%5�;�#U*Υ�/W�7M��ݢ�i���_>�&���J�ε���7�aA�ӲA����s&L�捪����mu�?���@D 3�Ѣ�Hx�j.�Wew���d���l�p�N8v4��{QN�#5E�)[��Ny8"�ҩ�N�kH�+ڠM�r,�&4���� @4\�Vby>J-cEÇ�Y��+z�;����C��e�u�9N�F��>�Όs���L����^n�j��b,��l3���Ą�#����J�A�'"���^iAN�g\����6��xp��d"��ٌ��gP��,�ƽL�[!��4wVY���D(���}�����<g2��-!��ש��3W���K�Rn �N��G���囕z3ie
�
A�C�*D|4\�T�Ѽ���>O�H�'���Y�A�M�,|�."v ��v-J
^B��mi��N>�C�5R����މ���x�Ç�� A��pDG��F�s�Jy�!�J�R|R��`��N�4V��atf9vn��M\)�����+�2�n����4��-ȋZǷ�ݶ�\&�!;�q����N��%Ho��/
SX��21�v*�}���D'"����27�=�y)}�\ ��L���f��	�Z����{�=��E�t�k=+�l�Z���5��N��{>�n���.��]��)�ۇ�s	�A؍��.��p�x�v/ܷ�����` ���:0]��F	�<|���F[�1
��,�S@1I��{��n�F�����۽�[w�<4x� Lya �4n(����8�s�{]��!u6x�]�&5^v R�7�X�]���&-S������x�K�b�Ac~N�1iƩ3��X�5�&{z�6����*mÜ4\Z���gn߽ϽT�/9���8h�3o���wb<��tx��Ֆ�^؋�VZ�n�俲gϴzc>@Gg�5�6:��b��,bW1�+\; B�~TL�����?�_������mer�5�����Y�.X�1�m��Ҋ	fZ�fT]�� ��2s����X�R$��\�	m2d�!����>?8��������Р��A]��(Z�H�Ye�&���P��І�%�!s1�;9�B$J�M��D���[{k��5�{�	�&l��:.�썎gZ�ܽ$�ohi�q�/G�؍��%�"�ֵ�m��:�ţq�v��eJh�av2gJVX&�"2�ia�m��KM�v�>�ہ<�۫^����"�ple�$�*Ѳ��w{]�r��❧�-S����G7�m*V�����H��wAڏ�U����&����z�6�'(ľ���_p�f��8 8\����|!�gn��|�΋������w����y
��g�[���Cv����Xݠ�z�Aï�2ʬx6��Aj��۵���/5���9HY3\8"��FA{���=���P�҅	~�X�7N̙�����s�hee�����\Ac��5��X��)��M��؋�#0Yk�C�^�A�p�f�C!T��/Oy����	}�\������S"�ΝX�ƭ8#Y2׆x!�0�/H��*���g���|���p�:������Az�6�l�i�`A�9����o]	f�=�Q{�τ}ջu���Fۆxm�L^"�ŊtY��{v��1�&�M����L�pA�vsT��R~���e��W��{ʢ��^���[����A�5NW�v�A؅���1������<ɥu4ӑ��wrv��j$2�I3^���p�C����˅���[Սe���ӑ1�NN�\�D���zu�;�4�-�ж�=�����sݶ���7��7�	r;ip �r��5���Q:���痊�N�ѝa�ˡC:�b��A�j��")���z}^��I����?eP^�y��� x� ���1As�]���ݜݧ!{wќ��	Nz�^k�����j��vWr�Q��ux���7� �|iN8ȠcT(o*^"�� �T�T�I �ˡ��N5睟��qGf�ߡ�xLv�����	
��|��Nq�7�=g����K<�4�ɀ�If�B�f��)D�P˻]�ux>Li,)�>����T�4S��޻�y���'�yͷ��9��N�q�O�U���v"��b��R�|��m�5��N`Njp�[�ܽ�vz����.�A1�A��Û6VoS��}��w�B
d6 ;�.���@"�3ɂ��荗�~uɓ�^#��+{��{e	��f���C:�͙\�ۻ�ܳ��Pm��V#�S���}ZR�n�!,�	&S��n��rҎn���aQ��"33&u� ���0� Yx��mᵫ"*;��XwcB���0nŃ[��Y��G� w��ϗ^��`�f�ss[��Kf^���ڎ=��Io��O�C�=׻���I����|[�{���o_s��َ�5�.�=�����賵����c���w{4��s�m�v0f�v��=݋ӆ�{����T�r�gioM�+�君�wU�'��)���1��n�d�t�	eU�9�Vk7��͙x��
OTJ�,�ͽ����U��[|��񕔴v�A�)�9\F+���κE�.ض6jcG�n3��c�5n*i٬��Zr���$oJJ֝���^�!BMָ	�M�'9��B5A8���Ϸm�FPƳs��;O)��[(a��;}�w(F��#�Z��3�0�f�'W7�c��x�:~��n@��vڵ�͙��Ƙ"�+)�鼙������%�y�i,�k�tv�y+馇�Yh��՘7;��V�`���8��\5|z����4� :b�a��3��.���>��2��;�Y|�֪P�JL�OWάR�7
��p��޼ٖs�Ů�Ch���j�H�o���l]�M��;�ٳb|�J���������>��ɭ��5�(�3�w�`�f�e���ZT"/2�$| ���QN��w���A�(�I�<���[��uH|#�|!̵�Y�H�yf���N�&���5Շ�u�gw
wF����J����kh���R��=8x���fc�^� ���O%"K��Bʀ�P%�,�:{��uәE^n|��V �! 7�(��!c��7Мw��}���闌�C���.4�M@�T5@)�<|t��㏎�q�q�nݾ;v�����HJ�ByWtD$	���>��$���m��㷏qӎ8㎜v�۷�o���'''Q|�������6�-ʹ����F�}o�ϟ=^[ҹ}U�͟:�<��wk{��/��y^o/�?�כ���qg��oR�$(�v��{�N��Iީ|�5�;�䭒�q;K:ނj٬l�,,�c�>�-���}�����ۚ�9�W��F5�~�_Us�ѹ\ѹ��w��Q��h�΂�?}�2|{ovܹ��㟱�u)�*�
�>[m4���!��չ�ٳ~���1�K�7��A��R�Sy��P^���5�l�SR� �v�3{���{j��l�h/��Y�6�c�1�,����ع�N"�_�v�Yуp{(��әs�=oo��x� ��Aݰ Ѣ�N*��s�=���
H��$���ܻn�+��]����G�u�ne"�6YY]�G%п{z�����r�p�u���l�|�j3�n���`��.-�z�z3�[����� ��N�N� � �{1yq��ݱ��`Ao,`.������U�/:��� ��ETP�9,�����)��� �&zTC�T���Y��\i	;x�NM��O���h��	��;�	8$���{�*EJ�BG_5�(T�H�Ƕ��^Ր����]�	��\A7��Ҟ�籔^9(�B��B舺�4��t�yu�cks�ڏ�"����cUi��vd�k����/�t:�YتvkK�z��2d�X����i�'j@�p��"� ѣ=X>[Mb�;�6o����B��5�3�}l�E�gkVD��^�Og��rlû�msƌy�sq9�6���ti؋��!�u�m����M�\.�jU�MgH�J�CA�OWk��%���o��p'x!A�o�tC裂f!@�2�;6\�T�3�H9�E�\d&��n����]�x3/m��.��~��.= j�A�' ���pj�m^ݦ:�?��u1�&gNR�j�Hظ��݊�V���Ez��|��2��F�t"�0�15�o?E�v1Δ��ԃ��NU'n�;�z�{�[�.oo8 y"���[棢v1*"�Ñ5� ERpANT1���;>�7P̋�������\A7��9�85I� �T�3�G���1ꨤ<���Mz��o��ڼ=���n�̴�ZR�6�I�B�PZ��ΝͽKs��f�aJ�ךj2_�BɣX����#����&A��=a�O���~�Ф5�ҽ��p��:�st�85@X��clOng�r��TM�n����y�a�ƫv�-�X��J�Gnݸv�.R��8�gv�Ň�+�ݐ8�Uv8 �D���A��qt��х�K�!12�-�$-3���K5vc�x�Um����5��x��.<v�v��Sx���x�*d�*��z+34�tQD^HiF?^`+��nb���2�:��Í/��to$�[���`a^�H����c2��Hy��R�R��-�9���6s��*��U��$����AȞvp*�U/MRv#n=|^$�sKѷ���~��w������؃�T�;VOo��]`�.� ;ɞ��"�ÁT�w�wf{ѽc�q���N��ӫ�,o��f����A�U�q���C�G&2��Z�ñ�Ȇ�qo�׏��F�������=���o��v#��b��J�҅�|�����za�M�/JՏw�޿?]�Ń�Rg�A�p����R*�Z&?���ڼ���� ����m�G�pY��%��.e�꘥�]C]bh}������ӎT��MR#�b^�nV�<LCv�������G�Y��5�ާ4�P�P~0���n���g��$��N�]ʠW��]�\������Wȧ�� \���i��ݕ-j�`�!;u�'Ηo�c=AP=�ndɓ��!�|������VF�\�a��s]�pA(0Ǳ"*)����nq��p{��Ai;X� ��&sT�&0��w�H'}��ǌ���۾oo3�JA�q�]� �ۇ"��@�ŵQ�~���h��� �U�}b�A�4y�Gv�R88�v�n1i�ü�A��>NZiCs&��pA�@=�� ��t
��93��sv���P��s������M�����Z�	��~����v�8H�DBy��ɽk��Ӻ�6N�:����J�PԆ6�u�����p�
��{M/b��N�u�,����V��{y��6�oS(X"��V��v�ȪA�Iȟl�7hz!��[`CԀ�Câ����a�#����\�zӐNjƩ �F���N[���2��cn����n��s��&x��{W���䲹)��2
��\Gz�uv���3X�x���m\|��w�c���
i��s� 4,� ��Eأ^�@�h�`)��	�&�k�O���P��sZ���E�v"�U;�b�� �8`���+4�=� �@�d�Ρ ��7I���rΛ��q���ڇ^A�&����B�����<]�-��^4h���9Q��Z��g��thO|��5xpp�C�W1i�����K�j�ozոr'�	�ˣGm��@��e��X�sc�eR�D��M�]~O/�Ĳ_� ��!|��ҧ	�i��߷��7���G��H �5��
,�<A�k����b�y;LI4r>�x���-�Yas؟����lښ��<w�,k�;���F�yϥu����y��!�`L.Av��ES�T]��v�z�e_�L���\���8=l��M�PA�q�`�ǀAcv�;!v��nѫ�s�?<��!�@eK@�n�r[��kۡn�=��z�sM��F����ڜ{�^�Q�>�j鬷t�'S0����F��{ﲤ�X9�j�9��
-��=3_�+�Udqpb�η53�	�yZǲ�5F����&@0���[�M��1��NA5IòU8L\��������mb��WQ��h����N�k�9a�����T������_��=�Olu�&��k���V{�7%y�١��M��\ۡ~>[���d�쑖�I�����{��z����{��8�G]6̦{M��8���I�� �f�6�'x��ܚ:Ã܃���_9��l��������Y�4��5,�<ݖÜ�4w�8��[2PB$�ӐXJ��@�&eB���X2I ��E����Q��w� Ԡ3c�h�pA�zc��4n�.I�ԏb#�r'\;TC���=�NF�?:��8�%y���yV�Im��k�!�!�e����~p�Ѣk��S��=��#v:��媲=�y�5���4D1�����b`�ܬ�1}\�����	|��7w�m.�{��Α�Uwc�����Lo/�z1ۻu˳H�1 1���,VĢ�t�;�Y�t����>>>>�SWX>"�f��G�1�T�J�J�
&�f��6,i��H��y+,���6�&u<ksm��p5����i��stMAS33KS�zl��'`��/n:��qz��xm;ng\�%�e���R���u����mliu�ZLmr���c�g/���O��M"mb�">6*�����%�]����dSd�N����]"q8��n*�+7wq\��C�f��6�P),�g�����g����Լ닣�M3�s�wms]/6�+:�V��w0]�>�K�XzS�A��R�C��3sM��N�~'��y�k�V��xM��C-�^�t��dU8z�b�C�
Q���a]ï�<)�VC��a7~��>~2:uP��ij��Il�і,�$�a��ޠ�H3^���f�{f��z#6f�M���x�sM!��{�bƩ�DSy�R�]�D�]Ӝ��r�݋�T�nnl%�ӡ߉�<,� A�A�>UY=�փ'A�ʐ~��@A�B�T�T��I;<^��Q�豣6%f�?��M�9�cRg�{�.�v'ط�*���Y�sn�1�n9��kV|%�;�OnɈ+��g�n���dax�+��#�R�S�"�9��=m�n��G*����4� ���pb��|Vi�`Ai�ݠ�9�Rv# �͒c|J�U�E�UXVH>
y�)P���)R��Ymv�B�k-��r�C�+-��*�RѮ���,�á�Kj���O(I�t ����� &L���gi(���>�f�]�:��3�p@�R�x�F�u���ӕR/4:����pJlT`�TೲN��R�2�!�M���u�o�cςB����r�!!�*��d�*a���}ÍS��9�A� �T���w9>�J�x�sMpn�pFl�P��L�v8�j�PkŪ��AN�ƩuN��j�ߘX�e4��|{���П��</X��r��� �T�BG(�豁�˻�t]�I8���=�������[LeRŮ�Ʊ4=z������6ӈ ߜ8U �ک7�"��x��<� d@ݥ�z,`{�QQ
�^�ga�P�Ct�RB��P��5"�o���0
A�nz��wJ�y��C��A� ��EW��Z�3�^�c�6����kS�S��T�X�+����|�p��m���\"Ŋ�h�w��:�(�~)���gL�d��kvhA!�3��NN���|~�C�}�Q�Ώ7/�b7fj��h'IaZ[�&L���$���t���	��3���ٷ#5ñ�eȪ@Uy��D�EQ�LG��P<u���ͫHv���O��%�@ȶ��A%9�][^%�������V�"�:� �T��0�H�zq�Ѻ,G8�߶�v{��<ɬ֚C��,�6�b*�؊TF����;��/dxY��)�1	˨��s>��ӛn���up�Ӧ�ș)�]i
�S��W��?���\�Z���Y,��>��{vu�s�3��ptMM���P�ٲ�*�8L�P��eF���Ok�b#;w	"�3�ZC��݁\g�p>�'�:���rM� �%OS�0����\�F��;!֠�P�  ��j��q^�9U";��ӲH����]y�8�2k:�p@7h9qñN��19�ڂ=��B̝PϞN��I�l�P�*��ۦ���=�:�9�ᘛ�R�m^���[J_���r��%�k3FS������P����B�ɵ�(�&�!Q>��9l}�z�W-�8�_i��h�G�q�|�o7G�N�
i�wG�o�\!׫-�9t�
��]
�R�S������0��z�.��-'������nS�ܛږv��H����A;�K���88��ǴO<�:�=Q�صbf�f�;Z����;���A��w�.�8��ӛ�=8�r�:��\R�W�n���g,מ|��p�������j�g5I�U'"��|��N��r[�x��>��r|�ӡwl��������(&!�%����@ߨ.�=�YM�E���4��r�Hsv������俹r����ɽG��=�'��� �d�7�Y��@�Zk��-�����M���K�ub�q;q�{s���Uf��3h�گ{G�P�B�B���|�¨zB���U���Hۢ�ʾǑ�f��wd랂�����	� [av�C��©�F_s_o:�h��K��o�����\��9r�8�Ò͗���I]�k�FdF���0,v�qs��efW�Ȍtjq��>ݽ�@���u_RΘ^VzOKN�[7����{sku)�,�ڪ,Wa�s�!��u�k���
�j��\���;�u���nP�鳛
�PR��n��<�+�N9���L�욆���!�����n�8�8�w$��?1w��Ӣ�ޑ�*ͩDv������{��;nl8��&�˻(��1WQ�oIe H��
>;�&e��hi�)�jn�n��O:���������c�f_#����jc�+�9����W�|
��޵�ݪH�W�&�\r���V�{�y���,�l(*TYu�2Z�Zچ䵀��]7c�L���wvIWV^1u�lvK�9f��+��"]kǗ�WJ�f�>#�,�|՝��� L
I}���*㓑�v薭n�¹���7���ݪ�����ͅ`�`�ե+ucܕĎ�bL��Hn�	Z$�v��'b�%"�WQI������Zᐈo{%��gHn�k{rTŻ�ݛ2m=m�׮��/�+7y6�x%%-���ՊQ���\�$!���Y��vV����&�r� oܶ���q��+!���VWV�ȎS�*��V����A0����һB�f̹{��켘�B��[���$@$����Ƴ��}�Y�U�t�*n=�(���b����̟>��+�_W�?Z���s].r�I!YT=UBH���v���ێ�q�t�nݾ��>>>���|{l��L�{��;�����B2H��$5
�cO����8�n8�:q۷n�>>>>>xC���QSt�1��ݒ�ۑb3��`�dƊ#yˇ�t�t�����r���D/�qJ_W��Ė{���|W���ε���{0B��$��nA�wsF�;����]w](��ұ����������a4@B`�(��'κ_[�"ɹ�ۘwr�e��ou�{�^묖���L$d,�D����-�$���I����i�{��x��x�=ۂ�5�מ�4Qs��0F~u��s�n������Ke��P�g��OC�%[km��:��q�Gg���U~�����ߛ7���ڽup�	�k�;'8G.�v��ݚ���sO&�-r
�ζ��ϝ=z�N�y�9}�����Gv׍�{H Ft�L����z˵��$��^�z֎�y���Ӻ;z8�z]U�C�"4�.�dY�ۦ�N1����lg��\l^�l�],��[fҧ ����;��]�p�jqa0۲��Z�wN.1�!n�l��[,�,RYml�i�u�+Y�116�4%-0[
s���6�K����6%��P�z��%��r��9�T��6�,��ֳg��]���a��R���[���m;�1��g8�ݮ�Kt�oh���3��m�g1�P.��n�W6:�ݓ]Fŝ7v�W����{bx偱�x�{�s�G��D�C����p�pZ3��]c�� ��$v�:d8v[��0@�6����Z�+s؝<�:^tG��;�l'O+�u�`�J�@r�H�mٻ��)��(C;��%�n�����%��혻64�+ј�����Z3cJ8�����jR�G;r�۴��0��Is0ʖĀ�V۹��ն��\uwWQn�'X�ފw�1�Ջ����,46uMi4�k�<|�w"�@��$!K��%�?g})
�Y�	]Z��usItڃs��c�{bۙ�o&s��u���&8��g`	����a�M�Oi��������s�]bZ�E�Jqc��4u-(ړJ���F���k��0zn�l�ڙ����,�q
��\ݮ�l���$��[g:�:�wSj�-{v�,��.����v��m�n�8���g�x�<�'���!+��q�7Z�:u^�8����q�\�lAn���(ېSk��&�{�Č��b�cKcW8w]c�V2]�p2�8����l&k��,�r��f�U-:�UTm@�奵�Wn:���}B�z!o��y<�ݶ���mR�[7/Vͼ�M�g=7�Q�Uj�I!D5&���D��N>֚h�𫜶�+Z�JHxv��D�	�҃��m���y��sjt\�x��(��5����Y1.�b4ɘՌ�ĉ�
b��+i[��-*16�51� B"ioj2�!�Mz����Ŗ�S��B�eF�)d!���#�FNf[�A�J��l�n�㓬��9�"X�R[](�b�;�	��մ�i�j!Yj�+7wjV^D4昡R7X�y���og�>4�~$uu�4�R�Q�7&D��m��2����qS`$�AH~G܀v�p��N�Z����+�K�>�!E/ug��ڠ�4��'b5I吤��cv�13�b&ⱹ�y�y �'n�Ƿxzqz�Vt�&��5���A�)�̇���x�6Bi	�b�A9I�H	��2��n��Y����Ĭ��}P���\E��v���n�rS�b*�^�f:�~�l6��A�{`�bj��������EG� �N. ��iـF>x���B1�3���=�[�]�-��
�R��\}q�Q�F�p�5ެ9���K�*����3hik�Eۻ�h�W��1�K�p�ǂ(C�r^ݦ�E���i�c��D��QMti+e���[?���A�?�B[����j�I�ssI��C�����e����3�c��a�B������!�B�������A�������Q}�W������{�!V��룖V`^�ڧ\������r0��\Q~����%E��f����~K��t{�qĒ_d�#<�ŷ���Qޟ��u7���m� ݬ���عxM��-�l���,n�rS�b*��U8�E�����H{&e��^���h��]'��w�5R�)�����)/�c�_V��A��g�uni~��}�Q�[w��!�F
�=.T�� 1�ͱA��r*�8$U'c]��.�-�6�Dyu��B���Tw�O
���+���8�A~�<��3��O�;��ݾ����������]`e,k��K0e�	�6���18�t��b$�%�BO�������^�x�8p�N�l߸f�i���Z��ypqk�b��3�mn��V��kQ�T$*�	�GvY�z���1��X5�ڙb�ݲ���k��-����3h8 �����B�FN��;;٠�s�E �����"�B�T�(Hj&-���6?���jJ��%��L��pcc�\��G�Vu~��[w�>p;�>����/�I��YإܝO�P�3Sy�ɐ`> 7�R-|��.��&�O��+�A�Y* ���ݦpj���N�<��1�����&�9rX�w/ES������1t��U�-��8$][<�����q�`��Bfa�$5R����?t?�}C!z����}�k��{�ͻ�౛A��A��
�BEN�dS�>���i�]6�!��=�Xâ��A�wfx;u[[�N�UL+;j|ɿ?8�t�"S�U8H
�(dF�����ѩ�q�eq���t��.C��x�Yj���A5KZk���B&x�\:mm��M� ���0�y:+7������s=�pH�L��U1���m�ЀcS�X�&sT��eT�@j���+���w�i�WyN{Ϋ���sn��Ag�WB�*�R�R%Ys��J,��|�
�;j�}��ݛ�{�ML�8�:�7e��S!�]c�P��/0��J����{#2�b� ��c['=}]oS�v[޾l^��8B�ܡE��.���v+�uz���K�<cl52dɓ �bך-Q��UC^{j��T�"��2�vyO�fV������Uן��9��8$]-�J�H�xxHj�ߧ�
�����m��2kV�N���{\b�f�M�!4���0�2ˡLG���A��NM'����Է�z��ͻ���׆u�y������j��=�t��BD2h@W��#���.�� "������[��{I����Pi�۟H�j�]�˥qGg�X�8�q0ql���p�ٲ�hG��8����rē���y[�]y�����t@��K¤T����?}���I; ǯ�4�p�[U�i3���ڻz�uy\{=|4�&� K���F������B
�UI�a"ͭ�Y���������W��Wb6�1���k���]�g08t+���������I���{�!��Pp�n�#�3���w̗���$�ʆ�{&a������1Fr���\��ˡ�8�G�v� ɓ �f�v/T�<��9A$�!��>�!�p�հ�<���묛����d��vӗ��cb�am��x��6��I�mͺۅ�t��&۠G�Ĳ\n{z�9ݹhK�#C e`\��c����O$ɝ��.���Wh�WϏf�+��f�%Bv�1q���J�amͩ��uaa49�g7���I�e��i��͈���n��Wm�O~m~}��]�S�U��%���AA�(hF�DU�T0s7Blح����5�u0��H�p�&��y~�^��,�����ٲ�.�u_�noW^xWY���D���Ezh������9���:\p��3Ң�'�7iȼ�|=Bϳgl�9���ƭ8�7������m�dpӼ4��9�G�U�c���18p��"�"�3�TC�f9��=�\�v��}d�V��K�瓂�85H �Rpj�պ�����N�V(w*O�A
x���s�sxr��Qu��|l�Ƅn��8^�U�@����VMRvQ��K�0�Qw��E�c���9gtR��/��N��;1ñ�E؊�-��z�ZnԿv��HS��;�0`��fy)�T]�v2����1�:dL!C�P�K��,����0p�"�"�݋R�����D�5U�c���G�g����|�.b4�l�� �'b�Ѣ � �z�؍��]��w�R�yWٛ�T��Y��Yq~s�{6k�=+��Yľm}ʕ�d��L˓�93�G}�K�@��!��8��L�2`��ށ���pA�n�ṿU
�]g3�3�.Aِ����2:���,\C�_<��j�sT��Gx��Ǖ/�� l{Ժz)�2˼e�Ӝ�i,�x`4]�/^B0"���ਜ�"�S�,�g�>��=*!�=���m%U\?Sm�Ly3��܎�����0�v �f��AΕx\9�g��ƚ]��W�p�BE]N����S߫9��;`��ܪ��T|0T��|��_��>�_���F>Z�1��F�3����\�Ƚk՞�N�=`W���:I�C�.|A�X1�EJ�X�Ť87i���q9zw�r��e?��i�p���>��pA%ÃGK�H8"����#�H�X����4��v4���3�<�IUO��m. ������.�Okn��ڬ�@{6�tJ4�O,��@����"�ڍ5��C>�g�[W���{��u��_T�+��u�<�Z�8r�k�Yх��\#���q]l��ə :�0�__�苕eEۇ�Z�z�\���=�J�B��O���0����_����gk8Z�y�����D85IȜr��EFx��i�2J��b�I��8�p=GxZe�9�T��;��k.1&��d�v�B_.�20౱�
��
�-�~x�3{�\`�홓0FlQU^��up�(b�rS�yi�r�E��&7�&)��d�;�:r����]�32�W<���paT6Y�L�f[\`g��O�c�rɈ�BeF�1���ߴnwOJ��|�\P�돵��-�B��wcJ�sT��^Hlͣ��g���a�O�A�K+^��,Rx����	�A�}n��E��Vֺc<�F�v8pEyݴ�rN���R�&�u���[!�ҫ�i�p,}���9��ܴ��k�>!f�3�{j=X�y-0�� �ݠ���~���yީ_����I��E^�A_��'��'�IǸ�T4]˄M��aޛ[N�������׎��x��OK�~�}�����D�e�7ߗ�]��5�\����SM{������|���T��Rp"���/�b��CH�3��~��_��y��H�T�����*��˴ uD��B~�m��#�ӻ�Y^ �#/d���q����B�jf�&s c�A�m��o����"93��ERgi��Yi�\N>�SxSƪѐS��);���(ӧ"��Ʃ:�9��Lm����S*������V�ҿ{/P#���l�X� .�-��6��Y�B�r�5�p�u=
�T(y�"+=td*����S<7���}O���.+�ؼ�s8a�@�P�(Wܩ �)�B*T��}1}�pT�zаEk��v���z�F�u������rS�MGF�����6}����U&R�$4�(H�U
��������=W~=y�l߬��z�"�5����A�C�j���c��v1K��wD����jt�[����>֔j��*����ͧa�����C��WKs _iM��M�ub�7=
��Qd�dɾ  H��ev��/瀮�%�;��t!;����`
ʕ`�������Z$�%Լ�������^�1-��tk���΄6�11��R�-���tu�ca���%+A�	�B�KuDm�K���/Qe)�E�T,`a�����8�*zx�U��73Eb��:N�8ps��t���RxnN=ٛ7<q�U:WV���#�'Cq�edP����ݜX�ͷZho�AI����~y��Իm��L�4�Fz�0��m���s	(�!�$�|Ac���Rp �)���h��-<�h����[bD�1�<&��aT��kvf8���ޟٛK���Ov8������5�%df�I���R�եo���w&�UT�X�=�V�=M���\�IͻJ�</ϗ�)�ݸ�
��T��n���J��\�]�x��UI������t�y��ު;�<��p=�:y��B�5U;
�S���I�=%�]�g�7c{�&���VF;sZ]�U�U͖���u޷&ko��J���a����*t`�6��Z��ׁۡڎ�^;E�&��|����<��7U8��܅ݛN�����ʡ��3����uh4ݽRj��W�!���N����+n�E.��V%um�l�ſ?��VO�����B��%�
ˌ��K��G����m��ϓ� �y�>���½PT�קM>���I�<w�{�߯^���w�4ژ���iڪ�Hu��p%�\6מ�5RaU][�ap ߝ_��$�Y$���q�N �r�����2�I&z��A!M�l[D���K7se�ru<�������� �d#y&v�@���U;�UNZ�`�8d��++0��W/�ϿU=ߤ�����nn)��XF���E��FJ}�V��AϨ:{7.�Pe�[����)�O�����ֽ�HUS�Dun���W�\J��[&�QG\DO��7oU����.����rg�T��T���Xv��F�v�S��3���v�׈	�ڷ.�^z�^ ��X��v��n����<����M�"�n�0G�Or".ma�E�wE���k���-�sT����u�%��U�;��̻׉�S4�[��Wp���MLM�ڳ��n��[�n�ٕ��k��+O*�7���n�d�g6c�(-�,�՛��e�F,̾To7�H�9���ާ`w;\�N��v�q�XY�w\-�s�En�r�W�sT�J��ؾ�u4VJ�S�2A�z�K<^���Y�:2fGMܼ[�	&��J-��"��a>��G������{@��#YTv[�j�ݎ�N��:wF�}�^v>�*��K�:������S7L�XJY�c5uO;���}a;�Z9C����A<�*���
��m�tbJ�]�{�1�J���f�<mՇci�A��̬�'2����n�fK�s��7�SWnL�g>�%Α�z��ZU�������0�6<�!]����jjL�$ή��W]kk���D����ˏ�q�D<��OG2�^����Hj��(
�S����//�l�k$�
��޹�}������R����PǗ��goLi+b���gC/����*�|����[��2�.��I\��^,'��ws�V
�m==y�2듫��#����ճF�,�|���W�e���3�i�r�7���������5�� �Ks�ݼCT�� wB�+{;(����}6q����]%�q�l��S7 s�Ԋ�wx(��nKW��՗K�T����4(����d�&�e�4 Uӫ+=��j�倛��IcG?Z�Q9tG+�FEwqˑ��9k�������w��z{||m�q��v�۷�����$���4y�ѹ��1�_ݯ�ވ�F���K����{Ω$N��oNޟx�8�8�nݻv���I�*��!F5*����n�;��R�r~��^�r�"\�I��� �p��2��wp�9��N<�2_�\�; Ȓ��錽�a�κi2�n�qEr��$ˮ\���.��hBn�0!��ˮ]}v��.]�(��wh��ӄ���+��&�]$(����ےA}�����O��.�p#��lg��qs!s�9��!s��aC �4X���yr��e�LFH�;���)	�n�s����A�I��y'��r�����$����dr��A�Ή@���]u���n�/81�`[����b��B$�J�Ww	�o�\ǲ�w�Mz���V�o�[}*ge�܃��8 ]ߚϮot��z�+�Y5����3#I���cs��p�U-��]��w�Mj9@�l�oE��^L=���6����.-��UI�U?�lo0{��9������1��
mq���j�[�uq�Z.W>u���O>a�/�<�[j�V�X�'v��=��҅R�
C�:f��Xϴ�<�
�h�T��9�=c��l�=�ؕo�'3�ϫ��j��YU�W�^s�/=_.�s� �y��tG8HUUW�������F�y14�������3���~y-x��0��{�"���&��|��&p�������o)z�r�7��M/��S��WO�t�c<���;�����n��`�_����˲u9�)���D�S��+/A�S���j���Z���		7T=���l����|��j䪜KQ�4T���ϥF*9+۞��rlj/ާz�VT�W��תMU�,�������?}�焭YL�R�.�&J0�^��qҼ�>s�U\rDD'}�14�T�7s_ˇ�t)�;=̧�uez�=�2�M���4���>&��H��ؽ�jh����#tb�z���n��<�vUWf�x>�Cumݴ]�=�=�%s^��E����w�%e��M�O4��%�����𼷴ѫ�,u�5کwv-�B9�K3���������M�b˷��q�"���*�'�Kߺ�΀�/L�����W��ظul&�q��t;uAQΞFTL=��xu�,;�-��HM��:�X�|*"����@�xWvHt�oV��}�%�d��/FU��Q|����|Z�3�;;9$�bƮ��YS�=�(A9tU��˗1�6wA7+s�V����<;�]���=����8;^v�ֺM�ƂY�SdG��٣q�AWrs8��η4V:b,����2�,��A1Q��@e�S�54���h[�/ q���"h�bQ��3q��sbѲ��XMf��R��EaMf��̮y��H�ĳiLm����=_~�֔��_[מ~Ϲ��<ؚ�5��cvD���-��H���anF�b�ۓ��I�����=�QB��=�nU��9J���dVMn`/w���i{���[�L����_Զ�.|��sy�����:`��3�w�W��8Q~���(
������2�G��!��i�2���z��Y{����n���j��2�������o-�f&�B��m��{QQ.��>E���ֈ�����-���5UUG��ۻ澇����5x	[�R���X혀�˻ɼv�RAn��#�	�(0xv��c�a���6M�XH(��B�l�g����bl�ns�摙�~�_^�z�8�z�U���?���aT���ݼM�ڄ{��.�3�]7���P����(ml�}W6m��A���1W?X�z�y�p�>���Xq��ኦ y/d��'h��zgC�)��g���$���oV���_�5��<d§�>E�ywk��Oш�H��p�T�������e��r� �W��ނq�QY���X�f*���UQh�|#%ĸ�������;��ڞ�~��7b����ݞ��e+�ʯ?[���P���U�W�>��,΁����o�z��x�1O�2/FܻtmW��l���9�"HL��B���n��q�\gz���!]+6�U�*H�c+����>z|�U�Kw�\�`�wآ�;'��QF�c6�U-�*��U&@/Y�>�]�j����\����z�w|���˞�n�eU
x�;������:��\C�l./ɮ�r��F���d�5�+2/F�}z�拎uƘ���r�ݩ�齙�:Y-������Mz��[1q핋/	dɓ&M�`f�$o<�ixx��U�1��r�s�v�UK=��c@�`�냲MV쉥}��k�s��QY���~挱�:�Wn�]k��N�H
�z�s�nהC��t��hә�~�\�p�C�UP��(�����^}���iq���;F�d�v�h�94�GQ][�E��<��i�#�]N��1�U
��]�����{`����}[�;� <t߃U!�N���4�>n��Ty@��m��ٮk�.}����s�USqW��%�������$|�_ؚ%��,m��.лN��ݧ8�O~) ?�5���7/���߇I�����lo\���Qݍ���CB�߮��||��l%\=�&-O@��|f�A�s��B��a7�]�$�OU>	�վ��i��p��e_]�në�R���zR�5��Τ^�:.��f�T��f�&n�}��erlϲ�q������,RJ73B���:$��󳳰q�z����^aT�UUV��/���>�v����^��b�e�r������?�������z1`_�f4\� ��ݹx�+۲���  ��T��RI$�Y��U���U>�L��{sj,wc蘻�˞�~�>��{�h}@���U*�UFX=+��9�>�:"��븜�;��v�Oz�	��ĵ}n�����Ҿ�6s��UOTr�f�):�s� Uzg�PW�F/;g���7�����N�fu�=|�s��_�~���{`��2�;g�:��{ �Ly���x��U8�v���:=�i�]��(ʍ����~�Gކ�M��*���������z�!{W�t�=�Rf��]|�V)��mt�2�S\�/:�tv��H:���Nwv]`�3Z%��0*���a>�+�œ|dɝ��<N�G���-LEUi%���F�롔���C���8���;�v�_�'�c� n6�؍�\��x�ݭ�D���ze�	��!���hY��b���M#YKq<x{#LϬ��y$��Ɍf\�B]���95��++\���:S��kU��q��7�p�<W{xiU�ر�W�pm�g�W�����m���cl��~���C�m烶��O�~���<-E�˭�0i���w9rr>ШRvxZ� �]�BP�\�	�+�~Jgc�n.���B��E.���F/;g����L�� ���$�.3W5fE�av�1ƭ��!�lOSh�ʡi�ۉ�ݮe��s��ػuwzf��Uڇz�G�|@v��I.�$�����`}�������=�9=�L&ŷy���ֻ�<�o��aZۛ�@{�mk��U 2�������b�y��\@�R/��a�R����vH
�Ut��)Dq����v�tn�>�|���:��UOU~������дiˤ���7M4ջ�	�B	��j�Ƥ*���lk���'S����
�©
�s1��혧��'����oY��Fu��>Rj�*��U&�4n#�4p2||��P��P>�V �Р�[����yB�[���p�2L.�i4en�zM��	U�0��Vֽ�`=N,��;;|ɓ �F|������_>��/�x�����q��b�tY�2����%���Z����Hsw�B�|����($6�މ�w�^}��s�é7r��aT��ۧ�]�������yUS����l�zV�8�<�wxD�=Ϸ0.���MIUUW����ː�K`��v���\��/\E�l�	�v�PUe*��￼���>7�1��Y���˭��jx.�����5$#��&�z�F�=�-��^�鱽�)��k��������_�bw86k���v��U;�����4O�nzDBiڦ�cc��/^���N,x3���8�z���o5m�-ۀ'1�Z��r�]k��x-0;���}�+^�M=/Z^y�ɴ���ꄑX��
,Q��Z��i��vDvR�+,Җr��i�/�����~�<Y2g��H7)����ys�\E�l��8��M-F���83�=�V�\�؛��^����ZSק�s��R�W�l�B��p6�RT�����qX�����tzｒ�4������8�R�k&_�O�y��d�B\B�3A,��%�9�AfU�����sf/l� ��wpڀ��{�{�:�'������E�;k���V�&��&��u8k�;]�ݠ,E����#���zq�B��T��:/8��y�87Z���j1�����t+	�p�H
����u��/�}릘Ow^���^���&<�m��av��}�<��S��=�܆W8�Sy�<��N2���-���x������W���Z�q滬	h�sy�}䀭��n�y�L���r�S�f�u���y�V>����۫�r��D��v�?��B�5$*�@T����0L�3���y����窪�9���~���kY�s^����\ں���M<����Tr^�2�y.%y(�t����RA��.p���;��BK�,������bS�<�����]�z��T�=V)�ט�^֑��L�]�`�3�b�9��B��
�-R<�O����Y9����gO;�{V@�����=��߯�W�����n�2I3�~��ק��^�n����p�q6��;�u0��vk�vf�UH�k�w�^�\{�iM&j�w���zf|+�z�9z�CW�l���&O�kp��"��x��2B~94��4�;�зvV@�^Oh�� ���U���np=F�9���/(�y�3�P���ɂ�0S���}Kݼw®����V;z����5�im8̕���GQ%�4��U8d�5f�0��EL�|vJ���]6��b��dhǽ�#�d�s-.�;�kS:�����}ב�8;���#�����Z����r����Zi��o�ck	O�{}�z���k�n�[�B���`y�z/�͞G�_�+�{$]ۑ�2�im�r5��ت2M��cA��e��q����:T��!��%�o��m��������][R���y;���ZRA�C�������fypo�v9t��[Ψ8��w9�/jT�u�j��`����*]�}��25�^��L����
?��X���V|������;pN2郢�nޫ�J��e��1�𬻻=��]<a�1�G�\U	-]1\�)[
�)\�����0%�j�.�/h>�k5
������S�tR(vw������(uѭ�`M~�%�p?Y�0ok](���ǳK=�2z����o�����*��V��^�"��n�nyN����st��Osl7�0K����nue���nZ#�ąQ�}ƴfwq�d�F[y1-]��9����2s��{��x;@�ͫ�3M�$x12pn���,r]x:�����49�!��]���%�۠���:�(ռw*���-��$	��P�t�$�<F�mD1Y�5ym��V=yqU�A �F�,�TՊ ��������E&��tӻ�\�-�c24j�I�P�%�R,$ vƛzx��Ǐ�4�8�ݻv�ۏ�Ƿ$���`M&���۔D��P"k��u�ԁuC$&U"I<i��Nޟ{q�8�8�۷nݸ��dj���L�\���fE�.>.�w2��6b���j-Ǻ�Iywv��N.lS
��1�.N���Wz�3�B(�wR�7�������i#x�	�BA'�l���g�W�{ם�CˌS�;��5��"w]�`���uo;+�ݯ+�Iwrg4W"����*d`��I^W1��@FC�%	���yћ~9��r$�~w~�h���~72S�� ";�E33���d���r�)9q�t�!(�s��ܮ�	�����(������~u����_����F13�&D&a�Ӝ�͂M��1{�&�1>w1a2�ws�u�m%���Lh�+�<���C.�q��s^n>k����t1�,�`̫�ߛ��?��+]pn.��;�w�?�~	�u��	I��m)�mZ+c���ev�k֝�<X�m&���Է眔�L��q#Y�G��cS۱����V�v�,�v#@�P�nۖ5�u������`���Zw`Q�2����=��O�F�Ҡ��i�Z�Gq�J���[�K	�f�@��s���{!�qÝ����jh�q��g�,�&@�焓��Gf�%�m0*�Tn�w2lW�gt�ݎu��.���a�����+\ˢ�!��yv���]��k��*��Y� �ܴ��F���#dK���i�Z%m%tц+���[�h7h{�]��R�Ws�Gh�S��3e������'c��5C��a:[Nk�+к���u��#XǡVֱ��[(�5�l��� \X�v�PmI��-N�bMM�nЋ���r��p��^uș��P6���� ���Ss�b�b��cu��>6름���']1��RW4ፁke���l;'n�`��h�<��3�Y��5�<+3��s�e�Yه,/`�v웷K�%�a��K�j�nۗ��k�6�vhMU�^̘fuMl�2�2�U��-ڹF����e�t��m��N�u��NdX�D�n�:8ON�V�ݏf����C�R���A�1�b�Yc����v�<�wM��v�;�nt�n��4s]nۚ�q��m1 �DҔ�R[QŃ3���y�r@�5���i����X6�X�j�\t��nf�x礎�vu�;�T�4��b��q�Am�ٝ�0��q�t7o]3AP�\�׬�	a�Zu��x��ʺnf������	F�9��Of8;=]���:��č��,籴Y�h��[���$�L��φ�3b*�ܠ�2���юs��������-��u�C�����[\�v��խ���c��\a;l��ۃ<���kj�i�j�mE�Ib49#����S����twXDSzc��͘�_~��(��-9,�aǬw�>Yn5j�_A}צxu�)�q�f�Ý���}�~���Z���}�V.b�%"�!�ˉhc��:��yi�����3�qI�U��[�7g����ځ��eل��ӵ�\�Q�^[��{�h��k��t��@E:��XT	M�ښA�r�R;<��ӵ�a7d瑆��H]b�a�G�b��&�l�K�i�8�GR�㶋�D��Ѫ!Y�6+&���4��+�:��w��J���L8������w��ߋ����)v�6F�Zm�2�6�r��](=��vن�<�==�}��6�{�O~�я�G���6gp�W<h��6u�/�n��/6]�v�g�pG�fMmdEgV���V���1&�7�#��L&|�L�_Ǹ�uY���US�X��n����˅Q�2E��|��5
k)���܈������K>wW��CjJ�г��e���M�c=�2JO��x��q�2�4W�Uy3�k�����A���ޞ���{�#��L-���
��ZW�^�������inf0��a���6N7q����5h�V��.H����Du�r���&W�������!Q~����!_�1cx�t��;bBe	P����Ծ��*�Y���_-�5`��lӬ�������n���ă�.vb��ދ�V�lV���s+y��al.��o��2glT=�k���O�e���F毐�'>�3�=xJ�ܮ�@�'�_L�f�f����y&P��X���[���a3o)���F�������]�+Ah�ɦW�������!^�g&����0f��׀�|�;S{��D���0&:��}�ޡ
�޵YF;De��oZkm�I�U��c�J�߸ǃ��r(r��4)���7�蓲�	z�5�m5b��5��|��I6fbg��V�zMxN�'/B`�e�VG�(�Ѹ�S�.&W	ڵ��v�2"2��Se�uY�˟/����:E6��T��_!U�n���j3ʷc�P�30&o�t�}O�TĽVz�������r��74Ƹq؅u-Z�u7g�.m1��-��}Ĉ��g�鬮nuk��(s%���ˀ>���@*$����>�}�r^���uU &S*��=��T)/��v{Si����|����jD�s5��'
b��c!zϹ� Խ*ک٪�5HL�xv[�wluƯ;>y����y����/;o�a���R�4?r!����!�E%ڴ��Zь͔�W�Τ�#,R�Y{JX��]��>���4Zm�MT�Rط�׶}� �Qɾ� �ܛ;��~,C�v�C93L�ڤ���R2��y���[�}�6��UH��Ng4�yL�Z���'���4B��q`jf�L����߽�Ĭ��U�U�o!c��^v�	������Bi�^�j><��wn����m��D�Y7�&��lNڟ��M��/��|�Z8+$
7�v2#s�`Cp��۩$��`u��8��Kgv��NT����c����{��Y2_�M�q��`	�2�`g��'�2�fP��f�?��P��Nf��@g)��9Ât�}���=��yCՅ�R�XQ�qmW��W���&+kwhVQ�4m�d�e	�=�c$m��O���z��s=Y��r��R�N�Hf�ԣxY�SK���r_;�ћe�q]�����ܟos��~B�7�0���3/{t=�:�T4e����I��X4�	���e�B���]s��U��~v7��owX�z�b���j��v�n��]w��&S;2�amV��y�z2��Y~��#(�MwM�7f`;L��9¸עg�,b�Nn���Y}��w4�3t�zg=�V.#�к��:��777p�d�q�X���7E�4a�����>�ͧp���1bɼ��ty=�_B}��|H�ո�&!�ke�lݰ�$,�9t H��6�^6Lk��C�x�oBq6�׬�{k�ukGg�0�g^ֹ�nC]����u��9��nE��h�_Re�<%�1k{Gm@�o]v��r�Mk�^г����VǏ����"���k��I��:z�kc4��g��i�m��޵r<�r%��#�K�30�Wm�П=;}���J젩z��ꑞZ�a�H���l�`+4���o<>��^��f�c�xH�И(	�<E�_MK�%�J}S(	�/n��<�z����h�٘�w�T�i��ۿWޑS�^f�]Z<�k\wMgX�z�b���	���wWy�ӽu�O�hF�6�L�i�ŧ�f1u��s��	w	޽Y=7�[�`��B��Zݙ��2H&c����m�n��A7c�����hǚOB�p9���'�+$D�p�C�|[>�f��J�8/�B/:�7�ο^-X���;o��0�rI��aG�����=JJ}/1�R�smY�E3����\qc�Yϣv:��p����d�@��*f[�އͯ{�[VMw\Nb��`N��n�ٳ32-���i���u���f�	k�[���2q���e�	�auu�{�_�K.����Ggo��-��09��խ�a/T�����N��J�+Eb5e
���/^�W�̓&A����S iNn�{F<Ҙ5�s5�W.j��S��P��t�u\��P*e	�5ә�m}��6ັ7kV)/���P�W)�33��4��<^h
˻^��������~�T�'�=9]y���?	��S)�SL���E_R�lc{V^uE���R滉9��b�&P5��cJ]����߿Ј�t܎��o���b�[5K�(�T���Н�F �����>B�L����ܑ�{�%+՝��Ӿ�.�,
�l4��4����)ℿ�t�׏^ޘ}��K�`�ʦ�@&ݙ1�3$�KlDkA��@L��L�2����C�f$���׳kmK���>�O��wwϬ�d67O��KC�J>#�f@͸�2	{xnR�?��d�2k�A�	�}'˩K��$�|&|���Z���`��vr�OF�@�@g)�2v�W��1)^���7�,��u���Z�S0�I@L��ѓ>�ȅ�����n���z/%ke�ʮ�7Hk�U!3���+���Z<�,r�'I?����B�/����l�X�=��ֽ�s���3$��d���{��iU&$4�k����1�F^��'��\ꑛ��W{-���|��5Ri�2�^�A�Zj�(����LZ�r�q��z2�Vv����Ux��w]dz��!Z��TSU8-$c�����/i�� �3�՛ϐ���U��n�gHUK84PǾq����}�M�2�۸�����%
� +>�#��u�d��Y֮^觠��YZ�O[�ޱԳ2ͮ{�P��4�N�6��wu����nE�oh�Ϣ���ƺpu������s6�%�*
�#vСW�Ks-�խ@f��`	�L�7�ʥ����yh�6hD��p�^QY�}���ꗤ���b���d�<��D�HX������Jd��%<: ������a���;�=y��{��r�e[_p��F����;�̰�n�ެ�(7u�����+gufU���bS���u:�(��$��֟&��i�*��{�F�3d��t�bf�S*d�ۣ��ѥ3�$�!Vr�������d!]32�ʍ���f�B}�`� Ɓ��L�~��sӢ1J˪g���ss������([U8�B�c�������<1�>Szw��+��9z=��ު���vP�J��Q���z<,�9d���S/qc�nK��Pܡ�L�2��=��k��EZ��(��aqĳ#�g�ٙ�7߼<=���k��ߚN���'�1�@\��Hh�lݓS���EX��B��RaF�%�����	rGI���6��i�@M��I��c:lY����PJb�/���f��f���&,�&ұ&3���:;���I��,6�1��4�1�GAu��S�� ��*j��{;��ù; ex�<{T烫a�c�@����Q�����?M`�7�XR̢o�Հ�`I|k�:�
�AZ�+f�q�j�Z��HJ��K�k.B�ITͺ��@��� �M��e	�u����0��՝��ލۍF��-��1T��g��D���7��F�Y���ђ��껚m0톙���i|���<��k��M��7_�lݩ�����^O��|rr��K_8�B�4�g����7��zP��i������9�����<��ϵ�����C��Z������m�����^��gϙR��lo�v��Ͱ�������ή(��F-�RW����mT�J�(yz�*��H?��L;冣-�T�2l]hK�v	��>��/B����zP(D˳�c��+�=V]�\�Z�����FUӎ�~4�V��8�O`�Su�-���'i'��������`ϔ��P|��\�B��ޱA����}���5|����q��a���ŷ��R����,��B�۹U*�qUo�'#�#�{���:�F��Uw8��L�2�fb6�V�˧����v��%�!4�i�g/D��M�wm0� ���{�9���B�[U��Ɗ.��_?uz�_�ټ��b���d&��&P�^�����y��Ʒרz���Ŗm*ZT	�X�b��YW��j�!hI#��(p��� �y�A~��*�w\�k�N��싪�LA��oB�M8�:�{T�i�����5T�'���i�g/���M�9Z=al�Uo�B�d�G�����zv��T�U@ӏ���<�ϒ�����}:f�zB#����=�2�v�M(WT'��"�楆�R����]q^gx�A}���݂P��fu���m�X;��W7�_Q�W�u+{ݖ�FRљ��g��eu>�?_����l�I�[Y�F����,�<��5�y.��Œ��n�2�~cܞ5���6�,n���ޥWc��,��b�i�//�e��|���^A9�iH�t���[.�w(�;�5�G-m����˵$+����]t�_�!#�)N7�����<HŤ]�\�H�oix"����V���;1*�*Ӳv�n���`���Tj��S�Gr�P��77""��]i:n5��:os����+�i��훺'\�Y�F]<��w��+�Cbb\� ov���_]���Ɗk��̫��$:����s����8_v^��)Pٸ��n�{d�� :�d��w���6{b���7�btz��֊�c'J��^�tgr���O���1��]�ʙ}¹�H��ُH�]�@H�OE������0�5���2|sW�c�l�dŶH̭��#4��D0om���2I�t|*rכ��l���uR��ˣw�;z�5��5c0�z1��ۡ4�t;���"�jX��]w0��o/�����mZ��f��
�Y��ޥ6�`�4;2����܇3#��YN�,5e��3v�ֈ�{��<>��V��=�-�W����x�!꽺��E��V�� �jE���v�]�I}�h[Fs&�*9-��t�&�u��\�-�1��ʹ<�nӴGfl噳�:�+EV���2��6�Þ�������I���ӫ[]KG
�N7[�|������޹_]5�|��!9r/񻧻guDbLww�����央\�� �����=;x��Ƿ�8�ݻv�ۛ������QA�Q��r�_�na˱�w@0�˻H��cF��s�yW��$�=�ۧ�o�q�q۷nݻqǾA�TI*����P���>k�@�9��oϕ��	g�m�]��ҹssd��1QK����r�[�L@��A�s&�_;����A_n�����tss
�(�dSI�bL��_Z=�LQE��`)(�wg��{�\���&B4��Wu�S�r^��׽���&�1QI�H���b�;$Ѳ$>u�I|\�w!��L�/ͷ]�u��]�%�u�D�E$����sd�(^���z����fNX�M��m��n�Ĕ`�f�I�LhK�	2TnV�3b�93η���t�͗74j(3�r�L�$I�`|��X���p�=�p��Wo���$|�e	��Ы�^
4V��a�q��m!Q��F�t��^��Wpi������na^�fѤ!2�P��&W::�hy�̀���=��sD�DM�9Z�Ѕ�L&]X�%�S�����!I�_�ܸp�/)Q��a��C�t�f.�<��6��*"
�Ov� N�'j�	�m���ox��ݾc��P}Q�t>��(L�2��"�*X��G�"��cz:te���Wp��%�Z���v����m��j�0����5W��PY��	X��u\뼃�߽���.�6i��5N�ܒIx�����B��8��!�1׻}�k%Z-x �?��=����7�N(nY�r����X�C^RQe�`+qE���jWu��K�����"]%��������l�|�ɦz�RMUQ6ΰ�G���Z~�2�����K��]�kꙉ���j�X="�MS�C���>�+#���[3C{>ݒ� 7C��OO\VR�{ki�إ
^fI/
/�5�l��5R/4��˭���9Z��Ĺ�˶�v�F���Be3��7����y�])�W�<�g��1׾m���3��/|��\3�����<���M2���B���(`�}�ӣ-N_���E�������Ww������ڛ��7�	�<+4�^˧���g4zW�Z�/�=��y����)0�L&y����7�[��������vtڸ�#��^�i�2Su���N��e���D�����ɳtԭ���ۣZ T;l�S[�T�l�=�0Ve�M��Ƀ7�*R��2����ْf<��,>���|��@�ߏ������4�֣��[�l])����潑����uxꐠk�sL[�"]�-��У��u�ܔd��#��6K���u�F�,�ca�Ƌq���%A/pjw^��;� ۱���Nj�v+l��g��rl�i�{]G�78�w����nOH'�/c��y'��̘��G���!t�+�������͚���-0���V1b*_��6	�D+�4��څЕ�čӕ�`�i6�v�2�	��u����'>��fe=��{��:2������f����{�I%�!������z��L�&P]>���t����ePsM��:}W(G+Y�Ѐ�e�7U�����C�,�s|��zSL�2r^�=�v�6	8�z�b��o#{݉�%5t�UO�v�^��R��X�B3�M���A��ܺpe���xWpoB��f]�cܝ�6��v�Aک�bG���һ����g���7��	���7]>�熺ϛ5����(�[8�{����Z�clĴ���gnme�Uɺ��A����뢝��('/L(��)L�c2�Q;;<��sH]��|�ۜ�<���N�wܳq�RHh=�� ��u�u�X|b`.��bN��r���z{i���[~� ���f'}�7Q��n�-
��y��j�`:�D\����|(@ <XCs-�(��O�~������Wy���dۯ2����`y�l&�33��J�>���Q7��_T(�ɲ�Nkz��	�Ž.�n����f}&O^��]��P�;ٶ��I<�����f�S�_�՚&�HL�(>i)�S������ѾY�ڜ��:2��z��5�
mתB�j�;�L�/7���JWż737k@u���F;d��N4��Vu�d�p b�E���N!©ت��-�;��v�#�&�@�p���FщB3#�ɚ� � L�,fPg�9���{j���ʅGh�����׈;���Ex%�7��G%��>�T��-��µٺX�c�S����Ԇ��YY}�[���I�)y3z�7�o/VVO�t�V�2Q���v�g%Xu�USw����X��^�����������ބ@$��z�&V���_Z�T���2������x~~��q���B�=��U0nT�|ɜe!T�ԇ��S/��G\H�B#�+��g�O�����5j(4�R����ϳ�#*
�<�QZ�c	�cQaa�X��a���c�*�,5��$�ul��)�Py[;�te+���ǿo�bus7Y��b$�)ۭ5T4ϘdS������}��C%N�����C��Y�:�G�nɚXN��U�i�um��M2��lU#^�vv%��G�@��+O7[��x���q�CZ�3��N*�O�v�K���&=v��xH=P;��Q�]��td�����hfe���'���s:f��O���3�p���;v+O�k���.��Hl�w�J����6��d��לI{�^,E�-�X��p50�S &i�ʙ���I�/t'�Vo�b.�p�l�f�MئP���r�[<��s����K�E΍�:)Mi6a�fԄ�H�R�PK:hw��+��!bf30&�nV�y{GHSY�|�%�P��m�k�l�2�e4�g���S�7�ᢜtE�f�Wђ�����E����^�%���?��=a��!����T��k\��w�e��|2VR+�v��ʂD�߲s�7�BCe���`��e4ʜœ9���঳w:Zm���3�|�1C�p���h6��G�f�>l�9H�+>�3幽�MџV��__��m��4�w�/�Y:�Gz��7�49,��_AP�mua6��ňab��V-k㛼���)���MNnl��z�5�0iP��Y�����oI�6��t�c�՘>yH%XEˡ*�a	�u�浬��j�ؑ�줣b޻��70Q��b��t+ŝz���Μ�Eڳ�#�֤A[��+���Z�؎�Ô�c��h�,�N����,��XbnֶĂ�/	����&p͸f�%�Q�s.v6�)��5qs� �\��z��v�W�f����ns���%�#��l{��h����~Z�燿{�ZC{&!�?�7X������엣�=Wl�\B�t�E#BH�
L����LD���L&}ܴ?�5:�x>�6j|o蕌3��|�3�&��u����*D��3�)�Y3�:=�`����7P �qUo���|z�M�U���L��e4�b�TMf҉n$�te��`�+���s_���3$���;�M�7t�<�	����sS���ǃE�45B`��A1Y�.���ڭ5]��T��j�gO������I�P��Ub#7��7w�-35t�0�q�9��O��$��q��J]Bjv::uk��"t6*]@��<;����[�S=!2�1I����M�����\��i�����Pi��؃�3 H&b�{��z�F���Tzx?-��{O��q�6 ��e���_v�6��k͚.�@���)��.�䌒���)�4꩹���\����^�/��r�5�y�虡�#�����!�cݻs2���2��f�����V���DnrD�f��V X��g(	�3L��\%�su�U����Z}�����]�E�y�Q�'�;�p�6ҙA�e ��S�R��"��}�@$K>!�N�����ja��>�D�r���T܉g��6V��B-D\9f�${X�7#KM�n���~��-�C!4ʙS��Z=ܐ5Y�����,�t�{��ƺ�����gq�"���X�[�K:��h�+zˠ;�m�Bg����~��ɷP�S)����
���s���s�2�����Xo��*��..!�'iu�	��a��d˸Hս�;����is����D�����i�J�z����� L&��J������K��YuK���6F�Ǿ�S��ȃU�cw�S1�H-�Mw�[[%������U]��ϛ+tꩌ<��I�>�2��.����@L��/�C�-�O
�� �:,١�\ePI��[��(�=F�޲���:�Qp�Z{��P��϶����'�c��+�A��s���l'�b(kU;
�3��&;�+��;����Q���U���dئ �MU��[w�y����r6�B�s]ٗ���&<��g�5~˸�3)]e�p�A�e����(L��/����8M��<�e0�S֖���_�=���h�!-5�)�ndЉw�ۘ�~�l�׷O����Vح\��C��/zܲ�봦�:X�Y]P�q
���˾Y{2j�t��7��!^?�DKs-\���u �HL��R�ًs�T����jMX��\�f+��&��t�y��S���M����߳G^�n�B2�j�5�[1�ͱm	!z��8�ce��w�������~M-X�T��@naɝ΍���]w�{Ub�Sq~�+����̳�(	�5:��wDMg5�*��yih��t����2u��\X��T�Q&�&DI�Ie�C-	�2�Α}�>�=�z�&��m�* �����+�UݬE���bM:�~��i��R������:��O���z4O���]wU��'*Ϳ'�뽰2���*�j��Z���8�y�y�>��tz�],���װo�Z�a4����!��f��H�*�+_�QQ�����( �lDU����""%㳪��Wem2����ke��e�Y[,��UK5��T�[++e�T��,��5R�l��Y��ke��Y��ke�R�l�[,��[e��el��Vke�R�l��Y[,��[e��ejY�����T�j�ke��f�YU,��Z�5��U,��+e��f�YU,��5���eT��K5��l�[,��j��R�l��,���l�[,��UK-��l�m�UK5��l���*����l��,��j���el�U+*��R�l��YU,ڥ�R�X0V:��C��A� 	f�YU,�K5���f�Y��kee�YU,�e��f�Y��[e�R�Yf�Vke�R�l��,��ke�R�l��,��ͶY��[e��e�Y��V�-��l�[-��ʩf�Y��ke�T�[,��-���eT�f�Y��[e��f�,��6��l��,����f�"���b��؁C!�ie��m+*�8[]e���Y��m��e���h1R c��F�E�E�E�E��E�E�E�E� ��mTX1X0TX0X1AX��`�Q`�Ec#�U�Z��VV5m�UU1�UL�[UK6�l�fkUL�ժ��ګ���S*�K-UL�V�Ymj��V�,�U2���l�mj�2ڥ���k�+R�ZYV�Z����##`�X1V3T��X6�l�"���
��啲ʩe�Y��ջU,��6�e�Y��UK5��E����������AAT1�O��+�����?_�>g��83������O�<����(�������'��O���G�����~��������������i _������ρ�@�ҟ�/�O�>O��
������}���贋^��ڜ�� �ȝ�
�����Q'ԑ���H ��"����H*�*,�
�*���
��R�E� "��, �X�,X ����H �@���B"�`��@�����T���B�b(��
� +*,����D`�"������5�*�[&�-�����������}�4��"�����   �3�>#��??���	������>�??��"*�+a�(>�F���������i������&ϩ=����4?:}ޛ�'   ��EU��Y���vh�PU�F�  *�
O��%���lc���{�h��e��F� h�j*�������Z��ޔUQ_�;<O�tNq�0��~�����X~�>!��0`pk�ETW������QUEv�9�C��)u�'>�%�i�h>�����`zN��Rw��EU�>��+$�c�ᴤ�4˸���}�����AT_�t�������?�g��}?��������(+$�k/+� ~Y0
 ��d��B��                                     �
�      P �       �         (          �Ԕ�H��UQR���RUBUJ�J�����$U	 �	% �(����A�RTD���D��  P�Q"�!UPP���>@#@vꔐs��P��y*�9wp �@P9�t ;�� 3���A�� +��Р  =�   ��}�k7��B�������: �·�  ���:4�`t[�U�ޤLz+����$dh
-�t�
��
    �  ;В(�QJT�$R�pFv�	��:6���R�t�z�=�СCw��JU�` �s��R$�R�\�� W  P �  �/@�־� �B�ޱ����օ������z{ޯi��I���p��qںc�c���`�   P>   �<�E"���Q 
�"�>��4כB�6TYe +{9 gB���F�� 3� 2��
�����    4�   }�����"�� 	 X��p�UD��$uA]� Gb���@   �   <<��R�Q*JJ��!)Uޡ[��T��+  ��U�(�c���l Y�@݀b��*S��]�{Ҡ ��   �;ϸ:����JNt�.t��!��Y�TT�MJ��Ҫ��Ԉ�J�[�Ԥ*�4�K���G��:�U@   �  �Ԓ%UAT*�TIUR�JCL�@w� G  �r�R�tvq ����� {�J� �r@N�  
�(�  �>@� 1� � ;�� �W =� �7` �$��os� �`8��`#s ���51��P��T�42JR�  ��U IJ� � �d�&$�   J~�%SD����d	53JR�� d<S��������ҷ�����$������ک�l0�=~9Er�m��!NQ���@��D�HI	�B!$��!O�!�  I!!����ת����V������ۻ+~�I����ǹ��:5�D��3��T�?�m'��z�ʤ�	pm����ȕ�P�6�SfզeCn����0�zk�}c�82�`�/t��v����-m�B4�ձ������[b�
h+Uza�X��Ì5�ʫ��ýv����&�&�Wc&�v&$Y�yxkiL��V�B����[[[���h�̔�"t��"�Gn�:�E���x6c;YU�P6�ۊ�8q�T��yZ`b���)x��������Q��uV�V�ѯ)Ę��J�6��"YZ����O>�%U��É�Զ�u��M�[y�E�"��gnR���L��`e
�d4(���r�Ie�ٹqۢ�S:3L�U���A@�Ec���j�M"K��o#�1�u�����,1[ou�p�{ckH�1��V<�0���b^��%^AVjI�ĺ����T���&᪼;�A�6��Be
�4���l�f�+��3�Z�+i�YZ�k?��"��D��4+� ͽ��+;m�JF��(ㆈq���dmES4�VB駻d��XB�e�A�ݼ�4:d�2�ۺ6l[ܣ1�m�uŏP[��kl;ݹ��̀�T��eVX+^T7b�2]M��m�w/k(��{�i�]�Yt����Y�H���m�M��"?��J��*KM���͜�v�[��P�J{������rQ�Z̅}l4p�j�����l�\Fu�V0lŸ�M7�wi�kln�u��mG3��"���y��IH�V��1[bk�[�U�ٻ	�n��r��q^�u�J��Y���p�k�Ӭ�Ӫ��P�S�ղ����]�ZӢ�KɈ�.L٪��!��C�Z8d�%���`��Yy��\i_Yʽ`�3M�y
b�θ��T����%��<�sj@�`3	�_]�obg/i&1���j�A*D�}��F�܁l!�c�����
�����/l�0�]����TǗ��A9[����Z�W�l�ƅ��o]7H]ڿ��t��/��,�,����@�Ӵ�n�[p+�����f�rQy��:��진��#V-��3/Z�V%Y���6��iTW�ۙ+��n�Bkm]�]謋oopAO�V)�giʻ�j���e���Z�^ޕb�r^D)hw)#�s�l�Ú�V���.��Kg*�P+Zv�HQѳQL�X�ȜGj�qͽ����2욲anc�@�Ȏ������fdٳ1�&��lj�p�{��$�0�_l�x���Ij�Z��J�f�6�^�wWhk���
7/kY��Sc̤WTZ��Uk��'J����0qުGs.�Fb��P�Y���5���YV�faK9�ѬA���e�LG��5�V��>����%e�F�nJܫm��f�i�L�^�f_�֣:�㵥(ZUr�.�p�|�H��7y�^%�UmfՅ2���ܑQ�����Zo�:�*�US�@:��o��:&�b�T�i S�ɚX�T���$^F=�`Ҭۚ"t�Yr��v��`�nQ4�ɬԔwo-]�舭��iƶ8�Q�񘢧E*YoT�㛧Z#&P�q�M:������]<�2b�6��)��T
�v�J�2��W�YY�@,�lc:2�L���y�*�4҅r�e�^sQR�2���F摛��b��v�M����ġ��W��J)��Ƒ�t�bM�黬�Ot��dE�F����qn����k�&�zI�wR�u/#�/�He�̺9���ڔ��e�2���P���n��ú��!�<��3�)�e�C��V*L��6]�呦]fJ��èm8mK����f'ܽ���[�vu�7�z]�������[x��G N�Ţ�tm"�5�<�����!ƍ7.��}LV�$U��G>GL�ӛ*ط�hʬ��L�ܱX2(�V7JU���I\{c5�:ݺ��;5�5�oFsq� ���&�������]�qř�i%=����d�՛���	��5B���:J]jQ$fcV,b�X(�R,�yye\q7rL�/˦U�(��N�ڻ�sinQZw���M��j����� ܻͬ�k\'
����Qȥ�b�㬋J͊Q�W�裖Z�!P����ؖ㸝��HySv��ږ6ѧj�C�7Ù�{ygT��^3���C��H��޺s+3lS�,��H��ں6����pi՛b�Ŗ���Go/l)�[ZK�p�����
���PGV&(^X���om�R�e7�f8����vvBb�4޽yJBɎ�A��ʪ�[3{v��,��5�V�Oq룥(	ƺ�5V��f�F�B�ձ�Բf����Y�"5CIzf&	���F�`�/�sVj!��wx�����*�|Ba�P�Be��K���֐����ذv��f=�aL��婧>uB�re���E]�D)y7M�j�R�V�̽�k2B���g]`P�6�P��W�^C.���b:�:��-뽩�A͌m�+�J�d5�5jͫs/^*Si��l*8L=Z�hf��7�i�@��܃H��V4�3��[�U�a	�f)WJ���U�h9���VAR݄_GW�����1^i�Z�u���
])/H�1�#�ͬSu��5/M�����5��8���9�J�^���L�nmmYr�f�ն�V��n7o*���]8�m��7	���E�fH�KRJ�n���KՒ��%ns}�B&݋2�l#h(�-�VjbK$4���h2�!�׸T��!�IGw��0k�Vf̗)Y�w�؇m�>�uY
iVh�ڧ��v���:�0�"��<k!�R�m�c�ݸ+CkE-�x��ǲ����M���Ә�Y�����c����e%��w�����Uw�[�@#xwg��-Ч�n+��j�Өk�VI�5c�nP{m�-���kM3�i�i�&0�ah���*�Y�NfP�Y2�.1�m5dF�Y�
��<;�0r͉�4�q���m̢�J˵�fZ�͍����S.��VolX�E+��p#h�(��M��[�G0��^涥nl�%���.ɗ/i�Mb괢�X���/,��U{��X�ӗGVm�f��U�P�e\oM�T3j��z
�Zj��V;�ܳ��Ճb�{W/
ݹ�=���7,��gq�jZ���q@�^��or�V9lEZ[����9��3V��C�@��c��o2d"�͢��nnf�Q����8��x�(j��b:7z/�)^ʪ�ueV�d����_�*U����4K�̘��O*��R�S4�z${V�am�đ�ާ7&j����I1��L*�Ɯ�o�
���ܽ���*u#mD�.��Sw(Q�9��������Ӭ�Fnkva�5=�j�>'sej��jRV�<��y�)Xm�f��K��4���͵��>��R��Om
t.7*@���N���5����UA��f�.�R�����1;Y6�n���=�FL���n��E䭭�Y�K��e��(2v�Z!��s7�5�֪�/a��ZD�����gHK��I��Zb"P�
��F�f�V��-�Tb�r�Wa�u���n
�R��ܐ�w+^��Fn�%cn2��@�ƌ�m-����c�I��X)�����!�bv�*�~��me;UY����QJPUV���U-ƎGg�4U^֢ͨ�j9&��tf���˩D��t�T��y�[9B�L�֪��-�c�w��I�ᒮ�ug�&dU�w����U!(`zR�"1<���,���YZ�8��:�+0@reU�UP��ڵ�����G2��ѫT�͚�+��K�*��<4���R���h�4�b8��v�5D�)K3IJ��o�Ō��:Iu��C7kv��[�D)��.G���rm'�-��Y���M�ʳO3[@��F�Y�@�W�cљV,n$!sn��+�Y�G�����Y~�s]�!aa�������q㧶U$6���(����I�)i���Q�uL�5��_��=�3���m�ꨜn�+u.f��'�Ŵ�^j�[C�mc(�ZC�*�h���R�&���:��U(��j?��o12mk�9J��i�KY��q�V6�Rìa#���T�ͥ��gr��y��U�O�Y.YֳseT��SYB�̦%�ә�6M�Ϩc������lɬc�NT��El��&��ݬu-��r��f��1b�Y�^d�v*��n`����u}W�뚥����C�/�\��Q�ojB�4c�,���[�p<��������ӕkoR�UOvhu3�l*��n�E6MR�k$�ʕv�mɹ�ȫ0�H�{����3��t]�u�{���E�����x�4�_�aFh��eJ('���WF٢�HXn���Ԙ���j�!��7i�.�R�,�r��t���t��j��U,#P����u*�ƙ��=Y�X\����Y�[ytUT�t5�B����j`�jG�N�M�+7sT��`��Opܙ.�l��6���9R����AQI܅�E��N�P��zD�R�ю��72���BYn�JMD��5�����R�[�D�UVC�]��ʊ)D-,��]�i���Ga���ޥ����������V�[Zcs�c��J�$��o�3T��tJ,�u��i����h���s.�T[4R�q�WoTW��ou���ySf˼ZL�)x�W� Y$���;��X��O!��L�
L]�0Te�V���m�[r��n�K��kUh1�_42�]�U��1�W6�X�D���{�!v�;�X����Po�5Om޹H�+~��Uhm�I{����&�#3(Ԍ]�f�x(^�9��ZkZK��d$ͺ8���V�UR���������6�SZ~ܔwo�swS�/&�L��#K�On�d���C���m[Pˡw���1��{���#G*�񺒐��ZP�-^�Q&"^iIc�+T�_f��j�������`���q�]cv,]]��v�{+���;2Wkʍ="�-�4e�1I�m��!]K�i��3u���Rm��o4��t�34"�eֹQo�! �I��6�`9X�anY�ӂY��Xd�Px�w�cR��U����׻W�HCgEa���.��鲦���}TQ`�NA���k���5����7W�iK��<[�+�ks׬̫�0�J�����*ӭ��yQn���r�!H�A��cn�Xll���f���a����$��5�]��S��ݑ����j��
ߵ1��<��M���;��W���H#���~�ɡ�*-ܗ��� �v�Vʴe����F�n�lʷ��oc���

uH �n�Ux��oot%��P�׿(��3#:/i�&<�R��Ƌ��U�x"7N�WB4��:t�7`�!ͥ�con���'r�j���MB��-��e��j;X�}Y.	t��
�8*�Ǝ��\o!���H%w�8H��b�-��M*���2)��7�(ҍ��X^p�w��u���v�q(woZC`&mTlm5*�2;�F��{K*�\�;6��B���C��Z��!4����ԥ�ev�J���&t�e���qk�����p�����S/D��n�)���f�����*���2]b@��F&me������w����GK���Iu�!�-�+� ���حgR�P-鬫�V�ּ�[	5�����[V���ފ�=KQ�#u[U:��T��2mYʶx2*���*Vڧv���:ts6�.�wu�S;Q=;3q �r��ɫ3h6�+r�v�1*�fԦ0�a��Z��a�Ӈ
���ǉ�D��4��3rc�����<١�Y�T�r����ݕ��d�d׵��CdVu%��j=�ff�wU�����߲�r���wr2����MU���F=�>i�������0�!_k����[���2AQYǖ2]�^��SuR�8�;�j�)��d���u6��w/qR8oiѼ뿪�%�S
*���Wx���ӗYC5
W0�#���f����b�/E��32�3�YH��h�h�f���ĩǵXҪ��]�E�{��f�
яZ���mn���y[K	�"�%c���\�H���fu:̝֍��{�z��sT�u��oT5���Ь��$Di�X�)ֽ�X��r�`ӥm����Ř��YW����8�$��f#/�w{�	����4��[n�2�Q�ꠘM3�(�fC�;
�Y��h���o)�2�pef��a�dͼ��*���#��3��zT�M@�2��-�� R�n�t��7i�֤%�����z�7��������ӵ���D���T��Rz��23�F�P�U)�G�7"�M����f36^�Ց2S
�J��Y���pV�Z��h���h�/c	M��V�S0��fV$�nGinIx���JT�8��{l��Eأ�a�5#fcn�{���yeeKQ�suM9��ܧ���[.�m����.�p�4����ܚf]��
1Xc�y���H��l��˖F�B	��J*ܫs����DjE=���4(��[O1"H�,�D�.�9�"ىc���ס�򛕘e@٦Իl�(f���3d����Zu��eR:�	��9N]��8]:Zs2U��a����i.^��{�����x�e�&H�vR:�oH7�p�OrA6�U�N%c+w(^�kQ7+��o:���sǮ�oy��r�d
�Z9W9�f�wn5"������&�Ȼ��6��%ԣN�e�����s���5��g1^M������ZH��L:�@��%��ǵ{I�j+�vvʬ1\�6���P^��gjf���B�n�H�E��yVp�{-M���z4:˗2���a��vݘ�U� 9W��G%]lZ�<����9�B��2�f��̭�N��/o4�
�����V!�+䪪���	���	joe�I?TD��7Miz�\uu{�qҚ~��dUr�dQ���\B�.�:֔��㼻����^bS�uN�9�n0f�j�r(u���Q[)n:���"�UfD�"��q�K)���u.w/nMAV���i]T�zއ��z��Wӽ9�������O$�N�;����J������� ���E� )E� �$��H)$��I$R �� B
 ��$@�!!$"�H��,$�P��`I �X@�I	 � �$��$��I@!
�:�㺣����+��$ ��`B @ �I	 ��"�"��X,!a �,H!�"�d"��Y@���H�$ ��(@RI"�)!$Y @Y @P�`P��Ad $	@!	"�� �d�(	�\u]QuwWU�Wu\WuD]�WQ�TUEu�wQ�qUtWQ��A� $���B!$�4�׷���f�?���`�-�ܛ�by��ܓr��9F6��"��wR`Jߘ��1a'�Q�FTG�ք����VP53����v��W�䭫z��&�[��N�r����²���Axs�[|�gmn�z���� �qԠg;��7
�ԖK�܊�ܭ�BK:M�8g�*��8*�)�N�Um��A~2���u��S^�(�k�v��8wN\/F@���(�]imniL,R��p�<��l	n�q[e��-N�)e��
���g-u!�t�sA�q'�ٛ�X����&f@��7Qp�LE��MO�۔��k#eeH�ޣ��N�7y)t��wI���Ʊo�L��Y��t��Ky���u��S~O����ǽ���NɕҁY�hui��S��s{���X����Pcͩtt�/�F�J�V=\���1t����X]ֲ��}�ʘ��t��6]�y���԰i�d=2���ͷS�]R;�.�6̺�]�D��9Z�$*��a|~L���j�Pf��\*�FTB��G�-��۬�U�K�N�D+zov��Cpm��;c�c�h�\j��^��{��1Yh�l��޼ƃ&
{�G0>������������v��5fg
8��M��p?#}.��Rs�����*�;L=��]t�����pI"W�b��`���I��yt+ZSss��}��s/�wX�g"�pjW�9�#Y�eUmvܵb�u��qsR�e����w���^��W�L��܇fY�T����{7(��Уpd렒6�T������&�]W@v�2��x5Z7|c�*�]��N��M���Mu]�^aé��'��ə"�'�$c]���m_R�3/1�T2��L��q9�u���K^�L�e��׵gk.���{$˔��W|�(��f��WOpc'mUD̚��6������W�|pY��u	"ڗA�DlR�]ży�;�k8c��Wvj�<un��tV-�z�x�:{l���Z�,�&]Vj�١���T�;�젹]�꬘o��ٝ2�z%��Ul���[e�n��ZHd�&�l-�O0�Sy�A����C�	���M��G�66<FmVQ�[�K:��|���Ժv����i�X$��i��F��mhjk��N�����!�'y�>����Z]����
dC�[w�,�8s�LV��y�Y4殼��k,;�E�oN|�^��lt�1�U��c��׃GSZ�ް���E�זN�}UD�v�Ɩι5�J���B��+%��B�^/����ꓝ��s5�t�^gv{�L��t�V��Y$��"-�a�%+�o�3[J�ֶ�n�3��y!�6�,�4�@��M��8M}�k��OU�Q,�	��[K@U�����&��M�s���+b�3.�A�x�a�e>���P�tE];�˧ٴ�B�>��׉�}�
���*V��v�ewFa��AI�#ޡ�i��/ �I�pT'�=��7b�f݊T�)fȳ4���mjt2�v2���G^����(t��E[ζr�4s4�Èl�c�BW���C��bt�!�n��l���{�;C���n���"�ڻ8��;��w�}��Vc�On��<���T�{�5��fqjqk�5��:�r��C�I��L5A���*Ɇ��X��\����쉼�ךU�h�Mջtu7	�2�L��ӥ���Ђj��9{�͓L���Ҽyَ�n���ur�:NX]u��v���ol���43���E��8ʘ�ǀ���睸�]R<�];^�]����+�"gl�!�%U���
*ޢ�Y)O�j;����O:�S8ɽ�y�W^j�١��˥�m+[s�i�����R�����K��o��Ѥ���O=�ն�p=c�K����h�����q����VR�$mngaY{���]L�I �Z�UQ��]�:ݓ����ڼ�mn�m�@����v�9����[a�fUP����ޓ��%Z3�a���ڨNxkl���{y����[��/z����M�x�ڭ�x�3V�%<�L�cz�`�91�^����vj�[�j�=,􀷺��vi�f��[3������-Ц1�s���{א)'C�+��o��:����ӲWVb�m��7cxA25�.r����#=g�׸�,9��'U��.U7n��:̩uz^��2�x���u�N��:�����:�aTq�VBkt9���(`�yt�\qL�2#ǽ|M. ԬŪ�q5�=Zރ6)eYiD�;u�Ux�mrɒ"������o`5Q�F���/����X$q�n��ٳ�,���
պg7(ޱ1�j�	D>�$���bީA�8u�X�UC����%�+�O6�Ct⼈+)ں�pvYЖfr�[T:�c]����K�$�/�;�ʴr���g*�BH��r�$������0�[9Z���56lC�c�G_>�V��vEX1M����"o�n��</�TƵ�~%c����3�S��W�֕m�s�%�����Wݽ�i�P:���L@/�82��5��,�m��n�h�KET�͝������FV_#�s�ܧ|����]ϱҽ��z��Rv3�,ͼ��[P���f�Uu#��@v�Zι�K�4 �w�[�҅�CK�<Uǻ7�v+��z�UD{Hx������Ul�-(6r��,u2�Q^m5�U�����^�t`�|;/���S�@�69�J�t��щu8M�F�N�k]�U�T�v�iR�.]]�]���Ust�]��(�j+�����D�8�o���Z�#�s���/j�&8��u{��������"9��Uݕ��=U�w%^o]*�˶�3:�*W��ͨ1gj�zMb���L���Wn�y�}�0>�pW�q�YZ�뙚�J\��BB�	�B�'��J��u�w�Hc���2�L�lL��-�2����l�2�k7�w��F�cÖ�P9,�9�Z���e�0�7����B�i�}uGO.�=�e
�L�VʦE<��׺�����e�r���hv�Q��6r�ۣ�������lɘh�[ݝ̩�4كf��y]�ժS1�A&*�:]����˱�D�;\���buw.�c���*����M�Xy���X�wUU����ͪ��ۿGQ33-��E���G`SvEkA
���N�3n�	�=���É�[t���c�jS��[�|�� {�f;��iDݺl�)�;s��aN�<Bx���<���g�h��y�d�F�_1к��W����<\wu����%eK�R&e��,�yW>�*�������sz�E�-�w�)T��j�p���WfnR.�׋Z3uw9�𛭻��)��c˾�t�ʢ)!�ydߟ��^���haL�Iv�tfE++kj�'BҪ�]ڪ�v�V,�5Y��9�nD��i�	N�t�[�P�d����6l_S\X��9R��eZ��zfT(f�6r���{�-�3Q:]��W-�1$6�}�iZǴ��5WVV9%;por�hURG��JLZ�՝C*��ʾ��5�QW	}��} ����z|�^��O^�dD����@a���ي\���ۍ�l�7�Ij��{]�&��
�w�[Tq�S���-Ӥ7L���b�[�/��㮠f$V���]�}�n�m�[�Z��������Oke�]²�Z*�G͋Ջ�9���r�MzU
L1Vw;�JZiފ�GF����^ �_m��{G����[|w�Yw��w*�q��}�*�t�5�hF�T�9�UX�U��D���6n�pc�����ǉ��뒹��9��'Ց�y��{���;���Ӕ�[w�e_�̇w�`�/Z/r�{ ��]\z�*5;v���ֻmus�R�;RG�n�p�;;{�̙���R�7��*���Cp�e:���4H�tL�w**i�$���ʇ����EU��2FJ��	��)%��&��#�Op��09����w���9�8�М��^h�=gFغ�x�����[�7z+g��.�庲[�s)�.�.5�z�0ӄ��9�����k'iїD�+诫3��JY4��)���T!vSV�a�[�J��9�q���T�U�@�9}�]��bՈ%η���yXk(���+�F�{�,���u]�WK���"��nwki��r�^��Aͳ�]Q�����2�y��h{��m*�O���]fu�3���w��E5���N\OV�a��곭�n����k(�˺�9�Y$�9�W���vd{���ǻ��Wrʮ�VB�3�4x�\Mͨw�R�r6�*ͅ��Bwoi�K��:�׷y�9�U<ӻ��;�h�e֝w��ܾg'ʱj-v^��0��Զ`V�,ǣ{����;�G{�7�V��%�W���:�W;�P|*�_,I�)"�D2�3zPW�P�i�5��/s@�bǕx/.ݬ�#,��z�5���ZQ	\J��*v��S�i��e�c]�gm�W�7�K�j��hQ�x.�W[ŉ-ۛ{�`&�E|��;�6������*n�3����)5NZӾ㽘gm�q�y�1�n5z/z��oT�+�}��ܚ��ڂP�>ɶ��V�gY4�q
5��ݙ�����jZâ�5m�m�lwjgr���`�g��d���aq�r�(˪�u�Wf�<���Qf+�������� ���x㽬�P����]��Pװ��Y�Y=����JJ:�vsXW��</s�t�y{Ys�ٝ��t�2�N��n�j��̩�u���9�b>�}��������eU�m�e�y��Vig���YѠMWY
�٧aX,��%v9պ���u,���K���:�U�.���y�D�Ӿ���5_fD�lA�kx�)d�j��W�MV�{�����B�=ܯ���U2�o��Eι	�uE+�nn��-��M*w���u���<C�Q�xh�K�|�V6(���+�Gn�@ӡ�R��v����Wo�:k]`�[�.0��Qᣗ ��]d����g�ʫ{Z��b��읠�ns�˃���t{-B�լ�Yy�TaXs�Q�ۯ�K�N�%q������r3�&�}Q�3;�7�U�C(к���I��R��t��%�Ճt��N�۾�R�t����X��JfG�MޱӬS*�����9�,�Y�;�����F7�JJ�9a�*L�H���B��β��O�[Q!'8�56����pUeof�e��=�n�;�cۤ��ף��!N�(�̡vt�fV{������V龈q
�ow1p��uYR�+]U�6<r���Zr�~ͲlmgP�v�sp�1��V����/x;�С��5xY��fN�5s��}:Y?*�x�M�uq��n�l\�d)��=�/�su�����2�֘Eҗ�U��sw���N��8+X�Ι"���S5�K];����]PǪ��n�v)h8�uj�i]����U��O���3�҇�[U܏�]��
Y��Y��]�T+�:��#f]����<�ͫ�̱�WtŻ�;�W-f��R�2�\-w���C��)(�fJ���3�M�`��e���L��{�n���wh�S��|֮�PgN�����:������̕���_[��R�B�;�w�y�Bľ��{5u�)]�������d�/#39���v�����w�u�2�݇�[\�Q8���$��К���UL̃j�Jy�7�{�4���K�u�(���%_�I���q�͚^��َ�М��fc6\�Ⱥ����/yG��)K��w�!+-��6gܟ
���T_q�p��k5ŗ��L��=�ӫ�Z�J��c��mq�pѝR�-l4������ΐ���!���ˣ��GP�{�XZ�$��((b�Ԗai�IN��;�曷6�[A�;pQ�UFʧw����sr�$44=�+[�ҙ�*CP�b\aݻZ-�p�i޻��Z���6�Npz�.���J�DUe�YM�tV�����ɽS>������TYT�Ewb�5��I��vb�;�d���m�
�[���;��wp[���A�r�QVh]u���:~m�\����\2��n�n�����lFT2�ά]ݬ՞��eؘ�`R��(�����tE�����	P���E�NU�vņ�����4x^�J��P��uA^ov��/4=��U�*��x#χ,�sJ�R����[mf>x{-;���T���P+�;t�s;Z��d�W�v�[�W�6��:�MŹ���]�>�0P��6��5ru�p`��z�B/�M$�4h����T���D�޹U�w
Qs�w+���v�wk����I%E�v̱9�̷N�R
���f��¹�]�E�ܺ�Q\˜���]x�3�u;7��Y�`$�{f�/f���r�Ӿ̲	�j�����a0���Y�|�L ��{Ξ�'�y�f4gnP���ϺfueR��se��_-�nK��(��Dݷ)�Xo���2�����t��W�m�W�y�sI�7k;�;{5��R�l�j��˙r͞S��/q�HXGp\�u���n�gmm�U���M˾60gGg3�-˲E-���恬!��zVL�3C{��f��)핷w��]X+��YctЊ!M�IT�V���}�B�,e��8�;W�ȯ��(n?���T�]c;�i���A]g�P�R�����*��D.��<3]JXEV剭i�x)uF��/4�s;37L�l�A{Seń*���.�VQn��*K4�\��cl���݄�j/�ꐺ]r��gd���F(�n�
�;�#��w1�����b��a�.�C��4E�j��%���6� ��E�lq.�G�k�ʕ��ɍvKd�Yu�m�7ۺr����uA��=�y�FJU�S.��ܴ���:�[���[˦����=[2s��I��e�y/1n��h��wS`��U��z���)/c��-u;�ܰ*�r�=2U\'��U�M�Cr&\���|�uU+7(���ͻ�5mծ��M�{�S�ʆ z!ͺ/v}�ZB�l���U�B����Gjv��]_Z����a�5��8�@t�X#+��J��g/E�)���9"�^��sw8w�\�b�U���g����2�gy���[�3z�s�?؄ BI� ��}���Q�U7#jVR�`�SԎ���cb]�ѕ(0��(�L�p�T��tlt%.���Q7 l�LӮ*ҕ�Tqpt�K\�2�,e�f��W��MGY��ά,*�4T�,b�(m uu
���b��Vi@�<&<�!�.-��k��/m�ݯ9����@�aV�ۓ%�q��;37Q��պf
LT�)q5m��T�R-��V0�W���&�6�JQ�-H�3\��B�v���1�G%tM�������K�ֺ�qya)CF���cef�"�1/Pn��U&crb�J��*��f[G3�j�c\����Z��,�ap�gF��aq�:m�e�1���`��h��b!WA�A�#����\2��� 9.hX7X��V̕e{6͕if֔��Ե���R7�+���+%�y�#��&����E�D;iIH�ZX��[&78�`oe��y<o���"��;Z�,vk�5���`,Օ�rճiv��$l4s�Vk���vA��LҪfk&�5�0����d��SLM�K�i���n	�)4ДPB�iԙ�%�h��b)�"K��Q����빢D��t]�snn�z�c�`�|�b����b4�y�K]�qG7f�(3aoai�-��W@�t�!�K������J�Y��Y���5��q�f22Z.R��\jW LJ❺�8nZ���l��^���G M�̩�`�%mήL�!��Lb�2�4�#1�.��A�2�L��4KY��̊an�X�WAŹ�\%�Km�6�]2%�qE�	�Ѩ�0��A�cBG
6%�u2g�`!�.h�V���bc��ufԐ�&�v�8ى��+6uŌʻXX�&V��iE�)e�Ŕ!�R&����bK2�`�	kkJ��f�pd�!e#��)���E���Зl�F�)M�4Ҕ���V�Fn�R�e[b8�H]��Khm�V`�	cʌ�^��pĐ��-K]�hA�6�܄�CpזުV�Ff��q�k��,(�X˩6�Ê]AY�����h�9qM�aز�Q�n�601�-�(�����n0��̴��	��V����G6�$ZY����e�9ĻJ���6���«�G�P��O�&�4YN�h�<�cs�!S�6���q[hv��+�e�B��k�qkC�.Ҍۗ$iTY��x/y7���^i��
�F ��Q���`E�jh@Maî�KZ��d�F��J�����0�"6���-��,͊��D4	b�/5�-�����Ѵ[]6V���H�%��K�de ��ڷi���n֭.j���h�b=�-V暸���0�\�5�t���]����V�Ĭe��M]H&�X,�F�x
ZCdˮ��ֹ�$�]�PB,�ZU�ji�׫q#6l�tĩ+c.�4Z6F[s�%{�C.X�&�`am�!�0W�+5�g�jl�eJ�$ -��n*˫\�P�G�غ�o6�\����0�鄦kc�hڰo\ٙ��0�"��]](���j�*�$�+��6�����G`dD�5�Q������`�,t��b��͢�
�,�G:R&���Q�;ru4�r�M����v(Jg�ͪx��kUn�Z���׷k�4̰�Z������F��R�m�)v����;�X�IX�ؖԙ�_�MQ�%�#uu�E3��u�:��b؎%����Z`p#��4-�r��EöM�ԩ(�J��ZVu�!5b̈�D��R9E�!���J�l�I�s
�0�Vوh�����"Ƙ����:�&���R�h�m�9�rcmP��m�Ij�n1Fț8�#,ئalT�ps�
X��\�f1�y�f�kUL�J9noc<�a��ke٢Ch���7b��g�e�Yc(���.�ج��1�0�6�0����)��.#�dX����D�%5���-2��� [��d����ʣ��o�M�K��VZY�Z�[���7eV(٩Sv��Hn�5����ғ=�P�ꕭ��Z$����Cch�.�����mт����Q�,m�WJ�J*�nv�Ғ�YJmL����	�BlE�t���5Z��Xu�k�0+��8�l-\L��(L2�B���CmBS�m�� s�0���h���<CT������c�B���U�"�ȡl����[�3.tr�q��*ŶL1a��Ɔn�f!�#��T�3W)y��([u�SF�H�fV�i���6�"�jM�:l�Pe�]-��̼�WE�i�ڐ�r�&���95���#6[c��l�m�k�^ΗC6�f^ٚ󗅲�Ab�]
���c�i\���Z�c+���.����ۘ�����촋�F(��F<�&����u�1-�S�B�*.�6Q�Mn0�sK*ee��EΖQ]*Q��ö���`�jL��лY,Ts�-Q�cD��gB�M��s��Jb�(8�bKM��ًWL�s� [M3zͅ�ҕ30�;.5vY�GS,���G��jfW���X�Զ���t�*8Ra�:��H��b�f=���4�u6kP ��K���W��Y��l&.� ����i�:"�-�A�k4��cU�L��b�=����pMp�=��ޮ� Y��T5gy��l��9�.�W�m�$lM�KY��%R�m,2�	Ky
�XJ�Gaf(�Z�1 (:����AB+���r�!lռa�c��ln��E���0��P֐�g2���Ee�.\�A�c6�6��X���]���"ZC9�ь�l�]��ČѱX�3f�H�m�/n�61���d13{	��-���t�f��\MZ��Pm��9#���f�\��-<���/��iV����kWZ��z�R.v�34F��1صڍ���,N�Y��>xkAb�ƙ̹� :6[��	�İ����v&l�f]�ͨ�^�r��\vs��j�0i5�ݖ4m��l�� %�n5���68�,�Lյe�ű+�R�\��al6��`fz����v�@#��Ǝz�b�nn�"3��@�#<˦�D&�[Շ$4�R՗F�� ͂�S-2��d��C$en��`2�q��l�M�Ԏ����W\��8b=FKM[-+�n��X�yv��"�Gk�ц��|��z�crԽ(�x�
V�Gi5�e�GYa�"�*[:�l�^1snLA���L���;F����Z�Kv5r����p�-�H�lm��)0�����%��HTh��Hhca�1B����i�]02-GM`:�r���RR�f�ధ��T4�e����ŷih/ ��V�u�L$������;P#���h#ZW��Q�uqd�f�u[D#X�R���Gu��.�Ս�����,�
�`�.�aFQ�7-�epu���p�����&(p%ً3��e�W��j�g���x�ڔ.,�S;J�1*�f��i-����]E��S[K�<�P�78lt�tf`.�׮�B0jCX�a.(���Ѷ�cn
���`D�8��)i���)���0��Tҗs������n�
䣊�j
�ٙ(cb��k���h�maz�m<�����vf@�[H�H�.�J�tVh�e�1�� z-�K��e:,E���kms�ď)��f��h0%�n؊�`��)�e���-`̶k�lضe�B1��2�Į(�\���JKWi��*�-����[l��[W S,5,�����F���a�j���BК���2�s6#.&3J�m�KS3�:ͭvu�T�/-&�J(c$5�H�]tAԔ��qZ�.1L��^�ڴs�e�8��rg��x��P�Y�Cs��#fUB�š�W\u�4����`ؼv�K`�:���pܻ�cO16�BP�Z�s�m�Ԉ"jj+�m+�i��b���i5��u������a0M����Rb6hк�[cX��f;c3[�� m��9��tr��/ZV�Z���!�S�pl��M/^�b��/m +Cg�5��͡���I.&�dH�K�i�B����#���t.(#5�ٲh�Z�\k�A]4t`�e�c$���SA��y�󴢨3B\WkiV�	TԖ�l���j[�����l��43u�,��
�J�$!�E�9�%��)���̴uFQ3.W��M�!lE��(Sˉ6�2R^���T�]Qfk��c+x�a��:f���q������Q!��HۥP��f��c`��ǹ�7W	��H5e��2�-c0dԱas+�l����%#(bh]r�������eс"��M-�k��A;]F�6.rL.��e�M�tmp]El���0Ket#�]+��ݱ�L�T�����8�Ye�a��1�@s3�v��A�Zc���S]�݂X��#��٢ƼFX��)�,�Bb�d��3�D���)[��4�*�3&����X����Ņ���[t���ͤ&�-�"k]qب��3����lIiv�JF�"kes�4BdՈ�	�]1n�V[��7��AZڣ��j��kf�XЙ[x��oR��K�SL�� ��]c1&�c-�h%]r���M����cD�]3JԪ	�J!�����ְ�޴)�Ggv)3�J;*nb;�VmhfbF�m؍qY��ц���J��;f5#W&.]K3��ŗ�WX\ո+�Tm��㴤[�Q!��b�E�V#L�Y�i��M���s�T,Ԙ*��1��+.�u@*��v�����Yc��L��ZS%3���)e°���-͙E�hޱ���5�JЅXV�i�-�mE.DaU-��Jl�ٙk��벥m]�]5����[����A��T��f�e�MkJ���]�[a���4u���t�	.�5iq(��nv�53�e����k����DG.n&Yq1���]n�,�]	b���pm���,[��4���J��a��]+��W�l�w2�����Ա�մٍ2uf��uV
�X�3�+W3eX��F<df���1�Ƭ�a� ��;�H pt���%��tGj�d�8��s��#��m�vv'D�B��6ˎ����G�Q'f���Rt�r�e	�pm���8�!�$H�ݢ�B�	r!�9��B(R8$�N�hw#�D�$@�RmbREVd�I!�JuĳDq	HqШ�^ڃ��'!"y�s�8J�("��Q�i
��s�ã��㈢��b!q�����s�8\��I��)N$�(���:S��9 �B��Qr�3�'
(�������$�$
�۳��R[[�qΐ�{�����,H�8H$���myX8:^ZD�(9q ��$�/�݇�4j�K��5iy�֡ �m��%�X ����`�%+�K�X�<m,�����)�a�W�.�i���0a�,�V�b<�7k�[F�հ��m�5Α�,�m��^K�6�$�knA��l�� �l�ns�W]`,#ef\,M��R�L�R�9p��V4�)ri�6��f��Lk�
&�l�3,�ۇ�&f�4&��A.��Dte�w�J%�Y�e��HK�ʪD^Z��4V��Vg�/�4o.���3K�Ѵ�ֲ��]2�h��r
Rj Lj*G3m�4a9��B�k6���0���^Mv҅!�W��[���F
S�[,S-��D�,�J+z�6���n�gE�f��	P�cL�ͬ�ؓml��j���iau�Dc��+mb��+�i,���]����P68	#v�X���Rf���`�b�iI��� څک��-0@�cf4s��6�-w둨����r۝��ΰ�ĵ�D���!��QA$4��e�3b�GJmd��bQ5宆��
�U4�,��G.��d�g���Km�XRh�+t
Ȧ�4*ue��Hź-�)I�JXiqW�F�,h*)ric!J�R��Ùf�1t7V�#K	�D���qe5rݜl�B�^���ei��9j�f �,ҁ�q��@��Q�A�X�Еe)k�Xڌ:��lˈ�J.����Dr�3c6�0Ip��.�1XbZ���T�F��U�2���&���ݙS,�2�������Y��n
hf��͠��`��h��M��.c����Z�K���7��Z[��&��ji���f���Kfe뚸(Zͱ[v�95��`ZuSD���7ͦʜ1օݸͷ��ҙ�ҮIte�`a�*
�jӕn�k�H[(7@q73L[a��.V$Fb�ZRSrK��YWA���-p�Uƶ�{GP{C����f����Дl�\e3��SMk:I&+���E(P�x,)[l����Njʌz���[t��Z+0�,��%!Ҷ�H,��F�b��NX��R�H�VXK� ��Ճ���B��o	d���YaJ��R�c60*�,�P��"*��P�e�Kq��"G��l޴���m������'�����h:(�ĺ����J�m�U!��S3L��2�R6Q�.��m}���a}A� AmU/�ɏ�5{��_ �*�/	��5Bͯ����%�J@$�B*���͖���A"JR^{�ul�l	������t���q�U�c�ޠ]�"@�g�}%���$������S9���}�8u�u����G,Y�� �%}$��l+�o�o�T��O+��$A^W�1��Ŏ�	�9C�qX#��}ۜ�3�m	��4�}�,%/�$IH���ŀd��Y���`=�wپ����'$���������\���+"JS=�|����y	����n(��\�&q�Gd�e�^\q�q�YFBdjB�]�;�O�/�}��ߟX��/��X��3���L��ks�X�^"����O n���I�X.RDȒ31 �9��������rE�Sq^p6���n5���$�b��/e>=�mqΨ��hM�_�y�^�&�O\P,~��)���	�sU����t���qc��w�P�6���L/a}�+��ګ얇�DGJ@~Kd���IW��^�M�ilTμ�oud�E�w?}`�[���A"�J� ��)�J����_����/f矽�y������&W� %/��a��n���Z�3�,��@�D���L�( d��Zv��}�UӠf�����v˞����w�y�������%�`V}$��t�FQ��Ut�e3vX.M.ؗ=��طR�ÄY�f��Af��3%T�ӽ�������d�A"JB\��S}#QMʜ�t��
�����V�P�	yA���P���	� *��Un�����z3��zD���]y�f�Sb���h �D����)�@�q�u�E�\��?IA"�D�3����OP�ӏ`Z{3o��;"�u8�f�y�pGN!	N�����5����kK.�����Θ�LJ쒂Aַp��.���s�W'vvɝ%cO��n/�r�I_`�X����>�G[yt[VA��سґ%)s;�q���4������v����P���$A|~�����dA��l&G��^��)v/�rs�y�op����<���+�#�,�H~"JFU��߰�
ڿ�6ҺR0H�&�`�6�vu��.R�q�ڋ��"�EY��,�����H��A�	�6V�n�3׸}�l[��dP���u�^k�"m��|��,+�D��>���n�B�cAݏ�l{�I�m����S�ru�C�렁�A"�qZ*YZ��cA���\V?H����$CIE���P�R��+}I�����F�"J@��fJ@�%}$@�kfܡJ�@~�_9�$AW+�I۲[�)���y(�y[���{i�.�1��c���]��["�P����:n�+�}V�i��2���}����n��4�J�a۱�ҙI�V_nŻZ��/�r��d���I_)%�J&Ay�N�E}���]{��t��9L6��wz��t.P@��D�mר�]w��{������?[����h�q2��ZTR�iW0�ٖ�]�2:UZ[U�!Z�<X��oH��e�w����˯v޺�Rlf[�.�H�_�mg}�V=��ʯw���{ԁ�)$����@����t�����nQ�r�{���-�;��>��	��9~���z�.�yz��^�=��I,Y�$3#��P��7m�^�y��p=:�".PFH��"�"C�{w:���o��/;� ϒ��$�q�o��}���N���:���|~��>	�<�}\A����I����A	��2E��m�[
���]����l[��g��?w ��%��Ic9J1�^�7��vbu����B��_qF�;ˊ�k<����=�����x��Kۊ������/`Ѝ����[LJ�Gh�2˭�%t��8r�4��۵����u�v*6�3n�S�MYkof#3c#K����bm��D,.�Q��#��Ŋ���.p˥��^.���Q4)r���b���ʯ�s�6��:�3�R�� Q�э�3RVf+��!�[��w�)�`@����@���`��)0�A��Pe�j�!��R�f0���^��s/����C�CSDX��%ı��Dt�v�em��s@�.����m�g����}]�=��IZ$IHE�����Oqu��:r��\<OEc1fаAm}Ӗ�D��D�H��
�C.�Pz�eh�މ|~��!�[[z�V���4��߈q$�A�AЍլ2)D�=�Au�G�+�"��q���6�^л��{۱l�.���y�����?I_/�����k�	զ��B����fJDD���wI��Oqu��:w�������^s+<-�JT,����"d��2 ��j3qVz]�y}�r���>����:��k�6��,)|AfF�ǋq�g�Q@��0a Q�D$!H�aTwXn%����j7krYr��KfXP�~|�������%�_��ݛs��_�`~�1��s�.GA�侒!fJ@�R���<+���bŲ����Ri�V����S�;��-c�ǟl��/�t�v"`���@�p����xN�n��V�����wTzoV�5���t� �Gu!S��Nf��s�q>�ӽ`�vP@�\�����OWK"���ǧ+I_	0/��UaN��.��}�춹�	/��{^ �6�9b����$�D�ń3=�?<��BM��%<����ٷ<J�w�s�}n/�0n����}/�|~�A|C������R%�%y�4��Ee *����fo�9GS�9��E���fH&)��bs�:��)@��D@Q%n�T&V2ʋyq��� �jA�9ܸ�}w��������?H�_I�:7�����3��uD/2�NX�A�� �yO�IH�%�&J�2�+7�C������t�ݛ���]��y������%K�xVd�٩	��K�"u A�IIZ�+,Z�y�������xhǽ��Q罵�uc��ẕ��lIR��B;×�[�c���bk��������<�[r�q�:�U
.c�7v�穇y��ޠA��$�}$_h���D��6��i��>��֬�9����Ib�F��|�o����{^D�@���iý�/,x�6��C�/��X�A�� �( d���]����_jW�wn���j.�{�<&�Vr�I�/��X7ǽ�1�k)�ͫ�p��	�h�̹�Vi�����2��q�T#��p.���oF�6-�����N������w����vN����НO�ww����0��W�'{Xϴt/�	�A�A�� �H��=���ѩ�`�~�K㭡�=^�Y�V��VH��2�A\���=��=H�Q��q�@�O]��A��A$_X����eW-����7f��E��}'�2+9� �IIZG�V�Qw��q���Ր~��zR	)|��t��f�oB[�"wz�eCӚ�q��
V�#���rxWb��a���}n�-�V�t�(��l�t�=�D�ewe�Ri�'s�+x���ٻxݙw�6��n��U����@�d�� H�?H�����Z�B}�D ��|�����;v �x	i@rX�%  �)�)�{����"b˦��F;M���V�$*���i�nرsuK�Nj�5Izk��s�C��Dy�\���2!��۳7=��о��JB��a�+�����?>K�$�,)H��"�{<��-rB��{�g�HH~�O�:N��}��Ty�N�}`����A"��r��Q���#�j�[�Ȓ�b�H�����]�����PGnw)�9��&� ��,�H�%}$��}��IC� 적��|D�%~}ݻ7sÄ]��@��Y��\�����}_xǤ�`�H�D��I/�+yе��>����T��g���9��Ȩ�����A�����!~�����YK6��T��M�첮��{��[��'7��;bՒQ�vL��T��#G�Cgx9>�~���ϥ�nw���u��=oX��2��Xv��C^�wXX]���@�����*����)����f���bM5Gi3&�3T�m�x�V*g(9��ۡ-�[n���SM����-��*�V��-��3�!�-md%��ƹk9��r�YqR�i����62�#�j�."bafz��Z%m�y�]k��U��Gi���`Cv0�\��e�a�jÊB`�8������})JyhM��L\�\�*��!X0���R����%{������O�l��K�����ǽ栍��\眃u�+��-կư^�#��,�W��$���`�d����k�g�wkgU	���d�/�+���ٹ���}'��E���I&s�GO���Y���)d�����r���S�;�wbm�����*<���M�h�������"w�[;ۖ2�L�J_�K��y�_I�vGދ�����9� �x��Hy=Pp��y��멪Ǿ.R��C��H��d�� �(#]�Τ��dH(MCj���ݛ��x.��(x|��/����!�
�����|���]���tE�JBSX!�u�.u�F�ͩ\�&�aIf�0�]���_p�Wpy}%i�)E���;���Ty�t�}a��/:�Ϲ>��u���iW�J�/�E�v����n;��x�yR�R�(S	G��s�um�#*X�)�ؠ�b]��VU�V����ˣ��&��5�_e<�XT�ۘ�
ʤ�RՓ?ւme��c]�n��M��Ac�G,Y���Öe�pz�n�o�����2E`������`U��_h�x���c���%po�����_ ��J�	%�2R���F���s��gW�$�"�d�fy�q;��e��?uLx̾��]N���j�?w ��D�H��� ~�����|��~�d���5���ȧN�i�5� �,X2R �D��g(�b�N���|��D��m]]
R�6�2V[V� ��[�nVz�]Xa�a����~|��=��i�l���+C��I;f;���k�x!W�^�]S9詬����D�2K�J��IH����yS�zj��% A��z�]�:oL��>ss���	�A~.W�D%,��3/=�u~�_ @=9YE�xfb�S&o�݈�b^�*�0�	ˏ*��e��!0@��P*�vdP��&�o*�;22�V��TY�&qκ��˭�9�(��:�+��_�:)�]�v-z��l�oJE�[�4��E�B�����+Wm� �׫��鹓��ʑmVEu�o	��-�	ᨏK�l�[2�K�%-�Ŕ�i��V�Tfu�,�a�*K���zW2.���3vi��-��@�4묨�گ6�:�3����r.�ƥn��k&MÏ�h9ݝwۘ�yi�hA]����z��=����iZu�J�T��W@�ā�xVu��n:��ee����rbm:A�wKܝ[�\�6#>��ǲ��m:)1��`��N�Aوt
�wW�)[�P�9wL��A~W6�޻r�N���hhv�V�
�۩v�-{����y7z�&���+/��r�:*n˕˓��:�*f�c6��w*�]���m�`W�*�i%)���b���E�ٳY��:�:�U���ľ�*�ȏ�
*q�&�Aǀ�Z�lNV����o���sk��S���Pn��p�n��.��l�.귴[���U5C�fW"K���uv�dDUa��[�ب�;{s��w�uNH�t�S�7�.t���p�*.ɵv�:um�c���̘]Wˀ�N����w�����8�BҬ�^�h�T�ɖ����482���$g^Աah��ݑ������k��� �S5,Z7���ͧz0֪�7a�E����M�c1XQ��Z�鬒���U���EF��uk��N!/�#f�]q�5�N�����ﲵ�TQ����]S����m�^��^i�i�`�r:q��^۠�	8f���=�%�G��tiYM{ד�[vY��*s���H��:	#�D8��΄��y�����8�9=lE�$�E�RG�'f�f�N'r�\rQf���G9�$�ÇN-�n []�"{Y*w8�Ȣ�!"H�k!�♄�����ؗ9
9	I.���9�tH�H�:�Jw�X��n�Nmd��8�;l5�bJֳ��͋��kZ�15T,Q�uC
�*��k}���k3�y����_���Qi� RAe��e��5RAaY��6�R
e���$Je.e��%$�a�;H)���:{w�z�f��ZA�D) �Y�@���)�}�3c%$*fQ���_�����������ax}���A^e��H)(B�o��i�q��P7��G�eV�[׾����x��Xi ��p5� ��높� fQi �̸��) ���������-'��S��N���)o��4w[�}���ߺV����I�g�?�
B�P�- ��Z+���SB0�ˆ��2RA@̢�]��o���{������~2�n+cy��YXݝ��@�s��Z6:�ۥ-v�$rG��O�tךO�H)(�~��L�e$
;��$�H+�p5� �*�p�>�V��s��-�~�]��3`I@���}�������>2N.}p-�RAa_�{P�AH(�- �N�̸��) ��ˆ�
CeP�ZA�D) �k���_�U{���7������L;���L��I
C��4�~2����_��1,U��H�m�~4�RP�0�}p�&�) �w�ZA`i����e6{G��_7��)�g.H/F gh�ЁI��K����4$��¦fjH,63(��) �P�\ˁh]���Z?-^[D��zSs�(��0����i!U@s�ZAH)�w5�
Aa��3���P3(���L) �e��i �������Q��-��w놙62�
N~�I�������kTAH4T32ᴂ��כ�uv�/՞�$�H�>��%/�p-	) �HO�s��Y_~3)���B�l��5��R>\����5�����r�M�N]sW7�����ت�.�wQ�O\�\
?iы6�^<��ԕ�|�{���$;~�� �fQi �S���hJH,32�n�
B���- ��\ʁi4�L32�$'?w��Օ>�a���.v����������}9� }� ���C<˄-	�� ��{`hs��u�O���L��Q��*\ks��b�+*8����96�Z�pi�en����ި��@��ʌ��TCI) ��������q� fQi4�$J~��|�I���m(�vb�>G���{ w��|	^�VQ��i�: �R����j�ЁL=��$����4�R
As(>#$��3.H)�߳�>�ٯ=���X|�X4�^�@Ѫ ���z���>�Y���Q��Ӫ�w�}E��
H)�*��%$��Ci����E��oU����޾��i��N�P-BRAa��p�AHl*��QiE���e��AM S̸i�d���D3(�~y��}�MC�^S�����,K���Ay��
Aa�e�L��I���M$2�ZAH:�̸m �`Re�@���뇿w�v�����oz��y��hi%$��P�Aa�?e�HRAH.e@I $��Fҏw`�*��|	�7��D���*�稴��D) �����{���� i ��
a�߮f�%$*!��i ���TH)>B�fe�L�I�2�$���P5������f]���R���I:Ǜ��O2�oΫ=� H6��) ��%?e@���XjgsP�AH(�ZN�Y(e9���t��{ދ�9WY�I�]D�8&����ͅ����N��(i{��u5�5�+���w�^]�uN��.��5Z��i��]
�ng�J��}��Z�����րU�"��ڊ� e��VB��C&�5U�b����/+�ƺ�+��y3/�V<Q����y�+h�,f���-���[�h���a��u	�!ųf]�0A(����5�dI(�iM0��1LHlB������gk�4ئ�����i���xl&�e�qv�xe]�9�e�T��o,��XX.ҧR)1�\dn�X��+�>������Yw-���b˖��cL�-	�V�Y�f�Mb��Mh��|�Xk�����
A@��ZA�D) �W}��SQ�fe�L��I
�fQ���_�_��{���}��nq��y �r��a�������ﵱ�������r�ú��L�I�ݳI������p- �T32ᴂ�`Re���R
�\CI) ��<��z��������Aa�� g�-&����L���h�����Q���^z ��?�~��$?U�QiAD) �}p- ���fe�L����g5��}&$-�F�
AH+�p- ��\4Ƀ) �fQi �̸��H���n~#�Nq��{5�z�y�8��c����﻿���O�$��e��4$���jH,63(��B�%�̸�����3,6�
C��U�{�[�w�߀��- �(�$��j��0��ld����E������{����s-�<�$�X~a������\4ɸ�H(�=��_yg9����A_ݸ�R�C��ᴂ�H�Zj RAeFJ\ˁi ����Ci��
@̢�g5�4Uk��~(��ंɃ)s��5�~�;�u�����}��RAa��ô����z�H:
!I�]��ZAM S̸i�d���fQ����?~\�g�#��YX7���bJ%Lâ��7C+7!��R7�4V��.p��f�6�t���\H)?S�ˆ�62�
O޳I���A\ˁ�TAH,32���>�s_D���7u���| ���) �>�k�{�{%/9p-RAa]�jH,63�ZM!I �e��%$�a��AHUP�ZA�D) ��r�~��������Cg9p�̬Q��^#�$�����z���%zz��v�,%�����l�33���� ���>��of�ڻ�t��)�z�����;�5Ӽ�{�@�����R��p�AH(tC=F�/_ϳ��;����̷8��H+ܸ�R~�S�d��H(��I���
�\צ����^�u�}| �{��l
@�h�ЁI�)}��
Aa���Ci��Re�HRAd�R�\@�s�'i��������}���_o?�Xfz��� �(*���- ��Z+��H)��fe�L�%$�- ��
H+�a���
F���_w�a���2}I�h�����A_~��R��f\6�]��}���~��3���߷߿@P;�-?D
H,�J_�p- ���}e]��{=��AH(����Y)����4%$�a�i �fQi �R�5�
Aa��1��v��}�O� x7�~t�Z�^W��m����H+ܰ�0�AIQ
a���I �g����R
�\Q �P�ˆ���{�Y�]mMSp����,	f�{G\j�6f,)V8��@���f���W@���O�YQ��|���RAaS������`3(��B�%�̸��k?{ٺ߿}_~�=�{��$���� �5������~�O�W�7tZA�!I��5�
Aa�ˆ��JH(TC2�$��W2��H)�f\4�R
u��:��}�������Ѥ��끭P�>#����>�����k�x�+>ߠ(��R?%.�p-$���;�$Re��s)���)u�h����H)
�@g�����RAjVf�ZAM S̸i �7̣H���uk�7}�(r�`���ڎ'[q]�B����%ec�e��J�f�ǸC}�_HW%�2���;�Z�Gm�b2���³��}���_{��o�Z}�q��<�W�a�i ��\4�R
��i �4�A\ˁ��R̸i ���E��) ���:{�z�"����:���높��z�I��$JK�$ �OwS�oT{���| ��?�A�v�R*���- �Q
H/�s��-�~��- ��
a�z�n2RAB��F�) �e��i ��p�AH(��i �4�A\ˁ��2�Yow} �T=��6G��r��c�W3n<�=�����#=H������D��Yvz=�Fٰ�� `�l��Y���sE1�ۡ�h[��sD׊��Y�̫
̓A_ܱ��=��/�H��c��m��3��)���C�9Et^, �#A�K�"�V Dlx�9}z/�H�Gu$��Y��fL�$�X �P@���!�yk<�u���9X@�"�|D���K�,�Ay���v.l��;ŋ��}�'Aw�X2R �D���l[�~޶��]S�u�4���[�H��^Ν����O3��<�s��K�Y���^�����J�7l���'���9d���C�M��f�ܒ��c�}Z��f�Ȯ�C�y�5b�~| v8��3��2R �%!�I,Y��ܻ�&$r^�W�"��duh�C(�<��z�����.P_"�$�G�Շ�v�
�e]���';-��J��Yu�n��H:`Q@.@�B�.�"��t4���A�G���$���V�ֵ�9瘱x[���FS��+��#9��V�	RI�%GUlk5R�{`W�ے�;�6#S�����5s9>r�����r�$6���K}�U�F�ޫ���j�{�����b)%_f�ҭc�3�2�מ�l3�����=������ �$=�)�K�|\���?{�/��X���9�>��ft����$gR ���p��,��� A!��K	�� �(/��Y�^���(R{By �Ԥ��{�7�#]�'�P���/��9~�/��K.w������c���Yl��F�v*�ћ*��t�ۊ:ZW�/��ź�33�R��y_}�\v:�|����j9���;�~?}��:��Bf�X���@"GJ�؅�J%�;f��I�9�fha#�*�u�L�kˡ]�a #vNlbV�MK��Y]�4���K0�Gٌ4v�i�F8b�a�%��	5��f$V�\��f�J�z�&&2���$�UQi0\ -��"��F�dn�f���V��0�L�@�V�bb�+nLSY�lE+�f��R��`B��4c�~�����+���(����U����u�
�1�����YM`Vx��J�� ��d����$���fxzf�2o'xX��J��P�	ܠ���A�~���Y	�ҏ�m����zg����}"��[)�Vn3�2g<-Ƃ	u��,X2T�Z#�ф<�G�X���L�H��"0Y��_��r���vl�<�6�r���VA��b��& �dH"���4��Rx-Ǿ �[H#����I���f{��T7���`��,Nx|�1��ߨ��޽#�Yl�n1���IA|~��.�����rŹ����������HzKd�AIY{Y�t1.�CV(�TMѢ֗m\1nK,f�#
۪���٘2�ܽ��/����~9�+�"�� ���o�ݏ��{M��y}W�%�v,�w��9@���Ⱦ���	Wι罬���U��[�_Cݵ]�v�HA+�M�,k�1S����U1w�V�֖76�����I�����o�ʱ�k�a�Щ���i<ˡダ|> ��۱�A�39y���V�0\�#gxX ������R���]��0K_������"D�D��%�0_q�G��&��\�.��'W�%x��/�+�%@D�����u�]��/�'r>w�Df@�6g5�z�m[��tU}y�	�9D9�z�����+�)�?V�d�@��D,�UOPGC#��[�非���`��CgxX'z� �(#$_\�.�}�yn�5M/�.�@�vU���[GMU��-N�c��n[��XK5y�2���t>���|$ϗ�D.��χ���ZS�E4N���Q+�;Ԉ#��,�R �% �]�%�/6n�~��Q�5Y{�_t��{���yy��U}oD�s�Qr$�!�u-���s�ŀzR �:�D,�H���+Ҫ3=�DSv�ڕf���Շ��f7�k�d��N�:y���ۓ�݋�����w�Np�Bg�o�,ʩ:�T��fݴ��;����7�{3�۞Y3�l��	ޠ����YPG�wp��ͯFʆ-����|7����N��0����w��8�!�}�������ҥ*/���=H$�I@ d���-��gWz�����ŗ#��������ϼ ��`�����f!2v�N�
�	(D�L�B�:�Xh�!(ݶM�nh��%4J���4(�Qt�}���"OX�% A"JIG=������;��5��mWs� {h {���?	_|~�|&H��~š�o�lυ�l�?��AE?Sze=x��N�|A"z�#�!fJ�Rַ��BR#�]�%A2PFH��F�3�w>qEM=��u�n�.�*�ǢA+�A�@�"_I�d�����8]�z/��#g!ԁ�)��{;�sא�=�-��N�@�v+N�V�_yG�Ǟ��/�"%o�k�3��mݎ���]��p�p�{{7�	[�P�4h���C�f^W��x�;��pR�{5��"��� j��辿�_	3���YH���b71�j����h(��[�)�ڧ�|����OR ��d�R��y��o��ύ���.q`!is��;-��\Mк�C3Q�	�LVjf�����������u}$[��\��?w�L�r7�o~�D��b���˔����_�������Ń%"	Rc�����evb�}H��H��{;��ْ���A���� ���/{��䖎��h ~� �;"��"D?H��D+�y+rƓ��}Zen���Ż�A���^u�2R �% D��U�&x����OP�ו����dA)~���;y��ϧ{�	�������鷙_��B�J@���"H�������v�m�,�=��{��PLΠ�xX �P(#$V2!_U%O�g���U��:�)�ێTr�f骄p�z��K����K�U�J��g�e���F+獥>��L�t�w^ͳor�-kt�WBp��.�Χ�a ��瓻8��97�e��Ք5ȳ��[,�	o�����ٳm��J
�)�V�a:�̚E�S����;�����]QR�^e.���F������l>�������b={]}3�>�2�ǭP�u�/�j���OWT[�v�h����pt�����e��NW#�mf]]��	 ��d���9��G�%'E��=��t�k�����1�v��eI�6�s�/p,��ԍ�OV�M�w�B
�/�Wv75W_9]U�]fK�#�f�R�]_��Å�v�L����G��ʷ�5�c-�+�p���8 ��]Z_P�5��{շz�t�3|L��8t:��{N�F�l����W85v�ϖ��V6��\(_)O9��ͼ��1Xj�kz�{��Eo��gi�߱rY\�k��|���j�c�)�Ļݔgj2��{�`�i���-����]�JE귫�����<�D��ͼ��+�7Ut��&dU�x7�y�{�u.�ud@v�ݺ<�XH�U�v��	����+m��E����3n�����[a4�p�VT�ՌY8,;�_A�A�A���Md������]hI��meg,�j��3�Z�Ƿ;��Ǧs���P���T�wob���ݘ���K�����SZf���2�J�C:��}���K�9K�����ܚ8Z��Ϧ;0CLSch1U��֞�
�Y��8��[e��
��h�U�$��99�"v6����mh��"� ��2�'),�iвΔ��� ��[��F�-$�+-f���RD���[�gZ�i)��!�~��G�3������z��8Np���8e�aͫs��[m�Ύ��̹�r'DEr�m�b��6f�|�!�N)�ք�m���3Nge�6�Nws6c;qe��I�iGm��������m}�'ygei�Y֜�Ґt����Aܝ��e`&c�M�7)�2ɵ���	e���6�2k[q�,�p_{y8��-�������iǶ̜�;Ns��z�Ro>y?K1sV5���ʴ��8�
�RV�����AB]m]e0�k���q+�FZns3��MD�	A\
�v����^`п���yY|����- ���f���S^YsZ�sih���ٝa�We��+e,��2Њf�/8$n��a�{^M�!Lڳ`�*��屘I.V�����"�3Vd����\�c`X#r�Kj]sYz�2�j1�Ⴔ����ؘ���B���a��B��1*�Wm�mP���KhRշ�֛ �.��j���Ńε�[ˍ���E�*1m���]Z�6Q��@HEu�v�����-R�ext�o*xV��3VU�����\T��+�*u���XT��X�&�ܕ���ݗhb��,��\jE#(�p)4�FX��Y3�98�Z�Aʑ�U�K672���Ci`pD��	����b�ٗ�hn���Y]�й�$��L���&�0,R.��f��u�X�&�-ȑ�L�qiV��-�Z �%nV�m)T���Fa�Jۡ��]�+�ԑxhu��^sf�)@c�7
Z[�LAL�&��9����F�s�V�`ԭ��"V&��G	�ZmXlLJ$͋���ilA�b��6�4�8���k6vȑ-0.5�IZ��ƐFK�����H�V�t46�0Z���VK�{lfX�mV��n!�km�����J��	��.n�qf4�Y�sF�e3��h2�mS�W5���*c2���,c�����fԹ�2�v��i �Ҭ\i��`�͛��J��tW2�نu���3�ÍK|�����0�i�@\���v�@�-a�J�&f�&ʗf�R�J���2ЖC(��EI^�1����usJ���YR��]�U+T���K8���v�@4ͯ6(�GP�ЌFh�ǖH&!��{aaLm��;m�u�,M�b&֩)xs15��p�c�\]�`��������f�iģ�X�L�*cf�-URն��ە3�73�]�9�eѪ	���b����&L�m�wI��y��n36�]��kP2g�����6p鴱b��T@�m"�;��+esJc59@v@��mM�V�-%���,�I�1� k��j��1���IX�*�Cm���)�j>
ðh�%+Ihl���R�� �i�bDդ6�\�4�M�,�wimm������	�˹!ٞM�tU�s�Y�jBؓXܮgY��t�
�
K��g��aiY�����쿺�"9^u�6��nfZ��eA4L�`�&C=\V��m�e�|�������%�����w�j	�A:�B�����`~��,�R��D��K	��!ڡg��ЩN����Od~����6n�7�N��s��3�@�'��;��U����6ř���_~�X�%|�"J�5h�;l��d�M�/ndPLΠ�z�z�?9A|d��E� A��t6�F�]���#y~̙�3$(��7��Q�1��8�[��ټW"�[�%"#�/��X�L��A$K5��;d�4�����So���F���_\�D��"�"�o��ׁ�����l���KH��6����j5q����蜱hǳق�u�pf�M=k�����G�!) A"J_-�������E�����hy;���7�u@ w�#�+ Ȃ �%�+�����*�1���,h�!.�����튙���`�d.�OsUˉ���uw��	��W)�&�{o#iv��C�`޽sJ0m�W�J.6mZ��:^k�}�� *�ó�_O܁�^o��d�g�1�8�A��ؐA�b�2U��1����� �Ծ#�!`�P@�d���~ �"��W�*}ʨ�w�N�wu��]'���%{�z$Vl���b��$�fJ_��rgyo��+��_t��Rn��gz<��A3:�}��z�#V`�nu}��A�r���2E��@�&Qw'g�U�����M�f4�t������4��H�h#���'+}���o�5���)`$5������#-[����ٷ4��nvB���l���߽��s��r�2E�Ȃ�̏=ާ��fo#y�� ����Y+m� �r��_/�����H������Z�1�ͤ$N�������w$�/:�}��PD�d��~�5o�V4��y� �+��$A�K�"�Q�ь��ۛRxU	;�[��vV(��Wۛy��-[�X����/~�C*S.�-�M��M�����6�7&g;Ň:	���"z� ���d�@����%���:<�k���J����"������{}6n�7�N��o���b�W{~�/����pHn�M����1�����N��:w����&y�#��A|A��_I�~���%ܟ.�.���-M�F:��@F�h˦l M�0�fa�ЊE����b$e��:hC�����p��d���b
��Y�-8;ŋo8��T�
�6�S ���X3�H���I.������<4I'�����F��� ���2?gy=��7yϧym�}s�_�cr����/|�?W�e�>�_'�d�,�H�%e;�(����ȯ:��xX?���$_X�~�|��j}w��ˤ9�ƾ�@��%�@T��ٖ����8�H͉#}����,��wm��0vVs�����*j����U�1f���6+z�u�Dvf���ڻjՍ*�o7~��ک�m߲�t5�y�T����}���ҿ�/��X�L��%��~��}�R��-��sfw�r�$o���w���A��?H���ĥ�V��!$�m��r)�JBY�m�H�Tb6ᖱ,�"ۺ�2��(�FĮ�yH������RKd�{�����Ey�9���޽���������Ȭ�(#� L�_�[��-�"��L�[;�,?��S?�AT����V��L1x�c�ؐAר s#�P�6�8��7�3)�.�3�"	��2EdI@�쭫�����h��>��{w.d��9�N�@�~VA�����%�J_u;�K�fu;�b���H���f�+u�^%��%N��}N�2�J�<�ު�>7ڬ��A�@ L�_�"�#���G�f�>B��_���Z�Bb�ǃo�3c�{"�̉ ��T���a��7H��_�����n��j~����^�:m���S��r��c�[U���*��=D�0ie�o3W�R"&V��&Ku��C߾�� ��w�R�ڮ�4؅���̫fu���
0��9bL�;'j�\���Kn�&�1F0���i(�+�!�F5�l��0�j�ơ0�`��hu�L�{[r���Usm�����
�-�)I �L�f��B:[kL�h�e��q�mWD��doVKm����r[�R��LLa���1Ŷ� ��V���š����󩝃&�F$
�7����Z)�v��B��W����"@��[	D�[�R�j���޵�41Ϩ�������gz��������ɒ7��}:����ul5z��g�@���$�/�%|$��9���S�K����J�rg{��Z�s֕8怾� I�A������r���LH#�D��2 �� �2K\����v�j�
6׫��Z���Ï:� �=H�w��d���$��X�3y�`��Uzg:���������/{�5��ۙ�&��s>��	�Ed<�'���T1w-a��}���� �%/�2K�2Wg_7<:{�z�o�@���-ٳ�y�Y�f��P��<%��+ ȅ����˾�Έq>���٠��u��5`ֹ�b䚙�`�tl6���'9��[=�~VC��"_IԻ'yz���çA�4�٩�Sz��&>U�! [� �D���]���;}Z�ݗ�}WOoS�����Z�N�Z�u�ȑ��o/i�j����=5��{[W~�r��s,*�0G:��y�z[��_a�8��b�9�N�� �|k��̞��W�]m{��eG�s>���7謃���'ځ��6wa����`�R ����%���HAU���Mk�6g���wUcs6�z�t��	ޠ� ���2E`�$_	0&�K�)B����
?<��3_R[X�u�ÇN�u{�	ԏ�r��.u���}_iԀ"H��%A2P_"�7�Q����¾�C:+��n{3$͏��};� A�E`��?H��I,q�Y�OZ�����*-�dk]&���#�\Ts����F-��kb��l�K4]^�MU���DNz��wF���� �(�s��}�Ս�����X緳�A$V  �"�I��+��vN�*�u��?'?Oƭ���N���:=	�q�3bH?n��d�^U�)c/o�|Gw���AJ�H�����խI귥�K��m���Cv���Y�khˍCª�P��g��{��Nk����t�F���y����r�_S��>�ﾺy��׷�+�Yn���M�V"r�I_`�X�d��x��z�uВ������A���5k6�kt�y^SN��i����=!�&�����=+�&	�+ ��?I�/�7�S��Q�o���n��,z-�Ɛ3a A���J�% �.��_��V'�aڢ��vV�݀GT�Q��ػ13[�d����7Ub�V+�s�X �Ar�2E`�$Aw�7d������N��w8z��߽m����@�ޯ��X�%|���"Η~=�tp�7ʲ�z� ��HV�������ܵ΄}�`����%�1�Yp`~A ~֐'}�� ��L�$�W�6n[�r�ٲ.��*�F{��� ���,)@"J@�%غ^�|�����A] �fP@���Ĉ.�f�ܫ�foiW���l^#�u�#xO8k��V�l�n�r-;snLN��ϨG\O�o�����xi�qe�sùV�^,r�3Y�k휠Vku�wow���I$�Ne���]�w��i�j�	R��$�,�_��C�o�UYT;�үv>~��'����΄}��%%��YPK<4ŕ��a��Vꤳ�t:�Ҭ9�Krp��@	tq� ֆFې�3#,�1�βP � �9">#3���{Wg�	��C��wr�JϽ~�^�a`������A��
��%�`�(Z��{1n���@o�X �r{ݹ�{Mߤ�3{J�z�6⿈"r��|��6��,Yݤ ��"Ib̔�a~�Y���ї�j�]�=���c�2�z�}�젾?>��2E��4�_!(`����+��t�����%��m�>�x-��n��4H͉ ���*U[e��mk���!��D,�A2P@"��{{0c"u��7szv�ߜ�3y�N�@�m�D�?I_I8�Pj����óf�	c�b���3�;w�����_���v�yo�kۖC�͵a�M���,]�ڔ�3�f��{3B��ݝϾ  =��H�*��
���.v��˥�B̟�8�1Ń�;@f��1	P�e�5��UTu�L]4�b@�o1m͘��',Q�Þc�\Z��Y��%K��J���Մ(�K��G3씅�KM����.��.mXTY����K���e�kv!l2!M"���PK:��Cu��&i����d�0[y�mL�eCE�Kj� ��M�MY���f���g���D����1)������]��X(l
K*�I�u���џ/���E�|��u�J@�D��k������b4�e�AV��g��?^S�� �{V���"�Ad��#/8ΙRq�fj3�<~��������ƅ�ҳ.!��A�ؒ�A|s"�U;g*U�5̆G���X?J%�XIB�LW�v�%'^�ڄ��T����qY�/��W�I,Y��ųr�>�7W�*��)�Gfذg�"JC]���^�3��P���e�kA��Я7e㯻1q�A�H$_\��&���������n��hO�U��chC�"�X����:F��[I�>���~94�Z��j�A���#z�1/v�b��Aª�p������C��4 ~�f>|��A!�v^Ov����/85N��_x��,�j�ւ?w��"�� %}'<b�{jӤ��35N�b'��*Z�f�㛛��u���@�]w}�8ԍ)�x��.�E���h=^hz=%!�ᙓ�7����|>�����MZڧ�A��A�)��Y I�A̋q/7)�ߘ�����VA �?I_)%����>E�M������N���R���%h �D���X�E�u�����] �~��9h Ȃ���5��m�Iy�,�w���E�c�m/1>?z/������I_!$�+m{e��ч7C���ݝ���n��Ck Ӂ���u��C�H��9o�=Ɣ�ex��6��3Z��2�cq]���\8�Jvu�Y�&�Y��_d������_/���S}����eU�%.bu}ꃭs��C�\�г�R�R"H��(#��p�tc"W�������5��n�I{¦};����_ ��1E9]'n|�݋9��N�AKd��%?�8��ozON�oQ|g��U���UW��V���4�٪��וQх�����|��NF���&�ӽ�Be����	�J�ě�O����l�Tƪd��"�:��#�Q�-V8���۴�P���Nx���b�]UTYK�W:�~ʾ��U�+���m��k+�u*��VFn`Y�hG��UO����J�R�{zJ|�rn���ۏ+�f�4o7(�N�u����6�U����s0ԭm���Ǡ���5Z�FeZ�B=!;Q8&\�ǬԄ�+�	�<����;1v}��J�vWV�꽥f��K��T��8��W+
����������T;��W
�3!�r*ͫ�t�E){�g��x:��n�U���g�ugv�/H��iʻږ�+1Ueօ��z��@�+.�6�� ��[T�N��%hw�7UU,����ۇ�i�y��Vp�O���؄V��!����d5�&]��y:0�<�����O��՗[��ʩ�a
�C��Y�r�}2�ś{�u0���M�{T����V%���W{ֻSzá�\,p�x��Tr�K��+)���\N�:�wWUQx����u�v��X�G��-�;��@]-��oF�gv�Zdi𪼷#]��������7���P�E<˧[��v��}�d��l�b�<�g��n)5]�E�ƠIF�-]��}.﯋��&���{�#��R�k`�*�J�z#�;�cS��j[�jZlp��x����I� ÔQ�qM)�����5Wxf'���f	��!�V�r��u��Ɩ��W��J�������P$�4����0��[X�wmn��ݧG�7hjM��;I��N�6�#�0JN�(�͒6l��V8vi)�8����Ф�f��S���$��2�֢
Aٶ�m�l��[�̒m��mjζ�m��[f�l��̷����u�j��6í�������VvwnRr�j��!i�p��G1�[y�=�lq�Yٳ�vڈ��L�8ٸ��qe'q�n΂464�m��c[[�4�'v�ei�-��̷"��Z��L��e���ݝb�#������l��\g[k9��c��.�l�4�;��m�6Ȼ8���K����Z���̔4���@��_>���W�v����Q߻��	�@"�A$_\�#����p�~���.���A|~�A}$BӾ��^^���"�c���g�&��}�TN�Z5w�jA��H��%�W�D��3�:�g���ٯ��w=2K�3��@��+���?I_)%��+6VjGn?�D��bV���9/1�S&u��tn��42ӕevB.�i��n�J��RS �ґ�_�V�H���}T����>l,�e=h���&2-�zꥺ�oh y�2 ��%��_�i~�21l�����Ծ=�b�N�>�yz*7$������Fz��X�%SͰ�Y��e�{"_PD%d��"JW9�z�P��j���,�ْc�S>�C���|���$�`�H�	nzC������m��#2'��l�����aޡ7�`���`���p�g�}� �*Y:K>����+�qS�ۭ��:��3�^Vl�R��eU�Ս�5U��4��y\7��/i�Y�yZe�[����*�ВH�Q����PD�Yl쯤�~ Ȃ?H�E���V��fW�� ��;n6w&�/ ���@����G% A"J�n�8�<I���j�7wQ�vW�J9n1ql��[��M���ș�nZ�i���''�	�P_����YH���݋7�&�|*oӼ���U�͐&����_��$����~"JDn]�P��G�^D3i|A#������?Q��f��{���A�� d�k���?_W�ܴ�(#�/��_����O_N��*�Mqc���#:� �r����	W�M>�=}->ʉ�@���:����{��7�k7�&�|*oӨxqYmP�����������d�A"J@�$�fJK�e܃%f��h���~��ϙ�f��{��] �PFH��(ma�*�M�-\VV��=�'?zp1���U�^Nھ��N�Ŏb�8Ҷx��)v�י����-)�=�2J���|�ݎ�D�!�@��36�K`0�n���D���&�*�clz���A�3Q�%%sr�]�e-#���)r.1��lg:��&w���<�n�"�9���;��З�P��a3��w&���i�u��h6��iu!sXb�Y���j5j�)]�ʌ����D�3bbQ�a���dq��k���,l�,��8��,��5	��0h�2�я��.����G].uh�b�	�a��]�-�»GVi���&��}b������`�?r�~��X���y�7r"�*�K��iX'��1����}�C�U���N�����Z5V$�ru���=S���g��\��l�1�N��q�d�/��J�������z�υ=�`�@}Hd�,)AQ�.���-s7cf3�[:V��G~�hG�QhǞ������l��"��`�+������_�_݋�m�y�7r.rj�'A��	��ٯl��o�;�舘�Ns���(,x���h�^�r1�bJsy�,��9�������֬~ؾ��۱w�nǹ���=���JV�@qIHaff�хf�eYQm �Y��UEV������r"	�B}�f��*��k������u�\�-��y
ȎS�;⛽�y�S�e�#�Yl�T�9z�s�k�[��x=}������/g.�/wTGuf�dH�U��5�=�[f�	U���;��ڞ����۸�Us̼U�c�?���\�q��#�O���|c^E�-p_h�|A#�@�w�u�-zrr�����	�A9��Ѓ�T8�s����o��_e�l�<�yUߜN���#��j�;G�U�m����F}���(������ޯ��/��b��Q��P�9�͠�"��g$���H`�VA�Yc9ENs��D�,�����>w��/����1��s�W�:Ƃ�3 ��k�e�Ddv`s+�g�ت�U����V$u�j���l��/%ui��Δ@��A���ұ�W�V������k��^�|����9N���?{fߺR}�f5���~�ۿ���n���=;V&ZШ*�8�R��_d��{g'^Ϛ�\D�����?x�������ߴS�~u@�ӕ�������fMϧ�����KC��V��U�H�A�F���sG������9����<����"�d��02�tk��W'�P���}����r.rn�'A��A��`��Uز�/� �~m��e�/�'��wy|���s�w=�T����<(V�ds�^;�昇��k���_��?6�X-�Y5�?_�X�,�v��O�k�kuq{��n� ���mg�w!���Z�����!	�A		-e2�.Z�0��F�#B(���jkkU*SrJ�M�o��2�"g,�g*Tg9����y�gj�v�bu}ܼ7<�o��A �ge/��6���A���''[��洂7�]Q��᷾�*^pk~�x�YF�?;�5k�-f����q�H��A�n���3پC�}4o�&{'�k�kuq{�_��@��[j�-��Ψvvr\^�x�Z����������wO�����1:� �1�-w���j��Dx�`0�3m�U�M�S�(��ݗC
���p���o7�fmN�t�N!�s�)�
�����p��������w��G�y7A A,�-�A7�������?T�G�77��K�o��	ZՐcA|~g���b�v���}��g�_��j�l=���R�]a[(Xn�J]]�0Bf�"�m�8M�Q:ީ�����++�"c@�~�9V��Yʗ�}����̪U,��"N;c�����G �q���ќ��P��.l�D����c�b�3�����h/���ob7�Ų)K��^��D?W�]�-�{�����U�M�4�״hc�Qh�Js���&���u�{ �=��7{\�yЭ��V�D�/�Ϋ��nŖ�z���%�&"� �yA"�Kwwj]�tɛ��M����8�Sx�k��[�I��ב>��(c�r�#�Yl篚�V[l��}ٖ,-�s�U{�E�)K��^ �|A�7b�t���x��׋����VW`���=�c���NE��z�;ɸZ:���}%�@�xz�w���9�������dj�WL����3]�q9a�?�ӧ~����#KbXg��	Uj�u($��C
S.-v�;Fip�h�u�$��72:�-�%&؂&�����5ͩ���6�fհ�]f�♕i�c�p#nѵ�&�Ԅ1�8�e��5�MLtͤ�Xl���E��Z�5��M\��h���\�0��Dk��X�X�i�[{+m�)*��F���.b͛ ���2<ejYs4Ԕٻ9)1����m����͎���t5�e�M3n���2m�A &�n#�t�h|����}�DAE�������xc�k�/:�B ]f�w�u��/��_Wʹ,�H�C?3YC����a��Hf�wޞ�W?i��y�|D��(|~m�x������ ^A��z+A�W�����˶�f�-��\����U{��rT��N�| #hYn���v,=��x�]`UI���=��������}�EyЭ�z�F���{��MV7-��#�w�#w �1��_]�F�y�b��	�Z�������sr�������x�-�`��=^�!T_�vc]B3?���'�T����c7h����vMc	���\m]�X1Əa�[̽����Ԣ/c�j>"�Ћ���#4��y�[�|���S��G��CLu�f���A�@{7.���w$g�*��w:��<�wD־���9՘����ef��᱓������U��]�Ȭ��I�E�(�}����|*�}u(Gd�?L����^�\�yЭ��V�dA|~{�xc��{'���|��G�[v,�A����i����:mWg^�g&o=���h���r�"�ʣ��#Gǜ[��#��?z��mص�9����SfC*���� �h�,N85��5�O���G6п�t,���}K}����l��g����{ż��*��[���`\A�_݂/��eԡ�G��,�h]-u�vΗ���[��(�4���Ņ���Ϸ��@����߸�Y���ޏcۣ/���C��Թ���<9CH%�_�_�7A����u������돣��栩7V�!���!���J�D4"l���i�HCܿkm��]5�	�{F�9�,g������Ua޹0W������W*5M��#�GV��a�RW5�(1t�yw�nX�C�s�$H��
�}�>�fN7���\�_��nOpn��JV�V�?P �����w_�v,�V�k�{�]wn�h�oF�~�K�@�}��P�j��{̌NF��	 �ȩ��8��"̼VA؂?2(�������]������jX��{_z��mt�eo1ҼA��hf�[��!���B{��}��F����a���MZ-�%-M�1V;b+��7l��waXVZ6�g��=Y�|%�߶���/\�}<�l����B,[�s�]:��o%d#A�B� 6�Yn�@�h�J��V6�D�{���	�}{u��mC��y�~{��~ �t�7m��q;��K���[A��};��m�����cX��!��ol�\�u��J��h���@��|Cnō�v]��虎P�A��k-��뙏����$��·��@��X#�۱�^�a�$��cm�9y����g\Cv���md��+���e�	GEμ0��H-0J��L���j�^h#�U1.�^ޚ��{��2��wڜ�|#�'>��r���V��Ԧ�CAc3=Yz���S�~�P��|,gP��-�`��+�ށ<�y>}6���e�+�*h!p��<�2�X���.��S\V�c��:�|��?�ng�ۧ�W�6�^��}�^����J�
���{�~����:�|C5�!�v��|/
'j���F�+��{�)c���N�~�X!�����dX�����+A Cm-� �e�FJ��J�8��l]mE9���7z Π� �|EڰAm~uAz�b�1�Q�1{> �H���A}I�[؇:�K�+y���4�^7tV�r�m AC@����~dQm�w��Жeq��@/fg��+-�IT�
�?P%F��A/����۱�9��g/�/�L����2����'�2'ݹW�.Aw�i�ͺ�U�TT�[U��v:��Zۣ[�q���&�z��ɤZ5]��YY�ףM�١���fk=2L<�	���v�XW�W�ǝ�8�V�ܦ�y�I�(��_VX����|��AT�e��r�RC��髮CFv�[K�q�.����}��i<��6]��:����2�����r��U�T-��yuF�g8�9ds��o�]O�|4Ӓm�i�,Ř����ld0�c/2��^nI�誶���$�+�o^:�A${��4sV�G�Q68�8�ۻ�+�UTNݕ��9WcU�%�V�'G��}+��[t��S6��h8�ME7EZ�2f�/�U��C5��xQXH�dK-`��U_��4J
�q�cI���*m�LB�fd����Х^Y�*�I�+���7�8z�;����47D+�i�d����I�}WJ��pU�RWU�.�^��l��j�6�6�wwN�?Wf��h�)�L�R.(�飃������ʮ2T���:�3�8s6�2��Z��˾��)�|'�ݵqłTxn�\�Ҙɝg���v�Z�\B��չ�:��&�+�m���U�Q�*B� �aj���j]m�su��젉Nm�x���01��iU!j��h�'�(�E8{��:���1Y��{+��UG��eѷ6C�*ن�4[μ%�9�ٽ]ծ����5�꽦s(�uimu�-vw0�*���nE��+�	����+�N=#6�^�ϕF�����4J����2�elojz-�k;u����(����eD��e�g��:����m���յ�Γ���[Y-c0���vp֐�m�6NJҲ����lG1��a�GZ��ٕ�XY���2�K�2�-�rM�8��ʹ�Y�Yͭ�r-m[���y���9,��[i��f�#��dfu�e��[c�3��Γ�k�}����쬍9mZVE�n]�6��lm�Kwfr֢̳-4���؝ͬ��X�d�#Jmݔ-,D��k��.m�]y�9�vem-���m��u�V[b���maI���mv����Qg-e�im���Xq�n�ʼ�^�6|�/ZmGYŧM���Lͷ�2#kq�[l��F���Y�h[�mf��kVZ]���e%�7�g)о|��P�3MJ�L��-A¢�cJ�c�[r��kFev��mF�Y�\��-�����i\��<��X�E,��P|-s՛��� �/T�liuv6pB:f�tce�R-Rcݔ�j��V�h�o�[�W6��ee��7:m0h��J�Z,��l[�.�+�A
�7@�<��5l5�f���fe"&��`<rV:���3e�@qZ���	�֢m&�������K.m[F�R,.���B�\����X�N#f�d��с��г ���vuYF�+�R�(s6�x"�Y�eYL�fZ�g@�C[�hگ��5i�{Dq��AB<����N�X�6
���yu�JY���-9)�oe
M�xv���B�[�[V-�^���Rlvm. �զqu�3`�jc�ZMLj�+�iXb��Axt�(�D��i�Г���\�Y�����l�C�e�GBb\5�+@T������%4��x6f5�#Ř��.e����5i�X�m�1�*��qp��eLqt��kX�6�Բ�R�w ���k4u�a3[�
ГfuQζ-Bk�vٛ���Ee4X8ƈg)�nj�1�ͥ��f`MبU%q��P���v.؆s����(mb2Ƥ���[n��`�JڠJ`�����Ō̈́R\d�1�퉉B+�cP�AIuu�FX��1�eHض���cek�e�X<�X͋R4��������(�CU]60C6RƶcW�,	��),)1�%h�dj6�fC��V��D��71�bX�X�Zq!Irk���{88�-MA[@��n�h��(R���u��h�ls`kp���FB��-ׇ���n��L�Q�\��&�Ѝ8����:���uĠ�.�:f�T�1k��&���"�e�$c�h��\����%��:�pK�m���t�-p�&���ڪ9p���r����Ɇ9�!2�/��[JjKDl+i���!���Gj��e�c3�<$!�5�ƨ1����r��cL������cǔ�b���E��%����ŋ	�(��Ld��,^�L2�\��x���4�t���e��Lx����F�3b�ˢ2Pź �g��V��YYt]*`�X���^��h�:`ֵ��`!LqWR�#�IZ�[��1�3KR�!��6!aF�+�qO^y��	�k���iWLF-v��v�rS;L60nnYa�f�#���i��я����	su;)c�bE֚�Wk*Q��BSJ������ ��5z�ݜ��"&4��4hyʴD�F[���E��-ʴ���~ײmV�_7F�#�g;{��T9��ܽ&{fJ�W�[u ~���nŊ����\������:W�C�M�,�WC�:�}�pw��k�76���E�@ڲ���1����s?y��ߤuJp���|�+ ��q��|@m��֑�mw��������7�?H�R����M�������_P@�:W{}�Z���`;ڬ��������n�??i6����Wg��=�=���{X���3���#	�:�~!�Y��|��.q,a����tn��*[t��!�����̣T�1n�[p2fEc/U������X�=Js����VL�����6�w�?}A�[HQ[`���(W�6�Yn��"Ce�Rŵm$�o�JQ��Cu�*�T4�j��m��6�J��Y��*�UacW�������jUQ�g}Zc
�q��{&�4��VB��~��ؐA��06�ך�O�����~�A�_e��h��
�@��P'#V-��?:������9Ѝsӻ��7S�Vs+�h�u�3@ۻ[�ǉ�yT,	� �r�7r#q*����s*"[1�^�%F�,Yu�=����w���/���6�_źΫ���wu��y'���X�\�uc�!�s�"����A�Vhp�r�T�J_�^"�v(����aFt�56��\d�,�8ڶn�e��Q���{��>��@��$�>�����ݕ{�\�x�E�+�;�=i0�^_�ՠ���B�t �4�E�~�~s�����]37����˫�5>~�AQ� ����>Y��U�����ş:@���m�D��[^�j@�>���**IAj�V��~��ͭǫoUDtt��q�����ɮ���M�5�sQ
˄H���ב�S��j׆QG}��������]��?c������H'H�n�~n�������u�gmp �' �����N^U����շ��<�0�X��ܼ��wكΤA3D6��A,�-����{wKZ�����37����e���+b��|���ݡ�ѐF^���;`�Ĉ���~��ɍ5��ԅ��R�@գ^p͡[��Q-t:�6��7�#����>�E����_�w�pm��9��L����a�@>?M��A���Р@-�`��1�aqc��G�7�!���݃��4�a�� ��,Yn�mW�d�]L_�i�����dP-�[A�q`�)�ۗ��w��u/zL�]
�+ �G�_Wŷb��D^=�y�9І�,���Է�vc~�wU!Ӑ�9����d�Kyx=�_xDղغ>�׆.�[��f�۫_zt�ZZ�v���.;�fuvy>�gx��Lw��|�S��=o�����^����~A�@��VAm~g����O�����ٞ�}4ni�^g24�F�A� @gu�]Uγw��֊*���)�[7.f�W*�B�:˝Xծ4�9�^v����	C�Ҷ,6���|[y�t+_gOk���\��)s�s�s�M.C���h7A�!
kwW���́WK={�޻�>�8/恛]�[��kW����`:�����>>3N+��'��3����=��b�����>&�GmwD>n��Ξ�W��R��-����ͮ-��u�������5{7~���3<�ۏЬs������m|� �W�zޯl{*��o��W�1i�V܊Z�����{�����,��x��g+��e͆��Cb�u�Z7C3V.[�ݍFPŹ��⺚��jw?�uP�R����%[MP:����iM&�[4�X��Փ[�^�2�Zf8�� �n΅ٚZ�Q,������Lƻ1���h��YEŲ�c[��pŹ��\L���P̈́����fm�Hƫ,G,��{7u��h#�[3��汴h�፡Dkj�*��A/V��U#��D��m�3s�S-(Z�Q��!���L��j'6����>�h��n]k�%�F���'
ǆc͌�6"ɚ�2?AB
3s�,r+b�.�]��\�-�2��
�^�kuNf�(���6���оy�r�6b�G�Ukcf/��������}�]��-�`o;��%�O���:P���7�(oEz{|;n��yq�X6�&9�L��Pm��7��.����u["�YU�뻛֝n!k-�1>w� �H[��h����wPm��t>n�o�� &���t6�ۛ�o}��R���%7_6��m�B�V}ީ\��B��],������:莚����xD33��LXQz�X��J�T���7�7Sfg9��9KF��'�{���##�ש���rm�����=�=8Sor5(�"�Z����k�����Q0"��p��z�
���&��ϐ�OI��^]*Z�M��������o�e�31)�Yv�y��|!b�]�-��t<+=ǳ��g9�&�k��-��;dBn��u�tm|��y+�v��u:��_n�f���]��\��/�����i�	efA��]ӵû�|�v��9��9KD{�ON���O�⟕*�f�ނF����o�{�(�d��������s���M����?m��"�"*�"��,P��Pi
��`1[�*7R��015�J��˹�Gm)�*�x}���ot'�M�8���\���|͏_�֡e��֏J)����p�^}�{���]�3�������'�xL��M���+)�`z{�4`�B�	��n����yZ�S�X��є��4���T%�v�7U:�ފPʥ�[�����u�al��Y��ۉM����c�!������ݮ
�t����9��t&�m���z���3��-�Ϲ|�:Rzo�k��.�J\��@���W�/W��n�m���s<��@:���g����B���zw��A��i�z��������%��9�EZS	�lc�Gm5�.qp5a)�j�4�Sf�G�r���U��q�����y����=�C��;P���5.{Y�S���m|�y��Q�L������X�������D��5h%�*�<�7g8�u}:�m���n������9S�7sw��\��T�vp=;�e?Pm����/�E����w���+��'n�u�=;�����V���i�8�����S3�q�&��][���yJt\�#Y�lt�˪�ב\�ē��ޫ�F��DV�m�.��a���3\�y���m��u�t۫�%?]����}�W7�7�_�M�R�o���tme���7�Ȓ�&��t�4l�*Me��8�Zk��-oX�.#�ŵv��-w�j�ў_�<��ɺ�7@{n�J�����|w{�
^���b�}���rm������տz��������۾�F��N�<����c�����r�go���|�owu��u\��o=5����딻<��#vm��7:Z��Y�W�[M��ͥ��mV���oB�=z^-҈^�隇�݆�7_7]ݛ�zpb�����N���5�ͮd�����n�ol���݇|FіM"���C�vX�/R\6���͝�)h%^�YAn���7:�e+ع�o�Q��D��wy�F|���:�%(���	-�2��3�6�^��ѐ#p됃fˠ��.f�Z�/��O7�n�3�mE�-��,�F���,V#-�W=��n�^.�VWL2�#h�avXVS�������)��2��M��/V��T�3�Ц����Ysm ����@i]���Ұ��V���1v�)%fjKl�P٘V��t�E��	C^%�K26�؆��m����F>��~��1����a�G�bl���!s���+T@��݃Z%L�YkT���}6��6���}%���v�k�yu�]��xC�֕�����;���@7A�����국w-������py�n�F����.Wϫ���IgfwN"�St'Dt��}��[f=Zk{׽�Q�r�ms'��_؛��|�^���S{��,���)s���K^{˭���Z��M ��3Лɺ���6�b�{R���(����o�n���{��\�6�6��n�G�����H̤��2���	�d	M�����dR��Y���R�J2�o��﻽~�����RN���>Rj��1�x7���Xj��C|݆��7SF����g�v���I��{n���5��0���CQ�ճc��c� ��$_��L�TkU
�QGNv<�)z�j�	@Y��Sy���w�߽QOK��D���[����mY�/�V^V3���}=_6�u�l`�Uy^���N���y�|.P|�Ͼn�����htǹY�� ݮ��ևI��N��&��鎑o�[���m�^F����tu�m��CՊ���k�I����)y�]n�g�h���m�T^쮞~y�ޯ��[��um�P�Z�a\쐣Q����⾰)M���+��]�N�4�����<��)��|I�ٸ��>�����m��Ʊ�/y���ix_��|��پ�G�MS��:O}{@tk���{�y�T�oL���t�A���K�,f�-4_�X�tx�ӳs�{� ����Y����=О쫵k$��+���H��z�M���3H^,�T��o�r딯%G����sh�ص�z�8�e��(E� š��آ���r�I.���L��㷽��eQWV�q��8���\�T���vٮ̣H�VS��T�d��w�r�T���+��k��֪o*<&kx����c�ث*e�u���Ѕ<ͽ内gJ�u��w�*���Ƌ���]�2�M�s:���':
	E�V�����7c.T���w/�q����$L��f%R��%k�Ұ5�sUd��Yw��ِب�:Y�^�Y�l���PYg[ڽxjVf�q�Cx C����ov�F��/EP���ԙ��*
1F�̸iy��e��')���r�*�N�z�i0nK��n9-�[�{�![�}��?���2Py�U�u5�fEƥ�sB�G)��P�n��*�AC��VIΝ�$���*����SJ����v=�Av
��z#�!�\�#%"KB�o*w�nWpɝ-j9�}������Z�K7�L�4�w��D�h%N�Y6��͡-��w��m�Fm��V�%׎���4t��X��|ڡ��Ӊ��+�Yoީ��#1_h8�>�f��������Y�{G��f*���>��^�˛��"Z���ܻ^��qZԁ�U��Mp���!}Z
�C�72�^)�S1z��u8*	�杬޿�ߞ7:�[9��}b_r���Xt�;Z����-��N�a>Y']�A��O�7���i꽰�Y���/lVJɛDL���~_��{�~�Kf0(�m��m�mы5����o[n��ֶ��6ݝ3[v��f�q�9�j��2l�e���̎��Ƿav`�u�g��#��ގ=m6�6ݜaY�d\�4�9d�6ݶmgN\����H��l��b��ݦ�kZKc%���&֔Ͷ�G-����Vڳ
��;8	��fV��ײ�[[��}�N;�Zn�k2Ӓ��ls�����ٸN۴�ݤgmj��6��Z�q	m��h��
Zn�Z8m͐,�,��޽$rq��S��#��'B�m�-#kPD�sm##PM�rDRfFX\C��m��.Vve�{��s�e�m��;B9���jm���o<-ي�k=�m6�ұΓ�K6���gN�a-��b.9ʹ�Yne�{zpV����lf�D۴�gg'�f֚nvn�:tt��m�4�۴r��̴�($X�TUDQ��ě�^�y�]n�ef������_7HyT��9���`o�|�E�����.ξ���|.6;۽g�)vry��M����m�Z[�7�6Oz���yF��['����n�u �?]���T�V�7b��S.i�k�
�P��Z� �n��m�N�.�8`|��&���o>n��)��K���t�=N����K�o��M��w�L!^]�#��u�[ps�{��1�%W9�.P}A�b�me���Dޗ��B�������ͼo��fEP��]���W�w9�I��v��|���v#H�����>����|�R�=/}"^��s+���vM���e�2M�����t{�9Wb+�}T�@n,��eu���]X���V��o�l����<��'^�F���o����Ⱦn�n�m��߯7�jYB�_��s��)��*��}r����or�<+�UFmhȟ�6`���%"D�tNIjn�UŅi�n%!AJ$��$���>�\���}v��wf�uUy���k='���jI�οWY�9��y�m�;)�����wa6����{:f�D�����g���|���Re"����>z�����'�
B�ra�{�j�",SÐ��|� ަ��������/�nlZ\�L�z�}M�;�u���{9V3�{����U��%��5��]=i����9������^���zKS���>�}z�����t'{�[{F��G�{��ub�z��hi�P��Yζ綮h��U8��mK�;�8<���f���g/���nǝ=͊�|�'S�3�Z�Wu���M�(�̗6�ʤY��ҥU�7���4� iPW��h�Bx����,,m��SR䕮Vj�n���ƥ(�V�ebSm+]kl)-Z�WK�P�v�����liIf�z�1��+V�&��K�T�X�V�X����"�nlB�;�Ò7���[B�8rMj\,�F\ۮ2�j L&l"�[�L���.�i�G1\d�cu���~O�������f#�R[+X�k�Ra��A�q�iX]T.�!_Y�Eh�6~e}���ۺ�����o�S���_u!�V������|�t�ڛ��%_H��v����~'������<>���t�1���.��YA���{Jn�k��t���w����y��(�3S�޿־ަ��i�|!�mW.�y�����|�T۞/g�_���؟�	v��ӥu��/�����A�l�|�V3��3rc���>����OI���tc	����O���k(��Ԛ�F1΢���̴4���#w3\�e��Q���Ut�o���e|�_7%.}3}O��෯�{r^OiR���~���|�A��6:�x�!JY�]��4�7�D2�ˮ�޳�-ݫ�$��S�p�I\{��t��*:��I�y�*𡚱{:����,u���<��(	ǵO�����LVpp��\�7��9Ӻ���|G8������|���43e���篹��|�|�i�</(}Ѧ��s�OC~ʣ�{k=�����~R��·���m�fZO�`�y�n�m���'8R�P*��yߴ�}�oŊ�N�ᒆ�6�����K,x2��po�}vn��(��8�b;u]�]��ƣ.�Y���B8��D*�T�7F����_�}�������y��i��=]�ǹS_gx��A���}��k���	yps���){zc~R��[������<���N_vWϫ���k��Y���P�7����Qwt��-v�q*t��kL��̎]WP|.a9�Wm���Yɜ�Z�]*ZҔ�UؚkY*�)�D>����-��}����N��d���t�ڡ��+S(^��jJ��=;w|�o�u���O��AT��l7A��u��݋]��_�'n7w���-��W�+�[kz�w�����>B�'�|�v����l-�,���C$��F:���Gj�(h�4,H��+6��޷��Y�4��l���{_��Y���|"�^rk��`{i�/���}�o���}��.j�/ջ�vM��Z����+��=yC��޺5g�gq>q߽���n�h|����1��Q{�������o�\Ol�|>�hoW��m��BƤ��-�4�����7B���8���X���d��/>��ާ�u�xJ�|:���kz��b��;n�3����Z���L�W�����O[	�a�*.����U�^��#�����O-����������.�~qwFڢ�\��;��^y�_^��L]w�ӽ���ɶ��ηnq�0r�1�LD���D)H��R�cʖX�k7�ce�iFm���/=���8`|��og|�O��ǿ.>��z�e�+Ֆe��#F����Ң4;����%ͼ��7A���b{d{���Hg�a��o�oi��=�J�z�pN'`�����{C��n�mގ���� �zr^w[ұu��޼���m
��9.���:��Z��7��꞊?dg��^�C=H���O/�܀n�n�m�o$���K���y��{��a�bt�|2Pޯ�h�\<�O�jy��g�l��L�a5�nګ7nv��z�]��&��]�Y��j���ϲ�(�.]SNx���W�$�-%q�W��+1�-9�t�����hcV���	�\�-���%C+)4�A�&��ں%kbgh1�����u`J����e����MZ�)sɢ���K��kV����q����[�ƴm`"u�G���B+���ra�B�F�H(�e0�T�L
M��ɱ���4U����Fʶ숷[6&n��
�$�e��k0�9*�h��c�Y�J�6f�JX4CGd,�G2���?Y���甞0��fRT4��T[f�fH7\�[�FZGF�b.�b�̿��}��t���?_����[�V��t�V�N�Q���|��A�����޼N��ix��3܀���foE�[=�Y<�x[hoSc��C��_c-f2�v��u|�o>����p*�r{�rN�����xd��M��t�3N�ԗ�����m�%�'?%�ֿU��];��,��ڢ���^kޠ�@7A�m�j�@�g��~����[�̓��n�m�7�|��v{��ｵ����]���D�2��Gjk(���n�j͖�@r�dKB`]"�Z){����x�S}�sӤ���buͳ]*�9{�en��7_6���)Q	��&�2昲�t[�g<Vc��7f=������r�N������O��2K�iHF�Q��곸r;�gνK�ﯠ���c����aL�GN��������c�}1�ݝ��|k���ֶqS���(w�6�y���^�>ަ�x�}(o^<w��B�x��oW��ov�d�LN����UF���������y�������79��Phf
NCZ�.����
_���� �/���k��u>բ�(��Jś�`b+��6:���Y�
ʸ1`&�gg�XE��&�ۥmf�m}��M�u���{ܡ�gl��������=7�s��ަ�����1�.ּ�*��s�%o�=Y:{��㉉�<:oP���pwdZ��ݼ��n�n�e��zR8��{*�ܯr���hɤ=���=�v�42����/���X�ep���)BؗӅς��+5�����ّ������)־5Wؤ�~�=��7M�]�����m?d|����=o{ܡ�gl�����@Wm�uW�K��M�����ߊ�V|��_�e+��*�Ot�q1:�{_oS~����=yF�������U]+�2i��\e�S.Ŕʣ�e.��t)k��?�9n��r�[..*��$�Ѯ/O������~���<n�h�d�7Cs��v��>�'<��(s��,�{^�ΛX�(��
�RW�:���t>o��T*�r��P�)·��:g�c��=�����n�n����mym�Y��kcw�~M��qQ[�!'8ު�9B�	?z+��" x�Uﶾ�y,m�#�M�Պ/y��lS����L�����lI������&G��b,ܽt�{5���*�yY{��� ��σt�������c��7sd�����/����6��A�m�c3|��'�{"��˴U��2RXE��4��$���12m1c��423-e3j����n��;��U�Ot�q1:g�0�TH����s���ۿ�h����u�����d���TV����������l����*�r�n���L#<
��_x�����/����hm�Ͷ��C[�o%�7��7^ծ�N<�e��Z-�߾�Ъ�|QnwM*�5|'Su�m����~�>�U�v~�y	2�<�z���U+�;�����@7@7>�,��n��î��u�v�uF\]e4}�!�EWp;%۬)}��>��22F�������l7G�ܗ�A]jK�n��%Y;������pc0�(#��^�S�U�����0g�i�,��gTcLo}�r�JXy���v~��U�vJ��I��KH���؍୲�r�w����͛�0$_cM۱/7��ݮu�L�����]�:9����!Ջm�\���2�a8�k�p�Ү`Z��m�[�*����f��t�67�<�����Ņ����ޙ�*�H��:��[�`�����f�ɇ[��F�Yg����wt�"�ͩY�f�S��U5ds�VD�*p�A���ǜָ�δ�7^�mM9;;:�J�;r���s�Pc"����A�f�iک����x��R�ʆ�w��k��l#U��w��:�lm��t�		��Ve��Yj(/�ۥ���.��Z�NT�Q�ݼ�X�evTW�&�)}Z7)�j��\�N���E-���)S��N��ݩ5�vM��=�3��o�K)p�6��b�������U�*���7en~4km�&�.o>�/f�Q�1��vV���	-C.o�k2��{�R��%�Ir�g/r�JKE����:�:j����r�"��>��/9J�y>���ݺ��\����l-�y�7�(�̲���ɢ�˓�3���wX�V��Yj3%	r.�ze�]vܖ)�ů^^�wu0�ͭN�5Yv�ݡ�mWx���wW�h?G�4�~��Y���O>�=[�ݹ��uBv��y�����ߠ�:�������nٻ�g7��<nγ �(�:�f�,��m TGD$\�h�t�1�:	�.�(�XJH��V�';۬��6Z�tN9��)���;+$-kI�KnӔTGekl%(������囿'Z�Bt�Ԝ��;�	$���m��/0����$D3S��s�"Ve�֬ٷ,����9ҝ�9������Ù��)���NkF�9�NH�:�gl�ӎ3G
+-:"v�h�;�Z,��f:Js��zq\��2��@R�6�NH���}�r���m���9Y�!���˒.S����gmc�fu��On�f����''��"�iG6���	��m��gn��:�m�m�˾�o�E!E��nܗJG8��t�=�B���K�{Ѷ�
J^��ޟ��LX7t5ːf�^�)*�X:�0��\�)�1.��=��-W[`ڌ*Q&s��d��	\�����Rl#��Y�ce�v�l�*�Q���L�;b��,�<��6�ɊQ�:�K-���BXV��x(-M���-a����u�%���M(I�nLpҸ҃�4�J+U]�p�.��u!p�e�e,&�HێԲf0�V�VXギ܍aY�1j��Kq�I��|%7ycA�Yb�*]X�@b�*�[�i+$��B3l�5���L�P,�7T�ui�V���#z�*�aYV[��0�9[ם7BE��Y�H�Xыl�6�l� �GJ9�6��6�6ǐ�u����^���F1b�պF�![`X���m%�*�:	E�.)�r���YdL�:�$��:�SeW9�T��ff���IZX�bX�2���o;�f�*�ѣ��]Qq��lSuKB ����Ե���] �;� �v��f!-�r���,!��/j�B5l5`����d�3��s�C�e��Hk�s��Ji]\�W\�!��6 ۬�I�6�4��Ƹ���
�sU�LQ�wf��J;����rH���1��KER�vs�� �6"�
09��ftYp��"Xb�S\��GL�$%vP!.[�	M)�"B�f�%8��b���A�(r��oc\`�Z54�Bf������uQ��@��K�H��#��L�,f)�Κʈ4��k�iK�*��t�͋����^ �k�J�Q��u*���JV��o'�+����iVĭ�Ђ��mi�Q�ĳL���5�Y++��kj�vZF�3�f��E�;s��7\R�b�J�XGbӒ�u]M�g
���t,Դ�&-tC��6���Qq�6�3��pf:
�͵p��)����a%�Ɩ�sX�6K�F�9�n�l[-{kT�PMo9\LY����Θ
�ri	������#B�P�BaIV�hҲ��\�m���Z�0%�Y���KM1��-��;j0J�f�hsB[�\�UV�cEa��$;i�u!��m&�n����I����\��3�jZbf����r�ٶ-_-3㲻U��7UB���a{&.�Fl!�Ț�:�b:����Y(JF[�e	�2�f�-���j5����͵����1B�IG�ҹc+�)��Y��آ��)+CQt3u�6�L��ntb��ᔁ��cbJ�q�w�.����²��%ҋ��?}&��O�J������Š��^�0Jƥ�B�jen��8`S��<�wr�nV��ד���N"�4V�D��[�κP�����].�������q��/���mf��S��|���}z���{n�n�z㪲���麎)�6p�mo�RW�;���=x��;Y}���sգ�&��;y�tY�Ȼ�W<�cn�������hs��t�|i��A�ם|����o6�MǬ&���7����cDөlj*��`6L�٘x0�b�AЬ1�l4ڻh�d�f��\�D][�L^:�����$�և5���GC�]�����]K�қ���v:s_���l�8^���ꓗ��[��J��P����+������r�4k	˹��=x�E}�$�vw^m[��*j�[o�.����=�Ǻ,�d]��<�}z�����ްz���߰	������M�jM���/Mf�[�چ��k4��6����+���:�_�_��|�C��coC���12�cs[>�n�Uyj����{��3Z�؅mOt��'��fE�Ms��k�|�|��|���eX���Eu��D���G�v�Q&��$x3��Aل��\ٰ��5aL��5h�@�?]�p2��Պޛe���s�l��]̓�������~8���Ɲ��9��9��|<�9m`�_T�������nC��{�Vﳱ*�v|���mY\�S:��p�lȱ%������R�ufV�yR��;��_ur�3�"*<� ���*)�UӰ��A�3�ea�X�jPˣïor,�Ȼ��yK7�sn����>��\�*���}��݉�;}s>=אvvO|�<���� #����k��=���� �%�.f�4|hXa��p>�r.��d垓)h%�GP��vE�J����A�ٮu�J�t�st(��vkVٌ�&,w�����z�m���=}��{2�q+�W�vr{D��%��^ϯ7��m�7@1���&&�v�n�n{}s�W��՝��=���o���2
��}�C��m�m�[�k���bYì�zwx}�@=��|�|�F��Beƫ��wP~��t/�g1�y~̩�J��/Z�K���V�2�<���;w��]�&�ۡ
�yg{7d�cWpQ����*x�)y�B�F�jU��Me�~����z^z^K���:��t=�� �|m���g�����QܬM���O�vM�Λ�������'\r�}�F�ՠn��ڢ���bG8s0Y��RT�4�ji���	��V^�(�[��r6������zv�Gư��o@����oם�O.|.b�@6�σt8gRG6�S��x�|�^���ו'�������m�>Oơ�N�]g<�r�}_���q���3�߶���8�u���+�=�Pm����ZÖ++�{f�˯����C~�ӸZ5Y1�ށ�旕����f�h|��f�;�s���`F������rN�Yٞ���m�뚦��c�y�b�w/�C�RxƲ:�]�Ǎ�kL˄u��飻�m���c9��%s�T:�������
*��g76�JŌV%h�{؈�FVG��8S�K�hY��)�k��K.r�]���J���H�!n��4�R��
��Jm)[�i5"�����3l�s�6%�i�j�-�aHJb�Yf��F6k�u�`�4y�0��"���\^Υ�[
���
�3�k`��Y��	`G\�vV#t�&���˩��ѱb[��٢�,�8���Y�g0�q
BW����27���	��*K]KJj�٠�U4��v�W�*A�+Yt"h, l�E]�J��)R4��s����|��ެ�c����Ê����ۿ�k���u�V�^��vgx��VLF�m���8�n�xį'����_鶀o�*�/#ʠog���xN�}g6N':��[�9����������v.�pj������Z���o��-���=�y��gwkx�~�M����l�Z
�Zȍ����=��i/Y���u|F��ދ������x��ƅ �����s�FVnxڳUX��+A�] �̖;Lpʭ������n���s���w\�9׾�p�����G���_7|�M�no�c��!j�})J����C�1>r[$�g�b�[Ψv��+<����d����z�fq�]�YB�%I�̺Ã�s����V":���g��e���z�G�Og����'9��M����o���e��(l�5�t��niu�5حߋ��r:K�����%|D��ڞ�*�c��1�1��u�h7}v�~w��q9��/��rUQ���u������_7���e-ʝ*�l����_��dއ�L��2��m�����OTt�0����D)�MR���qm�!a��G:3F2И�]��l=��bT"cxg�Gױww wy=��h�.�z�}����kl�]��͏$���������V��mug�������v�~����q7���6��[[���1D-�}M����^�5W��S��4g���}����X��<�D��۰��6�Wu�6 ��um�z%j���\���CΜ�
O�೷��5�';��Ӧ��ܦK��k�ۿ���2�w)�������Qu����d>����+a�S�&��Bu|�_7_7A�sv��:Ϧ�E�GZ��#�q7�޼k�t�����1qT�cC4\���`�P�?;�5�um�Q��Zce&��f��0����SO7���޽ɶ����~�3_�l�.���sw�Jo/�t�k���[�S�k�M��o.�'SR�2�u������M��3HP<rj��W��z�n�k��<kBz��+�7Һ�y��vw�Z��rm���Q#�����w���Zk_��7å�=�Yh��c���ߵ��g���Y�-X�g7ĳ8XC�Q�U\��u
�P�L��6���.c=�H���k�K�����Wu{��/'�7C�����Wm���~ź���K��0W����6���;�D(˺�Ʉ���l�2��\�bW�(M��yK˝�qia[T�3f]5I^^w�}�����3�rן�Gs���N�d�&ܫ��W����]������I�k���>}C��ݝ�����ٔ6Pm��O��{�kt��(v�|�w�m9=`�(3�/:t���3".ww�ݯ��n�n�m��ݵ�z������D�)ro�]���;�L�|-�&F��1W�ڛ���m��]��R��Qf�?f�K�,���������k��o�|]}���h൙��'�r�$GY��[$W�P���S�2��T&��6�B���&u7�D��W�m��C��g�R��<6�>���H]
�n����kG)�X��j�u*6��ĺ1�7`-n��]"]����
�� ���$n��aBܠњn{Mm**�ܱ�Bd4�sLl<���#c��J٦��,��E�j�jM\Ur�h�D�8��Ұ�2	�`�m�B嘪�[M1F�<�	,��
��]fܛ]hPj@�l�"�65��k�s� (:�1��3�ؘ)������4�5��"��L�6a���5��;@z�ff5�3j��J]RH���N�7@6ҝ���\3�D�c�;�!p�<OLo@����U��� ȂI.�JD_��v�V��o�
���K�"@K[��K��.�0c:�_���=FJ����g�c��_cо��"�ř)�D?d;�}_+�2R�瞎�]�c��|&�$����E�ȂJ����Z/�[�D�܉ �̔�m�I�>�������	���A��\�^���I�h@���#6D�$��% D�M��'���ʨ)�l��#.��D=�� �k2P ���#��fM:��+�xh��&�Q�b����r�]�Yh�6�mR9��,�ɣ�
��>���$��ّD�"w6��w��/�m��|2��AR�d�"��(�x�ِ��$_=9�iS��3߉�ۓ����[+:ą �ޅ��md�I�.���"�kx��B:���\D��j��V�]z��!5vvosV��'����ޭ��;>����|7{�����?=h#��l.�~��LSR'�3�B��D�Fd�fb�|s$Du�IK��W���7�7^�"���~?l��=_)��}&�������~ֺ@�K�د�9�$num���ۣ��e� @7q$�1��DX�Eo�_���� �d�� �"*��e�BNW�{j��F�E��V>{�?c�;܆�%|��?,�z�.�~׉P(U)�FƬ�U!�Zm�P��+-v�Vʘ`�� nuR��/;���X#�e���P�{��:�C�vd�:q�68�Ҽ�=��b�������c��/��PDb��{�DSإ���D�@���}�۾�N�9oFnr�Đ@� fe�>��D-��gP���@���V"D��@��߽����p��_y��iTc��SY����CG��YJ�f�r�]QS�w�Wu��:R�v,��y��X{�fÃ�s���NgVU��*�[��GT�Tu�s\�d�HQ�V��U�[\)�r��J굽�f+Q�����V*�9��7X��\ɿ���Pwp�ʭ�#�)f��v������5��(�)U��Z�D�K[����7YM_]_m�MlR�Ec}kג�/7DE���y���ڱ7�$��7��9�s�6�ń`o{��B���_H�0�v�<L����j�Q��^�3Y��eUW%�W{���Q�5l�4�nn�Od�'d��Ъ��x�Ͳ�Z"+.v����He%bf��Q�;\R]�ӹ�YAb�u�oE��+ ��Gq#\�ʼ�ZV���uXCc���;n�s����{�SԄ�7]�k��rVd�D��!J����˭sRfN*�eV�Pp�G��x�WS��.�'14U<JP���c,ku/sl�ڛF�1Pܒ�E�]b��+^��u]�U�U�&�=�f���юLW���9�o��b�b�N��C��]y�4��f�絒�X!m��J�'En�m��8ο�o�k3+�@�<7x�q:�ߙ�v��:_Q��{�n�X��򧗷�N/!�N��;�h�W4Φɴ�gvL͖଺��(KT��<-ov��R
�95��mm1�ڔ-v���=���[]u��_L�����j�����&�պ6���ܭ&դ�kX���=�uћi���y��
���)x�$�m������+;���@��ѺKm(�%��9�����)��9�Y�������[D�$E9�����Ф䊇$m�qɑgI$�l�$�:v٘���Q[X! ��6�k�⶷D�9g��gd���qDmے�9��V��Hs��lI9N�r)"qӔ]eh@��:�m�\�Np�����;qFv�NvZ ��C�ғ���m�-��(��9 t�
�(p��B'��HN<l��qKkrQ6�!�rt[$���m�ry݇QA�;�e�90)�"v�'%��'%Q�d�kQq8i�vd�e�۳�2΋���8�V(*SBU}��s�+5��k
/Y����\	��̏� `#3s�y����}����GfO�fH����<_��&�ӈ��c�&�%|B�'&�o������tpύTH ��g�ʐÁ?@���2Q�f�r�7�8]�ǝ]z���˟N�~{�Ku��D���"�`�{�����>_���i�D�&�`$�[�-�Ht&2���2$�\Fg7��&Q�*���{���?�ỈfJ\�V��Q},@���$_��4Ͻ��P圂=�$�Ff ���D�.F����t���=%���/؂���)<{�/�דt��C��MfJ ��D���m	�ڈ}��'>#�~@�ߨ AK�J��mn��Yݏr�Y�������;qo�f�@�r�H"܄�_��d���8��~A��Wgڱ}���l{�	��Ar���:;R%c����H�����LW��먪�Mq���8��4�'ƕ��'c�y��T9 :75�����R�\T�۠�t(����S��>�́ �%��J@�$A$�~��ۿ��(9��������:f!�����%��d�~�+�9p����CP(鿕+)Q�sw"j	[%6� 2̱�X m�,�ZM��~��o��I�!ȟ�}�"E���z:�-��fo)V����&b#YqE�D�7�����% AH���YKn�p����2�}��btv1�ǣw�r�H �7qs#���et&�1�O�2�J_d@I6�2 �����v�k={�۾����ɪt�C��A��D�H��I��@��I���r-G\z鍾�$�k���$_{����\,�����3dw�.$��<{�jz��������1}%`$VA�E��ZG~ygx����>����o����pTJ��v���!�d}?fHݳ��|׺�}X�ɫD#�T�������� .E`�܏���ļ��9{����{�/2��=W�mc��ٴWj��B�*�XB݋4���(K���[��p�F]t�P-��4k�j3�`�M���Vd�M�.���L�P�.�妛#/-���-��,ѭcE��ڂ��@r�٭�����,c�X�l���8�a4{K)�+�Vۂi�2�"YaVg)��6\�B\r��0�h�ڗ��i��Q롭.��WYQ�ZF4�<��8�S�P���{��=���&��h��̰��a�,F���Z9����n�,�i��B[��=z��ؐE�����fH��n���{�i߃���pt���`l	�V_���\�A�u���DV�/����W_��QG��݇���+����p�Y�qo�k� �Ă-��32�ww�D�����D��_As��?H�JD_��q�%x�.���ۂ�V>�;�A��B����"�$�Oϵ�?��ȣ*���H�A}�~Ks���ݓN���c� ��N���׾�,�����"�Ib�����z�aZ:�N�ߟ~��q��<qo���	w?[�32���H�WOo�fk�]E{�w�1�R����j�؋�X䂹��G`ђ�s��:�Ub�����?��r�nH��dHs2T'���"w�d�R��o��g�[����`����;� �� fe	̉{�o .:�hE@�U��� ���zqf����D�����e�3�_<��]����SF���=>Ί��]�^����NR�$7��-٘w9hó<8��K�'�;��ݓN���c� �y��yÄ����w�Z:�QR�q��32B9�$� ��lg�j��,K�/��M�x����߬�:D�$_h�d����ܗxB+�8/�I������=��&gx�LJ��H?px���4<��=�UW�DI�%}%"H%u��+3�ڳ�2�O��;)��dӿ%���	����#%"	�-�*KӞ��Y
�*b�i[m���2MZH9K��Vh&e�WZ�C]#3KY	B��nAl	 ���Ȣ̑7ζ�op�M�x��{�v]�(q��C�Hw�� ��=�����_)|A2E�%~�k�SlO�N�J��[�f'x�dEJ��}?;�$�A�������ꐊ� ��r_�@D�"$���˜�z}r9/D�WK}��2W�HQ�0�C�����U޺����J���8�E����"�4	Wu.5q.�7�\u�1�i�(g�<Y󩛾���3�bִZ���S�%���A7�(^HFJ�$V��P�0�j�zP[���(��d����op��7v���{���"yFq�]�!�z3�.���vD�%|�2Ed"�V��+z�׮�O]n�����".V>�qwA��A s#����{�Mc��UN��ɘ&$}��e�ghMF��bT]+0�-��qv �QG�dp��?�<�I��ِ$��cSS�r��C��a/mKΌ�Q� A� �?�_/�qY/��PDr�o�~�nG����({dV�u����n��odp/"A�nD���[�~��
��D�	����dI�3&yl�����y��J~=FS���=� O:���fGِ=����M՝����FT�#����'�w����w�~����A�'�-�7
��V$�=3�2(ҵ]:��]2Z�X�cH��9�~��ˮ��fW���N^�{b�h�^黗*��QV.�S�&�V�À<�A�g�4/���X�d��r�b|��3�wo8�y���3E���/"A�r$�̟�̐��Q;-W�M?�PQ	~����|`hT��t��sX:i�����!P�a�(��GM\*��d�r� �H��dI�d��_�V�I��.E���7���U�k������j}���iD�~�~2R#ބp9��a����C�A}�G���jp��S�a��q�����2"�V���^\
��I����P@�����d���K�Rf�v��~�7I���oy|�$n�32��+�+������I�G4/�|~��IwV�I����S��oH%�	G��@��s� �H����I/��J@��d���̾�CIM_��� P��;8\9ӛ0�����7y(��D��>?fd��U/��Ք�_�S�*׆�}"ʰs��P��w�����}z��Ϋ��v�s2ҭW����p�������ХϳYO�*ŕ{xe�C3G9wUʍ��
����ƺa+u��I���D�j`9�,j;�gp���+6b��X�ɶX��R�0��n��+)-�A�8ۋ6k�	��r��d�٫A	���Zq4m���Bc!sqXuL�:c6]�e��6��i�u�ꖎ�vB���6;uHikK,�4P�,�6!��6pP�!.���̱�����jj�2���x�-��.�rm-څ4c�{�'��ĹK)�#֙-��(�Yr�Й�첍!Z�CA��E햒�p�~�~;P$}�̉�M�X;�q��cÜ-� ^zo;32,��D�G�/��Ȃ2R��+#7ߤ�*�b�@�c���䠻�[�1�-N>�$��v��̎��Û�}���j��	�4l��`��W�P�D���$�7X��:OI�C=o��㮜نn��	n+ ��� �$VP\��d�p��P@�=B�>�� �"v�c+{��n�<9���Ȓnn�ݣ�?Uw���.���#%|��+"#�A��'�$��Aw����Oq,9�8�O~��A G���d�A!߳��~�=�g����]��i���������������j�kjB�����cke|�}z��޽����FfO�fHt���_x�������3@�ݜ����}��"�$_ ~2P@�g��+:���E׈�6JJ��5�)�F��Uo+��o�{U���ܐ��,�k�T���G��y���5���	ze�{޾n�H;�+���+��ķW:��߬�J@���e�;�W}^��3�A�yX@�H�d����m͡隣�~��8�g%��A2��AȐFd	 ��A
���j��ƹ�x�;�ۥ��2D�{��\6}Σ������B�A���oTp�Kk��K�-�XH�_IAd�,!L�\�p@��r����~��Y�g8>���) A|���"��������~�����?�}���]Qn���#Fֻ-��6L=�R7C-t˨�YMq\��m�?�7���쐛�'�ٙ('���<�g%�~���g6�}@�|�
 �ND��Hr�	n�"�~��N��r�����;���s5�%����7y(^H��d(��ro&{�"c����9DvH�~<�	�$�`�H�S;��h����:i{�2E������@���[-�j2efQ����Q�����1�eU����J��MX�X���gNy]��yJv��g��߬%"�_$_X�d����i��鄣��\?o ��PE�߶�c���,SK%����A���������'��;��#��I,X?)dA$� ����dw�"z�� ��s�ϩ�a�8�A��!�	9�􃙒����4���Ϟ�o]r�<a#Rg[ ��֦rʄa��[V�耺��U���޾�A�f�>v�@�D�̑"��[]�~��X���od&���e���B��|��2D�s#�3%QJ�x�gS|=�?@9�+���݃Ñ�����7��A���9�V�pZ�����9�${�I���_~��E���~����O�~յ��:Wz*��͟S��8� ݹD�2R�"�D�*�y��2�_���]�m@d�h/��}#2D�?WFWw\zq�'G8[��}�}^��u^A�{�*x�մkw:�Y_a{�2�,�n��9����x����sr�zg�� >��mZܽ۔y��j�{.֪����9
(b4W�~N�5�笷���0{�ބg{e�{
i�l�h��5�LL�W�Y�tr<<ٜ�|3{���B9�����G:����>y���cbw�H�3�����T��u�ڥWF�p�Sn�%&�F��Y��ƅ�*���-��_�$L�s��}�����}�8�⩚��G}�Ô��s����3%|Fd��P_�t�A1
�X���D�D���ӕ���u����� �D�E��'Tҽ��{���%���$BNdH?fd��VZ0�S���⡏c2�����@!��,)dA|D��s7r�Z��r>��"Aܾ_f@��׸+���?Su�p ��+� I��[=��r�ߢ�D�2PD%���N����Gh��WY=[�q�N�?��߅�%/�!��%��J|>��!
���0=�.r�w����ȸ��9��ʗݨ���]�����e�7]8�g7u_U�v���O��'����MZ�k�X �m��j���n���z�U�h�i��,Z�WZ�I�˲Cl�u�wr욪Ύ��h��Mn�d9�|�<��I�E��t�9����j���5�q��/e���f��v4Yҡs%R3�O�g�(&��t7E_J|ڷ�r��no*!bTF�QL�;E)����k�F�:�L����]�%�'Hq��'#-g!]]��W*���U�f�ݛY����y�,�����R�U�D0D��8VZ�ʛ�Ԩ��Cswn�ecr�!f��w��Ԃ�̙]�w)�ySPc�3t�ZQ��uf�H�M��M�̭��-}y7.��������L�6��+�6EY_Q�MS�� ��MvV�5���Gғ��nu�����W�Z�NL�SSuz�V�Y���,5��}�λjB��,���U:������o�}�ve^B��5y|�o)euA��3�d��;������ķW����qЉvEW�Lb����'L;����',�;���]�{��+��0v��cj�k�-�[��!���NS\�����]��Gi]��emM������	3B!e��]h˗��hQZ��!�S��V+��*{�*��d]�*�]>tn\��X�d&���m�z�)��ɽ�����qimUX����ya�ι�&bH�P��C���i�+����7h^;u�������yY��e�PӶ{mN�Eu�SgWU�옦��kJ,tڤ:<ӯ���;�J~EU`��FSH��)�.8�I�Pr6�s��K���% �D�C�tq��"fD��wfHG �tPM���������r9m�yjvem��98$���=�wfG8��G���H��vpW$ĝN�''�ّN	�A\�\w���kVtrRtf���gpQ^vm�:9���.*B)98���92��(�BNʲ*s���8Gq�A$�q ���II�I��� ��3�&�y�C�r�'��(�����B�.N8����%�'DPB�rĂ�'r3vX��m�:�>}��L�)5�6.��b��iF��[^�w&����a��]���a��0ؑ·\:�-u�f���"�%#�bt;Fmu����
VhR�Z�Z-z����f��h+1--js�V���	pXh�D.�]+����&J��M�uI�N�smCZ�)rQ�L �ո�sl��Y���ј�hu.��@u. �,�55�@Cl�J!fkV��g�mt�h���Z�����q\P�ɬ#�[F��i�i"f�Z:��fn�&��*͸�,����5�P&bgG5,gl�Tн�-5�r����Bk��B���0��+�ѳ,�6�7Vt�X.��K��{�g%/Kdf�gmÚ�[Z��j�cD��Ű�
0�aD.��m�ٙ��湙�#�T��H�K��6@���MkJ�e�L��q2��Nv
&e�5���UYuc�J�&I�bD����I�m���Tv�Pڵ[@� ҅�������b��.�ᘌ	Ukls�
�M�Ʉ SF�2�u����e�;.3���'����Lw��j�ˋ+�F�HW
�]g�]5���1�o-��4Ԛ���m��pG%�olͳ�T�]R2�l�7Ul�f5z��Ѝ(#�ڤv��6ZE;E5���&f4� 5�A����M�@2[����������e��if�GDb��`ò����B�sX�I�)5%�rbl�A&uJ�e3ic��K`,)�M
�jE��i�̨-v*B���f��&�m�e"�4�,��5�=�����-֝��B��{L�J�t�X����CZR�@�7���,�]�VqIH15j�9죶�\Z�M ��B�`�Z�ء.ZCR^G*W2�#�eP�ԙ(��qIl���*����4֔qhME]�t4)�J���.�B��m�\=.9qB��.Ҥ\R�e��lF�H ��ŷ@I��D���6ٱec	j@�bԽ��q� �g����l+5��:��jݗg4W��-��ѹ��4���1462�aJ٩i\���!���R�4J��vf��:�QL
Kd�.�UuK�\�&��ƃYr%�a2[U�(�,G
�˰��q�gf�,Ym�h��z�����Xu�6R.<���B�M��*d�l�U�mMe΄��UR�.�)2��V�r��)�n��cٛ�-�t�2�.���u�G^#bl`��.�l�4c����o��)���������YM`jV5�tn�WB�4�ʦ��qT?�����?�{�>���� �̔?{�m�=Įf�^|3zF{j�yU��`�9Z"D"Ic�9� ��[Q�@�؍�rt"+6~@fH���+���WM�C�q��۔C�s#-h���|�1@.Q��~��$�,+��X��mbSO*�ٖ�o���u�ތ�o{�9� �nD�Ff �2 ���gh�_!({+z���~�A�?̔;�[zN�+�C.+φo	p$�������Vw
>��^H�_�_)_$#��z���AGrw�tB��uƟpj麈{N8~7nP ��$�D�	��;|َ9���"(��`İ��mֶQ���Ia4�3pFR�qiP7Vǳ��o���'�p$�}!nQ7"E��غ��d[�kќ-���D)���>wR�;�k�m/�rn'��nP!{��c3���ײSȥ�8����O�у��։x}j����y]��}E4��X���+����Q[q}�|E���H��2�v�2�+�8��?k�]�'xΡ���ټ?p$~y����z�P�-�;�$��	�r�7"~6��܈��	ȥՇ��Ψ�E���!�8��۔A��E��A-�_�AVo�g
>�:�l���j�(�܉����]{\�V9�g{�}z��]�`S�SBA�?.�A|[�?6�Cm|�O-��]A��lh.�S�S�K�W:r_��ྷA6B/��nDk9���V�E�|������h���*�7ML��M%]Uf��ىW;L��U��$�^�]-|���|�ƞ��Cn~M�'f�mC��e��s��#��xk���Y3E�I��ۑ`� G=�4��ܛc@>�?&�\>�w]�.�[���o{���� ���^~{BdY��]WK߽����$N�� ��@�H-����q���F�F�R�U��'�.�E��Ԛ��J���,�ޝv�ek������p\	v��u��w�P�����8Tu|�r��h�����LY�*��������:�w�|?n ����(��$6�[c3���esƥ�Gt�v��ۑaj�{P�uwm�s��
�?]f������q�AΉ �������A��+q�����F�R'���]�pn�85�1�5�(��Cm/�ʹ��S����u�e����#�*:��h�*EY�+n��pV����\=n�:�[,6�����?>����Kq$[r��=��tw~N�:|3}� ��{�6�_l�j�C퐋�? ܀ۥ�n~�ҹ�{�G;*~B�PK���sì�v�Þ�&�e[h [����q�g�%=��_v��m[s�ȕ�����J;�+���ӃO�=�ƳeFl�!��Ŷ�-�՗g+���/'��z�n(~-�[�z7ǹ��:.m�ͮ_<���K���
�}��,�z0P;Nm����\���.�6��T����V�.Ї/��f���њxNVU��r�#�<$Z��u��r�?~V>�?�@ Am�܀�k�5Y��:���e�t��)ܼa�S� �r�~A��n(-���l�PI<�|	�������D�9	q6�6��ѲŻ�B��C4�l�17����H=��m͐Cr'�՝�{9��?8.�c����og����J|A�D�-��-��q�ܠD*^���S�>]�{��=�WNVލ�ͥ�m�ͮ�^@�A��p�״Ϻ�E���i�����nD��A|[h��6=;/�7�W��ƋQM�z�p �]�m��n$Am�6�C`J�4�>� �x��� ��M��}�{7��?8.�c��}�(�t���]�1`���-Đ~-�_ې�-����{���D�����+���qs�`soFmw������+�rh���+\gYѿ�֭%Y��g�#�)�`��4o*�:�"�<W�܏�uLsl?:���p�3v{9�X�֜���+�A��,�+�B�K���X��uL0L���pؓe֓E�D�0�U��4"�QW���%*ҙ�]IFb�Z��q
�Eݣf�n�c��^�:R:���D�.�Q��5�l�[���f[�Q�KYe�4�x����ற��;��R��FaR 0vD6Ir��\ay2�K,e��8!�[)�jgC�˩�u�aBl[�sQ�Xc���z����<��	��TLmC��G�5�VQY�\�h3B�7a,�Q �H�8F_;nQ��Cm/�m�=/ٴ�qM�\�dp"��ñc^E΂��n$�۔m�-��-�T���1���A�M�����o�~M��=��+e�$��Dgq��3K��~�:���� w�ۑe�D{�;����e�Y�����ϩ��N���R;����A۟��D6�C�e��o{}�~�M�b�/�H!�����m�Y��Ǆ�Km�=yA���@�j.�]n��������۵�p$��A|[s�Y§c�͍�[��/��7�ۈ���'ײ�/dI������U�~z�����}��g��;��(�R�(��eIP�f�Ε�jX�R���m�Z8�.C��~?���C���E��͹����q����sN^��pB��{Z�W�%o ���D�� ������xKN�{Z�[�O&Gfm�فgJ�K��f-��/�Tt�P?Mא;ǈg;[�Yd�{���q�ءu3�|hĿ�ʠQ7������4��5�{��E�n�\}�{+�1��coŴg�h=nW�nb�t	!�! [r� �#&T_n<�^��󎛼���7��'�Epǽ��l�C�Cm�nB �EscK��7i���Aq�[r���:�f{�4����v�I0^S�'���*� ^\��?=�$6�_6� Cp'�j�D�GP�Ͻ�<A:����
�]��e�@/6Qm|�Q��$vf��v�D�8�>�B`Ȁ�=��,�R�b�s%z�+R^iMZ2�CQ&vI�p]M}�H?|�����	־�7�|��x�W�����>�QQ�0�w4Ar$��_�h"�I�۔F�G��͕=�c�Ή ��w��:�^{�^r�k���Ff��-��a;ߪN�z�c~�H�Gv��?|s��
!�������<��-�ň�L�4�~>��W��������rV7��QJ�Ε]�Aә<|r��uJ=��D�r<���Y���}��k�����p���'>����y��q����F7!|[�?6�k�._��]>����@�#O7?7����q���_��"�c���_Vr���OP�R�w�k��?fj�A�۔?6�_�g��kO�:L(Z$ۜ�U��é�箫�=�� N�	����"۔AnE�uUk�����a%D���3B�Z�e�&ARj*�W�5��F#��flR�h� ���3`�/�m�O5�uϼ�m��Q��Y��{�B��Fm������?�t} ���H[�,T��G>T�Y����t����q��������� �l��ȐCl���#>���8��J!�!�~ �ܿw��ϟ�U#���������4�k�|�;p�jܢ� �܍��31�� �H�/�m�����}�s�!B�6y�q����}���Jz���F���zx�3a�pt��~�DЎ9�Th� n��Y�(� �]%;2�ח�`�u]��{���w�;_���3/Bff��, ���̷���Q���Y�%Z��뎛����<1�|���9@����A|[hS����6'zeJ�
eL�0�S	rmVaW�M5�Ҏk�U�Ś9���:R����������O����u��Oy�箫��k���(������ ��A�����I�͹@�*�9B�~������|C�AN�7���}�D���?G8�Qch/�qb�
��� �T��l A� ��Aܢr#�Ў���e^f�Úmϕ6�odp5NW��n��6�E��+tF:��꽕67�����[r��w��Q�8���z[�w��~#��M��u���>}"A�%�(�܉���TfD>�>����
|���_��Ļ��j� �=����@�A�>��ڣ��>��mҾ����HR�y���}U��j��Jŗ���Y4P��㠋����U����;�x{������o�9]Wv�3}��!<�~�۪˸f��¬[X�Bm�:�eʭ3�w15B�"D.�lƍ�����V--ZW`��њZ�0�]e�����#-e*�a79-�Vݭ� ��L��29u�� X�9 H�V�e��M5*��q��P�!.�õ�!G��bK��z���3��v�4�[2QҖ�g�bnE���,v7�l�Gy�P-���k*%"h���>[�x ̆
�Z�`!��*g\��f�^�f�]�)��!3�@�S��@��$٨ [r��K���ꍚ�ʛ&xc����+	��F׻���uH���������m���~�;}{���u�7P;�Wٮ�1��97�����|�܁?s5ns8վ��{ֺ��|���7��Cm��2;j�r�Vg�g+������8���f5�q�۟�v�
~S{�l� �٨"��Cr$<�>Ψ�-�Sd�{��w({�`�zy����x�ݛ!�I��m��q�Lv�b�+�s6��yr��Į��Ѳ�w�r�s��?[r�}��]Ӷ�����2I!爩Q�lb�YF�TR�F�ʺ�,F��g���пs��L�DG.�2K�{�����8;�ޖ=*����25K ���@�D�A-�D6� [��V#(�����{j���%�)�<$�秭/^�u�MQ#'+�7,�����m�*�ݙ$�����eSɽ�3s�5E���س��=�FW��d��!��>���-�SN�ݑ�������^�iW�������3�'_Oɶ�-���m�L�MnTUF���Sӑx���|5�@��~��@����Q����>[��22~�����!���es���X�C�}��j� �o�P#3=�d������H&۔Cm An mȢۘv���<�of�u�r��p����Ӕ!�!��_6�'���!�b�˨b*����|���%A�u�����
]3��n�u(&�3�ɄL2���a�S�� �-ĀA-�W��/�zn/%]7�Z��T�xo��/�����=�Ȏe�&fh���Duo���٘A��u�.��ޠ��\�;s���=�ٌv��A7�+�r-�vq���K#� �:�ʹŷ(��x}U�fFĘ���4�W]&��ը��&���	ٯ����9�n�K���E��U]���֟u�i�;�.�D5��u�n;dT�㚟$CB�GZ��qk���t�՛Σn;��Tztn๗�񫴡5H�p~k��*���na�b����Ѳ�m��:XL`�g����ƚ7X��'�O�]�D��4k�'Pv���wu�L�q�d�nZ��$�b��9iMN�W�и-m�	�Q����R5uvv� �t��5�J�Eo�i��I��L����l6�Q�����-c�6�k�MX幙���J�Mer��9�V[��۵�=ֻD]�U�e��U�.M#q�e�tx^�*���71��T����~�q��w����D��ϩT���$=s�����S�$K�s����.�'�>�Wc]T�&���}l�����˳��|
D�y�����d�}k���4dCz޴G&��a��e���q�L�)\bX���v˜p����C����'�Ҹ�f�rkz���:M��T�x90���r ��,n]?�̒(�]�h�z3������L��Ql�)^R��6kKa��W��M�u{�fT%n=�]N��[ӭ�Tx�Ƿһ�n�݃��]�*�[X�mу{q�����ӄWM��͖b�ʨ[}�
\���i'G+޷�j��I���싪n�*�c�-w��Fe��*�H��j���8����5ex�Ui<��IÒ�mf�4u�*�fZ��8+=B��JX�
�2��t>���4�G�m]��}�V�Wn�)���Y��>%� ���	$9Y�*C���+�ޝ�)�\8W�tB9ӑ�=�N:Y���;��.::8@��B�#��E3m۸���#���; �^զ�9*NB̦��tTGJE��ǵ�$���q�q��N8�)'K�����ggq(9���� �$��6�H"/k��	P����9�<�p�D�A;��'����t�8η��\����mv��E��9�ptP�w�aA$q9�Jyd�;7�i��aru�R8I�8�$3��{Zp��e�DBGrum�N:Ic�IDADAb����w�r�i�~~�bxf� MӔ!� ����A�H"�_���]�y>��7uwbH%�*�w/�zn/%zǛ�w���GO�f��mz*�9�+���_ Am�!������YPȗ�s��Y����/*��j� ��CnB-ĐKneg�Z����B`�hI��61uu���my��s���Xswn��d%[�>�{��	c��۟�Ȝk_g\V�i���᛼*��Cs'n��J���͂�@��|[h/�q �r����y��i�tH?_t��ܼ{�鸼��G���	y~ ����m�r�xa���s*�
��<�~n�K��C\�z�=��zh�b�vk����.k1�� ��@��q ��m�͹{[���?t��}z��!�-��κ��^~ʸbx7�&��۵b��c��;��}U{Y]���ox#������%#]�7Qއq=��d �=#�9��Y�v���ɹVҝ�8��n�3<o=UY�uÈ�d��u�-��A���|!��n=�F���Т�Ϻzu�y��S�w0�����?�'�ٍm��z�':�o"�X�T#J-���Aв��E�[�+��p淶ݥ���M
Q�JILmU���A�6D�i|~m��,�޽��P���;T}��=��B`ى��K �j�%�?6���{06޳�x��A�9��&�����u沍�<�_c��>� ���zy)Ϙ���tP �����mq$[r팬�1S��OM�ÿTS|6rG ^@�cA۟��D6�����خ�Ҳ|Aˑ$>�����P�no^��Ϫ��c�>�o:Q��7�=���� ���35[� �h [s�\$�����ڑ?�ݙ޹�꬜�lO��@�w(����_�m�σ�$]u1��⫇3�E�\*�:��<m�6�Jޣ����SF��*�r�T���J��[��u��w\�m2&����8UIV�um	���U�!�!6,�s��^�0��-3eL�*kj�/%Ќ�����<��k���1�މb�1Si`��<ِ�jقec"��1�A4�m3],�*<j�umDj8���������UL�Z6���Ѹ�R0�ɗ]5�,���V�\ښ$�kte�&l)�*�6�M��)Xi�\Q�$T��&s�����n]4*ɣ-��4f�t;8�+U91�~��'����m�6z����[{i�\�euu!�W$"L#wq�Q[��q@�[sx����髗�oF��*��$O�9�|�V�=�(��r$�H�nQ
mF?f����#7'�E�K/��s�1uqK1��p5�(Ƃ ���/	!�X�gT��v#� Hm��s��"k˙���;p����c��Y��og�ʞ �H�m���n$�Z]L�o���ȿ��}%�(^>�Ǵ��l��E7�gx Á �U�u���ϡqZ0�(��$�A|۔A����	�>j#��W��>��3/{��;�W��Q����@�m��-��?��Fw����NULM�F�ԉ������L[�n`��d�a��sj�+�Q3�0�m�?������4�#�W͹�AnDŽ睹7�^�Y��׼��&����ὑ���z�H#^��6�E��A����b���Y�T����Y^c�h����#Wl����!����9|C.��QC�	Ma!�$�.wK+����tg9P��Q�W��u�j�8ۉ��{:U��x��{�����F�|�7�$���E�'z��޿Y8#��$�ꐁ����Cn~_ch*��}]B9�z�k�fw�e\V{��}��t�Ax�E��-�D6�3��_�TB�_n��Cp'�yݸ�1g{ً"؞��?w+�7H�s�>^����r��A���| 6�E����1e�gtIY��z���Q�����U7�g{���A�k����܌鷢gY��K�H�U�|�Z38�7nc�)��g����]e�v0��RkV�5�+G��l�?w/Q�Yi��_6� !*�����ɫ��c��!>�rNin����~m�!���������*�(8lQ�ܹD��/5���\Ҽ�E�:5� N;� >�$6�.�'����;~���ǜH �sv����C�W�f]�aZ���ۭQ�Jj悌^�b���C��H7T�}.C���� �N^��5��MR����v�y�־�����=�X�fT��2�_4��B���l� ~9�$~�h [r� ��I��Z�c��3������6�P�gong{*��Ōv�>�Y��"��Da�S��Q��?n�@�A�n ��h"ۙ�:^)cϢ�`�W�r���9W�Ql-�� �__H���#_i��97��L�3���zW�&�u J3q.m�5��iP.��R�J�XĦUs��0A�\�?oj�H ��[�7v-{;B���l�*n�����Y {��ײ�-��[r�Sl]����ь����_m
���s:���Vbc�����~_<h"�{<�j���ln�W�vr@�t	�h [r���K]x�+Q�������r�2��\5���@m������}N�.��ٰ۪��Ef��͉��[r�߷7v-Vv�sM���́$O��I�8��{�o�j�������6����&L��T��w{Ÿ�@~R�(��Z�u1	:��,�F��_D�])�k�o�Ĥ�p�%� 6�nW�܀����<�����@B~�ǹ�N�Z��G��� ��s�m���[s��
C����Њ�"��Zn�&��`[��#�Vm�#�W%-��F�g���&����� Aہ?��-�_�	��O����^T��x=>�h�Q^�je�A�'�76~M�-Ă	m� �SY��ɞ��w��'7g[{�-Vv�sM��\'2�ٍnk)��䣧�_�D��@�ޟ�nD�h/�r#��A��{v�e�wj�^:;�?c������͹D6��6�3����v�*�B��9_[�0�����¬ʋc�5��~��E}�:]r��pP"������"�} ����_7	�ޏ=SQ��+���fwlM����M��\�.�Fc��-�D7!��*�:f�nla��_�]o:?��`������ܩ3f�gaa��/��ꇼG�P[�u���<�WΥ�hg>�qD��V,�w��O������\���#,��x��^�-��m-e����AKv���B)��&��<�p��;��^{+ĺ�C6h�ը6�
�a%�v�lFY� QI6[��^6�I�m���6��q���EHc(�R&�h��r3Z�2i���	F��uZ֫��mM-dk���͊�n��k[��kR\��t�v	�̭�k�"�k+e��%]]�)�����c	��X&i!�(4��WK�f�%M	�Ц�����M���4�C��!��$�m�m���^o�r��Z���G���98��d�k����G�$ s��-���?7�ϯ�F��;>���Ș��}�~�q^̨�+�n�@��r� ��$�����x�G\��%�J ��m��-Ă	m�\¨�~��f#N�W��]{;G��|��^4m� �"Hm��ܿ��ٛ^s�^H]|����k��nW_����t{j8���d�c�j}�tl͈��G���oJ ��@��I���1K�o_����"D^:�ڿw8����+���	�9__H�k�����`��mT�$�O�6�E�v��6�p9��&1��\�Y�3b�fh��76j�ۻs�������}�Q̩`�r�Oswb�+�������+����]�kN� �~���_[�r+�۔G�1ֻ�J,U(r�c�p�ߡ�=�nX}O'W��W�0y�3�J�<����I.vhJu�y��7QƷ>��8���2��EU���+���m�_����b�j>�V�����CdX��ǺF>����':�r-�@��W9��@�~��˩�3F������`W������Ÿ��cro�}>܌�����Gv$Knq���ث���\��up�|��S�Y��>����f��r$�H�nQ���w�4:\�d�}Q�iz�_]u�����+���V�@�n~n(�ۛ�W�c���m�@��o]h� �LE���ʘ]�!c�٦t�C5�eog䉉����>��vj���	��{v������m��d?LU�랺�}2��K �t�!�/�Ŷ���	m�!f�E{R�c��� ��r��6*��W-��\�.�O��4�����rr8��F��"H���;�(�	�����m�E�b�@�qq�>�WS�o��Q��R��5v>Wt���X�.x`�?Y��;�i�i�P�;
�l��Z���t�[�յ�l�5>׼�0w2�-ۻ���=�����r�A�H%�(��E�dȨ<*}��Ԃ=�~A�gv�]�y�˥lg{�r��EV����{��ګ�����s�n$�[r�-�-�x�t���ٝmo��5sO�:j�o]���n��]��A��AnQ7"�V�S�SؗM�����g���XF;`�e1����k��3ePv�G7�h��������}����i�m��m�JS��lg���~�"!ة5�v�f�]��8�~m�!��@��	w�y��?_�_�tw��ҁ:As�������]+c4no	�9��m���=�Y����~��� �q��m��q����gm��+^����W�X"�E����/ H �h [r� �"@!���4�DJ���z:h��D�Gg �!������{o�[�a���� �r�c�f9��Һ�z�)+��O<3!�F)�#ѵ_��V]��ޱ�궫IQ_���z�bW�S�^�盷�� �f��G A/�P!��� Kmnv�>"7'�t��Z�����ں���77�'����D�h/�m�a�E���/��1����毄r;�WB�0P+.΍Xb0ņUeܸ������嗥��㥗������(�m�����^�^uX������yk�����{G5��O�6� nQ�ޅ�މ�����ݝ"��v��R�2���8AZ��~n=GV�p��UeE����������$�m�m� �܇��{�캚��nW�W����[�s{��9_@{"A��?6���}�[��_�]O�����A���	m�����+3��]��|7W/ O�xg�}9������K �ȟ�m�@��nD��c��٘��us�Ed����߽�`{��ex�}�. ����{�� �@�I�@���D� BI���	%HB$��B!$�2�	'�!O�!��B!$��@���2�	'���I<B!$�@���B!$��	'���I?Ą BI�d!O�!�Y@����	'��PVI��j`�6l�` ���������        (@    �           
 �      ��  [��
P ��B�P@P �J�
�D�P �QD� ��P���@ �o��Q�EPR*���P��@�
�R��!*Q)Q
����R%P����J�UAD��  I"ITER�H 	� �} 3�:�7`�� ¢, ;1���\��; �ԈL à 0  x  p=� >�� :�U�GT ݀�<�t PTD�0 (���F � ]�zj
 Qy���)�n��ye]�t
<dD�P� ��"$U!RB�"��EB��)�K�@W�Þ*� �إ%� ���ڢRR�;�	�*�nn� ,��J
 K� ;�����h��P�\ ���9� �d ˹@+ $: ݁�2Tnà�)$�T� q�IE@P��$JE*)PW 2x�n���� N�, ;1�݁��@#݀��U� ��Ӟ��UQUJ)=� <� E���t�J�@� � � �;� q�H�p ��9 1z@���8� �(
I)�  �R��A��(�	H���>��@�`��@ O�� c� ��� � V"� �����(�/|   �{� >Gv }=\��J�ٌ@�p ��� j�*�V ���v�z��� �(H 	�   ��>	RT�J�P��	< ���u@݀E���^x�C �� �@s�:$<� #ΨB�#�;�
U(�P�   ��� z� 3��� �� ]��� 4X 6àu������=_CS�A���OS@ S�a%)P   �Ѫ�%*h  M����R� �$�J�=L0�	����Q�5*�� h�������?�G���{���xX���V�{�̱��BB�R����	M�BC��[Z�����ն��[Z��j�{��������_W�����J�9�*5;�̸,d��]/���W�R*Ɩ�@��ټ�XJdT����Wk�̵J��Z������Oa흣 �SX�&'��-=���7l#F��$��:�!^[�WEԷn6�;����T��'	���w������;s��`Q����Z�9�n"����^@s�jќ�?�D���˜x�8;���NJ�u�.=������M��w�X'~��	˺�ᚪ�8��U�ٻ��z�T6���#��l�6�ϻ�P��f�g9��ݺ��L���;U�����LJ,
�������	b��gƲ9�
��[�w�m�Z�OO�4m.��n��T�@TD|0uҵ�7@ZVh�!11wqGR��=Ѻ�v'�\���^���e� Eos!����fY�,�Uݏ{	�U�^�9=�k���cK3�#�5C�"�"b�SN\��JTSńGP���M�霯\`�CN���bdrͫ��Za�ö��}��Ӡr�vk��1��C�d�z.W�L%�cHq]�Hg���B��q<�����R�t{\`���`g8�R�ֹ�/6��I����7{s����\� �k�T�L���ʫ��ِ��p���.�M�U+we �7Ë���z�f�BYx3��*�<O��X�i]4�fuPG�1�r��l�q��on�}q�ّ�MM���ӵ�s�D5��v���� I�n��.��}t�y���u���$\��.��)�і²&5�XT��<��q��l��v�p�ɷ����{����r���]�j.���t�ե�3m�>�����0���6gD��wY"�5gݶ��Y4h�Wq�w �X��c�فv��ϟ`cx⻰n(Y#��Kv�W�l8Fs�s�v�,��7����r:J�[�Zw�]����+�c�������`pw���V�Ln�!.�3�,�ށ��F�>��P	�^t���3�mz-�ΰ��&�t�FG�J'���7wP}��j� ×����&�Fj��s���I{X���z�h�=[��As�a�ԥ<�F�Y��GwD�9u�u��2m�V�S�$^���eJ
b�'ght�0>8�Ir-�-H���us妣1�������Mł��5.�N�+�����w7�G<c��u<�8��+��:�ý��HrUf����}�)m�I|�cm��g4��zqs�M��w��@�N��H/慽�l�n*tτ2'��n���`\�V��r5��0UqWa�l,�r
9wO!ٶXؘ�wdYe���5.v�FR: ���u�"1MHon��L[V6�\zsN��-���7��\�]U`�HNbs�ۛ�B�oTTmn`_�b�^S��!�u�y��7-"�>1�+�Z�e�͢]�yt�oeL숆j������06�p';&�`H���S�m��Vhc�UoL��'6��sM�V�~q�DV#Dn;eᜯ,K��$@�����ǆnm{�K����vc�f�{y[3V���T�9	�
9"��)m����H�	���ݏL;��c�r/[-gb�������6o��+%=K;�~�U�b!���e�Yaʶ	6�"}�9v^��b�]�:��p�hо࣫�.�T�0��g8�xA7o��X-o*/>w+g���l�@m�.�e����t�y�����Խ���'��A�킧�G�SS�܃��Ր�c%'i#��3�"N�g*�d��};:�&Ǉ��f��v�吅�ݺ�wi���,f1�����%���=��.8�m|^
h2�edp"�{��&��M���:��2�hX-C�ӣq-/,U��l܄`�U�z��%�{E�tD���Q��m��*5�R{������%�u�u
|$e�6�߬� (��y�9�;��j��o.��m0��1"ni5����K��+N�c�>�MΠ��R��myħ��.�K�����T���E˅��8�x��v�^��w(��,CW0� zVjq8LT� �6K�[f���b)��8c�Y6�d�;�}���oC�.��(׽��._����k}uH`�{�ۃqtm혻��BsY��ܛ"P��-����=��j�S1KϳA�"^G��Q�t�2��K�"XfG:�/U�p�x	|��͎�y��J�;�z8�q��Pl	�ܜ�P!���c;l圲K6t�!r%�B֮�2\kS��k���iw��J�s���v�r�ؼp<K�tѶ����3z	1ͳ��Z�z,��i���>�5ms�;��3L�U�W+��e�W��H�5K������҂����}�T����8xb�r�.�ԼO��� }�h.���_o1�q"�@����)ۥ�k�k?n���Jͽ(�e7�r�+��Bj�a�w-�˃���ۼc�.����};(v��,��\���ƈ9Ӝ�C��� �Z�n�
�K��&�ĵ�}��â��@1꛶��9al��E�:N��^[�g����8�!J�q�߁�*�q��G&��`�wF�uV*^�ű�r뱽��7�t��k}���v/�:kn�/:Y�:RBv��>N�F�Y�l�����{X�rO]�-@�C����]0+�˛Ӵ$�nYrFʋ7s��,mb��v������;Y��(��974��1+����zvsT����R�#w�K����h�.G�tK@��b�-�G%���KJ�cvҴZr2`�ii=];{"�;�eR���5,�����H�M��9r�`����֍8u	�9a�J�+$,�N>��ۛf!N��7{6��e��R�>g��i���w4�Zá"�=Fl+]��������r���"n���W�en�]�u�����Q(�ݍ�.Ű�8h�B�d��US1����Z�����SK�[ɽ����3
'^�-D�	�R� ʻr�l�� /�F�� ���I���X �ޗ��b5����	�&����õ��4|*��%�,c��'8s�7U�s�q��fF��C/MÏf&R��s�6�}���_<��N���7\��l�(,�P����~:��LZ�'1١Y{���9�ӝ7�v���}���w.��:��%���弉�h뻧d�ٶ��
�%��һAL�i�(04�fB.�;�`�w`��폣�y%�qC������p�j-��@5͘2a�o`د>�|�=�{��.�w3�D=�7讎\�S�$i\�Q�zu��*u�dX��p����אf�*L�f=�{�N������#{sDF��� �mH鈣:�Mߍ�A0��ɜ�-�qp"��m͜����hڹ^�&�:��ȌxF��~���5\K�7za�k���x��ݎ�:�;�#6�3'$Y�l�ȀjsΕ;�	B8��5��6W���L]�72�B���:�>�~���#���(곇n
���7�����9��k�=�T'��5�E��K+B��g<.<y��y����Ɉ�b�F��-4G���j>�덛�5�95�C�����q,��K�����bO���u��ܕᐝ�����9�|�N[�f��/	S��j�:Mzw�.�k��@���jv�e�9'-ͯnn���.����֭+���Z�����o�gP_r]���C�Ʉ	Y����<�>�黇������yD7E���϶d��nw�AfD���'�gxn2A?Ve�.��3�nn�i�����g�g�bt��GL޷y.�N�׵�D��]�Y:ة���g9���2��ù�d߂a����g�=*�{.��ö/�lk%Ka�Nr법4��6nqӃz��.)�0���7����� �KZ�e� WnD�7��8��ob��ݼ_�5 �"��^����TL��S�9��)܊M��-:�-Xu���)c-�G���m�yq�?����"�g';�b���u�j�<ݺ�n�rk�J��$J���IX�0d�\�yQ�E�H]���quy�P��Xi��������m�n������<���� �٭s�
1ݫ�e=�wOi���;�BHj̕���ǹ��·��k9l&=��&]"Gf�y���w�;����Nb%q��q<�Y�w�`�;��ʌ�:�:V��BXX9k�w��� ���L�Y���F��c�:�_^͡+�I���}hX%��NX�M-�պ�B�Rk�WuLM�U�6\`��e"�&g#';܏�_��t^�8ށO;�F�o/�*.�۲�˽7u8(;,9Gnoۡۚ�*0<��&]����pX:�-B��w�j op��b�/�ѷ~���;��p��V��]�&&��*�!w`۝^���2�'�����o_�|�7؍��GU�Gqj��A��8! s^���马�oo}v��:�n�X���Q�`��>������.���w9u�m�A�\�{a˯���!k��t��F��uv��kC'3��q�ō׷��P��[�ӻ�����FIb�5�ٹm�x��{|�[�μG:��O���NI�m���T���^�]Y/x5�d��gf�&����g
�o�]E����3cK'���0�9ӝ���:�^���@�.�B$����W�wW���5�qq�/�4�+t�����`v{j�yvy\o�M�G&Ls8OUV*[{�v����RD`�j����r�Y��q��'n��+��w��!ޅ�u�{���*5q8�s3`؛Y�5^�2��͍'�vor����v8lQ�K��r=���:x?C���%�H��'rW�`�*��W+�{�o+�2F��~�؎��z�'iy�%E}�������v�mor,����ƞIr��;OJ9��34��+���ۃVj�F�عoo�������'!�6�k�q�붝�nY��>JL������q�ɫL��Q���鯫��8rnO�be�d�PQ�f���8�_�cb�Wۍn��t,�����s��I�X�V"ܽ�bIl's�R�s�w,pۤ�9-�u��Ǣ���.e�G�TGhI�P��U�(�{�k���p�JwnS9UA�n�K{KZw�k����ݺ��"0���"�c����®�0k3N�1�ԍ�]Ɖ#X	���P2,�|�����΍�F��a��moj�k��/e9� "\������n`��t��U(�kB^΋'��ӳ@�2a��@Nv�Ðf�o�. ��j7����K����ݤ�r�;/4�����p�5g&��ю�y�Ҝ{�S�U5ɻ�U��"zoό���?*x���=��E��&.k�u!���$6��ݿd�58�j�kiE�����H2��ը� 7a�ø�����^.�Kb0�E<k�.f\C�
C�6����F:��r:�3��qU�I�Q:N�����hv�	�._�_U��e8b�N0���vW��bf�J��`ͅ�{�d�t�#�<�^�y���F9�Q����5�Iq������ݛ[ȵ��������y��5Ht$B�n���hq�����R���|N�t�a6�Ǻ�Un���Sx�c��������ޣ ᶝۑ��+�f���!c\�խj\|;!.m�D���'�7F���3��s��ۢ��PT�YuN{:ݘ��y���Tq��M)���2v�s���f�۳q�楗���g�0j�ĢĶ3� �I������I�9d���"�[��^�擓�Q��bc�[UU���R���ף��;w�Yc�,���rq�\��Gmq�œ�s�`�.�LՒ�ݗ���Q/نn#�FLZ�5����{�E�әS|�i�aHwo=$T�RR���+qk�=W�Zg;룉o�^�����7��7��d�4�ү��S����6-I���;�j���k^ķ���[�n"������	�6_G,q��z�2GXC��?(�j�
��lF[��hM��a�&La�(h|��׎�`L��q�`��;�ǚfI�lMם���7w{�1u@C�N�%���K���>*ּHX�";ukZ�O��Ï�&�;`a7Íyҕ��nv3��;�W3���L{̑N@5:�Q�m��o+���Ypb�Y����K�aN	W��2N�s��QjXx~���Ӝ���LYK7m�0�oi=�����=Յ�cu�]���K�e����	��Kܼv��s�'H���j:��.����	ڇ�����y<��;g<��OW荾�x�t��u��J[Hx�ۏ
a�#����0׷�2U������gs'�{�{����L�.�����x6�����4طkT�S�ogu�����C�{Q��z���7�ݎ��:�I����B�՝�����(�a�t��a�0=�]����#�y���r��v����R3s笭LR@���:�S�.H�3�Ӭ�oX��vwv�	�;�\#��h��az0����R����#��,h�5�[��锁�ft��QA�^7"҆�]7w8�ٓ�v�t��ē Jsfp�;��m8�'/#�*2�e��P�ի2��3��=��d�d XI$+b��U�5F�Q�����6�حF�ڱ�E�mUF�*��X�ڍ�U�V�cU���EX�bլm�Ѷ�-�*�-[h�cU�Z-�Q���ڊ�h����-��m�m����E[l[hֶ��[�5V#hڵV�b�m�5��[lUmb�b�*�Z��ѵTm�Ŷ�Tk[EmT�XիF�-�k�+klcm�U���j�-j*�+Q�X�TU��j�[Fբ�j����[m�����6��X�صUF��mQQ�U����kZ-�E��!!!�HH@�fv�s'������D�W�{�,f�Wo2�Vnv�]����<�$My�n����k�e�0/]�)��p�c
���f�q�u�v ܥ9���jJ��XF�1���������8Vu[OU��j#�Jr�;�%����|���rW�75gf����#�#e8w]�r8�b5��]8t�Xb��x��:5��:�6�n��4j�6Nn�z��(`c�u�
<K	#�x���Z~�=�!��p|e,�R���J��?o���=���ʴ������^�0����ܞ�n��8�(S���sǼ���Rx�+zeU���Jl\��m���w��^�f�h8��l�Dx�_%����>=�+b;^Ɨ�<��v#���1_��&_'�NH��~���1mQa������n�F���|_�um��KˊW�����Aѽi���xu�Mè{Ǣ�O=<<��m�|r?>����9�i`I3�я����)���ǆɉ�'�o\�`#��vj��x-"�t`�����]�p�E��<"�'�h�wnno/,9ӵ�����{_l�˨4:�6^��F����!x&ڽ���ۏ4�oV�^ɩ�q#ݐ�����}��{Wnݺo "l�?>+9�]���GN�٭���5䙓H�YulNZ7uR>���J�>�y�9xď{���s�Tga|o�X�Vφ��	��53����$P~���r�b� �Wۈ8���Y}q%Rz�/yM� ��K/,�&#�+/���ÝkU�g�Ad�=��`|kl}ћ=��ڐ1.;��~��	.��f����;��,Ap6ji�/�-(�.PA5���S��v����s}b�V�\k�{)j`Ǆ�]g��[�>�?bZV����ɡs�3�Ơ<��ēyk^{��~�6&�ݗU��X%�qa�!	��gsnz�;���;D��'^��'��JX��PҞ���f��Q[�:��kptOW#�v�݆]��u|[�>��]�/y`�ǭ�ν+7����q�k�q�u���;8�o{�w�팘�ݓcD<!KR�QM<a�a�FZ��i(̛{Jq<zK���^�Im�D�a�&;�⦜�R��ޜA.� Qͣ��2��g���c�ѯ}�w�`��=�]����\��
����6�P��g�4����pV����L:�h�Pv�vbb�9kqJ�;"\��������{��Њ�o=���m�ROhWz��pֵ��r���hzŲ�^ğ,��D�d�3N�L}�1�4�i8�b^؝��t��8�N�����+���vYU���1P�JȆR3���#>�s_f���<^�y�p�qdw���Ú�T��ځ1h��c& ���T8B��������MP�\�q!6�1��\�W��xK�+Iپ�ڻ�H�y�E�{�,�Y�8���=�\z�5�P����}�13n_?�x]�o��sq���{�|c9����f���p��C�8�n.!5�B�Y�8�_��W���l�zq|[�&��l��|�����s5�4Xk�����ǵ�c}�z*�x+��g�������n��M�X!i�a���r�0�>�m3&:�Yǆ{�.��&-C�H�P�
���	�AyuR��Y.��O҇Xi��ۖ=w��{�q?5�ʖ�,ŵ,;;�S��J=���Y��5<�x��<@5��HZ�����rm� ճ�&%X���nv+�)���	�N>�r�e%�1I�8��4{��J}8lg)�n�^�b�{N�ݕ�<��k	��L{����(M�	@*u��l�[�U�7��҆3<�b.�������yq��!�Xi;�`�:��Ǜ�oYz�ܫuM�Ƽ���Ypt��j���UWT!{�ݏl���Ԉ�c�x�YDg��#.��CV�!2����k���O���e@M�{�Q��1�Ğ�n����ǽ�J�>~��[_�����1^��h{��&D@��c��q���r��G�x��/k]����74x4�ʲ�B.\Mfb�{�#D{6L�Zrj�>U�b;�b�2�۶��{n���X�z�Wx��+���ӂ�G���	ޑ��M��F��Lن������6�ڸ��G�;r�ձ��G�+� .�gL��<C�a�$c���������xg�5r�C�,�Ay�P��Wd@�޶v}ښ�><
���+�'���������Q�Ѳ>5���,��L-��Eѯ��I�bazQ؉�D/n���ɂa��ݯ
���7�~��^�f�|lfN6\�.�ޒ�eOi�%�5����1�l�/^�ǝ�:�u����й�x��9ձ��l�$3Dk�Bh�>׺��#R>��=0�s��yy骸61�t]�w�{�T�<��}�+)1!*��<����?k3A�v�RN>��bz�h\�E���N�U�)E�6�zuR{�cɴ��8�o��=���dR�-�f��n����JY��J1@Q�E�}�o����:;���$�8�^ʊ9|w�İ��'&��P˹0��J�$��\@���hc+��!@L�oY�x��2�xɵ�@��)�h�Y}�}鱿z]{���: �n�� �13��Y���s��Ư�^JC�+m�G��	O]�Τ�]m�y9�60��W���ԵJ�*����2.��&��gA�K.V�����<���^�N�I�K��׽���R���ٓd��'3�m�d�0����?��Mحеu^-Ը��w�{�=y�z��$iwk�;�5��|{���~%q�#ƻڽs�H�L�ʞ7���lF �=��$=�5�gv��������k<
��{��״��8n;բ��<ʹ��=E~�Y��� -����������g���,0ñ���ݓW���� �#�M���|.��#&�%���s;��>#e� L7�vy��+��do�g������Dr��(����ȈC�nF��w�6Vt�s=���NV-���s��Z�wR<&'p �_h+7�Ϧ�۱��������W�#��R����Z׸Y��{��x�3����C�3�"#4U4须���1.�R�Z��9����>�O�	f l�ҥM�EW�Ԫ�CGN����M�rDL������x�x�tD�g]�}�>�o��f����f���(��h���Da�s�n{�_{��^�s�_����V/.]PwwO�j��P��'(E)�wW�o�\A��gKp;��#XAg����-�gv�浻����)����0�=�f�jj�\;l^�t*2j�<�d��(1z,�R���*]r�=+��W6����#s���d��F��:�Ե��ܖ�\c �-)Zf�q�>���^�pV2;\^ń,�G�j랦������vr�u,3�K��l�Ϟ��}�ۄ�MŮ�����u�W�:��G��j�ù�|���=<1�M���W|�\/��j;f��xVoQ�vs��-78?kB�o7�t�}��_Pt�og� W{] �Coٰ��4��=O#�c�ol[��uj�JR�$m��)̫pf�ȱ@L��;��h�pb��[qD��q�):r����N���g�N��BG�����0���H����'b�N���h�MBW���,�0��9s���^Ԙɔ�?y0<
N��(��	�sT�M�]-Y��������v�����w ��v�W9�f�ɔ�=��D�u�8�A�Ĥ��`� ؟�RC�Z�kǅ���}0�����͈�A�
�M�X��M��0����&r}���~<�g���X�J����@���_��Qz^消�B���a�svl]f��L�A�k>;䴼S'9�?P���S��}�[��MHyx��s��8�S�����s^�V��h9P]�܄z/9�돖�ѝ��Fi��s����(V�����y�<�a���F�j;��vʳ���L$�����C������]�}{�̹�\E�>3s����8!��A�+�ķv�L�U�KY�2ga���فz��3Ge�E௷>�~��u��tK�:Qzr�p׻B^���܅����0��[�W}x���}����
_aE!KRN�n��Ѕ���w�wj"&��Si�%δ5�	��[sJ�E��f)���7,1ٹ�A�b�qy{C}1LL�g��g0����;�)m�qـ��W��3^j��x��n��2yѷEH��FӪ�4�sB�����hD�JcRͅ�0k/+���׷o��ˤ�7{���}xl2z7�-���b��>g��[��q�g�
}��&�+3F��G�)P���ݏ�}����;w�E�f�Չ>k0�m�nvB���DUS�N7�&��t���.���1㔘�nG7��z���Ʈ~�S�5�0�f{��	=@5�9�hx��ͽ�Ά@�:�o9l):�qyk�	V���l���̍o�3��i~=�sR�踱b��l3�S25`��{+*D�M��jY�S�~����mꠋp�l�Ņ�����D�S��=��B���SWp�k�G�=�=����'�v!K����{�T�=��ܩ��k��Y�n�ӌd��K�JvV
���D��3��0��e����0���'���Gӽ�i��͜�����nn���x�3*`���(6Z�G�i'�א�	�1�U�w���J����]�;�Y�n��]7L�JsWH�黻����ggcѦ�R =�o��8�=�o�91�zgi�aܻ؏�Z�:��r�<��8%}��m�O�����gs��Ӵk%��F�ʐ�¬�Z�b���҄;eE�"E�j��4��ɚ�f0�]ô*^7Ze�ܤ���/�l���4v"�λzL�w�{O��X�٬+L�����}�vU���eѐЇ�x�>nDc�Z���~=�?O$��&Y�}��W���j�������}Qy��? ���/j���zJ��\��w�V-���0�����*okz���#~��B�����%�&�9���tY�sM���|gM����@�GE��/u+p�/~�K����v>��R'uoƍ���{h��s�b�@[:$N�Frƒq��� ��!��Xnr������;Z�'��zn�0�Gp���
���
���T��g7Y��5���0BI�f�\��;5��� �s��饌��cB̒W�D<*���r�\�!�7ڥ��}�m
}8,�y>�T��:�	�w��D�:V����.X����܀jY��o#��2vh+�:3�y������G�X/�xC��︐��h�a575�(1�%TF��S�(��6�L̢75��I�a��*N��P�gP�%��|��>#����ل�k�Ŭ( @��$�1��fɦ�Kױ�V��Ln'����2A֢L�������Y�9����cc�����s4i�ΰȾ� ����;/������p��q�tڪ���?j��C']�^V[2���>�c�^|�Y�A������ A�x</A�^�������	cO)�^���|�U�W�M*��.�]�+�Iwxx ��c��\s�kY�JXF��L�q�a&F��Ɨ{��(�dVR�4�s�<����������쑾=H�'F;���V�Q�Z-b�kv��/Y5�(�H,��w�y	Kx��e�S���}���-�2�^�(���Ӽ�z�z��fk�� �v�s-���S������;�#T�������9Ձ<C+I�.dk"�r�>� ���j��jF�����yv�Ӆ�PK��.���$Lm�%��M�h]�#M�aqT�ڷt����wr������^c۶mY����2�N��ۻ���F�ݲt"��zq��]Z�x��&��f��/"�{}��<�E�3�0�8(
˻�g�^X�Ɂ�>4q@������p�[��w	�k\N�ZC�&n��ځT�s6w͸.*S	U�H��n��[4!F*i7O������RR�RG#n�+����T���Gm�4��r�B���a�U��^�#</��<-�oŕ*��;�a�������c�1��3/����na��7".s��)˪\7B{��%��;���vޙ��*��s�n!=�T�֎|2� �9G�t��$�hJ5ݍ�uM���"n\>(�'!�û"_9�'i�9����b��@a��ԅ�YJ�3MQ�̕����x\�Ƽ�^�^|Q��*��zh$1���n��～�ݝ�vP���ݥ����U��	*�#f�64�8n�*�5�<���ޯ�@˹�u0�kY9�d8<F�^�t��@�����a}N�{��u��;V��'uPb����u���}�v(�f�w5"�EȎ|��=H�y�z���"�;#��s�t	���rp�3��x��@2�p�fֶ��a���n�w�y��7��鞒N�*��&���{�v=w��q�N-�H������Y��Ls�����U�[QL&L����ع�+���ڷ�!�Y�h��O���j��֞q�_b����U�wop�/v%�p�������;y{�Q��v�y�x��)]�0�_E�����}�O�z�o9�g���]��+�<�x�t��e�x�
R�|��-�g��ݙ�A^nq��8�a���"vo��5<����{\�=��a��$z���A9�8���s�;��{T�<`�oڼ3Ox�x2�xg=в`�Wt����eHjJ���@��@��.�b�l�bYsg�O�\Ԁ��8�����l�z�t�py��Srb�2u���T�B'�z��(7^�X���̚m�k�#4���1YK��S���1s�&�������@M�O&�R���ջrq����Ǖ�0���\��8T��V������zٷ��HH@�h 
��m�ehB�1�	qZ�MvVf1�j��]�v�ba��1bј6j3X3gffSu���jW�z�)��qj��Wj�񴰍����ˋ)�y<��y5r͇�]����[�R�bU��Ɣ֤ ����V��ց7eqf�m%���$���\G6���&����T6f��Z�xxh������xD9�Xې��XQaBi��G\+ױ2�&sYX���гF� (�R�!.�L�a�Q�I�ٔ�uf�����r��ͤ���"D*�Y�[LَV_�K���.b�Z�P�\֭�f�kk4�hRi�,e\99B���jf��i�l��h�n)�Wf�qfʆe�j��G0�Ic����O!��W,�4�(��\�Fmj��h���ҀŠ7CB[��G2�
�0j�l���t��`�ƶG�+�%�`n��A������%KX[.���4(��;/2�f�i��ˆ\Tk*�,�j�i3��,fU��[لԭ	1�.��ڤB��)i���2�T�MY��bۊ��/�i��14�)I�jɫ�`�bB��L�� 6�!P5�nnf�]S)n4�6��-�1x��cd����&�������S��bkb��B�H�p�Zņ��KH[r�H9�X�-hf	�3,"׶h�u�a��۔%�X@�3��\�2ښg�V�!�&a +#(q�3R���S8�&Nn�`h�QNZ.�"�M���v�n��]�Tt]P��\�	�e���X]�i��,o,����YtP�im�9��E.i��m�&�/,(�Ɯ�]%z�.�f[�E"�t�1�ں�]�f@1s�l��uF�b��%kJ!s��eh�֢�3)Sxtu��w*��#�P�ur��,X,�]6�f�������Z�T��R�L��\0�^j�+�h4�R �"T���0��֌�,1��n�PZ����gQ6k�����$3���^&��/�y���6J��W�Wn��H���
������µ�Դ,��!b�i���*R�ڭ-�F\v��J�!���m-z�\am����:���(]bJ@��u�\�����]�����͸��J�hb�T�dV2*��n!o��\ �Y�w����Բ�H%���/U�5a2h4s���A%JSC�� #t�˵n:��# B�Z�+E��Yar�f'1�W�B�WT�ۂ3�H���d�,��ŷ�3i����B�-��-���X��r�l�(�YXfj����H���W\L0�ìz�ݦ�٪cjZ6���Mj�Q�]w�`�D�t�21��������6��&�Zғ*��e�B6V�KC��Rgj�%\��� ���5��5�l&�H� �&(ie����L7JfUƆm�����a8�k6�r�%�j���M�eC���Á�0��������8��k��j��"k���^Յ�8���b�,Y����1nԺ([m��4�:���DuU�MV����c��Y�\����Wk�!cm���;	̵�5�)�u���
�j�%�`{I]��ֺj$m�B\�m-M��-��Qf�L�(�)�u�i��r�da`Z,�u[�ILs�fY{\B�u#s(Ka��g�l��8CZʶl��IjGg7X�C2��X�M�LiHYs2-є��sl�������X5�X0�{fU�:�14F��-&u]l�r6Ы�6FgK֐������b�C8Vij�p��Z�4��1-)K]X�iJŎQ�m6	����V6KC+���V%t��l:F6p���9h'bZ���X+L���*:Z�Ңd+..Xb(�kc��k�c�zZT���]�΢x�1��Y`5u�r�]eBf
�Q06�>+|�z�`��L�Siu�1��i�M��D����鵁�v��i��$�0�`5����ƀ5V���y �\9�X�բlX�Wf���ˬ�x
@`)��]bj�ʎ�k�ٗK�%E�(��؛F"���Vj ���Y��x!����D+6�I��A@M"2�4��F����n��ܫF=��[�»E�sqe�CYs\����KEkr����m��^L�R��Ж]q�����6BͶ�h��<F�3�d��k�f�b�@.����7.�%�ך�-B˦L�	Ye����Z�Ֆlm5��v+H\$�ؠfLXl��C(�0f����b�ln���J���5����;V�@��9����VS�5�n8�J[z��K�rD�͖���]G+�vJ�nƁ���[qJ�S�ll��.-�Y b�9��chF�B��:��8�K�uC�	�څ�`�^��A�VZ�Qά��[)�P6����1#M.lu�P�M�1�jҶ5�t ��I�k*$�����.�X]+ Amn�̮�6k��e��1��9hvP����հ�M7A��k��j�R�U��ٕbY1ͨ]5��R��:�ұ5���L�7X�3;	�v�H�&�ؕ�V0h��{V��[`E��w���2�v�vykj�'\\�z�m�"�kh��.�ԡ-8�eH0�͖k��m���0���e<��,-5ŹP׭l�Ch�h�b̉M{$����`kh��ٹv��teᣠG8�����35��t,�i�����&�D��sΣ�,��F�y㥆g�v0Ce��+�ۛeNΤ��"!�d���Fk)Fۭ07d��5{sZ������$!L�獢��R^�D��t���$�H��U*%�Ж�d����	)��K{�1m�Ŏijf ��� ���S���\������4�=�g7�楹�⨮e]n��wtk�����1(˴�!�m�bk�Фb]�s��rB!Ļ2H+J:�&����kr#��Z�X\j��ũ�lf0���v v����Ka���ښ�d�4-(�!skbå��\���=jLL��Rc8����a�fn�ۗ(�x61�v����,j�N�ˑA#.��f��ń�Z��1)����!��W��Ü�m��h�Z�a��]Vm�f&�Xh�Є6V[2h��S�ـ�U÷%�v��v+	V�S��ҕ`i�i�W�s]�V[���])2�a@�*5%p�5؍a���0)E����=c-�;`)ImA�E.�ie�ζ9�Tnb��e*�f�n�ɣFn���a�Wj*�\�8Ѧ�V쥬�л��\�Y֙�Q��kk�`�иWa���f-�Kf�A�6�������ݬc���ٴ��GL�cR9����7W��`���4ͪ���m.6�gU�q�)p�/,���+@�-6TWJ�m�\9��jC8	b����CTav�du�@#�v�S�hq���:��	2K���ۺlPr]b�t�!����q��(ڑ��.��[as#�`c&q�*դn�,�Z��%X�K���1L6lk�˟��u��ƥ��wl�͵�cl Ke�ދ�����h�����6;]°rG-.�c�x��K�wV���� �k���B)�(�3T[���l-aRUn��[�Jd�2�Mb�Yej�Й7;7V�8��YUPmX5�L`U[� �i2ܳKs6Q���萵ۭa5���� T@KZ�lX%�k&�6�R���n��r�=y��1KQ�,5uذ��4ZSD�m�1.��f��կj��Ml�u1�k����)k�n���1�h���t�P+��2b����A�v
&�-��3u�6.hGPb�V2�W�%6����4�@7L;)������U�-s�:�nŬ�ii ��qd.�q�.�T�4)k�� -a��,tt��Í��-ҖhDHڲb���I�����&��4u��cD��tw�ca�KBj��9n6�`Yv����v�7Lǋ.�@�D���ΰԆcn��X��]mKs���h���iH�
�j�f�X�̴���uj��,%��4t�Z8��+��fO<�t<^#����:���/c9ֹ,2c,ʍp����Tl1fҠm)	D�:�a,
�J�T=^RF�mr	z�[6�шM�J]�0){K�أ�[�J���]�훞�^U��²Z�M�L��:e���J���VP�-��`*�x%���ڍ�\݁bF�U�Jh���S8�bZ��
36@h]��Z�Y�)Pl�biv����Ō�\YML�0��P����+.pBm�R���-#r�f�V�b�їZ��
l��"�(�є��nԐ�BDJ�z�At�X�b�Gh�4.Y�8��PXV��uWJ����R.\l�*S�������Mk�)z�2*M0�[���5�bR+k��q�\FP���	�q��@��{v��fMG+��)�Yf����b�H�TԤ4+GCh&�Р���<���V�M	�51[A�
!hR�L�	4"�Rg�f������Im0MK��*�`5	/f���f�K5�]�b	L��t�0ɧ�@��F�fX�E�k��s,��]t%MlR\̕��.U��4�\9ҍz��F6���0m�vh^�K������p�!n�i�q2S2�-͘��F�F	����eXؖ$���A]��=e�� ��<irWk���>�k��`��K��u+Tu�CK�d�lB�SV&��%�tDl��ko5	��Fl�R�4�6�c(��U�k�l�̡�l1��̣-i�tl&�6��ʲ��eЌ���-�Aق2%��(�lZ���x
�����)d��M
@�,�f�;呏UֈF��x@�Um6�Ζ�6��!��f�.�̠��b�[���WF��0L�B%[.�XŚ�n86�a��f����b
�km��qe�L,��!�j8��ukX�Tm4�ƙ��=m�ۭ��p���52�[\9/d07��y�K|Zf�*ZT.n�\����-�.��nq,f`��x q	�@���RZ"aEŲI0��I���J$$�"����Ƙ� A�0cDQ�$`@�3D�CRd�S&cEs��F���D�F�E�P�4�17w �3hJ2!A�D��)HLIR,L R���(�0X!(���܂%N�r
�H�I#fTX2#1`�`[ d(�@��lR�23	+���cL��QIcE-�wt�FK ʃc':QIb�f	�D��&�%�*!�%PY
�Iwn,IRTX`E����)����Б�0�*B0!2l�L��%&�`6J�ª�7��>���&6���۫�������b�mi ;�H*)r��Y��N׊��l[�I�W��iy��6l��3���<"���,	l;P�$�t�Fme�tHQy�6Zf�4Q�dҡt�2�^��5е����Sb�14�mu� n��[�u���^ή��r�]�#��m���^��`�y�֐�Wa��3U�KР��7F�[���W(�ٚ�&�ˉKYKL������+��kN кf]Bɶ��1��T�%�Y���SHYi+�X]��!`a�)���X�V�� 0Sc�Z�Z�h�h�Ks��V\�̰4�X&R�5��C�X֦)n%�^f�cb�2h��G�y��h���hLׅf��U�	�w6f�4&e�F�eғI��F��ř1E���!K�%Ś�� 2l��ԙ�����)�(T�%LK*F�d��Wa�R�-�WZS0*���^��l��/fW���덅�*b��/��m�W`٫ �I��i���W,h�:����m� �J@���H�,�cλf;K�I��1D�{WYe�Ifvwm2<��Tsf�50.�%���]�.H��;D32,hٴ�$i+[32���ZG0�h57Vdʴ���c��+WC*���`�p�0׳.R�A�:��m�m[�@l#���1��u�p˲�Ձ"u��hKә��:%��F��0�@.jb=iln��kH^e�.��a�)�/�f�yA��b0��Z���f5�i�&ک`H4��c�Bf�ֆ�֑5���,l��\,�D���4֭�eמ��2�S2���1Dx�s�X4�u�jh:+31)2<hA�B�lŦ��c],�ٱ4SiGAs��6�9e�Cp M�vY�jڕ���:��,��k
e6�jim��Fj6\H]5�c	�L�I�e��҃[��ll��X1[-�����F�+Cvc��Y$��&��R���k��FZa)cVȬD���"�:��U- ZZJ[aa`��)e�2��BB�i^R�РV��YV"�-KKh"�T����� �T	cR��¤:�BX�^�Q��Ћm�K,(��F�Z*�F-�B��U��Ycĵ��Z*�*#�=��G�X�[Q��#�c�QCv�4�DQwk�����+y�����{��R8��٘��i�(G��V��; ٲ�T-F8Ȩ<r$p��n��An+*�3ԏ	!�L�!ص�{������j8��k�Hv�E���&Jǳ��m��u�	݀����� 6�R����P���T4Nؕ� ���Aƀm�7��/���L�X�ńc���@����g2�1�NdO{te@���p뢢�{B��Ѡ��!��!���� A��m�
����$+��y��.�w�Q�5ڤGj�@ڞ���h~�65/���5��,CX�u���VQc�顮�:j��$J7K����Y�w��X�� >m6*k��d������g�̨�ذ"�{���p-� �[jH}Jg���Ô\�=U�q(lӔ�t�L��(EB����t���<�Oʇ�.�~��O��㙺��_zUR��Osn�\S����d A9���df�zj�$O{te@�r�"nȒ���{	�Lf�� ^�� �7���7 �8#�����e`r�;��M�Bq��w�&{W�sA� A/�my{��3���{4�ո� �Z�In�-��*���т�z��''�p�D��eC����� �͙�PE�D[jH!�n&�[=�[�RQ��rqM�Ö��F�D��E� �9P�	�@�Rߞv�������5�M������F�ZUS01���X9��rP�2�ٞ��7٥���A>A۟O��f�����p�{�Gq3�dM�W)���A�m�6�>-ǆ\ѓ��}2oh¢��;Ј{lU������F؜��Aw�1��Co0�B��^G� B��qG����E�D�fGޮw8��dӞ;݋��ؙo�R�>�� ٽ7�ne�"�K�J]'����U�)�M̋�S��w���ap�GD�s��=�cħb��k"��-��� �@@�3vD�[�A����S���쉥�"|[AE!{7��mq�
N=َ��j���$���,��/ǲ�󗛿 |p�$���G^���P�e���A�˚06Ĭ��Dc������7u���\��(GL���۲��.+�
��E���gU�jͲʺkVkA�Q�Q��ڽ/PE�@�mU�\Xٌ�/.B�n��A�3yX�m
�Aw>���@�܉Ÿ@���6趺<\��p�Z�z|Fj
)Y��yo��Rsu�q=�H<�E���%�3Rn*�ڒ1Ǜ�@|ۑ%�D6��v���i��^����Z06���A.�q�k��~-�"ܳF㷫���J�E�ބ%��U��F6��R#��*� NT C��o"�樎nf��A�@��mi���ݕ�l��+f
~~k���S���*�k=}_}�4�3�8��r�ۏ�7��</R7���ڞ���ڂ6�H%�@�h Cn�2���X����^�Vj]=*���)9��=��j�@��n>m���>�����޴���B�[c2�Slfպb��W\a�6Q!5&\f[�j��?y{~�|��{2=͠�EU_[9Gz\6����d�0���0����2��ϋh [� �����ɛ�}]Ń7K�S�}�F��fT��n��r�"3u	�=M
ـ���� O�a[@6�|[C$�ǧ��I�l�i�!I��1��g�z}���"���6�w9Ff損:�W�-�;�� 6�55}lD�]���%>.��ص��mŭY����'�c^n(6ԀCq��î��^H��F�)z�p(���ʑ��U�{* @f�yy�+�P͍bx�t^�t�<&\L�f6���I�b4C�n��ܣu�C�cb[=5�b=;����1r����U"!b�x�FI�����JJf�^T�LhP��m#����c��\V���a-�,ÈL�R����_<�ď�	��2�)�%�[��nÊ��a8KF.ݫ,��j��Ţ��`�pn��8�jr�����:�g�ܭ�,nԦإ"�b�n9x��1��0��J�^0��L�Y���������m�	���F9[)���-���Ŗ��	jPÉeekH6%���崊���l޽j�Q��51�|��H �B �9��m����UsEN눽3��sC�Hgnn�S�z���>m�6� �Ui��٫[V/Ʈ���_[5Q���6���}N�#۠^j��������Ȣ	m�7�p�%��I�[/b;�3=ӡC]�f!Q��]�9Pf�-�6�!�2ۻ��c+h.��� �������+kZ�َ�$���3ܧ�S� ��X]��7�O�n�n X���ʷ���	���cj����ײf�j|
b':A� �x���|C{�˰���<zOn�Z�B8�[Z��'l���	��l�p�Qo5$�G�!��>��w���� ��n��V�p(i�9�Tw�EW!�ƺ�c}��Ae�@�39	��A����An#*#��Lu����e��۞X���{ݾor���ß*��!2�[+U�]X���|��6��36��
̸y���-���ըq[3����M�֢�J�$�����RA� [��5��f�0���H����x�ۑ �nE����rO�یSk�!�#+��N=�-���n��k#o'g/{�-j�VF�n͵"��D4Ɯ�*;ۢ���* ]
L> �݅�h"s ��[@6�m�Gt^��
��嶂鹣uX�/��M ��^������T��\]u��L�B#f}c/3e��v�vS�Z�6j�5��
ZĉtM�6Q�~ސ �@@�3z|�X ��f�!�Bk\p�6Ħ�����D�lQ����O��A�y�S���m�#�C|{!x����].4!�9�Tw�ET�ʀǲ$��:dU��
�<@wjwcɴ�m������!�s:����0�w�g�����7v�^u���L��
�{��hv��*��5�u��m�3=��qG�ۧܞ���Zg)��+D�{�c�A_) ���q^ ���vӤ����4��� ��^�!�����V��P�	�H p�Fe�K����W��7W���ڟmpPɎ"�լ�V���Z����`Ә��{tU@�r�"1�p�9�۝�7��|�G�J�~!$0�KM��T�*�U%bG[a��;T.�X����3����O���CngŴ74g�Z��'�&�\� FͪWu�+�z�@�� ڒ^^n"�2�_G�wa A�!�u�u�&s6y7s�5��pn�kt�3Gbz;��Q�A�� �=�[�A��z�LN]eH�N�bX8�B�}�&�r�"=� ���D6�F,��JyU�J\o�#9 �[h!*���H�OB�ou�p �g�{��~P7r�����]D\�	������H�b���v�.�\��pTHY�ǧ_��Z|jK2��{�z`�Y>4�@7ܧ�6�@�� AmȒ�F��;�(�f�MՇ��Q��ȡ�}>ۄ�r'�͡}}Skޮ�Gw�xR�幎A�����[�j��ԻG2�;BҮ�v�δ#�_Z����H|����%�����ƤƗo��k�!��7��TQ�z�D���m ۹�p�:�Y�׶����^́b*�v�Al� ޼���RF���
�T���#���Z�^{[r$�[Cj�[���&-:�ݎEwA�}\�a&��8�1��m�O�A�{\T���c�^���#2�nڑwscca1���F蚏\��E�6mM Sm��,�Dk����Kq��۽�8��E�f����6��UU#��(W�b^�1�3ڤ�p-�ʹ�o�E����.I�X��~�w�W�1�ucrq'��*�H�Q�'q�۷�)�����9J��9GV���g*uoi�h�b��ke�Θ����K&�;A���k���)v��-�5i�\��#��&�թ��ʭʦ��J-M1�*�Y�V,� ��ld�]qZr�����lhA����cD�=\GKnP�)�8jk�CE-��
2�1&��f��-ɈC:�)������%xY�TK�e-��Vı���n��K�	c�&�32�\}�����6��۶ɠ��7(,]1n\��E��er��)P�c����,�����'�X�|p�-����ۃ*2��Ba'ޑ)[4��5�ۙ�� ��>���ȼjH5S]�wG�c�A���w"�C���F��	ʀ�A�D�����T�duo&(
�����t Cp!��!� a�қ��\��Gl�$�x��nc�|��p�@KmI��^��� �\�6<�AN�p��ʋ��P��NxH'n!9��J�p��cCޟO����[��jH-��ql�k���;�k�����c	�+9D�U�zr �7dH-Ǘ�B��0��N޾8ڢ8b�Dj	�	��f�i^X��j�U�Xk-ip.�--R;D�L��c���p�#: �ng�6�wT����{���ֲ8��z�I��'�/  ^���Ԃ��p>L�F�ڻ�!���oH�O7\�^h�F����5I�F��&��OL���$����_Hi��q8�UZ�g"�a� n�؜3y�8�� ��
WW˒�/���� ��[@6�6���b�3yT���ۏ#xԂ�Ax����T�-���z�c��,��p`n����r ��[�n6�}�VR��WՒ;��i��>!�]�-����&N�����A��$Z�Um�Z��@�G��jHmyp ��������R�+X�H!�֌�䫾���B^uA�h Cn}>-�T�����!|xlW@ؙR$��2d�U����3d��`"�Z:��$����
�����j?�>�^������ȶ���U��Vp`n��B*g�g:j�ntsP$EVH�s��mϤ[��:�̠v���dۗ"H�����e_�ɽ�`��Y���H��t���J.5� �J�;Rp�$���_�L��:�4+f��ܠ��Mj�f�c�	�juy?C��ջ`�S݆a����`:I��]_a�p�\_{O�ϴ���+�Ru��mS��H�IV��x{�1���f����o�-4eB�}�����<�rV{������nv�Y��sg�%�p-�Z�W=ӄ���}����7Nt��X�z�����S��;���w]�=gN=�e�]~����uQ��������5���V��Lj��SQ�==k��͛;o�mٹ�:n@�>^Z8T7)��+٧s�҅��ʱ,hnֱze���ف��k<�z�M�m������C�׳��piy�7A7�����'0�nM�r:c�zM�C�3�px��s�s�j����>���h�?5ۆ6�!�5�ҵ�*�\ݽ�;.z���r�o1ӓ�<trk<[[��-��z���s C��_ZS��֏&�x�<f:4���S��j"h���d�mttO<=Ъ2'ˌ��t��;r��r6��gg�u��,�fM5�vi	�ڄKЦ�ލ�������J���y��3�ܾ��\8�\���B�څ5H+�N�������~HG偮��g����"]�m�px{�g^�ּ��]�h���gṱm���Z<3���ݽއ����\���I��zl�r�1��+�vܜ��O{Rn��)^~�c��N罺�1D�~q�m��	uA�E�=�o����\���ͼ<=�W�����V�b��3I8��DSIsd|�o]���?�¥Ga���k�S��5	�^q0�$3*�LFF(���(ф,��B	&,Z(�FĚ�h�h�k���b��I�i$��-+&5	a0Q�D, Ѕ��!���FHƂ+&
@����2Z-cBb��#@b6#!�̢�1��!I)� �61DK&"��͌$��j"��52M"(�,U�1�cD�$�d��IELVB�ƍ�PIQQF�X��!�Y&b� �Q�RF7wRVց#h�@ɊB�D�d��DTUY�5�<9����<�H�	>	ۄ����"� FwE�e����.�^�[Ax��[j�*�镬3k��W |]@Dwja���<]cN\y�
6�H>-� ��^6�?-�"6�h�����`��Ɏ ��^�h p�Ŷ�p��՟'����0u:�lJ��ⴁ�6e:�f��F��)u ��͘�0L�(�/ϳ@�囈{��� !����{]u6Bs���B��̋� ��������[� ��HI�ķ�$�{!x���"�U؉��s�p]G�`w�>o�H���y�kX�� �ݑ ��D�@���|G�C=6��;�T����O>���&;��RA��n<�[j}�^B�X�}ĸ05�7  �t�: ���]Ĵ�+��Cd9���p�m��!���Qz7R���%_t�Ӿ��˳]q��e�O��L��=�iڄ�b2'df&����U�ث�4�/'����^��pmz�^n#+����`��W���WW�E�zf�4��3PG2 ��#z$Vv.W�礟�.�ٜ:Sո�h�������y��4�e�P*�"eD�N	�Dڂ!�3��*���Fru�D������#1��7�[Ax�@�Ԑ�8��M�N�ٓ�����B�9[U�KL]��]B!9� �p�#�����H�H]�}b�\y������qG͵ה��[ג�0�]�L4cp]w�>.� A�����Cp!� O�r"�a��0�!��Xm�Su{'Q���D[y1�;�H���t�y�8�Ō�C�"=ܤ���D�D��T���������1�]�޺�6B[�A�"��w���he����o��ɥ�(U!w�@{��c��zur��:q��/ݔn��k�^���C�8s�U0�Rc>��p�1�e�|.�u�7����ב'������XuN��-[v�@�g�HF����4�F��6�S5��u	��h�ݵ�����qF�#�f렄�+��bڋ��X�4 ����K�mk�8f%n"f��Ħ�vd��lS9�"���l�&��@̣�j���1�u���eR�ڴ���K�m�R��.+�-a���H0��m�ye8�"��d�FX֤���W
3׿��쿍�u�5�1hY�c
��J��;B;�]nͶ�[J/���r���|�Sws|t�·�R�:�]@ܚ��Yt��Tg4$��A�h"s���mT��f��Ep7�|G4*��QS��D[Y1���H:�@���v���׷l A� AmȒ� A�CV	cz��V�S�6��#g���^ �Aۙ�m��"'Y��/S!���m]�\t�;k�;8.�qwZ��b���j�������|[�&�^6����=������ʅ�ô����O�:�^-� �[j�d�7tj�a��bd��L�¥�pۃZ���W&�T�A��L�82� L��A�D�� Am'��d&�ҝ餆�(f���Ʌ��Z� ���z[^n=@�׬E�7J:Ws�y�Q��47��%��%�=ǘKw��ik�8�A-O���͔�[�ޮ^����(V���,����r>�.?����x�мA���]�]�5:?mFK����=��ݻ"Kqr��e�#&!�\�"u� �^!��~�7�,�sbp^�Gk.��B���t��A;֤Fj�@����ׂ{m�&�q�+��5�$���h*ޭ��2�zi!�F�H&� |�eZ�'�T�
o\����D[jH!�n+��{sy���Mg)Mg@յڢ�j;X&��]�϶D�� A����멥�#�O.��fɱ,�J��ma�v	!�c��E���Q1$f�	�<���mȟ�"���P�Y�J��s�U�	�u��`�|��ބA������	���X�R���7AƄ�u�ye-���5S��p�A�@��O=�s��������'�T�|��q@�[j.�i�-��z�m+��*�;h���Xg���8I����e�}&��sR�!�ۛv���l�N�2��@l�UD9�s�q�eN�J?xx
���]שU�Gk��]�D>�$����ӳ�
x]�I�71 �����x����F7v�emZ��\�Tj�d�~;���jHm �-�	�"An2b`�=�`�q�0\��.���9��
}��H)�yP��$g/I���
s��7� ���~މ:���?o����l��9�U	��ail$ηv��V�%u�Ze���[�W.q�~��Ϫ���I
�)7ܰ4�Ĕ�XT��$��9Vɡ��� =� ��(e�_ܻ�8��W+���X{�B�
C5�_>�����`w괂�`RAJ3�h�ld��B�
ACCr��XhaI9�XH,�e0�*����X�~_�u߫yĂ��i �|큽� �!ϪH)������~����u|�03Ul��I �����6���P���X�[#����ί�u�&�
"Rg<�4��i ���i�AHQU;V�]F$��s@m �l�Ü�ZRA`s�i��q�h����dl��Q��2���5��:��%2�sڅ����r��Xi �9�{�
Aa�T- ��09ʶi��
����~7�+�I��M��,!�JH,9ʅ���ݫd��H(���,O�����;�}�2�jؿ��|2���
A`s*�
AH)]�[�~��_*��L�H}��2�^�������:�e� ���[��9s�q �f�ѭ���@��.x�T������z.��ff��3_�� ���L=�P���P�v��Xi�$�9a�6�Rr�h��r��X�H�� ����D�r{�p�$x$��<	�V��R�?2M��σ.��) �PII��`i����p�AI�)��U�i��R��@	>������5R�� �p2�U��vb�Ѹ��̩���VhRW����\��2҇U�$�GI!UP;�ZAH)4g~�H,�d��B��JH(Ta�V�o��{O��)�﷭_�i5��:��'/�sW�M��f0�j��I�G�^�Q����l$��r����
`s�l��I
�)9�XCbJH,7�z_u׾k��� �~�H)G�#y������q��le���ϰ�,=�t�R*�s*���I(�w@m �c%0�*��sך浜����������j�RAO}��bH,��aϪ��������$��S���� ��9PI����b�ڎ�*�/���2M�]�][:�I
Ro��4�R�P���؅09ʶM2�
	I�r��`�Aa�Pi�AHy������
�ZAH)8y�����;P�=�) �L9��Aa����r����<�kW��m ����6�Y)�Þ�-@��X��Y��^�A`j4�Sϲ�ٺ ��ϪH)�@�9V�R
II�r��II�9P���B��*�<����|��a�  ��@	>�}߳�<�N^���r����Ptt�R�V�]F$����6�Y�d��B��II��U�v���߄���;sD}q��z���K�H����o57�1tn��)'�'���K�x��"b|;;�Iի�8�7ʫ�5�R���$�ͦ�M�6�k-Md���K,qe��ĳ:��p�2�+"�̎�mY�$	�FYiv+�5��[N]����,֥m�(tb�1.���0�o��)X �kw=�M��U��䪥^:�6Y�i�,��ͥ5(�0 ;`�����ɻ5�I���rq�k6�����3�R�a�;��%[�f�0�E�m�����m0�#���3/Vh�?|��S��i�6P��Q#L�
B�0��Շb�Z�t�%��g�x�S�y`i �~e0�@Д�XϯI���
s��6n�)�!�T4�SU���3|k�Y��s]�][:�I�3��{���/5��JJ��HdII�}�$�B��� �%'9�L�$��I!P���U�L
H)��E���yg���x�Y��L3�H)��U�o���yZ���v�Z�vH)��âH)�=�Z�RA`Q��$��
s��w����+o�ψ)�C�*H)���� �4���`i�) ��*�Rh�9Vɡ��P))7u $��~�d�ϣ���c9��)8��|�뤂���ʴ��I=���7)�9P���X�ZAH)9�Xr!�����
��Ϫf���{���y���^�Q����X�RB�CI4Ws�L�xWƳ}�|����u��
$��;`i����f��wϼo~}���q ����ղhe$
�����AH,9�GI!R�9V�]0) �s��H,�%0�*����u�����&�^դ��q����|;�}�^�]��
j���!���C)�=�Z�RA`g*�M$�9`otAH-!�T$�A��v���_I�,pG�Ĕ Il�F:,fք�ŹtmSKs6.Үm\�E�qs�5e�[�-��U����)7߬!�$��ßT- �Ѕ09ʶM) �P���,06{��w�=�n�2����*�R���k���ܣ�߽��>���������Ͻ�H,�%0�T-$���0�+I��RAL�,$M��s�@�J#�� ]}����h)��no��2m�������TU�Ct���9�{|;�2h�2�8�sq���׽֑�^�4��6)WP���P�S�o(�{��	_?|�R
AN{���
AitxI�љe�xK�̓{< ���gc%$)%'<큤6$��³높
A`s�l��~�}����m �RRk^X`m��þ�j:H)
*�s�i ���9�6�Y�2Sr�hhRAB��i ���鯗v?�d��*�U񘝏�(�Ek��m �Te0�@�RA`Q��$��
s��6n�)�r����@�9V�2RAC>��n��.�_��m;��C�JH,+9p�AI�)��U�i��P(JNs����y���~{Z�_�\�]�Aa���t�RU�V�]
H)E��q9�G^^��>H,�d��B�
ACL;��Aa��S����Ad��Ü�Z�����A`hi ��� ~|���+b֏G�4@SH)�r��������q_9���.�����P�%'<큤6��
3높
M!Lr� �%'9�'�:���|��
��9�7$B� ��Bݘ"�ks�0.5q*chÖ;�&� �XYt�Φ)��~$��$�P7ڴ��I=��I�)�9P�4��
0�+I����^{��|>�n����èm �V]{{�����M���- ���� �4$�;`l�RHs�$���*��%$(II�r��RAa��v���y��ZAI�
`{�ZAH(�I����~߾{;ǿ=�\�\������!L�	l �s�BBs�����������|��9톘A�v�,afXB�3,��A����kϣ�2r�����Dr�ǵ��QEu��g#{���7y���C
/�n��c	Z&�����X�����³��.z��g�Q3�k����<N��%�0E�����o� 4��Lʄ� 6׀ 7�\b��ݳ��w�ʀKaoۄ4!9ʁ`��f��\���|>�κ�n� k��$��	l �|�z���y˽<m�ߜ�I�r�e�I��L �˄-�̠3��츋s=��x"��y����k��{��k��$̠�0��~�!�	�P,`L� �g3���{����Sya��Mm������B���,nbM�Zk]�1TS�u������eB[w� ��=� 7  ;�.a��&]|����*��!^k�������p/�	�a{������C3.� ̠����P���5�y��o���`��Be \����N�������su�_Xv ���-��XB�3,s�/��8��M�({�@-�y��$�ܰ�aʄ-�̠-�32� 2r����E�MVS��[$l�-;�������̠����4�̨��2�,`�p%�k�y���`����	�� �`x0�!�P>���̮k�y����`Ta@6�^ �|>iLL��k� 3U���T��%��w��X�2k�Q�e��Z|P� �-�f���J�tE.7q��;�nu�����������&y@\`Ns� ЀfPX��̠�0�f\!�&e@֯�~l���C��  �����h꿄N�����:�@��	l �ˀ�`x0��q�>��KD��7�Jf!B�mhR��n�Rh�5њ&s4#�bqEt7ae�us��j��yA��
�ya4�ڄ-�̠.0�32�<�{3�)�s��ܟ�r ��xN��u��דS_xP	ф}�B�LʁhA� 32���
eB\a=���y�����߂0�g.hC��Ç���W<���o�><�`T�$��pY� �p���}�Bs���;Ac,��X�	������3(g�y��Fg��:ft]*���D�O� ��� o� ��L̰5A̨�2��g�����|��}�9���0���X�{ڄ��ˀk�;�:w�/;�s������e��9���p�x��@yP8!a�T �ˁ<3(�{��	����i�a~@�� �ܽ���i��+ǚ���b7�	�a�Y ̠7A�ˀ}��s�׍��f�(����s��_.�{ʌ��oO/�,[�G�Z��]��4H�oC�jy���G�L�l��/}��[{xg丵rV�PO2�jBhf���j��_�w�$T6�Ϯۋ�Q-�4��0h "N��-s��1r�)�~��T�H��T��X��0u��������T�!j6�g���o���w�����@��y*[��ut�o�d>s�w���[���ݾ΢x��-�-�������u�$B�^>���[��p����
�on�;vBW'�x/)aa����JR�8,�i�Κ[�X�;��v__{�<^�ٗ:��	h��U^7����Q:�Ί�`{	+5VHz�n���9_���,�>>�ם��gs����̺������dz��l}}{�<_�u�zoK���َhFb�]^���+���� ��ٕ�2O{;��[�����yy+T���*ZA%�0��n�ڃa��3.{�r��H=���<po��η����.o/.�O���=��r^��(m�a�Q��p/N~(����=��7ŕ��4$'��"�x{�b!r��9�i�Y��'�&i!o���b�N�4�P�,�c�5�k�×� P������k����U<��es^t�o�:�~�ע�ȖUHWq@��(���N�"��Q溬�����42}��[q��N3�~Ǣx��A�C���=�w���7}��xX�VW����w"��H��y�z��w�Ю�s����q����r�co|h���}�
IƍE�hѢ(�ڌ�L��3(�lflP!cRh����),c��,�$��(�ъ�&���+I��Dh�Q�b��b؋&(B�ѣY�Z#b�hѤ�b��f��+Bi�Q����E���شcQ�F��MI�&h���E� -5�b�F�I[mH�Ky���n�gUռ�.�eɌ�)^��!`�*�˭����3Fjf�X��q
ƊX/���x�m<���Rm�´-M�x\5�c�GL]s3ģ��4�˦��$%e�+��[UZc�:4�\2K*�MV51�BP�"2��)�6�`c
�FZ�7mCn�,�5�WB�cm[��������$0�膖���j���+4��\��[,�i*6�ڌ�)iy�L�X;Z����ݔ�L�cj���#Y�Ir-��H�:�0�F8�P���z�1B�B��h[����m,b����5�7!lt�4.U����^���4ˢ���t#E��&��6���K�5Djf��L6jf��[͢^��H�jX�Z�XK@(�1l��t�aa�
36v,e�������uu� �nJq�GR�a�Jָ���եں��k�	]�������1�K�	n�V��M[UCl��W]�P�QƆ�wh������k��e�鳦4��nj,S�tR�z�R�@�R������֭T��(�Fo��yl�B��n����E���y�N�gվ>1��.�vAD���,n4ɲ�3Ym�	qjvX��囨i��l5շ%e]*�V���hC�fvЈ�5(@���A8`�)�yM�kzb��XI�u�V��
m(����pS�q��i�Cf��)����ت��%�p��D`hՆ'�K�'��Ŕ!j�n�&�"m-���yTa�,l���m�fX\��m�v�Z�3UT���j׀X�X\]3]5��n�%�]a��T..*��G�̓MTL�9��s��	n��z��36!�L9Kmr�7[.�YCs�`+P���2�MccA�Wa�&�.�@؊�t85�r��2.�6RmW=e�%	�� lp��KM�$��cc�s2��֚� �U۬�v��k���De��[+t[�Yu�W��&���1�be�;T�pGD��Ŏr+06��kWl�5]�[)3��)�d��_�t���� 2R�hg,)A���GdeC.)�ԖZtڪ�2R��� T8MvX�ub�5��Ku���f�p�d�$ԙ%��1�k\HՆ��V�h�n���l638Cf�@�(BR�-!�f�$֣�kȒ�拹Tl�t%2��ՠ��.�f�s�R�拱f2�b��rT�k��(Eq.���MHv�ke5)��R��K�3O��?�ɭƿ�K-��
a��6���]�b�+u!K�C����[֨��� >��$���a��jЄ̨2�7�{��]�xo����7@�ã{���i�V��z��1�r�&{�	4�er�l ��a40���������{�v��� �<�\�;�?๾�����(:$�2�[w߮Є̨ᯋ��k�����n�>����@����%� �XB�	��	4�e@/�|��x$N����O��������x"7ۀ�B&eq�32�@3(-�/�+v�8��;Ð=�@;�uhB}ځbXfP�ϻ��]�|7�}�k����ì �yP��<+׾�ޫ��r�����|�I�3� ��Al �{�XM0��p��&e 6���܊��=����wc�1�	u�'<��A��y�ڄ4�̨̠m��5���7�e]�6�b�
�Ԛ���Q�PXq�p�2�t\�*^�Z]j���XtA@�ʄ���� �^��� �����p4����*�� ����s���\]��z0�f\!`�{���ˀj ��<��n< ��J�c>�q��?"l�0�G������AY���M�v�HTy��*�ݭF��^�����Y��4J ��o����>���y��C����@���r�=�}��?;��o����n��W�a�D������F� U̴_]ֿ�dx ��n L �s�XMFs.�2�����^ l�80T�=�g�>��p����<�$���A�s�@ʁ����c ��0�~����ǿZ��D�� 3�`x��� ��{�����}�+ʮk��A�Dw�	��������Wӵ���s�!��P�
�� ��D2�lA��!�	�P>�}��w�s�c��!C�@:��Y�[G��L��� G%�=���<=l �ˀ�p��ʀsf���~��/ϗ����k)v#h�LGjC*�Y�Y����A9�6�&������J��I?��܇N�$�>��a��B��̠-�̸��<�}>�������9��y�A�+���}�ܫ���A<a���D&eBKfP�3,5A��,�9���c�3��/��^3oM��j�6h�O��fQ;s��۞��z<?x��ݴ����<W���ߛ��>��{��|%��Y��U��I���{����'�bBgkXAk�{�c�q�rbE������W����?%� {��r���z���%�j�{w���fbU��b;A.��[�U�e�&���f�=��:���e�-?[R���{���ᯞxy�O�٣���82�2{WVb�͎E��zTJ�^�����K�F�����m2�f���F�\�[\g�7|�2��¾3nv��PN���x�Y���^�u�����{9��ٷ�f� �.�/9z����r��2�T�p�T[�f4n5����(��l�̡���f��z���:�S�j6h�|��3#33:r�𭌛}¥��d���
������u w���m<1G�����;Y�4w"�itӣ����x�[�o*�n����d�=�tɽ��=�@�;ڭҦ܊�8���0܏��<=�Oe��r���rәo�I͍��3��w9�<K�h��w�MpP=����fYs;B���n��Èu�@�e͔��)��hZ�P��75Z��
ķ���s=�۹��Om|j:�il���B��Ut�t�S�7��@fG���-���>��n�[zqvUÞHr��;���g6&"Is�y�t��]��o���,ےT�[�����^��T��e@���������hfWm�u8��pެ��uz��9:�����G��W�|��=vi����i̶�1����F�:��[vqj\T�D�.8��3Dҫ��u�\�W��X���b���(#�XƟ.oԀ�Q�p�U:��dӷv��ߗ_����цҏ\uC�+(U6&k�{�x{��e��(D���eKɪ�Js��&���h�Q35��9f�`L��X1�$�eܦ��]���jʹyp���d Ys,�Pv�cv��P^���eGi��gi�j�]����^�l)^K���O�b�d�����j�bcDҵ.V�n��Ui՛
�!� 4(�\��L�*�hƶ�Scn9����^\f��\+eeSc]P�&A;.�F��2܋��l����+Yca4tf��њ�+v�:�Z�)#����ڡ��{��xc�� fb���E��!�7�&���rXU��:��̌�C2*��`'K����]k���T�Rާ���Hj;<귬įWGt�C2 ̼Q�Ծۢ$�K�Χ�:�N��8�٘��2l�����9ac��ِ=��Jw�|����#\2���sػjɑGq��ݴ����݃���W�_Ǣ�S��ʍ|ܪz�Q�|�y2f@�R�~��I����o*Y�:rJ�$�]c��r�t�hp��#����#�>�9{ۙ)���&2;,���,��w���+��,���v�f^H���Ց���A��F&�e�`�z-��3m�#V�l;�b���ـٹ�w�d"N�6߀esoxG�1�՞P-Td�Y1�]���=�_}�N��Bjk�ߖ�q7��B���pn��edR���]��ffP̎���!ۂem�oR]��b�U@���-ǳe�rә�ާ�����)�������cV[�ʙ'y�V��ifEod��;�${3� �c{}�}>��\��^��u��B��Nn���6�!!_=1o�kPY��bpᅺf���ͳ�A�������Uj)�wI Q�*�Y�6��-9�����)ng9��U�L�������a��i�m�-!��R�<Ov:{�/��	����za]T��]��{3���Q�1[�?O۟Zm?[d��{��R�8c���w/����T��L�&�T��=�Lfy��ҟ���7}��V�©;���?Ezl-�.�����bb��Q��W�����[��3zb+"���SV@�2����uf�"�P\�R��t
ֽ����7-��1[���xS�#�C:R�"S�@�j9�~�Ne��m���'�h��/��<����[`{�t?^?[w-�;�O߾���o���CR�GaqZ��HRh�1�&���݋�kZ�1HŲ�����&��|�g�pf)��7�jEs;p�:���dN`�^���-?[vS�L���8�w���`���뻮ǔV��MF�TQ�O���ӵ(l��e=����o��-��Ȳ�9��g�L���׍�m9r*��X�P�GTԻ���3�����v�Ȯgn�˂' C=����H4nomS��6=!�b<�>w��١S��N�SYV��g���P�+��9���oj�;6%����{����s�c����k�N}i�m݄?�p��4-����We�MF�h�ާɸ���~���ߦk�o�ZnM+5��P�#�%�0]�5��F��1��iz�hrl-2{�>�}��??�s?z��?q'��D��f3H
��kXs�fFdfb�t���u�+zi:�yь��e��ShfLu�Z!�N[7ާ9���Zs�O�ݷp:}߸ȧ���7�ɟ#�aO~�9i��Zr��VM��'K���~��֟��@v����jh������k1٣����z����3#1)��͎�7g}�ڀ{9q7v�dO=�(�e����ͣC�tS٪l���]u��xn�W2"ؑ�pwOбáR�!�x��{�ZlY��@䏡�Q�����l���IӤ�}�=�a������q���7]ڰ �X�ŶZ:�Gle�tM��!+&ŖdXYr⋵��,��д8f��:<�346�f��l��Z��en�7��ln�
���f�����7n�4�;u��;6� ػ�3f�EM-��kX0�bi���1��qtMݑu���W�6��"�	p��K1�P�6��{&�Ə������R����(�)]R�f,
a�l����]����;o��{�}�m����z�[�v�p�c�g�WÂ��}�ffe{24]�2!�ѝ9���p��3y�#G'54K�-ǆ8�: .6��Lm�
��5���31����B!�Gn�dO=�(�z���ٙ����8����K�Z8�����o���We�GFº=>L_Xs���3330�u�9
n�p�sS@��n=���0�b��Y�u\���S&���!ĳ�,���0��IDf����*ܦ�v��|�<����f@�f!5]f4>�0�y�YFz�LE ��;�)����������?a���\��Ǽ�����{��3���^S�i��Vܑҏȏe܉�y��ESûI�9���M���αJ�n�@���E_� &���{u]u��Lmf}&vV��e���0]�;��N�1�������f 3#َ�/�qh�sV�F��54p�8��fdϷ���GulfoH����;�Jq=�T�Y\��%U\@��)�n<�3+ِdff��X.�W���];���gI�������fӖӨ^���%i���4n��sssA�\�K	,�,�b�˩�aB�9�l-���Bpw!���8r2kG��M���wf�vf?0g/{23#3��d��溸z�������%5=�Q���
mfm��{G�W1��� f@��3;ð����%^��+�^l%���n��aM�	HfBg�;�3b�K0���I�ٰ3Xwt.H��Z=�Ÿ�{8�^�[+�3��!6j��R�	����ƚB��;�{۾4O<A�#�rt��`�� �ǋd)�tQpv���m
A��4��C=��H�<׾\��zd��Y��a�m�Vu�[�gYf�����8զ���\�S�k�x_;WH_3�ʅ�I��-\�MU�X2�r$-�t���*|sA>d�y�7$�	!>t�&��F�L'u�ӞA��Y|��yt#��˵�2�v�}�+�1�jg��Z'-�=���v�
P�*v��#5����꜇�K1y�ѻo$se�Q	�A�
�������]����v!=O)=3�`б>^ PC�����j7���Ż��z,x�t��];�������^��>7ǅ�3��M�J����{vK�:�Γy��;��з]�N�,"���q���C���:g�6�~)#��Q��q��}���_� �H�b>���;N���������%�&�Bo���xj������8t0K�Эb�F�z͞�6��35�CI�e�e���zr�/$ �xV�w����F�a�=}��{�&����˾�k��8��j�}���l�����^�@�t`��B���gi[���imŹ���ORm�y��tG�OJ)>����ش �Rİ�:����X�sT�C��D_j͐����Kuna���)���{a���&��X�&��c�wos y�����=޼=�_<��܁H
�L
I)��j9͸뭋\��m���m�Y5�b-�� M���k���m%�(��8TF����XƊ�ۘ��ѹsV6Mnnk��E�\�ђ�b,[r���\�ʹmm���wR�Тܮks�hܮ�6�汮h�ʹh�lm̚�˖�P�> xx�_[��:���}Y�;�֛n墄u�g��=��=����=�g#$�p�=Njh��^�bL�l�b�P��N�@wFdffefP��5������9�1�wD���Ŕg���M�P̾��zU��y�n�JD�HDLHS*qFa�İ�����K�ED�鵳��1<7�}$���!�ڹ��`���Q����
F��ֆH���`�Y��f@޽켮1��� c��/,D���=��h�[ <��wd�&z��q���ݿZm9e�����j����ɳbSS�b�	�VG���̀33�e�D�ZWY����麭�`����lƋ=ᝈP���OM����&s����I��K^���5����#����Z�K��V�e{�x+�ÜIY��or�]�������O��j�{��xe�^j́�3��ړ���S��Mc�]M��=o3({0��Z#ntOL䨄,��^Q	7E�+�)l��WWVB��])��v�qYj)V#sfĪz��C�2Ff*�tc�n�MO=�P'���'b0
�ޠ332�"E�Y���J��Nj�t�m�`���r�cE��v!�~�O�����}�=�C�<m�i�}{h���>�+V(�<ghC����K��qޭ�-����3c�����n=�3Uu�ۢSS�b�	�w�T��e�O����w�mV�E����xw@�����:;1�ٍxe��n �̿�-L�,�}������\Zb'PV^ux;�g��S���Ywu���{9�ɸ�?�<�-�r`�������I�����n����#�ZA��)��`�a�����Jd2��9�$#Ù5c��h2�5L6�0B%.���J�l�{-�Q����]
�Mx&�mE:�%�B.Ҳ���K)��H�;
��@f��1���GT��\�ft��vθ�6�����a�*��/:����˔�k�F�	.&6n:�U�la�9mYj��b�ܗXԩ�{�?o�SR&�6����M����ʺ!6.0�t
�B�JQB%DL���k^�̟?�f,�q�읩�o�+{����{P̏fG�1F
���xN�n=��S�c��Þ{�Oz���7�ݎ���^} fFf!�̜&k���깵}U��Lp��V�o��_ �f@���+.��W�ƞ��}&����ȥ�;S@� �Pؼ�:>"�h��������m�o�kh���r����{��9��ȁ+��y�M���f{/0���P4��%%DA^Q�H��6CC��r�Ya Z7Y��
eDʔ�&d$L���v5��ݚ����-x�ٍw�CZx���J����m �{�'X�MP�ZJ\U_��6�DPr����\�ou��G��)�ߕf�,x��2\`F�P�������FyN�_����j��}&�FZ��R쭩�o�+uf�n������,���Cʹ��*��g���LE��Ý݌�=��m�p�[�����]�W�j*�Z+04�[�@�砨��6�O��m�6�n.���=}�Aȍ��kc/z���V��7����۠�"�_V,�0WϤ�j-��AR�b註kֺ��.uXD	J5��YK$)QBR�U`�����u5�q7t�=�%pp['�S�}�������U��ܡ�S�78U�Uk���3���e��9��%�bN�:f�j��nU��m�����v�Ԥ�N�\��5�m���;�1~���'`��E+�~x��R��G�o&�=U���T�d4%J�
ϼ<=�f������Oe��	z�ly���MǷv$n��X�*]��m�Um�G�a�n��븺[z����q���m���1Ptι��Xo�쪬�K�����g�W �鷊�:r��f�>|	�ED+�1U�hPMt���.�ʵ�P����(�l"iE�$B%L
5	��ש��n=�s)dgaꖻ.�h�/��lV�=��h6���m�62�_�������*���Ụ�s۰r�w�ƛqQ���>�������6כwSc6+��n�{r09��{��P{��Ǜi��.����A?z��A��9�Xs��K]�[4���f��f��u0�	�s�qGr���3��������1��F����󬰣�iq3[�7�w"�y�[f���ќ���f�1� =�֪�ٺ�p�m�sK:.��뻈a��.Wn����pƀm���;��̰n/���H#	���Yr�=��E6�vٖ$-À�P�r����۬��������m��U��Q[�09[,������P��^v�Y���m߃q�1�R�3�j�b��5�;T��t��_;��̀��k�����%�P/5 �^n �ٌ���Vˍ{t�r�v@5�˶�6כ�6�WV�����n6�mEު�f�Gf�Ƌ=7˓�9�5tRYBr=ۨ�n<�M�P�7�1s5G�@rͱ�R�fRu�N��l<m�0����\*�Wh��b�6�K'�	���şf���{�f����^�"�ܹ?9dm;껳$�ٺ*s:EZR-	i����蛔��|�r:���gks5�,�Ÿ���h�y͚řfI��8���ܦ��1n�*�l�B�%-v3Q��i��+	R���LD�P�6/i�Դ�����V���ZTm�#5+���K�Kv��������2��3^�����f�:��9��^3�T��h���0!5nH�h��f4-�T�	X�:1��W�<�%��3C;8�p���V�7{���.?�	x��4&�:X��+�U���5�WCV�\�\�P"d�|<��5�u�ښ�7Ƚ�g%v�9 �	��m����ӗ�� �6׃mf�Us�a�*HjbU跨�ڼ	֎�-�{��޶�u�z+2v!}�p��C͚5F�%�r��{N�fD�#}/P����m7�0K�Vs�"#�;��m	��|N�rWn�� ˋ77+ �0��ᶼ�A�m���7\��ebn'-�u��Kc�o�������{V����W�[P(��C���i�`�bm��tv���4�m%A�J&j�N����^oD�)�|2sh���6:3F��9sz0@ڛi�m��}�ޝ��g�]F������F��0�$�j,wD���FI�UK�-�߷Ӑ%��ۓ<8G����V�\��3��:̊#Xr�����} }ڦ����&Wn���q�m6ғ[t�/3��-�;�T�� ���n��a�imn�^n�óKc����ޯ7����т��8�}j;ٙ�����'1Vᓓð��	��8��of�:�^���ʹ�M�u]���+��S�W!��݂p�w�ǃƛk���ܒF��{#:�"�AE%�R�(�M2݈�����e�4���e�[-̰6ߛ��=g���������Gf��=�F�L�j!W��/c��M�<�y��ܻ�"6�N�^�4NeI��gq���}�z����Td�	���%nCz��M�m�:f.�f#�b@����Tr9v@�j��,tF�fXu��D7�0�4�vE�ZO��>��_��P�D�Ն-^���q3I�� �Fv��1۰N���4hᶽ��,�n���6ׁ�wW���7���
�.�-5B��tfĮ��1^͇��hy��m��WQr�\�b� *��Rw.8,�9[B넽^�kn�p��˻[�9@}3	$�L� ��M3�x�%Sk
��^΅�%�M�V4�ur��6����gr��5�q�5��S� �\]��{rmO]�����&ᶃmۿt��s8��5uz�9�<�N�We�7���5�nz��munEU��]��<5���q��zv��6'�����"kf�:^�fǆ6�h7��Lc�J�N�݀hMm�p�z2&c��\6b(�*8ۯ���b�R�6?Q�L�\�x��ۄ�e��(Ÿ��nh�3s'�ٸ�����J���6]�������O��	U�>���9������q��u6�Y��(FXe���u�َfw��]roW��<���
5(����\�D��0�ƭv6�:#u��D͖�&�73q���:�{w[w��Ä۠���f�E�q�,]A��x�m�^�������S��uW;�t�S]75=
c���m�}M
�At�܏e��c;�wv�����Z�n�g yI��er��3;�\p��ަ������^�U��n���r�]`���f�E�/��.`�c��S�w �y���k��q�\�v]��8z2�i2*;�� ����eoM1�r��C�}�� n�.��P#/ȨՃ{�*=�L�M̓�v�2h����������o�Oy�3o�8�K{ݒ x/k�<�l�3I%��WU|qw�M�{ŗ��_n��Woo?����8���ˆP"!b���;}�f�Ş�'���c��h���QM�wF���ҥ�zmG�����O}�m�?����菅�a����X���SE��i��N�YW���M8��$Z�ȏ�P��}�LC��O_�y���3�O(�O�b�E��be�$^��e�Cv fTC�yv75f�.�UP)��AӤHJ����b���]c��Vh�P=uS�Oz4����Mr����{m��>�\Z���}�,xCS,����N�q����f���[��!\���ų*bL���2(%Z �o�{�>�rgd^��3�dV�ЌL���ܜ�X����2Z���a3����e����x;dZ�
� K��fOu�O��;�1������h��tkRtTAOj*�kX/#=��<:��}<�r��Ǵr����ϧ\E��j.�Su��or���7�������ٳ���C�u�������NA�{6�y�톼�g��8������.j�n��yL��5��՛�k�zz=�!����zx��<6w^Zt�h9��Z�?O\���o��W��U���kJ�Sw_��/g���z=22j��f�7D+���
#�6'pX�JŨ�h�r��74kwur�wX�Q��s��ȷs�wusk����BV3���E\���sl[�TA���ث��r�wv���-.r�wgv3��ʎ��4W-\�+.��nk���r.WCmʸN�I�nwv��дU�u˝��U;����sc�����Fю�']d��\�
t�Ȯ��r�\�7wE�5ҷ*�夎�sEʈ��W#\����)$�y���������M�mB榴�c�J��Մ�.���.�$J]�yO'�K��@�0�Vl��L�k0ʷS&JBl���1Ѕ-�aF���MI��2�gd��n)�E,�G[Sb/ѩ�Hm�;XB�Z��V���pitY���]VkR���9�11��o<�V�\��i��.*isX��Uؕ��u�B�[�.rUX�� �nC���L��˝BfZe&ʺ��uص�[��{<��#[-��%y)��Ka�K�1���:b7-q�v��K.X�@Яb$J�^`f�m�H�M\̍�:V�A��Jk����Ĺ4l���j��J1���eG��k.�1k!l��E�24,F)Zg8-��n�8JXy|�,���\�����m�.F�-�1���	aXcg V\�7Lh��������SK�!�Y[lCe]��1�b��w Ю����l[1�\�[,$�n$�र,l��i
�툽f��ˎ ��Ѱ��i
&Il�`cV��f��3W��#a�6�V(��7U�Gl�&%�븍����DHp���G�slPE�bk�cZ�(�e��hҪim���gR7e	1r�����ғ)5�0a�e �������Y�BQ#�9��$r���m .r�k�h^�UKYH]��P��ʘ+��3���XLf�0F�1	�es��5��]�$Y{L�M�C�TDlnf�)-��"��6��ekv��%��v%�F�b6[�f�d+ٚ���D���nn�+WD͢�ku�e�rhV��@�h�ɐ,�R�,IR���#�2�[-��ª�Ļ�� ���6�v0�l�:�r�Mm�@��&��%�]��(.�oX��w0K]oW��."����!6�r�p`��a��4�ChKt\J��!EF!-Nn��5���Z���6��#\-�6:�l����n��|̵.:�3��n3̶nf۬�]
D�F�UIk5V����Z%�%e�c�U�k�6ۃ�p�������;���W��%��.��/�<<<4͸��JA�/Z�c.�^ĺajVf�sk�
D(h@�@��-p�e��<�V�Sd���.dY��6M*$�`&�*!l�n�(F�a�s+�"�1&���RS�����h�GJ@W�����mͱaP#��v�1�F�ɕĳ&A4�-رk�陭Ke¸���3j�S]3T.��[���,��2������6r��uj)1Yu����S9�,�2���U6`ͦL�W�:�zۦ��.�3��������q	���o0+Z��6�m�\�������iuݠ7�M�ج�+o��l�Gz_/f�x�Lg��ٔ���m��͹y�6�"�yN/�N�]��)�#FJ����m ���o
�;ׄʞSp9��f���#�m�s3�*�ּ����K�����݆����i��2���G��2���:=}^ț�\�l6��m�a��_M�	�3Lu�f�6����13 :!R�5���H���[K2\g�N�7���mJ���S�ppӣ$���ܹ�"5�r}���m�chg\�>���?]���xA��s�\V!�*4��5��-u���}�t��ǃs�~k�n��m�i���}�	r�0IuS0���3����>Yڂ����+nc�gt*���5��qs9�u۷ՒZ�l�n��}8	CG"��j���dM����m��q�.&0��w99�ٱ�ڕ]g����*�n�<��ZM�+$,�k�nmx6�n<v��]M_JnF��-�Q���U�/z��6����&�-��^IT�	+a�05�����s�EۂnW&�֛KQ�1�,�$fX�Q<�������f�H�Ʉ�u�["s�;�e�j'���Q��ʹpm���F�0��M��͡*��Ao����n�
{��ƛo"ƶ88����{�ׅ� �6��򍦥�ne�ʩo �e�	�d<}��;ݡ��aGzD����5td��q�-�qY�qpNMuut^86,�yTn��.t�,�ݜË67o!1N�9��
���/����m����Ţ0�]&�T�z���"�$����Ul�Ξ�\�ģ*��gr��m�6�n�Q��$�㴦uUh�<�Q�#tZ3����A��[Ù�O����)"K�ڗM�f��%U��al$ �jS
�b����T���[^��@6ע�.��ɭ�]�wB���.�'�0E�Wb{�ݷkN\���6�r��+�H��	t���P������c��T<�]��|�h7�QÁxL�
�yZ"�*�Wx:���y�m�8�ٌQWS�
��k�m�n���`�i�Ю;�Z��:�{���eB�B��P=��6O4�zP?ms.��p�=y�������w��E$9�"i�W{qf�<��E���ݼ��^nm�fu��q}{|3hH��
�=|!V�/�/��cʹov/ou�����vљ��CK���J�m��e�d)LGL��2&R�b`���� 3�d�[^^�Uà�����&��u�xl��j�T��������/6����&ow=����F�aಶv�zS��r��[��qw^��6&�3K���A�݄-�"s>!�-��r�t0?R�{�jcoD*��@�A2�I5y��mO�n;J�y���6�	66��Mh�vwI뤄��&�.�<���:=��ΟO�Ƃ-�����h [�R4�U0gQ�
��YZ"�JzS� |r����p�Ǭy���,�u��P.�
76��n-M!&����&�=;XȖL|�(�:���a˪�c��BN"a@������zڔ��J31&$ d�	����C.V���� �%%��V�&��R��[��@�b�*��֨�n�{)G1��`C[�l6� �[b�.�1���X^*.�#����.��t���"2�b�a�UL�5���q"J �p�#Jb�\�cr���M��JA�cE5e�&�p��u��t���%ƅ�f�ۚ��.	�m�.���=�B��d�Ȏ)����Z����G!H��@˩f]rGX9&�8�Cŋa�nlF�X�O���q���#��۹�m}u�3(�W�!V�Q �����j&1i݈ �	m� �p-ǐ V��@��M<챸��x��A�^T��r;;��ԡ,l��C������ȝ�u۽>"yT}zԀAmq��G�`P騬!�*�ƅl�V527��q��h s!�Ȍć����pg����1�#��O�h+�1�D�7��&�3P/��hY=�8/�㵍;��A/�y��Ÿ� ��>n�=��S��ʄ�yS�j=;���I�6D�t��D׃mz�^�~M���ǫ9�J�Z%$�8����k�+(itЂqK�sZs1V�U%����� � �n͵1wY�[5F�-�=�jڨ��Gc�wG��0Cnd�x�ٸpu%����S����Dv<.+�{˻y��F丑&�O�B~�����2s��ozG��(�_�ľ{��c�sۃ���3��'?������̣�U�p�G\T>���3PE�K��5�2�����uǗ�-�[�-�6v���D�������52ơUHqw�q�mȟA��1��
ʹ����m��lA-�"*��慢�vl'�q�k#Ȏ��D�ؾ���1�"s ��/[^@ہ<[.�e�RfvX��.�g
B����_)�-�D[k��FL�f��ʄFL	�J��ݍ�9R�"j2�f�1�З�J�0l�G����cW A�D۳�����T֎���Oz�K��t�eo�\�j"�iyx�͙�mp-� ��G��Fқn��  {5����S{	��;�g#Ȃ�ȟ��F�k���:��#q̂{�myۑ>!�1�+�s��K�u	�s���g)����M׹1�Mm��7��U(]���U�븭��J�Ӓ�<�zP��C�_��+�2����G�9WQ;=}�q�����}z��˃�E�c���̻+y4�hr��"Nt Cq�&��r;[������]WH%�/�O�!QOc�v�O��-�Ŷ����7p�|��j}qtፓZ;r��G�G����p���x޲T�dB�/T�1[(�+67V&x��nM]���ds[QV.Г%(NwH>4�G5�CngŴ��l^\��M���� �\z��I�<�F���A��݀�-ǐ#6Y��P��KGy��!	��wr#�t��B�|��#!��m���ӻ��������If�>;ܤ�Ygȶ�nD][AV��,�g8d���jl0��\x �ϛ�_�^D<s!��̛�� �� E�L��
����u	�{�)
ܩ��=�@>��=�fk�3�ܥ�ỗ�*f�cnL_v�ճ�.�"Od4��{x�Ţ��y����i���W�|W�n��^�6{�f��.��e^��xOg)7��k���j'0�VEK��֎���Wz�K��!��"�/ۙ�p8����6�>]U��!�4�f�����wWR�pQ�ט���0�ED��j�x��^�v��p��U���&�y�8�!Ql9�X�mTzH"�Ȑsa�ys ��.��T�*�s�Ȏ���
��W�&�pTk]L�y��nҳ�Cb�H�J�+R�ly[r$�my�0���]z�7���M�cP���AwXב�������,o=VE�mA��})�; /q��Q5
���5���q�Îeǅ"-�*�zg���弼w���ח�m�]�]W-�� ���Y�&6o���S� �5��YeKmb"5lI�o�<�!�����塚�D������r��̸�C6�p�tE�{��)���l�Í�๑`��ʬ�n(e+ӎ����2� �%%��W�TY�q.�ܕ��e��U�L˪!u�]�s�Ve&^t����I-L˖��&B�����)�"��Kĸlu,�#��S:�ά��8bn���4�P�r[[`صv��f�V�]��h[{Z�:�A���$���f�;,o.�
��Kmx"��cg�YmcU�����ljj��B,a�V�B��j���!Z�vw��~���ʎs0�1k��q��H��K.@�dښ9�,�P4~��6B ����y8d!U\/����
.�<�~�d��,E�>�=|������ �ڒ"%��mor�l�@�^r�6���x��q� MB=���/RGQ�i�r$�^ ��!�^�дy�5���!�E�4�TGM���Z�����R9�/Y^ ��RCh o��<v��I�xx� �y"N� !�"�tu�oK\��b���	w���^��7I�xFW��>�e���יd����0��::M��T0�x�d��D20�/�i��%D!@ �ݒ��X c����!X�͋Fj��2�͕l������A�AB6�|�	��W�Pv�͙�fO6v`��k�
85�~ � ���Am�!���q؎'掉�b�Ww�Q��M~�$�SL՜�����Lq�.�m;z*:2���+�N`��U�vC��B�d�Kf$��7��#��[g��{�)��6�]t����5�m�V�����!�?t��T ����,�� ��F��r�\a����0�a����p�!�@mؑ�ڑY/�̊�� �2�"|ChU_P��Uo����vd� �<���9�V�\O'xc���G߾�&eq,Fff��.�n ���!e�]��q��M*clL�H ��!��D6�|[AI�������|�_��lW4tVK�GGgņ�%]PX2RݹЮ��Z;s\���߶[���~��,��>m��j���7-���C9�����T�4F�}O$I{�!�^n/�ǃ���]���#�����h*��Yd�����̞��H ���Y��X�D.�پ�I�5�	�� Cm	�@�2�4HG�pv�sx'\�+:׹w����N��n4�Vw�~��o��{fi}3��>����-kHu7=��\��.zx;�:�S�6g����o�MVzy,N�yr*ڢ�n��9��A�,t���;�w�F4"%^��ͩ獓lteD>�~�I�&����_�^M[��ؑ�F'n+��/g8�+[���^t��$���r/S��^�X�#�_���||z�:�8����"�Pl*�1�ά��l\��ܽ��Z��~>u���wԴ��wz��;�F(ڒ�T�֣nT9SBEj6��
O)�y��//{Q~de�^Ų�=��=qx�#Y�	뙕D�by�e5
|��AyM�`�7���uվ%j�T+��&M��x�	]5b�ؗ���|�`[���^\&��M:��Z�S��8
��(:�bw�Z^��wdkgnL���W(1�vFn=��U��o  N]��W�V^nXF�R��e�Kwr;�����o�n�M=�^����N�c�.�Jۭ�0��C�+�B}��u�v�n�!�c����.���3��r��y$�Wٞ�Kh��I�q	Ksq�2�H׀�8�Z)�x�6��k���#��,�g_S��7�6|��o}�;��콕�[��6G�.��̓��}ヹLzM����	���%94'f��"X�*���=�{<*�;;�8�{;-Ω�����{+��0<��3�	��L�F� �)k�gjƓr���VB��gIYkFZ9{�K\Eڔ����nkwo0|ߚ��=/�=��rT�B�XRRE��Z�sr���r (����c���9�:];�Wn�˸���n�us�`�M��v��"Ɖ5BkF�����Us����6�,�̲Q���Mn�]u�\�s�X��r�ō;��slm˗.Z*����sr�mst79�I�M��#&�F@��J
�Rb�����ruɁ��A`ԉ��b,��)���r����CF7D恔����0�hLU�n�2I�4�5�ݻ�h������Pi$�t�\�I� � S��ɽ:�4�ؙ�	w�����יg�F�T�5Z��F���A �ԅF����7=�aƤÎ�@�GD,�W�&:�Wb�z4;ʰG�Ĵ���U���bfg!c��]X[֭#U�������.��𹭅�̞�ؽ9� Yex�[h�o�3���~���߳�8�Ѝk����P��;53��CM
P�5��)3��K�����O��@k��q�p�^��}��:4��S|$c�����=WB ���p,�� ڐFƑ��Q�@8P>תDѹ�:6n:�K��Ldr���"|[�)��A"Hݹ簁�m�Hm��uYY��Q#.糌�.ˋவ-vd��RA�AY���^�7z;;�<H��2D�eϻb�8d/Vپ�q���U�lL�	p�Գ������Vh�:��yw�ɛ�6�3$��0#�E�ǒ8�tƛ�l���岿Gȗ���wI��7���f?;Iy�7#H������Y@�[jA�e��(K7�(��Z�:6o��ri�* p4p�/vD��x�p��Y������ �=� �w5�B��;iF�]��,D�R�:�6�F�jͶE�VU����&� �2��m
����=gc���K]�<F�8���?}|�/�my�@��y��r:�唐��Ds�WY��oN���J�n	���@��y`8���m%�ɤ�8����� "�S6�TY����S��z\���Y�LLp@�Y^#wP��y6��m̌��b�9e�؅�������*����=gc���K]��ؤ��f�˙� ��D�Rm Kq�A�[��w&�o0�=uf���iV��\��Dב����6'\���]���.��]�
t������V�ѐ0��'W���=Sͺ�]�R���縬��΃bF��f�fÉ�6޸G����=����"��Xm��
�]4ݭF� &m��$�FĤ���^�쉥*�z�39�в��c5 qb�<�]u���Ɔwd�@��ҵ/l�]k/V��1jT�c�EF����u,(���pQb�ixu�s�..pX�Q��"�e$:��CS%���,�a��
�@�(�k�M
s�,K�V�Ά9�u�܆�ut9-I�SkJ��L#���k�]W���N��Ѹ�Jua��i��@�c��)hQ�ڵ�1gj(�.���}��g���2=����|�F��梶z�t���bc�rS�Z~k�E0�~C�X�㹃r� �܉�B���b�CNl���"^/c�~��ɋ΋����-k q�r�A�A�(YǞ?u5��@��͹p�ͯ%�wN�*�n�qY�d��Qڊ��2����"�"r��Ax�ҔI�1{yM�J�c�X�{KmHf곑[=Y�ٽ�bc� �Ǒ�:B�*�v9u����m̂[��� Cl�YQC-���a��к��5}.����;�u�A�n��m;U�m��z�!�[�r�͇I�e��@��PcT�%ط]V�,e�qt��&	�$�=��^ ��[�7��7�:йlY�c*�F��Us�8F�\0A�^Dol�>-�7�A ��i��:5�C.ЭUΓ�1��|E�˥3�{v)��A����8&2�l����>�[
A�;��zM�y��m:�l�GUm�����s�[C�8��syH�7U�������c8�ǐ �Ȑpêy7�L{����@���!�3����w�,����x2s��Ѱ]��ד���I���Q�my�fJ�����O"$l+�iW9�tY��+l��(cf;L�F��\$�!P��fv��N������>ހ�-�Dmz[^n��S:jm�{�U]Wr+��8#���(� A��"nȒ�"�k'?.�凲�O�����`�:�pR�`�ո�mU�X�v�s�䁁ܳ�?3?/��ϧ2�}�o6��H�����.�ikɁ�![.��D(ԟ�"�^�^>m���	n<�D�X�wag��=Ѐ ���W�����n���UސAwF5�mٕ�Rt���
���Q���k���A-��g� �����uqUs�)��E['K�� �ó�l)z������֗�j6v�:k�XI�A�4-�v��Ƭ��m��j#w'Q�j��sv|�X!��!�2$!x9ڢ�e(����gj��Sr6��:����n���>9\��<�]��;Ӱ�)6���ynD�� ��U��/#ˬ��j�(�h`�U�O�� ��yۙ���eT�F�F%�L�a\�J2((WQ��	�f��%�b�4�l�۫
e-��r���B-@`�v����Am�F곂[+���ܜaG!W��W$�y��7�$�B!����	n"Vh�4��ŗ� Ï"+�z{��AnWNR�<m�ד��S�A�jŖo�T���j���ZFb���!mȒ�yy�#�e�����Cm�l�A�C�ʤ8��!�������,���f1e'��X�����:t�KmH�7U����̭;��(�����U-���HdVD�I��y��)ɭͤ# ОgK�=�ׂ�[G���)��O{F�k4a2�1;��;Mb�5:�؅Q���CjfZ�8p� �q���%�@����rj��WR�����r'6�].�����g��RFl��>^-��&��>���2��`Ʉ&dB��D[�Jh�s����b�p��p�u�җ?���nO��!�ȟ�"�2*�O\vN�40m����7xp�B^9�7Y�������������	��#�W\�l��Zw+Q�h�svD��=�o(�$Dzݴ$�� �z����B�t���ZαO��t�g]�<A.�O��e�|�RCh!ٵ�]U��J�*�h ��gϢϛ����]��u �Y��leWH>.����a���#�dO��/� A-������B���4�h���f:e�8�bs�� yx���$�Kp2�)j��tRyw���]�2�DOV��ͼ�[+^�Dk��n�|E��\�Q��ny������+�{�瞉����������a�~�9�f�!�I8��
�v�EJ�W6�֐��D�\�J���66�`���&�YcT��ط����b[���:�bV�Ռ-��X:��yf*��^،�%��]��v��0-�`�P2�	P�	6���u�u,&-QsG,� �E�y�u%m��\B�ס1K JFB�)���c�-0�قUR��؉Q�
�	q�a����ev<�_m>��Yj�)5������&�I�:�fgf�)i�6�j6V�g�=~�� }�6�|�7"w9�T���7FLw�	Tdj� ����)��xKmH!���".OF]\�ͥ�Π�8�
�V��:�Rg��6��!�� '�l��Е}���S@UEKz��n�P$1D�VD,�0Ծ��t�c��̀�:�D�����@�����w]����@@��^��UH��su:#��ݭѓ|딟>�Z֮cH����Cin���4�Q�9B��ӝm`����L�C�ʮ�� ������{~Ғ񿥮�f� ҁCt�#四�m���Y�^�.aB�K���X�L�͎�Qar�<�{�>���#�Cp�A-�1WZΥ=��Θx�D�ESx/A�Y��	���[��m̂[�F
uvc��L��ݶap~�����'-p�AE��t;}?~ܼ�_ϔGU����듾;䙪�>fmM(r���{�����ꁀ��"|}�*�O_9��Q�^խѓ���栈n2��Bos��;�Ұ�p� �܉-ǐ-����KTh���2��:�=dP��'+��� ��@ۑ>!�qDpð3;�=��#��<hKmO�U��3������� p�i\��A@�^�B�n��cH^!�3��@�6nk��]4/ݔ��ԉ�{9�Q5����D���pe�A-��r6=|������o�f�-�g]��X7n�'��6�]P4+I��3���V�@��g���O>�n,|�U�h^��L��cМ��,}ʼ��M����5�sw̽���^�o�d���Sq;�6&{�kjlDw� ��׳���N��H��7�B#��A9Ё� 6�|[Bv��!L��y�މL4^8���� ��pfkM�Zg4_R�;ga�u#D��i;{������@^9O�wSƴ�y�<'$}���ot��g�=��{�h�}/��Y^ ��Rm {*��=KZ��\�iD0A�nD�q�ᐽU�lf������9Hp.�"�Ed�s�U�O�#+g�㺂�|�mO�n,�¢�ZD+y���ve�]���\5��";��@��dIn<�;���/�&m���;����\���a��u-,����(((Pd�3���<����ުf� Cn|'���AOgNj5�a���ڀ!�.�xЊ�i�J��^n|mI�	n<�ya�D�����A�k�
��c3v�3�.�9] ���c�P6�:�iU�q�4��	��$��  [j78Wm׹el�\nѼN�\5��"8 N�xk�,� A� Cn@�e\k�.��F�4F��f��m*�WsY�k�í�ݵ���C��/�hS��5���y���Տ�g�����7khA��2�ù�^m�cU�{�c�'q��T�����\\v3e�Ro �Rm	n<�-�p��ˀr�^@7�lf=�r8e���'+�$]�� �^@�܁>-�u<=�+|g�y�	tqrB��3\Z�]ZP͌b\R���(�K�F����[r���O�����`_�p�Ŷ�*�y���y���6�G/C�3�����q�r^�6��mȐAn��F,�Ӟ~!�O��n��Q���G�f�[z�G��^���rN��<���u�kH{�Ȃۑ ��#w�F*;-�̙��b0m��A.���b|���+�a��%W���@�/P^:x�KmLU��/�s��Ʊ-����:p��8N[Uc ���P�mǐ����An�6�H�fх��	�Vj�;'Q���޻(����$7 YeKm`utm�+�r&������[�v�m
��p*$Z�`��T�k��a�ܐ�Ue��cR㊤�di�CW�~���$����l�w�k�n��a�d囨�1��;@�l��_v�7�s_�e*C&;�6ж�G����v�oz�=h��iT`�ͣ5�[���`Պ䜽��xI�.�*��y\]¸�g�,����*=܀$��i���42}��#ß��v�!Z1����o��<�(o@�ud���<�@��}�'[b�Z�{���(LD��S#R%���e���C��hA�2+���*y��w,�����?]`�Wnz����)���y�D9#6w�yq��tþL����}�$�;�ˉ����=�٤ļ �8�!M�ŠW�#��H���W-4�u�͔jco���u�7��]O{�yN����٫��{��mA����+P���\T߫	\-P��"�.6�j�_.i�����*�8�.Y������n�n7��ղ��ʺ����f��ݍ˭,f��aE0���s�k^kx&��Cr�B����t�l�c�*�2�!�3�J���P��t�g�^�bf�����˸�����)�CU�^an�ꇆ�夳s6̢���D��� aư�:*"�f�FwJ�j݌��m�����"ɵW��F��T�77jq��t���cq&�O,Ryi`���JܨX׫CH����4"��U^�����q�
�c���O��d��?xe ᷹E�ż��l����Ĺ(a�����卤s����;���Q)ǜ=��=��v�"�YT�㷺aΜ6�\�9u>�; 64e�nwn�s�˦4E�99�+�]uq���1k���pƓC9�G;)���c����"κ7,f�P;��HF5ͺWw&�TF���ؒ����ܹ��0$�	����d�Ѣ�e˒b��RcD i���Ы��Lh4A�E��,��vۑ�9]��!��W"wvE�;F,r����'w1QF�Q
i��F)�u�$�0L.]0�`CX����C
�A��"�s��[��Q�aJJ"	3�-29Ý�dDGwL&!�.s@!��Ź\��I�a]�b�C"�&e�8�V@4����n���wq&Q ��M0H��.���ՙ���m�Tj9� �\f��m۴2ECa�*m�q٩��ۈ���M�qN҆lo�,LUք.Ҙ4qJ9��� �v%����L�����nVL�`���9v]e��%r�a�u]F��V4�pM)rT�V
�7��&�i��f����ѪD��#����0qG���6���ש�ZB%�f�C�'`*�ݮ�8ĥ�,3�6h�6cQ!@�vF*D��p�J1s*dk�t�؍��(�2平4���1��M�%�f�ؔY���h�b�t�)5�u��WHD͕flYJ��ь%1��c5��ц6dՍ�XFk��ƀt��Ri�vtc0�R֑f�%�1��%5�(�4�;�\�c5��NNL2�lZ0�eԥYD�h��5lf��Ib�X�s��Z���V6Y���f�Kf2�+��]ku���K���K8ˑ����%%�Ih�i��KiB�Y��c�E��$�Ц5�sv)u��5����25����-��RCm"a�)i�K6q0V�i.�G�D�]�R\���-��nP���%<�isr�U͍����c��ޔ9-������i�M�a�B�҅٘�!��XhJmz�X�����1[j&����i4m���L"���x�t�+�۩#��g)I�k���]�Lƙ��\��H�4u�ٳ�cVJ8���Jgh8Rk:�66�+�*	.�D�%�#�z�n�[p*U(]�.ZE��Ek2דZ��=�T�`�����R[M�FjJB�qHui��xB�Ņ�WMƚ�t�145%��ʹa�
���A�ĥ�0p��@ml�ZJmAVYf̭&�i��xe���]�.з]b�hucW[�4��F-�d̶��	��Z�D�J�M
)5�Ҍwe�]c.�V�t�����Wv� ��vN�A�Ж�Г65�e,�ں0]l�rGcD͔f5%�DH��6��Vm���S51��q�Wr6x�I��i�3]]B�k��v���d��kݹ���l�f�W8��,Y�"Y��a�*4I�6�tl�-�E"��]+�f�Z�v*,U3���+�֬׬��)��˨���SC&�SZBE�c�Ѵ:4*j��%(ı�ci��J�O>BQ.��!�-͵mm°��Uᕤ�ld3�M�X]F�Ќ�A؍��K�y��%�-��)����K�Nf�q n�L]a������F{����l���[��uŮ[3��b�c�ֱ��(�������G|�O�Yu���������6�U�l^n�T8e����	��'�YUux� ��!76}> 6�,�� �Ԑ���[��#��P�F����*�u��9Րֱ-����:p�>y�$��;R�"��m�!�&�� �Ј!�!ۙ�mɵ���]��y���b��ҭ�fOK�> �����G3/Bf]�V����mo[�I��N�H�@���*�����j��6��C�]� �qs�Nѫ�zG�s>#y,�-�$^e��R�8٨6t�@&w�tN�{ӝYk���!͑>-���"{9�;�	e�,!� j��3F�X:�L;b���8ԬMˌh�T؏����ߟF��Oll��f||�
&b�s�w�/K���vd�doGLjy�"Z�Aւ�(	m�6�%�B[�[;����"Бy��0��At�f���}t�=�bHk�w���kyn�U��s���-�����@���M@��2��p��8��T��l2*�����j����u��w}��D6̉8�ˍ�`�Af���O���P ���'X<���;��E����Z×�G N�!x��g���� 6��ǶUdf[�r<����؟�B&i^�do�S5���f�!ނ2��}����N6���Ŗ@A�>n.Ԍ���q�3.�_u��C���u�A.�C 6�|[C
�nO���~�p�x�V�C
GB�q^���؉Hֳ��3DH�Z3U�Ȕ���9�����$>y�I�Ye	m��U�m��YՍ-a�����oADaŞ��(�A�"An� 6�H%�@�E]T1�H����F�τ���!4�s�;��驚�vd� ��RA�2��мiOV���(�S�GZ,�-��qd2�"���أ�G���t�b���Z�Ԍ�ɼR[�_?3��}2�����9���H�����d>3�W�nzє�6Ik�I�/��C�� 3/���^�n{:ehZ��K�Dad CnD���E�}9���j�75h �h t��|�R"�3l�ugV4��/�@���!ڬ��>���kaFF�������!x������,�_���dӜǑ�'w(��׆O�^���� �mWv��r��~-�Թ��&�f[F�D+�r�3vBޮ&��2�fT�]*�c�ܚ��4'�t|[�A[�F/��g�`[B�t���Ԍ��1@�<B�ܼ�,��'RGNSP�Dm���G}}�b�5�>�Φ���
8 Aӄ�>n*lb9�uC�!Rl�w��u�ᐈmȟ��-TEf)��y��Y�7D�:34�p��@3��Ch"�(KmO�m1Z*�r�D����C�Ǧ���^���%����]p�;��;cw���"P��`�U��(AȪ/���(��]rve(}:C�Ќe�Q�EnX.���1f�:"��RB�kN>�hΫY>����j&r��.">�^�3.f@����J�΢�H`�jDV�u���m-a˰���G�{"Kp�Amz���V]:�7x����O��z%@��B�&n-e�j�ذ���cfI]k#(<����`|�t �9yx�܁>-��g�s���;{Ff��L�dѫɨ��{�h"� �ڟ�q��4Z��v�|1�!5�vc;o2z3�mU�A.�F5�ClQ����{�/7�;x�RCp-�@���OnW�9�=1w���+�kt:vp�� �{"An<�^^6��/qv�u�x�݁���ȍngŴ���`��.���=�2x�v�O�C�]�9��s�8�
:l�	��Hm/2�@�ۑ%���%J�`0�_B!Ovݘ�뵜�`[B2��]�� �!��m�Kht^Oi�9���4�"(e��5M\��#U�v�KEd�S�j�=���]ӮhT�P��dD���ˎ���Èw����Kg��߽�y̨@�� 8�gY4-��8ؤ�0�i�U�1B�5k�U��v�NE��!٨�:f׈6�И)��V��pf�Wqב&ؕ4K��v����!k��T�@3-���L���m���l*�6d�(`2g����.M6�%�\�u��8��s`:��J���m(X��3���+��ו�	rF͊��	 �9�)Y��߳�}�n�1��Sl*�B�]6.h�7�2еĦ3�5-ɋ��T�u������|�[�� �ڑ|����n'tl�
 T̽�����n�MǸ}���`k�ۑ ���c53�	E_�.�O�4�T�`��5�F*��>�v�IZ�,􉽝ډ�����R�^^��܉�@�"VD��t�k5�:3�Κ`;C��D�B6�O�h"�(B`�فв��޺�*@ ��<P �[jb�S���wt˱1�@��D��s���� �d Cnd[�Ap���.����&D�\�c_I��1T�p��;�H:�^,���m^�Q��ʘ��C%�PY�0��6��Zj�u��*���m,h�2�T6���aP�F"��&N�;uy�`�Y
jw�/6�uHk��krK�؈����8�E�L��ŖQwv��.����F`�N����h�."��"v����b��r�f6�ݎ���U��Ҝ�b5#Q6Y9�D59QM����1P"/dǴ��A �r�z����n%���T@���6D��ISļ�.��H�Ȑ�����B6�O�hM�F��q�+�a���w2�p��@3���5��,�-���z,ʺ�U@zf�(7�$�^ ���7�^��Τ�v�;�p����w\F�FS�>/�@�ϗ�mH ��@���m�#��R�ǣm|��굶����Tp^�dodIn<��GrSJ��nG��9�0{<�� �Š�	$��C�h�*��#.0f��ʨ��(MSb}߾�e��"4����h(����9�Q�pf^�=�2a_Wv�N�͈�ɕ��=��(�[jHn�e����������r�4��8uYз:(���w���@�2���vro�mהG��A�jH!�e�A�m����:�����S|g0<�}��m���麭3����o����n��;]�r>ڃ�Ε�x$���������������>�"���up�i����8����Q��͐��ϛ� �ᐼCng��'F[��mН�>�d of||�J�̞c�v�Və{�d��&w�����f�wi��s���|�cRm	e���"|[��tT�T�r`g�8�7$p�áw8�@�p�Nt"C!r'�6�7'W}߼���d��؋�õ�6�Ej"g8��ͨ$JͶp���M����~�|��d!?}A�(�mH��r����l���[������"ݑ>�yy�!x���%�^" �d�W�����'�8���Y�✙�죠��;�|A��-�6!�粤X�' &܉�n8dmGfW-8l��"�<'u��8
+��^ �2��Ax��mDe�h�A��gJ� ��F��U�]�޳-�������!��z��d�� ��2�}�'߈��I�xol�Ee*�;z��T��1U��i*�'z�V�3"U;��pA��ޕ*H9���w+"Awf�7-{6=��d"r$�\2�>���w!0�^#ϵE�s�
=�	��$�e�A��^9ٿr��J�Q&J��fe�b�j������q,�ZC)����[6`Q9k���3�D��"d!U�:,f���r�6D;BMŵچՍ���HDs���/Y^ �ڟ��Yomdm�2� p����*���뚻�⡭����6D��Q��WA�(��s�}��ys>-�H�⌽jf�b���혭�:�@���) �Z�Am�6��]�Q���txvoH��yy���B�N�w%�ȇ|$�=��n�,��ς�s㜂�n���q��UvVFI$,��|w5�yW����JŶ��.���>n,h��V���y­�7e�F���*����.�����w��γO�VB%��b������NR+�k0g�	�g�ܛDL������}��6�<&�F7�D��5�l�Z�l��F�/.�3@ UJ0�ee������m*����]sLmM.�	
M�6v�����F����s�qsj*���aV�U�KnX����z��q�ζ�h h6eqL��V��i���k6�"m{E��ځ�65#x����b�h.+-�Y��K)0� ��ec-���j�XXf�i�{�B��%>�M��P����#]2�Ѓ��y)K�4����&@2J|���^ʎf�/�^�6��ՙ��C�ȭ�:�@�&y�eDpmҠA���6ԂAq��B�j�/�+'rXgr �^[Sg��l���ܗ"2��.��ͯ Cm�^��R+l��9���> ��Ÿ�[i������F*f�닫�.2�m��]G��#3�H-ǐmx6�C�W]]T�:���y���h!+j�b�}��Td����r�p�S���)[���7�Hm Kq�A�qmE�s������ػ�4/��΋�����.��y�^��������H�o���S6.,)ֶWK��u%4h�7���£`f��;R��3�L���9��s���,���"*�ȷ��7�M�[l\pB��Z���hO�p�>Ƽv$� FS�v9�}��ǉɩ�t�����OU����p0fx̾}��{3�ԙ�4j���kbbq���'p:{��S[�pc�C����Bc�����ۑ:*댁� ��RA��鋗P���k�X����<�>mȐ[��m{GF�ާ�X���l]��Ȍ��K�Dc^�����ofۇ.�H���=��r��@�mL]�{�֯��n�ب�*�w�����1{84�D��!�"A-Ǜ�Q�y��Y-y��{����nD�{L� �=�A�� A���q�8�[;Y����ډ����X(�p�:5q`KV-�ZB�E� �BaDAS��B�n�-�7[=x��^��V\�r�	vk�-w��抮[F���������
 �[j|}�������v�㯑����5�c"�m�Q�@�f�ȋ�B|[�[S7굪+a�E24k�\�'����CnD��7���a
�/�֒�XB�ދ�(��+��*wp�L�3A;��ڨL�;wT�szf�C*>���睯T{Y>�u�����7��r�9���!�|�_?���\�^�Y�e�rp��
�p��A��[#�dǐsɳYua��;��s-r��
T%��=Su��8�Z}iɯ�v2�Ɋw*����aЍO��q����<�������1���X10)ޚ�9�1mm[�<K��cz�����G�-:Pզ�n�{���՞�7q�V�ǟ{�f���٣A��m~P�1�'!����a��aLe�L�PF����)m]6I����h�v�潇��k_9���ז���>�iӄ�3���@��uA�δys~7�X���ּ8��=@rlQ���_M�C������
���ӳ�*��(S���k�fιGH��qU �����U�ŭWI������`�ݭ�rlB��lf��՗*AH���U��![;��;�2�@�&-^���^QMe�W���n��nu��g7!�fuOHr����$!�Z	`�x�f� ��Y�^��5��瞂�n\Fْ�^���ٝ}w�D�K���W�=���E���XװK�q=��t�OpGD����hL��\Gp{R���/�x�p��O�}4���'��V���oɳ5�X�=ؘ�R֍R]b��_h�j�b>�o�H����i:|�Sg��}�~�8�v�2B�|i�V�OEc/83�W��o���E�jb�J���D�wҽ-m����w����[�VТ��C
3#wt	#;��i6D#��� R37P�)�!$ʁ&����Hbc$LY��&1�)�YQ��J%ˈ�D��2�C""���.��1�.�	 wn��'.b��"
21	�.]2&	�̊4$�$0RLę&J&b���.$�9�)r�q��)M@��FdR�*u�,@��hۺ�S1��BL����$I��H	"B�;�RDw]2�2,�P&�4��HS�&����]:br�F)JHFr숐ă CdѢwq��9q�%�L�%ݷ,"3$H|A>��}wU���;�9:*�9� ��R<�E�6כ����G�G�z�>���[^^���tk4hΉ��L����p�B�$�gw�،}��v�#9n ��Rn-��6&_nn�ڞ+F ej��է�mt���ب�	���B�p�ǦfNŷ�!Q ���zK.j�fk�j���¢.6q��Gr��ir�Ӛ-�ׯ�!���=ߤП>|_7J�����.tͶN�o�.�iUV�3�5� p��-���X,�'��5���2<���!�W��ѣ:&˝2_	��FB!�[�"�\k�}��G�(������W� ��M��-���ڣZp���m�Q�zM������C,����a�Wt�q� �aw�O�m%O[2���.tn�8x�{��futr�bU]P2nFtfR�kL,���Hkt�凎�M6A>�V��G���ږ��:��<藯`j��[���̛���7?�o)!����,ヨj���E)�!�x��Y�C\�9� ����"C!r'���lAɽ���Є-��V����HGHY��8%��9����� �YpĔ�H�����'k�`X,��[jDm�gpnp��7*�ب��[�L���3�o���O�ly��hO�p���O���D�O��!*z��t{�����8x��/H��e���F��b�H"�@�,�A�>n=nz&��9����P���Zs�A��>wrۙ�m,�(��Ko�.zNu,\�J�@GOA ����&oN�GFF���b��&K!A�F��X���X���Cʱ�C37|3/=�Ӯ����ܜ_W.ҳD^�d��A=\�� �� ���؅w�"��eG��q������Q������S��rj+���zc�	�A9�O^�`�^���ʛ ������啮~�3B�Ѝ&�L�l�����M6�2Aڰ1f4t�� ��]	���۲����
 �.��H($����L��ːƀG	��i���M��WU� �a�tĥ�Lb$��.�2c?�O<ǒ.�ց�R\p�-, ��ZF2�-�MW&W�HU�ˡ-v�T�/3�&�.SjR�=s�%t�Q�GX&XB��WMWU`�α"�L�����Oa����h��Z��*�5u����e%��M����2��r��x����|&!���H-Ǔk��7}sQ��C\�9�#"�H�0B�n�\��QDk^D7����n���בۊo8_P�p����;݌���Mm1Q� L����H�[��O(��A�/�� ��^my�^�Й��ػ�*��+�t�Y�/^3��RA� � /�^n��S[� �f���]�yǓk�l��M-u�r�L���.�,����L��!�H�v�E�|mH ���	���s@�&T�71{���aɭ�*9�� �-��@�����Dg���������>ŸNf�%|pOZ8RU,���TT�i��kp�7bR���ϓ�~0>����^@��ψ����N2_.�Dfn3�;�P��1*q��x�����RCiq�GU#����	�RB�)��/J�Z�����Ep�Q72R�8*��]^K��.��#��E/}���εZbo��+�(\�y���iI�	�lp6��6��ٻ���t��r�L������8�q�i�5������|{9I���
������Ëb�#���6zYɨ�-r�\y��$�n=D6�.n
��zݻ� ����y��h/J��+�v�����@k�H#K�qoK����\A���$6����[��4�b�dEr��mmjj�Ls<r\�r�A.�Ƽ����=�W<���q5�j60ϝ��m� ���..�ԗ	i�&�u��m;+f��oT�MW�z#_e�D�Yc�E��1��1or���ee�k�s4&2��ʽ�}Q�j=> ��"A{[^@���q`��=f:�hB��}���jJڴ�;q>����9� �RA�,�2:��e����A�Kۖ>:t� 6�H-Ǚds�m��`Υ�Į��C�6携7��sXD@I��:v�͵��M���y��z�f���s�wE��d��;�pn��umh�3s�2���s��Lk:r\�r�A�"����|Ch ,�'�4�/��ukTGtp�D[j}���ܮ��c(�P8,�DZ�:+�s�B6�H%�@�Yۋ浢��&PA���F��|+Y�ͶN ��RA�5�Y���oS��ew���1.�iv�f�.h������������)���jia���_'��hq�𘇷v|�X �׵]�N�ʘ�r\�rЛ9δ�E Ak�wn|@mq��Vj�FR2/*���|o5Lvb���W�xY���-r���[���Z�WN������"}�@6��!�"|Chdf��HÆ��Y�=���k79����x�r����,��%���
�FT2g�����>=��Ap�^�wK�[����%Ι/��]�i{��`���\���[j�$jI�����U�m��y࿊��ԣ�A�6V�/�&�RI��R#p?��2�A�����֪�z����ftϋh"�(�[k��YH]�;��{�j�H�ƫ#�����;��$:��"�In�p	��gb�ܛ�ޢ0�@�& ��C8��G�&5G&#�68PԆ��e8)f,��$�@��� mߧ�͠�f��C܇\5���c"8�/ܥ�ɣ���:��^�Rn n�;����w}���g����]n&3G�:d}>w�2�@<۞�=�H#�J ��y��,�A-��a�i�cSSQ}uv���;��%�!E�O��!�B!�>�G;��M8��G�@���>m	�&��ks|59���^1���nT�7tbމ��|�W��-Ǘ�-���n�(��۽*W��M�.�n�9Nt�.�A.�5�۰'�6�������Q�g����bfK��P�8��FmJ���j��H�:'b�cV��D5�gf�=轡��� ��RR2���Vi.&b�DLPa)���%�J��%���ʦ��ٲ�L�y-�5�$�I��uرu���&�62�m�&:�f��"䂬������f^ɥV���Y��Ʃv����BD��77�[,($v�˂Wr��XЗi�i�*��b�5�D1\� Tv��[��:�:�]@L�2���e3�KF�4;Yhv�]`�V�ы�.�k��>��~	�.i-��M�L����,cZXiY, ���(�D�{p��A��Am����ûUwÆD`��s�r2n'dDdxg�܉/CkȆ܉�q�v�ṕ���3��hN�7ݙ:��l���d@kyHs��p#9\M���F���D6�In� 6���D騺U�:2�Dލ9nt�.�A� A��CngŴn�z,�]�ޗ/)P �1s� |�S�ڜ;�W|8dFI������nL(w,Un��р�������An�!��Cn�qbU{,N{r�rg<<�9�7�� q����A�#��bk�zm��K�ؔ��P�vЛd.
�5�bv0�LD��t�`씹��gx�OW��ȃ�}>n,�k�uM�tm�z8�� �AnnL�,�vr�>�j&e�G2�\̽A5�z�Z�����C�0,ꛦ'Bn�+"+O*���e���9ŗ��N* C$�􅗔�����I��5v��V�~�"�&6���ƺ��51w�#vf���S��y]G��"Kq=���*�,���ɐOt"�^^!��!���wy�҇S�����\\�k��&���4nmI� *�q�q1ε��=���D���^@N��tm1{�e�� ���@���먾���:�D�����
��|��-�ب*-�ڋǧ����:����J�-w�%�yxo:D��kۼ��t�%.���
E�ƅ���E؊a�,e�s�Mi�����)*U^��ᗬй�K��ˉ��D�A	�ٗћo�Ⱥ�׊(�r�9T�A���j��̊#1���y��WlUwjsa}ܼ��n9m1*���s�A�C��D׃nf�O.DO�w �̀��9H ��@�Am���8H�����@���ԑ���7ט����Ȧ��re������ng#�F��}�w���r{8_�&���!��\���ٔFk��K�)�қ�/��K�'���Q̫D̹bcs!�L�gL�9΍"�<�G73��
v�ve�f��WZ�@�&���F��}�-vA$f�j ���Hn�n<�m� ��o�g�ܼ�ɝ�]LJ��2��r����@�kȆ܉�p:a�y��������͢��&�֘j�G]28��lZ�s)� �j�0�챣�F��
_�ϧ??n^��n @�7k�Vl�O��-r�εv�i*=d��>:�[A�B|[�GOu�S�[��\'�y�>�N�̳�Z��]ּQ�ռ���h"�A�{d�.0X9֤��%� �B�p�6�f�o<�H��U1jq���#-Ι/���n���6��Q���UDWL� ���Bژ���OUd���)[�� �.� Ee+
�K?\�'�8�n�7g�uv���v:b-��43�Yn�jt[P�$U���K(L��ݣtz&ڂ,iw�gJntQ�)�C��y{9CnD�n!���]��Ѻ�.O�v ���fo��>��� �kyIh"�"-��g�]�suSCUo!��W�!kN �[p�U�Bh�6;K)l��Y.L��!��	Y��.@����Ȑ[��h)ٓ}:�ʭ�U��A��YF[2\aN ��s>-��-���ԑ�Њ��}OlW��/@=��+��{K'�iL�P8P�"Kq����]Ñc�}w>΄Am�r'�6�$���{���7��n��˭x��&���5�E�@�[j|Ch!�sh������N\��΄A���M��w1�GU��A��q��mIY�{�P"]����"-�$��EJ��}~�b�O�9���+'�p�;��yuE�7!�#��}T�v�;mʥT�`���.��B^����8bNx���)�A5�ǂY7��������L-.�=� �u�G|�;ʗ��,qf�5V�b�|��<����}lȱ��zlk�<�3��}$��F�\�zH5������w{ٰ�Q�s��{�!W2��ؚ|b�����f�V-�wq:����}��B%b�x;Bӣ��
��a�~~�>C'�,�C�·�?l����E�~\�|{�|��c��^p'��Y��zV¦f�� �-d1Q{�#���K��cG��z��V�"�suW�]�=�X�-�y�=�c�}�r�5���݇��;[�I��8��O��?��x]ʸ@��؛t��ۖđ��d��w�I��ŋ5ہz+g+�F�ȍdY��r�V�l���Jv�tE3�G��&̕�,������Ӿ����n�3�y�v;��v�[t����o>��i��@�ox̳�A����!��G!o���-~�̘�<��_$H��}L���=��ҟ������O����ϕ+(�r�;&�X}���n*� �,�͌��L��T��π�,����PP�gy}��-:����r�[��\߆?/F��Ǉ۞��2����>��\���0��7�k]�;ō�{ʾ�Jx�݀�AwK�9Uú�:���d�Vo�,0�k�¹��c�es�S
�$��y1�����
z�g�I,g�%�NR����qЗY�����'u*�ճ���j�.���]�bɕ�4fJ��SB�a=���:\)	OO\v�4�h���E��u�J&#$����H9pC
)��);�L�S4�D��,$��n���I dbK��&9�bJ@3&c,D)4��)2%��2XĚ�B�dE��)���ܫ�(!�.XҔ��%css!��N�̑�e�$�DE�\�� ���b�2L̲ �PBa(�I�:�a,��h�F2A4X�)V6H�2�&a��L���\�Q�,�6;�W;�� Is���Ē\��I#4!
$%�sbLRd�("ɲẖE�F����&#d�͂�PD�b� �6,Qa\ف@
�U�S6��lՖV��]����4�kx�V��[s���E�q�ã6r4�����Ui5��K]�[�VˡhX�#5���A�˘�T�b%ҳi���vƷ+ԁ���1[[���A��T{%J��ǝ��+cb:,��	�K	H�Wj�M�5`��.�uQR�m"4΃��^6��pQŨ��L�L�ZZ�(r�,�2�N�@�3\��K&��TΆ��S
���޽�A���vA�i����iM��Ե�ؘ�u�vm�^\W�ln���`����gR�lJ܃D�.�yinu�f�U�K5�o��R�xyfq�=�:Q �M�/+�s-*68�Q�.��a���Z��4��V��L[IX�r��mq����͚؈B�a�im3F�;��j�)^��t��.��k��bk,��R����-	qn��kFfՀ�hQ��]�F#*�01cq��V�y�G%�k�h�Ƶ���a2¹63�c�S�)�̮�a��ѷ�f9���x�"eP���-�ǭ"JB�c=�BXQ�U4��s��Io9J\q��*����a[RV���#u��h:�6�"s�\�1�rf���K�t��n	��jR�6m���B%��ś0�L��!���\�m�CQP%K[�-C6���θ�x�(��hG]C�sR�fs���Y�:�0R[�k47n5YY�ٺ6��شJ��is(�K����%�ʎa�M���6�]����5��e����7% G)�cQ8eJdrШ��F�[6ʗ�3[.dX�H��\�0r4f�G&����!\)4��-�CA�%ј	t�]GR㵦��!R�\�.�M)�r�I�`E� c]��+���F5�]F0�3�M b��t��aSg�\l���F1Y���Mu��"�9�x:�!a.!Uu��']���;FaC��[C ��*�.u��i�y&�AF٥s�e�P��m3$Ve���r�jb����mx(͖�P#����m�kc���V�B�)(7^���s�fNYYW@����5*9jj��K�v&�nk�X�����
k����V�-CJ�l�iM��V�,N�hࣚ�,��ZXt�%YE
�n�Xݶl�&X���]�#�V��$�01�`h1&��)b�K�޹c6b�ё�]��EYubJ��t���|>��xc[m����3�B7h\�q�1Ä��k�
暑P������K~���O[^�6�����]T��Үr�^(�EqS��%|��9�"� ��Rm |pvdOeP��^ ��'fM��w:�U��A��p�A�h"rrz����`�V�} N ��D��H!�-���k�k��:	=kNVdV.��&wE.� �9[�A�h/�Cb�3|s.헯;#�P0mȟ6���녓n��Tc��x��w/Ml^ڊpIڄA9�O�m Kp�"Kp7�#��s�%��AxSR;�M���kL�V�p��mCn}>!�4��t=}/Z���B�$)$�-ʻQz:���cg�f��1(H���1[�_�{��=�R#uy��A��]��V�V)������	�3�JF+��� �.����Ch mȐ|[�^�Q��3\
}�$��dl��^��4�	\��ܺ��t'���{��=�x�^+���G(���L�)��K C�pW`9�
ˑ>9�/Muu���d��-���w) ���n:L��Y�/�9֤�� � <hX-Ǔh*���qN5HZ�������kL�w��/[@6�|Ch"� E>��!��ԺFeb�A�A��>m�*�)�Ë�3�)p@��"��}�hZ�^��#v m���D6� ��\{9g^�'�O!W�-}����f�k���R-��p�A/�Ou+��y�=����5$F��J!M�q��m���r�XT�&܌K-mm�.�u��Y���;P �ݑ ���S#�b;{jM5�A��H��0�uX2(b��܂���|[A [�%���ʭ.cn7�����K�R)\�����w�)����͑ �������wx���"A�<�Aۙ�p7fX\:s�b�%�v��	�#m�^���/BR$Ğ��w"�3��;R���C�!D.&�f�����>�S�:�uHJ��;�W�\�~E��t�������O�A7���� [�A �Ԑ���C��MҘ�� �B �Г�v+Gw-!�Mi�n��]�#�͊ܨ�,�ntP#3dO�` q�mI�^-��Q�s��O�W�]9�0_��[��y]@@�y�$��	�.�������t4)��M�ԭ&nI�ɡ2�fv�QF��.��@д�2&bG�bA=p�/PD6����/Ut�pi��|�V�ݹ�v�\w^�ufoVvڢ�Z��"��ݠKp�F��#�E-l{:<�E�;�I��� �������ClЋR�k���^��W�o)��^-�����Y�}s�0{����[��/:����$����A��.�z�w*��2�Dn�> 6��f��sג�ޠ�6�=Ʒ��Ml�_Q|NV�nGE�P�5A�vn�k g7wM;�f�M�n DMf�0�YH���&pDW���b��w�<)���� �%Ɋ�%�u���"	��$6��|ۑ%�\�M�U@k\�r��J����\v#����z��8��!��������o����Vn������[�s����-�v��S.�u���74����8ץ��KmM%o�����fkX��!#\枭����)�ڀ�Ϸb��D6П��WM�Y�X�x�����!U�Y�\���i�͹�[�H>�E�p���왻]�"�Qw-Ih G�l�nD��y�󒦕���ڊD�>�P�G<���w�A��H ��c�D6���Ax��gT��1h � �-�>m��[�2�{�,����c���5__�>�`�ڰD�,���$�[Aۨ��վ��ղqV��nE��Ǹ��4-�>m��]�۹d��CO(���ܺ:�F=������F�F������D�
��T�Έ�`�1t72�`�u;P�|��C�v�C5Y4�깖V�jbb������Ne�lt����(��f����Y�p]���׳�,��@��A��mҌ���%NWRM�ͫ�F4ڑ�"�4v4ݗj]�j� Z0�
=�tΥ3�B�fײsV0셻jW
j�bE�e4�e�at	\�w5��+)*���Jىk�WS�-�Z�K�[��`�Z�K�R�A2���ce�\;J�߹���1�c,��d��3mx��K�qh�˦�pk�-Q* (2�D���2�������S#�#4�T����$��[�M���AP^#^����Ax�����؍�.�\�Pfn ��TS�#4}�fvب�.�"�7b��9S�,H�A�P�q� �����p#*peB�ۭn�I�u��[��sA3ܤ����y��v�ɺ��w"7g���DA�>n,�Azai�9��L����$���.��p���y�)��k�����ԏ[^n)��n0����R� ̵=�aI|6/����&9�zП�"h�IK7�	#fA���qMs1�̲�0�KWj噶70��ɱ����R��!U����Cmy�5���0��>��"�nc�!Ul��ɹ�$3G %��ݠKp�j/�6n�32�k���rڽ!ٵ}����u�Șѡ�V�+�+;���֗�SW��K��6�V�_>T��]�}�<_wdnf��r�x��酧��Sى\i�ؐk8O��h"xz�G=��R�O�18@�m�$6�-�[k3���㯷�iI|:/B%����>�r'Ÿ^ ��D6�F���{c�c!�Ax�ݑ>>m5ӗ�c��u�!{�1� �=�@!�UB�}���AoT���� &܉-�)5�����^�HlA���f%q��d*�;�� A�4�mȟ7�	��T��I+~q�օ�)ë�Л�ܢ2Ź�n�눀Z!Z�*`�3T� �v�Iu8D�S��zeƍ\�'m��A6Xښ��ԙ,U��:�	;����@���%���rvU�1�02.�D�����r�{X���!{�㇏��I�n܆�u�]�d=A{6 m�~-�!���3����GKY�H�~p�ױ���We��0��Y甡�}ވ�6�;6J0H�}�O��u���0F��S@�=*Z`Y�mj���OL��MV�U��]��6��!�"|Ch"�"3�=�%_�7�/�G͵g�패�皂rvؘ��\��j�}�n������@�B ����>-� ��@�ߕQW�����go�u�r,�����)���n�m8ʈ���v��I2�Lʐ�6�v�2��ԍ�HGi���%�"7�"�,��$Mj����bG^�b3�sF��U��,+WE�Sҩq�3�"���������<$fǥ��͙�m��"-�>"�>�躞t9PsW��Z⎍�� d�1�.^�[�1�E�a��D�waCh/ۑ> 6�LL� ���c�����c�?0���?�`����C��p�%����U�D*�d����6�����q���4�vDVt��DnN�b��Q�#���z���m���dHZ٩��?t���I��O�aniUƽ�i��Tt~V�
w�]� ��3#�͘ǳ>/P@�@-� �Ax��Z�E�z��<�����<�3;lT@�p�7�"An6�؜(�13��`Tx�ߋI4�gg%T���D�.�YSv���9�3�΁.���Q�����v��v��mȟ�_'�Y����.��4{Ǐ�[�0��Oa:WWx�B͵ ��@���6�"��/8���+��q���)�숬���"h"cg{����zqz�(�������x�m8��2�U\*����%'��N��9��p� ��D6�}вT[�9�by\?{@�ޑ>nkg/���]��Vwa���RAQH��0�{���^n� �x�۟7"EVWu�s��B`uʸwQ\;M��v�,�q���6ק͡���^��E_L3.�0l�𑘆�kZP�l��KɊ�{� |=��q���b�+w��S�u���^Tz}{9CtI�����f:�zzO�ӑtd黧C8���1`'AKK��v5|�B\����F��p���mA�-)3f���ÛٍYuÒ=GM��L�a��PP�D#��\\E]2�Kl���X�΅k4�՚����k�ŷ�
[���X�sF�!�v%�Dl�!rH��rXi��D�1�]6��f��˴h�ua�̳)�3YRnIcrWC$�lT��q��a��Y����5���O��;1#e��v��\�)@���*�Wf&��+\��q�Xe�����ߞ}u��#}�篾�"�vfѢ�q;ldpCn���5�հ�@~ ֹ[� ���[�A�m9��8[�$K�� ��N_9��-��MF�lw� �r�C�x��P�x �R�Ej@�p�"Kq�A��#.b���f����
�C�]Ǔh"r'�6��n!]��"E*Eq�۬4���n�m]�]�LƆ.���ތ����r1�TF�*|�7�p�>Aۙ�x���@��EZ;TL�Ɯ>nP^��Ν�yo��kV�� ��R!����U�fk�5����~� �(m��RjZ���e���b�x��T2 0Y�	9���5)��pk(br%^��l����w-�:��s�� [�%��ƹ��Ɏ��b��̯�߹�{�گ5��k����\e7z�7a���%�^=��ouf�ȵqS�5ZkK}�o�4��Z8�G�ڟ]���34]���ތ�f��ȟ�4��\N�Y�o0o�A�P��ɴ!�3��0��Qʶ�;vv)���b�ե� A�������"-�$7 �3dCɮ���F=BOt"��OQ�;GeHٝ�S� ���F�����R�����>�c��nڒm[�;VF�I���ivԀ�_cS1�E�.v�dw� ��n��qd6��ΓY?���=���lGݦ���r�n4�u�)�U6X�,sݞ�k<թ>>�����N'��!�"||�^��b�4��m�ե�i
��	���S�h [�%���-��}����x'Ʈ�J5]E��9#em
�C��^ ������L+]嘂/�ֽ~m��"	x��C&T����?T^�Lk�݊X�h���K��#o��8���e/=�<�g��a\9_.s��ޖ�ܥե,�61��lX����>����G�����lp~:w|�n{ͰL�8��m�5e�@�L�]W����$�I����Đ8P�z+�<!�y�r�u��'���^B��$粘5���}��=��溽�}/&| ��g\�)�ᮝk|�&1]�ҍ��ۮ��=�]dm���z�޹̱�84��b�ޥ�o��=ٳ�xǾ�C+�6�C�!�|r�~�fއ�;���������3yI�0�-B2�֬���/-h��)g��:4_r�Nï^>ȼsKS��2a��bX�P���l*���.){�Xٓӌg���o������g���I{Ya�~G��&�(��Jm�P�3p7A���q.�)RB?s_(�x��-��=_�ao5�^���'q�k�����0#]6��u�.�y�ĦU�K_W��pp��<��(��A����\�pI�WN��z�-��ɇ6��0/lȧ.�R�HM@q��'��q�s��Pg����}��^�����y�b�W$&2P�sun�=A)�T�y`t��{�ݛQ6�@��Մ�w���S�ͭ`ae�Y�Uk����������J�j����.���*���#D,��5���:�Bz�?C��0}��n�����v]���Ŀ��AIc�P(^�f�7=�'F*S7��9*E�//	�9܌�y�K-]�3Y0gB�w���@�3���W8C��&H�t��n�dh�C��A��5G�B	�4s��(�4sr��Ln\,�#fI�84��df�Y4�	�E�r���	��Ƀ��i1�i�m��,���\�4c%�p�9E��Q&��PLɀ���gu�r�r���bD�̱̈&!�����s�qܐr�HbH�4����wnh��I�����`��$wt�4h�*	0���"@��c&�-4QD2E�%�&6�rh�$V1���n
)"�M����1DZ�nI�&�
L����$�H0H�)2)$A��Ub�W��k�\�h�W�Y���r#sW��7 6��"1S�鳐�9� C{>��B�*���M:�SZ����� 6\a�$�Fr�s�P9��݄	n �ۑ%�)YJ!W+���C5&U�u��:rC��++��]� �@6�	�p�8Խ��ʭ��F�dJ32�(�P�2�Ωpn�c�+�ژ��ɭ����8cü��x���[�A�m���ۅ'Y5}v����S���Nj���]��"m�s��p���d��,7�����ݑ>;�!}�Xsz�7]��kV�G=֤��-�N�>�Sx�P=:��� O8��܉�^ ��ݺ��ƙuE��9!����|��8�@���O�m[�D(�]˩]�H>�A�|m]�>��&o�`N��9P�<ͨ��{`��N������kͼ��Nl�ZD��v;{^7%��^��M�Ê,L*:�+�}{�z��uAI�U�"+(ڈ�ٹ�`��W�Rޅ��@6כ�Am�ms���t��ΫN9��nb�ջ��u�K�����_a	f�P��i�~~�o�+�].�;Q�/#������b�Rkz��m�0����n���^��F�~�f���mᰨ�Vڎ�Ւ��YH\V%�"���b�b�0x�Ԃ�#9ȟ��q^ ��R����`���Ÿ��)�V�b�L��"v�dr��nl�-������)��@��}"}�x�As>!��u.�|��O�v�)��b=��Z���n ��Rmx!KszE�TT�fv�����3vD�wcɴB�]U��=Y!5�2�.��ug
Y�>�AQ#�'�5y��A�����p}Ӌ8];>�+�_�^�6{H�� �@D͑%��mfnS�R�;�3�,X�܅F��:�=�#���uѮ�<N�#G�����[{�cdK����|����/g�����7���&��-kZ\�3e�$KY�Lb%�����]l��vYk
]p,�\�:Ye;�Z-�Y�c,eж3Mf1`\�K��Y�1��؁R�e�F���3�2���Z\���-U�B���*W��@#f���c������­��vl[�[v�t� ��,]y�-���#f�׌�3�ԙz�W5	(��;?g�����d�vJ��Y��@Wj�c-����J�n�XÊ��.ٟ`���[��l��������23Q����.��Gx��*r��p&gv�o�Ux�q��%��ݠKp"4���Õ,;��o!FraQ뭹�;�Mm
����"Ƃ!�+ia��'=}h#}s�$6��@|[j�Qѱ	wIR#;{lE��E��6�\@� !��$�"�Aۙ�*�l��n&�4�-�ٟ������;X�;ݘ�A���>#I��v��u�e��;�a��u�����T��[���$�a�]3Dv�) �ByU�twV ��YސK�^#m�Kh9j�]e��d�P�))�d�X����^\��ZAHcj.�;7P���FA�����n>m��V�4%�2-����(���5��|A��ϹǬ6�6�A�^"S�괍&n=U�o���~Uuq{�^���irwɼ��C�d������]6��R�n�V�Փ���d��E[�����Es�O�r^��ţ��յ���َ ���|Az��4���F���-R�H�܉-� ���ڝwsu�㪺��ڌ)��U�qwC۟	���8@������KT�6�۱@|[j�)�(3�M}Dm���rNxv��1���yO�@�܉���Cn�剤��`hW'#W㻱�aޭ� ���Au[� ��'{0��@0�H�ĉak2����Uci-�l�+��aS3�X�m�QŢ��ք��9�>n,��.�]j�['����Ъ�	�ޙ�}�b�l9=�d<s>>�7�ԟp���S.-�p�n�N��]�{Ľ&�΢6�Tp^ʀ���$��z �R/J����^"rА[�&�^!�"|[Bz�ENV�ò/�0]3,�s�:O�j�9����ɚ�n���{|��8�Ge^�" ��EJ�M�F��5몧i�n��-���X�n-���1��Ӫ2����Mw)n�^-Ǒm�!�����Q���3�D��B��^�U֢��w�r�����^#�;<7����nB�����n�ץ��qf���	DaJ��*|Ї[�GQx.#�0kC�p�6���s4l��`S��a�T�ک��lX��nZ�jL��b��,l΍\[iSD������ �A�^��U�7��o74�a�ݘ�7!58V�U;`/�D[jA�>��[�D�wW:��}�]j2��%�+h*�8��A�@��ovڪQLg�� �ބA�jA�-���mEh�T��-�yoG+����#o�y����-Ǜ�D6��޾��W!��Ă�ι��+R̅�s��f(f��GMw)#*��.b�$M�%	s�&!�F[����陜��Ե���ZP���L�;F�H���N^\��+aͬ�զ9���VE�s��Ǳ�7~@��|ۑ%���A	����M�ޒ�J�
��]�h�ψmy>��~���̣�L�iŋ4���e���44ݝ�e�13Bˬ�XZ�޵�~y����k�ڂ-Ǒm�j�#Ju�m�u[������X@�A��wamCnD��@���\&.�"���> kA
��Z79��C6�j ���v�E���ny��'�W�my{� Amȟ�x����d��G�	���qu�m�nV�U���^ ���ϛ�7�.����O,UZ�� �m{�(KmH�U�S��v�{ո1p@�P"��$�f/��j�Ʋ��!� O��!��m�ޞ��Q��`O��q�c�;�.(f��G��R퀁n� ��uK�s�\�鸦�<4����j��������/w��<�Q�W��]���4�����kS��3�#4�c��<P���[:C�ڽɌ�4�%I>^@�DTX䰖9�Ց�Kp֥�nL�eƚU1(́{l��5�0D��A�T�����qe�e4X*�5i1i3UF�&�-o��5�8�,�lajX���ZB�rcbf�ו�l҃��I��]]�&���(m�����ц�ۑi��P�7:�0�kQ����&F�����M(�+�nB���N��%�**���[����X++B�ku6<�ˑ�ųV6�[#�.v&�؍[�c;P �ޟ7�hi���t��.�V�S�$Wm�):{;���I] ��s>!���%���[��
���e�(�@�^�"�u�ҝl�+�[�/:��#��>n�#g��������������������t�ṏ�93ov���^��-ǐ���6�DJfv��u�vk�0.�D�����]�w���;�[ANw�p���bc�iS��`�7�'�o/7A������z��5]zf��|�
՗�T:�6�Wz��@����nȒ� AmƮ�7�H�
�!*�pl&�1Fl� ˩�m��h�RV�v��X�VS�C,	�A�S��^ �A۟O�h/WL��ѹ�����v��
��=O�s�7k��@������/896��;�§؄�umT�}2����b�)N'��w���{S�p7��<�n���nղ���a���*���pԽHV�Yi�yZ��@���7|-�Fr�N&6�����cA Cn4a-�,��w�����级��^��-��bq���{�E+ge86�Wz������9�"An<�
!�"Gvݵ$�fJ�v��խ��>n�##4ngp&�;ݨ�Mv�!؞����OffdOz�(�wyy�@��x���q�\B��و��E�F:�/g#5u1Bg�]� �h Cn}>-��،��K�����a�b��L�i�ܡ���5d�6��V����Ɔlt.i��%���������ѽ�jE�M�ه[�J�#p\���tnH��B�`+��-��@�BKq�Z��ʛ��-
^�>̀�Z��f����P�{��v��n6k$?B�>ڕ`��'vۑ%�Dз{:o"�+h/�B_K7qj�mRy�f�"'ix^׽;<|ޗ�0N������k�;��J���O�O!���s�!��
�~R��H����bY�	wF4n����-�!ghcX�:���A�A�@�[j|.�o�u�nܮ�7Oy���kخUy���ta��/۟	��͠�m�l�z	g��/�?9�3!��ٝ�6hc�ڎ>��> ��q�[j;j�7g�O���ib�h��W,&�aU���s�m٘��[X���1%O�Ӱ �͑ �h/t]�eÜ���Z��9�-:��\��kA�W�͠�[��jN^Ga]���]�
���{ڳ$�x$��[������.���$���u��S� F�H=Ѐ ��ۙ��hr'2��]�1Kpvgi�w�Q�A�� ���yڐCh!s�����ذg+%u��/�	�݄-����v\'��u�m�Y�A�"�P1�'Q1�f��j�'�kx�Q�* f=}��ۙUY�seQ��у, �̣C�F �����CqK�2U]��(9a饳��G<^�v��n<�m�#[�br�e�E��{jF����)��jf;ۡgx/:��9�"Kp�!��{jm�����R�_>-n���� �5����
̦�D)�'
�H0�mM�1�>{4��Ù��6z��|q��!��E��p$c�ڎ>���[����[����|�RCh/79gq�YP�jTFZd Gt:*z��_ub6ĬC�w�1��������|3�.=��oyI6��@�[k� �q�F��Ҹm�S1��<��F�B@-��D6�H��X�[]t��� � 3��>!�. n-f��@�1��G@5ڽ��N`{���\����yz��e��PY��5ʯ
����ޑ0�@\l��.�^�F�J�vО{E����D���	O��[Z��kmmj�|��֭�[[Z��[kkV���[Z������m���֭��mmj��kkV�붶�i?����$�HH@�T���$�Z��;kkV��mmj�x�[O�$$ I?�HH@�~�$��	-[o��d�Mgn_�ܑ~�Ae�����v@�����|���P A!@�     ��  $ )@ )E   g `ꂪ�UP �EU  �P�E �� 	(PU
�F}�E"��EA*RJJR����*T�)�B�R�%B��IEPTJ�"��  F�T*"UB���0wwQF��u�[���5�����)�"����j����>����֢��Që�As4��YD��B�}@9۽��� (�>�_)T���J�PITpG�2}�S{�UɢT��7�$�d�zb��<|��BJ�Wv�>���lU%���Q��TIw��*t��-�`:s�|�/  �<P �x |�z�{��=tz||$�:z t�}i���hs�%p�� �c�7�|�t��@>�P� ��)T�*IJ��R��� ��t= �{ x� pz�t]: e�:>@�;w��@nϠ���(�� �C�F@g�+����y �o@S��q!�7`#��;�Gv��( R� ��T��JD�D�B��O����N@|��误�T8>���v��F���l���' e�0A�!� {���|ۑ�[ʃ�dSvr��:u8
te	�$��%J�| �>JU"R�T�J+Ϣɔ7c����@�;���K-����ӹ%1��4�T'��=(x��B��J�!,8v t:�vuD��8X�#�ҝ4�١�`  P �F�JTD�C@�2h�`F� h"����T`       i��JaES�       �%I$� �i�� Ѧ�4@BQ5I(��2` 12zC&�Lj@&��M5=I�d��=SL�4	�z��>??��������C >߶e�����9E�ww�!!	p�8��	G�@�$!���I�z�  �*(�G��("(� �����������~B�/DAH��YD���a�)	L��$!�=}sU�w��A�}�?��߹����l^W���!����}�k`5xPQB/��c��׷ս����_[n�Uf�m�]e,t���h��R�U5\X����̋6o5�wy����ۛ�a<���Jʛn�n��%�[݀�i��hź��e��a��u��.�p�&����Wm u< ��LrU7�n�&f����#��!�ʌ	,�ºɏ�kSM�&��$�X�h��*�λD���aU�%&*o>mA����J���=4@{�/EZ�/���	{ 6�ư�[x@�l��[�L%Z��وqۭ�[+F���U���S���hP�@N�o$�d�3SY���49Y�I�*<�F䱔)��.m���8◇f&+WFHt`�`��D8�D�FR-	��,˫ڽ�˳wB��BC��+!�1��*n�6�k1ͤ���I�iݣ�oH���765����P;*+_;�"\�n,�d���+`Ef��q�Y�,|cK`T�W16�Z�(�sS�/q���\�Q4��M�6���-[��I�nхF��jN���5Mû5A�K�	;����!V,�Ղ�e��m���C��;4�/r��+j���(6�<�a:A�n��d�6��š���Y��ԳV��F�^��z�l�c9F�yY�t+&HT����Wy��f����*� ��[L��a��jW�n�bcU���i�`�lC@f?���;riڻ�� P�Yt���*r�e�J(6̭�[w%ˠjъ�6Rf�BKjYZ4ǫX��4�)�F0�,pC2��i\Z�!XkE-�0�ŋE�bX�xU1p���d�YY�%�Fp)��")T�Pi���"�#7PU- �t�Eu$A��ݫ�Ȗ�C
Z{��k�Vk�"s]���蹣v�� A4�i�R�n�����-S���PNQ����`Y�oi�C�
�W,��Ӄ\/�tZ@]#u�R8��bfFM��.\f:��[pI��኱8/�0S�Ɉy����p(��W���@����(&U����bVH��/�jCI	��I�Y�[W!��wk�[6�A�p]�`��c�@��1���v��$'F��fic-��i+ʠq\a�B��$1K<��fb�F@.�j.����0�8�v�"s,EH#Yb�t��ؤ��D�4*�z�#���h�`;�C
�����\���[�,܋0�����xn���d��W)]��f�F:ZK�V޼�w{�BX1(�g�>q
Y˛�Ob)���B�ƅ ƶ��H�5Ӽ�5��u������*H�0`��M�CO�Z�̖/[2�a�����S�2�ܭZ�+&eѨEnK�ŔU��e�X�`v�F�;0e,8��c	���%����5��"R�x�]H����͠��RY�M"�7l���*ȼ����;w�lXX�zM��p�H�nK�r���כZ�D��vP��,�`��)�1omfn7vK�5�ѐ٢�{Ee�7m���y�ث&�5�-��x��S�t"��?7�8�c�3�w�a�M�(�������s$�50�"��X�
�It4�W��P�6�	��Y��VBSRw+a���L�6��b�n�u��,wv>Z�Y��̫xF�͊nQ&ɘ�Q$�&pR0m[�q���MS�wF��ASF15b1A7����jԙ)I"�Z�K�ss�"�N&H݆�ӚC����5|��ì+F�LՈ(\�k���U��^���T�,>C�H5�Ǡ�B��xE_���ͱ�˰��e2ݷy��5�ދb]�p*�V��Z�/[�+��{��a]��7�w6,��m����!�q�EJ��m�6pGi��I�j�S�Y��CtT+,��Hޝ���@�r��,�]n:�0&�e���,,�ï2��RbuǗ��-�uԱ�0�4���v�Wn�	�t�6�eQy[��\y��b�����Lm ,��d.��4��heٲ� W�Ct��@����k�`�c+Fk֬�^�
7#�fSEZ�Zj���ك-6�m=���-�؊���&0��F�u�G/G���<e��&����պ�Wwl�.�Jө�4�{ZN]�����MڔEcP�ܳa��Y{wD�6l�X3dYY�w�ym�ɗF���q�-�K̪�������M��� �e^�_+u��ɐ��SN�X�1�e�o[���&�f!Z2��ދ���Y'k�{!���K�6����{"փOHw��L��KwA����6M4�k1j�;�e���[�[����[kK�NGb��9�8��S�1�b�m�i�K�9�r��{XE�sF�;٦�h�ZP��U�[�L
��ӛ��Yl�͸t�&�n�E�![0��f�	ּ&�I��R���h���^��T�TO�Miٻ`��QZA��S���ٖ�Ҵ��ȳ[Or⬍d����4��5^Hέ�ӵ�FK�p�W@ԎV�ʢ�m@4�em8��n-{�p�uw�3rPwj㨞�/jH幁jY��dr�7��`��ܤ�d:a����M�z�Q�ay�Q�P�X�u�tB�VDӘ��4AѴ��%�XL���9ɑU�ۚwmБ4B���W��*,&Y�VN�q��9�`��X��ڱ��dݥ��:B'�`�/p�b��.Jͺ�#�X��k����,hh�kl��@ku�cB�\O��ZQ�ԩ3�����/@��i�/2��sb�M���+��C!���ݤ�:��f�Qa��H&M���5YgF���;�tI1N�$��E3��E� ��"�)���@""P-۹k"��ql��+E2���*��wOb֔N��	�_����k?�7�+T�5f%x�q�ͬN]d{X�TNb7	�����F-˖���˺9��/����Z�A\�P�mc+(�W�5x]�&�&�$�uu�$�2^�ɠ�V�BLzi�J�>ь�#z��{�)3sf�m슬����$vq��6�^�l�݂/VsU<��7t���3*�y"1��k
m�@
`�9Y�t��ɲ�6 �yg�o+6��e���c��˙e�c�Y�z�l��&��״���(�k La�%Ѭc+n4e�@��x#��!�u',
����*X�+�yx*q
��<��1�J׹��Kٰ�P��r�($�ƨ��W��]ⷌ�+>(�$U2Qإ��
9EAX�e�-X,�wr�yR5r�P�uC)f�Ԟ���Wd��ң����3LJ�ׁ#{N�<��ö��b��˘Y�����j��׫s&އ��Swxa�F:�N���4d����%��8Eø���%����)�ܰv�yp�3mᡒDz�I ͉����4$�8Ϭb�5m�TR��ȓ' PCv��m�bRݚ�%Z+,�K�",�T�:Vz���HAag6��OVcЦ��Q�{4�8(U�$� ^��-�xtkB��7�S�C�ͭ�/v��Hv�LY�$����X�!�
L��Lsa��u%qڑf���ރ�;���ߍ�#�]f��QQ�
n�Z��պ�S�a|Z��SmБ��*��E�h+T�V�a��FEc�ͧn�X4�zFϬ֬��i�Q���^��,]�E���CYH:1�Xof���9.n��UŘF����;xȶ[������,��e	8&� t��\Bh&�N+� �)T��4���[2�؈Y5�1FAv�n���!��+�F�u��ØDᑖmP"�jɵ�yL]ڂ-`j���՟��)�/hS0d9$J���dk��nnv�!&�28C��Q�nm�,���N0F	���9/&������5kݸbF�ɸ6�U��&��5`2c̽�]�de�ٷY����0Z*��W�d����j����:سe����eD���m�hV�z0R�Tͽ�Tl�w�x
M��i8�"fF:RԻl�n�o7�Vf_׈=4Yю"�FX!m룠���䛊Rn�Äb���Aamkܬ4C�W�V��Y�tHӛ�#��n;;jhܒ5!i�ء/�-�5�?[��������+�\i�TY�sp�˫���u�L�(
��7��v�4��*�k@��H�;�*�4�$n��M�C�"Ȼ�cU2I��Yn�.�;Ӣ���a�z�(��us�[�Ȼn�/ɺoli��Պ��Î!���b��d�Q����g5���0��i��PO�,�h�m,�x�Aw��.�vS��Z�l��1��
�wr+�u:�Ol�U.�3�*�Y6M�iҴ*�1A�� _��k��7��4�b���2�l��r]f��acp��F��JtƷ/�z0���݊t�1L�^��u��"�l^n۩��x�*���cR�s#	Ȏ*8/l�Z��H�L��u'����6�^�ݧ���kvc�hV�]���ZT�V����I`���B�
�m�+��4���m�)֭�.�4����͜ y�r��ԇ؋�n�9��a,�$���:Tr*5��e
b��3,��(�D�ߢz.��9�kfl���U+)�G��(����,m�s�
��Qy,��IݵM����p�\������5( �|��ڈf2�i^�z������e��siXj ���tY[dۭ.ν*�VJwl��i��E�\����[��VCj e̸��/0l�[��%ȥ3P�E���
��Z�Ƕ[�9��<ٸ�gt\T��na�L��1�5棔0 .hc()b��h���&i�//Z�3jT�	�&��A`��9' ��e܂�@B����y��Y�r���0����nX�O��!P����X~2��0m�p�{2�6e�yvN�6 ��K����ع�.�674�=��̵Y��3z��L^[B�B�Y��K+u�'ԥ��A杲�,I�Y���VV�]�sq�Ɔ����G��˙	�6b���Z,Sʔ�B���)dT��%S+cp�GlE���v�Y��L��E��y?gɞ����?+RdH��xz�׼��=��������T��Pi�V�Ai ��V$Z@���Z�E��Q�U)�AUhPQZTiJUhDJ�i(R���i
�( ��ZE �( (PR�JDh��@�B�@���A���J)P�@�@��E�(�
P�
�Aj�D(JB�� �V�P�@�a �! (���z=�=z��W������+�K^������X$��>��hH���4��W������ZѪ��^��&�����54�t���lr��V��%��%�[*P�j:LʳM23���JŶ@��]r��ɠ��f��]�e�;�	�\��f]6އ�@u␝yv����u�dF�K��Z�s0Enx&ܪͼ��Ҁ��IV^4P���Rږr����2Y�9d"'r��Y3[�Υiz!�E�sV>���B\3\2�wE)6�6yn�-R�Dօ�h�V�[A��G�1SE&�A)�!�0�A}y�u}�(����N�:^��ƱU̷�չk09���m;�m�����vSK�Hl�<�����������ی
EL""}B�ʫ]�tn��M����\�9Z4d/����E��oD+�"F�N�
���K�rƅl�5��b�
X"��!�U���Q�v)S0Th[E�=v0�N�뾛}j��[q͔�;"��u��((t0�a�x���i3����Q�� #b7Ĩ���YT�㾌��,w*�A)Χ*�<5}�9�S�3jW���[S.N(��S2%E�3��}ci�a:�ٺ|n������LFf��-�a�,��;4�ڰs�,�M��K�����PK�]�	|�'5y��z�A�%Ң6!�Yú��W�+m"77n[�w�lq��V��ݍ��$΄��۪M��Ǭi��"��k�P�ivlu�@.S��R�ݨ5Wj,�4g:���Y.8�'���fnYw��{�550��]Ɉ��)������ʵ�Tק)�zޒ��L�vz����xm���1ָ��ӡb��U�p��K�y�sff�fh�|v�&��CΫ��f�e���f	����XpJO[�w��`�ݦ-wbl�w��zNR��]�(�X�n��V��/�vU�Ll���5��4W	Ko]Z�əs5��n��EU�3��ô�}���U�x.��7� q�l^8��ǥ�<�s��l����k ����Ww��?��xi�I��嵒ޞ�[��sE�J��<�vP.��v��V	��ݗ�K5�k)	y������-�yxM�K7ӝY�vа� �.��n��"��#4������.�%,J[�y�Ǘ'd���5b�^D�R�Q�,�hƕ�6jT֓�A�_i��5G��c�F�*����jv^f�o�b��t��̽��sbtV6+Ӄ#�ܫ�*Ҩ�2u`�Fr�G�v�e�����Y0��ח|��"�7�l����4���+:=զ��a�!�t[㺕�g1S-��:ŝ6L8wT��/��%uh;v�e�!m����T��ݲ��s[��Я3x���QdǴ��a�Ch�@��q�Q�Iu��*A�6��['��%�L��e�A��Mp��2��JY����5] @��;�GKY�ѷ�pۣ/��vilc�wfi�ShX�[�箥���v���;�]�M��p)x��L�9i;�� a!��i��{k�U�9V+�9��m�}����[q�Å�d�ث�f�_k9r������~���\H�cq���1D�gd�PaBxc;�6oX'y�;�HE���&��]sD�2�L��]� �w�b�A��_a�2*rӼ�hZ;2o)yس�G�.����-�(Z"�9��+Rךd�S��R��@t�\�.���c��U O*�e����̀ɣL�`�d!N�����p�6t�F�r642a2�=��2k��z��V�[�q�=6�K������;��I���f��Y�|d���2�sͼ��|E��٫sr�ot�G���J�nKK 6EY�j�������+tq�:����ο�`(@x�$K!��ǔ"�R ��*�P�}HZ{�.H�/��้J>�r�S얎�5XR"aɛڈ���s�+��r(�pf�h���-Eg�ܩ!F8mvu�Zl[b�d"%����x&��YUER«����x���z�T�IZ֜!��2D�ze���v�ޖU��1@(3����(̜��(C3jI�Y
ܨ�Kdn�U
(���u�+7��ɔ��a��pj�.��
�4����-����W�����0�L�]�_n��.t���%s�d}�ٮ�.�y�N֭�D7�7s=�U�Q:(\B��Y�o6�f��rl�Q93�״MZ�Vz��kM-4^N�%`U���1 P5/����0��8���ծ;߶��^��	�M_�a�H	�]��{@8�؞�Fi��.�1];xu]m�*���uh�J]��f��w�^�3x���u�-<���X7rVrtT�sBQ�J�h����]2��Q��î-Y��!�[@�����o{n�
��W�3:���{V�;����XGG;�Q+5�8wmpǼDje�O��m����)�,�+�.���",�3�ց���o=�¥���K�v�2U�[��91Df^\]Qk�_oi�/�����w�SR��Y����2����nZ�**-�B�}�r���u<�';���<�qý5�f�Y�f<�!Ǡm��3.Ă���}qܯu��YgL�N�4�:���Wۛ%��_֯>;�Fe���idc,�(�Y��U�bX�dfd��^g�&ٍڕ犝�I��7h^S��������"8�)�H]�nd�\��d���,ONX�SD;�˝N=���D��l�L�,�ݝD#��ˆ�[�lSh>��:�,^,�Ή������{{��M6�K �u)w�].S�����w�����9���*������΍�O������6����� r]��F����f��vq�jh��&h�l��@����Q(G�vJ�dц��������Į}sa��ų���l£��RU��K>������ܬ��Y�{��p�RC7����/5��tR��.��z��j�,&ŧ��)t��	���K�NE��T*�(�Iv2�⥉�d�����+kĘ�ov�Xǽ��b��՚��=I�kV��js����IR���)���[ �ctU�Q�nȢI�٢"��j^7���Q��bՀ���	��M�V� �5�C`ʕ������/`9�]_q�졺�ڴ/.ˡ��G�_Mo��#(j�X0��e��Y!D��e�9*F�HiQWxp��imA�ϋ�[�V��J�;X/*�߄������&" �����gNեކ�׮���1��ۚ���59�{u�h�F�^�{�G0�$xrr�u��e��rV�t�#j�Pk�C8r���ȳf������!�r@��+L4j�@�'e=	������m4㤴��6W|���]���L�z!���\�+1b���4���&3zMF}���e3+F�ܭ��<c�J�)�34֜k/�ge7�7"�R_>s	X#�{��LKF��������e�Wvh�J�ghCt�J�[]�W�i��Hw�q$��&�#v�!k:\�+7EG)�N=����;��#D(���VM�:t�mZ�ȥr�(D��B�IDl8�h��)�w]1d���:/o�V�΀�����u�͵�2�u�wD>-[H��i���/��lt��M�9O�YN�\WRj+�"�k={���+��.�B	��7��J�j5�T��x->fS��i��eQ��[��y,�V�2]	3I�ĭ!���Э�V*-��#qo?��4p���n*���m����Xwx2O]�s�E������e3-u��U�]3�Y�^���N��\��Z��*��у
4uQx.����`�ǧi����˫���Ê�3t��^\cf&3l,R��y8Ѣ��r�u��T��"��Ki��YZ#���	��u*�C+
=bJ�i�0�LRp��Z���$+��j�r7W��B��uz;kp,�/�^B�8�`������A��#X��,��ӳ���f���*�&U��}�
r���y�����sʘ��2���h*#wH�Gvm�BV�B�9Ы���`�
���ٝ�&3�6�)���^y�6VH�"���������+p�;��ܦ姶�ې0B�uؒ��]w���u�G���*ej���d��aE�6� >d.�������,���Y���LbK��� ̲�D�nTB�=�Y�ξ9�,썇Ɋ��̇A��vAu�S�[uy\�h�,�N}|�Z�qGk����"�J���gF�f�ݖv�p��/>��*��zC"!�:�+���>p)��
�Ba
6s*=ڏ�e��Sڷ}ûR����lX�]��	�nn����T	�;[˲����w&�K#���Wf�:�Z�e�m�$�]��
�ݣ������|b�f�bx��NA��%�([vp�Cɖm튡`�hKKkV�:�d]���r��/wx�3+�Ddl��\Φ�cp=�pr`���:n{,,d}'7��{8��NtA�sBS��q��A�Ix�7ʻky�����.Z�$gX �05���ӓZR�6゗�p���D��'M��ޛ�dQ���ɉ�[%2\D=�W(�v�1.O%&���W���8�{���yf�G���r�
���8����*����1�Ͼ�@�s��
�GP����(m&E��e$���^��$Š*0,ʗ	ֶ���O��⎺����980�ws6��oj����9t�]�?2�B���'[��2���[4�@#�Ln Hѕ2H!����lN��F��F���6v}���Sz<�V7ǟb�_0<�&�`FjQ�v'�_�o�$�Q`R�$C�H�T�ى�V�v�s/��}t�XU岌�9QQ�ز,�x�^f���K>5����԰��m��Φ��|B �ݕM�ː��Զض*�h���!5��ת���1v��{:vG�ML��]���ʏ0��*�6�]d;�0)�Z�&[ʙ�ً�0��vKj�7Z�}^�8w�z!AY� bI!űv�kʄNwZ�ծ5}����K`�4l�0���,̍쮛[���,љ�΄%�fЉ[��p:2��dԙ "^�Ld5uv���ݤ�s ����*�WD3��9.׿��E7���21{FZjĴ�L*8éq2����.2����2���[6u��1�3dF4�68�k!���2&uz��G�-`��զ���w]+c:����S0������O�mQ�^xawnyt���t6vvCH`�ȉT.��j)�2��jbC:^[aH�
�0��)j�PJQ��&�U-��=Lڝ�hA�[�2bP�
Z��$c*݄ �@]e���mܤڗ�Z�K*���ֱ�4e\��]������[YR�f3C1%4l!-�h��Ҍ�dJV�3	{PU%��]��U&cU29׌�i�X3KE]��%�a��+4LMv��B�R����f*�Q-Ò��C\P������p�
im3��j�a��m�6`��2j�ڙ�ŠZ2ݕk��f��nF�Ynk.c��V��Ͱ�h�Yv�k�m����(���	�սf���i�&��&��3D��v]"qI��a�\8X�W7	,-[a.8Ʊ��\Q�5D��ٖ����u���t9�!u h�,f��J����2��Zז3InƷ���,l;���5m4@���ۮ�k�gd�JM.i5�e��y���Zך4���9�6#t��Y�(�+-�Q
�a��F	]�,.����Mz���!�1&�I�E!f��FaC1���4iCj���m�X؂�̀�s��!h۰RRY_6�S���m�ǍfHí[J��Ģg3-���CK3Y\�M5���WF�+1v�j�z�ۺ�a0�hL�, �\::,"y�|��e�aJ������MQ]h�D�MN*��la�Z�J�"���),���V-���.�h�@��	k�&��]�2gG��-	v��pԫ%�
�׃Xjeړ*�Ņքh�SFƒ� �k�ic��K� s(XJ���6\%6��3L8+vi��s���EZhq�������.�)ڸīJ��/JQ��ĺ-�l,pcC�63T�l�)���LEu:��ㅛźmp�TwRA9����Y�,��l�3l��3�0�hS�M	on��2�h����ͭv�9�F�t^�[��7R�,��`��mSB�ә�PH]��!e� 㐣Jn��c7L���<���c�ܖUR֘�&b��i�� jb�s��d��b���e�V^�ࠅ�h��I��1���ϔ�1<�^�yՔt5�U�9l�]e*J�u�5��ٖ�.��W���P3�"g�+�z��5΃����^E���W=���� �m43��#�XA(��R��Ea���8��5�Èl�a�ƙ�J��Zܵ�fm�&Ų�tU"$u��&laz�&��Q$��¥�5��RkM�4c\�6f��(;Q�m	s('m0ne�Z��\D[SH�1��.�3Y-��l�M`��@-�k��cLQ#6�\d1X�Z���s�At6*D�5.�5���
(�MX�2g:�9�.�������tY��(Һ�X�캹�b[�b3mC2��h�-:�ڐ����"�mv��4хuԠ�ٍ.ct"����+v1z����J��c�e�vt҄-�xs�q�Ó%�k��m�QZA��!��i�@����v��h�WVb*�:R3&�m�EU����ٖ+���4�0,*�.�a(d��3&�R�b��
hǃ7Yn�>,��y,kO6Ƭ[Y-UvR�s�[Ie&m�4Z��ŃU�%�kY��$(�0�T,
r�./�n�Gn�.�[�6 KI���D�� ����Kt��*؉�)�E�nXհt�A�B��l�lD�qE�he74]�o�嶢 ��e��R���eubmip5��t���+kL�lLggcd����%����i�����T�X]*�
h�Kk̡nG)�5lѷh0�J��ת��ձ��\���s-�duu-�+*vahh��Xڶ�5M���B��&.��KpCM+D�C�r)
�l�MJZh�e�[��R`ݖ�4f���o��m6cc3�c�ֱ�"Z�t0���71��8�w��	����l������̨�[�#+.qH��f��V\��-
�#3������:�E65l`�QM��v���ƺ��6%�Ԃ�wU�BiN�i�PZGa	MJ�ʎ�`8�/bP h�R$eڋ��	G7���h�k�K i�E��dE&�Z����,]�ɚ�5-����[p��(�%�)Ki�"4�m",1��Bd�tîae-��@�Cm=[0��6���Ջ`��@�m�U�Dr��k�[����Y�	���;@ 3`�"�!jQ��.qa�m�Af�sn�TrЇ7]%[���i4�UY�еU�V�l3&+e�۹l
Qia�V�2Q��3W;�T�+-���ŕ�%Ԛ�.���0�!7�]�i���U���J@[�)Ԕ��4��!�f`�vr[H�U����t�ƨf8����-�8I���0��-*Sr���l �j洘�R�� �l��1K�9�Zl�چ�6��(��h�[�"��	i��� �#-�!z�)ke��f�41|�n<��mb�Y�.#��%Y��f(5����X̶�!��Z��\�DK��P!^�@]���
�5V������j���u��-HLۭ���&!A���m�D"�[��xet�!�i�Uڅp�n�B��r�1HR1 ]+b#";Ut�f�`����\��UڋF���Gk����6)��hLB�p۲���H�`]�a�v�běcl��ku�դ�:��a��"_<v���)m�b0iJ)�и�j���T�V�k�
]CH#@�$�j[�u]��T�.��t�y| =皮%�$B�����[fh2h̆�Gl���y-�l��U%K�J�v����2�\8�^�i��\���V+\kjB�h-� �X!A�*J��T�b63k���aQ����ɥ؁fy*��Lb,��qxM%ι(���emm����ai^� Zk�WE�r�h�D���]u!�E�V�.��L����F��9�uE �j�0�@�]��,#�4ε��L�a�9n����231��˦�r�n�eb�	P�5#��9f{Z��|1�f4�(�-G;V��ͱ֕�Z1�X#6�\j�.h䆙���^&��2�Sf�6�.b�Sm��clkLWm�˴p�+�s�J��Z��\��Z�
�4h��͇F��#�i�k��.�@l͌j�
��ʻl�mc���@ate�����i�n`ڷ ]��Z����WV�l5�<b���*Ռ�,n��L�k��ip���&-����h7b�)r�l���kS�J�+�#te�%I��A�3�K(�e��30ڴ�OZ8�,�:�u�KltAՍ5��*�%2V��#f���v%s����n̦
���6�+4+1��c���쫅��gi�f�r�Wװ����I��JN�t�	<%'0��I�N��9	��9۲QE76�4��An�vt�`<���͚�&�<�'��o.)�gV�v=��c�Ry�rNC��;w���&��׾nbt�Th�*9!I�͓�݂���I����r9y!��C���y;��.d�j����l1r9.�6v�^]��[.ݼ���7������wy��Iۄ��D>m���s�4[M����}��!�r�J`������yܚ(����r�h9/��� �PSHP�H�y	��h+��O-%�<���(���y�'���<��<�ŶJ(���p�
h����F�'���`����4&�N�@vݳOj4�#A͹�JRr�1�U#������;��Rb4Q��[nm7���U�9=�7r�~�����9�ϵ[�۵\�w�;r�;F�mod3�#�vb�R�2kf�R0����XR���-1i���g����) )5&��imh�K��	�AkZG�;dmά�8��.��K�5;.�nsn���2%#�k��ԥ��{S5)(	e�t��!��0�ZC-tn��V� f�u��`�-#t��Ys�Ce��JLdIz���	�E�S%%љt�w�1V�V�E���mKt:ۊ����M�2	���FX�P�6����[HH봖7X�{Bd��t���+q%���Ć���:�\�RU��j�[	vZF-��GRZ4��ͪ\��^�l]
Vl^���5#K��YfB0��YF��͘��U���Z�P,1�B���kq[ua��r64�ז��^�d6��ku��D�Z�#�p��(Y7c�K�L��M�mc��m6)]أ�4VD��6��ن[v7T`���+�U���uc&08riCn�Iy�oB�pe"WF��W�a���[�c�G ���Q;�cuK����[�	�b�GkS	oic[M��q�%�ԕ)��b����/�	���c��qA�sZƙ����z�\3m�i��R�@щP�Fl�gF�k0�Ǝ�L�[ƚU&�.����*�EQ]֐�+���a�c�ʯ:�iY��k�-{*�%�Jņ:�4��v	�i�D�Q]�wwD�Zyi)/ �%ZYx(4"^ �R�����)*%y�e$  l �m�Ą�JT UjXұ�`�A-#)�)@�X%��	U���m-E"�B���#�kj�/T�m`��VԪ@H�����?-"�ĸ��;���˜V�R�
�f0�3�f�����$7H�]�B�|;H��}q1�a��a�W�b�����ۡ=�Ϻ���z!��&wܼ����T�R�!�3�;������5����U!T�T�����ʩ�;��#0��&=�b��]d6>l}M��\)N�^���b�\�od�*w�!�{Cb��C}3�|��J���Y��Й(ȕ�*gF��&��5m��ߟ	���UY�����7�� �5���07�ݪ�U *��@�o(I��Nۜ����苦�N刀�}��tr�f�R��x��wJP"+"�+�10I#e9����h�R��=��^��lw������-M�~oQ�=�3=�ܞ�z�!���f7y{��|t}�)�ݦ{������Rd"��C���lWͶ��w�i������ޯfn��l}�6)����Ok����_a��itG;�H�BcT����niT�"�|~{���U*���|���e�v���G����m&��o��9�4>}��;����T�:@v!UZ���G���ІOT�:�m���T�����ڟ/c3�V�U*����R�R.^wW���x����y<`T�湚��1�9�%�5@��=�/�˚� :@oUO��R򒳳M���e��1j���w���(�,���͊lSr��auӭ�ZOڇ��T�߾L{[)�7�׽�����p�9dee�&��P��m�FV��thex0�����6�b�c\>��;���n�/Uf���f���%���oA���[U���t^��о��z�˃a�M�FQ��ɢp�:�9��Uު]�RUT�H^�˝v{��S�5F��p�9s��:��"�\p������ �%�R΁��L��!n���x��D� �c�Na��t/g�����T�Wf8� �����>���G���Wo[��ooA;{S�t�H�&`���%A43u���q�\�]V2ffz���*�R�ʭ֗V��n����p姸�6���dOp<�M��?=�W��;<�y���!���M�:*F�͊n��l�V�����+��U��6��so`w_�d�m�n��@{��y�lpI�7��xX��M�m�ub�
"f�y6�����M�g�Lw�5MᮅrwV�
�J(�3���!d�����ϔ@��
	��m�����|���Җ�Yf��0	�;����0�K&��v#+\��R��L��T�Ш����eu���ɴ���C8␚���b���j�O���'��®����(�c3�\jLn�GF�ZS6�I�%cE�������ۜ�f]�WJ�����5�bQv��4��'�|G�n�h��@e�9��e��I��y
��b������{'����xFfo�ۡ��Sb���x���wg�w=��y�ې}�v��;�o���l���g�h���׵�7N�Rb����7������n�+�zi�ܙ��{�{���D)l��g���g��l6>lSw{�So�U�2={�����_7�-��o��[��^P���cU�EW\Z�u�)YYxQ'0V��Gƛ���â�2�cwo���;���R��勲��Y.�*��b!�1H�7֮F�p���x���/epa�
�C�b��ꦇ˃o��L������SŽE�:�Z6�ئ�#��Ξ�{���~l}^��lSb��Bq�ϵ��)�VK�'_W�n���Vf�]��]��b��Tئ�H%���;��uL�)�K����Tتl�MF�+��r㋫CB�,5+:4��E*�2�e����l���5������5�M2���f�N��N��ݧb��35t��̻�kz��q�j��T�Sm��i'^���4伋$�>�lZRbr"������<�fQ�Ta��]���ޫO��k�o��$6r�仙{��T�*��e�U��
��^3�v����_�l���^�)��VlfR ��V���2�'�����}y��ײ~SG7v�bV�6�K��%Ȩf�)���2�7��<�٪lSnf���/w%���K��_�����m�^���}¹��;0o�/x�����
{�N��6*�,H�n���ɋf�{6�&잢�w�4�f�볻����h�^�UUU��v�����SHA���
�v�r:�0� ����4M���v�R�T]c э�7#C3���L�|���G����M��6����m�'{f��K�%��ǴSc��N9�փ���tp�De^VfP�4��aj��̻f A��0��H��M�/c��	�'�ʽ�_�ϱn��ئ�=�wB�i�c�I��輻�.�h}S�S|�����٭�M�*�Q<�s�;�s+�3\R��M�Λ�����gD�4��1���7d��6�n`����y��m�� 5�շ��z{w۞��T��`xfu�w�o���p�t��/Q�#�b���Q%MM�qnY�����m�>x4E�Z�ie6y�:�ػJ+�9�Q����Y�x�5uƏ�0���XmUڱ�u��h�cjFk]��MM�a�t�fԶ����fce�l�e2ֻb�FdGe�����b��aġ�������1+4a�0b�F���0�M�������� 8�����\�;0X�2�M*�d���p�������}Y;�o<��A��{��T�g��6�]?v͟8*�]%�uxM�<P��kWVڭ�kO��͇K�Dj}%F�]|o'#wq���5�ک�f��U`n������7���w��&z�Zbu{&䱎����b��/���b���L�W����(w�a��od>�q(�M�)��T��kc4�9ˢ�0��Ͽ�����������'��>�t��B4�{����<;Ͷ�]���6��b������أhY��1J�4�έ�H7�N׋��۷8�ǹ�X�;�7{�f.�ݭF3z�g���T����>�vAÈ����b��s�r�(���i����9^f_׷�P�l|���)��u��$�W�z����5N�`����f�b������Z-h�������x��6'�lS�w�;�˾OGy>���,�e��:W,	�a��fr�m���_G��6/}p���n��+q[G]vQ�|���T�T�R��x�t��������;���m�_������kX��Ϊ�?O�>�G�h���m~S�%�/�̣����%��nľ$��w`ǻ�j��ʎ�`�g�A.���a��J�{F��v�Y��ݪ�5;�2�T������]"�ٚ�V]�;qvX#y��]��鵳��dtV欷ݘ�ar� �������EJ}�f��Z���+�����ٌ>d]��*��U����w���d���E-�r���5��:��[��P#NnN��*�u5{Ԏ�C6�>�딍��J��ۀ��8q邦�%���C�E<v��;X����T�]��x��#�2��t��jn��u`�,a�>��ീ�`�W��:�g�	��^�������ꗘ��]��-LP�9�F�.��͍���}գ��aά�X����x��7yB�.�QVU�[{���,�OK`p{�"��֨�d�
��d����	6�	ޝ��gG;X%�,�G-�@�����܌��uLǎ�:Ƿ���Ֆ�i�Ս��p�o6�L�ծ�;�����(f�b��e
t;iJzvu�g�����y�s�����]��4��f
�u�2=�)Hڷp�*��˻�_�9rBvC��@s��v���x�{)���^Z[̎���f�܇6T���䆎\��T�!O6
h�R��q�qI�C�ä9>C��Iy�\金͹Q�m4%>sP��U/�i"<�B��-�x��9Q���͍݉J��4���k�k�K�tk�IN�.ӂ������]�lPPZ����ư�U��<T�� C�O���GKʃ�;͡u��T`��-��i{�8��N��;�PW/.A�9��hk�O�y����;�S�sy×��������G	��<����+�.E�<��G�����̚Z(v�p�k�ۜ��h��=�S&��VzO~]���
oԺ��l6*[~����@EwO����]�q�yy|>>t�0�D�A_V7R2�=v���W��1���U�>��]�lV�f��u7*bI���A�$�2+p8�A���L�X�(�$U�e��	fUj�� ���3�Ӕ�s�َ��ٌ���Dvwy��2��F�e�EKғ��}~f�U+�'HvU�b�ε��A�t�q��Q�QxN�t^���>����E�0d����nW5�۪'z�6c���T��䥚Y�d��R\E���]�SG�/�8vZBNȩD͌:F��kn�[?v}$m�,��۴.#���:���]��j��D�0��of`�]����F��dȉ*$��UP%+�lQ1lS37��L�ם�w��oE�V� �xF���m�3��j�ڞ������6c�}��F���^�@sp�yu*��qW�n���Ȟ��ۗr�
�C-���Xѽ��[���{fk_ME���h2�8Vf��'.�7b5�^l�y�c�7�K7����z�ٵ��0៚5ݵ����\�o)�%Jާ� qŻY�h�����Z�a����]�]��~9t2��\��[%�����%�1W)z��\31����Yf��@4(LP���Ӵj�貮XD1�!v��͵F˫��))���6��r�9�m�;9*�qtKq���;6�7f��
��1�B���X�v��l���h`͠�)�߯��q�5�dN�&5���,f���b%a�9޼��D��D�u��i�y����Y=7�
'�z�i��;��GuN�-��Vov�=��|7SyU�$+^�p��v�<�����-��͘���׌��kxg5�%���_����(Vb�����Y�o52^mҔ�抴#iR����+w��w�JY��q�ڵ��0 �D�s]̅���0����fcf�Ma�Io�]�$�d�����7�{ܥT��͘R�5gͦ�;W�*&J���t�DmQ��<s@�:[��3uu볅�a����ѳ;B�~<�3/�k��Z��O%���==��^�7ӵ+r`��=�6����z���n�+��s6∪A�����Y]W�1�6�wE�|"� ϳhCh6m�ڄ�a����so�n��C��J�J�U�e=A�\ٴ�]����k��s���C6�Z�9����y|���Կ>����������ơ���׮�n�:Y��
�S���z��\pm{��˴s �;�u�$��
��YM!l�t'����6u��lҝ��ѡj`e�6�MH�G0Ѓ1�lT��Mh�̟�����<�3/�-im6�c&.�]�|�������Q��&�{~���h6�J���܍����[�W��@v8o�2���,��c`$KaI�RP��!��&`.�ssu�*mu�3+4a�|�i�����i�y�}�Uj���Ρ&q�6�,�s�e�끎���[�/m��7Sml֝wSK���h7.��	u]���w��m��l$�9�%�����t�����ݞ(~���j�R�2&�$i�%�3Ы��6�`��7F9�0�Nb�6w
ˑ{�hm��#+r�~������m�)@�bq��s�j�����Q��=�*�p'~���Ŏ���V]6��&�l��.V�a4��r�}�~_�<����ܜ�����0�j�~����	!������9-w��M��P���\O�cw�]-I/�Rڲ}��τ���{�Gu6�>mP��U��lU�6�������97��$�)����zM;��n$~WI%Yz�c1iodho_��稡�]$��'
�Osne�Э����I�.�`��ގT0-�ǻ�Y� ���,W�LV�w����LJ>>BbĐ�D��dB�h,hP���df����iP�M1X�E�UY���k�5�n�Z�(��ؗ1ZJ��l��ф���6�Q !��[�4��-41h�u�[*�18%���������+��+i�m�|d�-Z`c��wϟ���]u[�B�L��g8X9�8��D�d�A�3_��L��t-f��q]��I�z�H��K)"�f�qwU�vb����6_{ͭ�ܤj9Q�:kg��ې�*�y�wĺW����n򯄵�!���##��o$�Z��C�v��oq���݄�W�my�lۓ��Kw����]�����p<�v2�=��|�z��/f�qt%��J9`M��ی(��ƕ5�~��߇��<�y��WMf�WyW�zw^my��T�vu���}`qʼ��*�Ú�u�1;:�U�Glփ0v 	Di�Τ򑓻:��T�K��]}�>�W!����;��w^��n�7�*�P��1/$2��Nj����Փ�וכ����>�RV
��u�HU��Ȇ��I�{�+#a�<)�U/3�כhbY.�d��w{��ޣ�܀�D���JAQ(I
&W�0l�Ql����ج�0"f$D������6�m�y�۵כz���Hw,-�,��-�IF�7�Z���]��z��>�"��pkhK^^"�F�@ ��/6���=dd��wS3��<묫'J��5�v�Hp����������J��cB�]�d��cL�{t��x8Ui��s���z'9E�	L�1�-����f�oB.�����d���]�͋�� �(#&h,�5�b^>����|ϛ^df(Ve��{��{v�8�E�
�	g�}�"ڏZ�P���F�%��)@9����ł�2��L�H11R���#����h?�q_i��q��H�BS4[����B̢���G@<�%^ư@�啕���7y�b��j��ڼ��ݮJ#c�vǸ�'
!�#Ő��#�S��n�ی���*�G��CPE��} �B{��+:qNr�(�x�Ax�=U�q��q��H�M��[���A�n����(�����#N�&��P݂�x�S�~�!��D����y[��<5�K4�����&S�l�/a2��S�Ub�1X�W������c2�n�6���^�B.=z�n<?o]迁	�[��J��u¤�c[���#cS�ͮ��� a��@��D�5�t��=�y����s=N��-sTZ�!��-�nwUg=���	~^�B6���9��n�����p��ߍ��lޯ`�R8����Ad9ˀj"B\�f�r��ܰ�5K���gɸC(�1C���A��0���]��i��| @��VX�1Y�@YCKͨ ��+u�1�J��w5��i�(w`@!� Y��ﯹ����ƂqV�D�&�A��(u��f��Ѭ�I&67�	+&Y���X�$/2��@�2�|�Z6��<5��Z�j�Z�{ݲ��!�l��J�},��(r�p溆]��r4&K}��mF�軝�"=��b6�@�U�Ww�GZ�j��%�5��m<�V6�/{�s���'Cu0q
6&�:�,�w��P��r�������l0�)%�����.���mw-��ͦ���$�guo+U�a"�!�R�Q<�($�']��*rU������1�K3n�kp�Jf��-�̲7�Pz�uǫ���CZN��v���| Zp�1M��V"����
������`7N�+��|����JT2_�7tje�V�T�g�9�D��[:##��ޗ�m�3�6L 2��YV���-��z��/�l�ce�c�M�網'o��uz�&*�|��һ5���[|��h�7Fv޽��W�-r�o&VE��se}{��!۾��f�=2�^ѭ:��q�г�ϳ�V������#g��b�^B4��3�uK����r�i �ۜ�}�6���rЗ!�j�r␧f��Oߺ'׫�a Q^���{���g�P~�Q���_"��k��'o��v^Ny�7��{s�44vu�Mw���mʎO9�>cs��1k�\ˢ�����n�n��On�򵣐�4��ru�-������ll,�Ŷ�1$l�&�^F$<���I�� |��DJP�A���P�+������62�5���$��n�vw<�<�`5�H��g��ܳA�C�\�<æ�`�=��vJj��B�;M����4P���I@Dd监whJ6���G6��p�CʎN`��B�� Y-��S�[&��������Ε�ȴm�a�������,�׍ƻivF`�ae�[������U\�u�-�Y�BWKfÀ����LDf[�ғl�mU����KK�5����+��lX:!2/$�����x�Lݳ6��#�6��L6�sڋ4���;]�J69����ln�Mt�������@�I��4�b���z�1mX���%5����n�3p��)��v�cV쑉m�Z�u��n��Ji�V%���Hb���V �]�m)#BQ0�����l-@�`V�����TMcM�VKqed��g��.��X-��̵����6��a����Qq�E���Z�8]�c������p�tn7Q� 3^��^"d�Y�n�PK1�0.�j�m��4ְػ511Ĺ3
��$�u�4q�M䤺YMƊ���k5�c�Z��Y4rZ%��s
�c)x�v�ጳgFb�em���h�	Vk)��˭�+�i�nTf�*�Qcu����p[T���+�,!*�$����kς��`���/%���4�u�sq ��-��ã�a^(�)�ڂ��&y˶B!���Ke���B��qb^\Me�uDx�m�
�a̳A��ԥ�f�!]����;1���GTf�8H�L+m���-�-+&�4�W]��VZ0���r��u3�Hh�p��.i�q�V[K ��vt^Mch�&��&E�e.��ƶƩ�rݗ*�	�w��y����Y����Ɩ8m��ńK���5uvL�$"�y�[1b�;�&i�e�� �j�bS:��9M�$ã0h�����u�� �Mm�F�i�n�kB%3�6�GBˉ����&�V��� J˺����6Е�`X+�K�k���i�S�{��4�J¬EiJ����6&U��"A��&H�@a�R�jJ#/~ſ}��+7,2.b�a�{��{K l/�20CK�,�&/��Htb�������*�@$2��k5�>�b�(��h����[�7���Ѥ{���	e� �&�""PE� �Ykz�ow+Ǜ��R�Q��NJ��������C(K(p �]u����cJ��Y��@���B ������{��%�1�ɁDB�	@�*(����T���D�e��&e�#|k2���H�w,�kn�i�A��qv�x�r`A|�(��@>!����:.NB�}G���f�o�j�2vw{	ӳJO=�k|+�9K���1�޹��S�݉���xM�m|}D/��~�W�7l>@��(>�!,��Z{n�A|��&�d3�;�����Ա����>D����i�و[�� ��jŸU��ot���#�&���gu��:ChAg�����
����܍��x�v��	�^�^<�Cp.���~���z~E쪱��֒��1�JD�)�T�9	��h��,��er˱W�V<B��tL�e�'�O�r� �ב�8Ǣ�JH,����9����;R
��BQ��(J�~��%���w��{z��<`yT����R
iA�	I���v��iv�k|ƻ�s�����
H)��I�J���	BP�y�)�]'���%	H{�	I~��|>��u���[d�Y�0Y�i�5���	�fV�Y��4��|�Ԑ�ض{�s�<u�s����$�:O���cBR��	BP�{ӘJ��rr��C-2̔�P��w��
�i�!�����~�;	C�4��(JL�S����[�;�v��t��\��{	Bcd=�%rCBQx}���^ڀ��`B�P1���&* a��o�<� �ϕ$�:ߜ������k�q��L�ɡ(4:>@h8C�)>���J����:�ѣ�!��������~�m��m"ܡXفQa�����v��3"�������a(JC�+������ܜ��t%!�*;�9�-����a���@��������z�n��%	H{��%	BQ���P���ܝ��)m>2�J�`4!Д�7񯼯9�[�CĂ�SM$��d��0,y��[���c}�Aa�Pu�%	H{hJ�!�(�p���d��j�/z:s��A`x�%'$Д}��r�������%!�w!(J�`4%L�*����Hhb_�M�����4��JH)4�I ���NBP�����t%�G���I�sAv�!�:�W�������Д%	G`4%>��>~d�RA`e�����{�[�<���a���C�Y �Te0�jH)��lu��
�RYy�~�k��Ҽ���/>��+r{P��D�ޔ��Y�9W�cZ��� ����i!G�a(J�{����%!{�%	A�:=�Д%'}�vH,5L�ּ����A@�)4�Lǘ����]5|�H,5��H(���Д%	G�	BR{�NA���̛ݡ)=﷾s���x�YK�yjt�BV]�뭺�d7WDʀ�}�,�ll��P��<���4%!��4%���D���B�3׷�y\����8�|�gY) ���~��[͏�������;	BRv��t%	G�C�hJO}�۩ �3T���
v�Y���z��8�Rr�d��X�R�~sv�9����AL��,�R�=��J�����)Z�`?���w���P������J:@i�P�%	G�á)=�'!(zA�=ڗ��(=�#�-������߾�n��#��
���%!��%���Jxˤ�ܜ��:��j��RAL�d,�Y-�oS��56Ú�Y �7k) ��$��9�Y �L��;޾W�9�t0<�Y�t%�G�!Д���~����|�n�H)4!L*�KFRA@ѣ�BP����˰�%!��%rCBQ��!)�.��rYc�p�<�4�X�RsZ�m�y����AL��$��Y�Y�hJCy���hJ=��1 ��jH(��-����+����\�ë,2ٞ��yu�ꓱE�H�;
��9��y�pn���<3W�I�_o�mp~Ա�9����j
��ن�Jڢ�A�P�!3�,�!.\�գsfi�^�m2�X�34;U�tcc�b�]�)��m�����d��Q�0<:��/e�qQ��3an����Kna��ak��apg�Fˬ���S�6�����'�ɳhhĊg�n��c���:Gv�777{���v���Д`4!Д����%`��B)�I�
`s^_gy�wn���t��<�Y �;�o\�`r�H) �����%'��NA�:��j��(��r���ܜ��%$���w��H) �3j �yP�AK���w�|�:sz�P��?ĺ�C����)9����J�iv������_a(cG���hJO�0v�%	�CݨJ�!�(ǸBP�����`II
fԤ�;�+w�w��gx���m �P�H,��a��9�Д���P��BQ�a(JO}��J;�=ڄ�/�&���K�RAH,6sv��=�H~�K�Д%�i>o;�<�g��r�d���U5JAH)/�\�;�Q���
Aa�ܜ��(?�?9�JNI�(�A�J��rr�hJCݨE ����r�{��l��]_ʅ�
sO/��\�t���`yT����BQ�A�	I���;	C�)��� �%&P)�ζ�s����9����m"�G[�cW�VT��]���C�+��'@��A�� �;T���SH���ܜ��t%��j�cz�������x���i �P�H,�Ǟx&�4���Y�I�Z�����(���P��=�'a(��=ڞ�J�`4%	^\x䑶���Ζ��M|��w"m�<�]1rp�h���_v&�-��kl��5�a-�9ݵ�  _��
OB��T�Xe$��@�{�����z5��~] ��*H)��� �Ć��~�9	O]'�����ٵy\������^Ԥ��Sht����t�~��cBR���)���s	BV`�ܝ#���ǂ԰Ş/�ʅ�|w/���) �Ԕ�@�,$��Ü�Z��=ڄ�(J=������ܜ��9�����c�P��	_����JxK���' �: �L3jR5��\�_<���s�i ��r����NBP��7�_�z�����S�-D�Ї���%`4��P�%	G���JL{���%!�Խǅ����'&�
AM Sx�4g}�Ӝ�}�Aa�Ptn�R5JAD�(����%	I�9�:�>��O��]��w1�B���+Ut��
��S���I���.��7.w��O��|�� �%.gI��N@v4%!��%!�BQ�
H)��B�.gn��]���^o]�*�u��
���9��;�-�á)7ϜN�P��H}ڄ�(��	BR{�� �3T�сI-����>c�޹�H,�d��d��XU)�'�ߞv�v��w�k���
e���)>{��cBR���)$��_���kѲ
Aa\�r����jxK�(4:=��p�BR{�NBP���R���(J=��~F����8s���ý�}f��ݹ�77~oUY�z�W������C���c@�5��E���`[oi޳�@	1�d滾y��o�WH,3�M�%!��%p�Дo�!)�O}��;��Ğ�P�%S(\B���7�=�76�֨Y��)~�%	BQ��0�Ah�jH)|������כ�@�ʥ ���@���Xw��k�����x�RpB��R
AH)�!�BR{�NBP��v�(J��9	O%�{�NA���<����a �7T�;�w�_��q��:�a���C�Y �S)�sP�AHR�P�%	G���`���$xБ�B��?��$Ș�Ee%�l�yì�T LP�u�ss���H~mO�t%	G�	I��NBP�!�ԼYI �P)��ofy�y�Zؾ��Aa�Ptn�R�{��Y�����*���HhJ7�!)�O�̜��)v�)<dД{�)y:�sP�Ĥ���3�յn��)���
x�kQ ���P�AL����wǛ߀q��RΌ��R
i�������'a({��j^Vog^s;}g��H)4�L4�T���a(JC�j�!�(�BS�t����t�BPbOy��R��Gќ�N\^}5���j��
#`�9	K�I�9�4%!��	HrД{�a(J�{��
^ S5K,��P�1��y��?��4%	I�?8������R�fRA@���0-�oz{�|�������;��t��X�R
@H�$uw3���P���S��&j2�q#(�!/��$��H�ơ�a�Y��橾1{�sY��c�!�?��O����v	A���(J�`�!)q:O}��Ƅ��R
AH)�g~t�s�	s|�����޿��fiA��@,��.��7G:)ۀXuy�����k	+f5�L٘Z�\���i�32�l<���X�ڒ��m���D�f����,������XE�"1/�,��(���oV3<�}�0A:VE��ޥU7!���:���B�yd#v��ב/�,K����>�x�N�f��Ew AdY@��C���Q���>�D��^gӗy�;�=۵zğL� ��oE�m͉�Vub��a�q��{�S���n��Ҫ���,�u[Q����r��`�������V�����UL	�5��|̵|}�-���?;������ҋQ�o��y�s��1s\�+��s��6YX�Z�V�HV�.mtؘ��mPx��p&ZL8�B�����2���f.��6��SB���͘3���&�]M��J5e���Z#�l�ٔt{b�Jƫ���%03q��ev����"�c�J�Fm
�,cϿ~���v(U$t���u��HFnƍ���ΰ�%��,��K<�h@mou�}�s3H�FL��Րn��3V��^ϛ�χm�b��Jo|�qא����ڽb{�ͮD|Ώ|ם|��8^���<��I��J����f,������T܇Hp!��mz 2'��T�TK!x�K�7Z���㹘4��^",�ǙwEL8��%a�hI��A [M��w[�☣�7�q����z�����}�����}�>��돐l0��Xj�XEJ�t�yyX��6M�!B�3.�[�Y|YŹ}�Ҫ��:B�JW�Q�3�Ã^�RAk��E�5��U`�]��j!�Kp�+/"��f�&b�g�aH�.#��8�Nu��
j;�V���� _{ "R��!��{��㹙�p>��d,��CԞP�I��Fd@ �� �-� ��ά���$WE+Ν����ڂ//�Ÿ W!ss�8 NǴ� �V�wf��L:�������D��)�~�XE"ڂ�9��*�V{EDػ��s��fi�h�d,�%��R���Qb+^2`tș
fA�j�(���:-�l�����b&Hoc�|���ԐZ��՝��;]�"��c�j�A����[��eQ<�F��n�2|���������SrtY�Aڎ��yJ��W���5�}$4�A{�F���2���n?w�P�^p*��v�2��t˲��;����m6���[G�\�����
���f����6�*�M���O��M��T-�������Eb������+_��7�}�/�i�����W�CZ/\;��P���0���f��B�Q�C9)a_��՚y�m84����\�y�A�� T�`��e��B�^��]&��u��-�>���dr���;-�b��k����H��.�	`���\���L @����Z����w��GcA�1�4��J;Ň;x*W���·(��
�IX�bth��g!�5�nf�`�i�m]��7�vd�yr�eWh�3�<���-P���;�|�(��m&��Fc)FJ�;:ۋ���S@�_�v�+V�G�ov�&��=�oc6B��;�^<��l�i�1���)=�R�J�4������>��TaK^vt=��f���i��uc�ɵ�sQE�J܁N���z�z=V�\��y�.�B>#�RÙ@Q���_�]O��/2��2:-�F�h
6�E%�r.c��k��EhtDM��Ei4U�4��P�&����N\&��!��9���l�Q��)i
R����i���sk����U%EQO6b�ӻ�DA\��m�()��J�h��F%Ӷ3,�f�CE�
�� v���@U)w��y��
����ih��N-#�M ���X�#%0�P�$�U��Fo�x��Ј�I�س��\4�ŋ)��>C3K�׺�ue�5���D�@�ڀC�;�4ш��^9� ����y�.��`I�[W��.��u�,���מg�gw�o_���/~���s��w�As��@�lÞ�6��;���6�������{��G���f��{�w�T�q���<���I�ChA����Y�"F¨�y�]@�v�Ϯ�9U�����D�L�v�"9��3�?%a(T��@3��=yQ5�����̻�a���� ��σh\����Y��8���������Vv���#�&�E��qZ�sw�a�q!S�%�`�J}0�܌�u�-bF�!,�'�8�\�`w}�g~� �2t�Tz�Cq���d/֟�g�����~����kdO ����C>mL�����V)W�fRs�t��G��KZT�9g�O��� ̂	el^mop�sl:�e��;��(�P@�^���PD9J-��h/;B<��oX���{��q�>́�t�;��{����=�/gc^y�A�^�)������]d���-�r�Q�ŋ8C8�ݭ�97�����ޭ��nC�8|���*wō�(�Q��/6�Ϥ�bchF�s ]^F�	����GMf!>,��:3i� �.��m��m��K�7�UaU�F�{L�P��!��0#�8&���M��geJ��0�b��om"���?��{�b�0���Li�<JZ`���J�qa-�2�E�����8# a���V�^6A�2�e͚�$.�䯒�o�P�iiq��Ɖ�3�m.Z7!�GW�4b���[V�XK������δP���@�C]���ۖ�k2A���������f�+�1Y���Ø6/h��u2�e��y���GR/y�Hyz��{ѕ�l�H�B�ރU�qA|��G�!2�/5��p@2B������u7!�z� F��h��t���7=g���5�k��^-��;���EDN`���{����]�IA�Cp 7}�'����/�^���Y[�Gf�������}8�F�O�E �wc̉Y�nDmE�F-���nC�8�ཨ/���4����O�,jؗd�����BY�lš��]*�a藯�G?g������>��z��iE;s(�58@E�n#��'�V:��FHX���,���$ոt��w�����Oh��f����`S�&i��-	�  xx=���E/!�=ܲ�~Ք'�8�KyP�^g�[3����m��|�w�P�s���osFú���|�:�-�3�ȟGOG�K��G�9W�^�˼#H ���W8�irn:,h<B>m	�Dx��(���7�gp�^Czk5md�ά�<�PG"^ ?7_��<�Ϟ�ً>\�T�:��ɞ�@�/f1j�M���U~b:|�	�d/,����w�E�M�u��u6qU�gÈ��ב/6���i;��Y᰼^@����b����f����^��Y�9�>�����j|Ak�9�L�6��[�:�F��=��O�.�6ə����༘=q�.Җ���u�J}4�4�3D�ݰ;1� x��������G���}����k̀�/�ʶsO����'�����QuN�:��>@��A��B���Z�p���>�CBah~V��t_P���;��,�A���f�tw]�0�TL�(����p��A)P�6�;'U�-\�˻��}���tO�k�7����+5�Ȭ�<�n�Jf(L�,�r�����X���a��y�G7!O,����T���Ag��"ڪv��#��|���ty9<�>k�s�;�8�mq�{�w3H��|��,�37�boR>�q��A�r��][��&k����{��Auޘ_�d��y���r6�(��*ʲ�g`�S��z�5�����0;N�� i/�[�{�u������B�~N&��V�K�#1�p��ߧMB̐��)��oܢ��t�'�A�-�!��ؒUQU�V"	�3���iB�5�\�mU�
	E��[����݄?>\C�Ԟ^�F�<�Ӽ��u��x������Wa>t�H]�c����3���o<�Nr�H��f��ݎ7�'��ڀA<B=��<�O�!�QDe�dbb�6'�+s�\UU��@I:�� ��!q=2��)m	��:B"����#6��γ�z|$�^���і ��DK�@ �������i�"B��)����upɼ�<&Z���CAx��TQ ��D�J�9�`�66�n�X��W�7.L��\�30ޅ�<3,/j;�7����?RI;����}��*ڠmt�\�s���mK�t��	Q���f��Uv��3N�E��u��Tji���\�^Y��4u6�64!�cF���-�@Q�k7���ɬ��+K��hRWV�vmB��#��CM]4�F�2��Xա��m��Z��}���s�hm�P{"�����+��M�S\��O�?
By�M!AgU����W�@���5�>	����yx���w3P9��
��� �彝t���ޟ	>���!ᬗ}��6C���gȂ�E���Aف�Ӗ���ɬ�$p2נr�4�p �ݫ7:z:��@ۏ2'���GMf�d�:���,�x���l�xd�%2k��4�ڀA�^:j��n��k1_f�=�;w�q|�#̉>f�m����ӱe��M��KfAlc4���b��&s�ʳ-_S����ͯ?5�6+"�gi�����;����}�#�f��/#���f*x.���ɜQ�����M�y]��H���9z�2�-u��ɖdd�l��M���� �܆p��>�v�;��M��o�y�5y�0s�	�ab�b@�����hEю��I���w�v�H�,�A�2�Q��کC�� �AV����EuN��<2�(O�kϜ��\����@�����Y�86�(gN�gV��p�gȍ>mzZ�
��N���A[Li�f�a?~x���)m��)k�eAs�,�|�s���/x���}��7��֑�^�d�A�>��,�.�0���cW�ڼ�*�oF��YByzZ�r� �tO�.�qk�";ibŜ%"����W6���w�����-�WT�]�]��Xxw;��!cv�l�#+���T.�bѭ؝j��� 	U]S������^N����<<����y����ϙ�ׅB�Ǻ��o;Y�v��,�F�q���t�!!Y<p�i�h0Y�4-�q�!q��+�:���9���g�c�w�������8_�N���3j�r�ޗ:f����c�5���4]�R�.�����!���{����t���ބ��}b��#r��aj�^�-�"���#P^3��{�=x���aA,�ly�}T##Jذ�mG��&�-�3�eSqM��Y�:7+(O/K^�^@�����Y]W�� �)0A���7�:�y'p^��táǳ+y;�eU���f����o�.��c{JÝ�f�]\}�^]��u7�a˺�>�x�( ��3�י�!�\u���Ҷ=����#��W�>�����9y��^����j��۽1��J�(��.�k��l6XP������@�t���<���z�^N�\7+(O!9���b��yx���1�%DGD��w�o�ne7���{/�{w�qw�;ş A��KL�⯟4%��;��א!��Б�*"S�V���F���;�dq���$�,�� %q�DY� ��� ϶��s5b�YByy� ��9p��^�F��o`@,��(����SV�wH��55�W��L]��ޏ3�F�6�Ϙ��8�!<Yr�9°��,ڊ�fM�+���꺆�ي�f�cջ�{�./f�Úd�2�ΨB�ùX�f�i�kG�(��[���-�Ϯ���)˙���>�ܹ�02��}fPY�)ͮ6:�Z��.n3r�!y�,�rn�Eҝ&L��N�va؍�d�J�D�C2��t�q�_R���]W�c�� nX���=G�;&�U��2b�D<n!�'���!�*9�W�gMu�λ�蘄O�YaI,:�Ckz�=�ٓA�6۹�MnL4	����g���������VC���+uZ��b��'�e�n�q�}CM�H�ft+������o�E�/OkU�@$�V7DU�m�9��璻n5�:�N���.�q*=�g'8�v(h��[�њ�-�d�Z5�*'Z�zkl�T)u":&P�QҮ�ǒ�ok�/E;4v�s+M�8�Khvn�j�F��o�f�C�lKY�S).���H�CX�_o[]��0��DqJW0Fmb9����BZ���V�������*M�:�f�9����'gzA\�Г����K����{~ܻ��L�ʍ)A��CG�r9,�`5r4���U�ֆ"fms8�b�1Ö��ng@����6�y�U�T�Z5F��Øt%�b�M5EDhv���DF"�%:�i5�\�-R�u72�<ڻ��Ud������iy.���Ѣ(�/6(;j퀈����5C�Q!CLL\�&bns����J
b���& ����4�w��c&��nˮ�a�5�\)h��6l����L��[�����#���]�\�I�5vDFYS4f���Z��lJ:	�.ͦ�Z<����&e6[��f��kL"���R��L�J�U��E�c`�T��j��3iS`^x"k��q��u��6못M/jʌ�[�J� y,;V�\�etF`�61�VQ
[6X��u�q��������Foߔ��X�Km���T�5��-�"�ֲ�	��c6��K���Ir1Qa�# ]i��Cc;V����$3B�fX�X�X�R�	l�׃�V�Z�+�A�9toP#p�f2h�����
�[jC-��P�t�#l�c��Y� �֭��\JK�Fe��0�@��V���Y�q�v�8���%�l�*�1Ke����E!�M]���4���f�i\K�����kaQ&j�F��p��l���m�p�]�ܖĉ��L7���-��L�fka�k]*%�b�hZ�WLM�;�U9ՠ.x�j��¤�Έ k5��:ƂR�,��u��wZ�c���4�AΚ��`�6��F��K.�),�R���)k�`���ʗ�`H�l�L�R൸��3V�]���hque��V<���S;��!�/
H]�mwqX3\o��<�yX;6�W4�쫘�.�TTiXͱ�������e�^ͳY�ź�Pp�X��X�4���m����Ll��Ӻc�4
����6��ehX �[R��)�5��X#�H���*Җ���l�.�́ԕlK���)l�$����hҴ,ۋt���v��,��X!��^�� �ݬ`�5k]r�%�-��
�5�n�����X�L5e��f��6�{���������n����Z9t�z��R�%&f�~�5��ב��'���t󽎳�VGz�Ҝ�zQ�� �	�1��L2�_�3��ڤ���df�VT�Of�\7+(O ���Ȇ�T�
�f_v�B㆑�,Z8J���+5�����Ԧ.�K�ş"4�[PAkȆ���={O�[�6�����n�k���s;udq��,mn���#O���'ş�-�}�af�@��s��c��e	���G/ C>mD�Z��U6P�%u55n%�[�K^;V8��*5�_��C�>~ndH ��d<�ټ���	| pze�g�y㔠^@��%�M�(�֢���i���̈́�x��"�tmN���a��=	�Qۮ����G�|��������̸�v�Y@�� ��$�a�Fb�	h"���w�n��3;��8n�P�@��x����^m�d"7`�}p !3W��o%1w_G��S�uܜ��D�A�^D4%���b"�(���*��.:��Q%�A΁�b/K0o`��%`S�S:ƈj��`�LlE]��j��|��z:���<���Lgv��;�t'��M��"�k�ח���q�@�YDF1�B�1���0l����*b���>@��ͦrLM?l]�H��"�k�^<�[ϻ��il�z�ֽ�ߟn%�YA��V��)���^ɾ�3:�z��,�qm�p�D,܋߀�s*�ܵ�y��:"�����ؾ1zs��Hg�K��[���9�wj�I[^��V]��T�����>n��^Uر
ۗ�W��L]����|�B-���2���t��T ��eJb���by�P�Ⓔ&b��� OԽ//��h@=����e���TG^����ǈ�^��l�� �>@�fթ�k�T����Iݫ�<�P#W�!�Rֆ�x�@�!	g͡%�N�ƶ����L�g#�n�7ހK>@�5y��k��^ۘ3c%b�A����� �u����v���,�$�����N�Q2vmJ�y�`����R����@8���@�WG:�f��l��`�ȁ��hVީ����gy�:�Lb����̘�r�e���V��N�e	�	mA|�gɸ������������=��U���n]U�" �fۈ�1A�K�D�{H��(_@�YK+�_N_l�w����,��>� �R�^D3�ԑ�F�g�y�#��ܶ���)u���82��^dG.3�`Ue��^�l�Zי�˺���2-fupΓ�YBx KjW�!��ЀY��y۹'�̍�ط������o���WFg��3"�wW��ͨ ��kv�g��� �um�ܥ�v����p��@�O�M�C�0�_%��f0��x�"���p�M�jnJK2O[}/�wK�h���g�s�P/9�Ԍ���d���W�f�{ ���ƍj�]�{"hG���z���55���5�+0��E�ͺ����L)kc(0�ѷ,9M��X�j�`B�۬:����fqec0�m�s�:[Lq��T��ll�-�M�2G*�J�YX9�[\�(8�,k��ϠoЍf����u��mM���Vj�Cm���ѿ� ���d/�Z��3����t(���8[�^����,��(��7mV�wH\oth,�'
�w�������� A�-��11���ğ/$#T�yח�BG���W�������泼c	�DQ7�K�ш�{�Ö��İ�r�����6��np�������s߇~c��7�~�;�=�ϑ؋�D��u&�Uu�z���c=�k�|4�e{�^����f =�P$Dʕ�KńV�En�خ"�c�0a%&g�f�z^D4�@n�����z��Q�^-�8�(�A��z���|�Ǚ�egsh��'�N���țZ(��F�>�ҏ�Y@��F������pvNh6�A�CE�mA���{��|�v��>��c�8}���Ю@�� A�Ȣj��uig�L{�	e[�2$�Y'j6pc��x��Nn3�n�7��]g�3��G/}翟|���t|�[B][����Y˪#�%�Eנ�D>�V-%"���.B8��b�~9�hʌ�۱q��;u<��\���׋pp"M]�{*$B�H��0&���1z����f�h
��3dQ�e!%�d�;����*�| kwYz"�i>}�z�^@�B-�!1\�f��M��w�\������8�(�7�̌}�T҈݈��-y�$�ޛ��A�EI�V��Z�����k��!�^?g����f
zJ3<�D���Ĺ�ŵ;v���4*���x��y�7�NUЯ����r�4�Bd�4�:�`�[� �R�w��_8Wp�ş"B����X����א!��j�"�[����32뫮+GY˺#���>ށ��%�潲b�lȍ�
����<Ś��J�\��,b#n��˲�毨��4!��~Yx��{�*2��n�e]
� �%�}\CͮD�(��bŇP�9畍ؽ�n��� �Aw;�{��+��I�8�iaWh�;k�kȈ>�Rg��6�ݍ�vu�n�Wiŗt|$�#y��A,��N��5e�i4�P-y�����1�t+��-�!c�㧂xu�Wt�aS94E�/�4-m`{ ��[ίp��s*o_m��9u�͜��y�@�9� =]��^�^dI�(��,����`��X:L���Օ�b��<ϑ�@��C^��ٝ1���tUb����ε0o�����(i1:�ݠeAs�=ý�=ޞ'y��������.�#�x���[Ӥ=�,��g�7*�����ꕄ^YSQ��ǣg*�>@�����^��N2"=�I�-Ǚ��C�I�m��mu�A��K>�@����p��z���ҥ�>�F�&�@)�m�V����B+�1�������1���|>	��m8l�"j�P������z2r���-�q���^-��액�t�����o\f��ƺ��n��D�T��޾��u�y�QT���*��e����N����(���{�ݷ7n��+vm�X�ՁAi�&��62�V^4�٘wXFkv�cf����\he��A���΍^6��,�0�K��+�a���o2��7jAh�YnưͶ��M�K�iQ���棴@+F&�X��uCJ�ZʭJک�qsm�;9����}6�_����.+��X�q����TM����>1��,�ۻ��*�E���U�J�bpY�FySX��qP�1���el_:���F\x����ᓕvG	g�zGg�a�x�� >���g���v��#k�OFNU�g�+�}����n<ȐDK��FF�w�o�s^�$��6.��o]p��C�>
��|(/� �1y CKͨ ���X�����ǎ�oU������'�;��D�	f�J+��¤Lu�lԒ�Ǝ�� c�X9�ՋA\�\�����>��/o/��*�/;�FNU�|��vE�R��k���͡�g�3���c�M0�����$���I&�1s�$l@j
�A��r'Z��fB�V�C�cN��!*�E�s_�xZ>��*�ﾹ��+�� �|�B�Т����V�+^DB@�6��א!���
o����[ENMUn]����#��Do!�� �����ɮ��R| Axը��b�����9Wa���	�J �ɾ>����D�2�-Ǚy����]�ݷ9\���|��E�5�=(ꭾ�����.Hl� 鸰*���Z��^�h��\e}Ϟ�����ϑ/7
yv�v�e�YC��so8X�q�F�X��&1kp®t5�b�5�>�O&�{Td�e��ڂ/ C�˧��n���!� B �����^b�)-�u��gx�홾�%�G�-��Y�����W�eЮ.>�>�K]�=�-�-��V�ь0��	�ᙛ����B\\m^q#�4e��:oU�iBR�&͢W^������;�x����в���s����}\��}���^J�Nʛ����u�uNq�]����������CM�Vf8�b�^�����&�$/R�1�����̝���v¹aq`��k�Ҡ�����%�fV�h�7Cs�ے��1VzZ���^��-:����t���q/w�Sإ#��ٻ|ܺ��-PC_bK`F�؊�ܕ%�۵��K�t�U�ηP[��jP6x�trr���h�r�-���{�����]X�&q����<7R�HJgV��9��S�({^�"�Ff�����n�Fa�s{1,�^����C-t���9J�&��^ڋU���9�9�T�0^8VH�S�si<���!+��$(>�1�׏.��XfcGV6����N;�b��Z�W
�m�؀_�ꆳ� j�i��� s��o������?mSTQ[b"���C��/�US%CT�PD���_ �D����e�Ѩb ���˗ �������JqDR��QLPPP�PDTCA�LU<�J�����*j���d����"����mMQs�j�lTr�UQ�2�$D�@D�QQI�(��Q�35W�&�<��kF��1t٠&b9b*�ӊ��-�F(��� N�[��v�מ�Z���e	� [^������At����^3�n_a��� qd�y��4�6(����Y� ��-�u���$5�[����#1�X|�񦠃���G��\wGQ��/�f���5���i62���Ɔ#�V��Ms��'��A�Ty� ��[Wy�7��]�u��a��PAk��E�=���~}Y� �uo;o��U��>g��� ���n=;yaeV�>@���z��<��i��Ӽuj�)�z�u��}a�����ɶ'H�C
E��D#�PsW�7�\hp,���"Iܣ���rU�.Y̽�5�ך�����������3UG���/D�t�{J�X����/�z��+���ϛLC^@��k�M�XP�j���;�^Y���7�G�!K*k!P�|'�D ��K�s#!R���r��+�un6`�͚�#����~��ʐZ�ت�޾�Ǐ2�pJ���Y��9xT/��g�s+6��0�����EY���Х�w�,�4���nz����	y5�� �בyx�v�s�]pw^���7�ydp>ex�� ����s�s2��/*��PG)z<זEe�u�^V<�|�p ��^g,���x��YAgɸYV�ֽ�U,n���
k�}�i�k��m�@:&Q��Q�QE�:�rK$����=[W!����}Y)��ל�o�S��su�k���3���J@�I����XL���������5��m�v���g-FQ-�f��p.1��dv*��Lf�Ll��j�W�G�o/_8c)|�kB�Y�bF�V�3ɨ↡ti6A(,#���8$e1��FC8�0m�b�,]��~����~���EQ�2߹&<��-��LR�@ʂ�X~�x�/|}$4�q涹�ٝ��,�!�Y�6v̐k��D�2�!��>D[���(�P>��.)�f�>˷�B� M5����c�ȝqsf3��� I-�����.�nݝ���v�'�#W�RAx8B��쭣��#W��^-ǋ�έ��7��d�X&2L�\�F�%3�D�-i�P#1E8�g/.c���������뮻y�_y5���CK�7�
-ǎi	Q�@������<d�����1�.�h�P�fg$��C�Y��Y͊Ӝw�B��T���� ��!�׷�3Bƺ�htW��$�>���Z(`�k����aq��Sq�����6*u�c"?�O��A{��)�oW�a̬�#�&���,����2����i�P�(����ᶯ����0�u��]��GMA|�iy� @�;������A��y5�8�_��Y����&:
�g�A|�i��!��[�/�z��@c���ÙY�G	��F�Y�Y�Z�=�_^�_�4npF�Y�f�0ej��#R]��6��Z]�O7�G��i[PAyz���u��U��E�Rq��.:�L%�ᐼCq�@�ϡK|z{���(t�'J��Ӝw����Y������"������G�-x<]%�;K_C@��:���wOd� ��z5+�Kn�
�g^@%lY�or�(*�#ӞO�}U�S�=��2���h�o@�Y�Y�hwoE��+h����w) ���Os6����e� |m�0�JY�R�dR�fG�|� �dl�]�7=�l���Z��A����w�:�-�3������=B�l�t�p�\��-�˝�|?~b��܈�'��4�V���a˼�#�틩��=5;'6݋ҙ��c,1�)s�^�x�:��d���Y���n��X�^ƣ�q�!����IeP���q!�>A�  Y�(T�]_*��Kkx�pt>jŵ�kȆ�̝�]�����͠K��՗�s/2��M@�Y�̈́`�d�wr�CgI"/	Ԭ.i�ѣr�T�<.o������%��t�">3��I���*ڷ3k��Wm��5o2ş\�#��!����pv+��䤠L̐T��2$l�B9�-֘�4v�,2ƬL���.��K+ʶ���ħ��+���i�����^%�뮣[n�Dbz����y�32�,�>��#y>D�������~w�"�{��OiZ�gj^�f�m��̱|��@ ��p�q�D���:�l�V�D�iK)V�b啽8��Y���u�5-9k�}$2my�x�"W��L�Z�8fe�Y�g��B "�="��'d^�u�)sH����a���+���4pI��݃j��m%��P7
��=2\����,M�<l͢�5�T����5X�ю�����CE��tZV�B[55��Mb��fevX�zf%�ѼjE�;g3]E�٠˘�IW6�,�Tfn�у��c\عͤ����A�t���Wl�P���L���Y��ns��7J�E������[�
[��$kWu��eUn-q���V
䈕3bq���^my�r��՝�o2Ɠ��l���Z���C6��b�0�hE@��6��� ��,�Üq�AN��3��m<�4�.��F/ A�PAx3���n3+z��^e�Y&� �� B ����+�;�Z} �1�Ak؝wmwm���b�/N/���*�����7�p���Qa��f�\FG��t/��݂���h�}�/���F�E��$�r�8�.�E��3o���|�5f��ma�K=���'_<e������w��dp!v���nϣ2x�Q� ���/0��j8
}p�l������zf�2fedhw�Q��n��[ؖ��ګv�j]<0g,�O< �>��P:����}��Y�y�/�>3��}$5V�7�Ϙ[� �>MǙK!gQ����y�S�u����-�@x8^c.����D^^#�n/���/���� p6Q{�Q*t �N��|�-y�rT�]���u����m��ٷy�,�-q|����|�}Ժ��RWM�'�֋��h�V��IB��s37'�͐r�@,�|��ӽ��t�]!��q���5���2mG��X���zB}Y�[|�ff<�刾����//K�7�Lr����
�C>mI�"�w	������RK�{��awY��$���~յ����u\/�ΒL}p���,=�]ZG�#D}��{9�����fX���qA��gɸd��s:.^v	�$�̐K(+�9�3��CB�D/wJb��0m� � 8-z <�9錀Me�ues���,� �eF�!�A,�_7�~�=ya�֔˭�冱���c�Ia�L�e��K���l��^-�Y�W�׵��,_ v��ёJ�9JC"���Ϗ����W����Q��;;�����A�E8��!�Q'�D�א&�A�!�7EΊ{js;n�����{��Q�A�|����r"d�D��U� ��D��u�p�����A�wÏD.�JP�*�;1YG*dT��F����'V_ʵgN���!S��HbӒ�q)�f%|��>R���	gɸC:*�y)}B����vgʸL��E���k�ds���O/���l(��m��`L�5�����hUsB�s�������A�/�@K*�:�����x�wr��˕ː}ŔCq 2���� 0��D�����wY�/�'��!�#2�E����qQ�6�D·�xoh>Tf�5W���;�Q^mH ��D4��9N��I�^^!��WOvWE���d
<��hq�͎�����p��2y�<��OyҀ0B�w���z��e#���q�|����,�+j2=NI��RR�0�s������CD��n�oU�����J�F���f��%]J#��v����4~��٦(�g7v��=@!8�����\j/� ��EAɗc�F��F��2m��;�n1>�)oj���,C��m���f��Qf�v	�����C�;{/{0����z���A���nga��[V�	�����`�z�X�\�7�X.�mAϴ��W�ϻ��-;f%���߳��?do�[��>=Z�'^:u�-iw�]��+�.�^Q��ڠ�1��śrA/�(����ψ�*o�)�����S�w[�`�Cn�bޕ�B�@v�ۛ�D��0Y��ł���}�Cu�ٹ]-mmoQ�!1O��Vh��O>R�U����;,euғ4�G^�xBnV�}{�.�W]\�7P����PVwMʴ�-^�~%/ձ{M0�L�|.�=q��jѺ��G�4$Y����A�z�ߎAJ��;�{ݶ�Zv;0#ݮ��i�yܩve�4�WX'P��;,CB��R���ܣ�Š� ��I'�����)�����Q[b � )��j��xq��"�tF�h��4b"� �֝G'\�4S؊-�TF�T�	�\ژӪh��ICU��Ո�#���㦊�����혢�	�)"�(9�LD�Rh5ٞmEs:k��0Tm�&�*)��LTT��h������5T֝U�CMSW1��Tv�)�3���&�Z"b(�����i)�ۛNة)�����~01v�:�^ʄM�b�̎Yy�\7D]s���LQY�\�`0��6�6���+o]�^Ύ�V#t9���J��lR�2�n4V�r�h�,�+�����Û�͒�"�h�Z=��G�e%+-1�e-WG��ܡ������sR��il�0�íp6 �6ճks,4��B�u�-I[]n��0Tp�(���T@�.�+H�i�����-(PdT���2B�8���s�,W�k\I��ř̼dͧT[��c3U,1uŉ@��F�k����i��d�ci�Z2�kk�ct���j�<-*�4�a��H��1lԸ��%�kGS(�ˬ�ͣ��KbM+�-rYz�,ݫDu��t4&V�m�`:��U��7VٓPh:��M �3�a�,W]f�!h�e�7���p�\��F�F�ֆDN��^�b�<;�R�e�6�%�H!)4FgUׁ������
�Hƅ�z�k�����B���eMYi)�9!e��p���
Sv��0w<�Zf8�Zm��4L7!�]w��h�)؍��E5Vcd#�kM̱�ҝ���fJ�:�!����0Y��2n9�E�.j2�ZÐ,ЇK�4�4Vl\��j-"v��ZA��p�i��١��MV�cWk J��S0��V�s�Ŋ�U�Wfm�ݱ��s�d^Վ��P˕k+*c��^FhG!Ck*!SvZP�Y��.%-���lRa���F�Vm4s}:W��VZ+�A�q�#y�\���'^�3�;@��y��.���h����.�����n�U�Ύm4�\��8S�0IMY�.4EH� .YM�i��x�f��)�34e���)Z��T�u	Y���n��o8����6�:�Mv�������W-+6��򘴬m�$��ez�v�2b�bf�� �(��d	,�v{w�u����0�3��������$ב AmG��YMy,�
��VOnWA��ޓ�G-���	�/[��æ[4\t�-j�Gqp(ԹWld���j�,a59x8�7dI��:}��P0 �#�WC�����Ĵ��Gȍq�yb��!��k�YTM��=@W���̞ݮ�y����>�BHeK48BIp�za��+V�V�De�ʳW��˘��6j��ߺ�KO���zK#U;�睷qY�3�& E@��@q�>M���!U���V�������+��S�^���W��o���r��ݲ�mU�ow7v�u�K���+s�p>#Fu��c�{���k�k��J9Q���^7�#�1zK 8͡��uE��$�]�v��y���@4}����P>e����P�($ ^/@,�T��{�n�̱�p-� �j�4{��gծ g�Y@�����b\:�>E�^��U�e��(����j���߯�x��V�Ʀ�#�kv�VR���獌��7��	] 
glB��7K�p�CK͡]U�ݳ+2�Y�a܍�c�P �3�� d,�R/��ڢ	�ا����w/2�ŵx�ۺ���1�<F�#�|�2�|�{Pݑ7�YQ����a��lfP@�T�Z�-��A��uL�  �$�\��e�A�ls0���~ ��ݩ�d;�"�P@������i�Ĺ�b�	�>��B躸��<+2�����?n�Ͼ�#�<�y����A�V�=��"&*��{�l[̡�%�����g͡�	����\��Dc^�6WJ`�Kb�i�Zf�n�B��r��I?D�혞��Ln��'�e��WW'Ï��Ay���*�+O1��E������n��Y��Gx�h�ށ���Wz/(�F���	h"ڂ^������V�(a[PA�/ C^^m��}�Sq&�91� O�+�wv���!����F\��\���f+�7�l�P����kvt#���eب��]�Ce8��rV����չ���Fk�׃��3>�@�FR�qN�̼�8����>�aQh�5q(�i���:��*�j
ⱶp��#u֋�?'�>q?�ʐ,�Q]Y����SB�"���e{{�c�8q�-y?O}���N	�W����;;Gk��v�D"kDe�ouo��Z���Y��h[���a�-�]اEf^
=��(���X��|��.{���q�����]Z�w�S��,� �Q�/"�ED�Ջ&E�B&1bɆ�<�[7�@�Y;�F���D;� �(�����Z��O���	G?$��qCA��/�4/�<qX��A�s>���%�{�^�;$�����<n~�p��Ywx+&�є��	(Sb&��^�0R�F�m���˩*���)*�[xm��%bF�G:�[]s�(��:"�Pt��
Efye�3LL[m�kr- J����hrFe���4�źY�ݱPme�f��1]�\�J�-�v������ֳ1Jj�bq5j	��F�W���0�v�~K� A�@QC>m	2j�v��Y����Њ�q'�:�dAg�Ȁ|C!x�<��M��!QYX�v����/�&��� 3�qǅ̿r�;��E�	���3�;�`�P�ָ���}��m�y��
=�D~�^y�^A�EΊ��+�S�,�E��[�
�j�v��Y���4|�rq���GH>:P6�dI��i㜚�272R� �	��b�����Y�MA��CKŸZu���̀�%)D��*TL�8�nTjm�c�\�!�m1��Y�A4|��@2��(l1y�c��TC��f5�QD���@2$�B�u�"�Z9���+pk�n���qYd�	�Pd��V�^K*ვ��܋�%m��*�0�25�D|F���!}�V��S���G���F�C9�+c}с���t� �D2-���&���+;y]��N�س�+�<���Ad�ѓ�����Y2����i��	Q�Ə�]N�=~T��-x8�Z�c�Q��� �G��+2�h�F���DͦnG��>�e�5��8I��5LG"�)��3(�s4�ÍWgz���@&ϑ|�����W\��g'yl_!χ���V��J��*3��]'3vӷ�iM	���+a�,��*�=GԜf1Yy����X��Cl�+3(L%��>1c��/"rLMTt�q�9Y��=�������H�6����zVd�S��s�w�G�����e�e�Q�  Y�s�Ҩ�׷g��� ����Ś�'b�r֨"nɖnq���\�,͛͋8JDp�cY�:уFb4.�i���c3BVE_@>4|4���g�����\Y䎘F@12�k�j^��<���d63-�13$/�&�z�^�n����|��^VQE�����hA��(��,�G�`��Qs�s��>���d��E�
Ё�5yx����M�m���Z7Jf���#�����y�m�`����	Yk���#P@��yT-m�7�Y5�CK�7 ����yYDp ��!�0m�:Iq��Z��������z��6�S���/2^!�E���][+qS�L��U�a�Y|;�+9:;B����8aX��b����g&j�Y�f�>Y�y�/�'�r�!��Cp3�sW[��#qG�A2�� ���F��3k�EHYL�;m䓤l���x��������v��T�2��Ȣ�ƭ Ȓ�jA=�"�� a�bU��؎yX(� �P ��C;+�N;���F�C!�k�"�zՏ6����y�,�W�"#�Ra�c3��r�l֨ؔ@f���]��.��0br��lz�h �D"^m@>d/�_�1=V��N��َ�yX(� �|��A��F\�޳z�2�) ���Ъ��f��3WPϚU���M�f�2[��ڴ�&�/5�;7>��6/���:O����C�,�I��ձׇi��P�KD�n��)����M-ٛ
���8%[����Tжݠ��Zm���u�ëF�M�c
�h)�J%���S���J�B�:�(�v�L�q�ci�T,GFQ�a����p�6�Vi� ��.Ev�c�`��Ͽv.�iTЧE�R*Q+*a�c�.n���"�g�I�g��;��[唫��5��U���C���؀�/�b^>��@��϶�g9�Y�Hw�j𥽼�.����[\��<�#y{- ȟ^-�}	�OuE�u*읜W���|YDo ��|��aO40� ��PA��++65��U�ő���9��C�,��^�Be�Q�f�U�M��^f�u����.� �!�/�2.�Nb"jC(��MZ1�����������]sڐ�.aB������z�q���h@Y���9�⼬{�T�3���	�.�Mb���hLb�!�������/}�4l��<�;j^X��aՃ�C���â� r�$��ִ������8>�z��}_}�����5 �x��.�riߌLaDY�h@��%�9���ݚ�.��E��j� 8]�V�f�Z�Y@���hB�7��ӊ��Q�|�"*��k�Xr/��>F��� �C^m<���V3,id/l_e�k;�G1�#�q�8�4�p"���Mm㢷 �] �����*�M�����Tmh�g1�Vz=���HO��d�etV^A[��+"�ю\�7�8� sAd"BוR�F������z�H�1/���M����YX(��>�BAҋ����K;E(�q Q��ړ�E��q�#,�'�U\��bIS�(qx0�v�֫�{vo��-6ፅ{�Jz�o���TcEگ^^�U�:�4�ghjTv]a"���0LT�CgpкYD�;\�a:��5���0�՚~6�Ӝu.�{k�
!�����-��㎄n�7)i}z��6��˯�[��Z���vɚK� ��[�ֳ����H'���͕I���l&[�����6U���mC-�4����k#��c�U�I�s�hr�.����k�X��#q0"5���w.�ʜ��Z�v��x��bm�fZ[��ӭ����v��>��U��X�hۆ�Փk�;tWN�N�%�,F���]}�n�LRO	����57i�ټ��HK�9�g�t�\Xw�.5�7��7�
����MI��osk+N8Tb��E�5mFLgj�8"ޔl[��5���90����e��Z&TS�r����I�����u`V���;��Gc�7]���޹���u�#�#��b�wN���X���`��N��M�lړ.���V��r��������x������̛Χ_W0����{��D5���DܳU�_1��)����hh"j�mM%PU1��(��9�DQD�%�h����Φ�b���)���&�E<�W6b*"bj�j"&*J�5��&��"b�h�v��P[<�8HDsJh9�����J�������
)�i�!AI��UJP�E1��y8�&���M=��r&�"��C��v�E@@��5�yna���{��E�( � 8^>n^#��yI�>�̟3U|ewgVE_@ �!x��7��b�)��ȸJB8�Y8@�t��0g��z(��ΌO+ �|��G�eK;ױ�y�ȈH*��S�Й"�G+���ʭ�:gFl756\��߳@��H}���.���]oF���s�^���$��Y���&�DY�nϐ,�?f]U,�!�#�j6��������H�PE����,�H Nb�� 3��H�;޵ۅuft�NV
<>,�9	�Ћ����-��];Ȧ��C�ՙ�C���cY��9�Yq�DH��5/�p4/s�y�`\��VdcQ���pצ�4�z|! E�u�S�A�q��!g���*g�,�T�1�bثb���=�g퉱r~��
���Hn<�������P��/Ҟ�M.-�)��E&?��y�3+�Iq�mv6Uߓ���L�;�����ܙ���]yә�}�5#͸m/l��U�ud�m�Uջ��Q̾%��MM��j��h��k�{��r{�sŏ��$�Ԯ�|b����j�-�]|Wo����>��'�تw� ��t�'Ƽn.�e�l�P�s��i�In�F�<-���4�����ʋ�Mέ����ʹDV]����[���'MŦ�� ]E\�����I��.!�ЋM���b�Fݨ�u��pU���ؠIHQ�@�����Kp8a:XrF���r��Z�M�f�* ��Yp��G<���d*s0���LK�pm	l
4�V��X'.��]6Ji�����n
3K���\�U#[v�E?_~_�����#F�S��4vb(i����5e!]n�W��ɤ<nC9QCzN�tUy4���2*��"m�ǛK�+y5&����u����vLee����N�T��^m���A�ԧ&��\gm,�앜��mяtb���b�#*(vI���-q���i�:���۔7�u�4ثh�f,��ޏ5�����%���+��홙�� dhL��%��M����+D�P���q���=Gͯ6�J�o6\oi���s���:6kv1{Hmy�#�k,�zF�8��D�}��}�/���u�Bb�-|�"l����u����]��,���~�Ƽ��;���tU|�� 6����!ꜷ��pqo�F��ů��g����U�Fr�2ٓ{q�j��>�!�M�Y��sg�HnM��zfc���k̆�{U*g\8'/d�oAUW�Z����<�����������c͛�n^̬k�����X@t����=w���=_<-U�L��=q��њ�LH�<�je�J�7�Ӛ��wUn�최6�/��C�"��.f�ZB�,�}��֐�Σ-ߖ�W]ܹY�\�W�d��.$9Bd� �)VH�9Y �m��i1ʔ������*��~���Gi�O;�'V�׎=�=�z��G7,^9�޸�im6�m��9���fGF��t��6�/���S>m�7���/`�0`D%2�Ab2���d�L65����[�(��-x2:��d��M9�<��~��V�ϾIg�����t��<F����Z��Y�2s}��וG+z�='��2m��T�&�z:��kx��_d�3�g͠��E^W������y'GoU}�ð��"r7/���UZ�����t�4;z�t�Ȝ��y���lm�/��p�vM��;��$�����Oxm�B�y�'��lc��3�\�jO<��g��=|���Wj�P"۲���ѣ���L��p���w��ͯ6�U�nˎ�y|3bcW����s�lZG���N!�U:N�ޫnz��J��9������A]%�<#]f�h���]�8]��[R:�^�����vu�qܬ�*8���-��t$�&�n l!ێ��.������K��w��������B��<�f��q��q۞�1�c��� �莢N��b/�)U�:����r&�wx0]a��j-z������B�1`IQ�Bgb��i��jԌE�
.+�h]�,�3Ukem��k��b�*�3��%Pk����1�o-�(	XÜX��1+3��4H�c��VZ�UQ\1#7a��
m�f�,2;$�Kp�4�����{��H���0.e.�5߯<���SCBjTt1\���ԃ��u�У~�[�	e1s�9f��m��Y�lF���6/;^��ە���C��oM�J�d���ې�W�/�\.����N�6�������9��)�;�k��k��b����&�_UZ��-�!�س��V�U3���c�nV_���u�7b��L T�!4��.����eL�"]r� ��J������B����N�j�yLՠ�gͯX�1�%Z莏Z}�� {�Ժ��-���ػ�=N�FʍˍX����:�būz��Uj9�}O.z����t�7��p�GtB��}1�wk/�J�L��ڪ5Xz�/�#G�����R�95��S�ם���7W����m>;�T��9����^�����|�@0޷��c%(�Q0�BE�,M1��)�3��4�_J�	����x����n�2w6�F����K��u�w���H����l��dv�C��5=I
�`1�pNte7Q
e��m��v\F�f�%�"��PinP��Cfnn�gb�|*;`���n��/\ɑ�YW%�1V�s0�U���<i�S�*W�B���!u������M�S����ݻ&y�exf��7�#�Ci�R��75q";���w%N���6�ݥ=G�0�%���
2R;h��k�f�@f�
]��{�I�6��V7c����gyz����mc۰�T��W�2sZ?j���}�۳}�w�%*�女U�>l6�،Ů}�����P�W@�l|�X�j$r��ؘ�~��Z��?t�u����a p#Uw�[&tu(k���Q0�A(��VPY���"6�{�\N۬:�5�L�WӃa��o�b�H�����~^��gǻvo�
��lSh��5�n�_n@*2T@�3
`�L�Q%��YX�0��*�L�3=��UHz�����w$�����B^Ul��h�,�6�L_=n��ܞ���;�����\���&�k�+<>�
m�M��z�=�0�s�����7�r]��ͶFy\��H؏v�����I��ڗ�{sO+�R�UK�U[U{Δ�*\ oxݞ����9��6ﾪ���,�sݿ.�dgq�:����K�t�+��M�ܾ��$F�ܘ2hi��v��Aj��"�b��.�rȻʹ�C ޗ����,4��hC� ��n@겥cY��l7�	�9}��L��Ts(Wb_jc3���u�[����v :b�5
�qf�oa�3�)��&�ڻ�
��3�e�׮�7��3]ƃ��b�$�݁" e�g7ܼ̈́�]�>��+6�d���C��Jnie�7F�B�K|4M��pl��{X���Q��Qvv	j������	n�V7�/�x^�}�CJ�p����z�^�)=�u]ۉ���0��k�ib���N._��.��Ӑ���Fޅ�5P�e]����<Wp���P�v���Nf�)�ǳl˛f��צ`�5��J�\��ސJ5�C ��s�V��o�1�7���
�G;F��K]���MpG.�=ܓ�[Y,����tF��y�?�sb�geM�sQ�C��QY7�:L���앯���ND�z�Ÿ�ulq�Lj_]��ux�y��1��}f2�Xȇ��C��{���uY�#N�`��"�FdΗ2p�ư�W(EQ4!獉"����0��t�q�@w;�<�^C����h��������;�r@�j���y&�W���:옚��1���m>IO'�h]��`�<��s����4�141U�ꊉ�O9�,Q�#��E��
t<�IG$�0�U�vtP�b�孱E<�۲��F��h9���(�XJF%�*!]�1%%4PwYu�{j�]�ĥ$UH�r�F���b����A�5AMTT��<�E5��jXa�SS��ߑY[���gVE�d�଩H�9�9ol��gL���WA����f�b��mb+MQ���e�B�U�B[�6hL�t���1A&(q�ttM4.�-�@�&Q��5�)��n�b�H��H�+ٷ�����v&����JA���u�(,�ًv*D�������3�嶥�fYX��k���]r�j�e�{bZ�*���,Œ�GC�0��S���h���"�RK��[�\��̣b��M�6@X�mZfDv�*�]x+kfv�`���-���FA���.�%ku�Hܕ��NhZ(�K��ґ۶��%��rM��׮��Gb����q44.@��R����y��s\�c1�VXZX#���I2�{uC����!��a��sY����T"�f���	v9ĺ��_,2���r�֌j"�$���؂G`��Ŷ�)Jk���qp�d	�eң��5��m*�TCm@�e�)��%(��Д����GTv�U�������i�F��2k��	�a��o�M3CkPA)1m�#�u���#{iu瀆L<�N�:�.�RP�̻e˥fc�˴�,.J�&���ȹ%涕��	�-,��^00hS`�s4��h��u�B�G�]���2��v�s1�V�p]+��Er�d�3-���s�XiZ�R�v\邎]�\ܶ&]Sf�l��M��.��3�̹%ֹ�`#�"�f2֊���C#Wa���.��#�@L�J�Շ7����c,�f&,C\��\�Y��Jh����	g�O#-t�qέ�Bm[5�qqn+��.,͕X*J��f\,�C��V�m.6���guu3e��� {F`��&�(�u�1������_��M�n����8,�f�A����N�½9��6=��y���������O�F>4����cO�`�M�|�'r��*���⛸�j��z�k��G�m��:�m�_��D�Ԙ�x6)���e�XS-�ǫ��a��پ��.��gsܵ�͏�̡X��B�0��k��n�K^�^�US�)��o���/�xD��jeX��y���Ԏ\�0j: �\鏾Z�}U>H�Y���|��g�U�QU-��PK�HU_!���ތ�N�����e�"��~��hF������o��`;��H̷��|���>�w��������k��UX��W9��2�l|�W��K���t9�	OW��4���l����~���ؾr�՛�O��LTe7z��������ոo�2�}��=���ݳ}�o�?Sy�����%�>���؆Y�ZA�]#c0�[��w1be���uU~y+��͖ƽ��9�W�P��zA�\e��S`K��̽��N��{37ޜsT�&*x7���[?.�|�l|�F���Q9Ș�r�Q
w�x����Iz��6��r�ܦ�ې�E:���g��cκ��n��0��w�����o�����9�����(g�F�lT{[�<Op�����������@n��T��^�ff��^赻��ޞ9�o�O
l|��ϩ��������A�3	4�k,Z��5t)���W;���{���c��;�}��{f����J�>Gן-�Sb�7��
�\x�ßV�O�W�S�X���!Y$4�lSc��}�/{7Ζ���d��NT�&*y��m��̪���=���ol�W!�e3(�U�E̪�b����'p��ln�v8����&�m��(݌>���a��s�6�EzR�G��&��W�Sō��M���R���6���62p�b����cm���o0���y�p��
�n���:=��E��7����=8gT���ER���=�&b�x��{>���
��}�]x��܁��R�@Ud)D��^�Ι�:�����ئ�a��2�W k�wŧ]�<=�~Qn��������`��͆�v��'����{�W%��5�}�l�ݖ��x7���h`z@1>�׳u��s�%ND��8^�+K]av!�T�o�e�ۘ|��^D��.��f����e��k���j6�C,uL1��G���fK�V�(��gY�	m�Xݣ,1n]��aب��,���Vhг�R��mڸ/cu6�*�LJ[X+M	���4�[�:m���ClcK4�gkmу2�r�ܗVh�U��z��Co��S(�[���MTX��"��S;\ˊ�c�_|�w�^��;�Swް{(M:�o�F�c�ol��֜3�r����x{�����h_*��c�"��r�]�
�T�V{HQ�ʮ��o��ܼ�[[ʩz�6>�/�+wN�MΗ���{��)�,!q��.�|�
���Sb��mC�����׭o3Տ3��_*����p&Cj�(�s�4�CXp7@�WGc7f�j��ߩ���עF��j��\�ol��Lcǜ�{���hm��cy�#��]��V{M�k��MetcU�j��ٙ(+�G��:㼖�V^g�9��S�ټ��K��˅o��d�=� ��ꭍ�8�� 0QC�T�R�ctl��u�_3Տ3���l}M�«y�ãH}���y���~^K���UD'\�$�v�TBF�͏��=��r]=�e����Kj�_xn*�Y�������~��	Ws15�2\o�3����ڝ�+���ϯ�����U!T���ۮ;���yI�j}���5M�+�[��+_��~���wm�w�m����%Y���T��Wf��9nt��D\�&���U�$e �tY;6{D��x-Љ�4Ĩ������x
�qf]����9��lUv�l6)�w�Bu�S����jA���=S}J�s�{�u���*�6��ש��['*}݉v�.�4{�=�B���UL՘S�{3 �*LyJ3�@���^��#.�f.5v��h�I9Σ>l�+v^����'8������:hv��b���z�v��Ґw�缯����AS�����"&�l6>mzt�n�{�h�t{����n�+#6�V��e
�R쳜nzw�-y}�ad�CJ_��aKU��\�y��u^v�I��nTn
�U�f����Nq�'Oe��#P��DT�顱�b�o��-�r�P9C{�#���y��k��U*���������U�h�����*�tҊ�1f:�8���D+����ϳ��l�6)M����0�tZ�tL�)z�������Doy]ޝ=gOt�{뷾~�9k�&+tS{^��+���KI>��l���<ZЭ��gyv=[�������a����S�$���+����v��w�.�C�=ELY��h��!h�l�b��M��,5}g8�ή��p�̪�U`xI݈W��ʧ���}���u�V�)q3q�X�{2�[���T",��\���ٓ��}k�~|f�nt�
.x�0ږ ]�� ��4)�YL���5��sæإzf�f8�a��4�V��
��B͉�����2�K�^F�N��CV���dؗ6Һ)�B�1��[�P�bh��wif�F(��5e�]6!A�}�����tјvq����9��(�M� 71j0����cm��[��;���n�����/�����c��b�W�c������������l]�o��y��]����M��m�`X��\On�kZ�:^�UK�K�HI�a�ҹr�j������.ǫt�us��l�K3������a��{p�u�}�Y]�=��v��m�*�Y� _]R����SүaQ`�������aDF"7DڻUHU,�9��>�5���\�c�����a�HEY7ht'���F���ev�^�Af��{�.�P�8b@g�O<�R����f��C��2l�Bױ�74�֝B���Cx]��ӯ��c��:����Mp��A`�+���͆�1�����fwv����3����Sc��~�|���T�uM��<��r��&>ͧ���+tl�e��q���'�_nu���z�|����n���)�u'��X���~ �832���&�#���v�e��'9��ͳ�b�Og=���7�]�yOJ��
�)��a�{��0|��T��7�ރ�~�1���x�=��+���������k멨ϣ�� ��e�3`�^3Y�ڗZM�j��c^��P�m�r��p�ׄ&#N�qŦ����gw�7�����E.;��Y��>͡p]�6;Xxu���%��T 纥�G0X=�oqM�H�����pPO3�b���,�ݕ���IY��Ȗ|��G\߶S�*ۤU�v�}��B�6�������ò�
3�s�2sD!�{��l�{p#`�h��H5zJ�b�ܽ5Y���+a7���L�/�n%�~�39)/h�Y�L��������)���*p7w�;ww[��t�;��7��q��F�e0`K�F@�p��q��,nܦGZ/M�^��>���); �Z>�T�]����j�f�*{;h���QV� �Q4��QIB.A�s�^V�1n�B���l*�*W���Nǌ Df"��0 V�7X�2
���E+N�}���ɎA/s:5��)�=�QÚlN�r,�̫�J�j��'��ֻ!���Jr�)ɹ�4�c[akV'Y��c�w��_T��Ĝ�������뮈����^�FD���9*h�{B"�wuf�]�7���g�K�}W��؀�I䜋aq1	�t���;�4i(���@P�&�F�˯-R�d��yrW9�iG���@r-/#����M&���yULv	88)�d��N#�G,KA�`�i�;ذkn�^�S�HO"�9b<��l>C�d�f����0�<��@k��i9U��F�)�sX.j[s���s<�� $�yx�<�RH؃�-p㻴�ع��r��u�vNCʃ^wRvO7y��>\��H^d�(+x��w�I��J���<��R�	^AI�9¹P��BkI�9y�9�syq���y�N�I�uH]�v1E�����v��IMPwj�d���������qz�|�����f�.Gv���v >�Gͅ�w���ۓ�]�u>zsފ�ow�6*�����m�ݦ��+��:{�k�����T�Tf��|�Q��L����F����ͷ
�^P%D��D����ᖽ\�R�R5�-���/^�#�c�:s�M�j�_mr�f�L�|��9՝���o{��Ű�a��'V����b�ȩ�:�V��=�9G�1�63�vT�4Zj��������ջ�1[�7V�3/�X����B�>�R3ެ�ھE�&�d��sY�2����Bs���gJ�hޅ�{�ll�b��M��������n�������.���m�H���s{��m����ѕ�R&�وK���G0�$�}U��[n��Ƭ�W��gwV�	)�7P�B�z� WNu�wO�u��^�o�{�Gz<z�z��ޱ���(����a�ڥ]3_=���s~����z!_o�4ئ�w�Ol�ќ�j���ƫ�W��UQr��]���l6)�M��3Ʈ��G���G�V�}I��
l6����|���pX�y�@��V��&�6f���M�m��ٽ}$s@�l���:�Wp�^�>�
l��j3:ǝ��a�i��o&	��VA�]�CYa����d�P	��X�VS��)���6:+�6�F��&�.���Fғ�2F�v���T*Ӭ؋5e�.[-��(ģ�x\$6
�]���.�.,p+SY� �#e7{��>}��k�ґ�	��,��+�R����^+?|�|��؎^��{=�:E��s��Mg�>�l66G>�Bc`��}�7�>�~����Ч�3���sf���^�*s{y���ũ�Rc�*����Q�����Z��Knƾ���ڷ��c8��1��y��ꩪB�
����xq��dtgt�w\*�b�B���x�ʥ;5p	�2ba�B Tٙ�K�j8�V%��J�̼I�¼�b��Vo�w�GT���w1�D+t|���M���Z{�� m�r��֊� ���ٍ�S�Q���w���/�n�V��r%����V�,��T��T��/{��9�ި�o�G���g������lK�6s>K}wo(>ك٭v�	ɿSb������]�u���?7O�s}���:d�&=��+NO|�M����l7�WF����B��{�����}Q
�
���p�ؗb�Ҥ�Դ�B� ��F�T�0U�Fa��	$�6I:g��6�w	�����~�ش�H�5o��o��6�o�9�VH���oڳ{{�Zd�&>�
o����Yc�Bpl6�b���= �3|	�p]�Јa����<�W{�q��+>C}�!p�[m�ha��qf2lq���GVnA���}��l|�"���#����7������&�M�(\���#P|���T�m�-���U��v��䎙=T������g���|����h���d�mTږ�p�U��,f(�c7\�o�6�b�J>�w�7Ϝ]�Y�|j���T��l6{:+��a�v��3h���O]WT�Wj+"n8B�}46�nŜۺG!���5�#�ORc�:����6U���:��z�z����z���\�y��a�E�#^�r�������Ӡ/���; ����h���eٯ�S����e�8}�+����T��UA�t^]��L(הc9�G'���t�eUR�	n�p7�(�"d��t6v.��S/��2��'*��3+3����:
lU6-~��{G?$t��uRݷO������F0{
�ԡPt�H��J=���|��W!^���\n���|�lU6��^4=<�;˽��~L{E6ݺD������{��.��9�#��U&{���!\��6M��ͧ�_�f��e/{�<3ϔ��5�څR�g�N�;��"�z^-���֛�Y�-y����-'�$�룥m+���E:�������i��^������9���B�)�2j�����p��/Y�t�0b�v1n$]��� Q� �eۭ�bь�]�H���I���lٞ�Ɠ*�f՗1��g	lQNjMu��[��D,l���L��ְa����H�u���J��J��jG	�Z����/�3ԌtcqY(�wm�6��AG/X$�^���|l����7���&�F��[�g�՗��E&�o�Ǎedv�>P8-{�o�s�ť�&>�
n��������rhU/U=3��~��&���'{��pl}�m�O��U�C�cݏDn��i���}(F�sw���
��lU6�T��n:�镻�7�9�b��LUw�6>o�~y�7�*bY$�a��n\,����R[tʑ�4�`���³��|M�rTz��a{��G+ew���=�G͊lSb���ڀ����1�等��Kj�m�ٚ��R&����:˒���콏^9���e\�ڑ���n��i��Ηb�UŰ�QL���0�h���6����L���;oz{1is�Rc��e��b������2��HUغ����u{�Ɓ���H<`+�=UHU!ꪫ�J&�`��;^�4���y���K�Qk��'cgc_A1�6bjG�SMb�4#�Q��dee6r�^$���y��lۚ�v����=T_�����b��6�|1Z�W�M=Ih��=3�_o�P���bL׍�l}�+��5M�ǋ�E�睪԰�����d�dP��.��ĦQ���^�j]ޚ�y�V��clY�I3�w�\��6>�l�b��{�X�YU&��e���O&���u��1Q=űT�����:$n�qa�p�����!^��l^�4�j��g�PE��0F[�t�6�ٙ�b�#	��	$�6I�k�٦�{OW^��\��޸��	��Sb�M��૳��g����q�v��<���V􊡏ۇܩ=<;GͶ��{6�]i(I���;���U{[?Sm��<�t��|��B��:����O���L=�(���ߑ�-�?[�}�].ڎ�Z�����/�NO�*�yw�*���y3a�wĊ�l��m�"�����>Ф�~����T��UH
�.�U�n�64BX Uع�(�ScJ�	fcf�e�xI�gS����b���Lg�����-2z�V��ql6+��n{!�O�:z���ѳ�[�^�>�u}5H�W=^;�rW��U{�-�nZ���9:�W�&����Wy����Qh{���L��z�O��x{'qs��5\�^<�K��T�oj�5��=���;�V�5�I������?�?�?���_��G��Z����aE ڨ���HC��d��!!�$@}��  "�3~B�w�X�����r~H �'nE�`���A�7ڒ\.%r��	�H@��?���'3^��q��ǿ�'a�yއ��1����B�n�k��oL�o�ac<��=�H��w�X�}|���	����o�ϳퟠB�0>RH���NI BB���,*KC��nD>4�H���?���>?�}Lǡ��(�~!!�?*�6�����-��@��>�d2ZQ��{|$����͐���U��dC>�?�Q>�~�~�'����	;��ݫ�s����!!���8�a9�Qb����[�M�`������H@��=L�)
����{���=����$�>��,�KOg�C��C��������_�G������'��R!!�f�='�~0���I�ϳ��0Z���a��P$��ϯ��ό�!�d����>a�{��'�������4{��B$!�'���"(~��̛�`7a� �љ=I$!!�ԄHC�9�'�����T�~OȯW�6bB{@��}�!!	fd�YTc��=���=����Ɋ���~������&1M%D����2q}���d��ç�����g���C����'����C�B$!�I�#�_l�O�g�g}��������K���G���-�>p>=�gׯ��!��[�����y�!!��/���E�HO��a�@��>R~E�0tX��O�s������O`Kt?f���"�6�:.1�,�+���}�>g��P�~�8�������3|����ɂ!!��=���B��yz��p0�}u)=�q�<PD<�|�^�y������ c � BB�$��ߐ>�t �?�����W��$�	|��a=�����|��`r&Ęժ}*�'����@�C��'��ܑN$&D�v�