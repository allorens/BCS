BZh91AY&SYz��֤_�`q���&� ����b@�� �	��k��46�m%��iJѶh45U��m�Km	�!R���m�T�bH�MT� �J
U
1P�Y�F�&�J�y:⦴b��Y�h"�Z�e*��$�+FSe��Ū���k,ښ�eM����E2��i�im�m�ڶ����m�am�� LS`,'�ޥQQ{5m��j)m��Ri�*ETY�EF�l4�m"�Z�Ah���5MmZi�0��Im��Ʀ��  �ڊl�Pi��U)R
��   lH����qT.,SV�ӻ �[d֮�m����\YS��wfl7�rJI�j�b�%��*�[-���X�4�7uV2��5(�5�[�3kjV�   �}��Ӕ�^�:�)v4��s�)PUg��!JT�7�o*
]7x\���j�Q����5ۻH�s�O+ݚ^�9���)J�S��]�JB��UX�@��̥T�6Qc|   �Ϥ��-�ؼyJ�/Jv�Nw�g
�ֳޮ�=�:]��^�T�W�;y^T�7�n��a{�:wV��3pw�Sު����7
��Z�{�	f��m��-��5=�  >r��*����μ�l���^�z�z�%\vj��/]���;j��㞕v����zy�7wiJ�WuJVڕV�<�ª�J��ǽ
��Ҕ���Ol�m��)!�[jU�|  u�ȯl�l����T��)������oN�ރ��J�z��<yzn���[�@��q�u�J�O{V��%Wl�ܥ����֤�u[����I��-f6Х-�UV�j�-��   ���l"�'}^��ʭ5 ��;ҥJR��=��)R�ޕ�vR��y��v�Z^���
����������ު{�=Cx�T.���*�ٓE2�LT��U*�ֵ>   �s�g��׮��;�)�J���n���ۭ<p����d�T�y9�T�m.ٽUp8T�K��{յ5$Uy�w=��7��Ls��<��[�,:���Ξ���BkV�LƖ�jƩ"�  <}V���[�랺Q����Xꆎ�`���y�A@z��v�UW�9^w@*���z;�W�����]j�s�� ���z,�eU���%)�   ��A�諻�� =S�t*�uM���<�^�����cMh=�[8z=;����z����:h��V������[[6�Z��d���Um�   !����Mրc��iY����ǭ�zr�5��� �=�Sq�]7a��5�^�������ѽ���G�z�    ��RU(h@ ��� �~A�RR�0#  CLL S�!)R� �    ����J��4  �  4D� �UOSL�dL�Bi�#	���IJ#�2Й5��FA�h�I�����|]�h���?-5<|~9S���������o��1���;�������y���  ��c�llc��m�������o�������}���0cm���U���������}������������?� c�67��~����������?�`�9���0Y���&��gc�&�}d����ɰ2m�� �� }g`�����0}go�C}d�o����}d�gm��;lY�����Y���l|�1����c�M��>gm�c�M��������`7�q��}d���q�l}dY��c�&1�}gccc�!��Ƀ`>��lc�8�l�l��`�>��`����1���Y1��M��ɰY������Y��� m��m������;c��񨏽����K�f�����u}�+zCI2X�Q�VT�ח��r��0"��懶j}��D�Ad}����4DL�dzL`�n�sq=�me=Vv�2e���T%�ȷ�j1������72CY��x�D�l��fa�R�gf��k9/kI�U�b�$��S-V ^V>�\R]��/��5�C��6��(A6�YJ]ݕF����I
KaBC¤Z�d.S0P�t���J��5�ð�i6yBX��T���z�i��6u��o^Û�� ��_�Bn�D��^�Ͷ53�����lӲ��n�e:�V�-��&ɵ���N��fv��h0to�Yvڪ)��@]L;���6�ܖ�i�<45���Գ�	5��L`�vJӁ�5�Tɍ��Wzh�� �C�C.dwl�&�+�"i�9�����̛q�ݎ4N}diE�
��rۚ-mY�WD����9��=kin��F�A�Ò�kfÁnQ�jb��"۠3�	���m�+6�%$5�$�%̹��aid{,�x�7X��`�ܭ�j9��K~%SjA�3p��m�2\�YM�ᖗ�tj����!c��Y[�,F4�B932��:�(M;*Zr=1ѷ�J@_�Wx�^d�+N�ä�[+-��oCf�Xt������ӡ�!v��Ò�uh�06kkي�5�?0H�*V����d�Řl�Vl�
��&�G��Y��N�������izT���F,k6-���R{{�'�ł��i����Hۨ�-<�7����I[to@���E�&]��Z�B��������4���Ȕ����ɾ���E�.��Л�-Ih���ɲ�w�7�X6�Ջ	6�sn$Q�J'!�K���m���w�i�.��][�4J�J�Ӛ�lF�,u5=�5{�*U5�CN�ۆ�K��f�ifRl0m�.a�w�3Ν�D'Lpv�f��h;M��#�/q6��ԋ)�u�,�TV��y*�c�RԎ��WW&6$����}.�Z#�tVm�\��LhV�i{�&1f�ְ֥�^�In����kq�/��]HY���mr�6L��g6�҄�j�nV�Kƫ� �&Kh���+�ݳ,�(��-YR�4�T���]�2:�ˉ�w(4հ���HKfCF���X�z���|i��Rk��0�o,U�'Z˗���p�Y\_*6�]fֽn�mf�|�rgh^�q���P=]N��}���֮�����o])���P��i�%����"�hDL�Y9�\wh��y�*�.����tu^���V+�	Oe�6p9u%�/m�pV�kf˥Z�G�H��"KiA���u�!)d�J0��\�2a�s%Р��{m�����ٔ�lV����I�"�.�V�e�A�ȫ&TI���
�lێ� �����a�ʕe��
��������i���6��պ�cT����kh��W�G[t7�!�@�f��L7k%��+v��4-�Y��i9Dfʖ+��vE�MPһ�y��DJ��k,�c�]�݁�"A�r�#�0�뛭���[�[��3��yV�ݼ+-�$��z�ѡdZa� �;� :r�2.X��r�	����D`v&�XVQl%j�7O
l�̓Dd1,H��4�RC�)K$C�]D ���8�
�u�̢-�����:��1Q��(f�7v��$D���&�i"��Y�Eo5���6��1�VK�&e<n�l|�u�3pC���۽�Y5y��su՜�
�c�����7�yn�"�t��{1��iW���cS�4	F�)ve�a�����ŗ aH�7K��a9�-d�v��A�YN����o��B�m\r����6f��1� E�^ �+*��齁�&T���ũF6�v���\��&]�eK�"
K�	qY�B���]@ɴ�U�fEz��l�8d��EV��DEdV"	Mi�ueVo�DPn⸷5P�Y��R�S%q��J�:y��=�����`�x��7�j�����i�B�$h����2�}4)YL'��9Y���Vlܷ�#��j�YZ�i�׎�ж&�!�-
���ևp՜-��D]�H��+4&Z�i6E�c�*Q8��a�w%멏n<ʺˬqԭ�m�I�Y!Xb`l�ukNֵ*�B)f��2f]�F]� 咖'A�D3@�l�flCi2Q�˧F��	��n�e+�`9�$eUː)x��[�׷��L�b�xU1�(�,un���rLB�kᐱn���D�����L��s	�;a��`�cޓ� �Ҝ�f����.ر{a��6�@$����Sɘ�iŘr���wRy'4ޢ(���	���b��ԍ!���$�rQ{ʘ=��mx�=n���,��� ��F��b������)���&�q�M��C���H4Sb	�`{0�xƉ��P�݀�й��W���pp�k-Y�$q��L�+i��[]�w���	�Eb��a����IY��L*��2�Ƅ����-�x�8��;y�]��P�ܺ�j(d�V:T��h�va��Ԗ)77b�S+9��R�Ҿt!�3)e�)ikI-��AWxq��Bg�d�v�0w�5��V���a0*�3�#Q�Y���+%����T�}�B^��F^�^��4E=�'$yva� ��[kL0�1F������X���,��tH��fCFEF��n��F�HQ�p]�����%�v�<i+>G�a�ǛKX�K�_J-�z1�
u�jؖVRC�Sm���wmLp*�
*�)mm<@b�l&U��e�ka��8d�0Љ�.�ݣ��jRe�(2��.�2�"MԬ��YG�����l�kY;�m3�j)ѻ��
˟`kV���϶gΜ�9W�鹔��.ldǌJ�W�VԆ^BJ��/�5��J���mh�9z%T�x�
b��m&6�B��CP3w{@�~�lgZeM�b�;jF�YZk0���r'u���)�?���W3>��yAT��	��nnS��ؗ]p'%s��a��n���6a��M��}�H&��K�lC�@c%A���iB�ٖ�KE�w���N�a3Zq�n��q ���b˨�׫�	�+@za������/�X*7Xh��n��9���ȡ�׃�_c�FVI���`���dB��`V(0ae��un�Nnf���i�m�
8V��pAB�ݣj��ķg`ΧC宒,�|I���H�n�ZO:��m����G-ŋ`��X��S�q�����Bǹ�E����ݥ*�`��T�*PVjx60B9\�i�֣��օW���%b�v�D�:��۴ھ��.�-�F�79Հp����T����V�E&�m,�"s#7n�)�V]��q\Z6��7Rq�T�
zڨ��������ܠ�P
nl�Í�N��̒����S�OJ%�6�f)�B�����ki�B�ђR�^�ŽˍA��n�W��<�-��:tJݺ%��ne� [�[ ˕� ;3�/�x��K��so5,*��k����;>
�,Ќn�3G�-��P7�^]2�j��NP�����p�d��\�O3Z	���,B3��!V��͖�R���u�7�(ǋaz�٢Һ;Z���׼�i��J��j\�e�Z!(� ��a��m0R�-���n��:�r�T%u>G6J��h�i<�.kU���;E� ����]�+P�
WQ�ڎU;2Z7y�a�bM��`�D�(�
�ʗhD��{5�F۵�8��e�Nb��ٳ�۹�IF�e���;�*L���&+�N�atY�M��M�Xǹ�.mm�^�SV�m4�s�-�H&*�<��cn�ڰ��2(A�.��C;u�4h��Q�ҨKh �hY�Ea��,@��%�؍Ն��6E�<��\t�޶�	��L�y#��@�pJ���`3`"������G*�Z�e �lh��x���1b5yX.���[VŪ��[�7�^�2T*yv�A�1adf*9�F�0\���}����j�]�J���㭧g"5��E�j�Dm�ݩW �Ȗ�&i��+"�h��(8�廡���Q�5$v��J���۵����9����[)�HL ��2E��fO�Qc6Ne� ��5�r�fT�n�hD(�VT͂����;u�(h�9+Ŕ�ĝ,�Kj�.t�����t�Ъ:�JV���NkyLe�����[�v�9&�&h<дWu��+^eSF�o^�3X��a�v���<tʏ$��Mm^d����U�N�nb8�pJ��˒��D2����R�Qs`:e�=�V�����Rņ?�t[8Cu�6S���$�Y��i��:/T,�'�ff�	يn�ܡ������#����MDb���6�a�e�4/�ڱ�3���A��j��F@m�P�	��*d��E�����A osu5k�o^i���LY��*T�9�ӫ`Ry��vB�2k���{�\��)��Q��Q�2���o3D���i��$�[Xm)�hh��jn4���Mc�VCdI�hCBX����#����A6�VT�#)��]�@�&{��`����6��5B�ƽ*���"�Z��jf����J�D SYY�R͂�sj���V'M�i&Vb�������P��sD��<�=݅��2�t���zF����JF��l3�
70ڥ�YZ2DiѼ���z"��K$��bԯYĄ�ߘ[m��R�;��:��8��1a��&iW>F��S�H�ny2��Q��D�۠�"��L+܈�`�f-fܹ�����e�E^Ax-�7R����by�h���fK^m
Ca=��^�Lb0�`�)Z�MLҦ��Ӷ0��S��aJS&]�s6�2���Tj���@��� �Lz1mn;�k����b�Z'.�NرdZ��U�"ۺE<�T2
���W��͉�r��#0�E'xB�;w�r����-V�J�������e5�]�#/p\&ܖ5"�B`��T�hǄ7�z���Ю
ER���Hr����r�`��ܬx�a��c� }��	Im\Cq��L�f#���q���bɤ�	$��,X�r%Z�̳(j�5�f��.��{`�Ҥv�z�IYWu�����D�M������/1|$I��3�f0�[:tޗ`b����'�(���V�b�Cnfeec߈�!�;�hJt�F\����a�pS����D��j���7�n�.���۩Jٲss2�=�J���������ӧ�XN�n��,����%�6V�mѣ�ؗ>F�mE��Ն1���2l���:�@���`v��ֱ�v��V�[��*�4��;RXv��aT�+A�[d
OD0�W�dk�8���S�*td�6���n�w���l���a㹐K[��Zv�n�m=��`��Hf��+OkF%�Ve���n�L� �x6��H�q��0�W����ն��|@�ݺFP����~�S$K�k�9�s,�ot4s4մ_Ҭ��޺29�L�-�GVV9��݀S��vvi7��<�L��K�S2�<�a�h�,ݞ�R�M�յ�,�(m<S	8��qK�`������� ��tL"`f�9�HXd�I������ۺͬ�Oe��:�M6͘0(hl���I�oc��ˁP����7M��)$��tn%��.��&��H���3N\�&	��j�Jrc���I��e�:���ˬ��KTĕ����[��e��Hzº̷��:3R���dH��1F	�e����� FV���W�(�)Hj���8E�����(⭽�tXՏe�K�L1� N�JD6���7[�3'bXJh�Ÿ^��sX��qk�%6��\������է�k0\ci��('�ޖM����������q�w�n^C�e��?E{0a�3
�a��եY�m@��f����1��߬�AѵK��AQ����
�,S=z7[oo@YZ.�E-r�`]��Y��Ԗ�l>0�����@�hti`��F�,-��ۍ`�X�x��si(e�xe�t�`X�qb�M:3D4���cO�¤X#@���e����Lذ�y��ˊ^I-�l�����ő{[Ar�Ə6�d�h�f���+f�l�� )M�Mz�d�46����1�:�*�ʬ���*�5i�t4KN5�͘�"�kJؖh��3J�ǅ�i�`����E�#�J�q,�i$d�)x-��:"�J�ۚ�i���EtƷX�����V̬�c*���WR2v�V�w6̢跻>��$�g7�+"�tnњ¬ʸ������Vc�DBՉDc��ah����B���l�wKd ��ͭ��hn�9ThԤ6b8�dI�'�U�]X�	��Lx(��Keĥ��Ч&��ol�ŒX�Rm��7�Sw�>k��Ji]��tɣ]F��l�8��YА��=��uu�� ��iC{�$f�d!ڝX�㒚��!V��O,�ŋ��\�j� 8 ";���jK�e���wwj,{�E
����꧚RY�w*Gc��.�����]�9���4)���G1���1JU�������
R�E��tIMm0��b�=��V767vLݎ�O(tj�݆��f#����A���eI��[�sL�Q����Kڂ�����b��[��G�ٖ�ʕ�<����t��.�%4Q��2����f⢖9@ p��yy��Q�
%�^�/� ; ؂e^ ���:~"2�Zd�VtTMr��yK\��ּT&��`�/C�Z���F�y��� �ن�Ӓ�w�q����m,��������v�Q;LF���C��D�82fj!e���gh`z�]3��8��5b��.���	bd���ɮNq]�O�o��5�Z��؋�}��M@N�93(��C��Ҧ���A���6�v-�Z7�����zڬ���;T����6�1�?��?�חm�� ��`c���o�C|�>���N�<�l�}��*k2R2U^���$mf[�hD^��wt���Q��l��	j-�j�Ǒ����WFK��!��e��3����ڰ{�d�s�;��2�ڔC�Ԕ[80G�|P�K�ʟ�Iu���J�ןoL�ё�ÎG�\*�"Xv�A���iA'Ȱ�ͅ����i����u�����P�T�i����ʕ.�>��U�>{�h�K*j�i��U+����r�F]��m9���Da`��0���( �R��Wn�]�V��ozi�FfI�����pY��ӿf�v��d��v촆�U9.�Į��.�xk�*�+f��Dַ�s���C����vf�;��0�逞[�������r\Y���a��hHo-F*�\�ӕN��5d
��̷�$μĨn���*C���YZ�6����w�+
 qH?v@4�����q��CZ^F*� �V�(�+n�����`\�ó5��f��飩]��S��13o�`|�%��)G*�x�f�`Ǚ�<�H\�B���!Ji���w�M��e��;��+���7R��<`ƀ�ۮ�r�u�@�_X�qŊ�g,���]"h��L=5}`�Rj�!���W�ȹj9�}3��:uA�;FP����k�WՉf_mM�Y�5�Np�p��u�V +}eb�o5+���#�ӥ��e��Ѡ�����@Iz�7+U��LZ�3�����l詞ɖk� ν�����2 b�s�*$�U�HT�l��Ta!��7z��W�E�)w+=ڃP��]m�u�F��\�U��s/9`"���Wvlf�ꉑw1�Q*:Y��M�Áu5.�wO���#���\��o򨷛w�)Ʋ��(t���z5Ӊ�
�m|Μ���#���j-;�o�TFi���g2�$S�G������.���DVvb��{�u�1���S�;��(�z��V�ݱb7�N7u
\��'�~�z� ��0P�PKY�]�;��X�v�PSv>�h��*��������2E�3-�LF5Ҋ��8�u<��-j�;�� YAU�o n�w�
�S��%�[)�0�����Y�NO�W��o�e��eo4�Z.ڮ�.�tWJ�GZ=:��[�'Y��A���v��ym����T��B��EW�p��w�2Z<�� f��_\&ӡԮ��⨪��'��V�t��*�=M���=�a�-�0uu�N�7���1��MҾ��BE�G��i�ޒ�*i��v#es��(+5�sȹ�u{��d��+��d�}/(��%V�n�ׁ�~_w���wtٱ됧|�o���,f��T�:� �)M���n 6)� ����Ǹ�S����
��n+��U4�>�@���:��J�ϑ��E�����ν����#���o0���ֲ��It�����ݓʘ)*΁���y������p�m��:�]�~n+��ݥ��,�V���[�έu&u�I�{\6�X(۹H��z���P�[�����b�SE�P����܎��G��U�7S+lW:�kQ�s�O-��s���|����&ݑ[�pA)"ꥍ�k �[h���y���� �����[7q����C�P��5!���P^\;�.��B�D6�H{�d%�w����*JiT��A�B��v�p�W4j`ôL��ʳ�����]$�|$[�J�ۦN;x+@�U���V��wkC��/s�G)�'�d ���Ǉ,��O���{�n�`2v��u���V��F�[Dm28�d^,�>XI������P�[��G%�9�6�i�J�V��v�נY�7�ĥ���B���l�yQ�|���5 h�`=�Y.�#�UΣ�YPC�k��4��ۍEq� }�*ޕ�N�H��3��%)�]�f��P)a�O0Ll�DN8���������-�*ټ�"�=�矵]#�n��F��h�C����4[��P��oKTd� �u�ƭ�B�=c�ɳ��i,�%*���S�gL*���؅����Y)3c������W�'��}�u-�Ō����C	z������[�b�bX]m�!el�*Nu�\��lУOP�g���^��$��J�,=�I����ق�7[�s�j�p�$���~��Êԧy�o�s}�b^�\���]7�
Q������t��ڃ��#���-&hr�Ä���;niF�@��*ɩ��
	Y�Qm>���� ��,ǁ��!��]��=v�^�(qB��w�T��)̢���^a�:�.��v�	[�+V��*i$s{S�`�8�ʘ1c�rT�*n�j�1��{Ǻ�����	�u	�dT�>�勶��P�M\�2�1Y��b����;���p�AnKP�2�+�r��c���q����Q���r�7���N�����C�ե���a�u���}�Ƥ��[+�d���:��eT"����/�z�4{���\
-T��l8�{���C8"�;�G�׳ 7��9b����5Yre�v���Ն+�M0��m�nB�"���T��~���@ �Wm��؅,�/�9W��d����g���#X1^ufd�C�)�+:��g3��P4ձ�nH;�dďWk��-�����G!i�/��Tέ
�s�V�[�[�)�N��jS������gl��4T�=P\WW@K��*�`KF��_s������r�d�C8X��tv�	`_R�|��!xBɭ@����J`ظa���H`MJ��q�q��ؠj�5���E�9����e.��
����Eb�:�rK�ֲ�g�m�ʬ�6��4��r��}��N��{l.�J"�|��t|�	s-����Ȫ5Z���R�B27}͗�����L�ܚm�;���(�X�I@��b�{���gm�1TҢ�,�>�+W����V)Q�)~�f�f _b�W�|�����I�r�Y��v�1�(&����{��H�\��M���K�9z�yqZ׮����8�cBЬ��nVd�p����x��B�&H��7��.�+w��1�6T��I����"hP;�n��*�UJ�\�y�{�@�V���&����
Y��H�g.��:Yջ2� ��vNЂˉ�u�u�+��v�!��8�3)�+V��1��� bKbn�f�\y-��k^)�.b#|.�n�6%���S&e\졑� �8'�Y���1�p
`OtRwI\wE#�Y�o㌴����v�XlM�)�p;܅v�bd�yZ�T�¦���8�t]�#��!�x�8�V�ŵ߹��vZ�f��\��-��{1z&m-�Y��������I��H+k0�:��o��
 �x�kn�p��'eE�����	Y	�[�Ĕ�no'y�*E�9c�а�t,���r٧���+wZr:�����uv�{	i9��	Y%ܔ�t�>]�c�Sʈ!��=�_��vސ�=��,ә6��.D�:�@�v��^p}H�����V2��X-;D�1l�K����cqmn�=32C��[Z8܏�ҟJ��F���\���{r�3��V8���H@��T/㑙ѽym����V��%�-Ώ�\�`iBЊ���1|�/C'a�7{^�q���{ �5���Z&wc�/�=�J�]����w�.��F�A��v�+t`�����|�k�N�p�7+�L�@�%*5����L�/,vy���w,yG-:�Q��q���w���;��(��a;��݋>v/��h[����I��e�*����tx�#� �*ֈ���h��Qf����yl�d��Κ{��zmR��ֽd�FZ[�����6�aX:���\�x�\;�j!SݺZBNF�u-��6��8��$Q�1�M$nba�qc���:� �n���)(4NW�m�8��m)\����pMuvû�B�_1��)\�d�}ɼ��"�N�EV�Gakʳ�^+��"���)��&,��Cop���=�}y�[*Fv�-�wิ����{(ϊ����1��W���ˑ�6M���D镁B��;7mi�:�q��T���VL�C�oNܧ��M�N��.0nd�z1�"��R�zTt�ZI�F�J�.���e�I\Z&�h2)+�O���y��癤7��Į�p��1��7(�N�Һ�x��T8��'�����̭�b�����q��V.���:=����\�ƺ��Ơ����
�J��*IngS �cf��"�\�yt�O �W
�j}�Mv�ە��\�î�*��HH�@,m��!�ǩa����znIv6ʁL���Ύ��1�@!�wf�U�R;�ݱ�vH��̐&m�Cp�E۪�(�S* ��ɴ���0#�����^bC, �����{z���X�9�WP�o�p'�ʹ�F��źinn��5���\^�n�{��e�ݻ�;)��!��Λ�-@b�Wvʜ�.9(O�����9�ΑJ����#@I�sa�ۭ��عQZ������!�ً:��Mt�(�t7��
����ŭW�j����HJ!(�۰���[v3�D��d70��3ے�k{����I�80�5�+�a���f&�ٜ�o)vܝ��I�
S�`\[�[Y�n��u�is6���4�	T� �E�t�P4�읶jI����2�fn����u%⣐n�e�bz���t�k�3����`�_o�m�b�eK��W:�7{0�o�έJ�۽�fL+&��������Qu����5֣B��f�-�H>�}Ql׃qf7��w2ø\�U}Q
͑L�[7�7]�) �15k{I�� ���b��\��s�5?a��XFY�ކ�p��/�W�Ž:�lZ�1\��s_fR}�,H����m�˶�a,��5��;�˾�\V�E˨-�Y\g^��iܸ����]�|��F�A�ox����ek"<�nJ�)o5�N�1�/y]�7�կ�`S�ùtnk�l-�܃��}g�����-Sld���mN�2[��<B=r��Q-��#�76^�]{ `�9CCS/,kwF��e�,�x��ُk����s�@�߲��+�٩�����g�(��n*��`xI��z����R��(C���oR��z�kZ����]��
�V�la�ľ�AY:�Cy9��%s��)���Զ�[���w l�X�l/&�����gl���J��9B�e5�+s�e>]a),�7�VG���"W	{@N�)1��ٲ��4�ʋa1��?+��s�{|��x�n�֩\��W �%ܓ�93�+K��Ț�t�0�Тk����/:���.�f��w^L28/"����;su��Ϋ�IY[V��+2���
v�wu��oS{�E:�v������bpޠ����{�'9SF>�����F��@� $Wv�:�;nf�!�jT���;��� ��E�WX��Ʃ������]9խ^롫O������m�;�b>����K�֤�ݎz���S��[T��c�1Һ��	�E#���U䊱wKP![e:���ToWr�]�}2s5��8U��pj�������l^�n^Y���(L���L��MШs�&�&�Pکψ�0.Ч9׺��}Z�B�7�T�|2f���u`�~�}���
�	Q���������f��ew}������
�hЙ�����t0�8!-vA7(.ky�5��֭5}��kSL���qg\���K�����s1�.�*/�R��@��K�33nɩ]��V�s�y�ť��s5�r�-��㕐qn�`%�Y�K�S_g4��|����܄s����ݺg��3u�!�8��y4;tچ<�l�M-o�J��e���3��Wޤث��[��6�����>ڙ�n�bȝ EoE��|��w�]���P4q��f$�2���#�J@�k�������j�v��3�ݯ��=�J�;�H���F�9�ne��EC��iG��
e�,"ĭ9ӆ625�B�:��9X����/���L)"`�W$�:�nnVg�-��'��T��up�bҦ�`��k����]�%�<V�]�Bڕ�q&��!\����l��mɆ�R��	+uj�Sa:���U���3��A���}�m܁JY�Y���d�����}�`�ԫ'AD�>]/��'���x�]�A��Ur�)B�uj����X�ٔgo�y��*(Vi1F��1\Q�/3{����J���YJ�Tδ�8_ĚфG�ӕdus�B��Ӵ�s]0��̠1eԫ����
 u.%"�ޘd�c�i[k��/v�Q=��w�I��yRS�& qĨG�	}l�S��N�{uW7]C�.vj�$����A*��٣k%]Κ��/UŰ�/&7����7���;3kx8@7n����������3�ѽh9vF�O�����]�UÎ��@V1ɡ�a�Q�zqT�Y«u	D�!�xib��#��hMw,>�����
�Ӯ3�5��]ų)�j�A��+���{���̃ge4$±�7mvw�:z�빜���1�G�H�{�VK�8!n]ń�N�N�W��6��+dm>��&�@ �F���:/��<�+����6!�r����2�Ҿ�ՀvI�5�$�r��v��"��{Q��S�d���#���쉔�ih�t�^8��x�D�b¡E�(
]l���·`�/�vKC-��nB��^<�t�#�^tx����ǛV�p��u�a��(��}"�ó��/��9���%����Z��J��;�����C9�
G����n��Sk�<.��h��9�/����L`��ꤓ��1��]��v�t�a�)�6��L:4l� g8s;�[�hn@�Zۭ۟9[B��}И�FV,�e�q6�ٹԷ}!Υ2������eclwwr廉/ɼ�b��⒬��6�|��;�͍�qc	�4w�@FJ���A���@�10�P�@P�Q1DŁ"�c�%�a�@���N�u����L���~�����6�o���l>���?����< ��������?ܿ�B������N�%���TY�cI�]oF�ԅs.X�����;���WQԻ�$��o#�!&:�+~�P��S��Ra ��v�����e������8�s<��P��"�SP��hq�혟Q��9H)�-�1��YgYv�sa���#�N^RŢ>S��8�k�@Įs@�S[�=�lXK��TN�g�|�{���{p4���r�v�m���j%85ָ����:�B];sJ��
V~���Y=��-��a'L�ٙ6���`htsV�fw_U��$A���Q��p	��#�9�`@6S��e�T�1�{W��	�a8y|�U
dr]���Ɉ���ǫ��˧!��7��ӈhtI�bgT�dfN��4�*����d᧢ʀQ���lMmh�cZ��CQiT�R�7�{��v녺s�T:55���k~�:�%1y*�I��d�+T�/0����c��7r�WY%t��wI���%����[򮲓�nI�I�h��bl��n��9�KW��B�9��Y�N_:<���X=�Tq:�Cȯ��"�pl2WPni����"�{��n��}\^����h��[Z^h�<� hR��=�=R�7i5TpZ���*A��ݶ�h�V��u����gV�e��\���v��*\˙b)E;x&���2�c[�e�{�+<bR�LեT��s+;(N��NQ�
���(v��7eYVR��gE"��mUގ��������+�4�A4�����>yW�Ǔѽ��-��R��ۍ�i�s��v�]�;,e�T�rA
��U�4�;��*����̝�m\�n��+OT�Gwx��J��w�n��բ�V��%l�֫�s�*��B�q�s��� � u)�V;��`s��G%��\v��l��Z)����Ƽ��
`�k!���fn�j[�:Nꢌ:o)P�����o(x����͝��Ŕll)�:�Q��vc�"])����bb[DY���6�V�U���g]�
�.�eۂ�Q��u��U �]���U�Z�Mν�R��4
�
�sslZ�7;O<��V���b�i�����+*U���c�p�1�u�ܣk%���8��ē�e��'a��i	{� �pb`�]8P�S�������Vk�b�)���t���;O3+��FG�z�=��u�p@��Lj��T��6��`�?_A�r#�t�J=��6����n�MWV��m���2_f�g�֮�[�a�f��F��n*�5����y�\:6;K�{�p	��-��*�ı͑]9h��ssPo�GB���^Jaf۵���4�d���6�y����1d����_M�D��6[$k��#(<��pJǵ�FB�|�<	��i3^���q������l�=�DU���w�2��Ì��T����b]�up	�emi��V�g�*F�뻔��i9O�rc��)�x-D�5۔�c�ɺ����c>�ھ�;�M4%��%�킆�;qAЂ��;���yϴ��]�Y7(뾊h�.��d�Ō��y�ݫ�t�zj^@�Vph�#J����b-�l��έ��|6��#s��n�mP��v�2�����#�c�Std�[L���C3�'1A�KK\bjʎ����u|7���e�m�m_`g��Ά�ml|A�)�W]�|�����Dd��5���w�z9�Haْ�i�5a����*��s���7ye��a��j����&���kb;5�tg7�ym],���a��{c��ei��t!�͌���G�����eE�ݨ��6b���/@�h�X%Y�T�ZL՘�B��fRx�j/Q����:6�b���mɘ�o ��c�%u�ӶT�8e=����fe��s3Q��C-.w��fb��`]�$�[�����#Ҥ߄&]���j5�b�׶���;�.T��֥ȍ0!7�K�؞u��s����k����\��cpNܲ�#���k�V�'��R$jL��̊k����U&hP�dz��R�g�����3�.[�EL}h�Ck12ە�\��?�]�.FZ��YRQ$]�LS�K@t̛wR+��h��4P̨�R�1��*�ե�-?"Kʇ$��;
EJ&T5h� �;;�no>%�aк�Ҭ���䄴Q�K���X�����"����Ev���͓9�ޛiPl'rr�YN�����95�� 9^-#�Fw����P*Q;�m=9�eݽ�s{���`c�(G]k��i�� 6ްJ W������礠kJ��6��k���/�lWe�HVtO��1`(pJcw��cu��`+��ȯ�P������*j��&3]�s�4�P����1�t�=4rS��5����� L��`�U�{��a����3��6�`)���triwk����` \����F�d<�Lw��U�;)�s�1�\=]N�b|GW.zczE�Q�:�)�9v�@��{c����Qh��d�Ov�:�[����h檥�Gi�T`��2Q�i���ݨ�]N�
��|��
W��oop�SL�\4��&_01��[��\��� ��k%	�����6%"�Ņ˷�i-�u��ҫ^��-D��/&n�ˬ�i���D֗jp]Z4Z�#���nѓ�+�1��o�D�h}yĭ� �s���̾��Mj|��bjX�:m$���t�V_:Yt�x��H�,��p�s#X2�d����̐Lt���T�K�VJ�(������n�BP�V,�}J���e��̐��V:з:�k��5�H~%X��٢���$���ՌN����ll���V�{՝w�,ѢFrYͳψW�+7����oj�F���i2��pjҚ[��k�-�q������5a��!�Qq�|�G�D��L]]�Sҳz�F�����n�)=T�β�[�f<�lj�9Eò�-��n��o���-���{EaC���bK��&<Ձ�r�6;���ji�zi�	��&9	�`���oD�Z��n�������n����.��O�}I�9N���.���kۇw��P�Q��B�.�`�y��޻�Q���
Z,�����V(2`�頳E"+��D��X�U���MbPvXi���k4��ʅaYɋrj����#e���w+S�S�T�7{��vfkYy�0�J�klV��'y͓B��7(\�+�c�w�1�JN2�w�$�lh,N�+n���0�;��;�I|���4�u�U�>��lh�(�����G^ܹ1�\��V�~�@EN$좪�#S�X��F�t��e7
�}�^�ݥ��a��HUb��W�����G(Ir���Mec��i�R�#s�ˏ�)��'i�m�t�
�.=�Ԓ����"�tP�ڭ�{�� �IEb�Υ���oU��WjK	7��X�pY���R�"���¯�:��J�o��GUgs��Z�Ŋ��c�C���$p�Fp�+6p��Ftp��c|N	W��ߘ������ �Z��_&!�� ����Z��:��>�k5��31�@c�V��W,Q����N�[�W#��g��[�1��GpL���X"R���ɇ/�X��P����|MLTw�����B0�GZ�*��>�o
bH��gu.��s��p�������y�λ��U�%���b���,��2���ph���"���x�Z�{ +!��a��������!��SF�c¾K@��:�����弑Q��<���῎c���Y݀�u҇/���T��hR�o5�3l���k[��]��"�AB^ݞ�55N��r�F����,�nX!4;�T�HqY�1���fV���^��V1�Ja���IA#畳sŘڟ=���x���u�"@�O����
����OKd�����9�5a�f�O��6�`a��X�*,�_r�p1]eJ\˥F4��6M���u�-3jb\�L��ꓥ��ma�&b��<��B��o)\�ky�oM�J�n�A���lI��p\���i�w�u�Vw�����u�a��ܷ!kJ��!A\	u���7]H�3l�2��A��r˿�oK�"����1��J��E2�|�h�CA[ݭ��0�豫4P��xE�3�U��a�˗բh�H0�,%Ϻ�F<�ױ8���z�L�-�2Y{Z�V�Jb�dQn���hP���]��=�A��/ �o����V��ޣ��=�aT&���-�V��Wx�i�h�d�l�H/��e��ք(k�JhS�k��:�3�e=7y�U�"����E�Nb2�q��1�f�G�O����qQN�j���+0vM��U��	��*Y2t�R�o��L*6ؼJά3E���.b���v�%�eC�L�Ƅ�=�8�I���fh�I�1�Cl_	�w���OH>\��wf2��|uVc�0F��qyW���1�r��V �Cn��Y+]�*a�Rs�@71�$3b�Ymn�3�7�k��+2�C��z�	
p�S�w\��{S2V*�6�V�D_92b�M�ك��kL0��}(X�C&�m��(W:�"9~�eV�T�y�Ɯ��Vq]n����`��>�v�G!O琊VRJ3K�̵C�p���V��fJ!n�ج{�V	2�!5	[ ��ӵ<{���Ae
�)[�n�,��wG��=5M���*o����_�E1���N�SHF�m�к��]��V]��<Q�q,<��v�+�u��7����Qb�cØ����c�HW��8�	R5��j�1|A�&oMWw86�2u�9�!,E��X���{$MS�ⷓ���gr*WvC0,U�qx&>`�Ʋ��~�s��B���-һ��w<�x Ȳv��1��%�,��A�`�no
�O^�r�mڡ��XU+q�mCw�Z�.���;[�+1��Ld�E�����v��C��!�j��]�q���ݼ{�X<{vm����6�8��G;殯��9�/5���޶i�*����.V]jt-�!�*��d6��j�ry��m@{��G]'Xk�Jms�))�9t[bP���x:��� 2� ���X��lu�j�[RGͺB��ۧ}�����j�;L*���v3B�Ό!PRds�3Q �hڭ��VZޮ6�8ͭ�"�[
=�Ist���7�}х�+���l���UN�i\3�Ka�αe��w&+	��P}��Y�-,��[T���^ƛM���8���v� �S��1b�z]�! �FԹN��+�����#���)�%��q
�uy��Bƾ�;��$�y�nЮ]Eܯ�k�ơ2�V4Z�;N�ˋ/�X�xă�5h v���r�pvH�f!�.�zsj�Y�V��v1Q�}ԹɆ�]v��Y@
r��M���m��eWaq�N�ڻFj�ժ�-ݱFui@��ؙ�T��q�f�r�_=���
�*�w�=εb��ֹh��/�;n��=ඣ�C�C�]l���+��i�!�8�Q}'n��)XU�E4�=Q��^����x�S6�>�:6��s���d�j8d��:�PS��匓OI&�r�C�BY'���ˬowI��+:m�	(󆮻>�A���Sбҷ]���J�-���6��"�7}��������Ok.;hD�ܛ�Q��WhH4^�g%�FG] �Nh*/9�o�j�DٷB�	�n]^�\#mh��l�:V�K@X��H����ճ�,����|�Z	� �)��H���\bH�`�jb�f�m`钣Ѥ�S���h���.���r�oL�����C�*b������ϗEh�Wl���-�l����k��Cz��s��5C �J[��������q :	1�s�����T��Wp(���n�%Vy�z������ݙ̎��9��Q��ɼ4:m���4gqiҍ���N�c�O���WR�(h{�GZ��P��6�V��2���Or���}��;���ĩ�s�\��r��$W�"*̢�*޴��ԶXv5����*^�	^],x�"�&��V�̽i4Y�%�:�jP62�u:�v*��RS��E ���H*��ͥ|���9���[8)�m��);Uַ6qջ��Lr�����6\����Z$�����P[�	e�V�h���4��I���w���SnA���β���:���b+��������t���5��
�VQ띈0Ź�o��Z;�������Q̫8wr���-�SL\]l��T�UJ�u����.<�(��H؛b�����!.���G���k/)����%mp)a`X����-�ky�"ҕ��:��(�6��t�(�Q�5[���M�ܖk6���r$j��_S r©a��;j�i�*��:=���M;��R�pL�F��1������:����ۻe�)�YZ�*��E��wՇ3�foi��l�y�̤��]c�a�1�{Q�l��n۶{��CCl�h�ZG�lܫ�EZ!�Ԥκ�Q�4�ݩ�N��mV�����$b��X�lJ��k<B�j�ܩxA�[�Y�&�;�Rf3���0�Op�O]ּڏ" �%V9G{��j����� �tE1�4N(����*�g�*���p�
䚶5����o6;]�����%��V��a�u���:�8#o.�e!3	��F -��l99	�cĞz7pv��<,T�aH֘�ͩ4�)v���j�C�+���!�����s��fL�q#f�>s
�u���ɛ�}>�&��'@�&LHg4z�;n���$��C(������F-���H_s�<��=���Y����U��3�7�$���9�U��iYpĤV%u�9�c�=�]Ae��Y�:��#�ᑘp+J�h�	�5`�.�[�����/-Aq�a7!i��#�w�%�r���6j��M�z)˞�N�F�B`�zK�&l���]
���U�4��N|ճVkX:�von�,nOYgP���&�	pA�L�DBsc�.�wM^���3��q%��.�"y��&�N\�x̰3K�qK�=���1;�<	7���W��Y���{��{���������߫��Y��^�=�}���{����7��@��{�|_�3�9����KC���̍�������`���m캝��N赡��u}�lA��V;Gqgw���ۓ�f.�6��� ���\r��8����j����0R�k�&���RZ8���,�+gג '\���Y��%�ԟV�\��S�nn��,N�A��K(]�J=��q���@�Lт��F7������N<�e�a���E❽%�*�:��R-��s�8 S��5m�I���➻�%;��-I��401���_X˅�-�f8 儥ވ����c�¾5U����<��K�!j��F7��@v�.[ڐ���(R��c̕���%���S���:i��5���h
�S��\c�*�:��Zi��:?��aC3(SC5�2^�M-�g
u��[YA�X����;�\b��<OiȆVY˲��62U�O��C���ŭ�t�i
�¯��7z�*���Lu�m+�|^�u43f�V'����jc�F�O��y��^�4fF�*:�Y��9G��-n��/�j�6����nJh�aZ�-�=Gyt8����ZK��,�;V�X�P{�K����Gk�3�2t��:���cum8$���n��+��le��k3����o+T�q6�����W w0k\���A�,���	�,n	����"WO���\�d Mi��� �ϩ�A?��ª)΄��UUʓ�x���2p�t�9�QW�:`Q�E(9���]F��א��)�/R��n�n��9D
��#��,�y�W�b�;�&I�[��qs�\��Q<3�#��(�
��g�R�ky<����|��\6���y8�{ۅ��9[H��dU�S�	QGW����D�G">I.�yB�|�z�ET^�H�""��Z꧓��(*���qɔ���h������S��T�**����:o\=__��!}���{(�T*r,����S���_'���ϕ���\H�]�zU�X{���YS���������F��*;�I�(��H&T	עp�ZK���O�S�w5Ԉ�9�s�A�CR��W(����~P*��HE_�dE̤���OQ:\�"�T\�"v$k ��*�cw��eATF�r�Qf�\��
)-�s�̈��9��Q�l�:{���EC�v��r�=G��{�ʫ����;L�ψ�Q�8�\���"���z���w�����=�5-���*��j�TN�s�gD��*�zv�喌��Ws�w�	>�[��.�e7h#�%U�2���ͬÿޞӝ �%v}�ϔ�/�4]S��>�}t9R�KI�	�;N�����b\�QsL�/�;�M�xvO{_�k��KJz y\X������J�!��*^ܞ��vLn���9��g��T��Ĳ�v����������1�|ؓ>Տ����t�,�\�����2����\��j��9�m�����gk�w�Y����侼�9�_{UWJ/����xEf_J��Op�Nr�ɉs���]�+�x�;4rf}\Ѱ�ýx�A�� ���Hۚ=S=L�!������'�h;�w	7�v��:���0�=���Os�S޵��jg��'	�%������ӷ����������F�R�9�O=��D{�=d�=��I/J�as�c>�r���E6�E�އ;�=ͺ�pqVTn�3��uIg�����ｻ3�mS���^�c�.5�h�X=OF�[Q\#r�r���vl�R�IрV_�&p��z��ItZ�Zh,�v�O0UՍ�RJ�m�̤M�/��L��q��om���B�mą͏6a�2t��y�����渺�|���m�oM:��qw�rG|�P�[�Nْ+���B�z_"�8/��'N�\��W�87�4�U��%����<ߖw-��_p5�+�^�Gx1����3��Y�G��Etʺ�L��^���S!�z��&���D�^���:�'�I�3���{ 8�y���vk/�vA���WDg7��׉��.L�y�@&�O����6@g�3���b^���,�x��z<_r*z:���0����Q������h^�<�\�jû�<6rQ��46z��v7�W�qw�G���x�IJ�{rOe��zF�'��0̱�M ���\���^�w�)�U�}����=��p�ߞ�y�%3��Ov-q-Ҽ�ţ׺ ��]W��{������S��7O�Z�ꋾ�A���Ȭ&��O%y�{s���s�$�x��~]��&w�;�q �@Z{�3��d��v�M�Y�/^0E:,U�Y�T[�"�vVMz�x<��C�[IL��s4�]j�[59�iS���M1���4�X�떗���
�x��Z��Z�Cv��2�9}-v�ziy�P0��O�k��'-��P&�ctf�G��b},�b�����X��r�m�X�oj�ٻ�5��>�f�q��ۤ����-3Ww��˯Mg�G;�ן5��0rN��������;��)��e7���-d].~�秧���k�'=�by�1���ٙ;�{�>�8SwG�fZ}��%�l�>���$����ec[/�H��s'y�V; ��4%����}v��1�|��j�F��#<��K�I��+�۳��xL�|���cϢ.����1r�A`��a���r��s�\�~�}��w�9췟{�C��W*�
��9Gؠ	�~�Φv^-�Rz��^j�����7Ӯ�y�h<�aO� o��6{*���s��eWxp?�Ϯ��g�Rٱ�870ۭ��_z��e�>�3���n�<t^{�r�j�x�\W�~ڬ�%f�S�� ����2ڔ����B�����gz�l�=�Z^:^V�����ܭ^Si�a�{gt����hz�{L�X�W�̵HVߎ֋!{/�Gy1�+ ���@�7�d��ѭSˎ�	4�^��6�A���Z��a���5�>e�����tj��bE�ˉ���l�K���_A"�1���c�fѺ3a��RV�e�U�hR��଺c�`�����.��.ui�ʿ����~�BUkΌ4;͙7˪���=�c^)�K���D������>]�ދV�%S����$�w�Hg&+��;��8-f��r�u��.��{��O/k��&��ī�,�{� �f,l����Ꚉ���*�v{_�Ct��ɵ彛��]��#���w��]�H3��B�C�>.�W�}ҟJ�oޚ$l����%���I�kڬ�z�I�[íٟ�Fy�U�m+�S���z����y�������E��=L�/{�����ʹ��j��yC�JU+�]�q���{�;'���;Ǹ�~��в �<�	�s���y��Q�O3�d�����W��t�;�^&�p�m�8��˸���>�r��M����}쫿ocz{�[�}`j�rA�n��D���]�Kk�MN۩�1��vb���[�f��F�Ё�n��Pv��.U�T�]BN���$N���烳���v����Km8�±�z[�Ź�3s�e�.C�r����
�����z�$�0�@�p��󙆱�n�U�҆+�M8��Q��g�ϩ�z�w!�1	� CJ��k���q�k)1�=-}���ٞ��~o�+��-��G[�Aɝڕ��Z�l{&\�W��y��H�	ծ�u��5Mx\����}I.o(�ďzW���ǜ��y���`ćCw��^t��Oz+�v�����u?p���bl�H��s�b	��>�ax�:Y����M^�	�2߻=���]������{={Č<�=^f��vv 9UEw��>���(/2ל�i����kO]gyc���O���{�����,g�v�y3�4{)�5�_����ܐӐٴ�4x��^��wv�fNгho>��+ڻ���$o;�z oR2�x����뭩W�q|]̩/�A�W:��������!�ovh�Md����eo�����O��12�<�X���x�Ff�[S�T�0v�;��k'��fף��z�0��,��v�n,o�v�H����p�u�I�zd@׏�p(�(��qG���o~�����ѓ�/b#�ٮ�e�ŅkZ"�Q�O{���t;�Ǳ�R̴�*,��U���
�u�^t�1�i������H���ƍ���j�7�QN�eu;1��Μ�Ds�l'Z��̫U{Zs�@-?IR� ^N�;�I��-�<�;!����+ƺ�q�g;O��z�m{ΰó���NI��=;��R�������s��L&pZ8k����J,mz�łǯ�<��+<ު�a1>��g���/��,���ٽS	<�-�����_�6÷��Q�Ծ���g��]�^�*o ��sS�[��Oclh�9e��*����o����gzg;��52����w3v�y��϶1��iͣ1���F����;+�+x./�--�}(7R
����c����i��&$�u�v����^���� +4�/n�9A�^{�\�g�S�'[�9><� �-!�X�Gn�v��m4���������\	���S���Z��C�>�t�A��Z��"^3 �W;��|B�L�o�ۣ�g׍��5g��>�p]�Vx�d>؎\��T(�f�,��J��0�	�]�{-�齛��27Yڇ5��K�0�� <�׵g�쩄�HR�nE׼俹X�ݗXog6�>��k��uL�� 1�����MA����fiNq��V)�:fjyi^\2v=ܚe7�����՚��#�c�WzY����~UBCW�j�^�_xUB��O���<3��]�.-��kS�Χ�޾�ԝ�g��^D�םn��W4vw����څ{��x�n�[_��d�����rM]P��cn�
�be_�j�47�׾�X�b�Y���kǤ7A9~�G�����f���'k%���RѪ3/���b�O����G������7I�Ǎ�s,q�6ksg�W��C���}��f���eY�*�;�>������� ��uh>���5��@O,��n����e:�����ߜ�����r܋}�J�gPw3���U�����q�j�7C6G�0c���|=���Ǟ��ؙ7��w��t]��$�o��o���{+'tz��OD�k��q�:���`��H霂.N=�}��rI鎧��}�{үʳ��PZh�~�4~3�k���:b4�k�x�,�w@��y���iJ:�A���'�m���c�a��CX���M>�^�������0�w�R�jV�!/�t$gV8�@|����T�恆��iC�.�5'�IT@�_^��K�O�o��e���hd��cg�j�!�Q&�\�]�9yz�'aJ�W�ﮟ<�L���5��e1��/�bL���uT�|���zWOgY~��9���D =�5'�WI�n��Oj��2���x1���EX���d���ɷ=A�欟*X�^�v����J�|ۀ�J�~����x߈����3i�7���� <dx5u=��73Xp����|0���Y����y�IK=/����'i��v��2�f�s`�k�	�p�3�������W	���Ov-���ϻ�K���;�{�E��R�y�Q�x���*�L�4�ϰk�gb��}�u�N׬�ӕ7�q�����[�.�89g}/���CM_x�pud�K|�}Ü��ۤ�r3I�$�i~����u��pν~��9\�]��쫕攥]�>����{�4C*e��PO�oX�&9﫧.Rp�ip	~��=[�l�gޕ��V�OE���F�mЗ�R�7M��v���n
'\^j��]M0-o��.f��i"���@1��T��/Q��cs�k�v)��bq!��D���^��tkI}ʰ�J�+_�M��I��3�2�pM3��$��/���e[���@��3�;�"�y>���w���h����p�#��*Ϟ_� �6����V�ZRPl�r^���Y[7�jzG�z�.����C��V��Z׽���#�j�/$���i�Ow����8��E۠M���ޟw����kth��
.yw�8u���C~�=���j��Qrt��}��oz>����7���6jq�����0`%�62�r������譅S\nےr�iLsw��k�~���>()`�7k��y.�wM/<�������uXco9׶C��6\�H� q�<i��t-�\�O�;۽^-��*�������K�T���r	$u#53K�|���6�t�X��1
�����ױ���^.�J?HM��>��~��R�u�ݎ�N�^�wMsԜ���q�G�2�g���;���ػ�L���v��w�j�o�gb�6iMΒf
AM��hV�\�o,�j�X����.��q{˷�����l���@�_��<=NA�Gobj�9gvf4y���m�]���}�"��峢J,W+�9.�*�H�9[j�V�P�ؒ$2u틷6^����	AR����Q�N��iV�NV��Y�ģ�<cv�f�2�>���6���d���c�]v�p���F���}�#fe�/w*�6�*=�J7�� �mq�����3�M����v4Iح�Z8�Eݚ�̇�krv�3�Rbo����p�3�]�1OG��8���o��՟{�ff��T��x/M�~hо�)��$~>��Myx��F>��B���E�y��=�����O�s˲���,^�7�}[�~�G��C�<5��:����[��{�2(Q����T���\��Ϝ�Y�>�-.��
���z{�v1��N;<�ܜ�Y��:)����n�0|���V��Ow�o�̔��i����CΛ$˫�h?J���?QT���3��;<�'��=;{ڶ��?X~��>�6	�i�v��E{z���}� 3�9���G����~�z�ހ!��eK���>��p ^��g��M̫|�<�v�׷S-��B���qu��A[��,�����Z��z�'���哛@~�%`6zt��&��w����e�m�I�	{�O8mm.ӥ�P�;Y�������p}
̮aض��k�,�܋���e
JC�tr��o$�̪��w� @���ӹ��X�v�&�����+�](rJ�����]JĮ+*=��}��]|s%�\q�R|�(��x�`���&��)SU&#{;�ـ��zZ�Slފ(r�'t�Z�Jʌ7��	0H{��ʜ����y�ɔ�X�Q�;�=���w�wn��x]{9I�4vW;%�M��5ү-�[��Y�:� ʂ_s�Y�I�Z�Fmc�8T�j`���κ[V�e�86={k�d4݆���cN]�t���1��Eq4]�����V��%�Ь����2��1��]�L9[A8��1ǒ.(�8�WW8<y�xȸ�;[�Ň�3Wc��R�6igG��i�O0�ٔ��n2i�]�en�wn��u��f��-|�r5MT��:�q�Ӣfa]�
�Z���N�UF��ḓ�mCy%�[ې�5�ϳ+���|�o$W�6�����IM�%��c�R���i�ۂș�� {r�dC]��Ţ<(��T"Zv=�z���ءN���Ie])a��"��/��wܫh=�V,� ��Z��/&�.�=)."�v4�\u�M��gl�:��ڛd�ݹ�w˕E6ӡ:S,���YG�Q��S��p�4(���2����܉�#�w�N�\څ�$�]E+w@�<0���[a�b�6��wl�(��heLwς"|�[ �:�� /���R�&��Ԓ�#4���9S*�ͱc蒴�9ҿ�L�|�����E[ę��Fo��®Ѽ�,vK�H��f�ӹ&�ȳ^
 �W�i.�of�B>{Z�|�TW]D��3��4Y�D���z���La�um��3�%��, Hb3nj�e"�bN��q�F3#���!�rn�;�G��@�v�[˔���nb�%Ӯ?`A�H΅tJ�fV���{I�Ύ�ӥl�UsX����i��`��Gm»&��Z饟k[�(W.��Ӥ�����%
7��ۻ�����LKT���'�[��s��ܠ�q�����s�a�ܦ�H��H���%h˾V��j˩��dS��Pۦ%��,l�b�c������	ޮ���@���� s:��Fڍ�4�u������l#�D�����7��jr��TW���B�IfR��:�W���ÿ)qr����7��O�j8ԟ]�r�U�$���\���i��j)� �s���2i�1N3OWF��X�[��pLx��ilB�.���U��Yǣ|~P� ��Jg$V�N�
��@��9[��lL���Ǔ��.(�=�}�@Yc���VR�^=�\&��9��'���sd�r�������P�}L�G갹�$�U���S�<��w�ܷ���y!Er���!z�I�,� hD��s
��D��=ݑ�1+3ַ'��f|���u	���d�蕮x��=ot*�e�z�U�(�q<B�9&=s�"Q9\�����(�΅p3#���Q��Sdȯ��>o�;��Q��\DȪ�Q��q�Wp��������L�n磔|��9Ou�����UUORg;ΐ\ �8�{���/��^@W�;�2(wJ�UX�������7�DG#��:$A�2���vBI�E�:EM�*�I˓�l��9�N<�Pj�I�QQ](�E�L.G"�HVJ%��=Ъ
/��n�UY���޴[�I�D�Qr�.�9�>P�����w(�(����HU9�ȺR��eE�|��C��VE�t#F�w;��"%B"&e�aF��,�*8DD:�/R*�$�I�.~�����ߋ�ꏼ�v2��	;e�#��G8�6�ٵt�mѡ*�r��a�y�����2�����PC�ǌ��P��T�F�/�Djw�Q����&o�G���4�
o�������ܙ��3U�L�����'� _nd��2K���O6בi%)���S�F��xE
8H��k�C�$� �Me͗wk�{u��󶓙�.'w:HynP�d��!�N�k�Z6����\3���^6`&)tcZ{A��|0��-�=�=q}�0�èbS^�P��d��&�0��w&g������D��Z"����O�U~2��-ʑu4�e��SȬ��yL=�ˎ~�j�9��D�01ͱH�a-k�Y6j�����
����Q`���P�T?Q"�e���~uba?f��ͱ���V-��K�s��.�NV����Sx�c�3c�x�)�`��쐟��C2bD��݋�S96-�6}n�>�F��:�qaJ��TZrWH��l5��nr9k�Ւ�����A���/���!����Ɓ�@��Ԫ\�����|��O`�o5�X��wC�它�=3;��(U,��;V�#�8+K�a�A\�r�nr�h��Qt����a{e%���tJ���wR�&�jf��sqX�GT��3��8�Y��jN,�Nʒ�[�IV����b��ϥ.��.�A��C���Zxmc�6V���op����=�&H���bR��ܗ}s��R�� ��5��r�4�c.��8��Y�w<(5��� 6�t���}y0������u�i%P8+�?s�O̮�������T-������ڄ�7'�6¾r4�}q@��c�<∉w��!�3��x�h1������;���[9y�wZV]+(]��I��gNE��\W��sVz�_d���)�
��e��*`�fܡʊzm�L/oE����N9iޥ�ǥLΙ�OlJ�!��ݐ1�[�QܚZg5�i��$CP��g�ݳ�I�(W���	�ނRXj���ۏ.�ڭ�'6歓/����ɫL��aX�g3�X!�n ��ݻ-�mײv���y]���]�^�.h��.�����+�'~����g�+��NQ�>7��1�f<Ph�1��Z2M$2�$jbVp,��F����ʤ��)�����c]S���-Awq
�3�~�|��vɚ� ���=|�P���6C.���آ�0ڢ�����[;��Ô4�˨a�j��x��i���~���fT���\���-zb�핔+oܫH��PI�ǧ(z�7�'*N�`�T5�� ca����½�&j.�8�<�'*WB
��3}��{b�� �JFʳG���c��&ٯSػ����yl1�tV�m�W9Y��j��
1����;+i���n�
��.珚[�2E��ԣW�.��g����Gu�6��y㥚��}�:�q�4[[t�^�������P���5Źw��7X�P�c��wlui�(���#a��͡'�R�� ��k�����/|�X�i7-���n�%D_ m�*������i�� �"\�]^ ���C4��(�ed`����q�����C�����u"�;N��mtCfGEl>ׁ�te���Zm���6a���dt�����/��:�&�Jb�tskƌ�J��:}N>ysN���b��u�_�q�9��ۚ�L�'����U�pї,ڮae,�9�a>����6KX�k�Ҝ�#���^�m{�eh	��-Bfs~��@��b�ĪR�qt�r-Gs����P�yu�6�bT7���x�Y-թ�͑* X��f�7s؇��E2���ޢJ��)1po�#����"�VL�Mч�s�D��}3�0���ކ0������dƁ�\��q�Onx4	N��bu@ҙ�4;�+^�l�0���v׀�ȉ��/B]��	�1���X?1=�=�D%I~����9�=�,����j�*f���m<7�GFq�o $l�c�:d,�e# ;��r����J^g^����<DӢ+�[����)yl��/�h���<���ս*)4��96�;f��M�&�5��W�jꝧ�B �F��0��&�-3��|������P�.�\<O�E�y�eN�#`�N*g1å�_:�����0�	�N����j-���4�SA��'
%Ŷ;PcO�N�RΨ�]��ahb'm���S���л� 8�W:	��'L2Wh���6K���KO�ڊ�餴b��'������n��˲�x�dE1���r�)@,�t+�B�=֣���n�L��ԙu�s�I�&� �ȯ9m�jY;r���p��Sb�*Y?j���OP,�V{�9;���z^+�����]As"��u�ݘ&B�0R"�ۘ<���Oou��2"n ��l]�p�x(�+�Kn���E� �ld��M��Ow��*�X����.a��u���Ӈ&Ƽ�V���$s��rC�G*%��bS�L&���[m�u�ę�|b,��'w.h�us�ye����ܙ��t����!4��y�gR���%=�DR~ktʹ���r�g��,v`�t�:��^=��M�l3��֡=��2%�b��?�	�E�U��(�]
$v�
�+�rKڼu�*�Ōk|]�e�B������g�f=��]�|�U�<ə�4{M�H+a;ɕ;s%��uogb��GN�k�,z1n
��q���&�(dKvr
�7��Q�%����+6��}�`��Y�7���l�NKk	���=���H�;��=������NP�[N���zU2�Swt3k�23p�m�F���<Τ��v.lC�8������g5A-��w�U����
.��x�_��X���9~'}���*;}&5ɿ/����J<?t͌�NO��8a��ݰ9ކ06z�n|.zʹN��ER\:�Hm���LeѪ�����?z���Q^�7-Z��F�;���aו����ƾ`e�w�GD���$�ke��VyPy�R1���{�yt5�r��3�4��VD�'sΣC�����s�,�t8M�	�֓�2{�)҃,�:�j,�C[G�E"�t�������̂�죅q�lA..�\Ds�f%�u���Fe�̷a�l (6��d�Zkc���M�Cl�WmQ�|�CHLܨC��:gۏN]Kdy���e�?��Q��mO��l6כ����P��[{��xs�qb���f������S��+Ipdߎ#�]|��*c��R
t�7!����:���˛����b�5j%�m��M�
�ֻ�`��,S�	8:�=�­�E�m����H#2e��&�nm]Zyj���i7��@�� �pe�ڬ�7�¤��!h�v�!�d�X�+�RG�9�4�F�o)��;�����,��	�����'k��Ob�`G�H�����vϬa��Hz�)���9��>�-i�Գ�2/#;��e�d�Ҩwi��5�t��u����+�\�S�["�))�{�T�k35~XMߕO�:�~u�T����N۫ɞ���>��#&�X;m���S�-�ǡJ���;��Z�U�ტ%��U5dJ��;Sf���1������q�K�h�Cn�<\��;�9�;�Sp����q���f�(܅��m���!^�5;?�ף+�3�>���C��oLO����4��mȗ}/��C�ծ�Ɂ���=���t㩥�I.��lV��.�?��O���u��+3=>;�����4�Ρl���.Z�M	�%��_���L����5���
k��-Y��K*v,�2�N�j�q�ˋOB
�TJ�*�4e�dx����:&���f�#LF3+%TU6��yy�Sۗ��#������AeN��zNc���3���F�����e��锞�EUV���r/62�ws� ��$
��>b���~�Տ�3��]��1)�[�x�L6��6�8`W1y�u��,�U43�	�%�av<�A�Zi���� ��>�wta:<�@�,m�՘�^��9���.m��֭T�B����z��ƪw1d�J䶈2��+����x:�:�CF:ꄗ`�������QΩ���i�"˴�`�Xa\����k_	�%���p�Kp�Wil�-�6�k��)�u;�.^]���<ʼ6Jr;��Yde[����Y;���q�m��7�`b憣��;v�&��MP�&��;����.���[B�.�G*�3j�r�C?�'!���j�E�"��\>�h�{�J� ��1N)�{N���3�� �QL-s����I����{e͞'�qX���\���{t�яT�D�C�ܸ{���T�p7�P�J(��VP��r�aM+>�T�{[�ߐ��^~��f�?Vψ�A�lx��:�L������}xB�	�=�QI�mȬ�rj�b��G:x,����_m��܎�CϝB,L@��*�µ�8K�(cv�؈�gVD,�������V�_^P��l=}w���'�T�=K�˨d�a��Y����V���������G� �es�	�ӷ�=����)�:*�����%��9Ah�<�t�=�M�'��U7#�ml�V�0�=���5t:�'�H���1'T[9� �A66mV�g��&�w7�m�9p��e-���X�{(���K���S��G����Db���͛[��߀��Y9s�>��&���oB-2�<��Sw. ���ĸޜ,�ߣ�^�u+k�X%{�Yqؼd��c��٢�c=�辀��3u�^�{��@��=�I@;�5����D��TF��W��ƚ*�%0������yX�&���44�錺%f���F�y��UW#��#�l�Z�����K���83
�8����Q��-)���^� �`��_�� +�������ճ��"�=�����)����-�'U)����s}7B�<��T+hdo)��'��V�o��|��'�h֟�b�����[&0T�Z�$���g�M-����A�*���ַ�\ϏF�KP1ba�{���$3�+��#"���+ns6��K�El�љAkIҫ���@������2!����\�:��xsCc������n��K�HE8�Nǵ���z�n�}�0S�{Q6�-#�6��r�hOC�]^`�cl]��Ws���a��KJpXO���5�/t�6��DW:	̲O�2|�CE�b�%�����������[�g��d�Ed��H7���lG{\ц��$�mMԢ
�Ϣ�HM��p�hk���i�Q���L!�{��K���"�}����\�;�["����+D��wJ�m"��Z4��gq������Z�^J$n�E^r���Y�\вV�&��4���χ n)ۘ3oG�b���AK�ԡ�d��w#��d?u��B-*��qXu���̘fk�ф���0Sւ�>P�܆�v�Me�8�N��Ἅ��fL�ݕz�'G��F��ǘG�Y�3��D��w�ƾ� �)�G<��w]���v\��u6C|�z��7�?{��yB���91����bS
Je2�*��s�r�n��8�J��@^C���C�j���h�K�p�`�M#�^�Ж8��i����������u]&'|��'������z.&�m���30� ��9�u]�/�\3��*U�	Mې8�-!�wEŹ�E>s��GE��zՉ�2v8՗��ћ��n
b������3���1�0쵼�����	�D����K��	1X�3��	͛�ч�SU��g��i1��>n�A}IC6�bCe��C�(�/y^P��\)n?\����y��Bn;��&�#s��ޏl`�c�`'�.J뗑���0���+݁�T����znP��� U�Ů��`��}���C�ŧ����Myͧ�zc�h~�����%<2w�ۖ��u��7-Z���dD3j6�Bº���X�Sv����2g5��7-�πa�<�qcY�� Iܣ#�3I�9�CoVj��7J��T�o5�"�1p1�c�q�p���O;�t�n�%,RR*�������#��2
94#~�LL9 (V~9���{�ۓ�ƶ�=��_e�I)�a��=Vw�s0OIY��#ҽ�W�x�(��ٵ`��8)�f.�N�9�u�؆��qV���a7�z�u��2���ٍ&K��V���y
����F��M��fd��?ԺC��'FQ(c�����{�)Ń����Jo2�E���]
,-�;�/�v6�V���͂l������	�F>�@�{t_ ��unD�e5)�}Y�zP��~\G���2Y��+�l�W$43Z�E�<�L���\ݑ��i��+���Q����4˰�n��k]6t\��ě}�b�J%�+�YT�~ҋmh�mQ�\E�&���NYƎ�� �t-��ZTM�H�-�bv喹~���N���6�`��>Jo���Ukl��skZ�M���O�;�ZѸ�?���m�I2�284vb�a~u�c
Q~E�'P�����V�v0W�	7���XswKӝ���^�C>��!���.����Ĩ���(n���r4�7fq�wcm���;j���4:�r;�R��Y��Ȳ�M֙��4G��B+Lⶁz
�s��_�lf�]�ʭR�Zy��m��
�U.54�i%��,V�t�}�0a��������S�������$ѧ�BhNWG[�x�B%�(m�$��p��1����W�����0u`�2椼���[��n�ù'U�{F��s�	��<�bᑾ���V�P��̉l6#;�Jٙ&M��=X��iuӷ�=ٚ�d�c��urU�]��LY4�/PBZ�����]��і�k�A#�eHmb���\�p�oO���MN�ɶ�C�����(�Ⴠt�4���L�ԛ	ך�$R�SZI�ނ����|��`���Qu�h��(աo�#�)�V������`�.��.���OB�l�G�:w"ȤG �:�yN�VlYSx���>|�XP7AM�N�� v�ge8�-���
0Ar�b!�b�*���ťa��}7rՙ����2^/��E����3�;6�k�qwNh�+q�v���4k�N�jՂħ$JJ�D��",�����D��;v'(u�$��5ҏZ�\�p��oxa���q�����X�	О����k��Vp�*�]͸��%�D�p"�F�
�ݭ� �}�ֹ�a�U6����ՙ���Z݊��Ԩ�w a��,���Amj�� �F���X���h��KǙ����.�<�p�Ut
7ڷ&_}%g,�p^Ǎ�7i#����]�D�B�sW<rn��.`�:>}�x��1�ZWCت)�88�}:7�ҜҜ]���Z�y�F���#A�u�t��4��V�m,���kw\qǳ�y+]N�k{Z���攻�gh�{LZ�3�S{8Jd�h	uu���'g�޵����B0KI'V���C�k�ʠ{z�ͩ���͂ ���Q���HuK�=I�Oh�ﲲJ��@_,RC�ɇ1@#��X����'�PXE9@�v���h��f�wVYd�EYj�d;^�M�7�	3�wk+KF���B��gߣ�ȱ����u�1{���W���	�5x%g;��m��Gܞ詌�n��b�.���Nm*�n��jn�J
!0��V�ֺr�ʓ�޲89��V���2�X��Á�yD`�`�9+	��rl8P]1���{t�׍>gH&�!����R�Q��3d�x�V���l����>��V�ŋ��Mr�"�J�� S��v�*z�*
�U�#��w�����)]�r����ޤ�M��N#�$�*ucїʬci�U��N6�_k&n����mK���#�`�T�АuY�)�X��l��V�#G9]�U�T'v��mW0��r�N���J�;ݕ���d�!��'d}!$'6�=Դݫ���҇㪻m�X��P��D��jT삒��Fd8&S⭨����<������uzy�%Y+Sy-^����{�XMo8��#1�B1t�q��b:f�K��2�ϳ�yv��� eFu"tq�͢33H��'*c���;�Y��Ӄ����)�̀�7�Q�]���xk�!qǔ�!V�2�z_iqJ)!�jV��
�W�;d2�=c8������=�Q{�3!�Xv뫞e4zYdl��l���6b-eq�%�ג7�é,4N�*�48�8^���ݗ�n��SN��޹��֜o\�u�36lr��hr������7��>��+8�M:q��I�	%�
(�EE�q2-���"�
"((.r'uįqp�
8�)9r�r����Y,�_Ow���v!UUr�VդE§A"(�s",�Ȭ��Z�.�z��Ep��um+�i�2kŭԇw����蜨�5(�
�S("�B�[���)d\��H)�����p�;�.˟D�m�\���Ԩ�dr*�Т�.`Q:��7Ps�M=���U�:U`T�"�Შ��5�䓇�G/�ET�ip)0��/2�L����&Dv]�$D_0�p��7���.��¨U�!��G(4J"�D�\���(2�yz��(�32���q�9�C_w����4��TЉ�Ш��e8E��@�&EOOwg �t�!*(�R��N��M�'Ba~8�"� N_�Q&�����u���n���k�O�Lғ��<��@qe�r����b��Ւ鑶_W�;��7[�yJɚa�aVԂv\ɽesQU�}_|/(gL��`T�������ߩ輀g��	T�m�gO^���f��0���Y�z��	�-��3��:�B���m?5	pp�c�~�2;|\Χ�#C��h?B��|%ز�T�h{�a3/�1��Haa���nqć���Y�܏gv�n�����/�JV�ƧQh�9cT��	1�}�.�����mx;�ϏZ]������V�2Ɖ��*�K�n���u2/xN�L/�B��~3�'}?OK�<�:���UJՍE�z��qȈݛ�pp��;ܛ��q-���b��N�¸�ʤ������j���yfE�Q����q��V�ټ���t'"ӌl9v隆��A�=jR��j�h>�I�j�r�6\��}�H�m�o��%='������W��íԔ�N:t�FnCVb������<���3TPh	�v��J���7sX6��[.G\�{��C�LϹ�y n�����c�h�ս�#Kv�����z����ir���[�$4U�����:�ئ���<�)��������e����|.��v7�Qw~�&�q���!�;^K��4�5;�J�,�W�tt�r��%�&oe�iV�F�ғ�w�D�Xnh
]�ݤAէ���g7G6*�y^B�Ic�sw6��H���	�C�3�M�,9R�a�۩+6㑑�{|��D�+!7���wж7oVO�� ͞�G>e|K��)�%m
��W�5���}w����||\��@F�����:���s-��?F ̀�ʍ=�~EW�yN߹G�WL�cGE\>ׁ�tA6)�O_w
���P�q�s�ԇP�gD�)�n���S3	��QR�vy�^N��:|L1��6\�`�G6�F^[�ΰ�C�BܷҬƝ�O8���Z��U�,��G�������e�b�(�������"iY���М�<�ɔ��Q��B�ĪR�7`ߍ:{��4��Fxc�=DK]nm�beL^Z��j�����|�,���eͲ�%�N��h�i�6�������<�Q���:dh�rz��7��.�zǆ:�pV�e���c� �'MML";�1�t4�J�/�<�0&5��#\6�<e$=߫��.�~G��~������RkQ8h8�j};�p�-O����TX��g�/�={�f*e1z���UɃ���܄�f4�^~ϸ��3ԕA�Md����s��V�L�^�)����J�`��Sm	�y��ɖ�:�u`�n�{b�G�{��*v�&h�oot�U�_��I��Z���vQ�� C�wDx�R�`�{f�%L��.����ͱ�"4�\3�Í�/��Y5��rd�\����*ا���ojo΋��햮���ÛZo��Q�YI	���ve�J�����P���~����]�������n7v�s̶5^�L��:�-"K���vHw��p�_sZ��d���E:ֈ͔S����X�e�h�l�Uc��T��V���z2/o<�4M��_���C='mj.�J>���! G|�J�i��U�����{Um��S)��I�6��j��4��j0:�aZUR���2K��d�3.�d
4D�D���uv���ݪYT��(�	����I���S-���m��j�1Qqp1�1Lhmd��#��j6����&F�n^��^�: ��B9R/nbS�UB��Ԫ�տYَ���?T��U�M��w�H�A�þ3��ld$�-�@B����ޕŨ���m�������fX������U��Θ��;ō��6���ʁ��#�q�J{=����=�u9��L��"^�7E����ڬ}��L�+���Ě�[P�ף\)SK�u�©�����wH�SwO{��7Dr3⽉�yI�jǵ'T���oG��t���qy��B-Rv7b����OH6ua?x�w�\�Һ��#�C2gZ�X�˶�$\�ZFA�EH�0eH��awy���f>2��\y��+22�nҊCs/e ��ҲE�Ֆ��-E��Z��R�Mp��[���@�����X�����,�+X�CE�wm��}��{�ܧ��c`���1o�#��k%)ѷ�8�S)���'x\��h��@ր�d:��F�5A�;�4t�ª.�B8�}�l��Hݍ���5��j�'ѝS�0tW1z��Q��p'g`fc��-����SI�ɮ�v�O|gq��Bu#¦y;�FF	S4���{���W��_�!��&��0�A�	9%�������u&����v��&�=�aE���-*���uQ̄���81l�����B��%���X=�Y��M��մL�I�ӻ�E'�z�钃�c��5f�B�꒎�',�p۴�GQ���m�W^$��*^��ޞ#��η���B/�G �)xx�HkF]޽�I�$]�<��Y& ��AFv𲋘BZ�T�O5�t:��V��	���IeP�e��e�M�q2Xj}~�>@�jַ�Z�:a�2�x�s���X����^�LRuι�?�E6$��|)�u�m�^����;<{O!pVk��,ų�I�-	A6��v>��incЧ�ߒzG����,i�P�4Ah?��s�����������P�T�[ƗI��.�'M��rp��ǲ�Wr|�M�鎉�$�)J���]��=R��!ܗ�^d�*�kC�g@Ӗt�й� (-��G׋4_S�ذ�h^��'�mu��ē����f�{���]=�V��}��7�	U�MC�A��}P��k�?!�~p�K]Ɓ{��J�i��1�ӨM��M�5x����aE��u՛��jD7/7@�����>��L�a��V �4f+(�$�O`��`�ON�vA�Z�7$���=�^�a�\�]t㩥�I.��lV�t�~��7�����cZ�1�}�k����B�Jy���8��7)�9F,�!hD���Z$��v�y�����h�y��J��!�E�^S��)�c�л �I�߱O3����1:��a������1�W�޽�S���N��}'���w���zO#���_�"�#"�е�m)Ų�J�_2N3��'_4>���ܞ�2��*�R�$B�~
��}���t��!*�C��up4j&tЧ�3]8h?`�3.�Ѭ1Urⁱ^{b��Ѐ�Gy;8�}{��,rۀ.O<I���%�5�4ij��-�D��z�e���a�]��Q���O��a�}�У��J�=�c�+���9����7�c����:�h4�*�6��*w#ħ�2K1e�D���ڤ�g�˻q����-8�2�`���;:�h�L*{�:4Y��]��.���E�P
�#y����| ���cڻ�.���}�jB	��]��fT<��L�Ϋג������|a��Aye]�ꯪ���^z�����-��x*[��������Y���Jm���l��m��ܦ��v��G18��Ծ�e��ʹ����t������W�`\y�6���k��2��QI����T]P��;rِ������ܑ��5�ڮ�{r��D�X.���h��&���171�h>�B;�	�����.%��꬐�ӧ������q��|)m���r1K1zvΡ&
LZ�f���X�#b�q�<�I��$v���A���ң˸��x�,&�6�9[X��)�>�!&�ǟ1�&z؀�^�WKE��r9��˹Hf����c���)�?g��l�f�m�3q����_#V��p�f�1��3��<Nӎ����c�y�/!�vL(q�LS⊔˳�ʹ�+-,��9&����R��4[���T5�'�luS~, :%�oj1�m�8hˊmW0�Q���s<���P�᝻�g�z�e���Q-`2}n�&#_���$�j=�3�
%J���E�F�1\�E��+5�"]�=���/�O����q7��c8:�O�g���K�Q퍞�L;�A%� ��~����'���z�ԩ��O, \�BW��=���D�s0�0�q�1�mMq���u�K�\r��݌Y�O�@�ٱ!\�ݏ����+9b��z���f��H�^�Yi:9��	��	�X�l�{jS鲒���fh�Վ�)��a���˘� �1;����o3�����6�c���S�PY�U75 T[Bz ��:��iT{΋�5|)��KFt��t�I�[N���݄t��E���k1Ȧq^����F�%y]4=9P��"4�����\�1���0�W.k^����ƻMsQ�Y�����\`c4�����ʝxb��ֽ����zz's�n�^�+��.-17	����c'�#Q<l�C�	��Z=�(0��0���Ix%
���:�	��L�l��Ʋ�W��(5r��4I�hk.�Ô�6��]2�Vך^N�pz�OgG�9�E?���)���ج~FVE\.~��ӉL��<v�/�Pǳ��7<�-���)ީi�X�CL��.a��6 �B���Cl5���擄��B���6��"+��.�6+�(���P��+�jYp\�5%i��2�仂zd�sǝ��G��Q�zY!�����xL'�̦Y� -:��Z�Sa��=�:�RqnhhōFɎ�Z�+�cn��:�"��Zf�0��6��q�����Sn�-S�923�]�B�D	:s0��_�C�z�!�g��7ch|�M���@ڛt9?x��-w�*�iZ��p��;��eW:G)���GG��l����/ܜ�|��҃�Eޙ}�@�ĥ7r�R���']��0�988^�]�tqS�����7fjn���$@��Kj���]@o��꯾��	��xo>�љ�b���%a��#D��u?�]E_}����_��ʂ��I����09�v,U�ܭ�5���c�`����Q�^h�v�Ȗ2;)\��q/";�h\��Wv�<ۘ�7�_/WiK�)av�6������Uj��@�ƽ\)���!�R�V�S�es���]��n)3y�/Jv�QC�sr���$�B�ۨ�f��45 wa�#�ff�o*���rS	i9!1ƽu�tw��B�h�mX�ψ�y>�P�=>R�bZ����,�϶3��bM�O|��O��[=G�5�P9���8��鍗3�R�Ϣj��(�e��=�,�-��
<���?������ӯ��밈f
�u�	
0��msG�I��_F�z�F�����p�%[+z��2zT�N��N���6
�_>���O|�u���H8���������F����z̶�+m6�]��7b���?L�gL�-�iqp�!1/c���}:i�,�؝U���ܲ-k��Be����ގa��kڬK�t�F=�I�>;�Nf��j:�1��;H����l���-�ϝ�p
��M�bku&~)ҙ%e�اQ@|rft�Sy����8ܺ�
ETs&�3YZl�����DI�Q�'��]u�GcOHᵉ��n��#!xXJ�$��{ݯ%q����C�k�V�q�H�wB�qV�ƹ]��_}_|2;����6ݒ�>�c|�k��Mz���ϹB)xx�HhkON��I�3��Ğ�Qj%-�9�]���B2E�v�1Q0�{1�Y��L�\!y�dm������v�z�:�N���Wc�^&FG�'!�v��d�V�u蓯`���E'6�P����<c�E��d-O&�mW������$ПG(#%�#XE���uB��v�!�j�ͻ�q�w��������R��v�5���ϻ�rĽ���#ǈG-��F�{.����ǝF���n��<�9����.������*�P�n�2���;ヌ����6��nS�_�� ��N���z�u�F�[3e�ȿ�ֻ唺��kK����� ����*�9�:�1���g`)½0����c�}#o���uB�.~
�<y�3�7:�Ii_�'���܋g�h��Zr����2�	�=�{u�`�)�:N�wv*A����џR��މк��)�[9.��oo�-	��(�Bt3��0[o�}f��q����u8�	ż�^՟ChP0Y�%(|��Wp��������mD�jO�VS����:�32�[�]�B���r�Nǣ�P���˯���z#�F㨷���b�K������$rj��E���X
AI�e�>v�x*�����pY�s���ܔe>�H��_}_xLk^�arD�o|��5�[�a�=`� ����cj8NK:ӵ����v�nMfE�>��Ҙ��P��U�v 걋�]Y2-����-
Y�(96���! �m.�OH��y����q���Jf���ק��n�`1:]��l��y�gL�%��0��g7��������Dt�¦
&Z{���^�xq���S"�¸�ʤ��)ʟk�bt��G9l�\�v�'�\�؁O*W=K�8��^���j]�� ��PCj0!���w�gbQ�T��!��D<��6vc���:�,����U����
��Ҭ�qL9�zS�>�/HDF�8�M@ާbm�w&Ѭ����w�A?Vv4���#�X=����<u���'�bn�pi5�f_+n��	�j�����݄��@�5ǲ���Eii+.Hj;z|�a�&q�[�eב�MBQmns�DF�v/���#�MA��Np��&����ի�a�����s:^��)c���K�'�yY�h6J!��4�݆Q{�ue���S�f�m��Y���� _�����>��sƷ DJr����je�7ץ����������p
}�*u:)��w�`cA�yҙWW�2؜6����b��l��ς�K�F<�u��랪t-޼ʫʂ�'��)v�;\�����N�'t/�B��,I-�'m�����ܸӫƸg�wVwhZ��oGe�m�Y;i���8�KP�{Ί�m��$I�y�݆�OJ�}[��1�6�%�64r���]�"LvNm?�"S�un^��/r�殻fW+� �Il�wN�dtg��#p6#(K��5��LgMo=����fGW�4S"���:[J�������h�LDg��H[�;@��e],���V ͥB�"S0��x�J����^�/U�(�G�v�ȉb��e'}�d�b�:\��b]d���Gǭj6ˣc�7`=�+-]�]r�,8��X+��&����<l9z��A8B(�33{��ŋp.��/+U�;MP�j8胆
�Ű�tl���{�(:�F3W�����0��� �[8qn��C�gf��t�w+WܡxѦ��7[�tWl�/�<������s�1k1K��7uo`��<����o0!��
�.�g;\��3�u�O'���r4t�ԗۑs���%��+��4����z*�]��SHfm�L,��W��&����ms_	.�l���	e�X^�;FL
�V6�m��+��a�4]�=ᴻv��S��<*��=m�[���E�jRoa���蝣O���(�k�z��Ɯ�3�ϥ��/\�j��ʆ����$=A|�5qN�v�ꊎ�d����ݼ�+Ye)�\��D�+���6�>4�]\�r����_ɃQ��א)�ݝn��+�p��v�=5��ji�磠����of�ܠ4�C*�ܔ�z�:0��,�w#3��r����V�P�Uz;h�\䧼{�Ԏ�d�6m�xejFjǔ:ͼѼy6�uG�0��8�+TQ^lB-x.IR�(=��:2��p}�*A�g.L����E��IxNL!�QK���ST]s=Rn��@�}fGqpp#$�s�*�j��{�2:cJ�0�a�`m��X��
a)�=e�$��W��09����SJ�����p��+Ϲi�[�ȘEB��e��2dխ��S����N7M	�z���fN{W���K�����M].�n�7���B�%)��<6鮵|�6�+N�Xs�+����l+��D��ENo���nuh�$N�b�^T��q��]v��;rTU�\˓�]�)Ы��� J�͠m���&��+��#sc'4d�o��1��:����"�S��'e�Dɹ��Q�`�;IG{Rc�h�h��ϥp�Ճe�ٛN�iήp͇�y�A�z-�[S�P���N��|�|��W0k/ ����t���ܦ�z�5��O���>� 3�f�g`U���
��'�+�\�v�I�_w����
���+� �e�}F9����gYEO�x��\-��dp��C�U&��EȜ�wh藙�W.U�N�V�9G�'s��/5I6NIG���I
��
.p�Ϩ8�I�9�wwe�/��y.�S�G�EQVp�.�,���u*�^Hp�f\���]H��0�z!P�t�s�9��!Rw;p숎�YGד�Q^�X�gN�t.��Ο6E�EuZ���^����R��i���O%ͅ¹	�nC��G9G.U�� �qQW\���c��N�w*c�T�N����H�		��r��`��B��\.�	r��I&Ry�D���N��*��6�0�e��������}�h������6�en�@��D�K&K���*��`�\�1m-��@�i6��F�d����e�3^ݸ��p�߼�<=j,���[�<�|��)�c�~����&��=�y�;m��FKr�e�(|�|`�	��z���љ*Ò��� �	�Cu�ۆ�y��Os�z�X6��P(�n&a=��y6sd�D�m��XdΜP(M���� ��ǘ�:!�#�����m�SU�U)q�';Fz5�c��h���A����\�@��⽨cO5 ]�q�<�0�4�C�=M/!H���J��^�m����Z;'T������pj1�b���̍ܞã-�0���	�nv/��{1��N,��^����sMr����+U�(Sz��Ƶ�{�s>=x�Ib�"i`/��p�M�����+�";E&u�Vfち���l�)�>�v�k�]�����������Y��!��qB����Kb Ѵ���|#!��,�o��\���ʇ�a'b���mZF�x�z��O�r�'�aH`�E�;p�zZ&�F9abJ�Q�㏠j�cC�����&P���xEN�H�w�Ԥ�ݖ����h�͛%�7uI��_��F���?	����ۃ�?��[`)�U��p�a[��#�աj-�M~��oh��k�)YW�~�[��s���M�wP�b ��k5�~ޜ��r�����Gʑ�E�J�ϭr��t"MuM)�g�jn�\M�l����'�VHH����&��۽�ps>6K�鍘��=�z"�wW��ߏ!<бHM��UB��jƑT�]x�p2lX�����PW����r����҇c��2����z�H[V�ǲy]ԊY�\�5%i�bn�5 ���\U=���W�_D�N��V�� ��쐺:$�y�jS.��L����hWXQ�06%"'L4t��3�����Ѓ�up�0.z�CN��Q����i�PinSn�U�ԭբ1m_?���/��{�����:\e�Z8:n܀�����i�4���6�[#31
"7�9�W�Iܞ�2�t!���g�EzS�80u��X��C;�8&6_�"X���r�՘MK�6zY�̈��!"���Q�8H�z���~r4�0��x������wC4Tv�fJ{�.Vk�?u�9��uӍ^�SbQ�@�PS�u�*2KP�.]��n2�n�c�,y�r�;՛!� ��>rx�Qo#��lH��S��6��Q�#�"�p�#y����<
�.�Z3�|��c:�>�8�oY�rZ6k�J9{��g�zCᘑ�K��W%����l�|�9�]0�ؐu(љ�ճ�ۦu������yܓZ'H�8'�
���{kv�n�(%0�T�8����ʱ7�27V��M�Ce^��}}�%E���ሢg�>���d��5*m`�d��S��p:��{��]�Wq�T}u�B/�oJ�A�}_}_}���~�Á��<?�D"����Qz�e~�^�a��ī
�@�E�D$�V�\]l�l-����;܄�����}��'aȽ�b�[�~"�	��O>ܨ#:�i6���m���Cb-��_'nCTCh�놶I�6��%������2�����9�`���f##,M�}ɽ>�C��5��f��d#.���h�AGk��a�cn�"+V�к�%��
��SQ�u��j����5����y�4�蝜�������JÅx�Kɜ�e7����9�B�٦.�$�75-ۚ��aL�O�o\��d�pW-���Eg &w`�g�v��o{%;�KׂhT0ڍP�,�삋��쎉8��s�kb���إ=�}a��fwE��'y挄�ۆpW�=����n2M�PFK[�m�X�ŕU�U9�v%Ue]:�Ŭ����%���ӓL5��ɇ���ό.
i�A�O�.9�Fc����m��E�v�;Qi��ѡ�E'�*A�VnF�*�C�#%��u�+M30���Lx�WەT�`׬m�M��ϝn���M�����.�;����V��Mk7����[yn�m;�ʆװ�+=��h�=�8��K������ߖ������Y��֬�R:�Xp�0s�����|k��/g;G� =����F����k|1�x��"oz`N�B���z�|�T��kI40Vb	D�ﯻ5���?����9;�<�ؤSW��{5	�?��[���-�|\�Ǧ���,�m4��[�[�M+$�L�,�3�hL{�0}+��zןGi�vJ��qG3����n�C>XS��`�\Vhǅp�݌F�<�V�ʠg�+�_q𿛙N	}�I	��#Rj�+3�U|Af��h>Ȟ��+���ԇ��ā��Β!�Y�m��%4����3t>�sPI��`����5ǔD��v����Ka��S�������խƸݝU������u]��[���vœ�k��oA��T!><�
:��Y��^��==]8�)�&&�	����EF�.h$k��ǂ!�q�ڏgp{=ʤ��)���í|ʚΪ�����1�<s!����z��*�Cq�S.sJ`�ǒ~`�#"[4˞'���m���V{��:T��j���������H�nn��"���W�ꕯc ��15gn��M S�b�D���s�k�ذO�!�
�w�\��ܽ��S��*W.n�L�2�>�Z=�2Qa�G�y���x���$�*w8�8�����f�.
S63>�o����'c�+Y=�r��9��XT�W������7�  ��z�=ǃ?v|y��$v����Cj���u�?JK0}g󢹁'�����Iwl]�{ycb�u�5�ap��tf��v���+����ܒ���X��gP���-��-�'���%e��~8uՁ��N%�:xQ��0I�y��c�yCo�m>����ZM�5S8���]o��
�x�PS��,�H�����}0���,���S�f�eGE\>�<1K?=(����X�C��(%�����>x�g�wX_��vx�.�a�Ì�b��(�L�=�<�*8X���ŚJ}-w1�}�h��D�/&�}R�[�`&��y�]ܢ��A��6��^	58f�8��L-���ՍƲ�X�M���bq@�p�Xᯃe���h��}>g�=��P��I��ל�~qme?bv�q�L�:��2���qCP�~z.�O��� #�i�!���)�ꇣ���!su�C�$pG�Aˎ#���ߦf�nOa��!��.��v8��iJQ��9�=T�d���L�J��Vŕ�O+vI�\q{jsƹ�ѱ`�M�xŉ�5���_�g��|*���k2ܺ,ϛaI�e�Y���t#+ ��v��H7.�@��n�ud��	�z��vrN��S!�Nb�N�-v��;�Xn>^�ټ�����.s��$v���L�����#�fĬ���^���bE�:(���Ĕ��RX�����p���W�W����5��.�p#�9+��ؾ����=�� �8����g�`c4�UR`$n�F$+Nv��[�.[ ��W<g%���-ExL���&�J{��?8���R�\�r���g4�2g6���Yو���!#�SAdP}3�ɇr�A�c�gs|��%�[׳L�L�C60�|��F(#Ss�"������X��c��Hhm�"�X����/Y�����^hRJG�/�k�y��fM+b�*����-@M�⮅cެ��l����B_�
�嵷��,�PjWU�F��S�*��D�O�n����;^���z�nWt�^Y�\�'=eG3ƋB�)Rg��V�AY�=�\�$�6����D�	�L�
�d\���WSa���q�V���n��?p{9**`-�sp�[�l���nC@8zX���qtPm�0��Ja� 8Z�0�>�-D�[�$���Qqm2���*�>�gCe��j��7zW��qI͗{wՂ�TۻN^1�g&8�Yϣ%�(Vu�T'np`����Q��a܅_����2;���6^/c�{�M#8�0�%f�KS��U�VM���ڰ�"2q���>���ݷԻ��98��x�
4Vn?��x��þǍ�<�m�� z�NE��:�r��n��}|/`��n_B-��~=�&��5R'X���;��#Ω���rk,�3c�n=uo<܁~� x>n��G����"�P���ܗ\E)��饟Nq�KYmi`V��h/���U!`��݃R��T����V]S*�)��%2�e�
~GF�~Qq�K��X�Z�E¥�ݎ������4�æ)�K�2�a%�����@��Gq?\ԧ�L3wL��ఏ@�5�o�uo�:y��
��A�U�w�>^�@q��>-gt�y+{�L��������[a���i]��������Fw�9�43��vvF���=,�n�T6ǥn�:X��@ܥ*�s�O���ƟlD�e�X�E�p-�~"�|�3v ��Tu�5"���A}��.���}׹�#����B��J)3�钎�'��Ǡ��"T�2kA��CѸ�qǡÝ���S���.'w:Hy�	�K.��6*�t�F��8�gÍBO4�=��MYI-��,�3��t2�}�yl:�
���p��Q�#<�$]{����䉵�����%Ч�5S�8PL�^sX`ꆩ��c�*AOY5 �<,s�d���M�� X�+��j�"��h<i��NY�(��/���AP����[�27]�顙1��ز�����8�݁�o��2�`����A�����ޜ���m�3^E��G�\�E\w����a�W={�¾�v�%�/�7�f��OX鼃E�|<�q[;f����M�{��<4�,;^<�Ш
��C�.Zݐ��!�A8䘤��uma�>c�e����G��h���Ф�1̵�(�g&E�BP�G�v)�	�#��
��kv�k�6;rI��gq�Qi���/mM0��qp��_�L��~B=~p�U6U�.$�1vGp�����X̼,��v���ܵ��	�S�#��X��B��[�_SDc�oT.)n�5��-�޳5����&���y-�r�mq�\�M���FxC�\��\7TI'z^���4�e.�ey
�*Ϡ��>�w����ܩj���'�tkڌ�[����|��1Y)���sR �L��ra{�#��t4�>�1�q�I�w��B�R�e��Y˟�3ŹR�33��%m�2ۏ��~*kZ������ ���:��>��|�!m��m�����-&wWevC��).1"�c�e����i=0(��@ \�H�Q�d:�5J�1��-Q�\7���앨��iFd�֋�>�6J��ZX�42۪"�5�'�EU�m9��}ݩ譅��.I�C�B��5q=V�bJf�<}�0_ � mt�K��YR��f&�S�\d��NM����c��u����(r��F�иAS�v7)��ٲ�vt�BBć�r��(�O��;霷&�`�顂d3M�K'�ʯ����V���i�V2��$>��ݦmc^�� �:���0���.�AW)��[:z`����'��焔\��^q���Fv� ���mxӳ��D{u��nG�����ܮ�4�q�9z�z�@\��x;��N.
׏6�˚dZj�"�촅m}�ܪ��� �^B���2@��u��'�W��oSP���I��r�6\۪�T��DY�M�pq�VT�
uJ�H�d�:&R��p��c����5�a�y���9�m��œ�:��u��_��C���X�zy�L� �fMfi9q]�S?<!b�t�FĲ����-]8k�B�C���H��YBDS.�� ����sn�AeV�j���*��?J�ۀU��P.)^�e��s-g	�ŎM`��S��SZ��փ��(̗�����H!���f�P�󙔝b�d\�dF�c�[M��0�7T���1k��tg���9C�З!����<�i�Xe0�0���1R�ֽ���m%u�¾#uP���,p� /y�,]�l�����o�a�цؽ���˻́�;��7�z�ȹ6KQ�C��D�|��ۢ�s��`�}++�OHP��l����R	�n�J���]G2�O�����鳠��m�-W�.�6j%:�8�e4��nR�3��n�u��XX�uc�YR�y�/;p�����	�Ff�G0����
z�;9g������R���i��}�/�wk����tKD?#շ>�k`w��G�Z:5ȥ��lӎތN}j;�e�8\P�._��]�q��4C?0f�F�̣-��O����vqg9�ʥ���v[)������R_ �(�;ܞã�0�����mn�W���-d:P�MȂ�o&����VZϔ�R�˅�Uޜ6�3���>z��kaz�uW��_0E9]��g�B{E�Gx
cCr�`�wk�;\]�����tw1V����\ѓ��1r��A���K���:M��ƥ9�������P�N�'r�:�/zD�$�P���:5����D2h͊7�C��M���#͐XH����Q��y����ف/W��ڜή�y���H����C��A!��͊l�+�mrEv1xÑ�L��n��b�/�����j��O64� �Z�l�����E)� UЬ{Ս"�T7�I�СV.��\�L߲���9zE���B*g��dVe_�_�B�j%K'V1�G6q��U�p�m���o?����j��~��Y��)��w���@����_E�z���tm��y�E�x�r3���n�I{M��+/f!�6��ބp�qY/vw((�WH�*�q��^�#� cqq���Ջ����٦���Ӆ+��]�LM�4�e-�b� ��k��jm�3�z�6r�v����#�6���sR��7cqw��{�9a��%a@��N))��:��΋.+i;��͎�l�1�J�r��tN8�9cl����)Mc���V��m9W�2Va��RE�bROkU,�
��P��.���ɕo�jJ�Z~�I��D,���U��	F��%抵�8�Σj�'kj��U<C9Ԅ�I���9���#xmIܫ����MtOTW�r9gy;�7��ΝC��y
!���>�ػ�B"�����ไr��gg$�;͏m��0p�O�2*'|��ӵ8Z����w�*�/�ʫ�mIa�3D�xw*���CB�J�[�=G*v���U�����(itH>�z�A���؅���jF��%��pZ���it��I�H�1��طXr���*�VuY���{K6ƉR,�{KbS�=c�з�!]7��C�V����i-v�k��vka7�咍Y�ں޾��BE�����&snw��}Sr��`�Vk� ����Jõ�K=��zur5���!)q�F��`��x�Ǔ�]��kE��Ǖ[�U�H�S�Wc�,����������mTB�@.����lF]^aQö�
�,������Pܣ.�E3��$U�f��H@Tiv乐e��z5���{ϫ_a�q�u�*��`����^Q@t�N�B7wP�Z2̍%8�-[ww�`aLu�{S-7)��\�Wvnv�^�
�r>��,����K��R��\rV)S:��G(c���c�t�i��!	Őn��x��a��{r��A���jC����p�f���gsu���5F��c2D+g����NJ�\�����ڣ��R�w5E�$w[{����<�Aqn.�d����V�j�x6����G,g�$6�2e����A�&���f���N��t�+����+�i���EN�ؚ�ANCt��)�f���c[��;b�*G�J
{�ݱ�ʕ��U��h�h��#z-A��F�M]Blo6�9Nѐ<�ڙ����&��[N����״#�5EZ�ݫ�,�>�Pfu����s'E�������F>(݅���I�6'.y4��r�S[��돖��af^�=,��BRڐ�Q�o:+�j��q�WE��kb����fK��S�����L�K��]��1�I�f0��V\��pb�2c�:Msڰqо�v9�ǃ%�v� ���`�����}�� ����p;:\ܠ)���]su�-'XQ�6�^�u�W%v%fi�r�BpK�4V;�=�I6��WۘE쁞���\R�_hK�5���b��Q�o��ܕ���V9Ɔ�3�z<���;:��#fv�����?>{�+�>���D�t�*h�3���:�<�� �#S�E�Y����u�dZ]wvQ��X�b�aZs):a�8����fҋH�jH�\.9Tf�����J��8Ihg��fP����<���(婡�E��/"'ZN%�]��ゕ�U@��Nߓ9z,#�uDP�>���T�QUTNZ��FD�4�RI	hP�J����J���}�Q(�@�#L�B��'�iu
�D�ft��q֕AVFi=PrN�y�=�NbE�MX&e]B�Q�s�����{A��QZh�I�6Uˮn�H�y9]�)XYӍ9qDOW2(�-\�t��J�g~"�� ��\��)�������r��p�t�ή�á���L���۽�LНô-Uc���cz	��9iI2S���܏$#���W��UU_}U���{h�/����&B�>���[�0�����C�a ��ȕ2˟��׉���+�^�UQ�Pz�V�r�Ɂ^���f8�!�j�,��C�n���jf%�A�L���;2���V�ra`�K��u�Q��鱐i������,O�<!7P�	�����$!��5���nWX;ST����);�8+���
·F��i�~~�I|tG�i�])W�ᶲ-��j���W�j�oO�1�G'��q_��n���l��k�bΜin�75�j��(�7��%�l�ɝ���aS,�����R�j��G7-��څ˷�F,�h�Ua��5u_i�lML[�A:�-BZ��47S�9i�T��LwL�U0(��n\�3ۛ���n
"�c�3dC铱�+�>��e�>�6	�ؤn���`�S(Ntؖ��wN��57=���C
�-����?=�`�@i���/
uH�yT�_F��msG�����隉fޘݾ���m�ADo;�F��
f�לņv�w"�X��D?
����ٖI2��=�����p}�������"�������I���.�m���n��{����ܬz7�:�|��`����֊t*θ�sn���H!�5ٱNʻԣ��ջ��5�p��.��2���Uf�R�d��m�.詋�8oJ-���k�.���Z$E6���_}��}��4�$?P���s�#i���,Ą�mZF4y(�X��(ߴ�8 �iq��l8wQ�cS!���f�[P��]F6e�	�e�̙qY�>��Ja����b�WLlsӾ�k���P�ku����=@���:�&�ƫۓX��O>�*Y<rP�ì��T�!�6����x�Z7kgrq.DB�{נ!����2E2ɀS>V\�Þ�0�sW�j%�h=E�j ���X?��O���R������Ć��&���C3��H���!R����<�zf�Y�s���E��)2/���Sry���e��&Y%7���c㚲B�h���S��IR�7g�q�iİmNl���H��E��|�6x�Ӄ?x������j�����ñ�g�a"
i�}Ah���I��b�Ч�uc��Ը"�����0P��>a*��P5+�lF�7tUoI���w�uc��O�%	x\��)��\!˽y"�=��u��gc���s���N4����n�(mfj��i�����#�ty���2�c��;>��QPJ���7���u���Ė�u����ĉ�y�չ˄�����;;��Q���m �wb����:eH�`��kf3�4hUȝ"�fqaK����W'Y����6��o]��]����_Qh�k1���Km��M8��"{%k��+I�A�9i!�n^k���^��ź�e�A��s-���Ӯ���ޜ�ۧ��)�O����lve1�s	�^����[�Q�EQ<�0��5p�w����Y���+Gi\�x�'��P>��k;�1���Am�����sq��#��6U`�Y����vz��u:�iFE�Z��Ҫ��(�Ξ�qC��@�� g���c>���
��ޅp�n�G6*lϒ�U����&8��3�86K(�E��4:��b�0�("�KU��3<D�y�G�E�c����{ �����s,�c6�^�L#�By�e�8;��,��\I��h�s!��3ӡ����yF=���B}���ũ�@a�\@�v@ۦ@XJv�wE4F�q���/k�f�9�"��^ߑփ6Z��d�����l�v:%i͌ʠ͇BY�U��3oo�]ƍ��� 
��mvDH��%UYR.�.�&ܸ6�YSl(�}r�fĥ82�2P��uh�]:�j)>ߊ��]��PJϱ�_�PX2����<�1�]���+��+ӯ���.��9�:f��m��-I���j�d���$5���#�+��v	�*���ݚ?d!%v���:պI�����u�H�k�ӾUv���j+%��aB̙;7�{�]�ɠ/������f���]���єF=@�7���ڛx4E�����WX�g�>�;ʎ-c��©`��vXņ�U�}_of�c>w�����[�c}:ɶ:M��e'�O�)u��ᕒ6��Q��uQ���T�X�F��pY�� BR���'��@!���f�ܥ�3):��L����,ձ�3z��
-݆��1U{B	�󽴁^���5/	�\��L�Ks�~��u�1w�S��P����=��ǆ�Q��AD���QlgO�Ɇ9��FY��k���4;!�f�i�m�a�x�"S��!E:#mnc����,��R��?�_+N(�.ĵ�����·d�;�����(���ܽ�U��J�.7K�1j{��ʌ.(j/�@�� <���T�{�w#щB�����z ����V*)����uX�b��A���*�mmF���D0�B8tJ�gf�D�Z3�bae1��1d:�l�\�H��S�|��z*}����<��ͯ\G�ԭbW���X���.Wwl��,�R��xa���{�'T�猦G�E<ݧ������*�x�kN��h��Bv�cn�>jhz"�ڭ2ϟ&�D�j��t���G1��nY��w�����o��[�3~�G��}U1�{?z_�V�nC�������t*�Em�Jyv������V�tM߶}�֎���V���x,~S˨7���k��é*\�k�]��h*N53P��m
s��fr��A����qyײ�t�{E��a!����/0a͛4
#�������A�M�G����0��46�ZF��5�Sm	����"[F9a}1�@�۝["y�X@,�9�s�aF�G>���y�axSS���,Y9�2N�)\!��M��T��䎦ǁp#@&�f�i�0�Գ��{+f�>��J4�ÚV�U��i5M��MZ��h��W�*�1ԕ��(�Q$9t��C�N�ιs��"�@�����j�Z�B��pJ�O׆i�b�of�n����N�*RqJ��u��.{�t�MQ��x�VT�]�S�*K���� ��B�L<穊�O���G�g��W�p�䮱�wE�@��sP��� ܻa����tϳ������.;)I�YM$���	U,�5�V���cFV�H���+Z:(c2�j�a+{�F���æ*�.����H<���f2Ef�׭	��R��*y�w�tV'ђ�B����80u�v|���!>�`���a��5\踒:$�>��@��rޡ���	U�ӹ.��;^�����;���/MZX"�&d����Ϋ{=N)z^1���Lz�e�F����R�
a�"J�m;g$�j.�ޞ����S������3��.*E�^��+�1���V<�.�z�\*f?�y	/���s|N�_�(��r�ҹ��#��v� �%]m����KV3�B.'%��ZfI���H�,s�Ml�[x�yy1��&u"V��9�خ-�y;u������X��F+�F��}_xsw6Z&��?y�Ph�Hy��^�Ɣ&ϙ�B�u*�ٯ�*�z	0�yo*i"�^hU�^�\��h�gv��z����7�}fQ;{E�u�1IfŔ�3
'LUY������)����O��� ���{�p��C���H�PQ��6]$lƍ�4��_{5�:�d���^�FzH��Jf��s�H�wq{%��G���+��#�F�En�u����t�ݎ�e���
fK`��������Mm�)'�
;f��0LQ��걖c���L=jh/E?q�����<��3&\K6�)!�B`=��HkڬK�(�em�&�n�ƚ�Y�5�a5���^6� �H�D�����l6�%��r���%<��Q��wz��G5�H��{/����D6q�wYON_'�-TZ��@�������a�4޻�1�C1���{4nZ�RW21uE��Q�\G����P�P�T<���R�[�+��l:5��7f�ݕ��;��c�LRs��k�=K!�\�(�5^J0c��rH���9&�{���ɵ���: ��C�!���%�V��X�L���c��W�+�v�߬X��~�5eM'�|h*9%��� �C=�[C+���97�������\���;��@��>����y�(�l6��\�ngX'�#��{��j�F(XEB�m���U)��q�%3n����x�z�w�	�:>��v1��?)%�Rq�%��]B��j���9/�@�{*�<c�,.�΁��rW�=���nɧ@;e�"7R��.PB����H:�,YC�\�b�-`�3���U�������ڗ��!�s���eir/oT��6�B⭑jצ]1����`T����X�ϵ)�)v�K���!��y�{�A~���O��?V�yy:�E�orpg����J�m2m��B�y�_�QDܬ\I�-���
t�]�*i\jL���jM:��;[颮�q̘�E�.R��Z���x��ja�Ck�a��}�����9S�WB�]�T���7!����9P��%��Z�my�1�Y'���$v4�7�Mo&�a��#7��tT<,	�?'T���<��6�	�ށRXm3I���s˾��0��w;:����7:�0��˱�� ��7h�8:<����~�υ�I�bJ�M����P^���ף��)fT~�Y�ㄧ�n���]]�اW��~=I��6�,).x���,�s2ҡde6�U���7u�L9u�ܦgjsz�)�_]��u�	��:����{���q]�ݔ������ͽ��?y�Xqb���lz�t�"���8�u��եЖ[��*�b�o'^�<!�(7:9v.K뜀�8I���3�b��G���^��6�b�������i�����?����Ņ[���?^�*�Z.xӔ�{�kb��5�b��u]��ٽg�
o.@���F�\��1���N�4��I�����C㚈��"�DY�M�pq���F'��κj��a��riPe�а�)�sԞQ��sq�T�i�j���ː�Cظ��i���ҰU�!b�GY�T�z��
ͺv7�	��	�=�O���*�U2ܒ*܌K)`)ޅ򃺅X;y��s��G�݈�-nx;O���jth�GI��̤�Tyw�ݯ�܍ؕ<��3�Q��]���
\�<KHn����Թ��H!�v�}ʕ=�0��	�BӹUV�LJ��l��Ӻ�w<�K݉�^���P���2��~�ǨHx_�ݔb��L&�o%+&"�1uC�d.n%*��;A�Z�3+->P�Ó�p�{࡮Y�A��?oIs)����LHO�7e��oaIJ�)Z�a|��tc�g��֜P8'�p�䵀�>rp�,����OpG<(�7��<�����`��Ak�,��4��-z�����8oH`b�>��anP�[��6��T:�wY���meZ�����̗A�%����:�u.��Y��C�˷G[�糛�\W� �ml"���Q�ˠ�kF!ղ;!�xL�Yv�uq��q���x*9�P䣲�s&>ʻ�;)8Ѳ�5+����ڭOL���� f��i�L�N�����wRomP�*K���ϟ����p����k{�I�A�����)׋���+a��<�pV��l�ܕE�([X���5��sd9Զbڎ�Wr2;��ƍ�\8�;�ˀ��׵�����.���0F7P���� g�ZE�M�g�4����b$^�g�sKP	�vg��=@r��8{���}"�Ɖ��kٮt�DvIa �d�8%;4��~�'�QwAtbw/~�.$��E�h�J�`Ԣ���L>:�t�4H����MV/j��R��9*hj��T�>n��؀�W:�y:a�˄8�b�%�zW�Ctk�D^��
�����t١��;s�+T�{}�0[�eL���S#_!)��-HM�UЬ}V�'Bܧ���p�&�]:�ҖDV^���LNz���b���S=�P
���l�V5������.��������'��}�GVQ�4�Q(a��Q�{HdG �&��L%��!�Y��Kn�!�6��Y.�%.�y���OoY,m𼵠�s
�Qy0(^4Rz��i��l�	��s��4{��oN'���U��|��Cذ�.Y/^یܻD�U�S��MJb�^=Gqv+��Oi�m�<�
,eY�	�x�Θ7&��w��>\�&�$>)`\�YY�1�4��mM��l8���8q��g�w����N�Ԏ��\�֊���<<W><7e�<�1)��{�T�ܞ)}�o�"��i����`�G��p�u=y��i��Op�*��^�2�[Tw�=*u&�h�d�Y�P�nq<�Wj{10��������OxDN�0p/F8G��������yg��S�ד�q]i�# ��㤓jk��F��n6�9Ep�XL��K�a1[{*e�@�%��jULq��G7-�
r8T��t�æ@�O9��ݴ""�Z��0vb��}����P``ǜ١[�1�b��s-�C����3�oD`^�.!��%��c�댴�����}�C��У�k��q5����uwC�	e��,g��4���r��O��0��;�/⟃C9��gdo�SJo���ddQ�ڠ�k�>ԡ�/����5;�()�OA�Xga>؇����	�8��UD�����cG�2~�R�ѧ����u|�����g	�Q�ДR,ODoL�9'X#u*� u�#8\DZ���N�fͿUCP�N�EI����i��;�|��O������+S��J�gc=Z͘8hX-!N<}mtk�ݥ����=�s���UǓ]1�f��!5�1D��F��7��o7��oE�]F!K�U�E���3U�
	�@����/;�]��2�N=�lќ�����: ݹX�h�E���-�OJB�j5��(\���V�ps��ݞ���}��b=�(
�,L]K������4D�G��I�t& �n!���j0��K"�;IYc�FnkX�#L�2�b7����4䨳�.%�|�?e\P��7]�J핻����q��o8_�!�JK���:�L�����K�R֭=�.Q7k�M�Tu����ū&v�u�s��	Si��
̘Fr�:Юpq�M�h�<zSg��������\H�Ԯnr�{��D�(gU��x�Ŧ�͐B&M̛����$�����+C9���<�����˕�9�x���n@zQ���|�ww���\L��T���	`Pƅ.{����X�ZX��xn�;X����Rup�Q�r� �,	���&;������\ї�u`P����ܶ�K�il�W����*l|�ɼ&�G���с�9�v|n����c��Z��u���J�F��%V��r�Xn�e1S&.��u��/�=�!c�]75@�{�l��]�ا	}G)]�t��*�D��qt�ޞ}��ږ]�������W'��ʘ�6.��|R�/�{���Z���F�]M꥖�a�p*���w[� ��1⩻ �j>"Z6�XiǙ}�t� ���c��O76V �5KM�\إc:����!�S��R*΃,�8���`��l^����6�:ԩv�:7��uc��8V����5j���sY�W��]ШH6� ����(_t7u���(7�(x;�y����l"ٴګ���ح����ҮWw���v=��Bp��������Y��O�ѷB9�:��E��g�f!�8�X񜢁챇�O7���M'��GD���eS#&;�+�����-�9"8�j찞$^_.�����R�	�d�f��3tHH�NCy�1��k"�3�7�u�z�����:锭-<�r����b#�jS�07mw�����lU�V�$tg�}]g��CM**,�b�:"��S��ӟ�vX}I9���n�����Wϵ'	�5�{ ��]^�Sys��%���I2��j9X�����-����T�����g�P4�
��u��o�3�#`�R�:4aJ�6lH�8��W,خ7��[�,f	pk�pVމ�vS��I�)�빲�]�E�+-�3X�[=fv�+v�eq
N�?,�V�3�Y^X�MZ�3-�/:��둝Ce��L�޸�[�4![Y��-�m�}*c�
fYP݉eL\*���dU1���gX���9�������<��r���V &�Q�@������T�(�"�I�~I���e(-*jlN⸬�$���
s�Ra$��IӡYPD��
�SN���yP���VReU�w;�O��q6\��H8�y��XXf*�;4(�Ly���W-���<�NdEAT�N�4Y�� ��99�T�bBГ���U�e|�YAuD����0��4Q�-�sм��iȾe��ףH��"����F�����㇇)��re�;���ד�H6�<3��Fy�uC��"���vܨ(��sj+���ܒtY��\�OC�>�WDWwe�Y�ܞK�X���������<���L���g���l���TE̥
���r;�q��TC�BH�f>"��K[΅�9�1ȥR��J�G��\p������^y2����}\�2T��-�t]܄/"C,�aR�����?_���Ď��G���s�ح����gM6���rI��L9cq�IV�*��C)ǤV���U�����H�6�%(A5���'^C�
i�\|^��{��&�vƥW����8b�v�M��K�����z}�;����W��~UQ�M�]H)�/,�<-w�]���4�wis�Hѷ�3�G	6�ܸ�ҵቡP:����$\�ݐ�=f's�����T@��$��֦��]�YH�)Z�W�CH�o$���6-�U�
�?��;�V�n�	�}�Ԋּ�|NFE	iNؽ��@��\��|2��
Q{�Qi�g�P��4�[w���؍�=�b������j����x�˃��N�#�O�>^˂��J�cנ"���}V�K�X��?NKBiU�YX����Δ!� ��y��p{M��"��#�Z`�l��R+��H��9��.������W&����uq�5P��[t�SmCD[�b+�]��馗��fk�b�M�`˔��t�Q�q%��k.��!���rR�n�Љ&��2�t1Gx�Ҹ��!\�DD�n��SDAW�!��5%�P�Կd�k�9��k�ۛ���Ҁf$���{K�U�>>Kl��W�j�������1"�CD+����|(��^E
nf�{�3Wwc�ayHV��Ց�De�%A�7#ʔ6L�]+�9�i��Z˷J.�����xۃa��z^e�I��V��9���
f����ۜp.��	�WP�6��;x���+�U!�g{�xzn�;�$r�c�y<�u��u8�	��#A��*k���XgO\CH�%�C�9���h1�w���G	m�(c�zw#�ݪ[��W�� r��T�Jf�����k�����i������2؜��]� ��ihcÖd3k�> ��f�cK��v����T�Q*/�/q��� �Z`��Y��OW�
�l�k��U:?KIf�ߣ��i[�[��K��ٖ�{՜���qhv�y0AW�6�W��5<39�0iCT��#0f�SP�[A+4�]���Ι�4B���H���a�RN�g"{Q&S��8G�]��G���,�*a��<Ln���澓��ެa^��ˠ����)�\��6���&�ù��r��n�.�]DZ���'�"�Fʗ>Ly���S��|^��k�\qÛ�-Yܦ�knA���3���9�s��������Rw�h�|�`�7=R+a�9\�˹d����P1���J�M2�7�tǔڼ�N9�����7q>�d�`�ݹ���C��q��H���6��8U��+%�0����WQ�=IZ�&�ru3��;�1�bӹ'�v~�Wϧ]m����(��uL��yb̫�eB�#�S�#��U�05!׫L�;bڃ-��a:e���c!Q:X�fd�,�����wp�3]����l�x�&@��GsL�u��D��s_W�U}�_k=�ޞ�|k��T���t�uK;.�D�w{ ��a�l:;W�\Ŋ������ݬ��}�2K5T��|1R��/��(VX���b�&���2�[�y�L��')̭�p�	���Fv2�ڮa`�%�`g�bv�}b�lq���'����� �k';����r���	OOL��rs~۟ƅP'U�q�����j;�e�8\j�͠��5�ar�g##:�kE�Zmn�4cN��C�9�QL�;���$ڡ�t��!�K>)�n��u�bxҡL�{��DK�GHa�]���^�y���cB�[rh ����:����9��Mtڽ���35�4A�\��b�gp����F+��2/���ˀ�75F�/m��jz����JH~�C?$bF�=�� ��4˹*�<�������>�ť�n9A�����mO����,�zܝ�]��ؑi$6��r�hOC�,�!����:��e+��k0ld��vM�v��]:����^��L.}��i����X��!�na����f;��������Gk����)u�`u|�'(�v2Y9��!�;	g� Z2��ɝӾ���������^� ՇkD��kҳ�v������D�/��k�ʜ�Z��.r��ꔣc�����!�-<��5�>T�=���e�5}j�����|�8�~����xmY���0[�FT���U#F&(f҆�L4Q�A�77��h]�"KIyYt�[h��6�&�B�3�.YH5>�nBn}�6�UX�G��:�_H�~U��6�.��y�5�J�wMP��E�Q�;��`��X�%�w��H!�mmb:$�i`�pꄮ�8�}�%��c������T�nFv��ܪy8�!�����d���3���0A��X���'j/y�~R���A�����E�+��=~��nc��,hK$�O&����4�A�;��@������ix�.ʞ.�����5G6ג�gC����-��Kv�j..//USF�X}l���w��Bqge��tm�q���sЂT�r�	ts�$v��-��D��ˬ�U{[�mj�
b���GV��O�l�7�:��P5�QQ�ءnoX�:�KC��W]��ҥ��˲���Cl`�wa����I�(8qB�3f�6�GP��Q\k�21U[���'W�G��n���\��h�wl�;�� +��F��-fQ����������7~/�z 7Z���ug��(;��Y�G��k�M���G� ��af�;���ԝ	�MPl�81ںX�OLlv�r!wݸL*gsx��s��������s�r�^�r�����p=6���&<�����N��������u���v3ߏ@|u���^�`��Di�HA~��TGsʡ�v�5˸�{�څtg�\��~���e��� �N�c.|1���L���]+I#;(�3�9; 0o��y���+2˚+��Y0�a�M�i��].Ā��,�C[$�~�(�qY@!nш�w�جAD��Yp������y����N3��}�(�	s���S+��D�遵r��ѧ4z��N����9�]���'�O��l�\M���%���y���/i�fC$�]���X�Q0�oc"�yZI�ߌ�s�ʡ��}{R
y�n�X7f3�4e�u�6�5��'��}�a��ĹC#�̎�W8*�c�E�׆&�G�T!��H��l:�1:�o39������W����1&�ɊG��-yG�;@�J*�RQ����!L����v"Oe<�,|U�Si6B�#s`�ц9��)T�zT�r���+�^ժ�LmO,Vq.i츗��.���4�|���_�C:B=���>������n�%�9���ҟ0�������a�h["�{ܹ��ϴ��H���j��]��o�2K��yL0X��A-u�/l���=�<�Y����{���.zcV��0���#t��m�c��æogV��v�wَ�uJ�WӅ쾆WGs�/J`m�}�e��e� 
�+ꪣG{O_��S�nT7��4F8U/���)��_��tS�ި��.����3�W*B��+�*�k�^��J�wuӎ�v�K���C�ݵ��6/�{�����t��W���-�:r��>���+ڪ})s�W���3�7-�d���	�O��;��Ɵyq�h��]Y��٭�A�^�F��'���;�x�~y�^׽{�ҀFO��A�3���H3�0�4KV�%Z$̨��^��Ԣ�='���b,:�m��n���:�#M�'�%	�s�Y�*])O��0����fm}W�e���������i��a�I�-�^2��<�LD�1Ӌy�,F������Y)��7�]������1C��H:{sk����4��g��'0�>���^�n��c�U��2*�:�ڢ+ҵ�%g�5��WT�����v���d��];q���]��Af�w�m��)�3j�r��b|�א�d]	�)�Seꂞy�ؽ��y��leR�T8jcIB��מ�I����{n�����$�z+��~�W_�[��5%���J's�%�m�2��:��{#���HxCJ�=J����pz�EN�J�
g���3^���`�k��A6���l���ދ�R�Pf��n�tK�W��M�Rs#��JTC�,��v��5�ܙ1jOi���[�P^W+Sn�T��ﱌM/O]�Q��ϼ.<����Q�'_��ڊO�VP��r�aMX�b@��G��(��8�$�9���V�L���C�e�]#s4�t(gs���0�k,�j�f�7��JE�E��iMD����F�C-�#���z�@{�	��<����Y�:xW�L���%>D����.����sW�2"�����\��od�60�q~7pǓ�.9�͹4�!��B/vʻ�'��o3�n���L�Գ_�x�<�T{uP��&o&6���,��%C���0�9FJ���!�L�6NF�vc
b�)A�)�9d�-�e�<6�:����90m�H&��Cb@'O�+W5��<+�7�S@�)�b���d˃�6��X4�G^9��	^> �k ^w��W]|�َk�Pv^�2���c��L�Nn�����%J�keˡj;�e�8\P�._��%�����:-���I�<��b g���Q��$Lisu�FOu���VP£��R[!M;�a��cu��d>�%�>�!��1v_�zǘc���c��ji��U�^0f��<.ۢNO-g̎�w���1�7���D���O.�����VCMB� ��F4�X��H��b���N[����T��l	�3F3��ۄN�M��,�U����
�A%�>��,|�5�s
c�9�Z7j��:�6��5L"�L�2��K���p�p���}�W���G5�Cs��7���3�b���K��������̟X`�&uѱha��n�@ܸ������t*d̋L���<� �IUJ|�fe��{�Y��D{`�"!F��m48F{�E���7������ɇ�`�r��m�"�0O��`�ͪ(:3��
%�H��΂��d��M庈���/9��g�{V���Чcv�8�҂s��
|�CEϱM��T��xF44)�4q��MUx�)����`{�	��+z㚧n�۵)���0�)��HM�UKM�g\"#i�ݛ0jsg%r\�lSB�1J(K�����)̉�mu;��r��E£W�V���w�;�X��r��޻���,�.c�l�FY�ن&B�0R"��;E,���<%���T�B�d;n�`��MۅU2.p.�lW1A��=\;KU�T�~�"�����a��T�r��G3�B��.�Y<���/)�
T��ª�h,���&n�Ն��:�����|�������4~#B���d�/���2���*��nf��GE�%
�
R���fv�$5���
�����d�S�7�or�h�!v���t����t���7*wQE��+�k���g���*p�����d�{�u�40V�Y�uL���T�*ًw�������F9���45޷�<B��wM�+�`}�_3B^�⾯���+J�=���������(n;ͥx?d�W-��^DH%V���]�;��LXU溩c)z�@�^�d�a���
���O�D&ޘ���ܥe��>�R�ifE��34ɍ��Z�����$�'���rKV�r��zC��!�8�(��0�0``��٠��ę%��՗���N)���5�S�&�g��:y��U���:.���c#�x����{t0ی���o,wiд�5H֠:�|�	�u�׬�5�jܶ�!�μ3א�����E�j��ډ����K��mt�H<�Ⱦ(�N�⌶2w�m�=0!��/\e�£�Һ��Ns�H�&�CE�B`���ێWW�i!%�GR.�2WkmJ*�8�wx`�95��`G
�Џc����������^��h�ȇ��C��Ba�"p�t�ז^f.%�y;
d
���t�p`o�-
�v�0���L���'�]�D��в��.�
E��Ѥs�qnxA)�4��[�7�dU�bK��o�#�]|�.�b�>�{�U�HkŦA,���4��m��\��lL���u�c���v��J�:��т
�:��o���v�����cb�Sׂy�)K�g��	5�	�CB��ދ_]s�j,\GfoD)��lV>�4%wC��e���F��N���+�T�o\v�ig�k4r
9a�t�u9�����}K�'�)f��~ĭ{�(A�P�ɶ�Kn۰,�j����z��
��f�x�l�*��r���/p�	��!�����n���ߖ�R*���.)�9��1�5�+���49��LZsM�yz���[۽��e�k ��Q�1�J.,9�K_�8�.�7�R�a��S����4+�_^�Zk��Y���4>��C?8G&�@ff�C�I��)�w��#w'gb���x����~�.�q�nM�04�_W�#gZn0�E��Z`���09u�W��N�%��#u.n���G����z,����]t�]���`���-�L�Gz�*Zt��7�@���@}|搖�OI���h�r�ೋ��<s�d����2�,����2���-�I�'K�z��Wo���]�h]�U&c�9z�|�=�8L���F���+�x^���?K0.܆&�>Y�_��uH�㔦�q�bq��	u�e���MW:OA�j�eB��Q9��B4b���|�A�b���]�C�)�C�sC�}���`��;��Z/�L�� ٞ���}�W��ʧ���i�^�W���]hO��J�<k\�a�[Ja����W2uB�O{��	�k'�S���Þ�[��E�z�'��è��+HCQ�m��^:��E��
��K��M�:;mrC��F�XӌQ�rq�y:ΌnB�h^Ӗ�Ch;��"�mᓢ�H�E��Jؾ�6��X[��c��s�|�����XIץc�{�1�Ǭ��٫��,"��pѣ{}��V.kwϺC��W������q��ef,[����L��Y0�-)�����#Ht�d�Ӯ�lYj�G�_*��7m������܇n��G�'��.�
N��b}�N)��Z�l�ے����]�D��FJˢh�&7	��[V^ud���Y�������J�kv�Õ*��¸��]���=0����Y���E�\��@�>�#%�R�)�Ǚ&����;�q%zí��
ç.;��]0�7��� vX2��Ĩ;kB{"��1�,����_o �bܔ!\�O-�8�JM+����Xln��F]Lī��[v�X!�]L�=o�[�;a��|9)���]il��4]`�	Lu>���i+�\Q_�]�,�+>�@�O��º���DU7J�G:#�P�j�'���=�ңה�U�ٕ��eޗ��@��Lf�Ĕ���-��Uo���e��/u��;�9BJ�5k*����(��.�ps}]@J�E�{�ⴡ�w]�B�7+�Gls��� "r9��f�g]fΩ/	wu����D��nL�*t�2���T�2�᝸�'�٪M���+�;�펎E��m��3]�m+Y9Sx�,k�Y�o(o^ad�c;�[F$˭j��D�q�軑�¶�l��Q[������:�\�jR���k�r�)��%��6^q��G`Jf�mk�G���p\�V�=�݀��S%�
hZ��uj�56=�M���rV+�EYڔ���*U���z�L�ɚ�;(_�������;�*d+���r�M7,Z&��*�qtZx'��Df��u�iDxK���u�ݵ:�#K�'A�N+�P�F�5�� %�O��k+�X��Ya�ɺzPr,!m�
Se��La�ǹ�5�6�w�����۫:G��W�e�]���v#�R��7���*�@�3�r����rz�
�u�d��ܳu�[Օ�$�0��G?G4Rn엕oy��-����5� &�C0G,���1��-(^�1X�Q[:x��k6X�ZM�P�WL)�t�WJ�vfP�k{'1$�d(�y�PI�&��XFK�5]m�k��J��ċ���W^���6p�Fg�
�9h��ՙ���Ύi��/\u�A������9���Ȓ9I���}Qgvν�m"���}1���
��Fm7�+o�dVf���vJO�q��	#d��F��˗D�P���9r8_V��5�Gt_B69-�<��8幋,N7���ֺcwfw['3+�>��/S�$1�K�m�_Gs�'P�B�>�5D�+w�;~4��wr~I��aQ���RC�q �C��#KLTNXd]�ULR�7��T^��s�J�a�dH��%��U(��T���|������d�4�*��uJ�P���[�%EW1��i�gHA4����*q<''#1+:�'Ğ~Q�OǇrC*�[��\�)J�5��sȢ�O:�q+�M�7*���=��縡Ⱦ�t�Ȉ�q�LSG�E��KHy�&s��B�,MF�7b�Dt��Q�I��Rg=%�㇆���f�S�fI:��Eʊ
/we�7K�W�aW�v��9�i����9L3�U\��y��讈y�=[�s��CZQ�k)R�M��w7�P\r=�)���!����|f�D0HU����w@��((�
 ���P���%���`�x���X�"}sWMF�z,g�{-��(���$��y� z��'`�Y-S�Ԡ��or�Pٹ�-�{��13����	�*����	/	�s�J�����r�<�Ƨx��h�|��Xٻ@h�ݏ?_l�;X�[��7a�Pb����=�}wCz]�i޹,8�(ߴ�9���`�C;�����5lul�����/�p^�7�.Uǳ�~�-{@��?�p4�*�{TS�-��&u��
�9%9���Ǥz6�v���⛖�����ˠ� �!�]1���d��;Ed��U%��2w��S���צ���=&��=�S���C�܇�Mf]c�^����p͗���ʱ���Y.���x�Й�]\�
��~b�e �6��Cx&e?#���AB�w:	���,�j��;�����ܴ%����7QkK�Hh�r;d=9��Bl8�cQ�j�`�m�<)��C�f�-��zC �FĮ��2#���il^=}yCn	��w`6�bݑ B�|z�!�o�+�./e t�ܥV^my����	sX�:�ͧ�e�����Vn������xe�E,��e3�ǝ�"����|�Φ�0�^��e��LS��aa�E�(VZr C5�ӘgccG��T��9������	L���ï�h�^������˹Å��&Yg�I�0�Yɜj���q��2�̷A!}B͹!��r�<c�t�c�y�E;cmq�6���J�+��ܼG�&p��f�B[�bf�<�����y?w�T��u���̾e������3g/��M�6�`k"��)���xL�����S��s�Z��t2�~�e��-Q�	��>��]�6F��ɪm	�NZ!�s����b�J\m��t���-|����*�Upt���`)hF
���ć�`�Co=C�s^��R#��x�j�������yB������H���JfF��{�����]�;��|a0��}B�1�S͜�6��RYnM��{�j��_�x��|z5RZ�]4=9P��Q���=��,?�
_�>lj��qs���![J��\�b�`�|�j�L�-�P�f׀p������Њ�1���s�Xk4J��%e8Bw:�>s�8�̓^=;��r�A��TP`��oa�o��Β����A�	���+�Qf���l9�jY�E�A9���{�.[�,w����ٶB1��۵,���Q�H�L^ǁ�4%���Ը��ʶ�Je��YBKERl�V��4>_��?�e@�?���4���֛0a(uÀ��T�uW�׿gڳ|[�� qR��/��.�o4�VmE�vlm]�t��{�;x_�a֓Rq��.#�U���U��\�ƫQ@%�w�7=+Y��k�u��t�Jո��������=��|)N�ZI�*�
�=-��r�׋��� S��ف��0[�~��%����b��SM݆m��
Y��~̃f(�+L����f���[�0�mB��E��	�[�$�M�#by����,T�9��m���W��ɁB�ʧ���<�PE�IkC�lQ�2::������B�e�d7Pw㔋�s�0*a6�*����K���cΉ�N^�'ך��N�Z�Ϸ`�L�l۲���,gz
5&ZN'щ:�%L���aӧ�?!�o�i���Ԭ��5@��;��ͼ�R�ѷ���ܣQ���u=<����m@9�MsU���x��?�;c@=��������f�]L��5��"z�*����k���8��已��ը\�u�d:��h���������cC�^�~����K��P#^���F#����Q�ҼMV�-��h��2"�?!�9�[�}���}žw�T�ڨeC�a�X��cw�svDY{�L��<�d�|�jk�;j<'X�<H-���^mi��L�D]ݢ�Yk}� ���r���R
es��3��ё�DJv�����=��=]Y�<^�����~�)"��j�үF$����]wo��):i�=�8���7���)�e��]#��M�&��B���盇5ؓS�k���q!7�sV����Ő��],�8g�}@�B�w=�����J��� ���h����8=�O5�#�#��F�v�b!\!>����r����0-Z��&���.巠�q�&�ׇ�\Gr���]!�8�t2P������~q`�^mϺ��.Wo��1�:;�������Z�rV0��5����[�
1�ע]K��ha�b��g�n�˯zn�o�k�7W[�؝^�"�.��0�%Q"�TԌIhd�#�]Q�ήR�P}��Vw�i�K�/���H�gK�A��h��Zi<.�z�F%Qbsϊqˌi��k�^-i%�,s݂��m�d�	�(~�F�[��}��:$��&):�\�G�[m�Ec����� �2�
�6�vuJ��DN&�FI�^��#,�f�Q���ŭ̪Z�
�NN�/U�����Jy�VLl�R���\:v}�^q�	f� �G!����F�S�qe��xq3�Q����ָn�W�V�4:�r;�]cM��s�.�[����0y��j.��0D�u�m�J!��Q}�1㲫��������zf�|,�]9�hv�K���G�m��`�t�Gx���}n�f�݁U�rG���u�Ғ8������B�VlBv�6�~\���A���ӆ.$s�+��s�t��Z�U�]-tE��y�B�t���æ[�Yl[��)s�Q4p+ ���G\�V:o�Yek���m�Q�:��/�{��
.�����;.�{\���M!��2%�_�\?ԟ���Q�e��tk�GYV�_Ԙ�7�Q3�����j�'�gW�	{��A2�Լ�{���ƅ߉T�m�S�x���������aݓ�:�Y�!-��+F2��=�e�:%�u��OѦGis:�hHȶ⌇�����v{�4��
�3��o�����ān��wi���c��oW���@����d_l��J}�=!sE�R�qpi^Qe�K9F��9���0��C���L�t�Wm3k��	��sd񎅕98��ӑ�w&���{�e���a��<�
3�'}
�������S�#����S>��U��e�Qv�Ƹ��d? ���2��r� �6��*[_�ǜƼ��d\uT��E
YX��c/[77��e�8�K�8��9!wq���,�a�%6J�h��~���{e͞����GZ��*"�d����?�+v��ˁ���u��a�չfPe/~/)��VP�~�X�mQ�MQ�����jr���r��vQ���Ǒ4�76|���
�t;Mz��0}�v��X֬�Ԍ��ս��LC_C}�=�i�0�V���εܞ<�\�X���q96>�ft ��U���GYBLk�+gb��zc�1 []x�Ô�3�Y���=���Zp���0S��uG�!�:���KȯP�rT-7u}�W��Xw��DM��/��f���N�E�;��m�m���0Ȃ�����2z��b�w�,����8�t\�ψ��F�ؼ{Ur7i���c븦���$*^r%�O����D�HDe�Օ��F�g�A�T��tS�2��	O�B��6ę����.�"�y�J���p�����u�[ʽ�����Xa��yc7ЃCoL!��<�m��FO��e���r`�������jFB����ǖΰ�B����wk1�=��Uv2⅛U�/�,�3�$N(�&B�?MS��*�D�u�S���9�	�.Z��2�����b�V��oF'>�ύ׌�j�Ԛ��h�Vfw@��U%�kTt���c;��vu�S1�͊�e>��[�	�C3U��m3h36۹����1H���UCD�'������3��s�[
L�pV�THH��lU�#���}z�e�<|���(���7L�	禇���$8Q�'g��A��/�&F��tp�-Ol��am`��:�ŜW3�01�J�C��r��{4?:���x�qRၫ!<o㕙,WMfN�z`�l�>+���+o��E�3	΀^"Z�� �$�)Ah��R��+̙z� �v���# ���r��N�9|�s,�4��/-#ڪP�2��b�����l��9|�˴��H՚���*�ĸD��q3�}]��o�jS�����329�0S�{Q6�-#����SfG\�r`Gfvf��8���#�L>#���E��$����0�a�P�m2��Q�s��Z���`�)�ԑOr4�`�/�������ے�]wʩ��
�d��ŧ��ys3�!����Ͱ��[(�\a8bã�;<����kű���=��l�G���\��*X�X�4ˬb�oiWt+̒�(�+L�{&=$fr&�؁�)�{�c1k,=�P�;���0�-ּ��\ykȽeu6y==�M[�/' ���i����Ҽ[tp����j�}d��͑ >�<���假gxܶ��m��Mm)T_CfD*x��íkA�0G��0k%�֭�cݽ+�Q�S��2w�tV'Ѿ��z/ɇn��s�_d�Н��3�i��/�gwGƸô7f��)���b�Q*�>��l$����*�a��Jp�.���p�q�K���|���$DBm�2۸��0T���1T�Aݖ%q��0VdUH��ܾ�Ǖk��M�EI$��ѿb����@ȼ��k�ڋf ��B�n�L���vG�g�{XK�D��T5{e���Lb]^gm�s�2oY|rō��r��\�f�CGq9���>V*)�����7��fR�2!O*�̈́��΋�����'�\��[
.H�˶р3p-�$���O�\>�9�KgGCi-peU�_Jb�p^���b�(ѕ�Q�ܿOЗ�7��-��8y�U�~=�G7gg�r41W�.�o2��Jrl��z/>�#Z�:m>a3��{=�MMz}�P	������U)��0�ƴ��`a��}��nt��A�-�C�}N�亂�'�u�"��՗�ә�/3��l$��b�[�N���~�Zߔ;n8��ݤJKd��d]���%���j蝂�W��._�W}��(::����&¡����_���C�<�����6%�e�i���rq��G6 6+Q���x�m�!�F*�T�gL��K�aZZ����{�l2)D�9��z�og?��7%�'�Ԕ^R�f�Q"�>�E:ϕ��M��G0��^���.1$�9]�5��Rf�mFo*����G�0S�`!3��Gr��9�Q�\Eڡ���h&y��_`��ys@�lBb��f8-�mmq�'ɊN�}5E�+�Kf�f������7Am`�ٹ������N���w�����R��m��a���T��-�לj���u[d��Mvp���,��{:Υh�\ ;���c����Oo�^�B��6z��`:)H�M'py������MJ�Qr��ε�Sk\ۻ�ZO��9hΨ�^TA��<]���B�*�Z�B���c��H�[�>�S��%ۣ#�);<�r9R�~	E�'���Q�iq�i��^����-ԹMCz���>��]����#�O�?��gA��HgL'�����k��x�#7��E�^2��YCoʖX���;V�0w���.9�� r�b�.t�v�:���C����P�)u�����k���]8�iv�K��
�n�A}ҝ�Q=N�a�U�R�ZqUO��H�c.zZ�k�t�t���-��Ԙ�9w̒F�B�\{��������~����>����ٟuKWqP�_'�xǥ\x�kƊ�(MZޞpIE�NV�§+�
�������k��~�>.����̮q�4-��F�Az�%��,�l���ʳ=�}���:� Aʧb��PZd:�=��<yX-^P�m1���g"A@J��X5��'�V�hl�؉��z�Np,,�_�ƴc֙�1C���y���ٵO
�=�u�j��*;Z^��0�a���njgK���}��^��:̓ƽ+�߸F0�Cx][[�A�w��d���Z��u.��'��f�O++v�:�V�� �ơ�����5���̠By{F+:n�ms#�E�Ƭ=�k���8��uk[�8�����2/�c��{�k��\�X��ڋ`��'!RI����`)?Wm~廩��7p)��X*Y�T�u6�}�<(Ø�j�z��i��&�н�5ܥ�W!� �2O)��l�ʝ�[lckF�&�r�w�y�V�i�1JU�K��߷���)9\N_�oY�﫲L���gl;�� �S{$�l��S�S��v�\����aS��`䲧���]T�Z�'#wrv^Γ���o����q�Ʉ�M��kJ	���Cj��8��c���T~��,f�Un#v���43,9M��!h��k�<��tR�/���=���܉��7�+v�[!Yͨ4���ې�0!��n��N���WОyG����h��$L����]{��M���ۛ+.f9�D�fCg������f�[��-\����p�p+�&=�wi�b!�o:�Hy��!�m B�p�a�撗\v����$����Hc������`^��&nDO]�4�.��o��1P�1Wg_QT�c2�G���Yb�dj��~�>��IUn۠��f]k���oz��j���
�"��K�Q�\-opU���\���iN�n
�֯����7v;��=^�\uF��-sd5cm����:.ے�)�ܫ�&M���H���� &q9Gx)��Xb�q'���V�-�,k)�D�nQl��=y�:h���M7�>�ruk����zU>=R���� ���`�3��S��:H�P�@���g���-J�>�6c����5ݬ��Y�G��S�X�qnoW��%�;ofb�݂�(".���v��e��<�p�nQti�V�u3�Bzo���=*D�����t��ҷ5Y�[e/�M�ա��uX2�u��\��B�Ļ���ʆ�+2=v.U�_�V��,u2�-�vc���M]1Kwl�2���5���w#�e�)�JqWk�;ֻ:�U�'�Ǆ �S��<����j{B����Oiԭ�>�n��l�sv.�u7��tXK��SE�\b	#\���nICq�B��M��2*p�w��˩��0� �GR���&�mL��9R�e�5m�����X�R��Ȍ_G�uwت����X鈷R�*Y��AS+d�/�^e!��`�|)�s��O2.c��N��i	�ԧ'T�yy�\��kDbj$,m�Y[Ձ�ޮ��
�E�.�]AD�g&�G�|Ɏ���:���4��B��³�b����̩x��9VN���Z}��tF�4Crĭ5�����oq&�vk��#����5��N��og]d� �Z�GkL����2W`�
ɶ5��7K��n�q��2������)���S���T�tEv ��{0�jMpY��2�ﷲ�k�zUe"�����.���ew�<�[�NfG:U��Z����[ݭPl]
mm[��B�W�t@��Ɵ>�}]�,�� �7�Z{��j=��̥�IV�M헴��9�+�����q$�!�+&Vkt�_N����������r��[;�WLՎ��C`^�oU��gAzk��Qu����)�+ն�3&��5s=���r,{pGX֭n�R�e�v��f�U�#�"�F/�f��w]�Z�8�F0��'6PF��CB*����,��@�h�O��\�J*-NO��wu�4=ѻ��U�����ñ:�ת��;0nu�}.��S��k�W{WO���[�j�d@ӱ��w���J��d{V���o/+�b3N�
�"��!4]��F���`j�ck�J�97-9�Bw.�ר�)u<&GK���^wR��D���W(��,��n;�)G���q�ީ:�"y�������R9>��iX��wv�֜깋�s�wI*�	����ۜ)uոlL4w	lA8����m�*��H�΁��f�,4����Y�� Lf��9:���J2�����u�O+T��U�N��R���-�sig+��:Q��xb�rU�X$� �A?��s�r����R�E�Y��5��Ӵ�:�{�����P!�{��H�vI��/[|�޹�I@�D$J�����Q�U�Ef�]+�p��459M��)�I#Zt�Ӵ�I,��J{��N��ܨp�(](ɚ	ȅ6�r�yY+K�b*G�ށ�#ih��L������$���C�'s�ZٵV���-3.��
ڣ.D�n��D��*]bnaD|�V��Iwp��QJ$��<���E�qʳ�!��L�+�ʵ2�U:c�^�ey�r*"�i(��R"��ZDE�i��x����������A<�ZćW%w:%���8�NK�p��D����7P�p��G��]�O5"�'IUM�Gy9AS̉�Y%)��硇$��w4B*�C�[w��h���PP����Nw����=r����{/K�Z�VR��ɕ��A��y�p�cy8\C��!8Y{�^���j:u�Lx0�I�t�ӐF9r(�2�����ݿ�%�H��>ހ���2ޟDj1
�9=�o��>6��Cj�ّ!�uխ7�2�W����y�L�ϸ��@qr�F�qiC�VԬ\�͵�9U�&�kt���A�9:�-_��i��0���?FpΆ-�.0�cG^�:��SS��s��4��Ѧ���=���q�$JI�?����'9ߕD�����������V&��#qH���[g�ILiqe��gޔ9�MT�-��|A�o-�Y�Z�Au�Q��<WR��΍}�28�Q��o<�I�5	|��K�F�]�@;^H[�-A{v�WE>��e)��lGy���m��+�]��xz�;��ꄮ� �\�V�<��,ߞ�r�{�k����x�2E�	7;���M����I�Z���6��Veb�|�[-v�b���u���c|�f���l���q3��HԕGV՝sK�ȧ�u�g��؏�ٕ�3F�]����5t����7�l˥ѝ����Һ���*N���6����%E;25\�%��k��������"y5ﴒ�Mn��+Y��K�.�;�eL�������]i�ZƆ��M�����f!���b|*ˎ#7� E��_v�4�ST��J�,���~}���9*���Ɣ��a�n��.�eϏ=ndo
��w�U0�Ӝ�Ye��_n�+�h\KA��2V]�'���Tqٓw��w?��8��]���9��0:ә�å)L��8�6����_osv��FYS��fv��\�C�"��.~z+���3�S����`����&&��T
�Yj/���mxrcR68���C�pj�&nkZp����Ţ�Ā�Q낪��o5�M8-;<Z�����oێO�+$6ٿ+���/�`�y����FM����k,ݍg�7�gda�dԃ(���	�a�݇	�ڗ��
1e6g�a�ut�\�E6&�Q�<̜��I@ז����t�|��,c�2c�'�B�Pp���'1>Z݌�e�cn�^�I�$�S����!�E��+�C�@k�BJ@��T/u�5�
mj��%`����;EW���*<��t�K�K��E������� kd��0i5٫��	�:�7�8���Ȼ:�G:�;�b�:���꽹s�E���e�����7�(�Ҷ�=�%��WThN{vEoH�r�j�j�j�Si�P6�l��$��RQ�`�gZI]K$j�h�Ԏ��!�!����|��Q���WU����]mo29�rC$Su��O�[���/v��5'��ұ]fd�Ee١*6�Ns�E*텕��
�R����h�kzk��x}�<��u�
�����	�
ކ���������q�y�G>IA�f� j_j*�sb���]F�lr�p_gH���0�HBqn1f�������wU�[��׮Vχ/'v��,9Mr ��r�4�����������י�+�ۏ�Rް^V����
��A����a�u��#I�5ն���ڑ��"",�h���oQ�e�j�}�#o����vYw�gޠyT�$��yn�%�Y�'=�eI��=ׄ�¥���ТЖ�������jj6�^��6�<�ї�hL%u3ͺn��ȭ�\Ɩ��1�k3�Tz�����u�.q����{&��t�
�����2U�4km���2R{zk�����بU�C&��7��q�9�CÇ��.�;���|&	ױ:9�j��K3ktRhoL@���#��S���dӳ<�����w�)ް�;7�����iA&X?~/_�1�H;���e�{���J���L	�m%ܺ�\����4�A���ް揹C�p�Ca3�
���Ǒ,�V0�}z��X/�.2p�a�U�G�j<�TҐ�A�L6�8d����+�H��B��kQ����<�$���h��#�m*�N��'¸�Ӝ�7kh�cq����S��Cv�Unl�{��IHd��ar�63�km�P�C�K=�کW6�\Di���wLY׋SZ�"�i�:��{�y7�eGv�z������������j�upM5�W&�@����Kljg��T�����os����ޥ9���U�y9`���G���|���u}s]�zd����v�v~�D�	Ou V��ɐ[)�dg�wm�D�dc�Z��Fc[���w��m~��0N_������g�9�/x�'?�L�V�Hl�_�k��z�x�6g����$�Hl+������7��J�P(��1�Qh�y��By�_����{���a�f�3�g���ݒ�PĹ�g9L I�~��̑N���tާO&�]t�f"�na���7�7v�<�7�F+.���Y��_d���$+��I��0�-3A+d+9���:�97���uTɞ9�����pB]7
Yv���Q4����c��.�R�2�9��::����u�ri��[�c5!�q�Q�W���O2.�D�R�Q:���[�ާ�3�Ee��oR^�-��͘!�y�y�#�zg%(����:�����m�\I=�������$�F�M�C6� ��ii	�y�u�!EM�k��=�U��Y�#^��Z�m�E���E���냣W�Íp�I�K�}6���jȉ�ts�Q5;���tv*r�}ĵ�3&y�?H��dY�'�*A�U��6n5�[r v-�������u���ǰIT���_��kȓ�n���-�Z��l����!a75���7�7u=r@�r	�m�ϑ�wj�?	=���#{����1�!���-°Dٺ}Ŧ�v�ϫ�P�"gq>�C~\���8e���e*��m�V1��Y/.��fk٘�^���bj*f�46���f͑�3�i�n�1�)��e��9\2�ߪ���͈���"L:2�87m6E�{r���V6^�D��(8�������6�]�|���U}���w7��=��m5z�U�H�ӳ��.1���S�얗���BJ��М�=�l�t���&W�����Q�L�P;@Z��f�O�]�ڲf��H��TnSV�j��9�iͧ�~Ʊ\'l��ok�h%u���sK�Pk�j�WNFdȞzݝ��13_C�k���!��4�����%+t���dػ���"%�l�ި1���4cUT�{��[g��l�坥�8�-ҷ��ƶ��Ȫ%� ̹���3fnoZ�$�J&@n��fa��pޛ�i���[ON�sk���ѻ��}2���o������[�fv��L����T
qƛ��[������5٤�,��v�	����q��w4s�3E��;,��/2b,�'^��9j�:�%4�r��q=�/|%��W�������Ps���\���Y���ǥ�yU�w�8�`��u<k�̷[	߮-hYBjVgBV�\��n��P��_�΄���^�V�ٛJ�}��ƹ���v��\ތ�����%K�`v*
�
��4��>�"�;���!Bs霱[��=�c��k��D�6u���_߅�Cȁ��.Nlan�XI�ơg�d��@���C�S�F�-�ɇ�����F���7��=��}۩����P�Y��x4<\=H��wOD�t���A���?O��ug �U�4�;���Rw��Ul')���w3v��i.�hql
��e����//�� Dپ��`����f���i�ؤP)K�'����^V�������䳋�6p�[}��"��fp3O�@�F�rqP�d�A?$�HT�{ؿq70w�{�qG�0e��Ck�T�I �]6B7���I�u}|�U�R��*�
�ô$����PƔ�Wi%~�i�d)k�\��W����(�Rxp�����]�����7yB^���qf˟�e�!��(�����������Z�nI�N��w+��������=�f�Q���1��w.����rB����ޙ��K�0�UV�)~ƛ_E���q�6�]D�m^�m�Ú�\��[m�vr�1i�R��!PZ�>RVD�M囵�a+웮����!���뛛n�O�H��[z�[�h^���;r6])�:���v�C�13�o����.q؞'�1H��y[�9vȮ��GQ�^m�:<��x�W��Z���s��IU�Y*E���Q>ޥ��j.m�#o���S�� ?;�<͝�����j�U�����VSvF���q�W~�
A��1W��C\��3��Ϩ�f����F����7ȫ"ַMۍ'LgsU*��4�A�gq�����Ag�5��k�b��a�Y�:[�_L�؝��hhy�kukw�6�3ҕ2;ڠ8���<،�����	��Ҕ�t)]��͙ק͔ǵ-
iHcA����d8��ǣo���-/&y@�6n4K��QS�Q~�"~���[O�i�m�]�$�d*�Pf�5뱴�z+��V��\3�i��y7H)!�S4{U:͙cp1�ö��h/�����SQO�i�7�^�Zhw)z�9��0�h��x��Kʕ7Tt]�j~ vf;8�3Y���O��E�'n��ǈeq#�WW�	�U�[V^|3}5��#JBo�X��-t�Nx�.u��ߠ.��Gc�9���K�C��:��k��d\�ڡ3����ƞ�;Fu�W^&ٔSe\��q���g����q�:�X��&�X;%���F�����'2�ޕ�fQ&6��l�7���[��GO�iM�&�(cT�;��rx��)�umޓ�X��I��n�]dw:G�b�Բ�+�]��XQV��Ρw�r�x�[gw�U*���E^;�r:zht�R<|��}I�k��ʙ~K�̊:��_�+z�j>N�75&]���`;"�}�����c	.�ۙ�S��~�x�u�A��Fu<\Y�Ǚ�Hg�Z��v���{�I4�X&9m1̵͠��Q��&:��L�˔����ge�Ý��ƆGG��EP�=�ұ<��l��2���m�� �E��fk��zzDAF�����4�n���0��6���|�����]���-��9�/��7o`|���oLF�M��i�,7'���[���/��R%-��E��ֶ�t>F�R��s��n
����e�ljAAV���U ��Yhc�����A�IZ�����g2J��ӘƤ!۰�N 
�B�2�wK2Np��"���i��Ω|���%b�����-��X��U��D[��s"cZ��w뻭|T�ن ��M��!�z���]��<��"�%�Rc�|��J}r��[#���;m#�5ə'�Xs>�m3}R��e�FE�{E�5[Ǣ�H�qH����\�n���$�	�3N�]ݠ�q�ݝ����H�j���h���vUxf����y��1EӋ��`A1'ox���4M f�t���K�G�ɘ¦&�׷���u"+p�d�usݍ�{��>�=	.<Z.}��?l������K��e[�S<��D�밷�m�k�fMWv�Z�AyRҕ�ڮ�*��,W<�H~�������gq��VVnp6Uȴ�;#����U�Y4�{nU�t���j�Z��s/m�A��(\a;��h�S�Wj�U�4>��2��(�'=���U��u��z��0�٘�E�S���j@l��k����8L�K��	WʗuC-�n��.鍈�� �5�Mr+��NSl�8-����GqF|/����������8�{ӳ�Xd���kN�y��b�#��0ͮ����첬N��*�	`S�DL3+6uJC�-P�����
�7m��P+�f.G��f��PG6C��,닶�\|y�A�۫9�(��՝b�ò]�����I��e��_ ����ƌݮ�m�Z�}�a�a�m+j}ia���AY).qΖ7鵔��
��f�j��ʽ\I̧�S$���8�畮��G�[�%G�q9z�;u������.�*����/%%�W��pHhq=IoO ���]j�e4��P��+�����e���w���o�����e�,M�2�Z�T��{�_7�>wÔI��u����r�S��T�:+��f��mfWl{V%�C�L8�[��m��A:���a���tIf]uhz� W�l���6&�Wjb� �0 �t{�﷩�nٿ�M�KF�ud�\;۩J�T	e,\M���t�s�;P��@ҰXJ^	�ds����梩�X�� c�+�2��E�Z�z�v�uvs79���%��I,sC>:&IÏ׽}����;WuDFw;����@>2�˭l�1�<�w��:ޭc��{��8JF��L��L[��Ĕq�:kR������ges��v�������L��*��'}#��Ņ��PÁ��U�K�)Գ(��躍���ջ}�8TY�����YF�E��>X�9�B�ٺ��1�i���d&
R�b��N�e�y�C6�\8��]df&u4���s&a���˼Y�h���]f�8�4�c�Ҟ��@���!���-3���[�D��>b���[���B�q�Q�{�gRܥ�+hl/i.��c5��E�O*��p�;���K�]�Ć�h�'>y҆�Y&�]qGu��_jr�;饑��9���@��W\��G���P�:�X��wo����[h�GQ���򺮼L�ӥ���+�[�t~�Y�!F("�gD�&�SvV�u��x�÷ƕfE���`�']1ګdQg*��rQ�gf<���J�败lYjr���r�yPb#��g	WgJV�tW�E���z�[�(k��cȮbؾ:���AE{��НS{��lB�,J]8!�dR|Fv������]�n]^���-R����kZ�]d�if2E��Z��Q�:�P��nU�m�̹|���կ%��y�/�n��k9&����EV&� N���ܸ:�i�nO�7{^E� 4d�{�@��&(�쏛J}ǳ
ȥ�WJ8�钯E(*�=��`z.���LWZ�����JԑuD�>�X��0r܃���t�rb�+��}����s���K����*���3��ܡ��m	V����a�6A0��V]����Z��*�ʐj�d�l�o�Ѹ]5l��=����oE_kŝ��z#�p���H�Λ����{3u��P�N�#<ۮ}�ar�"i����*w�7���B��SDھ�˕S�dj��A�I%��U��D��KJ�:a>2��wr��eT]!9��%f�ik��Dt�K�K�y����E��du���5ww:DZ�t�r�R�*K���.{�������'��<����<�(��ݜ����J]t�̮Ef���#���*�#��?;���B��:IEQ��M���㨤!�VV�$�ADE^yx}܊��;��<���՜��g�u�\(�L��1tK���Ѝ���rD�=����"C��U}^I���*��'w"Qc�w?�7f���<ÝDT����>|�vh��^o�����vE���<���
�r"��_'����bw2(�;�.�乑AqrC�*�Z���9A^돉/�9W	��w�u"�{�r�VANHG�]�h�jRt#2�=�US�$�	E�^��)G!�<��غ7
|�O��ާ>�{���$�$�>>{�P�y�|�&GW��hp�DZ�ww��(�ZP}Uud~W���S┳�UETE�,��BT(S&�   ݅���ޭƕ�'�bLSe�{�
{���m��x�]7�����]�Ԯ[|zQ�!���-��w�ܠ*�HF���Y��9u*�;�ui���]�1���5�,��͆��Md��eT2e�>^�{�&:7XR���)O���ܬ*�O3`m����K�,�u���d���p�dg0��/�Wa1>���]��Q}>�)�y7�vM��X�����.׾�v-4f �@L�{;�b�j��{�?~��嫽n��ɚ�pI�uس:U^�v�Ɲ������q�s��FƝ�?.~��7��gE|C��~��ɗ�a�{ژd�$ȍ�0�4��9i!v�K=�7�����=sc3p�؞��A��gc�pȼVfC�mA~��ݓ4]��������� k`~�v�-��M~sL�{a�Hx���"�2���q}�u[�}*:�Ľ�_�I&��@�r���hW��j����/pomOx-
�P�:gj�;/��gj*lny�(3E�"F�y�V�;�+�u������s*�@Z���h��#1=B�`�Ɩ�차�%]�1!�bE�O>��Ԉ��ΰ�CS3u��Kv������7*�&�J�¼ո��ʷ��Ź1tc]X�n�|�]eUͨ�xA�����Lf�n^H�=��4׶�<������wA?[��Ur�����? U�;%\�O��w�N&jni����^��&�ӎ�I�Hk��fA���n֖�6|aW�.���b''���w���$���yT,ǧ�u ��-s�Hl���kL�,׍e�+���N�v��v�q��voh��sN�]3�9Mr ���w�h�)/&��3�9����Z{�̖��Ϳ�*���n�z��1�w�9N�������M����1F��G��zw9D��"�:�֌�ב�铮�䘇�����X-&3���dC���Ʀ7m)��LH�I�]���L���j.������t�܈����@�f��j�8�~F}��c���-��]zmh�y��4���#;s��*oV��4�O���OH��=���-��.�?m��\-;�O�S�Д��{{��ٵd�Xq��)�J��j��ͣ�7�Vz�3n=��c;�.c[�p�惵�-���{�=pӥC�l�H߷3�G!m2�8�%��I��n^��EC�)f�R��授��o@L�ݷ׺�7����IA���-�kC�]V%�E ��AL��Œ2��=Ҡ߻�f�\QU8�s�b�v`���P����:��[�-T�6�,����g�+1vx2�iye4���z��d�s
^�IyO�J���ӯ-5ܱ�Ct�S�u���ƨX���W���0�zi���3��]�sQ�u��cǢ�x�s5�����;��W�W��*Y�C�/K3Z��dG�~ ��h��QiLM���t�w�C��Fmiw�,�����C�j�ʼ���i{� ��K���.n���K/�nn'�n����j�H�p�a�k�����P޹�4�F,w�t���]ǃ��Z�*,������mG6;;��b��6N_"���*�ˬ*�/ݖz�-�N͝B�9�v/���B��/w��^*YYm��?B�n�r��M�U��5p���U��񣲮�)�훾Z�^��;���3�P䌱���y[�$����j|`�qUOe���ma7�1|��.���=B�p���@���ҹ �Ӣ�D8��0�n�|�9`y�ޛ�;Y������݋�B�
� ��S�QL�3#:�2*����W� TZru���׎hK����-1�xZ�z��l���ω�۴t�6��l���	|s���)��`�����Vk/9G�	3=�~0O��
�NVC���}�U�W���X�u��L��/No	��K�Ore�؅��:����s��˦;y�%��֐��V�2�SG\�R<LeY�3Gue��P������ᴰ[ْn�UR��}ٵgo����3&.3J�k(�j�5o�����qa�6����j�C�v�0�N:��y�G?V�;��d�gh����|ˋ2��<�d�M���K�Czb�gu]9����/Ԟ;�f�<�����oqH��ɷ?}=+a�˭��؅�<"s�}��մO��*~�*����9%��9���L�ݒ�8Y5���5[�l���u_'|v��w�Cv�s���$j,�c�G�S.�Þ
�{4�sT�]9ػ{5U{[��mҺ��Z����m���:��me�O��hpTA�y��OWX���|to��8�#dK�A�#�:��+! ��X��Κ���mӼ/9�Qs+���lWmDn�_oL�89Pf��4�w���=!�zO#1�:���j��IύS��fŃx�ԝܠ��]rD�Y7H�1:�ˮ����z��L�PʀP:']��Èaa�t�r)��(t4�F�����U��XJ8Rv��]~Y�j��Q-�S1���Z�1f�n��j��*Y^�-�E������&R�*Ww�S����N�nO,�[H�<�վc�I��'�x�0c�3\r]d_���R��ȵ�sv���wf�`����N����h�^ȯ3r�p���pu�/�vf��V ��D�/Ӧ38[=�y�N�����vϒW���a��ş-�c�ӷx�=l�U���9�Ԏ�a�\�?v��0�~�G� ��"�ݗ���}3z$�kf>W��L�W:���e���1
m�ɸ��%��A�"�̷+�{d�nף��rT�g`lgU�Fj�SLq��EesҨ�3R�ӷ�NE���Y�+� �1{.�{+���T1�]�H���iy;�X������*Fm�=�X��/�p@K�R��l�U�>������@�_G�#<�������DfwMĚ�L�Nb�N(̗XU'm�z����csu G��M����Qy�p�V� ⺲����ms�;��"�&����gl�j� =z�`s]o7�Vo,f��ӛ� �������Wܼ�h��ąe��-v�ohq�S���$�Ysa�L���^(��f��%ײ���8�Kp6�ܥc�j�۰�7��Btc��Na�Z�~�ۛ�]�\�~�m�K>����f�f�9S��KbR6!���oy�YϚUHnu�M��ܬ'���P�J�����Rdڄ��1�'.u��	=�&��5�I�*��T�G�q�_!ȋR�%�l���AS�e�������o*����4����ƖP����_)�خg��Z�M��^�����������'�UrR�y��X��Ms����D�{ybV�Ps�}��ǽJ�RM%+�U� �dѥ�n��������	>HMTm\���(ǈ�p�9��Ǵ7%��y[�
�f��Pi��+.���7�X�j�<hӍ�a�g�ASp�o���|�w�q��X�ܐ����O��S��A���Z�NΝ��լ���c��*V �Y���y�(hS�*]*�L_���}Ν��<+<^�3��owP7E�P�v%nY�9�D����C�3��a�eەx�ưv�E)�W�Bt�ܶ�,�=ф{�!LU�e��i�Jc�6CM�S�#�ٹB{�UC���Ƅ�ǆ�UC�I��H�����LK�5sQ=P�:�sj�mv?|
�t`P�p��\dDr53��M��VKa�Xrf]Z�g��%=�*zG��l���׿f���o��%1`e�-�Q��?e�ޠ�s8�Gd���_Y��:��= %A���0���b0�b'�Z�55�2����\�X��{�HJ�u��i�{�ϓ�<e>�O� ���>V���N�4 �z+�@�R���{t�'[���Ŭ@�W�V�Ɋ`{ C��~�Y�F�=�	����:y�r|��jOz��5���|�J걦2�sy���2a�:^��N�;,��V]��,<;�����јv^&I��;n��h�5b����3`�N�f��1U!�JˣSq<�	 �܀��ΐGv�Y�#�h����Εj��hM�p�����P+G�#m�୻�P��ұ7}�%���}�q��t�׉���������U��=��w��L�)�5��g�½ڳ=��V��ӧ�_R΋��u����G�X���,��ɠaVا@ϋ�9	�W]�5\%�μ�I�jggo��%�c�����$o�:WPYu�
��;aEX[*�a��l���<�j.����3������o���:Pn�'	>LN���J�(s�^WA��\o*�q�zv.��u�/5qt�[DP��ǒ �% ^N��+�,]�L�aoe�ynj_v7��GPcu!���]�$wHݕ6m�l�D�)�--0��eftC>�e��spI�PS�ݚwΑ�Dr�Y�O>yQ�l؇z��s~��R��r�;�I�a,�,c-�ޘ��)=&tq��l������r��l��޵�f��+�B���L�ilS~�4��4ܷl��7L�Ɉ�jd��ʁ'�E��sV���+!W��}/�?�sn������:C�λ�xX�����2�V'\s�v��bu���~��ݛ]�_\��t'�H�4��G|��Ƃ^clϠ,;��ݫ�'[�Yc��8�F�~_�_f;�2+�:T��*Tw�]Y���\t�̽���{a�u�ʲ��b����P��1q<�[�B+ne�Z�e\�y�cl��I��}[R�I9�ԱwL��ib���1�2�=���m��-�\5Z0�]�7&�MbV��s�V@l��h�����g��\����Օz7�ٻ��bqv\im����Y���=�;�b8�iF�OCj�<d�_�y���L�OҜ�ϖ��{T��)�n��/"�JC4"�o����S��e�R�A֞]No:��yɞ��F�o+�Ld�~@�Kd*��6�r��KY���p&�͍X;1Gt�.���J���uzJjԝ�6��̠�Z�#��|ڈ�ws����pWezl�Mᜍ�6�r����i�����aOs]����v�խ�5�ƼD5��*�R�k�-�]�%��*bLC�=E��������ܐZ���Spu�tվ��=G����l��[��A���y���~�+"�����G	�K���&���:z�����P�8��A���D<�2��]���Xc���[�{r}�[��f�3XII���m^̫��L�g&�u��Ҕc�It��K(�SuQy��0L��@�v�k�PT�^��@b��'��U֮�W��&q�P�B�Z�]i�C5�5j��B^G\���\������ԑZ�
�G�]u��B�+�srvȱ�2����nzccm*�tg�Z�|V�����6�e<n�e�cكw�f�5�A�y�̉w԰L�{cz�wB]�y�$�3���#QU!�eּ��N���מ��p-���"�@v��y<������i�h�q�".mG2�ͳ�:M9���1�"7���ZF�fwe�/'*!�M��F�Q����[�8'��H��`^��
nwU�'wjܰkXs/��[J���!n������b-c���)�lR�����������On�t��e�,�L��E�S���ݥ�"�e�U�G*t�u
��f�{ޜhe�ᓜ��2;*�^�s�k;R���	�$2J�wW����E�Kt/�^_f U��-{/N#2�R��W)ꑺ������0^�����O�4�Hh�;�D�d�x�P�j�Sj��ҟ�*k�	��}� �<�}���>?�^=,o.�A��r"�KN
a< ��	�G3x��{,��GI��K���t�\Vn@�)���{����G*����&G�]�v�n�ef�cV!��;k	':d'��v��M�bn�Zr˩t���Z�p���lZ.e�xL�As�64ҩO�@�vͻO�0�T��Ma���6%�T�;�Z=��-dT��Ub[���њMW
w����5��} cpq���k{����v1˥�YS�p*���jU���X=f%c�Ï���Q-�J�/i&u�G�6�Z�(��#%O�R�]t��mG�u���k%��J���f�庫���)����w���P����#NC[6��^����ޮ\Q7S� q���(gjilu�
}�K�R���PDmd��sk�q�2�^ˣ軑<ę[�V���z��] �V<���Ï�G8�6�؝��I�Y�W8�52��:���@J��EjUաKj6Ow,������J
Zcz�X&�[26��o,=+{�T�1e��ɪ���	Y(KՊ��D�`O#��v�֬Z���M.0���&�7�#y�FK#�f)���ب�+����}ʄ\95�ۼ�,[ޝ����צ�ŉ�N^���U�9�Ũ�̃���]`� |F�;,�`�+f��f�	Δ��W�(��M�Sj�1�J(Gx��qU� ����݊�s�ַ6⋞��+s&;-F�<ÎwR���)�� ������V��z��u�����TՖטg�Ӂ��H��7��Rz&:WQq�fF�s�MY����T�:���<g����\�6p�X	��ԋN[;�.�:��v�L��(�zi��qt�e�SQcT�ν��L73�M8	*��}��1v�q侎w[�n�HZK�h�ct9؜K<ep�b�դ�Z|K�]��n[�eAx�=���
�2�(y��b�n�����]ք����9'e�`.Jͽ��#"����:�u�����qtVE|�Q���.Y����إ/�`h@m;)#CP�?�;�A�٢��t�S�v0/3jf�QNLd�:F�fٽf���;��X-�/���"O%N�\�v�n.�f�"�Ǉh;N��؋nĲ��Ц6���s	.%yc:�&��N��_1t[jJ�p�馕�ʴ-&�f%�Pncz������h1s6'��
�\���k0Yͽ��������6d'��#_ΧQ;��"�V�toX���T���5� E�Wmv��r�&LW��L�sv�}Ɉ���"�k��X`���m�Y��[�2�j��0$�����6�ͼ�<V��I}����鸪��Pٔ/eը���I�+��o�����k���5��� Z�<ÝAN��VͲ���T������0�ݕ8�ٺ�7i�xU��u����Pِ) Ud���pR��n;k��+qB�����|��'Y�W��鹌�8++��(@\9/�9L��PI�TU8�W��]��sR�
�!<�q��,�|}�wD�Tr�EO�9�R!�;�Tp��R�ιv`��dr� �wnxW� �~'�Ep�b�$ڴ�:�R����~z��Τ��U(���%��9�̝���/��s�P�}�8��A7�Q���y�\K#
";���P-I�2���y���j�;�EK��$7�8]á&���t�y�w#�p��ˏ���y�N�ruf��%]�n�Q5j�s��N��'�(��E/�o�#��Qp����CǾ{��9�\�.y	Q� ��/�G�UϺJ<����Ql���
���TBDD^���χ
�Ӈ�)Ⱥ3�ܿ�B�^H�|xDy��;����M�=y�صc�� ��*��'�R�k(��;��"�K����$p��F��ŪO��x�z!���>���r/�n�N�y���'J/�a=C�ޤ�$�"���<�0�9Y}��
��=0��Ŝ!�;��u�P�E]�W0�;4{ϒ�Sb�����<���.��%�<hZ��u���(�]C0s�I-p ]L��Aέ�z��WF�5�����:�c6k4i
�w{���ug����vJ���K �e�״�[��Ɉ��zl��Ɨ���{�â��w�r&X�8��74}F��G$����/fu��#!Z��ܸ���BL��"�ek;f%��%^Fe{����ܳ���*F<�l�Ó���>�~�2T��h�ʇB�@�EX��N��7�@�a5B�M�^'�]�; �8��=0����Sð��4�k�b�zwF�D,aU�}�ƛe�h�VD�X�0�>e���7���{��|ݗ��E�_�s�i0���ח$ƽk��+��-�}�ހ���~�X��I���������z����_�I�5�O+8��
:|�z���(5ۋ0k�&�an�n��SC�&F�$�r0�:��4qԩM)/A�0�;3Ou�@��ʣ|cg�!�<z-��X�wݤ��Ş�{ҍw��(O*�/�l�m�W4 ����,�AGc�|7:3l^IOuю�X뱱JT��c\5D[�xf0�G��������]��}��e>�t�G;e��^n�>�6D�l���r��E�݀o���!Wn��2�X�d�k�d ���rI,<���ް�Z���fG�o��63wK�qn�
AE]�����i⮷Qʨ}����ٔ���T��k�eLMu�e-����D͆���/�l���G�MG~����xj�h�O̇9���{4����U��U��Ԋ7���7v�+m:
4��z�U^Ŏ���r�/nH���LV��:2j�8�n�h�9�$E�Zr�MWU�9��n�"�:��K�M*X2������;�H��tׅ�I�tn�����H�V�n,��w5�۽�g5�Nq�~�ؗ�e"�?ɂ�}dm�k|��3�>�'����ϖ��ټkx�@��K�᭞�ɧ�p�qZ�R�D�w��З&li�R�����Y�3ѻ���	���C��8��]�Wgś6��$�bMJ�<���{�����%��b���0Ð����h:��u��4	�7ӱ��Ԯ��v��X���4n�����Zp��=�
��Z�7�i��50U��J��6i=��5�GSb�x-.���dk��#5�����u{Bf(*-�(��ސ�Ma��\�����6��N9�c�+tN<�.9�Z�u���)�C�z�'J�]��/~��)D�R�1�ug�N�M�F�y�40�߮�eP�ӏ9�7�XA0�P�Dt ���rŷ�_U�PL�p��[+�Ղ�a�[��>X��/�TꟋ�r�>���Gx� ��=�0�!�i��;M�o;3�i��>��g�Ƃe����~^T����ϡ��kU�!Y�Ik�?���ڨ-�2�A�5��dE�а�YSX.tJ�	���&��b�W��{��'j�����
\c�O�;�ι[��<,�yg?p�=P��^�}&Svn�K�zlrC��\T�zY_�[�gj��\�m�p��wlŃ�-9gж�{no�*g���JZUE��mYL�:��"Y�鞽n-�BFq�7fFԅ�)�m�
 �h�[�9��,t"���jz�h8��f���
ιM|,�R�A�8�2��5Ga-�nf�z���٬E �(x���+<��
�~��%mc��E���R�3[�U��&G�����!����(%�C)�PՍܚ��ܨq���Iw7n�q0���g8�p�y��;��n-}��ls���q�&b9����wSr�R�����Z5��;�?mn�_M�6�}/T���j~Kw�8?��3�ë��
�Y�����Glv��V]�M��ު��qʐϐ����+�Df0U��E�F��7ͥRf�NѼ��7.%��+p�%}P��n����2q�73��yW���މ��
�h�O}Wpf����+Ik�C�.IV�^<�ٽV�}�~S��7�b��Wt��s��Ll�26�EqN��6�Qs۷M�z�c��
�p�fr�9��HzB�1�,��'>�)�Uz����uO`�I�/�Q��\��nc�<�g�d%y(��}x�v�4O�E��\�vcz����6+6�f�v읎�ګW�6A��=a�|}�[�2�F#0�u�2��n_�m�m��Sp}����I ؚIHQ*[�2��ΐc�L���V�?c���=������0a���>Gg��M�=�\O�2��.���[�+x;�/T�ri��iZ{�6���Vs6)��γ��c�����qYѳl�
���tG���N��-Ƌ���wV�./CEŹ�wXg��ٛ1&PFkq�����������4��P��|@{c(��!�M�ý}F>K#{��F��/zn�$�.�����]���l�̃�����;�J�q�ئ���i�˾�� x�J��v'(�^n�To؇l��q˘�Z�q��Mgt�4V�oHP۴N��X7)���S�D���]l�Sk���{��c8rIOmqYX�q�]*�t�=buŗǔ:kv˴�ŋ6��i���Nՙ;^8�hy@%m�/D�y,��k,�l���}�M���6C���S�#Lc<����YW"�-��y;���ĪYv�\���f���-��Al����Cu.�7$��<����_��f�y@_�R5Kyy�7�b�L�$3���#LT(����g��q�)b�腇M�8�ȫ��dfL�ve�&����ݽ"���lm�5�LV�g�ۍ/}X�nDM�찙���	$��'��.6�"��y�f�����������шKє�nP��B�wGv�.�:�;Ɋ,�IB���Z��i�X1l�5�� #���p�[V)%W����w+Ҿ)�|f�,���N�h�T��A;J���3&�ݩ�)k��D��aEӟ�f���*��Ls�٬4�c��U�!���\�}Kv�}>�-�G{y�H�+��M�d0���c5�~�j����X'��s���T�}��Z���KLI�,� ��#�^�����C��84gm�����|��GX�V���SioY�u�o��u����eŻbx�j����nb4;� �����쎝.��xt��	��U���d>�kO B��|�ۣ`�/�Ź��v��ju"�N������;��l���9�M��i���R"k��9�Q�tl�ֱ�,͵�E]n�׬z���H�<��d`a�i�B5�Q���ӵ�������c㴧���a@�����MװڬV��-	��=5*՘b_*�tf4�A��=Fa�S�
�iKjԕAe䂪��diqM��\�K�gO`�����#u����c�d�!�֚���F��Dߖ�?���+�Ѫ='���Xб�N� :+A�";K����s�����f�8}ET��=I��ƓO��x'�%Zz�vV�dg�sb��6��mάWp@�J��R�T�9`;����n�RoxD)`5�1ݽsnb�&wN�v�N�ԏ+�c��:�^�n֙��{����,8j��*���]�����̀�͓�Kl���qj�ҍP�/ݖ�6�]-�Y4t��g6��Ď��znK_��F��\c�0@4iV��n�ٌ�������e�p˺�ZE���u�W�7O9�w5��fT^�!��������WqE?l5���]�f���/�֙���1�O���%��M�I�J�2�՗�ΡB/P���zVE�.ɵ�(u��WW�֚<�z@�͑cϕ��8��+�搘t䳇��y�b�z�*�%�q�ŭ��8BAť핱P��!���Ci���T�^����o`��v�>J���n|\��?�p�fDf}�3�v��������M�:�ˍh�^��#�`�U)h4{]����"�Ŕvð�.��9,n[��.I#��B����U�!e��שĶ�7p!�A0�'��շ>�]>�gΟۛqZ��Ѣ�G]|�����SՆŇ�DK��� [��X�b�=|��]�-��c�\x]��ӞE�w7��\U�v��a���Y����E����9�fud��[���6�Eix��d޽��2	|q>��H��2��(*�%A�:��׹�%��fi�˺0�fK��D����c3G�PP��n9�mD䋝���h~kn}̍��oܢ=\�y�(�y+��M'�v�oĐ��<���\l���'���"�r�A)�o��d�{Ԡ�U�3�m���3m��aIm��}v����UJ�BET:}r���R/*�N>���Ӣ���C���u���.�s���&�V���>�eZ����@:�@��ob��Ă�޻�����c�*�u����.r ޮy�Գ�9M�WN̵�齱;�l��[p��k���;�4�b���W� ��j&]�T-�Vz��T��@#N2��|�@ا02���P�	\�,�=o� �o�N?a1�w��3X��*���rȃ�S��Uk�G��u^+�Ӥ�7C�æ{^e�� �TD����D��3<���GIj��l�3���tH6�1y�p}���y7�v��� 
��3�U���`�5%��{�����ә+
;y��na�]DwD��j*e=7,�q�IQ)��D�f7�*��X)�"�0���A�˔��8Ҝef\؆VV�����`rie���-���ws����	�-�</|v�4K]��W*���n�S�ǉ�~ӄ���i>�WO��t�3�L[sC��c��s�6�*~�lqw-%���l�ѮG�&�&{O?j%>��Q�'�C�����c�wJ�iӳ.o������5(�z4���q�}�I��
�ä*��R#h==����ٙ�`��G�1�]x�7��n켎��ADd�e�%�i]��ۦ;�7WŨ�T��4�#Fk>KR���"&�DV�I�i@��"�.��5j����s� ��>��^�c��� �s�:��5߲|��X���koI�F���}d�7ܯئ���ª3֬����v.5�Z�3L�@�5ߦ�6�m��ޅ|�q��dݎ]�Fx��ZU\�	cE[-�{��sow�U�Q�gk>���>Un+��:ur'�Y@j;���Ud�E�\e�4pg�}\�/*�6b�L$���ˬ;��m^ p�:ê:�dS&jb�YN��B��[��B�zd���D�X����.C���0ɰ��x;u�o���l��<�+S�Rs�o%����w(U�]._P�ܵ"��\��Bz*I��������Q���;�Ww�G��䒲�wo�c�lo/{����Xc�Y��1=��ң�+���B]0Gl�(ؾ��m��[���7ID�n'M泑vVm ,�	7�]����g+a��S�RQ�`�PM�
��r��7fj�~���>2t�Ӽ�%��c3��e�"􈂍t	|��SİU���'���z�oA+qs�.����-�s��5�_�T)3��~�x�o띮c�|���-J���)��� �b���x�s��d�t{}�dRj2a&R�r�d���փ]0�^qղ2�J��L���r�p�t���7����4��|Y��!�}C?:ی���F_8Kn��،�u���f�N�_w�M[�Bj�托|��i��c����ڛh5�uf�|�tl�.}�
�eu�3����u�nքA82F�X�"����\�i��g���l�Y��}_����{���ű��6�lm�پ������������|q��g}����96�p`8��� rl 9> ` `!�&�|�!�o�}������m�r���m��m�s��g&6��m�s� s����M���6�9��g8�l�m��n�m���m��wcm����n�v�m���m����6�9��g; ��l��m��m���l�6�99  s���Cm��m�s���v0vv�Ő�l�6�9�m���l� 96�g8�l�6�96�g!���� �6�9��g&����3��ɶ6rc`���������>����_�c�`��� l �������~����X}�'�F�f?w���o������l�0��������w������������?��ccm�߆pcm�� �C�B�<[�������ك��1�����?_�?�{��}��}��o��1�x� ��[���`����` D�ȁ��`�`L�����1� ö� &6� �L`���a6���!�����V?���cl� \aL����o�������?����߈���+�1��6������O���1�����@?�������~X1����ۃ�1���~����lm�1����p~ܛ����k��n�m��6�`-�� �?`�n����_1������{6��?�����0cm�������~?�g�?h{� �a��~�q���?�>�cm��������cm���|�����6���G������?�� ���������lm�c�s��s�b� ������}oՏ��o�`1���������������/����,������)��a�z�EUl�0(���1$���ԕJt��6�R���B�[T�QU!�l�Cl�-�fi�$�&Ҳ��U"�P�J�J%d+f٥*�*!�P-`��$���-��6�&ʠƩ4��4ԍk&5Zf-����d���K##5S���V�!��XMkRm�5��ۺf�gb��$��[kZR�q�Q�m��l�Y�A-�6�m��ն56ͭ��ٙ��["Ld[0�#6�m���5�el-aL���-�YX[cf���ieZ�l�ٵ,�Xj-Y
ڭ�J�*�  2x��BCV�p����9�9]vw'ZV��;����3qwl ����Wm�N��XБDs�Uڀ��Gv���V­��M��3e#Y��l�M����  ������hP���#������űl{cCC��ޗ��CF�H����|=p�P�C��$-ב}wMUhhұ۫��j���r�)kmMl%����B�]֭��ֵ��wM5�S:��sik4ږ��ٱ�Y�V�   {�Ɣ4-���T�kes�vг����KZ�YmF�ҍXڶ�M)�F��:h
�l�jC��(���kl5�vS�S�`�iPͶ�R�i����lڼ   ǽ�AB���9���!��7:���ͻ���N��Rv���`;�'N�U��n*����6�k�P>�^׵p
�suil2V��e��U5X���V�   s�􄚆��P�v�:
u�v%��u��Rvt���W

�����T��]����@�v�aDɹr�#fͫb���   {����  5V���$vv�Q���@tL]�D�trj��������.N�EU���V��Z-wn-e�j�l���  	�P*��oEq@�ˢDR���V�R��(\�r���u˨��L]V�t4�v�[��<���K���K"D�-*V-�ū��  ����!}�����h%W�{�^��G��ozI"%G�)�$�n�ۀ�]�J.:��*{�a�T�*	���AkH�r��)�%+��ު�MY����Ԫ-�5��   �__j��Wq8�m�_wy���[�׳�UI"��׺�mU�)-�ꐧ����J��=��^��R�e9�=J"��On�x�$I��m���YI�2kV���B��   ��̌Iw>]ꄨT�uyޞ�lb�����z�nz���h�OLx�҅[e&׽w�Z*@�ާ9=m�b-��z.����T�D| ��T�(0� )�IIJ�  "���*����db0)� ���hL���2�T @�J�©@ 5?��������������r���2D�輥�͙�>��L���A�o��f}�gٶ�����6m��6���i�`�����o�0l�&��6?|����3����ṞB���(�p�e;tD�v2��Џk�� \ZXF�j[p��Va�!�b���ɭH�8f�I�ܷbm���M���p@͢dV�e �V�ŏ*��l��c`�D�$��N�f(i�oB7i�m��̬6����ǒ���ý5�#%���vVZ ��3Lk�g��
�o����[���Fm�4v�єM<[B�:^"�h$�����������4���LkmQ��X��(8]+8�XK{�d7��Pd�N:4�ۻLQ(����Ss� 9�;(ґ�H%����#�z�g$�B�2�F+�KL��\:f����qEy �}`�Q�xt��,�]ń���I���j�7v���� ZM�9�S���P_Pj���(�i��v��:�Y���$&���� ���q#���ss{;ڃ���"��Z��,[��hF�:��9;̌�g4��<����up�2]]�Y{cv�"�7,�ʍ�y��M�Ѝ��mɏt�@k�Y$VQ,�0cW>Vi����t�e�;�҉=!�s;�Y�7v�|��<!���y7;K�ؚ)�g/U�h�z��M�ݩOÔm8MR��4K�,E�uYE��,F3����Lُ�r�@m��	39<�q�Z����rk$�����U����[���K�"��؃�����tʗ�s�t�$�́.ɣ��t�wVR�u)rV�ݭڛ���P����:�Ub��+3 ���$��HT�K]���i�yCsu7�\�93Q*�B���/I�	(k*Ky���@ۆÔ�����H�9z�<x��gj1��j��4<eƢ��Z�Yb�,7-��#E���x�-Ր��,م�%�^�Y*��ُ4��A�,1qM��6�	,��z6��6(1��Q����ob|�K�D�ʾ�]h��ZW`$�*Z�n��� BZ�15��S�,�j�̽r��g&n� 1��n�TNT�xU�p!�Q�Yuq�En6���TO�dK`���Z	a)CMݚM��K5���1�m�JB�H»��N��7t6V64V��,ԄS0kźր��1n�D����e(ػ�S;���И�f� �!*���dL�;�8|�g,����GP�g
��"���(��^�wXa�[ئ��Y��	*�?��Ŀ�'m�;&�d��l;�<TK97�譎c�=���j�:�kJ�O[��e#��͵�2�`�n��;t�z�@)��Z��K��Soe��'Zzr����٠Ƴ���0,uqʄ����r���g�`.�+w�I�m��N8Z��I�cAB��W.��X9R�Bj�����`��Eӎ��U�L�p;t�V����԰,�n:���Ht(�L�(�;wd:u��<9vW�̭��4aB�j�4ta`c�f���3Q��e]�v�gǖ�E֨S��K�w6a��Ա�,t�C�,WOml� 욺�4�Sn�+v����MBK���.��۰�#)U�4��u�yм�*Ч�����C��]�Y��K��VU=�d&м���� ���w	��VN�H-}�9}��=�8�q{��7u>ߓr'�����t�]7��jѦ�:����+-Vt�X�%�9��F� ��/L��L<�I��+�Jb�������B��j��M&Qm��Z	���{�1.\t5�{�h�הc�[f����ݼՋuE �V�7]�R�.}�j��;q�C
��"`�麒�Ñ�i�Uf/����b��أ6Q�^�l��e,�0�x)	R�&���H�M
ڕ�Q9�m�DE���Ҵ�>ږ�yB�ˣ-�^#��R�ٶ��Hm ��O1<U7\�l^6��n�+n���1"�P�l:R���R�1ۥ!ymպ-��0��v2a�z��l��X�3�k�uk�SIt�-���X�����\���wX�^��;3]��q�[I��wv�ۘڼ:I`.;֥V$R�7�Muw�����Au6y`�a8wj��!�Ț���b�b��sJ@:�{Y�3Eiaװ$Ah1&��,��	��n��P͡0��[B-��;����Kљl[� cX��V�UǏ-W0����62�x�u���JЎ&���d�н�-l��1���9�壻25t��ytٻT�U��k��SƤ�+v�t(}�Y�*MI|��B��ڔ�s3G���i�ަ�gl�h��:��My�1ɍ�7:8�F���8��&�d��M��m-c帮�7&�X��/o 2���*r5&hQ蔕FN��x/���a�+$�:rMѬLs���|{.z%�,�*%[e3�5���0��jP�@��KVb�2�+����� �/V�C�XK�db1�]b;���LgU�r:w��ñ@e�(��y-��Wu	h�F�^CL-O3楋)h[d�W����Wۇ��ǟ]�޽T��ɸQ��T�%uĖ��JMԢ�σ��n�Z0i��P����W6�4�֣Zm[�Tn��c&�l��qfAnJ-J�Nm���@�N�Z����"t�s�U�����d�r���Cߐ��:E�Em��뽺z�)��0��k-����^��2��iU���kyt"/F%1���AlS��l��yeP�5�$2eօP^��u��۬���ܴ��j�7�CxPO43d.����i�3�CӖ��S��z��wP�g-[��ܖ&-����6�<�(�*�%�Jʫ�$
p&�����[��:hwNBEnP$��oD��2��
��Mf�(�vز�[2�L�ֳ��ֶ?�E7\�VK�xYY#m^|��C��f�����4õ��0�:ƙq'�ܢEm�-�@
q���VQ�� N�Zb��zah9FL���5��´v�q�
���t����n4Ɯ�����ؒ�ٚ��8ҹ���׷���cq"B�ah����;ѩ���0H0�/І�M	��)����p�u����Zvʤm�n�8P�c,d��T�쳻��[���n�#[�+iYfN�'��ñ�ڽ�%�A�-�m��0�ҁȄ�
�c{"I�3*�C.��&�+�.5�at��ӊcd�Lp�Jn
��7���$P��Ԙ�{�'�C3]M�ُt�K3�9��G'lTP���V�Pc��#F�n���e�Ge������:��͍��m��ӳ`���}��l��޷��m@.c�Pn�pf=2m7�1-��pm)4�Wa��(f�8�w^���� ;�([y����{�Q������[dn`�d�2�0��e0�b�4Z��h���������tq#X�p�Xv$
���� �Ac1�2 ��-��Y���K�ƤX�ϯ��L�因�� ��f�gP�@rfѽŲ�U���.�B0^Q�d�հ� �8Y��^AY,3D�(��-2.��ذ�L�Ô���[-�4$t��P�
˨�f�P���RT��pJ&���VK��e��Ou^ſ^D��D��1��kRv4�f}�ܝ�>[�@�|�E	�*j����P�l�˸cv#:��ܟ5-�.���l��V���Ҡ^�	F,��A�����,�>2YU3i�x$Ǖdѷ� �)�x����LKKy�9(q��#�إ&Y6v�r��zcYed�p��kP�ɷH�h!��ح��i�T�<{�a�gc�z�z5�d���@7��'Ak����9R��4�m���i��TE^�I�@hח�/V�k�f��婙�:��P�VD��+FV��gqX���Q�w���قa f�^兂���E�F^�)鴉z[��>Z&���Z�ĕ�9o4�������,s(��9PK�A,t3(��b(U��華7��9�TGnҸ��ţ�7*챱G�P7����<Yj��Y�R&�E��m�諰������H�1x�ݵ#�U�]�j��E���m�
n�{���L*���B��h,�I#B��=)I��E�ս���w7�@Z�f�.��H��f��֣CX��M�++T�k�Z����v�hܠ�4�V�:F-U�X�~941�Vh����ґ2�^�ݗ2¨P ��z��J�:����"�o6���9O��F��%]fޖV얥d�6�ux����)�*9�먋��*B�^���n���P�\W���$�ʺ�͹j��Y��h٧���̡�U�]3X�"D#�v��i�Z��\��P�ZA�!�D�sk.GB���lb��^kI�S��,�fnR�oh��%��G�d8���t-�x��D�*�LF�P	��IN�e��ua.�����$�n�q�Vv]J��$bly2�6eҊ�*�/�z"9�dxV(�-9;�݇���T�6��Jc
�ܺ{j��UfIz_��H��&�LI��ײb#�pÞ��F�9%�6�̻w�쭡��r��M��z�G��g���jt��/cw7s`��tN���ҵ[���ς�1��+3^h8�)���n���&K�)�0P���{Yt.�wA`n�{�F��=ٺ�F���G32S��x��12��"ӫV�ɎD�j�XP�j�VRm8.KiT��v��5�%JV����Sx7[z�H,(��
u�{���I��nj�wr�Y)�wX��I��a�h��hU�1�Gsr����AԾ��о"�
����X&��&鵙�:x���&��8諱u�M��|�Q;,{u3)�F BH)�h��`�`Z�-c�e �7LF(q������t���)f*j�Y2 �|6+K�i����z����r�u��31k����9Q���d��p�R�Ĳ���I���f��e�-Q�X�2�W� �>uH����t^h��U�ܵ���:ԬD&i�,�7w�ൗJ��j�wSR�x���*��eZ@��_n�����9V ��
���fTN��$���G7bYT�ֽT�ͲR_Xl}
���#�X1T�-7��0kcD�ֺ8%ܒ�c�[���=���*�=�hRJ����rn�q[ [ j�M[�1�a�@���L9,-Ԗ��Ϯ�P:�:)`��/�j���Bnm�i-z�u��j&����#�D���Vi'y��m���4c̘�������Jo�k
NSI�q{vS�U>�B�U�L�DVވO�UŃ7�U�cI-������w��[����a4�fhݺ�3�AefĠ��)վλT%��Cw�Of��P<xEǡ��Yu��%�I[�[(�*��#���`�V2��z��c��<l�E��ʱ��c�l��K�U���v�+���������ۗ�̖��:�0�����%�a峵b!�����³J';��T�ASج���f�6��aV:�m,={�p��Z¬HGr�Q�B�cZ�D��q���A��L�Z�`��mcл�'�n�4�-9=��1���ڵԫ>mdO56��w&C!����q5B��i�m &Q��#�e=5xwdҞP8)�W ��Ц�qa�x/(�G5����=�}x���z�%��� W�l�uy���Xt��D���B�3C+^�&��2*�jnIt4TYKj�sRr��Q�����vFc��z�-�� ��ne6u���dn��G��Ke�mKB���743z��v���P�ʭ�XXց�XD�]j6�(�
�Ä�t�)�Һm}8��X2�5��i�r����Ub˽����Ud�2�:��A��1r� �"����;J�-|��a�q��ώ��l8���uvӻݤ�n}+r�҂�5���K�캿�ת����F�CR7���A��>�BS[�0K���m]\��h=yPQ,�G�>�-6���6
�P��8��v���6���V�:&��������I�&�6;�jФ�+^�����a�˲PkC�vX�����M`�z�`Dk Sb��#j a��ٓN��ybj���V��.L�RWWR�	�Ȏ5����5��e!j*hI���m�ӋA�xj9S5�X]^���V��إZ��]�������bn�9��}0��,�kC��8��x61q0�iV�+��u���na��!�EBj�J�'\��#�Z�F
"R԰9Pdc��tc0��n���1��)���O�-���JB-�v�=̙zj�m�ٖmf�u�r���7���+H*�V�T�[{��M�1;�腢R�l��m����������2U���_
s1�i-Q�bf�%DN-����6�6��f�1��\^Fl0�E�����RKy�kS��r �.��St��ՒL���n�"�g
�B��[��$�WJ�������!�a���س��J��)�:k"�>�Z�I=!$�˫ʈLߠ$�:iQ�Æ�<p;�)�K^6h�;;[glZ���Scph��� %Z.�Jއ���]��E;{p[�c����&,&�O�ۭ_e�vk@Qu�C�l���n$Nț��8wqc6(H�hH�W�E��,�l���ω��(���cՍ�p9Y���Zq蕒ݫuSp͛����0؀#}-��]ہ��H����#�e�ldȴ�!�Z�0�p6�4Rb���*\:)*d�0��艕O* �%fc���� U��lNc̲��+u��Gn�Bw�Ӥ�rm�4�2��efS�[-���&�TX�W���۰ێ��Ekx[�6�j�R���J�ZH�:��%�,�n����ͺ��ef6n�]1I�[�G�m�m�1���/.;4ԣ��5-���i) ßb�U���F��>o�+tб�7a�S��R�5#O(�C��@F9x݇�zm��d��A���G�3�����C���c�c���e��Z�����\�Ц//+qjGY虜�l��pB�738g��.��Ȉ�VzK���>/�v��U�"Kc�az�\�\�L�F�X���\���!����nU�%���k��G�)�M�*ޘf�_Z�ڨ]��(�L>�9\��]u���.���j��w���ݦ�^��n�ۣHЭ:@^G��$TF�.j![�>���;��ۑ�A��u'��6��G4]�XJ��]t��U��gI��o�c��,2+�,!�ϟ+��}��Y���(\y	�� o=��vOv�u�]ܚ@m]f���-?\Cui���
�]M�k������u�Z�s8�'�V%"g���:{��|w��.7f疠g���Ї_iG}���z\.{�wjd8�h���sq�@՝YN*�:�	���1������e��}�l��k�%&4).�7�[!7�*����gt��&�f=�g]� �7S-���q/�%Ý;<���o���Q��nk�a")Yd_T�S��O�.b���X6�}���z]��.����`�`��b�/Nհ��6JPc�=f�ۤ
���������=����n��i&�%��\�/�/Mm^�')��p���ɭon��0���׈F�l�u	�Ğ�[���&L��zv��c��d�Mb���wi��D:���6S�б @h��]���3|���ݾ��z<N�q��Tx�Z۝���vm�J�v콫)[��w��ϾX'<���4Z[�g>����X$�x�gw!��!Ƀ��Z�8�m��[�́������&��bq��,vJ�D��Az^	ލLӏ��x�o4�>I���=Ѹ�^N�1V_l�ӑ�t��,�A��k������e��Hg!=��ݱ���7aG�D %!�9.G��VE�T�Ii��լ��z�49x1�ݒo��SWh]���Z�dV�v-�i>�����p#t�&�Q�p�"�����d���~^��p�^���19�vط�f�O9��E�w^��W}7h�pN�'�F[��,���]��n���ٴ9o)����"��	Ȳ�7`%�Cp;�P��� ���o�p�m37%���A���V���:N����{�!���a:X%yȻ{a��j����d��S=۔��n�[DX�M��@F6�\�Y�*n�@��Yz�ޝ}�C9��a���̮:�c���` m��a��)|��#YfU����"����8ͼ��p+%-	DY�u������3c�k�,�f`[K.��]�Ǟ�E�h�LD���..򎭽rYf��z�`@�I������r�L��Ev�E���J�]�L���:�[b�Z
nw<�5I)g%Sh�v�z0Or��� ��Wn���L�Cl�Y�F��(��E��~B�������իh@����蚊�B�7U�\ȃr�h���-ط�-�x�㛛�t�p��>�Ӧ��W�x��|e1d$�q<�}��M:N�C+]󽬾�����Q˻�:,qn����5��)*�X8�̝՜�L�o%&W��x���i��BB�&c����/�%�*��ֶnl����T`Yt�#&��6�dͼIWv�u��ŸkRB��Xy��ܶ�4�Ap61l	�Έ)֐��W��f���0ӝ���5���cfh

G]�ͻ�Z%c���f�y�����;40~d^��&]�t�n۽�G��g��Q.���kq�Z9_K�͜ɲɧ&x�M�GI�Ql&���"�Z fz< �X�h,"�+��WSp�2�7A<o~� F�t�S���]'�Ʀ�9��ﭞ��3��!�N%eg,�9n�Fs�b'HV��Fr�>;70mor�Y����R�ln�[���i�U������4�{�We%�|���')�N�+M��3��g��������G����b�s@ ��_t.
'��mf%6���$h�x[Gj�v$ХcZ�Í	�b��;���u05d��-���q���^��<1͎�PS�7;=;D{��[*���<����q�]�F[��έ����ŉ�:[�2�������&�u�孔V$��1�N`�G��C�\��=6 ����[rB�?tZ�ۮ��fY��i۹��vYډöoiRV��q^�^�g��[b�e<L��y�^G7�{�%+j^nj7� '�fdŵ���{/�zm�L!5�vU��� W�z>�X���W�sE�����@��|^̝3J����������k>مVtٮtz\}l�f#D�*�e}����ZMl[��}ىE����;��̖��;j�EZ`=�;�4�c-�o����R�Jt���[�'���F�|o[E*���y���cFj��dyV�w��{�ZP`�%��&��H%it���]�q.�/p�:O9�1�gz�o�k������T4�����fXӉd���8�6=���0�q��͡��K�Q/q�V�J�Ч����5��52H��D}[�@D�ǯ��;�i�Tm/��i�I��	G`i���}��Ba��{�퓴1z��-���e�����v8�b�Z�kq쇮�ϩH�q�T��K���	A]��x�`�nf-���Q���I[�n��P�s�����:v{%B(v�⫢@���/e���4�h�yB�l�t���B�M��{4��R��xH*V��x�Cv%���{3�.ҳ1d��M�:�2]����	S�~�ǠQ�Xq����'A^��]�$��c�S��JҮ��y���u����W��u�I��}�)	yyS©Y���m<������iF'K�-�ط;��n�tӖ2����y-�sr
%�h���f�=��Ÿ�|6�]="�*�b�\0ЛEWG���z�b���, �?s�w�`��B��ĩܮ�u����zJj�:�Yݧ�Hm�/k�,ތ���rN@ϻ��XD�'�H�Ş��Z5���]s�h���d'�f���H�f���4�=2�rk��1��Eդ�zk`v��w+�ߟ�e���x�pA�����h��ixv5&�뻢3/Kz�N�Z, ��s ���w8�X[�s>����7�{5�)&6�$���4+cK�(���Y�/3�U�b|���hV&ܷ�����YLf�.;���w�cn1���=A�����X�:�2��x٣orM<��1���dm�զG=4��v��z��;��MQs\ce�۸�G]Y�S��5�| ª�R]��b�3r\�v�m�|��K�7���#�<��6h��]��r%f��^���tG3"��Ƒ��顼�6/z���[�huG�7w�����^җ[AB�;�*
��\$��fo�S���٪:���t����E�PC�f^���i�Λ��<����eK:A�n"�Ŵ��Gn���S�eٍ��M9�������]��L�n�ZƲ���U՚F�Rdͱ�,3����.�;�z��\����*����1#�;�se)��M�UF��<���`�.�8��.2�o�����}�6��v h,�M@���Y�lӐ��4��<�P��0fJ��PN��4Q�C*�<�!�NȦ�I�i�yu�\�l��q�-D�xZ�i��Mr����Ґ�a�s�.�Րy��E\P�2 ���cD[f�#��7v��v�T$0U�$����G��.������x�/���4ؘoi��
d6;;��R#z����|�K��G&�Ha]��Kj`on��Y�6��YSlΡR�L6pdY�9�Lgj�}���4U�Τz����;�Z�	�_,F�1Еq����(s9�W����,v��Q�a���ܖz�
��tU{{:�g}䁇ҽ�����g���uO���O%��繾`�Cc��Z��!ཤq<Y�*��O�ӳ�\��H�w�'5ϩ�`ٚ*�	s���p|��{4���=���W�Z1��^
Ƞ.�Ǣ�k&c�u���m-�8q1_q�clgJ��d�WX�߼oZ�k6����)�6��t�z�?�ʾ�у#[vɡ��峁�YL�ח �L�kkH��p��ث;:��S�6�47ٳyMu1S2K�@���I�ܔa��5�=�D*�/�f���U�=)�"�՞34:� �X�c,�}ܢ9���Sxˣ1[����nvG��.+u�
|qC/po��o���������x22\Nq8D�Ŝ&K���V���6�A�δʺ�:�=�bJ�c��.�N(���l��p;�L�E�O�;������o�g�ʵ¡�F���(�ì����` N�|�.KԔ�e���h�����鋳ud,�[U�K����&X��w5y�|6��>���Ny���[7���w��ջ��YrxδEֵ�T��O�o%^��xS���m�5���:�g=��f��z�ٳ�Z~4���N�����1�N�$oYp���0���&��rv6�K�hֶ{��cȗ�����o�n����D�]Z&����I1�to�n�$���������Î�®��+U��E��Z-�@�r�7Z���@`����I�N�9*"����+��ĲTh�é!G3h&�cY���^��&C�������%%��i�h*��m3��n���q/�I����{I�#��-ż&	����*�2������.W,<�5�Ϫ��d�;o��-*��Իg.!��	����q�tdBen.�pdT��繆\ C�4#8x	�\�R����逥���k��ڃ�D�,�C� 
�������8iz�j4�Xׯv��t�ڶ:��P*�v������Ve2��E]A��pQT�h̡w�\��O���J)��+4��o����^խ����4&�b};,H�V��yV^X�.��Fq��Э.�QÛ]����@+��]c�#>��rΤ�kP�\FJq�*�0 �g�� ,�b���p_n
�z`+K!���D�Fgb2��q���e���&N��ua)�w4���j�����d��ǀ�<�<�z\���#�fci�O�aǝ���uUӺ�v�`ӷS����E�������z����1�pbT%���;�C�6����ӊέiD�v�1I�p��Z}��%^���b����*��}��-fb-�sKHP�v8�{�t{ȼ���C3A�Z[���!��N�%@OB��J*²;�H���Uj��tx�q�m�R�����I��(���U8d]��d�Nm&�ڳK����ȝX��|�t�hK���{DgoL4)��t�VoEO9)D���G��Χ�sc8���Ò��`k�"oM�Y:�s��{����=&��Zz ;\>3�]�z[�0�n��a��ZA���-*���Vf�d�Z�����oA��E��M��d6�:s������Y��ڸ�r
�{�5t��u|����*Ch�����o���Oi�|�!�qy`��7�j��]�t:f��'�,KQ��8�nOM@l�t-�ۅ�[����=�N'C9�;x�[����tsD��_q=t���1	,�MF��j���"2ɊJ_hDl�	y�z���\�[�o�e���PH)Lp���;��KH��d��k
�:��m���}����v�y$�K��Q�q�hJK��bᔮ#p�݃V�B�HƒU�l��?!0>���m`+�v��w7=�O�/	���D������]��.��ûyFp���U�޵:�A�4�V���sJ�6���;*λ�{f��k:�5ց��8�(���1�j���qH����\����t9\R��nB$������@���౯My����
>ٻ�(�ɒ�ėcᏔ�Ի'P�i���Em�*�L�2����r�;'qX"��ܪ�:�1��2�1���Ev=��fo�d<ft�����	�-��/1��=ү�]N�j�ozM�W��%볕�1��>���H�X�+�ti��@�(ى��$p�[�k��T(IByU2 �Gh���zn��\A�C5��t�����*��h��Y�;�Qj'�{�0���ʔ_��Ǳ5����t���n���K�Խ�>>��t��(�������"�NKϯ���%�td�s��ܮ��kY�q�[�Op#ʁ��ϱx1�5�k��7���x���kS�zv�����乐�
"�7�4
<_>�U�����;ݚy�`T�Zw3S�{/�U�S���S:�.��o-�^��a�L���η-�(O)b -�w4g0����_eB��V��1[�OVqa��bӂ��s�js@�vx���}�4;�N�@�6��v�r�|h�m�G9�H��Y��z�8u�=w}�*ji�96�$v�aA՟H]�_Y<ʳ��6���}җ�F��[�O��WT�����0<���9�n��4��e����>�0��lSY�tE���6_5V�K��P���d�i�b�Mvy-��i�mj-M���p��,�Ӻ�f�D�Yy��'BE���Ͱ�^bv��P;��a�yz�/_s��4x�;��eK���@
��̀E
7��m�1�)��b��i��F�\��1�����v��]Zu*�{l���_�~獮`R��P�:��`�Z��rZ���L�_�gֲ�%-��).In���yv�#ۣk�5�+�:D1t�=��\�C�t����̚�������Dd7���~��v�l�V��Ѹ��ض�]�-��rՑJ>�e�I�;�+Z��츱�;�֨�F���,��tz&��u��vK��q��+x�L�R�(G;=����]~�|r��#H���8"��".J�a.WJ��A�@\U�q(R9���ǽ��}����|>��c�ۤ#.�U�]��!̇�P��|�޸)�L�C�UԒ�8�R�֐�8��atJ;�~�CNY�v�҂J�]�D	�������/eі;���:齷;/��7+M�n�fk#l�D6����ɱ�F
I���f�W��p�A�u����1#��/=K�/K�Ū7h��0��DN$��>�7+�6-����qvD�����Z��7	=kXgWxz�{ľ�Q|;�:��Q[�K���]�C}<���A�����W�RF����-�]�VgD���fǆdt��ux��;�F���du�L�[�\!���̭Ht�+�sc�Z���0M<I���Ed@a@�������HKM��Su�C�2�I"\�Q<��7���0l�)*�����`B��� M���8���&v��l����?m����G�K����ֵ��6'�.T/��_´u��ee��-wp�Ju�C�*H^��.qo!�ţ�]u����նo��l��4O*dĽ�w��EN>"�7޵
d�{�F���_�����P�lc��^�f=$�s�����d�#��B:�/k���+YPW�]h2�Րq�*e�' ��ru�Z�)�{�1���嗤�$����m]Hz�^�tg�����t����R�^~�g_���(�@�Yc�IZc��'.�d�3Wi��K�5���8R��D�q���j�r��#�ss3��N�	�^1l�c�����[ùN_��38=�˪��
��;3��'��|�v<�����ը�0M�{�}+�AJ]w�.BJ�Tv)�����K�}/�q���n]�'0ǣ���-K��@����V�}w�`tFQ|�w�rTYc4e'd>��"y�gf5�b�E��Y;��Ҳ�P�j��j�ۏz�|�Q����k��2p��nx }J[�ק�Dk4�y^��{� x9瓌��|�������ɼ�J��{[#��g�֦����օ�YH;�[�_.��ί���|X�`��3��F��r��v�K�6��6u��	X��v<Q��\&�4�y;�.Rg�r�|O���z�~ͷ������bQ����P��Li!�Lv=�
����)��4i�9Jǫ��y9�u�b���ƹ�흁,˻�\4�;�	�)۔�%K�(�*�;����t���l�n��e?�qFr�m�������{���78��}:{�f�����z�21�_6��r<Q����ǪK�G�*�����y�{�R�{�5��:-LY8�	�M�{kR`#�(M������1�yGyܤ>�|@Gv��Ҥ�&���yI�\;j3i7��Q�8:��:��%�VbFPN�Hأk���N7#v/v��#Mڦ�Rm�\,]U�)�;�]��,WZ���b�ï8c}���ᮄ���WG��{;�M5c�;@b':���b�J��ٳUՍ�ƶ�O���5��UԖ�;��jG�u0,�w��nN�S-+@��,��o���fԻ%3���i�eP|�^n�������$�v�N�j�L�.ʙB��3s���1:9�I� ���7:�W`�9ƀ�u�+��R͚Ge�0�_j�x N�P���:�
1z�J5�dkv��.�9{�^�|N��/�WM9��nO�ő�xn�W1]�;���6-|��^:Z��:/7"���O[�<�/�Y��)��ȃ;���y|���ے�eu�H�F�)d~�����^���;�S-�gcZ��d�nG����=T����`ڲq��̭������m����7�h�+��Y��d�^]l�N�֮쇹u��t��;���&ٕ���p�oW:�
��z�5�dh< ��ٟU�{�>�ΙYAf�lsY ehZ�w��VR��/#�w�������.�I�x�`�}0�:>��nٺ�sUF��X�
���x��L�
�������-h�'(1�⨦lWVsB�/��`�=aZ��Я�zfRNb��qPm.�]��I�+Uwb�F$���A#vs]��;8�	Z����c���H���ץ�8�ol���On��"+璬�خ-��"��6�v���i,a�>p��w4�i`�+�F�R����M����S�R5��V�D�=N�
�o�5���Z�Kx֜��������<^��m>􋽳�{�KF[Wm+K#Oq��MZ���o�mX�t.ш,vs�ͱ 4&����>��׸y�tY�
wk�۰���P.E�etF]]�R+��J��[�U�mA�z�2r��_'����m�	��۳�ab>��.���1(m�
SeT���f��[v2�GE9iJ}
��*E��R���Vk#�mV�D��I�U��u�އ9]��=E� �:v�{�¨,�Y�o���]o�8����xw2%�Dh�����V�Ǩ�E㜨�C�H��;���KPG���m�/���F<�)��_S؎v ��� ��Gn� ǻ�O�s�>@�0gok8��Pq/n�u Cu%C������ҍ�'�.���Ww�B���r�G�����k��2�a�5-��흔�rÚN^�Է`�o�%oV'��f��<�n�+ˎ����F��V;����q�t��7Z+A��
7u2����N�`����H ��+ѳSC�Fp�̲sU@�[�	����]�ӏ ���s�4"Ć#]S&<P�ΞSb�MK �'��W��z�0�S]P��@oNGӯ	d�C=�λo�����3�(����	�~�B���OήG���ɧ��9��z7��A��h���@�-rv��L{N�����G����P\!��gL���H��ښIR"?��hy1�7ݗ�i�5�U}��������3��x>���9p-���(�1���qc���9՗6S�)�F�L�-�M��D42MIՂ��\�:��A� u�)�`A�vzK�AK��J�y��Ly�����>`ӣĠr�A�9�uv�x�n[��p����kMERa��-hͺ��,�8v:Z�@�����hU�$Vg�ڌ�4K��6.�9V�����1��[���	��C0�Wn�̥�v<9/ZZ��bx�k +��B�<��{���Q�p }�eEn��-`�A����7}����7�o���5���x�K⥦ ?P�YM:��,b-#��v�����[]Ӷӷ-�i�w����C(�r���	�£O4�'9����[u[�t*�]�yQ��+]FIpn[tmT#z�m�7ٍs���W��/k:�K�ʖ���2!϶���Pշ���Ѭ�v��]�OE���u��B�|xF�|��n�x_����#�j�n��w�jjM$p�5�{U��5���q�,��� b{�5�w`n���ى���XOb��6m�v��Ѯh<+��^:ǓT�sp<�&p75F�䴂339� h��-�U�nIB�P5��٢��eE����0�.�EG�u�9�7iE驡�4w���&۽Cq?_��T��bK�v����9�c�M�w���ԱW4Դhݏ!�	 t�6v��G\�wJ���һs�5�8�We�G"�+ltnqQ,�ӭ`�Xǵv�;TV�x�	�.�"�)��N;d�6�g���-~çjZ%|i�f޺^��7��f �U����Ʃ��fTh�\��O�|e��O��f�aɊ�`�6� �$j�����=vIFT咞��!I&��&^a0[N��
�ل�S�q���o9�o��cMk�w_�6Fp��&2Z�`>��ፀ��"Ky\�e,�D���u<1���7i���%����N�mt���ءcw��r�ӆ���Y��))�L#6C�<��G)��6�I��"_;��9\�����츨Mϋ������OM�oD6��;G,�vq;KH���13���n}���t�[[�5&Rۜ��Nv�۰11���|\<.�]��;;E�ukp��<��pX'9쓭�Z|�=�|ׯ`�f��_:A�Y�7�"E��GpB��T����k��K�S��c]�r��#WݿM���X�'j�i|���N�'���=�՚�s�u?�\	s��dZ�D��&��`l|��.��*���Ռ�?m����R6x�aS%p�W$��\Ӏe+7#�p/����CtQ�x%gh�5��߰��BR��[�^�k9lKj�]^iHN!�R�#��eټ�M�]��.�&hd��%e�^ݢzte�gh9&慭���+�v��U�
���ܤ<�SR����G'5�q����ۥޯW{��'�%�����o:�7k��E}w� s��X��i(���h��F�ه(`Z䗻`��}Ǫ�|ރ���C5��ѽ�1/g�� �{�'�y��f�`�#<�no`�݋)�vM�6vjR�Hp�ƶ��'<��L���fD�B�^%1�Z�p�����jn�{3^��&s�nD�`)d�Ί+	#����H[dċ�{�k��u+��tu�}����<�GA������Y�}��p3��fYXW��gC�y1pX���9���p��<����}w8B{f��UmqF>Z\��%Π8c�0�yxd�����B�1�p��'�_�5�R�/{	�f�k6ĳ@�/�+Y���,ſp����j%q�f��@a�oC��L���,�զN]��6������n�tŗ<&o<���m��W��&�k�ľ�1#ׇ����1�ގ6b�y�8�ؘ�mޡ}'b�bMҥî�虭E�P���G!�Xͬk#ݳ�}8���
X�G:��йU��}޲��Xr�{M�ҵM��q.N���ܯ�'�cX%�^h��mMݺ�����s�^1xA=�z��S���he^�D�5���a �-��RI��-	���iI�X뫠�0�bHY8T��-��=���GE�#
ග�Ɯ���,�ŽJWX�q��v���*�k��P�.͋���.ZH4�V;i2_M9����=�s'�pN<����'.r�(����>��)�&n]�A.�h�֟�����p�"��J��Viv�]��"%�ۺX��]�1β���{aN��̐#��Q�����2��1�=vW�ͣ���n�CwR<�-���2Ϧ��p_B�;��zM��n56$q��/	�FB� ���,>B��5*���x�ǣ���6+t��wP��^���+W$�nWo=3��M�y\^^ZO|]IX�gA+stN��4C��%�X���6��\w9O�`�����)>�#�lE�]��({D{hp�;4����%�.���O��u�.{/g��$�!��o�Ѕ��ӷo�s�t���83y�znwW`m���+i���bk�k����.xP��%`�h��;U�gwq� �t���(.��/7@��כ��?v���s�t��K�����s�(K�@�
ް;%�՜ܙY�>�z{UHQ'r��S��o��q�B�/]��{]�M�T7K5sW�VyeD�[K<�]�'6q��ئ��pJxh"@����>��2��Yo��8�N����l�TEs9t�x�&�z������:ys�	�v��Q����P=���N��{���mt�`���W�8rs���˗�i�&�_I*���^��i�w<�yؼ<�;����R:9A��X0��`)IQ��*b��=�a� ܤ���;��H��������N�A�=:�>V��4ۻ�k�f���f�"��%�>�9IcCC�__U����fJ�Ð�|.wi)=�İ��F�N^<k��w����P.�<a��u��L��Ka��Sa�g*ȝ�n����Dӂ��ip�s�ZD:����i��ZoCd�wVsu1��Cx���k�MQ�9=k��]��n�8��;�h��f����bt���zm��<3}�݋�����M��1�m$3�'�*.�x��{���z��#΄�&���ޡ��{��to��1�'��rD��]�{,����'�]76����p�(��ܬ��lb$Ӯ����lLaX�I�S�] ģ�i�D�N9�s���ol�՘�0hn��0�Ťw��(�mq!oU�^��5k�sxI��CA��äf:+z���<�s\U75hpK�
���\Gn���mZv�XtX\g���h'ٜ��7�"�-����<�lcx�+�=��ڕ���l���r;�gB�LKG�Z7oM�i^�}×=ۻ_a��A��j�y'��c��UnVA�\����$�
��]�q՘�����lĝ�d�7��M]�g���*ܳZ����k�%��m=����>�K滚ǞS�k|3v�f56�*|9Xq�joFy���6�A��O� Z������=cq!��FA����{Os��t�-b�:���á�ɗ5ig��vչ��n+��\���\�^��8֭�1ŗ����D��]����ھLC+�A�Y�z޺�-�$�\�n�`������Y���f�.�C彩or�(�E��M	^�3p�ϲ�h4:�[&��z�e��nw���Z��75Lo@b��W�;��=�\���[s�Mz��T�Jyi�@�vn%�QP�8�wϑۺ�X�7pt$��踍.���hY�jh9Ù�ZҶs8I��*̮�%r��/��gX�֦�M�:Y5�n`�}$xX��n@ʻ�d���(q�y�&B�r���63���<�_K ��ɩ��Ax1Z":���z�
-�^F�<�N�P��f� V/r���Fz��}���)z6֣�����[�N���=6Z��/goX^!��#�X�њ`��:���]HκJ5VY�iH	`��ڃ������Ƭ��w���Ҿ��꯫�ﾛþ dĽ��t�eմF�c7�Ru�~<u�6u`U�7e<]��іn6_-�=�/l�H'�t�a�}����c}Α�Cn�9��y���W�0`�f����{�l*J�4D�xuT�+؛f-�ⶅ�p2� Q��U�/�4jұ�'
U����׌�%?V�	G{�7Dͣ9J��N{צ��ώ1{��&u�������c�����K8�Q� yb�ȎN��˷-gQ���N���f�$p�]�8	�*�\G�(�\������λ���B]�:����n����9��ٞh����7�A:��uf��Br�s�%��vueV�Ժ�p�ݣ/���rttk�}�^�U��n��w�p�٩�"���%����TK�|�.B�Z6r:;A���p�<+p��=�B��{�E��VT�/������5��7)f,��=<q��-���,cl����/�����)E�:�{1�3j|2�	:��{�ٴE�i���7�΋C<��#�co%��G�ť�an�Y0o%둌_����#C.]�9�wâ�x>.�xM�yM���mwf�`���lw���_ ��&w֔xs�<P5Oy�?+�j����`'�v�$�Q��iEj��:��'L�(��'��)�]f젆u��s�*m��� �8�- ��@��E���|�O�I[a�a�]�X�{�����{�y/^�(9��U�"*����<��Nk�����\�70�WR��tr�[��6!�aJ�йN`B�r����F'�a��E��Y;u�=�t�:�0[�䴕=�ұ2wB9�G*���ʽp(qE�L"�g��&�ywv���<'"AL:)�Br���t�"�$"�e�)��q�#6\��衋M�̽��F�TL@�U�'"�J�wC�r��<�C�L��(sK2�ZT�JF$J�QW�\4K��� �si;���a��a�
�*2�.�^�J3�g��w��H�]wp����sԉ6��g��$U^{�"��l�JLw;��^eeEW����U)PEb�I�fjm6D�3H�"�!,�(��GdD�dm�uC�s�B溗�.Q��R�A$���a�H�q�Y�U��ﻐV�\��z�A���2���u�ft��I�6�|�y���KI̽7k{f�Ʀ���|Q�q�)�{x�o�3�ݞ���C ������VsšU7��"���u�u�mW,����PƔ�� �4��Υ2̻����Cd���A�!��Gl[���WECs)�"����m�Z7�9	��0�( ��q���D����VI<=.��^�5�s��P��
Z��@���\:���A�}�����U�u����[בx�Q�+�(=��D�tU풠�D����xͼ��7�a�~*v�mG�E�{�b��:b��d`�
���WO����+�s�[n���Ei�r:��t�7$Z���N�m�z���n
�hT3���t������ʔ74�9��ϨdY�
���(�s��Z�l�3�δ@��{������e�>��Qg[�Utw��:�xkD�oˉ�H����,�۩�o0�y�v�lW]7x�A��S�n!9c��<w�	��ۊ���J�-�L�ʃppwA����cy¾@N���t�)��qQ&4R5�2�Tz�$���y�\9�E^���K�ڗ#/�R�P�ɑ������G,�r��N�W�F4*8y���)�'<����ٚ&�>w�����'�� Ko�&���3�����֗�KG�;V���؀�㹧�Cx��7(��)�uynک�i���4����U/a��-ѫ�=��q��pEb
v������~�h�8��n_�j���������7�w:4����z9Qi5Ӆ�1���-9���"'��h�|ڿ^��ӸX'�ݼ�3>OsCu��-Yi���&dn�Umʲpt��YQ�F��i��p����R�C���s 8LS�BA�H�tТ��9�O�i�q%�&{�J1=�7�$��l?S����AŻ~��_wF+�zvM�2��0P�p�ʝÙ�S=� �4\��q��z)*+V=����{8��l���d�f �-=���"��
��a�"M�9բ��ī�m���W�_�c)������n|�ܫ��tI���7�1���]���R̺��OC�Kva�ä�C	���4��b���E�U"*��<�6��b{w
�u2�1�K�ܻ������8��iey����Ep��Xb��q)9Xf��#.�q��\���~rBz��>�s����:q�,7���y1���)��޶ �NY7�Nk����橄�����Vy�cuZ��Z݊�m�!K;�j++N��=���l��ʎ��T�����W05}zX~�o�m' w��ϫv9�'���׳L/�r�n�{�f+���D�z�g٬+3�$7�*+���о���[��k|(^9��Rl�;�s�����zyY�{ֶ�<ߠb����1q>;�G����q��a�P� �L5��OJ����m{��U���01Pƺ�鎐���S\sPYd����y^ْ��Xz".��h�*�K�*Zq��N�ԭ��ڤ���� �W�㛶��L��ct�7��o���#��hʤ�GPv�V<��˭fgA���l����LH[�4��{����Ĭ�i�2<>4�T�ۮ���7.�Α����!�Mގ��!^�ڮD�yx�h���,`�a��n^�5<�T�ړC/5nE=����XَnC��&#Q� �����̬R����1¢�E1�&�G8�y�6Y��%���*�b�$��wJ����}a#��\^r�C�3� ͐��w�­{�N�:��vip���866-ڹ
f��s��(*��H�*_�:�h�b�����6��/��9���]n����(�C
u$�\N���R���=$ywY�!������7q"��T��C1�+��;!�+s X�2Y������x���ܭ�n���_֊�EAɻl��u�q
�$dZ��}p�;�Cp�
14`7��ڢ�eCbظ�X� �U�V���,R��]��B�[zh���՘�j�Fs�8۹�$;Uw7�w��Ov��@2��_�8��/Y��e3��ԋZ���F��S#r�x��ˡ=68 懕�1�`H��V�٠�{�y���N�nʷ�~s�"��;��	�CL_��W�T�g�f[=x�I���U�v,8&�>]'� ��A���ok�{�sj]O+�=�w�B��c2酈sl�Iq�Ǹ'uQ8����*�q/�������x�~�n���t��P"��b�Jq 6!�ee�1:�Q9��Cog��Q�~�Ɍ�ț|.Zb��[\��{f2���b�Lݑ�/i;����(n���X�,m�)�i�u�Q
"�bQG݀'�b�y4�3*2;\��b�b �<T��B�ѭ�p��G�V)}דy�c��L��t'����U�]g�ԙ�^V��FD]�봨nc�\;�����VZ��ԀK�%�tO���=5P�7^��(����p��M_�K����Sc�u;��hn��*�����\��Y*� �<����W�8w�q����l{�6p�V�ke�d���Z�4��Y�yN�仢W�Ʋ�ݖOo���)E0 �~�5�=N[�w��3���1�yGچ�6�f�y[����}ϲ��㻹Lد��̐+Cuҳ�5c'^(!z�r+]y�����:��9C.E����g 'Tc�z�9X�;�F�"\�0ܞ;�#����V���)_�������<�z�z�w6�����wx�Ȏp�3�}�i��J�����.�c>�9�8��`�Et3�>1���lL9����^ƯƠ������ȍ,���"aO .I���G���'�~���[����L����w���=�֮B��W����� Kxª�l��j;s�A�D!OiW2�V���R��=���j4Erb�\B}V�jݹ#��v�/�#I�`����\�Y	�'���n^QQn�Oq\[>�V�z
��@❂K�����8�'��ٶ��ļ����Ia�
�@��W���2�	��q�j9�}���V��,Q�w��_�����s��>��-�T>��� u�����h��j����K�ؖY����!���@f���%d�^NF�"�=��.9��9�*V�&�����W>]U0��g��c��t;ΦB���OiV��}���SX�w|����H��<$Vv:��L݋u�U�By�U�i-�A��Tz�xy,���0T�Au�]Ho�#��l���)��n��N[D�5����䣛1an�x�|�S[vE���~=�F]��x��%Lko,Э �Wl�O��ܗ���c�z��6�o�Cb�ź�7��@YN��:d�b��{����t�43��g#�}�^���叶����%��)�:<��O�5~>��HRbɒ���#w�fsy���V�W���;r{t�(`�C�ǳd	����Ro]¿FJÃ
8ַ��Ӵ�޸�_�.��XzXL�/rcC�i���]���(ʆ6V8�a��ݮy��ܗ�"�UHw���Gh��8�n_�V���6!ۅ���#%�$,K�e��砻��T㊭�DƎ&��+WQ��h�q���dq��w<�an�CjL����m���x��f�k��1�gk�2��1��,8Lpv���z\p�R�woi�ܴ]hX�F�!�"�3���fB,�v�(C�����V�Û2����%>뉴xnU� ]�K�N�y��zFu��@u�
~�B�K�#).)ѣ������n���dWQ�wm�){qK�t�o���k��T1p\�.NJ���C�*��
sȎ������%�
�q�%^�OC�ݚ\�K<�*���o�
��\&��&����o2
T�!����'d=��/@U��=x���j�k/D�e��ϻ�V8�qX\�YAa��΃��^����d��P]'r-�yKup��#@��h��z���tnu�C|���ۃ�,��B*.��x>Fb����~�k�{Kgo��\7>|n'VX T�5�(��Dhk�5��L�ݭ��4�.�����cd�acA�(;�ud��*a����W�*��ަ��[��Tj.Jgoӵ�\�W0��k�ra 5Z�d��x��v�c�4,�UI�q<�\H��/0o�]00Ng�a�q�>�(��<�	���)�%�˄Dh.tO_<�@lo��F˭3
�a��lӢxO�pG��4��p�<�^��;Q��zu�M9��]�ɸ�Q��:��˪��cv".̥�����U�ܜ�ڃv'��zj}�Abj�W��3�\��l����;���_�e6"�w�6�3���J��V�R;1�Lp�^���9[u�d�E~�-\6��݇���\c)���F�sB1�Dҡ/3S��H�Ň��fg@���,��*Ks"Zt��2��q/L\7,n�3�5�7�::��qmt�@,C(��1��U5�k0�)W��Xp{BV���P���Qw�L^i�+�ڳ���gUv6�Њĉ#��t��܄�:o��ǂ����tXw���P��l�"��vv̲�=�	��هWJa2���[D8J���O���4`��3�h�S���j���d��*��(
�'"_iq�ٗE�����0�Z.�/Do!�_/v�0:���BS+��n�D��O���	���\D*B�[9�B�\�����P����N�G5n'z�؄�%Dk�(���h���k���/D�M�T���)�����k w��*�Z'����W�>K��e#X5���^�7�0H�i �5ռ�rt�GK�B����§1nr�L�3�����Q;�i'0�R��ӵ��ǹ�{��	�;�"Kzme�G����kqh{rul��>�����Ev�g'k�R������@P��\���n�u�n�U��5�HC��L`����0��V�al>�<�-����۱ ջ���AD��7<&�������.��{]�IIC��9�#�}����C��{�:v�ު�QΨ���������2�e���b������*�r����yܯk����Ҩ��N��D���U����@��)^߮Z:��=R,�&�O5�b��PtE�t�7Us��X�}P�S��t�t�X�*�w	���@2GD�q^w��aޱ���5��ٔ�}V+i[�+�A4���Q�Awү6��n9� ��K���u[��b��afˬK]4ĭݘ�ސ�=��镫�ڭ^g��_`�l[�N�mdE)|L�a��<�NӸ^W�{����;�X�f�~����*����F3�M1 _��|c"��4�86rs�P��^�n�Ŭ��{�Zd�X%�"(F��&jQB��_V��\
�e�bv��s0N��4o&:�$3\�cuw����۬���|;��?���>U��=�Wx��>�n��r��]t�+␌k�k��>[�����+x�w>+ �(���]m8s���}���<�myf�H(�p�nk�Y�l�!�o�˦(����.�^˷3ۖ�\�fF�Λ���k�N�.x.1p�T�g���$�#�O3���(B������w=�q�̞R��Uk���Gz�t�1���\�p��W���5����ȍr4�4"/�Um�}�q9���q�JG��UH��:锌n#:�N�,lD�����<�H��l���wZ�$q��D:�´R'��H�炤�^37Uxw!1�691ZˌS��jlK��].e�st�<��� ;|�!2Dg����<�[�����{���Խ�Y�yG����1xr���2�����@hNo�����@u�74�=$�q@F���_o�ǹ�pӵ��8���K�<�5�u���k�+�r�iC�A���V(��U�z_�e5�	�;�����m%z��/�ݙ�wz�)M�y݅��W@%����P�K�A1ð����ÍH�����$/��;r��^��r�ݡz����W���x�w�jSX��gz�f�34�Pw��3��<.UN�on��yG���jJ�g���S�o`u6�� ~�5�vUԽ|
88��\�/U��ad�J�A�"AD�S�c�T���U`�������9��'t�!�K|�)�"��/�V��S
���x��Y��>���
�j��$zv����s���x}>�ϖ�d�PՆ	R���}.J{�k�O�I����Dtܤ�YĆ�e_���<un���Ζ�d�����^�Ԑ��awu-/L0��y�s�4[�ód	����"��&���eE7���{Жq������r�X`2��7)���ɍ�q���P��x� C�W`�-��V��d	y����Y�����"���Ȁ���Ξ��ޅV�����LWn���Κl--��/v�����޲ɯ%�;��u����گ(��w" `�G�vI�YW5S�J�LQ���]r�GV��7�r!����t�"�Y��ps��}�\ 8���/��o5�`�:}a��7���ӭ>�f��<���-J	��ɲ)Ï5esg����|���. �6ʏ~�gd�{/u��<��15�h�Bb����6Ed��n�q�[:Z0?�)��ҡ��*')�\��V�iS*=����o�m�]LA��O���Պ�=J9V��P�i�����x��!8QO@�ձ$��GU�Sg(n��u�n �䅂�hA��
�%$_���&�8UX�Õv8�-ڳn9�[��H��{P �6*��VK�WuH��6�j�=ތ�謌�b��E%Zn5&�W�mp5W��%�{0��s0���یn抇���!�k+!`�\ȑ��"8r:�
P��ԭ7�����r
J�� �.��x����ϯOb�)�����O�p2��4/4^$�=
.��Ʌ�7���I=�JF�f-`(J��Zk3t�T�B��ұm+l�8�Mj��[PC��+4ä�`J��؀�/ڽ���,��=E�t�=�9�ddI�i��>{�?I�0n v�m������V�X�����'u�+yS�4���5��ڗ�Gd���D��sGN��1A��M_LO��J6���G�uZ��M�'��)4���y�:�	�P�D��E�4è�=g`�7qc5��+��²Ly�,A4"n�G�ۭ��<[��f�r���tJ��(����	�x�{M_
��vn�\=z睞�@�(i\���B�N�����v��b��q�ݽ�Y0�3OK]��M���(���0)]e�}��#�N�`J�ьZ�XyG�Q��͂�(2�^S��S���s��K"M�w���<�p�r�Y+Y��}��q/���_^W.`���1�W^���5�K�!U���=�΁�s�<��'��W�A3)j�Z+H���=��"_�Y��^^��mlZ��N�����jU���s=�v�܇9vt`�]e�E'���u�t�nu�Rm�&��"tR�C) r��x��P[NOV:��Ǭ���ƍ������ ��Y�)]n�s< 7��s����[�Z.�d\������P[⚩vm3��L���i�yDZ3���lb�Lǁ�[�x�#nƂ�7�q��c���Xˡb1�T��친�*�����ur�;��bW�v��p�]K��wmoZ��M46�kV��Ȕ��Tb�"ͷ�?E�0�v�W����t�jC�N��dWu�.[�J���}(^���.f�����;����)�á�9A9�󧖝���L2t��}���=!�yv�X�zЄ˰�iaz�M�\�Z�f���q�1�g��o^�jgoW�-t�<2�yr��N��qå�j<"nmm�0��aCI�E.�ӣ[�ff�0�6��j��SJ�K�TƬ�*%X�;t&�*Z�q��BjN4ͫp��%�q�L�p�m��(���u>)1��(P#J���,�����F*���\�K$UCZN��ieK���bQ��9��4�4���D��
UW*U7'vt9�W6��{tKʤ�\�RЫ�#��YR�D�X�F�Q]Й�0�)29y��`UU��"�C*��:�9N��6���DU[���(dz�yNs1H� �B��W75
0-hiP�g��U�N*98E$�9t3�9���H��BeFI���9�H�T��Q�B��YN�9Yi�:9�iiy:a	�Wv����BP��s)�L��BMM��R�Y��Q�^��GL�eb$JЫOC�(�R�
"L.�R�wu��4�/K"s�1��A�*宎T�h��zjs	f牔ANF�)���QsL�n�.狂j�E�ʫ����{T)�n�az�NnN��s�r�,3�]��=�*q#J��?"�UY�i��ܾ�o�Y�i����*0���w���I���z]%�bC�Ǖ�{��nNX��(G%E�u��Z�jܺ�� ��$�\IU��v���z ��?�c�=@©୑7���]�x����!�>���yw�S���!�>���!�{���|q'�?��|S���w�w������<~M���]���^�'i��2��o��xC \�����_;I�!;����������y�����aw��X��]*o��W��}N|�>8��pN������󿓓HN���r�����)�S~t�ݤ��'׿;����ڗ�vޟ�",����]�������'��Г����~�I��:v����� yM�N>��~�����{�oR~;H�;��ɾ�~��J�\z<_P�����n����T߫�5fBۓ򞭺�Qy7�����x��7���>�����U��������|������<�s���m�<�N���~����8�9���r�M}���ׄ��On��=x�;y@��@M!t�W^v�}�n�B��{I����{v���~�/����{�{�������o�]���ϼy�������0"o��s����8$?#���s�Np|>\��9>!�"D|�oV7qUz����4�舐B��?#�S�i���U�ɤi�׎���xv����P����C������������!�5�}��yq?�I�߾�ro�J�����~CҸ=B;>ߟU��Y;?s��f ��=#ޞpO�{BNq�ޓ���7;��{OG�|S
����C�=!Ʌ����xAw�v܇��|��o�Iτ=o�=��P�N/��Ǉ���z߾��>���p�*���Wj����ٙj~���Z�  ���0;��G�|`}P���i�����o�x�=��ӎC����ɿ����S���y�X��)�]�����<������~���!�� `��@�1��>0"�3&W��d@�$�f?E�}ꋏ�� ?�6��8���?~��0�;w���܁��y��Ǎ�w��������Wo=�����s����<!�4�'���ar�?�=C�������|�qj��mW5�>���zG��z"�� =�>��~Cӿ8��oZ��;��P�����nr�" ����� \�E���1+����>S�������������?�]I��mɾ!;�A��?�oǷ׿'�IK�lz��Ff��&E��'�f�<�,57XxqK�v�l��oU��ĉ�]�5�ǫC������T��2mߎ�p�ɠ�BA�G���tP{��*{�k8�vt�=��r�p�S ��2Ǜ�g�m�$5w`�oFU�����	�: |EQ 8qP>��Ϟ�ޓxt�����
o�'Ͼ������{�(}C�r|M�9�^�������r�߽�?!�0�z��9>!�%/��?r&7��>*���{#<�Ay۬}P ��
��d|@<���{Cˉ7���\{���Son�����o����}v��y���������oz�h�����z�z�G�\���w�_P__��>/�����&���NM�	e���9��y<��ԝ�x�㷷�n8�9=�����~�w�=&�~q��~�=~��n@���v���v�\o��"(C�#�O\m�Q�TXݝ�7��{����2>�����G����v�>Ǆ��o��
xM���M��90�����x�}v��'x���.�㓐�F�|w�;�oo��}����K(8`���q�~�=���X7���Y>��~��F =�<G��BS�"�C����{�SHH&�~��ɏ)�!;�y�w�1�|OE:q���@�w�i7�J��raCޣ�}Nq����^�cЄH�|=�?��$2����^���U����0>L���}�@����>7�zC�}C�����ۉ����~��!'��{뷔��'����|(������x}oS�*��V~�(���+���K�Z�w��h
���L|�� (�������<�����~��~OI���l���9��w�i&����~�<3��r_�޻P9'o|v�﯇_	��6�}HUh���v�D?N6?�篋/翟�r�&�xO�ly���r�?8����w���<v>��>�{y��{�S{B�y�>��=?\�&����v��<&�w��n������#r�o������#鏾0`�q�0��9an?{4v�����<�!��q��������������y=[��܇&����U�N�|���S��O���
Ǆߐ��C����ě����?;y�~pp����zǈ�|�s��ubD����Y�������}v�ys�M!&��c�I�Ƿ��F���=�8�����yL.���z?��{OhraO>�~w�=��9ǯ��q ����~���I� -ȸ����|��.=��<Xڱ�ۗ�d�/���301F�F��I�-H���{�2my����ܕd�W_
�����L���&�#)��j3I��>���?����o�q��1�����sc��i��M���#�P����s���8�I�!�ho��N'�k�^	)��7�nEӴ���m�ܮ<�&�����=u������������O	��_N?�	�{������»|I7 z^zY����Cx�Ϲ^wD�c�q��O�����8��'����&��O�<�w�׏߽y7�=&�����ɤ�"���ǿ�7�$������݁M�	��;�������!��^�u��2��(}H����þ�_�}|;�{��xW!���Ǘ�;�ɾ���=��9�rw�߼��w�9<��xhxL*��~���S��C�=o�߬r�&����x�-¼v����럧f,]���~��ohHyO��<y�����;���ps�����h������7�~v�||�<*o�J���ɿ��s�n&a�@ z P&>���@��� ��W�DH�#�/�C/�i���������/�N����s�o��4������a@��oI�z�	��v�ߐ�X��Ï
�@�俻}C�N'��[����I���>��/�iN��~��}C���p�=�&=B=� ���7j���}'UU���~��=DB��lG�B"=?o��4�M������+���{|�-�0�����0||���;���\yw��n!����®������7�9= n��{����OowH��q��׫��Ĝ���������7�$����󼫁M���߿�m'�ۂC���7�v��<;s�}v����O~/)�\��o�yw�i���>'�9�\y�w(d�G�>p���P�z"ܾ����_���=&OǾ�ۉ>���&���px~!��+�!��z�����}|��|v������'�p)���x<:v�_<��i�N=��	��;봇�1��7�%M���,�x��u�s??�� L|:>��> �����?{~w���]�?�?;�S�����S~t����}��ǆq ���?�m��I�w����&���9Ӵ��	��>����}��~����k����!��՜��_k��",G��~��O�iI���	��|���+�>��<&�/�y�;|t�pHxw���?>�}O�ɇ���o����A���p
�$�ǟ��)����/<xC���!A�Vx�:���h�AmA�F�q2-oV_y���%��w��y��@Af�-k�k)��9�-���r�`7m^aŕ3���-+��gi�o�r�_�5����w�R7��{��g�'Q�������{/0m|�pM>�Z��;�qnD�����T�K�}���z�7>Ӝ�Ʌ]����<{��@������� �M����S�.ߙޟG�|o)�!'�������W�����_�ߓ��	?'���v������c˧k�y���W�W3af&�]��^�p���U�G��7�w�~v�ii�w��x���;�y=G���!Ʌ�y�n$����_<v��}q��i�}��C󏿯���ɾ!=��U�=GW8�=�*a:��DH�k�I�>v�ӧG���Ʌ��'�Ε��C����{Nq�=o��	�{N�c���������|w�>'�9�����:C�{O�xL Ǡ���_C�;U��<��1�-$�b��L���N��}��}C�?��3~���_n�>�|BI~y�����zC�Hy>��<<�"�YM�ݷ��ׅp)��{�I���F$>>R>#�"�H���h��i��B��6�e�������oO&��~����
��'y�v��_�wߜ~ON�r��x��:w��n~�������Uޯ���7!ɾ!?S����u��H�~d��_xU\*-���R�ޤ��R����@������� G�~�a��1���Ƿ����ۼG���@s�õ�,y>�����Ʌ]���O�s��|?|��Ӄ�S��￾xǤ��]�߾��9IHUW
 
�>�+ETH7�	��Sw^�Ӆw>��
 Q��������z���ۓ~w����ךp)���xw�k�p|��!�5[x�������;_߾�7�yT������4�Ș�X{��\d|��>Y{_b~LN�w2�z��s`}p&�
~� �� ( �s���:C�?�<��<��w��n@���V?������y�yq8�������&���C�Ϗ�ߓ��Og��oi���"�<���x�c2�Jwv�m������E��d_XY��������R�s��ϑ���ϱ��]7�-={I��@UQ/Lb;����O�����u":l���tz����)x{�Yo�^Rv�u��s����r�9�1t	�{�������$͇B[d��Y�Z�Q�nL��
��K44q��H�F�w��{D;��|�։�]��5���cx��h���pcs�:٦L�i��Ug�Z�墫v�'���e�Ay}��*�:�A�ˋ,��{ǹ�[zǾ��F\G)v��3v[�b5�r����G�db 8h97�Y��]徕o�����gA��}<#�D=�L�D�V�<ܦR;&4R5�3T�G{$	��h���C2[Z��͝�=wt��n�:v�����R�w���lph)�8��^���v������O�"mO8��lG?8�F�����x�C��<�ݝ����l�{����0�i�o�&rؿl\s,� me�CѯTwQ2��4��Y�&�zN�G_\�Om ����D�Ǌ���'&�����(�E���1�UtТ��9�\��ף�'�״5���^��q�ˈs	��wXcw��R@E��(p�0PuB_��G.�
�O�(�ȟ�yh>c=�!�7rf�Q�1~.q$��9��Kf30���0�λ�38sm`��暮�Z��~]$:���׶�j2��]����*����].�J%1}�l렱�aov:�'"8c��]q���.X�8�F�Jӫ%�	S�ȉ+k1z��*�{��_X�W@��}t��ښ��
�i��1��Ur�|a�/&�{����dӸ�N:�qQ��9u�(�E����wR�C��n�{td��B�����:S�J��:����ie�P��z����-��x�'�Ҁ������p�+^������qH����Evk�+u�3<��:�������W{������i������Ou���#�D�NU����~ұ^�y�E������z���fz�� 7@ed�o��!�᫃����!�rí�٠8?	��V{��a��sg7=Y&�8'�+�~> �v�ws�>��{)��L0j�`�F�o!��ε����O�eZYʎyp��}kܝ�m�&{����U�}�x�����.t��ƛ�N{�K��#l?}����s1Qs8����J"R��7�����pKد�]D�{�y����5����J�S�U�}�8dzzk�H	�N�d�a�,���
���,`��p_2F�md��Mt]#˥�W|�l)���sN���:�\ +��2��e���ڥN�IW���U�p�eG��1�~�g\1���cw]�a��b�Ԟ. %"�ϧ�#�����q|��I�g77�v�n%GVuA��>p��q���n1��J�j��:��n&
TQ������bT����#S����GG㙸�F��}ײc
P믽�0]k4f|���O4P�3���F����	xj��GqB���;�І+]\a��j�w��*{��ݏ�ѬK4XM��+�Ք��2��lW�'~�����Orv�6�
��/�cBә-��i\M�L�l��8 ��I�2��8��_e����@�B�Q��T`�鉍˖NWL1����9�5����[��&��(���Z;��i�e�{�r i�t�|����^&�S�t��/��������y:�B$ȝ�˰��T�]�$_#���UL|�|��>�:�o0��"ꥮ���,,gة���,�w`W����Ɇ+��uA��6 	�r ����7<Y]*��@f���o5�8�����q@�L--���5̖Q�U�+ޒW��[6g�5�:K�ٟ#\%�LSM�~٫���G��:ߪv������1%�|�r(����og��h@���v�G�$wRa7���Ӧ�%V��"������+T�Ϧ���Z��{M>J�Xf�X��Sj�4����q8k���]�W�U��|-b���s�к��)⧧�a�+.t�9tjr=�����..�G
4��p"��J�Ƶ��Z�?��X���*.���Z��M�^������]`� {�'�=�"O�P�|^�GCe�{�B}��ͣG^<c�����%���h�ٱ��>廡�A:�m2�uk�+�:x�ue��{�7{w]?�[f����7,	���<�8����3����w��-w:���?B�Q�]y�{��c�дf�S�xw(�Գˀ�1Ȯ�`u��Ck�Z��W���#o�x�ʽQ�����3��
��
�To�WoٗהD�\�ʻ:Ҍ�4�vF|yf$<��.
R8=�0�c�)׹�[P�;>
�\:_�r��\��=v�k �~��zx@��F7�xh��N�1�:[7}�iuC]kk��.f�����(ʹ(80y����)����'��8T��XJ1��ƣ���Ⰶ�]��]�,�i�|x��O$�^����R��:ùJ�o�|M+���Q)�FPw�N�;"U�$Pfo�׊t�Nk�����Hn���1K�{�H�<]S�x̪�U�3�'�9����R��t�i�y�v}饐܁� uCx,��NH�&ޣ>C%�5�Jϒ;����ff����>�wRe��c�baTrO'>TG�O�I%�vo�P�Nla3r^P�N;�LM.��P�k΢��8�&��~O3=��GGC��p����(���.)��PUw�i��ժ,Z�:�G�Y��`�g�8�8�A�|I^I�&����[5q� ��۫G������q	�Z'|��y���/n^zOJ߮��=����1c��\		�ySΝ���N8��ѹ��j���ut�:�MiT����ޏD��g"�����w�>�lX�1N_?�R�<��[�cL!���eV��nW�m(}�v���.6��(׽y8*Z�[U���'Gj�!�gS�LSrF|�,��h:p�|���jD~����M��G�����_KU�y�$p�VQpk sօ]��*�g����OM��=��D�5����鈮��.s��D�j�~Cxog�9lɹ�J4'���%�`��[T�.�g'OJ��v�y��]o����:v�iQ<4��]"����}V�9���HCa3Q)Յ���ߟ:,�v���/#U@E:]ulf�4ts��{]sD	��r@�%�u;�M�O!ḋ����h�T		����	�ꬨJz��^��'�8َ���� omS�D�MDY�V��t���V��>����W�O�@��z�i��뗶#-Čj��u��@�A��̘)О�A|K�5�Й���6�eW��z��4H{YK�D'ԁ~@X>H?�qu���^tj��҄���xzМ��ͱX2�ҕ1��4X�w L����_��^q�7��Lѫb���֣��C�ڧ���4���rD�1�x���cFw|T��S��{]���-~�vU|�]7�~��K�_/g��C)R���S`����B�O�@A=������j�9}U�U{5�������'7���
�M��&!��:���[�"��j1.)ѣ���������y�,����4�3�T@#p�G&k�����"�rt7�Ib ∉&���ۜ�w>ި�����P?}�z�h�4T���:���zn!�&2�U�Ɍ�>zj%*��u�4������ݶ�$I~gI��H�����X�J?F[���Ud�l�S�XɌ2z�k+21I�t�/P�}�o�FA8-�>�{NE��8��t�U�/��=J�\ �����R���9�^��{��m{Q�=č~T��v��#�JK�䥎������RՌ^��t>���ew�Z ��?.'��4���8X�21)G\�1D�l�,�Z�\��:̐����m}&��Y��ߗ:ms�M���7~�Pʾ���u��D]���{�Mެ��o�{q����66���ɝs:�ν����k|}��A�]W�}>ԁ��YPAU��V��<X�����;qT���a
����v��Q=QA`-tCj�^�W���a^�����B��Kbjz����A\��ӱD���@
=��v���\�x�p[�Y�� _^�����:�yu|������x��ڀ���5x�N��8@׭�cVoEܭ|���|�Ц�죵٤�]�]�%��>YGdo*�Kg~~o����Ƌ���)ds�m��\�ņ���4�qq�k��ˁ���g+���^�a���<x�7�K������� ��{��
PN��"�i�ˠZA�4�'O�)����	�Iʾ�A������z(4.)C���tᬎ�1[���Vc-e��<W)a�����;}5���+n��(A����E_��� g��0�K�$����h��^�*��L���L��|��jろbk�Q*�wK*�%f��ޚ!�뺲��߫;�6C� '�"Pc���W�b�s6wbgj=:�޹:����^��؍���W��Nn���]0����p���T팧�
'Ŕ=�O$r6�l^�����&
�	+��G7����8	�w/�Y��r��L]�Y�z1n�>ӂ���c�'�Ja>R�m-w{����dGq�����F7��fp�h���y6L�古�n����4�N����]t2�.�g2'X�ƷS@��8s���{-�̦�*��m��H�g��2�V_/�yK�TB��>Mw��r߻YZˋ(�8-��NLu�* �]hѮa{��-bԈ��U5w�ߞ�{��&m�����O޻�)2��7�#C�d�Rݹ�1Y�j
V-�u�C�]�"w�>EA��U��WF������ۺ&D�f�+�S��-ӷ $�7p��4V���jģ��^(α�T��mKU���0m�����#�6��BR�)[��,��TV�µe�DÛcq�X�
����E�ӝ�#��Rx���W����ks;{�Q�ٜ�`\ ��<�͝� t�:f�cҹ<|������w�t���-���Z�3�.ɣ�L9�h�zxMk�,�'�U��������%Fܠ��d{lԎw/IokP�� Ԯ�I�e݂����E�;�	F�i�/�.����%��e�����9#�<�sw< #�Lܕ6��W8��t�Wc�����1��-�|�t鉥k�?���ۧ���V�\�<\\�9�����VrЦ"^<X�\�O���V�5|,�e+��쿈6����"����I��=�$v?6N�e�<ȃ2u��=� ������4�ǔ{H��"u)Ł]�DÞ�]Z8����<��^^�+�� �<�p9* :���vp�#ڷ���F��Omwg�Ʈ��Ek�j��$��p��&R�BۈQbK��=��=��x�O�(!�#㸟Q@��ޱɛ�\%�=�ݝsF���/v,�'-��=n�����
��c"e.��8(K���mx��R�`Bu2����o]��ɀ1���Sq\2�;��29�n����S��o����R1
,�%$�Mܽé��嚖]2'qt�%kK�]ۜ�O*���=N�=s�{����[��E��;���p�n�W��g<O\�6X�c�����8����{�n�yY�eŊ(��s7q�'V�V����]��fԱ�RWfx���wd^���9�IԮb���\�v��D.��p��%�s\\�N{�z�)&�m
���H��:R*�$@G��s�N�Q�J�ij���&YsZDZWR�H��nc�K��gHD#e����JE�f�$:�뻸�a.㺐�N�)Ȭ5h�l�(S��%���3:N��qe�V�`U���Ne{�����̢D��I"D��E!�9�v���J�&a���Pi��p-�������asN�TZF��%�sT�i�媤�.jF���E�E��D�'��7)9K%i��=ۘI8��ͪn����-�XF�"��3�t�/�)9sw��)�C�[��I����J�7��ڂ�����	��n	T�e���p�țH,qJ~�z=z��\�r�����Ҙˈ���]Ѕ{N�� ��>&U��.����{��-X^�F�nzT]�˯6ow'��e��Uw��lt�ߔ�SPLF��@�q7�<��v�0`0'ܔu��&Z�ã�vm��]B�%���`hu�G^
RC���������]D�&�{td�&WoTr5/�}\��Ga�"9����~U�"��� �����R�����r�h����{�T��Ө�1�k{i3x۸���	��s#���U�Y`-�9#Ue�X1wv��J%Ęcj&&��2��/�.��Ȅ�8m�vG[��1jg���$��Imn�
y��(�=�6���(�I��M׶���bFv�|{acY�bU'�{�Ei�̬�픒]����rLXt�*�%�})G]����O,E�\!�C�*�Ў��iV�@\�sɶ"�j@n�{�(`� ����6'����h�Q�s8h�Vu���-Y��>�B��g�̶1��e���wɳ��-L����<���o�#*� gi��Y-���J�)j�k��vZ6&H�oM��,*��5m�WP)B���2���{�]�v�o���"��&��t00�P���i&�Se�B�n�w�vOdNBq��}��%�rְ-�v����Ѣ�L��Ȕ�
���h�T�{ޏzށ��*mŊ��p��Yx���`?R�U����W�'`00����8e̔��{p4�bC�c�TNV��ʯ;(M���C��c�L1'�[�ӳ���:�U;iE�6鋄٭ H|��{e*�!Vx]��(n�W:�����%�<!�|�Ni�ݎV z����g��Ag�QF*�.�*��+%]�Ƴ�|}�$���2a�� +�ԓ�X�,�~��|_9��^��97��n �4xw"��K<��5VӉ�M�v<��چ��ew�p����-r��9�c��.�YAB�^}���<�l��(��s���[j��Vc}Z?#�������~�(EzӶ0ܔy��R����ϳ�p~= v߫n�,@��A��[$uD)�k�xٍ��\ΏX�j�ѓ�W��;W �GK�Kq{1>SS�h�g��0��-����ƣ��R��`����qi�{;Y�Y�\��b!O�
��11ή�14t<<Oq���y}U��!���|u���Q�ε�վ){+K�����w�ѴWg,dJ�<�Oa���Vbѐ�ԡq�1��֦�.Ar���Q6��ڲ3
a����|F
Zl��&�h�S�(�������<3��p��8� �x@��sNz�C���͎@��{���oXm��ї���=�b.Y(��V�A�p�%i뉐��bk7���W�@���L�q��:y�{[exL`���1p�U��[�#�
 �o��Ȋ׆h?p������l�!(�۱��6}�W���r��}n�̴�c�P�����mu�� k���I��3J�U�=��}"0D�W>�s��i��Τ�Cy���1h�o��M��p�3�����F9,v7sv�P�,��д}�����*�.pP��T�����1���Z)��<\�v�I���:��9"a�{gLs���pʜ�B�e�B�0N� C��`p�&��,`��Η�3ܑ�u�P�j�����:���@r�|�X�-ߍ�
돱��օ2���89��鸺��l�8Ĳǭk�M�1����E:�tz0_���":l���gG���ƌ�K�S۫�]0Y댙��Rc3S��xp�7.1�>6�)�Q�ٲ�����u�m�kjw-�c���m�ü�!���	���|K+e3�C���/]_1��7�����y6{h�Giخ��udЮ�r=�v�1���N%�p�t6���^Y�^̛힁R7w����8m���%�;l3���*���D��N�I�ӛ]n�������j+��fms���Z�^�z1�pm*�޿��Ͼ��e�Ļ���0��r騝�#�&PS���O!-�����8��wL�췏.�WU_A#/����C���F���(�z�!'",�S����+u��D��^��݂��w�ƹv��wD�:ۧp��g����T̄����A�K�
���eH4Ӡ�T�~+�={A��B.!S��Cr�l�cuHШ���:�H�tМ}VJ3��u���f]��wue��wr�1Q	�q7.��eG���[��d?�.Z��.(Ҟ����C��%q�~}�x��]�`�;�"G&k�ڸc ��fM� uz�$�V��Sy�5�aqˉ�b-����8ο#,m��c+�9���s���8�r�ڊ֬��Y�s����$��r|�`�M�l�V9���Mn�u�p�-���˺x�e�Hva�u�����jQN�<��?V=��"+�� W���_�2�{7��t�X��}8NfV���>��0���X?��ᒒ�9)c��~��U���-�E���b�6��Gw`������͌�A��i�/m�W�3�nl�l�W�{�Po*�~9Y�/z���&�[�вD3�˙I�;.����[͟ӳ��Nw��f���c�6�+`^*K-���4I���]�y}��IJ�s	�Jz���Z���z#��m%B��3&8~��G�OS (�&�9��j��{U�bW��L��Z��{��LX��k��.y﫷Ƽig��b��v��l�1܈n����lF��;�5�v�:r�;�b�Ǌ��`�f��ɝs��HE�u�r�l��i��	�V��l$�L,y���U%��ݷ'K�#��hʤ�a��NV5��k�:Y^���aђQ��I�$c;8�, �"�e>7�5�m�}q�c��|zk�H	�N�d߰�
�]�|�eeҞ�W*s���8�H6l=�C�
\a�g�upC 
cQ
gb	��^�@�J�� ,�3=ٺѾ���֦�v�tP�9��^�.��<�.�pX��v��a��5%�wMA(!%��[�����=��{���Ɯps�PQB���
]wn@�F�ح��&�^�~
��1f��ӄ�1* .�~�ޜ���3��u�&8{�}��i�4\���U�F�v��b}ku�
��Y,��I��11΢.���0��t��yѕ����[��8�z.)Y`�}�ʄ@)Z��v�:^��E�ZO%���<�P���3��"3`�<�Bi���Nu���F�(.��a��:��c���-�_<G�d�ju���[#8�ʓ����jT�z��[���&5ή�21�V��ND'�S�:�V��z=������f����l��91Z�� >^'Ih��-}����]!�ɍބi���=3/y��JC�QS#���3=�{�R5�P�>�����:�V�>��x7�5t���s<!�Z���ٱ/ٶƋN�1~
L!M��x��x] �|���.|T�}X��*�M�U����=ָ��3�ʄ��廌k�֤�9��0�T;�����#���b���@ӳ��ў{ӻ��m�#�WM�g''�f�L�LB�t���D�rt����&u��q�Uiͽx��ag�q�j�4[V�.U�+\^�=��9�B,mCڄ"��ֳ��|����\d���b�at�A���)�͓�6��e�½�W�vxKJ�P� _H\��j�����{կ��(@c��1\�ۆ��vy���^`��ɋ��f����\<�}�бc[�}��s���ꢗM����o��Z{��c��l�����bS�xo"���v,l)W/I��wΚ�΃Y�81�z��p�Ȕ���K�-�[u��0Nsg�VȬ�������l��ts����Ө�v�B���]��,s�Qt�m�e�d>��"�W�_`��Xoh�֝杋����`8$۽��{��;��{�Ae|A5`V�s�������=���S�H��;ުQ�o�)v��֭wn�Mb� w�.���U}���I��X����Y�o���Vy�jb��\�\<�2�g<vaӌ��4��'�!a�z����8u�!>; k��t*
� W�Ph��Gw�O��F8U̾lm@��)oE�.{��Up�8!8*O0{�0|��������ʨc3�,*���JȲ`�j3x����[zČ���r]l������Q���P�;��V��K�pz̮�H��t:��Q�����b��5�����u��zZ�p�����<�"�t����.��>��O���m�X{��;5��U�7_���p�LN��i�)��y +�ydTBrDo(�js_G[Ī��
�ֵ{D��C��[&��_G��M���͖Ԁ����~���@z,�ٍ������l����
uz�.q���35҃O�3��`#�Ok&tue��fr�y��ed[�� k®��
_�~4)!�+˥E*`�΄�V����VS�� ����{;��t`�=Q�7����OX�J�Z-ҷ\T>��}B²�9�^���mZ,�<�ft�N���t�wr:�&nh��n�x��[+
ڋx+W��ggMf_]�Cvz:�.��wP�?>���A�J��;�Ь΂���	�g�%�lms�\;�͈��s&�G6J��Ɨ9S�,�sG]/E���< �}�>���r�W93ʸ�r����(�f�p��'@��1X��O)teC޿H�[��_�6`�=��ߍ��B��_��v���V�>�װr�h��u�>��tɿ3�jx˭�q�n�z;ߎؖWٝh<�S/��D�@h�f?^Ĺ��d��R�زG#�U�N����v�:b;�`׽G�^S�.��2^�	���wy#@Xq�@��V�7��߲P�+�TK6��vK+�)�������X�W�L����������5�պ���@--b��.|�s�q���YU!�4�ρh��b�]�v�<cR{b(�/�Ҹ�4���1²WR�]@f���&�i.���E@�0��×�f�����&Y�gN�\C����`a�j��m��@�qU3#�2`�'��4��vg�����$��6+c�g8θ=O.8H�N��C}Hx�ҙ
Q��P�"7\\U��D��}vc�{�+���86��y����M��L�AyZ
�:@�wDR��Rp�8�ز`����Nr���,`�����9��[=�`�k�5�����������[2��PقV����kx����m]Ԗ_޼��f���:�WC ����(��;sC�:wa U�AX�-\y��Z�v��q�]{i�%��Z�ug|u�F�p��]Im!��=t��j�W}0��_UUW��gS�� ��� ����iWt�W��
�vvg=�ޠ|-ד&��f��Y��S�K#��j���c�M�}|mD���I_x�;fW�����ՎEሺ��vP{�N�9��N֭��'u���I���K��sU"+�ey�WD���%qۉ{���$+��!�G�9����9�>�sy!���W ��,1q
g��X�[�,J����#�O��9)c���uMڈ�Pr���<_y̥{^y�	�����哾Naq6�A�Lޙ�����ቶ�ØT�X�e�x�i�Ct��<2���KW7����@m��l��1���:�	��x�7R�iW�Å��R��d��E�������*���
�]{/����L��X�\�Hn���u9��e�@ɛ��-�u ڬ����_E^�v��+ƴq�Hv�U�Κ�R�]Π3,�V�ZqØ|j'��-��ϲp����U &*w�&��A��p�\�(Z����Kt���%1ĭ1~nX��
�	�cQ
g ����+���dѭ�Րu�ςx���V٥@����مW��2�5m>-�c}}�w=���n-�ݔ>9f����|�K����aW��	�<��������}���I8�{�Al�Vk�ލ�Y�|<4Θ�� u����l6���p��m�ea��T����ꯨ���3伥E�	s�_��}קΡ�"�8\b�zw#Z�890��QހD�ǁ�e�� �O%;OFM�ױg�{������.�(о��D)u�r�#��q8*ݫ��Ս���oUk�	�֣.N����"ʗ�/��7q�I��ۘ�����7]}���#���SП>V.��~�g�p;��O#�F��.���F4e{��:BwLBף����:������d�jf�.b9��r�:I��G�?��4���Cs��`�ۇrd
�v-�K�l�q�C�*9�g(��)��<����`-.�裮ص����Ŵ�q�Lv��E�Ruٿz[-+4��)0�j@{�e�c ��9<`6�1i��[������fi��(Uv�߳i�oLp�^��L�y��7U,�P��a���2�ȑ�"wko]|��������1��l=��ٸ9���ga����29W2��nN���{1�h)T�&Ʃ�绔p�B(��P�%�dЎ�\�Xn;Us����z�§�A����\�-��P��͛M�T�b��O%��<�G��v���%�$#U�*�v t���Y�7.�,;Oj� �*Tڼ��䆻[��t����VU��
=m�08�H�D��؃��O?Uٲ����; <&��eH�
yQ�b-ޭ��1�V�T$�w��Y�9I�n�o��c��43�_8���Gt���G���-k��7X/E-�{��O;K��X$��x�5#6܎�`泭��>��Wb�3W�%iJ{���#�!O���ɚ<�ݴp��^y U�&Q�1}�(t�����W��<��>�-�}�ǧ����\z���/6V���"b��7s)�u[����ޫ,9��i�f�R�˵�Fb<�Dv��/(]t�O�X����Ä9�b �"Be��69���:m��?,!ie���f�.[�nd��"�4� r�"3WK�쑅�Y�n]ۥa������[����ǐ�WW|Vi)�� ysÍ��9�8Ao�B�{t�~��W�x�10��:]�&+���ʺ?c])�'�E�����A1cq�É��'96���wWhА�����AP�7k$}J��6�奿W��bg�2��Ǫ
g���򌇎n�=��\u
Kum	,|�p��؛6;���̽-+�P_�F�C���$ӱb��k����Z2-�j�P�4P�Z��okvG;o��G�xְ
�f:OFK%�[�s��Ek{�\ ��������w��\�,(��s�𚫪0�[O�QB;{��@��+p���[�ƺZgL]��"�,Nv0	�u%Ƴ����i�����)�;�D�'DAVn前�7��췿��<<^�｜�Ժ�m��w�N�M�V'%���y���P�Z{n��K;jq���#O�Bp�~ ]pި)�4�p��.��+5I��cU]������/��E,�����廋���ј4�ڠ0� ��$����B��������k&@��2�Tj�t5������X��ޮ��gE2ɡW2����(�3hA/��^����j`�巓�ys+gK%:ub�^G���I�F���$�w���ɃTMۇ�򻛜�<����WY+x�l�ۥ�ήa��說}�Q��f�.�EG��~�w�������OW���l�;�f��
|6���^�t�����F�<[Q^�Ҟ�qu�#���#�g���yI�_!�9_�;��9N�U��@q���N��GR,ymgi���'u:��f� �B����׷�@GY�\���ڣ�V��lq�Ew�u�=J���p��绸�	�ZD�ީ���λ���*|\tC�;�$ׯ���,yN7�v����}�jU A�h|A4y�B��enw]������R��5/rJ2��0���S�U�\s��n�d�]�G'���Wuu�Y ��f;���y"it+�u�sМ<��H5�VWwwP�L4��%���k6f��CD�Oq.�g"Ww��L$1"����-���y���P�{�F�`���ғ4�$�SIwnz�l�Ȯa��ꪩ*��ۓ�n��t3L̲7uԣdn�D�r�r�īC$�h\��jkI��"��J
�3b�����!�1ұK�UF̑1,��֘�䋧�TF�J��w#�42��.��K9�!�s�+��eG"�ZrE��N�����r*��j.{���l�Ta�2���&y�I�i�'E]���dQ��Q�T�QK�VU��zd��%:B�R��绎����[\���d��L<�{��zes ���t��ǯ�q7^>X֪���3�y��e:a�v41J̗���5���r�7��#ވ��5e��[��ҁ��� ��ƌ���Ck]z�+���vxJ���о _n��*!�n/.�����;�R� �}-�TP͆��w���R�{�j
�IWx����[�=���v�V:%ⱪl��u��f'KJ�Σ��cT�z�v'F���$��ќ�Ims*�1r��~��`Y���۸L䦯�Ň�Dk��vT��B��C#�(���P�Q�3<��Z���I�=�Z��O�xS��ҫ�0t�O�B.�:<�a�r�R�x����M5��1�+E9��T@ G ��N�W�� Ve ьӣ�OQ<�$bj!N�7�xg<�V*x�.ؑea~*c+��k��(��>�*_r��d��G�i�J�Vj�鉭iŚ8�9k�w��4�޵�U�{�j
�ǉ�=�b��ut���:Ы��k�m�)��1����S�x8}4"�r�`���@w�q��� ��zd����i�.3��ke�k�j�z�=�zez�\6��$�h�7�l�An��P��d&H�w��R�(�Y�B]��e�����~�)8O��C4����^;}
2��i�B�m��F�{@�ԐJ��5oI�xzHN��XU{�ې��޳d���q�M}_�K��:�����[��.y��xq>��Ak,��}ũ����gRq�[�|�f��gFCY�t��7���UUT�����Vˋ�3>3�6�H��Z��]���9�h���F�th�5 6lK˯owc�oy�)ʋZ�p$=8N����Hc�ו�W8̌i����y���s����)�D�,�����[��W���ah��tmp�5vy���K��S����W���瑣����/hm�@�Ӻ�G�L�G��b���`�
���^�G��`�/^Y9�NA5}��n�P�ةJb��/��!�ѯ��!�W���`�=ʷ~7V�]a§gD�m'��ђ"�Gu;'J c�G�2W
^x��2�����r��f�	=�T
��o�[lnz�+k�~ۣ���C��*�g'OJ��v�n��r���[&:+7j-�Vd%mn�	���"I����/]¸�B�-�L�D�w��
�7)��l���U�9��)i���W�e���^ip����EzUHvӿ=�%������x���%�7l�p6�7	��j�߸P�#5D�#H�T��q5�<�ٸ���a�b"�=���̂��F�3��>�G�ӖV����r-�sdp�&p�%'���Ѿ졘z��� ܤz$i��vxh� �`m��Vo��y|��/:���{���.�V�Ņ�}r���%�ՊO��Z�秴L���G�":�5��=��">�vV�ɻ��ӹ��>n�C����G��$����f�)vy]�������8c��ᴲ��Yq�E*u�r�D��9xy�A���`<+�Y�9RT�����ӻ"��4(��ÐKGw�1I�q7�7��k� E>�&��������0��2�^0XTxxʝÃIL�N�rf��L0�.K/��|JgK��O>��w=N" ߼*�\�?V]!�rB�1�}1ګY�e��4Lf*���4�c��'���i�=0�|���\�T���<Nٟ#X<�M�m���.X�5���'[��bB���MIA�ja�2#a��;�WDZ������0�u�][��#]4�s}�W�k�\f��f�*R�jfV���>n����O����W��O+���e�ˌ¢�]z�y1���v{ѽl^�钙�8���i��"��0.��?hۥi��眜�!����Y-,{RR�q��<�^��ퟺx�V�q�����D��vj��X�..����;m���&T��c3vH�:�[J6UF���n���z���\��DKs��(��H�ِM�廒�œ�+��-�Y��mK m,9��+N�jyK�s�St�������Y���ڐ3��PW��DG�2���*1����pF�����>\������1��S���^��O9�[؄���Gv[Ԣ�J(Yq���ϼ�%]��a��8kÆį���G��mO.�Ч����u�J,[��:��T����|n�Le�{e�\d�0!��@_�w�$z �ƻ���}Ń[gf��1/�fu�?)���˺��T��(TR�;����ގhv7�}[8� �^�_�t{����P��K��v��a�$�����Xs��J�g��J�HY,�"�g�������=�
(bS��q�v��v��Y嚥0��j���IZ��L� �ܦ�`��.b@E�v��L�cn�ngBeT
��9Mu��$��}�7_X��7��>�!�I&4q��O���х���a�oj*7�*�qi��X)pL��0�Jio�V�zB��@UǴ�Q�������F�O��¥���j�����qi�1B0Trul�j���1a�s zc���2���M�.��Y2���7�����n����G&q1[��vgJ
h�A�@��Ƚ�.�U�}�\�݋�&�G��h��eL���~�נz{x
�F��&��%�b�1Ԕ�s�����3���w$ܹ�&��5��s��u��3w���J�wi�SV�P��>5��R��]w��G�(����n���>�T�5�HC��0Svi�a���Xi{v$\2x���n{�ɭ�X��j�>�iz��&���=�̩t7f4�e��UK(�GTF�n���3w`��+֙z�Z�-@C�?�a�%�d�b�/����;[7�(|�r#iTB.X�j(�F�媍�Z�E.�]h�<Xi=��C�J����AgYK6���s�P�:���t�f��*$C��pv��=Ƕ�Ph*]�!U`�A]z�9�u�+ׁ��S2�E{���v����X��L@Խ1j�_������F/قR7�1b4�LӬ�q+��\���Үyy�(�~閏dz���΅F2���:��鍵W~�p�
��A��=��\�Z��N�إ��0�v���}�]H�1̪��p�)���ia�����,h�]օo\JH��=�>��v�3܈�3e�BiL1�<��1#8�}P�.�:<�a'OKڋ�z�f[F���B8�R����"���\(:�����Dk�Z0,���	_�$�{DFFmv����u���73j\��C���7=0��b�p��κ�x��&��]"�4��{�r6��l�ցB4n��O�)ׁ�V4	+Hx�iv�q��J�C�����ˑ��I�5���wVs�#-�0�<d��;���}�}�V���\��<�gf���\γ��(B�*O�=��*_r��e��;f��	�(l���hS�n��μ[Cm~)mC�G��7��M�y���������V��PQ~�Պ-��G�f��_bW�=�̐S^øN�(���T7z�y�D1#	Zx���Jye���
���ֺ�7�wb5"�Rf�g�Utm�AB�Q�"��q��4��ǬwWr3�@q4vQ�p��#�֫d���P�Ɗ���Φ�����wX��3�*��wB��
k��,�fd�Y�!���g�+ʍ�bp��g{�~M���^G]Tޱ���UF�&'O	U7S�A�f�
��{M:6�xU��QXb��0f-/�� Uis��2�'�"��F��V*᭳�9��H�na�/J��'�4�p��lt��Ȟ.��=��F%�#"7�[͋�5���m�w��U���9&�6}I�nBg�L:�ǹ�!Z���X�.�g�\�T3��G;����E{����M	���&f��kD��	/א��{Rc�����Yq�0��E=z����q��␗�FA��*.�T�!Ҹ�KOi������3ݱd[����Yc\�^OS	���ftb�]�lTA�:j�&�]��~ϾϾ̪��|e�zy;�D�*n"�W�,�2�+*�"x�1���:!�j1ߟ�9� ���V�E��n����*� H�%n*���o�P��L�Jua�ʳ2��1'����t�O7݅P٢��5cB�S՜�q�h��@W��p	�󓇂�YU!�U���7*kq�3�	�[�5���\�e�W�=��p�pT���N�Tq6����{Wڷ�-	����k��=�?���_P��p��f���BKv&s,�٭W;c�GoEz�Z�_<ʗ�=�7��y{J�wm�`��BƺU"��Q�.N*�滅�K��u�tKݭ]?
��k��]��R;��y��i\M˨L�S��u�̸u�E#�V��,}�@X@jYrjeP`���xxĩ�9�e3�t)=�0}��C3"X������3M'[�����_m��M����g�0���n���/����3�cօ�d33^�����!5��x��[���ϗF�ã$�D��#30�eFe����Æ��Ea��b�iOVgl\�"r޳Nn�ArK��,�gO�j�l��%���R�o�;3u�vxNO�/_/=*-�f<'��2��y]ׇ]�IB�7+�1������7�%.&�en���^�eJ�ڸ���~�z=�c�Ɣ��y��(��e���,�
c[U"+�ey�WD���W;>z��a���s�-��f�'�o�oxS�T��6���im0�)a�j�WI� ��$H�5��^�``�'�T��rl��7�՞��亽Qy1���)���`)�&�[�C��|.�	o�;w��x.�^��}��t�x\�y+f��V��p��q��p0b;�;�6&]l:���r/g��NC~�ۧ�
��ٱ>\��q;=-,򨳟
�G<����/z�EMt�9k����q���;��3�_?��Y���r�(J���U���s{+��-x���y8}͋KrߦV_nh��/N(yO��Mt�U�v�d�0!��U 9�`Y;c�֑��"��UY�^����©��GL���;�^+�]�b�Eʲr��T�:؜�w��N{�S>�7v>�6 i	��V;�^B��"r"S�B��c������L0Y�㽭�=Kj���{y(�:S'5�B*\�}#�����!u�F��O�K�����H���sk4�:[��E�^�ޚ���r�:M���-����Hspo�p3p��#���	�<�\���^�%�:z4���ʞ�����78�%H:�t�s�	 h�z�i+�ⴛ9�16�A�_.�����������i/�ۂ�s3�̏	I���y��g�v��[��:����Wq"��e_DMT}���v��kٔ����8b�����;�󄦝�8�w�\.V���-n��ٵk�8\P��p�6��k�u�9�p��.㛡�/9y�}G֚^�G㫋��7��&��e��m-�w)�u����5�٘��CD�Z�J���4v���{9��b�e�[-v:����I�7Eך������p��&�(� �3|�U�8������4�E�:�{Y������-�\�Fa����'����j����?j�We���𼜫�zo��e%��$��hop���Q���I`��7(����>T}O�V|2��C��)�S����ΰ�=��s����]�W�s�\��f�5��3_0�z���s�孊�x��B�چ�����U��~it�ٳ���12�fa<�7�m��g	u�-�]C!�k�XS�vJ}�򮮯�F�s�;�<r;O���A�徺0?`�׏��aWZt,�U����v��5ۖuέ�2�5�w:V|yd�����/Q�a�7�,�=F��]��U}��V��S'^D������O!A�Yq���k���Ϩ�eCx7���:) �F�Z)�nwy�b�	�q���*[I�O������C��/P���F��wYƀJ�v7� �k��})1Q|�,W*�>u_s�f7��X��OX�A���w���`]B;�F�g`%¢�YkGD걛를H|�4�qj����R��F8ɧIX�z�Gs��{]�x�wl��=�<�%r�O)ݼ��F���~��"݉E�z�s��e|7n�ޓ�P�i߫yDk�sk���4���p�7q���&8 ז�k������p1+rw[��Gq&q��l(}^)G`]qW�0����O_u�� ����Ӷ�֭sP��%G*!s5x��`�&��E��}c#9u���	�c���Piu孼fo�^�N}F�����<�}��2m�Fw*Ѵ(M�)C乓����n�'ʸ=�X�"��q<��7 t-QIX�"���W��VmYH�.��쾓�rJ�!]Ǽ�`K�v�f0���K�KN�q��dU��z����s��=�lDա�/3���;ϳ�$:�Ʋ�ӛ�R�ߪܬxNnʹ�3�����&�r���_^Ӧb��+��.��nQ��2�S��ҌR�a�v�c�:��S4�!�a��kyb7�3�'�}�&��~WҘ֘�`Q5�{�Ejc��kʶqSh�1n$��0���=�Y��x���XT<�1:���͞��a##p^��o(-��	W��t4�Gri�V��/&c,p1�5��rh�"���;��3t�;i�z2.� ;|Z��m�*n��`�ٱa�:@;�����r$�Hw@6�]�(��6��7;�7����j��������p��t����$�5�Qo�v������$j�yf�q�d��O��:@�Z�:�y&wo�u+O5����z{_�[y���+���T�Ǐ,,�#�a��2��`t�{6��}���+���"����;9q�݀�GA���ʛ�A�G����lr�6�Y�V�8���Y���%��W����XG�v�G�.���*7�n.�e-��?f��2�1�!��P�R������x�k�F��۝��ˤ����;k����zw��:�'��<�'��	tӹ0�50�*���dQ�mno`�.�È1�����m-�8a�{n�:�v�n�i���� 릒W����u����ڟnɮ.y�D�m�S�UxNf�|7�;|���1��������w9�FU��]�t���{��/��p��У�K�7��^+Sr����i��"���ϵ�WD��	�9g w_bXj[!�kbUӴج�KX�{d2'D�Hud:�� ���׻ W|2���z|78F�uܑ��\C`�7���\I�d�{�����"��ń�^��5|�Έ��[�+8�5J@�2�R���:�
�l�k���Ɵ;7W��w�<�R���d	�-k@�\��6A��輟�#-��+�@�%/Z�W�L�9�;0�zh7OGf�i�O���i=����\�1�Wu�%O��-�%{��w�D*��W���"H�}O3�\����f�6�xٝ�K����^��5��oG=K�SiR�p�.�suN������08Q�ۂU�x�e~��稌������:x�ww$�-�k�VcΣ�k9��E�U� �]9vJ�e�x(E�u��M���Z�@�Q9v�Y�U���6�J5�9��0�sJ��G+$v�[R����m�}���l��+��ۅ�mZ1s�k�&xN.ݙ�7�5���y5Zg}�_,݂���	t��*;�n孄j�m,}�wR�����I Y�ͥA��}}ն�Y-ۘ��}M�uwV��x�\t�L|��N#0����,��sۃ&�7�=�6˾ż��9��7��hy�nn�;�2�D��J1T+��WD*�]ܼ�b�$��2��ݫ���xw\�2V��֑��ڠ�p�*�FjZ���EY����Na:D�$DĴ���TCS'Gg��\�''qwB=4'S�<�QT!�<���yQ����q\��Ш��2ԑ!tBp�<<�e�$TsR0�5Y�u3sKN�C%r��R\ΪNxz%$eh�*�4�S����%����4�lԶn�7p�qܶ�Ur:���Ri���V�U�
�h;��&�����J���p/4��V��I��<H�ӮI��#�$	Jr!��:y�XK��C�kwJ��L�
����qB�l�X�Z�	+�QDxG�Nh��Uwp�箔Uy�T�*�*K�DEU�H��9T���y9p� �EJD��*�I�B�_p����;�[W.��W:��8���ֻ�]AW)�ۍQ�G�F�W{����P�ĬC��i=��Wsk�NU�}_}_UQ�.pN>J����e�����Y�u�ᾅ�(�+(ȹ,3�s����vǾ��v��t^�g�g���r�����:-���+b7^�0�|���M.�G^R�������Kca=\/�nל��*�α�jl��U����n8������8���c�^���)�Q�yOs�{�y6��\�&^##�p�<��mKs}J��g.�:�97�9n
��0\���}��R�v���;{���*V�Q|��L'*2��9ȃ�7׋���a��&ksk��]���|�ʄσ����=j��>y�,O�
{�нF9��=���sg�z��;0�B9#x������ln��t�s�nHp�ksw�[٨<�M�����.����M?h ��Ml��'mm�~�ɘ�v;�-0��Q}���GJ��V���^s�J�ys�<�CۃhYt���Z�V�r�o�}� +J��,�@$��pG��;��K�)V�[��P̝�c"�"˲�ouS�ac&��6*�]=��]s:6X�C7���T% m�����lq��y���}���=�)��pBU�q	���uo��] ���D{�:K�4�x7�-�71]0��.�ѩ�kG)�p��R����{�a7}iSG�1�\��olNb��4S����������א�Q���J޿ƍ�q����0V�[�Q��V�3���KN�+`1�.e��
�:��g�������y�m�q9�Cj�
�%v^b� 6���p���iu�Uz��y���>N�:��*��;Me;��	��:�۽PΪU�)劑��7���,�j���to�j�kdwW��-Q\3�ƴj���n�Gj�p5n4__>�186�c�x����S�~�q0��	��m�~j�)�'=���+�ٞmZ�y���WW9�o�n������ƻDUȘ�Q���7�.��]���.�/�E��2�o�WΡ�:7�ϣ��X��W�T�(i�s�=܈W�^n�Om�u �tzt���vU��v�`[e�n����NҜ��'L�5��,UI�خq���<2�V��ߦ�~#�7ģy�#���Q��]�o;OL�ݰ����an�S9��B��N��t����>���Go�i�>ӷ���������]�O%D$��d�Mesޔ��.����{����4��޸v�i�9+~���n1���[���Ukr���=0_q�z[zE�J�Ȩb�j�/���;��N�e&�[��v�{Q
k���ެ��Դ8���L�/v�?\��ӱ-��_5��t�z��Ko"7��8�H�I���\�v��l��b;�%��|�Qk�Z����/���m�1P�a\�Ӊ�p������ld�R�jG�w:0��t�O����M%K'$7�H��2��C�\�ޱ�wW����EؘEoT�>��bV���#�a��*}v���^�r��.���wz���������D�c���PilQ\�d"�� �W-�t��D�	�~z�v"����;C�<��	�1�h鞠7m��aK���]l�e��Z�>�z�jz��u�m4��x��EU��5]�'2�h�W��[��p�+o �w����j�z/W���|g��Zu4�X��:�c�Y#��\Р����-�1a��"�56���e�.�׶T���*��g�nf���p�������3�������8��}Z8h��v�a%�6<�x�'���s&6j̛r}��]{픦6�k֝��83���~~�>ϳ�Hn�rը1�U7�v.�$��~YPq�����1>S�z�j�o_��v<�X���5�'��C��^o��jz�t=��h�G؜.z�ά�깶׫}ӧd-x��l;���c���KpmDu���V��U������Wm_(��ԕQ�1�r��޳����������[�nO`��g��)���&-�dx�ڜ�����CT��kn!�}��Қ��*8�����.��P�����9�Q:�g���K���O�io3�}�j�j{�������_�m+;�=�)1Z�,�������d��ŕ�h�'+���5��N����z����.��8�+i�es���Rj޻���kF�vm2�W5��q���׊��0��J�4cd]k�:��sslr�z�[H������-t[�(��[��ph���2�*R������86vJ���Qv&�BF��˶OtWꞎ� U��>�S[���|k[w�q�#��5W���Ҍ�qx��U���U�h���kk +��d��7��.��~:�;#�J��^�UT`�C$���~���W����u��g}��U}Y�/0N�:���՗�e��K{ťn��5
b)ؐSS��&��ݴ�Ks�	V#rx9{�Q��d#�^I��o��P���/(���ܙ�Q\��7~�˿.�[1X:����q<�7Ezz���oe��)z@i׺�5�r���c��^�����׌���{�i�{^���]�a�6)V�F;����9�����3�;72��y�p�S�6���z/yQ��KmZC��2_v]\;̨�2��ܠ�;�:T��c�n���n�W����]�9��l'��y���ӫpd�K� �i��E�p�+��õQ��oj��W�m�����ܾz��`�ޛ2/�}3�t�RzEp�¨q��=�oi�8�q��Q�rն�nN��G��x�)?u��;[o�w_�L�kҠֵQ|�B�Oe�6��8�Q�91��֝=�"����8z��Fv��+��L�o]�Q�u�v�|T��`� �f���-���6eu���Gzy��bSg8v���S
9�,�������C�ZLj�E.��p���sj�y+ךd�e�W�C.GG�G��OuBO��]��:��0����=ב���='c]zT�b���.��.ëz'+l��O��k/-ۆޣ-�mB������[Q��d^U�y�2v_k�����/pU��h�V�y����?cCj�C�.Η�Wt��I��Jʈ�2�ι.*�s��'���]� �� �������[�@Va��Ό%1]0��@]��>M#P^�d9��R�V�*��C��lv}�^��O�G��^0����b%ne�Ow<��<�]ߝ���q�g3'������7�ҵ�{����_c�xr{e��˼d\u�E�,^U��W�]�4��n�rf[�zʸuP�m׊�F�K�|0v+ 
i��-�\Τk�>�N��Yw�q_�ci)t�1�+��ݤg$ܛ9���z��c��W�3���f��TO���!�+��͆K�6w6���Fk.n*\DD�|NyOY���.ݙ��b�� �ˌ9#4�.���9Jōw�nJyjg�gW
��6cm^Գ������e[|v8�_��^�\�{�-�J��߷�k��'��fwn�&�z�	y���p�S7�Lΰ vy]\�ވ������
���P����]�e�W��v��9��tн��
��m�U��ڵ5��mӝk)c�͗»�t�A�u9���(�k�h�4�)`��%�k���ܿSK�U=&�^�&��ޡ���1s���'j�Jg�}�1ܜ�O6���&u���jl_7}	��.�ߝ���gzT�I8ػk�gj�Y��k\qk�r�ߎ�W�-ci�(�ok��؍{��*n���Ž�#���5"W!^�id��S�{���F�}��LR��Ti�4�2���0g?8s#cUK��
�����OZ%��g���N���iִ�.Y�D[������!%Q.f %½���w�)ww��Mn�l���^=�W`EzN�w����(#��j%5�>	��@]�/�l��Ӛ�9��=}!p_)�ڭ�ޥ�G��w�h����b��@S���}�Tz)9h�691X�����Aú�q����T��"���Τ�;�:#��O1���[LX�F����g��5ż1�C��s�51͈�\���}u;jB�
w���I8��/,�w+/�'}Q6+=�<���Ԝ��L+���uA�����|S�Dz'�'7�ͯ���MuC��acf���V��a1�-��@Ig��涽��g>���E������'C+��p��[��d�{6�0�i&������ve�����3mi�Ůo�=����!Kj���u�4-��۸��]��(�AM8`L>u�7���������'ݝ�Lg��qI������J��ll�w�_��-�/��{Jťw�%b�zuH�Ӊ.���s��㲱B��GyŘy�/��=mmE�qߎ)��;�7��:�H�m�հjy�b��{^���C�Z.ݧ�Ҷ������77'�I�i���^B��q/��!�-lB�[~���x��+]��}��;t�L���D�Տ;��)���<����b}��ڧ*15�S��v�4AQ����gR�}��_�����z|V�P}:�T_%Ki;)�1�*Y�{mQ/t���	�d�V�i�a���̅�N�v�
�i�v:�V���&��2�ʬ��u+������2Iv�B�K���xC����oC�0�9G*G��Uc:﨡#N��]���\���6zf�
�����jľ��X}�q�L�#��Y�}U_VE߆����_흎���+b��y(�L_%�YG��s&�D�2"z�is|�d�&�Y�I����̧�E�����ߏe�iZ�M���WV�'q�8t�횎M+����M:J�#�u'�Wv-���|�ֻ��cy궡5y]�j�q�5�ܕ�<Э�T�\q�N�=Q�L:��C}��^��٭{^\ٗSM-e��u���7.TB��א��t� �BwUD[L\Jܚ���ѷ)2�9�t6��obP�t�(�@�<���윍��cD�k��ڋ˙���>~���V�*8b-jr\>����jYWN��:�
�F�U�+�r�%��Sz�Wܶ�m=ѷ@�j����J�5G����
��a]x������1'2�E{ �W�E<ݕ�T�^6�J���p��1n������} ypZ��w0���KV�5	Uwoy���_����#��Wʗzv�VnQ7:]��eLaS1W�ǎ6@�o	�4[( FN��gdL��ɋ�%ؽ��;5�̥sFg�Ii�\-�����b�����K��I�N��|}_W�P�ޏ'ON��~��v���+���y�u6;��C�l5��둋A0q�����K���u�]��*��1E��qB���y�ɓ|4,���]|�Ԏ�TE�"��qoÍ��'���K�j�����Z�809�@�|0��:}w�����F�����r�5nT&P�lu������I퓷}�i4amw��Ogsa�ѹ<��ݞv��MvMƨ]�;<r5�zTeb�7���K�s�O3:�q�����|�ѥ�_�Cݸ��mE�n��-������x��O��kز��"/�ţ�[ٯG6������y5y��ĕ��5�>՜�e��#��ʢzf>������ܱ)uCo�N�k��Ȝ����3V���z��F��]�ٜO�ʽ�Jc(֩oYu[����5�y
�݉�Q�PV�A�����˹����i��`ӠRn����+�K������U{_�Sfo��#��'fr�b��uz�ʧ���.�'&�C�k_Ѽ�Ǖ��zxr��wb�,HW���p}	5�3jE��T��_d6z?`�s�V�^jKm�K�<J��L%^��yM�����N;�4��d�k�Jޓ���kv�)�_�����v��&����EY���J�9S_|k	$�����!G�N|w/�}����hrĄ�P.%�����7��ې(.%/2�w�ٔͅ��w�ng�N�Gm�H�Y�x^�ɋ}��%�wޗf��{;`���=\�mŋ�OT`t\�Oz�X���²���ݾ!�Q��98�)�5Td�6�+9Rt�U��p낻�_#RV�T�{N�s�\�
����{����}ܩ�"i�ĵ�ٮ�;ͱ+��S�*�n�5���+���+]L�F	 �.�j�ul��*�;.�s��w6^ɽl�r�T-��@9=
�x�+��ƺM2'[}����l��y���|
�vCJ�&(Wss/3���-*{��:�p�뀶����o(�wlm#D;��|����U��v��d�I�f�` �Lޤ���n�]�>T���21�M4�%m�0��}(�5�B^��jXp(N�eo8�O���0���4�'e�Nj�ž���-aᓅc����;tt\�.����Z�6����]ov�@��	m*�����vNZb��V��2��v���T�8x��0�Tk�<V"�J�Kz�%K��|3��IЈkz���Kú�.��d���K7r`���M��P�;Mԍ:���u�+4T6�^�g^�NdC7�7w˦�4M��3����ב~C�_j�%Ǘ{�pPiѽ�4��c�˙�"w��Z���ԝ�*�͑erw"�F��������8�=��Zm�n�Zf�xc_h{�n�8����Sj�lӯ����BY�7yG+;2�|5�m�ǵ1��L�;�̓���\�Z�A��s�ʥ�\���MS����X�n�&�[�\��]>����x;�FpS��p��B��b^���<���L��d�R���S;f�k>I�k��9�[�Sn�K�!f��͊�`��\w#�Ok�զ�{7��3pΞ�^�6A�n\��:�~o��u&�uq���v���v�q�vN�z;��4umuj���uҚ��n�ľ' �����<���;�Ѫ$��b g"�m���Ñ)/�se��J�O����u4;!�G���V��@N��:j�tM<�W%3�8�����U5��T�6��T�ͳk�[]�D*�lH}>�X@�t�j��k��xy5�'��`�Q���;�od|`�=3��0�hzn�룑�۸7������a,ڰäŦ����}��=X�����]~��#��L�K�0���
�1����l3�Z]���%h� m��s���J
 �9LX�c�F�*�vJ��j�JJEY]"2a*Q�	QU誨��wD*�E�a����EI�H[K2���вJ��d����DE�E ��K+\��SQK(�=���E3R��J2���U�/\t�HUIgMf�TH"*K��<�O�iUQ�J��*�2+�DaV\#1U
�"���FZ�d���A����뙔i�!T�E�{��Њ֜��J�f��VK)�Ҽed���ꙭP�Ш��i�EZ*��U���Z�f�Q
�5(��,�|q��>zy�\�,�HTχ��V��*��Qd^�ڨ�E�\����QiE�DT��wD�X��E����qDD*��3L��UR�:��0�TE#@�G�h��:Nuέ���8�)�O�����jf��vU�����Yn�[S���=�8���� ʱVwx��
�.�K*<������*l�S���$h,K�~�	Gl7`Jc����4���R���}/�m��������4�j��E���g&g[P�*��P���f��bt���n�ս]/���i�^-�ܝD'A�5%T7�y�z���Lm�L�z�EE��]��MZ����^{W���P������6fNp�g���m��\�]�Z2�}�սU��ʈ�O��s��ر8�<�y5=�{3!Rۃ���ۗ��T�M<R�m+�����죊1֑әB�˺��h*�:�p�\�]%��毦��ڎ��EXڞsqv�ܨ���p W{�Fx'!ڏ&�C��Ufkv������^*Ƈ��Y�"�B�4u��v��[��s���5J�:��>MnSr�����bUF��u�T	JS���~7�N�����RvS�z[��vᷣ�c%�����B��O���k/��N�3c5��1 8٥l�F[A����b"���D�*+�yS����T�LZo.�����\��ǩ���܈�p�,���G­[�����������ҥ�g�������Dؖ��'��]~�DD��Tn�n@K'��LnӅ225��K�g5��<�+�oQ5�E����}�Qie
�}��)�
� F��Io�.k�_��ܡ�����F�j	k�\^�w_���~�4��(�@��!,�t�@O��I|b�Nrv\־[����,��9�qڎS��w�rq����8�B���J�7VȔL��N�ҩ���Y����ˆ[��B;�ɮ�s���d:���D�8X�t���voJ]y��iu_�'���E�B�cy9��P�9y=ݼ��ym��]���hB`�bV�3������)<���5%��ѳ �|)ձ�%�|FF&r�o���C�����l��R�y��%V����rݾ�cx�f�4�Z7����P|1�ن��V.�}9�Z��}����nMx��Ӧ�m}�6닌]�����p��0��i�
z�t=����f��u�V4(,wF�1�WgQƀ�YG
6.F�\��%�6]?4)e'�y`�Ⱦ}��2�nj^2�`�-��ԞA��Dpf�C)W<�3;d[�d��¯1X�����Gm󑣂��Kr�[aْ+��KFƗ�.�C]*�U�w��F��V�*O�{�ە�T��3���3�	t�=�Z6o��ʈTk�y1-��7{�b����2�i:�<�Yz�ێz��=;����Êi�_Ը����6�C��r��Cw�u�7��0G&��a��z��(kV�v6����*���F-�hIſq�)�3T�P�ū�xt&�S����O����
�0zA�gP��*�%��AO�w9ܨ�1yY\��������O:�+�am�=>;�Q���_$g�b�*M�$��-Ӵu�o+���Y���no�{��oTD���u�ڈY��}�+��>���v[���gc�H��G�z�o���{�}'�yŚ��$��S9�;he��Z�&`v������kU���u�OPy���n�m���Dr�u�_o.O���7�5�V��+�rs����}N��T��6�j��9��:y��O�֬�:��C���Pam1r�3i������x9�7��'��Ҡ˂�1�>�+a��{}i�ǡN�e����z�u���`S�K�A�_�N{vn��AL�-z3�[��{{�
ݱ&������ZYkf���h{j�Z��M��-~������y��fzu[j��߼y�+ubS��4��x:}O�j�(�;����ʋtVj۱۔���Ci���N\t�P�u��J޼�� ���|);�Μ�I�$���_7Н۸jJ��u���X��:�
� ��5��V����C,=�y��E��[EN�_F�Ym�y=h_b{S7`έ�m��ͱ�1]��`�}�<���y�+}K���&Sa<Z:���p8T��?���I��N8���7peB��>�Wg�3j-(\�o{�Ws�V={*�!+-�#r{�RzmN�|ս�n+�{(��kޕ�'򬕵��y8��=v�z�O3�ޏړ�����EW/��Y�5��j��U� 5���]�ިk8�c�}g�9u����4��d�+޵�mz�잍|�� �\��b���C���V�Y%�|�Yq�����w��މS5�6�d H��	�q�J\U��x��w"�m�z��v��JMq�&��@֖��J��Qa^���t^�ڎ�o�yfg$�k�:�y�:��~�7β{;���N�g
BA�Mv!�#Wv���5�M��%I�lJs�����8G�M᡼���猪����]��B߇GmD��@o�_5�GL%���SJ�kʅ�4�b��#�v�٫�f�,?w,�R������s���U!�z���+�G�g%nN�w��7�>�L�"�W��F�6���/�}ZZ�CR������zYǭ��
څ4�J<P���'>��,��\��'SyQ'1�\�n��eM������C}N���U��	�o	[2Q�����쪵�o���w�f!�kC�N����Cz��s�V�|��3tkVvps�q�:�cJ�c�Oj/3j֙�Š�w'^N�h��m����m�^^l�C7We��+�/r��uy����f���w��MI]c�aܻ��i�N��=B����:i�����Ek�||�h�[Q��*z��K����y�<�0���oѿK=ֲ��ͮ���.�?]��s����W��z���T{,�ӞB`�d����i_���K���薯_�T�����(vvhl���3({���zF�ٲ�,�k&��8�8�ƞP8���5�۫�SF��Sw���U�p8Y�"+pwۅh���Us�3K�1�����%u�΋޹��G����v���f~�ģV��D<[���5}5�7�e�AV4�R�k4踩�XҞ�Y�8�8�G;����a�y��{��Ƕ6�n��P6�*o;�O:�ֳ�2���*Ӵ��������k.0�s���)��k"�K�-��I(Z/A�+��J���c3�Y)�OV���ݍ�H����V��j�4��lPX�65�J��
�k.����EPc���>wҹv�UgO7Q�������3��0�pI�T�Ǒw���K��GV�&���-���{�o�M��U��Ɵ��P��?�w/����r�g�z�b��J�MT�8���u�i��8u���n1U��Q�EoOj"�b����bH�����P{����;�U���M�r�js5�u7b0ӹ��W%颷c�_s,8-eA��C#��'�=ބ^T'C+ܝ;C��;N2�U�<u��Ê��y����vϙ�ةZ�iɇ���Oda���F/lu��1{���Q�q�`�`r���.O/�b�ݢ��:��fa&�JJ޵dgI]t7㯟:	m٭�v3�-/o\�woW�w)fEu�d�1��dpw3d�����8�OZ���*M��j�E.���.t\�+[�ژ�g���'���[y}�ޜZ�=�J���Whڪ6�c$�J|����;��� /��u������*�ǵ����8�{F`;��X�^+��Gk��n�߂�u��5zq�z�Ǜ�MM��V��5;�Bs^)��Y��󂮚��\��*̤�hw[�vꏺ�4�T�h<~Ev����ǳ��Z��9��Fsխ����\C{���in�����K+��s����"�.q�ǧbG�gF���w�	���ˠ�jl��5��R��rz6��6�{��3��ql�Tj4���7�e#�B%�Ӎ8ia�R}oiMv[x;�����^��FE�U崟s�KL�aP�����P�GZ@M���r=�5��E*�X(v(��]J>���ٽ}�w�������SV�|^��ޞ0{��W6kڇ4�
	tJ`loE�:@s�w'�y��k���D���V�T6���o��ڢ+*��~����u��z���X@V�c����R�K.J���Fvn�����ShgX}3t4��Q����(Y\��feN�cA��r�T������'�ۣ�&B�/zfr#��ﾷ;�����Ƴ���{�NsM���s^�ҽl.ys*��Ś1Ѫ�*Q/�]ىT.���[2����O�/W[y�^8�P�v^BÝ���ou�C�a��v���Z��fw��w�;��6��L�7������n+^�����r�P�.���^sX��H�49�s0rg�d;�����<�l�舘���>
���2ި4���u<+����=�;��}��t�Nz���w;~LL�6������`O���+]]*vVT{�gh\�٥G��w��5 �W����������+���n��b�X�b�ʽoۋ����s����<R���^�l��6Z���Y��S{'�7{�/p�7ޓ�]�z��-�O�lO]ƨ�Qz�c�����+؞���i�jRc�=���UD^lj��6�����wQ_9�b��gݾyZ��]\H�E��������=~�uu�-���o�Ϯ��hn��b7h�|Ͻ���fA!7B�tf��d,w-;��da|�Ѫ�FB2!.:UF�C�WS[L5if�pt��:Yc��+�Á����ݲ������g�P7/����s�?9rQ7��lO*3{I�⯘��՚�k��j5oMȻj0��;�+�z�=��y�͇�;� ���jz��K3=yt�};M�������a9}������oj�[�ً� ��,9��\�b�o�n8��2�
�j�(��Ek/�ck7��Uѡ��7G�ﱾս����lj�s	p�j������l����F��f��̫uHΨ���;�P��D�x�}ws���Ӌ:e��*�L�+u;�`�Z7������]#H�U�נ�S]0��ُ#���٫�����ƻ�ݭ\�j5�v���E�1	oQ�냫�kps��pF���{"~�9���zJ:�e�6���eC��Q�Lh	u�����67��暥\�l���a�ׯ���N�rfvP��Uï@T��b&6�c2˻u�Nu�܋%��6�U`*}Q�.��svΩ� �yJ�,�~���b��ȷ7q��ɂ���1-��h��)����^u=ӄu8{sy�확����AIq���M�lV37
���*�V�ԌWͨ�~�;pL����,탬
�-{ܶ;������]��7��K��e-�9;�Aב��3���dT��[}+��gn�����eU=�R�+�?K�������L�۠�j�c�Iۘ�@#�tl�s����ektWeWQoUz�s�=4��n�u����x���@l?s��1>|:ֵ�ԨVv�����vrq��{}s+�5�{��L���|�ۅ�6��*b��7��t�C�Qc3Gy+ݙ��c��?,�{�Ǿ��aU���7��بkC�����-�=���fubU��Zy��=�Y^��k�i���r�:�^��O�<��vԱ��;�m:Q� �K�t>������D�3��E�T��i�^��:V�cn��p�C�X]B)c��V���+СL��Ҡ�R�Q|�-���x���wݧ�frv�J��ݼq��7l��%C�G����;�r�q6�Е�H�C��O݂��	[�d`�����<r�j�K���%�a�b�׃����ȥ��ܴw6�ۑA-$�`5�Y�fͺ�<�gp��d� �u�ȑ}�(�{u��������l���h'T ����a�I<�e�*R���m�ܑ-���:[�b5�A�
)!.e���J��#1݃��3v���ZqT"y�e��;Inn����%	��I@M閯$�O�ʤ �>�j�rl5�����1	��؞�]����D�
.T*S��������a����Y��s��&�e����4S�pk�ˮh $��ҡ�y��r���Њm�y�sE��7r�t��ްJ�O��	o�����R�b���#���ot�0gp��Ѳ��C7�~]"=FT{�K<�w�=���>��jp=a^�F����V�[I3:��)��d�{y��:xw	��E�"��fɇ*36uf�($��H���b�~�� z�����Mo�X�څ�� 8(Γ9��F���ݳǾX�B!�����8YP}�]��Xf�yv�i5�"J�>��B�z��*�`5��7�dhI����%�盧�;�� `@Z����r�rzŎ�-��\�{��Hx�*#��tY$sI�`taV��Ac[͇ǹ#V�[wb w�>�w% J�����%���i���2�+j!�8�Q��j��#�
�7D⠃�T���c�(��
��ȍ���H���
�
��aw��_3*��ϻ=P1b�4 Ć|7o����]ZS�τ���$�ͫ�e����L����ᷚ��- 1e��c�n��|�C�;��z�v�}���S���j%ZÛ#t����]֨�P0�������RY�����1�p��`���,�$���DB���E㊻��?��R�+�̰=K�,��Eт�__<z*v��
�-p�灖�	�X���p��q�m"��(�=w��b�;���R�u�,�v���vL�BM�+Zܔ��y�(���� viO�v>�m�{���)�/(y�dU�G���gSnl���>���~Z�`״�tF�&ZO�η���/�r�j^�:�Ҿ<&n�Q������Z�:ګ���!�0t;Vm�����FXsׇ�85?5Ǫ{��T�F�-��w�"�;fL<\�gk{�!�j�9ٌ���`�.O_�G������K�3Ջr�X}%��8G��� ����a����55mn�1F�-6J��_	|��ӫ���a,
-橖2P>D�+���n����Z,�x���Rp݆T*ѣ��ms�z���ab>Ĳ���\� � ��Z���?d�&:6�+ޜΌ����A0�H777�)�5�����l�nt��[��_E@&����i}ݨ1�pA���Īv]t�쇻I��8�Q�4U��]yJ�,sY��s )QA�(�L+$W�s�XE2���#�(r*�e�U�#��;��k.Rn���\��!R�F�U�(�5�#�)ʊ�I2(�������$��D�t�P�D�+t,U�fj�C$ӭ4�#Ej���HE��`W�)!�I&Օ�hF�I�(�*ē-�&e%G�W�i�x9F*�2�	GZ��ES�mUf!\ң�e�Т)��W�w3dQ�㬼��a�c��eV�R)F��&Es-9L�d%"���J�T.�TR���O������㮲��"4SMDM�x�iz�%E|x�ǆ�U<:p������Rq�"�r�1B̠�
$����UDR��Y"���K��T�jJ<\�B�����q[���W�P �A 7��f���ҕ�l΃X=�l8�к<۫u�gW�傫�:a�,�4C|�%�jYyw|~J�w��EIYQ�X���Xʰ@��-ݻ[}9߽�:c�%6_u7�8��HmW�<�wz�[�=��D�kz5ˤk/we�-Wp7��;[�i�>�u���n�"�&�.�w��o�J���
}׮Mf����{^\qku����s�M@�f�Q��Y��+�ciE臸4O��%nz��]���$^W*Q���&�9Qqf�n�U-�`���^/��h���o=��4�����w��~F��Ѹ�/0�Xw��}�]s�a�p���p�2�l��K���8�i�m���d>u�����j�ŭ��������wN����p������6�1%I���Ӽތ����Kt��^5��9���nţ\�o��S��Mk�e���4��M��Vݜ{�*;\kΗ���Wk�k6!���;�r�fFr�����<�~vT���}s����֮u�[����5[�v(I�6́�)*�M��jK�ӆE9%1���2�Jc���|k���v�ڰ�w��݆U�"�e�V��^[�2����WVm<���x���Nҭ�=9��{M�[h��_���A����b�n֛�c���:��9S�'g;�{x{���N�4K���+�nF<m��7���8�q�
�In_"2&���8���K�RjkU�����x.㒠�N�|��D�&1􈐖>Z���γ�������uy��S\��9�u	�O��t8�eo���$�L�����Tr|���6��[Py:�a+���Ω��0�t�7����Q��&c�w�E���h�W�5�W�;U�8ɧIF�(
z��4{�'�ݭFY^Վ �U�9�p\���7ڎtC���Щkt�P�Fj�.]��f����2��_�p�j���.���Biu_j�1c�E�sp�i�G��Y;z�6���[�)�oa��LJܚ�O�����:�RV�j��p�b���N������B�@Lp��W�-�^�!��.�f����{������כ����mC�*�҇@���=����\w���`ҥ�Zt[�úg8bF�n��T������$dA�h�V#C���C�Q&�d;���3�n#��#JW duڄ>�"��u�v{�8�h���F�3֍���'�ה׮����S�}�[)j��$��'��oCϷ=\׷�x%��v�\���Z��!9�z�3æ��e�Ş�$��E��/M�){j�ťw�mՕݾ��.�jz�>��*4�����.q��䕭�mh�[T����Q�9¹lu�*	���j�69�w���ݸ�k٢�#�fQV��Tqq��R���'��q]b�v�{�'�|��S�{�/3nQ7�8����ji�}Y]��g���;cB;o�4�T<��!��t�[��;� ���\�U�ɵT�R���C�_m���w:x�m>�oQ��Ձp�5L�^��ji��3(�Pt����9��;�`�'�㔷��Żm��$T����{��q�w.�����2�W�e��V�'�&m��W&cck��s�9������r��Y�n�;�OL���p;�Z93�J�l�{�n����Б�=�� �K�����:����.�Ý����R�̠�/����{0i�I*�+��@Vi���v��b֫�6x��h���;��9r��>������M�|Ӭ7����8�r#��9�N�i���\����<];�}~�6���������F�����􎒣��oD˞�M-�S�ɟw�9�ƭގ����<+�oQ���bQ�.9�]�"UaʜI*;;o3�ܮL�7�����p��P�ላM��FLS���7��s+b�~~��g���O*����|o9���qyQiS�t��P�u��ѥז�-阼Zr|�MIW�c*�gl��rJ�&�5�]n��ã�Ч����y�bQ}N��N��Q2i���\'q�o��j�и�R�i��^xc�=�/���c#�tr��M�ܮ/B�lo��������٤���Ҿ� ���ta�a�`s�ܼ�]OH3Ժ�����9=�1�o��q��V��m.*�y�>ۓb��;���.of�:���q�Yɰ�c�W�Q�盋��=}K*ht7�0�)Q@�6�af�Y���T��s�J/V �QHqҐ2jX�R��0F�Y��E�`n�'s}eɽ
ޭ���o6��:���S �sv]Q���x�����><8_Dh����94�Þ���E�ԩ��ňl���v��]�E��N���U�XډqZ�O�{l��R�0���5�1�V�u�X�̺Ėr���k���-���Z�R���1|�,�����ա���vb��<ꕈ�q��n{P��\q����L���R��\/��*^Ѕ=�Ne��;��6�T��/���eE�Qә�+��7�J�\�f+c��`k��b�굚�T�ڻ/�GL+�R����/}N��Q��f�Ү�����)C!�:��k2��~���N��C�M3��Ji����;7qX1�`]����<�[ڈ0��W���kw!��&���v�+n�q��a븑YA`Ľ'N8�\����}^뗔9��^�J������r���y*��z�t����>p�ٗ�r$�u���u�;x��
v��n���:�v�'�-����P���v��u���ڢ�V�3ϙ���������+�����Q��_A0�ʋ>xM�wn"�1VǇͳ{@�1��6nn��웭v�L_��C�E��~w�̘F�nq��>��:M�z�o6О�xn��"]�����=te���8�x�#_T�ٱ��q/�)����;�T뜄��k�z���K,����}S��:W۸_cک}��V-*t�:����{ϥ��Y^e�׹Z�PF����\��\��QY����ͬ��E�u�}�1��Ka�`^��T��5dMc���iN�j�eo�%\���b�ZQ�m���D�����(j����v�9�k��c��U��Nnom��ά[�9���۞�s���b}���q�p��.�ݐ;J�5�+��y�ȋþ�������s�yA�_�tiO1��Nޣ<�PY�5�uJxms��P���.��~�����-��<��Tr|�8��-ۈƣi�ut%�T�5A��e��ٓ�]=W*=Ǚ~��=�G�ߚ������7
�WD�Ѻr�#�s:�`<Sp����,�pXs;�A���f>��\�kJ%4^�Sɴ�������q�Zpb�4:��� g/`�`7P�G���jZx!�kV�Wؐ�u4=XV, ��N�F����]6���5�+,�y7�.�Bh±�`��k"W$���33��Ɏl���'�������뵬ii�
|ِs��e<�*oV��p���kmn�.�V�dB(�����9��}�O���H�{D+��oo�y=�ǲt���
z��p�o![���oT[4��[��V�w=j\78���:��w+�;KeB�O�
���	�� ���ii�w2T9��c}<��~�5��oO7ݡ(��nג�^��	�C��n7��SZ��MYՋV{�U�8�fo�]��'v�+�I�o)��F�rGem�Z�-@B\.
���8�E�*���@�L�PR����kB�1y0Ԗ�6U��w+������T����o�C��iX�����}J��af{\}����v�\�D��fo��ZߪKj�C�r�.���5�H�!C��76���&<��u6�y�{�~�������~�lOW%��[k��EJ�~��زx�}�����{���j9��}�� pX��Y�+b����J\ ��[I��0΃�(,Y{}�@�3Li�w�e$�v��9�l���G���j�Ո���/<��!>�R/=�u�/�rTߧ^�_eE�������j>�l�S��$��L]�u]�s�󆨶�Q����X;�+�:gw6�s�m։q7ԵT_7^[I�N�k>MvE71J�x� $�O	�Ǳ�A\�$�R��z�σ�6��������ך|�Y�`��;aI�V��o�<Ԃ~�O=+����*���ꗒ��z��w+{*��Vڇj%Ӝ�c��r��0��nל�^�Ѝ�D�xߠs�ή9�VS�W�"���]Rn�b�Ѯ+���K����q�N���Ht�\�.U�3+ϝf9~߁��mq�*u������u��8u�����2�|�<�<���*�4?b�x���Ѳy���Ց��,�2׹3��S��3pU�T7`[SNi�~�y�8^��e����E�N�=�=�_b/5:�LL�}�ٝ�skne0�N�ki�2��.u��׍.���oN�/�^�M9B�:5�+��cK����u;����ua[��9έ.+ȯ;�{k�^�V9�L�.���Rmk��gn��8�*�k*fܺ��!�l�S��)��{GX$z�ג������":��J�
۹��[��cw�ci�+e��/q"Zt&��a���ެ!^��K�5��h�+{��3�M�<mAC���b<$�i�7*ծ����V+�����U5�i�޺�\t��w��OjrT�#naCњ�f����~�Qo�g��_�ˈ{{4����E[[�C��pb��BM�Sec�]Uc��6���P��w�Ux����7�y�����?p�W�7�vE�;��:�^����x�b�����.��X��B4�ٔ��o��+�Mɣ��K���:���[ޟ��Ϻ�1��A�y�f�6�_]qBi[����Z�w�� ����^���E�U唙W��R�k	�#�prk�#s��]����w��am�B����R��R�ʃ�54;6��:Ğ�yՕ���:}޻�ZW���8Ɉn��Au�	.7*���O�p�z�|��-�겝�s˝���wOw�/8��t�B<S{�\��Mj���Īk��[3�ˮ]lv���>tğ�W���쿛��*��k43�j2�?o�=�Y��YR�`M�� ��� ��m�'7#~X����K�i� �'���{jpY�Ρ7o�f�pA������f^�d�x�*�Ns���*k��i�n�˭�
V��շܸ��}a�N+j�U�J���v��UC�w߁�q,���G:�$p���p�v��DN�P�O��T����L7v��3۸�|�`/�L��Z_�� ��L�Q���c>MVѿ.��K|�|49�.�in����l�^p7���W�U�
��%Q�!���Z^�QPxl�̕��=F�wWQ��JjG>��S���;��X��|s��8�3��N�+Jܪ�8Ms����h�;�=��o=��.����o�{��e�����y�9��I�G����`<�������m�,��Fb���;d�]ۿ����H�{���	���b���ݏ�"<�;Ppt�4�v
���z,��ۙ�zqf����х��?D���Nӌ�����gyLG�m8�[M���ZM�`^��E}�|���[#�����p�G\_�	�7~��Ȫ������ک�� bкݑ�5>yo-�n�l�i�tE*%��+�ݱ�A\|��Ep�%)�,aٿ��u�v���C���
p}�y~��]��b��ڡ�ʻŀ�S=�yn6Ҭ���Z@+`���Kz!���:1�yr�Y�@i��u���\���KYRQ��gC�.gGש�Me�^�A��z�:�|wf���.(��g�h�-�U���Zn@�].j��TC��^���OT�׍��n[���_��Ҝ�D�,�p5<g�!<O��b�gƷc��T�tBm6/q��B>D#jsF���(oY}�ŜWe:�*����C�J�|7#�ևMov�Y�Y繵�u:�)�zP6�i+��pF���%zXkK�D�i���c�_N=��@d9���ӵ�_A�4ʠ���JGlFo�2���]�bX�&Y���1$te�tuPYNɃ%m>ӔJ:b����4����v����R��
�+��ٶ�U��v>��J�Q��/w��xr�X���gi��;>O3cW{3�l�\��5�y>�(bY��i�E��o70dE;�.��*��t��"�\Y�L��{[��N��)0�8�5ӝ���8��e.o���L�x#}-ŏ�Щ�h��WW��>��N����X�:F��(fKn�b�,2�����lŷ��ۆ��=����h��=��1:o$us���E��N���6�L^�ӆ�xIt�-Vq^0(�tSu�f�u���j�\˹ȱ!�l���<|{�7�8\��4���v���㯯��w�n��h,��ނl&��;C��m֥L�޵�N����\�,b̔Z�᥀[�{M��{κjb�= 6Y�)[d�U�1��S���2�vo	�7���.�Ҭ�J����w�W���wrc�>l�����$�댈�q�5�vp�f�e�tfݳw/�k����B�X��PHO^J��e��[;��P:έ՚�㵖Eu�^.%��im���/���}�V��z��ǛL���Pڊenգ ��6[p��ԜY��:����}λNpsWP��Y���F����ٛ��~4v�f{8Ï`>P�����8���[���_h$�������I]�v�k/�;�i)��͊˔X�*o0�8N
�P"H�M�X�.z���B�7�Rr�{+��n�/�՞(p+I�S�Ӑ.oQ�&���C���-\��3cb��Щ�:�-�N�v.�t]u�<�ǹ��.<�N[:a;�kt���,�
�{e�1��!X� `12[WӍ���浓'U�[3\*����������Is�!���ަ;�뽬2A��E*T�k�=���Hj�$.c���W�o�� *�;�%�H�}1;�.7Ǿ1��k�{l�D-[��h��s$�l�L��_]���<�9��W�쾋w	Ž�h ��W�nN��[�GKͬ���TY�0��]��1,�
�Ku�|v��2X��.��B�C��],o�={�tu%�3��)S�D����6�)5ҷ��f��Q����6t���e�7oה��9-%��9�~���D��φ2���+��[꙯�|�T�e�EkQ ��K���T�Iiu2���.V��L��$"���B<Ȋ##H��4KAbg(�j")eJ"VH���)u��;F���
�¨���KRE*����GCZ�xy�]3���*dQȩ�u��KR�LԠ�#6&KP�x�<��TO\��D"!1=���Rb&���5�$�UTYFr�����<7A9t�bbu(���K�DG �f�ܪ�­*���3�*��Q3�UUR�S������hQ2"�2��I� �J!ά��93�-k
�H墨�)lа�f���W��f&�`r���U��E%�R2�(�a!r-K�Fb��
�E��µr@�6�**��,�*,�K$�R�g+�EtT*"�2K�:M2Ȯ�j�ԁP����.sD�j��.QFB��U2C5Z�DW"�$�"�W�UUW
��*��|0�}u�Ǟ�3qs�HιvW:��?'��COr�ٕ�S�*r��C� $������W�C|�w3/���ea��T��i��rJP��w�T�ì�]�,�}A������=�ۘ��gZ��5��� \X�����3���ؒ�Lߪ�Ml�&�P���2W�3�s�n���:���t���*WTw����fY>g�C ��h��j�SJG���\/`[f:��΋��5J<�֥|�+�&\�>��-q�^��ͳC�@=�ؑ!*]DQ�]�>%qy�m�W��6h��D���]�s�k����'>�?y-��y����}�C,�|�&@_�&'���ӑ�Z;��d��$<��m	;��]�J�^c���U�d���9=��Q�c�0�<O��Q�lH*6��1b�5S�F2�.��[>����B���RǊ�q̯&hm��l�j�����Y&��T���Â�5A�{fk$�D����E0;�aU��ڶ�J\m�ݛ����7����9T�h�~����T:�ioξ�u���z���g茝I��v���L}P����5G�C�3:vcE�sA�5j�ܡ*�;�@ܣ�/�!+�$�v�jו�X�3�}���f��E ��q�"L�e�kq��o}����h�i�l��v*@S��	�:�}א���� �Ԝ����hԮS���������Hl��9Y�C��9Q<�x�s�M���=�u������a���ܰ:R:q�Z@�������G��*�v,Sοt����L%t	��
z�Dh�J _s'���D4�0]�������&pf��y��6�j��`��@w�+����TХZ4C�{���|�%}l����,����q��t-���p�O��L��ӂ����Kz�-/͍4�srѺ亩-?l��;(��5��vC��n>�ߏv��7��|3�Q�%.U���%�����Oݝ�ؗ?��,�d'���W#�uUǳ��z_�x����'�G���h;����س�S|�O����f9*
�����EŁ�)�[t��ҝ�<�x�Gџ6��O�KӬ*���	�p��n��$_B��+W(�쁮�R����ɿ��<���C��>.0OSY謧u
�uz�h��Q�ؾ�T�0;iF�to�9
�#
gI؍�tE R�&��+����	�{ەUa�u/w����u�1ݴ���OF�Ddkv��T� %/�fCf�Ш����f-���vq�<ݻϳ�'W��Ȗ{Q�����6�^�G���E]*�D���
�f���s��w��z��ՙ��P�7�xޞ%�ɥblK�L�7���ߪ!XǖC%�D��|��.G�w�]mp���#<-�7���g�C����%�o;��p�k>�3=��/G�"�1��vq/h]c��m1|_{Z���wP���פ�p�S�v1�"��}d#�{R�G��ً��{Ka��N+�\����qi>Ͷ�`���
� �K;�9�O�u�"\z�t�G|r<6]=;�����'*�G5)̹s����tz��w���ޅ���,#��hI�*���,��I�S��D�ƝY>���5p��lu�_�����D�OlV�[�~������]1C�N�+K�7Au�{�#��N#����c�[��57]T���y�Y����Wt�|ۣiUC�dQ�2Q�	���9��z��K��0�.�P�Q�Y׵���߲ɛ��T鏾uR�9�\5�˺�z��듧,L���Q����L�������c�ٜ,���}��Hyc%3�%+���/�\KRl��#t���+)��p#L\�����ۧ��Ule�׋���l��y�.u��p_���������ٳ����M���յ|#����K�NAٗ��Qd�=>Uа	�y��)l��󩳫a�Da �˻~}�cZ���z��X̉�&��T�}�1q�:������S����$@��������u^��/��ﲾ~�WhhϾ���ȍ�*H�%;P���W�8;�ʤ6/�܍�m�#.�su���v�KZ����V�s��L�b&9�]�]�bd]I�����y��Z޻->vI��	�;{[�G��f�Hw{�7XS"�v��𽫇i��� �tk0Z�Z�#�YD�Wn�;+��u|Մ`����/K�oq§vneww�}hV�����]?���ݸطV���UA��!��t�n������l����u����9����,d�=�{`�-=��"�#�y�#�py��Sv��(�WDG;7v��T�Y%���|�|�M̏�vZ&�'�;�}D*x�E[�}�6�W2��ƭڹ���$/�����>�J���K�_]E.;zUw��c��R\��Ls��V�j�K͊�S;}d�W�W��0λ�>��~4��%i�#��$M-��t�Zw��ǹKGc�~�G����.����y��w)�8'��!c�Ȉ��z	+OxM�Zlc�j����=����J��騪���䔧A�خ|g��/��
l1�~�DRrx���;��vnT$�ÒZ9��s��y幒ǲR*�5/M�f�XUJ6U��uA�rI�rx��2�|s<\����t��7�ږ��4�֯�R����ߺl{eq2o6T;o}���sĭ>�M��xQ«{~}��.�%�~��߿N�������~y��~�d�7��_���L��� ��;@��a��_A����z.WyU�IM8ek��ҍ�^���D�[k6K>�͑LaG��e>����d/KT��>�����h��{%���v�R���h�ur4��	�&�\��i:B}j%�n�Q��f��`�XϏ+�v�@����-��	Rir�������j�{�W��gL[b{M����c/&����֝d��_ÒU�ď���FE��Np�s=��d�	�k'�T�_*C���q~X't�D���P��ez�_�3�o��.�4�+>x�5�9�!����d�~T�w�/cl��60G�E!q�%)�,a鸊,}X������ ���W|��}�{7;+n��zꇯ��ӯ�3���#�I�[����1�(g��0���{izo�������@�6b.��g��am�g%>���.��9�R;�O�mիc�yָ�JE���a_I��Ov�ʾl� n�U�i����A�k�S}���'��#S�7����=�n2�T�>�u��չۑ�b�ft�0Al�����p��'�<O��P�_
��غx}��Ϋ�Y
�am)[b=���Z��Fh��c�]�"BT.����:�8J���m���^��~�n�����n��?�^�G���
�Q	��c�2��_H�H����'gIo�5�//M����>��C���lp���������DB��,���$��>�TnS��V�+D�{�a>瓦EZ�󼙻�y{�-���.�XNJ7{{N�7�J�����͓���a���f��A��7{��;�i�>���ym2�ZB�h4����*E���j��A����E5�{LV��ɫ��7�:`���e�L��w(a���.z��>A�nﺷ{=�3Z�mM����H�;��I��o�ه��/��I'�Oj��"NQ��b'w���1��7J6��Q����1_v��R�~<�C��sr/�ڨ}%]P~�wva��^���o�!Ld�8�+�%�v�(������rw<�`���<�\8����F�#�� E�]_ɤ��?B���Z.s\G1+�Ih�>���{�E��׍��T��m(���z-�������%V��v}c��_"S�3��]�E��F�w'd�>�>���Ǵ�{�*�C�y��y�?5k?]�]�w|�v���̣+����P�}��\,��ne��L�.4|��4}�/76[���U��ǘ�vlO�Dy�.wcp-vɰ�;�����F�x���$�vH�?na������o������? k�cj1Յ~ɝr�}3��Uq����������wM|9�cP��ꣽ�>�;~������N��R�����uS�纥��"_�a��G|ڧ�:��f+e�����u
5���Y�0���c���Q��g�N�F�J"��d�rR���ö��pS�y�6:����U��$�Y����[�gY��nS��.
<ۻ�[fq�D�u�Akx��s+[��7�[�u��eՒ�甹�������bQ�P�jc�	���w*�F*R��v[7�s���ᯝ>;�
���g���'q��9\�t7Y�B����7��n�OeU�!�K�&$c�n��+N��#ܭ�qc�aX�
aT�'b7�M:"�)W`a�W��;����^L�}>�O�z5������	�F���n�k�4W����(�$.�BR�fCf�M��Y���e����^u;��6��?@'��Ƕ;�U�w�p7��Q�1>�:��ry����@2P�o>��8�}��c�UE|T�9�Aq�������o�κ���ż��n��J�;����l+�����F?I�X����H�
��ĊS�>��T��Fv=ɚߛ��#~��U'��R�F�w*���K��}��9�s	4D�4����o)����WI�s���D3?�N�B�8�=�����#�҉���r�=?|��;��LJ�r_�n���V釟OI�s��۬���ՍT� �>��4ſ�����u#��=� �I�IG	c�N�/�nL;�g��so�)���Zin}�����L�Χ�j0J�YG�r��o��wQkdᡮO��a}����hܣW�e��U���w�s��'��;e3�p{��W���':����{{B����	��?=�&��7wY�f�eӕ�6œ��8�ɋ�ftG�Ͻt��D`�9R����3G*.幌嘞�J��og���n^p��Z�!Gz�-u��N�"}�N�ֺI�zi�f7Ț�����:ԇ��۴�Q�;(k����S���O,fJ���M�M�4�a�v�ͱ�3���x\c�,V�V=�F�V�q�Ѱu�ϧ�/��5��e��M�G�$�������j��3�b��nW����;��`��!�{&��~��߉�(3�U�*l��cιK��e��{�%|t��2��F��y���(�X)��/��/&u��+n�9:����/�k�[9��C�}oO�֩��\>�gC�<TvzvO������r����Iܡn�QS�V��܇٥zϟ�6�>8%>��.��1*7[��U}j0t�w�F��k�t��u�ꅩ�}�ӹ8�"�g�s'��zG��i퇟'I��eq����.\i�(��a�7�������q����h�T���G��������T��j�����G��g�]�q�������F�c���
Y,T<�	e�Q���⧰�wu ���.�9�����3�u�7����7����@ՕQc�iC�ba~�]"bb�W�qO��s���9�VՍ�l����C��g�I��.�#�7�b"���4&V���M�q"E.�QJ�S��͇�<�{L�z=�Ƕ���Ng̈́0�}��R�z��S��K'���:й�hՓ|��s݉ԘũPU���Z�����6=e�ٸXs���u�:� �0�VQ��ù�lx8WP*_�k��WG<ƚQ���+Й�X/�!�*�Ywb�I�k���Q��Nz��Ww������p��]&�e���Cs���4�ڪ�l6�!�ϥe�y�,�Ms��1ǢU�n��T�\��XXs���W�^O����fo��L�o2���vT�>ǋj�;�l�
�G60,;Q���B9�/��̿�*=s�q�2<]���_�{\��7�L
���| k��x����~�C�c>_�����2Vֿ-W���`�I����2�&��q�Mi\��{U�;2�8|�y�����ժqh��d��k���:�닅�wM�x~S0��V�N�\|��5��N��Qwu�.
X�J��y�&ו8��Y{a������c2Ot�Qgg�QP�@Vr��'��wn���5�`�]�d��y;\~��=�>��p��p��'QY J��&/��&d�浻S�����;L��>�j�E��eE��I�ɫ�]�g�Zq�7�}n1�~�F���9�o�><��񨞐9L���/�n#%��۩	?�����
wH���Mh�:FJ�S�\j��iԺ؅*��d��گxJ^|�pp��մ��(��+wT<�섑�id���|Sv��Hn��w����9�v8��`�E�[ըc��K�[�{�
[|�٤:�"WV�E&9]���v���W�;�H��̈́�6Cn���7����aՖ^�x�(���#@��g�9�Q7��u������(i�����1�TT��ͩ�霷�}>��w�2��pƛF����ba��T`'=g���ƫ/��G��}�۩�gz��s�֢�Ľ��~�����<��yFy�H
�D��;hL�}-S����v�^�����۫/�3��<�u�ϕ5yg^�9	�����ʅ��%�W�������֚����B��c!Sվ����{������3Cl7�l�j������Y'��}��4��wWr.���m�n��͢����\뾩�Μvw7�ʑ�:���ˇ��-@ܵU5�ghc�1�ű8M2��6$�.����dG�{5�6��������\����|�}�;uF��tG>�;j�M��x!e"����J���	������7��l�ح�Rh���o6~s���盎��%�Bo��.<�'"��䷂���c����myNCew*]Pi�|}�Qs��˞7�1���DP�퓁9�Q�֍u�P{�pu����B�E�
�6�6�e�>�=

�X��)�b�$�A0��5�wf�)�;�ϭtT�y- ��A�cλ�0m�;�}�V�U�a�ە[Xv�j�����2x�&p��L��E�#;F���{k�άF�t hE���n�b�'�S-��&QPL�U��t���_�{U�O;=�Q���FiU��qG6p9v^��}��'KřJ���� ���F8�н��<�ƟN59��wA{��ݜ�Ὑ�k}]��y&x��k0���y�r#]XKG�]�Mk�B$�c+6��r^G���*�	m�+�t�QT>T���?4�����C@��t�T�Y���k�������>�)����l���\]nV$��@P���{�:����ٖyo�χ���J��5)�Y�{%�в����u�;0'���]@[pSS�z���o��m��h�}��tLKtX�j��:
��/*���:�Z�(}���۽��|+�laC�X��dENK��]����??M��G���W�f{����N��9�m��bgJ��Z�,���O�6�rʻ�Z��}�m,�|�M��37.�r!@0���'5�̓Oi�8��N�Ű�ܽ�)<Y$�����$���8���C��.��P�*��X��LʃO�Q��BԐf�Gu{G/��1v�Y�Mi>{W)s��D:u>��쾹u���u�ۘc�Rt&� DB�e3X�s��ֱ-��Đh���G��,]nΊC�DM��L9Ly��,�\{uw����]&�����)�j@G��8�<�CsB����}� ��
Z�(�4��Z�;�A[9G�Gu2��_S�w��q��]|u6@� �ٛ�`�b��.��c@?E2���ի�L��f��Ùf΄�MBfZ��ͧ���Ι`3�u��Y�_ 8���˔U�۱#|�ye�k��5�l��]�J���h��o�τU�j�k?rP'ٵ;q�u�t����{�u��;� �k�M9mO*���]��wG<:��a��PQP�T�Vuիv}�'ry1� k�וm}���z���Ƃ�nW�U���0n��uhmfG�|����m"�S�N������K��
b^o�es�
��d�V�@K>Y�\�������3i���7�φ��RF�=w�{��3+��-+�����9�yi�U`E�Wf��`���hWb�.Z�a��׷о��s�Se�sv=�٦[a�����t���kD�0�~*���&4J���>�N=��v�ֺ�;]2�o`U��t�I�|��f���<[�ԩs8�T9��
�l�0ˣ��)��6AD�%4��o˩.G0��1CF����g�22�r\�(}{JZ6m�#��Vq��+Gĥ��J&ᗄ�r*(�0��rg*�s����˪p���:��gMք�҈.�*�)#YN�S#�y�-V%�!�xq

"T9Ars��T�T��qRdTDr9Ƚu�aְ���r��EE��ȋ���.Ue�`Gp��슢��$D+B)ͤ�G�����G�r.r�AU�K*�"��=wXDA�.������+�A�z�ID\��[��*Owsк]6�YQy������NDA(iQ*EE
�Ny9��S�4�\�EW����UZ��nuZ�W%#�s"�ai��DY�s���p��Y:iN,����*�V^��Ԣ5���*
3s9QD������B9;��$c�YDU�N���^��3�Q.�i�#�ER�Ӳ�eI��B�Z�T�x�8s�zJ�)��y\�i+�+F�EU̖]3�-M
�i,s9ziY�;�z!E��iнNU�;��TQ�8&��H�Az�`��p�_|3k��XF+��DKw�*�֛��	mH1^wZ��+y�Ky�����o+�I������p���y���ɭu6%���v�5�M��,G���ݍ��l�kkY���.7˫o�X �����I�n�����'�i����(u��d��?��L�O:���_i�O#�,<��{�F�û�e�ucͬn�R/��=���l�(�Oҁ�`Y�A.˘x�T;2���x�魈�_j�k���U�~Ǌ㱪,�^D����S}S��M�L�{w#��7����{�Z�	��Xr��~���Oi��Ҧ�(�Q�3�鎩�	؍v&�	�"V�>�=���ksig[�;�{U�F����19H���;��Pnݸ�nLm"CQ$[��X%�d��{�����"�9�x�ŶY�b�*w�[=�0r��\�%I���v�Tŧ�LGG���wW1�XF[�����9�*;������V&��݉�|Ni<o��BΫ�{���.���ٮ#��`)d�jOid�I���3���FT{���n����h=L����"**�gh�*��韧g V�a�ĢH|V��C댯�������p��4��$g�S�3�)WّVְGJՄ�;/]]����ɽࣣu�)K~�� o,C�$�ɜ#Q�)��*���-<�b:�op/�u�]k�<u�oe���`q��.X�ׂ����s�r�P �c��8�~���])�0�c*�e���gm��z���Z��\r����@�s�w@�ο�{��,s�p�}91=�3�Q;J��}7Am��x���:�4[�u����]�1�l�:�tPN�(���Y����]Ì+"�W����Tnx��fh_z̕7W��;�^��z�i����f�qA+v����pk�i��d}F���(��[�ˀ���s�}K�.��n���b���s��}���g=�.'�|8�&�}'ƃ��wf�Is��vu߻��s4Z1};;b}N2�Mx���P�Z�oӍ}@u�}~�kY�-=����N��W}0�;ٶ*�o��p}�}&��C�ɭ,^L���']C�}��ׁ{��W�V~�(�w@_]��T�����GW��a�Y�2��{	ِ�E����γ�Js ��V|i��޴�Nc�۸����ڧ�]ˏwʮ�=GbFჲaFl��C�t��4̊l*��o�{34Y>�Ef�͉Ol,�vU����=��0�J~�9E���	�h�<��EK���?fb߬��ՒoJc%2�z����ȺH��;�<���:p_���u~v�;�#�(�(�Sd,��A��#ݸ(��"W@+lvՌ�*����9ۤ̈�Y��n�!0��d��N��ۨ����gGs��d�K�/.���Ƹ!��A�������t�o��C��n�u��B�;�B�V��{y(Ϗ� ?��"~�T�&�P�㭪�߻U�\?�#��Q����[pg���w-K3Q#�V�W��RTY��J���.6�q�o~��|퉭Ѐz=�}����*m�n�u���)���9��0E�^<A��&&)�}��`  "q�n^W��PԳkZ��Y�c}�:�7�y}���1���	���pG7��zeH�9�s�nj��T~ݖ�[��Q	�+E�ul�Ū�{
n���9I�IQ�+ٟ.�F��/6*��y�خ�	��{&ǋ����t�6VhW˵�#�7Q�Ӫ����A�����+6_�y|��v㯀������l�vs�6X�2����7���:���>}'Nz��{ד`��}Uo:��]F���3��G���D�2�)��a��tV���w����c +V�r������4�Z�זt�'�O�٧���2���KGQ~��_�������ʓnlRR����Nr�B��H����p7[o��*-o��T��V�*� ��E_�1~����!��l�ۖ��su���1��Zv�E�B�-�%�>�-ג��z�)|󺲵;eH�>^v���k�,����q���{��fq��e�.����i�4M����@ʔ���-�ˣ�&�]~KޙSKw�t֭9�h��T�C�a��W�׾��}�����}����6��f	@(�ʧ��1:g��묟k�+����=�w�cldϺ^
�F�U������>{)���=����:�Lǫ�\���Y�:�����)�C��g�&�_�^O"���)�Lv�|�{N<��Q�>��@��!�0�'���_��%�����G�4.v;����ð9;�}�)V�|������@W�F�R�lE|����݇�r�!H�وޙrp��la�,��GJk�9c��&&%��Q�בW�>[�����Mgc��1�٨W].�BT.���λ�<ߔ��Ҧ���z�h��G����.�t�_�Ο�zq�X*/�)J5�_�\~����3�=����]�����E��� �Gw!���J�=��|^WA�<؈~���1���`�s��u��ٽT���.=B��O���-��䪻N.f�[ڦl?��rK����}u�<���Q�dz5]���u��1�ګYĥǯ�ݛ�.jG'�Ǯ�	9��s&��cY�s�����)NĀ�у�M��}�i�׿�w����Xlk���ݠ��FP�b�'Ρw�%/i�Ƕw�'�a��{m�3k�20�n��+,rCB*l�5b��Ӆ6���V6Veg1��-����p�j*��I�B\�UԛՍh�1s9�b��k��1��>�$ב���r_�&�:�sX�p��yV���P��D��=�K�~G�h�h�y�P�>s>�m��(�O�;C���{]����[Eg�	�e�n������+in����#������|�"�yw�W�ƹ:k�W�9P���~،�t��U���я�V����ͧ;w2}Nul�	��W�k�/�V�d��N�q�0�S���SK��Ł'�t.��¶�~�J���s����$���G��ƻ���\h-K5uu��Lg^�S��Y&��s�v�:ɨT.g��ݻ�9�j=�ӎv�=���XJ 9��w��}��|������J*,�����*�s�/���A��;���
�ϰ��FK�5�0���@}�t|�����::�ly�����1���*w�&�]�������U������;�Z�1#'���}#����_MTL��Up�*��#]�4�f疅�k�7�o��;�7���w��,{b��H�b^��0t}��D��Gt��;�~����'��[�W���ߦ~T��O�,Y��n�ts:��<-��Q�U�L��J���t��ђh6�o���p{�+ق|!�xz��x�uF�9���~ِ�O=��;�cT-n	�ԍ��J�ގ;�W{i�y_Sl5kY&�0�vkq�{��߬=?z�hT�B���������W���Ps=� �qN�LH�EmN]�t^�=��j3���1���(*���*[9�Tw�iL�M+r��9�s�O�����������8��ȯG�*J&�*�&>���f���FF�;���P��;�㧲���h�׻�����[m����!_ϬN�a#Ƥ/!��+g$�\=آ�+�X�c�ӂ���c�gM�����ڨ{%\�=�t`�r����}7P��L/�^3��5�϶ҽ=[���K�OGM���C�u�US��i��w�!ǁ̣9��&To��(.��Me�����f�?�:5�R{�����Q�_���T��>�b4����Q���V����|
��C�e���p�v�޹�ɾ�c�3�X����ߏ2��|��*~�{Q�ѕsW��~�Z���:m�7z~�\N�y5�^O-t7�Ȇ��9���'�VQ�������.�C����Hw(kMz2 �\���e��;&w�s��ԻS13" O���H"�|�5���]ї7��n�k׹�r�Y���g��^�,�ى�.�N6!��X��;s�払iLb�;N�Ў���cn;8��\�Vk�`y��2.f����`�cY����������a��<Z�L�P��`>J�;U��Zޓ=P��?�*_/�=�zw�N��jǯ�gH���lI�'fC���Ҏ��M`з�F{<�m���mP]�d^'Oŵ/O��)��ʮ�=�*:�&xפ��7�
V}���+>ߠ��_^�BE�۰��)���]?���� �~v��S�Y�{u�>?P��ߒ�ۍW�lr~���&�����_��K+[�3�{�;�<��쭟8�3��3Np��N;�_ ����E�F��U.�(���y=�g�h�,����i�!O�Ӌsv-��%^�׋��cƭ[�j�I���!*]F�.6͞�g3˩�����g3/�܏���;�}e���{��Q�=-��ۋ,����ba}r��}?a	c�K��%|��&�n�Ϥf���u���P��U�p��[���o0�Bpz��Zz�B�K6��m
κ��+�����{!�=���iLq{�+З:�p9U;ut	N�W)<L�ʦ5M������<�_w[��0f�F�z�ڟI���z]	K�m٠�̣���|rV]����d9�<��f뢝�kx���+��7s[�m�@i�/�`����$���"/C�N'\�4��Ge>�n>��(sܬ��d�ܜ��0� `����,q��y�S�{��%ّW��la��2�1OYJ��@U�����Pd|���o�bnT;�W�_�>f��J8���T:�`Y�r�.TG�g+�X��?Qk��9�~ʨ���Q�_�e�Ȓ�T�1��?w�tV������]���j_��U+1Ļy9���Q��"o���Q�Or��k,����3�}�"�Q�_��W�<)׻�ߍ4��׻U�h�`5����$}eq/���Ү��y�
��9^�f�� ͭ�϶�����q�%?3~�t��_�F�Z�`?K��s��������z+�,�MYϙU_(�7�|�V�շ��5?E�V+��&|��P�nu]���]�>�2��AD�O;$�n{g���Le�/�v�{�!�/��z�eD�}[�����.,-�L��>�t����#�c�����[���2����;l�i�m�(~��j�}�Y� J5�}qT��_^̮	I�{��C���P�5Z�rޥ|Ց�P��/����A��QG#�f#z�S�PKe~��Y��M|g꬘8�w�ַkQ�b�ױQ`rj�f�=���FW����䨑� �t��d%B먏�X��,g
�`�;#�������{F��r�f;�8䝑i���hJ�̈�8��RU�f�f������d�	ŋ��{/ �C=F��y����9�s�����v���]8R�2�z�r�HԳQ��{��n=�7�I$���e�0�M(����[�"�2�u)��Ϋ���������Ϛ�o%#��_������߾�8_���)F��W�~h�������}�rBś�н"Ev�����M͎\�X/i3砥}z w��,�q��P�;"wm������Œ�=��p��F$S��)�������y3c�>�e�Cg���~�&����ҵ`����d��ģ�cGTMWG�c�_\���U��R��ѡ�㙇��2�=�W?#�b��۽P�r^Pv!]k�'pؒ��R7.s_�.��u��z'�«��������k�^���C~�:k�X��";�U��2�jו�`_���6����l�w�Oԏx�w�Q]��� Ԯ&��QM��T\|�V���Z8꣇KdEf��W�%���c=U�}��^u��^�L�Σ��|�#G��#[�Zz:5�$�Q����f9y�o�f��K/�t*j:�}�5�\9�c�N�d�;�n�����ؽ���}c������]��l�c�y`�`��C�ɠ��X�ڮD��C��Y��r��j��C�QV�8ck��u��Q�YX���y���{S�3��C�`f>(��*{5�j���/u!u���6�֊���f���ǵgJ뮟�-1�����}v�Tc��ʬ��	�0��`�3�9hg��&��[�$4+�&o4>n�_�h��Y�=.�������F�.P=2�ȹ�_�mJ�d}?qS��{ۜ;���O"�gx��KFù^7�{c��F�'O	;�TFT�N�8�v�[�����;}��Ϙͻ|��q�l�~���u��k��A�M�q��U�<}���u8��8ŏ�4���|����oE���yy��6s��Q��#!:t����]
���P/}3y��ۘ��.�bfctح����0�/1m�ƾY�b�N��g�Q@y��;��ZJ���p6��5��}��G[���K5�#����+�������S([�7Ի�w�7��dz������V��a8Gÿ~�"\˞�l�������3�:�^�L�s��7Qf\�!O��ݑkc��m������u���E,�&������[e2D�K��S��U�T���R�S��=sn;��'G?��(��V�|����T�"�1(���뛨|�D-�'���E�J�i��yR#��I�����%n6/��Ӌ���F�TaYw0�F+��9�ҡW����,����_Wm�Gs/hU�z�m����C��َ,��B�)c)M�F��@���wZ����JҮm���Hv��G�����H�p�5�x�hu�H���r��a%�_�)�{*���i�I���B��_^ս�dc��v��̳��|w�������[�@�h���{��d9�J�:��{Ҹ�&�RU��)��8�Uz�ǎ��m���A�����Y
"�P|����:WT|��-�J���/�'���B�u�`Z��F�۠VLh��\�Mz^��P���y�[�����=�`���3ëk2�Iv�袷��]���AhZZ��L��nW	]�y#�h+}*�1�~ڹ\h��un�FA:��������,�^J��m�n���ɓ6��]Z-����q>ff9Nvi�8�Z)J/{64}k�kAƙ�ȗ:R��c����|嚩����Nv؃�k�r�D��2S���.gf���0����(a'q,�J�b0�K�N����E]�*&�9tЭ�m�OIE�'!:ұQ��5��ߩX,����(
Jv��C5����\}s��6��*W׎�QǷ�+���
7hC���CD�4�MoF��DTH�3��T����l�rG.�Rs��OmE��y�g{t͖�(�o�6v��n�b4@
�|�S�����/0g"՘���\�Е�XzO(n;��v�5
�U�Z�� &�Ѕ�{n��E"뷼9ۜ�(,\�w[���Q啵��ŉ@b̀�G:�����sP��n�C�׋x�wՕ,�o�[��OՀF|̭ޯ=�-���XZ�]Ի�z��[���B�m���%�6 ��"z�ق�X�3X�3Q�qS4�.Ŝ�[�=���S6�z���o��L	��g�i���V�ҕ�Wf[���[(̽x&��kk�j�> ���we/�YwR[��%w{SD�Y��9���wJÑ��Zк��v�w���K�fM÷�2V鬜��o�/b��R��ޅ�8:��l�K{8[ˎ��c����Ќ������iW�K��V�l��E5�����]d^*58v;�v����n���+7����j�4}x��A�כ@g�]�9�>��	ZOkz��.�����,\��E�������q,��ďm~	bæ�yH���ӛ�)��L�M��u��X��u�6�;�ڏ밪a%�*u�uj<��(\#%^;�����G�"��
X��Y�wE)��Z)gN����b��G��|רp�tDg����N���Q��]��J�:4^��홽k�9ZB]е�|9���/�.�r��1��|g^=�[p��=rfأ�qN���#��m+y��rL��U��nc�q��oB:���>7{Ըܚ�U{A�r�G(�a���.%��n��M��7&=k��T��(2��ʹ�LDh�}T��K�
i��(>��K&>gs�h �^Ь?h`�rr�w�C$*rYҋ�<����u�w0��u/SD�DQG!T�.\�O2#��ΰ̊O'tw�MiC��:X�8�����uZH�8^�h;�^�s�wnt�DI�J.y��2�$��)%�tp��s�
��+��r��'Z�S�\B�6Z�!�g��T�]��ݹ����W��������G��7*�S�����ȎT^
C�P^{�{�yUz���v^���݅{ԭ���wE�;���5�t�BJ�50����U��)w]�n�p�Iu�%*K�XwEE�Օ¨�+�#��C-Yi���G	:QP�y
���9�I�#)����QHG*���n�:�����u"�D�Ñ�B;��R�
.Z�{���G���Z�e(Q��RUFT!ATy��E�4�K�,��wr��]�"�Ad�{��8agH�:G%1�ηS��9iUS�G"<٢��9�t�WZ�Ҥ�TUNT��=^|�����6��S/�R)�7|w���ZέO%�ӌJ���m��:�|��70i2�H<&�pGv�G5|w����3��N]��[�7��{P��{��{�¶�fߟ��<�Qe���i�0T��f���Ŵ��v[}C�5%������2����+��e���j�=���3���Q � �����,�_� !�y�ѨkO������Lvj��u��}ic�G��̌�o~�6��>;!Qv�֗�
{Z��}�.7�Tu�����vK��ʦ3�cc&w��}�~������U�Z2X\��\n��0�����Y[��G��"���%a;2>�n6���d<�vwV�fh4�閏`���/>�TG���Ӏ=T���qa��D�m���ވl��uiw���=7�mz���sC�)u����U���&J}A�.��y�#��z8*��-�_8����"4*~ԆX���	�xs��	�7_q��v��x�rkg��#�a��A�L]R�n�~�R>�??�Pȳ(��f9lW�B��h��K3���Q�׈�rjY~���k�y����#�s5nՅ�r��X �bD����̫;��|s�c�"�1Z���0��5�7�K<ӻ�.���~~R�>�Kgبf�qw{lQ�s*��R���xU�r �����0�`��e�������e��L̢1���iorO����޽�ь��z�㇁����N���݉�iꂆWu�º�'�-P+�B�w�;�P�M�3�1�y�&��i�6>�E���%��J'�(AZz��$s�.���_�MЙr��R֪���aU}|@\s�	���F	}V�;�����!Xǘb"��P5/�����Z�1N�[�g{��I�'vr����[�v�O�\-���#~t��f�/�B�F�@����w+���u�gI�"g��h!ۛD*���+zZ?Q_�7f����ٿ�U��GC�m�G7=�MD�Yih���b�{(�A�Oe���|M�fևy���c�ͥ,}m�``��"�j��K\i�;�4vz�6��̏���0��xTI���N����'t�~��Zo5��g;�.�6�F���x�9Ą������r�]�5�eX��m�1q�	�7Z:va���X����]����U��\_��Q��n(/M�&1=����F��喅}��Z�;��g�9�O��U�zw^��V�V�?1�X�t���́>u�u�#p-�l�3�w�r9�{
?r��U�e-�8?3'�3�	��fh¦谫�}����	�Ϊ3�����K��؏���4z������v�랕Y`��,��M�v�#�:���-�].n��o�ݘ�2�t��f�o4l�B
{s���*wL}*:5���vM!�;k�ꊌ���w}n�W^�	�[���$ۍ��<���)�}�4.�g�Ǹ��e�C�8v۞��V_u�j@$���mV�
�2����7��E��ȸ�6�3`Jup��U�7]x&�'k�b�w�k�������Ѹ��6��^l�(� w�T�_Iܔ7�����~qyg���z�����]��i����:�Ke��v9E���4vb7�����[���Y5�n*Ǽ���{��6�m��w����}�Zg�����>��Dz��a�����@=�X��KP)�}߱�3��~����h��؂�'fy��T��4._ԑ�G�m ^F�`h���ȷ,� ��yWN�ț����=��W^5_g$���Я���%����?�m��u�/����dDv�}#�ؿ-�	W��B��^�0�.M	��fĂ����w�=��L�3�<�����)��a��� _Ejǽ)�����Ҥ�=����4g��!i�R�}�:0�nWi��5m8��K�oE{I�����{�;��	���ۨ���)�t+�MqD�_�n��ͽ�~&r��!�b�;ϥVW{��wXͷa��\[TU�cuS���ڱ�@yD]𕄇�6v�|���s�I	���?��s�SH���@	d궹�.�ܞ��q���.���q;9K�[u�c�����
�����M�k9���<�������10���pJ��(��rgxރr���r%�~� P�s����5鋚��ܘ��!�u{������c|�^U���#�j��ϵ�A��Q?%n�gˤ��cZ��UEG�؜��\�ǝ�ͥ���uhnM����N�|�PXo�[A�p��ge{��E�v���G�5`��{�u�>��wůsBzC쓧�3�>7;,e�m¸��\�,�y����N�4N"�m�s���,�]�������������g�X��z�!�{c&w�c+��9=�X�}&�0~�ݥ�Mv��DR�/��6wO���6�+����d����߀Qo��>�9���vR.����s>U&��0m�C���a����5/���g�
��z���Gx��IzzlU(�w�z�Q������זp�G���a<SO���n�<�����8�U�B�9
��S
�w�ǡ�s�����iy�F���DD�[���eym�[��.�9梜wxmz=ӧ�˥L��R���?!��,����N';bfc��Nj+�� n7i��luG"�*��_ZG>�B)�n}��z@�3���jw��G�}��"��%X0��s�V��x�����}����+�+��u9g���� g��m��b�P�⦩�'�,��b�9�9�>8�zb�S)9�㞴�k2��w!��}f�ͦ��W+ZU�4�!�Hq7�ه،�l�7�:dٶ��庙b�����������uQ��KT4����&Oyc��c�.Vm鞶+�O;G��X��U��ϳ��=9�(�P��m�B%I�|$�=r$s�u��:�G�]-;y�HW�@w�YڛϭX߭�N����D&v\�+)����v��a�����В���ס[�
b�NT�d_��4�J�Q~��f�y9�r=�ճ���W1:�8r��5�����.�:}�ؚ��EWm�s];�'��Mg��u�[����'2Q5!�e�8�{"�_׾���~O���U��ݺ�|t��P{fl|���B��������f�m�ͷ�n��t�Џ��z�䋜�[��OT]1c.M���Tn>�J���!P�˽8<T=�����Q����W63&�5�\��sX��$G���r�����m�������s���e��d֕q��7��q�߾�*�d�󷣜��G�B-�pl��;{ ?~�ƴ��Ȃ�r�l��}��[���P_zF�I�����n��k�юh�+U��s��/Kd�-�o�h�]m���<k�h]�U#�'sm�����W�N�?1�X�]l^L���]XҲ=�N֜���|S���]�z1�Etv�ޘ���TJ�	���*GQ��3YY��Gj�a+q ��\��d��R��f�Y�R�{&�zs�*��朗��N���"�;�b\^��Lv�t��ǯ�x��Z���g=��Cs���K�P7�N-�H'])X�F�3=�u�:�]<L��g�X[
���֖~r;d�،��q�ȫ[v'�V)	�o�>�+s�أ�1���ڞ�A���j���HK��M3��*�g@���D�T��O"���x�������F=/��ϧ0z��MY���}���a%/M����(�WF���q_]
.Z&������1�/��م^v�wv��z�cdxt����f0�;V��*,��]Ȑ�}u�Yu�̧2!fTL�c��޻Ś�ǳg���ը��Z�F�\T���]�<�"��H�0a}�{[?��A��ۛ}�Ǥ�����r�탰�']��Oʯ�~{l���ʈ���Wru����Yu�'펥Y~����� ��?Q�"�ר�����47��8��O��Ϗ΀��� '��C�a���������p���d�52�;3a��f�
����P�_G Z��ϝD�R�sfOln87{�h���V�cY�'^�Bѓ��#�S�2�|M�ևy;��|L�������ޝu{�tO=�F�Dn1o�uQsџ.��6߮��(ῇ��Ex����ϩ��zr�X�X�����I�Q5�i~��)]3�+��[4��*�x2{�K�l�0�lԊ��8�yz&�b�{��g�Q�3۹�I�<5� XsT��n��T�ut�����׊������u�9����+�*�Y%����(A;lW<���7�mnGQ=h��k�~�W�S{�o�~U�lk�F�ܫ���g�X�w��>>��{Ů�Jk�2��=-��Q��n"��[rc{K�ƫcl>�許���w��A�9R�n�çۇ�N��@�C�hez������Z�ݑ��l���w�.�Hw��5�E����n	��}\#��0�K>�&\aٺ.g]�cު�/ ��r7:�ǳS��>{)���T�2T��J���K7�ZX��avI�"J��� z⩁}�07%3�}t�9)�þ�Z{�uy��wY�����e#��#K���]Eq��x��o��S��7�#FG�u`�g���R�n��u����Y�ȱ�:�8Խ6�݇Y�P��BU��2���ۍ�B'kSܯZ�Z��/�#����u|���G6�B����:��7o�6��1�)o���ȸr�j���y�/:�Qwk���/�=�/�� ��G���c��EV�Fh�ƃ�}Q�Uu�}���g����BF��g�m<8J��`�A3&���/m3��l��6�c!2����Oh5O�����קrroӗ*���X&5�6&�,U=�w��%�\މ�#�\����Jr�V+�8oe�m���c��o��r�r��Z��S;���Dt�m>�dpv��A*nض�x6��k}b��� ��Fs.zM̨�6$���jwO�&s�W.sc�zn�I*8�~��iZ�gR��n��N|fM�� *e�k��K4f~��:�>���F�s���=��"ʨ���ww��gZ�sŭ�C�9ӛ�a�P�pJʈw
�\Q;�����7U�+[��V����q�yӿHX�/��L��z�Ϻ�:	Ւ��+/:<ꤎ}�U����'��ߤ�;�խO!dY�7�hg�\���]���y�#�ޱ���QA+v����u�G�����k�^�:����51��yn����Y�O�g�'�Ǵ窼{Jgg����E��l��l��7�u���FGt�����,���TO]��,0?Y���֊�k�u��J���Dm���'����'�^��߉�2jp#���uGq�⸫�ݶx�$n�s���nMixN�,(��L�H<~�3����<�JU��/��]�E�����<hY�{�ʜ��*#β��:}éS��>k��
�c�oe��8��u����G ڧ�}��zl*����7�?Y�2�D��R��4��{��k��޺ړ1�fJ�[oA�Ț#�xP\��7 ��T�z�e5�׸q��f�
�8.w�՛�2��o�8�vQ�[Hmr��R��Vӧ��fJհK��B���>�B�b呣p�ż0�����TY�+}\��M��L��?Z�t��ޔ��BvU=*4�Y��K�x>�8�A�l:�}�~��{氪��^p�b6#u�5�"��&��̯b��,{a�r�^b\n��FF�uq6A�o���n7PΧ�Nf���fa#b��QJ��/ؗ`�s�G�*w�O�7|�j���Rt�|0�=�N��2���%p %��=�T(�����K����d
����<�����Z�V���I�~��x�s+фJ���^:��#�_Y��:Ϡ�w��qJF���a��e:����;�n�r�g�Ȳ����Ȏ���1�Q;_ja�!��z��}p_ӽ��[�5���I���/\�:��ƝY>�����Ug>���C�0b�(���oq�Z�3�%��n�s��n��^�`b���/K�J�lXn�8��E���n�|�F�?��lN�����G�k�?f~��7��5�鉟�/���Y����e���T��B�����e_�����]|���˱���x剗�s�Q��/}s��c=)����*"@��9�k�?�ni��Q!k�DΣ�4�j���+w_Jr[�R��&��&���"��D�y�c�(}���Ns��e`C�'�Ph[+4A7N�ɨΊ�T:��b�/��i�q��K�M�Y�?� ���'��d�������ѵp��8��2���E�Bmlk8ʟ{"}�]g��N�ܹ�Ӳ���g�8m����0>����ڮkDz\.�S�^v�N3�:u�__P��}�xŬ�n$�?)�-���u�[7��:�}=ެ�(�L�lO�Dy�˞\n��1oʞ�W>�oΞgF��{��Ȕ����{U�_\�Z���x���&����R��dϙs�ˁj�O��;�e1֪�������sQ���V ����'���0��סּ��Z�%>��V��=ٜ���6��ysܾ�R>�c�*���2\g���LD�T��<�^���<��^��07���C�i���f���wN|V�4�����F�\����E�D߲X��t�P��1�s]�]W���ƻ���v��N���<hv�*�(���Y%S�Yv��sPgV{=S[��m���JG?W�%K��a}�����:5d;�#�̠ 1�ލ#,�
���9;|I��p��XLLWm-9�wq�P�$xd��o��>=���|z_{��>e��`���F�o��o��6m��c`	�m���Ƀ`���L6���6m�Ƀ`�����o�l6��0l���`���`��0l�z6��`�1��&�o�0l���`����6m��`�1��0l���d�Me�\}$�+~HAd����v@�����`}�T�D����*�* J��J�J(��(*� T�	P*�Q(U@���TJ����D�ۊ�T�TUJ�TJ�U*"����E�!U(�aUR̀ *T�RR%+m	T�a�B��S�Ī���T�E�A*U�T�����	
R�R���A!
)-���Q T�D�!J�%QG��R�  �)G2� `�fj���������hi�lQ�UR#VdR��H*�#Z�QJ�p  .)@k2��hm VMV����QJ)E(��b���@���
)E��W(����Eލ�(�QJ)F��(�P(؝Jm���(PG   ԪPs+SEj�P� �`h[0��e h�R�"�k
��%A$D��DHn  ��R�j���� PX�6�&�����P�U�*i���V	Zҭf�@M��5@\  8r�Q+d@ʨ�-�AA�l�&�)L2�i)X�V٠���MQJ��V��h�� �ha�Hͭ�����*	$��M   ��"�Z�h R�ʠ*�M�iUT�2UR3U��
�&��P���km��P�[[j2ڥ�B��U@B�� �p4Q!a�h�3,h*�AL�@T�l��Z�!��4 5�j(I"5�64��F#Z�mU�m�T�(�*���	R�8  ��aYS6��-�����MV�l��[J��T�C#Pk*�ڢj�
6V�
F0�6��l�TheR�T� �N	�m*ڴIX�I)UZ��U+*�0�0V5�֊�Z�(ڡ@�1l�M2�¨U�*%�T��  j�U 
�Vd*�3F�֪��6j ��cf�h�a�UDʵ(UR�T��
*0�*�2a��w�>�L�����T����C  � ���a%*I`L� �C�E M&CDɣ)�S�i䙩������~%R� ѓ  ba2a�OԏSOD1 ~� 4�  I��2�E &M�	�0��8o�X�7o�8Z��ՉVV��b��ڱ{��xch�^Ԧ�G�� A���U����  ��X�����c�?���@�}�� �5@D`���$" ��� 
$#%!A�.��,�R�}yi�]� �B�y�X\�_��d�����=�jYJ4=?�_�~��^����B�nL�r!@�W!Vn�F��jn:{S7�lZS>�"XL�ܱ��o�-�W����Z���n���)�X&2����$�U���v��@���m<��h�%˧�H�b
�u���[��1���"�K`sj:QG���d���f-�(�U�m�iՒ��LǛ�cUd ���V�n�4-i����/UX����[�6�FQ��dR�/f]��f�t�ʟ6���U(�9)�3k B���v�v��6��ea�<CZcd:�s"�,a��)[K6f&�4�/f2�*ԯi������--� �@�T.۷6n��9��1(��ZႠ˄�C難vS��L�&�#p��k�1A�um�ȶR�{i����;X�j�١0]@�낔�c1U�<�܊�b1���i�j���+$��kq��)d1����]�0������S,��Kt�����U�V�[5|�'u�4e�.�«j^��Zr���&���������/�˴(� �k���M`b74�u�U���x!#t��7�-M���v��s3�Z�h{���X�&[�*y�sJN�S5
j�q��)�Y�2�N�Ӫ��D���V`Y�$8�6����0ň4`� �k ��bi������c;Z�"sa�wilp����+Mc�ӈ�3jݭ��0q�u�Oe�R�n�3h��JIZ�٪Z��L-���tNdAA�DԻ�Y"�b�iî�]j��
�z �N+dF�O��[���kf�Z~F����]ݐ1'jbͳ=�ݝ!B1;�Dm�E]��gTG_��(
�350��V�)�u1w�>�?"�!l��r(f�9w�7xt�<�C⾵u���Ѽ�y�� ���Ӱm$3�lM/��a�X��wX����e���Su%�&�EM�qLl7[��U�ʊ*Q�f��C���f ����ni��v�ԀӷE��f��F�n$�v��2��r��뼴��6%ZT�3F�1�L�奊I�T�m�yf��{�j�iq�dq^�n��8�K�c^�gwD�*�e��BUT�U+�2�kƒ�c¢�x�if�1-G	ui��k0�X�qn�z2"%=�U��n��x�kI�-���e�\��]ֱ��n!��(�)J�̥�Z�6��B�m��a��<n�Y�RR[���Y�[9��ں�^kM]ڲ��`*����xӹv"5x�h��h�f��ꥎj�W�*aK0E+/I����f�n�[]wBT��#������L��Ӭ�5�PI$�o.�$�یb��]J���x���*8M��n�֕�$�ݍ�H��j�(��pdEK����3#�H���;xw6'@nUܕ��R, �M'/KK3EL^13]h�˘=Q:�RK�n�r���&���V�j�(�ܠ#fa�ܗ%����T,�e���u�3 ;Xp�8����SU�V\��YlŚ�z��m�r�<�&�Հ���W�X:��Y��=��ŋE5�"��ՊF�1cU�i��+E�lRu�('"{ B��44�蜺҄Z��Q�@n\#kV��bw(mnf;C0��h�:fҺ{�W�RRV���Oc��Ш	��F	����u�M�*M�3�n��u�%�m�[tKH d�T"�5�T�db�����z��wr��kH�D�4�ڻ��ԛrAtov�ۅ�F@T"�ځ����I\�����/��%:�[w���f�%���9p)"{wqAx�X���n��6'X2zp�;������L_�S&�i9���tS[m:	,�iV�.�h�&��`T5��sj�h	.��r�
�M���s7s0X.4�Kik�Z2S��8���ؖm�-+atC�J���uޘ�Y�fLk�[��S�D:P��1��.�'a[�-��a���۴�滱h�V+Å�`�]dћ12�ܘl)�n��{����\qma�6P;���ؙ�}e��i�Oڭ�!)����R�����tr�l#8�+�F�3.h�NT�	���J��B����m���]L�JȮ5��9t6^�Wi��&ˉFaҾ��!W�B�#ԉb�/6��3]˛���LZm���]=P�R�[F���w��K���/bօc���w*1�\�#vRV~��7���Sr4v����G����K2�wU,��9q�,�&��n&7u� ��͒���z�5hF�rꮯC�rXnX�aA�r��-I�a�B�4�t)e�*Z:Y��M�r�͵lG��Yc4�0%ZUeE�1Q	7sA�m�1�Ujn�1$�˼��husif�5��f���9yD�N2��Q��M�J�Uݨ��L��]�R�4���ժ�;��(k��m�Wf��N�f��Df=ܩr�O���H���,T�F�*��If��[�S �D� n^XQ<{v�*��6�Ԗ��ǔ[���N�ʼ��q0bd�֌H�S��[/盺˔����L�Ԙ�1!HѮr�VU�X]◊�Mܡ�m�B�-����2
���(Ыӏ\�5���F��@qZ�mi���14��/�N�m&��X�P��o$�Tę{a��)�E��^�ƫh�<�G���F�X�Z�]\�X�6�.�k>�ⱗ���D�na��X�=p^��P:@O4�Z��X�n(�٢�SL�S�n���:E��n���jV�"�%�oeX�Z�r����K�)�T�a����Z��1iY/*2ë� H�{�ک��]��73>f��{@�H,��ƦFΫea��"v�-JV�� ����te�e����`Mu��$��`�6�9V-��qc�l��;ۧ�m�H�W1m]�f)M+:M3:�뷼z�d���v-�e:��)��
Q�\O/l�*�O4%��p[�2�mܒl֭7c�l2�����O��fSE`X�U/�6--���b�%���1��N٦1`d@uй3f�"[��u]&m��jj-���`�g�b�囓>�^��FU���t�M���[���#D��/�n��g�20f�nd�4��n��}�5���ދ/iê6T9�;Ȳѵ4,q��$RQCz�f�TE�ވ��2ʕ�a2�غS��`�@���WS���
��4�&�م|��g9�V�{��JԖ�F�-�XĽ ���������,��V��2Iݽ����t�Ȑ��e�tI�CvU��Q��}�6��6)Zû2��!'mVeiV�f�H�ǔ�t�ȕX.�0��˻J(��+(^�j`[R�e҄��|�Mڻ��yʘ�b�f��֍�N�K*���L�b�xk�݂��4d޺�'�
 �Ȳ�{BGI�9����D�E�Y��b�.Ah�m��a�Bm�q�i��T(�#7�͋�i9M֓�/wf5l�n�|��hZIJ��6�R���uj� �"L��,b1�m)OR�w�/>ۥ�"��Ã��&��3S�j<�/�=	����*�,�2�*9tN�B�x¡���K/\6oQ��F>����{$��Bb(���h�r-I��2*���P "V�3l�E6����W�X�Ĉ�y��}3f�Z�a�ݑ��sDĞ��]QN%�v/�ʹ�r��w��E�-'�k]�o�06Q�(%Nܴ�k�LT[x���2�Խ�xp��
�I-NSnKי��AQYxD��VK"�C�����ޔhIf�a�F�*�R�q�LǓ+Z�'MŚ�±k�Gj�쭥��&S���.��#Ө1� !��Ȫ�V�U�0�+N|���跁�PĩhAR.Q�oa����U�Ȏ��nֺɫS�]�N����Z]hK�t�W�V� 1��A{|��K)�KN�:��W3w"v${wHӺ#,%+6�t�kRTM�?2޴�B�Dr���E���K�f�y7&Z]ZH#K/7����*�v
li ǰ�	��a���X�v��p9#��֮TN��R�Gg"��&
6���l��$�4�ʒn�bZ�l�z�I�SY��*ڽ��n*=�ئi�.�����^� a����z�l�m9����Cܖ.��,�%��W+戡��Ѻrŵm�IV�I��RF�)v�m\mܢB�F�^��-�CPнh��A���b�dʲ-S�td�"��LU�*�^���bd�7P���b/B�6���;��#�mV�ʼ��ڏ7�5��;�(5���T5Rt�w�ܱ�����U�kibE̾�a�6�X��t/(%W����[i9���k+0�ٵ��¥'��Ż�X 2����eKD@�Ko0-K�74%���2�R��B���1++�gM=;zpc��=M������ESv�@Y֨b��mް��X��(=F��E4n� ��ֶaҒ�e�v݇�K]�폜���j�2�	7aYx�2SPX�gb�AaNt��bst*̣��J7�x�%�j�[^;�%؛�SM���q|-ֹA��%!��-5�o^!H����hV�m�6��7)ۈ4�K�J�q��;�a[�$t+2��I���Ԙ�ɫoXQ��o@x�X�*C��l'����VfnE�F�1fc��2��44�A��Ci�^9-�"m8�M	�5f�y��/1,i����i��屧S��j/
����ҦY7��OR_H�%)���0���J"���/a�XS����wY*���`��L���n���d�����L8#Q�؆nH2�;���	��l�8� l�T�ɔ���S�>�e|1`��Z�R9zP��B\�=�%�w����"�82�hX�2��`�ᡦ� �5�CaF�5H,����Y6|#D�&D�\�n��
�$.��J�Q���t+�Zm�p7pe�ݼ�H�`:��[F��9� �ƍq��*��b�"��z�j�v�Dл66�@�/%n�AȮ�Be�:)����y@9��8���A��m��R]�r�TQ�V6)Yx���6�)hhm=h6e��pc_j�t&�;8�vH����j觗j��+�a�5+T�C�J�2JL9��; ��\nӔ�kZd�{bC$Ե�zn�=ǇV�<��	ɓ&Pۨ����"ҬD�^�`h�Xz��F|��Y����[����T�V2�H(񪘀��c9KS��e�Ep�@�<��۷�����fe�N�����b���v�젲'&VQy�<P����Y�vZ��boe��:�n��Na���+F�v��s��Ӌu*��[O+7%F3],
��/
U��2��ch莤�Tw���N�6���[����h7�3� ����j+6BB �Z�P�W��k��i�S�%��.�3	-�n57&ٓ^Mn�B3
ofb�ͼ�Q�#c,(�4��$�`�:yMQ��ua��C+Y�636�����(:�G�bm�Z�UҒ�n#m�0j9��3�v��N�Xtb�j5��J�ټ��I<O\t�Jz*��u�j��6�����|4�`A�{Xa�1
![>t��1�`'0�eî�Yux�;�1�Sƞ�&��U2�[2��u��NX��'%�M m�Ղe5#ĭ������F��p��iH�bc(XG�MH��m44�.n�$(���4�[g~�33r�Z��KTVԵm�W��(�]�7Aͺ/`&bQm��[;(G��J�wZoEð2��v��L6Pw�A	Z,B���q�\i�	v�Q�SD��(*KF\g0k�j�.���{iqm1m���g~��)˵LX6�yY�Ymk�{0E�h(���ttbR��� ��y�K���fcX���{�`6�(^��b]�b�ZV�Ӄ �X��sK�[U�u���^.7�[ˆ
ʚ��K	��h�Z���������I���)�e�)Yh�42'���_��ت�:?1�[?ގĉN/�*GV������C����l���L+Z�]��W!1;{��r��M&WGk��|h�C%�{ݲ��ɽY����91�*r��ލ� ���%��YwS�����T�q �a7�4Y�*�)ِ%��w�.N���#u�j����N]�ɼݽ������G�4���kɴN�N�m����tӟ>;����c^nG�x-���i�ޢ��R��]�OIt�#ūUi)�]�Y+�c3D��m:9OU��;V�<�)����hesxF%��}��,��WY�E���o�������[��ۍ�����@5d#d����eu�b����TFAܦҼ���f�:��l�#�عFkyǃ0���bU�V�*�ջ�q����[#z�9���wnpb��N�|�E�Lu^�L�P�ׄe�t��h)�owk��F�+ӵ��ʛ�e]gJ]�pA�:����&_���u��wMJ�����nt��b	"4W<W[G�|��rV�V��b��#���69ݝ����{`0�q^3-��d� �'Y�GQM�Q���x�Ta��N>e�*�F)�˫�X*����&i��`�R۴�LV�I���J��tF;���#-��r�\q��1�DÝ�������=J�7w·�Y��r#�N<�ݛ�3+~3�;�Ћ��������-���vv5i�wݮ�3Â�n�'4��'c�6��˖�\x�)�0&�wDb��m��C)�Ѐ������'Ն��ҡbRxѰ�@[L��n�*u����|�A!� ��b���F��#��t��
w0���y��,dV�R�l�V����z.�ջ�Gk�sU:͕�Ư�.�l2��F��0�L�u7�������.��/�BtiG��eP�[۽�8摔�`�e6��%�jt(X]�v,8�G���GVV���e�|�v���0�kQ��Ab�|�(��/���V��ޫֶ�}����`WJ�����uR��='v+�/�ٴz��q�a�A
1���P��U���N6mr�g�t�3MN�{m�q�¸=޾xJFS��;U�������V���r>�oD�kd�PF��O�,��p
�ʑ�uuchɎ1c�%�N���Uр��WMZ�b�LһB!�{��u�׶�
%r�w�M�����G��]&Ey��5���NrM���̋U_,��[�b&vX����\��m<��e��F$E)F�=�.��+h�u�����1Ҏi٪�c�O�5�v�O��^-�9�e)T�����e� ��p7':Y�u>N���\TL�lG��+���#����F�X"�Z�؝�]4����Լγ�����m=t��0���˒��o�ZLQ���ټA0����O7��g>��uM�ފ���I��c��*l4�kFn��j�.�7�����Sq����u���3��zF�y^S$��m��Vb��;P.�7��b�z`����:��]G���Ո�h�錽�Ko�ml/9յV��:��q �캺���Lu�
���:��8�^kC}�:�M3 �x5K�,	�$fc���7��A�7mo�{��αwʡ���X.���Oem���gnj���l�J��G6��/d�h5ٳE��9��fqE�Gw�`Z��s�rܣʻ^<s+'Dt5{�)��b����>�tɕ�GSZ��&�N�)�Zj�2`��|�7j��Z�K�^{C85,��'7O��u屠Vk"�QJͩs�t��q op��i#���8x7�.]��<��V���6yn-\stK*[��S�m���c�/�*��}[�ث
۶��-�Ǖ�QW4�"��u=��	�Sm,`�R�-W]3�����E��U��s��y��*"�X;�oY{MԥLR�0����V�ؙ�v�i��5�Y���O��Da�2l<+��|΀t;�`a�f�n+z��Sk<�fh�������v5�8��귨5�`�z��%��}ݢS�v�X�r�eAS-N�+kB9�YܠH�h�`7�@���7tU��q���"��[��/�/�t�Ӄ�^�2���%^�����׺�;wr(���^2k0��J�&Wi���e聎�v��l��5��U�t��cV��v>N�i�ށT�}O/v�YN�6�����QF�3'�,�T��JG����ݫ�ԓ����`ߥ��I9ǭYÖEЏ�^_�N]�U撢f���q�UR��J���Y+]����'wjqS��&gR-�z�ծZau�^���WO��Wk������QA���sfZUwc��_.��6�e�p�c�Cps�;n�Z��Pu5}��j6�-�n�&c����=z(c�\�u%emnp:��ٴ�Φ[X��j�"�=b�8V���6���q@Sʝ��[�v(�W�B��sfuB�t.YVu6-��-��M��͒������B�]�|�����qZ��}-�)sλg�xۮ�1���hN�V4�fl����Վ۰Á%@e"�(S��"�2�%�+D��3��k�eˬ�@�͙|����5��oD�5�B�]˝Y�30���C7���^d�B,-\�o��5�iU�Wa��\M`�U���s���Z�e�[���	]
w:�"���x�ڕ������y�F y�"/xmړS
(u>�ż��L���RF!�6�MZu5��̡#�vR�5�Z�U���S!�?sY�
�Ov�00���q u��­7��v��uɻ�w�VAnd睹���U�X�aɶ�7��"��.�|6R��81�ʺ�R�� �z�����qoe'*�i�N��&gl=���f�*����0��3`��vewƶT齶���:n�����ut2�8�̎��,8+[9�$�Z�;y���$9�gm��Effec�P�lE��/�[��v2AJ��Y�ʔ���õ�L`��6>��.�Oh�o;�c''����9݅��r�Nj�fwfĒ|���Y����Ew!{�^O���]]l�^�y:
v�p�!��<l�Nef�Qx��`΂���r��=��Ǵa�upV�o8P8]s�l���rK �uc��M�gQ|.�f�<�$i�/z�PX������]fP��mj*�Λ��g��qO�d�2�я�B�/F�}F�5ݑi���7Y���>:��˺��;)���9�˖�#����sv�N� ْ@j��'���]%���(H/v��Ƥw��:��޼��9ۓq���
���]r@-9�\
�h
��p�@��B_	�i���[Ux6��h��T�)��t���/X�Վ�=�b�P�{���}:e!0����\�&�Gc�5�7؎j��n=�X*&VVh�)U�βĮ9�}�c����lu��EW{1W
�:
��t�5�M�1�ie�A����p���os������f�&�Yǖ��:r�	;��իr0T������fݭEs��{gy�3�Q���O
��(F��r8lED���Jt8�5�-��\�:V�-���x^,���̆
�V���
����l<]f����K녚t����.n�VR�����)p+�U�D�H� y> w�ș��δ	W�* X4:�"R|�*R5�8)�v)�y˻��e�Ƹf�2/�_3*�N3r:�����W��ZY���:]��6�gv����%�B��n�s�ߺ��q.�
H 
�Ю�`6~�\GoPt��áM;*�F���q=��.S����l�[N�O�]�W��7VDAZT�),ȼZ��x�:Q.뗭�ڔ6�(n�
�\�ڀem<9�\�$�cJ��y7���&��Ҟ!�J�����㘰wC�M�}�g���
��;�<Ɯ4A��r�d�p��m	���dp���!�7!Ue����uc�^��q7P;�.`���ܦ�{KR�)S5�S��a����7\����h��d"�kp)+PD�GF��m	ci���Q-��h,l�i��p�}y,4T�ΥƝ��8\��z���$�nsP4�xxu�+.��
9�����ar@9}u�5�V��Ό��`�]b�uK'Y�_B]؇���V/d\X�)���������xψ�K��f��YP��6��2Eӱ�S����vk��U�l��k8�e� T0J��!m���,=}A�����/^��gB�-�W@�VyX�4�s ���d0�ْ���Kי[�m���hO���g�Y5�%h�4�mբ�e��7��Mp�I����r/w�}2���[��q�+pW��d�@T �i+7��QaԊ�he;Š:��#����9Xݱ�B��s-�T��ͬA�}1�U���VS������ͨ��"Ƥ�
W(]��î��o����y"�ް&�Z; 9��6��>�蔵�N��2��� 3Uuu�*յ�cB/jf�}2�(�o!�ʙ W.����'(,�˱ڊ�tUZWa��*Ge�LtxwX�f�d.`JK�t*tSs��f��!����Y\��ُz������EuS�'�E;��ʆ�L�_L�]6ɥ��s(`�F�TW�8�J����;5�/j�fP�0[5!TW� y��G|�)܍�g���j��w���j#�V�F↯��}�nʎ8cM�ɬ�<�9ج����
��C���|�����j�Q*���63EH��ސ��;�����R���;�݆�^;έ�;���̜X)�hlK�TX��D,������כ�u�|��ͧ����#?n��K�1SW�!Y��	�(2k�]��,�����i�O��f�cW�����+W��UoR��rj̚�Jb	ؓ��ЮE��������<���|[o���ըd*́:�L��E%|.evc#�������a�+��u'n����+�ż�.�|nP"���C�y�0r�$/T�g�5�ױq��:5���:�P����Z�h,RkɅ={�P�S��h��.��dT��2��11����]�V9"���L�S�ΞD�D�%
���/%˫\�J�.��OJ�V!��]��lͭ��F��d�L�Җ7��7#�ʷ\�C��9k�H�r���rӧ�v���9Io�ޒ����u�{O��4.�:谰���2��l�r�nu��l�|�I�Xi�JުZ\�%�[�J�Ql�(<��e�3��z2�GՁn8]e\E�/3��ᮌyo��vɏ.TZ����p�JM�V� _Z�*�>ti�Nʖ��.!4�b�"Ժq���;�	3�2V�M�Y1�s;pu�k�J�(*��#�ZHe�ͮ�ʆTR�j���Q�׍��|�}9MT����N�^ku�J9�t�,�ܭ=SM����&,�-�XJ����G�Y/b�j]p�Og%��'o�s�2EZ]�.��Jv���;�����V�4���w���4)"q����jbY����EՉ��q7N�"$�^A{�qH�h�l_!�V}(d��p��ky4���1P�0�W�e�$�Z��oz�ά[����9�g1�0+�B���qV��(Վ9�E�Zz�gF���K9��ӘU��C��WR|�uHkCo�.��̾v�kv�cB�����E���2�r��B�lq��k��9ϫ.R��㹀(�┸m*x%�L�+F�\`��7�I�����Wsjf	��M��b�&���X���vuI�gcZ���7�SK5�-����Ou�e��f����۬���v��s�!Kkq3��M�4��v�nu��y[����t��Nk-���
�jV�󴥮V��LYk�Ӆ������7%
$�!}��J!dR)Dvb��v�BU�pN�s�zN�;k���׽Q��A��רq��s,�7�)�/�[��ܥxPm�vu���l�]S���]-C:@�y3��9���Qk�v���a1�L���Z�f�.��Y��Kp�X^_2鞗�Z����Y�����z��l�"溽����}Jd��������{w5^Q�o.�	�5i�%3zmZ�Wm�7�YGu�C�� ��L��NF�Ʒ���O��d1����1c����[��0���&Ǧ��Nu1�Fyk�Wܢ�"3� �'��*��v$�I���j(�Q�!�˪]X�M6흯<0���Jc�6v�q�)�7J��0�F�p���Q�#�YO�:�B;�rʶi�&��K�ޙ�,�*�-Ո"Uv;kwl.�*#�o�I��(��n��b��+�-�������o4��]��H���钠���N��Ϯ�þ=�'OB�
���,U�s��l��6c�3t�{Bh��Վ����u;loAE��?>��L%r����
�{���C]�tS+i�>��b�[[]}ku�$ӷ�@�6�s-t�m�p�֢�M�� ��&�fd�2�6�
&�ޠ�pom��P.�5���K��ݮkh�ۂhH6�Bh-<ug��ʶ]���^�븞�ƫ���'M9�m�c��V�;}��eh(��Q+J��\8��"T{O8�Ɓ�څR�
�V@���8EK&1�Ζ5�g��Y��H�eow,�]�d�<��$-���.���p��Wv%�����Ox����C���S� �*c�Λ�e��Vf������o�R�yr{\[���F�˭��Q�����_�u�s\���1����s����r��g�4b0/e.Ȱ��3	�,���@����-U���R�˨�Sԥ�IUΝ�/!Lc�n5��Y�)q�3��;�T�5��[�E�Xc�F.���wO�n����ɹϊk�O�}�#U/N!5-7�f$�2�k���*v4f��i^�:^�[8vl��ֻfbL��Z�h*�K�XKsUw�k����骺�Ʊm��FP@0E�-�Qd�Ұ
���G]+�v��s�r�Sa�cF�u��*�c8(bA�4�:ZY|�k�T2�T[q��E[�[HSŔ����xq��:W�E88�j���a��u}��.Aշ]%���.�خ:�-��h��-��'��۽�;��M����9}�M�������4r�
�n]"v�="��	0oOnP�������ZW�ם�i,+�*s�#���N�zk��&�e�j@�h���[�j�e�(��y#a��(Ƙ�r�f;�b`u��p#{uꀮ�/k4���SY�( �8�.�-w��ge1��>�*��v����)�W�ـ��9�]�
��
F�����=��[T�
��������|����n���J�d^��`��|t�Yf.]u��R��rW"�-!T�%a$WL����rol��y�|��N�KU++^���\�Z�6��Yr�XOgK���i%��GH���@9T%�*9x���7K-�ւ,;+h!���%R����-]p>�>� @]���&�8iJx
X]Y�W+U�I��_42W^a��1�~t��y@�a!�]�:�0V����h\MӦ�L��޺W|6�4륾t�!+	r��r��g��]0R�u]��[C*ڴ�[�@���ʋ�f�t�L��Vr��z!4��vPh�E�Gm��tΜO��ÐgrPӀ���y�Ʋ��3
[:�����q��V�X�k�Ȫ�
�r�x�Re��!�1��%����`9h`�[\���·��8�bI��X�� ��B^�5�w� �o�GV���zo'l;�tDɹ��M��}�����]wVE�M�o"�N�K��]]�:����F��ku:{��k���%`P'��f���wN�NW�F�OGZm}Nn-i� �F��-�GK���뱓�$���������"�B�@�*
!V�q5��U:x�9:WN��8- _��h�1��
\���lU�k0Qh�v$/��E�;n`�W����u;y��7Zq8;Vӈ�nt.\���}�]����[�z�u]���j�춐�Ix�я�����jL�T�u��V̩��==�o��xjcy�����}S�$�'��"� ��!��Z��u:��m�_^E,���A����QT��cE,�]����Pe�щ�ˢi���s���yF6��#zv��BY4��GEޙ�b,(�8Bv�OV��� ��W�en��Kq#�6T�r�����fK3 ��.�*d���LA�[��BBq0Ue�خh�#,YU�;�"}�����^i;w�S�pɽJ0�Ý��
^A5�tU�ܬ��Q����%r���؂��vy�n�����%8�Uۼ��!y�)�[��ᘃ��R7�3�}�3�av���0Ր�9�*׏st��f�V��X�nwJ5�V�<���+mё� ��|�t/I�^�й�e ��=V��͜rM���!v�Q�`P��N�<1Vmu*uw��n��e��d,N�f�H���9s� t�kN�k]�\����V�\��_ͻկ#Ӷ��T_]9�@�k7�H;��[gE��@��/n'O��+|!�M��ż�˭�pHu��4^p���9��{����7�mmvCO�Ʃqݓe+�<Z�ᩴ�����-��ʄ���8ˍ���ʖ�5U����]��搛{�mY����Yy��:7	�4�ư�U��dɜ٣����y����_Z��|�MYKPc������*����.��s�,�锝�A��6��%�u�F���;�����q}�Ϫ�k�-glӶ@w�vq0�����
y[x:S�lh�]h)����+�{��@U���Zˋ�.��|;yl4y )m�9Yfg'�8�r�4��8�s6��ʂ����蝷kh�r��z�1�G4%7��B����V�ō��ќ.np�jr��k4���8Z*�a-���0 �Zo#Xq3E�Ƌ
VPw�u��;B���b�n�)���Z�����U!XE�!���L�Be$�Y�ap��� �lɢV�)�Aw,ܥ��MN��"��A��w�(g�S���k�n�u9Z���.���A�95h�c���}(�#S�c�4o��7b�򑷽L�u�B;f�jy7K��kU	�j���e��]�2iqCW�z�%�ٓ��C$�&7:�{��"�u۸ EgdwA�R0���7��NT�f;��.jwgq*��1�p�6b��43Wt����@�����0�ιu��%䉝[����Y�\�^˭��ֺ%`�GBKo=��J�/2�m����x�aMAB}l�0���6M6:�o[0G�n�s�Zvk8*���v������	��-��unY��_����b�1b7>���ǌ�e;a�9���㝊^�M�i�*�-+V�}�i
���#�;�uvVPLcqqXn���zp�u!�����%_@�wf���&]�G�n��i��Bu���û��M�� �Ckа�#��}]����-qN�rR��]=��X�a��j�%�A�h�����=����:����z��銲&!�a4擖��PѮN.�Ұ9tM�5��&>�X�WVǪC�w��gg�;is���X|�6�`n� ��r����w}w}�dMZ�e
�k���WQ�J�EZ�};VI�����[����Q�[y+©�շj��z�nf�HS"�]*q�t����f�+iV���p���?^0�rT$+��XI����vT�Xx�}� ���x�E����.�H�&_e��!�#
;�P
�����@9����n��,N�oNΝkp)4$w�k�\�^�ч�
�fܝ�Y��80�*��h��@+�-�8oL��#I:4�;%��t0Hѩ6ބ�ޥ��Ĭ��b�{�f�Tq���=R�%���A��(*ĊE��Z��نp{Yh:�wJ��G�+�Ӱ�6v�7�yD��%�Z�uS8�@rp"�7\�ej����ڂ�Iq֨�bm�[ga��b�.kA͜%�������JA��Y2���ښ�U۩�)e]��--�c�])�t�U���@P�����4d�Qr-�O0��Ua��h�'�X�u���4r��]�:l�6�efj���ss5�@^�Ģ�mvݽ�lU�!)PZʹ"��]-������T�:(>\�P4+`���j�\t��"웸7�Gn�D�s]h|BV��4���8������gqz��Uum�Q���%A1�f\��9��L�y}k9r���)*m�����\Vn=6��/��:y'}��^�PN:��rz�oY��I ��&�*ûq�QLLU�Eh�ډ�x�1��t�.a��{Z��k
�D�c^��-`��kvc�����Z�hZ�a��*'�˯wd�d|�9�p5��HM��V�i����=J>�h@-C]&v��r�(ԺH��o��6n\�ۼ@dJ�R��2"���8QT.ϢNfDi6�YMG�ݪ}�5
ʶ���1Vo+�R�O�1� �*3�;�}ǁ����,�k�Lܫ�%I��=�Qk���ww�c�D�:�ǻ�z�{Y�w%&����)U�ik���5$�����ʨ�k)�(��ms�Kx݇1�tpgE֍�y���*7֙�W��]��D>�w!6�l�c4'a�Rnh˺H53Fڍ;U�1[����ث� ���[��܁u�*�qCT�&�Õ��9�ʠ�o�_�7n��3��o���Ml�+�]3�],#�˅ѭ/�3��M����S5�sTp�����a#�ӤYVEmL�������Z�:Y�*�Vf�˺Q=���ȋ��m�C��_J�e�u^�GjCҫu$�N�6�4�5&Zu�[7z��⻳�ͽ�I�B��{�:��9��iH��ݹ�.���)f�uW�GDR&�7`B���mE%��쭤�_u�qL ®�ZZޖR'����6M�l�%�m!��<V��J��F��T��wα
{���z�G#+��e
�9��ø5k��H4��Ѹ��Tr��&�dM}�W2u��x%�X�������A���u�u�b��`V�}�u��d����яM6�eNY�b��.�d*�FN���l�n��Ҡf��hٕ�JK�!T�uZ�$��c�W�%l]6d�Fnl}�b[���}Vɡ�N������jy@��c�X�!�v��������t��Ȁ�\�IH�
�aE�%nVFm�8g�(3�Ѥ�*�$�_.�gg3l�u!J]m:x���SHJ�t6�C�b���&��Z��s5:�c�Ö��ނ�v���W0�Tb�J]ޚ]}ة����#C73�~��tg�惶l���,Q;�h��es�%���H0�ppںjг��o�|��vsF�킺�V檵]��>�]}���ر=�C�����tIb�S�m�Z�au����i����{���iVf�6^���eۮ��7-	�B9�f�3�f�X�7]@ژEҬv`�1�Mr��D�c��y�c����5+&����s��J���)�`/B;�)��$G%�tLNPehN'*���@�osZ�A[�mQia�:��+pc��cT��Ÿ�k-���B��dCR�E���t���BK�!���O��a��Ҋp�bwfݮ50ͣ[����)��M�s�g�dYH��Ż--��ԕ�-.��X�r]��xʄ`�:�N�_uGS���a�`u����J��q��Jj�(Y8��_[`�J��|�ܛ�E���B��I�o8��"tY:Q�T����s�y�$^.�$�5�+�r��b:`���w�yk|�7����=��`e�M�[\U������a��i��K��� �R�P#��,����2i� W�GP�f���j�B`�^Vcn�Kk��48_bS��fU�s����BK�yJ�����I|�`ס���πbЬ7Z�.�g�6�lbi������8;�b�Іq	�Ve��t�գ�VG.�q�GD�(R޽��y����C�]����h(ժK;�Cz��S�g�J����O9����ˇT-�R#�Z�s�2_!k|3��?�J
W�`����W`
�-
A
$ݪFL��.U�5mX�����	e;��,�#F�n�5�/�l73H�Z��B�-���b��,��:�Ҭ�qvX�a�}Q�����˒�ju���z���p�Q��eA}��|�Y�����eC�g�ҧ�7�;�Ū�!������i�B�uf�ٿ���	 �"�_ށ�d��� �|}�}��F~E��[;'5%��37�P�al�I���F�
M����ͼ{Vs\`4Wg"��Q�_l	�Իi��.#8d9,�\����׏N�zd�ש�䙐�l��ю�:b]QQ�3��z�g>��[�P[���\���T�z4V`Y���qs�l�2�=��ZK�W��	�n��ٽ��68or��]ǈЮ�������!0@C���W��y(�J�P'B����^Y�H?�wx�WP�\貃��@��3�\�K�t,]�e����g��}��N��C���-Y���=���	o�ޛOT	Ac���/e�
�¯)q�V&��r�i�k2�{�'���h7j�%�i���W�۽:�;�]Ы��
zs�d�Ӗf�-p<t2�[����y
Ń��R�vu��.�F��\�Vu��]��2��Pu�	O\;H�{һ��+����f]�`�Ӝ��V?�V�qd7Z�+ō]d�%��o5һ:�q��(-�IG�Gv��]���ֳuR�oN��a)�Cb��wtc/p��S��38�{�T��՝r��(T:2b��*�妲���3L�a�*j[���:� �.�J���X���t/t�Iq�����ݕ��/���'Ltq�3����l}aq�S]x�2��ֹ��]λf�#U�ϳut��,�]��*����Xe�3{h�M.�cF�*�`�bi�T�+��m��*�2�f�.������jюYe���Պ�q�3(W,��-**�CTX*&j�)R�W��Z�l��eVV�����m�*���-������!����m,W�2����,�ƈ��*�4��.�n\E���b,Pc-Q+n������et�1Z��-̘��V�l���W���X���j�-TV������jr)iUF ,]9�M,[j,X�[Yj�1Վ����m�֌UkE��¦��,Y���Q�1�t�c� ���.��X	+E��UWHTTETfR��*�\�P�QX����Z(�-��Pf�����D�i�*�EkT�W�U�-�����~��aͻa��Վ.r!I��I
�܏a�u{D�o4N��@�;D�:�;��j��H3��(��!��rܓ+��ͽ��P}=Rt"���p�P�1�h[�>4��J���wZ;����Lˏ��)s��Y2���ِ�G'{N��m��Y��A��+����״�>Y����7���ڎ{օmwX��^�K|��p�c�;���B�T��knʛ�Ȝ���ժ�孢�[�`�U�����W��R��ם�nT�^ʕw���=Ƞ�p�Ur�v��Ps3q5˥Χ��G���ZM����F��!�c�����e:Q�Yz�wV�ZW02��v:�	=4���'���T!���/7��n-Z��w�c�(�{a��Uh�y^iT4����=�O�cz�}S8��\��>��$U�+ټʚy��ޫջ���/��MIE}sW��T��x�9�R�up��at��pK6��r�#�ꕻ� �
Ѝ�9�5Zt��c�.�"��à��-�h�;�0�]-;�R�yl���8E��Sa��5 =ٔ�����]3�l�mH��8#	�wX���1�Mi���^�~v�Q�T�Z%���/;�(2l[U+��u�R#ԙ�Čۥ�����85�=�c�\K��z9^�������":xTF��+�n􈩧�m����%��N3��o-�.Ὅ+�(����a`ݩt\�y�'��q|�&�T��g�[i,��J^P�0M�Ddol��5,�ڻ,� ӎ�����ie�;�L��|�։2L^��{�F�7�z�	�Oc6L��"�*���r��U�d�Dr{ӝ�n�V�Wfs�:��8a�G8��ApxWP�2%Ys5YD�\v��sY��_f��Ճ�@��#�ő��5龞4D�]GN{3v#5b��m�v��<;欙�L�_	�kw�>�s6�XwSt��t�j��%L�̇v;4VK1Z�?2kj��ohPZQ\F�y"7�[�w]�F�V9���|yhY�-f��m����ձS a��R�PY��Ką=�L���7k�M�������{=Ƴ(#�q�ޝ��C-�vCU�2`���1�Ӂ�F��w��>�r��f�n6
:����JT�	�/2�ymEї���彸Cx>����G.}�x���Nv���H�^�e�l�ut2�l`��C\�,zvc#ۙ�������۝�OGfUxE�4�\!�������rRͺE�N�']��ߗ<�t�v�<��V'&i��Bo3]�O��]v5�v��[�aci���9��ís�'F/t��=��������cgoU�%�Y[=�K�v�H�Z�Pm8�Am@۟�]���S,�Me��d^e��t�G��J[MJ��~�/"֘hF�a��W�n,D��|vU�dǣ�ͥ�|k���S��\>LG�S��j����ѣ�}]!��C�img-��p�%̡�f�~�ٺ=΀~��ɏ�W�X��6rU�ݚ5��g�6t��r�͢�f��gd�;�W������L�X
I���o4�m���6.��%��{L�n���4�����C2�y���U�᳴z����W�}�@׻
xM��u�iM򬛥$Hm^P8a<��j�T��
q���6�mLjU��`�)�
P�8GO�Y�]n�1]Е�}�;y�٨~��7�7gDw8��*�z�k�Q0$+�����}d��i�@7L@��17�ܪ!�L�� �_�B��.��j�7��:�X��F�Ų��*��������+S5���z��Y�vdOq1�T���W.�E6���}T���z0�ۤ���u���,̗�F�B1���/2sh:�Ǫ�]��uͫH?f�3/b���y>�v�>��1^�D7}}Ks[u[ll�y�FkF��uϟX}X�U�"��/x�]�W"�剚p�3�$bg]��v�yWnjU�bX�#
���7n���n��^Jp���)�A��n瓾ά��e��;����ݜDr�9,Ջ�Kk���_-�t«��kh�5��N`�LC�W�;'�iI��x�����(s|�bj�_+�c��4<n/6z�d��p�ʉ�:����P�����yG���MJ�E�j��q�ۤ��u��
�^�SNz�Ws�t�սkv�+���!�����eN��ۙ��әP0A��9Mt�C�Qp9���ن��vb�[)��z,V򹴕B�t^���t|!�vz��Ͻ�!'�3,�rϜ8f���6��c��8̉�f�,:��7��gV�ݑ�/ũj�0�G�cJ��)�H�E1�.�͕T�q���M����ԣ|�:ۯ6*:h�YUPj{��5Q��q��b:^"+����Sa��/k�r�g&V�H��A��pe�Pw����x��O�6��D��}a��2p��ɍ.�I��㩾,L_5;A�zi�Pgڵ��'��n�j<:Ϸ=����j$�$b�+&�p��L\�]��g}���)3��l�X=Χ�H>iәÉHi	L��.劜L��2�3����Zb��j�ѐѸ2�0��nt���5~1[��ի���1�wX����c��s=䞖�����Wf*:`Nvx��hc*��޵{u�K�h͖(e���T�ך��Pj�d�VzOU�X�pŔ�rk�T1"�����W:���U��w�v�����H���kǢ_8��Hm42�2/�cpӋ��{��'"֏�S��('�Y�~[��{�6�u�C������O��K0�rr~�Ċ]g^PM�FU���B5H�݊��t-�l�z���)���xT�8�(yN��z�;hTйTv��yɡ5Uv3cWu�+�(H崒�]��B�������'GF���y��=��Wǹk�*�N8w��\��I��e�h$w�v�
�zq0SQ/��Y��Y���햺��d�N����w]�}s2�kK
�&#�G�1���,��6�̣�� ΘN�-9X�M$@�7�*�S޼�b��<U��*ץ�˷�mg;}���/;�f�I�T�Eڵj�嶀��Wr=�/�˽�;����߷�|h���h��;$G)����%y�(�5��3�����Bê;�v:�T�=�)}���B�9��i�ۢ���I<�R���.�����x����˱y���eN�%o����aQ�b�O	��!}¹�V�A�0��Fvq�}]Ozq����Ѹ/�eep���}-�U
��"��ꐡ�C{�(Wix��9<-hק�Ӝ�|s�^�i.���y�}!��-�B.������vv�R�2y��'*�-0�2���nF�ʨ�4�ΥK�X{֗���	��3�x�I%Y�V�����W�8��W93�{M	���;t<�9'wV�Q��zS����n�{���f/tX� v�>�/�a��;;.�=� Z�!aJ�ۥ�2�4 R%y��S�b&�Mt�K,J�p�	��L��Z�^t]\��Pe�'����ܮ�Xs�$��&��S�&�kJ���~���;jb�w���eD�q��۔�y̼>�W�S�`ƺck����T�\�yXP�+��Yj�*�Mc�iD,#,�� z�.v���c�C%m���[��kU%�4�ڋq\!�s4r�� �ށ�z9���̮�E-���nש����Y~~P���Ə:�V�c���ڞۄ��U�T�I�Tʂ8>�!yG'��E�
F:���*�ڹ�Mͼ���5*��~��zP��,�L�H����M�Ew19Uv�9�}`1}>��|��W��i��˞�m�e�a�궆��i����X��Qi���*;t7�ۼ��:WwC��������ib�	�K���^���,Ȣ7�V4�Orl�՞յ�,�\�=ˈ�r��{��W=\k'��+�Y��x������?\>����ۯz��~2'��:��v\�׳b:.���LU����� �.�T<-���_>��]��Wnv�M���>kd��>�4
f�@��lM�eGCNW������W�*9��Ρ�8�^ԡ��]�����R��߻�,5�b�t'�^�y#t�t��o�g�\s��2�4:܎�T;�Kj(7��8������OZ�}X��UTİq=�BV��S��������5:�7��8��絤�Eɘ��'FX�Ck9��R��/'�G*03�%�Z׽^Z����:t:F�����k�,L���ǫ��N�D( X8���y�#�z)���Q�}Nz�.2-�
��x�bs���N�ʹ�s��j�Μυ*��9l��x�����8WG��qt5{�lW%p�����9�3����6��^6�5U���Ӥ�MaK0o\��Y7�J�Pm��N�b�󫶠.��F��Nk��Tk|��iOK����::�0K,��Jc�۳�5�*�Ơ���AN�j�V��OO���}�*S���������t�6Ps��^���@;�oGp[@>����+Y��U�wh��_v�\�S�8Gy���ADz��!8��M�L_C�KJ�ħ�6e����Z����n��#�`�Yڗ!����������b�klQ�&��8�ezH����5+Whw�YO�|hql>�ו6�mgfrvx�j���=�A��Z"�xߧ*��b����w&�<�yc!���S�٠��2�1�T�Α����9
���]'n-Pz�js���m���|T�>=�S͙ov��:U[1i�uu�)�͞���nGj�����%��	��U��z�3�yY�"��FSsP�մ/7�SN|9��oU��4��מN�:
��C�˲�`����
��M	�2��.s;V�.��qU�V�[ԯC�p��	��μ�6E&{_���#߇�g�;�&f''+'G	�Ȉ��ɫ��1��O;��8r����jν�Mp�p�^N�A7:�l/�vLo�F:���]�Ok�͵Pf4/au������k�:X�>�1�Z������Q�.e��ڳ;;*�i8�g'�)W@ �=���7/yLz4�P�G�@P}��i��k���ťw��<δ�-f)'rr(�����@o%.��<	�����@Ԇ�ΪT�t;FR��(<���J��s�̗���zV���+�`�:�{r�
�,Q�y:�F�0��Wu4 ̷W���ctSl(�𜄢C�����7�Y�В���N.�˺.d��a��-�o��C���K:!��a_}*�
�{Md��%Ǆ��]������ėA�]�iZ0��G����䛩��$���V��1��j�� Z�r��-��l�ؔX�9�j�8��m��m�-W��P�����â}���vݜK4�����v�6�f^�@�u)��F��̗l�����VB��S
��S�X�-�je�v�}m���u�������p���zeĦ�Mn��z�7��+��*���7m����]���HV����Ò���PɆRr��XA@��Lq�#�b;�1�2�r�yy#��Pi�띚`��vćW3�S�HA�斥&M��V��.�t�6j�9l޶>>C����w왱q����o�´H�N�k��\)��ĩN��C*^��M�
����塶�K�͘qe�z�1q7\6%E��DՃ�S�0n��]�u�v���0w6%
�khR;ά������C!L�wYf� �L�zai7e��6�̨h���{�i\�PCr�T`����	g�T���E5��;�*���'-�*X�'��6e��1L��t��P,��̭۫.R����ƭ]qwv������{a�¨�aȰn�
�p�3�ǝ�2����~O��^�m�A�H��#�/��u1��2�m��I�F�2�M�;�����Թ��8��,�ה���\�xh��Rk��]����4�ɚ�j��:Qxb_,Ae��dY�\�M����Q+���,@/���,�YB�N}�49�r %G�[�	�Ѽ�K	��+ �"�.֡LFE:�z��֢;8w/T��w|�M�3n�#���P6�;����ז��:���	��On��e�MJ�T�qd}� �P�,�����}RE�H���F(z29j�
ǰ�;��O]�㽉K��Y!������I&k��i��/o�K��C�%�2ஏ���g���g3��l��VwJ&-��m�m��%��mDb1Db�"1UE]#eX�cdӓ��Z�F���(�EE5�X��QQ���
��ł.�2b�(�*1�X���KR��l���Պ
�MP���*[\J�Kh��F#i*��)Qb��i�dDTE-��EӦcUSIX*���QAU�EX���U�2��C�F�Im(��UY���FE�b�m@\B�ff
B�������QER��Q[j�A)QV���*��A)����QkP���1R[b�-�����T�K��&��YUVV�I\�ӑX+�����sT�Ę��ZR�3T�Lu��ӈ�֓MP�Vi�������֤X���V��J��et��k&2��U��QEef\��J��~��q�4�~�>yD`�Ҥm�VM�6Bl��ߡ�Ou�F�K��}`b%P�XVRF},��>��������
e:�[�-ag���kX}k��'��|��(���V��m:��m*<��2�nP��1��[J�[t�mmn��1���[��o%!^��>a�Fc����y
!~,-�}���x>��d�Ӷ�������!m>�,�[j{�\%Ʈ�oh��%�lv�Z̴�8ew+��g�K!�w	��i��<=\��}º����4\ώ��������Ү7�k�5��ck3_wVM�QP($aÍ�@J�����k�r�䡳��ƕ�v��jT����@��}\"�;u"�g�5��{fW�t�����x�b�VL���!�
��en�Tv��Ϫ:������N���.S
B�f��#ޤE�ٕ�K������b�踳ҡuCyp�����xc�]�̪T>\foQ�ː!Y��q]��37��Ŝ��Ys�{IN���{F!^ol]��4Ʈ(��ft9GH�pp��w5	��[�52��r�lmM�b�A ��h�z`�ǥs[��Nzu��[V̷J�e��i��ڿb��S ���x�[)�ʐ�o;*�����"%e�B��n���y���=�K�s��,�6��-Ұ�V�+�Ov�P�;-�S�������r��XT�صm�rw����JP�7_ZꨈڠU=\�3�]lj"�ucG5��|�8��y���k��m�mV0;�E�l������\6@��W���[k�Q����k���#,����q]U�� _!^�.6�Gq{|�<�*ɣ3�Y��/;�#�v�;#���� �dr�k�\�T˄f-�v%����\�.�7��Tĥ��/˅�ˍΨ�4v��
��-\��V<Ή��#Z��j�%Y7�RD���yp�y�Z���� Ug�VW7�欮�\�z���R�}�,9*�9DfpI�&`c��|��U�n<�o��`J�pB�Ҿ��f?)f��$����;VS�f�c&��Zt^�#*��3�2��9�n��9}�ʂ����5�x�)8�oDGZ�H����y��b��Ĺ��	�Gk�hພ���[��_��c=K��1}>��[�"5��<�������㪯x��a�" �6�@��S|�,���a^�EF�+5��W^�UJ�����eΉ� �o��;���@r��Ub�ٺT�J����f!gv�G"_EN�uz*���6�1�T�:0����n���u�"�����K	=4�ɷ�0(v�1�sgRU{�Rs9U���(z�{-�]jGj�X�ɍoheXͦ}���e�n/;�x�۹�Q'�ڹb}x�f�iU��i��YO,������x�4��Xr�gC�=H��S3�
�l���f��л�	��w����u3hJ!�7�Ugzޙ/���>fdA����g��n�L��%\w�-x�Vn�dֹ \��R]��]�W�*��O�,�1�r�؈���Ȁ�{��I����y��:n�W末�Y7ܦH�al���X�ߕ���sY�\(+���v��G���]�N$b�f�[��̀��B�j�S����Z�%����Y춳Ň��=�)N�׶�
�8�R�����Ҭ���)c���I\�y9��+y\�IT.#<��,t�sthL���If��ݖa*j<'i��N����z+���?{�0�;5�[N�-)�L4I�h�����M�Lv*�|������Tb߼�Y/oD�A�v\�k�9�tc���Ӆ�
��xN�}b��-sSe�gT�Y��Cs�|
�p�U\Ȋ��b�ɉ�	��ז��6��7XtS�Ѩ8�2|#�\���]�x@z�ؒ���ϼ=���[2z�$�`v�2qS�H��g��qX�o���l��L�>9��Y+&}{jI�M�2':�={ֽ����y��gZ�%t��0��딚C�'���4��G�N�8���RE&���s�$�:��C�=k!�7��� |��A��7f���b2b6�UA�?3/�U|��=�[�^��Y6���جdTl��vf�2���J�/c�]Z�b5�`���[¥F�Ε{�2�4gP����T�]|�E�O{yW�ʲ�J��(!������e�70gv�Y*n��Y݉R����>���>�����L�d���,�g��}CL�d�;� �'q��N�8�y`�=�Q�����a���o$_NS�Z�:>�w�4��'���$4�wE	�'ԝ��N��w��4��(q�<�2M�$�N2mOO)=I���Մ铌��\�f�mݺ��U��a���g����g���	�1�A��2M��E&�L�<a�'�1��d�/[вORu�&�I3�M�r�o��;>۾�μޖ�-|=D Ͻ��ݕ�>��>��I��	�!���RN3u��N�O��Hv��<C8�X�q'�nA>���g}q_��V�*w�&�+:>���N�Y6��`s�I�'���!5�d��i;�d3�C��`��<d���X�x���g�4��,>���\���-�jM�|<���9����u�I�d� q���=��I�������|׬�	�O@�;d�m���O|+� �����N���~w]|&*�ͤ��Xu2��5��ԓ�N��I�	�u<��I��m�鞧��a��u�m���{��$���*�M�����uY5�������
,��3�,�"�,2}l�Z�2k�u�O�t�x�m5�I��g��>�(R<	���K�{�+�EU���g��i6��9�jM��&!�'�����$�"ɻa:�|���5'E�a���!>`k�M<Bm�=�����Z�V����ﶩ1}����s�p:f�'G�oP��i���8��LE��!�J����6�>,-$̿ q�?2c&�����������{���\h���S�;����V8`Лa���B�ևvLz7MtK�B�M�CI��[���޶�8��f�7K�ܩ���uf��u��	Z������$���$���tЃ��Nu�clgZ���j]��嚺�U��D{�yd<g��'F�ͲJ�f��Ci&���i��Htsy$�gP�0�*7c�I���x�m�X �����G��FS���������z�
>d=Agi1��VͰ6���d��Y��h�M��8��,'7��[a��@�m���d���w�k��>��{�w�Oy�w�����rf |�l>d��k�	�!���t��vyH(c'St�d�{��8�$���8���sx���7�y�s.=o�{���{�a<d��O�N'Ya:gl���󚓦m��;a��gu<�z�L�G��)8�yC���7�c�>K��힕f�}���� �4�c�}�@���>�5g��3�'�XM<`vs��d�!�Y8���VM� ��Q���x񬉟�|���+����W��%@�<��z��C���l�2N�0�i9�@�'n�����x�t�Y�q�\����:�&�I7��빴v���W�������B���|��L݄�����7Մ�{��<}Bw�p� �k��;d�|E	��T=a�N��1	���A�fo�秙Nk�y��2s�a>E$�wğ2r�yI�06��7�8���=N0���)=�=�sߺ�qĘɤh�z����鍸�&���_W���x��>g5H|�L�r�$�'�o	�I��&�7lO<�z��;g�VC��Sz���@��Y��|ޤ�f!�[���O;Ο�ߗ�y�w�ȳ�I�Q��$+�|�9���=d�\�a=@�_d��I��N2m����6ä�o�Cd'3�ȁ�G�V|�����3�S�:f��O>����Ӂ$Q�[�|�uu��8#oN�U�-Y:��.�55�-u�T/�i��H��=����GV݆��L�V,Ey{+&�kn���$�|z6�=F	[x�ܮY{�S{��t|3�m��s��6U��3s��4����Ϻ|=����m�|�E��P�l�'��T�e���.I=@����3F���{��X��d 8��Q�lv����}�r�p;�g�����8�Ę����$�
�h�ClRv��g�6��dP>@�O��$��OXO���6q���g}+�m�qK�=%���<���3�ןa���q��ba��0���3q%a��Qd�fn�'�&���O��@��4���:xg/N�z��{�;ם]�x��=�Whgl�=d�3i��3l������<CH��c%Va��M�Y4n�,'�%�'�؏?�����ߺ�Rέ�)��N�9��$6ä��!6��Tv��;�3ĝ3�Y'l6��rf�'9�2v�C�o!Ğ2b)ַ���0Z���<�J���{��."�<I]�sVM���C�C����:�Xq&��x�<B�g� E��H�
�U�L����v��/��T�d�C���T=F�C�Xbz�}�fIl�{a�$��]�O�d�&3i<��
bC���0�%!G�i�W��oÖ�?
 �{�~��I�ﬨ2e�����*7|jI�MQI�ԓE�4Ι4_r2J�nɦ|�k��2q0�9��y����{�y��}�OY;W��%I�9���v������tsx��LaϨ!P������'�;g�O��4�I=�xx>�}������~Z���VO���3�8}N��'��ty@�&�8�_`C�ϼ��VI�u��8���;`v��L<�����!��;ghM��η��� ~'��C�|��j�c�t�r3�$�=�.���Q�јP��mه���Α��W��۸?������1�O�)�P�C����3-z��vLX���8�d]�Ғ�vü:�%t�ڴ��툪�ܩT��{�H��1@���kY'���&�qMN�$�'-:��v����}��� ��0�;d:��G���>}�{��<��u_֖Wk�}��	�'�l�g�C���׹>a=I�z�6�I��������l��ެ'HO�g�OXo�`m'o��w~cU`���3{�g�|>_O����ǣ�,�gia�d�3�T2kx�Ou�&�a=s�'̜�Ğ���dW�ϼ8�B�ߣLӹ�S��k�,�Y���a0���o
e��B��K�(���}E�l�!���2|���=I�Mu�!��9l��û'̟X��<�#�ڬͮ�104�G��}�	�!�y����'S��8��n��|���`��I�u���I���<I�Xte!�M�u��'������Z��u�9�����߷�����M��x��w��$���Ϭ������[!�%f����OT5�=a>CYE��P�-���N2p��{�|�����oZ�|Ğ09�d���;I6��z�����<������m��i��$�2b{>� (m��O��9�yO�V4&���u+��W_}�!Bp���=���d��iya��	�n�3��ͲM����~�v�:�}�l٤��I�:d�Y��~����}������M$�s�R�'v�f_>d��:��`q'OW9�M�:;d6����FY�	��ʐ,�Ͻ�a���!��V�4�S��;}u��<d�!�^�>d�&"Φ���B�ktr�6�S��5��0��'F�>d�^P�2 ��C���M��B�^O¶���\���%,X*%]���P-�ٴ�����6.	��;ݓ�7g���_3��T��4���0���ޅ9�-/Q�3�kz��N�vL�5�Fi�ٻ�0G��<�^:}��f�ݝɢC)rYS�5�76�!������#�	�������o7���X���N�c�!�
��m�|�ݔ�M�3 z��d�j�)�`O�:��;���S~�~�K�ܷ2����|(�}���� �Ȏ&�O=�ڲO��xd�7B�tɖ�7d8�XotXN2|ņ'���&|=g�}��d��m�wUo>���{՜=����Y8�$�{`)�"��)8���!�`>�;�'\�51�L�:7`v��>{jI�K�tq��cT��~�}������ɯl6�v�]o	�B|ΐ�N0:���'q�I;I���2��4Φ������L:LC���k7ֺ��{�9��$����&�<��!8�@>d�8�:a�z�8�!<}I��"��I8���	��{��VI�o��?N9����J�+��^dT}�ÏNoxz��'n���!�������x��6��Bx�`j���l�VI���q�h�u�'�2r�zﯹ�-�����%�z����l χ��P[>|v�2��=a<f0��2O&���Ri$P񇌜g�VC�4ɣ��OS���}�A#ެy���ow���_��8�7I�̜��������t}���I=C�sx�s��I�cw�I�	�u>�I�;Hk,<CL�d�,Y8�����*"�ȉ�yܧ7.�'����;��}$��䛶uBq���u=�$6�������i<��!�s6�+&���}�i��i��2���C}�v��<�Ov��,*CĞ����u���d�=yd�ݤ:�P�i:x��̒}���!6ɻ@�;d�m��0��+�ṙ��B�h����U��ޱ�nؽs.��S�P�a�	C~gM��H�k����rn��ڨ������SOs��
�T��·4s�Mk}�WX2��.��G��T:L�n"oM�u9Z4Y��tW#1UO_/�xxDZ�����P�~)`t�E���h��eh2h�ԓ�K�'�&��d�0�8����3����Aa2u�mRv�����o����[
�St����=���{��I8�a��Qd�C��mA`m���ՠz����֡>`tg0�<I6��x���d�g��﬷���Ru��r�;��{�ݯG��D��ܓ�tɈu9�	�J��QE�m�O-��)��|ԝK��8�y��z��2�eh��c|��]|}��!����&���ϙ'�7�$<f�;��tɈ��s$6�P��M���,�ZI�_�8��0���#�~����f��O����U�?{��fЛC���m�d�:5x�<B�F{��6�ts�2v��7��O1tkxC�*M��$�Qd�١��0{�#+�}��wV���d{�j��	Y���q��C�x�Lu`,6ɴ��I��g�h8�$ǭ�q��X��C�Kl5�� Tq��y��;�oμ�����a6�����Iγ ;I��d�������:N0:Cl;)d�m$Y8���"�6����dG�*o���c��Y�3@�Lj}Hw�a6ɣ���N��t��6�l��d�f�N���t��q��
��?Y"�9;v�| #OM��G�iM['sޗsoi���^��d!YyxVV��7i��T�Ţ�1��uT�x��K�V9�eT[�o>���dڏ����3�pX�<�f��]�eeґ��X�s'��Cw�EM���OM&Ծ*�Y��Cb��00�u<�D���w�q�y�!Ac���S������V���ϲ�ooF�g̾�Ǖc�t���2a�AL嗯�X[����Xs'A8� `��i������p;�Wa�L���Z/hZ��2�����GFnk�=}WQ�y�ke��8����üNoj���B�9��:�wPy%0	��8����x���{��Q�.��v�d�J>U٦ed� ��RU���S�s�7/}��v��K�s�#�vu���:h�E+���((�JtI�q]����&SŗusG%�(�>B8�U�����M(��&��o���r�/��M��F��S���V��:V+,��&Z������6r�|��]��̚�]�*\�ce�!��]2���x"Ov�Q��&x!۝���l��sz7�kkۮ�����H&ūY\P����x3]�};/��� E`��8N�{l� ���I"�k9�A� �U�p����Zs��W:T[�÷no^Y����>���B#�R�����e��B��e��z��dy��/�z��D�tM�F�;Y������,�w�Q[Q��T�Ϫz�9�u�N���%Ժ�˲���WP��'f��dn�+�1ݬ�J�%rj�._}*�N�Pݾ�V}z,r��N�>�����	6�%�ahj�]8r�� �l����w@>f��*RDR�Ev��mO�`J-��UH0��@�^�P�n��{l^J:�7��j�TS�Y�Q�k��Զ�v��2�\A$�nnXST#~�#���z�΂�9,K�eA�B�[ȍ������cX�fYH���d�aޕ�m�	Vu�Td&�\ˎ6N�L&��S���4M���g(��h��Yx,�6�-؊4k�s6���<���g]ʑ ��ǂ��s�%@٫]�Ku���׸(�]9S��R�Ѓtb�ɨ��wȀ<�����7����"Ǚ2��YyB�����t�fp�#�,�h�{V�R�Ԕ��X;�,@���1�o0B�TϮff�W ���S�
���rM��xw�#mQ�c��f&��w�)Xv�_������ ��b�u-�K�֣|��1t3�_[�O��j� 5ʷ�盽)Tt�L�;�qon,������wd�6�x�E&��!�z<��]���2�q��<��ں���>�~%"�ʕGmTc�X����Ym�AA`6�PD]]eV1E�\B頮4�LJ�"�������1��E%����V*�1�eF���9jf����TLI*-j��N�P�Ԯ�j���5*��i��%TUAj]%���\��b2,Ef#��#-���ƍed�1r�)S)A�����+`̹�q1Ʋ�`�)�.P���V�5�Um1���WL��5���R(*�R�0TFѥƎ�& �BQ*[m��C.8�e�*(����Qcl�T\�V%j�bX����E++2�V���MZ*�Ƃ����*,S)U��[P�VE1]%Ģ-E	SV���1+m30b��ť��cQ"�J��Q1���"1U�"k���6�+
�kE(Ĉ�T"&5ӘT���m�D�,U4��KK�\�IB�V
(1X�����kδt}���6c�e#���Y}S"��-ⵊ>��P����P���ʒi��u��VĤ��s������'����j~m�32�ڕu�y��*
/�v>�ί%�Hܞ��9'������J»ש�4��ך�y�8*�$l4::�^D�'�/.ES���w*f�l�}X���k��T�S�׎-sتl�;��&QwJ����R�s=#���u;	���������O�<���=��E:V��:{On;yrKz�����v�Ÿ�Gw>\
�U�:����S]=�+y�-zҞ/7N�B`���<�������7��3/��<��FLmM���u��NVD��;�oZĦ�}M��/,ي3�F�Jm���,Ff�'TS�k����PmV[�]��-];&*��i83t���ze��q龑��}aKv.�{�i���������L'Y��*�]��)�>��l��هLwBl�n��/]���_sHޑ*��#�(���k���y��+5`r;�����!�r�x3�L�imgZ����#�t �V1�ʯs��?�}_i3�a�A[��q|>ݐjy}^���ߌ{��hx��z�ztkcxE�K��ן�>m�a|#l�N�*���X��rͼQa-���)X���51
��a��W����%�R�U�C�f���z��N�+*��p��6(P;��XO��&����9�r�E5�˚ٛLE����R�B�Zf���U,ws��d�v"��/.6�q^�d��\�7��s����\����G�Q��쵪�{s���%�E\d�bb<%����fsZ�{&'T�u�u>.�*����'�bV#'��4�JgyNk��;�z�WEu5��fwc���V�X94��-� �G_U���k��c��d��fyU�2��;��� �)�����NU�C#�+	)3/��Z����O)�V
D�ԩu�ƅR�Y�Cuɖ���Zy��^��K�c�X��n+�Z���kg#-�QeϦ_Bsi�̧�s�V9�yk���z��{׹}�=w��(��&�������$o���K����go�7ڵ)���0N�
a��b���]X�L0(A�d5��ki��)^�
�Y+àtS�V�:n2��;�v
���u�i�6�k�P��/��MY�$�&�T7y|����y����JFB�a�gdOL������
DZ|�1�k���'Zz\ئ�E	L�B	ł4���K��Q��DK�iL^\ͅ\a!��?v($� ד0p4O)�b[oyuGQ��b]Ht۱�� ���vi��e�F��0�t���Υ%��ۈ)���ֺ�t�����n9�I�TdBj+���u�iCh��T8)]������u_b��w��[�9]ũ}�6�ݹ��@��)_�&E7"�Rs�Z������o6�܃�š�`���c���Nj���H5Jn��)�>�FCu�C4;ϸ�PI�}Wol���{�ݮ��i����M����Wr��)(������­k�+9����{Q! �G˟7���R��vw�xx����ObԬ94�r߽�WAf�Pk9�ߧ&}Hn��\M8�ηwk�/&�x0��[f��::���|�M^����[-]�oS}���d���hυ�U�]=ըOm�H˫ͤ�^��=�/Ч�O ��)���v�%.�ǵo$]�2�6\�;�E_f��73��2A |*7�S���t�U�3�،��zn1dCV���毘�¾�3��`���ձ��t��N#�,�V�7g��gZ��[P�/˅�r�X;ٸ�FM9��]Ջ3����<��sJ�n���HϐQ�G8��5��˧ܹ�Q6�:f�}M�J�"7`8�Ӹ���%�\���QO��T��F��F��c&�Xޙ�*;�q�#D:��3���Z�9�I��-��֥�
���+��4� �&�g_}(���Zjv
�d=�R��ۭfbc�bXR<f[�u×p9ŵ���Ժ;���$f["��'��n��9CSɗj͇ۭn ���Q��_�磌�w>p\�#��#c�"�o}!�;Yp��8��ܚ��N�33�]RÙŎ̃>�Y{�kQ.WT7����r�%y�3v��v���\H݆�9sO���ھ2�����qt{qk����/7�:�A�^�t���Ǵ����˜
+nۣ<U�ȸ��{=�n�x��b�U/�cfGS�J�ּոt7j�3`�}���{/��� ����L��H���z���x�tb��9�ӵ]�#5q��(;��(c�'Չ�v�_%�x��3ǃ�Ű������QJ����xyHl��g�5��1��;)Iz�^�uÕ�Kܞ]�*�ma���7�hh��hz;OUOLwmJ���yr�m&3\���z��cO��S(L���Sh���}���.\Ot1��Z5���|,vVH%�w-j��.6^��̻��,HNE׶��\���kn���I��
u��S�oK��pI��mK�����֐�J(���n��qB���N����P��"`-��g�K2{�w+�{��	���'��q���U*��uL4�����\=[��v#2�����0�uG�5��D��Y�j�*ɱJH��*���:�8+u��w9 N�,Gc���jER/��]�cn��|�^o5z�!: `�:,�"�R/�p����;���2�Ow{���gU��y��e�h��񩾐ܦ&�ٵ8"X�\��/��6��1�\�Rw-�!�d,.G	�3X�����9pc�%�-�����<519<5�D���Em�B��j��tֽǦ{ȥΆ\�Ym�Y��hjO�������8�PphG^��[΁Lbͨ�;k(�>�ƅ&w����c���cx�T�C�SP�,T4tz�UM̊ok�<&�ԏ*���Y�
���L��6x�!��F&N郴4q��1�^�fwK���+��9כƗ�xB�A^���S�fDͺ�s�׽�l+��������&',͔{:W0I�L��aN���3z�rc�C��7�:�t�^���_}�}�e���f��Ge}�^��<��	ٌ������;;�ջo��j�8N9���Ñ���BQ����x�q�h>�wܟqZ��z��|��jB�T:ך�!n�� �C���Bb�;��6�rNMUu?�:�сn����${�*Qg�#�Pz���i����WB=ׯюk���Z'�����o+�	*��i�t5	ɹ���V͇�� ��G���H����D%y�
�ۻp��M�-��ũ~�0g�b7���A��Z�}���O�-S��6��}ՏѴ���'p��X�#�Ԩ{Ru�c�v4J�n���s�[��ͥ�#RvT�I��L�B�UYw�����֓1�B�^��V!Kcy����pe�g�1\mT��kOFQ�r�Z��aOx�xk��م�,���t�DAqo�\��ϯ�ݢ���=鬏[ojt*�We坬ai��!��0�����|H;F��NCu����=���_m��jN�va*#fP.g>�*��V�tg�S�]�B��M�%#��}����A;����F���x߲`;m�(h�|��N��pyM��=��nw�'��������ӳ���5!��t��r��m����&:�k�+6�G9wQh��w�:��ي���W@]Sw��E�b��N)�*�*Iq{g2�U?g^$��|���)FF
nj�B'6�D(�ۍ6��R��T�ag2�|������ܻ]`�K�5�.G�Q�jS{uB�81��>3ծ�6u�'��;�)C}|���zuv����Q�cd
L�$w��P���mY��3���a�ľ�S͝�㻊#0��#���}oK��z�v�W�')�楔����ls�h �~�@��:}��u������wn�ؼ�=�h�{�jq?I�8�q��y3�zkg�5����sA�>��7�{�����RO4�4��k|��_��hI,=9��x��[�F�L{������Rev,]�B�2Txt�]�9S�Uv���4��;��=��o�w�c�J�/��H�u4.��̿+a�G.!��T�w�p��n/WU�\�\���9ޥ^k�a���ֺ�JWKa�a�F�"�~Ċ�Uԫ�����eo���J�Y�WJ���j@�.D�|xd�%>oL�0�t'*��cC:m���*Nb+��h��8�.�r�`�Po7%�}\�J��{���<�"F?�<�\C���N�E\��W��C���A��ˍ�֣qD�oF�_��06��E)�E�Զ���[���VN'Ѣ�1�n{]M,{Mf\ߟ�0.̝��/�r��7J��%�q<� U�+2/�%��r�2ݫNi������E�Ԩ�u�"�	��g5#�T�k׭ͪ܈�*5�lʆ�`�(X��!�8����ڹ}��=s�fؘR�4lb��.j�u�q4�\1k䵗��L�/�S���6�����;W��Yt�>�VT|�����&�i�����S���'vk��U��W^/� {�S�|Se��(�U��>��W;3��"��	��ԕօ���v�oN�9��v�k�	'� m�'�1Ȥ6�����Yk�[�kCʹ��Թt��3���<�ŦZ��=�7S��7��E�ݾ~.	h�����)O>8��n�
 ��L�3@�v�.��}��V^�}���D}���ʢ�ꎰ���r�^��]j�s|�tT|.`t��_��Q�]+}iVMҒ6�/ҊV���c*������}P��R)m�U	�u,c� N\1X/y��0���!���Q�\�Ƣ�2�v"rl�!z=l�/(�z�:MZ��$�zS2��7���	�����m������w,�Sɍ�N����9���:"��@�ᦌ�R�)�Ǟ~K����NJZ�;��3�-�8�f��Z��u�Yۇ��Wg=d$%�
.o�r7l�]$N�w+u�6	��Q�1)�f��@fh�6{2b���78]i�+UחN�Rx��y9��j��+{��s�;�V�X�)|�h�i�nm��!r��r~s�3���]���;bKǆ�N�e^�29�y)Y������
���t�nؔ1^f��KT�@pvv��U].	-[|����0��Du*�WY�h|l�>��kDw�\�RJg@Y+��U�Qsb5�r*E�T�Ճy�
�Ӳ�r����[�J�G���ժ�!�m-�3:�:ҕ��_']v5 ��4�R�%���h�K�Ч\м�T���˗�:`7�n�k䏖p�w�yB�kT�]��wcv�8�j�.�*'hat�u�L;�Z�Tr�m(�ڗ�3���B����z+YY!�j��:l[�OIJ��&�ڱqVa�+����$���svؑu ��X�[ƠBI�t������8����wYְДG �9�MC�i�!p�dEK�+gt�N��hi�p�(m&�}����QӇ^��:b۶�L�Ҍ8'�&�ԸQ�׆��C�)�����Dj9b��]����o̪k���'���=����q]���//Q<tLgː� _�A�>s�!��PŽ_��wV1�*u���H3��������q��N�r�:�*���-O,�M�Z'E9��.�G�R��ɷn>�*^�U�m��{z��0ț�LD�FY72��g�y���Q�� ���T�`�h%��C�J����k.މ*:g 7j�ʅ�5l�Zɑա*i�Rѕ���"f1�'�*֝.���p["�1f����l�%*&��a�ZT0^ n�E�|������ӳXӫ�R�<鎌q_ٛ�m�ۋ���*m��Q
#���/P�\e�T·�ٕ��%��יX�Y5��h&�R��\�,;Z�y�k7C�F"��ȰQ���r���9[7���f�Fѡ[)H�^�(0�u5���z�c�c�m^�$��l�u]Bؘ�v� a�5��{h�IٵJ��軭����bl�>�vtSr��mR���nX]��
$��3����`��w�Ѹ��IM�ɏ��R9C��ǭ�:���n�d���|"��;��Y����nU����C���M�ӷ-t�3qN݋�)݀�Y��Q�-Υ�`�A>$��>��0(�AE��*�TR,�kb*��m�B��J�UETDml�)�q�dĳ%���b4aQ��	�,���V�Īۤ�U����,���
0��U+)[% ����c�1XbQU�b-j�Jի�EV�"��bi�uUA�TQEDMS�)�V,QE��t��Cm%t���V�*�mTr�X��Q��(E����4R��[+�b`������1�ЕXj�j�(Hi�J�̪�1"����U`���I�2��c-�R��E���A)G.��SLF��m�Ʋ�n&:�(�YB�((�����B�p���ȉ�V�EF1�X����$U*,�PYY�麥�U�]f)��Fi�2�r�V)-,�Z�QB�Q	*�U�@��h�m�LC2��
�ji���L.JT�X(F�$+���0�����Yj���z��ޮLh,i���6��
=�G}��j+˸Q&����;T�w+I_�����ל����@j�����Ŏ�15��]��Ǻ��Sf�W4��lͧ��n�W'C.P���r�s6zi�̝�"��Z�0�U�%�wv�Fl���r�^4(^bf��b��K�V�L�y�v�/�\+[�t�sM�G�n�R5�Ȋ ��݃�5��{P�9����kM���b%�����l��z'�=��5wV����s6��i�p�b[Ad�~��ͻᵗ�^�/<��ս6����ֳ|��Rr��mwG:h�T�tOSI,���
S���u��3�TegNW�2�6v�b-����D/bb;̵=�yt�Wz,V�9d�ʖ��������N�>�B��}�>��(o��T�����=�����m���ȝ��V�B8�U���#3O;�[���C�W�Be\T(��������e����k�$���v���M�Wn�zu&�Lw�+Xޫ�BwBj���U�Z�!�o�5���e]�W 9��]�y�e܎�yӎ���^^�ϳ���bk�}_U|=v�%�[���o;庲e'P9��#����:�Z�U� Cm⅕J���v)�ms]7	��d!��vD���r#wLη�ʢ��l$�ne�2#[a�i�Bg��qe.ͳx��=���kn�ϣ�9Ub�b@����h�����5�d�+��S�z&���FriRoACx8���vVՉ���N�����*�D�~�f*��Ȭv�\9�lWd��3k&���v��s��Xd%w���Ű�e+���ٳ��2�iQ�X���O\Z+.��U/浻s~j�x�+x���}��mz_��C�^�an?9���f֋�̅\���ϖn{rᤷD��m�Q�3{���\�TK�!�O��p^.4:��N���O��qAU��;:���{n�Ru�2���B�g#^]R�$�n&1 �����Q�A�%��(�����&�a#���i.��,v���B�yW4s��I{2>�\�\��j�x{�{ѷ�ړ�Fc>����f�=����2�x��,MD���KrQYUň�^_�
xP�T�W�\�%N�UMV�!.�q��w5v�<���2�S�0@;h�4��N�E�ӽD�m�]�1l���j�[
�8���&h�Ml�3�,[�N+#7R�K5*{��]�v��xWr��K�e�/!�#���n�Y��n�m�Sw���@gR�n+%8����:��6b����;��=F��]��qT�U=�k�*�I��������Xh�����-5�j(N�-�s����,��O�dϩ�ޜ�(���.�Mꌮ|��}���3 !���x���t�`,s�iF���ˤ����ƍ�9��hX�+c8�`j�J�z����hJ�f}o6�'c_����rq�5(86{^����S	�k1�w�9��;������ru�᧮=:�����ھ���C���]M���o��펝��Z]�v�;CzwbT'6W,'tN��5]ڥn�_x{�����kG^R<�.8nj����9sO��;5��-Æ�SU
7v��sJ]��S�=�ŋ���`�U+o�̹�����9�mɸnƦ��?R�r��413�Ou*��)g�c4JqW%EK�ŝ.'���Sc��N���3��i�b��6s�"�Nݜuw�7���/��	ы�'������OǸ��!�d����9g�J=Fkak.�8r;2���q����"�wW�Pc��a��wKK����<���Au �(B�vn�]������N����K�A�s���L;ʕº�gFa�įx{<SOs����%li� �޿L�����O*�Kj�d�}p��㷞�L�*k5��X?2���ٯ���ڮqj�N亗�YL�m�y�5�H��`%��it��Zv����Jx*]�IH{n�s����#=�J��峍\w��1�F:��i��慖���"U:��G�i�Z�Ԧh�ҧp�6R�f����w�m��͞-\3��}� ���rUN������#�P��B!�j�'=6�䒫�q��O-�c*�5��S� W��Ӣ�L��J��/�z�����s��H�lgi���b�y8��7���S���ҕ��8�˙6��ÖɁ����˃-3+�+%���-(�����F_�a�<������rxk����|:z�8�gb����
νqW�WI�˔(^cb�=n�����]���O�����̋!4�P�m���ʹs�ƆRgG['�(n����1��->�y~Kj(7��8�d������z�����p���t�s�����d�}{ol�����2[�]�s�;k�;}x���͎ƾ9��Uˣho��q��Y]L��d�.jԈ���n�E��F`�����2�l���+��74'��h�?zc���I����/3�v��l��
8�貤�*T<��Ө3`�P�F����W�Pj�n��L	��e����_a.�/]P�T� b`��j�6�kHNr¯�X����+���˔�}�����o��uל>2��0+��O����k���Ҝ����\���u��C_
����|f�uQ��)9ӏr����u��^^{S��J�&&p�ZE��SU���r��qz+k:!0�%ߋΆ�y�y���O�.��p���x�+���j����q�%ަ�y�y�7��e)��� ?`F�� �-U4,�rB�+_f�b���36b���қ�w�h��a�guvK�&/6oyAJ�ڃ�}��T��1���sa�q��@�Ƣ��o8;�T	��AOP�
Ccw��NĴn3�A����ۨD<(��E\�{WM�!	jc�TI}^��u��ꐻ��q�3�Lu�;�"&���S��[c��jh$�w��=a�L�aG�d���mfVk&���v�!-���.�v�ih��٧�r��y�e����|hn%mJo[���WU����p��nb�N�R��:�Y�����<]�ͦ"��{���fl��R�c�EHY���J�\�+*�g�u۱ָ1����U+浻r�o�x���x�d�1źiI�ܞ8�Շ�;�+5���7��z�>܅|�IL[�5�]T�gt,�����Ȧ6Esi�����F5���|���3Q��.Q��%�c��J�F��>��PČۥC�OE��\i���p��'����w�L���X��#\������n��$7bvZQ՚�m������!^ƙ�$g�зo�h�����-���>N$:�Ҽ��r����VG^P�&h��"����O����AV��#8�����l��2����ų�^OtT�+���knn��e���*��[ҹ�Y7I�
���2�iؘ�Fr����{b���;�G�$�a��}�����Z1oeE��=�ͼ&V���ݠ���M���f�������a.��P1X�Ž[ �Dv�O��Df�4���Q��>��qH���&0_n�еU*�}� �"-4ѧO���1���p��]=eRÂ5*nl,5kn�˜H�zi�l]7�ֲzJ���{D>�F���O�����%ܩ}9�������|+�dϾ_��N,��w���:R�%Qٌ�v���aZn���AN�y�2e_�s�*� G:�Q��s���ŵ��\��������1��ی!��.\�yLT�cʺ�VX�V��]��<i]N��]��=Q7�n���ŕQnk�U�x��Ύ��M�Z�ozv.�Q*��+Y�0S_�=o8��hM�&ljFU9y[�=���ۤ�<�7�����|�JS-X���>���rE�6��g���=�gG�~���ܠN(:k�6����4���w�M�߿!2�:�0.�Š�'+��f��h���X�7�i0���ent�)�Q[���]B��^��;�t\6��-�rԽᱬ�P�a]��-}W{A�\�n>�䫎����r���_|\cgVN���0��ܻy_߯x{�˷�m�yy������v��B��GL���;F-�p�	��)E�[����F�>����v�3)7G�];����Ex�5�z�*U��蜗
=0��]my�XpTX���}Z�uX8ς��rUd��cLxW���R7\kY���\Ӛ(ફF㮷QM��ʈ~~��#I�eDoǗ��#��ib�!��GeQ�xG���F�-��̧�;6����P"�@dMwƹV�`�[�.Z$����|��ygy36�SI(O�բ�$�\�C�%��;����F��[JZ���l�"�Q;��l-�E��ƅh�dL�T2�,�'X��a��L�&`I`�I徦�7�W	듳|(�ﳒ4�qy`'"/y�
�u��fcU3Vg���7{�Տ{����zvx��]t���p�z�1l���499������hs<@�g��۴��"�Ɯ7����,Ѻr�mĔ2,��M{�e�;��g;eV�z�<�Vm{�'��`SX�K�8��\C�����3��ށ}�-�����jmN��%���mYk$��K�r+r���ݸ�K� {�G�D�jk�4yz2wV����~��=�yRr�1%��S�	L�Q�ؘ�$��@{+=}Vbο4��L0?{��~��d�.��$Y�`%�fo�֕}$������f�u�c���
�ܤ�~�J��WB=q�C����G8�a�"�ɱ�;U��ڪǛ��YrKaA"�mI��O[�۪,�N�m�#��QEW��GdK�Aͫ�t��%X`��|�gCľ�>LF�P����+5�#h\�����,���2��:��TF���rp������w���Z89��E�ĺ�J��*���SX
��/�o�z{�y�v�q�s��<�)'�'T3���hz�R7.mC�F�܊9VJ�]�dw7ة�Ǫ���>��o�G����U��(Q��|�����g��n�$�j����4��9�A�4vҦv�-��"��� p�D=�	��{_16�Un�-�ۊ^�f��zT�4tҁm+�2��3�&a�B6#}��X�q!t1]w�*�+��=N��|��T�YFZB�)���I+9r�7���%#]�nl����{|��pֲ��.wZdPqR�l��r.�a�f�u�0L(�飜��{�x��dg���A��և^iD��X�j*�і��s��fY1��r�
9o�̥�X7� q.�1`M��/:�u�uV���E:h�/+3���&XmH�[|�B�t�ΏFrMaf��$��ČQuI+)�<uVW΂��Y�5xb�9o.kS�"�,�˱T �0�Z�-�u ����8@�Һ��9]�R���^k�x�j��ݹ-bu4Ѕ/���pv���;{�5�i[#�7ȷ)�ӊ�j�2y�a��c]��!A��ݩ��Ue���d�w�ʽ&ӹC�9�q,����2����K
V����j��V�)Б�͌��A�F��3�a9�%gζ,tⶡ뺼�V%\{G/�U%��]]��aHw�����X�vq��$�[ް4�p�4��c��JS���w%]i*�������΍A�3����(�9ٜ�� %��[˽�ޞ�p���w�ت�q��xH�aj�!M�Gl�:^7Q�8�f�����t���v�̓pDo�N����w���Z�f�m�y]ǩ	][�v?����N��8;)r�]����Λ�2��t�z�	�67[0�]|��S�gq9G��w(�z�xGv�t@MO����2�kV�sM��j���'s2�Ϡ��(�s�]��3���g=W�#���بB���9K��Zev�zvj�2ܙ�u�e�9îP�S
aօ��z��q�^>˜s7��r���њ;l�	�i�%�r��H����Z�ީ[�V���͝�����
v��:��	t��f4�k|���s����� ��۸�E�ǮuoC/����D��sp���i6ު�Ɨ�t+Cl�]@(��s]o]�}i�g����o!����ծ�>��ِLo> \_<J*�puv��������|���yɺκ|�ogl��[!z�M��\��S&ʊζ���sxRw���i9x,b�	��I��I*����?�(.U��X�������a�$\ܐ�L�ʆc�V<DG�r��sr�i)�v��2E�[�k�_!a��,�k{,hز�@�i�9�ilw`�J�����ԩ���y��-}ݏ��N{o1gj݇��Bq�kR�P��iGA޽�Zv��w3F���꽼���y���z�߽���Fx�����Է2Wlm���U�)��`֫K�Y��14����B��P\j�����EVѥDt�"",��E��X�*�PDJ�`��H�Vж�Dea��MI���Zܸ�T�Q���T��X�fZ�X��(��V۫GT�����j*��Q�P��#h�"�JR��m�)��Nfc�)mTR�m)kr�Pi�\Kc@kt�am؉X[ejR�eUb��F�TU]f8TZ#��fFڶ4R��F[K-m��Z��j�EU��ih-J�m�ZP�6�E
�G0�j[XP�l�`���KB���4��h���m�)�-.�*F��E-���SI�,��meU*�УR��ʎ(��)Kk
��iE
ыZʈ������խ���7�OI�}^�����N�aL�0�o���VP��wU*�������`{(�"\�<�_�������o7��m�&����f�ђ�7#b7ҕ2&ê�i�{b�3)s�{�)������{V�/!��"D�0h��M�d�*)�}ɋ�\��7�Ou�Y=��{A#P=�	�V���N�TW����&|=�ue��P㝩���kv�y��"�'$�y��l:�88eR.�*�QS���|=�:�m�չh+D�aܒ�eTQ��lCP(��Y
�"8n���O*�y<�г�m�$�&�0"��FP�,��UV9͎nx�Á@�`�c�z�vҫ¹�f��+����n[����^��N�KU�4�*�[�[�4��61wPٰ�a
��3��{
�ԩ!�_���YU���<m�FC$���/�+���c�C8hJV��[�=����}]-���R6ΉKFu=<Ooּ<K�Ln�hk2�k΅��-R�a���Ã�,�eP�W)R��Gh�_����.'�x��!�v^��g@�����`�Gۮ�Ås�6��Ә�ZЌ��f	��s�l�������S��5�2'�uΛwz3��G�-X��gD����ՐM�s�z������S���<�s�I��E�ǚ؆R��s�~��꯾P���0����?��HV���\\�[�*(��D��i�q#��oqӃY��ءM�����Fm�z��U���/�FY�#A%�Ul��nE,��5�sԘ5U��6 q�]C���#����������ȜR������]�����^j}��"|�X����xv�E�6��4�ݲR��T���;�9�m�l�uV*#���F�L��*,S�P?E�f�s.�+�>*}���iB��NU�Bl�t(�"�p�(�����:/�À���Q��S�<���/L>K�1!�7a�v��8��Y&[�b�!���D�P"�)^C�*5���X��yLB�%('��W�+�:����V6%�������'��L��"�r���!��چ/�Zs�����=�l ��ؾ��|�ܽ���y(9�%�~��+���Pv瓧���P�6#&�#��71c�̷�- q�xQO�����z��W[�<�=v�˻~-r�0�����ֆ�y���oN��[�t͜\$��ڐ�ҭH��7�*u�B��-"lKs��ַDdܰc�
�Q2�W燀��X���������Q��S6tշZl�@���,�: ��ݛIVY��J��հo'�o���5`ϊP͝"T`#&&���l��/��˃.��4�}��*\Ud_��t�璫:^�fPwXi���2��6iS<|�S�,�Yky]խ��v��E�U�կk&��~�,�A����@[����S����r�K��)(�R���Q�H��؛�\b���#��p��amgWg4U��v�d)50F��28�Npd#��j(�Ɣ�"��C�.""*�G)+ҋ"��<\X2�5�UB�$��/Q��΢T�q#�^�V����x9SA�%�!b�|#�p��
�u��l�ɒ�y�m>��O2���3Pީ�������*N��\nT�.Y������fWEͫkov�Tk:Uzz���I�w�ΙJ� ����R��T"Љ���^�m��'�E�Z�gf��tN̝�&��}.sTY��^�I���ú��B*�$7��i����{X��B�G�{�k=�^-4���G{�dUc/��eGyeQ\\9�9��^��f�׶&�<��;J���*N�$���ﾪ��ϓ����#�hr�8�%����e	G|��l"럁\�4�!�h[L���!qrNX��L��e�i���Ӟ4�q��	Ȉ�����a�ٜ3(���沨��j7zy(1�`� A��0g���ʦ^�,E-�"BbE����]���W.v���:P�oB� \�o��fɂ��x��b���=��<�]��d���ns ˬ�G�����jq����~Q���3mPˉ,�����(WM��7���o�[V�����C����I��uY��
��ȗna��F��t��mV���0��t�l��»���G8�o�a͘�U�x�`�X���~ j��V�����[}E�BF<ۄ�{wT�����	�]�C�wd�UcAi�K�f=��T6�򉍩�%����T���=�L����Gzz��:e�k1YeiCb^^F�2��P�4��:P�L�F�n��*�[r�~t�ݚ�!+�i{�	ug���m/��}����c�:�(\T�%VF�3x�F���%t��t����y�V%��Y� �=|�[+	D��x�� G2J��]wl5�m�'�C�.�t�z�5�)ή`�[o�����~�����|�G����g��+I��G�H���g&z���Q���x���+��w����"j����ϝm��'�+���G<WEL+�d/H��@؟�h���d�>�Y��5��W������R�6���۫2.fC���/N9�.�2��{�@k�Fz����E�p�#MCUn%U��:�"�:F(93߽��K�=9���\⻬�D�4�Z(ٰ��g��Ud���1���=
��󆨊��L���ѵ�p#ޤ�e��-R�@!�
���;tl%܃>�Ň���)��Y*�J�y�������\K��>��>&���TU<vkƋ-ō%	���2�M��i)T�;vN1�3�<I���j �Y���:Ph�_���T��2�`�p2ǻ�w�zژ�E�gJ���wo�8؊	�c��{�`�C�t��fL<Q�'s���{��V�����X*�.��f�}>5���X�s��N�6�f�C9# �\ ��m:�
D1Khԡ��+�0�w��[����%A�V@E_'����:�/`9���� ����E�}��޽o�9��¶�v
�3)�i���K���1��gf�\z��fr�7��P�� ��(���?���ﾪ��}��n�ə1�~ ۤAbU�@׆F�fī����w��50���x�Bq�ޝ�#2��"�D�8WeV�5lO�, �����G�=�ֳAͅ^zlP΢}�M'�^�W���4�7C� Z��l3�О5�N!\Gp(��t��ko��^�l��E��=APː�B����3�FN\Ow<���w�jO���kz�?j�l�)�[\Q�.�a��1P�F}p@�#d k�i�7V5����|��m����T�;Jm�8Պ�->�8)7|e�F9��Y(5y0f/���[Fv�]�%�YU��OJ�k��Uټ���w:���a�j��]h���YX�u���"ƈ���g��_ �8�Q9)[��Ɨ���eQ�n�nRS�7����w9Z�D䎈ch�*�8I������TX���,mob�w;�=}M��Է�w�+�,��K0�����F���q^�"$
����lm�O�Lx�d�z)]�иr��0E��F���ͳ)3�R�̗���`����8e}�zuM@5�4K�����}������P�ON��Hߏ[��E:�=5pP*N�ZImq�7}׹gbP�T���I-�k�J�劤:�|V�����\�Rzm��<l����3�R�N�Z�c<�Hu�od+8g��s�9��s���<Y!GOB�=p����ќ3�Q��8{E�y&�,�f�o����b��מUoc*�����\�����p�[�d��K��t�����Λ;s6]vR:r\��۪`ٲ���Wk�k]�Y%?aW����y�N�Ϸ��yKG�eOL�F�m֛R���,�~��=^�-T{)E[�����H7W������q�A�E\��^
��V����.�xQq�ۑ��)�jT��ʮGbgϻ)~��s�S����Em�	H�,m
z�����Uu�J}�0%��?d\�q�yh�3��9�a�6���b�����`��`�q�rU,���O9�{�F֏��+�~�H�)F޺�#z�Q"wz��7E�:�GȎ�z��ЩD׭�+]����x�<0;�U����xQ���#��^ͽ�=m�p� �'��/6F_�����tۇMO�iV�y�&R�7���ggNaf���Qi��R\���^�z���lZ�˺��Yf�\����D��Gm�p9�ܣ1����Yݫ��B���T=��5I�D�Ȅ��4F�0�����7M$F�
���XW�wL�9��uo7*�L?�L���[u�X\8�������JL�&�D�r���wUb6��U{�Z�P"�����H�9$O:�
8�pɌRn��K��\�����ˀ����M��j$�:��2~�oA��T�r(T��yM�6�d�Iz��!$����6�D�6��a��L�)3�NF^*O+qJ��f��=;�N9��Ӌ�3Gc�1!!��4gÅ%��z*U��hD�%,o���S�0f��q.�,E($jbD�N��ކ�Ə8n.�\��m�>�G
��}�zoN�Ђߟ�n�N�`�a�븘��T�^�5{��ȭ��CJ�jZ�=���Fd3sD��C.$�殖�H젷oz31=Q�i\"�crx��X] ��Ž�g
Y4g[�+��t^�8�ͳ]�>��%�]�!䐓Ne�8Q���T`�W6���e�x��X��G�v�Rn����um��٤��Y����B�[�����F�"��������+�h�r�5����}{�>���j�\צE���Yyܱ~��{�� ��[o魻�"�� Ex�t�{����v�s�6�w�f��(��I���!���.!ug<��l������L�$a���y��5¥u��V��8�^x�9[�������&�w
\�B#�:�"i�#h\��8�s��=H��S�\M���t���(~�<C"���l`q�մ�����ϗ���&�<��'wԛ:���u]��l����8�p8�^�:	=��t#Jg���9%��Vs6y�nbF�\ޮ4C�Es�No&�ґ��J���T~�(a�	����Q�\�ݮ�8�qN�Y*C��bT��g���"�bC��p�D�
c*�:��r�u,�ۓva�#J��#���{!lT�OD��Eޔ���3l�4�X����*Bŗ�2"D�%L2K�1��qF�qN�!�.��=4�I1W�˾��̛�+���!���(�{3��H���U`d��[�7�塪ɒSv�[��v��J�G��KY4�2��b��o)Vk�c�8�؇���ݨ������u���r{in������h�ߎ�z����`�n�t�PZ42Įl���U�����z[{J'�� �)I�]�j���xx>���i��R4`��5RrLXP�,߸E(v&E�W)5�f���q��v���kjws�r�vP�6��N�`��,�)�9&�1��4t�F�XnF��z�u��71�r1C躍"�,oI.Gm;�6
q��f(y�A����vΔ\\�F�"��f�_����F����9�����;W�vk�����6}�FЮ�2%������l�tv2�W,P����di�UP���i���6j��Qܪ�z*��
vE���4f2p�ʭ4k�О5�6�'E��fE��4#�<�������:��V�u�Ζ�!�BE��/U:��9x����� �����S�<��o�k��b�V,��A�Che�D�>�����{N�o\W�a�&w2�0~��\/��yR�ǣ��~�����Q��"6Bs
'��vo15T.��U�.�FƩ�5�νVH�i���ۮ2��)�9 �0z��.4��W0tI@p�ݍ�]��2�n�Ĭ�=;��ζ�O�v��ԗ��X��:ٌ�A�x45W;�{6�Wd��R�'Yܜ}oz��I�qC���W.�"�*6�]󡌡|�4�i���0�}z�����v�) xv������N�&�L��.��O���*�Q�8٧����K6�C*T,�5�)QE��z�"V�BJs]evEy�	ҙ��3^|P j$+th�����ϥu�����O~�o1��]}Զ�-���[:����S��!2-�����9��@X,黒�fG]�&�4v�d��X��GZ��r�Y�^RH,���o;q_-��:���Woc�3D$̵}��[���e�3���8���;(6T[x�[+�쉾�b�;1U��o����;�m�>���J��W�.j��G��w�E=��/�B�U&�IPe��]..��L�q�},m��Da�Ƹ澫�#t�V_ló,�����Kµ�!�?���56������~ɵ��n]L��3U�H-p�\�h	nc�PcD��F67���h?��<;�݂�c��{ծr�xQz�Y�ҊCXhR��;^�����=v�X[k�֐3�l���2;{��`��r,i;J�̜R͘z�(;8�PKC��qs�㽊�e,}�ҡ��e����J�.lnĻ��z�gi6�?,|�O�M3ۜ��c�R��]���f6��}�!*�.\�(���m�<���Ih�V���
�5�w+��A뽬L�i��	��Wq":.��-�k��
P,!,1wo&�p}$�$Mj�pŚ��r�k#��w�>�ϭ����:6KA��l>�n�d� �\��r=ts��K��VUFw8��$�+�Ѿ@lzM<B��F�-��F�:�K'|UG��cd�>��J���[Z�{�ͨ%�}h�6�J�e�:%���w�%٧�R��ͫ��ӴF3B�`t�U���+WK���ѵiȐӇV���-�S���ǐbi��u��Uڻ��t�ة��^��kÕ�:�f=H�b�z���9VZ�+G%����\�F�J�_��$wÁ=�"D��[�T5맣7q�Ʋ�:�3 u	nG�ݬ�/������b�q]	,���-��Yw�Zbs�ޝ�U�������	OvĈ�����"��Q��s�U��^�ӻ�8 ���bM�go�a6M�Y]Km�6�U�HRZ8��./�o���e�C6hQ�F��|�[��W�.hw����*v��Q7�m�O ǩ�b�9�r�Y*��wcY/'<YG)�R��A-l����v+O)Cp�ۋ�y9G��n.{X��S���=�(WŸ��K�z8��>7B�h`��V�q�hڊ�j�[mmhъj(���̲V�VV�ʭIR���h*�YJ�J�S"P��ʕr��¢��T*�ˬ1���j2�mRҊe̩QJ6�X�QU�*i��-�j��62�b,��2em��4�b���P�m���Mk�n(���1��UR�A�[ŭ���r�Z��Q@p��-J�ҭV�jZ �*"-H��7\��e*jڬ�kK�T֫0��)cm�X�J�ҹi���b�Ҡ��#*�̴�7.�Z�2����U�s&*�G�a�T�kJ��Ts32�T+��i�kJ���+Y*"�8+�+YS.b�E��*�V��,�(�J�Km�ХmFТ�fS%̘!�m�-�[f8�kc)Uek(�b2��iVڰT�R�Qe�aU�\��j�Dĸ�S2��12��w�{��oڼ��K8�b�L4-C������A�ܜ{ܫ������H�=&�;j�H++Iĳ�UBu����#3{�+�t2@����&��*�5�Һ�����m��r��㌣��*��{��ެ+#����L��Í��qhat֋'G��P
�Am�6*7��m-&9���'��l*���9]G��8J�r�\c��"+��,k5���[�C��gB��R�󏌈ƥ� ץK1^b$.��(S�+),��]}�ԓ��w�z�p�鉞�
����$Ϛ�a���1WD�!3�βУ.u߻�+�P�R"�Uзna�RK(�QΔ�b3݊�/Ψ�[ �*9OF��5��&�M�����TE}(ȥ4�X*�662��\ok�(�q���5f���Պ�'�=�Ep��Pz%�����6ı�d1�(��c�w&�����W͓}�㠾�Mb����-u������,շZra����d����_�%��$�J�����霞y�b�~���/0R�b�����PDsm:k����v�y�z�՘U�#�1V��Ҿ�h�K��2�E��m�Hk��W�o�R/���}�}���U���l��z��.�\�k�V5�+�И�HKV�FC����ۧ�W�zC�s���}q%.��޶t�2���.-�g�쳶�Y���2�l�"n9T�LmF<-�ӫV:V�p�3��V�g�E��>~絆�T�-؟�$4���bC�Q?m�wKŒQ"�{�bF�<��1�5�R��t����y�t�+9)���^�7�
;\��f:t�~�
��`�i��ӛ(���"z�S�z�h���*���Yo�(8���B4:Qp!iL�����������4^��鼦�Z��PK�깋]!�s�"_�.��EDw�K7`,ׯ��:'E��3o^u�F�LXPˡp�.��Z-P��D`^�����J�6a㡌�o3�ʭ��,l�Cػ�.D�7QG�n�ȱJ���dف�A���nR�ӝ�����b�kC��K�d
J�=(�X�q�N�8�1@S�c�v�ݾ�n����h��%�K0f�x��FA���Uf��t��v�}�IB��7NVutk���3;\����+Ɋ*�U���#pw{J�Xa�b#�W��NR�0g�3�{]R�i�ٓ�iuJ��������# �Z��e�J�g^����b��a̜�t���+ ,aͫ���*H����y.�u,˪Yz�B�"7c*8������x�����6��#8#��p�B���m*
A�ZO޸�{"\;�̖}�j�T�>&�9��[v�m?j��r6Pu��@|4K=�I�h�9n6�J;���Yyʱk �����v�5��@���jq��#D3*3!�:Fm��o���g!���խ�Md95<p2p��]N��>��N�Fi�Et���8ʋV2�e�W<�x�Ӫ��ca��3��8��͔T_��aH�_)�8=�1C�a���L�^�o��b=J'��MROi�UP�����SQެv�8��R���7k�����m��/6�sK�bc�RZY� `�$����yŸ��;-���%��x�v.nh�2�,�#��W:�J��僪%��3��<M�CA�b;�|���;�o-��t�bYJ�F�b#���iL��niS.le���I�+Ί��b��"��G*���y��,w�O���~�(a���w��c(����];����v�Y
���,{�]��������3��@�h�Ьp��f�0K�}���z��Y9Lz��뱮Pq�s��w�34�s`�T��lq�]:��7�2�<�W��D��ęC,���>k�ZF��q
�/l�'�k1���3���d-��#MGM(*�=�N�����%�B]L����j�<���@c��d�lp�=A�3v����d3���s9Ruw6�-r�؛R�"@�>ԴD �mge�����d�7�[��6�A�B��zE�IL��K����]%R��T^&)g�/�$c���fVT��'��z"J�ڂ�%�{A�x�r]�Ƃ+wZ_��ir���ND��j�e�:	Xmz+�l��*��Q��&җ�� �1�K1�U[1�S��2�P̙�6����p�� wu��:��88GM�oL�R_�N�3��+Ur��2"�w�G��*꘱y7y���7m`��N�*�纝�\��.���Y�Fc'�L铢О5K$�¸�9�ٍ�p ��`\@*͙�7�7�M�(M��u��QŘw�G���������7��H�:�]+2f����s^|�V�:�����I�v��O�ޭ��/�u��g�X͓���&��!@�+���p��LՔ��	��R��׼�n5O����y)X��,��aWH��ٌ�f��BО4-K�Sm�N{w��UjkJ�`%��5����T��5T��p Q�GH�{���'�f���y�g6_��-���6�>[\QP�&���B2"�Qڌ�c*[�y�E��`�Y�ʯ8�Ч�:7��X�t3�Q"�ڳ�mWx���Z^nħ�r�溪P�
, eD���ևT�=+��
�Wf�����#��#�5�^��s���mD����Az�#b$J�T�1�Ƅ�mm�������Uz�;�W��V7/`?wU	5��W.��@��B6"@�,.1�h����������X:��{6bFВ���1�$�-C"�*X=@�^�����|[���y8I�On�܋���|�'���>
���U��L�9�(�K��p�������OB�8����wu�V�~ݑN�ȧ�f�^E��Bu�Fp�S�&��`�*�M��,���~�����%I�3�ق�`����н����`�TMz�.���1��u��"=]�#��sf�tji��Y�Gk���Pk!"oo�����*ݨ��b��S�@x5�����vn���� ����N�lvb��Q��eD�s!��;p��{]I�(g");}��eJ����Zy�Ah��x�>x��A���c)�:X;�D1�(�wO���0�M�������ʷ�ӌ�|�����L�)pT*�IA����G�)k��,8e,��|�ƒr�cT��z�z0>�0C�	fn4�Q��s�4.��J&s�������^��Ћ���#^�;�՝6�L̀��D�
�L�lyz6�(�Z���{���P�J���U��R��`P&�����(���[[���-����X�;A3S�U����Վ���Q��t
7�
e�K53]c0^�'��m�^�Ga��s���jd�5=��_�K�7⎙�B��V<{Kw���5qfTΑ̍�����(��ej�P�DI���/�I&�egW612r�Ib�U�":`q�2��Y�'L�J*"�K63*6N��}�G�����6��d�@��8��U�|uc7s�0����ݍ���ўڵ´Qn�26o<h2\)��i�*ݫ���܎��.Ǐ	ܚ1=���fR�/K(�<6JڱkM�W{�'>7Z6Ҡ�FYyHN`�9*Ou��;�rW����	`�԰����~��Ҷ>�����Μd"�\I�D�$l�뒋�O�ʳ-�6NB9��.����QG�����#�n�fz7��R՛�jΤ8GkE?U�� R^�,�[2l'8��E�-�Ut���������"O�ش�c�+�x�B4�ʉ*��N���>�c��l+z�y�=�
�/壁
��/[E�U�Š�O��>����T�E����i�;ә:������	��Z��v$�{�!t�������Yt �S���<�a��r^f���Z(8����DMxs�����ڜ����~Q��Ɛ��y-񭠔�7�jOn-Z�m����P7�,����.�q~{"�	��2�/�<����:~�������n�t]RQ����*2�˥#\#o�a^���br{��nx.��VRb�Z�Bʑ3LP�e7@��b��R�⍎�w�A��	�hV3�0D쬉� �S'Z�.�KJc���-i��W�;�i�up3���w�\�nuN�y�CN���ؔ��ꉖ�>��u�oe�д�5\����V�����"�$�KwP9G�v��
�4�vEN�/�<Y�bF8$l���x�r���uU9�Z��9^d�,B�;��4��mȝ2!N���y�yq>ɠ���v��y��QE�M�$�[#�Q8c��gb((k��uy@D=b��s�š��||���C/BZ��*�L`/��]e�Q3	�&B�������k}���k7�Dd����MS����ׯ�zaĥ���n�ȸe��H坷y�w���K�	1�	�F(Dq�]h^g_0�s�3xQ�t%��i���F�}�-�|z�p+�A]G�H��hA-h��k�~�&
>��gf�B�ί�U�Z��|F���_t���T��K���f�����h�;�ݛ1X��}�d�B���B��A�1�ˈ�!�B+a�ȼ������xbq�xõ��\���`�g\^����\����9K$��1MLDOa��4��8�y+2ӓ��u�o��e��V��AeKZ6k�er��e�����b��{\4�ᓗda0й �ƶ�2~y�n4+5�<�:�پ5�'Wm����[{v/�R�iǫ`J_L̚��o��_}U@l.{������VU��TC9ㅖ+��>��ypr!��2�e�n=�'Wz�zF��:z��;nE�UFl�f�5���Ѷ��\x>�Ե&��7�2��]
�md>G���N��:Gn����v9�تT�rP.������/36f��Ui�:�\�
����7��8O�,�a��
$�7���b��Za�Ζ����g��aU���zn ��1����%����ĥ]���N���J5#�(:�������þ�����f��{��J���*�W�R�g�Eb�˄��(Q�P��Y�~�"ymqEC��htO(d��z�E깺kZ�URd@=A���t��S�����Fu�eY"��a�\e��,�A�NWD��J�&�( ��p�I�Di�v qT�$NP�D��Ot ��۞�͵�;aL?Vʸ�J��O��b.T��G�ËE��Mh���@��i�P��>in݋�!�nv��#W'�Ʊ��k CD̫��4�lT�����gi�gl���]w}�.�������цTo/P�H��H��ɑ�㭫y4OD����rܓ�}��Q�I��ή8~إ�Qv$��$m*
"��3�p���q��O���a�����ۮu\p<x�Ɇ)N�:�؊jY�������u��pkQ��Fg>�z��v�1�P�05R5�v(�,��3�'���W�T����:���"C�;La�9O{4�K:����-�E|����[��;e�X(���"1faV�`��[�ռ��x@~͘:heNs6r���4�+��2��\o�]IN�:�{�i�����H8�n�bܭ�A
�j�3n*R:a�=�,EdY6���J�g2]s��A�^�:��Z�O�0�C��h�d�S6Y��� G9��dC"{7s�uի�P~��!E^Ԫ���{ӏ���wV	f}q�R�#$��A6���>������c�+��0h��,�U^�{L��8^t��
�1qD�����a0(Z�gň�K�{��]:R��DoC6�<�[������mW�3�2%�/]o�n�MN�;��|������Զ���;s��;��f���7t�|M�����<�����o�no��Vk0���
�7wQ����V���en%�'X�qN9��T��;��Ν��l<lRkv<�Ӷ��y�#ltu}z+��fA�6d����ha'@DC�<�eeAq�d�+�n��P�J���o
��7���Ȱ����{g^uc`<�ȅ�����MV���9��r� �аZJe:Tf)�m���Fu#�,��X�P&�v�u(�d���x���3��1Yf.�X-���W��棧�fY�]/W�V�ݞ >��9����/����L�є��;�.��������K�������X����)�yG��/��Kq^��v�;�����q��/ �1��a��x���<���c��ë	/Pֺ�,�'w ��:�w���\��sU�Չ\�V蕔[�tY�6� Pf��g@�(�jC;��9�ZQ��]L��s[�k2�O����b�[V����u�� �]i��;���	����|;�PF ʗ�7F^H�����<+���˟t�`'���C��[˰h�إe\�xuY9N��k �y�v�7� Res�Ո��n���}�JgfAz����*ʜڽq��jy���^�	�M�+�Op寡���9V�h9�%�)�4Q�(L޸�J�墶�nc���<cE���1��ٵ�.�k� '�Mo|*#��7#p(f���<U�w0eإIe��#(��]Ѵ��B��R��nҎP���7�C4iIB:��h�Ģ;\�.�`ն��w`*v�l���R���vf�ԭ�1�ftҢVCb���4X��y�b]\��P�MZX#{��P.�l�@��f\i ��j�7R�eռ4@E}���W�Fa��]${[b�-d��J�V�Mm���A�����HX/ � ���T���ʺ��ˢ
0u�f�J|�1��; ��F!M�܍啔w���x�Ma�9��)e�ydv�놴�\���N���{-f ��2Fȷ>9f������݃a��R���a��=��(��{�1���or��$er�Z���uLA���B��]n��ס�O��/r���(����ŔP�3�9q�YtS��`�����Yg_��v�n��t-�{6T��s�6�;xw����=!s��������U���B��Zf×���s�ʶg5H�\��[Q�V,��af	)�_:��S��V��#��m�H��RԶ�ث�.6�(�ʗ3ۍ�Ub���Tơ�Uk+P�-��Q�1TQ���V�1�V[R�UT��"�eJ
�511�[V��Uq�`�ҥ+Uc���2�
��`bfc�R��TҊK.DSb��ģ1*�+�B�2Ҳ�rڕh�(�5�0�T�31D)E)m�8Z��c�pQ1Ů8����Z���*f\j5�E�ʕ�Z�im�	�aJ�F���D�EY��E�F�FTU�-im�JT�kV��e-m)QaFZPY�qR�T1��,��V�QԨ���+hҲ�J��kU��iT�-�KZ�-2Ҫ�V���Y��2�Z"���κ�2��֎Y���9���
�/+O�q$P:hb�pZ����;�w$Ѵ����j[�xz�v��wÀ�/�����6h_J�F���k�q�s�?⾠B݆ۈzDٿ�"p�E�i)�h�0:��v��F��D��z��P��Ƙ3v��i�t��Vj�c������Ȇ��b��s�S$i��48�Nl��(DW	�b�5Bw��r��ti��,�W�Cb+�#!�g�ҋ�1(�c�����2On���^rC6�8{H9��W1j�\C���
P�'����Q�w+�h���or��i|�ȯDI�Bvx���%W�X-P�A�D/�r�:�����ۛ��בK�p�~�y��5����wS�צx���~��L���
���By+k'�E�8M�^��s@T#Y�d�@d&|��q�p���W����}�ÇB<��z��)H�ANֆ��<p����DA��fr�X�M6�1�r$!�w�[8f(J,�Xa�"��D��l�>�u��M8{�lY�*�cLk�}�õ�pE�C��&��؆�2$�h�:�u�����Y n�t�+�c��j�RĢ�Jd'���M�\�n�:���b�eb�o�k�B�c�t�EP�Օ��(�-䃌
��qwVs�y�R�d+��Rs�p��������D��َ̜Q�p|3kK,��*�����Г���gD3 (̆W���D�O���j�HC�����%�].��
6x%�f[�*�Xf�;S�N��y�{h���дi�к���̈́Tr��/qƃެ#����8��s,o�4_��;��6-�P�`�b��(�s�� G8J��&�t���3�%_���]��إ���~wd頄vEN�"8��ؑ>�$��s�b��+`Ν�[R�U�wH��eu�K��F��)�'IQ�<Q�uH��^�!%K��O�:�dI�4���W�
��U��V%��5��ҬuxCע<�U��	��7t�~�v�yO_�p���X�������=��꺵�eO<G�K����z�9�|_ƅxژ&�\���S���p�{j�41u3�mՙK�,���.Dpͻ�[CfL�`9 � ������YC����	�¬:��a'8���Q@�Ok��5��;�k�n�Z�
mѾJ��!{β,�E�Hh�!I�!�������畊u)&31��Fi�QAZz���Y�a�8AmwdNFj����I�y	���ՀΥ��o=�{�)�����sQ��V������3HF�L�'A`�qǁ��J5m��3�v�
���wT�6�>�µ�nP�ܽ�G��be�B/aؙ�L�0h�:('kZ�}X�t#�d�q^� �&,0�P-D���4!�El;"�N��b�k��ggq�,�F��ƈ��t���0qC$��T�����Xh-�*k��3��g������*�QS�zc>,�C��=��(�)��SR,��5|jy{)��j+�2%�4z�D�/�y�����۾��/=�J⊮���wљ�����Ew�j�4ġ����
cf6ܲ(\�B�/$ k#O3D7m>���W�<���v0k�����N3˺�̀�aDI����
�4jО4-���h�:���D�賬�Z�vC8dcΰ�&�n�=;ra���y��:�����n3r�+/z\GX�E�V@��r�4NS+
�t�j �#0H�l����s������=��Fb�Hۭ� �Tb���H�9WQ�K��:��T�i���uΟl%�v��Z�G^�L��]+��q�ӯ�R&����xւutErU�'M��=���s\���[�;���������﬩���yH�W��hl�\8��9��R���렶8���Lv���Q��A�N�l�=��e��WQ$,@�Lt�Ǧ���\Q��m�둝`j�D�}xu��0C�z��6g8�0ԐY�#A��I��裳�	�]��4��!f]�5ujwsc����X�$>�4.b�6D�T�~�g�F�L�eE�Ϥ��6d��c�v����n��H�LL��l=4���R��*�|����]G	T��*,S�7�k#�t_0���A>��Օ]��0C<��08����lE�A(q��\#�/����I��t`f].wqp�ȉ�H�����=L`�g��2�c2�B��]��HuR��O�&���3�DH��E;�J/ �5 �����7�gE�J����<��Us�?\DpxՏ���ƃ�p)mPf�2� ��*�n�s3˺�<}��C�a�d�Ь[�^�A
�Ơؔ�o�^^�z��11�>�S$�SL�]ʙ���w�syw��b�{}�%�T���824�;a��X���YY-�s����e��Kd���=��py���ݴ���'+�i� �s���D����ٛ����	��>A��%+�#��U}W��y��t������*_+�`l�=�U���벥%��֝�
��SO{y����Z�t<��26(��X�]Ozsϧ�.�,�!qp��+�c��������ﯕ�<��f�.#zp꽋%|��㚥��t�I�����/���ۊ�C^�F��#���FҖx�j�}ۿy��v������[ڎ��:ԙ�ܚ[|�S�č�8&%�1�M!#H�`v�k�oA��*�Ӯ�v�ǥ����,)��6;F��F�T"��0����hW���yP]����L�C��~� F���jg���F�p(�8
��\Y�<��e��	S�/w��/J3��v�I�SS	@���ˈ~!!tGO&v�jq�����p�L_���x�@å�GD��;.Nt���h��됾��H��Rl]7g�݋�K]�Rͨf��g�Bػ8\t�[�8�8dL��&�Z�*B2��=����ɜ&�U�Н�f[��̵�]�x��C-T�9WSY��t��U۾1�T��Y{�Uwv�X���Wtg<����Ҝ"�mvN)��o !�cai�:V2�]�]mvj��/��t��L{����S��ق��B;s��������~�t� 5��M�N�
t���(�ʡ�}}neOsB�;��/�M��,�~�2�-��]r����!C�~���`>�p�b�t���Ch����D1�Y�Xm�8f(J,���Y�DH"MN�2)]qά	��,�Ж�Ri2�����_��S&�*zb�u=U�Z�y�ڨs(��K��K��ik�&�r�����ɢ������[TD�/mn��StC+ޙ���a�Ů����B.c���2�Q��e���ץ�K���E�6�ՙrӍ�S���6�W����
���D�g׳]Q�.WU��8����Ue��8���H��bݾ�zBJl�%Xz���a��p��L�bF��ܠF�f41�"y�tr}��*\]dE/ٶ�#��ȟ;�UQ:w�GdP��(X���bE8$l)7Zo�m��ګ[*"Ν�#���;��#���*4�P�+G	�Q����X7�]=2Z�RF�ٗ�A2���I�7�]f��}L�9��P� ��n�*���;Lo��`�muBn�SS!%��}��B�-�{m����o��Q����-�Jƅ��|���"��y���|��˧q�r�7��#-W��7�[~Ju5���:S�<J�X+�ʥ(�k�\�7/#
�,պ�a�(}�\ �VX�3_Yb�w�JҨ{�֩��͕R��������b�CQ}辛p�z��(N:�U������g�i�ȫ[	U�Wn�/Q��J1>� � �F�]��O*ྩk���at�V
�ͮ���b�����rZ��4�ޙNp��N��!�Dh��`�9�@p��փA�q}�R��μJ֣�U��j�a�X4R�&�)S0k�L�HE�8��)R o�A]�GT\?{ع�瑉�\�����ާWƝ�C@������)ߺf�6����T=�Nh٢�qz"J:Ir:Cw�2H��q�Ȃ����Xn<���%o0$}�*�QS���Q�	��H{��(�N6 <TwW[��l���f*�#n`���K;nE�ʠ�͙�lۆ�Yn��U�uf������P;���=u��<!�l��Hp���[�Z�Q�l�i��w�3��+8��7��N}Wl��xޮ��'g�eI۬ٳ5oz����C�fs+�`�S`�{�Y͡؎-s�S��9�k1<]�\���_�UoF'<x�DI�X�dm�����y�S�/S�R�u�	��G�K]ԖŪ�+ȵ�h=�͌������h�38[�U��Z�r�8���3=ŧee}����2�b���}u���Mu�gKu���T���A��k�����=X�f��+��'�z���_:��FK*�T��'uP�2���KsgZWݪ��	X!Lp4&�Q�}nTB:��v�f��#��s�]l���5�v�u]���--�|}B�$]�C��׈��Nhu�;�2��ͽ�$9n�]DcO��&yn�-��^$yFOK�_!C�����U�]F�?:�[��\����&k�<�&�l����&�P���=q-K0y���lD(c����G�$�/?7;P�޸����tR�Muؓn�MąD QHB��R��1ڜl=�������/��iQc7pR�1�p&�PjYzT�*�z��u�7�^R�hb�z�8��y8�]��ЋR����n�0ŗ�	��LKu���յ|��+���1���;�sVf��ò��O����x����"�2�sK��Ep��(As��{2V�]d���}F �t����v�/e�R����
��9�9x]	^5 ��vE��༘.�}�*���LU蕅�����"�ȥLC�$�����j��֌^'��Ь"�]Q؈���_�ߴ�RY��V�uf�9�����~z�)6�"�f��C�f�%�b���!>ʋ=�f�y(�rʫZm�J�a�坨�J�8h��Yu���Z�|B��U���%fD�͖M��c�ºU�Z��{{t_T�hNmqc 2Ltqt�V7���:p�e�
�K0U��<Vی�[xE�~#&$R�7����E�_�����5�3���Λz������mBMZzM��UCM�cj(�FҖx�J��ަuԢ�͟-���ݺok�9J�;�|Ҷg(K=v8��"(@�Ǚ�����9��J�5;z�+.��qg:elM����r\#�H�@�:X�*�B���H�����"��>t�3������A��-�/6�e6�7n�L�z��<tM��a#omڀ�t#]&F��rk6l���y|Vwj����e��4"�c�L���'�k�}��GvvLƜ�ցlw$%�+��ը�s��Z�J���f�^+c��DBӴ6b��"��n:Qp!A��Ԟ�S5x��w�#�������F�p�W�7�G����8���
|��G�2�8S��^�O?+o�N�|!�7g�f�(�lק��"ױ����(:�
�`�%��<�r�/�}U��[JGqp�\�I���C!��'EM�Bv��-��ְ5��a�V��5�Ҍ���`AvM�B�C�(�B#P�G	",�dUӡQ�������M':l�ř��c����Z@yV-'kC�y?�������ܴ�G`>�q�HzS�-��1��Y����)
A��Bwϛ���7��\��d�CΑ,E($@��	�ʞ��r8P~��]�uZo�~V�{*��7�ϒ�Qg�����x��LV<=S���M���mmnԵL�f��ar<�I[���������mP���Y@�����].�C�p� �v�^��5ڗD8���fbF��tw�$�R������'7���\�.ہ�骟T���T�V� ����m���/1>�+{��$��u	U1���r��1�ThV�B�G:M��s�1\����X���H����q�h��k6�g
Gr�bVG�����P�(
�sq�uIZ�]�io���lŧ��F��A^�EM���Ӽ�������t����#�:��@�^�#XA����B@m�8h
��!�h�(�̷��jC�����2�mPBC�Ҳ���VS��h0jegjRb�hf�(���x�܍��?e��*t��)�ZL}�p�]ϫ.�P�<��V�1�q�����p|V�@��RǕj
Y���,c^�fnsB]!�Rn�̀:Y�����V�;~Ғ�+T��;���-}�F'(���iP�q�v�"�zM�kIA���k{9�&����&��f�m�~c"���2�WN�k��)���,�}au[Nʱжym���Y�J紨��SwDee3�*���d���rgV<y5꽮.�YRv�+�'R�.E
� �$��`������T�@��և�\9�:[���Z��
^|f�ᮬ��X��z�����	e�]V��� �g`s��T�F��ׇ� �X��ζ̮Фg�ګ=��;�"���K��r�������r�e�igmv �(:}o�����/�e1�[/R��}XjKSu)����D���d\s.��JWI���i�B��au��U�(�!PM�:�e��8nE�5�6��� jO.E�� KFV�(C*�PQ�����$y�`u\)^��j�S�Œ����5��O�*�ݒe%Xղ�Uà�`��";v��f�m��i��"�t�B�e*4�N5gV,V��eĶ��iⵕ�::e`��xjp�E���`��U^��@�s���4�/��$c[%�QV��3�,��;�J����ئ]#�赺�퉹� �L�~	��h2�'}7ӕ�������/n��7QǢ���=��^�Y׻J��*�E�;n�7�Eȳ�ܫ�K�Y!V>p��(.��겄��˻�F��[�>�}YJ�S��"����~\�s�>��5�9�����S��o�bZSn�s'lý���o-�;�N[�Gc��I.���x���gm��SΥ(T*���-,�>IfH�C�B���#%
��0�r���x��jE��wP2��:[����1�T��xTv�\��U��ҳe�S��U�;9�7SK���c7����Q|F�J����*�E-�m�UD�Q�Q-Z�Kd�DK+[D�V�T����FҠ�Xڔ�QF�T+*A��+Q,���Tm�%e`�J1��*��T*6�,m��XQ���
�J����r�(��[km�Pqk���J�����[nR�@kJ�֌hܳ�eb�m�,*���X�Ѷ��+*6��mF�,F��E(�PiE��j8¦%�[Kl��)lQJђ���IX.&(�kZ6Ҩ��hUm�Q��U�T��Z4+̠�(�\�eJZ������LcZ,b�Z�L¬Q6Ֆ�r�E���Z��YmV ��)J���UR��q�j��Z��Z�1`��J
��S-%�6(�T��^����3��|��������c�,6u��Ks�)��L��*S�#}P��f4;VdT�2k�b��׊T�.P�T�+3�:�樂oJ�B#p�V3�����.et�<��k�D�'��w9j����Z���v6r�R��}mRO���z�c����&Vxyx�w$N��%g�gU�̭w��x�9����A�ؒ�L�f���DfYƅ7���{3�a.܆Qޞ�T)y�9#0H�f�A���B��g:���M�g/�R7.Y.��MLz�[��qV��%���l��w/e�����xO������^S���U���؀/7��/��Z=�>�������yM�}#O�v'�!}(ׯ��3��B\���W�jH�ֽ1]�љ�T1|�̋�Y�rA$A��`�.�rᐍ��Z�p��������dTo��N�b>���?>���u�p���ք/�Z�J>ś���eES��^�N�؊҈v]U�mK؛�L�b!�d>���m�r͋���vޞ�$pV�w�M��z�wT�`���p�<�#rV;�,����"V�>�q�<D��{��漺;ׂR��D�K(��qX.3כ��[}���1%�ɡU�M;��8�I���[֬�.�4b�;w�s�qI�T�|��������"P��Y0�' �&,4\�B�7&*���7�z���w� XR�X�Z�z�@�
P�ȉ��5�E���D�+��=!��$4b��E�S��arK�12���hu�pxgȸ_���TT��1�	���F�^e�����[���>��<L�U��"<n,)/�ή[u�I�J�����ϋ��knh �ݪz_���K;Fߪ9�\�7���\A��*tչdT1>����qd��Mf.n��Rч��P-Ʒ:^��F��.E��D�9[��'.u4X��Y�b�q�5�wc0��]�$��8��\�jy���3k�;NS���vN����|Ӗy1{f,\�-r�=+��vi��Z6�S<6X��ky=K7��*5��U=J�@�b=A��g��S�����C4o�j���S�\�+M��1�ĳ!�� ��>�����N�uˮ(�q��gRW�ݧ�6.��ptD��[��]�#S��.g�JW����86��i�w#��3"<5���g4N�v����8�}�շ4�tfٸ����]p�\^���u�|;3lAK�u�#������|��h黯7�U�'Ze�(Â6�0dD2L�iꍘhK�aGdZ�og�Wd�_u�qP�:t�D��s)O\M���/ŖDB�z�Iөo��%�[qxX2Yt*YƖ�����)�zS�θ�������v Jx��t������Ⱥ³��)��*,k5��rs@��|�)E׹2 �,���<�DC��Q]ː�/ۃ	OL8�S���'"N�bu��`�*Y�gK���6�;��jb$���"B�5��g(n��P%Epf)%�ь�B�3sZZ�=̒�!��d��B���:����V6%ӔdS�p-ePe4k�{Q�XZn�F)pzp*�
01�TOk�4�������d���m(9�����D�^�]�)"¹�(�0l�.�]X���xεb3+�[�\�����GΚY=���MI�%�u��T�5�(��'z(�Jhf��������]�[��FT�(*K��UM�zve�@j�.�Ӕ-w��k;S���X�	R3B�3�qǺ����w�v�М�\!{%��Ϲ��F��]��
hboGM[����s,�
�Te�qw���&7k��[�)𷛽�׸��a�\~�����Wҁ��(���oS.&}��X�YӰ� ����;و��=��XU�V�9T�鍨����R�x��zYǎ�]H���ˋ��.��wۜ�N�Nbñ,�A賂bP�:E��4�0;q�2�tE���,CR=��8�ԍ�2�&���St\# �9
t�bd92F��T�(\N�*�}\�����b��#���:�
e
��1^�ϐ��"�3�0a�s���Ǝ�Gޙ�<z�Id"�fu>��y1�x9��Gl!2"�:��R�rO4�Q��W���D��j���<R�%ު=����G#�Ͳ�!��|�T$����:�˞7e�5pr��cb�F"z������M4�9��F��SUh���!�֣���	�(!��{ �2,���a͆�n��]˨}����t �������)5���!Y�\Y��*S���ψ�/}��P�m���Ŏ�
���R�ۍAGT�6V`�Ք"V������k4��
�Y��-�p�2�=�r��ǲ�a�Ed'q$ȸ�9ڲ�[���Ng��o���({/vWt�����z�]wr�}`v9�Ą�8�+���B��/�X�!��w���oo;����FU8wbT>����LH��醢2$�3Y�k`d�%כ��&"��i�� _=]�+-1�+�/�CK���	�D
�J�j[�����R���Ez�#�tx*�v|%#��d��#C!�l"�M���w��7�#�2��%\�]E�(���̈́�J�%��N#6���oh}~>W���BW2���c�dL�cd'oͧzF�1<��)5cb\="d
b���@����f�u��i����Q�C�,�V��lS�A˪'Jn#"J
g�;�����H��jsr� ��$��s��qn8����F�t��	�!�n���xVw�"�oE�E�LN�6�Y�
՚cS\�� F����V%��p���ųa��z
�]�T�N��><2�7�/)���)Ֆ-�`L�а*����亍L5��b�oVw7%{���T+'�8쀿�ޡ���h�V�L�+�_Yݻ(���X�c�vC���N���v�U:����ͳn�P��ӳ���(��5?�_Y��Î���t�U�#�a�wG`>�3�[>?JN-�a;����V���*��]/*�'��n<���z�9�=��[2�y��Q�����
� R7d�����^J3S{W0�;�9\�ᗸ�J�*F����*�2����0��1u�p�(f� D�1��g��<�O�fe�����R��2��8:�������!�Cy=����Ƞ A%���X2I��g�p(�""�{��S�̈j��]�x�~���E\;�ȼ�P#+j�E�4D�8���K$��r�U���C)>��������o�VH�_�����Lg�<=OPh�;����aS7�	�4�����G��tK���v�xT�<�Op�9'սO\Z�Q�͔�ʨ�o]oFtٰԋ5���;p�4�ۦD�$;Un�jj+#��ҙ�v1���M�Y��dd�*D�TmX��b���Zˡ���������45��<��䔱�'u���^	;�Y,.E#�`}Mp4ѕ74�݊^t=��r������%i�o��m��
ʀc���f�]Q�n�����vfT'��%��G/� �s4F��;�(�3�ΚN˸�c�[����2���;A��h��O|�|`�Mu�gKu��V+^fǯ�;��U"��)r����瓈V6Yq�EP��t�2���*��gy8��-{}�ܚZH����Ѧ%
S	�QV�Z����X�d�#Hqy����fY�R���8_�ӽ�Zc�$�(@��i��\���Tێ��i�/��Hb��z�/�^���R1NH,�b4�1z�.3r�x>���:Z����T6���NgH}�TH�RT.b�N�M�L��?C�p�K��in\�X�	D�ޛ��n?�������>GG��^����t�(����s���mg;Ni�)"L0++O�⨱�֏2�|�%��p��Z�D�F.���_G+M9*7���Us�)`�֣ſ**�����X�]gLGKem�%��Ǫ\���6��� *�\K���ε	��RV��D��DPw"�^A�p Zվ}<��,��ʊp����}tf��e��R�H4M%/z`�ַ�*��+�KL�T0;W�DN��rT4K�GwT�y����"b.�,;�`u�y�MȖ����&�]��ո�w8�����0'�^v���t��M��,�W~���6d:��)��6�����u����KG���ud@X��XӚ��b���;cV6%�.
����+�u��v��F�Ɇ(t��F�,�q��ʰ�B��Ʊ�6RPr����B�'�w�r��/��0�Y��R�ub��۟_������u�7�	|r�g�f�&9��7GK����}�,��!�x�r5M����>�0c=B������zb1bQ����dĊs����l��7��	ף^S8�Q��6^�W	���GiE����wXi���2�&6��n)g�(Q��t�o-Η��O����;�����Ӗe;�\���^��"�4���#��� ɸ̧ik{��O�Jի��R�&8j_`V'v�	v$G"#
6�n�ۀ�%�FeQ��t��$oJ�G"�HɌ!F�v3��[��k'v�p�3,�<�]��1�F�p�Uz�U7�Fq����fx �K��Uӫ ����q��q���2 F]�.���c�����̯{<-�ۮ�e�ݞ��Q��BK���-�$�t��%G��6��g��4��*�A1�l��.#!�7eKKI!��:8k<.�\��J^������J��3�w(�m��F��{��K��(yx8E�g��Տn�K���K�Exz�j�'�^S�ڼ�P���!�t׏�-p�¯=�7��ul^���1�k��gX���Y�Bu����~��ҡHA� =�A^Sǵ��J"�稱�i�������(+:�~l���0d,2�p�"���m�2�V�[G�=[Y`�{:`Ȥ�ٳ�%���D{u1b��^�51�^Ј��fz+6�&�,��cl�%R⍛2)�q{�E��XP��DJR���9E��7��,��\�_eK����̆ncH�m�b$�7YL�s!
Qhf��F�u��V���qC�a�}i���|:V�<��c6��
��"���-f�"�Ȯ��u�b��9n�#�q|����l�r�=a	����Ӈ0#)�G+�)d�@"n9ى�=�v+�_7j���ܳ*��H.���]1��u4�Y)�=[�|��Q�<K	3f���gIfs�{�ٍd��qzw�Bo��W��;������ͩӕ89f��$�|.��m<Oz����2.s��bU�C��Z���*x�C�����תÜ�'Jz2vh�>w}��WI�n�U7���9Ul�BDӒF���x�s�,�!OR'��k�#��C�nB���n&1�O���c��(6�\<��&
CF�51�k@��+������U�+��%�p9��7T$N�"!�#sҍ����a"̛�}D�S�1���k��U��������Z=+J���(Q��|�	�`���֫Aa׽VM�P;��hb�+^��-QL�F74dP�Y�rA�D=�	��9ي���6/�V����r{W�9t�Q��{�K���L��pb��lD�w��iYh�O�S;���DA�:�:��c]��t6":K��m�Q�6���r,�'��ý��������L� � ��,C��S����*E��
�L\���SO��ê#�À�Bbda�R"k*�E��A��	{����whX*�^>t�S��~��o�u�:��[��U�M�a�	y�����\��Xp��*(MWee9���ar�,�����P����r��#��vSyS����DPw#5���:�ą@4����p��|tuN]�y��\�M2�H�þO�\V�����P�5�j�/��	K�u�)���E5�	�k��#���vAE�`q^� ʫ�cx�ɉf�y'�;dF�"��+��ȟ's�="�gXɷ���+}���ƽ�*T�*v�^�YxS+H�d�V�;��ü�.C�%����5+Z�J�3��qw�ܬ��cV-or\aڷ�9��]m�К�ӴvmjA�嚻'[�5���M,쨀��W.��|�f���gq�:X��c���;V�wuw0ɕ`�V��w&hު��<��[o���*�R5n�ʸ����/���X��+��Ҡ�Ǵ�4�)};hꏅSq!���7k���؇dV*�s[Ɉ���)��c�����Dsx}b ��b:9L�5�vorL,�Zm���"]�y��} ��X�o7QZ��Ц�[�s]czI;{L�L�l�Y�OB��iwd�bІ����y�%�WM����9�k����4CQ�P$#��1_ve�pX���z����Vun�����-�L���"S�ػ�]���٥��F�4q^.�n��J3�i�q��`6���Ҹ�� ��G�W\!��f`i�Xh�M�-݉�fKU�lvU��(p�u��[���Z�+�Ɗ��0��*Usk�A�)�ش^�9kd;|r��tz���D��i���v'���U�;
v���wz�΢5}{�T��lmi�);�ި��[�^�J N:q�A�Qq�W
�ޕ��ژ��PeI������3	$
��Fܻ��o��������	V*���
�ҙ���n�/MH�d��㵕d=��-�֒��4%`��]��)��&(�ͺn��\8lҖ��[`c�c�j�g&VQߔ�U���izݰ�M�-���e6�e�;в����N����]�0��80��9.��r|bf��^�O��4�͘��x�ʺ.�C�v�"q�%�����[���oE���;���V;s�t�:܂�wؒ�Vbf�������={8�kQ�`l��Fw<}��LV��7x�%��{�&�bw]�z�z��qa�C`ٵ��h"GĀh
6�UF/y�¡V֔D��-����\-��֥LaQ��S��[q�C-2�m��[G+�0��+F�[amR���fZ�,�fQW�DPA��Z�fb�ҩ�r��1�cB�UU2�1�R�E��2��J5(�)j2�TL�&
-\l�q��*���cE���cnf�pQQ,��J2��AQqspm�Z"3���q���Z9�.5Ī%����e���9��0V�.��s
��`�kkjQ����W31fL���+��1Tb�cVe�����jW2���fd��QF+�*9W�Ԣ�LqS2��4k-R���na�*�c����1�0�QX6�1Qm
�E�ߺ��~=��㾮�u�^�����[{tdw0Ur�f�x����%���ԭ/�&�!�d�[�W��Qm�I���b���%����{kV(a��:x�|)���,Q3Oz���z@��u���Vؕ�-��UYj�ĸ*��mׅ@+�O^�^����bs}��z����[��l-u���6H����vN�A��V��庄�W�R�cj�X�;pˊ���ss�6*�ޡ�"�X"I�z82��}�^V�^�U����԰k6Y&�F��Z����ř���9�����:}=�vx/`/����{�L9�Z'���<L�Ls��C�V�	W*�ѬR~�^�����\�Sy�6��vӟR�P*F�T���԰9���g���,�SsC2cQsx�3�ҝ���=
ra�1P�G�L�$�0B��FО���%2"n���Mk�.��ck�;
I���
t�aE#�̆#A�,�^�Ⓦ�1�N8v����qq�������|]���t��L�ܶ�2���3,F��i��D�y�������R�B��-k"r��)U8�W,�$ԭ�![U��=�'��N*'�B��/!�95R��Ͽ
>�+w�ԋ|�t��F+��<�)i;9k����g���8�Sc*���(�y��R'^�cӶ���M�����pjQ��޹4b�:M�uㅝ���W��m�><�#C��Ѽg���]�R�0kܫI=�P����7�c~�0��xp<x֘ȡQrcE�^�V������F�L�f*k2%" '���겕��q>7Oʓ���_�σt|0D�-u�o��c�"����t?$�M��q�lHx��TU;|)׍.2x�F	w==�ѕǲ�>�M-ߪ�x!:�a�8f+΃!dAgT��7�,q�A{�"|��vӘ�S9����,N0jb�҆r"�qZg��$#�l�kr����y�M��Pz{_�xF�cb�O���V)'[�daʋ|dB�W>���o+y�.�,��XY�S�FT�������5����ڦ���e��:�Ry{}���1��u��YKB���Ш������
Z�������EmD8�]
�ۭ�㖛auY�al�������@�ڠ�6
d�t��{��5{UMu�*�ؽ:�*�M�8���a��u�zĢ����[�Xq)��RH���v	٣�M�k��bH΀u�77L�!Ɍ�=}��Q�.��>o��Rk���r��-��b�~�]��w��8���A�f��P�bxፉB ��T�,����ug4�=����ش*�yi+��g*�(�闑-*FP�F�"8�)����B�XO�k/�ԡUV�#L.2��qƜX�GЎ��W�ς�%VU����T�}��nvzOGQP�ǖ�`���Xc�����7��F �*���nI�N,�ç�fs�;����3,����P΋��I�r��4������:�K໲S��\ќk�4t�*Y�	W��f�8V�3v�ur�k3z��}:ȿb�]�ň������+���S�|q6t:��@>���z��3�����ï��ǦuP�;)C=�uX������AS8�<:�ڗ����]�l_M(�b�;�ŉNl�eXE�.������d��e�q~�j��b�l�YR-ܷ��b$-N�:��}��D�0G��H�ܽ�sR�%}��#AM�T=����f����7o�-��v��u�4�=n���i_B!��ï
�K��뷭�-6�&�����.-DB�ۭ��.�2��ldѱ򭳁S�w%bYG͹�5�Deޛ���W�.��)7;�.�4�f��bT�bq�<_yn_�S��&H�;�M
�7+&��Z�l;�=s��
.�R�9�e���f�T��[��l��orYs)e��J�u��Q]�-�8��;��g��fl5AW�If|�\�Cc=B��r��~�vf��;T��-�.&h�RF�ެ"�}צn�`�!�mo����ЍrǾa��[�M��p�"����|Y��<�V�����83���BJ�KX�Y���pw��3�q��F���ÂG\$c=����G��(����pυd_9; �,�-R'2(OM.g�5nQ�nTB��,�^�4]����8�"v�m�mA����ۥj�M�s.!��@����C�\:����<�����lv�]r�I�9U$���d��¿tO��!O���"1Q�@^�q�᜺�HrZ���N�τ�]ۮ7WϽmՙ�e��$d �q\b�@uu�S�o�M���г�\��PI���:��խ��_"/}��;T}Y�S[�W�j�fSv9��:���v6�QMK�NwAf;�e$��k�B��ׄ���N��C��f�.۔�3y.T�P���E��$���W��_���-��ڌ��Y�`9f%�,��
���цC��x�έ��؁�L��b,�\�)P؊҈��U��<�J�����ب���j��B0���B�5�g��4j������	�Ar,�����wW�i����}�-%�%���w20�r�M(�p�J4/zIy- m-ȭ{�Ö�	؞$��&3�*
�îz���_���..��}�u��ӑ�����yL;D�aܒ���١^�p4���2��Ս�%8�_�8˹�rY��l�~�Q�]u�^V���^vӸ�k]q�pٿ>�6k#=��ӝ1��r-6�&�����gB8^R+6CL�P�R��cW;�;dC��P5�[��$�GfÛ�6�
�4o��(`�ͦI��#
�<�`��dc[���v����\��[�C���<L:�KD���X�<K�5T>��J�Z<~7�3�sԂs(�b��x���,�D;��X�^��z��GN��w�=��l�2l��P����
,�cg+��y���Nt����(0����v<�L;�C�N��S�uf�z+/���֣bw^pu���M���m�ƺKK�2�gVJ}��{��y��Hy�x�#5�*q9
�WL��4�p���VS�"R��G5�1gz[�)���j�1�s��OE�;
ra�s�(B�H�Lt��.$oV�;�����\m�e,΋�/\��uTH����r댼
)pK8�},���W6���Hb���2������]j�B"",%=q;�)�4������^n^/OE\��6)Q���C�#�4�o��Ư��C&4Ƿז���'l���ܦO����_e%-^"��'��
t �:-���t�S��R�TH?F�vnץ]�/h��4��i*Ǵ���>+ƕ�+�U��w����]r�+�W%f�19H���`�͒P�,�y�:"�X�.$r�YH��w]T�n��.[Վ�,���5Ü0x�Q)͞m�i��!�
�;1�"(ݭm�32综1b]c�N���k�cbK:Aq:��4��������Ҿ'i��^�3�;PљL�<ثi].Wp6�S�E�`�����&?����'k"ev���c��"vbT�]�{k����.��ev�bk�H;���#�	L�ǧ��������m9f�t�ccb�mym/f�=�0�_ �h7�z�#��3�Y��#��w�p�ј�M��F�l�����Lns�/�9�߷.L}��1K	O�
�-%��ǥEx����N�]p7��43e�'4�:s�:c�d\������G<�c��[�&�zv�3s*B�?>��ũ3ًx=v��7�G;iD5��ںEڪ�4�}Zm�fñA�\��%`�C*�VD�^~K��N�ȿ?fU�ڈ��ͻt:z���S؜	R2�J�:$C9��+8@w�ʮ��6s��s<U��%q�@�];���J��:�f}sP�@5ﰋ;:�j�^�E�",��.�Yf���m4ti�:(W���P������ۼ��kZ��ՊP,�)�g}�p�cV�$^���b�� ��Fz�zI�ԉ��.�լt�@cwk�+�4�Xp�^�ց��^(������ �WN~uz�<+�e>�2.�jٺ��(7��.�<�Ȉ���O4k�Y�PE��ѡٺ�ykl����/x����U�3.����7�%w'�������Y��v��Q��h��渪Mh��n�O�ul�u��dc�ǫ�%�R�����~�F�[sG�8dh�H�z�P�i#��:K��(7u�V�����u�C�,��Xn�A�n�uX��aN���/�G��X�O�?n{�@y �q��ÚQc �	�r	���c�;�q�ᘄY�!w��;__+�pꗊ,h�!�(����Z�V��#���LH��^��1z�F�ݗ.�&8�}�참?���4��'��ʭɢ�,��)%�ݗ�WCg�V՞{q|D�Oa����ٜ
0�0�9��\��In+6h�'����3�	��)=���)q��ʨ���t��Fu�
�HfBͫq��ڊ�d=uCt�ч�j�:���uѼ�F�l�����
C:i�V�&��j���5 �k���jl�.k{5��7���-��F����,��62��s~Wg#N�����&���u�R���%��Υ��S�
�Wω����x��h�t��4j|�1�T</
λ�3pT��)b���uuZ�%��uy���[C7n��$9�>���� Z�r{o��!ϵmɭz�E��9C�7�k;f��pZx���3h�=GB���(�;lsӵ�xb�IfË��c���i���+ٜ�.�=�ZZ*��U~T��\�ڔ�������i���G�-���G�F2�r�����j�p�*�v�gb�#'n9;<ṃ�\���;wr�)�9���Q�7���a�;N#�J�_R�G�F����1�K�gO�/�d2M\�`���4�=�9^DP��g*0�sf\3�Q� �<WV�)ndgeB�ܼM�uE	᪸E�F3�'�٥q�n�l��8K�c\��#6-Sy�#�@��ELC�TF�k�MQ�a���Q%��K�n����HD�:�,]ʹ�t��p�f�F�'A)y�A�}�m�P��}㠞�Ot��z3��9f߹j����i�[	@u��<+_N��oG�xEe}-�Y��<޿,y�m�:��P.�U�Bh�B�íjxi��uܩS"z9R��L��o�Ք�:C��%
�I.Gm3$'сF^��0D�����b�'w���r'�<��.{V/��U{�,�ɛVN[�.�تd��<�@5��dN�oٞ����M%��)}�{^<�/4k���J-��s�y�a�Wy��φ9�Q�\&�s���ihRU;��1���ӻ��/w��o6��P�+*�`p�V�N���h�f�y��������rQ�����nk�U�=�cU�GNK/  {�3�)�Jf����uT���-��ZA=t�����O<�B���KZR1$=��t�nL\J�.�tl�|}��+��qR��DG�n�&�Z'C+!���Y\��P�*�*�6�.������j�;
�ؑ"̑���/ք�}.!/+ը�Q���y��V��c�f�*D�qG����X�<`�Q����c� h'6��;��6��j�$wB���N8��Gc�FO�k�\e�(�$���vBw��⹺���ݬ�$�ʨs�B���*i�(�ڬ�5[|��Q[�/���be�j�����P��dGN��,�'�23�$�o�e_t��ߠE�Eq?N���r���[ADWz@�D(e��&�*t`���,:f����^̭�ͻ���=t��s0��\�P�Ǡwr͘����fE30�9"rr���(�z���M!�Fx�&;MuJ@�3f)N�wWd�,�gJ�����;�#6���?�rf�Wso8��=�]�aTyҮrj,�.V�9���O��C�]'C��J�Plڛ�	����������������K�F�&sk�cu��L�[gf�9�'�w�k튺��Ձ��3���U�GP��XI�N]R�ԕ��ڣ���WRrZ)e��z�8��dܮ,�#�u��W����@�o���Wf�%L�4��V������Dx��y�Q��bd9Z�9.X�S/���q���B+i�uq�P.�3���v�<{]�w����2�KKn����\c�g%l��)�s�J�[/��7���h��;S9Qr�XݗHVI([��:�i�p���%��-�+s��;��J���)�(�����]Xn�}P=���բ-�֬��X[G����	jMJE(X�o�6[ܟm$���g���w�Eе����#B\VYI\����9+Y#�D��M+ ���8�;�۷��b �����o�:\U��invU^�[� ��Y}�<9Q@P��]��n����\���ܝHdݑK;����
ת�ۺgc�#dm���b����WKJ٧�Qe��:kr��Ԡu�����.؏��ڔ���u��;��2!-����K����鋳bߴ\03\e\������,�Z!Q���ΎuwΏ��z��i��=���1]����oiWN�ee5#0ağm>&ѝK�:"e�iEǑ�cy�Գ��F�)���[v�{iK�}km��<��ic0v��m]G��#N�<�`���QQ��ə*}Y�(@f՜(C���-7��.�X�]�P;�p���S.�V���5:�U>�[�O���ڼ��>��:��t@
]f�"2�n�n�:r�����Vd��kkGQۻ��� �Z��3O�&Vb}����<�s��Jp彂[��3O*��4��o����!��:���٭˰�
)�{��!V��tr^Wh���֭W��h�$����ɭ.��X���屇�7��/��;���t����dJ����)��g0�@$��p�ӊ���R]/k<��i#��<u��v���@扛��#]���s��m�
�9�9�d`��pli��N-,���ۯ�z^�d,uu'�����n���$�IN���I����f���L.�������$��^H�����ƾ�R�֊eŗ.e�9��0qLj�
Z�\ks�U��.d�\pE���X��Q�Qjʕ)��pZU���Q���l�
�kd�q�
c���-X��嶩�(ԣ��5*G��D\�C�٘\j��FƌV��Ym��E����Q��e(�����Q�f4E��r��f��,�m��]\ʓ�T����e�pr�օ��]a��*�:h��e���f2���QEC]k,�Y���Jʒ�U+F:�m��M�1H�T�SV��崥Z���LmՆ,WLӧF�nCL�`�e���\Te���U��4�
&�t�MZ6�-c�YtՅ�Yt�SH%�m(���j�WY��E5u�kY�Z�TR�*ZT�G1��sWL�X1���M%�5�KKk��`QE]aQM[Lr匶�3*�ڵ�c�f4���.���"�������h(��,��Ι/�},b:�,�����ZN��u�rJ���Ok��oLX�r]�lͫ�.�-��=��tX�=I��u-�]��%�wݢ�P�BV�U�G	є���~T�����/�C�i=93����RN�c�LO�i�3`�͒T�f(!'��G\�q<�Gw&-�"Y�x�mM���TC��ɈY��A��,Jsg3�b�D��<������� ���Ͳ�|q`�����3{P�518h(g"(>
�u�dvs�����x�d$Wg+s6r�(a�i�;s,�����=��U�'}EjqMf�>��u�sn����>�g�]�9�,�b�7�t͍�X���;�e�d`ƅw7ΩD%��KS{8�c��M�(�ł���Y�q�Q눿Su��T�9��=Ֆr����{���"�wR=���i���'6V�5�#fC91$ F:Os���loe^.y����u��"�:t��:F�&���f]	�TYbvie���Kf����Ɯ���!�P�H/��n�"�t�����=H�闑6V�ۺ.ڼTQ���T�om`�4�����������lv���]:F-�ʅ�
�'4͍�'8�kx�+9<��y��^��l|aՃ{ۍxh����h�X%�Ng.����u��=�}Ϲ�'-َ�9�A�5oh���bn��x����C.���˝4�2�H���Щ{C�<D��T�BbY����3ˁ��Ϧ��4Bd�t�,��Y�UH��*bK�G$^�'][Oa�'���۸n�rk>�5��	Z�
��Z�i]�ţĎ>Fs𕥊��L@9�ԷX#�h���Χ��꣌L���7�dU�j��a�DH� p���;z�.YUȌ�5�M��j�frE9�LR�.Ī�qG�u�EҤb�!H�8`Aq�����f����ޡi��˅�\2��܋����0�pNp�R�aA�D\o�X�De�������AV �HX����4ÚQ~�3��1!s`�b��2�=�B��k�12��`��4�2C�@�s�0f��:���ޢi��dG�1Cs�ҳؔ�[�U;7��\�z&!BE�u��eRT�t'yN3-1鳅�3R�����=��sm����;��������L�Ue��^R�M�xl��r|����5�7��[-�f߆p�q��-�(�U��XVZ��ɫ�>$g���ΧTX<uj�;�
;h]ni��dھ�%sf�������;�7���P�F���M[�{M�E�;�a�{Vn�>�O�Z���p��O�p��K��{C�kj��T�Y��V� �ځ{p��DU�I)����BH�5�,��+�-@g��^�~}��l|�J��P ������-��	���|��z�hp��({����:�6����cζ��&��Ѫ�w��]��6.���SN��plۢG�o��#�::m�0j���[�S��ߗt-_x�Z�\T��҆��,��F�ʈW�eQ%��%b��<�p�_#��f�~ٛ�g@@3�q	;P��;<ṃ{6]d��u��w���� �s���xw�VD�^���Q	���08n�z|�\���~(����2�{��x�!�1H{|�"+�r��Vf�b\�Q��r�귝7P�)W��ZG��3�'{�(*���sFC�L­���l�mM�r���b	�ƈ��vDkAƯj*���$��W^�r��n ú[k��$�R�R�%��a������]\b"�I�9,� &J��]^�L��˶+���r%�����ހ���>ȧS]kF:U�o��ө�v�"�,Li���R�s�9
��,��c)�ȕ}ϝ%
�q��� )�)j�FQ<6����h"�Թ��Ѕ�(\�s����랢�ַ�����v��pb�J\E!2�"��%V򢝹Ƙ�\^q�cOu��Y��[�AD�H�ќ�ԃ�d,�;>�G��پ�}����E����MFs���� {mx!�{�	�j�O�M�P��kʱBc�d�0o�������&~�Ÿb�YS��wV����6l>�6`�R;9f�_�Ƹd�A��3�FǝM|0K~�N�WPuw!3�aJ���u���9�F;�j�pLV���8���ÞZ��x� vs�>�܍�s1���ϫyŷ�=G����\�����"�ϸ�(��oC*�K."pH25�*�U��-�R�c{/���G�3�|S�1A�T6�H�>"3Ⅱ:]vC�ڨF��I'O/:3�4�r�{�f�r�yN�T9Ɍq� Q胢�rH�1����kSW@�9p��7��� (�=��n��td�J�FvL��FTU�:R�ҕ�C�[�%�C��'(�D��E�_ro���ã��"��Vum�&��-�f;9��J�`�i<{JF���XӤ�ݬ�|��3�� ���qC���$N�k5�C�2�yI(�Y�kE���{k�WC$
t�^���u�y+n�~.�Wl΀R�ʙ.��l+HF�7ٙނak�ew����{�e����L::�Q�h��[l>/��.�^O#��e��M��t�+Ќ�
"@�,�8ր`#"�YT qʈ���$�ū9Us�L3^�}���1��A��PU�Uk��Vc�z�Ê�9��`�6����fb����A�J�j�c�1��¥��3�����ee1z����Y�T��;^��lݪ��$�.,����(pBu��Fp�9�Y0YӪ��ݼ���0{�X�:�s�O[u�+
L�\H�LD�	�DW�3�v�/1:t��6��5ڄ��p`��iˌ/}3g(<���tݳ��P���:|�v:�]�ݥA{{��-��˖�g���}qkA�q�:!�"�)L�f�N�T�@f�,^�I-:!b�]otV`�\����7z�q�uf���G�'b�c�p��w+ �g,�B���ta��om�}��@7-VnN�R��m󨷶������ޥ�T���zV-����x�7L�&j�n���g��5>x�G�_,�;����=��jb�P�gǥE.bE7Zo*x�Ӹ�Tk���i�WV��/a�v��}L�飇��1Ay���N�5�ׄEn�Ý@efwvv�bk��˰E=�`��q�,�wH�
�H�~o�M�_+sB�N��if�ǉb�H�#+gb/6Q��"l���t&�bn"�RG2�s�E�(�ar#	���zg��s$q��F릅�q~�'�t"p�x�r!LZ�ꓻ��L(��4l#���:Qv&Q�tg�4si�3���Fןq�#͍z��Unoι%���Gb	^�FP�8�x�yxN>K�Td^��S��:X��]�p/���T�ȋ��^���H��Y�	�uxOlpf3i��\�Um��s��!�N��aq�N5C���8�#iR1P ����w5CT�����7�{qqr�8�(�c%>�n�E~����6|�	��Wr��l:�2�]�{�vѺX��ZE�PF�-�Yc�or����q��i���ҷ]S\ꜘ= �6&�`h�o.���p?�#Pni�W,��ʝ:��6�̫U��@�턙�)f�w	c�,Y�����h��\ҋ�1P+�1��g�`#�����X��3։��}�(�/����nF�5�"��[����0k�	�]��o�t-ȡ���XbҘؘ��AVa�Ӄ�%NL�bx�.�Ʒ��k�3�˽j��k �����U��b��2e���Ve�wa���{)P�Iet:��>s�Y>ɣ���/�����)�8t5�fZ��	e,ڷ(M꬜ஞ�k����5��+���)�^���
��JC:^���k�8Q��t5R�M��y����LC^��0�����i֊�@���q��:+����δ�,�c�ڨ�w�Nw��r�zAg��P��*#�;lO�$�ɔ�if�x�d�Su��u������U����@�)BEKl�(m���<�9���c����{���cΝ~ޡ �*{��:!��(��F� oӳƭ�#A�)踙���G@U�>Dn�E����؎��bX�|&w�v	[�IA���N�����d�'�M��1r�G5�����=�)׾u�p{���I��Zy��ٯ
ns:W�ُ�M_v>�h*���`W�Nh�{Ժt}�D椅qpl��ؼ �:���{�~�6�uiZ�R#����_z�x^���96�4U]fF�qr��3�dc���\F�J�ʊnXC���4X���̧��/�r}�Q$3���!͞��˔tT-�Q�ji��J2�Ʌ^���w��=#���$|��y�VQ�N�#e�Ab���x�����C����=,�s�uʮ������)S0X�g B4���"A�<dp����R�������osw�a�u�j�
���p�e�Y�F�"$VU�p�)W3��z�u���#�ȳ1�K���T�Y$SFrLPH*�îҰ�ϑ�cd2�+���~���\�	Ƞ�����%��%�m3$'��C�N��./���AS��)C���ʠȬ�@׍�p�ŕ#��'ݞz< ��v��t(������f^�e���vv��0�[�t��b�{5WPvk�5?].�~q"���U�y�L�|���ɼZ)=���"Ɗ�ƶG�:�`����A\�@y���
��㴓�#6�]ĳ#ͦ�*YS�k��4��7n`@Lm�R�#���-�q�A� 9.oz��T/�v���R���o�Rm��jL��8
�����ܕӒ)��
��g$zT�٠��|5�W1V�������c��\�"��J�l��������s��R,����ڞPm8�Am@ۘ�wa����;��}�-�ˑ�7���)x95��������������;[�ݬ���;�#���ڹ�C�s���:0�{�GA7��Ln���N,��0�{���J�_��[���V������B�]�]v��gF Y�*\G9�ʡ�uϣ�{*:�s��]-�cf�_wVM�IFW�`G>%l5"�N����/
�1��� �Bǔ{R�6��O C�,��.���+&{U^7��V\��݇�u��i�L��7�Ըy+�ʫ�;+>f�HP�)2��:f��m���b�`�G�N\M�ʯ�
�a"�$�.e�m�X�TP�}h懻���� 1�z:��k.�����>b�*�#u�N�[�rf�Cucݕ���xf�����	�Ӣk=IX���yBd��b);�Ѹ2g�̙gsr�y�㎪b
ȧ�5#�*���oJ����O'�l�l1#�5��T��=�9Em[�E\����N]!-��)7��U�"O{��\3��nm�W�����7�6�U˟^4$�M�S�:��X��XX�s����ya-���CC��ss S{7si��A�\�)���m���Lļw�}��fp~���b6��'bĢN�{W��@g��w3��*�]8���m�Ñ�FZ\�V�+�Rf08N�\�v��Ⱦv�TyOC��5f�C6-f8Ԣ�VC�B�X�՞4�ˌ[���uhO��ȉH.�2��a'��m�V�K�R��������W��?\?s�O�R�UUj��BcNDG�֒q@Dri#��>E��E������7����u٭���H�	�T׆da��ה? ��!od��u�Y,� ���� b3�I�m�/]u����wr��Jv
�}��a�$މ��ֹ �����c�E�K&j*�\a�
#�&����í�x��E@D}�b��i#�Y����S�o�o�����OJ�?���0��t*���@�~ (���{%������3�.3�[2�k"�X��U#���Y~��J]���n��M�D^5Ӝ��0ZS�@�[@Dcƨ
c9m��;E@P!	��N���zU���S��2\��Ҧ��k�<�dw �"9�@��[�h�q��o���H>�n�~���&����G\��٪-�3�sT!�
#���\��o�hN�z����-H��ޕMk $����q�[���"*�-@��Nˇ�\�C�o.^���s@Dv<Hb��8C��gT�ڷ�~)#U�������" �ي<�P{��1O|'9�.�.FSks� L������PA�X�8��p͙d�.:�QFZ��	'���D��|f���K���Sp�-i��%$��)y���PEŘv�9����7��"1Oi�6��n�7�z,�㑫C0>f�p~�D�'>[�:I���	��ּ2����)�!�mI��f`��� �"=GGJ�4�b<R$�>��.��@Dd��v1vg��=t��O?-I�3tf���Ԗ�`Caf�<zP�A5�u˞��>�
ۘ���]�>��y�8�
��u����T1�oޑ=r�d�v"���S���a���r�AdIQpg��P���uF(�P��h���u�Ԁ�S;5�d�!
�>�y�u,��"�|�ۖh壃��ܑN$<θ��