BZh91AY&SY��d��+ߔpy����߰����  a5�} ���à �"�@    h @.�ڲ�P9ܪ�H)QB�U%����QBTQ	J*�T
T�|�P�Cm��h$��`� �� (� P@P    �  ����g��{<�����}��{i�g!����9�w�}�}���z:���Q���r�{��o�F���h>�u{�>�K��{��*���Ϡ�;�v���󰻹@8  � ���^  �}���7��w�w����R�m���[���=�r�w��>�ϯ��_vP>���X7���k�;����Ox�"���AٖތϨ���l6������ � |�n=�  
�;o}�#��:�	�^�>�͎�'@������:> �= Pý]�r��}�m�Kݚ97��f��Н�}�}ۢ������>� 8���p  |QN�>��rݾ��|��>���{�9�T�>��LϷwP(w�a�=�s�/N�<��oO#�$=��;�y�n���{����������m.=p @�=ؾ���=��{����:��8�o��ýﾍ���n�ӹ �g>���C���}7�����C����}�yR���s���(                 �@� 
  ��MꔩTh~�����2h`A�@h������F��	�� !�0 �i�R�
Q� b   # ���J�F� `  24H��A0C@4��?SjhКl�OS�z�)���&�*�S5�f���0 ����1}-���cCi�_ha�#�J�1�HI ��_r-G�? Đ
 ��H��A��=tH����5?������/������Ϗ��B���g�І��l� @J}	��� ��Щ@�$tM$|1)I��L�$,ik�����o��~��������k��Rl���+�|�R'zn�W���%���ze}_7)Oe"s]4c��c����elѧ艷R�1�\����_�JD�r�8�R��c|����H��lKy)�Rp�2�o�7�jR&��H��WM�0�&�=�9���>�ےl�I�pܡ8�WD��UȵT�+2s"u�5S�$�cw*�I���N��U'�������Õ656jDjY��S���KfJ��}��!��A*�e%Y������>���-�{>]I��٫��d�7�]��'(���Gq΢�~��65�UtLwUã�ʡ�n�DsUI�2Iӌ��M�M���7"9:&��L��UXN�A�J�0r�a�����?'2A�H�����c���{z	��b-�G
gf������}o�����pb�=��Lz�������E��RR$�^�/bTOjY�纕�I�%��%�%��I�
���Kw�K\)t����=�t��t�7�AB�z=Mձ5b�"�ilNZL)��)�M�	��ƧM�96=�p�'��S^�SL���l�g�Fd������3���i�	�;�a���6WJ��o��Nٮ&����xr�W�oEQ��6�L���p�kD�H�>�Ө#7;'�&�K#�M	&�Q��d�!V6�p������Z��s-�FiY���r	ϛ�:��$���8Y1�4t��r�BțD�5(Lhy
nj����}6Ch��١�:"�V+"Q�`�D��H����ı��d��y%���ӦTه^JLd����١�D�$DrId�G�:�u+���D��R�G"Q��5rW����jR#ȉ��䯟��X�nR'���+�����D�YUGJ:��[ �6Q��	�ԤG�(y��>jR&����舺���\����H��lKy(�k):^�+���H�{)����vW��+f�?DM�����,����g�JN�nR'�"�VrW��e"k���-�KYI�����R&��D�2�h���4=�D�2�O���)�&�5�^JN��*����2Vd�D�t4ta6:=iH^A����b^�w=+�K�+e�cR�H�K5ȎN��;�V��������RQ�������>�Dy6Yoe"�1��W�Xt�K�i2]���<�G"?t��Ï*�an��G}�M}:#���8?t� ��l�So���r#�0�Z��+���D�ϧ~��J�̸��u�~��$9�9 ��(�f���9�Y���NÐ�����%�7aE�ä{�$RR	�ඤ�R~�?t�c�8�Yz�eIX��Iz$��Q=�Ou'����IbIy$�Ry�Of��qj��Ud�%�㹛������y��g=G�Z燺m����w-�C��s'V�üj�rsUT�-"�Z�x���ޏ��6��F��
«�ޘ��[<�/p�y.yq�0�(ި��h)T���Ě>�����$�Rb4N�,��D۲sBu�sF�'0�ɂG
��YtU�h��"r�u3^Ύ�zMY���	�c�<(��s�h�D�	��u0Τ~XL���:�I9F"p��;��&�J��nC�u�ʒl�9�I�܂_��Ν{&&��I/��I��y �d�Hu�u.�%�Ni��7�Nuk��vx:.o���i��i�H�5�l�*��Z!hZs�����l�V���4ɡ5���ʑ�$�I�jN�I�tH��"bC>D~ϒ��&%��d�>N"u�&|��rG�I��L"�N��L��'N�蘚/$w��᲎�8�P��dL)I�:QC�a�lѦ��na2�'xk��7�0ፓ��P�����DHu�(�Ή�R'o�Bl~�bD�Y>FB"QZ�8��LN�ĭ$D���V(�H��H��
�&�(LM=��6O��앤���fi7�0�L'�N"]$D�"LI�ㄭt�8i�>Fa6h�a+�)I�E}�D�")�|k�"'t�:=�(~N���LN?"D��Ɖ�dI�Cp�a�DN��6P�`�bQ�L�M����d�9:��I���D�o��������E��D�$Ha�L�Პ��K��%%��� hH��H��=O$�;��s�a���HA��P���NdN	��k��.p{�#�����N��gdF�wr��h�r�wʉ��藂1���K�r��Aȝ4�J5���b5�D�Ld4k�����Gr��YxhzA�e!Xt�bgg�t�U,�j�5��Y�6�J:�Hw����[��^Ҹ����e	d�>��H��u0s�r�^%$�$4f��MDwn��$Is7�eO�z&�ʛ4����'�'C���ڛ6���+s��m��\{>G�9&ƷS_']��ژkr; ɲSS��O�c����I���Q�n�᨝ ��8kSxH��6i�@A��r�'d6%`�4"�6i�AU43uA7;S�uUn�k|�e�u:A��uQ6p��#֦	LNuR�u4�����eTD{ʈ�d��u��c����A���r�	�ʉ�5�B0��H��I0�Z��5S�":�D�֥	�56A�"p��f�":�DK�R�2|vDHV�"�����9mM�P�|�ʨ�;{����;�=����6<�DMډ���Bs�M�r|�4�١ʈ��j"^��A�����Dؽ�B3*"rڛ!��=�P���Dѣf��b5̩�Z��D����9֣�+���|�K����n
��E��ۂ��C>�߄�I>G��P�K�fX��9D;�Qϑ���ǱΕ�9�T�f��Գ���	���ڛ(G�q��jlM�dB�gBBT.����~�G&hތC_9$'�� �|���6Ϭ)�A�thuu��Nv���,��t�87��1�TbRa�jp�����M�S�mʛ/�7%G�5!�ƹ��s�ܐmS�HjQ�O��6g�f��3���&̐Ƚ[=c=c=��#f�ԯ�9S[$���wQ��yڏr�ܨ�N��;&�e�����c��yʏyQyS��T���ʕd�	��闕��u������m�Ϳ2�C���y����O7�n��E�05௃<t��J%UbcG3�q;GL仝.b;F�Y��y�>�c�=�w�8��vGsCɝ���ܼ����^j�ȗd�M������{g���a�*�&�p�t�+<���c�����v+���;:=�`Ȕ�d��㩣7!���b$=>�D�i��q�������a:��/t�t�F8�x������%ʎDGs�reDާ��r�ή�|�8�6n�hA�3�ToU(n�=�9��Tjv�$NT�jt�I:�,�|`�"&�W~��֥|�D�O�0j' �{+��Ț�"<��ܔ!ږ%;��������E\D�e"l�:Q��Z�����䭚5�DM������C����R�5�q�{��~y�dPG�}p~V�)'����N#�/�|�����(�co�j!�6'����2����>�h�|`��^�}4��-�P�p��V�J'���y�q����Z�c7�v*���gwɇ~��E�������tw#|vz�5��ꆡy!�4��G�ϩ�ȫ�I$����X*+|0�I9�9'�	Xv��8^�=٦��\9=4b��Q��ۑzx��0�[�N����D�F�J7Y}�Y޾
I*��[q�^V�����py#�O�~�^(��g"����8"�f�B1����t~�X�c-Ԡ5_u�����-��r�4���=���^��w����ٱtT�o@y6]j2�e1OG@i�5%)���&Xa���9�ܝ�u�/
9
ny�ٹ�����O�a�	c__oi-녞�+Dfd%����&�l�l2�ca�ɻ�2x!D�nM�Xw8�m�{���$���m�҉$�Z¼*��h���=�������ں"�5P1�gHI�WrnR�L�J��s�
,%���I4��2i��v�T b%���DN9MI����;s��ޙN�F�|x>�7)�L~`mE�g����Q�C�!��ƌKC ��Ftd�rI,:���3Z�  t�7�����֘�嫢��@<c�EW��{��'�^]��(�}'��z]�[k� �.17螎��7g5�h`v_I�E�hld;&�ja��~��Ѯ �^Q�ݎ���t`$�s���{Wvs��;����~<�By�҉$���PǶ��4`��  ����{v�ċ7G�4aÄ43�B�9�_w��>D�lr� h~ =�P 9�����'��z���G������:1.W����t�l��Z���ּ��!��
z�i�A��ԇM׵�SaGᘀ{��+�5� � �9������n'�o��  k�n��C�l��zp ����(��=}4 x|ԓ�=�O�1N�wo����_��6�fиH��}ONLSe<�()���Z7�4�N�f>��:s�O[�xk�4IFx7�����Qp\�w<��4��
�%�<_��i<�䧁@��SY|ٽ�7�z�p��O������:���BLp�#J�b��Jv�3M7�	�Ŏ�)環Eu��wP����N�0bOF�f%F�.>r�R%�!����;o΂���%�Nss�^ ���Y@u��HjK\<�t��Y��!{�k9���Q�V�;&���A���Z_���*Z���1 rsk�3@�#(�i]�mq\٘[�Q�,�Dg�dݽ����|��t��3_��w	�-u��H���Ի�1��C�k�}���������-���޸Q�� �����}�ڨ�X�m ��Nj�).����޳�I�3نy����_O�0��N0:^o�ܩ�"�L�`]{{9�'gH�z��!�K�P���wvs֤�<CC<�����!�9\�P�M�m˷
���ಛ63�ޮ�vi)�o������z!|��׍��ӆ��N�;Ǩ%ݾlݫ� �/!�>8sڐJ������♭��K���f�@:e���tI��k���C�֧�Ů��'�L$�E9�,t��I$�J-���	�=3#z�~xɎ�O^�F�N����INI����n�����P�8ۍ��K�s#%�VG�wk�l;�9���Q%��qz���^M�w�����$Ie{[��׉�8Q�X�/: bٔ5�u'�|����Ã5������.�Y!�����݅$ԣ4Yo���ݜ]���  R�g���p�ٶ��v�4�D��%�kZ.��6 l|ܐr�� ���ڀ xz4�����͚&� ��3�-�1��wsg���4oz]}�L���dղ�����������c���U��,���S�w;��:@��v/fڋ$�u���q��l�z)ٯk^� �{Aewr���]擽B�`�|p�!�Q9ܶ�|@�����׹��J@z�1����h[� t`b@91o��h�Pr@��I86��t��f�m�t�3e��U[d���;�i�눛���M9zRv�Nt����z�w!�d��<�Ӕ��Rr�.��G�??~����R��0&� {�R����������gǰ�`
O���/H|z�r�el�������N�d�a���H )	l���D�>ǖ���-F��W{o|�+zp�1����V����ٌ�9d���HMw��y�i/�� �   <x�)�� t`J�l��`��Q(�(��i�k�?��"p i�Z��5�q]���������  ��y!�vS�m�O ���g6���T;�j���e :N��Gッę~  x` |0�$>  F �83<g�    �I�5gL��w>(å}�ϲ��$�9�8�>Ԁ hpz��l��'$ )�]l�έ��;����䩺}	��̍����� 5�H|R1'�Ojh� pѷ|S���� m�f�p`  7�q;��(�1Cƺ0 �',�u�gu  jH|,�P��=�i��`��w��{���:%�C�=�LP���i0�po�eߥ4����z�E=>���ႤI4�P��o� w�.����rB�h�7�t�խ�|v�9
��:��ŤY7 6�f�Z�W�[��~%��vQ�|��F `(��U�w�EcoѹMrCc cؗz��^/��ܐ}��Η�
},љ�{��M��A���c�ԓ��۬�x�h���l�ksO�A��9&��F4�P���QN����ON>�||^y�b�&N�[^�	6q��60c HA줦��� I
7��C 40R;׏�v���a�^67� c ^��S5���������~���l H6n� 0y9�+�2�(�smÅ�|yُDV�/��7�������2O�9Q9���V�ӓ\��t�a�+;��k�}:���{}�*ޞ �f�~+B߼�^�uf��5�~�BD<����d��Ҥh��w�f=u������ �](���e�J�w�o�I��m��)��Hh�L����b��;���.��O=�l�_�ɹ�ۏۏR�%w~�l��GF�>Hi�A��o��rѓ[��e( po��?f������F�w8��'�~'�:B�W&�浥Y�M͓C�-᨝���Xz��p��|� �޷u�Q���e�l�I����d
=�wu�Ql`��v�:0
1e#�f�llaye9�k��͎ ׏E�S���)�v0 ���̈́�MY�{�{\���=����_.�&릯�t����Q�[u�oRp�e:i�>����x��[BnL$����O+:Q��j =]}f�8tPSЯa,����hО1���Lp�o\A��'��c��׬��!��q�B^��x�? ��"��vۣQc��������H?����3���={���=〙���Z�W�~��n~ lM/�O��~C�>�[1E�&&!�c�q;�J���a��)��:��z}�zޭr�L�bI)ܝZ�(���X��y@д/'���d��.���؁����V������T���1u�&!4
�y��z��m���X�Q%r�?�1���k��v%D��hKhJ��J&�j�Y\j�Z aיjo	-���BKZx�^������D�8U1X�i�I�S. �j�=i�:�b�"U3MVf+�wE����,�dBb0P�h��'���r��%�r܆��ԓ�H�P�>k.���2�4�Q$��qU�-�cH�B��YɨE������X`U�8Q(��G/�hbLm}R��-�ްI�*j��\������J���� �����*{���OL���$	��G�,ؑZ��4f1D$`sV�l��ZZZZ<:�=�$;(hUTֵ\H�T �iֶ�k����K��B&`J0�@�<��c�1�m���gT֭�¼��ƨ�����D0�F-� ���;�1^�G�	�ς���p��ȁ< �NAD嗖Y켖�
��B]�x����nC��r׭&%��VhF�6$"��:if4%:Q�Ij�����)<�V���Cq=�y��:�W�Z�ǔ-��k�!��
����ʢc��"U&N&�0Ƭp�*E��Z6��}��?w�T��m�����4��fd��V�.M���J�;��]e�N����{�dm$����7�j��xr�hn�2$S�r�A��nRSq�U�����9�u煰ph�=��F�B��ѩ� X툶J����i��6%����[j���H!�kl�驑�3�����F�N :֙z�R�����������R�o�������C���f�Z%��[1������*i��aǦ6�M.1[+Q�8\�q	gZ81��F�$eB8���6�0��11SB�IC4�02�� �������BKy u�m+j����3���k�g4�x�֩8҂��Y�x�̢T�W�,�Zjw\��b>�}���I$�ܝ�l�6	�?��`A��}�a�������J�>���%}�>��������>���/�J��1UU�*��+��U�]*�[Uv�ګ�V�]����WJ�Ŋ���*�ݢ���U\b��V�Uz���U�V�]�J��Uz���U�]"��UUq���]*���WJ��UUq���[X��l�����R�b�m��
YVI-,bL`�6 Lm4�Ƅ�I�2�E���k�n�7P)Kd�Л$�i6��m � �D/�O���*�|ꊪ�������1UW�J��q�U^+�Ux��U�UU�Ҫ�V�t��UҪ�ZUW��������UUQUU�*��t��U��U\EU^�*���ZUW�����U^+�Uڭ�J��U�V��Gn���F��m	&0M�����Ci�ʱ"Ԋ����%X�b��j#�5Ka,�IlBضԶ�U�j���l�I���U�[j�,Y�� ���;�UҪ�WJ�Ŋ��������1UUQUUQ�Uz������V�Wj���ҫj��t��V�U괪�V*��EU^�J��[V�U��U\EUx��[Uv�*��UUTUU��Um\v�UUb�T��>��m��RZGU������4��T��Y�%�i-ȶ	��lb�؇��;���]�9�_8���U�V�]�J��b��,UUŊ���UW*���U\n*�W���Wj���U�Uڭ���mWJ��iU^���V�Uy�mWJ�Ŋ��U�UmUڮ�W�UqU�UҪ�H�U/]�&Ţ!�1�C�	m�-H��l�QՉ�'(�b�-�uB�B[l�P�Đ�6��$��(hI�!���K!��JM�4�4�����M	C@��D0P�BM����J$�.5{�|��}i � �&?��o��?�������>���}g�(�f�0�gDL0N�F�P � �"@�A(D�,M�8'��pH""'Dě �"P��:"`�����8YBB�ABh��M	�b'���&0L�""aӂh��B&�,舉�t�$4A4&�N�0D�"lM	�bl�4t���b"`�G
DJb � �tM�bX�!bX�CBQ�O�A� �! ��4&ć:t�f͈��=��}�%���]p��B(W�FE�Z�@������g�u�36lC[���c�:���K�պ�+�f��e��[h�A)�m0۔!6��̝u��Ԛ~o�͛�ai�k�p�K���;�[S}f������j�d��p�ho�|Km��j�m5�4�A��s�\�z��33f�,20���)Z롆�l�-� Pidq�((��ݦ����M��K٭��XCk�)bZ� Z]I�[5�����-� �b��eP�r�A����ٴ��P��e%�f�������K�t��r?��������	�����jK�J�ŪK�YM�є�h�m�cm�bX���ϵ&�f5+��@ItvW4��c ˿ǟQ�>��湶��>��Hԥm��atFe�����X�B��:�i�
FK�l[m�������t��j6�U�b�P���1J�h�o�����V�1[���*l��]���]�+Y��Hl��k���a0�w�'~OK���lmFḋ6���ؒ�ګ[���[s[yKbaX;k���NMM��aT`��uk]�J�y+=~�X|�m�7S!]-��F�T66�lؘZ�Qх�5ٻ .����J��ηfjQ�j�:]@�-����<�z b>n��4V��.QV��v�b������ua��֗���[u�q�/��iaW
Wg{6VЬ�\�)������nl�݊��ˉ�,e�Gm\J6]��A�.��޻X�fe��AӺ���Q�r�EQ�Nuqm5�U��.,���b���3U ��8]���a���Jf��DZ�U�M�j�_����~�= �oc<땦5�5�f����D��x���g�Y�S�r93��Yq� �"nN�e����4:QZ�S4�5��v8:��j�y��v.�wj��m����h�9-it.���x=�g���[�����=kfˮ�&�"�]DN���l6�nh9n)�u <�-̇]t]CXk.e��e&�)w&�5(��kn�mκr�I�ɑ��]��Y��#�앣*b��-�Zh�D���6՗��C�Z뵬� �h뙖�\��u��))b-
���[b�������Cp��Ll�0�)%V siA%����4r)$��0P�r���Kԅ�Vŵ�X��6"�WV�חZn�b��tЌ��$��%��5jْ�͵��;�_v�L��v���2�(k6*�/M �v����t��q��l��󐱳G:X6��]fZ�4���I4����Q�K�IXh�Փ�XF>=��#�uSfO[�z]�MF8Z�,MQV�*�#�Խ��Z�D��Rع��z�,ڰRF�̭�9��i��2T Y-b��]�z��ɳ��!DM6�q��=��<l��FR�5���gV��pE�JFX���SGCs�0`����v�Y,^�����Re	kw��!1]aP��k��Fgahb�P4s�lT܉U�W^ĵ���c�x_������Z���
��Kr� .���a%X�ЛR㫬?G���i���795���Z.a�Yst�a�v���t�� �,V�h���m���It�tƊ�H�~�J���c<5�n �k�nɡ56��l��6�t�+]5�4m�ad�IWf��V����������2�fRb��.�eff&e��w+�\�/Wn�v��5-��Ma]�94Hf����ڇ����Pu�:�Ш)Ym���{|�	o��c�T���%ݭ+.�뵎��qԍ���%�I�w���a2�e7KP�.A��M�և�6s�
5紥��m�M���@\%������o�;�ٙ��U\b�~��7��ȮffyEUW�߾������{�+���QUU�*�����,\���"���Uo��}�0�YD,�BhK�pDL�������}H��e�F�c�_���{i�!�e��,TT�"ƹ�L7)��Wk�6�cv�"ؤVˡ5���BB�J�!mq�[���)>}���x�f��^��c��	�����{�@��*Z|A�m /Z2�]4�6��9�D��-�%m&av�����]^�!����Mm�Ш�&њ*K��&�,B�U�:4mhh��l͚\�Y�]��)���2�v%����y2�8�ݯh��L@Q�̚�2��a�0��*Z�d�R�]u�^����+	��5d��F	7nf������0'��s�שt�dv�X��������qlu��s�In��U,�5K�%��P �N����J�E�T#�z�-�N �ⰝZw�[#̖� ����	��1#l���C�R6�V����_8P��6���l���m�3�F,��%	���iA�$�Ԡ{ni��Gw;n��@�tk��[m�5եDR���Gq�F!ڃ����\�3�/FT���
� ���Ƣ|ƕ% 9��UE��hUY���,���D�,�(�:�z����Ž� ��9�������$��(�of��ơ�E.�[cm���Jl��!�(��K)������kD4�7��ƱYGkZ�#܉v�L���>�y�Hb�빞��4�Y�'Uͭ�ym�s}�]Op8N�A�4b9��"�
��&Ë���6�m�ƕ�z۷�������a��>����+P�$���"p;���z��J��),�4Z���H�4�}XA��M��1˅!�K��EH�b��kp�������[v�r�^�/=�Gx;��m$��0)�!�M����f��8/Ed�����e"�#JGElw�҈�(�/��.���^�`��\y��tc���cֺ��m۶�p�J㍻m㎘x���%�%K*g�MO� ��h;@ËX��[�.��s҈��B7�(��y���h}��*�MX��1d���[����>.| ��� Q�����99#h��/6�qGij�}�Zi��06�cR&q],)F��z1��M%E�:��g>6p�i!ӌ���a܆�0�pѰ��Yf��8X�<pDL����Y�'3�<Ín� KSoKᨬy`�0҅N �l�����MB6��@ ��9*�!6�o$��$��\�Z�R+΄٥�>�\�Qp��i��.ҍ��e���v�Ck�1�㽶���lGGlSU��V�V�o��kf3����q�v��¸7��m��u�0�4�]Fh}�CqF��.�8a�Q��Za��4�bH�d�̼�c��޴�Q�����)���!#'�f����3��YK|f�m���P��I��&�*�\�j�����Lj�m��qc��\^*=v��iU��yt�l���vq�q��6�ǯ^��8׵���Ըz��sڭ��Ke�Z>�����!�Y�1q�]7��sd:�m����D��e��֎�����8/0�HL`�Il�*PW�� ��Qi}���bh��-h��!f]�E�10�b��';����`�`,#'�:-��B���]�'R��7mJk���:�:�4U�;�hЍ�)����RwL����n�6��J㍱��Ǯވ�&	��en��%h�kEUU���1B1N��R��D��$�H�4���3�5�2�H������Ƚ��*�pB���E�{�sw32����7�f���1N�
�	< ��8A�[S�ÈZ:�iR �o��B��"�Pt��kGwZ4o�\�P��5��p��h��E4�N1�7�4��f�T�IAD��,���"pDL�tL�ϵ5Ԓ6�E���6��I���E!h�7��\q��m�l��M��Y&�#��S4+ƫ�9�|�9Ӽ�nZӓf��5��m��洶�W1ۥ5NS7��m�\��:�5o��j	��B)b4m��S����gˈUq�>Q<��1��.�����`�kgb�B���	$�N�2�4x�����"`�'�a����E2_�>7,*h,%���݄��C��$Va���w�p̊l�5Em��@�&T+S0v��{֕�� �5MҎ�7�uV���Mf��\R�.�u\钛Yj8ז�`�ܻ��&����ve�n��*���וw~ǐ���k�3�Ǎ����Ohf�jՑa(�Q�wȈ�m7�H{-Z#cޡZ�����T�DG�'1`���ʹ��Bh��ɰd��qb�4ݑ�h)���E-�i���#��,j	D�4qp!M�����d ��V8���x��Z֤O+�I��=,�0��8C�'~�l�:��zu=v��n�(��h�,��0L��0��(\k$�H�s��oޮo4`��E���L�#���zݸ��,�Vi��J��,ݷGm�`��mQ�g:+���} ��қ�'��.��e�����,��F�-t,� ��>�jI;���mo���PJ-(�o�Y+���ܮ�%���ѲF�7P�u��*+�MᩅpJ<L=V������?j��ӵt����vV:kLյf-V�Ve��W�|Vԭ�4�򶯝��_;i�WK��^/o_n�ե���q��qq��1�\|�>kƵ~j�����_>�����/�j�_W�Zc���v��k�q�sVV-f��1j����\�V,�izV/��8�b���.+�[����\W��a	TO	_g�G����xJ<D�+�5���/�t�M���i���x�\\\_W4�ⱦ�[a�^+�����.+��1X�1��ݸӋ��X�/-Ƹ�k�qqzݺ��b�Ƙ��zk��������㶱q����.\����yn'�|���I�>c�0>N#�4|��UŶ�J�Z�����5kM5��[q��K�Ř�,��:q������o�m���ƻ_>N��O�3:E�_��㚷<+c|��s���n��B�������Si����g��w��׷U=H;�����(��䋥�"���9㵲v�D<Ｈ{��oo��>g{�r5P�|ֻ��w�59z�̯�[���|����w�0�7��j�6�YW��|��=���!w/�k���{��񈪪�t�7���������b��"��|w�̙����>�򪸊��}����2�3;��{����qw�N��۶�:WN�x���;�:xOK$��Z�j�������	����p�C���SAä�,a�4�i1[]]��0ĭQ��35�ߑ��������8��!��Ȼ6P�X��}��[4%�_��۵!ʉ��al���$�/�������w,{��݋S�M��E2�z6"H�h��T0�����Ahb魴��ʹ8�:S�����wxnNY!�qB<9B���F�_b#qeei��ܫ*cM'��~���b�Rr9=��n�n)���|��!�E����)��J��n�:Y��0æ0N���?v�T�_�J�L��ft{I�I �x�)D#���A����H<1^6� �Ë�!o�+��l`�������F���i&ra��h,��ZQ�-[���������!e��S���*�%_-���%Tﺡ��6��1"���1`�il��0������جa�F�E���I�2S��4x�mY�UG�\�]$y�o��kh� �b����u��Lj1\��h��<��Ң德�_�Vڮ=����b�PãN�)*L,e�Q��!�Փ��~SÎ�Ӧ�6����pDL��	�M�������7.��Bb+f�ʭ�\��|u��%�����(�]�N
�-^G���da!��'Đl��f��״{v��766�LMW�Ԗ�[�-��,����� vZ�:�N�Y�+q]�J8������ڑ\Vsq	��v&��Q"�)%�c����H�����8�#��(�Ե9M��س�y��+�t����uHi��md���q!�C0b���6{�%�*dPi%b�t��Rf�$��=q40�w��v�z?4��.�_C�ࠎ�W84�J�6�8Hq�I�P1������6U34s�nM�uň�P�,��!��DI�iK�!�����prm�y��jFĩ�ʌ��\����C4�E)%cn�����GH^��N�Ê�~��lmҞ�t��6�=z�oDL��	��Î�Z�5~��f訂"��,�I��H`lh�*U��[J����|j��}�@H�1ta��#:��h�!#؛��NN�(��h'���u�s��@���py4y�3��F"� f#/�ȃ������6�B�«�zm��Sph8��������"�K:��lk�).H2U*�J�o�}�L�����s3*������"�[ e!�ih��l3����H�a��F)^ hi���Q�71��ZܯV�i]'米ڗh�(��HK����1��R�����7=W8ۊtqҺtК?��?D��	���J����m��m�бr�LF!(a��#�V���1�4�dal� la����i�P���<��Ѣ�P�@��p)C<����C�D�h�Hn�R�����q��栨��ǾNY埋�u�f*ْ���~�?4�Ɠ�?[m�e<S��#���)K43��E����&�z�[4�B!��u@�cLu�^�[kn:��SQNEJ�V�?)�N���S�:}f�2�p�40�I�h������/٢��4|��!�f��6�"`��:A0�.�kw̭l�ǿ�"��w	2Vʻb��{z��gơ���W-�}�r�����r��ˋ ��5�V���Zm��m�h[�f/¨Y�29�1��'j�M'��y��0�6A	�!����L�Y(X��<�Za�)�n�n0^��'�A��ִ~�q=�n�4By��F��<�|S'm#�yښJ������G���1��<4�b���(�$!���:�D$u�(6@�̦���Gt���S�mh��c41o���g�A�/U���l��6�"�"$����J(1m��Kb�Ͱ[)v)S��F쎕����x{Zx���Bb��T." r�K b�|i��W��O:WN�z��:a����"'�L9�L�G��(F�6��֋P�k�E��h@�0RÇ
G�є�IM�Q�<4����Ϯ�t���JZ[m.]�mR��	 �	!��9J@�)�BJ֨B]6��e؎�:e	��e�b�/�(l@,ġ)�DF3����R�͇�Be$T$�(�zv��h���˯.I������b�f�ͥHg�������/T#�%1b4�&xe�M����w����S�~)>~m�J�Pq��i [Ub��1�xCc:��r�FYb���c&A�� U���(!T�W����%�rl�Ȃ�`͌����Bd1@�Ci�s���Ȉ�ѱ��#F_��_��B��]]���Umd�����{��z�y23����5��QǗ1�}���xs�k���4�X���
��p`lehJ�D5�l%���QU�_wۺ]9m/r�50��$Sn����j�[vӥ�"�S��h]M%,���E�0�F�$VX�6h�<l�����"'�L��H���&/�h�Jߧ��PI�IH咏��1X��)�l��zu�*G�4�3H��C)m�&�H���/"�&"H5�#lV2���v;Z�X�L h��Q�H�h��d���vheP��ap�K��1���F��#��8��"j���D��O3BOZekC�m'{"-�p� �Lz8���F��B��OQ��O�(�nI�J!X2�
Fn���h��F�ѡ1�K (f���<�Z�Z��m>t���t��ߞ�c�o^�D��	�K�$�]T���z;�*���"��#����Vmalc�zn ق��L%3�J����(
a�4ҥ��?+4�6��$\'@x��i���F��)]8���@��)�/�c��I��IZ���9��r~�s�����N�0P>���rx�x�r�֎]R�ōLiۢ�6��$[H`ڀ"�(p�� 6��/�h���Ba�ȄO�ۡpD��:1leo�����H�p���,�X, �Y�2�����i��J��oc�O�;zD�:tHa���S�����}+^{��h�>����?	PI�I y��#a�r�ͣ��H��3���GV�a��0����RRQ51#�����GT�r��1"�aZ��$S��(�E;	�E�i�c(aH�K�V��#-��b��+EP�m�C���h�`��Z��t�#�-,6Z&7�����4�L�D#�Zץ�i�S11��#6&��ўC^�v�*-��m)<ݜ���ԡq��R:8]b�����w�ӆ�e�|+�^���dt���GG��NCl_W�Ǎ;c]��mqj�Y-��uov�Z�+�-Y�W�+jV�i�MO�m_,�\|���/���]/��t�Y�Wmcz����c�X�����Ŭkk-Ʊ{cX��V���������O5ڱ�\_��>�ߥ��VaX�qj�}\Y�ڱx��:l��N>i��\|��]���/���O���_��ǭmq�L_U���֘��/�i���<k�j�.1��8��];k�ǍiqX�\V��.^�u������X���4�]���ݸ�-ƧK�Z�z\^�����cX�6��qq|cX������������q�b���f�4�Ƨ�k��N������Sv�[\oV���K��J���iWW�Ū��Yo5kK���i��\W�b�^�0��vD�jt�W��	�z��~�ק�C��,n4�%~5�G콟��Ҡ�$r?v<9��6@A?V�`׸r��YV|����B�q�p@Oĥ�NO��P��Ͻ~������|�ٿ;�$�[�LU,q�6�t35�͔�B0c�Z]t�������ʳ ���<AM�X5���LHn��@�䱣�c�^�3�2�sA!p��`a�y���C>{�t��lõ����e/�	�&�=?j�\o|-���+��M�{=�JXc\���m��?GLސ�hRO����L��Bo�k�ɰ�Λ<X�i�{�-!����m��YВ%kPlu�
���[hw���Y��n��d����%\�Qm̰�������)p�AԲ�+�t{�0F���z@WR��n��B�-t���Ê��l؊`���I�\3�1a+�1�_\��������o������?�{������Uׂ��y�Y���u������{W^���y�Y���uZ}�{��x��^���y�������+�fg�ffo":v�n�O:WN�x�Ǎ�<pDL�D�_ID�5[�FeJ��ŏ#4t������d����v�j3k��J�r6f)*��-�X�1��x=�=�u�k.	�ZZ^� ��۝m���K2D�940������ZZ�m����|�|�Y��4ն�l�}m����!˦&!�SKl��vc�Օz�u��%����&5�Ʃj�l!fz�LH����M�[{F��ꦫ.��e��Z����5���7�F�qn�V&�v��f}���_M�Ev�6�fΥ^e���1�Lb�\�3]Bj]���1l]�K1	v�Δ�Rj�V�JF��ڤ,5��J��Q�A��a��e$0*l0��F����>�w4�i���Fk�I���Cn���\YpZ͆�<>���~�>�DDI�&L��"��p�e�^��-%��m�k�.�s�]���5aT�f2�u�ٓ��фCeط��>Uկ>K���Cc�AC,J$�4��{k���ۈ!��GG�P�qQ����h��q��P��0�gz�iI�������ZR)/V�'���5�Ӏ\��!N����ȓ�5�,xy_� �Ʉ@A�m�/���W�FH�e���}�׳�����WnX��z��X������6��~m�]#pf4�sh���YK�.i���.R�����+������u8�t�ݪtqқ6h�h�����D�:tHa����$��}5fb�{��wǥQE8b��L9��B���G��%�J87h�@Jń�C$a�qI���9E�ґJգI��`0��2��y�R�=m�W��F@0�d&J�Ie�m���1ld��4Cl�(4mH�T�f��M�FB߹!~��Tu�Xh���"�>�fL��UsZ�Z�f��Z8`�wZ�vZ<����^dè�E&��6F���X���Q
��,
�=��YAhgu�#�|nM�SeB����ފ:I���2͐ٳBh�?���"t��~��1��T��1�Xп�<���jtV�Z�H�L7��+�dqmD��@�2'�-��Iu���9�1������k��B4��<��o�{��0��T�%�5�'@��}����Y���f�����z>��?>2�+����vO�pF��T�Q���]���P�2ƕ��"Op���A֙Ƶ �.��d�4��:n�4Aip�cs��*������Ն��a��	$N�	�N�n�=x�O��t鷭�~t��L�D���u5eV�D�\���c�,h��s5��X��u����R���@�Qd��J^���#f��o��u+G ���qA1��c�����X��\�.���l�"��/ $!N���B k��UX�� ��0�ы���-- �kK��Kq�
LD���J�j��h�Ҥe�д2�Bو���Pl�[�o�C5�@C]D()�x���d#j�L� T2e� 9<+jP�smഇ�k}��P�3C��ȥ�GJ�]M+��cǮ����N�t�4"l�~8xD�:tHa���kٺ�!I&-f\��dH�H�,l�_���"��7G�8=�i�ec$��v5�c&�]jӽ�0���$e�4��6&�uխ�Xl�d��Y
��[Sv�LX�u
�˵���tf��M.����ؗ:9�R���DU����ɴ���������+���뻻7�f�կ;vc����H7���W�c�6����������4�8iC�1�!(�W�LMQK�������M�I��ڥ�����:�9EDʻ6�WN����s!�H����`24�:		�kkkJ�T1@J/���Ȇ�9�z& s�PD��U`Y%�86:O�� �%�mVH�,s��B�
4n4iȬKQE'�<�=�3�H��<TK�����(��t���k�o�]8��tӧM�6������&�ӢC>l�������׵�/�A�u��{�4�}�^^ߟ]�g��5I����p5Լ!=�ӝ�Hi��=ML���ݤ�-���Z_O'�6�y�H:�_}v��ʏ���gOm9=�.����Zl�}��Op��~։]�i��{�voN��Z`�)�j����S�;���Q߳��>c4_��EQF0�=	䍧5��U")[�E��w��X�#��P�#h�-Ca��7Ǹm�8G�JL�4�MXVƚ��:�Z�<ۈ�D-����ֶb�k��N=v�#����ș�鐆�0��(���I$�<�I G����\�5��=:�ٹ�r��VL�r�����
��~(Ϩ?U�^�������Q�R�"Z\�!�!1��u5F�P1B��-myQ�@ic�Ȉ&tCpD7A$%y�ukf���ǯ��9�Mm1ۤ�ۍ����6~?<"`��:$0�-UU]��)�FB���1�I4%ُ����Icr�PX�H���W���R<l�b-
�����<�f1�֔+2O&��$!��T���
��4j �u�<ԓ5ND$�c8�0%�S�"������s&�v��[�\k�e_k�*���T�{4��ЀQ&��6�][���Q�������-��~��t����q���������4>g7}���$i�I$��D)�4a�`�"��J�zD�~�Cb(���
��F�~z�~6�m8�Ǎ��>v�D��!�C����RQZ���r�~��1�cM	C1u|��B7�4Y�A@3�v�6b!B����[N�l�ѝl|�Rv�"z�򿝵��1n�������;�'���y6>#4d��,�ͧ=����"�I ��G@��R�B�J���G�qf�A;��{m6k�zXbi�[& �-�B�
u6mYi�+P4mJi�E�ѥ$�����\���%\I�4HrE��C�6��bhlF�pڪEѤIa^QH��e�����ۯ~m=6���6�Ο>p��0DN�~��~�!>����\�Bd�'��s�5	.g�]ǽٍ��+.}��Dk��H+i,+l��\j�u�6=�?S��2�H����"�%�Qk֒Q�Ŧ����}=�[uض�,b����ցM�1��[t�Ć�:��-�7��V7ڴy+
L�hk["IZ���i'숆�^��uh|.� ���Yje/" E��F�{�y��qul�R]
D��6���
ɀ4i(-BZ%�7)I�G�Tb���HTO,�U�2��һ���K��Q�A�5�ٝon�S4������k
E��jI.��]y�Q�h�y���G��y��@3
��8�,�6-���x��a��t��߉#�(�#�RG��x����(h�ֱ<Z�%U�C�1�JH1v&����)Ru[�U��O4����`q9@��Zlm���R$�o�q<6���������ǯ�G���to��c�n�����aÇ1[GQ�UD��D��tc�I3��C�� �%W�d�zߦ���Kx�iPY
T��W(�%ע\���Y��(�!&h{�F��� ����)($�mB%`Y�q%IK���Ғ&�B���t�HI�O�Vb�2+B���X�pDC�4�v�^�)��M[W)G$	(�S ���J-,G|���-$�Ca=��pBdA�	��&��'Pbҥ����D,����#F���z=����>�~�+��-Ӷ5ں]�Kn[+�ڬ�y�|\+�-WK:W�VF�rB<8ᇆ��!Y�<iҸ�?4�\j�����n�X����+j�����c5v��q{\\\{�����ǭ3�t�;WK��nj�aYm��|�_|�~Z���,�x��jq�S�q\�����_��?+�c�ز�	\<RC�,�I<P�+�Lz����cUqq��Ʊ�Wmb�~_���������_+��qz\\W�ǭb��[����1{�c��.+��v��V���K��X�^1�\\\~cx��:kk�������o[�b���oLo�Ƶ�Ӧ5���Mi"lB�(�|��N�kۍ*��{n5Vx�[��t��\m����\^��M~'��0�L+	�
�<O5��7�k^�/��w���|z�H��;�+o���AQ$m�b��Ziw�<��ǋ�����yC x�T��ġ�t���r��P͡�i��pK�����7{�	��֩�Lͷ��:��/�6��[1'ZI�|��P��h�aE������~�e���R*���ַ��^������߸�*���=�{]��^ff�3=�+J���=�{[��^ff�3=�+J����޵��fe�g��]*�+����F��,��t���<l�㇏	�"t�µ2s_MW�U�rrP�1�I5:� ��P�k�'�m�b�6Q�j эB60!�l=:��l�%m�]iI���<h�Xb��G���m��Xs���� F����7���&�_��p���dy!�n��MS�.�D(6�=h��D�"��6�!���gy���#H�&��A8�:H�D�҅,���"���F��6k�ġ���2=ǐDD�ш��<��-�D�q���%	&Q$m�!��$�	G�#f�6�q\q��~|����_��^\\^B���m�>�֭��o$kM��41�c��5�h�����s1L�J	iF�$1�3#��V-/��c<���G�~�ն��`�RT�_.�c9w�	�����E��D�8���E#H�(����Z'��)!d"聱`ң� �bûk�"�>,�	�%"T����'�] Tice[`�)L���������1�`���Q�6��GP�F��\n�-�Y��n�t�M��znz�{qc�x����n+�ΖxM���D��!��2O�횇CTkb�-+��>�Yo����4�K5�3n��Jz�oDn��J�#�MSj���F�1��c�7�V���F���i��f����� ��֗��9���η,,�X6�t�u�[�5ن�\ٌ��Κ��rV��:Ҳ�\��o��m�o��,����zTpbepK���J#�Q!>u6M#C:t�QB��5�Ki\!�.yP�f�=�^�q�捦mw�F�FX�CP�g\VR�x4�hcce����q�t�oޕCX�RyZ:���z�o��������ֆ�-��UF����l���Ѹ|��puZѯ"�	�q��jt��!��/�RGĉ��f����W*�V9���zu�������ܿ�yb:W��H�T3W�q�'�T�eiL�g6qM�h�B�IC(�MQ�8x�t����ӢC� HJ��I���x ��
7�	@&a�c��	@! X�H���t�o5���i�" ���B�b���VQ{���v�qI�N��]�X�E��L�ɈڛF��6�E��Ţq�/���o)�����%�{�bB�]��!��.<u�`i���.�E��r��������kL�H��-PiE!֞���AY��4x6���Q��h�֕#J�B41a^��s.YS��ip����Pm'�!��]&�5�<4wd����06[ZF��i�J��F��� ���g��:5N7H��	P�V�@�Á��0 ��Ǎ1���n+�v۶1����ǏxD��!����=z�z�u�2�" ����h�ΝE���;/x8&�c{Zb�<��%b�DmC�-�e����Z�M��y`iH�����cG(���u&-�Σ%����c�&��R�ŝ��jv[�7V�$D�`�FV���wr����ŝ��U�cv�b��S$B�mo��V���TL�N!R��X�b�i2��!D*G�[i<�Fi��PA�7D�N�"����N�����&-A�Q2�(�I���ߛv��l|�c��x��GGr��cseќ���O�Q�NR����V��.~.:g�Q��b	""�J8R���\]$��ZZ���ذ�PO���<>�X�WK(f���j:dM���HۿY�nd�"�.�߹B��<n920�ۯ+s��}cݵ�8��I��H����X;8J��Z�<O.��i<�]ML���q������-`ph�FMDX�b�R��)
%��:�I�1�&��EJ�c\G:U��h�aSXݣl��peJ)i7S՚���ӓ�m�M�+n+�ͱ�O���c���ǏU���Pj4v���h�H�Q�A�~�ѭrTC�,�!\Ԫ�"͵5kh[6C2ʷ>>�b�X���� �@p��?�.�F��$���oy'�z�`ݴ"�ba,,׳ �,�|��Q�L���hkR�ĩ���&q=���Bo�܈#pL�����ј���YE���O
L>]q�c���<a�����J�13�	�e�Ш�jY��1��E���R:��Ƞ1��-�*����X���y���b�6ͣz��G�%)=��jp�"�-��N�ސ�ȾݿI�ج�>5J#m�qG���8/ݷ�p��&9�\a�T>X�o#"1����<þm�١IP�j�vPڠ����m8ӌm�n��v�<c�ǯ^tR��Vw\���^1Y�A$" ����![��[=m��F�']�����H�(�6�!���$�k�d�4jF�Z�4;GI0[4�uJ!�H���F$a��QV�|�|%a��H�@�� ۂCNyC-+X��\��_�tu�A�{ˣ:�6�1��f;�]�#йXDU7xq>��}������]���6�+$Vo�����qyl�2��^=�:6���of$2F��z!Lm����`l�e#�h�C�iǎ<m�����1�X��F�:��h�{��_��I�IqA@P:�<�iE44m��i�&q��J���J�#��"+%�xۣ�8��1Jj	������[���1!��r}j�W$�#���ziz�E���Ѵ12{y�ُ&p�����8����`�-�͉�#��~6�)mH��l�j���YB���u�{v�4M(�<�#IJ(+GSޣ����:0ۍ���6������Ǆ��ӡ�9��+���uEUDBPB�<-��#��R-��+G����y��ϔ|r)]�}zF�Ҫ܊:c���*ԁX�H$����Wau-�8a
�E�JK(TT�IH��C4u!��	���"�8��|4�M�ue,;�9d�3*����������Ag��0�	��p�0R@i�E,D�2Eg)H���+[4pE�tA�{ �dx�|4{v��Ƙ�[��Lx�v�]����XY�d��j��1kֱj���|�[V�K.��+���|ӥ�]>i����~^�k�����cx����3W�N1���X�7q�t�./�ݸ�X��q��yn���gK�°�.�%�Ū±j�j�X��m=��rޚ���t��\v������j~cO���f=|���>c\|�+�5_5�ϗ���cֱ�_��ⰸƱw���q�X�XƱ^�����cMz��V./K��ǯ[b�v��������ƜcN�����驥��Lo�4���5����q~v֟5���K���wn�c^yn�r�ZŞ��x���q���k����5����mޭi�*�kWUŪ�5���V�ƕf.�k���X��5���x�XO�T°�NW�TJ��~<����Y�����3X��P�X����������6z�1D� �n �A<P��ͥՍ�����
��|�(��Z�/��[m�D�'-���I���;swe�dA3�#��&Ai����d�*J��O�gi�������.99��C��d�7�K4�kx��{�ͺ�`B�7�]�%9��"�"�=cF��^K���#�n7F����-����v���5�\�|%�*e3p0eiu�ݥ����d�ٷ���J���c�	��lc��@pʪxy��/#�ZЉ�;��R|V������G*�ពz��26�v���k�IGu�}�~�g�ԇg���ݿ���9y��~ڮ�W����������{j�U^,Wۗw������{j�U^,V�w~�����{֪ګ���ͫL<6�m8�Ǎ�v�lc�1�W��ˋ�\N�r�G�FF��\s��Ks��cm�2��,[��a��]lf����6Ff�!�� �,n�����tDn�Kim�ƴm��f[�1մ��O3�M,��[u�5!��a3v���WSG�-8��v4edMEc��ٵ	�./�ބH�_gi����a�#e�me��d�.���䆭�ŻY]sL��;mG�h8�V�F�7^��X\�I-����3q�5Vi6๽ ��ҍ�ؚ�)u�b�D�5�m�0�����YN)�h[h��CA�u3x\۱���{&3�>��l�m���dl|;��E��U�;i]-F�M2�!��R ��[�c,��K��ͼX���L��.v����)i�6�m6�o1����9A�N9�a��6�T�֛�:�k��Yeh]��U�ͭy��Ĳ�)O!`JM*�%���b�������&����̲��!\��Q)�9���E�Ù�nf��H���Xh��*t���Z4�AE���oƈ��gVܣ�kg`�hP5�H�ICF�R�U��'E�930�\9��Y��=AɆ;Fխʌlv)4YD�J�jwv�F�!����;@��� ��|^̘g���h�6�l!B���%����Y�ۂ����xtR�kH�Q�x�x{:R���XIS��$�^:;6�m8��m�v��t���xD��޵�e/���������"!('��KF�@��,�I�F�(kv�E���w��FA' p��]o�()Z��m�!��AI�sh��cf,^�"��Ӥx�6܉�2($���E�b�� �}����bp!aVY`��#x�.!�z��/�����B�Q�2���V#l�$��R$[��8n[i��)1`�o\�������z4i{F������J6ӌq��;c��x�1��x��~�j�m �^�)�a��M��N!( ��&qB��P�	�P��3�6y��ċ�^�G����b,م�([7�ҕJ�H���kf�V��=��s���vO�'^��d��ʁ�8�2�f{y���L�5V5��N�{*��f٥*���DM*C:i@��"�|q����7��q�]0�:x�숴'hT/+:uaHfѲEfb�y���m�������8񷎞�c�c��׏%�Z�V��AD�%�eo�(��e([-����Z Vw��
bf�uW�9�a�cG	te��!�a�#rُ;x�&1��9��	�X���{�o&"a�lo˺[)&iJ�4Z4��}4�j��y`h� Y�1��R8J ��PC�y�H�>8p�]&�+�(cl{E�HѾ!��,=FiF�.�V,9��Jf���`p��tzm�q�8���v���c����u\2�!.��c96Q͚�Y�n�9H\Xݎ����l�(��"��I"��a�[+��"����T�}?w�$�H$��/A �1qG)�0$mm#�m��\��1����3su����6fцڃBmff����Z]]I4 :���D��4��>8����羾9����>�+�Y���M�Q]��
,�O4��,�`�}��P�4�&p���pnU�{`�[;��<Y�tl�*)O�����C��8�2�)RǋE��%#h}5����a��kV�k�"a�w��k�JWӈz݋Pd9l~-{áH�R�A�Ҹ��
�}9�~����N�xlzC|l�BGЯXp�ʳ��13*O%�9 ́�����RA�g�~~�t>,\�j�+��+���}�bC8Hlm�qǮ?8��ݽ�c��^<�9�=���>�?U�㚸:N�;ž�{^�x����/{_|�}�`?��	!D%-�J�D.���
GQ�F���KVH��])�Z��J�L�m��I⓽¶t0��b�(j�]=+�#�ŋ��m�n�M#�䍦�A���έ����]��NGD�џ������D9k��R<-�jD,r2�z��JΤ�"R �k�4�Z[6Y6��-��������nT�43��F&��x�ߗJ��ӹ�,t�n�룆�Wt�=v��1�z�=x�h=/�!X��Ӗ���$�H$���j@����J��#D�A�ZYh�P(8��*��)iɾ<R9����Tp�j��!�dPm�p�fHk��\q֘��(�s.!<_b��D�.��FRţ��r�0��	-���E�[;Ih�13K��R8^o��Q�Dt�A��^�͖��x�c�����&��]�;H��a�p�ΞL�L��i��y��W�6��~q��x��c�1��Ǖ|��uDD@�kF��P��Xm�rI'ZVI��T"��νbC��`���j1U��inVą�������";��[6��K
E���c�q��� �I�E�E�]:��=Ʈ��ȹg�oȾ�loC��!�E&qF��l���g��Ťt��G�.JE�#Џ"��vut�6������RG��x�%h�TY#0��n+�;q�c�o<c��xh��*:e�
?C�1��c�@����1�L��²;��bicǾB�ұ���a�\4�Sʣ�1p0�=�S���b���'�[P� *J9bV���[U]`Mp��*�Cm.���km{J;dK4�"���EL��21��YF\M�P�-?~�ء�,Y�'jVc��@��p~C�ը ��ZRJ��J�B�6ߕY�C���p���ܢ�1p������G0m�D��Ҙ���Hhb�͢Q(��t�f2Y��P�0�㨥��B:��94�����o�뙛1q�D��Q�K63fbU�MT,����� r����6�)�-���\���]��#A��B=׎"�f��d+4p�E2�)�n;q����>x�1���ǝ������)kO���4yr4�M��X���T���R%h�y��Exr�6B���x�U^GU�=*�l�70���Ҡ�OQ+�	<�[���mn�,��^���.������uJ��%4�W�by��?�N�L��%�����ʖ�4r
�xbҴ�R$8�J�5�"�Βb�A��Ԟ5����&-@r��!mR<Á���R3�����Q�<`~8xL:'���AC�!��E�G�<h�g�<Y�ƈ �"hDD��B�DK���"'D�6YB � ��EvD�4%��4"pN��t��0LقaB&�8&8hABhD���0��D��Љb"t� �Y�(��g�,�f�!�H"%�""tD�F$b&�M�0Lg8&ĳG$�4%P�A�D��a�4������ǯ�x����ᡏ�O����s�l��+�9�sq���}/��=�F�`�9�=���ŵ�#�d��{����H�:w���
��o3n9�t;��=��nfvd�b��3�N��k=��2d}%.����q��vk;�d�>�2��vY�|ܫu����9Ѕ)fՊ�3������ �混|/�o�tF�>o�-�d؍��P��r�W���ql���8��,���[�U���{��l�WAp:߁5-�կ�<1���z0�܅�IP�u���vq��b�d'���س<:(o;���\�]�7�3SH�B N]�-����+��LDn�z�!��k�Q2�!?-�պs�,��:y��*�^�<k}��|1�K&��=3s/��3�=��xMk�fo���l0@��A�v�Q��Aqǉ.TO;�-�0��ΐt�<�Ը@�G
��`7��]�"���8��Q�,��=��CN.SDR��fv��x����U���'������WMc���x/g�A>������HP���d1�ٖuN�\g"�Cp�ouniӯn�����:���(A�����y�oz:��7̪Itn+lx������t�ﾾ�Ý�ٟ)�������u���|��`��C�opLws;o�s��s3y������Z[�]�Y������U�Wj���������g�j���V���~�fffs=�*���Z[��(�����:l���<x����=c�x���/�kZkZkZM4ƺR�2�.��]��q��wz���M�~�{&�|�՞/�#���)]V���rֲQ�f��GH5J"H�:��?�c�H�h8ı�J
0FM��h�E�(�h�ajjJ��Q��Ņ������E1YO/q8��Ah�]�-֍��
F�-I��D���!�1l��QvAgT�wkHҮy��6��\�d�8\�'O�v��j�N>t�x��>x���x�:k�MB��-��e~̤3Q`��6�m6�4-.��R����cF��� ����6�x�D��!��k�F�横��p�!����[�4�6SZ���ܟ��ص�p��ak�Q�T*)A��P5�B+Nw�Dl],�6BF��J�TL�i�P��ב�D_2!��j����a$�몄Q�R�h�@Σ��\�k�g;ӓ�죉�N/�k�u@��#&��[Ӭp���J�6�61�q�Z!�1��oD�=���)l���<�m1��m\iǮ�~q���>x�1����W����s}�+�ݽzBL���q��͋Fiգ(��.�˷#D-ms��3f�������ֆl�sk����e��5~ �	 �C�oJ2�Q�\WB�mBg9��0ѕf�u��i�y�l4	��Y�eBė���g]٥d	��Si7*�7IT�2��Z���ú8�70��`8ظ=�?;�΄����/��y5I36�l��e���F�M��(�i�(Xb �8�D�T#������6]�AF��F�Q����b�v�⁵<��p@@6_\�FԢ����@�D.���"F�"Fl�q�8qF�D���?p�|=�����%�*�����E]קq�l�jxpd�<3�:�ќ�,g-xh(�ѭ�ե�)HQ��z���Ɯ~t���X��1�y|�^\\\�m�'�H6�I�X�m7D3�:�A�BM3����'F�1���ͫEv
4��R���6䮚�����-��cMO��ٛF�a�%,2�֥��n��V��&rU�M�����.f	pգc�g�E�5K.��+8�5�P| Q��
���Q[����w>u�6�3��rQ:R_���?pg>X�.%PYC�˅��f"e�&�I��D-�����!q�l�٨ Ѳ����4�Y8��O8ڸӏ6t����?<x�<'N��w�Vww�z�z�K筰�<
(x��6��HDAD��Rp��4�$�e��nҥ�p)8�F��#�<����	�z}<���f����3(�A�5
t��ռjU��gz��c%r>yx��q��{5�d�H�d���l��lp�G�$Ṁ�e������r�q砵K�Ҿ[0��7�E&E��ұx��Ka�$6�����A�T+ gH�W�4�و��Z(�!f�帘��i3��3��F�ɧ�6Ӎ>tq�q�6���x����Ǆ��:w�]�s��e����[�hkݷP�"���X��$9zp,GM�DA��C;�8���GS gT+(�voj�"��[��ZF��\���P&�O[��dCZ��Qm@�2MKKe"��Q�<S���n�4�R��c3�.��չ<J�@�(�B����o��o�u0����h<�&W�[Mב�KA��[F�8�u��A��ʀ�E!�E��0앴B�q@As��G[��w��k�ڣ�;l���rx�O��N�v��j�N;mӷ�>x~:t���x�:Kk�_n�(���]ŷ�Ŏ�L�i!��"'
Aoz����b��:�ٔ�+J����>]�M��M��y��ۈ�È�a��F�4��O�ү�|��[[��1 ɜ��7CD%������%�]���F)�F��������r\&���f���Bif�}��#�\��2��L�2��K/0��C��"��x�h�I.��'k�`I�P�K��D�����u�t�Ғ��а�b����MQ��I(�<�le#J�M�R��jS%��!`ͬE�YcDV��$�	޳$�F# !!E+Rh��'3��n��L$_���NY��vص�]�/��-��y%��%f�J��0�GgWq�n�8��珞<c��4~�k�]� ���a�b	 �"  c �Rx�PyrL7��G��-���R�	�����%Ty9�1U�#���W��s	9�oI��hk�Z]:�7#��"�.�P�\(pYI��y@iV�c�n�kez,�a�GV"��B&u|�E�}�43︬����>!3��k.d;����M(l7�o���t �B�Z��	X���[<�EŃRJ�äL��@Z<�L��1�[6��loe��{���Z��0��N8q�q�6���?>x���1�����ѣ~y�5ډ�q�q�d�g��" ��"�W��Xm+$X3E�ͦl���4iB1@QPq�������6m��Z��!g�#z��죧N���3���sk!�(EB<B��gBB��J��J)���:3�|�V��6L#�&T8�A"gV5h@��D��0�Ԑ�p8���rm�Lݒt�I~K�(8xC�z�#�ي&KzdDjSՏ�M|�nu����4�R�,�g?�<t��Ǆ��:t~�?ПT�*��V+��X2��d�1mNJܷW�D��\�qD�ǆ.}3Ө���� b�8�=?c���E�r&���4q�tQ1�qA�!YG��b ����&l���:ml�����6�G���3]��t)a'J��4x
3���:�*MzrO�ֽ1-a�cPp��-R3���@�%�rk:cˑɽLd�SQ��M+8Y�~8~4&��w�؛4P� � �ࠢ(��G�/ĳŖx�4""&	�A�b"pD�6"&I��� �!�DJ(��&��bX��`�a�D艂`�ı6tN�(D�"X��Ӣ&6l!bhD�:""U�
6&�6x١4CǤ�x���DN��af��b%�0L�t��f��	�(J#'�&�'H �� �&�	B&͈�:p�Ç��<'�(��E��ߟ��Y$�;Jd,"k���oq�N��2**8�g�m&�|�H�I(,a�1 n..M�X7��nmٝ|ɑ�سe$c����)o]�5dc�ya�{�Qdj�d��.��������C�Y`(�z�߳_ݏ��v�O�Y��%SHGL���ulX�њ�v�p�C�"}�{S�J�FI�w��pߋ�R�������5�m��׾�fǍOF}����|u��I���241�OJ6J�Ҟ�KC:����Yr�,��>�p"��B�A�O���׾�w�ؠMp�3�C)a�m$H��	��l��wP��(�K���ѩS��!�(��}st&����Ksq{K45#1.4R�	���W��j����K�#�7Y㯪Px�ו��_�N�߻��;����ګ�in���fffg3�Ҫ�Vե�ׯՙ����{J��[U�w~�Vfffs=�*��mWO�t���h��q�n�8�xǏ�=c�x�o�ꈒ-M�-����h]x7lk5M{���ձ#a�MvŚ���S�.����l�]Y�@eJ3Y�K@6��mj��鋩:m�SgKt:b�]K{BRU�I��H\�\RT��xs1 �࣭u�
�X��k���Vl:�t�1�v�%��$�k��u�,ה��,Shk[C�J3F����e.��iu��l������!�n�Jh
��u��]��7�.SM��+e���K3�6�mKFm�j�[�Ӭ�q���W�B\�.�Z�fj�B�n�e-m+m�[�05	y������-99��f������]*6e���ɬFmeCjKn���\^1�3��V�~!�b�X����C�z���i���&��P&�n�pV����a�`ĩ+Z۵���k��R�˻[�F���mf�u����ƍ�8��Y�
A�����MV��f�`ݔ�[V�Z��b�_[�Atr�I�I�Z��>=��#KƑI��!B8�'���Յ���45�r
V0�<z�����1�tQ��P!�	�06o�R#6���h�"�\:��R���,^��4����(�Hk
R`�(�>D��l�n6��tL8-��	h�#?}��T�e�m'���q���aytiĶ��y�VAD"6u���$6M/"JF��F4h�L6�4��ݻq��珝���Ǭc�y��L.��A��j	 �	 �B�J%�7��X�@`գE��%�L�����HÊ�픱qx�<Rᇆ5�
��6�F&�$����x����9�'}�#\��#|<��=7	h�s�`3za���U���(��W���:�<���O"͢`�$)�F#d�����[[yQ�24Z(d!i0���O#Z�N�h�l�g)۷�8���Ɯv��n1��v�G�����x`ѾXԕ>�Mc�9�Y�:kPDADB:h�
H�o�h�p�b�t�2Q�"�\	�M�!Fb���#^�C8�&B���{���	$���}�ɈZW���l��ȉԍ���4!ƂI��i���*���҂4ݮ�llt�`Hy��j}ʋV��|gX��{!b�)�G���k��'
5�[<���~$�I�7jÄ������d&� ck�Jh�GT��9�H�\E_�#F��.�8����ٲ�H� �f��g�����Ǆ��ʫ�>��?�h$�H$�A$F����,<�%
��.�z��������_��� �J�m~풶�m����t���_{/�^�~M<B�2��ŇVHRL�������Q����-�K��F�ib�$����D�f'�\�,���C9\qJ���8a#ʄ��֑f�\���t�	Z ��i��A������<Ȇi�&�3t�64�S$&�J'8��nm\i�m�v���<c�0��<xN&�
$ެ��hѺ�5�\�;E��B��TZs Ta��J���m��V����(��M�>TV+��_���~��5��`�Qa�=j�T��	j�����ش�8�D��n��X6�(K�V[���}�ꉶ�ǉ�P��CL�S=�3�����!�m=�ɷg{s�=ζ���`����p���#�\7GK��G��$�/޳�K�(62��)v ����D�,^����J��Hf(Ӟ���r'NJ��'�t��B���(�h:�2L��ӆ�-B6Qhc���CJM���T��k�����0���G������"AiJ 4k���J�DH�7[���~�޵����\���`�%�����2<@��IF*��D�cclti��G�㧭>p�j�N=m�n޾c�Θ�Ǆ��8t����ֻ̭��3��ɝ�sz�d]T�s7���(p3�
>ǡ�釡�Q�zow��A$@���I��%�m�ۄh��	.Q��w(ꍌ$���6h��lr�4pgT$�)Z��0�G@�cG���VY�A�Ѥ�zۓHa��J6b��ц��9{�q:E���-,�C*��7�R0�HdNkS�!�L��|q�fC���%�����u+c�)D2���gNQ�D�Fԝ��I<4�d�m+ͷ��QD����!�d��D�CH�l���rD�,񸈂!�h�g�A��K�I�D0)�q�6�o��x�?<c��^O�/�Fܬ��3�5b�X����A���Ppj�6�ƜD2 �,64ua%�qB%*Ԓw����)H��re�s�4jT��:3Bh6a/�"4rA�!��W#��a0�P{�	:���Z���9m�L���<�ƎI+VJ1(��D�C0�%�j��G=C��G�G	�6�s��Q��z���zn.*�1���p��f���w�S%m�2>�x{�7_��JO�=mr$;���w�`þ��d�']7<q����G�E�<��Q#8��>d�4�f�#exڣɄ~�u5�?=���'�X�m<p�j�N?6�۶?=x���Ǭc׏�暖�	q�FSfA ��0���F��Mж}^
� b`��1�B�4���S`�M6641�0����T�ӳ��.y��m��M<h�K`�D��8����r��/���5�V��;+jXVH4�m���!#L��������/d$9��t��iX�ў%[�nF.�4�x�X  p>��<���F�`W��Ȅ HCՔO�����-)PR�b6{��G!m4l�+��A�R[5���߻�^ҥ�,��Ġ4x��d�"��%aGP���~��cስ�@zd���H4PQ#(��Ƅ��<t�xç�	��t�z����J҆1!��&RH�1`$�]o����?,���6�.պ�6ٖ�d.�!�������dg�=�6�L��8K�+�jA-��V�f�2k�7m�跋��J;�A/u֓u�I/jJf�t��ɦv�C.9���6�d�u�[mL�c�{�s��2�*�@�q��(8���.t��ʄq$k
�1u+Pp�Â6�E/u����q�~���\X�cŏ��g���Qt�ڔ�7嶍�X)F�)!���LԻ� 9v�G��� fj����PqZ!W^G�_6C]�T�����ؔc'%�؎�δ��:̂ڐ�>�����c��S%�8��F�q�s�یi�Í��8�m�x����p��<xN�zL�~�,���9n����=��A�y�I�{���%h�G����p���J�Z!��H��X5���5GJ'��ѤZ���H4d ����%i(�o��m�m���;���^�^ګ&���cg|�qma�li�s��i&p#��y� ��zM*P�s��1���@4D#�j{o����Z���F���z�>v��>v�,��6&� � �	�
�UcLclm�t�q��DK�B�D؛����N٢�ACb�Ei�4&�M���Y0L6`�&	�`�&�����t�B$�DN��agKM&�M�����맮����ݱƘ�cیa�N�(A �"'M��8"`���:pM��e�I�4%~d��: �A(J�f�M8l�Â&	Ҏ�����7\�a�O'Ҍ4���\�$����\{���J(�o�W���T�bF(l�a��E��v3�<�7��/|��_òP��{&j�6����A�ZfS9�C�c8bOcQ�7G8y��C
m��~��,ߞ|%;�HmBK���-�kOۮ��~�����؝�{��;Rn��W��sٙ��}J��[U�w~�Vfffg}�U]�ڮ��׽3333;�R��WJ�n�^������J��]*��4Wd��D,����6���~v�=c�~n~k��DA�|(F�(��J��Jv�\ �ad��6Y��h��H�"�y<�م5�A,5��s/��㴅�7��{��ǒ�n~� �z��q(�\G�e�]X�H\'� ��g��yn��"S
5��+1@x�� �laf����Hv��L����/�����8y\WKV���R�B��J�������NM�m�][Í���:h�����<xO��Y����L�3e���b�X�I��{8�,�hF�ճ��-��m����[�&�X�|HP��z�jc��ۏ2����ُ��������7�3���="�Kd�qf�i�-.r�)���n��f�z�6o���3~7�ylm���g�
��K��h���k��mw�i��9�t��u��PI�
\E]��m��o���y�O��x�|0,�@�41��<c>c�1�����}z�ֺ�}mL��]�J�`��x�-"ǭ�qPţ��bL	2.�f�SU��4�ͳ-�m.�a��~B�7��sm6�m6�1sA�
�Em�m�X����Ա�k�u���.��R�gU�`�;���BS���;h��us��?1�>��H�D������R�\N����Y�f �I�'�-�dHa�:y^,X��Yl��בF�v��Y*B�\SR@κu��p��zE��C��]"�!}�R�k��Lw�L�&b_/���ѴQ"�q}���#��v�h��"�_�O�%$��a�2�.g�=���~�F�h��>ɬZ9G66B��??6�q�q�[�o[z���c�<'�	��r�E*�P�%" ��S�z�a�4i0��[i��b�-����v�UK���� �����(�j����H=f�C#&_Yqn��[E"`4�^8������8jGH���z�!g��}��TP/|�}&t�,
A�߈¿X,F:� �$��+-�I��XP�Tu��V"���R4��Q��-��L:���������Vm��I��cp�d�}jBP��m�8ڸ�-鷭���?>x���vǬc�GG��H.m����*	 �	 �xt�nъz=*F�E�CBm�b�d��%t�4�Kg�@��FP=�DV�m�ɽ��ڔ�����szdי�K:]�d}���s9�/
��$�8����ǥ=-���H�6��Ƅ��GQ��þ)J�ò�^�D�1�8� ��4a�m�Z8�[<� ��2���I�L<a���8xO��;�߹9��X�t-£uB��n���o�3�S�ﮞI�N���s�����S�ҊZ�����ݝ�.�&��}��}�(r^�yFF��`��0�J_�gǬH����'PI|�
��ղ+�A~�)8<���`C8�nU����^Т���PI���fԨ�z[ �Vu���l��=��!������֌G�r`�_l�$����ݖ���i��7)�qX���v��q��ŤI��h��#����%M"V^͍ϖ�{(�m2ËF�8v���a%�æԘZ�qOi�0��
!�)�TX��FE,��[�sS�����
�4Bʹ8h��:~<a��:t�a�B5��q��@6V���LcD3��1IȆ'{5]
.a�-��H��,i��l�V�z�������i��i��K|F� 9�Z���NI���9Ѷ�C=v��b<�]�ň�Z���a-�tܷ..J]��`lKį

L �
�W�/=Ϸdd��k���Me��r4�^!�}��~���T�m��Y�4��4������̴�jH�I��Զ�c2�MqR�Pui�\�i�j�;0�AI��F-�t-1���^C^�aF�Y.f�TA��p��Ӝӫ�h�0̔V���V���#���wj�L�:�G��v�	��(���6&\nU%-���&(0\gV��� �%�_{]ne�TiE���{p�nDU�6���?1��?1���^??[uB�4�1����b�X��Y�H��0�继��������^͢�jO
BO5�l�j�V�2��m��V�ð�)4f�j����2�/ͅ?
�vme^�ˋ����l����[@N���A���-�m���^����r�=�k̼qM�)8Q �Z���nQ�hp���Xz��2�p�!�x���#��Q�U��F0����8xO�WM?O�������m��CBҩ+����	�T��^v�n��vwx�l�Ch6J3�6�ӧ�Z]a��<6��J�[z�P�J'�0�
���y-C�4�����*6�9,yc��LĚ��Q�,�S��L��A ����U�:�#��с�%j!��z���K[%C~�qÂ��h��d��ilш��nE�^cd�F��GT�4��(���^�C	]���8ڸ��o~c�>c�Ǆ酒@�Z��P���J�QQDA|o��Z4�y�N��^^8վ�Y-[d�j��m��[U�0���5��
��2Y���y��g[}VE��0h�K8Zl�w��P���)R��י�x�:�N���qZ�p(Zꅵ��R�� ��}����֘d��LDDC$8���4t�羆�q��߲i�oY�Ȧz����51/z�|Ӹ�65Ϗ�+�o�v����<xO8h؛4P� ����aX�1�b�:q�+$6""`�(A�b"!�0DD�6&� � ��&�4hD�4"lD��&0L�"NGD鲄L(D�:P�t��Кb'DDN��NblK4Q�D�";�b"c��L1��1ǯ�U�ק����:&�٢Ĳ�ДFA��N�C!a��,6lD�Ӈ8"`�(�N޻�8p����(Z4�
tߺ�.t�4A�bB��_-�_b�.�u	�o�&�}���8���Yvt�ܧ����yz�U>��`���҇�v�\�4TP����w({�
�by쁌�秧&"j��Y!��5�DO1��6��޻q�q��h��/�jnH�T���8�0���Q��w��N�ln�I�]��7FV^6��e���Nl�w����g�0*$��V�p!8�۹��[�����s�c*9�JQ��n!v8Mϕ�z��\��D.�8� �U�N�!�vy$a�������HYj"���5�O�����ȱ�E���B Ya�:^DV�������M6�A?V���0�BZ��f���k���i��Q���h������+�Oٟ�z9��������WJ�����3333�誯ҫwwo�����g���WJ�����l�����z*��iW�c���mÍ+�6�<c�1�<tO�ǽ�7EO��/.j�{�3ѭā"A.�gY�lBމq/4�[k5O�i�SƷ�q�h�4-eP��Z�Sv5�[r�ɶ�K�W��X�/�hm���/R��3!v,Y���e�Ķl鍵ٷjJ֟Nǎm�ZiC\�W��4e�mt���a����������BbXmLl�,�?x:��ZL��ce��CKJ�K�}��-���Y�z��m��v4��m5�.�k�]P�u�m~�y|B���gY�u�P1-�̥p`�o�}�T���LD�f�i�Q�m�����6�[Y�K|x	��u�[��],��|��/���m14t�`�1�D��KC�TN;.�P�{2[��h��6�B���9���[�]���X�V+&�~R��]vjku�����X�)v�m����Dub��9���tɜ�Rm�L��#3K]X�-VjX��?[���ݙD�]���uݠ���r���s���k�hG����C4�Ov&���9��Z;���u.D6�n�۞��Ҫ$ٵh(�8�id�<������Vf*-�Y�@ы	[�����1g���7$�A���<���"���V��������ʞ���﬩"6�D-�9�M����� ��4yCm3�o��xф�@�)�6�?>z����oXǯ���ڿ�2i�)�S>!�M��b=�Q� �T-&��{m� ��+e�7F�x��"Q�uh(=����{d��R���h��������J��y�8]bx��S�<�jg�,q�eA��B"Y]2AP8�|��w�A�z{�����Av�%����|�731$�>E)4��Qh�'J�7n���zjX�:�1�n�4�8۶�,OǄ���<pO�IuP������l�6665��Q��Fg��m���TJ5�
:�)<QD���.�!��V��m��#�@p���yh5�Z:��v:�u15�w���3{�k��\�3[�;χ��Qyx4���k�9��'1STb/G����3�MS#ڥa������6����Ɉ dp������G��F�GQJ��t�#�c�K��?;X�~���4���i\q���pL<pOǌ<x؞<'L�&�cZ�թ�Q�5
���� H�*��e"�F"�
�i�hj�l�2/m�i�b6��Q���`c��H!9An�MYϸ'��~�����{>�|'�~]��~6h�fxO��Ξ�/h�Q�Q${�>�>���|;/`�媉E�-�h���Z<��f��ʉ4=���;�!�1h�$3:[\6m�t�mZ�FѪE���):�͐��ce�N��5��4t��^����t�~v�zq�q��6��1�~<a�����:a��Su��MU*��g��	pFB",�q�g�&d`�M��I��{�� �K�y"4q��c���[ @�9��r��-Ƥ�T�R[-iX���@�V&w�[�)-��)K��I���۞6.�pn���а4�,	:�o��T��TNmKՖ`��t��Ǹ�z��J�g=�x�y{�:�u�q�Z7d�-j�G��8�GB������y�ň�YG�!z�P�Z�N9�%�x;(�YGN��8��n�Ťl��z��(ڽK�=��mv|�%�(��B�� l�-h��:�Xs���+>ޚ���3���cn�4�8hᣅ�8'��<lO�;�݄�_�gd�aGH��e���=PZNe��xP�A���B7�vd84/{niEfۊ��H$	p|`7ߌvE�b&Y1;E�<o��k��ˈ������%�^]S�Q����������T1��F�G����ۙGW�Ի��pb1
����]��@� �,~i��ǳf`Y���[�*I2���d�Eۼ��Ln֑�NqyE��ӹ���<-t��cҷ�#s����o\W��G�:t�W��r7��鷧Wm���?>|���?1����M[�k�m�p�666����$��ш�����գ����&�������Y1���>i��}}���J�N^����uc>����@�3Y�"�Q+0/_j�}��:Y
�aD��p�y�[f�񤺈\F!�qz�;�z�!�����e�4���C%p�Z:^h�dC"!@���#h���0�D�
 eK��8���oX��1��1�������[-����(/���J1Y+B�9�u��n����MzմW� �y��G��1~������0�lt���m��qG�Hs�2�2���6�m�{�G�1�P��l�.`�+��s�GYF#���&B4�hk��O��!�G��4�<S��=x�F�M?=vۣ�*�4&��x�8'�x�<xN�ex����1L<(�n�A^�}!~F��ˣ�6R�>�-f�iD�pW�b����C�	]�UkqU�n�h8�mlƮ�2_�l��1��XX6�����mV���n1�-���7��Q8 �����s�F��%��?E���T��Ǒ��G�'��dt|�\i�da������[����h�I�-�6�h��h��n~D�����3��O�Z��$��TyI�Yf��k�x1�4�{K�l��[a�l��I�Ť��4��.s !BY�>?&͇
8h���Yf�Ϳ8���o���1Ǭc׏��~��nH+�1������-4R!q�jCzȈ���I���QGM3��zI��@͔�/�$�4Q��^ZU$	��`h�v8��!l͛�ܒNf��Ê9�ϓ�[y`�J��c�H�8La5�.�zG�����G�%X�ï��+�Q�F�*D���x(N���x��0OǄ�N�鶘a������U����clc�:q��cj���z���DDL�"%���	�&	�blM�(A
AD�DІ�2%��b'�'L
0L�0L����M�"X���'H �%%�"'N�"'DؖpK6'd�$0DM��� �Ԉ��D��8x������(�(��'� � �$!aԉ�ܟ':t�f�DN*�2^�Q�V����I�gk|�t������z��h0�$x�L��^X���}���:���Q���̞�e��C7���r�U;���IXRU��k��%�Um^���,j{X�w�lmncwP�|<�R�S�����9�͜}���z*��iU����fffg����ZUn��񙙙��"��V�[��|ffff{Ȫ�եV����6�ƕ�x��1���?1�=c�~~��.�ޚ߮�իO%uv����xzΣH����b,�a�F�4vב�˰�I!�$��u$��t�Z�E�� b���Fo4�l���4�-oCq������cm�=� È�g�tgBquY��2#�FȖ�8�a�Q����p�D�iZ4ӊM�R����ya�����J㍼m�?1��c�&��$�	FV��VrI$����Q��e�4�,�D�+	+�z"[��p�C�ڇ;]�{ś�J1XuI4o�:�T��h��coZnB��xS&�4�S4s��|T��w�z�\<�L[� ��,�{F�t�uN�8�gWm�o�z�;c��=c�=x��ǋt���<R"�x�q�U4X��"T����/̍���	|��Ы=_k��۬4u�VW8�����\^� ��ɬn�#DN[%��3SpT��M�
�Ю�#i�l�eƘ��4�l6����9����α%��ri�Ջ�&l���d{:��̺��u�+K�sI�Ֆ�imd���.��ͧ���k��L�յ�F�<Q�Mh �k��;����k�R��qQ���ڊ`%
CH�o���0�s�ߊ�}#TJ��`o�{xW�g�wsU�R���q��#����{ޙ9d	PE�-���*<���$��k��t�+�nMKs��L0��$�SJ㍿6�Ǐ^�c��=c�=xl��Ǟ���a�NR��R�Kl=����⪨R`sl�x����������puY��hy�C��/~�4�-,6t�i�ٰ���e��y��"5 }��O�I���@���غ)�v�le.�Eej |H�#(�du�g�$�����*�h�]m��,�闪񧎛xq�q�ߛx���<'���L���z�L���m��#GM�(\!<ǣg�!u0rl�DD8��4J�N/e�R��H�֊���)�(�"��ΪW��,I\2'rѓ(a�st@\����G^�?>ŵ��1�����!����
 �
R{PDT1�������/����6;��&��(�����m�U����Ήt�%--��p��!e�6h�b`�?	���	��w7��蹹i�۟wg}����M�͝�5խN��-�  Q}�&��ۈCቚ9�]d��H��7�X�h���i)f�%-Rk�@U�&�����S�TuX�.�DF�ތD���Sx!���G�5�S�Ōn�y�W�W��ᲊ�vaƴ���-Q��C���ϛz�x�d��,�:�dm�n�m�gWm�n�x�<'�<xO3�a�GꜷS;��MŚ��,hn��������c���֍�q�R2�V��Ǘ��� >������j]e��nB�mc�s��g�tر��D��4pC:e��&a��4��e��P���1Ǝ�8�����[��!�} !��s�8kj�X�.ql���Pqx���g���~~��)}yV�֜d��Ο�%ƟN`_��,[��%�Z!Zn;�ύ�3���Aݳ�XA-hj�hg(��A�#L��~�o���V�I�T��t\&��
�	`N|;�=�}����UPI�ݝ?�6a�ae���6��Ϙ��׏XǬm���-�����e�h x�.�OX��ĸ��7��mA�B1T�rh6�w&&a+4�D��loh�,�)C!D��#��./�qU�9�Io�/�P�[os�Kґ�69F(C:yt�� �#s��V�"i�)KUNL������q|����
�b����.]���m�<���d�QL�p7���H�H0��+�6�ߜ|��=x��z����^a��-a1TD���I-���6���h�qh��m� ��N�}�I4]�;�p�pJ5�~ό���С�O./�߮�~��ˍy.�� ��}�߮א9�0��ӆmz�\���xWT&��D�GF�%�h�[o����Y(p�����8Vb4y�O|�NO��1�����i\Y����x�'�tOƌ<aR򱞸"&s��Q�r[m�b�H��$��%ܫy�2�@ab�-���$������}�o�mΉ'�mO��ۣ}�	[a�c�:�*F��[R�d�xD1�����+)�$�A�:�ٚ�L�x�3Jelٜ �6�x6Je�vp�f�F�ƌ8s�P����:4�e��f��b<up�d�}p��/�}�lMjſ�m���m%HI���?��r��q�{�:-�S�rM���ѥ����Z��˵(���*iXY*�I*�(���&��UJ����b�J�ը��T���R�UIT�J��b��R�*��*�J��U*�X��Ub�UK���b�J�X�R�b��P�UJԳK���U*�*�T,UU)b��K%R�b��K%R��*��*�RUKUT�J�*�*��X�T,�UR�UB�U,R�R�X�P�R�e,��AJ�)U,�U,Qb�YQe
�ʕP��R�R�b�VR�U,�UT�UUK)R�)R�K*U,�T,�T�d����R�K)b�T��*X��*��X�T�J�*�*R�*���K)J*UYVR���UUP�R�YQ,�x�����h�T�K*U"�KB�YR�eB�YJ��
R�JR�B��J��*�K)P�J�e*�J&�*�*R�UP��QT�*U,�R��,�
T��R�E*X�R��UK*RʕP��RʕQ�&�J��*����E�*���IhYQ,RK)e�K),RK��i�),JK�����)*JK�%�jRY)(����II��%�����#h�����H�,RT����%���Qo�4�jU�eR,7R4��RYIR��K)*)*)(�Ct��%JJ),RQIR��J),Xj�h������J)-%JJ),�KiH�IR��%�Ie%�)(��IJ4�i))IR��%�%�%��)(���TRY%%���%E%E%E%�IQIQI(��RQId�������
KIRRJ))IJK),�J�
K"��%�X�
���%(�E��YT�J���(�QB�T(�P�5cUiJ%B��
*X�(QH��E
(T�R�R�R�R�R�T�EJJ��)*E��B�EJ*TT����"�
�"���R��%J��
�H�RT�*P�*YR�J�**T�QR�R�R�R,��**Y,�)*RT��d*TT���**Y*XT�K,�jY"�J��*TT��QR�����**E,�QR�J��*RT�R�R��X�QRʕ(�cLM14	�R&&��b��*TT��(�eH�J�T��EK*Y(�RT�J�"��T��EK*X�(�EK%J�"��J�T��**T�**YR��QRȩQR��*QRĩEJ��T���T�J�T��EJJ�T�J�T�J�T��dT��EJ��T�*QR**QR���R��(�eJ*QR*EJ��
�%J��%J��)*Y
�b*RT��QR��J�EJ��
��Tj�QR�R��*TT�R���*T�(�*,EJEJ,��B�%KR�R*(T�(T�R�(R��RĤR)B��T)P�
X���%*����K*��B���)b�RR��%))IK)b�Rĥ�"��%*�)IJ)d��)bR��IK
RRĥ������JTR*JRR�)QJ�������H�)d���JY
QJ��J)R��Ct��Y��IK%(RĥE))QH�JX)QJJTRĥ%,����T��J��(�)b�%,�J��B�
T)b)RR�)B�
Y
T))B�%,�)H��)B��T)
P���B�
Y"�H�B��T))P���B�"�
T�R)b)QH�K*JY
RR��R�R���E
X���%*JY
P�B�H�IH�)IJ��*JX��JJP�B�U�T��JTR�����J���H��IK�����,�)JE�TR�,JX�E,���E,���)E,R��)IK$��P�X�%(����RR�TR��QK%(�JTR�K%*)QJ)R��R�,�YJ�T�z�%"�TR�*R�,�X��R�E��R��JY�)b���QJ�X�E,�������sI�^h�JTR��R��)dR�TR�"�K"�)QK)QK��)IH����IK%,R�YK"�R,R��K�*���ZhX���YD�*��*�b���,R�%R�*���*��4,��b��EQebn�T���*���*�TU,��U*��U*�U*�b��RX�QT,��R�*���UU,U��e*��)UT,R��X��T�UJ��UIT�J���Tu��\�도ҵ�P8��O��0����&� @�lb-��5$?��c��?�o_>�O�>�p��4H���������Ϩ#��?�q����
�r�}h -�����?���}�џ!�����|�񯳟0�y��K�?���B�|��������$��A���~������h�
?�	�	S�?�Y�� ��G�_�����o� ��`/⁢��K���*�_�>���1�@}� g�y��$ o�A��������M$H�̄�������bB�6Ji}����!��F��1%
�������_���4c>t}r��L-�1����m~:�N��$5����G*$�� 9��D�T�HB-��"�H�e$"��&�6��E�'�����?��(^�/��i�+��F�"-D��5EQ�V$I%�YI KERDB�TI �U$���'�y�T�O�]��E���@}_���}���w��	������C_�����=/��G�� �H �}� �P}+����_�A��Pg��Oζ5�>_��?�7H=a���ؿ9�~Q}j����_�CK�a�&}�����I�;�?�4J>�~T�I @��1'Ŀ�ړa�~#�����h8[?F b>B��I �����$ ~o���@4���n��1~w2�@Z���V�����oI1%��>d H�K_�mW��۹�\,���@ j�!����)"п.�\.�PF
� g��ݤ�XS�b����R5,THk�T%t�q�b<,@���_��O�}���BO�ķ� � ?'�,K�pbO�#�_/�� �?�����׾�})�D���%�~��x�B>�>�}����O����_y��E���}1J��@$����Pć��@4#�~���H��_a�4~���7��h��/�|�x
�})��P}:B���1�_�`��b��(O�_�L~f�/���~@�=�D���g�T��P���i � 1�?����h����_� RK��E�_���}h�����#XPE�R�O�?RX�|%�hH�����d�PR}(41%���Z>����	�/�
Dr��~XK��zG����K��>៩ �I�`.�#_��?�rE8P���d�