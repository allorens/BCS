BZh91AY&SY�?��N�ߔpy����߰����  `�~wl(���UT�@���J`w�             lT�@���@���w��������u����;���^���zwu��k��@ >�x/�;�kB�8�ۥ�=�vƻ���^��N�Q/Z�n���R�}�^� |s��^�]&�jw���%��^�{Te��A�C���C��P�q�
v�mB�b�k�*@ �  n�]��N�:���Uk�(+�z�Ǽ�
��xz�ޣ�W^��[��hX^�����^����8  �0�t`��l�ڃ��Ѡ�ڍÝ�d���ףX�=�����y���ֽ�҃��y��  �a���zi�����:i��{�s�� ��N����έ���ӻƜ:=4i��>�     @  P
(�@ 4: @ *z�ޥ*�h� &L i��� �?ЈR�MF�1�MF)�����Q��A4hh�  �&�$�R�Q���M&!��`�dѓML 
�	�4MM��=#jh�P���OSiBM�*PI����0F�h=������&��>ci�޽ �c驈?��TU�   {�EE>�����0{cH���O��gY�o�����n:�r��A��Qv(�)	����a�U���E6J=����0Be*�O�)��@$;��g��O�����������[�������?������������}������4
�>�|f��|W�\%IX�Bu�vy��l���{���>	�^|W����_I4����1O�o<�����^}o�7������d�7<��m�8�����Ľ��ކ�������t;�F�h≰N�<6�<|�<6�6`}<
�x5 �.x<��A�������g�����o[�����\��8o�:b,���I4{t�g����S$D�3C�fh�dtg�5�S��%b���G��L(��jb�H��sZk9�����,I����<߽�w��{;����y8�g14�+޹��������'���8{Js���"�Ms9^1i����,�u�9\�_M�G9h}�g*���^1i���zH�9��\��}8�+�s��Y$�N.��+޹�ř�9C�ϹN�g���:s��\�r�s��b���#��I"�.r�k9�\m�ޱ_M�8BI�9��;�G�g9���c��SЧ�a�<߳<߻�Z�[��n�=�=� .���x������3�6� I<��pgdi��Q��N%=��+�3k��γ �9��></��՜֙C���d�+�j8��{b��-4Q��{z=�� ��ROcgNH�;�CI�5�z#����$V��Lj:d}�MI�M���r/|�܌��i�I�Z���d�v/E�#=�\ ��&�|��S��(�=�+f@���T^����S�X#Շ��C��U^���bj-a �����[QW8�����nkR^��Iy<{��{�=ҋ�#P����u���8�h�Ԏ�"��/G��mNx1<U?Tkuf���w���h}�M�۰W�9"�&��M�7:�*:9��E�*:��3"�9�o$��dy�W�E������H�=�|�_HI+�ЯAT�e�E�V�#�,��d�|.]�*H��mx�]ˁ`uv
����H������/Bt<s�=�;��z`+����&d��+�H���T��x0��.�P��`o��{�
z���U􏵺�}�NE�W4�H�䒤c����#$��R.��T��2rP�����Ԅؼ܋��OJ$G���^�'��g�NfCrk;6i"k\d�؞H�Ӳcy���M��7b�b��j�kD/{zA�$kr<6L���1�a�s����@��^���:����s���VF �$�7:w�A2�5�N�A�8�!�哞G�Oq����'�PY�^�=��Tr�S�Z����׉�v��	P��P�%
ԋ��f��M�My�&�+�q{��:�\X ˋ E�D�Nx%�=��|||�z�sEA��!�*'�O� �t@9�Խ��L%������5��0,A�� x�p	5?tyw dJ��Z�{�W{#���&#RJǪI�H�R>5X������r2t�'�Oa�Q�<�ѓ��k�o�:*2OH�1����}h�a��|g��[ƶ;ԏ�b�'(ϻ s�H�xl�9������q�����\�E�2J�Y2g��Ú��u>x&!�8�^V@��=��$�$z<�ROc���������3������ōV�k͇�M� M^�H���IX�&��}Rv�%S'P�(O��:	�O���b��qw�L=�J���VXZ��<��.�=k�ޞ�����ޛ�9N�����<٘<c:�8]$RpvM����3�_v<I��]���G�E���(��m6�fwG-_d��Nd�&L�.��0��7
�Z:<ӊ�ёhf�G�E�:���5�h�OE��I�9y��y��p�3��f/:�r5$Έ��2��&�Eۣ*�Ǥ�Ü����}$W�̮��ΣF��5��/s)��=Μ�y��ً�9���W�2"�ni$^:�Zy��D�39����ԑ_k2�﹑����ۗ����u�0�=��3��y�s����S8��ȝ�gS91��]�k3��&c�k9�Fj�	��Ok'�I3����a��=�g�9�f-{���U�D���E���;(N�3��c��fdq�3"5����dٗ3$=��6;|eQ�g�؋Tf�CG&��o�飢���a�FǇ_fh|�3�:�bGĉO���jc�A��&�H#�w�F�jg�a�3��4IO���\��4��wԃ�Ox�!�Q���]�s0o�dr&�NȞ�='��3X�c#==�ϯ�3���S�����E�1Lb�1{�����ž�3�gDo�b��b�ű����O�^�C��t�?�ih���͜���l��T-ї��2����c�gfq'1����}��t:}�z�����u�P�`y�/u����X�Vў���8Z������cȊ�A|zMo|s�|yw�m�w[����t��|wz=Ub�����p<���3��ޛ ���𳫆7u� �o���=�?��O��s ��?���	��C?�G/׃�������|$���tb1��B�'��?��_�S_���?�$`��nL�J��ni�����bǼ��uvlV�ƥ"jDm�G˦��0���r��z��r=�%���3h�;c��f
G�����vt��Np�?�T�`-W9f1�(\+����m0�s�?�L�0N�[ZO��~�'�K��I�Z^'�������Uy�}�}[�&ځW	�����ys���z�.�2uQX<��e���:����^纚��P�H�O�Y^ǠK0�rf�Ҡ�)M܃>ݱ9�p�l�X���6�9*'�o�=)�뉇J���m����v:��(f!��N�
r�1�S)��/\��!�MF������������C�[�bc� wqh�Y�:e�I���˒�����ї��jآ9{��g�Oy=��m54��-�ʶM��fW��ψ.�5�j����rN_�w����!V|��]�Y�2�i`�+�E5����x�ffBl �B(����Ŋ<�!gK+�o�a��Lu��[��b�Œ|m�G�岑� �2>(�Fπb�Uz�͜e2^��ؿ�#��}�����l�w9_ �*�O{g^�^�S#��,�������.j���W��bf�Ra������WlȃY�����\�H5���M�&\0�Ybxb��am����Nq��2�����=���F�on����?�[���Z��?B��>�1�<�R��Nf�_��s�qK��9������0U�9Dy�g',2H:��¬�m�mg�gg�L!׻Ifw&,}��x �گ3g�&���(og�w��g1���$.zE2'Y	�8�K(�t�1��0|���3��͜��]ۃx��d�ZX�׆����{�x%E�Ic����7�V�E����"\q�S2l8h0�awr���ʙ���9�Ҁf�|��8o2C8�|���wl�,5󋘛�ݜ"O�xw�ܽ�3����w�:�	soq���d�Μ�r���zz���[���f-%���qz��{��up+�'m�c�7���\����pW�0�.�E�{�d���^��ZP3��Zx����\��[�>�gkQ�{�=���F�N�m.&>]�r�{��f=Lߜ���|�ӯ��;7�|Z\�3�cE�ܲ��/�ǐksp�a7��3.%�S%�eWcA�����b�x�!�7��9��241�B�R���>��D�5`��r�����^i��d<l,�4m�m5\�n����>Ǎ<q�C]��Z��v�Bi[�:5]�Ʀ�"o��s�����k"�s�^F�W���T�{����e����[�s����#�!׳��a�ល�2I�K<3U*;g��:������/ �G�G��>��ڱ�e2������$�=mط[�z�M[�(ђd�Y3�)���s�o��]%�q������{[�i��c��K%�j��D��w�(�e�6#cg�|��O�<_]����]�#F���W����Rl��w"��%�Z�]͑���9�7���qv��v�����	�'+���_�|Y!�f���Nsϛd�n�Ns��&E��p]+/틻��:�l}��fu��]ս��7���$�8�a��Lua^�.��;�c�ǎ2����#��|��Nh��������$+E��'�ܗd�O?=�g9��[��������6zx`���5Z,S��I7��b��Z� ���vV�ݲ�k�g��&5:�kB�}�zW����'����}&��lO$`�c~�{J���,�8t��n
���W���w�����뻥��r}87���_�q��z��s%��OM��gG�7��4�	�Y��U����E!�gZ1d�"U!!b�%����#��-u����:�`sDqnkˢ�s����'ek��>��.nw���s���ruBq�5��fgx���s������M;_{5jo��3��������NrMrF�)V�&j޼X�=���@�$MJ��To��渎"G��t�5��i1�(\�d��Q���'����$��
p�c|�B<�&�[�zQj���f�U�ې�yL?-��Z��8'�����7!�M͕���#C��f,�7�գʷ���w陋�wg]��wG;��ngݹ�g?���r߀k���փ��g�j=ކ�ᄙ�"bk�9�E;��W�<׸�y�_^X
罸��Ne�	���P!�wu�^��s�(�u��֛s�8[~ս�߳k��Ƿ�LV�{��嘁i �9ި�1�[�r���9�H#+�����c�w�� �A�r�e�wr<2�j��8����w9��x�+Sq�8�F-�6�*ˑ7���b�5�qxP�.���]%Z�䘄?OMų_g��A�^�7nn7Qy�S�b�3n�ɋ��2��2�H\�ky�w��i�̻+j��{g\;�Ž���/[b��������ٝ�ǟc�[rR���0!4�śI؁���d��r�vNB�8D��1����ԫ�YM�m�����1�1ï��_�Q�������`��?����Nğ���t�#��@t�����-���L?����i�������,�a���2�e�5o��b�W`�S5��D��fe�iUvQU%mE[(�;��g�f?����;j:�>����,�|:���Ϥ�TQ1�G��F謨��Q�[�biJ�Gh��f�]F�
93S����8m��YqO�b��[]�pm�ٸU�wG���ʧ!�wj�Q%�(µ"����_�cL��L��$��#�Bh��j�c)�_�µ~�^�!L�z������+Sꪋ5U�bl[}��4xŚ�U�f�ri��@fϣr(V��h��������Vi��U����ӓ��B��_�8�,�U��F<�2F�"�m�H4�u�śƱ�h�K�E->q\B;��Vw�j��`4!eQ�vʣ��|�:���a'͑�J�aUcm����aM�/�̷��x2��LM\���/	�J��eX}��)��ym��$Fd�����D?�v�F��}3�N	0�A���f�"�v7sb���j]r��8��J�!��..*��1oF}r\�-!;��g5�j�H�-����V���P�e�����;�
���[Su{j�^�*P��Q�oj�X���&)U�,y>��͵k�^X��f�R�B�`K:U��*60{	m@X�]�%24�+ci�"���z��@��8�����P��6m�u��21���IT6Kq���FԐ�n4�cL�D^>��5�mH:���Sr&s!]�c���v\�ba~�P�����V,�Z�;��NYnvg8��̥x�*ؤ��TV(���>�MȬNȘ���(����vWodYc��+e�����9�Q~�O����&<�  ������׷( z���1`��i�����_��{>�yJ|�|�M�~����DDDDDA(H""""xDȈ���b"dDDDO��DN���:"&DDDD�����"dDDDO�DDDDD�""'DM���:"A�'�6"""'DDЈ����$N���DDDDDADDDD���sԫH�bI2�A!M>���H""""P�DDDJDDDDDA:"&�DD؈��8""lDDD�����"'���"&�DDN��4"""tA�&DDD؈��4"""tA2dȔ$DDDDDDL�����2"""'�H""""P�DL���"C�"""&
!�(�Q;#ggf�������"&�DD�����"dDDDO�DDDDD�"""'�L�����2""""%	DDDO���"""tDM��4""lD�""""$�"hDDM����2&�DDDDDDL�����6""'DD؈��4"""tDDЈ���B""%8 a�q�lQTY8�Sn���uuYgK,M����4"""pDD؈���&�M����$(ADDDDDDDDDDADDD舚4"""tD�"""�DDDO�4hѡB""'DDDN���"hDDDD����&DDDDO��" $ 
TAP;�� s !�U� biAhiS#�Q[\kpkn5\j�k`8�ϱ�����(�)�HE�����?�����c	�s����~L~?�7��x��hhhhhTk�NEr.�|+����t-=2�*y8�M�􆣅��Z�¹������oI��g��G7�		�
�y�zeq��o9ǽW���G
�W��Z���3�8p�Å��th]���������0��϶S�u6.�J�IKYIc��S���ݩ�6��Ϫ���G\�B$V��Lb�j��%��L�A�H���B�(�1h�I5���]ڥ���M�ac����Ϲ��8Ϣ��I"`[mR4�� �.W
��F*�����[ʜLA���*nY�E-#$�tWm!��9��|�Bj�JE�c��ۅ#�U�3�-q��}$#nѹ`�M2K
��'9���k�N,��U�M��l
RǮ�Y�X\�Q��݌6�����1mϡZ�2'+�i�X�f���"�%n��.%�_t�o&�k��`ݗWd[��H&�U�k�S�e��)h�5�sd� �,NHЬH����2��
*��� U��n���q�e����\Z���I�Zk"\�ӄB���$�H�e�$M��SMsE�n����!�����V6<l���"���8p�Â%�Ņ�Ye�Ye��""'8p��`�ae�Ye�Yb ���Ç8"Y�,,��,��,D8p�ÇK0�1���w�����+P�tG���G��t��	 )#��LG��)�"'5��y����f���\�b݅�刉V�U�>/���?��ܫ�a���ߌ�&�l&7�4�:B�!�2<;Օ�T�N�e/^������#��i�m�~{��n3��DR��/��h�^m��EV�p�AQzoN1�Z��m��8��'	�f����苲�h�:��e��E�����dct5)��aZ�\k���[�6�� cFp=�㽁 &�����-�x��Y�����,�Z$�< �1�i����>���Z�������Z�S+�lm&[�`]�Y�(;��]�Ѥ=��E{M�6LM���8c�O��E�Ẓ,����1�,�h��1�@5a!��f�.��Ѭw��	�ICR�{�<�4>J�P��\��%vJ�D�ňB�| �ɍ�B�T�[a։2��#�f�s����KLۍ���e����wY�")6��YYR��`�'!t,����ʤ�a�TUF2�lZg���[�[�s�V���9	\������c�se]t����:��sto�����I\:1�c�7J�x\��X�I9~[�ީ�=ۋl�k��`����I9�Ø]ç7��S�i���>�u'N���""�f�����j�7�'|'��������U��r7֚�aH��f���j�h|���{�?k;ӭh�d=�Mp�0˗1dv��yRq�SV;����C�N[��8�n�m��֩�57j�#y30l+n���7%M�J*[l�������Y�3M�h]�Pt6�mc.*��շ\6��UR�ə#�B�s������UDeɤ�+�M��iC�V6�Z8��g�I�<��}��]Z�t6v�a��9��t�qE�����Y)�a�?�����9q��@M�I��O��FՁ�SH�H�7ӈ��+ft�����UwEx�L�I$:x�DD���x��l/QA�D�u�m�W�hw�0�W��`�	�Gu��ZX��k��+D�ƙK��*E�sfT��!v���r)�X]��u�ƍ�^(8�)�m0��h�O�A$.x������U44>J�T=�c0�riwu�Dӄ!Bg�.o�w7�A����K�])f�Z&��ii���ʆ�v�
����'��������i�E����#7�-r���nE����8y�r֌o�D4x�Og��l�v������V*������J�16�g�!B	�g0�-{��1��HRJԉ�>q���e`���Ra��t�\9�BC���mӦڮDm-�.r){��~�N#�{D�P0��m��V�;5p^F�������W=�jb�׋�t��h|���sb�N#�x,n�8)���
����=&y�-�jd�6��fڔ]����M�jZ�]vT�Z4�v�Ɣ�U)����a,<!B6�׋.�cE�zt��-V�%B��稷��)Q��5A}�Q��$ȴR�&�Wþ�#Kh�GWB���o۟,�PUT>��\ZD�$r'�Da�[zG�l�ll4���zU44>J�T=�{vcPƠj`&$Lƍqsq���I$��x�0��f�����DV��}�9���K6Z�Q��{�M�oN]:��R1^Ѿr�ƌzE��,5XikR�U��V:�#�tt$U�(Gj`	����v���E�nc<�h��q��Y�ps�%%�G���e��?�e8����í�ј�����P>�����|��3�X�Fc<dg����ǅ�3��&<a�!��c1�d���Ő���"ǡ��f�c����;`�@�,l5�0�(c1��<��g�f?7������fQ�c3df3<C�yC3�6��a��n���4�Mcl�pf-AG��x@n�bl�����c6�d0�,f�a� ����б��٬�f�Fy�Y�C��c8d1��a�c��e̆3fCt���a�v��ح�3<��a�C�=0z��Q�0A����X�� >���Zo��|��9?��`��k�c�_�g|���X��qo-�^eo�ʯ�r<ޝ�{2��vy��}�tc�]=�ur�׵x����gj�wս�^������A�	�gň�""lٳe�,�̛Y,��(��DDM�6l؉e�,ɒ�,��,��DDٳf͈�f,��Y��,�İ��6lٳb"^����]���W�j�B:C&L�!BD��Ȓ�j��*�"�}ל��zI��B3��+�ٻv���9rTF�L��.�\b5ȏ�+C��J5ِ}t��.��g���ZRѥ�f\">�zӈ�)���K&E!$Ep7��Zi��D4�4��b�[Y�"E�/Q�d��7�S̓D	e!�@%��˴��t��ߪ���G��8P����h*N@8l2b`�l��~z?x��/,+^i�O��/!!������������	Ѱ1M�$�!�>4b l[kY�8��'R���e$`���;�8o0~@,3م����7K�H���j��>�*���"�������i�˶��x��CH��A���j���D5��;d5�0QL 5�
��ƄF�J4�4�A(�"��4
"��^�m�)1�!�G��:Iz#�J�&��tw◥����+,+^٘���ٯ��eN5���!u�ɉ�ɦ�W$�I]�"߿W��H�*��/�r!�i���)(�A�?�\�
 �&�h��#Yv�Y���興�����N[,�G��%WwuwJnHnI����z�i-[Ͱ��/%:H��o*=�Z"�9s��C�B��+�8<p�
󊨌L��I&M�R���>��zx��G��#�x�i��pd�&�0q����A�æw�6�L��׮q�$�MF��4u��ӳ����鑒�KA����%�$��S�	G	���^s�c���u�E�%b�S�曛�fs)DDDDE�L��0h;9��jwBK��2��F�A��ض�_&A�cp"C]A�r��<��SDTu<L,���:#�)�k鈗��\a�;`[I`3mN2��GUQ�Z���5�e�*���.|�H�AH9�[4�{�p�D���H��I>a���,z��#�]J�6�^�ɛ3C��ָu	�L@�+�W�*�%b�rV���sf?R�	���T2aj���DDDD\�����K���	����7�9ƧOS�T��w%�����Q`LL����F�+�*2!��p
�1(׭�F*G���!!bRb���T��&˔ف.ӀΒM��8�pwZ��C��p�}���Ie$5%8�=�U�ƍo�p>�M"&/*S��sgXTЭi���<3���ˠ��&.-�z�����ݳ����P��U|d�kg�$��Mݽ%�Ӿ	��������1�Km����m\^M
� ���1�?7��R��Ǧ�ԙ���d*��P�q�
)����-X��h�("��1�Mt�F#\q���]X�򤋯�ۭ�(�\h# �L�Q�H����	9���9#l��&$z�	�!�R<��z�I������]Gpy	���tԁ���Ruոޜc�F���3`ST��D<�D0v�|�z/�(�+Vd�Ug?o��ᙉ;-����R�,�u(�6��*�d�Dkň�?eEN����e�pP�i�[�d>�aS���������15$YM�OO
"""""���?��H+]�H,��gس-�Q��%��Ϛ�+�i=�G$zVԬt � D�Pv��&�d��8��+�`�;��.�]��:5��;H4������I���b�3���<!1h��"-�`��RG��%�-��V�j�h�:�U���4/Ǽ���]زf�Zy��Y���9�E��	������$��u�&P4�-�E�s��Ξ��x��p�y�R��ʣFp�B�!H%��t�H�DѦ�x��H�<�"X�rD�A<CHc�&�z�3�L����up��-�׾Q}s+�
*���i�rϊ:{�����̑��O�:�(Tn�z�7�)�vY҃2�J��p�|��L�k[,b�t�	q*k�N���6�ɦ@!}x�w�RR�`�h�K�CT�D!�G9���
>J�U�+�;���Hxɓ$!B 1��z%C[bGR4[r��}%�Aщ����}/7�%���24��%�gp����~�����ج��9̢�I݋Rp�ô��X̦�׆D�)�yͼ���D�5/:L8�����M���0&�2b�xu%�r�x|��L��8�#�b�!&Lz���'K����|���!�h�/0~w
�1�C`�P���_)螈�������;��)��8HW�i:is� ��bģIS���X}.ds����b�h�Fsmƫ2�\�q�MM��4���!H�)�ښ���RYe%�HĎ�HL���RL�<����Rk۹,q���3�U ���$���fSI&'�;q�8�3�)��f��H�7��mH��",#��p[��x���cǇ0���9/ �`:#�;���<@�;����4xx����`�f7�>f|C��5��f<td1�����y�|d1�2#�cZo!�1�̆0���3�@���b��7��Ͱ��i�3�ۇ�|�d3!����a�1��31�d(�c3d1�Ό�c@ð��6�������0aL0e0�P�+�N�Q�Q]H��[��S��F���=G<����<�t�ى��L��MOA��YFj��fC�!�����3!��2�f3fC���a��=@��e0�E�=0z`�=s�=DF1�6�l �b�ha� �d0�`i�?nC�Ȥ��[wK>]!�B�hO���X��f�&�x���(�>${�Q�YM�*)�[������>>}�c��;
3#=�U#�8�F�Y�Ӫ)){�g�T4��M�O��޹oy���r=f���;��l��iVL����+�+�+V��{F�u��d[̊=Y�>��]���Fƈ���}�G"���N�噾�����m2J��H���N!Ǥ�k�jV��SD��nH���b[V�z�UX,��ܗjk$D�m�^�:���H������c�Ř�0�D�E���$f8*IcD�z]j�
�V�-��vA��#��{
��kx�3�3u27gĴ�N����h�:�ݣ'9]XI2�H"�ۓvj�3�=��>�D�bj���Re�'GmA�@D� �"��b��n�	$�o�31�#M1w0�1�DY\��Պ�Q�'1��j1�ZԂw���C���&?����l�+qW$���5Fc&#�-X0B2�_��nq��L�����ɘ�͙��p|j�Er�֝=GM��~�,��<t���>�!e�Y�f͛��,�e�Ye�YE�B�,��͛6Ye���<"Y��,��͛6Ye�,�̖Ye�Yg�H"%�t�Æ�,��rx�|{�.�%b���7ܩ�:�T���'\A�X���X�Q���V8��SpYrL��xǲԩ�٘��-Lv(�i�M�̲���� 
�b'��5��C3�	��rA�nÛ�$�xx"""$��2W�̵dWbs������މ�1�)�a;M����X9�Y�Q�Ӳ|$와����%��N�)�эHq�TdtC�OIe7�����4��4^�F�DT�8R��)�G��P�rBk�s���8`�ġ��RLl�I�h�ɫ���iYf�h�H�B��qr�w' ���"���++�0�s���<���4Q$!���7��3w�����Z>J�u�Ú;ތ��!B�!�:��+��}�D�� �[`H����.q\;�Ng�rd��y�2e9�#���Z(�w�L�rza� �v���[F��$s�0�̼%���l�b��f�ǀV���"��j��!x_em�1XR<���#gO*"4�H�x��f����ͱ��z#Ǭ[��}�=�=�L��x��Y�9�~��B�R��ٲ�DDDDfL�gp��O�Rf��p���2z|�y���zʐIw�e/
5��]i%�a7 Lz$=�a�P���W��ն��4�]�,�L��M�k���&&ɞ���Q{���H��DCI||�>�x���ް�rzL��y�p�M�w�1:��e�D,ޟùUN�`����ci4Ѭ�iӗZxˑ�J�C�E��R9������o���3ǹ㫽g0��1��z�D/W����!B�#�_"#�|uoqg��ߘo��ٙfz���%Q���jUe5MW�Z,��5I*�m����u�:���oǖ�e+L$�2I�Xs�<&G��ۇ�^���0ck�\7Ѵh�H�5@�x �Y���S��ָ�㝾NӮ���')�gA��Ā���a�0U�#����|���z�l�RΓ��G�e`�-d2��܅Y��}D�-�,���ƚ�aZ�1����r��U0E���B>6K����rU��Wr��!�^V�����سY,���&���u��tDDDDFf�N�C[.��.�%���MXv�f�\Mm5���f��гي"�p�c8�#zO�i�E���ϑk|�q�F��H��Z�Tʪ;h��E�a5>F����i�|¶���\M[E!�U�	�V���l�y�7u�<�ִ�N$�3Ú��s�.l�����9|��B��lh�:H5G7�C�	�����3�O���|����UY��ϭ-.zx""""#0���������Ew���Е|�WIR1֑�ͣC�:�Z��dm���l�,��R���4��f�V��j�C�J�	.��c��DjM��ŴЏ��<�>q|}����5Z�9H���!Uʭ�
#RE 6�c�w�L��h��F�"�A���"0ҽxmwK���YN�O����A@b�9j�1�>�Ѿ�1uR��w���߫�%�~J�T=�6j�p�g��������t��.��QR}U�8|�IG���TYV�cWf�cq�� �4�-"��(��Ϝ�R�Rh\L5���dF��A�l��~9��G1"����G�֒<���l��7����վ(��A�={�ot�qX� c��փes}�;�f�]�9�0�{�Q��8���|��ۃ�&�[q��Gz�l������D�*WҍMRTK�kEfp	fϻ��fK�yؾ���c{뵤����㎗��q#�F��<�E��C�EO�c}W���h�KFU���Yv��C�d���C���KX`b<|����߸f�ÿ}�0�a�޳��	���$�4�ҋ�+Tu�ӦJ�
�Y��,b��+h�N*�v_D���ЛQ뙃3��n��"Z#q�*����I�f�-4��b7-�$Q>�����̏���ۼ�8��׻��2��p����{��$�X-4b��W�r�KZLt���I#�(���kkåGJZ/h�io��R��:d˝��I���9�8�}s���˱t�=q_Q�G4׸�D�U#�k���}�SNr��'C}G�W����t�J��v��}�����}�0�a�޳���6!�lF�c���z���Q:""""#3��|�p�g����|?qk������ɡ����!!�]#b�(�6�g�o�|^UH�� �a�oT���:dM�����+G��KK�w�>����?/.z������^Z�u�-�����h`fLT�D�K�Q�!�>�D/&B�%� \�\�A��	��{Q�q�flǏFC�!��c1���}�g�!�|�G����C�c�b�x�f�������[0f�l��a���ef�f3�!̇�7p�132�2���2��1��	��c0�,���!�`�kL_��@��o ��<"��=D1�p����lX�1�N�/V֙�Zj3�ga�eF�!��gHc1z\#c2��!��l�c3�y�1�3�3����i��L�]e�"����[�u�.�F�i���3D���V3k>����YK�r���jw緸y���e{,��U�׹�Ŝ�s�Aշ:���Ov�'���N}ܝ���!��狝�vqZ��UZ���;W�ӗ���^�B�j-v7��~ �GL�,��,���DO��8p�e�Qe�Y��,��:"&DD��N8Ye�X���"dDNt�Å�Ye�&�DDN���8YӇYf�x�|{�ᙞ3�]�9����	e�B�!B5���
����H��i��H66`b:(�qb<}�:�����]]4�A؊�Z;
E��������U5&MM�!�J¶�8l.�J75�*F�L�u0ё��#�BF��i��>��~0�uQg�ے� ��mTE�hAK6�]'ﹴ������\J��+�K��eb���Φ�4�iO�""""3.��I�h���.�tMT�z��qk�J��&rnѲ!!J�'�Kj¢[_0��2�޸����fճ��rI�q>��|�#�]����Mn��J��βiGO���1�6��[��=�o��o��&��3�_c
Ґ�Ჾ����K��eb���+H�u�9IO��y�WڌV���Y+���4H2�'$�X�pH��K`�`��4ڶ*5 B��"%ݑ�e$��KG*k	*\��X�tW�O�""""3;�����ʹ�*$�*���7"��ƃ��#��U*�|�ۋ�Z��8�kH�r�j�GJ�����}7�z���������:���X�`��:�iSMJTD������)QS�C��:k]f��F�>��q��9��w�b�,�ßp�3�f�<��stM�n�:B�!B5j|h>�ڻ��Rߛ��l�����m_QDi���/���|R��5M�+�5�\Mx�=�C�涍=/����m.���b�Y&�JUXE�/��(�a#�.�<�Ui��񩈻�>�=m77���ib"�M����St]�uc��wE�Is £��\�a������i�DHB�#['�E�Z�!������Ë��fH��`��_L��֥���n*L�9�k�he��l�7ES*���)q>�|?#6�f#����dqӕ$!�#��E;�E/�79GYk��~5I�M���Ү6ٳ��l�e"��8A���6fl߸w�fa����gwE׹z��Q���!B�>��R�4�eD^����w��ùӧ3�χG�ՈKwD���c�XiK`l>�����d>\�{���!��!����
|o�B6��o]MU�q-v��-wh�,�r#v���>ݭiqD@�����9�������}�Uֽ�ȶ��I���O��{gp����Ѣ��L�z������s}�7,v��B�p��}�CB�	#�4�Py�ѹ�n�t�!3H�J��m��Z�2Ev�e�Z�Ӻ�M0�!""35'b��[,JRı
�M2�Q�{$�W�U\��=�ZN�-)tD]Z����3��w���3!~�mVb����Do���?�\쒯h����Q����X�Q��l�vb{�'��}����X��F'
O���Q�4Fl\���1��Û/��x������
�睾n�o<Ӟ�w�����"""" ��
E4i���:�H����G���F��D�z-�/#f��φ�ӑqa����=)^�b�lo/�Z��6��>a۸|�O��6ܶ�����\��m�B�hױm-S�O�y�Y�KT��g��g���6�v]X�a]ѽ\��1!p��!B� G-uVtҾ��{��Y:p/zG�j�E��uV+G8=�m~��Y�p~�1����e¶���ۚRTER1�Υ�����:�m���W���i��5��:y�k8z�Ҧ�On#T�����?:}�?8}���3�^�9O���TU�C ��]yl*�ڟ`�SD�C興���:Ԇ��m�������V��"�F|ǰ�E��Jn��l�I*B�麓��?)k��;Q��6�T7�4RĻ�㋫�㑸BQo�6��E��}����������X[��Smo��F�;<2��K�28�x���~m��ǢX�`tf4���.$�@��pI���L\���2_4[��#
��x�.�W2\3d�c1�ì�X1�d!�Syeś!���a����� �a� k�[4����d3 Q��c:d3ƨ�y�w�Y�G�>f���>��0��>a�!�<ż!�!�[0f�0f�ap5�4�Mn���F6`� �(`ك6,a�\�hb�pf3�0�c��[��-�A���g��W�O���gHfC��l�d2�a�C���(1�2��8f�2���&��1`�F&ΐ��c1���c(a���c���3�d'�{��^��O����y]�loZ�W���}�e���蚥f�������ίG+���,�ً�̞��<R��L�����-�ܙe�'l�ڍʤ֫��Bn+��;���U$�f"��>�^e���x��.�����yݪ#��Z��uc~���l�;�ýS�o_y���X�=�ȯ|gw�g1�qI�v��q�[}��g{O�Yd��H^�ٳ�x���E,�~��v�٪�{�=�#���I���'#ɗ�wb�smC\�{ˋ#��7{�sݽ~xhg2��9;����-�Y�J����m��o%�'8����Ӌ����vy?j�>���jl�����Ņgu��3ʰ��ؖ�:r��X��ֳi�-�d��|���ϛ;�.�-�=����lÑ-Mw35��}����쫡}�9ӹ"���Rv�g�x��ݨ�}�s�O�O��N�o���+�G���p��o���},��cNf;1,(�w>�\�W�屮w��<2�Of���L�r{�܈��n�˙���={q�?��z��ld�{[kq��m]�(�9��, ���kr͹=&��O�>�s�Quv�W�����b� ��͹�?w3 ��˒U��~�Tk	RFە��K*�Y@��8J�!Id��ؠP%NF���ZyAH����&��bz�aid�V�qȿ;)�fs. ��ep�X�N�BJ��J7mvZ�|y�i�kˣ�7��Y!a������u��7���C/J^��a(Æ<Y�2"'��8p��,��Ј���2"':p���,��6""'DȈ�8YÇ,��,�6""'DM�8YӇ0�\.�p�8fg��ޮ���*��Ԣ���&+d�h�CTvՕ�ʣh�^��L#���-ڦm��LA�Cy�L����j�a"�Y��d��<{��8�nM��Ҟ����1�$:\�\���"Jpo{C����+�j��&7��T��6�6��u��yA���4qj׶y��6�.q�G�I�S~Xϋ�-M���"�Z`���0�K�(�m��d���!.8$�<ϟ��t,7FÕڪl,����;#3�|�?yL�p�g	Z����E#�fn���uX�����3z�M��E�2B�!?	�#kY����amv���]3� � �Ĵ�ď��-���ͮ5vm�mq�[�0�]�H�$cM�?���푣�H�9��-��$�c�����@��0�.oÇF��3�AT�&r`;VM������T7��Z^���i�硟Y��p�}�0�w��g.�=^���j)QU�$:"""" �0��,?K�o�b��k�#��j#�߶`�-mu�'8li+T�EY��gZ_4��4�(���j�!��ƽ'����|��HFI�wgȊE럑��F���2F�iV�E1gH�������L~�W����.ʺ�UC�����Y����=dCCD��䚡u��E>��h�6�~���Z;�%�ߌɲ�)�TJ��MDᥣZ��6����w�n��\ȋ�o�����Cx�8������`و��� �s'M���p�3���q:���u����^�V��Df��Dy��]hͣú�Z��0�v5�a~O����]�uX����d�p5�F{��&I���37U���$rYq�S-���76jr8���+c�)�ы3[W+�ӟcuf,�_�MS&
���F�MD�2�1@�V!��BRK��s�޳_&���٬��F�Σ�;E��ҧ:�Fֈ[� ���gl��ȯ>��|�����A
|E��b.��8�s��o���a�hs�!Nfy'����,+"��[����	<�q:Q��K���Di����`-��7�j�[� A/H�|8�3誔F���}��U�9����.ʺ�UC�іgzu��y����~��I>������G��(n?#��So�B�m�t)�?yeNh`�M�
G�����ͯ�m�af�B̅%,�`T4MB4�g�3�/l���.��ZC�>�U$���W�b/K�壁�#�Q��|��a}���|g��}�x�3���Y�ї�1ޢoZ�f�Š���!Ba�]M����ŵ�o����$X��z�?��f��8�n���s�
D�����Q����q�jjI-���dN[k#MD�e�9�'�˰�v�y��О2al�8�Lh�Nc׻}��5:��X9[��E�V�W����κ)�R�+I������p�l�����]�UX�����u��""""����կ��|������K��g��uy��U����d��du�ڭ֢���^C/�J:���cL��)Օ]�Б�L:t�'Z|}I������>I�ǲ���	�k�GH���g�s��O<m�|匦Ψ�:N,k>�7S��?u>�ῒ�j�P�t=���G$Tl������1e���-��1�#�����U9��z@�}FL��A�D8�A0OU�,l�
5x'�nïil�+e8|ug�ic4c��&#u���B2�z0I�o�g�c�C_.!�=wl�[�mZ���S��=h��<��kG;�?���d4���O�(��4 ����Ul+v5�c-Tl(�ː4܌�����#H�=��5gm�o_I�9�ɝ�S�wK~�h�ݥ��UB�y�&�r�L�,�[9ݒ:$!B��#~8O��:��tu�ߞ���-FG����ڴb�6�f�ɱ��Ç=��wB�j&�U�HkrKF����MV����F����*)���Ņ�
̌�0�p�.��ks>���4��}��N��:��Ύ�"��E�V4bf�x���������ѡ���J�i+ݭ�ʺ��p�]��u���q6�M�5+�U��8X+�^�B�{���o��	ͦ�>2���L8p�]l����{voI�ˊ��w~�p�Wb�2-
)Tw���Ç8q�Ø�,v;������ro�_k�a�C���{�^w#���ϻֽ���!m�����s9���qq�L�e���}�k��N��WÊ�����6x�g�l�E�gDM�8YӇ,��,�6""'DM�8p��,��,�͈���B',���,��,�8""lDDЉÇ8p��9��|{���K���}���i�����!�=[� A�R0�~/#F�v��}\����GH��i.�g�{��D���� ��V�4Z:��ׇ/]&]˧wEB�h�K,�b�l4�#�$�H{�������|��Z�n監F�c+�#M�v�}��n�����d}F״��{���zYo�v>��VOwD���g2fOi�ODDDDD�9���q��tM*u���Σ;��t�������Ԩ+	]��t!p��N���J���:����,��4Do퀱R���oGv>9$֍3q��:ً��خ]yz�Ud��~:d�;�:�xΜ���>�����aL���c�e�a�V�N��t����{UP�������v�#TVZ��Q*B�;��#�982��Q�c6[�]��aktr �j�Z����Q �2Yd�[)���4t��\%d�(0Z��DDDD��$���+uv�u������S��;P7�h�-�{\�O��cP�R:m&�����zO�FLW���냮M���ݭ=��Z4��-�R�w�bΈϤޣ[wp���+������z)�5��(h|�-���ܪ��xl��E�%�~�:!HU/��qJ6���H�qz��r->�a��&���G�=Ҭ���{UP������ηm������""""���{�6��ϣ=UUɋx������8s�	��`�m;�ϛ���n�U�ݬ��:7��%�V����`�|Q|��^��F�?���iE]]Cy>m��BW`SZY��&�3�a�RMy��YA�>����C:�f��%1]g��[6k���P�~/��T=O;Jf��H�YjT��E�')��J'�""""�9�~7!�3���n͝}��<S�e�YO�wT��¦����a�y�cm��qX�v�J�R\������$i-���}�vTa�9$ph�%�6G�������p���6�'e�M��m����*�ܡ��Ѥt�A������X����.ǕU
��豗��u1�K2d�!BbѡGŨ���Xv�|�:�Ǜ�1�)��8�P��UKL�C���4b�=xE��ְ�W:b":��ǋj#7b�ae=�h��-Q¹Zm��C�h�8$Qj��k{T���7��m>z��|��Z'QB���}���w�f����\ؚ��ODq�[g�W�I���ԑ�<��B�Lt�-��KP���5���2l���&:�u4��WKҗwf��ɔY[6�WWvl�sZCl�2��Ä=c�vv4Ұٻ�֠����_��U���5�,�G��Dq�,��$��Q�ۡ���q��$Du����>�QU�5�9Dz#+c)b�oa6e��\������!l����k��1������E�q�����V�@m�Q/{�}ձ�M��ћ�']''�I���5�v��)O��k�P�����3�j�6n�a��DDDDA�����/xq]�⩏�%�/%e�����Q��+��X="����e=���y���h�5�@�|���8�Rӱo������*�#q�K�A��K��%��K�\[}����n��;d�3Ꮵ:<�g4ih��7��������a��z�Û�znH���!B� G��t�?�.�Cw��⟴���ꍱ�8F7KK��͸�A4mL5���6`[�7�����j��kG��$"��J���d²0��ޮЌ�=z>k�;E|6�凧�]�g7o��0��[�:p�Ylc"3�~Ŵtn��=�J쑘�=Μ�g���k�P���8��$�#:I,ę �ͻsB�I�M����2d�{���ąM�cq�]+[G]m�;&tl����YL�e|B 6�� ���OI�&nܞ^�����\���
��c��|��UG�\���d.��Au6�^�5������}K\���Da�]dU�c��k���������H�^Os+w�_�8X.�ش4e���q6�M�5*�U��l�vuz-
)�'���v�8�L��f$�L8p�E|t��ˣܳz�Q�z�B�ݥ�op�دGCB�W�8��\8p�Çɐr�v;߳͘��u�2#�^��}[n�X��3��sO�-�)�؁�"t�+�?��q�ͩ�����Jg��яMƉ�E9�����T��`���Z������˟�L��*T��ៜ!F�W!��S���QMQw�E��\���1���K�����D}�l"��c�Iۋ�ߪʞ���.��ŰQ�� m;[��"vJ�7�fs+e�!؎�{3��;�Gx4d�����4�LC-�Y��a�xcŕ)��B�[ۺ���b=Ɋ�q�����ͽ(u���{b��kx ��V�c�jÁ�9Ky{���(r�g5g�6}��j��y�嵶۪} �^I�&3�lh�Q��C�*�5=�K���1dQ����
D�vX���PZ�E�r+'�G��#����0mj�
7q���A�G��D�#`��%��,!���%vˍ�����˓V��m��)�H#��>��\IJ�c�zg�ܢ2,��2s!L��ˊ!��w������ϓ�yEՋ��W�bp���,��,������6'8Y��,��,����bp�Å�,��,��,����6'8Y��,����Û33��}�;n�y����"i�2���&���1��H˭�A�"i5f�\7jSPF�m�T0��S��"H�;��׍�a�	��M��WVJM��vHKىa�ODDDDG���Z��E�g�p����▼����ͪk�!�������F��7�u%H�ƥ�G|����"��r)�0)L��熛)�>ae�˪��F�P��J�Ǘ��#�w��.k�ʑ�d|}F/��w����Ļ�T+'��ܛ����^�!B�""ٌ�V��S.��r(Á���h�fG
�,{<4mmqN*T��yb9ݩ������?�����$fF�f0�,ȅ���)6���m���g�-�]��G���)$�����}���}�}�>.�۪�d�tY��ލ���(��""""8.>Css�&O��3J���_�!�Es��ԁ�:��Ll����~t�+N����܍�`����C78�Q�=�s|��f��Ү.�	�s_$��N�9$���:�x���}Ջ�Eo���㎝�#^-�˱��Y=��vfMjk/��A:""""8;�{3��8�n[��Uh��4x�-JS�ܝ �JJ6�-�h�vUb�dsɝt9I��6�m�i|��XWj��\�p�m�����g�Ӡ��E�j��h�YgV����.h)�]i�F��������o�D|Y�w���ߺ{=��Y�st{��o�����5D$����<�e,s��ј\M��d*�[�j�L�]�R�1�$��z�2�j5d*�H0Y�HwSCMm����[R�6�%��_��"""#��;��B�E	R�$Tۢ6��ߝ�h�Gq��<�+t�qoG�
GW6���`l�u�x!a�;���/�9!Jo��jѵ�u7���,<��ø��-=ɐ�/�a��S�4�{�l�81�>�gt�4}~��j���4I!�,�!B���޵|V5�7�muEQ_+�q��"E�D5�FѤ{Ck��(/��-/���k�ɡ������{��­Ħ�;�U���<{��6l1H�El)Rt���c�V|�*�ᶏ���+������{�r��v�d��*�:p�B�!5:��+�ҋK�MY��L*��,��p��i�C4�v�-�)!F9h�&j�s�@�$��G��[ȭPy�O�/�t�HFFBl�]��XPV��J��z�k��&c�����(|Cɺz}^-���گa�y�'�}תs�������J�Ϭ6�)�^����pi�#�Z��jL� ����D�<-w�%���cW]���Ct��"�|��qn��H�{I.GN:�;�վl���>G�~���}*��y�%��.
�[�y�ち����������;�u�j���?��QW~p�6����[�W�4 �NS p�[v�V�W9y6I��C��R3;&��ƚ�P��8G�Y����興������em�Tlof�b6�e��*YJ9M����j���h�\V�b��X�Vy��4��Et�	���:�s�:�ܑƸ�ˈk�:�H�-Ur��R7�.iy����x6�~2(:�n��Nl��r�6���Шjo���w��rDD@��v�gx}���ܮ���;����$8�đFE�ŀ�,��BI�������a���#�\�Z��C�Y�zZuf�K>rDې-Ůy�h<�j�S���+M_�|�d�m��wqs>]W��ta-��P�L������qw�]��F�`m$[B7���$pn"�4r�.�޼_�a��p�{�C��Ш��'���Wb���Ӆ��]��XP�u8�Mѽ&��]
��p�|//E�E=��q6��k��i��L�3+�����w��Y�f��*�b�C츻�]�˻�wC����sYp�Ç8W&GI��j���o�ٝ���݋ۻ${s���+�sN�l]����o��h���Y��N�ws�8���q���*ڼ�]�'5�v>Os�F��FL���|&ns����d:p��'K����8p���Ye�Ye�'DDЈ��Ç8Ye�Ye�Ye�B""'8p�e�Ye�Ye�'�L����8p�Å�Ye�����ه�]�;8��B�!DmaHҤ�ф:sַ��H��@\^�l�&��y^{N���	;M��έ�]��	$k2���Y
Ke��q��5	A���!\_#M\�,<������F��ӥ~cgwQ���0��r\ur�y�|� �ma�7�t���Ce��U
ϧj�3��no:��d�B�G�_R-�"#�h�����U,E�����!
���N@G{m�i5�#R<���Y�ͯ����G�ߑ�Z��ԊBR7��|��9��u3^�s�6�u
����-}��h����Ð��7�`�s�F��}���ܮ���{���B�G+C�N��rV���"l�M�-���e9,#dr���k�ܤd��ۏ*�%�kw&T�?�(������NCfmmuR׫xBIKM���]6o�}7�������Z4꥽3N5E����,Yh�3����G<m�s��֖�#��|�(�Q���ѤiXw�WF��=��qh�]'���猲l뎟�
[��9��9Ӳ&���N:牮����ǰ8�3L�}eW�hl����Y�w�ϯ߰�Z\�6����DDDDQ�Q�t�s�GT�&η��V_)<���S��ͮ��{��4�N_��bݫ��"DQ�:�儈����F橏J�q�o�#�M��������h�m4am��f�����1t�O���>���ڪ�gӹ5�zfBLI�nl�2Cd�2I����Cxi��ߤ$����=�����;r������>��vn[�OM_]����Uڴ��{�{�;�φ��mw�kj�1m-�1N�ë�+9N��*�]�X��/�f#HΞ
�~*����0��R9Fz+��d�����>��Oa��]�;8�ޛv��8B�!Dz�����`�q���yNs�[�Ck�
&��G��{����#���3v�r#�Gʗw3�3�>b<��<�}F�ӈ�!B�x���ï��$���7�uYZAHh���3����>�Ob���ދ����qg��	�s-�Q��EH��a�]�s������y�ر�7���E�3����%���:4&������7�V�Z�]�`���)6�Gnr���""""8_!Ӓ	��b��-,6�D���$x���#��x�5�	�8��W%e<ӣ�8�0M�4�RX֓��������;���m�,�s�OsI�(}q~���6��+������|�/X�iyWXI���9�`���e�}��ߏ�������w}��㬒�=8w�#��]M���t����G*�">Ⱦ:j�okh���M��clcE�myvϔϯL��s���QȜ��ˁ�(z�C]�-y[X�U�����9Ŷmx7�uY�iە
�:�et��w�������>�]|5��kd��k�ΐ�!B)0�)�r�"}���!�Ų��F��I$�80�<��o�b�s��]3|>ִǭ��Q9�v��+㾴����>8�ɸ��0v�8W�-����۪�K������8vl���������(��}��2C9�,����Ŵ)_�Qu��T��B�x!"7�2�ͮ�6܁���������R��ܢ�n���-*��ʂ%D4}}i�2{�^���u��jJ%O�,M�%���pL�D��2!!s��E
���[XSN��!�סk��G�˼eR4�iZ�!;����s�N��M���cM�5E���9�=Y�W��}CCCCCCCB�^Os>9b����л|*��M�NhޓQ®�V��p�Wc��(���N&�zM&k�oFc��jaÅr>��s�ߋ;�9/B��
�=˅������,�rr�k.8p�Ç
�th]�����b|w�Z<�E��Y�&e�V|����S=�ZkP���$��n���uA7u���v�O!���:BWz�r06)%��ݙ�j�BJ8�[X�Iqŕ�|�r���ٕ9�1߬���L����k�lt{�*�!����'��lb���}�QȞ;�;w��>��n�ǀ�ɾי���ۼ�[]y�<v��z}2���E�h5�v�.}����j&;����ܓ�s�.�h[h�d��e���Xf���_r���1M��=0v=���xy��ۀ�-m���w/�bŧ�w�[k�-���!]�,-C"4�Zf]�J��en��Dv(��&�b�UK���r������1�=n�ۂ�J�i�Fw01���IԢ�+At>�ϭU��РO�������QX�D5,Oc-X[�YJ)D E-(|�{�Mڶꍲ���|4�z~=>�O��"""'8p�e�Ye�Ye�'�L����8p�ÂYe�Ye�Ye�2"""p�Ç	e�Ye�Ye�%	DDN8p��,��;G��=~-�J�Ҫ���ۗ�� �u�&g15�*�TmJƭ��G	[Z��ڜpn9���UvYER���9>x�pٔ15"1]1f`�<��4�M4�GgG���k�RH�H���SOh�]e�έ�����*�~:���^M�ԋ���QZ�+˾���c���U�<9�94oI���d��1'&�������u��K/]�z��f���D�=R+ʙh�yqr�E����6ăx#Gxj�^�*�J�W�w��^�K��9��h���!1�_~��h�ژ�/����x��j#�}4� k��l�ka��J׃Gʷ�H�ߟ?�P;�q��+��:�\�U0຋��NůuF�(,��z�6��K㹾.��63I鷯���!���kŴ)VzUB����(� �4`z�UT��oi���_Y�-!���������L^�����#lw�d�]ݲl�ى�0�S��a}΢��]8�q�ϒE/��UH�4U��f��6mN��9k�t��t6��h�4ZN���"6T�����9��=�B�g�T+�:�Y�bI�t�B��&��i���a�q����Rm'}�y����KD���Ʉi���s�d�ɬ�6�9��$�'�$�}C6�]�:��q�jli�A�D[ZF�"]�kF6��=#�Qk,cgo�Z@�Q�"4��(��|s8{�=㿗�]�[�����Ҧܐ�H�<�db��+�i��C�]v'�c���FX��F�dM�>�+��+ɉ�L�2d�{��1�?�j[-�lƲ*�º���K�W訪(�`:Q�KU ���!&��E?nW1Lx���j�� j�i��SR.#T�N�k���ȍ�M�"��lf�5�\�K��;v����]�[orHBlcLh�-5�#Dj�7�3突8�29K$(�h컌>����g�)2�IO��^-�J�Ҫ��cY�	ä �1��Ʈ�,��w�ҭ��/V�)��|�ɪ���-���ӟ#i����/���~:6�cچ�}�3�ر��܂d�63�R�Sb� @�����n�G�5�r���M�k��+E�EF�CZ�m����54z׏>-�J�Ҫ��y&�M{:4h��1�h����k`=�4�Q����E�Bh����X}����;A'Ԙ,Bf4X�jthΚ����v�lւ����e��~t����y{K���4u.��Ӈ,㋎#\��wmx��*�J�W�v�����$<QI'I�1����ɤ�$ror1�b�齫8�``��H�r@h~�S*2R"3_p-�6Y<�~0�F9ޯ-�{wѤ��.5�qq"-e�����|J�6g�ױq=��Z(��`]���������V�\�W�n�|-
U��P�h���s[�ri�B��a�r��yr:��\Q�(�C�(`Z��I�n��n��ܕ)C芟���M�)I��� ǵ����!B>[{��r�7�5��=�w��2��,�<�.#+����c5��[W�_}�I���E��ꨡ�tX"���
���R2�92�ƶ�*���z�����>F�4Dwj�44g��K6i��)54��?���T�{@�&Ӈ'ρ��N�=ty�/���=*�^���P��L^q��Lb8�2E�t�%mf����B&�!��{�<uk)��:����U�����⥽�G��������ٲ�dnHHLF�h����ڛ��eDP,M��k�rd�7 �S�D��D�-�D��U�4��ԒBF�h�4SG)�OfӃ֝&��K�>A�m,8�\IvW���<-��F���U�Eت��Xmv+ëB�����'!�e��W��r�`��z;x{���m7��e3�ƣ�Á��+��ŝ�Vn^+л��CܸW"��Х]�g��9��/�Ç�Ѧ;���T�u޺�8������7G����AXU�����2M���������9ܾ����j�&=|:��O{���{=���"�_'�͝�z�,ޫ���6V�^��gTޜ/{v��}�oZ��Y�.RW	�*wL�Ϸ/G���v�����]s�����,�𹙤�y�w׹����{8���z,{�鏸�Wq=�k�<^��qms���.�{�[�|�x'���L�>qx;�o�K�Q�_���˯�OF>�nw��Ԃ���<�g�_?�.o7��~�y��uw�{���+��w��9�G8�O{�e��R<g{Qϯ�q�<@;�.oٞa�\�L��{籢w���Fww�j.a��,�E�YBA�8pK,��,��,�(H"""p�Ç�Ye�Ye�Ye	DDN8p���,��,��,D8p�ÇK<s�{�~-�J�����iw�:"m�zA��<;�=.�6�k��jUH缹G��ʰ9��8&����w�K(->r�9F��W���m]k�s�ړ�Z#�Ѡ>%���������׾��J'�l�=���Sy3�����Хv�T������ьcѽwE�zl�`��Ո��R+1������\U�6!�H��v��b%n4@m����������m!^����Q7;����h)]��9^Ѷ�fZ�)k��xo���9�{�n�z
���;�`��<t�m�O��Хv�ދ��gߏh��º�*��:��ch�(*�L���q�el%,�YITr8A7ەɅvDUb�L��;Ydj:�w���=Y�1T�v]�兆��a���ܥv��HB��p�8,�f�
R����������p����ϛ��n��QDp��p��0i����r�*"�����r�O��<�g��i<L����p4����WXZ�i�˅��Y��=G4iM6Ym�E,����/͏b!s�O��b��l���6wJ�V���gx}�����E�E����qE�U����!I�7�FAр�-�4DTM���mſq��qn�cZ��lk�գJ.�u���k�ς�Q҄j5�S>����#�$��B��"-b-E�e6��{�+�}���PQŉ�:Nc�Ê'
���.�|Х^+��tr�H9�͙��u��3lB�Q�\�� �5��D}��8�c��cF���Lc�A�Qf}Y���tW�<��|��̌'��b��k�]lc�\��BI�#uP-G��{�J��5\܄��nс�/�\-s��Gͭ������ޑ����c��6��6)���^�*�^����r��P'$���K��1�#oV���m)��Z��z��t���ܚ-��bX�$$�m44C�G�4��͝|fϱs��c�i�8�4��$�Oe�1b2�Z8�p��O/��������`���Ǳ�dΏZ����J�w��Ş�X�c�������+�E^L�L������UV�mE�X�Yil�4�*��6�n7b�,�`�9ɳY�v�H�%r\��uyB���07b�kn)0�-�&�UNdiN��^�.|�}]mi�^�lͣ6�D^���/E�#�.k-��S���tkK��s�����Qմ}j3Jǲ�т���#+�Mv��#A,��\���CE��}eW���}��=��o�'9�s{�55�:81�cT�Ny߅���A�#�/��ľ�ĸf��d���MP�w����k�a]F�>.�u��/U.��0��>�d�]�kwq�hCm!��:z��fѽ��>3��0��v�խ�1�l
���UB-��к�g�������C���{�8�ٝM��c�sAlV����aߥ7�
^9�h�:�F�Cu�ds=���2H[I�M��
wR���]jޚ���%�MU4�y̟;�4�Y�5��m ؟;�Ƒ;剣�E�D71��<i��{�Ĩ8�	����h����Ŵ>K�zL��c+�6`�o&&�[��z89""!3�?|Á��=ߎ�Um�Z��[-�r[`�y*ȊG9�Lၟy�GW��?��>�oF"��,΍������{_}t��N�_�+��g���䑌�-|�`V�-p?��A/���CYG�"1AY�mkk���_�?H�ҝO�?����I�Й2Ga�p��\2l-����YL0�.t!������<tr�ޤ��d�Y��ߛ�Mf��d��4�4���&M&1SY�L�i3Y��4�M+#FM%&��%&��f��i(4���M%���h�5%5�J%&��M%i)l�"���E1�&�����+1�"�J��4�1���(ьN��Z�A��Ĕ�2E"h��cDR+1�эMf,E	��ٓi��1�I��+4cBh1�1&��V�4+�k�Dh�DX(Vh�`�edb*#AAJ��
�F�Y`�h��+�4,YX#@X4�,L7�TM�Y`ɂ��e5c%fe�Dh)YA��%a�4�*A���HfSl�����P`�nJ�~��6Kf��A�0J�h�A���уA�����Ɋ,��`�P��h1��у	A�f�I�f�Z�2P`�ef(0h1
ʃB��CB�A�������RQ�[)4��k(Mb4FVF�����YD	8% �H2���#) �����))"�@$�P�)�����)
�H���JJ��
J@$�P)���)�$YI ��e$IHR%$�0tlɂ�A1�P�Tp��)"�B��) �J� JH�C��,�+)
JH���2���)�%
JJ��$��<�`RT��%!IHR���%%IIBR@��%!	IR��% 	�(`BRD��%%IHRS�����)JH��!) �J����)JB�@�L)��H%#S	
@JD��������JR�JR�
RI32I�c3��3SRY�M���%iMIfjeif32eL����Y�̙�2��3KeL�e���f��[f2��,�Se�f�3L��3L���f�32f�31��i�3f2��ile�3Le��1�e1�a�i��a�s��SC0�c,�SfKe�f1�d�1�e-�c,�Y��f-�e��1�c,�Ylef2�e��32�c,ɚd�2f�3Ke2�e��1�c,�Y����f32[)�4�f3Lff����33L�2K�LB��,1*cT��ff��ɔ̶i��fYe�2��3&S�,���f��fd�%�&I�I������1���c334�,�����f�,fY,f[��ݹd�f373�30��3$�32LÚff�fi��X�fL��̙L���2�3,�L�f��ffY2�����,�̙L����)�3&S̲e1f��ZL���+LԚ�k��4��SK4�4�Y���iZif��54�4�Lf�fi�i���Y�i�L�SK4�4�f�32Y�i���3,�TI	!� I�I	&fHfs��@�a�	�d	��&YMRfY��Ze�je�Y��f�e�52����2�1l�R�jYK�,��YK&i����L�R�i�c4�if��,�w[ni��L�R���S���4�,���+M,�f��fk1&�&��3I�I��lF�5��ɦb��f�&�-�L�V�JŮ������<dM��#�8p�p����a `�B��M�G��z^߻��?a�?_���I߰~�	ȟ�#a��7���|���O����#�rxth�`��#��ߴ08�|��9=�?���t^��<??FOy��q�}����*l=ɀ��w����`�����O���ï��9� ~ � ~���~�Q�d�1%���H���� ���}"�p�	&=�_�������}g��~��>�����"����0�~B�6&�r�G��'���`����(:d�'ԝ�?����p�Y� "�����u�~��y�J���>Y]��l�"��~Ãϴ�i��|0��7��8AvH�e�A0���A}�d 
DQ�LȨ:����.b8��P��ɥ0t�ݮ���p�|���1��$
 BfD� #��*4Ĩ�����~��������МO�{�Z$���} �W���x@�0{��C�g�x~����?7ΐ�*"�O�pɐ=���89��t�"��~'����������Ѡ|َ�����)�X|�A�D���K��pG����������pz�������(�)�C鐁�_����a᏿�>���������@�9
{�xE����E?h|���%~p���a?5��T�L���y�Ð�����2t\�`��� � m�8��)'��V_����2�S
0d��>aʎ�?' P��E("	���@�@�B�(v&��N�9���"q�����	��UL!�>޾U�~o���z}}#��"� ��6��!X>����C���E���������?8���HL����S�3�����p�~p����������2�������?/d}&�aEOcߥ���p�B���~�0���@�Q���?����>	�x|a=���	�����)CA�����;6d�B�?��`���P�K��OA���Ԥ������'	�ɰt9���Q�I|E�����TbO�>�>���@4{d~#�?g�㧤�����H�����rc����' ��r|`H �S�9(�''X?������å�v'���}\qr`��Þ�6�}��)��0�@���p�?���.�p�!�sX