BZh91AY&SYHg,s�ߔpy����߰����  `�� ��@      �v�P���    P   �     /��)b)� �ǂ��� }δ��}�5�5��}��u֐���>���﷯�ހ���=�g�C,б�8�{�����b���mx��+��Wc�uj}�
������w�v�[շ�*���O>C4���ۥ�|���z��R�K������q����ϻv�]�����M�o�إ�q�>̽�e��}���cZ ���ݟv��=��ھ/�}=I{���{��w#8�W+�V��Ȣ[�jﯳ����>�ݷ��.����;o�����=��ݷާ�{6�m.�����=�K�2�����}�o]}>�{�ӽ���{������7�W]�;{���z����4�s�;�t��y���c����Z�k�{��>V��t*����}�v��#�;��m�g;���x_}��־��w����>|��ｹ�>�u�� > ����ϣ��q�=�{|�.����6��N��o}y���׳|�{﫳�G���3{�Uo3y�Y����<����ﻪ��:����                D�  *���T�H�`0M� M a�����A�&# ��` 140i�R�OJ�    i�   �� J�j`0M� M a@
��S=�S��e2OѱL����*(C�Td � �# #�|�l�����Ȁ@��R}b�`��~�!>#�pEBR!� 슥|����2��X&J�����?��������E��$P**��(�|���JP�$���  䈽�،%�I ��S6�A5�C��������������7��F1�Z,V�N��W��%h��1���lF(��u:">�C���R�4�R'_�%���vW���D׵+�m�M���2�>�&�"s����ߥ�zW����~��u)�ʳC����R�4�R'_�"�U���Z����H���pM������7�W��H�})���ߥ����|�OS*�W���M��܂q����2�~Aj�nU����<5ʜԳ��$)	�a��שx`Cs�`�7�SrljlԖ56NM�#��E����>�p�� �T��(Y���oR��_�M��ҬX�v��DH7r���zZV��v��qΥ�G���S�u줳����ǝ�B6H�>���ܓ�Y�d�9"wQ���bY�5U֪�d�E�X��xOn#�[!����7!ߑ��Ozz�=��%_g�螆�'�����pNA;�#�]H-K�bA2��O�'��J���K/R̩ �Iz$�^Ĩ�Ҽ/L�R����XI/$��O�P��s�,����I�0�ϩ�;O�}�t�a,�|�����|VC���"�ț��=���O\��[:=j��;���pR�/�q��3���zK���xj��Da>���g���o��H!��:��&�H����E�O}~$�֓۞�ݓ�����[��I�	~�;���P퉴�#e׉��V´TH��I�l�K�����٫M��ħ����>9��A&ӛI���ԏ���&��３�t��8;�w��_%|�+1�|��ԉ����0?RG�|�O'�Iicw$��rN#���y!�I��2N�N�g6WY;�t�5������s�a�FO�M}�H�5�>��>փHm��<���C����[�V�H�+I��8?vȔ��%��7H����i�:�i��$�%��J<��RxM7#�$��őd�p���m�����͎�;�(�C�G�%��W�?X�����;'�ȑ��<>�(NX���O	�Fl�?i"'z��IG>tO��=����#�%:%�8�#!&�DN"	�$�6%i"%"#g
�Ĉ��O�J�'Ӆ�#�}Ή"Dѽ�%��]I�;Ԗt��'At��H�-'K���;'��$��f������4W�DN�#g
���H'��,��J��8P�i���H���%Ĝ4;���%'D��,� �X��H���������Ȋx��6m���v{b2�s��
D�$IX�gH�7F��A-�}BB}x��$6�ݤDlR�<'夳�:%��T���sQ%�"��v�tN�J���ΕC螡�vv�GS����K:͔�z�;��uQ&�����ƥ�����A���������"[!��>�����J�d����D}�t~g�5Sf�U�6sep��S������[���M�J���M�E�G���*#~*�FҒx~�|8V�PMDy�����������M�f���y�O��S��ε8k��z��=O����������#���rC_xHH������Ty�D��:tuꈏ��|�5�����5F��O�F�t�!�ڈ�<p�>�2�"kcUQd��>GUQ�*"2'GMO{>D]TN��D{u�#���<kz�B:���'Jd�Q�j"mjP��M�u>N�E���Գû��+�O���pvH���I,�Z��uQ}Q,ވ�(M���ϓ��T�ʈ���&�Ԣ�":�DE�J�QQݵ4A���R��Q�j"y�N֧ȏuQ}Q,�ԡ;֧7>N�uS\6#7Q�����R�2|��U�(F]DN��g�����l�4pԈ�#�TEj'�8&���'<�Ớ�n����� �Q�{>Gҋ�
g�=�߉�!�y(�ܣ�%�Q�Dy4&��n�7%����+�G�*�|H�Fz�?"]5,��=S�w�M�Ϡ����w6k�ϑ���^�/��d�p��s1�b�'7Q��F�Z�=�D<qM��TG�rK7�ڞ�D�O�F��jy��jt�'�R��7mM���8o�9%*��j|�s�ϩ��^�V��涉&%�ھ�=�{�:=\��=��ۗ�3�.�M�v�����|=��Eta�]�Z}Z2D}��{����{ʉd蜒��e���F�'���0{�{^��������y}���͈�z�ӹ�f�"בѮ1���}�E��u=�T�ڕ9R�WD�:�Գ�}J��f�O_J�s��5���Q��c'�z{���8��y��I>�>úH��#��<x^$Y%�}�SC��=��3RvMH���q�u<'���z5yGFa�ĝH�>���:���8M'�G���|����r��|�G����f�GXH����cE2lE�'���}����^~G<��ʚ9MNv&�'=&�P���$;'��bG���>�i���x�u�g	Z1�Z��Cy����f����Pt%w�tٲx�%u+bl�#g��ɪI\��;�tJ;e�5\4?'�]�Y®%��%�DO=����}6&�{��"A)��O���L������MНd���&�?#؉ŕ�G��pu�_tF�Q��5�W���;7U)�D}r�~�Jؚw)��"k�+W��}�p�Q���J�p�Q�xP`�������ꑟ���8�L_�ob�ȸsp�	�x�u�l�s��u��>�ieq��&E�e������2`e��ua&�5�G�!�����U�6s��tޔ��޳{��[#�w����Q՘�3c$�a�x%��@�:aX?��ɻ�2k�I��|��c�LE2�)�����5��6�\�_2�ڮ�����=�|tw����ط!l��̞���H�*��G��:M?��܇5�R.Bi^�w~��p�P�9���	a'(�M,Y%���#}�W���f�%)�1g��-�����c9!��9N?d���Ņ�������j71cǖ۝/nk˃V�q����e� �����~,��z�z�<��r��͢���aU �K.3-7cx�����s*�o#�A�6c̮����5�f�Z�9��̫k���0��2��8bw<7%[�Tb��?At��z�/��E�V۸��'�ǳ�N��*vn`��w����3
�*R.�\�b4�A$���o�ύ��Б޻?e;�z{��1;��
�m�$�xh�Wc!)q�<d�ެ]��(/��6i,�Ob�����x�)�����DV���&`G�[s�&�ȌG#-�gq,����ꃾq�)�嗥wJS�S������:���0��87�!X]�ۏCZ�xK=
���/"U#f�K�en�
�d$u���1��ɏ��ȍ��~#�!�(o��W���6t3�I[�ЏR�7	�M%��o�t�e����<m���0�S�f�f6�rM;!בT]*mtɂKT�0����W^��a���q�%�ܮ��T~5�K\�j���	x���.1�����,�%��k��޹6�}ۙ}���U��|��2�$a��H������p��j$���J%-����b��Y�Gb���ĩR�G�'
u	���p���K}�&�P"�W��w6�u$XN��Q�B$K�}3AHT���HT��/C\��-�|�B,X�l��t;.	�X�>�K��Xn�'`ٛ�C�7�i͔-�Ch_ed��˯sed��������$��Jfsh�vf�d�sNA{�6XN��ߞ����/�dl��:�� �v�t���5+&d���m<�)"�fS�ǃVJH��߽��S��#�"O�㹹�HoC��`���S� ���Ԟ�%�fz��i�+�/w��>xsr� Ĝ�ʉ�FJa|Ac����AgMD�F+R%��r�|a���cbY�����Xo�a�)�T-B�ۄ�����;��9���D6���UպB�Y�ۃIQ��#|���K��Ȅ��{ՔuC���lA=>����zyѫ�Y0� ��bE�Z�ѥ��G:��1\ñ�HW�����v����+�15��3n�5�Q��}}�nN�2�B��n�6nl:IEҊ��U��1DQ�(0����O��Of.R	���md�DMjٲv:�Lt�	W��a������M�a.�`VU��6Pt�v�(���PZ~5��u��	̝{N���w���_e�fn	�z�J��}�-2	��gҹC1��NҌ��c�Q
5���l�w2(�Py�����-����8�I�8��?|����+A���ɗs�X#Y��7ػ__uǙ8[9�f���&0�qZn��Ǐ �%o>q�.�m�S7�#���]ʘT��W�s]�`�?{ڙ?zNڳ�~z�p�m2�e%�:�̂�9�]�z0�u�p������\�1�><,�es�6aլ�Z'�5����l�i��a�r��ͻ׏���Le�׵��&Q�eC2;ξ���c ��}��4Mٽ�_{,h�{ /���be�o)^�ǧC%�WMn{�������`H��2�_Bx������p2i>�~����{��Ɍaa?G)9
0��]d<��IL݁\�%�M����o0�?�nll�Q`��4���w�����զ�⯇�I,ȓ�F'Z��M����FTv���,a7���yI7*֊�~�<�߻�,�
}�e���\8O�κ�_D�"�>-���~�k5{��3�k�	�Q�'LLC��X�?��c�/�]�����o���<�Ik����UD�����y?�ߏ��~Ȧ^��Wo��o˷�����aZ�+�&+"$��Ҳ���n�Ɗ̅��C�Q�?����r5�W�&W	g.�dr�Nf<1�D��E�#�V�qg�B��F�M;Lҿ-�mМ2���T�ڴ?��ga��Z�!�l�Ö�X��L��޻�0�!�u!��-���9׎2[f�k#�v��7���7A���nZA��bÚ�W?��L�s{�K���5+���>(�~5=Zt~����X.manػ�3�	�t�)�UI����xh�3O���~ߞ>�'�3���t�D��z���=�ہ�4R����چ͇68ᅬ�q�
W�,)w�w�^�9\�Fe�r�i4�gϙ�����.����G��,��<)?�T.n�Aqا�/K8Um�&0Ǯ=�Uu��:n��&����<�ٴ)�
+�;�mW~+f5YÕ��'��=��{��r.�z!�zau�I�#}���w���:�]۔�Nɳa��bQ���95�>�%��bڮex�sZ�6�
��9{����=?F�%c�<(ݭ�l�d��2�Y��p��\�}�g_p������;pb�lV�u�p�N\Xf�+x�#�[y�̚Jt��Q��{ܹ�1�w;k�I��]0��$�5�3.&�H��>y���ek���N�i�E��ep��߯��aM�������-�i��h������ݍ�_�퇚Vc����w[l��=��̧q�Y�w3��o~��kN5�R#�;N�?�����%T?\�������������ǉ�c�?��}]�p`�?��$�?��N����	����"g������p�Q���J�]mb�h�rh���͟��	l��]-�66�	H�c���N"����X턛+d�05�h���zz\�y�2����53j���Z+��!{1e���IJXU�DS��K)(�ͳBƢ�4Vl���j��w���\1�������Y\Ak�er8)�Ի^Ͱ�ŎҖ.�5x���kca����m���L�KbŮv�����g��'�  iEZ-e��&.�=�4��K���u��l�Suׇ�<�Y�	ۂ(6�"JM�T�i{;.�ƅf��4""�m,g��K-�x���޽��N0L$�Z�ZF���)<�5�j���kl��e��@�]R1��`�m�j�۪��"�l~���z�6N�y6���y)����3I$l�ry̓d\݊5�[֔���TR��4�]o5٤qHƛ&�A,��B�}���_�T�\Ĥ5�]&k#e�����-Ղ���)�tͶ⩭��%AI�9ՙ����j���z�^��\�؁��I��J�Z�M����͞�n.t�2ᗈ�2@, O�Tu��/K�b)@�p�8)�B�P�$,2D,%�9��V#H��uդ��|�$�CmX �z��'���m�&kQ���!�� Ť<Á�N) L0dk",�2BV!-F`AzN��[��p'�nx�BX�2��6A@��e�2����$�o�����3�,��ȓ	����K8Q
FX�o!��A�g�>�b���������jHd2&�a�Kc�bDD󾛸t�	�U�$�����D�i7�<����KE=�������,c��e�s��9P�A���	�%�hA[A�Ʉn�I�d"�ěE��`��f�	0�H`K��kPG8��k
���`�R�;�O'��u%���ƕ�ּ�]v�tm�ְٳ_aÖkZ����0OI=i�2w�) *&膜�KCYl�n���e�)fl#��%����|��Fnt���>�'�Ϥ�]�+��q���3�Ш����nIR�!�>̧����?��?��C���$@��D����>Ϸ[�9�r��s�渴���UUQUUQUU�*��ťU��U^��U��t��X��jҪ�UҪ�ZUW�Ҫ�V�Un
��]�J��W��X���,���9�FU$��	�QD$@�7	��[j$�E�!V�"���Z+"�DcH�9�s�W���]��v��U괪��*���U[EUUEUVت�k�J��]��Uz��Uڪ�Wj��^*�Ux��U⴪��*�[c�UW��ZUU��*�UZ��|�Ё���
Aq�BR�b��[bZX(D��"���+h#@@���Ҫ���UU�Ҫ���W��Uv��Uګ�]*�Ut��X��h�����UҪ�*�UW�J��ZUU�Ҫ���U�UҪ�W��X���/Wn�z�"��Uk﨟||��i�K,��-R��*$��-��l�.k������sQUUQUUQUU�*��iU^��Uz��W��Uv��WJ�Պ������UUQUUQQUTUUTUUm���^"��WJ�U^���Wh��U_4|} }�>�
�Q0�\�L� 
f"J�a	�(�	%��B��V�kH F �+"�"�"�TX�yQ�F���!���m�$�5oE$Aa-���� ��9�B���.�g��~ߨ~�EP��F������~o� ��}?#�|�}A��i�}�N8p�Å��'�	�e	DЂ �	��F�M���'D:&�	�6%�,K��""Y�p�"P��8""'D�P��<"tЉb"xN	�6&�h��DD���bt�D�8"%��X��F���blК�pD�O�C`�hA""lO��<&�&�Y�N�D�ÆN9�
"cv/p������M^�����iJU؎fm���Ļy���%m5��d5�5�|:��!��Ւ�j浍!I[��Ȣ0�cBϥ0,��pC�m�~�������`�hͦ��n�-{l���j��-���e4��t5��e�m��F2�KmHq��SR�	s.~�������n4��R�2���n���5��4s��vμ�z����8%�K66���΍9��{�=<�������4bJm^<��7��#�,��5q1��IqbG����3qڻE���  �qҺ�����J�M(�.EZ��WJ�JO���찻n%��v�XSR�p�.�a#{Bb���@!�!���b�inf�P,ZۭѺ�[vc�"�m���6�bCpgjXY�T�M5�Кj�|��ϖ��V�e�"3|�M�,��&�5���qw���{x|��	�OcMt��5U�}��+��_ܯ޾�y�����||}���{��f*����g�|�{��f*����`|�{��a����s��<�$�9$�m6�l��n���ı<%���wӓw���I6O�U�,*e����ee�g�uҳ���e��բ�X��=�کٌ�f��[�����6�2�t�#�4�-��vd%x��U`�%�Te������'����?g�8{���C�*_���2]���l�6h��
>
>e���S-�V�j>m�_[K�s>:�I$.y��Äè�\��X��6�ҥ�#��"��sM��9�G�cN�잽|~|�m2�-�ۯ�L,K�XYW��W�w�I$67}���^�L�K�JL`0fvj�R֢�M�m����	�ӗxj�2�����S�4�̧<z��+sݕ��㬓ln���I!�	���h\}Kb��=x�2m���=���\c����	���/YB	�S�ON�N��bX�����
�������oVkx��w��<;�X3��G���3��a���Vw����fN6��^ok���m4dY�wIM��L>�n&�/���-���N�}�A��k�Q��T=��'џ|c=�_F��ͻ�ϞEg�������Zܭ�m�z�-2�N���\q�q�=�.����#���M��p4��	��9�_<�d��n�>j�K����Ht|l<=�)8%9��xw�N��>{�n�>�>���ǋ=WX�Y��W#L�Q������걙뽎�M;7m�V'V_2���,â"X�'���{��A7_V�k�Y|��X+�Wm#��M&E�����.jH��J�X��]�����-��;XhU[EaEK�0(&��5׋*]��"�ת7*e(��d��`�K��ո`���pLYD������9�4{UW!v�:)d5�l5�K&���m1��D�4��|7:�����7A=l�a0�.�D�Ȟ2�K��m�f���aЈ��an�J)�E�I	��$�e�Ļ�6�|jM2��'�u㞽���֚��ߟT��dG7;K���2-����Uǣ�ܘu��s^�!2a�p����b"tDK����>�IG�����>;(���GC�Ő�`�@��E�7����,.{��;/¢Tj:4e5�M77�Co5$!�����}fLI�	:;�z�cR�>u�X��9I�5�Y�u-��2C���g���2I"=`��J�VnO��N���ʵ�#�m杆��xѣ��6xK:"%�bxO��rId�6o�����0�F��e�Ï�uX��Q�N,oei5����)���Ϗ���Jr䵳�.�ZU ْm>������8aI�g�5;!;�x'H��)�ß0P�S��bXE0$}-%��8ZB6T��R5�(�V��a�&�F�H����5�ّm����s��*�;�����.p�ܧ��Ja��ı:"%�bxK�����I"�NT�B��M98å&��S�	��|�UF�2�����j���a�p��N�$:�v�˾,O3K��ߎ�p�.w�����!��
y~�Ig�ò�a3��U��t�\\�=u�x�+1溽���M6h�,舖%��,�^����M�ԥ:Z1��/�4�1IґzvH,�wie�u$����5� 6.c��E�`<h���j�Jط@�YC}�l�y���1$���6�UK�����ݡD�lLv���嵗c��7|�>����WU���dㄽ(���k<�d�T�_n�e���
�Lf[5�-�xj8�������UTD��\���E�۔Z�db���Wވ9��O���2I!u��+)�)�OM=<�"X�'���$�rI$,��\:��p�蹡o���8B���ߙ�e犌Ǳ�r۸���ի�3'������=�#N�f�HL�8�0O2>��uo�Y���YwM���2B�g�sã�	�3��	��v?nsz���G�t�d�}�WC��x9�W�B	��UN���Ea�0��V̩0�&	FRtºC�ԘA>�'>��B|(�|(��_,�X^���u�:ê�z�:���_����&׫��[^��^��(�$�(�$�	�a8�]�μg���c��?1�����^?1���0���1�e�:�^���}c�_��~u����~`�����/�].m�+�z�^f�q�:��+	��+�D��L0�V	�`�}I���y��^���r.������������`�vO�,X#��1
'���|DO�>!3�:���z�Xu\V�a�ir�-��/�~c�����:�.�g�����G⾼���lyV!#�3��1͜9$BZ���#S�g���@��>�YY��g�9{Ϧ|Ϗ���9�������*�۟}��{��fL����p�W{π���ffL�s3333{Ͼ��ffL�W;λ�����I���J�/�|��u�L0K��aj}L��������$�}��
!�t�2�`#����~(�T`�퉓� ��R�NWs�q�
U>��~��H�@Y�?GҎ��"5t�_�b�k���"�Fa=3tW�3s���bFc̮]��J��,�Z2��o�n�)�����Sښݘ��~�V������!$C�cU�a=�L�eOVC�9�t�4���V�`�-���̓R�����������3+�6^2�̼i�f,�a�,�g�:Y��	!Q����$2�&v=Y2�G �	�CȰ�Mwή{p�Z�롲)�'6�I+ќ����>�i�i���L@R4x�K�6A�h�K*���T�ɸ���ÑMG�~�F�⟙O,�x��*�Wһ^v�����a������^�Oi�p�IM��X�7n���O%���<YVVIȩtğ�W���柚q�^����r\�����Wڝ�|n���%�7�c��_z�i��N+G��d$fVJ$T�Ȏ)ɑ�I�JŔk�[i�]h�dM���aU��k-�]R6��M㴚�bM�mw�I$� �NRP:��x���5�=�=������a+v�r�<��SK���=�2��E��U~i�:Y0�gXM��[/���b��OX*,T�d�RUI)z�A��#(�7���#����>�T�<�'�j,a�,a׋�UqK�}�f.�x���dy"��6a�h��ǿ��f.щ���##�#X$`�A�e���z0���+0�O#�F3��{�׸�1�=1�G�vB��Ɲxz~:a�X�'�����3P�j������U:�,ʿE|��1!�5[��mQ⟢��"�{��Q���6�G����q9�f�+�I���1p�*�C+��j݅�svEab�h�����"n)�db�������vêO�S����F��LpO��^���'����ǘ5+oj��W���<�f�l�m<ۻE�B��)��ci�0�Z):�Hl�X��rM���a�a��U��[��GXFc��Ɯ�,<f{�V�q^EG��X���q�x�->i���_��`�"'�������k�*������
O���s��Qʟ��~�(�F�~�1�K�<Rrj1&U_����]��pN�7�I�D�h�A�a)�%�f��d�(��NX[6\�*B�z2�\��K!�4��Œ����^�5��c��x��gX��z�Tz�jjf��Frh�e'�u!��o�..=�O}�i�Ua����db+���V�r+���Fڊ��0�����$F"v*m�}�i��i������:��:�n8��9e��I��I$H a"y��g��˶�{�I�l��`i!�	�'�%+�@@��ؼ�g��^HUa8��płi��_MbO�U⊧�a���b{�i�s%TU��$!�(��YF���z�{)�v�۳ܯ�[pԮ)�['�y���T�S�#�^�L,W��SjU�����a�S�X}�u|�"���6<�C��I��:L���j,}S/�aǭ4�M�����X��ß��}_Mg7S�M놎k��C�fo)�:�^�h��)��TR�N(F����<`�n+%R��Ab�7�������"�1F|y��um}4�GA�%�J��r@d.%sˢ`��	�I$�� �� ����S8ps)��EuXQ��Jv��^��0�r`�B����e��)�dҋ)����V,�Yǉ�5�˶�Ǒ_�a4���+vM��;m��1%P���m\I5S�%X��C�&��_y���Ӆ,q�X������IVB�m��:\<��Q��"��~�<���<E��UQ觧���l�g����:a�"'������\�I$�D�g�>���$����3��89{� ��ib�.o���t����E��d�:�?gh�F���=i�Z��落6\�Ӆ^�&�΋�h.&4^AA�}���ԯ	�\�[�6�N�mc.������s4�X�Kvh�lRq�$���$ã�͐i�,�/���[ѣf�l�Y��X���z�ƥ��+��I$H#�_����>�rXт�7��V�2\� �n��n���@��	��a9���d{Z����!��	?(�*!F�IKMu��˽��L�p�'��o�QD4������ ��E5n�6���ɿ����=���'��3�Ӆ-�jbT��^�K�0��&��ɩ��e��6�N?=~u�ێ8���<�\~��I$�0�~�c%�M��{f��F�Y2���ڡ�lO�%��2�n$�zv��M,�sX��axr0;7xL."&S�<�Ri��&R͋��Zp��z���a��u�Cw|��kQwfWd2bd���s?
*������CDԁ�II�G�+D�I8V�!`�k��4���ufKD{7��Ǹ~N�i.�6]"]��}=O�,pե�C
?�??����a0jL"L&	S�Xz��K����ge�����*��WV�V��x��ut���ӬN����������z��Qd��(�
0�FF	_aa�D�D°�aI,�[0�L&�F�a:L&	�L**��0�L!�
�d�J�C�0��	:a<�;_�p�?��?������aG�_�����	��$�$åQ0&VF�åa�a�L�
/$�����4�������u���O�'��fՂ?�_�8(���p�^�]\+��ί�ں�}����Q4h�&�W;'c�c�>>�ǅ������0�AO7�.�,޴=S{,����o]�p6�F=g��8�|��Q�M�zRhX�qHdQ����n}s&�ۃ>K���Cʴ�l4�I ED#!D�}h�2R�D�A�[�3V�6cՇuS��/������8����a��v�i�&Ih��~�x�U
��$,D�Sx"���؜����l��2���u.���N1-�k)�Q�l[Q�3y}�M�9+����Ж�ԓ �J)|�0b<
	^A�8�}��B<m�c�!qgT�)cDA�ڂm�Yd ��	R(B17�Y)�d�,���A�!��S��ً�zo��˯�h6ց	���gk_}��!�����U��4��>�׮m�2E�/̰�6VI��8ƌ>m�"�&���1�&�d����3bk���E�am��WiwZ��G�Ow��oϛm�@�a��|�&X�v�b����=6��V��"m�V�jX2YV[,�(�I��ݼ���U�3�(�r$�ep�M�����Mo����u��Ǌ����tT4Q$&��up��A�-e6�π$o�!�������ʭ��������ffeb��c���s��ffeb��b����s332�U��\���Q�:l�gL:a��0��OON�OQ;�ݜiz�K7��֖&��#�@j�s���XL��B�;i~_5��7T�-��|Y���L%44J�!jq(�Q�baeM �D$Hڨ邨J*��̻1�K��^�gykh�|Vʼ��裸I"A6s��Lm�f��F�Vf�;��do�9�rDْ�S��6�I!��9<�a��Yy�c
aO�w���j��ּ�F]�3WEoc�9�b�.�����=	F���i��y�у�6���y��1�=�Ɲ$`�秓K�2_�:בU~NV���V7EL��������j}��<�U?G��5ϳ�x���X�:h����ǌ0��D��\I'�~�I$�9�a�}˙��)���tٲs�g&5$���$m-��}�a��{�3���m�ن9��߱�d�����3�}�{9ڝ?��9�H��N��te�m��*�Q�GdJNt4p�=����{=i|8�b6oڵkO�#&T�̮g�0i�u���w�z�Jۓ��e��΋^+�-����u�ϝt��<%��W���Y������(�f|>�9�4�X���C�޲*���ٷs�qM0�7m��m����M�����">=3���P�|�o,����2�qB��7�AJma�&?z�as�B~?*n���7)M9��4�����ۋa���l�<!��fA�f�{���|\p�C�d3�Ӆ2�ME���<�s��}>���#��7f�����i��~6l������af����}%W�3}�I$�L ~��a������s�%u��ME��'��O�;����țk�9z�Y!���@�s<�C�3җ���6Q���xo;8hx!ŝ�ڵ�m���Z�f��rvg��B�6|R;A�vQ}�d�f��i^��d�z5�j���-R�c�����Y�bR4�����-{�6�i��?<u���&�Å���Z��4kz�E��"R�&y��m�H2'5���<u�l� ��@�Y��9:(���fG��^�$;L���~w|W�u��]��G!D�2�1�b�k��b��G��Ж����s,��Ͷ�m�O-���u;6�:�$4��|/��~�2A��Z3����*C/^.lHĤ�`0Y�0���wR�5�IשG��n$K'�L�+īH�L�8�8�]�X,l�i��&eT'�`�fv!Ώ2����s!�#�>��@�90y����qIK�A��?;|z��pz�r1=ɷ�17ə���ǭM��
���6�oz����]p������"�!=���$�I&A'�ד��r2�M��ھ�1�y9��Pl٢KfL�%�f69R�����j=��*H0������eᖃ6,����r�$z7r� t!���؆��{q?�y�+���i��w���s���M��DP�up�i6D�-�^��`���W�$�h�eh��-�%��J��l��Q� twd������u�ﳼ�:�Ù�r0���J�m�]x���κ뎏��������_e��ܹRI$�F���$e���L�K��б��Im�&���PQ�r�b�g���ӆB��hfV�&�X�֛�[c�ē\m�A��Bl'���8p����h��.��nu�f���f#�a׋z���(�r{�~�F�
`�D�I5��ƽ6i��H\Щ\�዆(L�}��. B�S�ƚ���������Nႇɪk�䐴��IA�H�]���J���nI1҈l�cF��4d��Ǐ�&a�,=�͒V�Z�a���ꤒI���8%7=0��R�O��[���s�`5I`�Z�v�3�⪎�}�%D,0c����C-+!G@�]��V2KO��9�g����7�׭�a���x��S��'���핖~�=T=ý���&y���0��q�u�ΡU���tf��W���Uq&�F3~��ѭ.�]�0)`�D�m6EÖ������ce���)�a�9�<���Y�{�#�U�L��O�=~z���_��y�ou�G�r�Y�*�`���M*�A)T\���EL>	ʄ4�-�&�sn(�2���ʩ��(�$�DX�zp�%��\�nw���۱v�6�kqm0�#)yn��蛦�4���=)~���I&�c�m���2ZE��UM���s-�K=M4=�����:���f��v�I��p��Rd�c|l�K!TS��IU9`Bɗ��	n��&L�x�tѬʭkyM00p�GS;q��p��8���y���u(W4u8�ͼ��[�j��mޕDi�3��S��G	���4�kjԻ��>�3,�<�E�ZV�2Ӎ6���ϝu�u�ζ]��f.l����F�$�I0��g��P)�����;x�����ܛ�8uv������w��,��X�vHY<���O(����N�e��SEz���p���ek-<�W����/ۄ�ngG���[Ym����\�ƪ<ϖ4ׅ������e�ʯ���G/翝MG������yE4����!cJ3�-��g�h�N�5D�!��'�?�'L+	�S"�?Ǥ>�ft|N������|	�
'��Ń��4J$���]i��Xug��k��U��~�x�B�(�D�I�Q��0J�$0�D°�ȘP�V0MYf	��хa0�XL!��$�z�u����Luz�/W���]L�&�:a_a;&�(�0�'	��B��2��0�0��~'���u<a��~c��r�^�u��W��|���tU~'�J��������G�>,~!�n#��x���WV���K���gVu|~!���G��?�?�h��I����.m빽c�����������2��zT9ڢБP�r�Z)=]���n�NAw1/�/��TU�\Dqy%�Lf�Z��Nu����:p������C�<߮��A�nr�3f��Ҡb9�\A�tEE׭mf�	�cY�
�{�'���gq���UW�s��9���*�劼��9����J�Պ�Ü�333*�U�y�(�N�:p���p����ǧ���gǁ�v�V�!nߤ�I))!��C��w�1%J�t�F��0�D�h4b���k�-��eѳe�Wgp.r��ޖ��.?8�p4J�'���Ka%%��MV��>��B<�s�gyC�<>΋�~z�m~74�t݄a(2�4Ѷヸ�5��:[�I	4a��2�lN�4��(@��Ufh�q�re�=�s0�L���2��OϞ�?<a�	�x��+{����ܪ���0��<��[-���4���as�	��ۏ�;�9�/�d�ܗ��T���}��IL��H2b���f;v38�u�<m�]��i���[�b�w�1��g��I���7�S�&��Y?e:�!G=�#R�B��Pp�u;t�{4x�Q�,������6�s;)��G����=��|�Zmǯ��_?:�0�X^��=	U���ʕ�]��byHM6*��0��b,��\�Yq�[N`���JUZ��4�n�s2f��6uf�
J��ޓ��ę�k����"L�St���H0`�˓9
&����$�I�-5��mf-�Q!���Q*�����y3O���{��N,�p�̧N8tS��D�S��ĳo2�N�C��'S����̛i�3>r���;m�f~S4�N���f�X�c͊��J�'�8zd(%�6i)�!�K#����,������9f�ldmeU̧!ԏL4s�d!`��0h��������)qU�L�x��o_��:뭺뮶��ySu&n*{`�jj��ɜbG�3�H{L\Ȅ�9�s\�1CU��f G2�D+�f�D�P�#��#�oS�s3y 8�� gĲ��@I�s�UUUT�]�lt�i���=ü�:�_+d�X�y��|\Ц[�i�<�Me�m���t�=6�`�iRؖV���R����d��,�֦�i܄I%�P�#.\j�e�mde��B$Z��XLl�#1m��2��\e��I��Wr�KiH�5��lql��XYl��$�,�b�,�.Y���.F�	b.[#V��XV*���cJ�QfHF��FZVґ���r�Ȯ:HM�eI�D�-c�ۓY"L����.߭e�@ O�NɎs��(�Y�v��l�d��k۳��g�L/��íg�	��?%�j^�]�����tַ*C�+VN�<��&������ck>q��3�fN�a�㋗iԣ&�ʪ,,�:;$9��ӭV�Yi�O�z����]m�]u�OA��-��$�I�<&�D���9|�Z֔����a_��<�G��+İ���.N���W�1��d�#�ف��8'�';�<��f�QV2�&4�	�����j�H
C��2�g�!��OBœ5UU1�L(ty�҉��&�a�L?"�4{�=`�^ϝs������K��i�J
!�0���)��ؘ�$:���RQ�.S!�ƍ!��	��0���x�,�0����8*����$�I��{�d�Yb������]�$
-c���E��~����Ѡ��`�[�r�k�qɴ�K�$ae̇g�L!��{�C��Ì<bHBI�iw��(tt�N�ḟc��c�ѥTh�_0RF`Q]��܌8C<�w-**�AO�i�b�(C��is��|���D�x{�.�Bd7�N,��p�G�|��^F�q�����ckW��D�,���t�~<a�a�Y�^��ݓe4�tYj�QLhݥ��E�%�Y�����X�S��z�*(��g�4R"#�p�ĕ�w��rfˢوMq-w)&�6�l� �E)4M�����&�m�FϞ�t��Nd�[e�,��fp���p���C�C�Jf'�|C�Rs|��dS������6^ԒPCga$�]J=�w�ʩL),5=ۥ��u�b�J�	܂<�^I�H���;.bv3�?F�r;qM=���+�~�TٺSx	e�ͮ�\��	��TQ�?a��p�Z��||L=��I�!�h����0��������c��~�-d�6��I$�a>�y��53���)�{��Y$���̒H�=.<�N4��R�s6R�5%�J�����������j`�ԷR96�(�E���}$�IQ�T(ӺI��K��y孟x2�;�p�
ɛ�����֩��� ]���G��7	����Z>��.�M����=nv`M��CE;v��m��y��x�<q�m�/�u����0�0�,�	ڢT���>�I$�B��p��ꞟa3/�J�%4@��)�Y0���e2]6a(�Un�<-�97f,nY<m�ͱO�h6=e�).\;��Y�f��gܼѶ��7�A8/��H$0soȊ�{�������~DU�9v�sr���Z�5j9���@Ʉ�}���L)�9������ΌN�_����e��H���a�ώsO^�f����s��+�̿2�����|�0��0��P��ꪪ���4��j5���%ܖtS��p�X�����n��^sk�(j.s���ɗCG'ީ�$���C�ɚ�p|0�ZM�csRI1��0������!��p�I{���:"y�D#�78���t�ܒ�X�GZ>q��_��MԲ��Bx�G�L+�°�L<f�0��eI�Q��&�}�h�ҺWe�uj�WV��b��YWm�ۦ_k��U��g^�꺿/U�u������u��"C�U��"aZ"aX%`�����VXJ�aҰ�aXK#�����i�����}^�U��I��0��L+�'d�Q�NK֘�^�Xu��N����z�i�"L8UVT��0��++=%a2E�����؞�W�X�����&]&��G�#�~)O�+�tQ�'�D�(�?��?�:?�?/����W�����̪Ҵ�-��)>�����_�~���u�ʗ/��b���Kqn8p�Up�FA�ܶ�iq��� �]D�1�y�:/�����Y�B���Sc�mr�����26�˝ٹI�dl�t��I�t�sFy��+p��\me��U�^6T��'j�[���٤᤻Z��8��%� �]YY�v�5�qx[4�hV��m�����Y)�c����
����K2쒺�����G�Z�����d��� �j2�����{ڜm	����7�,0���c���LCT�Clq��d��,��c0�w"]xOWGL%�L��te�Q�34T�IF��:1��$p㪰�)4C��m�N"�^�}�|��f�ϐ+XY��GK>�j�(eB�k��Y�5��:���a"�i�\Gl�X��B*�kK��5���f�l�D\{]iRS���uΗg�B47dt	y^s����4!�0^�[���Ե�)ʳE@8�\�l��?6}���ń��ѕ�7Q��~��>�ivp��o&Ѝ�a�a����F���h�ӋDfG��Fo�<�$�,��^�&�<�e�j��m�х��ע���=������!o�8���4�*#X-y����n_~����9��J��i^gg9����Ҫ�ZW��s�����U괯9��33336��ZW�8Q�4t��0�0��0��5��w[�V겊ݨS�_W�7މ�6��9�AD�vSQ���Ig#k�f
��]�O����Vʥ�5�E���	����٩$�K�	��1Ye��,��"�Kd���B�zY(4e�	,� \�F\������~�k�e�{�����J&�����.���f`������Nw��͌��RI$�n�).Qı��4S�L+�ը�t�F�,�J,F�{v��s>�k5.���SLU����	b�H�a&�3�,��3T�q��g1�5kW#��+�zˎ���:��]q�u�؋�$�I&����Nb}��~�4�����H%��束�CèCRgXx|Ss�����ٷ:3�ψN��?�|����A�i�n1�$��2�6s	���N��e�	s�R0I�,M�͑2���=Y�GX��[m]'���o�^=111:��X��(�����rJ*UTnuֵ	"\b=�X�i��̽e��޿:��&	�YI���(��UUQUAC����E7<�i��}���B���9޼��Y�*�ü���a��t��
<;�������E���ε��	wc
�j]a�a�Üx��OU��&�{���p�}���v)I4�K�i+�sI��u�Ľ�=�n�����T��x/�搒�οLL:�<��'۶�fM�0��%i� j��5V�ԭX��(�4Y��8`�x�ae��kE�^�d�I$s�P�u�d8Aܸm�b�1�s�)�L``�o��X�Hɑ+��e�M���#��B��L��y���`d�_E���zb��=&.!�?8|~��0�>��w��/Y��F��0�.p/����L��&�$�4Qw8i�Υ��0��.�%�&�0�����[|���:�:��[��՘�rNݜˊ���(H�!ߣ�)I�����wy,<�c�D�vLd�8����2D�}A�UE*�!lVHФ�5aE�e�Z��y;�+�K��mҌ���k,N��h�4�6�Tw���I6�i��/ˍ@���]t(��Qk�t�vɄ���1;�ꚪp��A�0�G�te2�i�r2CQg���']�$�h}��5����߸���S�<��ф���s����#�D��:78\-��<�}� a|.<���0:�j8BE�J�!hHRh��$^���1����4���E��	N짧�	��&0��=�U^��5UUUUAF2��f��KB�{��#��r凸��QK�vq��*�ڒOKZ֭-ݔu*�G�a!����e���G�֙F�#1���*�(��L��zآ�_�-(�M ���y��V��k����U�t����㇍��dx�;�����,�an��a��4b��C�������u�񷱸�,+׬���N��a�a��YH�++Z�s_I$�H�9�(��#��.��P�&p�������kss�r&A�:?P�>���������G��=s7�0�js���1f����Ԯ�$��*2挧�l89�Ȟ`t�P��6�ʓu&�X�le�4cz5�#�v���F��\
�n�g�������Z��wr�i��h���Y�z0��LC/=��~u=ݶ�u���+���~m�Yu���믝u�u��m��$�H�	����ݛn��p�%<\�q�p�n�Hh� d���0�.7�g�������l��hɤf�[�d?d̹�.w�Ba����`8j��$J
�Qp�-�.�*NE2�!�XV]}3#�_�a��'�?+Y�I�:��+,}'X;�Z��P��묢��=V�Fgywqqu���M��ss���^�V�2�0��i�-��=u�κ뎺�n��:�=n��H�c���y�9�OUn%s���O�}&Ҋ��#l3��1Qɍ$R��i�S[,�0��e]�hX�u3��$�*��/�ٶ�m��ϝ�`7a�l�ۤ��ZtT�8L��O��0V�����%o��ڵ��S,�\�z��i�a��=�������B0���a߹3K��L��9�;j9w*�\����a.�tj��QY�s2|�"����cQ�\�e6��L�Y�7;_F]S�Xu*R[�j$�E΋�s�J8��&^4� d�XrI���t��g,��2�/m�.2��箺��L�,�U��Iv�UUUUT��:�8�/�I(�ɖ��G�h��na�Y�9'�ri�\�x������^��%QR�7�3� bz���c���X��6�<�(�A�&J�Vz�ge��r���$����L��:/��k*It��w�T�+��]4�,��"��rIW!�}�W��3)�9�U�z�0���&g��q�8��[=m[u��D�btDK:p��4P� �!bB	
dM��6"pD��xKİKı,K�K�,����:�Ƅ ��b'D��Y,���4&�١4ADM��OD�"lDN��%��8&��8m&͉�(J'�H@D�!�bhD��:%xCf0�,�6a�~'?{;�k9I����9������F��7����)-l>�(�RnO�N������́�;��6��D׾���=,���_ñe�\�ͪ�V��7��ffff�^+J��s3333j�t��7������*�WK��g�x�Əa��a�	�ǧg���{ҏ7�$�Ie� "h� \���҆�$aI�/Cb﬚�J0���\ɂ���zY%҆Y�/OK?ig3�H#�pō��Y���<c�yFm�m4*��Q�N�ü�(�\�q���������/"H�l��Lpʧ�o+cr�k��[%�m�FG�f���\Y#��8Lα�	��>�a�)0=��!�!�]3��<bm�L?>e�_:��^��Ŗe�N�UU*�񪪪�@�2aM:"�%�4���3;;��!��������y���l���*��,�ƺh秘�7&���y�p���CJ4��7�W#��Ʊ=~�'�|_�G��W��>vrfX�a�L�2�a���γ�$>�.|M���;C�Y]�׍0��_2��_��뮸��უ�G�rI�7&[�DA��m@�"IS�j���a��#1�I�/�T�6�iE!���nlF�f%�U�:���c����]vv�\j<��c�L�%-� M�Z��I C�=�ʖYMa�r#io/j��L����'��0�8������C�,�.x�t�$��RDpS�Ou8�!`(�d!AO�IAؓ4Oi0���~®R͠�;GS��RY��N&����P��|/������h��֟W��Ƈn3�Zz罼�P������ޟL<�`�c��3��1��㍽a����ft�tL0�0�:Ye����$�@��:�����/�p4A4�}����#&S��i�^�6F�d��U.Y4��n�*��}�g��m�isO��I܁���������ivѷ��M1ax��6�y������a;/>���è`�>���m���f�X�H׌�M�=c���'^%�c&K5/{/7��s+U��!r�|�%�����>���m����/��&dÝ���|���:�\��d�̤8C��Bh��0L0N�Y��!'�6J��I$�@���i�9D��c�ڶ��fa�b��u�ٙ��3�g��i��[c2]ڵ��;���$	� C�I�4���Fp�a(��#;ϒ:du[YA�e�C�Z[/FI���A]�b�9���a�z�-hڰ�;53�_ї�Oa�	���9·�Q7gxu��t\ˇ>lTY?�}�)�.e=ܧ�	I2
6�8MN��Hd�G�f�х������M��M�s��$�I�����j�g<{3���3�^��<�'�oZ�C��&��}az>2�́���<���:�Va �9�.��~�0��I	c)�"�m Q��ؑ����[ h��z]��(���F0�0��K�����8�.�E>j1�����~W�=i��_:������B�ha%V�[���<:q�fj�:�/�mb�0A��l��a*1 c`��.@�$F�2�.OΗ��ahcYi���vls����2�m��I�ԛ���wo@c��6����+d*2�D��v$�I$��2f����]%�a�6���Cd�#$�G��>�ϻ:Z{��!��'��<i/�j�T��!
$7�Ӈ�z�n0�Y����V.�~������?6z�/z��������a�܌ǧ�F����>�����O&g�F��B ~�L`�D��2_x��k��]Y���:>=?q>ɐ�����<N�ښV��q�^���G�4Y�������`�`�,��S�$�Iy�8u��y�#%e�i\��0�pܡ����O|����!����_wr�ɛ$&!�[��0x߮ͼ��U����e������9�>��=
�J�:�!C�6���:T��n�l������gx{8��Q��>�V���&Z�j:t�y�gY�iO�9�ޥ�������n4�<���a�_2�/��z����e���y�f�ڪ����
>�a��D�+b3Ji���F@f��[R&'Ftw3�O	��o���K�3�P���ݷ[DG#�F�nU/U`��)�g[����Ml�y��ԘNy�y�r�»Fd�&-h��ڍ�W��۶�Ϳ4����j�j]$���G�~O��^a�vp�襚?���舘&&�,�׵5�k���n��I$�\���~��C��6͆�����a�!��L&n�	���d���-l�f��̳V�U�y�CFeܾ�2/Ĳh�X�O�$�z�1)��1p�1 No�m_#���ߴ�+�ݼ�#ƙ2�S��\3n�T������i����S���ZK'�(0z�f�,b>�I��|��[:�\~~i�\zD�,K+���4P� � ��P%	�6&�N	gD��Y�<"X�'��b%�g��H%�""xD�H"hD؞,Ј�pDؚblК ��6""xD�6A���'DK�pN	�L������(J'd�>D��"wdM��8'D��	�Fl������o��o\�6>L|��Ӄ�$�a����wn�8�@d�Щ�x����^Ha%)yv����st����{���H� �f*�`�*���B�,L��yb7	�e��`p�A@�i�ֆ���Z�Vi�4|M�(ۓ����^�R<#ƌ�IBHʈ���ؓ�"p栆IK��H����!g�"��WP�����v��d��m�J��Q!�B���(�߂�1��f�,�m)��G�ެ��Y�q|l�I�҅�jD�1cv��Jv���$��$�c�T��G�d©u����i��r�P�Y(40�5T�Hc.7$�$�ӗ�"0@��Ӧ�6�u?1ש��%zI�����w�^�d����\Ap�����<Rk̦f�w)�d�m��E�-��Ƭ�6g�°����ځX%�W`�MIu-�l�۴ۑI�۶s�^9Iǅ"TjV?f|x���!�Rjc��1��F��k{�ޅ�5��bQ[��8H16�����1a���}�Q`N�ʍ�3⬢I��\��T97�k�!EUk�j��v�����]��y�o9�����Uڮ���󙙙���]��y�o9�����Uڮ��:QGN�:h��:"&	�	���������\�`�1+���m#��y�}eL]ˬ��R�@���Q�&��MN���йfI�r�=^�̱���{$�I B��YV�ZK%��֍��)b�駁��a�'�7L�a�A�	O.Fl�])�Ը`�;�P��di/�-��B���5���vг��x��N�O@���#$$9�7�`��&:?{'w�M�`��́v�qT�a�x~~>�R6�f�[_`��:YF͚?,��>��A���GԒI$�C<��8(���!�I<��$&�m,2�a��j����p�E���&盆���I����-Ui��0�p���������达T�-f�[��m��5�%^�$�J.ze���NSd!��'��9a������xp��'��E�x�4x�'L�%�a�hh�/�;�9�I$�H\�P��e&��r�#U�I���l��=ۣlMF\���M���Umk�{��^�p���R~�컥?:���Z�r��n[U�Y��;�|u��ʜ��K7�_>����TUJ*���{��aO�fS���;r��Q�UZ�4�喾�}n;&�<cno�|>xLO�~�={1V�x�����_���f`�<Y�����j�������E�'�H\2dvY4m)��Il��K',��Y, �ZQ�����w�G��C�7��4s�aA�?��f�ќ�������b�p0�2�;�I�wip�LM�UU��'�����N;MvE�c���---�Ɠ���n�r��rth�G0���0O�&'�V��EY�gE��!���l&�p��"M+T��(�n�ۯ��fJ�$�/�q!xY��;�㱳r�v`�B�e�Bd2+0�S@�ف�[�m4�[�e3-��:K�Ad7#	���I$�I �q�X�x�'v61�]�9�sqN���msif6h�8t���=�BX�=|i.��1���|.ZI!���/l�Vni�-9+��SNj��ֿs	��LX:d4x�}$��)�`��|�ޘ�m�m��ݫ��ˊ�~�,�ǉd�Y��-�h���,d�ft�<"X�`�4X����2I���[�}I$�H�i��u�p�$,袂�xY6��i��wNa2�Z�0�p�}B�����p�>�0^�g��y�>�g䟩q'����E65B�YS�l�+&G�7�C�����X�z���#G� lǵD�S.
�	p��K�3	שgSŌ�V>����x�ox���^�O�&'�{7_T��7������(��t�q.�N&�ˆ�%qO\���4��9a�wM-�abC�h��_>�z���G4b�Z���l%�e��IP��+�
�2�{�r�g}�\�=(�����1���HF%�-����$���C���:�9W=k�2��D\��w��K'r8��,s�ʛ��ļ[e����Ϟ�vCG7��1���F���ky��ɉ\���.%ob�-�ֲ�zٌ�dT�^m4l�d�[l��D�m����w��M[b9��m�5��6il5d��H���E�Eo����'˵�q������\ݴ�a͝n�4�K&M`�V�mҲ-��P$ZV�1��umz���q�'�Mv�:]񄳃-�)Ԏ�,
��C�PL`�|�c����>q��~u�̶�a7Dr������ɘk&��&�+���$��*H^H�kU��9����Lx�W ��%&n�5̎a��u*¦s��5��39��8a�*��s \$�*�E�G3:J�3���I$�&dþ�d��L�Ke�%X�[%����+3��$�#�-d���F��X�4豂Y5�B��e9OK7M"���57�j�e�ڳ����:��i)�|�L.2I$�
5{7N������nFFS�Fjr�JJ���p�E�4Y��'�K��}�$�MY �ݹ�Dw��r{��x�P�Rdb*lT�$�N���˛l5����C�)K�ݒ���7��k�}�Fķ2�S� �&l3�/V� u��Ϟ�O��|�$�I$ns�Y u%.��n;)v;Vh���>f��xs�>x{2�޳��{�pzz�|�S���oK���H���<Ri��&��;C,Ǳ�=M<���2דٓ�B�(�e4l�ً6r]�`�F���F��m�X���e��g��rh���3�լwqɶ��ӌ����a��%���<h�w�I0�}��߶�:�I$�@����'�n)���/"Iw�%p�CAcFu4x2�4s]��Tj�Od.m4����V��2.�׬���$!=(�U*�:E�`2d�\O���o�g`�g}�.��W��X���T�G�Y�����S�ޅa�_=�zs9�����)�=�8jm����l>6���N�믘`�a�%�(��4P� � ��P�dЛ8'N�ӥ�I�<%�b"X�%�bX��%��J!b&�DО6hA(M��$,N��6&�6hMD�"lDDnD�B�舜6"tD�,N��6&�2i���l��$�>A<A6h���BxK4xM�0р�GκӮ��9���U����E���7a-�j��$����E��'�'y�����,;d�j�KD�/r�9*;�&�9��H���3�#��oW����b��<�o*9G,����RbϪKy͸h�� )�ٕ�\0#���KA5 �j ^+x���oX��fk�[��FO��U����x��s33��U��s������Ϋ�Wo9�o33333:��]��9������|����(���GM:"xD�0�<h�|�I$�.aѧ|5M�,mdFÙ��\�űc�h�`�]0s�ìN�����8�\-?e�c�Y��%����[e^E�b�xuzÆᠻm�6�3�IکR��0�r���#6C�Xw�zy��*�W��LNG|{�������ryLM;�F����lчJԉ�<~:"xD�?'�;l���VS�{ܪ����z}�}��E=�ܠ�0�P�t�[�������P�^MY^$�����Qk7u���N<�����a��f4�4����Z�h�}J{7��HG[!���p0�盅|b���&�d9V���+2p����2t����`�4Y��:kp�ʟs������j��V�b�B?�hV�0��PR�WB�ʐ���n��-��~�=��n�Wifv\3c04D#�Yk�Dɵ�Ƙ��	��l��U����m��O?\8��mN�!Q(TL��B�*�ɖ��rDI-�;ϰ��?|����Q|�<�řuV���U����{���I�K�n�;=%SZ!�FC�R�$������'#�'�8�g^�����d���S���<�Y�xt�g�p=��~}�cu��21�M�)�i�\��J�KJ���s�|�'��zN�:�1������	���,L0O,�ҧf�W�)�^�$�Hgg����<H���_
�>�F9��M�cT��*����������ϰ�p�2��Z\t�����F�Piy��Y�y%�MT�.�#X}�����^��Gy�2p2e3Û���E�g�͊�#V�8r]�;�F���y�Yu�R�,��w;K�[\�d�LgRHB�>�Rt�x�Z�t<��Y=�n4t�I_��n~�u�<�l�e����8��&'�g�Ž�*�����g��?���Yi{��Km�!�a��N�T�w���<og��N|��C�c�k���%��L�ꍫGb�B�xT�F���Ns��G,�l׊ِʇ���$�[4��"x+eITU�;�i<蹢��Ox���n*���+�����4��_2V���'��<"X��Ƌ7���>jY�{$�I D�cS��4��~<����k��1H�M�v�W=�ޕ���9�)ˇ0��u����䝎Gc���Yu�fi����F�S����sn0�~����m/�
8A�9
��i��i4t��'�4Y��~:"xD�0�<h��RC)�h�H�P�Z̤�'�$`Hd�H0]�$W%4*Q��.���?����xH��.I��^CA�.J��c�91WFǩ$�Ii�ZJȭ��K����N��s�9�L�?i�g$i<�B�ӧ�;P�
<�s�O���}�ɀ,e2i�Y���J�ʄ0�N�:0�&B��.a�}}�(�<�� �?]�i���+͕R�yj�3m$l��þϾ~�jr9|��L���_����%���<h���5������������pֱ虁'�J87�i�\�QU_��p���[�;}b�ߚc9�!��:{dH���M>�����`~�Zϙ˻4�͗]�!��d/������C��i�o�UYlh+�
r��o����3���̚,p�������b~0O,�ꪪ������N����Ē2���flut�΃�>�X�*T��%8,>2��w�Kn�?[��qe����MiH�Юڢ�S^5$<b��,�=y0k)���P���N��N�w���)����s�zs�����w�^2N���"#�0���a���žllXB$>.d���6Y���<"X��Ƌ3=UUUT^������
ti:�8ɐ�{��i5�#ð���X�?Y�}Ws���r1#	%�U$\'��=���I$'�%=K�M��&�Bt�o��'2��fƤ��Na���7��~I=8�=���'��H�m���	�E}��}V�uȬ���L6x���DDO	b~0�0�8QF ��BhЉ�8lO	�4x�<'��,�ı,O	b"%��4P��<Q�Ј�,O���lK8'4P�$䈈�'JD�"lA�%�btN	�6hM2P�%��4�jO�C�$��f�D�BxK4xЛ0�,��0Æ&�BI;8T��$��	i�D�_֗�e�c/M�B��ɯX�J1��Nq��n@���#�
1��!���*m1ܪV�($QՈ�ah!0�E�����db3]��JZz��[;��K'��F�m'p�� �!H��o��FVI�J����B#�nC{-T�G�ԢY�S)hГlGS��uQ!ցS_$7����ʊH��4%G�)��U2-��IC���Pf{�J��.6}�$�j��I�T�v<���A�L�v�TG����Nb�D��e�:��c��v�zІjNibG �n'һ4�h���m��!
�%��e)�%a.����4Q(Yi�{��P�~{��9<��Ɔ��U���dn6TYl��E��+��!
���#�I
�(��ˁa��H%�V���B���a\�&�f;g]$�b��Zn�4.�ƥ����x�7�x0_ܠa�M�f��tiy��An3q��0�P@�חP�5� 4�!5xo�-�޷��y�$%�/}�pD���<��{��6k�t�8�=uA�C8�4�Lq���u��~��}�ٞZUv���������ҫ���6�ffffg��]��9�33333<����4x��G��0æ	���������ia�]n"�d�L?8%�c���m������,��[l$�r�-(��Y&:�v2 ��KIu�h�X�\�͍�	=�e�Φ����.��ݒI$�4��!�%��5��#�T!��g��i{	ĸV��{�Ӄ���d�ytm�Ju��a�42����?g�p�<=�Qn��b|k�	$a�?a���}�/fvx��=Z�b$	����gf������y/X�����X���5Z�nq����_�m�~z�<"X��x����+��|J�w���H�%#��L�����Ǹeцn�9����1F�aS���R^�$[I��i2�+ڒHB��mL��w�	��Y�wc%�RSe\e�݀�2�g�𠆔�)��R�4�u��,���J|h�g�0��O�"Y��+MT�S�I a0�����#���^\�ɨ�֞G����}+q�-F$�]���;1=7�Ŧ�n�<�_F�~h�ܽ���K�ྦ)�7؅g�Z�[�z�S�':�QI��/�UW�L�
5Úg���<�!'^<�$]�M;�ƌh�Ii�;(�xoF�Ə<agDO�"Y��Y��ݯ�b�q$�@�쾎g	iiI�M�(i�G�<>8xp��fʶM��t�'&��kk���e\:�1�mOg�s˼�?n���m�~�W"���J:�ɲ��n��Jl�.�&S�-�$�1`��QP*S����8)o�ѮL�ٳrmc���Oe�0�񣦌6'�:`�,D��7p>�1�ɂ������l�k1.��u�9�)5��3j�Lvc�J
(�	��S�$RƉ5Խ�$�뫥�;l�t�iI�v��K�t�S��_���J���ε�-����\<&�k㱩سe�Zm��M�����Q\LnPov�<`�R�A����+�R�h4�5�	!$ �sv�p�xw�;Y%Z����3������Ʀ���Ur�oYq��z�gL�%��a����k�4s�I$C�)��id�U(�{ōN�ĥ�z��j[og�?S�OK{s֥��q8�8�b�`�����By3��z���i���C�K脄(5�'�$��(��h�����s==��� ��vf���GͶ�ݙ�tN�\���?�7+
m�e��Z|�ۢ'�K,��,��M·$�H�%�QcI��BHGm̆�I���������0ŵq];6�����X�x|�����F�*�%&ER��������V�X�b�ę�SU�{���!�>���'J���m���痚�4�H�=�7KbjTd�e��H��@��L��<�p��\��u?U���>���x]95��0����rV_�:㌼e��O�O�xD��ǈ_ލUMԭ}(ꪨw�(���\�ӛ��@�M�P6,Yu�H�+s�I�K�n�R���&��;�ڪ2]�$#��4�<&���W5�$b�0`�Y����\3���.�gR�����J��X��t~=7�Y#�f������B�G�f	���O�"Y��7��s��q�J�N�)1F٘�&ȣ��eF[,*Wi]��&�Yzc�Sb�FG`��Mmq ��4�0��:[5��/���C\�d�/�a\T����0����.���U���!:�Kn;Kt��GUPH���wG���>�	�~r&���Z�ɘ�O����vۇ轞��a��=�߫��1<�j���jq_��a}z�C�����8ϧ�2���j�03�M�X vЌ����?f��S��}��xs���4p��gOtD��b%�x��5RI$'�'���cph2�H�"Mi������|��t`<�g�wF��$<�0it[��R���܆3$�?
8�z��Q~[[�������p҅:�N-֮3uUQ��!��8�Q~��I<a4�&�&rgG}8��p�Q*	���6ϟ4��Bt�â%`�<"X�bx��tæ ��4i�6&��:��<%�bX�%�bX�""Y�<p��%"lDDK�M	B&�D���D�blDẓDD�"'DK�"5"#���X�'N�blКIBhJ8Y����8	��DGR'���p�Bh<x�a�0O�֣F�G�E�k�e�ˋ�nA��.;�v�Q��Ǿ�O5躼�<�z�'KN�Ȱϛ�����+�܃����p�r�y����m���s���ffffe�Uy�s�\����̶*�9�s��������U�!Ҏ�:h鳢'DO�㍺�[}�YͶ�N>}5N[IUQ�WAvM��8K>���bꪮ���SMTN�\:���Y�Y�k�?C_z;u�$���{��^�ܧ��ηl���UD��!Ø�Y.[OO[sW)伃��'�Փ��)I���uI�!t��c�ב�_����Zq���>q��zx|v'����	���{��u�).��~������<?aI�%�I;ee���wĖA5d�$v��RJ��ü�.}���?~|�+��n���z�<zlr�0^�[`�i0=ֽRI%���(�T�ɽ㐐�X�m�<���y�[���u�[eƝq��xD��ǈ_ޟM�2pw�*�`�V�X֢�7uݤ`�QsQ��!�c{{�3=)}=��7�����kYɅc�s��V�D.�¬E4���RZ@�bWv��VԺ(k�akN�UA�m�X��`��]n��\nѺ��C�za3��C�=.ok��L/�7ECTQ��8\$��}ϛ����ƌ�ē5�Ӵ�Ĳl������:�ƶت%SET�0@߮Gg�>7;	�;U�:�%FA��ʌ�"mm�p����{$�m�<t;*I*����~,��E�<"tD���m����m�m��rrx�Q�������V-�"�#j0�m��;ھqQ��gl�y���q�:��ʑ�έ��]��7i�͆�(��Aћ*��q����]ER�2j�{g��)Hi������&�>��!��Kʪ��a�n2�|_6�[f�6��Xi����a���LY������;�,���s-�"�G��S���<�2�l�ˍ?>m��,D��ܪ��HI$�7�$�C�ĥ���X�8�˂��Td�EY�Mh�u�׮�xɢ��F�v��Q�v���6ĖL\Q�KS��4������k$$�p�u���3m8�g�a嚚���t����޻}��gOg.�/ӱ�a�GM	��t�'�K,�x��h,<&uUS��ϥK�zp�RHC>)����;�w<â����HĒt�6m�I�ڲ2�@�i��͙9�%��ɓ��L�|�8��d�D=*0���;d��	!�Q)�'��Q'xp�v�Oڞʹz�:h���U%`�%�16C&,a��N����by����V�Ns�1I��@R
���LL5��hC0>T}���䏰mI�	:Mw�K�k"�PGV�ho	)��omo�ݡ4�h�^�kK��i*MlZVͺBM"}�:����-��i�[�;��)���0��N��0��	bp�.W��󔽌�4t��Xi#��ģ�\d����N�m�I���da|�<ѣ�r�"�׳Kk�����-m��ASn=vm���f�>X��Ɨ��X8a�Ə<X�?��,O	�,�sf�/X�I$2��t�e>)���!�ã���s�'T\Ɲ�Ú�11�U�m6a8�K_r���)�,L����w��G~u�մ�i$����QJ^��4�"9�r�ԙ�h��°&'_,���\��wo�q���S��<g�:h��	����<"X����Ͻ���m�r�5UȘ�����S���֚�h�X��6��)4�{���O̚Ð��b#f��*�ȸ�W���N�}}<<�t��j��4�Hi.]����3�o���eǝr~�γ<y�L�vvv�VZ�x�WcJ��Ϙe�^2�N�Y����:�N^�N�I$�|��٨�*ծ��%g�1��~ߎ���>{�菢������α�dٛX��CӇc������;=�˴��:�n`��HB�ۓ������e�Tc�ITm3ITP�S�酾b���m�s�s�/��̹pѼ��0�M��7���Jzu"S�������ؒ$"I�I	D�I�*�4Q����S��)��I��,#����X�0a�$H�	$`��|�����S�,��b�""� )O��!��UR�UU%�UU,V��T�*�J�J�TQJ���UU%�U*��URX�UR�U*��*�KT�KUT�J�TX�UR�U*��U*�R��E�T��&T�UUK�UK��X���X���*��*�)T��J���J����J���X��TX�UU�X���J���X���X�����UE�UU,UUR�5�$ʕV*�T�B�YJ�,�R�U,U���R�b��X�R�UER�)K*�ʪ��)*,�QU*U,Y1C�Rʔ��R�e*�����������UK)*���,��YJ��e%T���e*���IeJT�P�R�,T�I�K)J�X�JQR��RUK)JX�*�T�,T�R�R���J�ʒYD�*�ʖRZRʕL*O+2�T��jU,�*�T��RUK)J򘊒����b��,T�K%*X�T,�T����T�R���U&���T,��YJ���),T�URʕB�R�*����,�U*P�,�U%�*�*J�eU1I���(��Qe(���)1(�ETQb��,QQE��)�L"�%��0,QeQE�*(�S�a���Vl[jԖb0)(�E�J*(��(�E�j�	E�T��QeQR�(���Qb�(�ET�ϥJ(�i1QE�(�Ȣ�,�*(�QE1I�E�EY(��QE�E����&"�(��(��(�EEJ(��J*(���(���(��QL)0�,�Ȣ���Y(��J,�))�&%�JQJ)d��J�QJ�Y�)E*)E*)E,�Y)E2�LD���V[iIQK"�R��R��%,�R����R�K$��(R��%*)dRY)EJQK,)P�%*),Rȥ�TR��E*�R�K�%*�)d)B�
Y�����IB�%,JT��Rĥ%))bR�RY
X��R�,��
Y
Y������)b)RRȥE,��K,)(R�JJTR�XR�XR���JYK)b���E))B�Fpf��&�a�JY)QJ����E(�E%�(��K���*)E*)`���E*)d�IJ�TR�)IJJK%(����J)aJ��K)(��)IJJP��TRĥ����K
TRĥE))IJ)))d)IJ����)R�RȤ�R����H�"�%*�)B�)(R�J�R��IK�
X�P��R�J�(R�R�J�,�J�,�c6LJJE*�R�K$R��R��R��ĥ�,�)B�%,��R�IRR���E*)d�E,�)RRT)RR��IJJYK)d�IJ)*JY)B��%,��)QK
QIB�)RR
Y���*)QIaK���R�YK)e,���JJX�E*)d�E,R���X���R�,R�)b���Id��TR��)b�R��)F�f�b�JQJ��R�X��J),R�,���R��R�,R�J���JYJ�����K%*RYK"�R�(��YK"�)e%E,��K)e(���,����K)E*)E,���)e(��K%,�QJ)b�R�QK)(���R�(��TR�QJ),���R���K��)b��K�J)e,���R�,����1�J���LPĢ����(R��E�IeE�*���)�U,��K(*Q,�,�������*�J��*���*��(U*�E�UB�*�K)b�ER�EQb�R�,R�T�,R��QT�(�*��iTUK)T*��"����B��YEQb�5R0�Qb��Qb�QTYJ��X�QTX�QT,QT�QT�*�T��IU,R�UYQR��U�b�IT��J�b��T�J�TX�R��*�I�)$�.��a�H|9�2��h�)��|�}l @H�BIPP#Xz5�$��f���������Rs��� �/��mXh>�����}a_����!��Ao�`�������}R��_�ڙ7�L?��U�����;�?*���?�dp?	A��\��{�|�U@�����ٿ��{�Aآ'��Q��@�A�����G����?��O�C��A��bP�ŗ��?�7�0�C�?����>���
'�TU�}H������0�P}&�,?fh���E�g��@h ��%��rl������К?��)�k��tm���I��`C�?_�d0���Z�����������tP��!���\�A�G��1BD��	�	�	�R4��*1�5E������܈4Z��Aj�M����.XJ����O�|���D* *�iU#�1BE�BQLRLS`��ZU$�!E%��S���}�P0z&Co���?z���h?4:��r�``}��P�?O��?1y���QU�����,'��2?�ɯ�o�@������?��A�xO����
؁����c�L������q��D?�>�_�� ����`��Y��'�ƨ��C�Ag�}����������@�?!��P`C����?�X�R�W�	�r��$����i`0�O~��|�
���{lm�X ёց�)QL8F�D���$��|��PB�2?����3x�
(.4��'��HP}a�Zʆ���O�F�nXL�CzG �`I���U@i���^�>��~s�@�n��U@ ��0��� ?:|ߏ�C�S{ }a������׾�F�|��K$�C�S���p�T���?X}���A�R
�ܖJ>��_�?�?W���EEP��]~�R�@4���ƨ��~��7�������6 �a�O������K�	���,�@Ic��>��x0`X�pK���킏�@-�!t�}�C��N� X8\����L�|%���۝��
��9�O���%䤍D���~@���� \<�X~c�'��۴��� Q����`x=?��"�G���)A��b����Pl����ϑ�}A�j �|��%փ�t��.C��f���G����S�$�?BPP��z|k�����w$S�	��r�