BZh91AY&SY1�b�S_�pq���"� ����bJ�|          {�񘒴�M3cR���2)�Y5��BV�M�l��5���(�h���JZ�%UB��F��T$Y�Զ�}���u�ַ�v��� j�MR�5k(��MY��Z�f��E�FfX�jJ�ذ[%URff��U�)V�e���-4�Sf�����ۼY��� �r�kM��R� v�U�jJ��7Iڙ�+-jʴI�6�T��kJŌ�Z�km��ZF���KVB�kd16I����5��s����ˡ   )@���Űh�ԫb�[�[��ͣ��l�]�ncT�[�;e�[J�h��f�ۮ���Ӷ�U+n�c��U�j���ծv�J=7,�3f5+V�؅�Ӏ  so�*�%�AY���s}ev^�����B�Q�}o�����'��{��{j9��w��޵Rk*}�Q��A�4�C}���+�Y*�ϥ������|�>�Ȣ�O*���V�b����(�U�   �y�� �۾���|�zj_V������}��N���}=Y��D��}�J-m�y�E*�ڕ3��z����(s�o�>�dW�]K���{�J�R�o�{|����}�d�k-5[[#m[klO�  	��*�em�V\}�=��UQoJ����L���Sͥ�����}>�R܏7{���2�����������Ͼ|���*�J����Ͼ���=Sܯ����wUkm}�ڙZ1J���ն�*��  -��%������i}�U|�}޴��U�wm�*�ޮ٭*}[>����B٪z�{ޕv���v���ϥT�^�׏�}��M!R�ܯ��O�5ET�}W��}*��F{���(�C����[R�  v�}���U*_8���i�Q�w��]e������J��*��Ͼ��͗�tQ�T��#�}��S��o�}R�RT�ϟ|���{��Jy��y�}t����� <j���z�6���ڍ�V�b�(|   9۾��)W��;¨:���� z�xq� ����@*����@rc"�;N�z뮝ޚ��z<op�C@s/J��Z�+��"��|   ��l:#)Mto9�� v8�C�0��Ѻ編 i�=�� (ژtw]������v� ,^��62��j�5(��L�@  ��|��i����c�@�� k��^x (���=:S���zΜ ����x ����pW�Gz�Q��m�̶��Mm`�   �Ⱡ �t^�ѻ '����;׮kҨ)�^pz����5���\ f�=�ٹ��z�   :    S eJUF` hi�� �{M�*J�      O��JUS�@�@    ��R��bz� 4`�L&� 5<�)
z��4���42 BJHz�J5<J����D�D= �iI�}G�{�����?WN�ԏ$$ ���4���bس/#3ex"��Ay՟`� {�6n����� *� ����QW��W�C�?����?�}*�T@`��UU���(���J��Ƞ*/�������|�F�0��2s���<��<��<��<�̜�2s0�/0�̓s'0�'0�0�0�4�0�2s'2s'2s'3�0�2s0s0s0���̜��s0s0s2p���̜�̜��<��rfN`�N`�`�`�ss&d�Na�N`�d�Na�93'0s0s1�L<��s�9��9��9��9��9�Nd̜�̜������rs&`�d�a�`�	���9��9��9��9��9�Ø9��9��9��9��9��`�a�a�`�fy��y��9��9��9��g�9��9��9��9��9�y�0�'2s2s'2s'0M�<�̜��<�̜��2p�̜��<��<��	2)� �
�ʧ2�(�
�ȏ20�0�����2� �
���0�L�2�� � <ʧ2��*s"�0)̀L�2��*s�ȏ0�� � <ȧ2	̠�� �ȯ0#�"s<�0)� �"<�$��2�̀�*<��2)̪s(<��4��0�̊s <ȏ0)��'0�̊s!2�̀�*<�'0�̢s
���0�̨s,�2)̀�
��0̂s�0�̡0�̠� �0�̨s"��2)�"s�əP�Q3 �ʧ2#�(��ʯ0#�#2�2�̤�2#̈� <§2� ��3 <ʧ2��*s <ȧ2	̪s ��3 <ȧ2��"�<§0#̂s 9�d0� � <§0�̠�(<�$��/2���(<ȏ2�̈��U�@ȏ0�s"����� �y�C0�s0�s�Ȅ�<¯0�̂�̠�"<���ʏ0�s
�2#̨�<ʆdNaW2#̨�
<§0���<Ȥ��2��(�!̊�)��̨�(�ȏ0 s(9��Es <00,�/0 s��0�� �
<ȯ2���(�<ȏ0�̢�<�/2��0�
s�2�'32s'2s0�0�'3���̼��<��<��3s0�'0�'2s'0�<���<�s!�2�s$��<��<��<��<�̜�̜�̜��<��0��2�s��̜��/0�0s2s<���<��<�̜��<��<��fd̼�̼��0�s̇70L���<��2s/2��a̜�̜�̜��<��p�.a�a�e�^a�y��y��y��y���d��d9��f@�^`�d�n`�9��y��9��9��9�$�72s2s��������~��<�y��!�B}L�#J�3<����D
ʻ�C&�V'U�s3Ee��@����$/{�NFF�U��k4X��R���KZ ����cŖ�E�]�.6y7�x�³�"3'i�#�7��\k`_+xyݑGKX��ʛ;�IR�W�oik�é����HyLY�.!�p�a���'%�0<��M���+��L�	Җ��vq+��\!�e�)�ׇe,ǹR��0)Bn�b��%�n�q�H'����b��n�[h�,��hKV�6�Ү�ԩ�Hl`�1B���ͷ��2flt^)�����,M�ߌ̦��F{� �tn+U���r���2�����4G��1��P%���Z)X�T��t&�B���KE�֕*[���ܭ���O0J�R�/i�jQ���p
�2�X{o�Gwj���c��lə*©�6������-&eLf�J��&]ȅ�4�����á;�ż�j�ı�;��I1�6٢�7E@�*dA5g��bOcoC��J�ϴ,[��L�zUMA�+�q������1
�aA��ݥI5!hU�˼�m.�2 X�B��B��L�%��nb��f��e��n�b�)�F=�[{GUJ�OQ�0!ĺҍ�n�� ��H��ѷA�8��	���׸F)�ZrI��m^�,Q�S*�r����D�+L[��D(d�lr��;����	��^���8�kݯ�;�.Y2T��P�r�J:���%�B۾H�)��]�Y�q�=�)-yD�z�<7�3��SXn��̎�b��=�R���B^&����=�"�,�@Fc�t-�[�j�)h�Yyj��X�/`82��øw!�Q���2�$Z�LrV��	
@��8�ҴӬ�&UЉ]
3N�#2X&9��9��;H���Jy�kR�9��,�QTv�3Y�Jiͼm��f�{�JL��:3n:�N	���5�e쬢>cTdV���V��<��W��1w[1�o"��t����V�uŨG��R�&���GnE��ĐS,X�(�eH��].�[��4��e(��6:�L��b6^�7id83�Vn�Yն���B���B�k׆�Z�"D��r�g&Dh��vd;�j@KF�V��*v��EeɓJ��<�+JZCj�D�jYk\�Pz����Ǯno״�̵ОQڣ�ƽؚA�u��j��6�F�I�u�vEjm4��C.Qglɵ"�w��Z�_��� �i��`��b]j�Plb�N�M܉�kK��Z㶫m���R<ٺ�����Er�,y@�B����GUu��R�ƹ�ڼo9�i����Qi����+u�0��5�����3V������	�:�kr�K:s-��3j`�^�GD'l�RCDX+V���1P��a�94��!K̙YT Ӗf���FE��n��cd"-�Y�3	�Cw�r��j�X��nV0&V]�{m���Ɋ��f���7nVؕ�l�M�k�5&:� �ݝ V�b��༢�̌d�"���[5.�7�7M��%̉�r��`{�L�� ���3���Kr�*\f�2�{��IM��ܥe؍���wS�I�%S�x^���E]�c2:�S�׀��@�ǵNTF�ۼ��uFۗp�sS%�՛bf=��UVj�cR+p;���ͩ[+���f\�l�&c�aR �)D��Z�e��SA�����-LN�9���jU�(R�mԨ3a��&Ἂ:�N�!R�m�D6:Xz�#
��q:35r�Dgʊ(��u�8IoU�K
YN�JR4�5en�L��PF�U�,޵�$�d�\�Y�n���Kv�5�6�huB�[>�)[
�	\�	aZ7�e-=ՙ�I�Y���D�=ۦH�&#��HՃ����0�;J��X��[�vcu���P�N�cqn�[�ͫ� ��q�j45Em�:Q�͠�,�AQX�j��jy&��(B:2��jڱ2e�(��ͭ�Gq��yK��c���P�����e9�B�fRҞ�[l����e����.��1��+&Y��).:���Q�{XMe��^0�^CC%ěՍh����u�J�XdmM�Z�w�ԤM0M���y%�P�B�a'�q���w70n�ˬ�Hd^�d�
}��1X2Ɲ%�u�����E��Y�A#G__n7o�ܔ��0��h�q��s��НE��D$E1/P;x1��Ӽ��g҆��6�hQ;Q��;Ŧ̩��L���A��W*��ti�`VK9��Z���0jx�1+]�Z���.�w&՜�A�I0Tz�-���`T���ź��.U�)�ܥ���ಭ<!���Ŝ��G�/���!j0F�OU�n�L�(����e�	j��x�'���Oe����[�w��\q���){v��[����������U"׹d�*`}KX�o}]�d	��ljn�'U���2�� �@ZF�D4/]���l_=�0Z�bDl�M�n�J��6ށ,)���v>9��3M"�wW۹�D$�g*�X$�W�,i3��#r�3	���C#��7�E�ok0�w�/k>��K�姣sq�m�B���`��n ��FM;�щPʫ-Z�;����an�yx	����y䆯v�fF/Se<,�����+ma�BF��MDk�����;�n�T[bE*,����\���k3s(.��8����{�I�Kve�Y	.�]1;N��Ħ�c���4�2�� �X��ңYu*)°���3!�AK�hI�'{YX,Jo-р�kq�&;�/�K�u(eG��2����bԚĘ^��� .���&�������-7���&�J�RM�12��1�ⶩQ�v�RÛ{�Vy�ɬ�J�Unf����XPʭI����X5��@s�zi���i����D,�Fk�çM1vsh��DC�m|ֺ���݁��.ke+��Ӑ`K@���S��V�.PF"�� ��la��r��j$�+�Z���9�A��f0�g	K)b�d�O)��rMSt�~-U�n�� 0���cub޼�:�oIn���Ye�r�ei����f��&CEѽ�fXz�h�NCy
����6��TLL���{{o��	�r����J8�4��.���wP�j�lxκ2�-�.��SɈ
�і��:C���e!U�Y1ie�ySq�Y7C'�ԋ2C��6���+� �\�w&CB���ăM2a�!�#1�-ɘ6e�8��%(UIe��M�Mvi��y�,m=I�����f9��wSkR�4��%�3 ��-��KuՌx�]2j�[���.	e�m������O�e��>�ƅ���3^4�"�ȭ�.��mȞ��0��2=zweK��j;��jsl̙q)�k5e��kiK�1���
��1��ٕh#{���4�<�|º��L���-DP�r�AԜ$R�I�:I��q�]���kZ��A��\ya��٣�AD�td����J�Kh��A*��!�ڼ"�h��:�d�D��ӷ���fWN�{�ܫSL3kIՊ������`���n�p��P��
�Ɂ�AD���:՛lѓ;(�t	l��,^VKR�o�t�)W!�(��A�٪�����՘��`Ƿ�H�#��iKBӆ����u�Y�a�Bt0�9#�se�C���l� Ae�{�|S���%f�U���U�u�Z��CLl�f�]���GXR���i7s�	��/0 ,�4�I^�m)@��ɷL� na��&�L��1e�lSoF2{���T,�{����o~xljs�����A����LZ�%YȢ�,=[V4��"�;���D3���� ���y.Īw3.N�ŰcX3C�ו����љ]�R�|B���u�E�U�-�����o��F�U@n���l�p��r��pfV�>X���խ�]��{{��t�A��w��X�{� 3NZ�Z�����A��8��3J�^���bJ��2^��F'R�Lۺ�m�z2C�
ǁ�j8 �D����)eE[���؟!����.hq�OF���-=$Y�t�թ2�gWRVήv.�/���V��mm��qϕGv�В��J�Cq%^�oI�y��ss�SAjr2�G7@1�`��a4]�������I��L�̋l����&����^Ǜ[v���J�`�[{SjV��^��A����Y�MZ��7u�T-��z$�/��cs	&�J��+hI	3�;X��A,�t̪�t�
mŏ�aA.�-�N���u�2�la2����b����h�8����F�˳0�?<�	杄8Kd35-�q41*��h���-�o���Uvͽ�@��y���im&s7v\!,��F�(�N�Zp�8�SF��V���g�j4)�f�Y�of�N�7/�d�e<�pEB�IP�e;���rL�4�WA�J˨�,7h�J���P�q7Vݝ�{�*-���^am\/�V;�.8�e`�B��U�ˬ�#X��D�4q��/65�U��t�M6zdF�D�w.l�A�{�c�r��OU��Y"�� ���/p�"�<��1f�|ͺI�°�*Qϥ!D'GKϊ�[���A�a�DZ�>N=�t���FG��^��l���r=�MáFV��f`��Y� �P�7+ѡ�m�Hs�/�d�H� �j����u����#������
��ِ"&��
91�&c�(�xЭ��C���;�J�"`�{0(��.�b6Ph��Cn�]�f8�gpa���TU��'6���Y�0�m���`"��k]��(^fc���]r�ۍ\F�!���E0ۭi)�H��1��uZk@���z[,ˏ��<2�u��F��c��yz�G�#Y��a��5C��"ҽ$��C>�l����x�Mj����b�WlM)�-�j<"��t��V��ט��e�$8��ɡ���zv�w�2ff���f]3�ۥ-ݬ[b�9��&����"�G�sI��D�w���n:K"��Y���AQhT�ĵ@KUY3vP.�]/�70�تXt �pe�Zd���F[���)�����J��Z���[�hV^����F�G%=4�@�����a���e.U�9��l���݇���ܒ�
��=��a�Ɲ��.l�2����;�w*TȦ�Y�*m���M����E2��V.'�.^ïu�Ԩ�C"������Sw)�gT�P��n	/si�4��D)����]�.d���jw�mn�t�b�{�V��䬱 ��2|╓)VSSE��At��J��14��-K�٧(�pJB�z1�7pf#j`2Ht]/]僋s�X�y�wB��`���ˌ��&{z��+���/�!�J-;���oTV(m]\��8´Ň��E
g
�*C�YN�_5b�葊�(�S%��mķ/\l����m�c�a��Ь���]L��WZ��i��M�2���2��F\��YBj�Z��D��n��4kp;b�=ٷ����/6����}�C.
r��q�:�<fDKTe���mU�L麈��6����ˠV\��
DQ�"m�A�R�Z�1�R6�q(]��9�/+m�E�t�za�V-���Y�-2+ˊm)�W��h���h��k5yW����v1TE۠�v7y1	֫l��b�靽��`�9le�8��Y�d�@`�Y�P�彼��Zh�S"��a��ű�f�ou�{��ϴ�d�A�G�^����.	<�e�����v�!"�%��>T�l#�Xt��	��^�m����H��P`;l��-��z�ƀ˂5��f�gĈ�����9Ah'.B��%%\m�HTl�wHL�p��m4Y�ƼNfec��[i)��pf��6omη]W��"e�h���nP��Q��Z��Z+øJC͖�G7v]�}s#*����Ql�[MK�P������q�|�ڻ�!q)WVm �C��F�M;�S�k��l���-�u16�7�Fn�N�=�&e#�Ut3Lf^B3��t`{�&��U��`�GrZŻ��4&�	�L��\X��ȥ2ti�UJ��"\�Ϥ�����TV �@��N γ/��ˣd-Z(+9���1oi���:v�k�0hD�R�@�ܘ�+��-r���bg�������*�E$M5pټv���$�K����|�����fA?�^ӿ����f4�!�Ϙ��K��Xc�����Ͻu*�	�}��~?��-=��t2�_<
Ty�3�k�]m,�KObz��w������Rm-��ߖ:ѵd��yp[�ʭb��J�lv!�:��+����Ͻ��g��k:ܴ%剈��j�(@�+6P�3,�V�l��@�731R�8]=��;��5��Ͳ�w�_�{3�3�,��^����İ��z�ؘ�cWnX�^yL���N4�ʳ����.s��H�'���)uggwJ��W��F�hw���޺kr��C�B��{z)"�/X�禣iP��]�"�{��h����8���3�D� iB�<;(ef��������bZ,x����5�\V�{Y��l��"��؈��d[!��������M 1���M>�������Ǹ������{ۻ_e�5��쿞.�FYz��2�f��b�{�W3|p $���[��j Eó������!g{�P��pz��38�R̹���|#�>����1[H�H�yY2�,]���:u�a*�^�w:c�i�=bZ&����c�=�c��s��>��i|Qn�F�����m p�� ���.R}CH�y5�]��C�55蒁ಲ�n �qB���4?�g���Ԧ5��i�V���f�4�e�
����Ȳ��V�*k�&�>NX=0���:ۧ|�ӗ�Wh���A�q�;$��Z����r��2a�Bt�S�}7�>Ncm�b�	{Z�\�3�9��l�!��맷w�r2�V<��r�K�,��{MvN���	�d��Y��r�ChL���t�ȫ �]�x�;L|�
A��އ�?y��NG��|{<��G��p�n���U����N�����=����,.]3��{@�<�����җ�ݙ|(���j��G��d@��=�'.>(�%1��`�e0�Q���������j�^p��3AU\�s6L��M�zZA���oݪn��� \���a�+z\�M9H}gv�:g��6e�?�-ٕ��3������Ĕiܧ�Y���z�6��+L�峣�˹C��Nh�a��f�gr��l �Ř�9�����^�c�%BD�\�^�s[�=/�MٔW=-�*�*g+Ю��F���EJ�r�ٙ[���s���V�0WJNq��;��W|񌊶G��lScEC�r���)�`^��qdz+v�v�{wm.W��X�Ώ��.�ǯ]Bz��wg#.,���etu�7�r��e��nV�\n;r�:-ۚJz��f]���j�B.X����syi4�.�"��C��I���
t��K�`�RL��G���)�O+z�8�8z����[��u�R���v�Z���%���I��n.�s��6f��ds���F>��⬥�o�pX8�t�C>U�}��S]���'�wؠ��5�r�#z��&+��L�L����ȗ���O�)�t�V��-�!Ur�X�Z=Ν�Ks6[�����dω �g���}��h�e�V��ڽ���胂_�ݻ�����e���;38��T뱐�
�p��u��|]N�i��rZ��#�3A�����C��f.����.�0t4��>��� �R�r������3��[�{��_{1��ǮY�r��t����X�	w�$T�ܡ3)�N�@c��f�𜮾+z���py�U�>ǫ��]5L��N;��s����{�f����@pٺ�,�f�BƲ���B��)�9e>Oq�U������)�����n�mDr�����è�4*�V�`�+F�A��$���cK.�`RXT\��YW+x;�K��+������
j��U:W��B�알+ v���z �o�ME�w^�h?��dk5b[N��)��Kw�C��:@+T�b��ߝ콗����b�e84,ݒ��]|7��STt]����v�m��V��Ф��W4tMj�vęV��&��ʲw<U,"�5�U��X���g塓�k<�^��> )�mԷIf��G �����2�>�vBzKd�ٺV��q�̭�cc�cwE#Kc޶ "�C��Bek��A|���'����k��x��3&A��GZ�T6�YG�f=:��v>}y��TMm�2V��/:���ݛ6ԕj4 
�Du�y3U�\nj�>Ĭ��B���*�vnԥ�h��[�`�v�Y�ڴ�"W��X[�B�nc��jv͊�S��=�m��l����̩s�Ǎ,��Ǧ`��kn���[�WsFp`�
�p��G���f'��+A�;z�v0��wV�G7JZ��@�BLF��n�Mp��_,(�;G�q7�cyv ;��?c�[0X˅2R�mIf��0�=��I���PE��|�
U�Y����.�b�:�V�
�Z*Q�-�l��u�m���c=Kl8v�gEtx0��v;d�����"]�]B�����{�_I�A�����t�dfEk�����g=;?m����ۍ��1m9]�yu��dVo<�`�(.3�9P'y�tnm�)nL�K��h�h\TK�d}���S�C��e�fv����@yK�,�+���w�1��f�^�e��̥o��B�Uˎ����ޕY7�9G:t�V���c��ږ<Jx�iܨ�f�\:VȞFz�-�b����)P���s��o�u_u_TUM��H{ �:�a�4[�˹1�ҧK;9v��Jc��4���m��,@;���0��xv���؎������b�.�ߊYo��ۿw˥��v�؆'���R�|�Yp�K�<�gep̹U����{�P�� �`�ţ�ڸ��4�o�*� zՅ�v[�p���]-�ѝϯ��v�P�Ĕ�s�Wf��Bol*��a��z*Q)�����tt;�4��ЪIo-n1���+��i�H�]�\���6��Ә�u(��gB�}um蒺U�	�-���1��e
�D�ʷ.I.f�T�&�w˳rB��d2;jEdYx�z�F)��*�#�rcc]��X�)�wD�v�1�M�;b�ʉ"�̻�%��r����qoa�K�\����f�sQܩd��把�(vU@��5��n�^Vl}��z��	#afd{���P�.2+��a�d�Y�э�(m��x����j�-zr�v��r1%���Ś*��х%���S#sDJ�*9wIn��jh�M�k��Cq������Cnj�.ͭ���
{m� ��K�.�M��������Cc�i٫}6gS��.a�w[��VW]j�ZN�)�J,Ҹ���\�����b�6�$qG�����n ��많���K;�՚�*#?m�wn�]�G�:�����T0��2��08��S�>yS9Q�����^:ݪ��:�^	�h���أu���7V�8DԮ�u�tܨ�ƞ\|��>Y*T�d�mnK�޽��<�Ո�U���
�֞�s���1m��t�(>��rG�C{v=�Z�C�)6�ي��9������S�l6��~�r�=�pl���V�]���	"$\�'�J�ލ�D*�I�,���D�WF�AЋ��U���ܣw�e�z/
�wE���s\;�ܺ���N��:�8��)���u9��kd����Zz�87��$kn��㌻��2�A��ܡs;	}awܖ�<�eݾh���|�MI�9�q/VI���'�%�l�b��w&�/�6m��-H�k��էt�&̚僦GM1��.�&gDh%M���=0�ݣyk�A��z�k
#����/��b1��3m���9�*Wuc���w���{��{�](�͈ w�uZ���M�������4]��pJ�]qPɋ��J�mӾ�n�Q	�x���aks�T�p�(%�5��0����Vp��.��v��������㗄gw1��Z��¦��7��']Kv�-_�M(�XcZ��rӄ����m�Y;��|�e���T��u��57Y���4&-\��lrC)&:�y��s����P��{l�XR��Ţ��(R�Y�2��b"���K��xGV*�Egm�k�;��Tѝ�X:=K"8��:C/ �`��3����<Ҷ��Q��c���N㘉K����DyC'��saz^�nհ���/Q/�&�A\���4Ac�*2����>WsUb��o�մhL$��uU`���)�Fxu�����)�.�l�� b��
>��ΫjJ]m�r��1��WR��X�Z��&��>�G�53"�tUDa�:�o�`;�y�gfPb�i��0t�p���v�$�M\�5��h���3c�N_e2�=zx;J���dy۴�7��:J��0Ǹ+%CZw5�����+�W���n6���{5��[�n�ǅ���Mu=E'��s��b�XM[���u�E��y�X�C�@�
���J&�҄}�Wb,��G�D��4<�Ė�gp�����q;j�o6\��ӕ�Jۛ�0h}̉#��s8˧ŀ7�ƫ�V��X��XKllD�}�,g�xUa/��y	��v�� � ����Ki���.���R3�-�S�vf��hқa*�j�\��������)֎J�YQ�q��c��.so��rKlT�Їp�K+8��R$��^r8+&k��"p*�̣���[�*��a�\F�>S��mv8L��U�L�s��س�vO�Į���-�ݎ݇C��w
Rm�K���Ys9ڄ���ij]&wl��C���ͧ�%t��hΜ䦟��*�0z8��ACAY�����f������'#R�؝`��[���Æ:�4��ٷ.���Z�.��t\���@��:�2-�6�OWX=����b��Jh�Ý
ႆq��tP�6r����(m��N倷�9̗�v�o#��N�V�Y+ �l�	;bTw����7�A0���vq��g4&+W�Ԓ��]@i�\'b�Uwbt�xx&��g��)=���#���d��t��J���Muw �<W�cd�Q�^ͼ�Y+{2C�u֩Cŕ5�G|���.oo���R�� �
��+n��I�]	+T,�Hh�)��r���0#��¯��܋r���ݫ
�v,��Q��sl��;n�l!)?��/�JiT`%w҇O��;��fs�e^�{	�<��M��FW9����tV͜#�T5���\�ZP���Y�^����O8����u����LiεnV�6m���K��=�̠,}�%d�8N8�Tuv=b��j'��t��pi�%���U�!������)_����]y�m��ly�V�{(h}/E��:����EQ��t5���(�ؙ��K�;���6G:�i�g�f\6t�1�bSi+��3�V�zA��q81���;�����oWX<������zb\�1� ��g8T��0;�I�U����"F�A���u$)�2�ӕ(��Ĵ����v
R䉗S%��������J���Ҥ-P]ٸ��9�WRĞ��3EJAm��Z�����$]��r�[y�t��ie�u-���5��`�v��;�,<1�#��Y6�#'����B���kP)(B�&�^*/w�;bs����_)q�7zi�n��Bh�a�K�I6<u�se�2�z�+k��H�v�ݓT����ʏ\�U�pB�A��+(�%�ȻsdI�GI*wV�[	Nx����_Q����Κ8^(��=�ۓ&��o=��Nlv~+��N��J�e�A]U�����N�+&�O��X7��`W2q�%b� ���X�>f��Q� �<��Sy�]Y�\�}�)�_u�D���3�(S�ؠu�z�Z:�1uh��(��ʑ�qu�U��A3����`��  �ɘ��!gu(Ӈ�ȴY����#2�H��7���I��D�p:�����'�h�sBD$�XIumtٮ�qt��Ӄ��3�<��u�'��\0������NE��X�n7��;�o�7��V��t�
��O]4���J��R!D�wR���;����*4��v�e���gʒ��.<��f�䇖=���%��-��.����f��E��%.E��# h�8Z�]FuəFh�9k�,.ɲf� rX)���E����n����\6�v�;�*Z�]�h�lnL7�<J������cM�,+9�0��s�R�\��J81�Q���b#4�vi���
v��ﴇKuB��xc��kY�k/$ 9vEF��ڈ��Arz0�l�X�Y�MܓV���Lš�����H+�k�k&|�s���4;���9Iosq�5��m[[�;p+�dٗ��1p\�B|��:!���X�.�d��,:Oym��_0 �W�j�7W]�
Rf
3qР!'Yz�Xr��m����XKi��SuE�F��B�ۢ�_u95�Q��ɴ��tғn�;)wv�:]��ǜ�H���X��̽Z�[A�����Iݔ6B�K��3�s�y�q�ʷ
�{1t��̵�jS6��n�34vR������hT�n6c]QX��0L����o5֜���k��f.�<��$�zqG7{�TT,"f:ù�f�KXۣ��o�v�=݈���c�ئ޽�$`X���y��f<]s6�B���ң�	�4gS5)�sD�2�n��kL�3�V�� �(;Z7+�A:k/	�3A���a1�F	T2sHє�`��58$,m��2��H4X��R��&�q��rٷ��Q��Gn��wz9���r����1����p����Y��d.e�J��K"�ґ�Wz2Z�b�8��7�A�7-I������X�qm��ʸ��GKs�wD1eǝ��/,tP���b��|���	�fd�ʃ��l8k�c���[��k��nY�6�۱]p����ԑK8�lo)԰Rk%ur��t�X�f��7i[��W�̂�ܶw�q��ڙqv){��p�gX��r�f�\�����s\9񩻴��B�6�sSV���q��Kq������qަ �98m��#:��Z�ܤ�E6!����j@Y"?�29�mlFLI��H�KҶU������	��w�)ү��|�ͱR������	bH0�]_[$�h%�v�`��Q�MA,���	pH#��;iĈ(�&BT��3�B�L*TA��A���A�؝ �EՆ؁Td$�P!K��)��3�JTP � �C���N@P`�\|cPi*M$�@��FF~lc7I�)��f1e�P�^(��YA	q�v	�f�2��@P4�8ٻ�����2ѧ%J:	Ӷ*��&��l)jH2�%
i�UŌNPi����JQ�J1����	�-ٯ�����$��DۄDJ�� m��N��(tϤi���
�L����A��(T�1P�ɦ�UƓ�j���	�E�����MQNؐG:ܦͩq��$i�c�B��gꅤ�E
a�?-���EL�_(*�U�#G���k��a�%�R7-=�FI�%G�ABH��F)���hD	Pq�ab����w��+y���+�w�*"
?�����~(������~�?�Q�_�_����Y�o����}���bU���V�N��E`O!��M�i��6�r�m	��ln�/���z
��mV�v�ƨ��BgYR��!�6պhIV�A1�e���3ӑ}��fCQ.[C�ع��E�M5u�[���5Z�k�w�p����Yǅ.q�QcȄ�{ָ9t���9X�Dr�q�i��d%�f�z�&�=� 80Ixv�V]�CU�=�Rq�S\*�k�Q̽��xcUܕEBˋ��pW9�t25�F/MY�7W�ݸ�9�-��^�=C�J��]K� ��ci��NbB�:�6��l����a0�\�*c�'C#�!6�1��,HU��n���p�D�ɠ�?l�Ҳ!ˍ��Z���i��q��2�r�t�Ms:Ѭ�K7A�N� M�PIn�F���s߲����oI/>�|��<l��w�[����Wև�2#m�֜��Z���X��@�bz4�V3�r����m'.��;��f8󻆗xw�:A��&6�Pq�ԟ*����Mo��20��I0Q��X[1�}Gf�Tt�"����֡l�dReY14F���\xv�ї�+��� *��9��F�% �w������yQ��gl̪n�	�6��^�URd��l=D�rw.�y����g���___������������}g������������y�ϯ��������ϯ����������������������������������ϯ����������ϯ��������������������������_______��������������>������������ϯ����������ϯ���>���������y�}}}}}~�__\�������{=~�G����{<�f����NLBd�\��mh�[`fu��� �k�kJ8�Z�j�.�a��a4����u�ӹ 
�x/�� �YW���B��v����n�9�t��@��"���.�j�<�v�c]ӥܬ3���X��m��f��$]w
:�͊�;)�P|�������K��4��ޅ�nJ�	��/�� M�g���sD?nԦ+1�s7��o\M	�(A1]��m�qX��������,o>Ϫ:�',�\b�J�{8��92�!�gs0��"
�[�q�lqqA�R�����4��and7.ͩ��>ǲ\
���δf��M�z�pN>�\��\�M�73����WŜ�*�F(�ۙ�74��H�V��4>��+�[+�ݦ���`9�a�R�ۭ耻�b�/E�#�c:�ޖ�h���	�vgg̘-8��.�+ �NA1hE�]�]/t�to*S!�X���]n��i�i�D�.��N�ͻ�*H���������gqL��б�����
a���2ar����ߪ�W�ϊ2��S�A#��ӗA6J�W��c�ƥ��E`��,�r�lͳ4�	w����M�B�����^�$B�r���L=9��YFIJ�G�Q2�pͩq�ك�V2emeHM�h.���5k���>?�����}}~>�����������}}g����������}}}}}}}}}}}_________��}}}}}}}}~�_G>��>������������������������������ϯ����������ϯ�������������}}}}}}}}}}a��������������ϯ������������������y����}}~�__^}}}}}|}}}}}~>>������{����<���
�F���R�piC��Cr�ǔ�T4�w>N�́f�Fn��C�����d2�������m`yl��i1nN�o_ka�Z�Pf*�y�O+�����c*;-=lLlV`u�ώ�q$��a�W{��M��q��'���-��xˤ3��K^�g:#��z�ё��T'Ε�\����������l'r:mP��B�2�z�ۏC�Š���Ҭ20ɏ+/��bR'MK����F�@��
�H�U�Y�9�Tf�;�'Յ��s�	׎�Z,�g�}����^s�Yi[<b��w}.��/�r����y��v��[t��F��(��kv�ZG�+�o;^M���FK�M��h-�.;w3w[�rG��N�qoL)�C��i�J�J�B�"�����4�-�����ut�L�X�"�5�����B���H,:\�\���%1M�NYu�d�f�����\�5���V.�e8���{i^�6�.Nr;��6��[.�{9[��"e�=�Je�7Sud��z�nP8d�˺�+��w��LΜGE+���j2�T�.-p�.�'\�����%_Bj�u�o���N�����,)l.�y�������~?O��������������������������������������������ϯ���������>������������3�����������������������ϯ���������>�����������������������������������________���>�����>�����_Y�����������_____G�������������~>>>�O�8�����gn:S��ԣ��U�>����������;�@�Z�3s3Xrlf��F�t7.�K�81h��X*Wnr�W���[b-ͽ �8��o�4�����VP����3}���M+A��f��N'F���Σ7���o��laFL��]WjoK)��:P�6��]�f���s���`�I�����D�/b�q��^�$�X�n�j�\�����|_v̽��_h9�ʍ��gU��i�ǒ�qZ��*�R.ل��%h�4I�S�u��>�ʕ���[��v�:��s�� T����X�X�Ԫ�:�KFNyE�h���o	X�����c�S�i��y�7�C.�0��0�E|����v�Q}b�U|��:�31�w��ąo���>;��ju�5���-'w3�t���Wת3�ӮW��<�-X������cO�4MKE�j�X�������%:)!7ye7�l���j���blW 4*Ĺ��"B�����%����.UtsJ��K��,�Gr[�:T���P��]��7�'�u���&��XA���R�G�C}6�14]�����t�?b8��͹7i�H�sz�'���WV�Φ���">d����G��=+}��00�Ra�WKiVo�t�F����3QS����/�]�G���}|���/ę�piPu��s���t�wo�B	�$�/�g*��3��tc��١ku�>���_o\��S��4�EvIHu3��}��C�[�����@�J�ݠiP�m}���!�Βᇸ�KFscz��̪Z�� �P���JQ�u��ѝ&���?��kb���f���'�m��W�J�Å�/�uFyڂv�;UT�T�ЩY��fJ[,��s9�����U��}�PK�i�����C�hI5�aRnl���:���w>�8��d��yMk{��g����ȯ����+�6Y�]ܭ� ��o���v��2�5@����z�{Rk�u�c�j
x�Zt!��T�}��is��W˸ũ�u�ԁ��x.�}+����4n���v�3Q�#��N�����H�=L3���he�����Mk�H�qe�$����S;y�:�m�!Cf�^f}(j�Ǔ�9(A�jR�����^cQs��i��zl�U�Nq�sb�����_+��婹�A��U݄x�_V;9�2~�:�۽����E�Νz��uILo�1!�,�{÷�6���S>5��Z;,e���J��)
�2��U#�a�wwe.#�bíb���������4~`rR��sל�x����U4m"���5�:�����Y�T$٪�4v�N�=�Ӯ�}�/��2�ɦV���$�9���Ԩn�2�|�T�����|ѧ��i�eL�;MU:59o"�&�N����B��=#ٸ�J��=��M�۾��j�7������S�O�`��7��ίAjɼơ�TyT�v��v>�;�Ҷ���uD��3Y��^�4o>�b�����>�F��G'#�J���j8��1T����;'X���1T�6�.Y��Y�q
��J8���"3�$� 6�"$|RMA3�eǫ�`�|5����Vl�Ζ7������c}KZ+塬�w:���cOS��f몝P��T�\+�ܻ�u���++�&�>dX��2�E9A���:�&k�FC�����"�)`Â�ޫ鴊K�����3�>	��@[J�6�4%ӣ�̽
Ǜx��:�5,9�-*�檴 4�x�����d�n7ںx�vxa���#%�$9��2&k�S�����w��K����滴����!ߡ�ހu����Z!��kl���JwSjT2U˘kq!�i���n&I����u_PV�\�"V�N������wk�Ǫ��2��P���p-r	�E`�+����V-2*�_LP���}p�ڭ��y�'h]��lM?��KX�չDdŵ����NIhJx�k�F������V3�i��f�n�\�EP�J�v���Z⻅1����Ӯz�c��DaX2�k��[S'ŧ*ՙAze�RL�Rv�`��p%�-�D(��.����EkSn�vMd䐃���f�L�u�X֭r�c C&��6p�ه�4�:�7�2:���v�8���ٌ�Q��fd�W�{y����Ԝ[e��3�I�'w���*,p1��;��m�czb�]]�ǯG=�܈�՝Zmm�V�\�$'m5R�ߝ-���v�Y�V�S�@ajV\m�9�X�`��4^ʛ�C1�I^MS���:�:��]���1ҏv2X�G��E�YrV�	}*���8u&�I�S&c�)��u��66EQ�M��ɧ�9��A��XWae���X��+ԙ�4�K�M����5�&��r�%���of&G��4�$��7c�����m;����.�����YYF\}8v��jo^vb�f�	�s&<ۢ�d�7�j�L�@�d�V��)q��P�������z��J���w@�9�D4������\l�[A��hj'@/{��d#*%�����X���
�"y��S�&��K"�ҧ��ꪊ1�Yݵג�qR޹2l��^ǔ�[[��Tr���r�UK�d�Z�2�f���X��I�v�����5�a��Τ��3>0���sm���]5\�&.w&i<P�r�KљZ��l��1��(�z�X[Y>�Ld��"��w+�ɑ�w0f��j\es�C䲙,�[�8�PWԩ��C��׷ڲP��nWl�f�c���>�P\����=�V���8ܱRNIW>)�u}�4�d�ڋ��4g<���Pp`͚;Cy����&r��Xr�A�ЩӁ�d�k�ҫ�j �=;ı�v��x��T���4f]hKs~����Y�
6�;����b	�.����V�;�rc�[CjJ���A�*��k�h�����,h)�@�s�WpB�l��]����p�噓E��/O/��2J�Gk5ZB���Tz����y)ӊ%0(c�ɺP��87]�B���D�--`L/�!gM)0J��*k[ZZ&��a�̤�aXc�1�Z�눊�۬c-i�|��}!�U=�53���К|�U
����HU��fN�����d[��1ƶ^ۢ�C�P|a ���ְ,���V�ڇ�z�)��zC�Gc���{M�Z�K�R6�b��,"Pa
���d$eɅ�˚����Y���)��6�	2�uS�]ۓ�F�E�V��� �c&�w�e�^�*�$.<�M�w[@�'�I��v�Y�0A������u_l�*i�w�i
��gPc�#����IW4c����_18L`'���vs7�g�f�.�v��Trgq�i�z�N�e�J��4nKK����Yi�:��;#M<fr�)&��f���x�3��X[Y����+~`���E�%�n8�X8{]��u��e����0�j�Vd}-���/V:�|�Y��Y�QXy�JI�<��d�T��M�Z��U�Lr{�@���U�BDc�u�7�'e��3Ml�,�#Ͷ+n��� �|sp�9��kJJ
��%��*�;V�[�$��A��t�soP.<�Y�^��J�S��ط��6�|�W�#a��LMm��22aR�8i�`�_VPg�� �w&,<̣�Y\[��v�=PN/`����F��=H�7�}��К{�K�8�X:J��Zx��A!�4S�ж	�G	|����@;�����G$��6Lp�ձ(�i�������wa�]p#�<�Jy2��o�'FD��۠�-��w9,�P�F�v�w��D��d,t�l�i�gnf^����QT���<鮜�X�Nf��"��Q�Ŝ��K1d2�S�z�}K��8}˟.=SA��`�'[�V<��(]�a=�{3$6W[�ᆃ���Q��v�����r��_�K�Wʃr�>���Q)ð�uҶޭlȷ����8�8ɥ������c{��)���$L����n���/��	�Wc3�j�@A�����o!���J����jj\�ARʗpY�~�]�S����QZOU$�NF������!�����%�l)U�b}��k(HٳTƬN�˱;1t�����n��9��	�d���ʈ�e`Z*vq��ͬ���y	W���-�Nz)-Ґ�Y�ݧ��f���v�߲vE�m#6.�7OF���dc�)s�|��.K$���#�Zsm^�g8�ٹvN	/"m��TZ�����$���!k;wS���]d��,3��;�'0��lS�Y.�k5t���T�������sf���O,rz(!.ȡ�dJ���)ç[�$�OMr��l�����\:J�x�(���E!66�$_�+X.�;�7�N]��c6B憅]�b�§;��y���qic
��4�o�q�-��6���ף~�v�ə$����Zz`8"��;x̵w,X�(Mf��YWQ&�s�ok&L�(��ۋnS�7��LybG;5��H\�>���n묇2���!ţ���Y�
�ZW�NZ��7/�K��� �2�YُPQT������
��;t�B�g�]V��%�Lm��3V�;zk��6J���M�k�:�저h�r�
�p>㵠,s�} ��*�����˫h�Z�ռҒ���6�&fp�[�%|��Q��ΚV�6�B�>���U#�%;X�T���s��ۥ_�h���������w��W�?����G�����wm�uo<���,���wm�]m�g�I ���)J�
���c((���?������ɟ�j~��=Oױ�\������-)6��W5� ����KO&���;wuĈ�n8�ǄbQ��.����%^�o�h���8�wi�Ӝ�@��o!QoV�5l+��v_b�s�ݩ�j��V�ԯ{�@�3'q��̤�G&���2��a��v1�loѹ���v�5&���:� ��0��K�G7^���]J��ԑ��ۏ�]�鮇�\�b=WoI7؃|%�Ѓz��;��\��k�I�����*ͥG��42��(
�V��{:���n"��m�WP�g�W($�J�MT-�4��Z���Mě"=ǋn�l�Ct�n�:VE���<����F������q2-�V��
��I��I:'0�=�bCE�a�|�hB�.�ǁ��'%v�X���ތ�[�	��ct����2� ���vP�gx܌$�*4� +`��^eՎf���eʃ��j��ٳ�2�,���'�#��I��{���9�K���:���o]��k�q�x[��+h�y#]��0#��zN�%���`�7�ɋT�{�5p)������CuS��P�s��Q�Ѹ���Ud;X�۾��5ћ���"�/�k�j|���
d�!�׍��Ͷ����W^u8��<��(H�KJ�h�!H��O�ӑ
-6��!$��,܊f@�bFI# P��jF��\��4f�	)���6�_ A-�	�b��D�kA���V�ݨ�i;��ݮ�5����m��>>�O������~���g?�~�mu����筧A��+Wgu������m�/�.�EUA��y�?O��������?o��3�Ϲ���Z�l�h(��Z4�N�4�MU�X�n�h����9�>>�����������fs��?b$����{�y�8�F��Uэ���yc=�o7��n�k��ø�xn�y�^b �O���]�]�%�F.��	�1ܱ�Fǐj�p=%�b���Gv^6����4QA�wf 5��^��:�쎶���+�P��l;e�w�ڔ�@Xغ^���R�!���w��y�o9�˸Mi��H]��/I��`�����ݹ{nM�s��o����k)��[l���Ó���$��ן}�#ш��x���K��3���ֻ��]�7��니����7n����GmX���u�"�n��|�ysk��+y���I�&�a��:?"CeQ�u����.��*�;��f� �(�<��&�/�-�'�	/�n�
Q|J'�	6�j6�KSy��ڧ��DE3m݈�ͺ�`���i�F��<���X��y�WE|ڎ�뎤ֵ�c�q��l_-��F6&6ֵMF���t�-4^n���Py�NH�rQUO�ԄlZ>l��w7��Vx���=�x�R�g�x&�g�7��GI�Qj��e�%s��;i+�� ��8�.�\�lmw��yZ�}_]���Ʒ����AQ�e$�FR�N+�^o����:�dJ�D'YQP�n�)����י]Nr�����4;��U�^�Nh58m�E�*�H��gn��z��3�����~��_��;�<{jr|���Id���=A�ۯ�wU�`��5�.�5{�C�>�H��_���d����swll�-9��n�
Ϳ{$��Y��������'��}+���v~~���Cܺ�@�x�*i����H�=����::���Y=h�>_z�Ћ����Mt$O~��{�(��C��?%=�9����p`���yF��χB���*h��'�S͎Ry�{}ǈ����Ņ��w�P/��
��V��+��K��B�2�$-|���l�|㜷���~�=�^W�R�;�gۙ\���􎙭^uw��䆳�^J>���Uu�щ�O�*C)����S=<�F��z�:��n��GV�x{�F� ]\�����.�K�"kI��z���m��7Ɲ����1g��Ql�>��XO�s�t69|5����t��4-��v��zV�s�Hqe�����`���*��1�]�:�>����g�{>
��^�)�<}�_�[|�ٻ>4}O��sޙ�槾��u�֐P�G^�9�}�_F7���d�^��,X�B�>{��p��v��25Fa����u�C�YW^�{��u�%�Wջ��2R%X�T�9!�K܋I{]<v^��>�����_�g���6��L�>�^7�#Ʋ���S˽@����۾�}s=`?s�a"5z��Q��ި^��~��ܟJ��g�/�~"���wq����k����2ȅ��{Wx��H��t|�+/~0��j���te��ޟ?>������DsݟO4]�X���o|������#~&�j����)XV��;	y�~�������d��ao��$��9^�|o_(t��G�Zww//}�[
=:����|q�t7�h�a��w�3z�(62�����~�J��|�>�&��Y��U����f�OݣGv-nI�H4�����f|`�x�VP�iu�-��C�D����E���Mf=�"��_.I��5�V1n�|��/=���{{cW*�c[]!K,��k��y�-L�j�Y�`��nm��k�x'޺��z��<�'����9�4�k��왨qQ�HcDY�ˌݫs��2ȗ=��<")��E�ͧu醤���^�~t�fs�M�%���+��'��8}�,xg:DO�z=��q�o�>)2�}�ɾ���½1�E�o��@�s�(��k(*q_���~��9��P��-�ggN��q�ڻ;�'�.w3�{��v��~����o�}�������/ʃ���r��UCϏ�'�d{9�L�L�.����\Fhe�*"�a���r^�T{�g��lϓBs�E�vh.�{�{+@R��~���.��Z��>��)�_Zٴ�=�r�{�/jj�Q���@�Yꀇ׭z`_!=�˝am����b���u꿏�7�S��<��vr�|�G+9VW�ۼ��m�����|��r�UO�.,���p��-�p��3-��TD`�߽�v���q~=,���}�F�;"�;���!`6#���E�y`.��wk���+|~�E �EV�v���\�kj��K�����P�Ʈ_,G�v^� �)0ж�V��S�Z@
֝WtM:R�fK}�2;�iƑY���?:gfq����̠���lg�g��q޵��Kٖ��������W��I4	�����9l��3����gՌvWS$�}��[�<��M3 y��1O6^���o�<�O>}^\O�]{��0����=����D��W�f����B<���>譵M��NY'���Y �ca�ч.�}gv�����,D�/�Ts:J=^۝>�S��X���C�ۻh��]Bq�����.�l����'����Jg����w?s���\�#'-�rʧ�/_�ﭟ�~�y�	�X���3�����W�����Q7tK�s�����I�rwx���y^���`*_�5�L=R��g�����i�lMǇ�3�{(�s4{Z��̯+�>MAӰ�RX9��K/�ՙ���pS��<�|4���{��zj�s[����Q&:��e��S�/PX���c6Z�r���8�᳍]��-�K�@u�ޡݻ>,�vF���t/U��8�F��I��d��	[b�x9 �*	/�y���v�yn*+[Gw���Iz��;ٶv����E�I�ʣuL�!/�jD�	ц�Q�?����.��o���[۠�%qA�!h�g|���S�{,Z����I���v�G�ӆh�8fT7���6�Ц
B��.���k���5����ڊ{����獠�+��}^]X��~�W즈?+��>�l5���ΙH�{�v����t���~��x(�)s�:����5jC<?���S���b�~��o{�+ݗu�^{�#�S�K�o��pR���a�B�s�g[tj[�d���|�x*?m�G(���i�ޕ�vyOv�i��=�q��3�Δ�v.�xM��5\|+��4���MU�ؽ�u&}����LF �D�����j�.V����Z���?@G�J����=��d�}+�d
����m4��2���w�VJ��js�-���y����j?��WS���izM����o�n��T��H|߼W��C��;��f}���W��nߕɾ�.�\�Л��-�N]I���Q��N�B�k���k�3l[�����|ѥRt�r���|��:�פ�g�J����Җ7D����eZAu�%��
��T� ),�w	���w����8��M!:5zG2l9|�����i�}X�'8�~���ͳ�:��>b��{��*+e�}
���d��yOx�bz�Y����u��b�O?K���yl��O��w����et�Csk|w):GE���0�㽰���ֳ+�A^rrs��_��+=l<�������f?�o�O�AP��K|_�![s��TLt�~I����;�fz[wޭ������<�yb^U�AO���]���B{>���nq��i���y���A�}�G��8�L����ڄ��&�qͣ�;ɫ�W���(W�w�އ뜋����t���#}��_���(l�^e�B�8b���j�y�^ue{_�;�?P�(M����e���t�����x1I�����]+��E�м����ꊽ×�����*5ڛ�4z{�XֆOc"�!��s�u�|��_ �wxe����NT���z�c̸S2���S�`C��O^��ju�)۔T� ��ŬU��k�6mZ�p��ڹnH��u:����C"j�Ts�
�r*�6j�i��}F��eV�YH�T%�wi�wyEU��R�u���a�S-��(�-����]b��=����������΂��7toQ��ٳ۽w��۷Cwt����5�N�~�fcu��Wν��u�C����o�-s��.O�'8�IZ:{G�̞^Y����V�ُ="pz��~"xf�6V5f�s���o4Ad]������O�H���Z����G���v\��V�3��EBj�kٝ�W=��䁿+��<7ex*�9�5n9���zC^�&��y�נE�>3������ϣ�3�\5���u�3��/���wu�:�Z����T9�7)�UӬ�9�Qǟ�7�T�"'?{ oݝ��[����Q�wv��}�G�����hǩ�+;k�4�0��ټ<gY�H�s��,G�ܺN�\��{����ܮ�=�N���ʪ-�{�$|g0�+>�j�ӥmX�=뮣/�7z<!��R�v�x���\D�IolN�2H�u,P�+��Ĭ)b�o�y/d�w����}\o*{�H��^�.�-�29�e����6!3{'<a�Q�4��viw�(i���l�	4�������=�^�<�uz�{�+-��j�<_�_-	��7ˠxT�~�p���\䘚\j��U٘��e�n��^�ez迪���;�,_1|>�m1�˗��W���w�����6f�A|�cA��;f��ЯL��u��~��c�����J��!;�z�rb^�b����K���ў+!������9r�t�c�)b���{<گ}��@���w�zm����������3N��R+��͝fT�L+�U9��)?��ފoE�쀪���/�a������G����ei�_������f��7;�����9M���v�� �B����Yp����*�߆�iO`�w��t�}ѮM�$�P�YOtƛ�,m߆.�/3}�qz�UT0Wx��"�o�v��a��z�0����d�`�nT]3[�F*������Ez��s�>��	M����%�4��h�B^"$5o*�*�<��}Y��WH�om��f�9
39Dq����<+"�2�nZ�`#�]��"м)��6�"��ذ_"�Q��Z=�cW|��� ��:_	]�f2�DM�P=�����$�V�3���;O����>��a��1'���f%,��Pg;o���{�QJ(�2�3ҷH�d������V�� � d�{ه;0O����b3z��vV�A����q���$��ݰ �l��{��<�&��+����u������"Muш�ѷY�#�Wf��U����<m�_}�7/�����׽�#�������꠽�j^����zv;�P��\��ޒ/�܋�?��s�+�Ύy�r����鲛���I���'��<Ip��8��ܛ����l_`�J�}��zX�od�w.��y��<�������z��&�\���毓��=<&T��0=W ��_9W[����>�� lAް��}5��O��OE���~��s��\�|�\�ԛ���/>*D��:�,N���M���3~��@S+N�=ޮ�*���}~Zhq�=�K���U ������y�y��o��,zVw�wz���}Q<�n!�8� �FfuO�j��Uܱ�h5��Ƃy�x�[T%��DE<I8,��pɇI���R���d�4K�{.
�+���}(�ghSG���D�Qp�3�p.����_�c��&�6,w%�O��39�2���@��S:����0+�[�_�f��}����k�㡿�}ӻv���[�v��r���{�_�W=i���H�7{�ɐr�g���dF_�u��{{6��HkΫb��j�Ǩ�g�데r���g��c�I��ׁ���f��rsk�-�:�=��㔤�<��u���
�w���g���]{��W-�l�y=~�yI�g�˿�q>{��|����=K��|�>1Y����7c�o��1����>kۧA�ͪKǽ�_�t��y��A�#���[��]���>��'G�٨zy����S�3N5����}�����Xf��d�Oo?������a�L����<"�w���R�����+�܂~�O�O׷���!V������};<��^���ڏ��Z~[Ur
�nGjf�h7�߾�^�w�/��G�������D���χ�o���߿������D���2���W�O[���y\�x�-��c�XcD�,\*��s�Ӑw��*�k&S"���yK{�u�@F���e���5�,_wM]�ܕ�r<k0�� 젴T���G=8Z���,�f�5�of�R��:�.�C�K��'\��;s�K{CA���S)&�����%.��HιI��	U�S��9L�b�Ц��zi�n���5�v3̉�h����X��-C�'���Ƨ]n��]�I��{���J�(z_4*�`c[$$�9�x⽚2��y��xל��]��?o!�m�5,����نA�eճ�
���m:�n;A*�H�����3Mb�*�h=B��{�m��`�Ek�uɃ�=,�0�*�b	m�$�ByZ��Cc�����6-�²��R,�R���o]I��]M�}��W��J����q��Hk���m�a<E�����O�a�:	�X5��\���Z9�R��\M���LN�u��s�b�f�91czq)��C��f�]t��ڟ6�� �<u�����Y��v�RڽѼ�ˎ-����k��z5�����.�2u�؋���j��tp5�g��J����9�٤)�.ڙc���6����3�4�zޟyg84�L��)��U�&e�ʷ$��[�t��]�����LJi�z�IWW.W�Yz�t"���c��"�S�)c3z�ڃ�"�����
b!!��X�c���2��uWT'�ҷst�"(�./5u}��mY<͠gc-�ᴞg�U˾KK��Sf�yi}��$N9���P�5�v��/sp�6�o9����kuje�ʃ4�vAo��������7ϫ�����Ԩ�m<���r9�E�0p6��o\teʱ�ƜtJ�t*�n3#%����@�;.��ֺuF�y�0P�f�l7����)�(�@��i
⪭�#6����ź�cs7I�nL��eը��+�t�+�dW� 2���N;��W2�$iݜ�P{�.�Z׸o4�yt*��U�	p�V[�Gq<�zD�䘺�Žu��e�!�o��Q����BN�ܨri?C64MvNY`�HDy.�S�!B��sV��s0�9����u��f�m�+�l��� R9V"��H�F�u�K&�ɳH�O�� �}�c��B�ލ�U�uN/6p�h-�i��eU�wZ��}�e�Rkõ��i����Ĩ��o�&�$G(MǎŽhd�u�\��c_J	�˒v���s����[���V�}.����p����\#0C�!� =yn���,��m-�s�꧖����K��X3!uC�$�\��h��]��5�t*�/d��V:(��((5iޛHgRx/�.�b�s�}~|�N�:�'\Um�����u�u�T�5�w��gF��7sm� �g��g�q�ny�?���������3����9������4�E��ğ��t�4��m�m���<�Q��lkN��?H5�k����~?�����<��~{�CEtkF�v;q�v��؉�������^kG�;V�A��c[��y����~?�������������_�b-�V6�5����-�UsV(���:��ƫb��tu��*��\m^X��]���h��)������+�@BQ���+11y�mE��qWN61]8��87o��6�cm�����.ڢ*��v17|��u�~�s�a��ۻowck��'��^~��Ok8'cF�[kA���������cl7ͻQjƴ���UA�]h����tM7�qQw��M%EѦ��y��]b��ky�^l�]����(6�1+i���b-����ƨ(�w8��tf<�]�QQAZ0�t��1�G����{fb`���փn�W��G����Ѷ)�͊�Ɗ��w����v�7�[�*4��u+�'JK�QW�^\��b@ɜz0gv��l��Ƕ%���.v؎f�o��+�;+��V�kØfr}�~}_>|���	��}����� ob=́�T;���Ҩ�v��!�卟t�bl�����؉�UJ���ف�����| @t*���-�7��nHv���CV�^O��H�(ͷ����Ob�^��@�N۴�Z��%`@xI҃�1��i��Wj�BD�[-ܟ�p���v�P�	�O᭑5�9�\�S��ϙ���kғx�˺��P��&&���o��Su��Q�Nd��U������+Z.f���b�r�L���WW,�a)wk ��eӢ����P|��UI��|��n�H�Lxap&�E�����p�4��E�ɧ��[� ��G:[&���M�ި�3��|���vb@�e�	f����ߏ�E�w�EzHv�r��G�~#�,���oCz)�Ys�]��b�
l��S;�g�l�V���е'����a �}���H�� y2�d���,����?��4���}��Xοfַ�7����y�7`�>L���T�^�(z��ϡ���G����/@�x���H=�@CW����dOݩPY�.�;hZ�����"�=���q�ʦH����8��Mءւ��9Fk�@v��'|�d��;f/
~ר*.�s���芡�SI�!\	��^锏~��ϑ�Ե�wv2�g�0w���W�ql�gaR��m�)�zk8G��:ݬ��)�l㲲��1�E1�j�PZve����Ǖ�b��K)�s.�vl���ꧧ\d\%ԧ&b�����|��8y�G����/!�3N�{�)�_��'Hꁲ��&!��a�o�<:l�ŏ����8|O<�s���p�}��zz����ꪨ&��m
���NP=Yӏ�W�f�X�k8��@a?=�B &����<�	5��70�9=�-K�u?�@�}"�e8[�N��[u��;IB��ĚX��H��UE2��(T=d�ZK���N�����B�������S�oi0-��Ȃ��Q�K�w,f�'��	�/H�=(�Pq}~m_?{�^����~�~��������m7>���/������6��k8�&*�]���{��L�u'O滐��?���X"�+�vz�h��H�{[ek��+���q̆3mf:9��	������Q ₱W� �_G��##=_	S�� q�g�+̴"}���~����MiM���q{Ѯz����v�F���Uӳ����lP��nf�B�ՒS�r��-��B��W�Z�kZ�^�h(���]��c`.� �l�`6���'�yI��T�7��^�B!'/q5#�{Vhu� �{#¦}��k�c�B�-�j"�턶�o)9�َY �l��7��9��iNb�}(�ArFl�!x���aܝ��Mu]f�qGs9~����L��9ؗw�s�4���v_S[�K^|�[�.�O}�vj)�E��O��b梊��Q��ke�e;=	>8ҷ�k&0�IfYgt^Di��H�c�޶��(� ,�@Y"���m�s�q�x_�����ϣ�����?�z�ߣ����?���>n��>|�=����ȩ�s6��M~O�kb��nO�bST�!dݬ��fC�F*�j�ڮ� ��`�'�M��)��q���M�fR��`P�E�f��*|�ܦs(�U���]�7^'^�:� �2�7�A9Q����2��J:_S�	�	�[H
ֳn�m�B���\��R��25����0��������M�E~`2ݛ��L�r��	Ot��\B�<����=�|#������ �y��Ic�>C�����hG��,]��Y@���N�N�$)�J�˷���<+��x��=־��ڎ|#�{NiT����e*���G[6���"�l���^��!1�nj���n�{�бݛ�og����O^��1(-��Z�Z���t�Z���0��"�w��������OϿ����c���n�L����;ky1�To��O�Xz0n����f��f9����4Ѯ�Ә�.�U6���`�$�x	����i+T{Q�	���5��n0`8@Y|�x<M	R���8�/A��5r�{tlRC���s������ȇ�d��ooS��>��.P=�"C����tyY��hW��`2�<���{j��NS�/�9��+��ds�tS�Gt�k�],Z�e��a�-Љ+�/0��̄��o�8��;�:*�;Ո=��:5�[�|cᯫ N2+xce�VKw��2J���;�^졂�.$�|�]������/�3�	��|?>���w�~�@4���>py��_)�(���:NC����Y�rk�>p�ը[QX�S�Ójx{�b'\����w�F�$��: �{��%d�x4�f���L>�o;CnQ/���k/!ܱ"���'����]����}T�R��M���Ӭ�� KH���m�>ۆ����O3�I��G������g���[���TS��*��{p@	�8�L[ڕȬ}׽~�~1�zu�9f�
���l32�T~F�J͘<�� �_4&|��C�w�O��@Q�M^�X���ȷɋ=�v�Vp4�>���P�U�=�r�U,��홵>B��.Pd�e����g��7yrX��vH9�o:;[.��| ky`�-sU �K>��v���q6�emkw����0+6\Pw��P-�p��Ϣߩ��Z���oEf����H��f�s�<7�"7]�ڭ����y�.M�#/�"��U�J.��n�7��p�Ȏi��RlMc�'���C5��ŭ��,6}܀گ5�{�� 25��x��_��]�z���������S���/�ȼ�6z�����=ndn�*'�x���@۾�o�n�`5Nzu�p�f�5�Z{�D��biZrv����ai�>*ĭD$�LH�.f�֟a6[����b?a�U�\���Q��Ui`�7��yŽ���Z������Pek���9�ؽ���l?>��>����~�#����;}�����( I�V�60���N�t�C����LL�ډ�K\ 6y����u�ӄWeVd����9����P�@�e�͛!�X'm�嚯Οt�ˆ�x93{V�nh�c3��R��[�R�SOY�3Lza��´�D�WS�����*�.�T�Ut�k�m/;a�˼��ն��yβ��]zk~�/|���'�G'�����x>�0�$C~�dS�""2ًd�k��~�����^��n�{����C*1�b��t�k�=������mOU�+/dE�-�h��^׳flMn!�xm)��҅�|�Tk1��.���m��瀛(���J�.+6�!i��U1��O*��U�`���Z|鍃<�ϟ[��ǞNj�Z�a	�K�|�ts�=Ƌ[H�}�2�]K��h�H�o����,�d��`�S�,�o�*��ya�Ǖ��h����эG���mx^*l�Q��x59O$g/o���z��%T�̤Õ"�U3��ۂ`ZwSAswu�g��[��h
��u�^�,q�f��M�VЈ�zI�G�f�EH�.nD.|�碞�&����ys+Bt�Ы�V�Q1���j"i���j��>��o���NU����cose�h#Rf�ָAJ����,v�zͶ��sFSX�l9����n"�/��J��̷a3t�ڂ��v�-�O��0��#y�v�������?�7����}o���6<���Z ���7W��i�$�p��F�-�O��E6PNcݕ:�{�}u�Voh3���-��1��\ScP�2a�c�h���8��+P�:n�1P�ŵ�%�Z
�84��M]Oל�W6P4���p̊LL{oqO�NȺ���}bǙ��Msخ�[�iZ9]�{��Ux�����!��-ܠo���H�/��@�Z�ǋ�c����O�C�q2VDA����\��P���y�ؼ�nkm%�>�I"I�a��� x漸|P���"E\�S5I�:�{i�n)��)�z �arY5�d�,cԃ���1��Ǣ�<��nk�*0rM�퉌���q�4{�:�Y]�M��^�*2���v�њ�zҥ��O��'�<��(Lf7���[.�ތ@�)�a�:�|�Jy8k�{8��`+�:Di���L[9�E�����v��"���6�M�������*�"�m��[�m!>$�lW8�G�x4b���T�T&[^����|��|��X8	���SHv�7�h��ji�p%���'����wz7pW6=��r��7߲��J,����%�9���㞷�5���ka���W�>��L�	:^��S>|��$
��n��đ����I	��w�"k��+Ǹ������b�5�Kv���:�D3:"Y�:�����(٠uH�"�\�V���i�l�A̻#*�e�q�xy��瑱߿��>�� �37�����^eA��]�����酭%r�����fB�p���D�������)��)�5�F�3C^��fi���L���X�Y�AWA��w[���9��<��̑>���Bte�:���qh�Ɯed;M�X���FQ��Z���q`t�㚈�W��7�`+:�W�sY��25_��_�P��{�5d6�ΞW��|�c��ۦ[MN@���=��4��R�ޙH�4c�Uk΀�s5��˰Ǵ�dǮ�4x�`�R|�b�ٍ��V��bx�Vi��[zG���7�N��4��g�'���=u\��ZK8�p��k���&�I��4t�5v��\�n?�qV/_�e��zu�IA�,��� q�N440�ٙ���9�����6����es�1L��K�`b�P�5�ɋ�*�%�q�Lp�l"����#b�(��И�\/�w�.��!v�{l3�M&�-���J*0GG7RR��*?8�>���/�;�+�Yf��JH��!0$��<�"ɡ@���S0�L��Zh���L`}ȓ�׿#_��$I���?[Eg;<6�չ�iI�_h�
���w�a��iM�t�kѿen��;�ͺ�n�v2ЬR��C9�vv�A����X�Tw_s��Y�a�k25���źéB��9Xv�\/���0�`],�o�
�qm^4ԏ��<}��<@0�!�T��>����z������f��eLBq>��.�T{`U�~���Ӊ7�	�w<y��RX]�>5\��,��5U��O
o27���8��q���������jr�z��H�&v2	�����fl���.�s���TN�[:z� ��1��X&6�C�
��	x �q
1�h5:;N��e-�NB�pK�R�<�U�=��`��G����<�DyQ���18Ϙ]�l]���`��=HY�(W��W���I���۔R_Pݔ[[�(p�d���=
/&��d4<������ݫّ�'ֱ�	���c
�kg�L�:z�ɇ�&��U(�3,��9v�vL�7^�A�8�C����O�R�%�+�M>ծ��xiqW�	R�Q=��MyX�X���0���>�g�X�2sS����q����Lf��L��ۣu�Sj>�������o����9RVbVlϗ~�Q���;��x�^3Ma7gӻI+kr������AD��_ ��Ve��-�xy�f\��p�H�/�3�Ö�_�z�㬅��%�j�>��p\�ŀ��tv⃣b�[֏N�]@)��r���L�u�0ν�����t��0xO���1y�CS��[�4��>[c8��l�4���͝X�u!�nVL�K��W~{�>}|����;�(��0�0�"`�G���=���������_�����L�e�
��:/ڢ�8+�a%E����up�4�O����.(bpn'��V�ù=�z9�"F�\��j�0��]&'B�n��m�
�6�E���-Z�ST�b�vA���[ ��	�#[j��}�T.q��x����؟��%+Y�^va��x�h��XM��/��r��a�o��qڴ�yc��1��k�����b�W'd���Y�,֙x��nۖv�4Me�d����B��ei	b���?��Ca�a���ø�y×��VS�qs49�m�f���::�,V�P#�FT{�QV�0�XT\2bW��I��U�f[�4��u�$��ߏ�����.��ni��m?�z�e�i�E�"Q�d+�	�u��TTQhv���Ӕ�ϓ�j������KuE��������o;�u]D�/�$g7�w���˦�n�͊X!W�*B�/C����cks��+�A���ރGy�?mDw�������2��"���<�.	QX��gٕ�������4q͓+��tr+f:��I�U�7z0]�˷Y4K]�aⱗ�X�v-Vm�Mdt�g���_i�o1��")�������|�{�����y�$�g�V�g�����3��ؾ��j8G�J��F;(Fzu�"����~���?���`��L0��D�JI��=�������y�>}�<�u����{�e��y�(\���o<�h3���?�؞�����E����C��ج1}���2�Җ˰-#��W�(%���r'D�TV���T%?���En�l4��Q8y����򴥱4	��m@ο<��C�4�6Ju#�{zG�\�����xOR��g�u�p�H*�ױ��1�d�n%�+Kj�m&�ׅR��xn`ˣ�Fc����)cS�enS���m��VFy���}���}�L��W�<����
}�]�꠹��z���V��\���|׈X�I�ܞ���C�}�`�TgPO��C��E��ffQ�P�i�G���;y=m�H��Y
�s!j�%뭽⤆����y]	l$�g1��c�㑋��֌���Y��H�l�4��r�P�'(k{A���z��
�kץ�ni��2i��ꆄg�R���Y3T{���u���g�;�^��q����� :�?b���u��WڂKHN�t�m�A��(��;���C��j+-oy���4�8�$Z�
� x7���<n�����Emܞ�`,=�2��)m��J�f���h9��w�Li2+}�X��Z0P¯Q��X�7�g���O-l��`yL��-w�m�å=8W7%=l�ͫ�0_n�G��rc��8ܗ�@�F�ws
�R�Μ�
M�n�hM����r�϶��L���qs��T
�>/.��9*�� �mi�s�b�����V��˺.&��r�L��"{�r9�hV�X�d�]�7F���w��U�Tf���<�OZ�]h�:nL,5ќX`e,;Һ�u�!�1C-Q��.�h�b�݁�Lj�X�{��u��I*|���Cv�WO	��%o@b�M�B�3�^\׉��M}t�1˚)�[N^������>��V�.����DE��ܰi ����F��Q���l⭮k�`:�*Elj������x�w��l�s�#4��<��5뙲�@�;�eQ�2��|pk3��0#��fVs7��+A^CXRFQoF�t�M=`YLfj��w;;	Q8�Q��&0`�1�cF�Wv��t��4q��d$g�m`7�Kx�ust��J�5H�X��Z]�3**�.��Pv9�Qu
�e@V�'s��H.�c"|�^RP����k�l��oA-�v�F���m �R9z�յ4�8,Z߭�(/���G�1�V슁ϖИ��Y�R��L����o-�}nS�]�,U9����0��3l���i�P3,/�ߵL}4���dۄ���B��r�6pƔ�HL9t��ҍ�!T9މP3%�K�]-S{ډ@bGm�I+6��#��{  d����W�����G�w���6V,8Ueޞ`U3��c�U�)��k�P�BO�l�3{���6��qV�2�C��nm����J�)
��pm)��AG�7�D#t��Bp��@䍼�z!ż/TWzǃ4#
��+�7*r�&�3L��\��e��X�s���5�k'9T(˻Ȏ���.��S/��"�1c�Q&I�g�?���x_n����v���%&S�`���p��^-��u/��v;;���n��\ڥhE6�����:t���,.&���#e��C�X��)���i�x՗f�>n!G�ݻ	ml�yZ;�BՊZ�Օmm]ii�1�љ�&\��k���PH�;����_�J@ �gϖCF���v�,���40�LVoo��ͤt��є�e�&�e7�o��ֱkvt��9J��!��u
%�#2L�j�Ṱl)�&<��80�@�T���ܒ������"[j*��.�Yb�,U��s��Y�/WP˭�Ő�h�s�J���5�e���5����1r���!���Վ�7�a��*FX�bI9�d�2�oj��=�S��S�5�:ڳ��ŝ�k$��&i���7Z�x���
�Ǜ����������ݕ���׶�8��3`�l�^����J�4��Xɻ���;F��4�U�N� B��c*=�t��g�C�|�4���K��ԥ�1
br�
��n�b7un�.�0�ь�Q��T�v5�h.�5��*.�	s����`��fU|�A(�\�At�'r�ՇM$:I�CulDF1�6����}y�b�N�:�d��Κ�*.۶�5�8�s������������__�3�������)ձ��N�j-�A���U�E�7U��{���E��h�m5፣M::4]�Z6���y�ǟ����?O���������s����tI������ۻ5m��E�UQ�;��0Gq���E7�4y�1�<���|_���~����>������?B��ml`kh���m�"��v,`��H�DAMSv�9��Ƹ�Qv�m��AAq�����:����y�&��k�GQQ�EV�[���Qq��F��b-d��=�/;�h�Gcو�������"���v��߽�%�8�"-t��F�mV1n��**(߶)�yۓc}�Ѻ����w��PLTߘ�h8"�6ēV7��*�����굧�ˊ��P�E�}m�Eu���*:���;����DQ�U4U֭f�+�b�����*��v�(���5�����؊�#���-�_6�F��~��N��b���+�.Ɲo/.�<�Z3QF��m��/|ѷ������.���L<p:xV�J�Sj4�Ω�ٕfܭb9L�Y��ө�VD�խʃy��U���'\��n����tÁqyݵwgxxۼ�b��� ��aP!�G��&�WQd±+Z����2S�/:��t��ނ�}8��ɥ�T/�����_׬Y{2��C�W�Z���]n�#�'ܭ�o<����R�O�p��d[�@�&E��"6�5Z�X�4�.�-]-�o:�?aQY ���Ϛs�3�D��C+~̏#8�k �rFwA�P¶)t�P��T�C�^Mn�<-�)�~(�J��)�"o]06�.`��8���҉����[�H�jӶ�fU����jƶ�c��������֒�G�:W�
!���dB{ab. ����.I���mN�z�c��7��ô]���(�mz%��tQ�wT:<ڢa�]����w�M�*� \\wv��\�:��qmB���5�^7�8��_�B�o46j�wtb���{s�Zr_x_j�j`��Ͻ�1E!�`JF	u/4�Ó�{�C(z9қ��$��yN653<�<��B73(ݨ�TwLoOC.�dt/�
�z��s��ߢ�ZW���ϯ��3ڞ~������S���g��r��Y����Ӱ��v= ��0�9�r�/	:Mx?=�1m��D���{����n�o�\I
�[xC�U��m�p{�7�Y�R�{�~��^x%J15��M��7���v2�>�y���N��#=gz�F�N]�v��;�g�Xע�l_�o�JM�vr�@<Y�-;"8�����{�>^�ߧ�>����AC�0��a2(�@U)U>�71gQyr���
���,v/]e܎G��E+HAu,׼�`2�YHh Ra�/ѭp9��w{���v�<�(��c��6�%�>�S�4�U�`�O.��x��y��>�,��<����׹��t]4z�>�L3����@v3	��F�
?��u(�v{�z{/�8�S�bt�X��紊@C�1��	���伋FE���A6��X,�9�`�鵌�Y~��Lh7ş��`�w����NdQ2��F�v���kdN���2[�:��{e�qFl��q|k�B�{���Z�[�΍�&� ��9C�^�,zCS���EPݧm�ήz9"��k3Q�lfw�;"����s����j+P���W��5�n!fr�r�g�lY���8�b6�d�'	��|�d��׶�A4=����5���G~�����/�S��׋-�P�'���9m�y��N��MLg*�c	�I�z�H	����}���s�vA��7`��g���5�A��Ϟ��q0�.���wI�ަ,g�K#<�4����/ �X9�%����٦/G8��Z��!P��s~��'!���/w$�އ�K5:wV8͎&�����nP� )�w�Щ
�K#�e����8���WZ�b��.��t�0�GNS&I]���P8�c�:-����`�����L�9eY�1"O�]��=�D_�ʡ
�
����  x��j���9:��sM��'��/��2�u���V�0��Ѓ<��3��=����!7��y5���$u�"��XS��a��M�����iD0ڏ)����Z�j��Ʌ{ws��_���g���Q���u�:4��,����y(�/��q��Vz�^��Rv�ʵL���
xd޺�7��̱v�a2�Ob��S�(2�O�W�(_Eg<*�f��d�pG'�3�S�����tS"c)�����M�@�>F)���Ǜ�	�b�{M�mO��D�l��c�h�����>���́.ʶ��ێE��g�f��ӝ�~gۤ�G.;n�$�F������+��H�[j�&��z�s���/}m?6U����7<���3�.�7(�J��	ev������Tp�R)�ҞoH��8+�G]ɷ�C���M!kQ͒r���N�-z&1�����<���j���#��l�~z����e�"�j�謵ͅ���/��!PaUCnP�^\ŘW��űq����n��0C�*S�n�_%��+>27�C��E��r,4ɽ����4Lco��)V���],���ڸ�˓�*^�v�-屯y�]�k����N�&���2��e6VKy�T4c)��y����7���>}v�ϫ��I���º),8D�!���xY�HɅ92�c|!)��&FP�{^M���uu���2���4q��(�W�ALZ��*%�Ons��V{���)������*������P�M
���r��`F���z�� CK�G��=례��%�y�
XG4��`ثU�T{�`����AgM�}7��������|���shCZ�[fM��i~pX�̍d���E���g��ߟ}�OA1��oi�nb4�^���//ʣ7�б���
)(�~�>����V�q�g�0ӂ�����	9�O�,eю�U���ν�mLԣ���'3.ɺW����
uB��M�A�Ă��P����}wU���c4�3�7!��{5q8�u��}P��P��1BS� �"1�D	��J3qS��Օ٥۶���?�P��1r��Sm^����d�~Eu�%]o~1 u�$ܣP6�����π�ڦ'4b�V۠K{�n��w�qU�1�+�pʹ��>z���E�ٵ�d�`b�M�
���ev$!�M��]�Vv���@hi��_���J|�΋�X<�¹�8��K�q̕X1�͗fS��N��ҭ`�R��!���y��Skfwh4ϯ�m*�3~��2�^J<��V�ƞ���{9�hL~�s����Ĳ�8 �mV��M�eN��h���z����|���EmBR�4q;�U3W*n�p� ^q�2-N#2uθ�>y>�wq�m��wyq�Q�(0�@h (@
 ���~�>���������?�Z��옖	0����\C�Gk�R�mߟ��Y����Ly\z�	i��%�{�����::o��vʊC;a:���)&c̀��Ue��\G1[�ߙ@�mNX"�<f�xd���6)�r�V=�u�i�ڝ�JB�΋?��Qѭ����=�!���5�κA�{�~�6Q}@��V_r.��0���2&�D��M@Y��n\�Me,���Њl��wfk��̎�	�`��2X��q��%��O��Ȫ��H�\�{-�'m�5����X�ǋW]N�����@Mo��#��5�h��q��4��d^�$�8�M)c����4���*��Lg�eAV�b �7���4$��V�0]+�W�^��"���N͂3�4그��;y����,6�>Ĥ6X�+p6��8�:|W���q���3�E懞�vZ�_�������K��	wgq]�%�ޕ��AU%���-�=s��GG���|]��0޽=�Q�_�M�~��.���:^g1po *ja��q���c�sF3IWA��^�UX�+�ŨJp���G�������P��c�B��*SM4/�ŰND����}���)s��랗I�q�s/�ù<d�T�վ�`�ɧ`Ī8�A�����-��j�v�M�vėgw6�3,3�+/w^SԞfJr��naɫDS�{���;�����<���?�!�A!��Pi)e�
B���7"��x��T]�Kո��o�j�}8�%���Ο7�[<\ݞjIuk�pb��X��q���%��D{��dUDZ�/��)�%
ކh!�=��}����z�wj��rݷ=�o���ԑ�jY2��tY᤬@r^���so'�a�Z�%65�nv�jВ�+j���鶡����܌@��qv�i�H��mT�m�ޘ�Q�����5�&���$$F�Y�*7!�ů5L���8ϑ7�V/^:��@Η�Q*�_����ij.x��J�S�v�MSn6J�fBE�ב��͋נ�2S�&)�?%�B���m��{�����@��]{���'��y��C�%�����\j�\o��=����r�_Ԧ��]<�A)Z�G44Ƒ�Q���z�Jv,4Eu��������*�sw=yOi@V�A�ԧY��z9�/A�`lJB��}��A�e��ťSk/c�A����Q�JЖf�X��B{`E�f��6a<eK�%�uĵ����[�zc=�7aF�8I����p�\.i�`$z��Ny�S��o>��C:�-�jiޮ�Y�D�z?b�/���"=�U󹓦�cx�e��Q�<^�מT̢��3���{G-S1�b�Ė�e��I��h��AK[���	�N	շˤ��Y�& ���%�cڞ�՜z4;����@0ʚP2�A�<=��` �M��K����+��ȫ0��4�ʊ��A��Li=����F��e��&�5�Wv�5��	E������C>���{'j��K���>� G�wU�F�����ye&/�,Gu�S�+�y��\C�Ry���p&�	�He�
�h�aD�;�7R�LU-�/��ER)ih�w��� ��"};+P���K�]"Tݾ��IƳo��׎��L�^�m<�)R�uj���
�C�	�����Cj¥R=�ʝ�=�a߇=Poe��e9���BE_k,�����G���^R	�l�!����g4|�l"a���V0��s��ŉcp����Yy��vh^�#W���cV��T�V:��0��ߥ�C2�1�!��_|��:1fJ1��Ǜ"2W���)��#��S'��,�ҭomy,�an���3.X��&�������!01^���{w��8���ջ�s�a��cx��\�SeQO��T^L�yN�Ow::�u<�4�4\��ks�����������!��H��_�K��6%r���oj�UŶ~+g:��1��x��w�Mv �Y3f��eC��3���^���cpd�G��G0�g��ӥ�����7	�6�4̃������7�f�Wz�#����N#�j�˥ZS@��L .'q�|�"��էG�������~~q����  ����G"�*�J R	O?~�ߺ;j�se�+�(�E�5���>n7~��NV8O7�Άj�X�����ӐA��N���"ʹ����Ơ3	�-�gf�f<����c����^��pՖT�������7����oH%.֜"4��G����]��ܠ�Ѻ�&�ֆ�~a�"i�S-��9�ƻ[l��Q�oL�U)�fCL&A�}(	���݇N5cyB�We0�_˭Æ�x��(�%���� �<l*Ƭ���y9⢵��T�P;���"�7^��tg�F��Q�"��c��v�3|���0�z��ؿ�B�rv��F��|��[�K�[�Q����\�#��~��R�����xC�"��t��8e��!�5j�Tu���CH���ހF:����qb����g����;�5¯�O/�[�Y͢�m����×-���v�Q;�j��W��d�ª$�f�Pkv�ɚ�CY��.j'��z�,��<�bt���LiʜL\?p4ŷ+'���Na��z�b�ȳۓ�y��:�2��N�Vt�^&_|�Z�K^���k	=G���%'�XR�Y���4��*��~g%����j��ᢝ,��y�=Ψ��Y֜�����*�+F?H|v��U�/�����;5F��:�����nͻcژ�9q��1n�Y�^���b��Si�1۲�7/��qڔᘄ���֕�u�ٕ,�a�R�q [q$�E��_χ�����
��/ŀZTF�{�y�Q���F]) �?zuEyT�{�b�6?�ĶPՔ���."9��L=��Cǭ��f����R�4�!h��B`n��@��[�� ũj��m�l�oy�Kb�ử�D>�+|�큖՜n�����z=Mj�ۡ�8�ގ�>p�/��=L����k�|��Sf.�P�ߍ]Φ�Z��2�2��h��2a��8��+�b1��u�g^�&�Q��՜m��3-��;X��j._6���7�����kY�Ny������q;�sm����@\bÞ�OݪG4*7C,u]b���V=;	�o�%�il=&��5�ŧ�x��wz6:m �-���zk�@nܞu��Z���܀���pm7��(��q���+{0}YՉ�ؕ�'�E��]�]�)�$`�(9��k�/&�ZH������ȅ��x�I;�KRQE��	��-ؠ:|]�~���"�^��c#[Sг��<����x�<���O�?:}~K C���VX��k��(�R�]3�y�n܋l���fQs꣗,ٖ0K�h�́�B���W���i�0�}(�»m2s}��+�.�Q�ë<㩲���y�i ��M�}�����n�b�`� ��J۹�%��s��A�>��r�flh�����q��~~~_���o�#� dC@%!�QWB) ���w��|~��_�~���.�~x�I\�j �d��*�"�D�uo��GF*��hJ}ktv�� r�PCoC�s�3E٨�1�\��J�����`�qG�.<�ǭH��.ҧ�Jw���޷�&}��m�x>�eH��fc��t���@p k6�zc�P�셛��E�ܩ���mO~���N�q�=�5� ���>�t��u��ͪ/!��OP�13i/��j�
"��%8.��4�w|1�Q�F�g.���A��I%��%�1Q�ky��?<��kVSc��%7~�(	P�f|_����M-�l�=�k�uHz�I>f�v[L�@���zὨv�nV���91 '�dmʓ.Vj��#�y?�����vҹJ"�I�sx�>k�n�n���\��[�4����zمc�.��oF�[L?�h��M����~�qξb�0#�̔�(�N���]��(s�\lw�N3��q�dWPN�mH��ӡ���Y�j��̕��z���~�Z�|��Ϻ�X�57��<=>����U�䁃<+�B����X�)d�|:�-v��k�h��I�hDx&�!n��������v��P4���-����f��Wm3R��σJ��N��WpԴ3̫�ݙha9�Y3]���ŗ�V��2kͤ*G'j"��Ī[�}9>�}c���Ƀ.r�B<�P��fb%��e:{�fh�zX>���'���7i|�;�ֽHnmg5�"�FfH�Nr�;mF���!����������`�yǚ�Y|8�J�褍i� �ֹչj��lyu7f�� �b���5b�VĲ��{Vַ�Z�W�������P\��at���9�)�����:]h���;�P��4�TU|1��J���۵s>0�3sL���J����G�e°i�V�ǁՃ�>W�TO�Z�(��V��:�x'6s0�29�p�c�ș�+|&�.[�֛;3�ƍv�s븰gV
�0��ͫIAܖŪmm
�짾8�=Z+{*��v���;bf���<�[�,u��c����k���	�O3W �PY��\	�N��c�ʂ���[,:W����>O;,^��
��95�F�I�,Co{/v%_R5��m���aM�=�h;���S�
��P��&�qb��_N�Nó���W
�s�� �sRT��X�����k�㩇�υ͗�G4q��vVb�;C�QL9M�m�\���d?<)C��*�L/2��@��%�KGM�������JـQ;�Y��4��*��)���Ի������\w��r�yV�
2��8��"����}�`ٽ�nG�@�ǅ��9�G�噦]>�[%I3*^���)9�'����
Y����2p��e��wv%�6�6b��z�Ro��Y�^�'6�a������Z�v*my��-�p�����j����0[u��w�&��G7��f敽ܰ�
mn�F}ǝ<7J't4�*��ɓkY���t e�r��L�!Q:���F��,;s2��5;K%H�bm:u'��r�p	 ��Y������l6|2󞼲�.3�Ţ�RB��[�pޱ��6j��R�J�	��Ƅ��x(F�I�fm��.���[%�iE�ء�2�g)�)�:�S���\?1X9�b����Q+�6ń-� n��ŀ�Nt�%�힣����Bk���p�q�7��e�Ա΢'�cD�[ͨU��>]l,Ks]<�wM�:�J}2�&b���5j�vL�2���s���z�d(��4ȃ�Qp{.aU���N�&��45l6E�k�wn�&o��0T��c
�vĺ�Ume��u�g_=�QE��5Vx��%W̬��^�wzf𛛋\���d{f\{sZ63o{�?��>n�`���M����[�q։�6ӣNƂ����u����q�כ�<���|}~ߧ��~�����������f"���
�pj)�]�[�1��X�F��*���<�q;��ɿ{lh�#��g<�~>?����~����?����9�}=�u_�c���kQE�S�QG]q�;h����IZq����Q�[��<�~?�����?O����������ډ��3�-���O�JQ߸;�"��~ƺs�f�H�ի�������۶;i�J��cUGY�"��QlP�(����k`1N�Ѫ
#���v�EU���Uњ�wwS7��N*��0USy��|Y�Z�m��͏KCu��;i�`���Z�w��m���]�h�kh�Zƈv�Z�.۸�bi��um|��F�Z�TU:,�6M֫c���v7b(�hذwn��|�^O��"j�;X�P���Um�Ѧ���bݎ��S����
�F�J:݃�~�>��k7�.��8cp��o)�)DZ���{��N�C����f��Ӹf��l#Hǭ7�k�ftب���r��������*C ����Gt����ߞ/��=K���g��;f�
��^�Ԁ�Rb�My���V��Q�:,�j�6c�b���Yb�>"���y���;5��r�}\�EV���πC�t�r�}ix��z����l/y��g�"uA�µ�RA%�5&Іf��9/�dO{T�p�2��Y�e4���]�]��ۈT���u�{05㦿��s^�wk�;9ꗞۇ��ײ�V�s���%�E��$П�������H����-�%j�A����h�`<h����UC��׸W<SV�����W���M!�	q]�~/��m�^4A�u�#�3���źrKs�[�d��p^
*3^��
M�-N4�EA������4���|=���Kɫ�57��,���)�͛%:~��D��kW�v��`��m�i�o�k�"�6��.�����Y=��L�8��������(�=��F�w�q_��U�vѹ�9u<��95Gw���ڷ��g�ÿ�@�zH'��d�m ��9\`�K{��#:s��$��X�H��;�eN�ˈ�,_=֭��-j0��]���ҁb� fQ����}��^[��fj�co]߁�hj��NS�Ĵ\a�-�-J�s0�x.�ȩ+i�]x�(D�&��x����Ͽ���O�O�0���V�) JQB~o>�������_�a�):�[ƂnU-��8�d_���fit��	I^��_<d��nm�6.�j�My&7��Z�6��kFGM5�,�׎D��	V���Y�.��<8-٣ˢ��Y[�����7�{˫<;�Z�)���a�J�U��S-n:<1w�����L���\��m��Vְ�
�ɁQ�Q�N�$꼱ќ�[�:L�C��Т�̀�n8v�C�!H�[����'�n%V�(��T���f���i�x�+n���i�rcJ��̈���nP>�S���B��79���f�:�0�x�ɺ�KL�b�}d3T�7��R禵P��������{呬q=&2�χɫ,�>3��WV�j��!{R����-�27^���N�5�V�����x�rC>͠ۦҳ�i�N��ʄ�h��[��]�(�Sa��{Qt�M��ZP�NS��:ȼJ���nSn�/:塡��ј�`Ms��o�j<�8�{.3L�'��b��ߺ=࣎Κ�͞�ǂ�p��ژ�V)G,�L8��[O*�oA�r+��nZu��Z��7P�pI0� i�q���bm�<XU��ŵ�\�O��z��5�a�>3�;�zȷ9�`Ѷw�ʒ�<%�s�<̯��ɹ�s�SUd!���.x8�w�f����7���+p�з�X|�15k��Ѥ��i�k{x+�m1��n�b<���]��w��ym����,0+���#@�(P*H��(���TC��
���,�k4Q7ŕ��Ј�$M�XDU��<㚵@����8��$�hųf������4?;r�=5�#�<E�i��<JH�ߓly�,���t;y��5�)�ʨX���{e7l]�wc���s��<�[�$�Πvr�N��*��Ng�����1�wV�)W5B��-��7mױ�K +0I��gڸn�#N��r����q�*\�m0�}Ġ����4L]�X�MG��)��3��1�➙����=�[.³T	ʘ�zǂ����/ܱ�lVA,�̍�4��`�uR��x�1i7ɱ�lԗ���[X35���<�RZĨw���������/G�L*���P-�����+�Ιw�/�b��о����'[X�hpK�=��ǑT��忖�)-�¼)`-���C�W6r�z�+hqQ����~��w��
[���ג�ĝT�kˈ�1�r�2�ӅIY��ZǕ��P�4��]�Z���/�Lc�A�L����[�����i
�P�5u��=�#!�e�~}ֹ��ׯ�'Ք嘣��N�i���>5Lc:���ヹ�	+*��co�\)����dGV;pNtS����]�I��N�����)}$�T:ju�/:fp܎�bm��hZ`�u�;e&+N�Y��Y$����5���������]��}��q�����eQ���(y������.��47�/^�M@]d�_�R���y��1�m�;b������q�F�,��NQ�6K,uު�)�Q�6��(�`���@ʹ,�#�n�!hEW�:k�� �vj˴��S����`-�b�C�19m]�+-�5�"����j��$�W-����{�f#qO4�Tu�~���@��3k��1���pb�9�����Kߟ�y���9.*�͕�a�*ɚ���y}�^���=�m<H8I&��Q�FE�>�X�o䔞!��C��8��@�~J�镑 �O��L��bc^��i��L��ŋ�v�Y|�Ft�������իw<�z��^
�v@���yC��Q����H.7���֒�@��_Bae٭�h.D ۓ��끜�|�7�z& ��3(��@8��Ư�i�{�h^�iJm�Q�w� �:j�}tyy��yLQv�=�R�n-��ȹU�X��������'z�~�mv�l�{lz��<�%�n�G��0j��-���l2*�,�
�G�^���P��אC(s4�^�񿽽��NOm1I��vQ���f^�l_��`q�:e2�)R�+Mt2��<"��<.Iy�#��MZ��l8��)"q�0�:.�XK�3�>WB��]ju!I�We��X�i$��+c����ҥK���!�e�1�~��������������U��!�)a�jFE�	�H�_���������~�����k���ؽ�:�榯a|����r��"2��u/:lq�Dz+��C8f�]���5^NN�:Ɩ^�	���{���j�^?�b�]������������f��b��8�nf��ڼ�[Zv:D�钟l�&x��Etؽz3(Q�Br����[==���1�w�����l�u`85�ӊ�����1L��(���u��M�F�{�=�v�FqR�fьN��4K�+�E�r[�9h��p�^��2Nj�-����q�1.j|��m�5d^NIה;��Ԙ�Qj��tŶ�m�N0�M��P"����j�!K���8��S�Xx��t�L_��8�i6p�j|��Q,y��f�y�<�˩�TL����k�΃�X2�]��Y��d9)�zS���q\�>��ͳ�Iؾ�@���fb��/��Q*iV�L�{4N�k�X��9��	V4�m@�*	�����[��z酖5�xQ�Tj����=��嘻�#�g�$/�4s�8�_ù�V'�Z9�UW���	�.�lo��&��Ԗ~�k�	ԯ�͸�f*ˈ��w�W�	4��˺j����"��6��R0��ѓϥ��9�o=������>��uKC�;��7s�6�DCK.)�d=�:���w(��
����H���ss�A2e� XN
yӼ������ C �"�� R�B�#B�^�>�;������������O�^@��!5�Qɩ��]�a29U���9�	(�tt~q-	�д�R��f�1�~�w��aB�۱@�i���HOp_mr���Y.���/��Y
�SM x@�i ���gɹK�8
�X3�Q��T�j{��r���5��qB���%���ۅv��?'��ǚFj����/?{��dT��N�~4`v����E[��bS��WS޵&�3���oū5�݇*�}e��K�'�)1�%5��my�-s:ˇ�`��@Ę�����k@i��,\�ϥl�Q��
ʑ=t��Q7�`�`l"�#:,u��*�����!θ@�-kc��x��	�hJ��z��)���a�It���f�U3K6��YFL�n(>���l-�F~��js���%�*�7wi�sr����x��[:ƀ�6�W%��izI����X�My���_7b{�o'�����&��~�_�a_�{%��מby�&���2 -�oe��F�v�?i!�������@UJ�� x$�Rs8��)�U��6og��0�Y*b;�p�Ҫکk�!����\�7Y����g�='���4�%e^�(�ev���sUq؍�u��T�Ź�K�ucl�����Y����@��E`�!�`��	�o�����P�!��Q(I
�R�;������>����?�=���6�\��\��Ur{u�J�J�s��S�����z�@W�C��&x��H��<Nuv�6��j��2b�^Ȗ��ͣ��74o6�j	�K���|j�0&���k�/*�m�����=�N�-�q�i���օ�)��������^�[��{��<�ѧ���B���1�<�Yp��v�t��Z�/�<�����u�]��i݁p����YF抓��iwT9K�{4�"i����o]�ժ*:�ցD@�0�M�u�ICY�}�n���h�˿+ފt?��@��z؋E2&��u���E���a���&��nI��;滝�Ǳ�׀T�M���\�%��"��8ep��C��xl�3�xi�	��Q���T�ӵOնS�hk�#��
��6�2�1����Mӧ�fա��uό�~ɣi����]P��uu��Zdw����U)�>aR���^�v/�3k�<5�Y~��8��6"��t�#bŽ�iS��~h�7�쪁&�;��a�x7x��̢i�1��9M��ϩ�r��B����	�=uc�3�ݟ{Іυ_#����P2����cJ��D������nti#!�z������V��Nѣ�R?Q���*�ϟ(�n��Y곚a��<��u��-3z؜�u��AsZ�����r�n�1��}�֏~���^�HE�*a�
S��������������~�N���� s�Rdt�%����s,u�5s�ǡ�	�9��qݽj���%�uhȧ�/щ=�o��QHu�<������y����H�؃�J�oG53b�,(�_�8��ʾ� K�R���mP�
\����o�kXs��s����l#
�K�d�m)���L
��ۏ&�*C4]��\�Ã<�)>�R5�Y�@�l*h��XQ�3������k���� �hބc�ٮ3��`�Q�F3���>H��nf���ʼwhCuå#F���qQ�o_�s-u�^����Z�M^>1���M�`�&�t�9�LL�'��w���z��4�
Xu�jH0�*�5�_c5Pt��S��+�́2T_��*'*$:��~�{,܋^��)���0�x���W��$.�����3z��c�DD�GL���r����[�@bT1��H��U�K߅�,���M1W��p���6���Rբ ze�����^�A�QfGs�|�>��o���a�{��V{9�X���`A���w����q�ѧ]`~`s܃��J[{�u���I��j��G+5��lX[��XR%}�3-npR�QU���-�0J�|�M	:�����{"X�m���]�49����YK�
k�vqjs��<���~������v����>�?� �F)+�U�M)J R������~������C�K�lcNͶ�᝞�N�N�Xǋ.{�>*��1{gNZ����DҎ^\�I��4	����� �v��8��K=僾K�&�%�څ��i����Y.7���e�l�+7���E���	6� #b��XP"�`��!=��q��2��+ ����m���0ms!mCn)%f���|�P ����C��f|���>�w錫�R�u=4���+y���o���q98u�v����|��
k���]W{��o��I�z�B_�?�������ǶY#Ոm�vodB�8���C��,˟�}�m���F[��Z�nVl;#^h��{��@�����6ڞp�lK��B���8�z�9r����CaH�)�BF��͡Z��Яr��z��za��E�e�)Ov�u��@�F�,!17�h���v؎O�:f�:tM����%��f��׽���0R�If�L'�RY�Ǖ�s����7���m��Sf9��5+�{���}"Kj~��Oy����{����'!� �-BC�mL��^�=F1/"}���|��@�H"���۫�UC_y�;F�N~��5ϭ�l��2Ӝ�M೶.�����q(JS�ec�r�j5>�$Pd��pi�y[��}�^h����w|̙�ۮD�$�x�:8)�B�oJ�ҎRbo�K�A���T�s6^
���?%�
�!�R�oy�� 3�y�T�]Ƣ��ܺK%�g����:qrD��������ޡpS��{P-5"K�ܪ'/i\��1�L659O���%%���V�,��qa��	`��Q
��V歘�ͬ���X�mC6�a�EuJ�Ny�c����E�'�gb� =I45���1�s�3�Pr�+��m��?'���FہSp\a�����Ir��E¦�K�wPy��Cv���r�>b���©1sG��c��ժf�t!�]�@�0�	vK�°z}�5�~�m�c<���{�dY/�fz�^�Y����?0�g��o��ߘv%G�bb�嘎 ���̞/�s4�k�<d;a�m1U+�p�@���1�G�i�X�Z%�-�&%�������cG���3�1���L~$D[w���ߞ����>|y��~cۥ�8�yH'�D=����HL�pU54�.;<���o4�'fe+�h�H�A�ns�&�7x�s^<��,0
�a�wM���)2S�qT2q^�('4��QD1~�s��44����v[�u��|U�aN��B y�T�]X�w��e�}R �.��)m�o0f�\]�'s�;J�T����#u�7C�7��k�U���,�|�b�֖�ij8/�)���)�ů'\<�r�& ��xV�X����e=9Х��bX�I�K��yk����B�T�M8�2^kv��v-�A"��]���FZ��Y\;*�ӎ��gs�Pn⫒�F	n"��G�㵊�\�o��΅��X�s�v�X�ov��ɖuE�U^;�+;5]5�`��W�%N��Nۭ��s�o9p�ږ�b��:m��MѮ2�pM ՗�2Z�X5��r�8�ٔ0�e��Ź����_Gs��S-vev۷$�6<�Uz��D^$S!3{��1U�n��
���Wm�p,��ھ�wl5����*f�m�L>�#��P2�1zVU�H��c!�U� rT�v4r|t�(�ԣ�̿�,x	�0�5;�:�e�똴z��n�����	E��d}@�H�ܻ��q������X��h�j^��U�����6���8T�����V*������@����
�gn�,8X����S�R\�^t�%�X�fN
�h�3}-�҆!u6�J2r��V�ט�����I�7\$�����|��?7�I��X-�K�ʤ���� (����;��Im�����I�8���J�]8�Bu��s0�xP�(� ��B�[���nP�:&VkwJk�x_r׮IQ�n?�k4,X�B�pT���hf�^`���]�F�N��uT�`��%����ct/;��a�S�AŐ���Z�ީ{ǈ�{"��h��Q��a�ݻ���.i��G!�n����!D�y7bW���_^��Z�$�%/�sY9�:��ɱ�,.ٚՌb����d=���.b	�a�$�N8i�	��
����W�t�o/��/��粐�;�G�C��wv֐��R:��֍�|*R���['�`��龵F�{U%��l:2�f�q�<������y>��ǁ���t�7W,O3xH�]�����ː�)���[#�[��oo��^�����Z�:T)�k�2 C.�N�Z���,�S�B�����PD������2�t���2���ѹ�}P��JMw�&�ݷ���˻�+�u]��%�M�7�l#ww���I��'+Vی�\�cv!خ+�6�vj���a���;�m��v��Ĵ�0N\��k,&,H����lJ��W�b�ә�)�M��uҷ����a4�2R ���� ��a���H>��v����q�[�A����g�!I��SS9���F<\e�+U�]��&M�����J�	lr�Y]ʃ`���a�^B�Ա�����{+HL􊷍�G��q��fS����W�t� ��!���]�E�o!���xE��(Ê�e�wI�� �FZr\_�0� ����Ln&1��(�$?Q�����q!&	JBdL�7v�'���B	I�dUy��}O�t]���P\&�����h>N�*�S��=޼�Ϗ���~?���~����Y�s?���~�K[w���|M�t4QQ��E�����訪-�b��c>9�>?�����?O���?������}���"/�Um��+Q�**�ulk�f�K�������������~��������3��������cF����Zdv�V�j'F�ڮ�6�q\WMwj.�5h톊"-�3;f&���*b6gZOmvj5��Th֎�3�;b�ꣾ��[F*�|����d�מ=SRl�)��ր��:�"��O���{�,[Q��u3F�����F���δQ��ii[�5]Vi�
�`��֎���v��(�6�D�(���TcL\Tւ���|�9����QZ�m&8�D߻�V�b��Ѫf�&����	��H�H$�p8�u��273<�Fѭ��-ֳ]�QwqS+N�ׁ$7��Rѻ'RM�WGR�Qu)�]sXķ��������l��iH�I_&�CIE$�$9�7�S��Δ�+���)A�(�����}�_���*��2&%}P����Q>�b~[������{{��b�Nk+#1C��UPاv{�g�D�`���[r3װ�\ǝ��0�q̱�7v��Z�!ޝ�`o�s׈�l�ل��uM��ʭ��N6��m����
4y��N��u���	a�s �b����Ov�+�[��wD�8�/l�F Ñ�����CX>�q8�-�t�76|cjq�����꧲/8�ǞF8w>��Ű�lE�1� N'�V1���5F7�b�sR@�dm�ԭv�|�k�e�����
��:������ϡ�Ӊ��r��y��+̥E�ܶ0B�X�#+�3f֔�z.�QL�����C�w�Ȟ��v(���Nl�jǃ���SYn����!���;i��*7M��l���҈4uS`p�k�q��P�Z�Ҁ�����#��fg�ф��;=C�Q�ܢ��l���%
TB�4$����lG�n��K��x���o��<�C����F����H�m�x�9M��s�yt���1d6 ����6���a���y��<��aȰE���]���Ѷa%��h�`=�����f���g%�[*��[�3c��3�N@O�ʾ���Wͪ��x����ق��8��ݵ����s��З��r�H9N����2�7@i!�]v�[�Ϟ'�]Wz�R �~�7�T�	ҘdHa\ �{��3,�Rp��,w�/��d�|�x�@��i��o'#y됅��N������I�sCS��iu"����vo*<;Y��-���q�H�����������S@rj]>�6+�kbeC�Ǧ��լ�m
] ��b��5�����-�16#}�3R8���4��LӚY/q����l~1M�DT<�.���T�X�^�H��z����X��o��N�~_��t��e^�ρ���L5�u(�V՗�j�_\�e�$�� w�Je8[/0!��]4
[#�s�Ǭ��C��닥M8�5s���~�t����0�ؒ��&��Ȱ��(�Ao!��d��������˦L��"þ���{���-�4H�,�&\P2ek�*4�B�ۡy^YQ�)-�/N�מ��5{��{���w��	X��)�θ®�Kzm�,+y�Ǖ��F@�1I�u�O������ۮ:̽e�`��\���Dq	[�܄�z���c��2}`�{�طJ�v6�F�%�l.���������ݮ�[hgxv�'#K���n*�����m@����z�)�$`�{�$nk��S�uavk��w]�Z�m7�{{w�v3�r8�}	���������+o�:���|*��|g��L۬3�5�������Ӑ�V�3�L�6�^�b�'�hN�=j�:��݌�R&7�:a�����Y!κ!�ʛ|�����pɔ�
���������"�҆��|�F0��׊<��.�0���#����*�'��Ԯ0���n�����G��������S緟_�}g�M}��;�둿8����/�_�aN9TPǤ�x*��S,���p��΂�'iuc�3MV��b�������M�R/�\�k*�i�����j��	��xǗgH�m7)0�BJ/�S����<�7����o�&+����찄�|���ݪ>�I�Y��� <��_�Gp�>��|o7���s<��!@��>�J
嗗5����<V�Nܬ�Ηt��Q`��3�=���sU=�H_Rp��~��|�~^'������V���U��q����yJ��w�l�oK�ш
S ��S?EV�����/��}��B�͓���(���y��ߵ|w��9���"�(�OL��û;5���:ށQ�j�a�ӈP� �=t��4V�R��F�ۃv:8��mK$M���C?dm�\�}��#:��������NM��5�x{*��x�M�����OL��s�@�,���R}�9Ci)�qn�)�o�VY���x>Չ�z\<�4��ڃ@��y����Ee�Q��'[[��7�V�a�L�M�	�דz��R�Z��1Rg\J��koj�҈ަ-lZ�ue�������_m[�����%Kۙ�#-�-��GwI��c�j��_�/�d>����(���Cs^����~�����%�����P0lI��0�Д�dL�X3��2�G*������]a*5�e�U��COy`�.�gnO�2`3F(:��
��\{����e�	[��TZg�׼¸;��œc,������W��9�jHɿO���y�ȼہ�|`>�&��R[���K���a��ܚ��-R[��Z⼦9��j�Z5���6�������U9xH��')PA�n�ٍ��V��!��sH����rZ�C���1��`�I-ȵ:gmqfO���C�:ritb�Ύ��&���="oc��^D\T��ي	Z��j&��a�� �qy{�&��隫hx5�qЙ�/�#'�؊�z\�Ud�~�P�(�(��؀mD7��%�]�Mܲ �]��c��ܲ2�F��K�B�P<�aAc��v����O�L�_��ی������|�t�E�Yj���̭:݂	�7ɘ��AaY�/��5�g(k����>�=��1T��&��;(Ual�>D��l�7�)�������s� ֻ�4�	�E =�m�.y���]$h?�Ư?M�1&f��[(o]ܰk�kN̲{�C����NT�yd�m���f��}��n�W-�_��ѹL1���+��[&�\�2���ې�+���9���:�qz�9R�a����Bd=!�B�o���_:;��#�6�7qmn�.����$?�)�2����J@�I{}����&W#��`�n�f��~U�m���2��`��Dy�!?��tj�	3�|D�E@�5r�a�{��S ky�{ҕ����8� 䖁�����76]���P)xr���w2������c��p�8��+����o,o��0j�$�W	�
)e���ݑ>�s��b��+#e��Ck%𐟂��^W� 8���,>�SMCqK�r%�ߒ�omx��� �E�4X�V�&0�U]���uԉ��J�@�����N| �=�>�9�O���y�k�h��T�ڶ�4��9�(�e�Q�G1rko�N��t\d
��:���i�A��q�S�K���7Ѯ��bެ<T�QJq���5<�`q�l9�IoL�e����}��7�S-�醮��Ϯ�<P9��g)�/���qA���s�ZҎn���~�ʠ3q=~l�����xx��^�yr�u����-�e���7��4"�U��Ds.��~&�棆=�f�/.߹3��h�l����_�F�]�,��0�!6���m��IǶ{<��p�Dҍm; ��R�{�5�����/�r����C�����y��u�{���D
�*{�|��R�{ٷhԆhk��H���j�v��y�-9�7Ȓ���%ލJ�a�A�`8K�2�����mP�m��j�v����>Nܨ{� �>? C'��C@0������ۘ!���0�Ms�n�-��4T�9�FFz�
9^�~�'!�	D������]��N�E0*=L�Kx)�	��w3Xk{�6���^�;�K9N���VFg,�fz��@`�σ���=N�����d��L���v�� �[���J0>���(=�u����2 ���ߗ��gzJ�7`�&��z�'��-��|*4#XL�����m��	����7t<�d���q �_���X��8�7.�V4$��'*_Iζ4Y}~�v5h��ލeY���O��]ônG��N�n.��o!��O�7*:e�QN��Oi����"uZ@�f?ɉ��(�o7���ȸ�t�"�a�O�S6�b[*\�89=��-۩��mN^�;�Q/�OT%qB��U/詈�o���>wP�څ�ŧ hjfnm�}KfUq,y�ֹ��[TڎH��n����A�=��p/���*�ֶ7���0f��E��nu����e:��M�����R)����S;�d/ S#��6��8�/��ܿ���/ҡ�ݎ���aj�M�y{ч����`Rg����v�j�?g�V_��t��5Ku����6��D���������7D3�@����{x���,Y�8(қ�U�Q�s���9#.5yq��4�٘���NWV�kn���jL���ϯ{�پ��_>�<?���a��,�7�x .�r"�"�ߔk���G���ڷI�gT/+֫kW,��:�j � �7���ڊ36���&��uR�f;�Q�a�#�1I�p%C�Y�j7I���l~�j�����%u���g���ݩ�����ǌf257�3����(0�_oN��D>\�A�O�:�fvNE���qp�:�L'�C
i��ס�r�5�6B�v٢x��pE$�]����ɼ��;�V��f�쐝���nm���pk0���޸��m�7C��Y��M���Ih��:������^p0#Jߜ��\�/�<�K	q��r<�_L�1����cZ8�L�0S��z��Ή���ZI�`�Z�C�� H�`V��w/tj�R�}� �.���#Kt ���Rq����^��1�{ �s����mI^B����W"w���Ԟ+v��W����aT���³�p�i��=����_|L@*��fOEݑ���ت��[��RY+�L,��t	�G�;�ꤌ�-�_����N%�%�)��o0�,X_
V)[��N�:���3"�'�1;��;��	�Q�:b��I�y�m^7��ԯ��n}�7��̖�2���*�̱O��*���	u9]���n��R�p�*�6��n��d��#���x�ߟ�~����������$0C��%�]،DFc'�o����3n�G�=|��V�T��:��0�"�ݰw����Al�.����;s��cu�1��p�_=$��� �;��k���������V}d�USc��;�m��sw����faJ�%Q��/cC(z!4�K(NJ��Ed1~�H�sDm�0K���+�{V�
#n���tby��𚚀܄�|/)��8�]� ��qv�;	��G�./���k��t�v�YG�:[E)� ���=�)>�J[�7�����f 2�H��E����{.��oja�Ծ�Z����N$?�9�9��N�8��sk��휜n�ō�o]��A��d)�O9�
�����.�݃G��0�� �1��),in6�t�G��(��	�;u���;�3��b�ηs���mJ8��'�A�t<y�G�����gMơ�q�zǒ��� pn�����=��t���$̝k�ڭa`dӥ[��$-����H�$r�X�٭Xl�<f��mOCuj��6!Q�z�XO���:y��2��Hp:̽��bV=��|�4]�Dm�������3o����l0�Y�60^\����yj�SOl�	�f>���`��&訫/q����¸(�ҕ��"��X*a~+��]ƴ�yWI�0�`vBu6>��Z*u��4S#Z��xc�׹$��N�<�[;P�Dσ��ؔ��3x0dH��-��L�	e|�����e!��Oa`���;��Mg#|�$�ݤ�'M��ݫTJ%�<�?O���C=��߭;��ܨ�^V⪲$���=Ջ�5��G�8M��m!�fr<%��p��\*��#ٌڡ�g��~�Io+����2��SXXv���lR=C22��Lp��H�l�)!�)9<�h[0�B+fK���w9ɶ����BIYkχ�˔�֘�[ަ��G=�ky]#K=*����r�ʦ6q���q���R�y�m{���O*�kIr�J��fr�sE� >���f灚��JM�ӵn�r���w!ϓ嶞eM��n�F�� ���{vF�<��
��R�~�n�����G���C����w�H���xů[�I�MЬ{��g���3�v�޾�Se_Y[�Γ�JM�����9��9Ļ��d��6Ѻe��9�R�ofXm=�Ű�ԄLU���H�||Ɛ��<���y��װ�K�f=��[o��^ӂ�`��3��2�i�.͙K��Ywc0�s��-����Θ�#y����4Z9"� �I;������������jBA07/������O�i�c���*�Q��rұZs(�Z��2�18a섫t(7�t���˾�B����-f0�iH����B�[{03ʲ�0}Y/�4b��k`�v@�:m��3�^�eJk����Cb��D�d'��E�{W�2�C+����Ͽ����ϛ�Vc��%����8��bTKaW~�l�3m��4���]#��!7D���5��fGIz�!L�U!�����{b��$���J�氪4�+��Ĕ٬����N�ծTF-�Xx	 E9�I��k�	f�Њ%W'�̺���F�����_��a���T�؅'�b���ꗎ!���o��	�_�=q�E!���y����
�}cL�C����yġ��3�a`��p����R>.,X�yPv���6P�hR� ��=��&wSn�;m��0��`�^H�F�3
&����֚tq�<���^u�M]��\�D�[�n�e�\��Q^��
�
���r���&�8���Dg�1B�<����H?�2�ټ�]m�J��L�i�1��;�}z{�����y����-xA��423�E�E��s�XӼ��ia��[3Y�3+���;~�$H"J�.�:|�N�������{�]o�m��M���Ns�gi9�)���	D�u�}����rE���	 ;���٫��O2���M�/�{�Y\]Y�R��s���X�D��A0;�%>�j�ړ+���7c#\Žk֫W3.<l�+5Q�Z�"�	\�-��Gޛl_��f�J���r�S�� �Dy�Vަ*F�:���"��$D����W5�6�F �Wu	�9n�/:;��^���R�tD�-�M��*�ѻV:U�T�X:�a��ꕇm�j�k��+�9�}p,���Zw@�D�p�a$����0T}e�:ֲL�U��f�׉�k�WGB�Է�-m��!�F£ѵ��y�������V�N�:��-�|0N��H	�j �	���v�p��d��O�ޚl�V���\�[��Q�0�u$Zԉ�ɯ5,#5n�����q�w�[�cA�/���s��Y&t�`k�\��{�0�N�h5*�j�j���;��Y����u�Qa�������{!�̤/y�U�elI���NVaC݋��GL��k�V�6޹�x<2Tq>�M�&۳�[M^�s&] +�Ҝ�٥�[��C z���x��/pf��3kmoaǛN@����Z��k�0�&�	���\��K�ჶ[l"\�Оm�����P3y\r*
�6�T������d�t�W��z�խ�,��ٱ9��s��b�����g4,�����hy�eM}ԓ��Y���
���!H�G���Iכw���|v1Pa��ڍˮ��d�gtc�y4�zS�hsklyi��	�WC��ȃ2KF��Gm�c&Ik��N�x37^�[������/���|�
�dl��v��_l�;eY31lc�Mc��
.�=��F�ֲ�jt��@��x@��&;c)D�&�E2ujrc�oi��R53,�Do�؞>J�>���q��ֱ\.mf`A#x�t��N��3�s;�V-�J � �#��WuˆU�X ��{D�b���\�o]�l^�%Z���ZI�枅��^.�����LN\% �U�Z���
m��g!����q���/T}Ǚ4�Xힸ�z�Ad= &�0�����cN�J}�9�Ǘ��K/3�l�D�Le�u��4ju7�h�yy�Wmf7X�mc�C@fQ���]	B�MHi��rJ:���#M��u��V�R�2F��MeWjǚ���#���!G��i�іU>̵�/W:�n�Z�J��MN�[���!j�d�w/Q����\+���C�TqD�ͭ�o�*]w�7Ul���䆈'���<���!�wսB[�0C�M�k2�}��\�)�}5n]�)ˇ�	rP뷐���P@4�Mksx�6:N�"ʛhP�d`MnJni��Xh�/� �j�E2Ve�Yݒ�b�Joj<��g0a�ss[�b��p��>   �Oգl�E��]�F�Q�ѷ]�0Z�1=�M�b�c5W�9���?������O�����3�?o��_����\Y�Iō�E����l�N�U� ������<���������~���_�g�~��]zGGF���]��3��,�l�i�<��塣�<����>>>?�����~ߧ������~��٨�b ��{�f�����TQ�ţS���QI�e+Dm���)h�N�y٭�����&�Z�(���GE�Q�cy�����ֻlCk$GY�{`���(���S��i�ƪ�:���u��F�]�������5S�<� 8*j�6�V�EQ@kTw���(<������֊�,�tז��ɼ��"1y/�j<�MW=�Fѯ1�NM�Tv��b�j�8����4�Q@h�v�4kM'�%�wd�c^]S ��H�>��w9��8z�U���d1����f2��\͡#"#���-.��ϿϿʽ����~�����Hb0 �#�w�>\�s?����񢝿�<7���("�}�|_�
$�����nw�7(څO��3^+em�)�O�E�pr���l5d���L�g*1�P_�un��b�D_Dd1���:�]�6b�ŉ1�3�޸��ⲅU�����Z1.�d�ܰ��:pc����Ǿ���b���'^2y�?��u��z:~^+����o���g������#Y����A��=A��ϳ3A���xQT��PdK�9¹�\ �)�j�"�Z�`�^����p,Fǝ
��P�+���g\㨎���kY[�`'��d���ZS�/%C�|��¼��f���^�ѝ�\��9�l����Sx،�v��#GL.rްb<�F�6Fd��Ɨ����_���D��3�^g�.��pRo�V�w\si���X�R���|�C	a�Κ.}�(��s�^��1d5,���SmIe@�\�C��׊ӔZ$���~n��>}���r�S�ʂ)%)�PY kAz��>l�y��a����T�y#x9�--��%�L��a��ݷ}���� ������5�P>�;lŴ�ȣ�ƻ�LR8����z�V\���6�ߣީ�fS�'k6;���t���Lt�����zN�r����!�f�r��FoX洦�'AE��t��Oh��� �hKￃ����G��<���` F3.�����='��"|7`�����9Ҽ�ʧ�|�+��"�I���;"5m+�z��d�1�-�vk�\�m��ݖdc NP���y�f�J�<�Gȶ�__�?4��?�]R�	W�s2pA�J(�9~	��H����u8p��R��ɮ7�� ��x��8��.����z:*��kV#&������%R�N��Bɮ`��$g�!"f,�*���/rوJ/��b�^�HS����D�������uF3H�W�z&q�c��F�yא�dH��Խ[�j��z�tr�a�*6vWf���,�J�n��3zHn������$��'�>�eKc�ަ �8�{5	��wG����y��Z�r�qX�n��2�8�R��5V����&Y�ReQ���/�j�!����y�{��s������%t��jO׋(iJs^��v�TNQVm�TSX�ݛ���� X>�Rd2�A�Q�,�)N����UT(tBO����b��]�8�}fD\��!j�%���4������2>=�$4z�h�]�#�ɮm{����0�sD���,�wS�<����<��#a����=�����Q��ѿ���ͬe�OA��Y]Y��Ko�8h%�_0����)�.��dg���.��Zȴ�W��jR�z܃K����L]uo5=AC>����wj�����s�Wպ#�]�9�eR%%D(!~������mEIK*����}3��7����?�g�?���/����w�6����ʅ��bac3^.'��E:�� �w���(Z	/��"Ґ�i��\:�o&�l.��"mcእ�uۍ�c����^a>���c�)H[��7�1n���	<Z�,���4����0��\Jy�$��S��q��:hr:�HY,�"�a�㝜w;��N��DF*����C
�Te�{5���Q��وS����!�8�Vfl�&�I}u��?���Y�ŋ��g�	�X3@{��O�i/�2y�8���O5��a��������������	EZZ�W����,��'��0Vg%�����PT��@��Y����.iOt�J��[=�p7�DzY�l)�L��+U���$_��I��t(*��qFnb���W�Sǁx�c7��\)M�����?~a�y�7�ߗ.5{���Nv�Y�3��h�Q�d9b��RZ*�1H�\g4K�y���%r�J�$Ɯ�a���<�^�i���)���5�����;�g*��-c]1���6�`�T_=$l:"D�:-����.�6���F�]1������U��v-Ǐj�d�NUa˻�]o8��rA5{�c���B������S���K�J��d|�x�g0=�DolP0kNC܌�1Y���ٕ��%������G�ϧ�߿=���������Ϡ�e�P���:�&!|w���x�K2+'�dBj�2mr�5c�խ#_B=m���4˲̻nlmf]*�H�F���Q�A�?��k��Cs��|�S����n�E�6�k����OX��Ke��l��u��'�)7�(ީ�8���lVD�S��p�ټ���J�6���9/��M���>M�p����:�f�5"��e��gz6aٝ"��������jB�Lw:{�.�X*�7qM���έn/Mp�f��E�L�gf9P�4��uwg�o�C_8,�6C�A��g��s�Z҈��	J��O��Ǡu�}�P��e�Dɹ�U��a��G	�)*[�]
�{�,w:u���y4�Њ�OaDs.�9���Tcs^��O��os��r$�+K���^�+C��-!��x�ƻ)"K�j[��
P*9�tG
���)ȸK���(0X*GP0�HCC��
8�y����Ьǚ����n4�E�
z\��-��֨Y|�IC'�Ӝ_�����	�O^<H(�aE����L����&�</��x9{�������X�%f���&�X8�\��j���ikF_�U�YB�缄�U���y�SS��Ƚ���� ��$O�������m���[�	4K�^EJK�V�[��ɜ���êQA�bE$��iﯿ���˼�>}����ߟ���?�0�2��xz�7�J5���I�1�Sv8{��{.�f0#I��4޴F��DW��Y�������a�m�`o����:F�'X������ף�����x"o~d��k�捕��8�;������{^U.�v`3�ha���Xn��/�I,aSe�9�t���u�?��F�]n�	�%G�I����f	����޿�|�^�c��L3����8��>#c)��sE*��4�.�SG!+��ʅJ�o\&�lQ�������tF�ޟ0+:'qA�u��7ߺ��X}�3<T?��ȫ�;m�_��<3��C,=�FW�F=�O]G��v#R^�+�ݷ��T�{�xq����:������ғ�c:RnC����n^AΙ{��4�V���-mK$l�x�}�,��lR}��E6W��ǻ*vO��;.���&Z7�'���x׾��0����X,Z�y�|u�26�l9P���B�V0֮Y9/��]�Ou��e�ڬ>������~�O��͗��R�h�#���vҡ��
�ݶ�ᕥgn������|D�◧���,ɳ{|F��*���:�^w��5�A��W���ǯ`�+
�gc�w���n�2EP>|�c�gf���y=������!�ar��2�B���'�ZF��1�u5vݐ[��1�ބ�)X���^G�'�?���2�d_�ϯO�����O7�~������v�`����iS�!�z�4�/醑|�W�w]"�d�v����2�78J�ֽ^��r�	�=ɼv�+���fTD�]N1��Tqͦ���9�����:�:ɇ��ݢ�{�UA+,���~@,�涴��K s>����:u�:��j�&w=z^K����W*���טn��) �Ҷ^HȫΒ�&��lz���}~`�|�<ų��᡼p��͵W�;fv��΅�4
Q���`Y)�h'hcP���g[<L[�j�8~�7@_�;�~����"���O9�E�o�zfP ��ia��R��m�,\��·aZ��=<���,��
I3�B`mi�SN&�T�9�I��G�Lco3�wC45澶7g�n�*}W�M���řZ�T���C&{��&�?<��Dŷ'�{�}#2�RP���Ӛ�s=f#�F�k�����j+(3zBQn����vO��4��݊D�-�WW<1�@�zH]��󞠳�K�K�VF���0�O�T[��Fm�_L<9�dy�h|j/�.������O�;"�%�K�q���G.�ꨇ+�m����l~A�8gq��I�O7} f�y+�ͥ�{WG��o���̀�l;Q�kK'5��^���ϫ[{��AS���5�'fp٦��U��ʬ�r��/S�g�l�י�雵Y�|�Rłh�c���
������<����`��p@M�3(M�u�3�yi�����t+z�� �(z!6�K+|׹*��6+�����k-�w΅�-���o��F&~M���A�MN�¶�N)oZn0`h������oز��Q�.Rw��*w.�s��d`u���dw,�P����r��*�nmx�H��2S�A�s<���t�H���ަ�g��N�Ve
~�S�b�$����Y��^uǦ;�W�"�(<�3M,��G'M�r<�9t����w0��*}���X��̈�qt�2#U÷b�HX)>(��=i66X{w4���%�%)��R��㚔�u�h��*A���/��ъ<��+��\ՒD6c�n���D4۠^S���^��6��X];H]�a��M&bđJ�7�#�Z��n&������Y��Z��~�pT{�֕
�oO�sf�*;�bPXrֹ֓��j��.U��h��::lDE��d�\ת�^�t�p��}]�P��Rb�Y��!#U5����������ʂ�v"�Yf�Nm��:bY��%��p��]Sg ���j�V��z���|�Y���e͗�5,}Kv�+���%m����'Qp4��7��X*�<��+�����t��sYz^�Mx ~Y��9�Xʿ�$��;��;�C�{�FylW#:��f��{m���sI��s^q�W),R�{����}�����a�~�O>{���������۫��,��j2!ۯ�3awfקJD���.���{do�N�j�<�k�Du�+Ǟj�q��#��f0�\H�A���#}�T�KJ*��7���nj�m����T�<�ɉG�؇���̋	��Vq-^Sy��������W(�;Z]��߇��~�1���SZ�����(]q~Ǉ~={�3ڼu�9Bh�2}�m�<��`��2p��nS��Yn��Q���q�V`�Kv(�r#Ú���>J}�"SE{���@��@cƽ�#���2�9�?`hz��~���,�$ٳk�,�B��w���??Ҏ��|���4"9]i����y�]�Hj�k��̕%~�e ��2K�u4Z��1�F㻄}�wW9�l�X�{�n��TȽ�QM�YX�Ω�E��S�2��G����A�iީ�8�mr�ԶE��K��aA*���Um�"�w�۾0�i�����Jl��,��т����j�!��{���k�d>��q!��W��g1��?7W��Q׶���f���{(?$�\"��`7����B%өSq������?@���=���a��r��^�Z���U�r��X;�E˪�6���D};)<��%0!�8�Rź}��Ӗ�ԥ�a�6�� �sx��]C6��?l����>y�}�<����|����F!��ԝ��ܾd�C3�dzb�W����[�)Ǻ7��u)��K+S�e��(�6>�(���O3�z�z��������!���2J�Ca�a��o'��m�O@������h
y��\�Y�StdX~��B��7z���~U�����h0\���C���h6a�P����	n_!X3�sb�F��󴞌m�-.��0��^8Nu��x:�Z|��ON��r%Vڪ�T�e�i��y/Ɖ���y��lG��[��O��
푇�~7{є�k��3�.�>#׆�c���U�TA]	��>1�26Cllj؎O�_�3L�.�^g���w�
�ȱ�)�ޖ���<��4/6@v�"�0��N9\V/C�ڽ�o+���^����Y�b�n�o����[E�9t-�ߚ_Y�	{��)A�+�4�����2���4+� ڪ��c�Xdt�1��E�fx�.l:�X��p��XApzO'�5��E0�c��9Z��Q9�TUWMz�M,�g4����ifg��,�a{�|�c�x�a�'��kp{6�O̾A#>���j�%iMsͽ���B>��4Q��e�2\�]�p��pQ)
�|�|��;�����%J�����4㬍my����t63�(_غé�']�bԆXrG-��z���Fř	{Ӌ�7(�8I��Cy@�+�3+�����xY��Oy2��O���9ɶ� �1кD�E�D��dc�C���v��u��ßTZ�qH�vs:���L��i�O��ҕa|���W���k<�O��\�+��t^�y�//�b�#��mb�c	���y�U-| ��L�fȬ�J��5�l]�È��2�qY�e��z�[���<�����a�ͪ���9t��wt��)�u'g(Kۑ˪��Ot���Ę\��r��Lx�f:/9�VX��h��w��+sUi^���|f�����C I�eDQu����g<@ͦ�DK�k�u}Khi(�����z��r|c^��~u��#[�:�A��>��4y�\��� �~[��߃<,����?V{*W���K�Yx�Ő�R*���C�u�=Y��׉�iP��)��I�T*Va��O��t�=\�m�����b��g4z�b�G�� �����)�ot�n9�#h�k��^�WL3�v��m��f�I�_'i�0]/�q�db���fs�s��z��Y;{�'�8�{����=�ӴE��!�A�S�rd��wy۬ާ�T�Vw%�LSVa�al�W�Jan�YP8�Pޞ���>EχpfUh%�z�]�$y�#�o�u<��y�ֿ��Q��ő���ݳ%N%
G�����
tƬ���C�r�v�/���m[�&�tw��O�� ��6��Q��ތ��u��BY+-�X��1��Ŵ�T�UmX��i�ݽRdx���EG4�]X�rzv-n�b�I�"��@T�z��x�9s�mT��O$�vM�i���M�[�G����-�4���Y��?�Ш
�n���i��
l�0�*M��fY�_�d�cD)����n͹dm�TAM��Kw.�=̉�OSA��[bA�*m'%b�Adǚ%Ig�݁3z��.Q�I��NwQ�=�-;�z�cd<U�\���{$/^Ǎݤv[ڽ��QX1s��y�4�{5����=��P���v̓��=SN�G��������w
�F� $�R����X�lߞ������cz*ł�,�;v�r�:�f�f�PV/_e�a�d*f�;�=�l�x�n��ӛ;|��.��!���[�<����^�04=r,�*a9ޜ�����&�z4�P��+���p���JpHT�_+��b�Q�����t��N�Kf��*�%�^�ԗW0_���E�^�������\������Ȃ�:U}��F��S����t��(�-����0�>��e7�)���K��CK�{Hh�D�7p�n]��S]í��(�*���KAWKK�Y{0��Ϛ;ȏ�L)�n��*���+�)�x�<4�g�
'�M�yLjv}8xV��F�J-�j� ���	Ug���8�݆���=�`>\˃6���D���Z��:��oQӁ;L1Zډ������(��];Su��*��DJ��Sy�z�D|��c�i�7���qR��wf�-Tޚt���c�e�$f�V���5�ȷ�WB�m�
����A��h��1��k��Iv[�#@��>�j*�j<�V���oaY�MM�'4�Q��m5���wE*jg4#YQ���B��	���ǩI+&��#�6P�6�U>�x���h�cE�j��!��)���J7�PQt8�����l��n$�+2��ܩO�j�%Ǒ��]�鬺���h^����+E���Ge��D��`�zʆE5�-Y�z��]��^-SN��Y�5��Ί�l�o�i�r��	r)���nqu7����֮�M�vsq�p�Z���@��A9OT��<<�\��^��(�d�n�nʱ�y'|f�IJ�+����wNOv��ؘ}�S�^������Uą(��e}�x�%$��*�����$M9�G&�ɀ��
л�8��n�)�_8;s�U�6�,�D�~8�I�Z��e�_�$[m��Q���å*��"���ܧL2�-lpƜ�r�V�8"�#����\�F�"���|�O���Y��i������v������y��S�T����y?>uՈ�I�v{�����T�Q��ͦ���%�?�>>�������_���_�g��C�"*���gc:�������"#O\Q4�i�����>>>?O�������~����~�>Gl��%���QM�ƻ�4��]��tI癮�G�{��>>?��������G��f_����q��KӪ>l����m@S�����@Q>G����o��b�[�ۉ�o���S�T5���1�#��/����vĄ��w������5�Om_}���I��|�Iŭ���c�U1�'�6�5���E�h�b��A�X���uӈ��-�y���$�]�;�KAם�>s�j��M�݄�lv���%A�ϛ�����"<ɹ<��I��s�����Pk#�<�8��ڭ%=�U�h�&�ձvN�i֪#��Ih>vf�����>q[ͦ�ܝ;m��b�(�6z�3X����[��󎢢���_2Q��yg�ww�xG�cZ�wk�x]��-���N��HT�YF(���:G9P隻�k*Ev}҆S�Df���p˚6�p\Ԡn�a�Ջl�q�9ө�ծ�����緛y��1���?D���_��(g��`ѐ���N�<�D?*���|�L���JqS�ǞX�8��曳Z�]��!]�����ǎ�S��YA^C�:��U�N��&zX�o�E<��x{nO�ұ��X���n��5�̄(�q[Й��ь�
�e��fm�Ћ��GyosH{R#ѐ��{��B��b�'j�C�d��s�v;h��Q������k�5�=$��� ��LV��|ܯ��x饾�9\%��C̳4��C�\���L}�s-�n7�N�����p췍���g���*�Qj5����'ҫ�Uk�3��m��4���W/�ɷ���)?^,��9�5�ykM�P��T۠�ߖtJݗ���#�-.���o�Z�!�q:��J��_�:D��Jc~��PI�*�o����C׸��b��vfP�ѳ
YU&"H�Vs�@��N4�oa%���2D�.�"^3��:�vw<�q�e�q)�HVr�٩���μ�oN��`��8Z��ʅ]�4�Yq��������2r���C���>�ςy�h��
��qV���!�;�w����?�s_X���Y9\�x-D`�MLư���E�ؽ\IO1�Hud�Pv�PnMV��0_[���̦�v�`P���ܪ�SS���W{<�,��w�ӕ��h�8M؝��NY]��7k9kW�N݈Yj)Q��Z-�*�0�O
NH�|<P�@!� �����h+U��Ld^�<���yP��(��mW0����g��s
_��ZG>��p�V�x�F�ݬP[؄3 ���1	��"5?K�h���<\P9�	��q�F�UE�����xݨv�i��
/�z�7�����38!��S���Q�m�Ն�w�S�S3�#���D�yVܹ{�7|Q�̆��u����Ńb=k��g�X�4�Eh�;�+w�d=+=K�6H2zm.M���s۲�b�c����c]m��hH�'�]�m{27�������r��݁�EN`:_����J��6����o�1I���u�����8����m7�CT�^�:�t6��O��\�ؼ8Y�k����řˎ�y�4� ���U�3ɶ�۳Q�׾/�5�Z4��J�$<`0�� ���WG�q6B}�-�27�`���kw&D�����6�-h���������Mq5��_Bu>�.�S��rh39�zn�֫t�3�p������c�N�+L8�k�̈�5�mc��%cP`j�a��܏��+��Uf��g\��a�c��<����7(��]]�0��Ӭ�{��X*SaT�C���%V�BX�K�T�YDVw��=��F<��|<�a�<�C-�Ņj�|���e{{>�%nݍ���UCu\����=�M���MQ��׌����9��`��V�8�,�W�7��H�5҆����Yl���3\Ӟ�C��=�����JNU.������W<q���v��y6A�HF������Cwڋ�h���G.<��%�),蛵����gp�.sz�jM]��0���'}f��%ב�2:)�I�7�Ȇ%r�������ٶ{����:��G;n�6!��儭��Fݭ��ِ��6�t�R����t�Л��>�h�]�S�T���7��r���5��;v�9Ǟ$3�=M�:��%{>)��sp9�n-lHkc�+u���nWe㲲���l}�z��&��n���9ԛWT����;3�����AE G��c�|�se2ff��VW�1��^]���>u\�f������!?~d/���=}H`�g�T�.�Q��h��=W�����*B��h(��	�A�t\H_�Ug�:mߥ�%;�W׈�4����m�������
�/	i:e�<��v��fg�`w��jɎ*�"�I]�ؽ���R[�v{�O K����>$y��r3<�U5S	��v�m���7�%_�[L�M�v[q�$_��t�nx����Qn�jxQ��Mr6ԼW�|Ξ �z�q���<ms����޶���zYz��x��FOH�ǯ=^v�_�.�����Wptܲ�1�f�wٞ�B�o��ɼ�}�^׶��x-f^�Q!��!�U#X�az��Z:��}�M?���{/�"�VR99Ia�W�v��娜���a{�i6�;z� ���c�5�����^rY�䜡|U�F.cKF��q�f8V1:Z��B^�W.�+������|�	e�N=5�S��\�-�ō�i|���dO��-�"�W�4�p[���id�w#{�
1���FjY�"�+��z��
���/�ٯ]蔋���ܽ�Q5�Q���7g�d�_:H��䄎Pei�=8�c�;�g�5>�q""�g�0����{C;VT╌6޽t�l�Z+�����h��bT;k�ǣ=X9��m���ʦ��̀�䪐]��t�� �*0+�#���0� �Lt_���Y;��{�7" C���}aU-_L��Yn�yD4�<:�a	����<ʖW���nB������J?(�J�]�G-XՒ8dz�
�վl-B�lݮ뺨�YꝬ�:��'�
�`�ܺ�Y�7�tr����\���v�k�#@4�� -&}�I�߷u]wF��Ͱ�17�{r��y�G�����5��+r�~NVߤ@Vn���h�y�c9kv*zEeX;�x��rK��U�6��:��p�<z3��~��_��Kuk��­���*�k��^W��Y���t6��m��^��$�冪���(����kƳ��@�{ř�"�p�
�h�l�mL�A���s�zp6�e����ouǌ������M����o(�a���(�GCa�r��v�{����|�L�=�5߀T��G��f�
��K��z�ƝT�dm�����f���Ν-�4"#���˞w�FQ�z��X�+��#��t�a�p����|�)���{��oia�u�a	5�=a�O��,i���[=�S5ge�O9_`�|��� ��Eԗ��"�}��]K����o�0t][[�� �n�o��9C,�P�
N���_}s+��G��=f��> ��H��u�f�٘|�>��n��ڻ�\�_��R�qA�Z������߉|����:�r61V�Ww r���[���Y :m��6ޥ9�{�c1�nݝ2��"N���U��`����E�0��鴛�o�{��y���ZF+;���_�+���H�T�����J������n�;�A�ƭ�Kz��L�����iupH����kF�>w6��Ty��۶Y��սX̷�h���^w�u��Ff�q�y�x����q��� ?8k���n��iő��g��g� ��L��R"	���'����]SWgu��z�� 4����\,�z��:�̭�6%"_O��Y�s��-2�;�L?v6w%d�Y�Kf��������i���7t�	��M���k�rz۷��]��0q�,h4[������ˑ�}얢̡�7W�Z��V�/z��I�Uƅ_i��I|�f�e�KG!�B2V����﫩���Ew���٢��34��C����("Br����<�7Z�t7��oT�iQ���EWͫU2�:�^�}_��Q�+˥���	��1������Ӽ��y�`�a0��M/<y�fD���k̼��|�|0TS@k-z�AE��WeS>^����׹=�j�INGzL������1.k���}ު�|��{�\+��y�Ö�I�9�n��S��aì�j���ƏY�x-F^��H{��\b��!�!\bjɛζI�v�>f��t�pr���d������7b��|!�o��J]��~}�3&��ꏇ�������%+�Z���5��V�^2�~�h8���h������2�gΰ�sy���{%�4�sF�{��׼:h��if��z���᧧��Lo��٨7?�z�t���`���h��ސ�w��V$�JJ]��#"��M]�Y�O���k��ĺ��p�>v�[�N;�r/b�)�`�\4mܨ�km��ۇy������g�U�-1�����!oP���(��:W�b7��
�ڼ2�U�3CBOb�Z��*6����˨�J Ir�"��w��Z�&�s4���L�V���pp$O ]2p]�=�)��,�1n�KHfp�?�ثcls��r}��2Z�>�5����U�.<@��HF��b��/z�[�� �s��"+/w�iSG��͢�8i���p��s��#�E�b��W9L�e�n)�"�˓3}��C�]Ɍ�;Z�׶�ve.�6�
N��ݶ�Oh�|�zD]f{'q�l��+�`�o��Y�pϕ�V�=<F�q�Y|w�\�7�!!x���In��hgf:���q�:N�ӑ�\y�x����7��`M��Dr*�a���7���;X��{!�E�W�w�&j�%dc/�w�^�Ǟ+�Y��~�l���>]n��ņ��w�U�G��S��קg�j��m�����Su����݃����~V��f����	>��jƾT�c���ӆ)z���.������+��B��ܪ�n�q�d%rh����z�V�<�(�ۚF��Ơ3����3�]sηټ���ta���~��׾=�{w���ٟ�)�������t.M[ �= nw
�ikI�J��Gq0���D�˨ǧ�ʲw�ݸ�,7q�z@ϬJ���Yj]���k#�򺼡m�f-B7� �<�x��"0N���|��Vݐ���; E�U׵���9�rO�K1��9�wQt��J�QL�DL�]T�tѧA�?�����:�{����boVݿ2i�b���@�~�]ЖQK�t����i�ڃ�o�}fҠN>H;�!�
��B���z��Kw��N�t��\�=Sk{�-��êzn��V������ǅx�oe©���W8i��x��҄��b	pyS����6�7�μ>NK,�{�s�=75�d��ѣ{�m��)O���Ɯ���}~�P{"�eC���Ӯ�1/Eo����8cF:՗�� �����Y�)�U5hB�;��l��0��>�~@d���bW]�l�dg�%>p�y�Kn����e��9��®��q7�M���'!4+����?�r�N�w�,z���a{��P��0%�oE9��,��\о��|�UZs�������sږ&���~T����C��e�5�9ʃ7j�*�i.�Z})>;z����p�� �*>�X/�BDA_�/��v��~��k�A;H.�Y{�����ϵ�˙aE��Qv��E�7Vg�iڎЂQB��9�����w7A}1�U��T%�W��~�_M3p�k��i�G5��Z��)7�WK+���j�� 6�ؒ�� k������"w��3v�Ci����1�gy�a=�#;�^{U�#,��`�ڌ����`�u����Z�$�Q�~�U����'�+�x�i��R�A�7�n��++�2�s�LB���R���c��ۅ"�X�S��T����ԅ��n�muu]��l)��u[vK�uKA����>�Ep&e�rO��j����yU�?��3�o���g�<T��,�d'���Q?y�z���a*"� �h�ݖ�F��[���g6��\�9�Hv��ۂ�f;w�1�n�E�%�b0#7�)�䧺�.�S�[����y��5R�w1�`#g���h۫�>l�5����`��J4���lb���;�dK�]����������i�(��wK�OlZ3#W����w���f\[�}X�rF+U�ν��U�/�A��wJ��YR�I��B�x���@�>�k~�R��D�Uq�����sx����uB���R�W�w!�G�6�����]�yV;�K1�䐼:�3��RۅS:0ջ�J]�p�.>'� ��n������r�giB@XӨP� �����&�l�3;o{���э���:g�/<~:��Ø���լ�V�x捩�G(�k�K�Flj����;³����{� 85`	�WA�֫�Y:KTr�ax�������JM	g�}���нw/��Ot �5m�2����`���m�a��]ż�U����5��p;3a�)�[�x'��tZ3�G�:�;�@��y!2k�'vR��"ȫpH�����q����I��C��8��Q����
�̏H)�'�b�=e�={W�J���{/TC(v�,[t���%n�Ao	L.t�z�ӕ4a�w������C��h/�=��䂰�1�k�-f��Lms��g7v���V2��
xyt��z��o�9��$��n؞ܙ���K �c�� �еo����wi�;O�J�']r&m�sXP� ��e�s�\);KRenY�����k	�Kb�E"��̷P)%���"ܙD���&���l8��v-�T��I#&����@�����q�Ǜ��^��)!:i�ɔ�9�����IC���݁8�p�;�:����o����/0ݛ=�F0��pI]-ԭ��ֳu�zA9"�:��%Ft/�_^o CyO�2SV-c+��w45�[�j;{+d�pT�Ӭ�����ͦ%��.0��uڷ�4�y�u��ҁX�s�[Ý���,4�w�aEÛ0o1��>qZ1��7Y�4{4�E�ʾ�f�vO	�,eLf��$�����g�]1֖���u�c&8�m�%�����
oZ��Z9u�<:3�*Ďۨ#�qdښ�6��]�g���K\�C���@�j����W� �[����k'�7�r����W]�[]y�nh� .�L,bY4�R"�,��r�`W����8V��vcCj���YѸ7K�0�Z-S�w�A�N�\��;�mdDq�C���[�� hL�x8�Ս#�nI]�γ�D���F�_fͤ�*c/2��w��m'���2�tGd�]@�B�-��<��〼�+' !�'e�>��w�\Q4蜹�n��`r�����k���.�h�Օ0XS�����֌nġ��]1uAL5"�k�f��6�2��t|������af�(��"d�!̐�:���T�k�v��6�K&���u{�$�+��xDe�;+m��iɆK�����cʝ
� vZ9:��znl)-�sogY�ˊ³�<yg8�J�s����'7r�m�|"X�хD ��A�#^�u�4qN�h�*�5��c���k宸�+�mLM$�=بg<��>>>>>?����������=�8�6�k:�TF���y����b{:�=1�5��h�ۯ;.��������|~?����������f}���:��/7{y�8��_��v�GZ�z�A�,�ͦ����/>q�^��Ϗ��������_���f}��0Q�{7m���DA���G����W��A�h�G#X���m���Xǟü�q�qh���8�ۭj��mwj:�b"�h�F�����mbf��Ŷ�cX��5T����ϝ�v�8��'lѫGa�Y�>m盋�v�DZ���D_'�������S��,j�Ѯ���<��>tq�b����%<�q��9�):��Tk;m�����wm��'j�s���w�4m��Z�X��;�;o;���m]�q�v-��1T�F��b�lEy��i�؏�Tu�*-km��Z��Z%����E���>��m�>c��mb���-MlZk�E�Ukn�����yn�,y�y:ӈ�4B@��P�qi��w;z���[�3�Vr�%�I��P��5��;�=k���ݏK�&gu��Im�vx�.r.�V
q��`-j�|ٲ�����q�\��}^�F���ׇ�2���o�-�UN�"�?p��q�n�Xa�k�m��ˮ̧�+Ya�OY��yWq��.;`�T�[�� :#Y�����
ެ�~��X���Ƚ�Ͷ��ο7"�1�²�*��M(�\vo��l�jׁ�c���dק��9��,r��'tl>�
{V�w��32�E��#C\�W��O17�Fg/0��(����C�'rɌ�G巫٢4�L��2�lX+�!�G��H��J̦�Xṩ�i����N�f`�>���:/��)�~�3�)J߬ȅW�C�T���ͦb�u]�s�t�(2���W���fM2�g�O�.�amA�����'�;]��whQ�O;�k1��nW:GG)[f+9]זAY����sb�)��;b�i����ȋ;�r�t-w�����Fu��<[{B��~���	�hzu��N�DgN����C"7�]��5��Sֻfl�����F��礦:�ӽ)\i��D�E�����oλY�cq�䦍'xL���J�쟫쫯�)���.b|�\����XC�E0[��O��H�X������_��4u�_D��ق_챒"H!e����i.��xt*MO����H.y���iV�he��Vl�sݙۘ�I�z�� �}�'�@�1(��%�L��­��nޘ�޲]{�Z���{e*��ՠC���7e���&����[ �٫�T^�H=�֌&�+��Y�Br�I�ga����C�fƭ��͐�^��ܾ��O�����$�{΋�]�6��w�N��٭9�^-�c79&h�ts�}�-5� ٛ��%��ף�bg0��):�u���g{����)�[�jc՞>q��v*liuf�فkW��޾�a�!�b���~�˪�w�N��8�lv�n_}�Ջ&���DXК+��gdn�՚mߥ��]�6�� �+�����9�Њ�CY��<ĵ�L;���b�g�W|t�J5!�):G)�Z� �����Z�5w�mY���&$�r��8WwUZ���w��jJ��*�C��	w�\U��C�7n֯�u�m�t���0V�M�΢�r&Qh��p�{��#wԋ����Yu�����7�Er���Fp��A��:.�D��4O��nQ%z�{���&��L�^a�^5XU3X�)1@x�Fk�|��X�e4����"_&�j��
�Vǳr=Y�<�Hd�|�[}8�#���������Ls��P�s�s*9ɦ8�9d�W�R�%S�8��Q�S;�U{m�Ak���׮X�+hQ�:�4��f�l�n���)o>΅��K$�Cx	&d���p�u=�vil�qf��<q⭷e���+=\8J�>���ٝ)�[�Y�ާ�z��� }�ё��=w�������f$�Ե�*��[>�]��
lz���޴"��)q�2�R�UזM'��Kg��#��w��qd���Vr���O4z�`n�޿s��vޤq�"l6NK-�y�i�\m�M�'7�1�Y��La3뎢����JJ��o��V��:��m��:7D��~2]����?�R�j�~�#����ã�:w�J̤��O�gU������e��B�4X��Y�#eї�VE�N���G��Tģ�Г�����jVx1�0�_���*�}U�ߞq�X���εғ݅"��7�nْ�QX�zu�K����<�#\Wp�\�1]A��ga\��	,Wﾪ��s�����_{���ly�d�	;Y)��aWݦ�.]�O�BX�=��M����������q�=6&
��r8�����_���l_R�9��Hʈ7g��ڴĿ�����9o�2O�F�L��Q��6&��UI���%��к��Q�$�q>"AT�1^܈�mZ���b�a���B�7sN^��0�JB'5>�d��,�$d�5��L��3�ÓJ��3��!���yj��-�DԍHd���/���k-Oa�*q���s�b.�w�� :�n5/f���{�*�ea�aq���Dhaq�&�m�2ՙ�}�WY�-���g�����;y��Ϯ��-�s`�1.k(�{�Ŧ�S�V��+��v�ot���j����"��xnֱ�̳g�،���݆��Dc�q�8���UĽ[̴[3�D�|VfG��6`;��C�]F�,`��%�,%�M���u�a:
�ph�k�vwaVĚ�
��̡�ec�ioQ���d��J|pqɽK�����$go�����k��Ƞ���7'�V�XܖFp޾�h���� �|�&jrM|̃U�ٿn��x���%t����d��5��1��ȃG�8\�fG�c�ڪʄ��V�P�˺O�y)�[��q5oC�n�Gm�V`�b�O���7��\+J{�Ǻ��	T=�v��4�:ip����5a�`�l�s�.l�t�;nm��5<���U�[b^oxi��~_ �o >m��A(�-n�F�g��Cg!�Y�����m��We�-kwIrYA(�";����Q��y�ۋ@l�$��{a��|5�@?0{$�a��u�w�M��˸�q-�e��4�}�im2m�H���������=���_y9�L� g�0���yC^��n	h�!�˘n�L74�M����P��o �ʵ3�<U�E��ǌ'g���bbb��{`Vj͓fpNBd���H>a���]�Jw�Q��Tϗ�Ŕ�S
V&���u3l��mi�ᘓ��1X�Y����[�oE��Fܺ�[jYȷd��۶\9���Y�Alg4��7�4/g���?D
xw����.������U�j����ڇ�ub�YG��Z��Q���яW���ʧT1�`}��kĶdq�D+�V��|_���!�}�*)6��g��٦�����B������9#�ɡ�-Q+l?Y�ߝ�o~���z�j�\�ܮ�i��f��������;��eqm�T��h-���j��	�Ś����Y�:۝ۢ��c�ЖRM�J�h���R�`d1�h��i��I���6��j���ڣd6�%`�]���Ű;�59���/��Ο���X 2���Mj�汩t�6����.#i��Ufh~G�4N,'P)g(-��[Y�[�8l�dR�Uq�B�L�J�}��i��XO/�h?e���g���,.��"�@Ԋ�Zp�WzH�j�b*�v�Ui��`ÚղqHM����@@�׋i!n-9/<_3��V���z҄���M�Q�n�m��w���b�
:����3��oG&��kwC��swmƳte��SU,�wo�XpݾV�D�7i̪x&�Y�+.��i�)���&�%�T�����%�g��@�ФAÛU����o3���%llĺv<sh�}�$�J&�F�C]i���mfWVB�,$h�Kf���O�f.����0e �0���5�\�����k:��X��f��~^ލ�hM�"�/?��;S�.�nᬼ&�7�p�xuQO�kzҧ�)�����_W�hO?\����ex������/C�N�y�������Yi�McĈ=Sx�)p�ݮ>�[�Z���e;���������%��p2��=M��5�̥[3W�xE����S|FK=|e&l� �C�D1��XD�w*Ҝ���ܭ�@����O+w���Ӱ2_:�k�D�GD=�[$���Y�C�^Jԯ}9������#{�Ԟm4D�9�ǥ��$�O2%7�tuW�䶮��^e�'\q4u��^a{�T���PYV(`_��y��<�
�:i��*+�¾���q��4������y���G�61V�W{����:6���%r}�X]B����QW�U�s^�F'�y�	�\4������}��ԃ`yp������Nt:�$5�,�8.cA�}�>t�[�X�����@O����]�f�1h����C�������Â���;3X�`K�E5ۑ���x��yzL�K
��F�G�����;'�^�y[}>l���-��F���f�܊����W9^Vµ�zn/eG����)n܀��~ �de�b������ؤ;�nXF<�ޛ��*f�zz�"����`���r6<�d'-}��=wi�\�X�л�DhO8�3�U�f��n�}�R�K����d��߮���*����|	;�1^kh�}U�Tv�P�s
���0��oTv���Z�u�t�i�G{y��KV*��#D�r|��wX���?]���=3@��-��㍯Ɓ�2�n�c�O2}|��751)��f:�{B�|۫zwf�=�����`�W�z��u�ZoS=��ݟ ~NU�1:DFs�ER�>��$c���/NO��x��U=L�Y�܈�<4�6F��oJhsƨve�t���������U�ߔ^]_��_~z���,5���H�uӛ;4�R�V����ЖZ��(usW!?�)���\��:^�ͧ���ϵ�\/� ���}��zEl��
�}�׺�ڽ3��e'��]��ge�'$�\OK�ch�GB�������$5쎶�������s�A{�dn�=��{>�<��Y���;�%tp��M?b�Ӯ�tz�v|g�n����m������4����ی���������z[*n8�u�<�^-yul��O����'��)��P.�STZۆ'��v��#��sc����R7�U�?a��}��<�N��v�1�bg���i��\��Sax��q��QL��m�Tsiw`K�ufW���f�+e)�����ޣ6(�X�}S��h�s�Sz;��sB�w"��ۦf�Lmv�g����������O�j��VI�\#>z:o�ԥ5CNlAhX���[q갹*ak�ڎf�a �i��GO�����Lo�ݼ\�B������+�;9����(����[$f��v�he�b5��3��ۧg酤�Ȯ��ז$�6p��R������q��1�8x��e����mֿ���ڲb���h����nN��*�cF2��~���Ԅ鴍n�	T��KgS�@� t��eh�S��I[�z�Nv�2��܈a�kQ�ۛ;"K�{�5�I�wq�]�}\�qN/��=�园��P,�����H�vL���>�y}2��Jκ�Wn�N��(�4��
3]��<����Nޮc���I��ٝ�����?82�Z�(�=5���"&C3��:@Ϥ�i�=���6@�o��x;������K|Ga"3�m�zՌ��Xc���k��`J�:¯N�^�|�,�\)�v���Y[���egW�{���ů�;�F��l���k��A8�O������ه�2-�ܝ0�m���fE�w�����ʆ�����<DeZ�Ҙ^1�/{`s������9ҹ^撱]� /�,G�
����-wl���i������K�_�t%�t�Y�SPN�T__U;Լܕ1
*���K=A�cR6W�ܬќz����ZT��KPb����d3�I&�tǩ�d�^K��yZ��� Թ D�WT]EAz�~��|B��e�!����*W.�Ǘz�Ë�&*A��.�M�}�ή�a&CLNucM�0�F������v��8$�Oum��5K3���Գ$��%d��ư��v�&{&+�I3 n軸�i��0�N"�R/�yI��=*�8Q�{*�c��"��N>7��+%�@�y9\��z�e�l����b�-lj�x��.8�Z�}]�>әA����tT�̝,{ώ�	��9(4w�v=iǲʸ{hjs,�}��I�������]�s �B��rŢ��>d���G���[�.J�/�g1855��/&gZ�'ҷ+g7�XNc�u�Y�VdRa��pqv;���nwb꺜�Mɦj�}�&b=uk�2���u�1��悳+:���)�r՝ @z`�hV�t~�h��m;n�S�b�Xq�*�H���������D�Gh��>�7s`�/$��kU���u��{@��hr���uѱ�G���Q�L9�E]<qЮ8�Ns��Glsz����.Lƫr�oE[��7�aM�;y�͢�5ʢ�'�3r��{��V�j=���$ֳ�R�����!yC	��T�3:(�s�cf���&��i���Y�;0v�ѧ���w*�����!n|h�6�r�l��1]�<�[\�ge��9KpD/�Kœ��j ��S!}n�<���l:)���.��t���-ܦ�I���r���Ĩa��(cO-�V���&�6�RSVY�jvƍʹ*�1	�.6
,�I\G+�*^]���=Pn�%Z x��74�<wl"�h˺�l���u�j�&�gx��J�M��ne��+8T�̝bȂV6s��'�${�F��3n�y�^�Q0���Y[��n��i\q�zZz�K�N�@�F[�*h��:��ʮr�d];�
L�cc.<�\1�J��-����]��� �d�
e7��S�Ff�&n.t�V}�S�}ȊA���y`u2��]oPdC����y�3%ѻSkO���.w��ym��
Y����Է;Z��k��k����s_.3�<��	!�ͽZ.��Ɏ劙7
��@�ms��=ؖ6F�-`x$����*l�;��Nܭ���$��A��]�i�g;Qq���Q���P��c�%���.��0Y�E��Ł+{��y�v,�GNl�\�f�j��iM���S�6ս"KX̩,mbȎ��@=x�ev���un���8���ۜ1h�j����WT�bۊ�-g.�fAKe$�.v��rI6��6)�A�=��q�ж�M�����W&a;Μ�{Spl܎X��dqq�5�V�Yϥ������-zk��f�C��������<�o�x�H����Δ��.�|٬�խ�B��z)���]�咷K2s���WovMAP<�nj�1��K(�(�!$"MBa��)F .Ȕ�lN�%�a8��@O/�q��G^m]�h�ڱv�q��6�S�HD��C�@���D0��M�#
)L���JO�
(b*��ƻ\v�.;��
�F�u��(��۶#��{���s����������?����ϧ��b��v�k����k��{�F�6����X���lb�0V<��kF�k]������_�����������Z��t�h*��AG�E��=��ݻ�յ=jz�ݿmxm�����y�����>>>>?���?��3������׻�ͱ���;l���t���Ƴ���w���l��#ʺ��]�ض�4�u�m�E�?\wmb<�w|��`Ӷ��n�I�T�V�v�w]�n�c�F��f��*+l��]��F���<��ϑ��[α�[m�n��:�J��鋯&��-�/���:�۫ͫ¦7��m��+���u�m�k��t]c�o��N�Q�����oq�}|�םƉ����L��7ߝ���wt�v�7j�ۣ��m��U�[V��g��`����V�oǳSQ��.�ݎ��n��ln3wti�?.�;����f64�]ŷ��o?��;�*�TQA�o7�\W\�/@�`���#��-V���w��s,��L-���ƻ�cXƔᵱE@��<�� y�wT��ԙ�\��� ��X��I�)|u��ը��
u	i}�"�s;�1L׭���)�VOrJ��ʥ��(�U6���`S��R.�^vgqu!6i�a/�;��Q�O�[�
�	Y��>`Š?pZ�������5ڂ���'��+"�l�m(TWr��mp��\��p�V�<3aߌ�1���a�/U�O6"\�_/�;� �����Kv�� ��ӂ��������u�׌�Qd��u��PKb7]�M��܈8��S�(a�.��r3,�x���=K�J;��Nݘ� �����":PmqŕGA3w�.t_Vi؞�9�o�U�0��W�'b�nw
�oKb����
v|�ȱΛ�^δ9�d��
�X�)��b��8�������+�*f�;��k��ޡ�S�*}��{/�$;�Y%[4x�<�+�ɫ3���7�M�-�q}<�T�s^W>�A?���_Cy����\=ǱS.T�f��K�2���]F�g�{�?�5�����٤EoX����h���l�f�u��X�.$<3>�qUL��adE8��{��B;389�#z;�4R+#ŝZnj'x%gA�h�l2A%b'�N��
��7s�_����I�h��m�>zUt$P*Jk����7�\�k�M9���2�_�s��\i����D��v�5�U 1����"�oex9"\Vn�W^�f��'7��5{yr��'2��ǜ�tt�2]�g(���iz����f���5?2�+��H7]�������y��-xUې����0�{{�(��A���)�F�_�6��d+���l���零m��"�;`����<��^�R.2�4��n��>.�qP{i� �(�*��JQC,�㾜n7-a����J�Ȯޟu�TWq-���'�5FN�)[c�\�	���Dh��`�eݯ0�$J��3:����T+���轧�Ț��zZqίZ��Ƭ�������/ڎ�%W�4̊��u^�}ʍ�'���+(�>ɝ�M�;�.2�ص�@:�}͊�@��A�|�?B��pV[݁�f��2�v���W��;1	dM͎B� �n�9�Cy �WQ�e0�ʺj]���p݈�E���[��A����%o)�'�g]��O�
1�ic���[$�N��׹�-�l�s�嫹u|����1]����$��G��ϻL��Ӧ$��0�;�􈄜�=��ӻE�6�-�1�b�n�>�/�F�(�nV�W��.W�Qo0�P�6����T���o.J���`ɊY��j�3�f�Rô�l�*_F�-�b"[�7j�5�q5�Wk݉�~�fތ���&�w�ơST)@�;C0e �e2��dM5z|e�K��*�=�~��@���}�2\L2����䮶{���g�� ]a�U�L��0\�a�'gw��oʀ�W:U=���-EwzLE;�����b����Z�*�o�1��_�p��uqg4��މq3Q���]eB�,.�	u��Y(�-gU����bj�NCp�m��'5k-�Y��#�M����9������g6���)�q�6�d�t`�� mH��w\�Ԥ�䧺��4���_��n���"
n̉gz6�H�:̵�Uƞs����:νߺ�༓h]-�1�)�z��o2&�?$�D�g:��q̉m�ᧈ��F�bz4���V_[o� I�;o��8�%��ON�����������y�Z��g��m]tc�con��\$�ᯯ { ��b��u�n�B#�*k���R¸���2��a�������=M�~.�(\&��;���d^<5N�>�*/]L8444k����|o��wV${�Z�HO(*n^U�~�ˇ��L�
�����������[~H�+h ���T���l?MՀ�����f鎝�,�K�d1i�"�pYV5�4g=�|�O�d�z���[�&q�O_:k��51�����_J����{=��"U%��7]����p�Y|2Cn���!�lH����yF;�nr���2g�-vฺ�;�&�����oM�[lgK< �+��%16j�秡0�G^Z��D>a�c�]לEX�2ƹE�$���֕Q���Q������D����:�{v����etQ
���'&P��]��n
��	&��U��x�p7]��M��t�5+Rn���<�)�eZᘺC���|��_\�{v�yh���)�N���CWHm8忉��J�Ђ!�E�IZ$��-lvڦ�wg&�6��ok����-�X���KR��v��<}�T5+[\��l�R�55�8����ʑ��L �|(�,��lX;�A$�׏xx"|.��pl��)ʶ)��y�p\������ˡ�u�_�)���'WXY�!e���v��� ׍X(����|=�ϟ�����O�Y�ǝ�3� gt����ob��d;��Vq��������C�4��ѱ�����V�R��v|��(k�׬x~���rV�@�Y#��w��yMȸh(p�,�]}��M@��~r."wi�D-�,N�7Iėo$�=�K�f�K�`H#��&��w��{���I<�/��+�>�Sv\���Dw�B�$�zQ9+0�v�δ�G��篢V��P��V]Rz���Ӈ��Frj�y���׸��s`;o�L΁{�J��!qh ��V�z�N&����;�U��$$C���7�����';ܣ�j���O�gr���u�5l$6��޼�w�]�n�i��ʁ�A�����F#0�ًY���CcK֖-�4���q����5w's�S"�\Y��D��.�eqb#zMY��Õ%B��c�C<���^�)_�՞/Y3��gd��>��2�"���I��ܽ]�uqT�vq邦��A/5u<=,���9{jg�M�W���F'��9�k:`Y�����S���U���x�ڙa*H}�aG(k�hl
�#�i��bg�\�<ԤUª��cr��3}�����J�p�H^{x,��� �� 3�+vV�E<m��㍝�;jqy>EH�FDM̊��q�w��+��b�Yx�-��j6�Sj�[�ΖÚ��o�K�	�}����8��ZjnF�����K�&���W�t�F�=>k�jtL�W6������{��9������{w4٥� Q�
��;':��W��V�P+[-�2q��^Pr��c�*mǁe��I�aA��]��zb2�{��o
�6��wP�Y&�m{��Iݩk¬��w�;\���[�t���9~lo.F��Ϳ%�Qו�I�wv-Z{�3F<�]i���������w��P�����H��{�s��v�]t\���R9�*N�ta��Y� ��Xvp(�$�;�����p��t�`���Z��H�P4��������0�>�"w�1�v�upa$�!ш�4]҂���L��`���/�C1�z/�e����Y\ܦf'�F�m9-x97�t��ˍ��Dfה0�Я����.���᳎�([��Q}�7�p��]b�O���_}���ϐ�a��{ Bޑ�5��&���H_DS�H����}�+/_I�W@%�wۈ��3�'���K���ޫ������M��?;�3۾&�N,�����n���q���^q�:d-�db?\��5�;0�K� T�En�ah�p;MN���f�2��1��ه��0�EvG&��t����r��X��v7Nm{����ک�r�\� �BN�&T��v<�"5�T�Sc��U3���+Q�q!�@�mT-5��w�x>G{��2�'93��g�s�,���������d��4��=����~ݷ���n˞"�fh�uNQ6��s�Y��S^rd�;�	�U�Ʒw{�D2�ʟ<��U�a�v��^Eq�&���qDz��oc�b�Xv���E�}.�D���r���"�����z�W�ɵJbE$��ЁӜט^��W��̭_p�gk�j�/(���y
?A�];��q�A���Cd�O�z�ݜhr���tr�3Jڴ���ۻ:�s{��tIP�Q��쀼<%Βtø�i��+R<vR� ��9l��Hk�Yа�Oc�yt�l�5xC�RǴC�)�����q�[*��ܨ�&�̙�+:�"cv75����uy�ﵲylY+�@��>m�[�/+wI]F]��y����e&�<�� �3�-~�ӊ%�9)�u33U1Q�w�A����R��]�����(�h}ڐ��c��܃H�FP��{��϶��Zj�}��W�j�Y,�+'p����c�B�ox��:0�t�:gm�� ��k32��k=�Ct�x��$��N"3��8m�I���B=�Z�K��=�n���^�H�V�Z����#x�>��xqv�Y�5`'���>��X����
D/7b������7����5�����5P��x���q/W��&��@c�h��3YH�}�5��Z��M��2�U?M��u�pZ���s�`(u��M�Z�Sُ������C�ʴ�d6%sZstw
n��MK����H�K��T���%���U�p��;L�]�6f!�'L4j�J �@�M���y:YKD���Ŏc���훉��0�)�����}jޜZ-��wF�<�������檎`����=�Pn����r�-�y��}S��`́y�	팦��x�5֯�D�9zi�wo4q���,�]�d���kЖ�M��+��l23�ٍ�e�'���՗����K\T��z�t6�x����]��[\fZA�+��,�L/̤ޏe�	�+�Q�1[E�w�-E�e�5*�`��&[�u��15��S(��U��:���]ٱm��jS�cw6�C�|�ɲM.�#pL�2���YK=Y�-��o�J�R�ֳj鷆�/��p� T�g��Z{�Ȃ<��5��W��s���a>ms���Z��}���<\���$���K�+D✀��wz������a�H��PK��	�z&k��e��wCwf�m�U�wds�-=]��75�S�=���g7������h�U�΀Y�9쪣u�2�,���͘��F'N�+��ޣ����o�f�K�(b��4�!\�V���;�=�f�玴;tfo0��S�+%S����G5�a�+5v8�F%��x�Tk5���H��O ��`9;Qp��Ѽ�eX���z���nl2n�/x�;�!��J����1�tD�͡��G��X�|m
��ی����y�6Z}1����}�T�W6�O�ʽ�Φ��9ۏ���Fasw�oD!E���i6p�)>��r�>��Vj&U���x��{Ꮋ.�����w�����0��DЍI�a:b�Ϭ��g�MtA��x;��u����H1��Pc�Ǖ�g��w����kx˵u7�O3W A7uz�+��r��*�z���t}m��M|2���h��郴X�U�Fr�yd�F�@٫K_/.h��?~ld����H(f&Y<�;�E����c�eg�ס#ӗY~jz>���u�����w
q���qp��"%����9*�㥬!��j�ӵ.U5hq���7�ՕNe���mY#'��`_��E�@)�5ݱ���@���@Dlc�ȊC�i�5�	m[u3a���V#���Iwz+�b�C���	��m��2/%�1����Zn���N��T�:x���� D�8����,�fҗ���gG1�|)���0�h���<�aݶY
���eX[@5l
a��ֳO�ї���F���#���p�(H��,�.���iWSi�⎹t ԙ�7��x�\�m���]��CWg`�^�`F8����<�їo%X��1� l��U��iKK8Ĭ u�:��Mv~rQ�߻^��ނ�Ԯce!F�k5Xѡ��vӢ���J�g�K�ÝK�j�*C�&�ë�]�h0D��\�YF����AL�v��cQ�.��M�-��-�k�����Yr�v�w�(�_7��Zu	@�X!��� ��>�����ʹ��bT��6��(�_8w�S$GƸպ�F8i��{t^!��ˣ��^���j��G��֠3�y�qP:��0ie��AV�/$��=š|L��V��[�Y� �`�;��0�Z������̫���+��XAq:3dљ�]Al�3���3�]��������f	3��.ſ��^��/�/h�Z����΋ Әo*���I��gLJ�Z+����b�jɛ�#�)���1	i�S�:C�E[���;�GR4:�d��vU�G�TԜ��ג�N�R�B�!��,=\X�tܭ�܁�?=��h]�IDB�4�D�GY6��@��ft͸F�ir|�7P�-�>����{�U���K���L��淲��&�?NJ�OLb�w��l��z��z���k`��("�Ӧ��Yײdڥ�[<'h!�'5�6��/[7o�~�(��$�u�\i�g7h��0bk��ND�)A>Yx�8�	����kBs��/�*�9ղ�;f������C��o[�n)YN��8���
M�9�%�Be�@^fn��^f��g7��|�=�wk��ժ���XZz>�niء{ݫp,���Y����xY[ܣ�{Ú���a�1W#�`8e�0Ĳ�)������`�@$��K��S�)7]�Tr�>=v2�cu�9�s�r��˜q	ԥ�O쏡W������4�j���)��;j=Q���u��t]"�Fk�q�oC]QF�i������J݀���V����V��Zm��N���i�yړ+����O��bc�\�&J2�K:�e�ؕS��{'[�B�r]�4�Jrg���6����q֊lm�8ȣ��]�Z�)�LZ�'�L��#�>��r��ʙ2��-KcX
���ˠ��4�.�ᵎ�܉_�N��Uf��U��| �Sv���w�e�^���l��QQkgj��w���%��;�6K�/��q�yIv��vآ��o���۸���c��m��L��v#���c��������|||||}~�\��_�H�V��5A�[u���n��wq�v��b(��]��M^j�.#�"#cF�;��Ϗ����||||_��������~���v�1��������ъ�̓�.۶㻍;f�_X��y�F�W[��%�8����Y���������s�G�����m���+�m���t�Z��]���ƭ�l~ܗ����v6�Ml`�#3]���t���v4�qE���o�����Uۮ���
خ�uY�mUWN�ڶ��g�wy��Y4o;Q��Iۣ����ڂ��wWRQ]�wF���U�'�:���6:�5��V��1͌h�C�ۢ;cj�Ѣ��uX�cQDZ��j|�v�1E����]0�]ܜm��s�FΛR�m�j�C6o�4uk����i��t��U�vz�q�mqky�DQ��bñѸ�L��PwZ���Wj5�wu�w���_�Eq�mO���F�Vؒ>EefHq"����g�S�@��r!��e�NeM�.��ya��FI������W�.<ʵM��CĎ���\����a/��QQ��kݝGn���J��cղ�_M\�F��WcV�a'�7�Zଲ�Ȝ�&=xb��+|;��o0�DD0��z1�jz5�Kсt�������a�L2�{���4����a;��l��=�6��\�N����I��]񝅽\�oۏ:���b�����}�7�S("�]!+��Ml��:a�:�IE��3{����p���� m,�l�oSd9PƬ��w��ogз���M���(��"si�/�g�����{T4$��=���������\�w�n#O<���q��Ƀ�	{��W@�3�M7H�a����h�wuOo�e�fl��t/8��XPİ37T?w��V״��}���#�N�(�|��}q�u�OM>kO(��P(R2*x��k�=W�+�.m��c�Z�(m�u�o�����<�5�f���u���2�un��x�a�+|����\Sab��Լ��o̽�/yt:�ݿp�q0��|3c(޼�2�7���ɩ�����ǹ��7�I��Ɇ�v�;G��;���h�sn��:�@l��\�8k�Yʽ�+-�_}��'͏=��\],/39�Y��/7�P���M��}a	�F��o���ys�ַ�� 6�`�*&wt�E5Xw���}'4o'���<�1v����\�e?@���2˚��2Lc���z��t
�f:�Tu8�d���t��
^{z�7Z����H��b����^ܹ��$�g6�g2R��9l�n��˨��$�n�l1v�˫S�vvgG�!>�W����s�IU����Uݝw�l��U��Ce���Z�4��w����śl�g۲�'����m��v�xk���qJ���oU�SK;��Y1^�
��rM�Q�=��zr��2�jjg3�gv�M���q��3A���Lj��=�P���kf����Cq� ��x�����4�����,�(��c.C��yF�@�����=�in�cF�֎��N'�ԛ�km�����Ճ��{�mh�=~�]2�Q�,Y���#pP��� �ȁ{�"ؐ�ks�c_v_j�����u;3�E���}[�K듍CpBڹ�ow��U�M�gT�g!#�����ܐ2�nm��A��~����b����q1-����ӽ�M�㺲��ؑ�+j�C:<3j�:di�^�]�7Ң�����;���XL�8��&!��M�w��7���6��p^b��`��M�Ջώ)طO��.Ly��kD��Ǳ�3���j��V�`�gy����'����C�H%�����c���W~��b����b��Q�nZ�v�4�.�����Y���E�_2�ʬ=k��Ԣ9��f���Õ��0�\Zj'I���!���*#�_:�Nl���m[V�N��gk�P䆒�x��<z�H-�@x`F5�o&����ݭ*���c��M6*��!'�!<�J�n/�h���]�C:�mp�������6��W�e �yKj�Ț'b��:��P��b�4&�r1�LL�F=�`W5�oe��y���v�nՒ-8�Xe��������߯��ݕ*lF#dY/6�F�����Ms=�3����.5��7,�_ze%]�"R���K.?:���)F3�"�v�-�q�]�Όr٩p0�O��ɏwQkQ`��j�ާp�ħ>�VR�����k�gJ4���\�"��cw��5��wF�H*�&�K�oy��yf��1���3�t���5.v������:\;5�p+��w��V�jm��n&C�V�Y��;�ũJ	&�f�O�V�7J�a.�IgR�����j�ۇD�K5���g�{:DX1O��Va��S��ƃ�Y*�O6�"�zڟrߑ�4�*����۲�"�;�l<COM��dRڝ��)VQ+,?4bm<��u��O��e����e��#̶�.���vc�����Ӯ��NĽ���U���p�B)��l�l��<j�'��������[���Q�ÙG5��Z��q��l�+!�H�
�Z�+�Cgw��G�p�֌g[6�����&��}y�=:�ٱę ę��]��C&3�-����3��I߉�q����ؾ��W�/5s�@�4�<���(��t�L���j�G玲������'�w(�ܨh�v.H��b���Po8WV��l��k��tc�a�e�.�/)�8<��=�T�2|-�x0s�f��fu�Da��c�v^��w%�r�jT]t��[5��[��FSt�Aǯ�U<z(��vڀ;}v�41��7K�[BU�L�� ;�d���Sꕸ���uJw���tު9���rC;C�M�b.�u����
�Ed�{�)�d�Pރ�#�{~���������Ȟ�-cWtf"Vǫo�b<�<jdd5�5 7Dϗ-�CK��ѽt��"�Eg[/��tI�Ue VeRX�x�3�KZ��!�槶wח�²���kFs����q��%���7�Wkhr���/e��s��p����t����'qO���"�=v��-���Af��<u�8�}Ƭ��9��}\.��u�U�4��1]�S}MZ�vV�1Z�dfY�0���l���U����5��]�ˈ́-l:h$�K�=3xСbƒ�\\�q/��o����ܵcVO��ò��oO��j�4X�8��-���� t"�x U����C�Gh���#T�'�oMl�\d���]bFO<�v�[҆�]�	�R�������zw�&l�j,|S�خ�z��mhs-oU��#���b'�owo�����*��eȑ��������E{u�81}�M3�/���@��t	� �Vw�q���F�:�	��̌r��\ڋ�:T՘���tiʳͦ6�M7O{8��=�� 4��Y�uECV�<5�1�o%~����e�NI��3D���*T��l�ŵ�[cD@~\����� G@�lv��hs�n}a�!�����RC��Ց������6���g�Y�|�fU5f�uHq�Nΐ)��_kPO58$�#��ֽd&�!�c���{Jbk���p��������5�"d���#׾~RkTzݥh�k,�9b݁X�eŴ3<��K��#�N�u�a�M(��xBy������qMb�x�m�}w͐�so�ט�7@��|�OtRp�n8�·њUq�JV%fIWu^9��B}��;��h�:�y�Kb�u[�F��>����%�	�.�c�Us�֚h��
 ���b�Ϟ^,#ˬ���7P�[~T�ۮJ�Hģ$nS�0fp�!sH!�����x�wl�&Zv����g@��\� g��s/v�TOIR�tR��w�䛺�����;�7{ ���m����7�fE��<tm��q�~õ�d�q�??���h���_�m��|>:�a�W��2� ��2I*�[�z�)^��.�_��/?{a�ߟ���Pl:��qK��ٝ£���@ҺM��(�y�ihN��e���E���K3͸�l���7z�Wib���[An�qAO4=��=��|�Ӄ����͹��1�p���4�|I��q��\uHK� ��>fSk�/��d��q�O�s��g����%l
�/꠸Ǎc�� ��ďykVυ��GF;	�ٱs�
�i�jX�~�Q��%Q8���Of�֩��g/99����h[^�O��o%�6�nT
���A�iW>�*ۨe��9m絘�'6���i7;���&}�mI�홀�ȱ}�94Nԩ-{�������fN�9;�t3ċ��f�����n�z� ���<c������7S�)�'�j�cX�B�2%�^j�w��^�Z���@2��l��=,�hu����D���z]*��:�)�c-�*w����0�O��_{yz`����VN���/m�-��k���ۆ�7\��b���zn]37�J�[�5�iCQM��|�38K���Wo���f��'+���&.tb�C5��p����&(�����1������'�P�}���՗L�-#��Z�3A�e;1��Py�W��qw�J۠0\a=���qG�o�z�{���s'+V?����\[Lu��=���;�rا�V�	j����񊾄��-�|�4�:A�1����7�}���~mX����ݩ����$�ο���d[�g�[^�'2�=�b�k�ʽx����[̤c�IG��V\Ы�KB�̇�e�^F��WeR��:� ��W��Q�����ycsuX�5��A��@�Z�����,�x_J�b=�����yPc1U�N�n[���	3ʗ:�W�����~�]�/�y�3"��l����%V��di:����v�:���;W��}RAޡ1��B���	�jEUaT+��B��M���`��c�>�[�댈��a���L����Y�ʆ�9�/�Ζ\�)v����H.V��'�16ëBTZ0c}��f˷R����>fb�\��O3-x�6$Mm���������¶m����~zE!e�J��.j�iw>���L�J�nc��z9v��^5+��,t�yf��m��W�W���8�g���ٽe�Yܟrk�^7^�h����1�MOS;J^6ߦ�xiQZ��-��}�t��A�{�ᅂz��EÉmM����C��]������_ú?����`3]<��2������Ɣ��o|b�9^�)��4ǯr0�H���Z�x�7�sm��&��AKw�h��^yy��~�@A|����>��K�h>ܝ�%{p����f�u��݂��&Q�!��t�8�լ:�vfT�/���HZ�]�r�(�݄OSV�R;o�m5��}#v�_�T���.���\��b�/��"��ǫ���9��`����rV��O��d�Yl���'P.�G��T�T��"�����ڝ6��3c�J�Px�*��VeRX��V�d1���b�4��dM�����B��އG��;�1��.D�^T���l~�����?8�����S�M�}�y�g��J����;�?M7�c&�P�;�>�w�
��c^�T�f&7>����q�㪛j��wb��=�h��R�ra��Į�gŢgb�ؙw.k,A��!��V�����EZ������/j۟h[|&x_��l�Fۥn�[�]�Cs�^�wl��� �y�+\��?���}�j����	���ڿ�娠S�&&=�W�]����zmI��&�O��Ժ�U��F�U�u�n�7nR������w.��V4�[c�vW��� ��.���4�f�m���}���Ne�F)�<m���s��2��3���V�g;�v�������
h}�]wi���m>/��I�����u�^�÷�óڳ�e�5�󌭑I%Cu�Mo��܇��]=��^���M�nh�pk�/}f~
#/�QU�n�K�n�ms�;c*2����\�gD�����7 6�~�m:�,�³17>�x&���B�nJ�'nrowv�N]�N�,q�,c -�^�=q�|�����?���?���� �
�����G�l���EP���㏡�'��o!|��U!	P�!R��HBQ!D�$�HBf�E%�����!�aUaEG� �"�B?L��
 v�UP�C
�wp�
��(�dPBU ��C�B � %p��H����H �*H�� ��D2(!*�B!�B�!"�B4
@���!(�B(!"�B(!(�B�! �B!(�@��B ��J���@ ���@ � �@ !"�B�!@$! ���B�@$! �40�P�B�H�!���B�+�	! ���wp!�$!���B�@�!
��C@ʄ4@�Ȇ�:!	P���BA!�eXB!��d�HT���?�A��}_��E�JTU&�~�������o���g������߄��������G�x/��~���W�������_������?� Q��eDV ?��?�����?���4��?���?�* 
���������$����a���0��O� ���x�?�b��8T�H��I `�Q!�HH� �I`ID��IYD��H�A%�HT�$	T�$D��	 ``@��%!aA!�H � RBT IT��YVP�d`YFP�`	Q��e�`�e�e!�bA�E�A�E�H	$Y�bfQ�F$Y�iF��hA)�ZP�E�T�Ċ" P	!@� ��RB	J� ��DL� ��A�"R!0	B�B ��J�$��R���pb���������Q�TJ �P�@o�>�������g�
��A�>��������*��������?����0?��1�?�'��_� ����O��{���@ب�*�؇�0���������@����/�&��!�x/�?�������'��8 �Q U�������� 
��i@}�׿���#��Ϸ�?�� ������>� �
�_��ڨ�*��?�����)?�~��1�`X>��f�O����>~����'��>* 
��&����D�� �o������'��� T_�0_�  ������}����pd?�?��PVI��p�MA��` �������ǽ�oEJ�/�J�B5� R*%�%V�������	Sml�P���ųRPJ��*��M!M�km��mIUJ�XP��mk+f�m1���!��b���m[i5E��cmKK[5�ef-���R̳lSak)&
��Sbem��)M�l�֪V���Veն�����\�j�ж1�J�mM6IU2�6�4ګ[Z֩��6D�ڬY�T��Tl�kTki�a[E�*V�ki�M3,����L�kV��Uf�mm�
�Ō6mZ��  K�*�-6جmm�٩��t��)J ۷m��d���6U(���ݮچ�Mf���ڕ�VwN���j�ݬri@�[]wCL�ET��sM��E4��m���;�  z��P�B�
(Y]���B�
(�A�;�
(P�B���燥٢���0jC�b������4�ݑնʄ�Uj�ڶ�h-7v"h��묭�j�3%��cY�����  �j�%��]��k@Q`m6�d���v�f�R�Wnt�(��8
kZU�u�-�4,��T���wr��F��]�[-���j�i�B-B��l�ݶb��  Ǟ�zi��T��Up֒��cR��5X �:����W ��"���]�	;wW@���l-��ڰ�Se����  ]�T�J:c� j��c�W@��qQ��7P���:n Q�ܻp�Pc�҂�ꎌ���B�۔�f+T�f�mB�U�hO   v<h�(/l���e,�2��\�P*�wj�)s��Q�:VѨUUF�m.���n��vi�Wa٭3F��m�HI4[m�  㢴TomU� n�: '8Ӡ��  s�� 
sW8 t��  �v� �[� t�3�ت�ٵ�j�ږ�QVF��   gx  �8R� �+ �K��  m�@ P'v8
 �� 
�� Pl�:( 'u� ݵYh��E�m-��Yljl�   �  �ۀ@��  �  ���P �ۀ  �un  9�  �� ]��  s.�km�fm6ڵ-5b�Y�mY��   f� � Mv�  !��  ����nn  �e���w  
N�� �۵`  #;� �S�)JR �Oh�JJ�L��LS�QJ�41�JRP S�����=@  �E$1U&���]��:2�q�,bRC�I� G�H0�n����v��-JڱC�������|����!I>I$$?������$�ԁBH�$�HH}��y]�m�0
Pd ��;K1+%�R���P�]�a]�b��´��qYInd�j��2������i|`��o˱B��*C�D.\�u@˜�b����.ِ|�!J찯�e(1a:�7�c3#�ꡳ0�$٤�ͨ����33hk�i�uښ3\)��Y�4��*r5��㬛����u�3Ih��0Cq�hcO/$nj����/���M��48^,D4Y���v�1��[q�SN�Z)�Q0���x*#��^Bl��rn����oq��\% �P�2��	-\��V\[��݈�`=[Q| UpU�lZ;Wtv�Tåb�!�܃d+\
V��
$Z�/P�&�[
t�ܗ{tq�f�i�]�h:ͬ�Z���%��+�i�F`�pH��.��or��)̐ �����8�N0u
���H�u�2��U��v�W�<	����z̓awF�f��X��dMr�9�bT��/*�@�7+)�Ưj�홷)��4#�[��%�0��+]�J��F�&�qͩ$p�wVl��T��bT5��N�P��u�X.`�ٍ�CkC�%�6h)�9�*��Z�V�$�_W�`�d&�@�uV]�	�#�j��66���5�sT�+J^:�)��	Ѐ��LZ�%�ɫ)��u.�Ą`n�T�3&�����%@�Kg ���-(cŌ]3RP��/:>9$�]b�v��ٷm�Ib�$D%Yӻ6S�K8�u�����u���!$�mٶbH�m��A�kpj�.�� LCS{C&�&0�.�F�i�%e܍���ҲA�2%-���ƚ�x�ws�Uhe�ש��-�#F��jہ�H��Sf\2�"��:�R����q��*���[�f򘹲�ٱQ<j���9I�7����cA�f�:mVn)�c����SW���mEr���b�R�LE�*��:��/FF�5Ռ5�b��K4�p\�����d���FU�rf���&ʺ�`�e3M���{���'��a6ٺ-�T� h0����C@��화�%�m����\c�b =gBt��"�7�p��m=H�em�TV��r
�h�[�sjL"�7y!��`��U�1�ش�bi�����*�J���^�[`��Cj�D���I���.�H70��yI'z��QKb�ӣ.ۼ�B��)^�-Zٛ�c��ɪ̆�����-�ǅ]� ���ةF���PJ�,��ʦ��N�oQ-:��m�eJ�fd |S�l��CtT`^'XȤF���q�F�n��N�9l:���(`əQq�V�/S:6����eZ{5&ۢ	���o��%����M�CU(@�E��T��=� 
�qkp��bӽ�4�O1�í:"�3dҤ�r��Tx�u�UC�-U�!����B�a.��j��jbA e*� ����I��.HH �76jz�e$.5AHZsꨅD���j*��ݫd�X$bLi�IՍ�T����v�`��
�m䁠�'E,N��#'5H�&�*LtBذ�t�Ŕ�ZӺ�U�FA�Z�F���K��e�<z#���"M�Rx���w0�����������e�z&F���Y�n��M�m�d��"#ZN�)�Ѫʐ���������lm;�S�D:J�
j L/!7/����vb�u���@��I�,	c2����ݕ+2cYVM�l,;�ٽ-^��TQ�MF�K�
J���n�DS�5\jiB�*�Bc#n���t�D��F�C�%���%�>ۭn���
�-�۶5]��yO �*l'��@[cq��D���Rކwmͣ���U�ѣV�Э9�j�˒��׵t�5�+j6�r�2gq�ʀ�qP�1�y��Q�\Sn Ḟ�Z�;23����c}٭k|���S���Ł@,;�w�@���R����*��LY�,T1�V �D^���,ߢ�c{U�v^Őme0%��h�P�G.�O�U,h����[�
U��s+]�8 �CJG%�6bfH�;�q<x�KnkjQ�z%� �1\����蚺�y���[�Hث7h[�-���ݹy�KV0�T���a`��B�޼��2m:�����y�z⭧t�פ%Fd���](�ӻ/�!sb<�h��zم}��C�
�Y���EI�豮��^�]e-�YGb��q*1����)�р��G��`P�o6��f+Ud��ٳ2* �s)]�r��%��
��aU�W{�#u��KYvc���:-G���ӷN�8ӕ�M��(��^�C�4���m�.&��S�_%��<V����k,�����Y7X+@�w�e�CK(�!�44�Q�OӔw)d�~Pӑݼ�V�n<��M!(�#�u�#���m���=Ƕr��Ȑ��3����8�c�V�`�&�b���~�ư�ea�x�gv�f��S:m�*S��T[nΕ�Z�F՛ؑ)SU��PmZMJ̘U�oN:̗���H'A6hɆ�U�`e�5�Re�̣�v�8�]ٙb$������SP!G�L����+Yv*e��Ȋ��k4%t�::ӭc.U<�Iݢtm�s(+��M��!�@�+R���QфU�з����s�z#>�܌��1�e�e9,l[�Uk�gD����Y���C!V^�j��$�ݬV(����Y"�N�Z���s��Vm���B*к�3t������L�����B�n�z����J�������8���ܑ�CD0P�X:ln�ߙ)�2Z*���Q^n3�����ή�͸�A���o��ך�E����Uz
٘+(��d��ռh��%���v��A�[�>I[���(3�%��
���,���ƈ�eź�v!GK�2&Ҭ�/e(�-a�"
��e��C�j��){�\��#q��AdYq�TX6[���m|�1y��6�H!��mb���Aa-����7B�е�qhRt�v�ն�
�����Uj�h�	K1���F������E-3����l���1�jG�N��y��!+�p^T)֣-72����mQ�/�R�v�n�N(N�:*���!{KC�X36-R0V�ɷ��F�]�Բ}*�����[X�f˦�0c:�s����t7�GpgF.N��{-�ū<Z��{\qӅ@r��f�)y��t�<O]��lԴvn����^",
�P4Sq'�)�kl���c���^���T�r`k}0��Nm+nc�>t�%�S��,c��mG�#�)�th�WGt�#RjRh��QL�VV}�7[f���՘��L-6�S��e��L�X1;Re�o2�
���j�'%� �R����&�KO�@��b�t��ْ`�ڱF�H�<N򍂪�M�4�j<sS��t�p��#u�#�y{'��r�ҫw��t�j(�i�nM�R�EC�0��b�2g)������B��5m����ŵ4�c5���kz�n����eB:���p���æ��B۫aoڶ�%�\������y�L�4�6xnD�P0H[�kz��Ν��]�{HeI8�3{�CH1�ڂU�lY҈(����j��눋�^44;��],�&���.��(% -K��]���J����,�(�ޅ��Nj[P�w�u�eTǧ��1F����q2�����@Z���a��0@�ԡ��;� #b��z7���̀ �;�A�+X?F�Ă�F��ݧq��HLB��V`�ZO2�y��46�j�;m�]��ɺK��iP{Kc�`�� �v4�Κl�i�x��d�J��Z��-a4Æ;�ʹ�Av1V�Mlź�p-sJE�5-V֦�t�5u�hL�}a�ŷ�t{�XrBS���(�ɓ�v]6F����RT;GiaenB�2Zٺi� �y�D$I��R�d�eFIH4m`��P�5ՕK\(�ʍ�;�B_�W��Me�x�ͽ��4�a  �ܶfᤡ�ٽ^�0,�4�?�`��7�Pir�XR��@���X+�.�UCs&�U%�A�	t&��f|pK���Z���&�1i�7�����(G�<&�� �ś�(�*���Z��ѰM2M���,k5%Q��^V��:�aFV��
���h���[N��ϖm
,ݲ�R�p�Na:S7�y�F�CN`�So�qP{�~*M-���W&��K�+S.��l�TKx~�U+) tT�����c/mԧ�N���J�ٷnй��tf�]eRST�f�&�bDc���N�m�n�ʌ�6wmAg�X����a�E܀\���"�����Pj�{Q$��Р1ڠ0�/e㻊?���P ���cy#�#�q�^�F��{�F�r܊�%�#;�n�Vb���{r��.#���TyE�Ki����tޭ�p�X�b�dl��SAjń/.��9b��dmShj�E%r-	hXK8]G6
� ^&2�ou�F��B6��y]5b�Z65U���ԒTvV�Sc�v��ܭ�X������h�C �N�)�l�,޳�dd� J�aGpJ�q��ݎ�ڮ�G����H���e
I鳧��ۻ��s"T 6n�u*;�$����'R��{G��#F`͐ ����Y��NM�r�İ��	
���.�7���=e�Fظ�Cg0�-x yI���4�͌)QmD �!�U2^���V�Q� /KB��q��u�k~��Ȟ�̼��oX�F�bk�i��>�Y��z���ݭ����ktP+M�9V9E|���!���{�z���r�h*�s%4�F�FB��ߚZ��-�5�
4�R����m�ר4�g+]\U�qff뽳z�v�)�w�LˬF�a�v�ҭ��Q^=8�7��b���n�Y��|�:U-\����WA( d��ck-��4��)H��׎��(� �ɀ��w8�֠w�ዖ�^�[��!B\�ek*7Cz��Gd:e0��qk�$.^��sB��
0��|�t��@'�H�u�%�����Tƥn|���9��q���ǚ�I���Z����JPG&�(�ܬ����H�Z�����"4&���Tv���-i�!Q(�:�c�<�x�^=x�-�)��|����$2Z���8{4�M��"���]1	�K�*;&]mz��9�,�)��$9R9�ܲe& J��԰nb�gl�v�F�4^\[�Ua�f����V����56����H�N�X�Lʤe5������5d������q;[Ge����N۬�eM�ݩ�7�\Ϝ�� �CX(�<��(,f�*�+20�W��u�`�b�F2�mnTÙ�BU�f�P,�wyz�l�t��V�VP]��YI���j� g(ɥ�B�Y�R�'Uz���T)�(�����;�%�t��RS�
:u��[z]�����c�W���^��K�T��ȱ�Ȗ��HC9L������z!cp��kZ�b��I�@)XآlfL��I��t�]K�m��2���:$�4�D؃u`�i���,
�6�Bcfݥ���v�E�eO�	�c��j�"��Re�����7��L�I���3فm
n�Q��u�5���9�`��MG�3�sfx�`IcwXH6�کY�h��Ƌ�;���M�U`LErcOL��[7�Ln����q6 Κ�����N�PA�[���lV�5���6Ru6�th��/�/��%`I��aVf�m�p�J���5=�/^͑�ȭ�͖�����5.=ZN��w�4֑���6�WqP�ƭ���\����[�Q�%U��� h�i.��Ҕ񣗛�H�M�7��sN��ވ�ɉ��!Xi[Om���Ve���@��!{F��ҫE�ׂ=���-��S��1k.T��+�<k��⎋ $��'�Iޅ���X1���p�j��&L\ن,�y�CU���mQ)�J��j�h��kJ9wyF�ŗ�e�$[ɀ[ȐN�l:"X�ʺ���W���`���[��x�l��iI���(�CQ�V;,j9�jjeC�hj�,�V������Rدd�b�-h�ՂIJ���J��Kn���ɦ�zCzp̵������[�F���^�?J�j��KU��I%Hjv�Z���.�)��Ԝ�Ԝ��u��i�܂�`�E��5ˆ�Kn�wt��T� ��`(0Ү���<�S�
ytB�:�4Z7*�+x�TGL4 ���e��t686P�����`����G��]`Uö�F
�[R�%�Ŧ��ą��K�AT32�G(Ͳ^A��[:N٭th	�P�P�tKOi�ʴo4�j��F˃Ʉ
�X�F�DF�̵��3+!W�,��IjK� ݦ�!���c#�/Z�p���a�J��U�ڳ�$0
�(��CtCpɔnK����F�e�S+.	BD]\�ݐ���ړZܛMTz)\�+�JT�Y�$�a{Yl*J��ө������J	;��P�ҷ�2����b~I�>�	/$;�Px�	�k#�Ұ#�n��u:[6�U�0͹�a��T�U��QRXm���4�R8����V|�8�f��/"˸.����ЭMѥ��k>Z+J����ʑ�n`m���L��ж�"����\F��Q���Y�T��71QY���.�LP�w��YM�z`H1晩�-�ƳI��h��w[kr�ò�R%婵D��&�/lm�l�"�`�Y,�(���#�7m�0�
����/(N-�-
\RhŌP�g
�Dڀ���,хm
{�fSyWP�>2��e�����i���,��J+���c�(���X���cin�ib�f0��3i����Cyj�]d6�i#W�}Օ�d<�u��G�x�#��[n�W57�]�}�|A��np5q<v�}Q��$�'{���ŴEې�J���WSz]Af�f�,� +��B`E�V0^�	[�	�M��uC�s?r�������h_okM���N� �]�/6K��WWO�����pV�����|�\�}~$����v4��n�r�$�C�XU���rcE�@�$�f��	QW�2�n.}]�<nZ�����O���4՚�L�,�ϓ�v��x��e�8�'�v-��/W�r)[�X���r5ɀz�B��6�"7dPÖ����|B�cb��X &9�)k�꧃�Z|9��=��YT4Ve��jl�|���<8���I�M@�;n����{K��C�7Rt{[��^Q��=��h�K���{"ܓ�;��}�x���ރu �r���d���2�JxxB�kq�-��N@]�q.y8�_l�y۬�Ǜ�$D�o�}�N�:.}�@��o �-�fнѹOe�Le&v �k��
/N9��3ލ�v��}�gzM��9DP7�8��j^����cfM�]�H9�E��i\���z�b�WZb�b�wZ�0�� ͜;5fY��Α �PÔ;f��t#�7�s��<n��W&pț�2��f*z[�A����]c1��c���������$��<FKwá	�B�v\<_�I�͜u����^
<���I�m�ض��L<֙:Ľ�
ۺG�Y�e��`�4��n�y��ed��܌A}�{ݔ:�8]I;o"[�Zʗb�͉��e�|gVh*�Ƿ��$sz��A��R��s]C%���ekR"��1�B��2�J������f)�����ŀ�y�v��'+n���6S������^=���9�k,[�9u3s-��,�䭽/�jy�i�+�`��z=�8�'*�)|�'�+ȍ�׽�8�Y��Y�=g�-��/gԐ��wP�N�����jo25pQgg�|��i{�4+��Z�]z�Ş�ޏL�-���&�����j�5gM^ڪ	�\W�f%�{��4ƤfR�>؆ѫu��7c,<>TDM��A��{7}��V�M#�-K&z�}z�sE�t*�m���U�\�E�Tr�Fw�m!L6x�R�2�8�����F���Fl nI��� |�N��n�{��#��\�v�P�5�3��o�u%s��V�j�$��tF����Z�K�ZQ��ʁ��$�5��~ۀHMt��=*��1�HS6��xǼt@5U�=�a�E}�y��;V�U��ո�tFE�ɜ­�zދ����2y=3KN�r`�)D���Z�5Y.�*-Ր�+0��;fho�R�����(�"����%rN�����������~�xP�JgΎu�B�)�(3��k �C�u`L��z��z�!���wa�A�t�c��xVQ���鮡���G���G=^� �mp�S{C-�]i$鼔��fC�
ƭp)��p�[�U�"M��Dd�4����>���XB��NV��M�٘�[�lP�:��[6�RC���14��8�^�!��uţ��N��²�a�ir8J7�bv_<�Y88����l���rg�J�\�!�/�Ĳ
��@^�O�E^��c��Q�,L�:j�cV�{s$�t2��էt�q5sn�ր3U�;���U]'�d�38U䥴Z����@z�`h�,4=b\�������Ȳ�2x��i�*�*D^����]]�xof��.�B��q�8[�ɳ5�@ڏi�ǻ�/.��ר�����xvWn�-�b]��x3�N�b�,�Ed�������en�O&:�$�p��cM��N��7��
Uj�,�t
:�G������ʘ&��d��Zx0!�^'#Hv��5� �E�ze\V�bF5Ϸ�΃��Y��p�_Pֶ�h��i�U�K�əl��V�X�@ˮ���m|��
VtwHc��X:&${�n��}���������]�d���H�Ǩ�lwj�Ĉ�3�-n�̬r֕��BN���� ����z��F�[�|ۆl8�V�C�A\����f=c��&���^NC�`�YeR�2{i`7��P/�ߥ���Z��g*��}|�E��O{
� �pCçus��Z;1�^+����T;�lm�m��t��3��>���	�q7�����/t�1fp��fu�l·�Od:4gi�z9d�O��aި)c��}�;<�^Ih=0W�	sN�����T���ԳkYj�!��w+���vKB9����/�ЏL%�)���b GGg�Pz:j�1��b�/��4:;�E�;�B77��c��[s؞(b�glSn��Pu�:bU͞�*�5`%[���F�p��.Lź,Ě��5͑��n�w�%�K_G�; [d��nZ�b�b�uw��7ޥ�^�����)w�c��8ͣ�6i�rK�v97X���M'�YY��.�Y.��W���LJgtβ{}��]�"���bdydɠ�p��4���r��� �á{��;���~�Dc�C2�ب��ry�*�3�3�N}���}��ė�v�]�sܭ/y$E�E��p��oGS��y�n]�t0ǵ�m�s�ז\�^�r��?ٻ�v���+�ma�'t	I��8N��*bt�jT+5���t�3:�~�Y�\�����6�f<�7�xȓt��M��u5�q��$��j�O�j�h�>ї�l�K��/v�bv��A�s�m���6����o���g:�+�V��)�lwz��.`���8�]c�-=c�y̻��v�����u�j[w�R:7&��p�7��ы+�T���E6>W�YJB3&��9��#p�9u��jzw+3�yC����e��$G{Q�)��'�.|��mg���]�|����WJJ2���ȱ��ѼS�;�=�,�98^2�P'��j�����I݈�m�ى���L_��2�+ͽ��^A�G��k��˵£��<d���{gg<r�n�V��Q`fѸ�ĉ�\����e,��F�������@Ea6�(Ŷ��H�V�c�|f���V���H�K��B{}�#�mz�ڭ�x\(l�Nr,9�
WgF1e�u�C+�	m�;�Gn����9#�-����x�X�+:��=ʡ��`}����JwxU�7�jٰȋD:.ͳ�����[��K�tS��]�b�|+�C�=�ݘuf��iˎ0tL'� ��ĮO0�SU��gq^zl�N?���Ӽ��ve[�Ɯ���*��0�#�4ex�����=�(���W���Z><7�M�Xl�f�3�ǯ�j<U� V��
a��SJ�zv9X�h�w`�zot������i\�]ʵ�g����p.�#=3��0�T�tu�pJ�롨d=��rG'	%�055Y�z:?�ei�]Jnӡ�lEIA���s;�R�ޭ�6$�f����W�%��>Y/}qև���Y���I˲e�2�͜�/���#�T:��'�^���{0�J�f��эB����wO��4�:\����tY�i��p�/r�q*X��i��CC��;�7"�`�Ot��^�.�L���W:ƅ�n2���|+��]��E�F������<�B�D�9k��J�B��{�3J',��ѧu1ֶ�̩��-��%��oP0i0bS�>%RCI�����4XS�AY�яGj�}��Y&��:��a�O\�8�2�橇�0����{*~p!�;O���#}�o#r�J�d�\E��UҤE�T,](���G�8%-{���NHO���:�c]�${��v��	X�w>�"ِ�C:r��{^A�ݻ���\ �'{�waen�;F��Pw�g[�A�A�f섪JW3�����=�-��>	����񼝾�&���5S/B��sӰ�������=��en�}�]y����ٽ��=�U=�T���eJ�\ܥ�v:}*�&�|y���S��DtLl*�P��2�Znð����Q���Hy�e^U��C�Q�E|�Z=�&�"W{:�N�V��-F33a@>DH���r+銢����r�������g
=��:�
����J��,~��;g��>����nr��+{�[J���wC�����p;;��o�GMH�I�<$>��k}O5��Jr�*�:e1 /묕��H<|����8�p	��+��P���[�d��m=wI�z�8�B���z�ʋ'��ru�B�SD�F�ʢȠS2^�0t��TPl	ݢ�{��H8.*�|�h�� ��A1�[\���}eD�x���K��'�B��F�L���7X-%{�'��%�* �/ޖyC�՞Mt������= �yHV�f�SYJn��P��Ǳ�6�Y,�H4^U��D'���xܶ�ɜ,C�� 5�%���5�~Qe�*�1�̿OB�21͈T�aS�0W�6��/�+#�X�0��m;a�5m=U�۔��ӕ�^�y���(�����J\J�k�T}(v�Q������k�R�#:��w]".XY�E����|��3���Ɓ�l��Q��v>w����i*S�>r�8U�b
3����qb��Y��M�$�2�Xg~I-���l{�I<o5����R�,lu����6�n�er y0^Jƹ�΃"/`�%(q��Lѝl���8]m<��������[���uy*�'4��DB�op,��ꄻ�6�k����8돠ȥ�Lq����;qu����Y����O)�'��^�s�ï ]O��>l�XH��n'�W[7e�B������}%K�!;�%��(S��]�\8s��|2�['!��ݕ���T$�Ѿ�ٗ�Ԯ>ɔ@󤷔�6v���u���Δ+�k{��.�r�x�C.��O�e�дDn���|��b�Ge�x����.w�%Pht�ǂ��5�EFíT�r �]|7�L+�ڷ`p[Z̑�F����Fޖwe�9��X+���bAv�	�`�qO�K��S�������|T��T��bɝ���X�ܪ�P1v$Y�/����l�έ��F�S�nip�[�[ӂ��NmК(>ۆi٬�4��cw������El�Qq��"�O���*yx�n���$�̊{�xА�NFh����f=���~pt����\�f=$���Ýy=i�Z��3���(�b����H���ys\+Lt���+ſ-����(�9�c)\�mXl�v`�0΂��s���W3|�k�m���xVw|fO��Z���cuI��Mm\��,Y��;����I��P�l�+-께,\���$����ĢZ!���e�M��^�1۟��j.,��;��z��8*�J��ʗݍ�SԁݩΕ�R<����s���u	�>jXC���s\�g�k����1zl��3�寠Fݦ=1�c~Wz��?R����K�`�NX�L�����,���S�=k:��+	��&w�(�L�rt�<�5��|��wF!cT>����=D
�'���}���eD2�ǝS~����rĕ�	�
����(O+R�K2NH	��uq�/�>��IY�4q��uM�!�x�z�	)R�zm<�d�d��S�}ic�S�Yt�J�iY}N� ne%X��F����6����ˡ��8�!{n��2�� �V�qDsgp��{�n�-�}��w�P̚�u��Sޏf�y���0��b���R\�������}��d�o��tǜ[��ɂ�+�������u;}�DŅ�C{zK���b9{�ԇ���o`���on'�y�9�=���oJ-�2��l�<�nJ�����)���x�h���!]}��^��g\�{��jݭ���j�4��X��<�+G-��raq�2�3�6�=	�X�O����s77.��|�4z+y=���w.�um�v_��Q��4x������6��wsρs�J�7Օ�00��ժ��[�����پ��zDb�����)�.h%�}����8�]n�J��cJ����=W=��*J��<)��&��6�v�&�0΅�ըV=���.I��S���-�G�Ƀza�S��D�8H�z���#�4(.���r����w�z��`�����%2{
Vr�Z��}f;B�jاSk�Iy-�90���,���)��r�:��|e	��[���v�v.T9OR��w%ǻ<�8;]pt>\��o���㫭m9��C��j��F��}�&�N�"�;g�u�闩��z�eH)�yV����WW�갫o�W,k����������n�m�Y|�\��/Tu�*}�ȳa�up 
Z6p�ښ��"�(|bd�2&f�kn;;k�v�n.�h��o��Ԩ�Sw��ԥ�U塵{v%5�Ց��bV4����y�xu.X2������+'Uͦ�z!eB7��]ۿ4����t�oVa��N�Q�����'�G
ؘ0�;b���+A��{qpd�=�()m��a2�y��C;C!�o	i8Uݞ�=�[�����Й�)0h�����BT�v��t"Ζ�P�q����
w,{�}�&V��)�<A;����cC���S��.�K2�5RR�VwP�۽���P6���ı��:�k�3�ѧ�e�ܷ�S�O<��Aru�J\��Ʀ�P�W�C�w��Z��b��G��_oDa���=�[N�zb.@���L^��!���~�Fɕ�+���7[h;C��t���� �3C�ʷ@;X�:��5B�;��c_T��-*��'`��d��gƫ�&���}��c�m�{!��6��)zܹu�T~�DVU'�ǮzYa���ܤ�Ҝ��Q�B��^Ei9Qv�n�Q��a�}#Ω�k'ӽ���{7��BI$���@!I?v��� �������߷:'G�-��;���D
Q��l�9�X�'\�Su��6-я|�U	X��F�`��ueڦ��y�O�Bbv���������2g���9��Y�+�k[�bu��	���h�&��MΎj�+�;���=�v�����Y�t[�S#p'�)׹�����]����B���ͧ+d|m��!H�mq��[3��%p
c�Unr��+�����J=��K�]�<�ZM��{�6eH�O��[s�kt����P�8q������;����(�?+투��0�����5(ன̃����G.���f���\0wC�ʤV��Q��.����Pt��Ѻ�}	�)�0ۤ]/�����ճf�ʵ���;t�ʘ&T�������с1�T�
:��Ok��^[�\�������"���c�Ud�v�(��c�K ���C�#l��on� }����dYIj�,��^�FV�����:�?OW;��C�3�����t��)�D�5k�o�+�����#�s͸�45���N�{��i�G�������:6,i;��Ci�Òۙco���*�D�Y�vP�{��O�i�9p�Iå�IxO<�w"{��Zi���
�o%s͟M��[���\X4�f�&侁�u`��ךlk�|��T�͞ݠ�.���gM�����[m�awƃW|��Es]��c)������v�i��"�uiZ�y�;���skc84�4�����lo[!q�V�gL����Q���mݐ���q����c���ƁFg�4v�\ɠ�v�,c, �ܻ�Mj�D�����˙���\훱�'rK�w�{ϖ]�˙Ǻ4��^]�9�{4@���W����N���+z�v��iƼ�w�X�[C�mw�\�{�a��_7	1-������<��lN�c���+���Y q�6���`��AZr��j��8`��8��w��<~���� �N��Cw��9n%������{����t�IP��^V�Kt[���Ʈ���\�us��[��g����ǈ.���GsM��nu�y�6�"�EtWn�^����*ͥ�A[���q.뚱H�'1�S����E��G&�A)q�94����b�0�V����xa�`�J���6Y�X.K��V��Jmd�N�U�Ș�VR�hw���s3Fww�^���_Il��$&z�Cn,�ŒyB�{��,w��;��s�[�w\a=sm�d��̋�6��St�}���l,��]�i�O��/z�[��u�}3�K-�k���Ё-ˡjB޽�vH
�D���{e� �V��B�H�1DSڳEb�{�X{��e���l�gv�P�nOy~6DI��;��&m-�gmù�e1�G�ً�ѐ�QO͉�q��a�5w�Q�ͥp���0�1�VǠu��hM���P̻�dЦ�-��&2s7��IO-ܵQf���\ʌd.ܥxq*���-���y#02�iѴ6u3�%-3 ']QPv�K0ӷ�u��ӫ��˶ow��қ��m�.�I�i�7��4mռ�+�<q_/:gʥ`��$��L�YY��]'^l�F�ta�`&X1�"���d��ܴ5��(�]l��ڊvv�˯w����Y�)ub�j͋�B��sy�0pCoC|�/${E<��������7f��bF�(ø��n���]��L�WN�c�Iٽ޷C��@S7ԥ�ْ��W����WG+0"]377�u�v����Ϙ�=�v˫r�Ns�az��t'�U�i����!���=ɇ�o��f{klQ�AZ�77x�	���}C���w�4`]յ�f
��$�N��r�N⻭C�6����Pߋ7�r �y�nخ�ky��W�w@B�T�,���:$�zWՙ�ݾ�j�LT-�u��0�1'�<.��J(T�����"�g�x�(,w�`6�Lp�|���kn��P��;*;�*9T��l�� ��ou���S���S�����.��Y��ƅ��A�ZK`�v���A�٧=h��BR�y�z|=�\�Vr�F�VvLi�:ܭkhR�ٌ�܊�n���|e�H�K{lo��_nܑ�Z�O|cS�=�{���=�V��V�ごz����ufnstc�Z�n��@�K,G=ֱ��䯱m,&�yR؎��sy��㴵n�n���u�SN�1�|�[�YM��x��m5o_l	^�;'g]3r�-��0<Ǡ:M�3U
��e0$֑���d�u�hj�Ĳ�^��;��as��Y�6�+�p�Z���eH�Nj��qrq<�7{/5AˤF�X���.��G�eI{I=���ܾ���������ݞ\h��=*n�G�;N��)����o^���W��Q�dw���
;]Ŝ�"f����3�#��$ ��=��ӛ�d�&��D��q�yL��Ro�ƨ��|�F�Xv(�삖��'n#�<���%�f�l���}}DC���p,O�N�Σ��U�o��8�Бert[�mc���B���|u��Ѥ����7�� [G{2hrx�'6f�˲�a�;7�9�c��MC�c�VJq�}�%ۊ0���U�f��:`5�k���k�b<�ί�߸dń۳�-Z_	��'���ac��Z��V��=(Y�)9V/���BV�h���7��z�qK�Wd7�3e�Wj���n�S�%B�1 �����NǪ��,�~E�(�
�G�����A�	-=.{�UP�|*y��\̗����t@��ʜ��K�ֶ��#�Ć��(�������e�Q�<@6uг����
���o����=O�o����쇹��%�����u�J+	����~��eW&vx��ܐzJ>���{r��7��K%[o�F��5��x���,�ONG��8u;��=-j
�eη,KG,��=u�Cr7�T~/1v�r��Jh�.��l��f�Ш��Eve,<��վİ`(��3�d�+R�X���9&���z�}z��Ū}1���:m����n	n�����;8���V�zH��
?p��8��N˪��{���;��A��o*�6��J;�]+G��/Y�t�fņ�K��Ƿ.&5Bm�dl���)r�6�>�HA��� �� ��N��N|y}���pH�Z�D�z&�S�����듰9"Ï���0���B� �N���.��>���~jxA�њ���27����,������滷�h��<�9������v4�t�����&n�v{%�+�Ժ�'Z76�:���D��t��C�Yn��F���p��Oj|�s�74���`�cwk��V$×�XY2Ԙ䰍q�p'�VRA]�Km.x3ICS�I���d{�L��ɸ���Y��-nDχ�n�ƴ_���Y�1���.�*BLM3ϔ�'���B6-���[�R��	H��J]����3S`�^����\��y���]xT�3�;K�RP�P<���I�>^��z�m`�P!'7x,)��{����ا2l�};��}���`ǵ�'��Ӥk;u�&_^���ӯbt��3�B�w�&m,ɯ��T-8�7U�C]�b<�_7����U���<�S�s�4�=�nM^#88�.J�^`��N�]��N�2���Mǁgi'��b�N�ų��>N�Vm��He.��TJ��F�IZ�5�]�=:�:�Xt �3�i*�h�2�ly�U��?/Sg��w���ҟ71.��܅�Z��l�ëk��w�g҉Gaܮ�����h�8w���{�Fs��'m=;h�[#6s��ޚ�>�[���z�ʆV~0�H��{��+�4�{��tN�F�AY<�1fpr$j��s��E[Pj�HԝU�z�%�Lf��;[�S|֬�V;7���}��gD�#HdRX0^N�20�4x��'õ��,�HJ���g�ȱV%����%��4�2g��i]@�-*�:7)B���3��z���}�q�L��g6�#�뀡�W#�%�,왻�{��޶��Y`���[�����i��x�
��.۹.�3(�Js[�.�>�ñ�xy��=Zg.9�3,�yX�=2V'�v虱�WN��z��'4�oǢ�|��	g��dûm�X�0�$tQ�z��g��8JZ���g��-�Ψ�pn�2�Y���=�pkb���[���jZtrC�&�+�:�4��57�*�_��K��X2N��X������ӕr����Pr뤻N@-*c']�Ʈj�E��C����t�{3���|t3�ꥴ�ge=ѭ�Q���z��76A�9:�:�w�f�<5n7��/i�u7��([yO��%���ҍ�bUώK��+B/Jnb����)�4�{N�[4�G�]il�$V�ZS	r�v����͕�OX���$'����yĽ�pL���@լ�D��Mӣ�ɛ��N-�YjS������a��o1˜շcI>���\����K�~w^��V�.�Wo\w{W�AlWcc-�ҳ�ul�*oo��a�Z�<�x���u�If�������d�pU�}0�i�i��~���rǫ�ce�[��b�n��GILľWd����Ky7�ܵZs]  <�*��pD�]5$ |Y[n�M%������K�RS&�gi��Ю�Z�ׁ��t�lᶻ&��N��(X}������7���2�n����p��kʚ2��s��ܖ�m��wZ͎d2<If�9��(��1W�-Z!xsW�N.�d	X&.�U����,� �9w9a���J���%����v�V��Q�x�V�<��7ԍ,[���>;u,�����>��h�p�2�j���L��J��ue5Q��j�^�:F�
��p�)v��ٚ<zޯ����A���=�6��|Tغ�t앙pTZk��v�r�j�{���{�� �{����;b�s���h��Q���RӬ�S75�9�L<�V�ݘ�5����ɬ*�&C�s�șT����J88�iV��N��4�wJ5�0�8,ug���)����עfD��uk��A������Qմ��Q_KW|��콗�z�����Uڷx-�9ʪ~#�n���գ4*�o5=�K!���%�ڰa}�S���|_sf��I<�]������uc�����ѻ��C�p/.9�MKc�CGJ�F̏M��T��� ����[|K����9���R�Oh�Fv��9Bj�y��O!��ڌ fQ���uv3P��\֭��#���\B=ܬ�p>�WR�E���Y�j��N[��C��=�8��j�̯�۴�ݽ��Y�s���n��٬_ݽ�l�S�U{�R��u1�@�[��Ʒ�S�8�<ūN�]�7���-;z��9�G��)�^�˼X��{�"=\��v}1}/�@���sr\S��1s��Ou>�L8����viʴ�멎qT��U���:]Mݺ�ˮ�C�]O{0E.�w�Puȉ'�_be��9@e��{���oksJ��v^^!�Χ����;�[� ��g���(<�U9�7SP?vƻ��M�U�E���2Z��c�Jѹ�u�dB5�)M�Qu,F�p׷�;�㧨���n�J�j�`2��j\��y�b�"����SM��C}ל^���娎�f�h��P��,+H,��|�S$�Zʤ%
��\fGT\F �N�y���.�R�կ4SO�I���/��o�t��k�7ΟC3��)[z1���3GxnD�M�SM�b|��O��"&�'&�7�.�7�]�1��|/�R�r<�n�Q�����@7�[{�4I�-^17M^��zp�>{ӛ�B��}z��(�P��-�y�6�0E��z�BU�C#{�A�ҩd��p�)8�|ksyöʏ	3�E�J
E����Y�ێb�T�}���ko����������e�U���S�Ѕ-ɏT9\wV������聗��8s�;q`BՕK�[�GYta�f�-0+�-�[MqNk!>�m��ϞEM�U�\v�|tA�l�Y��b.t�n�b�E�3j齽nCP�=v��[Kw�6�^��J��|���ں<�;/��T����z�d��4��O^� �8��2��f��Ysb�3ru$���ZfeJd]��J������w4�i�J��/�����@Ct�w����a���Ø���n����.���]k�{�b:B�	N�m|U��֢b㘸�!
t���m��۫����d�p�\|,ę����3��aRR��oH	ݒO���CY�M.���C� ��,�Mz����3��#Ǡқݘ����Y�n�:F�xH����u�䴧m����;'�V,T�jkB1��R�6�n������TCfج{�Tk���Y6��P�7�v+Y��D�X"8.�)�������Or>���˸S��u]wy�Hm�Ϙ'$���� u#�8h��X�F��c�j��]�vU�֔�\�X��b���\�q�LDޔ��OwT4[Ҷ5A�²^0� 07��Y��61�X�>-��s� �7����0F�M
�h9]�h��/�����q��V����v��M軅j%@�[ĩq�hV%� ���r��
Z��F����xTn����几��fEX�$�xj��g[��&,�z� ��G�W�u	�&����J�m��!���^^�[+��ɷ���	�y�l���׳l�pxb6+��lU�P��ס^��k�w�{`�V;�v{����{��C�^N��4��w���F"
}�ݺ .�t;-�u��f���	� ;^i��^Eݻ�Ur���5��0�B����ځ:��rx�8.���,�U����Y˜�6�i|	랪�?64`�F��>~!f�w��$�άnZf�����ޛy�O�̷��{�־N��Wǀ�B�跱����Ⱦ��>fqb�3�n��P�B���ސu
��9��Zý�h-G��꯫�������yo�Ўg�YW�r����n����9�
�h�O�ɡ�M4�Q��;��!���rh����P�O�$�p��A:�û��ݍ}� �� �־y�����1�t)K4N|Y�ȕ���3n�(6���)ݎ]�(@�s]�on��v�{%�c���e��s��}q���@����U�_�˒g\��)}|[���\��t{av�`%m�J���|��Ae�� ���}�9oX8�v]ǆ��P���Iv� ��!���@N!����9�u@:{��"����*��8�^�I^�}�5�Ӡ`�M[٘�s<���zdw���X˻��{��M�������= Ʊ�a.C�T�z�K��zM�鴦�Ւ�dƹ�C�,��}%>��#��[rq�x�����b�T�mҭ2Q��_pcl��(0�v������<m��[������/�(��Kr�V���ջ�VQou�ؙ	�7"*�y;ܷr7�U#D@�{�Z�\o*�*���_m�9d�/177~X���<�����d�l��
{z�D�wee��#늷�����6�:fj�;�G �i�i"wK:�V��*��`�w5I}c�5�I%#���g�Z��ɑm[mkFn�d�[݃�C0R�����.�`�qu֕���\���L[�f*n�Vә�ɳ��Y���տ�v���AL~����n�[�Uik,F�D[AL�6���GZ��h��Z�����Z��ʖV�F֢�sc
V�ڊQ���Wk��DEX��!Z((ʒ�VTΥ�m�*�YU9k��)keH��JԫiE�
�G\���#l�	m����k�"Ѭ-�aS5�*���U�brʩ�ɩ��KZ6w5AUs+��[F\�:������+kQm��I�Z�e�<s�j#JTTU�*-m-9lDMB�+���m[J*+Q��b������U�[Z(���ͤ�ը��%lF5���Vۭ��-گ*�Tx[[�ʈ��-Aeh���X[EZ�R2��Թ%L�(���sR��m��-h�Q������R���,�,k-�]Y�^YQ�<�0��j"6���4a����U,��
��[�j��+�X������V���Q���Mx�͂	+UTQ5H��QZ�"�֤Q��v�����wKu���[Mv���^�QK�k
ev�8M�ܼ	4��N!�q�v"
X�9��8�l�\Z6���|��<[��*���͆��w�mAY-	
�l�Zڗ[Q��XPҥ #/��[�I]��;����M )�9@Tv��wi����!o��d���*
W��r���� ��J�:L�.TGUh��Ӓ�T�6�2�~[��35�����c"�$��{�9��c��F�ʧe
�R��u���49�!a��ъ9,u�c0�}g�4.;� ��N��7E�c;z�C�"��=6�j�7�p�������MH�ӟL�w����\�_����`6m!�l�$�@����ߓ�+9�����n�[<�+�r
;���eu�g ��|�9�M���y�<�P�*�6�1�@�F��q���2�^ǓW1鎇s�^��֮r�'՞�zr�X�����E�� ��˝�3��ћ��s��\����1�o����ͮע	D����3Һ}iq�H�Of��YZ�Ώ��g@�~�&r���)L�v-�pB�Ů�(�{@R3������SY�/^レׇ*�x� ��]� � Д�m���\���ҚΔ#��nWV}<j��X�j��{ؤ��t���(��tY�/Jw�~#��[d�F��,%v ��#�Ǥ���p�1q�(��Mv���L�k��;�uG�D��:p;�,Y\�}�+��g4��сߩ�K������{
eij�����!��U/�B�D���|"�ѵz��׷���� O�����B&"��a����{��&��z�L^��=z�z=�z1�j�a�9C�Shx5�����~�]���+���#��P"�I�$��X�� �C���)���+eV<i���O穇V�ÐJGv�oݻP��UPك���|�O�ٕѾ���o�נ��e_%Iޢ�`�����;�3�S;�Eq�%��'����Q�x���Բ<��r�D�������U�r(�S�Dy�kl�lz&�}}��kݛ�j���v����ѕ�M�J�������I����~���3F�FD�u�ul��rL��w��-#_�t)5������Q�VJ�1P��LTcU���U���Gq%�K����+��r@}�M��\��0��8��@	�:Xb��dYa���uBDLu�9Rv���bf��Nm����t���t䥎�fU_��媰�0�voi &�"�`Xȼx)�fi�6Nj�3w�#Ό�0Nq�Pڼ�q�`���Ty���6x��V-}ᖐ,~:+=��2��	���*����rc�}ݭ�H��;�&�	��gT���ȗ/�R�y��^~brJ��b���>{��
�ȶ ���Ί�s5��F[�-F�f�s�}�u��[���wE�>��A�rê�^�(�e�@!�N-�{�*����,�:���|�؝�í�%�8��q�u���2S��k�}l��}j��<%�·&u�[�g�r̉M9kvo��Î?<ԭ���2�Ћí⿯��G�
����.�`��p��������uD�&y���\Vt�T3i��0_E�Ƨ��.ۖ~�{<��X8��y��bn����A���*kx���	C�m,(Y�c8/Lrr��*���P�F䜳�7�=���1o�s1��_:�s�[���6��%u�9V��K�N���^����f�C.�83�QW� %4�X������k���F�$j���C!��u�h��'vq�H�V��@�E`6)WT��THWd�����L����C��/d�����x�%����0��:=�1�8W�]N���l�/�������i�! �$�����P��FglÁ^���9�Ns.LGkypj-M9 \u	�f�;�j�,�cw�3"9�a$޸�h������u�2�e�y��H>�s�ݳ������T� �A>8K �֙���U�=R���k�"\*�P«:(��*�7�Q]������з�*+��篅9��Ր����b:��)2�-�}z�^���<LMr�����$B
!jw����! �w�l8������K�9��1�c���"�י���>��x6��;,X���!�mP��&&br���!�ޱ���|��q�`��N��z�T1_�MeqY�;�)�+�WrE���]���ٛ���:��ۧa���U{ߋ�����g�ׄ�q[�>���������!�n����s��Έx�j��@Ȏn�672~�o(ᶤ�(82�r��2#�T^c�gi���N��#�Vj�)j�3�Q��堯��F��Ցl��1�"�,��:{n���zgFv��+�ҽ)Zc4K S����ڐ��:��*|c"���oo�g=�F;%B�e_6�hEé��1�jQB��qɖ!^̄6��oN�se�N�u}�^�ŀ]�pn�t����#���er�(��|��Vy�BF�u�7U�o���>����#9��م���x�5KLs��CB��C�S�Dm�@R����@e*����J���śZ�zo:��.#�,�^�δ�N�s�Zz��e������W���Ʀ꛶��>��k; ~��Y������n�����d�߂�@�k����r�KTu�flS�T+I��QWp�� �A��Ԯ�E6�k%���Nw	���J�<��K-�%�
ډ�ԑ��\j������4�睱�t�VF�H6"�E�( ��K3!Pz8]gU8�U{��$M�zXcF���9¤�@��!o��:(i��F
hT���)C�����V�NC����B�%������g��{\T���wN����koK.n� f���m(����ci`�[U2bb����\c  �#�l�	]�������0��prk�Iĕw��;�D�l��$�bؘ��մtC�a��i��o��WC�Kλs&�w�\��� 5�����ʢ��������l�Ҵ�<"Ƃ���M!��+'t������H��N��E���'t�,F�a���+�g�q�[��U��7�����^�){�8;z]���`3�E7	�hy�7��j%�F.�b�ڌ���n�k�w�(�s��Tf�5H�R���NXxTͶ{̆(���1���X��1�Vd��s�%��F�J0N� C��@/������|�l����wKPDg�,\�F��� g���;����ն��j���tS��w���ʺ�f�t�*[��V��W1qp�b`�Tfm*I�T%�Ǽv�;[��v9,��X�X}E�ͮ���e����4tj�Bz��t�k���}���V����
�z7P�S43oEw�C|��l6+�O<�P��"<*�g0(g)�z�(cswN���է���B4�\�,}+���cح	��kW��W��P�2�/G����ؚ�G(%���X�<�k�x�Na�,F��(h��[Zv�X:��v۰�J�'���T�_|SI��_ݮ�U��M��\sq�p��;S.�e���] B&@ؼ�_E�e��y���7D8��X��a�ګ�P6WC=��9|Tۯ�#��WL����:�
��~�$�=z���=�����S��iO"�>�B)����ϲ4�|w�3�<� ��Q�*��B�-��;��?4h�e�U!
��H\a��2�u}Q�
T��r�k����U9��o<��ΞF�c�^�3�����*�bo�~��r}���U��=��=�QV��'o5#����=���S�"`7R���_A�?�����k�h9\�;�n��+ã;8���ꆺ��.s���/(�o.�֪��k�?!������F�ᄬ��;�6+5jf�WW8]N�ݮ�Q\���͆����Ѹon�-��@Ύp��
�X\k�ҟ2>�����١��̾�a`�<0��{z�����L�C8��X��|�+j�'L�}�)ӗ$ꇣ�%��M>��Ö�\�-�-j�­.<j�$��ť	C*�\�ԔW�����2��
��f?==�WY���K��B�����n5�WO��/<�;�K�gKU�ݴ��\��~��DaA���d�p�0��#��:�.����*|�k�EB�M��Ϲ�ӷ�_Z��5�k�r���/�WWS"K#�,"T���ZUB�3���v���ׄ�u����O�h��f(���̿/�4ć�qLz T#�J��|�23C�#�tw)=Q�6����2)��qk>>@m�J���Vϭy�Vj����4��y����q�.�';����M�+rP�{~s����n*��+沈�7T��`���'g�%�A�p����r�\��T��L5�N�����c�ۤ��yo��t0j��u ?Vyj�:4&���=����XjTK�0��\�#d���:dJ�l�m�h��݄n�O�G��݊F%"*�e�9UУCZ.cpMf��k�TK��곥���*ܾ1p���P�w1 BNȩu��(CWX�|x�:�a�GUVܥ�P��<9<�^U?-�7;jZ 5��r�)d�7�՜��h1�ɉZu�)�?K��rﮮ���ީAS��OkWd�+:����t��zA���4�*�Z���-�7��û:��d�v:;���9�;��[rw��h$_z����6 <�y��w{c}�㗮2e�"�;�en�;#��+����v��ThM�AU�>=d�ܟ�K����Ӏ�[���	�$GD��S
g"ehZ��_Vt�(����j���ʉ
��������y�>����Ǜ&�B[�_U�!�{�n�s3���h���*��V����n&���ɴr�EZ����X�\,�C���|#���r9�Nb��D�3��A��4�Fs1i��t*�3}�3�}i�J����xfQ�ts��'V�jC�BE�y��ٵ�ś,��.��X�������ӗ򎽖�}�?+E�<+�/6OuxW������G�&�������Z[��ݗX��8��7j�f�#���a�AT�Ʈژ/ �󫭽�T�i�#EBuX3G_��q�XnL1����ן�`;N^n�=�]7���=QeVDz�b3��il�6�k��n�G&0W���m[�k�0WMO˙�`�U��?9{�����pM��7��~�Q�ӜW��{��9�+R�r�zb���)�b�ŕ��L�Kv��JW��㽆���x�T7H�rT7Ձ�����Y���Bvec��[O��@��'n�UN$��:kN�9��U���G���A�h��N�!��b<���w�.ד�+1�&��K���(��w�V)�7:m /����;[{�{��'�M`��23���4�0�x��&(F�N|6�'���*��#���/Omu�����Uٞ�|�z�i��Rh���Ce�J��B����^ڄ��k�c��~u ���d��u�G����a�.!7A��Lp=���"C�:<��ڪ(�5l�?j��U�c;8v9�-�Gӽ��r�/�n�NP��6��ꠍb�!
/��Ј���Pv�S�sYle�w��*�1Vxm0*���c�)�GD`l��.J1)��-nS�0ַ������xD��Q2�XB0�vLl�Y_uGL6x[{\T��:jш�\]��) ڛ��ʒc�Į7�T�O�t;6J�`��z��_�e������\��;u�le�N�����Q�rb��Ӓ����>ׂV�W
U��1�{[G9NJ��m�8P��e)�����墶}\� 5׽p���VK���G<��S���|0�V�	Jm��������J��!��=�	]���
��E<3��=�����=4ஷy�sj������䫴�˶��u��q�z��V�����OBf��hv�6밎�,k�f�u��8��gln�)F�*�*W�;��{#������dY>W�r�h���-Q�t�ޣ�uuu�V�ˍ�;6{���/
uC� �s�;wF?
�>TN?��u��XT�[|ZW�\l���F�Dr���Lb�QGJs8@{DG��K��'����0S'#�%X�pa�68F2����@LF���29�DV5Jzq�������-p�~v��g7,�,�w�pO�,�Ɗ��l�!��b
D
���ϣ�G:���R��]>��ǆ=�{,;7�7��r%�A[O<��=j�)� =i02�G[.�3˨#�z��W�^�n�E|�e����WϺ��K�WT�um��O�z�i��-	�bǐ�:��B��V��a�ıM|ܡ��׆�Z�
S6=��S=+�4b�le����^W=��؇�#�f�����r�C)�h�Zb�9�z���ĩB6�f=����IT�{n�:������r���<�~[���w�XB�T��Ɯ�������-^��Y}@>��ȩ� ����U�m!�\������s `��渧:7���e"�hR+0�+�h��2��'mƵ���Ww[yH ����]'�W����myN�g[ *���맙!���x�mv�e:(V���Zuֵ��3�}Q�l~r;:���y�U �����y��c�(.�bn>kU��FZ򔄚}���ǉ���qx^'NAW���ӌK�U��϶�d̫�K�@�J,z,��٢n�� �)-�մ��C(_?K��v��mv�K+�JfV��^�JV��ԋ�u!9�k�XF :�,���2�N���)5��p���9(�n���xa���~�ϑ���7�����۸O�.�T�&�|^����މ�:�c��'��
+�$p��X�R���z�Nעv��9�e��ssp���="v�J.vN�d���B�7YښJ�^�֐�/^"Ƽ-�Jp��߶!H�<{�rZ2���$��ɕ/��x\f֟�ϏiON��'�{����9x�5`�=�'�%�̀�M�.�r�e�V9��it5�D��^����Ӯ�S$J5b�Ũ^��>���>�]+�d�%{����i�p{�Eȃ9�
��B�ى�S��䬎T��t�Yyp�{��|r�r&����~�x��ɜ,f�$�߽��� պ��ؤ��$u��1�q�앗�G��N�L��v�������>�����͓�$Oo�o5���C����u<���U�i'nQ����u��b��vj�@�anc�tބ:p;�u���0�Y�F=+7ܞj�SZ����=��3@�ӹi�%�S���k���H�i���ɦyv:�{7�ѷ��x Ǟ頵)�J�̭Ϯ1/j6���YZ6���r�n��a9�a]_d/����I/'�=τI�}�/���|9]�ȟ���?��U�xV�df��k���6����k��7&x��`~7G?�}�i��|����β;��i��惕q��o������̾���GM��>���ɚ�+ۜ��K��}Ʀ�[�^��S���1���R|�a�8��l�l,��lw	kd+X_aZR�Vf��-K�8�<�d}[f�Nu��[ժ�!v���c���7r�tm^�-�l�Ǡ���>.�ãC�c3i�A��{�YR=O�B�;sC�.\�W�䜳f��6��Y�6�
ɮ��U��sl��u籛��Ou���e�TU$��t��ξ��p�i�|
W�[�Dk�rP�T��� ��5K	V'v��ѝY(d
��r����{;�V���'[�i|hvY�*�N�:l6^l����"���K��/o\���ȫ�
FR�cmp/����q|5��E\�]3�i�I��-:��������c���`�@$�R��a�^ŲJ�+�{���҇lP�;�.��xYX��ct"=\[�;�v�0쯛Sٸ�J��h��g�.�
��}]֦vm[����|����gح.����l�'�r�,! O�ڶ�%lJ��[eV�h��EVR�Z9m�KJ
=���sAm(�J�,�E���F�S��:%V5�-�ͩ�5.
�QXE3u��F��cmռL�kV���-h��Yu�Kmj�U��+FѵZ�TQ�����b�R�PJ�UF

"�"*!hRҋ�U��F�KmX�J�
*�Yu��kh���խ�WV��6��Rұm�k*"��lh6����
�� ���m�eX�[A[M�V�[ED���Q�أ"5����J�s��X�#i`֣-�m�����Q�[H���P�V�U�D�V(�5+�͕�F��`���0��RT)iEKj"��Z�Z�1V�6��([�kUEFs�"-���W������AC#j��V5��%E��¸�[Q�
���Km�+*ѵ�*�*����E����E�P���d�U�|.��§&S{9^�w��:Xx��!/��
�i���C&�Ɂ3�EZ�[�x��|	$t��j4H˧k{k���T����
_����1PU86�v�̓�C?P��}O��t�Ĭ�r���:O*>�eC�=C�������������x�:;��R||O2;���:�v	��q���Z�G�"8Dh� Gރ����g�K��z��d���hz礂���C�Y*�p�U���v��S��q�Y�״=N�zϩ�}�3<C�d?0��� �OY_;�~?��ޱ_�''�M΀�����>���}==� �Ǵ���~'~B�{Iߞ���*��~��d+���3�,�gS�4�
����Y2A�gO�*�9{C�l��?Y7�E�_7�z2]��K9�z�C��">b?&ovg�>������t�U�^��q'�VSw�:�@�2<a����?'L���?w������2�$�+>�9�*J���n�������Qg2��C���gսǺ��(1�"OKb�Y<r�����x�~��l�RW��9��<a��N�����I��3>y֓���z�/�x T����:g��<@��=����"�N4�}��DX�DQ:C������>�ҳ�J��u�;I_��L��ė�P�¤�
��ٿw�|����%��8¾�$w�N%d����{��X��I����7�޷�n~���N�U \p�G�#�=�{�y2:a���!��&g�ẋ��r�
��9:�C�|C$����Y��&C��C��O�T��RX_���>�T��S��q�큐����qu7��s(�7��[��=��"S=2{���:d���|�JΕ���{ҡ�C�����`�÷$���8�Y�O�l=C�YΨ|N$��I��C>0���~x��VJ��WvF���c(z���U^��>�@��~rxϊ��T���8��+��&�=��� }J���9%k>�V��+'�+'7��J�2v��Ϻ�%~�϶~�Ă���>��N��rw���`�y$�C}8Cyo���>�#�>����-C���v��
����cƳ�=C'�O�{�H*�l*u=����7�y����t���Hd����7�{�C�K���rɒx�g�1�|�߀��ٿyt��.wf��.O���	/F��ۗ��c�W����=���2��r�,�f!�MKA���9�{����N#���G\�ڶڊ�%לN�z�=�y�D+��2&=�u���-uc}�<z����צ>W}Ӕw�z��7cͻ�ֈu`)Լ���RG��HUAU��6j�G�Ă��O8���8l� �������W y���2v��g������2=��	�Ad���8�O�fw�^�Tx��"Bzy��Ͻ��W�9ӷ1S�n>""8G�!�1�B><I?!���$��	�����~�fI����ON��C�<d�Y��4��Ї�\����|�vv4�̍���c�d����"�I��J���fv�O�Y�Ĭ��:柟d��,=g�%a���8��+�z����>yC�L�Ŀ;�d����Y���'n�U4f~0����@M���U���^�=>���$��7�I״�Ago�)�3*O�����eH/��S���*T:>Xz��7�O���Aa�����t�_��O����:�׾C���#�>�B����%{O�>�;�Ă�䗣�~�C���Y�|�o1���6�YXx���L�*VJ��`d�����i�~a\ï�8��z���������N�� �ز����Ϙ����c���2AC��4�!�v�d��3��Ago�7��� �ğP���~s�O��O���t���:>�q�a_<�3X��~C����Փ��%I|��w���VmO�En�St�r�����>��G�	<B�d�����z��!��i�Ag�|���$�
������Rv�O�{��>�C���~�2VN�y�'L��L�}�H�!�J�=�?s���u�@.���OKr���>b ��=~��I�9:�E�Ƴ�%~k'�O�bȤ�
�����z���������{N$�����d��x{I� �����_`��	iB{�1�l��G���Ͽ������8�@�S�z�W�񝡓�}Xq ���:��Rd2A�[�?0�Yĕ�l<N!�J�O���q ��oؾ�'�W�<Ǭ�|���$}��b>��G�#�ja>�����c���_�?~���Ь�%J���޸���}�C���l+��u����f��_��Ag�~g��X?$�8ua�8����_,3�
���!��t��T�P����$]�/^����+��`��wF�����n�'];���u� $:�GtjPJǵܿ�pC�S��C�u�$�Rec��퐂�K��'WC7~?Jr���N������e��N���z����vq��'�K�պ+yhWөev��DE*��v��}}/�
������{���κ�P�%C��~�Y*����d�Xu��Ğ�{�~O�����z��������$x�a��OP����ed��G�"�����N�8ט����,�} k�����~~����VO)�q��Rd��OYU��^�����}B����N!�J���S"��Y�^���
v��ζ��+�O�=N�� ��#q�y
��>Û�Cۼp��BG�|�`{��v�{�fd��@��D1��t�ω�'��1Ǥ;OP�/�߼���3<C'��� �P��9�!�����sXd2��%�� �DB�#�G��(t�}�㠝58�'
S��ykI�:>^3�K����ϴ񓖁����L�*V��p��P:?w����z�a��s�{@���3{��i�AgH~���DD�����1MI�����3�2�E�zW�IYP�;C3Ӟi9i*>�����T�'��8�?Y2Az�(xÊ��Y����
¿|����Hq%C�??�
��^�>�����Y�=���#���ç��q����A��{���糏l
��|��I��2AOo��%rO�:��qY>%I���8�|�|M�C����Vu�a�}}I�|>�fOYU�!�2L�I�����x}�x���|��f7��5X��E�G�X|eg���$������z����:0*��'��)�O�+>2_,�:׉X��>�������C5���`z�v�X���)�{��N���EHf�㤱��Q�N�d��Hd�P��<a������t��T?$���_xv�� ���ϼ�+I���:ed�_>o7Hx������}ꁙ�NVT� >IU�����N�z�����(}#�q��(�C�<L�z��}N�;Oe���$�7�*�����︆k
�����ޤ���T�f�����2G�q�VJ�����z�O�G�C��V��Re��'4�/f���;C�����;N��
ʓ�����ez>P2Nп�Vz��`T<g�Sפ��i��~�)<zI��
��%a��w�t�_>�:C׏�""�+'�I�y~����*��3~6�+lo�m�8���qh�bHT�dA2߄qܒ��Wh���yF�p��#���r��e�:��yd�����Ey	�_:�Y}Ic}���7�T�-���Mُ�=�vZɻ�XPGg��l�8��]֊���}�#Ca�>����>3�����Y3'l�ϩ��I�*OS��q�<d����5��Ȳz�XQ�>���ο���g��rdd쫭}J�bR[��H˗�+�C����G�	L�4:=�1�{Ӻb���b���9����۝x5���yRp�̘ʾˢ}
K<�j�H���&&)un��&̸D�y��#��:ۖ��5gp8\��;�b)@��w ��� �7a_p��O2<�k�f�ߓ��6Wt�@��fF��46.�o���vl���|�h���-]9=Xn��,!����t��#�V�m�ⵞ�x�ְ/�kF�a�<균�:�T<i��T\���SRI�����ޔ���\ض��dJWrQ���:����V��f��@LF���3�
��s�f�ڱO^�(1+}{��4l׫��e#��j�1_YzP�'b� �Ѐ��@��{<xpP7m�7P]�|��(��>c��˵��0k=��{�G���_X�i� e�lr� c.1d��ug^��@1�ޝ��|"���B�鯒�:s~^x0�C�ϭ��
��;�*aT�O���.�o2^�{�����ƹ %]�&D��t�_a�@��肝2���Ԓ�{��&�X�^{ �4s�7JR�6� ���D�m�7���o���G�[�c�
�]��p*W�gëЅ��~ٝ����'���r��W�;8g�G�����nS�u9#�1��+d�0�e��b5�/^T�[�r�'��Z ��PH�tky��+S*5�t�?U�\�Q��0��2���7�2�N������@�e�ԁ�.u_M�&h��`&��qv����U���1w������ʒ���
���y�f���b�M�\Ͼ=��n ���Ӿ<�
U���ok�ua���w�M�`i�V���o������?$@�
�Hce*D�F��&T�38�!E�M�����-V�g���N%.ꑢ
62�n}d##�M}]4+�)�A|pj�z?S}��� &�T����}���w�l�wX'D`���t@��$5!�7�����^g!�F�6��Szq��wN��rj��=L_��qrs�y@swDm�� Tt�����^�͚'�`��5��OЇ��"8,?[s� !k��ar�U1��͚U7�y@.����/d�ls����Gh�>��`ț��n�y�ሺ,x<>�\'���:�s5�T
l��[v�q���-j��}(�r5�{�} �_��fu5y�'��0&Vbf=�T��G�(B��o�a���B6�`=�*rSVj�:�G�*pRv[V�\!a�d;2��bo��A�)�ڴ��P���텷��")
��Uɗ�o�^��d���5�;t���Wf�}j���g,?� ��	u`b���SAF�9)��x���2�.��֦CP���J7p�;0��=��/'F���xcj��%e�o'���;�a��k��g0Ȩn@��'Lira��C.2��̢1WJ����$����U1T�k�m.vGd���ߝ��)��#B}'>�V��������U'��mlR�j��<�e}��o�}�_�+���@�lo���ע��O�ؚ��d�;�V�{:���z(y���1��J�ϭ/i��9U��l�q���m��%B�O,�J-�.��U>P��2޻�~�����C��I�*���J�8����<'�W��炑h��'oS�G�Ndb��k�՗��
cm�����06R�*��+6��`u�����XӼ5������;u�*f\0(�/�	d�6K����R<�嚐|���
Uе�3�h�����/���I�G#\������j�������0�	��q@!���n�o(��v�~���PvJ��4|������h��N�c�G>�m{U2�Y	�MU�wN^w7��������:`a�3VҐ��Al�$԰�C
�U;v��p���q\t�*h�S焙w81Vdޠ�ݪ�*��$����iY����/7 �O������b��f�=��T+3��i� �A��+��S����Z��c�����u�W�����65L�r��/⧰ňL�ܺ�72��"pq�Nb6�T����kթ���I���w"b~����Kj$V)cv6P΃C�ճ	��T��(�1U\�ոԧqɂ�������ߴ��}o	���7g�9�������ugL�K�����9A#{��fE��N�1f������k+�'����{�6�;�K��9J�|]�n�
d�Q���'U��#�6o�lL!�2��q&���(Č]�4��������M�i���F���N��F��d��p7*~�o(��I�sOd��9�WRS���V�%��h�(Bߢ��ϯ��)��UN����_��A�-E�U�Iмǹ��b�`�Q�9��E0a�{��>Z��ث�_D��_�1Q�@�{R�u�,�zbst9h��J[�݋N�4[׶�gܶ����%���IWCZ����ʿ +�bC���X�0�|y�/�o�P��A ��rԦ�A�*8NzB���>U{y<��ږ�����[|���w�;�������ٛ� *9�Y�cm�[�����Pu.�eM��Ȇ�T|:c���H渵�G�ö��J�Ӿu8�5Z�e<�՟������'py��z;�ɪ�6S��k�����)M���~�~���8s%'��<}A���3ڐ튭	�j������r���,`ڮw��DVm{�Ǟ�ڐ`(\�֞��B:q�3�:���*�Rgx{ Ć�F��W�-9~c����IV;b����g0)�8�܊�Ψ-���ܧY�O|��? �-Ƭp�;��'i�q���|0F	�iT8��9��fŜz���h��G�������-��9�S^;����T)�ǃy<T�%����V�v�8�d�;15K&��%� pY2����q�߁A�ei(oa��
&D�͌�Vm')b�n�7�s���Э5O���m����S�Yg	������4qH/pk���/<��`�Ѧ-��g �� ژ�Sy`�ބ G�E}��������&��6�>��81�PoD­I�ßkT��P�Kq�k�S-xU�t5����ճv��B{���8�
uk��]a��9X��5Lb�ME7�<h�T�O�'׹ww+�Q붊\I�FD�n�Ɠ��Z[��z�:��á�᠄�W��g��a]�wrb��J��ɮ�ۭ�|�CnM��u3w���{�m������9�փO��� �ky�!��-ަ{,aǅI����l�On{��#�'bn0��0� ��#�^��qh�lX�ǅ:�,^>*�q�1��*"��3ҧ;&bl=�-���c�O��-�Zد}�y8>���[\ ��o��< и��y�[CUH��@x���qN���w9��-W��؟{�=�k�Yȱ��j��=�P����졗��� �h�Z�c=Z��g���m7y�O{� �+"d���ڵ�����L�:EŌ�-�4��.8�f�e.vɼsv�"�x`_kʞ7v�1jg��k�,<�`ӷ2d��j@ŵd��Ŕ9��4�����g��sT�Z��e�$�\��uK������S�E}+�O���_���7�r��\75zջ|Rhd�}<a�������]�U`&���|y�>�lpý����7�\OK5k_.',�u mD,���
������%@YuR)J'p����E�������Q��lP��Ӥ�'�d�)�M�74�F>�s��B�u�J��_30脪�2�X�޷O�V�.�r�l>{���w$�ޚ�ȼ!�
ٲ��ݯ{瑹�b�̘�&��Vs����
�!Ԯ�%��r���W�{u���;��h�,�x3�1�/��\����ƾK��]
1+�Ck�:���ԭ	
�oj�0_"��������@m͠{f�3��?���ﾪ�B^���hg�o�&:��DL�d5:rvF���tE�\��e��As�x�n2�����ʝ����(|�M���<���V�M_�����qrK���!�[��(MF���V�O�rg���� ��(�S�y����xs~a��D¨�j��`���R�0L�VC���g��'=6mV���5�]&��j��|-�p������p���yV���gt��tŦ�����q�k�K��C�!���2�׸�ҏ�,�ܘzuv&`=y=����ElNruu�C�����I�Ha�\+�}x >�'X��T��⁷Y=B�gbP/q�3gs������s҇)�`c��g0ȯ��0T4$銈.@�7�䡒���Q�:��&{7&����hfF�۬b�@��e)��H��w���p̧��X���0����RhΥ�b�6F�a!A�b����caAن2�7�X+'��DW1��(~��s�����Ö�ȇxf��)]N9j�}��Z��!Qs8���/�ΙK����T���� �����9�:���J
���]_sS¬C���X�`*���R*͒��Ҁ4I�k{2�ۤt���!�4g9�����cKC834�J�ހ��\�Ze1o*�]�'{sx�:r�Y7��ו����-k#;��hك���n�ZqHay尥f[�|��4ek�ć:��=���>^>�7e�������s��N��eBۧ�a��'^PtUd��c"s��Ȉ���P޹gicO $W����d��f.]�>�3����E�9\6�ę��$&�h]1z�[[.�N��8�.%g3���C��u[8�thn�w�Q��'$��������/1�����xA��\�-`v����ϨPQ�v֑]B���[�q��p�G�u�{���oE�f�;6��r�Z�V����{/3�J�e�w�_fƷd�7�<��Q�7'�1��~'}�4B�{l����
�����(u�i��v<�3�4SI���m6�.H#X~�2���/3�j(��PYc�Լ(��Ňb�q�y���y�����η�#�s�;#���+��^j�+��ӽ��a{�NZ�m��>}�񞰚q�'����r��\��t,t���"�z��wMR�a��y���M��R�1r�^��s�56��h�v~��������E�h�Fh̔M�|��tS�+�6IP���U��$��'A��g�5Y�d5�)�J�g���Wb��e�9�U�WckxȯH�R��wd�33x[�{Yb����; �t���$���OS>ŝ��<�i��h���=�
0��9��E��c�C,	����3TͽP£	n.�T�Hk������.�g���Z��O��Э�aH+^!�+�5��<�J��t.��T;K��K;��t�]�r:ܡ��[��f�԰�͹+@ZYޥ7(q�B�Ze�T�lF��1���6�q�l-���C�ິ7��Җ�Z���+�#äz�~�FY�������,�s�V���{秤�;��_tH�wD}��'���7���wJu�˞A�ܚ���gkj[����{n��[�9�7ϐ��fGg��ãxlF�;'��#.�M��3g���)Z8q�z�w=�Alͫ�?�]�QΕ�P�F�P�r�7����>����hD���H�G�W�Q����r�T�yg�7�@T7��ͯ{�\�=�,�}����\���+�y`� ���MC�c�&��a��.��c�k�X��A9��{���&n�d�]S�,"���Ai����KP;1H�k����g8�5���������1��A�ŽJb�w�B5�1��r���}4)��N�v�N�� ��
z	�w��]u]��6n�<+� 
��E�	4:�r�9DJótb�e��[7L>P����T\�:t���p����#]XgB��%����e�η�_EF��ۮ6��V�H���&���o�����8�EMeUZ�j#Z�f�6l�ԱfJ�UZ6,�Kh��U��m���[p�2s�+ĭ�b��ʅ��ʜ�ւlMlm(�	mmu)��Q`+h���6��p֊1�cl��f�%�E��K)jѵ�'5NPQ�m�1�R��׌yL7he(�Qm�Ee5�댖�<�,�9Ղ������S"����ت*�EV3�\�[3*[f��Ymj�R�"�,Ee�V�F[V]D��R�P�kl����4imm�Q�U-�D[j#�1���UE�T�S��bjQ:�duZ�Fڶ�R��	*�T�cD�2,\�k^\�m�#Q^Zŭ�V)����e,D!]jZ4�J�����abd�N�Ux�5�EkӇ��]V��b[�Um��m�)�b�k�[U[AQI�]�j�UUB��a3TV�T���e�֯����2��y���X�*��jRڱ`�PW�c�T@��(Q&�C����;�-���s@����£�\լ�W���I���v+��hnG������T�k�����J��t�{��T*�/}U��}U��s���,�nceO����T�S�*��Ǆ���'��q��kKس�A�[j�԰
j����!�M�Ȣ�u�L.��Ud���|�.U]�|�]��Ȯ ����)�7��`�6����G\U1Acs�Z-�T1=2\H��-��ՑN�6Q@︢,����(�/g�[�P�����E:H���!3ps+��:ʉF�g&v�m���nH����'��j͸��h�!���|j������c� ��®1吕����5]{z��1�EUԝ��
0x,���)b�|T�� �m۞�1pT�eN���C�X���nW1;�*����O�@z���4~�Mx���mD��R���C
���Ռ��ҧF� �;5<���wH�"��������~Ӷ���o	�S�]��ޣ��� z�Sne��X�ȟUqb(SRm�P�:0 Rb�1d��pdߠ4����ӵ�{sIs�����.8�30Ѩ�̶3䪥��a�#�6_�a�ς�}�������[�X�>y�����^����z�-ޚz�f��18�b��ء{%�������c�Xomj�CWp�*+�i�[�;�4w���ɵM�W�sԝ%�S�<��%�r�iȮ�Y�*i��oF<��%����$.p��g�}_U}�@�I��i��B���~�����'��oK�y�j��@��<k�U_Ts{gL�"�k�YF��=N�7�%
I���*r�e�?�����3�V�N���_���o���R{�\]�`F��෥o�+VӘa��
����Q;</Ɛʾ@_b#׿gZ f������(	�ގ`�fm�h���Y��𶌾9&,GW�0���֨�/T��u�g.��
89�e�#��Y�8k��kN>ul���������Wk��j;���:�xt�[b��p{��v�H��L��s�ʧ�R��r���tƋ�KVpogDr�U\)�Z6�9�d%U��	�ծ�������N�'�>^��bB�[P�r��4��iL�
m�9E`oNt(P����Yø�W� ྠ�UH���@U��`C�C�����w�d8B�wmxD�E�'�蕊�q�Pn�$5��3�B0�vJ{?-�L><1�Zj�kV�9G&��Б��7-���n��W��&�a�h�L�1��vl��2��Pk�~����]o`}��H�ezڌ�ץ�Q�m�|T�bJ��<G�S&��f��̳)�E�ϫ����Z���X�@�V�Xi^hN�F�=Onn��ո�{�M��Q��9Y����D�r7�nNS��rr�d���%�t���7&�C}9b�֙�]��-V������U�=������:����N��l�}mdVe�[�}�n��]M
��v8��%�yy$����u�;�B9#,l7�l�A{LAF(��Xj��3v��_|���/�YtÆ$�b��DO}�Yj�����`v�V�� j�W�sT�b����,M�����T^W��i��cL��L�r�_W��-���h`�����.����Gy��]��<Ip�6�F�������*�p1���6�g��/|êC�wd�4���-��ؤ1{=�+{!�S�p
���r�
��҅��b�l�9�:�2�7\��8��4�"�w��ӁW�n|������^B�_1pحO=�Z�i$L��ŋ�N_0����H� G#L�$�SY\(\c�_T%�t�K�zd!zo����Ngv���c�Wόk5TF��T.猘�m�Q�[(`�yS������
�<��e���͕�z��� �zWKKΡ�o)��(;;�gF}NcG
��Ea٭vB*�үyc�1:��X�K�c��7*�-z��g%͏�~�+`��MaG�Vz ��[36S�F:�@ގ��*���9{���٬W�;8Y�G�݋���3����/`��~�5y�|����k�m�^�o���|n�����>��Q'�˦�j��	P�W(A؄��q{O	Uih���>���0JA�q[x�B�B��+L�t�scR�B��ο� h�#j�vn:t��0�
���'��/4C�e�Ů��2��*	[��q���Y k���U{�ʽjb
��������.�C�"n0������������aK�����"îz���+�Ɨª�S�z������Ө�[�̜���GVvipKgsg�:�j��l�yZbvF��RF|�$T5A�  Lo�]T�G&	}�;����G�zR9��@Vw�W��J��#2y����A��g9ַ�t�i�8��uy`��蛦"�#��R���WM
��nc ����yMW�a�u#�7o'���6�I�\ER�u�*�X��"�p�u���k��j/��6�c*�+(a��73æ�%a�3��B� �m�KND���M��g,�g֫�]Vr�RX7|H�A+��yd}��L�ֲ(hXhh{�E�e�N�uA�C���^��}� g� ����l�1c�������n	�{�]���;R
���.��A��ha�)�A���S�]N�ff��T����o��b�̍� �X�k�;{B*�*�o��q�U�H��`m���eR�3ZI���&�`��J��ȹ�NPK�t�XQj$ʖ)e�}��G�s�CۼHy�7NO��  ��}���q��:m��LN���u��� 6�Po�xl��wɂ����b:7�*5���gDE��T��VE�-�8��¡�u�f4"��$�ʐvh�J�iJ�!q=���fp�'�j��4|�"ά@���B-&�����`�
X��]�7�E�E��Ȝ��X팘�����FL�+:dm.����"��������t���)���`SU\�dZ~�����p�yJn �k<xKJ�:���Yϔ���T�����ŭ�t��3�%��ҧ���%{�>S�ʫ���J]��q�ޜ�n�����:�U|�Gڶ�_�UGPX��և��T1t�P %=e ��M�*���++~�z���l�ل�����')��S�8:2�!e��
,����V����5�ۮU��p`�r4�:�MJ�|d�״��p��;�(�[�8T=���{U�����Pb�H*d�)��
򫉟�L1��
��s˯��T��m��ˆ�R�%-���4�]ë50aU&�����p��>���a�5x��&�{�8𡐠*������.ʝ����]�B���]���ѽ6�4�<	&�Ջ}��-Cl�H7H˽�B��g��o	�z+i��/��,��8 +ج�fVQ�mv+Bs�_}��U��g�V������*�s�Qu9?"�X]�mR��5�i>�H_�<#
{��۷ׅrU�DX��=�%,H�9��%K5��US��un#+I�~�9%�INe6�nE��8+t�[z#��V�e�D��j�}���c8N %�E�R�n|g��X�44��r��_>��Lc[NN��>Ɇ�f��!�g���d��a�9Se�����|:%j�U�����d����F�c�[��qZϰ�x���f�:y���29�(�@ܩ����ֶ��=�\kSuG��*@�%���.��z��v[�������mG7���t�lي�Nn*}�aXN��>�9�'6M�� ]���W��;�������cA�lr{@yN禯2��� 9T�}���3.)�s��+��e+�s+���P�q��������M�%�U7#y[Ө�����+룼��,��*k�.s~��Q�'���2&^�j��yʜ� -."�P�s�W�5��NS1��ڹ�j���{�P�y��� Huy�^)~��4�������B�[y���6U�H7q,'pR�J4�Mԧ�I̥Z�^�
݃/6�t�Br�{l�>��VVz%��=/��R�/L��}ݼ��~�N1�8�I�v���<�LWt�oV�*[�G�+�
(7�I���}U�|��f{������U*�\�!3ѫjEa�S.9����
��B�r�4؞�O�<qv�A�Rْ7>�H
��ы0=i�F3�*\H�b+�+Tt�����+dEָWhk��G��ǐn�$5��;dp�^���g�Qn�9K1�c}e��j+啩��C5mqR�=:4b0�L��� hKb�Q�'C�pJ�QJ̅Ө��jX,k�:�1q
�����	ހ��,�̗Ӌ���[�n��҈v�z���h�p6����b�ڶC�bB�0 �����6f�spËA��[԰}"�˨��U�t=/HC4�	|��f�@4s�Y@Ed�@�Vv:%�
�um��U�IT�1��-�y�^Z�'Xxy�Ճ>�F0�D�{��fZ���q �h����MՄ��jFXo�/�T�:�1�UE�#Y�f��N�\\�fS��L3}ܥ@�����-�mm�1m ��G�mW=g�а����F��t�^��K�Z�(
p���x�V���5{�J��ݓ_�4��F˫��8􎥏OI��pj����,6y��&�7z��BѪ�PQ�JG$ף*�o��k���(�gX������#��nC��Kù�N��::�a����)���}+�q���u��&?W�G��˫�N�jx�d�i�+V�\��<W�o`���]Ĳ,�����Y�n�>�E������y�7�c@�k�z��i�����k+��zkꄰV�ϥ֍=3�:8�x%�	;�`g�[U��Y��Q��r7 �2����7�9�;s�h��P�Q�����8�F����9����^��+�Sp3d+ɝ?TY��o�SAX,<6ܦW�s2jYN�NS��{W3\�Z�ޯxjVy�@.:��
1&��Hq{O	�L�w��P6S8 �������Q��G#Q����J�p�q�#m��d% vkp�p=[��
�g3���O���L��u
����ˇ00�V������$y̨r"�F��J�Py�Vm+پ>�SO[�Å!�ծ����Ѕ*u�r�A��Fr�Cr�G-2��y��[��Ps��R4��89�����������P�T6C��W:�'��c��A�#�4,�0���ݱ���(80te>?K�g >9��Xy5_s��b�.s������`�k�����VQ�7}�y��pս�]��[o�k�ed�[;�@�(�f�@�^�k��w1����㜭lR�ެ�3�7X#Ǧ��W&X֥�β
S�T_o'�?I�y�t�o��2cå���Au�'v�V��諭����p�nr�� %0 �l��.n���$O���"��/L�	.V�V����9����~����A?cW�?#��6����B̘����a8�,c
�f8��d���Ko�A�#f+���"b�в�"�{��މ��*�0¼�zuD�G=I�u�B��M^u�/�Åv�8MJx�}���kc�zG���2W�:rR�]d+Xm9�����d�'�u>B��&0`�9;��.��qʪ����!����1*����\s�H�=�=h�f��b�uG�1�kj0�81L��_!-�vE���3�B6 ����6���{u/�{���,V����1t���S�+i�����u�y��r���^z0��,��Ӕ?�h��p��e/[�v��j��	�9���=u�[[�՞�R�z ����{�uA�Ƣ{�2�S�~��0��A"��	��e&T�pr��t�KN�J��^�V������WqNX�U��Q�����)r���B��g-J����ӹp� �=�̋����D��u���g�\mfZa�ps�M�X��^yG�7���0��c���qc�4Ic�aY/�	K.-�$�(!'����!�{��j�0���bp��]3�Stf��z��d�wo����#:L���v����W�}U�	~QtS{�Ԑ�e2�j��fU/K��J��qv�����	d�9 vk��9C��T�L8�O�%�������j5}��BN�:���z'E�V�|�	��68��쥳S5�2�p`�;TȘ=/�B�vK��0�'i�nc�!2�94�����~:A�D^�\O�z�0��:���ib�|T�����C/�nz�fJ#�ݴ�H�OfwG����+�U\ꧮQu9?"�q۪T���&'�[Q"��,n���eu�� s�Y85���S��*CS ;b��%���e6��.�u�k	���7�t��5�ho�����+WOu�oFKw�$%��򚡌�8 ��b�5,v������K%�Ψg��E�=]�jO{F��c&;�t�S2ˈ������׈d����le�أw��C�p�~����t�p�jeZǊ}��⓬5z��ϵMs dstQj��u���w\�R�z��y��0J���b|.UZ�qXve_!�SO ��IU��f�Ѿ�`�ؙP�E���Gcz�ixjG݅n*�L�N ����h3k�:+��hM�G��Le��^�梨�!y�g��7�c�f/I�;p�km��F�8ڨ� G�e�E����������p�̝���$˅�J �8���������;�S�ai;�4���V�v���$�0�ܯ��m˰�R'��]��rj����Ɖ0�lO���eX�L��ú�+.�޷�������]�D����qc����	si�v�Z�7W�VF�F���)�Wk��WS�����)�R���n�v���ڻ��SP�P�,��3'1�Mj��#�ws[׵�<�.1�������!�#r:�[x�n�ʼf&�::<&�*ͪ����L]`��t~c�6l�8n��8_h0���XȘ��{�8� ��K�{�(t� �8]�v$��]�o�rz,�5����S��Sa�P����䀧�y[��ɛZS&��J�I�=ՠ��xw�xmt}��/�w������FG��s�$�CL�M�Y��I��v��Vv�v�����_������u�Z�E\�'�B��� ۽�$�Ɩ�;�{)q��Qh�E�35RȘ9]�n���4E��ftf��ecRG�;7xi�!xݲNǓ�"��9��2qE�p����̮shktV@Xѵ/w��-��4�#����AM��Zcon,E����wo��_u���oV:}�K��lx�!��g��(g���c-g`�ws�W��^�&��Y!$�9Zi(���f�H�%����wept��V�*HÎ�m�X2�=��ӽr�E���9�p��93Rئ�Y��B�S��t1>?rܵr]�q��P�2��3M����Ѿ��G�<�v6�������R(钍�4����kX:�l\7��]���&��#��oT�Yw[N�\ٹ:]5ui[=;{T��N.P��7��c�й)�+d֎��*���w��HBk��-�|hP�
`�549S�i���O�	cVf�ν`�O^� ���T�$�Sx�u
4���7#/�չ�����5��>I����=�s���Sk�Ụ�>�8�a^Prs{t2)xa�aVjPڰ8�^謞��bǗuTgu�zo{o���2�.��v#�D�q��߮{<;�-��@��ý��wR�/`�Olad�XT�Ɩ�y2�:H�٭�Qδ7-�����G�V_5�*f�7,����E��S}�=`,�sR.�];���k�Bi��[�T붻�u�^l���;˺^|S������*=�8��ALX����ٲ���ĝ�v�q���7�3G���tJ��/U�P��`��Z$%F�[���n!�k�^l����ݿ�~������
��ٱ��1
�̴iYP[j��Ȗ�S�A׎Է\*$P��lPVѶ)R�[�iU��V�XjQV�+X��#'5��b#��.�UUU�MvU���m�F����+��p5�3��<Z,D�YF("#+kTZ� �X�ʹ�ĭ:o6��6F�[m�(�U���6�GmUMB�+km�������Z�sj�[�h%���A9�8�Eu���r�f����N�����j�z�fjR��n`q2f�T�*rض����Z)"��-,�֢Ǎy�\�,��N99�ͽlu�"kN�C58��q�������Ԩʑh�T岲ǍSR�ܵ�J�I�lk�`�����*u�YQUu�d���yn�q�J�r��6����+�q�5��%�����Pڙ��YYZ�)��^rPG�7��^:s�UAKj�K��Q���T����*Us�>����34~�T}�,�5�Q%�ݨ �Z.hG9��8�K ��v��Y��x(yr�^�@�^��o��'�1lYY3�j�
��}�G�%b�-%�ν��7\�å�"��3D�3�pw��U�S���E1m���7^�}��s��i��v� �.��ܡ�����d\~�Y��V+e%]�)àL(�OM��2�FM�]�ѽ��)��\��ϟ:�7"�h�����^�ˢe&,#�f*J�WcH��n��ot� g'���W�;��8�S1�R�׽��j���Ԧ��.���iۥ{Ki����.��(��tW)XbBf�mB��ʖ�1�y9b	�sz��M��Z��pį��@R>�b�+>�����]1O�T!=Lg�T����!\'�Z���۵�덳��;~�\��K����x��pĳ�a���2��S��O�R�Z{�[ю�N|ܳƐ�v�u9_?[����.�&���-mdͦ��
��A�б��Qf�G�OИi_�|+2/&��
�l���.�Ǵ���2�+�e���;7
n:�o"��!�Z�	���bh�eZv���Nt��]JZC����֭uD����9�87�T���l����E�n�"n)&�D�f��*`���xvDN(������k��j�^שD�]]@�	��y�'�7�ݗ�e\�a�]H���ړvDF.��݃OVt�8E۳�U����j���}��RGt�I'==^���}l)��1��*��LU5�7h\Q�����,v&���J�>�~�5h�#ѽ4��|�}�O7�*�R��vQr.�f���W��|���;��f�?2�:+�[�gX1�:]\�im&<��+9���+�l6�چ�*z7�mo��eW_E��?t���M�#p_���PyE�ϣ�z/�k��\l��s_7�)���^|q]F+���iN9��Ǽ�8�ު��5�L^����og��oT�ԛ=ϥ肄�e)�q�iT�v�	ħg7"�,Q˴��\د��۔�i�[0b�ӭI�2r9��s4y�x9\�:梵����,�]�g����ZS���:�y(����+�5��l%$���N�]>Uu�5�oG�F)��M���Y]��N;��{P��p��[�U�J��J+��D����I�R�����L�}g���[ ~u~���飴�F��ki����E�e��;�i>{+z�D�D�sr�w�����9��sN�4U����������g3Ci��^�����l��0NNI��=�V�V�y���ã.}���ct
��Ѽ�8�H~��ꪭN/g��j~R=��ܚ�g����s}0�F��������gZ:�y7Sv���Vo5���V���\7����(�7,��0���of&��J��㔓��UG���w���S�҆�4u׮�y�t��u�-�Xϣ���EUBQ�P!Z�q+^X}�p�9����~S�(�gqE���3�F��Q�ULK��)�c#�.�*�-������6���+@�-��@7���>����̍��Ҥ=ګ��4>�?	g3њ�J\|ê\���g]�n���Uj�蟗(�(�)�n\)�w-����4�Ի䞻���]^���O�E��bR�۸�T�����p�NC�:��#�®���H55oOC�n�u�o:��r��Q�:��H����2j��vn�6��U���k�S:�w����\��ط�Խ�>��uel���y�_V�w/��7�D����;Ҧ�Q��:&�.�k�n7�WCq���~������*@�B��H(0���N����Ɇ�z!�xّ����Z�������A�S�e�}�Q�n:�Zn`ڂ�Vwz"#��==S��mt�Q�6hz����o�/m.��Lyo�S�sиv�q \l*����+׋��K��{�k�Y�+��Y}J�-��TtsfrqV��,&_�+��������φ»�N��Ġ�#�MA�ք}N@��tn_Ye���֗oˌߪ����z��Pڶ���%ήNV��f)�I��������kn&�������UWu���gC�n㍄�E
��t\V\f)e����΢�`ܡ:^��#�.�P�Ƈ��Q���d�JSЦ'��в�f\D�G�KDb��y��@\������K�u/(�|��Ͽ�s�q^�e�?���p��W�#�T�1+^X]���۪���uS��=��v�G6�����x�P�(�B�a����&���-г4�ӆ(\	�5��s���V�vGS�H�o��j\)��o"b�3��_h�i��Y<��}���&P����c!8�Q�-c��/�|b�4���Z�4���I)!HE��3����%z�w���*���s������b�CZ��4�*=!��ǳ�A��q��7�*R��nݫ��*7@���<���4^u���o���m�� �+Ǔ�&�z�|��6Dd����L�着����sN�χ����Q��t�k�������Sơ�s75`��=UcT%�a_7F�v2�<����/3���ǀ�}�IF��@ڈNq�U뮼NkN֑T�\kSt1���o{�;�y���j�����S�7)]����󳷢��y��,7��S��rl�V֏TV�U>ڢ�m.���}5�{]��7�sU.�'%z���KU9���L����N���;U\|���W}~����~iM�T'�[�T���yN�(߈��=/�厨�²����
��<eS{���O;QˣJ�\�\C���=ڎx����[[�O权ϧ�m_<���\��,���j���a�����OvMfl^ΦٜHR"v�2v�ɣv�D��,���(����gy��\�R��sq��;R��7;�o����4��v��\�V��5�{�t��^��Cƙ��Na�TM7���izN�W����@;ϫ2�.U��_fT�L@�釡�m���Pg\��Z����x۴͇�nS�ͦt�/4(T<����TХ��si��.��V��k&��
�Qa�5�vPGx��(@T`.}g�;�������%R��o�s��pڇ-�e`��W+��	�z}<O*��d*�,_-;Uo<H:��P�hWFK�S���+���ɛ�Lw+�z����Gh�r��M�0�e�jc�R:�D�:�<�V�R(�G0�3�cd�ͦ�T�*��byf\@o2fo2�U4�d*�n�Uޚ�DĹ�7�8�e^
71�i�}h9��?bǷ^��P�utn�BX�,c�#����3�:�|.R���T/ے��R���aw�p�;�;Z�7=����Em�k���i����	�V�]D9}�^�Zؼ{�A"&�t^�eۮ��qN���+��1�͆򦡬O�۪��.;GϮ�Afz�t^�9�k=T�c\��;�ڎzz�L���o���Kl�qxq��/��Q�	vt	��4�C�;������\e��O%B{��t�<;�_n�U/4�s�ԭ	(�Sp2w�k�8�_s��Um�Q��Ǹ��1�C�;�"n.{��[�`5������E���5j湆љ(�{��54�\vmrӖ�����i��F�w��׎�GlJ���BnS[ �����Bq�#o	�������7%�]�ۄ���_T}��+,��|��T:���럮qXǸ��DwKۈ�lT_7�I��C��SXj�A����f�q��W��)`뚃ZՌ[_+�*�kx�!�"�SG��������5�����Ġ�#�5w�i�+���87Y�3t9�z�qOẻs�Z�d7�
n�E����8[_N��J艍ᔱ���qjk7�J;Y/���b�˺�>ע����a,�2��+ɫSOy��I��qg����օ���LEn��K$�neD9F`�L�mS��uTUa">�=Y��t��s0밻.����_)����G&-�E���X� tM-l!r!�LD�CU��YS�V���2���+�:����&4<[�ki��k<���a�G5=\߸xVT���lJ윌Ov·NEO7��\��í����]a(|�C߃����2�l�ʼ�s�H����F�R�P��ؕ�ھ�и�:�_3�N{{�dϐ BxRƫ���A��A~Yy~�����|�Ʊ��nq��&̮�vP��P�։��̫to��K궥�,��z·��9�p#&��_������:rS�k�����ݙ5�a\"}�a`�l��_e|i�:��ћ3���s��z��{j7��na+����ڄ������pM�+WL�Y��y��=<��{��ص���sÊ6��<�\dCC+�.�A6'�o�	��55C6�t���W�>�J}K�����8\��LY��4�����Ǿ�yLP����#�T2�b��{�ix$KѲ���%w^�|���_�zH�l�yE�y˛�_+��\D���Uq`�$��qY�5<���8����rx�>�ޣ]s���[���L�SK
��z����!W����ئw�S��+�ƫT5<�|�g��ҕ���ĥ�0Vw�7y2{{�uK'�)��Kq+�_d���}#Wr����m9��m����˚��7����le��5	B͉5?�U������n*��W��I�kޥƥɋ2bKaK<Dl3~(��װ��K����*^AԹ9eù%[�77Ik��vR>qһ�'�+7� �/XOV��yVX�����u�`����}:m����a���ub�sb��>��"k�ϵ�9*R���ϣoHLvI�b�f��ܺ�ʟ�}�}�G��U�\�R*�w���*��U9aО��O���N�Tu���6�w+�k��H�����p��;����_w�K�~*�%n����}�o-zӜ׭'9�w��O!U�I�ΐ�,��c��*����n���_۽�a\�s.��WW�CWn��T΋�e��ĄV�]N&d��g�-�\&�B�K��֬������TCjZ��ag��p����w�f[���r�e�k�-����^���=�q5��w�L�5���D�,�;�4�_J7v�@�˿��3�}�y���r���f#��nR���w�k�\jW��(;Y�k��SQ��|�|\vW�սUy9�-��5���q12�`;,	$|�{<��8��G�^�S^ު�{�����{���`��y���e����m�3�E����q��^�^�~BmrW��M�t�'��T�>Ktv18�=������հ\�(LF�TNCH�{<��!�'C��c�t:�����S*C���&�`iF�|0�'(�o��w�}��Ŗ��� �o��]�����ӯp�4�P�][0p����ٝ��/LF&B�����񏢲��	��������p�?y��z"�*�Qδ�\����k�i^��<�'.�',tR���\�\:��o+�=yǣ9ۄ�]�M������Y2�T�mNr�6r�Z�Ī���M@�+7ӹ��϶��Wϗ�z�߷��ts5z�(�Y���B�L:��#��u'��R�]�J�سO�.;���㏝i��'�;s���彎6ʿ�%C�eD��ϭ��5��b��ʣ�ݭl!9OZ���W�W;
�z2]Қ��L�Ԉԯ�V\�U7;:Vrg*���Wa�ˈ	��Ga掴�}oҔa��`�jf)�Y�1��R�;&�2�2�y��o2���[φ&k�v�ÁHa1�����WiG&��D��%�}l9��3�,{p���ã����Uκ]�f�ᴽW�Yݾ�FA�Q�G��ы�M����L����d��_�º�N��r��1ʳZ����u���D��C����&�iRm"ɼA�Z�2��*ћ��ӜGT����c3�y��$�=�����rV⎕Ƚ}~e x���ά��ɷ�}΁�9���$ds�������zU�'jR�)Ӻ�����i�A���+4 _.�a4�孳1��!$���iǱ.ά��޺>���	R���/jY�i����;[���(��x�sjr�����x��Zک\v�d�2�a�=%�����k��2͚:���{Ç&9u�W����e�������ϱV1�؍���{�����4m�G;fr�Q��v�H���۽�BAV�2�vr��6�b�Ɲ�^���]�3ep�\`��[�d5��ƕ�&ı���8���ZX�6*�Ѿ�B��+
��Dpx
����K/:n��o6l�:�j�R)GGS`n*��8�^�b侹E�J��b�KS,�8�Y5Ez����;�ɽ嘖�@�����1�56'd�b�N.ԡ�!���PV��c���WC�n�b�Gr�9d!ь�&K֐��aG0Kۅ��q�9�9��I3˰�	��������4tKi�c�b�Xi��V}��+��Rh
zH.%hJ�F����A��!@�u\Vcޚ��r�KB3f��A��]p�oΛ����v���ӻ��m.���Nj����T�CX�T�ƻ| �"��<�\2�_Y����R\ek�C�R.YU��p�h7ܴ%�q��m���\�cn
sv�U0@�rYq��Rޑ�[�v�r%�N�����U�=u3d�Y�B�M��B��C�>V�L����n��WsT�ӔV���:�	�v/?r�&��P�z�65U��{�4�t�u&�N͍�ĺ���a3xh�ӓU���:�	��+��X:o܊�RN�ga*�,p|L�9o�:�W;�Aӽ��R(:2S-ނ
����v�b�NKє��c�gl�܅tנ$��'C�Ȭ)26;�,��.���ش,�2��:��m�2�(n=����i��^���.ޮ2�	گ�'pt�_,�,S�	`A�28}�"�_.�٭M ��A�F�f�j;����cUr݃`7ך�Mv�`M�9�r#�9�l�SK��=�;���`����ܙd��'opo�����RL}l-���Wl�,�,�j�H4�$oea�I�����8������Ӟ�>������a��ڥ>`��@�#p�͸��7SqV<�ŭr{m�'������N�V��AM�h�����{Cb��}����u^5z��ꇱ��i���Z�����z���� +���n��뮸i޻�"���Wi��9��;!f(�%hWU�\�>Ur�a��.y{V�P�'u\����pSg�X2�wgq��Yq8���w]B&͝u��m�����1�s�S��zۛhњs���v�pw6E,�`��	�G�	�����|m��x�LP�*��1T���j� �H���"�9�2�"J�u*j6٭+����ڢ�[eڕ��Ʌh1�aJR�8�W���X�f�.��رC�����Z"�QQm��u��Q�x�s((�RŌH,U�m����m
����*r�"
Q*(�Z��V(T�i�.[g9G�8�P�lX��h�Mj/U�6�`�
��KciKTV-F�5U���͈��EJ�)�廍��EEV&�m*Bڥ�±y��j$Q֤U��b���j����5��X�cmw.�q�+)i\%E(�հU�v�!m��X`m�5�6��d�**���+�C[�U�!������(�QkY�����k�����:�L���li��EX�P̥���UTEkUV)q��*J�Eך�K��&J������1hC6,�EQ��
j�]�%{�v��
�n�]^!�]�>r��i�Ec��쳥�r���rr�u'I�q���>*�'��4�k��U_W�<��u��������;���|V9}�u�E�v��X���	��1oaw�j.qX�>���Q:1�چ������㲠�8{R^�>�]g.1�$�5?T����-�8��/�ޭ�<�F���o�7��-�+z^n�n��9��Kv�:��qT_uTb�tu�V�TԧښΞcaQa�K<+E�Z���ٚ'����DJ��<s�8�c���K�\ض��3�I[��'��c3�҇sվ�����ܗ	��f��u�����/�Ʃ[0�D��t$k;jmE��,�I$��s
kz����Ġ�"�͡�VV�wO7�:���j��ߩ��9��_TO/�p�m7�
o��GL-n��X�je���aCS����h�F�57���*�vG�����|�:��auŚ��fﶙ��;(m,k�y��~FIm
��1wV�E�7�ތ�t�	*e����Nfsh*�Ar+k����tM������.~+�����X�7d��+-]��M��t�.o��h��cN�=H߆5��8��e`̩Ab��V��04�������ok���|-����s�y�nb~�5�0��ep�]ıq��AZ���}��}�L�cGZR�������*"zd'�pe�}Y�R��y�O��=pD:�S7m+O.�f�SBe�Y�j��T�2���}�
�y�Ȧf�f�ζ��jf��7�����R,�t��f�[+�q<͛p���lV�۫/^��!'SO����Țw ���E�T[ykTL�oZjq��˂U��wN����Htڇ��
�ƀ�r�rz`����NH��m�����m^v��wJ��Ӫ����9��xlCVhĩ.���q"8R"С0�+� ����jv?S�ZXk׵:�	��<C�kTc;]-��o~�\V�tꏱo˩{i�,3�se�Y�j�0Y�Rq��`�^����j3F�{��"���9Gi˨��O,镛��
C�|��?�.헙�7��+��%}Ƈ��~�3x�Hi����r��zaj{�U���ԼM�f��6
-6\��u��L�g�#��8���љ���қ�~e�Ni��g�� (��7,;�R��:X�%�V�f���9k���
彜��9Cs��͡�P�;2v�uI�H���U�ȴu�����.2]��ѽћލ�]sw_<M�S{P�b܎{�gѰT�RH۬��\�V���r!��c^ŕ��U��\c�>������S2ogi�a�.�J���P����-D�>J�Wk�ù%������V��R6y8Cfn[�}_aa��Y�Iق�
��b��U�$һ�f]�܆\�u��b��,멨t�ta��X%�M���^�d�ڕhI���Y���k�C���O�{v�-ؚR�_��s�mh]��d�h^����v��h]l%1˹��z�;�ܞB�c)K1�.�0�i@�ōV�
s�i0HHU��YA��5�g-��+��]7��P����p�ұ��gꪨ�8u�Nr�ie�[�qc��qmDwQU�)�z͸Wo�hۦ�j����sS����k�l�ʋ��R�o���ݓ�r�k��>��K���:"��s���n�v�K"����1�/M�h#�@�gmGb�?$��NB��!vT�[�o9�
��i\x�Ϸ��蹸\rn7t��ţ�<�=��
pX^�7�n�wp3]�S���V�72�mZ�\�{�5d!ή�4r�}�}�ER^�M�\
��Ϳ��O�J��O�����;�y���b�υ�֥ 	Bgb���zݬ���)�����no��z]�ꇪ-�.'ϧ�b}�r��6�\m:��!�f&%�T����K��O9��f�y�[^�m߫Ly�M���!\���_w�[��7WR�<�}S�3��.��gE���߫��hrVR�|F)�w�:�ؙ�]�{��K��]cŸ�Q�eB����kr)��<[-r�Q2n����ә��ۉUZf'Z�ʬ�w�P���>M�k�k���*:F�S,lY���m�������k;��):NQ�N⳽��[a	[r�VVi/�Ku[��8��m�|�ۿ��[b�T��ʡ�Y['��������sۜ�Y�G[�[��m+q�)=JS����:�G)����7U��yeJ.�p�f8��]�b��U�)}��oFK�SP���Vk�>�%���9֤��F�hܧr������I�����_��z����;�B�Qь˸�Ǎk} �y!�[�j9�������pd��u[_�9ّ\��?KoC!�(�RQ�y-}f�2�{�9 R�2^
}�U�*;�Vۤ�����ﶛ�3 ������2�WpfB{۩t�k�����Pt&܊ӏ7ނX�"2��n{�z��\p��LW+s,'�
��o��������2-�詬8Ĭ���Lĸy�],��:"�M0��F,{
�z���-ȡb]P]���;����[:��t�)v��K����Y�w�����(����ls��omu����h�tf� PY����瘵	N�p9�]��f�O�M�F�*1����է���n�r;s���2�rz9W:���J����oMDj��Q}�\^�:�{�4����&a���7(ҞYȩ�Qx3k.q��߱F:�?Y�ʞ�x�����WlXT=4yȯ��g���;gy�n�8���r��c�@�A�ݞ��=nIs�9��Ojr�i�	�\���<�19�gP�,�a�\��=�7uΧ�& *С+-�N��Bq���_I\r����!#�'x�F�iޒ����/&�ǁӳG��d�����R�2s��������xG� ��S��$rj���<�d�ob������9/;�F̤�磌�2�-��xj�ԋ�kZ��n��{��H���w��d7C����Ǫ���{�|�s��Z�������oiM��am��P��@����F(��5�3N����Bm�>Jmj��*��1C�|6��_q���wڧ�I��#��)6T-"��˅DZ瘺oQ	�Sq����Da���y��G;+�����0�@�Xx��������H�`��sP2r�d�쭍NntW�z3�/�&)J1_yCU��-��Ƕ�|:I[y�^KS}R�B��x9���q��R�y��T7�b���t��f�T[Wd�Į����
�;zUwV끗1�ZN\>��Mà�&�	g3њ�dQ}��i�o̮� q��x��ד��U�N;m����+�{��Ƭ�t�X����N��i�|N�3Y�y�_^-נ�j�w�8Ɔlw��a���t�^�c}�M
O,E�k�M��+�&�{-�|rsWk����G(��a���{��$��tx/��VU��´\�]Ҥ��%�^�,��Xǳ�Wv:,}�7YI��FG��т�;����X�m�D�n���,)՘�8�8W~����d\��ݺ43�4]GH�8��*��r����ڠ�]7�N��I�S1��yٛ��/3._˅�@fT9*ȹΨ�9_F(Ǫ/�Vd���������]{��ݪ��ע��/ ���+l��j����sOy��&�I&���P�T'��EIצ{�����a��O7#}�=���Ǜ��`�7�5�=sN0�+���������)���M�Zx{��F%���� ���sNb�&r�^���dt���o�����gԜ�)�Տw�# �{W���KP�q�R��m};"R���\d��z�����`܁r�k�˃���y7����0�5�)p��5��kq ��6��d�VB�Vwy����'�sHNu@�S5"8s����U;<���`cG��Us��Qӯ�������V�FB�z�P�YQ�F�맴f�h�T�U�ao��;s�,9�f�Ʀ����C.(��ъ� J���Z�ʃ�z�6�*vs�$��[7K+�iaXYƭ�r��(�Ċ�S:s�!1��"�9U�.�k]X;�Bov�[�%R:|��t]��.{~̈�VPe�}�«��k2ƵP��9�w1֓�w����!f���\s]m{EJy.!�3�'̅[���S��8{M��>�k���s{S,���েq3���^���,sZ�c�.U�����6m�3��2yC���b�y��n�#^}��=��M)v�^K������n���t*�T,�k�$p����Jq�@X)�	_z|���j/1���b�*]Ol��y��UrJ��Y��֣�8�hk�3�7�+�|�Aq�Pq]E�U��ަ�Q�j�氐�y���z+���O/K_O9��f��o��m߫L�	K�jH�u���h��qK�0�<�iJ]�ǖ�Օ���*����=��#�Ǣ�^��6����|�C��r3�ϟ��;~Ҳ�syoS[�OvPjFI.�M�p�^ܸ�W�bUAWÌ��V�VyW�_;�*���4���fʠ�r�����������#c3��3�J�f�p\�����rɒN`�Ր�(�����xm��{�K���N��)u�PK�n�3��}z�PR5�v�<��PXu�{T�k��Q휦{nx�������%�����783=W�6�g�i[q�k<�-��rڅ+�Gf.{t|R���m
�++};�,�^&�R���1l�ʵ;M+S.v��>�MmGM�G���urx7u��a�����5wC�;[.9������\wm�ђ�7|m�xa(�W�9M.qsV�U�Jr_ǭ]���w���B�\�b�.��0����-���$�CFUxf6R\^߱w���'�]3��.̄�1qơ^p�BF����N�쮙��M�L�p�=���&�Jܼ	�_�\��˯�j��!1[�J�E�|��[����,U=)W���Z��������ٱ\����^�8Ne�'�l��4*�(}p����\L5L�٧�f�U�*���k��	N㧽��_=�
�ۯ�NZ��a�
�����ۃ�P�}8�k�q�f/W;���\v3�]A�n�HqQ���ySM`�|�ȗW[�|�܁jФ��,�ݸӄfu��;b�S�{��EIp>�NG&��4nsK�v�t�s�uw�;�����G#m���Ѯ���ca�iF��Hi��r$�ν*=�1�Uۮ�vymr�{B�����t��L���������+'?'}��gO>ߊĽ��oRs��i��^�oso5�~���w��s��>�� Jڠ���7�>��.��q�z�b�[ً*����N��n�`����3j�A���m߉����K�v���p �]B����V��g�o{��4���z{($X��MA�j�����t��zf^���N��c�+Rq�Tjw���)����d�7�!�J����n&�=aM0�\��:�y�;x���r�o'VW+�V�jyq�m��1����cB��:�	{F��fv�ht���yђjKq?R�w��T]ء�<Ԥ��]]c 8�x�P�p�5P�����^��F�L�:�'�K�r���QS

k��Sڃ�[��k��ܾ��왕}�M_DJ�g��i2d���P�;������y��͌U��JQ�jt+z�-vz�m߾��-�H�'&�y�w���BV��L mX3S]��oGk���'d��B�t|�'@�-������yv@p���Y�kPʊ���V�k�z�K���6��2"� ��k�b۳��x��pK���<�}��[@�Td�ܳ�o=�\��jXr��&vm<�y]=e<�[��h�DO4���"%��@O���Nf�7{�5*�C��*�����L5yž��N�N�l����_V�R�@zl!��=�9�²�v��p�m��<���}�n���!�mFM���ı\���KG٫"j��k����L۷�zY��c������ǚJ`�߃%�I�j�鼮�ϲIK8t�%`9��>�%}�mC{7)c�,= kiN��+�>�kZ�(cL&vq��ѳo
�P��c0Եc��f�4�l�4� ��Z��E+����0Cy�q?P
;�oƠ�9�]�e�����AS��9���_��c�FW�/��o�K;B<��ZFet�չN��ͻw&ƙ����-m�q����y��S ���bu)�h�}M�uɛY���Jw�31��v��t�k�����`�8�	��m�lgu�K��Gq�6q�N�/e�r7S�v����c"����q�����//Qz�u��|�z�˼��=�j�ب�겪	��'f�;ǨQ,e�Sw���BgoůZpk�ս�5��LN�Ѷ�-�1����x}+�i�v]d)%*���&f)z7:>����9U���`����ً}�����(.�9�</�Td�-����y7�^i�908lVy�F ��x5�	ԥ�a��/��)�{[�ӻ�Se��d���(fA�j�����{��N�jlYL#�������o�k��o�&��%�wN��q�n�QP̬q�n�;����֡z��'ٶ��Ew��gTTl��nIY�-u��sՉ�^���X1�3�k+/^̝59b�V�[�`�V�l���ޑ���g[����x���v�ðl]�ܸ��@�te�P=o#�[��u��G_]B���o�wR�޺#�=5'�;U\�C�v��tWY�z�O{kOdZ^q5 �^
|��㒅��i�ϐ�Hruq[�%֋]����.�M2��~;^���"v+���x��}YV��{���F���;K��	m�g����䣥�۳��M�vf�YpN�fģ���<۝��[��iP�P����{�V�w�l��Pϰiu��y��Z�pK�a1d/D��`Z	\�R�-��vuqTI�Ԑ��7�̕�zV�;���dy:���t�خ��2v1(QX��F��;s��30���j)��E8��젶�'���<��9S��*�搸��ް�	]0���{7�?5��6�{er�qZ�NrM�ghl����vx�k���#�NHΎ1��Ý�K�l;��:��\mM�+��Y���ݜ��kMl\�{���t�FV[�G�K�ic3)�gr[N:��mֶ�m3�36���mG<M�SF�kyL��JԬ�������8ػ��S5U�Db��;a���Ӕ����PX�E9j����%�������U�������eeB�/�Y�DV�jb"pJ+�UK��������X��.eV�P�++PDbh�3��V"��&�[yh���m�q�)hTjU�"��J36 ��#8�3u%U媂�J�[˒�LZq
��Z�gQ��[E����U��YL�1�<�vqS�����*�˩-�syl͜j��Q�)�32���Ռ�UyJ�����+���0J����+�b
�+�ЩEb�J�؂��6�J1GZ"�̣\��\�"˭V�W)+QCYUAb(d��r6���2���"(�-�[lQ[P)�C�h�%�.�C�e�M
t��o8�w�jo�#��P����Jt���q!��%t�B������*��Dϫ��!��DT�ru�ܯ諭�F����܋�ֹ��R��9�r���I����,���؍/�C��<R��pX�CW}/w�o��{����;C�Sp�;�����2�}�����Q1��Or���U�x�iǎw^oHZ�j�dn��5��bM\���� q������^=�Z����]�D8�Ɔ����F�SPj�Jd��a=D�{��p�v\V�W�˴�U���rޭq*yZ�ީ@e��OV�Ik�\���%{���e�k�Q�6��.�z�Ɨڧ>�q*,+)-觛�1J�����X��CX7o��󊬋��'�|Γo,�B�������i�օ,O�"��7���u|�V�0v�˻�ܚ�t��f��g}W;Ҷ���#Zoe>SZ����E�5�@�y��`˨s�Z��*�\��w�Y�VW;�V�S���v}ޜ�$>q<����δ���)r�ޚ��z����ë�'>�p�A��n�n��-3�8C����2)t�}�Ȭ��L�c�S� �w��1�S"B�}�RPS~�Zlw0S�_I��Ю�z�6>2�#˺j���؄���@�|�Y�W]�ﾈ�Tzw���=��0�������5蔢~��\d��z��uw���_a�M�[F�>Nvj{����{����� 5n$Ԕ�TZk/�\���5{*޴��p�N�\w+z2]�W��U�J�r��OI��ۜ^����HV���h!9N5)�Ы寪�б���<Ǉ��� �a�B�]��R�1�yT�Yp̸	��G% ���O!W��M)f*�g�8��X[wO#1��R�;&)�/rkݰ�;�i��}�u��j�H^��3Vz���oL�u�ƞ����,sQ�&#z������]\å�����u)�f��{0�U~Uݞ���3@�iK���\�%�����p=��U�x�����\:T:�Pz���w�&���_��)�����b��)�C�ƖHF��ơ�Ǿ}B=�_c��Or���Q��:�+tO�T�~�-�]ڶu�g2��q�ն�	i]Y�$���p����k9����LH��i#�u�(���l=®$7D|\��n����H]���+�X��V�4-!����S��;	p�eM߆�(]7W�����mXd�2�qϦ�1 �2n=�r�\��v�����\�tW_�}�|Vk��2uOu�����c���V�Q_w<|29���ީ��E���0���d��/���o7�8�wgvN��1h�T_V}���{��r��xo}�ZݗԻ�����<���q�Y}J�㨷��V�u�9��6[.R���u���+)�{�n��O�RC��5�W�yUQ�?>�ǻ-�g�Ӛ=)I�[���]�E7��^B�+�Ī)Bۚ���%��M�V����ʔ���39�r��n}��n{Jm���an&F��'u=�<�N��\�Nͼm���MM�.��������^�7M�e`����ے�Ӳ��R�(�I�-����b��J_u���ndúR,v����x�6p���\*M��r�ə|�M�H�Nc�U)���t��7�^q�o��n��U1-�	�,�sp�s�bV�XO2¹�e�k-\i��qؕ�j�Ɣ�5or�3�f��vT��W�!��T���Џ]1}u�CQX��6K^���E�or':���sѳ8Sp��C�G&�m�2yѢ��[�Q��mKV�z=Y����2�tX�2�t_������P��e���������<�+<+f_F~����؆R���S����J-	K�%`�Z�ge�M<���>���8UVk�넍�f����w��b���YƩ��6�$��~ķ�<��!�ɨ_s�v?>����!Z��潫��V��X�o�����o��7:�ʚ���<GX���3kg�����I���D ��Ps���^�OMF�=t����hl�2�bM��3��M�[ދ�"r#g�ۿV��\v�)�M�ԝF�ɽ�Y�9YZ{3�5P�ǈ��y��y��:=^A�r���Wg��.س��G*�nn��Ѫ�4������
��l����p�A]�3�@�v�ͬ�*��Z7�3yƩQ��{�l���w�����<��=iz��r��:ŷr���qO]E��U.���8{���[�8��x�ٻښ�gf���2F� �b'_
ۭ<o��� ��LU�	f�Œ�P��+ir~f`�+��a�ʽ���ޯL�(��Yt�=�Fr�|G/���;�6"J��k/��=pM�s�uv�9��ι��׋(է��zU�T'$�]٤"�/���Ib������ڮ��
�N�)z�{q5'�Mw58����]��OF�0�S&\��"�WJ�$ܿ��>�	O��5q&�\2-s�]�S}���p�d}�f^vu2� �4���ɮ�S.WFJ�rʉ�	��]�x�T�WU�E:��hi���sծ�K�
�5?Qv��_%y�ĭy�k��3�@1��qٳ�{[1{�3�z}��vs7n:��JY�!vi��[�V�`�����n뗒�S_Frݰ�c��I��5c���.vO���|F���>�]�}3�CziK���/c~O�,�T�M�|��@Ğ��mHi�U+q��$	��Q�ݶi�^b����j�f�o���/�[��8�1�Fe�/�'L7�'�6MCp�{.-�.;�����Z��m>�p���F(0��:+���~��"�!���ɦ�eD4�D9�q]D\�W�؇�W������x�wB#�rQ9�iǩ�j�%��_N�U$ܫ_k�(��{]r,��%\�� ���F.�!S�9{���}��%řN���=�C�u`&׫Ǉo+܄����VIC�w��<q�)�z����ڌ�<�Ĺ�O)J�7�#��[B����$��d��(ɋ=�Qʞ���S��xv�z{�U�U��Q��v3knl�յ��z�q�X�}��Eꎾx�)�}��rF���ۖ�u+G�)��޿�d(nk5��('���U�g�˴�\�������7���;�u+yL��Y�����h��8*�75�֬r؋+��]S���vX�
c9_nS�[���-d���m?�m�7��m��JQt�,+�^��A�3}9*�h��u��.㭞��#5]����e0�C�!S�B����t���O#ʸOY��6��R�-.v�U�w��ɇt�Yl��	TՕ'�nE�"��IM]�n�h����F>�ժu��{�\=�݉�r����C�S�ī�B�X�W
�΃<�\ِ������M.c��Uo�M�4�cH��UQ��њ����0�i+rq<̀�����}^���i�Ne��C����ݷ�ǣ�8�>B�Z���YZ�s-eѡ��(iWM��P����.x�U��_�}�����׿^{�wd�ep��ݵ'O�<�ʀ�X17g>�7p̥�sl�
�|o:1>���8�*�#6���?$ ��e�]��g���a��Ў�4H���]?s>�M6ܺm٘�<ȚT�WǗh�y��S�<3�k�9�w��u�m�/z��+��7�ݛЊu�Rʑ/s����1W׌�,�ԃd��w���p�ڿ��:����s��T?�,������m}y�u�����=1�=��%:�u��),g�P�z���\�:V�����>?>2��Y�ci�jX<k����\�k��U���1ꌈ�����Ƽڈ{�^ؽ�)�"�ݤ+�5�P+0ʕ�ʐ���q=s8��ڋJ�ˌ�J����i�n6��WF�J�)���k���W�Q}��%\�R�����r������t��+��eY��O�N���o~����$<�UB�C�鸭k"�+��V/�-�,�}�t�k:Ӂܖ�.M�Rs�)��Ϻ�o�ݣ���e�G[m<x�ICr�5-G��qN��j5u�(}��oQ��PX�*��a�6o"a��X�&�Z�g�b͈�W��h�W~y�)���ot:QC��-#���w������\c�4X����}�ka2p��ޘ%�2]�yk�Q�գ.a�-�ˎfȶ�`p��Th`�8h j�zuF�vX����X:�n_jZ��\s�~�|�z�a�3��}Dcc��g��������%��<u�M+��.�۵[�=6�u��vϯS�gp���t�=n�߰{�k�խ��J_u����c.�o�	�s&�7b�ptff=c�5P#VT���Y�]�a9�;uTB�n5�M���r��vNnpSk�������;�|D�̄�u|Wt���O�9�1<
�z{a���7\uCw��ϺB��-�?WaM�܍F�*�	駋�v6�����#ƻי��ݩ�p�.!�`�����\�O	��~׬�n�s�qA��Ec*��9���_�P7���`��骫�R��m.��ɾ�)M+��󰺜�{�����nKS%�ݨOtj�����2�������m.��C�['���F^q��y���:�Q��8o|��k�k�m�=Eh\w�mM�]K���&������e�����1��!�/^�+�39� ����_�� ���暝^�'os�)wEZ9��@T��W���V���}�ί�ª�M��jA��5��]�X��fwQ2��SB�l+̞��O�ﺕX��������ܜS�^Pe0���[dy+���]�B�W����)�c�k^W��؏���V�����觛P�-�g���Ef������~*��+�׳��z���=��\�OO�m�ة����[�<���%q\)�t�z�L���Փ�\��ܨ-y�eO.>��oM��VS��ã�@�g Q�x���p�PJ���J'd�b�+|�j�Hiuz=ǋ'���=w�|�D��Swl5qa*��nM�K���UjwŃf:L�2�ʽ�#F��n�y�N!��Y,�.���K��	W�9e}$���]�k��4bm�(���:�>�P�[��GZcE�IϚ���*�%�;�(p��3K�p@y���Z�͸
��>��]\s��5_	E���	l���t�`5�^��傥h;�/�ov¹��*�IӰ�>���:�ٞ�J���!�V�#��Ql�^�ك�ą=;O`Y]��7�ʲ�}7�t�J!��qǴ���.�훽t���U�X��i�κG�������>1s��+yU�hz�j�A�e�t���Ӛ��'��[�}������ҝ�o+\�tR�P�h7�5�Y���TH�(�Ũr�ǰ
��}��(^�hbe^=�L�����y��ޙŎj7�I[m�6�o���QUѢOt����fD��I����<U�h�=�󱋽��O�ڮs���0/�0��5 p�p֍����������o����f]������~^\�{f���甯Q�ʧd��o�����w�i��~�
J�#�g�*7*��y���ތ���Ms���p�k�?q��QSL�@�Ne�m��W�/}0����K��"���!��]�7�v��s�u^pf�p+��4�T��C���u��M�*�����zV�.o-�kr��f�ˎ�*.�tT����ܸ�RؕE_#sP~�j�*Z�j���Z�N��N̬�V27q1�����RCjg+��m7���*�Ӱb%(���a]XJѕ#�Ց��U�1���C�z��ͷq��W��eB�*����h�yV{�K:�g��ڵ%sM�R��`��Y�&�̱V�g<1\D5��n�Et6!U�Sܚ��C+I\�<3�����%�e���2��ysytގ�X�e�[Y�6�(�����������v��S�pS���E+�P@j�`K z�S������U3]CZI>���ds�>y�-��)@�M��=�e��w��1\����j۳��}��l�-�s��Z�/Tw�ݷm�Թ(��f��]�3J[4�(u��_�Jx�����N,��<��#�n�8����^����Nyg�w��\�y�s;�[�oj�GI[�f�H��٦�*\�g}��°���z�Tg�h��T��b�}cQ!�p�e��`?s��w�]�qԍ�3�@ip�/�>
�����L��x��<z�V��ۏ����\�(&�f�]�W��ގ�^�ߵt׫�9�w.�C ۾$=� �!�@��`8;D�p���ςEm�.ص�9`��ܢ�N��Y�e�ʛ8�Q��bܐu5.�T�㧺9��o9��Z�S����@MZl�?�L�I�5�y�q��\��7�ttdJ��xNE�.�"�w1�=��N��rH��ҵ��f��KfA�C%Yכ�_
=�c��k�-ɾ���y�'�����ٱ��u��7R��gY=	�����z�ʁ�����Z�*��-�yW3Ve�E��TB���toת�wz�lEz�"����H��;����g+^�	�4{U��)ʨ��[u��[�=��������[�9�y���座�#E����u����h�a����/nAҚ�O�:3cԑ�\��t4�w�c�{hP����\E&�Aiӫ�K�˦	�(�
8�rh��5�oy�$�=N�����.�Mյ�ychF�q �$k�g9�=��N��mm��6;���oR�{�]C-�͓��`}���޲��m�S��[��ʍm�����7�V-T;Nb$V�N��8��u�J��)��Es���B��ܷƻ	�dwy��^r�B3)I:�_��ԞX��,�J�)Zd�>�}-]୔����cD��T%_ 6��#�&v�ڝ}ٻ�g��7\���et��vhC�uJ�^�B���Cn���fP��=�V��H͙tfw`��U���P38.Y(��u�>ф8���7Vj<(Z$؊����=�1t�'������0SX/���d��+w��;Z_Jax�6rX#�q	q#�3��y���k�څ�l']~�;��Z��kri�լ=�����G��l)�0E�(�Ѹ��_.$�{�mº} �����u���{|[%E/	_x��鞋��7/�k����=3f<��:��Ͳ���+Bĸn�B��7�u>�B��?l�d�<��}��7���[��h�� |P�+]�S8v|�?_b��e���E���J�=K�W��.�U��,ܾ8����!��B9Ǯ�m1VH����4��.�tF�71{�p(VדwqM�n&V艜}3�i�2ϧS��}�����&����d��8��)w��(��s�5i�{�t>�ʩ[U�̨��AV[.MnUX(��X���,�c�fv�5(��J��b�\�9U�9�*<*�TD�mCl�S[���Q6�i[%`����F��)Y+�-f�֯g%M˕ffE��pX,���X��"�`����Ʒ2�a��X�ZS; *��E�P�d�f��m�+]E�d����kL�k`��:�.L�ȌZ�PΈ�����PYŹ9��"���F�mXJ��UqJ��*�E���c�J봱A�R�ef�*
��*�rJ�V�ZN%�1��/-�J��l��,er�FcX*ֵ�b�)��eDF�[b��«ZjsU��əR1�U�r�Z�P���W`�&lE"�Q-����ldF�c-(.f�3iK[�`Pp�!�:g�ڰ��)B���.�s[��� +�lP��l��	F�ou����zvͫ���1��nut�Q�tv��ka	����_j��4�1ƴ�^úHnW|!/�+�pz����{�nĭu���]L6���n�S�����������֜R��_�=j:K)�r���ʖ%��,'=��WZ��uBnT�sIN���f�<IX�l��<?F��˃&�2�&�݅Y�o��{��*˩S�R�^�[��Y�Yu'�sq��"~�L�A��%^^1O��5�O �Y2�V�}�&�玫�W�^��gt4��~j�Spi����T^b��e�ع2�R��1C�B�=7����_ۊcz�_ڤ<jjs��,P��,����U��<�m~T%�׷����m�Y?����Q�-��:��ZP�mջ̨������K]9�=�=�ڙ�����_�~^����跪x���|ϰ��wz���w�b�|T�=���]�D����B�������T���L�6ba�����>wx�WQ=�����!�bCt�
X�����h����3m��B���B����i�z�J2������}<�{tծ�!���_��X+��[^�D���۶a49s{��Gz��BNYC$��:�F}�l=�
�67�W|��|���Q��ːM̭���3N!6�+�G��s���B��}�Jˉ��;���ev�S���6�ٷ�T��Ds�u��v�pֿr��ϻ.�Y2Kͭ���M�mOW�S���Q�#]������3�]�:��0(��Y����]�6�\Î�����T�5'���~���#}/�Nc�\�a8���T�hk�c����V��`m̑^����2�#i�_E��x_����蔏{�������������+�ʓ��}>%@{qU!
�W�aωh�3j��o�b��R7�m�/O���F�3��:�Y�Nxo���]X=|j�a��6H��22��%���	��K���Óhz�_�����V�g���������g�ȫuNH��>,ԑ,�_�wO]k��f����V(����>����{=�wG���+�W��y���4�@���)�c�=D{f���~����z�uBNё�ݔ�d�Q�{׍�{�G�\���@y@Ty�zJ��s�z*� n)N��� ��hcw{����[�&�5�o`�i�KX�=�;����.$���m
�d��j��j�Q��K:iy�a�h�1�뙬�>�v#6�C��3�} 9u���N�r|I�ũ��H�6+y?�����H��N�Y��T����k\�3[Lz��Ud�q��{##��	Sl�>��� ��� �ۊ7y����z�Q��z�u�V�^m{������� ��~�����%g���s�Ċǩ��]��=��ǽ�G��+��!'�_Ψ��;P��a��j��i~=7�S ,�@L�X�{Ƅ���Q^�X���^���ؔs��ۡ����El��s��^V�+��,��N�hN�}PM�'��k=�+��`U�Y���Q�|��)���|.�#���kAYL[���("��w{�b]J[3>ѫ��:^��B��iM���T_�x��ߧx�Վ�z���Ke}-ւ���s�)�m���3��S��|υ�L�7�-q!F3�ږ��/��m�+�Ͻ��
�|���& ��ӘZ��Ch�}8ϧ*�	�����f�&X^Ȏw��)?g���=�����HK��]�:��;�t�Qsc}	�>��P�j:�t��]d����P�'IQ9��+<j�s7�=�*#Bu���9E��d77��r"�����q-nF�4t�W�זV�?���0���9��giX��_F�t��%0��l'�AR�c�?I[+���eo�\/�	�[�,�jLS�2+nؙ��=�װ��Yohѧ�[�Q9�2���ٴz�sꗼ_�5�Wy'���ep��k���m"�"�{˽|�7�^�F�g-�>�3�.�&^�ku���S��ߨ2�w�tW��w!�g�Z��Cf����2>��YF�B�n�ݯUUVY���x��~���}}���_�G�q(��:]�g�ȫuNHq>f��A�q=]o�&H�<f磧7�ؽd���KӰ��^�=��W�>�^������e[����׽QN-�t�s��7麎ی�LLSU�n5χtl����K�^6}���S�;�틫K۞��Z,NNM�zڬ�@'����URG-G_�U��^���/��r����s�>!V�r��G\����5C8����$����[���7�P�3k�z� ����g��R�x��6��'%�7�Z��Ǽꥑ{(k6�U���M�Q��=TB�N����NLů%���]弻����g��{-d6��
;Ί7��v�=���|Oi�P�6�'i���������9u�54�k��t��=<+N�1N��=��>�O�����sU{��碻��IL^Ϯ7�\Em����?UxeFMi��27�#�y��,U�>��p�{)����9}3`�:�"��P��R˼�?���ʏ%����E��g�&\@�d�q�T�>��4<fo����ez��f
vw�����+K����[�黚w�ޏ-�ƺ$[pк�h����T��wn�+�{����RB��GF���f�(Ǿ��W2���*��j1]1q�:���>	�T�9�W����߼W��Nob��U�@����o��}��������=*p795w��L�L��s�T<��
0UǺ*k�U��s��r>~�2�߯Ã�T�)�,�G�@S���r(�����'//7Ǡ-ڝw�^�}��G���U�O;H�<V�?u4s՞�qJ�� �G���*�dׇ���=�����=@z:P�/#e�}:~��{�
�9���mz�����ʡ�dF�87|:g%��~����ϼ^.W�i�K�����׋;(�q#����ˉ��������ڗW[��]D�;�����A��T�����8KGw#�,y��κ�������.8�����g=��Ϋ�{۹T_���p�SG�d���bi�m�/ǻ���{�F��)�U���z�l�3��#����� �����܁}>��6��!ק$�����)~ޒq���@K5c�>�ب���6o�t�s3c������>7^�NO��fֆ�וo;6'&~����F�Ab�PV�R"J*�<�815q��Y�:U��~}�A͹;>R �g�bڕ��t.�P�|�r l�0Pt�Q�a(�dõ�5����� b�M����W�:�/lSץbM��kB�Do]
�����t[G��E_lK8Ks����;�`��l���DnO�WU߹�L^��G����G�v��[+��?�z�~�Pr*��˙���߫c=�iW�N��{�`�m0'��#�#�w�w��7�{�gLUS���X��iB�V�����㞉څ����\f�i���뎦�d������<U���:����x)�=�h�f�~��X�nאկkƗ�?�}R<79�JS��n��3\$�ގ�;�͚ntw���8g��4��ݢ�dO�F�9XʌWp�&wӃ�*��m�n.������3�N֜��O���Gq���w��!�N��
Ȫ�'��\<o*+�/Ϗ�J��E8pV�<��nc��yzr9�p9״�/ţ�_��۬W�m�+=�3r� ��{k�����]���{"mnB��@��߈�����2��U���-�Ը��:S�Tz��z�1��F-�Bn}q�*��y�G�*���2��ԯ[,%���o�dU~�-����������Z�� ���V³U^����1P�L����n�B+԰��KGٳ/�븱n�I���p,�U��������30�_�T�lc4D��Bc��!}�VtƿOgy��{V[��S�t�c�bw�eL�"�^�	�z���.u�Ѡr��HZ�F���-�bRS��}cR��iU�a`axl��S-��%۲y�nה©]�o��\�w#����~��_!Og�L���{�F��Y~����5�G��y;JhQ}^�G3����\[�d�7���{�˧G�s��������\���|X�0|1�#"�����l�^~[/o�'�u�A>�\�����f˟3�9�W�e�Qn��E���h�c*�`����-l��v�:�����2+\�=��.��yW�&2=�P*m�=A��S�.���_r��~�Q�����7���en����8��=Q��b�\_�΁�顾�ٓ�H�Q��
��P�����~{IH�ُj���0��ͯq��O5Lʽ^ӻ�~�������فʢr���w�=�ES�/^�Y\C^�\�b
�jW�( 6����κ�\�-�{�n�{�z#�֢29��ݻt.#��Z.<��?��R��v��m���=��y�6M��
��*}*X�ʀ�o�W/\4J���|����C�#��yN��X��'g�ޟ
��3u~[�/J7��zb��Nx�ֽ�=/Ǵ׎iq�k���ܣC��[7w
;��݃�+=�ᮨ��W�e*ņv.x���1����Z]��>8*��I��YS�=�C}^��jZ�Y0'̩b�^�1n1���3=f��gvYР;��y�onJu2Ϗ�CH~�&��;��n�3����Y+-t�e[+��O1!Ѵ_f��t�FD��NM���g����]��V�~2��/#�B��^g�|�{Ƕ._�:�,�����apMQ�`��S��׎�G��H�\�W5<���a{#��b�����A�cj2:�q�3$��;O��T�_���<1N\w��*�욋�4�QjW��چ�E�j{�֭n���:��O [�+��{��y�a��+���^��U�YZNk�L�=�ȣ#t�ܖ��󷖕�;�r�35���������)��^��G�!�{�����.��]��6`�;qS"�ok�3B�2g��b�>�;�|�͟3W�P��{�x���7�>ȍ7Z.˒�2�T�w͝���}'Ӯ^G���W1����i܀Xʎ^�=��W錃�霈�N@^�T��=�WYlm�^^�j5QG:B�^*����P�ǲ&�=��ɉ��h޹����ڕ�����Cޞ��=S�|,��ڵxo܃G���\Z�h��=M�>��0�=]&��>����ʄ�UaI���Q��Ʒ���}ʀK�������Ĕr�U������ڇ�>����3氙���߳W���S���x�R�]\o���gle8�n���^w����C�9Dwf�!�0H��
�±��v�TxťL}ֽ��pf��Ϻvof���f���;�p���`0��r���>J)��Hv`�7c����� ���ǚ��ɋŻ�Im<�E^gu����ݙhgԕ����������<Cc�IG=2Bó��_�����fZ��=�+�F��� ��\�K�o�(	Yo#͙���E�n�Uǽ�t�>=:."=BP׼��_2jsj+���y{�{�5�^O�i�Fz{�,�O U��zx��ڪ&�=�<`m�_�6�|or�!�K��T��5��ɝ��@��R=��u�}�������ַ�hzE$4O�#��5bՑ�T��}�ۖb�{��9��VET{M}��ɝg	�MuHc��_���w��Fk��W �b��{ۅ��Lsu�Ǝ�ٴ��}B�ܹ����X�w���ax�O�5�����qjqo:���}�֜ex�ȋ���M���9E���	h�`>��`O���H�|�m=�U����.�=�M�}�v9�G5��\r=���o��Ч(��L�ٿK�U|���U/Gm{�+�^��
�OVQs���}�½���~�x�GNu�;���1�p�{i���W�֏ym��W�z}}�}
n�G�e2��r�s>��U��pv�����E�}�5�5'��nTm�غ�<�p�u(yP�A3}b��;��upgL�p,�Y�{�0r�$`*�2q����x����Z�YFnǎFg�<"�I���U�+��#6��5rL	�޼�FnNSe���Y\'����z��!7��ӧy�n��|�����n#� �w��Q��}�P��{��۪D�>�a�Z;�%�R���iڼ�� �w����w����x7���~���+���)ύ@Ϻ��=� =5~������&� ���e��V�em�F���Gź�>sX W�m�V�� Z��\�3c6�u��7�O�0Ġe�S���n�ݥQ�;��Y���Vٸ�~�
9Uh�|=���.��x$rr|7	�q{�^:f�Nfn��c��{�	҆���>�wp��Q���ĝ=?Uh�<�G~��K/Nu�O
 ~�����߻ٞ�o�����.�tV���O���R�dx?����k��.���	�������W>:c��]�>�����G��ŋ�٭7�����S�� b^��5����n`wF��������+���V��w���h>U�^Ac��_��.ץTܿ��af���nw��w^Kk���^��ޭ	�t��]�6�F�v�}HiS!�.&����yꛞ�êg��Y��`6}�L�m�7~ӑ���b�q�o��w³�E>�)�9��X�ᦣ����z�J��1���-A�u����r��)��+m�8��*��7�I�A���Y�K�����9�����U��f�ql�¸�r7rgo�%V�^���gR���v��a�8��� {#��zt�S�������H>ʉ�ŝ���x)��c�w`����Ȓn�vK����G�>���r��zzf��r�>�2�n;��j�e)@p)ּ�븭Q��cש����5v�<��k2^Ip��.���t_�j��Z[A#�AW=�f�}��h��zL���w�Kq[�	� �Ԍ�8��4�@�v�v�0h�Dݜ�{6�o���~]��!e�
�f��Q��b�ê���m���G�o�h���F��@v�Rf�gR������M`���vZf�����=�B�9������n�[mt��P�z�+�8H��D�u���n��q�c���\3��7go
�)>��n�pʚ��[jh�[K����޵8�������Ԃs�|e�;���c�˧<����j�,����|³z�b����A�j<��ҭ)]i�M�ټtּ��A��p܋� ���������5�K��^�W�@H�����V]m��%hZ�]EV|^�o�"�u��S�����_8Q�9�S�V'�0qIe����5������2Wl뾹�Y+�o���,s�VM�Ӂ�}�[ygJ�qxQ Z�qL�a0�LY� [q�Ýw��#�gx^�|Fs�/c����G�g���]X�v����$d�Z �7w�oc���j������\�D�����H5{�L�n����5���vEjB���1�d��ǵ�
/����6����s�����V��'\}�LFo
�N�����:F��T:$�����.��M�q�:E�ZJgG���C�)��/��O^*��4���D<˙�}� �Qt�m�\�P�^�xl�Xr}��ħݪꍽ���/(������>Ư�F�W��Q4XYH=��{[�mL�.���.��5�Ӻ���,� gA�5�s �����Yo��k=G��-�c0l����đ~�����Llc+I�n	⶚��6ٷ<�FH7�z�E�L S��P�n�8 #{䰵w:�x�,7&��oyw��t�$w˴�����)�d��6�j@A3`�9�[�!�ιQz�Q�,�t�}릘�W�^'a�N�*i�b>9y�&|��;͟�\B�~k����ʹ�ta؍d��6�dW���>���zc _���Q��}��؏��uf��IL��� �KcJl�k++�K
��Cz�Ƹ�!�{I�5|�S���,�il̘YH��4F��E��VN��;����n��͓�4$�R`,los��FDő�?G��]ǑDe�Ǻ�ɘF�n�L����X�S�5�P|K���k�W�'�;v����H &5�e��\�ZQiU�����P�sQZ�D�ʋ"��b֛\ZZ�a1im����.*V�6�U�2�Q�ظ�j���<��5k���]��*��9���V�)��m�.�Ա���ZQ���mJ"�vj��j�\�DE�-9L�W���X�[3UQt[e�-�jf�s-��������*�S]��J�bg52,KaQ���-�����9�ZPmlV�m.s��Z�ڢ"&���ӎSk�W;Tp���"��K��\Z
#cY�	��G[�V�V.h�r]-E\��b�(����VǎVZѭjQmh�,U(�F��*ÍX���-΃��78�v*Vۓ���j�5]e�U�m��%L�f��x',m�E��r�6�[R��3��Yu�U3F��m̬��YX��Py��m��YU8���\^l.TK�fa.�5-]�[�DEi�3�W�Tuu\�j����NYY��\�
j��֕E��-e-j4��S�m�+:�g6.�-��ݮU�-�T��Y�a��h�+�b�%B�H�]J�v���s�-��H����˛L�5:��w���[%�Ծ��s31�}�.�>�G��CN�8R�ˮ^�,�w9^ݹ����7INc�2ӞfCC�{NG�/ţ�_�A��5��{ٴEq��6ۡZY}}6��S6�S"�Z,\d��>@�h�ȍq�\q�}�������GA�.��Lߎ��y�z��[�L�Y-�-��m0�g���?:b�}�=���A�����U��I*dW��d1�J���z �k�zwR+Ҭ�-fmCW=Ō}KT�15�No���kf{�g��H{���t/ޯ���9PH	��E)�O��-�>Bu^b���z5����9����g�~��g�v����q�� T[�H�^����������R�/<���ꪜｎ�b;�yӟ��ܼj=~��Ϗ�Y���y@/z���u�"�Q���WE���51��>�~J�ꋗ�Eo��; 1*5b������&�z�>�4�0.��5��gm�*���{�d�G��oG�2|:Mk�j6��G*�X�#������>���uϮ�_�J�^��2�=�	Xm��Ȟ��_�[���^��<�� O+����HzP��]C^በ�������(�W�]���8u�[;��Q��jp[Xݥv^i��	*�R!H����N�/ҺC���R�7�#KՀ�Y�u�g�뮡��M����L�)Ax�GŚJ*�vp�3{o[�x�lS㒙c��X�ɞ�X3��1J�RZzQ�����s�/�^R�$���QGn"v���t�_f�i�/ǧWdz��/��t�/X����-� n�PNw�_�o����fU������/��ݦ��k5��e���rⲍ^[�s^=���烁�ް+�N�ǫa�㑿��\V�*x���<2}����{݇Ur�;D��ԮvUvj4�e\j����e{<G�?�bγ�Z�}�F�N��2�Ej��d�K��zf���P��3���3�^}�!W�g��g����z}��-����8�<6�ѕＬx·�T�Ĺ�\��<�~���򎧅����ѹoޮ�'<j;3�rW�+6P�}*�a���C�6\�dME���n���J�u�P�Y��	���^z��Zs��C�T��q>��dh�����b�����!���2��N}FFW�ݠUz���>�s�Ǌ�s�~Ԃ���5{¡�?RF��O�q�w���^��'���!�fgTR���Y���#c۝�n�����;�@>Nf���p��#�8�W��t���Yn��}wn�9��]q���sE*�(r�2B�`.3s�s��כj����&��/B@S]�;�#�u��[�1�l'=���B	���}G��.�;B�"�$����{V�3�����m��A9�q�C ����rc��ѴjZ����w�N�<��R�h�\�`gF8P}�W����W���Ox�+t�������S�����~�����!zǭ*!�Z��A�z�d�*:
Gn&�=ו�bi��7����τ��MIc[�_�,+�o�z��������z� ���n�m�U^G�蛨{��aߧd�/O����Ò�n�Q��H��w��=���� �u!���.IG.#�^���7�0�6��Wmv�|�`�?kP��03�M��9#�_GT|E暑�ߪ�zI��BJ9~�!i��c|o.c{�1��4����!��mV��<L�q`J��G�3� l�����n*���{�$�F�Rqқ����r���1^�z�ˈɭ.��b����o��-;�]>�N��~�F��\V�-P�ó&���؁�3Nxǣ��]�%Hë"��0Ζ62g|u�1���L0������f4\`&���ss'{y+|/e��7���n	lߪ^��"�=���t���Z_�{Q��e�jr��f?�C�\ܞ���׾�}���o����Yhh�~�H'�%ʈ�8����&+�p�0�e������,��Y�MŦ�V��h���3�2�܊���[F����}ט�Kr�@��^f��*�����-�C5l&�J�()����81]y�����f"ؽr��{��]k}��ت�P�w+���il}sO��w\��y�~�UW3��v�{�gѯ*�)߸��"�lx_α[��3�����`��Q�!N����zz�Z�en�k�@��S�zd4W{���I�r<WqzW�=~�(��4�\�A��(	���l�9
��3��:�R2�}^�Ph�"6XWӡ��Hǹ���}��Un�@�Xf;���U����$"W�Y+�3g�T_Wp�����E�X�>Tv��R.}�w��.]W���nd�}5��o��T���}^ӄ��� ��=������W�EAŽ��o������~�ٻq��׍��UE�쉐���}[F���{���Z�\q��˨�G�f��Ѩ����t׍�z��d)� +���QUW��3����!��ϻ�E���4;L��)>�:��|}��	��s��7�<�D:���h
�;�K�ɺ�\}ЃG�1��sD�w�o��y:��l�&N�=��wa�CuS�����V�d@{FϥV=�Ϊo�I1�;x���q��GOSq�Z=y:+M�����z���s��@��S*q\mug�?
��N��T�(�˿��x�ث�l���ZU�ֵ�Ǩ��⟰�A+�p�W��±�;<3j���Ή��m�ݳ7n��B�)�ā��T��-�֫�妧:'�5q ���C|�j�����([�FиY4b��y���{�wR�����~��(�:�;M�.B:va�ϴ�xg
�r�㩁6�����S�أs-ԟsQ�%~�=��ƪc���V���]�"}#���xj2���z�β<̬�����r�'�i��[�@z۬��߽�����w���h���ѥNE2��3ú}��<��ǞUN��źx�R��O����Xۈk��9�T�|�/����]�dG)(�{@R���
����轝tŞ�Q���H^w��g���^9�h;���}��W~�#:�q��ܲ��b��X@�� ����L����=�U`LT�"�Z,^L���^v_�������ޗ�`�N��$����&��3�\�u �ET���l�h�Ki�Q���~~vı�c^�`�~�X��*=�5��?~����#�!Nx�<�2�%@{2B+԰������,��ڜܠ�t=N��P���o�}=H����������Q�2<� �إ4+������ʧ5x�2�Iyo����0�]���_�p�k�Yנy�-̹#az�����~��`���ל�{wF��WRM������v�\&�a{u�� ��l�;��<��9�E���j!9Mwb�>�6�Ɏ=�#�fǩ��j�eq�x�Ɂ){2AW���{�<q��w�shh�
V�a巏]��͙�b٥�Ú���}���������Q�y]��us>����ߕ^���U��U�_z/$�Y�m瀞5������i�Q�wǰ��+5�񹋏y��u9�':\,��w5Gj��~�� }�V��s�H�M�{o+t����5�A�ܶ=p��b��\{ݪ7�|r6&�i5w�nV�����,Y��y�~�����k�+[�������`��]nE)���جk�u���z���U	��
B���9钎lD�C�g�����ʯF�;�s��}���妧������爸��0Y�fU��V���\���xvvX͕7�~�%�u9�[�56&�7T47м���s���6��vDZu�=[���#q��7�s���#�����%O�ج�� �ߕ�����ɭ=y3�cY	��>:׫��z�Ǵ��x�G���_W���p��C�[q[y�LӖ[8O#�{Z
ʫ�x��3��>E�鐨l����y��oq^ȡ~��S���#%��e�F�z�r;�e�Y�f��2�*�	��D�L��2��K���onz�U׊�^e㮱Qvl��F���+�ˋ�����+*�[�7�R�fe��T�H�Cꇱtx��jm#�J>A
��J򺷡�d�g��eMýG)���}0�cBvS�Wʣ��'Q��6ѝh)�/+���m�X�#�,�HVc��蔏g���������ޡ���D�\	��
�R�]B��O{ި�����w�-��8�]QЏq���G���P�~�
ϡU^������9FFxfkxgɋ�+�J�6�frX+���̘\}}�ϩ"���r=�tU��ȷ�Qy6Hl���8��89�$��vo�2-�Ndl�X���J�G��(��:]�ȹ�l�S�3c<4׮}V^v�Uz䀔����+"b�������r�!��W�>�^��Lv�6���޳K�f(��P�n���Ӓ¡-50�c+���MVѿ�ϸ�D�T%הX�O�}o�+a����R�H��P=7�=C�pyߍ�r*���D�C���0���t�O�N�|B
�����&��֠����8{�b������΀�fd_��G����n���a���ׄ5�S�!W��7�{�)O����L�mG��o2�3��x��Lr8�U­�6j<��r�TB�<�y�櫅��z��X��{�z�+��ٿ��������q���S�oݻq^�Q¾�~џyl��mO�6�����ٍ�����m�Ș�.om2��]�,�F{����:*���ռͷ��S��T���N�.٬q�ݨoاu���2Q�_d:_|_-u��pu�lW�u���鼾��C����]�#����$�&�'�r�Ν�k���5+%)<�v�ޱpƎ����Q.���@����ZxO�x<3���J���j�p;�g������R�~��7�F��V�vv��z7�|�dC�=��}#
S,]���d�����w�T�nu0���H�{VE=���'(�J{��N��{hw{*Q��%"�S�+��i�WL^L�7�L�'ϲ�b�;��T+�[�PC})�ӱ�׼{nX�C�f!����}�-I��j8	��\6��V����_�ݾ�v��(�Ͼ��:���^+���89�Lr���g�@S�.��_g>�^����>�IV��=��|���A�w���s���t<Z;�>�q�^*��(�5$��'&�9���3�OP�ET���S�X�>͖E�hw��1ޅ<��I�����:��VL��E=���3>��U?#�b��ѣ��6����yo��,ul�T�����B2�?�~�=?�ܿߕH�f����3���\,=��LLS���9��=�{�m��Vz�����}g���9mx�נ<�\����Z�-Od�ME�LM>����s�\ߟq�م���L"�X���;�-O��Uo{S	�7��;D
�s>cJ��CH�L�鳞� �+_2r�Mՙ�;-�+d�*/v���#�ݖ�L�l�-�o.{
��x����t�6m����-�U����
ϣSf�2<��G���/�� ǽ�_����>��c���"�å��pѺ�n��x������KҨ�i�V*?Q���<�:���h
���]݈�]���r&���~���X횤�����lf?��᳒5�R���ǜ������w>�Yۻ���}��ҿ����u>����od�^N��z��3Q����_�<3�u���S�Q�8o� ������?0s�8�ޚ�d1G�]�f��HGN�;ܯqb�͚Ӭ������h��	���M�����\@�{��@g���v}�	���h�=�s��:�a�ܭ�y��:�zD�V׭����*�0'��Cq�X�ߎ�G�|Ǟ�2#�����E�ȟV�*r"���W9[�7��y�r>���^7�3}2Ƶ��i^+i�n�B���È��Pu1e%~ګ���������=k�
�ezc	����X��y߸�x�Ƽ^��X�7s����8D�GIdקy:�����U`MO"*.|�J��^�t�tdk�R�w=ģ�kQU8�U�ʋ)LZ�a�b=J5�g�lQ���C��Ӯ��Wd腂�D
���¸����8�?[��{w��n[֒�/7�w\!�j��iv�obŁ}^��K--wgr"	���j$����SNa��aK��Z����qYWM��������p���v}�)ٳ�@>�"�l��jW��l��}\<<�yL)�b�N���-Q��)w�{�9]ǵH1�_�<8�5_i����=��T�RÄ�}�k����5u�dgh�v��r��c��z�9��ԁy����Q�tǽ�p�L�9�${7��=���j���C���P���}����Ly�]����g���\zp ��DS�rGzO��ᄮ�F��N�,���S�v/�{��E���x^^3�y]��N��9/(q�e���|ۇ��\j'/�֊�l��H�:jX�F:#�r�ȯ�\�`�cmu��ϲ�6=��H��Wc{�LNX�I��C^\�@W�W��dk���u�U���V�E�y`*��c��*�X�]�ꪹ��*F�{��s�'3ý���p���`yd_y+��螨�^V�y��=�����0cض���gݾY� �w�Ô̲0��/z�H��bP�y�<w&q����xn#=��'�_��0(�ȼ��A �ϴ�zo� &-_�Kվ#;��F�ݻt/�{�?{ӷ����+���:�x�J��-�3iਞ��gVv�xJ�#����6��]�p� �7^5;���ƚ=��ṭ� )��#9с_%S�ui�r��u��F�SУo/�(e��.vE���-� �u�7�-�[p��Zb�>��Y�L��<�U�zh�c��
DPJ���wW��i�͒&E�$zx�po���i󡩩p���1���"�CZ�����b�����ER?(�������u�����d��9M0u:۹ܲ����t�]s(LQ�.k��h��M������(�V��d�*��o��u�n��vn��O�<�P�ǁ�`q�Z]�x��Sw��U��snPUoc_,�޽I�9�5ݫw��(/3�)H�(�٪�����F^�b����X\�r{������4�;����M���톫��=�7sB6�iK{�5�7�:usw��M����7 y�
���{��OL����R>w({.޼��K۾|�'<�����z�w5�U��������]���݅�ɦ(ɞa��Whܢ^��Au�evZ���V\�4������p�Ov#����Z��|
7�^[=�lK&��=~�Wr��5�}F<p��(�9�͕��Ђ����-��m��鮻f��n�:�T��k���mL�";� �o%d��F7z�o\����C�{^�+��{��}E ���z6�����xnQU�R�t(���E�f��C�p*=m�
��j� �L!��l]8]�˻�]帰ES4�E���[B^����.��*��Ub�5u�B���\;�E�n���N��7�|����䊫j�u��)$"��˥,$���G5�f�˶u쓸�Ә��sox�����,�J�w��(�}������>i����o�p<���$�q�5�����H��aP������N��z�2&Q���nW����՛�}�o��j ��F��5Vh�C�s\���[�6�[�8���p|����ȭ5��j����N;�2a��(+4�/�T�����F�U�(B�#j��e��D>����u���i� w�j����Հ�wF��Ջ̐�������-� :/����y��=�:��Ee�c�Y�p�8�'
ɝ�l����Cv��E����i�`��B �x�jL�y��������cz��6z��ehf\b�P���w��ى� �v��D׮s}��x��@x�Y{�C�#B�3«����Y�M�&�d��ӱw
��nud�m�:�N����a^2����Ih*M�T���f���Z����sp:��s2N5�+!Ǜ�oY�R6֘:r�j1���h���c�E��g\�w+�]�Nw��7�Cy��}��������Qű�)����W7`Rʭ�sYZ�����j6R�cjL掷<fu7.�Ui��Q�Yu��Z��km���͋-US��U��ťk�T�����n��.Ɍ�"��L+kSR��-�V[��#m���F��(�ATK�բ�],�v�Xةm,kTv��͌Q��"Q��q���Z�a3Qj�Fږ�Ⱥ�#�Q2��S��Ykkcm��+Um�T��+EZZ�[%-5����Ռڅj�X"jS�8^Z��9y�X������UTQ�s�1R���nR���ة1u���Z�Nk����b��
�֢fԹ�DԻl��S#s�蹬mju�0�,ܼ�Ƴ���JV��Qj��io�s����h�7�#8���L/-�m�1�%�MhZ:�����o
�e��2�����b��L�S5be����m��h���0^Z1Tu��ٵQ�6�ˇ"��<��4�ix�5��6���M�4Qv����^[�L䵶���#Q�o-�q8��[eGl��km^5�FYkAB�
 #HW��ʺf�ǅ���z�F��[�����:Z�0�k�����m��ŧ�R��"���z�w� g^�b,�z9z�PM,���nc�����W��sq\�>�������|Uw��q��j��w�%ُIs�^�Ǧ\�^���}-V�����kK���L_��'7�ۆ���=O�qؿN�U����Ǥ�Y���jEXw����w��s�ogIl��/kAY�U�g�Xܙ�o��/>鐨l���w/Ey�MzN�vvT�Rƚ+݅�۲��:��I�{x]�E�碫��ȁ�_�3y2��Hg�YV�Υ��1�w�%�D}z2#TO��������#a�k�z��C,�5i����I��5�q�6��kwܩu��*�x�B��i�F�\O��u������d��,��Cs^�@{ӆ���H�w��������+Ҳ��O�^�mCF�/���νix�y��:/��F�Uz��U��UUS#'�:�n�9�)��碦@�|}����������i<}�|]/`٘�f����ψj� Wܢ|͘<��H��=�"�i��2�z��G���b�.fݯo�gxN����:����g��8^˃��$�P��dM�=���LLSU�o\�w`�1'~�vMt	��b����K����!̔��\x8o-�����j�f�	d�J{�P����V��hRI\��x1�t󟟻 ^�f�� ���7�ۀ�гV����8�����B�7�|��Ѻ���7�m.g���\5�WJ��y�#�(��u�et	�YJ��c&yVRJ��&���V�A��y�ě��p�x�����D�Cی����WIǤj��z'2�����J��WN�b��uG��r�9��^��$����]�l{J��X����`�鸽kRX+Ѿ}K���q3Q�ơ���ƪ��^��<nzQ��Qȩ��\��fT���<C��g�_��C��v�tx{fz"K�=���fw������n�Q���=��KR+k���-�I�W��}�I%i��	Cn'i��ɭ+����#}7Ł��@�U���>�=ei3}��}�az��g��W�*x�}���~B�u��n�<>�,�fy������M]��5��'�� ��*H�~�Ъ=�;�r�\=�M���N�+>��i��]1q�:��#�R���n���s֯����Fԏ��w�9�u�{b�^p�-��
�P�7�s�Q`RQ9����U�[��ئG~F_��esʆG:��)S��c��7%�ޠ)Ɗ'�GW��Nz5��6�����Ƞ%��Er��B�f��#�k���{��Y��.1��y��~�oP��8&������Ǭ닪�[S�_��҂}ꄰ��g,��ڏ��nn@FS��F7:�U����Zӄ*>��_oF&]+��.��,e�5m9�l�{�n75JȚ����.{ޣ<�"�Q�/V"��v�J\H��N�hex��x�fܺ�DUH��]0+�<��6XU�|C�6b�}C�����D8���ʛr�x���]uB��Ib�&%�p`��d��2�V.W�g�>
���Z�>����QZ;��3>\lk�����5�����9�^|ʃ�T��}>ñ�-�f��o.Ӊ�~��g�w��V�T����*���>��&+��WHnt���&=a_%bj��̭�dm�Е[T}Ǒ��%�^��G΀�fl ��[�\�*�Ѫ�p������B����P��FҜ����>�qzk�����fʏ{��9�=a�l)�Ȳ��sw�ڿt�^�u�x�䡷�Z=y;�5�ƙ�{c�fC��T}1�q'Mz�������g�0�QT�=�Mg�?@ݣg���+��?�{"'���;��:+M��;,�~��{
�^�P�.�������wnT�?uX��ʎ���z$�;q�.2�ŋ͚�z����������|�W����h�q���w�G\G�o�{�V��=�O�����᯲���R��:�W�Kڳ�o�RU��9��T�|l'o�ڣ��yV�ǾwՙM!��ڱd\�ʑ����Y���2�5G����#�����qiOz+ }�0�wk�Ҡ�[ԴN���v�P�����H����5��f��	�����l{��\y��5{����ƟJT����w�Zj�J5��hG�/�T?}�:�����6���N}���o��{h��Ԣ�j`�^��ح��T{�X*f�ȾW�&S��ɟ/O3!���q��~/�x�8�r�55�u?��ej��y�-�� >���
<�ȋ�"����U��KGE�`�oSKd鎏-�����Q��K�n��ϑ�,�f��fϝ �"�E��-J�u��ޭ��]+�h�{~�Y����ۿ����z=��ǆ)���d77J���!Q+԰�c�+O�^˞���#~4v��uG�]w.z�9��ԁy�����T=��N4��@Ogټ,ʛ��,����<w)aω�;�&�|������mp+!�g =�n֊��S� �$9��g��o���{Klc������1^�ӹ�/�t����]�Q�uW��}9��%\��I#�ۅ��]uO��l$r|jp�ﺨ���D�xm�g��T\�25��ހXʄ��;n�nc�r@�����5�	P�o"�~�4�U��ю���޽�Jd}�zm�R�5
��G�t�;fVv>n�ն�x�u�)�N���� /�4��5k�\�31�Yu�\
�ġ���x�:G�t��ݩ+�]`]?�y��-�/����p���fP��o^�=��2�x��N�3)+}���=3]>�k���`5o��-�_7u�*�]O���n���V�x|:OF��f�i�5n�*^N=l�OH�^Y��P�#��}�5���H#c�	X}'��VM�ЭlW����1_�gƿz���YN�[���ge <�ձ�UO���R'��#���Q�$��L�sgj~�ڿO�6n����q���i�<�M����Z�xDJ�o��~���eh�~�Z/�h��3��
��blS���;|�|�痢����w)\�i`o����Y����:��~��o�=W�Sɾ;���6{KS4|���;�Y8
�������29��#�ׯ�ߺ����,ꏍyMx�����g3Gz9QF�=��l������b�X���o&|�Ȏ���mL0�띚>�����qC���l_��۬W�{�g�}n\�.r�������ҙ�w��y�n�˯(ױ��߻�h�s�ף�<�(�~���G���q��.x�j.{�X�^B��f�Ӓ�oc��ҙU�چ�}~ڇp��k��=�{���z�:�^����;�Y1���ڴ�6r�� �VL��:�4��_:m���5Aw�_˴i������Z��� i�X�^�P��w]�{S�mu��}�n[s����ٯh�����t��W�wϮM%&���Jvڟ�������WV֍�Ӫ-�(1�Ž�c&�ʊ��s���Q��ަ������4j���W�l�zgQL����{=�=�W�D��W{fzF�)�����@���6`����?>����3e����P��{�N�(��Q�F�'=5[UW�\�{+��y�Y�$��"6*�3�tdJӸ\�hzE�N-u�g�͘��y����^�Ngc�8�;^�\���-����ו�bi��7�����u�u�Ok�\�(��Y�=������5�>t<�ɰ=��J����ٺ����a����(�i�z��pg�Gm�p�B|+�Q��PY�Uv7�O���Rx��W�ᫎ+s�pV��$o�L�����7�7�q�K����F�?�����j�|E���<n��y���5}��n��7��y<Y�D:����3�vrr{�,{�a���������7�K7��x��!ޙ���㕾�{�p���I\s��Cn'i��ɭ*���:��Oq`mby�c�y����o�%_.��	�Ξ��ȵ����S�y���udU1��ZX��g|n5��?�2T�S�#�[Y�Oٓ|��Y�:�v��� �-�@�\	�2�e�[I���K����	ZF̎{-(����n����v��]��X�э>��<]�i��r��S��Y���7�����#P7N,G|��VY�ǱP_N]�" ��N]mv��X� �	��������Xe�~�O��!��۔b��Ϥ��"�=�K�qC8�� a��s���>�<O^��_�z��=μ�m��:�e�����ES7.p70���þ�v�X�>���^�<���2���yP�:���J�j���	�-OQg�z7�"�2$�q�uZg�_xރ�`{�E��p*����!����p������}��\8�F|�u
���!�>�^�Uq�@l�ޕ@>Ȫ���W,yf�
��Co�ُdq��>um����|X��e�G�N��Y~�y�^��F�Kd@A��HU+�aϋ���ς�T6D����\�T����*�`~���>�Eϰ�=�{�+�Nnx����0P{2�����>Ɇ��=���"�>�y������,:�=���u[9�x��z���V���Z�Mș�'l�;<��{��ڽ[�P�z=�N����vTB���u~9΀=p� |��[�\��_����e�����m���W�W�3����h�V�d��^�Q�/O*y�͟y��U`�yѼ��>wR/B묛����U�����
m��1Ou>%�u�`ds�#z@)ξ�Y�R�9��+jC��\|����rF:r=[t��gj�9ՙy��M�:�$��j3��>��L��+�۹u��׀=�d���t�㓓��mhw��3��3;X�}�3!�sws�4�k^�#"�^L����O�G��ު�W�5F�G�Ie���?�{>��ï't��2tV��s���>�&P~f��w�7b�Z��q��޸�L��vՊ�{l��{M�>����Cˌ�qb�͚ҹ����}��1JE���/�J��`-�D�|o���_�~޾��=��}#
YP���|U�f��-L�rz�G=�>�gYuH���v}i�{��ޮ
�<����4���,��=�������}!2�uQ�ɝ��@L�t�mO��w�/�ݱu���߀{[LL�m�o���懐�����3���x���	Nc�&|�9�9��:������K�^nY��Wә�<�Y��u��ܲ��@S7��@>Ȫ�(�#"�ȱ���U��Dm&���E����^\P�~�m����įTz�NYf��t���H��l�Q�x��B6ͫ5��O�GZB�*C��{����D�{�$g{��Q�U�P�L����j�!�Dz9�ג�^%C�F���W6�f�b�pnQ�?�'�P���t���z��S�7�������a��ty)����\�OJ����(�*�7����=�gH����s�)k��TU�{��y�r�u%�4S�<՜�і{�:��3ա��SWkyG
�i�W��j���,\:�$}�q�,��=^�>3
�Rw�&eDuV�Ī'<`<��WM
)��{&�o���x����?^���/@�ߜ��g%���m�f�rG����W�Q���{�^���q�)�-�I}��vv�Wz�%y�^���V�\�
@h���1���=W+L�g|w�1*5�^�{���z�G�� �H�3�=1۲=��S�=����G.��񩇗9����+��:���Ŋ��
��3��X�G�Y,^�c�� ��y��wD���7�]1����0�켾θ��'��=N�u{^�>��(�@����UO��K'z=�"��!q�$���=TQ��A�/E�S{�nס���j�^mV��>�龦 ��n��^��޻bx��ܩ�!Z�!�S��x,C���%Rɳ��+u�{Zvx�P�����X��'Q�vR���5�@���>X<6��^�m�7	��r'�Z
�b���3����!9�����^�;ݚ�̚�f�ѓ�n����ۏ|_�Ye�=H��.xbV}Z�i:��l�vRgӤ9˴m�̫���E!v鉍���7�,�"V�w�}���$���}�r0����J�����}ռ��:�l+
�vM�4\���Co�
\l�Acޱ�,"��J�C�?��G���x�w�#�=���=�%����3@Q�,�e�L���D�	ʓN�,y��Z�O�iq�ϛ�3��|o�U��q�l����ES7�s�U`MO"�<��q�����䏡̠��O��}���=����n�c��w��W��r�|Ȗ�G+C ?;5Β���~�л(
�Je�F�4j��p�9l���������^nJ>�@\���y�W4n���bԲPg�FFTJv����/���W�P�z�9�S9�� 'E��H��v}���H�I�@�!� s9�Tȟ��q��Ӛ_���m��Q7XFz�z��{hi��~���%��g���+#��N���(�xق�۪D�=�O�i�Y�[~���i��s��ٽ��ު����W�W�r����3� /�	h�M�=��1�SU�C��������	��ܽ�*��U��|p��R|��������^��=� =�EUy�ux������_U���ڊ�1���95^�W�W���b����Q�y�L̋�����<o>�)������՜�~���d%����B��{u�l��L�a�8ox����KQ˰zq���@��]����z��~&��v������Cؑ{}B���ͼ1��[�"+�2�Z�;Z]w�t�ٍ*G`��cI]�(�f��X܂&�]v�G\�.�oGٮuX:�ܙF�j�z�������5���`��u�%�iL���z+��J�s���`�K��`�{��oF�f����D���.}4^*�u�hw'B�μ�f,���}�yx��+H�M���#���}����vEO;��n��՘��$<�8&����]����]�%^)m��*��ځ��
j���"����%B�3���z�`˾hY�rf��؟���p�n�0��A��4��n^���]Cp̹Wd�E��5�
p�@:g�{5�|��l�/�����;�ė��_� ����ݡ����%a�q�gP�KH�{�Mӥ1�h1yϴMm�c��[Qe��]�sns�]�b��fʏ�*���I.�Q���'W�����y]����9�
�����ƸӣRS�x��˭�S��oj����Y�#���J�l]��S+�bcL���d����A�V2���s�H�)���V���M�wwM��Ww�٤�;G���aMGa��s ���PL�l��欼M��60㚭�6,���Q�֠����O��"�t&��u�nr��]�o{d�ò;�����웄��=�8�5��P���:��h#;��t%����r�m#.���fnZ9u.�i�������\a�*���u����]�� ��J}Vq`a�g���tǁ�]���״13g��j���s���Xyv1�n*�<��SE�vnqF�t��ؽh�S)nhĐ��a���5#r=�.���{�.���o�ȸ�(=H&^b�'u�P٩��2A�ޑ��WfTH�@�<[sƇ�'n𭾚�N��ǐg9����#/�Ɍ����Y=P5�����;� [�e�����"%Z�x��Z�	�<a/����f��h�Gx+��Н!���/��8�u��C#ҍ6R������ � �Edo�!`̶q�����&��HQK�m�oZ�J�>+ ǂ�:sY��qK�I
�힭������06�=��,RO6%�f盁�\(�9�3�K�Bu��×A��ɹ�T��9����U)Z�17!�m���+.��:eq�4�F�ճ��X�
PpV�88m�}�cW�)6
d���G�
�]�����Gr�D}����Y| �Wbɀlt�G�NT����n��ϊͮ� �3(P�WʥBbΘ�P���N�H�{w������v@\��7}ں���т����`�]�N�E�E�8���b6K���Ѻ͔w7�5Ht�n�I�̮n�k����X=A-�Qݹ�:��v�,�>�N�jZ@���B��<�f��(�p�ۆ+�� ��N>[�糔#8���g�o�o�*u
wP�2�9��MM{5�s�T�MP��T��*Sk�*����m�&�nҺ�\6棥�j�jZZ���Q5)�]�X5��T5�ʶ�J�mjU�y�5�YFU*کm֌�9M�P�c�ĭ�jqR����<o���rZ�M
2��aA�d-V�[��ūnfm��y��NQm�X��L����j���-X�f���2��h"sҲ�^&�J�Z3Z�x,9W���ʫF�����k^KN]3Ɗ�r�DX�h��[EԺ�V�3��:ە��UE�̩�)Ym�)���q�EkR�LˊS��5^n+J�Z��Kj��Q]�ɩZ�)mhV�"���m֎h��<�]y���((�J��l�R�l��&r,TsMV���X�resmέL�5V�Զ�̮��q��]n�W&���iFjU٥p��Ѽ�,��ƥ�խ-e)����agiT\\��Ex����QR�h�ǘ�S��Q�V�Ѵy���e����Kh���'9^UE-^M��SZ��d�w1t�QT�ԫZR�*Ԭ�¢k1�lU�7*���i������e�KkD����Dk�KTڡ�B�pno�N��&6x��p�<�~ɑq���K���?uS�y2T�!_c/G0]�Y�VvSܑ{��y��@�����׭��������u����ݨW�O��q3Q�ƞ=���n�|E����~��]\�U%�T1�Ȋ��Q�Y#�=���rg�Nφ_ޜ�r�oK�u�?����g7y^p���:�����9\ߍ�y���t��zpzA�"v��3�vO�i��\���`gB�)yz����<�k�Wށ�j�j��:��:���%ǂ{M��F�X���c�Vc�C�<�lҰ����Jo�x	^�T��b� ������Ѿ�W}�F.��Dz�t��Uҳt��%��w�g�k{�VO�{fW��L��GT�9�W��s�3��P��m�@��u�R�ڰ��� ��;
�2Ͼ��b��+��)�ɖ�}��u�9����߯Å�:�l}7Yn�g�_VOWV[F�=�j���̊���W>N^l�h�r��I�\��"��!�G�N߽�S��n�e�i��5�TyU#*]0*.X�>͖E�hp���N�W��.칽�^�^va�t�/I���[�y=��,dF�Kf���U!T��XC+���z����7�<�
�mp���s�fl/X�]ǝ��޷�� �*��8ig�-�y�̌�o�����L��-�Y����+�k:�&�	�� T�E��l55k��V]�Ip]Kg+���ٯnxg'��ˡp�50jg�wȹ��"���0�*(�yܿ1߫5���^,o�Qs~�#����0*3P���3f�H�>)�����7�s(ʫY��:�٧���܁>��=4���V?^�����Qn�nª-Og�R��o���}�"��ĕ�
��h���h�F�x�A�gR���_�A�;�`̀G��9W[�E�:�=cw�"R�:�W��=���wa�q�Dz�ղj#K��7���X�|�F�{΀�-#�[�}��MUNg!�鷁�䁽R�����''�sg�ͯ	�ƙ���Ǫ9fd3�5��nT'w�Ƶo9��TǼ�(����{`d훏~��ӓ�x�D�~q��}d�7��3�ם�Fn1÷˽�L���y�����C!N��\o�Ǧ�ݵb��l��{I��ɇ}��,nǪ%�,�}�}��4=�}����@M���W�]����
��Z/�=�r}#�ço¬����El�ÿF��ʲ���u�u1��0�59��N��/���H%�\�>Φ���*���Ff�_'*|Y�K�T�QC1UC�ɝ��a���l5����K�}^��3���}����swcL��x=�h8�z\�F�f0�>�2�0���R����XH��F�B�ʼZ���ϳ��hځ�n�rT)�>�ez�Җ��[��ee9�gf��G2�&�����qxG�|d�`r�oQ�a��Y{U�����Ƞ,�8*鷊��[��!�����R���;��``��/�p�&S���g�ӟs�7�{J�>��p�^xȸ�v��KÎ��WD�Q��ܲ�=�3r� �"�����E�"�}�(yu�c�n4o��k�]��λ��l�:5G������m�z���Qf;#\S�p|��$V}2���C�9R�J��zk9s�}�v�X~��|<=�,g�N�������ᇙ���a�l�ĸW-Q�3~ϙ�՜.��c/+�(zVSß��0Һ�,\|�ԑ�{���F�[��x�<����fS��2sz��,��}�N|H�n�4(���@h�t	��\��nUz��[>� <����j��q�VZ�.��J�#�
G�����TDӞӸ��9�5�/�\{����W?N�#�˫��9�W���@+^���פ��U��R�lg��T\�2*5�xv�>���q��}5{�S��+��V�Ld?z�Sl���X�}%ѻ��(��������j={��޼�e��9[�/{���C�Ud��G�:���dg�� � 
��z����m���:��+d�����;Frhy����`�\PG��-�2��&h-�9z* hix���Mo���������|���&I�.�4.(����$�yd^�;Q�\^��8
��/i���c���1]���b�/9��]P�	����"hȶG1n�h�cI�\����ހ�N�cz�dBW��ƪ��o�9<���>�D{���z7����B鎜Vrul,|�z"v���醣6�M���M�0ڷ`_/V���S�ǻv�Nyå^�۹�c/<�����'N��Ti:X��ۅd�\�`g���\�	���<]2/}5�eǺ�6��q֖�q�}OVE����9$��s�Z
Ȫc+&���&w��'7�G����{' G�;pTmN`��k;�s�{O��;���w��F�Β�ȉ{Z
Ȫ�&�X�u�v�t/�E�Z�=��8>�y7ú�����8���m�+��z��r���Ѿ>S��b�Z!`v����H3;������8K	������ף}�uC�xuì��8�g�C�34�&hJ��T�	��w��s��1P=^�l�]-�h��j�N�9���k�z�LMF狀-�����D�v�W�����9�s,t�Q���@�d�}�Pѫ�v�֑��G������n�9�t�T�R�F�p�W���CeA��ۊ�\���0��l��~��J��T<��S6�L���j�#{*����������h�J#Y{�&<�VW���C(�;�Y��s<iWr���Zn7�}�w�49[ޝ�H_[�:g��l�F�4�-܋��^���Q������_to3ǘ$���&���7���P�ܭ�g����u�~�����n����|��(=��L�9��aɱȕ�p�҉Q����Gй�����A�W�3���ǽ�+�u�@��BZ;�7P��+�����,v��~��J�>��C���5%�ߪ�r�)ȇS�z���
���m�U�{'���W�R���'�
�0p��k���U�R�c��Z}��q�ᢢ9nc>N����=��g���4���=��m^���A�w�.�waa�ɏwٵ�7��3Q�ƛ̿������| �wb�&��|�{T߰?iڛ<�(�|�Zn'e��NQyU�����&�{cԡA�\bl���_o�H/b bRt�VTo��p�y�'��z���;LfҬ�N�F�Y��7���#���Oyv��>�j�j�zx�����qW��x'��D�FS,^�֖	'ݓQYz=����#���H뎩o:� ��g+�>�t���{mg*(�<B�>��J��0�w]�j��f{�\m�/]x\dγ����:�1��5���s�#��^:�CC�C�q�J��G�ئ�9�������r��h�����9~�%?]���$��ܺU%H���4!ى+�䙑��-?��B
Vg�wj���Ld\���b;�g�=��&:�v�7ַ��Y��8M�v�Xi�]B���d�{�r窲��R�_i�w�L^��z����\��-��}>���~�1@O*�,2���e����D��w�9+��n{C}��.�6\��59�J�7ж�="��3ވr��nz"��1M�
�Re��_w���@�I�,~dϊ��L��ь߆��Ｅ�u���S�Yydϋ��T�.XrǑ�l��#���꣞=}��zBy��1�:�3�#ǯ��h�r|.2b[6`���*��ⰼ��q��}��Y��]�l!��zP^���Wx���u"�>�I�ۙ+���dx����G�����'Q��=>Ǆ5%�o���o�_��|�S�|.!�U���_�q�����{�M��Q����DL��K�NK�)�zd����Vѽ/ǻ L<)xχ��^>���L̀i����V�ȹ�ʽ�*�����{v��H-�8<6�h�~���iz}F�Η��	�Q��l�(\��|<���uz�a�7w|�P�����?øڵ�d�x=*�g�b��ic�s���V v�FLdNb�,����TT��qG���V�C�4v=�K/ND���;k_�d�x?J�����6���I�B����~�eߦ�|��k������ax�H�S�AԞ��b��he�/���fB���ɮ��z��8��4z����Z.�p��CH�q-��v�G���}�r��gh���ʢ�����_Y�,b����pw3H��PVP0�ZK{��6�	��Űƹ�\��"�ݓB��{l���dR�I�v���y��~�t�;��/���Q��l֝D]�ux	�V�	{+�o���v߅�h�碻���S�=tbӏL��J���~�����ڏ^*�;�>��G��g;���U��^N��;���#��~Ώ!�/�s4|���ǳ�U�J��>�����o�>����cn��N{���W���Q�J����O+Ѷ}��ÖL���B��U���*��T=�&S���^+��qIL����:35w���m��Eq���W��i\���@S7� �*�	��EEϑbuZ����Z�#1;�e\���3��հ�4ltc�Wq���7�WB��\k�vl�P��E�wis9�g�w�ros�f���_����_�G�����+��d��pǾ�9�p��2�q�Q�t*��7ᓵ;+����U#�����Z>͘iB�H���M����=�F��<v�r�7
�y�?1�P��������Jl�ٺSB���9�&�.�n���}���r�vd-���zH��N�5i=�Ec2����Yx������������wvW�IHZد���Gn���JiKyۀ�����q���d����S櫟7�%*��m˼*��뇜�2�p�f�N��;mr��&��2�}��a8���]P�'��U�8�W�^{�E_��$Z�,��ʆ��������sA/j��z����`k��Fr͔�/.#Ni�>j@U�X�}$k�!��t��g��W�+L��s�<�t���Ѷ�`�5QK�7����Ѿ�Q�Ʀ=�#�>u9�P�|J�R}�TM�=������ގ���K5�pI��>��@�}^��Y>���F}�t9NC���j�#���z����{6�~��M˙7z�bp�ޯi��ͧ��;���Dm0��W���j�|E禎��P�^x)T�N�ګ��܅�#�!����t�³�b�q�U����znS V+v�Nx��z�
9���W�\�9�U�Tg��{����!d�;q>�1��c.#+n���f�K}7}j#9���o���pF�%��^��7�Wq�۞7�{Dw��ւ�X�����&w��';�s��\�U{��Y�F��\�����f�����j�(�<�R[;�қ�E���T��:��I��������h�8�L�/>鐨l����u�{b�^F�b����ό,�ES7�s�����?�
4k)���:��������-���y7�;zn��X��Oڶ�fKY��߹�XJyW�C���1��7�7�*�L0����J����V۷vJ�@;"ܕx;��QSJ�|	�h���@S�����w�v���YyE��ĤŲwd;�I��j�$���*��_*�=�q�,/g�O�~��B����xuʤ�:��=����vQ4�(�O!E���x��j.�tE�^.�j5~ڇp���>��dh٘l{�݉�(]����S�^�Uzd7>%힣#*%�@�d�}�PѾ�νi���f���+����k�:�h�>���fgn�@g�}��ә/�t:�o#m����U� =]�7�W_���h��x�q�N�y�*-�9 _�y���0P{t���s�:3+sR�:�L�oy)���\�=H�@,eF�xǉS�|�zg#�8����5���s$PZ=M�>��olyz�o�q�T,C1ҹK�L{ٴ��ڥ������~����|�yN:��=� y׍ w�yzns�.�ϔ���Bܝ��;%iz}]>7�V)��yݟ2����U����j�޾x⪮�&�'�&	�gg�h6f�C��������~-�׆��T����#,	1SU!��»�O���Z;!���~BJ9q����2�Ӂ�\�t�i~=&����6{ˀ���x�pt���q�{}�x��3����yv�ML���%���t�M.g5�m��{���^��3�
A�q��޺��Ղ�3���X+��pAU�V0�B���Y�q��q��{���Wm}_�}r��ɇ�ު�o&>rc��a�m��R��7����=��;w(�*&��yY�q�$��~�(m��1��UhX|'zc.j��-�u�}x2m�y���X_F%�*�<��:�\��*���s�.<�Wq��:�*��N%D�욫�����{�'<lyL���5��쾦 K{���\;ެ�7��Z�\=�M�ˌ�1�b�78b|�=uzfU�-�J%�*��s�(lFL��ς|�C�z��#\��r�Lu��-Я����<�'�/��3G�cr%ϝN�>��~��\<
e���s	��^ӑ����.W�f�=���|��u�n�%E'��=Y���9Gǳޠ)�L�"�Ȧ��'-F�����q�4�<�wݜn\��&���oN��+Mz�߆GNQG�d���t���F,��#���>�e��n-��ҕ�u!�ъ������ޅI��t�5�w���%��f%�p`�{qU!�������M��5	�;���g26|}}\�'v�X��}8vtjuPF�z����}����H��s�1t�hMz*�����-9�w`����,Z��oⲘ=�~u�z��DBO��@		�)  @?��B�����!I?�!	'� B������B����� �$�ЁBI���$�@!I,���B�R!	'�@�!$��BO�@�!$��$��BI�BI��(+$�k9$<� 
 K�
B �������3�g�(�JI!)4ʪ�!�JI���(�J���%�j�Զ*Yl�R��S� V�Y��p Q�����
%Q�v�UJ������[R�H�)�b� (�@h ��pv���Ι�ڦժђZep�t�%�m���(8m̒�fL�6�2j
���V�#V��kXՈGG�Z�e�����.��Uk[e�m�fC�    "��R�@�� �&�0"�ф��J!��L�2dт2a`20110�L�L���R�Q� 4     `20110�L�L�@R#E<�b���jz�Q�3	���y��[�_��5��@ B?{F�#���@	$�� BI�i "���#������a���u�i�XI$�!��� @�xhT���6"���}��0Z�����}6 �-�(������qƏ���CXQBn��|_�ޟ�����6��dܲ���,�!E�{�ڲ���9����"2�� ]CT�0jXMn�حV̸V�w3K�T�<B\w!G>��v�l�D%;�a ��Nj����LMca��E��u%��"�f��n@-��*Ͱ���'v��Kb�EV�x�)�iCs2��E�ږ��Y�J�Ԃ���l�í%����6%���:z-={��[��[�����ړ�*H/�@��zk4��JY���[v.2�8�i-A�S�bԴBɲ�Ju���	�5�u.��a��mGY��m�c�"�Y�e��P�A��n�ܳh:�`��t�d /TV��۴�ԣO\9��i��c`1�⭌[a:Z����z�:;3Y�U�e�;���T��х*x/X�CiTWx�����v�sՐ�r�iq]15dVd�U�R�m�qKna�X���ج��9��mf�a�E����+4������@�V�Xڌ��r��c+6 *�b�o7a�-Ƴ��um�� ���5Zb0>'2�í�p*�ǿH�C�[fL{e嗂��y�/��Lr�F;�E���ެ�kgҊ��FLZ��$�~zre[�˕��Yk�� N^���<j�LN1�e��4H��Wz�ܹ*���jQ�ѵ���_�
앚nJ2d�.`V�	c(	�j�n��mQ�N�p&(���z$�T!Y���[�2P6��%��¯Y�Wl�wr9!6�*���P�q+
�v�����c4�z���[xI�ո�v^t+Ze�8�m�M�j�*.�0�I@'K�pU܅Q��F��T)�Z��֚V��5��E��*,J����>����tiVmB���b'�[j�� ��W����c�[�{)D����Vh�@��H���΢�Q{/r�R[5�ðD�=x�%S5���̖2����C,<a|*��#�$$΍i��c6���j��u��P+s"cH�X0I�X���Wl�8�nb��ҷ0GUk]!X/u����K����ۡJVʖ��'H�6��H�`
ܦ�Z��15J#���^֫H̴�2#��^M�4���t��Z2��VXZ�G �nQ���I�j�͔�������f䩃q\Yyk��ba�\�������L�+U��3�C�-���A�4^R��� ��*"�:����B�S-��^�m�����꿞{���}�#!���؝�z��(g��5L��W�_�I�<��0>�=���h�(�/��c��n����/��Vk�ٙ�љ��o�1k\&r�.�q�Y�WSY�)c�[��E���esDv�7B�NsΤ���L��d������˰�3�|vݱ�ާ
��������1��=|�%بȜ�t�,+ۄR>%	Oc0�E�����@lz��c�7��3��INsμ-3��/y��8gQ��P)��]�)��֊M��W��`',��������.Vz�����7���z{K�6���������3gHo�]Lg��=(>݊�r����|�9k��Ev[�m��ū�W�e�EE,���=�.�t<Z}�1��ٺͦ�R�eΤ��n�n'g��44��(��8�/<�ޮ�V��J�4�
�] *�g��Wٌ���e^�T��r�t��j�劢_p���6���Ve]Jy�s��oy���n�j^�e�2VB �n!�))C��w�bv����[]��Z�1��]0�]v"{�h>�Sq��ɲ��W��a2��X��-�]��}+ے%�ta�/ L�ҒܿnkY]�W�!Vh-��:.�*Ec<gV�P�j�Ե�j��,��j�>�uAs;8Κ�S�:��}�T�c������L���b��= �AW���*��Ah�1Cū=�@��܎�|ü!UQ�������.=�h�6[�ef*}��ݾ�Ļ�f�\��>��b�[_v�-��ҵ�vB�]$u��q.��"�i���5�����6���K��<��17�`���ٮ4��rZi=�/�z�#�a��
rpK���F������FJ���Q��p�j7V��ܦ��o!�p�z�rڸ �ŝ	�ͼ�B+�iM�L}�h�:ջ����/�����A>��u�,�vuPbu�J���Y%ݙ����ڐvY�	��Mws\cGۀa�Ot��r1���[[j}˝�x�9�AmmG��~��]�4���}��u̴e�#8ڣo:��sgv�b#Vi�x̡��� ��+�z'.n冭me��Ҍ�LvY�.�d�a����H��o�w: ���!�N��8ح�����"�P�ݼ�U���1p�7{��ó�4-G�:��v4ΙN�&(e_a�OgmC7z�ZSy��+�=r�R�,#_�\���RBEΏjg{�>=o<�ϟ����-��v����1���W��Z!�k���>Ô� �{��kg���7���Y���Ga�Y��*dܸ?��V�}/��X6իgk��ˆ(�d#0����'�k%U�K��/����]�m�+�Ckx^�����E��&�;,B�u1Flq�]���y���dB�Y9-��~��"�g�hvV��|�����,G����1f�@ �[�;�r�R6ri��}c�8	z���z9s�5ɥʨ��L�ޛ�;��X��5yƚ*���3�y���r�Ӂ�G@�:���z���G4lyKv�t1���Wrؖƺ�hw+4��R��uݙ>�J�h��ãaz�����[�v�>�[!y��qn�iJ���5�H�v6ح��'�kB�c�ST���� =JS*����sOU���J� �#����JR���:e�h�ڬ�9"�W�tZ�.:��PZ^���w)s|�R0��BVf�:._\�+7�zAu��Gkl9e퐁w2��;ŝNr��y��� �v���vQ�‮�T9t"p)��Պ�Oy�N�USo��r�����u���(D�kb�y�Z�#VVC;�������Y�ʺ����])��dA`�8Ȕ�l���P�v=΢~G�e��.`�x������5����f���ȱ+ʺW���9u�LX����v`�X;CO��{��)� ƕi�I��O�]�-1��9�'�Z�q�΍�*�F��ݻ��u�p@�m<��{z�]����h&�m����:��T�x'�f�z�2��G-l룡.�E���9t�����黻ׂi��!xlr����[�msEƥ�4CR�we��9{�L'�,�Sv��bgC���ۋ'_^N5�/',�� ޣ[œ_R�Q�;��V�k��O4\՝{�p�Y��X��;NTU�Χt[�7��*�����0q��0���S�$������+ �
�-��+/����x�3e��R.��r/�(����uu�Su,Q54]IB =��ReУ��t��ӥ�_k�vY��V�y�o��kH�q�$�G'R�!+噔�����Ҝ�v���$*�K �]�7Gi��G!#�uS�s'�G���p�һ��0-{����u�[����K���o%�d'F��YC�A���᢯�qX���[�B3��>9ٗ���1���.�e��Y��T�{q�R"v ��ج|nA�� �;�C�B6�6����5+3��{���y�w��f<��I$�!�C�"��e#��h!��=y�_���#k/_���z%���?��K��yY��{��*�ᶧr+o�*���
�k����ã@���W��#^�Cb�6�h8rA�]�*2uV�f9�bH%v=�������e1p[��7�员�<�F�x����	��Y�U�)�4��A|�
LU)M*4Z����	�$k��I|EQ�����Oʢ&�%LH�6
�$"P��4uM�RB��dtJ�ܑ�n���P3.#c쪭���N׹7�(�v�����C�[����`ؙ] ��N��偐~B����H�l�X������n�|�n��(?5��.���	�῿�
�L5�{�e!g:J=��ǜ�M��Ł:�ݸ����yY�djJm���N%���c��,Q�i���	��m��{�߲�5�J��)-�J�9�7Cu��1���g����:%�έ#��}�=|�k��O\s��6�j�o޽�H�����
h׮��5�����*��!����fz��T��P:'u$Y׆WmWZ[gqA嶦�s�ܿff��g	�l�s��V�""��%M"�i{�s�����(GD�C9q��r�+�9o�mH�I�9���i��t9h쵗�>��$���#�~kϮL�.����ps����w���h���Go�BM��ׅ�
�B�a���𠌮��<v�KQ��Ű�R+�j�1׿c����nue�n���0a�q0�Sǉ�"���]@���� �re�$�J��z�}�>�� >�����v G���򛲊���V����\WA�k��ql�Ot�sc>�п,�s��c �c֪0�s=7T��c\u�[��h}��<������d�:vy[k�0PT߷B��;����<弞ݬ5��!��]���:�]� ��qU��N����{ޔ�C���5旺���hĹ��l^�ө�u]E����v���=����&�	��ݿM�o��冇�R~��E]�����2I�A���{����J$ӭ%��ۦP��]]�C"�|�5km��ջ��,Z�Y;u��/9Ұ`>s�����0v�/�a,ͯ����5�����o����G0�Ǘ' ��v^���:�]�=g9��z�+D��R�6��f*k�{�ٝ��*IR�����T��U���dH�PO%B����n���(bA�=�3V1��M^��4D���T�.6-t. Ll�VƔ���|څL���on��%@�Q��G����Z��}�ޞ����cW�GRP���Dc;X�����}�Sj.���_�?+O<50�C�e�j�W���Rs�3��f����ݵd��_v�t�Lu����3S<.f�1��^�NP����d�x�����}��;�T���=�yx���.�)%f��n�V]�*x�A��2	�B�d;'�@�6�˹v��MP��y1�w����r8��N�<�fYa�u)ӡ�Q6XpQ���W7Q2�``ms=�T&�	Z�J�n�9D����nS��J���t5�#"u%�(�]vB��c�����a"���FTwuW%S��UR.;��.�����It �
���,�b�Qc�
 R,uM��T���ېm��1�`�`�2���ڿA��?>kfup4[�1C�G$sw�+7�i�G��l�~9�}����s�`izW*h�����ko�˳�V>�25�Uyk�=��C�,��^/(�H�s�y��2��ЫMmD��]�SŅxp�bR�ju$'z���X�W��ʏB��k@����v�����s~����tϭcHr�^��>���/�<Y���'k�'T8)�QPC`ي�M[�7ER�fT�u�$��/�b���`�Wp�Q�K1@%�����O+̢�H�t-�4G�I�u�=�a�ͽ&�u����sr�g�[ɳ0\�i�-am����``��F��k0�Dy�زU�V*���}�zR<wt,[}�����4�� 0Ш`�n�<�|�:�J1q���i*bFح�-���`�wX`u�/���@�ᤎ�B� u�Sӵ�����:�g^��e�#�#�9��A��ALH�K�I�FX� �@�01��-$F-#�$SI�M!u����H�TJ1�^H�@a��xhJؖ���e��	��BAM,0A��4���6�0E�/��,Km*��q�#MQ�Zb
a���ZH�:Ѷ���H)�h����%�9� �ї(;�pg�{`��o'�Y�{�mv�j����W��S@�i�
b{���a��#6�E�
�H)�0�(�TЄ��4���A�����*���3��u��:����o̔��ώ_��K�j��F����]�tޞ�Z��Wi��t�,M�st��+u9gonR�(��ѭ�=yy׼��wqK�pK�w��|���:�����o)a�y;���=��ʼ��!ϓ�*��$����u�U�D��,R��D4K��{*!�6�m�-��:�ſ�<�O�R��ܤv=_��#;��;���Wۖ����Ee���Ƒ��p����5v������2x%���g�)�qǑ̽`�<��X�wH�J&��{������H�q	=��V�L������n׵1
�a��ҋ1�c��[ú���<fv�������xk��t9��×���������3or%�&].��%a�W�����S�{-O8���!�~q9o<��Û���-I;߂h��`g+��7�ӏ���_i����UT:��~�F<���7F��蠘��j[��$��G��{���^��tj��TҸ��\(�1�Z��(\�]� P�e�'��CԨ]l��ߞ��h�+1�G{9X^��}'����;��,Vb�;��5����$>�	V��J�P�:T,!�����4Rd1�k��]�(��~�,
���h��Ԩ{)�rk�T����ɗ_���/��;�\hg6����]�u¶��'2�ns��H�%���=��^Q�;��'.��BT�Q��f�څ��Z�it�u�$]S�	�֑:�ViRm�(��y�ݘP��Ԥ�mR�8������߼��H���+�]�'d^'�^k"�WA�`Si�ώY�2�(���f�!d4(���$�I�!��T���3ZF�w�tE��H�B�5��-�i�(�
N��(�G&A �R�����:����*(($A��K_2T�4�䡒17%�#e�r�wv���a�S�W��:E��(��(R��&X��DQ(|�	-�h�U9%]��N]AԺPd��UE���ը�R[�]��t���яz>3�}�+�\*��V��~Q�
�;ݘ���2��?k��Qm�� ���MՎ�o�rq�����M.Z�ٹ���_$��݃b�w�fP�t��4j[���&o�ٳ��4��u�wj4������k�r���GN迟}�}yF���ں����d���+a���m�s<�Y~���1�P-�G֦ͰA�G�YA�E�,&�B��{�|���7�$WY��旚��Z��9���}��U��?�^�6����~���yM<1�+L�B����f�x�8 8�Uܵ��Y��Ҳ� �}���J����Fj�g�r짶[=�;��(��Sm\�[�Z�^D�~��������W��*�E���w+<�r��L����mX�.a+Ɨ��۩A�k닟���B����h�tV�lk��Ocm�;�A�=�«ȫ�zm�eXҮ�}�c�ƒ���_USSN�~s�;k˛۴F�A,�6I����Ś9?4�M��[�||�<�e�(t�\��d�����2�k��C����6b���w� �G����m�\�$��ܭi]��"#ȓW��LSw1�ݟ{ln�M'QQ�&	�!�N%o�mи��͉O�;�C���/�W?^˝sƁ��+5�}�Mt��;׷�Q�� nbb�IMN<�av�9ꪯ�d_�Ȩ����e�����x�u~�޶8�	�X'.�f49��,//6����5���e���n*A㲆<��D-K#�s�z����V�}�*n���<S;�*���9�i��˝��}�U���H��|0��6�5~��!�TEG�I�e�Ү{3כ��S�Pؐ�jE\ａ�[�v*�8t�t`��ޡ\}@�f*�Ğ�n��U}��S�7T�}"�ǻ1G��Y�mA��
UN\W^L>c=k`t���
�9�ǡ�\���Q��-������%�j&j�tf#��7��#Ż't�I?W��V�B׿V\+Xx��H�w�,������nv�xj(q�xcD�Ht���1��uLf���C*�[,Vf=���e����[2Я�^$JS߫�����ڸ�\+��2��V�ר*GCz�5��XȐ��@M���>5�j���N�q��.��H �y4֮���g���Qf���l<�ah�h�y��kCeS{[��,�L`\�PypR۽�Z�4��������N!��(�/5� ��Ҕ�ݬq#�����`2��0J7o�5i�u���J��*����-J����,��*��Vނ�9�bE}d�qb X�l̩����@YL�U�j:Q��QS����\j1�lu��e�F�2���J��� hH�D�Q ��I
i*��`]9r\R�wD.��7Lu.�t��6��NX�U�r�HBU��r���bd�135Ts���]���4����걳�,?"���9n��aO,���YO]ۼ�&'"i��j�<n�iH�X�f�����v�Xr���"�aǌ��Fژ�q���n�Y�ɫ�h�]e=������2h���u�L�Y�F��V qU$VՈ�+r��M�q��'��sם�	������}U��Ƃ��3l��.5����;�U�e�r���i���B�7���f����5����=�^"�+a�)"�5J2gt�������*)�wqk16��1�Xe�b���_�f;�c,NCMe����j�rհ��̲<�Y|c�f/y�;��ռ�:�h�S~��S�2�c���^k�h��?����3L�Z�Xam[<3:�m�MSYh��
�-b.����Z��S|�)�t�i[Z�^+W�r���#�4��]D<h���)���k�Lm[�X��2̽5WZ\r���]1�Y�+i�Pc����5�>�m*���>9�);�%��Eꪯ��<4FF������|�Y˷�V�b�}f�Y�)� n21�����+�q��,�[�V�4ҍ�I^Ђ��*�ҿ���|�R�K��e�U�Z��Xsz�u�ykl�3���3���zh�
e46�w}dyh�\bU�b�yc-_K�]��<1�%�n�/{�M�޼B�r�L����6�n
\&f�)�xxe��kwY����L-�e�0���.�l�[b�Wx�Y�f��a��b��9�-*���Ŭ���_Z�j��:5L�<�V�S�+1b���xާf����zx�Fw��g9��a�֙��jS0ͳ:�L�ʸv��;{��m������;|3g��F'�HH�^C�(��-�j�]�Y޷&6�e8ճ</6[)��)���[���k�J�ƺ͏���#���x쵦�k���e��'o�'2e�4؇qm��5|k,�&���>sx+z��[0��\�{��{\Gq2��=�+zcce5;]�6�x��|��.n�������[fs1ix���kn�}x9	��x�yci9	�a����9�`i<D��鮼���9E3LlCh�`�����i�fy�N�����F����sr�t�ї���b��\�l��!��e��(ި��D]��n�6u�ਜ਼9����z�hN]f��}%�k��L����]-�g����3ƹǷ�����S[b����ll�p��-�%3��_9��A��4W9J�y�w7�am�kM|f^^�+pf�M�3��>rR0�6�e��C���4ц��v�Z��aL4ҍ�\k�l�q�a���I:rE�쪻}K�!T�*µo�y�zXgZ�/�Z0����<gm-5���)��12wX:ņ�5l��/u������Yw8���j���3U	Ƞ�ǆ��=^�phۧ�[��+�*v�1�da�MB�XS���k-6���b��3�.�f^Z�16Gx�������X���������H>׸�RSįl���Y|���K���Ȉ�����=��
`�S�G�q�3�5�Ҝ�A6�c-���y|f3�E<��y|��Hq���Ì�:����K���ta�kF��`�81�����^�1�df��m���^&8e�+y|gT�5åbY�b����,�`��Û�L\t�X���HkȨW7��c����L8먩�nik�[$<�W.��� w}:s�.���1�Nk��=�{}�%���ᴧ"�7��YNI�6a�8���r�E�N�!�ڳO��~ö)����pk����sz�G/�Ӌ/��`�'0LN\�ƨ	f�R�5�ӥk���gj{�(��'^�k�6�J��bT��c�ܽ�u;N��P	��u����k��$��޳2Wn�|ֶB�Q����ή���҆��bd�o �B��|�Օ@P	�(��8۷#%R�Q��:d�u �5ۍөd����[`�9����WeEM�E�[�j�n���Cm��i��%�:�K��t8�)7D�!��mI��E�h ������o|7�o\�"��H�^U��;���L˦[�E��43�Wp�!�ElV�#�>%�h�!�Coz�ޘ�����a*�����|�&����df�#�#��c��c�7��ZiFm����q�r"1��#0�ܪ�9�o7�ln0m��[�oY4<�29�MBb#�/�l�u�q�D�g+�<;��� ­g���7�s~B%�2�<��������Y��OLu�[.���׌�m����p�V9�:�4�Z�.k�Up��O,�M���ּ���7�me卫kS3kl�+]��E�����4�m�:�-S�p�f6���ݺ��N���HW�p�F����ϻ,�9�t]�Q�.��x��U��G2���~���)������R���q��F�����5O��/��ǌ�Ye��}�n��K���f�;N�l�<���d%c�i1t�������Gv��p�a+�K�C�=u�:�O������ܢB�V����DDD��T��~ﶤz7�@�D�#K�Z�fE`m��_vo��X�y��B���ǽ�v��W1���9
�Ν��p²h��Ld׳�b������9ù!�\���UU����*D?�����S}}ك�|w�lڨ��B����vGkco>⟄��^���J=D��z��9�3������z>�<\U;���HaUs���%<�g���ݫ��" �gؑ�ԙ�B��k6G���[������(u�o��+2�֏T��10zꀥ!<P�����J7T��k�[�5b�}Q�,=�h�!Z}���"���]����ʳ���A����3�5|l
z��"�I� �H�y.��T)NɊ{�6����²$]������McmJ�8��\��I,!���ʼ�CSI�1n��3{����Un����F�TV��xڕ)Yݢ���2ּ{E"ԛU�Ӵ�����&�ya�_v��\:ͩol�m�t�)�-�4���,�iw�:�I���E߾��'��|�߻�(��m���CD]旅b��K��{Xõ��F��$;0�t��0��l]���
7��og*]s9#�wr��e�N��yӢ��}UW�Q�����!���,��8��BbE?W�]Z[P���1w��ʂ�v�Rf���5�!l� �ץ+gy���W�c��&]<;(�x�߲(�R�W�:��+�.����q_f�aQ|Xͬƺ<T#����˜��\�VV_Z�p3v!��fY�KB*�+�8�T2K��t7�^�R�{劸�Tu�	�'ǎ#��,���Np�a���9��la��K<��ڛ!�H:���/x���K	��u�dy+��u޸�oRfN�aW�6ۇiЌ_dT�Ԧ5��愲����yv��Gڭ�]�]�Okaf6�U��L��,HD�m����d�v:p���d)���'cM��D� Ċ"�FA�%5TI$*U0�*�:Q�F�Q�S��8��u#��U5)�N�'RP�dh�!�rcDq�Sn8ӧe6���c���{�듂Z������򈈫)2;�)5�'k;��	��R�^l�˛+u�ovn}��w�&{K�2�4"�Ciy4�������V����;:U����]P����|���E��_y�	��!I���{���X�z�����GNcA��X�;z��XlI�^��6�VCFX`V��:��u�r�w&:'&�mά�j���k%a5��ܘ�-rhξYR�V�����}��%�<�?+��dS���j�����9���]�Ӝ���a�̯)��v���ʻe��	�[EU�e��;d���A��������9?,-�#�Ŀ[�����U~u�/�u��'	��466exJwK�I+�|$j�{%�߭rk�r�ט�g�*J�bzS�4���h��|:��Q�N&�_d���}��>���:��, ���S��܆�e���u{�X�y�wĿ�})����U��V�f�U�Ef3%oP]G;Ƀ�@qT�>+B��%�X�e�������:QN����ݟ�r����i��e�,ٵ$_�f�}%��v��O�Ͻx4����k�����6�f
���ܗ�=ԎyHw���7U��=R�w\g�R���}�j�l�\gS��{��R���N�I�*E�׿�Y�;t�~��w��n����5q�@c�[�x!]7F�o')��[���)�z�C�50�ufnD!�=W^y��k���~��<ðaLK�c����CN�����E�=�"�sK�q3/;� �1iR;*x��݀	�j��E�1��N�Q3�Z���|+)��r���&�w
�r��œ�{�h��$�}�rx~ͯ}~S)�N�7XZ:v�4�3��C��GW��C���y��۬8�y(�1��۬�Ĩ�{���0V�[�}��7Uf�+� ��<=)]����\7w;�<��$�rp�Y��E�Q5�` 2h�#��B�5�u�yYx�k��L�VI7��j��-�{��s<j�F�tO�e��5���*z(M��2i�iu�{��Ftب�֔X�hDʛ�^b�o����v񗳚A�kA��ܜ����tWRo�ͮ�.�8�
�������1p+�
�aum
]}z{+���B̏ୌ��1X�<�f7t)G�<)̼r�F�8��Q��j����0YX՚b(6VQk(�)�P�p�UJ�1i��Jm�YH��3D��pwZ�Px�X��J��a�V��� ��̏�tA�,%�ʒr9���ջ)�5���
���%Uے2���6ۦA�)��UP�eU\��:r����86B�UD�M���5N�#Qґ�ٌo]���R�I�	#\�\�}���}_U3��qYB']���B~��L�kB����̞�r�&y��ˡ%�ٲY�l<LKj��;�۬�gr8��^�Qwu?A5�������^~��i����U��~�xk��g��Q�M��[k��5��f���f�ux�'P'�ؑ�~���ޮ�;)�<��L�y���.��A�:�t���_U^��4W~�f1��+ZSf����j�Ƈ��'��	�O�DĦV�f���Wۛ��+�YZ6Y��@"
`I;������6�@.�l걺�k7��77;�}_|���?����g"���ԷO��G���uHj)^��Tʖ�o����PQ��զ�a��^?eA�h����*?)�3�,���t���?Oq�+�S�k�}��^~��if�P�F�����s�t����	e�bU.�Ow.K��V�=Sŵʴн��_��~�h �Y��P��7��b�f���y�N��WN����� 8�j%vn%^���P�k5mC�y⨨C�4Rݐ;��@R����^�w\���˯r��6�=�o'i�ͳ��>�5�����ʝ��˷���˝.��|ƒLݍW�P&ƝCm==hl����Īy�q��{1�q-���7ޚOee���ߣN6E^�v�Q}k�ѿWd-����!o��t�Sݍ.��sJķ���3�W�/(��J�cg<���c�iM���#�[(�N��)m�w��u��e�׬|bY�0�`>xV�����T�u�ّ�`tu�1��w7�	T�E.��F����7H5�y�J#�w(��o�T�/�����{X��s�R�JF�fᕹ��[ڥ���b��w9d�q�keK�`'S�k���Ժ/7/��^2Va�!5��z�"nrA�;C���ٵ<&�Q�Mɋ�(���+{��V����k�%�1��z�m��r���K�w�}﫺t�Qr��ۗ��KbV�vT���Z .�s؍�Yz�2�*�\9���a+���i*��WI���#v�P$5�L��釞��|�	����6gl�k3�a2��L��n�_`��K��Bkv8�������mR�b`�ɀܹ�U�������(d��҃�X.B~&YG�l"��@Ł��JD*$'kf:�H�ʂ;H���,jS�D����/MZǚ5iӫ�-5���t	���	�L�¤*��R#�Q�)�6��UR�m����*m�m���!uUppnFҩ܎T�"i�ۻ�i4ۧ#5U*A�m�A� �)�F����n+ow���	�^2gcd�[��Q�9�C�X12����|���Cd��vG�ί)�v�
��*8�]�*���yy`�,V�u�j�Yc[5�ʐ����m�]�$KT��h{Ӥ�<�ד�{������*ҽ��ǅ�~[�|U֏���w�WPƒ��U�1D��h7�vj�T"(���nx�[]��w��o��@�^c�0��K��6�D�'mѠeʠ�v��n#ELąﭱG�,�=2�J˿kk�a��������vY7{��"��������A܏B�����hV{Wϩ�w�/��-����}fռu��,�9l�[���=�" Ϳ8��Cc~�aً�T�^���jT�Y���%��Ȋ;����rK�p+�w��v���R���w��⛹q��k�]ﻝbo���J���[S��1>�;�T#X�m�����L��9i���h�
ݧ��	�	�-��%H��y�	�#X��ޚaeZ=P��
��Vx��P�{鞛����+=~Ӌ^z�%�Ǘ[mF�ݷ��u2�!��M��9�kV��b������K��wT�u^,��"Y��W�h:��C�ksŻ���M�H���YƂ��Z�+����-DA�:zw��X~c���K�WB���7O��>�g/���؈c�:R:���[<%�v��
^f���S^��i�d��lC͌%�>����q@�y^LeoLM��2��J1����U�������K���]٧�T1����}k�^��,[��fL����\��'��J]B���^��cMqj ��L��N茳��V&q�Ch����l�աRz�;k�`�&�nE���N버�q#1�36{$�]Z�!UڕaZ�I~2:w]�S��1�'�/.�ӓ��-�8��ٓ� �:c�ŀ6�K�;����Iu��N����Ľ�&�J�ڷ{�kðL߯]��|�[C{ �����۩�M���0Y�r��,�Y]ٻ��0�@Qe��)n-
�b�UF�Q��nl]y�g/{����g"����4�ѹDR�뛀�ó.��T�ced�L�W�]>��<���܆���7̫�����`6J�)�4�b�2�;Ʃ;�T@FTf���Ts#t+�g�n�K
���
�D�V�uv�m];�7b�U5�qǔTNT֝�^�"i�
$Ւ�H�j�N��$�qF���.���W��!wVꪙqT�c�weB5W�I!*"�
LQ�M"�$  RH)?'[��f���E�Iv@�K�7VM[J�{g�Uֽ�\D�;-q���J�n��2���p��+*�e��`J"�/�<�.⩅@�r�������f׼Y�t���5��4�Ba��N�;gkj�C�D����N����^V���fP�yO/_���hw_�l6���in!-Õ�{]�W���,��w�;��u�`����;�������ҽ~��v0{1�\�H����z3���)z��b<��]l1�FƠqu�����D�G�L����nԎ���j]�\9�1��0�SΙ����T�d�/^�I��5�^f�������h��M��[ݩ���%B<� ]�:�.���9�P?u`C�÷Hy�kKѥ�T=�V��/}7#�R�]v�F���$�Gw+ZWb�^ޑ�a8�]ň靯7��{if۶�z��j�r�wF�P�5����J��S7�X����}6޿K�u5Ё���s�?�l�v�߸�cѳ�m�0_wRȐ+&&�7y�$��K��뤽��,�+x�+�fp׊{����*zɈ��W_w��emڿ=]m?����ݥW��u���N������=DQT�)7�i#�1�j�9����6F��.�L��Ga��V��^:�^�������J\��lg�ĸ3�q��\e��ax���l��� 8�\Ǧ�ɸZ���np���ȼ�z��s[�M�(]\�EK�4RoN\J/L_*n����ąZ�5x훣��+V6Me& [��=�_�R���)�]��Y�dk�b�]�3{���P�|~6X��{Vmv��'�A����c�"�F/��L��t�5�xb������t�O!e�Pf$�ڙs����7�R;5k#�]5�v�W�$Î�V{���}����mT�i�`��f?��I#�c��j����������q�� �j��^��������+|��L�HY��Į�p�T��<wW����ͬ��b�a��%�86�t���!=N�hpcj�7�GP9l�>�O��)�5R��T�P��>��NY�����Y@��K�{��Uz��M�}4V8Wgh���g-������o�U�]�'sܛJ�s��g7ۼ �@�����/X}���z]�o{t���i����ϧ���(�ϯ{�c��
^�}M��^7\�l���mEw�z���v��$y���0HB�<M >�2�+�$)�Sm���T��U�:q�%���I#H�*7U$N��u*J�@�R�N���eT*@���e6ۻ��d��,�R6�n;�X,��*�j�HQ4!�Ei���z�ti�Nf>�;��Z�SV�m��It]a�5a�)\h����K�>1[�$�>��C��E���ބ=ks�l�B�;i_-ʄ���4��|W��lT�Jgn�{��=8����w�&zlOICY��Pk�5u���s�c�r��>�5����		����P%^Y���r�l��L:v�<w�xD�҄g)�b�Js�NIt}eG��o�c��}/�2nR����%�Ł����۷m������ZA���Eb^����f�7Ři�G(z=Q�h1G��y����ҭH��l���.���u�ї��˳�u�}w�ir�t~�^�[����gm�IP&��َ����\��w^Ic5�o�=>���\5{���X>�\i�3�u7��.e���vnʢ�q��C��1�y( �8�nf�K�Ϯ�>�zW��+� }��f54Y�����WF�B��6��z�����X��u�^�����fMޣ�m�: Q���pi������]5s�a��(R�Fl괠.�<.5�4/vℍ^�����r`m�<����=5�o�������>czU���}&�k��U��lY�!s]5��*VQ��랠2�Nf�*�6�u��e���>���^\7R4��f�R)A�k}j��+GV߄�wu'(ӓ����-J����Ztt�Fq�4�F�[i~��Z�ӴGfYqp��v&�����0�p�4��{�C�j���U�G;���W��y��[�"�6��a>��|xOP���]�ׁ��3���c��.��d�狲��cKi`.F�yb�Rъyҫ��Ǣ���M�OkZ���b���/�6h
�ޤ"���m��H�S�' ��*]�}tk �y��N[����:�������M�v�7H���Q�+��]�|�l�9Xҋ{�b�4w�>��}��}cl��8�m��މ  B)���� B?�p #¸~�o+�$MK"��[!yOU�K1���l "���\��i�0f�e��<��h5�ɫǝ!d0�S�?b=n�I$�p�ߛ�?_���g՟�ثK��+!�{lt{Rj�-�5�s��5��j���{zI���Xҽp #�#���y�~�?� a�}H@G�,�@!��&���x��=�=����A}��0C��V��������_$���  �o���ڗ��4��
�#b�F>�C�����z�C�?2b���a'�Y@�=~�����>a��*_�fW�b�/ᒀ B0���S�g�Y�I E���,,A���iȡDǜ�JU}����<������ �y,��	�3�G�ǰ����Z ~ό[E���0�"�y�$�����C��>�z��^�j  �c�Qv'Iz�G�~���|C����p�z��)u(Z��'���3������`ܾհ���������ִzϒI$���4���=�mO���7���?��Q��{���'K� ���ͻ��>0�%�B���E�F<�d��$�FC'��li������#b�z!i`����{hd0+�|+�C�GϽ�A��R�h5M#�1��A���������x%�G�$�@�C��LC�/��kG�~�!���������z��|����=�aC�>���>��~(�Dq�E~�g������I$�#�5�Y��&�HD������?�$�@����֞���G�s������u�y/@Ty���u�45�*D?�,cRT����b��/��が���������?�7F�:�<��焒I>��`9�{}�u�>�2���tg�������Xה5���l�X������h@G��%�=h����=K^�������C��d=��,�a<��ƃ��/�V��c`����A/��$/�K���H�
_�@