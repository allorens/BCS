BZh91AY&SY������_�`qc���fߠ����b%�          �                                       |���
Z�{        � ��   
          P    �     ���(�J��*�	J���R�"P��
*��%U���B�"B�� D %=��H I�
�T�J�!t��݇�w:]��J���Jy$����!��A=����$m���D9�*�����"���(   �O��iRI@�;�䯤ͽ�z
z+��J�ꪎ{v,��^Ί�j���:y����=;�A�A�G{�񵡣�;i��Δ<�s�B��   s�|�$  3��UR�%*EP�K���(ݻ�f��9��U�罍1��iT��;ƅF�=;�z{`�2��N��B^3-Q�t�EtzЯv��N@`   s�|�P 	�>� ><�{:�=��ϣ�{��n����3i���f{�=(��|$���Udg�h�z<�(���<}��� ��   ��R t���(
*�H;�Ҕﾀ�ޱ���*�G{=(<�rR�7}>��8�����^�/�7���_M4���UG�!��h�   }� 1�=���	�y� 8{��< -o��A���ǰ� =zo{��pJ��Jл���T�N��X�f94�8   K���'D�#��R�B�BD�u��� c��P����b�@t�gz��ps��=�9:QC݀�:�GTLqUR�N=��oD   +{�jU �����݀:�Ȩ��9E��Awp}���8�U'-= �`��n�ǳ���@  P
s���(  ����DIJ"�E"��;��J�
�`9@Nu#���4�9��}=�u:�WӦ�p   �Ȑ  \}�|�w�NqJG [8�7`�,���F��!N�&@�T�h;�@{�     �`  �"`R�5d`L LM�=i��#"��       O�*�?T��     ��R)T�       !$�Jjj�       D�1��$��54b4�i�hM4d�'����?l����-�_��'�f��{i�� ��� V�PT�P_��@W�������?����WU?� *��}I$��� *���EO�EQ������)�W�1Zb��3+�\��̮i�3�29��.ds+�\��W29�0��3)�C29��.as)����09�̦ds)���@̮`s3#�L��G09��as�����S0`s)��fS09�2̦`s)��� �.es+����0���ds���29�`s���2��̎`s3�L��G2��̦`s���S0��̦e3)�L��S2���a3��#�\��09�̎ds���fC29�̎`s f �!�\��f29��!�2��3 f��.as+�0��̬�a��3*f0���3�\���.es�\2���!�\��@�.as�	�̎`��G0��3+����0��3#���W0��̮`&\��G0���.as���29��a3$��2���.as#�����S29��e3��2f09�̎e3���G0�`s#���G09�̎a33�\���ds	�\��&S29�̦ds#���G23.as)���0���.ds�I�)�\��W0���.ds f̬��0���`s����.es+�\��G0ds,�f �.es+�\��2����.d��W0��3(f309�̎ds#�\��G1�I��as+���G09��d���S09�̦`s	���f�L��W29�̦e3#���0̎ds#��f0���`�s�L��2���e3�32���.es(fG29�d3#���G0��̎`s,˘��0���&ds#�S09�̎`s�L��S03�`s�L��2���e�)�L�fS2��̎es+���fS0���.`s��L�̦`s)�0��3�&S2���ds�0���$��0`s f�0d��3(�̮as2�0��3�\��W2������3�\�� �.`���W0a�� ̉�\��f@�.d�������.as���� ̎`��2��̆`�0��́�\��3+�30es�0es�	�0��̮d��3(fL� f ̡�c2d	�T̫�&0�W2*�Q\� fD\�©�T�Us �`� ��W0��\«�As .d�
�)�s(�`�(��0�@\��Ts
�aQ̊9�W1�fȣ�Ps".dU�9��a3)��2�2���e3���0dfs���29�̎ds+�\���2��̮es�\���3f̩�\��W0���3 f2��3�\�� ��ZaL)��*;���@�?���l�5z�_�� ��^	v�M��Ȇ:�D��*�����t��3p�XDC� YY�^�Ȅ�"T�x�;�q*ٲ�';�'t�����5.�:���v(� �{3@��/a
�w���H�"K�vM��3j��Fk6��ՠ�W�6��cr�7@���*��mm�1z%�����T����Wj��H0�tO_��)�$�0��,�[E7N0�b"����*ң�l��p��z�M��u�ʇ͑��N�10��tE�4���Id@v�M���e빩� ��o��LZ��T6�e��N�������H��n��
�*��,���G�M,a�ӂ]�oX�@��AM,D�PPw�Yr����=��cݖe�D�*?],�q����x`�웰p]ScA�9Oth��My�,�#�n�K��UҼ�i��)�k��N����ܺ���%&�5
#5����'t��2�i�1����qHy"��D���u :��mŹ�3Cwp˓i���NHnc{�ҡ������0�X��u��f�Z4-��ۼԚ���m�.�h��V��"�Rս%��͘�@[̼H�f����j�sq����b��7��䣐��q�훑��{�aT�$H����p����d�sr�f[U�zE�����{7L]��Y��ܨr���Xs�������Gi,̄i�vl�-ZhS[��#� �i���]�<�5`���:ԭ2�60#��
�,�+n�Q�B�a�[��z�(�#�׌Lt��j�$@<�P�>��؟��wg�[�۴Fh�"��T/p�!�{U)KB1r;Ʋ��d��=�{�Ww����}�0nݝ�Õu}�,��KTe];��b�1�jb6.�ʚ�`�n�q ��e�N�
�ٛ)l�ַ�X������ސwV蕆m�%cT$%[׊^ʷ{0ˬ.�'�j�*8]�Tv�6��TH�B��m���t��*�];�@�*ޚ6{�TX��v�b�c��9�Em�VJ�`9%<X���2��ɛ��Q6���fm!��`�P���ܺ�`����{n�j7!�,ڕ�C����F�5�lJ�L��ZZ{��qML�ٙb¥���cFo11]ݠ����{r�n0�ܞ�7�vu�0�v74�؛�wB��p˷{4�����MDԢ�*��oې;-��,�0mji�{Z-�Yۉ�9�u�����F3
F�̺�+^'A���V��E��Z�Ja�b��{[�e^Q�&�]�d��D�[�l��j��I�7@�Hi�� �VšK�5&�����'w�PSoe4�8�N�M����zQu �Yy�Lh��#�ݥ!������˖��<$���Mfهr�6�k���r�a*�H-�-�҆úZ�6��y��X���Y�ts]���6ٻƳI PI��+���e�F�L4b�j�<(�r�<4���)n���g.�8�����F�
0��F�7�V6K8�&wt�!�b��l�˚�׹q�ȵ�9�fm�Yebn�ݻ�v���n��$�cF�Z��`����2��,W-�@�F�r�F<0JH���ɷ!܅�)x�xU�x,]^�)��u1ܧ��[Ɍ�Ql�U��w\.�H,xt-ѹ�+��d~�����e��{��N�1��P�.0e�u�5֚e��9hD�!���$����f<�ˏ/��.�VP�w�
�Ec$X��Fa!S�qlf����J�/F��1=6`Ñ] �`)"�X -+(ĕ�4�횂��1�	�JVL����t�A��z�\U�n�ni�Ħ��E0�7�:g&!��")��;�s3h4Ƚ:ֆ��a�6`sP��)`,fn=Z�`mi��sV�V`�kI�X�oB�����b�B��g0Nލ�u#YC
���o�o.Vl�$��.��������*�]![�EJ����2�=,��7�-�=:�HC3���)\L�e��ǆ��v����f�P��T^f
'l�Y�;��(�ux�_�$б���X��7P�,TàO ש����dw�؇Vܲ�6mx����u71V���(���k�PV��^Ѽ�I��R3P�y%�ܺ���y�����.�I���9I�ۛK)\8^YL뺘�݉d����@`v�G-�Pc.�X���N#��	�15�໐�ə����%IH���\�U�Bƥ�`k�y�J9�2�J�wtˢ]�46)�Z��h̢�U�픱�����,Y�m�t�QLksP����fZ����&���n����k/X����>	+�J���:q�ܻ��+���N��ͥ����:h�#��C	I�l�enb�B��MD<�œe�ט��e۲��V�5�i&ޥY���a�S/Me�y`ۻ&;9��њ��V�;wx��Yaa����ș4� ��&�~��XN�/b�;u3*��4���"PɛM	i^K���Kŏh<��r!���F0��Vn]����!��{.�t�l���a#t�%��wD�
�Y��d�׃77̩��&�T.�ǘk+pX��8�e(���Y�PS4㷇��/�X�D��H!��D]�v�@B����g��P�N<���j��@���ΦT�˽�v#��Ҳ(@�^�c;�3{�h��H�Q�u��6`W��F`x�����e��]�	�/%K��1 D����n9��#�m�6c��3w���D��CY���j����] 2Mq��+��q��)4�j엥��\���UZ1b���q;�k��<5�]6�s+b�h��<� �hf�[ ))o�Yi��v+t�me�3\�l�+&����-V�o`.�a�GF�v�/.�ٗ���	��.U����ݴ1�ubn�y@9��v�.���H��	Yh��`�3B�z��q�n˛d;j�jv��e�n���2X�a��b�=�eplz�Q�-���6�or�a����n+=v],
]�+��n��e��*b�7�-�Ai7���.Vܽ�X�Wo�m�FU��֛��7l��� �n�Mmв&]�o�HQӻ&ic �c ���=8�6���i*U0�U#0K����<	�����Ԭ���L�KVX�uA��3凭��	B����n��*�ІY{1���xܱ�r��!y*��fR�E=cn���oġ�vM-�a���xmc�[Z�$��h+5�!�$c��b^P�T�y�4Y�e%��s��o4n�j�u�\�w�y�U�9�X��JIݶ �j��v�ʻ֝e4�:��4�Umh�UנD&@5]h�E1Hc�
�R2���w�Z��[�田in Xa7JJ-�ǯ)�E(��r����G$�fk4��a�Y�e���i����2��]Z�b���nEt�F[[�Xa�~���ي�������*Uo�7mڥ%�a (J�"�O0�ٲ]!�� �۠�eE{��N�cM��F�1C��0̠ �W��Qؤ	�z��`ܗ�0�ٰ���Z�(8 X������%ZLI���[D
8�u����0�"5�Xe���J�5��WU�U��Vj�v*K6�'@qӪ�-�):X�Ր]b���䗨�0E6�qd�f�1�4/f�ڽkk/+L{f��0��m�Ԕͽ���J=5$�@FTT�̡Mn���c3T�	�,��s
݄:GN٤"�w3*Ьw�mn�*���ɤ�fB]���Ĳ�b��m�!ûy�^Չ����t�θnG,�j�b)��K6̡ksf��ed�w�4옍h�uB��[˹���{z������;۩z�Y-����E=��PW��M�|Zi73�w(e��Ȣ�zD��w2j6`,����.C�fdY�=�n�;*�-��k'U7<�e*X�XSI�G.��������m;����]��y)-Q<�b�<��dǹOhŲY�˽N��W��5P73H�X7���r�X���a��YoA��� U�nb��5����ͼ;�]%r�	5��,t2�Y��3���CR[82��j��{�i�p+�r�̶7�w!���֪4���k�XE�K��33mf \ˬ׻�҂����V���t�0���wv��e�s)61LDi8��3���k.��ۗ[��,�t �:7u.�kP��%�1�O`�e�y[y/*$���5���X�����1=��5X���6�Ř/ �Qshk۽�1�P�1�(�Xm�{J�]��J4�SaGk/niX��b��QL�{Vsc�YAj�M����Q�2�o+eI�Q���E�����TMG��N����s&�b��	2Gb�媃q]�)Q�J��6JJy�E�P3�Cze�܌�9w�EC�/N�[�xb��V��j�dJ8I����$iL(9�:(,���|r���Ց%R��$�XV��*�b�54m�e��I����(E��+{�[�W�*d	^�����ݺ�Jb��H�����,���v$�=�Cv"K��)�E_�0jGF+h��*ڱ�,��t��3Z.�1��DؑMŹMX������1k
E���Ė 0ʿe�7VJ�[0Z���[.(4H+0�9A���H��$)��)����#������Q�2Ӹ�0�<�d��:�Y����m���VqfS�n���7�Sܻ���t�-aVn��PB�w��߅�3��ws.��B�]	��$WmG[啡b
��vk(֔5�v}[f�nV�АQ@��Y�&d��Jٓ	��������@��)f�up�r�m,V&�%���z���w���ѭ�!@�H��Ⱥ�4��Rf3�{[�C5�U��kl'A� ��p]�����f��Z�ת�f˿1&ٗy����o�����b6�jő�� ̳N)be���i�
ݼi�w��pKJ^Q0:�ڼJUʙK�
���
�w*����t��Z!�L�o'V���a]c��Ce�U"��l��$���#bCE��4U����6
6ڽ7\xq*�1m�+I'/0*jl.�u��7nM�-!�����*� -��m�^�j���=�V��� ��1Z���l�u��D��f٦�R�Ri!��������w�H���l2�9xP��W��36����K)A�Jdk7;CnZ��p�a�K���{����oA0���3-�Kti4A���fF�B�]e�ݵ���]X�0��ى�ٖ=36�-siCX(�CH-�^ŕ�6���j���v\�.-��Zeb�n��7�S�-AJ���bU�V��^��v�p�i!{7FJ����[�Z��]�zsp<�s�\t8oF��7U��CjZ��x�LmP�U���F��]�U�6�C1��q`[����q)omL��V|�g��em(�%e�m�zF�4C4H�%*1j����)��6�uek�l�����/2�U��Ŋ3o	L��ʀS;���[go}��� n�Kl���8�.Q,0� ��;m�6��]ԫ��r��L��A�r���U��*z�J�Rܼ�,^j��0�Wv����j��{���%���l�{��QF�/e1�GlR�K�г0eL"�bJMeY�� R|%�ںyЫ�dd*�snf-$70^_�//v��SQ�\˭͒hy7E��6�<��i��ճ����[5䥛����N1��J��w+ei�������3��`ؖ�u1⣩b�7�=if�"�ہ�^�ص�A] 
	Z(� ��m�j��f�
���[��֞�^�°�5��C���x0ɂ�v"���Y�����!���Y9+6d
���pؼ�D�Lч���
guv�\��v��1����̸4�4��[$I<
-[��K�!4EӺl��A�yy��`�pO"'T��[N��;Jf4n��I�oh�Z��A[{�[ Ĉ1��dP2V^
�ن�É�p̅��ShF��cqQT�sD����$�E�h�;. ����%���շ����B��D��2���ҡR����3q�kR^RQ[˻sw�.�V�$4e�W/SQ��2��	
�*�����]��;H�v�����vF�����Ҏٵ��i�^�b�e3�>�ݻ���H$�,���v9xoՕs$�h���	:4�d��r�dF���n�����p�*�P'^��{MnXF��+G�p5�}�ܨ����ۧm�.ɻ��ו� �Wű׹Yv\Ä�2�+:i�L>��gL��]8'v������cf�KG�GFa�\9�(t�pT��h�IV���ٺ(�܅,���ԝ��3��-㷵�p����v�k��PTݼ˺�NvZ�ͻ�2hz2����Za�B��(��zv�/�Ë���6�җu�^�V�7h�:���s��Se��e#���`�)E���%����QP
�ؼ���.8d}�Y	�Q���*�b�7�� g�/Tlaf��'Ot�G��ŏ.�6i����U�	Zk0�v��4�eZ7k�|:�`]�k�w9A�¾O�-�13>�<�fL�l��r�B��ɤ`��X��a��+%��v�TS�b���NfZ%�PP��>$��a�\�򝘠�9��0�j_�C��E��@5�Xhm��`��
��eXT��ݬ���eX�c*𴮕��8�L�]f^��b�+?9�C�e�(]`�,=o,K�3�}����m�H�
���YJ�;y2��]e�<P�򵆅c��/]m ��pf������p�ʸ!���e
d*hݺo���H$�iC��v�#^Me�ۦ$��I�# Gw��a�c1�̡��	kIS��q��x��f�WA�oV�0S���n\@�Şo<�[Եs黠%�8�ŗ��ʬ°�m��nɱpR�� �8�N_2Offv<���9.�˰�����ך�Y�jnk\i/InL�gH�y�hۏn/fs`����D���}�,�D]��2���V�Ӭ��n4Ҵ�O9�EbB�M^�qT2�&ٻ�a��m��_<���ye�qd7X݋b�z�zQ e��wwFi���>Gb��T�#�]�z�O9O���_�7�#����/��߯�wp�>�W�AA�� �(T(Ti �JPi
A
h�J JJ
@�JUJQ���V�Z@��ZDhAJDF�( �T� (D
TB��U
)QJ �P�P��
T��D�Q
T�E(���ZT�V��P�)T�U�J@ZE)Q�EJU)�JQ)EJ�$A)�(Z@JTZA(P�� �B�D�(JD��)(P)
D�JQ�(@Z
�"�� Ȫ(��5�뺝�w�Jy���	@��>w�&�_��v��6`M(9��g�W�ե�E���Q.PDx�$�;��}!��J͕���g�[��yo�E��y���Æz�������w[R���Y�b�#`��������(P�1,ީ57��yslu�;ZO>9��z�k����̇�^[+��Y�����Yu�ĴX�W13�"T��]5'��|�i�>�	��ˤ���=gŞ��_)�7N/�ɏ�ylf:�����<�0�f�]hC� C02s�; h������f=��x[ͭ}��1��Ծ��(fy.��_!|l���m�g��y-�I�l��_��.L��ߛǼ�
��b"Z	�r�c�$�V��K<��zЄ���5&�Vk�LG�#a�g���%�ߝ�����r��H�Z�X�Hffb0\7C(D�.";�}�ۍp�b�Y���E��b�=�J��G�^+�?�P!˯���z�<z�}���<^;|͞��8b��$�����6�����C,��W�`jnfDU��y�(�.P�GB�E7@xX���h
Fژ�D�e��d��\���Ԫ��~j\+�J*"#��C��٤P�7��?O���?������UU��Y�0���� ?�~�?�������D�~j�W�_��5B��/�}�(��3Aj��y��J.T�-�Q���2��8��S�S�HnJT�u{B�i=Wi� ����㍋vѪ��{s�"\cs��hl횀���-�������遺�:��ȩ��k���$-���X����5mݬVn�y\��]h�!3ꨮ��B֗\�$��N8-=�f���$r��1��[�U[�m��YY�(���+ [��,X��Φ��\��쫱�R��"ٚK,�(�.���-(�Px[�)e\�/6�;���J�^�*�>�+r�^MV�j[G��%�{u�Jŗڮ�av�u��l�/�G��
�s��Ɛs�������5X�Wyg3���/*�n�F��Y�8���F_��s[�xpӻ�U�����0���bjl	�R�s�CWXk����-fQ�YQ���^���)��;�juB�.e��*T���Y�z'^<���S>�ۻ�{ ���8@�d��2�oڀSz܆�Uw�v���:��
�����m����**�U4�%{��UWm�Kʫ%ؚ2�'d;����b\]F���
��j���U�3e���Qff�{MLFX���>!Wb�п�^y�m�B�ª��f������w�*f�c)��٤�poQ����)����4V�T�Wu�j��"������E���󶮹	.P�������������=q�n8�N8�8��q��q�qێ8�n8�8��q�q�v�8㏎8㎜q�t�8��1�q�q��8㏎8㎜q�q�8�N8�8�q�q�8�8��8ێ8�;q�q�q�8�q�q�q�8�8�q�|q�t��m�q�q�8�6�8��q�8�8�\q�q�z�q�q��qӎ8ӎ8�8���q�q�q�q�8�N8�8�����8��q��q�qێ8ێ8�8��m�q�q�t���w��nI����:sB��zr6�}z���n���嚣N� ��t2�";�'y��`uA`
��|�����	���>��*�w��In�K׍�[�Ep� ��t�ͥ�|�\F��;�� �{(����F^�٪��{[���1*����|fR�t�K�y��A}�V�nS͖<�n�ZZ	[rξ�{.\��/�о�:^���$��-+�pC:5����-V�e^{�Ve&*�z�U�5^Lʗ��W�߼���9wv!�z����Цz�#s['�A��o3v���NU��BK��L�*��lf�9r�1 ���������t���&�p��ר��G!\��q�x����Aˆf��f_J����P�v�y(f|�e^@�vz��x�\v�1D�Ô��*��.�u��E��*��jP�U^�+s.e���MTn�8�"ܹX�#`u9�¶tV�x�4��N��U����NYΌ�޽�{��z�E]�sT�*���)L0U�SK����b;,^;�]�ę�m�
�ot��>�M-�����K�{6'�,���(���N΁"�&�u��Ջ\V��ѫa��ѭy���%�e.W��	��5��eS����ހ���"����)-<=z�1�Z�շK�MV��g:*��lEێ�2�z����[�:hB������b���aw1�7]�֨e�����/�n^����L��n�cV�[��[{[���J:��9���v�S۫�/���^�c��8���8�8���8�8���8�8���8�8���8�8�8�8�q�q�8�8��q�q�z�q�q�z�q�q�z��8�8�8�8�=q�8�8�q�q�8�8��4�8�<q�q�q�8�q�q��8�8��q��q�q��qӎ8㎜q�|q�8㎜q�|q�8�8�q�q�|q�t�8ێ8�;pq�qӧN�=q�8�8�8��8�8�8�q�qǮ8�8�=f�����yw+^[��,�wwj�8��T|>�rI1�z�b��C=ぜ��b�y��Oe�b��{
�\,fY�ս��>�Z�uT�A`�	�?^+\��mFv�'oΆc>�GWi��'�ճs��f֎�;�iv{]�YG���*���y/(��Miф�o^��vo�=�r�j�kءM�!�%w��,B��UX�*��o(�-Y��|X��,�Z����L�����!m�A����W�"���os[]Z=n����f^[bûl�ޒ�{��@(;��͵�2��.�8s���WnW	j��[yv�CT��e����������Օ�Pn3 `�C4�xY�ē�ځhz� ���^�`4FZq�6z)������b�Q��8�v*��y�;��&�6du�Ҹ����w��E���:'��|�5��4�,��C��ǽJs�m�Werޜ�u��e�������OEU)s�=�gm�Os0�����O%6�R�J�E9U��/j��U�O5���<�S���Nx�x�o�Ih.��� k�W#
�%���y�xn�n�@��y�;�N��ZK��)�wҰj��T��q`|`�)���#%֗�՜�V�����PqWk��˴�sշq�^ҡ]����N�#}�K�zw,�@��c	��X�<����N�j�|��[Ը�\��*���r�Ց	���j
�˽�JVRw��ߤ�ȧM6��]b�\cCw�*�5�x��(��T��7Re�|��J�����;���{SP�[�����;��D�=Kڤ]=U;'�VQ'���oxP�N��c���{z�\�<iT��yR";ª��(f-�}}�ظg:�JZ9�+�h<��mXLt �s��˜�vt�z[n�>6���AV�yҳ��C�Fj���U=F�;h�<���Jja���Cr��np�F<��m�����3g'e�1[P��cp҂,��5ډ�=*&K2!�����Řjk���-�|��p�`�� ��Q�/G|���<�l���e�P�]���E5��$ �nt,+ѻ�v������5K/)%�%�oc��f4�h8/�X�Ɨ|���O9y�/P=����X,�b���6 I+4�3��S�1�u�!0}xއ�R:�L��:[;/{V��p]9�ˍ����!�+�슗m<P������b�m��M��]Wa��[����EEL�!�tT�V-��tN��}����ә؁�*[�@�zﺳ0���\�<V��I!CJ��V�;�����j�E��Gя����W5-5oknԳ�-]gX��s�TEv���;|�Ț���\19��6���Z�-�1�Y����(Vsep�y�uW����w՚�gOQ��,,Vm�f��|�Ga��[��LWc�w��o-��TD�d�K��N���ر��+��+��C���LF��hu��OA�K0RF���-�׊�]D�ͤ��ipS� p��+�|�\���5TEh�@�<����oF�z���kGIq9��y�TN��:�/��:(6C����҂-Z��u�(�k4z�����.{zz]����TWR�r�L��Q�m�۰�=�S�/yp@i4B����[��e&�b�W��,ݴ����\%NhN��v�f�v�%�WA�����#ʸ+:���s�իS�j�4+2ֺ��Q��.��uҬȞ�ў�F`�6����]8�'��գ{ TF����q�:�hJ��>������%�/�����L0-o��N<��5U�3N�Y����\=YYW�}�tҁ��E�S�w����i�B��y\��XF�̼�43;��е^�PyՅ��%�xV�(��Pm�d$�޻�#[�2^[׆J�+�����eH7c�/4�����S�;�;e��#�3��;�P��7�5���n�b��r5z� �V�R�r�s�{�t%�C�wr�i�E
pr���NٗP\�͢l���j!c+m�C�ֺ직��U�����a*r�^���լ�nq�9z�NӅq�qxV0��x��o]A�waj�J�]�srW��;�(gs��U���;Q ��f����wZy[����j��Ցq��T�U�q�Y�]�r�%r�л�S���8�m�*��ޢn����o]�z}��eQVg��e�Ս=�Տ�ș��2���7����3�$4������k��ǋ�D=����
���I��ކ��U�f���n��A[+|�@kw�՜�V߳*��m����l���s�]��c�IM��%�tD}��P��"ŗEm�I�yW�w�AU������چ�V9\�{�xN���4&�^U�z\wm��]O6�+���a�}�x�"M&6u�uUr�U�0��qT
�\�#s�};�IG�{Me�xw0���2����Q�}fwmn� ����#�u���N�$����L7���n�@gpe����uͰ!�c��J�?[�hZ�˾S���I��3:�]��c4��p(,L�jt���GRG��lxӫ]\�Y�Wg3�L�*ûb�B��6��ݼ���U��f�,�^��1����kf�ӳ���+r�
�2�YFU,)2��R��]�5:/p@[ɶ<��JGv�qft�����Զ^o+�����L�o�cmhn�-��a�J���꼴��Tl�y)bH�v��}��:��kd����㎧[>�g�F��a�s�����9�G���T�l�|�$}�VQLʻ%�w<K2���"�
�x�8dέׅۮ��h��	�A�������oYh�d]����sf�磭�W�0���+��{w�w�%p�/��>	-���M������e(���\Z�f;��I+W.�oY�R�q\4H�u��)��a9�b�tNX���l�C���@R�ܿgx*㮏�F�^Θ�eܥ�; ���<�������e�D�)�������z+��Տ(��
�6�����W�q�s_!f��­��KF�DX���^�b̥AË^����;�WR�*�yH/����sl	%���8w3f��8�R�l��f��a ᜎo�`mU�m����s�1����wC�MۦfۛW+�L�:���8�K�sq��}*�AUO�.Ĵa�%l�5f2[:��/m�18�d���4&G�^��v����7�B�ݦKm�]��9�;���{kT�^il]uyuR�������@;�%��2��`2�����ui�^7�r�f��ޣ[��g3�y�y������춲��V�CS���mh���L���ֿv,���yK�Gr�� V�o^��,Y�+kx�d[�ޗ�6�8N��K�l��-�O�a���ae�l��˽��2���W�`^�D*m^�[�W]�b��>w!��Y��nf�_YD�'s����ԇk5�c8��M�\8,]����CRiUfs���,�k�۫���ᨓ�]n�p�Q�eARBV=���;2fyb��;�{gk0�����B���2նb�ڨ�Hu���r7yA�cgSLŒ���+M�\����]��n�[��u�3�wCB�.��:3eF�� ��x{	ͦ�F��q'���YX5��S�@u�YBX�_w]�
��a��ҵ뫷�o]�Z�n����nq���Nfs�ԯ/o
�j���qvy�U���釖�оy՚�!_S&ƻgl%���� dy]����8m�+�6��u���}�o9�i�Ǖr��^� ���D,pQ6;$�UVm�ZE�Ve_������;;p���Vr�o7��J�A�¯N������ms�� �Yz4e���r�e�2��7���\�W[AYA,��z����]��m<�gQ^ugd`�[f��*i� -�7C�|��d���t�5��W{Q<��QUu�N��qoQyB�,��}h*�4�)��hu��Q]��t��ȅb=08��y.���/��C�T�~�J�^K�Op�U\ѹ{�*��F�n�̱��,AmqyF��#s
*�|,0�,�@�e�N�ݳ\��[�kX�`R�k�X�WY�J튵7p�붊v֨���a�.RV�o^��+��o��w]&�؝�'5�^cE��.��e�	�/'�g8��1�V�'�����q ��X�7��j����e���s��S�W8��%�j�1�:��$�f�t�v\�yZ�s]�g��W)�qOjb�&;p@!w���������<@�	PKK�ecvE�H��ێ�y�K;�́��i� �vv7"�U�ܻ�l-�3; ��ʳF!�+!�vw}g(�w`ټB������vh�e��{�m�4F���}��JO*��VN�����w^��v��tz������uQޏ�ʚ��U��\q�ɴ�-��K�@�dw�-��	�yp$:*�J��n�	ٜw�6$r�-��V��d���[9qx�Vd�1�u������ǻn�=��	�����p�zT�*3Z��7`#�vLO�ۓC�{�u�7�ѳ�m�L��1W�
FoV�u��鍫������ov�3[Ǥ4+��=h�gVs X�ݙm�{+=������yS���k�}��V���E�������q�Wm�նܙ9WjJ�i�yk��RNT�+`N�=�]�	��,���;J`�M�EZ��p���(M��h�ǹtm���+��+n�t��5��fk���:���r�����$�ı�̷t�f*��)�{E�o��]uƐ�� �)�9��0��(�����8���^*���=;���}%᭻vM;�Fٮ��p�	��S�\T��v�$��c��"3:K� "Ļ�-��䓝+֭*�۫��tU 2iJev��(X�S�>#{2��V��C�x@�2),�2�9��0�y8oqݻ��Z딒jiד��q�뗖�(�Z����n���\;�w9�9�ޓ��O�j9��v�����;i޽�oziq����j]���Y����ɾ����1mne��JZ3�{e ���S�� �hw^g;b�%ݍ�z�X�o���V�EyҎd�9=ܽ���6^�+�t���Y����/;f�=���˻ڲ�n�cS�n��)�²�U]�0�lK��/5�]��=9�J�ҚȆ�z�]G�Y[i�oLCt�]�M�+=w���s%���o#��w'�p]O3������?b� ����������G�j���������_Ħ�H}��.;H]ll=z��̹�2ka��<*�����K]w�ƕ࿛��-}�,����Ė�U��A+�$걽:׍vڙ`Q�v�۠q<�G����v��kt��3�m��ѓ���;h�,�i�h*;@��u�9crn_8ܛ�8z{�.47.�� �8��&��
�"�3��r�]Bd#�p�H[G���2��8����;h��;��[,.�=���nn:�S%ת��j9�b={=7b\+^v�����vSb���v#��\���lk0B@���Sz�<k�37c���j���#�Z�"w9{��[sG�/in7Od�x�7Ǟ��ٛv�9�Ι��k���0��2�e♀*ؒX���Kn�9�$��4:�L��`]hM50�7U��v	��mH�M��\d9���۝�0�I�����:���zwf�خQ�T�u��2�Wq`&�XL��ʕ6�&٤*Zט�p�@�����nFk[j�4�m�d���^5�Dq�G;d+1��!�16]4lsv�h�7f�3i�.xǹ����u3�q �n;\\侮��>Q�F3BG�a��V�9��m���x��B�:���5ʾ�yx����0
��']�Y���zv�L��O�P�ě�_ ��0`��P�;5`��驁b�a� v��\]yZw���q��Ws���&7��O,����:�Ց"M`Yr��2�Tk��PN���n�4\K�w��k/'77C�e���mN�T&�%���J1p��9ĎD��>�h۰��n@̻�E�5��gU�#�(5���7g��v�vڽ�3ہg�[	��P[u\�qGͮr�ȷ8��uڃ���g�]d��nw�k�����;v�E�W:xM�V[�`:�z��E�[�k�<ڠ��S�'a�8`�U�V�Z�]�͇c����P�����]�������v��G����7:��Ιv�H���*�S���D�6�b�6�����.&v]<���n|��޵��q�pmc�1̖jؒ�J�ef�y����&/!O&�|ݨ⩞�X(�t�6�6�q��uګMf\�SK�^wdQ˂g���н}�h�5na�Ce�]<u���_0��`�x-�1��������J��n���T��<���&"2��γ��j�U��U�\�d1��IJX,Z����V��VQ���z6v882J��۩T�n��@�cmÎ�1�2C���|���8'Q���E*��u�;�u�R�f�u�ڹ�d����e��㋞��hiar:Z�Ƈ9�e�Fgsҭ��r��u�2�9b^k���2-L;k�Gd��v86���ǝ5ŵ�m�2��"�H�	����t����f�Ktp$�(��\�Z�\/[��CԶ�����\��ĝ�����ƅ��C��Nܤt��N���3�Ǡ6����U���/X�b,:�Ķgk��hWM'�/�w�o|{X�s*��f:D�j،�W�%�`"hE	L+��k�u�0�L��Н:�ptuK��	��1M)��GB��Č<;l�O�)���<���cM�d��wRnЮ5�Ʀ�,!,��1̧=�^�M�����l�=��b��AG��iP�lԕұ"��e�D�ݸ;O!�UЗ$A�Z J�z�����3Qxx�'�l��|�r��-t��ޜv��Ġ=�
.:�0�[5�X�l	�Q�ڦ,��k�hPaP+R������l�! �����I� ���y۶Iz�z�)����v�����4���1oY���)�o�P8ҷ[��E�۝m%�S��eAq��^��m���`���+k�	�^[���Q�N]�.�zngg.��-u3ۂ�K�9��B����e0��3\�.��A�����76Da��pڽ�s�ѻg"'a�p�AҀ�B+�M-��DbY�`%�s�Sz�F$+�'
��6s���lq��|Z�ƣbn�%��s�q��J�I�˦��XFU��]��[��֚���Eb,B�4ͣ[��?98��-����WXJzr��7'e���@��î;	aה��L�BE�	���<f�\�x[h���9�hU0s��k���\O�Vp�PX�l���F5^%�b�5'6�#����*]�\b �\A�b�{bc:�ѶP�]�Q���囌�f�a�T���P�����J@ec3;^��A���V���og-��8�'�m�)籑��wgdwA���-s7	�G�]��h�u��&���Q�㍝�>���װ:�Q����bs���gF�[33[��nˢ"<me,�8���U&�6�km�B�Z��4�3lr��>�AN�tmt�H >;��*��P6�Whsq�V34ŵ�+л!�g���.�նo)cKy�	I�GqZ9/����9F�3t��wc����e�6�
]Un�f05./S���]�Ì��ɹ�h-�4�=c��A+a؍����L��A۫�7t����� ����n�4v@���gV���i�%b����@G/�i�\�w8S�u�z�]��71v�X3���f�h��7�d'�vx.'�����)���.�6����!0�{J .�ak��v��g�1`@��*l��2����Ë\y8��1'i�r�kq]���h�N�z�Y���q��ϱ�����!\#�����F:�g��5�)#�����9c]�|�nf��!)� Л���kf����cf�!q�Z�K1[�';r;�{v���*j��G��ԾZ�U��Ib�����LK�n,8cF-�zWN%�ժ��U̇a){k W�=�y��u-t��ͥ�-�ƅ�y��W,7*u�.��e�r�Z�d|��ͪiX�k4��݉��;qyҦ`� ڼ���	t̶�l�p��%�BP�S��6���k��;�u�\����$������h����C{u��]��<Sp�`�h��ݸGv�	�Z��f��ۋ��״���s��g�/N��;9�ʹLY�62SB�Jƕf��h���='�"��k�)f�ۈ�=�4�z�k�v�3t������� ��n����T�qV ��ˮ��Fb1�Ҷ��\�[Br���<<��N3(�B�[c�5,���{�9�搨hQ��Ԋ�श�6imc]Q��YA,����ؚ�H��eІMú�A�8�dC)۶����P�]�� ����)FR]���aN&3du���û8�ҳ��nћ�g73`�X���i-�扬 ף��<�u`A��*A:�u.3雯8�qh����<�A�:Yq�N�7n�S-S�I�z������["�Vz@��d ��a
�ir���:{Q��w㓔x�D��df�Wj�^+����'e��[��#����e�x+�\�V2��B�tY��l3HM����-�ba3(�ug[��l�/��/\\޳�"tlz����5����2�M�4�Չ�(F��ݦ��"i��&]����d��38KHh�P�1��H5eٸ�a�qZN&c�W]8�\�%�p����{t[��!Z:�s����u���o���Ab�uƸDW�.�6��	����Qѷ���V��|��g|��2�l�T.�6��l]|�atD��9�><�ĭy�|;�a<҃v�ٺ:F�e�gD��h�㫍;;m֮M�2 �dB1�ʐEJ0å�ܻt<v����ン�C��e�����]�`D٨��!&:-p�hM���}v����^L�-ٹ�Ƨr��8��D. ��-	[t
�M[;�Ź8��&�Ւ�X:��<q�a�5]# ���s�p�bh��&4.�d�(s�<�n�5����m	����*)t]R^͆)�He�x٘��९9���q�fU�Fh�p�]����];8AW�m[�Bkڰ�����A���ph:��붹�]rv�r����g��I�Z"H	�����& J�:h���; �w�r��`;����RQO[���Әs&Ļ[��޺-t;�a�V�У3]z��Ls5��^<%�0���x���!�]��q����]e����˥a�E�������v1�ci]�|��i'>,
:�,�l�gN�Z�NR�>b���iظ������{L�`�tp`y�{u�δ�s�����T�R�0%&��F�3��*�Άy��V7��]vh�oZ�떭n�Ӧ�j�����U�����������Wʪ���j����������������#O�c���,$ݗn�A�]��̮ JХр��Xi+LFL�-�؝/�5����C��Қg$�Q,G��ƱG\T�)5��i�X��h.x�I�G���������^҅~gX�uT͏L�S��K���g��$/������VhP�Ƥel�����8�OW�w�;]|�i��b�,�H�Q�טNSA}ڢ���]��V��q��UQ�DS��V�m���Z�-T`˶��Κt�ۏ^����8�8���q�N�:t�d�T��(�L�HH�v�3D��R�}Ƃ=�m�Ɗ�l[:1��I�S���iӷo^�q�1�q�q냎8㎝:t�ٸ���\�����B����_;��f���b�5Z�ݵ]�-QK�$D]�Q�OU�4�{��Km�����)E[#Hm��vLM��h1Dtt]��+N�m�=E���h4o�:����]N��;Y���f"�����`��IZzqR���U|��=D��h���f�N�HtQ���X�!�tt�kp��v�DUTh�h�Zi���P�;:���ֈ�6�&"�G�z7�}�ESE��Sh���j4�v����Jg`�T�M�,E���3=y8��f�;����hj�wY�>x:�����fb�����N#E{���8Ƨ��;���d��Ń���N��>�<-���f���v6p�8%�^�V<,�1؎�ʁ� ��.�:�t�i���k1h�����L޻V��k:�xT ��'X���5��Н!�z��Mrf�v�:�rm�!m���� 9��mO{n%�ݴ��5�H<L��1�B�\�a��gGm�zY�6oόǄ�-4�*��j7MYѽ���p�ǳn�f�Lv��l�Қ�P�f4��3S	����Th�lc��^ .m��^�pzL���h�ô�0��q��-��".���p��ٻsǞą:X�\�@nH��rݥt�bY�l�Z�n����J�ݣ0��1�M9���Sg�Wl�ͧ�v�J��a��iz�Kr�lVcM���a9�g62\Oҫ����n<������qU�i���v�a�<�x�qdŹ^����^��n���j�����\;�g�q-����c
��c,V��r\�qv�����LcFY��v�+�)J`5���v��r'�i�gY6q�ۅ����+�n6�� L��i�4eE6"�	oK4u��m�W\&���l�	؅�;M���aiD��2FK���v2�C.UCd[X�ûsx����c�t��7:�B��X95�Si���y�@��v���GZ�ܥ��7b����r	>zp70���noɳf̧gƑ���G����\�y{>qм�*�o1�t��E޽g�����6�����NrW����w��qۢ�
�K��m
���6z�#4��h�^I�J�4а��;��<�rә�v�v��!P��eu�����[M�u�J�u͆�Z������*vZ�^��&�8���,4��I-ap)�V�k<<��|��6��Z���ܫ%Qd�4KT`B�:����X��A��e����%�ؑF��ʡ%)eB,(��Э�)m���8�DXQ�KP�A��XKר�J ���!e�XŤ�%e��k	e%�`$�y#IP��mHekaK���-��a)(�YX͙�˝���y,?Mlk3s(�Z�o�`�x�.�:1�(� >v��	>xO�Gy��^�����;����ָ��;N��0}�Keg���3�Og��*����G�&�����U�V��ַ铯�L��kɱf���n�^4i�uz�5C������1�<�����}��}��9����=�<�P�vv�Ba	�Z��^a� x�d���B������G�b�Ne�\h�C�����F�n��3�T�&I��xL)1�%��U�=�u�}�b��O�r���ｨ��c8��{�b�ƍ���}|�����jh(���R�u��7n�"Sר2�pa^ea�������4Il�}w����ss�ǰg՚"�3E�S5]��Hk}"���x[z����뇪�=���댉i^e.6�6�1o�\s]�5C�k�ڠ��P7���)
m	��3^�,���� x"��b��
�{ۛ��o� ��ee��P�ə�����i���� ��U!�Ay{�~�G�Sy1��nO�ry�{a�ǾU��yC�
���>o�e�_?��@ ��`V�k�z3g=�&n��s$�@MyV�aɄWE{��n*Z|<ڧ�A�&"g�oz����G�/6=���nr���Xy�R)j�a1��N��N׵-8Q:=��KZXJjֳJ1��r��t�&`3�΍gdJ�\��n����Y�f�7>���O��Ne����u���>�5OMSe�O�3�����Y��.�/sٓ�3w9G2|��Rg�l��HV/�χvz^�q��EI�7�>:�������9������A���{Vo��^PͬY5B���C��s���O���yլ�E�,��u���z�'��CY�0Y4�����X m�י7�X{ӷ�}��̺���n����7Y��=;eSs{�w�'�ܦ��[��cpi�%u�y��yNϩ�_HA���D5�i�=��������'�!��;>o�t�����0
����#v}��Kf��
�b� ���-狴*�s1� ����M�yO�>�v}���2٪W6}��v}a�N����)�����ݥzrvݷ=Kϡ]�	�T'� �]c�������fE��N4�Բg�i�����.�T�- K�l�i�`f��."������5�t�&i�T٪l�y��d/����N[�&q4�2o}��������_R���/C���0�f>����p.�l�7 �N�B(�O�$�ƺ����5�jr"���Nƕ�c(���n��7�VR죦�ʔ�9kz�2y�3.��ۦ1��/uQ��l����A��m���w�u�+���w�b���7�nw^���a�3��7bE����}Yl`<�� A ����_�LŷJ1β��j���ԅ3��D���&�D*Uf��o���n�Bٻ��}��5��>�-��}9��}02��M�y���32��ey���
���ٝ>��;_o�������	 ts����l�����UH��̜���7<I���v�u[6i�^m�;��������{}�}9�/�]�|���6k��=���dz*G3�h$�H��%��;2��^�I���/�v��;�&j��n��_v?�>��������g��0T�;WV�"��NU{�<��f�� =����$��z-4�Yݞj�/�7�S���f��S���V�d��%�����֕R�Y^TQT��F�Y���^����/�!�\g;M/iFk@���[�z�H�u���;�vǁq8	�޵�c�g���ۉ{gqD bh4n�����]F%�3tv���d�A�*m�h����<a�.,��'T��n�y\ٷ!XF��.��v��J�������XJk�J͡vl V�m�٬Ѵ�4��X��x�������1� ��R�C�f ݸ.�y�=4 �[f4�"M��`�љ�6)T�����|�e�2.�Y���a5��2�� �Cy����R����q��{�f��͏�����f���ΌK���_��<��y8j�[�����i}3>����_o��\�^���*����"� ���"q3\ �)Ǧ�r�f}�y���m�@(q��V��>�S���'S$��J�^f�b[u�u:l冿4Ե{w'vlz��pfW���MSg͟y���M�K|�UQ|�a���f�2�K����- ���åj�˥�r�1r��7���:�T�=YY�e�E��^+և��`�n�ع�L����LCL�<�σ3N�LA�:}�5�}q`�ԇ�����+T��
)֨u�!��_u�{�%��T:�
�'����Y����gp����8˦R����k'*���xxx>x�e�@��ܸٟl^de7�FZfzS9s�������>����j����m���W#�5�JS��|�C����>�;�t٪mx44�֩�>Y�ߍ!l[Pn�b&}���{+|�.�r�^����9��� kn�3RcU�H	����nY�l��gw2��+�y��z-�]�*�U!2�|T]�`��J���z��~|�Sd��mnW�4��:�v��K3���AsK`�V�]Gשd���7z������3Ws����7����ٽ��׬�WY�j�n��j�
�n�����G�m��}�^�����}�6N�UE`�z!��!]\O���U!�f�#��_j"�����S��/�,ї���^�,��޾��[�v��A
�֬ot]�qC+jd܁;�;)��S�P\�F��xx{�]�5����׿y��^�ϛ-�~�8���p�3�K\1g�va6��(���ɭ������d��j�]�WI��ZSƉ�rmܹ��÷��jוV��>�ߍ�Y���/�ߺ*���-<iǲ
�ĸ�A,]C�Q*�;�p���ð�ŬdH�
I�u�`�D2�ɻ��|��{��O^�yUѓw�Ϙ��{�^�J�a�2y���%�4q�9��w���F1!㛳2ڡ$�y;�U��~�9�b�b�4�<E_��Rw����.Q&�`H�pA4����<(V�쯹Km�;B?+�g�u��������ܾ
����[>r�����#�;����|��KW�h����]e^�D�m�>Ek1j�	^� ���e�b=�9��t�ޙWy�cZTH�f��u.��JGG�^��;�iΓ���fՍ�%�F��m��檞Ё���߼���w�ӽ��9��s�`DiW��U��{o*�z��X�<���$����Ynu�	�2�q�T,Հ)4���T&����&�1ӋA��4�X�Vtvs�Ǜ�R�&Pi��j��V���������/�W1�{���7���<�J�������c��G���=�^6�+�*�V3���!ˮ����Y�^��������辳��d����Ǹ_޿[�][4�כ�7�U��.�:��o(�&�I��e��yUN^c�|@ٜ�h�6s,V'���tى��vH
�&r���V�{^��3����/yo��M�Be{�̉'ϸ8u�_}�/�U��7 {(A#����ڟ����T��s~������@��x��-�[�#�k)�ﻩf�-T&V�J�HU���.�}+ٲP=z5�Y�b5�-]���^�3�:�����z�Ɍ	4���=��p�m��N̛Enj��@cs�?����^�B����@F;�b��x���n;]����l��6�!�y��7[��G���-ƀ�9V�oJ�����\��B��ˣ�B�M��p-�R����1f �fj]�k����ӷ�y*6�=l��~�ϥ�4��E����o:$F����V���of�ND�B{�bHL��A���9��~�ż,���"v��rU,�r�>��6�w���Z%�T�3籺��O9��[�*�e�>���d�8���:�c�^ƶ�p�:jC���=>���~��7�{�����v����5�ϛ5M�^oK��ϭ+]�����A���=y�/յ��ƀ��ۗs�Y���7uUM��M���c�3�z4��Mf�ؼ�YU��Ş���N�*���[c�{�-|(AY�b@�;�d�:�k:�:��s88�Q\X�k�3`v�-����O~�|���w���fn�����tϪ��h\tm�5![m�@�V�N�T����(���2�Ơ�Ȍ�J�L<�;3�\�ͳ��������;+�卬4ֳ�9&��E���w��Z�g�Y�_x�xz�2b��@Dd[�4_�[X�kT&���w;7>q^�Ӵ�)
�5��0�I�y��ș�T�M�Gf2���ʽYx�Y�̶G�f�]
�CZO��|ǟr��@d�(>R�m�ڗ�̷��*�nc>Gk�	�N5�~_�⫆�l�^�T�N�����N�+��hzK!2������̬͑W�!��W:T�����^ڔ����6����,���dUb�ɾh2�fe��x�͋�[�>z��ǳ�ub�NUN^���N� ]8m�'Aӆ��d*3w}����WL���/y�P��RhNz���~5�j�����CN_���`��w7*Zx�2�T*F<��pJ��?�k(_^R�+ᝊݛb���+2�ǜ�b\�P�8d�3z�8{�JP�g>�,ə��]j�v��+�4E���^up��s��~h�U���61�ʲ���s����ζ�����7]�u�����h��5e����j��L!�OS��fl��E��
$�{}m���{W���[�֦�1�ѓ���+)k��1��P�]�M�%��t���Sn���+���D�.+p9Ղ���핖�������ms� 2`�^�Vd{pK̳pbԤ	E]�خ�cI�`�y�n�i�wU$�$�s3�X��2��X�;�u��\�y07��b����
��7�u����7s-�Cb������;pO*p���"
�(rC��5�]���͡��!��E���v���q��/;C�]]Z(�̺�����n{�L��p���H�B�9�*΃ַ���%����F�[�4����yoS櫥X��S��Ω��'M\�u�����Z�M�	`(��oeu�SK�nXxK�xWa+׸��U�������vwm^�'H^�K�����D��f a�F{l��7C�ݎ UZ�t������9k�{��ov�>vɕu,#hz�) X�kwU�$��[�[I�c��� ��GE��$�fd3����t�f�Gvn��&�H�˻��d�wJ ��*V{*�Nν���B���f���,���SҽV�H �u�A��7jͣcXk�@ci�#b�&8�g���5�P�d'���B��Fu������|;��#S���*�ɟ]\6�?��>y������n8�N8�������������y�����Af�C��\�$V�RE˾�w���ߘ��]��&��q����z�t�s��cS�&�3�8ֵ8M����u�Y�)����n�v�����n8�N8�8��X�����m���6r���T��tn�\�Z��le�6�m���mC�΍n!���u{�G�8+.�ƪ������mK=qpn��:��Fp�N:gRj�n��m:JP��͒,�yT�g �c,X׸z�ƒ4x��x7A_�������0����u`u)��{�!�!l����g-���~\GUI��E[u��5� u�F�X[��HJ�*qo$�pqjǊ^�ַ�=u��)���;���v��h�UMqb=��6�bsce���{�kqԔ�X��,k%�[z]�f�T�R"�4���=���S]��u������gmR2A���d����%�^�x��R!� ���Q^#T4�oi�:U�۱��Aֽ:���A����}��S�{	���������L~�Ay��j��ǽ���;�;N��"��l��4j�[ �b)���֪�b��������CE:�H���Ѷ�i��kAEm�����642�2�w{7�ǧk����j�S̢�x�yzulNr��2�v[�Bj��ٜ��ٕ1��hIbA�
c5�T�=&�3mv����v�'.Ʀ��R�z��_�6Jo:��N&J � �ERj�����@�Ց���f��n�ow\S�f[�5��ݠ�Ai�
��*����N��alL�m�?~�Z�6�i�h	��.�$ޞ]�f�t`�t��	��Q�>�lA3˘�ěƩ86�v����o�Nի�ˈ���N�������I����xד���Uv��m+�,��(�RC��3u�n�����x�7�&�3�v�y��vX w�� C�s�^�=(� <s��Y�U�_ep�&r�!�K��C����#��x/-�����ˊ���|���v�>�(S��
�*�wW���>[/4}�ʡ�M��8v�C]�hoNR�{7���V+�ɱ�/jq���^ݼDw+��u��o��GSt��dg_Y�\���*�9��<n/¯緹�e�A�� >���c�s��}z��M���}���o��gZh;�-�h�U��\3}=c�qLji�ǻ��=窻�1�-)��
�P�ּ�2�z��Ar��N��~���^�
�:�Zծ�VN�/��8�� uյ�)C��ZA|���t�5H8>b��T�u����|�les8��7�{�=]�I��Xs�y�y������pWN����9\Ƙ�4���v�7����^hP�[�{S�$j�� [�{{��i�n�W���g�rL\�����7p�[�]���=D�ly7�yk�{�U����1`X�8N�Ʃ;�N1���NW}�Iy���ż����˛�L�,�#*�7��.=Ֆ���8'->���>�i3m�v5���UJ $p��"��̇??³�R�U�ʾ�lf������3&|q��즓!2�J�W&�Z͗88L�ץR(�,-4��DedJ���fԢ<���3jm]9b�q6�L���!�y���)�%MT��C!�P,K�A"��|̡��4��P�f�h�_ӷ~�q�>z��hk0��SVQ�,��ZW�:�,ѳee6ۖQ�2��n�%�,���YH�K3��u,��K2�%j�z�[������;r��勀oX�5,i	e�¨%X��;\�f�K+U%-��.��]�K�� �Rٶ�J5%�J6e�����Fے����i#ґ��Z뙶i��xS�~�~�P���+TЬ K���2���i��-���R�B(�1������p�L��,E$��I쌾]��*��Z۴�~Ә���g5i��&�@xA�A���+��U����HK����È����닏ue�sE�Z`f�9M�㝻&�8���m��=��BL���{�x��'9^�J���#5~�����k�Yx"��X�7L�+�>{C�4s�Ϥ%Tm+�	zf���|.�/�'�Ƽ(�f|B�oL�"N�ia�
~x�|z�}�{Ͼ�x����\#�t�.�\d�‴���)�ƃYWNecv�O�ֻ�Z<���^c8'z�kf]��).Tx���c�w3'�}��s5����l���@UxbS��O{M����n�����Q��Pb�1�T�Z�Gm
 .�Ժ$�Ḹ�T�����B����^T$*��+�y�����>��y�ys�GTN���_�;�����,�w�\!�Z\9˲��� �=�~�~¥���kp"���h��hu3�yxy�4��0�����Cte�&飜	Z�=�tz�w�����v����!�^�.?��4�C9K�z}�9�DȞ��ռO���;aǁ�;3� �v(u�9�SPzx�m�� �v��Bu�}�n����(̢�{E�!������ӭ8���W��w��6�.3Z19i���\��'<y�l�\�"MN��}}_�w��M�Cp���~>�|C�Ŝ_����=��37�\������5�1���[��w �Hp ����i �6�.��ܖ"���w�#���m�уw#+Vp>���݄%����6ݜ�v��R��kt>l��BGJ}���������ԙֹ������r�䰢�˹�<=9h&!�t]%�hRZq��L t� t!��T�=�s���q;U��͒�[���|YTzÅn��g��;�i7i�`A�N[�5}sv}Ji&��d������s�W���}�A`n���B�/�9ss��� k{�i9�$�(��,�����-ﰾ����W0K�-ŉ=^U	
)	p��p��&�u��n�����2�P�ǅ���{�0�	h�W��.�\�˻��Wh+�!?��m�6�b��udV���Uw���!���#i3���9Vq�r���/U��ʣ���`��A�����y��7k��z�.3�g�i	�h���wu>��::���{m��F��Bá��!���*�C�[`5H�F�ͣ�x�L@օ�=��ft�y�e���0��� �:��n����A�U8��i�B�|�d6͙N�{h���u�md��c;ֱE*�Ѻ�*�@|�<�ǋ���@0�� ���U&���Y��ռ���;a�1z�����ñxG����~A���t�]� ����Mk^�5��=X�!���5�GU���]��V[�4g=��@��gan�/�w|��@�Gkf�"X_;8y$�L��)��@qx�X� 3��Fu�|�u�9��}�j�B��1��ÂRA��#m�'<>=�/��~�����#�l�n�G����(U�e�����aw�rS���6:}�����{���%8�4��Ѩ:���\�X��n�Y��t��Q�z��F%+��]�+ct��Woz?������l�r��S��\���!'}�q�eyNr��|��T�<����}�`	�5���;����Ֆ��ϛ O{E�&�e��)�<�3�i�y�9��i! p5n؇!�P`@� �κ�9�:��f�X۬�����S}�,��'K����I��'�3ݓ�e�z�^pP���N�."�Ѱ�!�B�EHv�zCYﺁ.3<�����lh�Ӵ������ذ�vq�	Ό�[��}Wy���(1Ӑ[i��W�Oْ�`7���#��NZL\�.݃����`}9|"�:�M���Ϻ�.3|�{9��(��3N\�n�9co�\�i�p�����^y�u]YJذ=���u��$.b�)<֞������W����C����7�y	����CƩ0s�5H��w�ܿ�7�3��_F���}1Wy���A�g�6�ga�UJLR�9����n�����Qal���*���C��J���ܡ��+�3;"�v9eX�Ř�T���2�avm��^r�T(ǘ�1xW�G�|F��l�qՇk)2E�o��E��>�mKm�Q<<��ɥڈ'uש�8�=�3pu�s��v���z5�������@[����۞�:|���ẻV�t9�tpָ���Peqv�
����󪆰�]�(�-��fe���E�+h�g���p����o(��]�9��8Ɩka
�ɝhL�61^ۇB�M�3�����7:�:��)st��[�w��~�u���k�u�
�c�AhL�
ʘ�&�e͍�M�3�'���8�� �)ܖ5H8,OL`u�����}�9q�ш�eK��x�yS;�!Y����죑'�Y��'�}�l5�o��Lt��1~�R�4����w�a�ܝ�/��y�B�A �'f L��Z�B/�4��zv�Cv��5c�}�����1�E�N�*|U���Zg�ܻt���^n�f�\Am�g5H3�T�[!vn�~L��ԭ������q��U��d4�b��`�u��wsS������û�rO�\�n��ݖ�SoZ�j`A�Ô�vsv���ɰ�<9��A�O��j�{������k�nڃ��ݦ�BA��-������J�u9%��������5-�f����%-���T���F�#�-ڮz
u֪T�ModM�:(�������6;j�i����]�L�V^n¶�L6d�ǫ��X����0���l�*�<�6Q!B�����;��f��#�I����n�dc�@�V�ͳ;�\�@{S�Ć�(�A��͟�0�1k��.�Oȉz(i$,/��o �0����lm��,|�n��~2���\���ws^ˌ֌Rǎ:al`��	�ݼ.k�io��.��>��
���
���Q'ݨ�v����ϫ����mڼСq��A��Ãv��ES��T��e�J2�`��u��2�b��@ ���ǘ����5K3ַ���������s��k>������k/p�����Z ݠ�� �6��7K�Z�LY�j�=={��R�^ˌ�VǁV��f�X� ����]�Ton{Nd7�LO� ��:�������Z
��&��G�WimM	��&�*hk2�R�Ξ�����Y���a�v^eT��&) �G�W^�����|��?0!4a�ب���>�m���;�9,����J���rPs�(o����I��KIb.���Aj���N��[�r7QYy���} 9���iCs�n�*�
���U( ��"j@�F�t��8��.�|�nH+O��81l=w�aK}'��֦̾q�z���'X��:��[N�)��u�:����.��A���>��#m���a�5V�eN�ԿW��5���e� �(U/R�^�yP��~�%ϟ�N)A҉�n�&A�g=i��/{qn^�ZS{Wo���Me ��WT���QF��aM�ZY�G�h���,*�+8mlwV�9�#<�vɞW޾�^������H)��v,7ɵ�Z��j6*��WS�kɂ$�!@rK`ov��ߓ�6�B�x�!qN�`3]�5!�ҳ*��)P��� *SN,pIPn�p�A�}^����Tg4ba�]�z��}/���\ }�.r�:9��U^�79U����[;=Gۡ��6P,|{��f.���Jo�����A;�����i����]����Ϩ񆼻HO����Ps^[5P=2��u��G��ٽ'E׫/5��\;N�I�T�E�I�Ѿ
�[�3lԐ�X�鋀w�T���W�=]2��u�������v�����W��I�͚+9.��\�*D�U�����fr&ɜz���V�X�������^y�f�~ ?>���F�cm����tu�o��}��M{Zd��NU�i��ږ�R5��}����0�S��벧ۗo��(c]/1ƒA��'��^3��ɉ$hk�4�܊h��s�3ff�/ 	�Z�&�Z�Q�eZA�G�z�޾�p����/
��UH��?j�'ߘ�D��ɴ��(s�{�>����V�L!�y��g7Vwd�����'��؟|K����z�w!�)41�x���]g���WD�FsFs8,sp*�9U�9�����K�cvJ<����g�vrR_�G�]��f;~"�u\���.�Ϸ.�4</�Ɗ�t�k�XNr�Nr��Xw���u���ݑ��h9�88�R�T��ެ��_t��^���W�U /1��n�?}O���p}�_7���m���Y����Pǖ�ȣރ�n��`HXQ����Q�t��sr©c��{oB��F߷�j�{�Wُ7���w�V
�#���WV��u}dZ8c�5���o���n��"�f��=[2�9�1��Y����紨���s���q��>L���n�ǬmS�y��/P;S�es�j��+v�{��^~�����6@=�'u�Ҍb��f��ӮF�:�[K(�
66�*��f�}R�u�U�nU��\��{�h��jq�Kn���_�c��F�d�Ni¡� ���h���S���úF�����g]��tT�9��ǽ;n�˓�#7��֪��C:��َ�^PwW�����|M�㷇X�O&�Pj��h.W�ҹ�A�zU�S�5���{L��/���|�����e3��SU�^i����R#,��$�S��14aW1գ�[0��omܜ�2Q����r��=Pe�(bIs�y��3Y��٘:�u�2�m.��w<,�֍�w�q�9k�;t�Ţ�Vƺ����Ψ�F�78��N��c���ҋ�"1Y�h��(��[�+U^����`��;6����Y�ogQ�]�x�"��f+ɮ�����4v`�� �U�Y��:jj��f��ۛx��^�v�t7��e@wb�C2�fGpv�o���*鹥��;���k�o6q����iqXN +�K��]K���,��py���3xa�y����6fQ��U^�m��Doj�f�v�B�f]�&�`��T�'h=Td(���B���ŋ�O	9��+����|Vc�&��������C��xSU����n������O�y��ٖg������n�:���v
���H�B���@#�b\G1��D��.|�c�6�8^���<���YY����S��i��.�s�<�z�Y}Zf�55�қ���+�Y���ӷ�I���`��i2��/�i��Vǃ3�}Ⱦ|�T��ͮ���6���O|����W���~��?�|ƨ.ڂ�*�j=��=���U�E�f(�n���<#,�
���ۧ�O=q���q�q�v�q�_:t�󛪓tW�X=�
};�N66�X���Ѥր�S%�E2%M˺�֝:x������N8㍸�8�c�8���ӧל$�Q'����A]i�I�
)(��"���Z�kl툊(�*>������:�TM}ƒ�(�Zz5���1��;C���"���Z�4SPPM�(Ŧo�f���N�����Z�"�^���h��IQ,��3PK1_'|�^ë,w*("
��v1Au�f����@P4Wͦ"I�'��M%��o�V��kDMSu��f�"�����OQQ���tDYŵL�35E5m�	h�	��D��d�����뱈�	'�D�{�Cl����C�::��EYű�5Z��M'c�(�)nƒ��ֺ(���?�w����x4��0-�u�gm N��o��������Y�����v���h��mF�z��40.y�q�ؖ�7[�`���&�q1M��F63&c0xml��˹��\�Ad�U����#�{T�}>TK�R0�K.����*b�s�ƛ#]fc�7n�V��S9�T؞ۜ��4W�8����VK����vϮǐ�8.<�ٺ��ȶV�A�-n�cX�S[�n9!<XEj�h&�S�f�=H��"Dw��l�ْz͇ �]�qSglL]1����k��J/z�.�g��Q�t8�9�uvy;b$B�g����b]u�`�)��6
�F��Ka�ݍ����'b��\��#��*���WPa5I�j�ē��#���,>��`w��1��43z,cKj��e�bӒ�%HgD4��Wq��bA�����sMոݦ��h�3��7:��8���囖u�M��e��M
B��X%�0�ۜŎJ�:��y���CO��g�mҖY8^����Hj���c�I�]�pE���	]�n��ӬhY1�f��e��]�VA�a�d�ڜh(�P�2Ш�(��x�{��yD��ίY. ݳNncj�dj��W%� �z7��:w�������aj��j�⬨k���S�ݷۉ8����Ex�#����+��,qb�n�m.M˟R\�qq�S���)i7#��=��+���6]��c{���Å�Ԝsq��w36+K�v,��cq	hGky���,����ϩ����x�OK�:�i��)�^7^1
iC2ƥ�c-��j3Zi��ݭqx(k1R͢M!�2�\4���i�J�p���.�]l5UUUUUU8gX��=��g�Ϟ��8�S�R�4��B6�!�N��z8�Slm�@S��I�ӭ\�,�õ�v!xۉ ���
�ڳ4ݙ`T����k`J8������xm4���x�[n��k�a;:L�LVgX�OPz5��G9Rc�(4ls�)Rk1�1�%�q�d�B�h�E�[n�fF�xpu1�ϣ����zz����1m�$t���l�j�`�)�L��������J[���>�??ߧ������7l�c�5�5n-U�GK���m���b5����n��o�l���Nr���g{Ai����3������B�#sd���n�O8s4��U8p<�U@pLR�������!�3�a�];;��q�W[���Mp�Ufr�����P"���'�2����i�瘹�T��_����q�Qf�����<��m��`q��q�TPh˭�z�fW�n�5�9�1b*�^p���f�^����V3NA.�l�1j��n׽ܯ/���r��DB�[|���yE>/7
�I�s�,�3�-�G*��)�r��Ѣ�V<��%7�fV�z���
�Vg-\X>M�����T�1Mq��.}�f��.�R~�3��$��%"vq��C!p��0���oW]D���������Y|�wW�5H9`XU8qދ����e{���3��{�>�{W���m�}�Osݖ�r��;����n��)z_ �5�����_���B}ԇQggk��cr���%��F�gnn��.nmk��wW[�����VI~$�_������h �Q ����Ր��j���k�Ϻ���-��p6�8 � �8pj��3�������1�DwPr�8T=R%���?14��_������IݫWA�'�i�ncv��&�[mx��~���>��1}�'Jh�6٤��6@�y����{��2��t���q�A؅}�wBɣ��$hor=���h�UA��Zi���� U�/������r�h.w�8,e;U =T�p����u��.�x?��H ���uV�;R6]껉Xk�4ə0��J�zzX0�	!�b���v��� �z�
�;T��`/U�ﳺip�Ufp�� ��^{��!�l]�^�rZЇ:y�5IȪ@U&l���ʘ�ImWHA5Ás{�ot��M��6��ì�i���O9�6Ѿy���oF��'{��=��2��]�<��g9Z=���~���EsY�@Ʌ���r��m���fT��<���2r�(m�`��V[ ���=����C���	�";c���cm��>�ܶ�����ݖ�C�|A;�m;U *��ݵ�ĢT��2��p�� ;8 15R�{/2=��x\L����Z|���Hh���W���ɨG���\� +�<�^�S�ȫ������X�p�w���oL���|�B��m�H��xH���wg³h���>��l�.J��7&�GdY��Y�d��4!�� �FÚ��ZA֜��h5�� �/{yn�uى��-f���8���Y���ku��ux�Fe�;G��h�4s�,��k��u�2-*��q���t^^�ߵvou5|����� � ę����~��燇�<i�W&��cLM&j�1hj���L��[������VǺg��^{M4k��w(����s�ly�f�N�x�����~f�^b�Si^b�J<wV��u��{r�h�.!��	��2�+��齃}YD��β5å0F� /fns��8�#�m�K�J*~ΰ���b[u�ﲙ+yU��!�.�%w�G���>���E���b&6>yI��<������ܒY���Mv��~3�B��'>�&{:�\{�&ݜH���_OQឪ������e;y�R� �z���O��tD2D�.|a$�Pn��~��nz�GR�Z�M�F�����q�s!�ݰ�(����-���Zq��0rN=~��w?�yNTgc����x�����3GH��l�'ym�C�����ވ���:t:j6�4ji6��<�1�@;L���1>�����\ŷ�9H5RO/7�}��g<��;�#9�d�;�4C�wb�n�<��a���;<�;Ӵxd�^h+�����Ψ���L4r�UlI;Ы�B�A	���;;�g�0	-z���T����^��㧔�Fph�׈8"�����=�y^�tl�=�6�aFr��έAݠ��n�*�v7�l>��ٯ>� �;���]ٵ֢c��s�z	� ������ ��c��k��vFfl��>�X�k������S���LJ"�"D�E�2�핞�͹��w�|9xU�{���M��9;<,[�M�]f��ļ�z&�.$��U(�!4ZZŶ�M���MK�:x��y+���~8Ǎ���mE@�jWhַ3�=n��7����ۧ�̲��4Ru�\�d�b2�F��QM�9\�VT&̛�� ni�]V����)���<��m�WZ�Ѵ9z鳃� n�<�n�NK��X��eƹ�xt��X��4�L�Xu�
Sl$pn�����ҝr�C�٭�/t��2Vuv���!�_<�ZFw��i��l�]7���3C0e)` ��]�+���ir*�\�}���?��Fx����2���"s�l�,o���}����<2r�9j�/�{#sg����ĥ$!��6Ͼ�"�	�U�h�Uē����O^?���ө�У-̀~h�7l{o��\�*3�.��v�R��ɞ��	�3u����!�6��A�E���R`�ER����c�F!��m����r���}g4L.�A�����������h���{÷�}^yE�y�.�b.�LԾ�m�Iѕ�y�-\A|���64��os�N�� ��]��׊���i��'Q�U�4kR�$4�*Wb)��K�}2=w�玮S��Θ�x�z�a��Ůݻ�|����?�)�k�yS���Y�;�ϓ���
����2�Yd�G�����seT
�R��������;׿d��8n�R�"[�S��;�/rw�ǽ��y�]q�j�=3:A����E�l��e���Y�����x�>Ǯ��h�K�z���s0L�g��a̼�n4G��r���DA��}7����v�0௔e�{n�ol�%%�S˿�v�9<����'�T�1�h�6��@ 5���}N�E㳊�J�>ܯ���ʼ��->NANZ:�8�#}�`7ya�� � �S&	S�J� �S�][X��c�nN=Y���3���� ^ *����;��(U8��6�n�y��9`a�C����?�c�)wX����/'y_����]�=��W{�"��`k�/y0� �y�AqI��`W;a���}�߱���m���v���]q���i]e^r���q�^)��R������;0a�w��7t��m����حl#�!�%M��,nU�q�5�끱V���z�=&�8���i0pj�pER�r=���������?�.��ͼ�b:��;�U ��[+��%���9��]�����1�m�'�N�v�߽����);ǝ:�B{�-��&�X�0�̳��EQ(�|��״\�fYp�l-�{oO}����}Q�wNO���/33�}�!�5L��T�|�v(t�YJ�|g��K�8�"�޲y�ׯ.gv�{_��.����~:cm�6��A@(~���׿}���ʼ��� ϓ�:�8�Xَ�18��P*:�	��֯{d��5�Ͷ��ȱ�s�T�=f3=�ѕ�*}�޾�@G5bJ�}]u�۩��N�F۳��*��5[��P����B޽�>e����s1\guǽs<38y����6�5R"�^�{���Ā���_���������F�w��"f�Y��X�Y�.�<=V̘��d-T�U5���zZBo�.[Ƭ��d9˱��{�o����M�d�j�3�!��q{�����&{VB3�U��Ig{^0��i-�G�K��;��N�O��G�Y~��ϕ�*}�ń��x��2
����F�5�l��('��%BA;�������g���;9�PЁ5K.c���%����ܟ;v��\�� y�;�m�D}�,��PXs�z0�v%�������u�_;F �v��k���r��ɿ��ﳸ��ɼ嫘�H)��NE_=������~Xg�G>���u���&�fm(5�z���9�Q�yz#���xbFᣵ���YGO:a���g2�g7�9�s��S�=%lh9AP����Lv�+M���Ah~�g���Q=�O��PH;� �A�A�"�ñ�L/��U�������Ê�1Q���\2�٭���^8�a��aE�gnљ�
_���(������Y�?&�-��c�Mp4�0,]�Kv��a�M	��k*�R��?�~�H�gߏ2��瘠n��v=F�Z������䡸!����}�8���d"s,�u�QdNr��U;�R���9��Ǻ��gH�����vq�΍���j���Sq�8�FS�U$��J�
]��0�X��p,w ��j�<�B��Ɣ35�?�6q���v�|2g١�|�pA�q�E��c����h�����3[��V1��g�]�$�����z�FwZ����%y_CLʢ�2r{���~Q�5=��d�b.�݊�3U/�MT�����󝮎`"i�����F�w+W�5�� !���A�vsT��J��������/�o�S57(����ׁ>����+�_���O�e�eqQ�h�=3shK3�ű����ʾ�v��m�<�_T�����M4У�Qf�UMj^��Q���بSlm{����oV�S��Gh��`q��p�8��E�ao\�u�s=���ns:.�u����ݗ�3s�������!��R��L.1C��� �!3/f�qj���D�8�㋢m��ǜpk���ڭ�X+��)�[¼�Ak�ӭ�;;J�R�ͱ�b��͛3pBmc�i�ٲכ^ދp�j�Gk��q��|����?G�-s��ͮ�҆�%�C�,k��^��s��$(��c8� �d� �� U �ôa�db�}�3����q2�H�ܤ�#��a�-�%>���ē��0Ҿ����]W�l>��;���*�wZ����<�ۙJA�v�L'���{gN��6�%�;�!�t�lzm�������
�R��}"�,�o�
חu�3��.^b�{�Z���嫀 � )' ��q��;'{V[I�ֈY��y�eo*�,�m����0�:y�hG��1o>���sz�8 ��z���LR~�f�M��ǉ]�-v�=ӏ1�5HÖʐ��F��O�9���֪���g:�|��j�3�Y;�,�EWn3~䧾��^Q��
��\�$@�F�p��4�P� �3q��X0�YA �I]��Wޯ�yO
�_����T�3<� bg�=��=��^\�r�����2�?bw�B;�!�(n�{����9$h��>��+&�p�B�"z\���qs���w��&Q8f=�^�F|^�&����hyz����0���,g��1�\��aL�rP�q4(I�S�~<c��J�cm�P�P$A@�j�g������S���~�5}���&}�޾`� j�9O>���{���vLj����A�qLa���M,���+���y
^7�g���j��g0�"؟ �t�T����d*�8u��=+p����0 ���Z��;L���lD&��{ӝ�����-\Ac^NXEj�����L島,��xw�|<D���H�	o�$_�`����=�k����������#�U!�"�X8��N&݊���ޓ���%��]h~�����B�X�����2�h�KoX���Z�pGp/�BQ��d��c<� A�p<�O�E }hɺ�9���5]G3��q��9�ٱ]M�Hq��u	]��9�n�11��3�Gn��)�m���sc�s�ڼ����2�d)(b[��v�!\�X�걆�u�
��g ��vj�r��S��  ��<��s���}*�`#ll��9�]r�*t�pV�{����x�V�U�n��J��&��9A������P|�Br�a3X����=�P�5�8±��a�����T�VW\�Kۺy�smWIꀬ��]k�����X�ˬ��ݛ�Wq̦YK�
̲+t�����#X���2v�V����7���w3��$\�,^��ф �S�w;Σw�R�<:����N�B�oi���un�Kέ�5����x�8��ҞW`}���Uͬ���0/^,�;�m�w��[c�� ƴXհ��2U��g�S��n�02����)�I�W�x��;�%�Sל��j��oK�o/��G0U�7W�hl��Њc��+
��ņ��u�p��U�˥.Iq���N�9wPN��-�;���htJ�c���/j@wL�J�kt�չ�@�e^��&�9l��8��ݶ#�*�[ʵ;MnP�s�.�W��%>\�n�]�k{�ۋ�Ǘ�V��|n��;�n��g\o���E�.cޮ�6��̺�U�-C���].zx���uӗa㚧I�d:uʸs:ٽ�L�=�/�w+�GҖ���'(���U��l�?u�����i���1-� ��j�e^�:��vw�����X��gNc=՝B��9���']�{��颶�^|`���ivii�O7;��x�*��1T�@�S ]��P$Iy�����I��P�\Gp*˽�w�e�ҷ퍌>-�ԥ�|����5��4l���X�6P�z���W��
��4KQ��𨐢 �%Q%��� ��?-DPU$E��P餮�1,�y�9�Ϗ_�����q�q�v�4㎟_:}x;� J��Q�)�J)�� �
+lgQ4��������|z���ӎ8㎜q�|q�q�O�����?�!��
��8��+������<��b��X��M.�j�ђt:5�U�i����>�KEWZ
��H���MR����35K�%N��D}ؖ����aפ����"Z=;�CEW^x������'X�u�-�M7���ƌX���cUT�GwLHT�Q�d��:��b�b�"Kb�&�����2cQE�4�ݱST�E�7m�?'��=�z����mf/�����m����뵉� ;w��Q�^Ɉ��F��Q)�?/�Q,��b6�M��H�系�S��_w2y�3�}���BZvB��*�8N�)!���H]1O��ɝ���8 ���:����s��t�Ά>�y3H^#���h�8a<�	̲�䄴�i�m���M����Ve�X��.w��<��/4�Gl�q�9�y�W���r��#m��
�9�R��r&w�k�W���@��W���f1�-�Ʊ�'<�b��0E�n�|��~�,����An��R�B��;{�{ ����>�g4�T'V
��! ���`����&��+�D���ܛ�{���_�'�=��T���j�mW=L�I��t�o��,�+w,\_�� ���w"2��c��
(I-�̟-�9����E����8���+���̛�Z���L�m�X�1�L��8"�8,Le匸�$ō�4���H8�7샛ձ�}>�i�8�z�0���Q�?��gN�g=����Nwe��g*�X��F���N
�/�m��'���];~г�_���umN[�\�vS}�UoL��k��|}i�6�M�����N?�g-��m�5�֠��d'{a�"�qU�=G��C,,�3}<;��\�w�_
j��3p�p�� ��T�"t��6s�\��9|���4B)1Aǡy%V�k��^�����·ڦe�˚�d�J��s!X�k~��xJ��GS�2�K���;8�I����u�9�Y�W Xy�0�ƌ7w	�]�d�֝Q�Wʹ��l������9~Ǭ%Xv3H9L@W�Fم�ձ�}>�i�8�&j�<EP�]rt�tO<���n ݠ�ZpA�tŪ�5R�����h��ឺ5s5�r�K�b����n��S�jg`jb���s��t��K����ؐ�L�f�vx����nwZS�5��[pF�#t���;��B���3��y��;|m��"I�Ps��=�5R�2�!����gelvO��k�wb��AȖ��8"i3�;(�ޣ��x��{�S�1��bmo�����QiF˘����G����,-O ������I>��R���o#�: PQ$��徳<����>R[6�Z�/;>��d�"�ङ�~���~������y�<(!H���߯�x��Ƈ�7S�kSOk�D��냒�#+��cҎ�r��i��]8����KCSU!f/8�׀�,�#,I/i�u����1l��V�h&��1�g@t�����<vs�Vx��4�Y��.��!l�;u�-1�1c*�RKtЪG�Z�I��9���V���=�I9�]��+�ke3����a�ԅ��hR�˳ 
��^ͱ���6�%���>�[����e���P�@��n�;��nӴf���u��9|�]5�#�B�1o���r�:@YE��l�����!;�z�����]��,{F�#ɞ��G��F�o�Q�ɬի��(r�b�n���~���u^�-����O� �ר=2��d4�=BEOp߹�a�~�οӗpǙ�|_S�E��h���ݱ�-�2H`��Yy��`��� �9�@8 �T�4oMa�u�M�
Pv<m�5Q𺜾��!G]�bŁ�v���E�'9eÜ��9'O�$��}a�n�}f�;۝:��Mf��~,	�NDbg>j����Y>��i�ƻ�
pU^��>T�-�o᥮���u[�d5�����ܱ.�7���0�v�r�q�M�dSYq:s}�k��}�h�^2�h�^]mF���"�<;�r�����K�k��	���ޠ{�Aˡ����m�o��nQFs۸���kNrg��+��⽭��f�V��g9�w$�-b���>k��'D<��D
� U���v�%U3	([�m�M� ��T ʃV�a�x�-�̔��ly��M�xz�h���,��L��%i���c�Ӥ�w����	6�M�$��H���[� ���v���Q�޹�ХP�p ���	l�'����>��4�|k����>U~=S*"��{����j��+�.y̛�n}\��_�9�NA� ���� 6�4ԏ�5��9Eʪ��v��r�
��ݗ�{���i�7γs5�G�z�Z�,Se�O�������o<9�aܽi��m�8�g+�f'S,�hcv�9�)�O�Pî�=���:*c���W+�k�,.�p�A�pz������V��pS�V�k�m�e�i��0P�����j��G��>zh3��T���T��:�7gzy���Z�����+]���V�c{�4tO}��D��_'*��RYƏx��/b�L胔���v���]�[ы����o�Bg����9e���-�5��ֵy��5��` ����1��,.�K�(�*��ڐ����<�WO������T*�Q]y6�jj���@�Â�S�+K^A�B��/�Ok��K� ε�:��{;�/��	�.���n6~>��h���mEVDIdP��~�3��]��������>�,�R!��-�����[B�>����ș��i�vw�����r�1���B��囉ݶ��k�NA �X�F�(�1L L�m���r�h��W/=�̜�8�h�3��ٽ}>�i�p9�9�*��4|*�E��zD;�/A�� �b�2�����p'���	0.چ�]t��pg��궰�������'��BQ2]-kS�a�V�&7k�v���/�����W0R��������σTjI���ߨ�$9�/�Ё�*��v���d{��xvv �N��vx��~�n�����jn5���"�ٮ�Nܩ�w�`9�ȪNA�U���n�p�B��W�����'C\�[���c"���5�	�B�@mC%6f;zAf*��l���Ƽ[�+��%N9�@��XT��ޭ�3�P�]��\W1gmm�o]�S��-��wP�^B%�u=�i^}�9��ՠg"�s�;Tn���i^YU�}�sQH�Y�p����m!���h�"H��V����-�ݢ�s�����|j3Ü���m{s�3A�k���.]�o�������ɬ嫈&��pA�vpj�H�v�~療m��:����O��-��i���8�������C��m]xɒ(�3��|?Ie�|A�#)�9�Aϛ�8�q\j�Ϸ��2.}z�X���m���;��/PUN����&�-v���J���y ���;�70̼!��n˸>b� M����a�������ї�~&yV�SE9�3�fQ[�|:���+� `fHv����hB�q�w=��xPr꽻���k9j���^]���B����պ]
�A~�5���W�P�A
�yCc/hO����w^�_�׭5�8 � �EE*��#&���ߒ���@
�	��"���Qz�7e��
ӵϪ�Lʎ]��|&1m�fvOL`�A؊�;����#�Y�r���EطFL�(���Ώ>]eD����3^����;���H ����n���s�;�l�a�U}`��X���to�acv�y��>4�cM`�ĵEL�������:^{��d�oI��
�~�~�u�o{{��&oX�=�-����MXy�(��ue�aV+IZ�����c9�,u6����x#���nz���dy�]�җ6�<����]9��.��&��,��^66�a\�h�1n��vj]-T�RL�fWtZ�e;bp<�kU�����G7=6�����%��l[]-��7
���������x�dւ�2��u��:؀S`���r�\v�݊Lc��g���gy�,�i���bN�3:����%W�Y�W�����xz/'Phc��D��T�CΜ��MMG��wE���� ��.�ǰ��n��^L���H�p�L8
�<P����ڇs��dQ�]	�ۧ�$>T$5_G8��p]��OݖfTX��|{�0��2`��pE��C�AN�Z�0��'��秽�}�+�ڔ4��� �束ޝ}���w��ɬ嫘�y9�o"�:h�֒7��༎���J�]���	&5H&��@�9[��6�7��p�f���%���
p���5�R�Q��~^#�����٦��c���H"]�
gq؍�D5��]D�n5��Q�+�s�׸~'޽-��� v�9�N�4��{xfTh��|{���Y���{hE�!��2^X�=�9`Eۇ�fC�cv� i��~�ʘ�/�w)kL��ɟ�ڙ�m����[�ȷ���\�t�τ�����ގ������{��s/�7�u�ڔ~���ZmR6�M�����������m�y���~y�}�J�&���,	�; �2��O����мw��<�gńw'#,t�8j�<-4\>� �F>�G?jA:�Wb��w�:<����zq�=BEHT�IzC�ˁ �I3�&&_mP}yw�K��.��@rN'18��mƩ1ë��祉y�Sl��;�MM�d�W�X��8�;��!w�7hn���>��x\�۳��缏vwJUyU|���\C�S��j�;�^#е�Z05Ɨ�P
u�M�����ӷ4��Fn[�5%��i\���-4+��&ւ���@�\�H5H9U8�9�2���=�>���+ެ.v*��#<��g(l�-��]�r���w��G��X1��� 3׏c%F��Ǹ�	�s-����Rê�lz������z��|��T��T�;U;vv�.
��䌠��[�d�Ò���Q��Ro]=�Ee�Ga'�͛��������7R��`i��r�J�!���oU>�P2����~(~;|i�d6�M�2F�0 ���~����%W�Wϫ����FS����Eq �pU��]����V'��a ���mbU@��;�v�z�3�>���v<�
�$����9�ϳ~t;�}߶ٗ!/�g�	;aWm�vj�F�3n[D/�o?x�׏Q}�3���L�SE �� U<1ڰ��+�>�wwI�=�s .��.q�Ps=��m��PKA]P��b֭vQ�~��~�K�b���f�MT�P��?F�sz��ʫ����nӧў�>n.b�vօ؃9�N)��2�'{E���y2��d}�ߔ`M����;�=��{�s�3�8'���A��B
cTw��d��m�v}e��A�NA�xb �'��g,��d{��s���T^��B�I��\�n<.�8�BӸ����%�=�Fz�m���}��N!
�O��7ۛԔ�U_&}~ ��� ��Y�7��aJ�TQ��#�"_⑾Z�_sj��YB����U�KM�s[Wu���4��:����PYG%v	W0���˼֗�:6ƵJc;b������O��s��<�(
�X��fX}�?���NW�Nr���R�UO�b}n<~߆�{j�&�+�L�ƭ��p*���n������}�4��Ԗ�}o��'��̷J���M�z�=����\�c��+����`�M��C��^y���,j��W�T�{ӯ3|�z�/��q�+x�Ӻ׼�C��)c�b�ER�0�]�7i�=~^&�+|���*�k��=3�������*�5s��rA�vpj���F{�]���>\	��xs��1f!�3���(وwv���G:�{*��&�+�L�~b�7��<�]�;H�vv5IȮy��S㶩E2	��lXCd����y;E����o�o^S��S�u�,��.Oy���ߐu|,f�Eϙ�B�!v� @� �A�p�U���q[_�ڽ���y<��r�cPn5�<�6���'j�`B������8ÿI����[�:{���T�v�x!�4$��[5p��ީW/�Il��\�J�T���+Es�. yVJD�.�NV�&��0H[u�{�U��U�-g��ǸK6\����%J��o�gd5h�ĝ�9#��C��rм͊�w�9�fC�;F�C�#�5���{n��ʱVȷ�\�k�Z|�έ�Y��K)����B�]]uJ�����C��F�9��݈ ��V�������.�lz.j�q��k2����	-=�4��lŢT˃N��`�������b���N�B��[�<�{SSR�^��o$�������(�_4n�
�;G)+F�]m���[�b���;�ӻL@�y{6A�ܼ�{h�`�4�c�8�b�6��n��hY�(,�ٻg�r�������\�麻
c]�Mm��ͯ�{�:��9g[�$ُpr �6o3���0{��Õ���j8.�����sc���m�:]��<���Nl�JM���Ù��ƻ���(�ݻ#�=u���^�nj}�;)m���ή��FOp���ܹ灻�M_kǱjU��ݩ{Y"3D��u����@�����wލ9�����^k�NCt�My�N<�,k��c��zadZ�U��@�8�O`� �6j��	5#1n<�W:k�<	[�(j�Ziqд��������N�&��:��#;���v��0>N�WF OT���V+"��U�0B�7�j��ˀ�n�U�����b�3��8j��XRKg�i��T0=b���_�l�:�u�u��W�G�#e�B�A/]�X-�Dѡ١��b崍2U�>7hѡ8�����-�!�����1f&Жz���s	�3_(S�o�\����v�̮ґ��]b a��*�[t	�R�Xv��[+��il��8��u.բ��5�ocP|�/M��2ٝ3x�g��7�3��ܲ���j)�]w�f��*Zb)��N�oZ��"�a��>s��Ǐ]�}}m�q�N8�>8�8�O��>��*�5(�ƹcQd�}��l���]�(M�ޓ��>t��㷯����8��8�q��t���ל�#������|����4D�=���u�$h4�M��Q���2{��t��mM�i����PDmM	5�i5����š�s���M? �E?'��(
*�c'�݂�~o�^���:[ƥ!ڂ>���IG-~�!�����L�hSUF�ړ�.�-�'���h7����	�-d��8�GA�b��AT�L~ڧ��z34|�(�֚4~�_#�-�����񦵍�����2�p-tt]�ǉ�h��`K��5�eѓܧ��y�8Q��]���t�k�`�g��c�Lu�ѬC)����،u�ढ�s8��x��lӬc����Iie�F\Ѻ��Eq+�*R=r���d���m�0�ó �3-��/6[4�k����� ې剷P�.�c�ӱY�s�`�-��Ybv%S)�uβG$��\n�N�mve�2y9���|�~&-��'V;�ݬ	r�ch\a7hua�.@�q6���Ҵ�[c6Ȓ��B0����"�<T��]^���n�ز:�Ħ5Z9�\:2J�AMNv�����Tb�n7^ݠ|��+Q�t�T��E5*�.⭄IH;��q�#oV�6�w񤀋��V���ճ\)�7a�]��lR��� �;��e��#m���S�1<�N�&7V�ˍ�k�`��/���l��{ad��v�ܜ����v�`��j�0.%�0��R;���d:i�g�v�m�F��Z�&}tt���ۜ\=���&3������:����ĻB�.��ځ,p(���.�k�Vxv��9]j�8��a,,e:Ʋ�/\��cfq+�v{&�n�]t�a6���r*�M.�B6W5� M#/Z=�!E�Y����Z�](WP�m1�{1Y�l��'[�@޽%�1�ݭH����[pq�bz�C3�,<�u��j�'X��h̛���"݉�Nv�m�	X��1Ռ�Z:ż�K)�FP0�V%�����K��%�����h���z6r�tn��p5���S��p��%�u�a�ݞK�id [Iq.�y�s@t�c8�9,�G\b�Q.�� ��qp)�ѹ��v5���Pu�����������ʎ��N���O\��]uq�AN.g�
ʪ���@���Є#m����E%��߾�ߺ�c{ֱ������xΗ�c���Fꬹ��2����H�Й�pܗ�3��#d��ZC fJ�����U�0Ж;0�$uWg<sM{o=h�#���6Ţ!���ǊB�5�D0�a�9�ʕ�]K�{�(N�X!޷.�=���	 ��n�en�R�v5;��B$�s�ֻ9	]�f�?���^~�p��^"�W�]%�紈��;��ے::\�Z�W��f��a'�QgZ(��Y;�.�چ0�����z�i�<��|:Ν_�(}![ʩxW�U�$(P�!L�z��gy�K݁�Xɔ�	�/n<�|�:�/D�p0�t�I`n���j���E�#�F����p�Y ���;^�偺p*�y����4'G��[�w'��U���&�3�8K�C ����H$�Z��}�e^�pɄ�H�v�Rũ!Q�sF{{j�&ޫ�L��M8�5t�~����RM��w�6O��'�y����`U-w�׺��o	�=��z<��u��O�|��c�3=ӵR ��N/�~��r���g����y,����{�͆W����\mOv�E�y.ۊ�F6kF:�uИ��������~��؊�v"��?��[����}s�}��쮂��EV�L�� �Rvz�R*��]��DQ�}uc��8(Ó��|z><����"�5Y�*�(�?Q�mh��T���#Gj<-���V��]���任��? �׍6$m��$@��Y!�1ެ�~}E�b��<q��?m_e[�sL�|b��x�}܁fA�F���R\/f����&�5R�ƍR��%�5I�V����s2�/��q�-t�
��2�P�*���ݏ\H���A)�<���u,G�ݟ�|��ov�_���WH��'�z���N`��r����
��!RA�c ��9�B�=o�5��na��ÏI����پɷ����V��n���A���s.�c�ۇ��T�:p� 3���{�B?���(�M�1��Gg�[�&հ�9���%9t�F�hk� �����Rr	�OuO��؇�̧��>\Xx)V1֜��}�:-�^�T�՗��~�?<��J4�;ñ�ڹ�?H�W�����n�^�r>�N_;F��r2m;5Rp�a)͊�*�l*�zi�B�>�$>�ɕ��3}##��3�~��Cӏ*�e.�L�\�����,�����G��>c=�?�<����)8�w���y�y��'��ƛH0�m6*E�2�F2�o:g���پ�9����'r��[��:���x�{ZH�a/}�	�k�xRA�;;��5I�&�ߺV�ofK��	�n9�����L�X����5���*U�
ʤ>��i�bT�H��%[��x����@���K�v�_�/�W2�����Юӂ��v�2��ll�8�8Q�G�	 \�S���:�n��rt���e˔Ҏ.����)4�Ԧ�<��A1�A�5�`�� �a�N�o�n�l�e[�sL�c��E���3sE�v˶9m���{O�;Q�=�m��}�8rr=I���vN�o^K�����d�C��Ì�b�v�{:ז�LV�N�F���չ�-����4�9�n�i�Ȭ��1��^U�����jn5�� m�[B�N�y�v���pD��T3{�����E�y7N<��ERo�f�l�a����6��=7�P�pȞeяp��u(�n;�._��H䣲�%+4ϯMʽͻ��-Z�����g�J��y[����[�2�g�_�cH��~>=hK�m6D��H@�D�D yv~C�tF~{C���^����Mv���w<i�78������t��t�rOz7�%��{ˈ�Kt���RA�vf���nS�]�Ew���%#�3WK��m!B��f0��c��*�9�=�����,8�A�́]��k�-u�V��񹜽�Rܥ�Y9H[��8�����M憷�Pzט��,@A���Z-��:����u�{89�A� e;��Fl���N���ޫ�!+�^Qa�l�M�+>�e{)����vY�)��H,��A�vsT��<��W����q?P��_^LEp���9��w���;�.������A�c�=�Z�P��"�݈�p�=yWv��������k�3�̨��Z���s<�VB�+}���1��r�!9��K/�<u�x�+#�'����M�N����i��p�(�q��l9�|O��OJ%��@wE���L�s9]37��b�f<%��N�����y�����w���xjw���W80�٭\�m����d�PuOŗ>

�5UDR P���!���`�ad[�/����9�b�y�<��@BU0��l�u�g������JݵCU�C{h^�K�Rī���E&X:�*�g��;�JE"n�Y0�d�ZT���.��݉��챆��uz��,�6�I�*�w��+t����O{��8���������QcG����P�u]�<L��c��j5�
��v�ǍR�q�c"���_�hk�Å��l��z�������G�v������յՖ�\�$�rqs�X��C(�Q�y~  ��NEj�x�;F͕�=����x���[zE�<$�B�n8s���j�sw:��A�zjk�{�݌�D1��2=u��w4Wx��_F������:ݜ�*���oЬ�s�E���
ŭ���8S����)Ѓ4�gb�RaL<ϪG=;���ɫ�o潢y�.��ފc��~���=�k���:�k�M���pU(ٲ��f�/@�&�A؋���1æ���� �s��Zvv�A�5NU�Ü�|��8�k@�vvڼ�x���73�ѫ��'���,�'b�o�3�� �Oz�?_�wǈ��U�W��h��Da��bͣF�s�uKb$�6-�kY���8��K'����&e6��ERg�[@��@�9�6{&�e�ַ��1�vt�t�F�ըHm�;��j�3���C^NG�*�rFTƓ��ط��va�B��r�.T<�Ƚ�g8>}��}�y���ӧty(�y}3�*��|��O>�'��8��$���d �����&��i%�όF�����֋{k��|~�_f{/Dyq�y8��p�/����ɬv!��pA�@=ۇ�*���!��>^��>�x���73����j�g�v�7jH ݦ�^ ��A���� 5�m�����1�R�#�s���l�˺���� �W�wUz�ޏ?G	4���|'�%xP��(P�^�	o���|����|sd��cߴD�-���
��	/
"�����s<�*����������q�4���Ҋ�t�6�M�5vE����(X޼gbAN5 GQ$����j�]�6�Wx��^��~6�"�Q���A�vsv���nӑv�A�A�^nlq��y���kPrU8x�y��{f�e�4?y��R"������,��gg�"��_9x��SB����'+¤2՝��ب�_���C�F��v�9��SK��_m*@7q�E��.�.\�7 ̾)T<:�-`\��Ժg
�f��>]��u��Lσѹ
�>��-��L�s�y%�X�����3��ˤ�{2��"W���1�Br�/��K�^�j  �F]*|�u��r��#�T�؀Ηĝ�v2�]�=;��+�oӗϩ�ח��ɇ9v������Z[��;A�&�@U!B��#y�u�Qj�>?���s�f�1t��d+ˮgt8�B������^�A�w�'�R�q��3Z�>O��G�354u�!6;M�[6@ql�(�h�j���?|�~�[�����̾�;C&�^�񷍳�{}�q�)7 ��|o6ZWN/������"E;�/,�*�'9O�W��{9�m��[b#Ӽ������9|���y��i�b�S����������8���#��L͞Y�I.3�$nݪ��� �8�lnDB�5�Ӟ��W�<����Z�
�ES�j��j��G#(V��QԊ���Nr�xX�U?�lڌ��{}�q�)���G�bB�LDz2�MF��J�c�۫������7�rƑM��,��(h���Jջ�4{�ۄ^w���z�þ��̮MC7\���F���y��2�7��r�0rۇ"�õRکÂ*��Y��م�a���	��V��ݺ+�kӗϫ�.��r���^
�T�b<���ǻU���&2��=��!C����8�:	��v�	2e5е�A8J�4��M��,�=�;�]������v鋁�;o6'�ݑo�<1�G3����L(.�����t,Fy�b/|�S�1���T�%jݲ"Mb6� [|�����I��fG�D�1@� ����v�y�ؙ۠�<)�E�ZK;Ti�e�f�C��������Mfwx�8�9������kәϫ�,oʯ���?	�
Cr�ʔ-x���-����6���B���A�-T���s�b{�������	�qP�$�D[�� }a����n���k���Yw��tߧznde���V^�1�޽%c����̏pyM�)y�Eˇ���j�lZc��E�{������=�ݡ�t��*b�>C�C_u!${A���ڹ٩.&�#ώ����}{�<�Yd�ϫ1W�UC���U�h"k��U�s�yI*
�dJK�3�<�V�e�k���o(��s��O�?���x���&���^�<�_g��GC5tb0��յ���@����ǰ��Ŗ���]M]��`�^(v��Ee���$��V����h�3\u8����(�;eN�ݫ�L��M�\Z��(��aeVB�Xi�uqT,b	i�@뜝d2i|��C���ΰ�7\q]�^6	v�e�g������l�	Q�������}����r\��)�p�̤�(��T��M��S)MXUnr�R_�Ya��d����c�r*�=S����<>nh��^��}M]�j(�*�x}�gm;A�V�]�.ж!6\�Y�EZ��h� F�����nnlu{7=o�:����6���p�EQ>���O�����@��x��A��w\q�9����P����;>y�Ib�V�i�ř9�:ɋpYH�t��YRA�H<73��q���<�.9�!!�ج�F�ݪ�8�_[����kәϫ�C�r
9\f��2�.��&�8��	�m�j;��p�AݕR�^�=O�pD��>_��u{{=o�<������S��B�v�{�s��D�|��\���~v��?F�S�z��T+l�$ t:��6��[�tC(�Q�m�W Z|�����Ʃ8-T�<{���;�]����yq��޼��xN��^�d�n�ŏ����y��E�K�)�h��r�yк���S�yOwX��xw,5n�u�vC�z,%�/��}Ra
=��p4�J�Υa�Z�'D��wS�h��Hz�!m��@�	,I%��-�������{>����G�������;FہT���Qv�9�>�4��Aĺ�AcPrS�RU!#cjj�v6zk۞�|��w�� �hT��P�~}�L��,������K�t��K�ݫ�A����.�~�|��O��Ac���<��'6Z��c�y ��q�..��A�mhg�@]��;��6�SA���=5���E�ϫ3�W7��6ݜ�' �Q$���=	�=���ĢJ����,B �p�,�vgp�p�[Q���F�t&0�hf��O���&�'�&�v)���p��Ź�5��]�d�;�8�oE�%MY�<օRf��zbK��Rq����=n��F�xk�ݯb/T?��9�wڻ'=~༛�� ݸsT���3�up�3v�:aÇgg�� �8pES���v��[��{mU��_���귘{Q�!��R�@�t@Xtc�)ZL;|Mw���烩��|����qF8���r^���6��X��k��Su�Cѐ�@�C�C�r_f�F<�ݜ.�E%�5���B�Q�/�)�,=v0�y��Y�	%U�uNS����;؎�+J�X�F� m��t�}9�o�`��f!�Z<v�o,���ɇ*��=F�Pe�qps�R��9����o4�:��F>��]e��͡�P>�;tF� +��-��WZ�`;q�_.�KCU��۷�U<��-�����5��k�\�)@���E�w'd��ڡݣr©Z�ݬM� �scƩ�S��:4�^�����7P�T뗩ޗ�-E/v�o��o,���Β����Ry����2��!���b+:��E�ܐ�2���J��.�V9/
�O>���6�����۫·�T�0�|.�uv��ћ��WN�]ٛ՛ʉ�m�PNݫ��:�nÖao�%����'7z�h�ubw�,��ִq([�� ��w��7Ed��}�Lާ��[A-w�9��E���W2��q�DK���/��/]d���a"��9ݚ��v�y��T�0�T%e����M���:k/��`�ٙ+�֛�����y�c��6����ŕ��fe�-��eZ�릐�.��(�/���O���Eߺ��~��X���p����>lV�z#���DS�����,)���x� O�)�݃DEKQ'��9�����}}m�q�q�8�6�N�]>��yS\�#ؒ�B�j1 h���F�����E���Ο�z����N8�8�q�q�:t��뽲l���!R�J�$�Y��M���� U|�"ѿm5��k��R�������W�>^�_�O�g߷���������.�'`��7c@W_#�4S�;���#I���+�(��ju����*�Ѡ�����/��������S�_�x�G�0RbB&��m�-Q�֚
5lRGͭ?}����tx���M��

��h=h7d�����$�:
i���������_gv}n�˫���'�>�X��J��4��F	�?ܞy�tQB/7r�Oٴ^�z�7Z
�[S8v�9��Ro j�b*��ރY��k����|��
1�B���7����k2y��3�P]]h���̭�k
l(ߔٝ�g���

�R/!!���=U[Dեc�uo�.��g�/,n@����u��1���݅:~O�	��_Ii�7r[�.1�A	K��+�ɺ��9�Uخ:گv�h�'�Qs�g�e�;۶=�#���ٴj8z�8���j��=��F1k��=Y�Eڪ��<=�P����r0l+�8����lv�rV�v�a���lub̞g~pA�CD� ��v��
c�7��F�����^b�@��v ���x�Ry��;�.�5��YC��rs��ˈ') �v�T�A��HCDy��{k�o"��=�_��Rg��x���5=Y���q�"tW�wqj5�W����2}�9.���$76�N�A��}[Iv�s6��m�6��!ϳ��oC<ALP]���N7j������4�4�YA$Bm�tF�6�J��i�I�,j�q� ��8�	��D���w �g�{f�f�,�k;�8,j�r�T�H��H�^���}w��^�t��P�=O�O�k�Zj�n��״�Z�.W��K�� �$MEWa�:yp ����n5S� ��T����6��{Wd���2��|��~i�1���s�m!��p�l�\�	i���V0ow�r48�n�Es�l�ŷ�k�}Y���ܘ��؍�v��(�C��Y�O�҆-�AȪA�Rꜱ�9x`fr��W��4�6��=����"�"����;=��PF�J��A����miu;=�4��j��A��W�}��s��ˈ�Ae�cX���q�H��A�"i��4� �(�A؃���Q������g˪�6�w��3�|���r��e���@U)��=B�������k�,GfWR�N��3nfAz"���p���C[�`:27����vn����a&(��k('�r�T�`���XX Ô$���ӎƬXAw�~��{�p�S�X*Ro{����x�����Y�YX���&d�i��/G��Ƹ��ܜkֺ���k,f�;fS;CV�P�;dM��41��ܑ�i��6b���A�f4n�J<)�[G6��C�7o=�1�Mf���RZ�������hU�8���na2k��$A�".�^���3F4�m��a�VL/F�k4m6�1��̬��������m���bif44"g4\$6�#��#�H�p�Q�)�V����ۇ5H9�È�U��4�:�3=�]��:�Oϗ�m;T��j��MRr�f��z����j-hz�9��W�;d���(�Ú�;=�g�#�d3]�$v�Ȫp����q��OB���)��]��������&��F�g7i��.+.]�r�"�0,<L�DEt��4������1qT���ʯ;�G���3���R���\����ǼLX�3S^�!�R��J���o��V����Ѧ�y���#��N{=�yp��A��A���S��Կ�R�Jw���M�l�X�-�Ȇ�ʇPsp�XֻII�Q��>�����,�}�������c���s�E��ͣ]'ՙş_�~pQ	|����z��5�_�?a�+��U<+I����}ڿw|�bI�%ȵVHյ_�s�goH�e���E��˽�{� r��aՎ�7N�+��Ͻ��ԃ6S(��Y��q��x�`����C������6Nw#��y������y�g�gj�R"�#�s�4뾱6H/��q8#14���U-ѓگv��xA+�����9��y��~&r�N�˜�'9e��.ϊ�.ר�:��
Nb	
%:0�ͥТ:P<rT�gb2]�z���fY�������s�ڙ�UA�6^�v������O��..�icr�yÚ�:;�xw!#<o7�}ã�����}H;�Ҫ"��"��k3�쮷�j�n�Z�/��B������	��I����ڀY��L]�
A�uR���g�vp�@)�2pnӏA�8��l����t1�&�l�����BXZ-Þ��5N���b � �v<Pw
�訆ڰ/���F�\.�̳=Gՙ���g��@j�E�j��Bj���"�5R�2�L6�+��v1U�;�8o�/5�x����쿾��BC�o-<��2�$�!j�*�9G�0T��9���-fM��<�nN���+���i.� ��������y�g�>�bU8�B@8v")��^!m��"�SCN8+��A�I�LٵX8d�N{=�yq������t{�ն�A�qET��y ���8�hײ �q����.�ޅ�����5�c��&q����'"��(Q����U��N�{�T{����=T�J9Mc��jK���T��,���)�Z6�*��1��`y�]N��9U8~�َ�qy���9���͂��@`�p�X妻M"]� �5���5F�~�[����=�l�md���<Y��v�'=�༹�����!���Q~�ç����~��|�lF�#-���v U;>��w}���K�=Ջ��������N)�C����NA�8{$h��{3�F�E�r,��v�Mld+p�<'/:cxG\^g��s��Q�A��$�Qĳ�hG��]*�==W+�h�z�p��e�P��3S���v&����9��>�qk,:���T���p0�<�Y7�m�."S�G�����k���&��9i��Z�!Y?E4Z��}[c0�{2s���H9]�q�5t(LU���>���}|��,Z�I .�}~�n[4�κji�1��Yi�\6o[]\�zN���v�N������z�I��Ʃ�/���Պ�I�fk��9T�\bɾ��[�V�h�p&��U'� �K�h�$���4Xҟ�� ���|'�6w�#.�3����	�A؃T���4�x��Co���9��Y�5��Jd���Y�OY��ɬ��[����s��ql��.]��"e�B�4c|k7
�f7�p����Y����|"�O�3�Qb�
X�ʝΈQ�|ƣ|�̂5��� �� � �f8�.ֱG�q������n��.�zw�:��2y���c�0"a"e��KF���+�>��=U/s���H��q5��Tr����R%{�����T|�3���6>e_],=q���NUxي���Q�BY���������¸"T�ZHFͨ����t8���-�����.�1�X���rl���ځ�m\�w<tmt�2��� ����n~�o�Ϝ����`��1c�f펴u���ڵθ�[mc���v�:9��Yx�c���a�3l#4-�,�e()Y���a(������׳����ZC]mb��ԗj�<,.v`�	\RUb���ٮޚ*ƛf���p��~{�����|V{t'�A�l٭��*i�2��`��`�x�~���O���6U
^�DgB����+'=�O'6$@�wx��7e��Qm�vY�IY��ܢr��/*!�F��n
!S���g�[������Y���繜�d�&Lj��}��ɞ���m�5_0�=����9�-��01��(�-7�����{�t��{�{��+�੥HS�����X�������# �)2;��̧*gc<s��Ed�I��%�v�p9J�.9�s/��j�l�7�$1P�M(9e��
4��b*E�?-�^�_W�^k��A;�Y�"�&�����n������ %��B��hK��Wf�i�na���Љ���U�7\�Qk>��m��X���A�>�L^IAi�/�2�}ºjs=̼���Q���'�s��<�*�a��[�]<�!|�x��d3;�ތ��H��z.fw*`��`�j����ХW�cReYC,ې�
���O�ѕZ�^�̀��|��#M4�BD�<��@���N:fy|=������p�����v�� w	�t�jJ�َf��w��))�N�5ۇ"�ݨ�MG��x?�ޙՑ���y>Uyϩ��g�Ɍ�g3)�Q�/��Q̎�nP���p�*�@f\>�^�l�WMNg�;���B#�����独����܂�3�M��U*H&����E2��ϑ�K�e�ٱ�ܵ�Y1�L~��i�B�g�X����
��J>�?�=�*���iv�p����M��ٔ�Q�4f�J,��CF�����A�}�ގ�~�}�c1=׽��5��z��|��_W1�H��6�j�ҵ�r�82�1�M&&e[tzz�m$�3�w2��·�Y��^�o�vD���	n�ĵ�(-6�[!�U�	exP�	�����Cr�Gr��ꗡeGF+�]�'y7:�5{)��T_�Β(}C��ݴe�v��Y�d�UԈ�C�-�HU�j�Hфa�\���Ɵ�B6�H�A���{??>���VLf� ] ?�ñ�e�2��"���\r�V�fx8Ld���MZ�΃}^Wyϫ� ���=����D���Թ8j�ﰔJ�bH�	n��K3��Y�@�p�w�'xWTNg����y����,&]���{M�n�Tg~����RYe �~����.�3n�8z���:�;fK�&����jL�&�}����Y����!�.
i)�&e=O�f�d�t������4�j�A�� �e��!U��d9�7\/�z'����of�b#�R���'�u���7��w����w��Q��|1-r�D*�WZ�Jfp@m8V<�(�A�BH�v�����k�]���ǉ��=ub��9��S���"˔�F�M�n���W�<�9��^�yN�@�Pǘ�j����m��ݵ���<A4�Pr+�*o�'�C2}�.&���}���ڝ�e�v��Νʯ�����[� r�T�R�̱�|��5�]�nn����5�s|��5D��}z��M�A�)���h��}ܒY��Y&�P⁧i�T�
���Wq�����e}J��6-u�]g>�b	� �E�&T1̭���Q�#���$�uB!:w��_����A4p[���L���i��6�P�vi2�0j���xZ �� ��i"e÷{M���}^��s)�p����C��b����h�2x��^B)9�XC��yvS�ޮ��R�:}�Nj>��]^Ɍ���Z���$H���{ۣ`+�M���;�$�sv\7��l��PO(�1tcؽ5�k���9�q�NA��̯42˧�@���O�>�+k}֛�������	���|36�_O�3��y�> z-C�����������<�ns;�41�@<�b�@̧<{��r������Փ1� �w���� L����Zg'�ûn��t�.�0�V᭜V�Y=�.ٛP�n�S���l�щ,�K&z�t�b�:ә���h���a=��Z/^�]��,n�̓�JWR�9��ů^�o�[u���<T�hf)ڎ�8+S ��
��kCKW��װ�T[*���:��^�x��́��Zi��{�CS�`<Н���ϯ;T �mYB�N���u����+�R��n<���W��T6.��Ĳ=�Oes�3xvu��ɺB�_K[�wՂ�JR�Ψo�OA렦�V��>������m^��QB�����Eg.u�.+�86�m��ԓ�^�������
o6���Fu�#k)���w���(��p=�G)�p�|�؄yw��xe�Ӧ�n�N�G2����Y�Bכ�m�n���e;:)�ç*ɠ:~�5l�ègyS���!�kic��:�M��^^�f�Ar��ss�N�m�E\c�FV��u�6�0k1�{��.�;f.�w^���W;j�zg7H֪�Zm]wU��uy��-'n]c�9���2;��_=.^��1N�Xlh����pn�v[���W���û��=�[f-c,������®�fR9�@ܼ�h2��<<��dL,�S�|�'ʳI�s8��x�2c��!�	����<�� ٙ�m��TC�s�hLV]v{��5v�r�R� kkLfV�w��ٲ�3�N��{�*�K�V,�n<���,tEk����XB�ƛY�������}=O,;I`����6��y�b�cp]�VaO.�4�`W��D�T����� 
��Jf/-</���lhK��||����@�9���Y�'iwŰ[�������)|�˛dz���}y�� ���⴩66�|�#� ;���`vNv�D�v#����%���(�g�>|�v��׎>��8�;q�q�q��ϟ?����g���Z��u��/��#���Ĕ�[{j߷�ƪ��W,�]�|m۷��}z��q�qێ8ێ8㎝:t���ݜ(:N��(��)���o�ܕU��7Z�15DT��j�sB��_�-���K���fĆɽ��U��DS�ڪ�S�c|�O��t��wv�_�!���>|�M^�	���mi
X[x�FM�^ؒ�D	z��ꅒ���dX[C�a{�M螻z�޹�?r{�E�u7Ov���X��t��5�����|f
�DQlWCZ���q�/��Xe<[�F��c����������7��Z�hٶ8�㱦���j5m�xv��z-1���ږ&�5��(:ޑ�E%:��I��Y��Eei��&l�-�\[3�|}-�a=,4�%�ʷ�W��s�)�5tAڳv�8��=��1a(��]S!��V��,s�*&sr�	���tZ�q���Yݡg)���P7G��mm�%���+�yH[T�7F��3��w]xMa����ۣ���>����Hk�v�i�Q�f!�LjC;m0jc��Z3n_q�]6J;4�����H$ũ.�:��dBb����=�����s(�v��Yh�i�h�v��i8�`�m4��@����K���{nqWc����snoe������763b�D˹�.și��Rtp D�9�u��ݫ{;��N����k:��kOB���t�._�Q�ʘ��P�EKN�t1Y����m͖�F�`���`��c�ݢ�JD�Ò���YZ)6���fĺ�͘hg(�V�e����݋۠B(�y6�lLڌK(�i��)@�ͦ-�B�[4�^1Ai�'#v
����l�3�K�Ȕ�$�v�l=M��<������[�ѷ)q�7Dbg�\B��.G��u�7g��:�j݄��Մ>�r=w7�lt��GF��r�<��{iӮZ�ڝ�l���ԫn��Dn�$��"f�X1a�7M�
F�SgB��;RRͣ��˭�Iy��=kp�@�jU�r̽�����&�ݵ݀�7Ű˫�ז��q���Z2n_U�Ծ�v�s�-��Ԗ8!�%50IPn�3Q�ZJ�.WLCq�s.�FE&t�Ƈ��;DՀ5�k&��]^�6H���ϴ�SNG�Þ�zD®-����!�+q^�7W���#U�JL��&��=��*�e-9mg���c:�\`�q"T,n�8�-��͖$�L��\�4OY��v���UUUUUUj�W8�X}���/�\\ؐ���6!�����o����WU����l��ߪ:nm��FO~�����f����[��i[B[H�Aonc�rM��s�9������qR82�n8qrO��{W ��>U`�^�3�a��ɩu��eb��H��3�9��s�N��$2 ;;2Q[f%�F��`	����-��vS��lqFu�c�Y5ۂ�j󺀣���h��n�V�f٧����v������}��y�4˹1H����a���hEqY��퉫�0�}����8 ��;9.�JbcLݯe�Z���m�MSj}=����6R�J�c�N|ǘӤ�Q�j�b��{�������L�B3�����{>��k)��JЅ�����y1:�e�[Jm'b(�2��W��.myo�mfܣ��y�x,rЂ+�9�B	�eÑ�\r�=N}i���K|I(xI��q���ދY~WYϫ�,c���n����|hځb��'b$�Sc2��1C�����������)|c:��wuh���繥�A�\KB�.�e7<+�t��n�X�$�ȑPD~��5&2�l/i[��=��e�Sg��x�T^ƷԴ��rJdfS�L�v��o9�n��d��<=:���:��s�h ���0t�A�qET� �Y4��*p�G~��KG!�\qS��?��Wgcەcڲ;(h�ڷ���^�hd�ۙ��^���!y����e젭m�ɛ3S+]�������^���>p�#�O�m�X���{�v:�47���׾Ϣ���u���1�}��Kڐ��	��g����.q�r챛���q����7=�)q�{ʫ���{�Oo� Ը��Be3�>bL`	
|�D�O�O �74�52�<X=R)K����ݷ��y�x�Z�-���\Ϸd=z��}e���,��*c+���$��jQ�}Z��¥#��Փ�o�gfk�n=���h�i� �fV]��=Ol	R�R�󼔷��t�5Mn���sm�Q��:G:��]�su��A� O��_�K��/��z�8�p�u���k�Gzo#�O8��Vd��ɲ~Y���o�l/Ӑ�H�J�@P��<��j_�0V�=�''��s�n��n��d��<A- �N��"�E����K�b7��x�I"h�r=*���g�$�kr�^AM�y8D�:�x�+?F���uG�-7�k��4v�V��W�3�|�Q���U���j����5��9��3��da�wt��u�����#���B�3*������i��R��
�U|�,�\)��y��8@����"��U�#)5�5J�`*��E&FeyǷ��g�c��c`���^��~����bO9h<���pd��2�o���p}Q����,�^=~����`�e��hX���s,-Q���1LR�hf�-̭frٿ��XK�qB�ÑT��B�OM���A��7Yϫ��U+E��7����DA��x�B�uv��K��K��S�o{ d�1<�Gm�ͮ��鼎���Bf�C�K��¶�f;��`Ҽ�#D&W$����,)�^t�E&R��s2��X��;�q/�p�=��Y/9�q�A؂Ӈ�{����s���f_%xt>�dSo
N,}�鈢��|���7=&�9�q���T`�"c����<����R�5�Oo%�"�e�f���~���n+c��W#L��ά`�Ju�k�W2�a�f�O���Zt��M?��r�<�����6�[E2�E��M����w�ײŌ�p�#sk��zk#�O��eIƴ*�pᨷ�L��ȷO^�C�����>@vԌ!������M��ힻ��J��[���e7��|>ϼB����_t��R}��6�g_�%�� ��>Z<s�/�ѶH04B��v�X��pM���#�d�9�A�gb-2�̊������7Yϩ��r�Feر7��a��-�H�N4�k��.�9�	��4��O{��2=U�j3�W�y��b���N-�&h�hjp*F��{�{���1���fS����_۳���g ��O$%��7��G����
�	�N3�z���xT8��	��¹�װn{��7�� ��"K#2�L�=�}�����9Y4��~�ʟ9y|v��"3.�+kL�h�D�8攷��T����4wa换��a�U	�f�|�n�q
�e}:K1f�32�����,a����k(F�>��x���'7��{/��L$���\��r����� r�C@om@'b��tb�\�,�r����;����t�LL����`�O\�%�k�����x>�����v�����끣d8xy@�트��{l�:�X�A��A�,X�I�뇐�Y^��m�S��f�KW0Q�u1"����������<X�o����_���ǭ�fb a�T�LZ�-X]�
��b(�x_?�/H8 ��hh�!�?��27w��w��9��1 ϼ){�p �9a�훦3{��Q7t�y���8�y9�(�-��z���t_�=��$�� ���x1fU��]�~pIqY��"���2��5>%w��\�����]pnw��9�q���bK#2����"���Z��7i�����2��G^���7sw�P�4m��>Ԗx��<�1������ڦ� X�H�-eTz�8X�Ǝx�F.��w�������Ų�rO�KB�U8�W�cI2Q#-�}�{��Y��()vٔ9d��8��`�v��6��6��ј�=z�e�����22��[����܅��Z���%ǘ�y��&���s��s�r8� ��xL��Rql��sv���>7ކ|u'`�H�B�!{��w���1qa�Α�v�"���Ouw:�o���뵅�Wy�h\���j]Օè�޼Fc�S�uUf׬d�z顦�FK�y�{�,�����}���T��4�j!R��&s���=趟&C[���0@�L�*�R&Ue�S�9�3��~܋��G�A�A�3O�`kA� �ۇ�$��9V�Y���$a vˇh���w�Ahw�/'���j�WA�N�>��D[��3�5���x5��$����N�"z�_�7u��	k�dooY{꛸���A"մU�X�^a#�Go�HrRp`�������H�ܩ���6�n��@b�WR�b톙*
�����5�a<���[[����t^Fy���4wϡyRة��'SL�;��Fs�"H����,��~|_IS�N�_z���B��)� �N������oc|�(L�&p2����=O�)9P0ܵ�)�ȕ�S���������0���8u��Wup����Z�ڙ�A"TA�����9�����39�$ �@<��d�vvL�M�xtvoY{꛸�_5B�L�Hk=�V�,|�|���������gFy��� �-���<�m(�.���OLA��1HL�o^c_�5{���D�����7����*frx{؄�H�TmS��q(D������N�2d�;��ԍ/n���b���Y��a����р� >�~���b��;	J/0ln�Y{ڛ��\�˷������t�PƆ��
�y��>��- m,�J�Ⱦ�y�Ϻ�t��'fz+�zc}�bv\�������xN�=bZ�S`�ff �>���&r�u������h�U�eL�撺���+��7�J�L�J3ptn�Y{ڛ��]PYe<��B�����5�v�1S�A���Et��Ŭ�/-ʊgXź�K)c�!m5h)��l��5�h؛����X>�?���_(9�Zd1[5���<���b�/���2ְ�47P�Y�SgS���x���n�8�����,<���x������j�N� J�BeLۇ����޸���z3r|���3Uk�Rj���qcN��<<��F�z�����������#���y��u�&���m(��V�9���Զ�������S(tȬȞ����7�6�y܏{�6ۜ���&gI ^�͚��Ñύ��]�8�����/{Sw��BLjNJ�΂���2��8޿*��7u^x|����KC����f��%�����᪝ߛ-��t��Z�/R��o�u?}{���xs�1c���v�#'%�s�n�9�ީ5Ri�x2T�uk�������Ͳ��7qʸT *P�Bf��8Z�#���.�yF��1���7���$���M|��v�δ.���EJ�A��J]�/�՗��=�����k��J�[�Ő��t(�i�X�_�{���^y����{,��j����2�e]Nv��M*�퉻v6SB&담�ܗI�x��5c�qt�=-�z�[�'q�D��e.���m��B��c�ҹ���]�m������0�Y+�Ur�h�����<Lh!R���-���v�Ѳ�*eKA�Rd��n ����S�κ��X�-⣊�Ɖ�Q�v�3Y�bΧ���/�+O��Jef%��i�X6�cq�<�;1�Cua�k^t'Q憳�oBgb��&j��������g������P��A�q��tY�,��b̆�C�]c5FmD�缧U{�j�ٴ_��xsXd +�L����8~���m�2���mہwW7gj����`��}鼴��7qʀ��R[��Re74��׏�+�z=ѽ�,�(�}��Ӿ��g���O�+�GDZj���@L����P��w/Kh�C{իw����q���k5r�@L�v��x�q̵��w0��D(��j�\�ihHd�V*ܥ.�3�;��I��O<'�d�L�������7���\{a�D>N��k����f� �UH��撺0�R�wyy���)W}a�O[�aR7�U=���1�z��{M������8x����o]^��0;\h� =C�r�;U<Ȕ:x��M?���=��Sezz>��ے��c��$8۸f|��\*'Гky�ssiq��q�12���L9d�˯�r�/�G0�>��S)�́0)��i��!��cœ�����
&��l�Ҋ����v�F��{Дѱ�KP�{�kk�h�g��꽁N"����l���������=���10�E�]�s�u����M�|������xؖ��;�٪��&��G:tn$3�z�m��(!?<��崚es���}���tèT	�热U}?V�?3M�!^myن�9uAc�/E�t��5j��z���m(�l�?*��j�u��wk����&���􀭪�5U79�.��?��_+j|b��-����rSO\����:��֭��u���CF\���+��ͼ��yO����aJr�����{�J}�]7��V�_WL�S����؛��.�v8�1�n��:����7:Vh���ph#�pKyc;��u�Y�f��Ţ��u�.udV��u��<�]��`5b����j��ׇs�mw�4������G��3_VNM���ӓ��7$�rW!xndcWWf�K;Տ`�\87�=�N1λ�H�-Δ�U8�z$
�]���I�\,���M��t[��cJ�^I�/�]^BeZ�
N�Q���s3+��<�V�\}l'Իj�,��N���U���	�O<Ѧ�sw�#����ln(�XvdxT���9���h����5�r�}��5Ѳj�μcѨp�e�G�E��&�|����y-�w�Am�[r��X�����2�L�1���e�Ӭ�,q#��2��t˄P\�*G ᝵&[��<�3Ҋ��8��g�{���o\��K�@�R�3���Y@��O�!��nn���Fv�Nܧ6�]N��5o!��C����{f�����oWgVY���u�c�R92��tz�8�fi3
��Y�Fv�{YL�4T��8�w0�T��L��s�^��J@����j��hSwq,������t��+ZV#��`��6�o-/���7a�8cz=U�<���oyc�g�[���u;�����!�S�������${HB�`y��py*�K�V��T�y`��<T$��e�^j��~Xdj\�T$�, �X���:2v+@A�&MyD&�	���Ile���e��oT-#���>ƭ�x���ͼ��qd�Ū���ÙIT�:t�����ׯ�q�q�x�8�8�ӧN�0�D$�x7����.�~X�֪��X�ĸ��Y-�ê�[ž���f��B���-�악�	J�`�U#B�U��ﳷ=��������q�qǎ8ӎ8㎟>|�����7���ӵ����t"Yq&J�8�ў.��k]������־��u�����[,��_/fP�ʉ��hA�(�$/���Xu��ڻtv���폶�;����g��%��=��u���J��BMر��|X=ښ+ףGm�1��,Bەv8u������������z �5�%cF�^շ�XV�v�Pw��uZ�Gݞ��f����z;�˫�x��}.��W�:��`���Nll����LPI�h��m��Zq3�Ӊ���Z&�l[��f��]EA;k�~^��x���ڍh�����i֍1A`ؖڈ�cU;`�DmZ��:���QUB��B����%��)hȝ48pQ%ck;; ɓ&��u=�{�����{�1T�T�28Ƽʕ�z��Mmcj[<�g�f�}��Q~�9�4l<�����������Z@�e0�Bgl�:�Z�VT)mEFWm���x���~z���t��
����9����Tt]�"������o�8��i�<�h��rY@cv��°v�L���y���y�� �3~�U���v_���}淬�>WQ��y�gR ڻ�wz��͆N�e	�3ޣW���uÛL|�.� W{�3��C`���jbfL�3�o�oΦ�}��������S3m�y@]�(�Kg��>�ݏ�ܸ?y\km����#˽����g��� �xk��GoOz8ѕ�Tۙ�x�㏾��.5���Z:��q'Zu:�B������iNZ�x�-�p���"JG�A��>����dɓ;\|;�P�)�̖��ݱ/�MHr�k˻�}��΢��shm����2�L��C��Q�("
b�{],,۶뫵r�x��s\!4Ҹ�:0� �?������{��C�O���~�ڈ���~z5r��v=g�y{L�Be�<�[�j��Vgc���d�P��8�����l�ڏg���1;�ǯ<n�f*�Y���~��`kU=V{'��l�Hݎ̌�:����s[b��'�j��-4~����Dz|�%����^�fs���<N�c��qY9��)/
��a0��)�ʙS1)f��'}|�q<��#۷�n��g�����p.�]��^ކ�Ͷ-����d����1۰�w�Pf�����M���$�H�����1�7QL��}�`�]s��9J�P�����g�ϵ>�l��qVR6��/0tk��D��mSG	�&�"�bB���ｸ�������<��BfY�Bۣׯrjz��.$Ü���s�ԑ2	ͭ�X����i�HL^0�U ��)�R�3V��2:2�u�Ж3b%�Xm���z�[1uG�|���)�/lm�HTИĺ*Ԛ�2�Emm�A�.v�B��Kq�p��N��k��O4�z����>�$͵��S��^��>~�����@b��f0���l�c�c�����ˈxt��~�F��&Pew�En�;΢/�f�x���6�ݧ��i�Ċ	]��|ıU��Su���r��w?N�C���?=t1k��L����o�2�mm������L&V�s���i����g������v���zE!���{׎�nf}��3��eg�Ew{7΢/�f�m��z��ӓ�ba6�f|&zfbk�k7_��!�˪r�d��<N�c��\Toʃ#���*�pLM`�_O=K��!��i�ݐ��m��n��P�c7�ӷV��S;�Bu}�=��!$
q=Fi
�>�͚�ˬ��{�UM���ڶQ���1�T婐4�41��O*N�J�xW:�Uq=�i;��{d��czx�y�C
p�)f�U�S�I�˾�n+�%���"�7�,��N��Mm_��442�2o���l�=��&�_�{7΢/�Y�4l;kFuz��[�m��qA;��v[m	k� Us=��־O�Y�Lod�ey�99���|�<���v�B����O�gh�!_T8A�h=3�T�~����Ou?<ï�6<bkzk�3.�2;�-���f����ۈ�׃��L�ʙd�z{�u�
���:���p�ئ`L�K�ث�4@%������o�s��q6IIiv�Ju���vA�O��'t\�)C{�{�PI+ԞSzT��::;jӳx���ܺ�#.Xg�3�i�g��m����me%�-7��'~s�7.�2;�-��M2}�Wi� ��b��Z�ŵ�UW�_���NQ�Y��[��xp��Y��c3x���+y�>����쨻|p:�|�8�
gw���{p�K�7ŝ��;LȺ�nè��Y�>�L/�o4U&zU�	����� F�@ԛu
cT�w{���cӳx���K_�uNz�>�os�z��&P�vp&u���W�g˼K(z�������Yv7�}��߼�zN�\�Р��O�T$�=m��X�����`��2�N c]��n�F�����Ț�%��M13 L��H�을�/�f�z}Z2q)15t6o���e
�VL@>�}���MW�9���cՓx�����+I��N=?�o�M56L�MU2Z&^c�':J�Ys~�Xܺ���-Q��o1��5S�vF�.j�Bi7r(&"f��e��BQ³s
b7�D�8f������('��g^�7�(������t��P�٫�Fq�%VZ�7��+�
�Vf��F]nC��[^�U�˕°���B|�Ɵ��m6&W��S��P�BeL�M�T��~��V���+Dz�o��\ *T�e��/Hv�GT[�K�����՟��3MUn�E�޴gLr6�% �V�
:�
���_5�y	�2�z��7.�2;*͜+]����i����A��kn�e�4T��n��m�^�������ÚX�!�L�C�4���C����&Ij }�hU!�쪴�����#�'��>�S��~W�dP�P�.&�f'ի�o>�� $�s�|��Be�7�[ި�u����hKQ�sم��OO�`k4U�ח�v�u�����_���Ef\��|+0����S+Z��W��L����0H��f�kg"�u�p�vy�ے�K�9����3tr�[k6��Z(+�Q�;-�t^�,`�yj��b�9�{�D��?޴�ZRz�JV>Q�1�[��n��מx�Os{����8֛ZF�nJ:�7	��F�Ϣ�����8�F�yj��l��p�|�|��1aͼ�7n(䋘G��P��cr)�uq(0.�H�.��S	�i��{�\ g�'jG]�Ɓ���j�#��֎a2K%��/n�K�G]Zݎ%���i�)���k5K`뭄�b����uv���!�],'߿�߬~�����G���%v�띦��Ah:�x��3͒O�`}�� ;	�&Qc2���_ݝE�jo#�����RJRT]��3i��OT�6�q��v�5�w��/s�7.�2�
��/�m��S������g��UL�ֆqw׫�F؋�}��S�'�`�Û�p3���P��AU	P�s�|�Ĥ׋� ��{���I�jo#�+����֐�>���Nb�T�UR�%2%{p�H��6�B�3��/�s+=����ZaR�SL�V��*7��!1^��t�]mr�ǖL�(n�	�v��=��{�����-��hL��v}��yy�I=�
�9���_�qȐ]7�UmT�ƶ7T���Mx3����9s��KJ����)P����BÃMz�r-U`������N۸�����ʓ}���/�u]�?m���l9���CU?�9�z7�z�]dr��!�|�P������J�cxl���<|�e2���8�FwkП���[�UR��������Xҙ��/0��>�V�@����S]1�p*�����rJ�\+0����MM�y�6O��z��PHL��ԣѭB9k哛����u[sYoɈ�g�
I������M!%��L��i����X�Ŝ�d�����!�]���[f��s�&y'�?I�њH)�KQ�Y�6���1eg�:[��OV�3���	�gVH5E�T��e��<�Tw{Qb=Ӿ�3��IW��f����gZ�Qq�'�w�K�$�u�/�3 kUv��&y���^!�=��QB�}Uy��-�]��S!N����:��]�r��j4������mXY}
7�ӌv�Y9^��˭r����n6�M�}�fy��T��k#��oBh�p�d��ē��2��O�"bv�4��댽�~�YY��3 ����S���fX��i�Й�TA��[r�5��lћ�rJ��k0�
��������Iߥ���}v�A*�Kt~��,�k�krg��K�Y�c�n.7��L��2\m0�=���L���j��w�޽Gn�ݏÖ������*�L�mT��T��T����΋���g9�6�j_�V{#�1K
S1؋�X���ẙ�T� SUW��7g�ײ͙빺~���v��,�`�L�a��j�I�WT��5���w��f�(o�r7׼em��{����6������bmֻ2��$/�ŇKt��!H��K)���M|��ā��֑G_wycn�"�8�U
�wrE��������yW�ú�����m?���m��?���
�©	����M4DP����b�#+=���	��\L�t�}עωI[#�_�-4Jr41R�+���.��`�(����a�����ӭ��T�j�3=��IW����CD	���Y�#`O,��(;L�@� ��������� n!��|�nw�m��{���qZ}��^�ژy�Go3*���P(L�����(|�*ʩ�����dwW�|�*�͟}"�Y��{2=�����2�Ƿ:�g�*�]�Ú�j>jH�qk�T��BګZ�w���!^/������u�����j��ܯ�Ѐ��v�L*��
�b�w!-g�?�Tj��� v^�H@�y�՗�D�DP�R|%߂l��uz'6�;���VnF���[�.�D�.�|p��Hh���s*�fd6��w�7����nFU�}W[:U�I0�.��:�uoa�u�Ս�zgn���>���2�^[�Z�(�<Ǥ��ܬ��;72�T�t� =��#�dX�9δU�'`�@KhO0����+�wuӴ�ԫ^��1A���:�u}�|��g`vS�X�>��y
wn�!�Q��W�(X;c&)J�N�6�S2���>�̙�r�u��v�ѵ}]�q�2�@��b�ǁl�Ś���e<�dY�q����ތW���y"ȸ��n�]Ų��o�Y�>��olG��q�ܒ���h������b8xR��]}n���Y���0[ӕ��u�B�����s.��z��Ѩ��t����C�;M,ѻҌ�%��T��}�"*� �Ј{���.9I;�5Gw�3.,��k9�
{����]Z*eANt۷�p�Z�}|�-�|�v�ƬV݉�3d�"�ݷ$*��� ���!�p:���ۇ�ʛ��bQ��j�K��&�v��ۨ�qW������	�r�s|�:��/m�
��t��(K��qs������@����&�I�sM�z`T%����Wwb���oKyi"s���	J*�7I��M�{l���LMEu=�|����h�Yb��vߴ=�t�b�����MU��\��x
wt  Uc��1%�zJB�^{��yy�B-�zL�5�	�z#�cÇ$4��&�,(��WZ3QyVUՌC.�^1��*��)��>R��R�'���0�|�6��#�&�u�K��;|�Oɭۮq���
�;��4�~j��l�6x���j��J�Mc��|�=<s�p��jȈ�x��,�����q�&�E�A!GG냦�b�UmA�;���aѤ�r�.��f�F25G��N�>�z����8�8���8�N�:w��WW6���61�f��4v�EEbŠ�PU}Ρ�������
"5��?��ϟ�ׯ^���8�8�8��8�8���ϟ�Z"���b�6+U�}�<W�����Eh�TI�u�Ek;j��$��MN��t�cx^Ʃ��fm�֭��`�w�v����᮵Wm:�RN�1E8�b>�vk`�Z�V�:�kZV�ڎ��h�Q]��T�;4mh����&��=kz�U�����UF�8�TTE�.5���Ƃ&���5T�#�A�X��j�"��OGu��m���ꎍ|B5Ӫ	��]b��mm6��*`�����ֹ��Vؠ���ZsP^�3}���_#?vf�;���h��n+��3lk��b���w��MUU�b&#F�Ql[6��Ehm��֫m[`�l5v4MM��Z*��u�����歌k:#lFk��Et榃X�������[N&�j��*��C��N�4B�� Ŗ�	��5�x]�qD��36�Ac�Қw ��D�.�s��4�l���w�e���C��F����ۗ���^\�}n���d���4�8狶v�C'��R��Qz�&�Mh^�.PJY����n�ή7Wjܡ��	n��/8��qg���"pA���$��6��i��Vc��Q��v�v����OE\ ��J���ݡ��6� �&"Nܼl��i��n�W]�n�7��Y "��v���:�\*�\��>���kpg�w-�p��Qq���6	�1̷�̀�2Ť:�L���1��+�����8�n�0G����jٓ��m��p�x��l��c��kK��y&u�l����+��ڣ%�q� v��K�']�E�����ˬ'd�W�V���/%q��n�n���Y�XF��K�i!�U�y��e���݈��5��2�T�tq��Ks�ƁjER�Qͦ�45�1RhF���T����0ؚ�����:�5X�f=tw8�J'n =������8��p݈;=q'>�q��n���ڲl��63�����3A�öp��h�/#^i!��^5��e]�(JhF�hgq�ì�f�����j:˼�^j�Ί�:�v�y:6��K1�t�b�B;:�W�ٓ���X��E5�>@v��m��&�KM]I�X�a�֡��р�v��.ӫ��"��pWX�A9=����eV�'oB���4Ѻ��vKi�:��㵶��ZA�"���m�b��в�	(�lN3k�SKJ5����\�P�f���^ϗ�d@��[�=�N�p��8�6#G.�1���۶����x��x[;��<��&���U�����\6�I.�n�g�>n>�d��֭ۓ���S3O�s��;�ǯ]e�V���U��-*���]�6|gv��Z��Ά�գ��غأ1��n����Fc6��id.%��ӈp�+m�lr�Q�/<��5:���!s(�\N�:$�;�hJFb�8�6�2쥨#�j�h��2�E�X٬�������Xl��S I�ۙ�ݯgP�5b��ѬoR�ޟ��狼�������U�f��LkH �X�V��Lb(���7�V���	���'�!��w��>�W;ޭ���dt?S�_�����eL�2����{����;ucT ��c۝y3�U{��a��M|��������U�֘�(y��w:�S/~�⇡����Y�[�^�9ت��+�M^�ekU8��2�i�V� �SH�!4�m�7U����FV\�p�mJC�a��uc
�t�̄�˳��/u��{kA b9o�o�fuʯu��9��+���*��hϲ���Es��hx�N��~:���kK��p�лX飲]&�����m��	����S(L�Q��m�Ȫ��*��xk8�g�ɞ�5M3� �Hk��R���)o`��y��.�Q|�f�%;2�޳�"�-���0|^È|ك�}��s���W�+Wo�^�T\��쩤�FDZ$}�;�LYů�P�te����׷Ws͸�T���W��5��e���8�@s&���f_��7�w���{��7���{�}Y	���W��U!.P�^��S���`f(�7�ӏ�6*�=ʻД�z��ȅ���y��T�=u!S1�^*�k��Y�޽�ʻ��n�@U!T�f�牝e��)am��>����M�4�FZ�in�Bm���bTf�
[��6Z�O~}�~�=���Jb&�{�yy>�4�뵘s@m��<�ks7��|<�O��4K�����%�|�y�g f���}ە#}UY�U��B�4ɍ]��$�5���]!2�SL���f����P:�c/+}�"j�_��戇s"PU�n	ݹw�Wy*Jb��!�Y��t-@�,�%נ+�5m,����̘�,Y3��^3;���&�c��T���&V9 �G.�۫W��6o��4�P9���sO�Y�5��(����$3���C�f�4ٯ6i�N/�W�7�q�V��3��4Fz�ܫ� y�)3J��~��!m�M�e�������A/��ɥ�y'�Nz:�w9K���LD�\�G8"a7�z��y��ޘ�3 _�i�zo.�n� ��AO���ck���:�c3�U�T��B��Z2z�TS8�B��]y�j:n�0�5�İ1�B��6��Y�R"��w�raU3�5��j����YӯZ#}u9�U-�|Y5�5ߚi5W�E���y�ۮ3P�B��3�����K{���t�ϙ���2���惠��o�,Z�٦����꜑��(��\�ɶ��3�oq]�m�0��7^���t#��,[���;˱�U;U >cv��,�lx���5����뚎���9@>����)�km�=p��Q�/6��!$�!�!"E���O��N�;�)x��Ev�`�L�g��%��_;�p�k{����GV.���u9�U�#�U�8�`I$�@>П)ɘp��0�}��T�Vwᱻ�r�ge�_gM�e�\�t6㊤Qh���P�#��wɝ��V�I�ޔ����؎^�{��չ�ɫ|Ü��_<τ¶v����ذuC�MKeCNy�c&׳5Wɺ��S��4f�+��E�ɢ�o�ƚpX�(cT�����A���Ua��6�an���e�]Op�z��@L�V�g=E���;�yk�+ �f-"��*������=㖭��_c���!Ŀ�#ڞ1�x�)!s�n/4�N����>�ݡd�Vn����8�j������He��YkMԧ�K9��MfbJxg�.� fC�=g^������[�p���0�����ʣq�K�]�H�==:��p�x�i4�,kl�l%�ع�7m�7b흛:�G'����e�3s��u�N��@
���(�H%��V����VgH�R�]�M�!�Bh��q������&�����y��h
�kQ^4srM{ad���L
]+%����G�m"U��3νf�9}������qc���۞���.4�4�W(�.:��2{\�������\ �HL��Q7�׏Z棦��h�[P��ZIy%�}�n�騙�v���<���x�=�hj !�f�Mp����r�;Ѐ�Q2�]l�-�kE���ҙ@L�f?<��������Uqyy�꺞ḪD@>i>	�y@��I�*�2{�S����ץ��2������\�tվa͸DV/����7�ܛ��'�H�.��gg������0λ3׆�F���WBk�&e�=��X��nף�|T<�_=�u?��[�J7d��+���V�@�]4Tn�3�"�� �Vp�@��� L�����~���F���Jh��v3*a2���m����y��7 ��2!�w1OJoK+�N����}cl𕀽����qڗD��s����)������Q��U{ ���[�C&@M|���Ӵ��F��|Ü1�&�MU�8�;�=9McΝ�1�&yM3�y^�o�f�PgM���ٺ��*��W6A�Rf��H4�b*󄗍��| YB��S�w#�3/�u]�-���;�O�{'1z�+I����51������H�7��=ۆ�����fۄ�ƛ>�
f;��?Iku�w0�V�Vp�`'�K�k��A�y�)f�H���	C:b3aZ��I��)�f`L���7�K�l�V{�Q޵����vH8�kkd�P�U-j�J�Q��)���7�5s����`��w�ܼ�U�_
m�����F.[O��:���W�[�[V�R۾��^�(��r
��m+?���_s���!���w���A��=.=t)N�����z�*���	1�����T��2�l�zp�V�~��9�<�o�fZ��5R��B����ri��q���7S��~mh���@K�󥶤s��H)W�Z*g������[�=t}=�*72�=WXݝGbhL�2�L��I A�z�qY"��g�ebpq�E��:����Q�]��	�p�E,��M7T[��8>�����ÿ^Y==۲,Sr����_��[8�SeG��}@fC?��_h��u9���?��&)�B:�}`-?<���"ҥ�d����m���2j�aT�e7�|t�����=�y�y���@6�K�̩�2�9��<W\�����I�k�Mej�^���sf�I�CJ��.K���6���1VG�i֨�}�@�Չi�e��,d&����-�
�\�5���a{Ŗ�/d����MC�?�ij���\���U3��@U?�-��8���UU͝��?l�V{�s?�\�MT�P�+c2~ڽ����{��j�i���I�Ԡ���+��Q<F�R�U�%iZ�_ޥƽ�7~Tݱ��ڮ;2�=Y]|(B�K�gu{ak?%2��I��sn+{�g�/���O�����Ú�0�Z7�������:N.��ͺ�T��%2���ˁ�U<
V�`acJ9���	ٺ��*��A���~l�j� {F�m���E\z\{&��e��+���΂���goа'şm����2�&�3��]3\�yjYwA J�?_�Hvej�^����f�v~��>n�}s�Քlt���z���7�G���Q����5B��='��f�V�8���չ
����h\�]w�C���`4ǆ���?Y�s�g����?��[�=K��<"�lS�y<�J�����g^Ϟzژ�vy�Aϝ[���5ei��Ef�[*ul:gH��H������68F�h�wC�n^^xk�t�p�u�[�������Z��N-@U��:y:57�ȗ]ϓ�ǭ� 䍔�ڽ�V�ؘ����oa��/[�2b�t�IY@�lvqŹ���Y���\6�[�G��4�oVd�7�o�߃�.�홰F��ors4t�h�8�&ѵ+��k�\%bd�_4�i�h����E]�\��;��r�
���5�A����6��j��tf]�����{컼��u�sH
�3�Lxv2�#8M�n�T��A�s�ϕ}�g��ګV�&��m�y�vU@i�o4�L���}�j�ݞKޟM7�͉���չqsÇ��7��\!���p-�����W��6���l�j��6]��`|�̵d'3���v��g+���N���*�3��/Q�j*<>�P�!�2��N��#U#Z�e�A���]�N�x{4E�m���<޿�qJڪ��{�dQ�"�\u��L�p2_�-�� ���w�����
�P�����u�y�I��>��ޜ��
t*;Qf�߻.��n�=�Խ?#y�T'�E9XF��
�wC�zxW�I^�j)�s�\�������<�.P���:�\��b�~m5L4ʙı��U�����r��+��Z�&�M2�@�2�s~@]��ք���׬������K�/'0-X���~����a�%13����Ǆ��c���G��]-�ѱ��7����r�D�-1�:���hyU�'�~]� ��{��Xf���e5��f<��� ݍ�kɮ���(C�	ӧ%AED����[?P
�T��9����W�쮾���>����Mܚe
j�I��VF�>��3}�wk�z�k������#hyCX��U�i�ӏX�p�?�[���]�<�4�4���}��V?-��[��7�&i .��r}�6���ҥ�7�l�u��7e�":�n�6��^V�:K;�83�zpQ Z6���,�Z^�Ἶ챙���J�|�r����D�d�����7ҍK�J��x��W$���2%�*VQn�#"�7����3U_u�]8nŁ;2h����t�c�
���	O�vN]��+;H��T�c��ۤnm������5�}� �l���ďS���%���V!l)�or���G]�uf�.)F�w�њj��hu�_J��{w�d�]^���>i�pޭ�A#��@�#�^��л��a�����W����o/�aճj�wofL��"m[C���.T�B�B�k�b�jvv�zrf���pW�:Vp���ە2`�;&D�����`�{��y�T��M���ru�'Z���Iv�gv��I���v��3N��r-ݳo)u`p���u� ٝ�D�h��uZ�h"%�����F]߭Ѿ���_)�W�C�߀n�ۗp���G�{��x�l��mf��NѨu�L
w�;��V��n�@�쾌�Yu�uf��$��i7a����P��o�V� �����'��k6�nf�p�R�蛽=`��m�+OM���uu�������:%�	���ՠ�a��v�t�C �fV�W31��h%����=j��:�l�&���4jWZ��Ӹr�n]s8xS��q��8RE��x�-|{*Iq���X��w%B��X�32�>��h:�ì��tH�ygi �(A{w�#�-4+v�(�S߇�dX�U*�~���؈� �mֵZ&?�2Dlb�ح]��t���7e�%ʝq�6����ׯ����8�8�88�8�ӧN��ү�m4Lk���p}�{z+vlf(��EQtbj����������h-������O�޽z���8�8�8ノ8㎝:t���n<nҭ��N��h�h*�6�{�����j��k�LSIQF��ӧ���ѧN�6��kn��h��������˪���5�b(�8 ����b��d��:�|��8(��i�6�6=ٛ��"b-�lhj/���35X6mm�m�k4�UDW��DD]b**kc4E���+g6��Ů��1m��&$�
6��튪��݊��mPEq�3UѶ�u������UOcA��|�tjvq�`�*
jn���E��z�_x�/1�z�\A����ښ���ݻ�A:�V���E�w���(���:��&�v���ӱ�gA1CM�cmV�ƜEQkU_pi��8�z�D�����*���J�H��zBz6��w�b������V��<�Ɇve �3�d����i���9����W�쮾h#W�G��[���kҎ�@5P9��MwTF�#{|<r�6<�;s��+�����1V�yC�L���.��PFC� �l�� ��=|�(_����IZ�-��3<�}��qۨ�:���ʝ��I?_�@t�&��A��Vz�v�*'2�ㄾmBB�#�^o���jt���5�3U�?����������=��k���\粺��,�~�*C��בޘ��7P*eb&lA���K�W���u�p�wy��<�i�2�e	��=w��z��r<�1��9���訜��Lf$�]�!"{�6O��*��g�0FF�0#<{o����h���&'Ʀ�f��\���ɀ���O�#\�	42}hMP�CX�bޮ{A�P�ֻ�v[�w�����1dp��+��__+*�#*~�_��CM����{�e�_#�ҴJB�}���U�643D��`\YX�o7�Uê7��y��g�f!9w������es�^��mm\?]�F*�OB�>SX �j\g,��eij/-G���\"�� ���p{{z�v��}����;>��B�N�`YӚ_��ƹ��i��n�x����̴{���hoӪ���]�ԭ���v��8�8�P��w�i4�i��y��p�wy�Y�B(N��k��{��3�7ʤ5!��*�{+^Tѿ_�ED�W\pad��4� V�~T��#�:���n�S;��v3�2��8+<2K��/�Q~���"���G��FI;1���+��Τ���;�R�򫪖��d�I$+[jy���Ѝ: �ٰ>�G:���sI�w�z���]
�7].�1���3
Qmt�I��<�c���F\�v�.-�x�)�]�nT��9�����^|�`y�@���e�R$��ݺ>�pP�rJ�g�ӶK'E\o<�L�٪�sX���R^��FZ�@oj
��DY�q�g��1�<cѹ��U�b��>3��|���ݣ�*U�nخΉv�Ͽo��8?��b3R�;b3�\ʊ��6��%��4˟&�?3����SL�q�=��v��U�}�����h�șLZe����]&�l��E�w�y]W�w����	�3��|�-�`�v �Bff����&��J��P����]q�4öO�e4�h�r���q�ju	�mOn�흫�FUwmWn;3��9�H��2��2��1��Q�6z¾$<[�Ǧ��.���:��1V��y4�1��=�*��\]ӐR�o�p�1]tŚ�a�\�Y�1��{k	�mJ쁮�v��x{�z�� �ʩs]���۳�Q7���S����J��˵v�1�Z��~mo��Ab�i���"��[�M���jݝ��V��hcz�� 0��;l������B�2��Jy�8���>���?=��51b�g���jwt?l�߲2���v�	��B�:��aÜ��wh��jj�&P�&k�;�7�t���n�6r�-V�be4�1g�@K�U�����{8uc���D��%�N�	�5:.�<��-���{��+����~�Urk�C��o��<�!\�e3(L�9�ʛv'7�
������~�ʮ�p��z��ʙ���{�������yJ�$$��5���0�z�ع�.��0��u�H��XQ��1_ޥ�o�zP�Be4E��ګx��ȥ;��d��{��=��x�]�]�5Rj������H�t�]V�a�]���=�^�^W[��W��vv���g�m]�Y>�
�vt	�2�4�=6�y�E�gM�	����f��h��b����؍ϝ�f�,���A��k�u�z
`>t�>��]5h�K/�رdr�dm�m�(�o��oU!T$h�xi��W���4��3�{�M�mU�{�1�J�Υ���(=)e�rI���M�Bgj��F쩾1}gr�<ޟ�~���ˤ���ǿ�^~r'V%���O�5�� �u�M��Qp�*X��.�Rlh�8�����eh�5��rHL�����c�Wrs�{z=�hy���LB@L���i��������8�Fj��ګx��ǥ:��y	��1(�0�Jci٩i�kg���k�|z�>z���X��w\ǯ��_�ے��y{t���]��U�As6�S)�{/����nq�g�xW:�ƿ�]�׃P�qt������ݢb�[3wIݻiMw�"˭4'f5����Y<�Px�r�Fj)뢢�"�E�I\�ň�T =��A�� U *�P��!��az�,�N��x��ǥ:�2�Cc@^oU��	�u�ٔ=�C�t�w91VV"���ܺ��5M��P�԰Ùa6���mX͔Qk�;���|��2��8�B��v��������k����~���#z �Ck]���&Vg?���]!�Z�{o��p�g������e!�[�:��	�v��U�}���e~�W��l�9D�lռNfcҕ��Be2�_�!Uߛ����y�$��CZ��/��i�ب�������z i�ô�z�pP��=��X�$�]�]�l�8�^h6��O�{,�1b�O"����{/��=\<�R�Be	��r��ǧ�3�zș��\mQ���ݕ�Og,,lM�f��xr;�ܨ�/q���+o��:��巠�U���4�톥�@$�U,"%�4���u�׬KA����^޼�/�٦��Aq�����lG���q���R��6��Q<��n�����6�K\���6�ƚ܋����Ü��%��KMlYD���!T������jG.����f]!�kv9�(5pL�s�Û2�0�6��k���tk�Զ����ۯO8�q' N��g���]&�ؑ��Ҧp;mڷ6����߿�m���UqK��W����-�5c;���5	�h�)�V<��>�Z�e�ս{�1�{��4C�X��nm؛��B�	�A��*��b��t�q�ݍ�=�a�ӝ�Q99]o��-ʪ�s�x7hsO��^` �fH�M�=��.�AS�(_��~������/HjC��^����$r��U�'�u�I�L����3f�߻3W�s<�-��מP����Z�WsUy���C�c��{�n��𴐛�Þ՛��9�]q��-�|��v-2"m�m-�	�qZy���m. �cWB�Fk1t���F֥ҍf\ �.|���� ;Tʙ]�od���o��=]�X��0���2����R��E�]=)�+1r,�Bܿ�����1����FRĹ���\ł	r���#��w���-N�{��d�CofD؋C1pI��-��X?�oZ��ǜ͚W~��y^�y@u;8���{&jt�m�gi�3c�'����7�t��v�Q7�=q-�c�W�&P�C���9׆��b'�::�&]@&-l5��R=��{g�~̊��2�\��B�O?,g�ܜuz��P�Bf7kщ"�L�߽�S��W~��y^�b!&Je3�㉊�h�꧹@�Br���È�l�(�����ļOLc���m&��ܽv������3�S+�e&����|�ש��뎀�{�jom��2�M32�V��>o����D��AG��x)��'�goّ]],q/2d���_<��=�,"�9�h x�H
��8�*���	���XrJQ�KW�Ժ�\��sҊ�������t�]ًu�}�^��1�.{*�YL�Jn֒����pw+ͱ��� 8���ň�s��W~��y^�yLT�031����ƥF%���$�j�ʪ������s���T�����>w���i��������ZM2�9Ѯ�l5�����};q�M֧����	��<����3I(�!c������0%��Y�Ɔ�D�h�Ԗ�b�١�M9��8�_��5��>J��vpɦPomFf�Uߺ�W����Ă���f&.g�ń�[H�v䯔?�{�,��>����kꫩ��~jb+�v��z�p���2��R�M�EV3ݠ��څnWK��k�z�>�Mdf=Op�@��L�.ĳ�$*�ez����jN;����x5Rh�Ψ��3w�Ǖ�`�L�)�o��]��5����.�h/�`/��4�n�e}��{lC
X��e����ME�'��^�s*/|���i����{�w�T��J�],>.9�ŋy���@Bk��©5R:�^��yl!I�����{z7a]�eu�;H�&T�ߎs�9���� ��ܒwK�g(�p�֩WV�͹ [n8{ ��.ի6(��5��7�Ϙ�0��)�&\_^v(����Ǡ'�+���b�f�t��M�lx�A���-��\$M�Vt�g	��u�?��z)0�S:'}��ci�Rjgm�m���U�W���3��cz����WuY]o���T��F�3����3�s	̾އ�uF�^d�3U�4�w^�C�EV�c׻��S�n���ںŏD������b5Și�i�oS���<g���urf������ͳ���A̖3?��_���{T��A k��Q����������

(o�88�0|����D0¨C�B�2,2�0�22,0#+#@�Ȱ�0�0�0�0,2�2,0J0ȰȰȰȰ�0°�0,0�!"�"� �0��Ȱ°Ȱ�2,!�
��"�"�"�"�"��"��2#���C"��"��2,2�+���C"�,2,2,2,2�2��#J0�0,0�0�0�2�0�+B0ȰȰȰ�0�0ȰȰ°�?~o����C�� Ȱ�0�0���0�2,���+ C�
�"��"�,2,0�2�0,2,0�2,0�2,!�"�(�"�
�"��
�"�"���`�dXdXdXdXaXaX`XaXBE�E�Q�E��E�@!�a�a�aVVF �E�!Xe`XdXdXaaXdX`X`�Q� U�G@Ȃ0(�(! !(�C���ʂ2�40�����C*@Ȣ��!��
���X�G$00�ʈ2���0� #�T �a�!�d� �``� �Xd U^���XfXha`eQ`aE`d aX�.U��{ �XQ��``��`dXVQ�p��#"��02,�"��00��8VVFFF@��n�� Q��?�QVDR0@30$���[������@��_���?����U�����~���Q����?�(?�*�������'������?̨ *� ������a�#�]� @X@?�����������"����~�����@W���������ρi��zp?���?�N�x��H�r�?c X���B�R�P �J(B(R��"L !�!�!!���* J�(�� �(�" J��,�"�$*,�H����E��� B"°��
�((��
�"�
��
,�"�¢�(��*,$*,���"��, ��
�����%�������
"#""H �������?g��@͟����p�w�@Z����~����ǝ�������ۉ���� �C�!������i�t� R� ��H~��!��Z����"( �� ���J������'t���'�6y���4 *�ԇ��7�X ��� �����������3��a�p?@��_��A w���?���� �����CA4R~�����?�x~�%S�?w�6�����;�xp U�T��?�R���|�a��/�ɞ��PQ`�A��]�_�ߟ�����)ܞ������)���u$�,�8(���1��               � (     
  
         ( �   Ƞ$(I@
R�(PP �J
*T((@ �@� (�
@ P @o=R�UR*R�AH�JT�
�H�I@�$���$����Q)Q
��J��J�PHUHR*����   ��BJI!J�
m�c� }I���T�+'Glh}�{����B��z�o�J��2 d����U��K=*�5������ �� |    ��h �)�  �(J���9�� {�r6F^v��Um{׼*{X{�RJ��mKn���̫�޼�X��떬l{��=f�*���  �*@��PI
I@�)AKﯚ�/y�S�U\�S�*���s��[�R��UJ9��J�f�5&���Zn����V;�W9z͞�޽-[m�ۍ��)J�@�  �uo�o^Ս�{����X��R��Z�o9�.�o;���l��J�޻��*�x(*���i9�f���B�k�7,��8ܛk!@R���@��!I)QB�������-J�ڊUy5P��T������(���EDwgD��:�%�T�W:*�
n�T�d� P*��=  �NZ�S�T[��[��&�)n�-�;�Hn�	p�۪�M�8A�In��R�� ��@/R��J��D	QJJ��;8�Wv ����(�����@n�!F bu�8�@ m�U�!� �����E@[�  �� t��QN 	����9 2;� �� �rA���� 9v �T|   >�R�@J"�EJ�T�l>@�� v� q��Q�#� n�8�� �wX �RB�����(H*8   `>� x�� Y�$� Dq ;�:�1 21 8t
p -�@v�� �b > 5O�%*�� hh"�����@  OF�S)P  "{JBM(  ?J�����4����j$������x����?�����I$�!��?�n+�ރ�(���Ee���H�r����	M�$����	O�! BI�$�$�$�����ڿ����o���o�o|ж�V$L,b��9K6��/2�ɻ�F��2��3M�Z�v����n���Z�5Ұel+r��	���U��B��(�y���u�b�.iO^�;�vU�˻�¦ ��kJ3t�2��+�VZ�,f���H S-5t�^�d���u�/�80���۠�L/�z1L�ݱ�XS ��e�eI�.�bcŉ-��pb�{X[N�WƤ��ɡ�I���o������ĩ�c.��+I�I�"�����G0f���$�ww[X/.��p%X��cr�е=����S�fj̱��e�9�;�U1����fj�����d;yxZ�Cs�^���K�W�����R΋��z�Y��u���>�V.����# �KT��c�k	k�2���L<�0#�۰�mZ�m��*�)CXR���;�n�����ʻ�M�6�Z�����&���b��N�[�h�����Q�NP�(��E'�مbfP6f�E`P �E�n�۬t�1C� ���i��a�y�����2��UǙ�!�ŋ-L�%��R5���l�T���V7��6�yZL)*W���8���:4�5��Y$Uz��a�mH1V�Z��J͔��ǌ�G�״*C��#ڊ'���+��6�[�;�#fڢ�R9�\�.��@�2��yB.���;�1k�1·J��6�!����
���l��i��ka��ͨ�\˶2�����C���D��q��/�4��?�64 7T$�H -�qX�A���C�/{�;hm���{��Zu��ĥ�阁�.���m3J��T>����mۇC�6��U3���KdK��,�s/P�e���Ա�hQ80RpQJ��F�N�6���m��@2ѹ�HR�OJX�f[�`9�J��V����ër-���ux���6:��^�v��2���M�W�ch�sY���^e�+6�Bڥ�L����Vd"�R�v��;{��Sǁ�3ryvCF�X�Z�ո on��ũ`�1T���H�GM���Z��Ɨ�3(7A2C�y{G+hnG����,Z�[4s]�ݧ/#�ky�hl�u`��n+C#ԉaN;�4NL,m����]�n]�ab��֙�5i�
���Vc���f+��V�[f�;>��h-�Qҧ��ڗ%���%��A�)��*���xh�n�����8�1�`ӂl�\y�E�ͳ��f���ӣR]Lq��)r����Ed�*��5eʹ7+sq�ӏf�R�̤�s��Y{�'-�̬7c��n�j�
���.��=F:k:6��Vym��5����mX,�'����.R  `5y�����[���w7!��=ȀJ���0XJn�U�B�]c鮰C�J܎�v�}q���:`�7 �h�՚l�U�݌�T�ս�z����3l]l���8��EYt���4���uzd�_ajb��@Q��l��`�4�������4jV�ӆ���>I�*]b���&M��a/E��mD`U8�E�cFU�w[q�Bv�E��1hY�Iww�Q�o��FV�����̡u�k�5^؟bOp�D���mP�M !ɋiU�Qi��(����^lY��xGR.�#Yͧ��:�V�$9W��һ�� 'U�{.���u�dq��،K�ku`:僦�����T�#�p$��9:�[&�o���Il�$H��[�&�/oY���E���*�eՅ�Հu�d%�B^��^ПGHʘ2[��.��әM��
�0���#3s&-Q���JŦl�B)��˲H0m�z�`u��,���Z�h<�Vj��vi�,���it�왪Z[)L�Oe�6�^"r�F�ܼWC-�2	��(e��0e�v[U�r#D��cnv:IR8k\	{��난�����b�Wsi�!!Q��@��̵f�GYEU�h7�-�Vw���{W�í���X���>��k~����[3oki���xJ��i�/�)�{�
衉���&���ӗ!�FP��P�|l#W��:�X��v�&���'̠�U�l���6&�i���FڬB���.jy[�7d�m5�e�'w/c-�b��Y-�������J������C�4�)-�����%u��*XD���ʩ�T�_)�˶b�	��56�+�d���k]�l�7E��z-�V���7��HM�Zy"�w"5c���7�7u�dRQ�#F5p�����X`�A$w!.�P[t/J�Ԑw�4�V��#�����Gkt>�r�}v�z�6��l���t�}r�9*�^='�ֻ�_��y%�uj��rk��[7E7[P�^QVi^���ң�kl�Z^m�V[�n�ݖ���wՆ]R@T�9jne<�9w9���ګ����&E��(8�����)IS�֋��e�`ٺݽ�Z�z/��V�P@��H��N�Y36-�N���p\;��A���vjJ�M���^Z���e�+h���-��#D� ��Խ�)�M�ú�QQ�S�&,�xZ�(�NY���_\�7)AK!�`:�Y� �e��Ֆ�kZ�e��kFV���ڋl��&Q{z�5O��+ ��^t�� ienK-��gv�v2B��;约��m���P\�tI��-mX��,}1�#"�XPU�H�h#�ժώ�M��Uff�K�[�n� �W/�Y"]�b�v���SQܽ�Y�
̎��0i�$�����Ff[�	 ���j�;���2���
�h$]�����+3 �N��Q�#l��;��bǬ��x.�3v���-��Z5`�[S]��H�+1Z.�n��B��:��ͩ�E���+�i��ͺzZm���1a;`��TݭMSȪqF�e��~%�$$j6�J+b����.��l�+'!w[��$���͓o��R�B��v������*Ւ��M��������U�Q)�Vng�����[/n��j���os^�����݅ ��&�
=˧q:��vF�6��4[˧z�Z��m=�����u�Ы\����Uŀ	��rk���%�(�N�m�oF\��È9��%c�G�k7R��@�1e�Y�t@J va��t��*�^�Y[��j�R�n�
6��A{t`1T�Y6�+#�0���F��#-|V��^��:�6Py�N���r:��^�D��vf��5⦅�I�!yB�&���5Eokq��p�]�2j�VՐ�j����J�+�J�+]"��͗��4��,Fێ��h�j�h�m���.���L}�^	5�ǻ>�5?�avh��p�8.k(���6��Q�O4��n��YX
p=t��.đ�x4=�J�@�ܼ�%{T����^�3æ�ȭGY�9�6ڨ��d��	f ���V�i[�O��(H����ܒ�n�����
IV[�d�۬)�X��!�U�i�ě�v�E��7[6+4�8������l9���؋,�:*Ӵ@qco*��N�:G�9�k�w��(�[��*U�Y��)r�tB���+Q;N��	C������U-9�@�M^=��E�������2�X\&�=U�
!�(� Z����0�zd����m:P2�O���'0Re�M��f���&���.�Z���
U��"$kv�7.M�w0Q��Dh��	��`�Z��an��9�:��q��L˲�u,�u{R۽h�hM�����o1X�,]ق0�f�h7=R�N�B�����fܻOHA�����!�`@)Z���KH��F���[K�fZYzL_dװ&��iʳs��o0َ��;��фHԫ�)F#r<*С�t�Ghl�dŮ�f��6�Y��J���U&֣�~�	���Y��j�<E���1q�@�x3�T���[�������	��CK,��,�dc#�����72�M��rZ�W.ҭv�eĕ)Ge��,�]�F��2A�)Q��{��+<�YhCN��B�w0VA�s2�`Y���`f�t����ѻh��T�˹����u��� �?l`�s1L�@�k�r�q����� �q[���=�2�n��=�������F�!�����S�a#Q剑�j]kж���Bd��u�wh�̗y�0PW-j4`K�$��<�grƩ����U�m:�-�9j�Y�@�/�q<��f�I�(&h���&F#�@e.�n�ܷ6�oN�lMY�T�,ˇ�ec��5�17"��S"ڧZ�3�1��o{��gF,iĂ�dm�t@�#3&�9��uD�ު8M�r��)���b����8k,��c@Y4Vk�D�"f
�l�	��$j���P���֠�=�Thf[�8�r̻��f��41nÑ��-ۻa�k@�y��Ūh�ͤ�ȶ%c�1�����F�T�+t���l�KH�p��P��^ ����
gV��E9��P@L��N��7q�/s7A; C�<��ʶ��0��� �G.fڙZ�fa�720u5v��N�Ê�e�+q-+�;�v靭��:�#y��!�SU8��g�ˬ�N�ɹ�tl������/ic����1@�f�q��*�x�.��2M�q��M#L�ں`a���U�Y456P����d�j���L{y��3EIYF3V�Ą%��˙(խ�ܻ�RKl�RTq�Z��:�v�[n��˛�-������\�dЬ����+ ��Ffm�<��t+5�"��:�>rn�n?�k>�&�㼥"�E�֐{xi�t��V�qa������(KYur� U��F��&*.l +"�n��b�s1U�_jɱ�@�Z^奓E\AV��Z��a%j�M��w~¢��AF�2�U��IE�zr]��m-�mX���%)&��:�(q��yB��h�T��(IҪ��c�u�ޛ�5�/#;����Nl�%�x��f��;�B�e�JV��H��7se����[2X�R�%Fl��Ȩ�82�3c �IL&,VfM(�z�,�IW��+sh�8`R�%wiU$/n��t��h�V(4"�i!�:�Ry���{�5�h������u7En��6�&o�qk�l�ZI�0(��kd�M����m2���fM�}v�*�Y�Ŧ�ו{n�K;"z�s4H�)�_�lF�ٚ�n\�:����24c�F�0��0���[��i�=���R��4򮚘�kSk�օ.⬃7e?�%��ҷhV�J��b�Rԁn�ل�fLu��%Č�D�md�g7+r�k��R�&F�R�cw�e_ΐ�i�TW��/�f���wp}&��%��Դ�3.�V:l�j�j��6[��Wd�6���V��4�]�XJ��X7�QQ����2]�9e�3cv��k�c*�����ۛ�Y/q]a���mGlMu��w���RQa��b,�������(w�C)0��Ǣ�����͎	�!���SB�*Y/Iu�2�w*��t���=��NiS\��^�׶m�XGd�1��6�W!nm�fD��Ө=��;o�N���VbE��Qښr`��.#n��ѕ���sU��7�TkV�7���G���F�~ͽ�u��2�Q<�pI;jg���n��d�ش�3s+&7�q�-�.�e�$c+M��Gʒ�4e���ytf����.Z&�L���)���i����W�q�.�l`��*Qh�z��l*=��nK�iX�+5۲A�y��m�v�4diD�re�g6�(nTV%��F����J�A���o4j�+�E�X���`eWQ�V@YxU��(��+���+�������4e�'@�32����1��������iZ2�I_h<���ۭ˫4�H�Ĳ�����4�Y�e@�����kn=V���V�ɐ��ՠ�$$ �R"�\��D�fX�t
����ɀ����l
B�M�z�2���cA˘���7t�dy�����w�� �$�U�`WK%yjA��/u�V���7V�$�h��w�O�	�0R��j�s5�/�f(�E�����(���ǖ&���9J3O(����PaF�-��mV4S.����ɗX�%��ݡQ�i{4f�0nٓfc�����/J�;�i�(V`���5+�����q���{n��%a�`y�yQް�`Z@b��Z�
�)�X�̀c�A!��*ʛ����N}X,=��E�:�b�n��b�9C5[�vT�ѓU(��Z������ h�g
�	�=&J��L�e�gsb�+;XӛLbJYIc+sme�˅i����x��z�9��Y+��'(�f��W�6����a:)�,4M�z�������"k�^�s4�ch훛��������B>Q�Y�4��ط����D�nۛ"��sv�f���V�C2�U�F�����^`��W�*P=�ܺ`j=N�ͥpY1����[��c-�6�f=��v���Z�VT�Ҧ�8s(e^�V�DɁ��z���ݺ�``�Οv�=[:���Z: �2��lj�/l�'0P�.JBę�y6uP5)Su�X�Q'�Q�SYb���;EBI���_mLOt"��9)fjܬ�X�2n��v���R�-kQ����i��������T�,ۼ,ȷ�HLk1l[ܢK�t��1K�%ިyHjdܒ���80�R� @;��J��?*9��߬ZN��y�hk5^m*٘C��˺ӻE(�
��ŎdG$[��Tokk29��J��Y�36�H�R�������y��;�.R�#i�n���7��ir�4��i�ۣ:*�6�:����G>+ͣPf�q]l� 5(J�1V� �-�&S��f�@��;T5ZgZ)�[Z���B�5�V�*��#CM�̵���`z�b��TYyYA�.��%�٬_f ��!�Y�c.�%A���hԖ졏.$d3]���7(؈���{|��X^B@I,
(HH��I ,��d� HB(B��(HE!H! I @P��P$R�	���H(I"�B@	 � E�A`
B@Y	"�@�	@�@$�$��`H�$ Y$E$I)$�($��	$P
�Y H� ��( �B)		 ,�a ��� H�
 	, R"� ��	"�H��Y$��B � ���YHE$$�� X
H��
 �@�)� �� ,XH
E"� 
B
I,d	``  	 )$�X �Aa!X@ �IB����$���!	O}���i�S������7UK�v06�����K�/?���Á�S�F*�lG��ɨ���3�>7W�j�q�f�ܳ���!Qbf=5��R<!�q��(s�Y��]Xb��Al1� ��"��XAimLb�V�+zl��˛ܷ����0<��O/����]��1GV�������)���2�?�z�թ*�:�!s���2��&�\;a1q��*
��bˆ�a5U���������]ӱWm�����.��̕�ݛݝ�Jr�w����m��S	S�����J���7���������[P��`t���`\����>�q��e,9p����>�K��[]B�Jړ'��KD<ɸ�������Imө��L]�4�x� ��ګ2�j�7�G4,��[Ұ:gq����3%�F���#��hɔ%	�r�\h�c)ANY��]���Ý8�,hD�v��V(D-��YPX�X+
z�J�����,)hu�&�h�w(=�o#H���f��x(ަ�=x�g&񥝢wn(�Iɬ�J�X.v����� �m<*��{)�[�����n���#��Xwj�:76�O�2�b�m����r�6vY�iL�#�+��Gv�Jvv��I
���݁Y66��L������y���F7�H^0)�s]�d��t��ns�}+zŠk�NN�&�U��9]�I�v�:��ek�ζY���L�'�L�����9�m�YQ%����X�O5���*�:ك���rt2\Q��X*�;=Y��]g�B��a-۲]�w$�'Qי��\�O��}�x�J�6v�3F�O�PLt7�� �����n�s׶�pNà����#���rv�
l��o@wC]9��D40*v�'����i�]�9\������.b}
�� �� �ڨ�%�I>��iGl ��<f�=M�ٮ�u�+n�JvA�3�K���+Z�K�Ar�6��y��R��Xl��/tf-쥰��L���)v�zM�7�$"�^5>˭�!]�=����hȗv��`3m���NdWF�K�j������t�kb� 	H�Kw�����S��G�>���섛��xNp�w���W�M�N�+8sS�eaVY�5�9DX���rh�Y��^�|�맃5hӹF&�4D)̗]p쬶��-���]])wF~�W9Z�]#5U�T�T����H�V�ь��1�fJ�����`�UB�N�^�Yh�gKX�cv�E�w�����;Xr3k��Rq֨��/.l�\dN\.N�=�N��+F}�]�j��n��]��Gh`C9e���NSwoX��m���Ti:	�6����(��wV�8� ��.���F+��I���n^1��ѐn�4#j�1i���J ��*.TU��B3���Yٔ��x��vMKd9W]��]�r�݆�n�BdT�ޭ�W{��L>��jp����Ȇ3v�0�o.����V,���9
Y?t��o��s��,�R�����<? ]��,��^��T��T�u;whp�փy��ZM]b���\]��7l�y
������v�'��!1X�[Eb�k�1��Yu�=��+4+�c��2���O��9^ik7��5:���ˆo1ageZ�3̐�$캬�2jRϣVU885��<E�*��qL�o6�T��h E�5ڷ%R�<�i@iq=�:�B���&�C3���i�B�_�1�(,Sz�u��+o\�nt���ܻ�v���,3r�,����޺N�Oe����%Z�7[b�_k�*u�䍩�O-��LH�d���U�b�x�=����w,TwWl��l���fQ�v�[z�]�@���Z����b_Y΍�v5�I&���U[�����.N�K�}�2��奖���+
޾ve�9Vpnt+�Z�T��Pu*������ս�9��M���9�:6{r�אd��S��`�M�h�]j���ffuuK�:��U�ǉ���ٺÎ^�ȷ�_Fv�pWٗ� 5u�l;*�n���"���r]��2�����;���@�.HfS��/qj��_�hT�{x��=aݢ3�,w�p^�zqi�r��siq��<(�rk}�DCY�����D��\:���:�l�(Ğ_f��qs�t�W{��V�u�nÖ>����:�ؕ	�^=m4���D
�����3�<��W>���{\�]B��+��
���.�oH�1���Ҋڼ 6�n�Q=�J�wv�N��)K��E)�s���V�n�B��!�%Q�/�lL�=�I���l���.�_����5ӱ�J���ي/���4*�YrR9o�.v�s5rY�V�o�c�X��RS������ԺKY����Pցߍ��QV�Iĺ�19*�Ps���yx��ƞ0o{3ku�(��n��2r����]��-kb*��S��W^�
B�F=ۑ[�x�ĕ�F�&�a�c����^A}t]�Gw�_U��l#,��od�W
��b���709\�0����x�`��{ݚ.�B�5W:�nf�	I��L�3r1(e�Ѵ��$ZhӍ5a���Z�+�ͪ���i{�q��A�՚��q�s���\�l�8��y��0�Iu�O�c��F^��_~�gL��ֳ ^؃[�k�4��D����m�y�:6vA��	7ۻ�Aoo^Z���ѓuƛ�K�S��r0֕}�m��wu����&xi����p���auݜ
4q'���.Ч�N�wvT��r[U�c�����s���ySZo�z�<$�T��vŽ�5�ĺ�`nV�6��\)�<Ʉ!���v��]�Y�n31����gd�+ٙ�
�E����Yt�4S�����y�6F��^�km���d.Ʌ@�F��r� RGm+w*��n[��4�JTJF걛d���JW��p+0���
n�53�ޏ �Ne_ӗV�T�t�|��׳�Ƚ���Ft�Bܳ��~#i�8�'R�c��<YY�qL�tHomp�<�܏�G\�g������MY�Qȡ�0e����v͂p�w{�)�Ւ���d�W��S.d(i��1�t.3$w3	���u!�#Un�j��jN���R���΋ɹ���]9���r�\iQ�N��t�X�w�&f�����"�����m��*C�.��3v���B��{)�*���D`Y]Q�oX9w�J���V3��� ���}�n��ծkh]����Q�5�G8�8�y��[�Y%��Kef����m�x��� ��]-˥ؖ����������`��h��S�pA��h%i�6��E&�m/��LKu�.�w����S���R�:Z)ېҮYV��/�hs�Qۧ�,���r�2�i��^�g�Ʒ3
�˄gV��}��{��ț�4Us���~{\�8);�ݸ����� -B]��;Ӝi-��aŨ��;�SҶWb3�l�Ņ�IBu��#�l�H��e�X��R�.kI����Q���&JmU�a�ف3Y3Q���"x�ͨw"��v4�I�"p}Ӎ$�`����Wsu98L�-���c���&�/t�в�Fe	j\"Av�)f�f�ma7-I�Gqd!�JD�z�;�*t��|q��A#3@�������
�`R��^�d3{7���{����d��Y�ۻ�3�_4�;r���\�q}@払���_=;AK4�]K���A��)�JuR�̫7J>C�2����faz���fN�U�-ތ��>���e<���AY���_-6#��AXIA�:�cyN�3ye��+�nu�nE�-��/D�5�t�1#~�H�;R��!U7YN���si��r�{\��b�J��d:�e�(�I��d��\��n^W+Y2ޤ4��ʰ�xn��n�jC^��@�Z����Z��j�ݷg)6n�D��ˣ���`�Rf�r��Yٹj���+q1f_u�1��`Y�Z:���ɷ��3-��	���᧮m��M�,FpR�X{M`����<� T�郺��b�Ժ�x'>�pg���tG,�z����Ĭ+"�׉��`����R��R�m�Oqd��N�VMlV���K��C�i�(������t���n�H�#歌���A9��w���#66XQYN;�zh��%��M�9R��g[�|��[���$����Y�}���}k�u�I7Z�z΄�+l���S�#��H��VLΜan�)����cir�z��_g��x*�����n}���PT~���sf���TI�zpʱ�16�L7�/������N�h˝y+1luJ�l-�]�vb��]��V��3�^m���v6��m�Ʒ�ۗX%M,��vZ���Gv�x%��n`�Gn���l�k��~���]D����c#�Z4|��c�f�6^�oz^�^�W�n�(k��p��j�í8���f���ᶇ^�Rp�3"�[Œ�uu����K��ڼZ�n ^\�DPh��5�'�J&m^�C:�sWw��Θ��r��j@g47�S�gw#�=��_'�mP(���Ùիyʷ���n�6h@��[�U�pA+J����b��h��p>���)���S{M�N�]�R�t��6y�Y�Peh�\�X[]��V�&�y�45�uҖ�cI؄�i�K0�R\�j}�B�i�[��ڴAc$7/`M����]�c�y3�q;w�͹����6�!f�W93��;��X^=��	нn�0b���LB6�mUkE�vbq��N�M9/.�tY��Q6����}7��_P��@��6�6�K���Э�V�M�:��ѯt��ar�q�D���
ww&��y�̴[�z�j��4�"�j���c0H���R��5�ν�&ԖF�"'��3	�Yc6]��7���gi#7g*�ߣ��m��&�j�a' �Ċ����I]`�9�j�9�e�Yws�*MaE�ӡyaZ�#N��P���2�<�t�c�����xC��"2��I�r�x��d��]h�Ʊ�F�v�XO&�A�r̸S��2+Ѹ�[O/UeV!ͫ܌2��Ύ�ր<.ۙ�%�G����N�Z��e��8g��-F��x0����F����-��.��e�#n�:�7Eoc���w�5���%�Ո�e�ۡ��},h�J�7�:�0�n�����V2�޺ΦM�23hU�F&p:�h��52��K�J�IT���F��Ѳ���f��u�C6A���ո���y��Jf��^�����:�%���6�e��m�Z1��&�Z:`:r���]�30�6X�̻�g�m�}��]��3s��r�k6`��52�m�t�(�1�a���������T��]Xo�M�����3_��vv�*�"�I��:à7Wb��*U����r�M��:L�U�ܫ�������vK5'e�4���6����y��P����f�w�V8�(��{��b��pQ���]�'̛� �V�d�gWgt��,�r�<D� ��bj���Xq%�L����oz��+iE șIͷg!�R���^Y�au�%^���u��=w�L2p7P�-���Ӌ��VT���o-���������n@�ta���j%��x��z69J���fbj�q��E�g5F밣@s61R'{c�*������]��T�DgJ��v.������Ĳ�̑ACI�R��0F�cn�嚐�0AZ����i�$�G���������5����\h]	��z��df�y�t%Vm�aؚ����sTZ��)z��ȹ�(���A���Y1�ެɩF�n�������k��YO�|�s.�Y�;(�
�1s뜀�]5���IR2�ĤF�7��26��ךuˤ9��8j���DįM+�لIK�n�����K�oP��z�q����'Io�;��X��H��f����X��]M�tcə���V�,�,���k ���phC������Y3.��Ԍ1�V������\W.U+̉�����t�0�J�e�NЌ��8�����[V*vb��K��_uZ�̵-Y�&hq�顛V��Q���(��A`5��ˁM�~ڧ�fqN
����%��&bw*��[@��Z¼�
�;�YO.]c�^�6��d&Y���:i/��+�'|�Qj�����c��l
����sˣX�ѧ_Fs�hVClQj�
�R�K[�2^�"r�{Vi�P3>��p����TIA���s���<�@e�]�@�LQ<��$�\U�C�	%l�WD�؄��Ws���`���.�K�^�u�]ݮ� s�Z�=X%pZEM��o�ރ�<�RU���N}�o�:�9n)j��k�����w8n\w�ݜ�g���%���h�NL��܂�cR\F;;�{P���HuƬS��9#1�3�/:�&2���ۡ��^X�o��w+;V��u��a��z�F�	�WV&���Cd)u����Q�qZ~�⛆�z�;5���t<�f|�Y
p)ڽ�c�9�`��f�ZY�bƀ���dķ������7���p*�Pm�B��7>�^�:�]�F]u'���
����F2�[��\�V���%����L@�X��p��q�7��^.VAIv�ź�9/��q=�˲��uV�b�r�C�����U�H��Il��.O 8�}o�v�`���sn��bo�f�Zsd��l��;t��ȬqӀq�U�����N��Vu���N���,_^��r=H��{,�$���V>�e�s`�g%�Y��D�f�e�*Lz��{�.�fYˡ�J��c��U���f�^`�釨1](���jK��WU�m��ge��Һ��\8p�����:M3�g`3w.ފ�p�!��\ED���l����Qǩ`�|��.��
;�ݳ2bR�,B��
�.8�6dBG�+�̵֟��&��}�-���]�M�5;z&m]52�N9cl�e 2�uf|l�z`;��+\�j��-h17Ҙ㖥�n��vR{&Q`򱉗�t�\m�b�V�ܷ��O��o݆�pώ�]&���@D��}w�pq�VE�@�4�v[�r���dD�3�Y���V�[{�y�{߯\����g9����$� �~�]�n��t!;����77K�.ۙ��E�����y3Q�M4�kd@�x��x�8�϶�oC��{6��0����R�kh�Ps��G��z����\�浼�g&�wpɋhd6��6�:�^�ҳN,���T�-�����"X3ktr��4l������ɳ�i��r6���$�ZB=���*�	��jV�����֑n3(�%�\�f�͖���"�	f�G����+5���[�C*���ڶӵXF�R�ocv���"vYM�tӻq;2)<�78���$K���[qq��ޞ80�a�D��{��=�M��'<�Y�	,u�X'Z�"�񜙍i�N��pj�[1�.bV�D��pt���#��X�k=�7�7h��=B�ٙغW4����CWMww0������i�-�r����+����J�A������>o"�v��3`����ɷc"��˂'����uJфะ�7v�T�b��Ad�ř�fi�Z���=h`x���Y{+��n^
�v��.3�ڞ�̫�<Z��ڤ0uˌ��2�hP���[Z����\��n5k)�۞x� �v�{d΂4m;8y�36��e��gfZ�P��[%�
�/C���.9��ۨ�I��UnoO,}�!�jK��D���]�u+6��ͳ�>ķ>�D�Nd�e3�؈hU��>�\����3Ǘ��3�
��.e:�ϭ�F����,�r�<a�
�=����IZ�.�sc+5Ա��a/C�����ic>�\���y��`J�[�t��R��nܞ��ٓ9�_>��8�3�9�8H��N3�-��xZ\;C�3���=AÞK ��x����,V���N���]p�;A�H�2<����)F�m��#S
j�m���ى㵚Nwb�z��v99�bMd)��ik
�Ye���b�8C�����,��IsM�b�c�e�̗3L[B@#��%gn���@u����q�1�i�m�mK��X�݃y�b�g�w>ǃ=�b�Q�ے��o>�\]+ʤ�h�:z���5�u���%��;�u�qN�][���2H#�nt��c`L9��VMd�[n�4����9:Rsq���8��x���V� &z����ɬ��a��g��m�C^��@B�ݚN4n܌���y	N-��l��)��F���gX��eE)��1���Ru��1t+�KXD5��-�`H]\K{Iz��ίb�;+c��M�Z^�[s�b2mr���F�Z"ڨq����j[���ʖe6���-X�S��vugd^<=�ؗe�S.x�u�#���$̮����K��l54v�J&�h������#ͭv�[`���vN,,,]�\#�H���S�����m��<W<Fnu�ث���-l �&u�*���X�ԉF�0��.���5c�O<u<���]b����YeEh�Sf�e#�uRF�]�IsJbi��X��2fn��D1�k�n���n�m��A�i��ppnc����.8�\¸���͑!��`�,�u�+6�2:z�Y���RQ[kfR� �˷i��N�����s��u\��Ϟ�1hB�5�\SQ����LUn!N�m�q���E���ͮ�P��v�=��^MٛP�	d�6Dsno-�ěY�(�eav�k��熗Y��n����Ū-�YFs\����n"ƹ�ۇN����K�K1��3S�Ֆە���r��m�y۞���6�;ygX�1�5�\��:��!6�Fi��7��nW.^z�<=��ˬ��:S��#�v�SP��`���lT�H���Q����fڤc�FjM�ū2@��.�k�9۟��E���<��VԺʎ4��>hl�Kll#���n��)��BCn���+�؄�N�!v��B���u]�6��m ��ac {h�s�q�����0����lI�QR�P�nMl=p�Nv�\��:w\�v�n�AuuФv��\��ȓ�{d��ha�n�Z��
X%��Ԡ�Q�pWr�kf�"� �ch�M�0Q`χ��,o$��[�����B�&ա%�.��XY��Y�F�I���`.�vM��M�t�����vA�Gۋ�Ӆ��u��Pח�5�l�΢���͠.0MKY��\�{]�B3��:�'%������BWX���H�p/0qN,m��<����0¢�݈5�ih@K�t��R� ���^̰�#e�N�n�+��9E�m8�u�F�ݬ�p;�Cۇbl��Y����5{\��<�ю�ŕ6pt�<g�b�vBh�F�8݋�C�b��p��(��cj�lq��ye��lk�U(ي��e-�\�lţ�a����1�+l�SA�x۲0�����u���Ρq�7�\�B�8�WV����toi�<�\qwip+��X�VZMCXc(����es�Z��MZۘ��z�v��y��b�#˱���O'�ٳ��]�=䛶{nP!g�v��y{e�Nܺ��o<ޓ�t����]�mu��G�`l�i�[�jE�cU�u�*l쾍�Z���NciJ�ٷV�&i��B��6�D6��m��pR�@텯D��gpW�v�)�{f�\�vr�|�;?n�N����7MF�W�^�v31��,e��cMu1�xO<Ѝ�����tf��֌����h���h��h�����#���1�S�\�M(�Y�	P�����:��ub�'<��V���lK��f,�B]�6�E4d4��hB�l �����['i�G�&��R��&��ی�d��ҔL]�:�����h���t��4Cj�	M���Zh�3(Ӛ\�ܐ�TSL�"�� i��y��y3�0׭f��<y�^q��7�Q�q�ݜYє:<vժH:6Yk���i���F�E&j��F�V@i�.�@�3�8��#��Ӛ<>F�Ş0k0�1��Q%��]c�Id���,�
�́��݃��)7e�8=���F�\�� ������Yn�X�X��,����T�9m,֡��ι�����Z��gq�YݤL��ok�^q�h@F�^�ӝ�9q�i�%;pn�*Ns��Q�;�(c���������G�d��s��J\�ǜ�MP�5�ٰ�Yv�aM�kaup`2u����.�f��f�5dҰ���q��2�[�T�]�6��0���L/9��l=��q�u�7-�f�bV8i�0Rl��B�N}�6��M�֜��y�D���&�m-5�Q�J�;���C.mgrW=x���5)�e��hEPf�i��7H�A���Ȓ*.3*�t6Xq���[
���K7�u�M���roV��a�N�c)��v��7-��g�<p�J��;H�Z�8L�1�oX뇸4�u���8ݓ
e]�nńe�jh��l�ff���X�8�� ���M�j���RP�Sm*c6�S;�n��X ���K�.(��-���l���#3tz������.���nA�+�۲n�=��d�v��;<��'NnrF{+�g�������\�[[Q��;�J����hܭ��n7E�.u� [�Z��ώ��QS4sl�vL��S�-Q.�ٖ��̳������a�l��h�fù�
R��<�+en+�F#5�7Mic��55�t���853Ih:P��(#t��(�P�"�L�-`L��x9@�WL��n�i�N�Ŗf��솻%�B��2D��b=���2\������ؾ���Wi����䦌�'Nm�G�����F
���0�ծ����k!tY4�3E�n�3��/��v�U�0a\E1�]��L�1tլD܋�_���O�۴�
�u���Ƹ|g��^Ys���SZ�E�4�PC/��q��"�en�E��%%�'�Ir��%8�=^ݶ��j;e�/b���ۗny����ýh��2�v��ↈ˶�s�x����BE���9�`y��ټS(���l��>�v�����:y�p]�D�Mg%� 2��a�6��<ݹ���4�뭘vh�ѰܕnM<��"����PwcsϬ� ���Y����eN�4\����	������Oj.76:J��q�k!���n!{M���՝ی���
b��E��K�pL�j�,�$}��c�jZؠC7cv�'\�\�F���n,(�'���,�>9�,qt��-uıCRk4m�7W*n�ڱ�͡���)#J�A��ݞ�P�.vq6��o���cr���
�E��ص�v[&���|}t!k��I�g��N6��ۗ��Q���t�O������tɣ�^�9e�_wB�QaVU�6��{k�
X:�+uk��	���h�x1$6��K�LO:���xcE�ۣj<03�^`�h�+�e��M�ai�����.B�0���u�p������S���^���Õ����<m=LRR���	ʔR�&�e�桅��T0E��:	��Ԙ�^졢�Y�99ԏ�//��n\t�=�͵��k�i�Ѻ9�"(�n�n:�ȁ^���/)�76��q�X"��db��U�!Ml-S۰C�dT�r��9Վ�����&�F�v����ڌGi�o!��e�Z2��6��������1�4kj�f���ո/m� ���g�w��+�����N���+���̪��@�5���kφu�����}�M�'���q4*�`/ѳ��Y�2M��dIC�+���#>�Yy��^qLl�A�n�7d�gȵ�-jy��8WXYL�X��2ll2��pR�G�m�z�ݞ~�l��4L{��h�b
VL�=4p�u>�u�Thh*:[��� ��[B��.�F0ލ�-��!��n��8�e��pφ9,k)Xx�S���6�5ڭŀ�z�����͝�۫rs��L��i���X5�@���jҕ��s�!�I�Km��%�n�k�u���K5h0�b�S;դ�z�;u�Kj�l�^��s����9٪�Nf�����;���Ik�wQ�Tl�8�r��1�s.�9j39������
fZ�W-�w{=&4ӭ�^�MU*�ƅ�Wkj�,Ʋ1]d��oi,�1]<��,�]�N5)�*B:Y��a�f�9ULҭi=X��0��Zt�ڧN�cee6R����p��u�Z{�3y��z�i���U��M:�-J�1�[\�����MMeN�sK����g�5�{-�)�5���s��[�fV��{zp���j�:X�=x��Xi��2N��X�f���=뷌���jFĳ�W���d�kI�[��憓iך�L�q��j]V��gLZ�͆�s	rq,�84�^nZ��Y�3�KN[G��R��R�r�:���SUEk6��&�5�K;9��z�f�qE�vi��ׅ�Z�i��Ѐ���$���Ķכ���� ��W�|��y���;[g5�	L�8�hqĨva�Y��k5��#�\Ҕ��lˊ \KP�G�nzNgvn9����Y�^�3m*Km�n��pX��h@�h�l�K�[
�\ܩ����	Ѐ�QVu���(���ԡ�5��3˱�<.��u��6�R噥�,z/WA���e#�8{f�m����mB��@D��G�����Nx�ǎx�^���� t�3��S�m�VՙW-��#�An�nYI�v٩�Iy�J)��[�1��#k�a��d%ַ�녺��ը�i雡�΃'</6/<��_C�����7%�L�TsKn�].��Ÿ���y�;3we���XRc�VScL��Z^�a �GjL@3k�Zٵ*õѕ5l�9�.ـ!/!�n;ri���/[nl<�>+�J���� �a���a� ݣ�:�R�X�f�fl�,�YbBme���+٣c(��l�AЍ�3���9v����X��7q�2�J� �y*�Ա���퉗f�6�3� 醌���E��g�g���n4��(Z�A�/�����n���%.�
�"Ce��0���燒�Ɠ%�)(��T��L�6ۚPK4
�]3 ��Vp��@����<f�
2�j��m�F�sa$䵄���lix�;qjۚ�h�0���"D���t�JB�)2ͱ6�)�-���\��ڤRh�6��b���vY{=�y!R����L6 A%�ˮ�č�Zk�h��9�96�ٽ�{#��k`�9�;&��p9���S����5�n����\Y�	����t��➻&��]�.OP�5[m�4��-l�B`촥�Q�js�k"b�8ԅi���vv�S9���Q[�� D�\7l\�2���6P��mvD�m�����3�� �l��n#z��֑m�S��[y�h;�v�󺓛v�`c3�	�͆I�Y+�c��r���:I&�q��遼���m�����Dy��w�xLc#��;޼�i�J�y<��:��6��hM7bv5mt.����糍���ɷaG�o2���m��G�s�¼{���9�v�ۍ��^�^�w@!HlM�.+ǽҭx����z�=�V/e����=�g����?���:�^�#�<.�)1���Z׌v�|����2���c3r���/~���*\s*�s,���f�߳�Hܪ0�"��cѿv�+�2c�Td��H�9�	)�(��H"Ѭ�7Y�;:��} ���݌��V��=�P?�A���%%;��saT�Y;�M9j iNBR$�I����#L�j�R�z�M�nl$z�(�?c�$3��|R��� $�P�誡ݑwy����oN
R'�ر�8��4n[��8�ٓDu��Җ�"�?��~?-U�Q�JP'��*R��	*�i�����J2˝[���l|(�l	�O�IM	H�7/�mԮ1,	�#^��بpjq���\���5Ql�Z"��4e������{\���BQ'�T*��nd.8}��3I�A�4{V���7�i�]�:�O�@�U@�R�$_e�e�+�f�0;-�>i\[����%�FY3~}� ����$�w��?t���3��H���N�HJf�gA���y�3g>�vO���	�rh��p���;
�x}�ބfz˂s�}z�yU�d��{F���� ��
)D�	Jk��f�l�s�r�N���{6>��`���IMR�$%*���{������ԉ#z$�BJ�dfb�u��w69�J#���УC��6��K�?j�C�����BJE�	 ����.NDK�z̉���cj2�p���;��=�4ށ � ��IqF\���T��Ӛ�ffb����❎"1�=MD畸]�,��\����e�l=S3J�|A\+�
)D�	J��%{���e��Z�z��Ҵt�qߍ�����~���|BP$�I����ۅs���Z)wm�	-~YW���QA(�wW�Ev�w���������N �#�Jp����M���7��X��.�Z�N��hܹ�9�j��Oz�2���-�"H�����f�O�O�x\�_D��e�~PW�|�Z��-G��nqؒ����ɢ7�I���IP��Q$v�cf\��#��)*��a�	��)K+!���{4>�A�?�' D=�1��ݓ@�7�H!(�A))�A�)(uϭ+�\E�E�Oc~.dw�:���
W����|(U4X����QJ$�
(�x$�蘈�1�0�\@��]���"yӍ��h9�����d��(���"JJ~��HO#��k�4jq�F��=	��ݮjo�˶\L}eFs�Ѡyʸ�Ǎ�|�W۽fm���$��,�5}���V9�·���a�{`I8�$|RS�)«���C" GD��4J�S��-4F�we�{�y{zb���m��*��o����i�(8��9�jh�V^���x���#�j~ĤH]��ӗk�k8�#Dp=�4M׻�1�뛩�be(x۹&���+�V��J���-t�vA�X���&!�x��������X���"F�&ݓxD�C(w�Y���B�Q$�2A	*R�!H9S�}�)�����ײ�Vt��[���0�q�$8��Jp��$��s幽[>}N���
���-����Ɨ�]'`�l:��=�c�i�]Q�V��g�NG}���e�2������v$c�ק�2�Q0��N��TR(���P��O��Q�%?% E!A���,��E����		��ft������;�@ �d�!t	��Rͮ���fw�t(�D�Ǌ?HIP��Q ��ErŪ//�[��3�V��P0�hA�P\�y,y�^�y�.'&{ףP�)/�v����$�T�$�U�]�T��I=�}��>�T��P�k�g���;�����S;V'9�My�-<���l��8�����D��x�Κ�Lg:1��U�A�&�]O�O���%AKL�-iVO����9G5
#��.�=Vx�Uf��xT�x�5w"ܻ;��iE���n��Z�2䦰mel0q�s$��q+��V�Yt!�@ө{w �i�잝��y��dSe�\�-��������3
&��i�{���Z�u�����G#�d�|����a�;��s�*77��N�c��U�n�B �GGj����2�qq��{DSy�J�c��"1��V1d���-K(Վ�r���N��ۮެ�`Ѣ\����k��.9n0�u��$�iB�����s��|)vv+c\�B�ˍ�c��M�;:Wx��5�;p�ծ�]Ѯ_kȦe\D�=��V�Nr�it��׏���NP=쭥.ޔ���������Ԕ�?%?H%%4E2B�$�B̫�^���nV"��X�On`���@���R�������FD�W�(��� �JJhR���Up��9��C��2�e�Όk��t�ٓ_��~Jg�T(�H�ӕ��;0UΪ�Q ��[B�(�HJ&��l��ncp�<�P0�������43%ge)���M C�~JD�IMR�'丱p�;�\s���!8۲�]^���r��o*����\Fo�Ѩ�dD��͡��#�������5�b�p�R%W]2Km�ʪ��v �v���+m�9������'�+�H%4A%"B�X�Κ�]O݀�U�v�I!���I�_�
�ud2�Ғ�@�?Q����J�L��k��&]��Zn��4�J��=/VX�z�/�k@�O�f�ܣj=� /�Xʸ2����P]t���͉��aj/��}B�%���c]fS���2�����G���JZ�ʎ�B�˧ݓC~�"AT����H!~��ʚ��nK�ѣ|�zǚ��r51�gb8�� �u
)D�Ag�U��wU�ؘE"AĦ� ���Mn#���F5��\ �fM|FF-`l����6đǤG��E�H%dRU�PD�d�F>߉�ß5����:�b�@�����$���_c�w%Nh���V�k쳗C+�fD#9pZ��<d��;��j����=��
랪��_öz���\�"�Ғ�B�l_5Yu�7{f:��G��6�j�O(��F�H�yG�QF@!%T	J�F�b�^taS�EퟫzD��n#���F5��]vd� ��D�B*mu)��$�^;_l:�@�D�Ŗg�
J��H?"�����䷃��J���TuRko-N�ʺ0��@��i:�y���,̓��{�\a)���:ΡD���N�'��7WYڹ䕫q`�v11@��@�^��
Jk��$"��fh���]N�F���Y�RT*�l_5Yu�7{g��v#� �(�sВ+OG\Ō ��Y�%�P%(AP��)�:�j��KѶ����1:j�1��ƻh�=�4B�EH��IP�8Wv��Ԑ������T��s<S��eh�Tn%����q��ڈ��
߯��A���B�"��(�A(�y��;���;���/�_Xׯ��v4Gtm��!�"G�.���!0))��|r�Kv�i�Azc�ϨP���VV����騝��A��F@ ����QM���8vE�Q��5�P%8����%"ѝ�Z��ua��U��t���i��OfMWH�R#�T(�~#5�X��	�#'J��/6��H �QFF=��K5��v1p�e��/`Iչ�O8�^a�:���i1��+�����v�j��+>Eq�������U��!-8�^�b����=dq�sD�$��H ���!)BQ���4�ԍφ��S-V�n+�9���|(��Q�;���(��ܶ8�ξ{��;~�����Ň:�k���:eژ�-��v��r:�b��U|��J��\� ������-��s��}R�T���g��To�w}���Ќ�Ybs��,��q��If�ˉ*�N�á�n���zf�ׂw
Ӌ�/���~}?IIH��/Y����D�r$�q��wT�)����n�S��?qm�Sq\A��~8n�@V�����Hn�P}$YV|�1O�̸�����jl��|���T��O1�o����]}�)��}�$���l��U�&4���52�9����_���Ic�ݴ���7�i���=�.3�Q��Ќ̱����5�W)��Vn
�Y�E��,�v�L�B���=���=�vR�'.̏R�n�[��sP̖ @��]�ul�L\E��$���DV��(c������.�C�V^�{d�"�&��V�B1xx)�Ua)jj`��a0lhv�tY��Ȳ�f�Y��i`݃�`�аk����0�\uF�2vN7� �z�iRcc�݁�+��Qĳ��\�f���,n:|�����6̤��b�F�z��D��a,���kOXIQ�]X��g-cd�J�M�8@�O~�u
�`�[��W�,�V��y�	Ey��!���y�;#��Z�"�}���|�O���wdP����U�h����LN�q	�=\L:ǽ3WU��O�}�k4j=�X�33>4.e�֝��%R� �R$6���T��O=.o�G˚��#hMpn*��[�O{WƑ���C�V#ǝ�]_;���Lo]w^�z1LP2��/`I�����2�f'�f��;�j��D�.�B7v��A�ں����S3�A#�U���:������b"y���s2��>:D��b]i�X���B�v�N��n���_���ow��Qc2�&fj7��w�uϯ>���q�@L�PŶ�C.��E���n�h\ۇn5�Ķ	��1���_�	�w���H ��-^v�+ׂn�!���/Ǝ�����[�_Q���P9̽��[�D��#2�N}m���`�_�h�+�Z�nܦ=�uh���F`O�j�p��s;���+y��a��|�������F^hz�Wk�/t�84B�����P�.��s7:7v�]D��q�?
~��	
��RS�it��r����B�Q���2��NUj������y�=�{8}~�v����}�ޑ3�[2�B7v������YD3�st(�D�H����r�x&�B�X2�P �5t+�_q��c89I�|so����}ƅ	%�
�Տ�=���v�=wOŮi�xfg��ګ���E8Љ��S2�#���}���i�>P���m��y+nW �O$�-f��v�}�I����㖔9�����۷��'����@�7dOr�F$mR�<��_|j���5h�'N۫q��&V	�pF&4���e%x�Ǯ����K#�}u��y^�w�\,}�^���'��wvV�[)��l@�"A�����˫��'�$Ͼ��R�޺���
�!2�3�������vY�����n�eqte��{JcǺF��ݧ�N\gRK0�歕q�+ݽ64��,%q�YCDB��J�^�d��l�}9S����D*�,n�tߧ��MՑ6���N���竪�2Svx�� RO_eޝ�E"x��amdz�;�\�[#��xk��(}��y���%�
+Q����.��-�x�;3RU(���	����%.=�n���N�Yw�v�Ʉ\�bQ3!ә��z%�h�a�Se@.���yA/�%�	��G%��vj�g&
: {3W(d2�w`�[J�w$7�K
���Е���԰����Vѻe�ά\�nqc} �M`X�p�V�2����&�..�(1�PW�o
Xgf*dL��'e{I��X�{m<�u�<��F����F=���\{�`��18Js�D��������.��Q2�%ۅ�G�cR������u��]�e��A��>m�[�n���4���A����!@�8�ʝ�I�j���_k�x�Co/=ۜ�
�Z-j�E��w�|�9`���7.l9r�m]�Sv�()���̎��&��_����K�O[��Cu9��#X$����u#������S;�Q6t��B�ݢ�5�le̡�I����nS˵%�x��Ƿ����4�}A�Br\u�hN��՜y�v��z�́��LGY��5��Y|1J}�ӧ�ē��Hi�D*�N�l����jeh�e��n����[Z*l�LWT(|�q�縊
]cs���������R�R�%	H��)�YN�sL�9�	��M-u��3�R<��f�*���5Ӭ�.�g����*cHa%[��Z�KkX�+��̮Q�iVv�u��X����8�T殀��f�l`�lt�X�vv^�m�̭a���J���q�8�Gg8:��Qj66Z���f�3�]SH�ɒ�,�w�Y����q�R(�ΐډ�r�a.*	c��ΰ�NZeʵZ�U֖�ꙴ�c�mWMc&;��t�LÌ�1��,�3%��Z�J��K363Ya�T�a����C8Z��uC��j�#3�2L�i�T����6�Z���8�:�3ek��NvV���YKZҕ���y�\oz�*�'{��ð���ʚ��M3���31��궩����.p���r�֡��j�H*ٚ����'X�es�s���I�M�h�.s3���Z�M-1��lcL�*�z��*��33��ڭP4�ˢ���I��KځHX��
�~�>H,>�)���hB�
A^T
@���Ü���AHo����]s�?S�o���_�������z�RAK@���3�d���!�Q��ÿ���Vf���}�޷�m �P~ai%��e�L����{�sy�z�?n�{�O�CIyP.]RJ�{����9�-4 RAe�����) ��s�����)���o�{�q��?}��Ad�2���=��_��|^�����i�k��䂐P=�- �RAj�\
H)`�L9�\4ϙ) �Q�Q~S�9^��f�O1�ߨV��du��
��UsQg�5V�%�9)�T٫ֿC�A_�8��
Aa�v�O�I�?Y����i �*ˢ
A���r��A~7}��s�^����U��4�ˢ�� RAg5�/;����k�w�ɵ�@�<	) ���i ������W��-) ��9a���RT9E�Q
G���4������1�>��?J�`2RAB��4�Xk��;¬���}~�J���х���0��p�'̤��\�f�Q�������oߛ���/��eB����`R��B$P�KʁH\II�9ˆ����Qi4!I �* o����;��￫5��z�7���i�k��䂐��=�- �RAj�\
H)hÜ��L���
!�Q���Q�$��������7�=u�Z�U��O�����M$�@��
A��9ˇ��w��g=W�ᙞ��Z�H�-? RAeFJ^�
H$|	���-zP�%�v�4�lTׄON+P�[�m͊�+�h�1��oy.6����C�Cv����n�x��v���Bh��{U���q��*�G���� g�-&��Y(e=`R�$�,>�
B���(����RAx����Xs��i�	�}|���̞ȷ�� G�>�	�V��2�����x`{{��� ���L`P��3,�����|7�������ߵ��K�����L�nND�y5qf����:6uU���U]�`|���i�I���HYRAaG=�C���9�-&����^0)��������e��so?����?G䂐���]w,�{��E��
H-~��R�
a�~�i �>�(�Aa��-�����.d�e$}e��fWw^��A`|$��
Aa���I�����9�^����U��4�ˢ��$S%=`R$����C䂐P9�-%W��>H,��z��JH,;��|�!U@g(���R���
Aa�r�n2RA@�(���$Y�~;�Y]Y�-�Tڋ����m ����R���L�A��P(��4�Xi �`]� ��9p�A~`R9E����z��?<��[�
H)����I�F��Qi4�$Je<`RϷ����{��װ��~?H,+�\4�R���(�����]�y����o~r��) ��
a�~�i�A��
!��H,40����- ��
a�r�O�RA@��,�A`i���]�3���z�������B��������ß���s3��}���@��i��(d��
B�RAaF{���AH(�����L��
@�߱��mC��~�s�Vm���&h6kةyM��EWdŗWcr�8��	uk�[Y��A�թVGg0��uٞ:��+�l���w��C� 7�y@Y���<����5s ����ь4�],fJ��\틅�i����E��5��]c�˻k�u�3lh��#m[�������Kv-&���K<�M)[��g�7m,7���.B�RJ�պ53՗sL����P�81݋�q�
��\e���d��[��#��Ȑ=�X��6��Κf$"tXҴ��Һ�g�����m��U�M*��: �볖�B���T�n�Y�G-�W%S�=������?$�U��ZAH)ԯ\
H)hÜ��L���
�D|	�W�sh
�ܢ�}��G�[����
Mo՜��~���p4����L�RA@�|�I���A^T.�)��.$���Qi��YC%/*!bJH,5�}��Nkٚ2�uY�zH,0aH�ZMD) �P�^T
@����y����~�m����}���!U@{�ZAH)T
H)�0�9p�/����~��[�H(n!�Ѥ��Q�$�@���Ц�~�i�ᔐP+��I ��@�� ��.G���"�qi9������:�+��2�� RAeFJ^�
B�%$g�j$
@�(��B�
A^T
@�) ��9a��AHUiy���^^^���H;(�$�������L7�\4ϣ%$)(G����͠h*�r���8>�a
���RTB�~�\4���H(fo~yZ;����j��I���
�P,� ��{�����Qi �C%/*!bJH,*�5��
@�(��}����Ԃɱ��P)�k;����l�}�w_��1 ���a�?$�U�QiTB�E~��R�
a�r�}) �@�9F��>���_n���e(Ny);��N7�;]u�.�.�673��1Ǭ��i�S�д���20����)��ˆ�
A@�ݳI���
�\� �
�9ˇ��w�oW�Y��=�٪��@ˢ��$]y��޾oz����@�:��
���|�R
�E��!I������q) ��9a��AHUP��R
Aj��A���s��Tjp9##��eL�,f��W�����1L�7���ռ4�"�oo�5j�m]���z�fW�����{�����ڟ%~�I? S~�p�>) �~��X{���c�~�+y���>��
�ᅤ���r�O���P+���A`j4�W��������t��XW��4�R
�E��) ��J_���%$s��>H,>�)���hB�%|~�T|�>Uu��-3���Q�H,+�X~~H)ܢ���$�������L9�\4φJH(��Xi�$�@�������;ކ�{[�i�l���\�4�Xi ���RT9�\>H/������k1�g���u��2���I�){P)RAa��Og��~9�z��)2�I�
H,��^T
@���Ù���
B�P��tQ
H-J������L9�\4��|}���~�˼�ɴ���Qi�y���U�������>��
���R���L����G�٤����A^T.�)�9ˆ������������i�Z���)��.����8Q�b�C>�Se�&�\-�ecu�ޓ��~��O��YL��P)II�O{�����)���
Ad�e/* w��}]���2<�#�O�;$d|	V��/P�1X���.�	�_�$��o��i�2RAB��(�Aa��$���RRÜ��L����������{�����g���$�@���nT9�?#�M����a�n�;�Y�|l��
H,�J^�
B���
�ߵ��� s�ZO�N�㷃_��� �xe.� ZRAa�|�i �>*���- �RAh+��
X�L9�\4ϙ) �s�ZAe�tǯ��;���\Մ�)�� ����+��,���7��oi^]�_�^yw>�v����f|e��f�FO*J�&lΉ���}�˥�NԶ��y�W����ai%Ss�2|�H(~�H) �*к H���J~~6R�\Ho���zm���@�D�H�ERމ�z)�Xc��^uq��G��x�VLkn�4��:]_��>�Z$��<�>]E߻�~��M����H����ޡZ>/���6$@#N����˽��t�6JR.B�^����<ki���݌+���0��oMmV�5�ԫݘ?v��C���s,���S�<�^�{1G@v��|���ҝGܲ�2����4�U����o|���y5�m��C0"i5��V�Xk����(t5b���ޒ�Z�<F�S�e��Oy����[2������V��|^�Sb�����39��A�B���PRL�݇!�3yy�J(h������"{{V�S�<�^�q�I��/>�!�wy@w�HˑWf<oo�֢��q]'�sU]�P����_`�%pʘ�ɔ �� շ�+|_�	�~g��vϜʴ1���_��T�b, �no��K�Z�a׺�{���,F>J�f^�fP�~��+�{��G�>�)\<g=K���6^Nsg۞+m�]��f��t.Z2��؟$>}��C���}Ƥ�^�tF�b�K���g�T
=3�Fc�e|A}B�)ĐA`��@��N�W�ފ�$ݚ��Hz�59Sڢ��xo���٢)~����tG^(�%B�� i�I2��!�*�A~�9��o&���VG�6p�8�'�?n��n��h@�J�z�s`a��[w��^q��$�Y������P\�w��Pz�->��*��Y�߶p}ڴbu�L�֦e�8�ݔ*ԅ�2�u��MNT���Ȼ5���{�z����
�fj{�}�st�s�+�\̙{��e�F%C'��j�i3{⑖������7�[�硇�b2�=���83��,���29lh�7,�y,�z�8}���ꯩO�b�~C�Jv �^���d���c�b0a�6��e�2��+vt�%e�)�0�P�s��۟G��8^Ѻ��-�ˌ��ø��1�c٢D��iIe�e��i\�S>ظ�l��=D��]�mvRR�36T�b5in`)f��*2W#���$��mk�n��!�2in"*F��
�;��˺LIϘ�Wh�lqhJ�u%����=�>�k3� d�\iZZXƜ)=8^��;����n�+`�5�mv_��'����0����>�W��K�Z�a�gy�P�4x�����u�~��fs��fQc2���٢;v�E�ґ�(G�f*Vv����#ޡa�P�+G���X$;e���1َ��O�N�5;�-�̽ ��vOS��]+�W�ML�ɮh�5����y��Gܸf�!��4�U��o~�7`�{B�ؒ	`Eu�1ӁּVk��^uq����n�]d����DC���1��Dfe�3;�Os��|����q۩T�Jؠ�>��� �u
��ĐHӒz�殞�t�NdOt��ц�լ���:�.=t-c�l� ���M����E�kV�?�����|�f!����� �Ȑ��jgz�*�����9l����~��ц�e��T�˙��bcT+�8���U�ա[%5~>Һ�d:)*�����T�-�S�"�6�f�Sn֋�l
�Aj�����;�K7FhG�d��M¨����o�X⓺
a�|>��[C�����E;�cӌּXk��^H�8�~�٭Q��7�s"Fe#�e�G2�Li��g���;�{�+=�	j�� �}C�E�{+>�PUI.��5}�)էpMJ0�j�5?V���D��unU.
�G��h��ģyM��L��F�yP���O���>���gp�g�`�_?h:뢶ݡ\͂�q�����@�� �r�����X��Ao,}���FN1�<]u��<携{sחM&�ZZuy�ig��<����b�#�%�P��O��urR^�3�O}����n��rҁ>̳@��b1Ĥ�.�����6�Ii���vm�|*CR��jgz�*�X���k�)�S{�O s��ϧ�G�H,� �ݯ�,}rxl�ݵ�i��*�W-�
�h�vۡ:\�I��Wj9���Cz[n����\B�@K�}R�̠��ow���w��w���S�f�����X� | s��/�Mm���q`ۑ� ���K�!��x,ò� �u𩦮	�Vfh�������e�}�-;�Fq(O���V^��.o�ѡ�*�z�&fjhG2�FeJs2�⹾��u>��~�}���ޭʧ�C(��S_~ޑ$i���I�5�_��1��T#��e�4+)�ݲvyL=v�����C L�G`h��ۖR��n�w^���JD�wF��WK�}�b�t֪����6�P�#bs-��i���OT��9zG2˂c(s2�&��֍t���"W�p#�Q�Vio�|:۱%%� a>���4(O{+�l�ov��?1R%�Y��Qh�Js2�3,�j���������I�53���I�X���^��z��L�Ѩ�U��wF��z� ��_蟈'H���5*��T��ݺ��>�V6����j���;�駗�#�ΕAT��c��ʔ��؆j�(����z��A݆]O�G�+�9��z�>�k��$�@������a�|A;�4݀4�}KÁ����ɑ�rJ�77�ә't]�&6 #�{�Q݉��t�.��P�ݳz�9 ��C#�Mp8�r�DKSvȅ�9W����3�d�5�ԯksS���Nԧ3/BfQa�g6����|
b�"�c��N����g�5�Yi�a��49�c1(��W���m��ۉ �Y&]���Sծqwkw����ǻ��>�C��}[yώB���mǜ��#3,�Ƙ��Ce������K�/vo�m+V/x��ᢈ�g}��[F8�f|=���Y���lFe}1�F����@�F���>1��|A)d�lQ�<q�ՆC0ۻ"��X� ��$Ϥ1e��c���h��3�F��<\�&�Y/ 	 n��K���>F�z��W��g���d�g`�OH�Q���y�8n��D52��j�)��gF�2�/S���mR�MMCs�^��{�:Wٛ�m(�ޅ��L����13�ܨO��zuZ<m�فe��֋�y�"T%�;7���Z�Ӯ�T-,Jm���sS�������5�ιV��M7��Q2���7��9��HYV78T�ʩ{v��b\Xvn4>�Fc���t"�9�í��Y��+u��Ef��-W�r
n��ak�ry,xq��X�҂ �a]�V��|󰑴1k�����T����J7�'p��|�X�����7:h�&=���gK{&P#e;��-Ր��,ǽ��Z���%:�Ab����z�Lêm����4����5��Bۘ��R
Y�j�$N8�t�e궮"�z���ڳ�g���f(!��Ȣ�Զd�'T��:F�j"��[�r͜�xC�1�Ε!4��W�
cE8�,���[+!N�ڵ�7c�)Y�gǫ+&���򛼡j9���RA��c���\�k`	Rl�s
���z�s���υ>��7�$^�j2O>Տ�T�;{�ݍnl��Vp������޳�q�:�ͭ�g&_A��J�Y/i̔V�#�-���6��eݒ7OE�x��S�A]�o��zma���j��0	��W�i�1�HX��[��+Hy��VN��a�5Zy�TY�Ԡ+f'O���adjP�+	�i��e:�c���ZjT�X��*�z��繷��
N�^v
.Ӽd**`�+QT���qZ�H�!����5�C�Ҵ�c%���u�idi����`y�88�1͛9Vq�Y����FWk�g%������U6�Y��^{85N�6�i�k�s5Y<��t�;6flj���b4�K��
���3�Ι�7qS�꣤��sY8޽�ަ���a�Ti,�Y����cu���U��"�ia,���f��lq�OX���f�d�o[O-o-�6o,��F3��q��;a�ٛ�[�{=1Jd��9(ɳ;���sM��yf^��bc�����<�{Y��h���z��I6�y6{X�C���� y1��c���{������35�[���N�w�8�q4m��$�v#;��=^pM�n�-��9�����&f�<���鬚uX�%4<�{� 5��{b�Yhͬ���B0�iJ�VɄLJ�r�{B8g�����H��p��g�{YSM!O	Gsti�&e6�,�d���0:��ؓ�<�\�8
�������b1������K�q+F��_�e������;J��!vC�qڂ+�����i8�x��@��m�ok;��Ƞ�Dz��P�ϰx��t�cr
+d�/������m��9��]���=�l"b�A�Xٴ��q�<��;�n]��<��=e�5�(�;U6��qE0�)+�E5��n�t`ܭ����v	�-�K��Z�%#�չ�H��l�,7Rx��;,�]�����=�.]�̻u��<<B�p��v��/��M�n��Ȇ�[��;ca�\�1a.��yk�p�T쫔��q�q�<)���:��ؙ��ŎL���A4�s��k)mb!�]E��!���3t%�mE1��z����B\�(�nرα�A�ı!nvt�ƅ���(seɗ���<�C����s�N }�6�ܘ�W��A�-+YK5ШA`�v��cS�B�a(k-�-�F�/:�wYP�=f�K�n����Q�=��<�0pb�]����v�!r�!� %rq;-�l���.]%�f̀:�i�a�˳�����N�L�En�n�e���-I�GIt9A�󓵎Y`��u�S�����MRlL����Y��J�F�^>�o�!�ײ�C\#�V퓰�7b{'/a�,n��Y�hsU��q�n:L�g�d%��<3C���8{�g\q�F�yق��:j�L�v��//dʯ]���tef��Ƭt���ևt�W [���D�{��tTE�;l��%�GY�#��$8��[�W��ڠs�g��q��u��9�����`�ֻ@�PHe��M@h�;k(��.:��%fU��{v� �K�Ð�g�n��4�n�\%�.��[0.Yh�^�F{N�na��vY�g�M��7j�a%�����wwN�om|ʅ�-)�R�;��vy@[��7r��a6�����ݏ��nu��)-� �$���8�����ܥ��ñԔ�O8}<<��q�H�0��R�N퇷=a5���(3E��3,���� ���u+��7�T,�f�.:ԃ*��n(@m�3�n�2t��Ƭ�H���釙Y��8�i%�b}�`�ns�AZ[s����B}�M� �D�cbd.�.�6�l�@BjU��9]�A���\]���~�c�r�&�E����5﷭�%v�������>8�^gY�Ш(v�+C���&fkBe���.^#�U�;�x%��A	H�]i����|1��~-���7�0�앬�_Ъ�Q݉��I.�Ho���6��=���L4���E��6
�^@��#�ݛ9�\Li,>��>��k/��ݲ��4>�]gؽ���{V/x��P(�EՎ4�+�}�)D�ǈ�7v��	 ��7vp��튞u�P�
Y{�J3��}<GS�*�w�'��TRK���Vy��WF0��ZiK�tn�Y�G����X9x8W�g�6T �����������B��}'H�2���Ѿ���d�)�����Cz5gS��4�����yB�ݑ �?A�٢2��ִ�K�z�t��RӓjX�������1�c�RQ%+���9R�C�܃
�x�7E���vJT�ʌ�Up^����A���>��JF�2{��j}���d�᯿you^#���Qݎ��J4d#P�	H�BJ�q@� n��vBa�R��9�7��j����{��6S�y�z����Ɔ&fh�s*�xƸwVxt�5�h�� �"a[EM龥��d�+;����Z�U��6W�,{���,��� ���[�'�4܊�}Aj�3�ꡔ��F��+xk}���3�B&w�49�q��ّ�T<�zd��A�" ML�Ѯj�=qI�d����f�Xx�7�Ů
nx�:��%����_P �Hg�wf��$T����˙Ǉ� �#)Y
�o����i���@�34i̩c�C�kw��6���KT �� �Y&z�*m�Qy͜�gP �$��@�=90���{��DƄG=��fe�:c33F��<IOLv�N�>R
Ó�k�x��P��7{Vìf�z|]ʈYR�3�TG=�=x[�v=�r�/wF��{Kuf�3f��U'���}�ܯy|bp,�[���U�F<JG;�ʰDq)7v��=�ّ�k�|�/���6;�'�ң|��q���<~[�@�	�޿}g��e�
lbg�ѧm�҄w�У�x.3 W��2{u�6��(���uzo�����3/�e�&��j�����翗�R�k�D�]6��x����Ȥ�D�\�[��.-���$p�,�z�����}ـ� @��.�g�����q3�C}�yi]�l�ZDWd��0��`��(w`O��[L��sIQ;� �Ț����_,��xx1G�٢���ָW�9.o�ѡ�U�eff�9�$4�������vdu�aɾ6�Fc�wW����{�Z#�3/Q2ˌ�53k��d���Oה(}O�V>�~L�K���|̬~�	�*+��v�9�<����;��9�u�X�cR��Y�4i� �7�0�[C�2fPD�\ó:5�Uq�!;2�������R/��RV�u�����| �}��3,�s(,ff^:�_�������Y�I:5�2��/��-������}��X^�e���B=�(�����=�N���V�;=0Du�,ui4*˳[�r;G���@�0!�c�#L	����F��gky@��Bb�4�]D��~� �9�@�K���&��Ix+m'�7�3kC�o'�c�;r�/c��������>�B�@@ �}B�;�ί�m�j��4��X�K�V(P���Id�C<�pݱ:�pa^\����||h��T�C��I2��6$��XQue�!��"�P�q$1�ʶ�+Wk'����^�@/`{�&�J٫ClYSS@�� ��wf� �Ȑ~ط�9���ڨW_Vc ��̩���c'�P�>��$?]
�j��%Y��Z�߆���J�nu%5X]�w.���-*z�h����蝏)�n�/�lmYS:9;�a*�k�T+ч��|��T>ߕ�y���ӻ�����֤3M����s��m��!�q�slpz���;�2�� ]vQ���@I��C���\��"8G�w]v�\�(��cu4=��:�R$c�y�e-�	��5,ΉY�N%!7�%&ήnnJ����j�ƶD�V�qV8w)���|��D2�A��!�jۥ�l��lƚ��V6�HكlvN`x9uC�y���B��VݭP���>����KW{f�/��CD\JY��,6�5Ê�n�YQ`��J��M����Q���G2�V���}�s(npb��:�/�8�5�:A�e��4�T�1������[�Qӵ��d���D+�k'�ۊ�^���(��32�ח���WӿQ��"74;�$�#㻴8C�[���8�����Ӿyu���Ƅ���G2��0�ڡB\����m��L@N��vEFv�7ۗ2��/�� ���>���Y��C2����Ne\E1�wv��3�&�m-�K�Q��s7b҇k'�ۚ�^�@-@�� ���Cv~5)oʖۚ�F�LX�L�}@MW�tK�Uv�j97]��qm�y��N��7j�^�=�gϮ�}	�}$�į��֕ʘ��ȏ���:v���;U
��A`�ݯ���	#�*�L']�]6��pZʻ�ݞ�%�ّ��#4r�v��G"�4�-\�:�m��zש}�<��i|;l`v�Q]唱�˩({�/�W�I;�?;���z�5{��u�����t��b��8�ɠ;�$�	�P�e�~��ލ�Ո��D��4�U�&=��������Z�˭���m�P/8
��\g��3/H��,fQF���׮k.__&�~�u/�d�?t����.�����tN��&�#� �0~gQ�n��j���s�bi33F�̢ю%9�=X�:��R�;��ȑ�I34o�Ը;�t�W�N�w����Q���������'��;ɥmqjʄe�F��b�4�ZEf��#f��]���v�������!>����|wbH �1�(����Ft�qR�P����(�ܵ�N�~8D|u����P�f^��E�+wZ�i����sU�^�ƇZVeJ~�	��>�w����Z�_k�VSvpO3=�/9E������3lo>��ڡ�R`g�#�X���e*�6<">�h��B^nR����!P���o�������N�E s4�su�����3[7O�������7d�Տ�?	&}!�k#��|3.pF�wm
�� ��"[�0���Xٹ�P �A�;n.i+�p��.P5��S>?I/	/��{�/��m��$uy,��6�p��J˩O�d���D��F�̫� �󹿵��q����n������<�\�hy F�Ք%5�n�ї�����f�������e��=P�hs2���YOY��u�N�+��$�iN��SŭKT(}���B~L��!��@@1�X���ܴ�:"� wb~ �8�Jx��<�;k7 ��Z�'�?n��׸�F�dH?i
nhwdI�b> n��ӊ�3EB,�ͽ�T؋����̪�Й�Y�̩i�&fh����/��\���C��t��C�,O�j��_d��ty(b��	y��K���m�dA�wk� �n��m���ֱh��x�v[!gJ�6�xwtL����1L@AS{�/gf��¥�\����߂	�p�̪�g53+b11��"�݁Т�UUɯe��ʊ^�1ӈ���Xٹ�P?�	����_wdN�>Ӻ�j��xk;�X��yV37VK���$v���Ώ6l��m�v��M�%H�^��XC���H+�ut>��RL�Gqx��TS�~�"B|ΙI�nj���o[���SbcI��4.�	#��4��)"��ɢ�Ȝ��z/��U�<�1_G@%�M|A�zD��{>���{��{5s�Wby�L�Ѩ�7�B�c��ٿlw���g���w�����=��ByE��Nf^�fe�S�D�����.
k����¤�YX����QN���@~(���k�{}s���s�h�Ɠ35��E�A����=�� n�4:��sc��ܽ_���<�~�Oow5��ٔ��N�����8��]]��J���2���v�Z�U�_B��j�]���N���O8��#D%�J�f�WW"��s0�Z��ϥ*�m?��>|�v�d�0�F�B�QU���gYNE�wnl�\�fe��P5�⍄!�� nu�l�2U����Y��|Ή��.����-�SVjdѝTsm�y���q���t�M��c�Sn�\�k��t��Z݁�{F�݆�q�sn0J�������q�@v�O=L�T�������V�3�m{Y�b��#v�&����e�{�o贮�\0�[t���{r7�r�d�U�N�#�;�!�+���|��BO����{�?1P7�{gm�S�,��Օ��i=9Hjt4�P�h�Cf�
����D���5u��*:�Z��G�?@Z�U\�����O.����k� ���\}m�V.ƞ�(�+�s(P�KDq(s2�"�y����櫙Fg�|S�����>�|~�w�*x�P}�$Ϥ�"5-�/w��
�B���A��0"[�eN.S�zٺ���,ۮ��Gx���s�\fT�̹�ˆsڽ|��L��}�Vz�?6���"B}B� �w���Cb���R�ԁ݋mP_Ï�N9�Z����h������l`]�k��D�V*k�ʷ=�'0���4;�)�׬��ȑ�����FTݱ����'��gr��i�Ql��ѧ2�E1���8g�39�9)ܺ��H������o9B22L�>lC����mNV'֨��Ч=��$�H9��2ٌ8z�f=��y�-�� >��}z<{bH`D��R��ٞJw�r��5��I.^Q�����l�e�3�B�9z��E�*�ff�K����ڜ@��� ���B�V2��ѧ2��Ɠ34h�,ߵ�f]�<D����1f��Y�*n�ൊ��@C���K�<(q���<���L����HlLhD��L��w����������{m9��֌�]���}@��	���<(�%�U%�(��{e1}ghxS�p�03^�l؃�M�"ٰ�BՌau�b�]-���tkK�k%�T��zFo�X�eff�����@u�)�=�"B}B�Z�\��t�)��@�A#L|F��w`Isg�eZA���~�"q���Y�*j�ൊ��=�5�t�6:^UF����P:�Hi�ѧ2�Lwm������5�:/�־����z�.��U񺈪�-Qe�x�rRǑpim;�.�y)tn��m���d��` ��Vg�yy=z-S�m�N��ǂ���3�ZBR�A
`�2�����9ӮH�|Gg(T�+v�$��4i�
)�ݖ�<Φȥ��U$AX����S�Fb�o6�무^���w�w6ŸJм1A�@;dѿ���w6Aٍ�k�s#��Z�:�u���R�ZY��L2�3ٲ,7�!Ɋ���{g%h���q
p��s��h
}:��J�fg&7��c�
��]�$.vi�VF9�t˚�Y�U��+4�U�EC��N�G2p�0N7\7�.�=M��4��(��"��p[[���[���՗Qx�r��σR�5[��iiV���Ff���bw\
�Y2O(ھ�m�{���d�}.�5)�B)j��A,�Jt��>q���ni���,e,��(�+t��ҷ�a�%n���F]�s',��>7��8�eΏ����>�'qX�P�V���/&+V�B���(s��-e�U8�a�S�%M�d�*wn���n�S�?;�&��MPWS�'�V�g��'�g^��ߙP۳qrgr�̐ԃ�սĜwX8>Ԭ�!�ϥ�עөx�2�5lV�w@]5�̉�,K�ihZ��ր�1���'[��Χ�L���up��v8U)�"?,�} {�c oE=�u�	mJ M�B�mP�b}�n�ӟq}���!���:�8�<h�X*&����}��]�ڗfZ�Y�鋔�QT���WW�u��� �?AA$_4yծ;��q[�zw��z�cɲuƘ�9���l�9��1�9�O:c�+��Z��9.s2,����˱�Ķg68f8�0iT��;T�1�k�(l�U�V���f3����Fv����F���m��̓��5���8Ã`ð�8��6��YQ��Y,I�Mk��g1���73ǭ��㶘�`Qs1ͫY�l3c3ls�'R��������z���nfvc�,y�;0sc�֫�a�ĳ�AS�ֳ��9���=B�	�38f�;9�+M��gc�CV�+H�T�-���$'w���{�Fs��qv�}@�R� ��ۻ6A�vE�ʕ9^�z�_5����ܲ�v�D̙V���Z����$'�>��o��u��s�qN����s(�ƍ	%�qY�'u|�c��y���u�����d�.���|F�М�%�6���n�?�i��]aB��F n|x��0n��ֻ��(�E���\������'�������VH$i��)�8���i�X.���g��鯫f_�E�������2ˌʠA�٠Gft�2��[c>?8���СW<� :���!>(T�S�u�	���{�����Ji=��4#�Qc1(K�BK������S�g�`G]G�}�3��x*{{��z�fQQ33F�̫?QL�g�~��Т�H4�]�aNo9]M8��
�(B��(y���1t)fUe]��CH4�ɪ�W�mI/�0��fp� �ۤ�*�ˈc&��+�ۻ�k{��L���~$�$����zG���2����ˆg��o��_�ކ�����B�s1T،͂�A�'�>3���	��+zi��D+<=�[��˗]2hsŕ��g.6��2���h��/E+m�<=��4#�Ql�32��t��\<���P��g�m����h`[���7�-���33F�̫���	��;H����+��O��fJ�S
qpS��ӊ�]�
P$~,����&p�ӽ��e/y�Ўe�̢�fY����XT8�N��$���G'v#� ��СS���$?]
�Щ&g�s��JX�����I�3��"s�p�[=�o���}�1��zNvٗ�Q[�����G2�1���L�>�~�}z�k�z%.���ټ��u�qV��(?D$�*K�3�򞆆/,��G�f��_=��7۩��e�gnr|e�c�+��]+��N�q"�[h��]+�u�ѣ;f�{�>�|>S(!1Nx�Y�G%�j,��w\Ḧ&}�ȗ>j��(�a��"v"K.�����E�jYn��i�6bg6Y
ibk`�ͣ�k,� ǡ�`�V��c���\�is�V��&���.t�Wft��w�GT�\-�͙�����μ�cv�r03t+LZ�m�H�j��Y��'��<��۵� ���ؤ)& a�f�;L��o�_����阵ԥ��yᯖ.�Y�,d*�o4q��`�>	Z�Pj�:����zD�,�c+34W�r�<\Dج�ˠ��p!)k0��Ӏ���M�lC���4 �P_}�����pP�ut���L8�է��������Yc3�������g����z沽kA$�X$?]
�7��w�Kq�+7���O\U�#�(K"��F�Տ�4g��1��~V�K��q��&
�����M���;z�G	��Br��绫��}�D�Q33F�̢ىA�٨v4ÞsqփLȑ��������55�B?{w��g���ED��
�6�q\�v�)BVa,�e�X�U魡��ͮB5�-�93����,�J�U�L?��!# A�
;�$0"Wc����NW<�5a���6�C�[ ~��c� �ȿ�К$�����*��ֱӫ*�{��N�0jYu�'P@�,�/���b���c�7hdo�!t�B*$V+�+����(�HT&��x����D~�}��U�����u
���x�Sb�f�gA݈��� ����e#{���f���WB����IHh`�W��Q@��+ϳZ����55��۹��Yc2�D2L��!���<B*�#���B����@S�"��Nss��Ց5�S��M�>�
�Ԗ?k/H���G�wf���~�q�;K/ 4.�*o0r���t��;� �C]C(HlP��˾���@՞��`��/g�i�Ss4h�ӸN�J^ˎ�ƽm��f�'SW�<�Q`�z�̿�32˟}�+�=�S}Ħ��]��or&���$H?tGۻ"�;�$F�!�N��U9Π�YA��"[�9���ٮ�Ë�@���^�f]����]�O���Y߲��1�ܽfQl�
�fh�8ߗ;����lg�,�0��f���a���Qz����=��I�o>�mR4Z�Ǹ;7���ԷW�M�0䨤�᤽«O� |>�v���f�Y�=�v#���j"{�ѧ2���ff�j�o������p��C}�υHj�I�0�2���OL�] �o�k�;9DWl�,�.���������hәP�H�f�eg+�ee:�-��N�N�w�}����רn���
"Ix(Iu�[��D�e*]�*�`-zͳRnM�Etٰ%`9�!��1��řCl�0�\4(Om����L?
�eg�R��tАy��	��ӳ;6�h��'���Р**I����V�唤k��nU��+���n�'�,����oAg�o�h��~ط�R2j]�ՊC��U�֢334i̫DLN��q�~���(�度rSƪ�8���(A,���t(}%Տ�5�#�o�K�z;ʡC�WC�>2L��)y׻.��<�D��P��c�(�@�랙�������մ�^u.�f����Nސ�yH��qiL��)[����YI���@�j�d���uN���Ң�ĕ)8~�}�� +���V"�j&fkB�Qh��9�o����7�]���O³FŲ^�_q)韫�����gl�eTL��u��0�����Ԭl\�QeA�.΂��݂9ںc���Ձ�]���6h�sk����'��	篬O^����0"Wc��ۮgv5ua�u��N�}�Q�^����L�.3(��f]Y�R��]!�1����hW�kwW�n�����9�^�D}�h�s(���[���v|DƄ�wF�̠��P	%�
IuԽ����vkl�~#�
�����=��ѝ�ٌ�34i̫��)L�W�A��(��_wFH�%�(�]��qWcWVWW�@e��Ng�����e�'�E�ʡs2�#3,�o!5D�	/�yB������5�\ʩ�N4����eX��۬7Ϸ�\�ޔM�x���:�s�P��f��;D��U���M�9�����'l���o�o(���2eN�ʌmKQ\^B�~���I����s[V�G7!����풄y��,�ظk[6Cny+�88���\ZSr���$�%�����:xw[	k��.��go\opm7FN�lh��
2=�t��������4b:��39s�����U��3Nn:�������%V�pWS�q�hN�2:w��)���N(sp��Gl�a
L�T���pw\�ccf�l������M.��4s6������OC��	���h V�a���P̤5���|��O�x��(~K�$��I�1_�{����]���a���_\���??P��s*�1����;r������z<�Z �0"{��G<�P���ʰ⺁l#���%��l�U�a�)�����~���IT�?
�ekJ�f-d�l�{j{-���:�W2��"q�����V�Lh��C0��1y�L\��A4Dښ���I�1_�{�-꿰W��y�S���zk������@�Đ4� ��
;����YX���F��2����ó=�^*�^X��I-|(T�B�=��o�lĭu��˻���ɩMG�������E[l�,��dJ6]	B�(�7sDi{��4AH�~؏�ۻBұ�S�m\�?x		���Ӕ��]1��{+>��hL�ѡ�,M}N�{�j_Dֽ����64T��(��;�����43�Q�6�7��ٓ���$�s������>�yޫ�Џ�VӶ��}�W�}�W�f�@�2�6��}�8E�'��z�~��nf�\79�˪��$2E	&VP�ت�}�s9�؄h�턝w��msՕ`��@��$�?n���$��ff��ɠ�8*�ܿ�"�D���Iu�RU�ٍ��A����h�_z��ٝ��9�9���H ��7vE|w`H?iwvs��2+�\�Z�#nJ�^�W��s^�}��h��q�U��ֽ�>�>�z,>@�E3]����i�!V�V00���ͧi��F1���Ҡ�lS7���	?�B}�_ؒ��0.����[\�eX.�l�[�Uҽ�5P8�l���٢�'����N��|B�����P�Pg��=�VaIW{�D�����|(
�hQ�{�W�v,�:R���M�-��B�D��	.��ipU��ch�zu��SΏw�X��u!��2Iw/)s��E�p��v侽�,Y�e�-��{.���C�5+=�pے�/R8r��g�^�C�;�bP�%���}^�=��gh�2�D��s*q�����u��У�'�	`}	�b'��[\�eX.�}@�V�%����t��ۚ�Yc2�\̽Ds,���y��~�{u/�W}u�)*��1�J�x��ԌN4"o��̭��;�泵��?sޮ���.��.���U���9�cu��2ڼ��.�����.z�c	~��!��^�M�F��e�ȭ3�:\g��}\ k���r�*�,�L��OÏջ�(�Đ4�����jíV � #üD���3�w���u�h^e�G3/0��bӼ��χ��h:�P����}	�I2��ϻ�c���{){�j�`��ʯ"�hG=�L��)�	��ї�[�ak����`Nk�싷�hd�Ε��1W@ �,�Ϭ�pܣ�)x��%�{3U,$d�,!%�CV��N�<!���Y�s�=��wa(��-�}Q�i2+�{��܎[4v��!o}<̪���әV�Li34i͍����8�D# E=P}=��ySK2Ê�@���Ad@;�4Aݐ��@�ԹB�[0�0EQ�0j���3USZ��֐�K���V&k@Ѯ��hJ��X����:�����>}uc�h�$�YV�*�vbm�'�����藩sͭP��V|;MСB��H��$5t*)Kk�l��
Ь��&�#:D���Ce��Q|.��t���&v˃2���_w[˾\k�Ѩ�*��33F�ʸ�Le���&��^�T_��]�ѮSK3���l	 �Y�wf�vD��#�B6���o7P���G�whR�J�ݘ�F�	� �>>��(��z�v�}���S��ύ�E���9�\����,hs"o�a���ۨ�k�MzT׷zD��1��g���z�����B�U�l�i�b��N�#:`�X�b{>��gk6� ˫���pz�L�q�)>�v:�&L�(J[g73%V��e���БW^����Q�*Ƶ�N���8έ�����_R\����pٷ��eMt��7I]܋g���Rv{�u��8룯tF�JAC�w��]:�j�Qv��$гw�`�̌SU-�e��}���7��X�̳�Z�̎�s�����_k��Y�\k	X���ѡ޹+vuY[J�+�����&��'���y��u�ѱQ�)�N�9���JV�irb[6�'���T��bRrI/GX�����3�9;���\�լ���-8/�X�;�əo�魨Z�v�X�o�}D�`r�v���Z���&l�,���n־�?��J�����%�����l�*�+n��:�"��T��'�Vͬ����4yQ���'/-�3J%c���ˎ�`ަe���S���;�`ŋ���ә[:4���ިh�u�� ���Yo�m>l����]�.��6�3�p;ˣJ\����lT����q3X�N�VTJ�xv�-��|OeL�[;�-�Ǥ�;��ť�:k�-�3NҬ���Z�sv���]��-��x��讙yu�%6��H��ne-U�i"5c��ʎ���u��۲�VO���zpAg/�����J�T֪9Yx�6\���Va�ͯc�� ��J�=���C����5��S:����˄W+�T��tW����OYU�A�2�q�ϵv�N
����ͽ0B(�(P���J"Z�P�t�3�ϰ�`���6��>��Z��������L��*�o��f*���E�H
��%�5�Euuj(�`7��[0��uGf6eC*��c�v��q��������t鱧N�t��wQuXlէc�;�R��j�9�9�ի��ic��9�>k;�k7�ז&���k٣�i�,s���΍�c��y;7�ϐKT8w����t�3�15�Vu_<�q6��+k=L�W�y�]�72Θ�WU�w6�a�k��v� t]I�mm�-gy�]f�=i��l�f��������:��g�֫<���{ic�/z�l޺پu�vvg�K�I����{�l���ޗ{��θz�cט�y��	)oY�=�OKmQ��&y,	bh�L�c6vq�Gv
H����*\U�
z��\hb�Z�M�5l�B���,K�K���!����`�g�(����e��� X������4�"�e��ݒ�s&��\����W�ۗ��N�X`�$��k[`�Z7b���Smo![<v��8����#����s���XÍ<�16��g�=���W{3y]Tݒ��	R��F��n�v��گ(&xy��omy�s�!f�y�;s�;�s�ŀ���t91�MrH�K.e;H�����nSU��˪;�FL�G4�O�7is�\H����F]m-���jX.�Q����(�-[q��U�;n�H�-�9��gi���c��#q�X�T��k-�.�D+�&������L��{L$	x4�e�������a�����J�]D�`��ۈ�l�&6������x�v�kk-G��5m�;m�Ÿ�2�&��rы�&*��)�fQ�U�T��s��d{��6N�����2�k�Y���%[`Է�M9����3DĶh.hyLq�u9�+�����+G�:�`�a��	�M^]����p��nXk���6�Cq����o'@t�s>1�vQ��n��ظ��8��� ,�q��Jq@Ѕ'	���ơnS<>�ۮE��`چ�Ʊ�ۀ�:��z��<�.��o]��Qqx�m��71nnn��|�����&�LB�g8�Y��kf �z��{�Ȣ���a���r���nRڇmҹ.�ЖnU۶`{/�7N,u�2��y^�1�N�x�a�v2�qٍg���,����z�cl��H5^�+#�3���8J�]�������[����:��:;k��%�5B�Va��\�쫁Z0l��.*�UnP�#��FC�[��N�}u8�\��z��v�ỔC����}���p�ބhw
i��Y�ְ�[�=;Jk��c�F�A�۱ �I��Ƨ��@�$j�VkQ[j�E_����x��8H��u�����d�; �8�]��K�����W����DѲ� +�y��������s���3r cu��;���p�OQ�Jgb�4��ݞ���z�!r�����UUwV2n9��p\�=֨L�D�����˛,җ@H[HK2�LMPl�:F��+v]�n�cU؉-MtP�� v�r<�>�g���}�l���qX�ֽ��ʃn\�.)U�94��z�K*�s��Qvp�sk�����z,!<���^��4�5m�E=���4�08���K���ýw7�<�v��/�G2�fQC̰��]�v�wYT>f�nV,��}يc7,Ox	�����J���[���:��Ñ6�_>ք��f%9�zD��bz��`��'�p�Q�й�{���\5�ބ�T3U��49�i�}wuV^�GAqP���I4�Rjێ�z)�Bif`q\(��Ff�fDv8�p$�o}����f����9�[3<�u�KUB���4��k"vN�{��F{}r�C���z�^���6n�ז.�`k�F�5�kc���,�-R9@�cYQł4RP�2h����ݟ�i�Q�rž�j���`���C��G�����Iu!�E�=���px�LNc#[�P���\��5�ɱN��GPql��tĹ6��̹�f�h�;���������t��0��t�*�������q������[ކ��f{��tn�䉛1Gs�:�f�=۪��~�.������:�W���nX�� s���C��hF���ggwr��i�Q�s���8e,bo�����s<}¶���O�I2��R_^S���[3AW��+�[ކ��fx}�x�$��8��ᶸ�j�6Me�9�D)z�ֿ�������h��;&�ŸN�����D�{v��K�-%_���nX���Ǘ�;�{��}|����C$��P������I:Oi���b��8e,bo�/9�@dF��ǧ컺���I"�B�O�R�)�¹3�R;n��e����X�1�ճ�m���"�Ӳ���?��˥.M]'/Y��# ��[���̃Y3"M9��cD����I�]���1���2 ށ����vA��W^�Q���?T����k"vN��i�م?t����;�E!�C$���⬖��x�B�vL[un17�gd�S���H�^hze�\Eza���rŌ7L�n-"���V0�
-t��5t�lc-X��"���d}ݲ7`n��s�1OC��X�c7�/�����N��d����I3�%�X�gǻz��ϧ꛻���dLh��t�ڠ5�pv��u�|�~W4�I$_I�<�N�1]�.�������쟆���wg��
��,��&�{��
.�3�+��c�o��Susi���Ե�H�j�YZ�Nq÷LZŸ�))�R3=و��>"vT���8`�h�ދ��kwF�T�ɝ��,�_������zG��UI.�C"��f���w�K�o���^G��ʞ�{馫��!����^4�\�ԡ��ZB:�+��8n�\��طOm�Anb{MW���Fe��uH_�_��'K<%����s#�����yڼ�Ν��%Ԇ�4^�g���PS�t�M'�f���α��o�6~�2M>ͮ��6|��]Hd5RA�N�{�R��Ul�I��#{�P>��R�H����:�fC]�uUH~���b�L��c�Qu���쓀-!f��9>�T�r�?T�K��i�PvC�vxsR���os\�?O%Ӟ�P���c�ܧ��@��Y�s3up��Cg=��u��uEnxU1v�%$Q�u�����iۀŭ0�6���.���{���.�#4K�Ku��+	A]�\��^�'�[���i�
���tQ��^���sXB6;l�=tePr�\�m�X�Z�b�N�Ȕ��[=��t碲�<M�xX�&g������O��r�r�:؝xܫt�f�iu�V�04�k*ᶜ����z��Z��y"CuZ�.6�ó���Pb�a�f��jm)]K�:dL�3)��C�'ߩn�XZ��9C���F�CU]B�[�\�p���Rݝ��O���I�KŉV��%�`ʞ�z�+m�>�&�]{MI$_I���Ũn2m�4�jt�����1�#�y�y�ӌ��z���2z+��x�/���>=2�/6�c��n��sf�%�R%x��v`�ع�����_ر.�%�`ʞ�{�ջ�N׆�5��^G��%����6׺���gg�z>������>����Ƥ�uþ�*h�;��a�9W���۵�!�64��4�z�ɳd��<4V��ĸN]����CR;��Z��w���پ�8�X�Z��3Pnӿ�`n��?q����w���F-���B�G�8�Ù���}~�-���i�n5(�i�a�r��oqzoC=�X��9��aj\�N�u��w��<��@�sWw|y�Ɏ��O�S��}! ���~���t���n�ۻ n���픺k�GU�=�*����#\�wdn��;��.�*�?|� ݇���fhx�Sn����X����˺��5!�IT�A�~�f��1:G���}u�K]{��\���{�P�o���R!��q�������ʻ�	�*��D�En�$�JN��.^v���j��F�ߜ���������rt��3}<�����������!>�_٦��I.C�b��:d!R�/���B������ۻf��6jx���o١��k��T�eI<[X�*�×�~�v������Y���*�p�`)�W�6����d�^����..�V��bH��lę��Rt��[��OD#8�C��ǻZQ[1�����~�C�ݾ��5!�%��B��ϻo����g�3}=KR}^����n�\_f>�UO��&UI.F;4����aK|��9]&�;y.��f��I/朗�Myt�t�-�n�����7y���YS���0%�y�auq�r�Q��F�.0���I���3�&+�*�9&;�~�x�7��J�tWs��Y�[Ƥ?I$[���Q�����ku�d�ޥx��������J��y��ޚ�馤�R@�-�ӥ�N�һ�uu4�پ��]HjCTՠv�8n���U��RK���`n+v�N���t��O6�T�A�Eu���)�� �8��nl�ﳛn��)�q*�:K�|��^��i�傜c;.b��N�y���I��(J���w��uVȻ���o�(�{ۻcv7cwi�^�8"
^�t�J��QY���}��_ӌ�Ou�kP{B�ꣅ=Pozf,�a�T��([���`!�lYi�P�@��V�r�fQ×xmo3U��!�Mҟ��)+u.��[7�j'��(��&�=��F��T��L7�<�9lܬ�ʜ{z�Z븭��:+{��֚��C&���}Q2W����I.L�57���%ù]�׳�Q����Uo����!�IuR���ӱ�x�O@̹}n�Jo��W:i��M�Z�Ӵ?<�g�u�]ƪC�I/�$��P��{��^��mg��
\v%N�'OZ�9n����R옭��av`�:e��d�j���4���\.^��8��:kq�4RP�)St"�[Ħ3�s��q��)y�_��������%��=f��r�ڢ,�_n�g�V��q�Bf낖,at]3fd �]�s�0���[����M���98��ь�[������Wl6�%� -�����ܚУ9���8����1��u��:�u[s��H7,���^�+�$v4��.�qw)�)��J'Sp��Ɍ*D��'gg\�G&�e4������A�.�2���vM4yiĦ]n��v�!�uEt3U�\�|Ӿ��{��ׯ[sO���\N�u�ie-rY�V������$���RyGKF�/���F���^��,��o��y�G͚�5����2�H�n��dےL�'�oj��]�^�{�u�o����w�ER�{���/���|~���Hj���6{�q+ۮS��?h��ݷ��G���!�IuRec�����c��i�����$�����o��͟��1���4�m���v�hXz�Y���l"�-WT���i���"�|,<���0j�"jdP�5Nx���wwn��t�qʖ&{�A��g0N?]v��5$��?#����zW�r�%�/s��z�L^�L�swf�-��g[����hK��t�u�F�ק�n���B�7�%1{1�#���G��vm�H	U{(�3��F�c9�;����	���e�8���q��������%�'��t���M������vo7������Ԓ��CRd��ED�*�ϱI�KK>�Xb�X���^w���;��e{�CRK��}��u����M���f����ܬb[����q�CU$��k>�ٕ���0]��ɭ��\
v��ٹ%o]m���/4��6l�'.�ut5�uR��]s���}�����:Ž�&k���������5!�Iu���s�dR=ˮA�A�}��]լ��oggb����q�ޝ��Yv�J�������}��#u�#�����*�ꑳ ��wZ�43	Z6��NKF�&w)�[���TW���lȊ��psd��#`3�$�5���e���']"]�hhd��z��9���誰A�1l��nыfε�̼4�EXvRvx�|btIlnwqs�n'}Y��(��'B�n��˥�x�V3�|���Pv�t�\�h�n�[�ef�<�f���S���W�V����x��W�֦�gi�s���pÏJ��G�w�]��O�_t��B��B�Wh́��8�L'U��ռ�UT:84���ۍ�Mn��]w3�']���W0k'��&̱FL�=*޸�m�+�g%bV�wV5ڶw<Tb�(6�n�\�j�f��.*���Lf��t�/����Q����8��e��㻬�c4m���; H��� 0��=6G�f��s[��l�b�8U�:���Ͷf�R�b[ʯXcn���'C�C��.rxNa���L����k�g�~��;53�g"Jfw2�TFqYi��'��zM��ᣮ7F��pk���	u���))#�̨��s;m#FR+�n����Fqmx�Ө"j �5	�Я&�����Qmu=��,98�܎jԃZ���*++]`��Uf:js���]���lJ�K�uۯ�D��ެK�.�,d-�iP�;InP;]�{�b��#���N�`��Q��K�VPǸ��̦���-W<m%�RS{�R���vuQ�W2�k�ɹ���&�MW�j�UQB
��R�L��C�� ���]Mp7�X9��9��o]���*�=q3��i���������-�1������:�Ek39�6��g&����޵��osk��׮��v������t �Yd��ks;�j�缻Gw��:�ڮ�/{ޫi�,�Z7�ff3g=Ykyᦍ�{��ʆfoFWz��ϬR�9�hǥ�����z;[�`6q6��;�ޏ[\�敩����y���31�{��F��<����j��Mpٍ�fw������}^F
���� @���V{�x;�}�]c�fp�`ެ�]`�S3fM3z�3�i׽�I��ʶc`�}k3fy����MT��3����V�
�a�5��6�޷��o���17�I&H���}��帥�)�r1i����~���I/�fW��!���{�eT�;�'�\�'��p�"�gzy���̇�%�!�5�����"_O]�٭�5nԹ0�x&{�/{�R������[�.3�1���
��:a�f�{<W�p)�+�r��j��^��T�[�$����.F�4�{�F&�&�FQ#L,�<b�g���>�Ir�?V銋�]��霗�{��\�'��8��vԚ��F�-voՆ�8מ܆�?I.[�ѽ���j\�sx=U���C_8jH����;.��+����R���ѫ'��[�
�}�󿊓�[J��xn&���J��-���-56�U�βR/�KU��tTlfU���N@�c�;C.�7�K(�%Id=cj����F���bj�?�^�~�]H~��$����WA���I�.~��G����oC�g�2K��U�9ۧ�����O�����|E28j��^:�﹝�o����.u�3[����WY��0��9��7��2%��{�1���F����Ovp[����;6��!�%�!����72vJ]�!���pJ�{Oֶ.���N������bQ���e����U$�I핗ꋅ&�������{�'7������E�T���^�0�Q���:�XO�w�8jIif.�ee��Þ���k\U���N[��RK��'�q�SǟR����Փ�z��g�s����$�(�֫��b�,k�q��x�� ��9������JOaRv�\��L=���m��e!ʃ�9:�m��'.��J�7ZdC��| ��Ɂ�1Q���H���۲���b��g��*�j!����i��L��e��̛ƪ��a�6���2닚�W�N�"p�������DM��u͖ �Z99��eq�W#@���)���z�؜�:Z��$u]Iq�\�y��Ȋ[z�6,�`k`j��X�[���q�vw0�����;q�\�il�7
�n�5�����P~z����X�La�	�i
(ARW� �[lf� ���u��v�֚�~u��v�۱��z��k��y���-O+��Yu�a��uR�Ԓ��/�oP�J�'rK2=�Ɠ�w��{��z����]�-|�ےeT���hF�Nw_���Շ�Z����|5��i��5$���w����F��M���z��k��y����|��xh��צ�S��?T���I���d�\�VNv1��=۫Ɠ����=U��t��j��M���=Vǣ�8�cğ��Vƛ�&�E�nў�t<��v	-�y\�ɬ�j�k�z|~�]H~��������:l��uLy�y�{�I��4ka��\�����r���_6�`dF�ܻ�i
�lӁM�X%�K�Hɖ�lc@��ļ�gHn���nCma�x2m��V����β�(wW���K���N��x/_n�qsP?|����$C'�_>���|�k�����Iy%�f�WX�{z覓��9� �(kT�����q���;��B+z��;o�^sVz�j���:l���C�1�}���� ��݀7vI8��Q����e<�Ě��w�:Q��5�6g��K��[/|P���v��B �=�d$U$�UT���-�b�ʖ�-��z�9�e��Zl�1��}w�~����맩.�(��Yfz�{���]^A�Sj�O�%�Hj�>7P�Յ��}<�E�ۯi��(��Ꞩ��l��UNsT�Q�=�Q���ͬ��w��K�CR�wE��0ź��;�B[|���ݦ�B�1�f��! �+āL6�p�7�����g	g�#rwKz8��k���_R��}屗�pQ�v~�� �5S�E!6>
n�{�a�.�:���wf�ml뢚n��A�;�eoiZ=�=y~�U<~|jIT��ԑm�0oӾ�5����یV�:�MpǓ���w[�����y��#q�4�`�B�1���\u�7=�S������ bvk�#L�sk�����z���W��VI�\g�����\��}ӶT�9U�O�ꤒI<���.+�v��t�n�L��`&���y�{�����CD������s���� p7`n��7tq���/�(C���d��/=��u4�!�Iu"��[e�(���W����g���lٞ|��o}>�ԧ���� ��S���J6&P��R��b�"� .m�];G�h3r���{��c��v����؜��?`��.�n���R���G���2yi���?���Ts�{3�X��=�}!���U!�J�']�r�����%u͗ȕq��
r�3R�xҸ\�=��&�9xh�f��k�Ʒ�����y���a�p��u���Э&�t�a��������CUR,��>�+��?l52��y.�͋ϕ��M���W�k��m�u3���e�)@IX�W�'��O�I9��M	��v8n�oHIJQ�J@1N(aTON�RR����Jj�෱s��gZ���H��ƞ�9�/�Ol�� ���;�N��=:0�c�:�)��kV�c�Ӝ�y��)	 �GM�������xW���˄t;ب	�������±��h�O��v��l"0�ܾ�ӚUp^q��[����8�����w��wz��4��#`�F�A�4�@����w%t����cOL�t��.l�Ũ�<����ac).���P�f����"l��1sv��5��ɶG>�nh�U8w4/g��}�m�7�G\<ҡ�Վ8�gd�ݷ1�Noj������q�����vP8s�`ڴ���TYk��j��嶸];��	=��#����E�vx�c�� ?�}��]��e�l�Y���|����WA�4�&f��2f�J�s���������/�BP>IH�k3Ԥ��̮Bk����Y#���m�.��% $��G*��x�\�Wg��c���j��'5JF&(�fJ*E���I%�"����-��J�f���p/}]%����ۻ %�G	]_NT��Uخ��@v��m_�ϫ�J�C��q�v��RRPD�b�gu�=[/��
܈��es/U�p�~�r�|��F�X����7�_�Yz���VҩFݫp:q�Z�<��u ��3S*�������>|�%?% *��=��]&���z�fϢ'i��mֺ�ӵJ􄔥|��n�*o{��K�1 A�h�ٵ6�֡�\�^��.�)[�A�"oj��EE���b�Z����zj���&�,k�)�
rFWDuʁ��<��t~�]�3֤�̮C�*NG��=�	,�#�xO�{ȧ�G�) $������w��h�Ob2۲���s<1��?������I�TGKs4�k���=r���v�[���N�;�o�{���o������@IHIJט7oC7��\����;A�o;k�2�>�OO*���v�i:���	WtMcྻ9ƍ�x`��7ohgB�R�����sn(��M53}���	)$�U��}�o��o%\�9�̧UH�ٖ澰�Ig�F��ȱ���nOc�S6;:���Z�{�7�=��%���󌩣X�۾ǻ�%$��W/6���k���I�+�n��X�jS���yƜ1��k�km��1���Nɴ�Z\u��D탁3��Kz����-|;n�Z���7����9��}��RI+
�uVI�l-����SWg��e���JɞM٥�GL3'�k�	)I$���!5-�0;�G'WѶ֩��r���v~�%!$4�y���]��<l@�$BFN.ݘ��1D�8u�	�E٭ѣ��3�(x
�&��>MHZ����b��]fW!յ'#�L�m��"E���۟��?%	)$��ꛪF�]�<��z~���b3Z�o%dO�䏳ZU����h���H� ���IT"��xzu�<��֎���v�F�w,� �g��RJ@J2�(�
A��4gM:�N~�$��U����{k�2�>�.�Nq�Vsr�;E�
��ݥ�.��;uϕ0�Z�.@��;Z�^<>�v2��:��;�(�I޾�&T��n��� { ��.�~�˼RJG�BJb��*��ݢ��O#bs;�G'��'���3]����t{3 Γ:c30�r��&���.zv��*�h�i�6%��V���+�߾|�z ���I%7.3���Zҷ�Գ|/���e.��N9)�䔥%:������%��ҁ��"��\�r�2�q��;3`�!%1��LCF��X��w�؜��$�$�lc�pݗ�����Zy/"x}o$f��䔤�\4�����RfFnN7?%VS��ǳV���u,��qY�aAȳ�.�CnBI+$�.�����1��z���+�n�o���S���[�u��������T�Py��}Q���Q��hՒ)��Q�-\�t����&����X;9��&�=�M��o��38u�y�.v���H�w�b��@�0���1�53b��s��a��v^޻�*���n���Ȑ6@�[Œ�\Bc�9A����n��f:JF_=��oj1�2�ˊ�w0�<����)��|���1�L���w�{P�-N`�N����x�:٦j�2����}�Gdc�b�!ING4��uڐ{eb���\=�.i)�0���N����p���o��ˠ�ܘ���f�Mބ��(��(�w��=Ѻ�I7%�E�-���}x%՘����v�E7n�ۥ8͗���iĔ�5���m�W|*(;N�J,�����\xᮺ�j�T���!�"��K`�5!e����NO�e�F,�ҥ��|n�+F��a��VE�n�)��Pb����@e]n���ngca�p�=V�.Y3r�a�p�N�#��캾Zv��W	����e˺�GL,Ҽ�1D3�]{Xf+�P]��.͍�vN��E(gJ����9Nt������{M�Ư3fT������(���M�T���T�7�fI�>��L�/�Vܵ�_Z;3�΢Vx+����#��)i�'�Q�(�q�ݤ��*p�b:��3�lJ��CV�y��DN*u�!%�����h�w�f)t(�Щ�˾�Y�0)5X��N��1
�m�<�Y��U�|&_p;��[4�:`"�h1���{ui4%��'�j\#bf����ʳ~L�1��^�2�6�e��޾���|�;Pt���U�O'p���ꊴ�ӳɃg:ҝ�cm�뫮o]gU�s3�ռ����V����fG�gfVlwY�g�֘���Y��޽�������S�5���Fs	fs���S'r�\mS}m*�9��}v��v17��:� t���ڐ��R7���}�g7κ�[0��oi2�z�yo�;Y޹k�0Ա�8ڷ-0uW���5�W���V�˳��˦��p��SV�[{{.a#1��C�{z��1���*�pg������oP�{��U���5�����N���oY92���{�oe卞��R^ 	M�Ę�k�3[�C�Z�f�8������ݎ�;6���U���ͯ���E��ٕI��-kz�W׽��3��Γ�V]'��k�� BYe)>���խ�� GaXem��^�9���`j�׭���!f�3�Y����3��x��0�s6�ȇÀm\�K�z�)���X� �&�YL�6,�x���n�F<\ov�R�8J^D�L���ʁ��vU�ջ�$z�+��Ŵ�6���Bg n�$yM(ˏ��u��SY�\����e|v�SSl����j���u����꧅;��(Z)s�� &f���j����QaWE�n�7��}��=�X�b97\!P�kي$��]�뫃Z8B���ۭh󀭻f��R.�[2K��\��Ɖeؔh1��6F��-4�q`�.�E�Ý���=9�a�X�EqY`�*a�[]/k,e�K���/bj��3�\��Z�Y��y��͠n���% \�ݥRWR[c��^l*$p."�n%�"�q�kv�;��s).8��/��=N��Ë�"��$wcW�{Vִ�H��7rm;��r<xx�=����)����Oru�ţOU��͆'<�6�&EzD��s�]�C���j˄�W��!\��I�/���<�&rq�"푫V�f�k٣4fX�G��aC��w\�Gu��O�AuvK��I��q�`��Vͬ��n�q0B�f�%���s�a2[Y�[�u3�%�c,�A���J;�.*V�GjF�ʘ,�Q��uvSn����t��.�Gt�Kd��7<�1���.h�\�(�����PZ�m�nZc��`�E�P-�Yz��5�l��3�ɹ��Wh�E�%ӣt@c�k�:�=pp�U�P�Ͳ�Ժ&�!�r8��<�P�Xl)�YvLC���3,�E#�cuHgB���)y�ֶԥ� ��v4��Ĺ�Nݖn68�i�;k��wR�8�C;�us�n�%ɨ�ޔC�s)���D��uF�ӭ��r�a/6�'ېF�v��bV)4R�@�M�Ia�楻�����H�m
qpݻ�:@Bװ �y��m��j�L�\d�I�V�a����{U+U]Tn�JpZg�k�9�)��(=[�^t]�+��9�4鮢����D9	������	f!^�^��3�7�b78�hg�K�0����s�=�FWM�^�Z���`�Ԇ[��W�뭼=x��pa�ǎky�:�������N SFi���ItK-�oY�&���;[��[+!4�\V��:�nO<��+��7�3ΆB��7l����K���.qQy��ǀcv�z��v敎�g�P�	�W6��3'���}{��I%�e�����\�'��'��ų\\y�
���}�JBJ~K3��쮵�wH�z����{�O6;uL�-��G�.M�-�Y�NBJR��V��2"������Γ9�ˍ�Q��P���|�$��q�DB���s�R.�8�v�ߴOs�b���|7d����j-�\�򐒟�Q�IO�(d�',�sO.5�n�<�\��3|즒�A���}���|�M��]L���.ѕƚg�����a�5�1&ew�ˮ;7F]�3m�������iXI[��ˍ���9ˍ�������7��������~JJ~�%!��.O���j�B�����2_
��5.#u��T=��G1f���h�X�ֻ7kw'�[��\͘��@�d�>ГT(�C_|�O�-�׶s&�O#����䁚�����_EV���ϒ��Ig�>\f*)M
��y�bԽڧ���wL�|�g��䔄���������N���~m߼~�ݿ�?s�m���f�sx!��O،^n� a�o׹#zR���PJ�ʼ�4�9��l���=�l>����s���Q��-��QZ�\naB������$���-�\h�$�D #%k�$��n���j��S�� m$���Y���j�j��,[��+swr�
p��I+	)IM��{Wݭ'�Y}"�9�S59����*8b��HI\Lio$���`(�]?$Ҵ�JeHB�n��4pWT�1ED��c��{
��=�7}�B�t*y{�1{z��2׭1Ab���]��zNS՗�
��ԝ�Χ�^�����7�p�y8�� $�X+����5r���J�7�gi�S��R5��1�"�e�ӟ�z~J IHIJFՔ;8I�������i�3SyЗ9̢�����������po1W��T�1Թu�+r���bi=#ue�u�p�9۰���a��P�3jjg��~ހ������;s���;s�g��BEl+�0��P��R���x���qsf��n@�V3���v��=)�#<���[�*:�龑�JBP��_X�ɇ;.��jj��m�]����>r���I+#�r̞��rJ�E휹������Ɏ��|]�p;�eM���\�<�qn��̞��g�_�4����,����u�u���{ZY���3���a'񙣤f++�3
���	H�����wm��%%?$�*add��U1it-G�v��=)�)��� 7$�$�޼��ݓ_����~!�n�x4��4 ��3���4�30���su�'0�8k*����9�l�w=蹕&�lc��]Yq�q���'4ā���wO�(IO�)�����u�}]#5�vFn�������Ɏ}?br3���u|�~�r;���������u��u�{'k���O)Lw�n��7% $�.oQ#D�g<϶wr�۬���o-g�n������,�A����{#�p�����$��ݕ[��S���������=�<��Lw�} -r���t��n�32���׵�k3��{!�����i#)�"_ j.<.�����;��HjQ�`����3L��e3fe�_*{��٬��s�S�Z%����`a���a	�aL[k,� �i����{@m�6�9܎ub�"K���+t�����u6�T�PMO/>Wgz�v����^���p��GEֹ���4&��rʴ�M��$-b��睳's��v.�D��%\Mp��:�"������յ ��i�����Yp̰�ue��a�HܫK�`����q(K�0.J�!;�WR\����|���I�:`�:��gVЌ��F�m�`������C�Xfğ�Ͽ���Gغ~IJJ���s:���o+L�u���5��7|s��-s�JR�Sؙr�_T����d��L�˗���ﻯ1��+���	,�kAQ	qwvs�Q�Z����A!�Dd��E��F�pn�����~ZҰI*Wr*]h��������jBP��n�ֶKy[1�ݚ��O� �/-m���	)I$���&������X�=�SSt�.nj��r��󐒑�Fk��̼�<��$X��&�Jg)]���W���YK�Z�vyi�Z��)����>n9�.I_�)0��ۛ�{�9ۜ�����2�W<+MXI$�|�L橞��b9yI3��.x��b�崎���}s�w��z�"���3ےf��׵��w�}bMU/�q���>��L_Ν��Zsp��%J��]�������Ɯ�5��[��<n�nH��|�vΛ�ZW\��srJ~J\iģu|f�8�SMTl��%+���q]�}))JS�S�ws�mM�[
�5&�ջ�\�Q��3�����Lp���>jf����v���u�JBPJBI
��j�M(�(�嵨ӉƔ.����ݟ�������t1#������߾ʙ��u�nm����cK�<�����F3mP��̬�G:����=z�d��E��� �������77\�y9����J���v��G��P��������s����Etp��p�.�
���+ۻJ������9����٢���|q׵1ؗ����}��߶���~!�"�-���nF|88�5�74ɱ�~�?o������ί$<�p�N���L����o�!�M�����e}	���/!��3��'��pZ��lӌ��'/]pQ>))���H�t+��n��@#��.(�9{y<�&~��q?�s��^:�W7]����g����z7�pY��CM��r$۠([s@�܉!�W
+�Ng���g��{B�{a�W5���r�=S�٢��(�A-���=[Ҿ���}��=�C�L�� ��0��9u��YD���<��g�<�����q��l�����ϟ6�[�!�u/�δ�z^��Q>�����8��3���t+�ۡ@�A����?�H�1=�S�B~>�H �}�i���.����V�������C}"�J5�ޣ�~�tk�3dI�E�� ��I���t)�^��*�^��c�4s/���Y��'�����q��[sD6�P�y��#�%����Q~鯈-ȗ�Iz#�u�+��ׂ��⒚#�cv��#�]�:�n�vvl�T7&�Zk9Ex�ø3Qk�bV]>4>[Hy�< 6B/��r�ƮC[�[z+���j쫋CF�̌RH��T�����#�������� ��P-«�.z(Red��y�SVo;%o�������	 �z�۟���Y9�����Q"������uQ�8od��6���ѻ@.���6q-�%h��b��p+���r$۟�6�W�61SG2��.]g�c�����j�g^O˽���0�۟�z+��O��>�U=籵��R���=���o�8�	z1:ࢼ(
[4{�O�6�rF(���}����E(�� �sDۡ@� ��'
�:�U�e���Y�y���x�
���{�B�nhnD�۪X��Z���[,����쯋n�}���AUQ̾�.��1�	�l�������a� 5��Cn~nn�m���ϡ��f]߯��ԍ����vR�N�lT��~�@ψm��۠ۮ�^�CޚFbZ�2vT�8��m��K�W6*r�[�dIyb�ɖ���3Z�(em��w,ݽ��,�_�(r�^��}(=�M�*ɡ��qhYy�Z�d� �]��k!���It��v鿻���)�i���A�ˈR�7 �"F��;�t�����'c�x.���pl�B���&�Y��z�U��<��;Vl	�lN;3r��T���F�M��6U�]����1t�h�Y��F�Kq��؍99�6y�CrK�<��rF���]3Ԥ#`XcjT+�4;��eLg�5E������߸�cC7��Ō8�(�!r�y�X��^�p�V�ڴ֣3E�>���=���|��FĐKn{���Ý�+����r��/dW���@~�@���������5���[423�Ƃ:�?{·������}�]gTǁ�=��~�����S��/Uw�^���tP �O��t(��!��ˆ�����}>E�:�j�+]�l\��~��H�u_6�P��#SF<Z�&�Α��W��ğ�s_{�\9����+�1W���
��^���o�[1p;���܉���P ���Cld��Ti�����n:�x*�7�������<A��hF�P��I���^���Ͳ��O�R$TѨ(Q4I��l��9����i�n�vm4
c.t5���Y]O۝�|�Hk��4AȜ��H�8�
K�V��ؿ
���H
!��^y=r��uȟ�MЯ�mР[� �ۚ#ʭ���g���h�Bb���:�b*C�$8m�K6:W\��ok/s7qw.�D����^��h%�VV�!�՚�d�1��ɭ��d�Y~������k��^^�^q���}@���{�B�-��P<�2$�������4!�mЯ�n������긽��v���u��:ީ����l����[����!�!��ׅ��9�#��Y���� �"s���q���V��ع-��W���1��ȱ�4��5�|_z�|[� �����
 ���`�����ٲ�W��K/uԯ8�\W�V@�;�"�nh���V�׌��ؓ@ə�t�9��r��e�[2�D@*X�U���1z�c2 �������m���nEv�䠪��c���1�BB�߽���s[<�l�/�$ۚ!�U�p$��Ⳟ?-���M�/�}4#�"s�9#��wᱞ�J�5�ޑ$6�i�,��c{�O�q��ޟ��ۡ@����C]��k��;u%�d�&ѺOFS<(�]��1P޵���;\����x+���{�cBɥ4N���������%K�/;��7�ub��1@�<r�]㡎���!�0#���22�Y8� �Yy[;_��[ه/)��I����Q�Î��p��[�����a
��ʄ[b��"WVRr��+-oe
����}kx�M1JK%5ܲ`�u6������e��-4Mj(l=��f���#tr�Au1e˾G�ӌ���!3H��a�٭S+x;�Y���'KZ�|�/�+{�f��=��'j�FQ~Z�yt��Ѵ����������u�V��"jL�/wf��,�ԛ{T����z�g^��[��ewJ�.��XMw<�o�),r���6V��^�.ZN#��$�O/3�'�z��L�3
nс���L1wf�ad���/�#2WV�W)��ֆ=޸CˈjYV�G9ͽ���8�ެ۶��ᦦ#�I�]�n�XfU�l<W-3;x�Q�A���7X��#�[�c(���%P��u����	�T]���ZT�#U����ӡ��on����9�>�yL@�-I��ЬשK"`����=�TӊJĔ��:�F�/rK����+4�r]��h���5�6z`˼�[��=W�%�ה���y�K/�_)�!��{��e��t��ty�O>�B�-=R�}��sOm�vR7E���U�Κ�v>8�&0W+j�̿��>c2�,	�>�+���j��rMU��R�#��Z�Tؙ�46�f�a�cvcTL�cX~|�>�)��XRʅ��iJ�>�a��o��Y�Wd��c�y�z�[Z�f�u�"���o2�'+�P��[�����t�`�Z�ͤ��C��
���1�tM����f��o�G5��o'fi�r�k9�MW6Ke!�n�y����i��s��k��m"�TR��5��������kK��[�o{�7���i�ƸM\�+K�]�IZSh�څҹGz�3z�q�Mi�˵�E[2���M�qse�e�������uٵ�0�M��f���o�&��fjc�Wy�ތ3&�AmhP�,�յ��:dkV���M�{��N�Z�4�5gZ�Y4ƫB̌�Fj霚��k3c;�u�+�1��"�꺧�ښ�U姛��Z]�2�kIft�beY�oVso.3k���mj�U��U��y����v��������E7uud�MQ��`��i�囉�9�3�	YA���nt�	6�
_�����G��?vl�{�B�?6�P���H�
�{�e��c�A�����=�h���}H��!�B�n�Cn����1�z"c�H�/{�q�x+�5z��c<(�M~���W͹[�ģ�=}��k��l�k
���-+��g� zwƜ��Wm�x�-�t�j�W	SG���!��̂��q �nk���3O/uҥ�>��P�}'{$G�O�qVe
>~��I��~-��^��Z�s��f�
��t=�{+LЫy��\���x�w�~��P��qy��UO�P>��o�U�z�ۑ_����e�"�v��g|�5z��c<+�h�;�$۪��"�q$X������3U<E�G�%�<�_����z�Z���~���B���>�����/���0�0ͼH
���`s�gwJ��dO�ޤ�y��1��VT����j-X�qa���j�D���X�� �"~6�P%�4n�Cn�~����/ޡ_?e�R��V�}�\��&<'{g���|�` �[s>�ݓ�:��?E��eE��u�e��i����� `�E��S9�P����r��Y~�>���>��o��1��ϓD7/�[���W�jھ"�f�pb9���"�@�v
��ۡE��-�����W�ʈ�c/�H ��5�%y�i��tM�>z���{�P�H�[sy�wJ������܉k�A�����H6�����.=�&g���ҧB��{�s����l�[����!�#om��{�� Z}B���-ȟ���}<sx^��j�7'+T�"'}:_��T�<�����H �[s@�n�|[��'V�ssC��/yw�1�����5ޠM�~}�m�[�$u�We[�ߡ�U�ҡ��J"{gU���=����ܔ��4�Y'�p�ef�/q�~wjRF�4J�֭�`m) .^4���w���D�Tn�2���ea�6����#-u�R�0XT��#���c�v5e���<˛���nދyƻPr�����I��j�;ָ(cu��l �ҳ7�.�6�f��/r��6��g��2�gGg%����y|X��z��*T�n�16�		8�0r��ݱ�w7F5�N�1����+�������� �u�O�\[�T�X\LX��نpo�!��3���in��*<�V�]�8�lG͛�==r�i:j�¶�x�sD�$���M�˽U�4+�w�˝މ����s#�¨��{B�n m�t>�An�������k��"~����f��X��nO��~+T�w�O�6���^!����w�~��$�'4CnE�I��4+cg};��D�f�;˼���n|w�j�C�H��nh��r6wg�sɠr�b�|��~��I]B�?6�Wff�q4'�yy������s��|pzkgUk��}w��?6����	 ��
�=^�]�@��y�O�;ѭ�o]�U�(����0ۯ�|@mЭL,�|�a�e���kv��	[�S���e�.�v�����u�iV�ָA�y~����a���������V��^]��g���5�'�#�d��M8�`�zE�hCr$�܊-���އ��40R�}d�8�P�M��v�P�Cd\n1ۙ�N�&;m]��3X�/o�cw�8œw;�)F��Պ�s�e�������3=?{�#G�3R�����y���LǾ ���������yu�!9�o1
���~����	mР[sD�Y#�Wu�~�2���aloi�m��S��π ����_6�WŸ�{�[�I�s�D=�P��O�����Kw��e�ъϭ��5ޠM�G�m'�ھ���@��nh�܉6�<�S��}��3��*�;9/7�����A�u
��~mɱ��G����oωcE�d�&˛F�Vm�E�!�e36$v���j&�D̊f��ML1�����{�����2�^��z7��u�|2o�P��>��Y���#\���?O͹[�[s_��T��`�Et.�D�J]4<���w���b�n|t�Y�>��3���<
�� �*���4AȐCn~��v֗rH=�6�D��gdI�쫟��|iO����bc�>wv�	�U�9��Ƹ���)P�n�aU]l��/k�uҬ���@�0V8=�1̻ͮwSM���Lǁ�w�D��� [�?6�!�_
Yڙ���9��]4AnD��}z:=���^����}_4���c���von�t���ߋq �[s@�ӡ@�vw�����g	1�N���yX{B�~����M�/�B�nh�܅t*�8=���GȘD�\�*q�n�kn�+�ڔ�=[��%g��G=�Y��*E	��ﺁ8�4G��s�nF�ٗ�\ULvr�7���"�}<��X��j~�{�����?6����H�}ЫH��X6�~��'0�h��F��=R��e{��h��	 ��ZW4��r�������
+"A��@�t+��}%�%dlKG^ߊU���Q�i��ρ���	 ��O͹�[� ��PK���uB4��#ޑ$/:�m����ۋ������szf>���M�ǚ�n���5QbE��4�'/V(����!����/�Z[[znKa&مu2����c�Y�mh�%ڽc�N�[��e��.��S�P<Cn~m�n!\�����9^�o'����̯
�����+�l}~O�п}�y��)�TB�ʱT����ۈ8�C�<�9��&�qu!����-�G������Ξ �~�[� �ۚ���"�+;D�7�n|_�	�ܣ�o@k�h"��(����m�[s@����i��a�z+����^���W�|����c��?k���W�T��&�	�P'��[t+�[s� ܎[y	���w������O^�fW���4�@�Cn���n�n0�4]vڱ�v$n���s�@��Am�zZ^E����Zo؜��@��H���zwÊ�}�c�A�?H�u�[sD� ��ٞ�P�v7�����B��f꫃R���^��c����~���%�74���W^zW��s���{faް�-b���W�g:��Z�"X�o+��[v�C�D{�b�q�Q�酓���[y���f(2k�!fP�Y3���F�v��v�;����X=�x�ZZ�''d��`�x�&���r�HR�����Sc|��ej��.[�iuca1[
��CU��5cK� Z��T��.�9��1���L3�PZ��˴�n΋H8�[B8��H�ۍnn-.�n �u����Ŭt]*�X	m�ck5�r�R��n��La�.;B��k���=����ז�Z�γ�O��Ӈ�����70p��ۂg[W8)��O_���B~��F>|��NNztu��{�=W��eH���W�=���;�t�#yЯ�r(���4	�7�\j�(���A �9�;Z�.��R~Z���H��6 ���(ܡ�T^9V�
�?��(_9�nD�u_�t2�����%�ź˸N��O������Tǀ �_��_�WŸ�� �����H-q'����� Aʅ'4Cp$d�N��tox����̩�?@ܿc�z}8vt�p��U�~�q �[s@��n���s~v=�{n�f��]��)����o�\��
�6 �ޡE�4A7 ����]�]E�5F�&� G>�R�#`+������/a����rә�m�a{D��1U��~s���������uU����7�[��{v��,�Ӳ�!w�Q�H-����P%�AX)�Kq�Kd��"���G���5�h�yAd�ʲ�u�n�ެN.�s9�(�Vv��Xԏ3�b�﹢G:��
K��r�����/�4~�?d�N�����6��w�^�<��ޑ ���w���F�1�[#�@�p[t(�A-���>�uHY1ڔs7V��ܾ�ס�s(��?~Ѩ=�oH��'{�/w��$ҭ�S����
���
�{�nOe�/=��T��-�h�ݿmB��Dh'�<(�ĐO{����-��Am�͹c6�z�\E,����9/ޣ�~�^Um^7~9����ސy_ۡ��6!���iPr�r��e������MX8n��XP���2ܺVj%�f8b����ֆmCo�<����`�u
��͹�"���9����\�
�u٦�>�E��i��H�BQ�Jp��3S>��X���
��z���qM�����8��� �ߦ��"�n:o����������#J�	��ۡ@�� ��s��w]��7\��:�Sw�u8ܛa���6nMz�X����&�@ǂV�J�x�q2ee����Yb�W9\$�N�G�Ù�S�܎�����xP ���A�m���nE��[ޓk��W�ѵ8A}�(��nk��)�75r���c�����$/w�¨F�M���9��}A��Knh��H!�gL
TxQ_g^P�/s�*{.�{���&>�-�h���n$�[sR){�����ɝ�UF&&�Jl[�H��E��q&响��-�]e�L�2�Vg_�מ��+�$w�B�nhnD��y��|��}W�u�u�-�O�;�A]�s����|Cn��O�nh���w����{��?r�y��Lo����0���
�P��nUy�=�\ZQѯ��U"H�t�ϧ~!�Cn��n�=�N�5�{��b���&'}�[�� ��P��q �[s�o~�G�l^���a1P���Cr'&���V����ׅ����S@�M��F�{<Z9&g=S�\��ݺ�KS�l��&U�XQ��{��֝����EIp��+i3��p�&+*h4w}�~�7��*:�a
R�N*[~Fv�|G.�E��-��r(��Qa��e�3��4&������0�(� ���P��nh@nE"H���l�h!�#D��Tjg�z�Xny��9t�sw]�V8$�%������>O�>���~��"@!�U�nGe��!b���r^�� ����9��A{��q�[s@��W���2���zi�(��A�s�99���羽���S����l�_�H!���@��_ݽB�/�AN~��|�}��熃i9��ۼ��OJ�����a����`��!�m��^̓B���<G��B~����˽�VMM����+{f>�o�_�RXM�/���An~m�Kp$[u�ns�^�n�.��#��^�����0��uᕾ	�S�|� 6��܍���z7u~���~N4����OstĬV�w�u#U3+��>Npu̢�05×vN�����7Gb� �\������NN6�n����%�p⾴Z�����g���ۨ�U��(��oX��sr�Ĳ��a�/fQ�Uz�W@�OkokFu(�k�$;����cHv��e�zn���F��kEm��wFdS��Ua��S��r�`6\��g��@�����=Ӳ��^�\f��VC�l�w��֩]�6���Uv�>;{���xS�
*�ێ`7��7�w���wQcwr>��e������v�{��M�ԧ2��T��6/�j�*ѹ��i�r�r��U�����P�A�t�3�Ù��32qݺټL���ؒ������1�5՚dѻ�kJ6m�IGu��^]`A��*���,*>����:7��T��g��>�9��f�%���FN�oU�7���^���wn�Yj�j�����qS"��:���{��'.�k~OWT4l���X����4�C�.�|��y�$왼A�yR�<OU�*����:wR���qԗ"�����CR�Q��6���*L���deh�륮��������I�]S.�p�3�)8��(6{_MӅ�g2[��0��xo���v�_\�E�t�gGa���4���<��ѕ���/E��P�J����S�kr�/���nK��pu���W:���wV��B�Kٱ���ņ�J���̏GN���!V��1��	�m�ˑ X�f�[�X�#��y�7��N���գ�w��i2�X��e�i6�����r#&�Xγt�mT�8�W�oH�r���,65F驭z��ޱ��fcJ�J�i�f*�d�i´ƫq��L�9�����mmS0�s:��Z��tX�4d�Y����fuk]��.�U�ֲ�'V�d�i���k-o,w��MY�:d�)�UV��0��֏Z��K��=����ՠ�ձg�͞��Z�u{�{�I��b�љ'Mg��+���)K��u�J���Bf�L�7���u�@�N����gy���^Y��4�fa�o,z�h,�Z�3����i&�YQU�oo&�ٚ�z��{�5u����������M�6(�U����vV�+���K{���b��f<��]����t�Y�f��[��*���ʝP��aða[OZ�6sz���ٚu�ֵ�jԲ�5�jB�ae.�ޱ���[�6�j��,��YXӈ��v��ظX���(��6i�M�Ղ��4Ԑ�v�ŋ��s����)�N��֤������fL�+����b�r�,�vƖ���5���5�[�	H[c�늹��l���[QR�GI��lp�<ys�Y�j�����V�3-!���D5�l5��M/2���XU�OSb⩽��/A�jm�uɫ��M�fkq!���ZE�a{9�F99xG���n^�{9�<�D��،�1��sz9;X6���~�6ۭ����5w+:�֔ݸ˷2\�M����@�nNH�d���Q����㮻���J�v59��r�*q�Z�hGbQ�I@��sΎ�����X��{g;����(�`�,!1�ErK���@:�������_'c�=�� �I]�GE9z�]f�w�6x�Y��0��qK��aT3�Ie��ხv�5pq���]{��b�0A�5��lt�X�}�|�>�ιN�ዴ��<mF�y0>Js�yƞ�L�����tk�rq���q`1��Kf=��ْ]�)�{I7�"����c��������m�wa���G4�b9��{%rxnͳ�n9��:�W um-��ú�V�[RYM,����n�����6Wq����WAvC�ݗ�Zq��WHP���Q[+pa1�]Ñ�10��oi���V\MM�nm�a����!M�����95t�u�YY�0�2AɌW\���G��
�ï<�\f\-�5ԣ��En	���Vʻ8�s]{Y�zy%���Rl����ŵ�B�`27�J�v%�����[�<���re��9��kI��8h� �h�,��i;���:��`���S�`����v+q�ԁ��a#R�^�]ks�9���,�՚[H�u�؍��0��84�2qÊ�[�ʯ-BmqF�R�
2��<�γ�5�k�N,IleBjDfe�.l��U��N-I1J�f�[X��Wt����E'a��b����e^E �e���nX&����b��Rb蝛$nGl��P����<�0XI��+�ۛ����ݙ��N�;�ɔ�Ƹ���IY�z��M��q���3Q�Unc��s^��n5lt-Łଙ�6HW�;ik�"�6s&���:,q��WLG��j���B���u�Un52��߿~��ತh�k��O �%��i��8��LCa�ƶ��T#mc�7��$!ǯ��?��q��ۚ����d��7|�<?

YD9V�X^p8~�:w������Am� {�j�0�l^�=7�+����VMM�K|+|�>�麗;�@��k<��Zy���vk�36��t	 ��Wŷ5����}�|�t���f-T��{�׆V��6|A�D�t+��n��H"4����)��Ԫ��A��(��O͹����[�7|�<?}_{`O�l�pp���V���S� ��
��MȐCm�6������������-�����D�P�[����m������èD�� �|fj@�5�gv-����c��\35�6�rB���a�G��}@�� r���;�7"FNg��1��a=���+|(f�Q�M�V�J �d�#���|۟��r�U�ym?\
��<�j�D��d���M]���Ucym)���z�|3Iv��c�m2tiƬJ.��z^b&©�uowEf������xƛ���$����8x��ű�ww�#������A�"�ŷ1�~)�ȏb�+�=��E�~��I���mȈ�͛��0:!f���j��jo��|э���� ����n0	m�͹��=��
�
z�_O�V�ҹ��	7�]ُ}^R��^[#ǒ�#�e�ؐ���Qj�}���q�	m�͹[��TY6(m�{����š�ww�#�s�@�l	���_����^������ӽt����]O��s��8���l+�-�^ae�*�ڰ&�l�j�D�W
��@�����iЯ�mЯn^�R��^�y�)�+�e�n'�/���OLT� ��
��ŷ4m�p$����"�3}~U;Lp�����"~ɼu����.^�u�r<%4A�D����f9�����*�Q �[sD�
��A�1jϯ��^?�)�Io]gwR٘���#��~�U�m�L �m4a�UR��\w7�4Օ (9��[�S�M*ޜy���_.۱3�j����Z����}�?C~�E�?7 6��e��{����jD�;�?Sn�v��� jo������(� �_���Z0��sF�gyD�A:�hӪ�H-�nn��=�r6m�/f-��+u��r=��S_C�!�_W͹	�]���ݘF�옑�p<�3@!֘�"㎞�m3Kқ�����7773��1j"���q�A-��A�
-Ăŷ4=�����xw��a�0�w�[�&��@߈#��P�u9��n@m��n~ɶ 7�?npd.���#�t+ۙ��D����1�%�f��?7[NNl�7Z���T���� Hm�͹߈n_�2���q���_�/Z�Ku��~ǒ�!��u_�
��^�3�b�`�Y�?P����0Am�{˶�:0���^��\�W���^n����*.��r���/)SO#cR�4�,?\�w�6lr·a�!UX��S���5����M��\���Smd}�]���^wޚ ��O�6�����m� �J>������*�V<��^�ow�7�c�K���P��I���n���<��	m�u�$Ѯ�������[�ql��G��۵u��.a�a�\�S�����,�O_>�@���ȑ��U�c�z�]-���v�CΗ�3f���f��r$���|Cn�|[�s��~�.��*��Lx�ď� ���yc�T�<;���|?P �`I��Wŷ.���r�_��O�z+}"���h[� ��_�T�*�x�2k2��tv����s{������l�}�(�O��nh��P�f��3\����E���~nA�z��{ײ�n�\7o=�~��-�C�8G���&�~���P-ĐKnh�ۡE�ظ�b&�� �ڹ���R�����������A���A�B�m�Cr&5�=�zv�f��_BĬb�h�7��/���kj�n)N�znJ�KOn<��W�`a�I�\BxiZ������q�f��k9�Vd����Pt�ܞ��1�ӧ5����Yw4ݶ\,��\n�;q��Wäps�n�����ό�z��ɲP�vh�[=mv�{�D�+�����s���IT+J�%
ѣ3�ˠ`#LcE��n ��m�|��1lz���S�ι�n=ri
��i��c^6���6�j�3՞���(W�������m	q1%9��������M�����|{mZ�e36t34��UK1k����ذ̲�>���S?UQ��	���t���_6�P��Ѵ�Ev���1�=��1�S�,�K��<�
+� �nh��
�]��E����W�4/�c�W�Y�͇Ku��~�A�SD�Con=*=�����~�?%���n m͏Y��{�����ri�ulf�����@�(G?H��nh[�$6���Ovd�Ms�}��nEnn�WQ�v��o���+�5��˙��cD����} ��m�p$�ۡ@������K�U溾ŝ��j��|7s���M_�O�6��m��[�W�^�T�G<�����,��y,1|�iZ�dl�.XcP�6�H4A3�;��MG?��q�Ӛ��ʚ`�;���|?P>�/tZQp}�(��Cp$��P%�4Cy����te{����6��ł���N�A�#h<+p�¨R�ݬ��r��EMTLј�����g�ű5jήɊ�'k<=��U���+�7�5�w7�o�ǈ ����k�-�y�h��u�����!�QN�r+�[s�p#;���1y�ܥV�s��^���o|(|���D�۠+�ۡ@�A'�Q�6���~�"ߨP>�A ���q�i���lf�a�.|(� o��Pn������l������(ۚ �܉!�G���퍜;�)����<��f�o�\o�c�|
Κk��� ۓ����xy���^~���7���J2�-��튼H�ї�ۄ.��pͮͨ5�r?�������A�P�۟��o]]��{N��i߆���a��|7ܧ��"~#���n~n�����ԃR�i�̽[���6'�>�M�_B�`�;���<�����E�=��(�]Wբk�������@�܉����ۑ�IN}~.�v�%���Q7��0��m��t�t��:��qD����=�y&�)������GNʹ�`�[�[gղ��Fl�\o�`�>#_��������΁����A����9�~ȟ��lS�<��OoZw᷾�>Jk����f{��x�yW��(��_'B�q$�n~�ۡ_�-X��j��
��t׹�B�`�<����.|(�H#��(���nG���z:��W	�d���H1F^czc�&��(���W&�+��cm�p�<��:�k��~��H�u_t+��B��3g7�.3�1�+%���x�ᑄ�J��O�=����?�����
�A���6��{{�?!�"a��C�y���޴��o}_y)�A}"@!�s��g��^�9��A�t���
��A�1'K��Ǘ�{�[�5(���5_�¾� �;�_6�~ ���$6�MO(��ι`�H��|��_�
y�5�ћ9��q�ُJΚ ��sf=�x�c�9?F�]�D��S̮zNW][,���z��˧;�W�.�!�R�3~�;F��e�<wĔ��u Wpc�i �����㞉��4��pnFۛ檫��R&;3�:�o��=�i߆�z�>Jk���
���4}y��6~�=�����˶�*���t��c�䭘�XM�����dɜ�mjkLچ�~�=����B�-ĐKnk;�9C�X�ZsU�x>��sbz{4���>�m
����_7"@!�T-����'(�c=Jo��"���|G��Yy~)��;��q�ُ��hF�W���~��I��y����4�HmȢ۟���5�У�تu=X���{m'~��%4>�$6�����P-Đ|��g�~]s2�/}B�q �ۚ�xg79%��u_��SﾠO� �q�8|��}���Y�o([s@Cro�Ҁ��ϯ68���<�[j��1��������x�������P�[� ������}�"rȾ�[�#A��{'qv'��U4��� �ӫV�]��%�`։#܄ ����hMu��g-Rg[�u�����]}n�Ohѯ�ϟ�{�������cG\.��׍[�)[�7|\g����<��n�9�<=�	����3�0󤃶�4��۱&!���$.3sS�L����1T$sB��h�K��A�s�.�&�ۍ�i�(���f��ʶal�d
�]��\�6[�$ٌ�Q�.7W���uuL�؞#wX[Z��Ny[��,"�a}i�d� ��������'��͈'�`�%�mȑ�Mv�N�$#Xi��d�c�)��T|7��	N�u�
 ���H�y�J��g�{m'~��p���va������ ����mР[� �[s@��{�/�ǝ��L߇��INhgxg79%�ŧuo��S��?G?P�ۘtj�K������8�v����B��������!�C��Ew�}S޵��G͜�綠y?xk�|�`?6���VƏyd�����D������AnD��{UK�vx'��wỾ��O�<PV�u�9�o|~O�P-Ă-��n�n:Q֣�q�ٯ��c�9%��ӻ��~_�e#��ѡ�{z�ld!�$���ȶ�U+ �.ŀn�Y�uee���!��ow���6�I2b~�g� 橢�IO�)���R+͜�}��/��޿t�_��� ��E��~-��u@����{�#�����F�k+d��^S��.V�]�A!���<�L�UFIs�Z�Ӡv��E����Y�}��j���j�ǉ��L���[��G9�e����/��I;���P'�MC�����Y�����ohP+"~ ���A�B�q Am�������P7�ӒZ�ZwV�����	���A�B�m����Cn��3�>nF�+�ץ�)~t+�܊y~AH�ѻ9��ُ	�٠��3��V��tI��۪��	��ۡ@���r��(y�xW�T���U^oo�n6�N���۳�!�D�ۯ��܏n���AhOT�	��B MT�U0����B�1/�jD�f�\@Cf]	pJ���,�X�����;���#�t��`nk������N���20�r[t^�
<��4!������5���ƛ���w9|����^�����"�F�������l�k�|�S�8u�͔���Ŵ>�	6�Wŷ4AnE .���nO��� V��p�L��B����e��L+�N���xu]_�L�q�Y��tk��u ����!���Ǧa��SK��7zu}ܳ��z�;y3OK��-�:j�(���h��fbA���
��gy��ۗ�w �����@j���+z�ԶM��4�T���[;�g����n��*�fЭ�V��M��t�1׈*gy>��ӹ���v���߉��a��
߭L<�b칕��+q�u����n�k�5�w�p]@�+��K��:�bf�Ҷ�v��͖�6n�����Zz��,�m,��E�(msyMa��)�)<"4�A��T�S�.8�Ƕ�巊c�_9���̹�U�("!�ҥI�ے�	) Y���h��vH��,MP�q�owsy�y+��-J��݋��6�r68źM�2�h�YX�s6���o���v�ѽސ����9K7��ذ�Į��_��n*�sghO��MN�V��nX�:ڻU�H	E�ףwzv����WQ;�tv�Ҷ��Ed�E�=ٜ8�4�����.��6<ލe�*pt�E8M�љ�-�X^VAzm���y3{��;�����89´}p��O殥=�z�ͫN�u��V2�i��wF���,�`҅� �b��hV�٪*��0*}:��u����a�NO�ggU��:�xl��qSH���L�UO1(�7;1ov79Ri�u����,��{�tT�VZB�<G�J�����޾��0TX�\08�}�,��΃���Բ�r�����~���ߌzU�vYt�3!�e���=
��Vl��:k9�k�r�Q�4��z�6{�x���Z�TT�u�n��2���η��U�����ؠ�����+�J�(^�������l�3�A�5�m`j�Q6�������'��,0t�'A�fi�g��f4��gW+eiPf޽��;9ټ�ڮ�,4�Y�¬�Sj48���⭎����,��{[�s36���5liǫ9�3�.�:�l�����^��fs{5�Y͛;�.8ڍ0vMs�q��N���;�[{��R�4�ga�Ma�׽�+�k5�c�ؘ̥rFaVt��՘������4׽y[���4�[-M37�O,��цs733�Ѱ��V�cj�՜��i�郧VӜj��5���8�fu�Fq�g�j�k���1 ���7UInަ�e$����P'�M~~� ۯ��܊-ĀE����� �T(�D�A-��3�3�����n���.}�}�$��o{ݱ(h;�?WϤ�P%�5���O�6��A`0n�R�ǽ���5!ލ��#��1�A �l�Z�B�q?Am�`uyZr�<Ll��S�(�F8�x��
87e��X��Ph������4�Z$���b��P?�$w�
����/U/-���l���{�=t�ו?gu�%��"H�:���B�n$�[s��u���C�������N���=����Q�����s�@�l	 ��
-��_o��>55��k�H!=�@��������܍g�{4����/���mf4w��LxN����[� ���!�B�����P7����W��M�5��ir��y��I���A�SDo G�����؏Y��zo�3�U���J�f�ڊ���|����F��w+��t�����U�f��y\�Ԛ��j����5x��|S�
-ĀA�4AiЯ�n;���BM�+�4�M�I�b����|9��� ���[sD܂���^�x~��Ծ�r�(KX���cFv8ݚ�m� �$x�:ٖЛ3\�W�_�c>���!zD�u_ۡ����<oF�����!JheW�w/)$��.ws��}"��H ���ۑ��C��7��ù��K���D�?E�:�^{��8�I;���ڦ�!� m�(���g�����t(����^��
��Kn^NGNQ���3¹��,Q�:�>���;�"�nh�܉���}C��vhnD��n���A�H�C�U|[t(e�h�t/D�����}�w�h�OFVG�g�҆���A;�?6�in�A��B�n}��޾�-��<6������{�l�����}@�j�!� m�|ۑ��3#��>��м6��
��e�I�
Fݬ:#E�v,Ҏ�1	�-�H���au�4;�b�Ғi+��V+�)��jfC֕=��|�����5͠�!m��@fr͝A�����hX#C,
���t�]k���m�Y��F�m�i$B�xQYѷ��ՙ(a �ǰY�4`0�7��xv+{t��Ӻ{h�C��K�F:ƻ/N�ۇBq�p/\���E`ޔ�E�eWsm=�O���v�PSׂ��ru��b�I�\�h)�UV���3t�B�#��Q6��f����7�g.xT�.WW:�8��'���,��ms�¥up�˛�d�6������|����Рq �[s��q��+�N���<?
��7O§\�p0oξ�ӿ~nD�۪�����>����޹�p�ޯ��P����T/D��ǆv�{�	�S@~�P��L��LW�{�ŉ/�4��}@���Cn�|[s@�܄�yϳW�7��	�Un��w8�I;���P'ڦ��D�ۯ��t(�A��V����q�>#[�_��=�q��+�N���<?
�`H#�/ʫ�D�`�yt��D�r(��?��h�F\�������PW���B�N�xb��l����l����
��@-�Tv�&_��B����}��������)�gDxƣݙe&�@��e��Zp\��VS9fS����!�嘇���P-��nD���UK���z5JN�l�8�]'u0#ٽ2��lCR$�.�_6�P��A-��/��]L�a�:������M�y���#�ö�a��'uh�l7���������È��u����J9�_Jw�ny�A�j^�nИ�"��A<��w�����Y����~����z�m������c� -���t��r$��W��E��t��!�Safн��bc=�������
-���m�ۡB��9VV� �wP�R����r��J巾^�R��7>�4Cx2�*���Up�u�z~n0�nhmТ�%A����
5Y5}���g���/i�0�(}�$C�P�۟�����17ȡ{��f&D�&z#�g��ȏk��q(z�s�����w33�����8��wH�m�|[t+��΅蝼��ُqC}Et�g�⥑�H�y�� ���ފ�	�� >��2�� A��D���U����z���<�P'ڦ�?H��nL�o����+��H �}4?6�Qn$~�3�����Y��WX���&X�e��XR�)�]�V���Q��M�-�ʪ�h��x� �Wq+��뵛�tep��ś�˪�3)Қ�mF��g+͜OO��#�l	��+�ۚ7Hm��=�Nϐ��p��� %���-������^���a^�� �o�����0���tRa�Q �u������ �t(��9�yŨ�ʇ7�~<�R&7ݵ\������������!�U�nG�Yx�}����?��3k��g7VY+ ���[�%Ԁ�m�Mwf6�(
�,��k����ׯ���?1-��~m���5��k9fl�ǁ��'��бf�@��s��� ��}@������P9��17�	��|~�z�}�����n��a^���o��#}��n.j�w�ޝ����\������۟�s��	νޏ??�)��;�^Wr�nnu�vo���l� �H��mЯ�r(�H�,+V��wQ��9�A?P���A��潾r�FW,͛���0�(}�$�ǆ���x_�y�ʣ�&e��b(
��hL݆v�+�Nv���U����kU�xѩH�\W��Gz��Wj���{��?wϤH!�_P%�4AȒyko��],Ț�N<�}�22�|=���V�{
��ُ�o��[�P��}%�&�Fi;�C���d�2�	ZYDGK�1Pin�)�Pi�DlK.Į�h�+4Թ�E�����a!�Փ}��Wŷ4AnA��^uW���N>{�B��O�mtNj�jvx~�Hݕ��B�-Ă	m�v�����W��o�$}�5��-��e��ؿ=�G�>�!��(��c��`m����ݎ�]�@�܉6�
��ۡc�'�^���F�s��kNEm�aLg�c�o��o�B�-Ă	m�|Cn���o����F{�(����Hs{��Yq�}�������
�6k�=�U�w_]�E����~?6�-�q5���9W����,I̹��S͇�/�f���x~	���_6�H-ȵ�O �3��9[f=ju�S�8��j�9�W�M*i8�����Ԗ��:�9Ⳉ�
 �^r`"����]_V�����,�̫���ɷi�/e�6�;t�nF�V�h�]��q\����"��hQ-b�����M'����>�]M���_G�K�4�1�%i���ꔕ�F�Uf�D�F�]-X�.Gn^n���H>���<	 \Fθ�qǄ�����hy�=���1b9��0��|���,nK�GW	�xU뇥���C�C�{�Զ,â(e4^����H��k��ݽ1�(����Ů-v�1�\���c�X$MU~]����MB�Cn���mЯ�^f�.�9��¼3�1�FG-F��7��)��6MH��D�A�����@��	(^^�<���w���4AnD��ޗXs{Ż�����_{v~~�q~�P!{ք�=YB�8�A�t�6���%�5���B6���v_�V�n���x~>���nh[� ۡC��g]�yU��Gt� �]_WŷB��4r��r�s֣�������w>�n�u��1F=���$�Rs_ۡ@��I�[r����u|��f��R� %\��a�y�-�No�^�����?H�s�|ۡ�����䴠x�"fjE	�R"�N8��k�Ȍ��Jun��i�j�o����q��̐�Ȣ�O�[s^�R�ggR݋���0�C����F��Ut�9A-��?Sro(ۚ �_fj�����e��.���ك�+h��x�����{ɣ]�A!�׽H�Լ�_��)�A��5,qz��{�Į��ɿ������y�<��������lǈ'9Oվ�
�3�j��o�.h���
p$�ۡ_�� ��G{D�zg��v��a��^-�No��}������
��"�n'�G{��8���=�W5�涾N0�[s�%:��Kv+�c�����1�룮���nZ�w�h}�Cn���s_[�$6�'�M��^Os��Z�P�X�]ZNUnz��lǁ�������� ���_�Ո����d��H�*DAKk4�ָ��h.�O�XҶjIn@��m�YT��4�Ǿ�$7�B�nk��w��:����wS�÷$r|�A�$���HO��_6�WŸ�	m�7���U:_[������)M3�{in�y�x�
l	 ��P�ۗ����������9�_��@�y9�r$���M���9��}V�����Ƶ܈Y�c/h��ƃ��y�'J�x#�v��]�ÙAѣ[H��N���9����$䛲��S��m��[��b�� �ozk����q�ۚ ��
��kp��}{�
��7"]�򎡙o=�����=�>ݚ]�{��8ő�uW�/u
��A��� �ۯ��R<�I��^\������{in�y�p1���H?wz��� ��JÓ�'*C�?@��Л�+��Oe܋��M���J�F�F�4���ъf(1��
�|�?{�I��mСy���탳[����#�v�{�PL�O��C/�@ �[sD6����ܵf���c��g�M}��r%ߖ#�3-�[�����@�n�|/�$��؊(?x��@���yP�mG��I�[u�q�Amτ�W,���L��g(�Kv��;���~ ���[s�p3�t(:����zp�=�C�U|[t+������f��z��G���@�}�/!݄D���S����M9�u�	Л�����c�r�yj@��f�R�@��kO��ķvK�=���g��x��y�X�̣^7�]?6�[�%�B�nys��	�z���\�y޽>�X���qMp{~�A���!� m��ۡ��Z�3�Q���K��]Z�uE2X@{�>uK,<�F�6�FͻVYh�P*��Y������z��$'���<|�q�ۚ���9G�-��=���,������;��P�yzh��H!�B�-���?
���_�� {ޡY��mf��z��G��9MF��(���Ցz �)�G7_W����
�4A���{�MMw����n�eH�w��nZ�u�	��� ��m���q ��׆�}럟��B����m��y�H垝[��{<w�}�$�m�qeC�>�VO�=�$��}@�ۚ � 6��{����=U8'�ML�����N
ʼu��yDp�������Wȏ9��$���!$��H��! BIA	O�H����	'�$I?�! BI����	'�$��H����	'�$��!$�H����	'�H����	'�H����	'��$I2�!$���
�2��Z�_P3�� ���9�>���`                                     �
 �          �                        @ x�P����UHE��P 
�)@��	Q@�R�HI*�Q"R�Q$RBJ(�R��    )JJJ 	��}ew�BUJݜ�J��OcR������ު��{ҫmr�;iW{t�T���Xms��*��K�^�;9V����[       Nuy�:0�rε�i�}	*�^l���ԩ]��E� �g@^�{  y��T�{������;��{�� w��    >  �IDP(J(J��H��@Z}���B��Wwp	^����-i ���7�)f gw�TOEf�
     p�}�q.`;�B8��͈��P��pF�"#�J�1k��a�KwЀ   �  ���$ �B)TR��$B]��������zaENa���w����hx��g��f��Y^�r�ԅw�z��M��*�� �ܕP��=���$(  ��S�{m}�:�ҕ���h���ҩVw���E�֭��%J�r4H�͕�� �u^�l��E�wW�4���J���{bP@ ��  |��@*��UR�IO���5�c$����JP��{�ZB���%R7(-ޕ���܅R�w��a�E������
�t�W�n���� �     c{�}m��{�Ԫ����:^��vն�۪R%e����
�0T�=f���el��UU*���5��v��h� ��  ��AJP	��(�A@UޥW�\��*���U+��U�{u^��<�J����\��iU��EOw:UBn�*�!��[�R�����[���`  ��    �:�f�E�u	U3�R7T�\�'���[�J^���EV�Ъ�ܥRWr�{���U��:B����)]��"� j`1R�@j��CIJT� ��U*T�&@ i�T�)H  )�����  "�)M&���S������~�E~��^8{�z��]{�^��y� �$�Fw�$�	.$! ��� I_�	!K�$ I1@$$��~�D������w�����C�\"︔���śx������=�/�1Ꭵ�%t]dʫT.�H�U�0��ս�SHY����n�J���N7Bd��N���
�8
�c4��qՍX�3N�,��R�x��r��b�F�n1zZb�7�)�s^�A�Z^�5Dj�۠H�B�L���[
�gCF��X�ߕZQɢ�)�kn�N��:��h��'CN��1�A['n��Y��[z��t�&��dW�C&Iwn�^�����Rޕ��wWZ#p*݉�&)�!���ɗA@�V-����75�q�3{d㷱�5�3�,ʱ��TX�+Yc,�V�Y��.�r��lî��W�`��S)�{�2jj����Wq���`��;���St�Q�F���̃�6��rM���(i&�R�]����$j5ajq�S[���R�iͬ��$j-���]Vc���P�d���1V�	��״�Y˷��V����W����9[�B��j�h[f芳�i.�n^�Cn�z��yF�`&Q�٦h7$a�_)Yi(�T�\
���ܟ9�6U%k�d,;B��GF�UhI�^$]��o,Am��S����4��ݿ�C]���a��kG,݆�eʪ�U=u^J����4겕�YӲ�9�v�u`�I䭫f�t�U^9w�����5G3�!t�"nʥ@±����������1a�e�f�:T�O"�+0V��h�R��m�N�]�q9Z�7�	+�R^��!���fn�Z��lОLybmu��f �������*��,͛l����Ѵ�<���7l�Ȃ�Xs�����b��(�C��IA��p���P����8�mi�E�ҔS7���ɓ/6�܂�ĵ�����V�j��q�[k�QA����vΙx�jě�Q��+s�ق�<)ԛ-`h��CS�[a��AAr�B�Gn3�w��q5V��Ye���f�����cM�t�a��ujd�Ť/A�rnX�%��.�j���Һ�!����q�MuU���бx]�g�o�l5�P���Ԗ7$(*hi����q^��N��������37r�EEʻ����ޗ���b��PL�Sw
�E��(B���vY��0U .n�*e��:���R�{�1U�6��4���
,��n]���f��XZuG�Mө��!/&죓;�C[�t��]��ǂ��f^���җI_�#�cX2��5a������u��Fެ�%�J�Q��Sm�¥��ɸ�
�sh���K���e�y�/.�2���mѰwr���@�YCtj��(+rM�&4dŹ	�f�P��0[ڧ[b�k��f�6��&7�f�`�̼#i\זb��Iudk:�UY�.
�w�+b�:b�V*�n5x��̺ۊ�����e�^�dۻp��.ɬ�\ׯc��k�w����z�w�Z3\����fTz��u���p`Z&nL%[�Dތ��k��0��ft"�2���vs�u>-]�r��ۨ%e4D�ӦX�XXe빆� �eVU+y�Vk��Nk�{BͺrZ�L���g+I�%��r�e�F������:t��!���z3�U��k��B�@o[�{M^n��]�UN�2��P�ʼ��m^cQ�$NjiTV7j�)t��I�N1y-�q�Y+V+���sA���B�U�b�M�@�1��$������TY�K"���q�̇T�X�!��{H�x$�C�UF���[� �PYF�*��I]	R�a�r��7/nfF�D��*Z���Ί�i�Y�y*ʁn�-���d�R��vj�z^�v�v��ѵ�y�%��&c�p��oo.��5AԘ�ՍJ�YF��q�dŲ��qҵu@��Pݣ�к�P��nc[d<6�%`܊C�W�j��Oo�49F�V�ͣ��Y3mi҂6V�ŕ�1nB��IUN�:�N
ɪ�J��	Xۭz��6w`��9��L�hj�N%�$�{��5ee�V���5
&^C[��ݬo-,C�$l�X�TQ���6-Yʂ�&ȅ�޼�VKҮ�r���*��"!�B�S˧��t�����fY�X��U�w׷*תc�H˦�;(��j	�Kie����W�`y{�W+Q�;��Vm��Vo4S�6�ULY̭O�Z�f�O�+�?�(��I�	�ދ��='2:��
���F�XM��~�wı�)IZ]�({�*U���(��VQ��ٹ,,�kLJM�T�=wy��x�,���`����%f��n I�Pn��"���,)���+���l�*�JZ�ͩ#�����N�[`��_n��o~�[��f�����Q��XI�UXb���V,&�ϛY��R}��MQ�.n2��V�zġ���
�+E�y�����G�f�tkna��w�i�ȫ�J���)�r�[�z�&����Ӽ�/*���+�}�j�֠s3VՄXf�ЖX�W�w��Ax����K�����UsJ��ʥF�6_c�(���l�w��!$�j���Ɯ����L[���;rTb��|�����HS��N�i:�ܑ�5�朗R�V�ɩb��ʂ�7T���{�.+ߖ#b��h����{{gt�V*����tE4�ԥ��H1ڙ�j��2k3.�]f^���j�_�.�n�/vU�:ofi�Y�tޫ�6�����;�,H��?��r�yY�56��ʥ��;��9��dx����W�����/6\������:N�w�!�P՜�d�\����x�9�Y�����2���s1Ŭ��Pw���#�� �ں���Q,��P��u����*��f���L�G��Z���u݋�fVf��v�݋�����{��6j�䷘�ܼ³Xhӂ	3�Nf+����a�4^�H�2����u�,�1�(�&�J�*̠QM�khR�R��R�{��6Q����,\���,�Q{vռxù��-���r�Bf�O�Y�tX��v]76ؗU��H7�O2�AR��kõB�S�׻2����V�8�����,�(]��u��k"�q����Sݕ�A��{��^G�7r�4��2��?4�2r�L��d���6�(^�W�i���Z(���k�T��ͷ�xK�paْ�kK���ѫkse�sN�(Ԭ
���J�ՑW�,:I���ek������E����ZڗU�HV�#�1�Ye�"�8������Ьٙ��
��u��3v��7%��Ȳ�F�����*R�Y��mR�D.U�W����W-�Ǭa�S(S�-	��]���ɚ�՘4ò��'J��eh�+��ګ�TJ�j��sl��z#��{WOoe3�֍z�!��T��8V:v��d�r�鵘EdR�fdf��d))�.�*��A횼.�$1�ӻA�]�L�l��J�Փ��6�X��H��C���+EVbn�������!���M+��Wm�j	�;A�O�y[[_7{�l9/q�vb�N��ˬر��l�1-I�Ö#tr'T��X�dڦ�r�v1J�LՉɱ]�r�eR�r�ɱp-̶Jʙ���2U��I�5�ޫ�V�h5�����/Z�0!Cj�йSl4�&�A��i��32�V�Ǘ�a!�(��QT ��),���u����;�z$�V�t���Q�wqa2��6�-�t,�w$QHv��,�(�L��e�����j��V�5:��.�ơ���*�`��/pf�j��{Xj䕃N��+Nena�[�]na�GEJ�v��Dibe���F��EU]�U-�d2*�*��1i��6�P�W+&]��W.�ꪯm0��}��<�f�>��R����mH7+Nfi��Z�.�P[.�k%��ո����l���u�a�*e�ٌ���cj,F;Kٶ�=�W�Y�P��aɛ[w�f��B�ݠF�U�b���D�b[���U��@�n6ŗzefF���̰��j�uzPr����U���܊t�F�\B��C�^��q3v�&<�>Y`ɸ����M�3_T�7nb.�T2�`y"�N�MVa�������,��-�{I�5������w�R�[��2mj�d��UCYI�E뤳*f��_�-�ZPU�f�Z*�q�YwwlZ��3O0k�V%]UJ�B��_*����%�~cV��VV����5�%*_B�ѦS�y�W�Q6�+ś�������V�i�̣�oU<۪�C�[.I���Wnnб,��*X�4��7��[D�����c79kT.d�&H����9��sP�V�W)EV��-�+�j�-�im[��ʤ�f�^;�Lɲ��Ѝ��V�	��ehH�c#r�j�;u���-�r�j���e]�����<c]��[�6w���y�/M7.�f ZJ�(��b��V�+J��U�*��7sr�kL˽����ZV�),��GyF���wv��A5���YiQ���E�yV�Ua�/r��
�r��(��gS�Y��q�(�-eB�k�2M�̳5�`�zޑ�%&KCNn6����y��*WZ|�7�E���h�*�;�ź;uyQ͸��/@qBѐM���Xp�WBn��k
n��70]V,�׫l��Z�5���ۙ�F�M�u�����`��1�5�|qf`c\I��&R�g7un��.���淛�PZQB,P�qayl��(����Y�n}�͹[�{w$̺&e��e�_�d�(鬛a���bEb񇕘,�����
&��hfV
�=UM�Q5,�!��4Z�u���b�K{g�pXۋ�*R�=��B{V�uU.�aW��[7�q8i�d��,L�T�'�<N���&�U�(�[T�my%�h�,�jKȩ�jbD��q�B��)r��J�]a�b�8�R��Wr�E,wU������ŵei4�b���u��n�5ؽ!�f�Vj���T�jhחNZ�勲�f�U��P�((�@��fQF)�
	T���MMԈ1Wy���uq�r�$�Z��4.�1���zq�{�7m�9hQn+��1L�`ؕ��%Z̲r�L��7T(�yV�Q�PH$?Eg���^ٗKuf��l�+~���j�/�f z�e�+/�c.�ea�U�Oe%C&[�FBas���n�'� jm2�r#RQS����z�0�NmfL���P�ܳ���������4BM�ώVng�N��R��
�|N	
Vo\�wN�F�ʼY�����+UaA4b�O[xf-��L�c�V�:���hiՕ4n'X�f�}��Օn�R�]SȯR:��i��6�Ӹ�td��2((fQ�FnV+RI�pe��j2R-jҍ9h�;�1*�Ai�M�
;3kU�j�K�"x܅�f��7h�1b��*��;�N�`�u_V�W0k8.�̂�M��F�YH�#�5Pc2�f����0�ͅ�,p�<�ae�l^�ٹfY���N^V�VC	��˼:��WJ}V�\:�ٮ��\{sorͬ�$�����갶��I-]n�ʼ;�0�z�!�t�Ͱ�d*GYl�.���5[V�Ct������A��zRw3a�n��sM�.!�@r^�srUS{zw4�X#�.h�b��)d%j�4UYj��G����,c��Z�[X����4sjhg�hfe�ʼұ���Y`ʚ��v?��Ly�K����ʺ-4������7s	2�[�Y8r����P]I1�=j��k+e�b#6ȋ�WV���$��%�l�8��v��T��qS7(�ART����4j��b�wU�����Q�i��UU�V,��)9�6��w��@ù�'ZP�Z��fm�Yd<6��ݴ�(o3Z�1��u[ �deR��1�t�ѷ{�-U�42b�xiU;y��7i�e�Vlb�Z�:�tQYM��J5.��!(F�6��M���^���*���;Q[6U7U��xŝy,ҷY`���ӭf�R�fmֽ�M;w1��\���¬�lm^���a��3S�^��$B�m�Ű�6���[��ti��U5bu���_"`��M����y�n����[gi5L�������U�k,�m�/.��w�]��r���Q����U[��nl �K��ALݼ9�6��u٫�g�4�ĵg,P��L�M��*�35=��6:;�3޼��mQ1�˅(~c2�&�;;���f�Z�ͺ[KHIe^n˽z]��m�T�E-ۤ�6]:�n,۪m���#/p�YD�mR����V�m��{uIC��� ��w.ۯ��V�^�a��֍��٣j��Ui^P�%�ՙY�������xi-ϕ�ʼ�{�aHɣC6�\ѵu��T�U]^L�Un��-�m�)'0�B�
۲��,ޝ�̃.kb��1U���3v��H*k
8Y��\d�N�����u�٩��M�w�X�+��b@�0g&7U�*j�\-���������̩6�x�I�HZ��d�wB(*�����E�OM�ú(^J�[�^V����Ϸ3�Z�7��ٷ�ּR�齕3n\i2�bnU��L�m:B%ȭ��+uL�&;�iJe�wB�i'	go%�1U�Wt�hʛ'��QWѻY˂��J�q��*��aEr�����3��`�E�mՌݚ�U���7bL���U`�bT#.�YR��N�Qڛw"����xqV��`��N]U�HJYB�3~�.n�H%�I��	�\%�Ѫ�R�a&�V�cef�9v�ӌ[GsCך�n�*��eAE�f+�2�**��XQ���^<�EL�-�կʘ-�c1<ϖڧ���L�{gt�ܴ�ʗ,�qTg3q�7�r��"q�ЁǷ��j��;��yV��b:���X��)�F���mJ��%TVu�� Y�B�hƨҤso*�!&�̗����:��eDf�WB���+�٣3al�C��Iz#G����d��c'j��UYT�W&v�ܻ��!^�Y�m��
=��!�j1^᥅��k橴��368	�H֎�֖�f��-mtu$�g36�&\����S���K>�bT�t�	��J�f�:�i\�Z\�K]x����ZCi$&���$�7t]�t]������\]uE��u�W]\u���E�Q�uT]�QuTuwTu�GU]w�]\]�EuGWq��wT]��Q�]�U�q��q��w�qu�u�EwUtwuq�qwq�uU�wqW]tWwu��Qu��$	��6m	m$��BI���:��몣����������룫����:���誨��������;�����+�㎺�����"��뫢�����.���ꈺ��.��:ꢻ�+��.�;�*���꫎�+���:����*�6�$�G��B!#���}�o���p���Mm�6S+%��.��k7,�7��V���ێ;X�us�T�\�7u�ǽ�Z���b�Sr]*,=��}U�iKO/��ï��
"ȑ��;�/����x��1Q�iR�as��_^Rd��Q:Ҿ�,���w;*�ige������8k��e؁���s]ثX�JYF�姝��#7�>�U��v�;�Ʋ����;�sT����L��F �<�Ie�J����i�嶶�������Đ��"M�e�3��weP޾��ߘ�Y�����;���wWnY$���}�q��b�{U��	�w\��Ga�WUk
�qٙxK3��U)�GVxk3Nj��xol����]w�ظ��JAKΧ��Q�ɷ�;n�h�H��~�wW�Nt&Vn����O�82m��{:�V9s���}���(��[�4��6�]�,�ʝv+��:�Z��ˈ|N[i��v�8_X����Gpr�(���ò���=���7U����74�����=�p�p���r�D�]e�er�7��eI,�lʬ�.�zƨ�z�stПk��4��*�,u�aݦ�oo�^�⳹õ��0�u�n��[���9�j}6���uvF@w\�"��d�W�_���*�������t��۱s$����1�3h�Ť;H��R���\�Hޗ�Jk�k��
���	5�oY��.g.��'3-L�C�1�#��6�����]�_^̜J�{��+���V�<�Yz�������eh�S)v���^*��+}BU�=�Ğ���5�(�Z/oo/�z�42�Wl.�C۳��*�w[��{�b��9T⺆;ʗ�f���$|�ʹ��;Q[Y�_L��쌬ђ��
]�yL����ͮ��8.m��ǍB��RKJ�A��Pg��W}*���U���j�n����eV�v)�f�C��Mcܛ��k+�\�o�Ү'u���0uǎ`з��R���i�&:	�qd��e[Ԍ=�r{}�gr�z(5Tz����ʰX��j���F�d")C]�� 5͜�t�ע}
�b�[��[U ���r<8õ$Y���6
\u;��BLTlq�����hͦ��m�CN�w[ZM�u�,)y��۪�W�t���on�ݭڱL�ס�GV4D+��;�r�7�r����ʵ�ù�j�uX�]��w2�껤�P�cr�9���Z���7I�q9[ՊX̨��B�N��A��ݻ/�F�L�%n)�����H^�96�ö�ҕM�ۦ�)H����XtG�m�lq���Z97Z+Fkʆ��p��'�W*�sH�k�HWi�ȨV^�%qY2��Z��RS��TCa-��gu�ҹx�P����\��W+�i鸐���\�,X�f��3�e+�Y���V~�EM-Z��os��*�Y�6�bu�ڼ��6.��n:-�n��ν��*(P."�ͮ6:�C֬�yX�^��T��M�d�%���
R0H��U�hWA��'��Y7�7;��_-��:�K6�m�J��u�;6�n��5��*P$��i]G���E"n��N3(b�ƈ�-��va��w:�;*XѼ��;
i�c6���Y�S8�I���ǋ����h�QJ���f��N�;%�!pଣx���ըląG��Ź*��T��돆�}�����5��sE2�����ڮF�:ҩ^�[ӈvq��,�w�����7*�����z+6���u�+*���	<v�ބ%VeWr��N� k%���Tɉ�Xi�]JSGd�G]�6�`�E+�̊����f�v�y���J���))��c�K+A��^;Agض�Xz�����
�k��)�ʢ\�
n�ioK���t��u�ø7���R�ѭS��I�L�ow,���L��6'J��f�������̨�Q�����0At�5ؔ|���K�G�5%yK��F	�=7r�;�V���m㗙q�v�^D�t��'�/>�ʮ�sk �J��6��_f�۳-̢�� ᣍ󬙣�vv��Z0�y`���ZK��.�$6���f�a�R�_Hm�P�[�k����Y�Y70o�;/uK9aX(�n�zp3[��"�#�=����oE0�Y�}�բv�;�#B�l
�oe�n���]�yW����7��<}Ƙ0�eob٭а^�d�4݌ݧw�1"wX�{5��(�gJջ]�\ݥ}�H]���Y�yx��F�oVpY@��=��޴�MEZ�o����}�nԴ+r�T��8��V/�rؑ�`�Mf�]@�a��^a�6�m�PeZ�������|ق�-���v�9���F�v�wvk��gsMB�<��-��ߌ7�u�6����,n�;�l7��}kFUH;��X�uV�=׮�Օb�,<F��7�Vx�fr��՚/x;�����6��,e�T�eH�bKtY���y���45v���*�:)n�]�gm�d����YЍ���;���)�Q��9B�z�c��7F���.VnS�=T��zZ����3�D�tsƞ��;��ݰ�u����[�Ҝ7(������vyZ����2ahQ��o�tκ�Z8�q=����r!U�5.U���<�tvVc�;dH�m��7����+��Fuʍe����EX�-*GVk"����y�!M�8�u؉�c���P��ާ��)�z��m���#�+��%�+�Э�n��d������%�i�aҖA�����ӡ��t�<�[F� �m�Wu[Zr�i���j����&q���4qt_-!jVMŮ]sY�IW�cY6��ʯ��.�]�3sg��v�Bk''öM��C�]�#[dI+.U]C;#������g�6w�8ʬ��uY�S4]��L�y�o6��4�=R�/h}\Tr��`㫡��a8�ӒP���g*l���%��c�i�a����̍�I7�r�mf����s�.�R��i�U5�4�(�廕�� ���Di$g7Z1�k+/`Đ�	ɒ�\ڵx�:�±
�%;��ӱ�-�{��Y����G�f��/hRݪ,Y�+��#��.�nN���R�
�E�X�4���m��b��wf.���wn�9dm�r�}�4�Y�uJ��P+�R�]%�d�w��d�3wE�P�M*#:�nmeQ�բ΃���Q�e�[�VV,oY���ju�E��P0�͇U(P��R�PוF���8vr���wI���ۛI�Ɋ�s+��"���n��-m�oLٶ!ݬ:G
]ئ]�_F	`�L�Õt��)�e�ͫi�FX�UN�9�ݭTvY^���!�,���]]U�k��v�fAA�i�Z�ʬ�nV]$�c�,���c����O����=-����{c�Rӛ}Y\6��p��Cu]��Le��}�UX1�et6���VP���#����v�t�:;�;�����o]{p�M�Q9)ug.f=��Pc=Է��bi�9������mJ��!��]R�dTԭ�F2I�\k�Ah�����ra6�sˠ��y�}I�wqe36�>]77��Т(Ǳ.u��+GG8�8>[}��7�̝K�g���؆��{��9����]�{Y{T�Jh����ofS��A����s�.��o�ۻ��"���B���e���Վ�C�j�.ݔ,ohr)��mt8��,��{UyZ*�Ť�L��#C����[�tc������]�S��X���q�C��[�v��n���9sYD]B���-gUAa���`5}w�u�A�z{/��{�j�A��;l�7nP��UG:���-�S!��),<k�Γk�ķ,�Yt;r��e��yx��à���v���VUX�ѯePW\�^���;�:�g�[U)Qч&]��ۜD#^��4Oe�2��/�mY����d����T�9g���f����v�Y�Ċ���eKʗ�{3{�x�uK��i�֕&oRlcLD��ܷ<��r��WM
�r����9��C�Zn*;����)��&�,u�ve<oE
�V�t̫�8Wm!j�e��;9�P���z��C*��Y,xMm�,+�(�.�I>*Wm��u֯Kw�3uv�θ1ә[+M��7X��0�ܭ�l���9���ʪ�%eU;�y��ZyYz�æV�d�U�Z�o���vmpv�b��zF��DRy5r[z9�r��wX�ߐ��W�s>�u.��w����|{�7��u��4��ķT�u�Ƿ�Umd���ˤ���i������*��wc{����.�$+��/-���UU��dgP;T��A��.Ǵ�W8����}��Tw;"U�2V�h]2�II���h������qD�]��V�b�X�lVwU�W�2�U�Z�U�r��Af^g��Rr��R�UW,J����[P���+������e��Z�h����DɵJ���>��J�FU�']]_Zn|e�~��êN��y`��;5b�o->_Pkv�{-�����Z,ڏ��E��;�o�^L����4G�n;o-U-[� ��$9���A�lj:.�T��%�kZGZ:���gw��gg�2��0�]�[{X�.Σ�xnQ)�pW�Z���5y0s�X��<�D�P� �)�I�]}��հN�c}݂�:�z2�K�ݍi�O�4ݶ;���%�r&�j�Z/�ܕ���4�C����q���m����
7[B�q�bRgs�$L�RIu��#`[���r�,��qO�P�	�/���Pq��uQ����|%6��Gh����Ka�������Z����A�7���9B���ʊ��u���&Jtv�Xn�3��ݧgj�X%+�h�5���n���ܭ��*�;�Ռ��k��d�r�k	�o���yY��r�M
�kAuZ^]�XR�ܬy]�����vd���b�xtז1j�l�Z_)މv^�F��-��=A��{X�ը�o$�ۋGuA.(3�,V
���S���he=!���*������O��=��a=1�y/�53r�ܫ�U��/�VU˥�0 ���g i�'y>��`�z[�}������4c�S����wK>�����s�b��P��믥�IB������"pwh-�W�˻�y�Cf�ъ����sg3Ugr6v��D�Q���WէrѺ�j��=p�꫷P{ugz�e��B��C[�����Cγ�_i�Փ
b��I�|�9�CU���U�R�hb���EϒW�V�tNIǴ�����G]�8�^�,�������su�w,K�ުN#�ݚ��mE�ޮ�,�3��9�D���a�wMb�⛹,:�T�%�M�F��SOr�Y�YR��)x�)Ƴ�("4Lɹɱt�������Wv�&Us
66�*�nv�ZBz�,̬8�9���n]c�V��R��h1afh�5��#r��a������ܽ���J��α5��6�+f����`�'��kr��*��{p⽙+�r������e�'e���
�Y/N�m�*�^>�}��f�J����O�*j�ʢ��l��P1�v�H:��κ��y�`�EJ�Jvg]l��V�xq���=��1]w��97;.�Yi��4~�v9��r�A"�O+Y�G�*3&p�w�R�0��)M���K���^����ͱ;�{a��W44ղl5�=X���[&�uXs��f��S����lM\�f���<����w�����yZ��j��e�(҃���;ժ�^��*�us]���w��F�*7����;y3ǹ<1]���od���͠I��D-u��kz�ڡ�zAqh䖦��X�=�ɮ��0�;�mTd6�i�F������
�˩��9������v���o:,�U��'�V�M�7qT�X
�T{ ��y[��v�F�VU�<�7��W+�J�:���u�$��|���,�`̕]�l��-�g:skPtw���\U���3���ѝܲ����S͡��7�%t�����:��_C]�u�Ckj��+z�J��uY�G��k�BK5kn^�@��;O��<�wuJd]Ӥ+9wUnЪ��y���E�U���I�����&��]�щ^�T��"��kv������q���|yPɵ׵�J��ut��M�HT�&��]���ڇ!�wp={NUq��&��a��m��V!\���7%l邧-��5u{ �j`r�81B�fU�*��o��a]"� ��V��<���ջǈ���w�ZN��Ov�s���rE.��wo.��Nay�c�6V
��.��{%�L��^���;���h���k7��9�tDT�;tۛpeWa�75�y����jg}o��Z*c5Bu,"�Ue��&�n��⮥v����R��`��16C��vn���9.�g?��y�X��^V��'�^�zkuXGN�[�k\5,�7�S��뚹RKq��V��U�N��HwFe)Å�qU��;:3����p�1�/8n�yA��{՘�倞ۭ�̀ۋ,�@�=��/6ʡ�8CI;$MN���c��hM˔���]U�8�Z�\xC�v�P���$��K�H6sFd��3ۖsR��=e1}Z�/(�+w���K3_��9]n��\��ft�o�4n^�{wA��YmTX*�{�J�٤rwRZ�,G68n�R�v�ލgO��bv&���˹����Auuس��Ӊ#q�%[�ي��nSB�Vt֩��4x��4e�U��UD0��ۋ��U�'K��.T�<wk���+�bM:��z�1�G��H�U��mc��y�##jQr����_hǝ��L��*Vѧ}/2�VZ�}][�-eK�8�XuYo^Ă�����U���!�S���"�#1�g"��]l���x�l�:�ŷ�&���wB�0�Di���YXܻ)R&$&���׌M���G/���/��&��!t�NЭPwt骪6��L߫�Y�z���EA*��p?r�{����҇�hO!q�
gO�3��do�믧Va����R��݃&ڥ���7N�vI���]X�G�7TR̎�UG���7N��w�Wf��?wT;���v����&����cy_H#U�t������gp��e������w×o�@�$� ��7EL�UO]�'��s��<^X�=tm�mn�Hn ��ˊ�Λn����qK��YfSv)����&�.�u����2=�Z�+��})�;@���qi�wG���Kr�t�Tq�!l���C��:��]��w`��6K4m%��6&�+,LQ̮�[1��pX �I���y�t\�b6w��<b�3���f�iK�&J�;>�C7k�g���;�����ة�\���\�R�f�M� e@6^u!� Ս�dz��:h��ol68�Wbs��t�;�Q9	�N� ͊��8�x.m�y� ��N}��\F�H����y��k�5��,\�lp�Ϟi�i��ס�)���a���J�o=�����5�Tnư���V:K�����هmb����(��ե��q�vu��=rv����=�$���`�tK���#���h3*����89�m�����1�� ��7Y�.���3�vܛHEЎ��k.�� XnR���O������pn�PҚ�<0q�2���um�%Ï;B��o���wRk�I4���g<�R�^n"kr�1��2�a)8%]��,�a0v�;<�ư퓈v��&�sF�X���l	�8���}mh)7 �mdQ�6�m��41p�h7ؚDs��+�Z۳�H�G8�j�����j�[ub�MF�i�LY�İa�A�p⎺�n#�k�x�����ф�{\�fݷ;u�Q��z�[�n2v�lpa�cp��a��X5�8���C��YN;8��ba+.,7��HB�<K�h��6`G�v�"����a$����z��o�M��ķa�N�ٹ�Zmh
DI6�۵ :�f�z�q�u��癇t�/��񽶋W8�t�۳�ܗ]qO,�YD��l�"^şe6��u\p��ئ϶�:nu�=�-']��o�w����f=�+q̸�I��%.�xXGa�o3L��pEƐ=<�	�9�k�v�+����3dv�,K�+W].!kf�X�@�vѤ;Ko!��h���b��Pa�M8z*�wi���Ō���phk���� ޳���p�^�(s�:T�&�Ys���bEĲ�֑v8y�����먮�r�ٍ:�z.v�G4��]�;z�q]}g�&1tDϷQ��X����f���
[����q����p+����2�e��Q���8�{	�p�1R�r0t��Y�V�����K˺�k�M�Y�c�mՕz���n�>�I�g�hF]Z}ɩ�Ki0F�kqJ�,�4\3W��"N4s�籥݄�S5$@���O<,y�Ҡ�{�W!�؟:�}��X໌q�Nϡu`v1�vL�u�b4J�;:��<rc$o)6�(��D�wSjs\�,Ic�c���L�h�A��x��wK�x�oId���j��#;P�x���s�8; ��~7]{��W+� �,��]1bą���3��6�ƌ�O珙�|qZBV�4޺ɊQ6���;@��$��Y���n���:��FT랪;j64e�тD���,HVT�DT�Ζ ˞SͶ��[<��@�c�n�'�t���.t<E_���̄!�I�V�Ш\jt�J3p�<���;ر�b�n��wWTq�p3qtO�ъ뱨�	x��̜7�LWbkd�q0��>�w�Fݶ���=������n)i�dMn����|ͲJj��hz㱩��ͻv��w��`I�.tL�m��.oY�m������,ACu�a�ż����GP��՜2q�X҆�/onu!�.�*ʳY��)��{q[�}k0�E�t�Cq<�t�E��.����ۀ�؅��9�!��3�$��٬&������ܚLfA�M�7��1�`�T���� ����G]�*�ܥ���8ّК0�M���4ḶM��@�K����6ip�Z�%!0��;i�=b4�14%Yi�ւ��X@��v�\M3��ip��1�-����1.5������z�y�BշW!�6���#������$Y�=sv=4���jM�6nJ�5K�K45q��%=t�v:��*���]hL]�����cL�3�����b����9�8Y�v1Y��2ؕ4R��%���t7Z����N��f�,Gi����D�n�����瀼��+�>�`➲V.Bm���	P�\ .{*�ɧb���l�V9��l��t�����O���k�c�8��眳fڼ���Y�'I=����;[zŻ/j-?f��NR���As��m��s��6�X�e�
:u�j����/7H�x@7���Z�ҊFnPS�n�)���n�E�f �'E�u�eҜ�M"��7a��K��4še��v��[bC�w�σ�8�1�:��ۆmN\M���lV�AҔ��ม��!6Wh����^R�u�<3�mO&�f�;s��ױ��k0����bKuۖ)/-ƏNVq�x]���:U;qtE�!V�^�fX��bh�Ɲk���O<�f���u:y�p��vx.ݔ�c��uZ\���o��.e^���=���8e����p���l[6�	S�y�.����W
������x�xM��4YvH�m�t��su,q�WQ��\e�������yیĆ�ɺ��s��q�m�l�Q�e��-׬FӰ[u(����vo`���W:�д(����x�v׊����u��`4v��6��(���X�pD�J����p=*h��h���%a��l����ct-�s��i1ѣ����<Grk��AȽ�Ƥ���q�0/g�ē�{� ��8Zk���itZ[4b�%a���iGv��trA��{z-D����b�nT�lͫC`�mm]�t�Jr���Ysݓz9�ӈn�G��3Ͷ�
�F�On�80/j��`�A�r���<X�x�KJ4���ĳƲ�����Q5��(D6��r��wh�Z�aN�{��΀8{bBj�I���,��F,���в�9�� 8�*��Vhд�u�J+B�6��aRng�ӑ�s��5�͐)�cvM&�s�tGb��
4bZXA�
�l�-��biD��v9�[�66��*��^��Z�ɴn���z�-���!��ԍ4���<��> 3d�=�����)��5�
�,@YcF�*��i��(/:�VL[�;nScn�v�]��Pv�xm�諷R��>_e�(��+a:�	�V"ºF�hY��5].�Rb2�c٦�6
��K4�CB2^ٍ�1shaG����h��tq덈���Nn�n��6;���^���ʔc����m,w3R�`eXPL��i��t΂�6����,��{v������ԉ���Q�fn�Q	�ii��ٱV�c����vx4p��@�{z���Ƶ��r�����jB�9��ŭ�a��Goy�ȃ���VPMtn7q��1�.�΋45ĩJP(�N�T�ɢ��R�ˎ�o;5[�R���bÉ�9��qG>�d��E�GAz͘�i�h����0r�κYd��hhҘy�5�LiIaf,j��][LSMCNN|��y[������,q¥M�	�mo\<���y����@�ru�pc�&�Q��V�.��f[Y;ixtv���e���ˌK6��1��D6��j����n�GH�K�s�-��{�]���^Q�B��eu�G"�A{X� k6��b�.+�琳�| �PSQ2ݛ�cԬ�H]�Z�#��[�K�1���Z��V���ke\N�n����|��/�v��9��7���Sl�7�f�ú�����=�sv�!��Lh{^9�x`�m�^��%����뗗g:Z�]���u\�1���U�Xb�
Lc���&���eb���).-�X�琞%�܊6P��L�\Dfh���lAх��a�%�5ɚ̪I�t�9���n���f��3[�i6ƹ%:����C�k�vԘ�n�f���Λ[
J���D���[��9�^g��=��wJs���x�E��\Fi�K��m�JM�<�Ƶ\b�(B0�S���R$t^z2��e糮K��N�х6x��V��闵I��V�6%��C��e��� ���*�GCfh�J��U�2�f��ֲ����YG�� �Mӓ��]v�3�P���m���Բ�%�- ���h�SM�(m2�۩a����6��͢H�c�W�u���b�I4ջCs���י� 	5-ִ���V_K�)�8�+g�P4&��� 	���MͰ5c��� ��]�:hR-]����]a�,e�"�F69.��p�EV��z6S�&Zj���G�a1��9:�K8��{^�8H^ ���u�xv'��'*��Κ"	V65|w���M��]X=N�1�Y�:Ʒ�+�%��ۮd�B&���M�#�e�.��4�m	Y�����{غ���˸/1�-t�yٸ|����ۥ�s
E�74�`,�42�:�Q�KO)w�4HK
8��oC #����:|'1��B�k]�Վ��WE�c91m��%��cKV�T��#�6mofC\d�I���! ;gV`+��:�8�q�R�w�}N��1bXj��Rփk���I�`Ŗ�ձ;>fV��F�7n�X@�6:�Mv��xN���=+'^�.�='�C�9-$�v�pY��jQ��N�6����WVG`�jFf9B̭��,�{1�& I��b�MwP��	ڼ�۱���Ouת�P��q8�{S�d`ɩ��'��w�Z�Mcq÷iKbZM.,�6� $�Z̷c�u�s�[\�j'H�<q��è4���&��pK�e] �fB�n�Zy�v�Ϟ�n���W	CO=���m�K:5���S�W8T�ܽv�sp��]qu��]6�ӭ�nKX�;m�vһU��;�8��㬐!�9Hr"(�ܹ,іB�n��r�M�΃���Zv֋�Fݸ]�'�jkJwnGA�p��#78�&�J�<�E;�]�,�[�9�W�\J��D�8۱y[e;:�Ge�.I�)�É8'A���V�s�P̔�����"�n��t�P\疜�쳷"�)��gY�w6��<�&b�3L��S��p^Vv�$����9Յ��qIm��Xٻ�mv�9ȓ��r[��yہ��zN�{kl��%�l�,�ŵ�,�zd�k�!N�D���q ��-$X��r�NGN�Np��N����kZT�!:r�Rx�b{ZS�I*t��pP��]��J$!��D��,�/D$�H�6�XN�r%��ޭ�v���G�K�������gZ�Y�Q$�e��D8��RH�|��M�5+̲�޻E�u<��I�&�(��t�z�u�ݺ�3��pu��p���n]�ٓ������Eư]�u�<��IM��Em�Wex�87����,���D=rZ�kG[<�6Eh��Q.�7n�^�0r:�y��4��xz���#�l�Kf;h1`��!-�l&ȝuJK���&2�; #bV"�k��7%s!j��&9�͝�l �ff�/(�wl1�ᓝ�����n#\�<Z�7]\GlzL�u#�±'p�dٝ�.�������{�hǖ�蠻c&6雍�=N{M1�'�vK$\����/d�$bN�<n���l��>N
��ݭ�v�H���^L��s�Þ#�,�Җ�%CR����2*�'i۶z��M�7�S�L;�&�"�0zm�C��rζ�6���Bګ^ų����8��j��X��s����8����x�iN�J�������Ģ��Jm���٣O%���b���1�<�g�I�ͭ,��'��\�W%�%\�vlb�4������L��ƃ�]�5��{���>3V$BV�2��64�F]lp��AS:�#ڙc,,8��!�>�l)��#�u�M/����etIe�4s�)Yt�D �mR���[t]�n�j��7f0�ԐPK�T!�鍴����	6�bX��12�5�p=K4�iF������ӑ�"z5��=�ج�aNvS��V�w9h�M��HZ�h���d��vwT�<�VM7n��yHk*yn��*�6���$m��SƬ ��[ n��r�YB���km��H���k�]�Mj1����Z����8#�o@���
�6�-Ny6MM��Q:Ǝ�nwn�Rb8RC���3>�<4+_+��HkT�lر�
Jk�u�� �$f�z�.���s����9�!�ٮ.��ck�nbF����g2t9���G����"a�JF�fj���]oi��i�l���H��XV�l�W�+-:дF�T��Q����Q����j���i)*BĶ��j�%�Ѳ�̱k
X�5b1 Kl�J�-cZŴkT��G�o[,[+HT��[i,�4`Tb�S��`�H1!�k-X���-��2^�-���ŬV��k"���F��k�db=��g������4�8駳]��=V��s�����š�.d�&�$m��C����7�2��i�N�y1؝.�K������_���H,�8C�a�d�A�!��L�&�������1�G��ϲ8�-WY�+
�Rr���pWjr�(����}ҀBH� �H�/$���P~���=��ŵ�f<x�b#�6�.�WUܒ��Y�f}Q�O[��<Ls�@G9� �M_Os7�7��gTq[�g� �PD�*U��J�;9N� =���,�#�)� �"I����z�z��D׻d+ǰ�)���:�aQ�|�_:G�}%Y��Y�G�qӚ���;���i��8�2��<���w:[�hV#��2�YT��@��Aӹ�d�"D6���A��jz�x�^�d����;���"Na�~�d���&ӛ�4Tc��P����ж���zqv�8����[V�B��W�j�^|ԋz�U�V��1cE�v�ʻ�6�����4(j��#a��������f�&�;l�KP�t"�(v,A2�l�1���H�#=�a�}+�(YF�"D	xR�Ҩo��\�%]a�XTj�8�u�j�L���J`�-Zь/e�*uP�����&�������/�(ڏ.N�F9��7�����`�5��PFJD��/�����aG����
Z�ٞ�<��m�Q�j���T �b	��(Jʙ3o�=��4A�A�_&J�e��3�U�	WMa��W7Bb=r�X5}������3�=� D����!����;ݳ��9\�}^��u��ݗ ����~�&A5B ���Mח�+Q��l��V�d����/�(ڏ.LX�F9�� ��^#Y]�O�rA�K�'&DhT>�$ֺy���@����9���{���|N^�������2�"7a�zw�Ǻ���k��uZ�ٝuUf�TKHޖE*nݧ���d�2v^��{��g��g�7�3% D�"H���<)��X{���s�ޡPv/�	�^�}ԑMqWYEV����u~��JV���A���� �2P@�$a�&ad_	�޼����J��l���n�T|~��`��|���L�$B۬�����@��g��7Rk)Mp��c,�Yf�H쒹��k�V�b��EMP��>�e�����e�~<L�G��W��ϲ{�ZuG%�N��6�n6�H^���.9�z M
�I��2R����乊�ֻc���#bv��(��+��k
�R��_:��
�hm�ɵ�^��a���"��� �F���":�N����'��݇.{�z�����)��Ie�Ҥ��]��ֹe8o������s�#�I�����	�έ:���'d?Ar��`9���2��˺g׻X�c�Ṱ��C�-��V�ܘ7^Z�;�^'������:0�����*U�Q�;ӗ��q���/V�/�X񽯔��I%" ��n
G2���3�*vI\���+���
�R�G��׬5B����x���Ct�o%E+$�����Oa��l�2&�\�#��ulmUK�̠GU�h��T���,� ���� �Ž'��f58�������iy^Ε`��b��o�.U�.$��i������(~Ȕ׸�Gv=�Mnui�җ!:��^���\;�%dUF�%�r���گ':2 $���Ȅܓ��F�Ԓo�9ruܮq}^�ߓ ��FJDd��D�����T���\ww��|A��TЀL���KO�x����`��c�L���8�s9�Jf^R�̹Wq�cw"`�$A+o���Z��A�N�{'d&�'���H�:�D P��\5�	��C t�Ćx��G�����*�2.ؖ�[W�_#�?<�/�1Ԛ��\�EneǨ�v��Q�����r�B*��/��ٰD!�O1�Ι��c�t����]�&�Q:�t�i\�[ �j@k:F<�3u���3e.�^ڋ,�@��9-��B�[���b�z�1#��۳pJ��8���ɰ\B&�Bku*.aT�;[y��G�]����n.η]�+{.�̖�1=)8lvsY{�����-�,u&�>{&dWh:�H����nrtY����������2X�k���5�sJ��x���Xy7�v����UEE)W}���\H�^I#.�Ut;�N���*W��QjX7�&{s����=( wԁ�H�"E��J���%d���v��SP!*�̴�t�}�Ê�&/��
�P	*��[s����7�D�����2Et��]g�' ��=�WJE	�(D"�@��0d��DD��2���^Vug���z�b�&�wk�(��)\Z3�E���:�ʉ���و�N��܉Lc���$J�?����vo�����V`�'Ci��}�KVgt@�X��t�=�	& ����k��U��lx�US͹���C�e���a�N�m'F��l/P�nuǍ�urd)2���rd� ���쉍��]��ܞ�+�"��6��c�D��a�u A �#��d��"�^���f�{Wn��S�o�ϳ+�deӣ̴,J��\��<��l�0n!�Le͓r^�b��2�V헻"Jwq	��h�[c�?y�������5�ǹ�Ҳq}^���/��܂2R��D�yw96�~�W�JcWwE��*�F���{��p���u4�Wf���)���g��	&?������Vs�=V]���9O�A&�;�^�����])'�\��{�.���z��	�@�T�I�d�2 �GK�oc�!�P���n�V�sɞ��+��4��.z�0G����H�d��8�֪e����LE�NӸ�{hc�6�e�CXE��;�h�Vf�a�
 ������9(�w0���"J�)���d��)����y��q;��.�E��v���Ⱦ��A�>/\3xR��˳4h7t� �&6�qY	���Z�R(O: �f��	��,|��ǈ GH�IH�("$���d6α������l���Kri�K�{�$RW��Sen(Bc͉]8+�k����i�yY��J�^aD_XN���WqKEE!��]%�Yf�zs��<{������� �鉐}� d� MX�hP��+�ܦ{(r��_���M
7���<��S� 5s��h@�/�gC#w���7��U�A2D�B��-cc��"�Iڰ�vBor{��L��O3���=�� �H�"
��e֩:��ƍ
��h2�m�,u�b�9L+aE�](@5����7F1�p�_���~z��4 BT(@$ׯ�Яvs�<��id.��E�Eg��1�fn�khW�'4 $L"@�%E��u��_@J��I��e���Ru1bb�%# z6�(�n��rR9Tߞ��3��$��@&�L�#�I�t�=��LξYBg��Z���tP��D' W�6.	�R��F]�"�ݝ+�_&a�A訶V�^�ӿ�2(v#<yW0��=�J�S����Ȉ���vI��U�E	gʍ�z�ޥ۶4���z����ν��'�pJ�9�T�ƅM�+{V�ײ�F����M��o���
�l�x��Smg�X��d�w*F;�]��w���!K�,��|�^��R4�X��(fd˻�I�ɱ�;&��.#�ܹ���ރl1�!fY����:�g��s�$�Kv[uU
%�m}�w��G�d�"ӻ��	���tP��Y"���1��Gz��uaPDI�H���r��9Rs���~�G*��q�Z�+V*/��_�?�>����GY2g����L7P@��D��H%ch���ҋ�F�V��R4�_�UX�	P� $�֒�p��Gd�~�T��n��ňNjBJ�;���䢷L�P�T�������3z��	-��w&?w �#��d�9ə�������yr�c��U{F�~�mU�mP�{�A��3��j�w�}������(:nf��=��஗�d`;/�����ljޡ5Z��O�a����g3����禍E;&(�H���M�AyR���������#c��cIi���C�����sv��1u������d�xw5�3��Vۉ��i�����k!Ν�y�6��eyN��������"�� �A����G>;�>�um���۠�рV�܂Q�������k����{m���k&ֆ�j���ZRWb��wl:Ν�I�EY����Qx.��qͫ�u#4�z�����­f�ͻ�\���aB.��;���j&��6��4-��f,��T7��fn�C��T�$�'������yB@f���܂bj&���P9����y%W8�\A][:��^� G%V:{����En�+��T'"�mX�IT�b.�^S/GOe�#+��Cw�41�Hfgi5��q�k��[#V��f��KU������Cf�<�R�fM33(��H�f�͗)�H�^���U��gU�����O0No&B:�-~�SS~�����[�`BSBBJ�i+!)�$�Ւ}Y���Z���J֍%ji�ȡV.U`@JF�Z���=n���� &z�T��a��%�.�V�dY�<K��l�jFJKUN�(��+��P�6�R�������(/OT�9��W�Tb���ل��Wuи.hG�UpWb=	H��*��p?=CC�c���w0gs��]�Q�[�u�9��/2���Z�lZ���/r��@�Ȩ�ɷn�KQ�
Rg�y�6�wc�H� �A)��Oz_�y�Z��/M#yU��P]35<�=/eo=�(��{�C��S̉��d����¬J�/��8�ĭh�V������,a��P�2i��JffU��s��8��(O������7sv=��;=3]�����{{�M��#��X1�k�#�[�T.�BJ��J�<�G;�����ٌ��4����K�nn�����`�;�ݏ���W�·+*��������CI����xk��v��v�$\��Uj5ٹ����A%M2;���>g��^l��d��%W���tCo�%�4��V�a���2�.̐-�_�u�����IU�
3 p��L$��Df������n���;�{F)p"-���Ջ��qc��y{jW}�<=�$c32�y�41��o�sz��r�t�yu.�h�*ˎ��F:�kv�e���@�L�;l>�t/T�?P��Q��w�x�4:�������rϕ๣���p0ZF����L
���U�x�5,n����uN�����i��{�\��S�Ӡ�+U}���0>%��=���V�>y%��7v��n�&���ڂsr������#6#{3�M�S�O�w\32�4z۫��W�A2�n�B�(��Ek��"�Yኗr���#u��s�7R���	�@����y��!4�Vwjʮ��u�9�x�vC��t�56Y��A�Z�[��Rȁn������f�+d68g^����2�OK��N��u�8r���|���2��6Ԣ���C�m��y�:<P�W��l��U��Or�<,Wt�f�Y�Y�Ԃ/ZuRt燥�߶l��v�����c��V[����^�/��ҫ$3�j�D:�?hY�d�ή���Gj}�0��ٮ�{/�C8�>�wY�w(7z��e����yf�W�.��T��%�$���޾{��|b�Y���Y���p1K��$q�Εj8%@�7sfJ"3,�
���j�s7����Ӫ��]U>�
[�a��Ių�Q.[˺�gSOf�p_=�B-Ǧ��mkzݳ�U1�r���RwV��w���l暀�>�~�Hj������3e�6F��UK��W[t��,�C��sM�ɒ��؂t���;���;��66�ֈGǑ�%�n2k�d�WY!��(��3���ӮA��V��.���Mg���\�V�s�(yB��z��!�ks!�e6o7z������v�:��
E=���rvd�
D�:m���% @����e`���m��6�t'�!�s���@�� ���8$�"���rBVډ�%��8G�Z����@R�@�"G!;9gkm�� �miH��9.H'vJP�$tS1RQքYgJ";�$\R;�B�/:����is��:'S�J�c79@JP�f� tRE��ć"9;�s��$s��"I8(��N�ȑNq#�]���ܜ�Ybps��%l��C���qI
\q�N!*J%$D)˔9$�Nps�j��I'�y;�����{��y?��&=����������"����K���JjBJ��o����If�%b��!�m���wd��[� |��[�JffQCO3&�<�%337�����ч��4SV/��ޞ,�]�|��4�vikw(��
G���N��ᬝG6�8��Gh��wS���od�B��;#t���D��T��P0AΠ� ��0{��@��	�-2�(���EB��WH�.Q�mW�*���	+	M!%W�0���Β:5M@�)WvW9���Inƒ�
��D7"��B����5����&�nuR�l�Ƴ$�feR�T1�9�'��kU����;�{F)b���CjŁ	M@�	*�%B32/���b�܌ sv.up#�*[����{�z�Os�_���/S�<��r���U�fŋ��)<y�ӧ1�![I纈�Hԭb�;ғ޺9,���Y�'ٺ'�P�����l>زQ��ғ��)�D�i�d���S̎���E�e����ը�V��;�z���Gr�$_I_>ջ����g���;ui����p͜y�aǜ�u��������0�J�.�7�ny���ɐ}�#��~���u�x�'�<y�]l���	.wj{�V:�~jt@�	*�	+��A�Ni���,�\�ӏ��I��I=�i6q��v�! /M���
��/�=��$Fn��0�ͤA=�O�%b�)��J��v��i��َ/����o0��(ov	c36�y�*�$��̥F��wY݇�SU� � Z�jJ��&�n��^uV�Q�|�۫�d�9��JF�۹���_N�L;��OuGw �w$�RMݖ{=���h%&�����3{�fv�P߻��̒Y��I��Dļ�7����Þ2�l:o!�,J�싼T�]qV�@��W �m�7�Q˕w�2wp�6�C�7a�<6���I��]~�$I(���)��e�R&�@�v�۔��
��ڻlQ��Ẏ��I=�n�Z�����]-Pkb�v�rFJ&�Y^y1�}�&��D�m�mz�.5�[n7<Gmj�C]a����4�+�ܼí��t�-��Т]��#s�q�%��[b]`w�K���
�`���[��F�8=���p�<�zG�юʹ@�{[`�FՕqqi����-�4�K�P�l���6uA��\M�{i�1t�]���!n����{�؁%~Jw� IWvu��mv�vIW�\�bx%(*t�sU�?P�b��y2�@wv=ܘ!}R^�T�����t[�����:Nr�ct�ꭂ�25�ݚ=ܢ��8��;Y�S�T���ҡ��%�3(��d�d��N�s"|2�n^�_��=p7���ɑ* $��	+�S��Z��힨o*�Fs�p�ׄ����}0��)n쒱���ȯG�Q�f͂�$k�G��@@IX���X��������H�#"��-]���f��;JΪ�*1K E�W���%:#�*�j��݆.��SB��v����ۺ+5�E�cB�q��&�knG0ݷ�ÍuL�U����A �f��2hcX�Uf�q7�7�zP����cv����{ڕ��5�$�ٴ�33(����g&BYW]=��n����@�ﰍݏ ���q�'��Շ)���7j_C���[1�ˡk��n���%��a`�uH���T��q�����~���HA_}W�ݝ��l�+wd��e�7"�G�L3��S��Y�:����l����	P�%^����mD͸�硦���gUl�ǭ:�V,Jh��ɑ��0it��D���<���1bUp!* ��/v�w��v	����R�T)z��f��������{�2���uja��F�9aV��s���l�8�h�he�����P��~K��@�A-�3�)}�7��T�@$(���Y�8z�M�O=9�x{�B��h �&֑]4�1��<���&�LD�#������[���=gg^�fq����|zk�RXj�Mp ޛMz<��W~JE�+-�
%�z�ך�7y�
���oJ*�A��܂����'ҡ_]�3��HL�^������y%F�C����<�b����]�[8���n�ߘ�(%���F�!EACs�,HM�WF��Y꼙�[��j[l��k[�܈Y3���}���T�L�8�t�He�޿7"���IMa�?�m�!�l��0��W��Gn3ݟ��m}r�`q2��fD����ٻ�LCbF��)�l�9��{y߸�u����!��ı�l>��ߤ
a�1C�'��/�߻ٟ���1�l^a��iSP�6&C3�)��p�6�ݔS؎D ݉b����76����J7vQL>����YG'����z��!��h�b���En���������}9x���l�C��҆���e���Ch#vi�m��ݐ9�؆���8�6es���ǿg���n�eu���͠�k��%f�]��sZ����Fx�����#@����Z��Cb;�)�lCh�}�#�Cb�h7bZT�1��۠ǀä�}3��'f�����W�C��!���}�r��=�AW�7Ƃ��>ݠ8�6�4���eÌP�6�7b���@�Cf��pq�lCh��E08�bA4{}������Q�}�bA�8b9��.@��73�b8���3����~�}�;π�����iC�C3�} S&(bG�l������nĴ�1��{<���؆��C;ې)���m��>1����K؆�6Q����6�ݔS؆��������RQ�KŒ�F���_wZ�x|��6s� S�_P�w���Ch#vi�m8b7v@��lCp0��G��0!�݉j�J�ý�C�Fe_�V*f��1�mw6��!��͉ixj�����۠ǀ�N��?|��3IT�����lD>�%�n�b-dN���}Q���V}*�g �����8o��ʚ���Eկڽǟ���������7�x��S^��.�'�j���;#��#�̯Gbx��5�����I	���Ck�J=J)���l >��b؆�ݐ)�m/5�(�!�mn�1��Cf��1�>v2�s-�C�؆�}y(����;�}������Ͻ1�y��wbZ��CaP�}�L8�Ch���q�lCh7bZ^j��6n�Mms��'��?_;G4v��p\�ۊ�"Z�:����b;Y���UTSk�J�)�o�Ζ���O��gKbA�b؆�ݠ8�6�(h��E1�l8ѻ�6��}�g�V�r��U�<5�l�nC��Һ�����|��h��QLCbA���bAN���d��m�(�!��ؖ�hC��*hE_9߮~��zy���B�	h�}(

�}����}���>v�'�	���h7`�!�{HE&3%��'�$��1���	M�.B�����SB̐D�3$
hCa����7/}W�	W�.:�P�8��`�� � |#�޿��T4!��Ѐ̄%��(
L3$)�����n{����/��[����`љ ��ݫݭ�'���3>@s�!�B���P�R�1���7ܰFB�l�CB�ْ 3 :4!�32ASB���SB̀>��>~���yV�ta\�(��m�����1��y? OnP/�A� �hF�JC����cFd =��d_:_��]72p�����V���2q���S.���>{�[�;|�un����=�WBK��O�.����U���y�P����M�X��]e㮁���+6o6�%	n�9D�E	\���1����1͖�Ji`JZ�H�J-"v�ֺY�ڶZ��,b�<g��e{V�ҙ0�q�Tҙ��`�b�Z�Xmp�tv9�v�<uwb�\F�n��8TX�i�U��aFhf�;[��fua,19��S�NE|T����Dr3;2�(��R�<��)+4������ �ï.t%�M���Z�]�[���E۷�r�R�ʵr��Iޙ?�ӥ�Cٲ�I�ݐD�,̔%L32P�����~�>Ꝃ��\����4���>����_&AkB�ԄSB�������32B���#B||Ne��6���#��{�J
!�f@Uz��x�U��I �� a��G��OԅCB�(3$
�r�~��!�����Ж�Ҁ(��B)�f@4!��(�9{ȿsO��mw"}����>��'�	��|І�n� �w)��^d���,� ���!I�����;�ϣ���e
��_�#B�~�(hCL32P���������ި��݀��*ߤ&�I��q�W��; KB͔&��4!�d����B)���A��G�b$xg� )5־x�U��I ��{�	]�(TІn�"ZfJ��3%�gٹs�94{Il��̲d��p�v�f�f�mrIW �m4�6�a*&���.���Cu�.�B��M��B)4,�Z�����{�dO�_��s{w����>M���ݳ�dDV u ������L����i�2fHthCfJ4#=�ڽ����{ن�h�����y��I{e���$rItz����e�2��zc�ޛ�V���J}�ss���"g6�<�$u���_�$���߽ ~4!�7~�W/������|��܎�ϐ����J ���B)�f@�gk,9ʻB<������3vP*�@�2��`�2PS@�H D�L.�96.E���cR��RH!����BW{(T4#v4,̐)4!�32P��4!�����}ѻ�;���Ͼ�� u�Y�(
�������}��c�n�~ �܇�cA����>>�99~�s�@͔6�� ��32P*�(T��3$#����Z�������'���+}��7=���v�`Vl���}��CB̀%�a������N�w�����?��mm�v"��^�y1�6]��8Viϕ��]1*�lj��G�Ǥ�zd�Ќܔ"�3%6�� ����7y�Fr�������>hC>3���3,W�@w�`Ю�@��0��@P��4!�3$�9���ۿDj�hW�)�0-W��{���+���[j7I�� V����4�
F�=ݤ"�����*�������*� onC�B��B�Ї� �����32P���oQ?�\�
ʕ2�{��t�m����u�Ѭ|�X�����ᅾO���8Ԯ�)R��b�X�u�*�J�ڡ��]��3K��yW=�VG8]�$��6{�ۭ����s��]����B�d&�?��B(hY��c̔ ��@���d�%�O��8�q� ���R@�]�()�Fd I=�ϳw��_/ޜ�|��!�B���B����l��}S�G>�Ml>��@P��4!�fH*�2�d?w��j�ev2~�/P�0��(
�������������|=���h7a N�� ��A�Fd z)�4ˇ������-|�2�)
%����.�up��竻=�s���.��2-�s���޾2^�1����H"A�fd�*L32P�.�w����ۂ������ٲ��s ٩CB��HE4/� ��Y�(
`�!Mmd 	�[����{�@��֏� $����ͣ�W�Ng�>@sޔ�w��M{���fd��y��@��a��@�036ARhC32��M2 ��J� ľRv2�c.��7��җ�y^}�[π'���hCh3`�f��C����m�#@fd�_wﰺ�I{|���zP�Ý�D�-ߤ
��(
��}N��}���s��>@w`>hCL
Ϥ4#o�xw_�4����o�I�6E���'�����)�����]2zV//��ÿ���[R����=�[��Br�	��̜!�s������K���#Z�@4!���P0̐���̀R4#3% fd������L��<�r`��}���_?�W�Ng������`]�
7d-3$
��(
������������ؗ4Ɇ3;M4+�#T�١�gvr�Ù�fZYw���>@_`-���􂡡��B)�f@�,̔w�>�����^W�s���	�>ϻ��7�$�ǈ�
Ƅ;�ԄS�l���4fB ��@����B��v�g՛��j{�V�8
�$
hCa�d�*�����}��ڬ�;N��v�1�Y��
_}� 3 ��~����@q�_nB���-��B)���AM̀GL����Re�+��e��K�G� gu��!���*��KB����fd�(h�	Mw��ϟџg9�F\��Ї��B)�}����@O{�~y���^W�s��@'���̀RЉ��z��������s�((`�4n� ����6fJ4!�H"ZfH٣��D�;@���������wݪ�s��5݀�i�Y�І}��M2 ��a���τ����ݫC�#�)h9�"Zs��X0�E��h�\s6ɒ��T�t���U�t
�,��*����-Jt/���:��x�fU���A�V���1Z�]�ӽu��m�L=��]�2��E�䬳�7��O�j�8����@�U��"�[�mVeV�˪�{�#=�kc�x���U�)^Q��ԕ��d������"�Yn�wZ�jvnU�Vvչ8^�34��6��XJr�2�]fs����cgu��.��vZ��]��wݳ���e���Y���f�jMm����7x�&��=�>��+��e�ws��X1��<.�z�	t =ȫ�.�^����P��o^����T2�����O���K":�,�e�z��^o)�<��v$ܼ@���U�v�I�Hb)��ܳ���vԼ�Xped��-���S�`۬�5�;C���v����m�,��Z���ׁ(����������5�]�yx�#��hwl̷�$��1]��+�a�U,�bu*2��5B��f�\.�Bn
���ZY����0O�q^vs8��&��I�͵k>H9Q,e�ϻON����ۭ�9&�qݷ*����2��m�8or������+�z���֊�V��5��UY��W�0�.uօ��F7EqI�<!4��y	���5|�U5λ��CWT���TN�!V��b����ۜ���/�s��}���C3E���7�Z%ejFn��Wpd�<�w^�4����4�pR\~5a��w^��N�,�h�����\vE���X�e��$NC��nG"��ֱ�-9���QΉ��99ܤ���H�Y	���"���9؈H�@smJ� %,Έ �t�֐;ڳ��q'D�l�N�:���� BDQ9�"
�rp[bQ�9�*��H�A.���n��Nq���s����!ܼ�9N G!$rq�8t�q9�l�(��*8D��$Y�l	8��J���ItT�C�؍!�v�;�%����7h��v�"N�、�@�$#�p��h�g��_m�������v��
l�f�Nc ƙ8��v�v��'���u\-�'\m��vA�)�	B �;.�\�����3so@q#�ng9�z��#u�=��L��h�NCCH��������a��8��w�nX�ݛ���+��X+��r����s����_.&/jf�X��%��u��jBŞ�0�<P�n�c�\��XB�F�ݠ+3��Ĭ@�@�\�ڮu,�4Tx#������#2�4�,�&K0c��;b�Ո��X���V��ͺ�O��u)�d��)/OWaa��|��S&�F�t�ڣn����|�z��A���x���i'Q��i���8e!��"[I�ƍ܂˝��t���V��4�lGuf���m%��&<M�&CԽ�.�2�m[͗�l;M�(��)0R��0�=)<宼�C�����5�m��]����3�.|��5Xd�窬]�||'���X�p��^5;�z;-͸x��#��usm��������V�/r�W\U�R+�����36��d��8{����կgu��x-������ːn�v�z0XRK;��Yr������z��rE�93qp�<q��[t���ւ�i�9�ݍ�Q�}�:�m�����jL�!qu�:A��&8X3�]p�	�m�h�[vN�m�b���S`���h�K�S��J�7���B����s�NL��;Q��P�+� M,�d�`�� �����(�6�UϦN0s�o]�*�CL��p6����h�tVE�i4�`����֋�U��&v�F�����ûs۰��`é�IQd�r#�ɠ��G]I��
��;��ۯ������2���Ԋ�og�g��rqIo:�H�df�1�{�d��1-�۶�c����jN@�sk�f���8u��K7$d��[L�	�+[�s�r�co]�cX��4�-%й�m�!(3����ǌ�;���:J�D�t4/z��'�����%�u�E5O��{������u��7N;a�øSPը��:�.*76lXe� v1�6��Z�\i�݃�#��Y�ָK4��e��#�#65�v�����U�\ v��v���4��c4&���i2�(����e0�]\Y-��cLM��,�Xznշ)��M��$��t9�K����B��.���t3f�Z3v^����f�Y���)[������C[Lή1a+4����q/8�%�؎;:���ɻ���Kq9[�3�V��ED�W�yR��6��Lϩ����AL�Fd L��켟������g�����z��GxFw��1�zeZ��(�l�.���@P��І��(����6j;ʞ��E{ HІ��e=��>�}�����O}(�A�@)���P�fd���~��t�#�} 4��4%���R�$(hY� P�,̔*���Gi��գܟm��ۂ��\����CB>�e��f@І0��@P�32B�sU�Nn9�A܄a�m!�]젦m�{�y�|�3��f{�}���1�w��I�ף�q��#>f���,hCa�d�(h�	M	fd���33)��� oӼtF��g���"z�(	�p�}��������	�>�ϡ N��C����h̀ܟO=�ʯ������@։�.қ��Jm,l�3��t��WR*RRX���胳Jm����?�N��=��B��3vPfH���������}�Xw7 �� �>�D;��]9 _����RMr���fJ�fHSBh3! s�Ȏ�b8�1�����r#��ch!x!�A��Kd�T<���:��UY�J.��
6����2��b�Y}�4N�1��~�s*%�W�� {��B?.��
`�� A�������3��gs!����_0.�P�4#vг2@�y_O�a��@P��	��M��B)�f@4!��(���"B��9��]���զ�[�ޏ	�ϡ N��LfJ
`��)�32B�Bv�;�y�����ސD����4!�32Pw{�~��{}�z�5݀���H*hE���_�I쭸�B8Я`	hCL.�PfHxhCh3 �B��B)���Aɸ���Ѿ�	���+�|�{�jSx����z*�nRH	 T�Y�D
�,�6A"��?\��O<-�A�]\�d�a���:.&��M��Kn�����h�2&s-���Z�[:t�wU�)w�m��U� L�h�C��)�sw�&�+������ۛ�V'�J�T	ݽ�;�����>l��ג�X�I����J�t�,O	��EI�X&1�8mR�x˾87�<�W��r�@T�m��s�㾕B�}=f�M
{�ӻ��� �mPmN�RԦ/w�;�y"Nxh�]����S���L�k3�k�����L)�`�չ�z�3�X��%	"H��$���T��E#�n&�s�wvJ��IPmW��I�LnwIO7���y�!�6�K�?�W��Mˡ��C*��hײ�I�U�:*���[���RD	��ˋ��-L^��u���M�.�T�* �Nx�V-����ƪ�";�S��ՙ�ė��N��0Tg0��x�{�Q��o[�ʮ�zE䁏+��	�M I6w�R7�Y�(m��s�wvR��%A�D���&�r��=�56��m.T<L�������X����Dg>��k(�=>[yv��B�Ж�*�{��Q���wpGa^VP�:���N�A��tt]���eQC��S�lK���R۵�*�4�}��x��ANzH���0~�VɆK�:�S&J���>�S�`��`>IQ&��w1t�uYߚ�9��Պ��]i�Z��gW����s��G�-'D�����}٨N�I+�74b�����T�$�uҝ�ٚU^�@'>$�&�2\�]�]�����ȑ�ڋ��=޵�L^k�4�Iǎ����!��4�d���$�&A�ڵU��@�뛹m��o�av*w��r�$�ω5�bb6�*�J���T&�v�#i���������QG���Gk��� ;'�*$ׁ$�N��z�:��"BYͩ�;�}܋���v.�D>���5I]l��k��#`��wX4����]�ko����Q�cx
��E��7�3Nlg���<�r^<��D�<��k�1��}�{�HH$��7$�]7T��SR�]OW��˸ݴ��*u���$�M��5lgt��p�U�g����W��ų׳ή�#BmN�c��.1q���[�U:����;k5��4%���A�vs\ы�m�*���;���k7A�.{[��:�?ŝ��~+J1u!�144Jhb����k]H6^{B��0W�i���B�B[�#����˥�i�|��,��cp��mav��"Cf� #�ˑlU�9)�b]'��)f;~���O����$�=�Ru�}��S����ݚط�?��`6�{ ���IՉy�9:4�Ἢ�i&5�{}�ۺ�j~]�7YRb�\ ��wh[T\�Mk����^��5Q>�\�H�޻IT^���4R	4	4	�y�LB�u4���t�'b}�^&;ev*w�.@4���ƫE,���dk�$׉�v$���=��8��>���m���v굩�tf�3�K�����csL��,i
��UE�Lq�,�-(��rR���I�SM�T)�MRT�gWý�I!�Yr9�;�i*��oX�f�qo����E%I�U�rZ������ڞ
���"�3�T�Z$�~�S�s���!]T����ٞ��hr/�q��E�&��W���28Tn�ӛ9��V��x���>���ꓯ���;̹�H�uX�-�T���y�Γ>$�'w޻�rU�u�yٹ���j~]�dMj�A�g��=�r�����e���M��/ww��#^��yhVV�hׇI$�hH�P-�����#��ּ���Vo�����Hٳ��F�3��v���WiAЬ����1V{��&7=��x���d��j��E�,φH�$�� �� �v��mgn,Z��(��t���GZ.A&�I�3~��y��htL�����*败�~�h�Q0�b,9z�sFd�u�Mx��%jC���wr��k6����r��\�C��oDKre�H�YD]4���.7^���+s��EIF���9�.k�Y~)���OWbb�I^����(�0����VhI8H�%���'p�o=�MS'�F�x�'s��LQuy��^�i�y�=y>|h�@� �D��6�"q),��s���wW��}�uI�gr��N5�%T+ONXKSE٥��M�B]�%�\뙢��:.5��E�B��{���y	+契_z�{��ޞG�)<�Ȭ�x�@B����z2I�hQ�	���������B��=�汛�Z�j`۠*&/Y��#37iy;���$�L��++��i��	���u&��%(vn���I�8�xۯv��R	5/^W-�����I
O?u�ѕ3��f�v����[��ca���(���혹Qݡ���v:�5j�|�:�	Ec������e���u��ڼ��Q�ޯZ�����~����W�r	4	4	�KZ>8�n�/8�]S���ׯ5���KS6�Ux�I��k���}{�\��HRl��)�$�fb�R���l��`*�nV9��;�T���##K�I�	���Ҝ��P�R��a�!mE����������f�I�L�h:4�\]�T�J��o6G�:��r�k�G.$*<��}�S1D�������u�I9�I��8GP��9d��[�n���Y�j`۠U�dhZ�X�1vg��,�����iu
 s_��Pj�כt�.5�g��^$��i�T��`�A�P��oR;����㤅G���`$�����F���3ׯַ�4��n!S��:������ڙ�T�>��&�\~�(�����[M�3*��V��'&^aW�+��>I!!Y���A%�>�1�ĻCh\b�fv.1�Ƿf�*����D]t�z�;V�ѡx�Xma�4���]���`�R�ca��3��8�!�%�L۬%��P
�qc9���4��t���s��z�q�(Q��&�E�t�hlű�eۧBnm�-�I�fl桖�ju.����'
\��t2�	X�s��͎�-h���]�K5R2�X��������9nԓn�;7;Zʾ�j�(��ev:�dy�s�ňBf���N���&�I�G��ׯ_Fnuf%���w���ڮ�rt	�I'|L��w	e*��n��o'/Ս��@�kP	r�����
������`f�$�I@I<��0iU�{-��U�xwJǱ��I
�?r9*�&��&�Giv6�:�V�jD���x��z�t��e�Z�6���F"�#&,�#��/��I_I�b�!yL����:���X��
@汇�%>�kĕ��D>����\��X��uE�A���V4�+\�%v�n�,�1Q��T�  [��"��;�}�$���+��gsǱ��x�g��r#%���U�z�{�I'<I��Zm�9NeD�)���Q�b���4>�����pvN�&�*�f_�<�j�,�g*�{;UkG|�g�,����o9t��0��  ��~��^��?��vs�k�r���.L
.�e�&�<�3�1�G������W���$ׁ:V��ӹ����ATm��[��KlP)3�\�u$@I��
�+tг-�N����r&���ج��zGi�����y�v�H�&�$���K��| -�����ǭ��^�^%��tˢdow$��[4�=��Y��`t��xzz�-�Y�](�AK� ��ν��8�n&�j����H�� ���D�Kԫb�HYֈːff�񎹫\�z@%P�&I4-,�=t�M�qX���P��:��v�!Y�5�*�I̱Y;�ڋ����dhx���u�_�{]��țP��V]�n��8���y�n��yh�$��3Z��u��׹g���;f<�@��KUm�XmLH���L�k_ݪ�ݴlfoj���iQ���.�Y�Sj7h^�i�O�jm�κqŔN5�-ޔN��;j�����WO�f��/U��ݰ0�꤮NE�\�wk1J��ƽʻw�;u��|:T��"��.�euS��Gc��g:��H��:b���'U�+�e��1Wp�!�|��ָۘ���L�B[�v
�E�0k8���ss�<�;�Y��wK�EHcXC]Djc$�/�����.�[賚�о��a��X8J8�����X���/�)����
l���Q��U�C����(啬��N8M"�T�+/p��:��:����ΪyW!ݶ�k��2-ڥAʊ����Gj�i#z� ��꫺8-*��h��G�_���nm*F�s]��.��2a��*�6Ռ�����'n^U�$T�wAʭ<��S��1�w�[�P&yO.s3����"c�n�ѕ|d�4(�Z(ZI%��R�=�xL�;[I��Щ;�%�5X(�VA�v��Z�C�>ҍT�b��ޡ��_=��s5�5�S��b�H;rԔr��U6��Fgۭ���2���mpx*�h٘:�/�t�����6<�����B�h�P���9Vb}mm̿�vc�\g)0B:N��]i=�Ǘ8�R�+�q/�ٮ�9�K����V��mr�*��G21T����b���;�J�봶�iH��&\���a���"�'���KH�J��P�H�:6�d�$R���3��JK�)�A.��8�ȓ�8Np�/0��^v^bY��2�P"$�%8p�E(G8Bm��Ift���q��h�)�r����qq�m�s;"�8�''_Aq�D�t9Ȝ�Y�n��V�u��Y�͚B�(��C������k8���蒒wͧ�B.��w�m���J''��pT��^��|�!"ڷ)"s���1���޷E��{nB"���/J3���mn����%��B�q� �>�ݷ|������1._
.�eQ3�I'Fk�J��M���LUͮ��Z�mL��~���1�S���gP�I�M I�qŕ'�3)����]����gq���
�=s�UhE� ���Z6��p�¦
�N�.�)wE�j��) 9m�#(���*V�����篿hdhhS�Lv�o�r��1.L]��.������x�I�	��nTLXŏ�a��j��R&�q�~��V�AHYךk�)�&�"k�P@��s4O�N�L�=:c-��Q��O6����;w�+�ƹ�k��$�W��)x�N�o���Mz��`�z�g3{/��mл�C���N2�p,reQC|t�����=�e9|s�a�E���d�T�9�J-��b�=���j���Sk�h·#�+n���
9���Œt#Ě���4uȊ����K�J�ċ�\��������/��I��V7G�O*)"k���$����qqgk8�͹cF��ۮ�XT5��""�w�44	�hB}�fK;��v�W��,E��qȪ8��=E�$�$�ė\�E��m��(�U��������+���*:k�6&qm
����q�hhg#�p�r�<Iܛ���:�eT���c٦����D�&m�v��IՆ��uP¨ j��2Y�}�;x��,{\�V��p�{R��k�I&��C�ω5~��å�G�M{/�S�^�����¹?tˠL��!�꽭ȫ,��]���:N̺����9�=�ӨgU��s�ʮ��yT)d�n�/�WAT�Wr<a���/F��dw�X��E_�;�N�������i���X�lu뙵�<H�3�C��q={'���a����;E��&6�n:�s����&M��wW^깞��[�ܒ�Ar��u��-e�
N,��6��m�����f*]��\º����`;;mL˥{lc�㬝�Ê:�עH����CDs�9Վx�ݵDq�<\rq��c81��!�.qW[��3u��u@Gn�2�K?O����X��6���E��1�SY���*ǔA]��L/].H; ������~z�����ț���Ӊ�{*��shv���<�Mdx�De.�}�/��&�#- �vY�gq�H��t�r=�\c}�]U��͜��ׁ$� ����fb����Wl�oe�\�6�@����[�;���$U�G@&/'W7N6�SE!��=L#��겧�;	]K+�Ȝ�&�I�J����W�9ʡ�{fK;��z7�.:�5��Mx����=�"��j`�@4t�XiA��)�b�KǞx{L������"b�M\կϺ�d�$��]�Y׏�w6��Ltm�q�a�G��ޯ$I�&�^��㪑e_��H������ys
�vŕ6o*/|�YJ�T��J���2��)��Cr�n�����jH�Gn�W]!s������� ��w����Nd���T�)������^JA'qzɳ����X9I��pm(�a�o���l�f�_m�	~�#��M{��$���spa���ξ�;�k)w�V�&�x�^�TD�A=�pA{e��fA�I�>$�'rr�m�s��EḪ̌%Sɪ}+Hus���p��.*.��d>����|�ke�S�e^�3�)���j�Kek�Q1�9WȒ�&�/ޠ=<�����=�=)��}�7�$u�Ol휶E��� I' $��5�=Р`Nm&;�ek�L���;�u|W'��sd�'��|d�oKu�̘:W�D$�N�^:LF�����Q2��_t�/���R�bwF�8=��ː'x�H�4Q�;!�F��_/ǳzk��q�W�E��<<=�6���S�X�����O�5�M L�l_v��Î[T1rX<Iq��:7�;ho(H���Ț�dp��\]P�V;����rI�	4L��9�x���ۮ�ɻ/��On�_Ɍ�^e����r&nVt��/M�æ�2�`g�x�/X��:�d�n��d�.i QN'������D$�w�{�6��!�Ǹ.��ޣFXN|�$�T� a˚F��,ٰz���Ѽ�m��P�k���䨓yWc�I�Z�<��>4<L�hH��q�Vԙ��i��;=�u|W'�e��&A&�5�Q��cy��ˢdM�������6�|����j�8U�Gk����}K��@�KxW.��=|.���f2K�{�^W�²�E�s� ���t�T�r�}(���p2��̧��qY�������k�:&|	4	4O��}�_mkȽz�Σz�7o;���V�5��I�8�j�=�n��U2h��L4�m���͸�q��AĶ�iU�nv3�l֦O߽~�����>>����c�Xg�r����)��=p�j�2���^MMx=鉞uo�N���y����o5�7w1ц�C/���jI/��
͂���y� �NxfiNqTՕ�o������G��#��k��&�"�g�HEP$ײ�S+S�7ۓ|V���u\�gm�*������=�I�IBH��D�uY��8q_9�� ���~�^jA&�%��1Ҧ��ۻ�z&ߣ�f��+`��J�p%�ە���gE��o+9��B��h���\T��]�C&6�rXaX�n||�y�����=���}��lՃ+�k@�r��]�v;M�Ӹ4� v.�a.ER��.ix��H݅P�n5v�۠-�2AVp�J����I�v�x72-1Z�n�4.�����b�\��	M�4���hEe�����f�!��3%�jY�ͦ��XtH	6�	v$�j�{v�8qZط����k�u�\�C��w��S�^�Z�K�hf���
�>��ߔ\M
QqL�G#6���ҖXlrk	��x����0��q[��{��F��k�w]�|����GҘ&�e㥖s����t<L�hknzme�E��}��������o�R���-O-׃j�$�#	�B�מ�4�$�LC�વ�>�}�����2_pk}��u$RI.�[�bG=�(��x�Nw^�|����G�:z(����å	"II#��^n
2�gUz*w��Cm�e�xj��+���[��>�Զ++2��v��&�Ef,�ت��S�"Ye�n��Eb�Ґ�]F�ۡ���M�D�A��⨓@"k5v7u�H:N����83f9�W+�Ms�h>$Ќa�W_Q�����n\>��i#�I<9v��R����B�gf�t���A�둽W�jn�KgR���K�	�e�b�cD|=����c�i��هY˦{(r!Lk�{��L��L��D�ԁ�x��$��̺�n+r��R�8o{�O,�Y��jyj��T	$�$չ�;�-|�8��Ϧ�_cwP�L��UV��� m�T1ٖ}��4	�k��J�b���z��-X�Q̧�(r!Lj�rT��)T׵^��&oC4]Q5H%LP`�L))R���7��v%Z��hY���-�St�I��*I5�Me�V9�l�u�qZ�VIʾjn-SSE 5o2Ow	�yt��
�=�u��$踬����5�;���c��t�<�,��a�d^bwC;�E��$����x�u���4+��͵��nU*�Xq��Ds��b����o_)Y��� �ݒ�XꉺyW˫+7�F�;p�ٶ��D]���� giOtۜ�c�!u�ᒾܤ�	(IRZ�@ߑ7C�.��M��ʷ<-��q<V�ZC�֎��a.�߳+�I0	(I�n=�ڼ��ճ:KX��7�Tc���`���I`I^���u�x<�aU*T�š�]�H�+%��S�v�6�ӝG`�
��l�3xrtL�M9�zw]��7r!,L��XwT�Ǚ��F�2	5�I��o<�f���g�$�e�U��l䛉�?�@6�ʒ'{,՝�#Ě$В!Y�w�4�����4Wg
�gj���u�_�E���9�7
YFAy�J�H��7�x��UȄ�=8�(ͻ&��e�;���>3GL�r�u��o^Q-<��Ŗ�n��ݭ�]M�Qf��4�7�)m�cUґ5»��1/����{���Ĝ��&I;�ҚȜ�ŝu�8���:1��q<V��M�&@G}T�c�CV��a�Ji�H���X���/X'q�sgb9(X�ˡrCSl%�V���gz�!$I�c/_cwQGX��W^��k��8:����Ě&A&��|�3RWH\�,��G^)y���&4��6���Im�DI9�L���k;)GOax����rH��<�^iP&G�4	59+dn���ˮ���7�� e^����bb5I]��x�P�u���Z����5��RW�E�)���Su�B���8���KV)y���&4�D��6<�j�8�9y�wT:�Fp+Bw��ݘ�jR�;]�8Mq��P��>6���[�6���v"-IK���=��gyoe����z��q��A�m�Y�d�{F�����U��A�嘷V�����8,<�%�6.�&�Z��/e,_+�;E�!�e�ѝ� ��3)m�ҸÝ��C�'���76����UU���5cI�j��n�,9�yM�6y���-IKK���Z2��P���S3�>2��^'�h�x���N�nv��-�Db�̶sQ�ovK��;KpV��qs|;��C�˔rl�{�eP�������3��g/��gN�U�������NN����W���ܛ733����7��,���N�'A����6�{�h�a����wvh��h꽛�-�l�X�f��L�ܽ6ڭ�}�2�P�ύ�cibvk��v�g-�T.g]L�W��>�,N�\�y
�W>&�Ms���o8�����]]��k�I6�97���OW`ǘ��77Z�̼w};�(�KC��<NQ̴R֓Яs�Y1�N׀��.�W!E�:���c�����n�F���N!�hNx E[��ZR�w�V���j�5l�s��*�w[�B]*�<���,���ecR�D5;i��yD����X�g��˂&/um�*��h{��g`A����^6�h5yׂ���>��g�v������8���}t�4��]h���YS�.�3�ږ��y�v[8�24#��.Ru�N�k���n��f�:�I1��*���-��C*�̮�h�`��ugs�H�E%8��(��@}n��$I�jzl��,�����]��!�{v��E�ko=N"γ�K���H�^�������y��G�[��m���˽�m�+-.�<�<�"��q^�;-#�;:�^a��$%%�'m��w��yǴڒK-r����r�,��gEy�ڊH���M�혀��yG=�{i�4y�y�u��zvqy��Vp�y�E��H��쓬��=��S�ܺ<�g�:�N���R�w�[nNYY��f��o^�Yy�����6�h:��#���{��>Lw]��x����Bo�e6^�,w\Q�3�).DK�l�exӜg^|=u=`�U,A.����Z56�m������x�k���LoӦ��3&��uB]1�	E�ƚn�8��jDM��"[l�Yvf�4�
�˨�m�B��Ĩ�=���Yq�aՄz)�d�ٱ��z�V�N���y�b�WI��k<��r]���Ћ�;��RJ��ت��0�2����lRM6�,��X��l ԓC$�r
@��kZ�4,�m.�nD�:����=��_-k���e�����綣M;�J�ۭ����|�������۱�2Mln�{�X��|4�.3��N-³s�k��,��w��֎�,><�c0܌=`{X�Jvͺ1t���0�gO���ё��rc�=�i8�n�ڢ��X�m<�njJ��J��̔��U2�ݖ�M]nPu[�b�+�l�ʲl�K���D5y�v����[�Tu=��sme�ӑ�]�'��C�c7M���L����Gj�:�%!�	���6�Q6B����y�y�g�6���lK�2�K�lA50�X-v����몈������!��]�=��Y�܏mͳ�5�K�<�1�7)������ZVe��$���J�۰nz����8}v��HҎ3��1�87$d��-��.Ԏ�ܓe���pE3�*
�Y�\ٵ��q���uڴ��)�;PqF��!su�I���Z4G	swj�KT[k�nٳ��\�F@܃�qO��=�}���7Gm�\Żc)n��k)�K4��Q��ґ�g-�m�i6D�R�Ο=e����)u�E��!�:�ˬ``�iqv��8ن.��:�n��6 �/]P��M��Eٸ�pRk��Z��)��c[/Dx�[D�B ��CB.�܇9%�{����`d�)a��iKZ�1�A�-�ub0h��]�vJ��p�r8��<k�/���C�q�;-�H9#�U�n)�h��^.�[U/���w��o��и���7F�b.����	41c��\P++
�]d"m��;SS��N��=��Jv�J�;������Y���$�Hb�%�K�ɚP���I�ݐ���E/�t��Z@1yX����t��Q��l��h�	t�,���,�P%��vko8�B�vTi�r��n�y�<t5�M��fڶ�Й� ,F�E�5�3M����Kt0�X�=������H�kZ;;�c�b�D���b8z{q�Wcrb8
����w/J�H�D�v�����Qs�j�Գdm��F��벒TT�Mh*�����<_W��&�]��]O���{��P�T�@�aq@rZ�L��ܬ���	(IY�t9�Z��v�R�^+�BX���Y'|L�hYr�\sI�^f����/<I��Z]���p�\�Z�����͋Jzb�4���J�JH��z��O�:����̋�����2�;���h��Lנ@�Mi��q�(z���K�B��BV:\��%+���a�Lg��M1kٔ4�h�1����>~��{�F�����@�Ƞ�7e�x�Ef+(�aa��gt?Gf�fx��i䠁�����l�~�&ۻ�;s�!dl��7���m�
�!r����:��9�,w}fb8GLΣ�.iiwh\ޅM��	���I�X��93^�Y��?Ā�t�g�%5�}4�������\��˭S��C�>��#��0d���,R�E ��4,���t�`�JDd��F�&�J����_*t�zr$���-��~�2j��r�)L�0D���^��n n� ���핀�%��3�<��\Q
����h@�.Ɉ��o�����^�%�q)�;��WrH˸�{cݟH��p���[}Γ�x��4U2�<{����Jo,X34��5�zŬ��r���a,P u\�Qى6�FʙtU4����ґ�"H�r!Co��T�ؔƪ0���R��=3j7^���d�\lh�;��eܒ6]�#'\��"c�M�[��s�W�)�3a�z��̴�
��Dq����Og6��<=��ו�A���ɐD�"$�AH�x�j�ۊ�=j�R��e28��ReU�ۣ�b�9Y鷇��ݶ�1x�7����l;�V5�xݵ9���⹮��1�;�7ul�Կ��6vlS��K���!����{���FJ�#c}��\�M����o����"c���p�xb�p�1�XΞY�2�*�� �퉂$����#�%#!��y׃��R-U�ե
��I�-�,@�3B���@&�;>-�9���^��pؐ(��6ԛ%�qML*tnLM��11iu2^�-�U0�l8/��?�_N��I@I^c���`��1S�r(W[��
�v���s���A|� ̔� ��Ex�x.� G���;�9����̷������z�T3���Y�GG�T�g2Q#y*����F2	��T�_L�ٓ�7��5�i"����H��$�����3{�5�1��A�/��HL�1y�p���פ�R��2x At#;���(�'��g�a�p��N��]34�|�{l�jY�I�UT66rܣ��Q�x��c+]q�f�p=u:c9[v�2����}1��	e��+�R;�%2��h�`O�z�%Уe��ٗnT�[��xL��{�@�)2Dxvu�	{7�>~S�����h�C6�t�*
��h��Ѣ���X$m:������vSb������'��Q�	� G�3a�z��̴�
�tz]c���s�#{�H���T�w!r��d���8Z���H�NLe�L>L��9EX��DR+�!�b�ϲ���H�{�%3��P��K���]��@&�(�N�̄��Bٕp�[�ex��S ��_%|��2$H^�G8�r�,�'�цvRd����v糽E]��/|�e"=�.]�#�[��<��}_%"2E� �VmcU�	ajƞأ�u��k�V-�9��$l��F3s(�wq,`���3����OԄY��a�cQ�AU�sn�o,�Ɇ�v*�-w�w2�6�<�1hE�5ǜ,]佻5;��+U�T�;��2̺r�[� |W�P�GQTE3�`�2�݌�D�r��᳚nj�9x�\j��,hԺ���c�������ËP.�@NZ��hL��ѳRV+�jRd�2ۇHD6���v#�'��
�Q�BB&�i��XL��.,��QɌ,fn�٣E��u�=[x��S���t�ʾ�ru��=�ڻe�F{y�f-Χg�T�.��.�W&��RkƎ����w��N��-�p�;�ohe�6;pq���6Ӓ�4)���R�һ���?����uD���[����y��f��E���v7Zr���Bs�I��"3�+�J]���b&<�q�^�1Y�����~�5�!$�~呜�ӹ������ҁ��H�0$U���ҏ�1m�����ڵ�b��a���"���	Ϩ7�����u�E׈� �#}���9ؗpҐ�v1'��6��H������Ԫ� ��x�@BH�2Uܫ��_! ���nƵ���Wą��?G��@������np�xgW�@�A�@��s��f��0�G2b:�WV��8X���q�ڨ`𞥗��^��
L��x�W���v�c�=]�r���u|�~1��1��K.�+eݶ	��ٹ�w��3�[ٖ*�i��*�x�r�Y3�Q�K�+{Nz<��,|s��o^�B�U�7%��l����΍���r���(��V읭���9�R�<OU��5B�#3���B�vf��k���tH}��|A�IfJ@�����[�BL0��*f��P79���O��	6);�$��>��f��6�gF5��� `�Mm�6��K��vaV4�"�����k&�c����l��F �H�+��5L#a�J+~B��p��n%�5
�@�'������2E��v���:Xϼ����UE1U�=u�^��f`�[�x�>ذ�X�R��MX�/7|���Ϩ@hб�z3�Y�㎽nn��n��e���Z�Z���e|���$��2 ���@�"s�����"�@�f�ۛm��S�=]xU�,P�d)=���w�f�ý�<7Ўn�'�}%}`�#"TJ�n�0��yQ<��6bb�u'o�9�)|�Ź�ݥ�x1py�%��]ʤ��°�t���Q<A�T��s�1��U�;���;�{	UĻ�����#�@�<j�5"�� �"`"r�*��#Tj��;�zR Ⱦ|ߎ�f{����������x�a��x��F����("2E��)��O��q���O �]�X4�BZ�W�@e_���Y��y=U0�~��e�#t�"^���c���1�gb���cla5^횸�����D������A��H����ff�;��z��t�pD���W��4�O�N��<�%��#��Wptwp.�=�o �]vK!��t�����ڍ�2�^C��X�eH�wg=��eUAR���A|~��2�d��&H��ޱ�[��UR��s�R�=]xU�3�3�)��2R"�$l+��t���p@�^���Я
��Y���^�!va��A;�20���.ܷ��9�������f⬠��k�φM�f���;��L���H��7�43�g�}j��$�2��3�y��T\�#�9�>õ���µ�쏽EU�ω�$߉�쭟�ւe�Uz�ZϠ�����[�e@�.��rwvR����Mo"돳�L��n|ܯ6���ml�'�U7�W:0;qurXb��0�l{!�<w��@.�A2(@�$Ձ��O�&���ׅX��3QZ�i�s�|Ջz�R/��?) DVu�Fe�>�7v�~&�z�7�t:��z�H]�d8�� 5^&Bi�3SGi��A�	����J�d�0��E��9H6��t
���T��[�e@��X��>�5^��>&@z��d�0�}B�Ȩ�c����Y��MZ�s=����Dؔ"�%�����ݞa��� ��&J@�a$���5+��� �W�>���q�!vdbG���TiL�C�۷2�T��X���U�"X��oP�Ԍ�w3˳�n��3�^����zU�
�4oʜ5�Ju^�]X�����o�D�.T4Z1T����UF��p��mN��ѱQ�h�Ņ����b���x甙��v��^�1�Z�45�����5˭n�ݎɞ��؈o13�˩8k�n&�m��ւ�;�]��@pr�X�6��ks�+i��jO7�$Iɫ��'����l�3�'fȵ�>��F�UgXy��������Q���6: Rb釬F���&;MY���}��6����]ec�n
��<�G�qÛ�٘H�uږ�k�O{��Y���� ��&E]�q��yv�P��7�e�"���L����� �"JDd��/�:;��uW��@*k�zucsR�_\M[��걥��P��b���993
���7��� G_�`�+��F�2 |{7G!E*����w��V�R`�,@�F������"$H�B�^�o"�B�ڨX��D"ꛞO5�͎ǲ��7�0N����_U�MP�����)L�2� D�v�ھW���vt��I�MZ�s<�#��#�`�H	�����O�{2��6hi�ݰ�ח�oQh�7m���)u�X�K���	M	�I�۽����FuD������wk���z�H[��\���������ޠ$�"@IA|�����Ǆ[���W>n�Wf*6�g.Һ&O�Vk4UQ��]\simV�+4���X(��1?{ޥ�>�SB<������y�-y�Ų��7�0N��=A|�^�O����ߧr�.� A99?�"D"JD��Vh�k���\��۪O�ծg1��]��fJ@��FǸc�i�{�s�}�HƟ6	��WpuOsR��/.�R��1��t���_����D��,����d����nz�D!��t�����4��-��9��_��D����wx���\fy��m��X6�n&�٭�x'gi�O=8�s����ėD��A*�Ch �rrdt����z	5y��s�2n�3�gU�N�Fpmq(����^s�R%�6�J@�T����7�6�����Թ��̇�T��;%����p 5B�1�Q�;BS0���^��@7"�G�6,�_/���5F�V)��ơ�v�ݛ�u�ν�[n�hԥ�J��+s/�����!F;���>�]��h�.^��/UX�w�d̒�os�2.OO�8qK0�55j
#�F)9����;s�!Vܚ6�������ͳo`�1�G�se�,��A��t���#ݨ9O`�#X��YB������0��2�7|v�q��7������M�ë99���.��X�{+:�q�OK��֋�7%h��Ȭ��#gY��Ʋ��祫�:�j�6���e$��ss�͒f�7[:����J�ɸHY`���ʂ�n*�LĬ���ӲQ���B�V��t��u%�JLU�8/��t���Uh����.�%B.��m��.�u���Z�b����Q-��SZ24��>������L�;��G��:v�L9�e���m�7`�!�̯��e�{Mj��N�7��`��Q�Ie�-�tե��F�җ�7Q.R����%�м)Nk���f���ݬ�u{�k�s����m�{㑛X�ln��/�:�9U/p�[V���(^����cx�N5��T��V
,s�
���r��#�Y����+���̬ۧu���5�%�K0�D���}���N:���n��'t�;�1��31v�ܙ���҆�9�TQ<o�-�c��!�3qZ����F��s��%eJ�y�y6�խ]�b1X��!�ۢ�D{;����i�[\������[B�v�2''������t8]:���ᆲ*���e�U��]>ݛ�g`�2�c��V*��2�S�}����Сh��å��.���wWoCf����UQUB�j��)h$�oM�8�c��y�o{/9ۖڶٔV��{cmm�gw�۹�m؏=�<�^ۦ�Em�mYƚ�m���Y��pin5�&-ɵ��&Sy�zw��e�zz2ԕ�۶�p�@׷yOI�n�n�į{yw����u�l�^��^��<:����׽��6f�Nt�[/;;̻�;��$x"áZ�m��K@�X0��-/"��J"�Z�;6{�sݭ�5��ܬ�sڌH�ޘ�±Ff��/;#k[Z��i'��Rێi����f��8�m�X  �)[
^u����;;ӣ�m��Zd��L��ֳޯw����1۶�!���8�����9���TN�v}q����`��� �P@�#�~�F�Do%����߻��A�A:�"fk��Xɻ`�m�V1H~-H�V^���_�9��̉cCۂS.�i�ı�%�E�S���s!��g�Q
�N��d�CԪTv��F�mP� 5=E�غ�Ԡ��1J�)�T
e4J�);gN7��Uv2��)���K6���_���Y��A���`) A2PA���fz�^�eqg�˼�(9~�k�Մ�A���D�/����H�J�B������g�#yV��Z���Y{l걉� Z���ta�%I��U�b����P@���펦7w���T�ܕ�\\�Wx�J�������ܨv�{^ ��L� ��� �"`��UY�y�(` �oX�*hG��t�>Ou��K6�J�gh{㲑�k��u�=�{s�IyN�nUM��������;�b�ԣ5\�fH��u��d���Gd�+V�w.;���Q��fi�JU��ٔ?}QP������aR �"`�("$�%��w��l��"^ѷH��6md��*!�A�F���JB2t�nq�ɿ3<�_���e���qk4���U��
{c�=�\�=&i��ni�&*e�=�
{p�w*�4'qq���2�R`Ζzv�r�J���&�=���y��wsI�r�.�"#��1*ά�RzPM��{���7E��R�Y���j<ԀI3%]ڞ��GpIG]/�'g/��"$�AH�A�X�����_+����}d��3���@��A�F�JJD��u�d�g��I�oH�����+q����2=���;b��Az&C���v�Q�O�F�F]/��"�JJ�$�?����z�UU񍬥��do�����7E��S����߮%�=�%2���ܞ�l����S{!�h�#t�8��XZ~���nK5ΪV�S��\�cZ��A
b�IN��沷0�x����^���sg�+���θ��}k(U�"�5�A]/���Y�]$/;��]��݌�nԐ�c0��Ny";\q��j;a�U]��;���RR;R ࡦob�����v)�����鸻co5���gl��=�5��;c��X.�F�]]6�*6�]
v�ذny��k\V�=��	K�9�e�1�bk����\@���;qg�8�;i�j�ܽj6�x�"�Rz��i���Fj�>�������q�,V�=��YO'����l��Z`�\S2�SFM�|�_�=��r%/�&H���ݷ�O�L�s9��!~�$�ؖb���@hͺY������(wp�������;H��9+qq���2�R��gK#���}�"$�����x�pW��`����� �`�HeC�z��vq�曃�%�M8��W�y�w�}\BIFQ�o]����uj�>�w�~�_x�`�d��㝷�O�L�&r��a���K=��<E�$����	P�$��;�ϸ��8�B�S\�E�C�*T����r5p#���0�fH��1w87A	��S�4ؑ�q0-n�`cv�.�(�&�2��(�kN�Έׁl�~�s�H%|���{��ڊ߯*uqqtj�]�oCU�AGy(�쫸-��#ww42]z3G��L>�i=6�2w\r3�<+��G|̂n�����}Y��̱d�Wd�0����8�^�^���f�g_o�!����� Ƈ�������|�5�w=�T11B"����ѡ`A3,c.�N�"��R��(~ؑ���,���˹ d�Q|��z1�*f�9��
�(d��%�7�Om|�"��ӫO�ֳ����y�T���Ds��z�)�7�F����U'�]����j�U���u��4 ���g*���z�j�E��o�'3T�d"Mˢ���;�S&g�*�{=P��ɧD�)"Z�F���b����P�kv�� ��]m1E���O�y�M-���@J|	5� �)��Fx_z�J���<~3�m�ʹ{j����A��?I�b�C���a��T�k+��H����{�K͒�@��,@�s�j�z'K�z�%��-g��
���@�f�� �2R �$N?Oe����J������$��l�Kg�Ԑ��0Ů������n�r�ǍѼݤQ{�`u�g���ouW^�ux�=֐��^��ؗ_wl�G&��C��RF����"J�#a�v���i��{k�� �~�Е��T��I�7e����C���kٶ��=�D��ȑ2PIfJ�X���Co���j�E=�5��d�P/���|ˡP	7��Ȇ1CwVG;S̻�F��??��*�
ק��G�F�ɡ��r�絎x�ñs ��k� ��_>� d���$L]���O��ʛ�B���jiF���(������"$�0@2P�骱�b�ۃ�b��B�,�y��o\�P�v\;�2� ��类��z�}�'z�IfJD"zb�i��;X���mT��*uqs�0N����<�"H��A4(A3�xFIt8S�2r���y���$ՌͲ���V��=�F)��Po�.���d;a�5�|�j���Ÿr�Z���v�P<�eV�;�V�v������7�/�q�hz��gc��"�A�a��O\/+;��zO�* ���J@�"�%!Q����p�A}ǭ֊�oY�
�e�G#W� �� �d�M��
�O��Wo��4��[D��Xn��c���m��l6��-���ή�g>m��<�@�2+�>W�g`G��Ae�֛�,��N�!�y��������ꀋ�d��D2R$O�������j�da��.Uc3l�vqճsOj���A레#�+@��צ��62�P&���o�1���{ԩ5�I���_w�E��>(�>��ΰT�ݗ#������H��H��f̪��q�t,���S�Р^�>�1��^����p^�WWb���׬��3�� � ȂJV����/'�b��v�Q�s%����{�I�s�>�@�z� A�7�g@�L�94c�q�X��&�7��^��u3u�fҳ���Վ;�\�f��n�b�q���ɓU��$^k��w0�RN����R�8t�L�E4�M5MjKJC[�02�w>�N�Bg����{^1��K��7	��g��:x�Jnkj�mu��^s�N��v5ӵآ��mơ��Ih�n탫�Ok��Dm<�l���{fp���E���s�l�\�p>���F��E���ctт����0p$�';���.��ʸ�Y��T s�LLsj�.#4�����.�2��9�`��O<�:�+�ݶ�0���3��hḂm"B��0A�K�r�#��dA��V��o\�R�vX�O&E��y�ڰA�A|gR�?��/���[�j"y�*�|+_�٨΅<��}��>y[9|��9�@��$k����&0h�"X�{�Cܒ��H�;����������#v+��{�N��E�����K��D���sj�{�PV�DΠ	[~�hR��V�p��`�Y�.G>��H�Dc�{�����M��*�	c�����N�ګa_��Ln�{u�O�_=�<sԈ?o�@�"�J�FV�~}���*�J��}I�p��]np�(�(�D��R�:-��읺���k��ܮ�f�3�#%#��^\}�-�U��ؤZ�go(��:C���~*w�D0% Ӹ����F�P��"�J�� ��3,����C��I˝(뉓�k��^c#j�(��Û�W�T�7&3s$�����u�FIטÀ��_*�=j�c��s��`@��u����Ũ�q�Ī�wP�%"�<I�IXD�������n����n!�1~�5���I�~&EA25|����9�� gP�ϫ�I��ӌ�X�r����"ӡ�E�[���_D��"M�	&���D��u��9��My�.�;K��ڎ��K7e���y��3�#�I��D��8ܫ2���}�3�¸�e��ڱ��mэK'\�/��4���-ӣE�D[�?������I"�^e>�l^�P/9سWp�E����/�/�Ό?��#%"	�&C�� �|b9�kpW�Ё���7N#(c���wŵ��	c[���9M��	��d�ս�P��ҥ{���]��P���FC�{*d��^�W-�Ǉ��X��tw���7���Faw���n��72������K����._n�|��
�����t>Σu�W�'sɂ���2D�"J�O_���O,z�H>�wX�nh@�M
���S�kͱ:����/��I��ǫ�4����?H�����&D2Uuju�=]�!�H�����:�g_���"�����_G��3%"$�[roXa�a~>߱a�� :s�qm��
{;Rb�`���Kh1�3&�*�΁4��vR"uD��� ����[q�ީ�	f��!G�D8��7$�����ʻ���� �V��F��8�%�#zj�,��}�	lnv�fs� F���P�I�N�O�cv���.�%�=��w���Ɲ�]���t�����/�u�OR-?
�}�a�%"�	&0h����2�Cf��{Dd��%��o���v��!,Ζ G����@n_D쭢�6vީ�T9�[OOI>�2�=�����縚�X&�������ne&������S��ؾ���ݪ��eMf�4z�6�������"D�J����d�̗t�"Fd�[�5���!ݸ
�w�#\�耒c�ȇ�e��vr^f��H!f4(ǗY�A�e�i�e���$z��{0�U��)��d�?"y�,l~�i��6_P}C*��_�����(@A����` �@�#�����
���Ϧ�0��ATo2���r^�2��ь~���*�";�9�g�>�R�2X#�	ޠ�H�2R"J��0i����Ϻabہ)|��k�Pf�$��<	�@A3�{$���}���U�3������f�����q�B�R-HqnE GUe��,3��-}:�Π7u}�PdA|D�O�Vv��uQ[�}�AG3��cڷZ��K3���Gk�!��&@$��*���U��+�k�1��c%���
�ƉGK�E����jVhɊȻk~Ûut�ܺ�Q�3M2.J�ڨku�B	������i���T&p,Q�d�;EۄA�:<v��m��b��[�.��koYݬ�6���9�V*>���9Bn�o&Χ��X�-�2��%�og{����U�t���:����Ԯ���֨���/�m4Խ���
|8&K]�ɂ1�wOg@�r���;m���sL{w(3]�[.���,L�o:���7s�:U�g�*[�y\��nw�Ŏ����Wr��V/�=�'��Ҫ�WUz��Fn�Z�[������e�j�wOs�1nU҈����3�e��`ۺw�{���=<)-�5�{��0�Ʋ���V�!�6��3q�\$�J�2���V�y��⭣��A��ѻH��ԭj�u�m��K����ڝY',K���N��b��m�nl�C��:kWϋg2�4��B��Q�*��/���mq�v�ud���A�z��d6k�	�OO1V�E��73�U��)�c�m�s�i�\ �󽪵|Q>���'v�}R�Vv����3�6��pm���L�1�إ��eJ_�WvN�á
�rul,WIX�dӝwӯsyZ�.��[�/w��ե�Vo����m��x����/�v�ko�\���O�}��!7�M���$ͥϐ=�#�a�Ḳ�}�P���l��3�v�,��ab�\#�5s�ssp���|�#n�^�y�-�ҽ�'!{l���0v��0���w������f9��e-�N	�ghF�,�ם�f��P�H��C�(ib�K 
L�v��͆�,\&�ё4ɵ�^�{�ݸ������ԅ��3M���hkm�l�/4/N�-�mi�4m1X�qk������u���5��{ր{-�n�.M�8rDY��[������h�'��6ؖ����la���mٳ���hmӶF�i6�,�f��f��
�ؖ�K:��斞]�y'GK!�Ds��fY�c��-���+���ۥ�y��ZY��Օ��km�i��i��V�k5�ֱmۍɖ�ڷ/M�im�ɴј5�Y9=�6Z��v��Ym�nwfN6��,ö�Vlkn٠V�&vJm�Z�i�����!9�9�5��m�m�m��v�lk9�s�b�!�qN�Vl�,������ڞͽn;A�Khu����
d�=ʅ�&��k3�{G]X3��h��3���\v]�rq#�`dC87`n�᩵�&����K�M,I�`�b1��sɮUܛ��)s��c=��[�Za漺ō�����C�Ү�c\c\8-ܹ��P� �l������B@מ#V8��y��"U�U���v��E���PM�X�y�^����a"v�l�6;G���v�ݸ��p��ŀ���5�&n�yt�GO�'r�>6L�b-��+WP�, ����<5܅��CZ��.�b�ru�7J3��aϐ���n[.�ã6q��Bm[p�v��}�^zm�u1��ݨmI<l�G:���t1HF�N�9���Fז�k&n;gd]��=�����<��t�s�Қ#'Aײc����n�
�uFè� ��a;q�ga��D���¬��䫫	tM4	�T�V�\k2���Z._���xÞ�%-���\��)A(�MJ�C/['D����̥�Yc	�����jTJJ8��0%T����j	+����޼��Ջ���n��4���e�ޣ8� ��4)��knz�73�����.u�UĻnS�nۉļ]l��F�n:��u�&�f� ��X9��S�q�ѣ�U����O<���u���4�L����Mh�p*\]�T�Їda�s3�����Т;�$��-v��W}��F���}�'���d��Ů���	ua�����B!m�+�H�Y�m-�F!�=�xyzۤ���m�ҷn4�f5�F��&c;��B�8��Bg��|���[�yk�o!X���
��p��i1S�$��6Ki}75�3e9Ku+4ȑ�Sy�)��OU��;pP[�U�[���3���������A��f#us�����t��y(��!ָ�B��մGMh��I�ۈ�t����n�b�!�p]����c	*�*v���=�R���;Xઍ�h����=qYp��7qͬθ�f��.\�`ͯ���VR;s�E�;uv�*0�8�\&nT2���0�c�n��d��r���M�B�D�Fˀ
�����	(�]JJ&��WA��Kr�f:��	�1����bMm��а���I`�+�lmG6�X�PU<a�i�۫��^���m�d�kQ�
�vM�+���(�⣍��SD��5���.�O���g��2�X���\�{]�N��y���ݫ^��Ť�r���6F}#�+2�;���]�)fn�[�x�v�JE�;�&rm�7ْ=u���Ⱦτ�#% AH���X^k��խD����5Ҫ�O`�Ny�x��/�>������d�n�߸�K�>=A�C�a�vR ȂI��hM;�����N�N:�FBY�,@��L}� d��"D��{�y���!@�ٶ,CS^�Х��z�����T��~� F9�p{Fl�hKw���w�T����SWw4�2�IN�:r6v�{�i��:�i�Үn3hQ�}A��@��A=�A�)@���T��C����|�=���]��n#�1�s��@��%C9��b��YBWK��-��o{�|�P�@$׉���y�;�8�]	ft���*������k�S����I��� oV��
$i�r�]N�oP.�+]d�P�讵~��ǼC���yE���F�*�,#Q��ݹ��q��T�f��|�cK-ɬX�e�j��f���>�7B����c�f�۠�{�	�R��JH�;T{u��w ���7�@�K�AH�,\���U[��<�fУ��OE���b�2W�H���#aҞ�s>�f]YZ�P4��&�y^�4g{g�a-Ζ׻��,wd��_m�wI~ؐcC�ɦH��A�����{<]y���:�1����q��n��]� F9�@>�	&?�� ^�Wa���j
�A^َ[U��qGiO%OWm�J��_n���&��{�PL�L=A)	�&/&��Jy�͡G�)��2�:�sÝr��0�3�� $��2R#�i��9��G��J�y�;״�m	n)q�֘ ��@*�;�zY�hxƟ�f���$IX2 DYXU�쫼�[]1̽�"T����U*�d���ڣ(T���w.}��E�kރjk�Z߽{�c�SRu�bٕ~]�M�$��v��ٞGeCVO!ۦ�����A$a�~���y0���6��^
���ԏ�D�d��=㘂�3�>���{5J����9��	�"$�0L��	@�%��6X}ݨ/>�c/RH��N��F�[�\��V?{�@�HL�YV�����
�E��紝�8�mmz.q(A��.�%�i��&�-[���M6z�%r���=�J�:Ʈ���r^������
�b��s=u�=��U��P@��}%}%@A��#�t�Y��fk��X�=��9|�v�:���F�la��Wq������Wmߛ�3׆2Jfm�C{p�rJe��&��NO����)�<gk���a-�.;�� ��A|d�?"`�(^��x{k�ԍy�b�%>�	�^y��K�6�R�a@�,X��>�����9}1�K����"���gET�}x/z�&��S������lT�v�{��t�������Q��{�d�ΥC�;��� d�A�� ��R�Z<�� �R]�4җ�whQ�E�B<"܊���a�)dB����V��ͷ��h�QO�Ӕ ��Fw��liy��a	f�X1�t�]�(=�M7��'}H��A$a�%�^��#=],��6�R�����`I9[�؞ń�A�D$L�_IA/�t|�V�u�����A��9/X�\�ܸx�� ߩ~�"Hz�Ȟ��n�����2��{��P�% AC[y�������ɢF�Rz�<uH��n@��ظ&}^�4'lH�M�8��z
� �@wLIA/^l�:����Á-�/�#�ڪ��ˉ���YX��yr}�Y��v&PFJIfJyW��$��BrFz�s\��V�U�T�����hNߣ���3�0�z7jX̔��X�vh^�{b��R�ӹ�*LȆ'#Nv�ꭺ���EX���ן#��.�p�bꮥ/f�'���[��k��7f�Pp9����ۧ��a�<1�,��c7���<����,��Z���v S���)N�(:��V�pvW��g+��)+�GMm��g�<]�a��嶧�t��}�]�E���t���m��Ի�%��&b�N^=us�oe�`�p:����8)�`�קV464!��2�1�v��%5�j��S��ce$.�$�BVi���>џl�[a�T�*jʌ��&Y�6͚)��pI�1F�߽��8��������?M���2X��^���
i�"���T<ו�e��8v�T&��$cEܒ�wt�wq ������٫��q�CԷx�])����RǠG���#�W����U��s]Ρ�F�f���R7�YwrP;�Wp_����Wg�s�P�Ԫ;l�������� D��� H�����uV_�E}���0 5"������c)c��<w ��u�K^�S3�1/s�21���F$�0L��"J�'�?O�n{���ʡB�������'0%|�Ǌ�@�5^��~2Edm1�n��7I���Y��Wk�A�b�v:l�9�m��\�]XZe���a�G�P+B�@�%#��`�H�$A��r��Zy�v�S�9^1����������zɡ^�f��j�(��)f9� ;c�����9_CH�ࠄ�sSD��onRF�f�V���SUS9s���G�^z���}FMض6
���^DM[J]Ձ}XǎJ@��&2�XÎX�"�R-1B[�P ͋�d��Ҩ�!{�8$��j���DHl�x��� ������zu�ԍ>�W����|{�0G��J�"dH�ł����J�m���"�/��+N��ӊ=g F9�[V�SB�����os�'�$���cC����]ω����-�,�_f�qK�dY�d�	L{��K��s6j�2=�ߣ�\[i��7ka6�� �B��o9��2��9�fR�[���C�O�?+�'�DHn�L�Y�u�l�1�8%���uvs�ܫܰ�"�H��?���J�kLj�RP�0Q;�̘�{�1�~
fu-�|~n!�oԈ�@IK���B�$��1�����]� ��X?$S�3՟�^����J�6﷬�gvf��T��M۩X6�ΑKK�}�nj���"��7ږḖV$u2/:�C))�e����{2��3�>��w�J�:��ܒ�wt���ka�̅�� jU��4*�wa2�r�	f�p	��� �
�<���v1U�wԏ��&D�d��"H�Jc����u�B���V]t��s��K����?�"D�I��"��}=V���.��=��~���Fyz��Q�N���X垦g�vu�q�ȍ0�6{+�~>�Lg�@�_#$OsN8�G=��<uH��@�R��$/�.*5^��t�0gRIA$ld���+יUDa��%S^��hP������S�����'� �(P;��V-����y�Y�z�CR*l0d�A!\�W�o�S�;^�^�^Mn���ף�����S��oԁ��"H���"%}p��(3�����V> ��9���ni���籷'���Ԥ?G���/=��u�u[Vwz�g����
ʡ}z��u�'>NRbm�w3]��܆��&��2��8\�2{��2�e�T'���M�eN����܂"H�`�d��PJ۶wh>u���.�E�U�ʞ��,� �br�H�$^Y��V��A�hf����֒;^6���Ź���j�V�K۵��Z-�Xv���oh A���J����ˬ����G����������g@�n���ܒFf�*N�I�Jj��Iq�]w��Ԉ �O�,d�E[�*�l�"��r*$lX�eW�a�ߣ�
����{�|A�DF�H��~���f�yͩs�J��-�>~�z�`5B���$_I@ןv_&�P_Gv��ޤ�h9�u��1d#��(�b�F9�w2�t,�/���=������ �d��A�}%Z��ܟmj�@9���lv����
76gP}���D�JD"�Չ�ھ�}R��M��ߎZ����l�뽫j�%��K�ݎH�u-����$�kOE������� �o�����7�`u:��{4�^~�e�w���y��}g��m�Y�\�LFa��]�]wiF0�u��҃!]6:G����e�6��M�;SZ`¢(D���Ų���rٚk�X��,`U�fb�ff�4
�ev5�۟ �m\��8�	Vvɠ�t"ӎ���5�m�<l3U��tG8v�y�*.������7-���F�\J�K[4�5�������`��u���z詊RVi��ߟX:-.԰��볓C#.ή֝E%��%��X)�4AA�ψ_������??̜%B�k�M]��I�Z��\�R�mz���<բ�w��LA|d�"dI^�L�:p��b�`��RT)��Ny��g	�Q�6ň�|̌�N��6�/����@�����2 ��� �%Y6�.����($Y��6�oR50���PN�3%"� ��!+k
r{7h��\5u��/��?��.{�-D��	g)~�3�b*����{���|����PFJ��0�2U���0,�2y�8m,t��c��'��z�4��)�ܒYwuJ���w|S�U�����-�	m4�,(���Bf��a���ST3R˵لmq���=z�/��],���=I��I��Nɛ�cd���#S�x�/�~�����ʇwq��H�� D���J��;wV=���AXw������]'�`jУ��u(-���[�ko
TEN������.���#���ڪ�f�+g��np�ߠ����J�VHKyK�y�5#`��g6��#{^��+�=�%szH�݂F4]���/�"E��C�ؼ�o[j{uA�9$��~kP�R ��A$��(`2R#��5H��/��A��zW�$K219�}hl�:�b~�[�P$�
Y�s�i��!�9Ԉ?lA$a�d�A!B&���Uj]Cٹ��Wm6L�ZS�p�����z���W���$�Q�b����&�g��q�M)چ8�1���櫎�o/mL��K�r����Yz��G�#�0̔����_���#�9$��~k|~��Z�Um̭{�#7��"�% ~�/�^VU����䮕��` �b5w�pپ�7(�R1:�T���2R��_���B��ر\���7�!�O9cw�ʣ�{IP�t�0�d��^��l������LV5{v�Ӭ�0UK�w�asظ���̧�q�ݻ��e6:�V��;�e[�\�������|r�_a�>��{{z���7�����c�LVRȳD�О瀨�p��;���t��{��W���ÁY\̦P���Nя�r�=GwE�ù�`��Q��uU�kj�楸�>��jh�*�j�M&Ԥ �]��gXy���++_9I�{B���yW*�muE�]��{�g�55U��ޞ:법�՗j��R��Pfs��y��⤁�w��8�w:]ǧ6f�RZ�fs2�H�!O*�I̷u�;�]�;��2��sh���8ffS�gS��g�j�,��FK�ܑ���H���q/B��[Ɓ:J��˺	
�5��ܭ年���ef^n���U�F�ǫ
�@�ޚ/F1�»V��p+Ut�޾S�^����ͽ[�{�r��C�[���V��B��wS�L��;z�u������x]�t��[W��v��b6-B�R��k#������]`������6�c�Z7v<6�4�i���Y2���ȷso���:�Ax��;�E�&Wr�U|�zM��#�$ʱ�֯p!�������R���//�iv�]#r�a��z�F�Z��r��1���P���l��Ur�Hʗ�FS��a4��K�X�V���޺�]i�G]x�ui�{	�i�4n�r0��;h�V��
�u]]+���.�9�\w;�h�Gflmr�Bu�(����zGc�n}XQox���rZݭ:�������nD�������_���m�3$�m�ڲ�u��)���q�ə��m�%3��:$lݰ�bf�m��#,�ہ)�KQ�nHw	6���l��m��e��۳lY�f�#�d���om����{V�m�e�sl�cqjIq�@6�蓋+M�f�fέ$3+kQ�ptA۶��I��$�٬I�u�7l��ۗf3���n�iv�&n6�[v��v�9�ݨ%��-67ch���B;v�3p��Yf�ma�X���M�%m�v֩5�m�kq���	ͳ�G��rH�1�Yyokֈ������gev������Em�n�62r�9Y��Ҷ�9#"t�[sfkkN�1��E�����d��\����{�n����vN�2Ӧ�쌳��܋md�ڍ���R����$GIei�ٛ���,�[Y��mM��q�����ɻX�b�ݖ�=��M�98䍻$��kDRt��zׯ5�1�ͻl�!="z���@�gh�	o)bC�W�����M95 hmظjk� ��q�/�G8�I�Q�~�1�׮�]�O݃Hw��9��&H� �@�O�u{�{V����O1�l�-�ˍ�Ρ���~�����%"�t�G2�������$�E���l�.��79�@���r)�Q,t��\f.���ƥ�}�����6_�QP	6/�4)^�2UA}`�	o)�o�Wc�=YO���k�x�: ��R �""��7����t�-�̚�Р��/�G8��{�{+��1̦3vI]�7!��TMJ��4=ݫ	�PL��M?>��r��x;���\onq=�@��A���H�􈑗wE��O�<�G���$e�QI�Я+��J�/�l ��>p�U�y��u�8W'@��cz�ln�ۺ�ՕAso�dm�{7X̢���-�Ho=�)�j�����7L������;�_A͋�3�	����$a�+�ֆ�n��AxB��x]'Σ�wq=�=���1�bS�2��Wr�j�noǇ��_ޭ���e`�4�1&�v(mW<[�'W^��r�vd�&�(��"�D�ۯ��L~�A% A2D��9�����{s�����~p2�T�A�d�2 ��6	��qi)\�81�����n�FX�@�iR��U�<�
L�L�!���Y����XE�	�@Iω3@@�	�d9x:6pN��i���Z��$�es�1Ϩ7B�Mx� ��z�,,�{VdAҐ?I�S���+8W�e@��z܁�<DYG�x�>��� D�d���DI4]z�����E�K��Q؁�
ҥǞ*�@jEA2�?Iw�
���N�s��e����0���A��x����R7�ə�JC���]�񜕵���
�P��{���4/j���x�LUPa�T�!�8�G��p��b�[8�Kr8ye��v��������nn8�5yJCm��A�!Z�U��([��ǁ��|d�ӻ>�ۆg�h��X��=k�K�bՎh7.��"c=y�S����UUj�g6����Z���7�r����9b�w���%8�8)q�铐2�v�^z���wE�
9�ۭ��M���[�O�'���-�3f��5�ؗ��N#g1:�u�,.��:�^�ۿr� ���H�(!�w�{�_���7�ص
}Ƥ��>�[T�țA��?��#% ~�'�5�t5��H@�F�W�Z[Xɗ�Zn�K��t�Na�+	~���8�|/��������@D�"$�?��~�Y筌��W�MQ���
ҥ�<U~�P�q)�ww4˸;ٜ�(�.l��̢���dR��tu��uzOQ�~��H�����d9Yʽb����W�U�A�&?H�2P���Uc������ڱӅ4�華��*�B �r(@���H�(�)�d�`9�(Sj���tww=���ӂt4���cn8x;)勷5�;������ÿ0~;)�A$�?��百���9|&A;'WǹR��5�{�� � �� ����A(��p*��6пڀ�MeZ)�ש��+U�<���[����cgB�V]eX�\M�;Gum�@��b���X5m0l;=�)�(�V#:jy�����U�<J�u���6%�ݒF]̛ٛq���;+���_1")2D����N�mU�m��%@��G�܊ 6����"$��3:��>�[wP�$A	W~�M
�y����[I��K��M1ܾ���ؾs���1�vheܒ7%2G��l�&�CQ��@����c}*��%G�5���}A� �w��(hZ��]o�J��E8�$�JPv��F�]�v8n^�V��F��L�5�	����__��������d��w��ޒy��cD�dN�U�i-1��p#țϨ�"H� �H��ڣ��\�P���_�*�w�*��`�0�)��5�p!�2W�����P���i��A� ��0�2R�_3^��R�(�#���r��1�i�ڹ�sP��v6��kY̎uD嚡�>���n\�5��E�W'�N�7(l�����B˽:IQ�ň�s^�܊	5��5�gڞ�|�vm�x�P�.hG�5q��sd�}\,��R0�[�B:�&�!������}�@7�DDI�J@�$A$Z�le}n ��g�TX�[I��ˏ<Ub3�gx�T��HT���~6tK"�ԓ�s:�eK��3]�l31��q^�Zi�[�#��߾���2R��"
��yK����ɒE9�ƅ���U�zW��@@e߯�	A d�� �"`�䪳�W�u��8�Ғ�K��7$�_���
�mX�&OL*�7��C(P36ň�h@&E���	�چX�C�vWcn�}�䇳�x�뉀A�A%"	�&�!T�ɸ�XI�0�D"]��1���{����u���5�:���VM���8�.F�
�������]�m��녅oF��J/6**�no_b�h�h��R�Sksv�)C�MU*�ȋW��������A|d��"D�#%y	=�w�R΃�? ��i��9�̗��6l�T0��P��b���"D;3a�U,��:��8d��E�0Ż4�b�4I���sy�u���[�pc����t��f�AT+�	5��4+��y�����0�Q��Sc�Lδ��}Y슄iL�2$A��[=��G�~=�Bx���]�Oe���$�������
	<-塼�곩����f�)׬B���$��1�J��gy�k��*��)�!�b��@&�"H���j�������A$a�@&���h��7V�aj2�=X��>N�x�d����|�H�@�($a������o�����B��dr��]e��%G�s��jy� �����ys����"+$\+o�%k�T��{{+��]�d���W��E��yt��AK�x����U���:�fM�ݺ��| �`)I�)�2�e��9R�E(��V�/k�k�q�sb�2{ny7\u؎լ�5�
k��p-ʶ�ͮ�A�GOkpaӺ3��B���Ď񎻱ۮv��/lu��0:s2��g�0�%՜ŀ�Wg�k7F�C�nٮ����i����J̖R���y�����-� <&�Z�tu7t;�/��ڝ䕌��e��~߳����Z۶
1.C���˹�<�"��j{V1u�]�۩�
3�����q��O�'�#% &H���Ovw���jqE9��Um&��k��f����D"H��K�:Wޏ�ǩ.U�0��@�B��sR����aj2�D<5~���3��0*���t��ߩ����i�A#wt�㩌���s5�w� �ދ���:�����˹�bc�W�A$a�D��*��h>~|�s��PF�z�"`��=���3����1~�u����n��l�JC݅7�H2��)�D�a#=T���r,;�JW�r;8x����y��g��z2D�ju�ܳBd�*�ѪS5D]��w\'�x�]�z�X�v�]�"�c"t�g��<� P����4#+[;I򪭣�o�{U�v��\B�9$���)]�)ܤ"`���ۛ��m�;Vg�b��FF����IWE��S������x�Z:{B�~���e��zw���i�ON	3�gqvҟ]�#�Z��J�x��꾳E`�~�n@mP�&d���`x��6�D_D�K�D�F/�Ȍ�T��m����ީN��Gd�;����&��$��� ��he܈'bY�[v�PdM��K��/��w�.�� �f���v���/�)FQ^�G�[@n��u��H���Q�T�p��XE�����~�9�z�a��� ���2W�D!M�<gu��]lŋ�l ��&�`����lm���"�z��xϘ
o�v���K�r�$��"	{7}��|��;�-&|�
��8-UUQ�4� �k�*� �@�ԁ;��̪}o�~s����f�Mf�v�Н;ǔy-��}H}� D�=;a��Q5i_��*9�:�Mx�� �S��NI�|L�lj�]{W�,2���qNl��:�%<nb`�sVm�K�����u�[��;��+{�Z�����i����o{yB]�q�6z�J�b�C�t�{�fJ@�$@I�r�V=�Z�M���**��M
��ʅK�)9Gx��ˁ�Pw�PӢ^�	���"D&Jd�0d�#	CD��-<��t'���K����|��c���KػY���< �WD�G��slh��.�$КƛLf-�ݝ�z4��m��� ���cO�١�m�)�ı�wsI�/�|�����ԭX��LE��S����lt�@�#`�%"=O����U�u�`B;^��U-�T*\�I�;�-&X����@��x��2Lniv6�}��vhg{!#�1�wJ�:2�D�L�	.�o,;&�VSb��yG��<o���}%���ZbU����i��;)A�&]��g���]cY9�(x�/n�Un�:w�*?�;�ըͫ��m)���q�=x�<�ʯJF쑚9�6�ݣV�K۞�q����S�͇�'ԬA�H�w#�U�[n��^"�#% A �I��l���t�~�­\*\ђw7�뒼?_�D�� �"�'ի���Y��_���5h��ƺ�D����
��S8�Vf�z��M6lk�k�?I�_��}6/�LЀL�[��b5Q˸�%��Y�w�Eh����J�����ؾr"D��Jww4ə4���-�^{�4�~KS�.v��B�C�r(@�ՋL�"�NU	0d�X�@��������'E�	��,W1�;}�4g���/Ѡ��f�͹$wq#����r�8��xe�Y�P�A��3�����ưi�j�<V�b1M�V�+|�y�F�d�A ���"�%/+��L����-(V�wv�}�K�Sy�<7݀�ܢ��)���Y��'+�O;��Ixպ�4�>� ��r��oo2�,��}4��Oz(��ov���x�����Rq��W>�ðU)�N�y���1T#ek���:���Ή�5L�Q.��7ܻy ��GGz�J�2�?7�mb�/ߎ��	�V�VnQ
�i���N�Y�L�7T�����H��_p��������Q���U�T_��E�W��T����Gg)���P�k��Jyi���˧�={��.�%Mfe�uW%s����&�'�PQ�FΜ�C�om��S�+Z����%��K!�j��fV��%��oH�s��=��֡���V�^���M�QW-�ɶ���f\��ou͟%����/�Ⱥ����F��J��7G.9x�hIO�khҗ��oN
Z�f^D�]��и�*�:Ý�՜/l��n��ַ����5�t�ۖ�c,�pυ�%�T�\�U�r�:�͛�G*3R��]�a�Sw�y�sa�Ӻ�����B�-�YZ8N剝�:�[ڎd�W��Op�Z��v��:�k�2/"S)UaY�}�sz�Ś��i��mna�%Sy������ɹ{ܮs��գY�L�a+t���n�.�.S)*�R�0�̵anދb��'8���HrٻW,nW]\x�Cʋy��8�b���]Xr*�8���s;����f�ʳ(*Te�f�)f�`�+2[.�sJ�����ʬJ�����ӵaS-u�f<�b�mU�z6��d�|��oU�@�wuSz^h��C�Ψz-Gsv���!Q�A�[����#�,CS�=˥t��u͛��|����}��H��,��:p�%��g[F �3m����3Klt��smf��ݖ8���ݹ��kf���o{b.6kH��g�
D�M�e�%�F��:Snlq�3�-Ў�ܔ��H�h�i6��X��Ͷ�{v�K�r��)#m�ٻv�ͱ���;�8�rS���N�
��v�pq�k[m�Q@�t�(�s�dI��$"���[f^xQԝ������ S��T] ��RJrHw�h�d�܋ڱ;�ڋH����C����&��gx%c�q�Q�$rm��"vj9JA!" 8� �(�
v��t,ks���n��s�-��{Y�ea�9� ���B�A�[v���Y֧nB�rη$�ےOl�yY�k9	G����b[Y��>h��0Ԯ�f&�tv*_<��͸�LL5��&u��!�
me��r��p]Ϯ�@��s���h�΄�pԷ]��$\uV�qݞ3���q��<v���ҍ�x�nF���6&+�m;KcR^�u�Z'���<��Yݰ`���qZ;!gI�Ħ5�Ǝ�'Q�j���rF���/K�s�y��؏`(:�	�cZ� ��v���:m�α���Hҭ� PV�`Ck�;���)����V�����K:�w������l�"���e��	��e#�®��>܋��<\��r��&z&8c�n��/Dgb��˱۬Ik�R�h���f�*�O͎�z�b(Q�:�/��]7Z����\U��6�w'���痏Oo'h��\q;��qǖ�k�m���7'<�gY��@��6|�W���t������s�*��;uO(�c�]�M���p�����Q�gJ�΅X݃L���ji��q���IB�ķk�i{'0�l<n��^��@�+�V��0h`;V�c�s�<�{m��>�Gm�|umV-�
Ԍ�BR]pId�J����F�{nfl��]&h����7y���[p�tqc��`�;L̙�-�q3�t"ꬤJR��h�]���v�c�4v��	Ȇ���wl8��+6�g��.��mk�1���2�,bLu� 9�2u�k4�零.m)�n�:�n�.n�1�|�d#�@������4-�tĥ�yS \Ÿ��i.q(Ԙ�c���.����H�M	t1�t.�Q����D:�:	v���ظ�l��*��2�ȱ��ض��Pn>o>"����q��w<%�)9*��qȧkp��ڍ�vڶ���֌���P�Q����N���<�[�I��v��u��LA,9�Uah�N{TU�m�i��a�D�F���)5	t�H��h�e#�vv��.���b��[ ���]�M�h΅�Ꭓ��V���*N��A�]wS*���vqNؼ�.��t[��/<Qmqv�����`��g���MӐA��j��Ļ��Qc+t{\���E&A��dU}���j�r��O[�n�r�z�����6��o�'*P��5�z�����:�瞸��x��Ԫq�u��\��A�7(�d��4a|v���`uc�<=�ǗrnC�G�vz1ԝt{CmjS6]ԩc���O��+aH\͸u�8-�7(h�`3dm�֦lң�\D��v(��~�zR ����D]���K�)�[��g��m�aڌ�g+ @{B��/�"dH�?%�y��M�L��4 @�B�m�\v�:��k"1O�5B� �mԝ�\��x����)@;�H�JH��^�d�Һp�$����=iP��ǣ\�^~������ D������l���U`"�'��СOY*).|����ƌi�6Q�Ȉ�׹�S�D���d�eľ�� ��W���\�ݘ��<K��) uq�K_�Db��� �E�DW��=��x_�UP!2ڣIP���.l��Q�� �L:�qa����\.�S3{�����L'�/��� �$L��ӷ������B��X�5��%��(B=9vR �Dl����s܍f?��uy�;�w��r����(�;�v��{���ɆU�)1����w�WE�v���TI�ҷ�,��,���N����B4%s$*'��sI
�e���zٯ>Q�J��;::�\�W�P_d�3% A�E�)�X/�V�5�t�9hSF5q�+X��sB�N�� ��@:��H���7�[����njxA&�(�4��r�oM��B5���@f��ZM�&�4Ϩ7B�X`�% A�D"I�MW�xO>ϰ
�*�y����M�$*��"۫!�2W��/�NF��!#��	F�q��[��3æ�&�ʖ��[���=�.�i�\h�OA��}}Ad��� �A{����M��T��v#�Nt�G)ϐ�@$t�˹%'w�;���znC�̂n��kQA|m|�����7�������z�P�b�G95B��ټ���e����7�A��D@�����z4�ǯ=�ޢN���'_.��֟l������oFog^4�Nm�j�U.�l��Oi�Pm��`�7n�7J��mS�5d.���!6t���\y�[4(A3B��H�C<4\�9�J��.0��5	�@W3���M�|�y-b��W�f��F��0ض8w��Gr�%"	�&"D�J�'�_;��c�/��Yo$��9W7��ʡ�@�r*j�e` �"�\s��[M�P�m�TCB��M�T&M�rDn��,� �>¦��qg���~o�>��h@�� I��x�)�DJK��gI
�%����]u�!��dT34&H�"D�Pmr�m�.o7܆�h@�T*��en�Y�VJ�%��G9@�u$��J������uY��dСϨA&����/'p�T��x�U���ܼ��dc��#n�;��˸%$B;�7�_dJ� ��������O#�u����]���������|�9õb�=wqJӍ�n+y�������hN�;x�{�w�N��w��vU]��Db��nV��Qe,�{*Ա!.�9Bu��#�HN�'� ���A AG��ݖ3����2���3hP��2�i�,Ϋ%W����r�#܂"H��ȅ�wS�';eUW�����-J�bYN�c��Q��WkvteS��m��DPu]ZA�����)�����.x�U�i�¨F�C#�8ɽ$�����u��"��0�2RQ��U|��Qӊ���^�#}KZ"d�3<� �^��ɑ҂ �F��9t��;*�F;�$c��Wqь^���\�O���h�,��%W�����#ܒS.�L��A�ĲkM�W��o(A��Dd��Y���񜫺=}�P�t"9�����3l���	&|�2R �N^�kr��Y�t|�GQD�$���]$*�x�z �2R �d�+�]�z�)�YU��[�V� ٹ��s�Va��^��2	�g������=�{�Oj۫��Z/I�ן��=��][���5��#<E���c6��we��&�*KK�h�Q3�2���.�/<����U�H�q×��	s�<����ӧ�GhԶWQ�a�&Ѻf�
D���%ն���eۭ�d��cN^.���1B��T<��u2a��hGYfS��\���.8ywL'#=A�A.�ʈe�3W��F�@�UZ����(-v�S�x��N:ꀎ������4��_�ߑ>�e2*�	u��Q��$�����܌#sl��16���:��_#��G��#e����pL��4*�<�ݧ1���%W��b�N��B6�Z���"�H��2-1ݾ\��޿1������gy��9wtz��9!�9 CjŤ��ܖ����Ͳ�d��ܕ�e�2H����L�5ms��ɢ�M3<���ۯA��0#��J��H�P�9�@��K�1�J�Gz �ߑ���4%ϖ�9�*Q*�WW�K�ʞ�u���ӂ�"��?��/����H� ȂJ��2��Reh�7C�v&2�I���˻�ݘ���G9V/�LנA(h�\E�׼��FѠM��5E�Js@�f��i��:����j�X�GX��6����-��D� �"H��P_.�t'i���͇��|��b�e���Y�� �P@�R?I��(#%E�fM}���Ϋ��V�v������~�:���Tն�ol_bL!G��u�8WYy^6��ͼ�Q/p%��۱C��ۛ�G�t�!:���v�ƕ��^+���sC7 �]ߎ�w�EG�sy�=��D��J@~2D��K���ߎ�BYƯ3��g.�vbV'��EV�J�	DI{�������ZF�F�/��%�=����:���AmՈ5�N9�����o�Z���]X"D�PD#�JV��cyXyPv$����w3�%_����sP 5B�	#�$A����G����I%D�]:&��8��`���m�u.D�8�6�̻J�����O� ��s�FJ@�d����m��ݻ�b��aڷ�i.����B�a��DIA$ld������ac�u��ЪD��t�t���̟1�\g�̋g�kޢ8CJ�@�T"9ȯ@$�`�H��h�z�v�'I���E3u>Z���-�U��ۡ��w.h����gb㺟5s���(Ս]���}��;��cà����+#�'�$���D�P��W之#����P	7~�k��z�}.���e%�ށ&���� A&��i-��.��vbV'��	��e6�5��m|�����#��� �(P�I�<�Y�2k��P��ȆWQ{7]�g+�� ��&G��J@L�m���y�*쩽������5�T�DЦM.4>u;�����^��ĖRh�6A������ї���+� 2�_���4(SG�Z�4��Ĭ�\�R]���s�B � R��^��������k{�T��H�_P��� S�{�+��ˣ��X����P ������X����B�N��MD"H���"��Ѓ\�_���!�^����Nd�x���
��f�@�"`"���j,WP`���k� hW�,�u�\B�Vy.��s�D�y�`�6��8N]J�r�k�Xi_/d̢�}��u)j��^�_CU��v��oݍ�o�7/:�����d\�����mh�#}����?$LD��f�r�j�n���&WC}�o/z�,��#�\���b�>�h^Y��Q������İ�J�8(b���Ƿ�9��g�Q�Ŧ�g�繥����Y�~�t_�B�3�Ģ��6�qS�,@��{L�}�{ix��1�/�#�$L%d�-A�?z��y�7��|��u���OIq���<ň�sB5B�	%)�癃;o%���������&AС��$�r�}.ai�;��\v�S�WC�z��s�J� $;�gu2�Q�{� j�{��hP�w��+��=kG=���*�OujxM�]t���a�H��(#%���~&L�v����9B{w�'�;�TA�K<�1~�5�� I�o���{��7&���j>G�����Z�y����+��w�\�BR��%1�{��]T]72_v�e!2�U��+�Ѥ��M�YƵ=�`��h����Y���U@$[l!�j��cn"�6� �t�M�*�n6hk����e0-��J1���X`hM5�rk��l,��$��`p��l��З�'�P�7���<sk:��mÍ�y7S�^8�O�h�V��R}��ػcb�H��K�ɋc�c��,�B��ʾkJ)�t2�S5�&�Ws4.��������VY�1)V�3Ԓ��ŝ�	���ڶU1rv� �6�"������:&A��d�~�!���!��W��V���B��%�lى�꧴4�lA�)d@I1���6\Z�Є���'"�K4�pW=Bz�o)�,@�y��2ë��"�C�cudn��2P@$A�%|��wAܣ�&b��-���Y�\A�K<�1b#נG��G���_)|~v�^k�}9`�jԈ "g2v�p��>w��ih���Wd���ز������A$A�% A $��!����$oN�k�z�o)�.<�W���"�>���^8���a��Tk�AX��6�e8iԡj1�U�^�+Oq��߬%�|��wi|AB�>��)��'rG���/+��l�y�_���{T���wq#�&R�p�%ש�&����P�>>��M��n2�hc���7g�f�I��H��"�z�WT'��Gt��|�rĶ��\�mӆu��)V��">ؘ9��j��y��ih�t Arj��	��u<������z�,ȑ���Ywt��	�LʚN�v�kd��<�1�4qR��~��`���d�A �"D|n�2r/d.�q�i4)�6��q���g����׵�"ݾO���ݔ��$��$��ʢ�U�9z�sN�r�`�n���Pl��Υ�Ec�}@!�s+�"6�m悦�MQ���b�S��I�u��p�u� ��-f�ƨV��Je����y9�zR� D�����V���+X@�݂T��#�z���q3Ճ�I)�Ħ1�ܫ��WpK9el��S\#'�W�I�PW�����qpb��K3�P��bS�$���p�T7�WU,�U�����4�]ʻ�1���
\�~����oҶ7��\w��/���fNʬN9���.��K�b�|{Pn�={������Ng1o5S]��輼W��&��ȳ~&U&��8��g.d,�VG"i��11�S��.��$��gϾψ��b�D�ʦĜ"�W\���5uo*��QktDx7�&�}v�m��rͩy�ڻ�%��U����zGE.gݩ�q�mͬ��\����5T�����:Sz��9�+p�*���s~���Ǭ3x/�Tpv�ޫ�����wt"#�v��q��}W��n���{N��d��<���6��P�86�o)ϰeiuOZ�'j��e��Q̺��U>�s�TO�,32��V1�a�b�Ҍ6��c�K��\����m�]����l�j�]՘Ɫ����ޡ0M귉��Ck/�of�au"�f�8[�p�M1��5>�̧��mϫz��Y[�U�=7�E:}���8�G���c���lB�<7ʫoj if��Gt�Ð���)�1Fj-9�9ƣ�ؘ���g5�R�a�)<f���ٻ+��#gtr��a�q�;N�

f��1�_M���2K][�,�G%a�4|�Un��d$�Z���逈��:h�.z6�]��v�A!��W�.��3�����u���]���xs�ZL��^�/�����G#�S:���;��
�ڂ���y�Tm&��dDg1ݺcI�uWV��-�`��O)�4P�5�%Ir�ۈF"хi��}�3����fk�|�8,�ș�y�p#�ӊ�J�ڳ������UĞ�u����Q���	��A�BlR�mξ;rJ�#��t��$'��T�kÜ�RL�)�sj�m�E�i ��K48��:Щ88L�9�+2��A�v{X%�ض��[i3��IG{a=���"��N'@�A�$m�@��qm�E�K�s����u�vs�qC��u�GIqE")ĳ�BH%�`J��RIݻ˱��l�Ӂ�BG� �t�G$P;��$DC�+p�l��� 9�dN�۱�\�e'Np{vr'�k-�Gs�[XRN�9;k';73[t���H̐��8'�Kj�C���N9�P"���9;���:N:$^�B����#�r��� �;�NJ�s��q�ppR!�P�t����;4��4Qe����s��ֶ�9@�^�ok��
FݔOk{vM�)����(�8۵A�K,D�k�}��j�y�Աh�t .I�r��u�]�)�wTF*�ۍ�Vo(W�]��Ъ�\]�Z����P�\���@}�Z*�[�8���^$�� �fJ�}uN����u��Z���_U*��J��?X��@j�2/���fG�Fxi`������uI�G+�Z9ݜ�;�ӧ2y�b�\h���V�����߾8��^��P�g���b�;j�s�b�Y#L�f�B��n�FWH����w�#��I)��y�W�4����U^.4ʝa�v��[ ����/�����yk���ߓ#ڐ'�@)#�J��V�_�ֳ.���J���w?�y�"� ��/��d�C�u�[�/�R+ �z�>�@��Աi�y�<qh�b�z�/b�_�[{S[��M=�>㘔:^�c�ӭ�1��-�>7t��ג`����.�x/�z0�2���T���E�ݭ��=ܫu�-���@@�q�	;~&P �_$��>���A+����sÃ٫6q���b`�� ���&lE]���^߯e�#\�Q(�O̔]U
�s�C��ӹ# ����Tv!nmLWEmu�bQ��$�}{z�ظ&k� B��>X[�<��ԯ�,���"��_a� nH]{$A%"	�&F�g�4��q�9�,s�N�F�(���y����V�D /ta�%v2�$���XME� ��D�����9�ʳ�	M���9Ã�Vl�ҼA�� �yd�~�'� �]�k�/:A���@�
v�,-�Q�f��W�zԿ@�mcۘs�:q�(��=�~�q�B	� A%?�2 �2W����ۼh��5 A��7�Hh�͌En��Ar(@�Ѱ̔�?	w�ɛl�ie���F�aX�����s&�<�������c�/��wj���-�ɆΤn����p�yΓ�0/��A��o��{�
�<�K�]Y�	��ѱƊEՉ�f��wh������7Ů'�s�ꍎ)ے��v�Р�l	�Tƙk�R��	�6�Զ���K�X��̽�Z�`:�hLښ�0�v�pڹ�F��s��E��]�ڸ���\닋�������.̈́-Y9:^<L�div�c�Vwmn;����L�$l�^ڃ���2�uG����5�y����S�&���+LK4�\�Y�u
�J����v�c2T"�nƻC�쯽�,�#�"�{�=-C�B���*��2v�;q�����>�� ��`%�֮�[�ᑻ4 %"���s�k��:��"�@7�@�=�"$��ɘu{R��V��qr��o�"�J�� �ӄm���Eݸ������͌En����#��V%D���}�:���p*�uK��#{��J	^�a�q�lY��J����ȴ��闞��/�ۼ���%?I+G��Ԭ�,�hP�d�I��g$�W����c����������.Y�]Q$�u�'���mOnZ.���]�z���7e���8��H�.����s�0A辒���2D3|qinڼ��V�~�خ��<`Ź�89�0vR_$|�2R?W@|֘i�S�N��ϼ�Wcl�s3}�]8*Ц�����v��9�:vIճ;�%Dӷ��Z��5��u��R\��5gUtUb:&3�5��B�v>1�C�B�5�T#>bڱ� ��܃�s�W6�N�W�$o��0��)�%��u5o�J��`ʢ�;o��Vķz����o!�oԁz �G��ȂJDA�=��޸~�Y����ޥ�X���A��W�J������+���׻�i��F��"lA�)dA	)j���k�֣w���/y�4�eD��P��D��׉��j��K�j=�������/X ���nź�Q�J�yɹRkcj�ya����qx�"~�ﱖ��G���_���4(+/�6䚭gd�W�܁��y��j��b��_1"�H��&�w��v�;���J_A݊�o>+Po6���ҷEc"�P �a�%C�y���/��͂gW�H���M߉��Z:�5��x��=�o*�����md��ghh�U�O�:^�,�v�I\r�2V4��Ni\�]@ъ7'�$M��[;���h�-�*�D�l�ҽ���� �� ���"dH���r��*��������IX��;/�|͚��˕�������Z��T\�F3���d��Ħ��U+�$�e��;�b�s�^�k��+Po6���ف_� �PDOD�� �"c޻���m/�
�<5A��6��j�p]�÷jس�u�Mv��]X5#LM�n{�>����e�>��Mߠ�����\�sx�FX���U��!���D�)H�P�	�^��N�z��0��bϫ�
��7�٩�f9r����b��С ��:�4��n���:����O��3^�k{*8��ӽ�ݻ���7��/��Ȩ6.	� O�W%S;�[=<�
����<M	d�=��C-q���J���&D�Ϸk�G��n�r����G�pV��i���Z^�퀉�X�(������50᫬�䥢��f�^�ps�Wp�̹��ɥ8�{~�4��L%����$�0d�W�;��uP���$��5;l�.W��}H7�F�P�º�IF�p�@@ڄ��469�]��P�ؗY`��ZR�ja�)���pnj���#%"	�!���!��7��/�Me�`��a���ڄ�@I0?��Ntܬ�h�a����h�{�pW�l㲀R/�P@�POQ^��[Z)�m4�{��ҀBH�J�J��T�r]k�5;mG.W���5: IFJ@��+[�yܸ�A�j�w.8�ov�f�J���At�ν�e�>�_=A$���	�^�I��2�����������[�Gp E�W<�
� h2�N�:!U~��]����󪪢"�N�Irː.�x�R M�J�j�P���V�`��	N:�i~dz�i������z��C����#ٍ�P�j6i�[�򁎍����\k��ض�F5r����w=2��9q؇it��T��U�u�b��"�`u3�y�w ��.<�Z�^�Ő�/W\� F�4m�J8�b�F�mn�X�=7�#�ݸ�g���L��z�at+kc)��å�%��[N�K�GZ^c��A�R-��V�R1D�4��p܏^sJ��uu�j�>����Hԑ��q�P�]I�J�u�s��ךI�͹��tV�Zv%[����z��F�?|�b���4(S:�o�����+�Iض��.��p�nV�����"l_IC��"d��ze�{f�G�����5~�g��ݾ�ЉY���r(�'�)�s�ۦ��b���&����	_$o��i���ߛu�=���ʷ��3�"ҫ�B	�P�"`��e��9�0�� A��S:�o���x�W� F)�&���f��PWwU'�$��%1�wr�]�@�I���ݏ�`ә��Y��x�ُ6�t�z� L�A��3% D����E��ɳ�6aͦ�%��A ��%���!%8ƫ on�qȵ�V����V��o#��r`AޤA� D�|Ĉ/���{һ��S�Tj����cdK�F�(��z��H� �2PD<ث==D/:�FW;O�J�		Ҕ�qt�l돨o){P��{ح�N�"�"VA54�wo�w|��mVY�u�oZ����<.���f������s�t���R`X�F9��B'���ג����S�����y|Ĉ#%|�2D���x�G;��{١���"�P lX�)�D�
���ޮ8��݈(U�� M
g4q%5�S�Tj�1�45�U���wv�D�^��e�����"�^ӝ�oN����A�M��7��#��Rb�z1�zy� ���" ��%]Z���[	:�F�!���n�)6�v�H冷ENgru��,:�&o��#�Ձ<�
�dMo�Y�qK{���+�`P�w�us�ƨ�����ψ��"H�IH��6X4��'V���v����8�L�FwT�������� �u%�p�j�x�ʿ@n��O�A$_IXA!�����o{���66����j�/.���M��.���6`��r��S4��(�T�F��x1.��y0)�j�WO�����oJ�]��Rv"1��hP�I�Y��*�p�\}�~KH#ڂޤA��+���-wnvhD�"�C�"�PN)�E��Cs��fψj�$�L�� ��y��{���zj�i�y&J�Y�{'������=��JD$F<��OϹ�����m�U3e�����ʛ4��.��b��Xc��&[3_4Z�\ߗޔ��a�+���esM��:�N�_�a�y���zr"�ےFnm�w$�����h��r���JŞ���lLmg�8;�ɛ١���B � G�6,A3��|�6�'���(g���o6�rJ~�)1"	�Y��Ζ�G�{�;��έ��:4�٤�n�#��)���w2w��m�9��a�Q�4@�v��SB M
�sM����NگO��s����Ⱦw�ĭ�Plq׳�"�,E�V���d�o-j�u�V�n�mԪcq�����Z�=;amRI)��o1<�$�C#�H�[�w�6R��7���o ����d��A��]�W�4��������;١��B � �pL�"3�r��2s���2�i�n���i�'�1����؃�H1Ճk\����~��K/߃e�B�Mߠ�9v�SI��;�F��B�"����i^J��Τ?"`�_IA��%�r��q�g�vh@�q�^׋�ot���Y�/�#ю���"I��:���c �A)	���H� �H�$Gc�#�<w�}6�-��a����^1B u�d��hTMة]�v�yʻ�g=�����Y4+�lqE4���[XTj�����n��5b {iA�ɑ"d��0�0=�h;=j��w�H�8IK0u�-���W�y�$g��נ���%�hB���$�	/�@�$�H@���I_���%�HB��H@���B��@�$����%� IZ�$ IB��%���%���$��B��H@�� $�	/���%�$ Ix��%��(+$�k%�n��|�k0
 ��d��Cq�   5  @       U@�
��@  (  � �@
   � Р
"P� �  $ H( U�(
�� 
(@��UT
(�� �@(J������=UQ��$�R�H�AAT��
��!T�
P��T��RB�%)J�@�*�P��Q(�  w: D
�$� �� W�J��TUwwT���*GvrUp�tI�(UwwH$��RW,�E��U`�iE�� P((� �����K�太Ң��љ�(͔����t��[�$��5��t�f�w�u	R������3�l�٢JT�J(W� �� 
�"�"*�G{�i��P/<� � =��P���  �g�Rx ,�o0��� z� � A\��  \�y
��   <�IN���EB@��|  s�}�zI����=	W��I��R�Nf��L�֐�;�t�E8tI=�S����i[�%)'��$��h	T��PP��  �"*@� ��� ����}n �Tɨ*Kݺ$H绉��Wt^��{t!*n�zl���lU-o;�*T�<+{�Iyj$"��P 
���   mC���/&�J��T%wT�\�J�������Ts�������PnǊ��`9��ly ��UJJT�   <��$�P(P�T*����!� {���(�`�z  �<�U���A�w
�P�c�+m� ����/g�`�(��P( P
|   ���@ww{
�1ޒ�� w1���� d�+���{�*��@!�!� �j@��JG{� <QU@J�(>   ���*PQQ)D�J}� ;��ӽoG�P<�vё9��p�� �= �۰hv8K���U<��9�
��*��v��((W�  ������%`������#�W:�J�ra�;��!� x�~�L�R��  ��i�R��  "~MT�4���  l� J� @��T�h`��&�Sm"�B  �=O��������W����]���}���&�Ì�Q���Z���<�HH@�p��$$ I2 �$$ I?�HH@��$�	#		yӷ��������dէ�7v��oQ߷TV����t�
ⵥ�!n�t�%�u�r8V�зP��K��da�uf]�i��J�{k>�#�H]*nЭ*!�Z�c
[����Yܼ�U&�N�pDS[���2k�ϩ��
Ge:[5<�ʙ��|Ĉ�B)�_$���}����XL��p@�`���3�n鬭�Al����B�������{.���{�V)�2UV��oo�t)ek��,[[�dp�Ԃ�ފ���kk)�eK�����jY���J���J.��Q�7BR�s8�t��ne���pf\y���+p9��P�d&%gm�S�,�2�cO��5�'	�-�(E �f��D.}u���u��kJ,9Xͽ�:�!Uc%U���FJbؕX�؁�3X��v0TO$T�Q�0b�)� VW۔�ZJ�v3u���SLh"��p�ʙb��N}n������n봚U��7z�m
�Q��hK����l`.+(^1����SDf�ݗ.��,]Cn,�5���ǈ�[� D���l��*�2���Yt��X�E;��eS�rj�\�i̺����b��h3�N���3n֫�{Oe��;g2��ڭf�ykFi��)ؤ��@�񌹻���/>�ɊT�/)<��+�ܗ0U:We6h�M
�o,��wc3a��M�h-F�MYr�짯h�zh�4��*�R���J'�[;�Vn��j9��"�-�[r{Or���0+5��۬�O��b�Zه[���/jۀ٧�iT��o�ך¤u�q�XU
�~x�	��j�v3r��R����Р��+���b��n^P�yt/����I�h�gCX����5g���vTƑt��R���X����E�o鈸�ӚC��J��K��%��4Un�;J��97,�)���wf�;WWjL̂�N芻Sn=9VEm�ƶ�;����mƥh�2��j��n��n]J���,�,����bH�-Z��ܣw��&4*�l�X�����6�e� �c�"�����X�4�ۻ�6=�g�����{S2�<U(UB+T˭8�w&�Z�
(iZ��{�����5��YB'�j&���C4�T�8[��C�cs.45��F��)��a5Yj��i��+k��Y�piV���V=�p��uZ���k1h"S�8��JW�)a��
�
�E��T�	]<�:�ԧvㆪ���ݧ����Ǖu[F�Y�U*��V,4���wi�N�HYe�$Z���c�U�-n捫ܽ�Vż�RhackW$SqU��eJZA��0Br	���eؤ�J��,iV��i+���/�W��4Q��J͊���%V�LYG��Cgv��iG���%���捹�'�pj�kwICe
ѡ�jn�t�
� ��v��Cnn�aFꂪĉݴ�ꥳ1�Bm
��o%���[�d��D2��uI6�p�[��Ŵv��б�.�9�۠�/�Aŋﰐ�-��Hӗ����FQ�L-���a[v.��9�m����ۼ��ZoqDa��ӉKu3��ե�V�5���\����R�� ���*��5�EaфeM��]�a�m�N.����N���x��rˑ�)˘Қp�XF�#1뢳lT��f9>�+2�u�"CAɰ(vU�mI��K��q��,�Y7yu�y�d��ƼW*�(7*f��7�-�n4�����(b ����G*[#^ܽڼL�`0fr�_մ�H�,%�boӜ4LΙ6ţ����B�v��ldr���7r��r����qb�v�뭇,#mbʲ���vJМ�U�X���6k�b�m'��y�L'0�N��XM<�LS6֬R�跛�Ó��-����F4�#X��d��"�XwV��Oqm��նn��mD]��,_Q���0��XȪB�jR\�`�Z�.f�(�T1�[�� ���ᥦ��7lM�ܦ0C��a2a��B�d����i,v�Y��%�J��P�o>J�f�x����K+6��E��2���&��+fn[��۱�C{�h h�F�]+U+Y���BG�"m��`�,ȧxw�˖l�lȲ����7WcM��T�&���e��$�h�Z���7�Ff�`ݺ��mJ�ڵ�8���:u�hP��v6<R�tVc1_��n	���lU1A�v[�Ix�n�{K|�1䣥����Q��zA_�`Use�j����kktl���4�Ւ�M��["&L�b�v���Xn�S�Xk��Y�*}oq��N�ͽ"kʤ-��c�ͺ��f��Cf^�w2�X:Y@ժ˴1l�_7��y��h㠆;9yv#\X�c1�3�\��!�4w����+K�ub��ːY�C~���,����[�p�r���ƫ� &�{�BhL��ˋ(�5hnL��v��#p*a�ٓ^6�q�r`���dԯ%;�yx-l
b{��WAC��ɋ2�̩��U�/]��ڽGc�,��5�b�#n㔍e�{+�#��fUW�����]���[�,�ƶ�d�F�a��Ac�'6�e��[���ĨU�*�5���-�#�su�����7����{��Q�$��V�hbю��c�ʍf����sFa�0�^C)�q�e���1d�ͫM �f%UY2�ܷd�5�Kf㘒$m��]E@�s4G2�ܡ���4�^��V�ݪ+ilҎܚ좳�#�����e.�;9Ye㲮2wwe��ǘ���Uz�<q]���Zԩ�dV�.�3a��[C5mUc�JW��Z�3jk
���W�
���@����03A��&��ܡ��]顂�m&��	IU^i�B�z�h���U:���,V���ʷr2h��R8l-��	��_)�������ܷ�4����X��+����`�úN��7V�oS(�5kif�g҅d�֝H��T�2�/MS*�P�96��++n*��a�,=.��mk���f+�Zn��!�&�5�t�l���L�T]��G�퟊RZF�M���Է�m�p?'U�Q�f	��^^uB��N��K���#k5�,�iڱe�5ѣI�ɻ�*V0���B�^�eV�P��to{��+���؜�UזQ��tj<X`se��B�R�,KH�r�]3M�FV�V;T��Ӕv3��v(,�o+&��+u:���Gu���#�6(�a�aجw�դ�l:^�y��%�)��$ǳiǪ�^L�ɷ.��Bܫ�����.��(f�@�He�beψ�%�n�5�2գ,,UO�Z����]��ꤓ�)ֱ��U-֮\{����u44��J�sfa�ŉ�O���PMAw�TH�������
���KT�Z�$*��V�U|����4*�u�̥[�����"x(n�7�F�J�u�x̢*�%�+��;_cT�l�o��X)h�T�X&�n����7R�裁&�-�TF�fc�[& �9p�/oa�W�`�ToZ����[x,m�=XȘ«��?�<�h4l��ڷH�6Q
l�6�C��wy��i[���#/*��pVR����o[�b0��W�U��tȞ깶��h�W��u]G�%�lf�~چ�)jƴT���I'2�]f^JueݚF�#sj��UuxdִlJ�n,�)t���qT�`�4~��-��Y�t��q�M�J�U�ܘ�R�9��Ӕfe[�h���>�&Y�����%�Q<T�k+l[��`V�MʨI���}�u@�RGٶ�CǏHoS����'H�e��;�K
���^��3-!����u1���q�or�-�jU��̭��/�[I�Kܥ�oB[-(V�įjB
��T/�.YT���ʳ:��a�J�"������q�X�H32歍�gMU�y���ɸ+��^i&��6L�ي��5�U�Q$\�qn�6�^��6��b3^�i(m�D±��Ƶ.f��Y�X/PҰ`g&�w�X�g]�14�������5\k&f��M�2V�t��([�{[x���B�_*�l�7@�MK3#��lYmμ-��L5b�b�C�D!���?Y�UF�Ψ���ckNd��������(���kT�e��f��i��k�;��+1�x���7U�Z�.��cw���3vR�&H�e�A�%�/�
�c����D�z�f+ܽ�9�/ieއAr$L�Ǒ؁m�nIot��iK���Ķ�@±VJC-n���ݯhzҺ���K5 �2me�è]FB�Sv�Ly���9�w�N*}�wD�T�f��%�ZíN��Uvq�j�B�ct�a�R��Ĭ��t��÷��R�oݚ���n�J��*�n7ZeJU�P�F�6�a5G�)���.!�(+3NL[�-�kn���W��%j�B��U��hfS���ޓ���J�wlɨU�n�bQ�v�h��b����PeL��p�9a�[���EI��T�%�z�\��aD�����x��x�\	\���lHs�j�0��g#��&����XcJTI��=�T��
F�^�y7Q7�u�(7bhn�&���I#w"���$˄ZT��[Eon����dT�G+*�T�����b��J��I�:�:`�r-9wUD��m�Yz�f5���e+Nٔ�:�n��ٺ��2�h��e�n���k�TN�ٶ�ܣH���y�ƅ-5jYfHeĻ��r�]Ǹij�!b�S�	��&�S\��a�O6��+2�S6�O�v\:���Yzv"VVc[I�m���F-���U��:�XDݩ�B�3HJ���*�᭷�m,�*��>)��[�.L�hMKvͬ��8G�-w�Ss�tBe���z%��s{B�M��B�#Q!gva�K�Йwa��c(Y'^X�\����N�m�YO%��˺�%
�/{v+3E���K��o�h��tX&�g*��o#4�jU��ʴ�P�f��Twk�vwQ4(3F��w4a͕IlO3v�%�
��7�>;�f��ÎƝ,��`Z�r7�������3t,AZj�vV^�@���l^�n�kUK��2�;�hkWz�0:1�F�K1��t�Ɲ����{Bl|�fP��Zt�W�)��d�jy��de�ݹz�RZg+h�yX"�OV=ʬ�Yvo\�]XWyOv#I6�m��W�5^:uoj��U��-bm�ll��7mͨ��턲J�U��x�uc�*����5L*:\���b4���x�U�aS�˩�e�Иsj��)e��<��}D�1��Q$�~��L�7��l��EZH-*�+S�����*{{0Z�P�抻V�P�Sp,��;�WT�+U�|2��J,��t�f^�e��0��̧j��&��7�W�n��ӺS"�i�.HB[{��CZ4�ӇLM��n��t��]卻F�+ёKэD��R9�ʄU�vh�f�b�F��ږ�k4]Mzݜݨ"^nU*�e,l<�w��n+ݬV��|�[Ӷ*������5��mM�wW�1zUD�d��	7n�3������L6)��ʢ�:�+�����������xV�A|�����-��j�����n�F*Xu�" N�5-�[&��
�R�]6&��ݣ�[h�r�R�YE��n�e#x-Rժ
-��(��w{m�༙�&�ȉ��e�RDX��2V5.R����E起U��A�fVoB��v�\Y����ߑ�
��T�u���Tdx��=�ϋ���)����i1onƲ���K�N�XX����a�+����w�4�&8����ͽ��'�NZ�2���Y�����6�q�Ь��=��̧]�YqE��#t�Yi�Pk�%�sqP2������r
�������R�MI��7a�,�����vwiij�������F��E*�U�мL�(X�M*�v5ԵݫGr�0؃O��5�b�!^GusNvZ6�
��A���:�FR�]�7�Y�XƉZH�K2�Ǖ��^�VG��n[pAv��mA����,�4v�߶�mʡ�-6�T���-Z�X5뭲��3�Ȱ3��+^�*��x��y�{F�4E�c�E��"�=6�ڎN��Iw�;n��L�,�6��:��n�/=U�	w�4k˻���j�,m���A����:��R�vQ�j�U��r������ƪ�{�6I�Őc	u�,Vź�U�qG��:"±/>��ّSՏ\�hM�x�V6���3�L��U����~�:.Q�2��n��^��-�b|qZ9a�T��G.�<5_'t���ѣ�)[���J�6��X�1��؍k�/p�%=VŔ�{��V����l�ź�Q$՜%�7&[��f�cݵWF��!��"��Vk[!�(š�F�n��I[��!R
����Jͻ�|�%՛�O�14Eڮ߶�2XG]����88B_^U���Q�
�$R�n���.�B�U��z,L���Uf����.��4j0�kvn<�[OZǣJ���k�қA)��4,V
X��\�օ)`�ӡ�7�����yW��R�+;j�fK�ڪ÷�uQdisnZ�t"��nM��D���`����8[�XF�m�^�B��Yu�bp9Y+wwfڢ�-e��^k�jab[���U.�_Ҋws*!�U�j�8KoN浯�94���uw��*�)=E�j��m#��н�zT�ylQ;0f����,�x��6��,�ңU�����{&<�+5�K
�m7w.���lVI�&$�[��Hر��tE)db
���=���K]<ơ��Y��c�0ژ�U�dK�{.j;z��<��x�P��U �K-�8�e�bmݪ��q"d��E�t�]*�"��t+Fk[7�fN���*��%��J��Z���*ċq�F��ȭZ�R����d���{�en�h�ƍ���Yka�)K�0�)��Ӽ�*4h5/1���J�{g��5.`9��S��[�� �`��+Fd�k
��%p*�J��ދBvɺ�+q�5l��2�h��动q5��(�5.�Q�ԭ�ƺ̼�j�����˵F,��E�Y��f�5����F���� ����$��$		 (I"� �$�"�� R�! RE��R)$"�H)!�@P$R@���HA@)Aa
 � �$RB
B@RBa�RI�(	a, ,	d��$
I )	"�"��$I� ,����a$��Id��$��I"��) "�@X��RHA@RHH,���I(���	a	@����I$��� ,����E$���"�  ��R �$�,		 BE�$� I A@�B@P! ,�C�p� ����$����?�������ن��˫Q�?�����+�c���8m^YƾgՉ��R����L�%��6f^�ҙr��&尞�Y.l�\�K������[�Cw]��*�e�N¨l�W٥�:���y�+e��8'�;t�:Z��
+��Mً/ۻ���,u��}���k����V9NT)�N�L|kV-Ai�tM�x���{/9�=���:�gG��B��ʗ\xǆ��e�|1_Eu�r���U��WW*���J�Îrʂ����di�Vt�#t��B(/�����`ۇ��=	�Y6c�ýB�wNFqt�{�9�yOb��8{�Em���q�.�:��1�S�qg��cޥ/;z� �Ѥ�S)���j��r�m��r�a�o�l���]��Jܽ�c*@��)^�!�/wu|\uX7�=�TVjB��������s�:.�"�˚-S'�p8������y��]�#�&��#+�z�G��Frcv�b�kr<:	�2�v*W���6R�ņF�Z�˞8����T�3D�/i���N3����m7W��^bل�^ڶ�Z��c��ޥ:_�c\)'z�e��v�)�����h]r;��_.T����-'�f�����J�(ӽW�.@��k
�v����L:Du���Jf-]Z���W���=US���ӳ��}օ�Q��g�dG��qk�i�x�h!V�yY���]j]1I��!�y��b���ߖf]nC�����|��5n�|��U�+t����^em��&R�Kr�Ͷ;�Q��V-K6�Um�÷uX���/eey5uj�wx�lzؓ�}ca��������[Ա^hm┍]�8��[Vrq/��_���B,6\y�F���2�G�2�;׵x��� �c��e�m|��`������5�V��7c]3+�uH̱̥�ێV"������J��d_̎8��̛q�)n\��F�0���Xkef�f�i��O��p�H�̫]�:J�ͺ�۝>��S�UU�*���0[w@ޝɀ����с�$��4��x�Sӏ�ի9Dܤ��p6�f�1J6�u�w7��r�,Q62�S(��x�b�e�0�S4�����;͎J��f�ۥ5V7���X~W�3>�a�cR*]_�6��*�x��*��Z9�,��.d���gU��jBक़9:.t�Z{�N��v���ŉ���p��M&.�n�)l�n��fq��e�˗�p���>j�J�\�i�8h�K�V�p�/J�s�����e��0���:�SNP;Pw�K_-4��-ZY�n�pVn������]��\6US#v��KD�!w�ӭ���ҫF\�Y�C]c��1.[1��E����P�deW�ѥ��b$tǊ�Gu�����נ�	]�Z��¸�e���X�p|�a��/�H��vFV��x�.޲`�uݺ]gdvr�I31��ȯ�����\�sm�jn�s!�+�ؘ˾�$�F���`2�y��2�nUB��j?`<
�8_8�WG7i�'��z�EX�v���eX�$�Ϯg��Ɇ���yO��:Y��/fG����MS��*�ī�k��a�Vh8�4^[���87��6/�i�����cvR/g���+��hr��p-�񫺮���m؈*�fҙ}8�+�uz�
p��v�v�a��V�
X��m��������5puD\�Ý'e;坼��e�Δ�{�6�{0
ޗ �]��Ԭ̻��V=�hA{--aeg���X�����F��xq�����a�%�$�����5o�K꣚�.����:�hK9���u9�j�-��|7�"b(�5�O��3{0jVw:և�r�9�v����dcF���UF�a���1�.��TH�5W{uh�uP�ڲ��3xB�2S{E����
&��F�_<B����kd�U����iU���z�E�c:<pEa;G�,�}[.�rHt�\�o-�dE�-O:p�؂�F��ga!�XoW�@[�m#��f;�e����e�Y�X���)s(�H�຋k�ة�g1�4��8)��z�ײ��RD�b�
���o(P�ب*���;��EwJV�wz�J�jT4�Qt�Cj���k{_[;bn��׵��b�;yy[��[��X2���pw*Ӥ��$�����[ާ �R�7V��2LOHק&�����ܢL�/��*�O�:ŁL/Bݎ"݊+�t�0I�ŝ�f`��+�cŗ��z�R�U5y��$7�t�n�ˁ�����^�0_om��b��Eш.��v�ھ�3M�q���Aq����2nP�Y(a{f�JcڻAtɔ��y�������[���;�E��9ըq�z�n�C���d��Tfd!�������`�;��OgG���x�FY�E�\�9=[��թ��wN��l��3��OM���a�f7F�v����͵k��9��W�f�4��MqX��m�Cƚ��ۆիqj�
<4��_�����.oԤ��`~�C�Z�]�|�]��yΥ�ݴ�Y�o����O ���/�.OU�{�LfUS��^�1�[�D'W�*���z|v�w��n���-�:�j�Neq�]��!��Spc��\�Ug��[x&>�`��1&������dṸ�g��LNr�Ȼ]����а[�KvK�R&uٻ�U��>6y�u��ٲ�`SG��ӛb,�l��T�e�E�z��׋�+)-�[p�m�7Xs�n�t�\�Ծ�9�/��Ρ��Z�㞞��ԭ�XA��h�Maӄ�U�M����žҵ؊� Q~�*U�t�
&�Kq^h'p�X��k�eֳ( ����)����� <�<N,]���]���ð�&�����B[��z���K:�=��י��]��a�˶���I�8H&�i������b��R��;��{B�F��mm�˟o�!S#�h[�[1g�L2��EI&��hxHw3']Q�t&�S��͏ ��mV��<�ڮ䠺���Q��JM/$�n�FZ�i�XE���6�P�^U�ξ�h^vm\f�l:�Z0g&��a�\4P��u^����a�Ȱ��d�X�����y�:�yA�K�m��v��X{�n�]�r��p�u�X���e��p�t�(�;���t:��^�Cg,`-��V��SF���i�ur�U͛��wY�W�}L4��Z:��J!��t�aK_?��I<��e�cˈ��;�u��-��mD�B��CT��Ǉ���u���v�q�n�}Uo
��tc"J�-���:�V5�Xu�d:.�_^���Ԯ�v2�&Ûqw����Re���U[��C�IJ�a�����:[Sμ���yu�S�t��ŕ�e�̾�,@Ւ7d;-�B�uM�8�5��2ӟ:Ԑ��K�u�?m��f��0JM0d͚8������q�U�a��4�8�Uvc;�vFEUr[��3j���KH�Y�+�o��}�8vo ���ܭ�x�Q!�b!�����]�u����Ao[ښ��BL��5��܌-U%�ج���������3d��n�0�UV�.鷗1���Ttv�U\�������K2���D���$����Y[���t갢��M1S��^_($���
)j�+�ʤ����:�G�jD�;Un=T0lwԳ+c����փ��.͆uUQ�ڏBmG}�3�W.��)���]��ٽ/cù����{��Yn��n��7o`햎b��Վ��d#I&���D��q�I�9�x�Ϛ�yy���zh#t7NS�u��l�Fb�
��oE�u�:�j�\o��EW�yyǵIwd�I�n�'7��v]�U1m��2U�2VmdU^s�����dշ��诬μ�u�B���ܵ��WQbS*����^�ʨ���F��h��,4Z����.�Qd�١{8��Ӫ�Gno+
��sm��\~�bhv4���c#z7�::��&;\�mպ����0�9l��v��e�M9w�c�se��&gi��uM�C��c3�b�u©
�EF9o]c{��;�?a#s̼�%n��.��;8QɎ�z����7�Eۮ��8k6�yE�gE�wyN�­ᰲX�u/rz��oN�I�ݵ������M;�P+�sM����6�LX����;EV-�:�AT��yΛ�gY�TqGVڬ	�Ԡ|��=��Ŭ����6*s�#3m�X]k�룋o
�M�*BE�I˥�J�
�z�ᙋ/KS�"R���6�s��I�'=p���+�ҷ��T6$73o�+;G��{.왆�]�Ү��N�m�5T87S[wF���Q����a\�T)�Ղ����ћ9��coP�@��n�D7���W�L�R����;�����ߺ��sl+R����Nd���Ɩ�ф�_���O֒Ub�g%� Wp����u��� 3���#/CY�ҫW}r��u��-����B.|̛p�����s'␳AJ��[��l���͈2fl�|T��^�g޸^�[&n��Gj�cy>����KH_hP��*���H�{���9��^����)�!�����3�c�R���#���Trp�r�|�V?�����n�h�٧ՙ����A�k�W���@�1��˼Χ�	��/|�ع�ԭr|N|�s"y3�n��6���nd6�xp�I�:��uZf�:q�UP��X��Nf���Zy+���eR���"�͢���պ��($�2�*���+ji�V�Ɉ�m����g�ڱ�u����\U��s���B��/��V�d{w��|=u� ���i؍]���N���z4��J!�r���6���U���u�2ε�F��O:���Q���vj��ꨣ'�����B\�w4n�^��e��O���S#��i3�n�%*b��!�b��9n����u��(�M3&>hw/��-Ӫ���Y�2	�������,#���U��y$� �I�q�y1X�����~�����^#l���莻����3;,��l^:5���>ޙ-�^<��o2)�v�*�3�^����P�%��n)��v*��w*�/���ߣ����,M�`n�����%8D�2Qݪ�JSW=Ǳ�w3�e�nŌ�������/A����"Xz��U�*������f��1�0=j��7s*�k?��[74V���٬5 n�$���	S����kϻ��[�7�Sfž��1|�7�`�W!t�x���]κ6Yٔs���J��ᅋl[��9����2�Kɹӆ?X��%�F�]n#o.c@��`�/.gu+㽣jĤDP���(��z�|���1�Թ�C����x{*3�VȬ�P�C �{]X�9\�p��r��GR�W'W���ۺ�_gh��>d�=]���ι�;�XZJ%���Gn�\�16���e^-��|�~]���B��j�}6�vV���2e:�t*�^uev�PL�A5�;��������y�:΄��T�v\3
�UX��*lcn��ϴP�
��3�XhG2�+Y����i�!��x�Ъ���-�$ON���ͫǇuŷ/�֬��w��U)��X���v�L���F�ik��!.ۇi˜���E�u(I���'rKW
���Pz7%�[�=WB6�R�Cy��M�u��	�^̀��ˬ�p�kY<~�H0o6���G_(�ԫ+�uo7r�d�ki��EUXΕ���*
�W�9�Ãz*�7Te̒��D{q,S3+vR o&Va/z�Uk�+���WԮ�9?����iZ��A�k���|�Z˭�\�6����X�eC��ʢOC�]g9>\K���S������\�5�{o^+���~�J��y,K_����(2�W�ȕ���k�;\
:g�Mغ����*�n�.��&� n��n|�Y��7�y�����nѸSl��U�9kn��7Ɗ�kz���s%i:27\h��r*����X���A�K�~�$PJc�cV��X�����i�m��:���%]NL�80�*[���I2<��lz����{Y��y����0�{nh;׬�(b�l���*q��ͺ1Z��!T���y�z��w�`���	Q���+�qU��}x���J��C�Jm�N꼊�%Q+��z���L��L��|��c���"^S���*����f�r!�o��ݵ��s���Z{�<I7�h=����FgM�ZwS�ee�!\v��S,V�n��]N��$��%�	O�ӊx��:!���GvN�񗼹Z�����;�%R(�u�3U�X�ļ�K��72m���|m=l3��b���/�*^Y�Տ���珯wj�w9k��jM�ڶs*u���^��V�\�齒�fsCM�#y�M���H�ƹ��X�����ܼz{�2rރ(�Ay��	�1�D�⻹�0+O��Mk��.]oQ�V��.DnZ��-?���e	Y�Y�I�0��su෥V�<5
�:�N/�w���Yh]�ŤxR��T#D��V��0��j]�b����8Q�f�*Go^J�-��\��l�y�ljHY���]w֖;'�U��.9�3ol�ޛ��Vʹ�|�fީuH�������a�����ʃ����]DJR�3.�����Vg��%�}�.<ŹW���%���m��cj�i��ͯ�Y9�Dl�wfg�g2�,�ӵq
�T����O�ùm�&.*i��������Jy����boVh��~�B�{�҃���j��;Gm�����F����r�'{��V�Q��uW�M���[�,�vx���t��N`�U�m=��`�Bh˛%
���F��sP��t�iȥ�]�b��E��92���w��B�q�ӯ���<�������Խ���؟�4��� �[b{�F�f*�)��;�w���}ۓ����6�nq_Kܻ8�������	<��jY��k�*��#�由�e6d��>��2O�N�O03QZ�0E����;��{ZW�{�^d�ThMɍ�J_f�׵Kyҵ��ˍ*�o��o�n7&9Ѻ5Z���8ݪ�}�+���jx�1y��BB��Nj���5�K��P���^���Ʊ�y����Onr��Vs�NxʃCd��fx�	��s7si�&]��ݜ�x+آ�V:֖w`�]]�3�kl5�W)˰]�mvH������`����-p�;9��ؘ˴���lXe��hI��l�0N�㓧	�8�)��-4Lt�!O.&���>�֎�?���%Ÿ��  ����g�F�s��h��n��l����F�m�{Y���i���k��x��#�'i�,-6̨ˍ�(��Y��Lv�iA{<���͜q�"�8�SLg(�3�et7Rh��/;�n^�>"y����\&���Z�[ԫ�@����mwSk�n�h��㮮Ay�����u��[�kE4�Ch]��[4���-
�a�&ˬ�X�E��]�.����G&���2mZ6aP0�S�a�Q�XL��-���l���s�э#h�u��I��η��W��MӶ�랻ԁe����m���v;/.0B֭��"m\��3���	���e�M�N]K�۱k���s�n_ ey����k�*��,62�4D�-(� �Ѱ��7m��&����H��jG=\������^xd�ɋ	�4�V�Bn��`�8�uh����cB7Zf� ����!p;�9s��v�JP�+�\�[uH\�^�
�����d�7�1?��ښm��U���E�����$CWJ�Mjk17`ͭ%f2��Z�������=�t�Dg-��X�&ΒR�V��b�S�n���\�*���H�W�1�r�;�<�h�F������.Hx�x�y�S<�a���6����`�aNG�ݫh���8��BR&y��Q�R����+�q�8��5-�:�Z��F�K.���:��m�E:�g�c�Gqn^�%����<]�u
�cٝu-���pF֩ݠGz��!��C��o�Um�6�]��u0���M*���n��ۊ`$$��Op@���{z[
�z�g#Jb3k=��j����,8ʹ����9p�
v��p�
����]��[�n��!�Ve��[;vF��somb-X��E�]#�v2������Jg��6y;�nn��m�4�c[���ڜ��^�t6�X���͕�vH6�74Q����]�]�ŻGOB�`q�q���Ӯ���ɶ�t���.mm�x�\��&�=���]<�V�5�	1�[��9�R'aU�1��,4.�,ie�e�)�2k�\�V;a�+�ۭ���p���e*�����)i�g�k&�)�gv�xbՁ�[G58��[��'%���F<q\u�]�)�sr������@��^�؛@u�k[O=��o�{}��� �]�v��]]�Q����9;f�\d՗/N6�ꛃmq��N]�!� ��e�]�$�v ��QK1Ys�p:SL�uQ����k�Y�c�y��4s����h�����:ɪ4F-g�7<tN��k����K��+��v�z��I�4�W/��ە��-�mX�^���kv�Kk�Ab��:�.�4���T]���T�pz�/n[[��2<2��7k�WV���u`�h�]Z�!�F�B^�҇��i�Cc�1�Ŋ�81����v{�#����Q���Z�l�qG<���ݮ;�!��l�%1�®��,����9�T��!��p�:7u��:n�wv���'��z���W-�Y����$a�f�Vb�!z��1ZF2���f���sMΡ��Gh.+��5���h1[���6�Y�啴BjF��l��������
,*�~��&O��rr�s��l!�]�  �2n!nj��6Sk5q7N�Հ��K�'����ʅ���dV��0њc	)�Ev����ƹ�m����4Dye����BX�m��kU��BiۦݮR�dø�y�&	�l���ѸՍl`����a�F���Q�RN��r(�$6J���hve�	2m�b��0�c<�a�F�s�kh�$Y��3b޳��JC�����t!�J����Z׳��n��hܺ�vb�t:�vn������Z6jٙ�̂�8����y�Y���dsֶ�ڂ����qd]t�a��ۨ�y��eFhCn,��Rd�����3e�]���Z+f��@�5��$gn�ȝ�Y��F@@Ln1)��z�;�`�u�c!U�G9�Er�b��ۘ��h��x�$���wY��1��0��H�b�c6W��>��yyN�Gnj� 1l�ѭ�̾X�f�����G����<B��5��Zuٳ�5�:��P��q�t�-��rUq�G����Gh[L6'2��m�k�`���K.�,�nGkdE�.��u���5�|���]�O��	��vt�As��_�󷫰N�ۭ��y�]�;)0�<�v��qvMqg�䌚xŰ�u�ں�4Ӌw";\h�m�2��͍Uu��Y��mgI�kҽ`;n�Z�|Sxqm�KE轭���5.�m��Ԣ�Z03�q���U˽q\�u=�9̬;���P4t�:b׳UuZlrMEc�+��ܺ����̾5�%,�+�Q���n�T���ݕ;��:ͼq�M��ǧ�
#<8g�ø�u�����+pʨZch8���h\uݴy��5���f��h˳b �]#�ƭ۱��t�Y�m��-q�\��p���� v���=����@�L�J��m��uƹhx�]-��c����h�&[e��u�����w`�AQ'��qT5%qp����G�ű���v�
����6	l�e#���t׍�;����K�1,����ؖ�q	�� ����g��� s˞�M��kZmĀSH�"�5���9�Q�b�V�ڹ�B9n��]X/s�]�]���lF��,Z%�hٺ`m�6d�E]j�e8��[^v�e��;�/WZ��0��L���:�X�J�A��,Wn{W.���[�Qd�v�^����lh���� ^sD��wL�ge���4YJȽ�plJsYKF�=�\�����}��ێ��l�U�U��T��ɣ���3�e�^+s6ȻYWX��a�lƞ�b�"�f(NS�<V���Qܤj�y՘�R�iCm&�yc��;a���h�0�ڞܵ<�N�;�-�-�[4%`G0��hC�]��%gq�zt�:(cZ��`b�s�[,D6�sr�p��ay&��MQ�]8�F6;4h;,�o-���$�9��7�g��=t�-�(�{l66���мZ9:��#�}�^�K"#)�"�F])��'�=6x��:<u�Ϯ�ԗh��\`��{]4�BP�c�ݲ�^�j�������-C۫��F��z虩ի�]�N��h�\ 
dFG�'���=N��Gl\�
��Dr�%�H�t��)��Y��0�x-��㞢K�R�2<��ƻ��q���v�F��&��nF��5ۋ�r>C%%�]i\�k�Ƅn��v7/.�u���Nzj�uqԙ�萃���a��qۮvw]5�D>7N	z-�E��� :�.M#���86��Ѱk��8rLtcpr��o.٪�-!m\B02glˊ�c5��&�����ř|g�q�8�\ �:���gq�f`Yp�g��Fe�-XlkZ�(M0��M�2d0: u��r�fǮ�˼/[�ٳNm�L�R1��&���J��.�iL���y��sfV63)��Z�^ִd[���{q�:�R�N�t3�[�b�I�g����θ� �]*u%m�G̸�F2-�n���:�z�v-�	f��In�����dʐ�9��o5�ŀ��-k-��=�نޞp�ݛcU=`B�4֨veI[l&�f�M�5���9���ʫۥ��F M@a3��մt�d7"֭N�'v^��Lc�nn��A�UȅZ8�i v{�sD7iw<sɰ�ٕct����t[,J�V���!��,���n�嚢�;4k�z��B��
�]d �Î�'�M�{t�q֪�ettO�cp�uWa�]��qO��T:z|[����utꅝz�ɬ�n�Mt����`�ؔ�׹N7��с��6镂ZjF�i�ڱ�2���c$l����9���s���e�GKF+���������]�����δ���\py�h�&t=y�tv�u��z���^���c��/
���W!����e��^]
�ۙJ��[�C�1��'3/�/5ܚ��^]� ���s�덀* �B�EF�Z���ʧn:���lL-�8�ȼ�A݃�x���ԙ����
J˷,�.��Q����y*�lgp�ַI*�\��k|(�&k+6|�am��Γ7L�5����5+gu��h2Ж7.�.zՄhVCMXW&,��.�A���m���cl��0V5��1B2���Vl�S�۳�^7Bۉܘ9�a�5�ڌ�qx��&�*P�{v�����ola��0��[���v��n#bw�ku��}ZݵN;\��s�w�7_I��m[ȴ����-cZ�� Y[�{<S�3t]��[��='q��T�����}����}��9��}���ɨ�;��zL�Z�uu Z��i.5���u�۵���-Gn��}ۭJ	T�e&�#.#��P�!m�/	�S��GlpY۹X�e׮��<nR5lm����v���ec�l3n�ڂ'Y����.�ɸ4c�ij[U�om����ҵ�X(ż��C6닶����GBza�ܺ��k�ĭ�
��޶�!�^��'m����5]��m6����]�t�C][�imxH\Ⱡey剶�8��Ob�;Z���"'=�4nmS�v����j��F���jb�O�=�L.�`�sq�۞zE�ۋK�r���t�'p;�4�Ժaς�#o=v^6�]�YP"�-�=ه�AŎn��۝�]	خ9��rӇګ��'BKl�_�m�e����T��/r	^-Ȉ�p�Ҽ�鵗%���<�e�t�RG:�H����y�^n��5����9���Ge����"��m�h�G<�$�x�9'v��!�A���� �(�,F�ÝNtC��	Ӑ�'KI��I�������m�)��;4۴㍺kr��U�rr�%�p$n�R(�r�n��� 8"Fݹ&g:V�V�m�Iȉ&V�\�
,&h㣑'!-�A����X�E*A �� 1� ���#��$����^]��d���.l��[q ;��7g���ܯ<.��pFg9�Y5-�4�顖�v,���ì3�m��vp�,i�}k`��r/[�E��2�.qruׂ�֑�q�����x��VH���`� ��6�e�#�x.�GYwJ�f�<�-�m�GpuK���E�{v3>��Ń8�)e��.����{g;nr���œsU�7 v۬H��ۓ��z���m���3JH�s-&�eҏQ�yT$e�4�ƹJ�d�:VT�����D)�{M<j���kyI^D'm�3y�vE��sv�;�E�s�+ED��n]��An{[�.;C�]u���x�'��=��n79�o@b�m�8�uF�ۘ%��Z؝6-G�im»�vn9�8�',D�鈴�Ml��j�Ҡ��e���zu<��!�hݲCa�+�s˳N��KfmƢ�`[�mFD_(�I�Ql�&�;s��<y᨝T��Yh��]��A��M�1�;Ct�ƹއg�׮=u�[��ȸN:�A6��f%Bk)�e��ajfh�Va���,WnY��m Xͦ�.Vϴ탭��B$&ڦ�Bh�>�:֎W::��֦cۍ%�LVZ2�hۍ6U�ln�I��f:#�ȗxF��;�f�sƔ��8��+�6����Z�NR]�K8秶��#@������GmUKr�,� f��60�{f�Ѕ�1��mc,Z�[w�_ =vܕY�c.�狴�G4n�^����ύ�<ۣ�=�8���������D<��G���*�3[��掟mЮ� s��Pu��:"K.،/SK����	v�:��뛺��ۢmc,rշ��;u#�;\[qn����*T�rڍ˒��j�[
����;��5�h���"��`�A�)�-�[Fxiwc���:���Pȑ����k �!���9��4�e�&����6�$��5� Kn�ѕq���7n�:�W��Q-�ZHK,KX�`EhU
%`P������kȈym��
U[e�i͂��YA�8��VR���E���+j��Z6����y�/Y`J$�YYjj�$�Ԍ,	e(հiB�#X2�!D���DR�QH���?��6�Kc�c�j���6.;5�hz{d.��4��"-�KnҔdڿ=�}�wߧ{�(}"��_`������|��~���-Z�߯�5}$�Ⱦa�%Pr�f!"]�s�jk�b�U�c���n��5Y��\߽�{�ޡ"�}��Cس�6w����:�k>�9*D$�>���Ƶ^��k��:�6��y�E�����|}Y��l��+�3�d�@$�$�.%~�:�ƨ
�[�7{cS]�)u]�j�f������b������;�fѱ��t�n��͡X閩����z˕et��eШM�����C5H��R�}�d�6>�|3ee��gSO�[Bu�����������E�]v���^��J�U���I4D�
��IӁ��!SM�[���+y3����I�K;J��U���'��tU���ǆ�w�v ;��uvm��gJ��;���w��9	^Y������[_{�	%}"I3��g�X��y�zN�����\mzj�5I(	�!*�&��OʜP�@n�j���hy��xڵfg�I]6���a��RJ�	�ٽ�ճ�}~�renm�d�J�L��9 7��}$��KYՓmRh��V�"�.s�|��.���m�J��=M�a����m�M2T���|�I�b��
�s��{e<�f(n��f�2/�}x�m	�$�r�%�T����?���|��84g������ͩ{���qz�/W����%%�α�׹�|ݖQxZ�V���W��&<�d���রU��j.�l�䪽�)��x��\I=Yg{v;/��i��~���]:�D�H��ren�ۺ�hPV;�h��9��}�	]������uL�/*��t�Xz{T7����n��6T�	&[>��p�Jz�g�)/=�7;9�
��R/���]*v�ۺ0R�n7n���9�rX
��J�6�[Vh{`B�G�V�$U��Q���������/z����E1Ʈ�����B�}�Cz�����}��]��8��s���.��x���u<��u�/|&�����z�H��Vֺ�6��CzW�)MH�����]�\�-{����5gg3� 䯤_H�����7C"w��؆�s��cg�H�c�xN�X��Ҭ�<>t߷='���۞��j�Ʋ���˔��iZv*�3ʇ�����^�*�������R��:޳�i�l�X:��%f-�̗�]�BE�IRx[�/u�ؾ^��C�=���vc�I{�5}$�a/+[+Z���+F<����c6�]��M�2�E��9nخ_K��]<'Vh�f�V�C^�@tR/������t.��:vs>���[hF����|$[���c8���
��n�����VgL��|6r�Cv_u�}l�������I+��I�2y�M��b9�𞞓��vb�	x	���$��BD�wk����%}��]�0f>+D�7������� ����]�����o����t�n���}M@׌�"��᳐�%�$��wț�W��S�P���w�GV�S�Z��Tj=l5��u-D�I��m[�m��V	�N ���[2`�5F�#��Y���ռ%:�IZ|�Ua����W"#�M,��-�����3��q�W4тѧ9�n�d$;���5s���ŷ2px�r���}�Ӓ�x s�;��;]�ܠ�<]zm[n7,�$a��W v�v��t�=\�FBtLtg�nu�X�����.�W!w.x5�a˼�v�J�^\s���S�۱GHVk�Y�����a`�n��D6ح��l&�����--���/Bmٻ۪X'1u.����F)�B�(�.��~c�a�����R $@-�߻�zf{���μ}�o�57�	� $���q���̡΀{��zM=Fc�I$t��d�&]�\������n�"�IC�4�2��=nht�z̧�}��d���Ӥ�$��P/pgT��k�H����;s:c�v����S�s1E9e�oP�����>ݭܾ�����#.���Z�f������ի$�"�{y����ZF���B3v�B��5b���+��r�T6�31a4�H]!S��
[+��ɚ����GO�O{�nԮ�\��G_
������5P߷�G�I(H��/�3^C��MP�|,:���c��٫L9��3�r��WֽS��a�T�ΞǊѳ��J��{-4���&
oYN����R�{�;�37������nm�&1U&����.�H��<�{s*�w,e�2_�oZ��������(H��H�����=��M}���7V�:��SO�����|o�VUy7���u�����R!$�(Y�v/���:�굑�鹏��ɻ~�M_f�$�'����z��ZdP�-]�T[��+s��\�+��ݫ��X[�2�%V!�h՛+�w���_n�ۺ��I4��gK,G���vg���m��NbD$�>�X���[y�pz�ͯ�op�S)�������(n�ډln�׼}�d_I$bF���B�'=B��`��oUpM��7}�FַG�k��*�h��̘�"�.�������`͏M�}��ѷj�u�W�v�;�nT6ܬAVj}�;�d�9't���}5|3P�W�D&���Y�2�JĻ;핝CwW�)&����e��'��s�A�3%���}:����/��k�SL��z�t᫆׎J��v׾������4�;g�B�<����:�֭�6==�ݹ���b�cqU��
���7(c�v��+�y����Vn�%�l{v^��n�N��k��I+�w�U@�y)}|2jt�M�ȳ��6L����$�'���>��L����H��g��C^�v�7M��%q�O����}�>@N���Jj́�k�:�P�^��oG=q��p�@ܼ=�����i�����)��u�ۢo=�e�/\F��}8UY5Q��m��HW��a��]㵵x���fm}�r���7kvt9���u=_:M�u5gO�9���d���l'�d���e$z���-�sʑ�\�u�p�]k��.+��4�G\�-�h���W�`�<���#H��{��F��S�g�5��7�d�רu�CwPݯ��t�r����W�;��Nw�	���͛�-��>����OT�]��ϐ�����D�N�u:��q��Ez���=R���ݜ߾�C$��$��}Y�gֳ��_<ktc���v�=��:1���tAd�{�D$_I(H��䧕Pkb=�sG�o��=���k�M@MRJu�>�|��1����V���BV�w7M�G�^���w(�ݵ�ˋ����w!t0#���c������km&��޵�۲�f��F�*"ҵUJ�]���Og�{Wm`ݺ���\u�[\�gl�\��ő����)۟B[���IԸ����v�s�tNէ��=�&Ơ�s�;������'�m�na�:�����fLg�0��S��m�&�b;��틋*d!�u�;4[[q��ݛAƵ�g��������c-��jK5�.�õ��&�3�)����eԺa��
���_�K��$u5�4a�4tŶ��3ìm��h�.ٮ�Z�����y��Ͽ^�b�D$�5W���]g�ݜ߾�9V�/��� �T�|qmo=Y�ʺWù�xh�:M�#};o�f�sFO�l��̺�9�����RIu�� �_����s{|#��嗻����I_I%�گ�OZ���{�{���樔�zm��A�7�7�{;�{���qws�5�E$��_�[���d�V���p+�`�u����������I�S��?![�Wj�ћA-	�X�F0:9���4�֭[k1��U����X�ؿ�}|���D�{�{<9�{�*�zka��'�F��g�u{Ҥ���Pm�TV�=B�v�ͳh��.���G
���y�R��ܫ%k�^y���E����9>�!����j\��9��<��;����>\��zm��@�oNo�^��J�{��?,����{^W���F$���+H�W�����}{����'I`I*D�to�no����z(����p����\s_����"�5颳s���}5	JI�Ѡ��1
�lT�շ�=�_�����7�z���_H2;�,�>�+�(�DRJ���ǝӄ�[��z�[��.�3aJ��\���u����~�}�$`H�wxn�:Op�����ILmu]��{,M>�qv�%H��ݧ�K�Gք���k��ݐK�|�d�����$��Jv��S����_I%�����2���9yN��f���
CZI]1c�V�������[P������`��*��y\����Ʋw9��;�:�n�!$������]��}����UE��;1�	�*��f�u��Yb����wj����Y}X�҉�L7g����Y92�\��b��]b�M<lض�l<{5׭�V5��Pl��Em���t�l��%b��ض+(�����r3��K�o�[�ɵu��p'*f�.��8Pp�J�s�UL�|v޷\���HE�ʮ��Ms�sf�|�P�j��5&!sU\hf���i�ߪ(S�h.GD�tu�o�������'�X�l���W�}]o,ۧф��n4�Ҿʇ�==L����{x2��e5��w�o�p�	�3/^=�X��v�0�V[���({�8��n�&�BX]h�8U˄h�{5����1֋��ˈ�����A��3t?%���YλoWuŘJ��4��W��v4�J�j�Z0�q�}{s�}�w�'s͜-�I%��Ѻ�H��	��z��=�ʹ_9oV-u�,�D����q&h�tʧ�.Qn�FG���0��룉{��;�7���Qۈ8(��Z5�%VE�y�7qmM���c�J��̣�WՋ�M�'�"��m�m�M�<ҳ{K4
�@���z!XN�͘��gU���|�j�6{�Y�:��>��h·(T��/xo���uȜ#.:���K��:5Θ���1W��
�5�N���F'��B�]>�;A��QU���e�ή "A�A QL�RAݓ�p&�����md��H'��(�,�Ȝ�m;m2�(���P"P��NQ��$��C,E��$%-�6�kq;���gpt�Q)�bqgE'6�:#�����K��Y�am�38�-�2�t\�P����k��Ck.γ��)�E�i4�;��.�I#;��(�'H���*��ZͲ����M�@Qqdtt��:��VM��.ěL��Gf��F�Gi���,�Ӵ�F�ek,�Q�vCm�e����;#��b�F"��������w����I{ӛ���H�_I+�E~�fi#2��[��G:p<١3zR�~���]����N��"J�7y�BS��Q,�܃��g����'�͙Vډ}]���d]XA]Ʒ3��9-�j�W�P��b�ـ���3�����6Tߝ���n�)rk�7�ѓ�;[��]�a��A�nخ��$RJ�D46�.�G�{�_c'q=�P���^�� ���!���/
�[�P�$r $�^�.u��LZ�vxl������5'���%"���vgd�v&��u�)��瑟S�߻�逳8c��w���)]j��W��(��1煊Y�.�˜����*EY}�f����^ј[�qx8~�¼�g��I!+�g﷔���H���~�p������w	܂��⓽{�{>ٻ`n���qV�WWʗ�p7i,S�3�l�]1���%��V-Rb���F�Hա�۔3��n�ۧ\�p�y��V���5�y����N�R�N���W�D��A����񱒾�W)r7�o�G�#���n�K#��r�ʨwr�z�ݡ$����f*i<6Օ�~8�A�|Uu�nx?m|' $BIBD��-Vы*����v�gvp����+d��=\�'눧:�{.{�
fn�rE����! ��ۂ�k��>�^�\�W<��[��2T��(��7�UxZ����{DsoR��]O�����u��K�w��[/��Aͧ�2K�vU��v_��}�;݉3�r�l����}Hsv��J���:N��w�=�����-�2�ËC*eY�cڂ��J�x-��1a���:k ����U���SSGWY���6�(mxn��L����ǎJ<��tTHk������eԮ��^`��u��b�P������9]�3���Ȕ����[f��ה��E^�-af��Ф�=��>m��,Ӟp�V��sL��
Y�����~���"7lP 6�Aͻ��p�\�j��ݰo=s�3��D��~V�SO���# w{��g�|�m�L���Q��~���ܖ��_H�#�b�-�w�;��y�to��*ww;{��I0*�N�+�5�{�Ջ�(}"�}$���s�>�����N+�;ZS�o=Z��$	�P߫ ��K��t_P��/�h�wb�x�ҋ��s�ғ�Gu�d��w-c����|$C�%|$�]ZTw�~��g�4z?g�����a�9n���$~�Т�u^v��W����n3�]��Y��Ƿ:�uΠcd-i�H����R�dP�7���ۻc��Mu͜2.y�mg W��\�%��n|'b���}�P�|���6�q�K���5w�P�~p�'��������6j��:u��2�O�V{(�W�<�M9���Z�y�)I�f%���ԋ-��wY�9������ױ7@��߳���c�N���w��_l��Y��Z9�:{����O��Qhk���E=�+;s��Ν��^����$��E��*�ʷ�ݔ9�ۺ�)sga��v�����
�7i�5��m�⏭��b�P�$�`{��c�}ռ�G�*��S���w�����)�Oe��Ke������#����0�㵬nf�sMx��Ex2���_%f���/���_}2/�k�U�������۹ӹ�k�J����xךZ}�x���4�E"JQ_mvR�!]�l�]];�Z��%#^�j�ww����wr�w�}�_H���y�Oi�*Uu[��!�0H��]�u��oՌ�BLL�5����e}W&�	Eob����e���gծ���[1�ݭX�g����yT���F����]�G��Br�$��_ڼ��������k�]ݜ��v�w�w;xNH#I!��R��m}�BD$�>!'�ct��e[�^���+����Wv��_nJ�}!Y鞹o+���/ei{���. �cu�t[�=kH�I��m�c��l��T�쯺Vhw;��n�tN���~��}r�+����.�>�T�H�����H=(}��t�=��Z���X��/�T�.��,��%s��|m|$BE��f[}��Xogo��vν�]�OիrH��$�uE,���Ǖ��=�Oz�ݣ�}�n#uϥ:��}��t��~�����]٧x��}{2c���և���o���aTr`��\N�F�[����b��.Y�)i�<�ړ���|����OHĒF$�����ƻY��v�%O�f�9����X���7@n��vz����G�N�U�ʐ���e!����Q3���j�[4re�tr��7�	���|�=��v>���^9�T��(��p�~R�Ք�/������FA�Ȩ~�W{4ɜ�Q����6���N����ܔ7�8�_"؂v�_��A%� �����:�D<L���{�o1���O�>�Ư&��G�8~��R!��_L��!��V�"�}�o����k���;
�㷗h/w�m�pc*U�m����3(WǺ��A�Ȩd��B��J����*q���
���w%�:�D��ݤ#u}زy�l��pMv�?Yŗ�*�fU�N:�4N�sMiҍu��,4�J���}q�\e�u�]�w�/S[��G/�h�~4�ո$6m�IelS�}���"����]�ZfU�f��m�;c��t�]����g]�H�pY;.����g/I`ӻ<K��P���yɶ"x�5�nXV�q6�d�|���f���w8�K
��o��nI�-k�0�輧\v��E��m��L��CPTMl^$#�X��f�k��ɫgu����q���K��é�ax#b4m@���	X��X^qK������H�Y���.���WA��[:�&���.���r���v�Y����o*�{r�s�\C����^����W�m�E�(�:�o|���w.堂1У�L����"�L�q(��������q���u��8����az�:@�����ԡ<П!�_v ��@d��A�A2$��h�>�7y�hPx�%�g��1]�!9��l���/�;��F�N�uٝ��������_2: �;�!�һ���X���s�O���"8�����2g�����2����?#ǉb!�Yq�+�x�c^a����!��I�O@�lv��l𦾸��j�W�IB��	NG35ec/�}` 9��kU���نց��խv�q��rTl��9гUM���=��__X��}� �dG=��s�L�{�W}�G��G�Qoh�"��mx��� F�dTG��b��M�#��^#_ax=X��oH��a3��)��יO�7,Va@�fQ"���1;�Q�R�R�t=��7�u�ow��5�/�u��@�j|'6����_ox��e���^��{ğ ����a��T���k��v��_k_i�!!_�!�jFקW�%�z+zv��9|�����ڸ�����.�9�.<���[�/�Qg��g!_~2*Y;;��/}5Uܔ7��_ A��bF�o�b��_	��ED+�"FX���5j�+���]
�rn���%gM�l����y}ShQ�
 ��V�u������>{�`��s���3�dN�k���N5�,�C���ڳ��QB�	�����e����A|wiwWɥ��)��z�x+����9<���}�c_"5���A�AA�QckFR�z�����T��ދԼy�j�䡾��:�_���Ƞ0{�S��w:�D%}@�*�2W���z�|�N�d�-y���;#�jad�`���R�Z�%��̯D/����n�xpMu��������s������Y��ί�I�f(b����� =G��ν��۞�7C��_R#]�
��"�$��z*��V�/W��_s�wW��<�pS�K�z�x+��k�6���͘�_�ͪ���(�AED%
 ȅ��Qػ���R���ܽ^���J�J��s�ᮇ�ݤA���;�x_�U�.��,�_�nҬ{sv�X�b�����sp�B�]eB�A�Q�E���X�}���ھ@���}���Ͽvt���$��Ή�<D|ʾORǮ^\7�r!_L���A�|�w�pD1��_w��5��s���^�ճ�] ���|���؁8�c��
ϐ�(�B�?ʀ"E�2�E�Pˡ_O��ڻ���:WrPܡ���������DnЗ�68���A�u|���gӳ���;���z�T8@3�|DZ��[�\`�m���q�%�5��G�s���Lw�C[M]��\�S�21�%Wvkk���NW���O;�SY�������$��͙����|D�@��AJd^���͙��	��yW�r���l���l�W�}�HvW�G�|d���U꽵Ws��uVMɍ�����GZ��>�mur8�S��l��T��`�fR@���K�ɝ���9�t�䡹�����{���\��f~���գ�\9���9V���}��S���� ����8s��k�Y�M�=D�A3�u��h ��JGZ[���[ڴ��b��,D�,��`�9r���g��cɄ�5��4u�w9ג��^�K����W�IB�2!D!��b����� ��A҂��U���%~��|�]�C�� N��3�xߕe���;mP ���"|A���������Y�_�'�-�����ˬ�nn�<
����ڴy�\y�-�(��i��w�e퍻�񌬷{�]�U��y�� �8m��}���+\{��g3f\���`��	�x��f�7q�5�0�bV�Ub�K(�m�+���i^µͧ;�Y����-ctI��k�B*#��h-B�ڐ]�uU�V�Z츟e�ڡJXSֲ��=��!�����d�F�ŋ�����M�O(�Nx������H�������!$��.��y���()/�m�nsc%�l�����貜���aC I�p1Ch����e)(BF�4n�`��"1�>�]ٹԋ�6Ŧ���"����Χ���W�9G�6�,ګ򗗋:N�
2��q���x�fWm�ɷJ�9�b��f���u���c�oKX%��@���"[̦�g=c���ͣYJ��q�������76��ͭgA��Ԓ-稼p�;�Q��y���jXW�R��w8C�9�xr�����J�i�䛪m��ϼ5k�	��P�#��E?g�ڮω�g��$����@�"�L�X�'hlַ�M|m�伭SNd��qR�Oӭ���a�#��;���vo���������ySO�/�zl�!)�O[D-���n�b�ۺ}۝�,ᒃ8��$�۪v�������ƫ�Y�˓�EMs!���Pe.��R+��Z<l-��7�*�$M�2k�9��`���P[�uc���=B������.��b�J�_*��UJY�m���9jb��鄅�C��6n�UWPJ2��z���!��7����J���H^w�H���e:�^hjy`�2��m�(�^t��� �>!$
$��?�f�陚�ce��[���cmsm��; ��5�E����؈��fvu�7kl�����M���mY)I�,�2�6��%�Gv���سm��kDCX���.-3���n�36�l�������k�#�V��3,�ͷGm���K)�mn�R�F\]�,�����N&��΋����v�e�u�Rی��Ⲋ¶�ɳ��kXqխ��3�v�+2���;.ce�Ii�V�gv�v-�ᖛ�tT�e�Y�F��%�ݶ�:I���6�4�;�:ʹڱ�,�::���7���|���Ĳ=�"�u�p�&JEH�n����Z��!<B���!�.er�@5�aN���a2<f���8L�Mlk�J9ꌴr3W̓lLʦTk�0+K�^��O(C<�g��L�#4��l�]��B3q-�9��Td�QN{;�W]V���S.AI�RP�T���֗]�ۊꖡ��<4����n�X�lI������`�e��p�s!�+�i��Ѹ��E��ygf��U�}n���Z�=�:�9�-��< �^���m�ݧ]��E�y�b�9J����=[�9���!�A�'�V8���9��i{n���'<s2n,�'��1��F���+�i<��`u�{>��lθ���#v��,����&bka�=�Җ�S4�<�u�&7Y��.�"D�j�,R�8��D�OW���K���K�1>�N-v���kX,Of�����u�o<�u���b9pC֮��ݻu��@yI��T熩�v�d�+�1�:�k)P:�h��v=�����W{�Pu��۶{c��wV8�XL��|7ګZ��Kh�j�y���Z��dtEh��w*�jL�n�d�+��<- �����=�=���ł�v��\�Փ��5�MP�f8��܇\s��F�6�6�B)��#�Mj�R\2]u�U���AX^�\K@� ��@ssY+�,P�7\i]�t��n��݈���b5�̇;.°%{c&�V�)�M-ee`�M-,y�6��-І�5+�6�kc�qՑm;:����e��u�ym툮LR��\R����7L񗱜t��<���.܁!Y�'9��]f+�d�"ᱻ�l5�FY��R�E����żrYZٗ1.v.�"� ��a�54h��l�2�+ j�L�������;=y:ȧ�.���O'�Z6M��=���.X�g�a(�V9�-���Bf����t�j�����7jN�a�]V@�f���{t��͛�`{m�B�\F�*ݍ�1F�������s{�T�]mm&I�qn�Xڕ�-��qb��c�xat�F�0��%M��-��01���̤�;�8��l;�j���^���.ֆō��9ャ���{%��ûzM�ŹN8#M��ݔ@*u;����=�lh�B�67�4�8�m{;�1�$���Ѫ����##��=`ު�5�ex�e0�v2�r�L��;�w����gA�`m�*!���N��p��V�=u�+ĚN�*�ѵV+$;�P?��9��D�/�,�w8K��3�s2u$���׍7�Z��˗�\��X�\g9Wl ��o>n����n�o��Q_�7�D��{���D���m�}�Tz�c`���!�ݤA���#u
KR�w��2��%�5֠���px�A��whPD(��}"�U�R���}_B��m"��]��ݵ/zO9�m�
T;㎗�#:�=V�=��<�_f�@ȅ�TD�Q�G�s}�7��%5@+~�������U:�B?}@�9}@��P2* �+�aD��=C= %^<1�˔���m�4��ǳt!.��-�]4h��GX�Ze�ݔ���n��ub/N����&�f��"W_=����(Q���AEDI@W�/���h����v�^o~�������[3��m�3s.o`�s�`�L1�s�e�u�5<��ͻ��[uѬ9��D���}��|���?*��r��]�������s/�WC��_/���#w���Xs��?.��u
�y}"ȅ|A2'�cV�?a㹗�+]���3��:�B?P?�� �&��&?I_W�I_Pͱ[�5�G2N�BcW��|;��!�^��*��y3&�f��?w���-�<�Pӑ
����%W�/�d�@Ƚ������K�����s}'l��&;��,U������?��D|	 �3���$ݠ0� ��H)�����>�8y��v�������v���$�>�;�&i�ηZ�nGq6�2h�s̼)�U����k:��P���ϨH)�sۆ$�)��v�c) �ݠ-���:}�����<�~��}�֐Xo�G
C;�?{��U{�ͺ�3�>��H.F$�m����L9څ��JH(Sܵ ��
n�`�$Je0ݨZ%$������~���I<��
AhC�PĂ�7�}���������7��x���Y��I
R{�h`����i&!L۵�o<����g�<~ͯ}�A@��;@[H,=�G
B�T�ڐ\`RAM��0d��C��P��w-H,C�߽��l�?���i�T�$�[M����vF^���]��h��"�W����S	�;�묚�ֵ6���L�s�/��Z�g��o�� 3������_7��|�����$�(?�1 ��B�
A`wj������L�
Aiچ$ȁLڶ`�I��<����/�I�{��Ĕ�XW=�bAI�
`{ڶLI��ݠ-�\��߾��<�s�zߗ��i��A�8�RU@�j��
H(���;}�[��_��*P�0�h� �(-�r�-�9�\a9������σ��H)�C�T1 �Nߧ��~���Ϟo�n��ui ��JO~�-RAaS��bAH,ڴ��P<JM��_�<5��w�]��`�fB�.���K�Vi��S���Qn�ΎF3F4e��Aa�T- �4*�s�i�$�hH,���n�-"JH(P�v� ����<����\߻��;�w�bAK��1 �{�����>�����B�>�I���i��$ݠ3(��ZݨbAL@��[22RAB������) �w~�;J͎�d���|	` Q��L��H)>��_<��{|�?��]r��ZAa���q �(*�o�i�$���1 �#%0ݨZ{������o���q ��aܬH) ��A��Y(e0�j��RA`V��A`cI7hH)���YD�Yy�T��=�7s?RsϞo����<`VU���I
II����) ��ݸbAI�Sv��RA@��ݠ-��i �ݠ�
B��7~?|4��U���S��`bAf�þ�-�) �@�v� ����}����\߻��y���
_�!���)�;P��R@��쇡�Q���c��f�`�)pdw�<}�[��˭�SS�2�H��U]��Y���v']c��F���C1��%�ؕ�e/ZB�q�Sr�e���|>I�
A`4�S��- �7�H)�07n�c%$)%&�i ���- ���ɼ��~����i����Ԃ��JO��-��Ͼ7�}�/��9��\��֐Xy�H)���ڐ\`RAJ9�
Aa�P�<�) �@�w-H,/�+�O*����4�ƌ3M�SR���F�S�+��kqd᫗ux�7P�6�S���1 �r�h��XmڐX4�Sv�̢
Aiچ$�[�Ϟ��_�c�;������Yv���I3�Ӗs���}�����
?}pĂ�)��ݬ��H)7h`cI��AĂ����ڐ\$~��˳̷�tH,�{څ��JH(S���}�~���ms~�������~H)~P|�$JL;�@Ĥ������4�Sv��ft�]9�ne�H)�yPĂ�)��.�c%$(II���) ��ۆ$��ݻY<I�)7h`}�o�립���2���w����s�ۮo|�mÉ �7۵ �����s�$`2Sڅ��) �7nԂ��$ݠȆ$O7w��|�������T-�) �+|�RH)Ϩ� ��ݨbAG}���Ͻϋ����{^���Yv����)>�����Xv�x��w~�|�����.�OFRA@������4�Xn�- �0���v��R�lH,�Ja�P�<���y��a���~򽯉� /���H��o�|������C�AK��$�ûP��I�S���F�
n�eRB�H)ӹ����^s��{�k��%:�;5ԙ��W'^�y��j�mi8ǥZ>�~Sm6�4���c�v6^X˟���].x]O;)�;�?������_���D^jwUz"V�O�7�{nY���8p�+\�3׻V\<��kOd�M-Gp�[I�db�vm���f:u��6]�7nD�4������F��<iP�s��68�;*�,&q:ɱB��R4�к-v���$��j��()�����n�0�%R�n����,o]Cɢ��ZD1,AƷ2�ԏ$6c�΂TԵ�cf�]?~�O�r�&�e���-E��V4.�LV޹�\��#�ֳ�ywM��]�0?m��􌔐P�����- ���i'��ݻR
A@�)7h`a�~��߽��g���w��R6��
Ci���<�v��
H)S�,H,�Ja��Z	) �Cܵ ��
n�b�Y*��@Ĥ���/Ϩ������|=��A`kI<��
AaͨZAL+~���}ϋ�����������R
AH)���JH,+��1 �ȅ07n�J�{��;��Y��A@�JN�i ����$����jAr0) ��$c%0ݨZ��
�ݢG�������շ�k?�xc��Oϛ�?$�(>C
AaݨZ	I�]�� �1����D�І�C
A`nݬ�
��^eg��k�y�I�<���8$��{pĂ�"��n�Le$��� ��<����/i��u��Q~�>q �(���]��$���^&���;���z�~d��P�0II
}ܵ ���$ݠ�1 �S)��B�
A`f�b�X�AM��v���_r���}�} �	��J�YA��^~�M�E�0+.�|2RAB�R}�hbJH,+��1 ������H(�Ct G�-��O���W߶Y��ʻ%U�í���խ���U���*L̓:98��S�8u!h��}�����H)j�w˵ ��������)��B�Ĕ�X�jAa_s߹���|߻����V��/��'�{Ν����+j�Ȕ�X��RH)�eRQچ$��ݻY�%$(II�@ZAH,9|�|c�����~��}w~����)�����DB�J�Zn�plK*(;��"O�g���4�m�~7z��;��k#�Jg����| �{��RϮ�Me$
JO��-��3��������>�y}��I���
B��s� �$�{`bAf2Sڅ������u�uzJH(~̵ ���$��$Je0��@Ĥ��ݻRH)�@a�AH-!�PĂ��i���[���^c�\+TrH� 0�ZD�� ��II�����'�pĂ�)��v����Rn������v�i!�/����3�����`s˵ ��$�ݰ1 �#%0�ꅡ�) �L7rԂ�%��n��k����w���C�AK�i ��W�>�sg�����5�.�~$|ƒ
y�i �!ݨbAL@����JH(RJM��Ȓ�
ݸbAI�Sv�d�����>�_���w��H(%'�-��w�O~�}���ǟ_ܺ�~���yA�q �(��ϮԂ��
V��Ă�d��C��P���Z�Xt����������RX�x3�]�@$�;lk�,]���nTI��U�::�ϝ=�����'�1 �mB�
A`a�f) �ݠ<2�)�9�H)�����^�\������
˵�2RAC�����;���E<�hx$���pĂ��~�Y0e$
JM���Aa�A��AH,۵ ���~�m����h�Y��L9ʅ��) �L9ܵ �����s���w����r��~H){A��Y(e0��-���b�R
AM����>�|���?o� �؇ܨbAL�0;��̌��P����hdII��H)0B��k&2�
	I�@[����[�o���\�������bg��0J���*�]�)�դ��ǬeM9��s@���X�#/%ߏ��*{$���;�X�قD�_;� �R�g��S�uzR��Q�͠�q �*�>�R��
T���Y�%0ݨZ$���ݻR
AH)�A��$M��W>���̮��;�@�JH,��RH)���AH-�H(��}_n׵�U�w��ߠx���Y��I
R}�i �������}���[��y���AI���jAH)7��
Aa�A�$�U@ݻR�
H)[�$dd��B�׼��O���=H(S�Z�XW������k���w������AK��H)��B�
A`gw1H) ��i �!�PĂ�����ߟ�(��Ϋ"�n�T������7-���޵n��gu��ɡ֍K�Bʳ�?07�ڐR
��{@Z��
>ۆ$��ݻY<����Sv������������_ܺ�~���͠�Ă�����{�Vm?��f���Ԃ�R
y�lH)�~�Z	) �7nԂ�R
n�x�$Je0ݨZAH,
�=�����]�{�RZH)�h2�)���i0��߫������w����k>) ����Ĕ�XW>�bAI��ݻY>�����|�� �p����24�X{�$���۵ �0) ��i�2Sڅ��) �L7rԂ�����~��v�~��~��"
_(>Ă�@�a�P�����A``�AM��
ApCv��0@����d����wǏS�}��r�"��@Z	) ��ypĂ�"��� ��� #������~���������~��RP9�ڐ\`RAGw����|3���i�-�]m�mӃ3�^���(S����Y$>맧f˻��x�y�hY۟�{����}c�^�y�<��ėUPۡ�&]���AEj��}����w�Ԃ��Jaߪ�	) �L;�����Sv��1 �S)��B�1) �+w1H,�
n�g�?��?�w�OH)�yPĂ�+����O}>*�������
˵�2RAB�R}�h`��
��H)1
`nݬ�I��ݠ-���z}����{�y���uTCS)a3��G�ҌԱ,r�r�[�ɨ�X2�\��'��t���gF�)��;v��Sݠ- ��C�%$(a���~�o߾�^~�s{���~H)|��Ăɞs���Ϲ��=�h	I�]�1H,i �;@fQ �!�PĂ��L۵��I
II�@Z$����������{ͅ��B��v����Iݠ-�������g�s��>�>����6��Ă�X��H.0) ������Xn�-=��<��}|~����W�� �>۵ ����A�C%2�s�@Ĥ��ݻR
AH)�@xeR� 7_#�H���4J��ӥߪ`� ��{��o�?0+.�}) �I)>���1%$s�$�!L۵�I ��lH,7h1Ă�~�j���wϹ���<��H) ��>�1 � �L7j�$���0��R�~����}�?s�����ߡ� ��A�C%�ʅ�bRA`W�W�ϭ��?���}Rƒ
~���(��ZC�bAL��ݻR
AH)�@Z	) �ݨZAH,۵�߯����]�������Ԃ@�3� G�6[}o�ٻ�_��9m�$�U@��jAq�I(���Y���n�-"JH,۵ �������}�ů��������b�W���L�,+9�}s���Ӻb�]enz�@�v����Ēk��^��i��DJI�.e�)��˜�|���! V��9e�9�fe]�9�kIo��%ѧ���<n�<v��Nzz+!c�.�Ҭk��՛:dG�w-며ۡ)0ǰE�`!cF�aik�l�9����]�0����ЖZc��gQu�ۜ>c�y�u̝3��>K7X��dI����f���P�#�lLp�]c��*�%�8ñ<�;�7e�0+I���kb
�K��X�����"�������3���q��,���n��{������Ve�m+�:�N��㦳��τ��� ��*�R��s����AM�&Q �!�PĂ�߽����O��g{����e�ϙ) ��=�w���S�P�RRAa��H)2D)��ݩ �`����0i �ݠ�Ă�����$��R�ÿi���甾���|� ��ʅ��JH,��$w��o�~�_?s�����o���R���!���L<څ�bRA`T��RAH)7h�Y��y��9o�R�g�H)��˦x�I
�)7hCRAaF��
LB�[tɌ���BRn��s���9�}�����y����9�������i�6�i!�U@�}t�\`RAJ���Y���n�-II
a��I�0�����$O+�'�{�{8���Z�) �(���H,H)��- �"�H)���߶�=����w����~`U]�AH(}R}�h`��յ�߾������'b����d�RA@�)>���4�Xn�c�!UP6�� �0) �n��Y��L7j�����}�}eU]���P�|�H,2���s���_߹���y���~H)~P�Y>L7�H)����H) ���Q �ݨZAK��=�߿{|V��~����k0��v���x�8�v�$S���E�<"�����[��.�X�n��JH(RJOy@Z$���pĂ�X[t��) �T�v��o�y�g~���~+�����i�6���AH{�+�/����ܼl���AH);�X�Y���wj�	) �L6�� ��aI7h1H,�2�n�- �	?��י�k���1����fYw=�l�OE�C�~�u��3v��.�M}��	�3KD޻e�Z&���1%V��r㛖��   �#�#�|�3���OظF8S���^&��u|�ƂN�e�Y����m|��}!��P ��y�ϫ}���9���nwF��k�k�P�#���(�d��Nz5�> ����| ��緭�߷|)s<6P͡����O}|�5֯���aD�W�ED"�V���;��Q�:�׏qp�:��1�~&�~3�q��:t��ݧy�DÇn��w����M�غ�F[sn��%����˗���Z�sa�pk0��S���>���y�9����B)/c�y�k���tkl'��\ȧ�I���Q�%
0��"�EK\W�K,5�6p~-���k��n�+��eg ��� A۴����C��W�/D6��&AB(�*�2P_}����õ�M����]w
����:J�wB�6谪:n�Xį1�ʰ�R�2 ����z[��j���e�w����֕"�vL� {�Mo1f^k5X^��i���S��V��Ր�o>[�'b�56�y=���0� Sm%+�U�I�Cz�F�Ӯ�y�q^��[�&�H��r��j��3�l=�����6���X���1�Tŋ�c�u�K�n�9��������V�z����rI��#x�эn����2�I4���^'1�=B�3Q?z�C7i�Y���R���X6^�v��ܤ��m�<\��=��X�v�P����k�Y:��Z���� �b�Wӈt���w�PK��QiyQs�ݶE�j��盺����!Z�-��{'��)�I���օ����(�yl��'i�R���c!.��L*]���S+j��I?P!����v��uw�'3�}��,j��խ橽"6��a̩��޸"=.��Q��¹r��>γ�3WZ��.s7!i:����u�O锱n�n�j���a��Q
P6j;�s���V�Pw>;C��"�si���N��.[�:��ܞ���4�Dl�ׇ���1Om���n[ۛ��^�˭�)GEk$l��6UDgM_f@�JEM��n�������4����7���i,�;��mI�|sZt����}D��1wv+��%]r�mu�}	�l�fde�w��umf��9�)��:�Z�i�ou��Quv�����"�DRw�������2J
�זS�ks?ws��<�*�2��5B�FLaN;������.��vgfm�"ɵ�k3M���δ�:��l��j�љ��Y6s������6ն�alՒR�����5Fv��Z���6��m��v�j�e�֦�Β�;.ܢHL�F7Y���ض֕�H��u����m�m;;Rl�6�;;�;lF�����f[v��ݺ�H��9k'	f�cK$���Z��%Yj@�,�����[hgk-�'6܄q\�����7t���BI���F�8!ö�2�L���2(:fI��-�;�n8�-k���we����K5�q\u8�bm���3q��6�mIɷam�-k5=uut)��/�����c��M��gW��h a��2*��*�log��h��QA�����'�~�?w�ޝ���3�={��C|ێ��<e�9V��a�����X�K"��_����q�^��Nv��{,G�԰D�[�U����^+��Q�t��p���J�@�q�c]�^�;n��rK�%k��+WX��T3=�ې'% Ak��_�������x<�c��M��fw{�C�t�"u}���AE@�(P&E���z�z���`�W˫�%��������<�w)u� F�yܖ)x�w�7����:X ��D%},��d�ĭH���fK�nd�]�xNC1|��Fr�D���"7R`=�����n���|̣����h����֚3�����c,f.ð���X�����n�I��n� �N���3�1m��0H\��[�ɜ��YG�V��`}ՊU�kU�y��?���uo��� ��D�@�"�"J�{E�f������k�'���=��l�����_�$`W�	(Wc
VX�Z]�H�h��Č��Z�\؍Π�Vj.�j�;��5��B�
����^� �����2*�����73W]��e�m�/=�^xl� ��=ʾ �"�W¾�W�V��Lĭ[GJ����Ƃ/�u�U��3��h�Τ8�@�Ӳ7:�^R"� L>"�!FE����4+3+��<��ol��*�@��$������Z�������+��F(��P���w4��^���9�
����4ݣ��E��b�	�(�$��/�=G��Wضu�C\�M/S�h� ��A��0��?X#N�a_F3���Y�1�b�N�7f����k^̲;�(Z��n�B�J�=��˦t�m���ҏ�狤��(6�ܑg/{�/)�\�| @�y^��]ӂ�yBnq�5��ҲЅ^�S��gDFs����MG7g�-�s#��\�^��Lgۢ�m*Oa0N�u�x�����P�ȸι�
���r&���������.�	��#��[W:���i[������h�W>w]����Ȏ"�p�ű��`��ٴjBQ�&���g�V�%�m癦q��L�6 �]��������r��-#\X�X��m�X�k�7A�g�:|ى2G�zա���p��zP�dTA�Iv�;�i�c�����Yk9��Y����.'��q�,���q�bW�J�:�CŚ ��S���sN�J��^���!~Ȃv��=��u�fO}�������W���DH����3�yo]ܥ�����٥K94�qOQ��:� ��t�@�wi|F�)P�y�H�0�}"`�a�o���Z����j@���@bY����l�C��|v/�����_!��:t�[�p���[��Z��oN��<��xo!�|��#:�b�:T���,h7J���ך�܏nCz�\�/qsg�9����K��Bk�i��f�� �����@�� �>����ez�C76)�h�#ٛ�q�n�#1��;G H��P?a}�]��L�*ʜT�m�˪�=���Y�fE�.���z��R������/�*v�F��'A|�9�gFo''�06A����?��:�!U��)��n�Ζ�tVp_n� ��$nމ�.�"��~�W�(Q�"x��ε��ziw��s�-K�67]��o¾��(s�(ȨDP�I_P�}Or�����.���!|C�|r��L��^�y��F����.R"�`�t��㔄�0��u F��}�H_�Aڙ=؇-*��=��Ԝ��z�
x
�"���$�_H�t�L�n_Z��.�Uub�]����k��[�3��,����룢�J�ջl��H ����ӥ�i��Y[yu�߷�#�A�������A����"(E$��EDU�f��U��Tʯ�m/��]V�����SN�ئQ�����cA|�+s��kul��Ұ��@��D(P2*#�t}�U��&kU�r�<���\��+�Z[�蚎Њ�l2'�re�֟=Y̜y�X�9������>�}��P���j�|�u� S�}�Qj�	��:t����Zh6=�{VF�0�;���y8?A�{�����g�t�yR��^�՛5Da��P&ED"��vMYB�o�h_�̓�}]u�cݩ1< Τ?cA:~Gv���(�=ِ�Dj�l]�V�?*����^m���y��4�`�e-)r��5���_��w��ݞA�dU�E���o��j�|�u� [C^�C39WTY�g�U`�+�@��.3������yʱ)��b���:���c�6<�_�ս�j�xB3� <Eu
2'\#�Su[b%D�0dU�kH@���v�P�5�D]��k��E�5�T��?N��ƂN�Av��f�g�7�o����hQ�TAB�[��]���NqH�}�P#Os��ޕF���N_���_mhB�ܷT�=#�1�nmg�Ε���`e���t%R�,�L]��ܢl�b���|m�{���WА?q>�\���e�7s�,�_a�~��`��F|�no�xE����xq<(a��gP�dTA���[����*�$%Q��DݓE"	����`�av{<��l��[Fi]��.�̸�f{���_�J_F�!|F�㺃T�gN����{�&#G�#s&.�#���6� ���GL4&E_%}_C�㹚�E~�3X�r���*�Se��]��ٳ�[������:�#w�!e��W��@��ܙ!Fh~2.����/0S�M���]�͂�C��!~Ȃ �0D�W�׻{ʞK�*��52(ξ[�5O�;��K��*LF�A�H���٪��o�&�6p�� ��B��@�%
2!��Z�����,�Z�($�d��������x�T:�E� ��O5��ӎ[ş^,ݫ�sLƆe[�h~��=�n=!�IX��4�a@l,gR�7&�Vu��]�dZ�n���޹x���G/�����v����h���0rsV�!�/����B�y�h2�7W^�h����]q�m{n^p(�]�������v��!�]�R9-���A�\c���]�>��5�%��m*y��9��b�����3��8y� �ܼaxe�%#L� q,lnB0Pe����������:�<q�g��N�����F���|}`1�T��s��1�#�zJO�������ɫ�Rlάm�R\�+240�m��͌������L���8��ڗ�,��o9W9��]�/GwW�È���{�`��4��D�!|F�_n� �}�+���/��A	i�owQR�Ƽʓ��:�c���8�D��R�ƚT��0����Di�u�O)W-���~�;+�ّ�2�5QT"��}"���}�����bN�ZD��>,����w�2�O!�|+�|B!��n�E�'cz��w�wU�DI}�5f���un}�>�@me��:����Nb(��:� �_i��	ݪ�컻؃HvH��Z�E$�ƣ"�Z-�B3�kR�;�r�Z�Ɉ�t�]�� @8Y��j�v�#kH\�I�5�}���OPS���WՉ. ��E|D��;� t�@Aݤ�b�r�#�|����r�r�c�G�����n�v7.�Xz�ò
����[�zŋ�W{����+)ȟ�X��y��K��(|���G�8G]lE�j��{��ݮW���^�G��|t���v�Ԏ��L�!�}@����"�/�Jă7���:�Fc��7/47������j�3ye�2ǜ��,�|�s�u����'�������֑*��8ƺzd�0��u�ܞ�굹��;�#�dL�K��cǍ��q��Ǌy�)ZY���@�R���9E��mU���{xW��� �P�"�P��yK�}w�v���t���$]KI�s�8�sB�������8��۷�T����|*������!�%W�!C�w3��5r�E���"�|G��a�:�x�S��~ �5}��wi|Fj@�:BO0���׾�J_��A��.us]�s�h��������B(���Zk۞�{��:k��b��P�a��?H���7I%T����Y��y��z�Y�z��U�H�Ȯ�F���aV���3�m3Sľ�9%T��U[���DJjvsgA׸�ۣ�̩@��������9^�+�Ès���W���D�(E$A3ޡ�&�;��P�#z���B���w��y���sG�:���6<�[�Ya�t��:@�ԁ����_n�� ��c��i�C��^�^�����L<+骁�G_H�TZT��x���:�q4ܚݳf6`�2�	1��ȏ�{],ݛ�wi,�����ӥ�v��9�}qv�ԫ}�!�B��ڈ���"x��Lb�P"J�L���P"���y���Eľ#59;��8]�����E?N�A�� ��/W��g���_wxP?t� �(P2* ��
Y�a�n3Ż^ǹ}�����f�C�$_!��N�B���'�=�-��f�ϵae;����>�]�z�o��#��}��Q4��k������gY�������\m�-��m�n�3�V6��5(<}Vt�v.�۷��Hg�ȈVQG:2F���h��ݏ�r��\E$��"�Qw꼴�/Z�y������뗚.�.b(�:�SP_:~Gv���J��9�ޛe+F��V�S^W�օ�M]rgv�]gT��E�J��{s��N۟ ~,��AȂ;���#�����5׏/��*z��U���.���"߈?D�Dk���A�J�K�;�-¢��k���>���Acp>�]�u�n�Fm}f�2 �;��U���s�]q�k�	�H�6��F��7P�}1�MFڴ�k���y���"���D�#�Jwi|F�r��n�J!��A�H�6��:ී�k�7.=5�C�j�3:K��oL8��#�W�u}"��"E�sQ{/�����<Ҹ�~�ۺзrFo	�WȂ2/�i�$_O��شw���S�����ٟD�ag��Y���	�Xǳ�[o2f^ժ�����1N���/w)]��ܬ�5��;�i����d����B�Qfw��q�'W
��mu�y������ΝB��5�gu��vT3n!��7zwITwG7���f<��L��"jf����U����7�r��♻y����aFs��Ue���k����b��ɩ�buF���}���ּcl���^"���q���	�о�Uv���R���}Ob�����޸o85bZMԇ��2��Ǫ��Z���q���=�ľ��n�ҷ�
�z�*�fMe�Z������������/}���P�HҬ�z��bu���X�,Iʤ�ǂ�%p�Y�V ��-�q,�Z:�l���rfG.;�v�r�SqY�f����Md���FxH|�9��?�e,��K�b�5Ĵ�f8"W37����r݂�vFA�&-pk���{νf�
A��9�K��o^�T;P��!���������y8�� ����#�D��Ιg�Q�H��(��ml��;�xŗ��;����{���jg�����j��)���_Vm1}.VP���]��F�%̿���7ڍ�*��[��sԵ�C��L�(A՝��J˷���j7f�V����5��m���8��Bs�<-��+�1_<�J�)�3�#��{\FER�2��N���I��w��Z�
S�}�v��-�re�SuAm���%5b��19��
۹"2���Ы�J;�!�8��n�q��ڌ'�0���2�k�f�+M�GqM�G8D�Ƞ��3H���mݙV��aH��(�V���m���D�������ۓZР�]��:�w2�pt����;3�Z�b�e�&�l��vK-�K)��j֚,�l�R;,�cfքN֋�Hm�6�&ݬ�Վ����������9���d��p�e����3	e����9���3Zˌ�JJ*N�D��6��ٓ4m�[X��b�D%��Z�c,�h�$ڶݜ���n�X8r25��li(rd	̱m��8��۬�����r�n䶲H6ˆ݉8"f���[ZvH�ciw�6f���v�Ӎ��(���NN[��u�v�P�β�:���z�g��5P�Y�a4�@Ual�����MSC���L���r���d�ѵ�f�׈�����c�:M�GC�v�L	���ݢ�d�q3�C�����Dzѥ.
��,Lܲ�6Y��m3l�zna�oJ���M'g��8ݮNs��i�7-�׬�i�W6����h@��XwFKM���a<��
m���p�n/T��/P���^:������zͽ��x<MS�o0���W40T(Ԕ�X@�g�v�]�ñ����㣃B]kW.�j����\<h/4����.T���Z�"���N�����J+�rpMk��3�͠B0f��,u[�	�R����Nn���H���']�^4�9^pǴ[Ϝh�x�/k%������ [n�WN��/�z�k��;t�����OgS�xy�K��hݺ�(�3p`�&9�t;�n'۴(iy�6�З�t�Y�f��Z�i��^�	�����jB���U��M�IZ�K5��}}�Ҁڲ�z��p��և���g�mj��v�V��kŷ]��}�d�y8�-�ҧciۄ�n88��,έ���v �ny1�닂��8ݻ{td���]��f�)�s���A��cnWsaKv	���Vk�l�o+���K>`�ȋ�m&���[c��h4�jj�8.�ı�ciXܚ�K��k�D�;(\V��;@r��/�!�Mq��X|d)�f����D����I[$.��Ι�3k�e�Hb�,�M�F`�:������2X�M)37bhL��:(���8�Rݣhf�r{\��.���qzb� �=�+���&6�Z�Az�]ۜJ롟1VL�Z#]�*���FRY��J�3uѕs��	s�%�%٩�-�.aH����T�n{1٣��MD��;fƌ,65�
�4c#i���"+����um��q��V�%�e���fb�%�$��Fֵ�X�ձ�3�$ް��nM��$�3;u�h���ki���>y<_(ju��\�7EBњј���F9m >խ�t	l��Ttx6"�Z⃔7qq��駞�g`<x�ٹ�e��G��vY�7�[���N-�i����<-�a�ue��5\�nx�)`֡n�L�3c6q�K�	��4UԶ�����$�Xފ���jBR��̙꽅.��d�8��Z����t%�K�E��w+Y����9���#�n�~���?���5�	�'���7c]���u�sH��n�%��2� k�|�� ~=��;��7W�㺂��y�Ӈ�^m�m��*D�H��۾�����"�G@����v+}�+��*�|_R����}.y9F��r��Y�o N�_F��7n���3.|��"����A�Jd@Q�7���w��USݔ�Z���#"/��_gP�����}Dn��ƻp���A/��o%��Arw��p�E��z��A�H���Ӵ�7�g�|�����ڸ'9r�9R�g5wiWi�]�}܇UB-b;�O�u���f
�����D�ꒄ3fs9��M����.��f���+�c��C(�%ܮ��͈�f���w0f�����G����2��
2%����O�)ARg#'����ݭ��1|�s�|D��#��E�ID�����+.���+���2�a[+���aE�ˣ'O�﫯�͋��o�u�z�Oz�\Hvmc��u�"J��}��s���Z/[3Ԩp �gR��&���
���u$;Ծ#����	(P2*+�~�����^�oT���{}��b�j�2W�D��}"dB�=��Z��+���8����}ڃ"Y�힪~�J
���2xP%�|�Z��v=7gP�#���	�P"E�"#v��
�=U���R�1zٞ�_+�3PGv�wk��y�5���Uݓj�|�J��'-k�<�[f-��U�.�������6��l�x��g�_Yo���M_nׁn��r/Һ:��'��x ��҈�6g������K㺾؃ ��zN\�r.���y7�0�W�{� ����}��������'�_Q:��_�����gl
�|?�9P �+�H����"��f?@��<��z+��
�vB�fjH^�w�=�-o�U^L�w�tWV� ��T%�X�yr��R���9>���1�:��ݻ�o�]m/G$R�1zٞ�@w�u A�B�2!DdTD�8.�Q�/o�� �����F��}ָ<3���y8��X[� N�@�{���w.�y���Hx����D�ED+�����r���U���o�!�jN��Ⱦ�_x��(Ⱦ�%}��pW{���e+��#F��ݡt �}qrQ�8'�9.�zl��i|���)����蟤��v�_�����$�~s���L^�g�PTc3�{h�� �(Q��~2/��wk�C��W�y�:@�#_r�ztuٞN=5���u�����n�5V:.(~_h��3h A-�����v���j��h-��η��$��Nظ��x��u
�Ⱦ�%}DI_Pޒݻ�O��m|�|����O��p�/۩�T8�gR?^�}q�^����B��v����cp��r��6�I\�Z���T$WA����U^�MU>z361@�ǯ;puaα�^�(�H�� �����A�N\E���{�m��AZcFl��y8���[�t�ݯ�#u/��Cϻ\���-��6��y�Í�9n�u7�Y��Naۣ�H�9�<.�Ξslp�ˬ/���o�}��Q�󔽸��6�$V�v��H���o�����_�<�%|�W��7P�K�-��:nG��3_d�����8Z���m��*өDݡ����#Ν�z�/�P&j�P���?� I_w�o��n�X�ޏ	��u��Х����I_W�I@/��A�A��Pa����[�� q�_N� %���7��kշ���� ~>��|5�-g��`�����n�� Ȩ�$���$y���W\_'T(K���p�/Sͩ�T8A�_/� �ݠ��v�|��wb�Y�:���
o��P.�/m��V�ٜ	��XH�^����S��O��=̽�ķK���P������.��|�����İElֽðO/��)�S�k�vuv�u���#F�o68:b�U�ӹyqA���'���n�>��W��bZ�k1�Ӻ�Q�N�xX8"n]�N��Z��Dkײ5�X��箩x�ֹ5/f���m%��0e|�Q�.�q���B^b:�����;=�'jcC�ը�p\.��ў��
���4�ۊ�*���ػ��G���~O�\�s��]��Gk�6rmn��e��V��UN\j�؆,���/_��g��e��u}N�&gv�+��1Yag|�K�o�[��mJZA}_W�fЯ��(�~�� �X�i�8aL3�A1��n]��^Yq�_n����F4;��o�8�-�#�/����'�|��_�|�2Pc��u�od�{r�C�j	rV�HtgZ?m�>yE���D��,���d.�d�㤾�/�����W�^�i=;��^)1��p@��ݪ3ȫ�@�{��Yq��,y�,�U��r�r�^�icҥ�x�r����YE��/���C:�|dTA�J�P'&뾢-��WZ�,#7[L�LJ�Us^n�C�<�uv���+��[&��*��P'5Q���}_IB��y���\�&���(��S�Wn�9�R �_a���P"D(a�(V]�}s�'����*�7j=.>�*z��9r"�w֍=b�,.��w����iۿ��e���Up�gG��a�Ο;��>�D\B�E̙��\����9|�"֐�#v��_u��o�T0Å|~r�ut�@�ݧ6�]Lq�4��l��ۤ�$�� ��؂2*"�"J.Q��*���f�����n��CԷs=����n�6��G�:��x�]S����V=�A�ŕ���@"0�(Q�M���y,?��!2wzmr�Rc,,����mi�_/�P]�v[���q�uEm=�쳆6o4r^.ܱ�&mf,V��ш�f�/X��-�fu�k�ږw�X��c9ʲn~��B�<�ԗ�:�=�|�v�9FS����:��C"J�� Ȩ������.���_��� :ּ�ӯ����k��(��Ԉ#":D�J��5��sʴ��X��Ա�Yc�U�9\F��!�뺚˻���\�-*�ԯv�����Bd������rB�+�p���aˬ7g��֔��cT�ϺS�9��;�7����wh�wE�y�٢��b�E���QW���J0�}����{�Y�;S �(W���U����z=����W��g�CYj��{1��cct�a��'v�mi���~�'K���:��W��O���;h��������0�A2%�z�>�[��<�V]�5�'a�㔕���8�zavo!��-�������!%�B��a}(P2*��"�/z�r�{k��\�/,,��Ÿ7�ٖ����ΤD�C��q9�-��\yʴ�3oKuǙWv 8p�GuW6��#��b�~�\F���:�@�ԩO�wƫ���W�@��JD���F�|��C���9=osv��ΒK��=�稣�gR�B�0�Ȩ"L�޽��o��|p�y�+��:Bw?���W��Cyb�5P!C���߯�1o`�`�}$.R��(3@��Ǘ�X:8xb&��W��vw�2Ud(9�ʿ7�e���2�$x#Gr��@�vEëY�qzF"�i�<���y˜x��9V�9e�x�Q�Y��i\�6�w#��eS�q�Bo�� -h#�_-�"Q~�
R���-Y������r�q��7R@q���Z��|��;��˅�fn؏��>x����y�=�{����������W#���X��Fz�>?Q�}"�"�?][̛f�x�0O��� ��Aw1跧4�L���
�TA�(@��L��c�>Ϲ��Yd��T"Ja���Ew����O_y�sWm�&n=ĽpG�C���W�MB��}QB���~���-c��>�!�|�?n��uצI8亿`�������@���x۞�A����DIB��D(P2+��{�<��B��Af1���4�L٧�ag N��miD�+�]�q���\�6�)ĽO�h��"��1e��fw-anrY���r�x��Mƒ�[7�%E�cffk�\��fL�S�w:u���ҍ�IA���nx��X��x���JQa�t�!�0�h�Xh�]ţnNݸ֑y"���&��-���ĉ]�&\��A�vp�n�Gu���m�W��	j���v�u]v�3�ӻs�.�{-�n�Y�;�qj�v�ƒ�糇�Z��^�AQۮ�vݜ�q9u�v]���]kƇ�X�n-�E`�j�y�,�K���e���"�M7�~�_���ev�hl�73Ne���\4��'mj&r�C7`�����K-���߬o���"���neӾ�Bj�^���&���;�ˎ��'�Nr���U���׸�"KH�_Y�S&��������x��@�ڂ:t��z]{��@�)$K�0�u�ݤA��:��ύ/\����q:�����8 N�D��Q/�J0�b�����eE���}��	ݥ=��]�y��|#�k������e�ۮ�k������@��PE@�"����QYW����B�s$��{j��|ѣ�Ǽ����@�҈#�Gķ+����x贝��V�6����Eq\z����s��m���	�`K��h�8պ�A:���A wi�H������>��fX�Aл��~�FTZ���BȢ#K���N�N�}cN�N�ȷ��.�����:U,��
��?T^X_�M�M���h��^e�	)ط6��'NiuY���*��.R팽}�l����>\�����{J{���]z�-z�G��g�@��ݠۀ��F�b�Bmx�(P �U�E:�D%��gZ���<����4|A=����5� �"����y�?5=F�>"sk�y?�E[�9?OxV��e���j�[r]���k�";����(�� A�u}�Kz༽_?�� 9�ސ�y�y�:���!q��;��:���Eo�eV$�){�P��n��Xxع����c��t�!�GG�6�դ�)����A�F�B#u��A`��w/m׳޾h���q&㙒�ϽkA��t��2*"J�@0�+�2�]���y��m�DP��1+9��lәae}���a�0�yϧ�(P6x�ܟ�(Q� ����|z�:�x�ˇ*�ͼ�L�]FpүWnr�=�j�)n�l^#X3#Riܦ���qN8S��hq��Y��\5�"����I���o6�U���X��mPo�v�)�ɍ�W#ܴ���>���*}����-V�ӕ6�@��^�=�~��6wvp�yZ���HU�N,�ov�qk�3sL7T�f����&�n���R�^!�(б�T�{}H\\z�X��ܕx[Y��K.�˧(�����*���U���cr�d�'�t��:��q�.}Z�l�� �}#��h���-�o}���h�Up;3*���k,wu��b��71�}�Ei��Y�:��P������bF<�ul�n�xa���8�"�)ٺ-w+yM2r���^�����3H�f<o�l�+�/��w]�M��c��n��G��p&������Z؂�waU��"��Osr�;\�,��B�=o]=�u�U\V���z�����WU[%L��xޫ˦V�!Ν0��r7y��`�YÎ6a�'�r�B���{�v�W��U}����D���G�#�WKL�{�Υ3b���V���
���q}+Ԕ�SQ��R�W2�͝�Ĳ�B����\�8�&�UY�|�R�#�J/^c�yؚuKuaL>J:��M�
�����WK��a��ɯ]�G�t�AQ9ǲd�&�|bz��ҕ\*MmЬ�J59HchEɸq�t7$�7^��w�l����=����H=Òj����Ή�h��3WNP���bT�w���)-�m�#��v�2LҜ�H�����ZNt���Hh����!!)�P�����ӳ���N��kqi@�A�rJIv�#�'6��!(�mlv��rɭ;n�!M��
f�e���kt��䳝9��R���#qmi9�8����!��b̛֭t�&�K�;m��enI�v���I�fYc4:�I��&m����9��6�G\f�v�"����֝�]��Nr�ֻ+2�4�@�Nm��X���m.���6�Ӥ9;lm�8����(H��P���p�Щ���LlQ;���K��f�Nرcnp���Y���ҧ3��j99gZ�p��Br��Z'��8I�q	�"L���Ŭ�bqH�rpHȰI>�kn��2���\CϾ_Y�Ƃ2*��"����vmK�+XE F��;�/�I쏻���ك�\�x�g/�Ӯ�*��\��~9��U0�%
2+��g�]�O|���c�7}�[ϲt9�+��P�#�9r��ʯ�P7H�7J�Z)�;��X����թ�5����Qn��3`�f�qd�AȾӧ�wi����ev疸��!���������{K�!�	��T���r�>n�HF�=���r;���E��`��=F���@�=(Q��YQ i����ȃ W�P����?E�P�~�����-��t9�)��r��1B($��D(��T�Qc�zׁ;)�7(/�P �� �:9{���nW���@��!|G{	�sn[�K�X�4�#�P���~��i^�`���(�s�Ҡn����^��X�b���	y�O�j��/A��'X�n��d@���]t����9Qx�"J	�QE�$���Α�)o�7������ѳ�~�/�҅|a҈'v�+ʔz��v��Ǯ�_$������TP�\[��\�8:�X�1\����8 NB���x�:B]�����OMx}���(v{��l��;�65�DgP���(5�Ⱦ~�����ϰ�_3e�=+��lg�����^��C�ψ�A͡FE��tr�r�a�"�P�{U@�_%W�J/��2�m���3v�����6~�:��(a�	�W�IB���8��^C|Q�_�嵤%у9�����_���� N�@�Z��^�Kq���o/���?�"Ja���TuՅ7 �YHlq�'^����^�,{{�6x�A��DP��i��$����2�M|�ձ��]��tsp�/7U�"Vaӎ�$ufEs���o_����Vߞ�v��v�Z�cwW�o����#��ARQ4��&lu�B�Mv�B]!��1��bsW:�N�)E��6^)�r���v�h�k�oU�P/���<Y[E���7ι@��qx��g�"LK44����IwhĒ딯	q�d5ۻFn�+;Q��2:��Y���^{^#sp<��Y�;�VN|[�B�J9J�v@��u����:�4f!�F�KXڎ�&�n6�XݲBo��~?����=q��_dinS����it��濘M�b�<�ԏGD^/���A��"�/�IC~������O�}ROY��^�r��P���B�A|af��"�E�0��"��f<�^���t�j]̙۽�?Oc~>����D��	'z�׶�g�s�*�@��D����P�a�� ��s��2���t�>���7u{\������#6��B(�(P��ɖ�w}���1w�XE'W���J�߳}�zk���'����gRQ���[ޟi��%�Dn��:t�;�#�BCs(9;�߫�R!.�N���~��~�o��/�*C�$_H�P�5�t�Z�tؑh�N�D^�%��:;O:�P]"z7V��M ��b�p��P �P�?Q�.��!��g�u{\���/WV5���SQ�QD@A͡G�Q(E"�D�u�M�u����_����on��=�uI���pej�`�S��NeKEC(ޑ�GR�Y���;ٳ�g�/z�6������ͻ~[YDqԾ?sC�y;���lFw�٣�	�*��E�0����Y��m��bξ���B ;��mi�K��gnym�lmkށ9�Ƕ�b��5xb�W�IB��
0�@�}��;\�Y^��������I͏���f��INoX�����([�>Ta�߳�|A��"J��TA�$���o��*}@;�@1[������،�s�G�{����|A�ȯ�3�(�/s�|�F����mcY��`9�d�2à��<C�.��u0��Kc��3!<��|��__��D6����979��j��/w�]�<��l�!V~�����Ch"�+�Ŷ��:�s�~Ew.��(��_s��y��wo\���g�@��X��tf�r���U��ڀ�#�#=,X �H��@m��ChB���� �n��pG�,uH���]�at�B뎫�T���x��݋;�\ј�YD��M�Y��̭�J�p�Ů�>�Փϸ<Ӿ��囙�)3`R��[��z�?p3�YyYe A-�`���w/�U�Z}\x�#=,Y}H�!�NE�ȵH�?
��� �H�'z���^^��x��e��,��%���� Ye��{.'�G��q�wt����7oѹ�}g�@��X�� Au�oxt/#��iu�I ��ʲ���A��Brq�suˎB�tWJ,��ƶ���M�Mt�.�=o]��ڱ�u,M�ɑݲ�-����{����mI�Q���$�u�������
 �[j�m/�d��]��������_-�"���z��j=��?
���	��A�!jQ�����*�� �W�6�������b�:���Gs�lOݼsFe�� �,|[�?:d Cnō�6�2љ!΍�i�L�#}���Ǜ�{��ͳy�O"� Av�`��(�LvVQ��ܧ�y	iZ�v^w���zj��%��nb�2�)M��ᣗ�՗�;4P�_�f�zO�Ŏ����$HWW}���a�,��,�VsNd7����J����mK�q�v�*ﾰ~1� �L���/��hSџD�wi�>�����Q�LGL����!2��1��j�@i�,̤���Vg\}F?�ۙݲ��[ �ھ����y��;�x����a�g����#��X=Ԁ!�B6аwU|F������WH?T@����!J̝'�1~=�<�<A����� �,���/��3��������$����>:Gl��x.߸m;��j_
�ƥ��Y��/{V&������,u�s7�M%��=( a��ֻ{����=Nn�9�3�&��n�WM:�f��:�a��-��L����*�
��v��	 �An>}�g���%����W�y,��mcE�檯}z�ה�^(]��������EnI��y�@�E�'��h��E��w�RSb��1��s��YԈ��]]t���m�}�>U��Ub��bZ��&#l�	+�큖i3yZ�\uu�E��&p�1��`q�8�b�0�eb��u�]+m:�6%��y��i�{V8g`ك��%!�X9�n73������SH9��J�lZ^& ��=�:�s2�v5:-�4Cn�z8�v֖��.�[i,����:���V��@)���۴����H��vls:Fj��M���������
�3RY�MLФx[��[ͩ�m�"»�Ve�Qv�.�i�ϋ�����w&�x��Bq�nԾ$�Eo��V���_�ʱ�u,N�p2n�c��Am�!y�\>uhE]A��Ҿ �7���w>����7S٣2�|l��,X-Բ�C��B#�o��z��L�m��m�㫎���
S�t�rϲ�T��?w�g+���QڰCh!�ׂ����,��e���7��|*9�݊���%}��k��=^Z`������:�.;�y־e�6s�;��b�������w{�G�S٣3����[�A�"�����w�yn���B��+B��� �mU�c���F3���y����R=��|�-�H�����m�h��?N¥�˽RZ(��Yw��U_�ڼA�� ����[k���,�=�T���۴�$y��JkU�ߟ�<���U��\�;R��,X�_uڵ�j]my7)��J|!�1巍7��Tt�����ݷpx��>!������	%zX��	�� �L�Cz����]��%-����0� ��� ���� ����o̜onS���{	z�=�38/���5�[���B���ؔ�1��kZ�A�Bk��AV���Ӱ�g2�eˢ�|A3�X"NO.��_�l�	���	e��?6�_ź�-����d\�<z���ē�������鐈m���پ����~oO�����Ҙ�v6BX�>��Y�-<Wg]!�����L&��K��}o�'����r�,���[j����{��x�o)�љ�3�o;����������y���L�m݂t�<ֽS~���a�=2��F��fd��a̻�r��{�Yo �,�c��{�gƥ����![w�u�:d7*��]�vUo����YK#��=�y������cL�g�A�p!X,u`Q\��r��JAS����C5����ڕK���5r=���֝�q�&)a]�J_]2!����e�:�]W��.>�^ ��E�(�[j�l��=��N���h��&�� ��{�j{-i���A�J���Kt�?:d Cn+3�q��z�7�*Z'�{�ed�z�]x�{�X#z��@m�����y%�o����=����$�KdB8�32�:�eI��b���X�rZntR�X���O{�2ο��2�޿~��~t�SfNmT�Ҷ&�a]���Z�<�ٴ�֐�G,���@��Gwnf5{�]�s;���c��Bֻgw7�~{	�����x���/��WY땎o�q���N� A�۱�c]s�ך��[�/[r��2�]ˢ�=ھ���,�� �Ր�b��7����LB�r�A�!�':.^pZ�٪XJ��%"�գ}✬�5:u���+�������C#S6��(��b�e����<F�՝�	����!I�m`�]vѼ�{�[6���:��{̙{s]g����ݲ�u�x��XlM���Hh*�X$����{���٣�C���/�#d�e�D2�7S[�֞�Q�Ӿ5@�HW��B�WVh�Om���E��B�bċ�wBuBqn�l`��B��_��:�t�j�mؿ�͠�����;�� ̻�r��V򮪁m���LGb��?ڲH,�F��N���P2}%}T#d��5���k3^�a+��H��w���^�I{��lό�����~mYg�[i���7�r�}b�o<�����^ձ��p_x�l��u��26��#GAu���ZE�_P����k�ݡJ�����/8Lq��"� A=���fU]w�O���Ǌ �ذM�,G]K�����JyW�7����d 37���{8{Y��K	__�R��Z�wrdݡ'��O+O<3����*���U����˕e�ћ5d�A#��9=Fdx�k؆���<K�oh��=�uukc��n=Ը��g��4�7���f��a�N�~[3|ݎ��[ �]���X��a���n�BK��u�����f�����#w\ö�ѫ��i��43T��� Z���*�D3����2vX�Y�����}N㭦.c��^I�k���\TS�e�2�N�NL2��pb-Tfz�Ru�Kӂ�����2�o4k��X객ܭ�2��3s3n��g�f��&��V*]�Vw�1�g7Q/���<[�Z�d���~N骹�/#���R���"s�nn�G��I<:�}���j������+b�ܮr��ٲ\cn������x�`WuQ?[�Tb�W�;A��ђҗU�_p��̱����9ཚ^������B��\R��S�RE�.�ɢ�9�����w&%��/]{���
<W��lX�%�U���jʌ�F0�������q:��s.�����b���n��Mx��$��B�7v����u~�����nU��5�Nni�8�Y0x��H�y{5��
�^K�}ngp�C�<��)�As��am��kyB��m��7w�r�9E��tK���S0M�����*z|ݣN�s�E銇k�ϒ��u�o�X�q�K�mh����j����+�zP��p:
��)��UdL��y��6�N�yon�Ĭ�����3��9�[T�2L�} Z�B굆�7i�&�J�裺��_��<�H�?Z�wyM-�%�ӻ�p�̦���H" ���E�\tGAm؉Ҝ��[���v�s�,[S3m����J� �N\gh�Ĕ��B�)��p�	�Y�'9�C�-m����s�%)�.�gv\�Űݝ�؈�r�f�̎��Ü�s�E%mZ�G�Ԡm�N��99E#n-NE̷�;;9X�3�k6
2�I8[&Y�2�)%"rI��f6ӎ�6�v��Fl�K��Ř�������!�ΔVv��L��)�i&�m��,�'��I��e��Y!��"qpI ��Hp�ڲp�����;;C�p�ru���qӝ��Э�-�G\��N:"' ���R� �8#��[g.8x��x�<��d?�Rj%U��N��aٗm���@��c�2B��n��c�8Ԍ6å�d��t̪\�L�F%W -hE[5{\X�с������WGn��H��ƣK���m� m=Sۧ�r=�q9Fy,�0��R��$�Ҫ����ոV{F��*i\��n+���1���笳�\s���n+a����C:�``d�vh^�أ.4�fFʎ��#Sn�a4+�J�Lu��ێ���v�-֓��y�k���`B��<DL���`+1��j�E��%�81�w�й��II��̪�� �]��i@خ���p��'�� �t��|����ѫ���n�V����ic0��F�<g�bU��tܙ7�!85��O7f�@���c�M`Oi5s�������vx���j��mM�^݈rUs��ź���7�!�q��{�6�a;b��x��`��7YwU���n��>�t��X�rU�{�'����:ˎ��(��W�F���Vi+5Z��f�,%�r���[t��m�k�K.�����rSWt�Ҷ�R��lqNI�	e�1�hD2�y�e�.�q<-۫D<��nŸ��g�cmRiv��N������ۧmB���2���=��;x�;c�0*�7K���lR�,ްdZ8��j;��ņjn�["��ɸ#J8�u�p3�m�{e{b�'�Յ���>���^�����M��\���:��3X����`V�x.�ݎ�e�ux[Ձ�k�.���B��T�1%o�7��!��>}����;ҖS`�ư��R�����mH�#�]�RO#���q�tp��`��q���v�`Yk�b��4&1�VP!31]�MmrYc]�*�V\w!I�ۖP��愎ͱ�7�}D���f��i�Ҏf[�s``��*9@�^��Z�q{8���rM���ŏ#K�6Ɔ,�2�&�LmlS%��L����TV�Ř4Q�a���	�Cj9��2ں�Q���{ʺ�/Us�ێ��a���p�ST6���̱����9֥8�.�F5�棒6�����b흗`k�]���˼�k�&ڋ��@���\�d��I��k�����t^박+m�[�����6MAXּ��\�l�Ӗ��dt�NS�ŕ&&
�印��F����p��l��k�QKџU�Sm�	\�߿���-�m��u��zgb����˘7�4�'K��A۳�ꪬ��?F~��"wl�]n";�~쾜���B�ܸ�����L_>�����t��L�Cnł[�GU ����%���R�~��� ����TQ�~��d��E�w��v�[��!_ub�wPG�!Cn�n���G�Vw+$�W_8��p�fk�,%k��e��m��[AY�r��K#�z�.A<Q����Ϻ�u���n\׃2���@������щ-�D��@�����At��B�н���Z�r�wu&�p�l��;��?p=����� YeKmn���5�S+r2m��WtAEݒ�ѹN4\�<�[6��q/�$ @�8�R���_�zD�������L�����)Oga�f�R�W�����,ͺ�U�A��H@��_X��,��?ڲ:E�A���w�[�#�%��o�ތض�2������/�N�wR.i�C^��XH\��i�o]^��÷B+�v����b��|��@OS��㓕�#�o�=[�5���8x����t�S�A~Ώ���Dfe�`�t�?6�@�݋����?V���iN�}�*��o��J�|A=����A� �ՂHN��z�����W�A����` ��[ӟ8j{3��5����.R!��݊�8����gr��A�"	m� ���г�f����s�uL�}��ܞ׃3�_oW���/�������c��D��~�}#�a�I��374
ms��n���*�����V�n��q����fo�L{ʴ}ۖ����~mU�1~}�y����qR��-ug���z!ڔ��<~m�!�?�|.��T�Ywi}Ҹ~|��9��O��-���X�}�������6�Sv\�V��PDd���7A�A���R��6���+o����^>�\�5j���.Lx���߸��a>��w�{W�>U�[�n�;��MS�:r)�\�9.Trmf���3������ ���,X-��Ȇ݋�V�I��:�A�Ŵ���]Ӆ=�Ƿԩ|A>�U��+���A�dVCi[�� �۱e����'C��'9����5���.R ���v�ChJb���8W�z�h�\=a����X5ݜfL1WB�X�l��&°RV*'@w��/���@/�m\�ϟ,��Ckr{^�Om�y�*��|4oe�=Ծ ����Kt���3��%]�nGWw��b��؂5�ػ��!�o��J��{9}{@�Chg~ߟ��xq�~���,^v��n�;�q�_0�*��Y=��;��lMur�W�e A��m���|� ~ŗ鋔���H/�@���ھ���,��ks����������XS⪯�/V[KT=�݃y�ՙ$���vJҪ���a׮KT���h�n�=$��KCҮ&����f���K���@�_7XA��m��{�W�lAY��rp�I6��~�� ��__�E��6o�}�|�|�@�v����SY\f\gB&VjGL%�su��$4m�J�7q�f�=ol�߇FO_e���H��k�6M�r�{�����)_sK文7-�R�L@��@�����-�D[j�,��w��^=� �y���>���%���z38 N�|� �2K��7~���:������H~m|����ho,�>2��'���y�y$u���T���r��-�_Am����7�xVY�^��!��g]/�-����{_
���1��b��N�"�uS�No����h"� �m������e��w����W:�9����e���z39�|�?�Ŗ�~m}��Z}<�3<��uF��݃��+�v�^tz->��M��f1GKD��f�]�k�����٩Z�{�?z,�g��6Y��]�c�� Х��4M	Fm�kt]��+3[�*%V#�nŀi�|:9�mZ���9X9v{u��=V����kZ���.��j��eu�6M�v��El,�7ePa�
A�+#����d2cmp��b
�8$�t5�z 3αS;��4�]��̖L��u���f
��fc% s/h$�\�yN�x��cչ;�^��#_�(X����2��N�]�}�֌D�'V]�f�YC�y�Y�ͫ���剺����<��/$���~��<i�D�u��ݨ#�A-�`���Yd E/�]~�*��s) GBޛ��E�f�c\,R����C�B6=���c܂ v���E�Q��ݭVܦ��sk;�*\�Mɣ3�@���D�ذ[���B6���ޏܽ:�ex��/��w��[A��yN�&���h����`�k��vH��Y��������1�����b:�\D��n��v�=���6��7rMn#���Ì�J�X'z�_:d�_���p�=��'��кiU��� ��6T6D�g����/�9[&g\���������?7�sAY����}ܲ�bS��}4np�����ݽ���4גŞ�@��HD6����_Y�	�O9ڧ�m�L�6����jUFi��H�ܿr~�Z'�澐�~hU�˖�^�d{ȏ��3R��l�i��.��C����,_��Ʈ>�S��H���訣�{9Y( Ye�^\�/�x��`��,��mز�/�.�f��f�s7xi�7{�fz#�j�;Z�wndݲ�,���\}K{ܙ+�<~�-�u'�}�?%==��F� �������~�p����O}y]�� 6�X �H�2�������®|��Fַ�S���ׯ_��G� �r�6W̳��m�[�ڌ~'�w��ǿ�v͖i��I�Z�];n96�is�|z;A�P\�jR���������b�u-�ܚ��t�Czs�|�{w��s®��`��K܆v��m|����b�!�,�� �ڲ=��F��Iھ��~���uǯ���ה���4nr���"��-�<|��m���Gk�q9�``�;R�֠�����}xj��Zڢ�Z%���\s��M��H�;��!���w��N,�(ʹLL��v�z���'��L�4�-uG�r��B�����=u�y�%z��]xA��`��Yd�g�n�9lst�BĆ��:�����d!�s�}Y[�3`���^��N�"
�_r'�ܾ��"�? [j�n�e�j���W�yw�������Ynh��	�� �v,�H��C�WU�Y��ܺ(�4����֍p`[\c�l������}�b����n���0c�*Y�jZn�dCh/������J����(�������msk͠��ڰCh Ae�,}�@�rU�>O�2�����}G3�M7XN�}`�aDC�$�+��t���3PG�
�ؾ��YD�Nko:�/"�&t�Tu^��-��8��#C>-��ya�q,�1ܴ$�����[Ar�;�=��N�_Z4@���8?o��h�����f�:�c����F{+V�w��~���#N��9+m���0zn(�(�C��:{=~˯f���)�$��Y�<��q}��&������v���Zk�+ϸ� ���m�n���M������H�F�����%T�����}��s��U�b�t%������b��6�ڬ�t�/,3���6#��WC�}^�/�^�%�Y_�j�K����s���Ynhܠ�����������e�D鐈m�`�K�"n��}d"/����A���;�8����G����#ZY�[�����dHY�/�-����!���J͗ƒ��_����n��m����ޤAm|������A D���4�lF����� ��F)�����zz,�4nru|��Q�I��?���#�|�m݃�n�n��!��Z�^��ϳ�h"��lw�͞�{�����W�kA�m	�%^�<�.������g��/5���r��Cw�}�9��:Z���M�tp�e6� 8�7�[�����QE�|�LK��_��g�韾��~Y}�m�"d���F7=��D����A:�+�L��^W��5���GS;a�����,q�E�,���\�w��p��%�4vފ��fۣ�9�[��׸�Բz}�^�
�Fy��t=�p�l1�d�{���t��5u�k��L���"�j�j�dR��8GPunW�L�qì�6 q�Zk�����ۡ�ay�M>��~}*�ij�V�Nm�Z�=d�ݳ�X��x�v��䪈{��p^����`�K�k�ofپ�w���a�����w	�{�)��/�̯��g����n���^�`�4��+�r�݋0B�'7��_��\/yOL�sF��@��ł�y��I�S����Fl������6����]�W+0n�)G80�ɳ.��6xA��d�Ye-�`��B�ksN�*���ݿ�� �2�{��w|5�Z�n�����̓�:[Wc��{��Fs�.:�b.��#�e������cS����nP�yb��߶t����~�nh�r!1��u�]2jW�?>����Y�V$�����f4/�4���b�3cɴDbk��걘Hb]���3�_�g�����-������p\��bOr]<~���ͽ�A��	m�!�Y�X�������^�}�n����-����0�=������=5I*��^�y*���oI۠�w�5�ʲ��x[�y���v���)=2���TW�����w��4�;����z��!�r���E� ]A��=ܬCk�Y���W�k��^��׾�O>�4�>�����@� ,nł�|��E����"#�Y\��X@�쿎���Ås̒�=�tl��g/�?/��xR�X��W��F�����![v,�G�}��j�!_eq$�b��3���1m�߅����i��`_�v�u�`�v���݊��4(-���Yt̶X3"8X�`iM��F�pnwX��~A�r�A���|A-�a_zI=�"�sF���J\������.u�;Ԉ!�!hYn�Qѭ�O����>"f/��a�zgwW��O�2�����dk��g��^�ގB���dMHǈD=hX-�鑀wA�<�{:׆���̸">�J�̘��mBV�J�5A�Znm���z�:{���1�t�,�GX溺�\���������+�^r'�+f�]y&(Q긳9U������'��Ǯ=Y���s���3�*�ʶ/0%�oJژM]�Y{L%؇e�w�(�e�ͥ��[�Ug�롃;j\B�j��,�"ɾ9�U��}pM�Iʎ�^u;�M*ͽ���;�&�է���/�7j�9~`^:|��/-f�E�(��L�7\��ʣkt]t�Y����X9��Ҷ�JZ*��B�����aM�i��}ٺ�	��)U�N��`[��2�a�}E���"�*w5�k�3&���r��L�̬]��+(K�Y@]C���]UQ��Op�P4��m�	�Y1�έ!��wRp�X�cK���G��j�Z�RU�+WY�Ni���8o�V��2nutgu�1�mm�Y�F\�]�h��Zq�jh��|�SX���2�q7;/W"�v�z���-�&�܎��36�����gwy4m&p��e)��jlʸ��ش��^ʫ�΅}6�O9��x���e��׶�DK�wZVuV�R�+N7t�΋�ȸLY�[كE�9�U�YQ8��(��'\��SNu1��ۙ�����6�<�
�����)1R\��*.5�J�5-�ue��^U���wfPÎ�5U�Ä�l�=c�:vWm�mh�۲��7��K}�]lE����d�W�K����a>�(�P����DXtV��i���Z�F��8���w9b�r{�{'���zR�0�r%�V{&�TF~'����I:����q̲C�� ����dI%&ۤYaC�m����9��IH�Ѷ��9��8�DA[v�tRs��8B6�"�Îɶ̂JD)9'@#�s��ێ��''I�N:R����)ʹH!9D9��99 �9H���s�H�G8��p$�(�����ڛfBB�R �G89�S��H�$��.��-�8t.#m#���8$%�� �D�$�Np8��Сӎ�m�C� �-�B! ��m	�H�m�%"�H�9���C���A�D�Y�Cm@JKkm���L��b�99�"r�t#��89$�%�r(�#,�.C��%*� �.�vH�)B�Ztwq\Iv֢��b"0E*+�����������c���ޥ�:d"k���,���q�i���J)TW�8�,ڱWޑ��a��wnh�P���<7���8כ����+��W�m���L�Com��+��V������g>&�;$8��e<'���u��e�k6͚�xz��G0]��� к�[�e��Ӛ�"�g�[m���֫c)]m�����y�><B ��ذ[��t�@s���U�\������o�5dc�d�a�g��m,�-�`����m7CLC����}�=�v��v��@� ,nŖ�_����̭ dx,%|�2o/���Ϙ�o/2̍넫����̣��'���G͠�ŖQ����T��u{ea�8�-����:d.{ݛj��o^9g)�����~<����Zδ�	Yi	����&�I`t�R�\�E��o��Ghu�+&��͛V��D��
 o�[�va��e�����ޑ1��Gz�ك���ª�1������|A������M:��ƫˏ�֩;��}�O��v��@� /�]�����դ{����#U��u��7�UY����i�:�:K���p����x��7���5�iR��˟��rRz�۱�e���ƕ��un�;��A^um��]��P��q�[ݼM�,A�R����{�����% D0����Z�������z���_C�B!�����x�B��%�|�@�
{�Y��̳�~z�f�]y�%��s7Mϧ�ܷi��@�|}K7p�v�FmjX���k��7�<���R�����_�����N��J�纷[���� �g��|3�;7�����b0{ݼv�u�/wp�ݦ���C@�d/�wlͥ]�7����{���z�� 6��C�N��.�ev�Q��*O*%��	�O��}�{.l+�d���Ť#9X2��;-�ŕ�����7x:�gc�zu���{��=z�~l
�SGA֙��w�m��m��C�vڂv��	�#)�&�t�c/i��3-.eܙc��%�Է��4l���7��Ȗ�cC����Ө�n1��U��U��"���$2�)..�	���nyz����`��Npfv,gӅ0Fݻ5v����d��b��7'Z�K�l�v;�#���9�.���"\�3�z������k�k���d��]����r56�z���3�1�]v�":7���[�ק�|�e�A����_}<v妶h��3��=����<aA���_��|� 6݂t���z����;���-��2 �=~������ɿ^̣��?�VA�E�zM�}vڛ^ޜ�������B ����> �dxQ=`��n"}�6�G�e������@��@m��6�e���j��ʑ(���Ye| ڿ��f§}���N����ǈ@��\lN�^H0{iT!ۻ��DL�m�������B�~9��.��W珓~��GA����,��[i�*��#��c��3�"
)R�|E]U1�Y]����#n���ۮ!��� X�7���W뷴���`�K��F���S���9Nǽ�"Vg���صs�`����#��7AY_KmX#K~ݣG�CmL�u����F�_oU/W����c�i2XmK!��-�he.�iq��iMyR�R���V|�J�v���
 ��}[�ͅN�����l�y��ǈ�n�n��z�\����.�t��_N�A�����������,g���)_�>M��`����V> �h Ct� �Ր�CJ��;�P��`�R?7Al��Ҫv�{,�?{�`��|������Dn��c@7^ ��m�����n��!�	f�_K��{ݛ
��?Jv�h���#�AF7b�n����a��[��^1@�]j�H����GV�M��Q�+L���Aثt6�1n�;v��������_�Ծ ��ۻ������:�~x��ق���49��C.�o��:�!�@��m�!� �� }0���b^|4o?����҆�u�*�a���������_��@�wP����d��7���j�ؘ �mY�!�@~-�<�L�U�)Y��z��,j�Y{�o][������zN���P��R��1e�f��yֽ�-l�
�X�nZ�]F^�*y#�<�۔ ���kf��G������Kt�)��D�ŭ�u�z���=A F7b�!��/G9�+y�s~[0VW|~��`������Oh���+!����"n�n�z�kǝ0h���A�����I��e?{�,�@�!k��0�w�lYY�B͋�����'"lfɨ����g��ֹ �n���t����ۮ��(�l�� �}�k�Y� ��W[�͝W�p���kf��B��׮M��s<��<�垽ڱ�Դ��0AݫF�b}�t#>#|����=~�u������m< �r�ƴ,�y������|���ƾ@�Y�۱`�K��EQb�O1�v��Дn$�x�����a��h�Z����M�,Mڸ������/.��EZX�b`�܂#z�?6��Q���^���m��^xP$?!Df��){�ɔ�G=�<P��Dj�]��E�=���	��O�qR�~�,���M*�ݭ�w��Π�\���y3:�m�pvc*^G�8� �B��۰A�U���t��؍�u����kR�����>��.���٢��Og+#en�_ں��]<���;�Z���M�UU�������sD�\B�n�d�ۊP�Tŵ���>�&�� tv,�H�t�f0�>�\�S����9��2�-�/��z���'9ܙݲ�n��c���0L��Eeu����@~9�Vo��U��Ju�G�� �v,�]:��<�U��߫h2m� �HKt������wO?M}��+��]��u�Eep��V#b����W��7�P�B4g�1��݋.WȷC�w����p;ݲ��6�,�_[U�9v��V��hQ�ׁ����h Cur��zc�>B�<��(��yW�xh��T��G��chX�_An��)Ȧ��i��눡����4��u�Y��)cT��;+���yL]f��u�;��EX[�\uǑ3E�f���}xD����Ϟ>;:Flk�� �����-�iS���u�λ9%�H#�iU���p����,�z8�Q*���z�i�b��m��oظ�j��s꧌/�zD����u�ŷ��3�t���g��U�[]\�0�2��V�uk�<Q�Qt�ܧ�s�9V7����8��4Z-��e���dSV�q�:���Z�MDM��k��1	��O>}�'ݣFի5��]�c���mRWK����-��;�j�K���޾n��o|�����F_���Gy�o3�EeqeHfJ�������#���ՀCin�#�c7
����x쯑����1����9^�����X ԁ�Aۍs��3��: ��@��� �����|ʹ7%��۷���\��f�o|��PDnŖ�|!�!ۿ�7��m��7|�x���/�A�2N��o3�h��	���!���=C�;�#��w/��,��,�1��G�
��\B�6��	�o
r7�����"d Cn��Ch[¸����]�cEz9�����=\Qyfg��lvq�ܶ�Ջ�%v �V#阬��e�� �[j�}��ƺ�fhu�G�����}U��x�A�Ń/�!�!h_ź@����z�/ɱ^^J�]���Ҫ�r����u�����p�|R.��@�Bx�x��:Uv�T�q<�X����>��kTߥ���-e���2�}�� e̓�G�˷Y��j>?q���;̳Y��ir���w.#ؐ �d Amؿ�t�L�w��i�w��'��#~��_�X Ԉ.������@Y_�p�����x[�Z<P ��WK};����l�f��_x�UFoxV�*���u2�	n��!|Cm���e�k�k�5^�|j?f]���f���3��F�Ye�m}n�W~�r��ٜ(�IU(d4s;py���ר�#Wcj]K��v n�DIլ�(�zX���ўw�1ݫ�R�ogcE���g�g���b�1׵��dO�+�k�i�l��\x��q3yAm���+�zD���A�V���+�p�/D٢� ���v,�Y�J���f�  U2��t�@����C��{º�~ͧ������L��粠V�kwmUn{mN����Hd�<��{d�Sk=�Uv�H����1c�*+˿���s�V�s٣j?g�[͚f#��fr��#y,�� ���Ci��{�U�O�4t� ���,�.���i�>9��������SxgI�];Њ�����ŖQ�����E�zZ5l�,�}֭+���p�u����_x�~ɷ���F�?t��0�}|=�>��<ww�g��s�X�f�{k��.��-k��[U��)�y�2sj��z���ݣA�&NR�z�y��b><B6F�wv~��!�\�������M۱uԸ�3�����g:_���y�n�O9���������.���
&����k0���_�Ǽ��#7l��[A-�s8�:�籫��v �u�����|x�Fk_7XC,�>!�9��/)�P���!|F>����˙8uKy�	����z���V~l�=j�q
��߽�ʥ�*v��ӏ�C��N���n�tu�i�{�Z��g-[��!��2M�R��syLIJ�Μ4K4�&�|F�ϗʹt��w�u[Y�7϶���Y>�A���:��z�<<���]�� Cn��Ch$<�cˬ[z�v����;RkKz$�8a��;L�7�GFh�0�]�*�=�A�ݽD=�,Mڗ�VW�t�pXΊ�4{9=G�	�(2�ز�� ��"v,�"+�Y]�e����&ؿ���\�ê_��E�=��z�A��� � ���Q�;��C����h AP6���>?7_w8k=���\��v.6F�W�^��/� �A۰/�@7^jQ���'�ʳ�����K�Ŷ�+ޝ�3����=� Ⱦ���5��Þ��v����'��m��	n��"{�#��v���ê_����{SB�q�g+���� ���m{���1Wu��+ε��7�g����ϔeM����,yα%5��Ҽ��:1���s�6�/�\��V�Y/�o��p����Q6����Mы^��o��^���cV���-�b���%3��l��ìA�`Okc�Ǽ1���CUQ����X�k:;�T�fNQ�l��"�oY�v����I�߼Ho%ǚ����w�8�̝C8ӥR�;��i=�e_�βD	X�d�2^K�H�<ϭ�N��2^V*�-�cyb�)0���G
N���^ك�碋P�C6Ht-���M�E��x/kv����y6�n�.ւ,B1G�����D-��^!#��l�̲9�ޥS��[���؇���Q�si��ͭg	�.Z	�YY���V�C*���Ϗ�|��T����,�A*��[�R��Ȼ_m�i� ������U�1�f~��ۖ�V��w�����Wx=F1D�+N�:�UJ�=p�t�e��O�a��P����T���0��u�)��O<i{�]G��*؎��2��8r/]e�6�J�a�.�]���]�;�)DhUs�دV;w7���o�'�Ë���T��/
aؓ��гt��r��kX��]LuA:>�����/��xv^����-n�]������}b�0��oCr��y���V�ѻ�ۀ�7[:=��~Wz}�z���<��v����hC;.��*�d>�1�RjW�7i��]]ܩE�+���H��:ޞ�kaܻz���<l�V]���+&R\h��;S�=/�V
G=c5k�t�Խ��o�4w3sj��雖3fk�˺7F�;^�nݳR�}`�Z�9H�.:��(��8�㨺J˳����:��i9qrNPtq6�C�Y��8���6�C�;t(�((�8�Î��m��D��\�Arq�,��h✈���H���$�!8�9;�
"Ó��8�3:��!՘ӎjr�$ ��#��I�.In�v�i�N۴��å�.9 �p,�J#��(�H�%
$��nrNr$t�J��'NI�GE�ee��r\P㙕�
]��A�9�Dp��M��plۭmv!ڶj��mݝ�$��������\Q8EHAE��9�u�GrEt��ܐ�N�QND�m��8��;���8�8 ;~�?�.�\>�y��Wk���]Kh�rqr��8�<���y]X,�'�u�݀�ԛ>c�g v5��O`ܷ����ͷ:8eq
�t0��V��!Ԓ7's���s�-�pOg�7eN�{&p炧Da�+��Uyx9IQ5i�px�-��)�Ӯ��e϶��8	ƫ�g+��1ۆ�f�v�J�f�;7��sX4�Mܥ��4�sc�����_<���<���,G/����^7��C]u���u�%�U�twMz�PGi�.�����C�1�{'�0In�L�3[�tȤ[�.V�irZŰ:�	.�W6��Ka��=Y�w^x�h�[��B�Q�5%�J����=H��lf�Vi��R��7/i�4;[vtZJɸ��CMml�ƚ��kIGc���p��4n��<�O>�=jn9b�`8:���լ"V�F�,���=f`�.��		t	�7"6Z��S��#�rg��d�;�^qU��m����{\l�9c��ƭ��_P8��� �n��V5\�w���7�8c=͟.�uvb��:z�pA��3�E-�콶v�Ź��<[��dK����us5�mZG�����vɸ��ɉ���1����3���=pVюf������]uZ:[\�������:z��Hq��@�ʝ��m��M-i��ڻ<mж�8�ݶ��,/Ԭ���t�l�Pi�E�%2hV�yW��f���v�aYbE��s��GYYe+Uv�F�I��-�̑Y���]Cv�/0�٣0,�P��-�#pD��۱�dD��|}�����#!;X�S�.ւ�%��N.�p'	<�X������:\���d�%��h�]��x�����C���N��֌v��r\N�OV.[�8��N^2����tj��-L�+ш��3u6��6jՔ�.kZGV��F'���s��N8�Sx��1�@6�
�r�͵�#�i���â�F���8כ��ec��wJ���W]��ٮȻij-�貎B1�טk
�թ�4У�j��7V��t5,��5�l;,i��G��ۮ�t�,n��������)\���I��4Q�,&%��T�A,4��S���nu�2�OcGG�j6R�L��[.kt�kY�Ik�������6��GupX�]�bGgFFR����l!����yV1��4Dk�Fէev��Qp�Ve��7;����vv�Y�\�lْ̬�J�	���P�&�Bى`RNe�+n��-<?s��Oݢ�>�p�v�C�B�t��.f���½�p�/��~���L�.��D}b�!�e� �Ղ3�y߭l��ӫ��Ε��Z�q�<��詳G�� ����v,�Wv�[SE�h�+�!:]�u� �d F�w�mC�c$��nf1)߷���{SQ������#�YeŶ�A���j�Y��y��R6E�g���Ԁ �鐾�绺np�M�<��/p�@.W޶O<5�Ka1�ޭ�F��ܾe�|A-�`����s���;�
=�XJ�#��������><B ���_ź�L�p�S<�cY��밍"R4��-*�������'����s�8�ǅ����B�洑ћ�ߚ[��?B!�w�t)��r����^�h��X��b����A�/�g�Am�!���G�"��JF�Z��ʰ]LMvy�s73�(J�9|�U���3�+�j��nj���#�HӒ0��k����!�ƅ��ƦIQa�������B�������6H�<<��	r���v#���-|���x�	͋���g��k��������q��C���jlљ� =�f��n��Cm	t4�mp�5Y�%�Ŵ�s�R���:kی/WA������;�g�x~N~�n�oݹa�E���`[�(�V������mΒ^�M�L��/!��H��n�!����_Vg�l0~��ϻ��}���\�vp�[�/1K�x\mr��(�-��jZbi��b+�P���,�}zq�!�@KmXI���y�Sz��+ʹ6��A�&�}����uCn���|D�>���+�p�UE�ؿ��_	r�3��0{�M{���p?L�w�_�'��:q:�'5���&��N����Aݫ��~矫3;�W�����f���HN}{�.܏�k��]y8Afwfî��U�mf�Ead��9We8V�Y����J���9�\��s$�8c������u �|Cm}m����à��/���7�_�"	m�	?8�C��d�٣��G���������K��t�%��Cnłn��m�v�Z����Ăw���~���1�F���g+#z�7HAm�}��Nxz�Gϐ�n?���^1���T��;u[���j6�E����Oc�]ee�s9b��E�y�჻V��AW)'I�រ�W�^�9J�B��j��F;�-<�ɑ����z&��iy?/y���t,9Q�����	� ���4{(q����Yn�J�OӃ��X&s�c�գ�,wna�|f)��]n�Fzw.��_��`��#��3��A�/�n� �ڰCt7˔=�[�:A�b�JG��/��s��z�{�����X'�|���u�����3��b���{��k�j�W篩/`�~.[4�WKSK	������5y�T��V�W��9�,����#=.�=@�"	m�����<�BV�2�b�9�V*��w��
�݀�����M���@����׸��� �B	�~�9�<p�9�;���(T�^7h�c��MkFA �ZU�*	�łvR�����_���]r{�g��=�3�h����y�z�!5mBjY@��V��,���:W�U=0Y�H�a
�[�&oi��$.������|A��!m2��3���<?m�_�#�{s�,u�D-����U�魽}U�(�jl����� A��n��2�6Щ�n��qo��U���#6X��͠��vSg���<^=�����9Y�+hy�xJD<p�	�j�m	e��-�[�ާc���O����}5��������_'L�m�����,���������ۤ�󲻼y	בgR�/��{����1X�i�|�UkmuRn1`�9Q�[cs��oe��0ɨ��+զN�b��X
�*7iR4o��{]l�v q�0�Dvs�t9���5� ��u��[+č�|m�47Ń֢7[��J��Q��FN����uv���vB�d�05��f;���h���zn�D�]�&����pg��V�$��p���i{2��m�t�ܛۃ�kI+]F�6J�L���[c�뿈yu�2Ƥ|ݘ܁\��z8�`�������z�\D�8���E�ݰ�,��h���]�Ʈ��a4t֮������{�K�+ ��e���Մ�ϟH�56`�����q��ױ'���Y�K�d"w��[��S���S�ο�n;������zW{:���݌/W	����h"����M�Z�`�i��۱��[ȗh�jyg��������xyZ���!�����e�|~�HUJb>���~�AY@��Vב�������������3*��a��H���mذ~-� �鐁�&���^3޺���^AVf<޲����_��h�� �3��� �����KF=�19�!���J�������v�q���fQ	�0Yf��iYV�"��*n4	�#�`�H�Y
�������nH]燕�=f���۫k~#��;�L����GwnZ��u�8�w��Yt��7�+'�����í����q�v�h�G��hp�J��;�zM�g��x�z@�^vu��v<�W�ҷǙ�Wپ�$W`�� A1򰖾�Ǫ���-�39���`�PԫM7���^֐�lv��DL�>!��n���Ck���}5����ju�><A���`��/�,�A �Ղ_:Dƫ�WG�X�ř)|At�@TQ�>�=��IY��}`�).�8��,x�Ӿ�@) ��r�|�m�����*t循��� .j��ݚ���^�)l������(f�����P7Le<�9�X���X�c�SV�p��by�[��r��}��;J�ܥ�Pe�|u A<��_���T��ɬ�}�S�ۢ���VR:��>�O{e��j�#��7|����Zy�YO*�����}ZAL�+�}ϻ��IY��}9H]2���_2�*�(�vEc���e��Ŷ���eS��Uv:��v�l:l����EkN��n�ʪ���/��y��m:�X~�;ᒽo�~<�ug-�'���n1ib��~��wv�fP�]k��|�><B �w�u��2o�?z����%BG��!�N��~�_�-�^n6��L�+s~s7�w�XcO� f������!hYn��~�u��b�N�)�d���e����#�L�����͡
l�-r�!נۢ����Onذ�d�-�1�&Ce:�����u��w�Ve6����^"wl�뭢�a&�=C�k��|^u��=�v��"sB�u"�B!�b��@�����=�S�zY{��]�ٯ=W��iכ����L�+ ��E�o�.#\������C��	��	�b�n� �dj�^��o���_�=�ǾW7dgs����L�զ��wrdwl��Y�F��I�_��b�~�x�mU;}�L2ìbZك/�!�{|�����
ۅ�M׽=ۼ�c�sr=�W�5͇/����H�����o*�{2u1��`�я�N�'�W1�b����dK&e>��21Q�\@��;�C�B ��U[P�j�ϴf �gvo^U��m:�q�l��=��?l_2ρ�wj�D��ǔ���H�B�U�b�	Y����s�7Z���֝Xjf�፶�3������_�?d�[�A�
�Ot}��znɥ�xy_X=�鸜tK�ՠ�!�.� 6�,�� �ՑZ���SK\��h�|p����u�[~q�<z��1/n`�����q��n�~�]��qg�԰L�2`��Z3kR�n�dwl�:K�|�,y��w�伫�i���ѳ�=��;̲m}�A���&�ŏő��b�}K�t�=R�>�z�7d��<<������.�W2{;G�ݑ�o72'���u�c���!�s]}������0��.f�/�Ǭmc���/����Z3��2�Zk��G�Tsfx^#��ʺ;'��uJ�������V���;�h�g�l[�dX6D���]Q��z�`0�o/��N�D���v�Յf¯�S�hNM�h��mc�<�s���4a���f5��ctV��]F��"l��Z�j[{p6;Aď-�����������"A&���l%���mh�l�86�A�\ם��$�\�Om� V���`�;���#�5�����1���gps�ٵ�M���P7<ݣ��=3B��V���68Pؾ�O��?b6�ײx�ruK�=�7(����]��N׫Z���+����Z:��B ����6���wn��S9m:�������~�d����!�.u��wv��#���g��!�t��[��gR:��*)�s���M�4��+C�r�N��eQ���X������6/���Y_�k1�2כ�;�ӳ��z��1�.`���!��e�D�2!�`X�>⛵�t���i�������ݺ�)zWiu�n��|~������&�}f}ݼv�uԴM��v��۲���r�a�<+��N��W��e煫��Z&֥���Ȇ휄��~��ԟ~z>�5�D�XZ�E����X"KZ��G��D�i��U�A�(B?I*�F�q\�s�w�<=0��/Kt��%�'y�|��B6�X?���Y���5U��7w��E�NX3lmf䙫֨�VpPv��e�ڵ��\d]����S!�.�Zw=��K=n�4�:7!��.Awqo6G��e���u
�w��6�S��.��ߍ���_X�Yg��R����+#�|��@A�b�t� ��:#Pi���t�y�c����س����\�C,�Cm}a�Ŗ~�>�yf�����X��l��0�	m�V���x�ʬ�/��׾���D\=4`�~�^}"�A�ˈD6�����!�ܯ����w�����n�K�^��]7��<A3ܬ��|�?x��J��!��nҳwHQ�m=�����m�U��v��2ˤ��B2��5]�I�y�����@�#�e�_�!T����<����Z����_�;I���� M��|��(��m��r����Y�+����@�\j½󏉮�˭ܧ7��w�O� 6�X�+��:�4Ɓ��";�ł�"�B6�����*���z��Y���^U�)�ݽ[��í��خ�hV�5��W���/<�WU�*��ɝ#K�o�Cu�e�Sr�bvD�����O.��z٩��B������y�r�:�����@��Mn,�HҸ��7����Q���7[l�B�cc&,}}�{t����-u�[2���u|j�#l�����.���d�Mg�"O���:s<�Ue��G�X��Q�o^\:ϯ�o6۸�7
(N�5����3�e�wb<��W�BS���"�����/\7�^�rߍ��)MO��,z�t��W�y��EBJ�WsI#�%�,����+gA8�`�X�f��l����
YY1h�顭	����	@�ؤ�W]���[L����m�ɜs{3��a�X^�&$�)f�vS����-me��w#y��X�g��8�J�B���ޘȱ�N� ��1�K�s�����������3�X>6n��7�`�%ٞc�uR��9�)t�8��)ot��a��/Q9�oMvغ5u�Q��^�z��l��N��mb�LKky_]-ܙ�5���(���齇N	0p�P��X�[W�C�W$��M�����	]m���GPyC�˷�H��(�k���;)���5ZL���Y7PRpEu��ʗ�ɵ�͡����B�<r::����GA�	����Y�Z�:M���n�>��՗G��r�ѬZ��U���ٯ�C6-�¡�c��r��헦�[nu,����M���A��C5�L�9���<�Y�U��9�E ��"*w��B'	�#��DS����G9�\%��ݺ"�S�!:H��p.:"p�"* $JI"p��"G"[h]"D\IP�Z�!:!$:$�:"$莈��;�(��#�I����BH��D�$�:m��pD$Nĝ�ȓ�q R $"��T��G'!Bt\G	��Y�QIw�E�I�HD�QQ�Br�8q)e�Yu�#�Bs�s��	�'9�G.AI3Gt�6������hc*�"(��\���5e/:�]7�۷s�~��߄�v��Jm�@I��m�.�l��*f�Ū�}���pmV_�ZےH���6�����cֶI��_���R�.�r)����i���#-�Q��,j�EGq�7�j)��n.�n�����<�=�����e>��a�.ʟ�����t?.}��׮��{��D���rt��WtA��n�j�傻ӳ|�����G�vG��jcrmE�K�W��m�'/L��>��_� �o�6�.T����z����o�5�,[�����@6�n�m���aw޵_��K��P�����o-^�;Kn�o������^ϵ:�������FQwN�U��|0E�'+a����[T{s���F|S��&������ENkZj��Z�ɐ2M]��߆��>��n�h6�o:�(�������xܛQ;��IC[A��p�����%U7<kF�A�N�\�ԝ�D���jv�詜�ϛv6�n���]
UvM�k�	���M�k��ۛ��r�OrK�Q�cɾ|�J�}��!%6�m��ѶM�����d_�:��o-^�;Kn�o��ܛ��u��ĵ\��yO��G�6�t>m�R�.�<__I���'��6�f�}�5�m|m�]������3Dt5�k�wno��X�䗞��f�m�Z�ob��lؾm��n�ʹhXҙ<zF�b�����w�|�}��h|�ݽ��ޛ���#o�+Gt�k�o��|��/���$Q����W9F�s5 �����Eᮝ���U�-P��{~c�.�����u��C����-��)�n5�\�kg�|r�����]��X�%�fQ.�kԐ�j$ƋB��L&f���0Lr���Nvuq;�O��غ�F��cc��< mչ�t�� Gr\(�M��n�\���:�f��b�W��=�ڝgBǜر��P�A����s�c��z��{]�$Ò@�<�����Cz�=������YPg�qt�2Z��)��+�qS���Gx3�8�*�}ub�ի���ݞ_v��ʹw�G��%͒ji�\9����!��;P�ɺ�6ַ�l[Mm �-�Z���U:���Iy�]�o!�m����7�*�	����	��m6�mK��Y����7+W�>�����s��_6����n�>+�ݽ�k~��C]���'N��fI54�u�{G��^��_���A�m��:����3�2Z	��|n��z�㗞ټ��n�͵���&z�x��D�뾎ڼvkt@�[���%q�Yڙ��F����״W[r�UѢ*���}���m �����y��E�nt{s������F$��Ỵ7W͵�cP�4��~�{\�h��OXZoP��^�w�F�h[.�nCT4���)�n}T��YS=����tg����NzVGJ��7�B�Bn���+7���ӻ����O&��p�᭠�~2s�ku��N��� �6�m�]z��ؕ�Y�8�P�[�r�w�7��[o��oWT������o/�r�>���<{W������k�ʅ���.�鴻��gD��m����z��L]���E�������O(��w�k��m��9A�7����T�l�ؽ�W6�\�a�Ŋ�$�#�n�stl�!XB�Сh_��ϟ�m��k��7�y�[�8�*�W60��_��M�6��A��h�j���B�leY��{����u���x��7{5���/��n��w��.�����������w�u���j��l�kN1RDq#�V4�/-�����a���,p�D��w_v����]�$Y=����w�Onf)���r�mM����\����w��m6�����ӯ��C��=��w ۦ����/�fj�b�'��$ԟ_������]�h鶛~��Qc�^Z�{_,W���ǵz;ٯm���o�6��[}��>�O�v]�+!	C[�suk��Rm�nkBWn:N��<R%RuT���{���]�m��}��t�޹=Qm�j^{��j���������@���İ�W�h'}3x�.>V��M�\���[_7������m���.Hg� ��m������ڿ�ʦ�]g���lªl/g��Or:m�h7@�N��fK�ɨI_��w��>����'�-�\�z�:�yϽ,������_K<2�f�}=��a�ҋ��~�A9Tn���Sޞy��>�����]����<����m)oj���/������m_*W^Q�ƺ���3�4>�\�޼��|=����tu�}9�7<�?L���������L/]	�����#nh7��Ie�h���v@]�6�@~�6�����W*��{]�Ƕ��:V��o���_6��������2�x�̩����:�6�d�Qm�᮵�����M��o���7b��߾m��W;��bE��OY�~��ϗ�[o�6�m/
���E�<'e��A�_|�}����Q�=����CW���g��kG�YU��	� �o�6�3�\�;���˗��S���'�M���u���m��E�'=Ԩep����ci.��e�˭���q�3��yXn�f�f�孱@����<�s@e�+�����hُ�~��+0�I����7ö�^X�1���IŌm�#���v��ƜJ�iX�&f�hy�˳ٶ�'-��a䌰���8�i����Yu�\��������8��6t\iQ/^��5lܜ��m�+E��v�@�����T�]��V׫�m�(m�]�X�f)4�k�t�d̤�6J�v�V`�B���㫵��I�-�FRp��_����~��nڑ��68M5�;X�9�X歶=�F{[�\RlU�����Bͼ�وl���>Q�n��Kհm�l�R��۫y�|�N�Sm|�_�=Ր�B;�����;�uu��w�S��9oSm�4?����߇sA�߾m��쬺��uk��`��mzG�Sm.�]����������&3*�JDk���[j��C[3Ǉ�.#��F)�w�)W��m����m��*_�ͮPL�V�^�S:T��ǫ����m��j`��Y�̿>S�~Qɀe�����pmt[�
jdV�1��@�i�f�ՅuF�_ ��ᓓtm�ݐw>�Ndwu6�� ��~�vA�����n� 7v�ؿq49�����X�;�����}7C�����k�=�q���rE٤�nU�5Z�6*�Y�C��_Z��~��{�q�a���$���^�p����As���V�ra��ǽ9m�-�s��:5��ޠ>m��7g����u۾v�7'E=�c��g/��6���>��3��i���m�}-wdϵә�d�]��K���Wd�}�6߾m��߳.��g��йt��}�{wܭ0����|�6߀m�c�w���~_�_�ɇ�Ta���
X64ͧ<E-q�[-s]��8^����v-!THWF������1��"�>n�s��|9:)�� �:�{�ׂz'P܀m��|�@���ܷ��W)����k�A��s#���u�t5���Z�ޞ�<���y� �6����e�h��b����eҘ�גO��nV��foF��[Y��|w�օ��ܚ��fY�_-Ͳt�Q�K���A)v*�������6�̱-����i�{����m|��m6Н<`����������7_J����W2]�;�L�������6���߇͵�ʹٮ�|D�n���7�y̹5��KU�ﵴh��,�<��r4n�WT4��.�Ø顋\G��W���� �6�=q�y�v{�3�s���I��׽i���ǽC��/\�	U]w��5�������|�t��}�����u�J��{�]p<���e��W��n��E
f��7�I���tl�d��¯}w����jk�VKU�c���͵�m���Q�������W����I���l������~���W����䔏v�uɵ.���,Y���i��!W�z�E<D��mޮ�ͬ�+�<������%Γ�S���.�c=C�&�� 6��T.Vۧ���^����u��OOE>�r�z�m���NyƇ���
�IZ�v
$|�3���Kc�-
M��SV�&mT
���.�N��?v��F߾m�.����s�Mw��j�ˬ�2]������鶾m���`���BlAK���s����vx_E���nA��o3�����؄����m|9o�%��c�Rp���L��6}�	��ޠh���x�B*�����x<�$��h)w�v��jk�VKU�t�9�H���� Q��' �n������(d�҂�J﵍�Ny��_{uNr�s��$$ I?�$$ I?�I	O��	O�rBB���	J�$�I	O�$$ I?�$$ I?�$$ I?���$��B��!!IRBB��HH@��$�	'�H@��$�	'���$��	!I��BB��BB���(+$�k/5�> �]�0
 ��d��C3�4
            @    T     �
   T@� �    UHP�B PJJ	$R�P�R�J�T  �	E@��J�P   T�E�� �P"��JT�QHB*�@*�
�P����T��R��%%QR�P�$T�J)T!R@�  4�"���J��.��J=�9(�.��	Q��
n�R� Y�P9����F�A��Ԋv(
(��B�� ��,� J���U���@w �}@���`�<��x��w"(@4�΀��� �U
(
K| �U�	ER)AH���� n�ϳT�z=H�z��/@��ĩ[���4r��­� {�@��� �g/ �h4�`2� ��C� � �}� ���N��@


x���'���{�M��l�h �`�� 
�Ƌ� ��礅^  �r����+�T��r� ���)B�|  �J����$��RTO�[��Q�� /6��r Y������8=��Ӫ^�9U$n�{�ZԞm*uL��9��
�  2��IH��Ԫ�M�s���Yԗ�q�R�h�T�wJ��O=J�=[S�����<�\誯m{ۗ�� A7�  ϩ�TJ�UT�
*�E;�U=�+֨���٧��{m�+��E7UB���]��J.-P�w:.��UCRR�R���T$�T|   �M$���@�8�T��*��uQ)��
���rV�H�ʪ���UV��\ڊ�*@ (�  �(� �AR�����E.��E.l@� ��H3�JV9S-G1�UnΊ��n���BX�.fU�r"�
 �x   l��iT�{���:�W�^�P�jJ�3���^!ݥ*�{�Is���Hn�Pww%B��q�*��rz6 5O�I�*R�  �~F�%)Rz�  ?L�T�ԡ1 �%H�   	OԩB� 2�&�)撥4�@ x�������_�������	$�xC&
cΈ�����8�<�X���HH@�d��d��	%����$$ I?�HH@��BB����>�����5U����_�?���u��.J�3�D"���xNN�^]}E�6�R�nTT�kl�3t��K&Q��{%ГsE�ش���2e��7+o4l��o�Ne���Ұ�y*�Rk�^�ȷWW��f�{ �sP5+b�N���������&����9�l]�۶4��Q�ŷ̥��	�B���*��g2���N�)�պ�9KXU����	�^���f�yj�fe�}�
��b�X��/^��ͼA4�b[��27j쫤ml;/7v
4�4+6�]a��j�B^���U�[�{��	O3a�mEI뚓�[�U���w����ڊ��e��P!Z��Psj�ݭi���i�n����%J(�a�Q�"��T5R�ڼ�G4s7�-�m���r�����5��]���6���2�AH݈5V�ڔ��X�w[CZ�ɐ0b3dnkW���{X!9B�m��,�'E	CD�aܬ���Yw5�Ę��H^z�V��z���=�0e�F`�lX��5��eU���cm�;k��6ŝY�hk.�ڔEJ*0�uӽ��ͦa��4��k$��1�N��+uG��Z��w&�0KݷW�ɨU,5��Y�f;O/]�;wCY���M]�����*�-U�ꁚڄ��/C'rC�ə��lVM�Yf��0q^n�]�{p;���cTF��/i�x���{��ҝ`X曁�ܧ��q��RvF�K����Ҵ�vef�i��X�̗%��ì���ɺ��4��uT#.V��7�yc-�M7k0=f-�A�j��Yyn�/���E�$��U�6#�-T�6��%ʋ�^m�d�Z!�2��B�T���pJ�fӔ���pe�D�<f�ݘ���l���3/HH=ۡ���%<Pp����oJ@��Z��͛��<�z����u"1Z�v٪��x��&��)��i����8��u�"������n�M���^}��2�?�ۺ�ٲ�n�ɒ�r��գ{��e+b����M�kN$�՗v4���g^��+�"(�R�n\E<v�f�Ȼ�%Uaї�b�3i��E����TqM�D���i�wKD�5����]F�A-�z��n,��{��6�Į��LV-�6Խ2��pKF�Q9���3w�K�[͡J�mL�D�e�~�:���
����bRB�̫t�D��cU54��%�3��xZ�,�ԖFd�2�R�ų6^av3k.ʷH�pEQ��ܕYr�V�K�f�<9z+
7I�(☢������llb�1n�0�M���jf�ݣ�f�2����v
�g.Zɚ�iSX�9$P�UHcM�%�$���{��^���#t�)^�Kf��[x�%iR�TH���d\��@,�͢n-�*��c��j�]`ڬ.�Bޠ�^ʨ��-��L[:�[k�x�/N����۪yf��UwC��e6��ХWA-�m-]u���(f�i��"�M'�Juj��V*���ev5�KkSu,�EsjVL�h]�
be��;X ��f�����]꺎M�*�n�Kwz���x�^	g(���:�f[�r��Xun֭�z,�hӦ˭��Pr���D�8Z�hk�uU:��q�+UL��Bu\�N���R�24ƑUo΄�lnI-7��-l�v��Y���ǲ��U�.�E��E娞ݝ��ԑk�&�	w�N�-eg�k,@˪ә��/�C�����M�R��{��e�# ��c����V�i��v�\�f��ǛG(�e]�ĒFn�P��lnd-m�˫�2���1�+C�]�]&�m
�UЙ�(D�VdTb��j9f#�^ڢ`�ML��j���L毉�i[��
ն�Um�c�y�t���y�JD,�2�������qe԰�B3�-�����3n�L�� CI������b@�+)������	�u���jz�רLߝ�Әu��y�y5iү���+n@dՙwKoJ1cM� �%놪���Bwq�0�t���cN��H3U��lx�Xً3X�ln&+f��r\FE>�/j'H;ڽWY�$[)\Am�R��N�Y�n���-f��N���T��ҭ�ˠl��`�04L�ы�Q5f��2�B�j�KC&MJ��n���/4ؽ.��z\N��D�:���p��;�5�dr���i���.��Q�9"�oP��e�&(��X�o(M�m�nTc��&�[5��ZR˄�
�������B�wSa�F�x�;fd�V���G��V��V����c7�zXlY��Ywb��0&0V�wf�(�wm��X.7M�r=�'�;��-�6�2��"����j��gu��o-Ͳ��Wf��x�3�Co[kZD�uCKen������+r��˶A���&+��2;%�"������q,T��m�ݰ^�#ϒX�E�!�ڢ��Wj�9R��{,���(Dt�$�^�v�����ȫC6ѕE��ͻ�]�k���6�!��Œܭߥ&/*SVE6�49,����!V��ͦ�;J����n��	�R|d{�fHb��]���ݻ��/M�l�T�~WQ˰-L�M��*.Ժ/3��6��f4׉��n���&��̟U���Q�"����vm�1�yV�旙�]!o2V0ѫFi���e$�����Y�E�Z�u$���z��Ŏ��zU弽f�\;d��d�E]��e��j�"�i�`[pB��Pn���ѐ�n;Q#�%�3e�>!�x�Zg�6��iZM�0^a.���J�h��S�E�Ա�y��/ٟ#���EU�v��v�%m�35*h!l"sm�0��0i%��Qmmk�]�%޺ZoC�r���M�5M�]P(ˈ˪�%�ԜǨ+�ehEDUe��g�f����pQ�������L�t��t�.,��mU�8�̌ʽwBj����#2�`�t~�%O�J��H����,�۬�F���n��=����[Щ^p��mU�*�q^�ԡ�f�ޭ�ܭ�Y*�۫e7�X�e��QvV��<�^V���7v�1��a�v������,Y��we��kV�Zc-��$�O5ؽɴ�J��sv�̭�.^9Jָ��u��7#�Z�fD����b���m]�*}�RŮF���!��y�]�*^b��{�։����2+N�W���z��M�M�{�3*��ܗ[6���Z�[	l��eq�W��h��N���k�l��q������a���$8kr����"�af횽u���F\���Z����5q[�T��ݸ��^;�0��çn�4��`4���;�T�m�n�ӼkJt2[҂r�8���]�9�I�ϳ
��@�A��%������[x���j�G�e��'2�]�J��)sz�Ӫ�30j����O՛Z,�Z�*^
��-5uor�:{�Ej�e�Ow.�Bߤ��}��Z)������iU�͆+B�a�r�k/N�;[w��`�Bn��e�UY�wb�t�Zwn��/*�R�w�V~�V��kp��n�4�	3�ER˳jf�<��)�s5��m,!�t7M労��;�FrG���z�f�koa��lN��ar+��a�E�z�2�nP�r���n����k$���u�s�h��Gҥa�g.E��GD�i���R���������ߢU���+�����7w(���ۉ͇%�Ѣ�FV^V������$�%`��St.d�D�6�jQ�cdm(򅳸#�;�^��;V���c.�~׎�ͧy&�c6�[Nn�.�Kw��`�iS�//,9��A�iy�e�S.�POn^1�6^���*�Ĵڲ�,���Ϟگ:x�y4f���.�ڵ7��@QZv�W�J�NY�"��^ӻ�uHF��]\�M$z&�����S��6�f�@Ph+Uw&�ke֗��;�f��q��6�.!�ߪ��c�Pl��,�����6ZW /A�%1VEf�&���
�&�[�8���N���rf�כ��h��R�UֻJ���ܻ������ɅZڪkCb��x�Xw4텬4/j�V઎�[Gfh�yz�m�m�Q<�H�~��eO3uf�kh$����z�M��uaڴtJ�ܧ(��.��*W�d�y�0�JlC�(d�%w��]9!��cJj�ݫm$jYj��ê��h�zA�"�PF]j��]/Y��>��u�7�"�����1kWV�9Z ���$��~J��3��4��� 1FFk�jõ�ʖ�2����n�wOuBI�k�S���2��y/u$�����omZSdv�
�V\xq;#sv���r��C�7&9BiX�P̭rj�)��~���e�3F]�3ځڶ#����[dF�]���bxఊx�n}z�YuD~Ǐl�qU3N�EhZ��Y��<�x̀��VZ���S�wr��+%\9�Ec҂�&
Fr��iq�Jf�f��u�ݢ���Ѭ�[�5۬�rcԓ��r��a\�[#��N�eGz��n�n�U�ج����K��Uk_-�"���D�ж��:t��L�)K��`jE��U*Y�e���d�06�B�\y�n'����&$������ޖNf���	V!�fJ���ww���h�H�%�a��9��t@�0�C~�(���5�u٤�	]\u�$��K��U(��b��z�JS3(^fjNi�Fhu��l�۫����ÏN��t�)2"=�	b��f�۔6�M��F·N<q����PЕ\7t���i��f���N� Q��,v�W�@��!;'��-F�ũ�U�B�iB�����ɵn�q��b��y77���V�XK+���Ok^R7YX�j�^7�I<yv�Y�J�a
=��MW�V�ͬ���Rxj�A�G.ƫ�y*^�Vn$��~�kC���B�4�V�����Zf�����9����X�y[+fe"�wWm b�G�nG>�cU��ڽ*;̪XJ2��70�Qէ"(,ܬ
�t���n`������v�@m-�[��-d�n+�
9TD�2f�n�J�zo�V]�ʹJP�&Yđ�B�f5��X�hy��/ZJ��N���tٔ��r�����c�߰Mٻ�凕K;Q,y���{{y�r�I��-޽�-�c$�n�1��09.:k1�GAl��cl`�ϴ�^���nV`66kV���1\U���A��^�@�[/
�2��Cl��T����UR��M"���6�f	b+�h$�6�c,����dU�xU�����e���b���m��m"ô��V�Z���\!�b��[��#�3ҋI� lmb�Z�ܯ�,Q3�Ղml�3*�%-�oX/wU���g.�Y��@�xww\���+�1[����r�#r��kon�J�T��x���{f�{	љ0nm�v�~�7����V�ۼ��j���*���ԑ���t�C&CkTGK���8ojhW#¤V�R�	V<Xf_��n[�@�wVAْ�SDZ��bK�wR��ʡ� �����n�`*��]�L��iU!6�փ��fJ�姖u�R��@�6���+�m��� ���5�m����0Ѻ3v�Kw�`��U�
�P�vf��F����ѝ2�T6�&��ʸ�`yOi8��Uh�B�!sN�	��*#ak��cv�Y{�W����c��ۥVU��5��@���C$��IRwm\�ͳ&����X�sC���q��1�`f!�dXn�e(�;�]L��dj�Sݻ�q�.�m�
��u�������vҺ����<Z�;��L���u��L���Sv�,\�. kv�嗺�8����V�ʷ�7�i�;�Vc���8iކ�Vj8u&���LNƅWT�L�����
�1�;�X�F�Mn^�V4�۵B�Yx�;�6���uL�z�6A{J���ņ�+&j�{r�5OY��52G�	Ѷ��`�$X��wVΗW�sZϖ��Ί֩=+B�����P��ڒ����u'�����hYi]S �����rc[̂�)���h�/6�ز��ݚ�4���{�R�e엗ӟ^C3�f�Jgm�d���᱗{�/ͧyL�ef�˴u��M烼��U��y�����Q������F'A��mU&e�1^��[*�^E�l��Zcv�<��ګ7#p�諹�Дt��#I�^�A^�n�8�T�ya`�;�jQ;��5Ud�ߌ��&�P�u2��#p'2]�»�fCl�D�˘��H�W�6:(�x%�=��6 ���ݍVۥ4��4,)D2��($�Ga2��UbM|�7j^�1��V-б^�ՖC5T�̬ݻ�o�/1e�lR���f�W�/�F�-G�V�\:o��!3Y��+��C j#n�]Q��
]�)<Ӫ�jاt.�em�F��ei�	�´{"md!���ԍ�T^`���9,:�{KU,��v���qRF�ͼ��+)ު�LHb'o,ꚨ�ݷN%�,��XY�I��UV2�jXX�f\6i5x����q�@�L6��Gle�؃X�sh7�*�%]��#q�����f��mP��P��E�Q�J���[2��,y����/p���Ī��
p�t3v�X����6sM�:�̩��_aTlk��M��&2�V/����tl�{g廽F��q�W��C ���t�E�Һ�2�:j���l�gF�vuR��"��&�"G���Ԯ���o.�~�K5[ZɌSݺm�GnB.�)U��Ecn�]��`i�Z�cp���x�=�W����K�h���nU.�V�Mx��ֶI�ӷw1t�/+&�xZ�uGV��������I�wf��塻��	����ע�UP�wUb��dR(�d�qe�����'�t7c&(n��Y���ڮ�EV��c��Pd�V�]�i#��Pڳv��T��Ы����m��؟=c��u<��Lc2��Z.�h�U�̱NkX4�T����Bvn=r)vȈ�IҨdؔj���m�O�0�Pd!B �$�� ,BH
, �HAE$�
I � �RE��BH,(II$X@��$P		 ,!�$XR@�!�@"�
"�I @X�HPd$Y$Ad$�$!	$P Bd$ ,��B
H��(Aa$�$!E�,��H) �A@� I$�HB,�B ��	 �P
(B
I�HB �B,$BI	 � ��)	 �	$�,�Y$Y Y$XABBH�!$�Y �AdY$I Y$��� �E	"��� �"��)	 ��"����@$$?���	'����׿�?s�q�i�6��_�呺UnĎ�V���o��XFe:U��kҮ���F�8�tB�y�����m�E�W�3r��G4ZSv��]�޼����Q��\�lo�$��0�9_4�����u�ۆ�5Y�WX�Ӆ�EM��9f�|r���v�P�t̬�����ҏ%H0b���ʩ��(>��G粍��֔d�ܾb��
��v�9V̙F��q�
<�T_.\�,�K���es8�g$:�]{k��ZW�-����M�[��e��vJTE����/F�:��N�;9�����;����'���ǭ���w�'	mu.5�Ue���|�[��K�]��i��΋���f.{�I�n:�y��yq��d
+9G.�r��x�-�:���3|�cG3t�xl=�\��t�y�fR[�Q݅��uuלvff�H�����qft��y��>�+�3T�Q���	����9,֚t�K��;�ܺ��}2��P!<��}�0ϴ�sS6��&;���2�^˭꿩�_�����(n�0D��%kRd���	��r'����C/b7>��h�4vv�nU��y���Vr�Aۖ�VK��^��U�R5��������0J�n���KmmH��㙒��ӎg�k�A`��Ӓ�+���,kME֤�z��e��=�t)x�B�־���x��3�	{�rs����\&R�;����=!E���q��1e����-X8�|�T.l�fTtqvc�;�=5t��۳�.�T#k��U���XB�����i�W�M]y���W�Ж�����i�u��s�-ffC��F\�ǝ���R�Κ�k�/���[|���n�1[%�����Ht&���^�͵7c�Uļ��~>g���l5�ĺ���,KN{_���}�P��>Å�?S�8�{H;�ޚ�����v�v�ݯ��ӗ7�q����J��T����!]�-	��0����m��լ�d�J�[��=��/LfvV�Չ��)��h�Xi^f�̎Ȏ�X�o�T�=R��c�:�QV2��b�)ңug-`a[n�[���B��I����[%,�������3�J�Q�V���{H8,ؼ��.P��et���8t:D��f�[wFS�v[���ú� �5��ŋ�?W]UJy"���gr��3\޷�l���I��5���9�CP`�T�9��:׹x�^�>��,N^� �x�E0+i������mǛDt����,�Z�j��e^���$��Q��W�ۜ�f����%�'�ί�!�6�f���!�t�3�V�q�ϔ�Q���[��iDvRݣˑ��/�kU��K�(�<2(�4��%A��[��=-�hd��Ǽathz���<Ӗft�O�.��V���NT�:�Y��>�0j졋㺳\3%y\����f�E��5z�É�&�V��x�[�`k�]��-�����Y��+4��60]v32lA�eVm�Fȵ�VB������6n��;6I�Y�V��)����x���Z�y/�9K�2�F�2ƶ���׌��0Ҡ��gM�՜z�}UѴ����ԃ���%q=}9]v-���T8󎳐�cO��N��i]�"B���<̤�ٷ#4����n��Pc'�9�wӫ�A��ʺ)�̘jb����RT�/pP��n$֥0��f��ea̻���Vc����t,Vh�&�:�LJ��ͽd��O;*�;�[��A��u�U��%�
�d�;��	i�F�\���Yo���=uy�ƻ)w������4��H��i���f�,KP��r�[Pŉ]�t�C�^���w��Ȫ�		�Ʊf��	\u�k���õ��$�6��C��X'�t��ڻ,?(�n^��z��^:�T�t�{~��� M�ʵoY�ͽ+jR��)᫄��Y��c�Zbv֛c�I����uD`��1����*��I�Z�L����77+�;tɵ�'�t�Cq�n�BR���m*ܷ�%��|��Yu/���V�7i��֜tu�/�Ƭ#ִc��d�Ӹ�f3�Z�}�TMb�����מiʩ2p�S��	��d�9J��_$:�473]N�c�wr��g�ڝ���*����	V���t�L���_R�ӓ;���Y��5m�r/�}�3��8O��d�8%�ݒ��d#�\魾-�%��>Ui��u�8v^��<�+qMN=�yG���˜ݣQ�=�knQ�B�x�ۢ/�w^԰��FgedՐ[���G,|^9�J�62L�&���ŜWW6�H��!J�!�������+l�f5����q�v5�[��V���Re淬��o��>��9�k2��z����\�ˋ���l]�8ԝl�&�P�y*��2��tX�1�g<pV7D�7�����r��	J����-qoG�{S���P� o+��j	�Y�<�k|��ݻX��@��o���qX��}y'�CԜXObUw�{�Tch�o�R��-�R��%_Tʤ��Ow��ͣ����-�H��c��oG^J�V%�A�d�{��XJV��g/��ݛ۰Y���:��d���tty�"X�����*�t�u�/q�v
�3�Kn�$��������q�"9�i�z���(˺�T��YT	{v�U�-5f3}A]P�1��-����b�V8f-��ف�b��(Nݕ*�#��"��=�9D�!�0o&�zt�%ߙ(�����ߜ�x3~�j���3Ϣ��Gd��4��Ƒ*u勜��3Q��ۜq�#��S�LHA���y�;7���Y�2�ʶ޼Y�F�^��z�k�U���|�6.�Q�7���Y��:��1���*�{���NQ�o.=�ɛX����Y�q	u�)Nԉ���g��N*�i��᧍H�!R�갓�S��|��g(3�����k(�-�LBJo]��������;B�,���Bd��ZUe��6�W,`�eav���.Ǫ���ݵН-Q�ԩBw#��+��0�s;�2�;�{�c��5t����r�]��������b`y$�9�4M��ݓ��b�*��թ5�~d�s�����9t�e4�`RXC���9Ρ�L��:��n�+z���
����0Y{��.�f��ӄ���4��˳%�6������H�8%�)�ʣ����G2=�;�f�{�-e����m�Cf.f�U\{������lnu��[��s��Ƒ�Y��uTOށ�^��HZ��Jfd��4��+�em]�ڰmWp`�p,2Uضu_�#1U&�b��j�<�.�[�4�eX�$�/ig*�y�u��+fusF�l��y��Z;f�5���A��	:떽�Ѯs��q�צ���ܾ����z���2�iu�Տk�p�*����Ts���WNU�Zño���*:�Z�)jU����M*�J�5�y7�k��wY����-r������<�6��LᭉϤ-�{��\�\8��'&���u��GL����+,αmV��[Vz�L�i��:T��Y`Pڎ�3�AK���G��^���B��x�Wi\��
�i�h�սz�;s76�s��g䇘����xq��jƻ5��y�2�)D��;V��G�vo"���r�+�-^��j���BÐ�XNUڡ#��$nh�ݪ�ՏK��:ż���y��x{S4��I=�
Lsxdy���4�o����!����6���LZ=��T����-��H׍��)r�*���'���:פ+�f��Ù;>��bUK��VR�<�ZTF����i����.�۠�q�˳���B�LUt�暫U1pf���%�5W+9���6h�0n�BҖ�JIrj��@�h��\qJ;b�;{�Y0R��LX04�����q�*�R9K�v��N��MM��u<�8�Jw�fM��7]k���[Uxe�5h�H�kk�69��yf6+�v�y��>K�^^.]/DwUY��P:��K*v1L���7�4Q�fȲ�����n�X�Vw!��]d�1%��t7wz���*iT�/۽�V�n��DTo��W���Շr��u��&[�磀��������ͫ�Y�����e�e��[�
��Y�ώ�`��#��ϝ��s4Q����ׯ�p�� ��#������8��D=�#V��o�]v޶5]h�5�룚f᚞�<�C������1�pT�!0m|�6��U)W�y��R���m�ai��d��x�2�If���ً��<�^�p�,����`��P�N,���C4!&�]GL4z��(�`�T�Uu��7���y>���e':6#�X�󲳞�by���]}S0�F��=�a�9��D\Rۗ}��3n+��kR�L�
����s-���,�ʛ{UU�C�O/[Y#��%��]z�3^��N;G(Ğ߫sg����N�Π���b�\,p��[�Ū3�x��0����r�kY�wj���\�n�
��2��4���B]��(rD��]��ԭN�1����w�rj8a;p�6^،�&��3w�믚��7���4_N1E�-Au0�s�YW��]��т��`�b�A˝ܑ�&w�{��xw*�U[X��g)��z��Y�fխ��ơ��O_0�د���ym>;ϰ�*��ߪwlx�(�P%�FZ�����zle�1���߁w3,`IO4����3�m'�瞵f����ۈ�;PB�W&��OjR����seH���`×}z*�H�Q`����s�|n��r��O��K���Zז��Χ��+�y���:��Xm��֬]VV+�G+��A��k��v�eZ/4���� �t�T�'5#��w�I����7v�]�x�+����t5ᢌ4��r��P;>�꠵�eԼ^�pa�j��2��Һ�n+C��z�u�e��-!��̊�����	Uh�U�fQU�TR��)�Ӗe:J_])Iz�c�U�s׸4����ȭ-o��p={6W켨�;�88�뫜���":õ;�_3n�h���N-�+m�	��2���=f�|Ek��o0��=爕wK�Ո��<k�ғ[��|Utx�c�֝]��%�:�.�D�ӄ9�����\�"����A<k)o�QPXT�YUy�<���T(�L��]�"�	�5N���̊����ۆ-B��9v�y�~�'.�q]L�k-ٹ&T���m�n�^�G7t�땳r��L���Eu�Ӄ;
�ʣp?P��/���ad�o33,4�w��T.���8hWq�k�M���yv��&��3yVZ�f|��X��D�kY�$W�n��d�`��7׃"*��5ʼ���Հ���A�Vs�*z3�j�����m-s.�ް�UVV�����C��@�%5�(��c¸�K�f�2��<cn��ŉ\xfM�}2a�^^�͹��kyS�VU�ϋ��fe��Q;�9�,_�����b�{2�h��M|�+�yR��T'Wi��qn��m�p�Ͱn�4�1Wcۼ���V-!I�q�x}Y��mn��H�sq�[�$����Z�
zs��>\혴hk��͡;"z���a�cQm�`�B���l���(��꼡�R��3�t������Pu�B�pSv���LX挛|�i��:L:w:|i�V���mvmc��M+�I��e�z��e��ɱ%�EE����1���p��C�򣜗M9�.Q�}�vu�S7k�!y��7}�e�0T�L*N�狐瘿&�M9�4����x�g�n�f�oɧ0�ov::G�{)S��K���s�`,ztz�䧍�e�!΁�&�����(��p��:���MT�,��ol���Du�|�-��w��5x����k(��T"�& p�����Ն�Ap�v�-TK�q���ڕjb��V�ek�5���澬�w羃3w5(V�yX���=���=[T�Ov�֭��D��B�:��ͮ����dƒ2�v]�Y��3j�ͼy�F,��F�+8Ǡ�9�/��t�w��n6(�Un{�*��	���n5g�ZXMe��LQ\v[P����Ç��R�t�5ׯ2���o�~1�Z*Y��9�wd�������������yo�ڝ�X�#�*yԃ�u�e����hO+c!�0��Y�I�tq��!?us豝��h�&(P�*������B���ZM^�8�}���]���мu��V�����<��Ƌ娡��]���
�x+���M��3M�G���\:�|�U��n��<����훮�)V:[��e��l3%Zvh���9wX�r^i����:�\���.|\e����X���9KHu�\�;����֝��(n�.�խn�r�Ҿ�2i���x�kYYV�pr��H�dZ�(u�}�g����[�U���Y�y��.���{����|0\��d����iPԻ�ʙ ��P=i�W��˘�F��3�|�y�S�y�A3[�v���S�֪�GZ��SU*`��.��l�2�G����NEx��GR��L���ڡ:DWI��֋�2b"Lµ��)�V���Y>��pb�W�"v���85Y1�u�.s	����A��MǓ�E�5f�ӗk�*1%�8���ܼ� ���I����Y2�fN���0i=�y˩�O9�����a!{�Պg!&Z�c�I	�:�q�j��a5t%�7o�����n��\^2�f��ǫl��,HJ+ɚ��:,�Ѹ7v��΃��ɥa��z7ԦF�HST�X�]�+T�P{(c��ݳ���v�-��C50��+u�j­--�=Y�wx��-P�=��j�^8'����Q��Ñu����Uf:��L��=��v4d����X>�PV�1����҂Gzu��m�0{��Z��[���*MV僎P�W�s��u�Nu�li�ކ��1%^Ô^A,dÎ��5���v�$��\���j7C
���R&�����<��o|���l`�G�mc����9+${w�8E^-4CT�����^a:�����Lжi�ƥ]ATw�u�۪pʻ��rBB�� 1�0GK �ZpB��x[ᰖ�6�\ob�����3�:��*y���U�o2ܼg[iu�d�M�KK֔4e	�-�v��%cGZm���YJ��� �l��B2��*�T0q��Ы�	\��"�7� ����ܖ,�h���n`Svu�ۄWdOdFpWO����vE��=Sۭ����Nt����5<�8����r���Y�r�PE����P�-�y�mÅćm��e�ʙs�z��;����*��q����	Qc�6צ&;��;,��7.%�n�S�.y0��bgJ��ݭ��Hb�n%,k �F����֕�`�&Zqc��o'sZݍq</B��r��[�����YmO�{I[�/ZVնY�`�Yl�Cj�2� b31]q�[�n�;E���vƷj���eە1C�9���Ci���LK!k6&
ةe7k���Pv�w��NS�Pݮ ��zD������x�Z��g��M���m���ۉ�:� F-��d�n�G�/ �s��<h����UD%�m��ͭ���M��ͩƺgY��"��e�%�KfƖ��aH@��K[É��X-%�u[�t75�ԅ6�z�(Ń�q'R�Yv����Y�H��Qn2lȔ[
��G����5�[�'G��[E�ւ�B<��-���;E�v����n@m�{-�뛀�v�u�[d*��(�]]s�k(�kN�7`�^_k��]�Y�z��!�>1�x�yr�՟:�0�p���
�4�#YL�h,6��$llk��١�.��L�lqF�N�M�Z��\��)Քxs/�*�h�em+��e����3g��PXR˶�lAͯ(X��nq����nIWD��;1"���qfyޥ;�{��su���!�j�,�+2U���utRnH�i�;\�ť#)Mf���fb��M4ѱ�5ko�7m������771��܂�y��n��虨��fSd���x��'^%T���vB2�2j��5a�����pn��C����CQϓ�p&uo&Cn�RM��(��).��������qձ]�;���=�y�W��@�֫A�ö�c��B�ce-��v��]�˥1�q`ܕ��s��GJ�R�L6Zc7Jd�ݰ� &f����8Ɯ	��$)D=����qR�vjJ6c%�2��{g
%�;S3�;����'\�}��D�g����k�����0[۞:?_/}�������پ�㠱��.�ĆPv��۩�yɂ$4��vz�'m�ܑ�u�盌t�.qXgG4�Wkp���sۭ�*N��$`�W<f�z��N[sj�r�6�˱Gi��Cme��q!�⎰�p�+��Q�Y�v���R[�p#�w��;l����z#�պ��D&�"2�BĎ�ޞ:oi/��n̺]i.
R0�&*�+��&�C5���dh;RS�W��u>���Ɛ+��^ٹy�˹��Qf��N�!n�wn��M:n�F��ۈW�u�W��C��7(�\S��.�YK��d�መ�/��,pJ�&�]�TRX^H�����$�U�KS���u���#�Bfj�t,��O$%����Ii�1n;GE��%���&*�9�TF���l�s�hz�L;�uR�=�V0p�5*���{-c��/�\�$�ܐWfx�Ҽ���N�6�,
ְl�Fڬl�T��Wv���C,I��u�g�G10l6��SQ�����sn���Y��YH 32��8.�#f�!٫=�o�wa9�-�8�=�Bvw[��z`��O3�Ƴ�W8â�,S��b�%b�&�ݼ]��(��C��X��y�v-�+�包yظ14󋁰�溵k����"�b����Xl���Ը�Rc�r�랷�x1ΗS�ޥ։��*P�`�\����j2�׻[��On��k���tE�����8mQ�z����R�ڲ�aۭ'���B������-w�む�iz�m��ͣ;�gl)�7d����������ǜk����.�,��ӼՍ�r�&8��l,�/PM�%�pMfe�<;�ֻk]eZ�۞e��k�[�NP�"DG2牮]���`4�%DeY���M���rJWP�-%��͈c(��c.]2ξ�f ��g����ѵ�草�m��<������7�m��`w[��D�Z�r��FS�z�~ܿ	��?5�jn��7`1�Rn#��5��������A���ސ�v.{�D�7���]��{k��:�8JHG����zs���0k�CP�XR�F��B��%a��0P/"KR�2B�7�����7`�ж�а��a�,��]Ij෫5,�)P�jƹD��W>	� �s���g<�nmķ#.����Kz^�͝Vj�m����fЖ4u��RQ�ob0�ͦ:���w���)�ɤ�ۅ��'*g�:�<��*�pB��A�L��yv����lA��f�^�+��%��Yl����`�;�eL����͔n�=fY툜��uiCs���-Qܦ��	z0cs!F�\[�ׂD�����3د���I��o$ct.F
]�ϗ[|3-3R��֕!�n�bfE�	��\p���]�:f3v�
ۑkF����;$!���i.��H��l���m���UN��W��GL�0�v7�1���<1uQq��[.��3��KPQ�6�����B�u�c�s���nWW\uk�:�x�&�1s�Ҵ5%�F<Tﺾ���b9C��Ζ{��=�>����m��{QM2[�Bn�1^��q6�&b[��-+���l�Kk۬^`M��t�8�����v�.^�E�N�׎�:�˥�#c�;k���sۭr ܻ�y�=n�#us�o��!�B�(�Kf�P7&�b#l���#և���u���/7�-5�[%�V���5�yێ�����5c��E��j��a��j�`�6�&G9Q��r���ۡ�F��i7Mָ->]�\[���l#��C���Ź��e�l�A٩}A��;#V��K6��03Ռtz#D,�3�j����ve��[��I�pj��Y�q=��{Z�+<=��xW`��s�ky��j��L=�:.qF�hv���J���`�G�M���-�h�@�^N�����˭�
a0���l:��0�e���L���K��+Qfg���n�'Wk-���a��If�� z�Y�snm�l�շj�<
���3�"���.��eڃ�ΌX�7/Uqϙ�	�E����F�Z�A<4��Έm�H�zŮ��@�7ƜU��D��۔�; R0�۝v�+�89^#%���U��x!-J��剰4�F�Q
ڄ��qq1+�T��h�;�,]0�"�59჉����Mm�H�JF끴4*�	[m�7��'ly*��;�t�u���	8ݎ����)��g!�7	^�1��6rLR"Y�;�K�+W�����μ�v �����T�'5��s��(��SP"h5�I��6���dA�kR�g�k�3��'���g���ug�WA������)`�+1�c�k]�m踷Vے�(&e�棡�Â��%��.�jU�u�1�K�D����)
kLlAu�j�26��ڇ��]]+ۇ[��{jL�V�ne�aaf%ù �����s���Y�-&��F��YG�u���d1L��X3+`2�,�L��d9==b3�3��wD��弗]O\Rc�p���%��ae�`�s�)m�32h`ݹt�{iK��^Y��G���NGnٻb�M5Q8�p�B�č�<��j%����y�����XI�l�|]k�p;�4�����X�Ӻ���ed���ۛ�B�㖲���e������g�.;*�=� f�W^���һr�q��Z�ˇ�.��,ngqW�<�^�n��e��,a�(XU�s�3B2��i������ٝ�ضtŖ��n��/2s[�-4��ۀ��n+�ۧn�7q��X���0�n����s��:̹������4G� �X�jW]/�Gh0i�:�x����׮g��F�+ў�1[���9��}��H=]��:%T ��.�:�����jV��,͹���e��|�H <&�r��x�!����w<M�C�8m�\�JB��.s�s�v���Nδ#���&#S�����҈��,��8��GM:f�cb6��ţ �P�M����J�f����v�t�����b�=R�i:JlA�%LI�b��5f���X�n���n���+8��i��m���M�H�i�M�s��敩��3Rbit.&�@&����j�9ܼ��g�ι��a�Ӻ�.'��>�:��H��h�#�	u)��gPݸ�.P��4�� pÙ�=u���["I�!F4ˢX�
+`��Q���`D��m���s�� ^8Ę��U���ΐh��=h�1�����n��Ȍ���V�%�	
V�P��ł�vw��g#V1m�*�R����\�S�N��9��qq�[-j���1��8g]�S獫Y۝�c+N�A�=g���{6޹.xa�]�x8�R�u�[�^���q�6
{D*:�lp�l����g�+n����_�����/F*����+Z^�hH$�c[	��B���Sj7\�����
M��]�۞�s�V;Yu�<RՌS�@���i:f���*ې�p�ٙe-�H����
\`�!)�4�V��$�ZX1�i�Z�GE�8<ݽ��箃Ӿ��!��lՓ\�2M�Df@�Y��[1cr>.8�2�����P�������CdY���4Y�JYl�cK�5��\vH���h��p=V��p6��d(��׫m�<��K��[)x��M��cN�:{Z�u�\v_o\὚�-hq��=����:��8é�u�:�kpm�^p���;���り��Ȏx�Ͳ 袒J""��3��,miZܲ�H:8�mEBtq9�AHvnAD!ppt�gi�չS����mvt〜SKt@q�v6�"��p�")�p�Vd)��RJq%����L�gb	(6��:p�L�D�$@Λ+l��:���+:'̋�)���Ef�:RttQ�9Ip�Ͳ.$���$�mdYi:uQ$8���gFq�Yg�TAr]�Rt�%J"8T]�ICk;�m[i.�*t����ĕ	N�fqj�.����ת��Za�&�B v�l΋!f���)��8�Bj�-�m&�Ҏ�I�ka�b��V٭��q��'�.nw/$�t��o1jbRj��W�cf,,JeWP�
S����H�+�C�y���h�k��ۄF�5=\�!��v2�;�;m84�F�7nv12i�Jm��\�s$�[�������[JN�\c��rcm�I�����7EӷN�˺Ŧ$���T�3\�ݐа1��	(�r���Y�is��7��K��Zh^�^a�kR�$ev�pV[��<������i�	�J�u�����/�y��|i5�C�քۍ��K���Ł5�l��Rz����B=���6K5ĨH����b)���Ѷ�Y������m�Y�V��Si���rQyp�7\�XUR�1F4BƃG�bRU��cX��xu�F
��G���T�c��ꎸj�omvv^(�]��N圈�!ݞ*c����-�M�g^�葪���\n#�ˁ��Q��h�+���S�ǷL�;0��qv8b%�ly����1�6�1�]�%��L\���cq���#��v��
,p�ZjMs��E�VaoG�����֋[��] 62B�a�p�,oi��������:h�	�#f���a�θQ�q��Xx��i����>5N}�5��麱u&�i���*üg�P��\s�oDm��N�Ɨayn_B�xm�#ņ[�^3��wT[{vp!nt*��y�lX�2��]��x5qy�,E�L��u����8���m]�fsn�<ٌ��;�(��N��n�8�׬�Jr�֗5�x���r�vO��ѫm�5ͅ��̝�{�z1b��\�%��5�I�sku���c��D�Ҵ��D�iH��X�\�:$���j�F�� �K�0��ʽln�д9n�n�W��Ѭ]��-�,�
]s���T5��c���<��yNNq퓸��+K-AA�X� ��Ӛ�1cR�e�I�b�J,J��F�����($ h��m��޴�R�b� �YKc��<�ǃaUZ�:ӫ-�R�U[B �`6[k[,���Rť���+e�JU�����)>�?�4���mZز�懭��-��jBi��i֖Q�շu�����X���7�Ѥ��"�Ts'�C�%m�ƣ���g���^ �a�,��[�C-@��Bȧy)b�w&�|���:�Wq���jgT����A�X��n��Ւ.wy�u���~�~?wR!�B-�	�^\��]x���s�[�+�M���7��9څ�PE�~A�`7A����1��5֎��u�#� �~y�z�5��˱��ׁ��Ol��䯬Υ�?7_6��2��	�)�cG���Y�}��]��<pu"���������euT����	��uv���ұ��������2�)*�k��X��^f�ZM�:�-go��w�|~�_6��[��a~ʭ��׸�\�޺	�\�@������ #�~mؿ�m Hn���Ʒ�����otf�eoygv�JBG9�j�d��R��X0�ۜ=_09��j�Z3�����ksE8kG�"u�1�V��A�wkJIS=[���}�� 쯛k�p�[�؝��?v��8�F�u2���n[�oO�!���i��з��=��?wK��|An�-�d^L��L�i�Nuv5`��n�p�8����׸��޾@��@;��Ol�|�-���|A%����!��!���܇�X�h�^̛�z��ҒW���~� ��m� �[]ޮ��-��PI��P��UV�(X��PF]�'$��@���,tحB�ԉ]5b!�|����耹D7_/�v,�w{�^A��3�Tз�SV���t�Oo��A�ز' �n�-�`�t�#�I�״�U�}ϗ�vS�g��:����~s�]��s����Cu�I�����zł9��"u"mز_/�n�GE]��huA{���)�"=�.�1�g	-
��b�y����U��ˍVpy������/pU��V�켈�g��ơ�_7�ЂMiI+��|�A�R[j���/�͠��w����Z���A�H�۱���/&z�uJ�P�3�t�O���A�dK�w� [k��D�[h��{����yV�]�0�R���?9��q�����!��B)龃ʳ+�#.Wƪ�)+ �iq�8);/^s�TN��@��� Y��Inc�_�c/B7)Gb�!��
�9!�wkU���1�Њ;���i�A�B��U�A�G�����Q�]�W�0��K�A��gc� ��{+��w��� �:X�n\�v�������yA�X�"�B-�`��n��Û�Bs�V:��	�&�O�xY�8�B�w �,��mذCt*�=�gP��:A�ő��,�o7�>B�iHc�jW���TC{++ȯ�˧苽#�x�U`�r�5����]u��/�&���o�͞��k+.����y�S��ܔ�6�2V=g �\�h齯��������-N�~���5��Hk����@���^��+���,�̃޹���C��A�,X!��:dq̡&�zU����ڧ�,��v]z�Hb��5�&f[�p-����ue+ �
�
5^PO�"���}�uPދ:��y�;�{�,߂�t{[��+4FrAz���Cn��Ch K,�=����!��_CC�8<��Ґܞ:���̤�͵���mX����	}�Y��W�۰��*����ՅNf�4_��rC0e���(�Km/�t�͵�9�1�s��n� C:B;����W���Sپ�~s�#���,�5;�Ug��y��<||Q;�_�7A�+�m���w+�����ő��t|<��Ґܞ:�	̤�@���A �GȦ��Ϊ�j;�r�:�,��]J�Z8��2�+��k�ަ��*�>�l܋���X��;��Ĵ]��Wϳ�4Fn�ij�yo��	��_���E���������'�z�0�\��Sj�\E���YJ]jMu�۴�����U:��As^�7\u�͋m�s�nqt�w[��T 1.�u�m�{,O\n{q`�s�t�,�!yF�՘���P�8[R��]ӄ�&����j�J�;J,���k,�n�WK�]	]�X�\��0�:��[vu;yf�4���տ=O�"��],ک���p8�b��MǕ+e3��h��V�-�{#�
�2��W�-���5�}h Ye�B��c�+2#w<s��2���p\�1w���`��|C�B�ڰA��{���<���{yX ��@y����M��]�9���Nv�.r����/,�X�vu�{@�,�A��_L�Q�������� sZR��Rޮ���͵���"j�'~_�z��B�<�F(�۱gY����s�:�/���@�s���Էי~�=�}��E��~-���!|[izu��{n�m=ԅ���Tѝ���0Y��~9ڀ�9|�>݋".+����{(z�;��xk�³�*��ϖoe��nz΍c����m4k����Y���_?��ϟ_L�<��py	Ǜ�!�<u/��:�{u�)�~��{��?7H�Y�[hY��*5cԮ��F���fp��|ì�_	Y��,=8��A�SC��v�$�UkxY�l�N����7���Ükڨ�L8���J �'_��c��Tſ�#��!�b��\��wq��V��Ed��D韛k R��J�9}��¥j�k��v7¾���YenŐ�
��/ǽ�e�����#3lY���L�=ܐz�����O��A̤�m;�ꮿ_����A�K�j�m�dA�0`:Ɗ�]س4�=1&.x�	��|p�nX����e���@�z�Y��l� {Z/n;J�
]a���h���ך�V��Q,!B���O:�}�@���[��ʏ�i�}�/?l�f�P�K��Y&�$,���Ǌ ��Y��,��!��d�;X����}*��ݐe���\��Ƶp �e  mBm�X�osY����q
��Yg����i{���=#�Zq�5�nq�2Iw5R�UwR���z���:�����JA��E�+�M�9(q�&���"���%%�5�,���y����U�y��#� ~>8QG,X!��:g���&�3�/�:]}֐��_X-�����Ӈ�/[ف��B�!߻˱][�?d��@�Y@��Cy��_�ηO�U�ft���G'�+�Ƶp?{)�P�[j�%�Yi���K�n۵wيO�¯])qns��&x(Z�}km�7�]XD�!"�bͅJ��Ú(s���Y���w�c��cC��1��>�%��� ���Y��鐋mX?7H<��畨B{U�A�HzLؼ6��z�מ���s�:�e��p��XA�b^]��C>,�DnŐ�_L���m^��oo��j	$ˋ�{i/��+�6��Ղź��B��۹�H�f�}����P_a@[w�zew��k%���2��,ᯈg�Z�d}w�n�>�{��d+^R�R�W��%�h:$�m��U����l��x+^IZ����|8�Ѫ�lx�(W�r����Ku���?6Ӓj~whU֌�����k�o��6��`G�阇|A�_YDn���ưY��:<.�&�����5̠����n�u4.��a!�P���Bŏ����}�(�#�`����L���d\xt�./I��.2!ZqʄZ~���t�!�B���v���a����:ŇOz���Ӑ�{88Ǘ	�¾%��vG�n�J���� w5}fJ�L�[h�T��=�ߕ+��^�3w�>���P�A�rY@�nŐ�>�$Yc8���zŀC��L��o�%�	$Y/�f�_q�R#��%L����G<��̶(�B��
N��n9�Q�U�c>���dԺύk�׳��yp@���KCi|]24�m�R�����|��<��~��{:Q璴$ ��`kB��z=��ܼ�]=s���4	�m�R�/r������f��,z�[׉
��Q�eS�_���)�j6j@�Pκ�+�K��ٌ=�c �ͭ!)4��J\��l:�=��V��SF�t^�NWu�ق�4�CAű��bf1����A��p����.��ىm�����n�*����Л��Cūq��4�U;z�^Nݸ�wQQh�we�/\�}t�ŏo��{s)f9�=���9�ۤ��;�Rl]6��j��qGk�����Ag�̽�l7` �t��F�0��2hӘ�R�lF�d�p��(�j�'�_!�_ڰA-���طI�X�ߞ������q�*�7�'P_x��!�`7��(���f=�F4�2�<��b\xt�d�9�R� �)F�!|[k�_^h����^��H���z�>mYe�B�R�T��}�e���׳��yr?/��x�.�ڰFw+�lVb+�H2��#Y��y���9'mc7og`��ϲ���%*�]���qgƁy!�����(n�n��>�폔_`��
���.���"��9�R�A�K�ڄ [j� ����]��u���v�]�D=Z�)����Tu�=\�X�<Y6�8��TU!V�w�b4,�� ��Xt��|k\��c˂��x�u�9�x�<A��X�A|@t�_����T�K3�9�b�����6������|��"S�3#��%8�ٗh�w�����w���=P����s�7�zH�X�*@�h[�y�ClŘ�i�ޯ��^��͝����فu}��Yr��",��'���XMA}��۱`����d{ؼ;WwvQ��O���q�S���{�eW� �_C�{��W��H�Z�&�>��8{ۜ�����A<Q6�[��7�Ẓ���\��r�=�a�uX��x�m}`�HC�B��Ҿ�sү���j�]!�&�z{fuc*��������jD��� ��yeM� ��UUj���\b5�ƺg��my��Gڀ��{\0�ۮ����F�P�a���X!�̲����'�V���~s��t��x.�>�o�D�B9�� C-@�m"�(�~���gO�%�dg�ߍf�+���<�|p�r�nޚ�����
e�_����P��L�[j��T שuֶ�2v���)i�kl�/e�/J�7)��_L�vq��i)���3'��������$.�څ�^�X�=˳3RcE�:�	Ia�-9l��y�f�u�;��ٮF�+�tK6�2�ɑW\�3ⳍ̷�T�R�gR��.��foP���E��X�m:�In-.��tr��06gV�챘ثKx�o�yrӋ�(fX��U.�7�=a�Ǚ�{J�f���ss)�	t����fؙPig3u�%�[w��^L_#%�T��t��v�ٚ��l�t%ԥ]�)���w�ҫ���$���b�Ԣ�k:�Ѭg�m�8++�V��Ն���S��F�W����}��8����w�}L���Z�}�>������L�+1�[6�B�K\6z�K������;t*3�-.��T4e#�}af��n2�l���l�X�_�,Cb�	���0#=��d�hmy��S}�Wb,�1���.]O��ng�3�{K�^�Z��^���=���n�"����l�e�B,V���n� ���U�^U0�2�0۔w
�1H�[Ɏټ���J�%\��vw[�ʷM�͒�e�
�NW�Ιq����׺�"��]Y����gh��g����,�����ɲ�������n=�FV8՗�a��W�=Y�^X߷1�IZ��K$My��s�<�G�V�Y\m�NӢ��Pх4��:&�,���9�t�PcyQ~�bJ9
�=m^�X��i[xu-7o/0��4��h�gvح�ʈYX�`2K����{���*3�e?��].��N��}�~�:F""��L�P:�wv�v�mqև9A�q�E��pT���
��m��:����m��q	u%�	ӜHT�Q��p,�&sZ(����;K�.8��".�
8$(�e�rV]�B=��(�k���h�D�"�EY���!�s���6隠�U��WGGp]��;������k͝��NY��.������Q��ZQq�qݝgvu��3��Y���݅'e�u�ź:�����✩:�v'u�ArY��7whT�pS�@�	5_�V6k�^e^=��P �j��,�� �݋ ��
�)6WkO�,C������Bsd���{zJ�~s��e"Y2N�����b�.R!���B�n��f�Wh���G�A����
��PW���yp|p������L��}�7���P��6���n�r��ɫ���U���mzY��]E�P�����:_F�mg���|-�l�6gW�V�f�p �W�Jgz�߈#܂=�6��[��y�u�Ϧ�{A�4�������޹2x�N��K� �e|�ؾ@�ԩ�&N�;���Dy���вh/�t݆��K3���)x�b���ʇ|}��b����6�E���C�'j�WZA9|�}���|��g�LٝXʷ�0_��';P� cϔ��μ��8a�uy�f�r�*Բ��Я�4+���x��F5�`\���c5�yd��1�.��Z�Wp-������<�{��X!���~mذCd~g���+#�W���5�[<�����B>4Fj�����a�}��*+��YɌI�فhPz��7vcj)V����p��&�u���E�*�!�?� �@X|���v/���U3�Mg���Y�s�ܤ|;��� _7_/�mY��"+]�����y%N}�|��\��a���:����0_���j�r�y�({:������ő΂J�۱`��_���<�޿)�5���^��N��K�����b�ڰA��_7@,�g-��#5}���6�[峁�X~u<�89�절�S/3=)��{ ǋ��-�g����� [kO�"��W�4�zwq��ǝ��[ݘ/���s9� �z�wv��.���_�����V��V)�Ƚ�֖��~���}F�(���U��^Jk(\���Aԡ{���ɦ��im5(f�|��]N}��}��#�Vϴ���iaa��Hg� �pS���$i�!��f�k�wl�o�<sq�q���;6����)-\���4�4e��D�ES�w�8.9��vج�mcrZ��*"k�p��;X&:�ع�ϗK�m��᪗�)\sGI��a5#����ή�f���8�W7W�@�a���ٓ��k�潛���a�q�2��Ҿ���h~�����3�����v6�Rm��c���,.�qTBA@���P@�;zŐ����nd����_��Z���:x�E]{��͏�� ��|�.5��[�Cu�-�,���E�k�:6��8i��@��|���z���[��5r�절#d��U@��~����+?G_ 鐋mY��{��5��GCQo�{��u?y>[�������}���YrY@�v/�K��3Ջ�H�߈?�A|C�B�ds%�;m��0֮ ��@a�Z�[����6��gR �Y���k�Y��({���P�X�&.c<�Z��d|(���b����L�ד�>[��ޟ�+�d9�2��c:2��*1I�f\�đ���\��2jS����|�"�Ŷ�Kt��J�TǞ�ҷ�0Y��G�ie<�uC�b�؂�? ۱`�Yd�������>K����X���]���lo�t*��h+}��ٜ�n�ͅk��wӇt��o>V�'�gY�%�ڮGx�����UP~#:�A�#]�ޘ�a����0֯��R �P�mu������wX(� F�T	�!`�AY_Cn�G�w�U"�M��U��e۳�̃o� ��_vK��|C�B-�`��� �`�J�_p^!|ج~-�q��܋&g&��s�p�A��,�[v`��o�������v,�_2�ʹ0��߫��_ґYs�����Cz��j�A��R!�Bwk�u-��Uj�L����GdBn&�xܕ��6�U�EV�5��� $K�t�6����h�YeCn������y�w��m�0eݜ�3�,��L�L�鐇Ŷ�ź@�#���3������� �vS��c2,��Nռs�w�	�rA�r�ϻpl�^��\�X"D ��!�b�m/��G3nfxe+��}���Ռ掵-ކ�')؝�]��l�w5b�fv�줥h;^Nu�$��U����T�ҹY�	2�+N�.#:�u�nx��}��|>�z�z����޹��}��R �� mX ���T7����k�����A�A��b�����;�y�w��m�;6&��{5����Y�t2�c�m� �� At�@��j?;͙c�r��汹)dΧ��9�ϻ����,D�ŖQ6�S�N��%[1����DO���!��M��羑ף�T�e;0w�t�m�S�i*�����~�Ǐ�Έ�|C�Bm��o�����^���w�"�����~�Ud���d[�e�_6���k�/��y�p��g�N��43�)������@� ���9,Y���[B�{Ԥ��*��_Y�� �d [j�%��Y���Og��u6��,����,:�,��6��%N9j���o�^>?`�e�#z�A�!m��w�����f�*W���"����^�GN-l�,��uf�n�������V;�r�	B[,����∨��M0ڵxVe�5-�  |k}O����e\N��B=�l�!�����E.�`?�X�S��ȳl3xl�.�(����?L�{3O�~y���ߏ�>���L7����͢�������sZ�M�\37Zc&ڣf�0����β���D�B���[��}�IȽ3�Z�74#�ަK�e^ɚ��;P@��!��n�Y@�7�������:�O��=}
�|�ι��}��D3_�^�����~�b|W�|��A��d�̳��v;g7'�?[����aSr���E�|Y�>�/�K��B���پ;���l�+�֑���25	n�t��Os�u[��Q~@���`��%�9g����Ʒ�6a܀o>@�Y�6�X!�W����~���ƈ��vtT*Y���sMj�~ܯ��B��Ղ	n�G�u��u�u�4A��z��R&w�������vn�z�K��y
�����o�5�����͕^����v�f�myU����e|@G{���W��uW'Fd����Xmؗvm��p�t�4�jw�~;;d�H͘�L���X:#5�n�� �,��B3G=����S&�S�v96;=c(�ە�<[��Y�����YH�Ĝ�J�r�5yp��]��,�%�]�Np�� n��Lv̇l.�Ȇ����7h ����;�S�C�u�wێƈ��i,G�jſ>~%��ϰ���ҷjCrcڱ��0؅{$	����R/�4Y�RF�ÿ��bC��(Cn�=�/٪���N�A
qr��V3�T��^G��!"�3�m �0A^4���C�F��	n���F��W3�b�k��
�9N��,����xy˕��h27R�|A��b�!�_ZE��V4�nY���n�H-��\5�5��۔��!�W� ���#���7�:�u�A��, ��q��y��0۾n��"����x�lZ������՟��e��k���w}�w�7�j�up�m�V�~�4#�	�rAr��|!�cH4H�Y�>���;F;�� 2��iI� �s�����������t�T�e���b<6#3��I�ܿ��"h7�yj��^z+��F7>;ެXB;���n��+�����}�{<���.T����yo�ݰ��q��9�m�^���Ѥu�:~�G$U}Uôn��ۼw���"�Ix�X����Z����*����G�����M���n_5�dp@�J�܅��u����U|�M|�<�X �Α6�_���n���-S��OZ~��L}<�U�ނ����,D�n�۱d6���E��9CH?<v/�;����k��)BQ�ep�4֮ ��/��MײS�tg��W�)�|�m �-��l%Uu����t��9~���ʷ|֭�E�}�A_u������^�j��^UorUIE��d�.�Cs˘�sk�v�f^��8�qy�k��b�Y�\��A>�D�����t��{-�vf�د����uN��=ΓQX�dN���A|AmزH���ٹ�%y�����/��^��(�2�l�U��?�D9@6�u��N����@��D��@m|�m��}w����o�G�5��7��H-��oe)f��ۆ�21�H��l��P�َ�*����z�쪵V���ஆ�ʶ����������|>�|zn,���ml������rCh/���-���
�P}��߃�_z����[��{-�c��ڗ�sB�p�g!`���w9��y���PD}b�!�%�[v}rh�SB��W��_t��}�8l�U������ڲź������/��S<iA�q���Q��Um���h����CŦ�B��czj��]ữ3߲�DL�=t�,��3g�.�����\x=<=��[�0�;e�NA|Ch���~3���Hb���:��`6���^>�!�w�j_����~��9o�E�z��J��z���`j�n	�ACnł��k���y�0_N@�ψ;ۙQq���i�_p/)���-�Kt�n��ўWld�f"դ!��:�w�w.>��Yb�Ӓ]��PD:u�JI���x�WVe݋���Mz��?b�p.d4��x*I-:qI�(݋��A��9�b�r�b�;�nz?'z]�V˶o<����@�
�|�z�{�,{�ޢ/{R����[���
\���Hz��_q������н\A9���_ ��nƶ}�>����>�[�Gs������)��ʽ�J�C���M�bbͅ�߽�����Y����͂���L�{p�4֮!ݾ��:���̒u"�_"�VA-��׾ �[h`��Akκ7�OΠ��ؿ�w!�g�z��=�$����#�X�C`)��wS�\��;��}�:D����n7w�w�׬�{��R��h^���rA�@�A~mؿ�m)K�7.�tOk�/��	����ɲ[�IU^Ü5�5�� ���ت�L1���95Y��D7H��m�ͯ��[5��>�������޻Xm���j���(�{=�Q;۸��;=����z�0��x��Q��	D�)x���:�vtJ֣W��MO{�\7z�=˒�EV��xcwS�lTX0�}ֆb�XG
�FT���F,f
�5V�ժ¡0g�aa��T'u�8˲x�nZ�Y�ܑ��ۑ�f�ٛ���ڵU�v��{����9��ּ�v�r��y3��Yy�3�8!d7y���wʸvh�������Շ:�!T49���5�k�d(U`vb>.�]�$6�9Z�y��,q8ݓYB���P#�ȯm]�f��/ �Ý��AB��F�o42_Z7`ٶ�[YTP��>.�v���h�Y�����Hú�7O����jG{Ÿ�Tz�$�S����s�J�eP��'w�[��SYvo�v%�v�*fQ��u{Q�r��G>5��u����ux�1��ZvM�ks�l�Y�ev��sn���6ژ�������a1Ֆ�3 6�L�ښ�C��� �36���L����/%(���e�uK�^�X̪���+a,�h�1��$�f�n���O4M��g%k�6V��w�����o#�G���qdk���`���F^P��囕e����o(
m�fƘ�F��Q9�����s^��}{G�.���xַG�L�
�)����v$j��˹�EΙuNZʹg3.�q�F���/W�ߘؠ�5s��9^�[�b�Ê�#d�R�t~�yy5�=U_Nt��Ц���&�:��j�䚫Ӣ�Y���rΖ��hL�촲�8V�ޫNf��f`#��T5��&�n
]�:�=Cr^]�oϊ��G��t*ڋ�
aa��
tG$weg\Q"\A�q�%���9�AQtGtEG\\qu��EQqqE�gY��WEӝ�VugP���GR��ԝ�GP��"8�Î������Vgp��:��H;��Y�wv�"���]�w9t�tTQ�k��˻:� 
��#�"H����4.��Ê*.#�,��-�twE�ݕ�QY]�k���N�(��肣�:�㢅�-�o_vO>���Dӑ�m������N��R����/�f�ۡ�#^K�X)��y�z���M�CѮNє�r8r���l�p�v��K��<y��Wc��8�����H�#�M��s��E�l��i�k�O9�E0h3C���+T��U���M�s�n��w[�-]�U�3b��X��s��Mt
�����q:���v6�梨`t0[HZ��,1;m����]zʄ(y��� ͫS�RԂ(�c]�����SB�]��-�t��h��ݜ���D5"�r��Fv���n��!�قv5�ҘB�T_/)�6A���cvQ�\3,�91�n�mصq0v�h�x�'s� b��3�<O�9�nS�S������u=�On ��{$����;sGX��G=��H�_X���:�nu���u�6�&ݠ���*����Sܻ�%ם���"Թ�l���b^yq�9o.k�Ǟ��A-<�X�l���-Ɖl,��`�v�54�^	GZ�����
hv�\ڹ�t��j<�q4���#<-��`Τ�M
����ŁZa�Kbݐ<��3��f��M6Ԫp`��@��6x*�%W�ے�C��]thi�Y-童rix f�=۵	�0Sp�/n�7�㊂�dء	Z�T�a, e�)qubj �qD��M�qw�4�q�" U��mT#hӦ�m����:��Ņ����h��w'g�a-�>x�-�G�h��T��ĉF�h,S�K��N��ڷY.q�d��;�aC��s�P'��Ht���.���9���r7g�m�7`���î��#�=7^��-�S�׫���\qn'�n��R�vQ��6�v6�cf�;��=�m�k4&�Ѧ2�(��h�5B��6�E�I��>�u��v����3r�b�,g�Pn��F��s���ڛ8V��<o�����CRce���v3�P��&j`wX��ut@;6@ui����%[]�o���p f�n칭�B�0mq��ՠu�6�o�;�N��y���[�pGa�-��!1�S�9�\�,A�L��&��A�I��&m�Z,�d�3F��vxN�����A��VmۛzD%Q�֟V�l].�k01z��)4e�5�C X4�l;�c��}Y)Rha��W�zz��Y�Ov	�ֳEj�p�m�PuP�� ;tn�m����t��VeFT�"&�Ζ�XĤ��k���bc�ϳ��i���N�B[0�J77L8A�&ҋĐ.�u]G%�-5�}�<�|AؾE���� ����a{��~�4/W*r�p�a��swn�П@���P_[v,�����W�Wv�q7�C��}ܾ@k.�H�EU�9�\ڭ@o��ȶ�꼞������������@7Ct��M�b��?rBv^���2���5W����/�A|[_ [k�4��n?U`#ޯ�9"��n��ޖ��w���I�e}��k!K{G��oǲ� ���@��"�b�!��`����U��+��U��*"��p�V�?<�. k۩�y�{��@���QJ����b������Hlux��J�..4^#�!�Y����e>x��A�ź�B�Wuk��3)p��{wJ�k��
������'g�����Kt�#r�ϖ�+����y�]��na�z�z;Ld��&�e�i_L�{nm�ڤ�=������6��ܧ�wa����R���K+�5|���k�S�	$����~��H���^~��7?-�=�hY\ �B���C޼̾�~��.c�=��	���0���_`zv߳�Q�n���mT
��5�U�� ������-�d�}��e�\�,�˹��](BΡGem�`�C�ՙ��l�W O����K�t*��ExO�쯔���m�[��͠iö��4���K��>��3s�Ҟ�4,�?^r?>A�� ��x��zX�f�Z�D��Un�:�����3�hۑ����f���B�b�����{�Cu����S$N��a���b���=�?l�D���^�;ڝ�m��l�g*_
���<�-��=܆5sq%�d� ~>� ���_�7��xׯn��eP�0A��H[@6�Ku��+/���� ��U-���ڵ9Rs����w).�O�½�.cʧ%�;f�SG�׷Y$N�>��\�6:<6�ne�fB�n&�8�˫���> �ݍ���>��Ol�W��rA|��6�X!����=�<�vd��!�X�9��6�Z��!����������u�+�W���/ʈ?��/�ȅ�����/-�١_��_r���U�d�w��A|A��o�6�'8�����������6U�2h������::�i�܀p�M�tYI��MJ}_r��ϣ,�+��-�`�[��v�GfmM��*{dв�����_��F��n�n��"�m��8�͖4��/�Ú�k����fp��\~yK�./���}�*�W��R#�H���_��h/�t6�k3ی�ev�����pm�6A�� ��u��|�|����	�J�z��h�UV��|{�X ��;���Ȧ�v��rh[_p󐿈̏�>9�6��Q��ܬ-z�ޓ@��
��F���my/*2��PIc�-[����o���?&����		3<}v�?~�,����tvx������ ����WᏙ~Ucs����w����8�@�ՐAn�x�^���=@���!d����m� �gF�L͌��Tp6P-щN�l��ʂ�ip�'�G4-�@�v,��f���\�k�w	^�P�{i3�w�/?@]�X�Gr�/�ͯ�-�`��"73�F��@q�A=Ծw�х�M��ڞr`[_p7���_/���:)M���X��P_l��6�Y��?6�3�N����h�`�(��z�V7 �4�.���>_ [j� ��"���wVb�C��/���6�X=܆>�R�{|���5rJ[����1y���/���[j��H��k�mJ��
�Z�|�<�n;��X���\��E�?�@[��t<m�ÿ^�\ߍ�^����w��j��1x�w��8��eN�a�]K�]7k��5R�p󮘻hb켙n������,��:m��?�ӭk.�kx��s�B�z���U�3v��'\v�q��^�/���\�y�֊�MÄ*�Q����z�C����we"� ˍ�z�h��I5�k+�tekK	��g�!�Y�tbj�VFb5Ɣ�n839�c��xpM	���]���Z�����к=C���j��B+�;X���ŮݮMt��jwV�c$k	�.݆cK�0Z�ib$:�6�bj���������m����v��5���Z��`��Y�EtvQ�F�:�5j�7e~�3�.#��ѡ;ڝ�MΝ��l��9cs���bU�m����=@�x��_"�������-�,��Qe��n�"`gr�r���<�)����\6A��@�/�ł�ɏ�z'ݰU}7�1}`�R ���|[j���+�p���D��q��<�����y�Y��"mذCk�,f���|��'eq��8���_/�n
�!�r���q�b�~yH:;�U9�B�B�U�	�H��	m�Ch"��]8ﱎ��,�Eǧ��{E���5w� �rłK���4�_�����Qڸۂ�U9+8�ua�k3a��n�Q<�t�m
*�]�f�ت��P�c��b���	n��[�S���������;�[��`�5gP@[v,A|�
"���9����Wf�T�r��߸7���w"��
����)�v~�P�=/�F˾�N�Q�{���_�^�wu�)u�� �s'޹q=�GIU�C(��7\uX��R�������\l@i�#r�FH��m[���c��ezM��M�z�J�h�A���� �u�6�@���-З~u�6�7Qw5\/��s�X[���0��u���8��~9�B�yp;�l��-1�@��lY����Ah_�7�ř3ʯ%ZZ��K�����%Ue������^R�����[���KA��U�$Qa*�t��P��qp;5���ư�H��a���qp��Z ��,\A� �mؿ�N]*/[��=^������e�@[�в�v,���k��m� �[�����7/M����;U�A]'���,j5���8���{����V�1r���ŀD� Kt�Ci|�}�T.�p��G�4߈y����9�A�2�'�Q셙�[+^Y�~U��X������zZ+�z�k�o���'�����.�z{Ȭ�<$�Բ��~��-����|��]%]ۢ�P�A� y�@[v,������Kl��́�}r�	d&V�U�c��րm���� �E���u��ܧe!��{eV:��p�n?��~7���_/���ͻ�9p�*�ЏX������8�ȥ��s�Z��HF�VY�9�Δ�,�θ���\?�=�x�n�A��; p��7\f�p�`���R���j�|sb�A��H������*V�n���L�U��Dև{�6����7��@� �� A���Cy����;��}9�>��ߚ�κ_�|�-�dub��f�fW��U��=6[��mp ���/�P@�A AmزA���=9doUFv�3������\Gd�7�M�K+���E�3��	kb��a^̲�9�(�_c��[�L���*�J����y޽^���O%5@���Ly�[��F��v�}������X �ߩ�"-�,�A��^�:�� ��]�,ˌ��|���o'�pw�}����Ci|[_
���{7�y=��|@���ZB;Ld��s�m��o�8�hn۞ {m��E)������W��?����ڰA �IUc�OG���[\G-w<����{�{5�t<�b�m|�-�G�άaү��_p`�D���_l.#�	��u�U�� ����_/�mk6�Z�*�E|�}{^��sZAm[�� ����=�N���Of+./7��o7���|��A������ [j����yנA��3k�D|��[���ڔ�p�n?���{���۽c��[�@ݖ,�@��"h_�7��^�y�p�~��|�p�GdA�7�뒫~/)�y �Y��Z�0;D��g��g��~i]SEA�[.�Ռ���*����R��꺛��{���V݂�+L��7OY�����@$�O��*���6�z��.˹�S�G;�u��j�@.���λ^�v��\��\W-�R+��٣,#�SE�k�B�	,t�K:��ۜ����c�.9�˷HtScs���-�H��v���r��W������(��u;�r�H$�O�Çw	cm�c;%��;w[n�c6�p,�T�s����)�IYu���q��m�y�K��ߟ����X6���m�tf뛵���"�C�x��R�h�Ml�[���?�A>|��A�-�_CnŉP��w�G'�øm��cr��A���K����Kt�"�or�Y�U�f�{>�rj�:�z�u+tp�n?����7�Pu	Y�E�׎�p���ő"d��6�����e�Sg����%9�e�����	yH����_X-�7_xz����ɑ �A�!��������f�;����,��~��gW����Dk��|�E���	n�A��-�z�v��T�+޻��x�!�����[���q�[\'=�X �� t��b��e�]X׹�g���@MJvz0#Y���}�Y�Px.��/�sDv!.Ú��ؚ�?����e����k>|_�����H��0`��q�U����[��.�A��` �� Ct� ���ċ{f�W�������i���*���^ZQV����Ⱥ�}�'��o��d�ü��q��{��H��D�`��V��N������k��������<�L=����P>��i ��>�+�v�߷Ϳ�s��<�S?P|��%����ɡ��P(�{F�cI3(�~��{u�f�AH,3WpR
A@�?Y��@���S>�-$��³5�)&��̳L�����Q����o?k,�����"����y~RC��G���ڰ�$�P���H.�$��XH)�
a�w����P�32ͤ��S2��H,��;���_s�����ɶr�'�) �Q�;�i��i ��@h�RQK_G��a��It���㟀@]��'��YL�����JH,9ϻ�sXR�}���)&�)��d��H,�2�2��%$�pR
A@��4�R
ANfXH)��L3.�5�������u �D��~�^�������9�~��� �~��$Je0���MFRA@��m �7H)�@jj�)�$K�H�:�PY�����e��-j���n-�\��9�y-NԹ�u�h�j�y�,:p3q]ij���w�4�D
H)=�����XT�kPR
MRfY���Y62�2����������>��s���v4�R�w�������]�ݚH/F$��XH)�
a߮�L��P��Y���q�$̠�CI��S��S&�I�kgU����������I9��Q �!�˅$��ܒ��+�x?����-B��$Td�����RAaGo�B�
MRfY�Gzݷ��s2RAd�R{T�hJH,;]���AH(�Y���`RAJ3,$� S��RAH(i̳i��������;���Z�V漼�A���D��t�s�X��F�%���Źh����
oԲ��.<s72�X���s�v5e�6�a�.�z�X��o^^���WfKB�Ui��BP�����;��H쒮�E���2�G=p�wBEc_��|��)�8��+.�L�p����.�w���,)�U�zjم�o�J�x���R��7��G��<�>�h)\�q�݁
C���X��q��̽�o������ȼ�gc4�0eu�z0���TdL�S�J�/��M��"ZxT�YR4n��v�����9���[T1�fu�*�;f�9WN�X{��&:�tu^���cuL���s�ifM���u����|�d^N4�Ŕ��v�f�e�B�!֮ix�be�ߞ�I����o�-nb�N��|�����WkZk�:��D��ɼ/jb�����FnЋݥ�i���ƙ����^���[O��[T����l5r���Kk��,W׫k*��R�l$��t��7f��[�>OW�75��K�,y�R�O_�J{v��V�aUgzL��c�O��ܥ��v�ά_k�dF�	'h�;�][��Y�;��C�ݢ0�	I��$�m0�=4�z�V���t=\1�D�9�f����ٴ������M˕�m�w^h-U��m�.ɒ����M��2F"����D��7+���Vn��W���\�v������M�j�O�-�d�U�GC*�=G'�պ�
o��Wi�(�GQԝE����㬬����(���"⣸��8�β��:�����ٵ�K�2��ᵶ�N��s8�f�;���;:�8�����Λvt���R���8����"���Y�sn�(�
3��ӻ:,�uQ��n��Q�Q��gSnZ֗Y�eM�㳬�m�C�vVY6� �6¤ʲ���+Z�a��-sm8�͛1���[l���Y�E�ɵ5�:.&٦�e֘����q6��sr�ٷq6�Z6G�� �u���l6��.��r������so����C�3��$Je0�_\)�Q��P3=f�q�����D��yp���)3,�AH,׵�����N&�@Z����$�)���d�) �̠-5���/���p����s�����
B��7Ϭ�Av0) �+[�wU�u���
i�v��S4�I
�}f�
AH)�A�CI��L2��L�I�3F�
AH)�@z��������o�ޯ� ����.�SS}��Z����}��w>�|�I��I�2RghCQ%$���RhB�32�2m��Y)����{����;����P�йA*6�]
�uf�=��_mWk��\�����PطVkP�q.�f�:[����ͤ�J�?{�i �`RAJ�XH)�V\)��) �Q̳i��Ͻ��f���߹ό�<�S��>�Ad���_�������N0ʻ�$���|�F�cI>���j�)�V\) �̳I��(d�̠-$�������ڮW�}ϝ�/�Ƿ�) ��Y���Y<�N�h3|Ϲ��-�8~��o9�Ă��v�I!�P��i ��
H)Y�����@�Yp�f�����ʳ��>���A@�uf���S���M2�z��L�I3,�A`n4�S2�֨��Z�˅#�H������u��z��N�x���?��;��
�Y���(d����RN�څ$��̳L�e$J��̠-II�VXhm �7��ϵO��s�Y����I*~偤��@�W����P�̳i��Ͻ�޲��_�s��bAN���CI��)����L�e$	 .�����,n�--��p��7>�n�k9���Q����}����`v�+شB=�<̿��5z��·?����� ������"_��I4 RfY�؁I��I�@ZAH,2��I'�)3,�%�y��~����ɶRot���p9�}���N}?G���-��"
A@��Y���
H)F}`i ��0�˅3L��P�̳i�ޛ�}x��]�z߿���с6!�pB��,�:�["oQ�g[�[Sh��#k���ط���8S5@ZAH,9\�S&���G��H,�$̠55D�ЂK_G��s�.���8f����KP�? @G���s}�;;�;�� H~II�N��AH)4R�,�&�RAd��L��4��Xf]��I!P�3,�Av�����	]�_�����+ �AH,9�,�2RAB�3�Y���ܿ������������C
g��4�R�]�d�) �Q�����H)�@}��?k��מR���j��@��Y�؁I �z��4��
�֠��B�32�2n2�%FQP-��������?��G�k ���$�v$�B�~��$c�
TϬ$��2�?��P32�$�) �e�4�Y9���_���2,;wpY<���]��H,ƒ
}�i �H����$c�˯��3�~ q ]��I�@���)=���II�7�̷����y �����f�6�H,��N�@ZAH,3.���AHPU��i ��
H)Y��
i�f]�eW7�9�}����� ��Y~u�q�3��Vf��?|S?P�R��'�) �W}�H,�$̠- ��G��;�xN��a#mzLٯk�9<��}y�w�w/���Ѹ��V�d�5�&l�pt���u�]h�[{��B�k�=�pM3҃c)l`���g޻��~g�<����;���]�u}���F�sɝ�5�u>��h��3Ɏ3��2�	f�K�r�.�ȗ��[��Zm����+:�N'�5��\!��ݧkX#]]�]�˄ڗf�F�b)���A�J����p�B�m!�����H����k���<�0[��#��y�\��*���V����2F�Û@t-�cB���֙��Y,3[F�:a�=�������6m�oF��(m��n:m�q�7&�ظ^�����v@�f�� RAe2R~���JH,3�) �fe�d�e$J��DI@@���G;k?���H��w �<w߹����7�^��f�
AH)�z��AH,=^�S?��P�̳i��RAN�i�L�Yp�MFRA@�����~}^� �AOv�Ѫ �����>���/��3�~ q +�f��I�)9���JH,+���I&�
@��4ɭ}�xr�=�4�Y9I���R��Ѵ����9�I��
fP�R��S?FJH(R�f���^�;�k�MB���7�NŒ�Iþ�R
o(>4�Y)���}p�M���S������S2�樂�Xee
j RfY���Y��������L�i���В�
���RAI�)3�4ɰe$��( �Ĺ��'"��Y�l���H����
C�9��4�R
AN}��3X����?�}
p@�^�S4�I��4�R
AL�i �Te0�˅2i��P32�$��S2�﯇����r��������]�.�p������w5���q~��s�<�w��'�$S%'=@Z��XQ��P���HRfY���Y62�2��{;^�~���w�Mi��<n��ݚ�A�c\��݃:Ӯ�B��	Ye�d���Vj�$�Vm ��}f��$��`i ��)�V\)�d���D32ͤ?{_}����9����}���i �r���}\��~j��?0�r�L�I��Ѵ���H)�P5D��+.�SB fe�M�
H,���2��5�#�O����;�V��ߺm�<�1g%f�����F�<�L�ne���̦�C;]�ju�U�w9&\1���}�
�a��&�w���ug5��w�|k���������P=�٦O��H)'� " �='�2,�՟���#�O�;A�t�RT?}f��$��XH)�eB����3��H(��Aa�aI=�!���X{*ɨ�H(��6�Xi �e�Q �D3*H)Ͽs�����>ų�p^~�V�z��X����(d��hCQ%$;��I&�)3,�AH,�e&ehJH,3(4� ����~6y������,d=�B���m| �~���7V_�������@���>�}��;u��T:���q�bA``�AO��5� ��3�$�@�̳I��I �ehj$��³.H)3,�&���{}*���s�H,�)=��?_�ߎ��U�k��3y�H,?v�i!��|��$l
H)S>�4�SQ�fT-�d���!��m ��{�5^����!����V��IZ������%#�\�\R<D����h9�\��h¦�t�t�?dCI��L3*ɦRA@�}�H,��S2�Ѫ ���#�H��NW�w����G�~ q R�,��Y��������}�IiߨC�JH,(�높
A@�=f�
AH)�@Z	I�e�$����i �`RAJ�{u�������뿻�����)��P�j2RA@Ͼ�I��{_{�=~���o��ό��
g���Ad�S�T-�C) �Q�����I3(�\�5��f�AH,+�B�
A@�;f�
Af2Rw(H)�eB�
A@��4ɑ��Y*2�2��k5�kC[����Ւ�����!Ok-��=[�un���C,즄�V�[{7d��>���w+���Z�0�P>�%T��v<Ī���M)(W�|>����;.�fp�sH,?Wn�R¨��4�]�
H)��H)�
a��
H)fe�H,6
fP�Y:s��r����0�j�L��I��h�A`li ��@kTAH-!��
G��	�>W�w����G�~ q %�Y �|2Rs�����XW�ƽ�s��w�����b��޳I ��P�Ȕ�Xee��i!U@fe�H.��
fP�R��S=�~�eۯ����Ă��ڳI���}�>�o�k|��|g���Sߨ>�i �P�a���S&�RA@���6�Xi �e�� ���˅$u�3����oL���Ut�ݤ(�l�]s�/J�_�Y��[���6n;4#��U��v�;���l�z RAe2R}�����
2��RAI�!H�f�6�H,��̠-Y���t���U�߾9���H,?Wl>m �>�w_����_�4�^�
H)���
i�ez�L�%$(C3,�Aa��$̠�H,��a��
d�e$
�u�k�_�z��ᤂ���TAH-z��I4wٞ�m�o����7�w>�|�I��I�2RghCBJH,+���I&��̳L�ޝ�~��e�b�R
{��hJH,?W,46�RU���H.��
T̰4�R��S?��$�x��?��J�5������v��{��a���
{�i ��z�L�2�
}�4�XH)�@kTAH-D2��I4�H�f�h�Y�{���'�����%$��P���HR���H)�l�̠ ���1�.��?�3��>�2��H)���I �l�p�$��*���Ņ)�/3��ݢ�P�9ws_Vav�� �;�ﾗϩ�;!H����h�ۛW�.�|���������䂟�
a���JH(P�{�6�Xm�$̠�H,��a��
d�) �Ws4m �7H)�@��/��M�������>��N�I5�{޿m�{�|Ww��;��
�Y��@��ʌ�����JH,+���I �fe�d�) �P�L� � �����o�WY9��U$�Nn7Z��k���7푘�<���gWQ�y��5���m �*U�9f�
AH)�>�4�SH�+.�2RA@��4�Xl�}ϱ�O��[�s�>��
{��H,�ϲ�{����߷��Wn�R
���F�cI>��
At�^\) ��)3,�l@��ʌ�����JH,9�~��7[��W;
H)4!H��4ɰe$Je'}@Z�5��=?g�U{��f�������
B�P��i ���z����@�Yp�k]�ߌ�~�������~H(p�e�H,6
~��$Je0�z�L�I�3F�q�����Q ��^\) �f�����;���S�ֳd���? 8��,��#�ᒓ�@Z�) ���څ$��RfY���Y62��@Z����+,4�AH].gt��3?t�3��I�`RAJ3,$�@�Yp�i��
�fY���s���~��=�:޻���6�Sߨ>�i �S)����I �W�����?{�R�i ��@jj�)�=yp���P;�f���R
fP����XQ���$��RfY�L��s�ou���}���zRAd�Ro��h�_}�}3|��߿|s5��8�X~��|�AHQT���H.��I>�i5)�V\) �4�fY������~����e�z�r�"�Y��%qoN���T�f�BW�K�u[��i�ו$q����Mq������p���;�3_�)j�A�*��������V(�~�BSƷ6��=8L׷q�n&��6�ڝW&���a���i����1��Nu�w<Hl�
����J�<<l��sƮ��T�2TB
C[.c�hb��2-��5�&�6�c
9K]vJ�.Q�GHn:;
z�8�]�P�!�/^��1=�G>���`&뚹v���[���:��.Mu��l�-աlE�ǿ�������7Mȶ^ck�����y�-��t�`�j%t�-���AK��$JS�n�R
�w�H) �e�Q ��˅$�����5���|��o9��@��O�
H,��w���=�j��_k�I�����%$��B�
MR��4ɸ�H,�I�@Z�RAa��
H)U��i �`RAM|�_��Ԗ����AH,=^�S9) �w�f���{��gt�{�y񞆒
~�i����}p�MFRA@���H,��S2����}���ߺAH-!��
j R��M��YL��}@ZII�V\) ��B�32�2m��Y)����~���~��gś�����y�����3Y�����ͤ�U�}f������z����)�V_¾�$�dH��ݬ�c�_����=�:W�鐀~��/�t�^�Mq���A�_*���o{-��_0{��T-�,����7ww�\ڹ[��ue�>}��m�{�{�!��|x��X�Ch��!i�nWu�hT�䬧3������n\T���-��q�lKq�;b�z6���Q(~yH]q���A�Myƥ�۵ٞ��:G�g&<�k܎P߈#9|�> �v,_ K,�y�}����q��gV�(��	���K*���ؘO��T�ms�U���2��A��]�D�&�Z�s4�&j�k2�k� I��Ϣg*Y���|w0�ￜl���_q�Hv��[hb�$�^}���"��m�d�E�Q6�.�u�1If#�1�|:Ym��A���<P#dB���!�!�VC���/��� ���o/��N��Yg6�g�3��@�y����``�� ����Ci,��6�Y��w4����L#�c��K��䞍�k�JD�Gwj� �Ո5w�J�k��g��ն�NR��mU`ȍa�]l�8��Pm��"֚KG��_<�Yl_2ρ�b��΄��{޶�D=(e��GH�i�x�;%���:d"�_Yn�&��I�nc�퐄|�Y�I�>ih�wg�7�#���e��r}��Di��7�Y�,6�Y����!�c0`�(��9�:�W�R%[^��kMtҴڛxfH��l�� ����n��������줭j�YV�PU�Д/���L�s*�%�b3��g	�-���f�Mq������HF��m���� C-
�s3ޕS�A�:և~؂���~mس�Ud>���J�̫�������� �r��W���D���Sy5,{L��ʄ��z��w����`z�A��o�,~|�-�@�v�mz��nY0j5g[����>P�;j玱whspt��/[nt:�ݪ�� N��ł��m|��=���p��ϧw��A�J�x�{Pg>��2r��-�2Я�h_�{پJb׾�fh��,���#Գ�n���C�><P��U{5�/.��U"9���� �L��Xͣ�S�0y5ɒ��8f����;������A|����݋7A�
k7oԃ�a���`G�/��B���N��s�d��}�� G�f�\����63��4y�W�������[O�ѺF^����xkNm�*�⥯MLʼi��s{�N��_�ߠ@wi���oH���u���{f�g{e��ֹ���۫��|��u�Z�g���Bg|�Ǌ �,X!����L����~����UU�ʛ����r|=���8h���R��lg�����P��z�O:C������-�^��2>��	;���x!J����W{%�d��|�>۱d6�%�Q��:��/ۼh�Ƃ�����T���ĸ�6Hk��|�\B �վ��k�;��㊁=܅��Ye|Cm
�oX+��v�2�*�����?G�,����g��ψ��]����z�B9"��t��t���Ŝ7d���(~�,���:�0�!��
 ��,��e��mؿ�oe�i�5���=^!g��WC����~�#5��%� A\B����n�����y|�)�5�㬝��}�*��osr�M�]Uj�eM(��;�-)eP곕ZMf�����[ط\U�m��:��Tz��d5J��&�^�vR�n�܁FzCLJڼ����v+��ں|p��YR&����(�_tp���۩O����MԳt�wL�Ɏ�3�}���8�ydUo��m�j��>��lfve��=�PNw0(P��(�u;�L�3f}�b4��Ml����jJh>Խ�\�d�^MP�����,,��</+x����Y���Tʵm#�%�^�z�]�����jo]�Ҝ7�3#�gQ��gZ9���̇���G��C���ݜ�0�ʮ�[�e\0t36�k0&�[R�pw��;��#�������FZy�ĢN�ŷ�κpν6:�Q5���W*�.7*b�g�L����ћ�Q�[�5͈mn��[�v!���ǻ�w�A�kr�R�<*��{ojċ2b{X�VF��S��Cz�e���t%��W�]�te��C��t������<���S�����v.�GyJf��S�ul�d��1-��h^�E�7UH\A�J��ca��ҭ�ry|�[�v�6"�}��T�j�6����_m�:�ż�Ua��Q��	�Mu�J�HR��̼�,���y%Aq�	�6���0e�U��늊�2��G��e�7^jy��;.CH���fz�"d���o��q��T���WA};����Suk̪��z߭�,]Hӯ{s'u�U[��Y�\��t��YkWe��4ZJwl��`�B�һf���@�3A�O�v�u*�u}�Yw�=p��Mf�F�w��U�����#�A �8��2#�ٙ�t$e�9Y�-�mf��VV�I�GVu�H$���qvRvve��Ʋ����ŖM٭�6܍�t�Xfړ-�
�-:SM�t��[vYc�+Lmvq�N���9d��l�E���'s��G�Y5��7����q�݄��*M�e��֒%��[Y�j&��Y�c�e���h�+m4۵�im�ƭ�kI�F� r�[s��f�2�%	9L�8�HR;0��sf��� �6� K-r,��eM�˲��k6:ma�'"�5���4ے�gv�B��X�C;I��&����Kk�[+��)��[l�ΐ�Hr���Ç��)��� �lN��#`׵:��h	FP"6U����JZ��:ٍ�X���r�vpmԦ�`�bf�`��03MjcBӴ9�rv]%�!s�.u�h�`R�p�1ڊ;10��oR��z����zr�\��[[(^�g�t�ڵ�0�fb4�az�f�R�#	�����VQ;����v��Zk��)q+�aE%�*􌝎�ѣ��s�����ϙ���<��{�,�p�>�h5�:�e�}��(T�Ż��z�.]�8�^źQ�z�.���Gxx�:�:�/m0�)�YM36�ڸ��C�c���F���a35��E�m�2و8��V����mP���:�Ӿ����D�6e�PK���ckXb�[��&��E��m�	�#l�%ij�X��ͰB��E�GZ�:h�[gd�9�u����GCQെS�ŐE6�c�Rsۥ@�=d��a�@�����*b]cu5�XUP΅�	rKơ��A�,ҹ��ҏ#Î{$Ǔ��A��oF��3W5�b]a\E�4l֤���XS���n
�e�	����oi�O���Fy�C֜��N98_�NoVM��"!��ut�;��_'�	�y�:�l���h:2zv���!�!gwB+l���X͛��$�s����R�0W�7�XQ���ts.���΋((Q����AKc��yzv�xeN
�@2�qX%3��Y�-h�V�+���Aã*��%!�u�M6e���c�Tv,Rgn`�5�"�<C�����ێ�Ҕu�����d�x(쾞;v�y:�籔�n��6�p�`k69��=�.	���ڙω|�y	��z뗗�\+F���R�1��G&����N�r��H�J3�6"�60=�E�,�ɻh w�P���7cn����r����Y�ГO8��X��v��)9��6�;WmX)ƞ�Ѻ�&�3q�Oi���Y�}��}��z��
X8��lR�%��4A��n%GD,Ip�5�\�J@�355�W��P���.�@pl�6{\�0F��%)t�1a�`��3O9�������\��]
�-��a��o<1lh�tuɞ�=�5�8��#s4D�����[����`�-�t�mݘ%[�J����æ��ĥiF8�VG����͸$��\o7i�	�u�f?~
@?�-��͊�67lF���ۅ��׮ՙ�:Z��n�t�������LB�!�ŖQ�yoN�n�o���!7���fQGH��,ܗ��!�VA��򥗷��^�Ư��~�+��Ŝ7d���q�r}AY=}���C�{���x�Amز5Я��f���q(fY��๗�}��i�\��4�Ŷ�n�e��~F��6�+hx���g�����Ħ�Y>�y������Z�-�������=����mY����G�-�H�;~��V��x'����'s���^�����|A�6�p��˹u������Uf�;M���9i1�M�j�r�����p%t�-	�ӥ{�x��d[����o�#7�9�b�B�0a�]����0A��+� C-Wʹ,�;� ܽ�w�It藸|ѩxQL{�U��e�y6g��oX���2�?#�:�g�U��{3!�g�y��drжc9�5o�>���8�!g��¢݄����!��(D}b�n�\�Qf^_��N��W���e��m� �wT��T�N����,�	;����ߢ?tA|Ye[v,��/30��ǯ�����C�|�"�j1��*���+W|A8���ws;�c#���zz�^�(G���nu��w��_��#�b�2�eAQn�}�����|x���m|�.��+TR>��6��7�>��*��2��8
��C.�Ѹ�f ���v��a �M,*JiG2`���,�������-���[��I�=Fߥfpݓ���Cׇr��9;��l�X��GK(Cn��Ct�Q�eu�5�r�����#�/��-�F#q�uA�r9�j��:@F�!|[k��7t���g�@�_���"�(��B�E��Qh�,�{�+�,�g��΄Mm�����E��M屌
8�/43<vؓ{�t����藬��O����m��_�s��?�!���(!d7_2��-��Պ_�K��|�`ad#�����*L��6�3��2xY�+��@fث�
w����D�Ő� Ae��mؿ�o���t�e"��T��_Wx������Aڇ����k�U�~���M"����M�
��x���(r\��<�	S�s���j�mF�lK���B� � �,��-�꽒�Tˌ�7ègz�G{���>�px��,_�H��:d"�VA-�"��T�2����W��+�G�����ӲL���7腐~�,���t'w�~�Bް7p H�A��b�����m�u]*�9��m71V� ��� ��m�� ߐS�f�0�q�dM��#�/�m�c���G�ˌ�c����ʈC��9��C@�������՛w�9���}J�Kz��wb�W���K�y?avk$.��`��^�ma!�ys@��� 적m� ��"-�@��˧��N�0o��*��6�w��;#���ވ_�"m��5󝚘��0/����Jt�EB�'�J��nͦ-��GJCM��MK�l��*�5�>?̟?�~�,��[��R�9=Qu6�̺h;$�	��r�tǣ_X-� �Y��B�^�琹�j����g�>B��tv���f8"���x�ΰ]��V�t�j���B A-���鐋mX �[�f�YA����j�z�i��g}@�}耾��Y���!��絮��V�Y���b�_'L�{�T����u�v�]E�u��)��s%l#~;����e�@��B�?�E�}g+�n^n{�D�cM�tw�[`�3��><Ql�z��ZCp�Ǟm+~�C����g���e����'s4�-qI�]�uC;z3�1��a�Z��C_?Mg���w�y-�6{�ܶc�%U���roT"���	��le�+�9��JX���B��/j���o����>ź���c���P�cɊ�W�ٞ�l�U�6����v2-�X�0N����=��q���k�y�jМ4ƳK���9�hå��d��wg��$�J��\Y��I�Xl�gl,;i8�
�m��:��O:��ڵ`㎋sV�u�G�4����eΩ5�h�M���[~��݌R�4��0̩pU��-�U�X�[9��S�IUYT�T*�6��vW��<[j� ��]$z���Ӵ�g�3�[��7[��^ �f�m����ٕ���g�n%�B�R˷!���ۙu��D�E����ě�b\��j����5�@��v4}]����J�X���.ۚ6��l�oX�DA}"�2J�F��g����Z���ρ�.���w��vG��ވ_�vϥn�P_:~��CiYe|!�b�!���3�x� ��|'.[W��g?f۞�����@����� A �WY�`���q)T�tP';��a�9�4�ڧ�ݱ�:�F��3n�=v��2u�Bȇ`�~31H��P!����J<�?1^�gC��C-
ir��;��K,�9��_2m���t���o��w�nG�ޮP934b9}��e�jv`+,�̝���e-J|��5$��yVi�TI�7�)܉�c���Vޜ���V���5`��*���U.�i��gP ��� Yg�;|��*������0�Amذm�,��$��Do.vo_�~ͷ=uN����"�V~n��2С\��͢0/w ����> ����� ��J0W�:������u�Sn���p�w���/�T!|[j�%�D2�E���Ulsط�����U��������vG���	������|���%����7�N	F�!]�QWwh�W`�m�KC�y�t���]Ab�.!d&-��SX��={����P ���n�e�퉫T��0�_W�]���J�{{���:��j� �H�!�D[�Y�4��"����s�M�^��b8 Ah��v��F\����B1�}fr��!%Y�E�ݬ5�{����ʏ���e�c
�UE�٠�8	�ZR̷�S`A�4����RmW�Ѷb��U���[�m0���Yv+7�1u�|:ݳ73�޲��G��Q9�Y�9�,n������_���E-P?HW�<�s��N�_��2�f�t�=���{����`���i���b�>��[���I�[����.r�8�M��@/�:E�}y�dv�*�70:�c5]�E���s�����N=�5�X06�Z��|Y�wW���ҧ�ehR��p�q��Өxn-˜�g8����QQJD�W��P#V�F[�g4<G��CԾ%�_-�\d�[����qq�] A��wuB�kWeg1r�����ߪ�j�G��4#9�,N4���f���GU�>���wd�d��TF���L�Y��.\G�C�r�n��ї�ϕ�P����V ����{�%��nc���慑3Ee��YЅd���	�1ք%��S�1=�y(�� ˫����_WuؼJRȼ�q�E팦8��'V��w���(x�A�I���~�X�$���#����씫s��4��A�H����(	�u�i�>����(�tPA�rq�r��,2v�c�;n��m[����~Dx?P��(~�%�S�}��hu����?Wͮ��s� ���X#��$�����&;'|����+�Hm����w~����r��_/4� �x�\ݫ����ł<��D(d��_��/*�>o��p�k���n�6����n� �"�� �dTЅ"�n͖��f�l@������=}��B{���G2�F<��>�dw/����L����IX<����uy�.����H	=�=���A���r���V4/�A� �_wv�o�z�����Jf+*��<k(�4�nޞ[|��^Z��U�M�`��.«�:�v��x��B^U�mBQ��c�g���U���?��DC�u4��X�z��C��n��!.�
L�����Gl����;c�n�Fa��4&�4&��V�[�ó�q�q*�HFx`eD�!]5t��SW�A�*�c�����K3��
6)^� 03@�ٱ��4�Em���	U�XT��m� ](�c8P���`řfU�y�D�c���լ�p�]��02�)7��|�d����fR ��Xԩ<�[p�ׁ���h&�+:V�Tn�E�Օߋ'Z�����|N�B�p��ꞞU��ښT\ٶs�4zOz'���/�{����@�$�d[��'v$�w�2� �����h�v)a���j!=C�f�� 7m��㞖��=���#ޫ��s��^r��_���l�ݥjl��~�@���7�a��X������L��A�,����"���uL��7��4���uDe��JEeI.ȳ��	�d�,D�(kǯm��s�rV�ɑX�/�Z�Or��A�F����.�&
~(V-".�)��H!�J���ڰ�àj�F9��\�X�2��������}�� �%X �"���=�J�xZs\?N�0vj����X ����$�`�(P �P#3ΪB�����d��^���74�V��wA^e-n��VK�Y���1Pҡ%���j�7���hf��TI����� �sv���U�����_�"��6��L����ښS\A��Hǈ�����;��ⷬ�O��f�P��r���'ݰ��޹���.�{N�o��mJ3~�"u��ܳBs�Xq*<�/Q;�Ib�uWKk�H "���VAv��n����g��5���ⵡd!�'��b��W���QΡdIT"2K�}\��k!�!��\\�5�ٻ]���&:��P;��~;�bo&3z�Ͼ���������>�ۖ�Y2&���0���`N1���cq4�JĆ��lИf���wϞ2i��(�QI,X�]��>�����s��^{~�[�x�A��/�&�|~0�d�d�� �<�F�y��r�A �K}۽�ڌ�&�~�@���-��!uZ�u�K�b��`���X�$_W� �����N5�E*7k��n�{�4�W��k�zv�<���p8��<$0�å&%�I<V�ޤ��n�V�n�[�r\������ڼ�s�#���]�B:�oi��~���uD��X������I�$(x*�o1ް�ț���o&�d�X����SZﳲ�Ž�W>�љt�VgA�pU���pCԅ+�V*�Lj�%�C&����	s|��a���U�yW�AgM�(7"ҵQmeLٖ6�}F*�[I��rśx�L���xVB<�rܛ�V��6�����lxu\�Nѹ��#Rf�zT��}u�yݗ��*���]z�❷v���˛18��k�5��v�_k[V�X��c�p�'}-&�v����6��'��mE�h�v�:;��ø��p�n���`��}[N&];��#�/��{:K[�`�FO>V�����%��&��}S��B<$Is��;����;���h��y�M԰�kc���x9�Z+r[�[ӷ���:`��@p��]����=�;�(�k���i�������y[5�a5ݫaN��\�@�$�:-�1���s��kv�i�.+���>7�S���*��Śi^LY���nJM�,��I��5��]����B����{^���%�cUB붻�'x��ʍ$����5��_�f
���]�օUnX��D�K����o(R<��oTX4�*�ח�X�z*#n9�gS��lI̠��l�e�@�s5�ʱ͝k �J֝�F݇� ��(�����6�mbc��֛j�3\�V�S�q���"�R	�A��H'�lڱ�s6�p����;���I� e��ݑ�V�۴gv�;s��;13S���[v�Gf�ZtFՔ��E��6�p.[jr�m�n�"Ln��"(r"�B%f���9Ŗ(���qm�:�m�m��δ�t����(Ns��`s�6�Am�ӹ�NGm��9XqY��:�s���am�9&nN��[v#�Ck8$��Dp�&�s�md+jԜu$r��pEN�J�������̜�m�"�t�G�GG:��Afp���YZ$��p���m�n��5m��@�ڧ��f�mHn.��c��Ǐۺ�Av���!l;��y��� ���3Dn���粮K`�;�������|�[/q�Xdt�_����A�Q��V��w=�n���!q�|Ǵl�ȩ5���_-�Y�
 �%�����c�.���,Y����ݫ	fL��1n���[���
�v;[#��|����}@a�nző%W�E��559藓��!���79<���[K�S �a�;���	�Q� �2J�X�*(U���4?f��8��y�Lvkw(Or����,!��I�fX?Yd/�fՂ	�T&���A�a��o���^�ѯ%Nk��)�,� ��D��,�ԅ_s��-�j��Ә�Ye����W�EA�5<�Ksٻ]�������Ѫ.ߝ���;]��KF3h��c5Kcg�PUO/�|�ƪ���Tٛ���n��Ն�4o��&��mV:1���I��1�t�/�VA"��H$�d�DCA|�C���lw��=�wmm�0i��n��8�hDrő������y8�n�I
�YD�z���[c�.�7b㤵���2��a.�גZis����U  ���??I)��U�7�86a��p���MC+-z�bC�>�#�I(	�D+�"b��11��ʱ�֐��h��+Ͻ߳��!��~;)�_�^X�wa�ƶ�?2(��(Q��Ia�.�c��]�oM]w�U11�r���f�}�dn��:E%X!{~~��,p��}1}���{�VAv��<�hׇ��5������²v�j�";:ő" "��,7x�,�+���\���a
|�{g���v6�7	�H~<E%}`ȃ�5[ly���-�>��Uu�\�zϖA=2�"�wQ"@[�����cօf�@�Ou��mUQr��6�-�x)PS#�dh�8MU*�mJ�#g.h3]����֐���q��s�E��#k�F{�Fр|q�a����m�n�]d'�Z����ŝC]���-�����p��nϘ:�i���m&�*��X7%$�שE���C�Ե�m��lʬ�)��Y��B��U�r�2�M,Skr��t�V��sG��#iY����6��nb݊	��K���տ~��_��Sbf$�#0K,&�ٲ�4[lㆶ�!�8���8��Q{����D�n��>�Wm�h�z� �!�uV�;�i�P���b�̹q���r��7�U^v��^-�`Ǌ��%o�y�7�^\�ЎH��� 4��7׃�{%�"5��(D�ő%
s�>R��o��cVg����.���x�;���"��v;���Pdf!_
 ��vŁ���Թ�G�k�aN@3�T��ݿ�t/�'U|~:B �*� 	��%g�IS���{������0/�p��e�,��h������{w���=����$3[��C'�I��؈v��ᇚ]L�8�سC^G��'��:{�#u|�?�PX3�>_��ܼ�7R]E��zm{�a�u��@�5d�� �/��J���^��W%�f��þ=��=��m�=]C���?���Vk��̪KZ�"i�ws4�U(���rvۏ
�Ȏt�u�L!�A},^g[�R{�g�k�aN���ő�����3w��M_欂w�����?H��n.�)����9��}�;���B=�Y�Oz��#>��w��r��{7�4A],Y���:B�����ܼ�7R]E��K�.Y��u{���#ϙrr��}K�~�	��,��� �8���3��r!m��jOy������
p@�C5�l�,����ݞ��|�}?i��奧�ؼf�
�ΰ
�ۣa�:Q\-��2��l��eBn�3ʾ �� d�d"�������A�y��?N�zxt�ŭ!V�=1�V  |� �4��,�� �4F�𜥳�a^���,0F����ȯ��ϗOA�y�n�����G�"���X6���ƨ����.J���X��4n��q�~�{}�6Ҧ=�Y�#���ϧ�;v��y�|��
�׎z��`�`�]T~�~�ܡ�$V���<�rM��y\u��`�s���9Li�����%G���O�������w����?<�0AEQ�����3�y��?N�Aw�����Z��)��|G��X����$�dIm�Κ_aD!�n�Oס����k��W� �* �|BIW��D�]~>���=�>��2�fh�^�K�D�:˜n�]-��,p�ja�-*�l�eU�3����GjD?I�xfu��'��b����;�;:Y��J^|D6G,쯈0��U��TE�o_Z��������K};�)M����!�u>.�A������<��łP_������/��2!��W{��uz_=���jCqq�?I* AD�8Z���g^���44Fb�4���xf;c9� ��ɷ�V�P?�|G��4��Rs�f	3N��*f�Mk6R�MΠ�R������`�NR���*�̥��ׂ��v�,>�l��8t��!�r�<�T��U�A2*a%y����W[}|WP�wHzI��a.���?B8��`{�(
%��t+ϖ1R%���뗴�Xۢ�kfi�f	4�W;����sfDB��nY��<�:����7Y�P_t�s[�G��^�6�7(������v�~��> �"���|�;�����\�N��M�#|A�b���c9� �}���O� �hd�,���?f����e����A8B��$A2��gp����c��vO�C1<7ܳB3޲Ӎ	�r�s�Y�b��z�W^���D�ő"�|A�)nlu�cޛ�}�Ԇ�� �R!qT�����S�e�"r�����g9e�C[��|�b���+�٩�.����[���k�$�Xn���z-�����-fv��x.���u
�ގ��pۘ�|<�vee��1/��H�wʣ���,f�����wd�iC�����#�l3b�э[�sNS�kC\C۠������i�KaX:�B�;h� 7gH�61[	r[�uy2�79���H��)a`���{����6��T��1x�&�&��a�A)K:�<c[����X3ҖuEr��� ��f����nLj�i+���<v1�q�ָ��6���[G�VY�c��K�t� :Y�kq���v�O�g���ܰn��w�+��� a3MY^�MN�+�́LQ]�U%i
�_�b�A:B2J�̊��&xc�(�%�!�p�U�e�{��~@@3Pl��@n�@���#W���9ەW��#K�x�Fo:�c�Ɇ�ͩ�J�?�Q��V��.�oQ���*�1)�2��X'Ns�l�{}�ok�\ǝ8�g��.���x[��FT����Yq���r��\5u����Rމr��(	GCGl�䵓���?N)��v)��G���$ϨW�%���)��U��*��E��uzh����jCqq�z���P;����lW�Φ��r�~������!�@��vۻhK%��iG��,v��u;l��bR��_evPǛ�G�YiƄC��f7�fz�a_�]L�!�溧#oƼ~�_g_ȝ��i=�ď����"�i4��OVp�+IbCP7d�d�>[����z�L6g��9�����9ud����7Ж�];ݼ��fp���,�9,������5άA�F���4�Ng!�p�~8��� F�<���{vL@���wlX#eW��<��^xv6S�[��~{�Cq���@����/��T��wW��u;��H��H0A����ݱc3{أ3�&���`��!�B��{�`��}���@&xW���*�~Oۺ�3�m ��:A�篘�v��㹌�J7ܰ�{�u�9c��,�#�7�V�@�¤��"��T+�(�/�y�<B8�nom��M���h�Pu����&{���j"o;�Q9�.#ī��{��|�y2�ڐ�\Eڗ����L�_�X��@����5I޽�a�e�X��O<���2�:~����<G;�b�e����|C��|Y�����B �*�&E�"2��;�R������TF��c~��r���JE�w39fSL�G����.,쓡R�_7�-�iS7S!���҅�N+Y/8w1���r�����DNs�4'9B���f�H�B� A�ؿ��B�&PIɳ�ٹ~����>�A~T�6_��>"�8�W� ~����Dm�d��z��4'�,t}�*1��/v��\��3@��rX�F��|N���߿\���Lf�I��i�`���5�s�nTph{kq��X�E�|��~�/_��/���A�F�l��k%����9��d�=]q\��<z�!DI(�@�������7�Po��u�:E	fO,���Ξ��o��g������?+\r8&Vz�� � !�;ޡdH��� �����L�{��`���=ދtc�Kݮ,;�!����,7h?l���2L�X&�߭{��?d�d��[�;e<r��}���G|S�F%ާ���[E�������$;�W؁B��˾��ǭ��v�r�tVZx`���<*ı�*�I�7�f p��Ӂ�g��~���(��hМ���i���xea^�d��E}�=�yL��Onw���yQ�%X �"f�^���hp�*K)(v����6��`뗣e���Z����3b-�bY���sY=|�z��5��A��#wl_ۻ=�F1ߒ�7(n��Q��A�s��_FIVAD8�7=_g��g'P�����'��x9Ӆ|�@_r�{h�qYae������X�u�9�Y��.\G���]#~��1��y��n.w�O���L�	a	���vr�]�]�P�!�(�(�%	&��tfۧ~���S��4]ڥ[1�Π�2/����P2J�~�P �a�*�����K��s>o�z��!�u
��{�l�$�4}P���+.0n�#Q��M.�Jfl���m_�&<��:�Zr\�f@���̢������a�!�y_]��}�q[��+ee�g�6]Q�{�d�wIoU�]e��P��~��8;��U���q&���x{u[Ի-g-�[b���*V��Ƙo��E�8n>m

-�֝����{�}6����.ۻ�Ν�@�����a�Y��J���M����}�:=Y$���y���̂�)�㘵��%��wTL���ޙw-Ƴ,ev[{�;q�S�??C�5�H�a�kM�͎��\�껾���'��)
��T���LYUb��ȫu�l4hac%i�ז+�`"��ә�I`�3��Sv7�5Kv�v�����F���3�_4�@^C�ɑ��X�˸��č̏�����v�jz����ћ&1��陫g��w����	u��(]�5�^�NZ�󐐨�[0m�=�������y�g-��:WU��u��$���Ү��+��Ms&��yz�ű�f`Wz��!G{��wm����`ˈ-C��PB������lRa\W#O�Q�wU�ah#�gQ�oV=��iF�����Μ^4๎�s�˹���A�n�Tۼ�mm��WiUG�}�,�2���R��}W��̬��ٞ�1,5�w2���)W�y�ٖ<ވm���i�he����e<ny��&y�h1�1���y��r���ۈKixed���TH̘�ע[�����7��Y��m3;�ʣ�����ڜv�����dۮ��1�ڐvv=�U^�1�QE"�UPf�.L�8䃸����	nH��� ٳ����,�r.6KI%g�JK4	ȗm�f�nԲ���5��$���K�fu��k:��4��`��8�s[lm���(�vvGfft̄�v�FY�mim��m�Y���	��֢BI'�rG9,��#2[g�D":H8;l��-���Km#������Yc�#��� J�Lm(��S� s�f�:)t").E��A�Ĭ�ܔrS����u�	�f��Ӆ���$�m��9��A� R$@,�	q�Y)È����N'r;,�25"�٫P��������ŝ���p⶚�ݠtvOoJݼ��zo/7&������O]v�g�gn��]$ �m�c�n�mi���,yi�ѵ��3m9��k����>>�^N��]�,�	��6Et6y,i؅�� ,9��k�b�h�<O�n!ދ>�V���lH�;�V�:�M���Q��K����h��u��ɮ!l6�[����$�Ã쪯Fg���nY��C�8-���7G/&8��l]J��,�)dFcm�"�ͻI�=��'3(�6tm0d�`�:�0뮉��\�ɼ/�ĭX�9se@�]��m�'u6}���˵.��b%
�+�`�{�v�N=-��q��2�]�D�q)�SUb�.�	�`��YD�����b��2�Ѕ�V�2�mjS-���I��݈����
��Z��>�7>_z��v�.Mk,&��˩*��h�ե�>���`ܼ�Eۄ0�ҕݬG�.��!�jCk�3r�����H�P5%�����[�u�l��c���\져4c�A��#�������K�8uE��c]���i)���,tf�%1��KUc��.�Ǉn�U&0)��Jɚ��̵�v��-6��t��S�`Rն3�m�cc���,i.�Q�Bq����n�C%�a�Ո��i��SS1��*�p۪9��mF{"$j6�u���=;O^��ù�c�m+#q�FU�u1IOs�^�r�[��v�K
�B�x)r�;n��3��x
�&Z�d:3�\�ö�]�Y�Ҳ�6w<ud�[���l����ʚ��n���m:7[i��z&��ԋ�>���c�sp��]��sMV�:��=��.����`+�P�t5ϵu��݈��ӷ�=\�����e�_VTc�.3p�Yrێ#aC��P��ۋ�͉@���4�k��sg�uh:��l凭Z���+�-,���]Ў`N���r�mn�sV���j���qbgc)5�K��\�j$.�!��%�M�픭�vqq��֧:��G��z���`�axl����jvι��g�J��W���n�8q[��n��j���St�o$�鞟Y̳�ŭۏ^��c���m-hN&�-�l��9��mә����:Ѹ�j,��uif����hX�]u���3-�-���v6�)V�N�1�m��٩;Tv�W�����q\j�I��Y3w���yf�2�4n�h:mS���YYrC`��w1Km�4ݵ׍G�����u�wG'{ͱ�]Ӆ��,S�B'�f�s�q%p���O%2vb���\E�A��g���!���EG� �(Y�r����^���7�����Lu�~^��,(=� ��Y�|�d�c�|E }z��������W������:C�4Ҥ����OA�t�?N	R ,w �ҁJL��oy�0y���=b��E���N�^~r�����ez��~"�wW�r��� L�����=���]����`����y1�c]�{�$�9��!�b��/���̿{����[}���ɭ4��d�n�P��a��OS�`�����.@� �C/��=*<�FIV&EB'���ު�|�i�D=��	��i�3}�h ��_q��bȒ�!|F^����l��f�����F1�s���b��T��}y�gb�kٷo���ˮ<�]���+>�^$���9��������J�t�Ǿ"uW�W��#3�Ϋ������7�<<�X��y�_y�=�k�ܫ�"ٴ,~��@�$��[�.������*1���ޒ^
�� 8����$�#�չuC�v*#��ڳ��!�׳���k=��!�?(в.V����'�uK�}=bȒ�a$�/�D�_%T��2�e������&~��8�^����yW�_/����;���������a�E.YH%�"WFM��`�Nrl�HV��Z��qd��ha������s�+�I,XK��oV�����/§!t���a[dh#;��7����%YȨ'Q��0g��9��A2R��r���g��r���A����U�x�=۵�P\ݱ`�� @:@�ݱdn�� m}����<h��7�5b��F1y�5[Z�nX�0D�r,5��)�p�RK�e�!zW��K�ˬ�n��nv7G50+�9}ozb�{��/�9�b&T��9sC�U��@&~^���t�-C!���A�wl^��Ɏ&5�z�d��S�"��/c�h��*��z��v�|G���*��ED����<߱iч6�n'�6�y�NB�򚅐GE��,n�:��j�+v�X�(IŸcn<u����'O)cӮ��EV�U�4m	��WZ֌��e��,�~������/�%�3����1l��/���c�m_�f�|�#;R����#r�8Ќy�Y���:���/4z��<I�,n���r��׹�s������$~�NA������T����c��q8�y�^�#�PYe:�%��j��k=�Ӑ�{�*J�#܅|a�KD�(%�CM�u!	�`gg���$%�a���zb��!�]��Fk�]&+���^�.��WsB�������&��v���hUu*�g9�r�:����e��am��wS�I˅M\�����^ʰA ���Q%"E�"�f����Və��Z����O8 N@�#�`�*��UOl^q��T�(�f�+��wV9�G��]����<E�U�%ķ\5"Dr���W�~ �g���2J��EB'�Y��k=�Ӑ�xs8�w�%ٝ��Gu}�X$�%
��f��Ke������HK����y�d����A3�|A�FIY��Osc��E_4�A.z���(���O���ߞ���m��ky�ޯ��A�ő%
����*����f{���IK�g�i���;���άpֳ��9g�MB����ғ�A�n��H��"IbȓzV������d�xg_z�������&r������";�=o�)�Tw��q��w;�4r�_=�%u��.~�\�'�ڽ�e9<5�rŬW���>Ĳf)S�1k�u�c�]�oQJ[�xV��>�b�y���>���j�3p���B��5�uY��0fļeĝ��ѫ ��_-߇}��w�X6Pp4�ԑe	���X/^����qd��s��4�띦H�$*�,]����'k]��!���Ԍp٭.YL�I�B*`ٳPsZӰr�H�aM��.�f����2�Ku�m	hB�t�D�Ƣ�i�b�%K�ۗI��wLطnd�v���z�Ť4E�Y�-��2���ߜ�����#��Ԡ�㋖3qh�гB�t�2�1)��ht��oW8�{vhD=�-�T#wP�����RR�~�c��_ ��p��f9	D0A��֗�~�� �� D��:����E{�� �:��X}�|�g�չg�*b�:D=����i��{�ł$B��"�ł$�_t���n�(3ʍ���$��y�C�ӕ<BIV&D��=�q���_r���Gݱc57׸����ꋳ�;�E�X�7��Zu��~y��L�IC�D$�T�]�~�%��8����{][��SJ�v��wkWO����Od����j��&e��Q6L�7AClدZ����	Ŋ��U�6E�T����}��9���{�/�m<n|;2�Ve�V���}���"�E����>�x��C��"��/�/Q�5�ԕ�F��D������39ty$�!��{v�
��S4�y�nV��%��^�$��3k$��]ʳm��p�;[�@I�u��Ջwhf�"�I_�F������U�y:������vW�ܤRI�W�k=#��W(z)���;��9.�7x^�}�����+���g�܄�	%}"L��<1�Q��k쏜�j�g��p��> z�97}��m���﹮��6��f�գ��H4�a΅�l��X�*�.�yu�b�(B�`~�������߷��wk����u�38nz˞�מ��n����Cu}��F��'3�<Eҥ7U��e�}�#���m����1М���o�̫v0���WӤ�H��x}��)�fwP�w[�����	���d!����;>�o����ڴ<D��է7�ҿo��Zŕ
������R^nڬ�#<���qB��d�s`}���� 6 ��$����h�`R/��1$�+���g���jp��:P���ڌM��{��v�ݑLT�ۥ�����rwno��nY}���7u��l�q!k{o-�����b����tW�^c��'P!��У&�d�8�6)"�W-����yH��W�M�]����1s�7��p����_�yCy}�H����I�z�]�������5�mA�o]φ�P������t�cީvuÙ_lC�$�"�A�f�"�4e�Mޙr��w��f����J ���N�lĥ���)%���r��=�y\��C�L �K�� $��n�,�o�'{ۂ,�ݲ{�O`�P�K6v�
��B�h�޶0�=f��x`va�
왗�V��6��8��{V�f�Y�����]�IBE"�O/k����r��38�^��u�n�9���_ۻ`�B�\�n��]�ܷ�tt9f&��A&9���58�R�#���5��M�h��6|��U�Qp��W�{��v����OϺdu}�z���
~�Č����E$����m�{�/|=ܾ��r�����o�ON��rE���u�]�rWr��$RJ�"���]����=�ҫu�:���̞�(}�BI_H�����*�s���w���sA��ݽ75/G�Y}�]\���u�ޛ�e�}�%�+��J��س�oq'��mgf�.����o�Ol�� �Cu�g�ԱX'�g����ʨ���g�q
���:�k�vK�o����>�g�\��+8;1Ǜ�*5`�J̄�M��2����+12��x�t(��64vD���מtt�H����TΞ6��8(źl�rU�����H-�����&���`�@L�p�JJ��Q&��3]a�I@wK2�֨Zl`;X�5�a�Ev������2�7�4jk�px��N��v;i3��FZb��%�кB��QL��`�t�pT�Mǩ*��XC��ֈ{a�T�[���*�Hf'�JP�~� :����
�nx%ݫا����h'ϔ:�w;�*�T����!�RJL�sKӱE�2󷥎�g��N:�ƇrI/�ct�{~��7����w�K��7��t�7v���(�/u��_oz��H��<ήW�S=X��]oz9\�����ݠ7kwP��f��}S;��־ݯ�o��5�emt;y��f����m��K}	έy��I>�|$�!�0f߶`ysR�'&��vf��z��y��Wٺ��YX����4�*wT�Ջ*�&���ShG@�E���˴�nN�oQ�㝋q���������_lBE��J�5z��u��L�����]�+(�o�f�D2!$�$Wo�*���5,�N�.�zx��t5n�i؛x$p�Y�۰��R��*?<[Yu�¥�y�A�,=/{��%�X�Wu���==;:�nge��6����'|=5}�I�T��\�)R�y;��?�/��$@I:���Y�ʉ�����2Ysf���P�?�_H��ε~7:yo׫ڄ���QKإ�����B��u��`�&��ҠIU��RJ�H�!$�TyJ��{�n�G�e��������Ε�I�L~�<�ߩ�y=����d��8����&41s�^]՚Z�M�%�6��B�%�C�H����ٝ'f;>Ǯ;���[��Ul�>�C3k��	%s�^����zN@f���ʩ/b���կ��+�1Ż�+}��ݵ�N�;��!$�&�g�N5�9P�?Y�>�UB�q��X4��Hb��y
���Ѷ�̭�W�'6:�hy]�g�Wk��z+/\s��S�|��-Co-�(=�g�n[Z�����mŕ+�9u���Y��*c��6�v9l�VPSv'�ܮH(J�5�t�.u���5����^�
��N��1����4�R7Mu�V�^��3е)ua��(�z�*�I6��L��aL׊������W����������o�-]3��C�W�M�ڭ�����/,��c2Od��^�UK�!4�@�W�/c��obwl�v�V���ܵy��vM5.�t�)�x:�n�Z�e�}�7�Yh��I��m/{P��Fs��s�C"~�/mW�ʳj��VІ���P���ܙ^�'�%��x�����;�4�����ݪ��Tt���.Q�B��t*�ZO�:U��z���p�ML��/i���)ofu��%V7T���Ǫ�d秉|&�ὖ*%�Tuv8�qu����|�ܜ�V.��Ɏ�T�o�;��V��{�=�P+�1o�:nE��p�[������T���尛��w�Ƣ9{rIo^v��fR9�s�r��n���8f�T��B��K�}��kG\��yM���'2-���s=y�0l[0ǃ�m���t=a�T��>�ԓ<*�`7�.�����J��!��3��(��5�.�3��x�b���K/5`4*�����E����e�Q�U���=N�r�P�4��@�s��[mJ9��#ι7��VR�mA������9u���r�Z[t�+O�v�ǯd�����emݒ�� "��A�Y�a�����8�KD)��J$%�egv"I�֣Y��J:&il�9�7:,��㣧4�8)"�����Pt۬�6�"���nB����,�.�tQ�� 9#[I�fr	�m�� [VH6� �;3�(�;�;8��(�b)"��m�e�Gv�˵'.:N�K���:2��֗d�A�u��ufִ�Ӱ��	!;�l��.C��H�Ȉ:�v�i$�$3vWmk4,�f;�8�D��N����B��:e����������\PD�Rq�q�՗b�Fd�;jАm��L�APwE����fqJ�����Bq������\ve�v�2NB��#-q��\f����tQ�fSn�^�y���؎p�����Cڤ�1"�=6��,t=�H;�C��u�'}�vc��z��Wի*�5���o�߫��!$��BGl$Ķ�]�Ra͠-��_mu��E�����V�Ω�K׋e{=^<�$ur��9�%4ٗc!(F�fє�ͣv Jh��V��J�"�+Kn��>�BI_	�%�X;�/���yt}Y�淗�J�H��^�x��j���=@GC6bN�9ِ{1��=� 'I8uΙ�Su�=� �H���{)�uܶ��]o}�}�}�]	�n�ݡ���v�,�9��"�n���}�)ɤ���q��&�r
b����C�[�DXC]	�����yy��G���<N��Zz��.f�MӘ��iˎ�b���
q��td7_J���5�Ω�D2JI6�b��X��$������g6M�}���F$�j�����W$�#֝!@�UU� ��sm�٘����hیn��W�qm�і�o���y��_M���w�%�~�N܅���j�ן	n���D$��罺%��I�F�|��C]`ܾ���յ7n9��M@s��ء�[�h����I@H��)��UN����㵮����>�l�x>��gI �K�(ym�������x˿����$�5r�Zߺ:��㾦�o�{ŝ:���/��I_H�RN��.�yFT�Z;/6���Qt�����t��C"�HKuW�=ՆW�w�4v7W.G��S���
�L���Ya�Z]�5C,��r6�U��V3��Ñʭj-=�vq�&���(��O���ס��j-�#���ԣ�51�h]��䆍�i�d��wm�.A� j���F�r����W�|���ҷj�2�=��PzÒ�N^e�v�����p/A���3΋�`�wD����L�kG&z-�����۠ܧ��]�� s!R��@��[<о`z�Q-5,�K����ݧ�g��3�XJ��CV�,N4�n���f�S￶_��j�E��ƅC"O˯�^�G ��u��:��ґ3�֯�X���<�'��=��O{[��'���M�=�pzp)W+���c��N��$�����7h��g޵����R����K�NIO�]lCw{��E��t=�_7_n�Uם�d�0Z����x���/���t����J���G�UX������q�I���i��s�����Q#E'���@H��P-���������Zג��鋂���e��k����/Nw��l*9��4�C���N9�.C��#�$�m4�@4����-Qk6�U#sj}�_�$��B��b�g��WI}��0m�c��7��ޏ�ù}�RJ�	_�LbՎ�z��n3�=u�L9YKi���@��Vc��JZ�z���Ju��^yF�Q��w�	*��u�[�*e����7�����$�{�&��u���j�L���μ�|+���g�|$BE�ݥ��P��� ����n��?(�rJ~�_9�"���V���y��ʬ�;�H���=����;�Wk���ۺ(��������"�}$�3�*��/s"U:w�;k�x=���1&���7�}>~�{~� ٗ�K�؎!X;bM��D�k�ύ�v��h�U��T(]���D$���Թ=sܕz	$���������O��k��$�J���o��4{�(K�<]��qu�7j?N&����H���(<������D$�?��;��x4�]�
a��[��[���>���ȭ��5���N7��-�8F_{��������^����yͷ� �w{(�IUu����2ܛ�7���$bE"��~s%��>���Ps�mN��~T�����IU��̪��<3{���mn��H��}�p�+�a�iɰ�
��^��"�}�J�ڄ�Eu3]Ǌ�6�}��;��l�Q�֬f
�v�Tj�i׶�yɍ�Z��UwJȴ.�[���t�H���u��l�T�&����Y�%�s[���C����I(T������{>Jw-S���%^��/{�r-��8tj�� �}$��$U0��9d�H��r꣹=]g{b�}�I@{W�)%Hg�m�-�UM���Z�W)��n���_|=+$RE���V���pSs������+5��ܼ�G��ٓ_o�N[�7��8�ޙ�r<�e�g[�jl�*0�k44K-v�Z��W�_n�"J!��=�]~ɠn����Z�v��O���הfN�ᖆ�W� $�|K�v�AR�{�.��<Q�Z�;���s-8^�=n4���[{j!�m/]x}���)%}"�'�U�ޫ[�gk�W?o�0r	�� n!�!$��L-v;ꮍ,�|�����]3�{�\���|��Nz����!<����@H��/\�1)��5�hյ��W�]���xe��ޕ"�E$���6gz��z�܆�~ݕ��9]=�c�麉�V(�U���d� $���J�y^�:}]�:%ٝ��s��d�\=+��_݃�z�G*���c���k�w-U���+/[�/�Q9D�C{�5B��y�<]CZt�J��Q۸,�m+[�n��./_��u����O�p��n�u�'�ָ[�����$�@�[��kx�<X��V|�!�a�l���m�C,��"�tV�\�qY��^Q��0�v�wWT��a�;[�h��0��sۗ3���#q��-��t�iz̓����
��&v�H$�T��8�155Jc��+�[+U�,CM��n,q��}������]�!��[@w7�t�#_���?��iqh=e��ФX옲RGA����ct�٬��&� �b�5j��~�<�@I(=���_/_��d��9�{����7�gپ](	�P!��^w;�ٽC᜾2{.���z�I����ݒ��H��0��za�U�y ���ջ_n�J�:� �;c��Ouu�I�<ڹ;��|�|;T���H��ӱ���h����%��{[��N�8̒�u��.�Y��{������CsP�ݽ�甩Ë�<<2��7�����6i��}7P��큻�=�|1����'���ɮw-k�@���q�y���^��2 ��g1���]����������I.{s�]Η=<�\�����Wm�ߵ`������_�I_p�����v-j���A{j]��q�SW������73̱��e���As����q7Uv{���r
�ʺ��O+�!"M�:����̇1������|q�'����=�y���I�	u��R*��/�_G�V�n�w��堓�*�n3t�{z��{o��IC�%�%	�Ȏ��e{��}�Cv�ǒ]�����ݓN�|�,9�gK�rʢ�z�J� $�?��/=�.���ݬ��έ�xӶ\�/<2���E#�|c����<.�!�n�rWM�8�%bg0)8�;f����)�T�;Y��g��ܤ���M�v�w�W�v��Ӗ����1�$�$R!�6T��yH��܎��oݰz��_�_�$����Ǻ�%�|���I,	&��UW���^�$[NM�w+������Y|&�7v{G��Pn��̱u���>�V՛��m�5Y�O�*�m�vw���N_�:��䔖��8oK�}��=#�	%}��Ã��N1���_-�xn�};�=�c��=�2��G�Q�-�oz��H��J
�G������uv�o�����s�hGBI_It�z�ڄ���BꮊV�&�:����M���u:���Kq+Yt%�YI���}��'�g� ��}��T��U\u8oe����򳓕���!$�$MU�a�X�����:{^��wu�f�s�_s��H�y��x�[��;���P� $�v�N珶�S�/{J���g}q}ڤ��H�����N_`8�0N@w/�����RS�i]�������/6{�o��fb��r/x���cP9�]s,���;��n����s��Iί�={3�1wR�E��R�^>Rz�[�R�����t����3Kw�b�$�$R/��Ǵ��i�V�d ��=�⮳Ϻ�׳w9�_j�}2+U��|�ǧ��ե,ݞ�71y�\�Q�]*�V[W�[�7uh,t[�u�ZOC̝����O'��3Wn9�^s?{}�|(!�>�C��W� $C�%|���%}0��|&o��[�b�n��f]�����I��R�m��K˅�O?�P�I#T9�P��
y{����:uw�������fmڤ_I(H��^��嬆\À{b��v��&'�����8\@�N���y���2���m��E2W�J��^�̋�˚o���}�U�݌˿x;@f���)4�KW��rA!�,�;3��nu]�;��V[4����;�r�En�'ne
�Ɵ{�v$�����z�%R��j�5}.�c-˼O勞�+l�1�}z�k�VЬ��Uu�n�c����5X�y�������Pwx���ǛM>�vkT���/��Q:��e�,=�Z%�;��6(����\�����V�k�M��R�ٶ0�֢*2	��X�,�"ծ��ӪnH1��,����}Me������JEkܪ�1�Ϭ�bm�|�n��j�r�)U��Ox7�bg��#�[/�z."��*n���;��WI�{.�	�rbB�g���uaK)�m�ۧ��/��,f{�g�/Z�T�஌�>��,7iů��iu�Z|wB���b�U�o�1�=h�ƌ㘮�%�6I������L2��2���e;��Y��u�zn�(�]+��U���(�N3��&c��Q����eu�G�A�ɣz�|��V�F�#�P��s�^�7�1N�Um�Tp��F�!��ꑪ� �iaV�`�&�=����A::.t�SE��2�h�']<��r�]��²<]Ńg���2��M���/G��wV��wf�Z���"��h��/E}�pUsx���n��q�,��Ƿ4֬��;�sDu�|������TgNq��Ý+'�yVq��ZM�q�M�3�g,���i轎����tO"N�a6��o�� 5f�@�_��Q&�,Q�c%���SW-n.��U`Ѹ�,c�U�!B�g����@˖��iR�s�7�Wn�p�;�_�'35-���g����9���eӑ���6�� �B
D�+kE	m�lm�:���+H�:'.��B�2���FVm�Γ���,㨲��;��N�θ��%��Ř�'A���Z�����⹵�Am�9*&�q��'Rq��'�%`ڎ�m��ȻmvV\%ڳ�r��.#�����8�(�8�����B��ʲˊ(���m���d��*��B�"��:��
. �qTtN1����㣓�q.��"�*����GQӔ��THRt�M��"8�1�D�eۤ���qD[nDR�"�z[ Ym���H}}� nFmW-�&���!�	tJ���ٴ�ܖ6(wTg�IX�/�#��^<������6'�;cϊ1mg��+�V��W+�Ř5�A��n�0�-t�=���t��������]nH6���q�'�e�(�ժ��mYy�A��*�mM�!�f��b[��[�xڶL��T�ˁ3�\�D2B�Y����9S����cY�fv�y�������'voM�AG�-���(7L�e�Ύ��.y�fh�u���6^m�^8o
ڶ8s���u�pՆj�k�#� ��+����a�L�5�TF���D��In��P�NUM��'���X=u����3��X@4��� 
	tg�],���6M.M��\YV��i�0Me���2�X�=�!N���j��Ln�э�������9���ˢ�vx����̀�!��p�h���s����w$�m�9Kj@��+�3+���y,�_#v9�f�. ,Ե����J�[+鑡H6�A�u�ӟhx`�x�z�;�Mn�,�u��� lOs�8��ȓu66�R��H�u�Z]E�&��MQ3�h�u�m��#�&���c�u�!�lA��-q�ٓ=��k1v�<5�:SQ�m��ۛ���	(�9ے��y. �ʜ�i�&|U{xf�ݐ����S��wma�;c`��N 1v� ��kM5*]���PGm�ղX˄)cv�IA�&�h`;Yqe���ڋt!I-E��{%��[�Ӫ�:)gA�WW"�RJ�lP��8x��q�].�6cZ8��"��E�,v(^��T8{B�u�yۇH���:y�t��Xfn	��(��[-�фq1h���(d*�ci����z��207n4O=:8y���Y��mY�lҚS#��n�`�R�o	tm��".6���Iv�-�ɫ�2;^�ׂ.\��[S��Y�L����hS�b�4�09oVӶ���=[M��on*�z�ua�k�R��)��XѬ=�Mť��`���1U�7N����Яf��Vm��)%���ɓ(��L7��e�]]�ĺ�ճ�K�P:�C�x���n�kY�\u&7S�Iw��X���w]��)����mv��ヮ��Z�6<Y�7c��Grf{��Qx㖤'l�a��'�
��	e0�[�m܈z�9��T��&���.1�]���D�ҭ�����U���K���/Md�����)�yG�A�mi��а�ժ\���z$��I*D:�4,r�{َ����{�7̰����c߅��BIR $B8`�iV��ו��2W���re�C��:�m����!�j�K=5٧���m�z�J�H��$�g�Z����c�=�7v$�=v����$_	���������[�:�k�1��-�y����������g���ϯ+Y� u	$��J�@�rҪ�?����}�%{�U�����m�$��f`k3{r���(`� ��/����{`�������j�n&)�˶"�2�`������O_I��>����1��λ����~ዺ��pI+5}$��"�;U~ �'طW��rn�\*�]��z��}�Z�d�@�h�vե���w�&���P{wś}����4;̳oL���׳U����1��r���]�H-ڬ�ZC�)�@f����$��&]�M�;=E��Ƿ�>3o�����_� j�P��&�OS����A:���s|�L;�U�Y�p��ha�Z�V�|&�$�$R!$c�Xw���q%&�j9������w8��ݿ����ϝGA:��S7��ٚ�d�c�����z�5��d��r�՛D��+@~_fБ}&O~��}�s>Z���v��ux�ۛQ=����v�ݡ���H]�jx�/�(Ƈ�1�ONWj���.��z��7n.����JVD#o�ݨ	����i�t��}hF���X���dv�@�)FR��Z�P�U�{w7��� C�j�R=۽{��;�39�V�8n��3*������-��ۙC��$_I$#�)��T|�`;cL��v��Z�ʛ��x9�����{����%	n�Β��L�n�+gCȹs�~�Wufgi���H�Q�|�W�|=��&A�� /e��I�T���1;<�������l�j!�)�I[]�y}�BI_H�[�:!����{:��6�4��5�Sy_�}���F$\sך�����=���r�������v�$=��[6�c_ޡ"Ȥ�{�5�s����꺻S���~��N��"I@{�B���
�ݴ$C��:!����t;��=��Y��jz
Pp�g���i�uS��yF��!Z�V����S.��{Ut�	�c��اU��ꂥ]9�I,<y�=Z�]z�x=_=��_	%H;��[���]<yYz�*��˛����)�IBG���Oy�]�=ߖ�<Rl�n׉^���ɹ��λr�������F��HU��>���tR!$�l���le˯n���ޟ,s�|7k��@n�V�yp]G+�=鞮�1�}%;��Ɲ���٥�w�x�t7z���gי�5��5� $�1%(h��-���+�L������h���w��|�r�I@H�ݠ����K��=��n�z�A�ʮ�le�^����8����ܡ�pͯ��G"�I'qcYϸ����gg{e�oC��s+��$C�%�P�#K��-�2�N�P^4��a��]�u��G�=ޠ�|�}�u�;O|�k�ئ�L0�����X���]r'������vl+<f�xм����P��:���lv���3���&�cXi��[&͟���ǆ��w"������.���hnʉ���4������!�0l��qɭr�>;=�"�N)���v�j����KGG0.uV���e���@a0aT0�bm.�JǱ-���-���^yjޮ4rs���ݥ�`���M�鬱�Zf��:$f=��ԭ��8�&�΄�]F�PSm3�K&HJ���c[�v&f��&`{��q�H�/�j��o��dy�γ����{�����[n@$@H��P^}��n�U��d������򻪝�k��h}$Cu�R�g���@�7ww�u����R�նO�|��9���<�#�7hI$xf�U��y����b�D2�l����b��`�Yv�r����3�X�P!%��[��=�b�&����/U�V�;\��m|$��K���2�_����ٯ�\x��f����7Y��KZ�#�,�&t!rio*$B*�DR��UJ��q���$_.�l�;2s�X斧���;|'���{�وw��P!&�	|2��]���|9�W4Q����˺�eA}��^�/
ɹ�!���۸d\22A٧h�}�֗aO(�(>�n���5����"�o)��|<̹������	#��˯N��Z���"�D�Z˴��ӾO8G\��85�^��W���h�@b�����ϱ:z�۴��d����mc�Z���'n[~���:�öP�	����m�s.��'�kC���z�[����o,��$����%~��Aq5��G�{r�����N^�qW��7v[�q���J�9��z�Օ����:���C�n:���i'�+��Y�9��@n���rU�s r���N��9��5����H��ګ��|�%k�IR/�ە�]8wƳSe{��i)+��\oyٖ�Y�N�����Wvk������r��R��k1��XpU�K�efV�<�I| �7yg�("��Jߚ���f������p�cs��_�q}<���	���إ�b*Jn��g-�0��)85�O�^'T.�^o�;W��I+��A�)Uz���gx�'v�N�{nr�x����$��o�N���mRn�wVj�j�\t�������?M���;B͜�Dx�GK͢[3�n �hH��~��WV��2���~뗵��\��&J)�P����SʹS*��B�sC}��ڄγI��D�/�N���I^��������y	J�I}N+q\���X�H�'�vw�n^���y_r�$�ը_����|_�;��ݯ�oulU$�69�|>�z�񡵷`���MV;ȣ�z'��S����������[4����;v�bQB��+afx{�fcx#��v�:���u2���
�4[w������zP�5	�J/��cl�uQ��J�3�ڀγV�֥{��؆���w��^���΁-/��Kh����:n��u�����d�m�\��vĨ���{������{�����A�������m��_	F��}�D����j�IBD$^��PDM.a������������+�=���[sO-k�}��ڐ�I+�" $����)ogT�M��ZK5njW���vn���$��=Ī�&T!���W�!]�i3���wx��/��؆!���̼�3�Z�vm	/��G�嘇�+1p�!�g������+�졽_n��w�Z}���̕Y��mi+Ëp��9���*μ���3o���=�B����Q�'s٫�+++e���t㋫���AƴU��������Ix�A"
F�n2r�h��ҵ�Ӎ ����%cfcC+�k`vv��F�Z�6&��c�W`Q�!���n�$�s�eZ@ʊ
\f����ݘ����8^(lIP�:a��b[^v�'V��']p�6x�j�q�4x�lƭ[D�^��u�"ⳗ��m���%���D񻪭��p�h%jd���[&e�=j˝X�{�o�߲G&��3)�ݭԛ�kcj��h�5�6�M�Aj��t*|6e}�|$�8��qN��^��x�~�+�3��܋�nT�$�$�o]5/Vf�6!o�Y;�������<��=׹�#b���������p�]2uX���sts52v�����P!" ��>ڑd����z�e�KI(G���8.�{���~��?-�W�=�^��:)%}"D$�v��H�� �c�_<�u�s����'�<��:�����b@�o�o�X1$8Z���1��@*JEG�X4/(���_l��}"���0<�͚���z��=�{����� $BI_Z�).tG�+����c^A��uYLJ�$��l��1ׅ*qm�rE(zk33J�ME)e.Q�7K�t�^(duKۚ��Y��%|H��$�Tf��V�3y?���T�P:v&JQ��W�5"�W�C�;��7�2�	�"�G�y�;��s+ھ�	%H�����!��y���7h��S6WY�f�.ｕ;��ӓ�\-no{�E�P)�<��]�Æn�����}Ś��'	�+�eN�E���w��/�b�.3�#�AV.�L˩Y7Wie"ƕ�&�@!1F<g�`�a��<���:�b脒��/���r�G���� ���\��2���ww�v�.���j�<�y� N��OK��F�69�|���RG��O�҂D-�:P�E"�d@��8j��;��*�Ž��Y6�����޺��#V��IG�2lݕQmEY�=n�.��cxgWC�*[c6��)ybP�YU��Ij{,���|�׏v�Y��f%q�M'����+�P_L�Rp_�O��h�W�$ԂXۃ�c����Z6�8����U�+��-��f��b�v��J�v՞��YC*fSk�'2�vt��դ�����y�ot�f�:�`����>��yU���-�Aֿ��r�N���gK��ҭ��f���Ы��,��*�6�ob�ŹohQ�7��/�k�/3�tގ�{�tv&��C1gT���W�6m��LET#Xc��ienV��M����Ud��K���7U(�f�9��rv�Z�ܬ*���9�ѡpe�ǖ��+fH,�������e+�m?WR�qPV��]PE�旪�Ѥ�̸]��N!W�Tk�Շ_K����O@�Z�����t`۲.���>�K��})cVk��M�ɔ����V�]��{�U(�+i�ك��kB��{���j��K�jY���B]�t��CC]U"�w�b��֥[5�8
Ǆ>�Brr�H<T�6���7�qUf,�[��w���:u��ӝ�.�䤷jq3��m��F�«�Z�W�O(*f��.ΆȰ�� �WR"[�.��B�5����{7n�D���p$�`�Fz�c�Xŝ�:�1�D���]��vVWb6��S[[�˥Nð��*U���J��S(UВ���-G,�O=���H{�w��CR(GJ�����*��	'yx��>�:��o���U�ȗG[�mgևP�fQ9�E�PD8Egu�wf w�%[n��;��,�I.�����u�m�(��;��8�.Y�:m��f\EXZZ��t�Gu�s��ܒ��$�4q�6�Q*.I[Y��DF�9á��IЉ�ۉ;.�9!�a���s�(�)
;�P8�8����Շkklt�9��j$mݐr%�Rf�v�2���������;m	���j8�@�)�1:���쓹��kqݝ�q��p!�'B'8�Dq�Z:�98��l�!��fPt�@Prr6�-4�:)�fqDQG᝔ts�BF�"r+mQ�\�vQ[�C�������乆j
N����;�DC�Q�P ���R��_j��h0Ar�����k<�����d4M��>8W�c�c���ǈ�_/��dU�"�P�2-���;u����{O���L�/�����6~�P���~�aTܿ��g��b�Ĕ���x��<e���kە����]�74����s�gB�^ha� � ��/����c�}��]E8]9�������OtZۯ��@���7;��qshѼ\�GǊc��83���-�A�D��A�#wf���;_?� 2'��T"J�����%��w}s�����]��osc�
��(/�;�Q� �%#��}I94�W-*z�4h��r���N���v��J�)�ښ���W|F�uK��f"��C*���̍����Spm�c���n�s��Ҟfe����W����}ǟhpYݽ��5�Mf�8�)��6�T9�kj���L��0�d@P������=�h#;C����9��=4M�� ��D{P1_C}�=T��)p\�]%f��ml��ŰR��kl<�s��]��o^�Fln�������Am"�d/��#��-��꾿Qs'o1F�Ϫ���%tП�A�(���n�GN�E�|Wh�G��eAdw����C}�_��� mMX���� �@ȵ��_c��z��8/���D�Q� �%�[�]JQ��Q����&�_x�@��4/��0����[{A�o~��|�x�u� �wi}�!#�W/���nxY�	�PD��]R���yL@ܯ�j�7R��D�� ����R�pV��{o�oP�y��|[0R�6�,��AܤA;( wiN�D�i�i�y3ݕ����y3u�����:o�?t���F����E�.K�M�{�/v���_���	w�2��nҘ�t�z��z/5��ZO��K�ƥ$��tK��
�[+{���m-0��O������G��/WjM⸱Ѽ�M��;�P����ܺ�oc�Am<jNۣ�k"�0�q��/�Hq��\[�j�O�"<͓C�7&��;�l�nѓ�C��tɴ�l��z&�zn��v���gi�,:N�j�B�fQs[5�/qbpֺ"���PuǊ�7��w'��g�p_������?n���Kt��s��bcr�ݮyg&�A�5ɡTV����uuZg{�X���q喜�K�� o u�����ن扼���/z����ws�X���e��X\^r�yʶn��K)l�ǽ__W�����G��w�9����P%�y"��/��Y�ݗYac�*�9�sw�q7me2��o}Q�)G���+� �)�q�� Ȩ#Yz���lW��A,��#u}{�����=��3��Y�DY��g^���v��}��Q�}_|AB(n�A$����J���$��~�U9����~�Q�_C�	(c�H.z�Q�5waO�YWT��P�:7/;��P�(श<�CpO?�� AӇ�5���kH[����HxT���ŕ�EW	zż.�*�J��@�"���D(���4=�aR�����Yi�vy�Ak�'�Oi�p\�1#"������伻<�㝊��a�&��p��I5��(C�fZ�P��
 ���������=W4d���
��4���ޛ%�������'�Q�(Ⱦ�dGk�8�AW���0>*�>�}�*�Ľ��7¾�PD�Fk�$B����M����⏘��L�Gr|F֑��=漢���sWA�R#�����K+8�sk��U��d@T��0�YY�y{�~	�|���b<:�f����8QsA�_-�#�c�c{}Fj	%��1Ϸ%�
�	t�;c5�%�@ӌv{s�:��۝�m���k�Ȍs�X&>K�9V"�g�#�W˒��{<<o�{��d���T<D3��ϙ���Ӝ�b<x����|8���7����E9�}����ŷ�X��x�b�(ȷ����e/�(�'|�~���A��������em��~�q1�D�Ŵ*U�Z�ұס��{��邯��ұ���K��S#3Z9SeD�H�PԖ�-]
)�c���ƌz����o��mM�8?/�:G_��E��U��v��<��3�P;�dPr�ȼ�ʜ鳘f� �B�����Y+_i��P"J�~[�"7`V{���#gN���p1�j��b��⯈1q�� �"UI_�7��_<������9�͚Q��D�nucyW�����SE%�(KK����#6=O+g���e�����?1%}=Wޱ���K]�C,g{�1=��0��@w�|b�PE@���TϬ/7ӏ��A�S��ȼ�ʜٳ�f����B�>��w�eP�_�Zݖ&n�c�6��Ybs�,�q=��nwq[�MU����[;ꃸ������ ��ꋈ�"�AE_"�j���79�P�A�A�#u�z3s�La�}{SG�/�t�F3KUn��&[��n�d��0�Ui�s�������R��"j����ȷ��P��u#0+[*^�1ɕ�z�A�+�1
�ǈ�_W�|E2/�(Bv��d�����B���]X9{^��߾@�^ +�B�0�@�%}�θ%���)��c�WlAA���yI�a�n�v�s)[\SZ��hum�i�9���_��7q"�9�l��F�r��b����i�j�!�"�EG���2!@�~�ߥ�*]o���=C�ŔA��[f��y��>���Ӑ'�J ���m�]i�Dd_C�/�2.�0��=F���-X=Nl��� K�(��_aD�#u|�6��4Y�A�����嵤/k�O�0N��OL9\~���sCS\�8��R"�/��E@�e2!DH�4(y0��Z�i��X�ѯw׋�|��0��m
"J��"(E(N�:�����-餵cw��T�ҩ�����8D4S)�l�g.�y˭��g*��-���QN�[�T����J��5ھ=�CJQ�IZ�<��,� SS�l�rGI�#zn��9.����ѕm�]�+l/��⸇&O\�s,Ƴ������,!�BQD�h:�؈G�[h^�:�'����Gv^a9�a�����K%�
�8�9�܈�k�v[�N`���o,��P[5ǔ��V��usq��mh�U��N �c����d�����5)��֓y�����6\]��F͟��~}����J��5���򻙱T��:���N��㜨��ŧ� �Oƿ٩���͛��7����Î񱼄 ��@��D$�@"a��M��V�6��_n��.�on�>0N��^�r��ڠD<~�b7�↕��q�	�@T�(a�$B�ɯ1^��:ƮǆW�\��~n^T����G4����dU�2�^�M�k� E��QȨ{Eq�Y��sf�0��	x� F��7|�î���D� F��:W���n��5��7���'ל�L9@+��B����Hg��Vy_�L�"�E��YJ��VMUY�9���p�J�/a��s����%5��~�~��#��ӥwP@��`���L?>��h��/�-��1�t�D���/��+�"��&D�T5�q��K�����sc�)��0vIU�%eY�-@�8�p��7���S�9�;�H˝�r��뎻/[�t��ͽHb9/���p ����:�z_��������dp�Ay���:p��k�C������(�(W�E�=zoO�6y���#���k;��,^ �mP �\~�2	ݤF�_

��4�7���w�����
[�����N{����Y����L�Ļͼ"��դW�E@��Q�dJ��+ι`�ֳ�(o��q�S�79�o��^��X(G�K�ͻO�vG����A=v�Om��p��6�ը�L��A�[Hv3�m%���}����MA7P_�#s����Z���&�h�J���yq��s"��H��E@�dU��_H��w]�;�Ӊz����|�?G��^�f.ǮϷ�5M�8���sA�Σ{�qyՐ�JDyQ��QȄ��Ӷ��ig��a*�i���>��늅f��;+{i�nA�h�SΚ�+!ڪ��7�]Ppu`�i�	���ProQӤ򦍻���w]y7w9�o��+�Gj0�"�(Pgܳ��|��� �eF��?mis;_��b�.nW�� k��q�6�4aU��՟=���P�
��|a�tY��꒧;� � z��vf˯od�4^��G�
"J����{g�>�+��۸ʔ/�Xs�:�6�7f�7nX[[v�����q�H!j�"�h �����(|AE]�Xص;�.Y���7�<Q~oɌ�}A�~�t��#u�����ҁ����%��6�df��Jd!��_����S�:�4׈ j�8��2.����j_:�U4� A�B�2W��ȑx���o���}IM�6��\���]�b��qvˉ�\���%�9V'u��/ݮ�u���ȡ�T?��Ե?w�,��O#���X�yu?E�W��-��n��f�{i��{��ހ��N��Z�>���}R�� �zák�ѽ^�6���[�M,�%���3�ge� �z��}0�%
���:�����R�����ݻ��su��]���ڠF"����DY���_c�/�_'����:l[�m�v��'�rh��p��퇣ZYiY�]q�nO'��K}�#g��GN����;~�W۵��T�����/!��aG�|;�D>��֐��|�ب~��1ь�֙�r��=|����VM���/�|�_v���P�N�Я��!�a�n�7}���ir�H�=��
�nM�UmK�M�]pDu���~�KyʴG���.���oT��x_]eP<�<Y@��㷸�7y�b�uʘr���UcdoG{ �l��Ι�Ղź_C�B��>�Rt��g����kU}�`�ħ5ՙ.m�pDw��Ўv�x��9��BB��D��	'�!!!I�RBB��	O�$$ I?�!!I��BB��$���$��$$ I?�HH@��BB�Ą�	%$��!!I�		O�HH@��BB���$�萐�$��	NI	O�����)����t�柬�8(���1�                                      0  ��                                   � ��H��IQEJ��J��(U(�"�UTRP��*���U *�@�I(�R$�����ER�T���  ВE*%$J*T%Q �W;�HR�n�	W!�R�v�}i�<zR�z�v�Ugw/YT�l�R�o'vRA窔�t
Ww8U*��J    �   Yҽ�:Uݎ�R����
WvtP�n�PU�p�9��[�J��%Hݎ��Y��EV��     =�  ��U*�JJ��URO|B��u�W#!H�c�QGw)T��*���{jW��yZ�Ms�
E�R���*D�<�T9�J��D�K�ܡE  P�  v�_}�zT�OT(G��'w��UyhJ�{�T���yU(��UP��I�G�	;�tx�

��Ul�� ��X���tR�*�   |  �ԐJ��P�T�H(TBM�QJ+�n��)O&�WL*[��E<̮���Dg��J�4��B��G6*�nD$㒻��Em
  >   }���>��l�8�T��5E�J]�	w��pD��6H0b��������      ;�)IP(* �$D� ^���AVa�m&lr����w�kR�k�Q/{�б�;��B�7�c���{���{�@  �  6�{�p��B�C8�]������{����=�� �{m�*�
��QU�t��j���^�*������;��O`   h>  �UTJ�UJ��yJ�� h�(Q��_lr�U1�gA#w��Z��]
���R���QUCrQ*��m��wT�.����  @=� �q긌�
��r�TOz��/{�4��n�QS�ܡB���J �Z��Q��ʪ���(W��xQ�W6H�c�WPS����@h����IJ�� �4�j��Tb0 �a��T4J� 24 %?R��h�`` j��*U7�F�hzj�������U�O�$����������_�����?~�I!!I������$�@�HHRBB��I	O�$$ I� {��������r?h����q���;��.�$W���h9	6f�G2]jØ�:��T��ΦE��T�.�B�*M�6��:J�V�Ǫ\�?U)���¸���I;f�VL�{�o��ꉱB��^��8��B�x�Z?�t�3-�e%�U���g��ifk�"�5�Zyw��'iȭe�u{q��Jt�q��:��Un��[T�	֩j�dL݆����7�7r�׎
�rL7��$ �Pb8�-�Oou^SnI��=9�/-�5�(���6�&�2�+1V|��+Aک�YB��${�7�G72�f��n�r�գ1�d�Ui��Bv�yzDZ/r"��t�kV��h�6{��+y`�v�bǋj�V̭�/\�Y��%iR��EnEon�[�&��Uf��~��!�6k�7A5�4,�A#g)J�
��bՙ�.��1l��U)`�GN�&toE��5=x���K�����h�vX�yn��U�`��i�e�E�r�RAA�EHk'03.E���E���:���[�w�/M�5��{Q52�����B=�	�Y�r�����U���Fe<���-짪ӥX����������me]�U.T�Dâ���t^��"Sۚ���l"�DF��l���[nL�B��ј$��M��7�-ԣ&L/�,�H���Ъ!(����Vl����a�N�rи����
ަ�a��F����jW��!��N���G7�W�j�עfKB��/MT
5Z��b�VP��O4`�usVVo��r�V'DVEHݱ.1���Q	b�c��z���*�+j3e
əf0$2�LdŹ,P��JZFi7�ֵ:��oDL75;Ǡ�sI[�ފ
�QB�0�V(�t�P�R:�f��j��fI&��I�"�b��[��J�QdUf����0��I,,�6\7ym���H��,r�`O�C�*�R���ڦ����)��oi��[�V��.����𭨑��M�d�5S�����bh,ʷ2�X&�m�72�5m]f�3&�3E��U�+e+�Bn����J���f�MT�ɕYN������^�Ж��Ùw�D
�V��v��;��c�E�����[�˦!xomn�T9Y�1ӊ��U��M��wu�j����M�ysl��C��7y�˳��V�����UW��Q�VF��ii�ZZ{�*�f
��Xs�h���t���Eh��^3��XSSji�q��˰�*�:�ki
�[8�\C���.o�U*�:7�`T%L�����ջ�"�@��*��4є�b���6/ ��f���dL[�ڃ>��Uz]�t'cM��,��ݰUK
���E�����mP̹zIU{Ml�z��%2J�M���z�_8��Nw|�*T����o���ъ����ީ��Y������7Hsv�cM%��=`޻3$�p��1iXAڒa9&-��Rff3h�Փn���P��\Zwm�4V��͘��J��V��+73�ݴ�*��-P˱��l�i9�	�W2����64�3t֩��Y'rȭ�CV�'f�.���5��]�%
Yx��*��L��ڡpͱ�V�����UMm,"5EnA.��S,Y[mnܷ�N�)]%Zj̖�^��Z�^�oFm��)X���m&VfQҪ���qQ�5M�Khn�w��U����ܧ�)Y+̦	VC��n�n�q�rY��õ�/�4����H�,hzu�Upح�Y9l�Cv��ڪ	�kH��YcnD�Ԗ'OT�v�e�MK�.�P�6�]ńeL֛��9��˹���JeK�r�dǙ����O�r�+h�kiaɮ���hǛE]J�J���T���U2���*�+3e����U��ri�+
ڛ�-��=���į&VVh[�T!��Y�if!e��77C{ǃ��X�"ˢc�/rɤ+3����fP�E�Sé1����]�����9�֞c����Z���59���PYyzB�F[��nU�Tse�����6�3 r�M�dV"���V���l�E��pЧH�Q�*7�6m�T�g̲oC��
��t1iկw0jӷ��%V���.��(�7��n��n���rA�5��	�X�B�(e�;R����O������w��Q'a��q�rU8�*�R����Ap��QS
[JHx�&G�}�-��wq� �ʵ[{E֡o`���5W��ެV&8�V�"]�hqVn^S-b��X��b��Jn�#�GT���bM�s�ƣXP��*��݊�2���Le�L�4�#M^q��c���[��i@�ҬSw&Q�b�n��,i�7�dL����P�h�)\9�̷�(�@��е.�[9�aǯ�kpIYug�Yzv�J��$
ʽùZ���FY��	�(�,��k�W�ͼ��l�b-:��^<�m\��q0�j���D'���y0�Ν2�!0�ݓ�7-��r�;�.�%`�u6����%Lі]�a�&���7C�n'ASt�9%��uj��5$f�T�3>�He���q�ZX�)�)��Px,���n�Z��un�'���ͳ(�T��;wr^�1^�Sj�:��w�U�kaU�!F�l�Z�c��x����[���˧mc`��� ���3��k*	T!V6a�k���#"��*xi"�Y7%T��b�06��L*Ä�=W���٦�6�0���W�'nj�Ż,+���f��ҁ��2ݗAYD�+-n$Dȡ��缭E������V�f�3�{�	�tZÒ���m�&��V2�zn�&��Y�jD��+f%��P�9sHYbVf�����������)��Qݕ�؁h�S��8���Z{f��#zն����bv�cͥ�EyaY{��jjd�Uj���nn�u3f�niP�/Cm�$̙�(UkT\F��t~Z�B��bN���kJ��Z�4[C%��n����kn�K!�c%�W��N�����Ӕj�7H�ԫ.17{d�CѢ�U7��Ź��oe	/i�6w���ܿ��]����Um�Q�Ⱥt������N+;3%<��vر�F�En�n�I��n���^]�:��7awd�2���I���gZv�BeGFKcf����`�Cm�m���"5�r$l��7,M�nڬ�	,���V�ؾ��9�/�;U4���෵#Ъi�6�j#.cH��Zű`�YI<گ����U]G[�
1���i5��Jw�L":�2����2�0\�6$6��+��,�����JlXu�]�i��I7s�K˫FL4��.�JV��#v�լ�sM��&r^��c5��vs�F�xBՑͣ�CtZXxT���)T�D�BT�V�G�G�A^�]���nV�q˴����N9�*�q[��گ��{V�uo49N�Y�ut�5���a�ݭ�:�J�NUr`Ҫ����y�cl^��ԧ7���dsBt�[W���Y�T���ZfL�k����Б���{�y�Xh�L��w&�kF��w2R��w���c$?�N��.�^�p�ݽ�wrV��z҈J
l�t�f��EO�7��^�*-1��o7LwKu���W�M�M�GT�Wf��аn��O�Te�oղ'�ksv��d�;WHX���Ԁ��b:v�#�(��P:W��n�!��[��j��t�[���'�@�DƪYF�W�F�+:k�Ɍ�V/���7�����^��R���ead�j�sm,�^�NV[��J�w��uNVRG"b�Ҷc�����hM���Z�%nb����F9Nͭ����[!�&/�
ZX[I��+a�U���Ņ
��R�%�T�o2�EU�wzw��Re��`�z2䱗a�(͸֥Q��v̡�������3.l)mkۣ.�i��tF�	��?h�ĖT�I&�s�D��j^���8�7x*:�*ŵT�[�5U��e�Լ5�[��ٗ[�.]k��
ܛl�{�w�wNV�:A�w6�*�j��Y�75�Ԝ���#/ku��ϲֺߛ0��[�6��9pK-˘u]	y�OF`�Hv�Kd��N��Un�4Y�y��Չ[R��R*ãAi��V��:Z�pa1mF�-d]�.�N��K(�KŊd�W�ONM�Y����GM�&	��D�
TWicx�l]a��]ѻ?^��LDf�c-�s[�2�h�{�K�E�sv�n),*ˌ֚ٴ軹z�-XE�R�ʙ�E�iE�I<WOH�����X��+v��p��7��wRD�ʧZ�͸X�^��@MF�ù1DB�Y�����Q�wnB\��Ct�W]^��]D���זr��s	`�D1���Sӂ�ޜVt�UXE74m��v�V~��[�u�U�֦;š$�M�1	�h�t�
����ƭY32�!w�'2͌ϲ�ڤňB�eĤ*:��L��r�P���`ʹwGfK�F�e6�m#G�Mn�$։�y���
���&�-�e�F����2SUDm��`��ףvK�"��SL���V;	�45��L����c4l=�C%|�
���	G5,2^`�����&�2h,���-�gd*� �ԅڭ׵KC��C�FmY��:N��7VI�*�.
�ܺA�7�-c�W�&�"c<6�P)AQ��sk0��#N,��i�b��UÔN��>�˺�K	�c\0�Mf�
eUf�/5���x^ř��PQʨ�h�*���mA��U��6Z�ࡖwS��Tr��r���j����v�ۺx�TȬ(��U���n+��%I��vw+wm��3�w�/a�ң��ӵN�#2RW	��ܫ�����T�֙xBɑ����5S��l�3ǐ񚸷C�����y[2�����vwt&��p$2�'Z54A���d��f��o�9@�Q�Ӥ�C�r���l:���X�.
��4L��KT��Cǭ˫-J�ۻB��Ut��R�6�U����2�c��w��i�9zFQ�Z`�4�&h�}J
�.�X������X_YN�Gz���L:5N�⢨\6$�%�-)4�{�ݭ41c�Zۼ��ʭ7�Z�c+ScZ�٩�F�ڽU�n�e*��]�];�������t~�CV:J�Y��Q��N���S6�.2Y�k]k6�ƂK�*�=���ա[A��P���5�0�S�>z!%Y�t��ȬȒ��1^\���c�̔�
�kPWf��u�WJ�R*�ǏkV��d�WU1��oNnE������6�Ѹ����`�2�EUlV�'��Sj���cr0-����&+P:t&6����_M��Le
Kn֗,�L�q��m�1�u���H�#R�&5�U�B0X'&^D��o�zb���P��-*�nT�3*͕l'���,�/U'YfZe\�S�D�Äh����cT��-�әJ�5-W�J�ŅHͫ�*��,c����7Y�W[�m�,IG�NnU��'m�g[B�l��Q�&����N�h��a��e�9�&ͥ����@����Q�;-��V)�ܷ�fKM)%ѓ�y�#a!�oѻsn	��,�Z5�bf�T��������wj�J��4�")�j���Zj�-@�L��M�;����Aޔ�U�Ux,Vչw��nd��v�T��3TDT�y�ؽ�,�j^���Q{��UP۱���o���yM�*))ֵL�`��k廷�o�*��/T#uEt�P��Um�˸�T�;W#V.��x��m]l��c��̠ۭ��,�lӭ�v=�� �r0h�fF�)�*�,��+=v]�tv�겆uҋfA5�WNl��ͱ#��``��hn
T�m�t�Gk(i��xD�cL��"��Û�U��fA�e`�T[	X�0�{�N�-�ٖ+B���[v��T���:�O�۽�:e۶�'.G�y�ݜ����9S��������W�L���Xh��M�f)�i����[,Q%X��ayy�ӶէQ���S�:^ڸ�)f�p�\�.��X6��yx��*)�4m��Va����+�є�]U
��n�<����eA��F�T��Z�.���mZ4x��J5L��`�ǆ�x�T5C�W�L*����0a�*3�,Pk,bߖn��v�CX[�X75D��^'�#E:u��Z���Q�B��	���au�U��ȑ9-4ƌ��Wu��^V3+IKZ���Ă���#6
���Yy{A�g��wZͳz�VU�XFbx3Hh�sm��%\̵O6��*�`(�0���͘5襌e0�hD�}U�)!�r��˘Ȏ�sj��f��d˻4���4d������+]S�N��bջX/4�*G�lۏ0]�H=��45��	�W�Q�+k/n��v�M�Xݻ �*f�x�h[�MBA�/+C'V�l)��r�Y��eT8s~Xj�E&�b#V$f�#��0�	'��ܗ
�����3HB��z�g2��J�P%	��X�b�V(��"�AwX-�yP��Y����j!kj�$�[������s,8k�w��ʫz�^ԍbV�[yzsfT����S�2ffkA�VA�ӻ���-�͕��uS�b$�̹�ݛe��&�K)�YH���h�Mw�/-ź/e�B91Sٗ��VP՚�a����D�fڪZv��9�e�ѳeɻr�PJ�/�y�b&��vF���B�X.��8�ˠ�;�����M��۫-�C\12"uW��B�A��)voFA1ɖ��a[�N�f�n�ω�Wx�?"^lb�x-���*��E��UQ�#XN��YZ���N���6��kj�Y��W�mLIm��ZNfl�Z�)�%�X�x񼱧N�Z�=�s��ܔ�e�x�t���{t�w�R��+t���-Өp��J+T����R�]��(�c���k�r��/��.Ң�K9uUHKve=�/t�*���c�2��jҤh��N<��n�����MR�Om8��+�)K�&��%-��+p��i͙Gsr��÷B�K�v����{-��	-�y@�R�Ò����<���_��� :�E	 I"� , �H ����@� E��H@��H,�F 
H�EAd ��ȲB � �B (I`I"�"���B) ��a  ��B, ,�HI �`$$�	I RB
 �$P$ R��!HY�a�@X@��H(I"�
�HE�) �H�@�I�!$����H�!�d�
BP� ,I���E�Ad��I$�R�AI��H�E$P		 
H�$$B�� �AHH�! R@�2�BA@	��,��/�a!!��$��l�q<�+?�����_��w��+5ݪ�;�r�� �K{��t��Ϻ��Qi�G!w��u�+����3�ɹ�Bb|��;o�:��桛�8��IV���4/0�w+�!B�)2�9}����b�m�-�F�M�L��v�f�ݹ�A���]ɶ%Y�܂�L�[T��&r�w�����xN��j�l:���D�7��������X^n��·S�Fq㦆=���ܥ��n���:�0���<�1�y�'U
T�PWSC'XT��eX;����ujW��m�p��r�r��a�`�	˙}�g}bR!;S��P��j�9e���Unگwn��zV��ܲqd�;�v>�6��L놅�B٫F���_"�2-έ�d��]Bq4ӽ7ׂT�ڝ�qï�g)����ݾ��n��&���6�A���b���Fl�U��e����Sx��u&+��j*j�ki�W, o1x`w�,n%C��Be"�݃(�skl_�ħ���T1't�Н��N���X؃�uS�-��+T�|��̷�f���;��Q]�����S6�,y���ewǛ��#�� ���X_*AJp�U�ۦ�j�4�\���Ѧ��:�*4YY��#��u@��3U>�Ԍt�:j����1��XOi�ѷY�s���n�[�#�ݵ1��ngv^T���(����
uX���+H�Ϲ������]m�к��!x�痼f[��mh|�/{��eX�&�Wf�	W�s-Zu�F��ij��ޥ�0HB=���;���5�{��9Qʦ�F�BYyN9��=d��{+n:�r�f����]q��g�ie��8�г#W�oCz�RU9�#��3{;���r��s��R�/�L����6�W*�RMG0lCfS'qI����wA\uv�[*�����'R��*�5a��4�5��}���9����T'�����]�Z����@��c���Y[��.tu����#V�N�uκ��ؗ�L1�:��_^;M��d/�r��J*9ҵ���;��gnΪK2n�x�"�sz�em޹Uw�/,�Uؠ԰��D�tl�H��W�{�W�1w,�֏\�a�
]O�TWWη�fi�;�{](�[�b��y��q�����n�,�UM���g	Ղ��훥��즕uóR�˚v5w���;�����4��S]8F�y�/MiRa�,\/6��WTqұY/z-̽Ҍr�J��m�f��ԧf��w���Q#��,��������C*�NξUU)_haTKyu��5v��6rhik/��5m�i�7:��J���ۯ3�\
e�Tٜ{��̾]��%ő"��r]���$��۵;�u�jB��������zuRm���P���)�S�<k	�۵�qE�J�z�J���/���i�����.��u�٘�feK���ϲ��#�C��uf�ݗ{˖iֺ�Ė��є��5�g�Z�ۊ�A`5Cu9JS���tS��S\�,�D����ч�_Z�겚����e�N�0�k��6��\W^:8�+n�J�r�7yvd��X��]�`hnd\���$t�εˮ�iw��w����ˮkx��)�v�底�]�K��޽�c�]5!�D��c�|"{;6,Ydax
8d�Krl�K�Q�`������dE�[y[[����-�uz�d喗<[�$�90Ku}���M����q��d��Y�N��{6�� \�������w}�����cu�Ba��H��u(�x����˫������*z,7���TW��5����̾9/;�z%,U�t��]sX���9F��_;���So���0R�n��^�=4��4/*�u�|c��IK��`G�H@qR��uFM�s�u{}�2���ݹۇ[=�V����ꢭ��:�a�5�,�Y=*�i���}�Xu+fڧ�U��8w(�4e�.�e=کSH�����Dj��{-�L�#�����6��qE����.-,�YCy��_qR��Q�6���Y׶짲=V�UFvb�e7���R:�+z��s]��=F�=�WN���72挍�AW=�EV�[KF�B�J�P諏����y�*���{VѾ�z�Ł�':�X����]WX̫���1��;���޵�h��]�2.�Wp9UH-����*#�wF_]Q3�����S�k��n#�W&�j���&�IT�J�#f�5�2�;һ����pr��+w9���[��eƲ�F�;x��Gx!Dڦ�[T����8�c'��x�V��*R{,ƴꀂ�,3gV�2[:��'��:�oR��uV��<��l��=��(3�-�;�{��4��u��&���ަu��Ux2]���N
�*��R����p\�v��M�JY0\����-ǽoXI���^�;7{e�5z�n�Dč��ysq@���N�gm�{M<�q��h���i;K���j��r������fռ�{f���w0���r
���çљJ�>�m��QU�az,��*響�ѕqLxNu�X�Җ[[�ő:t��ݺ�:em��7��B^���ͤ�v��wPuwa��zWa�Vv�ck����U��rF*u��d�Z4�W�t������:p})s�*��ou&nζ(�nV�fU��o�7����Ut�@�����8������qr������lfn^�l�7�P�l��N�}A�r���!S����.��m|�7y���+���ݗ\��;Eo�vmq��t����JV������d���ٰ��N�S92PUn���^F!SfYk�$�(3��Ω�q�����\9
��5���A_nmwAϲtB����UY:Q�ц�`y���556�%��:"�m�t�������U0�3��j�V�
��32̈́��%�I���¥��,N�2�TvR�o_b�Y�����)h�{ѫq���-��*�/�@��0�ol7�<�����Z�� �;����dه�+�m�����*���"�^�Wtq�[GY԰����eJӫ3:��;��cR�`�z��W$�����`�}J��Ǣ�	]z�Ի�$Br�vt�2�����7�r�Z]S1ު�@\���u�{F���9��Y�y1M��֫�B��e5�P��_}�r̋�vK3s���XtQ[���/0�\�j�`�oʠj'�py�Z)V���0[�9�g3�>��t�ߦ�ήf�eeuH������։�rneuV�UU\f[�3��݁�zh槺��j����w������S���tM�b�@�άvq�5��-�"�4-Bb�SB�L�2PA����moNl'��K�A��eP�u/��n���uǨvk��&���،�W��c�-�����e�q�csG��jũpܼ�p�S����Vm�I�Tx�m��
���|v�ûR���]�M���>8�P����/v����W{sg�j1�j��O�ͱ;�F	�79�����4�̥8��k�,iCk3%�EUV�����v��ҕ����f��,�ߏw=�jV�LG�+��m]��U,�ok���(O[�{�GHSM�u���j�����ǝө�>�T��wa��=���a���e��y��T����G�+n��Y׍�e�2��>�ow(tk�^�B{C]�Mml�g~HdG�VN�]J��c/7�ݷ+sO}�h#�6�&���'a��Tq���]�Vua6)��]�T7!qp�s1=�斜٘�Q���@�Im�\/�o%���5�@n`�`��n�
	\Ƴ������ƖN.H雗@�6U�:\N2w�gP�Gh�t/��+kf�c\�����!�k���N����ak�nۋ��������+2Z���ug����i�S�����=E9�h��;t&�:�3��چd4j�N�e���^��0�"BV^l�U+Ag6<�#\c�2{a�C��I��df�y%wuUe���*IR�]�@�*����7�:�V]�u%���ֽ
�VjB�ňfR��:i�g�9����3T6�]e^�%�Bd9/f���5oc�n�+��LSB��N�ΦpiUv�)!�*��*U���z2^��XR�om���C�����Kᖳ*�Q|�J��|�Ȧͱ�WI|��H�6q��7&-�c�`�+X�W�2�T�\�����F�ܬ��	ޡ��d�W�[��l�<�J_V`�ܭ��^�
�\�hԊpu3���{+����
ץw_q�x�1����[�יY������7k �vL�vR�4:�u$/]旜jul�&��Y�3U�
��I*�yf�]��N�}[��M�M���0h��kvn�4n].XWi�g����Y:����t�r�X��:QS;W]�۬������}转W�ա�dj�ܬR+9{�
��6��s�r�T9�]�Z�N"#�j+��B+����/Fz���\zw+ͥ��14��%�*�i4-4��L/�u��KÎi�Vs<W�����v�ҏ"�a]{�Ֆ/
�3�L9�o��]���7��W���i
{���9��q䪾���PYx���J1���Xh�Ѹ:=f�ou{CQ��:�*�U7p��S�{̗���ٻ�t,A��c5�#�J�V� �� ���:wW"㲊;$=��i�f]7�FG{or����.��>��+^ʵ��h/���7t�"�/v�޻�C�7�@�{3&M:�^.aW_L5]zo(�")�3�Q	�y���j�����6�0���.ݩ����y����FDB�9uP�����N���c`��0�oi�n�vvW^����[Uڧ��u]�j�Ƿ�Z���IK���v:r���kI��.�cz\|�y޶��*7!���V�9���=����rt�fX���h̏�����jQ�d\��[\���v9)�s7�Cm�\z�o:κ��,�om�"{�Au�����e.�Q�tUyw��\Z�2��ŨJ��XrgL�*�(�`�b}r'��2�v��s;�ǹ�k����v��>kv�wg��4�;y
��n�����o�ժ#�I:�ϸ��Z�����m�U�D�w����/ L�c]�Q�+��9W�'w�l�D7�s���L�^N�o*;��97�8�'n%]tH��۫����N����ݳK��bz.�M��M2a�"�϶�m`*�{Rҵ��f��Vvq�Ӯ���U�e�tm�g�.�R���Ź�ֈ��x�vt˥����F�ݬ䷶�C��[�^�g��­�Պf���I٬��v�yu���O�Rb�z��7Z��;;u�����W鼲�Z��[I��E$��H(���(��T9���׏*���xX�'B��p�w�-�_T�����*�uҫ��%:�k�k\w��� ��-�vEs��Y�@����np{F���w�����38rw��4b��]���3�lwQW$�Uѵ���A��Ev����mU�<�v:ό�2r�w3n�q-���,���nd6�F�h�c�:�$���'��;X�Q;��VӨ�����mwY��¸X�ܡ��ѻ��������M*�w*��8�U��U����͇|����D.��gHx�3(�`j�P�j�<n\�=V�:��W��@�1+W���vc��B�*d�nZ�0G*$�쑌�����nG�x�����n-���b�;���Y��:�1'j��{C�,�c��6sGnTu�zi��$��u���պW_h�"����w��bh3�Kځ�ԫ��mEZ�k\�;�kn�;��Wv�Y�����1ڷj�\mf����n�Y�ԕkf���;t�X���z��\����9KY��.=��>��&3�ۥ2F�CB.��*�դ�����N�|I
|ˬ����X����S]m^n��P�J��Q	�{�vY�縑�{f�H��ת�9Z�nj�W�Wn��o(5�O3�=��>ɢ�<�v7����󴵉�L?m�ɵ���3��p��V.��
9as��H��P&�����l<�k����˔[����IJ�-�Jt�&�1���q
�[�xi��U�L�:�3�+-خ���\7Dn�̮���b��-��:ŽS3��i�Y�@x<�J��h��8��eSyy$7�>��w�V�ٝT�en�Wwd�uj'�̶��{�e�0�]>]D_3{)��c���8c��oN�Y�A�ׇ�Έ�+��h���u�T��
O+��,�}��8�[۹f�l����*�}��ͼ��U�Ӹ5��[��a��!r��o.�p�ѝW\e�y<���
�8o*�E1v�L���C����!��N�=}��ef)ָ�k]�z�kE �l�q6v6��
�`�t��Rr�u�/�3M����v�����m���Kp���ޟ�L�]�A�=Q�����R�-��wF��^��;Q]Ս��9�|Z�Y����]KԝkD�[,�">﶑��7���q���Y�<�̮#Y�U�u-!��[�L���J����
�����������u�k5CW��w>�ȦUv��Co�ݢ�ޒ�!���������:��p�D��L��*���3M���o�=I�1ݞ�b�N*U���an-yUS����,=��T���,_m:���NĝX1��t�32XUM51=�/���V��\dE�vfޝy�u��%��c+�T�b�__��ۋ�jT���k�k�>��4��+y��n��jsӟT^I)��I#ŘS�=���т��ͮ����A�ԙg���X�LX50�ZJ�|����*�S�,�n�AR�����Vm�q��]��SU�ha5M�N������EY��c�e=�F���<��\��;�����sw��NެN���-�2���n��U�a�L�o�{�P�DdΒ�|�vT�{��v�Q[l�ښF5]Y��n��ww�ϓn�e�kjc��t����2���s���(�u]ah�̽�n�*PKs�S@��T�����M�������[��qRn:���]1����{��F�����wJwXt�*�z�]V4�)]k����Y�(���)���b�_n�������v��n)
I����,���[��ٰ��=7�B�:*s7Z2�~�{����I'���<��&`\�hlKI�.lrA�m*n�f��a[��]�0qF��u�X�K�[���-&�J�cՈ�ʽe���	s���F���eHeu�6ᬔJj������;Z[5�&�`[-�W�����.��ǜY��GU�Ԛ�L��:[y�Ү�f.1�M�-2��d�t;:�ڬ����w�ꌥ[ZYT����Ye���,�����:3��饠R�Sm�vR.6M b£�,F�$�B�+yH�k2��5-�6pT�t#m��5��N	`[N�����\�Rh�C@�z�1���Mvi����9{;ma+����˴��Ys0J=�2�,MJ�%�/XL+���Kca�T�t�v��0�(�T�8���t��2�3���D��\Yi٤�Gf���J
ŁGX#�,���jh�d��@ᔺYo1{#���,ζ�k�3B9eq.y���ʗ6��al�f1443�v^K.�{Q��X�E�;XSB5�R;�̚�
�qenWYl%�����������h4܌`DۋpR�S�Gg
�[��94r�M�AFl��a���N5Yt*V�č惦�
kB�T�en��q�X�]�<��8	k.��[5�[ ���4&�W�CGj���k�lG#Bhj8�^g�K���ʓI��%W;;i��E��Y���mF�AchJ(��έ����K�V�6�u�7h����d��F�X����]vq�Q�^1�6����ΕW�v��#���TZ��&�H�b�
7G1�hRP��3%�k.a�m��٠������[I����llɘ�l`lq�%+�M�5�l�)���c��Uܗ^f�qL�XM������
�],WT
iI�u�=�m�E�ci۝2ۃnEn`ݫ/f)rm��.�T�b	���ƖU��n��jG.�WRPv�����}6�V6[ rՑ�*CV8��714÷R��Ԕe��&�����m���f&ٹJRv�i�kk] җ��DQ
B�U	�$�TM��c�+ΔQР:��:��-�jĭp�q�s�i-Y���\��Z6���l�K��+4*`���A���ʸ����SX�k4�م�n��MVb�%�HfmYsUR�4���c��X0�Z���X�!�S;\����G�--�Ė�5�C�+\�\��kX]&,t.��Z8ٗ6�j�kH
�]
��i�X�M�a˥�@\Ye4uZf�cY�X ��Fk�i�b����bk40�X����B�1d��f�G:+-���,e�E�j���e&M-3m��%�����K:�)F�8���:lA6�Gu;=��ԡ͍I[ttt��\^fk�����8X٠DRV�R���ջEp�i���bX�v�Ų�3����T�X�QC+n�0�J��&6Ķ�:ͩʗ=�����dd�1U�۶��b����U.f:�
�ZI�6f*�\��J�u������%�5D���.n&"	/5�V
L"�md�v&YS[c����Y��ZZSRm��Am4��t�B��W[B�B�)�K�ʢR�4%��]�X�*\��Y�b�R$���yM%�u���du��R[hKZ�3��/h iNƺ[���0��٪�2%�����J��4��V�ΰz��R��zn`0����4Rٵ�aCGS �h-�7
�Rb�0��:���mZ�
�I���v��fH3B�����j��R̊8�`[{KE౛4VݥHB�h�M:�QҶ�QsBV�i�.Z�m3vl)*&�5�od�&���C��[54mPÒ�,#r=��h��вV��@�YC��;c7nJ�SA�V�Q^�	+6������[��+����ir5���[l�])�B����GL������)-�,j:5�@Np[�k�-pd=e�}Uc�)2cA�ٖT+�9��[��F�!rR�yöx��[�i��-Դ�rk��+u�t��i���u�y�m���P����	`	.�,Wb�Z�E��꽋�at]R�5�sx)�dQ���]ـ�{ss����R��%��K�a�v�)�b!v6WD�]��t[u��K�j���QD�9�ZݢRť#vD�zb�s�R!��E�\�҂W\f��yv֪82b.��	�N�@ˬM5M5��XOy9a=�Ʀf�A�#qt�C4#��\L�Ùn ��L�=���<sVPIF<Z� WC0�-Iu��lT1D����9����d�b޳9���+�٩LK�u3mP+2���ˏo5�$��g���1�
͠�N2���^v3	Dd�#+5	D�soh"�YmLi3L��x%K!�au���=sT����kBkeΖ�����&F�n�h���% !x��lr,�����mա`#��&%k5�iU�J�Cg!3^JR��U�gJ��PԆ���;=�ƺ��w%�Yjp�B�C��gLW��^��͖�r�7\F�$��rj��!u�LB�W�β�ԵD����BU]I� �a#[jGLlҡ��3M3S�]vez���V�ΩrEe�x�i��4RZ�J�bkXz͂���Hڱ��Va�W�S:c,f�6噪#��(�Y[ �a֊=��2���8���Y��p�ke�WVU�A�[���(9�9�R�5�-�P��5��6�� j�\D!Qs)��6e�wv�Y��,�}�o.�]�F2����BY��1�e��(5��K��T��6}t_j���RnF�(��!�ie
P�И0�ne4��n��n�A��	f��8�앶%����d�,b����`J��&��U�ؤYv�s��2B�ۮ�C�ЬZ�,DiVҨ�jkwKG��{�V2�6�T9�Η�Q��-���Z�e� ��"�,^F�6@�v�������Bf�)�ɫ�u��M/!V\n�$lM�X�vL�uCM�kq��D��)2�Ǯ�L���ne�qt�0#-�ᎃa��ѹ4��� �d�15�Rd��b��TskQI���SV鸘e)�ՖM͌�83��[ۈ� f\.I����+lCJ	!����U3z�![0`�J)�K�l�C�\���\K�X�m�[f�8tp�	e��&mR�1e���0��%�6���u�)%`��)
Х������Q�(&�YWf9%b8�f:`3K�mWB7e�J��)#s`k��6�c��v�t%��X&.F��i��3��ڒ�kY2[,����i�U�q� �am���&�T��qqYw���c�^&���B�{Ȕ����Mu3���s�4�K��r�AlfָƦ`�k�2��h�i3��C v+���5i7.^\�L�i��tT��L�3�z�c2r�JhQ�	2�k-����2h�(���Vb�G��;J9l5�Ґ�Z�56�#��"��zd�e�rL1�l�MH\3;ެ!A�MuIcB8k ���EM57S z�4&�b:����0�Ĥ�T�!K����1�C4�A�qZb���	�����+ �i.�M[��˶�%�\�Ts/1v��.�[�3[
'g , ͫwo[����J�б�
���E%��tI�P��%�9$ZĲ ,+�yu����Km��[��v-y

��0�5f���ѵΔ�dҸ�,WnKc�����;�f�m�څ�B�Vb[P.���H�MA�6Af��ۙI�E],0�J�v@[sU�q�
!aVl�HZ�3ڇ�}ea@J���Dڐ���5��(�٘`�8V�k����n���̭��Em-��Ye%5��2�4�������l&)�G��1�k�;��:쥽p�l=a-vm���#Fm�X%�CpQ�D���%���-�D�ۮ�BR��X�ġo%-Ж�M2͘�:���[L�<Gt��ݫR�i�e�;JD�Y��Pu��qq-u�5��3��5�TvX�J�F��M����a��R7MZB���l�n�h�T�s-:�=V�6�n1r��ܤVW�2����T�R�3��Y��\�G)�T`n�����ҡt(<ˣ�e��P����T%��q�Yl�{Vl(G���pih�n�e�Rfe�[o[*��u ���z�R���YBʻU��m.�UD��̶�;Ds&M  gHj�3n�\�c��ś ��Ûv�]�s�Rh�f��e�ı���ju�ȭ�6m�it��J��b��Ź-��hl�cG�6fX\1�R�ZM�6��u�޳Xѣ%eT�3�\0���R���y��h�ͨA���K��hkM4b�%����[f�LbfB`Nh��X�FD�ut/%�z�ku+n���9f1c�m�0�$��b$%�85��H�i�v�l�G/cF
���æ@3+̰*m���V�iit�� 4�"�1uNW�GZ[2 ��i��1m�`�Mj��)mN�������Q����/3l+5[G'n4����)�1a�:�p�]5h�-�x��%iSMf��)HiB�nXKjD`es�hX����6������nj�ٲ�*̖�ˍ��Iib�p�Pn����*m��l�� �ɳ4KU��)^f��� ��a���n��VbGJ5�n���,����d������0Z���Tm�]f�o&v:�mvT`m2�Ze*�9�m�ꏒ�Q6�9��)��nJƥ��ܷ1SJeK.4�&���@
�v3Vk-���T�0�Mbl��5� c5VU4IvPJ�7�4�]Fh����լǷ��z�V��[���.���n�L�+`��Y��W25�1o%*�D�ڵ2�g5�Ci�v3=b���.vS)���%&2�k	b�۝�����͛�e-�m4խ�h-�6��Ŋ���nL$*7�ՙ�B5��],A�\���\^!��(��5��2��
��gK��5S�a� �e�2�-�3�4u16�-,�We����Sh�P�]E*�[tP-�nf��2�=�Ꭲ�쫵�f.ՂX��Q3���齵r�ʎ�3;(��Uj�V9C?�!B|v�BBwqɶ���ɚ쐲"12�6��#KV�Λum���wgn��+ӳsM;3��wee����oV'B(r�X��[�(���촳R8.:����
"����H�wvt�f����gY��Z���^wZ�m���2���D���ˠ[v���E6�Ȭ�vnٳ�ٖ���[����<���:�:,�XtI�%vv����zͭ�Yq�fvYg8N%'e�m��N�ҷ'�Ev\�vBT@t�w�q�2��6���v\\�-�m�JQ�l����X��󴠐"N�*r�.��bw %A'kM�i�Fd�R�R{h��Σ�"�mgtI��t�	���rp�[��)=�'��_�T��F�.�L��ː��cX=Gl)3�eyx�Ÿ	�0����3fsu(Y��M�E���#bm��!&M1]v�f�
�0۩3�l̨�2c�S��Syu]�R�f��k.�0P�B���S%����r�t6�M[	j�ձ�9�1��-�GJZ�X*�b���2����^�itб����6Ҧ]2:YHV-q.�e��l1EG�Fۂ	u��
��f2;gn:�QѰ����4�V��ˊ�F\j$%6����Į�i�l�(M
��3c1��Y�	�#�)K����D�#[�F��1c#5Ҏ��&��m�X�	tl�hhl![pM�Ͷ�����3,�.�ta)�!)�En��i)�9�����ك4�0�V��Z�-\R�-XA��x�Л�X*@���IF�����X�\`Ca�R��n��.�h-�R�lЄF\���%eީ�oLP�
R�Z���-����a0�����r�$��a�Ø-l�&��볘M��]^�ɋ� R�����4�ə��r.�l���E�ѵ��h#!6�i��4�l����Gbi@�Pb�6��Pu��ƴ���[ꪹ�%���û���㇕1���kkrj�P�s�MF�K�$��J78��{C\^�T&u�d1��5⣨�]��&�;B��jG�⸁rd��WF��K��\hֆ��X���0"K�]^�j&6��Q���\�obe���ԁf�,ҹ�٠]�6�c5jPZ��G2�\�x]l�jW�DȌ�`lhd�i�k]��K�0u�4��4\Z�l��*ge�e�d��sj�i8��Ҙ�l���-������м�Fj ]m���)m	�∭�j.&�aՙu��5e֦��.��6��2�]*!�J��� �4i�e��-���4Zڧ�95̴ҳa�(�@��8o �a�"�Ub�if�glY�P��5ˬʭY$�mS6���Z�[
um^G�B�p
ʍ��8P
=m$��un!K@�o ՄK2�ŕH�z���[e
��z��@�����)�<+VR 60i�=yb�Im�:��,���� %�-K 8�Aj4�ڼ1�-������Դl�XZ��Ѭk�U�J��������'�9�	���h��4����+JV[��mA11����t�vb=v��|� �n������,�}"��ћ�0�y�6��8��΁H�#c��d�(Ⱦ`Ș?Wy|7u��vI䥃}�U��.�"�$�G�"�� ��9�ɒ��o�l0D� �y�R0�0�"ICw�J��Xm��X��};n�{���|��P����dO�D���j���I����(�x�3z�L���}��M�`Wd����:� �,ϊ��-��a���w}B�2&&DȂM��;��ZʃCL��3(+d��]�������=�Gr�d���~3���2�ibSG�m�tH��ef��
��K�a��U�����Z�i�m�������YY�	�^�M��W�CU/b(�����"�T=M����x��Xȟ�I*�2 �q���<l�������Ur���II�h���\��O:����W`4��Q�]_\	�9����Dxe��Dŵ,=�*rV��)ԋɡU�64B;V�t*�(��F�l���T�qt#н΁ $~OPԾS~_wB��LA�2�W�, ��|rm?
Ω��.�g�s�how��L�0辒<#�$a��ϫ�|�O��z��F(>�i^�jj�0���r��b�48�y�����'���&P ȃ ��H���#�`�:�ɴ:������M�֪�O� MU�	�P	a�$aZ��(r��ϻE�X^��E�����dI5.�G2�d�e�Zee�y�36٩��ި&��ޡFD�&DǄ�����w6�c�b��7қ���;$l0f��	`"�$t׳�ˬ����$ذ��z�(��j0��K�|�"H�|dS��E�;��.]n
�`���2��d�ꑌ�Qj�ͦIG3�K�oC�$"��soX�RNP]�1蚂Vn��̎��nR�Њ�M5��g��$8IR��s�{�.;���6�ڹ�[\�h���{��؆|D��$b�2&F�J)�պ� sv.9ϨA3L�*�m�sa%b,��G���*�p�okv��ͫ �9���� ��D��<,��L���ر�8ҷؔM\5Qݹb o�"H���dWh�m�W�nM�<���a�[.�hW�KIG@�3�3[�a��\*E�$P�_�1ц��@H�P[7�~���+���amY|qo�3��\��w/���|dL�dL|G��M��R�n�p�1|�;;s{����l$�E��� A2(�B8���>��g���F�`��:�da��z	69��mNE:�Ü�k �u�^ �o� �( ��F;o�Z�{�`i �y�g��$A�[&5����T�j��^�!��1/:3&ᬉ}�BVH���GC�u���Z�ή���k��cN3��7	���ifj�zuP-n<�9;٢�ͩn4�����a�^���(Ș ���$�(ȕ7�.�;Y���Z3t�j�3���X�	&,Dq����v1�n��\=~lWO����&�ې(��x�鮋��Rش��o�L;1�Tɠ�������~��H�z	6A*�n#UXm(�s6_�]c��v��{����ňn}^�gĝ"	�P*�N�U]�<���(ף��z0��k��m�j�\5:!�W9P��(L�U�U�yʱ�*ћ���Z.��޹�ES��GZ�u��X�E���� z?��#c��*VFk��X��	ez&��E[Ü�(b9�.z1Mz=�[X�U���F���ͫ��0c�E���n��5��WE�C�PS�5���8�h��`�{��z0�7��IC�*jv�|l=��زg������K�貎�CdYf��c����ݍ�H޳ٵx#��{Y(ՐL4:Ӣ-=uܐ���#rS}!��S&G��@��TQ�TC9�l�d���(g`J� iu�[�/�ke�	ʷkF�if�VWXL�D�tȰ��*T��d!P�J P�X�@�̦r�a�:f3V܃���I�.K6&����32�n��W iZe��I�Lʉm��hڊ�1G%�Eq �:c���SX��{[1-�X"b䈢]�bƮ��[���F��m��9J�1�>��/�2̶]X �c��e����p�R�g�lV�!�8��d�v՛����}��G�P�dL	�>sgu���o��A$�dЋ�V֞�*H�
��΁ �7���"�fW�I�鬧�%½��a�$��,�5�K�Gwe�>�L�1_��:F��z��">2G�Nw��V�n`m�X�7=��v��<{���F7�$ظ&h@�
BY|�(W\rt@x�_���� ���]nw7�U���v � 88�C��a��(�u�*�@&�^$���hTi�7GiW��.8�y�mEe�����}\M��>�A3�g������7��f��0 �u�4M�a�3bp�ir�K��GQG��9[
��ￌ8����4�	5�Р,Oڞ�M�$�\11C<�Ϲ��m�nda��/��`2'��"deU��郙�t�W0-k��a�N��o!2�Ef���bĜz��^^{T:� �m�� �`WV�<Z�B�f�ɘj��"﶑ŕ��ٺ�>��4���V\�w7Е���b�G ��?����f�Pf1B{�0GG��^�hP�MW�ěOI)uFfj�y��[QS�^B=�,G�M=�ظ&h��푅]W*��7��0�+X`���2(Gi����I��bb�Cj�R��{��[��7�=��3�$b�&rw�W@���c�[4���^d�s/���bw1�� ��3$tD�U�N��߿__�ׂ�~�Km�mb���,��,[.��.]�*ŕcc��CM2M��o�~���e��	��x�b��V�Kۉ�����b �C���.�/���`���&}@�`�)d����`7��[P[��^o�'TZ# Cj�h_T��Cs��{�ν�X��\D��0wh7h�Ӷ*�^���u�}V��őΙ�$]�u��W+
�^K�G��2Z�Fq���U�{��}/Y��FV��DKZ7k�����WBX&�I���"�<�zH���	-�l^wM�F�T`�������ow��������?F)��8�^��{���CǼ� ��dI+�Ȁr0̑�?���}�*ЮwV�d�2uE�1?P�mU��T+�	�P$��;��z����YJ�A:H��J�3+
�r��p��5]��B�+�����!�Xtz������-ϫ��ň&k�"	����Vd��/�u�������^*��Ob���w: �����Hv�!�N� �B��lZ�)[�/luV�-vX �� ��W�)}�ŕ��"�"fР@>�D�0d��17h�xd����#�����Z�@��\�* ��$��_����)��X�T��|w��x�aof��;|��K�)PpL��ǜ�u^ڠ��u��Sʗ��'����se[�W�� ����S	�����4X7pkkK�}�V5���!WIh�{��=��:�}/;0{�yΈ3�17l����Gv�u�ͧr���vp,ر��}������'e�z�zJ�E�dO�/Tmz��l��]$�YR��l.�%s����V�i���ݳV��`I/.P ��2GDt�Hu�.��Jg�vy����*�T�
��D�\v��wp��ՌݫΗ��gj���e��mdm�+�+	��ǁ�A�a�d�����ے
;�B����y�F�H�rJ��Z*��N`�d�F�V�w������� �$��X&DȒ1X;#�JN�8��3$t�H�^�?{�q��(D6��)������%ܮ"����W�gDx��M����;��7��!v�J�r��i��D�����|D�[����]<�{t��WF�1r*.��پ��Owٗ��m�qa�yU��㴕�z���u]V:��8��g��P�\E��V&��т}�����,�\��F32�a��Ҫ�6��n�v�u��j�k�]ma��faZ�	f��Q��#*XA�34)���M.�L�b1̣�q��sl�aJ���%Ю������Mc �`z��[��8��^�x4le�l:�P�
H�k	\&5ٷ �e�҉m��.ɡ���c����m���TKe��v�ĻK�v3R�A�\˼��|O����e��mUc,Ұk�m�S�WQ�t�Bi�U�Ih�C�sΈ>�2$o����vS��Y�����z}u�<�ӛ�P =v(� �"dI+�_H�"�j�S�ZH@�΁�:G$;����ʙ���`�{�����]��ߓ�7�ܙ��2JdLL�*��UU��V�7��^��d�=���d@>�0d��H�"F�[ක[�z�A�;��att��y]خ$ϟ��
y���s��_0g&F(Ȁr0�2GQ�D�{�>?n���sx��{��g$bb�ګ��B� ��M5OXU��;��<���m�Sd,&QdA>dАpb.kUٲ��M-ɓn��˖�u�h�K,�}���͋�4 D4[���Eo2��49'b�T��c���!zy�
�N�@"FH��<`��������wk<j�n1w��uk����[J�T��Ώ��U^U��e�tZ�xmg]�2�i
M�uj����k=.�QE^����>�͋]%><͍��b�$ϟ�Ёd�@Ƞb�p\N�ƃZ�mP"8�Mx�[�M���3�]^V�y��̇;E�/� {�F�"��(Q�3��l�ZA���P2'��$׃{��[̽��MI��z	�.�ך�����Z,��F� �#�Ш�p͙'�^u�DrO�>��ݿQ���7"H��` ����/'�>�8�]*�P�m���j�CM�!ֳYu�	�	3�5+�N��UH\.�
5 ���d���B�s�F��[�P(�H��L�y=�������v�ݸ�����IB���~�?�;;���ʋ5��>��'|��ٻ����e�%�hjO�"	���	5�A���.L2;�`��Έ20ȑ|Ē����xIm1��/7Z����6��:e�J�3�U��E\՝7[z�+�T=]�+���<68:�ua���.���^�׎��*�'n_V٢�n�Ǵ;+UܫQ:z���F4��X�fP��g�nҕ�S{�,�d��U��J��
�j�۳��-o\��1�5������u¨��▾{xF�=��88�5λt���VU���6�\%>�B�~M�3�R���9f{�X�»�N���6���ꈽ�w�n�zU�ӹvv����(�O�;v�Yм=z�z�r<�hp],���]��5��5F}�u�m�����Ǡႋ�mꡙ�Ɗ�쪨;s���̏��rT&w˳��v�u��w+ow�8](UjDj�qu'�{�x�WU]+��;������eJ���-͕{��ΘƵ�e�6r=��wb�k��/�'�䣯ǵ��g0��>x�k�aly�V#×J�4�ZMK|:�����p��m�e7��LŶ�j�橜0f���HI�F_����IJ�
�x�s{t�e5���7�B���$iv�j�t��!b�K=�ԙ���X�L��]�o566o��g�b�������q*�9��%:�ԕ�t�Ʃ�]�q� �����U�.2s#�h�2��9ʍot�(l*�r�(mue#�i*a����0��:w52h��o��9{33n�*ô�}U��ʡ��Ir��}�%WN&�.��bk�zv(f��uhʮ�%Eu��ˉ�S���t,�+�ʻnVďZ�v�Ӝe�Vk�̎|^Zg1�������*���@�8*ow9�2��`u������+��g/o�^��<B�)U*���)9ABn���"(fBI��Ͳ�:J$��ˎ:��4��7'$Ng7d�$#�*���Ar��䧷g�I�v���ĞVe�t��P�d�	O[�� f�{n����ҳ��Y�f�rM�1Bp[b�66�ۭ;�7`Y-n(��A�gH)4�N-�˜�Z�l��b��92Є�M{u�O-�Y�[k	�vQynݰ�,���.'��{�9;�u8��ZnfRq����m�Rk[�˶ȝ�������:���o/A�Mkm�TA QpfNQ)E�]�A	YFt
Qf�r8�!���S�:9F�H����q�
���Vr�e��pボ�ۀr%#�q�ckH��:D���:���*,JDEo���{�?s������x	��IB��|��0D��N�Ѵ����r3�q��o:��	�q�Ʒo[�*��H����X\ޣ�
�oٕ˳��"��vP����2/����N����û�=���������e�%�hjLX�&@�hW����}�"���*�9A���A�7m�aY���I��%�*eG]0�sm��#�y_l��A�2$`?��{A�������o��l��,�z�Y;I���(dL�#�C����ӝ��"�B种vv7,UIZ0��Cҫ��a�$K�/�fK��t(�ɂ;ɐD�� ����;$ЕxWL�=]�-��MI��&E�kĚ� � e���k��w|��A0��?hZ���q��Wc�K�� G��}��D8��fB)۪9Բ2}�뮈��{T��!�x��S��SU��۵Ow�Lݯ������O��n��g�C)��K�/
�گE�8��?w�"H�D�3$x>�4Vg�z߻_l:F�x�y�e��' A?d`m/�u��kڿ�:=�T��F��"�(U^���/b͐kE��K���#�l���ׯ��_03z�"d"c÷p΢�=���a1��z��r9�3��@�.0�w?�F?�?#�G�����*A�棆�y����+%>;��:�B\L����n��&wv��7�����##���	�°�7u޸YwY}Θ���3��!���9PX��(Ș#3r�?W�`"O1@�	���`���k\��hjT�#�67_Oz��؇�t?w�dH�A&�� ����h��X�#�ѕ�,&!���=Ί�u	i2��j&�L�Ȼ��*=*v9�k�?P'5z��^�Sx�ޯ`�(f]3�L߮�ûn�xe�J!3�q�z�V�����M5U6Q8w��3TE�h*L�狦�:貗qZm�2�r��v�
�34���J�[4�v��رr�%���\���:�u�����Zd��ʓX.]����l��[\	�t����{$K)�L�sh����d{R��Σ���j5��!���+���!���eD�h��5�/i,�SC���KI��Xu�׆l6�l�[���f����K����tXK6Kl-X����T���.���TF��4��v��O_=3�K��цd��"F�we=�^���5�bt7�`�f낷������(@�_9%}"�2&F��P���2���v�@�AR��ݒ�'�Z�-CRv B�0GD�??anꕝ(W���o�tt $��J�S�}�<<�P���{/����>]�/Nrd%}"���&}CN��^Yyz��l3=�@�b�7��8\�N�Q\�&(@��\�@��=�jz��=l?��z�"d%
�ș{��I`���On���ͭT����1b!��@A&�@�c�^/\�mucGΚ��-�%4[��p�#FQ]G�2i�.����9��j]p�0y7ߜ��tG��l�v�'{7.����\�$^��TmK�r�+cg'�"�I�#�L�����^��o\3�1�!��[�w�2��Tm��_,���ݮ+����x�tН&�>T6;�"�d�s Ҥ*�a
�u˳L墶�9b�`��<d�P#�Ы��6��r�:qEr�?mW�o0�"K���&��]�,�(�LO��I_H����>�N��P��s��T�g9���@�� tI�0ȑ��I��K�R�砃��#�W�M���S㷯:*����ˁ�Y/
u,rg�P	�H���?kt�s��(z��Ff�J@�8����D&�ܤh�M
�M������R]�1�Sd�E�Y�L���{V#�6P�	L�X�D�V�� YTIk��f�W�!ϫ^� 4o����A3A��M��Mj��M��4޽�!�X+�)� b�B9��������/�4�u�{���%�(�+��ذ�G��.��\�J�e����#d_B���v���23r����da�#�"F;�NNyV�V��PC����6쎕[Rw��n��u��,��v���X�5^�i��E%�p�3jfF����f��ç�cw�������x[��ICW� Bj�$�H���(P2&Ewcl۾TGtb�4 D5�wA�������T;�	�"�<�V���bzGD��H� �D�2$�Z����_.ڡC���L]�5=�g�E�A;ɐvJd_3"
c�]^���J�T�AE�(2��,p��.����u�ƃ�54��ŬM�j����>D�A�w�`��F{�\��A��S���uw�M��:�35� �0���"IB����L��=[9s��cc�Ё�`�tR��\�
�ܝ���d
�̖��p���@�b��k�M N
�x�b�b��vJT��&��=������ϟ������3��gĝ�2�w�%�d��"�@�B���&���4��1q׊(�S�y5W"��m[Y���s��V��u$��M�^�]UN�}J�pJ.��,1�5	�2eo׊�]��N,���ۗ=3=���]�;O� w4�'9w��`�բ;�B&�L��vc��sD6�9h��՝c7�+�0A��H���.�/;ݺ�P�@S�2X4i�I1T�tat&hnvZŖlF�Y��nIW&���k��$�����y��"G���$�C�5K���:�g���fĕ�^z{��x�|}"dI*�2 Ț���1������#���4��1q]�$�S�Bj�xr�@�=�b�Ek=�~��У�� ��0A�I_H��dKk�euR�"��1���Y���|z � ��3$tD�0D��1fI�R����|�@N��P�ä�f�GM�u��=��M;�1�5){q�W<�z�F��@��5 �~�� �#$m��|&m[��L��\Wb�(�B&��@�B�i�D���e��,Z:�4�W���\�K̵,p��j�rb�Nb)56	�)oHpa�s��Z�쮭�Y���[��FL�9�mH3�/�,Ż���������݅`����\�(��B�D�vI�����j&v"�le��Vk�ir�U�e,o&�95�kcks�%��jLB�8nF93��ZT����]��d�b�p�Ҙ&�X��\����0��#c��E#�X�Иr"#Xl�UR���v�-�.�Vh�)�L�`�M���z�{L�ݢL�$��M5����5�y���?��v��8X촪6]��KaڗhY��D^u���IX�=}��K,���,�>;��wAvi�/T�B�o*h$�p�Q@�a����	dH�$t��Ϙ��oƢ�wR�a�G�X����W��7��-FX��j&Ł�O����s��� �G����1���+����O��{������w�?�: �0�"E��IB�3P/��*����V�H� �~j}�Lט=���`�]I	�ܫǤ8���Ҿb|j��w0ȑ�2G_������@��_�m�ä��(�u��Uz/A�L�6JdLL��+�pՌy���s�^,+�L*N�M�AT�(���H�09�n+�lSg�7�,!�!m���ߝCߖh��$x�A^�Үv�V�|jp����{z�uoJ�~NA�;��$�FD��&�/Gӷ��V:�����wί��.S�;;�{.�{Y ��Y��x,%Kۛ�`�Q>�}3���p��&���v�v�^kn>��w`��k�"�@|wG��s��HM�ňD ��0d�i��o�6���49`����:��dH��I_h���"�>��d�P�L�{�?A3C���$���,ݵJ�{948��/�X�L��9ƙ�+��Mb�(�B!5V ���֙�6گB*��	�W���Jd_Q�Uy"lh>�c�����^�����P?F�: �$c8Vw�9F'L-v�9T[7Hh��q��[d�3X���u(͙�6�1%1q�l{����t�A�D�?���}������U���t^ ��筊6�yQ��Q�/�D�J2 �"�N�}��FC���0Af�� B�c+��xW5Z���w� ����	=H�Żv�c��W��&> ��}$c>2&AEi��L��6�ߛ���Q5�I6��[�#u�(9���vV��Z�bh���;�	ث��ɼ�O�	�sa�DXJ�6>   `��d�kv�c�|,D"�ta�$tD�0D�3�Wu�#y V
�M��q�Ʈ�%�-FX�A��!ؾ&�u\���P@s��$�@�dA���d�75���}�`��_^s�7�X��:	��9P�@%��2J����z���*�
/!��X�^�vչ�!��vsn�)@����3F:/��g�
6.	�"	����s�/>�n���j3�ף�BFy�}���0D�?����=�-+�^�<S�M�|#�8gUo�]B�e��g&;%
�Ƚ[^�
��Y��.�g��}�A�A0̑�_	�5*���Zyv�-s{U��?P�,Ոʅz����"�E\J�	3s�����6���T,�p�g0V-����LX������n;�zo��k_V-���_*�ׄ맮j�kq�[�0W[�o%��m�	��ʚ�oEk��������Et��Lb�4�mP��������D|#���}�2$ld����"J�T9�4n(�R���8gUo��J�e��O��B������v��op�����\i��G��0��.n�Ĥ�`2���h:�ŕ�L�`���xP �Pd���Сc+��<8�^Ub��LP7��J{$~�#���$��X�&ݱx��L�Z�n�L�������
�KR�(N��b ���
�M[O�G\��}r�P�\��Z @&�'+��M��V^���b��[|6�U+8� AS@�1FD��E����ʷ�i��ц���:��~�}�V��N� �G�z�i��k�&�
D� ��IB��h&�W*g<�Oîw|'�����n�}@�"�F�:"DuO_WW�4f�!ڼ������꒵��U��E��%,U�W��U�����\�L*�wu	�1p��U�+����k�2�m���S�%��Wiȭ�c˹gaR��/���q�5�3(C(4{Mp�;�us���g����Vn�����]�[J�m$Z�}��V,�6�]�K�{��3w3wu�-�iݢ�h��%�ulW9���u8JK���\�&�b�*��F���˰��E���̗۟#���*���bwR��V��f�6�m�u��Y�3�J|�w�Z�Q*�u����&�{��,�z1�jЫ�(�U�92��[G�Tc0Z�Fn�q4gZ����c뼪��s��#��Ǚ`�[�{0n���;�bm6B�n�U��<�ےoG2t�-a�[��u�&^wJ˧(W<�\H��a��[3���e�v��]ji�u��r�Z�'hl�;�������V���y׏��5F�w]��9]�k�j}f㙻\ji�F�����b�����/��f��z�wp�Vx�r��"U��>�ʆ�j�lB���ܗQ�u��!��ǧ���emUV7����)u6�|�%W�4l]�����線,d�i%GL�d�j��੧���v�ɼ�����V�z��7��]��}OH6GU��om.�)wm��QYf�U�s�!̵8Q�W�:����ܫNu.����g
	*���8�����.�lC;#Z�O�=x;�˱�����ö7Kw`'Dwg걙�z��}�v�	�[����e�s��/:onb���6/�mUi���ԥ�����+D�8��Is���@q�$���v�絳�v䒇JN����nL�s�JNp��D�H� � ��Gm�����#�VP�\i��$S������K4�$y��\:ʹ�G'8)NB�6�E�S�H�"D�ghm��9%		�P�q�2����)���k9�ȹ'%"�B��y���'DZ6�G&`�2�w(�D[dFՒ��R�h8�q;����$��3m[�� "BF�:"�-�$'�G8�S�mh��Np{��tЖvDY��&�pq���{g'N$<�rET���S��4D�"N8�H@B���~�߻��A���Z֭�镫)�i����k�]�b]E�p�R۴�ы��E�-��K��iFh<Ո�i���L\�m�Zʖ`� 5��a�H���&��B�^��h\J�(�6ʰl�!T�0jYI@�����&]vu�6�b-[�X�;Bmi`�WBj��k]"�����ME36��t�����rZ��Մ*�����j�M�\a	`�!��.o�<��i���ƌ��"A�1@�,�\��i��١��lw:�6�m0��B�f%�m�Z٬��1��B�KFL�q�Q�f��lMDT��+e2�vm���g)�]f�rTl-�,�e��M(���ڒ�5v#����)��ٌK�Z����zܬB֗Ui����c��"˕v�3B��\U	kMus.iTDno"�´��� EЬ�(JZ�2�Վ�;�ZEb#�1.m�1��w:��B�u%5�*�7:�Z�hh`�RmZu�GL�tM4a�֤e�,`7*�7i�ں K��is�f�$�&v��q�m2�i�˺���

]@{XB�df�\�J�����]��ڶXڵF:3aeJ��ږ������,J�χǵ157�G����\K�����ԧi�MSl��i��0��1&� Θؠs��KB�&��e6Qܧ
9v��V�������+�T&e��Ga�l���]���c�(i�Ta��J�޼�iS3jK#��]����D�.���i^&2B�K.�,ntl%�h����4	�%�7����k�{XZ�i����#p[Z��ɝc�&��s
�]�Y�,vn�r��aĲ�l����kq2GV0�1-�ٶo7CPB�\-����&��sx�Գ2bk)�Fj6Rhm���]5����[��IlkB��4I��R�ƚn*�0õb�ԨZWY�(JܨQ1f�9����H���lS�˥ẛb%,�WYcy�5�bm!/j%ل�G�r�V8� 1p�l��ƑU��Z�����wwt�w��W0��"�+5�)`E�Pv��&4�F�ڛF]�AHZɵ�!��p0m1��$"ni�b��V�&�&WM���R	6�gm)\�Yj�hg.%ue������:�W&2�)4A!qXLj���n(�9u,� �B �kƆ������oM�i[)x�b�R�ŗ2k��u��I�ho�S���6�2�m@c t�sTҥ��6�-ia�(i�����?���m؛�[��t&hjr��6e�]��\�)u�j`��2)����tA�0�/����j�����R��e�q/#iD�y7ݱq�@&s�	7�Ȩy�N���c@[е��B���ǥ�����'y�g���a�$�/��o�
����=��%}"�>2 ��5sB��ҿ���jpV7g��A���D�2$lo��B��Ƴ��U��a����lX\:N8g�
��J�2p��6v��\!� ��L$�Q� �a�#�#3���h_׍� �:j����[u�8N�`��胼����I(^�ק��������WY�q�K��v[ Z���PYk�.�eZ�����WK�������������&}PL��s8�a�]e	��X�~S2�������A���da�	�^$��ͮ�W(^�=�{.'�퍰}��w��L;ծ�(n��lr-֐R�����q�Rٟ*>������s�<��S�}�;���.g�Z!_CC���&>��W���p�9�3�o�it�gq���ر̓{�]��5'�����܃ ��0d��"F$e��S�S�WK�i��U�(�}�7�`�$�FD��ΏT��*�������o8�A�j�\�n�P �a��D0q�Cc#���F"E�_ս�^���������V��.���>pTנr4,A��AE(�W��L�a�
QTNo���W;<]��n4ѹ�9Uik�0�b��ѐ���_
�|� �0��?�Ccf�w8y�u�8N�b���ƞ��E��qF���$b�����~���d]�
�<L�{9�Z�U��	��_�ܤ
�5�M>��[����
�Bq�_~��D��D���U�{w�ޝ5S}Cf��lc��u�4+T�m�{��.o+j*����݆�<|�njWu/.�f�n{^}��=T<G{kسv���M�P�� {�Ü᤭��ғ����*~{Ҿ�g�"`�#Y��͏p^�7��l3�΁Fcfsw8y���B#��p[	5��:�W�aV,GG�;��GwX����,\^K�B�A�2��Btw~�"�#>&< �����K[K�Oi�uH ����f�)��8uѸ���ҁmЊ�V[tԃ���M{�E��$��5u{ff���){������ٶj� ���(��?I�"�U�CNK���xƀOmz�T+�2�UXP��v��S��������6��>_gJ��'y0D I�b	�T6�F�1̌�Fe��J�����w����_H�H�[�ˋ����7`���IB�h�X/{���Rs�� G���e���|��_��	�cU�0��'e|ι���_I��e��V��j�Vo����Jw�}z�'�yU՘�o2�8�W�B��i�9������b#���S�&P&D��$u��w��a��27s��>��w� �GD�2$o�$�T�̪�=��U^�m��Si5e��F+��� �SG[Z����k
%�u��t�޹>��j�����	�Av�yh4�y,�'Gi�K[��L�]�H�#�<�Bu~� � ���t�l��n}���|:V������2�x��y#b��Ho^;��m�e5���9 �a�$tA0�����`�ѽ�O���'!tGD"E�JdL�EP�_M�f}̫�.}^�f������i�R�����w�dy�\���{�sT-X�ێ�؃H�`�#�D�Y��,dw�tزGK��[]ќ�JY�|�4?wJdL�"U��ugu�[�g6����H�w
#:^T2"��wojV?i����8i=݉�OKPf���ܠGYY�j���*�$I�r��)yߚ�߈@	���{Ez[w�iX7n] 0Z]1s�T���[j��1�s[�P��]cv&2P.��1�7h[
R�(]*�5e+,�9��!��GK]�c̺��M(YM�X�e�n�6��
�dr�K����@���P�[a�Ƶ��s2\Ԛ�K��m,�H��[�+j"��(.%H�\ͥe�(�h�("9��)Z�h�����SY.V34��?��].�k[��A*����K�q��]���Z8�Z[�Y�}=�����@1�a�d��"Dcg�����.��
b��3��yqth�N����2=��%
��"�l��r�l\%4����Z
�T�
��hx���$|�Jy%g.��w�J�K6���b��/"&�v�3wp�"ݮ0�S�<.t������T��e�3��ь �L~2&D��t���eN7 hn�F�V&�C�5Xa��T�;�� 9ʂ�<E��Ѡ��~�P�"`�"$H�[bC���"M]E�a.B�f��"� ��?�����u*��{�i�%Jz�ݝm¤�Au�2���t�:�fYFe֊��CGU�ۅZff�lc���9�\Mږl[�Ұ6���j�,�>�#�5�{ֹE�+�:��a�L�~2 �U�v�fN[u[�}�Q!�˵�)���C�Qw6��O�;��A����F��v[Cf�֨3q�9�{vLͪ٠������^7��ǟ I������;��1���p���T�;��=dBk0�s���~�;3>�M�LЏ35l���a�q������њ}@��fH�d`IlU�T{h�1����x�m
�΅z<I�o�J��S�;9�If���}�c*��ReOh�A��O����"IT�D��F^�%d�Y����4*a���kw�Ě��΅�=��Am�ݲ㻸'���mo�����c��N���
-���e�T��XPYj`�(kD3R;��4�]-�@����AsB�: @�e�ݰ�VK*&R�/Fo;E枔�2,�ӑ� fЯAn�x� �#�I���������X��z=�X�å`M���¤�T�@��L:1_a�ĥ/rҨh8�"�k�� �20��:�"mp�-����J۪��|�;{��+�ݛj���.���s5�t��Z����|M�Ա��j�|�2�t��_m��[)gS�Ss� k�{�@��ߕ�8Ͼ�k�p������: �"F��1FD�~-?U���;��+�� Ș���s2V�z/y���E@Q��j�Z���P	�W�5�&�&vȦ�����س����U�;�If�p#��Yt�@ȟ��(���OV,�4�K�b�͍l%4l��J�uvSL�3g(��bic��Th$�-$;oEf ��2G�h���W]�NZ��N�r{uKs;�����2;���%
D��D�/X&�akD�c75=�0��Ő[Iwd��}@�w�0A��H��gc(����0Aގ��%���P�WP��E����h\]otcRW�X���s�
D�&D�"l��m��Qu�NC  �0���Dy��箲�mY@����ǢoT�Τ±h΍�`�V�F���_k�]�ꮫA�~�7�FQ�)��/�m�W�s����V��#�S|VK���0.��x >D�'6ˎ��`�ճv�7v̑ݯK��U�yS�:k�������^��b�;��3$P���R\�缴�T����r��vF�h\��2�1:�����`�(8Z����B�t)����	�;5�[�	/����J��U�шI_)b�@���n��b-�b	���5 �~�~D�o��c���U�� �0�`�Uu^�-�%Y@��!�С �P�{�n�V�����c+�+�ؙD��$�@Ș ��f��Er���V��Ja,"�gs�s�BkĚ�	�	�@���6�l�$ؼn��4+�	�^�M�|9VӬ��`�J�K �w��m��{�`�_39}$�@�d�a�#��R��h�����!��V���nJ��N�z5��23��M��[ϫ�j��{1�jw^Q�ʹ<�m����Bq;E!:��qX,�m�$��%�h[N�ܵ�����X��Сz4�V����I:I���m(�f P��&m"�֕-��1�$ʺs���l�.3`\�A4��#�����O�!2b73M5�/X� �f�(��t�4��b�䶴��R��5��U
<4��2��it���	�(�Fh��-�m�l�m��T�u�VYe]e�k�m��w�{��C�*mb�`��j�.�k[��vY�m��
M���/l��&aF�n����/��lۚ�c/�V$&�ڄ�m�L�@�y%sm:�x6��1�%���z���b�54=ã[�}��,"�v� .PV���+$(��#�׬��$ld��w#�<G=�Esn��r�	�Y��`�J�K� G)� F�~�n{s�h?&��&�ڠL�da�d����x~.�l�7���]`�<A]S��<s���%���P2/��V��q��r�ϳq_��h�f���>�P�z;����"�gS�^k�
���f��C|�"F �|������X�lYA:��u���
���`�z&#;�P2'��"��хc����,e����m5�.-Y�2��9��2�L�eeb�P�J�RIU�0�^mr �=fH�2.4qw�z3������!Ί�Ӿv�A�$a�D���așv�{�n�-���o�Y�zv�Ǧ�=�z궞����Uc,����@|�����vr�L�\���&������-jjz�^c��d|�>�P�zu{T�>�I�r^��Y���#��΁ ȑ|Ē��xgΆդsM���{Б���0U�iK��jT4A3B�2$�C(v<�=�;�5����CB�΂U���)��VPEЁ�X�R�ϯN̓lQ�糨Q�|�2&D��"���X���N�Ix�x�n�q�"�i���2(@�r�k�M	z���%�>�&`���K�i�=f�.apF����EiYa��t�՘e����G#�6�{e��wl[�ƱC4��%b6���#����u��s;��&D�F(ȀO}ʸs��A�:f�I�0]���WT�K":�9P� �}����o��f�y0A>��#dL�� fV��F��j͕�����w�3������ҷoWXU��So�og:yY��eL���1�벜����WO���l��ޑ��;���k�=�n�{V�VU�����<���n6+t�}ט�w]��۪t��y��R��"�����u�6�l�8�Moh�-\=���wM������zo�r��]���q�s�+��ƌ��cuLkzZOC����I�����W0K����7���7o*�GR�7%ݓW�؈�!	�Փ�o`�u,K]V�jyY7�@�Ev�M�7�-�<�d�pe��,�i"�T�78��^��A���r�����qi�W�V�ٷ�}F�qk;�����Z�'�|�޷71�����L�a��*m#�
�U��F�7�-�ӹǩ����P%L��d&E�R�{�m�0�`̺����C!"ج�xTI��%�Y>�靾\��T*�^��y�p�\;�ַ4o����;-]��Y�����6R*���Baw�a����݆�QH!\��mҭ9ӧq4���
d9��B�r��y��~5.��/�Q�Ia43Y���p��VGmn�2�&�3��ۀ�t����zSǵ]�{,![p/70E�a�[�vel��VfM9�iV�+L��x���Y4�,ɜ�ݡGn��ýS+QՓ[� ��s��
+�.���x7���x����p�El���SH9uw�tL�rS�)�o/1�΢�hZܩ�R�a�ɂ�Jb�n��&rS-^s�Y����o�Tݗ���U_f.�M�;���c��;}�;�
�.��%rv�^h9]��[BΎ�V��z'0��7�{,�a��tJw��r$�M+?��D�'^֓���H��ɲqӡ)9�D��j��i��#��BYg��$	G.p�Ndr��
Di��"q6�t�]�[�q.��' �۬Egk�������#�z�NQHgfn�J��s�Ӭ�y���m�r:�D$Q���8䤜Yi����Ƕ[SMb�Hs��'fs�8�	�:)ޖ�����-�ۤB���M��J��hP���t���`۱ТR����{iM�r�s��݈�������ۓ��3�D��("rA�M�NKm�{d�D��r�93� (�#(j(�  Ow?=yǛ��=0�7��y2G_D�	/����8�cv��F�Uz	6/�h�X��b��IX�җFk�u�TN�wC��?tL����L�0D��#9�wv��Un�z��XqH�L�,~��>�`Io�#.�3����aW�3�:�.�Y�����s����f���Pt���+0n��G������*�g��M��� ������Nަ��ч���U��}�:���aW�`��R0ȑd����+�#��*����Au������.A3@@�w+ �\�*��zwF�㿏��y����� ��	�3��e�������;7�f2I�����o�t� $_I�D�#��ʝ7�I�˕�r�A�ȸnm�[1��.���؁Ȩ{�k1�Dw�߮�8����)*n<,�3��Y	㣮⒮fΣ�����(�Y�pP���t��Un� o6`{���yuk@!$�t�~��ȉ�,�ݻ��x"{dH�jz�e#A�l�6	����~آ�s�� șъ2'����}�x��[��m��lS�M�a�h�&�qv	v�h"���.�h�V�%@��>ɥ��� �?��20�`��p]������B����7�=b#5.w] ݠ�I۪|A2&A�H���=9������|���;���-��j\V����T�0�����b���a�D��;��##$����9:e�`�<�*�}�5�����3S��("`�"`�%PSmP�_C�!do ��t&EFh%gh���E]�תLp�y��n�}���"��dLD��"[���
c'n7�n����h�|�o�)EX��}@����H�����R��~���a�f�Ќ��G[�mX]hr2�������aa���5k�jVܞ�m�"H3����M�{5r���t��T��^<Q����	�����+fh�4[e���U�[�4���*Y�w��G<�5!,9�v՚�֣��F�P�%)�4#�5B��f������3�Y��ٶ�[]2�陪�J0��d���D�2���� �bK����hܱ�vҩ��A�cZ\hˉ�e��p���"ps0�j��0嶳Z��eYR�ts5e�nQ��1s3&��u�@��F;�?���"d�3[6�l�Tˬ%\�I��� C�2�B�"T�t�*��b�鮁�?�����ŭk�����[ڔ���$�G�s��+�&��2>�Kڸ&����\ܞWGD �c���	:��(8��P%��\�@���rzV]���4�Z#�*ћ��;�`����t�g�i�V���ٝ%5�o1�� �;�3$tD�	,0h�U��V�= �0�"s%
�dJ����ի{�!tׄ��c'���:6���ܘ"IB��A��d��'���^���E��^xXqH���P�C�_P��"F��1C[��e�G�Cw_1T�ͰR�˅�[�du
V6⩫�f�B�+i���S�x��1?�3z�|dO���ò�p)ܝ%�53�w��GgR���dt�::��#K`�d��A��xd��پ�H�����sM��&3��^��;������6��;o��;'oh�|�VE&]�Z�-��X1g�/
�{���j��}B�4�L���׸�� �b�R&ň&re����3�8寺y���D�0d�� ��-Ƣ61mL.�_f��n#-8� ���dH��I(Q�}�e<��~��mi[�E`�wW�Ǣ绛4�F��`��8�i�{e�ĝ���t��$a�����'���^�n���/�3KL͖����]eO��Yt�� Ȃ�|��peQEQ�et�khX�D+Z0������������2�Ѕ��`��}@��@o��G20��z�Y��e��L$5<ꗠ'"�4�?I(Q�3�F���v�f]f�������	9�<Y�3*9�`��s�&��}��Q������';ξ"D��IB.A��Vo����E�USC�/:1t��Zˈy
�G2�m$VEX��D-뾵k�H.�Z��(�u>7-S2�-�Yչ�I#�  4;��L�ox���TT���%
2/��D�"IB�z����)�B�V��9�P���2u�S��Z��6x0A�k�Gui7*x%��H���=(Q�0 Ș �%
D5^
�H��΃�R�v��	�ږ�BN��}�#9�-���nه��<�s�3���z���tLM��"�E�3Z�B�j\1 t�-���j�cQ]�B��r��~������?4�&|I���*Zfl��n/�U>7��P�[)��x�x���(Ș"$�ȃY��Y����{�3Vd�Ί8��fR(q���W�� ���Z��蟚��u�
 �&A �L~�P�a��L���l�Ú��z�r�z�K\V�{�+��~�I$A�#1eS �P�n���A&ŇÕ-�6[�7٪���3P7���e�c�J�1�����-OQ�w6Ⱥ�ו���z�z�cVЀ+��s[ؑ�[���\q�V�����x ���}���9�'E��dddh93�-�f��[�U�r�|�9�g�'��2$_I�fv��n^ㅺ!��)�U��#Qզ�]3f�҃f3^�������:�f������A�2��
�șȟ�uh�&��9��؍�X��+�;����m� �#�$0L��%<�%�Y�1�� wUz&����(j�-����IK�������׏�[�X��_WvP"�Bx��&��&�Z�xb��;/v�'���W����}�� �a�F���lX�g֚sGjt�Ol\�����}PLט�|�LYzy���9&,D%"�	��p�<-�l:;�\���P	�k`@Ш�fLv7}k�^�Xdlj�=��Gn�{�A2���6J����0X�S#�#3yk���<(�͵ڹT5zz���V���Jp�\=��R�q��8�ת��+z���j��p��L��O�$�$��.�8rL�a�+,.nLY�lThq�t�b��-�	�W�)'c�ܙf�Z1γ5n.�KH��X�B\b�Vh1���2�D]e��q�fd���&�Ĵ�g�1����lM��0�CA�j$���:�
ք�Մc2Kv�[%dF/vЋ���L��CX��0M���.m�K�f(�M�v6#R����F�jJƎ���Y��~���G
�JbP��!�i����1�uf�U�����v��y����_H�F�#����KΫ�U��]x�	�!%K�^y��ov���c���IB���D�!�|=�yp����2�юjAs@,���B��e�����x� � �a�#���r�)�5�:�����H�"F� l�6���h2��U�!{�^�;w�]���e���(W�v���!I��S�T@Ȕ�Xs���>$���O>Qi���׿\H)��}p�z2RAB�R.�G��)եV��igQ�������}bAIDB�~��H)����կ~���A|�@���Xo{pĂ���r�L) ��)�*��) ��������)Ƕ��S��� ���>�n5c
���̡��t����AHUP��r�RAk���S
a�r� ����[���y��?�~_�;gQ�A+��#��j;a��]��A.��tel�	n�G?�~������a�%S�ۆ2x�H(�,Ă������
A��ī� xDc�e1�R���qٚ�� ���+����{쟞�P-RAa�{pĂ������
AH/9P-�Xs���� �*U w ��C����ƶp_��~�l��כ�J�^K%d��uCu>G�[B�~c�=�3llGF}�C�q�-5�.�Lve'tv_r
[�f6- �f���� bAN��}Ϯ�R
!���H,2x_��ל���y����Ay�F�RP�0��n�R
��1 �0i ��@�;�8i �P�|�x�R
}��� RAeFJ{ʁi �Ü�CĂ�P9�-'��R�T@�߹�o�U���?JD<��|�Y��:��AHT����B�S���S)�9ˆ3���
�9F$�TH)7�W��i�y�w6�y��~��d�) �Q��bA``�Ayځi �C���Ă��A��K��e���d �P>����S%<�P-II�߰�g>�y�{�u���AH(v�I��R�T@�) ��9a��AHT*��(�������\H)�Ü���;*��ﯞ�iB�Q��O������s<���u �����RR��ݸc'�e$
7�bAH)�*�AH4T9�\<H/{گy��������/���3�$[�CCa�[U!lM9q����&��b���t��7�6|�$(d��j��JH,(���x�Xx9�- �Le<�@��z�ȵ�w�F�D|:�G�N��ѐ<!!�=�^�y����w�- �Q
H-wہ�0@��.�JH(R��Xc
H/9A�1 ��
a�r� �T�{��}�g�z�XH/�T2�)������A|�xLr�_}�n;/W�  ܊��� &���@�2$��s�
A JE@���dU)�	�`t�x�%<��Z	I������ �*�r�H8Q
H-Nr�bAL�0�9p�y) �B��X{�~�~�F��9��[��%�ջ�{gn�
Z�Y6:�et7�p\u��~g��<���������SgL󹵕�R�a�Ab���N�b�������Í���տ��2<Ay��1 ��)��p�OIyE�4�^r�a�AH5P�9p� �0)���
H,��|�<>}���J}��Z�) ��?nCĂ�P;���
H,�O9P. ��z�k>���	:�Ă�����H) �����=����~v�1�s{p�yJH(P���H) ��ц$��0�9p�O#) �Q�Y���I�*ok���sߩ�� �B������e�9�'����_x�r*�$P2S�*��) ��{�d<H,<�)���b�Y(e=�� ]�I���Jm~�}gQ�H���]�ƥ���&n�j�Au���h��B��VVt�Aa���k�AHUP�- ���ѿ\H)�Ü����I����y�o7���{\�y��C�����Ry�+���_��m�<e$
;�1 �1����i �C���Ă�0)���) ����R
����y���^�}_��H,=R9E������
��R��o>�[�#��<!���� �v�H8B�A��H)�Ü���/�]o��5 �br�H,1�$�h1�$�!L>�.��2�
Nr�H) ��@��AH4T9�\<H	5D����,o�,�=�{f���߾;�->@���)���%$=�2$)���b�Y)���
Aa�r��� �;�����������}�ZA���Z�끉0@�s�3�JH(P�9E������VU}�u+Xh���xDj�>a� ����1��RA@�{��{�eN��/a?�u��wHT��g/�f���
�Wna:GS��z^�$oM�D��]��%MhW~מ	�I��᭾	$���x�R
Ay�@�(��j����p� �0)���) ��%<�@�1%$s��x�Xx9�-'�~J���U����|�Y=e>yP ���"�}� �,GàxDx���AHT����B���H)�9ˆ3�d����*����xy�o^����o�4Θ��Δf�IP�k��Kv���W.���mb&���$����������c{�B�ݨ��`z{%�Q_qݛI� ܁�xx��Z�/�g�mp�D����O�P��� �a�0���A-�}�Ͽ|s��gs���;� �n���&�ʯ��n�? t���{�z�\xxg�pv�ww�釞ns�t!l;͸��	� oj�M���Fv��#��= > Njˁ��^��.Vo���ك���ф����0�s�[	��0�!�P@7h-�;߹�+9���@����߮�	�T
�< �$� [��PL+qخ����G��@ԏ :ne�Z���*�o���&�@[(s� ���A@ݨ{�X�n����/�/�<� +� (Xg��+����Xh� �0�����La�n�&�@���#��@��>�4��c���b{�ܜ'��c�d�c�B+��$�*�Kv�e��w��9]���)աW�ʡ5b�OtZ��^^�Uw�e����������*�3I���Q��v��-ܻ�*���ܵ�J<re��s�3�Y���u7���]MU�&mk���^91���/��ʪ�ϴJ�gv�H@�ݻ����V�f��P�5�ܜ]֮��Mɺ���J��KjB8�{j+{3Mmf�n�w,u�.��0���]X�/�-��NL��^gP�����2�}�u"��@a�[WwR�V�ΏrC�^�WT����,f^t7�3e>�_p�ݙ�Wݡ0��(����|pV�k^ڱuB�oN�T��7Ӽ��M���wo.�gZ4�	]V��9o��������5��_k9Jln�z/��v�mԧ�fkL�)ܬ�/x7�}jwwW)�B�6��J�8C�t��
6$}��
/�9�!��d�WU�\��;<S�{4N\��\��4nK�c�j���b�X�Q����q���*��Ww;y⻅�c{t�KF��ٴ�s1DU�
�WK�_g+��巳���Sm��!XN��a
7�ou���t�B=��jmHj:�Ī����D�9ٚ���%��^�-͏���ԫ}�å���T�v�nC�R],ww[���&lb�����l���e\����>�";7%�	q]�`OK\�.�*��{F8{��{ss����[��g�IY�2�<�����F�[8<�('�{�v��b��:d��r9T�*Cy�d����x��
����:u���5��2��s���܈�Dd��~l��w�	H,�?�E�8�.:t��H�s��8���ݸ�ˉ@㈼�.fH�R�)N�/;s�̐.R�'9NY8tE�:tp��^���8���nB��p�w"�G���!�և��xYi����=�8�9 �\�S�A8�� R"�
=�t	O���୬�PVfu�]9Om�;��
u�}�u��9���s7C�ڜ����G]����E���o+/O�����:�t�֤�%Ͷ�}�q+I9�:C��ޒ_-8	D�-��z�Ƕ�f��	j�V,`�MDc1�{�W/�
B\͉tɚ��;Ev�-	� X�,�0,�[�YE��%@��^S��knb�STim�n�SL������y�7,"m/�4l����i+[l,с���6j*�p�R%Ke����(M�a5y��p�9,B�4p�1ښ/A�+V��WA�)uH��.���ܷi��쭶h�8�n�C�k
�˥����y�H,��R�fع���s������6څ��3T4+\�[�1le�ˡ�ږ����h�\�!��m�+�h�nљ��3�4��y�uF-�&�l��KhS�H٨����EF�f�Aat)�D�"4�Zْ�.v(�&��f^��u���[v�&�۰.�`�ٶ���R]&�f%��P���b!�����F�ը�ƨ]�,m�¢B하���v`Al�n��)R�㍵؛Ws,nZ`�\��D����a1QR-%SRlR�R�&�Q�U��6��\���s�ҙ-�$$*;ln0�!@�Z뉶i�	f���i�GP�c0XF�6aB�S���u^�XD�YU���`8�hF� �a��m?����V�%��L����. �-CBS]t33K�nX@��L�.6��2K�^��x�
��i���3��b6ҖwQrf]`^+���6p�-��$+r����4���uu�jJ��FX�E2��ѕ&hiX�d�����B]7\�M�lc]p$����R6YpB�k��f�����I���6K�,���j���f6�P��Z�-�E�-p,E���!3��4�����]i��Ҕ��Z�V]k�8�(�/k�qG��)04�4Vm���49�1�3�ܭ���E˗L����7l�+)�vf�v�rE��kn��Ŷ7S��B��s�M4�W3mv��ֻf�M���x-�K3Wd�׎WP�S:���9�F���+H܎�a�{Lcg��K�����k06�Ύ�:Z1�\�s���s�wN�%�=�&�K�]56.����!P������6g]�� d3rf���,8�ruѢk�L�J�Ԋ�me.fn��\f�͡Q2���[-"�Y�4*��u�Ur�B
�����b�]d�dT �-��Yn�t�0��p��-�eIy�%����A+w`����U�*X�a�n�1�+����]�bYr�:��{In̫�hͿ����.�.��m0�V����	�+q-�%�i*Ұ��f�q4@���O��'�����Ka���M��A3� ����/7�[v#� u�<�ޜ�F�)���1�L�O�����w넙ݨ�v��X�a1�9�پ���߯~���'��B� �%�v��"��W� 7> �	���l!�&�����n׍��f��̨���$��KCv�a7v���
� ������V�U�/>�j��I�f� �����`�	��!hMځhAa���v��C����g�~��ф=�n 9O� ����|B˕��AVؗ�N��ayA,a��>������|���������g�X0��� ݠ� �ݰ�Cv�Bn����ʾ��L�>���)��0�;�+�e? w�0�9P�0�M�r n��A	��h�qٛ�����̰]�e�U�Y(;\��2j1rP��Yi��6�[,���bA���m��� yڀݲ���3��ue}%%m�? ��'��[��r�'ф�n�&��X���pv��(�@;_�����3�G��9�wm�����z�R�K6u��mO_��rݸ�����B�N��������RMVov��"=~��G�P�k�>�Be_�!�	���A�� ��=��p�W~�}×�
���ф@�PK� �X�n����/p�����T�{Al ���r�c0ݸBЛ��,7v�/�|��w#>�L���;J��wl�� n@�G��@ڄ�M�p!��ݠ.0���@-�n�0�)��_�{�}�����m�{�B&��0�ݨG�۫������p� �>�{���s�w���ۇs{Z��Ba��`0�a&�BX���.<<L�3�?s�W���� G�]7�g��߾ߞ_�+�� ��	l �[	�� ��P��U�~�[Cכ����;CG�j0X��F�X-�M\љ.Q ���#�J���uy\ �ځ4�l&0�sn�&�@���`�t��n��1ݲ�������
O'k_~��}����	������'�T$���@.0ݰ��M�	l!��`l�?Eo�x��� '> }�w�՟���W9�o����|����c'�p 	�Mej���Zql
�t "�P[(ڄ�ww�n��z &| ��Re��Vj�3U��tv�B椹�]�����*`����T�Չe�/�mda5M�;��|�v�q�h����:[w�<�����g��?sz��¿��l?�$�PKa����	?n���a���+o_��kl'A�\ �j�An�gޞ�8��s���O���} �h>a �>�}��rg�oi0<8G��������7v�A7j i��&�~�J�<�ߓQ�ϼ�π4=j���|��\p� ��@���W�v��MځbF�`�߽N����lʗ���nPd�1H�QL�4���ghEp]4G<�гJ��3J����ٖ*ݯ�I	>ޝ(���	`��}�M��ݯ (<��8̫�~��b~� �@}~����9~y����[?}p��'9� �n�� ݠ�������v��Z��̿v���P,@��G�f���������c���� >�|�
mBX��wM����{����ϳ�CD/ʀX�<��� ���X��\Mݰ0a�3����T>r�U]=�N�*+@=���s��LA�n�&�@��� ��7jL��5~߽��8t@4����(� �7j|���9��/>���9�a_@7������	l!߿w7����ӝպ+��~�+4�rn�wv������/ٙ�Q^�����Bҕ�f�.���vuT׍GfU��uX��&j:*L�u%�����g燇�xy�#"��Ȁn�[#wl&0�n� ݨ���^��B0�ܰ~:��ۭ�=3ի� �� ,� �����n��
� ��{��<��������v��*�N��[L:gs�Ay�,bkF�[vp-���4�w�|���$�쓾�}��Mݰ1�ڀY��7G�v~P��� �>�ˎ�s����=��	���,Bo��n�d`�X��P�0���e�}�=�~/ڮ���yP��!ߪg�{�g:����{��_��l>ayA,a��B�Mݰ;�p���!yPܠ�c���ݨBЛ�����0 3�V)�\+���u-�����w�0�3h�^��CM��ACv��7v�Csλ�֜���	�w�,a>�n� > `|ۮ�U��	����xA`w��L�!����טe���~�!���*Ȅݰ`�D� ����n�\��k�mc_^y�'�����?[�&o���CX�)�q�L��ܼ��ׂ�mU���,>�٩��=�wp����MEb�w�O[93v�Mcc�g�m�<�=�����^�+j�Jc���㊯s�,9�>���/����:h��sՕ̖��2��m
D*���I��6�J���e�)*JgAB2٫Y��e�c��R�\ \�ѮZ]\J:�6b$35��(��n��w8&���z�kL�pB�8ë�� ��B��`�J�n����vu�"7[q@��4uhu
�M���m�[e�	���$vfMHB��6K4ۮ�u�&�KG�\pۻQ�m�J�t�6���1M�[�e��������f�p5��h�JX4h�h��6��Ѧ�Gm-Ah;]�>��<ߞ�����OF�Z����GV$�RX.+2��f�1O��������}�զ��U����*צ�$V����n6V��s��m��}�d����~�Ǧ�L�Jo�J�ܒ��
ݜ�$_n��[�E�Ƣo:Tb��6��;�h��9�;��MbI�[4��9�HS�d�n��wv�շ���Nb������0�Ea�`��������Q�����&Żja����c�U#2\if������X��8�k"�H��s�O`�ܯZ��n��K �%1b���׃��:���;���[ʔ�5�Wy��VT�.y8����'[X�Y�5ڜ�Uєtһ�����r��37=S���l4��Q��S������{V���yo����l�)�W��I1[;�C��9�fK]U�nY��r;���wD��M{����GA"��?����wu{�W>y=�p���3�绤;֬������;b�OÌ�Pq���_r��9���wWt�艮��ޟl�<<a%7
���x�cճỻ����f��(^m������UUH���m�����c�vU+u���
K.��jA���R����RU�Q{$V�Mߑ�J��Cb������&Д�pϝ��+�����;b�OȪJ|	5���c��l���9#!$�]�NW�z�͆�1J�äi�����|��Ú�p]���4/&���e'���غ-�� C�M[�)���f�U�7��sdM��
�?{ƇO�9�w�i�;�}Z�c�?�_I׎8�]���*������^$�]�S�%�A$��3����lNS��ϝhx��$�&fo���ח�357��m��ؾI���I���������ؑS�uH�$R�i�q��앳�ZV�aq�u�lP)�m��^SYXl���{ߛ��43�IZ6H,��װEⴹ���zF��,��^�2I�I����o(<t7^��R�u5(Ii�~8�q�oй��]y���5�Mx��U�J���;=kvꭞ�h��A�&�I��*:�mj��� ih� �f���f+I��
�Ob�<���-��T�8��;�bzK�s���]�T���3���ջױ��xXOV�˯3�g�����8���2`nmq��W���ۤ��I�Mx�Kg~�1�ܱk���3��ԡ%�q���pf|����Bb�͘���W�f3�\�5 :�
f�ZcCa�im-�"�6��>�v/���>+�շ���c��/61@v��@$�h���wo��{zm���d�њ�[���'�����"��j�HE`�C�>���$`IC4��
Gxv%�ζ�J	-;��Ɓ2	4Lh%Vo,��̙>�Ǜ�]{�v6���v�ڱ�0���X+��/-�|��&�&�'6<��P;D^	ܬ�g�h�E-��V����D� � �uJ�F�vt����u#��ɥT�%����miڪ����i���ڷv+Z�ܛ�f[��{Ѫ���g�9gW=@ɑ�+-���}�k�E�j�:4й�M)m�i���-�EQ��3��i�����[C��1�M?��_@�p�ՙn;-�9�XM��fG�,����(���9����v�4��:8���գI�T����P�BZ�u� n�����`���Oh-1�n%�:\��ʻj��� [��M�cVksfB�SZ�.cCD�/jM���1�K6r1�Шh�i��4��S&\tͤ�����������R�܅�*V�!�$	�lֶ�U4��"�P������xkĚjTΦ�J-;e���u��h"I�Mx�&�m�:{���+َ��r�EmS�}�t���Ә�RE�BR�[Q��d`I�D$�me̠�N�U�=/��Awԓ�d���&�$����nv�!5D�iTηJ.5����SK^'A5�s�9G���U@����1��ͫ�y��]v�I�U{��hM�{?}�}��f]����D4���.n[6����*갭��4��)4Rn�|��%���D!5�4�,��j��V�(�7�m� Xi7^&|I�I���1�Cɕ�g�'�,:u`^�H*���n���z�N��U�]�OD��\�V��7�i�x�=�q��g�i���#���?<<4�߀/�v_v�O ��㊽�ƼM㙝�x�Cb.���hh�j6��)h���̧��c<�9Bw{�=�l	#�LB}��(U^�>2I��F����X�j�~��g��ي���ʽ�R&�&��2	$Z�b�wo���c7Q�u��y�ִ��o�'Sݱ�~�2��e:�*�	�j�ak-�3κ]�\�n���\��Za|��'�}~�P�r���˫���;c�bwN��U�}�ӫ{Z6�KI�I��<�e��b����<��j./m38�&d���D�\ol���f{]�I�O�����~��/T�XF����ۡ�suQ��u�.+4�W�zb;w;������w�e]V�`�����+� z�m���=ʫ�َ�t��(�9J�.�V�3�4���W_:5��R���]����k�vbʹƮ���q���vI��[��Ow�2��/���o(u���Vn�:qX[v»qlm]k'��{�Mq�^_bQ+ݳWP��4�~��+eӊ��8�Ua��YZJP��N�؛�xq��b��^G��t7�Ê�],��Fj�r9�{l7�VM�o�->2��n��L#����:�E���7:���ػ��,0�bˬ���Hn[����mW��2��Fȁ�)u�b��!WZֆ�8Oiq����n�o�ڷ��n�yTƇ3��뤭�-�s�
��b�Y=���_KZ0�퓪��ˣ�OOyx��4�{f��?P���S/�]�6�Y?M�qk6���Q΍�|�)]Q!P�{����eT*�r�E����to$ƭ]حεSEop�+0�幝��o��+DVd���VmtG�hg:��߶6��%
�ߋP��B��w%�q]�޷d0��ʰl�3c�vWw���쎫3c|��Y{׊`�oB�s����P����{+������M%q�:�b�x�*�[���֧]��\��؆n�꾮s��v]n�_ �*�ܺ՚��:�D_c6�]��3jB��Բ���.�h���3�bmf�+�f�޾��j
�;��l��]C6���U�|3Y#Y%��?n�:i�X6��'e��)�k��㚺��r��bd(��B�L��r�`->D#GP��9��	ke�E�b��C����n�;ڷ�Ǜ�����B&;YY�vg 'NG$s��O�X��dw����;��%ǖ��9J�{w����>ۄgk���sk^ݨ�8���3�Xg3��8B@� ���G98����]�I���r(8�vb���'t��8��؄����.��ĸ{U��)�hr�G���jN�l:t�n�_4�m�De�۱Αf��	"β�gft�b6Ғ����qw۶�mۜtB�3kR�g���	B@����ւ��9Y�f��G�^Ť�3	�U�6��K�J�i{d�[l��M�[V�2Ѷ��$�����!��i���aeg첔AkUM2
��"UT�����M;��6�画�X�o�	uĜ�$����;'�7�}@�x���%��v�`��⟑T%��4�W�z�s4L�Mxk�-K��S���4A<娨���Lⴟ�'I�I�Jz�/+n�Z�]b�J�`�cE��bŲ�����[w,��+.2(^��t\X���s=��xr�I�k���\����a���;���Nd��\���@�@��z��h{�s4An�jE=I(�W�8�&v��U�3�L������dT	$���:'qbqz�Gg43Y^蒾}��@f�$��"H�=�@��n!�M-�N��+oS���uH��vJ`���ڶ�0�B��t*�Ueʈ��#Q+�]����8/p��!�<�}x��E����N!ڱb���ΉYw�*�,���G?����Q&��h�c믲��疣��m(�W�8�&v�$�+�hwT�	��.f�O~�vp��&DkM��ކ���jb�fd�� 6n�!Ι@�-����0=��@I�1n��ؙ��T�����V��Eo)%^�&�IݚV��oS�͍k����b��X����^&9ì��^:�n���I:<N��h��Xb���ux�&�lrL4��dI'A3�weF�5u�7w�y	#����eV��|�~̑��+{��rà�Nxh��on�V�o�ov�f��*�㦀<\��$A�ٛ��M4�6�"�r���}�U<�X�g���l禫@���wԖN��։��-�K�Rޔ�T�:jbɛ�����|(_Nf�Фh*�4����,�]lGM�n��!f^"lִ�W��e4��D-��\�e��]vL2ҙ�%p�͵�1t̰c-x�Z�/\�uf�j��׬P�n!W]���c�똶�q��Y\^D��ͬ3I�<������i��B�u��FZ̂9�$0�^��@�We�l����L�X�Z��jˮF�ف��KZ�r��tM+���!���ز��u�F�b�Kr`)t6�V�X�i30�B���>�h�C���PV���MN�䛅� �՛��=�Ɖ4L�kj&6�ZQn�y�t���D�.sJ�y��I��c8�����T7� �D��_�z��&�,�b��X�2169�Hđ���"�$��^���g����YœS�9'�ҡMNcx��:k8���P<��I�	4	Y]yT�8ɏ]iɮxP���\�R���g��1'�^�{���O����N�]tԱ�tj���K�cf�Ҵ-ŤWe-�"��t����̒kĜ��l�9����d	��m�o�O&�4	���D���~]��Q^cw�r�S�a��B��b�����]wI�5e,F.փ�0㦢\���]��O{���l�9��<=�%�4�Wڒ
��ŜYꝱ�6�xq$���aޑܨj�{�׉$�ck��e�aJ��V�	����*�$������I.�9������4	�H�F�a�r�!_��z��G	pju�����x�^&}�Mz�Z=Bo5y��b�Wu���iW��hl��ϳ��������6V]�ifΕk�:]��VX�,�%s��*hfin�h:n3��~�^����&��=]d�3<����I?.��=��o&:������{��hx�=SV�ݨ�.��40.H�;6�¾5�#�&�H���L�D}M�>� �@�D��E&7X���*S�w*�6:�k���Ԏ�g�l��3em�J�)�/����[1��ѥ�~o��Czs$7U}���t�P��Q�o����;�X��s�8��T$��&�2=�e�Y����ĕqkʛ�����M���@*��vP�s9y�$�$�1�nۛ���m�y�A�f�WƱ��P$�2	;��N��glJ\�F��<袪�: �Q����q�;jjd�5.�h㉔�dJn�0Sw��yP�ݠ	5�i�IEӼ8R��S���0t�e޳�.���I��y�W6썠h<:W{YXg���2� ��ROٓ��$���H��Łr$�@$�����b��mK/�0��cG�:L�I:/b1�����m�v�sK{�f��P�w�]�卝��������:����&dv���;N��JT���/Eە�vw`�ں�k�O�f	N���щ�jmX���(�Qܢ�p#�Ӊ�g�{���|���W���M I�O�oUP�#,t�4�C�2���&]aeJ��̟k2L�IB3��z��6����M�@m҅r��PS��T�Z����� �9A�������hs�M I�`ԓ�M<7�ʾ5�bx)G�xf2��@k���G(Td�AY��'k�����xR�]7�8��{����\4I�kr�8��&�&�$���ۻ�4łٰ�������d��T�I�y#Y$I� ��;'&;���ʼ	4e1i�g1�NS���.��Tg�G`[ $�@>$׉6����k���-��x���U�6w��`H���"|mYQ*�V�dm����y�v2�{���&ˁ��f�Uwp�;l.����+Y�v3����%S7f��KU]뚌�ӊ�"�r�lc;� h���U2��	L���(K��S&b�mcv��Db�5���e&CL�-�m�(�g����n)�v�۴�5��1u�e����;%4@�m��m�2���:1m�rae��Y���)R��M4LJ[4ceі�r�VQ�t�էde"�:��4�p�X״�pR=�a�c�Zf�^�=|S_mSi�RX[Eu"�h�l������t����S��n�gr�`U�ّq��(��¤�L�^�<��Sau��g��=�4L�ii���X�tq��&�q3���H�J2�:�2	4&�R���qy{| ӝ��M֣X5���N�b5K�S�=CĚ'�9G*]c{�̻7X� \�kĚ�2D°U�3��c%��uM�)��^�ph�j��]�00*� ��#> �AꞞ�\L�:��4��e��7�Ƶ����6)#�I�D��Uv��+�D���,Rqe�g;UJ=��G���3�M����ۓps�(�X��2��t�"T�v�\diF](0�0䋙��I�3E��.���}����$�E��mz�٪/68�aA�#�'_o�H<�Ě&I7P�Ӝ�;TN:�2zR����fm"M�o]M1�[�yR܋m�]!�^j6[�5��_-[�[���0���o�w�O�|��OOY?D�XYF�����k����:�DFՌ�J�I�$��pjC��՜�+K�-+�ˮ;Lz��3�MS�{h��N��Z��D�b\Td��_f����%�tF�Ny]u����	�MxI�Y�YZr��դk�^�秞�Ў�J>�e��щ#pG�S�6���.�����U�Mt�,�j�BͶ�L��T֣X۰��[�Wo}^�Ě�&�a��T���h���Kg�`R�ջW�ƞMhdX3b�����c\Td��K�an�� q�I��sf�'�nPm���&I!��.v�n�=oVrs�×y9q6ww�{��=�w��V1�Trȏ)����.:�޸n�??�Ӫ��e9�}���u�}�BZ��=<�T�WG.��_�'��x�@�N �9ۉ�4�<hk6b�t��\-wu?"k�z��ʍb�ޟ6�:2 $�%���D�k��P"�c�l�Y2�9��po�f��I5�i>�4�������h��-u34Yt�9hf],&\.���l0*�i��N�[��us�f�|���:�\�/g7���O{�Y�������o�2	4&�_F����۠t1��b�t��\-ou1�M x�$��Q���[��|I�M{Ĕ�Ӈ���wvD�������04$׉4L��2\��pT�/W�*����:�^���o{q.�- �thLm;����-�s�u��"�����m��#�#1]7\��z���p���Z���Qa#�/Z�N��$��D$�$cb�H��˥��ά�i��,�I^r�k{��0x���7 �������~3�b�F�,PDv�b06���J�S@�Y��uE!H���%r:9#�2+�%�6N�.�ܓŶ�����6��{7��٨v����@��|m�k� ku��O!;����F�,f��hI*+2l�k��U�>��)#Bgn��r��bo�1z��y�E���&�&I5�MzI������N&�	* ��hS�M�]��&٩�8K�����sD�L�hhԌ�	p����z��tl����@�D����ק���Y�N�Ue�ө���P�Gw-.,�Н�TO9�۶v��g@��,������Zmo}����`���z�r���4��{}��A��6��B���4Z����]�O�u&�<TE�N���'C �G{A��z^l��y�!sJ�tҜ�>$��m�_U]�Qhڻڰ���έ6Őt�̢�����q%�aUGEk����mTv���R�8��Þ5*4lϴQ���ͺ������[&C��.q�!P�o���O��־:��k�(�v{��튔���O7H9�w�HlT�@o�Ul�V/hwf^S�̟=[�Ҝ�)-��//�uU��Ƚ���ګj����}�.��;�-�v�B̓T��R�&�]fnVv��w�g����	ou��1cj����g}̇�j�6�V
�״{L,-����b��ƭ-�-#O��WYQ��nq���5]D�V�@�Y�l��ל�"�L�ZqK�$!�SYE-�O���^�o�v����Y�X�r�K�5�nH^��agnҽ���{�������kE�������{k��e�>Rd�ֺذ�'o���w9���ʆ��7u���m^V.۫[6Y��ל9C;6�V7+,bX��Աi�j��I��]��2����ç���}o1�����w�X�J�P��C1�;��`�}b�g���v���n���(�:�â��N��˸s�#��|)�5]�ݱB���}7�o峯�%�дcʼ��u��7�P�/F3�Y��&�7R���fv_U�Nҷ�@>Ͷ��8袞[βG~ǵ��GNP��I�L�E��wδ�_}��amns�mݶζ���Bp���-��� pq%����d֢f��y"N�9���^e ��<��9_-��;�.�k9IB\-�������:@�>v��ޟ=�ѵe�m�D�	}�t/2�A>׏v_7ky�D��S��Fk�/Y��G��݉�l�[v��l�Ŗw�nr���ͲFkf�,��l��6�24�ݔ֬@�ۦ�2�Z96�ldNt[j[dD_;;�+mcN"HM�]��!|�"���)�h���`�-ƁGHggY��ܲ�:˵�5�#mם؜��^q�V����:7���d�q�v�;�����ז��%�����V6���Z�Wy��:����w�f�[��EС�#�t�WMl�`Q��3Kķ)��lˢ�D,ʴ!B�h�]J������\푖�q�+
��f�Jّ1����R�5PcI]	ۚ�䘛)��b��m.����G�K�Z�3h�f�J\v�
�5�D�X����8�4%a�лkS��HXL��q�Y��%��X�A��uԑ�W8(�4��h�
u�ҫq.�2�4CP�8�is5Ś�(����T�K�Q8�n��m�;0�aAКmqP�앛A`L�1��:���%����l1͑�9�-��\ą,�<��it%��b58��X;YJC	! q���z>��}�6e�Ev�:�cVY�Z������"f,�Ys����!pf��#�[aT�b�fj�6l���A��H�ĳ��F�[|{��Y����4)6Si ��E�\�v��:�ƕ"Ǚ���ڕ�s�����2--���U�f��nfSd��;4W�X4؎i28�R�����k�kͮ�CB�����5��"+)�P�ڭ�Z.;5����Ra�d�T��\G6�رM,+��ilkJ����Zو��mn��X�،΍ժ�Y�6���5��;QڭŹ�б��m�@�R�2�K��[4�FR���1��5��`T�����@y��iCY-k̳]h \bk�m�)�,�,��9�m����)KV�`xH��,S%(�[ ]i�[�f얓gm\YiQnΛ+1	K�(n�3��s4F6hM��n��V�5�j��h����`����FiR��]��=�S�x���k9˨&��M��esI\j1�۴QCjV��Lk�Et�+��)������ó�� 8�4��s	E�Υ�*���KUtٷx ��#��c�37gJ8lܧ.� ���)j#���j�`����t7Vg]�cEF�Vh Pf�l�K�39@p[FciR�Z\��b(%�-�pCm1f��7V(<��X�\�kma�������uf[B]��\�s�rZlX�Ż0c���ݲ�Fn�-����Jb-�rc�b��af�A��]-Ұ��ıXX�.m�]�l���r���T��mP�l貰�!F����
�ƅ��Vb��ֶ�dFi�fX��K.JB��#��8�,�̼A���ō(u�P��-[�h��K5��0���%�X�f��)1nalҎ*�8�2eaP~����4�|��M$%B�mvZ)�hk�r��qm��qFlK��wݎ�9�&�	5�
����y�E����F���+oc8�*I4I�LŠ���D^��r�=T�+
&Ч|�;��GrM�^&I=�Ө���mN�P�>�x�ĈI*�+�6w73A�pһ����ڤ;a�:�Mx>$��x��նF;�}�S�P�{Щ�jSw��,ޮ=ͦ�\	9x���]MgĒL��ۚ����P5O���HS�M�]��&e�"�0$�ޭ}z�J�P"�Y���d;(/&z�Y6��f�KL��2jn�l��Wk����ǵ��$��=d����C�~4F=*�XlY]�I�I�Mz���d_Fe���t��VV�;�ekLnJ�Vm^������3r�o�:��#�]}��^)� ���ѫ0�ڬ���C�p�/��_��7�9G�T��S�r�u�a,ޭ;�47Kzvj��\v6�{�L�I�I��s�..�Jub��Grh�I�6k����&hmLBpa� c-�&��=d���j�C�`b�+R�z.��uUA���<���$`H�"v�T�+��m��Ѹr�u�A,�y����RD!��Sd~�A?U4j�,6-	�u�6��#-v�J0��rG1�F�a4�jn�n��b��׉4L�VTPy��.�]õ&qY�����ג4&�L�pD��r/:�_6�t�%l�N���)�WhvB/���z�+g����mkh
��lH��H�0--����[?��j�<'�	���c���m�~qY~���yy�5*�I��b�h���=��5�˽������(i�9·E�#�
������~����d�D��c�]���/,�vP%�3Xzy�󱲻!wԟ�f�/��a9��H��^�I�I�I/k��:}����%(��|�����E�b��Q&�3գ"�iC��X�c_Lj�E�+�J�9u������� ��K��Wl�W\ٝ���� ̂Mx�A�B�-�J_@Գz���hqj$�5���3�t@IG�����ȇ��Hl�R+���+�p�I�٠I%�α^R���o)�j�	4	�	5��u�yW�WzAj����RX� kTI�x�N<��E����ʼI��*n0��K7������ﱎ�,ZR��]nկi�D.�aZUC���.�|e�Z�b��w�S�X���\5:ɬ�����.������RHٜ�Iy ֞�<�{ܾ����dx�^$�nčO����n]s,��=õ'��{��$ׁ%�E�jzr�*�,k��f�)�2ն��ָ�[,�֑����M{>�y��II�<�H<�e�5�ا�
�2m)��6����$׉4(nRFS��3�i���A�Bv�:��f�cq���":M��w]��Cw������6,��6�ٹ�v��kU���0d�$� �@��$ӮQP�pv����B��d��e�*��S����;�aU����	5�I� �����5��.bf��[ʎ&u����}�#/�������l��9����#8�g3,V�y�=9���u�ϵ�]r����j��*B�5Sû��r���>K0kCyb���7����7���u���[��V3&����j�`�AF�øG]6ں�6a��`�h2����#�m	sy:�Z�30��fE�KA�������4�*�1�pBj(ݭVW�jhiq0ܩ3j(ض#)��ă�a)n�f���-�AsShs)���K���5ՀC�Y�]]
b�`�:n6sB�L,� V`6�d��b)��ڴ�CP�o�g��_�@WJ��i�ci]F��]���M+�C64�p���(�"���}מ�I�����ȥ��wԜ���E����r<y�$��$ҁ�3��%
{��7'ڝz��|a�u������#Y�MsuT��&ۯ�9�MM��2�Q`�+y�❜�eοrY�X��^�I�MMqX+�f!B7���h�L��:JV���n�����)a���2�\i�&{�/S?�Ҿ�aȀ`I(W�b��L}{�؏A������Yܮ�rB���.����H��Աֈ�lu+��20���V]N!��Q��ٰ�bک��+�R͔٢a�
�ᘾ��u�z0ȑ0~�1Kz��	��:��ܗ]��|�TvLe�g�n;ʸ���i��`��\C�;�TM���\z�]fzS��U_�Q��*�6��4t8��]���\�kV^K�Mj|��麁���\�K$e��,Thʟ�G��B�zK�s�g��=ѐo/ǽ|A��H���S��Z]3���-���+ě ���N����{�jz�N���o:ܴr���m#�nX���Dݲ�v�3��Ҋ���U A�#��rJ���yP��c�,������dT~{���wc��ӧpQ�����$�(d�(��A&�<���\6ygT����Zʖ��R��R��H�/�"5��B�e���%#�����5|PEwES��.�+�GN��Kv"��YM�y�0sm�vڑ�A��7� �J�E�"\�wka�e��{+r��eZ��w����D4��0lW�0ȑ0~�: ��1�7{j��� v�G�2�=�.�T�W@K;�-x	� ���Y��N�[�
�m�۝���r�ݼ��G�{��ĚQ�(��*�g^f���]f���N&w�D*�z:�R�ô�fJU��ٮ��70�㕄Y�N�Ф�Y�ȫ\v�_$���H�,G�5p8Ȩ��IB����sn���yo.��P �~�Fy0A2 ����݇ݙ�͙[��=cǢj�d1�ď|��Έ;�2	��x�W � �9bo
����qO?%��k�W@+;�v\y�=�ؠdLL�Z����7ꦍ/�"f��mC�Ě�����b�c��c�v�Ĳ��oЬ�~] S5��j�A4*�x�w�ɮ��0d��"���=w|���a�'6�wwڸ��E���{��zg����],�K�2;�;�u=�{���e3�MA���նj���)��w4!�a��L��tA�F�H�bIA}��+z����<س��׻y��D�v���wp��ճv��ܘT��ȡt5�5R.u��kubh^oT���A:7��p#Й�L`R��$f�^�u�
��uAK8]i=>� ۬�z/����9�P���w||���ܸ�eQ�ZD�3:�\;��M�ggf<��]c9���Z#�E��wp�A3����NDR���)����ם�{rB�v#Д���� �^�My����?'�4&kp��5��ݲWa*ۙ@p��$4nbݳ����T�St�U
����@G���$ؿ=����} ����p;Y���^ʺB*s�bρL�L��{`�:/�0�(��C�V�P���*�f�h#gF��>p���hTef5V0��}����N�Q�LOr�$�+�"g����t"��w�'Pv�]��3v��ǹA�|�fH�$a�D����^����{'�����耲M�h��Roi��;7e��2*��=�:�������I�2 �G�I�u�	��l;��9���Sv�5kA�7�����ƅ�G�ě��d@�U����'�A�'d&��E�xo���r�Y·�uq��5��+&WIb�8�ޫ�N��C[%����+j�ĭ체�v�h��& 7jm]ek�b8�,ڱ�]���V؜�����̅b��e4p��F2�m ����YU�Bh�X����jhj�ݴ���^2��z�̌�
M0��ƃ�mβ:����er1r�`����ݠ�����Yu��# ^���a�k�J� ���A�ѧ��l]䙵�n��e����3e,%i�=Y[n�������?g�J��ǳ�3\�Ͷ��^��-�EZ[u��8]��uO6���h���E�dA�s�S�ݫ�{s3l�z�[]w֙G%l������o�$A�$L���M-���9uܘ�!t�C˕��Z8����}`�����dP�I�~L���J/{z�#����P�Cr@k�M�IPڮ]���>�ڐD��X��yx���i�A{��;�q�z��zP�s� j��n}B	�XTt�pMt����u�_��^��˔�����o��By�D1�����$a�����c}�mX�]ӊ�v�XK�srX��A�(P2&~���=�~����ۓ�վ¯�Auti���
�Wrr঱픎F�a5��z�3weٖӆLj�h���|�#�u,wMX	�Y��%c�]�Np�	��Ʈ�O}F�� ���i��	%
2'�� ��{�W��X�YD����֗�x�7��m\�w1s�Eco-ˆ�Ut������8�twg�4��o*�����w�.v��G{��ml��#�1�r�5x�d��.V��
�BŇ�0G!�::���2!�}$cm�PW��G�����v?V��̼��A>�0A�(Q�3�?��U�.��	�Upqu�'���&��쒱�.���7��bB.����[]��W�v�~;҅|dO��DF+�"7��{U�����3��{����mm��#�1�rw��d��20�&���ׯ��d �a@*��H�مAp����kp��3�؄)6ڮ�c�`�=�>Yn���B3^�$ذ�qwN(�����VZ� ��m�?r~�(���A�$�(dA�)fTt���Mp@nEgwd��q�(��5K B.�{`��;T2�ϱ9_^/�G� ~�8YHgO]f��Хs�PWY��W{u����w���8��a�u�b�V��kZ]z[���^��ͬÝ@�����+��B��Z�j�ڮŷ��T�Ak�]��X*��t�k���k�9b�4�0��J�t����u�t�q�����Bu)f�\᜺��� �!a�+e�N�>�T70+��,��[�������ss���w�;x�S��{y:ͅk�)���W$]� ��y�}��2n�#j���jڼ�8]����u��rK�t{Y�ʱ�v��w����}oF��5Q����֝�����K"�P��˳��iK���W&���N�}�B�P�2�h��]�vݾD�؜��Y��I��C�0�5��VfóBω�Ck����,T��N���ћU��	�p�&j�yd�L�Udy�Uy��o�����hUֺ��U����-�z����cV@M�6�t_��:̦qu_J�7�w*y��S۠��j�"��Y��wq
��}{��TٝIG~��" �D)��L�y����N�Yy�h�{H�d�wo�j�����w3ό���
n���P�|��V)��%,�w�4�7{�K`�������	�5�3.�3�u��柶���K��nV��-s#��G��F-��O(ږ�N�T����hӷ8�h���j�o�^ˏ�����-�����̪�Ԡ����ԭM�(*�z�B[���l�Y��^VJ��ee����Q��qLNܷNn��I�p�/,ə��K89�I�jͱ�a�_Q�" @��;q�Y%���XfVm�k{zfVm�mzvL�efM�(�,�mg	�M���Ӳ������d�팴��b�ʼͱ_+9�}��z����M��,�,�[�+Ί�.���.ƷYfy�wy�J�ٻ(�$�vtt��mͫL��6���du置�[[�::�n���0�㎶�'m��f���Q�qpGg��.�ˆh�:�;mY�Dsn��^qevP]7v�;��Λ��.2�����Ҵ��q�V�yzu�f�ݔ��+����ٖ\g�eYYV^ۉ��c{zu��v9t�w�ei�M6��gV[���u�̝�W�k�ݝ�y�w�6��Ȼ.�N�;(��3\�$ʺ�=p����<�z�H��0$W�"Ȗ�X�7�.�d42xlX�t���۷�,N����)�6�y[>��L��(dA�A���2G�c����ªJ���q�+�p��������	����/3��za��7ٯ�e������Y��`�Ik/+uue��
��pXK��a����~B��f����0�0~�s�'�;�<���͢:g�'�:�ni��0s�����"�A$���PYq�`���zfŀ��C�^��R�6�'�ގr*6,A3����X��R(@����r(�k� �^&A�2"�Ů��X1��Y���f����O: ����&~2J�2.�9�R���@�8��\�_��L�;��=������m۾P �A�u�����C�&!�B�.��cr.��£�:f�"�h�oUC�����R&ӫ}t+K �q�E�m.�]�d���8^w__ϛ�,k���u�`��#�����$�5��O��*���HE܇D�wz�nm�K�9Ȩ㲅�����1W ���͠��0���j�K+a��X�42i^��kcT�:�-�U�٥��S\g����d�����z�.7�x.��+�.����9�t�	�`�D�� ��2��pv��KlXA;�;�������d��Gf�P �A����#ɾh���4u6�N�P���&�M�g�p-2"���c��Į�J���^�A�6?�XA�ȃ �%
t|,�a�#�|�3���;�Z'VVYņ�o��!^t��1��nX?{|� �"�%
���|�~���r���k�w��\��T���$�!�딫Y��yͶi|������5Oo}���B���c�	�KL���w�5���Ƭ�Į��[z�d��l��:l�d�J��J���&ń*�g;��n2�W��P���ks��n�"���������K�����4�e��-)�� �L8͊2�A����b�Ug&�s-�h�C�I���Lf�Ue���+��Gb��7LU�`<�����۬`�I��Ud�XK���]�v2���6� ��F�fvhB�U�c��SA�i���<��i�ڳ&�l�ui���WV�8�f+l�q�10���q�ٱY��������t+�	��@$ط��rq���J�ڻ^\�ؚ4��P �%
����A2 $�@�g��K��{�X�����#�С�o�w���y��t�$����H��S;�t�Ϩn��`���bI_H��dC�߰onY���ӯ�8*��6��	�������d���$_s�en<Bfom�#9Gr@$ؿ>����'Z�Vf�d�=�P�+�Y����g�=}7��{>P̊�I�@�d��uO+Ѳ�{P�ީ��ݲ��Ko�p],G�ub{�
	��P�=�^Cr���{ZN��ٍc1��38a��e��X�n�HM�и�ͦ7��~A�A�~ޔ(�ȅ����}�
�9͢;#��W�H2������#�G���gp�A'�W�q���v-
�z�5V�95T�+܌A�֒���^W/Xy=�2����ط�M��W�c��{G)�3��ֹ���q�[�!��B<ڡo�.�k�����v�A|������v�P��sP`�Ρ_O �H�fH�����;�q���^�-'���Fp=,G�u����q7j�;��;�b_S9��|�t��4��B�rd"����}ژ���z�#�����C��]��@��?�	`"L�� Ȓw�n*1�g�vX�B*�iy��������C��$��XA2!����9�|Q��R��X���R�KRc[v�5�J���Cl�K	�2%��F1�������\�A���	�{'����g�%�Fp=,2/o<���vA�a�F����(Q�0ADU���s�LC52=b���݆�����z�#� W�� I��&��i�T�	�� Ώ�0ȑ3��IB�ɚw�'�va"��c6i��A��d�Տ"��r�GFਜ਼�F�Sy�Y��sw�.�޳��L\P�u�GI�4�
�����͋66m1���vv�]�]�D_{E�3wp�v�F;�X��c�P�+���Ɛ��?����u�i�{'Y�im��K���71K ��4W�LL�Fl�@ȟ�" l\7q7�i�T�~��W�R��>�C�U��2:o�9A���̑�H�b�z��L�pP���.��t �6��ݢ���b�a��6f�[Ec��`��=��&�΁цD�����h��b���]�3o2\��sZ�@�kϥ����J��Q�f�Е#��� �m{���Ξ5/d�=�b�3��b<��XdH����!R�?�B��L~y ��P�����D9U�qzw��0�l3�Wk���3�G���#�� H�H�#δ�x*�5ϒ���#�:'���(v���/k��gfu�U���`��w�l�Mvg�0e]�4����;��Z�_#��n����;��vʺ�w/�F�M�vf=U\*f'�v膸��W�[��uN/��"��3o��j`����$�d��-n���UW"�}�˜V:;ϵ�VFp=,@�	�����'�?%�;{�l���cR����̺Ɔ��R�R�L��ڈ���k�RS;.�i�B���C�#�(P2&A2 �l�\98e���;P��f�wi��¨���X������X��c7v��n�i�ۖ��A�f����h��xc���v�ͼ�bG9�	6/�L��y��x�K��:9����>���̑�F�!��{���Us"�w��c����v\Ubxq�	�?%
Dț9xx3��LQ������2+��6\U.��~�
�Q��J�U�W����:�3���H�"Ee{v�V�>�3Ę.�`��oWn,�˗s�Be
2&AE��G�Q����<��ꬫ��Q���kw�1uk�}U��Z����yUA�[��G�Q��C�d7K+7���� �Z�Bs3)w���Et���ͧ7f�-�.p�6�	��3aW�=v���h�`Z#z�k��|>�+sJ`�6u��sm�mJLݔ	f�,�-VG�n]f�0��.�iX�h#[k�,6z�u��ejVi���dq@���Ƣ��cmkh�V�r��@ЛZ�e/ �9�)�(l�L�#+�-VWJnk�]�M
@@�!a%t!�� �M�c����_�	�Ŗj���3�-q�2ˢ�sf��T͂���n�-�*���~����#|�#�DhW�N�����J��e���*����+�2�٨��J�|̈?��ެݫ�{ ������A�~�����k�dt�=���#a9�b��7���d{��A ���lj�k#l�TJXk'0�۾;�w�gn�^U�� ��A�d�(Ș"�$�(q�����W�ds���s�20�L{پ��ި/D�� ���q�h"��2tף���~&}�d%
�ȩ_�{krs������;��sK�e@G��G�� C5�Iu�	�y��~5��,;%U2j����#�R��W*�m1��qf�ͦ{Y������6��O���a�"g�$�(��ꬃ/�[ڳo.\{"�6��������У�L��?��1FD#F{����k�s��n+����5�{n�$u��K5��4^'q`�pn�r�v�i�&�	u���?v��Ԙ��P�ٌ�ڍ=Z��5����U�$Nr��n{��-}�{���"E�K��i��y�0���Z.�;���K�<~�8Fs;o��u�qE�}����x�A�G���d�� �&��$�A��V�]��#u����(Vv��{]�x�9f�\��T	�}���gK�4�&A|��e}"��$z&jR�XU�����8&r�o[y<���rz#oo"3ݲ�v����.�z�9}��Ov'�n%D��4͊Kn��2���[^ʑ��Mɱ�F�S$��.m( א}(Q�0A2 ��=Z��A��uB;#.��u�|��6�C�r: �������u�n��h�n�nTz7���M;؎v���޼wK�w���_H�mņ��^U�}���{�/�Asv廻s&휾z]�,=R����S:-����*{EiG�Tn�w
��d�Çh�5V��)@��!��ٖ�s�sp[�ۮ�ef<x��{[�gZ�p^	k�OO:#b"g�$�FE�uܨ�ݏwf7�V��e
y0A ȃ���V�;}�m-�K���"� dخ��>�:k�����C�0~�?�FH���'XϷ�͋/�R���o^+�Y�w,@�� �_H�L��C ��(B�Sx�c1���"�p�k��[�p�ŕ$��;f&�-����wL�h��ݹn��	�G��:m��k'��Kl�ׅ�WW����]�1�?I� $B����<׆�A��2	��wع��o���kj��@�"�<�z��	����{��C�l;��Dy����-7j���y^b��4o^GK�Uב	�}�7�u]Ϙ���6P�dL�"���j�^yff^�dh�n�BU�Я^Q��=og��&��%��MU��"�iN3]����8��z�|�Ⰹ�����3����ej�}Q
���'|�ӌQ�	[i�v�]��k�����,���֏fp�r���=�dLL�2$�\/6�H��r�]T��9�ِz��XZ����73�d��`� A��p�n�}��a��m�H�
mH�pQ��!eΚ�L��b����y��tT��l}=��!�/�X�F�@&j=���ӽ�i��W�׮�xB��ڦ3�\0�F�1@�O��2$���ɱ��X��=����@��?��Cjk�.��#�0K^��:�?��g�2��t^U[[��{r��_3�ŐD���a�Jj�_�S�פ�v���d���S5��2�3$T�2$_cz*ȣ��N֍!;��z&ō}&��COZ��ws�#��"9V������[w�Zn�1ݢ�v�wl���.ݼy~o�	k�<�S�fG`��?�: �a�$L�$c@ m�f�gD�f��r���	�'�S�e�m�&���!Yk���̫���x�nfv�Z�Iס�85�;�
���ֶM�W-⭆�ioV5��m���]�F��i�5C�2�9[��j�4$�yKn��Aol�Ʒ�k�¶���2"�t �D�������K�ۡX�.t7�e�
ܮr�O2�����1��)]�V�x&�ß-�)칌�����˩b�Wv��
7Ԯ�=�O@�=HY'h��d;�렬�1ct�W�L��a��!���I�vtd�U��vb
�u25:�mQ�L�{w��^����:+Wl�h�eʖ��:�[�;��覅�ա�M����y���y�0��d��b-Ma�ӏz>{����7�?��y�Y���Wen��F��L�:}�>��7�҆n�Z��n��8���sx-��(��",�����_l�Y"N\k%��Z�UM�{on�ĥz���Y��L]�X�_P����/6m��Wr̊�	�V)���Ud��=ɋ�P�V�s�J/�,M�T���v���)y{��{��ʪƌ��r���G���A���=d���ٺɶ�b{Y+�=T��Tե��.����q�jk<�e����A_]*�|�Zct����YǙ�8_m���蛕����]ǫr�����65-�B[���K�g����r��}Xt�̡�D>s޼�UVQ�~�oR��nr9�:�8:�+�x f�7�{�yb��[,Q�z1�i�b�0��V�͸�-B��'+7ʨ�Ɗ���\m&�;����" �kk���y���ۂ䳢ٲ�:��9��.�ku�g�!v��ӊ��mYVIY�gQY�5�dq�v�ם5��Y�e��F]`]��Xtu�s�u��F��QF����yX��6�;g-�Q6��0���eaNe-�;V��Vn�G)�Nww����n/;��f�m�eGe�;n�::��y�ve�(&l�;#Y1i���kQM���ն�26Զ�Sjʦ��P]�Z�As��Z�E�c.�msj��T�vsn���j�\t]�w6��ٖQ�M�8��3���8�+*˓���e��EIHEnIկk�2��(��(˰�dVtge�mpeXqdgq�q�^]��9�wkZB޲J@��/_�o�}�wV�d�R�]��e�L#4K��Wn6�lXL��5�s
g�q�*��E�NZ�t%c�a��V.r�t���&����)�w�t(���Wm� �*ˀ��l������T�[��{h�gLvllQ�����^����COi�3�eYs�-�RWd�e�U��E!��E��[(f�K�r�-\$Fi���KC4� ����Z2ҕՙ�7�-��1��e4�A�� �2d,��D�CS@�fՋ-�In�q�0E�ѭ�B��uν���.�Z�4�Vd��:�����-!��	6H�MU���M���֥�\�'j�Reֲ��9�i� -l.��SM�u)-v:�� H$ť-��:��ׂ�E�\��L��4�]��`G�:���,d�W4 d��E��W5!����Kt���ik�ItV�YV<�Xh�ĥ�@���v�g�i�H��h�e1F��ZJD��]��v�b�J���k1,���	L�s�J����^6DGY�ɰ��I��Y���تbm	v�
۔�S8�����3b�7X��tc*�AL�.���X`5[K���Hݎ�0]e���c+�HƵ��`�+����()��p1���̸�SѥH�-��fa,��4(����j�ڭ�IIL�i�6��c ��Z�i�*b಻2�s��@D����H�ֹ-b�	,U�bı��-�6Yq6,��2B<ښ���t[[�6�9nT��d��Y����F�Ѳ���3�l��e��%�Q�.�]�1���n3	Ii��-A.��r�Z��h�$Yr�Wk2p-B1%ʋ�q�GD� m^!uh�	�� fYl��-,�Y��d�la1�(�k����{��m-��\:����lAqm� ԁ�c�ș��K�c�km	Jl��t���N�MMa,��`�ד]�nk��!�9�����j�c
�#�C:q�c���n�F;c��^�#kf]	���Sd����v�$�ne�(P�!��V�L�j�K��\�5f^v���)e����[X1r���m3.�L��Ką��;��n�t�� �<�Yt��і�j�Zr��jm�b��y�+����Lu��E[��^a���^�ii���-93�a;]6Kv�t�-KpT����lA�@�V�w[*�l�lŊ���Φ�4�
]��"�Di)3XXJGh��R��i�������n�K��u����R�P�r,�Gs��UpJ;"��m�|?Ŗ��F�<�曯�}^�dV!��PX��WU`�`_�wk^�*%l����{���@�#��#����Q�r��`����;�^��T�a���grλ�~"9���'��m���i�ڠA� �3$t�դ��xr#1����287Gd�MW���@&hG�5�g��QT�i�K�u����P�{ɂ	�=��p�P�9��6��<�@���t��R��Q��A�0$V&H�"��/�9l�����yA�X%���������A�d�+�"`L�]�+��w��`5��K���嬄��50�v�¤2\��ڲ�X�a2��$�j�����A�w�G�un&d�=�=G��0m�|F���4U5~פ��#�3�J�E��A��VV>���	�z�G_o[*��	1��Y"���LU7yR��U�z���Z����v6f�S��1���}=�vP�v�x�'��A�a��7����O%s�&�WӐd��fH�L�{��(�l0Fy0A>�:"D"D��I(=�=����E�؏�vmWn�ʪ^���A�D��|dO�	��1�{���څD�� ���:�3'��u���\�&���GF^I���2�|~"l�FD��"d�(ȍK�
�k�����Y�9��pI��I�����fH��fW�˽�{�.�%�����j�:�yz�6k�c^k2,ҍ���(�,��.�6EUP�Z'{]~�a�D�$�o�V8��޻G���Z�'��Α�4<��W�r`�"H�|dA��`p]���� ����:W'��<�FF��1	���4*2�K�[�7������w����@I�"`������2��=��$�]$�3{y�\��TJ�"u���wV�S	�w��3�!�j�꽪��M�5[6w���_u�I
��)u��Y�Ϊ�����[�9��|(w�dz/��?�C "D�"��/�Ѵ˯UĦ{��fMp��D�4ؿÍND6[��]ԍ�O��r*�6�l�����b�%P&D����?]y����|��[E5����=<�G`�^?t�؃H��$�=���.���z�.�Z�+�k��V؊+��=UI]S:&D&�P���2�M����B���FD�ȃ�]�c3;̷�s�2{�_5�*���z�Bk��;΁H��_����-½�!�R.6,>jF�w�k����b� �������=�#�#A�� ��d��6�ݹpwv�v�.����OV�R�!5�$����tvK����~��H�?$�FD����;�g�z��=z�<��Y�x;k^w���r�$c�� ȦU��]v���:��ؐ5�֙�.Stg������"�O�ә~ �Sa�vf��b��s產WFwQ��s�[��0;���F�H� �$tF,½^U��g���}u�,���4��Z��n�_���r*I(W�D� �mgv�*�y���+
{�j(k��ەkZ�V��2��an�0KL��EPu�- P��x�}�#�D2�������G��n��A�U:�Μ�OS�n��� &��~2 ��ӗ�X�*��yv0�& � ��9蒦Zws�N���_�H� @f�PI�V�����|��L~{�ꑆ�0~"C~fL��*��	���w#UR�y ��dLA�D���9��.�VU:h�<�`��|D�Y�7>�mL��=��\����̇6�RR� Fjg�7}_H�ό�0A�P�d^QLִ��!�P���;)�M�:	/�;�����#��F!*��n���2����!T��q�t�np�"�E�'���wFt�ڭ�`����P�����X%�u>o̚��هMK�����z�����c��F[.aЭM6-��ԙ��7�v
�Ĳ�DjM��%��,5pDam
�&0�b�BS���&v�Wx�Ys.CF녭�I��f�IXkQєM���Ć����ʖ�0,�0�1.Z��.�����fx�͗
45C[h61��ҙ]PW谦���ĸ,R�!���lř�W����\-��GP��f���s���O��e.� im��am�0%�+�6v�s�`��k�[4Ѥ�\^ �ky���0D�������lj���z�_ލ��-�K��fN�d���ߚ���dTM��2(@s�Z�=>��~p����EA��.��`�^ �{���"�fv��v���$���d_z��Q�wzF�B<���j��X$�x�G�H�$`H��e٭�����(@*j= �b�59ͩ}����8�"��*3Xhdguv����s�2 �e
ȃ"E�2G��A��O�Xëy���ܗk�0m/	��@���ƾ�1\y���4[&(��	���hQ�R%3+z:�� h�D�����k��ĻK�L/1o��Dx�e��ڰDu�lj�ZuKڛ�*t]�ȬP�<b!�XC�o����0��?�j���wKky7��En��l�'Qd�E3��p�!��GG`�OTKWb�]��Tr.;������w�ܙ���}�ɘM�5|�:�xW����k��/χ����>��uUK�2z�&��3x�47��hP��z�_��B0�H�#�l�;�!�t��C�i��Wk�0i�<{����2!�|D���`"���V="5�#4X��FD�����w^���.zn0��Ib��Ez1p}��|��s�\]��;�x��e��]�ZUlg����U9���4.��w]g�[I��c�V#u:�s���d}g���,D�JT�1�@�7*�i��R�0ņm�J����3M����@=^!�����#U�97�ⳟ9�M'�bw��7�kj��4��} o��ǌ�
Н�|c�"8[��oV�>�F�+F<w�0�2F�W���+���l�5��C�/"&�]����;n�m�cq��}�%;�ٻ3X%��R��,�zq�}���T��.���RM�f87�ܝ�[��Н6�K�7��2���mi��fp�ٽ���7�,D7w��\F;�������f�G�fא�r0'����#iG-A�i��T��7,@�B.�@*�:ؑe�D�`�w��ڱv�D�ܛ��['���Ɓ���/o'q�}���6z�b�E�2G@�#�v�7/�����ߗ�XϢ��4Ԇ�۶`U����,�̡ARW��l��#rm��<��B�_2C��tdH���(P���Y������^!���_���C~ ���(�&A�ȃ�$�@�"3ep{�&�Ň~�YΈ Nb�(�(7��Ƨ>s������bD��,�@�Ү�y믷�DI(P2/��N�ygZ��qP�}X��'��S��b�dTe�̑�BFH��-7��g�IU�;/�8t*9��x�b��Ƨ#S�Zƅ����ǱȨ�(eGv-��3`���m���=��%�}�iW^��}�=��=�/S�Q���� �W��ErQl�2�� �z Ȓ1FD��̑�����P�7�h����w�$���*���B.�@�ƀ&pG�4>��>m���y�hն&���X�f�L����6�KZ��l[tŰP�9�߼H�'�,���(ȟ�"���]�'�Ed�bl�/e�\�7)tfX��j�P�� c� �d����g��\�B��B=�o���N�k0�몖 @�h0A�(P2+,�)��暎��,��doy��!�$`I~��LM�N�[r��:��~��8�	K����(g#�x߉���h���� {b��2�D�=��m�q��+'+F�2(@��4CE�Ύ�h��y�D� �$tD�0D�v5��9Hn�܈�y�-X��¬��L'��.��~� ߐ�P�"g�� ���i_��+�s@�J܅u>
-�x�ЫZ ��T�qŽ|�p��� ��rm��%+�p黨�µ�"�1/��n=�g�w�̑�qv�F"r��3v03XR�)�pJf�ĵ�6�B�mS�����+��p�]iPH��۶ְ�����1li�ˣ�\M�أ�cV���aÅ���clu5��-�K�A�`��lXV��d��flK������5!Յ�u��Y�m.�ڨj�!U�+�u�!�h��&��.�..�ɢj�fɒX�;h����Q~�f��ֻi��e�LV��x�hl�5�FfM�4ˤ%���c�� � �0d��F�nNt�x���Y��n_��JDvݑ�W�M��M�\c��c�V";�������*�V<�d��a�w�n����[9X�z�;`�E�2GO8��'J��T�`���N���"�%c��9g�o��e#4B}0��R��h�M��ڴ]�,����p�ۇci��=Zqj�<?\0w�tA��B��t�x���Y��nX�&�����W>���C6���dڰf����;�q/�Վ�S�^�_OoNc�H�*p{0c��pFwnX;�x��b g����Yg��j!l 1�D��Rʍ�Q�P�B�H�
Հ�����/��L�F�С�݉�8)�8a;S�u�wK�gt�0ݬP;���0D���dN��p��X������]k]�3c(���jU�{��ŀ�bW��]�w��wT�^��x�ܙ��Ʋ�fFf��L�b���y�&�mЯX�1�&�*`�U�����t؃��*�;�TG�=׉yyeظn@jF@�I�pL��dh�^�T�vh/r��w����đ�����H��0D��Fjˏ�=��s��2$L��vȝgX�
�ᄮ��ԇy�'������2�A������."nܱ����^��u%0�BP����i�x���Z��)xO{�~���rJ���k}���a`���&�X��&
�U��h���VW�؍�b�J��(7@�\&b��(Q�8 ��7T��� �t�I�Vvem�˾�Hq��O: �$a�"`�j���:4:�������$�>1:��'i�rv�k���G��k�i�y�2�kn�nE	�$� "D(}zR����* ܯwA�Yu��FP[+MM�8U�`�[A�Qvfv�}u9�6/�e�۸��}���a�����TԳCGb�)72�k�q�����&���҈N�Z��5;������7��)��z32�� �fVw.�K˛t���	wMf����b��f�0lC�\%Ȋ�V�"��`�+5^�Y��k��q�z�1�ѵj�2����~�5-�嗙3q���c6�_��E�n+�WٹyQq�yF�[8%]�Gq�A����nӔ҆!��/�ϥ�)mgQjA\ql�a�P����u�u�q��8;�e�Y�v����7����5f�lMY�n;W�;e�[��y�����&�^Z�צm����yeOYϡ�[�-�R�@�QW5��k;�nYSۊ%�L.���F���6�w�ؔ��.>����o{�+�P�8X/7j�޳_\��v��b\���T�3^
�=Jw��U볺�J�j��[w���	�Dt�%vd���/wm�Yx�k��I)��Z��}���qoj%q�b�����UM�g�9e.)U�`��T��E]3vW
ŸxZ��cp[yZ5^ں��V��M�x�8u������i��N^��"6�*�|�n��U���u��9g�QOS�Ќ{S���wv붪�2]}���7p�)�Rn<�w��ɛ4�p�i�Gu��	�g�V:�ŕ�,�����2f���Emؽ��!���W���l��՜/*�,�4�!g]�$�sf�_���y?"1����UKUH
4W��vvs(�2:ٳ��GAqЕ�R��YgXv��w�í�Y6r(�2��[j4���3��-�t.,�(�堓�6�b��w�M��j;7"�ַln"��^ڼ�m[mmd\�%�gͻ��n$i�Y(�.vі���C��m�͒���yW���99��i�gdD\rI�ܴq��Ge���w���53Y��k�L�&�v]���dSl��+n��lu���Ή���%�k�޶m�����[��+[IF��	���5�h [���������m͸$#��-�m���[�������.w��v�ʼ���۫l[7ggv�i��{^Rw�d�I���L�CX�3�k$mj.�-;+m�D�HD�_� ��
��;5�q�\�����tA��H���$���Wy��\@T��|A�|39n�;A8��,X�F�7�cp!�J_p5� ��$LL��F"jz*;���PJ��.k�L&;Fq�k��o��P�"�B�X��!w����x��vq/mr0"�"��hP6��s��+IH��B b�kCF�?Gןt���F�>~?���F�nG��~������~�r����u��?�v�=��J��A�Ȁ��UꙖ�~^c�9��'|�Cvt�b	�J�H`D�,DoH�@�k�����{S�ҧVGz���>����#���D����J�к�;޶|=�tf�ڦ�����t�("`�dA�$c`���_�_c�HX#b��O:��%<k²�r�]�ܿ@�MU�
�l�)���LDv�*&�����䊋�d�6�y3��V��i�{�mX�2��P7�yE�L2��*�	�[�81�"�7�VgQ��P3]�<F�`��:� dL��$�@ȍ��37�ggpF����Ռ7�!!���`����?�H�Ķ�p���BS_�+0A,�]��Ֆ�"��B�S)ieT���ԷU�e]Zff���������v�0�B�����&;��]wR��b�dh�T����_N_`2 �"IT	�F]���	[�����ڏ"=]�9��g`7,@�	���43�'O��u�&�3�0��(���2;�b.�xDdA�y%�5E�!��[	��A���̑� �&��:�L��� ����ɟ��J;dN���c�o�u/�"1ȯG��e��2�v_�P	��J	�D�0d����e!%�b��
�]��0��K3�t"U��@>�M���vMܰ9N�D�^fL�,����+;g�m]Q���k1�7����h�E.�s�����5E꾬f����?�~>|����u��~!6�s�
�N.�9ֆ,�3+8+K�e���e�ָ�63z�PN
U�I�sK-ŋ��h�2�����)�� �!r͢K�l��Ȑ�]�v+��Q�U��nm
[��"	3���e�̌�[-�7+֖��\;B���X���sD����v6S��)�ɭ��Ƅt5%8���+1�,@�L�a�ft�jB�\�Y���}���O�kakc�ʶB,�,�\0Xa�I`Ѣ#��&�1���2ܹ[�*tsj�����Z$wi�܌W�'�rC%����1s1!D^ ��t20ȑ�L���{��DX�����3r��6-q5X�
a0p^�mU/�����@��5���ǻ�֤��ر�@@�M
�j��L����=�lY��0��+3�as���3ݰ��.;���X�tT��t�@KhX�נD4�f��q�'��C%���@$��]��������#$t20ȑ�u�r�Z��z��cuX��0�:3�뻖 A�&��"d"ŷg�Q��;]�F����Y�D�-6�b.n�2� 
85F��M��UAS��H���(qAц��dPѶgLö�w����q���DѰ�y�������$H��dL�r룦�y��s6�
T�t��������K:�5J�:�]GkK;�Q���wC�<;3�6F,�}Vh`]wf�8�9�dы��F:i���?{Ɏxw\o�z��BI��A��a�Mf[S.����)�y] �
��kġ�#%������\��</�x\7��UK�����c 2&&D�J����&��E�k� ��0g���A�F���;;n/{J���&��w���\�-�(���wu}"��~�P����tޥ�p&%��'Ra���Iv F��ω5���#�k�.���/�B�B`vm��(���h	�FX3�8�T�f��]1�ۃ�����}|�����9^$а�ɬTb�V�Nr]wr�y�E����eǆ�qt�(��ȟ�I*�2 ��3�G�"_�~p��0�tm�B�����q�	��8СI�t��������` �z&A�+�A�m�˾�ܐ�76�(��
ʳ����)�)}�1�����,��+y췹�a��ϲ�<9�t�yҴa#��͛�e���0՚ ���w�P��M���G���H�"D=*2Ot6�ނ/�dto�$�_v����:��^�mU/M�?�O���:�\�9b�>�� ����#dA�������R�ӕ�����F0��+3�Cǧ��D��~�P~X�S�O�a��f�@յ&&q��b͐(Q�+Li��u��k,���K.�o��E��#�{���	���'Q[XiB4�c���.��B�uڈH_����H�H�$�Ws��)n6$�5Я@-�|dժاFy�H�ܸ�9��ň&z����#��[x<o���c� �`��/J�P1��7v��H��s��fv����]z�Шϫě�3�\�C�Ǝ˓�{~*}��f���:��5ma�P�<v ���y��ȫ�h���R乬}�s�RZR诉��Ȑ>��6(��Χ�%�yZ|c�o4J�zfi7uk��*�
�r�F�O6vZ�[�ǽ��� �"G��D�?��g	
\+��G��mU��T�P��+��_����$�@?H��^�x�J�=���F�+e�Yk�i(m�XIv����f�́.�n�T�4������: �B��m�B��s�,��u��ut��c�����#�22&��a�Y���P�hG����6�Z����P���A�� Pf�I�/�vu���݂�
��Nt?H�"F�2J.�`�'̋og+6�d�A�W]\���5 �BûR��Չ����q�(�9˜�_�G��WѶdiqm�gj[�����O�2��{X��|�6/���dO�A�ȾrJ��x|	ۑ���i����xj�j�B��w�2y� �^�hN�71����VS�(k�<�f�2�n�C�]h��뤳��Lˬ#�UF�����kdy+0��s�`�f�̓E[�7�}�kR���Z���[H���,Dfá�PiFa��:ZRcV�³�;������m��{�c��b�h�2���49�%��{F*�ɳt���`�L%�b��۹�P�1�-M�P�"]�#	������E8H�P�Q҇&�Q�h�+j�-����dW$��C1GB�ae��p�W���4�cL1ڀ�j�s��*�"�~�O�t��ҁsJ�s\<b�U�p�;u��\]3.�[v��7Vy�4!���0����z3�M���F2N0��+��\K�z+sQ���e
 �_0dL�%W� �\��K{|Ay��'�|�i�24�x�W-��zC�� q�P	�w�S!,u�z�����P9?{ɐI7�g`D!ԫy�b�b��ھ��ȸP��<���#ψ"F7��åI��ŕu��P�^�I���u�M���vӥ�ߗ�h��L����Z�	ؘ"H�`�#�f�0�2]�ød�2{�����ʚ&��{���������(a��>�/-���'�����)��l�i�a��%fnج�S����%Qt�yW�Wb.v�'���wjX�fi�K!way�7�³��uMy�_{��A�F0�2G@�oChy��O���	�9�Y��������e��sP�����z�uY`u�Vq�)�oBUWp���ZOu��ޘ�����/�<�>2j�_Ls�B��W>?_&D���ȟ�5㽿*�>��#�hP'|�H��<�뮡l������ի,�<�B!5W ��I(P2/��̭���[��VA�����AD�]��}n�nz������A��ں���}y�s��y��?�?#��20�"O�|�О�28��|��z̚{Vf��+��_�G�����` �"雕w���
+
i�11�J�FU�R�i�-ͮ�궖�Ck��3��B��<�����."sl�wndݲ���Ź�ի,�<�
wn�-k�����'0�"I_H���N׵}�·�pP7��	�]M�Ҫ���r����@�� ��a�$i��!SE��sa�X���tF"E�K�E[��,3R�Np� ƮV%.�U���YY���Ÿם|�}m�}��\��ǻB+e�����_�?Q"{�L�
�J�n:y��ܺ�&A�it�K��|�#7wwjX;�i������CyU�Q�1W�*��B����9�]���<���@�Y��i���9X�&/��� �dL�P�"��z�K��;�y�����Wqv��64�,Dq�BS�#��0�b©���yM�@��5�j��-аw(nnɬ(<�[ *fQn� ��=�>�U��h
�x�b��&�ݘ��صӶ�/�I��̂3w�#��}(Q�&&E��}"�5�u�[z:���^�u�!:/��Gt��:)v��A�Bj�|hP�HP2c���}��\35��'�I(Q�22+�S�������ɛ:�N
�������A�}�3$tF?��pL}e�z���"s%i���h;��mt�K��`�R��Wb �~�hA�ͥ�Ze��U9�]�,�B��-��CU�VYˠLV%�3�򎸡�7+�ᇷH�����w��0�?�C/���:�Ea�B\����Y�^��W�Ji�,]�o">�&�ˌ��8�\}�o����3�0&�� ���pDIv����l9(5��a��eN�iR�Er�'�?�=�B������g>��Ξ]Cg0�
[���|��A�?�{�D�	,���
�\n9L�Tn����^��ذ���dAa�F"�.��)�&�L�g<A�֦G�꯷�`�$I|A��.�gᗑ��6y��Q��'�s����F�H��IB��2(u'&��Aѱp���49�UR��E�T�X�{�dA���i���%�G���@��v˛�x&����Z�גּ�3�+���ɩ��\~��cu��d#�����$�ܐ��$��$$ I?�$$ I*HH@��BB��$��	'����	'��$���$���$���$��$$ I;$$ I*HH@�~�HC��H ��I	O�$$ I?Đ��$��!!I�d��	'�$$ I4���$���
�2�Ά2-��������:�������   Y�p  ^>�P�8�O}�z����M w���@�� :��_ <� =�}���G��P��>�}.̚i�:
rw�疂ڞG@P>      ����S �4    ��R��h� L�2��UUQ�  L   d`j��T��I( 4h     z�@"Q�      A&Db4h'�O=	��L��:t�S�v�|R�8IA��d��DN�� ЁtUz �%�/�Br�YD0)+ۃ����?���\5C���@H�� �	���"�'�.�KŨQT3���V���c����=��TU׵�,Kf���Ҙ����P��i`����V��0�7S���_Z<~b�*��j�cD2�Q�CI7h��b˺�(�5E�H�2��q���B��eU�*��]���W>�yjY)���h�Skv�hiVUɥ\��ZF^T�b�4�-e��bff���V�N���3 �1I/6:���ʖ�wZ��z���f�$&�]�� ��n��R�B-_J��V�4���Û��7+d��*��ƈ!Z��s���>�&��c."Oڵc���I^R��ZҚސ���ۻدU-�Rtv�ޕ��Rn̹MV�v��ҵMwPVV�wIf7/MU�4'���Q[�I��MM"�/l���[TM��W���]
["C	����B;�i���i�u���I=�A���w2�pB��[t�9j
ښd�ś+2���ik4��t�;Xw5=����!��#�E���lJ�-;M*�l^��oM]*�������^J�6 ���6��K�7)b�ۅ�r�)KFޟ��]\��
Y=.�1q�5�#˳gX���b9W[Uu��5��j�-#�PMXܵp��V�ZǺ�-:o1��t�U9w�Q���XY5(YlB�]˪w���lCs!�Ut�1ʣ���d���БMU;���'�|J���H���2��A����^-n8��*����z�멓Cs�@;`�2 #"V�ڣkk�Qkb�F�H*y��t<87�s�n���_�!����8Hb��l���=7�����܈T�QG��POQ�#��m\O\ދZ巵�&1.t�*�$��uJ�Tև4��a���|��;�6�|�̬��z �ڵ1�bX�X7a٠�_.w��d����{u��ur�j�\�Ҹ���I�/lT���S9Z;Z6]�,|m�xTL:���CF/��wn��_hSJr��r8^I���#Du���S.o��.�?+��6��mSx�J�Li��tۥf�u��|�.c1��=ۗ���ЫW�2�
<��ڽ㲻^�r�]�3"���r�-�cx��ݙ��e�����[�+�0\��f�i٭�Z=W�m7�N�n�g#CS2��w���R�ۙ]׶�����T4�Fq����aY=�)��.�]\e��2�[	
�[��5�����{�w��)�����bf/Tch+�-�y����(�]$��ܡE$���#�T�r�պ��
��4�X3k�����"d��U����+sS;0=�34ͷuV�,�y��N�����ss�j���ح&����%����qmܤ]�Jȹ�T�]����-�{]l\�6l�&.�;1���r@����v�*OD^�-ͫ7��srGwx�?���y1�s���Q�)5�Ҫ������}����V����j�j�t��ɧ�g|����v\n#p9 rH\5�6���&d/e�m�lh�N]�0�6E��z��[1л^��o9cc��<3p��a`��MXY��#�Ũ;XJ�n{�uX�Ƣ��:���"�Gc���z��qu�ڪ=<[���Z�ٲ[��m�M��;V;dndnF)�{�m��*s5ɳu:��[:P�Y0*^ч�sy���m�6�qn˦�b��(���o��H8���[�v�Ƹ��=�nQ|b�C˃Ŭ9-�#��`x�cc�V1Z�9m�����эū"�u��)N��N^m��TxԶdjwz��q��/]�M�rl�zL����ݭ��a�!����Ukɖ���.t�݃v9�x@f��<8�F��7e!x�b���^Mci�a�3euӨ��\x���.���Le�Ut�N�z���7��/܄t�)���3R��#b��FIhI�&��M��]�s|^�u��HM�.�lKLK���v�ͯY{s��m��g\��"�{^.�m��y�v�7�_YΤ�IH�c6(�x�m!��A������]-9z���`��8�p�*��o���{�'�osm�A�Q	Ƶb5+M*�:yT2WE��r��X�~*�ba5��-�C~�a4'�$)k`�sd�z�8�I��-#ؙ$�������/P���w�7c;=p�&Q�p��� F�ɭmk�jG��T1�vB��P�ԡm�o�a����?yqr��a;����w���j��iR���J.���m`���b�x��I���@�U(�(���T�3�3i2;�~��v�q����\}>謄p�^}�:qՙ�@�q�	�۳az�u���A��l�L��I �&�+E�Hi/mf|��/�/�q����*��<�<5=�!�jL�8E��������I/�	
����:����硙�Ŧ��㒘��Xl�a�(I�o)�v6�7�b�?\��߮�̐���Q +A��5���;L3F���?��<��A6٨;�Ү���R�du7)�B���f*4E;���E�gg\���xJ�;���[�x;qV��#�����K6U	���?}���� 0b�
J����^m����m����|=�� ��+���'���A�}5}�?,�l��y�0_+e0����_�m�����8ܰ��d+-�hq��(��Y���nu����.�`��q8�mƤ�
�ja�3Ϗ>{h�����&��QeLs��F�E^֓s�8}����~��� ��}"�/�ɭ� �.��1H�7�C\�L�ۤ�,d~����r�B�ۙ��%���n�Tw $�3PGQ��D�'1ٺȷ�����T�w�t�3��M)�+� �qSy�X�����{1.��q�S �
*�PS1(��u�=�>&��D����K`Y~��l���R��whj�����^�~�(k��bb�(AJ�_���NV}�u�gXG�2	
A;��~��,ג0�b�<�1H��iz�!{O����^�{��Y�O��1՛^�b����y�ɇ6Q�S�o�?��Q��������w��~���%�g���L����-�ޒ���͕ r�u6B�z�_Z��_�pg.����?�~�/~�Vޯe�
-�Q�! ��"#|g{߂Ĺ,Z�W6[G`khpYc�1kß�k�3XseY��m�<!�[�2�I���[Hu{N˺b��DE��-V�#\�ʰ#06+�k�4Zj��S�#-H�L2��7l5e�������S������wtA�=!�Ƀ�� �ߩ�N������#����{z.��:�o�D��I?�@�kuA�pFԪ=:v��$�����ɵ���^n��&. ��2��gk8si�;c9|��ù�ge�n�e_�n��b�"Z �i��7��$�'6f�y�P{��-K`�����a@� F]��u��b��i���e��d���2�ˈ��NP^�����o
ڟ� ��?�q#����7Z�Xּ����0%[��F��o}��J �ΐvל5&>x���^'��Y�綥�,��L`yNqE�2񔜬'+ �yk�	����e,̠FU��k��b�ߜ���-�NF�h����}��'�$�}j�Q$�Y�l�AD�~��f)3/n?Pb\���V]�:t4�aΔM�G�'�I��\��Jr��|G_�%LJ���e^��a�4g�I��5E!zl�ݩ%�<����[�%H��WX��9��B"n)}0ǋ��;uV����F��h�SE�IX4�(���BLv_����ۧ,�>_�#���&���?z'��>����'J�E�z�Ȝ���M�ٗB&��L�CT�uN�\�(Fձ
KJ%��]vp�1!-8Jn4����2��L���R�<O�?���ju{�A�>�)��b�a���ݮ� '�gR;�͂�� t�[�M�U
&_Wk�Ir饌��x��D>^��:z�����=��S��Y/�;�����Y{��~V�b�;(�H;��{wI]�U��5�%�W�&7ѹ2V�(��ң���흝�*��?}�<Ƽ%���".���Y_>=w�q���~@� ���3[[�	���ə#)IB��pV9*�|>�.�1hV���]�a��(��I��R!�v�~&6�B!���Z}��|>1��>?�#�L��3�JJ��M~;��i�ȝ��X���,T٧���8��@�]�T��~P.0�@r�m�zK@�;%� 2i�m�S[ҥ���E����x,��7֗�Zٺ镛�k����^�jQ�z���'&�]�Ӂ{VL�3%=>y[ۘk�9rJ���}1UD����>.�/��{�&DfĒ>$�hv\�LD���"�Q0��I�u8��ח��x�1���j�ػ]NnF�b�v넮��c�f�9�S�e-�e��1��܎�P�5��[��8p�'�'rE�"�;c5���I�":��������'8-�m*ٰ�U#h�W�mp��จk�CX�ZR�f��8%�/qm��9D6�����$1S�	d/�H�q{�I�J�I�M��E/X��Z�i�[UU�H,�ؠ���)"�4�6S�P��U��oki��I¹������-���kY� �x�������^&�B�I�#�-��M! 닪oY��B��]t�{k���]w�p�d^"D�ZB�Ko|q�^�k�B��ΰ�EMj��C0�P+XB�
�首q��ccWk��|/eŢ�h�Z-�A��Z-�n-�$H��7�c{_loY�+��[Zr��k�k���m��5k㮼�8�����E��h�Z-�E��h�Z:w残E�Ѽ��t۪�h�Z-�E��-�E��h�Z-�E��~�u�E��h�Z5�׿MuZ-�E��h�Z-�\�-�E��W����Z-�E��h�Z-�EMk���۵�wmZ6ֻ��E��h�Z-�E���t�]��(���m�A?�W�|�r��$BS<_o��$cx2�#�v��������j5�!UKP��L6ڗ�~���Q��NN�D�I��nv����}��S���ނI�n�[IIVv�q�l�)��������߀��+�����)�F)�O��2�t��Y(7*�!\�8Vb���9�"w�o��
ʺ�4S7a��Tŵ;��`��t�{R���/N˰\([�t���\���7�',�����r��>�?1Ĝ�t���H����<�s08�;���2	������9<{��*nb��^������U�2��Y��I���h�XCDkM�H�xg.��ww�㷎����W}ᤛ,ĉ"�QL��s��uV����{K��l��L�H�m�Y�ڔI���g��Q� ��T�
��ߚJJ2^\&���'�$�E�ښ��ʺr�κŧ])���9뮼d cQvr\5��"m#�w�b�~6~QOF���DE��wm���7���d���6��O���>���	&?�@g��ߝ��6C��V��>PUvl�	�d�^؛eC]���;m�i�I�oHD��j9V?"S{j�"FC.�q=V�s�ݟ��o�N�d���fK��~�g��qנ�c/��	�U<��~ �n�(Ҏk�QԩEѴT�<x��fٚ.k�6��k�=�M��X��،`,"�%�T��9����S�x�ĺ�I{�w�F�|�z|+W���yS�0�ۦ�:�;���\.OW����5JU6�Wt�sj�j9��ݧ�>0�I�jЋ�^��O-���:�n.�,���n��y��8.��ꊁ4�e����Giق��{i.';[�Đ�[�7��o+���'�x9q��8W��ȥƹ#�'9�'!r!@H��QJ��F@���qE�n�G\��Њ�Vg���ˮN�tv��s�:壡���᱘h�M5֥�S,�Ԉ�n�Tܧ1����^��7�mnbq�v��W�������j�Ӗ�1���%"�A���f~��\�s�O��O��7'>��V`-,D��/�}������wn�؟��f)+�~_h~{�M��U�k~���}�g'��S�E^�n%���/u��%�%��[!�\Cu߉l70I������^�|�^����@���M�l�37��s�jK�=�W���p���1����:����C�{�	.g%՘�ܱd�µ�J�����1�Vo-�0��-a��?	*����e���T�ߢ���qf`�_�����cX��!r�q�o�j8�̂�$�b0�e�&)�^)ko~z����޽v��G�/vH�:w����qm�>�1d�,�]o��%��w��}����xLfZ����:��*��8�U.\��-T�20v�#�Ly׿�mн��c�j�'��D\�O]�F���#-UxI��H�Yk�O]z�ώ�z{�ޘ*.�7\I�C�����N"EN@$I����,�)I�����K����`�3]�C.����<�b��}q`������!Z�i����wuO�%��B3��\Z p�������F�9�h�#�--���9�4���w�cI��3����H=�.�yu����_m��g��'Iۃ�o�{i\&3(c��_\A����=����MJ��5[3әJK~̃:�pG��C��C��Ǉ�{i�������ZF)�e�����DxǌV�&��e*�N71�K큙��x	
�!�.T;�F��q�y�-͆�dM��#l�� ۮ���`;��/v3�c'3 ϘM�M���5�'؃?t����3kT2q�VW���̳���vi�m�%�ڱB��x�:N�e�W�oMX�wT��]Jy�oz���逾�p����c��e۷�{^=]}Jd�dȚ4�� ��)��E WU��LB-��-��8��Ǯ�wa3M���n}j�rZ:�N��8mŷ=`�!�/L�Fn�m[nՎ���3Ք(���`VB�gu���!��)^���$n�F��v���&��t[:�0ۅ�ʔų:�SZ��=�e��~7y���ֲc��{^�b��kc+�$@��](n�����j.�U-L�K�Q-/9&�:�q��T���я%���6�:�<̖����5��Q�y�m��O�ނkM����-�.BZv�R\Y��ּ��6�|���@;��*c���c-IO���}���xu_5{ �Y��*�c�1Ic��^}OɅwm;��G���������q���D��i ͬ���9���Sc����X���[�B)���V?~&��^�w��e�G��Q4ג�������pq�S���VEb���j�$�������]�9\��v���;�j��߱D�̶ ؀�R�\�a��M��ʶ��A	[�4�K��$V�(�.�{Á;(]�̡r�.�ټ@��Dyl�(�RT~z;wz��Ϟ<�׏l�h��'��RX��[),H �H��@���_~�&\��M~��ߗ��b��-WE~�a#5�O���ێ:{��_?�/���5�W(,!�0�?E��w�y�4`�	-m��5kw�s�˖?4,�����!���8�E�0[ͥr���;vop�+_u&k�i��D�4�HO}��e��(�)4,�ݦ��8�v
��̥�����N��f��,�B�7���{p`1RL���{��J贌�e�p�&z��.�O��n��w��;^%p)5��i��Trן���jDOI�5�J@f'Ot޻��w9���Z��;k�%jf�۶���0��j�u�ReMA�����:;�zk�C��I'�B��_n�����=�)+<�H4`��F�Ew��vP�KR�~����*<F3Q�	x.��^��V�RM�6��>G����I!�EJ��HH))A%��/�A>_(vEPN�}X��^=��6�����K�Iy��as�㌗܆��b-�~U|����la�
PKD�LPP�f	\�OM4�c|�9ІCK\�?rt���	� ��i�5��Wl�f8� �l��Ԣ�G��=�F�)Ժ�c&�t�Y��Z(r�ĕ���(	b����77@O��y�9��.�� �tW�@? ��("���%-�����'#!��O�|�����`������s��9�J2��*�h���Ohw�!;]KC�A,�`���&_h��9��l�У�%;�*�eX㳡�������0�că������炝����z��Z|o�X=Ұ
��".̼� k����F�j�`ǰ�尝/>�.p}QT��L��E���{W�=��;�s�����0�`�w����= w=�c��]_�7.�}��V���+ᧃ�����ƀѥ����s2x!����C�����G���Z,;�JS���įw��W��d�u\)�_�P>A�-�_s��x������PN��"�k������������u�����;�B��	~h��Y���'��z�6`�b�R�(N��}�A��qu�0��P	�¿Ars�("d2KB��f��B���G�&���I@"'i�\����`f�* ����Z|ЊK	���sV̚X?�	�`�Ǵ�7D�S�A%�z ��"���{�1>���?�r7�r�����ꅀO/`v�"�3�ZX�O=|���O�|�m�N�_��9&���
������C��I�B��_/��&�=�	Kpǋ4l~��_��@�>���sC���1=�zn��@Վ�����r� YKN�ĩ���_#�nP2JnG�T��q��A��/Ԝ��<�&{���Lx����X9ׅ̦�<�
!�<������QEw�u0%ՠ��=�H�O�ѳ�6���z>g����xtO�<S�D��9C���.0̴.�C[�d=ֶ��$a(x?�<�9�����w$S�	�5�