BZh91AY&SY���~<"_�py����������  `���)��/� �t�w`��gU��K)jբ�/y�:R��P �
� P J   =  ��
(P��G� �{�hz�N���gBN�� sk[7٭Ǣ{מ�ZY�c�і�&e�dZu]Ӯ�;��[PL�U�  x��n�ݔr����f����롻��ZD᧳<�{��}�׳��a�ح��*��s9�u�.`� �  �c�5���kCp��j�\f��nի�$NQ����y�sw]���͸�ݝt�2ݹ��R�z( 	�琗F鵮�;.�[�ҝ�ٯ3�ýɢ���]]:;a���&ۮە^�  R�;�xwd��������gN�V%��-�9��y�k��v2�[��]��ݹUu�    @     * P(���L�U(� &��  #	�jx"$�H# LF#  &�hb*�FM���`�2h� 22da��@��Q�  �   L��$ �2LFF&ML����2C�jjx�*$@Ԫ��=D�SF�0!�`�����>�̽!-AxQ�%QP��-y{ի�u�FL�Y�w��H��Y^C���4
  %O�C����  ���P�G��aiAp�B�u!����E��ŽS2��_���	,G�I<,���I$�S��U �C�����?J�?���F}��ӏ���a��-��(���4o����	�>�����;��o�﫾��j��6A�$��'��V�e�|&u`K�wN�!�e���9�=�q	���dDhlD�Z'�l,��Wcw9m�%��S�Ϭm�<��ov�܍ݫ�;��S�W����Y�7��#�iO�U��p5>��r���=�W���q^���yzY3�l������m�X6�W^O|���E����ַ<�b�۱Q����[�%�SCu�y{����;���o'M��]"A`�-��<0���C~3�i��;}�����pߛ
@��N�Z���4]9u�$=qs�H;�\^��_x���xw	��.�3�p9E�9S�w"�+}VÙ}@������/`�!�Q�����|�e��с��T�gQ�KG�NA�]B�p[�+��%���@��O8/H�\%x�ZT���j>Nb8���S��0���W���{��
�9d�*@��K|��/6�,x�O��Z��h+|ؼ�k�`�ŏ0q��ߵf81������
 �q���I�a�� ����G�J
�*h�9pr�}����pg�������&���<2-�E�՜�z��g|�f����z��&�4��f�2�}�x������j�њG�����Y�n��ޒ��Z<�<��7Ŗ����3�y��3~Bpڝ6+���dFY��m�2�b5g����능��u�Kq�6ud��pp+8�g�t��O{ҟ�}F���8�$�;f$f[;�Kً��!���<��m�q:m;��w\3�p�.���z��ѝ'���|��yV��B��t��!�o�q{��Ot��&T���&tnŜ�����^u[	t�غOE��xFK7�J4_N��f�ӣ`48�z�Q���t��P��\3��g��2���o݂�_����xJҧJ�����#�؏gD�8L&p/U��9�4|5�K���.s��� ޮ����v� �F;5�sC�`�1ݻ���-δ�xp�ӏ��a,�@'A���v���⦎sC=0�����9�f�� ��B��Ɇd(�c<2��j�j�x[+I�3�w�3^{~`�S���H�mԞ94d/ ��7g�s��O/�Wf���=]�=�;՜����+ǓǓ��'�:��]�{����|f����bXK4^�-}8�8��_N/�����ح�}�6ud��pp(&vw�:8�O�'�珯zQ�ҹ�R�4����G��2�=�T!��N�i�l�&w�(�^γ��$����t�>6f����x<����R�I�|{��_�x]��b!�!�S��k�D�A�qU��/_du�=-��ɕ��m��>ܖ{��@ܭ,T<V9Q��Cb�7�o���I\[5�Ƿ�Y�u�������Ә�_F閧*Y*�/g�W�V�����V�G����d�U����U�v:<j�ӣ�i�za�=G�ȝV�t��͋�+�ڡ7H�V�u���]�7S���aR�%_�Wr���z5��em��i��{��x߮Mw���vN󣶏/��]v+�zx�����������)�S�(���ֿ/��-yS	]��g�ڟ;a����ᵞW"2��/Y ��a��O��Z����:J��!>C~{�aѺe�*Y+�0�����������ѣ&���Vj��n��e���k��O�>B��=HӁ�/Exq
��#�b!妏1I�٣u;�+�.�_ÕX��.��P�U0�L�����u�����7���y��[�ֈ���T
eE�8/�ߑ����}�\=d=��X���0��o��<�ᮐ��ѭW�Bb��O>��bb��"������+�Gf�G�<L<f,�ȇ��z��<>9�^�ãg�l�����Խl��T*�:��E�\��
}p�����?%B��o�uj�7L������Ũ�j���1���hʽV��Ծ��ԭ��?/�O�(�W�<���Ǽ�vCF�g�0�ȯb2��v`�N���K����GY��VG$��*yD��=����,��R�m�J��E=�3�B�2v0�+~F�z�0ﴻ=f��wA�`t���|�|�ޞ��4��G��+ּ>��M�|Nyo�]h�Ș�m��bt��Jd���ׂ��	�](���@�<_3���:F�fJp�b1�/h�y!^�*%8>W�<0�����Z>�5��V�������s��`��a�O����,�2�T-S���B�B��)��B�	��Z�y?�>�Z���	��^7�;�5l7>�Ặ�'�?Ƞ�ǒ���Մ�N��-�����,a�,rG�B���yW�o�;�YH!�� BF��i��a��Э���o��c]��z{73c7;��j��[80��\Sb�Եo��"ӑ��?7��4�V��焣��i4�'��8N�Ƶ��k$���O:ugn)�1���������
r�ۏ�5�K�x7S�٣燲���}�{�Du<"t*�ЮN��5�����ϦZ+�-���5K�J�y�u��w��<S}����<��K�0�)b�>̝�Nv�g&�P�۲^��רq��+�����%D�>m/��s��7����ex�CM��|S��2l�z��qo�'�YVj�5��DU�8�����]o���[�S��1rzc���}�,;{��;
ƚԌ���y�\s4Ϫ=�1��B	�*���6}{�l��};�w�C���Mn��=�����Vi�;��z������t���e)u����\'���u�[�=��nB�ϭ.%�ǽq�ͽ��7�qԡ;���������p���6�l�������\.ń�>*��}������I1�w粍%K2��~k7��D<7�����J=j�f.C����їNTWϽ�2���w+��{��3
B���3.�+����	�Q���������׌�{=��k���Tm�uD_���|(P)u$�����z���,[W���z�z�؞��l�3���]��W�����e�iu��n*�-��	���~�����Z�{���D�g�!�f�=�X��#3E�nt��zg�t>����`���0�n,A���b�v�|�?9����m�;��[�{5say��Ҁ'��.�r�Z�>~��zW���B� {ga�|]S��^ā6�q���^h�<{
�c���O��C;�s�y�$(.�<ICX~��ıl�L�Ϭ�~R���RyY���}~��Ƃ��^2}�Ͻ�c�vڜ����ꪺ]:YۑD��V;�Ii��kX�-��j�)ݔJ��z�A	�|y�G�v\��Ǧ[F.ޒ��}��I)JW<Ȧe+ѹ���}*�`�3��Tc��KX�Ψn|F|��GX�W���t;-��WtˆwE�S�C;O��;��>*���~�W�w$�_E.C���"��_�Of�
������y�7�Ϻ{�M�9EU�/s�E��*��[�n������eg�B���]GaM�=>�ġx�w	ʹ�\���/��8L����+��ȅ������^���Hn�5���X�����ӽ����Yi�U�'�w�b�5-{�1����n7�I��twО�_�)1R#K�t���=3�^���^}�	ӛ����YҘ��y�i.�o\R��F�jvw�O=ǥ��y���ë/ʪ7
6���[��f�:޽q��u��O���t��j��0f%z�d�0�aV���m>��RA.�39�c�t�I����Y�l�=��i>�~�tc�wM���C��ƐC�9�@�A ��4�^�w;w��A����s�G��=�N�e�����w2L��p]�Z�ً��FMݷ:v͸�=���{�����rkJ��Cum]�_� �v�1h�D^*�v����3�ۢ�س<P�{=�d)0�e20Tz��[�.���3���#W��|����a:��>]'.�J�~~����^�OOU
�S��	�*m�4�}�R>E��t1�Ԃ%v���=��D��}���k�ϻZY�][7��}�^��;ߚ�l<C��g�i���V�i ".Ѡ���M�����fu��L�Y�{��{�jSNs��i�e=Ǜ��\T&��������ة��!�̅����7�S�x��RtP�� ��P�S,!������t+�6����z��ġ�2�IӔ�݀�������i�juf�gAQ��S�Ӻ`u�+_j���M&B��+21 7VN�,^-�J���s��ޞ̙c5�f�_w�$)�������g>��1��qH3ɿ���S���E9o�����[��x�O1�ҟM�;K.�����uE���VH���p̄��f���'{��4(<�~+/"N"�9M�MTeO\�uƌΨ���F�m9և��4"�P�%�v/I��|�1f$]*�i�r8
5��;��z�eh�5����{����#k����ϰ��,>?a^3%���褡�ξ���`ON#:i�h:Y���5�-�}q�h�\��Cs�xJ=��`�rL�H�ν����,Ab�y�>��gw1|偏$He qxv��0g{��7�1э����7�����>���ӳq��-�c�3O�9���N=�N Pk��OH��S`����y{��cn�$O�ji���Ṣ�Ɗv�^I�����:��Sز�?��Z���N�F5ܱ���n���id�)�`����F�՚�(꺦3:hɕY3*���%��K �-��Ƞ%�b}���rR�<�k;Y\�۬�v�����7{&�^>�S��d�^�p�����Vv�7:�#�=�;��A6�j��ip ��� �B煏Yǁ;FA����L����4_�n����~��BB�)!o��;�ّ#�O�)�͛/��$��A�O��>�&�f�Q�1��@26��D<��Po�Yיg�V|A�:�\]�`d]�2��A�P�Vq�PmUcr��q6���p�M�q ��#��R\`�q�d0_+
OSq��d��Q'��#d���YH0V��}X�2s��l���6��������!9�:�+�\7�:��� Q�K�(��@�1������" -�M�R��#Q�y�;�*;�t�P�M8DC�DG�Vd�,�Q�nV�s&д5AI���AD��%��\O���0\�B�F�Q��
��p! �X�;Zm���!��a'M�J��+5�o i0�B(RD���D�h��*�!����5���m�r4����D�>�Ѻf>QlKL�B	2Ԑ7"����B���h���2�* �p�=a�����V4A50�D�Q"�A���`��@`E9j@�@�$0�AE10h�P<[�#���!#@�"L�u��q��0آPF�)�	`�D
�[�6��e��k�0���ۏY�4�|�B�J��������1��O*᠅-��F�"��9@�M��L��iTP�5�D��`D�Gs��Z	��K���dY��B�(ŵ�7��z固�����}L��&�Q�&�,}� ����"G���1c`fOH틅��,�$]\-�ֲ���A��1�I��a%!�a!�D\Щ��*%/E�Q���˖�@g-!�LPPCE@a2X"8C"zZ��j� ��@� �s��!���M[(/��?p�e�z@{��!�[��
{�.�ކ�y���롡PN��<P��
э�Dc���1�DC��(P��ep�TšX�1[�f�w�c?�C�>���-����#�{��J��A���\����?��A�?��?��=��� ���Z�/��f~��s��9�s� ��v0  � ����< H@@  �  ��   
  � ���w@0 ���
,�"�� �峜�Y�9\�8  �$ ( @    � ��  x ,  0 � `x� ������ <�9�QEI� yV�s�_� �   �� �  `z  b   `@ P� P  (P0 4  ��<�[�ݝ9�r��9��QzF�����ށ   `� 0  (@<  �� X�    H�� ��  k ��&�����B+��/�s��8����b(��B��c 
 � �   �� �	 � X� (   h� 0  ((G��� � [����(A�/��&�K Hx
 �    `x (D   �  4` X �� HB  4`������	�$�^Q�	D>'���UD�I ���������?P�����20������N;Wϕ��J��Ο<l��ǌ8h�bx<<<%���+J���+B�!Z��Z������BhP�/!
P�V��Z�
�/)B��֡j���Κ<h�Ő�bx<�Ѣ�6l�Ƌ<Y�	��`x<<'�x����Sg����&�.>l0ҞN�/]��T�2!%���JR<S�m�D�<Q��L��Z��I!P�%�D�vYK�����3�C�~P�mI4Ɍ����|L��dw��A4g������`CCf��@%�	��@��L�E���I�Mq�B&�kb�j8 xAH(E�xC�m!L(�}���`�;[R�k�8	2I(�!>���7���)B"�cv˅�%����hP�^� �(�b�M���$�
"|I0�E��%�
�\5B�CM ����FBR+����I��3h<�m%�k�h���k2a�$x��K�X2&d�"Rm.8#���ȹ����X\�G��$�
��f"Da2t��<	��|��+�ə�1�7�K�I>]��33<�8�$�s��7��|y�[���y���S3<����K��}��33������	������{�s}�t�h:((!�������g���T�l�&�B�6�
ղ�B�\8㎶AQ�~b�nc�GZ�X�E��q�� \+�8�0U�Av�� x�rv'!-<P��@�B��.������!���T�"�����T�T�I��^�V���0�.��ݤ��[�j�
�a2�yWF�>�e<c��������q!1[���"K�LD̔���v���g��� Cb"t�HH3�2��6����7MJ���yQM�c3��o)Gz���q�u��0�hټc6�tb���3�(���#�4��<��Er��,N� #���:��F�$X0MTTDSU��L��g)kqi	7V�Ru�!B@�`��<YC�m��b�1���+��RRZ�gG�d��2ކ��蓕t�d�`Զ˳�e�#��r˖�H,�]tQ}Z�YIĎV0K6�$��㉳�B��v�#%�I�11�!!�Aw9쪒��O�����M�z���4� �Am�!��[�ɪ�%n"��@/>%�㩦��6�f0�D�#*�\�i2�8��w�l���$2�-�6K�t�i�LqI	�������).�F\�R��Y$�����M��)�c�Uz�1�k��ұ����/:�$)�T�HcM�Pw
,�WU5)	C&Y��d�]lT�!ZB)ȹ$U�FFQX���.�F,l���ˣ�4���`	�;E��eE[�q�[X�&�4�K7s�7�a�-Z���A���ڦ���Q�9�W6V��u�b܋��\`�cm̄W#���ʛQtgg��ݜ�p: @��D��B�|�R�n.iļ#�Q�yE����cx2w���d�	$)�X�;.Y��{!%��K�L�(�S�y#ԥ���g��z�a\i���B��%���������lDc������F�Gѻ�a�����!anr�b
d�F¶HU֨L]FN;F�tk�T�D�*�j�Fʮ֫�	�R�ܲ-�e��9��Z]���W�J��}�t��IQ��osQ3�mq�g�����Ǔ���陖��8or��0�a����Re���P�)�p����T(�,!]�A^Ye��*��ԉ$�F�]��b���Ъ����=�crK�7tY�(�r۸ܻ�,af�Q*v�U�}G�[��k�Np��83���H_H�b';�ɔ�� Am��Y�	V�%E�&Ό0�BH=`������
"а�hƈ���G]H�Jr�ʋ�)�4�HL$��
gup�]�
,�FT1����YV "Ht�8�t�`@�-2�)n\T�*��@�!J1��	��m�<���3�z��E�e#�t�v�a���[�젽%47���)��M�o�X���/�;G@������[w�v��b1 be��0,�vpv�����ZX��&��,��;���[dK+�$�M��~:�]�K��*�����\�^'�EW�en��{F�PD��#�w��nn��|�96Ы�b���\�u6�,�󋚩DaFX]���8�Kr���IbA�Q�6C��'�#��P��ū�j���W��YW�~_��.N:f/K�q�8�+���q\]/��x�&/�
����l��cc\�TDx"p�;��.8�8�׋8����^���|�W��x��Z�,�����t���<W��UUx�G��I^&����|h�î�'M���|r>'O�|'��	��x~<O�$��c��a�p�m�8�^-^���v�k�ls�Iä����}!�d ���&��t�t����ҺI�s}疐�;��_�I�:H)w��^׷����KM�2N�ut��t�s��0���eT��<�%����#�"���j��m�g���nQ����Ys���N�}Z��*�=�v{5�\Z���=�Ws�C�|R�3~��4d��R(�|3"
�������� ���7��O�{������}��33�;�#���>�ꙙ�ϣ���}��33�;��4�s��Y��r�s��s����Ϲ�9
rr�4V����Ye�{ҜEQE��p��O�:��q�Ƚٛ�V��"Kц%DL0a�(����,��HF�^�P�-�R�vsL'�����	}{�6}0L�m@ⴒB�Y)�D�n��:Z�1�T��S�=`�L�B�T$��tȋS���J�裩a�I��H>�ʪe]�`&
��!t0A�͂%�0ǌI�QlS����R�Rd�QJjun�+SV�WF�a�:�(�����H5jդX���bq�Qcu1wSQ����.�*������6�Wƨ�����T`�Ç�����I@OR:`�;���E$cȎ��c�&�
b�"8nkȩ=����ۃ��"���t�Q�I,��Y) 1 �L�C��ơ��/���ّS�r֔�猰IA��JN��SB�0Rm":c����\0�J,Bm G��0�0�?|�&�K�I��Q	�S-i�P(L�5Z�&������H�.6�I�D��6ܷr���Z�u�1�2�9(�����)bM4��l$�Y$ls�S�M01M0�yi2�)�:i2�� $Cݫ�	ۑ�s���,n�_fd}f���)JH�� 	��w����7�6�)-�ٰE4ĉ����HB%Y��CfZ���b�Ɔ�ZH(@�p �ǖ�۹%�\���tTh�G���P�Ћ	J�r9�wg��$gK	�����&���i��h�Y<�mT��Ks'Z�Zs�L6�(�V�%F��Ζ�r:�6���00�,f�D�)w.B�L}!$��$���1 đ���x�0�[BBȑ�䄳��������x}��-�n�j��wS~nfU����dd�����9�GVQ� �Ѝ)����,%���%��A�
Zi����J�$G���`=IQ�����)l&ؑ��) `�):Ǆl�Mv�Q]�D��b����ಌ��L6ڰ��;1��i���|Z��Z�VI�C"�f�m&�ו(�TK�i�	�'R&��H�;@Y���S|e,9�R:���D���L@�C�Q)"���W�P��*Uꤴ�^SyrI0�R��H����ɟ��s6��)N0$��t�����Fz������m�J$����-ĵ��i�t�u˟C2��%��lP��n���p�j�LV��8�M4ӧ��u��m}f�;��lL�!! ��߫I���blT�j���9�ؑ�R�mˆZ,E �Z�̷%�E�&�u.��L>bOI�6��I!O����у cv�5TJ��D����ˁ���l��o'.Rɴ�W�R�*O��;�tf�Z5�Qh��א���==�v�~���s��ƏVa,���,��,��}]�2G�KAb��LL��Bc��"�b!�Uq���@�BG��n�ul1!v�,���ړ��t2Xi��l��|Ir���&�\�r�.*�v�J�"4�t��2Hr��c��	��Qh���~K�<�x�7952z9͐n�|s���Ӊ�'(�(]���N�L��p�֭j*�g)�@	�C���?k��Z�(թԉv<�:�0�7K]5p6�2ٖ&R��,!� Y�t�e�Yu�� �D'�"yYA(��D�P8/��s��t�bL��㚰�x̦�L��Iє���)t�s4I		f�L7��R@���۳�"�g%��g]Q\�USb�&�o���Y<�<q�UUJ0���H��6J15�߯�i�#��g�<qP,�Y�8p�!f���d��s���m��]�:�G����I���e.-	����ҧ& �n�u�p��膠	������Ze[QnU���E��5�(��<��=961c�#��K5��;�+���l`
H� ݞwNd6b�0\�:z�4�i����Ɲ��E�Dn��[�U�j�첨O�&�cR@��-@(p	��٨&���n��a$��HAH]��������e���6�8�>��S�(�t��&nbT*ISM� �R͘�J���{�ԩ+{L[6MvI��:܇HȑkE����V���:�2����s)Ma��؛N�-��E�讷�	I�Q���*�D��
'�𥒿
?
�\a�;k��6����Y�q�W�����������~�(�~:A��U^2x�x��l~_���q\z���q�8��g՝�c�W���^-^4��ݷ�ӌ�̷���v�|p�O������5��t�6x�?��hz~'�x~����������y��׍1Ƙ��x��/Y���pp�>�d��v?hfŐ��A�j�j�/��q������;~�����k�h���Y�����s��t%��l�{2���hV'X1��P6�Dm��5	=@9��P��H9軻���D����XT���/*�+���d���Τe�OG��y�@
I[-)���^bB��h�$<F�q�U�bPJ�
J��<�%��*���[�v�u��s\E�����B'L�J��L��%Lf�v�-8�ֶB���oL�'�!q��(bG�q6�	��auC�9�Q�8�{G�1��냽�]������Ÿ�q�|���d/>`��,���{.T�|
7d�0K��FK�SX�E3���Z������(�i���)�-�M��aA�GXaǒp'\��W���Z�R-�7Q#+�AM$��LTca.!	�+�'<�"ce�.���ra�p�B�%��8O��q�0�"@j�$��"H���b
�,7����k��
A��c������n�g��8���=�w3<��p|��;��꧗����wU\��p'����wU\��p>��˺���C�|��ɨK�V8i��4߮:��x�y��%�Q�TN�|o���H��j(��$��#E�D�,�y��L�B��@උXl@��!�S!p�0�X���텶���T�!�)�m�{���n�IV2ˤi��R�4��@,�q�d��[&2��i����3�u֥P�*QVn���.��Ik�L1,{a���7ӆ�
+��a��)�B��͊�ZKX�Y�k5�ˊ�ӱw�~���?G�cD'��bő�`k�X|pH	e�!�:> ��u�y��*,�6������Naӳ��u6�@^%ʖ�!$KZ�\�k.\�"��IXN������#Y"r�;�U�朥��}���#[���ʵZ�۹d�$�`�e��I��t~���R�F��2�|�K�M���I�Io9JA6d
���g�*ֳhQc]J��f�Q7c�aZi�~4�� �F�m\ک'Sgx(��󪖪ې6֛M��I��Z����w�B�'��%�P��c�(b�~������p("D� �K�~��+I-$�lM�.�NvS�	�&M��Q�6�"d�	y%�_�tǉI�4�i�䎑��I�Y1�/�6��j�e�I!7�,0ؐ�!�g�.��>�;jV˚�]�)1�JM�'zi(��/R��ïv�`�B@�l5���ˋ$���Q����5��o��ԧ]��#�n<���N�Nb�*Z&���3���i/�7�@�6�t�n��	p8Fm��ؗ�Ǎ���N�Ig<f	���Ā�Yl,���֧-�e�������x��۰*�*w���8�EŔ%(�Ua����bmc���`9��PS�V�ht�j��nq0v�d ;� 0Ǖ�s2"x:��vU˲�mջ��]պ�r��N6�Y�6x�Ni��,i��w'���Ɲ�n�Oy�N%�7�Su�m˼#֓G]��ZJ�5��F8L#��!j}l���dsTS�X��L�ś�ٽ�!{UBe��kғ�K�c yla�_�8o=n�n�zW�a��´��ӊ��5��������Q��DB�r�IӴ~�OttٸH�,Y�/��4��6m���[���~�yǟF&�Σ�hk�s3Z���UQ�uԳ�tQ`n��f�Q
�o]F6�W��Z%��u��J�p��7�s~Lp��0�6��k�RT�[*b�9m�sY�d��2:�:�����!�8Y�����l(�cn�v��*QFS�N��$��L��!��nѣD1�$�,9K 4��7�@��1D�PBِ��lNs�Ut:7Qa��T�q�2",9E\��N%ܤL)XJ1p,�[<Ba�}�S!��[����գD��bD�L�@�M�N&�Ν7C����M�v�+M1�M8��NǕי�ޯ��Wł��O;M{��'��^���y�^^pO~��:�)���d�����,�Om<�2��[Y۰�Sr�p��Kד)��{t��%��J���l�>�t�$�P�\,���n�3O�$�M�}���1�3��cs}�VV���gg�ޫ
�La�g��g���.#"=�ш�0��l�"$(�0�lk� �T�9F�Aj��e ш�rE��1��fD l��"@��p��|s�@�}�*���8�$ī��)�ee��]k �e�󺤒���%�D�)�aa�])�i�a,�H��<�L� ɖR{s2�P�D,T4����M���\�m,�2��dOi����NO�v��%!��M�8H/������ʕ/RN��u �=r�Ӗ�N� �:"x�+�G���Kb䄵Z\v	g�����8���p/��*�ӫ�}n����;;�;:�^�O�*��������Qwh�^8�����_�L��вADd���P��k���@h�8O9���I7�0�#��p3����tː8�[v�b�B��BaUv��+��J�WʫŪ����U��U⫌8�q�^�K��\]/3����Y��}V:f9���՜+�W�W�q|~f��H"t`ä����8?���x�<g8�>g���=Wjۙm^-^��j�t�+��Ӎr��(��b��Tr|���!F��qt;�/�ı��?�|?���>ǉ��w�6&���C�#�W����x�<g�1ݾ��m�mx�^j���\+��x�1�P~/������Ѕ��7�资a�#&X��MhU��cx�z�Byc���9g/�5G]k���,f�MI�Z�)OJ;�������)�G&_���!Ɩ{=�Q� ���;u5ww���Z��%}�44oq�C�v������QKzE�Go�v��#�K7��q�������E��˺�~���v]�W.�w{�.wD@����YwU˻�#_ww��.�wtDk���ue�W.��Jq�aX�8�ӊ�4ֻ�s �AFD�N^׽.��˷F��h�p�P@�!ld���@y�#Z:��>U����~���;�v���FU�V.]9��x�,������:`Jqt�t���d�(��3��I�5����##�B�̟��q�4m�aX�=U,�����e��.<
ʮQtv��=�lt�W57��G���c&���C!HF3��>����>O� ^||��a�U���uCN�y\T^�E����KP�0�/Q��f�1z�{^���c`׮�.��Y1�=�����4��@Pq:��� ƊMv��.�%��Y�{I?��W�⽓qXV+N�ZqDt1J�lx~�
yq�\I�Q-/����	8���KY�2㿢8�����g�F��wcI�T�4� b��֘�c��3�ݡш���7���ͪ�̎��=�'����y"Y2��ԭZЫU�&@����×�3�!��r�Ɗ���Oi9ր�֘��w��*J�T�NS�fӆ]$��i�W�QUE��.�,��3W�� �0d$~�-d0�o%�$/R�k��ә��O��(�,;mXV+M���U󙙉z#�g����P�铷,��e(ޖ�w$d�|�:�i7O5�UB����ˀvPJc��z^���'��).q�-�
5�6X��\��K6����~�Q`M��/`2�.�mۦ��������9�m�}������)�J��K4"Y����d{��B��'[��3��oQ�{,B�
�jf�d�ͤq��aO8�5�6�$!�jD��tG9��`��8 I���t�_�*����~5'��"�Y�tx�5��w�h#�@�����K�ET�n��%�!g�Ԅ�:&S.��J�Q���Y!��`�	f�,����a-�Nf�8�{%�'�/��K���e՜��8��/-�Yt�kb��֨�aܢɴ�#���pܔ��!`�M��=TIR��4r�r�ևM�qO�$�&Lt�r�`��IOqy!R��)�B�ɽ'X��S|�nA,�K6"~;/��]����������t.-p����XJr8h-#Hf������p��H[�"��P�E�a���I8-a0Y!��
£�8aM�K��b�@P�$H �r�[nty���0jl�p�R���H��o��>i���馬>�N@�QM�L]����@3�x�zE���o�p�p�����8 �3�s�X��" �2$Q��\�mcXʭ�dc�JWqY�b��Q���㲝��+�j�:Q:{��KC�V�T�@���2j�u��oi6��A���v��<,|��`�ʸ�Id��2��k f<��`<>3t� �q����,�)0� �o��PɌP@|k��4��p�B�%e������u��T�� D��&�n9�瓣�nՅb�mU����A��q&�`k,�
6q�����5+���j��u~���-�X�o��4��PcӍ�޲z���
 ��5�l�g�T�y��G	����ɷ S��Ä�&�%]:��"DÑ���v�%�%ҀۮY2�l~6�p��!A
x@C �G��d��?�"F,�Yc�2ɫz{C�$I#�Σ�]r�� �eTV��Ky�9d��[2��j��Vi(mL��%12�)��o
K��	��bx���a;w����%���s��YjzTBJ���-(�M��<���bK%����јI`.�|,�r�O\]��&+�v"<�"|	b��F��	��"�*��'�O��p�:]/�x�Ǚx�׊��c�=yC��'�+������O�:*�*=N��t�tOÂ~å�C���+���C�p�=&���Q�Q��آ|(�5�|C��p�<'���|x�G���}��GQ��������'�������8}��lp�����k��?����(�:NO��gI��yk��m\]/5nb�,�\/f>'��'œ�4A}�;٠��XsYp� �V�yL�L��؃e�Ҡ�p�U�&�h�l���w+��]!�h+M�j*i�>L`#ROQ�{�,�C.H�D��5+��i%��S0a"��1.war���Y������P���e(ܝ:�n��e,�b�Ȑ-НcE��T�d�l�LSbc,xs[��k�OwѾ\��V0� RDJ-r*〥��WDzhҒ����b�)2�VT��<(�)(QqU�*�-��V��M1[�NG����u��
4xȼ8�a,�����D��wK����ta6hp��������M�����l�솮��s��i�9p��I���5��i7���xQ8鬆"-3�+�0
��S\�6A(&�m@V�If�3 �j����$]J��KI��%�1��A%$DPD%DP�ض4�!�Ą '�@h)��#3!p"S m���#&;R��Vp���1;��
�-�W-A��IH.9i��XYpğ���w����o��}���z���s�z���z���s�z���z���s�z���z���s�k_w9��ﾸ�/3�8�+�m8�|<t�H@�yU�Xy�i&�V&��#9F���bJ�T��)AV��|a���q��w�
!x��@�R�$E0��4���q𖳄��]rV@�:i���Cf�l����{8rGS^,ʺ7pv�(x�1kT���۵<��䃼�����z�bٙ�3yj2��9C��ʃB���G�^2��NX�@q�x%��E�P$���!t����QĊ�_A81:���ddlf��90�M����GI�+sF���R��kZ�UP�8ˠ6���y�w�F���	�'�@}��ATF�d���^O7K�⤼�)<�e.rS���t]�D+�C �V��~$$�V��GR~�ѣ�oXcᶟ1�l�+H�%&�e7�ѣH������$!.<|�l�|�1c��Cθ�K�hh��K6�[�,^����-�kܴ���M;���L�����}�WmV��]�S�zsQ��-�p�a���Ebw��UQ׈`Ǻ��0�ݰ�+f�v�1ۿy��M�^ V�#d�f���I�������J������'qmo&e�k8�tՇ���sX��BHMc+��L�t��z��$��)���kY�I!$�]&�%�<<��ni<�
y4�N4��������i�T�0ӌ1�ٍ��c���_�"��e�0Y����TZڟ�:7�P0���Z�Ìj|k"�#%R� 8[@� �!Y	�q�A��� !r�B�%$A$Ih^>�`�l�E���I���V�X�B�k��7�B�lv��K�ۦ�i�f�*ɂ;�e�Ħ�+AIm�MYmUa4�h#��K�n8v�k�''�K��c�-!�T���2��2�S.��%C���|��Q��/ʞ�u��~ʪ�٣��1����<Y��N?�ƥ���9�]I$"[^�H\=l$Cg��R:-�*�yD�O�Tr���u_�TXy#�oOX`�����K�$�,D�ԙ!�F\R��8�%6�ˈ��1TV�F���Q�=���-v��ne�m���l� i�W� B	�!~9Tu�)�I�J��%�$���S�+��&��&���I��w��2u�Z��7���y��������e]�(�g�n�킃ǭI��.�N�f����G���o�ߕyש᭥qm�����í�q��{��;x�����1�]7]���Aɩ�c��9(��XO��b��Ѷgл���Kc��+Zr��Yur�eex��[��%�'M�T�B��p0L��\2�D6�$d$>�r����J��6���c&���<;��W.H��n�9�����	�9j��� �!�D!�xW���VJ�B>n)K�	?����+	���!-�C$�1e[lƑm�̅� d�6 ,��N@ �2��F���,�!M �y�l�V�!hl�7_������������c�6��<r1ì�������QUL�t�L��d6�፼�E��7A����C�J%S�Fy,a���0IoʕZ��7U�I%#s�ˉ.%�a՛���2C�F�[kN���u�h���A4"CƈB4�W�]��\�)]ѓs�n�G~��e�Wcq���e�p1����	��q,{q�"_Iwɴ��a�I�ͯ���I$���P�2z3Wlq�#���×?:֖��Hi1Y!���|�W�!!	��&���lK��x�7���,�7E�-+����4��&G�"|t��%�>|"6'�O��oW���q�q_.�ծ1ӌq^8�Ǭ��8�U����U�>"'�O��U���x%�,��~�~G�8�>c��q�/��x���9�Ux�}Z��Ū��,�m�8�G���><Mǈ|>:N���ȿ!��|)����x�������>7��|66}�p���¯
�{i��3����-ی�\]/5nc����1���~\~g�����Du�Fc�����|��B�6�
#J�mY�j����;ٔ��B��*���L���N<l�=��Cw�u�L�>mk�%�8ERL�mv���z)�~>�}����S�<����l�K�0�*��/(ywE��~�x��N$h�H? ���|��`����\<������˺�s�x���z�.�s�x���z�.�s��o�������w7������.�s}������.�w7֕8�b���]��yZ����: �;�>Ua��lMu��d���9�]�':~I�{��D'�n�~.t$�B�F�a)���%��������'!��Թ�I�铽�H�9�2���w��0}���������v�'HhD�l����Qn��,] t�h�D�d=u*��6r�9CE֎�v��2���id8e�f��i����	(�IN�_�r>`d��3�I�/$(�]�g�%��4���,���=��cc!st~��档��c�*�~Wov��BPIp�R���!�Z�L����Rh�X(�cF4N�-V�E1���CM�ޙ�-&X˙d�1�bngl�S�ȅ5\p��N�hSo��)��� B�6����JE!�IHCu����e1X�7^4 �*�tЃF4�E����Q%5�gGG�S+�2Lټ+��NJ��l6�eя�`���q,��U�6�Cҧ!�$<d�����������|VN���~ue�0���p��6&z�M��r�^7Y��/��Y�r4�oM�j:���G�Ɠn	�s,0:n�9p�`e%f~d�e7_�W��}jE�U$��w��7G�=X|�"z�>�D6�U+xI�T���UVo������� B	�4pMqy���hP-Ǩ*�b��V�.2U䙗��9#k(��Z@���r{I����`h�`o�5�G6�:���|�i�����FI��{i�e4��z�G�B���(�3���ѣ(�s|��Y)���U�{^I�A�%���G_�f��]+��t���g=�r_��[x���D�G(�Q��`�/ײ�$e�,[pn$����p�pn�Q�5O)���l�wZOL�a��SIs�օ=^U4F���&R�Čdh��S~�/�J�}�~j�Fraǋ��Ƈ��+���S�K���!r�,������g�;+6�kʪ�4����^	�
J �4�� E�8��#Af�eBa��ڶ+1ˬlI�ˈ�j�M���j�!l5�m��JC��5!%��n���f�Ćy%;<R�!a�X�!%��1`�]<���3���#�p|���D�hH#�p(2w�׾�݌R�WX�U���)j6�5$��b�@�^�s��6pK�l\4�q-�Q������U�Ϩ�؞��4>�>e?!��=�*W��ҚC�K%�Ԡ��Na����Q7Lt2Y.���p���m�c�8��K8M%�{m���z�
tY<|�� @�!q:A���W�N�^T�ݻ'��h�fG^N7���9j��������[�x�4�I�Y��xYv,1fa����Yf^Y�lJ�"]W��ׁ~��1��S����	=
�d�YrrH���۞n���չ�9��	�O�$4"|h�է�F=n�n��95�*�o=���c�s=�˭D:UHP�P��%)�����)	Z���0ڤ�,%�a��c	�o�	��i)��BI�P��2��B9r��j�!`�{&��M�o��?h��B�k���
6"z(�DD���NplQ�|~��	�G�	��2z�_��ӌq|q�����>!тha�T~~!>�_�G�
���W���	?��/�����?/�X⸿8��^M�Ϣ�����Q,�_���N5���3�2�<g�>k���:N&��~8O����x�|O/���<'ǉ���>7���؟f8ʽ8g����/3����\>&
|K����Q�S�|3�����o�v��f����Q�"{+6��h�3���j�#ɶY���׶�Y��\#q��yL��n�w�L�t�ҜH鄽�;cf&+�m�=Kwi��^��j�u��?�}���Pډ��*O�S�)��g.�.^-ۺ3�Bi��*$Y!�&s0�Q��E�A/AҎ������U1D7D=�ŞK�=W�	t����a�XīSX>�v�z��0}��mֈDa�\]��Rxi⭘&9s(0������	a��v�ݺ�������E�f*ǐ�L��Mik��8��F��[X�r��Nyk���ߓ$� P�*T�9C�l��&�Tw+.=S�*��A8����,PNb�Zi� n$S���"�A��0ZN�W���M�EKقD��I�|Xy� P�C��͉�K����Q4�7�	7�'
&�2H �(VS�H����1�Ғ4A�P@�IHX0b�Z���1k|)*����
�g�TD �2SA�����k.��[��˾]�����ꪬ����[��陛����M���33u�����9��{�q�[��8�q\Uc�#�ќ��Tap�����B2�F$�r$��\��$\!8H�p@$��dK�d�tB�j,��Yv�-�.&B5�2�FX�9�N�o�x��t��'\!��C�a��:l��	�I��	d��x| O2Ic�9���c���ZZ�v�W���t��Y��OF�R�Q�����B]��m�3.c�� ��;Z!ٷ�˫�2����`�!�գ�J��4����]4�M�Hu���P�S�J��I�,�n9�JC�N��5Br���Y[�]˶�rԲۺҭ�kq��9�F��'#S�L��Bh+����uX|��-��ˮ��=El4 ��$4"z�|NH��)!�V�e*��N�h@��v�2�D�#�d��S�&���oڢ���I��H��XL�\`�>繿�Gx��ľ�$%���s-��E�I�<���:n��c&%@�`ᤎ�Շ������:"C�&���z��7p�7Ƀf�s��7��p����.��Г��ݗ-��������ke��$��o�L�r7�B�.�j�}^�SCG�.����;�[v��cO�O�����=ڔ�CD8B������Z[��Z�~�Z��-V���0�2r6���8�-�cN>��J���
�0�J՜&(l�Z%��b3m�PLXp@¥��`0��s�2en&h�A7��pP9y�>z��٢y66[c2p�5=&�D��/�$�Ih���J��C�����]�4�'�?T��}$�%����˄�wd%�;$%�87}�0Q҈��&[�Z�����[S�=c����V�qT��*�h[�+V�Ӂlس��W���}n`�O�Sٮ�-<X��#)i�i,r�.�����_{���#�t䔅�0�cZ���%��%'��W{k^�]L�"e�:�FG�\a╥<c�1�Ͼ~a������	o�V�]�]s���~�D����"���0��a!��ê�G�z���ꮷ�?��cl�QL�%h4`�s�R�����>5��U�7_VQtz�eW>]���UYtw��2��r�yGL��,H�3z5�O��(r�b	���C�i.ն�R%Y��]܃I�E�:qD��MY��Q�����/�m��/.�'��_���j��F[\�d���a��BI'C�M8�A�����VO&��⃌Mh��_K7��Z��{!��;c�C�� ���av���Yh�4��mq[�R1.e����"s��҈�C0�$>0J	��!���+M��i�!�R)qF� �P�E���@� �<�9�ę5u�2I��r!p�dR*"����w��l�C�I������x�U�{u�J����Q���Z�QIX �z�q��#}1S���%��"o2HI8u6�7��SXK���}���ݶ��fKi���-p��Wm�ض�L�&^&f
���n�][+�g����jQ���醊(�%�\����к��Ǭ&q��3m3ҺCQϭ�V5hd��\ꝱ��W��b�{7cȱ�u{���wwL�ԅ]*�����G�']Ŏ݄$&K%���B�FG\ǿF:�tl���U<?�W���c�+�Zv�n4�/Ǎxzh�X���	���l>6v�\q�n8��x�>{����O���B�HV�,V�Z���/*B���^Z��Z���<h�Ş ������,���:h�Ş!x<�ǎ�<<<<,dq�YE��ViE]���v���Ha������I�VF�!��cv"�g5��ƅ��ݓs"��'ǻ�dɳZ�[���A<'۳:��2 ʱ�;��t������;��t�w��u�4���A��^Q���%Θ�+֚�˺�8Z��N%[~���ۂK�U�.z^t���r�o��wt���r�o��wt���r�o��wt���r�o��wt���r�o��wt�����9n�)\S�q�c��d�4{�w���8a�]4�ѓ-���pL?�r3���~��&_�ځ
D\b�-[���7��>���?�pm1xH�S���*�M]<x��Pp��������-1"m<x�/FD���⪼c�1��ZKd���B�u�S.�y��-�ٴ�R���Z�%`��7a�Q=��8v��-&��L>��ۛBm2�������mG�:��,~�S;�����U�; ��42�$�q��Z1"$��Q
�b q�t�<&�L�LQ�(<�i�0ڥ'�&	/j#�0�b)E' ��~������fU��'++��>�r�G���Rg�(��w)�/Na:T��ԃ������R��%�$)6R���8?pQ/A$��}�)�?���ffA��/z�
�
1��QD:B���ǒ:��G��J�U\c�1�������!�jűA�#9Xr��B��l�~?{����r��D�p�+���la�Nҵ�OUi;��_�����ݫ��J��;e��2�L��	�	��;���{���ZM�+�I�ٕϹ��l8������!���wvke�̽K��{y$�o�Ovե,o�۸��!�{O]^ �Oլ�5G8��S�q�\n��[%�T�G�.�����*HD�)��T�����U��&��R]3Y$$��=oi*�u�پ��H�U�+�c�1ƫ�5č�u)�1��.Oo�E��S���G�z���C�z�g�$ �RK��-���JK�,QG��n��9����~�#a�>LL�u7�$�-ҍ9}I{�hÔ{W����+ه�I-�HY<�)�N�\l�������$O��?�C�w����5��.J�1�H�CT�u�"
,M��m&�������xXM� )��ei@RH�Mc�jb����L$x��XeS'�Eċ,�D:8+��h+2g�IUX|n�1/�ر-����<��m2X�����&��ɗ=�%UUQ�ӣ��g	�*��i��K���5�����-)nJ��D%����t6{�T�:�i"a�,*�N�&�D��<LԄc�X��b���#�G�4�T���Qv�I�ے���L��7�/S�K�s����`�S�����t'$Q(!�*�� ��Tگ+�ED�xX�x���KZ�Ѭ��Ti�bO-F��w6�Ut�~UW�t�1�C=V��9��pw֋�-��k�V'�
�ēo?|���d������\oy[���;}��n?x�H��Z�g	�%��@���0Ӥ�}�Qp��IR09���Q�$N��!t�޷e�e<
����1Y��:�8�Ý�TzT��ɴ^Q�դSU�'KQUj�k娶�ىr���P�!5Y��L'��6�.�95EUT�R^�r�(���Y�Ib�\�,e�bI�����p,:W����0�x؞<'����|�\qǏ�8Ҹ����ϕ�����N���8��x��4x�<tO<"<'�x�Z�J�!j+R�J�!�j���O<t��4x�g�<A<��h���8p�f�<Y������z�>:Y�Ǐڝ�5��s,�eB�1�"m4df�A�Œ�۫�<3n8�Ȋ�.O��.��I5��:d�"p��(U�B=���n���E0|y݆�qU��z�>խ(V#f�٣H�����JF�M8`������-l�� �k�D=�SY�i���iIv�J+�ތ�f��!H��5�0��)�7��j��{�D��*�#;F �e����cnJn(�</W��N����{@���̣�*��_�^��A��8�g�!-F�-�d��j��=Ɲ\P����_6$�J��R/�7ﵚO�8"���ÂY���1��
��s9��-?����N�e�I#������{�6"-��M:�SE�4�/��zFnT$i06*b�H�M+��hs�`�����ҮBڕZM5�k��J1I1�[b�[*F�B|�VU��*L�SbI#�q�ʉv��D!
a�._d�I%t5&�Z-$��A�jL*�0�`��D0�28
Ђ�� I0�5AI ���AH�	P&�<fAq�"�e|.��D������MS������/��nywwt���r�nywwt���r�nywwt���r�oܻ��ffy����9��{�s��8���Q>!�C��f��{�ɑ��f^`A"!I ���*��A�m�E-�$��aĚ���0����0��a�Bq�+HQ\% �
�A	��H��BOZ���%&Z =�=���@��$�JL'��i5l'��N�� `�,�V���^ч�9<�7d�bHHI�����=�zz��Qb���0�|i�I	����U�k���mUҕ�Ux��>ye@R�@2
д,w�\M�$�T;����� m=�=�'���������y��2c�ε��d�K*Aa ��$ժ�������Q���*�7N�=��]��;Ux�v�����c���9�T�:�6���)�%�d7s�B�q��E�)���ժĢ�X�S)���Z��H��F�$�*�v,���?�F1�!�?iXW�'��`]����^�L�޿2C95���!��"a��:Vb�r�ʙ*]Z�Y��Q�>��D�[��P/mp#$L
*�I�{����?I�TJ.m3O}�|��e��N%\$��ΓNS!�vgn���&'�{�f>�G������5�q�UW�`����!|x���Ǳj8����8�8��'T��%�c@r��[r�0��bn5 F x�1�Җ"`<:p���aBxB�0�Yq�����u��1��<m �D�90��$�_�'������HU�*��2��KT�@��=���=^,�ʕ�ڦ^f���t�c	�	��z�©���&S$c�RBv�iÇi���H��aV�V1��D����h��dt�?}o�N�S��V1�=UWLt�1��^�V.��G�߬�n7&i���!!%&\d�Ixi��i,���ιo��(��D2�R@�I�G���!�u(��5ߤ#"J��,�<:U|�ڪ�ǌc>ǻGj�C��q�Z��<bC.�,�L�N��7L	���Ķ��"cͽ���D���P�B�$6P\�xt	��ޞN�	��m8g���H\L��SU�Ǻ8
]���3��*]8�K��!�<B���o�@�J��6�5UT�4�4�w��И2J����.��3#j��h��tz�l�Zk%D�	\�Q�U�z�E���X�ђ:M%�H9y��ƛ�M���!$ca���ۺ"8�<ZH�	�X;M%b�鬅�%tDM�C�������0q�P�E�F�+EB�|,2� Å�$A�B22!�H�	%�HuHD(1CPB�\��C�i8ÉB��rX���a���J�
�82☘L�����q4ݸq�D�ÁDNDd$���M&�:.Tnܷ���Ne�L&2�c��Ĥ���=�Otf�U[�X�9t~�n5��۲��$d����\��>�_�Ol|GQƝƎ@����>!l�A�gaj���j�V��r��&�V	�K�F�Ȓ�6�]l��4��zN��-�2�����ݛ������r��zQ�Oa�u8t����R��.�	���xaٶ��Ç:T$,B�+^��"b�,B�b�/*������>c����o�Ǯ��i�=|������ �Ѕ�!J,B/,B�B�K�P�+B���Z��Z��Щ
����ŉ��x<F�4xٳǍ���x�x�<�	ㅞ<x��{Щ�he6^B;(�V�O�e}�ås�ּH�ߟ�V���H��H"�V�Y�sn��Aj;�c)mم��k�d�+���y�z,��ua��u΅s'�W��D8��ѵE�m��g���?������p�y}�Ӻ�;���p$Z���������O.��·˧�wwL��gC��˻��fg��������33������9�o{���2�͜8�qU\c�cnvN��U��o4�n���N��<;Mo�b�^�V쯧νF��e�g�\�[⑗.���Q���fQr�[�6�&M&����D��y7(�i:&�&���W6ې�9b�*}=4xm��U]��1�xZWh�j��ŋ���h�a,�l�m����b]2��6Z֖���R�K95#	bRe�v����S�%z����׊.�Ӫ�c�馆��jγ=�mzb~�6�Xa�TD��0d,���2�aq��ЕPmD/k5r�$�!�1#��90[ʹ�V��A�i��
��"��<�j�o1�p
$a6�4�C�2DI�1r��&	�t+R�0n�.˲\����v�ZC�-3a4�N#�j��V�&1d���ٕ]M$&�%9JqwIƊ(��c7r�N'����*�����/����FϺt{h�[�˲J�㉕vYm������O��g�����*��v�1������f��;"�g�����\�өc��R�UO]��7s��P���{�BZ4�p�:��$�Hi:�3y$�#ʺ,hh�щ�_��9rŗm���\�"��>4DJ=�(����%��luc�nc���򪊒�<���!�`��!���5��7p+�4M4���կ����!t���.{�rY�#'���E"DD(�nZp(�By�i�n��^&=�$�5��6e��B?Y$%Z��[����+���g���N�a�8���c�Ī��m[7-�g��Q�����$�9Lgn�B$%)�d������)V����
l$x<3��G>h�wu����:n�]�I$EҎ�4��a.t�2�$�JK�tۻ	�6��6|4w�g��r�Q̤��<�a�>UWLq�c޷���D��#"��(��"�,�E�2�H�7itS�+s$�M�Ht;��USb=0VW�RK�m��wwv�K�]&�4Ѻ5��l=�!$!t�v����m6i6�_����0rBF�%�k<��k:ro�\�[N������N��*'QmR��`��Ue��2�u0np@�-6�l7� '�)�����cڥ�XΣggL0Ǌ����%�n�3fZ�0[P�4iO��8�v屴�p��ZwI�K��=6�4G�19C��8�֫E��0�E�-��f�U���a���A���Q�1)8�0���A�8B���K����f���3(�(�z��z�/�HΈ2q�����D��K��t��[3��f%P��+P�TV@�A"d�ƫ��%i���Q�QD5�g{GI��!!��x��ʫh���r���GS&��a:"&�C�5��M9��2Ք�Q����xy�Z�AF赚*bOh��-���K+�R4]&�UU
��M7N��):���=/�V� R�Ξ�	!$n�������>��a!O�HI$�HEUD������?�s����$����lX�!�  ��
D�G���_WK6u�R�1b����(��DR,���)!H�"�DR,�R*
E�*J�Q�������*H�(J����B�$(�%$��,IIY!E�QQ(�
(�*B�"��"(�#"%$QQT�E�X�E�J(�(J,H���X%E!EE�E�J)V�b0kXF��E��Qb�EZ,XeH�E��X��eQe�d��-(�(��(��kXF�(���-(�X��,�ʑ���&
�YE�-(�X��xګ����T�R��TQe(��[T�J(�E�,��(�X5H�Qh���,��,���YEYE�P��b���(��,Qe(YEb���YE�YE�,��*(��X��X��,��Qe(��X��,Qe(��(��YI,Qb�(�EJ,Qe(�E���(�E�E�,QR�(�as(�E(��(�E�QE�YI,QE(��(��YE�*RJQb�(�EJ,��Qb�)%EQE(��YE�,��$��(��(���YE�Z,RKE�X��,�����*T�b�FH1�`���	$%��TKYE�,��(��X��$�E�YE�*(�E�,��,RKX��,Qb�(�E�X���,��Qb��,��-!b��X�b�X��K,TJ*X�b���T�IEK*X��T�-K��)QKK)h�)d��JX���7�Z%���Qe,QJ%��YK)b�Qii%�X�R�)T�K�Q,R��)d��R�R�J�X�U,R�K���X��R�IjIb�K�K%,R�K�R��K�K%*R�J��X��%��)d�E,R�JR�XR��,R�,��J��X���Q--,R�QK�X��KE�R�R�R�)TK�R�,��K�K%,R��,R�J��Y)d��*�(�JX��Y(�J�U,R��K�R�,R��)d���I�X����R�,R�K�Q*�JQK�K%,R�,��D�J�--X�%,UT�V)j��UX�TR�K%X�%X�%X�U��VJ�UV*�V*�R**�Y*�UX�d���Ub��b��b��b�R,U��TUU��U��U��d�b���,"�a�D�Y	H�JE��"*K �*H�X�DP����T�H��`��	H�)I��"��,�a�a!H�JE��")!H�(H) ��"v&O�p=��1r��(L�� ���b (����HH��H'�+�������7�����I�������_�>���9������_�~��q�p}iF|�|�4$��>��ڙ��|O��^�	���f�%�������7S�������N�TO�_��ߏԇ��b��'�	�� �A��X"���D�VP?����?�\����}��!�)���%
R��'����?�_�c��'�����6TI�	�����_��$-e
���-��7���Y��&W���%%'�M������9ѷ&�}B}��~�6�\��\%�X��?��5���7�A �4�aP�TQ[W�
Z*��-����m�!-���pJ�6����4�W�G�����V�%��Z*��Г(��U	h���X�O�����="m�f~/�����G�8*S�����?������E�����-^ߟҐb��%'��������O�.�ڸ��i��D��k���M��
؏�G�}O�2�X�0�&���C���_'����?�����~�TO���8���Y��_��?Æ�?�͕�|G�.C�?TO���ެW럟?����X��a��6�� �H)F���P��p�;I!�6$�~wH�K=����d��>��&�1�n�a����Қ��&D���i�I�6�?��F��=G�����t>�O�1��}+��EU��&��2}�C�j�C�������s���[
w�Aj�h����'�?W�����R
9G�#������'R誨�"����T�+��r��*���0q�h����s�����?�>g�~
|nW�r�0~\}�v�,���m5$ļO���)�)����D�� ��]�0%���g�l`��ߨ0"�����}�_�[�5
O�>g�����/�>V�v��|i�xM�"����p���2t�'�M�|����T@���S� C�]S���܎S�6((�>cu����%.O�Y�(~��rO���~"�*�,�)��>�?����H�
����