BZh91AY&SY����O߀`q����� ����b-�               �                       �      � �    . ��Է_xy��R�Y�}� K �� jp5�f�mPP�   X� �� ���           �׾�$(H�R�QTQT	�!U$J�R�%JPR�"�H�R�
��* � ����Q�=Ɠ� R*J��E$�P]���N��k��C�\�w�oB�y������j�s[w�R��8�J������@�)�4  V����4� �v��|�t�R�����{���W���H� �|���`<�p/}�(��� ���U^ l<��`}��`�1{�     R�zy���l�E��T� ����)� w�0��z�K�p�>_]/������� y�|����@���1� �群��=�}|����  <�}J�����^G{� ���w)> >`}���;�p��s�^iz���l>��i��� |��� u��� � ����e�^�l�}���j�H�TU�͔I� 2>���`y���/G�� �����W�Qk`}�G��;����` ��_o��_ 3����x   E��}�5m \���ӽ� ��o
�y������c�}��z����n��ӥ}�����>ǽ��  ��v��s}���*4W
���U �(��� �Z ���v���`��IH���y} ��^���>gy�����R��6>l�� �s�饶���� >�v���=J^ c�a����`� �xUt���`/X����N{��   ����m��{n�I�Ģ�


����n��@/{���;���w��>w�CΔ�� ���)�`{/0 ���� .c�{�  Q���zg��J��}�=����"< $y 7�rhr�{��A�yR�!�(�{��z{`�� �    �     �A0�JSz����F��&A��)�)*��4� �h  "~�T�&�h      �ED�)J��0�42h�aCi�H��J FC�1#�T~�$�aCL�(h�444ad���������5�̀" �2�
6+b���ng����삠*���� "
�(�����A_�QP����#����?���?��������~ʟ� �
���U~t
�*�����B�H~J�/���?��O��'�Y��?��l0#�XA�LaGA��aP�@;ed\a� �(� �(��ȸ�0���)�)������*�����0���v���22.0�2xʘ�<`\`\e`e�̣������g��q��q�g�c8���>3���2c2x��c3�c1��8�7Lc0c=��c8�1���g1�g1��q�g�q�g�q���:g�q�g�3���c8�3��L���8�0c���Ì����&3�q�c�q�l`��0c8��c8��1��8�0c8�g�q�g�1��zq��=���1�c>8��8�3��1��8�1������3��7lc1�8��o`����1��1��8�c&1�����8��q�d�g�q�c�:`�q�g1�xq�`�g�g`�q��1�c�q�g�q��q�l`�:c�q�g�i�g��q�g�1�g�1�q�g�q�g�q��q�flc�q��q���d�q��1�1��c�g�q�cx��3�c3�2c8�3��633�c8��c��0c8Ɍc8���c1��3�3c�3��3��c�1��`�8��0c8ό�2c62c8�l��1��3��0c��8Ɍ=��8�t���3�c8�0c��c���:g�q�g�1�1�g�1�g��1���8�1��1���8��q�c�q�bq�c8�3�c����3�t�1��8�1��c8�1�c1�����q�`��q��c�l��1�c8�3��3��1���N<1�g�1�c�1�g1�c1�c�1�n��1���q�c���c�1��q�c�8�1�v�0c�1ۏ�c�q�c�x��q�1��&�1�c�q�c�q��xc1��3�c8�4��1���1��8�1��`���3���1�q��g�g�1�|x�<g<q��q�|x�`�1��1�`ƛ�1�g�1�c1��c=1�c�3����1���1��8�N<1�g�1�g�1�x�`�1�c�i��c�1�g�q�c��x�3�c�1���c�1�g�1�c�q���1�g��3�O1�c�cǏ`��q��q�c��1��1�1�c��Lc8�1���cc1�c�1�c8�n<q���1�g�1�iǎ3�c�3�c�61����c�1�cc8�7M�c�l��3���18��q�g�q�g��c�1�c�:q�c=����q�`�c�c�c=1���1��8��0c8�2��>0��)�*xʘ���������1�q�1�q�{`�A�Q�q�eCD�1�����#��#��#�!0c
c� �*c � �(� c ��2�2�2�l	����#���#����0c�(�*c*c �
c
c � �v�2�2L�� c� � �
c"c L00.0�2.2!��c ��c � �*��8¸�8�8�8�0&2�SSGSGCGGN0��8�8���>0�0�20�2=�8�8ʝ0.2�2�2�20�2���)���)���#�������\`eLaLeSSSS1�&��T����D���ʘ��ʘ�>2&2&0�22�2�0�"c"c*c �(� �"cc(q�`d\``OS<``0�0�2�0�2&0�200�dLeLedGG1�fT1�q�q�q�1�1�1�q�����#�#�#�
c
c
c*c*c"xɌ����T�T�A�A�D�e1�1�q�q�q�1�1�1�q�q�;leLd�CSSSY�SSSSSSS�La00�����������Ɍ����������c�"cvɌ����(c*c*c*c � �
c�ʘ�8ȸ�����ʝ00�28ʘʝ�.02&2�0�0/��+� 1�q�q�eP��@1�z`La	��΃�������Ϳݷ����	�#�$�y����ͥ�>�B���6n��&W�ռ���x+�m���j��]M�]�A��;;aܑe�eĊ�x��,�ǣF-h�4���t��N�����ۡ��^�V�oR0a�Gm���1=K8`�C
�PYi�l����Sw����%f��������� N;����\��Ń���}�����ةx�����.��%c���ܷ<��Ďsu��|���Ό?��,�:��Ҫ�Ј3]�d֝�q<�e����\YteAJjH�b�T�`��������]�p��N�{�[1��&7.���Z�l%����<Z9>Z4��ܩˣ������n�]����r�H%�4$�.�Vx��a�ѥ%�x{�ݤ�	vG�����鴻��������$ڲ���Y���9;F���peM��4��0����îoB�|�{��^3��2��3��vk��ݛw�R-�bM����w"c 75M]e@`�r|�[]�9=��bݲC��dN�5m�Qr[��/
d5�3����e�ӳo	�,�3
���f�T��tOm݂-�*��I�>���G�B�w]R��$ ^/��A�A�f�^�/�V̓���ˆoZ/od��k	+B�a��K��ǬݕEF�=Fs��Nu< ��&��6+l�L�����r0U��bPV��J\�,V]әg�a�u��#y�׌��jü�X5ܟ0'.�-wKm�\����OA�BL�a�L\J3h�@E��S�ι*goek�v\F��Ql4yǅ�b���;�۝�J�F�v	���K��r
�[�v\e����g<��ǉu3������5�獫�g��8P����y@�9wy�Fv��9��Ǫ-s���k�u.�f(gvk�-<f����e�A,j������۠��_��t��R'#K�w�b#c�g6�i;�Dݗ;X>��X�q���^6J�S�:Ձ�/=�T�����^Ld�R������W� �6H��RR寱p��D�(�.б�P�gi��X������n�9�s�[�Ý����x�I���gc�A{n�]\�NvWݠY��vrq`���)&�����8g#�ۼ���;��^���vu�r��	ͼ��2�>���kZ4l�Z���9��N����f�owH9"�8n�y0�=��7�R�=�y�n��U���l�w`�s�w����������p¨]ϕ0��p�ʂq�s�K��u��),on����$z�7��;7(�p�:�涻��9t�2q�X ��ⅱ�G�{���خ��/ ��k��-c�A�sA]��;�:h�Z�U�\�+e�Vr���P;c���bɋ��ݧf1WX�v��z�F۸�v��EYg9�s��A��:��N��+�oB&Ʋ]�����:҃؉<zO�����ۓ��d�r�6�Lx�n"��߬��N6��7��i��Ĭ�q�(��>%o>T��/��rל�<;�tV�w�3:��9b�������Ӑ�B�F $Ā�O%͞��Z{���)Ď������P���z���qǻwf�r���l�ǈb�.��i�ʡ��$�r��Y�ZI��'�q�����ƷR�k�{x0�������ɲ�8�Km�zj�:�p���G=�GX'20�������ٛY��9�JU����rU��,�@e4(�;�E�(�s�8彁��ZN�- 0��Dp�-�*P�k�	A�I�6R�^��M���_w(���/v�μ�$��ΰI��N��-Y����3��F)#�\b�ś���m�Y�v���y0����l���_(.\��]xhʖ��M��9�w'�]�V��9���]����8��;�퓵>��]�����I�b�Ꮯ>�-�����}qLT5�vq�'Ŏ�x��a.T�8�r���t:wy�w����&�b4`��`r,O�5U����ٕ�\I��$��0vv�ar`�	`�v�qv�ֳS�tƴ=�K"B/�ٜ�?^�U��A��@(68G��هy�G&#U�f�؂�&�,\L�g�-�W���C@7�$��Y��.-m��^�}����_>�;�[���a):������Sv�=�����Nof�㮚ٌ���m{�;�i�M���V�S�{�{٫����M/�e���ռ5l ȴd;���D9��E�(x0��)o�҇���gs��E��+=���իy]�{	n�k���V^]��i�8�]Y�m�Ǯ.<`�en�$�1�][�f��ӽ6�չ5���FLi�J�b9�f���PNܷx�a|�	�㵨�kI���ri���6jś1scLI�:.C�^��+
��O�W��ID���/[�q���x�]q���]�!�P2�Ks����m�
�ez����/�� �۽gr�s���f�u4��û�y�7���I7���]3����!I�C�.��+* �ݝ0u�*���pWN<,mQ^q%�7�)�{^o0��ܾL�b 7��V�WԼqn�xY�%��ç�Y��� �u�^�P��4<��9��;V+��Ϋ"��;{^�2�&mz,�xͥ`!�]���ex���P:�2گs܍�sX��j��}\Ǧx��t>�º�ۧa�`z�[�kdeS�w.Tr�X�,�9���sw��i���@�����r���u`Fq͏
sh4��p%lW{;kx���tnE�1ܺ1ɂ�����7&��Oc�^ �W,�g���(fE��b���1;i[,z;;j�گ	��B9�1�K�ʖ���r5�4�;�؃J˒V{�0�P�M"v�w���Cz<x��KS��Z��9�kR��t�@��nk��8����M�.ޜ3��N#�\ըj�
���Mym��*J_-#+r�s��|t,5sDC�nRgM��2͡�ޘ�f��o+SK����E��a�
���ɔ\�2�yGݜ�[z�i���=9'��o^�	�Õp��7�6�V6�z�֛�[3[�h}�X��=>P�����H��Z5���O52�Z���_>���<x7 ����r(�]܄��	�{F����d�œ&W0�Z��8���S��w���^�f������]i��z��\��nU�����e�݀�A��P� 6�޽�w)@f�+���a�i���H:��=齿9�r5r�U�T�zF���Agpk�1j�O(�~=�r�X�u�(�DrHm��'���;��塾C����8Χ�ow�[����k��wPD͐�i���N���R��ǂ�h���ׄ	�y��J��T�)4���ݭ���5bp1/%�xM��>��\�#g��NZ���u���� )��!�q�*�h=ܵ������\;�ݸ�=2�s�O�,fh8�)�r��;-3M�;�q�Y�w�U�6����y\,+���N������uf����
.�F�u �|��;�^���]�����xբ�f���O�wI��5��z٢��ec��K�6T[�t)��]0�w�w��8.�`�d�5qY���}�Gۚ#��*��;y�����c�Le�����E��;t�dC�%X^P��*Dv�]�l87rȦP��	S��5��kq��]�P�-��N�xYG�����6&���T���v���N�J>�����c�&L'6[5�N5�9���S��8𗺱��s�w�+z��]��9�ރak4<!��K�8]�gL;btgF�ޢ�<Vn�,�q�B\J�c.Re�8j�Ԑ�7�3�e�-��M�I �9k�Pkr�
���a��1��x[�+U�eqզi��3oi�\g��%���pN��#�Y�:����I�H����V=��9|Z�B�%ڵ�)���z�[��9�1h�����ܓ�ۆ-ɶ���g*�|��*(�DK{ ��NM�
��zʝ�;_m�X(s{w2�C�A�!x0G���Ӭ�*���/*Y�H�㋣͎�:(�f�<vM�w�C��λ��>A3r՗�q9J�x��I���,�((�fX�n��ȷ�ܾ�7}��x'2�kss�������a��o.���d��v�sen	��H�ՃFo��P3SM d��`�x��Z��nn�ey0ZH��2���=h��"�l(���8�\�'l�nށ�F�2WS��C8Tw��K���j�Zyۢ�bgb�v�bv�0A8��2}t����i�q�]S%*]}�X��h��-�t�`߹����w��'0�����^��7�uh�q �)�7S�Աs|S�8���g|���C���#�E6�!NO��t짔ŀQ�ʢCw9�[4�ǯ�1�b�!�n�x%Q{�b�x(�S'�s�W�5%u�x짋Vn�U�{�*�.�Oպ�d\�׸���<r����W���ex����Ш��-C$*�G�s�d Ʒ�
w�f��f���z��܆)�q	$��\��-�P� ��\Bz�@�0��ܰ�|��^�*��_�j��M�	0U��د�Ѡ��.��9	��ݪ�oix�
�"�ǎ�u��k�`0�(�+e'we���B����N��0pJ�sn�[����q=�ت�)dYrw;�Hټ�n�C�U�-�L�� |;��F2��1^���;hs��!�wh�$I�v۱v;yf�@�Cc�;_������0:�=%Wq�Wb�J��{�h�+A��-�زr!�:�N�:b)��j��o���j&e���\-nN1c�r�u�[�"���л�^�\tp��pG��ݵǼ�h9"�8�Z��
�R��\�no>B[R�6qy�:^Ӌ{��Q��1>[�t����uW��@zi�2�^:f̍<Bj�1Z2�.���49	�k)*���볬���N��P 7���.X8���z�wq�(�j�g#��jv�<}('�;1esK��7�s�>�����-YY:��}�R��6a������L�����S��ƶc����K�ʧ` k�2�s�XEo"d�<�w,��î����a��N �@7\���hJ�$7Txr��W�֧��TE�@��D��t#��WAV8�����!��$���f���O<J�>���Ŕ�����t8=硓l��ż��`{�����e�S�j���5w�qR0�F�A��Z�h��o��=S��𷫤�C�x8�Y�(,����W#�7��f���s��g�mq���� �����c܄��B;vX�Yw.�˒c�2�[��ɹ�i'�9w�.��ێ���ۢ���h������3�A���^4�0��x7
:a���m'�n���O������\/���f�^V �nW�%�f����s���q�Xk=��`GU��H�$]bF�A�@��RR�>�_��<��c���U� L�X� 	.aPu��&�3�n�M	��p�#F��ɣ-�SQ)qˊ���ϓ�J���.a���1{*^9�:�r��=gz��/�3&����;Fќ=����%?I2,�#'�sr%�b@���<�����-ӂoVI�ޯ������zV�&����ưa����CsuFt;��_U�_^Sgx/��yN�ĸ�OY�9���� �<rG�o+��~�c8n���hä{J�o-�|��xa����W$���.n���m�3wa���&�m��K�K L'�z	F�^�A�pL#F���4�a����I����YW���؊K/�!-��|m�є�]�R�?L�Rq��&OV#I�D�R�!��v�m�r�'�z�m��<��bg����s�d�:/���$���>~܋�s�:�n@���D�"a��pd��a����^&�2S ��Ԝ	A��=��LΘ��熦}�Q���f	�t��:-w��0g�������f�麱̈́��@x�2G_,�\�)�r�zs��sN��݇�ڐ���O�F�i�l��3���	[���
87��r�O�۹��~�v�� M�3�Yh��« E���z��f�BY��#	@��sE#0ώ�>Ӥ�$���M�2l���2��GZ�S���]�o��93Iؽy>�@�W�7����㲭�˖��@�]��|ϙ���D���R���^J�e��yݕ�c	����Z���v���,���$�9�2њ��E�˼��c99p������|*�8S���z���7�"�d���� Z�a\Ə��@͢�V|��
��4d��:�ތ�x�������Ni������r�2 �t�. �Q��L����ha��P4� 418r�z�0gg��Gv���9�42E��#��8����'H^Z�����5K�c:g9�(�H��<��rE��D>$2�#�Z�ہ�g}�(6��ZH�k�Y<�ب��{�N�V�ƹ�!�W�({�����&�n��\-9gs��a�zX�� ]{c�6�ޞ'Fe�G�yt��TNS$��� ӹ��7}^2Jj�n�3}�K4���	�n�D��A=�A�q�V�z���u't�����f��8U�,ᝰ�=48��@{�8M;!]��>��K"�O�=SЄFyuŽ�������8�4iKgI�{Gr/�;5L�Jǖ�ڸ�|��?D�00�i9�#����U>/�+�&�Nwa��N�:2��?tb�/z�L��'6.�x=+y�qXB�H;Y&H�������9]1Eˮ��������֠��.�W��1��=�'�xB����fj�q�Y��-��;Ї�&�g眲���r�L��5��6f��X?�"��[��n��u��{��y�G�! ���V���y �B��/$^H��)�S��$
H� �@y"� �!�B- �P((��^J!J��@��J��(�4�� � !B PP���	@� (�
- �д�*�"@ R�� Ay�/!h�U�IH��*Ј���% �� C�(�) y*-*(Ш4��"�"!H+I�@NJ-*R*�'������w��8;&�$�����u��wj6!9-��>�$kbmݩ�_�N>�d�`�<.ǻ�m��ٍ9�2�Pf�N��>���M�*�ED�+J	���Li�x��w{��qXA��c$m�I%��}=wۮ{����5�nƍK-�c66PFk;��ƭ�P�{�`���bc
����2�����l�ڷY�m�\��l�H�IZ��2p����h�bdV6˼�4�����E"��5AH�Wɲ�om]���5���E2D��@�V\��R�'F�qÒ�@
���j��՟���nm�{�o���!�e���go�t��e|��n�b�1nu���a/	��)!8�r��թ�N�'9���A�Z�27���f�!�!YR��^v񓺵u��k����S�g+CAڟd��+�'\���Qq��"�H��=������٧~'�x�<W��$A��BT��L�ո��H���*�|R��]}���{4��)�{�r4�����"_pwN��ֺD�r!�Pn�U�֟k�Z�Q�S��3GY�^�zu�N=�ʖ��y�F�k��H��پ6��0"���ϘmB�1c���q6�H�C�'�$At�uxT������mp�om�_�X�?Y�H�&�;�Ay�TN"����Z���P�-4�u���ٹ_�N��GJ��?y(w��k��W	���.��U<�������+�h�UT��?/0�Z�j$Q��pcQR4�O��y�|Aȟ���v!��:뒕s�������<�ޫYe`02�1" :�������A)�YƂK
-����G��q��TR*�"j8��[�z�{����8���X�	+Z��N[C:K��A��w��;J`����S
�����D8��9;�Ӻ��X��)�BnƍK-�c67���Z5�w�	�.i-�  P?2Fل�8�5Cw~�&��QQ���0��K8���o���;�d�XQ��1[S `,����ӭ��Ac,�e4�,�I�!�m���k�:��G���{���T���~���DO�����~��?�����W�~���ÿ4�/���/�%��E'w����_��è������u˼��NpH^�ۉA��(c���$$�����ޝ ��ECv�K�K����y���ڱ.�%��>ڷ>��M�ܮt�~>�b#��`;�L�ޫ�f��ׯz^&�����5�Sf9X��}:m�g���=�+b�ܴ�~+p�N����Ž�0�vwxT93�=�*Ǉ<��~�ǜ�瓼r����tN7����-�8��8b�Oz#������6`��x�@8�p��d��\;�Gײl�{D�]��9vt���S�3y[R����q.ͨu9,Ԩ!�?P�~s�^8m:�ɻ�h�<w��=&��#f�����7�acޙޭv�gp���Y��aO�9�I�a��83�k�j�xya�k��q���M��E����ݷ[���V����M��;�b:2���#*_�{�����/-[�;�R5���FhG�.Y��>XK�T�2q�+�L�v�s��z�+�}+��K��p�:n��>�ow7�}��k�z,�{�_M�7���T`��b
Ħ����iimho������뮺믎���^:뮺�뮺�㮺��]~�_�?_��~�]u�]~�:뮺�:믏�n�>8�뮺믎��n�뮽�뮺�뮼u�]u�]~�=�뮺뮺�뮺뮺�u׎�뮺뎺�Ӯ�:뮿u㮺뮾:뮽�뮺�뮺�㮺�Ӯ�뮸뭌��."=6�<��UD�x��[��M�}����쪷\G;9���>�R�hy��[@+�_z�ttN�׭`�����m��ƾ1�1�U}���~Je��7Æ�e���À�����.�߲.mT��|Ȉy �����gW�{�����ݞ[��؂�x<�=ݚ��u�ԗg/*��=6ww��QO�7��w��n���jK�w�3��5&z�갾T����j+�h����;����>WL�s�/z�s��0{����t�8�V���1i毻�0������y^R��7�Bǀx4(�o�cT�2[�æ��Om���f�L�{S�k��=��`�G�ϰY�mY�/.�ӦO\�^�}MA�����r@��+����y�śl�l�x\��'�]���fƐ��g�������mJKUQ��:���ćB�s��g5@��d��F�q��*@��E��������ݱ齪�։�����@��3��3=D�y��h���%o|p���{������"����!�!�|^f\VM
3.���y{�W�6DrE��D�*�k@�(�0DІ�*.��ه��SV!f��2��&#�Ȍ���5�47�|u�]{u�u�]u�]u�u�]u�u���]u��_�������~�^�u�]|u�u�]u�_��������뮺뮸뮽:뮺�㮺�ۮ��Ӯ�뮸뮼u�]u�_�����]u�]u�κ뮺뮿]g]fu�]u��:뮺뮿u㮺뮾:뮽�뮺�뮺�㮺�Ӯ�뮿>@��>����u�D�zj�������]��g��D�y!�������揑Y�gW��̨����p�A�Q~���b/&���9��аdfx�T�g3��u��}/6�wֳ1v4����y\�#���eV�G��/Q�� ����<i��tKQ���)}�<��d;6.�!��v+{�zv��E�1qxiYˑ&������@}��m�Xp�F���g�����z*ni���Ac��!dzU����� ,��Y�y�d��|IG מ\1�3�Ϝk� y[��bK}�oz�����}���pJ]'ʻ��U|M~ ��Y>�T=�˜p	���0Rr�r�"KF^zdf}�ƲCfW7_7@����c�v���pJ�����X��'�׋Ώ9��{̳y��藴�}�c�X�j�|����⨭m��O���纶�^W�'���?H<r�j�CaP���M�O:׍&A�b�%�׷�E1�ᝏ|��8/��T{��}f!�|������ �e]�Ք�[�G`�{�{Ǖ���y��x��.����U��x�̡m�}=�S|uz��P���w�;�[h&�WS���,c�>�؝�D�7�f��� ϝ{ܝ=�'R��p�:=�31�yy�fD;��q`~�]�o=��ٙ��Y���4�Ly�^�~{��n�ؽ�7}�}�>�2b��R:m�>��fb&��R�"���q3��W����~��C;3��/	yV�U���f�m��gu';�X�Y��)��u!�����>�e��ܸ�v��
�'��	���z� ���lklllo6��u�]zu�]u�u�]u�_����]u�_���������~�����^�u׎�뮺�����Ƿ�G]u�]u�_����뮺㮺�뮺믎��n��N�뮺㮳��뮺����]u�]u��G]fu�]u�G]u�]u�_����뮺���^:뮺�:�N�뮺������`
0���� �iT�������7��0hψ�����K����ov�F�`���<������q�s�=�Y��r�}�zA}��� 0m�.��BC��n}��xRe��,Drz���t��d�}��>�q�|���Q97s��u#D��O���?������ڎߠ���\{��{����x�_x��v��糖����3w�O��}ݗ�}�����M�;�ֽv ����4�0]�C��ܸ�������sڷ��޾�b���tiy�e�TNf Q�䝶k�u�Ú������]%G�!ן$*=�U�{�~=Ə!�/�PE]���.g{V�{�N�OS�U�x��!��vh�������n����No_id���gK�k�h��Mw>\�d�<�����	�$��C�OX�3��T�s��﷊��^�w'�>����ӛ�ϳq<��"a�G^���s}�Z�vfg���
��afs��׮{I�n TCadM]��%N�|.ޘ@�10�m��i�����l�΢C���=]�L>��\|����#���� ����U���}�<��٭Ê7z������vbK7�M����:ߙ�v����BI#�2��id�ǭ���y����������]u�^�u�]|tu�]u�]u��:뮺���������~�]u�]u��]q׷]{u�]~>>>>=�:�:뮺뮿]u�]u�]~�κ뮺뎺�Ӯ��n�뮾:뮽:뮺뎺κ뮺��]fzu�]u�u�u�]u�_���뮺뮿]g]u�]u�㮼u�]u��:���3�A�d���/�/Ʋ�}��)��FouK�x���o���ڌ,���ɪn��+���&�%�~�9�~�G�P�э�==�2�!G̈����}��;9d\k0��8{���uX-�=ݙ82��S}�>����x*��d#M����ǚ��@��u���kدI�N�w����B,^�� 4y�=��c+��j���]��}Ey����рy�hA-.A�F-��Ӊ��<_l#7o7��t<�vD�N�c�L#�z`��墊g#�Bΰ�{5�;���d�6��)�����G�vU���[V���w��Ì0�w�vp�~��x��iL��;!��l�z�xb��t��O��x8W�e�
>��˪�i�d9���M�����w�/���fy�����	��1Ƴ���r�B�<Zw|R}��Ww?��'�p$Fqf`|��{�g���>O7o�N����nul�a�_`�ڙ >ۜ��7Go��[~�J�k����Q��|�܅��L�}흗GbGݾ�ؼ�LYī�w�=*�2��Iݯ��_�^��>�7˻ϝ<u׎�:�u�_����뮾:뮽��u�]u�㣮�뮿_���?_�����]~:��]u�^�u�]{u�������]u�:뮺�tu�]u�]u�G]u�]u�㮼u�]u�\u�^�u�]{u�]u��]u��]u�\u�g^�u�]|u�]zu�]u�u�u�]u�_���뮺뮺�뮺�u����}��x;4�ޓ�&v?UWD��|�o�7{�'tt�͘�� �7^��<~>Z��zB�����B|�.1��:��K9u�����΃;:{��g��X�3��xN�&<2�p=�:ZLY��>��U����Sd�r�N�ơVƖS"���x��Ɠ��⳼���,�+��դy�o'��;���Sy��q�۾�TJy�U�:�^S�ɯǒ)f�a�����^[�H���z\O����.�;}�9�9,�øi�I�qϼ\-o>r�ݤ�=��A���JE�Q/s�����_L$��Xp�v��������ޓ���r4�,�j6����5����H�wײ��MY6v^~c&��'-�'�K��7����1�0^xE�2��`���ldL��{W9�����i���c� �\��My�{��qc�_{ʁ���bEҤs6vz��0k�L^F��#�X7ܽ�R�gy^ �W����w��8�_���b�)n�r�����t/i`a�}�n��|��gw>��ѹ�:_%ݗWvyvn�C\�=�{��W���]��/z��<�8�d�"^D��eT�Au ���u#1��������������;u�]u�uק]uק]u�]q�Y�]u����������뮺�u�u�]u��]u�������u�]{u�]u��]x�뮺��G]u�]u�]tu�]u�]~:��]u�]|u�]{u�]u��]u׷]fu��]u׷]u�^�u�]|u�^:뮺��]g]u�]u�룮��6665�5������[����ⅅ��U��l�_*_{��+���6s���϶;�5`N�ߜ�|��TqJ�~Y%U5�\���oK��Qw-K�|�|}3����W(�rN���z0�븍�ϯ�H��2{3���Ƌ���:�{K�弄�8,�8�[��=�X�P����x��[˔z�{�zm�ۗ5_ ����.n�xڼs�{۞�j�F F�}O��{$]c�O
�N�{پ�{�A������TT4�L@����}u��O���<<wl>}�j��H^|��w[���:{��l|�^��Ș�=���U����s=�f=�wK�N���\f˺����f��]f�s��{[��ӷ;��:��4�\�?.�ޜ(۸�G���g$��ٻ�gLG�k9��uV'=��b���u����]�ړ�1��|u��_���#g����u;��׫p��y�<d�t劎��À��i��f�ʵ�a�'��D��{��h�~xW��=C+t朶/p.]�=sE�tC��x�2�H��?n���%����
jX���o�c�35����ˑ'{rԓ>Hr��D�����'�����Vz�B�Lo(�yv�k��?���b�k�h�g�{��}ٳ^�����L�V�����-��U�v�w��X=f�33z6Fs\���q~��;�u��� ��x{��S��:�4����q_3��hS��?/,��t����wN��u���!�<B�>�3�Vs;���dG/?Qa���
7�صr|'t>o�o��.���Ixr�	����� ���q=�߰m�R�bd$1�!�M�|8j�pr�q�oS��N�5p���I��Lӽ�o��>�4������i�9xVi�@j��8�b~����T�}�xw��pj����j���x�NC;�oLr�Ǝjj+J�!2��	�b�����O^��&Ӿ�ؽ��2�g��=x{�[��w7�I�I����r�������^W�z:'�g�愈�p��G'7�^���Ë��wj�^w��f\^�^�����hS8_���{7_K��ϳ��M=>�ػ��8⯅Yvh���q�?G'|kns�
�94�.��J�k�+�Oǅ�e���V��3.d����A���+���r��w��Q�=w(�cbxM�7�r�@�Xzz�ET|6�3ϙ��ʀx՜< ���x+�c;�����+�w�*`�>Ӹx�ǋ$�׽<{ck���|���F��:��{�%�h�-�\�lw��������ػ�tN�=	���}��hΑ!$��7�u��(]�P*|i��>���a9��%�wI�'Z�7� �d�-^�M��v�H��{4.�<�oA�3i);콺#���.u�[�b~�/^䃧w=����T��-��z	���6`����f���f{�Xу�����M�k��zB�Mj�F��
qw�㳷9�}=8A��ܝW-��o��տOw��V�_��<Y�>��6)�>��>��Oz�Π_vj+�n:��\�a��|7����L e�w����� �S�/C���'_hX3ی��S�Т�N{p�Jh�����hҷ}��យ�>��ܷ��W���{���K�Eמ�:�}ye~�p�|�w}����绬n����G�ѣ.�7̲�\��>>�h��'&��nC�h��.wyoz_�W��q�^�=�����r�H"V��a�����!E?F|Nz���RҸy��y����� ����bVF9�Uw�����{{�:yL���CLn f�vfk������ӛ��ڸ����};=�W|_����p|3�)����=[2�w���L��6�K��lܝ�9��S�2Vwh��_W���"�:�z"_5blJ+X->S�����ٯ)`Μ���l�=���w�*�tq�A��"�,ϳ�_,��=�/�{��pY}����l��9v�f���o�a�?�Ok~��������Y�U�rzo�v�S(R��=�;��{�n>�'��x��.���G�!$��f飀���<��z.[406���j����[qň<al�����jлqn��쯫����\^+��d�m�x�zfH�|<���i^ok�s�x�%6^���{�����T��W9����w��=tٻ��W^��v�5u�u�f�=����[o]	��{��}�x�x�`��{��2�}���= 5�k��5�"��f���<�*����v�}U��e6��;��Oo��q���E�*Ӽ��Q�q2Eשg�~����f�fo��o_����v�����A�W���N^+���?�w�θ�=����:�sw����TkpYE�(��x��͑l�O^��t2�V7�\c6E�X��;2������ɪ)� 8���u�6&����׫V�뎴	"�YD���9Uǉ�\>�Ӝ0c$�☡��C�ZQ6�5�W�kS�յ�)�0B����sui3j�s`�MOn˻v՛�]<�B-Vk`1����˝�i�21���q�i���k����:n"��ͧ:��WDIE�;y�hm�!��ÝV���,�����3�]��=y���nͫV3��t�:����5��%�2ې�Y`3n� i7\+\=r��-Z��wl�g��;:'�.Q\疱�uHevz�v��-�Gn���r1�	�ma��M�oZ�0���v"\��t[`���t�]�onۃs��69a�LQZ���d�u�J�f�g��眼�/*n��Mδ�����A��Nb�YI���4�fC�@���R��E�VY�vM�iF�����V��;K/;��`7���Ek֠K����V�5	n;/.���g�lf�6v�bX�����F&$,�c.�Ui�kKfi��1$8K4�1����ݬ�6���968��
W�^�y��ŘF��m��䥱ֹ��=mq��e��/&�S�{^�Ɋ��U�$U݌Ƴ$إ������H��oi7l�N/==o��c��^�Ly{t�"G�킵H�XCb#�.¼�7FR��2�.�i�ff�
KX���0Ř�U�խ�`A#q���x�t�-`D�lX����Zh8���w�uѮ�;8:{v�N]d-�8��]f;jW����ɻ>�s��9xxqA7]���N5m���u����If�NU3A�b���^��Bg�ƇAg��cts�P��]m&rK:j7c ��J��t������X|u��!��;���*�������P�]f댜�u$��lX��X��\7Gp�ĸ��l�!%�79.j\�ޜ۸킅��]ID$iR���Mrbg�ѝ��;6�j7���t�[ �Yv�nE��U\m>v�Wg����&��ٳF���	;�.[\]�m�F�P�/���nb����lh�X�Y����I��2�u��Nɺ��ZGi�r�WF�RbG�1�\��ݻ*mpˎՎ�k3��-�M��Fm,��3�Y����]��#؎q���9�X�%�.@e�1�cu�©��/Qm��<���O��!θ�v�6�rP��wf7l�����Bg��3��5$�	����9��x�2lɌ<*ݧ�=�p��=gv�5��f�nNVP�c00ڦ̀�j����E�]rӗ�]e!���F�s=
�MȀ{b�u��ֵ�r�Xyv�fxܸ�=��=U�[��닷�ǋ�f��.���rk��d��ɍ]���gy-<��uBlp����=���ne7:*��`	l��A��:�X6G��]�����u�9�۞W]��� k���,�[]��ێ�#�'�Ld�X���nnݽ�Ξ�q��&p��lűɱtF,ζ�uXT��`��!GG��g���7�V-���H��0]Q1��݄�0��s9�a���
w%�,s�3ڂ#�n�jy�[]&N�wb,v��07�]6��-��GΧ�����w.�`�l]��L�z��k������c����m��r���(�료�gM�lY���e�絻k��Ρ���t��]	�*tf"Y���P�phl��\�he�'� ��;ێFd-��VQ�<�ܻ�Ъm�U�+e�CSK��И��3���X��j��3t�T����o����T����\M�;1�s�ܡ�[�::|�Z��z7i��9�g�Wk�X�5�¢K6�K�%�9��^%��s����;���eXҔD��g��1�vS27O[Q�5�x��ۻn���F'����B�!�lB0�v�B����D�N�WB/9��n3;:�z�0������b�]F��d�X��a���Ќ,��2�tpv�F72v��V�i��c[u�X�H����M�]\�Ws�k�+.(1"�dj���q\�����d��&^���_L<��9�&�"��f�)�6��l�R�W!�u�Ğ�iq�cc�Z�ն������t3"�WOl�[�[�=��:��ҌlX̙�i`�)��k��eb��GM�6+��L����+gH��e4s��Isf��.Ѩ��
�A΂!Vd]���x-���nX[rnS���ågs�Tv��:[V�;Ek1��K3H��sy�7@��\/(�k�{�I�3�o_<��n��B͑�lXք�m�4H�ϫGYa�۴t!{<��p��C�����Mk[��.��u��6��f�Y�F���<m�km�]�Ś99ᡵ�d�\����@uku�X���X;l�W�+Xs�� ��;�_i��Ѻ�A�����.h��խ�����uM��hdus��J�T�:��cړZ�2S��sI#�Fl�`�KW6���;Ny��q����8;F.�Hk�\hB��
9�^mu;s����ȓм�kZ��.:�-���\&��:����O��;�>��.�V�K׉�V�ZhM,���V2�)
-˙c�vXL��jVk3h9���B:X�Q�4�<�ݸ+nw6L��I��CT����f��jǄhy�;�ֺz�r�)��5��t��"�n�)� ����Ζ�xY��1�s�x6퍜fɆ��Ŧ��zi�X\�-��Qk+/Wl��Ė��b�m3Y)�y���:����E�s�=�h�Yx]ۓ*��q�cOvg�̧s��^;WC-q��{p9p��/h4��eխ�-�i���V!�h�.]�u�vT���M�uE�^�:MW�F��1R)]3c��1�I�+�m���1���Y���Bi[2k,�ZɫGT�PvƎ�x5w&_Վ�{c۶:�g����:��'5-��IZ�ع��ѓ9���ƌz�6���r���s[S��yA:�%���&�j�SJqv쎺��L�۰r��e.nz��y�lj�]+sNK��ی��Y۠T�`U��N�6�gL�=��uǟd��P]�;T+�"g�����C���l��jh��$Щs�m���U�;�M��k�R�>,�G��]��ڋ�rQ���[{�R�z����3��SLX]s��On�C�SJx���簮KA���<��ִs��u��nMT`�6�u��,-e4�L�vz��!.),q�]gY��1�Y��U�V���1s��<\]�r�uw�j��w.�m3lW:|�Ц9�6;;�Qs���.8�a���ԝ�T��[�1-aK��"�dI��n86B�i։Mrq.��;NmM»5�����Y�w ��v�I��7nR2�y�;8�g[�ۆ��0�9��j���'�۬�X����DN6]1l�:��#XX�4�^],݅B"�]t*����u��˭���,ʶ�շO�De��D�lkleQ��ꀳ�˸z9sѮ3���-�kc��aϢ�ϝ��L�x�V;����9#�	PZ��CW^��b���h���1�<�r���iø�7n+��sxG�;EO1q�	�R���1'%��l�m�2��^�G�l#G��K;tg$��Ѭa�f��,�n&�0dR���:�;�����ӬN�wh<݇ї<���h:�F3t'�t������[���p��=9z��ݝ2-���:�D����=<GF����n@��Ϩ����Y��j�`�uu�ke�m���4޵�V,=8�k��[�:ŗ�4�Tlmnnl�,t�����q�#���=t7ny���x^��i�I�z�sZ��&f��X\v�8"��j��;���f��g�'��%=b�%�:. �^��>n��q-�yW����;��/a�X�E1��䂊�ǞH�?M����6�Ef4�jى�gP�-/�R�V?�co˓[��Vt<���_[��"�KQ$��mS����,;��b|A�T�ǥ�n�o��M+���\2´�~��֎�?H�4���;tdM��ȫ�
���Z�m.Oԉ1�x�OT!%X[�n��(H�	�u�8<�q0�Hzځ�Ll`�~,�y��5���;���n\�r��Ԙ��֠r��3U���D鑑_�@�HJq#�	��'��;���I�����:�����n ��A���`�}}fx?�����Ƿ������:��j#��y/S�@
+���P�*Ns��R-P(W]rˀ��4�"��^�8$��'ww��%������ܔ�Qԇθ(u<��PN!����VB��K3;�D��9ؓ�G�wx3�x$�@���t�V)�"O�IЋ)�*��15I�uE���eϳ�0���?u��������<�8p��Y!{�ӘR���ye���8��W��ۦ��0���ҐX�A���OŁ$Ȉx^�L��/�@溺ݫ2�n�wo��D$4�v�*i���o�=�s�0Ƴs�g3��>�˗.\�]A���o0�QS(���5�'2'��0rD�O�'˂:%�^�ٲL�NHbvJ�1�,�=ϰ�w�s�y�gٹr�˝Kt�\�JrHz�D�<��I�/pD�C��%��͓�MX	 Fg�1Q����#���+���u����?�=�s��7.\�R�-Z�chg\��-+<<�$����B2�)<R�#Y�XF�ks�{q0#0+�'�0��
R���^X�"+*C�����3��.�Ç�l��Lrs9<,�hVI�8*��3�8"ĉ��Vb!$����$��s-cD砘���'H�t��#�qց�$<��;Y�|˗x�I��3�Bs�����xI�ӈh�I,���m���(�G���a����{���ݞ:�����n���t&��2�ħ;��,0\��n��7=�)�㋜qYv�,���s��{g�\z0���4$5�
W5nJ�g.�	�K�q,�eY]�c�;n3u�(�&�s1?�yt�>X�Fm�C��.B�kVܞ�k���ҳ�ͺj�f"��c3`g���mET�e�4ښk+RVn�]c���9����[�Jn�:��tw<	�\嗜�e��{g��Ѡ*F�%�%�n�UF�b<j�;v3�e�1�p��(5��rK���F\�\����U�Ik����.�$:�Cvo!u�n�s��1�j���\�M������]p���M.��7E9��hQ�Nn�/P� �����c����Yj�R��b�"������[Yvi-Ve1�Y���nK�nxl���'v��]q�n5�)�Z��SA�0��\jëͣBť�S���X�U�QC���Gv�鱣��`�&�V^Ex�=�8v�U�Ǟ^��{k=��O�Lfsk]��n�0"-'����#�K)�g�xq�h��o��1�T ]�aD������M����	��r_���V�9�&��i������L\6��@:x�н;���ˁ�h�˹5!	��f�,U�u�e�iݹ���N��yƎ.L�7]�wcҒ� �J��K��e��2֊eK	����e5�㶺�2�n��<��	v�BsW�Ս̦GQ���S��t,�-����!*T�e���ƭݨ�H�"����;��g ��a��������%�F��y�m,h���%�l�lI��j��P�Z�Z��ZIU�⤴a-�2�R��	e���H��YX1DVQDe9	U�[Օ�إ�KZ$mzX%��z�,,����ZK�ևT,����׭���B���U��X{��)����o��{�t�{��H��	ú����\����i��K�"�{�B�eh�s����ڧP�7�Q5���rIkKL��(5l(�[��u��s��n���a Ӓ��ǀ�u�E�}1�>g^7��` �m{��Ū��N�d8�F��1�̦m`!�!����t�� M��T����Nn�Z�M�Ԃ�ǢT<K(q3�tAP(դм�
�x9�{��WV�o%��ϟ��|S>�JW���Ybh�=��|?�,�"H�M�1'mL7r�՗��4`�\�P'x$���S�5��V��q �P<�����}ie�x�vi,R�C^�K��|��]�*�z�M��ɝȼ�p�NE'�X�Zq�G�?ߛ������Kg,/.��%>�=��.#z��=�VJ|ɯd�X�jK� 6�Ć ��Z����p�u� TNd8�;S.��<�+�Z8�����Vx�+���l������8�2E7�泈� ���rS��B{��:�'�Uݱ|ovB�E R�&�5��%�d���toZ�p����O��w�(4�Ae��L2@k/c����>�Tlh��AW�FA�MO�.�y��x$��������}v$��Ky��O4t��N�]�ݞ۴���d�\���8��bvԝW��@���0��``��c����ۯ�㴰0�-&�Yx�jkĻ�
���k����0�����\�	��m�;�!2���8b�\ϧ~zDy*�;Q=/�m�Dd�[��f��Lz^�lԌ����|�X��r�:����gj��Z<p\�N�>9���槊3���"���޹g|}�;�0�u�y	!� ɖ>V��'K�h7b-D�{w��x1ܽ�>1Z���A��h����,3*�A��צ4	�����|���c�o�3iǝz��h�XP|��F
=�1��S�3�X�K59�A��H���%G�~��M��{^�t؂
��ucd�p*����5�av{P�$�u���v�&�Msۤ�Eb���W�'-��g>Z���ܹ��p�)����&a�_eCF���ظ�h9���L,���rf�]xF�����>5�!��%n��2CVjf�qs���|My,uw&K�Nx9C�Q>x��֘I�~����u��@QZ��d7na1D���붏Sz�N��AD��m%OPDg�HL�/y�X��"�>ڧiIm[)�Q�����AH#��b�����@�8۝J�����œ��]�ӊmT���NfU^	9hc�[�����,/�h�
	ֿD2,Q �LF���i0���D����J�O�#���I��o��=����ɯIP$���HI��L�ź���O{����¤� �E�����\����ݞ�ۡ��M��x����o\�����~�|�Kq�e��/�x}��#-�Π���U굒F#�����)4�˫�S�����r����|����w՞O�L�#Hx޿=t���]Bsq�0��}�<�C<4�l(d��._`Lc�::fP�d-�u'���@�+;���Rbo�iT�o<��1�WR���ϡ��|�!�+vY�#Y�y ����Qƽ��Y�8��W��r����ê�J;Q�o�����n���z�ߝ G�vX�-P>��{�Va�N�L��C)S=^,ɜ���m�9�eпgoBg�>{=�/75��� �{�W��l�rO`d�0��31�&��JD�ݕogk�1q����kU�.o^� ��KD��⁛ g/M����4�~��!�P�]��&�k[t.v��V$�ٳ��d�)JƄf�v�p��ֺ]�A�7��x\�f/�~��x�g��e�y��;���d�GZ{d��6v��5zd����s��{K�vm�N���9{�'<�.��w:��J��M�hAv�f6�`s��wY���"�Yx�m�&�z�'���
Y���<�
A� ܬ�[��y������?��Gc���/.A�옢�y.Lh��לe웡qj׽uz���.�F�� m��L<.��B)Ey�������}N|֛}��N��kQȘZ�g����Ң�W�z�E*D������!c�p��6h3p��Ig^͖��@��w���\k����.	/�������uB4(dP(?���fܡJ�Ӥ�wN��2CY-Ȉ0�)iͷx	Ǭb ��L}��[��F��ex�[�F��ƭˬ�M�bA��v-7~��!�>�`{s�o��M�$LC��l�V�'^�u��tU�+����Kk�W :��|^�m(�D�w�C���J����2�߰rog�T-��>�{&Ô
�jeTq�c�o���!�U���AH/�߶/�/�Ot�[c����$��q���Q�^1j��Wt;��W�]2���,BY���&�s�}��=��༙�}�)=��)�b��È2Dj�^T�G8��nu��͜}�W��Y���tA=dF1v9��,�)�s�As�!�,�x;{y"�z؂H.�޸�@�c���X��0HL|؉ڷ���W(/���t�?
\܊w���^�o�U���N�0L�{2)0^��v�GIG0�y�뱛�UӫP��j�+I�y+��U����{���*v*Tō��]���	i[�����h��5H��Y�^~�2��,[w���=�S�uS��.��z�D�m6�<���m��2)�ļ�����q��6Deı`��m󾵨d���7����D�	$U�B&!���[l=j&�,9��2�򲪶�W�>	 h��E0�*�w'g{rx�2��?k�=�ܷV�y>y?~l�(�\f0�JPb�!��o%�i�-.H"
mY�I� �cs0X&Awpd>62��Q��������S)�<��B�>���2^c�ܺ���*� �ݚ
0�	�=�iA$c�lǣ�	yhq9V����Ǔ�6c� N��y��p�����|�]n��cv�T��ˍ�&T�p"tl�vJ�$e<�HƣVy���A|�ƚ�g���R�R|S7�i@,��Ǫu��k��Z�_������֣c'�Nu�Aj=	��L��2�u^�5D��lu}o�#{��}���\��~��%�����Խ�	����5�5)Uﶓ���p���������v��������/~qK�kqY�A �s}� O� pƩ�J�U�dLB���>:伝q��5��~�Ng~�c��Z����(�3��a�Zg�4������,�Ę��{�&HN
�9��. ,0��h�w�>��ߌ������f�iJ׈�I�pY-��F-�l�XՈ]߷�-߼"<�"	-JƁ�rJ�k#�������kb��m�h�n#+�l��FĖ��=��=ݖD�>�۱��f��J�!a���(ڝq{:��b|�	:�_�ݵG���|�ƞ��'��UW��}�����J
�ja �isU~(�7v�M<�A�N�@z��l���C��X�F{�k|��s�nT%�����ɨ�~�%�U�<�먼��wɜ:���=�D&�N
eo�L�I �5����A�ɓ&����U�^��P��J�1���[qo,	��i��{vh���F�s�����#((s�F�׼�%�D��������~QM���S���'���I� �3gWݍ%�ڗ��UU<}�;�%���ƴ�|��b� x�
#Z\�@��Z��	��H�[�FF>2{45�g�8�)LpŦr�L�|��x��M,3����|��Y>��)��;L�˭�:�v�l�b�,��s
���U6ĮY�x�g�S�lv��ug=Z�;hx�I:a�Nܛ:N)�9`<<�%�7��ٸ�s�BQ��4Ð� 4�ۑ�+0n�6�[���ɗlq���9����s�((i���f�sw9�b��l�n����)ۛS����ڻsٚmw7i�v%ҭ�tB2������֬ 5�T`�i��^�������2�;��o�cX������M���"k|'�(�g/�oϼ�%1�Ф�.��wc搷ϥިP��A�KϢ��;�5�&{��ǌB�ʄ"M��uꭥ2N2��޳��@ �a�ɐ[ȷ��H��>q\wߧ�8(}K@Kէ6C��T���	0�n���y����EL�c�[u������\��չ~�-���W1������ H7�	Y |�Ɖ$�;A�N�g�lY�A�N�W��출)6�>nC�����ہe��&�q��߽�$e���y�A{�ܹ"��E1�ב�L'��TD-�g�L�/�p )�.��8��
�ه�n|���~���k��c�����ų^�\r�:��r��3�D=�G�g��Ǝ����f�(\^B�7�u�d^y�aIɠ�[>����=�eK݁ �-I�\m���MaA�vq$LD;�=lv�ኲIN}�L� �q$����[/sm፳�K6��IL���XP�!m���c�;��9���o��	$7��3Lxe,sO������'Cm�;�t4��`��c���ڸ[��
���6���LH/t�2|e[�Q ����>��;��o�>	"�7j
�S",��� ���Mt�@��eF$SAfBSi��6ٙJ�=����eTv����@�7�l��Zc^}>�n{k�C�� ����L�B}���� l�3�0�*��^��Ǳ;��l���3����z����Dp�{Ҹ��G�N�<�*g�7�,$��9rd?�Լ1%5[�A`�a�'5��wO����]�y.6���I��w�w:o�y7���JW��Q��^Y^L?vw�/w1��%�e����_�5;�v�b�Z9��f����^=>�5��=I�����{��q��
w_N�3�T�oNܸ�kE�ky8Z�wE�]�;�|�B�����0v�;�Ǭ���<�����>��5��;|���n��㳞�|hS��+gQ������z���2�Gb���;�Oo��{�c�����&�=�Q�9���!����L����3����u8¯���������^w�z;�Ȩ�%�q�w&�~N<��+oj�ҩW幫7����{�=���̝z;S��[:�}�`�X1p>��a{�{���0<t�s�f�%��5x!���tc�x��%�MLm��ݪ��}�b@fL#��x���t�$��S�g]C� 3|�y�o����[�y��L�>O��-�,YUy�����;�%�^�x��o='��՚��t�5��wQ����:���iɝu����^3ػ/1V5�3����+LѾל\��2��;������v�����13��J�+ް�^�2�Ŗ���Z�3T�!���t���|�l/8k!��|���^a�'�k�j�1=�-���H�>��G�}|s� ��ڸ�0�U�.����#��*��^k�B��?��{^��F00�??��8wq`�� O��Y����_�D��ȼ��"���$�$d3�P}Ό������Ѕx'y�Y<�G09�������韏���믯��ooo����E`JO�P��s�䒑�# �-g
��o0���9u`�{u��==3������nn\�rT�$-c�������wq �Lu�}�0��M�s�
+�Tu'#��Y�y1��gq��}���.\r�q�&��|;B�0���U^�y$�3��2�8"ID��i�{���>�3?~�~���������ws˅��Bd�RDNv����f0}ǣ �Ax��"<D�;�~�ǌ��g~<u���Ƿ�����G.s��G�����	ˉHJ*�h�U����I4��ﳾ��|秏����N��������ܔPy�%$D	���S�Di$V0��AyA�����9�ws�,9>يH�(q���lD+8;�JLZq8��N����"�%#���l ��@���`�$b�c$��X��%�p�c&�'�U!��� x0N�u�8�1��	1x|��D��Xa��3�0�_7���!�]I�'M�-��;	J��=]K����c�i�1? �����j[��#�f�P����"fE^�f�[ 伌�����d(펥�NC��GK �q@�r�"ˣ�2��-��fgz�:��g�=��߾t��X�� ]�]P�	���f �;=�/H,F7���H���ӟcŐ{Ѽ�݆fBɀr�pIX@��z������R�gz���^���T�A�Κ���5�~�_ל�) �����u����E�(�!a֦�[�6\d.�Fʫ�D'tI�ӌ\'n�5�X"6q�-�,�:f \�?m��p�bM	�� ��α�8]�0Y�!��̏����!�-�>t'���]Br�}� 2"Hkb�qz9Y�%p\�A8��IU�A`-$ ��󮶠44~}�Ӥ�A�����'_w����g��'p��v����z�İ�����1�塘	"��0�-�0�l�w3��/YX���S�D3JL���#������X
��1O�xM���
�v�8� b倂��3�/PK�ǀf4,�A(,}������	_�]M�)$F���Σ1^�z�-�Ĉ�~���4�inb共W�7z���z����/��}��&@��A�d��ާ`����fk���w��9o~��h�
�í���<5bo�(}<�����r$C��I��r�b7�x?|�N�?�Qٛ��y�x�0�3<��'P}a�^w~�ř˂�:D�-ݗgR	�BC��7����!i��v�P�"����I �z.����A�g�8�p3?s�ǰ�_e��٤� ��5φ7_�zD��K(��t����sh룔4&�1�z���{whnڕ���:b ?�x~~+���?!���ʱ��!ș
���]�`}n�����D.�A�4�!�0Cd�G���{nW�6�o�("��s�}޻�����t]OX9���p �� �� �,�5b��P��LIrO�zd1'�g�3B�����a%1`��0N��;��[%��X���KsY�����_^��t��41>e=�- "A9w I�̓9E���Fy�'{D�	��E���BL��D��jc͝��C����5��?��PV<b��x�SWy���[�BR �Y�"HʝCz&Qm�1���@�$�ߠi+e8t�~��a%����'b�nHIoc�#�s�b�#8���JE=�5S;� ��S+����J$/w������B�^�VS�w-L�sJ�LV�1u���o�@�9[C{��W��3N`��>�|�c�\�y/g���/S���&�u��y��z�ᗿ��1aU�����8���&�J;Pjl�ؠ(m��]Uh��3͹^�|����n7ķ}r��?f�a��Rx�ź�cOwv���ۖ"��bt-���&��ugp��2kY���ة��9��۪G����1������+�]��K����,Ԗ;!z� e[��ܛl�5�ʓYz�;��u�#&��]tf�en�k
�X� �ҋ%mB�h�v�k��}��')�옟]�強����|��mq����e��E$�{k��:P����,d�MXE"����ҊxPPq�'"_� � ��K�,�%��&u�׻�.�x?�}�n�oyᬢ�An܈ n�K���N�&�<y\� ${�{�0fj^�@%��@��M��SHpj�8`���0��w���.Cyx���4�j�����=>d�I����pK���>�s�g�%^�)����	D H>�pIxC��&�&����;=��z�����)��!+ہ�3�:C��Ii(�޷7ot��^쵟��@��$�U�� �" ��M���m�����H�W9�k�L���� �K��$�bi��ϼ�@^n����^y¥�Kh�z�?��煦�1]-4B�5	�)��t�m��٣�a�4�Q}����
ݥl<�w��Q�"A,orx�g�$�3��R��Ť�����x�zA�Z�"׽es�3�p��!�-���S(�bp����BJ2gtu`|F�9��+��8^G��~>��%�e��z�x��]+�9�v�x�w�/��%�ǝ�u�������a�f�|�u����)�A ���$�$Yyw))(�x݉.�K��)_7$H$�'��K�0�1�0(�y���p:��P���@(y�H�U#zr�I �x8�Z�6#�*� g�f�9C&{̀Q���K����ؑ~�]�m1�l�~٩jlK;�z��;� C'pn�2wۗ�%BDB>���y�%��q#YK����B��dذ	,���L����x>eE����'�N�x�Hߣ��]�������iN�f�����ث:��Ew51���5�i�����PK��I$}��R���]�G)�(ў.	�
e�] ,J[�"�]�W�̤:��@��Y������pdlj\��K[<�Gb�����-��=�.� ���		 ��?%��J�}\���&o���7A~��x�8���3���d� ���RJ	x�/F�ҩ���}qK��G��w�����j�W��r�����ٷ|���M��8����g�Vy�t�2j������.��~���O��00��ԟ��{�����*A�w�㒔�ǩ˃�
Ay��=���꩙�D.���	 �5�<��%$:c!y�8	w?J�E2����7Ig$�q���w���:D=ݲ�\bBI ��ĳ��j�yC=�@I�xY$��>�"Y"i7tt)	{�d�e���mT�!)U����=-ٲk����㊥��7Z.�l��"�H�+�͠�Oߟ��靶Ð���{5-bA�??_L�4�0-���L�ҫ,�'�ٌJ�	�@I ��% �H9���A�Ô��ę��'gCB8yװ���>#4臾gj�d� �di�`�3�p	��Ф$���q7p��ۭ�����`��Ӂ$IH�:���%�������BB;�gz������S8	mކc$;�$Uȃ�'xpC� X��?z���3p�i�߯�@ c$H^t�$������>޸�������������w���ݩnYҒ|0{�_=�{O�d鶨DI��ɸlg}�D��E�.gxc�p��b��|����c�h� ��c����ɒ	ٙ�y��E�#t�pSb*�$Uu��2E��S�U:�\$�}��E:&�{k���n��U��d�z��&�;"�w3t�8ّ����<3�X���	�#��s%�V��a��e�|���&
k�	a�TNx'��mk\� O��,$e�M�k%��"���imd����+1�o�9y�$@>�ɐ@ � �� Hb��x�Omo����ư~�d�"�/x���Ɠ%h	��@"��E�8W����'V�w�$�$1�� ���Iu�5Le��R�Kb̎G�)��gH=�2
w�~���1��0�	c~$���,HvݿI'�!tn��$�O�\g����{�1�d���ZB�1��Ћ	v�G v����wq���7.ft�D���U�YO`�z��5������e_�OD}�	Z[%�gTPn�y�Ep>���|11�� �>巒�D�OS2��8�q��p��A��a�x��S�b�3�2�3ia�����|g$�����7aم�4�#�j@nHQK�Ke��t[a���*e2D�[�n����ֶ:��O*��Y�+X���L�v�	���N�9^�r/�4Vw����d�0%@��]��\�Bݳ�Hq���Z�nst��Sc�B7�D��.z-n]5���r�[��H>����\B����iAڼ�;�t�$f�Z�a	�w�vrЁ�[��f@0$y���Rh	n����K�`���,�`����A A�2*��H�"<#��`:E�+-����V�I^ε���ن8Đ.�,s�@��S�B|"k�HS����s5����z ��(v,���2�mc��Xݞ��2dA3�ښ��
l�CY {�@�{����(	H�2��3���bۘ�A�Y#�H�(�ϐ�j�������������-)��I�wf�wF�# �7�I �]�p>FΨ������ �k� H�Ɇ^��L��nu�G'����͡G:<�U
O�swf�;hTZq50�y[��&�)���b�v���r���4q䊈A6����p J�j͉,1�9�/,�\S�'�#�e���9��-��ҩ8�T��0��@�'=,���?Q4���њ'x����z�
���t���֍3�~�y=|��+���p!N��.z,�`*�3����M��,�Xf`�c��� �-�|cG�@O��9��9����O�O��w�H[���}�t�E�~x,��$�/�����ϛb��3�"H��Ǜ-C	.�ݑ6�/{A����<.��V񪝿�] �I]�.�ʙ 	�ކ�P�@�y�#��1a-W�0�(	{ź7� �; s(��yz��/k�5�&�,�%� �3�CIz�EDG�+��Oz�XBN�D �?{�Ю#���,k��,�,�*������"� �ӐWټN���;�6|�҈.ŝ���@�P��2�3�w3�zEI���$�w�K	2e�_�b���;�K��<���Cq�NzD�1=c�b|Y���p���k��J ����!�ѓ饝'�M�2ݠ���X�	C�T��-
.0�A ��}"e��@V:�}x�S�z�b�^EA��}����n��r��{�Yۇ�n%~|}9g�%���Q��5L����G��-�oO��s��!�"�̵��Rػ}����I.�����)d��;�*wk`_މ[w��I �.�>�a-̐@!O2@0�w@��#��/�ōtz$�$��uчxOݭ�3�!�R��z�$��r��=y'x�S8�ކ�I$c&���U���oY���0�rɩ�N̢��I�'��4chGC���J[����Ͽ��a(.��Av*}��@�Tzy�� ;���E�{#+�K���L���2@�_SP�X�h���Rwr`82��G�[HX����T�ck���{3�2N2`�nd	ކG�����CY�'�
:��.�$b!�B�qՂ@&���&2�!Кv@��� Q`A1����8�s���d�D���8K�y��+�N���$��X��>�������β�, û���mK��	x������]'��&����y˞��Z�y.�^w�����=����x�tMu�T^��Ec���c3ᘡ��7�ZN�?��gjY"�X!`���a���f��E}"m�&��R���g�:PS��ǚsa��ƻ2%�*7+��N6 �+��$C$�q,�����.ky����]fgL\��S�݊Ɵ7~{��_����ک��K�h�(ȋ�Xhv�b��j���;�rb��#Y�\Iio2pq��2 e��tQ�hoJsX@�L�cR�m�0�'��N]]��h�D%�$[ty���}\�p�15�r  �-ΖĂm��!0=��0h\m��&� &��Qwr`841C��� N��A�@>�ؑ���e�E�Y�}��	 �n�Kn������������ �m��'��g�Hc�Q�Vt�b��Bgx @ D= �H>�^D�B%��hF�L���X�s"z���L�!���_eI �A|�&f.��}���x&ŉ6"-�������>T��d���?��=���Y�q�o���/���5��x��:����'e殦ŉ�.������v�{s�N�ɺ˳Wp�<\Y鐝#W{ٸ����!�;��w ��b�T��v�i��&n��� �~=i���<�{�X��7��1�»���<[��;�Fqx�OF9�7����3\��l��wޤ\�!9�Oe���3�z���7�t7Nl�vRL��v&�A��7���)���ws[
�H[����jׇ�Z���<|��ȓSB罋s��Sڙ��x�<1`C|�n\�5v��s}��0-=���C^/:���}�p���nn���]��`w�#7.!�K>fy��<=���xy�Oo��{�-��,���6f���}%�s���xf���*;-.�7&���O_N�^zs�X�SFlTok�A%�oU����:-0��eW��E{��R��[$����U������w�L�>Ώ��`3�W����a�]�sƬf]������f%����W���S7A�}� k�,Z �b+���n�7�y������瘸�窘yR�E���}�nI^Oy�u����^��ۢF���<4��#GF�.,>�A��K(��#���d�sб�-�6ir>�� ��gң��ђ wsi)!� ��u�=�l�ʬ3�<���8n�� j��mJ���	.��f��fM	كe�
���R!:�>�6 `�"�a�'E�vۥ�G3�Q��7�9��(��F�i��e�33\ٻ�[������^̻��� ��{��l��z��:H�5�eA���*�x! ؔ]�T���K��m����ҡ���4^_�|�����Ǵk�٧ľ�Ś! ��刉��Y����/$�I�'�ȣ��~c<k�sC?g��W�M��y�S,�s���"�]�g�`�NKq?����K�~�a��Q�4�m��ꊢ1�;vd�J��q�wv-�YW�6�[-�u�ˣL�ۘ��֟<g��ye�c(65f8�j�3n	������?I洛��3��ʎhy��&6��
����K�u������jrGQg9jQ�MHD
X �2�m�	�-R�*dR*�wvrC����~������*D_�Y������sB�?q�Ӑ��)�ﮎ�C�:��<g����grg��~�f�˗5j��d !�,� �# ��"H֪�09 �9�� �VD�\��}u��<}g��������8�����ċHE�8��qLt��:�?T#�Vu��H$g������*��V�I����<}g���Ӯ>�㏏oY�wV�#�R�܋�iʠ	�/2���-�A}������F
pBY�>�,b|��}�y��ώ?zu���>>9�yr�s�;N���byYOVK��R
���^`B �H����)� �%�ӈ wS���}x���8��������||~*w��	��w$�J���8�,x��z�c�y3lH���E9�ryp����<}g��ק__�>���y�{��c�H$X��b�C�z��ypB�I<���Ŋ�P���~>���X���wB� ��@���Pb��0 r'����Na���RU���[b@R"����ŋ�R0�C	@�ǈ$�$��&^�@�!Kf��LAC�|� +�PF5BY��M�X���'�{�߃� �
'c�;X��4TU�jw9x����w5�	�<�l7"���=�:�]�.��GMl�.�:֙JCu�,�tmԅ+B,Z�LQ�@cT^W���m�����!�rY[�9�㧁x��v��Ivw��p�[�<exy6x�6�E��m�X��k<��W6,����s���y�8����P�C
i�T�.V �竪KG0�0ہ��'������;���85�oG�g4�a�Y4�k�uƻDpx�f��a`��Zւr�s�����uyc�$g�����S�����%�X蹉���ܮn�v��=���E6˝ĈȖlBV]�lL��Vkf1�ܻ`v�y]��^մ�:�l��ōs6��6hB�f�����SKjS��ll�=k;��o���ՎvY9��'��-�ef�k�����#6�ۇtm�K��=P�&ܭ�Z��xW��G��,�w\'j;OG,NW�y�s��`u��%VË�0׶)禵�ݮ�v���E���K`�'�`ݑ�����v^_5�KMtg��r�Gp/k�(�td��Y��g��Xn����n�	�E�F��\u�7��ۭq��Tr�v�L��b��t�:��qڸ�_! �'3�v��ncesC�e˫H]*Zʎ1mf�l��E6emt���6�K�t�B�0��g=M��vns�I6u��延Y�Kvl6��-el �{be%�M���qZȚhQ銘�u��&�˻R��{k�n\j�2+�q�U�f�le&å��:.�;\�i8���F�lL�lRk�b���d+n���j��Հ	o�N��8��q:Bq�!�a�>�U�O}|��u*b'�������.�[��5�\M�dƣ������h�in�5pPΉ��0M-,8ӱ,���u��-�z]ó��s�ݹ�B���1`�R�,,�C"�l��|�ȭo�&�潈8�SM���4�v5��i�l[Rx�J/6�nѮ��Xz:���s���\0�渳@����Z$k�<���k���
��w4��@����?�����LGI5|��	p�p�	��/����3�E�C��q��B��}��5O�V�me-/��$o]�����(�1�ۙ%��ޤf����kp8����X�%���H,A�y�B�r��4�^�
0R-������4X��.ZK�drlצS�30�O(	d)��ސ$-�"%�%�n݋��0*!���X{T�Xf,]����{��X��)��"��g�$)����*���jb7,Cy1�*Y�dKy��D2y��7=R��`�����{a�y� )�}��)�1���$�$-�Z�P]����i1c3v<�/����?,V|smLv���\v iy�Eh����La��f���P�/�����[��h�ِ@2p_odH �G/ra� S������>b�HLB �ṯbXli)~�l��.�`��]�M���;��k�w"����ʜ0e\b���-�6˞�23̰��kx��hP�|�g�G.x��C3FF~��C\��3�B]�� �Rea�!�HlrOǴw���@ O��I�b��LY��~���`�=���A̽���1��S��B,]��$"� ;�7����0���bI%��Ł�JS"��&�kl^�@�`/c��/OfiZ��H�}-Լ�@;���*d���M?foK����0�KDd�,F���wr`8>�]L7�vd~A��6$��k���M@�[��2~�A`s��"Ҁ,����$2w;<�A��{Jka+Y��k���Q��W�9�h��I��s�����r��C�i��d��e��CP4�=��IleO,��=��(�-N�S�����6�T� ��%��`L]ҤN�w
R9���멐[����n���{����4�� V+��bx2 �z$ ˘t0�/Z��n�ʐ%���y�����e�!�@E�̺� 
c,Qb���%�7�f�֎�Ϊ�>�R�רl)�9�X[�k���z�Y�t�x	�)�L���
���j$&*��&b(���y�I�G3�:��/�eBP�E!�d�	��y
��Jҿ}�zK1 ���@�@�Ho�$?�����1+Ś}�9��w��,��0�'X�ٝ�D� �/�p�5>r�ov/2�$�2`������b�x/��hi���bv=T�؀Yk�2� $^F�RbS&D�c�6������x$���[6�$7#�a��R�������k���R��ͷn-a��A�!�~���0T�E2@P2G$bH �@cډ�,F��[;	-��7�t�$aD3�=@�e���05 �@�*��yL��Qb{�1 �4��׹�� �V�;6}����ɷ�h��mZ'�;��df D�l���H�p���)oHѮhaB9Q�Đ@-y�2I ����W�����xAb��[��*٘�6���r=I�혐&�NAj�ۈ�G�Oų1�뜿�򰺷����{�jٺ�v��Cʲ�&*O�ޚ1��N�2�!$��2R30�1fY��
r^�R^G�����qfD8��kkfA ��/��"([Θ_���ɍ&%����+ٞ�4OFm>�c�ِ$:�p�/���
 �����	7yz��9�_��ܓ3���2�.�T�amo��M��W�8�8z�yn3�5��㦬�]�R;M�.�iWX~�Ͽ�1� �o���d�E3�ݩ��F���0ť?��Z��s�l[�I�����UH=�N_`���������X�ήj��fz�,�Y 6����@T� ���j	����N�ǋ�����y��nm��0�@�P�.��H-[� ��	W#�x������ 	 =f�L���Ѿ�LY�j�A�Z69(N�-vZ=ճ�2��v 0igrY�z=2I����b����̩�x����L8޾q�����;�J�7g��ۊ�<��׮r<�c��t%��ȶ5�Bg�8ɡ���Z�Οnv��t����*9����]��������c�׵Z��S��)���7xf��bқ���������N/n���j�b� �("�I�H�۶�5[�d�n�n6�����sW��p�%0_ksD�T���pB�6�o��xO���^���v&�}���MJ�N��N$�N;��$N��C(!�.VC�~��a.eo]�,�z��d23������7g`�5�˳�7`W8�����W��$�'c��Y�el�Ļ�s1��,�V��ܤ�(6D�L�����ґ9�m���F�=uǸ��vR�:A���f��Գ.��R��=���܍�1�( ���;�m|��x-�ǭT��L��\/��f�m�2�t!��y����K�F"@����y���K�\� w�bXw=C���f�:KKgl0�el��脌"���E5&�m-M0o�3��~X��&"�.�KHD�����>5q�f�����U�"V�w	��(� [Ӎb2��2�C1���ow�n,0kl�� b+a���bl�S7�ü�% �=�K�9���գ'O��V��	{^��,�wL�L��TK+pVt�v�K�Y�z�@87�=�J�%	��ƏM��${f|��N���[2b��U�]� ��\� �K�t4�v����b�N��<h�K�"��$����6�!l��vm�'ep�w7MV�0]�nc��֭�{0SY؄%�IϿ~�2�b���	N�(! ��\��pɂ]����_?r�<=���{�A-՗�o/�xE�"��&+�"SW/gk�'�2����
}~���e+�#2Oo,�c�2Ps���f��D�`��囸���D+��>�������go>~��`HdW�B�!�P�O;��e��D�v@��Aw�;@ƍuG�7컺8w<�An��`Ð��mp�y�O1�� &.$I����M!{
�r���5��$b\�Qq,Io7��r��4�۱ ���Tż�eʝ6Ϸ�DD�V��Y�{ I �C�2$%�������C��`�X����@�e7�*х���T����؀@�83����,@#��s����8S{�1�@�ǂ|����w��t_q��hY��J�T@��c滾����ɍxhNq��#�]2�QJ�\,Kf�����O�Bv�&[y�)��,h1��v�+�u� +�����2�������-0'�R ����v�xq`c��� ����O�|� `���.�bjݙ>$��_�5$A5���,��e�j�6ٙ�<#�<x�"R8�3,YR�1$�2}��h�Ǟ���P�{oA�7�0b�$�kL�k�������7��L)%��V�����Y��=eN\u����{��Z����?������!�dBP�P䊟$S��{���m�lY���2$1|�@�d��u��"!�P�6�ދ�z���Fe� �7>��2"P�!�~0�̐�o�Gf����v�<�y�Iw^��xb�I+�f����w"�a�S�7 H �w0�F�&ݎ�>���J���s6~r4�ӭ&�i�2{�?wv�M�hi��Լ�p��a%h��̨�������������Xq����	�~�a������[��Q�8�?���r�Ȁ��z�@�
$�}~��bP�D92,���nd[)���\ǝ����$O[�ZYk����1� C�w�A��0a�y��k�N�C�q^b�2��O_dH &��`�T��A�D:@]1(�
otm (�&@&�]l�-q�a�A�t�^a3ۏ�Ѣc�u��	^��$igp2��	�	��.���ǙE�@�y�qy���q��}�sw|�E������p����Ny{}�K���;Ꮻ�;=�s>y�ߧ�K����vyp�|����~��82/p�'C
���2�C )�@8������xOV���"��7uz���M���GV�s�Hض�:9���_<�	&���q�� y2�醑�b�r�V3���E浛5n���$�W�'�5\l�ݷ̷A�ܷ\V�]�u��:78�������5|�1N� �E�+��,i�2gz�X���^g{cj"����0X�x A �L�{f@,ǚ�|:ф��6@��L���®�c�h`|�B ����ۛ2i�&$Ϻa���U^b���X�.�L-d�T0�tD95@����b1$	{��@�.�y��d@b-�Rr�d�$=�0�E2Ot�U6�o<,�g�0��/�m�#��9`0����1D$��d�,�!�6�q���?/3S!��-i��aY~�
xw�F&�����S)��W�l^Xbm�!oސ��/�XK2�ANr�hem��C�U:��6����[ �D:M�ϫ��1��(<g��'"Ŋ���5��	��_%{}�	t�:��ǈ7����|�I9�wݜ�DLA�ozk��U�wp��Щu��+/ۓ�\�(G��D�z��upeP!�U����|�u�n9�hE��X�(��Z��K�J��:�nЃ �7oc��7T�d�n#�.���E�M�i��Q^�5a�3]4I�Ykh) n�g�rز����g$A�z�Gh�d�Ŵ`�c�Q	p�*ъs%B��7������Jz�����`n�1����P�fq�"�7��-�h��v.}wf�\���)�=����|7+ӍH��U�Мg@9>�� -������@"�����3�aY- ��!�9x�MPuF->��^�����A'��Dh-⭒)�e��s��[4� %î�8�L����!���`��@Q �s�$�cZ�f ���B��U�aa�_\Kɔ��dA ��������b�5w���R�}��d�F}�"P�b��RX�(���@�7��'� ;8���wV�� �3�aw��$�U煞D�C��Y��&X��q�v\�1b�d#���vEKNwn�{��ȿ}|��D��1шq�b�{|��dx7��f[.K	Yb�3XGٍ�m�a�[�����BF*��6��X�V�� �%l[��|{�"�_u���,
I�n����M��X�Ҁ������t�ϖg#�j��M(ɪ�
��nF7�zv���C�)���;��9��s�_fVx!TMڭ%M�8>��zanԜ���î�{���s�������'�S�"0�ԃ��JA�P0g 3�4w� �@,O[�@� ����)�b�e�g��y�0�8��� �ge�AÕI�|	�&��)�T��%�ڝ-b蔻��8$n��"��X����3�d*}���'������Kk .��!���A��X�5�bC���ۙ@X� �,�Ő*:��/'k����G0�������zuVBO�w��,$�=��V��0v�(��� M�D�2DL:�j>��W��>�_c.�X��P�n��*�̾��Hm�����G�:DMZ��@#�x?g��!v���c��8��d��������@x�Ig
�����XA ��uQ �o]ޑ��A
5�����-����W����F�K"A=�XS ���)� ?r��Lw��/��^�6�Ҁ��6j[�\���E�2f`�0��׸�b����A�E�N�c���]Y��	�ɯ=~q�nOc���Q���ͳ������]�0�}@�x����r���9<tl+���n��̻����B؞<'�n�/�x�,��~�Y��Ќ�|���75Mξ�q��������-�{7H���[>���vw�ޯj޼��x����g�2���BIlU=3�3��(x��HȌ�����O8";�<������ڳ�H�vv"�w)�睓+�}x�^g��zl��������>�ozyv�@�zh����c ��9�_Ssb����W&�Ƚ�F��u����%ln�+�؞��^�;d�O5�7�9@�װ>�^>N�1�L�aY�S��R�{轀��w���z6SP,���F|V{O�Y����爬�o��G;�n�2�l�
[�1��o<���a][�p\8=~ԡ���O�~����q᝛��j�����{��<�7�B8ڑ��{�8rաw���0����S'�)&�ݽ˷���b���x:{q1䅯��OG}��zf��᷽���ޝ��{�7������0E�Ѡ�`�-,$xwnM8�ڍΘ�g�g -=wo@�~��iE��Dy����~ɮ�޿�Qp�v/2�a5	��N�֛�qM�~)1�{����e/bvr�77�2\j��u������|��-��:{�93�3ͯ~�TpA%ʑ*%�a�^:����ѐ�:T�Y��E�kZk���{^��R����H��&I$D�("�N��7��l�2lb��lkglmn�3���ܩS�4 ����>i��E��z� D	zN�ke)I���?kI1|������}���~>�:��q������q�sy�a��ZT���*�U`"u�:[uG|�G㏯<}g~�]{}|~8㏏�x�s�\�9�p): �q,!�J��z�^a�b"���G��׏>��?_^�_�w��y��x0D�&%*��ƌ>�X8〓íd`$(�'.���׏>���㮽��?q�Ǭ�*xt
D�%H�@����b�!�,z��>ν��^3�?~�_^�_�8��ᇜ�y���$�R��!N�	�n��H�$ �H��#�A�I���A��
��DL��2� @�*�!QBO���' �����pcĒ�1!X�,$`+5e�	`㗔�"����p�|��I�O��;���
p`P�`��"��"�M�����ƠH�M�?T�@�@��&K&���t�1��Φ�� [HD��:6/��i��\N5����q��I���"6@�>��D%ۃp"�!�%]�ث�,.�B ����r���a��^���(b���\��r�mu�l�H�������:q��d�¬�>ƣ����tg��n��:���X�ffط=�R����'$C��p����X�
��	� C�[�� o�*�Fu��ϥ�u� c���$�𳌃�!H�i����,�f<�<.ك��i��$��	�$@���F���tF�.��5���'	�:wYwxDN"Q#)�cX�O^<1�,����~��>fleq��X���X���s�om���]P�{6궎Uk� H m�L���<şA$)�s���ڽ�{��[ʉ�W�_/3�FL�s������Z!Oc'���z��J��Kۓ�ތ(}��Y��J��p�[z8�	di��L��!�R!���Ȭ0
�z��{כ�̳֨���;�b	6��`` k�dH)����+�,]�K65I^�bǻ:,������Dh9@�r�:Q/!�*������mw��]�Z�:��䐥Զص�NK�-��ֻ�ʌ���E]W���߆�0q����$��^�4����t���]z�*�a�����87y�z}Nx��My����� &������2�&i�O�$[{:d��E߽� �>�������yc2P��e�L����Ld0��m�z����Z��$�v�CS$7w�Z�i��Ƙ��C�#�ݕ��5:��P�tSq�ji��ɖu� 9}��Dw
�xb1����捺щ!C�"��l̂n���t�j�9��pZ�n.NG�X�$�{�@�秨I{�;��qO�LeE���Po֫.,�yY�+�TH˼�����X�Y�2�N�N�׏<�].�����S��_6��c,~x��ץ|5��A{���.�uLb�̈W�5��.1�)��y����lۇ���׉�m�k�IX��[vl�����O��	����*�`T�Gff���Ye��㨨[�r�tO2v�����]��U���ʑ���٧pg�����On���L֤����!e�vQq4�, brn(����s�;��^��;�ⶓMj��wj|\6�4D��Ƭ����5���;��g;f�ޑ)5�un��G�-��W�S*[��t�h�]��[����eH��m���c.�"��?~����A� ��G߀m��E�
��&�|I1�u�4�u5S;+�0�wج8Y� H��,u��P��"�T���.d�e�~D9~|�O3I"�v?@�4�tv^��۫�z%Mk=C��M�OUy���ɻ�ۙ��\�.�M�=g��bX���'��.Ŏo\��W��1P�#�1���+����3�{�	ld�����$�mޑou⽞��1��a��u�18x���fZe� ��q ��GW
!g��[R ��L�b黮D���}�t��x����D;�:pY(rokɵ�9{6�[�Xi�ۉxI�<DI��$�@uWu�zD�X�{"@$�[7�A�:w�jm��ץ�YK�܉",�d��`t�f���禔Av۫�IΔ`��vU�픣��<8?���h�~�q�;׼k����?�@�}߽{�jK����p4����� 45��+�:�����!"C x�ԝ' � ��(��  �tuț�ֈ�>�$����h=�ow������'���
�K��,��LEr붦����xF�<��`�;������~,"ޥ���ɧ~�~�Ӓ�+��-%��נ4�hd���:D�e��8rI�sg�]X�y��dKT� }��W1P�#�M���.&������ c%��<Ɓ -|0��*l��gM��j[9D��2>y�q��:9����#�=jek:k���Bޯ8�쌕J�0������|�����xk��KE\Y��'=�"W��[qٸ44יr��� �J�}���F <;�}�Q��2�����͝�E��{b�+;��;;�SL;�_����P-��X�'�rà��xc��x$d����h̲LhY��q�05$��4&x}3�z�ÚN ���z?=�����}�1��>��1UH��x�,�0337���@!�N�!82�����DG�x�w�ǜ�w���/�律Ж��y���w ������w�ٖ^jh~������\�o'3� �j���b��\���97�8^�����J1�2��lާ�{��m� �[�^d����SLy�4!3˿TKL'�:�����$?{�I��c<m~���;Go�}��ƄwN���޲��9�亸٫m���������̺
�}�ׂH���hd�$���]��7���#n�ǁ̙W�"B�I$s���@N� ���+��6�|�E\������,� O�:SJ �ވoU�u����@�P{�woE��@xwJ�[k��6�@���i ��@���F;G�a��4n˄�"�6q�N�S1<۽�2vxc�O�s5���$5�zG��"��Ɓ;�*��B��)��n_����R#���z\�#��t�;�E�Ur�w6{9ַ]\��.��� �m��p5�&�r|�"�|H!��x~§��|���!��Hc�(peT���5��ܜ�w �s�ȒS%�e�ݶ�%��y�r�$Mw�@$��ݑ4���m~������z=�E�.��wg0ЏR~馳��JJ���0�Rb�t�Ip��+Ee����>%ȩ�#�����@��V���S$@=��-O�{�C���R"⮣ȂA�ّ'��gڈA�
�s�b�?�����X&��f(d���{&A%6w@�NFʢ:X�?��$������ ���c��v����@PK��}�e��I1�I�e2Q�I�{�Q��*�sznoۖ|g|��F���vtA�^ΑC 7w��:�#x�G�Sj�n�bq��,:d����^�,I��۷>�4�<�����I\}�.m�t˂4�����kc�dN���(��o����iGLW����q�*e������G�y�؏\Z7�xn�n�=�3���i��s�������^���kj����:����ÙI�3���kg��4����c�W�-C��%4iޭ��d�>� ���3������*�ȽH�/C
�bf&�ŋ1^�o:R�6��&�Cq����rr��g�>�s������+��;`�a�U݅!	Ff[6��͝P�IJ��ښ�����0�!-�B�Yu���j��/�P��;G��g�� �d�6^�<'j��m�	���Fx<����\m�Nsn�n�nF�8��7)1bB��G�q�	4n<�H��LY2�pZQ�:|���y�.���l��Ȓ<�^�q%����hɤN�o��9��&�!���st�K�8�)ylth%�x)R�s^�k�I!o@�m�-�,$Ύ���[&f��D�s�� ����}�D�3���I�����<<ܒK_d&:�A/�ʨP�
�:;�T��j����#�N9�֦<K�xo2�=䦔I+{�c��*�P�0���N��W{�BP�"!�fd������򛉊XA痿�Z݁"c����_L��x/�3+;��y1��\=޴`��e���QՃ	�9zƲ:�4v�˼���RPR�]Wn�tp�w�qm(�O�`O43�\�� GU�W�.������8~x|�wz7�<)�����@�+�Z%�q���c�TܢB��k+�x_G��w�5��zs���7>/��]���
�rtB{�ӅU����x��Qh����Kkc0.C狆2�p�r�����T�ʌ0*C
���J'R�(�@`Y�m�Oۛ�L����@ k��5�Ϋ��=~�O�
�5{�<x��tb�~ikC�ߔPr�w^
���-׻ ��"YG]ԙoM���s\B�7g,���n�-?�y�~M��|z`���&3�2���'�'##v=�=�<��c6xN��!�CB��w�F:�A�����]��뻩i`	cmy���vr�l�1@�onf5_�<u��G�~O<+�|&<v�nZ�Ts�
Cy�ۍ��E�룞�]L�m�ˢ��R��$�X?~~�O�C�xw]�Ӟ�nd�1�ؖ �[� �o�ʗ��d��A?EȓH;�v��3݁hOT�e�O�k�Go�<�d�!S21�m��,s��ƒ���O��|��E���ńu��t+ ]D�Je����9$��ʃ�C{�Ҽ�^*,���٪�" ���?�sq���^⏲n����Z�th���q&wpφ�i=�_��Tއ�ܺ�IQz��߁Q�2u4��~�D���dRA�Da��+H����?���BAib��>$f1$�M�?Cø�]k~�����az��v�d)��D43��2n�`2G�:g��]�b��/�+���3�q\B���Ds�p4'*��"*/;�$�e]`k"�ot��k��7�
����skb���N ��g�c��P���-�	Y�f�7<iA@zJN�+�%��s
�h[�ʯ��5,e�u���(=��0G<�Wn�\�cX���F�U$�s{��w���什"|�l�����j�N�m>�g>����������?6lLH�� �.�,)'hg�<fU4�qW=��@&����lS ��!AEgoL�Y�)n唃������e����>�������d�y18˙�&b:G�U�;�4N?�ç����r�ы��ɗ�*s��4�Ϫ�+����7x�����޷<x)�;��n���n�ߪq\EDA�.��]������i 0�,�C0��a^*CKB! Y� 0o����2U��s�s�(w�%v�=3�gi�����X��fv�	;~J,Nu��#X��H����
�̜����w�Q5vx�l�rQKt%^����P������P���Zʠ,^������U����N��yA��2��^��2�[��vL��I������Z�D��7B�~���:��� �I޸c�z�v�Mg��Gv�N��ww	��wy�~�&� b�fH�H��Y��
� ���E��$L���XI ��Х�ă����I�0ї�:���km�6�<�/��}}������6������n~�����% �( ��x��$���/Vgٯ�YSu2H(��&A��CXK3�P�[��w�eމ�����E(����@v��	t��l��Ϳ=�Ҹ<	�93�6$����� i}=�G���p8;��
ܵ�(�G��1�w�Qo6J����Lq_N`6}��g�A|;��~}2og�Ӵh
n��=�e�q���W���7���/�M�ӹ67���޽���5<r�g!̍s_xM������!|V�0�^�bN�׵�1�������ܳ���d`@G� ��i:��Uv���˝�=է���@k{���� �������pm�ҽ���C����{m�/�q�	�s�]�O훇ۼ�`���Z`:���xo{⶛�hO{q3�b��rb=��z��`���C�}�ݤ��7��c��
n�T���z�x���/d���T��_�ê��}S���r���ECs���<�IR�PN'�8dӜح�p�[����������?'v>���gw��%�����l� 7y�{�z��%ݨȦ���zo�������Ȑ�����6{v60�����]>;0p�<nOnU��y�n����1�$F��tV�嬉���}��k���y�V���=��GZ�ii���`kJ�C���)�s>�5��WTp0���� �|�;�L\[�^��i	�k$V`#*0�&*�E۷-�8��×uȃe^8��"��1��K8P�1k�+���sS7i�����]|w�LGM&<p�I��U(�F�aH������An�X3v&Iu�E�:+�O�;^l���/w�4�h~��SG�X�!�&Y�@�^�xpzt����'c �)�l,)�"�=G$�&�K\�[�g� ����uB�1���9}<��h�F���˽}Ś�`�}b̍c��~�0��竛���?|��g���@U�x��c�<�Ֆ�3[�Ņ������d��q��@0��fTe�Č�&�V����[���}�N{oI9���l���+�����2�����N!�8��T=��u�?��~?u�����>9�sx�w�?�����@��h2 w(���s~�[$&o��w������o���q���9ȮG<y�����:
�+Ԑ*m��k����	���L��H������׌�ώ?u�����>>g���MUH$�N"ȁ N���x�I�#���w���~<g�q�㮾�>?q����g9U�{�M�8ա)��c��8F\�p�2Uu���q�>���㮾�>>?q�2>p���Q���J�A��ϵ�	 ^�!~���8��$d�L�Đ��ű��-mm�������8�DC��#�ۨ�h����|����Q#u����x�Z%5��D霒cB�H�A �1y��^Ձ��1��>�wz�a�O$� @��O�i�,�,�F�f�`��B>���o�%�p�,~Ò���hN��FC1�H��� @�!�5�a�i��T#�":��
��Es�mZ�7�;n���	�'n���sv���Uq�먝�o�p�.��뷭�^TڬHmh�u��Þnwn��S�Z�@��l�.�c.�k��Ba�.��A�usn��ݡ�u�E�A�V/�p��L\�o���˾�q�K�cl+Aj�� �Жƶwv��Q����v��C�F����gv:�v����^wn؛ D�NFm�GnaFԹa�˳jXCH��ؕ4�]��t[6�Ћ�+��w7L.�e��`7j�G��ჲ,�óX��]�*��a�DlrI��1�y'�բL���eV]U�����4\܅Q��� �RI������*.+����2�v�1O$��r�zŴT��r`�'��3<��6(y�7G/
�S-f킈���4:�9ͳ�ڶ8X;�Z7n!��L�q��&�#{*P{E�������j�A�2�@h�eҗ6����ʉ�,�I��S71h�i��q
�R��nhu��ҁ:��q]�d�����ֹ\���t���[nMǍv(.��kv�<��L�Fx�4cX��ƥ�������7��;7M)6fa*饅6��䉵)E��PЖE��������7D�32�0[.���z��GQ=��g	æŢ���-���b�N�C�.)��V�;�m���-���h���f\�IB�.{3�3q���v��a֍�a%��|��z$%Kz�3�f��a.�e��|'�fT3��ԯI�b�X.��P]V��v��:��M�F�m&l���,\ʗ\#��r�2jq�2��Z.���îr�s�~��`W������ �Ȅ0��� {��ߓ"��zś���e�oe��=Y|�@����൝ޅ��Ӟ����k6��˦-ƚ#�j��Sp��Cyy{Y�s��%����`=�d�Y�*�k8��]s��<�N]FC�Қ��v��.��̃K+c��c��Yfln���.c�����}ɨ�F�c�[��s̝h�*�y6�#Ɯ�ܥ������?�mRF�~����t�L�1��%73��ܝ���mv��޶�ލ�$����Tꛮ0�ҝ�9q
Eك���|�w�:16����,H��D��k�a�]l���u}���I��I$��w��`�fz�fX���y��ʈr#�;c%��1��L����JrA�^ᄋ����:��F��z�z���YQ�ݙ�)�&�~"`e�f��xU矤�dN��S9�&=�gU���E��e���ƥ뎉b�T��hoA���Ijǳu�#��B�����\�]�M�Y�ںݞ���fj6玪��x��痞ٵ�zP+��';�Wd��#[�����)4��ޔ�g��|�ra�q�c�5�0$�TM��%DE�z#�e��+��9߷������zp_bH6�kݜis�(����GحW�u��E�ܦ"�Nͱo�kį{�r��_�$!��W�y�H���@�u�`VC��x�+������ׇ�]��i�/�O;��勫\ʨlʺ�0��q �Xѥ;�r�`�x ��v�ēL�����4�o��l�2	g@�.ɑ{Ӭk��8����E���O�d�ۻ�b$Ť@ ��9ޙ�ߝ���O��A��1Ǆ�*�3��B"
��FME1�I��[P�z��㳵>�b��DF����H�����,P�;7o����sk�ט�i��*��u«�uP�n��r�7W7%DDQ؂1��}��D8����5��B �KZ��4	4R��v�J�r(\ͼG_,u��!��̙%�}��I��uu�U��?D�;>s��?��,�6w��Ko��d��o��c��b=�!��,�� �V'�`DFߚg��SAk�Ĥ�z'zT>�<b����Ë��:�|.��kZ=�t��r̒�O��2��.���:�[ʪdF�p�Oߙ�^p�}��ҏ�ș	��a�a�Hd`�����LH'�ޙ �.S�4��X�;��(R=�0�������o8%�?�$���NKSr-�']��_]�,_�c��iT����t^h�|a�cX���R�2� o��42,d����=��	P&�M�7Ͻ�"��VMիU�d���#�lE����VŴ�Kt�Yf[�Jܸ춨�[�|*հu��������d���ZH�$�1|�`K$�݄���U��0�t��͛r/��\�_��hsD�~���bH�)��fA�N_�2e,��=��z�TuY/w�u�)9����&�Q�A&�t4���9��6�w��,�4�.�$ٯ�"��I�{A0Fd�zj�Nz��d7�1�ڵ� �솎�����^e/��gˢ����/;˴����ɺq}7=���B Qw��~Wf���Y<��ȉ��ߣ�r��))|���� 8�b��aXeHnBQA���\E1����H���
9�>S�*:���|���nI>h��$�mÅ��2q#��L�Oc�q�2�ɣෟR�eg���D�é4@��)���������73�^��g�/:� ��+�aqj����߫W���.�[_���L���ey���Gtdɰ��^I��X����"Wb�e@����H��y�5�$�)���OQ�ڊ	��]�9U:b�{$H'��)�U�6�b�L�JH����ໂa�0B�Z���5�1�J��ܞ5O���;]E���N���!���o�U��PATXч�=�!�����m\��2���[� �wc��&�֊s��e."}����0 <B*�vӹ����\t�P�v�)����	��d7���;"��|��
�|y�sO�����=E?ܬ�qё�D��� %���r�3����z�T������.���\�@w�v����<�?��j��ҋ)	 �\��N�\v�[���ʩ\�ԭ���I'�8���Ia:1��Be��~gϝu���y�RX�2�֦��M6��ͷnL��S���o�YS�j�-(\��z�VXC�3bs a��m��=����EXݡ�9U��n��s[���`��ok���k�j�#�P;�	b��۝\u�h���{)u�w�g"5�b��S��]kWepw����B4b���䦣!�Hܚ�UKHݼյ�n��S��3˖۟nu���W[�Y��ޯ���@�X�7��E6Z葌�� �m��M! ��W��k����û[0$� �g�'K�� ������H��6�;�3�^5��p��FNԂ �z:f��_�{E`H����I�ۄB��-�n�x�D2GޜƚX��]�8,[Wv��ziL!�[��1��7y�4�)�0�#t�3Ѩ�v�G]�a��k�]�r��1���$<�y����=��$��:J����H ���^"��^�Gn��� F�t�1M����*4�q���4}]�1��o_�Ni{�����&��Y]#�W�&n�5gy���p�j���F�EdR]��%V���m
���z�]�-v�y�𬗘��g�>t	mC�;6 
X�,h:���!�W�[�W�x2ɖ6�ޓ��{���ʣx��vV���A\�����.�w����������x{t�� �0/D��1�F�����?�d��>�!� ��٨����	��w� � ���u��/YD��rN��F/#��U�
�%�7f@�7�[~��|ٸ��[B��H�b�'|�@�]��v�J<Bp�]��\�a�D_h"�W3�H�2{�1�W@����9�T�w�*疙��� �ɒ!��Ǵ�I�0�"�ʣ �%�s� Iɬ�H� �����;P@��� 2	2�� ����vj��F�A{�^N��Ce���)1v���[ԯ:�b�(�[]s	P��(wr�$SF��)��t ���ٚb��֑	n��M! ����R޳~���9�cS�җ�s��Uaj��{�{ӬHM,�"�6�Mz:��$�Z�b���&w�ޜjeN���m$^��-�-cĹuQ���׈�̊���,�r��_�y��@�+C;g���z2�p����Mۆ������<k���▧�y±��E$pQ�4�nX CA��0����*����8������n��d�M���$�QF/ X��S��]��Co��Z�-*����i�D��1�RO�����Rd���ل%	<D �6��\[��z6z_vv�7O�5S8[ٱ�T�K&���S���ޯ�f1&���W���y��`�Ye�Ŷ��x�Dc�p�*�~|�߲ű�Ѽ���XN{"[̄��ހcvMܴ%�ؖu�> ﳤH꒐)n��N���P9��}U��u zN= ��oq\c:0� o'�H%��df�RO��C-��*%h ��-�qA�똖<q�C�-AS2�Ǆ��!�vF�H}�0�-� ��xH�ox�s��d̍�!���$&I�����,�F�H)�f���IMɁY5#��y�q�Ճ��B�:�ڲ�ܘ}�ۧ��+�<�u�xS��������( ��0�4�;�x2r���0rJX�Y0��F[*g�lx�"�R	yن�D�j�࿞��>��&*2dI6��D�%��%��<9z:/L~�a�BA���S\�-	n�i����l��3����ƍ�	ܕ��P�T�s�Ǐ=����ށ {���}���-�1�gj�&�"� ���p��g�. ��P
�!�5�͒��x�I��m�AxcԳ��Ex����84^�� ��
c��![��dQg�W�HȎ�D��DK<�n�y�[cL8�{�."x^�멌þ�˽��W�q�AC^\� �%N䷚��gtϲ����4�q��D�bA7���.�����xb%�y�k/Dٓnnw��A,�"�IW�U�y���f5{{1U"����q�P��2׼���BҨ�en��枞��7`�;�g�<e�� .�������B�$�3��z<��<c�ֻJ������]���z.p�c|Y�me�
yS{�x����ta��ɡxZ8� ���K��X���a��d��C�gϜ>\8]usV1M�[hk��$̺��R��ɸ�ti���v���f����˂�:��$��>[n�Ĝ�l	��֍M	�o+[-�<.
h�5l�l���{/lM��wa��y��ɣ<<�gVF��ܝ����lvxE���v�@��\.�¥$VXM��]���]�e��5�)�d�E%�g�q�V+9�mi��ZŎ�_߿��O� ~��ڏ����A���I2������ٍ�md�vNć܆��H>�p�P����깙 �W��^�>��e�-�;Q=��J�z�_E)�qZ	3y��8I��B$X��O2ûb@>gdm�-���=C ����P�ީ�G6�xu�%�<}19�7����'�vESy�vN^��p���h@��@���\n�<�຃Q�1��2@����N�9�B��@�M2j\o���K��u�����}�^)����k@5`7(c�<A�M������k�*���_��|}����~�Q^��)7F<HԹ�bY\D��VĺoG�ı�*gOѓ�A�s�i�Bֱ��e�ˬ�#��Ml{���*�{R!=�3�cC�3};�jV�R�rC��p�f�;*N&~��X���ә�s=H?B~�y/B�pnGBD@%��e���� �̗}�KH>�����C�iv���$ ϗ�,�TB�y;q��{2Ab�;�Tn'��X�6�>���AS%��.Sc]��� ��\��AL�l�D�HL{���yޑ���L�w�F�e��]�D ��r��l�4��c�,.����UL����H;ǜK�:us��y$�	@�]�V��k[�c��7%��V]9.�;�p��HƳ��ޟJ[$����|��'���֔�;z6��G�r>�J�A6C�z@�E��s�-�I"�ǎ2�����g��l��ۙ��5׏O��Aԅ�[L��=�6�@�Wk����L�$2�-#��; ���BWDN�Yh���a~�P���#͟��z�..~�o��תn
4��>}�H�=Ç����>�t�;-�eQ�)ɻ�E�z�=w��ӝ��4�K���d3T�T��z{Pc��9l�䧧�R{��~��m7��6�NyQ?Pz}��u~�W��z^��F������GN`h�2���|��c�~�e=y��C��[�f��-C�|w�>�rM�4a�=����WL&g^k囫�j�7���[�"�#����>�{o<E�;�R%���wR�o_Oy���l�? xo���k����;�,�9�Y��PLG8y#�<��ף���.?���E�ձ��?F���� ؇8���[��)�6L��3R���B�_d�|��YKg��=���~rz{������z)�m�(�9v������^�D�	�ިts@�&T�Ō�g����-zlW��!c���Ǚ����q�^��q�N��{�qg������^�-r�!��"U�!;/��.�طNB{-��gA�[�z���K�'����R��ݼ�j�����d�*#�s@$Q��%/��Ģܽ��mF�Q��g�s��{�^�W�'�w���K�毬��ɜ�qx{j�K�fs)_�����̞�3}w�<���%�\K�Q�?y��zC2����Ȍ�4�T�q#L	�!d��h��f`�속��}��i
�=G�t4VŃ*+Dc�j��˄��'����3������&�z{���n��M���y��{�cΊ�chMc���B�M��0��Ĕ���<��éml[1nb���kmmiiio7��{���%#�X�!q r+��e��� }��@N,�>��}g��]}|||~8��|:�8s�c<9�P�ǀb�Ɩ��(��^yï8p�q���}g�~������q�#9�X��˜i�|��c��U
{�P �����p��������q�믯����q̞�EYÕ�ː�Py�MkthXa|II�Ϛ���\fq��~>�������qǾ\_9ӲM��E+���+�1���82�d _��
�������?~>���>>>?q��K�N?X����'?�x$���;����!���r�a $��ǂ�l"�XO'����<�����T��(�����ˊ��`tH�	4�Y��#{ݻ.c�@�bOa�C� �YgN�c�+�W�e�����p�Z��I_k�Ʌ�FES�<@$�H��H��9�.~��������8��S���	�u4	;���,���Y@Â�˚Z�� ȍ����mmkh�^n9�O���@<���sg����TOx<������<:â���#�eE�,]�S��)^烼�{����$|�<����'w�����J/��Jg (�匢���A�i\�փt�l�����	"tvA��￑'��*���9�w�\��Ixh
϶�H�ޙjT����q���NVϑ�yby,^;`���m�"�(\t���dW��ڈqw�iɩ�T{���~�t���g][KP���<u��('��Rw�����L�2�3F�����b<}h��m�WD�rsK���o4�x�d�7B��o�>�N��p@)��Ω>nCW_����M�ǐ.�yx<��yQV1�'���ʃ�ɏ1$�zn6�g�O5��C	&��
n��U��%�D?��`��<.�
���;+��Wp���ᗽ��"i���DC�j���g[y���.�H${����ށ/w�go����ߔ��m�@�[H咶n���]�ף:[���J�UK�ة��,�����E??~��xr�;�驶�d��{) F�< w[rx�yTEk��X�Ajb�k�� �興K�r�li �zx�^�l֕~����$��Db|�u(��wB鐗3��'�(�*��q�"�({��ٖ$�쫹�P��9�k��y�}`vIܮ��(��x�n�<y���B[��/~�~V�V,��.�Ȣ�P'wb=���r�O�>Hsߓc/?U����^ĉ\��{m�I#�ߙ��.ڿE����A�6�^��=�ϋ�~�2g��m۪�uV���}S�r��Ū��y��Z�t{��	x�.����&�{n����?���s��������X�#$�&k�z��.2o���g<�|dl��X�u�����G�U��T-	|��D�G�I���,�X6��a��c�|���gE2-�f�p	Chݦk��抣f*�cL��H�����ex
͎�Y�����\�3W2�,ۊ�6�&��i`nc֑�h����B���4.c s�eKM���U�sH�i��l����.��9_j/���rך��J�[1�l�X׃Z��شrm�}rҸѼ	uv��J��.v뙶��ر@�c�ImQ�p��~_���K�W��5��X��	�\4�Iż�4�S^Xe��O�DOt�c,v�"�	A,���0���g6�����|��2�DL�=�HvH�c�;)bY��1F:�ד>����� #�y�'�e��z%��~Ɏ#G9KJ,}[U]]1�P��ǲI4���xb!��WZ�Z}�t����:�O���3�6��k�DR�&��H�Qz��IhHj�C�4���Q�|�/�f�kwP�l��D k�u�.�t���c=�@�r>����e�Q��0�u���?9����LM����ʕ�2���[�z�qY'Jkn�Vݰ,N0��G��>c2�S�^��A��w����Sj��[ޣ��B#E�v�i������d"T��f��|���v��<mŢ%_�Q�C�;+2�Q��`�A ����������S�n�o��I �o^�ב�m���c�Ϋ���Y���Ha.����42@�Yɼ�+~���w7z:�y�^Cwp����.#�oX� ����M��u�~��3�M��RH�F��X�&X�(Q�z�l�Wj�d�ܠ	뼐$�A=ܛK�u�tW
���P5�O�Ӵ'P���Ŧwc�������Kk7�Jd�P������w@��=�!{l8Ff�rL ��
������}x�x��:�`�2m�ݪX�N�aM�~�K������~Rr���:����w$.�3c�]��=8�<��U1�-�fX�TI ���-N���H�7\�� �7��FȤ���/���Z�|���")���~����=�J	os�d���z�X��H:�<A"@ڬ�z@�y��}��XR��+�ȫϨ���� ��+�D'��1S�<3"�Qv�tzyמ��kkG�x�@�]Db#TT��<Hn ���`�9��$}�~}z�A��%�<��n�M��l:0�q^o���pa^�p	 �{�|�"[��#�ܯ;S�I���|��񚽉�k�q�+�@�]v��\x���2]���	������+�N�~wg�>�����;�Z��:ܱZ��f3m"Ж�ś8����27i��8�����kh~|��?�f�Ww� ��8��I<��ie�-D��7Ay�� l��O��$̆��w�D���< |�c�<�T�j��ս	�9w9�$%܀�S>�H��4��Ciy�����	[���z�.N���n����A,5��|d�Ms�����8�Sc�Y�"��˻Y�!�H3��4��9P�C�`v�ʯa̕��>��d�tDH'U�@$����)#М�t��?�-1����Gu{�ax�#�����{�y{}/�ue=���쩽~���������Ü��?�a���@��_�|l�yчx�U�`�yA�}�'5te0�z��L2ƾ~4H9�p��9�
�z)H�V%</{eˣ�p�~�xۮz�XRk�6��X���ˣ�*A�DmYbFi[��61s�~G���P'��~�T���D�Of�Ɇ���ng��MxX#h�[�#[ɲ�[!>z�wp����v���>�wT�d���*zfd;���Ap<	��t��>b<��>=NCc��+��K�'����Vņ��
����ZE�6�t�$).��e$���
h�E �Y��^	0���[ݷR|0�Զ�<�rr�H$�v��ѽ�sO
И�|{�)�J_��0�)�7]�V�@[$5r胹YQ�/W����>�yZȉ ��KHtI�ɵ�y���0E'E��=������ط��~���Їc'�;f�w,���QŴm#w{��r~}�-|����W�2�7[�H�����#�:�$gx�5U@��� ��N6�l�$�D��ͻ7�wyg��x����ܟ��xX߸�Q`��4�<x����vYKu�Ƈ�^�t��Ѓ���$�@��zlh�Z.�v6�M*rf�� L륱��c�K���8�������V�٣X궋6��p:��+�^���/;n]�fW�n��q�K.��1��ю�����$�7v��{�A�A<8Z0��rX��Ӓf�9�ŧ\N�LZ^l�U�t������RZ�X��`��q��
�%�s�ptT<�cwǥT"I�܉��������O�Օ��~eLH>��<	/��<TAxK��� ����*M��`A�\�fO2	����2�����Q&��轤�	�'r�+=ޞ'q�ʼxb�q��WVݻ�ݝ4ŷ{#�Pon]�_̞"R.��Y]^�py����z����w$[وL��ܟ"<rW�p��:N="��:���ވUL��g�:m�[���XDv��I$��֖R��:��]P�=�^�.i���F4oFV���i���LG>�5��>�4�ޥ���T̰C=�~@��O������ �]������������E�?�@~����P�
ZI9��B�K�%���ܗ��V��[P�?���<:7����>���|���	���JA�N�.\3W���`<C<>y��Od;�~��7��:�a�� 9	�>?�>�d�<�m%����~^�@�ѹ�/�o�Gev�\�>󾶣�UBut�m�1�p���kV�/�vtFuUbiD����Ŵ�(&*ד�r�~����	�'r�rTl�fwQ-�μm�R�~��|�&��� yd6;խԖφ��g8H����uD�N�*{Sa,D�\I�Õ�yjFͨ��hո��"ݝӍAt��=��?�_����5�]i��k.Z݋�wU�WU��M����[��UL��kW!Ӷ)��{�p�:PKw3ҹh�$>����d����kG��7Eh�M2ǽB{=��t]��P�s�,E2zt!O�Ȋ�����7��@$��ސ$��
��U��/�D���`.<�W����)�u�D��E_*�a�:��U"¿6�8���rE��K+�:����|��t�hx�u�A�^8{�w��n*���,� �$V�P_#0�C�/�Ì{���0�W�����F=�ꁈ�ʂAk��&fz�'*����gv��b���'��&�ra�-�Lx������̹��c�y_���2��(���@s�ƀOy��O��_��!,g�)��ĉ^�e��{�2	�[=����|��N��EYA�ɇ��Zuv�+Ǟ$q��r�����U��,t05�������N�.�t9�ݸ��2�v��)p�����h^�{s�$��R ��Z�����-Q 㚪ܹk�̗�A�tݜ�1����=�e�T�/Ш�m�o0���!csf5�\� Kc?1;��+e-�{hwe��x`չ�Aͽ�'yܿD@�l�J���� �8�N��n�<E�a��?�	d�Y׆ ���{�L�| Ϊ�r5�xzd{*^���G�ݾXy��wH�|P�����W��H�aָ��mC�C`ޣ
�V��sx�">Y�	���X�R"��>hjg�쏍7���'J	���x��Q0���A���1���L��fIbOo8�t�(��uotu�r@��肹���&���bs�뎤�N�2�X�v�1��ks��'����ejЉ���}��Q�w�S+ K�r�^���F���WN5)b�3$�L�zI�y����!����Jwz'_k"�$�~؂N��	���Y�Ӻ�p���V�7b��w.X��g��$���-�i���v!b�/�}߱�I��ye���}��<fpԾJo6���ׂ$yU�c�׻���#�{O���M�Ή�Ȍ��\(�%��J��K�}[�.�G���hgz��� x�+���楀��0���~.�mFC���	�L�Z���/�x|Ϸ��vnwT/��}x���ܔ���yuBs���{��'�K��{]��:|F Z��ù���ͭcAz�n�wv��v�ɷ�>�S��*Ŝش�m�83;�����H{T�tPq����B5����y��Nr������ug�l��^��&l&��\?~g<�j�W�JN���v��Q���;�?
L<�0�8��[�p��=��G7���=��r�o��{q�"�F�d4��T����n���>�[���I��Ka�i�F#����c��ȕX���s��|\�L��yh�/M��CݩdU#�X;����F��I.��B��w�f����5����&w�}(�^��j=�}�O�+�ǻҧ�ɔg1��\EA睦�G��ru�����Hʛy�=t��=��>�7�{Պ�|R��K�9*)�J�>Ջ���c�����6��g��|F�<�������)���CB�J=�J���g�{ڋ�G�g�X�D�C�N��������i���u>^}�<�6,P���j���E���՜~ȟZb��M[d��y�ӼB���˝�<�<���#��q� y��Z$ك	���7J�o���z����.D��@�q>�uQ�wU�VN9c�D
aΐD�;��b�/kЎ0���(`�R��T"y��yy��������l�`QR�x�k8�&��ՓN�`��䦑�����҉!|w�"[S�`��S�Jo� 1�U��!j_R�r|��N�,�Y�aу|"��_S����,
��uh�-؜<�K��ܨ �K^�"�����9i�I�
�%�"8
�V���<�WKw�}��>�.1��+���_��n�I<�[��>&��)�����&����jz�K���m�v���",��:�x4�N%,Ev���=mMm��q�96��r��B��V�£SA}^�}�������X�1*Lk��~�9W��Oѫ��D��mC�Q��*@	�Ǳ��$������0�<��gs���__�8��ƞ���9G�X�[@�+bG��Mz�tƃ!M��"��ָ���}}g~:�������q�2�9���+ ���L�ųu8����=V%�����\�n���]�}o�ξ��:믯�����|ʐ�\�k�'�E��φ���I�4�@!�'��-� �;Y�������ooon>>�~g$ˠ�ZĖ�>�Ϣh33��7DugGY�ð�*���}}fq����]{{{{q������r��s. �RZ:�?/�D�,<m���UU�9�����}g���{v�۷{�{�}�"B �"Ϯ�8ӕ�R��ٻ$+ζ��,�MP��)<���m<8��\�A�jV#6+l��lD;Vx`��Y	�;/fb6��1���N���#�a�����BQ���� d �H5�46 ��5�hDg��l����C�@�fж&i��e�Mӭ�6�C�9�����ރ��U�n�z�r�`�^�u�n�α���;yy�OQ�gvrR��Ѫ^cb�w[�����#%���$�����^���kmu�\�el�5�X�dΥ�N�����v�.-�glǵ�r����4�WBLa�,ĩ�b�&#v�1���n�]׶(�E�%�L�(�"�2��>�&6�� ���qL�B�t[mɆ)Y��Fb#u�;m%.�ɝ�������ЫZ�����(��-��Iwg�;��9��K���ܼ���WYaEч��D �vp�f�չތ�o$<x�mI�P:�9�K��-�8;Z�C�����Q�:b,kW��N��#�YҎc�ց�e������Ņ̣l���7*��3F��9n���$r�MM�J���7%ۧD�����q�z��.nܦu41�y7��}\���FW��Z�n���<�jM�%������9��a����h�ͩ;z�mϰ�g�d�{���ӳ��LS�faLt�qvX8݁�l��\#�t�X�=Q���g�����1&���MmXʁ-�y)�;Nv�vV�a��X��s.��{����9$�q�4�Td˩66-R�L�+�#�n��q� ���������)c�))�2��Euf����5��큛�9�,���*��Zm�GE�3�p
�f1mm{Z�í��.�5vѸlѝj�t�ڎ����S�n��0s�8�\:���g���4��Myz�Ol��79Visfrl�	*���Ȅ��A6d.��?���g0�$��5�΅[ѣ�r�� XGGJ�^��dKlrg�� ��z��]�y�Y�TC�E��nޯnt��n�K4W�[ ��X�YfìX�fu�J�y�;��(��}��[����R�4��v�z�J�mѻ�����q��*��}�=�n~K�i�;]Q=�<��'����wv��ő�L���F;�3�[9�r��=�9�f�=�<1�zV��kb+=�%{��ND9���� ��h�2�p���v��!�0�{��ű
�ڂF׉E,˽	�,z�l���;��
᠂I�g3��'�����X3�z��*Ul����	<A#���!�΋�H;>4%�:u<W�lgrG+� �;.g�����I�	I��B9�ם��okeG.\C[;���X� �xX�Ǆ�4|}(k��r��9�r�B����%��.W Gzcj�h|�@�ڡ�1�݊$��p"^f�+F�uy7ܜ�ߤ��,M��@]��F9�\v�ɹZ�NQٵ�,�TWKHF������5�GlQ<�'6�Hv�q��X�y���zT	��S��jx�"�@T0�"�ہ�'kOz(��z�� ��ggwyY���t}uT4��'ov��4'=�뽲��{*�r���/��b�g6Fu��"3�	Ĕ�Èu�>����s;���i�H�����:�b�����uZB 8R=�i=s�J�� tS,bbw���N�ݼYVg)$�ι�%�9�m"H��D�!èg����tDw�����;ՑD%�놃�5�s����h�}�1�e��v�Ăv�|�߃�xF���$x�C���	�flܱ�@�\ɖAw�3�ɵw)��ޢwQ�Pd���#�(E��+��sDF�x��ܻ<vuq�rbP;N�W#�ff��;Ð���R��9v��q$��1��1b꣫ީ%�=�;vx��������ܦ����æ��^��6�{��mgyd����A��D2���&���:��{�a�4B����&�l8���Uʪ�ȑ~�xv	7q,���Z�����œ'��6m[�SU�XY-���o<T���]3=׏qE+�t���~����8pd:�b� �^�|'/@�K����dV���\*�h����5��ɂH'���_wR��x+��Kn�֭��ć����ykb�Au�D���Ҽ1n����]6��(�E+�2�f�P6�%^�]��D �'.��9r�3ts�vvsm��]��K F���rJ2��	�����w���!���7��e�3�>��}�^��c�㻠�ۈcF��K$�#H'7z�wO�`ڜ���팀�;�L]@�W�ܫx$�/b�J�J{��M4����-�\��5v��^D(���ll�C�B��C`Z;�#|�����i!Y�SL�$*�'2kJca�U�|z��뺧�Y�H;(=�r�ލjH;�7=��\϶�?��L��9e��p'��>�;tтY�p��i�9s�u
e��`��9���ם9��NO��A����	�`y��Ώ���(�{'���.�m��O��/ޚ�T�K�s-o-�%��n�ݼ�O��{�V��O��ݑ��"G����~SPuZyJn�$w˾rި��p���_jwm�
g���ÉC?��&��K@]� �o80|���ȴz�쌞b�$�����wȅ�DH��y�n�U�'=�)�Y�n��8ԉ"�u��Sw�yVw�8U﮷ah%4O{ ��N��{�}]T(d*�`	2�N�rb�@2b˷:(�7�fx�PbDU���f���De�WE@�4	n�1v29o+��{�6�H-M�W4*A'=��!�Y@�ب��]�.Ew�ϵ���zd�I�d
������ݎ�O��ެI��z�jQk*��={�~����_I��w��矚YV�vw���{�@����ċ���,���y������}��U�k�������[ZUI[��Ͷ7f��0��?���!9'+9����,�����������;M�nG��9�G�	b陝�&T����p������J��&�&n��q�Y�6��i�g�S��ƣ�=6]��G��n��%�՚UH6c�;3%��'k��� �ܜR�����S�]�����r�K��VBW#�[dpF�ipmv�f`�r��L��o-	nVm,��j�Վ9��X���Q�������0^p�pF�M9 ��/gH�d�Κ�q�R|��Gp�=;�e�̦H���Akn�y��$�3Ȼ��.��N6\��$�rIÎ���t��o3�E����\z�U��^Cy��E�9�+��S��)��"Dzy����%���&..A����[T�zԒ3��J5���:x�
��~���\�V�l�f�O_��;:6�Ր��/:��sqܗp� y����=��:�!)	�^$�z�LS��H��k?d@�H2��P|�I%���k��{�6gS�і��pm�*ڵ*MԪ�<��9�f�D�30�*8�vt�2((	__` �B��>�~$�݇���v��a.�+�~#i�^LC��PfA.��D�x���F�����>x
�X'��-�����x����f@ߛ�w�)�̻;�L�ͽ�y�8w5��}�%��G�
SR�D�Ȑ~P�!��NMpy�+�Oo�.����e����$O�t����O���i�A��KW���;���@4�m�D�N��]�yڏfA��]��Dg��H���I:�%��?�c�O��25!�
�$�>;
'��|ɂ'{����MY�b%?(8�_��
���B��@+0;E�Uc$��ܬ��h�(�@^��l��	v1�;�&o+��E�BD����h�C�[����a-(�U�n޹�x+��MVZ���>�GJ붿ߏ���[vnω��kΈ��p+�d^v��gOJH �r=��$�$���H��+
��8Lp笿d�n�8>�4k�E1vAS ��>��]��R��A��6�0�8^�ڊm�΋���d��_���r�
�t��}�GH�7�PJ����/�4y�������y{���ꇘʚ�_����-C�o�`C2C$7�p`�����9�ǜ��x$bȮ�"@��7�\�y�}-kǺ������S&
�$�	'�A�>gw�]>�{�wp�_�@�SO�O�/�:�]�@_���$�ˎl����ٙ��";+'��2
[����<H��P��ݚlY������j�T�6̱���YtT+�M�K��˺��R�1X4~�I�RJ��˛�ۣ�o3��Z�$@ü��e���]5=I'�ȏ	2�V��DB�k�T��M ˶|�U\;$����=�ȵ8��TF�w��́@W%� �Q��I6��1|�i�	>>��H�W/����9�*�<�!�y@�r���T<9pe�ݵs��O41@���x�($�}�7
�뽾w�^���yWg�/�q���d���Cgp��s_�ZaaD7���/��܀�k{ǅ�>���;.s�~�a�����0�C�	1�p��޿��s���G[^���#�n���B6� -�bF2��M^�D�FA2���Z���9߶�>���^�n���4��;Hܗ�j��aަ��]�v�#`ncrIs�[6���BGp�e�]��z2 �L�Zڢ���AS$WGL�׽�Tnc��C!��̑Gܠ-���A�� ������.�ޝ%���o���׹�}�2E�ξ�W���y�ikA$�g,!B��x�B�uĎd����4�g8 �'UʂA4ɷw��|� �ۗ�� DJ�`�9�ॳȅ4cVy�cc@�|��2]�1 ���7��M�LI>7�H+X�Y*4�xe���x�^evU
Hq�:D�ߧwx���֪TIk��vO�1o���O"�\ȓҽ`��>���[ʙ���uؽ��h愭S��X��p�#1n�r��y��p�ެ�0>&h3�֫�),!c&�E~��L�B&�^�K���Jƺ��%�l��M��w��I�1�81���˃,=�G]G���#>|C[cnX
���[MXYF^�і��\9���n��g��gc�gq�n�m[Z����Ը�"�s�ŜHUt�u�udy���ȁ��CZ�S�-n��4�Lq���TXչ�� ]��g�8�4���l[Ĺ���Ґ�hP"��F^���t���m��S��u]�Y.��t��a��3cD��bl*(�3߼�߀"%���i���Ñ[s<�';��O�}�O��Y(�n�铍s'�(	��/�팽�G����u�.A-)
��v���{� 4���%����$A���B��A��O��	zk�>�������t�&�y�������3֠�9�2� �9ހ �A)٘pD@���0ቌ/k&4�)�ff��/�%�"� ;;�a�Ǣ"�k]����ڷf�D�I����b��x�}����?4+05�e��R5.�f�K]�ò3����[~���>���\�3n(�Eїj�P0K�X覚��GKt���J�cY��^zU� y���9�߱�nw+:�Dr��u��Z��)�A�'� ��5�/�#�b,}B��._�Q�Oޏ#�,�B��X������y�{n=\_/�+���K���=��^��w�����u��q1زZ��%���&&b�j?�ņ��	c�����s�$���D�Fs�a��Z~�w[�c�$#A%�ʣ�p�A� �v X;<��W�C��1op�x&��h�$� N����Aڽ���!D<��c�}:�=^蚹.l6���w>� �wF4`�b��8%�w�U% R�g�a�<A��t�(b@ v�D��NTz�DC[��k�D; �.�g����a�y��)�S�~o߯��i����Z��f��!�3+H��k\-Lۥ4�R�Z#���x������U(Ӌ�?z��$���e9)��Wus����VJ�����V���$��B���tT�,�������7f���	mU� >d�����)��W�w�a�+�F�H���i!�xexd��>3�ƀ�u�%�(��ɧ���<9���94�x5��/�b؟�ХٶAk~�rk=�맧	�K���ΏK/�y�����M�(W��Ȇ�{c���vﻕ���x8��~��گm�5v�r�����=���K���ԳP,,X�M��*����nm�B��� ���M��q��6�G��@���t��Ǝo%�c�0gh]��Y]��AᤍK|����/T [���n��F��N�ˀ�G������s~�OS�vyV��Y��+ʷ�)��.F��M`���p�<�Ff��}�p�nS_m�ND��5�3�]��3.m�G�/x*�������g<��W.C}ty{�3{��tM&�Ǟ����Gj\��}��\��[�A��-�~�k@�4�)�r<��;}�l��p�b�[<<����J��p�kb�Pw��q�c�@�Eƅ���]��n(������=��.����{=� pr�m!�������&������y]}�{�U��2�v�^����&�̼�!��m������|��st�n��]a%��B����%�k}�4���g��{���wb�R�m��0�N��;5�x��޳�?�ܳaB��,ÍR\};̻q�ϵ|E�ู)q�I�͛m�
x�:tvՔ�#�5��y��X��1FTc`���!D6���i��:~�3uj'���/���@�.r�C��z���"��ͤb��P��uT�炄��t��	�{�Y���H�>���V@H�!�}#W� HH��l#��~�>����㮽���������3����=������Ԫ�9�H�clz�oc��;�~q�}�g���>ϲ�˗.s&뭑6Ƈ�3��d�y�7J� (�Fb��^�t��D�@$!	Uz�>��:������������ǝ�x>#W�	�*� C.'�c�$#����o0	��tt���~>�>�G���������ی�P&0I@�lL�`  &(��b��[{�}���g_G_���������捄VqH���eT
��� ��B3.y:~�
)�Դ\O�m�B;�Y�w3��g3��}ｻv�۽��<�C��# 	�E�x=��%�0��)��� p ��	H�U� @�V<��.�<�!��8#l��k�H �-z{Z@�1
��XD�F$#<m%�4 V�<� $;EU��jS�Ą!�wI� N��wmԇLH�h0Q"vPD��ĐͰxXC��Z?�44?�s�C�GI<��:n}�r���%���F؎O�&E�}�{��������ڱ��I��<��.�a����55��ܯV2�����"	Yus �N]����A�N���~Y� �J~{�v2H;��O�Cת�J@�)%Kb�o�ô]v�X�C;�\u��n_>��:�C�s��%c_����W-7��.�=�b̠PJ�g��b(s%�	�����vs,�+�E�K^vM5��xK� �񽣘� ��u���rkt��os%u��Y�ov�5�8�5�tϲ�l>۫c+��r�v��䜿w�dI��h.��o����ˣ�.Ajܴ�x�{÷+��b�<o]56�������.	�_@��&��nmωNI9�� ����SV#�
Fy��\�Tze^�葹�G|+��*6�^N���t��ݴ��������N�כ����f��/`�\��̋7 캧�V���z����zʻ� �@�^����R���kbgP˱�d�e_�a1@��0c.���{u�?�f�I"k����󪝷�sGV�p�|)�q�u]�g�nxf@�ڡ%B���'�%��W����{�|X��Ȃ1�Z��+����׎ő��c�~��G|��겖Wm}]�٧��Wx�z�[=�NZ�"m�� @�J�.���e�~����N�X���J�e�b���<����.�����[43PX�)��C�^�t��C��Rf�ޚ3�l�'�$�ݓ��x�u��6�Y�OyY�I1-ݽ%�^���h)��y���SS[9/�W�3˹�90}s�V���ش��C*���a��ɢ.	݉�|"X�]�2Uٛ%m�rt�����.�������tn6ǹYjY��ox�Q4=d%W��~�Oҙ��V�^	���?`����)��D��r��D!Z��(y-����E�v-L5�æ���m3a�|�gF�k�5x������kK�K7i`�Y>z���_����7:�;�����y��'#4��w]M*��Ǯ��)Č�ГPst�W��k{\ѱ�gYݕ���4� jJ��psX����LsQ�8y}DG��M�z�V��qn9wcۃBm��Y��W�fpF+C�۰���p6ľ�zn�[��x�}�^9������&�W��0!�5��V��S,E�W��:H<�	rE}l��b��~j��DvwU1��:�u��߭�Aݿ�j�V��" ����t�T��D��7{Û^�`H�|�Zԇlt���'z�W&�=�֦�7��4��	�ٖ�z�A'3�8�Ϯ"9 ��'Q��7ˌZ�K�ޏ[%���V�f�"6�Y�;��+� 5��& �+.Ј'ٝ)�� �xN%},�9��ɗ~0LϬ���9p�w�(�Q�M���W"K��������<�6�<�$[�̐N�@�{�zK�`!�TD*��Sw���:'^��9�K5�b�K�����?BH����p���5�a\��o<�O~��^�x�v{P�>�6��u[�ȵ̑l�肉���Mq���ę�T%�ÎO{}��-i���٧�xY���:s����N�nl�9�\cGh��F�M�;��y�Q�<ڎ8.x0�@D�@�X�j 4���
؝$�r�M�&���ZA خ��Dy��,�O�wd���_Y(��E�f;fA�q�ᥒ5�
r�|m�� �/dH sz��s�l�ͣ~����_�����&N� ����� ���d�2�p9?�[�*�f'� �g7�x�@��?�&;���t �d-���z���L�ϐ�	�\`es���2��I:D$yP��g>��ݫ�:3�k؜��Otk�/�����JC��=��L�+:es yq�q��y�r�����j2X[R%f��$^�H�r^H��t2�A.�}�R���ܨ�O$K+�i�Im�� ����Dfd��ή�R���H7TI��H����,a���!�*��o��GL%���8s�/�,��ё�|����Hԓ,Ԏ���~-��[�Wom�/awc79�%��2+Ғ�A��2!�	!����%����6tq*i[�%��7�*c��3�n��UlAme,]�Ϧ����1X&�Y��MMKl��	�CZ�U�ِ5����4������S��G��K�V�7�(��Tr������wW��%Q��n[$�і�0y�qι�[4�]S��q�m��:�c�߻�*�A���m�5�d��ZZ�]�+oY�zں7H��9塤�-��_���46߇���B� ����gXaܥἺ��T%���q�S$D�t�2M+}sDk��4G�I(�	�a�'�(A]�'���m��gAg$=D�v[�?b�I+��H���O�:�#޶]��>׭�K:��	��OP	����T��4<h]�����O�]�������[�>%�U�R�<ef�=_�>��o��|�1>����|k0�X\M�A���p�E�f� pbC��bb;b򸌎V�Q�͇��cG�߻�wu��kė����f�;=�Z4����Ӄ�X8<~z��1<pT��׊�k(jy���\a�\������{4��	��@9
y�2�ƥ�Y�D-Wz��s��gl�R|�
P���@$z�'wwX� �N�X\���-	��}�u�؜�R�s#dCi]�i�{6�L��a~��a��P��C��W��>����$�x�w� Ke�u��2	>d��"gux�� �z�:����L{!6���a$�����@���`���@zΚcB�����&��]ػ`\v��/
s�D�ûI���d-� ��=�\�;�r�y�s.����,/�A���M���u��@'�w}}���f���a�o�+���AmPӑ0!lL��j� 9��]��o��)��D��uw��������K/�W[�;'e�� mK^`�ь 0'����)I&�?�=Xn5�o.s$	�ܑI-�;�WXH#��K2j��׵eb��Y9�Ӈͫz�`���1�ٵ�^�M�m�{s��`��fs�t�j����݋��l�A�r\O:��kbf6k�%��#��8.�[ù�{�5r�!a	������-�64���:y7�\��%\9xܫ���Az�^��q5v�r�;��,gh�Y��t�3��n�}��D"���9� �K�����F.��0Л�wd���9�%�{&Z��#yj��$�����j��m�;�՜��{SlH�A>Dc!�r�2�^͊���1,��
D�{v�`8��;�םh�(��r�Y+׮��xA��v��Cs8{~���'bYc�)>l�
�S�p�
�wz���*�ėx�M�I̘�L��v��|+����}O��^�,1�QŹ�K��D�g0�I�sa�Wi W4�j�ڊ5M:�i�Gn����C�=���t��<_���U��hG$QEi�ߘlC��B�2�8,�u�����7�U��?��!9Bl��qز8r�A#{�KK)^��e:��s��a�|������P2MQ��B0�����$��@ev޹Hk��;���^��Ti�3������ت^ 5���U'���</���	�*��=�뀆�ep3�y&=�؏?f`a�0�ݤ�H%��֨s��:Ӕ&�=���=�I�7N����T=2�Lv���i�3�^�e�F��sx��R�M#�x��9�6	0@���k.���p����8ָ��d���)S&��ɐ�:�{Z�bhy�,cA=��)�C��^��~�T�@�?>4�k�:ؗV[o/bH�^L52�3�#���}>�pL�4�i�ϣslN�p�3pn�tx�Qn����k=�MR&ʊjȎ��D/�J�=_��A�AScGdM753�c)/8�� �FE�L�s8C��PI�s�VH5#�G'd��2�l�bUf9�;�4 �0m�xq̔�m�ؠI �dE1F�X�[;*��RD��S,���j��D<DB/�ޘa�7����I�[���}~ݎAL���O}Jr��z����g�~��^��K�w��w���8`��u���8;a��ݸ�6��� 9���� �-��b�VH$]�Hb�o;�NQ$���8!ʈt�p�_��rs=�yr��[�u�'� J�c$�-�.��7�zv$�f�.链wg80'LF�i�>90�;fo,pM�L�At��b����6/g��'ў�����o6Q�٣��K6�*lA$��Ú��n�;2�u5fEB%�&��q)�s��rvD�䗶 G�#k/ _!Fv=V0Ǻ�@$�[��\��8#�%	[��7�6MM�ꋉˉI_DMl\��P��~&��!gXК.�d1@��"�[.}�0�9h@4�կ]�ot4�2w�8�ż�C$��uc�0^!��v;�R��'2�KR%�͈h$�Աט��3z&�鞍5�ޛ^y���
�K�J�:�����Ҧi�(�ܲ��_\���H�;9��k'�JE�r��J�>���#N�၆,���l���,�Ó���G�~�{X�K��.���:%��[�}�x�V��-29�'؄j���飑��°V��ߢ7�;v����d�N��]���vLHt�션�6sXX���fl/�~���?̯��K�Eo�ot ��R[Zc����(H��oz��I�(F!�ޮ���1:vk.O��D7�8'|�`b�ޙ�#�qxM��~V�����H"o[�1��0�a�\`����$^�C�:��y��/G[��>b�da9�0m?���}�~��W�[{H�+�D2z](�V��vg�H*�������XEJ��CUj��`�C�N[��w�A�;��W�ˤ"@�c:��c�}ƑdtB ��G!�7�(�/�cM/�k{��'%�}�R3�C}=��63�{%��/i�rf�k�#7��>��>���wnW<_A�Qz�n�Q;�<UO�lv�θ�fr�<rw��K��3E�Gq�7炇Z�w�K3����/w�yvC=_ �����k�w<8����;Lj���M�VS1d��`�������K�ƫ�NNj?�����,�r���#]ިc'-�'�sl�u�w��
V�n/PwN�޷W�&2������6�gPCk���d���nx��#�>{���n����/5�+G]�[�z�w�f��[�sx������ɞ���R�oj�l�{����T�x��Ճ����mf�yA[;�O�{��m�+X0�|.�k����"^%,�qY����wQ���m�P�����](�w�4[���#�٫7��	��w(��_PO`}9�Y�W�3���'r�v��Ei��3����U�-y}8g]zwl��t.>���}�d.�{�g׳ß!�|�m��bx�K'�{�m�=�+��q���12m״R��b�s��{��,B$����`�Þ�@(܉uJ�8��{ou���,�~�� ~p���oM��a��������r(уHغrez�J.��]���x��ܹ�83ڃ|R����Ӵd�c3}������ǡx~۽�Ӱ�\���*�aol2-�y���MWNE���CB��J�s`�+<;K�����|�|m[��ុ�S�g��lgn�;@�ᛌ7���w��'�3<`�h/,���{�틏k�VA���
�"�d����S����oz��@�w14MÈ���V2ayg{��3�0qa�YS�Yˀ��!�c����E�UH'��]\���@��}�y�	l�z\��@���LO�ioh�Z��`{VG�����Ic�7'[����88�"װ�f�5�m�\{v��l�Q��{��y�w��N��Y�A c"��
�����>Y!\�Q�jӑ�����OwmSx%W/m�i|'�>�atO	`@8�w�2�JW��u�a �r���΀.㾸����?���~>���r�˗9�noZb�'�.���dI��`f0`3�S�i���\��}_Y�����������r*��ֈ2�  0 F�P�YxTo�Չ�y"��BN��Q]��]>�_G��3���~�__r�˗.J�C@�A�A��a�b��|:08HU%��X���U]�<~����=>���������۹۸9֖ ���L�zG�}�P����9��ӧ)�2�������Zرgm�����oooo}�MU�O
b
"b��"H�"�BC��$�!�ʙ�A�7��|���2g���]}{{{{{z��<@����XU��<�!��ց<���� ��V)01��	F<*��Q!dYf�!�pg�� �!�@����;��]|�A%�2^粘��<�)��}�(��
��x�@(��&<�(�g���!	���-�o�Gg�p%
�ح���2n�Z淦v[�8�&�id��]Z5�˗g0�AY]7��]dE��kv��b��a�t��̲�&��65[��-�t�p��6)���Ƿk���]�k,�)�%���h�hDۗV�Dai5��:wJmnzҐ��6�Y�C�p����4Xxc�n�\q��6Q���٪7h��X	��+���r�JʹRI�izv��Ň�V�#5��l˦K�q(\V���v�z]s�'hv�7=I�1qr���Q���<��Lp�k�������!�`��(�k]M�a�b�Z�e�1ɟ%e���tW3��ۥ��ev�9^�܅pV�k��vn���+J۶�E�J�[R7JԔ5�8�9r��6����u#�v��A,S���Ū]�Yq��&�z��;�ѺN]�Q�r��;�Tc7%��8vlWn���:�msZǜL�g���R3V5W��񱦱�֒�U۱��r$�۪-��%rs��/��1��r�7=ͻ1���.|�:�\v燃Y�n�ka`�1���de���IH ����14�Xan��V0�D�J:4u
hdWF��y7��v�[[�z���2&�1V�}�i���g>)D���;
�tZ�Ob��7 s]
��wSݮ�K`����j�EfF: �y��%��&�6��TIWl�$�V�سˁ�9꺚εth�X�5V���I��C]	t���nk��3�ݘ6`��\��*�+=.��Ƃ��z73�%+�u֮��Ơ��q�F��M�n^�ኻ5�pv���9��㢵.O�A`��z�s[��X��k�K��hCV���]u&�	-R��9��m�l޼w��������^���q��}ɴ���;��J���]��cy�y�\A�Q�5���,�@j:b7f1�.��冫��nt	���yC��c���� ��N9���k#�3^L�h.\ݛW�I^1�z�~g��)g�[� j�ۍ���z.Vay뎰�^��s��t��Jd-�}}$�[�3�z���ݨ�ML�c�m2JG���V��j,;B9F��l���Cq:��H$V��	c̒�k�M�BA\v��G�hp{.��B�b�2��X�$;-�ȀJ��x�>�(Q�Ή�HV�o���g0�%�<�f��wk�4�RЗm���KY+͙�%��}��G�tG�k$F�u�;@���:�lJ��ہ�z��Hu3>��>$���	�\@$�n��&.:��Loy����p�qű4�g:��pu��F�5ځ�,�Z3h��i���v�n�I����\j[*sV��֮8�@�ݙi$�����ϲ��=��\���]	�W �L�`��D9J}������ݩ����C�r=�C����_kK�W�²�����:D6=�O^5�s ��"n�f"%Q���!���K`%���Ϳ��q��-�Nط���@�\�+ݲ��{�%��$B(��` Ãz����4���g%�2����&Ưw���IbN�;�����$/��
ͻ<�B�b<ީx�5���u�V���k���C䂜v�N��L���u�����A*�k90!,�d�C�@�}�h�{�;]֛�q��5�$j�(�d�ս<��y�E����#O���vE���-ս7�S��\ڣ������K3����c*�����y��W"u��� �n�1�A��v�T���j��{q�U��!��ܹ���l;�x���ͺ+=�!2@���]��>�űD�@A�C�뷹�I>YT!r�ڜ�s ��]����TC�{�1X��܉'T�[Y1\+TGg[�M���<�F�w��|w�)��0��*�b����e�
p�!�to�\V�-���y��=����4443��ǽq��ڀa�bٽ�X�v���pLYA���]o+�t�%� �ܹ�u�GWA~�Y=�,��g���n�sN�A1T^_�k��f�vZ3�$B|�L(�o5{d��r�-�N��<~~A������	Ŭ���jh]�����ۮ�̽y�gb�p�4�j�5~������5��[yf&�>�tILGw<�e��NQ���R�q�Dcgv��mT���5P���]ez}�!m�y6�j��`@=�q%2T�{��ћ���,����ribm<+�$�Hn|H�現8G�����;Qڄ�#Y.ޙmjz-؍��!üD;�6`<kޞ��*��y�ȃ{7�"/p��Kb�E`^�����EaӜ��}=�����o;��[K>�F��Tl�������9:����v���{�����8{ggu�!S�hB�އ��R#=}u@�l0̾���c!P�m Ig�A,����Ի� bd�^fz�R@����܆vz�ا�۸D ���m��}Vd�yjV��Xc�tm�Kl�;m:%�"�!�U޳��t����=��2(t�<]�?rɦk�-�Z���m�m�ʪ$�n&$`!��rN�$�23�1׷}������3-t΅�Dl��)�{2�E����^���ofA�!�9/$x
b���p%���Sg}��-w�sc��"�$r�('Z�����<C�O��m�]O����m�Á�9qZP�w4ܧP���Қ�n���5��H0����	�7�e��i)�؊� ���b��B�/O�Chk��K�Q�|���@�}� I�=e�;��8l���N\	�[>L��ܓ���Y���çp[���>�
���݇�>;��V �K	x��9�����s8h���,�;�$���!m�
!;IKL	*�bכ����BKТy����]8Sk���ui�k".�KS6P0v+�h��p�!3H��:;vӎ�F㋌�R�Y��ļ9��-�]Ye�YQ��M!�2�tr��2͵��fE�
ī����vɒ̈́n�X,����g���Fx"��Ųe�X�F��5�T���1K�)�۵��<IٸgTr���:ړSn�ƣ��=�d��rҪoQ�m�r �B�(��o;���T$Q�(V�	��$��Zz�ڡ��Έ��K뻏���Tdr�YĻ}��w��)��ؙ����� |ܕ���;@���P���;�y�����h�8�>PHw�����y�!�y�����cC?��9��C�A��Kܠ����r����!�9/=⻗z)�e��C8�YO��[�ɒ9���H5|�4\{r�/C�G�@�m��׈p�?�=["Һ����7����z��5��"��I��L=A3q�L�B!$�o�WO�oQ���Τ�J�26��Ѱ���������0���(w�MT9̗{r$���i��۞zk��!$���a>m��v0<R,yF6H�Wr��J~��hW���WG��M��j����S��?~�����'��ٶ���Ɉ��{ʥ컪A�Ywx���Տ~@�vu�2�̓n����
!�����rǘ��6Ƙ���Le���8{���g�=Tp:t�	�^����:%�����y�z�֟�T��5�͍d��9�!��I�.f����x���pB�tK���� �[�ޏi���=٭��$���[��"g�I��95�xq������2��~;��/��#w"A/�A&[�ܤ��0X�����m����a�������u���4�(�[�ո�]sf��{�����W/
�sz��2T���G�$�3�ż�nx���p���|��,|˜n<@�n_�è)�;ׁ�U�y�v��]vH��t���cc&�
}	�X{��6.�z��y����caٽז0�`x�[�'�I�rh�g��΍�x/�M�i���pڻVi����@�gG�+�q�z��5O*w{5�{��X>y�o|^�����)L�v��,޵�Ć ��#&$kr�J/*D�%��J�K�I��M�wI��w��4����E�Z��ǭ nwB�"��{������yި���������ɍ2}�q&#ǒh�=��3�%݉�~�$�D5V�Q]1�si@��(�"�����f��0·t&����*�a{Mѷ3f�
��+>�~���q�KÎ�>@�b��\ �1��D�1��t�s*�0�� �mD2�sR%z��'�r@K2r�d��y�V�A:��Ů�Į��Aѱ2}���y�'�����x���T3������^*�{�ލǵ*}���#��yh�foV�o13dZ����c�/{�\��͈��ɦH�t����Y�4q��.]�m�ϼA~&��x{�^���>��R.�(%=}�e>���o����A� ţ�.|�1��bC��՗�6�ç�Ḭ����A"YV�4L�mp���[��j��6�ɀ{����׾�?���r��0N�h�Y�����z� ��n\'9���\�. �~���8+���D�r	<շ�M���$h��9��R��z]�$��/Za,s/�	��6�8����QΈh$�ب������!����wL���d�y�<�>���K��W\��=�h��r@JG�����{�X�E���Ě��C��8M^\�md7��M���;��O��Ɔ<�M�)��I'ݲ�,|�N��"aW���o,i��l�{��Ѝ�^0�xbA�h���{,�y������b���=�O��h�>C�i���b�s���m~�+����}o�o�O��8�~x�P
+�}��x[�@��!疎�>s������Ĭ�VQ!�J��J ��ú�O��DI��� �+-3��䵸#�=t��f����sӧr���y��dS4b���I�4�G-����=��V�	�t�ع뗋�{v�|��\[u1��-�N��Vǖyc!+nq�fn�e)Ncn'.F����!ft%�2K��.�2��Ʌ��9��,7<ˈ�c,p=h]�j��יr�FѫՂ�G^u�9vs1�su��,Ԏ���֦�v�޵�79�-Vce����ȣ������@��@� �$��v3���"w�c3_]�҉�؂ݠ�������������9�W��jߢI�C>f�T�!�u�P	�Y��y�'���f�ԁH"�߁�!Ƈ3&ߧ��H7��.]�6f���s��������"X�N�� ��g���(��T�t�G�yl��vI_<7���\k925�n����YYgx������5d�{٩��!=�6j��'��^=Җdн<8z�q�p�Hj�Ph��$��x O�׹�w4��w]Ƶ�"�X��[)BA:S\�HF��p���ٱ��l]�78���|���Z��w�ҳeȦH��ِc�(��\Ŏ��cx��w����Б�2���AYc�:Tl�JT{ҝ�{�|�Wzo{���>�s힗�@p����o��o����=�߯�پ�u������}y�O�4��@dCAf�y��c֨6ƛ��&�v'�*�鬓k��A$�^v����2=���PƘ����^%��&	B�ѰJ����>���[7z$��^&×<8��.���3��.Y��#�[!&�C2�wS@�X�ͼ>��e19W�;~K^!D��ڷ�B���O�0��H5[�n=�ls�ʶ�1�e�N��M/T����gen/}�o�ۮ�c�e\�k�B�s�U�ں���V}8�t��ݗ���Rx����H+��.f$y�K�=����f!�ܞ���ޘ��D�70�a��T���T�d�� �A9��$	��h��*7�:�J���}�R	��4�çP�0��ʙ$�	{��D������b���fF[�Jd���W��9�=}j��8�Ŏ&�K2n?�#������o�pm����+��N}�|�~t���̝�}k>~y�}�~t�Ay��4���P���}�>����b[_�������Xݽ�x���$�c��Ĥ/� ���w_��}�ܺ��{�Vf�3��o1m�[�7��1z�Vxa���r<�����={^t�i��]�K�P=<�b��G���:��4`ɞ=w=M~@��촏��auۆ��l�xC�;�>�� �����9�<J���8��87��t�<�װc�;��cw��wh�H�i=fDz�G�Q�Gf�rzҺa���˻�g��H�;jc���Ӣ�{^��)��3�8͛����L9����<��iGC�o)���5���D����<l�&M|'C��( ��~�{8��G�{���yf�ؕ����m���ܞZw `Y�ȏ{ڣ[۰�pڗ�����^�eW�,{�G�ë���}�FW׼�8����v��흼�X�!���w=A3��9ܻ�W>;����C��%�X��6�7
M�T%��E�?�^��I�"�����_=����CU��q��ξ��w+�ˌQ�~ |i�^D~G���4DB�y��~��WH�F%�:���}�-����)8�3;ҟH ݏ�-97�����}�ϲ%���	�����`��zw�^�z6k�/��v������ѐ�yw�j���w��Q0�<yǕr�Rlo|��� T�� ��NG;~>�g����q��u����������E�<1! �NP8�F��� C,L�	 BBͬ���ֆ�������������=<d}���!$t������2�@"�$V��(�!PE\���xϣ����~�]}{{{{{{{��(���}�:�5�x�SA��
 ��T�Uc���G׷G��_^���۴��2'@�	#<e�0!! Q� ���a�RE����>��o���믯oooon�3���`Br!��d�	� @���` �N0hm�_g3�x��e��0���}��.\�Mؐp�fkhn2*"t��YK���xLwX�L��'��e��h�=S6̆.Y 
�@�81!>e�+!U`p|�	�$��+�IT�а� �`BQ���	��ȝ<H��2� 	���<\��tyH$)>}�BU�y�}-��z� �m+(�1@������"��Hbc�u�\=�3 �$]gw5O5v��-(%��,���`:k}0�V�DQ-L�<�MA�ܧ�i׃�w��f�T"���.q�֠�g��,�y�F���^��i�� ���,Ί�g�;�~�����}9�7]����V����;`�@�U%�mb2�IIi3�L]
�Ai�r�'��u/	�R;�\zcUc$su��$���P��ѝv@{���8/���n�@��OWG�ߧ�	��?refkm�M�$e�A �N7:� ����p1�c�:ı���A�h
�N�G�憓ݮ�9�z��O^�'�Q�ı'ݑ��ܠH>�m���w��S]�7{�QÎm�: �8$�ӱ  Y��l������ؤ8�*��~��H�*C�������}^��I��l��~��~.�N>�Q�[�/��'��uᰀ�0C��H�C*ؙ�Eewy�-	()�ƥ�!�5ݐ�L�*�A��千c�?� �ڒm��ސ���~�bF�×�F�ìu���{�J��rk��wmm-]c
^��"�F8ۭ
6��^٪������������s.�|j�:��4H�a����xxg/f򘬆�g1OLd�P!7���!D����c��2��c�>_� A$��v�md�Hޙ�#�0kz+[��< �H��c���Oc�ζ�#=�H�C�%�lϗv@�H��P��2i�;�0�	T���?S�D��U�AӤmdŔ�.�g�H��0ӏ�0 rt��	���n�AzҖ4ە4�wI��@X���I�}�q;<��oK&��\�c�}F�\�;"a���O���_�y��f������-��ݯ
���t��:��w"N�e��`�z^��Y�1Գ���s�`1�c�r(���.�k���b�֨����x��:�7�����e�𲩬�l��K�Jڕ�X�Y��$s.��Km�宵�7AՄ�GY�Irag�x	n�v��.4+��KYrЏ8�]"ޞ����Ð�c���K���'���n���8�Rő�9�te��F�2X���!l���C�df��K�ۊ�$Y�ɳ�2��!�m�Wpk^�.͵���ݱ�'��`��	�͛�K��n���u!�EHhW&���e��	Ȃ�0��g�FK�ŵ�z ��8k�c�q��zG����A���ܕR�L����W�"m�\Xp��.� �K_��(��>#J���@r	$N�L�L�No;&��=o�ך�Pm����u�	�Rzz�0y�bX�"A���x���( ��I=��t7�z;�w�
.���\������kϼӬX�%���W��Q1]ym豖�~���ػD�T�P+e�h^أ݌���1�����#���e�,Efƴ�@�O�г�������Q������OmX��+��HuΎ.�1�M�늋p���s=���Bw1���˦A�\�6��Mi&���x�� s _5�|#=VBQ�H�"�yw6�>����\m8_�e9�7�A�mb��pa��Ǿ��\o/���;�߽]��[�|6��=��V)]��K�K!0�C�bC Hh6�� �,M]�L�$i�lq�L�Ё��.��Z�f�m۲h9q��É�a<\7�U2@�+�N�-kguy�R�j݈L��� ���Ea �����D'���o�:�c�/%�`�/�)�2
YG���Koz}2�چ(�@&�������!����^��&\����-]��O2��D0�v�$*Ȃu*w�e$��"�h�w�	�ĄCk�wx����S�H�[Od'�l�;v�JK]���M��}���_���y8�.�q�__�g���V������ @)����e�y"��.෵t�[!�;[�3}�m��طU4�����2	O���ttAhj�PG��E/x=�62�wG�$���r6Ts�0܂~ѕ�i��SsN��I<u�;�
t4�^1{�M��{O����h�����Y..�G[�B�A�۠ �0� �! <�!� $R�PH�,��w��p=P��#�j�����Ӿ#��_�30��d �^>d���5삆Kw�þyN���{��I��o�!<���\
l{��)]�M�Km	�Cmo?D�.�v����U�:����w]�@S~z�u�	n����^�Y�Iq�&��)76,\���t�w�Aw�0�aF7;r�D9�k�s*`K52;��F��A����p����D��6HN!y'O��]R�p����� � ���	.���zE�I^k�I*���t]$T(Q8�ܪ����>~� �*����v���^�q[��-d�c�4���!��k�S,��I{��t���� �s;�\���/H���I�Ӽ����K?h���og]��<�@�Hs�xmC��g`9g�[=�w
w�ޤ��:����7w;�s��7{u�D���j ,t�� Sy�h�\s��p[�����0I;��Z+���g��7I*n�<	>AwC��\Az���s�>�l9e(q �˭L���^#����hȽ�S��,������'���h�߷}�t�˭�A,�~0c=ru$)��A׺om���ຏy��L+�uQ�g��ȇ-Aa��1���85�E�G��!�r�j.^㻪��LE1Eb�LJyJ�^oF�$ʭ�M�"%A��~��5�C.{�|����G���z}�]���͜	 ��p�$u��;�<�_J�s^{�1��e�n�aL�	(p֣е�^������2yNo�0�ą;�F�1Ơ���]�͜#ޗ����K�6�0Af ���{l���1���A�B�~���W>���ga�6�s�>�a������]-m�P���"������i.�|�Jd��Sq2���1��c��M�XA���|�h�$Z����X��[l#��09��v�͎��y����rK�'�^{Yŭ������wP�)q+���6.�d7��J��=qݬ*��8�肁XT��:*�뢛�f�l�f %�%&(0��y��c���m��=�.A;m�䳨bV�o,��F��
m���Ǖ�Q�����F������u��#��H�IE#���|�E�^ā�gD�w�rۏTȱ'��f�,Ӝ�˞��YL��A ��Д$!�%芸��5rOz�4���48
�����<�M�L�wl�at�7!����y�:���/!�\�>D1�vdQ2�z��nO���1����a���Ē��~����y�..=��"5x�G2�|��ȂX��j9�3]�	�x6�_&���
q#ئ`	������9pA��)��WwF��ch���_�H}�y�9������ ��ń�%�o��n�Љ�pQL�B	t{6A����#m#(`�TC��cjg�(�W{��]�d�V��A$�ޖ�:�D����Oz���D@=�����(k��q��1t6ɟ�뮷����q����v��ǯA���w�]���W>���٫�ƅ�c�����샮�,�oc��{�-��]������B��tH=ّm������/} �D�??	�4��٣�aC�	+���&�(e�L2~�7�f���#����dȆ��oDvn{����ƃ�t�v?�}��s�W5�Ędݽ#b�Z���y�� � �/�:�r�f
I���T
�z3y�ʠ6:d���H�z�������;���y����?�D��߈r�ݼ���`���eጹj�d��2�����|���>�Wh��H�6��^� {PO�.�8���Ύy۩�ɢA&���@��-3�*E`Ʈ�g��Sƞ5���K�,���h���x�#c�;q��t��F�xj.P�u�����#)Y������%2󰅠�M�L甏fDC={�yb���V\��"�͵�/�h^<��d/���+ו�p�3� C�O�$��,Bm]�	VH>��:𒻐'�^�8_�6��oߡl�@D��WkoCE�D븼'����.�����රb���zn��>���Aϕ�O�ӽ^��2S7	�M�$b�P	'�� ��༇ȑ>r�@(��� 8s�fׯv���ɶ�Vɫ�B��F�D��j?��{�!�Ь}h�g�%���@)����n����W��Wy�L�D��P	����`�D:N.ۀ��f&x�ֆ��� ��-G,kdb;����2W&����j�#?:H��Pz�4�q��;���L����~��m3�G̛��@ybE�Co�d�� ����!����*��1bU�&�[,�M��2	$���y��Ws̳N���;j��!��޾��o~�x���wZz�=5zA���FuT�;���i�Q�
Q$-��]��w���{¬B�B"[s;��{�{c|�q3��g���*c��C?uM�����~�s�y�wW3�a�����ȥ��s�Gk��N��Z��˕Gml�(1_�矂�e��j��:f����Y"[�r��S-詽��){��	bi�o?d�I;VP�D?�HtS�������p��� ��g�t6�'�2	���P(����v3�&Z�p""!�'Ι��"�������ޞ;1�n�ꮮP��ٓ,Q��MR$�g�Ias�-�����-tĴ�|ꘒAv��Kr�J"�p^��{�$����:C��ځ(>�F�n�ƶ0����)�����+y�ux_������+��?�@U�H�"�������x����T��t �`��8w����J�*��
�Ь"�!(�!*�J B����EXB� �%U��PE`BV$`BQV$P�  B@@�T%��z� C� !
�@��	�$J��!"������@�0�)�C���!*��G�� $B@��B @�@�@���
�$@ B%  BP%  B   BD<�*�� �BUX� �	@� �	@� � � �	@� �} �J @�(J @�B @��J @��J @�/L��t�P$@ BP%  BP%@!YUa	BP$@:��@� �	@�@�	@� �	U`BT!  B�TyJ @�(J @�(J @� @�@���!(,B��8�||��_���*("�2(*�P���_����߸?���?�������C���� 8G����@~��!�����_�:��W��?����(��_��*���?�?�~� i������O������W��a��/���I=�z|�����9���?�~��s���0��" 1 *�
 ЌB+H� ҤJ�D�@�"1 ��$B�@4�$�J1L�̉B2@4	R���� Ҥ4@3ҩ,�2$�$J2�$0�"HH�L��$�A(�
B@42$$P�(D�@3�(��"ģ+ Ь!Ь�4��+�"�%�#@3
̣�J2B0J2$+,0��2,�$�,#J0ʒ	"R,�
�$�����0!(̋�!�(��#!(�(Ќ"B��0�@,��1
�J0�����
��(��"�J2� ���2�Ȱ�I
�"�(̣2,��0H�(���+$��H�"ʄ�2,ȍ ��̬�3ҳ2�+BЌH�ҥ+(�B2�R�P"Ј �"�J��IUy(*p������}ҟ�AQ((@hTT�P�O�>���?��?�����Hv���O�}�'?o�@*�a�|���?w��tw�O�b��� ��1���N���?x
������Z?ǯ�L��PeEW�j�ç�C����vt
 �����^���*�O������k���s�a�����;?n�;:�����<�V�������/������@T_���9�>}�q�o��g���;���A��~�O������W��#�?���*�����x��{�i��p>'��?��������$���P|L��>?�@���������_��~������ /迈�: Au��������!�	���
�2���ym�#��� ���9�>���� [ �� P � @ �4�    ��     5@h( )� _  �� �@��@�@ Q% �m� (��PP��@� �� ((B�	  |  �      �T�      �      �   @   �       @ )�|:7���i�����U���]p ;�֩ͮ���}����֭�ݨū�;cT� �9��)���2@
  ����ZU7Z�l������X=i��u�����t �N� @� �l-�����,�C�t���y�����;���� �����  �@     @1�E��`
��y�� �v^`w�=cC�� =�vR��73���u��K�)g<���۝�*P�x �S6��J�6�k ���|  ���S��v�Vڶ}� {�J���٩W-I��ۙ�je�ܱ��} ��T���3*8�$��rԪ��҄@�@<  �      �=
K-y���j��j�ͷ;��n ԒVZ�[j�ĺ�[�Шv:u��� �]2�wKI'-R�


H��  ���ԩ>f�b������uX�:��!SN�J���P��vҕ\�H�4�Ґ�:zz�- 
P4/�  x       zUL�\١.Z�+�suЩ����Ng s�����tI'!�u�;��SQ� �.ƶ�M�]eW*�T��M(��  ǫ�}v�7�j�i� .�{�/Y{[n{��l����	���%� -齛^]v���]����-Vi�X�%I(6�{�  |        7���^w��[��ٝ5�u��nn媦7 εm���z��Yzuz����z4� wU�r7}�z� UB���  7^�����y�ڴp ;�E]e*�ӛzx]V޺�v�0��tv� ,��V�nժ���L�m]gZ�';t�>���JR   �~F"R� 0'�R�Jj� �j��SAJR   J~�%A"   j &�Jb ��������w��T5������0���a;�����$�	f��	!I�! ��� $�	'�H@�Y!!H��x{��k����s�?������ٛY9$�X�Iie�F��iՌ�V^亸�L`b�{��k�RV�tO��^)����uG��b�ʦ�֎�.��6��An���%����Ϯc��j�1��"l*f(�e�GY���ٍ"ګ��C!�-��4l�ٶf��`��n��Ֆ��v�Հf�Fk�d�FfM�uj���c��t� [�gNQ�\Q�ߎ�[gQoK�W�l�l�Q�w1]2���X�n��J���>�Uޔ�OY�1��A�ri7��u�48~re-�k)H˙a�n��6��I3��iT��R*�HS�b�σ���U.���
	լ4�)�u6M��:�1��Z��˄�d`��!��[���x.�3w{|F�D&\�[�ٔ��+�K*��JH��F��F���8��A���U�)�[��X��,*�ݚDS.k�/
ؖ	`e_ٯT��'�ޛ��!z��+vV�b���r\�Ub�hf|tV3��M4�X�ܴ�����v���ॶ�Ҡ�b�;�� ۊ�������.�O�,&�+n�I�ؙB�^�Ǔb��i�fme��@�;�e�ݕ�����O�q�l9Y�l�f��@�#���'�M"����x�r��V���c��wb�l���ݠ��h諹n�iP�ʇ�E(%f����b6.[�Db�֌4��Xk(rr�Yv(̻���J�;�����Sd1Lɛ��/���g��\ʣY�<2�	�k��l��1�8�[�<���r��Ƒb\�֝]��p1��7.����p�3+rQl�x���Ip��wV���n�}/�e�����ۚ"�����&Ӷt�hHŉ�N
��Kn�lL��-R�Jm\�4���ܺ{��r�G� X-���݇�Y�[�e+�^�".���\0��U��Y�T��λ�O�����ۼ���vtM7��aY.�kȉ[�?+ي,bK�%^����e����$V�N*�F�fXÖ���%O%ǵ	����֐���kb5�JԽ�ɹ�H�r�Q�4�e]ѻ�[2&ʫvk��rlMh�'ۻ͓d.59\��[Dܷ�(��h"l�H��B��n+��È�2�V�lZ�V	W7w#�=�4�[È�[N��8�YL���������&W��b�����&����[J��
ܚ+s�ʘ���9�b�[��rbE����j��/r��)�����$�Vn��Y�INƑ4n��,^ۗ!�`Eb�gt:Y�bK^�Vk��n�F�dbg5�V*�!h�S&kFh9zr���+k[V+jn�ܑf�+��諸�Ck.cN�����g�4]e�X���%����;j��I��(.��[jU�V�VP�f�&̢�G6�[-{�x�/ұ5<�	Ԡ(���#�.j�׸�L�z�Qq�+P��1��إ���8����R�ք̼����Wt�^�r�"�e��a�0��7$�3,\���o[7N�eeV.;�2ŭ��+A�ԑ�ɺ��d���*R�Hm����p^�ma��(�K0T
��я6��ͽ�QQ�T�Df,��a��)0��ӳa�o�in+2�8�9�"����u���G��ɊXNs����򖖺I���Q<�Yy�ӧG^�`�Z��ٵp�w�e��e��7^�^4�z
��֌�6��#��|b4���`,�{�gv���*��n@��t�]�t���kV#��X%���X����3��m�
�hҁ'W�[P6��X�,	�����gv��NQ���G&ި^�%Ѻ�p�a@���%>�c@p�I�;y3�.�7��%�ͱR��2�:��a�EF��UJJ�QkZ��7�L�Zv:Ú`�j�ʁ�湲�V�Շk
�v��7���0��IDazi�����q�hM�0G�EmK݁<*�/5j��b��I� �Kf8y���9�o�3S�
 �j��m,�jy�V�۬#������.�]VI��KR�M���M��:{1^�W�۹`�c*m[�(���lI�xSRμE[��V�嗊�nJw�z�ӂ���С��	�nD켰4V�y�; v�q�V�U�͗v�c[���:&�y����x�ZC��Lxoq�"�[%ъ�@��,hڻ#6�l.ཻ�ީuH�5t��Pb������Ղ�e�PN���v�Ė�d�i�B�:Rf�[kv �$�\�U�ڬB���6bⵐ�$FB>a�WV���^�775G�8����]�y�u͌���R�ZL��V�3+�ڕ
Ϭm�^t��)�:�ju����V]Gxp]�re�T\�YxK��A��<�*�����/]�����k6ݸsͺƵ�u�!ˬ.W6��IywXXͭc���`j�tqcٲ���EF���#Nܼ�ek���F��+m5R��7q�q8Kr���`i���ۡ�i����j�Y��H�.lt蛨*����R��f�K�"�3T-^]�{�S�n0�7j��Qb�l��]kȖGW�
�
`�����nm,ʲ���W�1e�8�����'7Qу)�T�֬���b�٥�5��[3Wf�AJ�}`:8�	�4w�+6VE,G��[wsj!�Yb�����Q�C%ȶx34�V���6+����I+cZ�eϲ��ڹ|ML��P2�����9�1-��5nZ��֦`�e�>�V�8U"ʒ�Z�w%��6`z,��v�jFMm�mG8e{�7���l]�5x�ʌX6@(kR�Ŷ6�\LVm�˳3�b��ٛ�G*�.��1V�4�zc�1��{Е:���*�`blL�p�-�+3V���F�<V���y�u�cҲ�,hӉ-͸�%'B��,v&���V�y�e�<ջy���yN��E�t1�l^LN���u]@�$R��Zq�4�+�Vh;;&h����3�6�iDj�H��[yb�g"�XP�T�V"�"+(�[{�⛗cn��	�2mK�z/7N֋�W�Y�Z�hI�����.K7y��Gn�0X"��a����c7a�z���,�[,hV��'�S�7Q�.֒3.��3���/R��ى��T��x�N��18�$�"��J͈�e����Zv��V,	�:Ag+b-L�L��c��Z+Q�9�e�I����c�j,C$�謰�(�m���r��
�c�D&"S�j����k$-�5� ��n���N(٫.�fB��6`z�.�;�Q��D��*�p�����ͣ�+"����q���1�D��9�xH�xs6�m�sK�ެ+x��[�*ǯa�}f@�m�v6eP���u{������wD��])X�w�+ň���8�k����LĀŶ���ki�R��Jb{�1!2�X�"X�v^��n]c�R�Yz�'��h�ڻ�-���X�H.҉�P�c2�F�khmn)��V0�yw��h�(��Pj�4�ov;��D,�2��AWg
sqbͻ�n�Ӷ��v�U�P��陌�Z��d̺P���7pj����\t.��&����3)-�E�tq�-�7�L��vʚ�GFf6��B&�4e ��ldR;͊�Ո��QM�d�k�����C坰����X�+ٕͫ�h������V�h���[��f�`h���3_�Yn��19��K$�
K��B��^m[���!����a��l^֓+5Y��Nb�[��-c���	�]��]�Dn`�{� y���L*1"��9sH*&��h�z�*jv�}� �q�`�ku���K*�7Ѡ��Wd�Q�{I�re^:֣Vdmd�M贴n���y�,��u��k�Y��kvj��f�C 5��X���!c\�wd�r�<�xv�ۙP��yr����kkV]'�e\W�[6[u���Y�&�Uz%���"����`W�	#[��w��^���:�j���{b����ot�v؛�b�ĸUec�	�(�ɘ�l��k��&�N}i�I�wX�ޅ#�*+"�õ�N��:-�V��,`��њ	;�H�/�(�P^;����n�G����6͇EnG[�}n�����c̥v��P����T���%�-����51��.�Iɵ�Љ���ɾ�C6,�a�����N���%����q5Ev�U	�H&�oj�
@(�%�L:馕���rWp��N�f;Mj�1��W�y�M�l��g"��F
�H,�`a�q���l�^�}����h�\e�|]����֠��yx뉔��Ђ^8�D���{i=6,;��Dsl�~����siޘ!�3%Z�ӣY�M�7tn孧4�oq
�2�Ei��:i�ȅVQ��e����證��$�"V�4	Ub��%;���Y�S����v���`�l�b�%dʍd��9�
bF���mڔ�	JR4�8��J����ͭU4=�Y�l��c��rf�^�9)�h�H��6�$�N������Y�PIdM�Q��:N�ןR�in�tb��cY�Gj�1���M����5b�Q���;M��HF�2�Ve�kE֜��;z����l�ؖh��e�P*�� �9�yx/5��j	6Q�G��dB�#S�P�ѵ�/u3�MU�V����Ge���&�0��8p��k�c���4���l��9+m�:���fe<���^r��sre�8	N������'�{^�^U�V�]J�a
��F�#��h[Yp}d���E��ǈ���Q�K��-�*ͻF����l��)n��� ��Vf"�kN�%˽RQ7��u�b)�5��]S
��5kr9m�j�0Ֆ�<On�:�w��ùR�)�{�����f�H��epIW`ь���I��	Y&V7tt�x�՚�V�a��(���oNɮ��U��wWyg&b���V�ۍ����Z��[ֶ�������rn�33RS%(����m�M�Zv�D�I�.ƜVoYۺ'5�=M��l�p�V�]����ҹ{e崑�0M��=n�Ԗ�22�{wCen�J�1�j;�8 �t�[@u�^^cX�ǉ��N�5,����:M�t]A����ӗ@�L=0����w@�I$��J������ڲ	/j5���Ò��VTˠ���j��OA9u�W����8oLQ�۹��^���C�j�`it�P#���V�����jTz��kX�fЙXU<j�A�r�+"%��A�o+7u��w0�R*]Hww^`�P�5nѓf�[Q|@��g�Rۢt�y�������7G/n`����Q�L!w})����$���:�tȊ���VL����[F�]��(cU�1�3��Db�j�Բ\h�a�B������9W*dG.���-!Jوw,��'�캊HX��U�5,$6�4^e��u��/e�o-k�8K�¢v��y`f�o���5��Q=����G3"�^]����K׈�x3w,^8��[�s�7����X]�Qri�I�iN;�]��Ba9XM��í�[YtLE��{�X��q��6��ݷB���#���A�Re1�3Iٵ��[J��mMUfVaku����k0�*�b�^�`^]M�̛H�������vXkYrd�[�m]!�!v`J��^]L�g��c׵�##�����#�Y��r=ImՔ�!�c[�vHҴn40��J�ٽɪ���EV�hfQ[{e�"��t���p�E��pYYFT�vazj
�+��h�9�,�.�[8N2��@�Y/eJRB�#�2!E��>R�Gy�櫚	y�o���h��>
�gR�ϞC�R lua��R���Kf��t�yw���
�%ʷ���h��w�*�TI^&��hkݲ�עU��t�YkW��X2�Ź�]��	<���cώ��f�bL��.-���ѭ�Z�)NM�V� �WI� Zr�-_�J��a�ur��D�̇3	�&c��5^�;0�"^���l�ۙ��)�n�(�ͭ�6���tfU�~�˛Ch�P�kv���U�"�����b��,'���w]�Gu啍���Ӱ��N�k&�&�X4IG.emj�^e�l�{�d2XI���2�65�\�V�;�Ojb�X~[w*�y�h"Ճ[�f	N,�����4��TyrΨ�f�B�$��w���U��fSD*�ӑު �{o2e��7`�n�/-\�R!������{�����sʆ-gV�$N�Y5��i*�2�>Y��2��  ;�c|2�bL^�t�U��Uv�S��!Zj��Q�m[������
l��7^�eP��3%�w�b��dl�{kQ���1[Z07B�:tM��\AX���Y7
���ώ;��u���4T�8��ң�Z�C����:RهX�2�;(<���o,g�c�l7{�^:P�]�%���x/BU�2���Ceʹi���	"��Yv��L)97Z�⮗��u�C3�؞�ݛܩ4�ú��y��s^�O��aѱ+M���6��Ǝ��M^a���^�T.��}+��V@8�g'Z�7�d�%3{�왶���ݨ-�iJU��(�i4�YY�U��ރv�0ր����f�ۆ�Xѿr��������.��ʱ��pn��7L�4jwJ����9���Rml_An��wL©���w)�d�ī��ˬ��xʊ��[���Ho!36��2��L�y�r���n���J���<ĳ2#(m�y	{x�4�B��`Jʌ��$��]`#BS��P.�v�mVɑ�N��%tԪ������B���YtwM+
�%��x�S��I�8/]I36�{u���U�J�i��mސ��s8���a�rW�y�l��7�b�.���TN<OeB���ł��&�T֕� �Or��0 �nE^�ۯ��ʨ�c�u�d|�����y�w]]�wu�u��u�Eu�E��w]Q�QW��wuGwt]u����wwtw]��]�����;�軮��:�㮫:�����:��⪊���룻�.����뺳��.����:���N諮;.���:����⺻����:.��Ϋ����쮪�����:��긫���+���㸻�����:꣮���Ϊ��ꋻ�;������룺�.Ϊ���:�:�����κ�����뻋���ή�;�.ꣻ�������꫎��*��:��������뫨���꺳�����������ꨮ��볻�Ȑ���	!!�I	O�0��2d���/>�����BF��i	�UPF(�Y���%��B���9M����/8^e�*�к�y/X�K�0K�yg�pVM�w�s#;�����f%���}�Y1�����b�}������c6�ݍ�������J+4T��L��osl5����nv�#�.�j�"_j#T�[(*N�	n(1�9�rָ�	W
7(�^�.�(�[��qiR ��@�yה7(r��n�U| 鈧��n��"��X\�޺Osh�Fks'I[*�۠V�*�}4�|�dJO��(�RX�7݉��ZB}����s$��̓5�I�����������m�f��,Q��JVk���)lk*B�P�;u�A=r	�e΀�bn��w��1��� ����s���=�8����AgC/-6o`�X33kJW�67�����u0���h�P�(E�vo)����v����=��R���\X-4�y1�����y�V����N�;�|�]Z���������O�]RIv��es�w��h;����K�Q���F0N=wCq�k1N�4���Y�Z�^ޫ�xkz[��̬L�9eŨ.kn�pw&(��w���=���ϲ���a<{z���w�t60����2e��Y�*�����2��QM�Ю�s��Im@Wm�#���i����V|u���^��j6��5�1�vD�>7
�GHŁ#���ƪ``�a2rk:+V-��źq^-�o]nҙI̸���W.�G�����7+���2�4��y��7e^܂�+;�r�|xU).�s��
�F�`��n��V�^tĴ�����K��r�0n��u�[�.�����MՀY�j��G��KB��GWk��oYD��;ܣ:��[2���Wt��v��;m=��.��h5�c�J�bN�[I:IX���V���%ǊV�'_�,5j�ݐ�%.�Om��3���I�U�
p-���6��o��(>+3�������\#y4H]���nr��y�5�Gl�/���R�|��d9K
y��B�	[F[��/��8�p�%�c&�.�X�v���Ü����̋v��5�"6*�g^�Ow@�b�A�K4tj�)����%RQ]Bo!��Ѷ�md�(9*������j�)F1P�Ճ�y��l���vg)1���.bX��]b�K80e��ݽ�.<b�	9�VJ���2j�#z�k�79TmS��&�R�B��,�;�;�ޗt(�Z��9;.k��z�̕}���o���7/o���U�Zޫn���n�"OS�n;7t��0���l¯	.���A�7�5�'�z��"�!4���|��4�W��2��6�n��Qs3Fi܃1��R�!2�e[��B�+u��9��7�lwV��wv!�T��U���!��(�re^������� ����b�Y�u�n�T�9c="�\���(�[Έ��� ]��"dRJ��bn�D��{S�D��@�@��:��U���	]t����ͫಓ�}F�H'�	A�r�Z�Vu�)�����\���9��A7���{4��i6w���VՔL�-��g�Q��qڏ;���t�BuL�x����tnn_�tu^vs�Y/����Ŷ\F/�^�%�e^��>¸�[���ޔ%�f3�̔5�{J�s'�ݕrv��A�$}�Z��yMmLc��}�Զ����wl�U����Jތ�c�ܺqvS����|ru�m�{o.�DLB8Ujp"����xq�J������q��,�U�j}����~n�ZMa��L�����n��]�w����pwۛ���˷k&s��E�μ�Sa�m�ij��͊pf��h\�����b,�[+D����`��OKKbj����`e��w�����M��Ot�n����ڊ9Ze��w����kD��E�f&Pob#F�I+BOf�%�������!��2(�v��C4MԌ�+��T�'�k���˫���3�={�gm�C#�$�L{WlS�@����x ֺ!�6��$���mѸ��;=�5,Ń�ne�s�=Ɍ�T��i҃���2;δ(!N��Շr��d��NkO�R��ִ�e8k�V���e���yF����^D�^�b=9x�˛q�VK�!��$�o�(gc����OkJ��n��Q�
��tTӖ���Mu�n��ػ���4͡��{:ƀx>�t�w�\��������Ak��q&�lϳ+F��u��(���Y�ݘ��+�bk2�Q��J��U�k�O�� �n[+������O
����W��)m�ƪ�gED�p�@X�R�x�½�v�a�1�)1����)��f�u����%N�v��)1�{{\���ʧ靹�C��oa��k���E��3���w�eXֆ�6��zVz����f�`�S�V����C*P$�kk��_=?Sz�'��@����ӫ�fnE�b�R�����E�l�0dG�)�o O� o1���kN]ɑ#�c&l�ֱ�q5�-�ض�%�tWa�p����y)�fc�J�V���A@����O��Jjsh�=ܟc6�݉��fbv�p���Kt�@�*�>y[XJF�jv��v�LF,"��\��T�rrk�+mU�p�6�\��h���rL��cv�q��b��b�k�M�5�1	�v�죢v�ڴ]�޴�EM|�l��]�(r��N��h�T�� �:YBs�u�Z��koc0����`S�t�����+�6�Ú�i"�q�P�Wڗc��Q�ˬNۼ�S� �����q�A��-`��ݾ	,�h+�&2r $�+u]�)x���+3o/t u���g�t�'3��K΋��[j�4�m��C#I�	T���tb!��b���ɖ�YG��#=++n��޾y62���n���v�\1�cX��-���P�(���^�!t�L�,n�~�~��욚���/f.��J;c���E����s�vТ���71h�q�{�`Dk���!ss��>4�t����*�k�]����NTå��ۓ/u�}����:�;�C�ʙt�>��j*��jر˫���DA�(�ݛ$=*f2vZYFS��S�$5�z��ZrKܴ�׷w/f�;
�:ko
�@��Y��;wu�Dķn��n!��U�A��s3�3X�5}�u���w�ܶ�n�����hb!Hs���s�e�QU�G�pU�g�/�o�����]֓���ōS����(�3�+z���$	����cV�j�0<3Y5k���e�i�f$�N*M$�W�,L���jdM땩��Cf���7��%����Ų�]�X]f2����$��2�|��� �L�|�����9,�oiɜ]G����k�8����"\���n:@�ѓv� �y��"�c��Mwe#,F�'|e�I��!B.������Y�Vb"�Zd��d�]��ף�U�^�t�$��1YJ ���@,�(V;�#�s�5�y������r�� �U6
ߐ�r�(�
�>6��0�W�s�\�ӄ���C����yV>�����W�&�^��
��c��:�T$XĒ�#j
±�Z]���N#Z�����p��xh��;Z��(%lt
�����X���m���.���[��ֈr�K����!eR���K�2v^8^�1P��ٕؔSnњ���6��]�ikF�yVvbK{���{:�����&�Ik�߳>�;3_]�4���|^��k��D�6�L��tN�#���2$M!��jɸ�!�Pr�E�J��<���jp�k�G]}�gWW*G��m$�"�;��*Co�>Ed�+u��sU\�1��]o:0��1�f����8��u�Áa�{�x�:Au�m�HEk�&���zXs�A��±��y��m��X3j�*�[�^+ji�N6^f��0��Z��ܥvv4]L쭠����N�Vur��2��ƫ��4=Աd�{pv� ���{���K�u��n�.�D�;�͉`�Y����t�=gn�}t���N�a�`�d��I�.�ƕ��n�흴��S�cA���8���|��Ρ�4n�Wҟ]q��ɧG��bKv��Ӭe��\Û��
tٔ�����ќ�
�u7gn,7�$p�h{������x�g_n�:;<��!XC(wEl����Y/B��:�c���ՕJև	�6"\�,�7T�Ë�#���,p
�Hl��p��y׼(�L�A8��f��S�8��,j�	�ЧW�����f�{vYϭ'��e�*�ѱ8e�.�)R���s�VI �̰��ZZN�<��ǖ)�۱����Xo��8��(�
��x�:�,��ɭC1���R��hH�=H�x�\�ۜ+	�'3�r��<ͺ��M���^�y�bg.K�څn����!n6s���
p#kE,w@�Z�N��Y�⮭/T.�Y��p��{��	�U��[wd;�V�8�4��0��$��ݓ�)z(j�t^^۸��BUڣvք�W��БP֍�whP��S�e阝�݊���F'X�����΋�w����5u{G�<e�֤B�5_k<4�zIU�u*��Z ���th_L&^%��&�Z�vʏ��`R�v.T�ʈRp�Sx�\����P��μ�ͮ��DgQw���Wt�@�V/K�&d�M�"�[�$��D/��78	��WY˭�^�15Yu������rm�yՍX ����O"Üi�ٰc0,�4�J�o�C:���͑�
Y�i��%�{J�Cqp�7$=hs�2w�2>�"�nvݧ��u(���:F��s����XQ.��K��x�c�u���Ch��&_\��.t�n,��a��Ӟ	/[��x��ܫȚ�CL�D�Rq�٘�����d����Ꙃ���o �̛�h��erv2���T�{n��<�x�Y���W'څ�n��b���̛t��ƈȖfE�n]��4���/�1���ʇlf�n�k9���N��fΝ���We	����`іv<�����%Ҕ��o�l�P��Y�G5=@�����{�G9Ɗ���˖�Cw�o\�$I��e�P�
�g`7ۢ�QҩjQ�˅S��g,,7W3>	Q.eGE�G�r��[L*��n�C���xz���Q�)A@'}۳	܌# �G��o���ɷ3��e�ӂ�F����:7�
�\��R���l�C��3{����:��M}sa���	�I���e�s�
��VL��;���b��y��}�ylR��p˧sbo3M�Ώ8hq�]n���`���w}2Rv`׵�@��9V ���&��ˣ�u�Os^��jѹs�C4����fS7[ۢ�#����S�[��β*$/%s8��3;V��Z�H�5���{���-Q5��P���RC:�n�˽��ك]' �'^u_)�m:Y:5p�˩|�R�I�p�=f�U�ٺr&�R��D�m5��wh�ۨ+r<:���{�U����f�-��)X��I������n�퉐�R���h�F�ŕ����-
�׊��L}�;o��Q:��5�M��ȏ"�9��b�inKT�Վ���#٫X�cu]��ܵ�����M+�v7�|���.,�1景>Ʌ[����v������_X�ʰ�Wú��xV�,�OQ���\[(�{2������<��}&�kW��N�j�M�Om��1��*�m�j�	�Gt��4z︋��3�A�\q�0�8ܬ��C�]�����t7>A���H�h^<�jɭ�|.�j�C�x�yᵥKwJ�uC�y�t�v�1T��iu�Qe�Y[RZ�;����[�[O{0�Ȃ���cڣi��L��%Z�������{���E.����9}��qg!��"��/f^k�wl�]����*b�6n�R�zWW��L޷8�}�]>�#�����&�M];`f�D��ŋ�ǯ.Qz��;d9�si�@\��\�۝��o,�VQ�z%����f>�3I=�}�[��C�3hh��TlRoD���`���{j͎����m[޽��H��}A�2r˾�@�2���7s%۷+��uh�Zk�b�ty��,�Zr��m���%�t6�l����u�=���Vj뒯��4�1jۗ�s���4q�k��̧f�#�{2�KmLY�˷���u�%xE����]:	ѕ�RB�`�܊f�;B�{�r]Z��n��֫G+�:,�8oP�M�8�סR1z�IcuI�S�I�dA�4�ׂh�'7-�R�nH��u��9�f��,w\��w&VC���J+�r5�I}�GMݺ���8��|Eثkz�;Kc�[�9n��
�/6o� �;F+2�=�\�!��*D0¡�KB��Լ�8Kj(J�(L���
6&mҤ��6���$4���j�}X����+��tC:+J�4:mt��0�-GB�ˁ-��*�B�����of*-����e�6��g��#M��z��j	�I)w�t(v�S����@�:���ĺ�6����ݴ,X��7+��%_%������@dǜ�m�
iTu����];v>w���Wϓ�\t�%h�s�y}W�s�E����T�����Z�B������)Qc�ڈ}31J�73L��{��}��X�O�:r.����xk�����4�ު�b�6cη��u�VK��u��.�(\��ő�ō�*i�}��R�ɛ�$�Y�엦e��(�gE�ѥff�l�*�ZX�q���}{�sfZ鴌{xܩgcޗ!osd^��*�fb}�o;-T��F��oV���[t��l]��1n'��:��Yz�gq^<y��3Z���)�7��V���ŮH�F�������G��'U��wN��+�5��K9mkGH�����n���칦�q���jIN(�.��F��=�]�,:��G��O/v�0�b]ˎB�Kܹ�w��ZH_t��2�f�9�6�m�����q����&�ғ;$ӘS	�(��t#�@""�--Q<k�����$�$�߾蘼aZ�5/i7J�f�k�%�KO-�f��
�qdn;M��������4��m� �k�q�^��-�jz�l=�)�	�챛*W��뇌��z�\�v��ʜ��mu�vk�8yw���m��n�vܺ1X�*�z�����넆=�Q���nx#d���B������:Ay��H��n���]��j.��sǬ���`'q����[Y�^��g��ף��bv�l0��Q�BM������$<l�x+��5�Jq�U��'������z;]�e�}64r�=�uk�xzws���[��دXv�p�
��v�ݯm����{���:n#<��.7FO;�t���[���ZѸ�ާr뎒V��2]ɗ>�:Ϯ�&�.�NWf;�0l�;۵:�vq��$A*b��R�*:D*	J�n�Ske� .�`�5>�l=�Ļ���G[n��!���ˬx�,��A���r��؜Q6}6�O'Q��b1� GZ�s�vݞ̹!�R�LĲlޞ52�vf�3{�j�퍛���=�ú�
��ڳ�vwqn���sN��]�WO.k�m�=���3�v5�\[�WWi���uM=�5��{8���[,��{d�:���ɡ"�p����x5t&kA�㫻#������ͣ^x;P��)�Io[sv��S�[��<R�K�^�wG-�΍�$r,��� �b��v�۶K��흇����,���r��Y�<�!�)��,�m���g�9����v�la�7vN����y|f8���7U�u�vSX�8�F�ۀ=\U�>۔4��ع�MΡ����;9��r��F�뇷#����w`��K��<v��V����:�����`!��q���5���
���㶮�:�`�����Y�=�]�Z���/\竉�<;tc�%�jD;�k��n=�����vb�<<�gm�����K��[]�7S۝n�����L��뭮1��q��۵Eذ�6k�X�{r�u\x�,�nOW������;�:zBcj|�۴�ѻ;���]رv=��積uF��l��Ͳ�F�=�n�v�#8݂�"�&Q�k�(�P!F+,��cY��6{�Cg	�{k��lպ���ƲT��mk���@��G��J�Z,=��2�(�6rض���ۮ�Zv;yN��ώ9��q\O��r��q�DxqM�=�bz8�շ�e���M��ܻ�uu��NF�sv��T+c���mv8�L$�k`���:�ׂO7g�r��3��6�cv�>.,Lte�>��[;����\�7Xv-��6z����{co�˷:逮:�s6Ym������3 뮺C �w5hy�s%��p�i��=���Tͷu�,��@���L�Y��}5э[����6v랓��<���	�9�3�n�7U��0 ;*�2m�p	u��`^�W]�$����ݎ��l6d��\a�<�gV!�M������t �˴�w�a������KKﶞ���k�$�z�ez�x�!�3���w/`�ܤ@샲�$M�Zp�����(�:�-�ގ�=���n�ӛ�|�|��[��%6�۷;���;>�>�o}l��z�;f��������٘�vzJ�q��8TW���hW���6�k�LF��.�v�<zl�ٝ�B�ǥܧ'N�����`��G�%�\����B�粳+��O�2���ύ\:ۯkm�oZqJ�N� G�u��M'��Z��T.Q�����筍ݚ{��^���>��6�ֆ�C��wn|<�H��t�S��l3� ����+lu;g��n�.=I�y��L�Mvk�&쪖z�f1v�8Z�PГ���q��ާs�¹��j��Sʶ��xG�Vn{��9P���f��7"��Ѷ���.< &��:��n'����]�z��ۛgş6�BR��l�@����g���v͗ �n=h��m�b)��}F�A�t�ךu��˷>k�y�÷��C��d�����<ojCuf��x���ț��Wh�p��:Λ]�wU�u�ێn�v����5�{{V'�ݩ&,����]�*g�r��/m�7v�9�ʧ��K�V�{����L�wj���'b)�k��<�j����rv�
l�=r��5n���zKOuvK�<I۲�ڶn���t����Z���A�v��;e�מ�<0a6"�q;OX�&���H��9쉹k�.�����T=�]�JeE�g����:��2��z{7]��v|s˛a�mr<�ZZz��[�R6N ���ۜBݞ݋ϰ��U�O��n������s���+����Ӏ���X8������ɞj7�͌�����}���n9�
 �s۱p�:���v��`�-o@-�ݺ��l��0�xc����Ϟ�U�N�wv]qˑ�wu��|ggZ��Z��瀶pnn5�S���.Հ^�#΍�9��^�۶�q�������)�f��n�zf�ۀ���]��<�x����ҳ�{����׶۫�1��pcqF;ikX7�jx�2�������ۖ�r��A�!�Q6��<���Ti�s^���	��ڻ�v9�yjƶ�F ;Y��6�U[n��.{s���I�svU����6�g��u�<v��:�tƷ>�}�V�rt/WU�%٭�9<��[Z�^3�'V;F�١K�2���N*I��k{�����7V���L�s��k��y�۶�i1�X�6kV�jȸ��0箁��]�[m��lm��f�Q�\w.�7�.z���)�k���]�Je[8@�m��t�m��I��P���x��g��[�KrA��n��1�Ο؋�4X+Wg��.8���Y^���ۣmr��S�C�pm��^���'\�)���)�O��s�K8�ل�S����N!�ca�܊�1ֹ=��)���0��X��1gn�moVY}k�ə�u�1�������s��ݝk&��ݼ�S�ʧa�#��z��c�B���;ۧ��P[���nf�K�����nՆ�C�OanXgL�݈�v�q� p/�OB����*�z� �x:'��m�.�3��v�>�5�x�"\lpK��O `^�w+9wZ��ٸ��[=Jٍ�]'�k{Z�ʳ�v8�=��r���f3��PqϞ��\=�ݩ�G\�O<��t�Kƌ�O����kuÎ5���<�pz�)�`ۅ�r^��H�c�s���mv粵c�gt�������5�<�DS�[��Xۛ:�	wM�`��Z�p'm>����[k\�t�ƅ��_<&{��Nh���nG���r���+�npvgs�H��4ckvݼn/j���룷��'d.Z6����[m۞�7n.���[���u��ܭ ��&_=[n㛜l�2�;uz��gZ�4z=��g	�}�����nۮ�Zѷ�F2�����s�]�������t��:����Ӆc����T�Gn�fg��v뭷[������';u��bp����y��nIqWm�������k^����qB1z�F��^�QݴC&wEc����zwF.n7>v�M��'����r��h��r��������[I}x��%cf���&�6�����m�=m8z�/Wy�!u���͗�;Z7�g7nQ��89��:�6��2�mp�ӻ�y�9��x�۩v�:@�r���H���K���R�gs��]s<�8�%�[��wWX.��W	t�8� uq�1�
��m����W������g�m�lQ��5�%�U۵b�5�8ν�r�d.���ΏLύ��óE�a�k[�mۮ6��u��ۅ���=�7��^��r���v�/m��/�R�\[��jh��l��G�N��ӵ[�Hݷc6�ɹt=�k�������6�u��V;E�e��3�d�{d�֍�d�D�ڵY�C�3؅ݮ����g���T�%{K�xL4����]g�:��}kwS�1��kv��ۛ]V�ui�htw-��^.V���;kx�9�v�{u۸6뭼�X��nʁ�ug��0�a�;ru�8ۖu[\�j���xv�۔(���Z�ݹ�S7�8���X��1�;p�:r�Eu��uӈB獣q��̩�;��}��x.x7�=v�s�ֱ���[8�vںDm��	@�`�;!�ܳ"�o{��k�__i��[}�l���6ym�u�m�w.�t[I���<m�y���Xz6�!fٍ��Z�c���/O:���V�o-�ݢ�)��.��p@\������mr��<����M�ͪ���Y�8��.�!m��7e�J�������M����k�y^y��W��ƺ�s�Dӽ d�N"����˫&�mθ�w.��؇M�jnBn=�!��񱃰v����]{��S���a��r����۴��c��8K�m�F���̪����-v�fc����-�vcr�S�4��KA������s��C�G=X��2��H�6�s��ۮ���W[����y ����V�Z�:���;sb��Jhxm�wr]^U�X�@�e5ٺ��[nBZ��7��G�/'(sa��;u�rO	qvF���,����e�y.0�
Q����5�Z��J�s��CS�ʯ.���]�:��H�ɦ�b�.b޽��
^�ˇ[-�6,n]����>�t��gݼ�������oL��پ�n@:k��:��P85���u��`��.������ǎ5s�f"�v�b�,�n��n���]n7n�x�A
������3��t�%rGj�)�Lh�<�T���eq��7Qٸ�xrm��ʯm���Ȯ�L�pW
����lt�s���`r�E��ʋ���s���^3\9R69|��� �m{��.z�Wu�\����KV�ѵym��{{y.q���h���Gr��q��������!κon
���6����T���n�7+��w���sTK��Lq��޾����|���}������e�m���J9㣨H$�ˢ�A�"vwd]'Aݝe�'t�n������V���օs5���q�ݝdGu��gt��E�qS�VgM���ɶ��M���8�"�]���!�w��yv�$��eagۋ3�;������=�X]�Eͪl�v!�Kk;����ՙݶ㢴�6�r]	M��;2m�\Qpq�[h�ʲ�4�쬃�kQ��j�(�;���	.�:8�(���+���e�'N���qY~]^q�i�twG^�[k��(�����;�ٮ�(�89�Ae�7%o�;�#�,�����;�^x�wf�O�]����{�>}�|���ݷ���Nɰ�jb��@b��E�;��[n*�^z&8 u[(m�v��&��������ō���@�d�,q�F봱.�J��:�v��v��(cn�	�8,�
��r�`ٓs�<늜ݧ���b6�"��8�g�n�c�np���={K�EY{v�sݼ�K�5czl����;&2�����x�i]���۩̽���:�:��糵Ɍ��ڼ���m�[�9�$u�m���gvϮM_~_9}1��=Ӹ�WF:n4G�'����;WVN:��7�m���r5�;�	q���9�{�\�g9�ntY��LzbM�4eI{�c�n��5ˍ��ٍ�=hq4{Dwmk�x���r-��YWq�4qٮ�ŕ�zZ���n7,��7����j�Ŕ-T�3���c�:�wș�U"q���Swm�Q�hLݳ�M�q���ݭI�W�*��4u���՘����U��ǜ<�N���!v6y�z�71�J��d뇷+��Ki9�6���96*�f�C@n�2uײ9D�ݞ�,$X���kc��a�բ൶�<޴���U��qs�㶧<n�[��״9�rpt����Z�<6ٱŲk"�.#�� �l1���,OD��:��ݙ|�#��y��튶��ָt����A_��H4���#(l�_{����ש�÷<�N�n�N�[�\]�սk�1��k�m����Q��8�3�	2��+�C�mP��fQ56�t	v�Y�
p�����k��N��K��n:��算��������<z6��;��:�U�]�¤�u�x�M��Xy��ܛ�������>�n�KG<t�شn8���v�1���:3u\>��n��<�\���u���D5����\�۫:8��n�n��uCڮ������l��N�8���>�CWd���<���+��>`�t��S��Y%����h!{dW�m���ٳ��{׽�޴�s�����vq��<�s�E�¹p#��;�ceM�p�gp��u��������^��/f��@l<����_/l��a�T�r��;
)����Ǵ��l��������6NKY�M��=�=���מ^\�o7����sm{hk�y{׶�{ն���o-����^<�3��;�4
@#Q ��_���_�P��p��MW7̙E���㘠�7��.S���u/^_����)CC�y��d��`�t�gu��l�,����U��� �6E��UqfVŧV������|H���4f*f���Y$��n�M�Umo��4�fIJ����߻5���3k��)l�]�c��;z���m	T,��@�udX%�r��[�N�zV�>�yal�d���2r`�32b+0���$uf���\�s�<�T� Ou�ThP�~�ZJL*)o����A�>ӏ�彵��LOVD�%��W>�sٽ��ewY�1�HcR���9dma���,�w����%�r�"eFMh����Zo���}5���[z�KAl\����y�-�L����Lw�e�b�����]I��Ԥ[���1�1���R����^t%^Ή��q(Y3�M4k�T��ʖ��x�On�Ē	�Y�H�Y�0�NU>ET
]�����ș�
�*I�ޜКys�ϱ-/f�bY��ȭ��_���#�ug,�H���Dp�Z�����Z׻�fsM�}3PA���Ă{�ث§jd��m��\T�+F|l`�VEa�j���e*7�WX��t�B�p	�ݘ	'����Qq�tN�<f�����M$��=���>w��̘�8,�?��QX3�F펐�S<��C�c�H��ϓsz�6��߱,m���
So	���;�������6ŝ�����^��KM���d��;:�VΟ/v^��	� w;�d��#N�o{�s�d���^���H4X�f��Rw���u�'�e�X����G�N�2D1�X��1�� 
]�z��� ���y4����u�]☏�fqV-`pߡ��e�b�z�k�巃<O��ذQf=�7ꈢDP��]Ҫ\ۘ]=����a;��	�wb�$��r�h���뾞@��Ow0���$D�L����9ъ���X��^�3I�Zr7���T+}�Ѽy>�{���7�ɹ��q̺�Ury�p �9�i}�[A�t��/NzR��%-���9���:������X	�wB��:�~4����ŏי0�/7�m�W|�Bv��Y�6,�t:����QQ
넬�Wh���/��͑e���n����ƎEWUv�@�:]�JH㤪��մ��oޚ�4�h����^�v_{yӱ`�
�7b���S�Pʭj��7�9��u�c榧��� �'6l�Oe��8-�SH�w�}�>Ck���i�,A�=ڛ��v�pV�ӹ*rӖ��J>�M�syZ�(�{���M�ߨMy%PW�M��m/[�-|ߏ3�>��V04�*�ٗ�FM�\�謻$gt݈��_+�yBc`��p� �R&d������mD<��J[;��=�۲q�d�+����r�I�����Lԉ���+�yX�I=�l�$�_,�Z��[{��%b� ���/����yW����0l��m�6��}N�S�w{A	 ��XE�z�`'�U���*_��B}w,�/.ŋ8�~�E��f��{2��64��c	$�s� ��s�����kjǤ���G���5��K��Iyӷ �cY�$�w;���	��[_��,�!Y"Y�$E
h�S�����Y��F6/����8C���?�{��C���ދ���좯6!ׯH-nk��(�Hm�]�):jX�W�*���o1�6_�<�}���;v�2��G�L=
��$0l����td�sm8��^�틥�c�OZ�y�q��\;;/s�s{]<�v�y��ۙ�0T�K�x<S]���<s�oXy�I�W���˶`6�z�ð���瞥�Ƚ�	�98�l�l����H��:����Nu�8��W�m %��9b�R�@Ḵ����Z�k�"s��s�ᛧ������RY=��iݹ�͒���S��ƅd�W]q�8ܸh�gy{t�Lv�,-[gvހ�:z���"����*]����wᔊ�����!��˞y�> ����gs$����v ���s1;�w�2K!\,��gޛ斓`�%��:�n�Oh�Iu�� $�]w��{�Y-]L��;]5pA���+3	��}�Po�R }�2��3rA�D���e�AY�0�K]v,=VÒnr�Ԏ�'��y�.6��w�H'�����J�	$�)w0]AXg���\�=��ϛε�f��-T�K���d>r�%!�])�^Z|H�z�	��� �w������լ}G�K��{c���u��5��\��Ӟ��F��Ok9�X4��>�;ݾD#��*���y���şs��B��o�6g$ܡ�{���$�뱦���|�U���>�s�Z��\��3�R�i�az��Φ��X��@�VB�湷�Ճw=;�[���שfz(�N&��gF��t���/��w���n�_�$�*�{Y�q6L���j�׻�$���k��^ii6�7��	��b?P)ޑ�OW�`U=�|�=��|4�<��815k�OS�۝ߙ�n��L� �%B���7�I�r��9����T�5R+����o��5xrzv���{�&o��MI F�ذH$�Ҭ@>$:�Y�;C��a�כa�*�R6⌶!3���[}�����=϶m�I뮮�a��k_;�����+mP���ز	\�X@ ��r��#x\��<.��U* 
�z����V��Z�U]fc�/;�b�N��9}5��]u�$�ʑ�I>u��	U��z�kko����*2�-b>{s�h<^��|�G2����R�Ht��{22R�YG�	�@�c�y0��P)��]�$�j�i�3�i�Y�wջMs�hj
��+�+'x�6��{8֛�׹��W��~d��e���n���%�]�Z��� �낐�x3ďoWX�e���D���l�1���0�UsѱB�粕 ��9�.�lK�bz��IV�3��ʺŝ�ќ�Dޓ�q��T�@J�q����z������nG��1��.s@2�؀�~��m��v;6A3P�s�n�=W�	�]b�q�sƛkL�Z'��G�ػ[����{,�$��ʬ���K7������cz��	�O�[Y�$<�œ�Q�竰�m�E�L��֯�kR����O������]�j���`٬�F�I��0-u�c�4DMQ�`�l�{]x�of H�n�`���R]T*��W"�Zz�]"ܵ�G�d���C�+����"^[�����qg.:VLz�
u,�ۓ^kC�GauI٠�UZ���f,=Sw}�$0MJ{�	��H�u�IT��z��6��vf��fᱛ2{',}U��0���	� �9�|^�5�o�S�D'���ϥrڣu�ϯm۾��{ݯm&;o�^�G*MB(�I%Q��oɇ���Z5�����I�}^�������$б�<7�,���9D�"f���:B4��r�v`I�V8�O��~&��[F�ǜ����9x�G�~�ڞ�p$%rUdzF��-|�o���!�I����MC!v[�I����Fs�5Ręv�MQ��E�<��)��Q �j��ܫH��O��T{P��es`�&����B��X/0&�|�����}ΌP4���8�Y>!5:E�G[��.@�����NY�˓��b�]��إn�����[�ᪧ���I��D��\��v����
j��p��ٱ�Ry��Z�����0�/Ī;j�����u��;Zb�X�3��q������]�v�uN���Ol�9���;![�K��Tm�Z���[�݃��k��Zv��x���<�4s�۬�zx��C���;ybA�n�ڎ�O>_v��v��X��gR���k�`ix ��/�js��u\Ol�㵊��ݷ9�϶:Z;h�Uc�:q+r�ӷk�۶����u��a�{@F��8:�J����Y;n#7Yc�ȄH82�b,��}���Um�����,_�$�9ۏu�����V�-�uu�a$��N\$ƲD�F"",��"��M��T�>�`�A v��d�Gc���6.�H�v�T�6�S8�C����}��������6ؠ(4��y�7�	ɟ*������M��﷘�َ?G��*�7yꮴr�9�Έ�'�g�\	�!c{�H$S]ct<��{�u])�OKu~34Ęv�MQ��E��[��k��K�Y����$@x�s>&���w�*�жg����\��!ɞ9y��,�����.:8��ix1�eB<�$$�q���>�<���k+����s+�H&��y^㺅�y�gǱ��'�4ߢ��
�����7�X���~�{�-���T���^�څsە��4�N���ܶ;���ʃWM%��	���V��9��V(U���\҇X�n�4��õn.fqWA �nsY�k�W��L%�rsyu���D���1B��@��w����/đ"󳫚�V��|��$��X�zP!H�jh�fj3�{\���r��Lx�+� �I����<�ʹ�p+6��l�[�)�c�"�D�TUI��~���d%�W�eTr��;��H�癄�s�O����V{]F�dZ��k����Hi��5ah��\p��5֑�jH;��^-O9��9Z<�����ɝ�k��G�/�m�a�[΅�H �m�zpwe�y�x�f��h�): �����3Ub,���'��y����&[�H$x����_!��3mm�w{ߥ
�� �fo~�-&��y���?��&O:Ɨ�B�25�a���cA0M�)�2�f��,�cjf���C��Q��Db/E���z2e�+������T8��p��8v*��n�����S����ϴtǛ�G
O�}����z]%���ջJly���Q��٤�Vt��6=��Qt��^�^l��Bۤ�bH)UN�(D!p���SMV�a�u{���د,u��V!�����h�mR&�em��q�S4��ي���*�P��F�7�]�mB
�K-o^Ő�3��Τ$�j�s����u{.�i⺶Q�sStze>)ζ�.�l�Ti�r�o�O���Ԯ��hּ�٣Q���W�������İD��;�v���WR j^fv�By����̠��L�e[�h<jA�%\���6*�aɽCB�
�_5����m]��zI���j�
B��TE<�%ގ5�J�$����=�,��Rv�G�ڦ1��2�*��3i���f�<Ó 5�ћ���>��J��qeY���A$��H�yrgu��+z����h�es�Uͬ<^.�@�;-n���Y��]M[Wx��캼MQX�փ��aܺU,�g*ak�Ӆn���l���YZOL�Y�뻔Ӝy�5� 6G�ɰՓ4_>��)ɽ�%�¡<{�VȺ��a31t,��P�x�x�gV�eo$�Y}��R���5ܭL.�[�9��l�C�<'D��p�9�mHlcN�0�9��Uf�]ۘ]]*��;�7$Ȭ��=��f}�f$�ܭ|���y�t9��-fua��b�V�P�u�컝�gG�'�i�wv�""��[q6ˣ.;8�8�Z��t'qНE\%�]�p/����gq�k��Ύ����Z�N�.-�\|����f��H]�k,�+#��{vK���Օ���W��@�D����6�E�w���n�n����:r#�2����%tGG�REy��ڲ���c��t�W���p��"".)8�q�*��v�Hy�m���|י^u��yו|��3�V����[��\���7qEH��Kk"���N輬���_.��3���ݒv��gq�k���:��(���Y�u�ky�ZtOϿ�}��T��`�Ŏ���O��g���SUB�����������в@$��b�>uܳMveFR��'I!v���2x�l5"������m'���,�D�.֬����0�ӡ`�G5�d__,�k�gֵ�D���(�o��YZ��)d[�Z�iq��OG3nNBy�R�E�:�ԯy�v���W�G���/����  ���n�fM=r�l+�łI;��*m�11�T*s	�-���iЈ�ϔ�:]�9v���H����I/��0�-�B��iu&��[l�c�n��}��6�9��0�4ݥ=��hwm~��»;���*��NU�=�P?]���ѳr	�u_�����-u��0�BmOW"_�-ٹ[i����c'W.p{u�j�����)�s0��
�E��(o&����0݉ͱ4�N��� o��
�:�[@]��P6��$ή�~1������ځ"/���$��na$�*�N�Z!�x^\tV���*���U� H'H� ���pq�������*`�(�
�;����;>�KNy;����A����IˬYfg)�n83COg�t�M�y��x�fX�-��,�k�e�Ќ��)nu��0��|�?����Je2g�vs�9�ԧ׾�0�1�����1z6�X{}�Y�i!EP�~�GE�(�$7�;�����׬��
N�� S*'�߹�m�) �Q}�k"��]�n߿���������6���_�Y��u�˰���G�È��O��jͳl��@�J@���Ф�L
�O��o0/��w���x;����{���`SF��z[��pb�����i9��Y�2�Je��ﱼ�d�9��÷��6L!Ĕ{<ޡ�aL(aH��g"�B�Q��Q������g�� �����9L��R"����n���!p�SN����ެLǃp8/i��h�n
O\�3	���i��<j�k->���Cw�9mm���*�A�iR+B��*lN8)S�"uێ�a�����=��Νr���sn��]��/\��۱ΠN`��5���Ӝcwmn���R'�����{q�O��&;Fp�WL�T�t��&������dx.2���f��ϬR�2s�n4=>�/��Pq����%�C�5ʫ�����qc�bx�˗��[k<�����<��]Q$u�p�ەŋ���{m�^EE���ٜt>x��
ڞ��0���x��r(8TRJ%m���g:���@�4�k�߲v����U�w���RAh��{��&����:�5��]��g��y�m �l��!�}��(i%0�c�;f꒰�]��P��)���2ZAI[ϫ=/�n���������4��%0*% V}��РhJ`Ti ��q���tA�!^Ѿ>Y�Φ`Ox^>��0�>G�jKW�/V.��BK�~�E4 RAH/��7��P�IL;���wWo��^���C�aL(aH�~�E&��C)��S��̚K@��}����/]�j�[i-�?��w����>�;�!�L���.��_��_�����]mk�ӫ7�s�@��@��
e	�o��6Ϲ�����k�L��HR�wY��Eo��
�X.�pb�B�i�=���!���P�$��0޽�2lf��;���/ޯ��(�(��Ф���O9�o05�B�}�{���
�z��]��ѿ|�V0qV�X�JE��ݳ/e�� .���v�݋$�D�������m`ض����wzȦ�
eFJH.��o&�KB�R��W����m ���;�w��������6�����Rh�Je2P�{��y�BZ�zUk�l�c�V�@Д�X׻���M$91���#��Վ�B�����mI��۬�]��ap�Uiә��a���i�N,j� �t�7���W�M�iߪ�H>�����o0)4 RAe'����6����Q��~���1�s�4��_8Q���J�1xŹ��laN��s!���P�$�
a�����6�L�
J@޳�sy=���y޵�|)����Oy�o04]R��w0۱�N����-���p�.��BMc����Zu�u�>�}�>��A�u�0�֐P�%0��ﻨm��S
aI(O��k"��p��V�w��7��&FS%��������G�s����)A�1m��%0�}��v�R*��w�r:(����R�ث��4���S�I��IH�Og��0�6�I
�{���(hIL;�}�����c����\Gn�%��vyb��oC�7��7�����71��w��ӷX���j����aO;�{0)&�)%S��w&�m��)�� �9�ـ�x�>��M���G^_[M=���0) ���w0۸���������V)kޠm7{�޲)�
e��gf�x�ƴ���-�X�N�ZRAa����a�TaHw^�E&�)��L�����������X�d�5H�}gSr��Fb�%����}��$��P������7}�fg�(ԩ�;s$R2jAlŕ/��3n�*�w�����p�iK��ݚ�ժ#�/(ܑ`�N���U��j���m黨�����>x�c����ٶJe2R��g"��JaW���]%Lc�P���:�9����T6�/G��x�¾oli�d��@���D����(J`P����W�%K��k�Ȼ��x�������巴��ź�7bd���CP)4$�s��)�
e2S)����s0)�����&P�S{��0���0���g��%$Ѕ2S)��N���_}�5Kҗ�}��yf�B�vOLn�[mYl�+���tv����N�Ua�1xw�o���w�c.�X��_� y)�~﷐۶$(���>�IAD)���~�7�` #��Oz�`�� i�;��m�d�P�HRϳ씆�S
���7wV8�U�ZA{�����������/�1�>�x������a�O�)��
1����Xi�Q�~�7��������㷶��gw�f|0)�}��������|��5��k�����-e��-��B����M��BĴ-жVq9��z��5��Yk}��m�͡l,mII�}�䤚�IHRJB����a��a%���U��UV+�֋I�ؖ�y�=�3;�o�xj�����w}�M3Pm%�wD����rV���ܢZ�����7�iM�hZ\BжX'�����������e_�������`�:c2;�� l)��dwے��pn,67�A�1�����Հ�5[�9殶;h���y�g8\k�!�xhZ����g%!��-����ٻ���q�V��m�-ξ�2v�Yt���{��^���tZ޳_v/q�G���Z֊II����m%��o�}��Cf(��]л�{����x�з[���������IMR��q+a�	&;f�F!{`�{pt�=���xk?���>���,��W�������%'�-e��-��B���o&�m!bZ���l,>�����pmag���o�i'��oY�I5.��Sq���e�w��a��a%����n�8ŗx�P��I�ؖ��﹞!���6���ǝ�~�9�~֯�i5�g9+Eл�KB���o�gz�д؅�i)
e������ghZJB��]o��f����R��g%$�)�+��k|��V8�U�����=���!��$��Ir]��ﳷ��Kle��)%&��g��կ�W����BZKe���X�����Ca�%�I)
������8�����ƠRR���|��5�k���Ҥu���}����C�a����)�y�d�6�����ih[����q0�hZJB�]џ}�䤘������e%6�Im����=�m6�Iigy]ߖ�c�kE���^���������Z]�=�9�I)
Ӫ��c�h��X�:�RR��w���i���ihZˉ�o�g�q�e�l�Z�Ĵ���rRKB�s[}���j��L�N��|.jiBy8�|���ӱTh�ٽy�d�w�z���L<D�U�c���'�\�g)I>b"�GY<0�Ђ^^�h>w����2�9S�11�¸�Z��A<<lg�XB5ݨ9S7���_���ێ²�n	Q�<�7=��\nnw(B��8�6����^��a�7Wr�
�9�����sۏ;�a;�s�[&�1�����݋�x�n-���q���X���[8	����\Ib��(�W:�m��B���#�&����f�`�*�r���v3s���][\vL���#����1�x깮٠rj�d�>;�?;r����h��[�ib�@z��_}��G�t^`�h|��6��ױ̆�0����.��{������$��ZKB�R{_g9)%&�����|{����g�{��a�7�%�WD�-�;���������}ź�)9Jڕ�ϖ�Q����ZЂ=>G�@���[�y;��q���ǲu�CZZ���l,�����a�ж6�������rRM]��'�G����*VEʃ�~���m�i���oY�:�k	��}�Q����s<Ci)�IhYtKOo��JԢZ����Z�x�a���=�^u���������-e�����8�2жX�B�R{g9)	h[(����N�A�\3m*�[N4���_i)�"�e�g:/_8�`�H��'���;x�$��i-,KIi}�5���BZKe���X��w�6�U�8�3�S����M!I)
����}�!Ĕ�<߽��%-QKϐ��_~ߵ�!��)%!L�-~���a�-����ٳ~α�д6%�l/����JB�pmIwG}�g%$��ZJle��WΕ�aH����A�um���f�n�5����㶐;OjY�jM{�ݯ{}o��=�n�ĒU�K8��h�*��Q���棆���<g�Ke��Ф���3����h]�KB�R��w<�6���)9�~�:��8��hi���o���8�B�l�-KN��g%!��-���;g)e�1tj����o��9��t�Dz}0���g�������Sz�Y+iƍE�SD9��_L��$*�Iw.ڣO��e�u�G�s�E����>��RP������$;��$aJ��7Xm��j�u��~ay�go�q%��IibZKK>�5���Ii-�Il�6���s��b�hU�KB����^0����mq�c�ϳ�:�Z��o�uw�q�Z�д���s�����q����h[�}���f�����ih[���u���cz�o=�$�)%!I=tw��rRJB�S�ZKle��q��mm��ѩ�l��bu��:��4���o;gq�f��MRL�i-�D�Ƿ��KB�Z������P��Bд�-a�}��hm�w���}U��i�l�-KMgZ�JCBZ�����뎠n���-�ҏ��}�iI�t���[{��v�gZ�W���|]]rq%��i-3�g9)%&����m%���s�w0���Z����}���<��3��5W5��m��{����[���w."�n�l]&PF��ɹ����C_��}}�&�Y���v;���Zo��rRhBж[-e��-߾�rlf�����q-a�}�ސ4� d�'��]?l2� iɀ��g%$�t������;���I�L$��+���E�a�VKI��[���4�A�H��,B�TN����w��҉h]�-IHSg���P���Z���l�>���x��Z�>��6�FܭN��v�~7��+�۱m-aw�z��R�m�	�Cl7B���s!��IwAi.]���w���q%����%���8�Ռ}���L��b�j��5)�s��A{��@�Z� �)�f����t�=[�&Lť�nP�j��p���s����i-�IhS�{�4��Q-
��Zu���<C�#B�8k�i��I~v���J5��k=��!�g�~�󃗍&/`��q����h[�kd�f��%�i)
a��s�6Í�l.6������Ʋ)��c�7��4������-����M��KL�^j�Q���]-��KM�l=����Z���tKO{��GTKB��~ֈ��l-l�w��B�qB��-e���{�!Ĕ�3�-BĴ�:���IO�gb�gUd�_Y���{y��@��}xn��M��Ǉ��L'NE���\]�}=m��t�����+}�c����K�Ai.�-�>�{����Kle���������E%&�-%�w��[�~Y]�M3q���9�m��ZtKB�s�������m�ۭ�U�b����)������E5�-%!L��Y�[ǫ�iߵ���6�����ih[�}��q%!L86������Ȥ�)%:i-�w�f�3}��n���qDzH��#g�]�X���ZM���o~���9$�X�KB�i����tQ-IHSl-u�Wϝ����w�wX����uN�Z�!h[->���x��Z�e�h\KM��k"����;f�)fbMQ#�@��ն*x3~��]W|kǴ�Rz]��)�3����g[l���$�߽��RRi-%�I)?od_SI��Q�~��J��Z���,ʨ�%m�W�خ�e�C$U��tRqIB��/Y�`��(�Վ��7lO���Q��7�I�E���"�_TY��P���j�@E�$	(g�.f&kƨ�Va�-%%��g"�Bд��2��@��um����(�ۛ���X-@���0ν�ghm��h[mIwF��Ȥ�t��#-%�O��o0�m��ѧž���k9������vҰ�c�ݟ7B���D>�Yk�U�luº��o������sux�QkI��[��s<g�-��KB�i�{��h]�-IHQ���� I@�;4�9&C��s��8�3�1�o��ghZJB����ﱬ��h[�������n�wY��m�o��>�m�Ip�I[q��9��8��a��}���Jz�Iiii-,�}�hRRj%��X�Ke������i)
ܢZ�y�x�����V��mڿ��A��;`航��T'oP�6�BӾ�5�MZ���X�B���o&ٴ0��hZ%�l/籎�7����ϸ��|6����-%���k"����閒�n��o0�lL$���:&���V7��m6��{�=�38��������I�m�����-7�c9J%�i)
IHS{�s�ChZn!hZ\BжX'��>�Gǈϭ8O������ �DI~��C@�����x��v�+wV^&���h[���d7���Ai.�-��u�GȏIKE��K^dzȢ$���{�օ%&�-%���[,}���a�7�%�VQ-a�ϳ�6�$�{���韢�n~�V!���S�]D��s�#]����n�����i����8M���������h=��IVmP�0��z7��C��{�n��:z����Y#,�wϖT��h �V��.P$n`�b������2�A�K��gVJj�6����r1'ͩf�U$8����Ĺ}ݻ��}�%���y�6t�slV�aVn[ƒ�r*:q�V|�Jラ`��!*�%_�����PY�	�e^�ܓ3`�4vW��3����C8W�+.��j�:��얄�㣬�s7n��<��'3�P��2:�zS.U+Ӱ��qj5ɗǻ��,��+]za'���ڧW�[��KU����D����.�P��4[���o�]\�����砙x��9��}��\��tQ��"��G1��L��P�$w͌�A�����Z/��-��d#�Ou��i-+��U�|=�F)���ed���lwm��*�p7^��wE?5��H��|=��\�lw3c0��Ҋ��UcLBnP�	Ғ�S��vjk�(���k���ggqt�XȻ���]��,쎲��|t�پ6��1�O�Խ�(KWsW�2���Ŷ��ն��f5���S�H�:oZ����6�����5[b��iK�l�mЫ.�Ǆ`�����Ƹ���(cvF.�YC��Ʊ�	V���.��{i�gf(�����_| ��U`I�	�LKK����lW>�{3rKx)[#M���G�A�R h�-9�/{;�gc�qÎb��s�g ,U@U��LG�K�I\t�%|�.��$C�[�����pqN%�vI��ھ�IIӾ����^[�E���k|9���������:.�ҥ;���Y�'ev��圯�we^i'Q9�\W�-kY�rE����:����|�mGM���7���o�hr��{7m��Z����y�J6��{��:#��޶Ok�b)�s��7AE��dr\G^efu�j.N�

"/4"�m��qm�:�����ٵ�g^��*���)�:s+�����B�:K��w�q'^YM-�e��v�IPֲ��mѥ�v{k4��jN#���z����e���V�޽���}���M3�:��{q���- [X��Y�o1�k:���н\ʺι�K�%�:v3d��J����3��'=�^�9��m�f}�C��Pq��9>������I�{��o�z��[�]���=�ӭ�x�Uv��nc]4�ݮGe%�{=�Hc���uz��h=�i9t�[�L�����An�vNܹ���v6���������n�9�3nn(9x�OnN�{�W1�m���;�Fӕt��=e�Nvv�<;���Fݺ�Housr,\fM���{N�6&9�`�r�$��[M��b��X�DM��p�շ�C��V{'Ic������O�[��z0����O/�kls.���q��Vc���&Mɭ�E�T�خ�m�"�G��s�Gbה��|�W+���V��mT�q��b��HS��V�m�;h�dȮ3�����]���N;;��I5����ն� ����u�e9��6����k��^֔�t�[Ő�������Ms�:�vtj㎦ewcqE�qq�F\8٩f�)�r&{cv�5���'K�8���\9���reŢ5��cɼ�c\/q�������& s�c�<���>K[hwi�<N6�;Wq�f��@<tۭ���G���n(���y���o.�057�m�g�ӷq�;��H�w�����}��7���m���[m��;҆�*s\�غ�#�9���ջi�ègӑ��Gn�9ڐ��L<s��<�\�@���M�9����Ŷ���ީ}��hk����q�.wm���s����y�8�::W�l��u�#�N�� n�=�g�����ۻ&�e��ת�^.<�4���v�:�v7Fg���ڍҍ����q��r�
fK/Snr��y�C�'6�N���8ڳ�Yϛ�ۘٹ�krm �v��p޷�����ss�Vp۶�6� g^�����d���[)[.⫱v�豺�	��Z���8mث�ًUȞt���:b�q��q���Az�̻��*۩��Yݮ���iy���=��tV�;��Y��u��dݫ�G��k����]x��5m�{<W�Y�Cu�gv��2*Q���l�COM��������¹�ú=ںx�V��z��=y�ٽ��)
�K�SPqs���7b&��b�pZ|�ۉ����jۢ�:�'n�Hl/���3u�;�� �(Y�sc��ʥj��D�7}f[6�9{sA'�װ2"g�!K$���t�<��;�C�gqg��q��1�{ǩ�]���*��uO�!i�{Ȧ��-�2жX�B���o0���д--ag�{�k�q%!L>�y��Cvs������H�	�$�B��oy�o0���{���c(m��KZѴ�M�����3�px��q���4;��n�>5~�����s��Q-��hZJB����a�-6!hZJB�b{�s��3�-IHR���SMo8��>���E%!L6Q��o/�L,�m��i߹}���ҭ}i)
aϽϳ�6��2�Z��a�gx��{����%&��[.6�Ч�}��Cd�Ы(���C�{�g�q ������)]��|��5�k���dSy�U_��>Ͻ�����Z˃-{��f��JB����������a�6������^�Ȥ���:e_T+�l#�xI�'�o쭿M����/��Ԕ]Y��ZM&�[���x�[.6�в薚���GTKB���|��<��f���-���-�{�桴-6��ihZˉ�}ϳ�8���q���`�����E%����_�/�d����*���H��2}!�;��3�VK��į<�%)oձK1ʤ`�+�<�u�T�m�x��:�͡n��s0��wAi.]��}ϳ���Km��Ф���}�hRR��z�V���o)-�m�y��Cx�ZtKB�{�s�����s���|����UjB�b����E4��i)
f;���_s+Y�ho�1����C�`�N*�xWV$����R�q��g��I�F�<�vF7*��\`�n�u�T�q@��Ѝ�޳5�I?JCs�}�iC𖅡q-a}��w\C�8���д�]��5�I��-%62�[�s��_�>���o�cy�д��ƾ�1�P���%-d�L'"[s�s<g#Ė�Ih\�%���g"�����:ah[�s�}�y��q~�>B�����h[,Nw��x��Z���--5ﱬ��(�Q!{��%��!�iG��v�����!����}��͡ԗt�ˠ�w]�;x�$��-%��-%���s��RhKIl����m�;��B������{N+�����T5�o��x�4����boh��:[\ϐ��[iF���9)5�-�2ж\e�n��7�pf�������=�9�|eIHS���;Cl>mam�i.�׾�rRM]���i-��������	-;�{����u8�o�O���3i�)mr&(�h���I�n�o0���z�j��DNZ�J%m�ͦ�gF�0�Ť�xKa���g��Ėˍ��,.�i����Q-��h[q��l���xiH��$��v�J�$�&�[>L{��<C��-e��-%&���%!�-a^����i��L�a���c������Ai1���W=��]
a�w�ghm%<i-.%���]����Ri-%��IhS�w�4��D�*�%�~���w:���o?!��#J?�[V9��ݪ��Xҍo�j���JIHS4�-�2з�}���6������)�$�5{�~���w����4���keq�y�J��U5�V�.�jcKy��h�6��җvf�����n�˽ЩL��m��:�7�l��������C��ж���^�s��j]���ZKm���w�m6&�Z^s��x�,Kj�ZѴ�M�l=�}��Ӽ����s	:���.]���s��R��h[l-no�o0�M��������{���%�y�;Z����<�,�e2�q�.R�߇UN�h�s��Ú�q��G����� �Ĳ�K诲;ғRJO���%$���m��[o{��CstKB��Zu���<C�Z��<�����-ۦ�"Z�e5T���y��l2��&���`�(��"cQ���V�\ufo�o���T�����_w�ִ��4�e�жX�B����CHn%�hX������s�6Í�l9�;�ư��p�5�k9)&�����e���o���M�m%��J^_�ӊ�p�E���������Jg[Ih^��{��]��3�w����9�]
%�wD�-��ж���Ci)
IHS7��{�!�q����Z�~��N's�g%!֣J?�S�x����#Km|4�������K�IwAl9�w����Im��Z���x�^�	��\c���}�����$�tm%���}����tKB�(�������hm�0�-�p�ғ��ݪ�|�ҍo�j�ZC]��#a]���$�O��'��� I��pf��%�hX����}��\C�)
a�mIeѯ}�䤜����~J�
��Z�x�f�B�Z��өZ@ڃ�ea�YA����C�&|�I���㒍��z��p8K
�+�������>����V~�	
�IO�-%�2���;�m6�Ii�ﵜ^0QmU�+Y4�S{�o;g��Ke��Z.�i���rV����>�����{�I�:텡m�^�چд����h[,N���<C���B�c-BĴ׾�rRKB�w?k���w�ͭ�EE�1V�ϟ̒�S��+��vN-3�xB���o�mn����?'�#����w~������ǲ���]���������g[c-%��ZKK׾ִRJM%��oY��ox~�~�=�>�N�����}�m��Zr�h]��_sv��A
��H:TLH����!����u�����j2жV��w7�~��fз{�>��͡�.%�i)
ag;��\C�86���д�����JI�����-%����w���|�-��˭{�_F�+����������m-���}�3�Ė�m%�e�-5߳�����J%�i)
w��y�UO
�1�a��Bд�-e�����q�h[-���`�����JCIQ��������+�F���i;kl��T:���_�& �= M��u��oĖ�2�Z���ߵ��������\}��y��λ�g6N![�Z����������m���kJNHJ�v���J5��j�ZT���i����h[�����͡�5f5�_��zm
BĴ-��Ͼ���R����.�{��JIHRJt�IhS���4���uzϚ�j}�Ug�+�������M���Ԩ�%5��u�K)�i���f�_\*&\��UN���l饱ӷ(+�7?<=�x��?�s���vx,�\��<�]��G�.�|����ۂ�ma|�6�c���#��<��7&qlm����&�#dv���Ƶu�{A��9�<���=��׳v�%��2v8���j���vϔܻŸ��2ua^{'Y�;�i秶���v�	rZ�����E�8nT���t��YN�û=�*��s%�m�[;�`�g��#6�.9��αn:t��6-�ku�{n�#�S�Nc��18�`ۧFƚ%s��r�����F�_�g�c_V�D�s��x�[-�����^�s��D�-%!M��-�{��B�pBд����mgA�6������>��-�2д--5���JCIh[�G�L�J?��q��z�Im= Q��$�U�q�>�����$��ZKK�Zkﳜ���BZKe���`����6��(��XQ-��t�x}w�l��zq�0��f&��[Y�!��O}�g%$�)%!L�-w������BĴ-зó�ę	�7})M>��$�A
IwG��g%$�)%:����o�}�a��L���a~�/��ݦ1��m6	l7�s�����s���)�m%�I)7�g9)%!Z�Z��ж�=�oP�M�hZX��l����s�8�S���׽��حn�7�8���2%���5�4��ҏ��������6�ch[�_9��v�R]�ZJA����JȏI�쉶6_D�#�F������JII�-%��Il��z���ha%![(��ܨ{��s�8�aQ�|�s�2�*��j����1_pi;p �7��x�<[���f���Y��w�~v����*��P������JMD-e�-e�Z����m�C(X���dIO������FH|)v�����I�tc��rRMB�-%6�Im���N�_-��_oZ��,�����ًmL&��w����8�%���Z9��{G�E~0JL˕��[��y���T���t+e�U�⽂΍�M��e�Gj[��u2�UQ��4K9Y�=�=!7�m;��9+�л�Z�B�?~���C	�-K-e��߻��3�-e�-C��<w����㉿oz�[j4��C��q4qPnKl���ch[�_�fC	7.��]�[�n�z
>�=$#�G��2�ͻ�5���RJN�ZKe���m���y���JB�(������hm�B�5�5�����BQ��[k�߹�i{7����M�]�����Y��B�l�-�o�ɱ�C(X���ih[w��v��q�-������>�rRNۺ�{�h0��2�Z�W�s&�e%����Rb���I6�Ka���g��Ė}&H�� �Au݈��ʥA����m���HZJB���}�Cha%!I)
fӾ�{�!�r2д��$��>�r ��� I�v9�%2v�>�s �� T5ڙ�,�g��g6ԝ�:8�m��׉�Z؝���H�1����&1=h|���_^���v�R]�ZK.��{��������������9�I)4%��<�}�V�����w䖅=����Hp�Ы(���P��s�8�ah[~�%_n�mq�Z�д�����JN���>Ń�o�z��8�K��H@�KBд�-�������JB�q�-%ˣ��Y�I5t��i-k��>��.���?31����#�C�דdI��V���lKa���3�6�����$����䯊%�wD�-�����9�}�訵[�n쭉�S}���RҐoB�rpDMR���<�9c[5��%�݈���W��R�nх[V���$�s��C)�B�д-����s�6�2ж[-II��g9)	h[���6%p�P���w��l7з�Ͼ�k9��_;��]����{��v�g[l���%����=�h����i-��Ke����y����s�Wz%�X�KB�k>���<Zٯzmv��W�S�SZ�!������JN�-e��-�2зu��ɸ͡�5��;�0gF���h[�{��\C�86��������s��h�IM��I�}'�oo�H�F�j�.q��&���l
\:��h��a��a:��<pt��rbq���JI~_���޶� �\�f{~�=�o���_ �x�3.$���<����x�}'��Uh���X&����v,B������H�h�+�����o���� �����Ϝ�V�7�9ÇPs�>��f��*��X;U3�g�� ����$�מ2�+�����߾@ 3��z_ ���33A�)��FD���������u�WCU�d� /���K� @.��e� ���]�����ݡ}����\�*\�R��h g"�4�X�J��F��Z�T��\2h+�8��	��&z�i����LZ�����6�bc(F~xx{� T}舍wz���Ũ�b��,�ho�=�^�7����Y]0�mF��=��M~�<�(����-݈��pfX�S��
��8�չ��ǟ^�ĜΌQ�;v\�W�3d��cq�B��[FYϸ�[��krx����� 1�m� 5����R�ݢR�.��5^�0ogs3�z'���P�B���O�$���~>��
�����I ̘ۜ����s��� 5�kcy����+o4�Nj��Ƹ�<ox��M�v�	$����lT껳e�%�xs���}�o{_��DN@v��U��,�>�]�7����$�N��[$�j{۲BI'�;�X
��z���s�?oy�E�6�u�-�
ja��# B{ۘ u��m-�Y��:$�I�w�d�~$����{ҽ��CG�|c�G2�ee!z���c�
g�o׎�֎�)�ܻ��4_DU�������ea9*�K�4�M���i��v3���$�Lz⛫��#vcki��>6ś��Hv�,G����ݶ^.��j�;q�ш��j�Ɏ��p�%��\�c�;v��94�9�&Շ��E������ݛ��vj��;�8��P�����h#��9���4q���B���=��CX�c�lf�c��R��>+��Uq���)������{����
wk]��XNy�kc�T3��r��Q8���]����p��UC�/Q�1=��I�6ᰦ0�~�O���#��-�h����� �=�f��N�R�)��������mI>�ݒWuS��̼6A�o���  PZ�kݮ�MuF3y�I����$�G}�$ ��_���g.|=�3����&>�Q2uf#5�����{�^��6�i�n��3���M;ۭ�	4w�c��.O5�>':�W���cʯ���v'XH��� $��@"I$�n�����F�]�����{i�"m��R����zσϝ�f��ܞtO`��:f~�[$�I$k�` *$��m�nϵK���l��&욥���h��[��f�fR��m��h}�p��M���]
Yw�{�¸�J*�5<s|���`|�w�$I�ݏ �˧�w/I����% ׽������A��Y�|�ŧ�ˀ"1k���A�:�X*�vc`�������g�Oo*n�{��c���O���=/�����{�`�wB�^K���<����\i���+���|��3=��� =�������9�y�fgG�����{������֑e�FA�Xg=��@ �vs@ ��ä��g[��h$s����G�o[�j���	|0�"͌���};�b&�>9}"� ����6 ��^a� >ｾn^9�G�V����&&�"a�<lhq�R�kfzo2�������S.���s�|�`
� 9שՐ~$�{��	_������
�ٻ4.�u`MтS�vU��;׊�7<�{q��=t����9�����u��R����{5��� �{9��$��M���?m�����X	!����S=P��v�WɈ����{2���O9S����j�؈$�MR��Q ��6@!.K�X{�=^͇f ;��#"��`�K)�<s��Q�oݚؔH\��g�a�L��ͳ�Ͳ�L(��+
��cgthN���Ux�UԘy��"��y��W�����:�CM��ՒS�*�A�Z�.�-���A�\.��N������wf˼��
6Z*+|]�ײ�s��sRT��l9s@����-p��'_5�F��[��PV7�z�g���a헑���9��F���й}�s6ˬ��E���a]a"�TCH��Ѻ���WA˻7c
���[�\����$m�-z@X/z����/������+�~�|jq�W��� !)`�Lsw6�p[I]d���u�B/C6z��fb������i��5^L���ީ{�q�4�_Z�u���Y�`CF+d'��$���	�g	�uW;�;�
��Wz�o�U�|����\���Zk%��(>\��vʌ]�gsn��>}�(�͗2�[��ؚް�]]xc���z��X�&:ugX܇������̀^X�CsMډ�P&��Y���W���u�]A`�����F%��N�-���A���@q�9��9��IG�f�L��S��qv����C�LF��iG�c�6��ݚ.�x����Hɫ�"Z�bY�ۙ����5*���G+z�eΨ`�ۘnA�0�qQu��%�AWV]�܅�C&H��T'�[\���a+ZF���Y�e_l=�n�.P��쎸E������d�r��;;q��$�(�S��1��7��(�\���n+�N��BZ�x&��A���b䱛�5t̛4�u! ʾu��w'e^W�r�by����^t��䬲��lkl�+N3��/N��zW�XV��&�*����l��:��6��Q�y�Q�^ۣ0�y��m�Yה�Ľ�7���Ftv����y{�M����m/
;m�V��m��Np�޽�{��h����(�m�Y9�x�l�m��;.M�m�%���=���Mj�2�+1�K˼��o;�m'y�RvY��z�g6�/{e�jI�Y��m��dݢ����+&�
H�m�AMmif�k.���f����Y�4�`y�m��Ai�Z���ޛX�M�m`��,�m�����mm��Yol��d����%��5Ė�l�,F�=�۴�^=����AkZ�Z�����n6Y:�o;�"?�ww]�^���Q$�Gt��XA$���6I�%�}��AeDd��;k��ض�n�����'�wJ�l�I��M�Q'�MtX9�{���?'`s�sxI�x ��f��fStW��! �Q%Ҋ秳M#�������$�{}6ITI$��E��ޭ�;�������X� 4DY�u�9����5�����q�t���¶�aj�Y_<��G��h���0���@߹��7���� ��02�yJ}��5=�d�I�qb��q��ژdč^�y�ߴ�Z�z��Oğ��6@'ą���@�o7�~���{�53�j�AR*������ k޵���@��,�Cg�^�B�����D�wM���wU���#"��q�IJ`ߺo��Y���n��Q$����T&�4I�ܐ�@'�kg3vy�ig�!��ǝ�q�f��Kq$�BB�c�w�����u���JF���8�I��i�.kvmXxS�+2wYɥ[t+�xx{�����wDDo�co���A�?n�� 7���]�����3'�@��t�J$��,�A�M	��R��g��;�շt�wD�ݑ�t=u��c�m�;j{y�66�+Y�5��aϺ����AR���$Ѫ�[��ѰLDZuF��$��5�uD�t�J�$P�k�'��^��_ ?>��,�~3tmm��M���c�����M^�_~$xM��	"���Cr�we{�����Ŋ�m��V�#=�^���O�tm I=:��ޏ���v�k��J�vׯ�� y��Z53�j�X�$Q�99���{_C�/b��&b9�P  ���I�w���+�6�ʢI�֫����=�!j��.��֝h����=��������5o���|.�������|�����MB�Q��DnRUFW#��� ���}=��Y�M��RȾٶ�&�ҵ�u���y�b�o�iuz(VL�=y�ςHI7:�)utx�Xo1�i�]M�W.qk�s�ˎq�n���6���[�:v7e�&l��+�}��76{q]�������+��n�/�ێʭ]z1k��yF�;`�=\��c��Lޓ�M�m�< ZQ�9����s7r�s�#u���Wn��tv���=s:ܣu���r>��xƎR�X�!���ϭ�{����rW!�/Dv�]�2]�9�q۝���)�+��,
9llvN�#�{M�B)�l��~�~��9�M�S>~������ Y�o3�I?{�6@3�=m�Z�>���i`TK�{�֞!{�c'kQH:�Y������|�w����j��r׀|�� �F�&�����$��W�}��͉:��C��]�m�|}#�q62�f Y����Q'�}��B ������z�hԝdOw��	>�t2ƒ|rV�&"w5_!Z9�kY��mN�`�n�� �&�� �4^�`�V)gyv�m����X��K~"�)�{�$��&�}����!t����_�u�(�3W4'��[��O��TNy��޳��
D3u�H�L$���b���ݶ��YKkzL�]u�L�P]u�o�_���ߐ�uu�oQ:7���'�f�됟�?i���FR��W�QANo�A'���$��X6ܩ��>g�|�'uu���Ǟ���2�u�������`]�a<��T.�n.����js�I�޻�'3�엠+qy{8n���[o�0�����J�`����1}t�7�g|��[�gh!w�MOZ"8�v�v{]�-�@ ��נ> =]��z�o�a�ܓ�u�����{$�O�y�Z��τ{n&§~5�5�v'��Y�'�]�>�d�ĵ� �$�R>
"W��ux9h>�RI(��9�+���J�2a;�W�� �GΞ^�yަ�ÙD�KzHH��>̧ٜf9۩1�yE�D���᰻Ɲ��P�g7�a�t���ѻv��'���P�{�u�g��*⚞;�{{�� �$�~$�^�l�����P�*8�vg s��z�sr\nB�0�q�V��==f�zy��M}�
���&�����A%��N���y�@%{�k6�A��a��U����;�Lڛ��滾g��݆�;�ފ�m:ۖ��NLX��ą �5��d���U�a�~�}2Q������ݍ�T�|;wR�9�B�^]���c�<���z" ���z ��9�Ĩ�x��u�յf|]{;��w~��|� s�k�����v'��[�s�ZPܔ�ɟ �{گH�o�kj&�/�1aۙQ��Mf�lf@��{�p�J/���jNHD�M�����ܽ�$�o7ƱyY��h3��jD*�գ�d�v72�<k�8�Ơ�[��a�G�7�u�-�՟���~�RM�v�E�Xğ�����?�ݭ�$i�t�)��H$�������Ga��mR��3���w��n魬{�-�o8���_~ �}�ǈ��n�A=}�<��Q%�L���1��0��;q`|���c�@$L�n��W�;����D������ �}�o{��mf�66<�������k5-��I���ɢMQ'���	$�.�[��'^ޞ�.�g�����&;Y�=�t��{m���7z����ɓhwu-v�;Um�����q�4�ڵf�8B"��������ހFwܹ�����%�jڱ�w߉5D����k���]����D����$���I}�Q'λs��ϳK>ь�x���	+؀��	~�ӛ�X�q������<��S�:�~���}��H�����7鎙5D�����>��&��^|� }���je���r#���'G/A�Ga+tɈ��W����S��ˡ9̾��dlk��f� ���
�cE��6�)��1'�F�$��dM�>��%B~$������I'�.k��~���/.�Q$�Qo�ID�$y�`TO�U���4,^e��8t	�ΡB�}�|�绛�l��� ���b�3�v���ݒHI�������ly������� �8wy�˲�ǵ)=��TIޛ�!$�G�  ��z7�xW�;��4�X�Vl��X�����im�uk�D���E�6��Pn3�9K7�ٌ��}���b����[��^�_�	 ���ؘ�${[x�]ps����j��Ev8�-�6���n�O^�ɻ�v�tn�;����<{;Wk���nΓ��z�p��gA�8�B(�����^}}�N��{G����ɧ���gn-��y�:
4v�k�����j��(�l]\n�K�����m-��)�9��p��ݺ-q��W8��(g�òOH�Z�u��ZNͼz��MAڧ�r��;�
;n0���]�x�m�ӎ�8\s���[�W:�/?���5m\�Z���h���D�O��v蓺���]x����߽2��oτkj6�/�1|�t�$��8����w���6:�4I�숀O���ȂM��w�؋\�����Zs��J��&|g��������I�&��������wv��Dv���w���b}�=��e��3��q�+��p��D�{�Q$�O�譒I<��&MŚ�멄�7D���4o�je�jKPh���xh�"�kc]~��Of��T=;�M<ƈD��MkxA$�/v�*��\�.�o��o��23Dv#�U>�6��#�m�ua,;$ѝK��9��(��{| �cLQ���r��  ��,�k�����~��6W���<�}��4 �N�2�8���h7mY�ֽ�������W�oŋ�ڰ!+q�M;�!Kt��9��,={wGa�F��v�
�Q���S�lE�p�&��-T�����K�
ַ�R�Z�V�!�J�������gj>��N�& �~�?s{�@��I���4�95�����̍s��c��k�������!5D��ve＾L��wĚ$Aݫ �}�ω3�Y�;����0����;���߻�| c�,tH�v�	?j��&�P�l,�zU�#�y��@���|��u��Tˇ���{[�;�h0���I��=�eo ^�����=7M|
y��w�������ԏ;p�"扖ݩ+�!^���N8]��2���8�0�|�?Nr�V�A���{3G���c�=7G��^�j�Uݹ`��2�50�T}�sO�X �T`�q���h�y�y�8}���&�2{�$�@?�L(�h��ea�|R�)GI
�ul�$����
�(Ӷ�d׻�[ >�r�  ��dR�{��nӞ�w\�������W�,��ޛٽ�������R�8��.��TKV�Ѷ���僃8�/���<rޟ�L>_-�""��i �p��~*�ߦg�ݛު�t�߮P���{7�@|�����oW�x
�P��$���I(��I�u|����ML;��7�o|��%�o.�ĭdR��{��$�$�p�A��d��b���:{o�y���}����R�k����y�ٸ�nn�M���Ɛ��ƛvQ��o�߮?P�!��V����w���� �)����MI��_�I�qV��ʅJ��^��$ {���@t|ơ&W[!jw|��n�%W�݁}�oj�4H�숅�'�D��D�Js����w�}7ޟ��}z�J����_ @{���$�F��{X~��]<��8�Gg�^���߮7�����
�4�%=���U` e�� D����$�w��X6�Ԧl�m����T����{�T+*!Ѿ�U[Ζ���Uf�n�x����W2!t�����6��v(��VVA�B����*�����+K������O�)���Q�f ֽ��` ���7���p2�|��zxB���NxDC}�w@���|�S�P�DH��I��"U,@m��z�񎱯���y���#���:{C�)�
��t���wM lA���� ����{o��}�L��@�399��-U�kj�у2���͠�.2��;�@UD�w=}�x���b����;f�3�ă��N2]l���<����Yo~���I&wJq�}��r��BI%s��7��{���q�k '%(�<Č�����{�K�σ};�YD 繙�ٯY�_������os1P�������4�1��g��5D���TO��v{�o|L�r�H�wkl�I��疉��j��^�1
�®�Ʊ�(�+��Ĩ敤K��O���0`M��I�3+V�"Pj��F�ι�u=�Ծ8�)v퇯u�GXoj���6���4۫�����Ѻ<_V�U%n��-k��܉�x!ua�����n�c�-��*��@u�q�^-�f����u���+'1s3��em��&�*+��+	��;3MЗ|{�����*���8ZW����J���N<��37�ON�g��֊<�����n�ml���qp*�v%;�/M�xI]��9�N̼r��U��4q��QL�i�{�٩Ym�R�iH�l-bI@3�n�@��+S٧2M��Oh���Co'^��0f>�+�Q���'!�@�ԷX��� Ѡ���|��h��E�ea$���Y�$K�,d���#X���oi�Ġ�Lă�4�S@�T�{&�:��gh<h�FΞ�\
v>�nm��/�Vn�'U��x&�Վ��}t	�0Z��ɐu�gv=6#:�ե��X$Azt�Q촙�'�k�f�1�yK��`�SY{X��
u8k]Y{Y\��W^�xV���$����d�[f��AY��"�*���9`CRh��;u#p+X]lkuV�[�-�:����.��[[�}Ե�Ng.ezW<�Sݗ}X�`4�ή�c5�[����n�gWZ�2�A��0s����QP�X4��Ge��Zz��`�W1�aIEp`�ar���>�Kw���|±����4�d��+�
�4�@�w*gv4Y.��K�3jq�ײ]�Hb��UQ������Zm�����v�k.=���g;lS������9ȶ��^�^�[rE��RXyy��G2�-�Yl����z���KM�l�l�&�V��R����;Kmڙ�v�Q��{�dv�ͬ�����dY�����I����cg�oZ�Y���Oj�y6!��&e'��M�)mq��{׶ѦۛYnM��䙋c����n	�fBY�����=�g5��d�{��Fͯ{�ۈ�����qD��Ѷ��D�f3$Z�V�w����ns�{���Z9����w��,�Vٶ���ڷ�v͒	�������;q^y�t��{��/K���ュ���[hͭn��(L��Hrf��tS,�ǝ�e�tmۜ�㶱�$  �om���9>��R�{����Nn�V� 筯n6x�j-�n��i�������>sf�-��ځ�c�L�e\G�E�<p�t1tF�1�t`�Z�tWls�D��&2���흊y���g���+r�;���fM�
Iq�Ѷ�u�.bεv2.��u]l�F4��;s��yX§>N���w�'��J� :�9}��.�`����u�'$q�ϧ����u�5���Z(5��&�7^vD���p�:�v�I2��=s#��s��fɎ,i��84Y�\��^�,:��J����:����;G473�i��w]�6��s���F���n�F��`�������R�Z�\�Y�Gi=]����n���*vG�K�����7k-��j�P3볏GW�ö*�3�v{Y��ǫ�1q��4{vMGC��B-�88����xp��ri^(V1�!�s����q����8�����^��
�ʛ#Y�&��l�G=n}�Y�rh������m�T���Зe���N}sY�\)\�{:�ru��w%��;��r�J�:=���tř�vӻ]�㞵���v�a�7K��N��W����E��Sӹq����>�c1�.�u�/=^��v��獻q�::�u�m�k�ݸ���p���v9B��>6�6�^k�uc��v��1�>��s�a7�֝�'z��x�ϱc���u͛Ͱ�0�<�1p����G,;�V���Qd����8�M��+��{{�lE3���]������'=,ҁ��8��������s��{;����t��l�!��C�|�Q
P�;m�&����'vwd�v�	ʩ��q-V�����6�y�O/Gr�؛ٗ�]�ս������6`�&�O\+���s�l�C�۶t�NC�8��E���s=��q����K|)�K��g�.��c{m��W<{%۰�1Z������.M���)�5���;2,�q�uj�9ڄ�k��J�֡9E)SRJAY/�_}����!���S�D���Uu��n�*�b�ΰ�����Еn�cЮ��c\��8Xy�x��=q�u�^e�jv�Q�4�{�\`�S�r�-Q�p�vu=�y�-���13lU�ݕ����g�מ���,c�[|!qWd����x�t���l/0�����j����Κ-rk�v�m�]eA]���5��0�����d֧pkx-�`�G�p�G�B�=��݄�Wd���m,`��~�?E�_�?�]ަ~繬� �=��H:yJ�aǯw1-~�30��TSp��0�\Yh�N���:��P���4I?�������e� K��]�l��y����^�b�n�r���7����=�� ���[u�q�f���l���fg� ��պ��0&���,c��C�1�2�+�@:'�� 7�j� �	��f����x��<@}=��bc\��R�Q�(��� D����T��sdyt��d�s��ğ�?ܳ  "�ۍ���Y���=*(�H8�(��)����k=��vƖ���i�/-Ȟ���_���Xn��D��H���`k�����5�ܗ�����O�)D�M�y��G�"�������3�{���;���B��a�4JJV�<sU�<���pm<�Ӱ�di'*�VMO��;'�i�묇�uJ��4�=�=O4=ifZ�#\���K���﹚�� ���z �~�N����(Otu�!:�DE�&�;����L���պ@$oݹ�� �q�[��un�3} �[�g�${=˘�ZB�xVG@���3�����{zj�0Ď���$�$���&�?{��$O>k�m�����{���^���
ے�\x�f��t���i��|�_~d�IK� ğ���ctH$�{�n��]={�8�����~.;r*0̎��P�Vw:r��J���͹2�qI
r뾻����E3b@���뽷�y���������ă����.�T������A��� `���0��m��۶��%X�^k� 4�i��-��o @��o�ǀ ?w�����D���z�y]tb$�v���5S��3>�n���;�ŀI�}Y��O*��fE{$��1�0�c�Tw&+��ć�lf&��[(#�kU�[�t�,N
�${�oi'���j6�Y�n��L�;� <<S�?����鷀}��s3�c�,-tɁ���\߹���w�f�{ 9�v�� �����7�e����rݜ�m������,Ӈ����`�w.#��f,>{-o������E7؛L:$�i2Mh��RCt���Fs�Ym��R���(�5�L��$h���\��~���n�K�ݯ��ZYK���� 7��������=�{��3�ï0�{��	&{�l�R��,�V�Q���{���7������wC���6�I$�<�� zcsգk�Q>���O@���EU$MQ̉�y�X6 }�[� 7�4��PZ��w�� ��w�� �z�����"��b��'	�̮ۺ&�i�+e����B!�Zİ��5[z@#��.)9�w�����B(�Gv�`ʌ��x�� ˒�5V�&���n<ׂ�ۮ��V�&��t�,$�m����9id]�00��> {�ğ���	��u$��6�[Xdo�ջ�A������ݞ[���ù�$���� ��� �_%W����o���KQDEDT�n�fx�v��Jt���S�^9^�8�v:n��px:����J�Sk��H﹙�,��و��&��^��`�z���fG��b  �v�$�W��L�ZYK��/�؀:*�=^��Y�=�|��	&�gu^��{����n�\��gM�纃�Nq��*���m��|����0=��|7��T;�{��	{�m�1 �����[��quW+���	�V{���/w�C7�ĒC��D> ��� s����y�W5վ$�[��7��"r4�S��1�N�3�M��M����@]��l�$�5�|I�C�q?��I�����/�}����s.��ff{z�K=�3f]Ȗ0���� �E�z/Mg�ܵo�ݳi<�"�p���7��-��ֈU3�Kx�?/�����pG\��β2�	�kz���mrglSF�^6�2���A�Y�;����n����q��`ø�li'��mڽn��su	�Nz�c��pvz����.���q��[#xM��%ص���8��Wq�&凗��� ����vn���]�d��,�p��<�m����۞s��-���,�e�b����7`�V82؏^�l,�l�����v�l�v9;�.ǚ-���8]�	�&�R���r���ߟ��93͈�����n� 7�M�� �}��x��}�N���N����d��d�p��J�Sk�s��f}��Z��Y�S�.���4Hw�2� ���m�I%����ԍog�!'��F��v��R���vw@�=�f 3��=�&j����voX��<�UD�B�Juy���Q	�K�6��Dy�H��N�&�3��~%�f:�-D疂�k�� kޞ́�϶�����Z�{]��  y�[��j���mm�����j/�=�g2�$�I�ѶIoַ��h>�I�e��ڇل,������|��9-��Ս�]�%���:�������=�NT����no2  �=�f~.y`TJ���oNy��6��=���}�{y���U�~6"��& ��W興���R웋�`�;ݢ6�a��"D�
�6��I���M�Sk�΄�+�46��3]n�"�o�*��t݀M֭C���]m���" ��9�=�b�A���H��s:���3������no�Q� �w.�{3���ً�@4O�b��vL��9�I$��s3�.�n�_�'6:�$������ވ�h��[����""v^ N_j�$w�b͌o]2wN�>�wZ��[u>q�k�:�C����l�I>������[��H�~���Qg�f�1 {^��@��W�����wϟ|9�Ӭ�fս9�<�u%�o��osf��' 7#�#l��Z����~�nz�T`�|�G������Y�>�;�wX�'�����{ë�` �_�-|I�q4lρ��� ����2�e�^{ݫ�N$6�$����$�9{�:$����]��z�R�y�"�X_����0��cz@ ޽ۧ�;�;Vw�nL�{��ݧZ/����랉o�*fM�N��[;&�U(#��S��jE�֯�ـd�E��; ��ro�	���5�=�gz;�$�Zˮ{� �9;����ۘ֛��ȝ��;]ˈ��d]ק.�l=7��g����|��w���r�-8c�E|I�.[����mou�6�VIm.<A��n,�A�O�Fe�,���-�I���d ��cq�}ٙ�"�;�V,]&�	1 w�t��8�c���a��y�]�9��\jv��k��WmM��{c}�r�u<znv@߷َ�?I��$�H�{=[�;��~�j� ��}����#�kU:5k�=�s3���^��dx�j���zǀ =�{1�c��-�Þ�T��?���UR�����s ׽��σb�{wՖ2]�Q$�F{�0$�/y�@%WW�~�6�[Xd�C�!��61�u�7d�I�'��6@$��I�h��3�����A�U[����y%�����C�>����2�R��]�±\�����K{t��"���1�0weә�o!Z�B�� +?DG�w���-o�R��[ �U�{����@��u=���S���A=�]<@$��{1������t{��*k�S@S�D D#���b>�Z��ԩ<�>1�Ϭ�ZHo@ug�ߚ}P����4��Ob� x��f 	$ߤ��x��5�;�,z�ze�@tI��z�$ԩ��kWꊇ��C~�TkM�����nro=�ky�@rw}�� >5�iQ���KP���{�g���H{��1+ֽu#�~ɋ �A�M}@�.�mɮ}���v�$�qN�$���]�[Ǐ��X���6E�<����{7�P5��`�/'�b� 4�����=7�/���\��y�������W�~�b-�20=��@���y�Mi7��������޷0� d7ٯ��������.��u�����_5�K��I�_a�S�i��5�ZJ��Ny[�0N�ĉBoDؚ-��Kl]f�����Y�z*�P|<<=�z�H2&[���dM�g�����׮���㔧v��m��}���{u[Z8������gv{i�V�X���S������p��0�co��W���NT]zl�����r�g�p7j�f�͂5]�%di.:�Ѣ���dθ���յ�ۢݧv�:80�b�n�̎��v���6�g���Og���횭c:i���z�/u�����]l4��˷vm���^;vɃ�.1�뫳y|���l�6��v5��������ȝ��u[��;��4�����TI��O\E��J�WY�޲~���>@#!�M*u?V�8Y@�;tK�_7f��u?N��� ���h��( �7�4�����d�˵��U����4�}�0�9/�ꊇ��C=k�&�?�ێ���ؘswVU֕gw�7� >2���`ߦ�����"=^�9�3����K2�;W� �s&� l�z� ��p��w���6O[נ�s&�,���6�UE��<�N�m�Ke�\���X�]�]��5G���Y ����Ą��d���٧E�DJ�W(���f+<"�^ɜmkp��<*GP�,qX|5 ������:���ñ��OQ���M�C�����5��.���l��J��{���Jַ�P����*-ɟߵ�M�����󑳬D�b���%^^
�5Cs"�24R�(p'KU7�;M՘�6�x���4aj̤*N�x"I�ƈ�0�aT�#Z�)!.�^@��?����eI~�I?��2�Mo��CtI&���`M�/��K:���?,����GeV`tK�_"�;��?�4L�:��u>R��8+�7/�$�6�Y�[�Z�ǌ|��~�TD<���\�V՗\�|s����\Xg��q� 0�+������M׭HR{���V��z�`5�V`n��^�?~$3;�}:���W�� ����� ߽������t���Ϋ߹�Mh�\��D.:9�;��[L�n���l�'+�[�n��j6������7:��u'=�s{˧� ��$���D�}�h���ճ�{{�5��@b�;����T^P9X �0ɉ5ث	'���!�����l�h�Sܠx��0�.��>�y�μZ������C_KIQ.LG��c�=�I��q��Lo�7�
�RR�)���IaN�a'�J�k���ʶ\:�ӸO&%����^�w�g�o��h_M���E�w�cJ��(�*j7wU��s����)
�Z��/q}����y5LM6�X�u���p��TE�5Q�9k��A�ݼ좻M�kޙ�V�h�m�]��B�c̎�9]z���ٙ��.ه*Ɯ�i����R�ʬ�����[��h̀�/�e1�m�$�F���ht��B�4�50�}yKn*�V�XC�Op�엖]u&
�����l�571�9��4�}����tU�9}:Di����yl�s�ޜ��j<7ca��x��Z.ߝ���&-�o�e��!K+z�c� �	n�qߖ�
��qd̥W��w�z�+$�P��(����ɹ-Z�5�.d�/_ef$bpR�.�����(	�����=~��h����Rݒ
%=�DF�ŭ�b%�ӱ����Oj�
��o9v�jU��졤>����75<��n�W.���0������V�L��ܡ\y�˙�ǝGC��3��1#+��¶�r>�V;>�/nM��,�!���zU�_����{'�˷�C���
�ܶ�db@8:�ح����pH�w8��칕��ϝ�ajY���6.:θ�+�&ܪ%���MMD\�A���=���3�;Ǧc(˻W���8%9#qʫb���2�h���Z�0���m��8Z ^Dqc׵-��Q��Ӟ�	�[�+���*��ʒ�R��U;1�c��!-��g)[e�t�X�-f�����y�5ұ�nlY֚D�(b)T�h(HO�SڰE�h������(�ڵD��m�������l6�;d�d�-yf��KlPY[n�#mI�X��Q�5���m֐[c��kt�:#��-m�;h-���:δ'�{���M��.ˇ)�Ԣ4��kteu�E'����/1���+nӜ۬�mX���U��N̝-�8�:--[gq�Y/m�Y�f��$YXk�8�LmAt�{�yGf��h3��pE�������{b�;���4�'�1�mN[nm�:9�m����+[�\��A3]�ge���ڋN���ó����\�i�Zp�3�[V���6�I�={޷9k���Y�m��Jw�c�PS� E��e0�$w:���U��ۥ�UUY�s(sI���-R�)T1��w�驙�G�<��x�Pfz�ŀ� ��l� ���w��Yt�Ch���#Ҩϳ�tB�&nX_I��dM?2�f΁�{[y� ��ݱ� �s.g�}�kW'�t�>� 8�1ʚ���[��3��ǂ�݋�!�ą��]�F}K(������vO%+U�c牝מ� >����P@ 5]<���ef힘���\�M=믨}8'N+D	��{7�0>'�d�����%���~dHGݖ��D���� v`/�p��S�)��1un+���C�t� o� ��=�Y��0��I��y�1 {~��@)S�(k�b$�Irb=�k\��ִ�� p箕��ؘtI$׻�C�	�
}�ͬ�apέ9�zJ��z�1��E��pa�m,X1���2T�X0���`ܛj�a�(i4���,�{sN�� ��6~�uC�p�ڶ�]��3��s� >w����hk���o��f�cz�ى�	'�塁a�]#���w$�_?N���˳٦���-��e�k�Gvй67��N�6�>�U�Ƥ*ͽ����~��|�ws�P���X  =�k�0"޷f}4X	Z�d =ޘ�Muiۻ��X-�~^ �10��ݱ��&�4I���}�Z��_0�}��=�(�[�~~7�d	������> =��=6��Zfh��>���lG���m��/w����b��P���F��Z��9�)�>��s��ϰ;��=` �=@�Z����sw0	���U؛%Ara�sX�` =o֪$�����e��>�mQ'ʹ� :��P�z""	��WY���4�U�ZTR�X���^˧2r�ũ�F:��:�$�=g�>�
��ګ��VH�v�����.�	��i��U��U/��W�j��S�ts�\�m��Pݏfñ���M�e��W�.����猕�l2a7K0�j���6���@X�Y��]�Ө]˶8ct^}�<lh+g���r�"v��A�����lA��٢��uۛJ���W8�z��;j0�D�^C��l�X���l
�ˎ�8�pt����f�aX��a���؅Bȝj��n|=q����LM�sAgv������m�Iٮ�CDt�y���^o��e�J�-n�K�.�<�ZA��&���s�;뷋 ����%�e��>�e�w�&w��&�z|�*��"!�#s~�_ ���׋w����k9�I�MN��~$a��m�6��/B���i�n�|./;i��WE�{z���n��� �fmM�K����9���@{��<ϐ o�hm����lVQ�&7�c�w��9�/�7t�H/7q������H�*��@�t0��]U��~�OP���߂XL'�S@��v�]꺹���-�@k��<� ;��i =����5IO,�}�[w����Ϫ��[e��e:&�A6��^�<�'�ȅ]�Q�*m&���>�ê����;�k` n�N�P> =���S��h��ͭg�ט ug�t�>��'i	1�g�ۋ�%��~��I������׽Qq]g��+S�Ha�Q���YfE�9;w�Qwn;�$1*�H|Wm�q�&g9���[?x{�[N��d���%I'���YM�A���[���m���q����Uw��'�(	 ���.` ]�K]}<N�� ;�8j���.bˇ;%�R�QC�|n������L��:k�  ��k$ ����ˋ�*2�&�(�Wr�
���A��b�O�١�ϩ�=L��N+�%�3���`D>�F�D[�Ҟ.KՊg����Z`���?����_X���y{���{��vT-��cdΊXФvW5����;�K ���fJ 7�r���{\y������ڋ�ά�*�4I��t��T��YH4J���{~�<�H9��o�{c��{�6�$���c��������~�g'�}.�wkEe�$ǁ��n` ����� ���gr�GlY�c�!�#Ysu��	`5wflt����,�t�.t�������T��p�-t��ܻ���u�i���~K�}���~�s>@ϐ�{[y� �>L���~P����^\�����ϵh	���o �{��� .響꼟t�뷠�v� ��{���S�(f|Oo]y� 7{9M ����A4����"�e~��L2I'���I��rg��p\����4��h$#�Q�+��k�K�n�����|���݋c(��r�������gh�R�����{{˘�{��zm�Y�j=$Ys����~��]�%���g����o��~��w�������u�$|z���g=���ݺ|H �}v�� oz��|����'9u��}��+"�J�p�=�cİ> ��[D�����!޿?��� uk���������
�V��|����랼�~@ ���� l;�,�@��G�ӮR����i^��v�>��N�xp�7���a�La�{˫�f�gۿ��M�(�͌T[�짹T[������5+�2_˖�ַ��_.���{�~y�-��J_�r�o�\�b�OĒN�@���*[�-{ހ.s���@|�ֶ��>����F��a�֑����r�HR!B���P��3���/<�,�@���@�p�[+C�����lqI��מ`|���Zށ���5�BF���e�6�;��N�UX?q��VT&���e��;���;��v<>���  ���*$�#���� �4����π����D��vU��J��`MIP �w�K@ L��>Lz��#w��$��ي������T<�C.Ń����*y=|u,Vk�� �;��H��=�n�� {�P1^�y9{{�H�1Ujd9sB�U�$ǁ���,��뷋�+��{���l߬z ���d����e$�WY�i�m�@_������ܙvĪ��ga�3�RSp����FZ&i�K�:�\���7��R���zR&�������d���kv�z�� �w��/�ӹ�kh
�uE,jEaI��w�wl�󶸴]>)Ƽ�J碙�r9{<��e�P���ݜa�۷Wb 4�<�W��4�)�����@�έΤ�m�dmV�l��ۇw]c�yG�R��w͆Eu�!�u�H�N�n�kkC������ۄC�s�����6��x9�@�&q�4˹�7^�-�F��:LW�뵥�nsu]��^�籉�J�Gpk�{{)���=��畍�x�N�2�7Y�t�ES�:�Z���z���~��R�"�����l� ��7�6.����H-�����&�ᗧa��H�;���}9�#��*�1��^}��s��瓯o-�2e�(���� ���.� s�N<����l�z�/�F>u�2��	�ٙ�D��o�� �k�oj*-��c�$�h���{6�� ��W�����J�Y0��fV�Ý]����o:kز�߽����~����mz�5� ߏ{3��CQ��2Tˆ�k}�
o�7g����`kb�O�[�`2L�($�h���itӣ�ﻭU���{Q@hl���U:q�qz�W�r�u�c�U��݌%�?~���4*ZBM?�{ٔ��]���Me�+�ac7��5Q���a v���me:d
���c�H�߬�M���wy�kޗ��ᏽ�擓˻�2����qw,���/�y���m�gD��F���sN�QN�o/np�W}�>��}�5�?{��t@Y��6�V�����h���g�#��ߔ��`��Lf�z�����?���Iy�6� �r���$)~���ߑ7+bS�&7�]]\~��;�ї�� �p��� O��{��閆\������il�Qz(�߂V���v�5 ����Xm`}�c�������&��������g.`a�R�����Q�(��L�)��+��k��j�3���ۃ�Pi����ˉ�>���w�E�e��G�v놞 h���� �k��0�$��O���]���Z[�Ijrri@��U~��;I�{|�S'�{�n�a�s��tI����Fހ=���@�sk�{����8��Y�������f�� �=���D��-t�+���wm��8����O5gv.I��J0I��KŏK6��~h*K)8���5���9�v]�����ݩ��7a�}�=s����A���߁�����}f��q��)1����xpR�P˫4  ���c������V���UO��ȍD���Hq�e��\���j�� ������/9��hw��2�Vj�'����b@/w5瘁t\��<���<����P\Q�"��Q��� }"p���r��x��Pp�NDj�[]��e�%n.�"z�4�@|�wt� {���^�k�އ�yFޒ�7s>+~ɨ��#%b������$�^��OH1��լ>$���9�c� {��<� .��s�a��zO���v��Z��Z;I���2�w�x �4My�=�;��j�@H�w��� m��|����M,�����~�*���f���P��$��^D�2߲��g��Xn��6��B���̄��ї���B�����c��Wn#u�f�@����k-U�|N ��P���7���ݞ}������[罍h��^z��c�����_ϋ o�7f�sy�U_I}��	��� -�5��@�ݍ���.��8v8%\(�H?�Q�JW�n�P�s���\��ʊ�J�J�j���Y�~�C����<�g3.,���,���編Ie�s�p�Ćz�!ju��Lwc��8ߪ���%n,���՚ *ݻ�;y�]^` ��Y� �����N��~�]��y}k7$���vh�9+r�oy� z�bmbr���G��� x���t� -{-U��I�?�u�I���k��.}� o9�����rkڏ_ �w�9<�HD,�@mQ'�SΛ&Viʄ�%��X����s�l�yq,=���}��.�w�Ř�@|{W�m�{����^Y�7�� �RV���-�\���(��x�	K4*��4T4Ve�уÛ�GN��[� ��W�,���޷���>���n6���`��B�}[�l�WF���<���wfٚU���c5�;,�fXC�Pz�Ե
ئ���73���%aQ��+/��&uI��,�ʆ9{t�e�x�S���)M��M]Fhui��W��;�:��.��yw6�kM���;R�����K��R�
�3zl9��)���|f8�w"#����hu,�{r�ITp婖�%d�PU������g�>�ܾ�C�YY���^���k1	���CD;AUF\�T�^�-n�y��,�r��Y���HML|%*(N��輘�Jn";y8�9��YѲ��%O]��D�n)Ui�����9Ѕx�s�M��fw!�qmX��坆�s��֮�i��&6fU�mբ��ݥ*���n�r���t�]�˻�ڕ����mIx��WS��w���-f4n�#K���ݑ*1J8%��c�S�������5�Je�}�r$�)��`�v�uuj�p�����E)}���(�>�TwU�!)p4�U�� ��L=У�,�-X�bʮm��s��~,5��y��z�t���h\����wH٥��6��w{f�>�4S��9��m�g�ܓ =�j�A�2ݸ[�f㛮�N������ur�����hl��K��+4���;`.����i�膃c�9G5���ˬ�^�4ͻ�mW$���tvM�����T��Pen��R`*Q歽&�'7^* �|,�'{i�	'k[3���ӞwiGgi�^Sf�Y���^^�c`�������%�d��e=�;��v��<��2//;���:�����@\�z��������/tv�M�gyy^e!Ѷ��;H��Y^W���6���u������n�<�H�c{X�G��擄w���{������Ǚ<�޼o5��{��YE�ۇ�k���������f�â:\�:�B��t�ZZ$��a�I$f��N���e��Iݕ�$���ͬ�fn��NI-3kmZN(n�J
:B��e�w��';�,m֥�hr������{�K��N;,ζ�-�͙IE)m���m�	Ŷ6�E�2	2Ј"����3��jgj-m:�:miЬ���{ZH�;nȤ�ܛ	�m(�[`!�J�#b�����N��W[�X[�����wj:�]t�Gk��d;ٰҲ�ͷ\ڷi�X๝�ܛ�u�v�&�y�y���aA�6����� �/C�&y�v�'�Ji9�y�-`kۇ�p���\I������c��*c�l1ԁ8�c[c^�6�w$��s[H�ݚ�9�pV�'fېG���:B����Y�u��7D�}��WY�l �Ou��[�Z���؝&���]5���p	�ϟ�t�_��!�/Bmȳ�^wU�X�#������9X�]u����>�tuMa}���qW%g��%��g��v�>����9`-��n:K�u���rv}�Ÿ��Wr��Q��|��ǯ�ݻ/���>	�9O'�,�����y%(j���O�ݷ��O!�I�u�.�g��.����m�9NG��i�v���BVz��{a|�3�uը�Z�m��u���5�=�fGsݎ��>>3��G�חْ��3�z�y�ݷ�6��������V5^c���4ۮ�n :5�O8�^^zm���vv,�i����5Z��f�3Vp��[�p��ӜȘ�gh˟w��ӎ��A�,�k[�������ƞ�����C�.ݺ��<�ݷX�]x�_^�n{8{dݰ-n딎G�Q�y:�p�[Y<
6�]��L�p��y��p]��s�������[���oW��k}���:�J�6�k�f�{kq�63ל^�؄�6�nޫm���gU�0�:ڞt�.�5�����H=0`&.5�(�ocD���9����֏˹�&�϶1������_�2����m<�0��rv�8xö5pc�-j�ޝ����"��^ܸ�@���zV�n<{.9b���NI��q��v�:pc��v�8��rԾ:�� �n���b�ٝ�8���Nz�n���y݌N�3��˔���uǵ/AW;ƣ��ø3��"m�n����/cF��lQt4w���z:�9���\a�y��{�6�p�r�=�7Wb��[m��j9�8�:v���q�xFݞ��h�ɋ-��\i����`��MB{[�q�m�U��X��O�&V۬k�U�Yo*�A�����<�N{6�{��vjY級�� -�j�&�{���oik1�}ͽ�o�ն� ����i5�֬�\1}k���{��GN��A1΃1��[�j��ڃ���BFq��cq�v�':x�3��n�����]n�]R��r8����*^/���������D���>� =��k� �{��<�8vz,����.ob �e�4��Ƿ�8�~,�V���˘wZ^��}���m2h�I��D"OĚ=��`Nۧ�r�^������/�J��d�6�� �=˧��o~&��=劦�I_e�Ď�n'�&�g�$�؉Rᇽ�b��&p| �ˈ�H��S�5D�?*^m�u�gV�o�����p���UN�	4���N�g�O�N��5ܵ]��%�D��� ~��@tI�?:`���t~��m���W���f�m�]m]��u�����7�W�F�u�F�*���x+�r�լ|���  ��9�#m�{��Y�:{���x����ؒVuV���MJ̘�4�hWQWT���w������V�go��0�:�+�8��!DL���эόAm���w��{���|T�Z�ț��n�s	�MN��efOJ�x�n�� ����o`6��;����|�G��c�n|YF�S1��n�Q&���*l�~%,齊�{�8MW����Nf}������:��5�%�2bAۖ�l��jo2��Ozfd> ��o`�[��1b����n>�.�32��Yd��2:��J��I$k�b�s:��[�z��&��Yd�j{���$� OL�TLU�w��{���c�O$�!Ϭej@�Ϯ���uavlk��ON��^5��۔��M�����c�PHI����=�d �9�oK 6��B%y��F��*Sj�b��Y�>�F�>@mk���P��X�g�n����+�+ �]��u_��P7D�o۷H�}�ys�s���]�=y�P;��]�*�j�3>D�k�>�@홋�$�&���y�`��{s�>�j-�Ĥ��F�YAPg��lV��x��V�͸�Y;4zU������t.P�mw$�d��R~���I�{߳oX 7�v��>6�����Ŕj�1�/ż��nOri�D�3�d�LD>ۣq��J窩p3�ΚFb!���π�<�j4����̘�[� �=���\�/34��_�hL�I������Mx!]����~W7� w����b瞀d�K����n� t�:Ov���:��/y��EP*�C�wtl�� ���DG�	�ҖNDpBW�77�u� > ;�[�5ך�Z����â}sxh��{���V�1�L� �^S@���F�fK�n?���q�V�W�!
�k� �N�} �g��Vρ8���k���y����҃ H��s1PB�s��l]ef
ʻl�����b�G��l��z@��M�& ��=�y
md�ǧ�a&|ӷ��η��@�Ӭd�o���R����Po�qU�V�ln�LN
0f��S�IM����L��,w����<�	�����|�W>,�����gu7� w�,5������,R�ր�SW���$�����|���tL٤慽dWb�]X(
9t���Ϣ㢞v\;��Лt1�9c�u��"ݧ�C�O�@�ܿ2;��&��$���t�I��0���5�J���(����� >G���bמjY"vGU�?wwO�` �Un��y�2vv�$��"�$�|�`:$f���J�����&��<���B�lrLx�OfA �<��-�5��;��rȉ�{�����o{ݸ���ൔB�jZ!���׷ԸR>�8��7$>:�Iy��٢@��0�I&_�� ������w��̀���U����j�3	�� Ne�z̼�w|]����NmfA:�`�I��/3)$멉dt�f��yt�)h�<�x�:�����8]#+m&�Q"��bq3V�W_;�o
Ω�����3;+���˔0�5[���v{���C�[O#�v��g]�糫�s���g���n�;y
��o.ō
$��n95\u�v�Z�^ǁ�m�y]]VEm��M)l�|㯏a@n�۹]�A�;'��˭۴�a�eZ<��e�<��p�d�n��Լ��ې��
:�nzp]i:������*�!��=`���=
Tꃱ�t,���� ZX�8wE�꽝k��������DSWJ��RS�5HAAA�T�Pj�&���tT����2)KϳܜٰH'�w���Ȉ=s�}�ӟ;Ig�˺��!mx�R����e��Me!���oϦ��sc� ����$wo��i�{7�F_Ow7���cj�b`����Bd�sGI$W�`�I尺's�V{#��H'�uY�H#v���f�|j�*��3;;4�ݷ�����z���	��Y ݺ��/L��ʩ�|-@��@2k�B�{�`�A��wʻ�g�\V��}u�͂	n�z�#�5g�dI��y����Z�q7QX*@ZO}���/�������e�"j4�b��������t%p���,���\A�İ�J���T�בΰ߉�>:�z���\�T��Q5�Z����S �[�����Xa�+'���S�f��5���l,���3T�js;���]�w	4f�߁;#U}�;S��	[�ƶ��U�Wf�0 u��h�
al��AN�'��bY�+g+tb�{����D������1^��Rc�͝#�5�0'�d���V$��j{HM��g9�J��XA�䃪G�쮰�]�Þ��q��5�X0���og��TjV/k��Y�$����
�TDI����ڭ��H��
9��:���U�8�H'ݹ�0��,��V{�����gڜmdn
2H|��\猝��:7Q����	$���UF�,��kt�\؟|�b���	��]`I$�ט���]bδԬX�У���5���LMT@��YE?��UH�ѻ����ցS�s�O*�	1�w�`�k�戢s�����=� �yӡ`�P�J�D����;izu�a2��v�f�)�P'�����k��-�3��i��m��G����tA�̰��y�t�WL���y�'�����'�8�`)1^�Rg0y7�R�ճ���$䛦 ������<��A1��A{SN���X.��WvFU�^�* V�lD�ݮ1C^ZL!��fI	uY�	9�;b2�Hb��5,D�3���g-�k�cvlB�vp�j�X���TT\W��7t�@�4* �T�����o����	�Zl�
�!�>�IfSsf�:�5d�"f� P&�Δl1B�ˢ��v�X ���7�I ��-9��o���Jk=�c��߀��VQTk#:��O� ��n	��Fh"�_=-7�N�Qi����|V�~p�ߙkr�i�;��{5�.a�y9�O�$.U��/�Ջk�v�;�6A+�z�N
�*����C��7[)a&A�yW�(�/7Q{��V#����E�x��ǯ��˺�[��mˌ�H�6Hь����]��lg;J��퓛��b�u���b>'�&����.�#�ufR��rkd�:�.�q�$�"M��"H(,vx�
�}s�z������_�qZ� ��|��$љ�4&O(�s~$��p�$��Y�=�s2�TB���5��U�pύQ����!1�͊��GP�� �|�P$��8o����K0�n�zݣm@\�.,�ܭ����?g�46��o��`�	���|�b�Y,	�eY���9��o����U�������n�����R�$�s�,�C<�n/^���Z"s:�%�BH�$EQ5S������@װDϓv��Fu�{���H]�fy6t �s��6�.�߷`�Kk.4-.��K;�<�{b�eνA:���Sn
�5g��
ɬ��{sU�\陕�*��L���]�yy��\��&d殚mi����ֻ�t�@�9�s�鶍Sˮ�g����\
#�=mƹ���V������pF�:�k� �۶�xx؞%�* T���wgԎ8���N����[�v�\������4F����lս����P)[�;����>e�\�3�e�3�.�'����]>����U��n�=n݌��9�6�u 榰8v��&s�\����5ƞKvL�m�M��c�JtH�`AF���:6/(T8��uN����O-j�A.9���]��!dW�k]Ճ���`1����H�3Bd�RF:L@�ຮ�n�A-k0H�ri6���A^���i�ov�iz�c7���cll������|���L����>$okY��z9��h_��3D��|�h�؜���lռ�I
ɲ|	��졶Y�70��ui�����M���[��
�*�σ�� ��ʰf�vO[�qk��)}^&sdl
��;U�$���� *T�k5�\��>��X�CjS��!EA͕��=�s��r��^D��Q�b���Y��/(խ����W9����9vU�A>��`�}��ՓS�9z��'��eX���1B��3b]�o��s}�4+��㚂��1^*�qMDϊ�b����*{���?*t�=��1`;1{�nZ����Y��Q%]�>1.�ywwD]eE=�XA$6�	����箸�V=i��ں26�RPzO��_��9�m�}\�+�L��y��'��
O<Cq�0s2����Y�~��dw�S޹�6�Mr�I:�X�	�n���g"j��w*����ȓT�M��Ug�۫=�(V���C�1ˤY ��U���u`�����L5�c�ϱ�R@b���:�\e;8&�x{n���i=22�D��m�rʂ�~}�eT���!tCޛ$��eX'Ă{�Va�q�0JAF��&�>�ݛ���_��\j��UV�i�׻ŏ�/��є��qԚ�� �	�߯ć٫0�ʹ�[sUD��gVy�1b��:[&c��[�A��g�xވ2T��:��\ݘ�W�3�.���8��ɼ44r͈9̜��0�'��Ң�{^�6b.Ɗۨ���$kj���0�a#^[��V��Ս�	��9W//E�a�Ѯ�[���N�B��B;YMɗT��w����ׄ#}vA�K-M���v�z;6!�b;�e��t��VR�.�f��]wJ���C$�a�}	p�p��!�!����C7�,gb]u
&�0�����eŻF�ol��[�7��RE�fI�������h��9�Ү(���^s۾uȣݻ�Wٲ��:���--CIwt�>��\�pW�[�ǤI6�c���fiW8��v�'ƗRkZ��dn�Vζ�TA�YV�o]�V�*�	���N��9�*sC�͘[-^��jC|ݕ��Z=]�nJʼL����oM��L�*&�74<�ݵ��b��ږ�_0\�w��nI�;�v����N�LqZ4z(���3Utģ�f��U��6�w��W��M3d�0���{��3�P
�;j�V�9�h����0ݓ���PSP�N�IZ{�t	ƨб2�R�VF�ͻ� ��p���6��r�z��K�ؓop%60�#"�R��7���b%�-n��V*>�U��;gw[��S^�ӥ��k:�z)#����ͣ�$O���-rRNb�rŭ�rn\���+�N�|�n����aL�ӀV�IV]񽮬;m�@�f����͝�z�;�h�Z�z�nu;��ۆ��W�3ګ1�N���u�ql�6�gmT���MJ�c�ʘ̳6�%Zښ'E��@;��3ƴ����X�����:�w=�w*"[*,P�*"�d*��6d��6�HW�"�4����)(v�tq;Lviqm�������9�M�rk5�Yw�jxZ3"9#M��q�;-�[n��β#�Ұ8#��wg�ܳ8,��v{�;ð����hJ[YӜ���M�'q/l����
H�e�p�qݝ֕�Vp[[���*<��坐\�B��:Va�f\R���t�������۝�^M���mg$����6����È���-���:�$Vv���Ygm��8����Ru�Y�ge�l�Ό�"��9"�����՝IYiEwkrṆN�+���tV�V�]e�Xtu8fgcn�{^\�Dru�fwY�nݵd�Z۬�3�����DT��T���{vG�vt�⵶t~�W<H'�7���O�f��X��2I&b���FS��W՗\�$�'B�ٹ���|H��s�cN,�`�mvU��Y�3ڏ��o5��i7��������,�N�v>o�� �y�::����ήh�e5x��\7�!��P��݆�Z޸]�tQu�.�M��V�2D�;B�$h�\��o˾�j�	
ۮ� ��Ճ�z:����{����G5�>�h�@�a�Yy�fx�%VC���!$`��^~%�ט>$��X1,�uC�
������+����`�
�DP�Tfl۷��đʝeV2��^k����"�}��Z�~��\^��ťTt�Mq��̽�8�8�9WۘA$r��$o]g�=1e�Fr��e�y6�<�fV�e���W�뵽^O�px��W��z6��/~sͭ��uڞZc�k�u�����ܼ5e���0��@���n�f��]]�H�&jLA�^S��H)u����]�r���g����q`�u�n`$����m'���ۚ�f�뚏W�ƙ[���ù]v��k�Uj$r޸���Qc�q��r��t��K�\MU���&���x=��;���H��~9"V��U�S������-{I��0��d�B�T�&�JuT�2{�X	>)ӫ�o]_� �m,.D-G����߯vy2�(����㛼i�w��m����±����A��������V_ξs��J�UkrM|����g3x���B�>(�9Ak�X �ݛ�&kOk���y�'�贸�� v��̶�v<��y�:��P̩Pr��Zb��
 v�eR���b���܃��
�;h:M2��p�Ǌ�۠�!���S*�Qι�ަZ�v��v&�%;\6�`��Rb��e�k��M��6��5�d���$�Lm§ES�Z7C=��wNWB��qrc�v���%;;�����Ů3StmI��z�Z�kO-�]��o4[9��CK=nu�mdx6�*��6��ZV�qc!�{XM��:�XT��	����I�s��n��[���k
	a�8C��;&r��J<��D��a�j���i�ּ���kD��k�F뛳�[a����֖𺦐!������f�^-z�Y1�ٹ��R�krm����@����,;����!$W�jA�s��>��ՒH'�7���\����|U� =3�|=�Kj>���Wܾ�ћ��.]f��y���U!C��t��{�m޼��APs+��b7�U9���EW��|֕�:�'��IN�X �;�{3��6̢��k���۪�Ok�ذ��<�n�>$�y�0�H��~&�B		�P�EsB�=4�R�X�=�� ���`��h�L�D����Ho5�!zw��֮<������u�*��]~9�<w)y�n�6�[:ڣ��
�n8�VXk|8)�A��
���Ӭ���o`�A._X��$�H���:���H����v��UG,`����i���ku���Z��v�r���/��H��:��̥B5mjB��oy�F��
�{�RFN�%B�����h��I3�P oI������h�fvՌ4�9뉴k|h�-�O�U3 7Ԟ{$�}B�><;�t��R#)�Iw^�������50�b�$� �ި{Ƿ�j��A�K��
�sʐ�~ˆ��N�T��(��L9�	�UP^Fr�~$
x�ͩ|&�kEn�@ˤ� ��VlIݿ]&ɴI5���9ϛ���*�X_�M�������l8:�;���=.��+�.�oF�:8+��}�y���,�-��u�E����Ȩ�k>�ȷ�\�}���{�0�ٲ^�t	��bf�B��������m�ħʷ�O}�O7VlH9����Vvܔb�m�s;�t�ݬ�j��Po��i��K���MS���óH� ��y�"U�nm���)��Ш1f�d[ɪ"̝�3Sb�ʚ#P9�bZ���Q��v�Ӯ`�VQv����P_�J��wf��ͼ߲�9�腖�)�-A�����3����L��/oă�R͒H%��I!�j��q��%vr�l�a�  ��t�>�k�ϊ�>���$ZU��n��/��f��z�OJ�F���=8�
����w�����)6�n�>����r�.6yD�Z,�%cUo{�<�W�GmGmq�O�\��_f��v�����/����Msޙ������>�5�q��{�AQO��d�T<{�:x�
Jp١�s[��x���{��vz��A�B4Y�A�ϲ�e�;H� O9�� ���#�;[���bA  p�4���kt ���D��	3B`��4m};��{�P|O�Lw\�I�{�0K�VSS����/}�î;\�Y��-{�˫�Af���o���2#ݘB��v�������X]�����T��kn�%��c������J{��Ni����f��^eYl/R���|_9�����[5 �n,�Ov�fs�6�d�4�dV�0}�ȅ[��C�Z�(���=�����֙��i1�[)�kb���2	�I"�"	$a�}D�ۺ�<Gt�� �mAW���r� �[�,��w�6�����cj��D��zs��oBw���.�#PL��I)n��l�M����u���M��T�B�Ǥ��#`
ܾ 4{�]Z�լ�B�׃<OuS6	k`�&k�"�s����u6�e�	7ϳ0�w�Y�ӽ|�^�-n,��z����f������4&	��\l�Q]r��D�x/f�t���2|���$�9Uq�F�y[�]�ֶ�M�j�E�z-d|��$�o��O��^�WvmeԠ��9��ۻ��bي-R���9���u.��܄�r��&�&���uZ�j���oP��������ŧ^�����N����(���k���n�]�'`;�F�E⃶Ŭ�=37�[=���]�8�Y�ݤ�#����k�9�Ł��ӝ���oq��a��W��m���O0�@�wi� �oi��j�	�v}/V���w2�:$q[=p�8��ؗ���䮱���q�υ�6[�Z�]i��;��ȶ7�����f��+vzz�m�O��֢ϫuWWq��]��O���^O^�0�|_T�,�FF�͞���"f��wz�U����ʜ�8(�����G9M��)�ݽ��a� �M��Hýv(o]%PC���5I�H�G-3Np�m7�|}�Zm�zix7�%�@}�Z��U`�6E�$@�2G]ۜO����qH:�,�H$l7sd���KD�<��{L��mx$X2J�Lǧ�֕6���VP?#�o�V�j�;�(Pv��SM���f/��Y�v��"!����c<lI���:�b�Wp�[���s��nN'�����?y�

�B�ގS�|���ү��}�qf	��m�<�<rq�`u8�x�S�ZI��~�w1b��ssO���)%�ZY4�k��U�l�L���|��M���L��e6v�Esζ��xj���w�ٛ����/���	��E��<p�!�604ġ����I �ݓ�Զ�>Y�i���6��_F7�Mꈓ"7�j�GĜ�K=���fz�YV�F�Q�9�/��(X=֕�>�zX�ꢕ����|5��X���^�3Z���mf/��-�⊒����Ne� ���T
 ȑRd�wn�Qn,�E���ޙ���^�OmA=�n,���P�m�=��M�I�R��j�쭏��a�_Oc˺_Q��v8�AmY����d�:;N��ڮ�#���I��n/Ƈ����`�t�Y35�����9����cDL"����5��BK���mm䔅 N]�/��	�5Xk{z�Ő�4������2��y������� > T�t)'j�I���RT%8�s�Y�;�-��4		g;�wZ@Q���v;F����"�!��;.�����^�n����̴�w+�I�<H'��L�haȌ$Q��	�j�*l9u%r�Gk�>$���7�I ��`�J�cg�ܝ��=�wX�;�TtV�Q����h���UI9|�UЅu�fx�9<�g���ҳ��	ť�k�~^EMG�4ڧ�(��[Mn��97(���qj8�t�֕ʫ�.s�S�F��2$T�<m�;��˲�,dr�`����F���T�z�6!� �/uA�J�1\��"�ݿ1B����;�b�1�1^
��v�0b�yX��d
��;+�o����i��U�Af���Y�O���~$�M%��Ņt�FԴ�1'��&���;'7����NH$�8k$_���Y����k�v��A�Id �Π����$Dn��={���'�d=>-0��Kr�Sj��oC:�A�E{s�q�2]\��L:m�ժM>�&@��} �
�7F�UC��mA��uM�2����#WV�=�t	!�j�~�/uݗ{���wr(����K	\�(v����ۤ8]�>�V�/��>h#a~%*�ߗ��Nf*&*B��k��|H(��|O�٫0<l�o���6	$�Ֆ�8�hБD���f�簛�Ia��L�������@|�̪ w��� �L���~��S�|M�I��0Y���]� �yf�t�vJ�ɬHot[!����٥M�پbŚt��TU�Pzά��nA�{MQ �Fu�$�7�� Wz��tg���@P�_~�i���&�*s
�}�|I�qe_e6�Jy5&&�~$v��H%������F��h��~����u���g.��3V��*�����ŗ�a�VM�R�U���bI�i���'l5;8��ФΪ�3��9{��5�J�i��{����)[�B����mMh�,�����d-2�ZUsלv�$B���8�Et�j۫�C
�@�]cgjh(�=فg��0̹�]��6�I{��^b��Pll�X/b%3{�B�ɳ{&%tw�H�J�u٫Vw6�4.��w'�{��=/�Bg���f������-HBR*6�n���g���9�x�D��khF��D�Vh1��ˢdUe���K$%�kg, �Z.YՓFP���h�����O�Y��j5�)۹�*���*1�nD�Qj-h�M�4��	�'����C+y�!��ʈ�f��n�o��A�Iˣ�S�U�띙N�E�0<�-I��T�LVF��w�_[��kwf��s�Ƀ6�Q����V��M�u���*y1�o(G)�K�P�.�A)U���n;�&�M�@/~�5��Ԛ�Y�;)e�ԙ��Jˇ$@7��d�ִ�N�e�]k=�j����j��w/;��sx�hF�_AMr�N��͍kw�J�f��aK�q�D�T�G:j�,��\F��\vR3�uS�!cI�g�D;�d����c����N�{/Ký,�仑�~�ә+m<;N�!�ס�9meʆ��%u�����Z�V�e���MδS9Ϻ�@Tp��\Cw���V-`�w���0T5�� jf�jQ�WY��Q�o�/[y��֍ju'X�Y��g��{���S�;N�.�6m�Vu��+[q[n�;(���v�'��"N�,�fu���\�rtw�����]�Y�l��8�C���(��2����,���Â�//r��2�S7��6�݇��� ����v��Y��'�ڊ͖����"������j ;{w�E׶��^��I�w���3���9;,���⽬�v��[n�˵�՗ۻH����;��:;���eݦi�NQqm�B$����tqr'E͢�����<�+�lgdQն�j˶՜Q������mY�wyh�]��;���va�f�\2���˒����߬xܘ�v��!�Ë��L�4��vmknݸ��औ��K�[�oGmͫ=��4<&۹���v��]6g�G�.�}>�����ݓ[��8!�b(�Qf��ކZ3g��N͹�\�v��n6�,x��Su��hƗ'Sզ�<8p���cZ�2��2��Q��Ƨۂ�P{�Vtr��Y�<�;���Z�D�ưc�����'&z�d�FVnx8W@K0���2r������d˞w���ʱ��.h��<��� ;F�qq��FmB��������G\p-]�轋�zOe��ggѻ�;���rn�7C���|lVx�[]ӳ��ӫ�V�3��Z�;b׼�����}����}�mm�n�wn�2�y�2;m�d���i�.v�����ɓZ�s�[ki�O*D����c��o\��ۺ��I��8��7�rs�wa�]��#�D�>=���=��v��K��ŎÝZ.���m��X��cv����ZE�l�ŧs�*�'OSܖ��	�mx��X��ů0]��Xƪ9V��0v�N�	{��	N}�����#�sryU�qX�m6�6��v�'owN5�����ؼ�:��x9�Gjţ�i��5��{[C�b:�j�x�S��;���	��vv���jݞ�8�Q�6�nVD�v���ϊw[�n5�{Xq������o7��26͛["�0��ʌ�z�sº=�͚�;iļq��Y�/[�
\���˞ڌqk`�ي&�;�Z��^ܛ�n�B�=7Wc^mg�y���8�p��[�w<n�ݬ�\絴�j=�y�Nر۔�糃O.v�rry�6��/��=��7n
�yz-nn�|8◍����n=���եw���76�g�a��a��ݶ��C��!���z4*��'k��ݶv;�[������{O;�\��n�l�in��T.�[-s]s!�孽s�ho44�ו��<��M��el4���z�7�n�f�l�fK�ε�[p�;Q�2�<���N��4B��ێ"�n{m�Iq�g%u�ψ!A��6��J�½1���x�q��X9ǫ�nݬp`���M��e<㮔���d���0�n�G�N��=�� �nL�6��>�%�ͳZ�y\�;v^�7ms���wV�v^<] ����j��x�۹hY.��y����7���݃�����N�t��t:�f��̈́L��3������+>�)��Nx뱼v1�a�E�*a.����榫����-O�����LW_k�Π��������L�|7 ��#B������s��td�Qgޛ�z��_�3�To���89��0 w:�d��V�U�Ҳ	wK4hO�L���S�z0w��A&7sg B�_WI8�,�A��aP}>&�Nad�n��h�6�yJ� ���I���/ĜޜOB�-�����ʕ���N����L�*�"��W9�4
]8p�+�KB�Fu+���aP =m<vlY���@[���8;[+ť��Om��k�թ�gtu������+j�/3|�ݵ�l�^O���}��{��H$�ެ6c �4�a��gb�$�p�-zv	��Q队O��g*�;�Q@�s��/e,
��۪�ydę�Aע^+lD;�,��s7.�k��4�(�y�qۘsM>�g��W��)h�������x0�I�XE�A��i�;F�,��̙����p�����h����Ѐ���T *O8hM��6fi2�Ն� ��ڿQ��E	�͑�f�^o���Y�s�-�  �ز|H}�f���2�e�g�UZl�/��(��0X8��,@|+��������qNI�6I{*�$�cY���׺��Q5��ҦX��e����&�̕���]���DDYcu0~�!���O"��&LT���,�$��eX$�|��@�~���{�審fbPk�/�4�3D�&�jo�]���k!ٓ�N��@�O���-�r��(B�A3[7<t��/T���)�s1��eTu���iή�36ټws,&���/�r�;����:�7�)�ip���B��ݑ�j̸�4eْwm�b��p��7(�b��VSwBhk5,�#�����Ovr�M����:�Qoە�.w}��WδJ��X$���a$�<���t�K.�A&w���/Ң�zfb��}N� }B�߂�a-��PJW��� |��`�jx��~"a�����* 
E��s��w	����V;��Fv-�g�vݎ.7�s��l;��A�P҉��$������s1W��R�b�'A�/����N�A]�)Y���5�ii6��{F�M{z���r��g�X��ܬ�&Ρ�OU%��EPI����iݲL���	rk{��E���d�V�,�H$O.�d��NA1�EO�ǧ�Vs��U��I��"|uVva� �\�X'Ās{)SBu�u��+�!.���\�0�<�����A�Yk.�w-rS}%98`�n���pX���DћOoܩ��I.�Jڧxꨵ1s���C�s�]�%��U#���3~ݫ����y�I�{|��,�0�H�w*T ��}.j���b�c��\2٘L=��ء�c�6-����|�������P��R���Zn�m��j~">�,��m�� ���,Iw��P�9��-ﮓ�Ӫ�>3�Rsc(�Y�S��� �\�x�O���fo0I��;��dtk3wE�Q[�g�>7��,�V��,p�5��i6��=��I%�F�ۦ����|H'��_��n�V�mL���l���,�1?e筒����f{X	�;Ԩ��/��O����f�ee�={�~�\��q:���M�:�|I��y�ը�2tv�\n���X�;�U�Iٽ�D3'r����{K�Os�1Y�2+��h��Δ&W;ձL]q.�8�D<�������t���!���᷻,Na��,�w����-j�����[TXX�/y�i�����bu���ч;y���wh�8��\��m׶-�qo$n�#�=���:޻=�.3�^�j }�hy:M׵���Z���k!�s�����[*���eqO=�W'/Z�ƭ{R��T�.r������d��g��Z/�[��ܦ�Lfݹ-Z�޵�e�+tnz4[nGQrh"����:'A=8�\t�W;l!��ۇ�l��`�.�A�+�cUs��=Jh��ß��v,O�W,�`�;�{0�s'�J�x-��~'ă��X��0�r�wxN] ���c�Vߩu�b�A��t�	 ��d�ݛ�3ǜG@hoV��՗�^��A��#����y�j���D������\�����s18,���M6���~���qK'�����TV�Pec�&��, |��Pk��'�ˬl��O��1���˫�6��*��nR�s�s^��{��_?oE�zy{=#k�T(S���|��H��oɟ���δ��j��-M���j��R+��%�Ð�k\ϳ^3��
s�Lqssֿ�]�}��"#���]V	�����H����E�L׉���ݺ�i�PM	"*I�J~ؕ!G+H�T
����' ����Ժ�Ku��z�U�Ir%�8�Z�wW�7|&�6�e�|�M��7ҦX�F��H璐]�:��ʺ���$����PwN����k���I�Id�33Q"�m��A>eu$K�"lQݰ�V�	;w�<Ir���U�:����Y�����v�n򬭧�w��O�[�d���ʄt)��r^�޽�ϛ�����$%�js�ZI���x�N0Q�X!n����<d\� l�d����DY�̞|ua�V$H&9'q�[m�����ιն-�����kv��6����Tz��P�4	�����c����]B� I用]��z����#t��O;����� " Q"�7�аm��"x�C��{�'��	��g����w=�7�w8"��*u�b\��X ��y^�e�����䛈�Di��k��u���,nb<K�sB��(�2��z�͙����wJ�]�<	hTT��z�Z�\���CN(���S���2*����dx����uw���7ֱ��W�MF�&z*���� 	��,�Ov����w�KsDTc�M��^jtc��Ex�2���~��s+4���� �ۡ`�����!�g3FM�{��4��9DZ�XA����q�s��յ��%��F�Kj�U`���������0d��-;�~$�����H�yد-4֜Yyh�-��`�|S{VO�V���Du7iKq{�{���z�2nvrۡ��|	�5���/;g��,�����M�����X�Q ��}K� I'3��O�.Sx�uJ�a>$�`���س>i��BH3B0��皪ῥ�������� �ǋ0�]
���p�S����9���Ef,SZfGͧ�o9q�T���HE�yi�S;uF� nム$��id���8�
�8��X�yb�_ɞ�X�Q�p���*����_y��Xuuа\�kى��(�2��Y�s�k���wp�����I�Kf�(0T)msp��h{W��nwhx������t]�*��C�6����
O:1�a��O�z�����q��I��X$elp��"Uh �}�����Q��I��L���kKM���&6���ˮ�'m�h�I�`$��R ]b�z.Hd�ɞ^�߀̧�<�jhA����ü���H��B���nb�M*��,m,Y��ˮ��BbA�",D@�$��˷..��"���J��I%��m�oc�����&׽�d؋nU+��*����ڢE������ X�6S|�  �UW>Ҁ�f�����IM��W�{`̎��皱T�����3���7lÏ��=�n�Ҳ-��i�^�>�8n�d�[��'+gE`�*�Yb����}c�v���/Pq����3g;��.�i{rY����۳m�-S���1�y���{b#l��'�=@i�.�t�b5Ǜ�(לv��h4vwX�_n�"��u�F��v�H�۶�R7�����.�Sr>��ЂE5/�k<���7q�zMxR���[��+l�ś8������
���R�ۇF�/���N��\�.�/��ݎ��w-���Xy�p��3��;8/NQƫ�KZ��5��޶�"��r����$_*�d�T��'�ݏ0�u�ߵ�k�I���8�y�?]�i��QL8�k/��sy�]u�!�{ޟ{r��z�z�quk��(�S)\ꆒH9�v�v��.n���$)���]�$�_)�@�d��P*��������!�r8Sb>3��,�I=��� ��X:)����9����I�"(D@�$�ۗpA&���ё;N]d��� ���l@>'�ݫ v�]w��}ߛXv&����!d-�82��]�m�����/�V���G~����'�Ȓu��b�� �PI�o7R��4�ĭ�زI)���!�4�"fI�7w��rR�,�)ʝt!���ףb�G2��LEJ��2ƍX{�Ų��ϴQ�3(�99º�+�������a��Qаb��m����>��M�m�����Ob]UfOf=H	Z"'A�LMI�4s{sv ����y�Ff�Rq���o���Zo]�����5�	
�b�U�����@�͛7�Iۯ3ĀHu�F�o>��)x��;pg�B�U�����:��a$�
��*x�Шz��}� �k��� �t[�_������'qFN6v��S:�������y��������l}��K��I8��y�ƃ�:!
6�������׃!���
"�ػ����G��rtݼ�� 9��x	n��/���Q4'<r��@@ �ǽ�	%���S��g�}^c0��<��_��GL�L� �7�0��vWP�I%�Ū�S���+��{k'oU�L��*��e.m8�Į�x�:*Oys�WX���d�-h���+fĬ��ޡ��e��Mc��Ga���hfmv�^}Ll:Z,����{7du�����o(�{�0�c�@u�ɺv������ye�Ů��C��y�7�Ʊ�ۊ��5��]Z��Y��������c+��*>���a�;e���*ػG^��s���C6vŃ���0˧Z�jv�������7��,��DQ���f�5�mP�l�)�ٻb���3��]��4)�B�ƛ�ۜo�HG��Z��6���\.�5����0�
�6���v$S9��9Û�a����E*{���L:E�:��a��Xk:��	Da���p����jT�ɸ�OP���&D`ÒĲh�f�t����]���uqP�7�j���:̷Q蕉�̕B�պ�y���wjv9W���,=�`ݓ{̺%�ۗTB�����y効��p[2��̰fM|N>���^ �{�̵:�?*+q�$�vdS�u�j�Lí*�dڊp��Uľ���Rn��Ef�������u�7�4�VV��n�
�*�B�l�SIM�J�t�u%����n�kf�e���V��]�&uvQ���I·VlO6d�1�&��f�L�kE�wܫ�s3n������T�Z�I7x��A^X�������1�Ն�fꡑsf]�/����a�eJ�I�o��!�(.���s4y0n��zu��=u�u�����E6C�XSГ���+^��1��0n���bP.��H-!H����Qe��vE��tGg�oj"�f2�.*;.�mu��y�7s����9Μ붷Qr%�n.;�r���9�3mgA�e���;:�\r��Iq�$rڲ2,�:��;���3:̧+3�.������D���VqY�On��ˣf��:�bR�苳��:�貰��I���#���:;�l�T��r�IDGr	�!�gf^xqA�qt@q�Ӷ�#��gBGJqQ�k��%�.˨��A'sۢ����܍�(.�²ܒ����λ(�����9;���lq	�ClM]�$;;Vat��`�r��N@yVj�69�^��܏1��O?��@R݋$�V���&uŬ����ڶ�����9��8�S)����i6�y�9b)V�cΎ��ȅ�Vg�s΅�I]�����_W��L�@Q��$��
��0��(.9��0F�#f�G�3Y��H�����~���*ѩ������a'ǧ�$�W*�~;J�oM��Hӫ;V�|HS�ŀ_{[h7�У_vw�y3�%֟���V��z[�`�H+���:���骹�]U�O<	�7�4�1@�&�F`�b�$��d�=��p�$��ky�/NA9�U�S��5��̎q�5:'*�-:MԹYP(L��,��6 ���q�Y��������]�^C!��{�km.49*W����J� �Z��_<g)*�-6��9m���;QZ~�P�[�\l��+��T�w��t*l�AJ����ֆ׳y�K!�e�o��	��X#R��=��0�dJ�&/�x����6a$���" ��kf#� 5px..�&�6Ltj���S�����'*e=�_X�H#9�؂	��(�e���4��Zm��wٽ!ޭl&0V�,�˘���Θ�[g��S �n����	.�5;F]t��(�*��9AEج&��dRz�Q
~���x�v��e����'Ϸ`%��H�b��T�3��P��OϹ�z�kns�6A��0*���Ɏ(��I�r�! cd��R"(�ϫ�^�'���`�U��K���p�$�z���]�3�/u���e)��D"(�����љm�N-J8�+o��9p�nj���̱�ͩ��5u��[�G�]mkIM��Z��S!:U-t"v �ځX�;p�<�\<8�5�B�=���q�\�c�7�;��9[cF۶qq��8J��a1�-wT�;�S���1�'#����=v���a+�_8����˭�k�f��T:lys`:� ��1��M�qܳ˒Ҿ'Wv��lg�b�g<fu���0r���Qoknt�h<���a�g�&r�
0��:s�$G:ɩ�lĺ�[z ��A{n��˺��i�/'f�������Ǵ(ցq��߿�}�g���2`H��*vn��>=���'ܺ�X83��(�ڪ4(�l_�wwBŜ�p���*@kM���NK��	#:����_� ����t��>��2�vһ]�3���{>������m�c׋0>Σ�}z�$���X�H�QD7�^����Y�Ӝ��ۻ	�s��J���B���${]����%a���o�m>�z9į��+v+V��N�M�$r�������6����$�;Z�Ѕ�I^����1u��]���y���j-m��"�R�؉bNޮy3Ѿ$T��32>�ٙ��j�~$�s��՚��`�t���}��I��͓��1:��%�⹉�nkC{ߑ"���U���T��j�9X�X��2�g"�\≝��3tA��ݙBE+SU�c9)�|���S�|ʸ���d��G"��|0�Ot���H9�v�k�Z�B���k����zRH�!S)��Oh�m&�?z� ���<���Y8�@>�~E@��w�̳x/�C�7�ظü�^'�n7 �p��z�Vh�5f�����oE�f�t��4�G�N!�}-A���l�ӵY��uW:�깿�A��n�v��1Dm��9�gR���n^�[r��8�a��Xһ���v}�94�S;k��������V2Ƭ�����A�t�'��v����s}W�Kx;_c7���^�)�V�jrb�ݙ���fa �n1Wx��������Y�%�1qqsiB,�Ϥ1\��ܬ x,݌lz堨�6(�=�������-�º��U�ehsAJX3�XU-H
�tn�`���^,ɬu�Ip�
թ�-v<��+s`����BnQ�;[qy<I �s� �Ge����������B�SKG����s���W=t�D��s��>$�e����A=�K��_u:���m?os�H��=�+nҒ�boj��>$�]sf�;���@��S T�������֨6ב�=MC6}8�B�6�(�0VQR���u��8Mn�^�	��\{I�[��K��/4yZ6���ϙ��|2+/�>$�͗���wA��kw�Mi��k��~�;�"�ƩIl5���`�E�>�����6��H,�9�MJg���۪��A�Ɍ�K�H4fdX�{0g�c�X�@'dv�5���Vv,(���f\�2.{a��M����a��N_��(]�u3`��o=�ēҩ�$y��F�0:s�@�F,�5Ʋ�^�tr�Dh�c-��A]���V���9G�+�2�yNX���U}&q��-LE�8���!{ە2��'w�y7����A�B�SZ��zm6��7q[�4�+˘�T	�s=����~�&�����ѩy�fߜS�*�GoPll��Jv���ki���rnL"[���̦1���`�2�U&��LM���` ���`�>��'v�hi�����`$=,�*��F����u�HA*�ͼ�j,���o��*yذH'ǚ��@>5��}��JOo;�m6�;�B �)-�{neh)�ZDP _$<�w��6���(,P���2*��yy�"}խX����32,���}&L^E^�T�d�A#��6!�cȷ1�N�GQ:��d�ud�D�I��=��$4׵��fl�vZY\���Y�M�~'��g�Y=�2,(S�m1��qh�j�ĩ�E�4�i`͛en��B�S*��8�*�>�ԋ0k�~dc7LՒ�;�b�ܣf���9����ZDJ;l��Y�\i2��;V`��[��ўwA(�gZệ���n;n��8���s�qi5����J�m���:	x�$��ׯB���;����2b�R�\4�(�)�:�\%p8M�C�U������v��wt�8[��]o۫Ab��W��q�����<-㌊[v��`���͢�lf����ɸڕ��78��3�����s��uEm��q��<�n��8�oa �Wj�l�K��%����������*��o����tr�����Z�=�kJ���~�k�<�P��@�Yf��{usc��w/KN��P�	�	t�Ogc�Q�������
�_��Va�,�]�ਓ�|��I4�#v:�g�ı��ZYW�M�\�qf��u4@����1{�֕.�,������y�* P��y���]~')sSaamN;� �����LK���]��=�1@P���T6oe:��D��6	�n��@'�+�Xƞ�\��g26��kc&�;eV���@sCQ�gi��8}�G��1pX=_���ߙ��dT��������$�n��|H�]b��X�V���
�>���0�9�Srd5	ce5�ƹ�-6�����
�����4z�Rz7H��Lً���P{&tl�8���T�U�2���D*A��c����Ŭ��1[oL��(P��fH�]~���릏=��{V�e�QM�Z+	��7�f&��v�|�m����)+�Ή���@�R՘I"�q��a��>�ǧ�zw	Ï�]��{ك'�t,�O�s���5�^��#Ҝ�����
6NX��������*T>�Ӗ"�E^rD��v<�|as�,�9�ײ�e��?w�)�?'kTU��c�{�b��:���`8M��=�q

H�J*XJX䪵V��� VQI���f,i�o��I6��=�a|��_<���7�$��|�����=�t���H���6��;ט���C��W��H�����yW��/����}}�t�L���B����F��-|�m<����ڛ+�38��
��U��"bd�&ITL�Ǔ��J�[o��ӡr�E&��s7()Νɐ�C}py�\�#F����q�2;�]�5��O��;V�i绕i^����CcE&/���ޓ�`h��
�E�P/{) H-vW����tLWD������[xm�a�EX�T��o�y}���?>���[�f���%'�~ �z�{0x�&�ɳ��o�u�F��Eb�`� �.��v^�S9��Xz�"[j
H��ȋ*�{˿,�Rjj�{T8�NsʰH�����sz��J�wgh/	ֲ�ĀB`�H	��5wa|�j��9^�&p[����I�)uaH��y��ꬍ7���O��j��-7���Y N�.'왾�I��x0��*���:�X�1+�<禴&�}��$�}�R"4KFS^��`����N9��b�x�>;[���S���f�c��yf7�E���^=��ꢒ��e���b�enh�ۣ.��r�t�%��9*��
��yj=� �����p��X��ۡӫ��|I�N���"��\�l�~���dev,�I�f�s�s"}0��Q�p��^��ي�`.�#��О��'Q�X8����ǻE\b*������^�a�{���)�}�v]%P1.n�;���.���9b��^fϷ4R!����ru ��{׀�_U3`�W[qr���#Ȫ�Y�>!p1�Ѓj����ƃʥ�'����9Ub۶��i�	%��`������Hs9b���Y�����=��C'�^%�I'�W �Nn���W�0�6�-�cԈ�v��s%��~禴��q[�Vb�g9O����{y�^�$����$��HH@��B��HH@�y!!I����	'��$ I?����$��!!I��IO��$��HH@�x	!IRBB�D���$��BB���	O�$$ I?����$��BB��$��	&������1AY&SY��R�K�߀rY��=�ݐ?���`�`P@�P
   ��U��EUU    P� �JQA�}�J�"BI�BDQT��ԊR���G�W`V�r�]��l�t5����z�8��vЮ�nm�����x��P�N��]j��iE�M�4���u��A��zU���scv7a�U�h4n�b��xyP4҇z퍱���3��5�rnu���< .�6���d�]��HQ��-5 $���"����AG@3�u@tiw�����CF�tA�P(�x�ȡ.=�(h���u��\r�� �t<��: ��5�U:�|     jx�R�����P�#	��4S��I*�M4� &F   F&�i�UTj�  �0� �5=��bT�       e%P"�M4i���&�42 $�dI0�F�
m&L��Mjm�<��G���PyX���@=?�d��P@�?����+� 	e?�,,������?��(�����ǘb@!P4��T N�6H�# ��� �����W7��3�}��]��Q ���6�N��ΥG��Q��p������P"9~��2�
�.��J.Ë��,Xnc􉦓B� ��i�@X��Q��rt�F��j�y�xEP ݜ1�U^Ԙ������~N��5�\����d���x�i���ˇv�#va(�r�o��Y� �bL`���V�ӹ/+�#�W��{�nJC��b�*���ӷ�ŗ��8\)��'$����R���3!e���n	�ιp�dįpֱ�z5�. �P�t�hr�#��!ba����@�Ɋ�ǔ��O���z*8we�3��b{��@m��C��o<�w����ȝ�q8���s��;�E�Q3EI.�{tZ:��/nIU��<��=�_�]g]��ۃ$�3�ů�/#��W�kgs�A�On�-�:#�-�d^ҎF��N��m{�ͪ�m��N�F�a�;��z��vν��K��h�پ5
M5l\�Ɩ2FY��q0�T���D&�G�Q���hH��&lחN��g熉��ۄ.N�{���7�ނk�)��hՅ�d�j����9:Q��Ӷnեs����`�L!k�0׫v��	l�=�i|�y;;n�mo:�u\{�w 䌱�{K.*����Yv7���[Cy�Of�E���p�,,���6-lc)�=̳�Ǯ�Ѹƾ艹�шlˮ2kÿ��Ś�s.t���9�Cy�μ�PD�Y�ZHz����Ȇ_<8�wq˯F*H�e�e]Q-,��u���R+0��Ő1�Ni�P,B����i�r�q�nn�ɠs~9HKh��kK�)�a�Y���N�Gl��$2ޅ��&�7x-I��Zs�����.Q�]��-u7�u���r":�!Q��q&�96��4JR�6Vk�~���	Ziˢ࿝k�-�U�K2⛼e*6�y�d����U������%��w`yY��M�ٯ�n�.�3T�>C�k�a��d�VgE2%����x;ԛ/7���ۀnPk��9�[b�;�#���,x���j��;:�O��-g�DWH9ͰFI�woR{�r�"<-.n��j�e����'�rX�FYǳ���4�7��B��ށr���r����,�`��o�VT1��z�qM�dMQ�#����m�j��#bws%c����=ڶ�&��'~w�
e{㝡��gGJ�\�Z�ˆ-��kE�qA�� �����@2���;;��^8�4a�[T��k�1��êI#�t-^,���s��Ɵ+rIq���.���s�H�x�M'ZOD-l[�����j.�@4���K�N�4i3b��1���+M[^��&�j�0]z2`�l���$гe��E�����4g�Qֺh�
q���nB��'��̵SѨ��'L��¹>��op��{W�N�t�`��Go@{�t�wV>aGM���i��J�W��s��M۱˛0����қ�޻;k� }�d�Y9˒�d2d=r�S#c�����ќÚ��sc��5]�^6����K�/m�{��"9a��G�E�S����&�\׺��3I�O(��W��K[����4��L��F�E��1�d�0u��V�Gb��1�9j����د��q�&���I8��[Q���xe���1bgk�� ���S�Lb� r韤F�a�������n-Eȗ
�j'pmʑ1D��#$�G����s��=�Ŭ�I���6�T���%�L��,2���o�8&&�$�1t�&
����a=�v<���O������n5�u�u�<�0ΝqjQb�^�of���ml�:�(���EQy('��wu�&v>�j�U��53\��</;�M;Ceѳ_���/��D�ϻ�:q��-Ab�{�o�֚y��-��� (X\�"ӗWA�F]gQ���X7�/`sy��5��Y!X�m��.ni"˕�t��j�KD��eV���p��{�`;0�xTDvLzc���	w鿎NOGRœ(͚7����n�p�ڇ[7�Z�q��ۑ���i"<%��{���K׆��Ě&w����]�nMh��P���;ܻ���tÙa]�m�n\;�Q�09��)�'�pl�Y)�v���
i�[�`�Iڋq.�VFU*�-�)�`	(���b&�,z���7��oei�mrɇ�yy��y��c'����9݅�:0�3��DFL�m���6mÂA����4� %�/�okq�9P�}?U�8�1��E}����4����(A�I�I^���,w��(��V�
�*� 
��! *
$����� B�5A� 2�R�Ȩ2 &M� ��`2����q�C�m�.�(vp,�H Ƞ! *
��#�y���']���X�N��  ����n0�(	�qd@��j  �G���_��W�3������K�n�D��cVdn�9vz������4���D�7��f%r׏�M�m=ЃŚ٪�ЭZ�J/�BC7�֩�04y�)���F��\��st�}�Y��7"<�ۤw��:b^�k�rm�P��c����BpjoQz,K�V�T�UM��[B2��s���{݈��}���N�+�0U�=<�� Ѽ�g}�q�8��1N�l^(��5�W��/<����e�|�o{N7=D��6Z���0r�K�Z����e�l�}��os���K�á6����J���"�-^��6gt�n�Ӥ�[}>�����`��TS�.	�h���XD(�Q2��T-��ѼBpQ�d��T��'�@���#�죙�ǒ��>[���<1�����V�ʬ����\�S�P���Q���nn�󉄎'�vV�.�ē��2ά�2�
��?{)X�VA����ׇ/0��od�N%°�ڍF���^���o� <}�P�{���Z����A�T�u��s�{Z˝�]7}�e4y.Ζ��?n>��ٷG���,���%;ۓ٦���L������)���L��A��h�=}��k�e��A(��{���3��Z�W���&�����}�ι��,�L�׆=>�s����_3������w��HGy��b�����=���^7�=�%���ץ����C�7%�{�=Z���	�:ĝ�b�������F��Ş�u�Q�7_bч�]_� �ǯ�-����qo����U��q<��)���Ð�Eoٻ�;�����#���<�C��W��z��\��瓧����%&����,t84�k�hRp��eX������%�=8�pz�m�]��n����s�o���m��:z�61���c��s����i١����m�m���=��;�SpV����V��9 �u�.���᜷v��\��g�Xnz��;��o��j��-�uMm��,����_�u ��:�-� ��Bi\p	z�9���շ��@ɝ��Ãk��� �d��c-�w�V�����ڡ��f������������??E������2'zas/����r"�-A[�I�w����H�5�+����ԯ��Z3�榯+�ay��<X����l��O}��<�JȈk�׏�Ob�;<3�]��W����M���T��ڿ�ڠ�Fv#.��L��\�:5�4\I,}�y�1xA�@�}R�ƶS݈���ъ�S��piޞ�HH��&Sv�X
&�x]���������<c��+M�#�˼sq�� ����{�}�5�F+�r��ZjS�[�q�Ir~����
��6Ks���E3�0�[��L-��3Tu4v������\t�pD�U�'�q�g�~B���U8��ơѽ7��v��01pţ��۠6��{ݯ5�׷�G�y�~�9�:lx�ܾ	�
ս�����6��`Q�܆���kx"����>���I�a@�\����.�f����*�����n�4�'I���:�W����NN�~�z�ib�^=
h�@��n�T��p]ES�����7Ͻ<K�#4��Y������>����%�;O����3ڮ�vi��4�x�{��8u�����u��s.�P�5���+�q<�j��e���+��� g�M����bC ��YY�nA�g�r�B���f�+bv��������ӭ�q��A�Ź�c>cfOF���F����N7e���;��Q�SO�W�}o�cb��A�VUPٻ��$����K6�	/Q��;v�6t�+f7��	���8j���4�ݱ�3�/8*��cp��5WA��[	��˥S� �>�����x�ѸZ:�J���7�y��~�m�"��C�<�6Bqm��m�0��8XbP�a���ú�[�`���k����Gӎ��b#P9{
���ٳ���z�^������^��-�S����/P���HJI�3Z웅��K�]ZosW�đ�m�+��T����zC������/$��V�͊�N&�19���T����	����g���V�N7��}g�ꆦoq5ç{}��9Lc�_����G{���qњ�H��
�2$�uh�RС�YmC
.�Ӓi���a���ޏ���y�ηs��德�p��C�e>��.�g�Ʒ�]*���������}�Qd�ׯYA�c���]�o�+�Ūp��%���xs�ϣ�{M$b.���y��,���l�z���s�|�  �!"I�!tSr\dJ뚲v��y��kܩV�jX:�k��3kt��J͞-{Z�3�l&�8�FK�,pXs0�6�����[q�CSe(bs���ט�V�
6��d��c\�t*]�Z�����=i�d`Թ�{^#���v�i�.�:���IY�E�P����mÚkS����j�G%�f10�nĩ)��#	��.˶�0MɗSh� �tMe�Jj-mѲ�P�&m�!L��C�5����J7MP�1As��-��B�&/A���ڮ̭�+�P�7Q��d0�
$c-��,B��.u���� &�S�msj M�0p��Li4��p�ƴ�0��mP�L�dEPr��x�a4u`TL۰	�Y�E��6`٬�䫂��X����sr�6��s�Z��V��{CK������j��0��lE65ڦ��lnj˴ѱu�8��{^ʹ\k
�녚��&`Z�K��1.6̩ևdcقV�H�vXˢ�˛�/]ZA֤�h.CT��R1��k��G�AGX���ݒYH,���T�L�]t٤�%���ms�����6�.]�#�b��h�H��cu3iA�0F�2Ł2j�����"5�ں��ٲ�eWM)5%�i���-�KW<��`��+vh۲7v-y���[eQ���� R�j2���8���)�9t)��u"�5���ZL�\g�a&&!Yr\f3Zb�؊g0�Kc���sP�7v�u�����z�m��t%-4θ�	��[lHD�.�C ��$r�&Ե��`ɴi�բ���:��0���6�[`!�(���tÈ����K-��u�<�
V�mt�h�&{0�T�/:�%��Y�����c,̰�+��iV�[��	n�΢�Jgk�P(\hȕ!�
Yp�nN�v�lF���酘��K�RY�4��.�j��a\h��r�J�m��iIl���i��T�-@��[*Ļ��z WJMZ��#�B`��[Y���T�崩����b��kn��ԇb�eH�G�����v�_'*SA�^x8�R�v��D՚0�G7���9�Z7��)���P�[H:��3]����5l�+l�irT�6����
XL���X��ia�%�@�j�mB�U)p�@�!���0���kx֮Q��u7e�R������\����b[P!+X���0Pʳ`i�b��h�ģK�ܷR����.�i�anVe�3��4�Vmq�7=�B��ɵ�A�;�rSj-�U�Gt5,���ņ-Ŷ)nr�� ���6٢:^%��Hb�nnB�f�G�r)iԡ�=k��er����[���K�љ*j0iIk�;]B��k�f��j5IHK��e�k�FY��]9N&�K���h6ݰ� ��ite兲9[&vK��J�Z����F�Z��5�����l�[�R���5$ɫ3�5�����m��P��D`�Z�3˦�6K.�V\�K���Qsiu&qe��X�Qrb���uFRݱH�r�������v�ȱ�-��Nf[v�%-���Pn%7,.ᕨbPK]Aj����j�-!e�����Ȼ ՠ�K5�6k�{R
�:h�̱�*��e�
������nQUUUp�3��l�	r�h`͓%hf��T�2�˹k�3bh�@.ר�0�"�"m(���o�6���gO6ٯ]����U\�sFP�*�2L*�Z�t筢���Zu�2�T�Zd�U��r� �J��(�H�"�_
AN�H��.ԑ �́IDP�j0�9DN�r��-T�f�hY>�\#�m,��Z����Ї�#�^�|O���Ӻ�`�d��2P�]6�X�b\���iDʄ��a4�	��G��a�����aMj��ZjT%c.�gJ�O�޷�P�q7h6�mn��Bכ�3�E.�i�X�րؚ��u��i�e�nlV͝)�ZbV�@*镊Rb��n�d��Z搗8�5��Ʃ�\�1R��"s���cBgk1iRj�H]K\�����%���Q8��F�6�ݵmb�a�j���]Pe���Mk1	aQ눱�m5]jg,�j0�V-�ѭ�[Vmr*Ŷ�u5�"�ه�sH���qLD�[-,:�V][(P�\b�Z3mj\a+�q�X�+!�E��ûϝw,r�p�.s�n�����W�K9�X� XJ�JTkE��%"�EKx�YH�e��~ǟ������"���|��$_�:��u����^z�$^0��N�5ؒ���a�E�g۶Đc�Y��;_�������8�d����fu��D�P0�IH-��Ee&�Da��a!P�3W'��Mb�b�ca{6�'��)l>���~h�yؖ��~�2�8�K|���N�s���4�!�����4�1X �!��E�WZJ<n#R0�Q 宓b4�x��o�N��D�Է6�Br�m�{ǭ/����.x�n�16YQ
��g��AJ �0��@�� �95���:�'�uL�&	q�ϓ'��l�
��?i۾�[��b��l{�Z���A�7{}z~�A�����S��\G��J�3.�3D��*�Q+>?�,fÛI ZJX���3>c�f�5���uSh���}�}y{�L0I�c++e>�P^u�^7αI9,3v���cM��UwjӚ:�~�A�H���$�&FbV�P��$r�$����[dEOD��8�S�c��3gga��Ń2P���=�͒:��UU<��]�����B	�a��d��ق�bж\���]��y)�e7Hh9�3�Z�ú���	9F�ܻpC�O�G sF�~�86�p-' �Az^U^^fPd�At�.NF�i�$��'HD�8�ILu�	C����h�#��$�Kً�j'ѓ��틅�iлEe����;��N��MA	,b2�3B�1T�уA1�6iİ´Jݣj�k���jX�]�)��Ky+��V�DV9���b ���7[Qhq'O���1X���>��	*ש��$�D���0�.����	9lz� �sP}M�=@�3m�/�~�Q�*Q���X��:׫P���9 H&5�F�YJz�8c��,X�>���m���0���5��d�ъ	��UT������pp������r���(�y���� ݯN�%ʢ�E@���t����c��%�P:Z��=i�w����f������m�I�8�%D���p���D�r��@N�f ���0UVw$�3��G2���"���E��T˛^t��) 8ݨ;����G��J�/��wר��=��jv[��(��^�1����T.�2A�l���V"��j�J�$�L�M$Eҥ,:T��	9�p�F�躀��$.��U��u�A�]�Q�
�!:��u����(�+Z��b1W]�:��Ij�@���(@5P:鄡�h�����}ul1��
��:�uFN���Hx����rݮ��5�x,�FVV){3cC�V�R욺-�@� �Z*<r�&��Z�#O�W�U��p�Ow�~S0	]1˵��]�מu�����b}�޵�����l��d&�5�D� ��:��˻䜍HY�L�^=&���	�	K	�1���Zg�I��#��U��8�6���5i�I�YY*4Aw��{�sr�Q�`ⶉ7?��6=e�"!��Kp0�-+�K4G�6�U4��Z�lEΚ#-��lK�H�F�:�ױv�,%�u/D[Q��6ꦙ`Ã
�8�P>+S#iA���jșL�����:F�7M�sP~"�G���!lh0��l�% NJ�Y���J�Nx'����%�s���B)�<�hvS	C��(;m�I���v�D{��#�u6ו�C7���S����I#
u/v�B �A�X1㊎�",-͞��b)��$�Bx*)T�R�)ek���/'���A8Q �ΐ�iږ^f�I�H��$f�
��!������&��Hx�ƞ��p�껊uG�rf �H�2�#10Tkߗ�x13I@c�X�<���v��c�#�m�"I�c�t%3�y�vQ"�2��v����c�p2F�`�L?�%{��[�N�n�|K?A���~?��)<{�>����"�ߚ��
�uoM���g�~�?gv��Ε7g��طa�N8�T`�f%��B�ܸ�TE��h�WF)��x���{�׭��wg�Pxͅ��DC�}-�Cӱ1O����N4zvt�T]�^�{�<u��O<��ҭ׽�.�<��������}��V�3�:��7��y7մ����=��Y�cހ_?+�o�zr�ah��S����}�/G�n�̖�6F��qW� n���JK�
'P~Qp���G�T(TtIL�:vA�"UM&�� ��	5C�T��#��eP�QG.f����hp��P���s)YGCz��D�EI9�8G%L�*+�*"���P9�P�*#�(%rR���k�J�fN�L�W*��>D���*��}?�?��ϔ�^�pI��F\9m�	�LrD_�y�1N��e�K����DB�3$�JR�	V&�D1q�v�΁��:�����y�#A�5J"���a(a�T�&� ���"'BS7:�$i�jU�gk�L�5 ��<l�f��1h2$Eҟ��}�H ��K������������t>>�V�bF��7D��8���_��w��g�\�1jٴ[*ۗ}���:8T�I �^�L��p#�8T�_�x�m�]���0I� _{�3_U�K
Q"1�B�,A|��w�%S��8CH����u+c�`�dǎ�$m'�T0Ť5�I�bFZS��x�j���I`��MLa�4g��E��K.�B�۶�Z�M�%P�D�jl���V�m/
�0T�%lt3[F���ּRMf���,׈�Q��bĬ�q
! J�,��o��NF�NS~�L���t4�3��=@�<��'c������,+��L�ٗ�:���cS$���&��j�=V���Ȝl�r� ���v�έ	UT�aE��Y5��Y�|Y�vz<﹄*j[.x������2.�B�c��Hcߧ`;3�@�|����5y������W	�/��� �ּ�� X�wUP1�p`��O������g��ih8|��V�6�;Z��?�����_��EWLֵ�]�￳o�������wg���D&3��
�ሡ.'�.��S�;��+���SF(�2*+��ʥ��
��>	�f�Z�G׋�w�𳙕�Nm'� 1�������;����nɳb��͹_=�\��H��q3���+S1�:U,�O2���29::�J���Dι�u�g����鮟S����>�8df<��s��"�G��+V%&���&�N��Z2�;�ق��f�@&�`���I�%��R�5eK32�1��, :�˼I��lb���]�o�!
ϲx��#�	Sϟ`:���Sy�Nb�S�3LV��sfB��;����u}-��-u�^R̎�r]��.���6�P�J�n	��Ě������ձ؎Ը]���D����z��`R�U[Q6"`nr��W>^��I�Fe�ٞ��B;vc�DR�|�9���u�����x���6�~��뇂�-vC�~��/:=O{;���Ϗ_=��u��I�j�1*���p)�\�/�T�%= �H�է��X�����k1���e	�<wg^߶��������GU�;Ᾱ������*��^��j�6��xL���d!�P���̌΂;�87!���CpZp�,80��9%2x4`U��S�cR&)�}��ה�oMI�!ֆx^T�����ؑ�D�>A�����򯦗�}3�����#�ߏ/I�M��]�.Ax��L���^ܽ�,�%�j!x��m_p�{��F����|7�IL������L��Eַ����<�����ͱ1 �]��!Bӕ���{�{L.�~���}콩�%�&��uc������"�3�x_�5�s�]�~�ԧ�o���%��֠],Y�`�;>+�����O/$a�wX�e�E,˻��Q�Q�^�^�7��1v�k�N�u��|�y���L��^
:A�<�t����O��H�-�L��ݍ���nhi�ʆ�=�
'^�MC�����@���{���Z��i[���L������V�;�gx���g�~;:E<�i�8�g w�����g�S��Bb0�Sd������� ~k���Q�a]8�ib*��
D�j:^c�p'��^Ӹn_4Z�P���S}������/5��/~�t_���>��;v�[�tG�c��3�Hs�7ݮq;S�s��%�#���x4�N�[��8�Ǝ���(���M��#0h���`B����'�b�r���8Q���"�Q��k����`�QP�W��"�X�*�H���qP�
*��������E
��9ȉ$#0.\N��>}�Q�(���sD�
D$$r.h��E(�Р��\�VȠ�W"��e�* �Rg*��*�Ro�x{�x.��X$�0Zm�C���h1
Lv7\�vz�
;JH���kvDإ�Gi�-
�^���XR��h�8+]�qFi[�A��$�a�4�L�[ST�pRm��յ��T�咖é�oZ�ah�\�1�fҼF:�3@u0La�P�R4�VZs�lX8	`<�c�[T��oS�l�� ٶ��Һ�K�ki.��Q+���kx�	ke���YE�h�e�C2�G3�cc!ĥFXZC8:rgDkq���M���H�BGW[f�ؕ��pksl���������+u�	HV(J��x2^XQ��a"�g\�9UPs��m`� �~;�}������CW@���*��
�1��K\SnL�Mz����/��9٠]n��#xͬ4X7~7���f�a�ٹ�Wie�4w�y��h�$�_�y�5�Ӵ:~¥�TW��BH�.������!�\s�uղlc<w�Ib���[�]ع�FU��[��]��˪�x���Fq�9��P���Sc�]�/�����z�'�����'{���Dr��GV�fn]315���섶���� ���wÍ�c�u�T�/��?Q�C��>ǽ�~8s���?RL��A��I�ǟ�^=��|��,M*�2ͧ���������[�1k�����v+�^���6��':���W�jGZ�'�y77쏷"�u���4ǆ�m���xx{�݈\�,9�@����I�k��眬�9������Ԯ#��$"(�O�@���orK�/\�G������W~�r��M/�m
ug�yیW�bNqE�\��WU��]/B+����4ow�EP�1�����u}�K}���V*���!n�5ll��(0�E�
0�(�_VGU��:A�5"�'։ΚvY2���gt�=����3�3��m¾x.т1�%8�?xG��I����<?k9j��{6��1l����y�"z��]�t���}�2�lb�s�(�f�f�:�%&�:[n.����ks�f���3vA�b2�廮f�)/SR�5�Tr5�$a3��0S-DG_q\�N�e�������U�8�{�7�Voȧ/�h��.��$N,ĳ'�O6����ER������_y�W*��ѱN`AB	f Æ�G:�(����/��x׎���[��ka�0,��PЫƧ:�Å��"ԓ&~��t����b��ۗ}F���4�M�&�E)>�>�����#�wu2�=��}|��pd��ǣOۻ�h8˳���6��]u��z��{�z�qU<SÞdF,>���-Ps�K,��g�u˭�_,.��c����mX�#>���>hfY�ef9��wʳ���Đ��Ou��`cY���Uwu�n]�����av��7j�����?y$�d�u�-$kvD�W������
�:�auJ��1d8��) ��	h���P��q��p�箵*�@�Pqq��B"n�*�X�H�R��$ q� X�=jVm�	��N3�^9�qA9� �0N3}���~��D���:3%(1�;�q
3���vT��C�)�x;�	��Ah��P�����^�%��R-���������̽�
 (%2��Aj!��j�^����Ut�7H=@9�#b	"�@Muő�P�:� W\g�U���DL���Z�I7�R�C�A!�X�kT�V�Gl n�@�7$��y����Ё� �<�V�ꃎw�U�9�nԍ��)x%HE$5���~���ΐq� s|k�Y�D�Z����Lj��w�LZ�����zqx<�1+T��mu،�����y���X��ɓs��x{ށ�}Ĳ�j��ce"�)���3usi[o2����E�\]���Ms]uX�0́R!6�Ύ��Z�g�����bܢaY�R�\��"�7�^��\�Y���CP���9���P���*�����U���1�- �*	":�"�\qp��
�|tJ�9�; �x��8 8!�I�5�@�u�ul j�1��"��B^"Hq�!�u��;�PI��%[*f6���C�;�{��dKE3����-�ct�]M�o��U�^�h%])k��뿿i��$����s��Z	"$�6Dָ�6랴�PC���H'o	U@ �@Y��#�/w���E:����y]Q�Y]V��S	������Hj��"LfȖ��t�|K멄� �]��U��+��4���)����&b��H7K�	mk��V��n��p�X�M�&��%���L�ͮ�}R�8:�`uA���H�aPI]c�o\�MA%^�Z) <n��Ex�I�?]��a�hAM+�͝�w�UV�j��	5H�	��&�VGZ�Z�o֥b�@�^b�����D�)KEMA
�jל�5�@��ԕ�	�6��$"��g�����:Qk��W��v�N�̪�*C��؈8T�P�/#"p:	�3���\�a�g|�k~`C�4��tor%���:3��>�&}(֖3�iW��@��w͆���G��ǋp(dYi�t#N�N��
�A�t�z��=�ڇb�ޘ��W�ɬ�eŞ��^ăǝ���8��
���{i�9�&�>�uV��e�7+CQ̀?ݹ�P���}e'8�W���#��v3mc�k򼙇���v��q��F߮'� �1J��$1?�	#�9EE��%��Qj	!�#���=3�VZ�rE��9T��ҡZ-֞E� �]�[�$��*�s��$�\��̌��"#6Ge�h���IF�Rq ��'D��$»��$���2�!Ge@L�t�h��������J�)�Z�����/5B������K�[�5���[9�*�@� � �����m͸R�No@�fTW\R\���y�1�{�:͗j�Bm��6����;''�-Ah+�DIά%����\`�!�[�
�窫esJ�A*�E���x M��҅��佃��1��U�dLŨu��HA9�mβ q@(�H���q��Y��A��&�VS1�j"_�h$�ix�󝩝T��-��흆$^D���u�Z���q��&��Wa�v"��^��rVT���-$�Ё�@3����=����/�P�.B�	-{�J��V��}IV�p:�H��i <��G����B>�d�':������l>��v��\�;�N/�yi�_E�P��'t����d9��Y�
�vlY�V�E*�wD���ֵ�=��]l�(En�y�<<���	�%PZvk�X�t�A,u� �B���$Y�J�i��bQ�m6a���l��lD�`�6�oSXq�b\�lq�ut�l��nN�w�}dQ���M�S�wi~EO����f�|w�c�~��(��|N�x�^�~�&r3�q7q�; 9����L�=x����Kf��1������;�_!��]4
�N��QlԼ������kr��m���x�8TH��Jw^�A����Q̓r>J\c/i��*�]���8�$��� ���a�볊56���񞷓��ӈ�Z����C�#�(Tu�q�;�Y�
�\j�]�r�<r��#b0#ٱ�$����f��b�� ���C	�2�N�����+6/�^���+��������[�Kf�4Z��Ѫۚ�7��'���{ِ0ۜK��*��]a�X���4�ǧ�2lna�9�
�ݲ,	"dj0�Q��A�V�,�p�!�	���N��~�| ���S��g��ԙ��뮆Dnɍ���� $��>*8i�+f�@���4��ǃ>3�a��?���'ۍS���=���0��͹�b@�5wP)m{ch��9i�2�~�ep!|9T��5� �;c��]w����Y�4C�v�M��ז�h��.֓V�hY�+GE�ֻFh��k�*	U���rK^e�d*���Hˡl�4J���Dڙ���j(P�۝Ĩ�Q�^������Qu���BEQ��]�=5�:1L�I���u��aӌ;G.������yi��%fJZ�B�
lD�P"7
^�����UP�˪QQ���e�SʫC���s�N����t���� #'�Gr�c뢣(A�ҳiA�9��ӳ|�F�v�_z�o�*b}��}Y����x��篌�iH-(ʴm^��ω����t͑'�N���Բצ9�3�r�d���)y�W�FgP\x\Pͱ���mT�ġ����ߘ�~*�l��&Ϸ�X����G���?Ɯ��}���ξ��A�1j���R��G�>ݳ+J��ӊ�&�Aۄj����XC��5'Wt���M[A�����H�q5��S˺�ءGr�[
u�
��Q���	��u�1�y�������TEZ�"�PT@.�8P�(kr�jtxI�u7jl�a��O,|]�!�O����3�+�ɖ'�*�U�u��ot�����?���8:�(Y�&�!�� ǽ�����&v6�� �> <십8=qn��g��ۏռY;un���ndnBJ]0�z��2��Co=����h�	�/3��4W����b���2X�r��sb����+��M����C�~�w�9�Bj��ܽ���G��(���P�ɕ� d����{� ���N���ټ֊σ��)q{X���al&:���{��+��e���w7�o�"�E\=���8�F��a
�e��4���S�t&�wy6����B=@��!E	%EQ�$��*���NiV×ꯍ*�r9C�
�L��Y�(�+B�(fDh���$����gIZ�B�����J-hQ%�v��K#�*������:����q,�~<�T�:٩�D��M���MX�RZf�f���0�S2l�9+̸[��Yn���[M�CFu��������� �%��c1b�rR\ZEL�ZL�*]p�:f�W��]x�l���M#���nZ@td��a���vŏ؃�W��՚;-��*Xv�\	SB�0�R�-�Qꔴ�����3[�hӳ��k���H�R��x��/���g6t2Ӕ���p�]v��Vh��l�*WLbhc�Qo2��|^�rx���NS�n�Ǐ�dњL���H�e�.6�V�Z$c؍���nH��0��9�2hPNlY)5آU�ePͩ.��ʪ�iF̉���e��çwJz�Xƾ��	�v�:k3b>O��m�ł�sM�v�6�ȐE�(�GM���v���R�(�-�Z���%DP*���7h�W\��������<�N�꽲Xi:��᪂8��
}:���1��Տ��U�Q��|� �ӞN�g�;M-W�'�K�+0��33�'Ώa��͉�m�-t�Sϟ:���z]��-����yӚ;>��h�)���=�(�`�،�Ybn� Q�\}@��Ӛz��Rd�ԋ��j~�<1V/걌"��tݠ��	bDa}]�,�Ѻ|��>w.hٙm�SQ�:&׮���K�/��rU���=���J>���.�C;w^]{���6��MD"�}�]lMWu�B��D�.������i=g_ֺ����gէ��87.1ԫ3��_7G~>��<ָq��@��Lhm��5���C��M�۠��+�	K�5�C�v�@�hg)��(;Ci
�`�Dݚ���:��·9��r�b�?_}v�7�DR���15��5h��T}�w���К%��cPK�I�z�B&<�A���{��|��Y�*��!��x���
cõxa�qf�n��`�+b�.*��YJ��{�Hq݁Q��I� �}zװ��n#x)���(�u�k�n�"�![��˷�x�A���9ɳ�Fť�櫨SVj�n�F�⃠�-�#m�3Z�:�8ؙFG1CmZ�v��c�Bh�PElѭ D'J��~�y�)!$
��v�`v�U�Ov�uz�Y��^
�\H&��=��� �w�N��?��v5���)�5�v�۞�c�x��)���Z����u�>wgX���
Z��Y�gs����`�9�y�չ�TV^��Okp��g�d.̃D쏤���hӳ��+��	c�,Sˋޫ���=�E��ڤ>�f[�J':�r��L��d�-@�j���J�tj��"wR��I��0����#2��r)\��K�.�O�`���ө�f칍�x�=��nv�������g���_�1���Q��X��t�&�zO�VVQk�L���<�����|������,ĦQ�\IN��~XcΌY�uiN�F�]�˶�Qq�[��ݵ�C^�7�Y���x�7�j���s�-����n��xxT���R1/O�DA�G>~�Oi��J��RL���U�>�����B���*��f��{�#�J�p$Lqe?(IB��B��Q�<�g#�v7����p<.}�뤡�ۅ~�N,r}�}��������rz8�J�5Ou��l�ܩ����ߏ�7��V2��̴�u�1�D����Dc�q�fd�	Bݝ]%�Q�V:ddlٿz�z��e�m"Rf��#��U��[������'���<��E��̱ٟcܕ�&�T�p�CWM���5s�]���j0Z1!^�U�\��uF�zS��c/T"�c׹�L���ƠUقo>}����+S�b���u���Q��n:0Oa�m��O/!���8��W�� 9�T��xe��c�h����LLb_ATf����PO�^��^t}���!3Ǚ�fvF�0��佃y�B�. ���AI_���d�r���S� c�\�7�@�V�3�Q�U�4�МBml�ѧ���������|�:!��䰺z�����`���u�[=}|�y����������Ok�T����Ǽ,���]_����3�ª�/Ij��Fd4���ȉB��k�8#+*p57.�k�%\�&wΫ{}�s��;}���g�,��q��$��qu����#6�2���h��+�S�f�`�_o&��qĻ9�	��!�}�ݡ�$�ND:6ɆF�Lp��qd�be�{��xX��^�]��&ў/ݍ�<��wD��F&�	Y�;��*��P�w7[|�L���&N����S��$����H��Mc�{�V �r;�zQ�r���;����,�t�d��q�^��.|{�W=L�r���r��:��p�EʠI(�@?���O��uP�,p��y�B�8��-~��RCh��eU)���#�8I���@�S���p�`�l�dL��^[��<�4ɭ9.8��b�fNF�n��}��Z�kx�	"gt��q�5[�3�b�l�[�∁ww�ﲬh�&1w����0�ԃ��	�\$[dD�ռ9=g�{)Uy6���Y��ּ�FR��^a��)�d�͊�2S")(�ݚz�/�EA�!8��x�����"�B�H��rɜ���4p<���pI���p�����bX�����U�M���H�����k������!7�Y�..�����g��_Ŋ�Bj@�h�2���8��L� D2�!_�8/��j�����x�<|<�z���zbґ_e����� E�v�d�Nq�yH�V���Ħ��r5!$C����f�G��S�'ߟh�h�m-�5�m5`�>z��>�7T�n��n�'F�#�8��5�Y2�"e�7�\Jگ�(�V�|8��5fC] Г�l���Ha�F��;rL�}bS*YA���=miyy?^�}��{Pn��S:ƨ-�w�7���H�F�TVF�\�ӇW�۹���<��x8)3�������=���̪*^Sj����U=������8��5f��N.e��V1G�1��&��_g�ww~{�=�t39�;R.����w��U��4ka���e'��w.'݊ﻑx����9�NzL�2tZ'�7/��bjr�ڣ8�l�ci9���0�¯�&p��}��7E�{�|�}6��Rdjc/]Q�.o���u5r��P�᫳(E%]\S�Q+�q؎c�˸����1�G71�΃ۜ����̞8��z���ݗds@�f�:�P0�1�k��|b�!�ܐr��)Y
����ހ���QfM35���v%bg�v�QI����3�W�YeTt
@ZB�� ζ$��»	6B;����@�vmD�Ub����V�p ��p��I�f�޶�R[�'���;{_�/�c�>�$f�틎C�ש�"��'��NP�B���t��c(N ��6��!��K0�A@��BI�Nn!��;4�2#�Kx����9à��i��R~>\�Gތܶ�d}�����6��|1վ�^+5�};�N9���u�N	9��'�p�d"U���	�y�q{Ϋ���iB�	�� 8J�.|i	�;t�FfN]H�͋��m]{�*�wl]��M{hq��iL�]nӎ��Ek��_s;ޮ/��>�����SW��?���ދ�Mvމ����;ԝ�#�3�]r����u����ޒ2����dLu��O!���/%9�t�d���1�N�9Sf�
]���ᖅWH���&��<zE�S�q��/F�,��E������}ĕ0�Ք$��+,[E�(�w4��)�TCHD2�"����B�I�#$8Z��&߅��-7�R~�	��V�UTuP�U�������̸U�ﲴ���=�#���3h��Q;�t����y�҅�]]y寰�&�	O��A˸WN����q7����0p56�\�9R��[L˥���3���0C8��D,>�sc���W�mQw�Ĺw�>�d�$�2���C�[�ys��=�Ϭ2ab#9����k����җ��n�Oi�t"JS�<��u��w{��̹��Ut�<�N�n�X��	����/}�;�e��ξn�&�z.�C�f� �q�<8�#�����N��3��r��=�d\!]�S~{[�bb`��~�1E��C6y'����D��$�a�63�٩W.��(����rWv�4���̪��w��%�L�Nu��;��BЫں��W���+S�%Jn����w�*�D8I�G���eR+-s��֛��U8��9�*�r;U�ܪ��.�|��i�J�a�4�5J췭����ձA-Y��s�����w+�-M\0�e�R�f��wmn�� :V]u��F�H���.�e�V�A�-�6�K�UtB�6���齞e�Hxyy��'��GA:h�(�\�ZA偋K2ۊ��9e Ã�
�\=L�B��'��ĭ�Ԗ�n����ue�D��P�К��7YN����[؎�c, �]�qa[fs��,��{a��[�ΰ�R]�q�X��b�Z����X�m���7P�%5.(�AĬ�8�tq���mn�\�&�W0�6mn��r���R�˭�G��Mn�GiR���i�s�U���iV�ͦa����4f�Ǌ3H�*��˓T�B[3����j�L0,HІ6ZK)i�cR4��&֜�k��Q��kʹ���ڙ��J6<A��.�����}�Wf��}�ż�.�bOo.U@�
"uCf�
O��/�~�7��?�+	��$�'��Խr���L-�
�������_�����Z�SMf[f�6���|��֖����@_���b5�DG2���9�]B���q}Zn����'#H���9�l����N(U��-�{.ҷ"�q����9�^�WL�a4f�MDe�B��iy��C���?���d��!������	A�{꾅\�}Y���n�;���LW<!f6~��@V�ҝ`��
��S�
�q�M��B��"eu��u�jb pa74`(y٩k�Jm,&��QrC���dy>Y��w���Zk�ͯi��^8�զӫ	D��8�;�<��8�~e/�f�.݊��%�;� ���|S��S5 A��,�q��F���ય�����]]�7ޝ+^���ET�9]X���Ʌx����s��k�M�c��#�״�sY��]�	L���3���ۖ�FȚvq��ʀ[���OJ:w���{'��}��5�JM�싴n�6��Gl��[K� mi���f��	-]-���,ij��5��Bcha��F�5��2�U�L��V�ډ)�w��S�� ������k���#ܘ/0P�q/Y|�zex�G:�4#��������H�LNctP��:��qY'u2A'-�$��5��ms`��X�;�0H�lE�E�V�~����TţjhZ��C߿_>D�p*����6Q��{�w-��u=�9��^v��:�0U��K���u���Ngj�����
�_��Dp|s$+�`�u!��(�nF^�@�&A8Wն:��K�j	:}v����0H��J
Q$Ű��\H֬�$�1AU:`�Q!�c2��&x`����~O2��l��Dv&���(�(���B��õ$�يu��q-���i���/g	�1��V���12ۉ�'>  y��@��˜!����"�2�D��L��}u���j^�X{]�2����x���-~}�LfT�rۈ��'�wpZ�<DZ��l�
�0������'PÀ�ZP$�ݠ�TA���*�$��1��Q�m�Ӝ���|������߽���<�o�i����ʄ,G���ԃyc�,�B���9�x�Ql0E%$dK
�B)��00�8K+��b���⊛�sQO�E��e�"˹F1z)I�����%9�/�uY$�H5zI���q �pJ�r�t���
��a9�7�֓�<�"y�-P��XDX��ŉ�u��P	A�V��w��m��
�+h�[r
(���mVS[KrY��iB���kR@��44b�^a����"���1�.�������&��[�UU�מN���pKz�2Z���!�0,�U�8�Z�uI>$x�|$���`g�+9����D�#��=��Z䛖	'HG503���C��?Q��xJ�I�
�s��R��wS*B�5j	(0�e	A�\D^�rOx�D���9�Kb�A�� *�BY�l3"�f��=��Κ�B�#U!�v��1���ˬ#��l���=m���΁����~�B	�a�eIon7<#�2����N�#�y�Z�L�v���Ooe�`��E�p�y���ɳ���S��$�{!G12sGH�sռ�"ϗL���n�$(�(� ~¹�o'���Q�����M�եw�PC�֯{x?�ͨ�qCpa'��x�)ڪv0���R�BU�جE�y�SNc��'D�35� �U��HN-����b{׃L�������p*_�w�_n^oӗ��~��x^�^�����G�#�xq�͵l��b�3��d��T�~Σ8n{�S�Z��4>V�&��(���ɶ��u+(p;�b�f��v�$��3Jڻ��hY3�[��u������lӻ陀E�		ż�,��RV�[eN4#lKK��P�ET2�Ԫurĕ�p��䜵�*���u��z��Jr�93���D�Er�8P<��r7pC��3	�gM�Hs�YUsD���\M��|���B
.�U�'ǡ��ߓ���o,r·�{9z��mͦ.�	�E��J�U7`�d�g�3b�i0Kn�1D&��Z�5����V�$aD�|�Ӄ��;�0S�	G�/C�iv�i�
��<{�0�suG���d�J���	j�*z��m+��DN ��{u���J�o]��;�WQ�e��z֐��mU��A�d���i�#T����/u��H��Pb�vO}μ<�}�������l�o�O/C6��/Pf�?bm���Q�V�'%3�Uo'шQ9�7�ړ�:�r��jg5I÷��}���Y�m�D�FK�^b�y԰(������;Z̵v�e�z�۴���z=˾:�7�A#7j �]�b�cY� �a�6+��mu��@�Zk��ۢ�j�֗NXJ�J��l�M�u����-f�֤��Z.2A�̨���!P�w׼V�0MbL�?�����G�C%�N�7�� =������,�=DؚZ���z��	�l�S�	@�o��U�^ $��*M��h7�G��:P"�Y���A��þ����_~l�-Li�r���`�e  �iq����L0Ȅ��p}��o����pf���v��K�L-��b"�J4��ɝ�RI �Ax���0�3	���HD��2�	"ϕ����'T���HgӪ	�l��(��Q�(��d��ͪ�QĈ�̿>3�}�����nL֛9� s.ƍ��NFr�k~�A�Y�ڒ�Gg��;@���I�Wpb����"� w]vw30���+V6�X[f�C&'|��h���4{�9���;��e��n��
Ԟ��xI�~$�3v������Cp���6Ɉ!2@i��:��G�s��d�l�`*k�S�����B��oW�UI��;�L����U���6$�D��ك5\}���:���@��S�gA �@Q��D�,��8:l��ھ��o���Nb�+bp-0��ܩ�p2U�ļr�)>�����߿0V�e�,˒�E]���.$�#|�V��[�!���{2R�t�H�nײ^fV�x�u@H\�'S��DU(L�ͤ����� �0����^�N:�ؐuzu0�@��+�(UEE��w���9�:��uk����2n�f����/5k�٣aė��{Mp��1�a-�e�GV�;�4��lLu��l�i�Pcn���Y��к8�J�Z�Ks�X' �CW�qj@����C��!�)��N�D�T�O�-�H0UY�Iu���%Dd�#NjQdd/f �t�s�fdT�j`���$���G)2V`�,�@Ar���3H
9q�'nX�fd6��@�����K��/�{�#�4&�!&m
4-B@� ^!ܢ�-�����٣,�	�/_�k����]	�� S�'h��(���ֽ7M�I6�n�5J���HP�>6�5K��� ��N�X^�n�y���}���y�����5u]������9��5�K���Mbf@t�;pDfw�8�ͱ'�!�	$�D^/n��CD,�))H�~`��NW\5�k9�1�{p+�T"�A��Y=��$�Kǭ�ݒ�M�q8EA#H^9+�1��Ep�U����7(^� A�b�A�o�B��� �c#Jm��6w����=�w��L���d_O��R�H�s��#��h�9)�v�D/T���z&����y����G��#u2-B@�W��U+$�TL�;�T�oC���~*��m�G�B�Oz�������OH��7���}��^!�'u��S���}.��z��13�E�j�sYP8m�v�CT�!@�&^�NF�2��^r��ϡ���p�m/Y����Rݿl�i�W�ă�9J$��d��r��.ʡ���� L�v[�8�+lL�+�"y��W�i��;7��C޾=�;�Oa�'��HK�h�m�<��A���oq���=7��S��!��Ӹ�W���wh���͡�����Fj�f�N囑ih�*nl�&��Ϋ=�H[����ܛ�&i�	0��o�v���� ^;��ޕt�$�h�����?��M�İ�u��{���w���^,�.8�:��� MD����8���a���u���&jKӵ�VlEm���m��>Q �A�$H'��(�&\u*�OVNC�$�
v9��E��ӧ����/PBwH�(++�r8QC���e��A��ҏZDTZ�
�{�����wG�&Iv�L��L�s�#���l�D�z�!�.<2���&G)!	�I2��t������{�GR�\K6��a�.l].Cfc"�V�����T�f�2y6��5�]J��e�֐J$!Fj�&*��7VS:�cM��J�و�B7�&tT0��Y]xh��,5[b����s&5`ɖf�dְ��
-,��ٴ�����[�ke�Xb�c	m�rg^��@����lCѹ.����VǁڅG`��+HL��k����3]KZ��ԯV٬R͉���i�!�X�K	r��!�kJ��m�ΗaL� U�)j�%ĳʖX�!m���Xh������Ax���`��)Mn�NhQ���.2�
2�����*�3VW*h��m�)��P.�k�
�h�8�i��ZDY�k�����2��f��Aն��e�i0�F��Sdn�!tq2"�M.(8�[n��Be���N�ow���F*���k���e@��z�B�0|��3��ЇY�󡶁5�֜`�ϠM0fx�f�ɢ2	�!A ݫ�o1�� }����}��|q�q�|�=ᳮ���u��t�V��R�+���D.�<�.	=)�ԙ�q+�V`x$�1U�p9����y%X�OK���+L�CCg#�Gd�^��LNR̋gݫ�K�8�T�p��N�ȝL�׷"H�^�R
��y���C��܃$��G����&Y������*n�	&%��{}�36��:8&qL��CcA��$e��%MC��$� �Y�I(m`f�od�>ؿ\
��VS��u���*��s��N+\���[���N=F��$�� �sˁ&���e[�Mb�&�$�Yt�0�֎N��f5�$��Ϭ�n�Z4��lC�&�6�n��������-�<�Ȯ�SYWK��]�����6��4�L��d+�]l━>�TH.�y�$�^�L����=z%�Q&HE���nl��jȀ������Y>�E���W�	Eض\	�~�C�����`�tnr�P�#
A�

IB�b��'#�.�ɼZ�F�>;��&�l0T�%n߮Ԓ	�Y2�ɫ���^�^�|b�ofj��K���)eur�G�{���ݦs�U�+P��F�=�Z󥄒��K!3׸���D�HƜ�{��i����f�Q)r@�	�-'�f�R���W^ƹ�:�U�-/][ٙL���ݥ��\X��)�ֺ0a
�DQr�j��k�YV�w���T4�$]&IZJҒ�l��✍6
�=Rz�>#y0AW����\m����D�:�A@��t^�$����p�Y�E�F�d���d��-��,AҴ��N��hcqX>�� �m�>=x�\͖�"�r��ϳ��yX��J�-��B���e@�m�q�U����z&��J�:Ƨd-�8˘�o^��8�l�H=�2B�U!e���q Lj��8�b� �^�A�7D�3m��E�0�A1��u�<���������Ejen��(��� �&e��0V44��c	��v<��<�EJ��l��b�v���;xO8��8��I7��4�$�,�L��T	d��Ϧ�f8"�Ll���Ɇ¢6�X]l�o<{:�L���z���3��e��Aj�3�L3V�WU�Ш֠ɽl�t�ۍ�xܡAj!%����(
����hq�L�I�.���^x����)h�a�0�&}��M(7�'Y�X}�۠A�~f��2�����^�Ѓ$(wR�y��I����.�4e��)�w6K�-\\OjNFgi��/�PE���5;�-" ��#�ڨ|��ݿ���%��̊ށ1,21wv����s>����	ܰ�V� 
��x��AĽx���:̝Q�Q��!��>�ANJ*���)sJ ĶwD�q�����y�F�	'��[o��y�[�OX�d��ba�(�K�5�^��b�f�n�9�E+��`��L�����o+5�e��mI�h��7d)M�	6@&��6�q�����<ȑ���$���]�I�}5�+���hs~�2��^�L��?:w>F��1�"�FT�]b	�a�z�Ҳ��|E�&�S"���~�B�xN�G�	�^#a��00���f�q	�C����c�z���G:�z��+h]�E�
�u'6$K��3�N"{�۬�軚nU+��ġƵG%������xg��I&
��6�o�h$�S�a������Fr�x�f<��D���ҥ�e#��a��w٪=��w���q!�ٳ�А�1�s:iq$a��aY�b-��$<�� �l��Μ3�a}������C��N���/}���k��}�yN�y�&���e�n�=�n(�'���.�[C��b>S��P���������f�v��M`�{�e��f ;����;��3_���M�m�ms��pէ'3�����zq�e-��/@���N�g?K=�o��N����s�ǗT����%��>���Ҟ�/JG�]��#�̕�2����yH�9�	�[.����i[�wPba;{ǃ��{c���<��ҩ|kݩu�^�������m��3����rz�xH|����4T��S�"��7_�}V�|�>N�4�Ǟ8C��9 =��Y�8	����	�\XW�0�rI��'=%�I
�}J����Z��7��
%����e'�=w���I�Gi0""c�ܳ[*��EH�QY��)�-
��p��~p}�S���)�&�� ��(�r�T��T	������X�AI��{٠��;m�oݷ7=H��e�SC1��c��"Ds~�L�"	�cz�k2uaiQ���'qy��躥YU<�� �A�����h0H�a��������I�oӈ���u;qwL�f�EjY���u�D!��˩�a����Fzb	�~y,20�En�9��M��7@�6��)��w�O;�o$X�z�p�S�l��-JrRC{�/x��рA�0 \���1�x�Rˍ�H�~f�.�J�r�۱Gi3�(��x��%X'u��/�sG$���S�6}9�O;ְ�����)���+r(fL�ٙҫ[b�o<ծ��v�ɥyc����[�,nԩ.�z�+6��u� ��
�X���e��˜XM4��iv��m[:�*)j��b�t�ց����]wom���e Mrf��|�BA���XK(tXdˢ֯I��f���J��8Dj`���K��#�@� �zN�KU��`?����3X���%L�*��3��}�2}���wP���ChAE%(��e�$�a�O0Nj��d����Gfu���x��}u3�U�*����W����j�3�ڙɑy�uK4'{��TrS$�&I��	�~�R	�S���+�ɐ�c~�L�n�z�q����Š�u%		�l��Ͻ���n�w]�E*;%�]���`�nr*<g��t�$YGM���c�$��o��~5M�� -ws%Ԏ�%^02@��>����}���.6�I���|b%��j\FϺ%�	��VXZ�l��L�����x�=����CtQ�b�@�	$�@�� 8�̜!0�D
�C��Ý;C�:B'���l�N�
{h�V����@\$I7l0DU8��Г�8�$�6I3�2gy2H������Y�lfM@@�����VR���P'�(�ڦķ#m���v�:�ˑȭ�vω5��n��CH�g �6��=���	����P�@��s���>r��O�N�@�����P�l�g������y�$"TN$�IX�9I�I&���H�~�Alg�����������'1�v8C5��	��͙f��b�I8E*�����Tٶ��]:E���ß'��8� LCSZ�L��Yu����3����ġ��K�Yt�gkl����+FSc�k��hۛFh*)��x:4˶e
���V�>���S^�_Gw�N���u�M�ҥ�L���
�6}iL�MA=��Ө�d�A��&L�ؒn_���I@�U���A'�c����0淂N��m*2`��l�e/6�<�7�3.rt@qv�מN�m�|XȒ�"���� $��np�!û]J^��ߚ�^����Kz��{�WO3��ekPf��\���Mb�#C�$d�$��"rؾ�\Ʈ��g��c��ya�ȣ)�u%;A��;�X�5z1z3'���P�HA�Z�\���'��/e7��;|'F�Dp�7y���<����?�0�W�#k)suG�z� UE�G���<l��n��^�[R������0g��z��䭍�V�$m&H${�gĜ��p4꧛�u.�!8'��u���3���ߋ��`�e�!i���RQ��'i2H"�7�NbrPU=�'6x���
вw�>��ɻ����!�H�	�/(@5k��]9k���R��0�5s��]J��յ6��?w���_�"�.���E��p��&H�m��#1��!�"�TE�6�f!1��sz�Υ��{<��^ό��e�M��Q�E%���0�1'x�^�av��q�R�sy\A0}����a�H�(Y��.��3;s~Ӿ��V�j��G��+lq�D�H'��~'�yP|����I$�I�J�A I(��U O���D ��}!&_�TƮS\Wm_3��\��c%���`����QmQ��B�v	��������0��4��ڄ@>��ӈ���X��3���m=r�*�c��䱵��ӏ���5֛�Rh8�
Y���&1�~6� 	�ӟ��o���~ 88 '�9D@�A䌉Kc�u�������_�~	��G��m���=�Os�@�z�*  �� ���g�댐z���hl	�Sb_kF���0�i���Ak�/p��[(G�'����ɩ�u�nXf�� ����  �x����]�>V�	c�z���5�JDK��/$�oE��uq�o�郀�0���s�� 	���^F}�����/������Ӥ�w~:�;���K��y�Ə���Zq�s�h���( &=�<�,��'v}I����o��K���͟
��������g��}D�O����m��n�{����x;�r� '���#5���������ӇV$?�(�)�#��E@�,�T@>���K��=�T���D���tp`(��2~��d2y�$�`��f����N!/����甙�J�$>���R�g4|6�T�����A�K��m�{<�i�ؾ)� 	/�=`~ly�o�(�C����ρ�������X���צ~G�,OԾ��o���O�C�;�ߗ�c�����(�y�{���x ��J���}�4��Q ��`3�f���C~���\��;> �����g	��d���ܰB���^��8��������?_����?Q�;�<w{�(�z�'��߬8��In��\�h�À�m�� r���G�zs^:0����w�  '�`�1�z���W��<yz{�=#�z�� d/�!��P����DC[�g�k`�w�@C�(_o]������w$S�	��f�