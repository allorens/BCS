BZh91AY&SY�%S��߀`q���"� ����b>�      �辚��I% ��ŴH�kJ)USA���$CfY�

X�U%T٠ ����J�����
"���(KYZ�֭`�z�Xe �k6�*�ŭKkdY�-1f��im���#X�B��*��Th5�2�Zɣm����L�Z��5YMIհٵlk%��/4�F��m��vT��m���8�S[6��������2U�l����m�6�mm5�a!,U4�kJIl�B�f�4�M�X��E��l��M7���c2X�m�l  .���QTnî���;�1�5T��[Z�MhV���e�) �P���֫�U�t�����:5ҕZ٥m*�ͺmm�Cl%V��*ҵi�  n�}= ]�w)!�h�:�p�U�{n�
h;^�yJ(P���Щ퇹㇠���yZ  �����*��֍S�}KT�df�6-��kTж�� q;� iӾ�Uw� 4���t ��e�����43�� ����΀z�Gz�}�>���wM��=���W���&�@S㓍@eUZ5k+l�m��%�  ,�� ����O�Pyϼy@�;x{���
3�8 � ��pև@z]z���=���� R�z�s� ]�Mޚ=��F*h�V���3$�[>   ܏�C��o ���{�5{�{��z�.�`M���A��x�G����Oz�o{�=hlo<�ʨ:^^��Ʀ���i��k,�  v�  }�ou��: ׽R��t ���  =V�˴@=�۝z��v�i��^��)�եt��r�E):� ��е�Z5jֆ�ٮ5Q�lƭ��� nϭ� F<�:t(e��Ưn�q� �^׺)����=� � Ʈ��.y�� W��h 'J�YZVض�ֆJKSi
�  ���t� ����tovW �N� �s�� h6+�@(	�� ��L�Z�s�Fθ( #�M��54m2�Z�5Cm�ճ� r^ z��w�S  pϸ �*� x8@n��OG���0P(3�;� �stw@
ѝ�PKM�
U�5�-�5��g� �,Рup �
t�4 >�{�8( c��4Q�s�  ;�s�րm&4      �   S eJU`  �`���%Abha �2�JU(�4�� O	�ITPM     �15JF�P��A� F��3R�'��&��=ҁ�MC�S4��Ϡ?��D��S>���\��=�Y�Z�u�6{�N�|~w������w7����UEw�E p��
��D U���������	�3�� ����S�QX?��U�@*����T�)QP���o��k���fC0��̄��L��29�̦e3)�	�2��̎e3)��f0L���&d3)�L�fC2����&a3	�L�fS0���&`3!�L�fC0��̦a3	�I�g2���&a3	�L�f3�f09��&e3!�L�f&a3�L�f2�̦e�3�L�f2��&e3	�3$�f0��̦e3�L�f&29��`s#��L9�̆a3��fC2�̆băa3!�L�fC2��a39�fC0��e3.d3!��f�2��`3!��f2�̦`&Lș�0���#�Ps*`�(9�G0�*�aĘ9�G2��P�#�s�d� ̢9�2��ʃ�@s �d�(9�0�0�ʃ�Ps"`Q̢9�0�U&Ts*a�(9�G0��Qȃ�s�e��0����s"e� 9�0��Q�eFe���G2��D\ʫ�s*�dG02(�P\��s.aE���2�fA&�#�s(�s
�dQ̈��s ���Ts(�d̨��W0*�P\�eQ�Qs�d 3".`ÈaP3
��D\��Ts�a3
����d3)��fC2��&`3!�s!��fC2��d3!�L�f1�fC2�̆d3)�L�fS2�10��́���S0��̹��̆d3	���fC0��̦s��L�f09�̦e3)�03	�L�f0��̦d3	���fC2��̆a3!�L�f4�fS0���@�8�y�˰G�?o����ǆ�F{��M�Q�1^&��ZB�s4܆��Aƀ�P��Ytӑ,�w�!ñl��f�n��$�2�!���˱��%�մT�4�̼�U(���`�P@�M"�P��{���fӛB1��%Z�ۀ���l�֘�#r�20uZm��WF&���P&62˂*%C45 ի6�^L�x��n֪7�	8��Z��aX�|��Kch$"o�Z���`Y)i��va�Yh�6��KS�EQ�����&�j�����f�A:��ceэ�T��d�bS�����g��oNܻ���7m9��N*u�ADcH���ǀtv�g��@�EC!�{	�Bۼ�.�S�z��*�9���n�[�j����VC�l�Z�f��qY�dk�%�*B����-b�sL̦)UдkX5�e
s!�S��F�8�7sFm�'X�B�R�*,�!�o]2��-�#j�n��O|k3���t· ����t02`���fB�UsgT�[ �D����3D�[H���©�	�MҸ���+.��4��2M��Q�--�Je͠�ٚ^(#���dg���a8���٧pS���4m�V���� /rB�թXY��.�,����u����ko(�Thj��ڈ<�%�3Dflŀ���(�@b�IV �����r�j6ٍ��ca�͛�(n�]9N��9c�ۑ�	�N�&��0i�S%��H��b�1Q�ixP��h�t����09��.�f�="T:lQ��Tm��6-�)X������T�ͱ*+d4���R�n�y�3��q�R�+Y��uyS℗����թ�E=פjI�86����7��Y"ڷ���-�N�[z�ղ�)T*ap��Y�d���L�u�-DP�ݩB��4��-�
F��r8�0U���H��!q�L�؅m<�nBd�9`; X��Y�7*=��vݺ�ȥW4
��Z6������L(+�Y܉���Zh�m��V�6��a�,���[yk(l��`��*rnLe�G�rU��f�EM��p�n1�ƌӣtՀ|��
�kM�lNi������4�Z�㈈�7j2n�و�[�]6qk/h	�e��M+(I�#����5m	�[�֨�T�d2[�D���3����P41�R��W�d��� �ַJU��kB�jU#�,e圡�5�jD^]���L��e�JkՂ����XYt��VZwD�_=k����hsD�֦��U��ت)i���t������:���nB��sk1���.,0�T#U"y�9��ڽh�v�ct�ebʽck��e�7��������Y��L{`X�V+`b*���ۚ��سE;�ojm=ɦZ�̬�L˰���1B�����Xd����
#M`��;�����Ě���F'({2�v���n��
d��U�s"M�PRD���Y��F��m ws�s �4b�Z�L�i��� l���Le]+�j�',Ƣ 0�Q�=4���5r�QV�� n�5=4����tἼ�5��A�n�F޸쉺j�/N��ѭ%v��T��l��N;а�ώk�Nau�J��36չ5l���%]Mn%X�ta$�ڡ�2H�U�eh�'�p��f=�{Y�)S�	̽1�[�r&ۣ�,kx��ҧO��46��S6�h����g��m3��e��J�����m묨����@`N�]�S����װ3�N�(R�r��MFP�ZČ�5YD�VZa�xg��7�K*��p��+�=�+we�QH��x؃���͹�20ӥ��2��F
��UҒ�Of��.n�W����b5H�kw�4
l�u2;(c�$r-�[����Kr��ïAf��9Tc���z4�ŰG+7O�W�Ļ2������SJy#c�Z���^�854Y&�StKHu�@��x�R�KfFthC)ѭ�{�uD�
ViFS��$�f�*޷�������t���x�@bf'�5|��Ysh�p�M���l�{{1U�<����0a7�xt�V9z�)�d���:��n��0�ʟu�u�eY�'�ݖ�%k�aq�A�(%v�8����o4j���GwElY�<��H��̉^`�(k�v�E�bU�D��i�Y�r�	e�J���Wm�����ݰ�'�=�bLk�sG^��oe,cTג��1�q��n�c�t)��%�yt��lk�$�F��y���^�ڏBAt���a屆a'V2t�M.iն�Y��Ը��ŷ8k�n����'�w��ò���j��a��&1���k00����,�N �^�X7BҬyv+F��f�b�)�Y����mfӭ��0YpU�Lt����X���f*lHq��*SW/�� �p'%\ӊiܧ���[��ɍiH%Y����[��#)i��v�� �\���.�����s�.�ݡ&���&PsZpMz��I�6�Pؒ���=�v[Su���E�T�i�[#�I��ci2�H�e[z2!�Y�)�P�4U���8�U;b�4Im�4�V�X�D������.�9�X�ݧy�d�7a���[��.˘6�k)�{Ō��b��XS*"j��س��T���"�i��S1��^#B)�ڑ�(�G1hE�ٴ��E��{p�,�ǱVz��c[�����2ㆳE-S"�s6���A��qE���[�J�NZ��,�730]mH��܍[�gu�ΪVS���V�-]��$�v��ݶ�fh[[V��]��@�Y��ҧ�UQ�cF&����%��1���C�D@([�7�q�[KR�4QޗI^�*e ��^���Vzl�.��2+���`]�+6�h0V�-�����*����k�x:���+��Zh=��]�2Q#S&
a^D�af�dCS���@��ܬ�cCl���Ū�̛�1A�늕b�-��1�bI�HF�T$�Y��@X� ���+w4�eI剢�A4Uh5�E�޽�͍X+b��V��u3���r­+bd�̋
o�@@��b�%�P��y�6Vb�m�8��D��l�2VCN�<R�]���G�EU��鼻��8'}]������ٵJC�Z�1�.������݂�	�������+3oХzl�G���X� ��	o=V��.��ڣܪ�R��"o}@rcvѠ]a*}{����s1Ż�GJ����
gq��tҀ�{3v	�]���1��(P���h�C(OS���+(6� �5���h$kI�:�3Ah�j�eU�C.�=��Aa��G
�-��J;��+�"�1�Wt�n
#�4)�Z�1�q�x�f,�m�*�ĩPz��@��],&�L�N6ɫ�Nṁ�R�`��M�+0ʊH]k�u3�:7&b{C挔�ڑT�#���X,���݇()����z�ix��f�����YnP�2�Q�B��+ZXUA��b����3i��n�hJ���5:�n$ȼuV!�X30�̹���5+�z6�'[LEb���������z���x�A��AÜ�3lX t�n��s���:��z�Y����q��T�u�c�V��a]���X�vX����}R��h"˺˭��&��w.����wz���,�n�I�V5����������G,�*9zL���I��:��� �f�Q��l��v���8�V��1hu29� P�ˑ�H�7y���f��e���7w#y��r93~�O�+c��޽l���ݬ��P�D�^�S��/pJ~�]�-���ƨ
��s�2l����9��?�vb��j�B�l��&�h��A�R����[`�un�^��!l����ayX[Vq�.�eV
 Je���cH�^[լ�uVE�ݰ�� �]Z��qk�r����!�,n�d��@4f��^K�(*�XorȔ�D�u��`DV�z��°�n�J2d�1���O�9'ڝ�gI����۳��VsYб�Z ��i{Vei��S������ۀ�om���W#؛�-=gk4��@p�!��"c[)P�Nbɭ���nFt�9V�Ү3mM&F]�WN���V�-���$�sU��|0ݒ��5ݰ-{�wY���e���ơb����f�!�  �f
��xu��e*Zbu�5�� �cL�v��R�V1��xaV�A0�Sۙ�-Q�{��9F��&�@��@o2���x�%�+q�t�2+m�%,=�[�F�A�LgsQ�?mh~NQul�j�4���+;[Y�S�8옆��¼�F��
�yy
�+&*CRɨxK���nU�W�$�7L�@E��6��Р��r%���K�]l8�1k��M\�ue�M�n w`�.�Ǆ�u�tV��?^�+d���⸱�6�a�J@mm-Kx�V攰�=sk)��a�	�Z�lw���R���[���V����΢�S�!.�u�S`,��u6�!@��P��C/�R��o�"�f�*��� �^�3o�dӀV�.�aޓ#䥸�G]�ݬ;�j��f#�[�;����Kv+w�7uݢ�8�L����^V�mcB�\��ɘ�[/$�{x�e�QN��*�ԙ��0�nfa0Hפ��U�tĐ�u�A�Q�&���Z��f����as
�z�յ���.�,d��A��ͩ�P����!�b����Z�x����&L�Yb,��R4��h.9L㬛���Ei�t%��^�����h#6t+��23e���-a�hba8�к9h��c
���9����W:�[cF�[4�5-5��n���Z�Sf���Gti�ƉO�&ܺ����p��-e�6��A��ͨ�fiq�썹�X+|R�R�m [�-�`
�̱`�4���.�^��z�������pP[��8��@24��zܻ�{(^�١�j#�ŢN��IT�Skr�6�n��f�Lw�b��J��oҞmm��؞���������z�ۛ.�Dlp�Ӗ(7u�qmf�bR�u�y�v�cN3�;7�f=����վ���e%wI-y����s�x̵0��F�6��?ؤB`y+6��ڎ׵��l�ԕfTSB�Xe��X�E-Y��CEy�[�vZGR�Z��|�L���5X[��G5��Z9��:0<�zĵh[x1Q��Uv]�Lcl8��0�D� *���8�9��qBn��fVn�u��IEˢ�#kX��Df@�[����C.^�( uk(8���H$�FY>v��%J{KQ֟�
c+^�*�jT������Jcj'�����HG����o�;ݬ��  X�����9Q b���l�^���呕g1ܡ�8��J"G���'Z�\9���U93�Q��3Z�F���R���N
�TuV<l���f�;�ڷ�>OM�G3B�2ӥ1���u��h�r�]M�Fã@�Y����%�
;��	q2l�^Z��b6��Ш�4����W7DVVҕ)j��*��v�c�����n������)m<��՝�7�LP�m	��G6��O�/��ܥ1��q�̬�F��J�0^]��HƮaZp�ޓs��cM����8�1uJV^b� ���*�Z�ڤ��PY�r�)�QXbŦpa�D�����ӲN_���Л�Cm��R!X�m<��.��
яb��t�\�e�J�z�5���밫�$��-<̴U ���mT�{�FA[cN�.f�7���j�<xv��
�1����R�R߅=n&�*�`!y�&ލ�VR��% �T������emo�%s^ؽWo�J����bԨ-(-�uI`:�dmZ�LSØ�6�۵ZH��2���擺&ֱ�v��P֡چ�{�vV�)�n)W%8^�^�(n�]��e3�gjP�pi-��Z4�S�֗�r�L�����oF�s3^�,R�Pڈ�2X��V�Of:�/j�\ܦ��\{�(�Y�on�B�`����
^�6� ERl��@��M��z�Jbw`݉C�R�Q�6ɤlef����m5:f�"�����i��<�r���h����-���xq01^P��!������n+�X.�l���((��#Ҧ13f�̺{E*�G�*7ov��ӵ��Rɬ<�\#34�s6:H]�
s���-�8�Z�Y5f�k^$3� `�䖴�bmj�[f�YW2HQm;bI�fRg�3UfPYm5rem1@ʈŁ�z�`WA�j�i�['
�6Y�ojRU�Z�8^&��kfah������XzK���b�����)5\CufBR�1�*�#^�1#�k�A�I35��'͌ĆROCE��U.�3&�y#�ɒQ�����4��mE.{V�&��l���;=AV:!0 ]ƕ:SRd��!2�=C��<��|�ݚA��Éе˱�CE'����u���ĳUc���v�ek�6����S&�G�xVg/���e�F6OP4"9��y� ����ƭΈ�b�+�D�\�'hK\�t6��dR�7�Y\)%c`;�	j0ka�G�c�5x6֊�G�3�S�NiH�N����V<��\ƴ52�<�� #t5-i� ���{�}ņ�j�o%4�d�Ga��a�4i/պ�F�91�p��}dP�:��7#��mЋ�N�i��t6/�@�Lyt�<
�݄8�M������Ðtr�CFH��m^i\�W� A�r��]���`<d��#�L�N�o%/a�E��X��2)�XHC��'6�^�KF8�h�����d
E��
�ݣ	/2� �=X�Iw7�<|�����`_R��ῄ�^)����C����Q�>��Ȟ�C���Y=ֻ�� ���.�E�
=V3�42���;[��@6�ppB�r����V֘Z��9hj�f+�áMs�X����ȃ 1�K���8�!|%+>�s�H>���������|�����"u�_���������~������nx�����#�=8�J`_�Ω����
�;��fp}��Kn�!o8�
��Uy9W=��kb�XX��9.��݈�Kx㙔�s�`�9k0�c�6)�Z`3�<��e!Y����s̨���#�P���r�T�~�f����6�5%�ڎYrև¦�Ά�\�N��;��c�%lbb��K����U)u����Ô�M�f�Z,,G*�b��W��o<��-�U�2"��_b��2��D�=l����_2b��6IX�p��fr:�R���fǻ4>�Agk"}�	XY2��Z�b���}vyA��ӷ�]��Y��W8ކk&�m�����;�Zd������]$38���(Md@�하�+Ӎ���n�|\��ծ���:SS7�V����w�����O+\�`-�E͈C����%�y�}�E��mfj;�ݤ�q*���B��ԑU�xo���*.�'��e����y\{����J*��Yx��}�dl�r�k>�eV�3^Iܢ�����}��Z�8��s��
$X�9v�no�V��ǛHU��g���������z�+X9�fpǀore��l�3k��eru�X_A��L�p��3�������90[�C��+(q����PΚ�5{��=z�x�ZΙ��j��T�}��8^u<\���i��hq�@�jۣ��24���ʔk\�������=��U��d�� �_�-�:�]��W��p�^�6�<�S�$���������;t�f�`�C�NB�L��`P���q!��--=B_l�sFVdI]<���v����UqX�D�wy��f�f�V�k�f��tbAX���yI��W�$ǰ�K�)�Hi��z��z���Z.@����E�Ajڏv[:;���xL�9aS�iY�F�*���7p���t��KJ�j*�,bb�R^j�x�<[y�r���r��.i���t$"���s.�bz��}s}~��.� �啫 �v^��bn�O*j�x4g���1a�������R��o�S�����U���PT'V�����e��ȉ�]�:���ޮC���f�Z�Ag4� �
��l�@g��G7>�"&蕂\哥*��B�W\�.���d�z��}m���N������2�ikf�7Aޖ�_�َZQ���m��\� H�ҹv�����⇰cE�fWQX�!َ�@����-L޲���4��a��P'
�|]��V�RO:��ԊI�ǌ��o�m]�M�/��1�~a�i��5Z���XΉ���r�>�1jg?s��P�5qO�<�tj���
��k�1t�77hq==vZ�彬U�l�f���lf3{��h`Oݰ	��y��E�}����4���aZu�^�&�w�xV������pN�K(�����q&����R$b����aN�ŏ�ZW9��^����]�
JN+�e���3\K�����%���]�����t��ޙ�D5մ�i����ֵ���X)��n
���j�Tq���ۭ&��b�α��o�՝5������j�f3X�c�R�/���/���p����e)Vc���t�!CJ�n����,�(�f�5�T���g6��}�>{[ �z����b�嗎�'^ʶ��j�jd�Ÿ,)���9I1L���;��(��u�SX�jQ�8G�:�0�)���O.cB��\�t�1�V��n6�z�Tq'�%u*ڛat\�]�eu�ޛΩt�v�4s5f�ޒ�6ʼ�+o{�!1>�v�u*�����u�q�=u�lIL\b#Z0;����)3�>o���:E���7�_ay���v�����1�,��Z{,�F�t
��[&�I�+/M�4+�.١�caL�˽٭��4S�F�5oo� ��:ׂ]������1�Qź�B)�nN:���>z1ƙ��X�2��X�ˮ�k�F���7f�h����IX]e�����4s"�^^i#��,+�c�+���]��a�ͤbg\d�l���j��؃���6r7(� �܏W)�%�/P{�+�!u	�\�ل'zM%���ST���R`���V���"Hity8-"���uuI���W�kc�:VR��i�pu��tf�f��থC-�Z�z<�f�Q�B8:��`��Q�[�LjU�>/l�������+�=�E��mz�#�*8l2�P�NVH�'ǌ�����w]IF�Axһ��&|�J��m�?LYvA�W���+M�$k����c�m��D�n�B�2�Mrd!�M�nw�s<;PI)����ۘ� )]�|�[c���Jx��y��Ǹ�#���6��f�=�V����6��Kt�*Z���wnU�(X��:s�9J�	ڹm=��.�� ���BՃ��S�l�rv+�� ���������B���W+jU6� ��tu4i�A�!�Ze��e�D�=n�c�Z�^ջ۹٤�o���(����D���1hMl_�%�mn���e�@�vrv�k���P��rPJ��r�s��t/n��U7�i�;Y��F�V6K⽒��>Cԛ��V� �sa>���XŁ&p���A��Do�͒붧`5B	d�q̕Sz9��&ѻ͏^,�y��������ã��9�s*-O-'q���_��^q�%��[i���u/Y|(T\5�� �����Tmľϭ9��^%�K�+�袮1d̮��x�>0���G�uP�6wѼdZ�k;&ocҶ�/ۋy���3���v�#%s��4ORU��H��΂��Ia��AñO5	s�n^�F���� ��ҫ�M�l$@���-��h8�B���m�f��g����cA��%;���nR����lwm^����6�&˸��M������ -��%+��MH��[��l��bf���9<�U�hLV�x
��sP�i��'s��m�B�y��w�-[��Y�ի6��݀&������b m�;N���7��h<z��e���3k��:R�Z�0��I(�&[�cuլ�b"���F�����Җ1c�{��-�]iYQ��r%i�h�4oU����S��ߗ1�Ԝ�`(�NB]eZ��˼=�-[B�`PB����Y]ۙ*�9��b^Ѥ�hx���z�ݻ��.�C�6 w�Z"�/a�ަ����z2�El�%�w\g_=�r;T�R�e3.�l,e���J�����Q��8��噮��)CF*g���}�8���#��}��!Ͳԏ0�������뾦�{�]�]B��5å�X�^�U��֍=�M��}���R��1eK�^�W�����L�'��}�;�$�UgYF����ڱb��v�Pm��҈�D��k�yS��Ȟ��P���N��p��%|�ѸN��]t?�+�����Ȟy/���	(��\��*ɳ������������Le�&�<Z�㭝�8h}8�#v��x�cy��*����m�"
7�k�,��@93V;R�=�[ڈ8�H̦Q�j�6��襖2����nvMn��r�5}�e���OQ�p��n�}�^N��E7i.l�Zɘ6�>L���Q'QըECA�LJ9�b��Y+t\m��|9�����M�r������������o:��x�<*�[�b�o��k���-��&�:qM�L�]ɵ̛a��ÒS���v�hu1�'�kF㱠���F��h�u�o�{�Y�����D��n���̧���ڍd�y�혧ww
���k�7fh���q>I�u�W��y4������W/�6h +���a�s �L����w������+�^nF+ߦ�u�|ڲ�8�*�ofajʌ�;-�l�7��$n����나�tZv�+���qR5zvue+��\����/'��x��0p����l�4xP���G=|4<Q�N�)^c\Lҫs��,�x���D�F%������tA˧�$Ы'`r����+��WvhR�]�Τ��5������?��͇U�����k�c�b@m�|���\�����6��ʃa��:�@+��0��=	vU��GW"�ժ��5���r��^� =;sb.��<2�R;���,j��t
�����3���Gc2�����@I�:��qj	���a��u�H+�E��0+tv�ͬ�;tG���NQ&��@�..I�\����[�|�Fՙړ���/��+Q�w\s	�7]�ŔF5vB9p�v�j���s��5���IކUpGZvL���-�s
��<ث1��5:�s(N4�γ@�w8��)W�_	+D���CY�xB@�y+x��&�#u�6x Gp� �E1	2�Q��:�=���9�Y)+���^�Ŗ��M��u�雾}��%E�'2Z�N�re��`�Eq+]��;�39e��_3��֎�E�oF��v�.�
�7�{5��6ML����	:S靈ڸ�8��)�Y�7,T�*֏ip��hgF]C���KV*ظˬ��΄un���u{6���F���2e`|{&w)��y�'�z�f�7���mH�bu��N��n����Ii.�n,hJx�u3�(��Œ0oJpT�p����Y�n�9�G��D<�v����θ���J�����J儓�к-ͩq��Z*���n���ЭQ���6f9ˬ�ӧ/Z�+0���ɕyn0�Ԩ9`��;�U����nM��Y��R�i���QNH�p=um3F�v";t&�A��+�+pf�Ah�:IݯH�$YE�Y7��v����+k�U���|z>���t�����v��u*���t�m,�Z('\	8��)V[�	hP9v��8�jrP'%�CV>�S����w�pS��e���f;��{O:mh�v�<���e�rk�l�įr"�c˜[��HVK�w\�F�I����8���^lgs5h��.���j�\�ֵ���"i���y]���(���H��ϩa�:�UXZ9X=�V�cV�[�̤{9ލx���T���[u/�2���� {ƭ6oKt�����U/yՠm���%�T�w#V���|A7QS ,78wW�q�T�P��n��櫦��[�������z�]�6LhC�)[K(팷�.�u�]ә[�8�>��l��`쏨�t+�7�$У�-lb��*Æ��!L��e�:�-uD��W���o2f<t�@Զ�;��
�P\e����n;�]p
Z�⋚vE8M���ť��H��M�V���n��h�)�鈀h;�0��25X�*x;R(j��)�[}p��]2�RV%n
�XV�.���1�:A��`n��)��7s&k�[]7{�B�2L�|���cE��3��8�`ZeZ�`������t��:�-f0��^��:܇���8ջ����7��·��3l:W�\���'�y^����y�ͳEX���
O�b���ueڰ�/	2����ؗ<B�����3�9Mm�W>�TۮT�kR��Sz�nf�kEn�N͘���{N�0n�CLbX��������o6�����b�|i�p�_p���v.�n��� ���b��oR�_ڣΜ� ���)#��]�����:U{}�i=ڔ���RAL�-<wԶ��aGr����+k�X�R�N��[����X�m�9Y� �ו�S�]�Q�� ��V�iXT͌7�T#�K[/�:ì�'%q�����Ɩy��6R@|�4���uxB)Ƈx�L|���ΐ	D����IiB�>K^·{
vZS�:���V���9xd�D�k���%�������^5:\�xˡ�4��h��*�*����0/���z�L��ȅ���J����3;���J�I��x2ލW������FYE��.Ӷ�{�;%\�t�΅T����G���y�vJ��.�b��=�Ƌ.�|��a̫\�v4�4T�d�eo'b��ӵXFh��d��%��ѱE�t+i��㥂���]�~n�S��Zr,�^��]��:ҵ�5�x�@��>���P�}�!Eb�9��6���t��t�\7$w���WjX�S25�;�N[���
�N�CqnCEو�5�-�1�*�,�ĺf�MY���v��x��ܡ�O�MM�w�4u���ۘ�LZ9m�C�s�؍�5�y:��Rvn�l�d���=�O.fh�ܭ�ۗ%�.EE�N��v<)�V,]pu���Z��V\"���}RRF��
ݬ�w�r����T�K�;3M;�n�ZE�K�}��-��-��x:@�]���Ii̓��v�	gc�Ѯb)W����Q���*L�c�^�W^hNfi�Zto�%��� `{���	�)�W��Y;�Q�n	�,V�=�j�\"�(%9{��kW��z7(w���$�������@z�j)Ϡ3l�1�|@g^wWM�&�e�v�`9x�H*�"�y�-�O5�U�V���bF����Ѝ�;�[#��^lk���K�ܙ%A:K��I$�IP`�q\�y˕�*`}%������G���M�w�h��=TF٪J!���=K��7_3�S�{��A�%�U���a���cG��GZX+^�F*�4�2�
!��o#�ƪ�㾲yrOwP���AGR|�����t��_;�=��������u�1�>���)+�3��ޡ�^g��;��J0�U0(��(�+ 2+�`�p5��گQ�W��{��4����ee��$V
�j�xI�LxM�U��T�Q�%��~���jz�y�s�H�{��ι��^�󿇞��[�>�����D�?3����U?/?8�?��������Q D/��_�|������?w(.�=�XuϿ�������{��Mj3s4�ҝ3�s]�[`��H�ZD���j�+;�d�#�a�� ,]Nɺ �@�M�&)iZ|a������c�}�	v�a����Q��SN.�����6�l�]�Mn�(n1�[T8��^Y�éy!1�ׅX�)^jB�T��8[�^��yu�N��[Ͱ�U�7�ᐾYrZ��~lt��oD�լ���%0+�ЩX�V5=4C:�:.��wh�K�h)\&��7�P�E�1�t`� �Kr�W[�������Ͱ��e��2�%�R3�vq�d��Uרʷ�v���%3�D�1�N�}ۅ�8ɣm�=[~7H�ܗ�Sl�ojh�V'hm`��loaUe��_X���*<*!��O�/U�~�MZ�;!ǘ�f�}f#td��dC ���dX�c�9��'�w�;���.���m�ZPţ o>�S|0�,��^:
��Y�s2�d�����Y�[t��m��$��b�x�����oE�K�ww�'y�� !z�;Y����LL�)=���eerp���P����Q�T�d�R�W/U��D0�T(�i��1Ubʁ�x.��9J�3U�5��W	�����}$&��{��Z���t1��d��1H�6����W���6�_*\X��FpQ�i���Ǵ�@��\����g=�9��c��������|x����Ǐ��Ǐ<{x�<x��Ǐ<x��Ǐ3Ǐ<x����ǧ�<x����ǏO<x��ǏoǶ{{{{{x����ǧ�<x����Ǐ��<x�x��Ǐ��9�Ǐ<x��x��Ǐ<{x��<x��Ǐ3Ǐ<x���ǎx<x��ǏǏ=<x��Ǐ���.k��O���療=�F�wG��� vlҨ�(�v��Z�ɴ��n�2�}C�GP�Wfi5}�au&�#vV�+�xި�XL��\����orr-�wuճ����M����uj����4
�]Piq��1_n!݃v�7w���޺<ָ�:p�Xvyf_Aw�����G�����d>�:,͍�e�S��%ZE�ם�\V1t��n:��Ya�:n��]��g)�X: -)ݱ�f���.�oD�v�6��b������i��P!�[��ejen�����v�����Ьڕ�1�\z��LmܩI�\N^��%��]H3�]퐦���E=��	:㲦*\�6Iͱ}�i;ͻy]Y�ݼ�+i>����3�k�p�?at,	4�� �-��S�����Q@j�:Ʌ���n�U�E���)q���
�ePޭ�K�ʬv���F��ZŴԢ�FĹOpևY��.\�J�2Z�2:�]�[�)�y�k+�Jx�o��[6�^T�n��ռ��)����b9:��/p���r�P39�y9(�q�*ꏱ��o�Ar��MI�2�*&DH�ޫ]u��]A>�9�3	XU����x��w�-.�&�N��cBv���=4U����є(f��h�u��摨��^�{���!:�K��!v6���a0v;'��۴ݡ�l�l<�ZP��V�^��{En,���{���w���x��<x��ǏǏ=<x�x������Ǐ��<x�x��Ǐ��9�Ǐ<x���<x��Ǐ><x�<x���Ƿ���=���x�����Ǐ<x��ǃǏ<x���ǌ��Ǐ<~<x���Ǐ>�<x����ǎx��Ǐ=�x���Ǐ<x�x��<x��Ǐo=��w����{��*�d;���(
ת�[�N���3/R�n���vY�Il3+kELA�n���
���]'S	����^���[��[kBč��Cc��a+:��[3[�����&>���W}����#����<R���S�<s��-���E�t,(�W�Y�	N�wb޽�f��W`�]Uҍf����A<us)�Ͷ��Y�d�����y�feM�a��E����E��Ж3���^���;��Φ��a��6ʳg
(ѻ�t6�rT���^���=s"CJ��3XI>e�C]жY�Z`
Cb��-��&e��M��L�Q�ѕ�xХ[;2l8t=s��1 0�(RF��ژ4�0�<D�J̏,�s�u3�v�[s-*'sC{׻F�m7Gx4<��e`����']0�,ن.�*��C�nn�{ؔ��?Zʰ1��ڐ��:�:{ ��M��؟�Ջ�93�Wm����F�h�m�ʧ�,��<{`��: �V*�9i�xP��:��=�Y��7�_X`wl�z>K4)��-8��)�b�n����D�N�ȫ�����+�'T	�zI�j54���4}5�m:����9���wd��9S)��&Q���n�c/��ZA�v���l!.o�;/y�Y��77)VWA���G��32�)o�^�4�[4�-r¦0�ot�r�u+�˶�cH�ZĲ��3a"���:�'-�qfu��v�ك������oQN��i��єy�Z�L�p��Gn���V��+��|���[y2�v�vn;o
(�OJt�ڽ�"�wj��D�)=����)��y�:i:�]ƍ<��ͺ�;%ܘ�A��@��"\T6'��0��J79�ܫ�,�g	�5��:����Om���s��� ͵����m�ʬc��mU^B���gE3jο"�n �_9*�q����s�AP�r�h�o��"�
+��v��]{�ݦ��]���ǀ�J�Iw�h��D �+�S\L%���m|Jƫ���av���<J���s�J^�Q�X9�P�D.����m�֋�R�(��~�]�q�gʅ`����\�LV�.�#�+�烱�N�×��Ɨ��e��'�B����"�n�UX��:��,�iVB�R�ed[�[�xI��s맙z��p��ќ�C*$1�o����&�.�(ɁRaJ��u��N����\RN�k@����9��IV�z�>Xs6���s[���@�uP5|���V�das��۬�Sn�RqqC�-��wyY����g��N/rM�+�������U�b���ױ�%��R�x�^���o���J�p��9إlT�k�봊����t�*.��1��u'L��,�5._D6�����o�`�C�y<M�۞�9��H,;;����=�秖��6m�ܭ�*�r��JvH�1�ո1[㲐��c�r�J����6�6k>{F�����	o�BC�Wp{%�EAG�}|u��U��`�YE0�g{Y<�g@�*d�"
�&�U�[�fJ!8-�d�� �q��Zt�����j����sS�e�Wd�V��'m8�iA��|hX�Itc�*��ӡ��9��`8�Ŝso띕��IWQR���9C�dw�u�W�Y���I�XQăӽ��.��vg[!�Υ�]�;�t�S�ӆ�ޠ���;j1��Y�.��6iV4rE^���h��ڇm�����V�5�R��`�(�
��O���6E�O��Ԍ[��kݻ��V�2�)6�=�pe_`vw�B4��`��԰�v(���-є��.�����P��P�K<�C` �C���=��1u��U�z&�S��b���.0;���NaL��CN�W-�w)���E(��;,��H$�An�js79\��w�R;sP2l�����9��%�����M�n��Ƽ����)����IeN8ݲ�{&�xt���Pm�dq�Z���/Cw�� ��C2��jV��ɓj1����zZ�SY��W�Jw�3Iһe��y�N��.��&+�����Sn�m\��Lo��n�͇0j��k}y�ZN�u�:Y��JR��[�d]jnp�X��u^����F-8�*���x=�ENn7wJ�"ꗶM̝P����mo�	��']�J��[L`mBs:ѷA��r
ϥӣ��'Ľ׸��Ky\��B]�J��{��^���n:X�y�XE������?�ܺ����mZ���}u�g��0��V�7.MEuE{M�������\;5�U�˧����	�yO�7+��]�`�W��G�n��§]Ջw����cY��cy��e���YŰų�KoCe]�
�-VC�`R�.|(%g,�w�ꋚ�]֩�g475�뢂?o����C�έ�e�zp:�p��Ƕ��b���9s�6�K2�N%�#��L��WR�}V��r����b�z�f4�_h��_
����R��Yګ�2��解��\X�.�и�,�,���w�I�
e=�ِ�W_q��!0�<Ŵ�m����K���ok@"=�B8cd�!˧��)X��Y@a������}�r�5�J�.�j�#YEMו>$#�Ô [��5�R�gIU�������w��vI
�I͕�Ae�����ݍ�S��T���VŎoPo��)�|�ցKL��c�ܮ�T�.}���vS1*�����v.�Ot�Vm/-��M�q���C��#��YxUY���@C�#��U��-Ѵ;�����q��Vo����9x;!F��:WZ�w2�a�������KE,��#5Ӷ��ahvo/��ܣf�IB]�%.�������'��ϻN�,v��c̛�<=I�eͥ��wB�)��U���U��Ӛ1t$�و�����5i;O��\��;��`���Ȗ���Ո]�n��-�c��� �%�7���ɣ�Ua]�ӌ[X\��h@.�\/Gmaa���WVB��Q�֩�x�x�c5��X��ufM�Zn(��F,����t�7r��K9Z�P(;T �
�b�]<��x�D�}V��)��
1�j����L���Ejw���lT5�������zG0��|�Rvm�(�s��'�-���ut�7�v�)�m�jb���6�:ce��]CI�B�ggN�#�B)c��` V�79�2d�V�7���B�6�ܵ��(:�Ȕ[�;#� �Kwu*��-"��oF��`44(Hr����=���w�����yJ%���\5<��d�37�l!!��Es�R��>�6�l�����:�zc�ggX-V�Z}�/�[٢Yę�Z�9��<\�|�U���z�51[%��*��wz�J�F�D���ub��X�BG��1��V�f�J����'b]c"�l=�G
��h�>��q�e����2�m���Hc���y�+�.������Iż�w^�:�N�v���I����e��i�4�,��Fk�:�����Va���)�ݫ��[�ނ�.���9m
��ף�	���E��3$ݵ1Ү�
44y)� ��� ����k���7Ƴy�#���3F����2�޲1���Q]$u�9�j]���6��b���Miޱ�6��:��e-���3%��'l.���+��J{e��ro��Eu��@R�F�us-��t���^R�cvqT=���\0��^:��g^�i��X\Y��R;љ}�:���kN��s�^)���,K;�,A�����-����k���Ro1�t��s)���
׆g]�T��P�*7���u�3�}���M��Y�AK�K��Vv��dZ��OU��X�M�CV�[M�]:`�嗸Wl>�J�v�.��Jq���7y���\
����1v"�m�Y�������[<�ʭX2k0�-��s��c2��Y(���uՄ�A��c��s��ܤo\�^`�u-����R�ѓ(��튈�t�aM���T�dn�>j�z�t�܆��)�LY�Vv��޾̭.�\hհ쪃i��R}s����X�\(��3��]�6m+/� �����{�^��s4�Fʄg;]�Lv�_Tk�tc�k�.�mU�Ӛ��ͦ��Jr1��
�3.nG�Uj�m�c4Em��ч��0��sB���7.<oK[,r<�vYZ�4�e����OL	��j��:�-�;�e̸�:�q�p]+���]u�,kH�L�vx����C��e�ُ{��:��]M��X��<"(����}| �J�ou ��X>A�DVfp
E�o4��G%�qV�JBa�v�`D�.Y�+#�W�q�-:r��C�.Ѣ�ʴ����h�tW�H]ϩ��FT�EX�ή�ˎ�*We'�u�;��3d:��[Gpӝr-F�����:0��\fʀUDۚ;qܮj*y\�����v�	Jǅ��q<�����/�f��^h����HF3���z/z��s޵�̃*��[�+b	��%!��}�U�SNYO��U��bɫ!�����y�M�q�8L��:�'3却�U�%���X�pҗ��d;n\�JŬ��X5�Z���v�k7�%ϰ#Ng]�tʪ����r��p���ŪR�[���7�e]L!p\��Zj�$*��A1i��N�?�#*���b�eG2��{ ����`y���s�y{� 30)	�3�e�9Z@��.����|rNz9���u�"����1xE�*�v�o��J}J��S���"�ȯ8P��c.�.K������9M���e����/ֆ
+e�nZU�l$�9{ ��Wn�=�
����1cf序n�a&�����oh����f��(�����5k��*��6�ݲ.������uw�rv9'�K(4K�^uI����l���D���-�5"�P��*��j(�a.\�nv�Hc�L$ٗ���R���wbo ݚ�h�X'ZF�޲w��c��q��y�r�9r�P��Өkn�tI*{u�o�!UE�`@�%ʤW�����Um7�$��3|E�gu�n���2�����i<�)����̻�˵VΖ��6a7��0,��2Fӫ��X�Vk�xs&�b��4F5�ز��U��)_o(9�<��t�qڼ��R�<�F�$��:͝-e\|��ѻ�M�����_��C�[��77�=��;#v=؄qýDG.��n�)��[V�N�u])<���g(�8�&�Ue�T��oo(aN���Yb�A���2����2��w���8T��m�l$�1�;y�B}�[n�����̔:n��x�����8wX�ç�����x�	+F���s��t$Ϸ�:����ę���=��s�����}�"#����O�~������gD?��IS�*JJP2%~��Aπ6��vKA��`��!Qt���@T�3i�v�Q�lդT�2�����l�\�N�		T���K���Ɉ]:UA#�ulx��l
TM|��˰;���<1oS�a\E{�V��V8�[�XS�)�ﯬ�r�@��f�!�PW��p��Nu��:L��KZɵ�'�k:���&N����N���x�Vs�:�⨁4* gG\��W��FP�3�*ׁL{�z�X&��X��Nk�O�J&�x`��c!De�_#�ʁ����*8/�Σ��>�X�)�ť���%w�{�7��Z�g9s�x��|,�t)��J44]�3Iza�$��[n�񭗩_^m�R�n ��ˁ��V�=;6ܑ`�R���)�J��&鐲g׹ɻ�Ť�.���S&��2q�]<�7G+��������.rwe����|L6��{�G��ֶv��IH :�;�)��+�]��~j� �19��IkĻ�	;�&��M�vlwv�X����ps�; �^�cH3���<���gT��ua����SE^����.�����!�/��;K�d��mFF��p�A[R���e�F ���o�N�VO:IU��B�ޫӻ4`c��y\#|Pa�΁�z�H�,����/��g�K�X�p�)ӏ����7�4�ؐ\�k��]D)�k0VJ���ɪ�@,T�/_%+K�'h��[z�mw�5�LIp�,��"�ã���Ko���R�N�Y-���F`N��:�Y9���VL>��C�tC���$� i� �f��CM�VQ�@���( �LQt�A�T۠�n�~F�D�J%��=�Y��D��M���Q�T|�5
�E&�E1I�f͞�jʳH2�E���i
�.����Ѡ���j��f�FA�$���&ǝ�H$�5`�ҥ@yr��][%����.�����@�HH�]XUn���($(&�֝آZ�`�t��S�W��PC�:
�)T�=IMW˨�_W�}3�����|{{{{{{{{x���G@:R�;�PҽH�\�x������������ǃ�>%t��	�!ԫ����t[%:�4��4#mJר���XS@u&!R�h �:�����Z-�4��t=^B�R�)�.����I�z���^�]d=������u[QmCX���TG�4WVY��O���A�ڵU-�w�I�T���M��u:���1TLz�u!���DRT��g������(��4�SE�CQIPMMQ�lj�OQ���Q5E�4�Ж�!��TTA5S�E�ꠈ�*b�o�к�E�,]��B��T� ��z�nz�`u-Z��f�����Y�[Q[y+C�ѹ�*RW�Ս����eGϵѸ)�X�$ӻ��Y��#�S�V�(_�T�*hRI%M��M
�)�6��/]@�R�}R���v��7n=���� f�����
�����*l=������O�	ʽ:z�Z�gwMC9z�q��Y.ש�A�ʞz���'���Y滣Kh�	�[��ծ9�H��9�D������/�G���Gu{^8�'��4&5���/qg�"�v˞�ϱ8>���>4�s��YT��x�t���j��{��������dvU�.�^2d��D�27���2����6�������{o��cvC���{ō�����|��W��s���k<�@Ǳ�31'C��}�}�79�M���Gk�t����~"��}J������q�9�}�۞��Q)8� ��s3�?�6雠b��y��j��g�+ao��_H�"�kӱ��w���t�q;��I*=lԗ�2��rv�U�u:�qˎ��`�r*��>�Ŷ+K޴E�3��&	8�f�$hZ����ތ<b��<u��R���kZ�������{�����Z�v��2�"қ���Y��8��Y�N�6�6Պ�-q-i�`�m��jg^T�;6r(A1������Ӗ�77���/[SQ`}�m�M��Ĺ�:�3g��U/�7N��^�C��a��2����F�"��B��oqo����u��**ٿk`'��6�����x4j*��"�ke�=��=���	�lg�*J	[U5�EO,�p��q5���[h��7
��}C��W���Q�}Y�ǳ�~����.�~\X5Xn�6�޸��{%�Z�^i`ه�#2�����`<de��7] ��J>Y��<=��&���1-z��UO�s�q�:p�FD��I�<���pŷ����~$ݚb;��8�>髨��u���:�X�����p�;�A;t�_<�{�g�3;}���w����|�3~)٩W�TG�?l���7�ӫ�Ʒ:������ c��0M{�	&���"�m;9P߽M��,5���Fj�ɓ��	����Ii����o�� �uR���3����>B�hςw̆�c)GfR�s�<�L��&���fy��Ϝ��}]����[g��MT҅�k�Nu��Lz؊�M��Ѐ�=:���P4+pgm�W'3bbW��.s*����==�!�9bæO1�_���׺5�h�t[O�K���}[(n��P��j�V+���{[�e:˪�_�i�v��'�����ͷ�]��^o�|�e��,B|cv�>�^�=&^}��u�r��^�/ϻ�=y@�k=��ON݉�5���by�Lc+��P=ң±�v�=�un�mV=������Eͩ[*j�N����'7<�-ӫ��'�ԩ�W�{*�77�s�����	�.B����.Jfw��ՙY]Oj�|���;+�~8Z�}�i�������ʩ�A�������'-��1�����)S���r<�Ȗ�\}�O���Fo��T�c��G6J�[%L�%�U�^p���t�gʌr�7N�ɝ�?gp�}F���ъ{��΢��?����z@'�N#��f��ڞ�f�^!�=��>5��Tz���ڼ�H�#v���;u=��MW��VWDz������^�+�*�2�b�����m �k�:����&F���u8�ٯg�����x]O�K8�I��^�}ݤ�r�/{��I��@�;�b��>ղ�����]/�mV�t4��X�}ˋ_�w��E2��vϫ��uݎ7v�oi�4��˼��e8E�U'n����S�u}�Q|:�pi�-:��d�e���Lru~�3N�E����<o3d�$/�\EƖ�� �2M1%ǶnחU���Uc+�'��������^�c��2"�h�����g=��y�T��w�}яg��Fzz-���܏Io-�1/e7�J�+�K��Urw��$��q�^���8����wO]�c������f�C�F�y�M�Ϋ=���;=��ޞ7���Gu���R��c���^/j�{zj����un�}��.N��R����9!oQ�}�xTt z*l�]�Oq�r�6ڠ0��0`�s�����K�G�uϼ�Ht��}�zo���{W|�N�w\+ғۦ��=�VA���W#$y��t4���~��B����p�(��N��5*.�+z��*��^_{�z s�m3 �z��oI���7���$wF����m���Q�;=�ϵ����4��>\FX޽1g-�V��������ѷ�<�p�����	t&��R:v�T^Ĉ�Z�3�S��E�N��9
�ȁ�B��끙���'A�F5<��]N" ݨ@]9(���e��s�lݎ��oC�/��%�Z��T�C�|�P`I������}�lꆙΛ�|���T�|����c�wd�1�d3�: �����s,W�=;>ˡm�nj��ٳηJ������*�1��}^��O��7�-޾�������4��Su��f�JM���YN?/����J���ӳ�%�y��p�oN^IG\p7�z'g*�.}�w�Ǫ��{�q/z;�L�w}����m�%7<�����6:E�DS6O�,���6}��ޒx2j�Wnd��z������5�;C*��q�j::�Ke�}��A<��;�]7e�k5��c���j̷�&�'j�"mWep����^�f�s�8$��;F��z;�5�'	y�I�'EK��@��'_��3�{NÐom/	ޘ�r�������x��l�a��ٵt�^�Vz�·^e��Z��ý��G��ED��ى��յ���X�����xC�i"��ǘ�['���p�'������ݱt��#����#���{���*_LJ��mr�y��V0��Y�9����������w��p�*��	W}�H�;)�Q��?Q��Zd��4h�q�w�g����l�N��yA8�s1�_���{s6>�s�:�x�Gw���� ��0�}-�#d�&4���[��=�a^9��"7(��U8����;;|�o���<i�8������
��b����#z����\m�������y·n�&q:���m<8{���-��s)�����)׷3;�.6Wu�`�I]�y%�kۤ������8*�*�����=P*� �tȷpn���1Sy��R�v��y^����|���u)�qV������G[o\}���z5C<'��.=����d�c���_{�[��ZX� p�mJ��t[�L| \@��s���$Y�r9ͷ�}=��m�}D��}�T���2����͆�����l�1�V�k?� t���H��#N�9�5�x�5�_��g�d<@���� 䥘�I��1%^jJ�.T��}���w�A�������D��j��DN)����g�}H���4;�C�W#��7X�iw8d��&s���j�s�Wh��������PF��������R^��~�=T��P�w>�x�%���}�Ԫ���qK�u��)�s���u����z$��ƛj�XĶ�@�c��MnE5��[`��G�f��x�e��x$�reR���������υN8�]ϓGd֠���^�W��zv^'�ު90zx�of�7�I�l�t�W?Yc�b�{��w�����=��͓B����:h��my���F�ٞ���S�!鸲$�G�Q�0�b5������t�U_T|�'{6D�W�6�h�S������^7[�z�M��+���sʨ��Cu���}�i�xt�Mmr����D͞*{��¦���K�)�p}�Hz���5�V���I��+=�<�Y���^^�O�Wd��T]O*���v%z����B�x�t�S���VS�\��~����r�߫�=���W�Z� �U�^�YF����7.bc�R�zԭC��m��j�Kx��)�H�f�f>�N���0�<�@���F���$F��h��wRq����m4�P]�%ʺ�����ǌNy��V���_8��irvܢF�9a�;e���k���_g�m;�*�hNf{�L1&�o�l����᭓�����>.r�Ӟ8'���P]OM����N=(f���d2��C��b+��4��r7+�tS��K8��E�Ty�cl^d���_ɾ~�=}�s{fe[Z��ٿ|v�^��w��^�Vv�Izo����K�N��#���z��"��=���~�ޯZ�U��ꗾ�Դ�sV�v׽}&p9����n��d���&���*�f���^,ͣq�g�����Gy���f���p�[;�I�s�&�<j���M<I����zB��F�z�Y^7%p���_ܳ�6��o�*ߧ��6RD7�:��Cw=�c9���2���dt�τp���=�?l]�~���,��s�u_�O�I���^}��ʺ#�W��l�y�8�zz�\k0^��P�d/G4�V�K��Z�&]�������ky�\���1�y��"�-z�sW�Բ��0P�-SL��㇁0��ks�8�cn�zb�%�+3��R�t��|��n�Hf�v�_l�d�(�v�G��FA���ge�� �:�#�����	����y�[���=^͞�����s�TͼγR��͊\z��^�oВ��y|�g}�YE]y)��n�?��Y����9��Lw���tO�gy�����>��OE�'}0��S���F����Ɏi���'n0��1�㻦<�EϽuS��?^-�Sud�Ү�r.������+�������j�{-�i��+@pI�k���}Yzs�����{�u��3/)��m>���ީ�J�φ�@���*��y�0�l��{����`��$?'N�v
:���:��>�(&�;��i{�_��'>����� DH��<*���9�����#f��&�����HÏ�r��y����k���vڪ͌�Myߔ8~=�t�(�*�(��{k�%d�D}�ŏi�����L��I�;�x��˽\�Eż�f�z㸰J޹����ۤnp2��K�_#��7.�l#U�n�vOS���ǚȲ+:z�o3"���;5.��ǳt��C�o\���\��z�~�/���:��)����Wo7��|(�Jn�z�">B��p�:���J��xu��m?SL��]X�x�*>�{�^�Ur	������CQ�1fb0d�_�����9�@��RDM�j��mQ9+ٶǼEa�-�'*�m�*��jޡ�;gK$��x�������d^rvc��v�\��?z7�/[���mҞJ^w��'L$k�O��}����a��a�����"E��!�u�՞�s�:����>y���y�����"���뽠��z�ڔ��T�{���H���FC����73�|�V׋�wI�^�}��roq�6� T����ó���Ϣ,ϣ9���{}�����-<0t���)�i3�}���4���6����5��c���`;潤x�f�2z<[��.���__�j���W��;9�k�U�Q�׷�n
����mn/�:�oD�=>��6�'��<���
�bB
ͯujҫ�����Os�ش"�K�5�W��=�W,]�I���XaN�����^
��u\m�m(��^xIp�{ܖ�o_a��b�ZT���|�������Yz˱{���Vilj������V�a����!���������HР�����h��
��ـhˊ��X�r�^�h����B��J��#&��a���6�3�h�y
 -��m�#k�K �ou���Å���u���.�m^i)� P�����{M��PeLyX�%��l��t	���l��M�]�:M�GW*y��87�i���2�1G(r
��D9����T��|8�i�Tn��y��2���-�N�$��ǝ�w���O#9����:���]Z��|^]�T*J��-�;Y�'��nl�1.K��\��X}��Ek�op���6ı�^e"�[�j!{J��Y��	Ck����
a3����r���e�ZD��;G]�T�4�*�H�Pb�]nEY��R=�3#1u�7)mY���?bm�<�;lݱH������ɴyX�*�S�,�@�j�X�q�fj^�!��PՒ)"�^�aϣ\dR��^r��r�����wh�B(�H�ұ����. �����N�ꂖ���ܽ\�N�P�^U~�V�1E�"=���]N^8���f�-f"����kt�c-&rE��4�҆ �;6���357؋�ڮ5x�gm�S�r�n^椄����̰�0���^*��UW3[B�s%ڽi�\���U���xǬ`Ul��5{����F����縰(+����_$�fLQs���:��v^��9>�4!��W��te�Y#+BU�deJZ��� �s�ɵ��A�E[�j��X&��/y�h�ؘ��kBh�庫&�ސ9yZ��1�r�����ihQ�lI�[��w=u:�E�i���^s���li�a�G�r��L]�GW2���hڔ�r%2:J�h�8�)��v}-Z�9\k�+���t���^b�hd5Q��6���cc3u���D�Wm�;Ly�:/:ݬ��)��V�:P��a����[g�S�-g����7H=�z��o�H���W�n%�j�����Gh\ઘ�d�Wy�#z��ԯc�X�rZ�y3��ޥ�tȌv�%6�xgXj�a�mJ�,C�!�m
��ʛ�kn��K|��'��V)��a����fV]�=c`��5�zx�up�(�x�y{��[
�㼮Ĭ�Z�.Ȧ��ĩTY/5t���Ņ�^�N�X"n�"�/jV:驵08;�'�G��\l��8,�W�h,��:��er���Ԛ�4PL���vu$�Y�{�	���x�P��(97	���י�|㠀 ������SC֍���,��/��Ȗk
�@�FF�y.}{K�u��fg��bVe�lT�]8͔�Ug�B=@(�F��Q��(�JB��F`�����*�:Ӣ�&��('��(K�=>�o=��������<~�����X� �{�	�C�ĸ�ō�(���O�����|||{{{{{~�G� �e�.�SԽET�=�z�)'p�(��Yh"�_!��U#�����n����UI�:��z�4�%RƱH��#��JZ�J��
��u�CI�z��B �� )u��:
!���SKE4T�M#Mz�T�g2R�4�PPRU4{ڊ��ݤ����I�����T�
&h����*�"� j`�	|����-í�x��w61Ffd@�ʕ�h&̾:b������I��=bV�]7��/��CMu�uM����B1C�}�����������%�T���]+ޠ�Y�(i�K`ބC��D�=N�O�苏>�T?VD����y�E8���,��^Z�pU�
ʜ���K�q�������+(��s��)?�Z�^L�	���0O;=�k�����k��,����&}�4&�FFS���s���!rT��A��lL�?#,�J�ݫ��${L���g��T�>uʘ���r��k��V0J��W��%6�mkx|�2/9<,�=G�L�g�o3w��$��L�
�1���o��w����0D��h�Hu� ��rN���(]u����P��s^؄9�%Ƚ�%4��Lߢ;����ϲ"����h.�u7�!J�75{Y�[�����0(��|rO=���$�ħW�E1����[X�a�P��ȶ�2�t{.������.��p�PP��q��������^p��^1��F���NV7H��y�5^O[��zR��s+�o����a�����B=�&�������0�vA�M���-="<�A/9J)�#E6�+2��<v� ,�7Y$>��F�(�b���rv�o�ثl�O*��^�/#Z�cX�ہ���*���n�7�6�O�1nu��e����7.�_&�_mp�.�l-��֫�B��*p�5C7�������9�;���F�)�:��V��5H����hNL��y�.�+�2\��Y�V�Z{���r�:m�������̞���Q�P,�YK.1�t���+(�h��d0~�vd�qɑ:ꧤSw�+(j5B�����Qև�_���ϭVO[�s{����U �3
�~
�a�h��/-�]6���g%��|����d���Kxu1����Wa������E��(&&=��ɶA@XXWv�����]��&���w�y�D���[�*�١[�i?��s4;h��b�-�-��;�+W��m;�kUΧwo�-�&v��S��`�^O����O��D� ��vv�0]�ȼ���Z�U�@Q?����]�y�0{�����H��X@�n9���%
ƫ�n�Z:<����	̈́�������הV>nLC���cPm݈d�5��P/6�k�"���2�cxC�["�&��^~��Z�w������g��8��VP�2�fϡ�!)?�����={6h��,t�X��:<٥��@KUK�N��U���/�s���uuEn��7�����R� K�[@k(���6���un�pP-�q��Z;8�ԥ��ע,�ֆ��̛8U/b���98�N�\��(�U�R����Fũe��7+�|�����U����5�굆��e�1`@�Wp��@�ݱ�5�vj�	+Y�uyM�Lc���w��R��{�p�,����{: ����x;�� c~=��](�]@�IPwe2%��!]����1�fN�v��iY�:��z�d�����������OVq�ah$���f�A@�{i|+��Υ���D�Vzt���D&I˼'<
T-\�)�-��"�^�!��,�����C�W�Lc{$a��e��oz]���T��1UM�kF�րK������Cĸ�tn�J�3��>|w�v@�!	�'�pG>_G���|i��n�F��,e��֜ٙP� zA��� ��5�X��H��±HL��gBo"���^S��@S�a� ���h���G�o8/�����,.�N��j��;>>��_RP')��F��晻!C���u��3��=��\h.W��,`ۊ��Qo
���c6<�����}j�p��l`�8�jۤ�ů`4^�(yx����f8*}#���K��-б�p;�)�(����B���u�x�����7�:"���T,(%sO����2od�{%���	�k�(vu^��
M��N��@C�e�[S.04��a�ɑ.�G�c02"D�L!�6߮a�'U���s�Kpb��T��3�S���63
<�j#�a�c�H̻H:"����^F����,"�F�yO�(EE�2]�Cf\��V�qX,����Z��j�]*^mw~1�0-ȵ9�Oq6�+��@�u%XK|��Է�<��P�ﮃ���v������9�k��i�{�k�&c\v�E���gq<}�ul��[�R�VИ��{	]�kn%�yd���������<��;]�4L�C�Pi������ou�5�<&|�Yq�hC,W[�H��yX���g:Qi�0y��P��9��B9�[�z�6����7���r�Yh��/���,����>����&��L�[`\d&�5��eK.��gU|��oN7���]9�/L�OK�Upe]١w�����ј�/����Gw��}R���%0|�&K�N�)�E��m/.z�om]�6���{մ-g���cռ4��;pN�a} ^������>����L��.Z�4��cfԭ�<q͸���	�Њ����uw=��ׄ�P��x��4���L�dy�T&]*�z�|^sB�-}������2���YT18�=>�{w�A�8�.�^�,١#̜���s�W�ul�n�g�lP�3	�2]�_EL/�J.��	c�z������wV����t����X]�]?ǈ�	vb�8Acr���4��5�p��������Ƃ�0�ԜK��HɶD_;4�U���(�2��=�لsk9�Y1)�	�-�Z��.��0����ʑ��Pv"�u�l�q"�d�G?H+��s�;U��+��̢�K���{r�����9�kH�SR�zd[Y�Tʌޭ�x]k]�X#��������Ƨe!`�� s�.yAI�#��p)]h�ͣ$��)�k^�pMA��,]��5m�?xxx{���gq_a���:)R	��;��1�L:�^��mW=E����ka�ac����%��Z���ٻ<�k�K�[�uԒ�c�1� ��-�C�*h�L����զm�In+����Vw3Y�C��5�O��?�G���;2�h���c �����{�t��W���F��ȡ!�NX�<����l!�fw+:|�@9<�����^��y���� ���!�ɉw��0�Rq�
�f(����l���++�C\�ô�+��{y��b��C2�����(q4�>��o�s~�����fڠ�gl��$<Z���`P�a�z��^=��:��W�d�4��ë�e)0���6)a;�m��춭j�ԫ�)������ɑ��J�S����W�|���T6�A���
�R$<���$�E�C�_XK!g}�a�oN��V=[¬�c��kG�8^D\zJ��	d��d�Zr�8�SWfo�<aC�m�Mit�dԱM'�Q�ma^=�Bޭ�[�����>���$�* �+L;����ǁl�&N�'��(�E�P�2�&��Gc�sS;y6Q��S��b﫵<=fB��+FR����~��C�� �
�k��-��	P��,�
ˮ��]27���؅�8=J���vN��:o&^�Bƨ` JkW����1��+���ҕ�p��x(���sսwNəi]��+!��4�A[�x8֓�r�������_�o���I�Z�x�k<�5�0`gq�p�;$�׺"S��c���tޔ����$�5����ȸu�ݤ�1}͚���k�=�x�T�c�9�&��v�v�����oI�]-���$��W7�6a+x&�����ÔG��מ����y���Bm�1��og��ŬaR� �&�z�����1
Qi�L�v����/����5.�`��,QH.�5ٗP�1�gqs9���«�����D�1
�ޱf�(D�4�mS|�7�1sU$3���:<����L��d4ug�"mj����2.ծ��=��ؠ#g��|��zR~l��o6�� j�e{b�ٶF��� ��񆬭b�F)=Q�A�n�=�����ټ���T,�s%���Ʋ��G�8�s����H�`�6�)h���y3��x%hkgR"ذ2��ߥ�>ȼ4#s����0$8��	�������5���zR�-�vK���|�#��Ce2�<J,h��!��^�K���J��^�>U�N	�%5�%ŏ����\ڧ�����{��.��4S����@�q���:�&-����= ^_P���<#A��)r�f~17������h+�#4{�8�q��p`�0�v�Uʘ�����Γ��7|�^���thS����\�ͲD���s�C��P��p+Ax)R%D��X�7�c�j7�:���Eڤ;]Z�N��39�v[�{�At�Wo�u�̓�mĳ3��=g�F��)���P��M���oWD����
w����B1�[�l�z0=\����KC$]��C���m=����d!���\�ԑ�g���4w��J�1��8��S�k����gާXw�^���O�Nχu�EcP����@t��%�;�*+Y��:����Ϳ�4���So%Oo`MD`RryP�����ezbw�!�Ɍ�y�N�/F!�{��Z�B��TXS-����ۭ�mۓj������)���Tz� ��t&v�{,�&�SsWD&I��Jse*��N�8���uSOY���Y."uŨ���'v�:u� H1��qb�S�.�E�K���T�uO-1��n����>�����ڵ�+��EXNb��] ��-�F4Ð��� �y�%��SgpeqW1�;-0��/6���yk�a��2&�{'��,+��` �kϡ�n���/���uk�놭�<���X�O*��a=jW<5Z�IEg��,Qن���|yS�yck��& �5!� 6��n.�����"��̜q|_�K+��ͫ�a)��Z��×�M��?[���6�Vs9nhv*��Ӱ��<���s2��E/���U��g�	%U�Fk��A�����zZ�_�����Z|/:֦ �E����۲�g7V�j;�[J�K�*����d�im5���%q�._kyqX�y4r]�n��]��1�@�{�4�z��`��1n����p���eH��f��0m�q~��~*	{hO�N�qnh��T���Y��DZ���WBW1�࡚<S΢�\�s^�fY7ԘkW���M~y ?z}�|��'��cy�0i��w;�R�RŨ����a�9�^�P���t�u�\�K��T3e�vI��B}�^������1h{��0^J%=
��]�^�3.�3D[��_Z�t>�yO�-�]�G:x/W)=Wf��:�!����C;�|��T����\=2׊xc��s�`^e����JbEY-�GP���p�Q��sQx��3cZE�$Z��A�W!����6�e�7K�:�m��i��15)\��X>�P|`�:.&.��_{G��[��H\��0�*Yt+<q+�p�dl]��E�~\�-���t<�޼���scN	������m\�Ly����M��&*ZY�Z�uDI����7;sY���z��M:����3�iᶞ���,ҜI|������7�y�n�'ܣ�t]Yרԇ��D��Ţyͥ)�<{���]MR�Z�OWM%R�Tƭ����?cᰫ��2�*.����x�Sɣ�w��2�U�Ќݺ��hʻ�-���w�H����lS�4@�����m����� �&�0e^��F{ H�$t�|-Z�Vj��#�5���Θh��{Ci�����Ѵ(qjd��Cޙg�������_U)NC���T���bD�>޺��I� ^%�u��c^(�aO�\ᮢ���H0͒e���2���c���=��'^�(^���E_Qw��������9��[���\����.)�XsK 'I���u<��@H�fM0�su	����ƻ�g=�I�Ux⮗�Qi��rĮ��I�z)�����Fp�2G��8��d���֑Fk��IuRe6{<�}DH��ݓI���Ҩe����ꮝ�
�h��n�9��q)�5 ��=8x���a�G�2��xl[;E���5���׌��_�ڵlo-o��1C�f$�c�ܼ�ɅZ�$�W� ��$c�x<�<��������B�a˶��x���&-��]>}I���>�t��@;R�hņv<ᚺ����款v���i��V�L���6v��dq����@c����^�"�@����ų�C��tK���x�#�׭Ew1~��=���5�ĩ��%�+��6��4��$=qhO�i/��ʱ�i�#��Up�;�����=��g�3Y��SPl[H��I�z/��n�i�h�-�n�V�@F�����ߠx�2�ev]?�4kWL��=��]�/(P\�
�r��.`�B$=z��9<s=�uk2��b�9-]�:���
u��`
���Z1��ӥ���8U�N�Qr�A�v�gD����C�/!��/��8pG��uꅥ\._2�No�rk��
(B J����%C$=����6^�^n�[ZY�sK�6��X*���B�1�ȥ�p������q��BC�^J=6��q;A�6q=cռ*��[Xd^�=���
�X���oh�\���oX��VjP�W���/R� [m�(2e�%? ��Xz��P8�� 5_����e�'�����P��z�d<Xa��dh��k�����(�E�$��_�Mw���{�Ξm��i}#��]�;$N���z�8��N��7Q�:s�'�O=tD�I˼'GT�cIMl�q�/r���;wV���ns���-fӄ�L��m�·}�Y��2���q�Z�N]�>$�Q�=�ĶaO,TE ���|}_<𢮽�*�Oop<�>h�G�9�h]Oܨ��.�rt���R�і���t��(�`Cǟ��W��)�qyT���=�*�>��#Y�K��1
3�W34�:�;F��1E&�2qx�n/���q���\�I�iF:(��t�ò~3U9����:���N9^��M��]V��>�������x�[�Ͳ6"��r��KҨ!z?/���Ϝ��[��2sQӋ��)�5CKm�r4Y� |��!�0�(��2龾�fI	ݘVm:+%Z���xT��:h���|`f�k�ڙ}�6�4ЉWE�w;�F�j��z7c�|�grm�rHEb�ue�/e��rqKv�7���;�j�G��8o��Z��씋OnvH6먢q�BR̲ԛ�3���M��ʽ�|�)��B�7�E���v�
��ھ:��ۑ�8;V�4D�d\���88�u$y@86쭟���7gsKTyg�͇)��!|�(��X�V�s�u�H��֞��]���@����l@�[�×I�E\v��yi8�b�����~('5�d@V,X�[�S|*aΔ�U)h-
��u�>n���T�����.���Mwvw��bM�Uy��Wr�i��WB+2�CtsV�-q&evf^�K�Y�o��Z�݁��)��(ٓ��K�b�j;F>�6p��� |:n��k�亏>���œX�2�@���KK��g�=/,��T@�;�̙���FPe�vo��-�z�7a<U�J�YxS�Zx����k�)u'i�hw5�g	CK��K��A\�.2��lf�t��@X�;���IJ��{�1��L�˾���G�
,t��9��uȄ���ˡ�+z� �!f��uڋ��sVM�ᚨ���A͂��RB:��-��BQwCH]�V{y�/�Bɠ��[׀轒�hr�D��m�J�j��n:�{���cAԶ\tAt��ܴ�}�D*2�����R\��,~���G�4�<��]i��Z�i:1:<�ݦq�{El�Y@nI�[�{J��b��LYV{�ӛpGA�2��Gv5κD�zĝO�%bօ9HB�=�'���b���k�M�;�6�o@s�ByQ�b��֟B"�w��uu�iQ�T.e6%W�QS06�_h�mL���*u}�k������R�"�P&�L���7�=)�wZD륍�Q��;m�C׫��d�i7r�/pT7���:�� ��˟ f��Cg2�S�;vp�-ug15�B�V�K5��K3X���pc<i�'m���`j�A53)L\�� ��b���;��wR����4Ԛ�.��ZNZےP��v�p˾?��yЊc�[4����팫t�:V�7�N��^�])M�r6���v���Y��¦j�FN�E/��e�gi������975:�Z{��_)��9��L7��c���_^��ł�̗�۾1V^e*�_C�Mq��L��&�͕ū�Ւӫ4{��+P\�^k��	GILd�}��Z�/�twL+R���J��o!ިmG�b�M\��hf�"��{x�s9���lv��t��6=�69~�E�#����Y����G���3�Ε�NՇR��oDM�r�&��#XNn-��<���Zo������T�����HUy[H �b��y'� ���t���X�T�.���fs���������������~��r��ITUM͇Y���&&��("b'Ӟ�O<x��|||||||~�_�6
�*��"i�QEy�UUT%M�i�$UAQ%!ME��6 �H����R��*�b"������(*�(H"�"��((}C�*�"��QE媖����oY�SPD�A1APLD����H��)��"���
��RUU%U>��#�1h�gTAETD�U'�5RUQMDDͣ��IM�s5LTTE4�N��;+�X)�N�	����枩�I-W 3j�6�#)S2���4{��*If����8�\��2��S��В�+�GbN�#tݮͤB�(x ���0X!��Uv���:h�(4ix�J�����~�����ִ�ћ�����5fj��=����[��;c�xfO�zk�͘��W���:����۵R�k�}'V�g0�����U5a��ΑɃ)��:b�!���z]����F�Τ��%�����1\��بҶUvڮ3�D����^à�2�,(�P��Mm/T�Gw�W��MfLIv��_�L���c���'N��UWg&in��p�DZz�x5;B�� �4ds<:N�L[e9͏>�?���Y���m��	B�kl��>�n^)K��}k.y���%�уA�S�#XC�[aw0����]3;ol-���>:�Ƶ��A�ل���!������β��l����ʴ��;������%Ї�z`�p3teEcWt ���A:�e�׿{����V�v���!��g�8Ob���#DN��xN��:ɨFB��t[���XZ�R�TXSk�nvU���d����b/�?zZ���,y���kҨE	���a��_JnnwL����Q�Oj���R�#��Gv�����6@�')���M`�td�B��4p^�7��ýq>+��
��h�~xQ����f���L�mS-,�;[��4m���O.�U��븪o�
�V�}�[�_��Ν�!�U��ʜ3"��f�wu&-�n��QZ&��(�hfy���-�F��ځd"�LT�vɭH��:`Kt�����(Q @;�wך�V����<P��y��\h�?�l���<0��B1�r�D9�e���lv�S.�C�wc���s��Z�I�S"�s�e�\�6�{zX�Ey��~a�K�~|�L�-�t��1Χ8��\�'�
8e0�es�W�\��`�,kҎ�0���L8�	�|x�f��h�C�Y��N�����8p���`�a��5�[`ۊ��[0�]<�oԫXJ{���Na\�)�_�v�W4�ép��p|e��� �c@Ll��B��9��:�_�k�PK�"� T�j�'�z��0�/�d����#�f�69��s@L3,�{I��g%@��F�g2N3YvuN��k��R]�i� #R��z-�W�NA�N�\��7}X�*7^���_rs�ے�U����;�]�����/@�f�z̻I�Ž�)�|c�]�!p&tFP��v:z��eVI�ݚf^�!��ͧa�-<�ސ�z*<�]��D[*�D��~�������� �m���D-��P�/^j����5�myѭ"�	-B��%r�gͷn�}�Z4����6<�ԧ\8?5Y~�/��f���O�g٨&D�@��N(r��55V����]n	���n�슅?luz���9����N!�N��ԡF���l[]�/f��u�o��J�])�u!��:��O�L��}ē;*����=z��w}z��w���>?��s�!u�K]�]#�"��â��� ��a�8{���/m=�U-�K��υ�dBˡF'�-T�G����˝���o\:ӌ$j��,�~S_H��w����Z�ss�	�us�9;ld;�4�5�أnr�S���K��]��O���ebϫ�i.'�*`��mB[��;Vje=��;��Rv��'�/��2�&��`FNc־��z��4�[Zt��g:3���1�&7ތg��]O4�Y5�1:,�˸xA^/ʖL+ϱ\��a=k�gW�5���c�,��d͊#��.Ct��"U���E��t��Iu��@1[�L7w�u9l�}�Q��fnV$#��hup�5�pP�M0D�p��_Mk��qG�TpZщ�^�,fX���E6�N.�͌�_���Ѷ¹�l<����x.����-�܊��Q��G:ˈ��Z1_��ͨE_�v�ڐ~��ʗ�(JF
��������&�o9����������&Ţ���)`���{	A/r�UԳm�l��à<�!�kJn�}}�;=���<kq;3v&�N��e��W��:Mɳ)�'�L�s�����-v�((��ۿ��\h�ܧ7X�3N�C�}�v��ss�N�_ E�o&JIf��ՓL�e�̛�s9&.Z_@�iA�4�:n�0A���Y�C�{�3�8T�p�/~s��~=����ߟƼ�����c��q���׎���}�_���1&,3����぀����Z��O۷
�Յ�q�{�n}���;�����Iz$@;\b�t<�l�X�c�IZ|g�s�/k��9���ԺC��=6^���A�}�XV0v�oA!��Z�ǩ�+]�	���)�jhN1��"���D�ǈ��҆Ai�=�O^��z7��ӛ�@3MvIa�r�Mƾ8˷���օ˜h.��G����E�а�Z5��;���X6e/�;X��DA����ɒ5vG)d��)8;a�jq>4��ΑN��-���Eǧ����^c(䶛����;L������%6�1�{
�u�x�^=[ռ��t�̢�a���r�nέ���/D����:�:!�D�/a%4�ģI��;���_�4�Xs֝-�˝�X�(���pXu���B`�S|$��H��ޮx��9w��	nIMm�'��wvC�®��/fY=�����8�{�1�J�n�L�>���Iw�e'��NT��N�|����I���jذwA��m_(N�N�a8�R�	y�j��iJ<&qۢ7U4M��I�*���j��Ҽ<�`���k��t(�ee���]Ʀ2�&.����*��g_ϹTkfm�ч1u��3!�R���2>�+ݭN���W~�~J���8Q3� 
z��ߍ�5����k�����
���XsR1e��<�>h�B=��sd��k/�
�hv���֨���O
9 Ze�;�N�	z\^GR���{`o�kL9�C;-w��E�C���K��u�1��֊@�/����x��t��;E�7�s;W�@@��1���Wk�j���p��Mވ�BdJ{�[��k��I���o*��T���wf��荜ոۚFe�2������ C�r^��Ȥ|bK�1�e�c�O�l�z����sx����n�M}�n��Ļ���'l�`��Y�3<!	�L>��.|�6�r��JpStK<H��r�u���s�.R��{�GU�<	(�����S[NpLm�[����:��1͊�b�S�X�}��}ڢ]���2i�'�D]xŎzǃY"]����i���_�-���-�4Z�5����g��\/Y�5�2yڼT� ��˴�o�i�m��ȧx�d!���T/Z��v�O�[��'��J[9К��m����R�(8�����!���=��U�-�<�����e�
n����Z4�݊�Huc�J�����X1[=qu�uo���if���1#"�\.Y�� �Æ��B����gf��-��͛be��E*����ev��8��w	��/p��gYO���]����4��O����V��"��\��u��P������P{���x䗕#���B7^a�}��.[��@.��^A=,�,h�Z�~��)s�c�dvs� ����C�w�T��Q�R�eLO;.�d���D ���q6�b�Jx5C�t�Bݝ��Uwj��h�w
�S!ݓ���p\c<"z�"�L$�7���o�75tBd��hƛyyU]ֲ��c�ns/IwP�~��q��$vE�*8ސ_��&�[p�����t�P9�۸��W{9;,T�1���K�x@��eٲ�X�#�!��G��e4;����'�ȷo�nz��?}�i_W��v�}RS͎Sl�Ŗy�i��i��3�,Au}~��W~��P��Ư)�Mg��E��5��uc��\hVޚL*�fW<5Z�E��RX�GjJxw�m����N��wm��K˰b܃M�H�	��	y�Q�Ed㋾*�
�y��*^��	�lMe�gK77���b��qu�dhV|0����5��5Q�4-1�n8��ǿNI�MQ3�w'튻;�e鐝�öDk��C��D38C���|.h	�e��Z|��[ָ=���h�r¢u���٘9��*��H���M�P�e���$���+)n�u���w�Q��vw*K+�^i�kz;����ӷ�s*r�r؃��������o��M�ۼq��+�fnWa�AE�mf�rn����Y���Ϟ������U�p��u��~"���}����O�X���hR��z��Ɂ���x�	�<F��;W������c׺53qzZeح�,7�bK�0�q����iD[�@�r�5��'�)@�h!�-}y����u%�
Qm��|���5����o%@A�t;a�ʺ&��m;���.��W.�̮��A�����@�'R�}���+껗fE�����}sג�PE��;�
���mjɞ�sF5�5���&��RXT܎Ьf��t~�=�R�"~��Xڼ�K���xaO�V
T��=m �xf�~x��u};��zq���Oi����&Ƒ�`��q�_(Ɇ�סL,K������|�ኺ�k@.��ib�I�Wm�zw^�=[�S[;X@Ŵ��5�!�xizh��Q�ۺ�'1x���=�AL�L��Nl)�jU�wWYq/Z��8�m
7l߰0���w�Z˂�p���q�>�5�脝p/Ⱥ�s�1(�aϱ\ᮢ��f���"�J���E��,�t3t�!0<�.Cu��/��υ�Qt��ʥX9��z����/0J��i��f����|ׯ��Ů�8��3�D` �7��.���~�=;~�U-�~]��{�3/�DPU}�L�d{��pb�����o*�>��[��F�0̰��&>]��	�z�Xh]i���۫ayK��3/��J�L�X��e`t?��UU�!D@�
  ��ɽ���yݚR~p��頃�� �M�$�LhaT)_�W;����^�E��Y���:��2aM(U\�����wI��f���P�\>��@`嵤G�� Iu^�X�a9B�?4�;N£��h�i�j]{�	u3��6��>\Ae �4;##q���ؙe�)a�S�wWkU��Vmᖶ(F�c
	t�{*	{����<���k��?I44`<�<^���G�w.��6��vd^Ej�n�G*Lm<u>_�O�^����0>��(��*�����Yg&_um�xаR��4�z�����S~~��!�gݒ�����Iz$@;���v<�LZ��!��4��qMG{�Dų�`R؆D�ŇL!���E���t�d>�M���s�ϸ�54Ѥ�������������V:�c�[�rS��dΊ~2��%)��l�m7:�������Y��k`�(a��q�%
=dW?s�(:��^��0�W��:X��ɯ.7��(��a���^�nq�B��fӰ|��q�j	���8��=[ :Eg�0��,:.���D����Yf�P�W�N�ov�c1�/�bʑP�)���ߠ���
�9��z����e?��#{��� �C
g=Q����v���������F��Q�3
k�s�,��P�y��Gh��9�N�4�q����xNK���s��VJ� � (�@�B��;ٻ�:�;7oq��/2�������w�\�m�j+���o��ɖ(��૧Xz��oV�^��;�5���.̎T��P�)
,#��{d!C%
��t���%�:	d�+Q��~��������x�cՖ;��w��Z8�'"�`��1|�"B��-�nw��?a���	e7�\��G��v�v��A�f?��(���^gJ�D�S},�M��q#{�fԼ�ȼ�5�z���֧m�o-��A��8g�Ñ�>�p*p�.����K�a����Xkc�K�\��z���Vtu)m"���v^&1�������	z���:���?	p��)��{n�#�2�k3��?�&�%R�jZ˭�4�xMs]�R��Z��a�{^b��I�󔋁��#E������9�5���u��D.rzE7W������)?5��o7�s��FVŻ�k�֧0���G9v�V�����vh������;'��%�_$^���a�Ʋױ���y�>z����Jb�p'ʱ�zE����e�q�.�;l�`����LZ����	vO�/M�ԓ�i��A?b��7�-���in����<:{u�v37&�EX���GL�p�o+�ĳTׅg���8�LUm��jB�ܻ��K{�[��K�+!�T�p{�m��r+Yy�:ZwS�{`�~����W[Z,C_�T}Q=�WE)HC�Ǐ���?��f�ݭ��&D�f�x|��?���r
��D{����>�|�����M~a��1�5���{��h�gl	�_�ac����J�m׷�hW=i�k�����{�dJJi;R2�ZG�tԸF'-�K��-�<�ç��,�K�'��>�P���~���
3�{�7�@��A�܌�[kR|�x5�)�0�0��t٩��7��[��	��W^mkOl$Pa�J���Q�g��6ʽ�-�;Ү,��pz�+�K��X�"�<ֽ<�|Ǧ蛚��QX���B~k������ƽ�ֳ�y�Y�q�F������}W������G��%{�r��b$��]Es�������>��A�=��Rt�L��\V�V2�@��Q�]u�)��[`���sB���D�E�	;M�p���ǡ��R�=Ik�oV�i��x��T-?�J��[�[����8�|�Ƙt���!��|��¿>��7�w�d�y�� �J����|��-ށ\h�ύ�!K0�W��K�~�����3+���]w`���}S�/`Ku_v�꒞lr�d]`c�}��F��vn��k����k-��+֙W���V>�jmn���T��"�s�O�;x�[wi�6���7�)���kR� ���ToI���#�1#t:�v�9�=��9J̡W��v�wm�ݩ;���R��`�CG�:+a�f�n�}�u��w�o�����F�`�ݩZ�Z�֦]a��]onaW�L(Z������b�3�`�XB�9��!m����p�7ʃKt!˝t	�W��vb+њZ׸4������p�j�]ɬ�8�0ŧv�/uG��ra�5�"����ٌ�
t�rv��bL�˕ǵ��\r/غI��T�뫫\-h5���r��:m���/��c-�\
��t�
Ǡr�*]{�)�kZ���B�2`(�_<�XF[�VeH�1*��q>8d#���n��M�ׯ�h��Jp�' ׎i������t��{��ܾ�]axy��d����ۧ�XA��s�}�����uѥS:5YeU�����>ĞM�Y&m���!�׃�{W�v��7�J�jAU��X��w���9������θx��>G]��NL�D��y�&��r�#�Ă�39��^rN����T��ɹ��p$�S}�bz7)�U���p7Z����.���E��nM�;N�[DԮ��Y;&��i�Ki����f���*\�����w��"�j�S��v�qY�^J7��h�Ǣ]K�Ԟb�a�w�^��x�x���{���������P���ėڲ=�_B�>w��j����d���`��(���SB*Yu�xGK�P�p��#ᶺn����ֆ��E���ԉ�w�1��Y�kb�PQ�e!�x�ڑ
c������NGč�t��ν}}�n�Զ�w3n_X1h +b�(u��h��ܮ.5����2���1r��j
�ޡY�6Y��L�����֯1Kth@:��z�.��B�ӕ�ID��Brฬ��,�^�KB�P	��R|�r��#F��]�VD�{[��r���˦�zv��y���X}Z��X�2�	
����/em�wy<�i0z[̶���ޗHSܻ��=a��߮�ƟQ��b,��%:XI�<V� 58"�ѥ��-���3P5}B���=
jY�����蝻��s��r��vl�O)�P�Y�ЦY�fl��ؐ�u�{/�Z�Mm<���"Օ-l�q�x:��*������G#�u���;戭&�ul�l�j}��%[c�2�J��6��wK��0�ȗ^Iի7],���)Wke���e
Q�e�x˼�3�N��6���;�c�t�_;��,ň���T׀v�Zub�J��k���cQ��o2ԥ�T��a���sN�^#��_'|Ty%b�f9�����)</t�t�����.��]D<t�'l��F�E\�Yͼ�ݰ�yo TivIs���Y��O�Ļ���gX�a��g7�����/v���VU����������*���*J"���� � �������Ǐ�������������������2f��j�����j�����Ǐ�o����������ب"i�`�����(�	���*��14�u0TMU4T�IDSD�MU��E�˩��(����E�*��)&�(�j
i���)����6�J:ƨ<�&*J��54R�PIPV���LD0M5E�D�؊��b�)�j�.�UU0ı�5LEE.�(�����n�-��PMC3E1!C55PTEPC%QOR@F"&*����cQP��EUI3�^�
���w����g�9����e�e�s���1�S�ˣ��g����:,n/������QK��{�nf{��w��UY��(�s�@_���~ba��Y�:v�����*]6��y/��D�i0�es�U��^o�W���>	9�,* �ݘcq	n<��ռf���X��×������D�^5�Ow���s']�����c2�f�:�i�!D��͓ں�|�A�#qoU�F��� AC��-_a�<k��@�0Ԏ�pZ�2q�d���l��kC�Zڞ���R]-�OmbQ��Bu��ÿs�8G����0��/��,"��k�F�ֽpi��Cz����5�c�<��o�Է75轃燐dK��tƌ-��f)!��!N�C�g?,�v���-�\a�&(�f8��f]��D[qL��k˺�%Im�8��g����h�%P��z�='���ͧa�,��@$? TG.�iD[*j�m��rL�ͭ1�
��f<5+���@�ˌ�)<K�=5��m�Z������B�{�51�����R���◙�t��ê�E3�[�'�X�/�=�U-�^\�.sP��к�n��܎M�2;Er�Ԃ7B�Ru��ޜa71P��3��Ƽ=K�/5���|�uc)��7|.#V���,��M@3��9�&���]q�MҔ��a������)A�i��B��N������JQ�o_`r�vޯ�&Bޠ���i;�K�Z�p���U���@�����꾤���K�h����߾y���O� 7 .s�=����շr�-��5��!2��Wy�<����3�i��gb%�/}Y��H�,�v�_��w!�/n׸5�=ϣ����Y�:+e0MBT7ٞ�>��~ׄ�o��V�#�6��g�Ahm!�L�����|k��	:���u��Lhi0�خq����m����S=ۮc^��HP͒"�^�!�E�*�}E���a��@E���9t��o��fM�n�=�����|��t^�@;>(fƐd�Lo�ۤ�B��4��Q�].ρ�vh���5״�G]���A'y�>k�)1�a\�c�B�fC����1%�H�X��J�5��i�Of7L����J�;�R�/��O�P�zY�}�e�l\�VFt�p�me�;�+�	[��ݞ�e��[
��kn�B*���
SX�o�]�:��%�X1�c&1�A�{%�P���綔PQ.�;k�vf�{��7��I��<u>X�>�~/;;R�hņv9o�q䛋v�;�m��ye`<!����.��E�l��E���ƪrC���+��&-,^C�)�:�wbw���=�%
r���LR;�v���0Mc#�)���W+˕���%9W�P�:wn���6��ԅ�t�Ĵ�p�pZIOX1���5��U�`^�n�ktj��G��K���'7#x�<���Q�M�&�p�D 9!@�� ��F����w�v�0�9)K��I���7�t6o��)1�x��ň�6^��+��g���q�!ժ���[Sf+VF�M.�BB�Nӊ�TL;��YI�C��ɑ�����;�����k�Z���7ő����Dn���~�LԼ	��PG( �p��I��m�^Y�X�iiABi���4̹�b���asQX��t��t7����4���`[R;A�ٳ����o
�N� hq�<];�0����b���d���5���n����Jm�`e(2jX��ڮ�a@�^=[ռ��-�?8���3��Vv-w^�`\�p�ar"��l�+%W5�B��rxeO�%4������o4ѝw�pd5,��}�9���K�[�c���Mb%;6P#/-0������~z�Jt���|~�o�U�棫�Cr;b���@�.�I��F��P|��\�� ��cT��m���/��)���],��(�ͨ�,��,��Y��U��E�%�c"�W0�LYz|�(�i�A�(Ba��&86����o�ݖ��YC�������i�i!7K�zOȄ�	z�ZGR�@�GSL�2(ֱ�7�m���Љ�B�j����`ƍs��P%y7t���0��t�#Ko
 n���k�M��AOδץ�4�u�u�-u���O��5�tj$%�,?>7+L�68�]t��$�*�Өq�e'GH�lZ�~�0�ͼV�| +��jw��o}�����>B� 
� ��v�<��oP��i�O[]4�yʹ�"�J7C�}�@'�q�K�@��v���mC�T-�ݚ'�Z֟6P�(���zE7?t�V{�R~lF<�� j�e�Y\�R-��ov��R�lC4K�d8>�����!�]�.��"�д^��5���]>��U���l��r[ٱo�~�;(��/ՄPp0>�����Fzs��ܑ{$�����a[�x��S^u�)`��i(�� ��Kǀyt$,�������8��H�P�Sk5��f�nF����ݴ&���v��]�q~w���<����.�0v��v�?G��ЯXVv�2�?[�ne޽�S�Nsc�R���+����A���kmjO��o��)�=K:�y�n�ӵk�c'���Wyz��|�nO~����l�,t���g���ɰ�
��x��Ӭ���'��µ��u�&�:+D�屋�;��(Ċ5#T����r^m�.��^A=�%�D�K�kK�i]�wҝ��3�����2�����f�]������i]:ɫѐ��e�4?���,��D6Y�w��������GKM�[�i���6M� �k�w��Q�u�ґv��kB�]R!�gw�r�c8fC�\6r���96eغZ�f��� �oS�U��x	��^w���,�9��.{� @q��DB�
 @'ܯX��{�c�2V�����
Je0��-�Ʈ��uB��D�(2.�0���3p+ue���l�sg��e?Wi,YdB^r�&;�I��J����`F�0�g0�ƕw8z$Ƙt���5�.i��[ɺ�(oK��b��FS(�U�y^�W�6#���w�xa��
�}0TM�4�_\r���b����0��|�hʯ�;O��Jy�q�dW��1��#4����ܜ�!U5h���,��8|n;����BpУc	��~�U��b���T9�v�Sf���27���j����Ap7�K�:�&��e�q[�Qa3�Z䷻�j���cs�5J�XH�}j���C4,>�%�x}�,Y���MJ���Gu ч��}����]��˟3sdn:J	{k��NНnj���0��f����9|�霞�IHVkm���L�V�kj	T��5�c�;N�5-�yŗ�^��¯)�!@w�8������;Z������;6�͗m�۔XW��L3zfa�lU�#��x\×�T��w��4��/���:�P���=,�ˎ}6͌y��;�=�-{h>������yV��f"��<������_�UuC���yQ��c��t6ePJrv���}ݡ�Ij/��{T���YJt��t��[V�ǣ�N��`�k;��.�2k�� �� @P�����rz�����HP'C�|�<����G|3i�ā�^���	\� �9t��j�_t�<���=�K�؈�
۵�Q����2�Yp���Ľ[�nlkm���3=P�o������':$TncyšA{:��>��r�:b��xtS<`~�BE���U<��Q��\�73��"��X�ڍPo��3l�|�㡻2���QJN�|ض똨s�,�&�т`��~t$[�*o�ն�n�5�X݅���;Rɨ(BSe�,R%?J�vzwC�i�b�~�UuVk������N.Y;��=�Ã�_W�4��<�Є�Vħ%B`��EP�Ȼ}l����� �d�፽\v�g`]�0�^�$>C����8_��BN��K"�<S���������S�7�)�K��s辴���q��r��"U�.��%��Qu��7��*���n�Lz7������A�-N��ޚP͍1�uz`&�ƅ2�Ĝ9uQN���cɛz�A�;�ʩ�=�-�`%��a��q0�'`>ȥ�B����Z9��(T���ӻbVk?�֜�k��S�3$c_�����~�F�:{�P���J�����Z���G�OJ6��&aj!0���;nΘ���ʁ��݀����u��=J��L�
��F���cQ�P�1p<�N�^6k���]�V�-�gy�k'��]��K�26��
@�iR~���w����t�&�p:��Ŏ�5Uo�쭁k�����ʎ�3����\�c�q�)��쌒1�U�8��a�����vs��hQO�bY�I���	�a\zV����ڸ�w,�C��?O�C���;4�0�����u�!����ux�4M�r�����4�J�U}�B�N��9��jY�����׷��CǢ��f�:�9D�0����R�گ&N�������E��x��$89yݻ9��ia�l�xA�w���!��")�\�we�zj@��p|N&$͗�/x�^�����T��v4_�e]�[gu7�EzQ-	���h�����~ǆ{�&%���l�{d���ޒr�,*0�6MM�1Sٚ��v�O\s@���y�hp��ٴ��.���U���������;�?��<"Vu)��5>�{����dN�1#�'�$v��ŧ�z��]"��u����v��K�{�vgB�z����5L���j+�7����d�,SI�WN��멩��ݺ�6k��;!�׻@m^��2pD�����.�Pɯ+��'<7Hı�����:���?J�v�7��͜�����G��MKx�4:��+T�ne����)
��v���u)Tt@�\�G�^Uz�A)�8��}.�d��z蘔��X
j��=�n���纸c*���.���]�+�Kl챂�y۳}��ܛ��Ȁ&>B!B�� "��m\��݅���������x��bx.͙0�)�A��<�:"S������z����c��>�d��=��-hi5�����ȸu]x��۞���|/��.�{
z�;���r�Y]�����"��S��t�5�U�9�b��|�>��c�A�=M�{����\�nu]s��ه�-<��i9	�^�E�匤�5��İ���!��n��\A�9O�j�h����<7k����ʹ��E��c�*;��N�� ��v��L6��K'cV��r�vPQ�cLK�;'�^��u^��M��4Ճ�R~k��y�+�_�rjNd]���z���!�n��!CA���C�y��/^�m|��BՄ��&�(�z��ѽt���M����W<�r�9w3�|��D��h�daaxLZ}���]��ޚ��.1��mi|�U���e^g��S��J�H=~I�Ǒ��.���N3��5�ȉ��_�t���Mj����A��CX�Π��xO��v�2�Zx�;� h�/��v;�!��Ә)D��Q-��|Ɲ+J(��mWQ�.���]!��}zL�8��9�}��M�<�;9��{ջ�zNL3JR��(�[ʮ��^�#�5[�6c{��u�Mdk,�^�t��Ԫ=�j�2`U:|��2������X���e��W�G�@@P�@�ܽ\׫�}��s?\Ŷu�oG�6�	��'��8�5{��i�Z��<����1?ncM��ׯj��l߳�����X����R1A��?_f�6���4�5�y+��Q�g+G��2�z7Z�X�����kӼ
H�<��=0���M�*)��K����0�	�\�h������5�H=e�M�M(yfֳюo[e���ոf�P.}b'�eLO;.�d�d.r%�����*�4���o"���w6�P�>UE�6�e�6�8��m:��x��ގ�dL+vS�itgm2^��M�[�hf&�!GId��	�{1���W*�qw���H�m
��ZޟP1� �Ns�A���8���Zy�cu��a�oR��=���K�+�b:l�6S�	�p�p;�����BG��{���P��ʇ��v�_T��|��n��0�NA������_E7m��3y:��nK�~u�m^a�NKا�~�2$��I�P�+��j��Uӵ����Wj����w��kM�K#F��wMR�AQ�!iĆ��:꧍6����l�2o���c��^9�AghTBW1���~�ߊ��ھ�έ��˖��{d��-�\[�WAZ1��2���]XA�E.��v�R��}cY�a��p����D
ѻ!)��c���D��e�%�ˠq��י�V��Y�[+����������{׀�;"�2��,:�9��*��U��C����䐬�Ǟ�ry5���d0�N�2e5<���y��������{*	{k��qGlM�o��<u]�t%g�~�%��U���#�����t�����	�k3��L5��9*����׳�K�uy*�-K�bz�3�D��iLt='nss]�3f]`��fBD[x�nna��U�.�#�(��1%����fA������p���|�[f`ZS[�);��hu����|};�U��͌���)�;l�j42��M��f��΁��G=5�,��3?���#�)f?ߊf���ա�_}E�������CD��Uq�M�<�0�^��W��M�[�E�����L��XXd�_�K�ʴ�&�Z���=�h���v�Po��-�g�v��2�,�o�Q���=skb��M�8&9�w6Y�rK�7����}n�'j[���D���&T~t���S�r��8�bX�'o��1\�BѦ�T,� �ħ�q�0_W�k���Bc��_�J`���[ʅ،��@y�8�ԧC�b���k�GV�H�g2*�lʔ��u�{s*j�OdճEEױ�xuwlz9>��(g'��Bj=ysxʼK"�����0�8sm`�}�Mbm�d��@+;�^��^e��]�-��RP��Z��L��q��̉j�t���f����e��gRd=�Etm�wW,���:�ɶ8,�6*��F��f�Xv�.��;jU�R{3��-ۺX�-�0�+ߦ�j��=�7���뫘�L�V�{� �s���:�uuK3
4��M����������p1љ�I�:��#����Vq�9e
¹�Ld���
�)"�{�ȶ��4���TVU�q�dr���nS�7�m��a
*N:ەӴ{��E�S�ú�a�mi-�K�𭾦v*�q�x�<I���EY�Dd�w}�i�`Yu/	s+�S�ޣ�J�� fc����7�) ���Xu�g��C$�&ܳ�j޷���Su�U�UZW̋aēo�\x=�Ky����#1d��1H���Μ�ћMPu7�D�<��.trX)t�p�PEUg���̜���~7Г�M�|pݷB��Y)�^�Ch�/@[��s�LQ��@�r�C�{�(׭n�d<�n7��m�9����y���	�bW��o_m[jRkܷ\.]m�s{�j�)�vR��^��V�Y�J&�ͧ��4�2(xFW���I��쮖��}��?�u�9H�:�ܡa��"|)��Bs�^,*m�b�t�������΀*�|v-��{��m�!�e�.���l�(�3�b5��wk���15��un��H$��7+H֡��A(�͜�Ia���bvk�i�\ܘ�V�ap�r��W��b�9+�@	'*�b�7wE�]v��u��+�xn���D�b�h>����odW륶{Z7��P��3m�J��˂}
�n�hY�y�*sw�i"��tZS�h_�SX����+#�l�r=؏�F�T�Y,dQc�Y��`R�!J�.Z2���Wgz3}����ۘd�`hS;ib�ǟL��a�CI�&��H��+^0C�O5��܊7w�v�s��i���2��K�o��)+���#l�4(�&� �h{�!�I@�&w��9|I��]�8���Ns��5�"�yp�e9�Ӯ!�ַu����WK`��qH,^e��]��z�-���6Ln�PݣZժ��WSDe:5�2���JH���7=����uO*�5Rv�J��3����v]<ԫ�-�x#�Cy�Q���Qꍩ��Q�w&l�Oin��x���`�Z��R��M������f�ηyɈe�);�.��И۬hiu����\�T��^Y髡�H֧;��kK��|�z���������D4Uuh*j~9�EPR�OV�hf�����9���~?>>>?������������&e��������4y�EUUT�IE�j���1�f�}�~>ߏ>>?_���ڊ���hh
.݉����TU%D�SDA�,��*�+��#�b�"�
(j��lbY�j��U�������
�j������QZERTT5F�DU$lb	�"���蚢���8��������b"(��_]`�H����Ph�
&
*�j
�(��&֡�&�*�� �H���:bH�*��LBLLQITRF�B�6qZ�AQ%4KKz�AMC5EQS��EDҔ�QT�4�TE^�=Au���j(���
"� "

��
��˳�Z�|S�E E?"�H6�i�I�A� 5��P4;x�{�e3���]Z�5S���_��tC�EV�-{>�]��z�"�q��j�;宀�aR�%�	D�H�4ۧN�ThQ�d
��T=E
EФf�-�4:_A#a`(P��LD|���ԓ�ͮP���4�3/3!���/	�>��[@.�|�&<�ƀD��^�oL��Ĳ.��X���QP���V�h�s��Rp����5��ۑ�sѦ��$M�Iw�y.�R./cP��[��!�}�����E2���9jw��M!��#�&�7H�4(�۷\V��Tܧ��.�j.श��j-?5�%�.��CP��e��Hb�䐴�Q�6qd�^�Y�{�3��:�V9@MJ`[��Uv��;���v�,�� �8~���aۆ��̇�������A�p�]C�tt��J�a\�V��Jq$�S�{m
�n�W���{jߓ}�,���(�^�ˆ������� 4ux�4M�O+'�z2U&6�S����u�sW˹��x�MѬ3.U�_!�_S1Cb�;-p�D�}�ߡ�_ߥ�|�hNHv�ܔ_��IuN����i�2�(cE��K��j�f��:h�Q�G���K&��!��ý �h|.Yxj�K��A�ƳY��S	���ڊ#���,!�?䳎�P�_E�����L�ŝ^>t�W�OVn1+��&���S���;��?X�?os�5�w�%�|�fp5�(���8e��sn��R�I�ځ��f���PZ2�����cF�zD�V���&XF�:Y���� ��#(�Gaf[��;��Qɳ�d�����_P����y��7Ƥ�K��V�Y���CZ3s��wݲ��B�E��~h���k�<̽N��<�C����wD"�.G�,Tϧ����K4�䩛l���lh	���8��1���!��ș+&��9=��^���4/B�##�Fg%�j+���%?1�{�a���Z ��T��2�u�V��m��0<0� ���FB�m�q\�Y�lb�qawt�*��|��%KTn�jB#��s�9zkw�HQ%ٲ�| ���W÷�Rc��oy��u�bt��oV��\�(�N�T�cIMmb7'���gG���J[lTpe}�`mw��~��g*E�+
d�L	ڹ���J�|1��n�G�n&,�>G�C�
A���34^'Z7w��m��6��K_Ji/xT�O��L����x�R	z�R:�3L8~�t��W� �UX��=`�L.H��@��xe�^��u[E��\�c��BԍcS�:kw�x��Sa}�n)�/�'B�{'>�v�����l�/b�h��pL����8�G,�����O͈�����𻙞���n�2[^�~�c��W�{���0�`�[ę���j�BBU;Yۺ��{G#�P�*��ΐ��9���]�(fPu��}�(+�s /�_ֳ)$�)�U:���?�Z%QWh��A��$}Y;k�6Q|�k��	�T7��(P���Ǟ&���/}�U ҋwf�������C��o�v������XuS� �Nw&Bu��\(��P�].��m��i	<����h�q�V�����l�5�^�C'��c�N��[E�����6w\��i�D�\	��_�9b��p6m?�Y�Y_�����]��&�ЯaN�/Lbhf�}|�2'�O;�^�}���� ������ŏ��(4�?D�/�~����C�������ٳ���&��'����A���i�ִ�-33p�!9���[�+�N}7����om��M\����Z��AŗA��+�ߪ 7��nշj"�X�¶u�6ǣ��Q0��wϩLH�*E���� �<܂leEc.r��q����m��|�4+F���]ўjc~&�Y��|jQp�3���Iq�5�v]tͳ, �TmE��U��p��yx'�,�^|�):���%2XKo��䇡^扇T.1�C��yA�{����S��5f��Ӆ�v�7	��-�]Y'�b%���J��RS�|�aò-�W�q�y���R]T� =�x���<�ǝur��þ8�b����f#����n��T3 O�!1[�=h��d�����w�,̙o��W3ݨ�Q�P}\�!�ko�'B�����g-�� �`j������!�k/wl�0:a^C3��}N����-/���@o���7�ڡ����7&�����v^���r�M�˴��T�`/1\�$�[�8���v��J�9W���z*0#�!Ƒ�~�	�G<��ΘP��2���O6T�"����̡�FoU�}��8�'�~g�m8Z��r��K�~��B��4�UfW<6N |��[	��VEm���Sw׈���&���(�"u4��j����9�Ɯ���6���fj�SWr�Ⱦa�鞽�e�@��1ak����*��>�{p�3����`��� �c�$DCf잋���C�d���N8��V��*	|k��H��+����`��#�ӱ}(�S�m��%��`���/��#wط�kP�J�M^�}a�v�5-�G�ay���O`��l�q;C0҄kv��:"w�~��d�P͗m�v�8ė�L3z�3����l�ջ��)�q��1$m�Lt�S�R~bfï)N�a^Ql�l����ސHse���25	gz�N��+�ڄ��i�lkâm�����(=�����^=��Ӷ�[b����,�~\C][�ڣ?Q��
���5?u;�N<<:�~� 9���bi+v8��9A���t_b���W�Gr���WP��E���Y���(MA�9�>��>7�q��wo�p�Y�&ؤ�U�Ӭ�j�b�/(I��u\U��+2�zG%�W��t�Jq� �9>���x�VZ��A+��F��.2�5��u]����Iň��.l���2[z��6�c��uc]U^��)@\�����Q�
j<��oN0�.vm�=z^0!	��kRm�u���n���`����#, Iv�n$	ږ-΄&��&T�P��+����Ƕ�xl"ܠ�W�'�̥�~�{���4R�p�HB��C_(����xNx1N%0L���:����<5UfF�a�f���A��%P��Ǿ�-����]S�y��_������*����"�4`vLA[j�a�KR�T�S�W8k����� �6LB`��n�|$J���3�� p\F��q�w݉����<��jK7��l�uچT`Ӗ�p���M(fƑ!7C�LU4g�Q��UĶuJ�I���C��]�PX���֢��ZPX��7'�����y�kVo7_H�gUkս�9��.�;r���|�&m�j�.��*T:���oԨw:���,"�<��y�Ae@�IN{��I"	jw����:6�q���?TĶ�����L�= ,}��.���T3df��{��d:ڝ�'v�t��'��!�
�ن`�y�piꎕ^"�wm�Hy�"F"`Z�r16�mf¶M�ոjk��i�N�cg�rCO���>� �|��,���&(R�t������t�2P���B���x�2�4�y��l��KsGX>*�AC����)Zd4M�O+'�{����O���Q��%�`@Õ�U*��_Z�od�o|�(����
l=��ڢ�%�>ȼ��nB/�Z����&��l�m�~�Us����zi�� ,�z+�tE1j�X�c=�,#C�p��焽�=�k9=�TeF��0wu(_W0�I�:	��Ӵ����b*�dK<!���υ
��2Θ7��Qj�-^ͅOi�sdc^Z�i��L:��PFL8y�i�Þmᵡ��R�MwFr�kB������jd(lk>>K�i���Qyѭ#9*fӦ�� +gX�$���ŧoKPm���j���6���̮^M@�u��m��yq��5X�-��f��o��t��kC&|)jI_m�˕�3��RaC��# ��U��(DA�.�P*��tB	��5#]�e�w0pf����O��O�bX�)Rk����9z1����A��Ivl��&r��5�fp���x=�s��+8��tD�%�DJuz�SH�kk7'���ɶ�Sc�^�y���ù!iड़���\rͫ	p2�	� \������ޟѿz��y7����2�ѿ*s8R����\�k��y�`V�|X��]7�q�ө�Zt7R�Q�n�r�u�ndb1�
�+ovrE!��gr��GI5�v��k��Ͼ^o0�D�I�9�l+�Y�H�%�HޣI>I��H�E�d���z�Ϛ-�=�؜|�x�F���}[��6���R|*��&�~OG�R	z�GP�o������F�L�Q��GwB(0�a�(�G8���mt߭�<'�s]�2��R5�=�GsʻѰ���k�56r�qK��"��D8�lzA1Hh��pL�����띒q�d�߄��:��|������g���*���-&�Fыwf��CA����]ٵ�|�7߬2#�C�F��/�K8=���X�5��WO�oƫ�A{�Q9����`�S����U��V%u�3��R���sSk�/v�ua��Nf�W����1\���,Z��`���S;b���!I�΋�Ub��1��8��ٴ^s�К�јzO�ۋ�z�v���O�𭉛�Ç#n��L:�߫��(��?De��?o�':Oy{����r2��t�V���fZ��rL6s��FE;ǰ(�
�|��镼M@����>[fnf �GT�Yy_~��r����D� :GJWkUzxc6�;��~��e�}��%�����+���'m���}��{W�T��A�N�����8H��~�N��\>	�W����,m�ˑ��48VkȭQX���^��	��7z��F���*������t��k{�0oyy��}j��ͩ��R/�����z�lk [:y��-�)^�	<�|Ǧ ��Ec4�^
��5�Fws^����DS�O>��,�,h�Z�_��eEÛp̂q[�%�C�;<�sNO3`��89h�Ѷ_-[{}.�B��r�ʇ�*�ʫ�g���nq�^�����x��މ��!Ьx���M��cR��.���$_Inj�'�)̀Q��!IN.�'n=4-u�qeriL��`�t6ãW7����_��}C)r���^�ҩ2�^b�s�"��+�
ӫ�ӽ:�'"&#�n8_%�JЗz�2�~�3G��jƔU�bYPƝ��IO|��TO4�Y�Ռ��'�����'j|d_#��Ȣ��8�A� C��0�1�t�|dIц�
�Z���ub�,�T����2�ە΁PO���268SH;��E��t��x�~J���z�u*��>�c�s#m�$��������"utّ��+ �>
��Ⱥư���Y��5��i�	��Ϭ�l2q�ҵ����U���b��y�*�?f�>�-^ �B�;HwM�����w��[�J`�p�H�LGo�=��3}��3�m�gT�$�<���*�49�<$�b��5��K���T.�5:P��8��89�z��ݛ����;wt��e�L���U`y�{o������c����~��3�}���a��b�%HM�8,�}�pq���<��܌�,g% �����	�&����R�^��l#ݼz��?HD7[�����<)��i*�Ɖ�Y���j��N��{M]�������W��۰���6�F���^]ぁ@�B�%�,����kS���ѷ݁{b6��x��{}uo��?K�q�v8��Z|U+;l�h�bF��B@}y���=3�sE��=��V3������ ,�pyk.K�W!
�y��-�P鋇�k�<X�a:N�M�k�h�L�F�ݒ"�z�g:��;}0�ˌ��A��@�Ru��Ű�y�:6)��b욑�r
��Ф!���)�8�u���N԰��%6r��+2#�a}�+Ǣ��[�#���ߑ�U��FŴ��Z�DD���}�T�^�BSV�q4�`W)�b���yw6��º8����ڳ�Oǖ`u^@t�\=K���B3[�_�Z�(�E�oD$�:v�%z,��2�����C_�ke:�1������c��'�p�X3C5��_�z��+D����6ȴ��l��h�LZ��(�U�������3��2O^�'C�F�*Λ���c�<r���+튝��|w�:�=�����s��	>Β���v{E��X�Ь3C�V��Y�t�s{�w)�Z�'{�7�諈�K�X2��v�oj8h~�o0$�a�&r�IwCTQr�ҩE�y�)�-�7Y��Y�7=�E��a�1��؁[N�C�L7=̷1c�dOY���=/�����?7 I��L!�ݱ�A�{�`ݬ���iŕ����ώ�S~YC�sBvKj�9B��Uz�X�C�����@��pN>wEgAσ.�sctm��C�P���`�\ؘ��^��L�Gu[
�V�NKԹW̋G"��]ju{����m:!T��A^Í,�mZe�k�c��Ӹ�Fg��[7��M�ؖ��z*��uzq׏Ai;R�F.�M�J��'�f��(꩎܇l��|5M32梜'�H���1�����ę���x�2�����:.-C��G���'p����ۈ������㷣�}�k�gP~�5�!�z D=D<z���-�#@�ja��΃�c��#D#R��-��ۃ�34*e���^��^mz/-S4���@���0aƋش��H�������N���tZ)"�]uB1��B����rj}<�/cW%L���S�W�Gh;�:�t�쑵�E�{�3%,*���dh���y��.�)�cU�v��I���hWJ&���<k���N�����S���ѩ`עVJc(L"s��;Z�O5ãy1Q�RI�%�P��F#-;���uw�Íe=��hRN��A$���]��T\J� �ð���PUj�_T���/hu�����P.�����^Jb�`ht�;��z9K2H�P�S�
V$���<�y��ހqXƟTIޚ{h+�6^3����384f ������g/�>�.V��S�Q�״n����v�u��ʝ�Z�v��e�}�)���ޠ3K�(�p�6��+��n�������ax�)R'��ET��i�nTM�a�h�[�+|"���\�����}~��yIvRx����(��A�	�c���7T��gM�K��4��
�g�v�vU�8붦r].�:���� �堼�\O:��f��)�Ff^N��Ht[��C��7e��5np_K	mc���:����{�S�eu���b٪�jh1�Czۺo{�.*�.�~3�u����f��`��(b�l�>��<����b���kE�2&�S|�0�������G��*��院ʠv����N���J�ʏF����4���Gm�TU:���o��Ti�ҒߏL w:@Xy��n�q� 6�jt�����_u..*�I���*	�^���Vʾ��'�NF �ל�z0�$�J�7�|��?��ʵ�n�A}Y��5i�]�%LZ��!���!���䀭��&T�����|��X�;y^�u�,/��]큸N��q8X6�]<d���{�b�'�^(�z�n]�u2p�
[\���0��v��Πp0��u�=�S�TV����[Y�6��]�����t�*�7VލU�>VI��/:լ����l2�����F���j�p1A�N#�Y�}OՅS��9�k-���VW|��K�*鮥��Wk�9#�)sE���ǈ��X��
��e��,:���6�pT8�ѻ��@WTPңZ�tΫ�(�BlU���t�|�	�v3����nk�W��m�6�[.VQJ�Y�Ü�6��z�#�\�s+Қ40,�\̑b�.���}�;�I��t��lfr��5?�����{�l0Гh�6ɬ�pQ`s�Yַ��3+��R���U�m�N�~�b��6����P0��D����2�B��-�a�0�����Jz�+��&�n�[�����1zK�m�A�w�[cw��,�g^�š���!w��l���l����%l7W�0��	˷L�#��X��A�G�E�(Jx�kgt��uem�<8��ñc6�N���,n�uɬ�!�2�S xtأ�DR³/*�J�2���8��P��W�Fv�vf)����rΫQv���+���x[ת����>HE@Tl�ES1��T�1DRPU5ES>߯o׏>>>>>?_��Ry�
��͊J�
"�UQ#TD�TQLF����������������������SE%QQ4U4Ɗ5�� ����<v��S�)��D'P��U1QE����lQKLT��CAIALH�P�Aa���:�EE%P�D�LBP5EDDM�N*iJ"�d�(��K@P4�a��=Z��
(()J���h)C��ZJ&���Z"F�JH�q�h(j�h�����+�z��u�(&(�bP��
J�h��R���
U�	AE
�|�]��}p�z�@�nم����-��n�w�&�06U��{�/�]�P��wv�a���dݴ�������/������m�5nE���^��zY���k��.=2�m�7��\D���)A�6I�cQs..g�Bl̹��`���7��6�Eǡ�P.l@�����l�@d��{���#�4LZ�m�XxS��x�Si{)�W�F�W�v>5{���ϩ�� �`@Y���ba0X��_T�,~�}+\_g&�k5�!^�'��$����ʑx$i5���$ȸu��`[q��m4[+f����^;��L�U��2���Q����(l	�3�5���/A�<���KLZ|�Sm/w]VDlE���<�>�ß��%=_)v�[�I�&y\������<�\�6��9����R�.u��n0�^���l)�j�C�H����M7X�T*��\�B̄�u_"�C�f�,޽�����*�\��cSH�-��<)�qHkNy��k��w\X���c��ƞ1>{�~�f�p��Z�a\�Tכ}�����N��ma$>�1t_'}��%��Is��Լj���]���B��#ʙN���]>�36dyWB���� ��ӄܕ��kw3��V�ƥ�"�5�q�v�z(�66����S�V�z� ��V��d�����+��F#����^�uww\�D���H)�
���TEJ�&gN��
.Kюg.���+juf;>���樆T��w�Ѓ"�'���]�2��y�?��bY��x;��­tz,MgJN���a^��;ha����~��\���S�?{q�����i��[�w-�nB`J��A���b�K�K�i	G;�O�r�r�reo3J޹�{�����ގ�;B�~ʋAD�gyjNtfϢ����ޖ��j*B�2-�i����4�,ݛ	�[��/6�l�g�d!��["�5���e�Hq�[N�C;��Zs^�1F�X�R����"L��ɦU�-�<�zw�a�y��zaB&�ę�;-G7U&:��s,PK�bt��%��k=�q>��M˛��
�"u��S��lm�\�)���l���^���]C,{�Й,R%r�,)���7K�<�3Ȓ����x�/�ܓ/3��f��������i��'�қ����=��NJR�����2dQP�V��}Ϊ�m�=�0R��$��5�bC��2��v��{�'zSz�,�&*��Q}I��ܘ�sw&z��|A��GaWT�Qv�ѵQG5ʁ2<1���%��j邞 ��x��R��uІ�Hڊ6��fum�.�+�4m��� ��I��N���4�w����R^]O����Q=E���+�q�~'o|�&����ͫT���5�a4��N���3��U�r���uwK���N�u�Xq�Ո����	*��U_ړ�moe�y-���#�X�PB��/9�7c�e�qsH���zs��~y�/}��=z]7M�GD�5]/s+���4]�i,
*u<5W(�����ơ�'S0
�}yp㡃�l�o?�{wy��{�Z�0��7l�r��qA��U�]<�n�k	=���z1�����+x��$�Ôٌ~/g�u&��N6*��E���Bչ��(���S���Ts	��\�^�͑W�@�X+��;���rǷ��{�`��̐1�"��̮r�&���~O�c���jw��K���e&��N���λ�-��}��W�d�4��
F�Q&請.Ӥ�3a�dv*L+�I{�I3t񈚫�]5K53M=�D���tg/#�]�����yOl+�Ql�{m;�=d!�d*ۖ���~�ڇ��%�.�Pz�0iz]���x���p�ag�E�n����!���酣]v��r�_^G���yʨi��!q�髦.u����:!"�ip�}��[g2ln�n�%�fk��	��-�]���s�aK�����-�C�?VpE7M���15��J�As=t)�{��ݷ���\K|���!%��T��k;�������]`��I�'�Fm��m#PP���r�)�Y�������JD�[���ˮ�&7�V3+�\�����&T�XOC��4��rVU�{��R�^" C����}5}'�a�t(@��;|�%ħ�Ѭ띩a6879�p��b�)�Wm��&T�ͽb���5��8m�t-��i흡�iĵ� ��|CW(��Є��r�N_���o[T#{KU�>r;ݼ���cem~����l���
bȇ���I�ݍ ���g����S��W���=O�'�d���)�x�I�>�s��{������a�����kԸd��=�����zS��@�ƻ�TRtÔ�.�tS�ޡ�r��k�w�A;0R��NK��6�To_s�k�M�L�ok�ř2��S�����pJ�a��'�;`>�aؿ%�Ď:�vq�3�JY4���z��ꧤ�-^�r��*��z�k*Gs�Y�z���M^��ѽ�ָt(�x ��2�`ʟ�	�lQ�%�Gu[
�V�����e�n�?��];"�{�1�-U$����,�r>�a@�4,�D����9o>��V:U����D��sq�mJ�^�d���k��Oa�����=1���Ї����vO�Ns��g=f�'�M�F��~4�,Xѫ��nCBn�H�3t�^�2�\`��M֋�,�"�h���ٸlK��K��0&-*�2�w�5I͝��.�s���yϞd�#�t�S���A[0�����!�7�<i����YY6-Vk�=0������o0��7[��#q�}��!��oN�O���V���_�(����H�ZS�Oߨ���=�� �n�����b��kw/f�}������H�dq�v�_E���a��&��6?;p��pݽ�6�-C/H��vM��Kս��Ì3W�@+(!H�M�Z}�tS���݊�Ѭ��P�e�����B�����V_�*f8�7rS�Te�3�+���,E����_=��^'
���%VQ�%^��S6��ʊ��"Sn5����+;Q�׌5��4�=^�ON���x�oV�^����ق�wb%�H�>f��E�!Mmt�j�;�&�hU��T�ڋk���Y���eȝ��Ơ9�<�ۼH09vkx	}]�vkSR<�ر�]�G	�'��C�$�D� YR�ނ@Mm~��c	�d\:���V�zj�S=x�'��&߸�;��2Ճ|�Hڎ��q;ԩ'.�A�EW3�����W9�Hz�STwe�n�<��@�#�M��O�͑)�9��ǆI���S)�g�H�`����p���&/F
k��t7�G�6�E~P^^��ܠ.<��6ŧE�Z��Ы2(��ii�eE��b+�K�4t�V�/�������9��9�Xe�8_d `RRuJiv�w���:�Z�]�ۗ\9��6,*�2���ܗz�������W7�e�t1a�a!t�"ˉDkH�!��C�-z�|����Λ�_��� .��^��Z����e;�j} 9g�Gc��>;��ݣ��QE1r��0֜�&D�׌I��-��9��U=v��ܭ�%8\_��}�s�~U�Iu�ӌ$��������v.��h�yqcWX�iz�O���a��\��_���c˞���(�l�|�>On�#z��X�*�-?o��`����S��XP����΀�n|��ChgJN
n�.��22��6oR��yt�|�I����Ğg�����h����N�;ī����~�Ξ�|E�24>:+��-|)�5]�ᱸ�H��u�|gɁ�
6r��E߃!��=3W�d�I���u�i�{�h�yz��r�c�y{��Y�\����&��v6�H��*;��j��}�~�hZ�f]W{&�f�Y�FC��+�3���Hj��i�L�ta�.+�Z�?~
���:����۟�%ϻ�^��)�}na���ג5��c����C��v�����N^��]s�-��iu�Fc��	��̋�S�.�+S�ϳ\��?o+��ŝ��|06
OB���3NRJ]q�o<�^��b]v���i��շO���yJA+
�V��0&w_��5�^Ψl"�9SI�i��f��VOc��F�P0��/���Rڃ ��
}���y����^��[�kt�ڔk��Ȭ!���~X�=tA���2VdI3:�Yx��5{�,��y�A[�����s=�e-9����.��u1��	�8H�����	�{�3I�[!
Jqi�T����7�D�U�w^>��S�&��Fq���3�x砠�9��r�CO�����6�p����g��2���?i����3=�_����#�	��H��i�I����!�x_v�+7i|g2�T�L��wfnF�_E7�m�xȭ�"��qXHM��!����*�h�q\��8����޿X����qܞa)d�yj�r��PX��P�3��@�
yt?[d�ٟ!nz7(���P�a	yN�x�5�2q��@IaKc[�R�a1���Ar� �wg�jM��=�e�F�B0/��&1�2)k�8�=+^�PK�B~a�hN���c��>��F-���O.7���C� �p�4k�¿(�ey�Xќ�i�k��t��[�}f=MV�+d����62ꁜ��g2�g�`<h�� x����<�C�N��:g�HF��^zr�z�kE�ltP���˱�tYDֻ�vo�B42�s��D327[�twm㟷[�I�x�\P3<u�^eU��:	!O��bW���Vgf�9z��<,#��/�N�ѹ�Y��f��63��/�Ҁ���-����e�����{�|�i3�8�v������S"N��<����x���S���F��tc[;	'O��ۚ���lkD�#�=`�z� 8"�	�OՑ����B2\]0�7��N�';k���}� �u=ȶ�1m7��<�_A碮B�F��q�黽1r�9��߻f�L��і��OPE�C�{���&�J�ږƠ��\��0�*.����͋a��%�$�2��6+�����+b��8��,l&�#�N�2Q�0o)��HL�b�I�iHd9�5w{M��ő�@S����Mـ����+�#J�������<��Bh�Za��]�oY��B�Pr{��#oK˧��3��V�Ncֽ����{[&D>`'�ƀESv����o%m�]nr�9y{�.S<2.F��%L9�+�S��'�p�3[�`��ٙm�����٩���;F-Q"A�jS���酎U(������u/������;�t�2��zu��gGuՈL��>��Lm����y�`<�^Å�/���Y?2NX��L?5'�Zw$q���Vf� t��f�vXxK:e��h����G�~+�,���Xm�t)[9�牌��P���bw�^�c6Á3ɬ([���Y�$\����<x��!��2��Hc�Fڕ"5Ҧ�����]�K:j�:.2Q��]�U��ê�U0 Q��5� �g3��,Ҽ�=��k\�	�lsm�YB�F\O�c���~���<?a5xQHg�i�W^ފ :����#�:�ꘖ�S�)�Gu[
yJ�^�]���=����M\dG]��r�.��F�K6VŰ}��3��n.�l~�X.�\���9�/��H�uf��8��(��`������Գ���gn�����I�[������}ju)�ף����3��(gHvٲޞO��]y��v^�:�c���B�(���
�F�2���M�6����S.��E�_���m��3�Cf���`0��O�"���^�]Sh�j�q����
Z$8v^Уa��z��z7�S�/'��k��Xu��#&c�\m�WP��}�lNxw�����|\(?|X'������QR{�Nbc�ς�1�rT�^97_'���]A�X�ƻ����bC:��Q4Z}ǀ��Փ(	������~X��PW�nZ�fO��!c;�n�qT�g��������,x.V�0'���z���u�v�����1Q�W��Q�~���[�ϿP0g� /70maxև��[��)[�3)�,:��ޭH漵ْ�3T4��$�[�֬�QԽ�uX^vZ���8���Dj� 9��b���qۉ�CC�����躾+]�]���(�5,��n�<x���b`�����ꫢ���MAD �P垚d_�m[,Ut*���Ʈ{gO"����$J���Y75Z^c)��{؞����`gעG	���~��)�{)͕"��F�[X�N׋����a��=�1��F�5�c�$lg=�!�2��v
E�󸑽F�r��k�W0�7 �n%�]��6,�
���y�t[p�C�	��86��/B�K�ۖI�Z~V�X�p�/F�85s�!��-#h.�a w@~�0�aAF����H��=|��w�O�z܃����}�9��89�F^ݐX��U��{	ZAǓH��҈�H]����a۬5N��7��U+�������[#z��Ҕ�U��/6�|�`f�;�g�;rX@!��e�f���F���e�bhz�B]1�YT,��ø1�e�|�}F#[��i�`��.�ʞ2�Б��n��S�����A��->�M������޺ԓ�i�i�M������[��,�O�j��Zn)h�D	ggC�&v� `G�![�p�<�f�{|�24q�.�8˷1��⠅�W�����H9p7u�m��9'ɛ�{�� Bɬ���������N�cEa���L9H��wBu_3�YOP�����"�֗H��i�U�'yى��������0|�8jc3U<�	:�!؆�v0��u3�!��ZOn㷏b�2���+�*3����������3m���eN\��22�{|�4g�G��M���è�uVV:R�8��p�kx�Y����r�]��{6�޴��w����9e�s�uk��#�t��6��S�,o ��	#���֒�<��ewX���t���i���8���˓�MR���!y�NIr�����B���=���=�0:�c��ܱ�t��x��|�I�(B���W0]�v{8�%�F��^"�_<�[�k1)��է�-S4u�S�0R�dcY�w��_c=X��'(;�؀��(U�Ę�ںN`r�:����m��x�%�;"0�yH+��9�2�kڮ̕�Z����/W�n%s�)9��K��i[V-�ض�����H�4�����M��M��,�C�M��Ϋ��1�#ጴt.����"$�D+<)k�M�v�h�w'2���*�;qJwȣ�����]�c�X�_b��p��lu��|���bf�ځDڡ�����y���l����s�pH����%�Ňm۾�qӌ�=Ƃ}��n��򎛹ѽ�Gh�vT�Aq�D)��FX���,�{� *�^��d�m���X ���ݮ��ng׍�7� R�ܕw�k�6�z�C�nݫ-<��3.�T*���0n�Dh���@�7!�$k�<��a혺��%����[������"�[|kk���噅��Ѐz�Z��ڇ��,��5����[?�^�vԤ��d{�7�׽#�e��N�=m�tWV��J��KuA��m(�h�+����N�O)	YX�+�Ë�"��m��C-��]iɰ�.P���rW4,�%��αE7Owot*�f�j-����YX��ov�V�u���ޘ#ʅj�]^V��;;YZ��o�`#@��ʊ6r%�{���L�S8���G�����Z��2>"��i��k��W[0�x�c�r��B����KF)9�r㸃����Q�)fdޠ�'�>�9��%�F�P�6�	Y�ۡcg��-8�:�����fM�9H�aY�nҥdk04��U�ſ1,�j��Wl$��7[��B՛�L�_ ���c8��E�9��sB�[�:���ޔ��|�: �,M��w�kޞ��e�^�*�m�>��rJ�H�7�(P�Ph�Ej�Y�����L�\��GK��L��,����;�S0;��`�T�ѽ��j�0�����h�[��es�o"YV*={�w4;���g+sX��ޥi�t����5�ֻf�/�R,���á�׺�l[%�Hb�9%�Q�MV��Z�NW��{6�دv�s�ŕg�a,�m]�X0�~�	R����CC��y�	AT)G�T�O�����������������)���o,KAI���JbA�J��hf)h'�����x�����������~�@�5GrK�ZZ�JZ�����h֚�)R���)
������d�����դJB��Q���:&��(h�������A1RW�T��4%&�((4�JJ(�(�&��A�-�H^��)�
�4EV�Q@�6����"
���s:h��]Dz��z�$)(ZJ��&)A�i�)���鴃AMU�=��F�)�>,�����x�Cc� ���a�V�����j�-U�n�_V5-(���+w���w�i�[��V^�s�}EP����bZ�Y*���)�fł�B��K��`�MSPA6ҡ��(�D�+d��1�"�<��9̧.����0SҸ�>�}_���,��q���]2W��F�eC֨���d;���j����)I�)��!��6#{gmD�"d ��;g��Z~h���l��J� =�ǟث��b-kn����|��ގ�*e�0x8�oA�A+��FCH��e�)�?4Ϣ('i[�������],��7���<d�쨬j���a��qw�%�|Μ�Ϛ��k�l��a�!c��s��E�R)�v���M^���C�e�tܠJe`-T+�0�9Qm����q$�~�ܓ��΀�f��.`n��Z�C�Л�z!2O~1��)PXe�'j)�q�ܧ@�)���aa��&��S�E��] �a�e m˱{�3zM&Ze@/�q��Z�������p�5�O"���!��_����	2�i�I���}YZ�ZѦ":qwu[��,���(e�U6]'�W�C�d�������i���{�CK�`;�~��$�b�]����t�ŌV�G��es�P�r�ߒ�Ƽ��0L��!��È��[�P��T�EL��Zv�<>N�<e9ȶ=�5R�8m�iz8tׅe�C�b�]棾�[��cWc�-0Wb	�}���&�U�h��ٹ��bQ�9�s*n�rl���\�w:�y�Ej��`�ȡ>}ƻ���[b�;R]*lvCV���y�;L���`�4�lGqj�e���SԼ����p�����­t��ʝa�������j�ˌ�GW��Le����cpеnd��ז����B~`�F;�̮�"9n�qX�0(e�{w� (,fp�AiS�3u�]s�3��X8��k�7_=�p�є�3v��k�jX�x�����+��J�aXZAJ���wV��.�˥绎�6B���Q)�3z�2$�b���t�)��,4>D+��˭�[z�����T�S��?vE>��Ti�@��h����A7�l8"�Y�����0&����˅���N�3ݸK��	ؼ{l׏c��$Z��z\�9�h��ۦ���xZ�v�M��6(~�0^E�o|�̷�}?e�ʎ]@��L]����/j[��!s�t��Jd�A�S��3wY�~�濅����1P��,�>ki��Y�??�����,'��Jl��Bd#h�hk��3��%s?Y$M9��	_�r��kxi���1l�C]�D���/�������t����/���P��E&�ޔ�+�qDo4kvs.���w���'�Ц��v`��ܩG7�=��R;�l�]��O8�u�'��޾ymԳ08�r��}�!�rԶ�Y;aZ;e�n����]��E�v_��i<6�W�o7�xbA��J"5]�����<�Ҕ�5EP�Ȼ|׶t�On�!ŲdC�8I�w_8�ݞp�Q�m�l��y�^ͪ�����G�d�q�x�}i��E������e�H���~�w��G��R�6������#����<�L4�r7�Ζ��^��Zøjx6�á�*���z���d��YP�f�F�Âۂ��R�(q�k�K�zO̓�r]&���xf�v��=j����vd5��s����cDk1>�.�jy�5մ.�J��Q�a��u�0�cFƽ�q��.],x�j�
��a�C�;0F8r��R�gCLO��Cl�X�{����դ
�Tc�v#B��%��)�]S�UR͕�`��5:��6�k�f�~������]��tDZ���Ӛ�qձ]=AS(��`r�M.���Oqpr@�	@X��V��Ur��WNMN���X�K<��ns��B71ܝ՝�q&E�b��Le'�E��@���᠛R������1´*`��q"%M��/��{6���X����?}F�{Y�{嵇�1�jm��?zΝ�~��Mx{y�>�뱑l]ݑbb(�T�v.w7I�8iû>Vrt`��w�W��U����\���V6�P���$"�7�����]{���V�u���[`q�n�:�1��m����Q�(��k���T#:������U�E{�k�See��ˉg�3�4,�v,��[ѱ�^�y}Lӽ�qYA	�P�z����+[*v��U��t=5�<j`ԣ֯��T��=_.E� �*i}��Þ�-�^X�ڣ ��v��5��0�C����q�H���f<����EG�TͰ�4es���W
@5��eQ��^C	�ҟЃ&*�K�ь�[��x�/V�3:
�xag$�;d�A5�]r���!׷L��g�B2�Pw9D�.��dB�B�.���5s�:y�̙tS����ۑMAz^�m	�a��D�_J��	�{"S�H�4����#rEއ��q��U4�A޻�z�]�j�y^���ڄ�i�Hۗ`�^�_�oZ��K1V�Q�cy�)s�=�W\�َ�Hŧl=��a��"mLpm�^Ȓ�|��{ �����I��lZ�6��ӝ�y�W�HM���=4�}��XE����i�#�H��Z���M�5��|��l�U�]�'���(��Ũ	�?ΛF��$�"oH7# �kO��l��~��o�d�aՍ�Pf��Kz�+Z!���U�[������鑮	�g �ǧYսVt�P{�ad�kH�"2�ڇ�.�٤�#\�������w��E����"�Z�e���4�������e�}}z�2�3'T�n��E4e�r'��� �� ��Q��d�O)gp�V�Nhvm�S�A��+����V�{�S�]^U@�2Wr*��n�ы���?0�h����#�6����O��t!�\��[+L�DĖ�,~[���ͺ��C守��ۖ=z��_��gr`�@p��!6��rĽz]��鑻�)86��L�A1\�Ԛ�J�7����+���R���je8�xF��)*~�)��HfJ��A����1%��ƴ	,[�m���d�⚚��N���c]��v�����sdK���4�	=Mi͌���jۖcv�|ұtC�m��(-���� �˥�A}kO@sͼ�̀���C�["�QIg/K5edŦގ����4���8�r���!�d4�M2����/@f�����Ku����6ɕ�D�.�Z���ͯd��r[^� �6�+�u�U�K�O#3%����$ق$�bd ��5�	�k�1w1
�.����3���Î����;E�44�Ĺ�����Hh�+V�IYxD�q3 �ѡؠ�K�A�����-=@��M
u�o�r�P��j,���6�V��WL�J��D���f��p0�da�q=9ƥLU��oSy5өS{��` ��U�9ZἝ�E(�0��D�.������v�s�� Z��ˬh�{%L��d�̻�u2'�:�0R/��"��0b!7�}'v:/�c(�?y�z��v�ۖ�y��w`f%�0A
=���2Ǒ�h~�ݽ�u�������.�W�����7�v�s�#d:FD?�n��6��t[���o�]�˝��R��J)�2�잞�c���-�l����3-�{jv��1ְ�8Fp��tdՒ����T�$�J���Cn63��C������Qm�i���Gu��8���T7�+]���{\u����|��5��C�(�0+��m�D99>=�+�u+��C޻;��B{ج]P3��4�����6�0OoC�LP��� �9#�w3�TVB�V�o�;q���l�,4�$H��{06�����0n�3�"�����7w�� ���ztۙ��E��v�C��_2wd�;6"�\M{6���oy����D�惂�k���2�:�D�#T~�g�J�'_���b��N<�JT���
�vE�U}\���|9���l�!v�Ԣìm-
u��BYr�Ϩ��؞V4�U����@^�O\�*<�ai�ىWf�KA˦ܫ�e�z���w��T�2*^vm����2�� `�� �H��*�||��;H��|r�}Sחw����DH�;>�DN�M7���k����<����[r����P�}F���r���PR��O69oV��Vɹ�c�ٓIe[��A~����FDa
��Yb�&��^�P��9[j��4�h��SNf��WG&��H��B��gb�a��u5���f�8�/*�)bd�l���P&��u�Dd��p�.���/����}x�w)ޒ�gG�Oq�'I��ykf���w��kgHa\���tN�͙N�<Hn�y��݂������s)i���j~��?ן��_�1��r��U���8ɇ4�T��$L�E[�E�sM���m���@�M)���R� �?�r�;�s��x�c�u�n=���?��3���z)!�{����9�7�-u��#ec5�O��~M�ٵw�����mvyGg^������+Z���� :ך�DWPu�Meow�ˤ8e�s�(��ܭxZ����[jھ��/�qt���NW�,�e�E��q!#:K��H��ڔ��䖵Z�p��B��	5f�s�I�+���0�${��n�w�Ux���{k�Q^T�3"��I�|7�qm�#Kv��=��j2��h�����=,uej3��=^�� {�5G��G5rQ؟f%_EWuXyj�P6�>H�G��K�[y�4s���:�	��K
j�7��{[N���gy��@+�L��x$��۝�;�"|H1�Z��sh�����E>��g����?$�<U߬�k��~ g{�|��*�~�#//0X����=�d9K1Ь�חW����S�"��e�����~��^�(����'
�^���q�smH�e,��d�E�"���K���ػ�r�2���R���3��f�۝!�cwq��-<Ĝ�ӸZ�GvﺲOH�Av�)OL���N�Mc^���mvl��9�`s�s��jZ3�=eb���P⨤T�D����9��5�e��/;ݹ�
���J���\m��n��/�徺~߳���-]2�N#�S��	�c����t�/)�M�wJe�t�39�u�!�K��ʽ�Ca ��\�3��ڐ�X\��m���ir^_8��.����L���\C�]���1�Y��EW�oG���wі�%@��~
Sj�^�oBKG:�w?}��Q�ed�f[~^ɷN-��{��l�f<xm��Ӑ��������M���:�]�S=>���v�������T�7Cp[r7��p�R�ml�ەyۍ9�V����'^}\���]һ�q���`�:��~羐]WvV��։�&I��E�T緒�Kw���U��z�7x�r�w�Ͷ�Y�z�ڧ/�؎�j�3�۬2���S�-��=�; ����h�iS��H(�V�>��N���Zr�.��*�7h0���eɦ��f�U�a�Pe���u]@T�䕹p���|�7��m������R1��ߥhE�c!�/���M�e�ջe�y�[��J����V��~�����Z=�mP�:*��Q�*xa��j氎~7S������K���u���qz�H��`��~UٽX��_#L_@T�q��;��㛒��2����Vv=}�\[�1I72ri6�0C�����-^�u�VNt������eE��	�G%.���gYYl�j|P�I��@$	�NW�wg�� �]��g��Y�u__��	]��g��N�u=,�k�[�(ތ-y�=#��fd��*8U��r[@�	�R:���cV�K���wҵC�����'�~��p�~�%g��L��y�W\��fK�#(M��I���4�l)^�藡4�]
Ȅ�o�gԛ��R�pW%/���d�[8�zd��X�bԍ�u٘$[�$�[o��.�!\���h-��
��_gl0'��t��y%q���R�o15���ǽ֧�ZKUdm�lg2��a������-�J��W��S��==,1�N3�a��P0GI����UaIO��zq������R�����R3lz7�s��/�J�n��a���D%>�&E�����U���c=;���F�2ܵ���䉖�:c��ߘ#��w*NO�j���=1���Ӻ���
W[�!賲+���9������"^�F����^:�'����c�X�5�b�۾.�Tԩ�%9CK��P+��H)me�5���O�'�&1�F�p�jp�̜ڷӬF4�nV�V\�؏͏��إ/J'Q�Y2o^�{V�J`�i�{(�7Jk�D��W�������s�m�J7�^=�6��E�Pͼ]f��3��3�)�6	�خ�������Bf��WܵX��ڬv�b�/&N�-c�����&�-��J�I��*��F��$��}��';v�L)�z����^P�O,mD������TV2���&��p�M���*iޤf�.'�9�]����OKd��8�35���aXn��ѡ�X�WfΚ���I@�p���x�k�y��\̬�׀=N��^�1W*��8��4Pu|[Z�gu{�,�����8ژ�2e��Ტ�J[�uЗ�#b����_v����h��l�lp�*9;�դ������L�X3���٢�C�M���we�}��2w'{�KL�au@es[�)�NI�N�&g2�����Y�������4�VG[�4�ڒ�cp�*�#���K��Rm=/��n�Kase�?H�SrзuƸ �T�~IU����u:�֊���^��/&�]Է����q<�Y��vX�Z�T�Џ�\�����c���̨��C�s���5�ԍ�f.��GΑ��*��V��b)�:��a�'����@�s���o9��f��KѰ��]v�e�I0�~�m����������Gl��X(����k�5"���	\xX�Ԫ��v��\.��V�=��T����EO����sL\2�i���ѬAVZю�VՂ2�-�)ϔ���Ǉ��*�67�Cк�h�]jJ�yD�ݠ[o����s��QE�
�:�g�"+E�ed�^��
fV��<�+E�R�d��iSw�jٷ�֩�!	`��A�v��4:�s�g{%㠔s�s\�E�|k��hh唷.Z�,��k$+��3����)bε��\.ë�����o$����':��*[v���}u�8������H�N�T�o�� �&,���t��:��Z�(��H������귖��z7�t(�磕��y���C3/M�Æ���ֳk�n��>�7�.��V���䯎Qݥ����<��`�
p�6{X��s�7Z���[))��Pz�y�.���s�v���Y��R��ϠT�p""r�[���:aw��f<�i��ƕ�%����~IVR���0�B���m�u�Jv�=���k6���o���e���n�IK+��.w](�^�l��p�LT2��sy�.�C&�2�F��2��]��JB	��ef�ƺs)p��~�Z�p���5�f�@֙�����0Y|	�[��;��������D��RЉM!AM)��%	K�Hғ����x��������������_��D4	M4R��4�4QJ�r1�z~��<x������|||~�_��f"JF�(�bJ���|�"K�t�WVJz��B�����*�70���q�8������*��+��_r���hiR����h�h
���JZP=m����4�R��4�P*���444i�T҇�����Д	Ԇ$iB�O��(:� �RJ�	C�a|�^��P4�uh
[�� �)S���V{����ђ�_��n�/N	�Ī�s��՛�4Gu��"2���q�4���i����{�Ss7x��[��6y����37�k&�P]U�ܸ��L�9Î.�+E�
�
#{/���}�L.6-�{8�]u��q�n�����Vt�c �>c�}%�2�.(�}eb�\��S�]��ߧ�IO��Oi�9�΁��YPZ&G*9R����t/D�����h�m����� "H�͞8+l���o�8'�.�p��1�g]w��J�Е���uכ�xH��q��DN�L(����a}+&Z�7_
�^��Nr�J�8�|�9kb��Z�P8���lDT�.�p���Нȝ�cyj�]^�8C=p,#z�[�p��ɐ�"�����ܝ���'��E������;W*��ճ�k"؟X~����Jn����ּ� j��8��UA��e�KX�ֆ�z�,XLMUYw��=�m��R7�%~/�)�<W>�W�=۫�;�4���~�Ç#�*��2)���EJ&�i����z-�����T�x�1t%é)�-�o-�x
��HW(�(����^ң�I7�V�WPR+�6�!++7&����oyl�:�)=��+zƤ����o��w"{�����d���@�^�����ࢸ�f�%c�"���Eot���/��U7=={���q0Y7CTz!��.��ˤg�)�[d�B��4��+�P���o��ϼ�$��}�����WC��6<�T��ug-�a���qE�+S)�?u�Er93G���k�)�e����î<�oH��!�7f&�qoJ���Y��!�iRIk{��	ɘ����e'��S�#��`�q�=��oz��l=$ #ʹ�n�b�*/x�x�g��n�-j��Xb�r�-uXׂ
g���%�ϯ��z�~��m�ލ�vǚ�R���<�M{
ъ��w h (�a�Y�E�xٗ�� o	��+�7�Ow�{g;ȴ�c1��'��n
\���w
�邥B*��늺�̅o�������S�d Ix�e)ا3�qc�U"����Zx�y�$U��Щk�.�}���u�G�z=�<����)ж�4t7�Y�fWqx Ĵ�ְn�h_q��Pr��Z�/�_Ks����cm�u��Y�^Pw��ƩW{��m��y90�i�Ku��g�۬�5��Z���gq72��������f���o�3ڙ���4<�7���-�6@&Ѥ�ߞ���%�����:��0�ӏwwp��ճ���u�Jˌ�W1��6׹ �+��;���ˉst*"�{���0��.H�$�ݪ�n�i�9�(�75�r��_g>�;?g������u����:+/G�]>�H�<�q@Q�
f�p��צy{\rcKwG�ݮ����k��7rڸ^�F���j�� g�otWbw�C�n�3�j�h��Ѷ�!p��4
��hL�-$݇��&��3�����i*o.V-��[$v�����Am#z0}d��uU`շ#*�z��Y���o\�x� Wt�ǂ��mq���6J�Tl���p��[9�.�>���_���_�A�7��-ރ)%뽯u�����W_U�W3|��m�w�rH.`��ۏ
�J��ǩ���]��}���o�*��.�!�s52��,c�<�bc3.�J�gF����ի[��5,4p]�m��q:�뺥ݮ#���S˜�`R4/4T�R����t�M@b��I��*���Ž��,a��H�ۀZ^�˴u9�:�s@m���%v۟~�������\�{��W�Pm�r��'����=Zr�.-�� �[�&��`V���v�/M/a���d1�m�gU��+�������;φF՜�ܗWs��`���O6g�L`d3����qzN�^�m����ݗ�&�^_F��J"=�Z9m�zpsE��h�.f)�1��nc0���[Q5uW��˼���A��E{�^p�f��N����L�l;s����v�%`;U*�M��dŮK7��j
]����-��e��u���2�X�1���g�b~��Ѩ���B�����EV�ݽ��8u\ğGj��y�Oi�=AA�d$0_w���ȥA����m�z��Ӫ��^8�I)sƩ���r=p�ݗ-�B��BV�!�#����Tu�B�`o'��?Ȯh:W�����10��{�ʳ���;�����׽���ᴱcz��}�|/��@�7u`�ʳ������N<�`����}]�ZFߍQ�ab<X��e�|��,k�F�؃���fE�KzԺɯZ����RۄU�J�;�Co_2�U�_0���^��"��y��*rT�z��WIU�W�j2��gǧ�0mSrwc";�vl���;��	�������z�|�U��4�K�N󩹰��N�/Q9��1Df����0[��v����IUL�=uCyt���q��	��<�]5`���a��q��K�P�v�8C7�,��Y�iS��j�6V��Ɗ��]<��]A̓J ��[`m����ƽe���Q��5������d+����6��n䣛��)9��r��NǇb�h1���9gSO6FR��+Ȍ�z*�q����0I�=��?G�=\]f���H���Pn��qV�ҔU�Y��/-�7�"H�<������vyB��^DI�ǎ��lw.%z�>��{Jc��߳v��ʈ�z���yf.#[;4�Ec�	��>1O�%�P�k����Q[(Q��}��(;7��W��f�y��@������8��)�7���L��̜��)���]�hZ�L���V�cS����꬧rޡ��ы�%�w
��k_"r흮�
�ߡ(�M�5Ҷ����1��]�T�f��<��y���R��6������S��,_>4�'V�cH�����:�-���Z��a��q�#�T}y?T[�g[�~��)��I?�b�J{'�j�'}�׌�G��d�����N�W��%iz����OO9
F�]C�J�YWo��u�g�ڱ�_5��E2欽�rtX\���q��@��;Ғ���b���p}���lTXB�u9����Ι��w�)��~���N�(ţ6y.R�y&�0�G,|W��wO�1J7��������ݹų�Ⱥ@�e^[��.g�߮w�b<���pF��:'��3��W�!qw�J5�����cp��̚�wHBtL�tk�v�Vy�f{;z1;�4s�G���0~�p��0އx�Cuž5&�󲸹�Ⱦ1���io�
 ��6����g���9wP��隅9��A��g)6⳨���ث=�NW�� t��r���m��55��{����䊩���p0�U���Ƣuۅ���I����p�@�y�H��Q�d%;��CM���q�R6��
�tG�����#i�>��ԏ4��c�b���e����Nl0�kT�y�J�D����j�FŎ�D*�[��Sr6�����uW���ek�ּ��廱�gްn�=5U�?#��a�Ԉ�/�_�l��ߧw�[{4+wӰOЛz��U^��޳��#���
�z-)���7��!����ó�j;��S]� ��h�>U�o��D;�+���*W&��,�S��6�U�]`�f�J��{iQX���z�W�Ng%�1�tϐO�Jm�Ku��j6��ݰ�t���HgD�,��	�Cg��5䎴�ڐӺ}�z�)��)�@P��*��F,���� NM��ɝ�P��PR�;�Z;W޹�2Ԛ�i�[�}�D�i�8i��Юjڰ\-�5�*�9J4
�*W�&Y���%��<�"�~��c�����?�~N1tUk�����G��k$w�[�̊f؎���Ff��=�����V:���c�p�A��i��(H��.�q1&�V�>+���_���=�Wp&���6��!p�-~}�%�'EZ�q{�b2���41'�������g_Fܣ@�X�oO�v'L���$�_*�x�[ɵb�}��U����j�� M&Q������g�u뀺���|�p&94��ܰip�����b���І4��i�l��V���nf��;�k��_��RO��T�����d���T�h1�:�ۡuT���Y�G��k鈘w���-�o���A26zz�s2+���\��w.��]�m��.��;KZ��r�}֓톻��Z��#ƪ�~��O�n�P4�Ue���q-igC[�h`c��h�wC�踍��a��Ǹմ*�uȾ����6�$�4:��HR:�v�E���.��E�����Ǥh[^R����S�W/1#̵'�ödu1�?�
s��8`l����f{�q1�dm4e/y�is�A3�����D�}�y��k���3��<2��{ڡڡ�mE-�A�xF�ȫ=��< #�gr��?f����ܹ�xǼ�OGI1{�4"jꀼÄ��|GJTD��@����7�<�y���uء�C!��j��S�k��1r�-3��w잺^�W�V-z�˯�
Us�z�ӥ���Z�[x"�3{b���,�B�t��N�U���_;��x�E��P[갅��0c�����{�+b�C/���P�yO1`g���뽲Z�Aɬ�^]��f�w�r�Y���O�"[e�o����	��3��w�K2���D��bh����-��O��~G ����f^�)eM�Ǖ5ۤ�������w2zh�4΁�Pna![�ᐺw.���JU��p�����t��xD�����[��{$_zR�iF��PÁ�sm�+��5�EwFlq<��<�q�'e���v�}7%�h�O;EEB��0���>� m�U|Z+��eq��eo>����U4��Q�&j�D���Нs�>x��!t
�=^�H
�esϩR4�v7�Q���M�s*��L%�,l���a��z�AR#��g��yrUU�lX��r��Vĭ޼��9�G^ǺX>����`WHؤnS\3	DS1h�5�7��蓙�5�����韞ӛ}{���g��b����g�=ZԸv^�oq����%�~��5FOv�a�h1�8��o0B�k��O�L��ޱ:>Kv�7�0�H]�4��'���LR��,��`u���+)�zZ��W+�a���L�&W��E�XDt�M'&p�δ�N���sy͋�<������W:,���S�h\�C��FuP�d7���2g{����|�(���k�8��ۊč2d:��b`��NY&KY(h�|�Vn�v>�\��m�m��|��� �q�*{#��)<�d<MO�����Ǘ���pQY���g^�֌NL��+7���R��gf~��g�WT����M#�:�[��g�Lqf	�d0̣q1���Q�K���n�f#k�͖ r���PWE.��^Z�����As�X7��B縋�i8������cc��iIPX�(����K��[g�.)��ӍUS�ԟ6�vN��pʼ샮;�|zy�R5B�JT!T�w#i�m�õ�xt�7zKa�clq#��"s��.�,��hb��<Uj�=LA���G296[�	���$䶽<7�^�@�-��r�V�Mzq��b]����F���]}!�h�����յ{�l��
v��M�L7�v�c��U)Уښ�ˡ�ihqn����c�B��·�v��WC}���V�.F�G�,��3����N��_�s'WKJGLu��v��s� ���-�溒��Q����`���J�kV�^�)+��^Sw|�ʳWJ���m^Pv���f��wZзA�j�b�p��(rR��HݺW����n�Anm�Gz$��h섊 )Q�V��6�f1{�՜S2^�LQӺ�,�I�D��3OiZ�:�Ӽ��n���5)|C<�r8ުW��ҏeZiL����i�42ȇ��ђnY ]�Ԛô�wX�Q�ԣ����[���.� 8�������3,>�uk�/Q9g6s�Ɨy�V��(U�;�ת�����I-����灀�b9�T���[y�-�R裳2��se1ئ���m)+yY�K������g������[�D��]n�>���F����^�q�^�Y���L�[F�Y����jŬ���S����b�t5\��O��7��U�ȘVJ�5��Ue�>�E�A�CgPn���z��M�8�-bfTʮ��bH�@�OL�V(\���B��y�o3t��q�:����U)剷�Hd �h���Z����}|�u ,N���v�Ū t&���%x�ph
�ˮH��5���pDs�ءж[���#Mfej)S���i�9��|C�
�����9�r��A������4H�O~��>RmY��~S�X)����}�5Rڭ���[��o颱�b��2��^N�����%c[�n�Z�&�Ck���"��h,��.=]h�'���ӷ��RIeeI�|;H�N�N���9ӧYD�}��զ
˷�3G�0>f��I��u�V����7���!t��K��
5�-�ǭj�d��X��kAt���`��l�B�|�NV�(uwf��R9�-����v�f=��/�ݬ�?+&�@����*���۹z (���@�q�R�޲C� u��!���=v�I�������oQ<�����^%}���"��$�!P���洳u�桺�WR�W.٭΂�9:
}���t%cc��$i:�c��u��k��v�[����8�]]3E[[��Bh����oH!R�S�h</V�l�K@硡uf܅Gz�h޾F���j�m���`�X�IY�jιH�	\�7���*��]�����'��{b�Jc{���',Q}-�oeG�2&�+}��\���c�u�n�u�<6e�mR��7[�ϵ�V�+!�ܟN��[�K�k�+w����u9�*=�[�Z���Vd��src��Z�F���em�G���m�2Z�ַ�a|���y�d���g/7��T˱��9H.������$�੟M̩�<��Н���V�U; ���5�?��J4)B�M#C��:�)
�����|x�}�<{{{{{7�����~����(|��@�1JQ�1-*x��A��������������������~�����
k��4!LAB�䁠)(Jj���Д�R����8��eБP���:A:�Ҕ'�t4z�1{���O[�5H��{�-P��SHA�P�	F���u&���Q��
R��4���t!�C���(��o�M*P>�q	KA-%�tTA�"i�{cH+�R�PS�i4�HQJ|�*{�5����=�S�P�>��B��RR��}��u�kz:=u@d�H2�4�+9����.�)=lC7.��Z�Thb߄�8`i���Vu��J3fN�qS&�{����p�|V��
i@@~@
��m'e ��W��XD6����^Kހ�ZW������^M�n��O2"*�w���
5e"I\_�#1����זW��ó�OS^ve�퉕`�tn�Nw5n뢷{o�i"��Z^Jݐ��i�cJ��zi�O�B��}Ւ�ۣ|m߸���}�[�gMB������(5���D������V�fS�lY/`8=	�e�gR���Cv+Ң��x�co�r�V*]�N=`k"S8�Y�Fl�u��^�ź3y�'��H�U-��C�Y�~����A���������/CY�"��/�3
y��>��(�я������c��݂U�b=Q�CL!_6��G����s�����$/�ğ�bY�$�(�����S�s9-c�@A_�KV`M�f�xD�@�ׄ�<���hn�h�H�H͵r���e�&�O�Yܻ��7?n���3 =�ʛ*��d�!mPJ�9��A�����ImN7O655�P��LC�H�(uc2��{�Wj+�O-M�vH)7�+�Zf�7c�}W���pA�� y2�N�����Y� v��R��d�7���̋!�Te0�&���/�*�]��2���������o8�rY�:v�sl��7����ַ���&W�hʠ��&�ڦ�l�Ur�JQ�Uj��U	vvl����vl)ܫ�j�2*��'9��U��f~��A��!U-)w8�Iu�k�"�~��*�EO>�uө���ä#��~]o�A�������s]�o������㫉�����!p�-�wD3KB�?���f��F�Ƨ�I��W����(�r��~e���rw7C2���_��eoh���״���==|�Erך��˱�L4=N�Bn�e�U��=o�����0]�3ȩ�GT�-�S��M-z(�ʤ���-����3z��#�ꈪ`} ��p��F�z�ݮ~$���-}6�w1&g*�)����HF��FH���m��S��@Y��!r���2�߁q��ֈ��g�&�����L�]J}�@�g9��0 ����ѥ"�r�-l��r����7|j	��� %ӣ�"�  8n�Yup��5�E�O��81`�x�M���W-��t�OwZ�9|���H�ek/K�*ˬ"���k6��ɴ�5�Q�c�zykE�%Æ�M_94o^�]���x��tW<X%X�g0mYc���c��ͦ@'��3���@��=�ۆ�K�;�N����p<<q���a�]�f4�Q4�G�-�]��Ƶ�w3;�{AqQMw���kK0m���U�)Q� �/�:��W���1�k�+~�k(U<�g��r[|Aȗ���s�]�pӌs_�ոWKsI7^��XY�����J�;��Y���J�k6ߺ��=|&�3O��5�:��ft��� y9��~ǻ�������M�9�*�.�E�+|��ƨ�S��u=�E�j�4���a#ZDζ���G,�������>LW7zO{и����No��AS�����n�Ø`��;��v�.��h�t�Zeq�ڌ����!���WN�*���}�7���K�]���!t
�=W�UY\�J�>X"���{�$�C��BU�#+��V��q��ť"��!���I�\;"lu�/c�QJ�}+Q�<�g���W�,bb��2��.��7iյ��T�޷�n7]ԝ(�*�CE枓r���fBnU�R�I+��ͦ�<'�M�AQ�`��x,W)_�s)�^-������an�d>��*Dq ȳ�Y��&9�b5��6p���=	v�^St��+��`�m��3`0���Dv+F%�^M��r߲��72+��6����$Ұ'�<�F�S��|�F{�0�%���,�1��ۙ������+�9#I�&�Td�l�f���=��\�Qt�_�؎����ά����.s6c{�9 q�� ���f�F)�}㭷f����N�4'_C£QV����{����f�0ԟ��E�kO0��\Vk�s�.-�ͦR�j@������ɵ���ćzm�}v�T�;f�����;O�y��"F�&�^ڞ�x�g;��=ܚ1ɋ\v*�Wv��il�1ٜu�]��[	@WE.��l���-~����VLy�e�Y��{�@7�܄d�+�)BX�r����y74�V���Q�
FLf6����6�s]�r�&�v�z�<��}p�`���eRL("b_�0��]����T���
��m���(�:�:f����s���������Yz�+�y1fΰ3T"��9��=�#�ō�`�ި���ں���~����B7�Ǣ�����il4����
է���q�\�ʟϗt�F1�"S;3B��};۬��@W�Lu]��V�ބ��F�)�t]Ý{7�(sM����F���5ӝ��:+c��:�o�����7��x�z��\�)Z������zGf��_H�c�O��,�F���3��םZ��6*+p<W*�E���>��`�eq~�f<u�Wye��)����YEL�b�l����1G��{���Y�#��-t�`㱝�F�T.黬���ާ�!'S���&eK��o%�wL 9�������ֹ�c�U�6��y����p�L��gRn[�دJ��Ǵ��Ѓ����M�:��.�a)�p.�|��3\V���x�L�+g��6,�発[�o�HE��Pg�us��x[u���p�T��m����|v�=^jF86�i�es# l�I!��������)3�h���Pe�J�+o��������I�7�вȭ;��fV�N��|U����ˎ�$`0Y�/�s�����c��|���[����\�]%����]�u\��·A�������K��_��-�^�d�7��K�(O gO7`�â�dd3�Ю�H�-����M �{3���x��͓|⮶3J��X��^�U��s d���E�%�!1fMI��6:��S�/1O��'�<��h��Zٴ�]0�v��4�s�w	}�b$*�����Sӄб,# ׾E*�q�'��4�1J�K:�O|%���>Ϩ1P(B�<b녧��P�(�͏�`^+��M��LI;'&�j�3V� Nj|!�]Jό�?�6�ͮ��q09�i
�G<wW�o*)<��ucs���!F�6<[��׫��Dūa�^2(7�9��I[r�^m���=ʡ��-���2�f��*aؙ�F�x�Ù��Adl��F�-�49Z�a������*G����O���R�,��۰Fl��0,ǜ�S�vzz�F�-y�H���c��a�z�Ö��2��jԎ�Aw����r�*4�.���@]
���K �q��fZ��#B;��vj��:�|�tK���>,;KZ,;	��"�b�t�����7��.����p�F�+�����ـ*�B��}F�O����[�$��@�K����|��[W���/��ds��]���cpEF�Y��%�S-3�Sx8��(oC����n����ǩ�v]��5�ї�eKuoGgh켭�� _�ss!pF��o�@X5��^��'�*:�nO��[ah�ݲLt��zCv����.�#bZ�?i{���4Ȍ�Yܼ3[b�΂��0�z���~U��j��~���l�X�-O�Y][�j;B�!�]�Һ���Fo:��o
#N��[h>,e�W�s%Y�}��˧�A�l/J�hעj�2�GU�����5���i��v�"��݀wg����:S�T,R���7<Y�1r�-"������z��<9�t+��Ư���TK��A]z�g��~��T7;!�Λ4/#��v��6��I�fMA�4��d���5yР�C�WQT�򌵸W�q>X��
�^=Wzת,>��k�8�N��<"��7.�c�� ����������oX\�t�0�|�pڗ�pC�ʭ=����?:�������I}����Q�WoGu���N:c��*��l���߾���o_�t�!�̷xG���k�J�^���<j��庮̊�0���MD���g�C3�K��0l��Eo@͂��t�惠�2�:�ӭ1m��v�S�=��'���6�$-��G���#oۆU�`6�J��W��|K�O����Hľ�O������m �K�
��3t/�����[c�����x���]���^l��d�R�q��/�����ޯD"8���3�VU�SQݹ�Ɠ3��ѧ��Z�/+v|�`t�q�����vp��zu;��u��I1�}öru�2Һ��i�ӫ8�J"S��i���L��өd�n���������2siF%���3|��.^O�^��{Toge��l1|[�#�pL�����a����pAP:��(mq���&|H9>�#m��Z�eCY7�Niavm[�;PB�`h�xUo6����nl���T/3ŊǶ���=P'L��{^Z�����{D�G���e�I!�aM�Uu��Rv4@��7`��nx�����3\�9c%c��c���YL�kNŖ�^#�[L�Aij�D�\!�ٜ���o �%����.��������8>`����zϘ�m��|4�g�R��|��v�U�V<��<�� ��0���ܜ�n嶡֫e�k��fƌ�V��wL�'O&�{jG�)�D���~� ��Qu�"�8��Q���>���O�X�+�)v4����ӝ��!QH�<[2N�#wN��O�n�o8���A]x�g�̓xڹ�MD�;e�y(��ܽw���`0Ɓ�|������_-�t�P����//͝ɚ�(O6�b}�0FC͚�1�jw���<�T%�������	+�K8;�5o8��Q�8ޓ�J���k�[A����ە������{ti��r�7n[w��)yu��2�w��<Ŷ� ���#R� 7u$�I��WKY���=�fku��oV*�^�g����u��W�XWpy���䷹���.��N��q�˞h�y� ڎa��@�-���>�������i\�i�=K=۔��U��U@��ز�>!��(�G�ׅ5o۾�i�����^�V{��zׄU�9�HV��.����wshL��� U���#+M1;%h�����έ��l}���R�n����[M\�*�KCk��(a�r��_�ϯ��܊�o���-B���A��	���Q�Vpr�����?ZQ@Y�����c�G{�މ���I����Z2�Vu*~[!��\iS�M�䓵�3b����3��9�#�!�&}�#A�̈
ⰾH�G����jp�q�8�ξP��E�;E����ƻ:q��³Qi�$L^tS>6��l����n V�(�$����`�;�#!� ��U��B9�T��ݢ��Nj�S�����H���H���{�FK=`kҨ�EJ�֝����)�7Q�5�k�5�j�#˒ZM"�c�N�r_�2L����c�_�U+?|ɟ�n �y�g�=�	�٫`�Խ�����=Й�*)��W�
9�h�@�r �]�,
5��*�[��A[n.�F;�L��������;y<���� H6�9��S|����eFG����F,�0Bq鬕�U���c�ō�W�� �*M9�R���1�Zҏ�cX=�W[q^u�	n��vƧh�e�W��Az�w-��*h�(1�{\Q��i�˳E����vv�U��]�u[T1�1)�0¦�Lh���ɘ.]6";s����_s�x��P�J�H�e13��=�d��#-eF'����6f�09%vڬbДvP�c�e[j����Iٺz���AP�"���֮�#������kz��DP3jt�i^���6|�r�Wb��p���8*WM�Pa�+e�`�����H'���6�`䇫�|���g|A�k)�$�ʖX�خ��@��d���%5�:U搲1�������Z�2�;-A�Dˡ�PJV<����J��e�جѲ.K�[6NVE�6o��5M�����i���j��ؓj��%�u׳ �C����1��-t0���`�@�ka�h�Fb�ZcPJ!���[&^9�G�|ss��*�w�ǝ1̻��[*�Wv��In��QZ���S1��@:�g�3Ϟ��gh�m��\u��#���e���-��{ҽD�-��fc����������5[�\��y'u�T
�~�E��Qi�F#���bl��S7tG����t��)�[k;�S$��ͬUi������F�5.����n����R�d��	n�#����Ǽ�h/r��w��_$!<�\U�E�8.�ڰx6
�ݙU��OKr98Dm-�:u��os\�����Q�k�^��]e��׷�G\�:'�ްs���_\�ÍA���f�8/�Ʋ�^�Rb����7��T ��f<ߧM�ծ��ZƲT��Eڼ-���G�]� �$˻y֕����Wq�k&�����<-bo
�5Ys�$�*�MRI�1��ށ���r�SiV7K7�U���s����JZ8g�W)�e����9ۤ����U���|y=��z���h��%��8�s�nu3`ݗ�TpLP�y���]dI0o1��3�����!��9G(�[�X���@[�4v�Ȭe��o���;�[��Ē���t�^P̫�݋��-+����x�gs�1R��@p�S�V`6�0�N�Ӡ�,:S����)Z�%@E�&)���)������,_Cϰ己��W4�Q�og E��VM�x� 9Def���#o��f?Y�!��^��@�`��E�Ȼ,ܤ� !"ՂF�6��t�GO0KX���R��tD�ӮnH���z`�A����;F���WVl�nVCϧV�{1�x]' m��V��!������bLΦ.��iE4Ldi�k��n1-|ރq�+���s�g�h`_Q�S&a�1P��@���X���Eu�vT�'9�@�ڴuj���Y06����������E1��hʛ.���(k�Z*��U�Ey�8\���<�ЉH=Jg�����x��������?_���	O��Kԥ���4�����������������~�_�a�@=AIIM	@hЯD� �JGԦ�:$wY4�ZІ�OQ�z���'�C�A�:�:�IH�iJ�z�5�8�R�PPu*���R:J(t	�i�j����'��=HkC��V����A�� }�@u-�CH��@��P=H4�P����}�C�Q�� �]`�qiI��z��b+-x�ۓ�i����⽽�wҋ]Yr^.VF00�r��Z��j�qy��;}y^ÊAT�}6��i�g��y��OX�n��a���;Ŝ�UH���q�N�K�탥�n�w � ���1��\1�N�M>����ƛg�q���l�Ǳ���蕈5��Q�����i�v�'�]"8l
����M G^7ʔ��2ص����xX�n�Ά�ɼ�=�F�q�� �1�v�3\��1���pbXf�Va�N�tF�e�W'��w��1�su0�d�x�%S���<��9�[⫵q\or�N��c+��&�P6�'i�z��`Q�qXiEh�O%�j�g33M4Y��R�_c�:�K����a�2��c<�o��C�7���'��⥪8�?n��{�ݙ�8�fϯ���T97l�v�u1����T�%�3��Nb�݋��`�|χ�f��������.U�:�H�+q�:�G]G[���m������a�q����y�/��qDH��:�:�s����TEI�m"Q�\��h�S���:,r���X�V��=�=��җ�Om����G����-~.�������:/+�๧YN1�T�ij�T�+��1�'��Tp�V�7�x�J�F�7����i{R�h��Uy{O��v�y������7����ſI,(��{�j&��� ,$u�9pw�j��߲8 V.�ٯ�Ά�T�M�8�|�t[�,�@š�fGx��2����;�K@n]:�u�U�u����O���&�:Ǫ�%����k��}�]֌�v>·%��h�/�\��9Jt׹#&̚�����.Lbg��>#1��_�-��)����b@���5q��{�*V^����v�K ܷX�����>k.�gf%��H����"�}�7�%e��J��m|��=��U4y�9�`㰻�^�r4d9]>�6=�e_��Si�Ņьk���f����򅘞5�OKv� ��?κ��3��N��X���h��4��C�o�ޞ�"t���N�ki����`�3��ޡSp�.5��U�x�c[����Kͺ$�6��T��
�kt����<ն�m�w�)k\���r٫ ���Uz_��ǹhv��+���n4 �l��*}�~��*' >?Z�M˿A\=��~U�U2r���D;3��8���{�����_E�.<�q�T��-� 2��0��v�t-syC���ԃ�r��xxx�=�P/_-�~=Z�������o�?�����&�N��=Ԭ*�6����Mn�yZه�2d�Ǝ�d
0�t�1�}�9,$'5��2A;ب�BE��@���`�]�j|��6����9���<d瀔
�v�h�&I ٖ��&a�\��1�tgb#p��;�r}��ιڐ/��:��H�kl^G�#o��^�h�[QwG��l�;��;��^_���/(Y�=% d���wx��P�?]*�Um��VgQ�tG_n�6D���/ms���e���d$Rp��m3eت�����ި�x{�6ǹJ�P2����\ә�hݛ��q�:����t���enAQ��B�JIb��{�s]ų�+�֮�� �٭nt댘u+�mz����A��_.�t�O�Ĕ���>�/q؍\��{b�˹M�L�U��6<%lDm�x��$����w�1�ᙓl��D�����l�/�p�1w�i�\��oU_*3D]o��a�<�N����}���Ӟ˵��~��e���]p�i+�Y��m�)���VR����C��څ׫.��~�A�u�V�X�I��<���{S��;�7��y�vɷ#����������8��Ϸ����O��'�·��[�t�,���|�9[�M����6d�'	R(t7{������^�җ�M�n�ocgv絖��;�NP�RhZM �ؑ��ys�D���(�w�a\;�����=�b7���j�t �9:����{�/ R�y���O�0j1�(��Aڪڎ���b g�K��>�R#eH}ڟv�[eQ^T���/+Z!�x��X��.d�6���R}�� �p��#02���B~u�G��r
����m��<$�Ѭ�<cǤGHm��n}�yA�.eg>
��0ؙ�]ucPGI��:&�n��YEw6���7�WgPmf#��a�Y����7�T�O�Q�	^�t+�ؾ��Gr �b�y�v
3�O���N������<j k{ͮ3������|譨��W�t��I�+�K���#b����]�s�?j��#Z���K���N�\��w��ŏ�Dt�\7 k�_U��;r�3�>9����%�
��m�@��m�܊��/�dp<1.�9���1Ƨ)Fޞ��Q�5��gӨS��$� 4/�����W�˹��U�{�5S.̰����z�/��V���<-���D�/l�OP�|`$:���6�$u��,h���%ߡ��:��p�zqXu���4$K�#��a����[^E�w{�c�K�^��#�M�y��^H��SAR(G\���M���۬�����껌�b4�_	It�IB�9Q����W	�[<�'50�xH��枙�ɘ\:�1�7efךd`0L׹ץW�T�$?\t�F����=��]���W�6�hÍ�.�{�zRC��I�^V{�Ǭϛ1��"��xݑ+8�Й���+^֦�%O)K��ص� �.���sD�ܿ��&;'o��Ԗ����􈅲6zz�FW-sei��Y,lv��Z�C���%ii���q�w<�f7"o�pP�jg���uk�A��e�6g���Ex�U9{Lg�͐F�1F�m�*_3�����FJ �R�G�yQ���}�;�`|��o#��5r�ҡ�ڄ懕)����F[50ih:�(9�:�_	$�c�l�}ٶ��vV��f���d]%��7��8h��g�����\ܶHo.����d�R��zu����������;}��ΟVΥa?-�'��{g��N�l���o�pF#F��J�b����n	�5y���jbP��j�仁}�ɻ	}>;fz����7�A�1E`Ί�1����E�5�!hf�ǯ��� w2O4fe@�~ގ�����%��3R��,*���
��F���'x�7�fv�7p4d��uE�֘�f��c�l׌[�,�B�<��7X����I*i��5n�6T���n�C��WGU:���`���zb��oQ8vY_?��1܎꛻p��{��=�VH&��GZA맇40��p`���j�ݢ6��e��{���;�F�r�G��.uN��gD�_��.�m���Y0��'�[1� V�Z�5�J��4
J\��ݬ�C݋
dU�zߔ�[d.��}�Y����o�����$\tf�F�:EX�Q�|��f�f
W��9���qW4�<���nn��ru��k2���@��5�!�����{0��u�� �2UИ�r�?L���2��*�I��a��kz0�f��c�V`���y����+N���[[@����	��\���G`�ս/�V7��'�xxy�|sE�a�����hn�Kf�m�)��_�l��̞^���~E�m�T/�G�����	��"M	�،��5�:7������Gy�A������H��+��ޑ7���[h���E%�'ԩ���s��)c��Ü55�A�p����{�_�s����ǯ>M:�E����<��q��e/gH4�݌#�gOt�3A5�l�>fN�<����8ҤEgH�4�ɹ��Y^��J�tx-��u�%�_��4�Q�do_7����~�@�y��D�r��H���;�u^�B}͸��#D�q۫�#o!��(��<e��mp2�$�,��5l�1�{O��f�^��{)yUo�<��t/��<*4"�7|�r�\��FJο]�]8f���۷xȎ<�pT�/�/��1B����w&���ʝ'��y!���8��;��f[O&�����]�wU�E�,��\[ ��:�>sLI��~t��裺f@:Io$�¸��,�5�t{�[�����Q����\���}����0��6�"Ŵ܄�Σ8��q�N0!+F����3�=�ǫ)��������/�w��y��(���stG'�7^���V\Җ�@��Iv4��SsN\�Wk��4\vf�I]��H�;cΡ���q�D+q�%K����;F��|X�����Ik"r�٢l��uV�ӓr���"}|�C�J
=cT��~٘�ͻ�6x�U��6�}*��j�}���1�/�x��	��S����*���[9Y���Mo�����U��r����:+jx.!�.Y��]���.�;��@�ց�IW�T�E���4��H!�	���F5�nOn��?6�q��e0��M�:�$�ˋ�^5'Z�;A5ۖ�]V���
�Ty��u�P�T���wVrڡ��Y�vM�&�
�k4-�����'1��h�,9@p���>������gMF�4��v��X�ս<��y�4��o�^�C��7��e�gR��n7t�2������b�/wv؈&(h�����^��#�]B�v-3n_	c��zr�86��nl����o,{3���֕�K>5���>i�`i!9�M�+C���$ȍ�.^��ې�y�-�/M���8�%��͢W��J�ڥ��/b�e{<ޞ��K�p������T�ˣ�dt�~���@�������@��G��Fr/���ʧ���Mr�]ѳ��}#�3��0�.2��Z��1���p9�$F�H�l������ Ǵ�G�ا���$�eW���;C��.Q�WF�k��D����	^�/��_�T�U/}�dn�ͼ��*�u��^j��v^���C{�4��g��.1�?��nx����3h��r�A]�m����&�c'ˈ[Gf��wug�-��cjv����O�z�WOpc�UA����ڏ;S��Jxˢ/sn���v��u����1����U��V�v�]9��y]�t��&/s����e��GC5�ӮQ�x���Q��T�V:�ԍ4vB`�V��j�HF�Pk^v�NS%7��В��מ�<��Y�=v�U�6n,}XW�X>�nZt+�g�1P!Qɻc�!Q�WL�R_Ye���͜�C��I����y��G�w.�]B�f�Νk]���e���]�1;\�>�mD��/�qU�; ��	N9�+n�:3�*�R9y�|�Ƿz��Lt��S��"C!��r���n��+.!d��b���4{l�<�Թ[*���N�uWM�]���1����T������F�����.u;�O�h��g/S���;[���5(+� Ǐg��Z�]�u�}�4�5ed(ۆ4b;13&�z4�;�(��W�(UY#i�瘌�7�D�;0�	�N����Q�A���y��c�՛�]��I�2�Pm�H�1��3����Z�z�����B�d����6��nق\OQ�9^��N��-[.�;4U�,��f���k��mA)P�m�_Y-���ws_D��������fh:&e�f����y�T��F�k�9�bx�/3Z'#5�t�^)���~91]� ��?�lzs���'�"�=�/s`^g.�w��R�d3�_k�ƫ[K��;A&xa��jNr���=~����������?�n��ETW��"���y��������d=ϳ����P�Ox+ C(ʰʰ�0�� C
���0���C�0�Cʰ0� C"�0�0! C �2�(C
�(ʰ�0� C �0�*�*��2�2�2C*� 2!�C*�0��CȄ0�(�2�>�##�0�00�2�20�20,220�0,#�#�#� ��� � � �
� ̠�����0�>�  P P L��p 2�0 0�0�0 2 0�2 2 ]t�S
 C( C* C  C �C( C �C  C C
 l�i� &�i� &�ba	�@@�`dP��z�U � �@�@�ffdi�di�`Se�0�4�$2!
M0)M2��L�"�½u���C�0���C{�0�����2�2�2!�C*� �0��w���{�>_���� �*��(( �'�������;�����ã�?�d��'���|����(~P�����/������������������Ȋ��@����ȁ�?�d����~�����ETW��������~t����v�����z���b�F dP@%@ �ID] R�  P�H��$�H������� #" B� 0���"H � 
� � J�� B��"��!*�(Ȅ$ @H��@��,�B*""������?�?ꠈ�҂)@�P (�� ߰��g����=�?S���
*��?��������������#�{OA���������~�截��ڇ�'������'�
�+�*��އ�!��(�+� �����UQ_�@g��i��}/�>��0A�����?1����?��=�H����H���航����(���~��C��i�Cߜ���	?���������?�����������~�!�)?U���~�X8�������^�'����h�����A}��d�=�wA�����N}_�DP����:A���E]��'����P�~����d�Mdy�ל��f�A@��̟\����}��R�
���
}� ��4hYm��MkLJ����Qm�l�
эj��*QE4Q%)B��%-4�!R�ĥR�i�l��jd��m�jU�����2�[M�V$����KU���`�J�fY55�*[
����֠��@���Z�T�"�5�X�������V��mi�Qf�k6�[K�UL5ff2�J�ڛҭf��7m�V��h�&mI&֭,�4)6�il���X+-�IT�=��Hl�ڵ� �����5L:`'ir�p��uNZ�uҩlU�w���֭w;�9�vN������ݴv�u���o[�m��[5�޽b嶴��m��+m��m��4we[��T�6ԛ� ��=
(P�B�����C�Р�wy�B�
(}
��xt(P���[����-�!��j�v�t���]sm��.�m����h0�-���]���Gn�:����Vu�43b�M���f�fɶ|  .�x�i��.�}�q���WU��٦��;J�N�jt��ݧ��u�/^m��t��jW��4�7![ki�Wmu��*�V܍�����W�OF�w+�aJmm��)�Km�l  ���f�eNq�6���=�c=��T�t���u�L���w:ۂ��F�3+.ڪ]�+�Ur��4m���p4�Uk6��!I���X٩0�� �{Z� ڽ�����Yڸ�U���k��t�wU0�Yٮ�M�]�wt�h��@��r�(� ��@)̤�N��j���6eY�[^  ޕ�Ѷ�`��wAʕ���k�܂z��UEU�w@v����OP����
.��UV��Ӆݎ�U��kccb0T�6�ְ�� �
m�8�A��u]j�u� �QN�MB��R��<�iJ��MPҷ�t	RM7�<��)J)Ku��zP��Ѵ��[I��V�SMRQI> n�|� ]�\�;��hR��^��X�g�o=%IJx��y($;�V�O	�=s���+�Gt��t��T�={�m�
S��,�4̶�͢R��1�j��^�
U*��w�J)D����E$m�y�:((�����PEAU�L��W�{�J���랤�B�<���M�޳���A*n/-�Tlm�H�je�j���<}}i@y����ԣ��.���[y�R.ڪSp��JG�����=)EH�;{�z�JI;��
m�7��ʤR�޶��j�Q_ E? 2�����~A�RT� S�2��   �~�R�� � �7�@�J��jF@)1����� b���?��4?��?��º��J	]o���>E{}���X���
�VZ����}U_W���\����@�������0@DW�耈��EaPUE?��.ˮ�_ʯ��NKT�Ge��%���� ���l���*�V�@!A:O�Y.��J�������E2�MThl4Z_1v�4�eTwXL�"F�0OtmM�V䀥�R��>2PMJ�/3%�Y�L黣�Q	u�����A�a,��]v2�Th���d��	OYF��^O��^bOm�w��PM�b��9$FG��=W)��ӕ*��]6/v�n�˗b��)$ q�c�*n�2&��(Kb����DR�6��8l`,�u��[N�Y�槤Ո��&��w!J�U�q��xPں@@�((-�jh�7s�AMִ��&"�3K���kEe�[�S2�s+m)��n=x�he�n��:3)8P�t��F��y3^��kkݙN�N�k�&+�Y�-5�f���d��l;�����寞@v��l����+��l�r���t)�r���QͺOi+]��߆J�f��\�1��Z++,�KR���Vfڶ\�pƍv�e����R�`;Z�2	v�^Z��n��n6�7(�b^eF34 q20b�{T*Mn���D�����M#&��.ʘ��5��Th�B^�F��#.�r�%O�%�e�׀��[(=��U�y�&����K�4��O$EkYL:Um�8�[m}z�F$�fܨ�k���U�ISMf ��}�kOL��e'�m�8�U]˵i�%:8L7Y#uyx��k�'f���Z�2V^�e�a	�n�R
n!t�B��ƛ�T-͆�Ԑ�wv��8㕏2@��9�����J�)��i�A 3K��3�A���Ǹ���u���r�ʤ���3q�o����9�H֩�a�J^=�uYq��!ShԨ�;��<�v� E���F�N5�+d{L��W�:�䥫`�4�4
��( �u�S�m,�W����Ҋ��M5��˦U$���ӼL��,/$%�u�-�.��;#Z5w�&�q�Rt��3����XK�Dz��K�Z�ݱ�sg͗u�`��]�ل�c`�*ُ������F�I�R{b�m�2�����V9d��u��=�:���\ܹ�4Ў�Fm������%lQX�u�[ڏ)nV���M�l�xVu�S�m`�%v�[X	T9�k�9�T~�P�mQ�7��z�7fx6� ��Y���I�M�&��J�K�4hX�fHZ�{{�Z���GCg*!�Yyhc�9�+j�2��6�K.L_9B��!�&�a]�"����%Zĭ���<kh��F�z+Ǹ�n]-F�m]�{�z��k���O*]�8��:�q�+̣��-�h|(\�2�/s%Dh�kw��(HyZ�^�/3a�F�Y7��1�1�l��Q�m�P5�%��mc��2�;���[�&��	���n�h�%�F����w�W5���9�:
�vk]$�7�G��+Q�N�ek� $��gEaV�Xj���� ��&�Ո2��y�޵��7/b���r�5�NEKH����5��bL7�%�@vF��e7b�0L�j����
�ۉMG\�
L36Q�o^QW@���1�]�h����Rͤ;T�[w�Ʈk�M��6哔�n)��31n1�(���Ulԍ<����a`���n]�b��l�����U�P<
*��Ӧ�ccI�9b�b�!�6]l$_�V���Bԥ{/.Iz��{tj�Ԛ�]���i�@E��r+���2���Q���Wt����%�z�-��v�cf��2C+�G*h��k��n�9N�F�n��V͹�/�,K�t���]�aS��8N�*T�E���H\xz��Hd���.��ZeE���P��)�Q-:6,y
�C�(�]�L}6#z��������J�AMXШE�׆ڎ���ʓC�*Ӑ-��	%fQ�OU@l�G镦S��7^lU/q��!v�GjVʹ�e�i��q��,3m���2&9���h@��ct�v�y�oR���ںˡ-�b����4q{�;\#�5�
[h��׻Wo����k��t��M�nЗ#ɘ���6*�'�fd��nؔؽUx؁�^<�pҒPT�O=�u
m��Xr�K�O�H���[u#�@Qd��&�l�dU*���ї }��nX�*��Feꗮ��kr�}���B��0�S������5(��X��%�D�.�kvo	5�%c̍^��H���\��%I%1W+�0@}w�w�n�ͰRRjb���vvms!ͭ����pJ��n�elz��0m���&[fC�ډ@O�ML{(E�U�X�ѥ��"^��qi�ݭZ&�A4�E�޳j,����m�]�!:!v�9&�7Zp=�S]p+ҝl4�^e<t��B�F�C|��%��M5����i�@/�ٲ�U�:WCVP�lY�m�2L��W��]7a��6�@m��K+f:�N����[��T���s��Ct)�o�̾�˱�W]���<�]:_%�`��yIn�"�i���V]��NK2n�M��f���=��+v�K\�aȵ����t�hHF�Av��{�.��dU7X�E��Xȳ3ibJl���n�)
�y�fehl%#חLn�����*c�m��<���^�څ�[#��H������e]�X\�S1���ǆ2�	�pnѤ�^E�pn�#u��U����0�Zi�����d\�1�X���݃s-��j�p�V ,�"��:Q=ʘ�+c��GM��W�j��*㙊ٍ��ʔ���3z���o[�f$]�z���Y�^le�[����2�i
cq��-��ˋ&�ԨV�ss]�W(&�&p30
T��z�է��j9W/H������ՓM���oV3�[���C���������%ԩQ
��32�r���G�]3k	�1�����p4 ���#Bʵ������"��]4݊Ǆ6
õ��oF0���B9Q�1�.�![qCY7��!0[�˺���0�VJma߭�,�j�kv�G����Lbi�Q'(+[����W6%B�=�@�f��:�+��a��$j�y�wt�lU%�3i�6T��i��r��)�L�8^e&�Aj�����e*E a�q��('���{W�.:�������U�-J95���L��])��M�5u���{�A�W�S��GM��1�#�4�4�
��.�r�CL)f@� :q�e�3t����M�[ A]ff�(�b����s.�f�3N�$9q�7�m�ug1e%���(c,��jt� ��Yq��� `5��Ta� ��kB[L�(�4�1˼/��qEN�t!���Y��Ap�v���5��EM���Lw#�i��j�f���!�{�����r��ܛ�vC�+B� mGS09wE35)m#y,�5p)y �cP�Bl;q/��/����k��DP�*��4��gm2)�.�@�r�,޻�vޓ�D�y��=?b{�S�V��HWIJ�$����������$K}��+-��+ֲ\�tֳ5nk���O4ZO@�&�-䳗����ł̅12�˰�Y7�S��i"��-՘��s��%�gNGr���Ѭ:���abe|qnJ�R�7�[I�cU� �9B���M�*���Abk�@7;o-P��r�I�D�z拇*�;@�� *[�t��*�:a8f����:r�zp�jD�3n���T�SsS7e]WJw9M]����[�& ;��S1n�)O�>��QbA蒍ñ�ӽ�lܰ�QRvvci-�����@��� X��hj졪 ������`mAzq<����D#�7J�(���~f*��T�&*{�؍n��%����8�\Y�]j�Y׏*4S�l d�İV�����i�fVd.u6�(W�NK�t-d�2QU2�^f9*U����Y(L��qU	M�U�0V6�sm�laW��1�tNۃ���۬��nQ�'��{���.�6w�Oǘ^kуR5��لV���3Uh曨�;�.Q�w0��y�����Q k���Y �5��~2s�fk�Ҍ �v�pJ˻��[Җ�-b\)������z��{�P5\�`���Q���,#cS�ϕ�%t023�����.HVт�L�l��hZrd�w�����*�T]�jØ�b����j^\�1C��12d&����������2��1���ͺ]�Xd�˩�SsJ�)�.]Q�hn��BT$��zo�u�1��*okZ�X��-;Oe���9v�Qi�Y�O��4�V�ѽ"�v�e��S�H��LT���-����B�1�t,��Ś&�-�ha�rR�HP�u�j���(Ŧ�P��n��G$��CD);3B��t�Pa�q�&Č��QH���6	{����+bTv��"Ԩl(�YP3���طj�n�`��*'pmh��#6�2WN�x��ՒL�Q��5ֺ�۠�6қ2�R��E�U�Hj2�b+t�z�`��l��;��G�Agn�rT�.���[F�����hJ�U���d�+B��u���T�O!x�	VdRM�-��%Hv�$f�[wr��t\���a�/���53�K��:;�=Tv���%7pT��A<hYg��g�#�n�ܤ����N(f<�j��zR�I��p�˳�D���V�d&;�RK��4��N�h8%q}.�:L1m�cչ���P�$Jk���O4ؒ;�{l��dm�[��Ȫ�tRv-��G1�l���o��2�z���a��{��)���!�EU�iY�9%����GS!�����	+%�N�ړH����qT��YjC)�ϝ�M�͇OV3��Y���}�	z���kLm�TC� ޯ�t���;v�4ia�Y��y%Cr�ID� ��I��E;.��d����J�1f�5��HL�F^�������Tf�)u�4;y.KG`,ѥ����g!������6�h��G�V��j�|��@f�8����$Sr���B�6"����%����D���H��4�=[-	�n=2큘�|�R�l��p	�/j_��w]9��x�5��;�A��	��Tw�5�f#�eh���a��ܵ ��p�c�u��tͫ�ȋn���.��<��(�\̼:M��1���1ٵ*����+XŬ̤a�2	7,��ef<P˻��a��(��f�H����oATE.�k)ͶI����F����fm�mn8���Kf(�R��Д.k�5
����5u��%1��Ա(��{wa8�̬�TE�U��U��N��Y5�9�m�z5#�+ru3T�SJB\���mR�g5�*��ōf-���2� 9vh}
��;Wh"�eaco3��1�!���7pi�,�y��.�c!J����6�	jy���cw6�f�2��W;x�jڼ(fXbq�N�(�:R4F��ͣ��M�
�^^AK��71��GQ�Aϓu�������&KB��uf��JV	yhŐZ�ި���&�&����"�C���X˸�hJ㸒͵�h�k�:��ÍmХM�F
S�̉m1�m�6�`���������Q�S�6⿤r�aՆ��j�Q��j�ӭ�gJF��`����oi�U�P�+;�̓FlhyZ��M�W��d��K$&T�
�*|Z�%m03 �'�"�Rix�\`�{WcP�u�pbG,���8�� �faNQ�4)��̦�V�4A��֛u��*څ��w���n�BP�ڼ9��9$�ģ�U�O3wX��z�Ya$�Ϯ�Cv2�
[�%��Y,�F�,�.	NhrԂ͔qKi��5Ѷq�Q�6�J���C�Dڑ�Cn�y��j��*���a7{F,��n�9�ܘ��;�Z��+ ��A0��)Q�V�m�͵74�� SaI�дQz1kf����D�xc�$W�V��׆��,梋��ic@�2���[�5��wZ�փ�]�yd���j�e �M�Qƕ��^f`��{���p2h֭�t�ŧD�iHm��I�q���y��#R֬����I�
(��13fa/�t��֬5�+n����a�Ekǉu�C׵�Q�W��[8�sȫe��F)"kd0�bi��v�K��^i��%:�nHU�PstW���KJݨ�$63f̺�"5梬��t�[؜��>�fU��c$;�5�Hݕk�Dc�j��f��;g/X��U�,iIB�m�"�՟E 9@�V�>n����e�l-�����I�H+u�J�q�w�9iw0h�7|�h�a�2�уw@M��J2�@p��I71�RfP���+0 V3Vٱ-��Ƣʵ�x���Y�8@�73@��V\�7H`�W��}��Ab���d{�YW2�@�9j��}qZ�
�U�ȉ��*[���pAA輥(�j��h���gr� ���������L�kf� �ԝZToI�!RGiP�V2�9�@H��M�@�'n�`���J��#bR���u��� �ݓq#��J���)`,�scS U��ݸ��i���Jn�t�� _Wp9��Ol�^�,[��ɥܗ�0.h���ҎlGL�َ2i4t�h*'
���[ӑ:��l,z�e濱Vy�&N��̰ܼ;��q2�[ג��� �bQ���3��6l�����T��Z�`4~Ӕv��1���26n�:�dn��LJ��T�oKš+h�M�	�lͺ�.��92�Y�n�M!�1�3[(*ŭ^��B�ns��(��,�ɩ��C%�[M���J*��6�!y[!�͡��{���ǅՋG35&-B�&GZ�P���0�y�� �rVK�Y�\�
���*¨h޷E��)�m�4M��Uf�Y	��we^�G,�2H�ʸ6�d۴��ң��#y�����-
�F��y�9}7ZP�e�<@硊j�K�LR5q_�Ex�nAyW�:ݕ'w#�e[�Ə'I@�:&?k��-$+T�&�]�	S;m�����o>#�F�ܸ�z��v�L��sN�m×¹t�%�4i�stwo�!���$�x�+�ޮǚ��m�{6�-�ţ�[Z�u&̉�Sx��^
{��ע�],:}Zû�Jdy�M8��Z��b�h�=�]���%}0��Zk)�Ƶ�:@2��)��[e},`�3���=�E�QUY������η�!���X�y�ނC������h� �M��).�s|��[/��������|���c��W(���&�ҙIZĺ��d���W��~�q����ǻ1$W���'��/f���
��մ�c��X���O5
'2�d�fMϭ�U���/���N�h���V�(�e�Yh��A�����--E������]�8��;-u�34�;X����@�7�ϳ1��bsw
��� PXe+��}�HJa�
��2ZZ�4�O"�[c�����,�'ܴ�7u�PQ*�m�����n(ub�����s���9�D�&T;���S�攁�x�`pu�eVb)*��*�pvf�>fSN`ܾ�gN򬛟*��"H�hm*�<�(ʹz�ٲ�c8��Ҟ6�L�Tn�j��q��p�q��o.��ޗ��k*�.��;
kԱ1F]ͻ��4SR�' �˾�1˻�V�P��r���x������]L�L���������뺥 7s`
sX�C(Q[�;�e�C�ۅ��lʇ^Ʊ�ڭʈV���v~8g�w!�ԧ�F��j]��h�s���ں�LYݛɌ�,"�@��]զ�3��&R�@;��u�V�ݸ	��Sj\�@��O:^��af0���Q{��:�4�B�p�ut��j�|�,��dα0�,�e]���o1ZǓ��������8fW���=e ���� &ۡ�Q��ޤ������}�*��z�^
�*%�2�n!�ŝ-�
���0Q�M�BV�)��Ӻ�N��vA0��$[I�# �hʖ&�6���D�}Y�� �jt{��Z���K�e�[̋�W
:��ٟ��g*%��7��/�&�\�=)�h���o7�z�qq������0���X��:��(?I�2^;�v�#�t��1V]���貟Qy����A���rRJ�2��*�.�uiY*�*3]�Ʋ�N��WJ�:�L>�1o!�޷n댬2�ձi�R^�_/�Lˑ�����H4ha�ަ��u�9M� �;q|�/��
T�H����"jVq�]�|Y1Уj��]�a�3���k6�넍���w*Lq�̫��v���X�{pc��c�h!�o���H�"7�]��v܉lT�["@���������]�3o	<6&�՛�7cFj���%�r�'���MM�T��z�\�崣"�q��k|�ӵ��g2U���9��7�]:�F#Yp��ԑS�W�t��ł.����$��b��{�ٛ�a�)6���4�s�Wd2�-�r�4A�<�Ջ(�ꕘ��O�Y�r��"H
&��f�Q	v9 ���aΒu��ll.�(6�[�De&v���1����jp6�e.�>{kk�]�&M���՜�A�(�:n\����
Z�J��L���sf�R]�n�j� iJ��MF��Xh9���b�dWP��Y��v�Fx�F��ψ�9+Y>�!��1rtU�j�5���)���{"�٪rs��vP�x�wkWY�J�9���s$sc}���;��놶J���k��%xM�(i(˻����VXy��p�P�1ge�/;�2�`��|c9u�;� f�.\4����j�Bk��#��O7�(Q�Ez�B�٭�&N�n�����
��k{���P�*��n�b_|������dP̺Zl�!��j<�f>=N���uX�Z������N��׊!��]X4�y+�/��}oj2&��У��׌�m�+���N��b4E����pS�y[B3�Ͻ��B��&��A���d86�&�ĝm��9�%wS�Ei4.��Մ�5|�T(
9�F��=����⾔�*�_#:a��@M�ހ5*A��-wQ�T9�x_)����
��֧�'w�İ�y��м��B�Y��o1�9nev
Wy�����9o��ySm�˜�=2�%�3�Ǹ�<�:j��t����N�<lW���B�6�V���mk�1A��3ܒ�20�Fd{{=�Y��\֑�����]�d7�)�$��zs,��"�:6�3--�/�Yr������Ws5daiL�1�]`Sk���"��|�Thoi��u�ȷ�{H+����|9I�i#��U�X�څ�]�ST�&�*�P��Y�G�`�'q�6��w��T�0���ʼ�S�H�H]�)B��6�� [�`�b���v���[�2�	H�{fcjIYi�˱]|]��[�*���=x2xsG��]�D83p�X�l+�M�z^�w3��o���<�M��l_
�.L%�&l)�ׯY�9�mI����=�iz����-��Ի��7D�t@�'J���\�Uƛ�P9�k�4�8�2��𽺈'�ȅqX�Å*cot`i^��A��F,U�r^;RX��g j�i�HQӨW%;�K�8��nf�qN�C��c��e�r������6�(�V2zMo��wZ�E3.�{��꽶m3�\�q��O��Ź%�C��}�c��"%�	�)Ey�����ѧC�Lp�oTgG3Z%*V����fS��o��eR�&T��Fz˽�Zǩ�{����R�YǓ�F�8����}x�9B�i]-B��O�ӑfM��k�j�[W�����K��dd���o�2�bqU����ʗ��nZS����H���[�2ҙ{�/������ۗ��	
�����Q��y��%F�55�"�e�W:Q��W/q�t&�J��lU��v�;���\Wa�]v:�1�󳌴�r��C��lK�����	
��Out]V��-�suۗ����ܳ)Y�2VQ�*!�A�i��Rgp�g�^�W���V(����\<��;����\��o#@!�:`2=vX�z`yF��ح��� �Z�70c|%��yn��o��+���ث|���bv��NI�g���+"o+{l����j̻���a�e�B̕�$+ m���7{Y�O�s�Ϙ�2X�\��gV��寋�2S�jӲ�lm�3�Z�g���"�npCMGs]�K ��(Y�ev�@��2�w�-��{�;7t�yKi�����r��m�	��]Y
T|L+��;�q�)M�lȬ�ښ���&o��i҈�v�<�Ut�9g�ș��T{��ڣZ��4�m�1��wg`��A�+jn�È	D�me�Y4u7�ͽ�$q��-�-�=��m�y�KXdvgG{;U���������@���;/Qk�;K\�[1��{-�[o9>ڜM�{W����?+�n�3�sxܓ/1FU�v�.��@Y�u��&7�]�vN;��*q�1�0��ۙ��c�ޚ����0����ykY������36��Z���RU�ۚ/e�V� L59��I��ۧ�6�]��ؼʀ�m7;N�R�Y�A��R.��w;&�#�����ػ9��3Qj>�:V�f	X��A���ҩۊ]p|��u��=�5���kp$�r���Z�{4peBEnс
��nd\nY�y��M�]r���u�M��� >���,:ʩeK�7;t��H�3o���o�u��T�/��f�4Hˇ �M�rݩD-��AH!غ���,��JJ���\�h7��Ӭ]U���Bkϯ_GJ��WXA��`�D�H�U��]NV� c�R����usy�ToU7� ����]�B�P�s�d4r�W�:�{�uەpu\Qnv�g%�=�r��5hsy5x��s7�̀V=;l'���c�����W�/}����뮟��iɵ�t�Yu%gi��
�u��mc���J���-[�ce�2�
@�ި��S@�r�f;q�c���YS�ҷ[ ���]HGn0��]`�N�̓S<�,�g�<�n�9�U�3 i^�HOC9�_9Xjl�cB�n�#t��k���R��Y�n4=�H�#�=�q��g�4�S����6���(���N�W[�5eI�ݫe��1�N�X
̵WO
ZV{ennFbm�e���N}��	�����tjG��Ƴ�����3�ߴm*�L�/���k��<凗S>'#��H;kf�������t$�o�^%s@5V}[؃Z^1?Y�pˌӥ/��J���u���W�,��6����ݮgR���U��6h�ۀ9�� �0uB��r�b�}M^���Īu�3����ː�L�&_cx�@s����L��"(�=bM�G�>�\�aZ�>��8�*�6.Ә^w&�� ��_���i·C�4pp�N֢�N��c�#ݢ�mm�4�gP�ͧX.�NT)�:��������¡�U��	{��c�o*]t��[�uw�Z���X����?Fy���Vmθ%BD�)���.��Jy%r����P4�<k��׫>��3��󚌴:$�u.�Q^�)-\y	2m��b�k��u��{�ǔ��r�j.������ |�EE�.���L�I���Wh_b�������blW`|{t�iSL#���蝂�D��GI�3DB���[J��+]�7��S��vy]�t��bRp�H���Iܕ��W
)jS�X��|S�nnk3�Y}�*qf��\Ω�\M�4��n��Y��9.)L.Mu�_	�ppiT!�\g�B! �Vu�}�7Tr�*}�u�u�H܊I(��uc���j�u:�5�6� ��'�ɚ��o�n�j�"e>7�u��`)��Jx�s��#�f���8N���g4=�� &�b)十h징"�@4GS��*���r��L�|q:
���{�<�X�:�B��>����XU�q%(mqh��h�E�A�)_T�GggG8��W��X�ʛ�k��.��<(�vUA`d�(��U�&lw3��W>;q\]"slsô�]'jò�3b������G��=��*+T�]oK	����	E��������<��n�ĜVH�Ru]��d��I���K�����E�P���%��Qp]K��qf���������1�t&����
�(�l���l��)-�l��.�s����A�������X����xP������F�� ��w�%�=Mt1S{β^��e�H���2EL�v�&�����V(�f�����q�&�y�*�}�h�H*
e^e
��>Pˠ2F����lp������i���"F�<��;-WX������b&&:�1��F͎N�l�#%s�����I� Ŗ᷒�+v��u"�O-���``�z���{q�L�Ȧm���;�wj���v�ozVKgL�unrM��N��f��:S�fɷk��%�. �+]7OnI�+����8�+�4E>���[�!�^�-ʬz�;�`����*P�pN�05ZZ���gYU����w�6�[c����07�tri1M+v+y2�3+�*Un}�{�)L	�LL��j�v8��;�^]Y:��bV�o�j�	[r(ۀ���GFb��q�A������j��l;x��z��dX"��"Eۭ"�VI}j�Wt�5�n62 ��ɩs����q��h/�Z�s����+�+�/\iL��K1��`޿u6y+��Y����ja�-*q鋩mY;]�"�[hgaz$ �)�r�	��x�\x��`|�l]��LU\��w���u�ͦ���2�bS��&��ZPVT��;L��V�i��/%7�J�V�K�@��i�����{�2A'$8��0��嵫K}V�:��j�ݰW"ŷ���V�Sb� ���Je�
ٜ:{���j3����y�R�s+��0�"P;�*� xZ�Z���ʔ����6�k����mۛ�0�[���m��N75�ɓ2��̂Fx�8��ǔ�=�Vf-@c��hW[:�QX��[7�fG5:�z�7�c����bn�V!V�md�wn�i��,(���N��Hl!6���=9]Fk�X{�V�4��X�=}J�u�u���	Cc]�4P���]�8mJ��ؤ$��9T�8b����RZ���CӺ��+��(;,�Z���6��}���{%�={5�K�Ԩ`JV�^��HA������7wj|Ti^����ҽĝf�J�A��a���m]���q��70gnǃy�5]��V�Q-�[�X�J*���P�M]�����g���S�D�l�)]�$��	0b���߼��y�>̂�*h,.��Z�9v���nge�O������J<�ŷe��WHM��e8{�]���*��c��*��:C���N�M�6��*��[J�V��;��TYGT�+��iNMksx����]����3GWs-Mskw��k���{A���\*nӬ-}��b��ha�r��ɉ2��WK����\�&�2��ˡ[���]ծ��-[Y����6[Aۈ��{�S��U�	���n��ܻ��ww]�*��x�V=�1�bͪ٦)�F�Z!ܚ�Ej�nV�ߥ)\�K-�g�ً����H�"�n��(>ڻB.�n�б��6�Rb��yۍIh��D���kł��W�d� ��S�k���_Nv��I�\�ث(_���{��J,Z�Voaǖ�"��O�i@�{	���2����u1�q%Ֆ�ڵܞ�*P�;��L\&�d̡ǫ�r��H�9�Q�jh�]}|��7���V�CbZ��ѻ`�|�3�Y�"bQٙ�S��ml�2�t���]KN�zp�0GY;wuD䃮��ұ�]�9�ݫh%�R�2�Ve�]�Q�j�ʓ^^.�4�\�qb��)E�Gؤb��t��9��h�q�2R�fNT��1��̸�6{SRQ�[��5�@7<���zf���}��ηמ������)�����3y��W/	ۼ��FFxU�O8>�H�#�(HW`��]R�9
T�����.�p+:�\�ݍ�"�5J��a�ѣ��yZ���,S��\�>b��Bg���mͼ�KX��=��!��u@�褦l���)�^���԰]v.u+2�Z�S�m༭!ϒ�[N8�t�ʆ�@����m�v�2�n�iXӬ+$���uj�`T$�Z#�sr�g*��y�ʻa�*�;5�]Ƶ��۠�T��iin��a�׸�븻.$a�{ ����I�vĉb�.U���Ç8���9+�PW�j�Q�
[ɜ��Doa�]YWVm@�v"i��$�5dN�ߎ�t���G#�#ep�5u���j�3R0�:*&M*��Q�3n�[+leY�Z��.3�vN jV���i�J��:��ֳ[��[g��������ӻ�Nr�\&b�6����w�L��X�����dl�:"&�Y���jXC�t��D��֏s�P�J�yb��$�[a��=��l�\�^i�#�#��u܈W#���4ްx��BC���kWr���n��F,��:��k���.�̺e&�5¥�\�S���y:�j�dn($�{������ؚ�]>���r��7ׇ��@�DzM��Z�P��7:+��듷�Z�#�#�yo���[qGc�Fmei��'>�X֜�5�q)"���D3�dS��V�M^0��<�Go	11�"p��.� c]�n5��ɖ���ʌ�M뤵.��.M�J��m��%���e�ص�Ǎ�V���6��\�p��>҅�{"N��ҳ���jh=�jN�k�@+<-�Ph�\@o6��ʲ�U��ۯ;79�����ZAFb7R<���0oH�M:��E�v���Ǧ-��Ł�Z$�n��|e�(-G���VA����f��f�,ݠ����6�@e��p��#���4h@h��9�2�\��h����;;q�{s��>SiTM�S�b�D9ޜ=���A]u�޾�%)�@���)�g[Eɉ�J���tmSؐ3#��9�;���%%Z\�
�dŹז���k�0r�㋍8��ڏ�vg�$�Y�����ɬ���a���tq	(�o�ʖ�����;�3���F=R��&������9:�$�En�
W�f}����hV�E֦����W�ڒ�kn�{�ˣ�\o���]��A�*һȻ��b5�����ʺ��1��яc��`�]�2���R�A�s-�5� ]��+%�������}����R���ıs{�p%�^-e��{ս`�ٱ	Y�����|��E�5�f�YM=1�5��mǷC:nT�5�7$��0wcj�f���[��sFS�ɫ
��L]��k��!�����λ���sM�ق���k�#W����8�)�6���N�;�P�m�/6�0�A���ڹN��2u��b�,��s���oJ&���ց�Ux��?
��8{�x6�K������i�s(�%y(a��֭�F��*
�Gx��4�w�u[=A�f��u�+R�u���[ڼ���Vm���"N�� d�@��I���-֦�[�ri���y\ToL\p����yָ�ѿ�K�yV�R�EF+H��� �4M���H��^^���.��n��=����m��U
F�n��/GT�d}��DD����Iڷ�t����j��R��ym,ŏ��*v,ˣ����f�Np�վ;����-sV�ҡ��;.31pU[�2� ��"�����<f���E�]�����j����٢i���J7�v`���V��A;�]�
����E+194�q�
��W0e%�#)Z��48���m�D�H+8^DK���Ib��K!�X��l��L���[��fm� �T���dn�>b�ݭZ����qv��}���ݖ��,"#��� �7*���nT{ۚ�4��o
���Rxz���˕����L(E'O6J�KM���2FV}�n��"�3w0+���^��O/j;����J�V�_B6�Xׁ���y
ueFf���,s�}l7�t �.B���;�6���ٻ���dÑ�U�;'�.�W<zĨ6��l]R$�N^)�u(�`�ԁ0f�.ٜ]v3�$�T*ĸ��t�i�')�d�e3�[���)V8���^Nzְ=Q��G\n�N�P��Ř���#��={��١�F�����8�+;��6o����h���4վ˻��1��9�y7j��I�|7MZ�(�3��c��w{�;}�R�s�[���z�=�N
V�+�_*�J�?c8mn2cu�l�.�k^�K��%
<^�-��V���/m|�/C�',�1�v�r��>��N�˦
S�����De�k�����ъMza�����BzkҮ�ƃS��엗0��Wg8�����[�0=f��hk�;㙕��T����t�Gri��nv��P�o�<!�E�Vf�N�ǻxrVΜӗ���s��\!����N���T��������I�je��ą��Z2�_S0��D�I[� 误�,>�/j�ͩ�/]���x�4.H�2����6����帇8�`Z�F�����Y;�R�ƚ�-�hk
�r�R�tɔa��O9�y�c
�:���K��T�f��x��Z�Ǣ���obY�J����]B٭��F4����+t���m�F���C�n�����ʈ��;�&qj7�865�T�!�Gu�l\�u�������H>%��v�Uxtz��dBޗ�R�)���PV��MճDN�@lο���"u2�vˮ�blѭ+���7����Ls�/-�1�QQ��%CZ�gF6.���>Y.�=��kr���V����:����3�%1�L��r'�^��B����]i���h�JT�Wn�9k��e�t)ݱL��p8�.0�\��'w���'D��&�+�S��v��y��W|�WwW��T����aQĜ[S\]Z���2p�T��zc�6�� ݰ�f��&�yF1���M��v�G�����p��gV�r�!������B��l��[��S�V�G캵�H��k���% ��Tul�ؑXy��RZ۵�T�븷:F�>�5�r<�v��ڢ�'1nݣ\�^H�j��3z�O)�Z��#w�R�]1�u�/��ۥ��mU��n���i)V��YT�byrN�7'F�ѩe�y(�d���1V��6��av\��t�{�[�V)$.���f�ŶnX�}�bfe�z�t�I��=��VK_fJ'DIX��r���S���Xث��J(��
�}���c\r��}ѷ�4�T����ٖۧ�E��̬�#�&�L�v2w��C�%�jOrLv�s��z
�]m�́�d]%��Y��
�չ`GsU��o0�D���W��ϐ�
�� �N9���^m��s��CX�ur�f¤Vc<TN�DT��v�F� �����a��骗T:��{�[�Э�	�kcG#�G���w��slR���21�����)�����/1f��5��f��!f�#�k�s��U4�m�c	���qo1;Y�%�ُ�g�|�Z$Q�x�
��͠r�"a ��Y(Қʎf3���$L�m���U:˵� ��;��\t��Z�u�`^#VᮼD�q�x۳�<洃�%��Y��MT<���1�jЪ�3�0��_r���]�Z�0MG�L�Z�	rU*�*-L�����Ed�-�,f�g|�`L��/(�]�ӽ���묹���`%����e٥{�$a����!E�H�'��;p��3S,"�χ�!�,�ÄU��{1�r��e�8v��SU%b��%sr�m.x�l��}�h������� �J��+��H>�\r��$7s���X�q������1�	eU� ��J���e�����,m��� uҲ�m����r�*�뮮B�s��s�f���3$Z�f14{�مT k��gPr�NX��=��j�)W�/m=`�H�.�m=n�]�����*R��p}�6�X�U V��c Y6Q�:Ō˩��pl�v���:�[���-���V%DP�k�^�{h���^����׃vI�3���U��Ej���,���¬Z�v�NƷN��R�y�hyX{���@V@ b�.�9�=�R�ɋ�&�.����z�ް�KNʔq������t�qv�
�)f���k!Z�
'�\�55�x���Z�e��d�.eo#|�A�0��K��,��m4��uʋ�=enV.�m����n�hv���\y�w�,߸�p�	n�Tja�weثެ1U��ź/'"`�`��h��C4��B�N�U���72��w��5��&������>�eL�݊%q��`��N=xif�԰�AL�$���7�<��#�P�ݥ��q
�ɇ(R����9O��,�sV��T�^������\-˧�[wVi���vPkuu#1���{���'^\�n�Vx�B�T2�X��3��+��@��;i99�g-ݡӻ٭�>�н�[��T>F5o�9ƛ:�v���bŮ�[��iԷ-s
d�q��]tu�=z���{^���W��,l�U��a�]�Ø�o*{#<78CN��ƺ�[c�Ю�|�j�[��z�V�\�����ԟF�t�`N��&����>�ga�\�;�����!Õ�.:ˆ�Q�����vP[���ר���'��΃�2[5�'7xs�NLKt>r�e�d�B;�֙CD�û��S��{Ϟ�7)d�3\8�Q�i,;��|����H�6N���%Ӥ��xU�F��R����5���ԝ���S��,s<����\	����J���8{O2ޮ��
�N�l�o�r�
r���ޥ�y/qH�Ҕ�E��뒒��av�ӞtbR��J��-Y�5�wSz�s\���Q6�f$ML���SM��u�h�V�B�*ˡ;��j�=���:�vN5����%z��N)��D��9�$�	ys�F2�̒�eX�!Pۮ�9�Su�CY�~��q�l�mc�i6���I��!�U�v*�V{+��8�/���p���53���(� k�i31�]en%#%R�L�e�S��k��n�d��-�f!��I�E�,�}K��9����ǵC��x�CۄV�0����d��N�g'q3RZ�C�x�9r��g�΋K��!Ԏ�v*lwX�#䃭�ӆ[��&�@�+(�]k�.� �KC�T�\�֎M(eŦ�-��볪�-��]�����71j��V��i�iB��+V�lѐ�'׽y�g`,��l1�kvwJ�KT�������f�4p[K;nW-�V��M����u�J+cM�R�Y@-k�dD�r�$QoV��0����ѣ�`�o6}�=�Ie=��
�,�a�[�s8.r�t/��'0mT��۱O*�-�~��[�V(#i�V2�Gh@�*
�:�0���cw2�/��<9�9��w]r։�!ԟ`U�m���Pi�&<�EͷRj7x�	G))J�m!��Fqa�i�r�a�+]N�uz�^�nλ��֥ӻ1\*ҹ̘�옴��W���+�X�ô�Q��uJ�&ek$�����t.o>ɒՖq�[�Ms�j�d�9�.��F�JR��JT:3���.�}��c�jC[���R�Q����d�+��j��O�W069
��_ K�많�m
2��`n�����)��|�#}(�ju��¯D��̫ǟr}��dGq�%t��c��w��u�����sk�F9J��p�����#�J?%K�rB�s�nܖ+���W��.(�މ�C5��V�f� $)�_�s��-�B����,��x�W�NzXy\I�Y��Aޫ�ef$��(���$��\���������Tv
�����݇�Iq�C�<��;b�k�L�Xo����3R� Y�*�h}/2�pГ����#4�g�R��\�ӥep�9wWb�J.k]f�ڵ4Y�>u�BȪ�ƻ�i���p���bn�茡�d�j�&}%�j�\�o��\�F�4^귋6��3%j���u9�e�W[�v���]A�:T�L�!7����ϳs�����lN.����0r����Dk��#��RC,��f�;sz��`��sV
f���"�9l4�X�����ű��JR��]+���ڝ�vH��y��.l�owmU���"�J�%��o+/v������L�յ�E�_\k��)�]k�άaw��)%����YQS9���RI0佺�x���v���ۧ�/����#gM�.��&L��(r�ՙ��{��X;t�h���g]���+'l8힕9�Ƶꐍ��(hm*;��qn-��\��ՏR�ۅ����YT��ڷ;N^vlX&lFN������h��̫ɦ��;�R�;G�쩌s��c��[j݃yWmk��d�0�A�qo�b|o�.���]iяE����ڣč�$�u�i�yҙ�rQR���nw�+d�ݡ
��e86eK��4�m��I]�J�S�k.Ԣk��>֥�E�80���EZ��36gR�V��m�Z��v.a�(�ŽH;���klP�Cg �[+'�28b��:�n˂���'��w��"4�6��\����O�,޳�*�7�e���lR����XN���7���R6c16ad�ۥ�qV�W�>�8?����a�Z��]�Ό�oV�t�l��jB�P=v��H��	.��|��{WN����Vk��6[6H{C6�5cA�����x+�ʏ.eH�g25}��)��'+3b�o:����.�|m��ӍJs�Z�l�kjS��O�ǳP��j�d���R�;������׬
�{�'�R���r8.���Vo[���Z�m2[�B�����0.���k7)����qU�Yӱ�Kؾt*i����c\���]MA�pae�}]zn>]ձ5r�t���ŭ��_����:�^�ߕ�]��E{�棫w�3 ����D�}QL��6�'It:(l��|�>{��[k�i�U�WƳ&�����F�]���zk�o�8��-oY��˹�m-�\�"�|�R���u��[�%A�ޚ4��o:Uj�z�!qw1�N]zs�J�R�[�q�щ�������a��v'u����|)r�gRt��֥���k�.�Q �t�����GF�L�h�w}
	N�M�TT�nṭkj�I�/z�V@��T�����]7 ���j�,��v;��D8��V���X� �G9��trtޥ�e��K㛳�bA�̊��Ɗw	B��ȳ
��`�{#/�P�wn��w;��wNS��e�Dt)`4!�$�8E#���+q֐`��-��&m�w�����
��,:k����\�Z��.��w�k�X)0��˵�}�>�aM��x�qY\���r�40���mY!u�6Ă��U�z�{�P�ؼ�v@�R2�mene�&�s8r竨F�-�µM���6����:�C�TԳR'}+��-��W�J��$�ϖ�r��Yit��N#f����K N��Rlɐ'��dOG=�P����5����ާ�nԨ�-�;9s�qf7���+2�*0):�7�*nÛ�٥�%!0cߦ]�y԰|BX�E��S}�f�a[5}�耤;a�M��mp�˲4��l`�s]T�F��/���(� �Z�r(��J �ĥ��Z
��(R���ZZ����(��iZ�)��h

B�B������*�J)�)�B� ��(����()���`��(��J�((H����bR����b �&�J&b\�)R�
���,���(" (����r*2�p��������c1rR��)�iJX�
)��Z�)
����#"���0���2*��j�i2�$(��J�*_P+�fIf�ֹ���2ޮ)�
�{��Ce��/�%��M�X�	�����i�+j��q�o]�j�w5�Id���Y_��S��WuLq?�-!��w�5^Wv���[[R<��L�Ekn�4�eD3��a�C+����^P?Dp��Y�H�-�ϡU\k��M��K��xR�#�/��M��_ڝ ���,F�7�b���˃G	�k�X��:V�25Н8�iWѺ���z�H��__�򙇦.98���������8�&�A��u����(�Y˚ʒ�sޠ����������U�.���I���j��Gj�#�W:�U��Ot�<+�UsXo�@1xa�1ح.'�y��T�Y����O�Ԥ�oJ+[��)G7�w(�,�Vg��:!��TX:�1��F#�Χ��uŬuU���I�A�9rs�V_��w]Hۈ��N�FqtW?�#^��i��E�κ|'���Atv��TM����M�c���9��j���P�k���N����u�M.?:֠񚝱�2�z� ��J�J:P�-��9He�ϴ��վ�B๶^��JY0�;`��V��~���З�Z��7�/(u��݉Pf�aQ:�D|�fl�(lT�a��F�X�PI��Ś�����$m�=��7�7�eG\�N*�ouJ�g��+·.Z6�N�w�R��swZ ��n�����}��f�ȵ�0�ٻ��j�0_��q�&��?:�g):���X����<�ê2X��!E�F�ܚLc����B�[v��D��S���:��U��e�N��������N~Y��ր��XT�c95p	@@�bQ12�u�p�K��pF���V�9t��`D���]�໌��J�˰=��h��>�!\Y�;Xc+6�߼2��)o�ez��d�2�ؽ�l�^�q��<�**���Q_%�Gx����=�����{ҸјS��N����8�7�����#�=�x�e{�`O`�cn�*�J���0�<�ja��]ӛ�y�y���i^Mb�(-5�.DrwhƳ�'��z��]猺��T.�M�5]�����X��ncSz	���n�1S��o�I�ݖ��������0��q���a얡���c�9=������C	��q�9��Zt�0��@
�uZ2��^��M�Hյ�3I�2k�))_8wu"�s4�,!)�ы ��sQ [;Y����'���Z/��
�q�f0�u=�#��)��9O���	Ҽyu	pf��\�0	�*�Ɣ�a�R��:&uN�Et��+�҃��8j����͚��ݥ	>	CEAP-�����=|�^9]�Y7:��־�Ɲ!�քI��s����4ے$�<��{��;�v�ՏƓ4�k)߮�xj��*�B2=Y�@n�qw��W+�+�2JÈ�p��aY|cq�p��jh�t�i��N�Z^�P�σ�c����s˴���&s���H��Eal�yү��(p��� ��e n�J�5O3iԫ�P���B,8�tū�T�>��&�k�>�������j��Z��,B�!b1�T�{�%M��j���V�z�*�m�t|�����R��{M��#ۘ�p�����c�eG���!n�����V���P'�i7O2���W�_\Uçq���&��69U��\�%(�ݍ%�tGg����L� ��U
����b>�"�9]ώ܂t�����jw1F�qΈh����&�@�uV"iL��sG����0S�{Nw��̵ҟ�T�M�֤oj.D�S]n�f8C�����q\H�sTp�J�Ά�L� ��I7Sz��v�!�ǡ�����Z��0�td���F�
��]�&��t�Z�93Ɩ�O)�jӕ��t�����j��Gi+v�4:Z��ʦ��ֹ�r!��Sd=����z���@���Rx�%�Nw	2e��1���{z =8em9�M7u�%)Jv*���E��e�������jd�{�I(���N�'il�m�<�$łʳB��z��/���h��e�%��B53tZ����@s�ǟud���9���Y���B���Ϳ:��X�J��Z�3Xg�Λ]�C���ʥs<����(W]Ԉ�,��l&ne�(��M���sWx�ǯ�(0@�� V;��N�#�K�}HCG"�������Q�~�eU�ur�����ș�`��Ơf�=��=�=�x�k�d衬�j���zP��*#��1��Q?m�˩2Ӽ�>���\�P��`r���M����N�0���}Y<#v��b��`����v�T���RA��)���e.�tEmuV}f�Y5��Tb�LE�)��u��L���:��ӵu�,�X���vZ>�4!�M�B�g�ت,B���.�kw�#\L!����z
�C���(���{.;��+m�ꃦt�'g�=�Fȓ�+)!W�b?d���� G���*��E���F����'��=���a2;Y�T5YB�+��FM.��Ì���WBlH�mD���J��`m�ͺSiʳ�1�i��r"<�-{D�gy7o�>���Vgk9�u��>|��]jr1��b�.}\s�s.WHb��Dþ��%>�,��|(��f�BI��$�����̔ff�Qe"�.跩0�rfe]�k�[�dJ���}�u���96�x�F_��ѤH"3��=S 9�I���]��7'#����=r]�
��}���b�m�ω�)�X�M���ݳB��F�I�ZK�G
������"<�O+��\#�9�����~'�Z��A1��a�Њ���;4QYJ��=R+Yfx]�t}��BYu�3W�d�J�1pT�Q�2^@r�כ��#���o�y�U��VP6'5T��y�Y���u®�}���ݜ4���泭��z�z>���������<��"�1�?v�TqX�����]�Ԧ4t�t�К�bn-��%*��O�]��\�F�e#m��^��b8>>}ů\S�z�1z�&|����ګ�%Ύ�Z��:�@f��3�ȫ24�⌋:H�#}�g����#޳����;b{.a�>�'��]���}s*���WT����Mp����D�8����6���'�����&f4Lh���K���	��Zi��C��^_HE��o�d�='R�X�؞�FX����0v��+�E��('#6�
s\���n���t��і���n:��zr��� �6���Z���q��˷Bmfty:b��Es�|�(�O�ԷԂ�s.jF�d㧱,m�h��p�mΈ�uݻ�6��IId�e���23h
�|-��@K�uPb/d���<��Z{.�Z���i��Rb��3���;~�.�_lY&��q�񍟧�#�Ȳ4x��Hh�.�Db��9����Nf����<��p���j���V��h$�L�'�������0�^��t�y�Y�=Mu(p�;����2������Ͳ�h0��@b��yj_*�C�YԺJFS�ڰ`W)��N���Su񯜱��=v��FY,}��V.J4_x��!�����b�<�By� C�E��Nd@�B*#�1�W���(js�OF6���.�Г�*�����eG���1�(z:I��8�������w��e�&�y��a:�\��Y�����!/q@=��t�u���tq�v_���M��JC����u~-#�������[j2K|��� �P
�Q�jg�&j ��%m`�)��1��Ƕ���p7��
����ͪ��y�E� k_T6�b�3�L#�G%���c�ܷN��~�Q�+Žp�IF�-B�yR�;�gqي�_r���T�,�,��\�"�o1�[����>�}a���	����ȳ�P�Ndt	�f�ԒfǶ�z��	eI2ީ�wx���KV);��|p�YQ=�W.fEW�05͈�3׶�;�
�"�w"9L��C3Z��g�,�k�#�omNs۰�/_̚�y.�{g��6w�0E
�x馽�皶�����5��}xMf|��F�#�'��Օb��JfMHv������M�Nc���fySMA(`9q�hW����g��O��T�S���g>�U))Lj������6�wQq;�EWat}��V Ox�@��="��[���#�˧�֮JL�}���W�s���A>ȵl��0���U��=3�b�;J��2��,81H��]]��9�,:K�<�������fs�ࢹ��Cj�Y&��c�JU�H�W	�Q�k��5;�ܘq��I����P�H(V��2�:�9L_G�gIHx�U��%�]����t�^X�Z��k�Z폮Hf;Pڸ|�1l	qڨUHr�.��x��`X/�T��W]Ar���
��s�hƲ,�˪�z�ݶA}|�s� �k&R�ìÔ>���Jd�N��gw�_�?�}.����P�Vv�ge����,��r��j���Y���u�\Jz'6㳝	v�}��#��<�E
D/�m/��!D��"v�:�`��6���pљ��3S�r��2�)s��DLf��ӌ�'a���Ǻ(7\�j��Luȉ��]��X�|�s���f������^�{ d���tGc�M)������Z����"�-�]�в�j^��E��]!7��:!��^Vp���uV"j�(WT��a3�/9�>ݒ�.�p+�h�q�-r�ep�tq1{˭ѿ���Ys���VP��"�\��Ff9�L�І�i�G���W��ҩ鹆$P��b�ei��R��Rb�N̖�F>
���/2�vSSf{���u�n���{�g�Z�],�^��Z��uGl��N�GB,3I�M�ݲ{�3�>�GW�h粫�H}\���W���~�s�n:�}��lh�5e������{j>}�xzK�.z��!~�*b-W�Ucn������,w���]s���,ڨ*SWx���{޽�/��wV�&�t8%�7��h�S�ۜ-���~�e��uW.�����G��Yau�pʍD��z ���:�bs�#��S��_�Vq������8J�Hob���g�^tc��OU%���,���%+���C��}YlR[^��i�Y��_d�6e�ղU�K�d�I,;#=X���~��O�eFݔ��=`h� �ʅ�6��Y������+ϏWMC��׻��|��6�ɎI2��vD�1%�BM�iԡ�[|O(��a�t�cׁ	h������1���w-'���܍Q^R��1wNl��x[x迪g�Tm*��!�5��Wء�')�ȧ\u�;i�
:&��uh5.���4h�q����[JCuA��]y&����w��uKp�lź���^���7��}v����d��#ĕTW�~���2��ɗt�n��_3�D��9Z�b�-<�gea�!ǎ�zn!��g�~��:L� ��0�K���Nb����*37,5�A��t�\M��{��sv�N@�x�E�;�F� �Ϻ�$�g�P�{��F��=앗�`��h���Êtـ+qq�`���Aˇwl�D�xj[ZΈٗ�r��o32Dla!�o���)�2�t���<>�]L ��(�c*�
�(s�'o�hSk�j�z%�*N�	�j���:��NGm �#R�X}S�G%L��{�'+'#a�uD�Ƒ�X�_Xc�����a���ӥ�k��ˮ�{/��<�����Q���+r�-� b�nX^42�.��c����M�������k���\�4��Zd^f�w��m�8������0�vrC�P� ���m�9')ࠉ�3I��=|��@��0��}C����S�����5�R����jl�R��^�bh��ya��J��g��O$���|��6侇{Y���0�nV^S�֋�;��qL���e�ʴ'ru(L�=U��Tq�a�\�F�Qb6�۱|^����nX�?'Z��l��]9���e���0[��d���l�vڿ�L���Z�s���/j��`��0��ԥ�~����Q3�{+Gx5[X��.0����.����dڭ�]�+�����=P���lK��˅t��v�3$Gqb���T����H��<�c�L��ϯ���P��]�2��:|����gt�d�h�%
�G��ų ���E��5��рq�̐���܁7b�W�����\�����kI:]Y~9�^g��@��m�f�Y^ᴱ\��P��a�zs�?0�Bf�Lj�pwd�㠓���G]n�-�lE�Q\�ȵ���]r���?M�9�2��i������\�/�Q�P@��&�`��BA��Yu�?�K�mO��)��n�4�.9봎󑧯%���uP�+͇��}�uk��ђ�A�����Eϧ2J_bu�C���l��	�q#���n~��&������kC-��wj�W ްb�=��jl=���A�
�u��3�/:�Kf�Qx��^k"�]�b�<�����L�?�JX���}9�v�yD��MI�R��C�������]�Q���{ċ�V�k�6Q��<��D9�nV<$�E���L�y��{���)vɋ%]`��M���hn��T֎f�WbWt�N;�Wx��bYNW@�Gs���˫Z���$�����,:��q���x���/�0u�;�:�&s`�ҷ^P�e����4	W��t���i�	�3�l�l�\���JA�Gt����03j�h@�����hVa1�Z�-�y��GN�ڎ"-��]�7ZQʃ1���u�3�
���.kXҎ�b��ui�O5B�&b�Z�6� ���*�^g`M�M{�m"x�\�^�����s�=�0]�M��Yl�Z�R9�����}�䲦X։9�T�(��2�B=�g,����.�'�wNι�JG��1s�+ɣ�Mћ9�;J���I�ү��d=����;��J������G��0ݩ�y�z�Ȟ]<)e�9�rY�q���Ss^�t7CV@{����W�MJܔ�q3��ȓjV�qԏ��놮���Dq�L�C�̻}G���*����;�G6���l�-��y� �� sWtr�`�!�W%����?�o��֌����5�'w]���o6Ȕn����h��{����XKS��e��rZ /\��$U_6�n�)@ڣQ�C�a��њ������}ۑ�x �'
���F)j���ɽ�l>�x)W���@b�9C9>�x�P��El�`��+S�3!�y/7��.�`��NB�49�#�zvj�k��Ew��Q���r�*�/���i�؝\w����X��Y+8>���O
rvȮ;뜔�/d˕�=v�QiQ�6���-����z=v1��)�I��͠X��0ʾƈ�C�фt%KfS�w㱥�WU��ax��*�qB�<�ѷG!Q~�eB0��of1���z�c��������>�w��)�vC��m�l=-)Y�S2^
}Yń�o��5W@��Z�8f��6�{j�˩�:MX��J�0��
?t�6���2ɜ�{�j�댰� �a�pH�����^^[}]ip|�_���9��Q'�
�q�2��î�d����t�R�w"���\�?-��O'<�t��Q���S�y�*���bVq�KK���(i�:���5�6���2�ci��7Q�l����֙�;�D&�L�r���A>O��7S4Kۦov`mb�p�u(w[�Z�l�-��pG��d���e�7Fjח�H�ܶI�s�J����J���.(�7���Ã�Z�G:d۠�K�wH��7����:_r��$zV��;"���WgJu$:��B�����(���R����1(�,()������h(��rɤ�s0�
�()���2%���)ʲL�0�H�*���i����Ci���"���r "

)���(h��*j�%�h��0�j�)
J
i(�
rr���d����J��)���bhi"h�j,���¨*�����¢�&"���(�J)��3"X�̦���JZ*$�(�2"b�(��*"J	�j����ɢ����
jJ�j�0��
���&*(�*�C Ċ��0��&��j�*����������j("�!@UP�ܜ��!���Ә�3��eb�\�K�M��w��k�&'rN	�i' 7�,�G���ԧZ�q�P�n���Kml��Wt������xW��>�+_�]i:��p�G�dPd{���Zr~���0�亍BV������������%�`����u	}������K�FG^�ͯ�s������5��A��Q�F���!>�DH�9pe캍s�НO��c���Gp��:5�k������
���Ѭ<�z�2v��I�r�P�u���=�Q�Og��J����w������K��R��""�}�}	^ƹ�R���r:�e�c��u ��s�˼�@d=�����:����{��~�nJK�K���OF��Mԅ&��G���ΰ����^�E[�mk*����`��F�D1Q����7?A��{=��}��J��9϶C�2C��k~��F����9��u&I����sC�=A�y=���]F���j�5/��˹u�a'��Y���2{6�v�77��z8|G�.C�ìw�����u���w�gX�5�'��jN�>�o������h�N�`�%|y��h��jO\���1i���}��������x��b"D�c��f�f��_v)y�@!s�f��K�I�a�����ѣe�jK���zA�亍T��p�\��oFw�d�\�ߺ�y{�)������?Z��y��HP��>��(C�/��gڹ����<c�#�0���7���`�}�I��3P�O�~���O�j�ΰ�5��]Aֵ��2K�������?A���G~s��(yGk{^Z��d�;�����Wq�ϴ-��O�������1�)���7=K��ƿ{��N�B���u�p�X=��ny�Py���)��W�a���*�Gpj�d9�}��5����Y�d�}B���h��Xf�������#� �<��\��j_��4%�9/�����w�a��I�z�e�;?g�o�]Ϊ^��5'V��������SѬ7>GP��=��#�:��W�y8�&'�
3�*�䫵��� >����\�4��ŧ'�3�\�Q�~�O����>O��P�G��s\�{�/0�}�U?K��~�cqܻ�>K���|�v��j�z��>�� �"�w�2�G�U���&��̏I4a��Vd���.�Y��I��9�+��n�z
^�;�B��\k�J�>6ce��+���B��f=��EZ��Tt��u��Z0G�:�ͮ��Wٙ�$i7Kxo��^��*�\�*սΘ@YZ����aյ�%ol��F��>c����1~����w����;�4���p�>�~�a��.k�_k'#�5C�5s����䚏c�w��w	A���k�=�R?f���kQ���Gu�5��g���9��e��7��&K��|k�Zf?@�٬5/��=��C��{��������O�i2>��{��(>���������]\ֿ~��5�*z�qM͓�g�>c�HW�Ub��}� �~���^���c$�8�{{.��kC��}�I�^�:�������g��\��gu��''���>����E���H��s=��{�������=�s�\Ó�{�sz/�L�C�������%<�f�ܚ���0(
(<�g-B_bӑӬ���%�j�`�}�.���~�Zz���s��u�
�+������`~Y�2�r���>�{���O�rN}�?��伵>I�s�:��2�]F���:�.�Û�u�	�����WѸ��S��`�jky�P�s���|�5��`H����H��Dޯ}R��eL�/Dʍ�}���W<����MG<�݆����~�ǫ�>�R��4�����_�́�:������z��9�']����7�V��2��:�q�~��=�1#��>�������I�j��xb^��^y�����:�$8�5��������t��}:���{��j��u����y=A��s[��2A�ٮh����\�����ђdt����u�ϰ:�V��5:���������]��s\�_���o�>��=���>������� :��6K���\�9{���{�p�>Z����l:�	��{���I��5	_}��r:�V����pPx+����+������s�~F�����|�s��:�.�QØ��b��N�?A�J|��1׸=��K_h�]��.O��}�K������!�����{��%�e����o���sk����1_&���ݔ3���hl?�����s0wj?}���+�������\�G��ѩ5I_�P���k�~�P�y�9��~�Rv�ޓ`d5��OǞ��������or�Q}������ѿj��wnOR�t�K���u��n�e�����^fN�՜_��+���1�L�:���C�ǁ M.bn�s{2���/�ە�J���=��#�7�<cj��F$�4d�-zs�eD�P��X�|���f����@Z���:8^O�}���P����a�d�����觩r9�-�sRS�rc��7&�ʓ�2�Q�;���w�d�'Q��F�)���OS��Kۮ���C� ��*��`��j� �}�|��q�����}'�����_��:������9\��5��l{��Ky�w�O���.C����u9=�טnA���:��iC��j�a�7���|;�P�4e�g�{!t���!#������u���9�W�j?k���������%�_�u��O�!��u�Й>s^����}p�G��ϴ�~��@w�]�ܺ��.{�r5��C��x%P��{��{�ݾY��H�!��f�ԅsѼ��z�~�2�5֏��1y{��4;�K���ٞu����sP����sX}���=�Q��oO����G|���>�P��v9=�{(��FEO�&��>�#��O3�C_����&�=����0���]C�vu���3$)�<�O�u/־��g��R�r��y��%%9.]?��Q��NI�=�sC�X����z5���8EB�����I��`�?A�p���~���J:=�`�=N�jN�ʓ �|�k��ki�����'q�5�˩<3�u��9_b��uPd%�{�sk�0}����B׽�W�'U��T�Ķ���Q�/�����4C�g1|��滩
O������^��?_�1?[�S�j^��u>ɨԚ���f�*��(�{�/�;�N���u{.Ҁ�>����F�[2\̮@�U���do�7	T~��]�����}��a�uS��掠229/���y��z�pe��sA�wR< ˩u��}���3���t� ��.f���� }SL���uό�^
�������/�o����>�Qï���;��q�k|�j=��5��U<�/d����y��ב�������|�z���uQ�ju.k2B���#%�(�Of:��L�v���}8���|��.G�p�=�������3P�=�I��U���Ơ������2}��������B_��{����?A��`�;�$��k�u	k�v��s��G���*�dk�0'Z����Q7�Hl���-��X細�V�T��2�ȉQ�8<�:g��n��2ʣн��{�=��bTRp��݅��������z� ����m_]k*n2]cFE(�}�P�B��&3��.��__K��}B&)'2�2{fg1I�j���O����x�I�jܺ�s���+�J9�Pd{�_g����˾�~���r]��C�y}����nT���{���A�`��r����5'53�������Hc�m5޶�7�+��[׾u�p�KEǚǐu	o����|�� ��w���bw�o��j�7�K������]}���s���29/��S�rA�3��lE >� H�@Z�b�>&
[����`����y���4�}�3���u�����`r�hJ���&��X� �3o��?I��Z9�������:� �I��MT��I���#��]�
�\v��I����'���׮�ܺ�������s���� ��|�����CsԹ��`r�Ԕ��}�p�5��+*B���5���w�	��i�:��d��-f�ivw�T��Qo�_��������.t�q(�7�b�ٜ��xT
����ߟ��~�Ɲ�vq�~�o�g�m=��g��x��>r_'̭�w�'Fi��b��B�ܬx ��73OmRKa"cY�0���?P�,��^���DK�q
f��J�sT���	s�W��yxȋ�v�^��׌�5�+��;O���\����o��ᲀ�u_m�5I~|�����$�e����Ōoɬ�v���6���ʺ�G��ϖ�N����%����x���+ޒE��N��#[����ʲ�u��ukI:Z3�_]#^���
a�=�-b�F�p���꺈���Dj{���U�Ƥ�j��M���V�EdH�T�h�����8Ћ/rR�H&��Z�\T�)����S4����wI%.�fޛ����:�#���%����\����������Zs�)r�f����*�ٔ�z�Ҡp����ʁΞ����1�&aD�Ln*���j	+��}���̞t�w�s�v�V�L��*�<j8�5��9�2�柘ڋ}p��sl�� ���Q�F/�*���|[��8 0���w��u�I�����|�/��H�s���#%����[f�'�0��i�4#��|]m7�*�I�g�̪p�Nx`�M\C��2�,Mp�ɤF�,������5��}ptتS�|�g�"���iR�q�+G�j]׽tF�4(��|�3^X���ql���Mxxp��Bn��n�h�f&8����Dĭ�FGC�����̯5J�g�w���������Q��UM6�y� p�(UH�|���,���z�w��}l�}|��6n��s�ˁ���Y�غ�w��~�4��M��� :���I��G�Y��:�p���e
���ݪ�X��+�Om��:��W�9;�c5�̗���ߡ;�:�f�Ƈ"�'�Ou@�X�>Ei�x��U�tA�^�����&�ً���c�g?L��{�q��P[!�f���:�<��^͸��Q�M(D>�NK�a���ʚ��4��;Q���K=����;�D
J�A1�Ы���&�s���*k�[r������+,k��Sv
����_uX���J>��fD�wϜ(7�̬8�Cțy����j
A$�������ݗ����9����Q���u ^������N��.�f;�r����c������W��eWB=��e�E.�;B�E�Db\��W����A�_{l��0�,�ke���mep�7&6�'�\���+]I�������L���h{H<�b.�BF�ʀ��Yd�%<�퇗�
ϡ�۞���+GE�z�?r]�u�1�Q�^��lO|��T�ت���#O�}� Bg���t�����} <�LK�&�J�ɨQGج����(1Pm���t�NZ��ik�>��HfA`3�@��4sX���č)�Uk1xg�t��*BC>U��������,D���5Fb�'�̖��4Ä�a������p�If�ѽ0f �� s*�#_p�v�Uv�`ro�P�b�p�� ����t�p�`�fB���ϙ C__��	��nGL���[�����W�WA�x�\k�I�G ���zՃ�y���^�H��G���ܺT�z&�MX��:���ʕ�o\���\ffY��7�Q	G�Q��3�7Gl�Q��Ѵ$�q�u)�y�\��{��G%�S�f�>�Bu�gr)�!͇�WRU�]��aՎaj{�Q��rh�sT�\T�qW�E]rk�([��<#u���m>y�6���B��лE^$�� c0�%q�����o\���nc��2^@U�#(�0-�M}9:�.6V�S�wFQ���y�R�?���Nj�7U��_���N̛����ʹ�k��DGu�����MJ(Ve]{�Z�d�W�%���	���u�����ppײ��S�v�.�Ɵ�$��c����������W��,��别u�Af�yH]k\+�>���Z�rݳ�Ί���]*�����Z�3K�1A��f$lu�H��;�ݨWYMC�d�F.��*�d���t`��jR9���;%�5LCG����=�j�x|5(�e���W8|竢��\�|�7TZ�O��_�׽�4��N�(k=p���ڬ�q.�`�Ds�/�X�J)��{m�Q�Q�2�A?m�30�Ӟ��|U�&�YU'jM��)-����	���Jڶ���&��4�P�#+��:xcKµrzP�ǖw��1�Xۅ��)�O3���_/J:�3���Wc������C��=(I=��U!_ԕ؅f���°�^gg�E�����b�Ɣ~c��Ub��z,���uk3]NJQ�����9[��G��b.i	N���Ks���[�f+�7���nf���+�7�;nN�_L<- 񼝯'orڲn�Z���P�&���.K����?d���*@�@2���v��Jn;�U���N�q�?T�F:��w��q++��%G�*��F���t��2�*ʝXb|��y����8����~��t��9��{�!mOn��I�, �� �{�	��7Z��T��v>�uƪ���j�Q�{��sv�N@����e��F� �i���G��V��W`�L�u��!:�W��<"���ò"S��ZR+��0&���=t�m<��]��TNt%���$|\h��j!R3�b�*�˨W�_(>�S��p���Y�w�$j�W�LsV��yO-ʼ'=T9�KW:N�v���t��"�g���p���C���sf��ms$ˁ�5qԫ�d���d�X� W��'QQ; ��>/**WV��0�N��۲���q��
T!�-MUɸ��&X\#"�g�=,��������kw���fR�*`2`���_��YH�c�ܨW�N�ND.t���m�{v/�/fr����ix��q���o:z�h�_F���-���>�f��K��5�z���O۴YCQ�+�߭h�C]�5���#eOu{*5+髵�I%�,���}\�ru����7��;B�+���l�L���.˚%��;]q&�P���F	����>���shk��CWa���ъҢ��K��F/mע8�3��ﵴ�����\Z±�|bA��&2�hQ�E�������/��y��>^�uL�|s9�e�MQ�&�����]<+�m,9�K*�!^��2�G�P�����Fk�h���bo?T�r.�8U\��u�鿛��{�S��R�va� .sѥ9t�;���Zq��Ah�$b<��yLG_Ϋ���/�]-���'N�<]����w���'@gp�Y�6�cd�0�k��@�ON��v��p�����ȅ[|@6LJ:	;i��IEB�}��ޝ�U�Y�d�g�	��[�s����3����sl�`f�4�-wE�8�T{�6�l.�P�4
J~���}M�ƾr��]�w��=-T��Iȴ��Ho�����}��
�P�0�Έ	�X4��D��́҄bs�|��}��bLS΍�ס�F�����wx���p*����C��P�GI�<�2����]ɭ�����'����7W8Ġ�9s�r�������D�����F��+iч{��o*���tI0\KΕ�����u�Q��X�cD����o��y�9�oU�8�Q�����Qsj�*j4�oM,
J�!�G���]ӻ�婨���nE�ӏ���l�S���r��ǌӸ�qP}�ؕ�j�U�
U��>�ɰ�#\�j�zʯ7!Q�������\��8]�o�u�U@w���^E�F�RB�7��??�]1WR���zWOk�m4v)�Y����<��i�O��a���_�{��:�b��5g쪗��/ �ZuU�-�N���?2i��Æ���\�eļ����.�3��F �0���Fj���(4v�/�T�!͗�����r�ur�Q����ki3�I����k��a�'�9� o���H#wA�^I�L��y�gJ^�����9��.�E�d�i��n����MA�Oy�k$�`��Fw���|��� v.�6y�6NC����&�E:�K�樍]��:K��:�\T�}ث.��*F�|ڞ���;U6�!P\K,����}���a\�7y�!��rP�z#�Ɓ۵��SǙ&��=�ao�v����`�Q��t�рC8�7)�������5�/2�N���7�K�G���G�� ��p�*]��n�)�S|��\C��q�NNWP*1�V��79ۨ�̖�9���Kw�.�{i�>��d�rr�4�r�~nm��Ml�v��\�nLR�D���5l˖�Jkf'�Ӌ�Kb�i .����M>�E���ݮ�0S�G�D���cJ��|u��)"68��s�s���鱑��&(�yܳ//���q����Vlά��חD�e�>�%굸��bB�L�q��e
�ì�w�k,�V�n�W�,�������(��f�E�]�ښ4f:MS_���
=v_+��:���)WT��C,�L��c�A�~G���}]������ʛ4�A�H��u�ի�OkA�x�;�y4:B]�[�������I��a)�ǰ���Ǘ7%'X���;�u�_nr�bv�QZT�t�6�ٌ��m�*��yX��z��E���b�Qټ�ι��M�I��	�>��6�%U�"�L��RܛhK)Aj5�G(��0[�FJ�Q��)K:[�;@vKxZ�!��K�p�|s7k�)���y �gc�k��D�om:M>"�'��.'g�cz�-��Ʒ��4��v^G,�wg�m	�P�c2����_���	Q�(R�Ҡ�Q�KY���X4f�<�pn���<jsy�����[�V޻� �����;5SqP/NS�a���8^%ٷ������hZJ�����;�/N��P)�fKrHF���6=��S��qbn@�T&<4oU�tnn>���v�����c��w�p��.��K�lwZGMroN�O�-� �2�P��)C�ԙ��f��q1)�XtÒ�ЮvM�֙�P+h��5�0
�o=VjuL���/�+��sy�n��+{��/����YZ+pn9��+co$��q�(��ӬF�R��z�$�F3ǳ�]C Ȍ�3�I� УS���e�b���˜z�\���:L6'ٯ��a[��Z�L�̝k���x�X��w[Vی�Ɯ����: !��̚��~�M�.�7�@S!����Bq޲][}�㠻�ۘ+'1I@�܆���*�ݡ���k�iK�|%1n$�Z�mui7������42�{�$g�vc֮�n��I���G��:�w9�е��ӣ��
ݕЄ�tg�n\6'e3��yH0l�/���%׀+�m��PP)\�Vّ�����;�]����pM8SU!�����w�ͻ�2��%ڭ��]�2�[ދ�v��m:���X�Tҡ�����.NTA�����f���-���y&�*� ��3������2��;D��Lu��f���ɲ��b�[�2%�yb8��c���{%G#�̾'a�Rܻn�Ej2��V��腶v�\��&������[P�/�}��c+��o;���-[K�Nr�^i&.:	ܡ�sn��)��<}r3�;�R�kY��t�7�x��6�k��\�^�Y������Ґlne�(
_� P���-a��8�DLUSS4�14FFL�A0�DQE$SDSP�T�U)MLUe�MQE�E4D�PL�SVFf�2E!L�D̕I0�UYdQ0SCT�MEEDQ4QMEE6X�QTEIQ4T�TQUU$UEUDe��aNQA2PLU�dSU1E,ES1TQ9SLT�PD�QU�ST�2DTD5UQ0EDTAYeUE�BVa�$UDL�Pe�FMe5DUTTYeDL�RD�AT�31TM4UE��@� 3T�J�më��q�!��ލ�uiw>���v3K��]g&�:N��{�F���WF��$u،�Rr'&��}��}_+~L���a�d�lK���P]B�/�.��ƣ/2��+$�,,�F����]��?T�r,8�ٍdY�cA�ΕBc$�C�ޘ3
�J��'�Ym�nCs6'^�O������p��p�9O��t�=�#��'P�8�I�=8�s��ł�;t�G�>��X���9H��D6C��u�zê�Jd�60i�9���6��ִj�) ����+N�)��-G.�Fۘ�Ys���`9ROj.�Ї����tx�j:w�[�bE|�1]���F���1\��G��K���ٳ��;$s.#1�:�z��L&h���}f����^����b{�A�֡0���Yշ�{��ܑ��S-�`I�jb'��U ��,���Ln���?�ָW�@�)Vkή�^<|#V�4x>ULE�t��s��Bs:�dE�NTa27f�F�ޣZ�E���
��˶o����󥣛]L C�k橈h�WQ=o����]GO��!ߧ�^ffέHl�su�P�9y~nc��z���蓣|�x9�j}��4b��]��u��u��r��^>Iv�NXWXcv4��������ە����B��&̕9���w3�7�35��M�%*��3^�Wwq�|S{e��Nrt���a��ݚ������������_uFieE���͔��'Mp"{\<U5̲vg�W�57�#k05j9�mZ�U�{������#i`�O�&Y��QɃ����JWU�چ�Sq��~���K�+]m������5x��#���*
l3hF�.�)\��A����7���`��f���DŤ!�g��u��"�Ʈʔh@�~L���tҐ�G»��n�ͯR=N�>�n
Yb2U���&��@=�n�znVW���IZg�!�x�&^��W�v�>��o��/в�'��W�~EK��s��n9��{�#m;���6J��Hz\�xnN���#�Npc���
ꮨGi��UX\r)5q ��B0��p���ԋ�wV�(5j��)ڇ���4,A����*�P)�p8.5���dJvٌ&��C1b-Ҷ&�c����w��ި�Q�z��b�$x�戨Ƣ#=O�xdç(>���~(�XrEEI��Q�����ɌD�
��R�p�Gn�U=FY�GG�l�4�G��_W>��`�����V`
���mHq�z�m+����Qřz)Lv�\-����{�_��At�v��Wm��1�1��w��}%+����lF��f'^O:�G'`��)�d�9dXfkOU�|� 3fu��C��/�����I�;|9�o2g���������W�~���A�;�~�IS%�r�ׂ��%:���(��������E}+�����K��Ռ��k��7�C�y屉��8�健�SC.��Y=Q ����&;N�OEכl��37Thw�.��j�MۦY�Q��bo 9��p�u��z{�3I�'ny.ܾ�1�f�ñ��W�u�:�q:sJe�ڿ��=1|�W2�9���
qt�����|���ų7�PV��(9�jY��O���/���{�x.��އ�����.gy�K�91CQwb�A�+���f�a��@1a�\�cj6�^�n�sAb��W�n�2��}�m������g��:��a|N
���-6o׬��b#+����dL:��/�)�1nuC�b9��c:!V_���m$�#�0xz���>�:��&/��ʃe�̮t��i�����3�KT�⭾
^j�^ۺq�v�oB����ǦS�a�Y��X��G��c����lN�Nh��*x����Cw���$�z��ڍId�*��1r&�sJ8�ĩ�*��tmV`#u߻������L��$߫o�xɽ�y�j�U ��wgT��\53���CggT���5!2	jf����\WEZ�Ȳó*Qf�h\�(���J����R����������[bS��n+3��� �b(�w/��Rg>�n�5�8`�z�"��:F��4F*zn��s�j��q���(���@y]��D�E�B.�;�7}uINM����4����,n}�	��޺:n�~_>48�(t��-&�)�xv����G!�qe�'�-p�~�G���Rͨ#�&��.�1a����h�~�vh����u�w����d<�|YY���#��z��*5#Q�	T95ۮ�L���@�M���P�������j�wFQk�{o_�-�q�+������A%2h�~`O`�c5��.�xpe��Wt�d�i�Q�c�0K/O��ȷ�:�S{ag'v�g���M�5U���̈́fB��׼[]Bש�V�&�ҙ����~\%A��Du��b�6Pw��6��t������q7�vN����.��:�3���ƶ�3�������k�Z�a�% aD�Pg���� 4�޺�,�;Ο9�jhw�����u"�"�;�Uv}���*�v�OD�킰c���|g���!��� �J��.-��D�,��Y�ʛ��^���V�Lz���'�S��F�4��&��V(|(^�YLg�����/T�]��Ws�/�ɛ��x��r�V.�0�*L�%�hQΫ]�{Q=�r������\���|>�0��a�ΜB����'�H��c�"��u��~��&��[��o;�5�X|KC��%��<N����(�*�e��޹�h�� �%#��o/�|c3y�!wX����W��f�X�T�M�G��&�:<�	h�iz*׳�ʊ�u��+� �q߽�2�4�;~*��'%�^3������`������8!
���m�:S��(����ۨrp�
p��O+#"��pX�����f/�ᢠ��Iy���"��\o��%�B;sR����EܮQ�
I	�X��KF�v�����!��������6Na��SBF�J�PnwR
�a]�~A���p��p��c�;�]��~�Dc�c�rG�� ��	����Re�<�m�9�e�8��`���+2���.5�NR(������`�N�F㶤>}7�bЛx%�L�$�HRV��e3p7����u�7�s!�.q��ͦ�A�Q�irS�2�5��F�L7�:�U.U���xL4�ӳ�w�����*Ϛ�'��{\:�����HS�����Jk�.��0���.7[YF��hV�ۗۆcO-�4�f��GV�Y��ҝJ�)�Y�|h�}>ǜ���y6W!kR�� �1f囬:;�Xfuq̌�0rxڳ�+Nfv��g t�*��3�K�ﾈ�菪�����嗙0���U[�C�]:��(�_k�3V�n�.^��!�&o�r�pQ�p5�{�6������L�',	/ܪ�o�@���u�U%�[���OA=��{DR��]�7�.���ƻCE��ťT�\-t��1A�����
���U��4O�ǋ�o<��_Gv�~��-���f�0FΖ���[�u�b9]D����ق+(:��ςީ���Z�v��!�m=�SS6Q��'M vb&;\<U5̲bF3��}�Ы:�UvM\xo`G7�����0�k��	Ch����a�r`�*�~*�������w���>���뚙~�9�Il���GAG(W�7�n�Q���`��ᩏuF�~]���<��-s�����=Q�!ܦ{)��#8�.ʔh@�G��EG�!���u�ek�����x]#B9�Wb; kw�5���@y����ܬ�
,�v�J>�8-�sS�	��JN�?2��g���>����?aϣ��m���23�;���6J���\M����b��8�	7f<h�������jq�6���U�ӑ�ё��=��x��w���'�x�;mLU��ִ�{w����ݒ��Ф��]�K�o�R|4���N-t]59Zlm��\u�S�7���$�r.�8�dR��jĈ��/i)�lO^G������>ȫ�-����}&��b$G3������Rj�l�-�2����=`R��{H�B@�er��ΥOrmU�9�Dl�d�
`%_
�3�.Ʊup�N�0�H�i�c�5�G�)��ܝ=r��!^���=����|����*1��'�aq��P�	���=��N�v	�9��Iߖ������Y��y}Y\��p�Gl%S��O�ty�CI�b��nr�Dq9{�A� �ПК�C韷��K�XЯ�޺���ˠP�_���Zay��~�TНw��'}{�uk(W�N:�W�o�����7���健�SC����d�	��)I�8�����ҋ���˥[��ۗŢ�����	'U��:ѱ�X���۱�X,)Z�خ��Gil��ZX)����k}�׃�k��t��]�q�j�D���W2��ܕ��Mc���喽�:K����_�Ճe��5��p��K?_�i�1�_t��+�V.މS|r�7�|�ywD6�8�V7ew=�O��\h	/�*�/�{O�i�k�������^!�.�r����#�R5çbz�����퓣:��J���U�*Pj�Or�z�-������q�SBi6]*[���<M�bdW-Xy._1�'noN�%��8i<Q�u���g�+�U�4B]G�z ���5͎-Y+���IǪ�fN������D}'.$�X�p =��[N�	�&VS��Ky<:#{jxݖJW~�$��l�Y9W���lz��VK�Pꠄ\al�Q�y��r�j��pcr>U���v�?��N�5d��9���O�[�d>��ψ��|�:�n���y>a��p���j��9\uC{�]l�vk(�r�S��i4���߀��V]��&��ꡁ��{�����x�������&���)q�9���i�U{����Y��8 �����iO�]T�Ȧ��N���[�zH�<Ȭ�˔�2n-�H��i�,}{��J9�@ޯ�������y���"�h�
j	5�:|�ҽ*N��6P��t��n�鉗?p��B(tai4���1�=x�=K#S��lX\Ѩ�q��ɪA�<L0�M|���;����?.&�K�ARȨիM��1���C�ݧF�v�����H�^�UM6�x0X��(�[�=4:G�v��~`��P\�%�`��l��zW��_�	��ɢ��5V��H��f˽���zN�4��ö�˵�]�$�wFl
��i\�њk4%^Κ�*
�^��v,�j�w{�+ި�z������B^��U�mb��a���g^ݜ�'k��?�:���t=K��)z�=��Q\$�;3��]�bU�".�y{5V����U}���}C_���X���Œe�3�PrX��>��?W�Km��:�Uu~��щY����n�B�=�q��O��X��z}
��5|��ATtk��z��sA�0Z�(�ȵ��[�Hȱ�+n�As������d�ä�2��@�k�֫���K�[�İ�М��A��x���Pţ,�7Ο9����q}��e�!w����z�j3f���nZ���MsǷ��.U��Ka3)��ΖE�)��Ϝ����MW�k+���9& ��o�_u\�:ﲭ��(�8�d���.:�!�pv\,��S̾�y1�_K��qme���*�bp^�6�z+�0n�I�D��N�Ɨ���|�4�}���@"���y{�B����5Z��4�7d4���x�z�:�+�_�\Q�Vݿ>O� ix�~�T?j�u�����B���P��,u�P���^5X*��D���]�#(��3�㠩�{n�2����=�)�X���T����F3�r0���84����2K9_�;7R�ylrq=���Y�.�j��c������	A�,�>�3n���>�tt���D+H�Z�u�>�Vf�d������I9��}ƇR�X��O,ʝ��Y�t���a|A�omZ�P����.�0*�ڒ*΅�8s�`|�6�[�t	O��$�IKU*\����W�_����ܒ��;U�}�'K��nr�Nxi/h��.�R����\�� EМĝj �D�Z�+K�?.=��}_$�"���l�������V��'�&){����耠,{�
#�pfP��7���:���l�c�a�uS�&���6wi;��B�HεGK)T���5ʼc�a���af���un�����t�e(}��R&�۳F���p�*3eْda�pQ�ǺH�ܑ^:y���Pj<q�FSek�		����N��,2�`���LF��'td�t���`�E_����qa���T�B�O<8O�Ֆ.�b-k��[���fṊ52"�
'#�sJ�"�z�r骬I���\u
�)#f�0F��L��S
	���v��Db�]g����Eᩨ�ߨ("�~��ޗ�@<!�Vvb:r߉�F��+����x��7���b9擴Hj��_:�lEٌ�r��	B���~��G�TNA�@+��c�)��]�n�����]�r��`ʎ=������{M�Fٗ(�uW�I�������_���!ZT�|FI[���06{�u�c]�����j��7[����af.(����:��ok2vUtل2�CMތ9��u�������)%�9��U�
tt.ˍ	��{��h�X�J�,ўL�s�u���[��;o�sn��X��Oww�]�㢮$y���A^F�pִ�&��gs4�,�1���k��^õ���Q׶ݬ�|��M2E0BS����i k��g;7Ki���������Jw����x�'�
��� ��ݲ��y��I$��VwZ���V�VU�8��)k��I۱)C��:֪f�2�&1���Au�"bm�byĪ�Y"�ٶZ�ʝM��a�bF+��z霩�+ةG��Jo�4�b�볭� uy�ث��c���B������X��|�Yl�.7um�×�Ƹ��"X��qċ�w��`�����\��������������F�7+�P�<3]�yd��<��c����Z���t�6z�sPa2��2"5��=րf�ٻM4�׮�7�r�l���ŷ{Ά� ˗}��̓�4ɏ5'��������5�M�}A�j�\FG{t��};6鼐]�Ff����Ak�N��T�zVeŨmu,0Q�]ч:�wqW{R<�,��9M�.��6Ld4�Y����+�hm�1�9����R��>wһix䭚�*�p��sr��ϜS2���n���b��M%�d,�y�:�EWr[h��!WΟc]�7�oJF�����V���g����̣Y�(�sG[Q���ލ��r�cfm�Ǧ�,t��P@9H-Tv��VaMf�
�V�d6u��.Z�p7-��5���S+q\7ce���N��Q��S��f�N0ab��t1"�W��j�&Mj���JZq���u0��+(̼��L9<�i�dM4d{x�t�ƍ�uyݯ?�^�-��;��\�4o@��dƠ�.��+f�]�l%� �թ��x\J,��`۲�����h�hU��-�e���5�P�	F��V� /zfv���`R�������,)%#j���c̤�ݩh����%�j+M3[)S3��L�L&e�S�GhY���\��t0�qsY���ɍe������`��vv���9[����- PY�]J>�hE�T��"s���8�n��Mz2�1��h���n��{Y:�$(M�<a�`vd�*����v��[%��<��vUe����f�d���u�(���wͣ�*P����i����y��h��i��
�(��%�v�uG}ۺ�-7|�4�^x�d��X�0;!��^^��bf�Nw�l@dF�n$q�z��
������e�mֿ�D���wYJ���:{4	\���23\�%�]�4�F|��/i�-�6����  U
( �DQAQ^�%�EI@PD�3fdIR,CT�ERDITSIASTUP��5DQEKAQU-L�5T�,I��T4SDMM4Ԓ�fa4U4��DIADE4�UD%%4E�AQ��KMfefcUHTT�%U5AIAK0SE-AT�MP�1U5$�d3IE%DH�AEUS@a�15$�LQ�D�49T`ATP%%P�%4�@��Y��SYE�MR�U3UAT�a1Q@RR1D�D1EM4�ETEESAT��7�o�u�׊J�o���'��k6S=˩
�����	�ZD5ƶ �zfʻI�M��9]�g��KIU�7I�yvH��f�=_U}����_sbE�a�u�#��1���5+M��Я
�����𶗅=|�(*Ȣ� ��"-���k��9�d.��q�1�r��u��D��0��Qߢ�'��=(\��򻲎1����*��*��kw�#\L!��:��w��r��(�QCI+�
��U E��U����ţ��2�����xR����xy��b�@=7z�m�w;�m�"�܋���.4M� oK�,f#6R������{F�["�|\��I��'/D�@���oR�z�w�{���$���4�Iʇs�P�>���l�ԩ�f+&j��t�ַ�a���<���\1�*u-��4.�EI";*��/�/��\5᪙�.˕`b�Kf������P��%���,�5�OX���r�I¹��U=FY��ty��{]p�$~�����/t~�T�}S�5,������0�DON���Z$��������vc�Mf\!�m�MUɿ����4�
he�g��)1�u^>�:�t{V+���̾c~�N�A����r��Gu��%׼��P�B�u�4w{���Jz��|P@#%w�%���ES�)��-�n_�ֈ�(���-�D�[����Z2���!�wZjƆ�\��U"�)��!c���[p�W��}_|�ᾧ����?P?k#��cĎ���>G~JcE�a'w�:ѱ�X�κ�t��esgmR�U��vN�2�g/�T
������eԷИsb��m��^�\���]���lo�䧐�o7G],�Ƙ,�a�j]�����k��>'.k��r�1ޭ���w�蜧��C�1�P�a�&hO��\5�����$������<*(gf$�����]iIZ����S�q<�φ|�+")�ۦ���oeO��J��c~W��F�]���u��BpP�j�,T��-�1nu})��3��mu���k�3}O��۾�\N,oB��4I��Q�c��Fa�#�������9�ӟi�����3-S�ɘ���2N	�����75�hN�b~Ӡ��Ip���[K�ε�0�`a9�C��x��I�[
����+-��!�R��\��(	<|J~���;u��p�etl��	����(X|��G�uDd��S��!\��D��TPTv�=�޽m����4k���6�Ƃ�ݜ�>��I�o1���<[e�wn��qb�7�0ɭ������q�
dr����
b[3z4����oW:&�QL��i2fڼ�f�;V��JS7(No_9Wܒ��_�*↙׶3�����`��U��ﾈ�2bz�b��m`��=
���{(g|�wx���q���@G>�"yB�?F_���氦Y:�KL���Ȏn8�%z��P�V�9t���1��_&�@sN� �fMX���<nn�����\F=Jy�n��u�xtjF�/����-@t�,!`ZW�N�n�ә����W�U!ό_(/k\T�v���+��$����U,)�F����]��;�ˠ3uC/�,�xŇ
t<,y�0���߃;�W�vCn�7�1�-$�تż�)gY��S�&�K�;'{f��8x@aoX9ѯa��_=&��C����	�WW#�D#<�448�O�3S��/�6����[%�]V'1��P���2��1)�l����
�3϶/�p0r�����e��>s���9���ݠ���0�b�q�ug>#r�����������){��Dx �t�.�O:l��?c鸄�p����^�Jb��[[�J��z�ݹ�C�a���o����R7sѸ���+�Yd�r�e�����l.3�~N��́p-�-f�\��X��`,�x;�*�+�Y��b��@�:T[�����'��ѧ7gN�l�����>7��R퐋��X�e7�(�Jn�FxvSn��V��3����讧w%>F��<]��N��@�"�P����Ln��2���߾�����4#��"q�B����E�`
�Z9�e���_GC9�>ae; È�Fh'��/[Hy�s̬���5��0Qⴐw*����Wb�[^}5�]䇤��Gn
Q@���c��T:C2��������~�!	��K�p��l�+�^�:9=�<d=,�P5լŻ�r��,V';hԥ,��3y�B"���L���P�{���I�T<W`�-����)˨��9�|wS�8���eC�Ko;1b�T��#����3< a��IN�iw�'�Ɨu}I:H�s�8^V� ��ɀ��ls��v�uX"j�ԉ��4EtM hw���{N�=�o˩�R����dU��v�qv�47eAPx��L�z����Sn�9FG���W�xL4���J�^{R�nW�M������%���Ra����nb�����ϕ�HBZ����P>�c��|�<�&DN)�n_���a�.����p����c�5�����/ؾ�v��gF�M�����Y��4)ƺ=�n�6����b�"AKI�)5tZ�v&vuܠ�Q1�Z�(;b�b��a�Z5�H-Z��S;h��]�tM�򌫨ԳΚr$�x'D���5Շ)�C�c/#Q�Aȶ���);��]���a�o]m::�����9~�i3�9�m�W���������J^��jS����:���;��:�"xZ���Z�����Q1�M���9:��wK�4����j�������qS8�t��=�~7�]�P�)���p1D�|��B������/�(ƉXRэ��<�כړ�F���Q檁ͺ��,.�k��^��S;l[��51��9m�1�A�,�]�m��;,w]�:�K���P"a�Hcs{�N2�98��tcc�Cx�z�_=���Wˬ���6b
w۲�[j�w�C/�tU[
��N�R�qIR����8k1��m=����
3��F���BΪ���0�[Qyu��Eҥ�P�<�b�k�r�@M�v�ʦ��I��8�T4K�|���$��^���.��뀱���U���&�i`)�K;Q���v<�^UB#�>5�$C��q��������cJ�4������L݊��l���靯0<M�:L����u�j�e�%�論����}�	k*y�{})�A�wG:���sq�D)�Ȩ�����!>�	��k4v�c��K.�A�]e��]iԩ��G�Lj�H�9�G,�|��N�;k��+�|&�<���\�D)��.����}5+^,���\��:�K��N&�P�5l��W�J�x#� �ӓ��E63z�^j��٬��q<�j15Z�u�MG4ÿ�7��%:�����u�3�vr��*�/,�>�L]�ٗ���Y�w�>MQ���n5�6�J�.;qB+/a6��}�Z�P�ys��/'Mŕ�:l�͵��od�i�ln�OP�����mmTG,7_k�b��yQԴm�f��<��;�`��j_:ĺ���sO��G�e�6^pn�u����J�s�|���vL�7��F��ՉÙ���n�Q�uۧ��pwa�^r�Г�*$�eK3�7�*��\o\a��|(�M�t���۷�{՝gj)��ib�������r��П��,�N�j��W��Q��܇m������yD�UM�;�H��JżS[--G;��>�א��ڲO}�4�:B�*@�����kZF�iss;��Zh�	R�W*�s.��W%c�V�8�������gl�ѧ����u�(��-�lqg6�-��Q�����+u���n�8P�2��^iH�T��^��>�Q7`)�}�W������yW�%�}����Z�F�}��i�/[u�z55��3m(���o��߆	q������8Ӟ�o�������Ϲ�Wc"���Bڋ\�˶��_oA�^��Ǔ�7���&e���J��8R�	k]��3j��R�}��a�!��z�#�5��g���r����'����ZW��OtTE�2�S��B�fp�d����}�;xz�^���e��*���W����+��C2���z�h�7rr.����U%�;�Tܭɨ��_jG*�4�����k�*D:��i��u�����p�N�<�\�nMD��Q�����MQ �Nu�xz������/��]�7_k�'��e������_g�����$߰��*{�$e)N7���8f�8;I�V�7Q���g?��1w���5�z��/U�虙��^��;y��������M-4�G2\u,�YaHT֐z����[ć�x1���V�]gH�e�_:ގbz�BIԨ��t{6�ۑ�f�.�Y�޼��-)�'v�c+*�;5ɋ��]���v9W�g{cd��}G�:3চ��b�����ڷ%/q8�l��ڣN3�eA�)��=��H�nev��:�������k;�S/�|�5]����˳j�Lʚ:j��Y��G����D���laQ1ظWǚld:�֚��w�5!�󅭥���.�����˞�P�p�b��7�B�[P�`�͹R��UKV�Ov�s�sҳ
���*eY��Y(̪��)9[\r�v�����NgH����m_������X�B}�Yn�J��yʷ2�67w��ө^����{;\5���6�����@那h�ˬ��"�PV��W1����wETJZiJy|���q�o��t݋��6����E�KC���Y�����.�Z�j��-�r}��3���[��	��wG��U-��7��$�T��r���)&�;���o��'<��z)ҙ+n�8`H�H6���z���rTJ�x(�՗�6^�WnE��@�_N���g:]����+)'C�oGe�p�9�z��(�ڍ�ۡ��d���=݃'6z�5F���.Õ����@�C�,:���v��:�z�����}_}T��oq���y�dTtڔ�����O��ne�N��ĵOjѶa뱏q��Y-�aXxÿ���(Lu#�9�PX�K�<���+V�5ܹ�Ht�|��o�j9&&�q�Fk�'�و���#�te[ZF;�6��q�&����j�u59�M�ڈju��h��B�����"��b��sڮxjYs�yy�~K�|��u��ÚyNv���w��%�[v���*O��oEꋷ�o�%`ʌ�����R�_��֭7�W7ݕº�uq�cW��ގ���Ϛ�Zj_�o����o��j��kfu�+�r��j�)�Ƙ���m�毻.�syU��Y���j]��P���YUsu�T2��	+�H��io��*��Y����x�(�ւ�1V���:�ݕ��W�bo.O�_=�9���38i.�i���P�ߴ����YZ��#]�y![�#�mi�j����dU�86��匏�gR�s�����a9W�ؒ��}΃0<�;b�|]������.ʗ"���(��*$]`�Ӧ��<dԚ�8��j�ۤA���2��6p���p\)�a�]=�:�$���\UbT����X޶�qY�+�gV����h�-������Gs޺.�R2�<�p�㇆6�U�%0O,͉H.�ic���x(��A�n�c�e>,��1�L�����j��sq��fզ;�s�h����xБ�唚�'g�:`C�=��`u�D��-,֧���U�y��61̹�D.��4<�s{�wTu��j���\�����ڸe�w��ĩFx��9�R�C���͜b��Ims�j_d�n�Z�����}�0���;
�'&�j%v�5����`���\����Y�o=i�=��MƳV�]d�7��6�/�.ݦ�ȗ~;ٗ���ڔ�:o�{a��߬x�ټ�J��a�=��ۭ��j�����y[�)�_#��Ae˧�/���X�%E�
��><{mD��A��Z�r��#�f�uw��Z���L�ڙ�Zu��yd9��:�K�k�>�˥�����\��p�"�2�G7���k06�>�/rj��R�U�&�勇��a���k]Eg�$EnZ�@���t���Y���`mJ�rT�ζz��Ow!�L��b�㤧V�)gSGfqV���	Oo���a�x*���y$�d��սpͲ��.�9��f,�Ѵ����5�hf�Yħ���.&=��G՗}}Nv�֗=uΠ�JN��A۹��%L�����o���́�����݀�Y�htT�j]
��|;*��p�R�zamʇ��tn �m>y�9��������5L�����1�3^�pLI���XlJ�v�<R����V -�9%4*�-�DA��˄M��暵�y���ӣ��/{rܴ��c0��{��q�"Vm�Q&�C��^ �bUHtB���Ly3��ɩXJ��j�M�8�q&�qJ�ν�T��-�(�9�+xu�	�Ph�J1���:�{9�g'{s� �ܒ�d�w��t��1r?%<7̢�yύ�ٚ�[��N���𱺧N�{cL*B�׵Ι۝��d�'�΢y�M�w]Vɪ�D�}�e��=���U��,�Ѭ�hu|��(��6^�Y�Uu��`�b���&���o�$b]�L��<LJ��d��(�DM�8�ʮI�V�.emͱ������̬yi�v:.N����r[�DN�1�}-��or��	ݚm��-U�4�u);�J��t�ze���#�3x����F��;��	�{K�|���J�iۓ$J���D���[���&�.�r��妴������)&�FF��-���Y�յ�t~jn'Z8)�,S�$c'����K{2�a���S�Xl�k[���	�ߵ���6Vo巫A���jF��I�	ny]��Nt�������[�ڽ&�MSF���:�*�_sr�(ڭ#H��z�,���{�r�{�t�&9ue!�X�:�p7��r����ʬ���i2��{��1��̳�Z�m%�if�VQĭP���wAlu'p*��r6_g(0��H�*�+�)q�w}S���휍�۬�ݦP�y��n�q��s� ��M���iuӯ�2��M���e<2P�j'>��*Y@�x�c�\�$�4��u���D�S�����/�)B�kop��	[w�[�7�wE��]��7	gk������NW�*�"O�rae!��C�X�߳z7���Zr�e��Na*3�扯nYA�JV�c��B���E��]��=�o���u�,�$��g�U����%�K��wѺN��f�H�8��7��Ef��)p���_RTZ�p�4b�#��I<�[)�jώn��/kp����\i^��f2j�ٕ(>g��ʆ����V�1_�/�:vs��E>� �Uk�]�w.��̎���+���כ��﷟����3E1$ADLU��4D�R�҅��SM$EDAK4	I�	�Fa�@P�KUJ�3e�R�DEITU% D�-449M5BD$E�Ҕ�%ICELKMd�4QKAI2�TADA�M �P�PTI@RQQ%%NHQAM�deDES44M#@��@D�HP�%% S��-	A�A���%AddRĩJd�4�--!YSUQ4�%$M D�BRda4&Y5BRSE%4��Q"D%RQKQF`dP��ߺ��s��1;Ѩ�>A��|�]�����c6�uɦ��5��*�}�3�e�ǵ��E�V����ד������{7�����ױڵ�J�F�{i8��}Gj�3u8H7҄�ߦ:/�t���w���3�ί:?l��d�ɜ��4�t��wG��C"��n��ٵ���vo�,������p�����}��'�Q�gzN�J��ĵw�c��P\�KX��'z��`lls�����0u�fGwl��j���q��ʝp�OĽ��=���[���N^-
&����n�����Q�Mpz�SD��W�hy��OLFL���ڐ��/�>���m;P�zq�r���<��m�v�����}�*K����u3b���Ô������-��=k�5�m}n.a:J�XS�w�����mtf�ub�o`��	�}����Ʒ!=�Qm��uFx��x�p�o��N7�j��~8ƃ����8����k�W�w�x�n�镍���!)0+����C@�,lh��u:[ʎ�=*���#���O[H���(�91�!�2��i�?(W
>��ɽ���Wt7�4��|.�k����n�4��/I�"�b��k�2��5�H�'��-����)i�+��τ*�.�żx�FZ����菢8ڃ�Z�uU(<0�����Q�Σ��\����֤�g`z1�F`��s3=C��j�?u@�|5��3���؟�;]I�q<�:�f�̃�m6k���4ۍv�k�oTez�]ϝＥ߲+�pf.plR���#I�mZ�N�8G�pv�ʯ��Uo�Tk�fAG-�moV�Oӕ+�����y^���m��T^ջ����bp�܉u[��[.�h��??9��ww=�y��Q7�_	X2��c�jeฎo��j���-�HhU���d�8y1���Â��	�63�������D:��LM�l��K]кC*�>g�θ�$fG!�PU���TK�*o�uF�WJ��I�u�����{�)k�W��+���I��K�bT�Ȑ*%���p���\�E�%���-�GM�Gm��p��|�1������i�"nf�e���;�m�GB9��`0Ǟ�,�Á6q֝32�k0�0m�S\�y���(K�tom�9,	;�wSy��
-�G&%��˫�]ӻ�������Q9b��7���+�l�b-�{ 0ef=�k��8-b����2��3��������6������Y�52��֪�ky����6��X�P���٪)��:κ�w����+��%-(�{ͭ���ڋ|19oD�_t�+�w�.}A�/��Hl}|�c�n_u���!<��o]�L���j�8��J:�Mi=��a�`���rv$Қw|C322ej�b���93WkS�*9<�snk�B��B�4>ҩL�V��8�w:��(�Aן�j\�j�w:M�v �;�R���GX3Άڣ��blͳ�r�W=`/d���[R���ռ˦���䘯���+��p+��ҩ�ӆ,�w�Y-H��eĮɨ�ɍ�j�u4�Ú��m53��@; �#�]�mֵ���O�\���Dm-}��j7++�����r�\�`ZT�h�z^i�S[��zk�z�_M�ʆb6���g'Q{\�.�
�MMf�%�u��"DS� y�U�,����u o��*mH;�$Û�j:+���u;[I74��q1o�L+���Գ=�O�)y����}�zhvw�L�]�ܧ�:�R%X������vY�q�O**'%�Ҷ��/-{�e	2���nWj�}�E���\�3��/Gu��3����M�ߕP�:�5.����W��]��K�����/W[�ld:���oϯq����|Y��^Yj�;>��	Թ�a��nL$�>��Q;ڐS��bo&/h�Vx$KoA��qԯL��@�G|"�N��%ce�������_ɧ����]gq��S�j���J�N�e��+j$�W�L��1*V5��Z���OT�c��c�3i^v��Zҝ`�H�D��~yg�d7�G=���z �˟Dmw���O2�YSuσ9��ެ�m���TDfK�z�Η{LbS�<��G��+��g���o[�ζ�T:�J���0�KD=�䁱�Q=����sl�X�p�-����<�By��62�uNk�D)�]#F�`�fTڴɧ��m�N̸�[�;��Gsj��ö7��&�<Q��%S��Q�d= ��Q��m�ݭ����ܤ����P�bUg=��fd0rY�Ӻuԟ1��3H�5���k(~��ܧ�Z�n��jۃ5�v5"��r\䦽s#�vŲ&-�*��ێ�r�gPu+��F1�y���+s���^wQQ�+��W�f���}�k��]7��ɭ�u�K\�rL;�;�
�*G��k$gK3��o�W��Pݭ�{%�w5|����MQX��0mӼڣ�&㳸�u'�y;�d*��T/e���K�E��7V-�X�4�Y�[���c�Ikst�8ԡ�<gjʭxn���{?�-�\���T��3*��H���K&I}���vy�_�0�}�waf�v���gK�~����<��nzx������4�����߫$趤�[UyUۦ��7�͉���bX��|���79QS�:օ��c"=��v�ޜ�Wi�$��q���m�錎��%N�ӽ\j��*9�{�;o�q9[�<���$�1�'z��g��V�]E�]坎�ϟ�Pƶ�CA�v�w���n�&���'ϯ�d�ߌ�0N�f}�7�.��3���X[�^��m[0Ya��0�*s�W��Re�+��*����Ab�Ӕo6��V����RF {oo�d��>���#v�,G��r�t��&��W�35Ř7�nZ���rLsV	�M`TUZ�¶un^MgqM�"Fdo	-\��&�T<�7��)��&~���wH�BqҪ}���TE�yP�-���.RwF|ؾ����}I�vx�����0������)O.9�]��6��\�IE���˛�Q0"�!"*omm��n�Ar���_t;k;�OtT[c)��:�Ec����e�I���S-�+]�G��.:�I3����ҫ�FY��}Һ����i#O僁��..����ўq��O���7rzsF�*�n�%r��ں���V|��勽�7�9Zjvӿ;�8)z5�i�8��5�I�M�>
�5��൰�����>Ax��k@IԹ圻撼�R�-��UZ���ӄk��N�]�:E-�q6��|T̵Ӷ��yʯ��N�������/jݥ/o�[�uNve=ӽN�+>�#"�y-%�<��N`]����V��5������9��g��rc���z��oD�nz�io� ��oRBԷs(����*6Dh8�qc��6P��;�f#x��ɔ��ܹ�����ˉlW�a�u��]�!:�9'ڪ'�-�( �+G!���{$��2�w-z�5����>��p�c,*��1P�ʕ<��腞���͗u8Ig��ܨ�w�[�M�[=�_6�t�#c2�\�;�s���Ji�Ó�}'u�U�b��0s����^J�uzX� j��ȜLN�ZM�+��B�$�,j�v���gQ݊�����C��C�W��{��.�R}������?p�����m>�������Z�tv����E�����5Z¬r[S*VµK[��p�_���|�{pV*�C��fx]��B��K�[�D��������KMD)O/�[c��o�B�c�B�AتX�OB�X9�A)�<���G]���zJ�������#
�*�s��,��r��4�S�oϻn�tb���/E�ٝs��Y׭Uj�p&�����ۚ�.��� O�/��n)���lv��,�ؗp��:��q�
�;�R�Q�@ﮆ=���oZ�X�=u�%I=�0R�_ex�`�o_oJ�2'�l�I��b�T�
��f��xd��)M��ts ��T���E&�3�c��>'GYr%j��<8���o�h��vJ�-^����[�Z�(V�ّd%V��:G���o{�I��I�����
�o8�S7����eW�:=�>~�i��b�q�¸�N����{9k�S��*�D��k��PK,������j���MB�Sq������%Ń{۰�3˺���u�س��2�wu���n%ױI�{K\9u*ﲦH�I��.��4�.��mTr�z�E=����W�KF��w�͌����OF���e�kRތ\�}G��w�h�}�fQ~���nr��M�5]lM�.����p�oCZ��Sa:��	�����˳��fW�\�|���p�R��a�J�'T󗞪ղ�J_L�-�SR�r���¯�$2�B�dc�N�甧��`��s��Е��j�6+7��>�u�o�7���m���ރ��w.�)�X�s ��eA[�R�������w�}�o;vǮ�NOC��)��2K�7>*��!'�%%J��rz�F�@ubu�}�Ae��Z��2!���K���bP�=%j	v�r�2��8<��\5�Jϩ��T�]-y�:aw��)+m85�=��v3+�¤=(�C�%��V�>��g �c$�3���e>��������j{�m�	u��9��w6j�}��th��OW-�GQNs�w����'uFQ��ݵ�?�
�[gg�j��w�PR��:[˄��ȍq�Qm��uIX���ޓ��-������3���b�̧�
�\�w<O����<չ	le|꜠'S�4��[�I�<�����w�*㝬�KxmBM+�������o!�;�ٮ�R���T�z钠f���SQ+rwy��v�K��&�;��c4���.��A�業5�z<���l�וo�y�mDo=w	�1Wr�U.�B��ܚ-���H_�t�P���R�şo���eWd^�J/#6�J����Ԡ�E.\��V�p�C�jʨ׆�#X�������y�E��/w	��=�mf�`��*�ʷq���q�c�:��>�vo+���
����rq���m9����|;i�WY�~�w�tML屧�͗��a��Ab�����3Y���6�|OQc���^�G�6����Z�m\���邷���=�t��'�-���Y�U��Ԯ�9��UT����Μ���=֭�z�v4F�����{���;��J7�/�8�� �@f�Mu��hm�\,l��.nJbOQ[p��nr��:��ËM������Pwi;�nS=/q�)lv�Չ���"�쨂�Aޯ��WӪ�p�0�+�7������霮��jJ���g�ړ�W=:�z���/��t����y�o�\T�λ�q�D�Xj�JgHx�m=N�ۣ5�|fUbY�~s*�z����hmu�Q���J<��J��y��p�\F8{P�{m��ZO�Cv���k�bEF^8�-����N���R٥)�<kq���*��XhG>Wj����D��
���������+��N_u�X�s��E}m��:�Un"m(X��K�C�����-k����\v�i[9�ͥ6���%���&]��r�z�ϫ��.�ǟ�yًw�'���{(�D�щx6�Z�[��m�������p�Ԏ�<���5/b��<�_���ti��BPL�7�6���ȃd�زe �a��#2��m�&�}���֟e�R;h�]7mìrLs4a�Yڒu2
��1v���)IW+�Ũp�e��+x��s��k���X�*V�bn�D��:��K]+�R���=�2 �TjR�6"Ɋ�<����F������T��廼�:�5��I�6���*�u��G�u)b�]���E�j�t�ۄ��׶.��JTn���Yg0�/�as���.nZ��3_>[���Ё×�$΁��nJB
O��n��qJ:�Kݭ��:@��-�k����`�I�v�2�!o�aL��8�	{)$Ҙ-�x��C�tv��Mf�XT(9@�T�O�v�I����K+iv	
:vS����j(|}t$��h��h4%�3�r�����6�����inC��Ĵ�9�)��B�ĝ�wVx����A|�r�v:S��[��նObK���mejtW'B}�T�2����l�.t%�=M��p*:�S���WK���4��5���FbT��y���*Z�L��9����l�=��Ţt���'��or,�%�z9��__u݆[�+�� �e��]�2���&�������u��%�du�kU��/,ds%��U�:L.w}�k�4f�)N��:D��(���9b�����GY/��C�zo:	��R�o��]�U(A�h�tu�1V͆[�t��ee�,V�}t(XXӢJWh�r޳t���EG}�WYП9S�CWI���*V�r���l��0��ͷ;p��S������m�ٮ�K��$��|Gb�0�.i��V�q�vɥ��y7N�,u���)WZl9�~VVc�X�Z�|���[��T�vC�&޻4���,�ϥ�Feǖ��Sj3���7�VI&���ى��_��S#�d�W��މ�dl��X��s���NLA��H����4�D;+]w7w��<��$o1�&��=[Y�7:�n;�����Ԇte�<cV�u���U�Zg6��Ȏ�tv>)nLz��E��M�+�t*�Ɔ�p�޷Dp^SO��#3�tVg3����0]q��8���2�eԫ�KC:`�QP�\Y�k�(��2X�&mЛ�qlw��VOZ]���ib][Ӵ-�LJ�t��]�Y:"��y��͑��l`=�V�+z�)�m�[���s�n�>,�J{`&�_d3c�f����R�js	�QJX٩N��Z}�w�#�L�D��G+l�Y6wct%]�p]��8[�7/e�S����=�[@p�&��3y��v��G�7G�YFe�E�nXb�d�ᖪ]c�VY�I,nM#��謽�Y1Ι���cb�n� T�袯�R�r�Σ�J��ऱθwH�*�	�7nl4�s�u	�Bq]*����Q��+*�dTP.	��ռ��9MvswX��4�d�O��t���N�Aڵ<t�Q�';�ǈM��I't������ hh���n��h)�J������(
����h��L���)i�*���������
��C 0������
�*�p�����V�)�J���("�����)Z(��
����������hJP�������D�����iJ"����%��hB�J��
�)Jj�
J������J��J�)V�ii"�)ZT�
ZF���V�JJ�%�Z*& 
����
�(J �*���w3��]:N��B�`���7긪aZ����RohZf�A,�f�S��^��v�X�АrLQ�+���̏,�*$�Ԁ�?HĤ��4��n5¨��DO!�kp;d��ᚸ��q�|�y^���3fӞÖ�"����Uk�'X��o�a��f+��|�1{��+����/j����Z�ʋt3��'UY�E��Զ�ѷ�d���bm���9:��k�x-��]eil�c�t��-�Ʈ6�⮻7Z�er#g2�p1Gc�[	�N�J�e�,o�Kx8U��]�_]Y{��Ity�so��,.�n!�����}o!NCy�#�N8�
k�齵]�m�γ��v�p5K�{5�5)�kL��5��\FS��l�@��E�%��=�?-�|�=3+	����F����[UӮN�N�����j�kw���:OB�OV;ɺP*%�����;�S\�TIK���)i�)����p��R��SQ䢏|V
���2i�h>�+\���e��dڒe��0�ʼr�Xݓ�Y�|>�|���S���Ȫ|���乱���^a�Zy%��V�N�F��ĪG|Lߵ�gL��e��j�B��,��n�`jCX��K���ZT�_dC'\���.c�*��;(o��]O�Xs�ࢂLPK��wB��P��u����	s&�F򩭝�mFmB�r��)@,�﷤����	��×_6�M���\W��wW(ĳ��n�<Գ��6�9�9�1�F�<�Ovn�R%�ډ�Yp�S�5ֹ�����������+�;��J3Q����(yr����gts��=�,�9���5��jE�}S_rL;��c��&�)��n+��
n�'�U"�CvG@�a\�{�q-��,؎��U+9��k���B(¶z�s#�$��a�c{DL=?{]�/2�)k���X�:mT��ݬ��,/{�WW뤞�o�j�E隸�絺��6��	W�39��W�KF��sM7�3J��L�Z��YT��y��>_>��׮���fQ~��b��ͻ�i�ɨ<ڋR��q}�!جR�k�M�u����v��ue�ʎC2�*��<H^`m�X��v�{�7|���n�\������h��.�YX�m�I�3�-yh�I�9�Y�[,�4A��0�N��h��:�>�"���ڔ�vQ�3(²��[�B+���(k�-��]��.�E/�E��$�,wB�[�Gٰ$���X-�z:U��2��8��4��n����%#���k`��k+� ��A����	\��ፌ\�'i�xem\�>��η[^�+�����i��uEˠ\ʳ畴��ĩ_�[��dOh�eF�مR���Q�F��shh�
�2���eY��T�ʙ2�j�u<N�z4�s�R�*ޜr����ڇ���/���0�ޓ(���]���z�V��j>|<����\�)}��Z��\f���ʇT�PY�oLu�:��fȇQF{wc-�d?�7�p���m�J�<ո�语����Ȏ�T�⢷ `�x-\�מ���`�8��.8�P���$�a�j�)7��gR7���"�=I��L��:r�]_�5+rkw�jGi.sQ	�v�g���r�P���q�ø҇1�P6�dS徊oL��zoBg�Sd��b�E���?H7ֶ뫽mϖ{:����`�൛{���<��ď̛�e:�yS������:�������UڟQ�1<F˺7�2;i�]��w]9qM�tti��Y6S�[���h���Ǽ��ǯ3�i��ܧ�Ϻ�^�Z�^�<�OY���Su�q$%��]�7Z�C�Z�t�'�*2���\�p���a����p'�X�9΅���N�>�˼���}�BNSo���Y�i���;r��ukq��nU��/�k�k!���J����b-JY\�C��*���MNo>S�ʫ԰\��TԬ�?:�~�(�*Ϳ�oKڔ�Nv*�	B��e�?���I�Z�xK�Ԧt����M�U����܌��=��odV#r%����=S���k�Q����ܱ �%x���N�n1s����k���~�sҳ
���*��%��=���r�Uۀ���o-4��'�W-�� �T��t�Jy|B��K;&�N��Ꚏm��k����ڄ��*۱a-���l��^-���bؘ��-�R�\sֻ5�k�7�	�u"7�+�`�.�FuƓ�
J��Pw��fV.w��D�Wr�� =S6��Zϒ�Y�Ԯ���ũ\��X����"=Ff_8�e
V���X?'����o�	��@�c����PLW�Q9YK�Kt9�����J��W+����̔ը�o}m��b��nM����Ch?=�f>�e���\��!=с�$\���F(֣6'�gwr�H�?����T^�L�ў���Y����δ��
������wv4�n
I�S�s_"�4�}%m�|7�p`�O.Q$��@�h��r�����M�w�F)Bc��y�î`�s��<��V���Is�3uư�ϼ߇��;�15��a\Lk�'���Z���z��
���9��N��j�\FS훌׵��_ܝ��M������vE鱣r[K��ڮ����'��>̾�y��{W�n�J^��j"�'-�uq[��Rg�ZI˜�z�ۧ[�r����<�J�����sD��q3I�c��A�j�rz����3j���3n��dM�T	�:�b�\T�Ǝ0��<[��8�]o���:�ɭ�k:���s�U���W�K�?F6�cbl�)j��:&����qc��	�z	�|��bxNw՝��Q�ƫl�Շ9�w�w#N�n�.\R�� �ݬhFS(TT,�w\�儢�-K��/���W������j�b�K�'ս�K�[����lK���	@[W
5���t����<d�87�2��(̘��l$.l_Λە۶���%�o�A���ty/HS׷�u��뒝D*p�����i
��K.O�%��S�_.��-����E�|�@m�N�8.��VԞ�ڧ*ժQ�ݸj�B���+2��v�[fj��0�bÝ��\��B]�t]D���Jy|�7�+v����*�si���m�heG*n�XK����!&(%�}K�>��N����r����S5�r�v��o�l������7�C[�j�B�M��x���y�%��$��+'�qC�%r����Oxc�~N����C��h�z�]ۮ�΢A�z���#j\�ܿ�4���ܹ��e�w�
FB�x#�wSd7��l�"��"�Wt�锺J���=H�o�j9&��w�W0�3��;U\�<�^e�O��o��펠��g�M�͎��U4��EOh�wb��E�yIĦ*�v�E[���.�Ys=��C��\���|��w\xr�+P4��u�>X��
a5� |�Ku�����f�oK���j��{+��$�ߞ�f$�j�M�+�ȭIB����x;�2�گ�Q�f;Ԍ�k�-�m��c:�h�m����f�ơ)uw~��Op.��`�y���+�ȼ�����Л��YS�����F8����[N5�sO)��{\�ֱ�OP̙{�Ǒ�����t����.�Z� IgV�����N5��t:��]#Y�f�Y�k3o���Ե���B�wFZ��)���Z��:�}}�vr��Ӫ|�4.�k -�y�%Y�lJ��1����|�H%�����{�!��j�[y�����**��R�iBQ�������!�}�`��ߜd_Isy�1�,�Kv�N�y�*�/�iAU�+�]҅3#5L��[\m�HȾN��-=�+9\
V��A��TII�IE����"a�A꫕��:UM��ꆶ�=y�:���_oO�A�w=��Ҍ7��OgQ��yil�<��r�/�z�f�ͫlc��P���g]Ct����&��Y��];:/v��*�|fs�I��8��n��]�r���QV]�ئIz�7R�m@�k�%��F/m���܈̧�q�kw ��d�Ne���vm�(.fTi��P�q_MX��Բ�Һ���8�۷��Iu��=[h�T-=f�Dyȶ��	x`�n�q�t�WZP�Vr{�����:�@��h�S�bR�䕂�oO��R�+]��R��6�i\2�;Ƭ`��ץA
0Ff�jG.<�W���Yt=)F/^\]yT��U)
��������.����t�;�:S~j7�p+��Y�b�ʉ�Y�~3��]�3�ٮ�dvG0�S�JouM}9���k�
n���H����x�D�ۗ�u6���\�׎ܴ�ګ�/W\-p�8:��F�7Qú�X����3K�]�����׹�h���曎R����IΈ{�_+�f���۞�JW=�Y�#1����e�j�����L�����Vl�S�$����z[J�û7Q�`Uʦ�*�5�=J�v��^�x�G~h��b���8y���{����J���|f�Oo��ԯM��-�@��.�z̕c|��k]�iq���2��F��r�Vsf�����ٸ׬?B����k໵ޢke[͹Z�y�q��m���NTd�Ϸ���vl��JL�x����tLD��Y���/r>n�^ԗN����v�6�f����_J�s�/1��u�����9�Na��{�+ޑk���]�|�Wѝg[�5|g���������xh���Ή�qu0u�ڮ�ب�妟9����>31 ���z<S�������������aU��ڙ=��=�ۍp�\F8{I���V������doV]��f`�|����>�`N=�x=.+R�_�]��6�q˻V���|��=�Z�s�q�	��Te!O�1�t�>>n����̭A�����}*k�C�|6��=yP�t��ǁ�"T"����}욲T������n�R�Vb�0�&�+��~N��Qt��t�s�:����#o��=-�}JF�q�k������<a�@W
P��Ghu��1s��2Ö�_n�7n�Q�J��j��D'�k�bjq��+��DO!�4��yAȳ�t��*�Yr����/)���[Q��\G'F����ߚ�')�0n[Fj����]�А���1��dA�L ��KǶxӁ{��mf���t-ē^ �XbwB}�b�^�]�R�f�y�����Ԧ���މ]̗##U7�/I��NZ�R���͡�@^Qa��������7��w�J�$��έ��ZR�dN�E��t��b�B�k3�vc�k����[H�����I�����49 ��^U}�f���_*���+^ru{\�*��uB'tQ�ܥ���d5G��{���\k�\���mc
xG��M8<I`�����Zz��61־�Mw[Y՗g+�̨*�ov݈���jv1mYnF�j9�^?��޸���.l[���Wn�7����;_S��ۚ���.�(�^֔�s�S�9�=	w�g��Ж\6��9Np`�r�����(Ԓ�;63�A�Q{�e��j��5��ڌp�\��y=PJ�߯e�o�g7�D��wTes*�v�v}k��r�H[{p!��?p���N�#7�[Qk�'-�
a}�?LW�.������v\N
�O%(R�_�)��,}��f���2����- ������N����>�5@)%��t�Cu�/;jc�Q2XS��	�����.�%��6Roa̰Q��jvj>o/�f�I}(ݟZLT�*�н|���P��v��;��4����;�Vw��_QD_n�Ȅ�E�9m����taj��*��U�]���E��>��y*�U_��lR�`�d�U���1F�],Sw;�,��ܹ��aui�ۻ�6�;ZPb�o;2a�j�b\\����S�\�L�خ�yt��&����)I�Z��3���V���3m�[�ҩ�Z�����q8�KfE��y�u8&��IF�T�ٺ����Ee�IXe�f7���O�:$�^j�y�>���L$�@ʎMn�S��炐�Z/r�w���F�9/)G������� }1g5)�6&��|�zM �����1֎T5p�*���oq���[��pm��a���8�svY�+H+ib��7n�g'Vl�O6_5H]%�#]/ns��Fo��y�!K�i���7�(hya��C�*�N\��R7k%�	T+w���`�������u��bN�i�:��{��A3�!EP����/�r�s G5DR��Z�j�I����*�w��c�u���4�,m�����j�O�j
�e�yYfi�(�%�vR]��0�&���'��k�Zi��K����cB���rϲ�1���k��Wm(7���x�H)^:y�xmƣ�FF�
2I����D��5n�u�yR^�B���m���}��\1Өep���d��%��P�{il�)tǏ7�Zv���F}e����SMgt��fd��rEBcL���ȌY�(.�N����y����;���-����+����`�������4�_IbV��ov��|̆��,9E���f�:�͕�n[E�	T�u�2Z�w��3�o�%��K`�q[|��;�jT.̀����8"y5=v1������l���)�K�c�nH��Y�HV\ê��0�Sr�Q��V�m֬Ȏ�Ku�7�N��S�;�8�6Ĕ��z��i�1wnWbK�j@����f��X����J�ufE�R:�u��I@�
.Аlω��棋^��������@��5��dw.�'^
�sr�;�\�9m�Ym�3.��G��ua����^�sB��%AjE:���Z7���q���_�0WZ�+wm��*�^V6z-�.��M���߈�������	�)�)�&@h���t��6��)��L�o=���X�N�(��3B$�󺛗g�]G��������uW�7\
P��n�uwd7[s��[�)k��B�u;+ϻ$��vn���*冴�{	����w+-%N�8�-�M��.�gh�G �f-��Va9Q-,���Y��yQWV���9�t�Zy��O�e�A�k�ӻ9J,�n4�噖s��V����&U�
���rZB�o�������+�����8�p;��x�\�QA�v	�)@��il���l	�6��2I����W�"QE)E�@DP��RRP�д�Ҕ#@P� R�P� PD�)@�U)CAE�H�%	BR�MU�JP�5E%(���+J�	@P41P��%1+IAB�҉DM	@U�HS@R��T4+JR�@- )M*RST�R*�4 �#@-�A@
R�RP 9�7�z��y�<���Q�� 2>�X���7�v]!�{w������^�߽�N��!a���r-� �igeJ��u��]>x��NR�ùTF.�-(w� �&�S�sQ��Fb����ښt'�3��xx��ԮYp9��/��q��P�2!J=neC�
���D��B{2S�wa��^�+�s�:�R.��I���0�[P��|��Xk�xE�`�S[����yf�<vک��

���ڣ�����SMS�4�z���!�.�וW����/<��nU2�2;!;��/a�Z�)��4���Z��<�;i�W;7�v�}P3}6�'�{�u<~m�3v�>�=�nH������;���7��{ٮQ��c2���,'ʂ0�Q��\�N��x��2��Q?e�w�M�u������vs\NT�v���q'�ĳ��\���T��W��ҭ�c>v�1ųU���&�dR�r͎:wcu�X��.���*��uT���P���j�cb����V��oI�as%%���d�Y�RٛR|4r��Z��C�&2�$v�Zّ��]��&5:!�vw� ���_k�~����Ч�pk �ӧK7��;�E �<����O�1���JJ��'Y�WA����L�����b�VF�媸3���q%�Ú����76�k�J�Q�y���#ҳ�@+�/�T���<�d�2�L��z��<��Լ�޲�S�Z��7��>�i한��0�����ʢJNm�a���������qs�8t�j7��p�/��ڇ���n(,����P�1;���\$�QsY��R���\F�n�[�N_e�=k�#\fն2�uI\t���*0���	EoQm�ٮa	蠟]�]��2����Ȅ�EE�1TM�����P�pF�zn� ����f���.#�T����ahM�0��/6h��r�����>y��Ϩ)��\]5��#���T�12��R�zw�u,���ƻ��B��6`��������k&��˼tr)�)��s��]��3г��Mƻ�)���dLr0-mn���Rs0�^��Տ�u�)�\�u�p�ヴ�V�5��v�07#Vx�W&��d}��R5\�M�Of��ڹ��3����v)�̊�G.��%�=�ƴ_G���C)����|
q��dU�ôa6�����v���]]��y0�P�&D�2)�0�U��J{7�9�9S�+Mt�4/%<������w��;�A7��ʷ|���\sX���ܣ�h-�p��d��iFz�	u7���TAn(��|���ijꔄ�����L�R�H.��UDeٺ�C0*�ˢnr��;��\.Qܽ�x\IF���������X��]��u}�ge���*�ީs���^�*�g�m�+�5����o���z)���7���v���Y�v�@�=�
qn�9�Zt���ި楞����5�Qn��4��xom�U�i���U+1S�3����v�/��Gu�g�Tq���޸k/=��Щ��q@e\ՙG��GqS���F�b�I�<�-5��㞵ٮ3D�yùwwI;=΄�ݝj���'���m��+�"1>4��:��� �<�P��A9SY]���Lk�S��1�.��▊]�1�Վݙ�=&d�n�
�9�X8�i�;F����M���w&�zӄ�6+&\V���t�]x86lI���NTP�:i밢����S���!�z�L��׮S�]1�vZ���N�!���J�x��*cw[AE�>�M�(�v�zoNX�7M�L̫���M����?{|s[σ�	��sNk�B��]CA�����dN�]�.pX���.r���xÅQ��	�Gj d��H��Y8�����f��D�d�r��'�k�bjq��
�c]�8��w+��)V�[�9���W�}�e7�y�j#UZ��:5)��q7o6S�.�BT��]����+�H��3��y�Ե�}������%/i`�y�e�c;z�:�f�t����.��˹� ��$���A&����z��rmc�R�J�8&Gާw�N{�ƨ�C��Tj��3*
�D��0�m�׋i T��~o��h^��WO��ԙ��:�֚�vr���*��iӴ�;m�U��&��NT�@��끊:��+�6-�{D�ݶ�TgY֡+Gu;�[Y<ݖ���}�Ye����Ч�����KOTK簖eR����p�QYH��)��-A����ު���o�+,%���]����I����n.~#\Tˡ�	`L+.��FR��\�E��t3�#\�n轎���V�N��Va}c��ɵRQ+6�_j�IZ���+�d$9�����l�N���eJ�ǹI�=�/��Qr�p���c��J��7�/8�5�=$Y
��u-8N�YＣ[Fs�CD��tes"J]q�Eԥ�ʓtF�W�9��m&5�S�6�C{�w��eBt݋	}��T	1A.¶�6�أ�չc���Y�®SJ_u�>܄�5�7���"}��b���0^���᳠*�cYI�WF���W楁�
M��uNi��p�<wO:�o^jfD��h%>��Z��5P��%�&_�]�w�"b��YB�K��B'ZG�xÌ��ڣ��k�'7��"��\���KY����Z(�=�s.2�{��/'�G���Nv5�n�	:�ʫC���i����+b�Mq�.*n.su���*>��=W�_����Gz�<g�NH�n�j��j;�w�:��ͯa��c���3��y��!��Q���V�m��뙿}��Q�����PŃ�^����B���'좫��i���O��xȏ0��Z�{a�{�7y�Y��)�m�$JC���^��h�B�i{�Č���SkB�Wl�F��C��D^ȷc�ng!B�D��ܼlZ���.�N4�Ïpv��L��r���[����,.��w$Rǀ�+��kۖ���d᯳!񬝐�GD�"��'����^��ޖn/��~3k:D���QY�����߃\1�jY��7�D��`/�<�<2R�x��2�须�y,�
��`��x`��/;=.8�œ{��R>�ZD�ˆ��k��\탎�2�{�OYx�5��N�y��y�ÛQ��Q_�'u����s(�u�����=�"���a*��Aݛ��`�}�_��!��<;>u���=��b�Fp�u���&�1GG}�)t?q"�n�s�V�<<��s�r<^�o��Ϝ�j�^��]9�I��e�0<�Z�zX��ذ�Y_X<(7���>��O��S��߯�X�i߸�zG���={U��>���@8. �F��q[�<��+���X>���~5��;�NZ�_��x�i�q�8����L���;
�'�����g/+� ��2�o��%yN`R¸��C�z����c_�t��L �+�Ȼ��}�+n�c&�4Xib��L�>���D�]u�����j|���R"2��;��E�$���s/:n�3u�¸�|yc31��;�WV(��i�6g�[i�S�yk���S�ܻl��gR�m�vTX@.��)�7&.�En]�Hg_k<un�9_D����G�Sb�N�7�mֱ���u�&5{[w�t����L[a����ع��M����~�>�5`�.�h�TNÙ�ʿ��ٳ�D�/��n��q��08
���m{��EG{�w�R>��I_���ޤ�z� �g��P�4��¾3/�q�_N
�-�@��DY�^M=�N�;g��w!�ݩI_m�dѸ��@w����t�&M)�T��:7ڨ^�7=���ʷ�3�;��6�օdwKr�:��KH��Ĺ(;����Z(atb�[m���CŰ�'S�x"+��t+��i�p�������ʫN��2z����ʬOndg�`�w�N����S���M�Ə6�0i2[߾0ם����mփ���`
��+�s>��F�g�<�>M��X�=qyi�(8V��u�.��9�f���\VUiX� �j~Kxo�S�Up+ww(X�������Q�S���甂�9'�����/|g�ת�����v;���`��3�3�q���NoF���t�gj^����{=:t/����({)Ùͫ���{O��^_����S����%���U��;��s�<}�G8�v��WǦ����q/%���az���<2� ����ޏ2��!$�wPˈ�V8���~�0��κt���+C.�U�S��j��?�B���V���lr����ln'h�7��&屋D��#�0WS��vg��$X�d�j�J4m���v�{v󃩬�ڭ������N�ȥ{��~������Fժ�W޿������q�����m���fUcqV��If��%і�)*��9���>��?^��{�̫��t*fs�^��E�9�u1:o����'ƙ9T� 7<H�Z�j7�k�ƩSrFz=�d�Ƚ\�%~��s��؇�C�������ݱWd�@ ԏ:[���.��C8�T��w�kf�	����#�k��q���q^89�~��̦etI,T*���Fz��}� 
�QS>��+7I��,	�f�t=���}�E����l�'�����X2��\�ɧr������2h�o�_�߆�
�rѡq^���GYϷ\�4=JZ��%�ǭ��H�-o�i3ݐ�r���5��#�Γ��Ʌ�%a����dm���ަ:��2�܋{��{�
8S�]�g%T�Ѽ�^@Z�_?܆����>w�fP�:)���)\�>[�Å�u��7*f�9�ܱ{��ּ��;·�_��t�'�b��ɏU�&�x׷��G!5/Jc��(o����PL�-%n�/��K��=}�s��ڹ�n�4�b����D%'Y���b�&��y{�E5]�[�g�6Ԣ���{��:nw�Y����oEOW%z�"�wLJ�&�ɹ�y�K���ZS6�� �o�[�&꒣7 �m�� �6}����uU�&�}/��,>R#Pyu��TY�͠&^>���U�m������T�9�8�Ϡ���������e���9���ȅYư�&t\/IӾ��`f!���ic!��'�ti�C�rπW�߁��x���^��j�w���a�mV�]q�2D���ٹi�,��o�G��.*g��[�ˎ2[�x����?�汘�92����ey��^a��!�ژf}�����=���n�����x��<����T߽UT�_�ލ�jәn�����P�~�=�>�����Y�g�*@08z>�Rc��}���r�3[�6w'\?AK�����r<�}@{��UHۇ�`8K� SRX��-a����6�siH��C���Uc�qߕ�_�Z�4\[;��Ǭ�1��Ԯ3��񰠎*��q3�C�o�e�9������ �X�����T�c�[f2���qvJ��@�����ZZc��ޚ�chOv�U�%�#{�=Dښ�x��)�w��dm�j��O���%�TU�8�Gy��]��v(�����e�:�3�vӎ�TVvm6i8[Ô��t�l记5t\&�-�0���Z�n8��b�w�����*�gs+cP�U-������,Pe�yǪ�ު\�.�e̟9m��ӹ&��k�%8��㠙n������0)��Mˏ?VP������v]����/��v(��V����w#��UT&6�R&]zNo��,��=x^� ���K'���}���NE�y��㮮��O���62���ԭS�<���~�P�~���̎�L����p.6vp+�V��_*eg��Q�y7�ۊܣ�X}�}�����Zhv9���u>�ݖ/�}�9����A��W����[�a�=U�}�L��w�C=�uxmº\N��_V-A�0����=cH��՜z<m����T���oN�ۤ�CE�zg��N��9GE�iW��]L
��,�2�~�:�747u,WF�G�~�����q�K��
�e����f=�|��ZlӠ<���k�����=Qh��0kd桏��k؊U,n�7���ʞ7gĥfaᯌ�C�L��n�n:dx:���Xnq�-no���Ԧ�ft��}������exyz�N�ж��u��'�G�W�A�P��3�ob��г;���[�^��aa�Hm�r��>g����b���e}/m� �.��O�_|:�?���<�n���(#_SB� ���.8o��V�Dfg��rEIDuQT�}��6[�*���aO��K];�5rك]<]Dm�QI��*]v<՟3m���0p�6�]-d�W�V<�?.����ylE�HkZ��]�k��<f�U�c|��횎7o"�p�Gn�j�R��S$�j*nY�ۼpݺ���Ε�ү��/�S���n�(;���87u���ɂ�_�
��<��Q�*kaW�*k"�
Ad����8��v�fS����wz��԰�&#����m�*�����W�D�Z�����
���v���G[�U���
���E���օ7��j��*I�lQ��z�(�me�.���VƛB����7�{�O���k+`EΣ��Ǜze�1b���:R�o��r�\&9r��znIu�v��-�j���.X�T��N֎œ�KP��j�ʳldx��ث^]�1�k�wّ.�Ӭ��A�s��T:^�k����B�╴C�m�˺Vu�|�X�vC�,�KO"��z�T���gn�K���P�0��₭�����U�\�c�v�����{�)|�>�V�yY�)�2u,��,6ȭ�%];E\��5#u>o��=Im���aPR�'GO�,��g<Y�:���8�]{y}>d��0Ɛ�N	]���0+vS��r��έŦ�/P7.�=YB�=X��*�-(\Lo7��0{d����f:4�m� ����MƉм�U(F��T*�0Pkj��=�}[�5�^U�f�']1�1	ַ*�	����7�2���0����MɊ�ǽ5qU�0���$օ�\�t�'7X�r!�&��/o-��3���}x��T��P�jg]�EVm�k���S��n�����"�&a�2�v]{v]JmTðJ�������i���`���0ǀ˩�TK��ƾ�7�!fF��tލ.����Yb�I�HB�#��f���sע�&;���{e�*4v��za���C�Q4_P��C�c���cB�ie[5�����L,/������0��e��Ey�
�zޜ�A�,�Rz6�͠S2���s��~`'l=יY��v\`�_l�#��K�mB�3QV�Y`90��SVY�/;%aQ3Ӵ:/���D����A���MF��	6���3��Kl�w�qw.��Y]\�c"u�<��Q�A_��#]HAy�����E�2���ʙV���.a;��2��o7-��(ꊥ�A��}�;�w�[�(*]'P�q�Qcm����XW�a�k��>Nݾj)Ձ���W�4
X��b�OD��U�
���Į�a>��W�v��2����M��m]����s�؍�U��7Z��wWh�E��vi��+J����Z�I�|�aN�TEY�N���<��*NI�,���Û>}��T3y3pv����n}ـ�[��Aٓ���;�|j[��5�����%��������B�F�j�)Q�
T)R��B�(@�J@��
(JR��((J�B�hR��(F��iB��h�J����i
�����J�(@�)E(�Z(J
��J(�i�JB&a�(�
��)B	J�)
(J ����v����2�yS[y�(*$�B�S��k���g)nɗ��(�i.&;ih�H8+]5���յ�ݍ���p�R��+�W�/�L�J캖P�+о�����g�зg���.m�CƼx��7��su�\�f�0kKc�.�C���m]?���	NZ�_�x�i�q�8��ֹ�>�QQL�Ѡ���ȑ��,�=���2O�GA�A���I /)����q�ևr�w�������ں!��EL��U���X��(j\����z|=�?z0�1+��o�/��	��ϖ�7���,M��7��)��z]j�h�ޗ^%�N����:>���jϦT#�/��n�����p�o0m�Y��i�k>�y���W�7�z�>�O��`�4��¾3/��NČߜ�{����n��Q�/K��nM��83^ �7�I]q��(6��y!����5���Z;�h_Rz�~�t�N���E���²7���\<�ii�c䯝��C��z���(�h�������dz\��n=F,�l���P;n mh��O��V���c�;n�xbu呐����߮7����ʎ1̈́��[��{�F��n�F�5Dv}5/
}����L��\_�5���{����Gv�?�h������?�I����qT�"'��X�&^ecõ�|�e*�rGh�Ż����;>�S��4K��ë�S�����Op���1��eAg�F�[XG8�.���;�n�Ɨ�k^���G�7�ǽ7y�݁�c�_+����ʻ�s����B��ʏR��n�G#@�9ML�_1̝��su�����
{����/ޒ��Q�S�?:Ay� �T䞻���L� ����T]	��#4.૞#�s��a���.Y+z5���;B^����{T���ֻ$�q�y��Ar�o\��~��&X�����R�.^�h&;��n3�<}�����+��֢݅78�:��L���7���g�i ��AH�u*����F�Z�/z�8dyS����� V�{�n����>95]�9��� ��#h}����J�,	�R$�ҩ��M�	������aD�@�r����j���o�ǽ�==�'M�����$��"*�0�L뉲W����j;>��N�^�+q�7�'v؇�N��W�/NXnw�J���:�wlUÙ.P 5:}$L�\=�K��ɛ��s�=hW�^�j7Ѩ�;��5�-�/&�Pڿy2��:d�*!T�Q�MQw�Vl)C{�s]ZϜ]�����~��Ce�2-ojrW��D�����X9�H}��wc��V��w��oG����p�G	:���}�.�\x�p�F�.7���{Ǥ�!YVz�\3r���FnL6c��ry[��1�-��9�7'��K���A��gZ�tY*���']]񒃱�����O�*�R� �Ij���S�|�r�w�!��;�U����;���_�y~31�cՂ���и�J�W����~Ԡ�5�FJ�{�W�
8j w5�T������!�''��DTvڱ�n�ƻ��\��0���U:�.檻j�33^���O�Jz��4X�\�;�O�T2a��	�0��[��\�>\��EW;=;�W��NǯG>�*�����ޑ�W��g�?uX��R3K' X~+�P�'�ѥn�s���=��/�e�g��-��V-O��2���_E��Dj.��uDF=_�Í/C��,��V;�Ź���F=�1=3�|f3I�@�p􍷨:�����+��Y���7�2gB蛾~��ʺ�o:�5���φP�C��Q�'�<�a`r����+����u��j�}�A�9;�2X�:�b�j�vC쩎(x�� �c����7��2�t�����"�ǫ�}ǵ�~�y�q`el�n�Jo�9�^��F:ʖhq'���*���H��w^�-���o�)�A��wm��-Οp�6'�;����SҾ����%�4���p&�C�[+h����uuUө+����v��6eȤ��gp�;).\�	�5�<}ٴ	Oe�O{�lU��ⴅɈ�\Ƕ�S�F��f_�T��{KX����ܻΛ�G���N�3��u��w�x�ԱB��Қ�s�G:�M��n\�nv��t t����G����^̈�ݐ����/sB8�q`K�B-;5�<�2��>���������%Ӑ)!�Qѻ^Uޖb���QP���>/�gUt�==/dN���Eų�ls�Y���R���ę��~�L�+ފ��������āހ�\��P�
Z7�!��m�Φ���%7@ד�c���hd�u�C�g�8��A>��DL��кs�;�O�����m_�=E�Y �1\�������n��VM�t����"F�pq}聬DTvO��k&�S��G��Vxz�`?��jz�z�����>����Q`k�܃_|������@R&;&��u����G��NE{��>�
�&}�5�Ǽ樧��=O��4��o�� �)�*�������]��(d#�ߵ��ׯz���67a������7�_z@��������g/���4������{�݆j�y�>�%�9(f��q<s�_��Z��K�����Ew���]�������ӱ��m�Α�ݎS�M��t���L�t6t99'@�>'.�nydxc�^���eN�}�����k��A�#��z�[5�OUD��f�J pGƘ�tƲ�Z��Z	syƯ~��vk�l> ��	�z�U���M܈�pf�Y�52��|�ap�:Yf�����+3v���Bn���H��O6��Pϥc���e@��mcÙ���jY.��� ���O�ً�ʝ(2s6�ʁ>E���kM�t�l�:�@���eŪS��dJ�J䥾@��/��C�����*x��)q�xj�C��R7���HϹ�]�GDץB:-�|��>a���vE��Ol{+��#�hxvC��.!��qsĞ5W��cds����V]\��-o���V�MI�����$:��˳l�����=�}�^W��]9�I��ϺP��~���y�i�����G��)c�]O��ubn9����=g���Aޡ�EͲ�ڲ�l���F��q�E�K}`��u|�r��[r�Z�~9�Rq����>^�[G{�4�����W���q�^��vc���Ww��2K4��ʾ2���,��9�K
�_��;`Ё�ͬu��]Uy��Ju���w	U�e4����:|=�k��������܋�o�joG�.�llSp�q�zB�ׯ�>���>��%�Ӏw��P�}2�����2��GׄG:Lex-�5�g<�ߕ�^�q�y�1�ڿQ���HdW��s`k��/��(,����N�����'���ڴv�ʅ�F�U�\�8dOB��TL[�ՙ�T_���i�;��su{Œ6�(D�ՠ�=�`�W]�&��	����nb]�P8��nf�|2�)�l�}(R��1D�]�]M��(�gk	=7rv��Ç-��I���((����-͝~@�^�^���v�r��)+�5�%6���^�Z��d����S�[Y�I�`҃_��G���V?k�.Ufߴ���:��y��P�K��wz2��6!���ˡ��'V9��;F(���:(�����0��V���c��۽	זE��wORc�%'Cn��\���=�4'}��b�eN��ay|'tÜ�q���`�?9�C��勉�dgo�u����u��!�z��r��h�;�uS�,��0:��^��53f&՝Y��7$�mGfh�}D�'���Yz_�%Ǯ�|�� ����B�NI�>%ٗ���Uy�>��ͧ��ᶇo��)�x۹p9������w���t�ghK�3+^Wy|/b��FW2��X��Y6MO��[Jsĕ艟�2�\T�S�[�._zh8�O��g�x�Ms�gj_ �<�G�f�J���R�c�ޝ>���>5ă����b�U!�S�s�<ub�!��Æ}�=Lk�mm{��MZI\"�3s�Vw��^��`��!�O��U`H)*��9j����"����%ў5�<��b
l)�q�7v��[Y�����@ӥ�B���Y�]��+3,\�Q���ؓ���������2��.gS����a��jD���$�,�ꇹ��v\ÁmEko;R�yC�hTD��#;�&��X�aJ�w��Ns͛X���KN�p����ߌ��z�w�g��@�Af@����08z =ӄ�N��q�D��®�@�މ�¢��3�m;���yb�k��ǽHq7�Q�b��sP��$%�����P+��v��.�����V�Li��o����k��q��e�ߊڿy|�S2�D�û=��_��/�{w~�mMxӑ��Dk����5�ds*�L�[ڜ����P};�}�XҾDVx��NF��3�
��s�����;P��za�3>�v�ؽ�·\�>{3f�hɽ���:TGY�^��s����r,NF��Y9_�}�c"Z�Ѵ��iGu1��;�Z��y3ZpLL�*�"�ۼ�+�����C�7�O���<�b��RGO�U&\	�0�+պU�����"�\8Uڸ(E�c�ז�s>ҟz��^z�zz_�h+��xY8����C���wQf�ȼ�,���VX3ɳz_�-j~�������{)�<��r*
���f��a�}�%LV��ɟA�ѷYU�Il�>��۶�Pc�zKg4s�7i�+�~�~������)-�dݐr��.\uj 3�
�oZv+{��]w���Εv�8��.����z�6�Z ��O\�O���{I��m�E�P�r:��RΣ�q��#�z���RR(�Y[�N�Y��	Ϯ��ֹa��; -��;�;JZ��N��;�x�^�ߑӷ3�*�_�.���N����`-�F��/��6nP�&Խ�6x�3��_v���]��}��*xݖJVe��g�O��rNM<��"_��Q�7;^گ8�7�Y|�"b��Ny��z��c��a��f���f�T��S)��̸�+������R���@��z3��|�����_�l{�y(8�Y3ĕFa��>U�>��R]��1R�r���_]TK>��B<��gϢ����
�cր���p�N@����7�xx��cэ-�p�v�E�*��ȯuG�#��H������=��H���V�G7�n��۸��VF{�{��3ꈙ���~(f|�n>֩�u�l�A���t�t����	ȟ��g�q���Xg�"���كh��<̂���ŅP���IS_�C��Z��7=uE��p�ix�4�%B���Ө�F\��0�b{T��Q�-lծ�=;��x=9<j#���bNCI]ж�x�G���C����r|����݆���vM�;&��V��vP�\�[?4�zȿm;��c�\5K��{�I%>�s{w�$w(��s�n ��t�Y��b�I>�e�����6�D���$/iقCo��V��꺵��,��oO\�탑�V�Qq*emKoa_d�}�5�R�P��H�oW'�1�|2�$�=6]z\{��^���y�ѷ��=V�~���w���>%T��ܬ�e4I]v�XxS�Q�f���9�9�vn6��R;��7�{p�]��>��>ڟ
��d�*� "u�}���=�j|���Ƣ�ś�ɩ�Z�j��p�ds+�Ũ:�.���[;nd�s��*(�j5*��e�>���R?��grsbe�T��*r��*���_F�G�C�^�� ��Ϙ�f�a��5,���^�V;���d��������^��_��;��N���L
�%���Q>5����#�=���;����Hw{%���E���92G)s:i6�-�@{�
��k�J2��'�����Q�yλ�{�]���:�B�ʑ�sĞ5W�f���]b6��.���uh*qޣ/�����}�#�{�4��=v�s����eGZ�u'�6���p�'/�4	/�6�:��S�Yu,�7V&��xk�q�{n=�쎴ps��4�褼���l�@8= ze�?(�7(e���^�!7�Z1{�m��,T߼�.�U��_Q��`c��`���5��	.Ӵ��=ckzw�t]��ĩ���9����S|:�c�WH�M�.����܅u��(){��2�Z�"��!��`�e�W]Xo��2m�>{+�7@�tKN��'�mIj9��N�.+/cM��v�hjI����@���}$Y+�ra/�_��^]�o<�ͺ�%���i+��q�����2�M�0xΟv����k��t_m´���].�W_Y�˖�K�~�k$pOΘ�sĿ@���7���.=~�W�%�=�4�rc!W���d:�Kd�R_�u��7|s�������|[������ �X9
m��W~'aܼ�g[Ҧ-N��sŚ���~�&�zz�}���L�ߺ�Y2Sn}�t�g�5}�ʬ ����p�ߵ9V3q҈/��M|rP�
p;�Zt\m��
ȍ�|o�����v�c�Ez�f�{���������
1y��d	�u�}�a�7Œ�d�V6�;���t\+u��Gu1�ڬ)�M�?N���}>^�K�ѭH�+�Ubz��z,_��(�g��_��#�j^�ߍ�4��uݟG���[��F� ���3�^��/K�갑��AF�T��>'v��:2�ל/�1�@/:��1u�N9�V_Ƨ|J�(�|����~����o��?:Ag���$����6�!zz��r�mmt?5����7OfS���5Kj�هgh��Bt:�ɹ�,��s��	�M�a�vY��V%PӺoE��h@�!�	\�u��Y����)�|�n�r�m�KZ�$B�F"�Jw;��w�K���dP8.^���.��/Zi��z���;��n���ƩT�{,��nfX]��n>7v�ۈ��Ţ4�Z�D�������0��0�m:]��wm��ī3H=rﯘ9*-�[	j���	��Up�.�aD�4�j�t�NZ��חi�׭�����|�h֭�1t���O��mr���m�L�Ux��8j��M}B���.���oK2����f]�J��J�Y{��R�����0�Ȯ��ݷq��8����Jۋ�N&��N?�D��qK��o.��qi�Ќ�M�Խ��R1Oz��5y��5=��j��Zn����k��\'AwwSS�3V
HȾ�v��mg/u*�}b��x��|R7��H��I��c��<̝wiq�Y>���<��m���v���vy>�>0m�ۺ�t�J���0:��f5t�iQ�M���ܫ���k�@���&�	:����i���-sx�nZ2��͠�Vʐ���ܓ����JҞ�r��3@=ݝJ�nʔ��wwlRֺ.Ʒ�.�y�*�ek����u����qb��q����'�$k���'��ת%��#Xz���跇0_>6vȽ靬`�ǥd�&gR��ggun��(���� ���,Fi�[v�E�f�݆&	`�k��w=fE���è���PL�	���m-Ӝ��z�
��#���0�n�h%�֖}���ADv�W���a�ʆ�K.��R�B";y,X�t|�54e�Lo�cwu��j1�ٱj�VƯj��ƚ����r2��w�����q��n���F���f�c;�qiʕ�ޓ[�ي�<�"3-gWl���{8�M�x�r�O�sOI굅�7ZM�w� W��qcz��hM�f��V#K;�N������x4�Bo�E��(���;�	�C&
��
�%e�Yb�|�n�F��NL��+|,CiU�99l�;2���
Y[m=�q�E��uI���rL;����0��:�=�ff�{y@}˞a�u�/���4��őv,��;�U�AT��<w��E���v��w�Z$m+<�����n]gWvwr2�I-{�F�J�N��f��.8',e��vˌ��o���(Jɷ5��J�,�"�$$�F ̮_Y��r��h�B��>ڳ���@8#C��@-n�e��>��ʺC6�O8 r�<ê�����H#�,��^�,�9]8nC��:Vw�#W|�'B0a��b�F�s+E��;u:j�`�u�.�3ҁR"qrz�+��l��B4�D�y��:��H�גu�bb�{�6��9\֦t���87F��Bx�V�©Jܚi��D��Z�����?v{﹞~��}��!BRIH��	H�P ��*P�� (E
R�J%U�4#AM�d���!J4�)BdD�DR�
P�d9JR�*d�NB&BR4	�*Q�P�% ҹ	�ID�Qd�J�K�I���$&[��W �ht$c�{�uj���J���S��9s���d�R��j����"	����%8P"�dY�+pJՋ?AS��U���ǟ!�r�咷�YxԆ�t�C2���-�l��ش�w���Ϸ�%�^I%TL����>Sn���}��>Dg�x�N?K�V3�[-Ǩ�9�^岥)�,��kQ�Ea�k��`t�X��T���z���V*�}���R��B�SPn��SG���mϙ�ϐyG����,q%��R$TKjr��X�wr_�c.��yOÜ���u{ס��3ϽCN;��QϹ���Tdq��l�= �N�BΘ�r3-�PvWr�mik�#Q̡|�p�o����,7;�%ۈ��JئIs����=���z�XH^�l�����`�^g��4u�1�߭�N"�l���A���_9�ff}}C�%lx��^�p�X9$��T�SI�[��k�c�����ojrW���Y��|O���&�س�C�v�f��*���Mi>��#!C�5鎌f}��{=��/Q�~Wra1�~|�|�uo��^b�fn��,���t=�,NCF	���������K[z3�^�Y�Lv���g��]�|
��0����Sz��~��q�E�j�hV^Z�f�ȑp�[��=W�+��R�F c�k|fxNbw�B`��]�t��Yȩ]����W4&�V�׶���*U�G�-7J�ԯq�Z"��\�U�=h�ee�I�&Gct����hM��HrO�<?|�ۑo}A����	�;�Cc�� �t��C&X��
};�wz�e�� �
��5����U���[/�������z��\g�ǧ���Z̩{,��p?4����tv��<�՘�?��>��M��YkS�|��Nyׂ�:��_{�8[��9����>�d�g�w��_����=��#�}�&�l�u��Q��o�=��Y.M����%����R�d����(����3�3�}�:v�e����'�ti�C�s��W]��N����V���Ω��}�9N��	�ew,��La�2wp�P�bI�;n�.8��⒫6��H��_SP�9�#���1��?>��z:&��SR8I�3&6{�	��My����1m��ѻ�����?�_�e�X;��ё���;���~���9/iK,i%#0�;J��d|:g�� �8�t��*{�_t�vu�>��-ϼ��ǭsI�׍�R2� ���ޑN�D�G�� �}' ��W`�q��4r'�Jr�鯋�gp����q ����YN�31^O�t��r���iF��Sڴ�W����q��ceD��ӗ���,���y���zh	޵����DAM�+���Yk/�_�^#5Y�:�$�)�@�j���N]��Ԭ���)sp��ܨ��m�vGI���I���랒Wr����7*�uX�r�ڂ-��9�^���Dqu2��p0��KF��C���#�w���3�p��sL?W�ְjn�㞿g���ꪦhk�,ҩ!�DL��4.����@S��*#8Z���u�rsҫW�h�z_���N���=Q�)Ө��#]�2����'��~ckh]y@�q>�I�:}����r���wB�u�}><���)��A�,��C�}�	��_O��u����\B��G�rm��.��+��?S}*Jn}�(sO�����\G{.A�S�TO�o{��U�[��黴���3�986���۟q�:��7�{p���8����j|+z�,j��%nt���g^y���=�_�Z����6��R�hj��p�ّ̬��:�/�n+�ZQ��ӕ�,GX��S�7�]��?+�P��l���;;L�~�:���J���]L�+��%O�A݀�s3���.� }�|V?U��*�c.�p�E��;�>E����pi�^�0�����;�Y{�a�^`z1��E�����v=t�^Ez��9�R�g�Y�)_�f3����H*
��"�ZS�)$!Mz�.�"hZ���_y��N
�Y�.�x��zea��v^{.vb\E�b��y%����$��v�f���1��f��-�rZ��-E,g-
�k��^94�鳭S��U>}��^-GX���ۖރ]���ה�9u�&h�/����|��x:�0�4��E��W�=�{+��=v��gβ�j�GQ�N��q�Cj��S��i`�HhI�±F�G}��c�f���{���3�>�%��W��9���>�����N��I��*�u2��b˩f⛫q�߸���z^�C=�9��<��$�#����Y��g�d1��.��@�|v9T`L(nP�WO�+ޤ&��z�Ѵ��=\-���z�t����}������Ps��v�8�YP Ծ2� �H��W��,,�����]�נf�"{�ť�=���#ӽlv�?N�(Sh.eȞ�<ti��l�0��r�����N�}���yak��'z�H�pߝ��z}H�g�ӣĿzp�_�&���e@!����28��Pxk�f��mw��]˒���ns$6o�����S��nw��=^ w�́���U��v�����Y�k��G;�T�39�˜�:+j}�ugk��)+�5�%����fT�XIӬ�A�پ�y�n2���Oơ�/����+N���Kz��yp��W�������SN���Sh�6�;��S���ܨ��*n��϶w�v���|��ݫ30�ך��Rv.��@��ʗMa�4.���o1���);e�*���e���Gs���R����剚��z��t'��3Б��,,ّMݧ��
r�g�M÷8#�I�5�엻=�jNy���Y;#��l�}>ӡS�'{�����Z�u@]�{���̥�=ޯ,�ޑޕ���u��D#~�j��X7du�5/:�������\�
��oRU����U�^�~�z|�^^��ua#�ym!q��#.!O�ݳ0��Y�����g99�z�v�x��9S:}��J��LKZ�.W���v=u�9�:Ady��z�$�oO�ȳ�d�.���,�����?�6F/�ft��8y�r�+.Y;�Yw�:A����C3}�i�0jT�,pX����iw�;"����$�L���qS>S��K������ޯ�9�.Ϯj026�����9fe�wp�o�9�;���#�2��5ă�e�1�>E��T���u�s�X����<Y��C�ۺ6�Z��·Cc���;�*������G�$�L�%��R$ԉ�]�꩗p�j7B���\��=
��Н�㝎}g��(��A��AfGfјp,��a1mʟC�ij�������;T8�z{ȝ^���E�Ӗ�︛�o�G\z�ث�̗:��K9c�w�9�|ʻ�����e��i��g�-���=�Sz�}1�R˶�d3kx�d�t't��)�L�;%������q����ſ<���V,�2ml�7.Z���>��{/X�ĸn��\G���dȻ�G@�U��q���Ti��ٴ���4��^��|}��4oZ57�l�w��G�p{Հg۠zM�.+R����G5KH�Oy��/a|r�����5��e�2-ojrSp��n�A��v	�������f���
�H}k��]��s�ה�X��iw��
�O��G�f���!:Eս1Z�a�h�C�1�u�b@�h�2�'${&X�a����m9��+׾�S��on��Ϯ�1���E���M�O���<�b��R}��U�}bwL.P㽬�Y����1����W;������yח��{�|��<j��c�ӏ�V-fT���N���P�)��ˬ)mUVwz��g�F�&�t��hؽ�g.v_��e�4�_��|�by}���ܜ�<NϏ��C=�^�s��fЈ�2v/ܦ�l�N�t�Q��o�=��Y6�c:�	��u<Y�dyU�S��\έ�Wyz���9�:/���ۉ�2��u>��K��=��`+�K���.�b���ۨ�����.bEy��^��9�.�B���("��@�z��x�u3�o��e���Mȱb&$�g�E��2��<]��O�ᗁ���&㛙w�ʕ��#����6mվ+
��=�dY�,C N�er'{�kqb��#� I���{؇Y�9�Ƿ��yf���֋�p��:��(��P�Z�e4C����W�*b�:��k�B-�w�F���b��~*o����mLqA$�̃=�7gC2l��kIt��OR�����~�lC�v��w����@G\�"x����{}���:��S�y��8�=qF|�ϖ]����M�Ĺu�=��9��7���{1�\�~p=��a̛2]W�{����9�>`{��nl��V8�����H��ZW��4�~؍B�c}ב����g������ ��(�@n�����n#Z�9ϩ�4|w4�e;���KW��׹�AS�M�~�;~����©!��u2W�и�=�O���v�����3#�;�+W(Z��ڟ��8z�4�d�yȡ�="7Ǡ��&azY����%j�c޻�Z��������{�^�����*��n�O���g�wC�܃_)d�!�{9%�����<\��R�O�G�o+�r�Gj�nK�~�:�7��P����}����J<pgv�%�7a�[�O	���#gg�;�~ۗ�Ȥ^��{p�]�������xW*�:=~;]�=�d��ڔefN-l`J���}�2^}�	I���nT��ۜx$�A��˜[�%by����f�٤}��ٕ��i��:ZV�v�;�U�3��5T�\pҼW�+m������!@&.�VĮ�i��[V�H��G$Czg�O��v�O t<�~�C^>�=�j�q'�s��?��y3��
4rXW���6�]>'�}�/���Ǳ�׸���x����}N.�q3��c5 qߕ�A��(�,�Y>�᳡��:6*�N�.��F�"O3�ՕG38,��^c���O�ڛ����Vi]Tŕ���FT���Q�1���H��jN�d����|~�|��\�?g��]?>�7OG�ԅ�ڞ("��@��>�}ӏ�	��bn�ދ[���x۷@72<�O�dk+ޝ����<;!�Z�T��=�(zH5�GI�J����t��FL9���_b�=o�dp�����ж�=�������pd��G��;�>ތEߵ�%��{fX�rKs��.���n�M��߸�w�x�*xl{�U]K��d�[F�A�8���g���� ��Te��n�r�}j���W�HK�"��u~7Ri��1����7�����mi����%��A�D�� �7�6t��>��;��T��{�6����@�����9��M�l��hOx�7��v��ф� �g�gsf�F�9�5�ٱ���Z��mY�fmv:|)a���`�h�N
�
��V>�n�ݫU�[h�-���_�8d�͡��% 0��}O�1@f�KtZ�>���!6�gX̷K�m)�	f�VI�<@�TsW�a��o��S��Ĳ�!��RO0�o;�"�����^��k$poΘ�sĿ@���/ޜ�~��O�T���9Z�\���_Vwz}b���"5��BOz�E��w��S��s�/���|`���[wu�;��{)B]>�}���΋3)���uh����u������L����Mt���#"L{$��x��u��Pێ��&�Ǌ����G��IXpv���ާ����~��ϯ
ɜCs�۷Ч_"��\���b���P��������\ߺ�^��t�=#������#�ds�H���w]�c!���ȇޠ�/|�����Pws6z4��`�EY[���%C��켼���������i���;�� *"���3�U��qz��/~�	�-�.72�e�����Gncǲ�Ƒ���v�W�L��~��53e����̿{�6�Q���H��M������.Ѽ�L�7P�Z��_���m�É`#^�v���(xmR.���iJgq�Cev�a&7�c�(�zs	/Ew��g��rxt_I'�eBg���򘾷B\�頮�`���sF�wO�|y��Y:�1��#І��M�P;��=��հ9�H.�d9��t����YV����]�~��=�v��[R����:���f�����mw|#��[��\�ܫhb}Xҋ7����c�{4��X�����p�+���nI�sĄId��B&��{ҼVEy�{�!�j7�+�w�A���&�,\T�B�����ֱ7���"n�^�J���o�~3懩�����G�G���ǰd�j�J�,	��k2�x.��{o��i�~L-�v����>�~�.?^��{�̭�P���'M��~��|2O�2 r�kzg�4J�(�y�mp��r咾'��V��v=BS����P����ﰕ�1�_���"�����a��&��~�/�x�9�|Hu��|}}�CF��Q�߯��kg��{C���+0�E�
��Ž?�w�ު�k�%�$��H/�½R��܁��n#Z5p��Q�yz��� �/��lrm�Y��D��� fY#!\��3�V
�=�B�Ҵ����6|��P�=Yd*��ɠ�x��ܘ^~�'~n�:�H�#!���O�=P;�: ��ב���ױ�XM��j�r��5�S|��1���E��So��'��'��#�n8(����f�y��"�qy�ʽ�c=]^�j��Zߣ��pΫ�n��q��x��������*Fo�W���s�u���1� ~�4T�yn��,-������W8ᬩ4^T�J<+��h�oAB������e����/6��:�ͧL�>��X�ĒG�٬7�.�Vս�7F%��]{D���+w����VA���W[��ti��G��uA����!a��gA�;f�>�_x�Å�PXER�u&k�]���ap$�+��v8��J��ݢ�u��&b�`���R;��DIU���w&\�[x� �Z홮ݪ}	���N*�%���b�82���$���p?�9W��%%���Ғ�������+�(�찬�(6���r�kQ��J��6��+�����|�ׁ�+r<�HTӦ�M�`��m������i�z���iK��<�P6 �3O�ĺ�؁u0F/���~v�:�H�(B`�94f�����{�aJ�:ء�0��8��p�K�u�ժX*_5�2��j���f�=Zor��n�!DY2)���V�s���u&�=f��K`��SX5J��;��|�j�gv
wj����@=�� �ǈ���3���T�5o5Zn����a�P8���Pě���y㙙)X\.�`�r��*�d�i��}������괕IQ�4��S&����/��T��p,��Z��|��ݗ�¹�n�gJ�#�lA�A�X㒉��)7S�IG��)�ׇ�H�	����vQ@vk�WCqr�y�狚\�R��A�-��@��ipr\�O&K�͛C�]��Ǉ���A�B����î�D�����%�Ҩ
�B�K�q�|,@rA�x�r��j��* 7m	͛F��y^i}���++&};�v�1,���_��[cD����WYR�+ɤ�
��i]�{����+;"��Y�Q=AV��_:��*�%�ǂȋ�L�9�WEN�
�78�:b���7�<�E�!�I�W!��䝟�����q)4Kv�)��J���K�&��t�o�ۄFc�+`���2�b�{�� �vN�zJ�aխ�};����j((�x���Eu��w-�؛Y�-��9�s�.PO�K�6�;hh�����%�w��j�Cx�ʛ�&�aYN��ؐ��-�͡��kw�e���idL
e�wq�;B�ة��Op������W�1�M;��v�
v#�S��K��2�ӂ��o�	N�g.��"��'E�;��#vD�z�ܓ���{J�,B��{��J_+�#6�����p1�u��a��ٵ�Y��ڷQL� ��Z��>����Yc�Vm(Vs�i�:��X���Qj�V	
0w]sJ��5I[z�Gf�-�R�NˬY:el�Q(��^ q�y>Ւ�.=X�lWYFj �s^�:EWE�B�\Qu
���9��^"��t��M1��ZE���p�gp�,fe<BS�Y����k�yd�r!$�\�;2�\#.�ڱ	�r��]FI�k�뫎�_�{^��~��}�Z�D���$S2��$(����
@��2p��2��L��C!2F�2�J
U�i2h��J2)��Z
�rV$V��L���lŠ%r%�h����
���X�����
@��JJ�R�(i��
U�%��η���o]��!��K_�_*U3C��`�݇�J\��m�Q�W:*8���]�@�=;���fJ��3c�V�;�^�w�wV!��X�ڏ\VSF�Խ'N}�_��ڿuU�'<��y�ǝ�JB�C����s���IKC���9q��Ӷ^���r�jg
cY:}g��m����Y7˴���9��~&<r�SIn��J��\.��<���`w�p�>PKG;_��t<��*�Y���b]�ܯ��Iyf1�nm��A��9Sچe6��_^�����R�Ȁg�3�G��ޑ2V]�������r��c����k����_��9�v���<��`�)$��f����S�m��U�*�EL���K����{ף#}�w7���=�c�r^� d�n���u­J�����ȓ��@�Ū��2�J�|z��r��yzG��F���������~������J{��� �.��9�����
#��V9O��o��H�����)W�2r{�d��J;~q�T��+��s �J�>����`?/�
Z:ԡ�j WEǦ�x{�D�٩�r��k�͂��nA�3,ϸtA�#f�W�O��ܬ/�c�3�6zmԒ�_e�M��!S��&��I�i7$J)F�M�u_��k���qVJy���5�ձ\����`�#��o���/�wu�at߰��rwM�1_�h5�����Kdd9w�E㸧8)W��M=�yݫ%쨶�Ѝ��1��;c�Γ����#�ײ���Qf�.-���"�y��|W����PSoz��\�?�Xy�ò�Y=��+�5p���w#���wA7>'�z|�>� ���z}Gݳ���rW��B����d]�zZ�ӑG��\n�>6���3�y�ѷ��=O��4�40��y�g��&z��ѦV(o�� �M�5���j�������7��w�����/} :8���j��M\�Wz#ϲŢ�g/����l�wY^q
��<sz_��vڸ����x��w����I�%�f=�qK��w�����ך_ߋ�P�����I~ˡ��Z�p��5k�<u�ha)��Kĳ ����>@z{�<3��/d3h�7V;��F6�E�x��`uO���H�hUƄ��/E�69W{4���,�H
[�`��^~���~/>�R�=�/V��>% ����]J� �+��x�c�R�3�}�g�}C�����Q\�z{}���z��u���JL�C�=����>��G	<H�|eT;�>F�\	f������W���G�ܬ��߹zC� ����U�w��A(�����+�)��O�}�E�\�~z���T�y���m�v�*�:آ�-�����SNi[.�wz�����7�K*nr��è��
�����D��U�:6><���`RW�ԝD�L'��[]��\�([�ǒ�咍Ի��*\w�_c�^s��İ,yT;��[��ꢍ�Ub��߸��~��S��\��g<4�Cr�z�dV��"�Yp �X�j�r�*��kk}^�^`�9��[���OK�0{������Tg�pv��v�<�%�P@����;3����1����/�y¯-r�Ok�!�z��.�w���0�M�l��M	C�24����]�F	���ˌv�g����v]Qh��j�k$p�o������>��%�Ӏw��>s����
B�k
��Ϟk�u2����DϺ��/���1g;���r_͹�?{������ʋ?rˬ����K������q(4��QدȿM��f�{�׈:�L�RL����{�?i�a�gK�s��Ԩ�@uCn#��2iL2��K6=�R�轷��Y�O���^��m��q�V�^�݆9���i;�%;�=�բ��1E,��T���!0�ߨ-}r�{E�n
�koS�o�T�����'^�S�o��J�ڬ,~ǁ�m&eV'1����	X鉂�Ϣ�scdF'�]�����p��������!#���f���8T��=L��\U���J�{�r��g[��!Iӕ��s��:���2�(��k���M/9º��Id�R������w��4,K{Yw��5"�ҥ��Y�*n�Dzr�sHk�Ud�"%N����*/|��W�A�^�/K��	���B�2�b{�RaMt[��WyuX�C�{���|�X������N��i�*�d�~�����y�	@}��MeM�<X	YC/^m>��Py�d�Du1�5}.gJ�b�|h�ǹYrɿ����u�Oފ�OL��󆦗���N�w�}�^��<.�I=S(z	��)���B\�2��~}Y;�ܭ�h_O(Y����n|�Y��ڗ�<���+�ю((�1�������>�Qd���]욽���
��>�:�K�^=�҆{}CǬ7�<�E2D��8I�����-�"a�<��Z�\ǻ	�}4�`�E7�$.�j��������/���,�i��%�ov�4���Va\��w��@�>�q(�gj���+���������/��G{}R;=JW����M�a����=�����O���<� *u��|}hL>/{L�C���A�^̻8
ű�ev/Y�1������ߴG�^�j��s$�P�KS���R_����kF�{��'����u�����N(�ě�nS�-�fL�U�L4�/�Ñ�W5���nv��{�*�gfJq�1mN�yg��|s�����u����x�q���J�	�6�����1�Β_e��D��9Y�9ӫu���h�G�c�<�����շ��ˮ��"�qn���{���ql�_{���1������F k�#��)q�eAwm��� �WD�}�� {ɟD&�C�~Wrb�����1�u�BFCF	�<NO�`-��,��'�۞"̭��=\ya��	��׷kî9]�a?UHP��M���	�;���S3��':��ܞ~wZ�JW�q�~�9�:\��W>��r��y~7U�8��<k�4=[/�4�A[*hR�X��&�Tv<2��Ɖ��{8��܇O��'
�/����d:���u��E��S�.�k�'����]��w�VnM��5��./ܦ�p�f5�������m����T��^ڼ�Ίu}}5�%��1���!�@>W�Y���-plڈ�P&G�87����N����z�o����~\
�ʻŃ��=���w�Z�-YS��ωJ��_<X͗����U�N�h*�}�_�2�t�n7��B�_���3��;�:&����Nt���&�˘�f��8��`�K��q�t�<����w�z3��O�܍��A��xk���N�v�8��;3w ����YW�R���چ6�c|����g�ob�;�n�����q�A��$�8x��xh��Ǔ�P]7�$Y{��[{@u�k���ӧ���+�L��!��ʉ2�p�M_f_�9m��Y�/
/D�j�Kt�vlL�R�AM�-����:xq% ]0�Q���Yw�qM��ۧ~Ӑ�#�{#}@{��S�,^p��ނo1z0�}#=]�(O�!������u�H���V9O����Og��I���(J�csnp�9���}r6��ճWdT�lL���p7 �3 )h�Ä�w4V8���%���8V�c:�"��]�ˋ�W6��UW�Ig���6H#��@hQXċ�٩"�Ʃ��k�2���5�^x�I��ql��9=?t􈟴�A�聯fnr�<Gg���^$���Ǿ�������Z����w#���y]д�x�d@���@wD?]�>��ww�M��3Ӹ3�/'����g�D�ɻ4$�nn�u����樨������>�Qk}O)��CMnX�˭Lx��I�5�q^�.n����;���Z�:��Zcs�n",Nm��g�ڪo�
���u��/vXC�3{��Q�9>
�l�wY^j��<r7����G=�`Lǹ�ը�I���S^�ߢ���� q��)��(����Q߅�F��?���b����է��9K�u۝�TX�ˬ�Vz�_�O/4��t�Wye:X�h�ϬL���r]ӎn�����Io�2������n	Ѥ��s�����D������-��u�j���t�/5�G�'o>�-�dj���|�H��D=�����pԽ�ߡz��dx+�C��{��V�w3�B,����<������"�U=�]w~�(z)�q��U �i��L�+���w�O��z��9�R�jp�پ&�g6�������9����R�F���@7��4��E���{��K��3�~��
�Zن����+K�m(�kQ��2 �6G)0���8z8�/�!��r�������f�M���S�,]OJ�@�����\���^��]9�I�X��w�L�1}uR��4*3},���R����x�۬se���/}n=�/<�a�g���f���A��(���r�Ǻ�\�WW�]�����T׬�%����������1Ǭ���i[0� d�iA�A�={CR�{2��T�u��u�a�T��}�9�>
�_����y�Oz�������hOx�0rb����b&.d�i�E�=H<�$Т��r�n�Z��<\�.�����@Ԙ�ܜN�Y����u���O���DO�c�J9��<�%	=��}������#ڜ�۝�r����A�ϝ��k5z�Z�ч���{�e�$@P)} �L�f��iS��10��fS�{S~�^��k��d��
߻��u�f�n���,ز���5(��v0��S&��|o��;��+k����a5Yҋ���\�;������O� ��_V�,�S~��fe���N�tV�K�+���+5������֖8,��3}�M܁��P���L�S�{�^pr�{E���8ӎq�jӏK���	{���-q˕#^�KH��%�N�Fs��x]��������7�gcfdW���C�ku�]��V�'}�^�����u呏�Azr=�Bv�ދ
�f�}���Ll�{9�F��Ub�G?	�c������Z�`
�/|������z��/|��G<����?�����C.���2�ׇI�fѓ�#�S6Q�~%di� ���d\�S���z�7�}֑@�GC��Ee���r����=�C�}߱�:�Qt׉����\����p��_�=�˖N*	�&���Bz�\����ҟ�\/��qܽ���T�}�'|�9��1` 1t�::*�b�"�g��/yewG�p����C/
�����;�v|����Y�� �|e�0�b���x�����2<�}�-�Z��P�e�z��,ub�z�4(�!�cs���y�{������IY�ع^1�x�
d����jt5�b��d�mGE
��@Z�qT���-����6�Jl��SrN��^l]�QӜzm��n1u
c�sEi�Mw��s6�-ܓfU�\JzlKz�;	�j��D�|�e����S2�A.���Y6򔁜�����YK��� [$z���E��>�o8H�Oף���߻�4��P�=����l*�sޝ9�j{�Jْ���p=��@^*������yb��OԇUM�
���ܣs����C��
���.j yM|H���k4��7�`_s�ӎ]1eP�C����p�fS�;ŝ��7��y��3(tA<)T���=$L�Ru/���/��[�a���c{�ۜ/t����NJ�Idx���
�4��\���^�62\c3�s�poAv���f����Xܞk��_sԠ������c�t��тfd�a��n�:��lTϧ���η��&=y�ѕ�Zj�kï�ކ1?]�{��C��	�<����)�S @{�ą[X�	������Bvn���/r��u���{�C�P��ՏWNÜ�������S��-gW�{�fT��(����@���&��@�u�f���e���3>�r�[�R��I��Ϝ���n}�u�npvnM��8p;(�t;���pjW�G ���� �Z�`��w��[r�z!�V����wQ�{Njl���Rt�˽m����)@2V��Rӯ�{)�%��lނ�êNu��؞�<HmH��U�����D�ݥc�yf�y�H�0N�d�9,�u/Z��T�	���)��3���w3E���bs�˓l���7h>W�}g1-��9���0�uM~gF���3�j��ۋ6f��:��nO�s�>����ʹ�;��e5qݑ��|�\jʞ4<J@�pG3>y_Ve�C�ݚm����L�^��P:hy��_��k�W���?��CݑkQ����gJF��� �V��3�}��������!1�bR�O"���{ף7�>gs}@{�#޶=�ͻ�����*&v�:.�g����8p��G�\*�Q�:�����7��װ��:�v��:�8n�XG1��^���N���,��9 r��KCu�H�ǕXh�7�Fk��29���j���q�Y�bڢʜe�l�:����f�̂�|��*�dHn����~��QZ�G�;{�R�o�v�{(t��Ex�����9����hlC�,ҩ!���AL/WK�F�V㡶�s�4=��;�O��|��MW�/���J�Td.br�:��N��j�-H�g�2xF�����6rJul���jW!���W%L��3�E��"�������� "+�����E� "+�����E���@DW�A_������ "+���@@DW�"��������E���E��d�Mf��0O9~�Ad����v@������o��䢅
(T�@ �U �
��U@�T�I**�T�"U�*"��� E���IDnpE�	@UP	 "��*�%@ �(�* ���tQQ�;D�*�ٱ�͔�j�BѠ��+k0VcB�
j0h��	J� ��]�����JG Pv�@ X �Ll)@���!V�-"��[��;C�A��ѭF��	Z!���6�B V�� ���ʮ�X
يZ��# 1bR�͢$mf�IY�lEV��6���ѡA��+�-e4��E�SY[S$�-�����d[+d���X�	kF�5��U-V�Ep�j̆�!�f(UV�C6R�Lm��6#2ٕ1�K0�Y��6���@) &���ٛlƱ5�+M��֦�YV�j[43[J�X�Cce�� ��B�D� ��h��[Q��SIQ6�leF��-kF�Vƕ��)R�L�S� a�m)�-�c56�+al����1�B��Em�UR��J��
س"�5�B�5f���J-�lRU�6 x�@%
ICSh�H�m@�    ��0�*QF�d�� `�	�T�L��z'�4ђd��LC� 6��~%J�D0��A�M4224�ɓF�� �0F`�@*�����CA6�=5 �heѭg>[z/�v��g��°����/�RBI����a��"�����8�mQE?X���7�X���Ҩ��
������_�o�������)4�� ���@x	�  ��"i$����%A^a?O���q�����?���w`����A��փ_��?|�:^O���e~��&��w��~z0��l�)L9c`�,���:FeC��&AF`�RXa%^Xb�rb�����{P�-���yNl�s1@5g2��欽���>tk� S�i����+i� �8��[}����`.��I#ufغ���٪X�U����&��M��	*J�S쬺�X�B6Y����b�$�.w,��Wl��"����1��f`e(���`����!vJ�n�5PY��+(�V����S/j�;V-ȍMݰ(��#V�ՋJ���D�Eh�5����-5�	I|̃��� \T(n髃����WY4�xr��
���AGU�TӢ]�c.�+�n�v�ޔ2]%�ͼ�D��Y9�i��m���ـc����|�4�25�������YЭ�YLU��kqb� �RΗ&�����@�����wX�v�I#�v�3�Y)�4&���6�R������+�ʩ-S[�q����g�^V��
��M�QwՋ%pYifs8�,J`�PFn���.���NA�袴1�n��Q\+-U�Q2R���ӅT�M^:�٨�D�%�-�iYX�a�{�f�A���On�Go�d�֑T���L��U�U��&w/S�,�LWypn�mX{ V���.��tܬ���fl0F�̫	�we͕�kj1�ћ����q,��H��)| �hE׀�Z�a��Z�),��Zy���+�Oh��M�93tm��mVQa̂�F�fϥ��RT]�<j��%;7n��*�KFM������{�l�Y�K�t�AnA�>gi��i9��2�B�*��X#�y���
�r��x�,*�6Z�B�M��x9�^a��82�ʺ��#1�tTŭR��Z���E�ٍK��H����+ܺ�vZ���f��jf����+k�4�V��l�In����M83$����ה/V,(SxH�x�;���T�Rә.��>��ٕ4n�
�7�`z��-P�����Ԗ����h�O4j�Ue��֐���C���E�	5oJ��a�J�����$h��[ń',\u�.�l՘murTw����Vlc��+7��A�p<�.i����O�1ˠ�o,fivM��r�2�)�-�F˅Q�r����2�O&���ki��X�n�7j����v4Pgyf&�Ύ�Z�u�x�MW:o/��IS+�<�id�J��[#�,�J֚��j٢���S��/)'1�ȭ�*�]ګ�"�G�S�׻u���d��x��@�ft(�8WD�g����'}�ad6�Gù��J�V�J����,S:,m����뵦�[m-�zp���αv�[�E��*{�У��U�"�)j�w2�E��ZMX�1���˒ZPSW1+��n�����+&!`�c��o*7�,b-|�Y�y0a�vMҩ`��ʂ\YZJ�����W3-RmMN�Y.e�+f�E4��z��c�T2�cة#]�ժK��*̆�:��G�d"�͇u0�vY� ���fb̻�o
�x�X�,�ə�i���|����j3�X*Y�&F�mى	wwV��v�A4�V��{5tu��&8����
�{Yr���Z�k0]"�ڌ��ic]��4�)ۊ�7ak"?�Qz ՀM&���9���(�8"�B@�{�/Z���/`�����k1X��v�m]�,f���V\�n��.*3FJ�{�j��G�U�5��U	�j�z�;�vp���-���ۺ��Z"[��=ј���^� �y���飝��PV��1�<�G-$�E)�K<;-�v��۶��d��n�A�u�N[O�U��d6�M`\1�%�B��gXf�ðẽ����M`hG[�W���L��(�a�xk.V*M]�S2��UpmY���9�C�97T�vA˸���h��eEIE�kp,�1�"P�/5�n)I��+.X�҅�49l�y[4+�³2��ѐ�ڼ =�E����	C+�3�&�)轣��p0���V!�������^��h���Ih47i亚VSF�K�B��攱�,V��*9Y�2�L&�� IcF^�Է7-l�kbr��Ԭ���b�oɲ/B̓^M�yS+e��:e��XE�y��luбԬ�
c��g��Af�CHWZl!H�Ҧ�U�9`�<N]�}��`�����Q	����mi3(�%6�dYA�f�V�H��9/�i/	��zh��ɕlvp�I��˺̔�F�@測!X2X��i�iV�b����-hy�tc�p�У���d�⤬0�:�Fr+�׳f�)�gV1iͻ�ӎ�<�i�֬&�z^�Z�uekJ��[�I�%����ݫU��:ּ�kV::��D���������m�BlRM7��u�<�)��ڻ�71�����+)G73F�kW�����9�)�E��\Y��_�F2�tz�9�n_N��Ԑ�r!S0j)�9I|)�ݬ�誈b�آ�ד)�"�4f)�?\s6�f��	�'u*Ĭ�n0dV�S�w�!v�޼ߦ�(��ϭ���w�ҤZ�c����yX�@n	���o;u|�U���d��@H*YIR�,\��'J���Bd���,���֔j�iw�u�T�iX[T�dH,˖�z�b��@2;��J�5nTۋn�]n�PA���!��G�f3D���/kr���ei�1=�p^�c�c �$L�
mڷ����z�<#ø�@:���i�GBLkU��Y�|�ͮ�%VӍB曩*v�4���*�VU*8�n!4�=�v�1m�%-�`m�iH0F�mX�bE4��,Ɩ��Y���(к���L��M�V�ю�+
�a+#;L�te�kGfVF&��,�&[|��ƚl'�c{[�K(�	��%0��ؑ�7{WW�+N-L�VZ�i����訋�M��h����[*Ȣ%77�%]���+���{�c: �4�yS35�N%j�v���J�����ˣa��5�+�[�՗�Gi��~+U`0�y�:r�G3���G���2C೐��ok�e�33ni����
�ޝM�C2�(��
����I�ْ��x�ڋX��l����š�V�#J�S!�i���jԕ{B�o@�N�,�(�ڎ��SR�i,1��8�ƞ�*� �D��B�ս�p�V�[P�M�bJ����q͛V� "V�_Rkl��P�n��`�e�_5l�I�nkэC����Vͽwu1ti-�ىK!�e2���OE2g+^Kw��!܎��z�e�N �3r���Ki��,:�n��&*a;�}[x�i^[�d|�7�H^!�l�'e֩�<yp`IFKn����v�XT�U�[�6��SZQ�?l�DRJ�:Ӽ����)�5�Z����:�J"��h'��`�B�Q��Dx(�(ؽ8����`��!6��06Y�ZshC2kב�d��5{g���W�� ��O�Q�ߗ��zp�!�?���/�Z�=�:�O�	#���4h�}S5Iw.�:�(�*q_���  �G�����;64����V�/�X���.e��qov�0����L��;YЦ��!@讜x�J� ,Tv�s{���������cE�X���2�%Ӻ[]w�R���/1RWjU�3�m���SA@i��-�B�\�[L�`C�b��mJVGv&�v��T��JTޞ��S�[ܡ6���/{)AmoR�4��.Ѧd��fR�n�l�sE�.Q��/��K����������h�p$��`��2x�|��S%�C=]{��__'5�u��h�z!=J�j<���]`��7��i�%R��{2��KɅv����!w����Pg/c!���Ws���B�	����ǵ�"&�!�<�E�މˎ��B��N���Ϧ8WHlj4��Q>ͼС{x�ǫKB��ꛑ[��yױ�t����iU��}���v)]��^^0�m��;��å
�,n�oe�]�Fp��$�⩥���=ʹ�j�a�&Ҭ��
���з�0�T�kH����̾+ wZ�B����s30,��tw����B��N�I娨�f�
N��0$n�<�O�un�FH=V�Eu*L���+�kt��@�yz.,ܱ6�0|N:n�n�yn�y�ׯU�1P�}Ô�n�8���K���: 8�yQ�ьc<�a�:���o����=�z8�i)�Hb�JL�����`%\4:�w|y�p�Q�;�ӡ��g�G�� �ܸsu<O��y}�����YyJ�Ed����<Ol�]�ur�:.jP0�&�`&^��:ư:�`���w���R�6ok����^��X���F���)%�7��������n_=�`���$H�7O0����HӶ��Nz_]h�F�����29���D����vu*�\w�d��l�+3t;*.�s��]\�4R��6�+��(*�nb���E;�έ��ydܷã��L4��L.ҥ֎K�D�*��pR��&��#%B�u�ʆZ��F��4��� ����J��s&Ü�Vӧ��RvE31fK�H��H��ҕ���*X;c[/9"r�IM�/���o#��xi�N�Ľ�Y!���u�i�ܷ/ ���ډ���%��5q�H�¶Md�h 4ܡr������[Y��"�&|�h�jQ�"�IT�w+��J�ۺ���p)ji��}�H�#�n��B�H�rݨ��ʓ�,3(AF��O�'�\Y����6n�[��tl
c:s����t�ɸ�$5�8��Jr]t�/c����VEe��P�y{����/qfh��)J��gq��˧E��e�C���	Q��(����+��`�RP���5`G';�,.��ZH�]�ݝr�A�1�#\:�U�n��a����ݥ1�V�l-�J3���Kk�g'�еS�q�:S�zaͨm�z������U{v��R�S���fW^���:t��z+�ٮR��j[܊�����5�Z*$&+�f�x���{y&����C�D�<q���JI�-�lĲ�w'�&���S)�];��/����Y�ѝ�qW ���{;�z�]q��!M䕃�%�,J^P�[ /��,s[�]��[r��e%�F�
��mX�mJ	��J\��Yb<"�-e,'k�͸6��7�.Dݬ�Z2;xޛXz�D7'LR����w�B8�mh�t%�=&w,�g��+�=��e\]8��7��uB�CUa(���ogY\|�����]�WL޴��U�ǡ����S�>1��`y�|�E��+dˋ3��k��k�u=d��[���Y�mHP�f�jc��ȭp���w]7�㒻Z����+��MQ�k>9�[����XsRs���9��V��m��R�<�f��~;��T���~8�;�:�x/j����?��ˇS�{��Z[��Q�+���lW`7�j��=C�X鬎�,���CW��z6i��M�=fCM`㓩w1q���hų]�Z��dhl���B�X���re�Qk-S���5J���Y�h�[�tX�C:�n�w}����K؇'����uӇ}d䚌�Y���ZNd
����f�4�D��f�J�2$2���W!ImsJ�<��]����6��Nn����5�>{c�7��*���l�+TU�l��O7u�Q�2YP�.ڥ��up�:����-��Ɨ3#m����F�^��F�t0a�[�9KѶ^[�w�`E�gɶ�Z�y��C��Nd�e+�e�(���uG�H�����U0�2��+�����.��"r'w�V.�������ԁ�+!�׳���3Q��#�y����em��Ɣ���%a��k���Y���Z�7�<۳y��Rc.ֻ�JT)�y����r;�7��g^^��&[2!̢�VcG�7v_#���4�S&Gc�Z6k�k������7�k`6�� �S�.]�9�ܾ��lb�X�qvd[8[Ø�*����YtV�ޜ���oP���	�3B۝צ�d��Ww�P2��"H5�Te`�-v��}t�]I�-���[����*U)�;r����1�o2���7L�����D�U'��פŕ&���U�V�� =�����Ar\�4Ƭ��Ŧ��B�ٖ��FZ�v��OnI�+i�F��ZI1�qErCۂ��Z��Q�A�Fk!��h�a�g�v˽�s�s�
aΩFc!�}���Db|�V2�*qT[ٝ	���dn�ڊB�2�!\�Քӝ�1����}�S�Bbn���q�)VBE�'WFu m_5� ����cn}�R�>U/����ؚ���.����u�(�9G�
Ui*��+,��*F���PZ�R����幠B��V[��]]%��L�؃ѫ	�u���'-���Tl���|��G����Ʈ���0̵/5�o����;0��s���Ў4;:hc���2��`eO�}�c�^�e�<RL�qQ�ܠQ�쮜�^5������z&��d�}P�8�m�s�:��=��̢v릚-2�����k�ΐ�y�y�V�$᷅î��Cْ�R�b��G$�"��I$�I$�I$�I$�I$�I$��$�G%J�Z���WC������ˀ�������t0!D�m���/j)�&�<�D&m����1�
��i��/	�j�����n��+�C8�����vӳ�J��e5Y�V�Q�ܟb��1��� kAɶ��gcÚ�\��ͼ�@Vwd,���	q>�g\�[@t�u�U��U�t5G�թ���uoa�s7s^+5���t������[��I�ڐұ�0�Ag5n�~ý^͈�׳79׊}��������Uw��B��@�Y���G�=FT����,vVC2�}��텏2eK�ļO��:�u'<�I("N�v=��7=5��nqy8����'����yҗe�m)���������.����?��^������������A�H�z��A �Ш��=��'�ؠ�������߯����W��k�����6�:�u?[�i��M$X�9�6�+yX��k�^T� ��wm�gg�:�	���^�s��9��/�̡� s-����Es�<O�N��-أ'6�7t�e�i���9����|�Щ���+A�,���p[\�'6�����t*���#v�`ck��WY]�{٢�Z�)�5.�
�q*Ѭ+�aX���<4���,+�v���bY��!2�Z	�Pj̇���پ���4*�i�=�ض`�7֕A�Ң���-1��啸��]f9D9اV�0��e^�%.�D�/�ꐉW��̽���,u��]��lP��x�ڝ�\�'4�r��%S��C�Ȫ
�U�t��ヺ�gtDEz�✼Ŕ�<hͳ�F<՚��_>a��+���֍�v�a���@BUs-*�N��)e3G�݋�]���h�)��'���^�j]*�#�u�x�L��a'��J�vm�yݯ	��uJ\y�)L��1qsV�O������mγ�$U�RT�~�j�'KR��U�p�N�]��|�r\ �G
����Lݚ��hu��h�i=�{(=1֛s�̥�����Q�����U�ﲢ5�E�N��%�����W���Տ����Os!͹��MJ!�+��%mM�p\����:G���(CX�.��iL�{�;"�Z���A������*T+F �P��3e�Dd`wA��U��f�uv�8zhã�����ձ'IAQ�K~ӷ����x����^[<�uQ����±�S��p�зh�cU�;ʯ]��n��や����x�ҥXB�� �u�<]�B�*��M
K�݊�$�<�n�!�RrF�z���~7J2 �l��_"��/O��9+x���){�7V�6��ҫ��=9�рjËMb��` �n�A�m�������q��ٙ��C�)go�X�ǧ5�5Gdl����3�v��|�%�E�<���ϟV^=�S�	� ���Y����U���4q@d�V<|4�۟��M�؍��I��(��9�0�>�Q�k�mW7,	S�{�����}ݮ�%l�d`��T"���Υ.�u��-<Mb�0��&S�U�E`l�l��X�#��Z�.�\����땀H����O��oh.j�����,-<oP8�	a�uc�q���)�el�ͧrnh���;LM\�V]9�6U6]�.�QW05��py]f0��a1n�'���豖���=��Ԫ,����wf+�N���/b�I��Uw;mJ<�cG��vH[��a8n'�%bW�~�wYt�T�KiZb��L
�&�W{��e3�2�2�\�h�S	��<��>���N�m�j�������R�Dd|�t���嬶���O��QǗ:�);��f�t��]K�k��Ya����M��o��֜J�䉬Z�DEv�	�h������}�3E̽zr�������6S�_.�,sn_0�*T6��~5&�G3r�9u��4kU�<d}r�U�H]����u�I�e�i�R�̳��}[}�n����>-�7z��J�Y��.�����*�V)�D"�ٛι7І�ʭƛ�L�r=6��:yTj˶��Mۧ)��ݧM����o��a�F8j%O����`&jްE_Mu��VS�vi*��]6�[���Z�[��m��y�5*}�2'I�MW��n\�w�Ƌ=.p�2ƺR�^�(��T.�(v^H,���7.wP���a�[98P�n�X�R�&Y⍧u���U
3�u��h&�Ȉ4`�{�W&�>�e�l�u�!�%�����ٵ�s���T��ea��`����rt^9e�A;-\ɪ��w�d�"�{�i��w7Z[��&��d]�mXJ:����**g:��.�J5�X���hU�9M��z�:��ݏ�vl���1�(��%t!Zgg���+��5������wK���	H�=��jv4'�Y���Zm�+Gۺe��SXw�+��Ct��uI+�T�70�w�2Ɲdj�n�j��y
j�uH�iX��&EN�փR3�ӧ�M�{�h��y�]����iX\���`�nr0�ۮ���ܦ�6�;nā�Q\G�YO�E��;���i�N�^>g�}�AF��T*M�w2G��0�d��]k���K�p��a���s<뱸��b�L��2���].���']�� �AyZ뷕q}J��N��� �n��lp�\X;\��퐩s2�C����4�c�[Q6��$��'o0[�x��B8�Hw���� ���f�=u����,�����W�\�-�$� �bh�_eĊX��S�*�5�[L�.pP�\�N)���[�R�Sx�	i�̲!����s�0�6��])ՅșCiR7!��"zwlɓ��#��VQ����Xjv�����j���{�T��9�2e�����7OC��[V
�Y�N��]�I���v���낥C�ƅ 3���.B�C��s��N�V��ם���K�u0ԫ�����V�:*um:���S�faۡ�SY*u*[�^�5<�ˏ�ŋ�8(��LWF�͇t>�S��^f�8�o�\{/���c�t���6�k:�4����pT7a�<�Wf�u���.+36_'�/Dk׶_=�^Ǭ�σ<v!�uӽ�{b�Vҭ�fo5����.�e^�vMˋmWA0�y����,
��rRD	�ݺ�����]+9C���]���j�XO�CE�ma�*�2�-�|�N
i�hT`	u�|ub��P��W+2ܺ�ۗS8��nT�3f1��Gǡ4
r�"x&tܨ��Pw7�����A������8�t�]�G*a�V).<E�zd��p�VW��'r�t�у5 �0U��.gK� ���0�)*��r�G��� ���@e�9�/w�!۠�)�m�xp6j=��Y
i�V^��z��{������@S��f��B�'{k�w@�G^�f��7cU��R��L��{���ij5�S��H��/47�fZA���(�V/;D�34T�[�e��p��aʗ����L�D��b/:s�[\�S��p[R���<X���J�VCd��'bGv�ѹJ1Р�gG�蚣V+<5����Z^���ɤ��d��͗2��p���NFrFm!C��(.Ԛٶ��\VѾz���2O<�D�������U
��(R.�ڽ̩Zʺ���̸4�)�}xL]j��RO��g�F�p�r�}��ؙ2ܫ}�>����N����"�Mw^A����[��-e�=4'R���I$6��%-®ˮ�Cp�m�e]�Um�/R�;��"xf�X�5iwbd#G�>b�j�Q�-к�m=�Ŝ�z��*�14��zn�Z��c�sr�5F�Ku�����Y��1*wTޗ������\�6�R�����݃	��e:+����%TA\�j��=S�\$B�#¿A�"<@�M_���[Ξ��@����_'�4�u%�9u�S��ؚ뼚!���[Cu�"/%�9G��dg��6�>hˬ���Ƀ ,�[�O!�Rǳ{#��2���AO�Z��>i����z(K�!�7�q�1�:�'�kmC���U��9T0����5�,�	���1��t�ֽ.���6��n�c�XX�^�WQU��7��.!Pt�|Nأ*�[�u�t@J*�VԬ!f�9cܭ� p;�������b�X��P��޽�Y�WG��8@9����vT�q�F�uҝ-�:aX��w��Y���2D傥a$��]�x��0������jK�Y���ѐ\}_���l��TRju����)��{kX��2]2ji�1���l�j����2ՖF���0�#&#5���fj�5���5��j̭f���9�xQVf��Σ.c#DP��QLJV[�j��(�E�Ġr�f���իDӗ:��q��դ�8�5��Y��|&H����'�����&��q�]Pt�zJ�/%p�h�R�V�[f�2[�<%iZ�+�߇����BV��w�s�Tt|�/�'W6 �aM�v�:t�v4+s\��> �dI֥�Rҝ�&7�M�{	O`�:c����T�&�ux��/r��������.����+<��4n��s�x��)��n��f�>b�e<7��`�\.����ꚭy�S�3hyq�%nf�}ե���4��љ4�>���	-�4�7]{�������{�54{��7�uvb���RB�U���J�W�e��=�k�fl��a���S�_v�
���J'ں�k�Ҙ'+ �n��[�[Yy~#<&�Mjʽ�OOK{Ҭ��@��B7Y��3X�NL�����=<�a�K��>7�1�T3f��W8�d��4�Bn�8S�q�)}�/e���ohip�J��8�Ruz�������֢xUMj��/�(��ޕڭ�営�z]��O Ӌkݾ��P6b���ۆ��x�]����3s���-Ի���b� �RR:8��P���%�2��� ӕQH@xz���K��EV�M�S�.]d��	ɂѦ���lL%�t�j��زT����w�r��Ql���k2��tSwI�7�eǙ�?]�����Bc��<&݇��v �u�ɍ�ܾ*mT[óϯ�\����7 �]5�/�짗���z�����c�nΣGD���䃬��W�[W�0�Z_�F��n{[k�����I�b��5�9�Q�����\�3�<Il{+�}��z޲�,��y��V�Etܴ�;8>��\Tr���	��ϵWb큕xZ�ϳT��zn�${�s��R�҅N�(h�V�UDb��=mh%l�M�Ɵ��$ZdFo��v9r�\�Lk.Z�v;�wF�s�8��ʒC}6*�n��c�&ĥ�����+�SN�vIw� ��o/Xe5�6�v��XoV®��j~�����>Gi�x#�1��RI9�Kh�Ȟ>r�	�o����T�*�d�q�� �o��U[ם���a3��%<fj��sI+�Շ�pEc��pS��j���U,w�	�"�ي�.\&g�����N����r�kZg�	����K�����X2����	��������\�F��W��"�Y�q*dy+��m�7ι$82$ȶt������N)�s[~�Ssc�+�mn�[ZD'�8V��'>��p�x��gt������H<h�gM�\�v�>�Xn�yx0���n�}�W�`�w�a��]u8ޠ����UC\�f��-���4��8�'��x?Wې��!kVIo(�RP�ڽo&�p��YU���k�%\�͘���F�p��+vvJ�热�e���^���C�[�`�G�~��i[c����C�G�.�
���V估Ne�vƩ�6�S�^6�3Y��R��*\��T�UkjA3E��\�-r&���x�t��b��(ݮ�m���长@�o��ӟb�����Y��^Mz]��F����,�۾g��(;��A�a������ۭ���7�`���c8�j�i���^�o}��ӝ)&-U�{�s�7��<0����ޗF��rb}�M���*f��eru
�"6�B�3�e]��ۇ�m����v呛7��qΣ��`7�6����^�������+��^�8L��>�=K�C�"7w	T1|�h�Ζ�� N��p�7(��:+uϢ���Ŧ�� rN`|�W���u�QC���v�>��u��X�J��o�.�X���V׊K<'���+:���¼����rz}�%9
�v=u�z*jѩ�׹��s]�Z��=4�����G9��ken�IM���+3��P=�=�i��^���UM��be����'v�AN#&'����=��cM.f�VW��34J�q�EBc����;8���vK�.��K� ۼi�ݢ�˹J+�r�5����CP!8���*�9���&R����}��v�dOn_@��zK��jk�x����b��x1�{�&i������jG��f�w����Qӽ֜t��WA���
�5��;YikzGi�09�	]1\0O*i��ē���X���tEj�7S��ɋ�ȡ|�f�m��U�=�Ϲv�bEJ!��$.����An��^$�D8�M������r��1��.�"��]X�����K谳�0�w	�m+B�`�9�w��	��?��;T�Yo�8jQ�I�W�k�iف`rva8��Î�s�\$:��<�����ҫ:byɖ�;ޘ���(��eC�+{Q�>�"`�G������ɭ�Aժ��V�6(��b�x�T0x��Z�u�5��4hM�S����=��k�qSv���L�1:���X�+
�C���'/B�_�g���]����j���R��F��+��ыgO]r���~�\jV�+[�2�+�q/�n�Vp;�/G��A�r��k[P���k�~�i��i�hڶ���;{a�+�M��fY7���1h���u�{�kE&�"��tB�9��B���{C�z�@"Okwp�H�7|�L���E�'!�B�7]����P��W6�Y�-9i�u�;�7y�X��^���L��i��u3VC��xopb't��j����<R�א�O�6�W�kFc���Hus
zqA�}�fgޮU�6yL�dC�8���S�ú�.�����o��)C�gK���ă�]�;�۝A��ɺ[��P�� Ǉ�G�"�'��^�j�!G)���P���w�};����WԷJz��Д|GA�S̏b�	���n��ӵ*��tc��c��;����:��YͲBY���q�`�C.0�J��3m��w��ˆ�ՠ]�HV���$���P���Y֬�����)ZD֭t�gn�L���ZZ�l�o5���	�K]fh/�Ų����8H��ۨ����|n�����r��Gtv�He1{���:����xF�5ǹ^;It��G�҅��N�"�S�J����,�W�So�_t;�;�b���;KE.>�r�U� �҈a�r����	{�[$;��\6���������L��΋�sN]��H��)��E<BN�j����̔�YR��,ęhsEH�fU%�����M˽��r��8�VTwNU3�fՌTq�َNh���W'qs75&�#i��]�Ҳ�k��Rt�W|�>���K���%�>�\�;�I�̧�4�3��I�R`��K�+�c����N�F"U�Hz��i�'c, ���S�Z@���})��n޳c�I	v���E��Ƃ�v��Fk�x4v��s`&�&;VVیR9��b�
��n�}Ky���5��2��BR|һ:�#�SU�ܲ�ޒDؗeCi�h0`6E��JԻZ�P$��ِ����S����춷%Ԯ6)���3�j�hq�;=Ju2{��C&���fk�וyJ����rSB[��F�(�,0�y';�~�:��ɦ�c���fa�es��ڬ�ݨ�1�,�J5���"�fAZ�іe��*�*��
�aQLTT�f;�faL33ŬL�Re��MfD1SU�d�EGL�URU4n����
�*)�7UQDM4�"�j��)���MD�L�!IDEEr�(�O��YTjJ�9d��%j��H*=o!(���*F
��Ԙ�T�ծG�d����+#Xc��
�STQ����P��9�c�1��S��]C��G����n>��V�܅�g�Umn�:���xk������ss.�ղ�����e뇐U��Fn�i�v}{�OP23;�۩�q.H)������5�n5n�quͭlIr3����8�n]j�=�71����M�]��΅&'�Ѵx��ܑ)饙��x�'\`�B�м�A�JT(�W}ɀ	�){׫z]>��A�5껞qh�KԘ{��rJ�q���/�kʸ�[*�@-9������ȼe�b��>T��t�٦�\�j�v�3R(�w:��@��$s����fA5P%�`��m���:���޻��v^�}Jz�w6�J�r�:vՙ�lr̭�}�������>��Inc�n{5��u�R�/G|�
:���A�����=�91pӧ�i�_?Y27my%�=�>-��:��{��M�7�o�3�,Vy�zSl�������n8T���*U��K�IF1��6�ftV�뤑��_j�\e;O_�}�º{W_�l��)�<v�H���!yѼ��|˒L��$��OԐ�����L��s�:��vx\�t�]�^(��`"����G�ŷ��|����ȳT;�֭W@�ÛN�d�e�Ax�f3ͮ�L�,E�5V+Ӻ�x�g��Ұ�{��_OK�:[�.jvl���@�'G�o��ü't>z�ް�T5�˞����z��>F�穷��t���W��ډ�����N7���|wѓpk��r-�>�^GH�I�O9 �-A��Y�;��>�}2���w��sJ������>G����'6;=)f�3�hr�9�#�2���7M+:,���`.Z�\�'pk-��nm�v�j�p��u�[�t������i���>U=1�3o܃]��~� ���0�c���`D{�w� �R�>�{��z��>�2�)ϸ�+��9���7��k[��y�~!Ԧ�����]���� q2��%N�8��M��})�0���5�f�����_z2�<�GX��� }!J�'R�R�/RH�/�ΰ�5��B��:�|yk���{��>������x�G짲�}#�%��
w��>�G��x	'�b��z�o�p���~�q��P�!��!�C��8}"}:��
�!N�;�7��g������G�R�'r����L5��!̧���/{��L��(w�y#����=��}����J�O ?[(��Ǯ��i�t���2�d�4o��
�nN�*^L��2�dUY�ek�r(����M�E;�����8ߞs׽H���>��C37����L�9��;��!�<�Ԯ��D������}��?x�2��`��r!�ԋ��ǨB�}����N���M���k�7y�Wu�}���{�%�^���D�ĩ�y��Jn5!H���0�w (b�v��^��y1���D���O$��z�:=�uq.���W�SdOP��|���^��<���7y���羪j�)��%5�S�{���P���G[�@��	�s�#�&���y�����8����R��G��VA��짲��d�x{ܽ@sy#���8���WY�o�5���� ܧR{�/�/0�b����J��_��T��ĉޱ {�=�������5/��s�w�z�3��z�نw�;�o�C^�� ްN�~ֳ�w�Ǟs�]w�ԉ�<�9 s)䯐zy��/2��솳�_#gx4���{���\�޺�λ�� �ON�S�:����CP�Jw��*w!B�̜���.G����}��)��O��9%]�����k��To}F�>L/p/3���r�W��I�~Y���{�Ws�5cI :dU$o"=�Sq�J.��kp��(�>���S�C�8��]s��Mw�A䧓���u ur/�o�s���>�=���^%�=5��k[�7�Ԧ����d�1��M��{�%��9s��������뾷ঠ7+�	���%=�p���7>�o��N��W#�p���!�'���������^�j_�x�0etB�B����ة��>���2S�x.��OeH����x�x�}��B�����.�p�t�����/r����O��0N�toP�����;�����~뿾�C�9�5���	�pCϘ��/�.Z�8��B��w�:󳞼�����y�~��=��S���0s&B�܉�s��w�
j�.�x�8��� /�dl�}_6�z@@����
��S�
y�{Ї2ps���� �=��d ���&G#��S�����Q�S�8.�4f {s�)�w!H{2{�C�<�`Ms�R�z��������wU���{��p<+�x'u!G��ђ'W[����)��q)ܽɸ��۬㻒h4�e`l�e��_�:y�0Q��dY<h�sz�8Т8�>bn�.��緩�t�9ݸX<4j���0�����77��Ovv� Tl{  {�Y�r���b���q��~��x����]@����:���83vwߟs��|����/P�C�]}��?K���1N�u>A�̏rxx(�ã���}յo��6 �#�s�;��;�>���G˃x�~�<����B�\`��ם뾅���v������@�I��q��}����Nc�$8�Ԏ��{��O%!N�߾{�o�{�|�=x�}�����>��C������A�p%y#$M�؇��N��%��^_s�����P5���� g�>@s!B��V�z��O w+O�v}��q���Bv{לk���z�Ġ�G��~��;�<���=�7Ju)�=�<��}��Aq��u�f�޸���c���)=���_�K�^�N%�C���Ww��ΰ>����}�?s�ރ���{��5���אxG˵���|�~�+7�yY{��0���;�F�y�2���Xe�3qE�ޚ&�9�*i�\�U}��'��ח��C��*#d���U���p�������]�\�~�3M� ����9�!Dk�ѫř�2F��J���+2�A|��i;�ȶ��׵9�}A죝���oͣ<�%r<;�k��e|�~�띻�Ng�ko�i��,\�~�zo6�&+�S�<��2�Э���=�n��n�J��t����9wYi�*��i�Q;��.����gGNPY�ї,����F�X�u/�ެ��z��**�[��>�ؽ��b�/�S���Wi���÷2��Z�F�;I��W_�z[���ɰu=U�c�4�)+X
 k�H�r���n'����_�=~�����Y>v��=�6�]��b�l��T�k�S�h����J�O�d5��k��{b����2ӃY}�-�h��l�M���]�q�\�4��~NΔ9b�zct�@��q�`�ǩ+&$*�1=y�����f�^\�s��&�/2���kK���ї��i�kVrS\P:�&��<0�\߂���˓�k�t!R==�gǟ���ut����o8jr뙀��B��)��6��n�k1�f�v}�?�i��gc^\>�y|�L��]E��D��:�Ym9�}_Wդ�#�~��S��cr@�5��IRV���=�~�3��*� i{6�TQ���)m4����ﾓ�ut�����T���ϓ��vqy�#D�{b�k3�u�-Kկ)S��Ph��ݽxR�V����/��%����v%�^���۵�{ o��7�c# �L��t��{N$�#����4�\b�i�FL��w|�+u,�4��Sy��9�Nb��7�OR�X��6�c���Y���Pޘ����t��˨;�ЪλC���lr1V*�w�ۦ��<��̗��2�_b(��B#���Z����Ltn�g�ވcux�c&�̷(P�O����;��`�)�6�\�̓,�T�:��m�è|��s�,@��B"s�um�8>����|θ�hmL츭�F�0����˵s�lG�(t9u�ds�n�t�١����-�ǰJ����L�s�H��	�D�M���sqtox�6�o��:uĥٶD���Ōi�H�{֠�%o)�6���u��B�]3Z�K�K �Ž��Vv�:����M'L�v�F޾�{4���ƻ�y.��&���S�\@�2���
=�ĞvX525/.�+kI�n0VKS�H"{\;d
X�P�B�U����%��3�'߷�gr��
8��hv'�lI�M�]�Z�W®���Ķx�J�:����8�����Q
�����7H�Bg�VUp��	���c��5�Z�_��N�u��`=۾�Q�E�_P<m*�`�� ��*F_�2�s����mL�r�ob�L E��-7l})O�tø���n�B�Ô���N�	C-�ʸـ� �宗������c�R��Z5m��X-�vu�n8���� !�26r�M��͏w4��X����k�qgT!X���{m���)SH�p%
O�s�xMjL$r��9�z����^5р����d]|��w�	���8���z�?�~�
*��>̨�(��3 �J����(*��h&"H���C��AT��QDDT����Ƞ�-�nM�$CDI0[���)��*� ����1U4ĴD�F�(
�&MDR�!Q$�TUn� {����Y���C����,��5uo��j�(�)P̏]Y�w�bn/�W��i����~$���|�̅3k�f��������sZ�v��\dT��-��M5u9D7A��M"ѼQ[(7M7��n����8g�k�V��Ūgm>r��e�
:�^$`�x%���{�~�O��|�s����w�W�jKm4�SH�\b�t�؃�/15ҡ�h5�����
|���{<#�d�'v�xV
~�����w�ێ�4AƋa��[ϫ|0�!�����eeg1GUg� v[�����X�L�Mn
'������g>o7��?����6���eME�����ؾ:�zk"�!m�����z�W�+0e���������qs �ެJE��`�ͥDC�U����+3����uFՌ��}���Y���u�ʋ#�\���}�I�O^=�L髯�G@��v?H�>��8tq�z&���+�{7ܥ�>�u
ʻ��dY7�B�s�[������Y~b���b=�����T��]~q=�z�+�y������I�������]cNW!^�b��*Z�^�N�ege�&�"Ɣҗ��@y���z�*#��빢�Z�
��=^d{2�!�J�⧻���3�e	�h���W����<=O1�T�/Lߨ�nu��G���3M<����+t=h�q�vDZ��q7|�\Wt
�u�˔D����5i��wq)Q�f�O��_s��2��7s�t��^��x3�.FEaV�S�ñء�׫UKl�*��j@���8l��ĥ=���3sgFm3�yb�C)�֬�l/oƜ���t��o�nng���r��K>q�5fOR�Y�R����Z�qo�o��9�t q��+�X^ڕ=.��5wJ�R��L3E�Tѳ�]�?�m��y����Q�N^Xc���k$�	�}�d``��K����x
��|�ॲ��K�ت��+̩������o�ұ�\D����^Lo��&�K�ۂW�7�l��
��E3��w�z��(AR==�͒�����ѕ1ׁ�C-�E�p����eR��\w�]/!��b[�&��>C�����,�(��-sN�	�u�/Jx��{�|����<��J����V�j���[V�#�fZ3����ճ�k�?R6������r���ƽC���z�S�d��71�&���[h\�1�B���-��ED��&�f��`���X> x{�|����,�ؕ�g��N�DR�Uw��t;)��K<�|��h��Օl���Ǣ�Kp��ݪ��F�W�R���Y�l������R�{y�7��g# fG�f�
��(���Pfw-�t+���n���������/�j�%u�"��ދK�vm8k0�-<���W�f�y~�}x��F.�#����\�B�MI��啷��=Ӝ֚�=�������j�e"�!����N�5۸��@�{�3�m��-8`��I��@����(f�z{	��z9'��x>u{��}h�}"(����%�p=B�p�O�Xs=1�O�)]N*�8���bM���a���F[�$����Eu�<��=��b�]�39C�'=�=��ޮ���[�kP�"]Nv��}�ރE@���ywv�Q5��Ǹ�?d�F
Λ�&�%p�H�D�#�+��Ó�X�2�7ү&�+^���iX��L���:񊾡�^ST>��~��׉��"i�u���s\�Vs��ቮ��QD�S�dl{�a&�z�#/Y<Z�ej���o^+���;l��ʍ����������暜���}�=���D"�޷�Ln6f�ϊ7	�]=�23�}A����n�v�λ�/��[�W�����5�/K�}��)���������{�L������ϷÐ<^հ���硫�"-��/&N-����tD������{{�秳��S���cW�lY�?�s���CW��h���.NY��G�� �@�=�]�Z��k�L/�{��a��"�/�O��mpm|wy,�ok�+	���xeA-:�9��Ɩ��.��vf/#��)�)+��n�����ݦ�N�s^�����N]�黝�s �=΋������5�r�+��ʋLJ'��WbOSp󡝸��Ʈ��e�j�v]���c>����P�J=��E	���Dp�ݽ�XȞ��t��/VV]`���k��P��~Jm>ܹ�zs���ͣz2��5ә+`V�3��S��!�!ߢ��p۸�nx��I��G�xI��q�C�yOwv�v�b��;ξ4x�m�3���R�.��ѹz�>T�_6Qb�M��h��r���p X��<2�m4%nQ��%��� 	�M�=���}�w�bXeE�lZ�Z�j�|��>q�ۢ�
��-��F����j�Gv�[�"����<��fB�h�C�+�T��뻞��7�B2�/��QW���u����!pn�7���S�i��$A}ou�S�^�O��������dd^����D�c;oX:�m�R/=sn[1枽N�#����o��ˣ�u��pSX�V�ǳ�'v��Gye��1N��>�}Y�H���!�A�ѡ�r��vS�4z
[���Òԋ:�wB�s�K��-$��r� <��%�V�W�5��!���6!mR�n~�;���uL��<�f�k[��k�r��wc��*'��F�p�FtS��3Nv~��õ�3�z��omO|o��mVl�gʹD���';�,]BK��t�Z�̐�\���K���Ђ*�I;3��]�tnyѥ�{[���֬���ܑ�C�
X檩��.lj��c��7+-�����	���|���ڱlEs�X76S���O�V@�yO�&1\�����4���D��μ�v]Gǅ��n�d�����ˤ��r�n��4J[��Uܘ�+�]������`�f�_Ö�����E�w5�c*U9��X���'����6��Չ1y��a��2��}�����bs_kU�}�8�^�=Ν6�]��*��g-�
����G?\aR��v��ʵ��-�oC�v���(�2��Lی�6���LX�Nt��_*j���T�%Vnt�����'Qэs���Ya���2��"�G�
�R��}�`�����\�U�;v�M��N�:��� �[�t[���u^WH�<��@*�Q>�pu)���khͺ{�Jb�j�eV�R�nS�Ɩ(�Ԁ��H%Ev.�*X�2�YX��UO�^�sg\��r��'v����v-������rU�7�aRvԤ��|/,�x_]%+j�R�.�7>d@��!(X���F��M�8:�ŽpU���՜bH�}wo1SgT\�^��>�XXp��uI�ޣkL�9^�}Ҝ3Fm�2h�#x�R��gn�`�S��::[�p�c���@��X�7�2�	�z1��A��o��k�]F3��=�13};���]���E,;%��^'קd�X��(�\P����e�M>���H57J��N�q���
��B�V���(xW��%N¸�����3���L8�<�X�.\#F�*N�O��U�T2�&��[�p1$9��A����ՅP�DKA�dKO&8�4���1CTST1$JAn���VU�r
��$ȷ�MR�M��
�� Ȫ"(�(���*��uc j��AB�44�U%�!�b�������w&�CM!BPnSR�)j����4�T-֓PRD�%499��~����ܵnr�6g2��tG��pE���ű9�w/������i6��Gv}���/��2�.���r�N�󚮍"z{q{k�e;�_�djo���P=8%H��Y![��yu8�uE�>�,fLz1z�<��^js�nK�-��yn�P�>�nV��e��z�[M��M��ǣp���d��ǎ�U������]v6��X��Y���q��]\k/]r���4ͭ����5���p��μkFkr�磏3j*��4�6�c�� W+��Nٖ���V)u���k���g��Z��`�5��Aɏ652�X�BR���y�l�8�������>�o���w��{#c�`�1����td�r|�uW!Y�W���(��34r�eվO��y��'Gf�^m;���\��f�[��ᢻZ��_P�r�|y��P/'�i[�-�}[]����V��қ{5O���~�x��^�qZ���1Nx@�ǝ��U�.���7x�LX��R��T�yz�����,Bj䌖�.uo:��FQx&��+��a՗8]w{Y;wW���ҺT�GLE�E4D]c^��^J8fu��c����]�+��ա���f71h�76�u�������ݽQ���w���|�j_e�jl�M����f�͑Y��}X��S���x�}�k�F�H�*�{Cc�1�o���;���nWi����QW=��)di���x����"�}�ֱ'�\K��Υ�����F��˧�Gms��7v�Kk������<��<:Efv3�T�RReM�Ɵ���*U�����3�c�����r<�������(���z2�`���8u�]Rf
+�X��#���xP�tx�z���+@�7|7zl�3рl�*�ܒ�)F�5B�MbI}�=�2�[O�Ǭ���c-�%�I�Ʈ-XW�UdI.�P�B�k_V��x�^�ַU�ى�Jks�;�}�r�:nvD�+"'��Fib֧����;����]\Ո	�P�7���ڶk�h�1�g+a(���m78�=����"�����c|S����FyٚB�����[��i�:�]I��Ks�$�>/+�0�8��Y�5��tDjTD�#���Y�$R:;,����w��5c:ᨫq�ʔȵ<��������+i�7%v�iq��s,V-�ǯh�I���vqR~�����(ߍҳu�:=�d���;ϯ�b�����q��K�Z��#��r�6���1fg`�޾CHܥ���`Ed�
���Z ���g "�g,��9�R�~3M���6���1���t�ޕ#"Ql�'�-&��\E�O�(~��w���l� 1ה�U���::�L������Wb����%Ǽ\ȹ=�F��t��� 7r�ޑpNR1�D�n��E󷶚��\myϱ:=J|t��b d�3��r�85���Ҟ��.����o+�[	�{��}%� էL�0�b,
� �O7��t�Z+S��4�W�������	l�\����:����_xxxAT�c�}S#g�,G�
��P�	�Y�ʆ�>Z����ep����ɮ�@O�v�>,ո�R?I&z�^?v�Z2�~�54lk�8pǲ-�;�΢�jt��H�&-�䍁�&�q�}1+$o�δ�pCg#`` ��8++7Ai�e�뛾�����%I�2�|��8�
#�I�q�"=N�
���\T��Nz.#m��C�8� X>�_��7�>�~K�ohS.q��Dl8P)Lc��u��v$��C����>�\d:3d9sИ��3sk��\���B:2<��$���@��j�{-Kɤ�G�tj����`s�WX��8�ek����}7sod�`��fPy��6nc�/T�=Y@v��ZH���/Qn~�����s���~Y�D�������f�xK�;��(-�o���Dd����C�	t���A���=~�� t4V*���}~6)�Z=gF���Q^#[3=ޚ4X 
�}��3��B�Ї�-S�������_�Dj"l�O���$�q�	�^V^��ZF#�"�γ@���c`�8Q����i��!�: 0ƆO�)�N�D����_gh$���(q�y5V��>V���ŏ���o�o'�*�����&����"`t_��:��F�Uo���I��&l8Ј��C����l��űs�U'�!U�͓'Y!��7�c�i��D���g��`��K�=�x!�v��sX��o�2��ȭT��Yl�����V�K���=�tC��EB�eD�����Ǒ �Ï$}Q���ؠH,�j�"�A�~��;$�y��a�8N<}�.C�j��`MA[n.vmrg��}��`!T��@Z��5|âlyЧqsիS�1I�B�(�D��T�U�Ѣ�`�_�� O,{��>&�p�)�K�����4xU�&Ń�a����]8�f�ė�(�9�F"(k̃�^Sլ!�ș����I.t<:)���c�:o{ԙ�5��a
���N+Q����X��ޣ���w��=*iQ\iF�@�;Dl������y��|�^Y^�7Ktc6fv .��6|:v��K��KDSa|ޗ����I�hêji�wTM\�8���qV���xY[���__�6:��}to4K�����~�� ��M�*D�<w�d�u�t|�_e\���5�ѽQ�PX ��6Hl`��o����>�#X��Z�^�Z��
�� V�@`�cC�t�z�Aw�5�ȕs02���fH�=fv1�*aSSx�v�rѬQ�6GIp ���@�{s���nt*��1ן�xhU�x`����ó��s��ʠ�Bx��i������hV{_����|�jC��V�V�ɘ���q(�_R�N栗j���0(h�(�j��
f�5�P{ƛi���g��=6\7`D���\h���&���&i�{�f۵a��|��K����C��9�Ma�.7?W��[ƛOD�>֚d�; P�K��ca���r���S�$�U�9��Ѩi��	�TU��x����Ǽ=�@Q`׋����t{��־�Z�GW��~�\�-5]u����YB����e5PQ���Ã�0*r���|:����F���p�.����,�5Lp�r�oPH��q�1H��@�jFwm�^�!aL�#	�����̎T(�;�'jw�s5I���*Bg$��t���AP�M��vU��Ģ��e8�m��
焿]+.����1J�^�*����������&(�G�>�X���(	�S�.g������p�76'�rF�#u��j�:�F�{hjn�9�Ҭ�7��eh*n��"��OakV(��c ��9tu�D�x&v�&L��y��5�y��|�8�]mA�(�O\�$Ý ˭���:B����3�X�JCmu�O���P��\�EE���1A�G��]�����x����۵J��/�f�
��h����t��@�Z��s΢\$YnN��ZJ�f�'V��<����eD��l�w���(<�C�U�x�� l�?d�+%�w;JŨ�m�1h�sE�vjP��cc|<ȼ�v��>;�)�̛8�o����^���2u��Z�{x�c+��
账3������P睸�Ȇ�'q�hwj:0̽\�[�K��`gBz��_�]t�7!�ٮ���
��Cr����W;n�ޫ,��(��{Ne�I�8�>f(�L�/�7��R�T#~.����~��{��@gkٚ�����F�2T;5���y�C��%oW�dE�'�N��R��nCQG�(9:�4/]�֗1�]`l�
��Jz���Xܝ�}F����m^�1��y��7�6JK�5y��֙ji*�=iΥ1�]hewnғ�m���R�uJ���u�;���!�ZU�Y�+N��ܸ��U4r�%����\�]�Oy~+)N[�)bU� \f��uY�a���ȩ��!�X�MǂE$��8�⃺��x�����e�71�.�{�<ymŌ�ˇ�G�  ��
���$MD�PqTD�4�#N�\��5&J�E�2$�X�h�ܙ д4�	BS�W7���2�)�b4 P�0*��"��)�!PR%+�!*��7#���(�&����[�ˢA� �EG��g�T��퉞�쌾�˾��j��R(Z�{�A�]�~�� ���Z�1ѲL���*0̋"l�$gEWHQ}�)극*�����ѐ�虩ˁ\I7�A#b�e��s=ϗ@C���,W�k#კBT5��;}fצv�X>�*涇����k� �ƟPD
gb��́���o�cɸ�s�f#����u�#g�Q�H�������3��2j��ꊳI;�:�A���U̝�1���"O�'���<���58������瘯o�B����Mn������ �U/�of����k�$��]��
�g��(/�,�Dt ��_1c�N��.��7T�z���+�o�+�x!T��EK�^��3���oyu�{k4����mq�d4�Z0Q��}d��:4f8Gl��C�0�Lz5�V�:ġ��X�Y�.uѣ�q�
z�v�l�m�͠]��3�@��
��g�1�R^絡\|�<��V1��*��0J�Id�.^_�tJ�C��!Me(������`�n݌�X��Pv/&�v���[t+�6%�d�̅*(318�v&�V�b�� �b�h$؂�b!��>,!�f��:_u�`
�b�
� R�p/j�:�4z.��,�e�������!E��5��q`�9h��<��>�������� �〇5R��j���W������$�e��ax�ص��¥����b�h�o��5���|=��@�	����c5�|i� ;<4W�ȭ9��´�~�f�g�
����nO\�-<7Y�M]:Hm�x3�_5�`�O/��76�K���ݰ���V7S�|���v>�f���u!�'+�՜���2�s�����I�8U̜�v'K��z!���v�����k���nj�Y�g�p��M
Yz��؇}=,�eGF�q|k@H��*U
�m2v�!Z9�OX
�py��6\.���Ό�5~hH7�=k[QN
� lv ��v�AW[Gő|p�N#�gr��~&㣢��> �	dt��**6)�:H�k*�8;:"�f�`U��d�qcV<(�!Vm`��O����sR�@�>�1&v2��L�Wjmd3TE�B��f�Zz�@��dnƅ��\H1>9��,�NY�Ed��b-�n�q���)�j�1h�o+��Cn���VQ4�W+������E�]��䭓;���b���_x��o-��5���.��ж��X����i���3��5�p&�׃񺜨'.+@����L��.��7� p8f�\kf(ȫ7��F�嶹�a�p*2EmW?,��5ᰱ���49ϓ���Փ�D8�.D�ء��r&d
�(᛼�v��b&&�,���E���g��hU�֫��Y2U�6���6���2���h�R���:�ԞI9�\�Q�5b�o*T8R�J��*�Z٪��1A]2=�w�x�5�:�<�e��<��/���%F�kuZl�P.͊Ђ�~�CUF���ʡ񯰆ySl����/��O��;ܮ?f�-�.B��aT�L?f�73�7�v�D<���j�2�KP��|������ڵ�Mn�����:�b�妢�؁aȘP����Mk�gɞq�\}��*Gq�oƴV�xj�(ѭ����/���\(�|<<8u*F�i�3�ά;����LD	E�LE���ȅ=(��{�^��֭&#t�P�
v�[�C
��J�4��Xe���� `�~��h��Ihj*�|)=D�tFr-	z9�o�uһC��nݛ�L����0�aQ�v����j�Y�<rt�=<���2����z�Or�{jCb��k?/�jk_*�ƽ_k㨹G.��$6�V��@�+.F�bb�eb��w�A֙����~��pO��)k	ʜ�(>[�{9/��o@<;�N�r��Žz�W:@aI%�;݊l�J��vy%�f�j_���wm�d~P��O�K`�ªi�J����;<�Ꝯ�G��LV�`@
�-	����eDǳb(�*i=�PƑL�##�zB��2�~�B���>��<g?2��y�@��q��`D,�4T�$��1����;gs��A��ur�\�Qٲ4
�Ɖ>K� =�(����]��)^���8�Fto�f�V����o7Z��)��V
��z �!X)W���� �ڸ6�1��(Ȃ���|�,/�)�9pEI�n�*�{Mpa�K�'�^Ȇ���ySSD�y��bQ5� V��U���=� ��L�I����:잵mn���r�����Grn�ӵ�Z��TSC����̾��{d� s4@��Α��A�&��ңhw)���o/9/���� ��VI�;"�B��Ď1
D���MZ����q���>�q����%A�d8�1�t��O'Gz���d�'n�9���i�/�5���\�
��8��gG�l`P�k�	�Z �ȫB�Lhh�uM�ʹYή2ە D.�f��n��q��ġU{�7��H����3#�Y�rDi؝*$Hg�V�[����3¸T�ֻMxX�VoW�B�K�x����#��N�\S.2�R��F�q���� �6,�b�n˾䉏tH��!B������#p��;7Y	�.	��j_Y��WF�DDj=��������:�<Dc��b1��m��
�u��,V�&��C���$�EU��o�"դ�ɷ�ΗZ��cӋq����U}9'?T���]D.���ЬցC?�]�
A�Q����p��(xW��UV��/���2��7��&�����l��!�k��O,f�:+E=?�@X�bX.�R놷����}�U��]�+���G3Z:�X�y1��fph�~��:�~?3C�p�ж�����ݕ�:�۸�},�3�\HeD���L�5jDD�"���O�u~x�z ��h��=@�p���jH��H���m[���j�G�8� D���ج3�<0�C͎���v7H�8  Ԏ�ҠdM�(��n��7�E#����=lp���٭�D��
��.���e��ж�@�;�h(- �_��Z�F罖|^�~�M�I�{h3�!F�0=2�;<^���$�4ze9 �cj3�mG�6���
�j��T�N�D���Ǣ&�a���R��OC�)Qx}p�A2�1:��1�W��t�(����i
ț@�F��Vw��4+��҂�5�Z=�_5�>�M����!����j���l�G"����	ɍ$�"B���T^�O�:E=�DS:�"0�D-7N���FS��g�s-��*9=y.��dv���A��G@#H��7���c�v�=� S���"�pv(Q�6&���E��!�%�Y�!�Q ��X�rb�����=3
Bꓹt�ڴ�y�q��*:I��͘�6D#!�2d_�u\HOw�1eC^ p�x���cؖ��u�®��IұQ��v3��a��Ad��P�w�t]��������[�{�lo���r���m�9����=�w;B$B�M~{V��R"���Ӱ'�f|H>��ѐ.�i3X">��w���۞����ܺ�JУ|2Txэ>��e��W����}�c�5<>�o����Q��ꁹ��s0�bY�b.��$���4���SB\�y���>�M�@�N��X����M�S����d�_A�;�w���:��hOW68F�P���ۼ�^3�����OdH�D;8,0��j�#�t�)�̝��w�Ay��*
*�i�k4耊�x�ʶ=���y	RX����6�����9N��tF��*
E����� �܈���b��]lLtv�ب�?X5E@1zOh�?�f��
��^��4hU�$}��iM���fj[ݠ')��P:r��/V����Z���X]��7bu�i���&��,�}z�·,�'��r�z�u�ա-l�g��əE,��K�'9�Fv���N���O+����u� �,N�)�9�S�d�e�E��2�2���.a�٦��p�΢H�Κ� j�WP�ǘ�����I�^#r�Z<lur��Z�Q�]y�똷:	�;���2���\tO�%\~�Ot��٭��֭�;�b
�Q��N2n�z�d[b�EvU�\F.��X���Q��2С�y��[w�����W_dj��H֎�t.��`���L��\�F����*�wة0�,q�[O��^�#Q�X�b�Z��B��z�宺x��B	wԓFW�yjPA���*^u�]C�:8h�P<�հ��#]�$�NA���T�=x�,ZY͝V�	��NP�e�P����N�����.�p����+�aʵ`�I�wy8�h=�&��Q���H�l�
)k��� �ڊ���V�O.��޳+JVم��4.r�\!wc��gFӬ}B���ئzV=[}M&JL�v7j@�ׂ���)��W5��pqRNx�;ݓ�P�q߶�+����ŷĹ��32m���kwW!�Σ#E �q۳:e����=kDq�fk[Ѭ�M�S�x�X'���ۯ� �"(T(=��( �,�b�#)M3�����n�r�@%f	�Pn$�59�
(2�Cs�'$2̬V�!���eR儥e��P� d�(䚴TU9�U!�$���&�i�)�B4%&� rAԥ.�@aF�C�w��tk�y�9����y����mV��'(��Q
#�U�[����0ݽQ�?tn=���!����Y]	pv���x#g���{�
�숝���|$LTS=����1+oS�ɋ�iP1i���xk"�*ۼ>���y����HO��
6:.i�,�H};H�X�s�oi�:>�爂����hp� r�h����3�lft+�\��2�	���C,�"q�uDV��k®n{;[��q:3g?��z4�/(� ����{^{iV�4u�p�^`M*���"�
��>ʽ=מ� ��0>�΁G����ǁx^���o���{!RΌ�BP�f�ł�;/Wu���Gܾ(?���5l�B��b��U�&�X����ܭ�M�!'��J�Y��=7��BJ�I�w�][�۩}��W<5��>9~#$d�"�9 dw^���Z�}Ȋ�a��hp�x�h��^���\*�O��zY>ٛ[u�t}�Z%#V�8�����2*ͽ���tN`�}صÇ'�,FG`�26��Ar%��ѐ��(�01�[Y{ݞ�	�D2v::2D�$$bAXX{F�f�&��%���� �U��(K��L�g3-����Cޅ�РTM�$}!��A���A}�b2:	r�;�kr�5��|bh�C���Ĺ����NġSmV�p���FLχ�|%x��yp�h�0V�\���MK�a����;� �p5ʥx�ƀ��@�|-琹��I�u�����^G8�:��L��w����IW��P������Ze&Œ~U6��Z�Rm0�/%^N r)��C�q�W�]�����V�ܫw�~���xu��o�/Hl�1�g� &�Hh�ed�r����Ժ�w7����G9���R�g�|(|�9�������(u�%�*b̽�ʨD`�]t/ϸ�1�i��YTa�Z��G!a�b�OC�*/��n�v�}�~tB�Rd��
�oqV���U{Z��~}���,b�AZ8����[[C�ѻ'�y/oT[���W���ST0�@;� +'L������}��K��ƈus�E#����Q8�cD�;�y�<0:3ּ*Y�R�Z�[>��U��:�I�,�MP��|�3@�zt�)Axh�ӶM�ڬ�����w �<e[ݕ��Ό�ɚ�U�4��.�i~UT�~Zȡ^�j�v�q�X+V�GB�7[��\Pc���"� <6������-�V��}y�� ���GI0-܍���E�+Ȯ��x�m�z��}���G�`�w%���q��
�dnI��r����!l`�F��X=ܢt�wK���q0᫗=
�aԡ
<�%@��9VÍj�y������R��E��4�����>�t���ՁG"��+`ML��
G����A�|��R��=/�a�W�� x"ex��X'�>�*�*�R�h��o%ó���N����p�� �b�������MǤ�^J�s�̜�	:=�.�|i��i�r�߆���ld�ͬ�3Y�7��o8`EFEо[�f�wZ��=ټ�𷩷�j>�"6އ�i�f*����m5L_;]�=��{р=1|�g�?s�*
*�i�Y�A�l�5�Ɩ�-748�HQ����a���o�+�gDi|�r�hV�/��^��;�p*&���������X2�GS���Z�%x�q1���Pq,�NކM(
����ƬyM������<����Ҥ~:3�>��23;�8�g���8	���`N����C�����Ѵ��}�g"Qq�����B��<W5=�R�/�Ce������,�����1
@�k��B��z��;"�[h�������ƥx�P��a��ޕ��B��K���^D�$r�g��f�s�r��a��н'�:�az�����Rz�X�#e$�*{{��?Ui�7�AC�>������'tt��P/���;�v�R��5�����2x.
��z��%��ژ���K�(ٻ�A/�E��
8+�Q�qRt�/Vd8xTu3#��d	�1��,�gw����u�jo�!�K�p�2� J#$b��~6��|e�U��NwR�5�*����`R63J����Fϝu^�K�ԇ�֌Ɗ�Ec��5��4�K��<��w�z�X�E1�*[�mhV�Kd;DR�>/�g��#���>�$�H��#�A����	�%W(sM-X.�P1���Fa�V��}�D@F����[FBE�%.��m�yF,�j�T����{o�j\��j���گ;���޺��Ϛ%E�ɐ6�n��A47:�v�$������_�E`Vm3UoF��Z+�2��I����@�&=��;�^�`(
��b�b���EDq�d�V��eʏDtg�_W(s}}�
Ƅ>�2�
�Y��*��x�4�{���#���m�f�ҷj���w�%��#�f����|R�\�����D�H�yB�������ؑ�#5X����`�X�y�hR�U�a�q�8�콹��'����0F��ZY�X�v@����pV�.[�]|��fOH�F�עq�X9�����Z<3Q�8��LZ>~DtQ1 _�Ϝ�2�t4z-X9N�fC�`�^��#{��ER����^
�5	����F�S�W�c�w;��ޥ���W#�0%�k#�V�$���r7���{��u��VP_Y��4���X���p�>�} NL��a���vj���V(	Bǅ�X���z�׳,�^r���d�3β)��D�|�X�Qt>sԅ��X8�;ʎ����7%��#�]aʺI�k"bt��b]d� ݙؖT(;8T[Oz]:K�6��
�+���2%m(�Wj���\t!6Ӈ�_���V<�� 6~�Ǒ�ס����<D�_��2�Z}�L�c�S��A;8��ld==7!L;­��ǋV��I=,�
c����ѐ-�4���N�g4:��j.fʃ��rP��ʆJ�h�-���	-S�=��R��������h�N|+�yCr��.�����^i��t�u�	;�룽��P���K5r��:�i\��z|�	���ѨNgɋ���#m��E��o颻(O��ɪZv�*���C�w��� �X�a�8����F�*��>�=V� T7[�[�xv�ˊ��*j&:�P���*c�y�=k�����Q�r��誷-��J��*C��prɅ�o8��k����h���u%B`\9;����t�L<QW;�^1�2Ld9r'�áѹ��U\�Σ�$����|EA�O�;Qg���_8�!�X+�Ar��@��T*N*�|+G�m�z �!X+�W�V��ϯ�1�j�_qᢘ�<p|�`�[J�,nRח��<���T�'���;H�w/���;=ߦ.��Y<e��5Q���0����IT�Z��",d�j�ME��y�+���K��׍�u��~���c�1�9DG ���� Vo͘�OlQJv��hVWy�,��S��v��ܖ]�ୖ��T^~��M`,���Ȃ�Q���[G�� k��oI�w�C��x`�%y�Rg��P#A��!�D���ۼ���|�P`���W�}��4�k�m�{�����0",w�k�>�
MxA�8�xX�]r�����ݫ�M >84k8,P�0�Y���}�x��Yܗ݌w�xh��t�5�*Yт�(WŚ0,ꖚ]�!츭*Y艩��q.=q�}��\�EmV����C$-��@�]1�E@Z��F�qh��{t���v��n��?!�>��p��M��0�)�a��kx�L`,@X�k]���.��4�cyl�� ���N7���[��	�ukӉu-�P�;�g����,ޱy���9��e�	 V�-,G�n5Ƴq-]z^
k~F��'6�YP5�L< �ٳR{qna���n�](���Z��C+y}i0$7�Α��s����D�$�V��4�(�fE��k�:*۲ӻ�ϵ�ε���E
���ݍ����q�s:�e�`A�Gs������[mk��gm�Zn���rQs4<�1\(+) �����X�ٓHWJ�-IU�5�jԨgQ����)���k45�1-���a۾C6c�ċ��:����
�e�r��j_"��,TWk�VU�;���]�Zx
{�*3YQ�N�Dt̷K��u"x�F󓑅9�9�I�y�g��"�s�5*\�gN6+����M/���#z��
�(�<�7DP��@Wa���׺�MB�%��=�DPNUԵ��N�t�2+�%^�Z�a�`�)���1II�ϣ:���:���7y�̣ӵ�	���jBɭ�]);�tr�ݺU��ճy�nh�_�.k�X�8W�u3����SD���x��ԙ�x�� �y(u�ŗO�'�EG��|�Ź�����)��s�ذ�O�hj��}�O(e�G..۽�p�*�ܨ���R�"�x'oE}Y��r�Z�ZYR���j�9�����ι�]�O~o��� �Jr�30�r'$�+P-4-+��%	LIM&K�`�6aT�����d�K�H����SQ���f.H�ӖAE��YE	�V���hL���������2()+&�iɬ��$�"W"��*��0���30K2�Ȋ*+,�0�k$l�2J2S rFZ"0ʣ#�32�ɉ݁�2
�0Ȥ�(�������֦�Uڥ�K]�,�l(yM��"HA9X����#y_��R���]�5i�Æ�Z4:��Sve�y7;H$S�%���+�]D�Vx2����M��5^_޺�!QǢp�� �	�dt=����u�2H;uQ�Bp��-`�����+�u���m�ΥC��p���s�A���3��UKڇ����x��s;N|d��<!FH�0%�OB6q7���8�v'ئ�b��!K���ط&��yu׌f��!�a�3������*�3�q��G����������D��ae��5�y�<}\�xn��#��G�(���C��s�|MMVi���,���32�@�>$H���W]����hZ-^��,���-ꮍ�;,�kF��P�s�A��FV�Ub�����X�<qH�}�(�7
����":'#飰cfϖ�8�w,b�ևf�UbA�U:�i���l՞�=�
����*�磆���>0KB��'?�y��7������Y# K�
��b���S�ןV�o�=ba���~v+	VPVk�i��MV2���ӽ�׮�����#��<+�a���m��/9��L�K���*�Gg���R2����������7ͮȪ��o��p�%�E��y*��ʑ�Ӕh28�yӣG��t�065�]�v�WPǇ
�B<(�j^��Qp�p��DH�I��d�����5t}����7Fdû���6��k�|�*$�;|��jR�'
=�j�����F�Z�q��.$�U�[k�~�������������##�,�t�AW#kf��4n�������D�%K�q��UpTNA��%��;�j�4�={���&�I2ȃ둱>b]b��bރu�E<)�N������,Z
�¼�P��q�w�k�Ro�b�-(��W���(d,z��� =k�+*���g�f�f�MO;x)4����Y��bg��?f{�+�`�,h�������\h��Vl�9roow|Yd�WZ��شh���1v`A]���F��)��3��D�W���8�q�e�*C���
�q�鷝ݨ��R&6")��E�ԁP��3���Į��=�.IZj��E�0�Z؇6�qβc��)䰗Fhf�.��x��A��*����4��.�w\v�-���.QVWR�I,&�g%��ޭp>�F��B�����[.��ۗ
;6F�Q��Qqg)���d��"�I���`H.x8.�8�hؕ���Ȿ���S�0AV3�Z<+m��ɥ#��F�����Y��e�3�D�2 ������&-��w���C�p�ܑ���fc`r*�F�����ySI���SѬ�51dL<<8]�J��+FU�@}�Tٳ�{_T!jv(�C3Eň+��NATtu\�T��E�b�}���w�@߮�}5���e��0��A��)I��}�@Q�W�������F�-�~)�:r��p*�B
���(�=
&͒(p8��Π�r��nB�{S�d��xt�Z�q�^��ͪ�6���@91��p���nf�Yw(`(DС3v;<j:��bUfr_x	�M�O`o�#bQ��ǆ�[�(�q@yڑف�rtN�`��xm������U�;?#MD��&u����h�򡧂��4��
a\Gr=�ۧ-����ў}r��Hmʁ��5����ˎ������Mff�o��ϰ�
��T���
�)�و�ʎ����@�OAW�^�Yvw��tX�G����*� *Ϊ}�L����
�Ef�z��>W1��e �۳t�H;}2��u�`</Ċ�\&�`��xJe
�:3�����]���c��*�3cE��vH�Ʒ+�����:쌻��^�1!�%FXS�$��8
/D�,�Q%(��[�u��q����{c�Qݹ�[�2��\��yS.�c��ozH�ϑE�}�
Zz�<v����Ev��U{9'?U}��b��{�ဃ�+Й���b��D9t�d�k��,��X���X ���&^"�#b�
�,E���:��b!���}�^ 4!X4c�c�:<>u��n�7���Q�p�^�R�W��Æ� 2u�p�ɾ�ƚ	��V��6����K]8+��B]G��qw��>xW�Z�)�,u�V�bA�U�{M�'T
z���Q���a�*��=�@Ql*��T���&�c��K�aە�פj-MX��Pp�/���ךi���0�_�إ��,W��գ��x�ypA&����P�V)�=��e�UJ���X_%�ٵ[@�;)�1=�� =}�N߱���`W(��yO�����I\]n�{������tq�V�%_rK�{�ԧ����&c�L��d����LQ�p(�QҺ�poa����0q:�Dp�0��Z�K?%ʶ�:r���V�:�sc�"��\w4k�@�)ڥ^4�8<8p��~z­2>�b��64p�B돂&��ЩH�_J��V�z\t�V��C���FCcQt�xVX��ogf�(Pf�תҩ���
$���\tg�c!����V;����I�$���4T�0�K�5�|q��xn�u�^�B�{�P!�G2��v��@��P��E>�l49j�ա'6>,��_`�)��졎��x�>�@�틭k��s�ϐ��:�@ד�4T�V�3�K���`����46�&d��r4��	�=�QZ
�����w|2 �%��I�LX�k)���],£tGm������h�ؽ#�2㴱��� 02xQ�Xk�_��{�«a�y*U9h���a-�� �[���EiP�b.d{���dV�0G�Ea���K���uP����jR< ��6<��:T*
VsN��8J�5x���+��:��H`t��}����܋Æ�*V'�I�Of��̱%��P"p"j[�*:�3�k�=9���A��<W�B��V�_�Һ�C#�'��+�����\�MA�8�=$�=Ȅv=�@��Ocy=}�i��8*;
6�2@�*������9�Pc���D�c°e�!�4p�0%J��Z0h�*�������m�e<�A	���b9z����|ʴ����T:��p��;�1��O1s��ט���<��p�n��������F��8~u��ɣ�3���W������V�N���3����]L��ؘi�]c�>A� �[�c�s��eH�o5�7�;˩^��=㔹r*�\U�
�2�Ϋ��i�-�'�:9��W:1�J�Ov7�Ŗ�����y$18�;r{�W�ĩ�U�c��Y�wF�ٶ:�C�k��WKށP�6DxwK�iɥ�;5�;y��e���T=k�� o���w׉�_)��/ʄ�ǟƏ,��]�f	>�5�qc��+@�,����1)ZA[[�Ad�+{:�6����/'R΂�;��Z�j�nQ��^���t��<��{����e_J�{ox���޴"��<ĝ��1q�|Gl�dTS�����[m�7�-s����P�W��a��@��"eꖲ`�-ԛ����r�A�嘯3Y�C�#	"[���%����۽.�hL�r/��W�_6/G	���:8�m��J'zY�ك)�&%�ɪ���3�(j�.#�Wm�.�\�M�'yY���z-�u�:�ʝ�so��3]߿�b
��~���n��T�c�AwH��2�2ơ))�Ys�[Nu�nʓ�I�9����>K��@оx;=���*�o��hІZj$�V�۰�f������#��Z�Yg�'-�[�V"�|��>4)�3�@_�T@vq���D�CM��,��˧V�-�Y���wq���`
����s�
����M�~�^#���do)��[�qx�om���r��ݚ]dE���J7m.ز�n����ٺ��i��c��o�͸��5�vk� ]wW�*۫�M�7��,C��ݎ�B��MJ:��F��zk�U�P��j��hD);)qQ�͂ﵤ�l���������QMR�u�ئIn��q��)Y��B�R��D��Y�7�`';Y>xt32Gi]��,@��'�)ӄ81�L	�"XeK��Q�u\"�j����T��J����5�@�Y8d�D��NK�vx�xn��Zq�<�F5LM �F���j��ṿ�a��DL��S�:)B��b�zXVu�[:97��a�n�\*�R5tVY�U��)T�E(���5�\4,ޥ5�cUdu�4Hr*���1P:���(��޶�=Ć�}���NN6H���2���	���|r��S����o�9WU4P8�+k�o�͆^��u��!2T.b��Ψ��"�r]��  S�%gP��Hv����(՜ܹXn�����볻��O`8 ɳ"�2'' ȉ�$�i(��32�r�"�",�&�"�l�!�2�"�*��̨�3&̭fe��5e�TW���-e��5�e��̊�31���3�0��̎�Q���,�
�-�Z��&"���*#&+3("��̃̨�Ֆ���(������h� ��޵̳1�"����"
l̢ȱ�*�����³0��3#��)�ɋ Ȣ� �©�� '*�l�*F!�bjh�ѽ��������I���Y��y+��q�\�����
�DE������>��� �s����3T��=�h��F��t����~�s�ڞS����B��dC'�6��}��rqu��{�Gt�#�"�ޏ&��xK}��wU#ZKU�߹Ap�e�%� �O�zC�7��}���WD	���+��up��rb�M���(�K�ۦ�������턺sh���%�a�8	�cշ��;<<�uۼ�t(iވ�7:��>�j���"�<�j>�R�������&�8ǝK*��ļ�������Zec�)�.�3IㆳF��[QQ.�T5¹N���W�����wn�I+ݦ���һ J��쭬����v6��,�t[��B�tP�\�=5�k�k���Dc� ��óT�*�4�qs�Z�Y�d��#Yʥ�O?n�����==
�=���֛�g-�̕iO�kg��a�tɚ�FD0�A��wm�9�Y����f��f.6��x��ƌX�Պ|�Y��t|��񸔒�MC�P���Gc>�2�f��[�s�W>1�r!���&;�6̣���
\���U`޺Ǽ�3K�/� 5�=�s��=EA�2��{u:�Ҷ�ˠ���otAa�p��gV4,���v��8Ĝ�T�<+�~����4)�+��~ivm�;�g%����1z�w]W��yàN6������^oupo����>�b�#m��.�UVU7���͹���R��K	W����\J�r��k��U��=�J]!q���'���3�Xg���bVm�᝺��|����K������ц��twn�Ĺ=�GW�tc�*�7�q
�����so%�rs��s�@��x X���IŌ�:�������	��:z���wF%S���㋩H��Ofk��S-��T[�-�Ĕ�N}עy�^#��,���}�&���L^�iYG�WI�x����R^��#�����4�O��\� �t���T�����ۋ��1x&�[�ֿ_/�����p�!=~N�49M7�,֓뽞�=2�qP1�;��f��%�6��z�&�S�ms�{8��Ƥ�q�3�2�$�md��Ů�7��t�_N����K�������t�m�����!.T����jܗ��L�$D��V`V�A��"|=�v>�v�|��,^H�S�{b�J_lEfݩ�9"�(�ٻ]Ct�'k͍Eۋ:�{c�:
�Mw���Ȯ��%����3*�b��	�j��-�iP��77ەN]ѽ�Bˇ|�����s�H����}�פ2gv�����O(/=���f^����Z�f�8I>�r��Ӹ3"쬚|��Q�>g�ѹG�=y]4��y��o5̂�ט'͝�ҳ�R"rE���{ȯe-��J�����h��sf�3�y�1����#qоw��\O�I��o6�9j�>�ж�:Z}���+1�u2�-��s��,��%�w���{��Ěʜ�X�w34�^ʷ�c��p�e�a�?y��m�t�K���=b���/9�s�:3T#nF����փuV��&�o.2����]�F$�v'��T�~��M��U^e����و�,L�G�4mv�Dh뻻ת+��x�I����©����Jz�M^c������#i�F�S�v6�6�^��X!O9h�1-^L
�Mn�rǬf�fm};Z�g��C�ȩ&?I�o��Š+0S����	�����f�7�g�.�9��]�;mpaj&����%,����b�qc7�j�{��q��lQ�N�l/s��r��+�W'�S���q�NQ1����B�5���S�:��(c�q�B�:jﭪ�z��O<6��Ov��]rn\�����Uo8p�缽sP��I��-�����m7�F���Є��A�t���$�t�*a������QNF��z��f�F��ẇ�G( ��t��m]�	������U3�Yk㮅d����/�tC,��cw�+7�.j{L���t���$Ȋ��83}m�
z���ԯ5I�Tå�������qe�ɭ��Υc[����r�:(�{�E"[�Έ��7��J��O2�ɛP�$�/��w9;OX�0P!�ԻFoνK$�+[�JЫ"jd;�k��CO��c����.�m��:���+U{�i7��q�n���}MI���a��84M��\�!���[��>͵�:)zCX���/FO'6w�59�.��w롚�6�Y�����5���Zb&�/F��aߢ���~�v�y�0�����T{j�V���!zD��V"�k�`1��2H��y�Kj+���8�/��[�����t�N�r�T�����{��qQ��ni�fK�B�'�u����$-Υ�[.f��Ji�tyW�Ks�W��ތa{�Ngİ}��5�0�DK�H��+5=�7d4��VQ"�4�.ښ�S��mr��eJ�{������Dd)�S}٫UKr�h�ˆ)5k/owCq��$��w7'F�BF����n��X��N����
�SY��<���B��.|��.��u.���%���q��x������A�^t�TS��ZS�v���U�R/4����\ٽ�����ԣ�6�7����o�+s�����s�M���+��W�G)m9�-��g��,��L�ꍡ%Ȧ��,Wy�sF��ផ�Ĉ��:h�e]	��J;ϵ˅��e
ns\��V�fM��+��vE�����&�Ӽ���hXS~�.��?r�Pn������m�]�N�W�[�μ�w5�1��o=�~�g�`m�hH*�3�.�*sn�M�����7�m\ِ5�r�揈�i�49+g�K��3��miRʷ�T�l�F��k-�N�E�Ɩv�8Jsq�e问MS΄>9WZH1�ČO���t���&b=�]j�2�m>�3���oc������Uu!��!fq��妓]�U`�a9�ÿB��P �5�T�̭�5fa��d�;��a2�[Мo��֪H�M��n�ܫ�������k�n�e�6�M�:9���.�v��z�V�1n�1���+�]=í`͕|�@(��9-�P��e*����J�k��\=�ң���?�-p��IX�j]��q�e�Y��8��;���p��d��v��cr����=��K�$�pQ�S��t��;�M�gk�����Š31�luu�>Me���=�T�r�7�76�'ˮ�Jw���m;���m+�7AŒ��?9{A�Hm�ű���ZM-���[�\��t�5��d��sa�2�zL�y�/D�#*'���X"T�p乍����Z&�duX����)��]*�qH�Le��W��,�^��}\��cq���*�h&�
�LM�3g��|��>�u��[q�"K��]m7�`h؛���uv�_�*��7�M��Wr'[;4�[9�d��A�3���d���QAZq������E^��=���e1]N\�[�^2�����,vg2��:��\XaE�V+��h����V�@Db�w}�m��G�[3���>��N�3Wぬ����4�,�2.�Q�Z�i�o�sѮ�p��Sjc�2����rp��JrM�j�~����kʦz�[���w�9��wd�i� (
� �>��(��ĉ�����,������,#����f2�l�Ɍ����ȉH�Q���"��
���j\��*rL�#PaSUY.A4D�f�UVXUDUU%D��Y�1��"
i�'b���2ɳ0���%�)*h��(3�2�*�1
��X����L��F� �dZ��
,�ƈ�"h)*�$����
)��J����0ˋP�xaF��1�)�(*�FPo1�XeDIYFY%MSI�M5fdk0����4`f�ȣ޽ٮ�������V,+ѷtɇ���[�R�6�\]�'(�?��k�;b�7��C��B�b�i��}S���g��_�񙧒S1�9����K�V7EM6��g�57�-s��2w#ZJ?_�`jݎ��]f��򄞘�Kڶp�]Lx�/��-dJ}��n>���#;��f-���k�6���b���$��_����mK����J�~��V��;���m�������$�}�����Hc8��C��-84� "`�-��f}���������>���&KSm뻳����l�{��b~���ڵ큸�l-I�����g��d��@�]L���*�V���a���Q˖�hY�CV Xՙu�9�ц��p�V�����tD�ю����󓚕�Xu�k���e�:wv�5sw����u����ʲ}z�=�p����_�{�V�"�N� saē�^d`����&
�F7�U�D��&��T�ݠ��x�@s�P{��4����:�Ͻ`��WP��ˎչ�����O��޷OenG��&�h�R��)�)��.�
���0�v0��^�^6l�ͩ0���-�C^s'y;m橱�]H�s�Β(g�SF��o6+0�s��d���f�+;�;�{���b���_�l��Ӝ�����eh6ߤWb(>���:���8Gᜉ>ⵟ^M0���6�ܹ�h7�[��zj�P6.�|DeˀD�L�$�'�˻!�<�}��%C�'&�gs��z}Cj�GX�"Z�p�ͳ�n{gSҖ/b�yA�*�9ZWY�,�M�ml�	xQ�Z����<'έ/ywE�� �������۸��u���=��qR��S̉��-��c�{���I�/�E��3�a�М�-9y����on�WM�U{R�$��^�0�OJ�KB�G)D㐼�p�u��B�}'ol`�WOf��oe٠��;���'��}↕����l^L�C���}�n��dOM�H�7�+*�I��wy�M��P�T��R�O�,�Nnf��T��>mz1��ֺ���T�Nv2)6�D3��p�K^:ӏk;y��:�s.7rE^H��oF���b�^�r�`��8����۫�VeH�}p��c�QqGNӻ�����Y9�J�%�j��%
)'r�}����Ūɻ��l�`&��܊lҔk��S��~y^>Ud�@�=�)�r���W�|+�p��M�y
J��s�L�jv"�v�au��y=�3g��<�]:ܹ�k^����/\g��F%@�ˉ���8�6�u7�h��;�u/����7��V�^�t�l�b�jըI3垽��
�rv1���?N&���$�xۋ�P%�#�i�SZ'�_�n���$���w�a��3����@�doY���;��2��*6^���=G/���ת6f�m���J������!ޥW�e���QR����-*��)$�c�w=�/s"��O�N�I�7[�/;ݎ_���yb����td��h����5�z�Tv��|k1j>m��u��6>�=�
2���%e%��(AQ�_F�)�d���̒�.��n�Q�_Y��}5�2�m.Ʋ�����XPs=�%7Ɵ)�[���c/e�ޯF����%p�7�yy�������A���i
,T��}4��ûXd�ƌȤp��˹��U�\.QX8�4��Ot9�n>2�澸Ɉ\���Fji�Z�ueaIv�36�,�:�Hxd�HDݑ��"�sF�,�+�fU���$���o����ֺy}2�z�v>o�����rŊ�8�8��ɢ�-�
�n�>�E�(U���+N$O5���V��� f�7�SM��i�a������rs���f�T�rT�9���o-z��Q�r�{�6)�̹�S�o�ל��Ηˢi˨�k�64�o-˼c�nM�st�lgC{��7Ϝ�/v��|2�ŹS/d��ۮ2�v�q#��-��5]��ʝfMY����}-��t�N�{��\���\B��\��Е�F��.A28����i�z'���.�ic��c�byOރ��Q�'�ִ�bNjd�p=�A���k�ҦkEv��{��3�e��E�罒(�Z�N��	�R�ov������.u����U8�sw%-��읮ĭ�g�2���kX��G��R2L~{ ��y��T�V������t������g�]�B��jr�)K�>��c��f9����gO4y�K�nJhs�֞큚�|�jFm��X�`��+����PVnk���MdU��E\#�A@�"sʀ�I�����3iA��NޕG��1���y��oL7�����1�'��V���g<������w�c<	����;����|�P������Q�ݶ),�;�f���AԴ;0�C'7�\�8���/Z�8ms���8�m\h�Ѻ��E{w�12��+��	�Hɸ3|��ۃG���b_�9S�T�f�U�{ʊ�Ef]��0�:�}9�_q�Õ��P2���ߐ�%b���ǔZ���
�:�9��g�eP��zq֪Om'��)X�b��N�X':iv��Td8>������a�.(��ݍ����~�AS:�Ք��'KXk�1;m��9��{�W��nVbG�睴��چ^λ�ή#rrcj� $�RjZ��^QW��c�:!	齇[��t�/j٭��>���R�ӽ�{ṗf�շ#r+�s�ѵ4�ʠ���K��72K�:�m���3���-�mY�o����������'��RZ���������1k�5}[N����՗��2�7"�ກ�T:a���^�i����vfU�<]SH�J�*�n'S͕`˚>�(��:��ϭEVZ�J�k��K
����+̑�fh	w\��YE��I���C�6�q�8 �[�u�Qn�0mI����j��.���
;����%��:�3��j��6��Ǒ�n*���\�#�j�CCz�D�/o��l�&ʻIT��o_q�܏n��a���c0;�)T�K������-����ن�k�[/*�Wc����η�P�lKzwo,�Li�S��
X1į�[��O��}�H�2�Q�*�݁H��� c��[�O�ݥ�SI�1�L݌|x�@�����,�%�8��0Y5p`O�W��b�v#���D�&]�T�ǻ3���zڻ讗
j?�6���^&͆ �Ƽ�F���ǻ�����A׼���I�y���JR�o�au��z�|4ڭ�u��)9�^�l�Osiϰj������:��[i
����]z2E҂�Z�ͥoV� x�'%1�t��yC[̺w��޴�v�"��n��Ւp�k�teh%$��d�Ŕھ�ܨD�5��-<=qAV�eK�*<��r����JU��YZ�2��@CB`x���ųk� �X9�{�X]�;d��V4nBpt��{�L��|���{��}�GQ<]��H�Jg��33L:7��u��ئ��n��f�z��5�7�u^�*��/� �}�NQݑVVf^o+dP�Pw&q�fa�ta�Q�̌��
r�jR�r2J�����kM��k��(�ffkĠ����8�ތ

��F�����E4Pn+-d1�'Pe9�DQ��Q�̚232��'Z�:���Q��֍h3Xa��fdf�(�*�,-fpiw�浢# ՚ƌ�]Z�DZֵRRS�jƻ�%��ϦP�{��B�U�j��*�{�u�D�h&�p�(��X){ʍֈ��Q�,������ӡdlRH;��X]3+��uic[I�*�`�kF�f�)7�c+�'icH�.�<�,L�]����Cw]�K��o"f�>����\B�ю�D�0�[�w.`�q�eu��]˜�֝�V��(��,V�Zw[D�ͮa��v���#���o���O]ڳf	����{�&��;���UhJɝ����,%S�!\�<���By�$r˂�\6��x�!�V�TaJ�.���6y�����0�:�As�Q{y�J
�n,�Iͽ�r�n����J93d��:�zۼ�*(����U׷1�s!�H~j��1p;�NO,]�tnjs�ƮF���"�GD��G^�ȷ˛�F����`��e�2�b7���ʬ�	�u<�'��s�=�d��pxYӞ[Sd=(_r�ޠm{���,��*O7���햻�Ss����h*[��e���f�콭z��ڮh,��\A��r-�����o-j���7�G��ٽ%4�x�L��B}���콋��QԾ�0R�H��~,T�w�^2˷�{��X�{%ޅ������W�ȭ�{�ջ�)asS-�pehk�n��[&ŷ��!
7����yk���q��wz�gf�+#'ψ�R�gL���[=M�s��vr�]����6�W�fPw/{9bnvϖX�0x��.��\�M�\��}�{k�o����R������"�n�\=��+v�y�G����v��l�+��>����;(Y�Wz��{S��(f�����>-{h���I���'��ۑt2-�R�1S������Y}�.[�:�P�ޕ��&�r�c6���@�v'
��]Im��*}�T�ݦ��6U�����mQ'�ڲ#��3*{G��J�����Xf#p�f{��cd��.���5}�&�1Yug�خ�[�~6%=�&g��	�zFq�E���ʺ}��}��G�2-�l�cǩdHg5��e̵�!���Q���_��~O#u�Jx���Uc0a���1�z���p�e㰩ݍ�D��������f�ΫN�2ŧ�������ֽ��#��攞%��������1�X�+l�lG7۸	��g�=t�=w�N�׭w5J�b+�9�;9B���}*��r�*�$�2�H���2;rk���K������Z}g_�[/�ENW��'�){���u�V���y�v,;���[�P�=�ٙч.S2+oT�w5�c�DO�-��O,U7��L�N���_�玢t���h����
�:��!�}\B�piw�%�ܻP���b����P{g��12�� ��^~t��2����5��8�P�d�k�b��>��ݬ�ⳗ崣�bU�J�Z��b�*��D󭥏9JOݍe�z	����p�Ɏ�]f��-v�{0ٮz�qr�E7��T�^��V��u䮥�������=tyk:�U���<�?7���xWV�E�3���Ǥ;��9JV~9C�֯''f����e���n�"�cH�^��pgp{7=�g���3�n�ex7��_r)�=�Z]���0�<^շH�~^������z����+��/�c�����*H|�نZ[�8j�wl]�׻���0�͚�}gGVou��FQ�)�ea��9Qf(
Vy��w]��32��!�r v�[�4���:i��L�.�[�e����2+U"��T�f�-��y��FeKs�E�ovj��]��9���0f\�UL�r��_b}��O��	�]�\׷b�9;s�:3�q�a��foa�X�'���jv3|*F��ꉮ�3q�á����YB�;�Ƿ9�8���`i�ę���{�OM#����]&t��Q���=�����2��p4o��y�ߖ�ӵzA���*�rll~�pM�0v�'G�*���0��j�vCׇY�S)�5�{���Ja�������v�Q���ʑ����Zv�:ﳢro>��yQ�����mʭ���:Қ�m�҄Z�Q1���>�	ߴ���H�j��\���N���)��.�(>Kh9m��E��G���;X��~d��[��ش�?@=��*��k,��Ko�cK�	������{���GoL�|�ƗTM���s��(��5�7��JY���-~��Ѧ�c��3ž�c��/�<s�̖to��pS0�ϥ�d�8������Qb^��M!�Û��1ۃ+FU�0�>������4��#{�`
H+��
gQά�f93�<��R4{�ऱ{�3�Eo���\��9�����=�^*O��U�5���kk��`3�W�-Vpf��ǵ��H�;�^cW]N�'&��2����]�f�����+���ϒ��oL����8�
��]%Z�α�J��ctY��]�ջ4����ŧ��%ݝ��!��z��꾞yI��|��{������ėT���>�&*�}>ǭn��-�(�/)��w��H̩|����{�¨�7r�׳q���F��������E�X����.�=�[P��㱽r��Q���c&�5�W�NP��F'0?Wk��	)�"�ГոҬ�}��FL"������s�m^UGTƫY�k	3�.���ϯ�����fl��Y�/OOk�������+�̭��g��Yt��D�_{��DT5]��P�9j�e��^�7��
o	�3M_����owd������]�C�9v�o�����#|�u��?��G��߸��0� ����1 PV�a��� PW���L ~��'���i���`kGZu�rmM����6���c���E TP-b�(*�,�ָ&�:9������s��?��3��?�x��;�������q?���P �����u�9��~�?��	��h=���ɄF�W���[ ����[0;6'A������CN�4v`���gK��&h�}�pqӰ��AA_�E����oGL��}D��8t�$$���BI��dETY%�ѳ�����a����dy],|1���[_�\m4��*���P ��a�
���!����4���8?k����@���ߘz����ÃP��{L��k�`���惘�QFz���i�yK�ҷ�?%� V;?.}a��f�#W����A]��_�c�_�C�G�aԅ���pya�fFKƞT��1vBI�K�^�UU%�r�xȝ7�s.�Ngk�E�e��^��'"\s���T��S)�\#�s�v>���~}��}����;���$$�oK$��l5�di^܏��CW���ŏe5�b��$Xg#ӹgf�����Ure%����X�In2N��w{�gs7�BI�U%������9�����q�j#�@�=�p�����)�� V�  �����Q��H�#���?�cX&��7$�%�9�aĦ��F���� *
���� ��@Ӣ��X?���ė���S�?Pr����{��	9�Y�!t#�(�i^yq�t!�9�x�;tU|��{W���h��nv�k�#d�pHI+1\]I>E$�e7ꃢRy=ا�ţ&(�M\}���8u��ŚįE(�Y:I��n�8TxG�%���#7��1�f���BI��2���d�΋,X�o�EvBId�����C�r����5#�����۟B3��:@�$����1���p?��H;�����Ƌ��4(�{������3�#A�%i��i�Kv�F�]|]�-ٱ*�����N��~����������Ʉ��_���;8h�<
~��O�*I�[8�Gv�rQ#����S���(���t���)/L�%���b^]t����>����*~)LAG�Ď�Q9r���.�p� �X�