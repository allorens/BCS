BZh91AY&SY�%d ��߀`q���"� ?���bA�}T /�
 ��P � �  4   �� �4�@ �(   �
� (   ���]�E�ٙ��j�-��6�j�I�mMkl12i������[2P�X���T[6��,m��2k-�L���VQ�l�L��R�6q��l�ٳ6�m��YZѶ٨���4������ԡ6�[a�kZ�[[Kf��F$ʩ����&ŖaT�E
�k$H�EV����:w6�J)+X�   `���֫7�Ī�;�:HUUSN�� �n��n�B;���T[::��؊s��B��w1��U�T�]���l�QIi��)� �)�   ]χAm�
�:�hKl�����-���(;�k��ً.g�� .��(R���t�F@��硠�JN=Mej�V�I��Vm2[mm_   �xiT��v�]�P�����ƺ��(h�=8�ր�iCl)s��R��k��A����JQ�;�( �V�B�@�rkJ�*Ĳ�Z���#�   l��J�������E�.-�(&��F��Ҩ��GAE(;��T�ܮ�)w#p P�.��1EkCk6ֶC�  ۯ �*�0�HP\8�@hR변} ='��4(
yGp�"JN�\�
K�պ�Π)B�ݭ�5K���7�� I]�d�S3TbҨ"�  ���(
����T�h�[nP����@js���T��{n4��R�N���L�]� &i@
�� h4h'��(mf5Zj�UKO�  ���*�/rۚ
U�֗N�P���wT�(e��RUn�  t��W*R�FuX r��:��p(���gt Εlj��[a��m����X��   7^  =ݭp (�v� �j�
�P:R� �����T�c���i��gP:K�U]H֊`P-h�j�)��  u� �4 �b�j�:�(��pP
6��  n��@�� P�p 2]� �ٙ��k6fՐE)kTO  ;�h5M�0 ��s� ���[�� ��� A�� 7=�u�0�� �.�( ��  � ��M���� �  ��1JJUi� FFC	����bJR�i� �0 4��T��R�      E	���қ $ڛMLF�=C4�f��)%Ji���h �  ���ў��<��O|�o���8ֳ��m�޳l�Y�sճMj�_�f�\��F���1TW^@�m��m��6���cm���q�6½B���=��C�?_���>a����(��o�_���6��;�ߙ�+�Q[����0B�s!*@��!Q����8� ��A �8��������!�~6���v ��?`��c�v���1� ��p`��?��c�p`�l����� `��? �`��lc�M�~���C~�����������7�m��dpm�~��߂����������!�6?`7���l ~ñ�?���� ���߃�����C�;~	�߂ ���v6�������P� �D��|P����o��*����H*᱙��^b��6T�[��O7�˻]}%*��P���)st'���L�8櫽�tװ��@�5�.)%�z�5^A�軗v�d�V���݆��)W7�4��Ro��X�2�g8�	�/�j��Qe�0	nc��G�r�����y���s"�1�7��Uf�|�6�x+�݄�<����-��&f��S_h|��ܝ���>4��Uڵ`O�T�����e<G.ZV�x�sP䢃5�i5���pO��X�$w�w��l��;��Q��ѭ��%WWP���2�)�> 1w9$����Y�0��i\�SC�RO3N��Φ��/�\������'��#��0a2�6�����i����:�
(�% ���A�G'�1o��S��U����.����h������Ӷ\�p�C�,�웝:�{ Z�6��ׁST��Y"��"2�z��r�Uf�Ū��(c=��f齎Ȧ4�������On��<J�B��G^�$n<R��&.��S�w1Hq>ţd�7N).m'WK1h'd<:g�r��|��x��8AH}� r{-�a����a�p��ױ�B]�G59U��������`Ԏ*Xd�#dW��]M!�_���,ˬ�5R��;����CP�6:��6~�"J�s7PF.��B.+��#�IN�U{n�;�+�i=t�'(�1}@�n�pw��	�q�r>�ria���D����h�Yn����N�W
h�u�*�n�ۣ���˦ұt��vn���mN�Wi�qԉ����v��	�.��`���q�>w���a�5il3�H٭��R,۔�9�<�9N��(�^�u>�)-Xם���b3�tM�ü���wv�1k
pK�U��nƆ���*9-z�IO�� q}��H�eI�i�b���ĩ�s���k�8��#�6�s�z�5�d>o���]׵%�ye�C*�F��N�6��8�9N>ih��wuJ��e�&�{
�FB�oe#-U�d�;�g��_�	�tr3�Ƃ���mIwt�|��jq�0��,P;xi��k��˦�o��'b�.jp��/$�Wk�ڌ}
���F�[f� W�oʽ�8<�A�\6	���>f!F�ẋ��Z��61v���l���F�ͼ�,r�dk:ƴϔ.t�]&2��3aH�ÂlLV�\��.Y�YOY0��
;���c�sTT][���fH�j�gmt�gF�%,܃Z��=�sZX���w��2LK]�S�B�渷�M/�Ĭקh��j�/lٚ*|��Ш���]p7D|!��p;R�˜=�̘��C���Wfq�:q*��!��
�ܽ 7�K��Ϲ�˿�M1&N1LF��&����{����WE<��A�9m�t�㩃4S�q0���$��d&NZL� Di�h�s#zEF��n�ݎ3]�pXwm2r��Ol!H����ϣ����B��P��$ �iΥ[�B����2��ώ攵$�od�V�lfv��ܑ�MZlG����#6w!��r�YyIE����q��[\Ç8���Úե�)F?Fv���9�cf:��%}���>�A(#�\@�yVKi2�ŭB�jmqY�9�:�]������<�[��l]ٹ�����:KӴۥ>��X����s~��{(`�=�s�q��B�4�c�p%Q�[_[9G�Tn
�o�V̽8�qhӽ�[�9b,m;&5��t�cU2&H���T6�-]\�%�!�%ۃJ9��|�a� ��u���G,,��v��>�����vqr�n���,�b��0�z�A���\���c�[�(���<�lj��|1��sF��=fl�79Q��W�7X|�87
�of�ޛ�������HS��Ս��"Y7�[W"����V�@��	��G���0�2p�S�{�EXޱ��+a`k�?	��ML8tf� �R��tC���MOov83�d�G�qH+y8k���w~�ojEU����q�:Q7&ʩ�N�;���gwn��`��%���/{(�. m���|r�s�R�WW9�\��Չ�U�'�KQ���n�]�v��ڻ'kG^O��B��θ�J7X�k��$L f�E��KFn��X<�k0���0�zr2v�#��)�2#mX�}�O�s�T�mq��cB���C�9fޤ���m�-�Z�@:Q�����T���<�sѲ�FRӖ�1�[�C�&��|u+W�<�i/��GfZ2�-)k���(��KN��n��U�̚7w�7IbK�(s4ŋ�M˧�B���F+���L�t�]x���9�)���C�٨�3�Z�d�҄�d0݁�	�8U���}mf�+�x,d��$�2<�ˍ�"�/QGu�.�lu���ǹq�\M%�o�5���%�`ه��ۂ���[�"����(VL=�ʰ��Xp���s�󡺞3��څVNm�*ejݼبف���|�����Sy#�_Evv��kDs��Xr<���ݤT�f*A��g-��1�\��\��3q`���{ 9~m��{�w�N�g_�g#�7�-N^9tnwd�J�<�:9�7��_��wZ�7���5R�^��Z����Y����7t��-4�k�^k�p�!��^��;�̩$M�E�5`̸���S��'���Ւg�=xl<2I;rƓ[&�wy���I�f�s�
�+�#�k���-=�ݒ���e�n˒
^n'��7CGb�S�0���1r�2q�Yrm�s��'r�^�^���޷@�L���<K=�n��g,��&�<�N�TN�������L���U�����Ɍ��\���-�Fq�`���lo�.|R
�c=B���DxI��E:�2i���Ի����Cwu��AtT��K�#{H�E��4���Zz��4�����\��[Q��^p�FA�mQS�JM��>k��S��Ӑ�������>����Ћ��`6�\zD7��Ql�a|�[�,�&�pƫF�1�8N�����Ty״�ﻪKp�I�է�>.QB{�=4����E���8ܴ���%�e2������-ߪ��ƀ2���ܶz0��
Ǡ���M�Y�q��V���p����d�����z5Y�%�&�ц�KĹ�/U�P���1
��K�^2ְ��	��פ��\�؉x�����p��}*�w\PR��i��ӑ�r�q[��)�y&K�Å�o:���73��V�2=�#�+W�K5�*�`��ٖ�osx8��: �#PjWt��紾yϬ�=�����`W�U��c�~臫�d��k<8�Ǐ����	!�sel�w_1��wr�햓���R@p�����3��qN"f�,��!n�Ą�6��a�enV��b�-+~�lcw�]��=_otO�=���6��Z��o` � �3��%�{�LɎU-e擰d��Ve��pj�+3N�G �����f9g';���7��[��+9DJ��X�h
s�ovv-��G8�i�aG�oڌ<��C�ڜ�׈r��uZ)Q�1D�HT�ݻ��1� %�;%�}�n	��m�Jz"ݧ��l+�-��GN���0�Q�@Sm�%��y�٫��F:<��އ��U�Fm$�8��eJ,��Um���uol=����c]*�q���h�4��kA�ު�m�t��ƈX����߁�$�mzا$b2����w0A�{t�g=#w7�vm
o\eω7N���!�5�j��>��aK.hipݍ͇�筕ɵM��$2�*2��D<��G")3U�u�U��[}��n�n�u��e3RVS�z 3\�j���xp�HΜ�f�wy���HƸq�_�J�Q���j���`��nL�t�ݜh�:8ag�2X;&ܩ����Κ�ygi�0^g;!�h�xnJ¹�qL݅�X3K��"֟���KXf��7�_K���#F�����\yu���Ks���TB��5�1ǁe��Ҟ�Lf=VK񡐕X���&���  ��]�om��ܺ�rq�jv(oe[nr�g�\J=&�}{�r���M72�#4����em0r�9���v�-5�\�iӝt�s�����F!��l�p��z+�:��;�b���B�B)��w-�D�˗�T�f�I�L�Z�F!SS,�$;*�Wtu�U�n��u�U���S75��^
��ܽ�$�VM�ll'���eԤL��D�7�/���
��󀳇�dĦ�3O�%��$�Ϫk��v�k�%��;J�lv��V߲w�n����=�{6�
�c�@��"xt2��2Sp=v!��W2ޠ��jK6]#y.\{J[&��9Rj��^����D���-=�8�W*VR���/[9f�\rҏG��6�%÷]2^�m����b����\h�H�Q�F��v��Pڊ���Xt� r���Ta�z���3B�&LZo*�c�N�H��!����wn�y&���zq�q6r>[��ɗ)�	�����A���nd�ۢ3��ǝ�_[���Q��jb��V�}�m�1VՖ��>��M��ǲ�#��z�q�s��I�\S{!��T�:{F��]-+e3R�L���}��vN�"�h��8�9��
Aw�u��s6<{vb��X,���3���$���Ú1n�,F�x�����D��9�������Ea����/]mΊv�ɂ���L�CO�&�n��f�Ś���Zw���t�Glð�E�$wiY��!T�h������H��l{���l�L5 ��'����D�ƽ(��$��"-��z�7�Fk���{HE��6��U�ez"ʞ��R�\��:�|�۸th��'�n�FzN��8�t�8�k]��-�qgy���g��u��m�` k���N[M�H��y����C�g��>����b["�ql��@i}�;�Ȑ�{L�~��K��&��ܘ�8~�_Mm�fsL�z7��h��ݷ�ݹ��ib��q��ׯ�AA&^���U	�ё���v]���8��μ�GtD�[(f�|��Gk�&����0w��>���3� zs=q,��Q��������R����V��j�GD^Uq��k���1K�1!'L|����nޘ֍b�d�U����0�u������G`u��ԉx\.�%�qX���WJX����4�e��H��H)�#\�Ǚ{
���E䙭l�G�Ov�:>t���K'�䡄�hO�{^,ghG�ݺ�d%y� m��`L���1wr��mbl�<2;����o��=p���!��zv:��7�,�A�X��vcj�A38f�@nj�9�wؾ��K�X�4;4��@R�{����A�7UY�U�۵>���?JW����/F�#;S��Q��6N+,�
���
=��q�;�
�T�\�Bv�z���*���zD�TYE�i��RM3�n�o�Zuh��.��u;VϚS"Gj
:���t �K�hg�"���$^�=}>bb�F���*�,�$�{2���[�Ѷu��M�h��a��i�;7����I�1�UE��@��ܷz����+y�lЁ�UJ�J9ūs���L�n���Cs,���}�"�4M]��E;y�"Cŷq��{W¥�{������UK\�X�oIY.�e[�XhŸ
6$հRq]�R�ҁ�+������I�x-�:��<�4�)��hn�Y^X���ΐÂoom�m��t��OtK�A[�:z��Yӻq�iprkh���n��6�݉G+l�T�A���2�P���^�G�����vn>�p�r�]K8gf�������4x׻Z�<���D�IaVLc;Q6�Uô��Z���W��}��N��}�)�aU8�'�zN��DǴ�aP�h.�0Sp����*巅f�"��ʺA5�܊v�ba�3�M��2�a˚-�v���`�l��\��e9�dbސX%;�Ƶ�qt�v�c(�ᝫ���j��^�����*c����v�/;r���@
���8��RÖ}%��X�cޙ�v��l�f�Xu5*�9\z�sY�r4�s^����;{v��q��E��=��Ǒ�	���ƻ�3)/���_(��!��M��%������v*6��w�7wJ�}��3.j�R���P��F�ԁ��>�	�R�N+nNݰY��˻�P�`;ðm�G	�����1�ZI�3�KȵRD�+�%�	����/��%SeD{ݹ�=���^9�v.�/'1{�g�!`G��l�R�a�.��h�r�Vv/~�c���#��u��n^{5dyy>̓�I��*wVХ�˟<�$(D�dI��<JmիCi�s���#���{[�3x�i�;�i���!9�6�9��.���w����ft��'�]P��I�.��;"���ra��0���w!��T�n�i�%�m�Ճw`Z����Q�j�5��Zu�s�
�޺j����]1���)��km���4�9z����3A��2�2
Zkd�57\�TTaw@s[��pK��_3KEd�ɐ$PGV{$v=|����fk�8��	� /��*u���7����0kF�ɑŇGJ�9� �mt��6TGv+�$�hz�w��+SM9oЎl�R�ܛB�Ͱn0ރ"@����j��Ɛn��p_o���0�b�7%Ҡ�%^�Ϙ���f�LS_��z�8sx�����pRp�m��b��lsw�bst�ע��I���ϗ>Y�%���I϶p�tc�n]�:RW"9��N�9G����2��c���(����8]ٵ��'��a�Ь&�{��m���~vQ+���C8C']�`�l�tp8����+ө����X�ǳ�ҶT�u����CS�����}g%��(%���\Y,r��6��Վ���t|�ԝ}�I',��c�H�-��p�+Ѕ���_q������%q�qA�?~������ζ�ɝ�٭�޺��r��I6lED�2�.��ݣ�ɼ�j�;h��z��V��ػ��&š�}^�܏J�eF�GK�hl�[���:@���X��e�{;flT%�*�բ�+#R�<,V��U{n���[f�n�q��u�=�>S1MCtd�h4��ܫr^���̃�I]��ٸ4��Ef���b��l{:�C�uՍ�W��`w��$Q�v���*�;��U�8�շ��w&<p�;��q�ոu���F�ȭ�7$~{�7"�N�x���u�\�ۙ�m�]�X��)�S2jY�;��0^�/j� J��o���)�}r� aג�N��i��^���J껶�)*.9�:;�Jfm�}�c�����J��r�PwC�Ej��ތK��n�m�X,���Hr0�H\D^��?B��$��KW�*X�{�Cw�Q̹��Bv�����Q~����*����׏�l��zp���i=�w�k���b�cGRa�+��`L{K#�-���}��xR8��ЅD�էx����(6���$��l�ORKe^
�j�DY]�ӡiK<�����#�ȣ�OWe�e�m��{��m�(g��v��2�ю< ��Qf�i��8(_V-.�b�Z����J�\�ӹ�2D��w�a�ܩ����PN\�qx��Z���NZ����n�M�-��_�l�-��5�.��k��Z��1s��98r�F�&<}XnL6k�Mf��K5)&��,;؍9Էd���%���j��e�4c=ܻ�5��{�^���( �n�V��h����,���!��w}:�RA�]�7�e���E���y�_7�ײ��J��W��h��XF����Y�G�9�3]m�fYS����|�ٞN��3Z9wh���r���:Do6��l�����p�(�N��n9��m�R��^S��'�lޛ��b����S̱�����wl�0�vA�cꎬ���ӭ�i�Et7���fӧsE�I/ʷ)���^�{Ƿܙ�]P\R���B4*l7n����fc�e_,��2;%_L�:O:�v��o�y�GX@���{y�ڋ�C6lV���[{h���[�]�T.���J�h������3�� ����c���ٽޤ�Zs�[+:�����i�"����林0��ȉ�����M������*'��f��5WQ�*+n��F��{��@tpU�tP���m�7�W
��:�{��=Mh
d��~�ז&�X\cQ,�{���E_75� �ؠN̉��nl��U����{�[��M�Lf�����/K��]u����V���:Vh��r��jp֭�y�N�>�5��]4 �k��{�ҤB�Yk����"u8���pP7�u��y��J�qZO���/��h�F�`�,�}��{�_B�=��R,��l9�����l���G�cW"�R��6u��s(R{�&X�p��M�-�ؾ ��TuR
Ǹ�[��f��t9�zL��v��w@��Tr�L����FP���HrT�/�^���5k���JM~=3�L�g_�,�\����q_HF�qmmf�WV�QbW�Zv��C:ի�9\����ܣQ���K��t� ���)l�H����*�>���N�n�gHe V��9��wp�J�z.X��o���k�g�>O�[#@l�Ľ 3x�� ���{2K���1*s]}1��ӧN�Oq-7(:k]b�V�[T�V�@\��K�{t����v�>�tu��K��
O{M �O��r�fV(�������p��%�_ݶ���(��r��j�(1�*,�-W�)�:7ܮ��:��l�]��ϖ&u5Y�M������fڕn��ǽ�v��2s����[}{w������X�'�s8�ᆵ=�:)��iͼ��)w.���G���F��b�D�9K|����]��"��ҜL't��.=��jӂ��u�WQ���v�j�c6X���ٰA�<�Uuhі�#��s~�f5�1�5�e�xY��v��̜"�/Г�^���O���Aw��B@�,4j���T>�_hF���Ctvu=���pmX���e͒dO/Y���Hwc��s��܃S���Y��`w0��qϲ8X�J�*I��ћ��SGQW�7J׀��!d��!N/�r�}��i}�Gv��>W��kQ|�������6�gn��C��f����l��h����*JC�t����s���G���4�;�0�vG��]�oUh2aYsl�齎����C
���r�9�"���t�ң[b�-e�쌼�Բ5s��W�� �1��f����^�ˈ�A^y!�{]�"R{v���Li��-�K��o�7Z�Ty�Ä�\�^s�Q�>�z�FH�u8h'Kn��S���D�4�{8Q�9��A�2*ڎ�bue��r�޽�����Tȯ3Zp�XF��s�w��A�jN ����ZFf�䀽b�u�v΅8��.�0gl'p4K�v�p�b��.R��.�g��Ǳ��]�����Pf�ͤ��\�k����S�մ��(�6N����<D�)]����`��l����kN�35��'9]^VR��-�9N�ڄ�1�`��GAv֧#|ni��+�����R&h�p�m�x��VZ�B��z�h�=�\���%6�B �;��E^);L������~�?C�"������C�TYw]�Q%�Y���F�H�<&���-�@��)��~���G��K�7��>�÷l���l�X��I��e�Bf8��)W�2b�gL��*�����	������ABh���qd;:��>F�O�[��{�:0)������uR��.�v�dz=�{u�gc�z��B#Xج����ג���wG:�!iK�����5ڇ�TP3L.���-s4{�{~���W�^M{�e;77�����x8��뫋6��y}��7!t�h"N��9C'�L�W�l�S��7��T�rt�㞘����a>He���,nz���ʠ����VZ�.��"mPc0,5��t�w�s8coZ���������έ8[�X���zuܘY����r�M��W<��*�kov�S�NP�Y��f�wv6�F�{q=�b����q�*��s~�g���'3��]���o�f�*?*bO!{��ܳ�՗5���%�Zӹ��fu��5��Fd�;B���;>Z����6#��j��7~�]��ą2u̓r�w܅C��\>h�@�<�<�f�n��s�9�+��yk�>�OwQ��O%�!��6�r|�5�/m��r�s,r�L�A��(��uȮ��ޭ�M��D�b��rt]�J����|%#Y/q�*��;W��]t�L�Ƥח�#�&Q[Jû⤜���hvh��Qp�?�B�i}��s�3�f��߻���{���˓4A��)��陘��!j��CY�:%��g&=�e3f���s�����}aC�
[�	uQ�o+�/DX�ԟ	�u��^m�� p��ȥaŽV������d�+ ["��[��9Y�Z���m��>d�և�d��*B��v���1U�-g22�_iW��U�/d	Yk�ݨ�L�����5r�7����`�;7��u�_K��ܠM����'p������c�\Q��ޗvI�;�kaWc��k\3�Ges'��t���n��cJ����6�!�ܴ7���ũ�ո�$w1�,d�Nt�z���d�+ʍ���S�w)���=)�xz��w}ޅox�֌���
�h��/?r�5��}g�V��Ks�x8��ם�Q���8��%��٢�����9vT�� �XR�15"�U��s�.�s�ޥ�tx̞*��w���5�^՞�k�tey{��tx1jW��n�͑�Ϫ�nC���RY�oȪ]W	��3Wd\U����Z���Ҭ�ഔ�b�t��7Fj�9'����ݔ{i&�Xۨˤ�+�)̺��"E��n�闭�P>Z�,�Le�Z�W�-]�s��P����ᯍ���tN;����yy��;����<�i �Ȗ��K�zF/S�3���i�0d�����E�6�����<}m�����+Fg)�5-� ݂�m���qK"v,3rV^Kw�v�ԭm[I#�X�̵-]�Xi=�"̐l�q��-DD,T��(�ɷq}v�(�[x�uY�,�ɓ�Q3d����:G3��|�[u5?�-и��=��<�~=��ͦ��	y�Ydi���2����)�<�A�Y��_(xyU�:��\�NK\4*�/E�(2Ȝ�,eGB���h�㽹+]��8��^LѯY�V��b�(���>��nk�~��� �$gӵ^7xl��	��9����7���\}�7�5_kj��K"���{F��8�8�3璯c�!����+'�4.a�I���c��A�LGҁ�J*�)C{N��pw�(��åY$��L���hX�u�vP���<���B�f���(yvY�;�h�;�ɛ�lˋq�9�w:[�,�ӱ�Y��c�ֆ�r�����#���Z�H�p�U���gb����v����rV��A��0�C�v����������ek�j.��v1NA��`)u�0��Z��.^��׉R7;T��KaQ͝�+�(9Zo���G�d͛�IQ�Lw�]!4�7{ޤ��&�9�Cq���H����6{N���+N7É\e����3�E�$s�o18d�=�0��+\w[��tt��h���x��	���+�#|�Y'm�(�ug�b��t���<Y��{��R/.���:�T���	�7
=;��3'QۉLz;��{�j+�I�7��[c��L !��[��s�b,<�-��<E��Ύ|��g����T> 3�x��%�&��HE��ڛ��]�2��.t����`Y~�{��-�m\Ҡ�든ƽ�S5|nx�AJ�c���u�p_�r�-eb���)��z(���$sY�;#�����S���#�D�;/s88���}vx<rw���*g��Cޗ���*���¡���ir٘��r���
�W1���h��~T'���} !�%����gsf�\̳��gw�k�k�۔�J�&~�����/�[�����3�Fױv���gy�/u����&Jz����m��;���Ƅ�rlCr�.�͋xh�J��/a��Ri	.<X�8��W<͑Y�X3'K�A�G�S}	Q=K�?�/�����۾��M�v��A�
���>�c�t��y�s��f�I�E��� ]O��Z|��P|ŉ�/g�e����T.w3�j���h0C�O��\+U��p�w��;��cp6�7n�&�#���G�z�d��o0��{�d��{7�3��h����$���hb�%|���D6kdC��R��+ev�jΏn���n1�:����3����K{�!�%�½���,��d<�p����8t��B����Џ �u'��	Bl���tm�������y?W�XSh~S������.H�i�rسn���~�B�F��0m���+J5,������.�V�Lܽ��j��ڳ���X��sאJcT� ņ�v����6�G�uc�}�8�Y�;�
�v���Hk�*eV]��8g��'�B+v�t�f�y	H�s[�B:���/")Wn��d���h�FԨIBuѹ���;����<��p�o�^�ن���n�=7v�o����j�F:�����nR��oE�Ni�,߬�=;���&�ku��6�fɷ����(��V^nz���)L���(�/1YYA�֭�L�(f�ɲ��[q�N�Az��{w۲Z.��vp_-�i�x�:QSN�c=�.�A+,W)�^Kf�˸
�"���A`w
_C��Rck�@kc#�1�k��� v��Q�!L*E}9�ϫ1Q�*��E1����/vָl�w�2*���$K���|��3v�^����5<0ŕ����p�4��h��媘t�6�F�Y�hܮ�-��z���R���8�X+���$�7�Z���k��,7�M�ۮ�tx��[wa�9�$�5#esy���b�Px|�gy�����s���7�;�N�V�C�k{�Ӷ�nX����{4'9 �z�z�����̯i�Cø8�=�98��❾�>
<c�lYJ����m����[sub5U��K���N�|ޢ&��$$��4:6y��)7g���� ������^���6v�¤�ml���Z�_(u�;-[;`q�0ќ3$�x�������Z�!>G��C�|�&��e�X��"�o7x�������u�@�\��aŪ\�i��/t\���i��2��j-n�Вqn�k�{XZ{�M�ߖ�Q�\� [fsKY:ܣ����'yд.�9��؎5[� �o��-�}��k�}��Js|�I^�R?rT��x���+v��= ��ԧ9;�F�U����ʚ;���M���!�7���m�}D1r*�4���|xn&�i���þ�/��2��f[�JOr��][�o.d���F���º��7D��%ڽ�����L}��YlM�LᏲis��ۖ. t7t�]kC�fK�ۙ�oS�����v�z��jjU�.��Ps����7+33�Fj����/Pn\Xo�OqN	���1�ٷљ��K��%Xv��t�U�SW����㇜��ͭ�npZ7����~��˒�v��Y�$=P��+d�H�F?F�_���I9J5�Q���PH(B:��o���kH�V��"�h"$+_z ���?�J"*�x��a��������`���8�Zy�{z��Jt�o��z�)z�1���z�/zɢ�֮� }a�w�]/h���p�(�A"l�==���e�Z�ᦕ��^r_'�8�!<]��K��&	MN����w;��[n^r���Dm��D�gxrp�]hK/��3�QaE�)q��:�8�W,�,>�{�p�Gd냳�U�ǰ�5��у�\G|o��%���YO�]���S�W�.��8��GDT��VX��5�<����&榨~ms��]�!/�[�P᰽��s5�h��:�v�ia��啙dT��u��M�!��g��xc�9�s�q�KE�4�kח8py�o^�:��Yc�N���wXܥ�漩�tx�R�|U}o\@�N���rÝ�)b�oHg�L�oa�w��®�[��(�!��Xu,��Y��|������u:��=��P5��|1#�V�W�FNG�Ǧk~
�I�OzWQ�*��$=AQ(V�A2��҅���ф+����-yeG��;H���`�^e	,tS�ݰpGUq
r��<23��F�fp[�s4s�*gE���Y�l`�-r��,݉�5fO���]��ҩ}akC�'���F��m[r�jlq][W��È��9Qt���{�c��rFo�Kr�����'���U9̒䊠��"�����%J���Iʌ宖��臥sM��e�U[X���"�Ӻ�MX1U�{��M^`�,n�2��c�A\��A��u��ͷ�iW6C�*�}��씿\��^���٥�s$�<��)��6iEK�<x�}���_l�5ZTY��:�r��6�=9C�սnЧ�&��η���SBr�]a��ɪ��2!� �F�s�LfM�X�r�vh':��V��~Y�4�[՚�?x�~��	�+F+7��B�r��A�fi��u�{,��y���=�%>
�h,�S�i����zJSt�;;F��~Ԓ�;�lE/�\�k[R�a=�>�W:����Q�D�rB�C�9+�V㋍>��H�ئ&��w`��dvz���敓�47ޠ�]�tѮ���L�h��Y4WMU��Kq��f�S���Ѡ�br�d��w:.��"7�R���9�{�0h\�[�9y�WسYoKKS
2��V.-!<	D8ź�h��0E�ι��x���'�U���x�t�LV3������	�\�����ɒ��rCNN��la��pL���N�֞P��G��gjS<�� ����ya4�dP��d&Z��^�gN�5�0T*KGOaL�SM'����f���uVc;�i�P���5����ZW�7��V�1�M&@N�%[�NM�p�y�3��۳g���-�9�܇%yX�Ӫz)	wLu�OE/��B�Fbu��'��'�s����QP�yZ��Y�	�G��4@\��s����Vy]�t�6��9쭒����V\<�c��=��3i�j1�-V�A���D�ܗǶ��fv売�ӱf���05����鎯�6��*]�^��V��כ#�f���f���{�}(Ws;���O�����G#�n�&k=6u-�5й]ZQץV�C��,YB�u�Oq��4e��)P9�Fu9��٦1����:]���(<�rfCu�I����sO.h��Br�݊:q�a�w�"�,� d,��.]A��,�wto	�[���Fh��X{(��Bw-r�&�5����ʅa�%ў��b�lfn�ܫNN�պy>p*����,�X]��R�C&��}К��w�tP`��vSi��R�xa;hTm�˗��:s�ݮ��Es0�����ǚ� O��jͻ��
b�RJ�f��\���ڣ@�����ُ*��p�y�v:�c� �ɼ���>y�vm�� 9t�.���h��[Me3 �+I]���Rn�&p�].ǯr��>��pj<����C�^��18�݆A\7B�'���o�9��UMpI���z�
��}��恥�+�ؽ{t���Ho{I� s�<�S7ǫ�kfu����r=�0��%}�	Z��^����ҍ=�^��^��{�]e���oBɎ挰�Rj�bܷ��L
��+@�a|�z�5p�N�;����2�҃7^�R���S�|gZI=3��Bh�!T2�RՉ�:r�5���nP�5گ��EOj���Yk�'n{��i�2B�[�5p|�=��m]_6�˸z�¤�蘉��:�{���.%=!��?o({���b�e�|��PlN�kS'K���{�S���q�C��sGVK��rۘ�p���镺	Y�W>e�NȚ�.� �]ɨ����9�����������@�>Jo����:���2d$�u�I�շ���>�ȉZ�6p����[��o^��^�Z���R֝��������[B)>����nbwC�\�U����En����U;
�1?xt�{���g"�,48l���V	\ip���[��4�[�I���-7p���k�)�f������������}F�MN���<�K��c��Y>(�g���	�͙�)�d�����!/-	6�_\��Q��4Gu �Bˢr-����Y(�]�Y�x���6�Bs2_\�ԗ��pt��� HG,O�.����;/���ːC��H�H%%�ݹa�V6;ln-}�.�}XP89'�7ye�O8�R�#ڀ����U�PC��U��Fw�T|v��/�OX����gS��(Q�R�c� l��#[8�m�rEOc��Z��;�"�+�k�y'�tX��y,�@�@f\�T�;3�F�i;65a�1���"�v�B�A��oa�\X�i��N��W�y*�NN�ƌ�m]өy���� a���˺�	 ᪔ͅDUAAV���h�ܩ&Zȏi.e2�l��M��E�o���7u��LI�B����b��}l�H zm+���XX7E(."������Y]�Ǿ��[��ok�d���t=�Pw(�3Fn��`�}��y�y�4tW�(�X�<
�i�n�.��X�Mo��UF�p�׶]����ގ���p�js��8�v_tlXt.[c�,.n�mN�g���$:wQQ���XH��5W�SM���q<����XTh� �����q.�p�H�gn�;�Ѭͣ}���,��S�������"��VL�ten���}.U�ِ�y��Ң����Qw�B�TF� 8�a�=��qR6�-�7.e��E���J<j\|1Ҡ�/���ke�F�-��G�V�?j�x9܇�����i�>�,�	��pʁ���=q#{�z�c͔$��!�wu|�ӂ�%����N����Wٵ�ِ�c2芛��0�n��Z�Y��	k=���g<ac&�ꛛ�UӜ�Wc��x�;)��uĮ��k��u�iH^V|V���hi���N;��v:=����{ZB���h\�d�J���|��%��5.��tm���+�?:�6��Ѽw�C�I� ��m)����M�]_@��L};Z�9\*�{&�.���5��jgkb�rq�z54w����&��)�6�0��0Ö��gF�Y�}�wW�"�x7ч乮:��b{��F�;n���=0�fWh#��!1�t#I���a��)&�&L͡*+�p�L�t����G �WL�ۛ�E�_C��Un�`�TC$�����-	�e�Ϸ��ĭ��4<�S���w���ı���ڃ:� ��T|���ܧԕ�܆���C3gpQu;c7IQu*�c����v��ot��#�i:�J
��|3�S��~�D��=gR�A;�I��wH)��vK&��j�_�?H�F6")��z��nr����6g���C�.�es}��ꚶ@�<��G2���&��Ϭ�ƌA�Ƙ.ĔF�8��/��{][�!�Qj�ǁ��cq�Y��z�;��9J\�� �q�ɏi�=�-�|{�m&�XJ�u=�B�\�a'�^���s��QG�h=�e��M��j���ً�:�;՜�y����ىG��&(�
�����HJ�*�(�`Vj"�{No���h����'b��{�ho"�ǵ�we	*\����^k�"�<��$"������L�H�E}��U߫/wa���Wm�+��<��WV�P|�<�ao\_����8f��#G�p���-�b��\�/4r�7J)�"C(�S��
��|�J����7m%���c�Q�0��IV4؏a;�ktMT��e���F3N��(v��+�܅�]� T�������+FjJj��8�#g��{L�w-�ޒ��Ey�yk�����h���l�Z�o��&G�nr�u���ur�Ͳwzd���xw&>IL�*y<�S�C,S-+
��-T���U�y�u��bQ0L �fsj]�lB���㥓+;kS�AWR�ۄ��}��dY��Y�{�d�L��j�Sou�	�B��XJ~��7 ��x��� �һw�Q�2��l��a�	����5�Oi�Q�	W�����<R�ú�9�m%���i|�|��F��������S{Ta����m�6�?ϊҌz�e�4�n�VZNdݫT��.�r �������엯$C����i��z�[;�V]���+T��9��6v]��qA�(!s���!K]�--����݄�so� ]���f���+GW�*�(����mfh�M�@*s��EAl��=/�9��|ز�Ez�ջ"ibM�yI�; �"��a��9:�thS�G���)�����x�:U�x��z�ݲ��ͳk6N�&CN�T���U����ۀ̇<$V%���h��]��7�L)v5�E��@�ڮ�����rԗ6�ۼ��O��9��us]$��N�/pn��+�n�)Dָ�L�/��2ݑ�Sݼy(�6;�Qt�'��t"���M`+�����_#ӡ���Q�b�	�8�͒���.�u�N�B���q�S�Lq�{-�y����rS�Ż[�ʅ��K���hc
:o�2A�0�=JY�q������q�n3f��8X�l���/˛��G��J�\#���{w�D�J��aQ��ư� Cf� �ǣ@�:�����c��Z�:��[^wN�ث�c%_UwZ��VF��I����S�����+ں�P-m=y������E�-��H,�����m��z.J��;�<�!�F5�-�8Y���{��c�^+��!7Ս�.ҡRT�(FTͳς4�$kc�b��v��c�έ�d�z؋4��:F���WHm��J�E��{}��m��GY��Ǝ�v���jD�׋|�®�y�oc�_��$���W!.:� ��+���V >�1.��s/��1qG̞+�DY�.?�@��H��[�-��2�h��%T�Q8����H�j�m��&�.���+ip�k6z�`Ja�����-첒G����*���/eYo�
��2V��s�&��nb�N��c�l�����}q%���iw�	mᩢ�um��R��T���C��:��):8/3�5t0�V��y�9�pw��x��p{J�4�U�����h\%Ն�ٍ�֑N�^��ɬ�[���jQ�����h�V�h	|@��F��q�7��^�|�pgnv�P�V�):�ijEV5,�3A08tK�/���k����댻Ҙy��Xٸ);�qԍ�Ǚk]�s~BΪ�C`�=����s|�f���}�·`Y�2b۶o�o��J��O���k;�ﺓ�u�)>��^�!V�V�Hb��ç6����Y��N�N5ś��:��0�YV�r���?uc�][�"��C:G����`S�iH�2k�}U���Z���x�:n�͈�\����:Ҷ���=���_J�lT��>�%�#w˝7��<;	S�m΃.�q����*�n��__ɫ̰����(�)BэQ�/{6G	�[��h[���}�s��I���<��X�际�6:�֐�d�IB�l������ͼ���9n�Է9l�*��ثer�'v�T)I��S�yf�x�m�C��{���[�r�:"ͬ���˩9����2N��G.3���q�,�⽃)q��W@G����[�7wY�����8	9^���Y��Fz�qBf�p=�nM���0�.���n������ю��;v�?A�Y��t�q�"�Z!��#{r	Qq����|9��SU�4��
y;��2�r�
uiղ2V.���z�	;����N�;���[Qź��'udHc�o��U���@݊�&�O6�uF�,_~�;i)ݒ^d)��*�ի �s���|¼�+����PO��ף W���F3�P=秋��.q+���#Ɵ���ն�>�����!��I�����kf.L�V���FY�m-���]&L���f(	$H��cgr�	��W�);��E5h^���ݴѽ��0n?���8�m!Х)�O(�́�:�E;�k��*��mj3w8���Ǔ��آE�[و�\S�橝]�
�K��A�S�PUlH^w`N\�:�w=;�R��'rCG�cȃ�V,+zj�J�P��=�xV�ഩA�&)��Ν"��3�'�a=��Zx���J��� ;��S8]�n�}���_G��/�n�Hb4��-(i�6c�v�`�Nܺ7ۥ�cSי���B����ؖ:���0�8Ş��|���/9q�̵�m-v�����;8Pw��݀*O� :�S)P���l܆�	B�ugn�U�wy�)wאhY�;	�@īߔ錛=a��ak&��˘hI�m�$���t��wv3��f��2O��s�2gf�],���8�Ҏ�ܾ��nWj���f�)�ڽ3������d�硕%�/@��>�O72��U�Nؖ�mvtkfvH8C�	��>��#�)�[�1������݌��Ǎ9��{,�N�'5�&6q��S�ߥ�C��67�鳋�	
�j$��am;\rh!Z��HG�]����a��ܪj?-�ڃ��[fG@:�Ykn��v5=-�����_�W��*+�g�����_g֞	�u<�C��}�) h1N.���@�s��+/4�;۴�����R�nV�k�-�E%�pV��Mo2�7�Ŷ惎��R�V:����r~���8B$�u���M��L��=�a�:�v,B�}�T���6O`���c~�V��)d=���ͩ�:�x֜_*����`û%Aè[��c;/s�h,��G��f�}qΩk��,�t=Sa����i���-�ANA�U�}އ�SAap���m�U�/�G8�oV�3mG\��c�8/4��lR�A����;�Ad���n�oU+��L�^�rl˦מ�k����=q�gN�e�*��M��fB�������k�÷�����no�.��"����⩦`MB�n�����yy��T=PJ+=c����6��]���оwA|"b�sB����啸�3T=Y�K�\�N�X��à(B6h��x&"QY�wgb%x{�8��e�D���U��,���������kՎ��!Ԑ"��%�^
��®�p��n�S�wt������Rl5u�C�ǘ���7˚Gg���7x����.V��̕	
�ΨH��6��u����3c���`�\���/�W�_;]'�_kf�n�!�C��i�v� ���g��k�� �h�4]�2��ʽ��/&�����u�H�-ҥh��{�۵�ARK�C2뢧�^���2:�{%�5n)q�B'0�:aI�'E��XA�ӾD��	����/Ѯ�QO��jYD�RluܽFI Y'y׆��]QK,�ʋ����֩�K�E˺�Σ���V2̵�B;�w@�̨�֊$O����<�"��Np��%@W�z�|'&���rP��#"��t�9䇣*���I!�J<��=Qr��^�99	���m%J�_W+JI-(*�=Ľ��MV��.�ˤ^gl�դ�O2ef�)�AI���:���n�9�P���
r��$�{�y�Fr��Ȱ���$��N]���B�IȠ�̑���ʯ��=|zN=�w-�X�Z]��BV�x���3��=�9^h����t���F9�z����uU=�<���(�s��f#.Z�VI�sB�Ő:����$�$Na�f�瓞E*�T� Z�P]^nҲUowM~��w��}9X%��Qǭ��Ւ.��}w�ݴ�QLi�3!8	P-{HvȠ��YKa��5�\Q��*�fm�-��_O�W�>�_%	��Ŝ��&�'k�RqƜ��2F~[c�_g���K&g�Jd��`��*�"���z��Jܒ+U��4Lioi�x����oӦv��F�W!�G�z���{:h�RY�O�*�P��Y) s������/d���,w��(m� lv�;M}�F{���<nh69;5��s�}�z����7���
mJ]}d�J�K�;˛�v�{����TYv)=Ll��a��^G�Jz��]c���6:�0���vZ���5������t�Ë�≿�����Ì�D}�n@��Oڈʋ��+�4'V]��ޝ'o�Q�[�o �����n��]z�E���L��|����;���g�P<��w��m)Z��ˊ&��o��m0�˴_���r�ͬ��Ŏ�o�P@�Y�=���A��ʳNB��ԯ�Ol_�	��k㢒�	Q~��{G��L!3o7�b�{���"}��t:���oR,wg�z(��ft��М`1֩T��i�moi�N'�ۣ��An�!oF���Kח]$�{+7ma���b��1�B��e�S����mQ퍈�6���J�c���o�J��K�ӆ%���V��G�B��w� ���+
�8h!��4|(�`�@uD���5�kN�o%��՟H��6E7ȃ�e� �uX␰S��*9T�XrY}Pmz�^��@qy�<�U�el�j��g|�鴚�e���KP�L���ud�bc.D�ؓ����!3��;'�ٱaOޮ�|���鿒>��}�{�1�<k���F�$�I�="zm�5=��]L^��Y�Jx-��~^X��L�I��ˮŤMǸ�qD������/'�3bAkE-�������Dǫ�l�/m�	�%�ׯɟq$}�-J*����\-���W�h����`�����5�F�"9(������i,��U������U���2��=xVY�ߐ�S�eA�$E�YлL���i-3h�6`f��_P�0E��^�a���wf��0)z����{'�^Ts�I�����5I��$�V� �2WY'%�2�n$v�Ul�~Pǖ;r" ���SO;=��φӿ0/� n�q�Y�@���R��ڐyyu�Q@��v����n��w|������du�*p�g���Y��GT�+��㋒�J쩌�=�pВ=�~�[�zry�:��]#�P+��3̽�g�k̞��O���]ڨ�@��4:�װ��|���C���HC�}�㣮�g��ܓ��{��U"^����W-|�<|=.9۹��Wz�f������z��^�)�ja�<=It��R�`�������Y1�f��{V���y��L�J2^�K�]̯e5�of�����eXґ�F��U�+8"xX�T���U�A	��۝"��Q�e^�|V�ӥYVB	\�(�a �7����fhW��y��2�g�O87xߠ�����-��þ�[�\"��H�KP�H#֙��"ʣ�aw��PA3\:��Ц�ڌ�|.��z����� �{)���l����k��Jr-�G:���[���4%C��b�w���a9�����撎gs�*��?y���OG�~�	�����&�8X=q�z������E c|J �����:l�����5����;X���1�R�dÊ���q��K��](O�|=Y��+K�jc��K�_?׬2��7YtZ��׏�fF��S.�|�Bs��u?V*6
��f��7������4�����2i`�^�o�k�z����RD/+X)��o�%^lH�W#�؅ҵW���B��w���ڝr�z/��F%. ��)�9�v�F;�HM\�^-�+v�ؐ��$��pW�Wi�6�ߌ��(�%Ĭ�� �u/���iCʷMm(Y44l�8l�~� ��+��δ�Ez.;��;��������^�o~�H� �ʫ�T�<�Jo~���jol5���.�[b����Oo��G+{龯zM�Ao��SV���˯<�yͬz��8'�G&ER��N:_���ޏ������~�74�W���n���I��I���o8_fp��Q�jص�S�-+�,JV�A��
'3�D��u�h�#�6W�������j̧���dυ?{V׍#�q�H�]zt�*��ŧիr���W�%�ٻ[��a�Y��N�ns�e?�맫#Z�X?1��|[Oi��f�(v�j�h�c���f���Υ�F�h���Y��,��sX8y�=���]�]�6�7[rջi��s�um�w�@�,�=�w8S�\�m�{Ú��O�f�����l]��
�����Caq�^��XIg�:�ӥHpH�{����D^���o�?n�÷���Ụ���Yryj��6_ޗ���;)����eS[+��^����~b*�u< �h3����J��~��ϧJ#�GZ\��p�.��Լ��:�KG��/M�]q#�
5��M7sʱ����q��;��7���^�Owl5=�&s�&�ۧ�l�	�W;ÕY�H!K������ܛ��"��o���h��/-~"lF&�G��U��fO�0z�TF�RC��}ں��Ԃ;��$RYq�K��z*v�]��㗱��H}�\&�z�eN��Wm�m>�(v��I_A���o��%G�GX>�f��Z�*��ΰ#2W��P#a.޲�襧�!LrPmtOxO�a�]Ƹ(K���Oq�5����C���]�<|3�w�#�>��v@]���r�AU-�M���;��JS���E޹F�*���&���<EY������6���{����ҧcM9�H�7�M��y�JL;�s�����C�g�T�9m���@ʆ˝����g���8)��81	ֶ�[�D�p;Bmg_Gs)�����#�3�y�����7��tj+YWMה��ܼ+�(�U�N�u'��{7}ޛ]".z��K����������/���Pb3���u��K}WP]yM�n����<���jzC�} g	�F��)W���6���_z�������K��g�{�}~z�{�]`v��ð.��%H��������pA� $x#[W��ޫ
;���/w����Fd�H:n���fEFk5q��NUӆ{��[s��5[է�m��ʳ��&���I	+���*9T����z�/yW^�q�<��x��Vg�s�|W��`�6�� ��������ʯ��ۏ�O��#�y~�3(�Y[���w#���R?E�����Ez|�=R����I19�_+����2�q�ݾ
���W�<$w������܂�=�Xo�oI��oqe^}�{rN���o�7��a�ܽ��(�ę��-«*d8d�����F��ߠ�]aOcx�;�OHu�����CĎ]J-�WS��^��:�ʐd�A���u��u��v�o�h4ά�K*�Jm�;��p�Ԙ��p]}q�ίoz��y*�2���Kn�!��N�=;�L/e��!EK�.��c�1��\��k"��w��D�z$��^̐���n�H����+U��&����4�|�̈́����N���	g�u���^�q��]<���Q
��y�򚦇��F)�M�^�{M�>��_}�vH9��F}��z7�$,L��Y}�)��t�ȩ&��=�m������2���M6����.�����q�k����x9���]t^�}hm�Ԣ�I�>3K�1����E�����!q���j�����Y{=Ub��K�8Q�I(�9x-X6��v@�w�u8��K��5����6�'�݋�:������߮/q��U��m=�y�]R�r�z<�f��P�=�������'*OW=zR9� �ʣk�+8"z`靉��K�2�/f��ۛPK6a��s9ci[^�S>�t�ޏ��wl ���l���\�3F*��λ
7'�Щ|%��L�oEx3^�	��omF����!|	�傭�����c��ݵK�m�ݸ�S���N7�c�{=q�kȱ����ż"�pۧ~�j��㣯��tv�*��ZAP��G�T�<��N�}&�M'W��;�,WP��]YK@��ãܷڅxrDZZ�U�g)�4=݁�V|ق���xG��m��U_!�S�����ޭ�������"-f��]�3�E�-B��{�V7!W�q8�K@�{ط�%�X��&�d�T�����#����Q��b�f��I���5�<���F���g-�>����!w�X�'���i`^V���^��[��C������z4������
���+ ̈́(v�t���%���QW�����^�g���Lz��=S�ez��_�]�Gv��(��[�&+d.�Xr=�lY�V�	[��ḁRB�� �1o�^f�`����^�or��JRA���tv�E�7��on��z`�7��d�rt:��=��S�bKN�2|Ww^V���p��=S۝\/TfWe�@�<�c�V���vu�]�/y:VSN�1�b�ݬĈk���i'{Ok_�Lm�MC�[�2�7�w_pX�9����gy,�4��~O6Y浟�/^ԜD����9�����u3�m)�/U�l自q����&� ��e�j�]'�^x<��N͞^�mk�U=[Z���PN_�o���ר�=|n���R{�jd�\�| �2Y1	�K���<�SP�׳ɚ�������j���*{���O�ew{\���ו
��Ǭ/X�=zR8!u�Ң�`F�=+��hTY�^ĵ`���	<�ʿgo�$�{���\
����wYن8���U� �|�EYޯ<k7쥖+�3t������N��o<��Vfi�� �"��BIzw�|1X��6<#���0��C'�=�|{+�IXm^]�_/X�(���,"E��Y*�\H�R�JF�]T'v��E��Մł9z�4\�{�Ҟ�����z;��!V�;y�W��Ƿ�7��y~�M��X�׭�;�`�ѱ�J�9$�R�w�ݗ�u~�^�^l=���������,��
��ʻ�3Aܺ�m�0��*;e<���V���4��{{�����s�;�/N�˘t8���$�+���	��.��0��:0]�)3mS�um���굌�<_.�	��C�:	��MǸ�i�ׯN{���6b�4JC�H���J�KæM�WN��|WZI���}Y��y.NĊjRqD+�(ӢoFz�LJ���-C��6}Hc���}��v��${iRR�*����y�/Ok�ޓ�k��ؐW�@��a��r�V��6�z��fo�+��Y���kkS���j��D�}�p)�ºo.(��
�H>�NX5;�X,�/N������b�g��M��"\��ni�7���*��\�j��=ۻ��n� ���B���
��z�W��|}�Z��3���u|7��q��[�i)^������ΜHC�H����ŀH�1sXiTU�駴�Ǟ�ǁ��r9�xE^f��B> ��8���<�Ѱ}�$R���j���sjt.ƅ5���DY#�ɪ>�����D���Q�%EL4U��z��g�h�&]��5؛��L�V��':�%��:ӹ�OtZE7�����t�l���W����8����ޗ���=��Q}�2Z��`�a��,Խ�36�Nњ�t��D�����<joq'���G[�byy�1�����C�w}�x+��#�2����n=�����y�}�Ր�v�Ec��vˍ��)���r�N��)��4�V�G�q��=�(KЧ�7�C����1=�-l�Iվ1P�����7��Ea�?+���s�AҎ�=|������(L7c����I�j�n�ܱ-�Ӹ+�uk)�^ȳ�X���z�c;�{B�r�5%Z��Ϯ�-H�k�{�v/7���"����N�����j"���A���q5�Ѓh{��ã�&��/L��4E=���ǲOy��4� �[;�r�\�{Է���p���v�}S�"[慭;vf.�n��ٱ���^^�-c�ؼ�M���ZR����2x`��dT�ayu4Ղ��aԬ͑�h-��ܖ���l-���{���;����D<)����AZ��� ��Y��D��=�1���Y8�Y�¡�q��*Ft�J���e/�(�y� ]e�ϭ�p�e�Ρ�S
��|Wp��jwg���v�TJ	Y��x��o�â����ӷ����G��&�'�5�/��fm���˸�� �p��هV=b�6�z��u� ��C0,I�R��Z�[��K�����)Dgp�;iq�\1�PL�9B��˓\���ZsaA��� _�#�������ݗ6��Hq]���;��q�e/鳺�鿱;��˲�Y��u?��tb:Br�������v�0]������v���c:�\�CB̫��m��(-�
ɐ#wWg����%Sߦot�y3�(�b�h���KZ���׭���>Y3t;'�s�^��ٛ�DjWWM{�[x��]���bh�pE����|{�{ʬT���q��"�ĳ���[�1��"rA��k�u�v5�Ou �T�=@�jO�\�Ʃ�x����~ ��Lu=�����Ǯ��w���R�=�b=����6�B���E�i�ׄ�i��6��j���������aݚ�D{�Щ��YVH򲚧���c~����խ4-�@Bo��Z%��އ��{�d����)$���0>���YV�^̵��W����R�зk��!�Q�tޡ��Gw �Kc�՛M���J!)D��ae�Y'3�j;w��fX{��W��K�8��i���E�|޻���z�ACܸ"/��=&J��v����0��=;<�o(i�poN�w �;�p�
&96��#�H�TpT��X�ؼ
�:�;ˋf�I��oc ��NA�'�=zz�����:�V��<�{=�l2�0��n��#�Vs�������M'ݜ~:E?S����czi�i��f�G1�)�,7\;�:�;���|8v��|>����r��*�����r�U��(�*4�:��F�&�I)W:%DW_�=3��)�'�B/:��g:t�$T^����*E*,�9���$P�B(��l�uE�t�3u�ʜj�Ss�9p�:�ep��D�)�y�]:IP*�$GH�E0��L���W*�WH�A*HH)��^c�qΑ�����r��T�B�$�S�U�V��U!�8��b��B�ui�v�]f	��YQ�GS�'<��K�UN��KYq�:,�t��)�% ҢC�%!��kT©X��r)Q"�dT�W:��!,M29f �[,����O/�]�(���Na�L���w:q
���DTHPd ����+6Bs^�9�%B���¢�P#IJ���N�*!�� "R��Vθ�����U�A'_���ֿgoFF�z�%�$ۋ�s�|��-��rJ�qY���X����&:��3[Fe�����Wު�bs�Y	zp�z~�;+�[�+��ݞ��J�ĐؠŖraG�������\I����N�O����V���lm��[���{���V8Q�q��N-�ժ�67e�`�s�_)A=����^��<֨�
踶8��_�Z�s�S���0M�Gj�b�:�]�ޜ6�K���\���M[��)���6h�0.g~�Z%���{���3�7�՟X�Ÿ�͘n���.q��	{��G|#!���������*�����U�I�y��`p�c,{�Y^��W���@�Tvݩ������20��jw���:j�a��O�>3�.g�V�������~�_I�r�����1a�>���]�sભ�f��#��8�c~}f3��m�2'뜖�Z�a�=է;�u��M�1������G����c�<n}��)�����
5�:����!����yǤɾ��W�����F;;,�9���b�\�ƪpjpZ�9�����K�OX��Q�	��x�w�.�<#߼��_Blp���r�xcuSSK����?%������t �7���3�P��j��z�!��ND��r�F[��n�\�����:;ۆ��R��ӌ���#�드oVשQ\���օ��Z�e��]_���R��6��J�;o��떠�D��N:��+��5
df�^��ȺC\�s\��{��{ʯ��P�ʕ�JX�ϦvY3񮉁A�A\	&lTÒ���^���\���G���{3*��*߇n�W�~��]H�F�FE�#�_�r�:.t��!=��3T�J�Bٗ~���tݓF����^���D�pU��:
7�v����h|������A��B���~�I}�i�C�n��9Q���Q����f�^@z�X]�:����F	�"��#�C�>��[��we�٦�z&(x*Q�}+�9`�z8��7��3S�s���>0{������W�~vp,�]n�Z�W������`x ��|eJ���|,ߠ����o��E�+Ncͩ����nT_Ԓ�J���ry٫�fY�e�n����x>b@7�iSɇڰU\�]���a�{�b��7ܮ�u�$0�!�7�B0&��>��}�������P���M͎��X6��S�MW���5�/+i�[���
��h]L9�"�p	��N|���=s�+�B!�#{��R���y/&Ύ�z1�v��fb��n~��~�<]c���������,[R�M^��Df����ϫ ����y'd[|�j��9��yc����n��/t��>���i��]�mb5dV�9��{��/���H���zP��o��2kh����zG��]6z��ס�N�\��/�2�h֔��o[c�t�d�kW�R[�����+f9���6H�xv��
[?_�J�7�s��T��B���s�U[��n�5o����}�j���P�׆��_NE�����ڔċ�WR���B�T{�X���SA�~�j�s3�}��Ff�U=�����O�Z�����@��A�B#�u(9&� ��P�x�ʈt�{����F���]����>���װ\�3;^�G�6$O���ԡɹ�*�X�6�Y<��3�)�����<p35��5p�i���	�����%��kT-=�����x�C��Wg�=�.+��k���5h�k�7AM��/gN?U��i7Ӝ�����X�]���;`i��V��jB`@��O��P0H�,�վ�B4�Jt��h�IHg��ϛLQ��vu^<�ߒW��+���}>00���ˈ}�x�c>�o�f�ғ���0;������� �ϺC��?*ӀΈ�j���	�ynM��>����G���NGZ�D'S�c="��3��f��%s������|�V��hlJ���h0�_�,�����4��+�^#�����)�|֪�A�P�z���!)�=~9�(��-f��#N~Z�+9俰HS� ���g(ǩ^��ű�=��Ko��pT�Bnh�z�q;GJ4*m�0d+�u���jE����2=�e��"����/�<��17Go��ev����|&�q�������u��[ 5{5:�D��]�Z�l�Hj�>�{X�/���E�ŊX̭s��l[3�kX��z�S��Xa�GmvK�S�/Ʋ$��yPǾ��vwz����18�]/{5���1���3��N�3��b?{-O�<k z�Ǖg����;�j����L*ȟ	Q��¥��H�1�^����p�1n=�a�~v-�y�鮃�+�,=�:n3�f�v����T1U�h�F�vg�!>0��>ϐ���ٌ��L[�@�o:?#����8��N�ͨ2�x7Ezf*V�~Ukb=��ಌc��@�( r=퉑D�s����7�<�o�l��p?A����p0I�22wn��	�
�=U8�Fg1�X���;{y�E�Ƙ�o4♿��9p4�Կ5G���3�>}K�4�Vs_�k��.)�ō}����D(u��;��k��Ԍ�ON��&
t�g�ک1�Eș{�s^r������he��%8�P%G��1]>�r���Q�K�n��T���L��x	����[5��W���������2���Gv(�R$�0��/�y�]��}����ϳ�w�a:k�ٷ�Ј�qٗ�`�X�&�Jr�VS�2�+c��Ugo.�<�燽3�YT��؂�;a$#tc��c{����(�I���΋��Jr�݌��{�K�)>�Ï�E���Y�!ฏ��c@������A�Q��;���LV<�n?a���w�x<2Lx��˗�q���A�[R�A���]�����m����K>7�+�*4{1�>�z��y�!Ү|�o>Μ	ݨσ�w"�0�P��	��SCin���Q����jHz>u���s����&鴤���Bq!@�>	V|�NB������%@���\ϰq[�������o7� ��e?�	W��@w8U6'>lPb���������UeI����N��NV�}�r��K��qq`hT���`��5�:��,p�8��"/>^�`o���R'���u�x�3u9���yY�~�^��-3?b�1a��?|>~1�L������ˮ�3�y�<���y�\7���{�>G֯��M�;�7[C�'��I���h����+2~��#�z��
��3�#jۄ�x��̚�.�q�}�q�?;�:�}���^M)����G�xU�~υ͆���\=M{t�w�S�Ӷ�����`;X�L��5�7(��O}^7a�ņ�++�
V�/#�?�~�:vs���:����;h�WOX	�IO��6��boV�o��^����#��N�,�8��>R���.�A����&o߼���i[����8Ѹ ��
�f��-���XZ�ݙP3P��;��WΆU�G����3U	��N���#�|��ξ�кWC�>�E��^��,��[��>^�_����5V��UV��ld-mc��}f2}[R���4[]����<wgx/�Q)+�9�dCϗ\�k��GvԵU�&b����1/�#|��1δ�of7M?\�wFp���J3�M�l������n'�uPF�pjJ�r]9^�
2D:����]���'�X��7��0��^ؓp+���_�(�Wɽ���xcv�����l{Zoskg���w'�Şk���U�Y���E������}]�~h�+`�-�N.�z����ox�`�
^ln�M�&7����n5�=���[3l��$�b
�~�^c<�.AS��r-����/r������K� ���w�����(��3�P!�=��)򝛛g�����p���8ڗ�9P���X(����-������X]�:��q�t{'ޒ�]&*�9��3�	��5X(��0�Ł��]+�,oGf����jw�cw�������{�}nO�u!��V�s�٧�*g@BEEp�1e�/�o�vW =�yp����F���˛��_1�x/�k~z���^�?v�S��=y\j�dA���1lu��O�w{A��F�w�
R���B���}�:�����^|��{��s�d�pgd���w�͑ף�Wl�P�.��Aa�%�����$����3-�����7$1ۂ�L��xp��#}�d��C��l�������-?�l��u����>�n�z��+��}m�5�o������z��߭ϓW���{�X�SPĪ��d���ܗ{�§|<�i�޾���p5�՛Ƙsѫ��9���ϓ9�
�ϣ �Vԭ��{�{
���p�5��'�3�XɬS4�C��jL��<]c��ض�⁐�kbR*4�Wh7�Α������DՊ.��J�7.i���\�}n`5N�UV��o�{,��n�����O�����H���Oݎ���a�����ƽ��z��dP�*��ܱㇻ��=>]���Ċ�}ޏx����=�9�1�|�Xѿ)��M@�<b�9>, �P�{֢-���4V���f��]A�������j_�&8����l����G�R����A��R�>M�*(�J�e+��"�z��g�c�ؠf�ݚ�����	5�Z�(�/��\�������n�鮏���B���V9J����J��7Jx�g���,�y�m��1�'�ĉ����e$>:���J�o�$��N�h�۱*cƇ�G��(��z��Vs�Ή=+�פ-�7�q���ۨ]f6dB���P����n��EJ�.��q�z���Wy)���>m��m�oL�\�����]H�����m�X6Uǫ^���7�M!�߄��bLe��
/��ˠr�����4� ��3��S���%# B��Ǖ}+�-8��5a�5:&M�� O�W��Q��+����@�Cɼ3W��z$;����$��L_�	��0Ԍ�����s4T&�S�+j�'ò���70{G�%-z�����>�J`�x�0�c����/N'wQapv~�b��O�TH��t4<�SS��q-܏���?~�~[	3O��txP�(%��1F�	�~5{5>����b� �ƧF�V��M�$d?��-Ƨ�/��cS�N�f��5�<b�8�����3�}��.0�mK�䍯K��/�&�x�5���Z�V�]"���i��v�j����N��ߗS�?{-�#"r���Z�#Z�%���e�R����O�VD�c��R��H�1�^����p��-Ƿ�8y�B�r2\�엱��Oq�7e�Gh]��n���2��_��f!>�Q�60�>B��
}�6w��.c'��a��c���Н�2�x7k��N}�ޗ�V�(�+{��4����k�a���=ݰ��J��ƻ�Cy�2���{\�[��8#JIˮ�y�*�.�]�l;������\�~֮��$Ut{�,V=�p������̸%��w��Ef�s����ť	�^Ƥ!�s�YO�]N�S���&ayE`tѭ��1^�Ϳq���1��,��]�/�j�~�YX�A�2=;�Npu����#Ȍ��������j��Gn?W�VK��<�ż�V9�k�^[R��B���G`��Z��h4"�9�"������}�43\�t1HS����g˽���R35<2*�j�rcBt�`ک0��s��l��5��2G���%٠'n|���B�][��,�@Q�K�n�S�R�$��s�-^E���K�>,U��C\❑5���o�}R%��켎z�Q���΁V���F�����]�b��)�g._�ի���p*���@�A������FN�=��{�GO������Sr���x�%�F�5�>�9��C9Q�h���Dg�*C�5>#�1Ѩ��rY�i]����P����^�jHS�!<���xNB�tT°j�[j�O�ޭ���.OVr���"�!�ŞRnt�l��ݞ��p�nDF6(1`�Ex�&�l���K���������
�cң�.���[ӫܱ��"/>��,o��5��\��.�#�s�r7{k~V�A��-�G�3�c׀�]���yָ�����$�,��BIؤYߠ����a`�g0w'O�z��X�g��
���wa޹�]�J�C����͗PF��Ųîy�Z4<�qa����_lnc�Ǧ_^�Z]���^�~\]&lj�1a�a���X���e<��ԕ�{ɼ��lz��{�ׂ*��4#j��K�����̓k�7cU-3D�%���8����l�n��3/E�Q^��D�o��?1f<U1���xo�3�k}86sf��>��X��I�ʐ��3z3�(��b;X�Ϻ��j$�0�0]\5:���s�W��oqa����iu����U�����!��*�� ��(�(1��Ҝ5V���LӖ�f�Bm[��G�aӛ2��y"|+sw�Q�ҽSl1_O�DlX��#��Ȇ����u"�����*�r�����ٖ3�qž�p5��G���<U�Q�n���qFr���
1�;��ͫ�5gY�#��u�����ԅ�Ug����IU���ؐ�c*l��W�Fě+��o�?B�lp���������= b�Z�9S/�X�3�}�=4�+�RT�.6g#����5�02�I���%nQ^>�AU9G'���߆E� ��}Vo~�mɍ|�l�k>��.#���A�?1& "�<,`"P�B7^9��%{��X�����,�J(g\@��#�nkc-�7�f���c�J<��������ծ�zwV�d=`�����5�	n��R�=z�{{�0��c@��S�p�����}���ޡf�îV�c��]F�=.��T���7��7�j��a��1���假S����"huw�3�n�GȽ؇i��ҷڋ�_t��+�	���TsR���	ߪk�q�L��|	V
mq�o:Wٕ��Fa�s��pQ=�v���*���&�gV�iݴ���-�z�khehSk�s�6%��on�C|�2٢5Z��e:.{���Ŋ=��^�od�J���r[�/M�Q���z
1(�ٰtF�4M�'Ez��B
��.��	"b����f]�uehÇ;{�261|�S?t���Ϧ_G|��};]\��X�\Rg�g)���no	4u��sN<���d���� pE��+:L��y6�β�Z]�����O	�}v��w��(�ݑ����q�1ڐH2�d��3
��S�H��W�'hf�?��
s=꥕�Ӕ5LG�e��j��WHq�O$S�����ڱ�Y=�:�:7�R>Ův�H�)�l������;������-��f��M�ým7�*Y*���Q��-U���ݦ�7Fi�/V��Vq�5f�]
�"�����Qj=�������sa������ٷR��a�<����|L��/,m�zZ�͌M����7�X/�ORF,ʱ�#��{�Q{��fl�vĵ��M�}�7_U���c�s_�>��ݜ�.��W%��4`�'	\���XR�+I[sH&N��3.�m7�qq����o��pG�)@�����C�l��,���R&��N��@�Oe�����uM9ĽwK�*v�V�٭�B\yb�MG��a.����:�p�4�q�j�/g)ݵM_�s��.x&o�I�(cWo����m��M��׏"�yw�,�� $Q�Z�P�3�����ݕ0�}=��ywC�`�.Y*��_�#>����2�6|���j��w��=��5�/$vs9�sF�\�;�N��Q87�^]Q�w��Pdtx�ټ�_l�9�u���s[��m������6;�z�U��oiX�SZ;3`FF
�o�b�Ho�x�٫<�$�kw}v���>��pZ��m��P��Y��7D�B���#�ϳ�I�FgC���U+v��j��8nw�/���՗U�8{:?%�j���3����t�9Ft�x\-m �7������Ց�X�ZЇ������6�y栚�O ㇏�NS�+����6	�����7I;y�5��Dp[7����`��fY�j�Q����3��B��]�����o{#[�*⮮u�� ���m�N�)���ޱ�4�@R�̆Yu�Ҕ�����Р*K{����
�p�ʃ���߷�AH�H?�h_�2U�C�t��9�8���"��)G�"�Vja��D��V��%J���\I(�]�dt�a&WҲTBN��VX�Ђ"添�\��W��*�ѥ�<�P�LɗB�Q��#�dSB)*��ѥ�)-Q$�5Mj("T��)���I%E�V�#Y��

}�τ�t��us�DS�)҈.-[*8�B�E
�ʈ֪d�;(���!K��Ar���$�$�$��IT���rOo7Y*�DV� �"�uiTI�hv�R哒�T*U����\����EMʍ��"������aEafGY�E�ɚ���Gy�p�*��m,�B9�s�QDQ͗(�bO=2"�T�;�^��'��8fȊ�9�4�"���Ut��4�!��\�C2���>w�o�����~Z�b&-����¯-� �a(�W���S�-q����|��Q���wV��x���ms���9h�"ͧ^��V� z/����k�pun�
�N�o����a��Oh����=�tAU�3p�i�Q��0��M���믜q�*��X(����-���ӊ�'X�g���/a���xfx��ނ�yXHaE@<�/���=�x��f����jw�`&��G8�î�^�l�	�p��5!p�s�f�i��"Lx ��o��Oy{0������XqR��}�~�HA�\E����n�����ߗI��`��|��<����Sw��
y���g��5�{=�c2�?��3Y������P[��	�؞͖}�Q^Yʒv>c71��u/�~��v�&_�6��v�g`.�o#Í0�WSs�t.�z'�F쭩H���Y#=W���No�����h����ɬs���q�-O�!�t��/C��x�dF���ܳsq��u���κ#��G�N��������M�?9��Lv�F��s�*�r��OW���e�ޏNo���akq9=[�������|p?x!A��P̈����>j�X�}8�5�]_�Sª񺵨��8�����=���1�ȇ�;�K�졓9GqO��pA�71X����5�GW�Ŗ(����o��౉��{[����R.��z]u<���;/2��i��:��#�!Ѱk��ӯ��7�z�=�,Ɉn�$1��1��}^�6d��ߌo�GB],�������NL�DЀ���xc_.��>)���'9؞v{�\א��K*,j�Nl�Η��&���l�R�7�r� ��	˺S�~��{�eUY��c�^�Kܬt)���#�fj�f�vS���?{�D�i��*��t�{��n�p�в' �P0��Xe�Y�5B��S�oWA�W��;�z:j"ښ��n��x�n���D��	P��1b���;><�k߃�} �m���)�k1M�U1��הh�_p��GNY�z���сN��B�+�u��+>츇����o�ŕUI���W^}�݅��b�:ڹ��O.`f���:"Ra�_��OC�ܛ����'�^���*~ѻb%G�Jq�Usߞ8�)�J��
����V��hlJ����i0�f\�.�߸?e�ƞިO�%Յ��@b���70l�hr���N�m�\'!����,B!k{�.�.���/qWٍ�)}I[W��8-j_3xƧ�N�f��5��aK{A�K>��� ��b3���a["��n���*֛�������q<,�xg�8�@���߸.��5O�F�x����p[�V��s���w�fzv���������i���1ܔ�r鸯
t������V�e��'P����Z]Ֆ�\�嚲�U�{��� ~�^�sҍ�ԯʲ&��Z%9�z�K;�cV���Ϲ;�WS�?{%{�U�\�G�>${���$������O�5��]���0G�H�1ν�}�
�N7�`j��ʣ���ʻ/?�P�V/��$�����������H�'�]c�ȁb��Q�Lt��{┼���OP����u�w����y�/y�fs�����4*I�MԶ'��<v��/V�}�׍�|ō�4�g�>�7m��SW���Y�k
���!A]��Z��խ��� �������q�t�9�Ѕ��b�X�l5�\������d,�y��*Mʎ؇ޗ0}g7�̯w����~^-,P�'L~`�9a�]�-r�u#3S�S�qɃ�t�.��ؕ��F4;�]Ԙ"xȞ� Wʾ�*:,
"�v^)z_�(���OL���}4&��u�b�	�7��f����Kjrq7�h�4$��N��Ե�D�����9�(�l��Ѝp�Ѕ�ql�{��y����KN��nw�j�g��q��*�V D�A�5�T��1���3�͎3��n��"׻��Aw�w:�ԕ;�C1��yۓE�����܄s�w����Ҩ)}��ؙ���ޅ�+�,�������{�#,e���Y���Y�u�e�9����$}��z���]�ט����'n��Mmd޷PƬ��<�S�,m#r��k./����g�o�s���{i<p��o�5B��Nvc;qh��aP��	iF���i��Q9���Y�\��r�{�Lu��ړ�}hN���*Ϭ.���Ss�U�{:�u'׼��=�"2�)H��Ǟs�r�e��U�vz�©�8ؠŖrbƭ�dʵ"�#��4�PWz
_�J5~�
c������yX�zur���"/>^�\Z�.�����r�xovxP��>h)��_*�-35B�������:ɖ��U?NT;$�WuH�@�����T�A�\G4�o�/���9������< �ɟ�Z�տSU�U�dU���g��:�j�O��u���v�>����]�3[�s��@\��I��ZĘ���8��B��1mg��]3���G/᫬���0�0�`.��	��{mc��흏;�C�v�Q���������aV�`��1�sF�|��c�npUf[�|���f��?6��ŏoE�j�y�=�����Z��ڗ����6/�i�AӖ�v�0�:���7>UX�9�n���y�`��������L������E�]j��]8z�P����T*�27-��I�{b��_��B=v}�qfJr������iG#�+��u��ݫCCI؁����J�oHnB�ha-7zv��6���β���pWS�p�'�غ�ǃ�4>�����'L��`R��W��LPc5��Z*���`cW�(S�ϻ,�8_��S�.wQ�w�C��z���:��r��5��ޭ2߃�	N|S`�W��&�
�p�R��`t�3/pCȗ�y;���ܠ����7�7G��
���i�����_J�h:H�zQxs
�I3��D7�+oY�kۓ�5�70c��Ռ�)^F{��&5򵳚;���BsU$N��dt������'gM~���8<��Y�SZ�*�����!OC��F���U�3৴O���l{3&clPEܿ-3gPs�D�bh1J_��9N��rpy,s�,nBU�i�����z�y ��ߞyYV��g�)����/��<h$/�)���E����|n���f����+Q���ׯ�_8��q+��Q8�T��V��7�KX��H���m�����Y�A�G}���sw=q]�Ș�.�W��숼�h�bw�b3�}��ߗI��$�`��<O8����B�Ў�t�"JPz,���/3o����hߟ[bF�X�7�BU�;��dy�+�~�/��i��*	��*�f�e�;��J~�e@l��o�lMlɅ>�'/vu��2eD�n���b�S���v��\��:�,���hQ�RB�XyU'���l����=�U_(�m�u�H��q������w�]'*ɋ�zf���]~UÖb��3�1Z���t��;f�f��a�F���s�]�����Gg�j�׷��P_�n�&����FDF�#�V�Go�5�c4�C���S���};�u�[�b�`�8D�K�~���wx���ӵ�I�ڕ��,=?�Bn�O�F�"<'d�����}�{4�cD��nvG.������>�߃لA��W�8>�׼����}SD�����q�x�w)�Uڇq7�u{^SA�z��9ͪ��>��')2/��a�x<3�_.�ϓ߹��uv;=��k��$"y�/M���*4�77�{K�1�b�.�3f���Xf��-�=��{tgz�h����8#�qd�9W��`šv8�U�5����j|�e@��b��{ؠu�ُ|m��*\�1��	Q�!�S�5�^��pj�*�H�<P�X��@��W��3�Ӟxg٤�+�����Tr������b�����������][�afL��D�:����΢cJ^��}D��tY��N���@�E}?1�b�,����'۝>#��#�����+�e�~閩�e�(�_�Oj������X92VQ��F���׉?{6��)�|OS�w�w@Hӡ%����Pe5�J��ڰf��=P�I�_f�_>�Ȭ2m��U�k"CTת�gUܘc=��h�fQ�|�]U��Ɨ�>
�ա�Գ�k�Q�����e���=�8��Aw����w1��'�
1���V�\�	��Pڻ�I�ߒ��}�>��|c2�Aq��z��<��V�1+�>�]�Z�[�S}72N��5%3�����9EuW��/n�e@���R���/P�߹XHIr��E� �V��j�j1���6�,tG4�\�/X� �^	NG����>���ޝ��j���q���Xa�A�<��3���j����y&��jNՑ>�f�ND�޼R�ݳ���#ܝ�ӫ��c{^��q}��,{kcI�;����9b2'8�.:kծ�����2J|h?����A{��\(���a6���^�����Sx3�XP�?<�E��G�(�t��W��V���j��	�Y@�=�ѫ�5���ɼ��|b=^xC�V�!n��r������^��R�v�V�~W�c@PB�b�Ѿ՞����������n.�pE,<��ݷ/�j�`��?6���"���F�z��SL�k�MK��ڷ9�o��F�f�eDlʀ���!.��j�3cMc�K�jY��G�3��V�xs��<�*ȁ�7]�v�a]9��V,�c䋸���S�4��.H��)���#�Rv�e@)�F;�%��{���{�7\��L�s&^�`���*r0$�+�4-�w6��q��n����g�Ar�ۗ�ޫ���}�v'���戴\׺Q����Pۻ�"�\~C�#�$J�n��}�,��c��y��8��j����}���2xUq���z�����Y��k�/������GL�t��/�_�(ϼ�`����LD��.S��yE�KU,q�2�q�&s��eFH��H����?l�y'e�sj�jЭ��`R���Q�&�.�A}o:F�IN����1�Q��q��*±$hM �0U�T��lY=��Cu���w��;p��G'�Wճ�]����BS�&�TGf�)�㮧�J��u�y\�Ø��c���<��Ò����^�jN¯�	ϒ�*ϗ	�QR������nB��|��4v��<�xS�;��9�ŞDWNW���J���@w8
B܉��{�ϧ�1����;9��}� ��F�
_��ktרc�1�~0���MYn{�5�:��(���-�K9>[x�g=ޜ#}�@���g�Z��U�z���fP�,>0�??:ɖ��*����M�	������s�ܱw���a�Y�[������ȩ��8=9�Lй��D�?k�r��t�q�~@�{h�)*��3Ή!н{��,<��%�E���a$�s�4S��z��x4�^<�;�XOGN��zn��s��BJ�`M��KA��R�a��v���CJ���1np�,�=Ut�O��y��Xf��Խ��ZQe�n��:��H�� ï;�kil@�/���}�_V}|X�.��[�s�<7��w��U��,,��ʞ��ۃ�'���m��r��Bt����� ��jH	��{���6g�v+�C�JuPt�����z�k�+Kߨ|��79���Ȱ��%<U�n|U�z���++$��11�5>�s�la�O#�'k�ϫjV_MQM�Gge�\�k��Gv���k����o�/C�|�Ӻ�lc��`�k�pO���+`SW��D9;��B.�F��[�Cy,s�������Q��~s����S�2��f�{�lI��X����C'��S���j�J[���Yv�S��͚k����1����g�g`⬙��&|���};䭋�{5��'Mg��*c$��1ʥB�p��ctq��ƀ�Z��u��]�{V��u<�� ��;��k�C+�9ؓ�	Jn��8T� ����8�U��to����a���4V��/��{�β�Iw�~����D�%D�b�(��u��M�9$y,s���Up����"���q��J���e}H�jv#v�j�v9��p�N�ټ�罯�g۝������!wd�8�cˁ���5*C�6t�b`o����)eu"��l�d�v�pu=�.���݋�Z������s�뀩S�U�-J�}FkN�vb���75�;�2��NR�F�����ǻ�5�L��}YъH�q�)�2(��������E���}+���&f����T=���t���ҌF�L6���I�Z�������%�B0h�Ɯ~����^�gۓ��+�s0�ؿO����w|�t�;�1Һ�=���,c&k��_G]p���+`�ͯI,�_ CPW^����ޙ��SbF/S� oք'��g�1�+�]���Α�|d��Um󹖂�o���fv��=�a�F�����\,L�w��S�*�ߒ��|h�ٸ79S�"%CoEZ��&�Lf��q�]5&e�~� ��/b5���享��y�${|LOq��=�y������S_e�)���??�7@D��w<4vO���Y���GԭJ�sO�b0r_�UfZn�:vT��V�V�<7���!^�-�u!�}�a1>�i�FM���/g����}�`�Ԫ����g�~SA�z��9�e`RkT���@���+��B�7=�BSʼ^���g�+�Ne�AK�\,�*,i�nl��j[�)�b�������)�+���B��7������7�F���bg�'\y7�Iz��r#����4D%v+umA�ݢb�K�Ø��]���LI�Wv�8ޡ��c9޼lHS�Ê��]^��,r�lcy@�SVvr���좆H����EY���;��2w\��:c�|��߼��� w^���˕I����qm��|h��i�L�՝ʮ+�<:��3�/���ȦM���
����&��>�aљ��k�ջ��~�:pw����Q�/6+��x=�X���s����~�۹�M7Q���I�e�#��g��N�,�1K͞�4=����z��ι^�\S���Q�Sx�J�����L�B��+�ݥ)��h���:��]��.Īf!�P��q]Ie�G�O03�����{��]�8�}4K�M}���pM��9�-������&��1OM�j������]�Ä-����n�3�ʱ��E<z�@�'��۰eL�ԓkp^��)�cp���y�9�.��ͭ����K��&M�5_ w毮�̎~�f)Ȯ3�s�)珆�6�l��8��MF6&��Ka���1pX��L3����=����v���s���$�Z�n��ԫ�&ICU�yb�$�)�-M7�2�h�v��wؓ?i�}�s���{Ӵb�E)��Y���/g��!��d�c3Z[u����GsTؚ"�7������v�<�0�j_k㸱%G��H&��Eυ�Մu���WX(e�;d��n��N�O��w���6f���gv0�u��s�%�������r'��z2��#�O}�1�8��!�zx�ٳbm�~��o ;FZ�ےRQ9��������!���_}�ﰅ�F):N<���CD��)M'��p�:�!U,S�>X�i1\�AWr7����N���L�d�!�:v=5(����c령A	��u�g2w����k�"؞>�
 ��.�@ȇp�����X����rvF���߆w�vh˛�.�r��W^�^F^]k�(�%1.��ڥѬ`��y{�L������:%ognR�|m7p/(^�L$]pd��ڤ����P`MV�d*��`�� ߴS��,��9ݹ2�Q���5Ec�i�Z��t��@]lkw76T��}��8k����ø�&��ȸ�ۥ2-��w�p E�
]Ñ����tɘ��6=�kS�{��su�(����H�
�i1�F"^Y�ܽ��RR��M+=3:����3m�S��9��~k7˛���*�N��b�]�(�e
TWr-j��_��R�^�\I�k�k)�M��4G{މn�S�n�v�h��X��fn�Z�1�y�X�ǂ6%K����}/v�]ڥ�õ"�vѻD�gY��5�/]o΁����vZ74wJF�ܸ��)��v�|N�jS����W��N�0K5:��'ol�v	FoLЫ'9z���I.�TPA�)C�uC� }_®A_�z��9T�DTQ*��GSU�+�QTc,�y��\�>���
+���r����FV*����k3g4������U<�x��s��np���V̞��Z��e�U���l����DT%�Y�i�fa����Zb�h��RH ��*�'�MSNS�z�6p�WNUP�AQʹ&�C!
���A�FgL�J��"��ŅÚ�I)��Y�˅��Z�!QF�Re\�J�G��;J���jaE(���\�"��%�Q$ChI
a\(��EEÒg
"�.\�IUu5$�21(�@����������E�%p���뜂�B�:e�Y)�8]�VL��ʫ��W+�*� ���1	I�H�	����jDY��!�
�'$�'���ʮz����֔b�`���Rr�P�c�YU�J��}J���@�3&ny��c�o��,����7�]�g\$�C%ܩx��ׂR����;)\�b���s���TLw(���������8�5��T�u~1��Q��#ةB�+��g�b���fV��b��s�v�c]�����,���D���ġiy3]3�& J�UN5�^���U���S����,v!Tp㻲e����핂\`S�'�@�bz�z^�v�oۖv y`׮���C��؁y�4�V��8O+	S��/N�9JA��c�JD���"X���_d�	���)��x�!��w�:��݄�����0��o��zW�����<�Q���*0D�b�h�Bk�8I�_p��"_�ͼ������=t�#'�)����{U��J��Wu��|��Sc��I�k3���J�+0��ij���y	Η�X��4Wm�5��l�k�V��#�F�	�v����L/�y���|u^��3��l�kx;�*{����ޝ�4�p{��7�^��o ��Ay�'�9*���iv����?�|h~���
���C�a{�O�3*�^۹��{�������7)�q��^��}���#�{=	b2'�lm�T��Ța��19���}�;���p��8�O�����띹�t<�	�nw�	�&zz��tHd�8����ٯچ�!WR�3$�@S�s�n�K �W+�s9���#�7�<<T��ÚiT�wU�L��qq�*�޽JL�.=)�!Ö�,Q�w�-��{���}�|.�-��)D�o�LY�h*Ç�?<�E��7~F��>���E��LS
�-ȴ'��~>J�G����*��.#9�����E��f0b�%NY�;pe�i��<y��C8��~��GN��C�M�N��,�S�O�.�
p�(1g�>��ݷ/�)����d,�p ����`��\�ٽ:��&*è�L�ώR�.��[���9p4�Կ����	Փ�k����|���s��y&"k�D�W�Dz$�|$�e�{-v:����vț^u��G�&�74�o��V�C�C�mT��"�M�'����t`�+���R�e�����9�*�Ԍ��/
T���cW+5-�����3��4�)�G�H��`+�k�>��U�C��4����٫���̹8�&��@(��)�S�:1�Q�?m�U�%*#��Lw��}y9N���+P����2LY��^��x�Ô��P�����^�UF9���V��Y�?�K���߻O�<�Ce	��R3z���r��u�����Rw�U��8��|���4{�_�ޅ����FOz�#,BO��z�^�#T����K.S�C�����HM_�%�}���{�|Q��a����wF.�uG:@�']��*U�)w�8�7}OQ��d[�9�W�]�muix��2&z��k���(&"�γ�f��Qm[q�b������+F#�����깚J��<�o�yO�W���J�vz��U7B+}��%p��3��4����Q�Ň���
8!��ʛ�긚�!J.,=J,e��sFs��z��߃{�GVz�Ex��D�-�����R'��yΩ���n'D���C�(�\<.�C��ِֆ�<�.�K'���I�Gh��oհwɮ�9����Ui���)'�d8���q�>w�Y�G	��{f��:���g�ŋq��p���.�l�N�C�u0z^s���s���/9���S�R�ۯ#�Abs᧬!���F|j�r���5W	�kh�\���<�\���Vi�]wޘ��Օ�+J\u'�M�O�z�>���Ҝ�ܷ*f������1�xQ3<|x�q��}f0O�jQ���
�6,SwI�vІ�L��H�j��F~�yӵ���?/�ɾ�X����hY>� �#^S��� V���b��B�w]��xm�q>]�����j/��n�5˃S�Z��39�l�0.��~��@9}�mN���*���NY�y��dۣ��"��;����7�8&u�i�p�7���&h�goE:�B�M�ff���]<Va%v�n#G�[Ў����v�E��w����dj�"z���|V�{��&ອ�s/�(ӏk�[ٚ��+�׏�>����7G��*G�2��Ӟ��y�F+ji��C�N{�����Ss0g�`3���B�'������l& N��-x�2�Z����If���m�1����]z~~�	�k����R�7�e�ԑ�1�.DV�P+�%)��-O�ʃ=�X5�� �
�N�Q��@�~N&n+=��U���u��u������>�ְR�߭J�c*xW�~�^<��0لG�}�@��X}�'X��6\`S�dW�j&�
11^�z��J�X0ޜp�^�������.��=/���Fjw�c>n��˚>���@r���6��A��E�3��sɊ���R��x=I)�a��Ib��e��7�{�vr�f1;�1�J��kNyW)i�C���֗cL���s>r�p�<ح�B�oa9��Ưc��#��Q��ЌM_�s�/a��~{��׻���w>	WO1�*Z�������{� >�3�7�՛��L9�],9C]��*�y�xV�9��~�7'�<��Ԭ��qm�`�>b�>^;t�|�~��|q�|�/�_��'e�_��K�,"��o�1���z�Q�I��YY&����8*�jLzrl��=J���͇b<.בp){T��9:C��j+wa�/x��9:�9��Zz��Y�r��<����Cef	��]�$d�7*�˕��8��0�^tPk�]�,��9�|��VfG�]k#���w�e`�bz�"��ݜN��[����	� ��#���<�,��uW�P�=�7�R���êpT��r�o��9����>��y�7�����z,T�$3�h�~F�gknf������G����f��N��p����6
o�pL�f�X=CK��D��P^�=�k8������ ���y�Gi�noAW�Կ4X��y�_�]#*x�V4�ߏ(=F��J�$OEh��f�d�۔�{-������^�np�j���^���=NT�޳��h��E�r�u���.�}�0fC��٬2���V�V�F�)��gq�u5s��^gY�
=���DWAi���ZA~�-=?��N�c���vP��3�j=7	O�\j�wފ*#<��'�d΄�)��n����
0L�"_D1�c(O��d@�9+s)�Z�>��@���8�zRu1~!<�P̌r�JAX����BtoJ�����^��:�/�#�PU��c����n`��^�
�S����U�E�������{/.�N)��^xo?g)�Ƿ�Q��Gԕ�;��Hv9SG`2�eT�|*%r�6MW����8X�5�[
o��>\�����9{ٚ���#�1eʧ��[@�Nۨ�(r��m��ұb���%������ X�J��ˏV��+ﾪ��{+�]
��g��w���ˬs�+���s ��jY#����	�b5Q�^�����xuw�P�q�0d�yMd�y��~��$�B�d��
�z�����T3_���^����5f������:<9��g�ck�La�ڗ��'�T%�<̫�{n����6_��_�7�慨z{�̝,.��!����#"x����_h�E?�_�19�y^C���*4������q�`[˅�q�*Ç����;l�Ѝ�NNl�X�ؘaN�+d5��\yH�ƻ:�Ǡ�hM�@����;1���~SV��	ۀ�)��v�~��v�9�����oû�!���Z�{j��e�#6n�!>�"��>>�Y�ϸ�7-D�5)�5��6���_�9��uf�����#ϳM?\�9T���VDz�R����B�u��Xҗμ�E�ީ`�n�s�j��0:����JQ��Ʌ��J�dGMH��a�G��pp�	vص˱ԌǱ�.Y)�/au��Y�gս.5:P��R`��A?����s/3�����_/�u~.�鈡��`��B�$�5���}�j�ܦ�3����^�����s��J�u�z=�O�nM�͋�$+]�랱Ї����)K�Yі�^1E�݀
�u�������v�iɴ�c�I%c+fqv֪��m�t��&^�t^b�,�R�E�i�ͼ�K-���ni���  �|��z�8�BlY���}�t�*��L�я3��4� �dM�"�b�@5��oo<^������B��07/!�v�!�w�z�IRL�ͭ�7޸���`J�bq6S��tzz]b�^��|�NH�_~���U{�Ϯ��a���5�gN��D'�+�"s��{zag;1�e��h4&����u�<��*���bc��RL*�М�!@�ɭ`�P�{��@����P��F�S�5s4��	�~�y�>��x�~`��0�E:���'&=�����ʗ���|/���b�91jxl�c����j'C���cԢ��a��f��P�(Y�7E��f��ơw��=��dE�^�`o���?�ofyW)i�5B����?xy��L�X�^>ӵj�n5���B�9OrU�}^�ڬ��yں؇���F&���]�P�V���AI>�����'�����=�C��\?��s`+��#P��0<�}}Y��,[�h.؇�[����k}=~��v�/@�>���j�<�f��&g���®�E��OXC=z��SF�p��ɻ�p=��n
3G�o�du{���0M�=��Ϧ�̬���,���c�w����x���Y}��*�@n��cH����w�圼��W��3n�sD&�$#�R �`���9w�a�c�<e�����7�@rpV���M���`S��\[I����26#����������۞7���6����
�c��յ�?G`��1�.i�x����4U�noԷ�Q�ut�����Ϻu�c!�l��=�֣'յ<g�
b2=M�G`�!������R�u������p�L�޾����UX�?|f�,}��ה������|��	B�s�.J��ܩǾ��t���t#^��c���_ک��ϊ�r_��Js�j,td
���&�l��ʳ�N�32�o�֎�������T3>9��:<1��mM`�:�虠<�+=_:H���|4���ޯ���W��F_:���`�ہ+����%`9��T.RY���ۓ�Z���蟽��ұ~�i�tY�q�V��.��IST�KS��3Ǖ�eո)�~��)�2^�P�J�qz3���_���C�m���=2
�������t�rp.X$��Ǽ��xϬҘ:�HLAw�qAx�X��.8)�2LO�_q�a����;��5��/��:9�X���=�\ߗ�8���n�Xj�B�;�qt���`�?�6w��U�.}��/�~�۹�X�3]�;�Cx�q8���So\�%R��k�G�I������u�l�7��V�|��W����L���*����=�x+T���+mM����ƄF�9�;��G=���K7�������oT������J�����}���8��zMr����OxZ�A�^o�}�"/9Z3�N�F��ltc�|f�iDa�q�
p���q�Yz�̰��z%@ۭ��3w���Ƴс�6$`��(�����D��q���ZƟ�6���s����W(�I����]wN�w}a�/�68�}�Õ����"E�-�'��q,oь.9�
��5�)�^�l����aϗ��'_#|�릦�8׬Tz�[n#��D�!���	J�%��=��(z�r����^��*>ϝ+��R�µ�Fg�7�y!zyi��Q�9�<�B�UJ�
�ܽM�ע�'#t
��>��x�>�W�Az�L��U�A�k:{s�(А�)x}sE�;��n�2�p����[*�2���!��t�Z4�=�������Z�oX�0V�Ԡ�`9a8P�k��;�9m��W�Ե�b�W_��(�vH��z&�e��"�o��? ���W���8r��W�-p]�gڭ�������wa(��c�L��5��	��Q�o,���%�Ʊ@�ð����cǾO����?8�~��q������p۳�1�m��|k�IY��`8u�tj�M�<�GhɓnCWd���c[ݽ��j�7)�[��<�v
�%ܕ|��Jg�v�f=&&UU�I���Gu�`w�!^�\(ؠ��1���`3���'=X,`��<��N{(��N�x�=ѓ�s����|>U�#PW���~��fhǝ��	��;"ht� !=�OA���X1�:���c]xu��f�E�[�@�m���)��t����W� ��"�F/�y�z惫,�R7�^��K�xC˟?e�>ϼq�1�y7�l3y�^N�3�<�Q���8�DJ�b�aP;�����A��u�����p�%�Y�Wkҽ�q	�����{@�S��� ���p��襶z�����/� �g1�>�2nf�Ш[�>ˬS�]�����jy��Bp'A��\����U:�3[�@�P������Zg�5�P<ă���J���,�2��c@�Ӟ�lMǴ+��U�g(wغ����kC%���K>���n���5�5��(�[�u�{5Ḳ�����؊O��&�����o��ӿ.�!���bn�H�ul��eJχVD���x](�Se���Y��m�޳Zj;X��zl�[}�
�N7�V<~x1��=�u���/~#�Yھ\��~�\g:�S���!�7"�I!!�}�1��2�8J&���Ļ	�ٺݗ���4dn[�����U�h��c�tD����n�ӶeH��Y3��.o�)����ɷ0�����5�OkV�HaQѷ��X��f�u�h�s�����n?���5뫡�7�"o1|�4(�nΘ7 ��h�q6{Y[�7�%����d��3�D��rmm Tcq���Vܿ�?�/NK��B$�7����'u%�: 2��s7�<��l��5nz�Co�g���zݨ�!W�I��ƣ[��D��t��-�}���.�D���iW]��C���4�a�x�G�˹e����JQ��;{�Ϊ�����YƯ]9�o*􊽂�J�R�<�/,nϱ�b����'�*�]��rnӒ�QXu�6MHX�WZ��v�97�YH�%����Y3���O'��T ��z�חI����f�.,SNvGx�eU�`�e��9v�@~u��3�ljl��J/6�IOx." ���M©8%��`�蛏{��l���y{�����\k��E[��v�oNR�/����x�7F_'�+�R���;x�z�}Ӷ�{�mщe�[-�|��r�N�-�u�@�ow.y���s9�K�~�#�&�Ȅ��dV�G�����5��3�\��B�8N�Y��ܺ���v9��Uw4�a�ڻJ�e��[�1
���Ӕݗ�=����1g�^���X��Z<S��5��=ݪ�-���K����j� z���C}�M��Z�t�
��ĺ���������w��5ej�݋�>�1�
�p��v74���Rޙ�8h!іqIT�Xpn�hएΥ�]`������}�3�W>��%�r��|܇/�K�����:���=����V�I�����r�u���"��Nht3(�=|ڀ��+�6c�_j�o���<^��k"��l�D@������Z"�K��e�u�]�3Qq�u/*ۢK� ���_fL嘦���ҳ���Z!an�7y���E��h��T
�XW%���;�w���>�8��rn2qÞ.j:� d�&�m�7�5�8�ي�nÚES�������'l�ǺeΗ0�n��'�2!i��q��~ۥc-��i 1B�N}�lo1e�=C��㹘�F�#�,:޾�V`�6�iK�"86�a�¯=��HiƅK�Q,4��}�twg>܊Y}p�,ū�7���z3��EZfvR�r�������С7��E;x1[��Y{*CF�w��!���9�r�qh�<8�u��az�շX �q��ev���80���S5\{��kV{H��� \=���t�)]��lc�B��|;fa���r�C��E�4]�w�/�L���M�a:F}}��Lkg���ɃZ�&�JjL߽OU��.K�㤔e5�&�!U�f���em_j�ĩ�v.�/֮����<�PSN��$�,��ȼ��Vk�_5���N�
�ӕ�d�����f�w>�RfM&��2%dpA�U�B�� x���G*���+�}B�<2<�y盜��T�<+�S���gU�{��&f�Dy���I�	]�\�˨ R���(��r���*
*��ETz�$�!�)���r��k*�����D��
��8GU�Z	UY�U&Ur*ʔ�_X��Uף�U�����'��s�Q*���
����#0*�蹶r�YE2*#R.ʨ��DY��M;�U���E��:\-5���d�ʊ�Pw\̹��G��E~���
+�eVvP�Q�3"�&W(�#����(���AT\�Yt*B��Pr�� W��2N�̫β�n�Ql��r��W(�G��*��1*�T\%o<�t��C@�΄��W-H�E�T��E�����iUQe�+��Tp�)ZP�m��G��ir�u��$�ZP�BeD\��uy%؆@@�H$�$4'�({���}'�ԇ��[���$�^�e򜄳ݾU�Ռ��׭�gT�%>�O �U��(.z��$��Z��eQU�}_|>l�KęG/Z����S�$?MԴ'¤ ���(!g�>���vܿ5pܰf��V1X���'��;�i�*��F�R��@X5����fp�!E�z����X�����b�{�s����	�^���C��*|���2#��NED{�pY�3�,]��iu����ʋ}\����c�xnsUk��t�P�O��^B �����`��~|�_m�����ӏ&+�7�-�"ˎ�����hn�
x�q�����3������zD�?P�_h���t��ࣅ����z�8��N�^B:b����t(�3�'IN��5j0?m�
���sK~�kqem�c�-� �5���(Gˌ=��5��Ԟ8[�O����8Uه;�}⢉�-7�k�^ǜ�9��`����!�BxKS��ΞRna�_{�Lu�6�ᏡWք�r�Чu^�Cޫ�]$�|�1γ�\+a�0̑uZ�(�"�x��|���V	^;cح�z}����B"5\�����lPb�91ih����]X�O���� ���_�<>�������5�x�N=��W^����ﳝ����o<�?��|Q"}$���$�)��e[�D��q�qx�-t�f9���.��ǧ���в�1�A�1���57�ӽ�'�W}W6xL���ꊥ�>l xNi�ڔ��r�ms@�۪;g#3k{?����?���8�^_�9��=߃X�Gvfr���Y�e
�|�W�������B������^q�C:s�4��h��զ���̿��|}w��4�Dv��؆�[Bg�%{�\�6i���|���{�w*��.d���OM�����;���zo��-Ƿ��q�o��:�
�ܕ2 ��~�g��ގ�Μ�����=Vq,�s08G��P{�s�=aS�SFWN�����\7�^��[�=f�l�^oqa�ܬ���i8>~;A��'(D�G�v>�d�MQԵ�iw�Ϸ����fN��2�иG��8�߅w��zr����ATFŊn�;e�!�@5Ҧ=
����Ƌ�Ǖ���շ$*�r��3c>� �|�����C����������&��y���Q�r؇��ъus���U858
�r_��	Nqv|��
���;u�<����^G�����2�L �uMB2A�^Aߏ,1�<���~���q:&p9���<^�/Aq������?�f?]~��CG���7SJØ0��j�B�If��Í�&4>V�r�gԷ����ˏv:�#S�t���Oi����[�pS����v��F�iVZ�����o���x5�Qi���G����W/!��G��=�h)G{U�����7[���[m��,�y�W�s�k^Jj���%��u����l���jی�9�d��$�а�?�����%���{�qO�Wql�B��%�0(!%M��KS��3��^�� ���v�d��t���,���R�J���n��)�������AZ�^?��tG˫��t��6/�Ѡ�DTٶ'���a��8��Bl^��#%�|�Dȣ5C����z��/s�<�1m�u�?�����t$���7��3Bw�a��q�Q���;�{4��\�yF���[;�k�)j��!��,ete]/�ߠ�}����Ց�r�f0'~�!�U��F��5�A=p�t�<ٮcld�}��.د@������3o�;�Y���ؑ��bc~�"2ϣ�]V,�7���<i�K򽅞��%Aʒ��c����U��[C޹���i�=˟+ �1s/�$��#�Y/��. QΉ�Ggу�[R�hDO�:cEZ��&�Li������e�ϲ5��bgq�J�B;��mJ^V-R��{jϺ������c��M���������*��|}9��g:ه����Pc 5N�3NY�7�^���n�_�X���)�Gÿo�Iy�����~�]�ť֎ĖZ���g�ґr�X��� �R���={�#'*l6k=����2�L�0�Y)G�Q6�Ī��d��u:�5�Á7������ǹ��9��_|P>���r(zQ�q�C�!�73Cƣ`�����DZ�2f�Ç��Np�b�!��;����X�?4'�lb�l�~�~S��l�1��ǻt:7��j`С��z&R|r�
p.�pם�pӖ�ނ�a�~S@�]_*t3Z��#�B�C�;�7��D���O����B	���c��lZ�c����fj=W{�{t���r���e�M���q�;�6���f#8��ݒq��5jC���ٗ�f���Y����x[l)S��#Xe⁁�م��w�������@t�(OA�;�1!K��Q!Q�@�^�����9��G�Ұk���H!}0�9�%# gE�Q�exB�C6/��er�\3�u��	�/>Yq��M�Hf�Ҽ��gg����*0D��Lo?0�l���f�.���lm	�*m]�I��ܽ��Y�o�@�UZ�Į �p���n*���9��p�Dr�=G=�,�STK��>R��,"������Bo9XHM�v��bb��w�ݙ�d��,C~WQ¶|j�h�Z�+�I��� ��^�V�;���� D�}���]��U�]�y5�feA]�vʼ3�a��s;:9SB.yj�ws*?ϚǇ1m��h�z�����ep�1`gϺ���0�S9IR}�i&��*r�8I�3��ݽ���%YJ���������d��HY4=7}=�5D��w�>�|>
h#evIB4~HM���8߬1�,�,mvK���m'vuKD��N �rw�*�ů���)hœW���KzV�C2���o.60�a���!������Ȝo�6��h긚W���a�ڠ˸��4g���ǆ�J�f��.��p4Ÿ��a�O�Ź6�`�F��>���Dњ�d=M{ζ�Æ�����]�g�!9��v�O
p��5n^���%�c�{��Ic��^��J���ؙ����i��அNX!O�ݧ>�X�JQSW
;Y��-g��C��7;Fg���~+�ZdF�R�p��¨�X�p��!b�o Վg�bT�f!�u����](;2`1ݖatMA*G%D@��q�:��_�E88��\M*�tK�e�TL�/�<u#3���5V�1�҅��k�y�kg�G�>�C׫G��3v���=��(:�=��/@Y~�� \��)�����z1�&s��g S�&�P��2��7��+��N�x����럘�<��ݗ��ݨ�g��YF�N�IN���ը~ʈ0<v�/��=�T2��²�`�����8<�a���s)Q�BivQ�y���h>��u�8����],��l��4n������Gv�Ս!�n�t��{���(w�FsU�nG٭�����d�]����f�0�E��Mq��\��y�u9H���o�I��kVFjz��U}U���^�Sޫ��#���/���:�g쌝�W�,�'n��o�_��yo�B��/�"wA^@ٟt�C�ۈ��ֈ�V�D�M����t�|r���=�&:ƛjM�����5�9
��+�����˅l(�a���~��g�c�����O9{ٛ��×�G�<�|GiGX�o�����lN ؠ��Yɋ
xl�c����j'X�ǩC�(O�)�.kpl��¶,̊��:_Þ8Qǝ�Y^�c~���T��u僔�����[s-;��ft׃�u���8~�>�d�^��|�vIf�o";B�b��	�X��c�ӽQ�o2�J���mpj����m5c&h6(h�sc���г:z/�>���n=���>4/ޕ��f���௃����[�ow�}��d_*�FRx�k1�xU�~˛���>��0���="B�9��}�r8�z;e�U�=�����͞4W�R��?��"q��=�X�m�2�5�Q1U6A��bf��KuV��UV���c!cklmw��zr����&���:D��X�>���ׇ3��n׹^ϫ�:�1�7V�B��,%�&�_~a��mR�&�^��_�y��ea�G��] �M���4���r��������4�D�58F�KWʇs��9^��ѵ���]�xN��uG���)�y�j $�}y�Q�l����� ���u�B/�P�������H�8��U���~3c|���PX�-��dr��t��m�/��u�%�g�lWG���l[�\�T�5<Uk����S��$3y��\a�VLh��:M1��į��1�WE԰dX뫆gA�^Aߏ<1��mMg��:�rL��/�)��|3����:���gb�5�1@z�&BߠI31J7b̵��%����&!�W,4��w#���n��Q=��S���T��H��d8.!��EM��c���r��`<�k3�������c4�+������J5��ڬ1�Oh_��X�ACB��?����ߗ�o	�<�%���|��7��T�=������%�7!h�� =	Ņ�u�3�$l�A�K����o�`�������?ܭ?#
�G�1���_�X0���&o��bu�`���8��ԋ�j� ��ҊH`�9�޶�7ˌ����`!"���^[2�f�e��Yy�ј����i]G����'�
s#3[�%\a�����%��:�8�Y��U��םY���ؑ���(��Tr�\5�د^�֥��%���3!��zNu�jt���B	 ����P�^�3�]�K��MOS�ov���Y|n��R]=1oɕ]LO\>���#�I�5snܒ��;���.�����lǪ�܇��y"S������;�jg��:��7�wE�C<#�&�꯾���5��_����_�\s:��3e���Şξ��X�4?yO��=�[Cޱ5՝�5�>�k�@�_y�'ZzT��~�p�3��Q��g��_U�Jb�'���T��gxU6��x�L��Nwv�"#�j��úJT��%͹L>x1�P23�޿F��/>��MX�i˭�ʾc���8��t�lE�s�sY��1��8nt*�r�������'#w������)��M�꾱�s��v��c��[*R,WQ�\�g��/�<p���f�)����ڧ�U�ZhB���������%�L�0c���]JN����*|�TXӖ��U�ԱYꞩ�(��,�{�O�P�}�:��+����Q����?��P�t�h=�1B�p3���*��C/o�r����~;|��	�*����ީ���'��\�UN}f������b�cg_u�{�4u�\�}#t�@ϟ����J��9������@��O~:x�j)�>�J/�v-qS��ܰ��<�k��} �#l�r��+t��gE�Q�eyP��;��7n3��{���]����(˿��D�,uC�m�ļZ�J�B�l����V��i��?.��T���ߓ�ޛlV��<� x�HK�RMT��z��O(�`瘝�ښ�+ʄ�ܭJ��p�Y��.�;���#�qwN��/�������zq�fs��[�'&#����%	��y�"p�� �&�-�����b�Byp�>f��N��L+k�ݘS�����>�B��q���X���E��ld��ټ.�_��@*iL%Q�b��z�.���W���#�]�_�3��;9CX������*|+�o.�ϠOet4��}:�ߞ�ܬߌ<���y�v��7���X��`�3>����9i��k�1 �+~:���"s���ߞ}���l�X���ߵ�����p�,)-���K>���^4:;k����``��N��۳|��5��ݵ���#���-u1>~�Zx���7�6�*V���1S�gO�\�Ն�)��N,R�fc>�}��\(�1n=�Xpߝ�r~�{�7�0�v�c�x1���MϞl�3>���,9��>����}�!��i�p�M[��ۀ�=�+�9��lz��mW��p��3}K�g� `hg���j��ud�'�A8���}Ʃ�uQ=1�y�hs������G.���Sp�ͬp(.w����hZ`��x�rؾ��L�OW��c�]��Ī��D�B�w�X���S=���R�&�r路�o�_1x�X9�AK໽E��]��T7�˥�Ӥ��*��a��z2�shw���*��2�����DnG1���!k��Ժ����y�N�`�Zh�X�:��U�����Y�\k�����-dO�%LO��g�]X��ߊ�j_��B��*G%F	�0#!�1�Q��F��*�w~7n�\�F���8]j�b�}r��Z�ƀ�(Xͪ��\�]"{D
���WN��JM�����Ք/�h\���T���2�q�&s�c�4Ω�u����%�=�2�X��`m����/�`켎f�FC.�tfw��%;s��;*e�"zhZE���z(͸�`*�lu�?0hM1�ʜ0e�T�O���R��J�{{=��tƼ�%N{�A>_��n�0#��*�
�T"$�M}��ΞRna��P����ꀴ3��'��iLk%?��ք�HP>Jo�¶g�EL+�e�P0p�)�ǞRt�u�*jx_��\���9�)�Ow��	�cݞ���
���lPb�R3��E��[���¼ś���4�{κ/R��u�0�u��v�oN�r�
3�<���z���c��R&�����[$���ׯ��p�����Φ���`���d�]�S��]�Y���'l.�!�~�@Q���2�$!b�![��u{�a�7�)P�y{�}y1��Q|#��3:xvs�1=c�)��z��َ������4��E�N!��VM�uO.�U��u�#���FKu�qn�y��K�G,q�E빧���+���`!LƎL?	��]k�t��ٮ�3�T��ѻ�]J�*H�D?�t
�Dոo��ؘa��*�zo]ɖ�m��6`�o��;�*��sL�ߺ���*\��i]2ۼ��;�җK���V���bMFSr��no�y�s�/��zh�G�ˬN���j��;7/�(?1��hJ<��ݽ����=fc�F�	P�h	��,��6�Fz��!Yk�j���q��nYA����)
�<Tl���M#n�PN�e�^J{A�n�o�OBv4F߇Ec%���Z.n]8&l��t�X�k����s}�8j���z9�=��{�"\V��\c9wwâl�T�=sQ��Z���GNn�N��Z��c=�=�ak_�f�tV�a �G*���-p��k._\��*�ږ*u㺒Y���Y��gr�/���q�!6��$Z���G���$\3��{��h�Gv0��z�Mi�ɳz��=#]�C�)�|���?U��#&��r��J}z�ϘC7�u����q�\����>������;,G��B+�
�3�ws��ZH�,D�y�`8��U�h�r$VO�����n,�`��+�SqGH*�X�t�L�ɦ�\;�Fḱ�t\��n��L!5�����V�0XQ�Wy{˜e{����Ѿj7�i���ǔc��=���a�s���둲wk��]'O��u�4��)̾Z���P��ea�X��:��,\��\_h�a�[� �UL���]�,�ě�C�7�Q�P�c9P9Sw�.��r륋�{�����d"��R�����VL�-��;N�!�nn�B���sf+�Zh��g{o�{�E�Q�Ĥ�w ��6e��W*x�;(Q8�a���<=�������22A�EF72n���㻣��I�%n��䗘wi����D]Lzw$�!P�(;�g"�S�]T�9�׊��C^�_T�ߺ-�]�d�Yx2&�A{�>خ��.6���tD"�	�s�N�Ի�U+�D��0�6ۻ�rvn.������k���}�o~A��=[3~�:��7��+�j�]-���Sj��KS���d���s��؍͝��o<�D�E����V�.Z��u�)oI���~�L��߯ڴ+�7���HZ�^��>�u�){E>qx��$�C��"��h�|�KLM���n��P����,'���/l���f*�Φ�3b�j�2jG��6o�����|_��W�y�oz��6&c=�pϲ�Y�U�G��V{d�qe����v�8�ޜ�%���ٞ��t��Xח�g\C��z9���}ť�S���U���y7�/#ِEw�:���UɅN(Ve*مs�z/�
���9TETr�y<��"$���#�SN���"�\��'.�D�`T�%:j�$�B��8\�D�J��������sԭ�<���4@�U�TzŸ���rS�p���5'>C��"_v;
�E9���qA)�W���WGt�]g�Ի|��r�DE�uYr�\�G�V.8�UEE\�0/<�W)Շ�a蟺ܨ�
���yЙ�'"#�\��2� ��	�E	$�*�:�9FIPQWL�Dv��R'�~�"9w��C����TAp ��w���	��J�EÔC�YL<��^�ް��EEr���K�����ȭeˎK���T�%�s3�P��O�ˑå�[��{Dj��ٮ޲ku���"�5�λ�sP{-]lQ�A��G����6��x��C�^�	�(&2k�ƫ����eyO��^2i���6h�$�,��P�?W��#޿�kϯ��[�iv�8U�Eu�D��lo�K;��k��#�U�Z�OʿZğ�1�\������[������zkkb^�5$d�Q�Zn�5n2g�;r����V�/I�����n}�/5�1�u�o�Ǧ�xi�e��Rܩ�r�;X�c~�����mKύ}ALF��+��?w���^����1��b���ԋ��<n|���f(_'�`�k�r}_OlY�e���>�=>���,O�J�u�x���+�Td8�
�r_�l%89��}�)zx(��n�P��~��W@���>�9��r�>3�f��y���mM?P�w9��b���n3R}-TW,l�����cMtL��$��SJ7b̺T.�loE�(��������t���`"�l�㟟�BsU$N��A_�?��h��ʻ*�d�+���r&�t��iLM�a:��8!WC�ߊ7�v�j��)���0o�2
��q_���5�kă當�?U�z���.�g���Y���YgJ�,m��7Õz�H�k�˟� ���M�_�௓����)�	����C�#�ٽ.�
7*1�3�Q׼6�l�kv�Ht�ٛg��xX�(J�U���q[څH�W�c2s�d^����|>:��Ez4�ȿO�eC��X�|��D5y�N,.NmG$l�ϔ�&'�Uu���{>�Xr8#\�>��ҍ�0ߺ�����3Bw�a��p��HK�j���Os��*q�q���=���i����ʕ>��N�{ex7�o�dE��h�`N�G!El�*�勛���琁�N���q�s�7�O�D�~��$�xC��|������u�ڽ�"�:�Nu<}f&�9�~�C=��s����}0�͖}�Q^\b[c�2`~�ַ� >���F5V���uO<�E".s|��0��WSp�	3~��Ggў�ڞ,ބD��չJ�;����3��M��^��f�����&��qꔧ�S�K�r�Ϟt�@��z���ڗ�^��M[����b�W�\���{�a=F'�ȱ�1g֠��e�r�i�)X��������=΃�������r��EY�����E����t�<�0�X��/�<p��p����q��n�Ex��4�d>Gb���~3�g�5�z�0�z.�'>9a8���^wQ�鹸��􌤯���¤ԍM��j�1O�ϗf�T�Nva���Q�6���{,]�̸P��$���DƱd��J�75"r�G����i+��\�|$sLca��y�d�����ݛ/�l�ݒȂ���K�;��5�s�&�K�yzA�6s�5�}��}Eg/9������h������0m}��J���~,,x!�S�B	���c��g�b��]+;%Gg���:L���/R�/m�9�7j]u��i���� ��!x�lx����9���6��{cm_:���1���U��7J�z�h|�Gf�΁a����"zB=�|F]s�>��_�85�]����z��H:!ft'INƋt�*謎�)�2����1�����3��Hd��D�aQ��/��츇�<q@1�ɼ3W�����v|˅Ǻ+�mgH���=���0i�����V:������)������}�q��70o�/b�TҘ�|�)���=Ә�;�3��}+[gþ�0��+�ƨ�1'�>R�c�@�]��ׇ��r"O'�sB�ػ'���!6ҰX��17Qk�l<�f�gP��B�1Z�^_����$��;����{:��������R�����b�0���04�豵�.NT�7�xR����0p��LycJ�!����{7�pݳ��.60qvJ�b����]"HޘD�鯈��
"���+����<h�7�8���(D��Ӳl�p�� [>K�x�O*]5��7{�/ouJ��,�C��tW�<NK���
�*b*�9}��Hܬ+Y�Q����ݏU��ITQ^�Ѽ�kk.��x띺F����Ōr�T�[7������G��V�;��`ǅOF�^�nc9�Cz/��Fb�{~*Æ��[�l��巜)t��&�^�"�g���f����V��L���h60������Fb܉Z���c�z�Weq��\��x�����?P���f*��q>Uk��b�׼Q�|���A��g��ʯ<�R/��Q�*�z_�ܙ ��3�t��r��j�%�!J�?*B�Ȝ��G�t_�����q��nvr�W��*��X���^[R�f�>9Pp*9*3�0#"�u���i~G��G��a�~ �ucrÇ�.�Zc��y����ɍ�:P��mT���\�]"{6�Gݛz���->�p& M�D�*;��KK/�.^��S�S��w�g�i�����a��)�{۾Jcw�H�,БCE(�?d�}'>켎zb����t�>��˚rUM�o�	�Vg�WC�ۈx�`KP(H���T��1���1��񽇿Rx�v�N�f�����g�d���T�U�~�	ݘ���B��DL+�P��	�����~Z:����>��Ąb`��d�n�~P��Y�!�>����{��_�uPb3x���sɽT{����m�.]2h�Zb�!+�XF��s,ZۜH9�j���F
�r��Qf����D�<���у�䜒��n����{�=��Jdl���|��~K�'$���|��[&��c<�)L�x3�s�M�~b`�޿ߤ�~��	HH;�*Ϭ.�����s�?�hY��}���|9:�{*ǭ�}8}�=/��岬J@{�����oe���i�#%���Rԝbi���\�W�M�ӵ��z�m�2�a��5�:��(�ǞD^/[������j�H�޽r��ڰ�׽�;�r��垚���vg���Tɖ��U?NU�%�w�	ϱ�	ml�
My����M�#��O������V�s�Yb���?Ӱ�΀߾�����n<���\N���\z��:�FCf�ʳ[�5���g6_ʅ�I���2`p�c,{�Wc{��3��{�}G_kǞ/Y��)]g��~�SF|U\5:w��[X�v��>�3�-AJ҃�������wՙ���o�;@�蠃֔�5V��/y��X���F8O�j^q���u�Xv}A���y����+:�;Z�u�k��E�8���)��61c�0b5�<2�t�J6�ߵ]�}&���Ҿ�@z���1�;,�8_��\�����~!V�O�9���@�ŧ�}s
�׳;T?@�)s�!fk�&�־f�Ψ�Ng�j�B��7Ne���{(�2od�(wQ��E���@r��}�3��+`�n�������ꪶԹn�T�g�����nM�Ƅ�kSA����r����O�Qt��Έ�y̶,l�cܯ�������}(��� QT$�zP(�K(uR�3�� ��7|���ts���sk�Uy�G��\��Ss���+=C�I�J!�c�]�4|��9���c!c��T=@�ͩ6/�����ǘjʓ�|�l�w�ʨ�t��Gv��Cฆ>�P4u{�sx�i�W�'�:�_P\T��+�4����,7��}�_��/��6g�V)Ж���;p�"�/uC�C�Q�ʜ�R�T98,pycr�^@{�N,.��c�6\g�t@�>��¬�H7���#���@��j	|���v������]&��{
����:��k5��+��љ�Is�^򖞠�X3���S�^�ӧ��q��}�"/9Z3��F���Ym(�8�т��_�=d�d��3�
����GrϾRS�:�K9�(���P����ݔH��!!�DC�oք`M_�p{e�W�b��$ŏ���X6=�dzY�Z��d���c�Jo8K�=S-��`L�D�Tkk�읩^B!�"����Y>���%NU�X���9瓣ۃf�W��cu�ͼ��
�Gnʓ���ߗ�Q��y� ��4�_��K��. �'8t9]���n;T;p�o��&�H������Ѫ:I�uq2L;�De� ���쾍gu�CnAd'Z#�ʚŉ[5lB�G�� P�w{���>�����5�����g�����}%͹o�ŪV`\?�z��*^�v��򙈻Y�z�o�"[��Q*y�{j`�}j`5N�UV��M�׶�97ͫ�^��{k���Υ�ʋ�vz��!�|�vD~~��8۷���<����f�S�`�==��S�X[,x���~S�>٨��P����'�)��.�5�õ��I����DSFm�^�r�c�=�����)�+�����G�_�W 5��^�7a��Ȧ�y�bh��<p3�fj1{m��	څ�v2 c�$ObX��aǲ{��*w:�~z}ry���zk&ԧ�,��%Z���@��f[���w�a��=S����	q	evW��iB�.?�p��v��4� �Fٝ�:Jv7�t���c_�d�b�77YOi犙��bg^P��~����+;.!�P`�o�!��J�	��u^�>�Q���~=X���f}ΣѦFz_�tD�V.f�T&�?Ź7`ڄ���7�=3쯈��m�e+巑�n���j�cV�(T1(�Ґ�m@%����طml�r���n
�<I'2;8����m���$�s��=����䟴Ayy�VǤ��~��K����]�1�X�d�b2<�P��K��Ң�ӷkH2Ʋ��n�4����.��<}~^��>�i���t7d^E&������͕|�^���s����u����sW�j�x|�B��3�.:���v�CY�������ev����|&��6��#�7Qk�l<5{5�Do�
��:�u�����n�3�ZGK�=8k)b�����3�{��7�����E���/��ڗ��&�2|�j�v�b�f��bqȰ���r�v�j�}���}:�������[�dO�Y#Զ�N��b��3Fz�Ԧ�"hxR�G�K��P�1ʺW�p���xa����f�:��V��7w�f��4��{��Xe&n��~V|C�+��쟾uф1n��I��u��;��nw��>]Ӭv�8�i�ݮ�zs���s����U���ts�Ex�ڠ��y�u��C�<;�L������2������ ��$֙�T�Ä�P��#�T�3<F�D��Yd彃x���B5���}����9p7��ڗ��B|n����ɑ4$NC�\)�f���C���D(���,8K�Ů]��f|�����\�NT$�Rc��?::;I¨W�_����ү[�s�=W^�>��u�EL�og�:�ɜ>u��"�$u�u�,�v�Y͐�.
mhެ<�TT��)���N�h�x�wdW���N6�G�Ԑ���Z��iA"��38���u�J��5��3)�Ky,��moR�叺d	q��+#կ�}��jW���he������	Q迩��8;/�e��\��ONk�eތx	����eLhi�t�s�}�G�o�0�\���XC�qX#�������t�>���(�2�6��y��G���t�)zr���l��TA�[U�bI��QS�:�fFN�ޖ}��Ŀ�3s��o�R����i��~J��IUF;���B��DL+T"$�Bk�5>���S^M�V`�qT�?9�>�s-\:�>�0�i���_Z�
��U�Z�[&�S
�\�1*X�&k��!�o=�{�f��W�T�r�e?|
�*��g�<�*[�6(1`rb?X꯲����-��ƯVE����3w�bP��S�˭��~�[ӫ�r�
3�<���p��`c�R'[�F��U�Nr'���/2i���3)�~0χ�ƞ<�����r��,���#�.�!���3������q}!��}��/�b�O��J�,��)�'�F�΀ދ�Ͻ�̺��y�D^�z�H���aBkun]�l�o�6sf��y,c ���X�����J��;�yT�e簱�o��jD�U�%F_UB޷ݻX��z_
�����%�,oo0�l��� �G�����y�*J��{l��'5��#1�pT�Gu�ؖu@���8��F�b�;�I��B�sNw5�w3�$"ӥ������� :�x��!���������r3�]\5:�����8�]��`3�.ld��XT�rf'���p���z�Af�"��4`5蠇[S��[���U[�^�v2|���w��zr���:3�ZkN�gw������u�b�����ȇ��`;^�R/�<n}��)�61c�1pby͓SYB������~�K�����!_W��dvvYOVũ��FÎs���%�X5�*�؉�ߢ0�Tf�'���a�P��7�*�6$؁^����]JE��W��sאt��ؐS�.Te��d����6:�'D�9���ϕd�Q���L
��$͊�rV��Z��'��ў���k�ĸ&�P_¹���ܭ91����X����T��k���D��\C�JX]���0gůlY&����P�v1���pS��=��s~�Xc�����S�5=�����h{��83�b�X�ӎrna�+�	>V܄���qav'X��6\Ww�X*dNV҇��b���<+}C�2���,��ǯ-t��a��L��^X�7��\�tO�~ �C��0`|+k~G�:1V�����fh��]�d�@,ӕ���Z\�2V���{�n��䄗M�Ӽ�t�qׂ���T4�%����xL{�$�%�<{6_�0e�����"�6FDt�#h�x&W�q
���pjPZn���W5�ǧ)��%��;�7)�hy9�֠ܠNa��`vS�x@�^�Ѕ�n��S�է\�\�]8�pD�:���2��0��4s�y�ִ0o�ǃI!6A/�}��ݡ�n��4�o��>a����VP����o�ДN��(4�i��e�k��H�p3GYj�6�N�:N����{	q����]�
��F9�vm��k�EƎ���]W )2�6�l�s�֊� ��w��lq��I9�s罻��qX��r�P%s/_6�.d+�r������k��6m_�J�]6kxt�Ճ�h$���%jM�s��;X��;��ݚf�oi���9P�oK�T�ҩ��)�s�IqYιq��A�n�x�A�&]wO��Yӗ�qgv��Cx�بW;} [�+W,��6��S��7����`wt��noq�*���[�zn�,�Am��}"}�t�Q�p����!�%�j�q!j(�����L���	Z���@��C�sނ�1Ϡ뫦+=[ʱ;�5y�d��U/tu�z,�޳d5�[�`����6z�4	67W���C�roO��p&�Vv�2d���V7hIz)�cd����{�eYθ��o�/��M����oˀ���W��������#U��]ղ�J�4r���Qש쓺Y�ߖ�髼U�m��T���?�`A#Ql�gx"�Ih����1���v�.sMk�N}N�J�K�iL�\���Ia��v�2���xwoy�h�=˚\�'=��U@{��ٗK����}2�'����r� Ҏx���i�[\Z�$�.�a�{||��!	���zVP#��-�
���n��v�Y��9
O�ھ�]Ս�g����l�ς�u����P���6`\��[Ľuҳc;�[�u�t�AE���U�d�lt�i�	g�G��f���NRE�Y��LӨ��{�Oe��,ڜN-��>���*��A���+&�U�f�5��q`��*[�����m�#��ӱTz�@���|�A,�9�q�KU����1��hm-��v$$�u6$�̢�M�@�)�p�GM����91{#!�wޤ[��/*�ej1��[�z�g,����X��"��OSwV:<���_ء��xv����W+�d)gu�G�L
�E뾛(X�Ov���f�5��|f���j�*��v��ǊW�/Jo��0�7+����՜Xb�<������#9�D�E��m��p�f�x@6�sK,i�o3N��f��&|���^�Yhvo<�79[}�}�st�z�B�o���!����TGd��77��Cs���bڍ�a.�W;hf��\�t0���agW�Nɋ&���������.[�^˺烠��3yK�����LV���r<��z6;�O��+.�E���?�GԮV�z2G�"r�9%���+�~NL�iETA��IU��^E��W��BeDf���E���"��j}�׬\��w�u#"�S�qʎ���5��U�(�D>�}��^c�N���*�BL3�}�w�'�9_P/ZZ蹎t�����j�{�u����11,H�������z�\�:�;�q����Вy�(���TG�ۺ�O�+�**��s�d�z�_U'"�tO��E��È�n��^��x9�u��z��O'���'�Uw�sz��t"��EDJ ������:>y<�좽B���Er��Uz�w��Ե�Ҫ�E֙Ҫ.�i\����i�Q�Z,%�{��L�C���nyWo'��B�7}�>F;�Mq�{�P�󺴒|�yq��/Z��G��̪,**�9%�O%Ε
,�r
1՗�<��ⰼ�D�����˕Qy�PjEUf1IMF����P���Ք����=��]gU���n�<^`פs��Ϲ�2Y�p�ۗ�Lw��<TnY}��LG#NǊ^���򾯪��w�z��`ަ��
�;�CT��C`�|Fh��T��/d釭}������ʓ���l����5���F|Z��g��qt�ٰRO�����GrϾRS�;y����'�Z߳��]��&^{�{[BF/S�~�#j����y���*�70F3F��,�Zo�7����g�dQw��fm�f�4Þ�]L9��B2'9�8���0{+jV��Ǡ�.�[x��^�����p�-�b��"Wl�����z�)3,C����|�c�o��[xʕ�m4;�wQ7~��6�5���y�	�?y��ǎ�~-Ϊ�r�7�_.��NlM���Z�.y,���JC<��D�v_������^�B�HC�}s!ʪ=�x��=у��ߖ�x����=�9��p$V���N �ZdA�c�ȼ,5���|>_b���Jk6�	��Q9��M�]C]��ޕ{K�S@ŏ3;��7��ę�$O����ةB	�B����OX���W�(Es�ϟ��1�]�gڭ�����7�����}�ȟ��H���(Xt�W=R����+�8mЙ?��s[�v�>�(�}�[���|�^�Z�
g���O{�L��w�YȬ���F�3�o����������2�[�����D7y�I�e�~�H�X��)���&7����[6�o&n��XF�R_cj������G����|�^�p�P��P�&r�c��f�բU���S����za�a�+AT�B�8}��{����De�!���b�Qb��X1�y`׮�􃰍�:�%;n��y�Uw^�[TO���I�!��2lu��L�F$G9�}�q�����C7��b#���pڌ�A>q��Q�hп*�X+�iW�0���E��`ڄ�����
�d�����g�Ԧ��թ�J�� *��
�X�Sc��k�>bhY�ʎ���S�Q\"4O���}s�XoǼ�'&�jy��Bp'A��ь��Q��Zg��	X>b.9�a�������+�ܯ{E~;���mҙ�O�[pW��8߬0ҿ�'�.:�*^5E�<7.�TQ���o�İ�(4J�>��٦~|7lƭ��.68��@]LC�����FD��x����{��yb��*�l5�P����Á���br5��}�P��1n=��vLʇ��kn_�I '7�w�1����������y^�gE�"ПTHl{�}�!����LV��.">X�c,��.:�\Pڐ����pص�)]t�A�lW4���B�19!�ﷇr�L
Ole���O�K��|\9��$ͼ���	����fo2�o;C3M[�`��GbM����{�Y�����K����1W"�=[5�A�]���v���k��B��$ѓ(��c?���/_�zx�~��.���@j�Oʅ�I��)��x,��y?o�����f�����ס�M��]�/�j�~�d&ղ��9]��CB�Ȝ��x1�
�V�c�{���+%��b|z,[��u:fܸ�3+�n|r��TrTdȎ�&C�Nf���[�������HS���{-]��f��T�:P��U&���nODg�a��${b���ȗ��������є�t��/�����g�T��D˿r�ح�n��=X�x�*�ꡮqNȚ�H���\_@��w��9�9�6�ǽ�}�8�P��9ƻc�,$���ʒ���j�?eD����� D�s	�>�F�/pU����&b&�yq��$|f$�5�\���z,��U�l�Wfʈ\h��*T&�
jV��.�ӳ�e\zc7��/ѥ��z_ݕ^u���6ԝ�_Z�$(g�V}ap��tT¿���WQ�S�r�6�'Ս�`!�ŞS��-�bR�g�;���lN6(1e��������ތ�x���r����BQ�M(���
Mc�H�(��/eϞ��ȱ'��}�m۽��6�S���,r�/��㐡��W�2ug���w�Fsn��w�&�o$��[/@�g58+r��(;�m�M�.�c\�=v�\�m�h��ю��%�5~�3�)w__��	��or�]�����+�����Tv}���z���q�q@^�`o�[��we�3��i��k���F��z_�>2�9J_h���2�~�^���Ϗ��1��#�o���T_�sv\"`���bB1�������AVl�*Z~��ROl|�/��N�x�A�7��e�lwy:�"�7�����U�3[�s��|�o�b�?�K<<�A�ؤ<̛�_�G��90<#��.��b;X�Ϻ��X��a�ϋ���Gɻ�{mc��*���ό�KPR��������]��=Z�3ߛ����/���%<U�n|��/G;klOm�\اqu��ܱz�|d��/�6�}"������#��ȇ��0�:������Uc��f�/G�]o��w�!2v,�WCu�8'������L!_P�8�DG_ýf1N�wQz����]�G�\Z���{��x�$���nl'89��}���t<#�G� k��M�r�V����b�C�K7R����μ</W~q�������s�'DˏL�73>���H+�Lة�%H��x�y�K�M@�c8��[�T��+�>�ޚ���y�=�����A����Y�G[��g���M.�1���Γ��/y PV�J��쇛}-�w�fh뾮�Zm5wN�k�.�NეGy�l�̈c�y����v�sULmk*#_�U|�2�w��U:+�������+67�7=����h�S˸�t��Gxu@��	03���Q���J39�epJ劘�=8r�!GB9�^����t>�(���j��)����v~�=#i��j�����^O8�\K)A��ӎ2na���byycr�W��bu�='鼪7~xvw=���`�>�����i�Q1C�R�U��\r����	3~^X�5;�0=lN#ê��w����$�p�Q���ˋ���B��я�8���:z���o�~g�f^�C7ٯ$��q�V\�7~�#J�,l�k�of�P���|ğ��w,���~��:9I��ߞv�����^���Č�z����k�}0�6Y�!Eyg*I�1�>R�9pb�=kƱ!���w�`/��^��͌i�=��(?P�X9�8���YN��Y�Pk�ٙ��3ww���'�|9����;
�G/���5��~ڬ��/_<�[�"y�,_�9CՇo�=]�u����v��o
p=?�?Bn�m�w�`�>�0�ʙ�.c�̩��ꋕ� �1X"��pP�G�G0����݆�t�A���Ύ-�����.yx��nA�Ō%�I�h�W2j|��e��G�_R��Z���_\�¤s$�����������Zw7۹��(�IV�[�f����HTz4����V.�|
~�L��w�g��]~�`��)`7�����z,T�$_]!�����]A���4��ZֆG���=H�R��s1���f�)����Q�)�3횁|=B�b�R���, �<V��}�:�`��"�y��i7PƬ���{K�S@���b�.�3}TbL��F$3>����^�ŝ~ �^��X�����5[3Q�/m�9�;P��ʀ�fb0��Ӓ���˵�(�}]���C���'r�0���a��g�j�V�F�)��h��w���pOGT|�.D�~�\b7yd�w"`�	0bB�����z��H;�3��S��މk���p-��i@ٟ
9�H`j�n0)�2�P�D�Lu'�Vv\C��� �y7�
�^�Q��F�{VUv%S�=�)�]�gbyp��/ʇ��_|�J��Lh~!�nM�ٹq�]k�*i�fP�s�#�'�?��8�S��NwQap�����_(5D���M>^����g=�Ŧ��p����g 1^�p߇���&�9XHJr�h�E��.M^�B��"=�7��_'�1���a���Έ�Ԛ��o�E[ͺwսfW�se;���t�%�
���;V�p�� ��8��9J}�6����+�F�Ek��=���!�=�c���:�|��Ԩv�f�4vғ�V��>��X��'�C����gk�&�oF��͚}ޙ���}�{�師�~��i�c/���ו�;�H�}���`^�����Ϣ��%�\{(c����sE���3ҍ�ԧ�ϕct)U��O[<���v��uk;}g��ӫ��x��b�t�z��+E��.�s~���ޔ��}0�.:kuB�����#�����o��y�g���ZE��ϭx���/�Y��tc�r���r7�T&5i�6Q����'�*&=�]���T�lm*D;��2bgm�9�1j�չz��SO�Q�zx��Ӝ>I��b�{�f�[��s�].��=3��b�����_����5pܿA������Mi��N�Ӝ�=����tx'��=�0o���Id<[������S�JTr�FW�3Y��X5�bY�+�>�"�ެ�\�o������y��6(�Ö,]��u#�� �Z��r�f�罫öv����> �WRc�4����C��!|t����jW��>��(��v�S�S�0�슄����y���)zv����~��qNȚ���(�_�>�ò�9�1FÁ�Cs]�7�B�|���>JZv�$���鹵�Ɯ�Ϣ6��q~�P��.�{/�k�*����J }-����&����XHapw-!�;��n�H���;���o֗����@�x��`e��2o��G���Ths4`�>�n��'X��Z�N�����Y����EDg���?�vL�N���߱�Q��n ⭁*±2%�*}S.)wwza6NԳ����K>W����D:9>j���]��;q>U�&�B"HT$�xI�7�^{�ϸ�:Dx%���})ϾYP�{�Lwi���?R��ڂU�.���詅��t�Y��[K/��^�w�fZ�(h��_�yɹ�-�%�vz�©�8�YɊ>���̡��Mj�����c'�3u:�WA�qqa�R�˭��ΜG�8Qǝ�Y�z�ʪ{��ǣ+'u��P�|�����U�ZgK*���"|<�c�yo��UOӕ~��v_�Q�^c׼�p����&��߯�`Mv	�u����<�)'�,X^�A�'���������:*5�՘���w���|R�{⭈q���[no�j�����6���N&�ޘ���t1z]�B�����Wsh�w�r�K��գABsWX#����FQw���&�!�V���O���s���/�S[;QcӞ'�V��s=ix��I���>#ݑA�ZS��[��Lӗ�B�����6�}�)ܺ�hS�X0^Ά;ᜫ�d�=&V=ӳ��o�b=p==F�D�!_���G����@�w��@���1��I��Jl�T�ˆL�[��0/S�+wTX�f��W,BJHk�}�c9�An=�'o"�x�����{��c7-9 ���Sq������u�!�׆���t�J��#�##�'q��ȇ��`5�u#��jX
�����^:��Gj,M�3�U>�����(
1��W��N�a��҅8�DG_z�b�Ϊ-�p�����'����7�A���t���Js����ѡ;���*P2/��h\Q��[���Zw(d~���xcty�SX���s�;Jtl�g`⬙�=4�I�lA]�B>K�/}~�z��⦼�0c��Z���RY��8�rc_+[9�����G�rf#����Q�hǵ߫��4� 6'�A����A�<�c.��!OC�To��Xc>S�'�~�G�^��z)��cPf3�9�c*1�*'>)B���G)ӕN|�`��X܅��������y�*���J��1���VVr�_Zk����sB��O�~��f{�,ox��>^V����L\.�=�{Ư�ٱ�fBY0�e�(*KA�r�S{4�u���D��&4e�/�o�vU=�C���{tގ���:�Y��ev��z�"/Fc�C��u��KO��)&0|ă��*�Dl��_}�eH�>v_�q��o�7�
�*t��Y
��'�ye�;���}	�d���V.�I�O�'�V�Aչ^>��U�P�u�d謵t�۾r���1�^�^�fD6b1���\�����Rz�����(���"�Z�'it���N�����ﾴϙ��;ٟ�g�����;|�=�� �S���j���g؅��$Q�|�����U��^حsj�v���}Y��q��j�a�?P�X9�8�D�3��Ǜ��k�h�^I��mװ\�3��[F{�]���%J�ꇯ�Nq���7x����o%X͉�Hm�6����h�$�n�g��Ӈ�v=ۧ\qe"��]���XC�-��փ�}d��5�k}�d�����J[k���E.=����\=�0ǡ`tJ��Vv�ೲ�ov(�B6�/�j�|��n��2�2@�1�Y���7W|��{�#xy-���N�Wmb�����jfl-��d�>��>�1M����{x�}0T���6W��x�,��^?�-�wug��LR��������1b��'�p%�_q���G�Xܽ��B����$AC�G8������y���Ą��z��7&nڭ�]�咶 sZ���� ����)���ҵӭ�:�鳍��l~7#���g���@s�]�`��.�Gl̘5�X{�d85�NΑ�d�tpL���
jN.�m�1A77�gQ��3t`f��>Jm�}�
�o�V�%h����otR�vކ&�F�|�d!�^�;N{�>H{=�����\f����J����yT��D3�A:t�-��;P{�����g�v�v^!��s��l�Gjt
*p;omv��kN}��s;'_J#73U#�]��Ar���&w�.=����Nr�]֗����/�a�Yt�[VgL9�
"�!�V�)׼����dH�A[���n�r�gs*�F��^uƸ-8�8��
:#�y\��iR�3 ��n���RK\���L�"��(�B�/�oz�-��3�t[�4M���Ġ۲Sxuч�nq>䝚̗(��.tM3�zQ(�U�<ʺ|ꕶz�Tj	U�$*����ǹ,��8��ԝx�}<��d��{�`�Z�;��b��b�1��y͇6��
��G�줌��ՖB�fon��E��4܊��Y��q5r�y؅��Яν�$ߟw��]/�N��Ӊ�uY=	���Vv�gt�n����xv�W�㯧%reM�&K���ҝ彦%:qvա�39%����i�v]Cd���2�,�uV%n>.q�Yց�o��߷��Ǆ���m��Q���K�iY���9,��`���*���E�����ب�6[��{����5ǉZ0V)3�Dd��%Նa��7����/��j��C\��Cn��D�p%��{��iL�js�SN�&��{���r�D���m󫏤��nd���0 Vt���y���������`�G��L�h�u[��yl�� 6w;�d���dp��(�B��Iq��C�fp���kٱ�δ�~{n%±&�R�9p�+ugQkt f+��ۜ�<����o����=�5'����h#�.ݢZ�D�2y�s�����u2_b�{rf�# �v�u�<,HM=��b�-3.ko�2�@��kwB��ΆS��sM�� :һ�}*�$����۾���<����aK�]7*�PR�/9c������:n�u�V�!D�6��:���v�ܬ=Œ��Xn=���ے�3E�+�D�����b��`N��<�O6�)����Ò�X4�\Z�~�2z���k���u�G]��N���t�\޳њ�`�s, �<���'S�|U�=�s&oP��n��q�����5�K� �ʽ��8tv_N�Q��nT�U���'o1IQ��4�8�Xux����y	<h��eG���Aqݺ�N��N<f�ؚ��n���ٛ��f�]�1-�7�l̩w8�ev|���8V�VT��C��}	�8�U:�z��d�ؓx�gR��Kޭfց|2�(�;o�G�����G/�
$�QJ�?]���p��q�GLӕGHA��p�HC蹳��w����A]�v92��ʾa�����DQDu{�QG��+'�Q.{�'���>y]�������y��Ĉ>e8��J4Q�s�'�}��z>����sG�"�;�=����TU$e_::����TG���u�˗��|t�|�$�HN����=�^��G�\yR�/Z�7��}вi���Th�wr)^�U����By�Ow#���jʤ;|��Ǡ��\��I+�z,�*I'��][���M�w�"?Y��<N�Ը^Av�o*.RE��/R��{�]c��������RE.��)�g��Q< @��Rw�
��Z��,H���ۅ��*�a{���i�_�!�֑N�r��z�i#��4Į��ɸ�\�c���*z:�R.NN���*��we�''3�|F�LUoq.G=/��<�GWLR}{�u�y.��8�b��]"������H.�E{�r]TR��-���}�����K�).�"����Vf���:��\��@��,瞌=�=�7�J���WL>��亷���l�CJ�����S���ѐ-��b��M���7��of���Q�'m׻��8����
%�5#�_ް�cy"����F��޸O��yD�+��V����}�h-�T�ǃT6��M�{�9�O\���9����;Ы�:^|U�a v�*����r�W�T C<��t�h���gx��8������	���X9$/��!��\1٦6�߹x{�3b��ފ�b�r���PН]n��y�;��7���V�l%�Z%Ňu�e�=G_����&��
�z�q:��:�{؟�;
�e��m��aڨ7J�^Sڙ��lot�}���=��m�q 0��R�:l��s��R�#nKU��_LE��DI��y����|��f�m������C�-�s^�cvo=5�o��W�������4�$��M<�=�}�^p��� ��~���W��s����V;`����SM��l$S��e��ࡏ����a1I�cv��U��qǺ�{"����˺=�;�OM�v��N'v�i�\�$����2��Kj�Gb��HAf�JL��J�ڇ��$gS�Y���ȯ�|j�]����/���{�6��@��vl�=�z�;�v�b�>%\��M�s��u�ӧ��F�����
��S��s�'��i�V���18vo{���[Z�q�[HC���`�X�-b�Z��7k_U�8����rw=[-��86�C\�����3�ԅ��4��G��b]���NdM�2�^���1zx�_ww*�-wZק���'�Q�,�C�c����{���eg����M<��/<(�����l�pu��U��)��[�ocj�ˆVO�(��lY]�yA&7�,����p]��<��,h�ѝ���[#B��Ilw���:�z�yo�a�9������>���᫒��X2n�.��W��3�F���~�͏=�Z��oy�0N�[�)�a���Z����[��2"v}RL�|e�h�ި���5h�Zފ;ؼ�o��*A7�m��Vxb�/�����z��:�WTg�Pa�[���,L-��z�	�����;� ��Y��M�nQ��E<�قN��5O���[��è*ˑ� p;�Jv�o'\�&M�!C�S@,�3���4&�Jx4�+����d⡚]��=>��*�W8{�~�s{�ܪ\,���el=}٨'}��=�E߆���^D{�
�[���G�߆�K����mL齋��_�熍���}gh�,ӽY-g������ð1�X�������6:�]]�Oe{�Gg�'v��R�
|s딆c%����R-7nYW�}��g=wx�XY�g��9~{5�9lOu-<B|���M���u���}~Uٕ�s׾�V�5z����7$��4�[}d;>��y�6�7����_������/GN� ���2~G��{����@J��	�Rs1��Mb����&��e7Յc/\�y���u��`��`5��`�[��v<���8�mϯ���Z����Ҍ������gӇ�W@=C��ꑝ�w��p}�v���"��n��E�ϥ-Ѻ8�p?%��m�od�>ѷ18����Dew�!Ά�Heٰ}�V�I���|
';~�G�g����M����u����ի�Z��Z�#9��ve%N�6s��DL���$F�+�����8����>��ۛV��Fڵe�X��x�2^hԃHU������8f�oz�x�*3������K;Of�,gU�K�b��&ѳfkUβT���$�wטFﰑ�j�a`��Q���Wr�a��;SD�F�p{ܗ(sʫ��Q�D1Z���xb��Q?$x5[V���[�8��v�s1�G�pn��gQ�<l���BSh���Y*�����u�F~��h>J� �����Lӝ�����X������}��᭚P:�~��OW�/��Cy14,|�k�J��Q���y�~3��������X	����{/FD�ar��
*���q���@��oޯ{�ٜ��������%��}�����.;�p����]8�a6O�O��A^O^8an�ox�C;��j̰��o؊�2�.�"�+����ա�>}�nJ͍��:ClE6/����`�UK����+�����	BY8���&��Y�}�϶]��XC���R��WuHus�
5ĬXs�8�]Ԧ��փ?�{�V�G>��m�߸z~a�)�S���\Hݲh����C�m�sjR�����jЛu^m�^����p����ЪQ��}�k)�;��P�JB1�;���n��g�59��[|��N@6RE�-�w=��O�B����Eĕ�2�B��G��OvW^ok�%-���=�Q�|��6��]���/9�6�gܱ��\_��^{2ݵ[�[A���g�y���$��n���l��y�S2�۾	�h�_W� [��2�s�9��pѕ*T�Q�/��Œ��^�U��f1@h}����p|eᰚ�ހ��Ƥ6�u����>��vz��q���Y��1G	�P�'�i3`�*w���A��dĲ�[w�.�,�G����I�|���f�sB�T����
�T�ǃXՇ&���1���d5���C�X=��4�xU�$��T����[*�T)5�ۚ�\Կe�a�z�,��!�@]Y׵��h���P�䐰�b��y�G�t_ӭ�鷋j��R��y�$xuS�]n��U��6=͊��R�:���E�j��o�ٓƜj��s��N��z���>��Y^���o��|x9�_�1w6����ۮ���7n�&�V����K��/?{�)������:�2�hϣ�lV�L���὆	:8�j�yg�x���n�sG3±��ma�ݣ�s��
�R������x�ݔv9t0g�Ic*�pE�w�9��wE��5��,׊�/$�HC�ќA�#=�^��eZK�;u��K�{��M��6⪕L���ӕq�ޙ|D�o�(v��?;x��1v���J��b~am�Cђ��*w'#�c�,�aQ���ؽ+0�D)��|�o ��d����]��ѯ�j�f�s�k85q~$��;v����j%����H��t��A�J��y�Q�z�ӳH!��6g�V����u$��i��(�2�}��8Fy��d��CU���ف�=>޲�.��^sv����5��lp��q�Ԇ�3����RZ���?>�8�]��ޥ�bD�]�<���;�y*b���K��]ʩ{�}k_���'�X*�T$>&<Z�x�]9���(6��Lv֡�q`����>���[&����� �ۨɚ���91�}2u�|��a{x��)�Vx"��
�2��,~���+�D��4�5��KrݘcS�RP�8�t��u �f��v�Ӊ/p]�^9��C��e��E���olj[��\C��8�[�}.U�r�S��v-iUc�tVWH�:I�Q��K^S[����d�]n�e�Ļ��)�bv�eaᓤ�8�]P�˓V�0�=ˤ��1��ڷ�u�o|��KG#hb@�ң#}��y����;�L��b1z�P/���U�-���7�
le�#K�{q��~1��'������ud�Lg�*�ƫ����[�ȼ}����Zp�O!Ċ��O���Jc��wՒ��V9�{�UO���S���)��[����s+������&=�0����G�߆�K��0h[W�F�j���-z�#w��\������X~�
a�5k����^[��_�hg�tJ�&3ם��d?;�E5��89K<��>.��ݼ��X&��ᛵU9��{��nڷ�_ٱ?P'�,n����@�.�l���\�@�o���=]v�~�?�~�~�S߉�v���V*nL�W�d;��O>Z���#���~��H���g�����C_��#�{��������@�a��(>��
�몎M~�ϩ���%���*ו H�c8zt��u(^U�޼����kȔx��`�Ʒ���yv�'���z��ГS�����e0�ljjX���Մ���oSY�zj�+]h�8b�|��X�L��G3s�3ZA�ľ��u���aF�B��.ȅ���:�����SCf�>D)�#>�V���06:y�Tz$Ӥ�? hK�o���>�����_;ϓ%�NWGi�~ �\�}:5Y�k>�xd�;��M#�޻�Qx�,�-��7t��3�f��Z̙=����p5}G���J5���o���\���D�"��]X�o�s���u��Aߏ�����T6�r�l3/(���R�GF���Y��f7��^0�>��+|1��:58��m[�޴[��U
�݇p��?zV�tv<�H���		𶌫�ܮ��ǳt�����;J�ƞ���|5�)�l?r���V8�UO[U��#��׷C�z|�8�`��?ug���p�"�[���{���l,�+��gb���N���=�����zy즯���W�	׫��~���ǋ�|���K#��e~_:�e|2��|:D	Aov��+sqDJ��K�h��n�9ʵe���㮞��P;9�TTQ��&.������W�(��o�����YŞ�=�A��s�r�Ϧ�%��9]]�[��H�u6��c��8t��>�]�M��w(�y���r�A^+����O�shZ����~Ve���۩^�:�����n.F'�՞�����ߦ��6'��Cv)��`���Nz��ތ��<LL���5��m7|E"��]���ِ|2�/xZ̮���,��V/J��F03�
�3m=���'�:F��:P�!�3.��5�*S݇�R���{����o��m��X��e�3�]Sp���2I��b�}�ETm��P=#}r�7�k>W�s���53+m���=#v��?QY�L$?W��&ߞ]
N�Uҙ �	,�7e��^�}�tqx�U_z�;����0��ܷ~N��g Oz���Ƅ�Վ�{��/ޛ��2�����3��_G.��m�l�*�-?G���s���e}�)jg(�8��-�\��f���~*O�=x�B��(p���f,f�#أw>�����pr��1�!��5�n��(�-��[R��:�P��v��"�wJ���ٱ�k+�|e�3C����oB�N��PVi��
�tc��%}ko�ҏ�|�,rl=��N�� 4�q��\�ve$�ohd���Y&.�O:�2�ߺ�o=��4�xU��9��X2�*3i�����Sӗ7���/o�w7VG������z�y-���B�$8&ز�#[&�F�n{|��-�M���_�O��.���nj�g�Y��lU�`�頯`,=u�Y�̯_��P�}a�����`�K�q�-������gb��a}����Y$T���*�:Z�HL=�X=�@.R��,x{����['V͏�2�}V�}�����*TL��qm����;>�پ��V3b~ao�ב'ʧ�U����bV����J�[�4��Xk�8M�4�=���υ�,L_v����BA�!�$2�B�J�M��o~��a"��y��e��;��!�׆���~��pM�ߎ ���S���}�i2�������:��~�JR �C�pM�ٵn:��c�$>���.���o��aE�4j�
�ǶN���H���	�L�6$��N�2mμ5,F3J�'�YV�8�J"z�9���Њ�v4ji��6�΋ޕ�HWC�q�&��,4
���˳٧;�)��,R�g��hm��R�v����4��8s馟D�{�e7�A�/z՚�٣ţ<�\�|=��%ŭU���*}��6��
a����U8�P�=�����|_P�6�jI� �w���v\퐴c���-m
��%�5�ޡN�]+x5#C����5ox�K�{~�	F����w v���J��GC9ǧUe���6g>��Ȍ��gn_1;+�R�Wy�s���R���v4�崮�ٺ�id�r��r�Gs��Ӷ3a1�]��6R�qFfnө�\2���1=8&����\�<fV�3���LQ�#�h�Z���"&yM'�m�	�m֕�J�ULPY��a���(���*h!q�y�Ḯ��#\hݙ�m�*Sp��c0�V:�	���.V����|�T�k�?����;s3�Rj�c�Tь�� ���ε}��,�����9���W��L����OS�7z�䖴�,�;��wuo�'7"�C�	[mh��%d��v�W0j��]m�RJԀ�p���NЭhS�u�����}�.�l �$w��P�M��=�'V�%>�-����R�J�me����4�l�M���~�gvc�)��y�z��Gz��zp�E+"�漯�Dh܇�^]P�;�܋<��g=��vw��8�Ƹ�J9����+���u�+�2`3�$��y�'�h�!��:���j��x��!%3��g_{{����~Z��lU](�vD.���;�TYs���^�Y�p�"BE�ښ�L�.��;�Dy���%I��c��
_'��u��Pk���@V4��� 1s��F���0ܬ��|��y�v�m�,��9q_�������0MO��v��Z�T�W�o�Q:�]�ۋm��ݤ �$���Z5�� {$�y\6h��s���W2���N��
�n��ܵ{K$;JbKi�ґ�]�#Ӓ� ��ԇ)j���թ[b�\�Vi�b������OYt��a���K���I��t�&�t��:��.]��a�{019�3�j��&�+&ݨP��OWX�s0oc������\���G�g��׎�L+�yk��X�T�Eb=-�J��.�ϡ�gm���|�1���S	��N����3R����:d
m��:���IF)����,^�q9�����h܋�J�s�f�x�ԧ|lp���9�Bhr"=;kQv�5��.=�=:�B���xq�����ǖYW��>pLK#���@�4\כ*�3�nL�c3h��)r
c�PtZA�[��SU���Ւ  �,
`�7��s��2!z'^����t.��K�x����p7@�ȸ�Ȟ{��P'G�1w���"� �[̚Cq ���(�R־�RL���/�݋zո�@�*�.	���C���TN:�D���x�U�:��4Z�9z�&����|�x],S�{�9&~y�n�޽�r���Gq�����h��>q�^n|���q��B���Qj��]�N�Y�QA}�s��N��WB���;x��������>Z>NQ��n.��r�	g]]nn��y�Ot5炷wu��s���,�{����}ˎI�('�__{�z�U�.�I*k��,�z�j���N��OWwoE-'���p�x~T�yz��79�J�I�%�J'���'�|�ETS�e0��Wu���;��y�Ēs�sw]�3���𓔊2��^v�I�Ģ�?u�����*�]@��^���qx���r�N%UB�t}{��纙���ċ�Ҋ�C���zaPS?'���������*)���Dy���n�w<5x���y�r���X��T��ʟ;�8Qv���ywvz��众_!�9�%�z�?>��'+�JIRڦ�=S��f������f豱`�|qN�-w޽7�]M���1��i�+�aO��9͡��L���!ݵl��'����r=����7<OW���I2��R5tu@�_@}RG��wz;,z���0��G_1��`-��}ʰE��Z������)�ݓ/~o=��y�nOEN���#J�%��_cie�M��:�8�Z�&�g�ٍ�K��w�P�p��_H������8M�.��]�
�h�B��t�m_���kL�Ԣv�f��U�}���S�4�pB6���-�[þ�ww�����(�z�������%C��z���m|8����� \O��Ҳ�z�9���h 5(����c�Ւo�)cW��ZށG{�����z��tk}�Լ��SXߘiL{=���o\N�T�tm�L�u���ɝ��~�.ݜնl{�	n5ɮ��c����Y�g�W�������׊�;a�j}�#�Z��
�u�,?g�0�]�ן#yzi�ƽF�3쏺F_�rl����s� ot�߮Y�}e��,]��m��)�K�$[c(��J���� ��� �sJ`���;�B�Neo�f����ri��'ԭ�a�7d��E�
�H�o�6�����-�s���&TgBIuO�G;hd�zֲ5Kf���z$x����Cc�y�i�,'��i7O�lDF\���;�}���ȳƯW�wo�{*�bh7�CoꖞB�W�M��Q��
F�U���]}�b�<���'�؍�|�
mK����=�~���)�{��g�n����m���6���f��3�!�O{�!�6��I����~���U�"'�b��X;�p�k�X�ߜ�c��_˭Մ`�)"�y{�̱�^	��J�lyڻg���ϳK2V�w�2m�N�W�����5&/<^�2�uCC��ԆU�_9*�	Ks97��N^Zk|!�'"��_׏�ܵ�Y���������*��j�6�w�5)��.}��i�X;��^�T�i.��>>��'��bX���.���A��5ݻ7��R�:l��m�NXN��o�:�����o�2f:�z3���{��PzP5b<�����Ʌ}4Eخ�<����<�d�XkT��cX�v+�x:{/[��:J*D��o9�%H�p`�̥*���H�c˓6�͐��3��9�I帷��򎳸˅�S��0�-ǈ+�A����q�mn^��cFqna"~ĿG���|^!i�4f���5��1��J-O�v�
3��X�y���+����
�$�5�>׀��ʣF��J�e�ſ�a�����F���s���(��J��ͅ��&���G�y��;hܣ��tɬ��y���t=��'�����fsy]YcŇ��$��.w�5W���[Yѩ)����s��=x���x�����I���ѝ�zڊ��s��I�Ȃ��5��I���yZ�H����5r�6(#��ۊlF'��s$�;m(�W�B�M�e��Kd&��"�2�a�d� }������&%�佚�na��62� ϡ�����e��6�(�g#rTUN�Q��>[t��W�xq.!��`����5�۬�2��6<�s^�[v����o�Q����w���[T��j���6n��{g���S3-��{�ֽ�qM-�w�C@��m�q�RITȜv��p�z�Ӥ"�@��;�G91m�v�s�^�S@�,H�5�Ӯ׵�;"Eq�����܋�˱O��A�x�g�<W���Fn}����7��G�e�9θt��Xs�7��I*{L��<e�����=B(G���$�Xn�ϕ�(Gn�n�^���W��}��ޒK`J���=���$h�(P8�V:��?%Z��ِw����Af�/�K݀A��
'�iXg��B�~����)>��?��o'Lܢ��x5Q���|���f�sB�eQ��=y��
�
����Gh�p/2sy�?��;�z��R�������Gpӥ�Hr@�SG�I�Cg<�Ӟ�P�gr�'�*'B�5躵�Ev�\`���W�$���归���k.�g��$j��}Y*��G��j�u���W�ÿx�~��!᧼/����6������"֭B�����d��BY��� ���%�Yv�.����?<�{�%n����k�0�{����cݮ���V\Khh�T������\3Wd��:��Z��+�a�qm�~v�;>�پy*��$�o�޽�X��-$���2n������eTx��������W3r�l/ GP;v�%߶�&��z�o��.)�!��{�t+�J|W7�	5��lRv�k��B�ԹA�,������c����r���)��?ou�dj>N���y0��p�ߣ��u�5ol���w��JB��|��j�2�X�%&Ц�G�"khC�^SU��\xz�y����f�;A�\�=0�9{
\���i��GY#0wW����f�Gc�ĭ��7%X��F�L�A/D��s�'����q��^y�3-�ғ�q?�7���7;��I�z�X�ֺ�[�r:�=~�d��1~ٴ��0��I�&ڹ�:�i�B�(�2�T��
2\]��W\H��[z�.]�MM��U�Zק�`I��G<-���;���cw��U�bE��R&��'[���ie��d�X�nM��u�5"y��x�k]���FO|�C�~�L��z��,�#�
����=�v����_"�o����[�jq!�85[W�Z:�7��OX����#hT7	~�P�ƪ@�ժ���Y�MD��-�[�5���-��{o���#n���v�p��]�`��}[��3����֡Um-;��~��m�[�a[�\$Ɏߌ����ܗ�-��W��(Z��y�2�'W��'K����=|��`�#q��-=],��4�ѕč{���Ը�j�o�����;ݺr	�<Z�E����}�>�$�c>aU5\�n3�|�g7}9��z����`�7���U�u5��14�+=��VJ������5舧문��9vL�C+�=�n�V�-�a�
��X]`��\�(�(�WY�.*r=���ʶ�����h=_z��cE�o+��Ň�v�����AF���]�@ޚW���YHu���lI����\�.�������	�v��7˳�LfW����{�{�����d�v�=��A?X�Cn���B�U��c�4N㴻���8nB�ݛ⇓ō��'��nK���m	lu������v���}3yz��7�}���i��Ͳ��ͯs8��ǽ=@�a�H��g�ok3��<������Z
��g��f���rO������F��r���s�n�Qk��8�^BHN�]��|ol�>]������w��}:t��}�u��ۆb�ܳ��^8������ ���7{���o�M֌�.<��*�)��6>h�^�\�L��b�5B�?v�Ԥ�V�Dz��5�ф������!m\�����w���nL��-Tj�����+��={�����_��m����G���2�����V(K/�ro���N�����x@g��n)�̯M�,w����#��`��ycR�q>�1ps��]Zf,��%��^v�n���X<�7����n��Zl25��.�d�\p�
�7_/$B4�8]a:VvpC�j$p1?x5LGU=����{"��0�r�i�_��K�ƭN�#��m�\1Y��c��xd�l�S�U�wh�ӵ��c:���ܜ�D{��P�K�	��&hc�jr��[6��^X��BQӽy>_eƏM����Zۼ�5�|�X�Vޠ���Y�����'�\!����+���u�����39�������������=��.�����Ǚ(�b��z-�y*�CsE'�cϴ���u������}nb���*&w}iJ������E�����y��r����S~�l����W����M��7u��۸�=�g�n��|,�"hF^�=S���wZ�>��V����K�{��P�V���fV��u��6��2=�vWR���8ͥϲ�t2b����Lt��=�}�i>˫���f�N}0�j�	r�E��w���v�)��v����?|}����?7���1�r��'yOU��EEhlACT���ih��i�j�(�:�7�wu����Q�
���m�>z��o�g��/9���u���a�'��<P���ԵL5�_U�&:���l��'���U�|���̹��ˋT�I�o|n5-�L��^*�>�n�G�@�PW�YX�y��j�;�h��>�U!}�)S�{�oīB�u����w�y5WNe
��R�oL�7�Sr2LV����j�0]y�X�O݂>�Q8�[J�8���
(>�'����K�8R/��׼Y�ͬ��kB�d*6=x�B��]��^y��B��Ct6�������CN��h$x��~Z����F�^��ԁ�B���>���U�V�[բ�zڑ�o�
䐟��ٽ�z#jo2l�w���x.��P������o�:t�5��';���d�����t���]c�&��w����ߑ��rܽT�-�o�wr��l��G�;[n��}Hˁnq�]��G�_j;�6\u|��nC)�F�g^j' ���U�=+�nӕU�ӽ�hX���χ0Gw�xg�-p�f�yGx*cUNc}W�þ,�˧W혤�>�v<{9d� ��K�OikcK"��٬�f�F��Ct=^�'s�b"a�	�3���|�ez��`M���k�w�ݵ����ݮ��U�Ā��
^?B���Z�a0Gy	�hyqk��.�y6�j��Y�gϷ�6�U&\>����]G�wws��\0Guv��
�ŝ�Z���|f�yM<�C����"�qoW{���׆����9��PgИ��Pw��B�J���z�lb�[�����3<|q|7�x$�#rWm6��s�Y�z)�Z䪺���Fuo)���f��}]��aoLڷ�Y�Q�������~U��d��G��\d:�+���0����7�8'�����]3�D�Z��l�׽����K�k>����Y����-wZק�ziN��ba�׽j�+^��v$�ґ�v5ZC{C׌�=�Z�]E 8��.��p���a��]���!Q`��膹3��B�����ֻbsT !���u-��V���M�?���wm�SY�^��)�Ͳ'�����p���㋷�K[��i8�zaظ��ac��������=��b�җ���һ"�6�z4�n&+��ܣ2�M�Y���Y?P����C=�z�x��0���Zo_�vy �l�Tf���N�壍�^N%��j��z�7�S�4�jO��oQ���3�Ǽu��t��j��TD��\<��o�M�6n��Q��+�"�������3x
lXl1\���Y&�Q 0���m����.:v�r�V�]{^-l���1GSM�Jb��c�Ւ�����0�ߛ��#ݸ��iP[���]�նlx��V�X]��[ѕ{ڜ������$�n4=��:�{�͡^����1N1�Y�#��ӵ��=^��\n(�zs^�O^lO�=�%���FCe�t���gv�d#��9}��R���n�=�f��O�&�������A��
�A3P /x���vuݏ?b �e��-���*�m�Eޭ�=w\� 6x���7�� {����d�ەbb>OW�qa���x���nR^8FGM
���E��8U���dhwF�F�d���\��ad!_��ݕ���?wN��ʁ|	�����q�m�މ�O�f쮬3���*���p�9_�����s:�c��WQ�:�^�A��zrd�F
�Wg���UPb�E��3,)[}���X/���N�&���ܡ��^W\G����&s}]��ᐕ���!���t��nUB��J�¶㧕1쩝� ƙ�F(�����gq[��V�����d]fmx=%�4jy_���Y c=d�U{�C=}��� *�H-�����s����s^�C�[�';8�M<֓��}�(���5�Lmq�z.��[��U���w�8N��+��x�=�(�l�v���*R/T�;R���V9T;N,0���I�ZW'z��rKzu�OL�lnŠض��m�?3.�4�E�a��4�Q�Aӻ�w6f�tx��������l�=j�n��c���=�ɩ�C�J��kIk����׳kS�`}vv�i�Ď� ��w���橹���&��,�ݥ�U�S���q��v:��]��P%�s������F�S�2���7n��Nvŵi](f]�%��=u����:2Υ3,�RȺ�=����LK���ܫZ��V��~�D�L��<���A$�<��я��q���z�k4��s�Tl�GU�Ȁ�Y�D�K���j���ۥ[o{ArG&˭� Cr�ܴQ{�����ɻK�^�j��Kۂp�-)����ޢ{�e2�@ˈ�׀���k�ڦ�䏝��x6�)z�.޽j�m=1���q�viR8��Vq�5�蜦7X�q��Qd�b�����;��7֕�%O�$��=��?����Y�I����z�����s6h{z��j��d��m�(�����|D�\�I��_90�kzi\����i�K���H\�zR�~M8��ltԩ�y�Ǳ�a���΢�v��Ԕ̏�)���)7J�C�w3R��z�t�櫵-X����ě�"�*��œk܇T����w��G^0}�N�`��&���d�[��Ff^�]����a��!�ҋ�n�X�Z�{4�s��'h�Ā�Co�[���4w1�|YV��x�gp��*��9x3mu���}��r:�X�d���<}���	�c ���l긳kU�w#��EG�
�MWC���cݤ	�-���G=���8�T)�s��$�T���UX��D+�����{I�ù����AK�D�A�Ì�w���uK2�T͉d��u*�Su�4�F{ؼ��������]��Gc�8G�w�M�_mJ{Ӳ��v�]P�ԯ�.����X��)`��m����13����}8�
�R	��<¨�݊����;�(�N�=���⃝�'��G*�G�$���ާ�8{�޲M�����;e�/�)�	L(���I!^Nr���w���\���.E�7\�:]�*���Snw]q��c� �QI^x��@��n	Ӳ�39VE9�W��6��s�/qY�r�'�624��'zܛ�4�ΐD�0O��^C�Y7;�9x'4����9�7ռ�z��ܩ��Ӧ�5�[)�RI;u5D���I9U�I9���ҡ�@S(2�*�F�
��*d�\�L��d\=d{�x�U&j�����t�s�2�I=�;+��0�ӆ�Sɏ>G�ܐ����]��Aʝ_tr������Y�O����D�*.'l��I�Ą�"G�_v[��G�d�N��1W� .���_�����ZiZ[��wW+��Mf:��,���I��o���N1�Ԅ�8f�do7+%t�%���X�����v)��;�r]�(-��:��譞,xڱl��/=
�!�1gCw�>SC���Ͳ�tٿ�^�p|����o���դ����g��p���@�>�x���٬ �e�o��c�u����7��؏}����ԡ��ʀ}_J��d�Q����4�+_;!2m�m_�"n#���}�@���>7~�GS|N}!�b���_Z���Z�[�G�>m����&o�G8�~���On��T�h0U	Ճ`���,k�3ݽ�>�_�)�f�%y�VR����6g�/�}��i��h���A��]˦EvÈ߶" v�w���n����i�iH�#m�NXN������r0h䮶��|4e闩2�ϩ��5�8����e����j��>/��vњ�p�f�V����|Mi��=
�����ul����/r#}�W$G|�w�} .����w}^���kyRu��:��|� ���G����C7��H}osz��u��G����t���^��c�K���؂ߒ꺲�E����\�B���Y7�/<��7�66�D�uj�;|�pz m>�룝��Fʔ1�1��\yt���~���u���<nw[��5�\�X�5�Z����7�&=�Hq>����gk�f����>��{޲�3������c�w=�.ٞ�&`#���-v�&z,#C776U�Q?0�D��\�8�\yul���\��n��iXR��t��yZ�E�����w�A�Y~��j��gR�YּzH��X;+�u��ډm5i�H�τ�]��NB���ַ���'����7�6����Yϡ
~S_{��a��M�`�ǲu���ҥU�^����[K�Y��P����(3u�l+x���m�r�R�q�Okw��8Ԗ���o�y�ͪ�X�A3r�7�iVQ��x	����c�c8MN=,w�ʳ�G������g�YX�t.�������y�z�:yO/g$[�ee[��Y�ށ!5���Ԥl��+��_���+�R8Z��;#eI�%��k^��U��*��u�A�:���ʅݢv����M��tOǵ���v��0e��}��bm���v�dYB�o�d��#��b�L��*xϤ�j6�aֻ�`�_�u����&����#�^Cm��v�t�|�� Q8�[J��o吨����VM{�)o#��(� ���Fx��sk3~ZW��.z��~��
ez�y�za�����ݫ�����G��4
�/��f��E]h�]s���>4��{��D��j϶�����ВF�ʉi�zg\p���&�)�7��@jlZF+��(tܛ�LHaU5P����}�^��^���ߙB���KȊ�u-B�D�������:�G�	��oӷl�~��~�짱ą�f�ϖe��VX��h\ÿ��Ϣ��]���}p�7���k�u��RZ���#��ӿy0�&�|��;�f�,�H.���H���y��&����O:,x~��
���!��e�c�3�&�_wx^�Nm�w��r,��'v� Ыȡa��hz�Kw��B�iW��j&^,b'"�b=�sF�Ta�9��FfpRѲp��V��Z����U~t�[�=�Z�Ŋ�W^ʙ>�c��b�BvW
{�<��'s�Pj��V�6��q}�9����[�F�Xg��SI�n �	�V$�e�[�xh2��o{o��O#����M��VFJ�ɳ�����kP�n$��^�{���M7��d�2}����}>�N�~ɐs�'4qS~����=m[�u��w��?5{�O�{��ζ�}�r���lq��BiX�7�W4O޴�wE�t4�q�-��LP�L�!׬�<�
jH���+�ֽ+ x����3ѧ���&���=ju!�:�|n��$�ϸ���Yt���w�ܹvov��3b��&��`��BG���޾�ǀJ}p|�j��F����r���& ;�f��G��'���0�|6��:�C>�<��î�spƯ5�Tf�(G;XTXJ����'�%�hx5@z�����ˠ�J�S0GJ�3:�z���e����V��x
l[a�>���d�z�~bdk��?��5 7o&?��?��}��ſy:�b���5��1m)���}Y+�����w蟶�6;F&��f��Ú78��Ė��v�K{/'Td;���b�YH,�:��*�ӟɺ�����nf�b��{3^�@:Ek3,�k�XR�Q�x0��bl���L"����<������G�����Cb�"�{ڳ��?z�}��oDn.{4��9�V_�*���3ݷ����2ذ��䵬�4����^�\�f�]�	�͵�~��AT=^�-���z��x���w?g.H�VN��r|���~�#���_���\�0�ﶙg�{z6���\F��� �}�ɀ��,׾^ݾ{.�lH���3*Zt�y�.������b=^�4a���Y�KO6�g���}��T��ݏNyMTΈCmP�޳�w�|��
����r����+��^|�>V{Ҟå7Qmx���_�xsBéA���`���sC9�XV2�9�k���;Z��a
Wfb�}��8�i�t����4%W��s�{g���l�n���;:�dF�Z�h�>3hjv��ޏRj0ʞ�dQX�Rܣǽ��,㮲w���KI%w���~��_d	�>{�!Ƥ&�M��@�zH�a����tl~}��}r� 4H�!Z{�0�I���ݿ����():@���.��G��B���HH,�[�5��-a��V�<�t:�^c��u�)Z.(�Z��Q�v��)_�{Ψ�g\��z�gen�T�i��t�+�;�6d�{�\�>(��D��`��~��g3wga��m_Z��Խ���K�����]��au����	Ұc�pC��D�W�ދ�F��|���p�H\���߽m7�8���e+B�@��35��{)����~�{ݱ�r.��WQ#�cU]Yy=�kG�V�P��B$GI��B3�Ң��ݵ�dxԯ��8ke��ht�-[�U_��yz�6I��j��+����3�E��_(g�s�~��HФ`n7v���j�'���|)t�=�"�7�t����K�=̛�U��Ha�h��eU����h����+���6ݼ�zҰe��-�U��� ��5s�^Ed��+�{>�.θWk8Ca�%!��v���SkB�omؔV`��5B�3]/��T���f��V�Z��!�uP�SK~2�{��k/X���vk�fe��mk��HI�Mh�v���=�=}:��,gzU��H�bH��8���7���{��DN�D�S;J�<+o�],�AP���YMݚ�ڥ��7�7m>�h��5��括/��%�W;KN�b �_��SS*=�l�F@�ܑ��n��s���٦R��|=����R��o���r��mmK�O,{%��W#���������vj���$3j���yP',������K�eL_��|��,m2H\e�`��F(A�`�(�w�OL�k\�y�������ֿ��^��������t�����`�@��hT�?A].D��>��y��;�u�pX�:~�\��m�i3`���>ȼS��ENR�gW�� �������Ĭ\��ߖ���U�!�����^�;;��4���q���{O�6��=_�^hC��d�@R�����O�y.��Ky���HapՃjޭ��kx����T��V�B]� �����:nM�*�5P���V��]x��ڱZ��yZ�|���kY����qc���frt�H��g��:���8�o��ePgM�nV�M2�˛W���PѶ)�yXB)���\�BZә6�o>G��WJ�=��O�w=*�[6��z�3sʚ[U�S��6�hEئ�rP���j��'�ε�Ÿ/�^��*���֎���I<�`������#�l/��}�|��ouXl�/}���W���#�{q�E��{�W*��G�`�WӮ��y���ɇ��rm����Ӳ+���_n�nm?�����Jo�fĄ;h�߲��g|��j̰�K7�r'�n^itM������<m���b����-_�-��=�iSK���7Qu>�g�
�����,u��"�}'M�ܗc�	eKO��y�vѱ��apR������C��e�M�fՇ��������?0����3۷\�'*�rɿ0lN,��|�֗��'�|qs߂i2��R�GT�ݟ������ؽ�����B���I<�|
jq�O�k^����o�b���]��7}�zP��2;�!��o�S��>G[�m,��4fw�+��#��ty�p|j��)��`?1�R<���;��o���Y��T�M�%U/]�X_Y�c�3cR��g���t�.r���w��:�>�F[�r�
����'VmFWwk`gg{��Ks��֓t���?+�,⨝����[�d�X�17�dǂ_|c\� 蝗Jmv:&,�9�5ϫ�lUWU�/z����c�nP���	�������F��hG`�XA�_w������hZW�z8{������}�߿?EA�*��k�O�0�9���T1GT��9��|	���^��i,��u�)�[��Q��ud��QY���T��k��/�.�o~���|�}��*�$�z����c��+��r���QӤ���O�U}�MNcUF�V�-�:´�����1������J�O�CN��:�A����ǿY��]|X~6⟫&����wT����J�֎o��U��(`���\�0�����}��p�r�#;���xU���yL����c���٠�ġ��rlL�ts�գӘTGl�cL1G�X�ma�KO6�d��ܗ|�F����%�t.�<��V��`aj�v�v|��+mɖW��y��'��cm\×���йY�V��� �ܖ�����Rm T�5F�zc��`<��M�_�i���ir��m���D�j��%�-��#�{�����$.ջ=]k����q���e�C�+�pدX2�oy�t��!o�㶱�Z�Ԛ9�7�+Tլ���|=����MO�~c�cjX=u�l���u���g�c/C�}�]���+ў=�@���XA��3�J����'λ�/������+��z���8��l��>�S>�G��4%�b��ࢱn�1�$=.�:_��R1G
Oo�g㴶�����_�q�$&��Ppϧ<\�yT��Uu-+l�d�\�
'0R&��`��~���7ޡ]�}��f'�P�z^�ޥ�54s�]mjp��N���g?P[9�h���o|q�!U����$�m4�`֭O>tE|H�e�4c)�o֫�^���}�A�B� �=@z�B��M�7���ܷڅr\�X�"��쎻��ʈ�hX@�M�I����c�ֶ�=�����N@�dL
���9^b;x6Oii�e/-�b�`2,%S�|�������~3"y�QQY�AA_��g���6cl�'�7Q�-�IN�0� G FC � �  "` G` G` �>�<  ��� lG��m��"  �m�D��"m�țm�&��;lα��m�Gm���dM����D6�#��dv6��m��Bm�Ȇ�dq��m�Gm�Ȇ�d@ 1�Ȇ�dM��&�Gm���dM����Gm�6�dCm�!��m�D6�twc8�l��m����m�&�l�6�"m�6�dCm�;`��;1�8&6����O?� `�$���D� "C�vr|z{������]���y��O��y>��>��8��	�����?q�EEru=O���oP�*+�� 
��?hyݟP�G0��~��k�}�(���<`�Sb�	��#�|�? (1���=�/q���;	�`C �����6 ����c&�`q����v !�q�w�r0����ٶcl������z���|y�b�v�B��< ������/��'�9ؒ�Z�y���.�sAS��"���N����+��TTWb(���� ?8%E��G#ATTW#/w�%��0K�a�3�T���������������_ӻ��*+W�L�����3�vr|�������������:��(����MV�@t/XI�1-�?oݔ+��9�0�qTV���/@�z�_�ǆ�a�5�������h�oaTVc��N�,�n��������)����6,�8(���1$=��EO�Hڶ�L�f���*�u�-�JZ�J��jJ%U*TT�[b�U	[5P�Sl�P֖�I5��֔!E%MR�$�B�3M�5�ko��OS�;�N�*�Fڍ�ȍM����$l���j��T��kCV�zwj�m�U���)�w1�5*Z�+�km�Q���jv�V+Z՛ �j!�f�l�hԢFMjͦ�,�iZU)�66�T�P����Ij̲���� ��cX��V�X�j�IKJel0R�m��n��[-
c|  ��s.��Tyޭ�tz�=b�w74�z�v�^xg�OZt���ڥ[]�N7^���P=iÕ�{�5����w���t�{�������ܩR�h7��h�j�����[S1�յ�6�Ud>   }����СB��{p�
:�l/��hP�B�cB{��xW�ͬZƙ��&���{g[d���v����r����	��I��z{�����n����k��M���{���m���-�jҵ[cmVmY�>  ;�4%��t�=h�w���som=�޵穜�ny{���f�v z�\���w�٪�{v�v��Ӡg6�P� ��랪��޴���Ǽ�o{<֞����{�kf��j�[MeE6L�   -ާmTo��Y��mCv�O5t����6k׻ݽֽ/]4=:r��jt�wn��n<��{sOM����^Wm�P��]8�Kmw��yTu�ZS����fɶ�V�&����E��   v���%ќ�p���T���-��ﻮ�(P���A�5I!�{j��{���!A����TV���y�nrbDkV�kTM����   ���i���%�m�#U�)�C�vr6�v5ջn;a'[��uPP�;����Y����j��:����wn�@'vɵQ[�.�Ղ�cj-��  ����[wu].���UAtd+]w!��m���gCA��w��wA@��*Ma���F��pᆁ@s]�c��飺�K�5��'dڨm7�  �{�  ���
 ���n ��0 ��w ���{��� ��0 Q׷���)@y�ۏN�ҩ�{k5��l�VK6��j�ڍR|   X�� �aN�@�����x��  v�s�PP ����T�hc�:h���zWz��ӯJz{� ����[V٫P�`�V�h�Q6V�   .<�4 ��z ��{^� �;�@ {t8��z��� �{�n�� ��������  ����  |���R� �)�b��H��4i��L��JH  "��4��A� F�T�� h&R���� j�����m�6-���Q��Q;�3eG���ǰ�#^�mLURi�sYnE|��f�3{�������������6m��`�1��C���l`�cc�����@�~�O
�By�&\+.�.��m
��h8�S4Z�����AKTޢ�#��=��b���xLfՄ�Е��@���_���o�-6��*��օb|�U-`�RK�L�I�M�F���tM0i�*dCH�Oh�f|r� ��)1{3v:A)
�H�y�����54�Z,��m�rێYJo j�f��X^zF�*@UF�؃̘�nQ��KO��!����*��f�m]���ք�u�Hi��cH�zq�RH��G%[,����7ŧf���5��v���2S"ܳT7�@(��VCW�D�z��P��&+��#'r���nQ�W��ۉSN�B�7�މSHْ��� M�O������i��S/D��4��b`���I|e[Q¡jkkJۺ��%��
����NR+f�;�dH;��=�+�#�vj������ѳI��֤�
�Z���x�+��R����2LX��dZ�4��t���<p�������6��+�8� �[�7R��T-*n4 �51�Ј��ȋ
���
���˺�`��P����0s�U�:]A�������N�#D�&̭و\{C`Lր{��*�Tu�W�Ulf`�@K�[gV�/�Z��v�$��d��V�s0��B6�8ay6@l���D錺�U��B�e�-J5v�:sJq�/۷�S$�N%&;($���4qjB�$�Q��QՑ�`�D�f r�Z�8��/�.�ɶ_c�ԫ��sf;�z�5eC�	����5�a3$F��� Ae`��%=�lS�7IFP4�Vr�rhWZ���ޢ�۰Jݏ@��n�76\-S�fh&c�h�������͏�����ef+SJ�e�ˤ�uҽ`���%hZ��O��Df�N��*ZT�x8m�E��ѯ>����,˅�0��	�����K��jQ�"�z/^�`ٷL����,#!��5�a4b˻������RۧK^ L��Q�Q���"~`�ʹ�tn��x&���/5�=���h�1)D�
��`��q2nVl� Y,7x��[���6�Ѻ'6���l�/�!ʖس�p�Bimu9̖-�e����M��d�O�\L7�:e�4��֪��Y�2�U�/�f�م�̰"+2�ZK(fT�F�Ĕ��Ƴo�Ay�6�ڭ�	;��A��n�W0�%d���D`�d��n<v(S��2n��ҭU�Y����:ᴢ��lXy��V��HlXp����tE�Bҳ����s>ٛ*1�v�"c-J%���[���'sob�e�.5�uu��y���{yp��	9wM�k�D*{��4_�RT*nZ��nԀ��9���Y T]�A
�;D�Nb9�A�3��0ٸ���B�?i"f������{Ked!�T^;)�T-|*�W<���C�b�J�`M-{�-N�
�Ja;W�*��D�hQ�w�̈m�%F��w��m��{%^
/%*�}s>�]pԠ��:JAp�%e��&����.a� H�#2�J1f];�z��aR�oD�h�.�����tL���ˍ���`�Է�����D��+� �zֵf��fnʑ�B1��5ݣE%�K�v�:���R��(��З�2�V��r�̔�[d����w����*ڈ-�w]Ne�ˣ�]-D�BY��gV���إ��2�xu�u�#��*����5��NU���9��SqA�±@�3A���ͤ�'�!ִ�JdYtnc��1�޽�y&���R�
9�ڧ$u�ͭ��V2�cn����g�
���21薶�l�F�D,���;x
�1� �:0���n�e��) 3h�Lݪi�Ը��\��Ge�[�D�6#-�,:4�U������ǀl7��Yu����,zO��F�5�sfF�or��a��m��Bb�$ݼ�ҥFe`�rkrf���ł@�0uZ	�c*�̏(���Y&�"kC-�vo�(��:�2�^�3Oc�L�N6�5c&7.cץ�%W���V�YCuc�s�N+�tZ�["Z�3tj�Pn�d��/�Y	@���-�A�e�vث$�e@�����Wx/��3r
ۦ����sbB)�U3�5��Uj�ӛ#Չe���f�e�WpB[#CYY��V��--A�ti�?H!�����0���cV��N[,D��[�;����ͭ��Ә�dMi$�WQ�+��E�]�m�c,����x6��hX��7� Ӽ��r$�%f$�r���5��
�6ͺ�-��{B�+X�f�3`F#1Ä�(���6��v�m^�v�ͽu6[�`��%$	�G,Lы����*X^Q�o ��cxn�7L�(�*���K)k�k���bY�m��y��u;ӆ��Ɯ#�<+�+A�e�D�̨�xM<�B2қ�7�4P;S��m��y�Fぢ�¦��)n�@��8�׆�9���a\w���mK�Q�l�S�lҔv�1�յ�H�kJ�WZ�(�K�X�CW���q#�K�y��	�cMڇ42�[mH��(
)L��^^*f�Vu��@f���2�۵6��!%�:�ڙ0��ԫrnǈ����N��/m��V��VMlӔ�Х����R+�Z ��Xd�K(
ɽ��rջ�p��!q�AQU�Ϧ�^�����f��i�YS)'B5�M]���j�\���͹�������ʔ��޻�4�4Zq��@��47r�s����7]hp��ɓDe�����Q꧵�N5s%,-P��m&Y�j
0C2�#YD�]�$hZ�b�sU	�� b��ܺ5�MylYܼE���^���DLv(do�֜��9 MY��*�fЏ���mVC��/j-��&f\�y1l��3w	[tN���{wN��`1��4X�;B��L^R���{�mG�,�E�8�b"X�Ae
z��j�C{L�Kr��Ċ���@���[�wZΧ�Kwm���f�u�-%F�İl�ux�ML�X�͌����m��] 6*Rڡ��}4^�40䲦�v��C/vku&5WI
V2��9��Y�ۓ[���h�JX�� ��N��Q鹪f:4m5C7b.&�v1����n�T�nC���F��(��,��M3\�J�V�K�B��9S2�Vw^�i;�H-�3�S�^�۬��^Ӹ��W���`��٥Jm`ǗhX���z�뛏-�w��V:n[��d�
o�n%�v
Z��c
N�P����lG&SLNMӂ���P�D:�]�r9�;Z�[��l�du�2{u﵋B�n��JsX�y�՘m?�!�m�anL���UMݷgiliT#f�yTE� �/+C��]bڏswQ��bII�V�omGB:��Fi�Mjص�Ef*ON��+C�)9(do�*FU�T[�6Cj4���f(�UJ��Q����V� ��%kƦ-�;�����N`�)��p��Q�ü�,�����1��8��)�U5�%�ي�nǪ����˂� 첞��L�M�D6sQ5�k���F��e�b����̅�(l�umF�n�{[NI����D�Α�d�C%���ȹY�3n����j!�b�f����^�2@�н	;��E��+ W��l�f% {%������sx���5f?��W����4Yxm���j�%B��Q�6l�Go$����Mhn��U�#R`����L�j������Ș�3	en̼lPh}�@QF�@�6�X�Y��`h����[̫p<�E� t�dّM���8�:[�r���A���Q��$�I�1I����HH�GI{�LB�b�!"7/5�l�$�:��6�H/6g�2Tt�jXk�Z�;�H�ḏ�����e�ux ��\o���\�q&�#B�L�ڽ��Y���Y9��Y�˼�6�2Q��2bfcWN⼫,]�&җd�˲#��,�L�y�C�^���Miц3�i�cCyč�sD���,̍�յj-�EX͖���su��j��ZEdW�:B�Bکj��-�.��D��Ln�Q!uwo]�# �k�WpZu����2��wX��+Z��gf� �+/H��*���7���%�3B.^VLp�L!)&���K�l��Z���L�u�m*9����p4�xv�me@n����w��,:�~ʵ�E%5����ڰ&n	�8�	oӺd�`V�jҲvSpԚ���)7w[e�!E[mB�ڟYR�7�Y��f�c�eXW��ɲ�[��<;� nd�а�wR�fH7�o6��4��#����ӊ5th����Ò�+1�i*�&Ŏ�z.�X�K�R�wv�a��Лy5�5�p�`���E����>w�N�6q[�2�̽��(6�	`OKF򶴧����I��DwYj�Y��		f�o[�:ˉPI$�,�wY�i�7A̦N��*3ۗ0�'�]���)V���̴���l ķW[7i^<A�ۂ9�˺W.��V^�¡f�8�N�׫�bO��2����OHd��u�k%<r�:d_i̺%��q,�q�6��cw.b������.c�8�hy��OY�
̴T��V\M�Ɓ2Vf�M�e�&�YM�5�Kpb`k١����Ӏ�f�H��)HDLV�=��D��mFfn�gs\M,�V3C�b��1� S���݂V`�Xf!"��Lͭ'P��Ҩku��)9�B5��"Yy3'�S�����wIc�����C�+�[�	E�i9�k0k�khfV�LMyH�d��>jКFZ���P��<�aU��ē�f=(�J��m:R#!*�5cI5�9�m$�qg4k)u.z[��]��D�Lj�B���2dU6Zv�%-3�bH��
���t!zb@	"��"�����6ŉH��Lתe�y&5�7#ҠnLy��Cyo�����F�妮|��5<u��'A+�v̶���i�0�+��K�k�(+���Dmc4�G1�b�f��d�n�)I�fZ�t�08�,�$��n�״�P(®#v����n��ݤ����6��[�L\��M�Ʈ�Cj=�(�7����Kj\r�������
d�I+e�]��E`�9L;�и�q^]��~&�٤b�MԚq�w�`�����rմ�����V:Śd�"զ���$�ˡ�@Z����y�Q������9��+0��S@�;sKlecV�p����vR���LY�(��;�.�g6A�� �wm;���e���O����CF���fe]���.�-�w�jn��m\���Ç%cj�͛�����Jb��W��5Ū�-�R���%�
����R�i�B�kr�ݡ��6�h�t)�e�6,Ð��%&쿅`�1�nAnl�Bmĳ%�CM�����(��:��6S��M��(j�`�ѧrk���%VÉ){OW�ַ>e����
�#��3�6;�.*T�
�rZ��D�q6��M��ۡ��u_�ig�v���zSjn�ku����B��1���b3,=��e�n*Ҩ�7{��~˂0��Z��"���]�Z;�?#5ʋ�U��/�����5XmF4�2��%L!o[(昵CC�@��\3S݌����)��͏k-�p�{I�!R��h6�t;�$�Im64�jL�������Jf�j��j�dt*�V�h+�%\a��d��	r �:(nCM ����)�Vu	��O2Պ�X��u�j7��jVeK��n�۰���XE8_^ܠ�liv� Q�R+�͓6��HE��of�9�$���+#�25�]-B�L�s$+%�#JA�Ci�:�fVJu��^U����F��dh��&���
���7S@�����p�J۹�x���@Z�T8��>�*��՟�ԥ�	g��Lc1dǒe�/VAm�N�����(h��Lŕ��Q_Kh"C3d��,�ة0��ӂ��P�.#b6����N��JEk�t�Qnѻ�"cv��R+�W��S��K�[w.�P����&�y1�ic	�j^]'��	twHj�ɭ`��.5iؼ���i*su��ҍi�T��]�X�?z�m�cZ�f�_L(ΰ��:��S�(�����A4Rт�Mdaۚoh����֋�m«�kCQ��[Q�E�&,����NFS�O��n<�`� �-iR��qA`f��n���s���y��5�4�e�W�\���eB֝�s5�{M��%��A(U×���0�B$/f�H'L���V�1�y��q�p�I��lHsS3)��$�՛/�Y���$u�A�B�%A6%��3�ݚf�����6�X�)Qm$��Ǥ�t�;�,|�Mp|v�Gi<��e�u,⬀�僰%�|D���yCWz�J,}�S�^^��$`K�k
"�S��ӹd�z��"��G*�47�2�ۅ<F�M�H��2�����&c-<���mbzj�9����!��٩��`��v�$3�*(v�7v^;�]�6ŀ�j%�N��ar&d,��on���)�\���d��������nC/o-�d�I08e�Z��b�ղ��)�Z6Eȇ{eD�%M6���W�XfiV���W���C���_l�-�K�E-�f����˩W�I)yi-��5C��0�nQV�=��P�&�㎶���]-�iջ�*����b.VdNQ�5�u'&�RY�5��jv�H&��nV^zf�6�YQ��I��3��zN8h�Bn��P�л���VViU�{�%:v����e�;�EkL�r��zh�H�5�z7\to?���(����w���+�{�JHd�Bʕ1ּjV8���%0�]"�{�tnK�{A:�Y@�6��[V���O�T�(��C�E�7������1-1t���K�e�Nb�4���Җ���ݷ���Cu����,�k������ȡX禎�,=��y˵�U�=גq�:�ٙ�A�`:�5���O0+ķ�4��Ã�k��l;�Dn�I�!�.�t�.�lk�+����4j;(�9DV���;����8f�V��V�Il!*Q���ÂV4�+/y��G gW:t��V ����9�|�a�XN��^N�6:V�X���Ptzk��n�s1]���ۤ5����f�rT��bB�Lc
O�Ì-���r���%����-F��)��z�N���*�K�l9��t��=ϴ]a�RF�:9��u�Ý��q7�m�V��6�]��K�Ϊ�R�u������>�\��o�s%mq�ϊ��^��I��XI^9-Ve�>���P.���U��L#�n�[�lJ�"�*�=IS�m�8=�,�C!)��Hӧ����:6��u������p�����A����)u!��C�o\�$NN�O��=v��#���Bj��N���m+��ܫ�6q�Wi: �/E��Y�DeJ�2��.L@���+h��![��J���w-��\�С��˦��u��,Y�Q����1=�=|�K���ɵ�@B>R�=���z�f�k��^Y�Kt���Hu� ��-}���]5�H2�����8ˬ�ѷN3n�0in�U�;�uh�g$�M����@v7/��G{��*��\dV�LC���k0�|�z�q㊍�V�D��Y�)k��G%�j�;g#�{�(k�2�Čɛ�`ý�����MF��,6�c�O��	�̵9;Ŭ���v���s���%�����E).���K��8��j*�F�BsQ-2�6�jB�7ݷl�M.�b�V� ���9�R��쮗�BL���I�Ur�#{SNB�lT��4�ɖ8�I\��L9N!i;9 ���*J��́�m�:����D	��b��	V�3k��|�\���>����o
�b5�`�ǀ��)����u�������#V����6�t�!�Ҟ��1*a)��t�����V&��O*�F���5&�gz���6)%	ר���iɝ��% �[Ua�c�s[̺������*�������|MuJ�7�.rK�k\%�l#3&��20��w2����0�zd��3s���=,�Q#���WV��صfm��I�4Id�-|��`<�+]�5ζ��넹�Z˾|e������]��D��)B���u��>�L�ʈ��,AR�l�r���ςz�fj�9�A^ImEǢ82�V�1(��a
�{�l���9�BES�	J�}2V��}�ԩ�*<�Cq��o���C\L����.�#%n5��Y�^Gֆ��­VPB7ҹ[\�1�1����뭬ض�hi���-��r ��e�t:�%��G�J���G0��v1����:������s�>�z�ס4e����ɻE�}Y�R�\&1̷�N�f=ـ�gC{��
���}CS��dV��WԱ��(аԚ�-Bj7|�aym+�1:1V̳x-qH��t��S8ڷ��7eC}]�S�;!��4nҾ"�m9ҹ��F����aʺY[�0��T����x/�h�	�:k��ȵH�o�>+ph��va��{�X�^��w�t��.�ժ�Է�K}M\��]u\��7���d��7%�17���,�ss�l��q$	˻FU�h����5%���\�qہ�%�x���v����$b�y��nʹn1����xg��0��p�B�*�N�cʹa��As��mVJ����l�[\�9�Vj�K�Gr�V����ݪM���m[U�,����E�f˜R�{y|eh8���`t��{]`U����(�AIJ}I��$�P�K�좒uy:֮�	�i�������sd�����&a%����m�t;���,t Kot�m��bf�d�'�����Kz��	����
]]���.阤�ʬӝEϗkz���o�Q���(���%]+5S�>���i^;����F��U�u�����l��(C�.��t�4���BHO7/���ƃ����
���7�`�&롤2��ɿJ�ĵP�%,����k��fK�ݨ:�(�k�퀲�H9��粶�i��s�AMi�tBŚ�īN,��_U��H;�C(�T�9�k�汵�*
�3	�����e-�JU�(}n�ɶ	��s؂��a��8u�%aV��m&��ݎ�,�<5ދP�ףz�C9�Is�$��;[���`U�:�������hmM����&�;]zb�5��F%#"�]���Vjî��#+�]`���P;ƺ�1 Z-�i���WW2�QR*\��S�Į_S�k>���v�I��v敆L�9�6V�5��Y�Q��fe^���hiO;����*n�����M6Z��c6t\Iogf:�:��ҷ�2�s��w:j*�I�d�sPK���	%�f�h������lu���ZUYF񋥪�YK>�
k�L�fW ������|�,0��sJ;gr�j���q��kG�w:�%#��w+��]�`��N���ig���n?������);cAx�'@�L�Ee5��SGs�ՁmV��h��2�u� �g!7il�.�k_e�Χ@��$b��ጛP�U!�C(q�x٧yáM$e���60��]�h�*����r�V���6�V���Ik�?
�X\hYm��m;�
�΂ר���B�7졄�}���*�s�G�������Ҳ@�,�|�|M�'a��T(���l��P��.S�v�Vbo ڲp��1�<��hv�e��K⹷��:I�����rl��ǰ@�/V��v�b�"���Z�����Jn�n�|
Y�%�Q%����1�z̄�.WB)d��y�f�iܡW�ג hQt�2�^���/8oTP�ڱ�K�;��v��n�EY\mruul����EӰ����rT[]��������c$���В�=�;2րv�-��D��M�Y��rnn}'[�୹(@G$���侦{��y%�+�eZu�L�願�j��"D+=�u6WTnEn��QoB�r5$kJ��뻙.,��/~q ���9���f�ۓ-UnD)�W	N�7&M�y����	4�XB�Lٽg	U�Mf�h�j0��(���T6��o�<c���5���L9����Hc���9�bGr�Te��dqNU�]OV����x�N�;Vi�0#&n_��&eu��W;d��av��УO[���3�1wV�>��"mU�	+.5�y��N�l9�째��!�TL�9\%������`�����q�0AIjR��V9#���n�D��t�sK�b)Č��#9i�pzf�+F�ȫ��b��}�����=C0֮�84���un��;5��K�h���h�]�1��M���@�0,Y{���AW��L@��s�,�DCwyئ�`��\��]�hܦ��ɮ���i����9�xq�cQq���yf�fD�i�љ>�D\n��p���oJj��jZ���_&�U�ᇥR��aj��� Ƿ: ���A�Kp'�*h��O�4>����-[��j�Y�}��ފww�_7G\mK7U���{2\@��R!��u�8��Z��)V�"�w5�
����K���Q�^�H^��]<n���L�`RO�je�x�S��8k��w�*�Nsj0���둣�!�h;q��u���KW��{{Ҵl���)�۵���3t����\��(Y�����^6(ֶ�b����Um8�Z�XTPͮ��ƌ�[�hè_ϥ��k6*�	�6��ҎL!ե��qDU��*��}�-C�ĳʹL.��*�ѷ��{��p���TU{�b�~�M�J>Y�O�Pͭ��l��^8�e�F*ɼ�
�H7Ǆټ�g9�tFg� V�{�H�ݫ�6�ݡk�Q�t��,}���ɧ�Z�bk�)l�zN�O��$9OWZ��}d��*@k|	w��2���(-`c��d+8��h�ɮ	 wm�C�t1�(eȘ����j�pU�R%����4����
���'z*X�$.JQ때Mu�!8�˫���mk�1���iXR��B�9V^�9�� 㕝wxk9��Q����--��*�_�)qޑ>����3skj���v����)
�0� �(�����k��SE���)�o�����GW}`^��CN�<�˧׮��&@�#b�V��=���#C���I��ה�WV*�ݗ�j;l�T��NQؖbu��nW@�:�e���0(cۅV�a��}6jy��0��zo�JOV����No3�ً�u�P��u<�햭wN#DZk��H^̙��]N���G:����֝s��\�Z�r���b�@�R$�����j��]=Y0��*�x�]Ws�#o���=��=t�Qm�nw���(�)�@�[�+rfPW�tp�9�kX+)���*��;���)��KM��×���v��H�+[���qОϺ�M��\��Yz6*��9����{�i��,	V��1:[̫��@�WL�BuA��=����5�a�0�l�;q;E�4!�dMi�3Q�Q��=ެڄ��6�J��y�d�8�Z#Red�VGF��q;s��x9v�hG� SF��[r����Zj��":�rf��H��̤K�Y��-�nE��	r�DƤu�V��9$�����x�\
�l�B���:�Y]�����[��2=�O2Z`J�F=OK��q�_4�T��q���8����wU�U��W6P��kq�Klfԛ��K��4�qh���Q�Pv����ܰqT�A��r�֛�[��M�u���*֙�#4�z�2��Ҝy�V�}�З��S(��sY����GP\�!Q��T^�4 6�,Fж�bLծãr��r��}GEt<Rt���n��]�F��sXӻ��f��C�]q�J�\q
W+�T�(,
���e�=�/��}�rl<��p����p{��jaR[�
��i�U�>�{�_��.$�=���p+��ҫl�:�m��<7}�-�ٲ�^J��s[ة���@�
̚�7 [����1i�(ʰ�g0��Mp�h1mT{w��u�I ��[�3��c��y�����v�W@\՜�Bx20�u���윮��m'�]�����i���+�l#Mr5���hԕ�l0Ĥ��vG2,��	lZ����lG�*�G��L���rT�����v$M�qX�n�Ʊ��9)Q��F����^Tٳ��Һ5�[�KOr(��E܍wi�]�4И�d�֜���2����G�(c��Kvb�;����9�\�Wp�1��u[�F�ީ�Mփ�	�+f-����3*�ʝ_6�+Ǧ�@�f�׵�.�uьVL�5��c��Q��$�q�+��F�{K&��\����J+�U�t�m��bʾ<r��R�iST�C�j,�{]r�Q�X��X�R�� �:��)Iot����$�����6�:f)Q/J�Ρ*�7�L=�(���Žz�Ṁea��ѽ����J�a@��7X��B��������MX\�,&�)�����t3xȨX?���\Cҏ��H�9ԃ��c7�����	�5]q�P4�V��2�ؘ5�ψP�s9De�ڡ��:c�%wY�om�9Z�yǶ�U8�wl�[��\yO�t����'��뵬�2:0�K�KL�����ͮ�݇�"@SS2S¡�����Ω�N�s$�;�(j�v���u�"��e���Uf٤q*���Πu��&�J ��F�g_=���`��*f�}��A�����;Z�WU�>l��f��OO^����|��8�ː㔦�wʈX���\�W�N��m�ʣr%},19�I�4Mʼ��n�.�� �x
GXwjl[��M��N�́ޤ���=����ʾ���ҭ�8qn=�0)���ݧgoM�h�	�� ��ڻ�4û�QcE�k�-f�w�k�����X�E�a����� m���F�^��yS�U��w�+rM�k�dV���_W:�'@:�,�agж��k���F&� �R�tۣ�b�TT-��W��I)X�h�B=Ccŏ�j��Vi�tz<A�E�^�f�Y%OR�u��XVL釀.�n+$��klQ�sh��.JG�o�����D�*��X�W�u�cr�4L�i���w2���y��b��M$�6sI��闘�4 ����.��wOe����Q+&����h �]�1Wep4zd�	�s���VJ����Cj��ܑM����eo
Ӝ��{v���u>����xd�y;T�N�wjɨ�Ĥћ�7QG��%�Κ3OE�Ül�����4�sb�޽�nkk�9�x��w� �4Ȉ!�w��n%A�a�h��^%�6�Ƞ岭����<�T�j^:����<�$�
0�L>�kZ�kb��B	�y�e�/*D6��Œ�ۯ*�M�j��H8��e�@�5k�i��I��h{Z�A�L<�]�vo�ښ��*;�OG�s�r�K܅NO+t۽����wc�A��B4o#s��rT��^�ȍi�4ޣ��=�l01��d��m��
�����P�����.��x��A,,C�Ͳ&^��E�g��k�v�$�7 ���T}c��Gr� rl�A��K(�Vގ�c�J��1j���U�3jWw�X$h���W�&W1PK�e`���g
��:G�"_u�sI�KP=�
R}���v�������B��5�����V�,pќ�v.�(<j�^�H�5:Xc�-��eL
�ڹ�R0������ *��qK�hId��\�t�A�9�E� \h��}�9b'.ksC������`�33a�0�i{^��v���݋�z�n�M���8wb�¶��tM�V����3�{ҭۦK���qT�3V�pRIl���:��R����!�0�U4K㖔�eeNh�Ԟ�YRbP��<�x�͖rU�� *-91r��ME�:��av�5�5QBuF�k�u�͍�ͩ���gv���jDRvŇyR'���ů�b{m�Va��.5H�PG\YV��h5ܲ���M}hQ�sk4=��;������R��KUƌ$)�SX��3�:�:�*
ڝ1�N�{�-я`N�k��6xm&z�i�V^��3�đ�`f�Ɍe��i��0T�UN��n���wV�^��#e�������ܴiƲ����j�PFoK�d�G�8	�[�CYv�r�ݻ��t;ϊ=��>O��-2�1��%��^<͝ɭt3����"���T�36Kk�D���=���q��q� y �R.�r�2�=z5��YoE+9�k�X��h��Y�l����ZZ��-a�O�C]t�P��W�^Hq2����CT��9f�腵%���:=�fv>�W%�6��5��T�Y��z~6�(6>]�&���F�?���S"/5������9=7��p���nv�^���z$��� �C�I\��T .T����k��T�n�5��b��f���%B��B��*�G���DjaD:Y)�Y�u5|Гe��462���ȋ����ѭr�]qR�>����Y�1I���V6wiMfQ�k�J �k31b�B���6����-G�˴V��̷�����qb���9(RN�37��WYWWz^D�D��لˤ�^�	si�XyV�ɹ��^w\��p��9,k_��9ٓ�Bl`б3�<AvL�e_W[�Gi�L���(V�������k�[N���	)DD�����6����A�ʏ9�*��U�oA�1}�C��Ĕ/�8�.�ik!��boM��G�cyQ�k�ju-)�m\�l�̭�Z��Jq�R�M]1i(iOAޤ�*���1nb�-Ql�OB��4�;�������d3�N���u26$�s(�@��WZ֣t�ú���U\����D&�4,((He���	ֱougw���fŕ����8tM�?��72�dաٔ�N��<�N����ս!C��r�h5q��Se�9�ԫ$���r�i]��{���������,�-nK�^��䩍�Z%�s[�2>d՜a��a_cH47��M>l�Q7����ORԪ�C��1�����<s&�{�ֆe�M�w�I��pj���Ta:�c2���(]���f�.b)E�5�?J�ۺx�tĻ̽�)��v����9�ˁ�r�Kz���ͫ\v��WL�#6�h�*��Ov�nfGJ�!<�T���9<.�:���m�A֥�*4���[�O�`a�}�̽M�w��}�*cl�NG�&��9�;:-�0�+r^0�xjd�Ep
����̈́��ݷ'Q[�����C7�J���м�%g1��( �
�𠦴�Y]�(�vW�7�T�r}\if�F&��)�k�9�Ъ�,,^�J˙2��4T�_�a�6�JC�XZܭ[jF�ri^]�C6
l�U�R���GzU�Uu�,_Z��t=��
�"մ��YY�	{%5 ��R!b�Wrw�v]g
·熵��i<��^�y�3�-�4�vDɏ�9�V[����u�'�"�\��M}���q�'��R�Ft\ҭ�,�QQ�Z���.�o7�[�X��;*W"!G�ci�T\;͉�-
]A�G\5�u�x��1AŲu�Xnu��K#|�3F�@u�_B��G�i�u�p6�"B���\��/E�Ӑٸ��q]�퇜i6ڬVh]]�c�	άdb�mG�Δ!�[QD��	���3�N�r��V^�^�[uͪ�P���#��>D�5����P?�Fu24�o|G3���!�nJ�Ӊ�zj�	 B��� V�LmV��H��U9�0 VJ�k%�XU�ۙlr��{8��c`�[:�����M[�4��WSCy��f���;Ҕ�r@���P��)-"�{0Mp��:�8�T(�����{IO��N��;WJ{�jI�$�+d\�w�if3f�<7��D��3Si�h]p�92W `��X`=a;#�D����}Gr|����S8��z//'s-�tYo�p�%t��6jQ�y3t"�ڢ;��z�@�h�n�B�hK�z�ɤ4��k�hn�P�{2����,\,���bY��LZ���	Y�]��C�\�ظA}�^�er�yZr
c�1�B�P���95����Y|����`�y�{�R;P�Vh�V�r�A���;�gUݼ졚��7L|�8M2���5�;���ӌ�{2�Y�ٚF���32��e��H�Ϸ�ؙ�8�FX��J_>ݹ�Į�T)R9w�����Ǘ��z��S(NU���;����)rJ ���C��1�]�c�v�jUñ���r�Cy�5 ���'Y�1�국Բ�]����� en<p�5ڋ)eR�U��re4(�Ց-z���
���s�%i�st�ghϭF�!M�ˎU�Ү_95����%X�����pbͦ�M�:�s4�����Ʈ�swZ��	���o����e64Yޭ��-�t�R�ì=3�A&N�a���]�-rB26�ͮ�*���^��r���7j����fI�]�&��h|bp�f���|�WC�[k��OmN{u0�����6�PK0:�X���s:��WPc'=G���I\D���}l>�]|2��]y�Vwd�5����um.� w[��u�k�ӎ��Q�X](�Y�ao@i����<һ�W�#�£���șD,���B43L���Mf��qV'KS@�	�k����YЪ]9h[��u�&p,jjL��:n��F��5;i���K#F[6)��wS&�XA�����N�W�w������ ��*U�ˠ���g����;<��4�L$<a����K(RR�nk8�܊d�WG�T7&vm�Df����wi0\ƥ�S�@��l�Ěp�l��U�ʽ!}ɥ���n��ZaMY0H�&�W�˗���P�kh�΁��ՔrѶ�� ��$�(]��q\�\�-�sc�*7�Wo^�<�V3��Xs&��	$���H�6��y�m:�B{OA���;m��NA�q��Eg|�l�}ҁ���,�駘`@6����'vd�vu�A��w1�g��Rl�E;���C�(i<;pn������6�*��9�ì��὘n�K�������K"6y5�s�9rԫ�*0�혇LՉ+�I��^)�nj�F�i#m��:2[�hMװv��a9�q/�r����_g*[I����Ვ�-�!�X��+��['�M�d�ա�٦і��Z�*����Y�Kˡ�m6��-n\R1�tJ���9p���ϲv	I����['%�:v2���U����g��WR��Y����l�a۵�^�f�3E�(��B��jAi��H-��0j�����T%\�G�nSy�`���V���,.��L�}ԙk��r�Wђ�5�<]�O��F驠�_<U(YY\����Ť��i��]j��z�*cY�s��w�{d��*ٶ��t��9E2�96��{��2�m���� 1�f�'oc.��*=�� ]���c.q�d�hfv�������;���9j�v��X���W.�2�� �8��Ż�^�-�}0uq��:�
k����]�|zL�PZ[u:�M0l%v/��n�\.�
ޡ��w�*�t�V,%��ѥ��iU�5�̾y��+����)kY�R��˶��* ����iCז�<6E�,��YSy;���;�q3����4Q���K�m3��ɵY�}�4�{�q�r6Fhuݠ�n��7h&�n�Y�y%j�H�ehi��[�y���,ܱJ����;1��RW!�=�DsT���{�-�|�����sV�rL�ޚ"�5Ƅ���i��C�ÛMK]1�T5�!U�a�����v�MNƏ��n�ݮ+�GF�oc� [�f@��ޅ���|�e��ח�V*ֵ��\+�X�|%Lb�B�� Gg�-Su����ƚLM��1W����}�-��Oe��Y+�޾��ae*8���tU���Bng�,:U����E����6!�P-�&f<�#v�CB\b�z	w������D�)-j�j�^V�ԟE�J�� M��5�^�p%Xz�g.�Ev��S�V@dZ��v�S�x[weX������ذ#>`L�T/d*M*G!��X]���:��vԑ]�Rѝfq��m��&ee��T�S�k��S�m�+3�FQh�U�3wA_�_���ef��=b/����HAE�X�QYL;/(>��-"���n�յ�0��]t9�N����L�1�\y��<q�[���᠈8�᧺t�[�7{p*n#�N�F�>[�x�[!f7�i嗶Q=�elM���t�驫�O��0S�����-�֌�0B��`���F(!62�q�=��W;;{��4��J-6K�ka�r��T�6�t��$Oo=$����?��g)r1N�,�úk��G���E԰b�/WJ�`����rT�יb�gMv�����j��h���9����wy��1d�WW���Ȏ3�nWeiԳm�2$�p3�\���Q�j��x�<��樭��k{nL���n�-�(��.ݘ�3r9ٓ��k�[*v�+�	|�%�-U���tq �5��p�����"�>jk0`o��s*�>�W+�hd3��;�^SC��Gn�QoV�M[�t�Ckq^�W	C�71��,���p=71w1����/L����i���ɗ��ngK��ff,�\s�ˤ���VJ�@)2�V=��v�P�Xq��ʁ�5%�7�OB�՜��*U�7�%E)P��P��B��ٸ|y�;c���6��:�R��V)e3�L\���݉��C��m���/u�8��s��e]�k�uX�n��M+,NX4��j��r�_"*+S]����t��Ù�N5����w_Ri�ڵ�Y�:��� ������ܱ���Z^�^1�H�PS��ke��������ǥ��*�c���-(u�+��|�Hj�����QI�b��+s)���>q��f����ͥ�ͣ�S����d����M��ڄfY�"V�s<r^୒�C�y�%U�Ԫ�8mmp�Y��h%�
4����2HI]�*�On�¶�tw��M�V�W��]����L)��&s�+��$`��[�u����NB�w�}ǂS{�8�G�Q��Ǣ&L�A76^Q�����������R��s.�(�a�f^��#G]i*3�Ԥ���ӫ`b�m�Ps���Z�่�D�R}w6��XR���voq^����&L)��=tf�넷|9U�S�w��y��a`v��%����jiF�L4��갑ݛ�&���f�՜r/�Z���X ��Wϒ�f_�ռe���y�u�-��ɺ�,�pd��ts�Q�)R�4,���wBfs�3Ho��SS�ˬ�ʣ���qP=�,v��A�PmHu̱����m����GrD���WAbZ47kU��]�T�
�g��֦��S���]N�]�\p+��NmA��F�4���)�E4Q����.x,<ِ^�-�R�m!��M�8��~�`L�7�K��{]�;-�i���ȅ
w�˖6<q�o��Y
��̎=�ֲw,Ȋr�<B]_R"wWJͩ�b��I��㉻y���p-G��X��l �6�{J��Ʈ��W�S��Z��v�.���9�����m�ۑm�b���f9q㥶���r*�{bٲ�<��r��8B��u���
�Zr�*��oJ͗w1S���)�/t��OC+�!��ʁK�� �M˧B�!v���̡�Ak5^�gID(E�mu�7�T����6j���d;�Z!�Ζ�ځgR�O��l�pi�,�_ag�˱��X͓DP��tj��u�yt� -���o�S�5�u�h�ӷ!�P�'��G�p�f�6j�YE�o����)ͼ����t�Q!.gK�sk�j���[��֬!�h�2�Ȍ�����]��^��i�n��ٰ���N�݂X�+�js��z浏�+�::|0�#Qū��{2qbgC��[�(Fm56�*�[�47�r ��5{`YyX�5�qN��5t��ݦ��e���z��
5��ާǓl�+j�[��p'�O���r�k�yu�M����U�uQ��u^��-��]wn�����Fl���p0�9�L./r/� �ۨ�2�٠s-=����넢�]�N�q��o1���l����:�4�ɚ��IN{�!2��;+%gL�'j�z� �P�1�&Ӻ�7՝Wq�_f��J�vA�KW���(��zt�Tۣ����ڂŹ$����@�37]�]����}�C��E:�lQ{�&�s:S��1�̱��t4��#[{.��F�u�Ʉ�XGEi�Y�^øC�7 �]̰��/��)��ᢺ:y�ݻ��X�*���l n^���*�޼QRF.*�ɣ8����X�c/�!�ʾk�l5�<u�M�4�(YT�_[�D�LE����sg>�sp�S��
�s��X��L��Ljv��1<��Y���Q[����	}�%�u�e>�W)v]�yS�-ʇF�X�R݊���e�Q�GH2䨔
\�a�iL�r�C�=����q��t��ʋ�en;�Rq��T;tC�Ȭ+�r�2f��k-rV��; r�02���ě�^�3�`��[fԍE���Z�B	6�*��<��Ώ+ueCk#S��o��;x���Q`X"���P+Y�6(+{��S+�XWq����CG���k�3�����Qp�S���j��{��ʹ6tI�� �f�n�Z'�^Y筡�^���y�_[�#��ߍ��֖���0�ii��{����q�wK�xM�$�N�*�'�̮̘���g�����;�-��t�_-��4������P�+�<@t�D5n�z��Au��q�������I�6RT�OgE��qK�+��JJ�v�@�\�jl[|�K���I-цaj��fr}(�#D'";�.vX*+��wN��]��;Q�|����s�i0�$�۫F���l�7mٓTcp�,#w*�G�m�/���E�:H�;:x�X���f�`9n�k�,��®3��Z��̺s���&0�&��Z�=��cB���_9X�hT�6��;f+���OA��Zӊ�ܧn�)��j]b�LV�=cz��q�O	痸2���΋]�U2���[�p��٥���j`�$�ZŽ��;ᑧ(�SpV����i��ŵw��5w��t;D�e�R@7�&�t�qɄ���Q�-Х\/����z�c�b��c��^B:�Ǌ�N���H���u�1�v���=P�ȈAm�j �K�	գ��w&M�9�Ym�&�1ۮ�)�K�^t|W��nS3�+��4����G`a��	NW`=��2���V��nE�1m�D��.7aJ�8�z8�N��:�����V�\ ��d#oLsr]����J�����S�����=w�\e�3{�s�eg����N�{�<s���J�t�r���Q�dIZ����Us�qG]�Zy�å�*snU8:�.��J���ndh�����]�-qs]ݮ��;��J��\s�����S�y�����mwv'/#�W�#�S�{�8��HI븺�^y�Q�����By�rw0�8u��M�uZz�����]����n�p)uː\(�9����Q��u�˹���(����$�g$wC��9N뫐.��G�y'�Ƞ�P���#РN��2�2��.E���z��a��N�]K�w吡�:��t�=̠9��	�D%Ҫ��=�@����=-��P�2*��Vl�Ť��7��<��q=,��S����1u�h���;I�Ҋ���.�r�';�#�g��DB���B�rWq���=��.֎��Fݓ���IST�0���pD�Z�+T�k�{����鮫{�b�m�(S|�.&��ͩ�8��[��q�sh����x#���*Mv<ÿS5��̺��l��	T/�VG��%
��W+��'�C�ݞ9��d}j/���F"�=�]��<*Ų�a-vJ��͓We�,�^i]΀t� k?e�݋��(�p�Zᮄ_q,x9�;:�2[��z���oW��=I���^B_On�}�c4���(سQ�Pa#'G�O���`}8p��ṣ�:x��(���!ӨbU^��O��+�sU]�7[�d��GX�z�*�G�S�U��zB��a�&��3#>V��/�uM��W_n�GET����Gmoq�����fg p�ixێF��*�S��=2�4{�t�M�l<�#�����ͪ��K+xhމM֢�Lq&�|�LcS&����xL_r�Y]=,��K��[*/�]kPq����A�z�Qo���#\�t�	�>��R��-�,��ʤ��-���M-/'[4�	q���r9He��!��p��h����]$�'��|R��b��N���=��m�V�c�|�0�ֽ�%hv�!<�z�`A���ۀ�
�&i�R��X�|�����Ӆ�Me���]��+�u��r��A��|ĲԺQ�MZ�53)���C.r��#��(��rw�F�9q�Ra�E�E\�F��%聭#V��C�O�7���n�5���=���CL<�*�Q��������o��6�NN�ۉ��D�!�\�s���놌���p졹�u�M�u��x|�����l��v��GK^���U��T@�LL�]G����3�ڮ�\��2 �H���ńHw���gg�7j�҅��5�=7�+�(��}�F�2��Q���H��+���֍F_�T9!�F��˕MTR�f��'3�X���/��G�P�?mP#�Y��V�oCOeҙ��el�מ��J2��:���M�t6�8�g���u��M�I&@Ӑ�D��{s�և�V���Q���^�]!�ԅ���i�w�"wh�>�����Bv�w,��S3��ߦ{c�kPD�?1�Jޞ�tD��	�UϯI�U��y�c��9�g��(*uz?��vs����O9�r�MZA�쫄���*CZ����7����Z Wێ��E�Fm:�bښ�����s�Ws�EO���E��'v�����\� Jd�����sU�)u�׍���{�D��΃�V�P�{Ҵ���s���>�듵�64��Oee��GW��ín�����Ɖ��'IAn��;��o�s���<�;u��4�"��t��h��W4�z�o���[�++������&Y��殬��};�?�j�M��[g<QC��8�CuEe�O:�;�1.@V!��=ɇ��EG�y�)��8Kݕ������xFfê���pe�$Ң`�	h�zߒ�W[f�X噅w�
�"�W���`�+�r�N�}�b����}JH:
m���'^D�-{��$�6�,k��Á�E)��S�>�P�`q�ڸ}�q��P��Jׂ�_q]n�����x+$�3�O�NdY醍⺂�"��.%�.9�4c5�ì�6oYf����jo�V��˽�:C^p9���&@$s+3����Ė�8w�]��2�'��Qj,����8,�����F.�@B&�A����ؒ#8�b�_!Nv�j���_�2�%�����9/~�:�V(��x����l� �}�wF��ZN�|���z�[�O��*U�E��c*9��-��"�/`���W�*��9�]�Щ4�����	v�3s$<:;L^�ZoS���PB�ޒ����uS�����I�W�H�z�!T��`�-�r��q�v���,&Z*o���B�>}:��ˍ��"T�����B7�ޭ�8�Wjڂ�5�oD�м&�(*r�ǜ�F�2�t�����,��{C�˔�Q��L#Q�EnȰe)���
|e>.�$�\����蛆v��I��?w�,�C��4dN�zo�6�U��\$��\"�S<�ȑ�l}w|B�wz�Z�p�6��u��Hb�y�1W��[�旞aιB��cE���b�U1������CE�Ͳ-��!�TC����s#��;�
���h�Ʀ4F�_n�[	�4!fd^��QX�):�wL�����L'���o�D=>��̪?�T�Æ���y9��jnP�\N$�v!�s�L�<O"+M�v�d�EYN:H�Y�hԁ� ���l�W���q4�j�8ƕ�6] �L�Q�S,�t��<c3y�4��`�
�^�3�:t��o�N�o��E���[J�Y]XY���Z�(GCr��w\��0B��,kI�d�ީyJ�s��30g�	ٞ�=�Y��J�B��`Z�a��B٧X���U�K�^v��Oډ�������u00���wAZ�;[�"8�=��-S�J��L֒�
��ԁ�c3$�����ۮo�t&:����@*<�¯ჸ��bi�����De��J�fq)��l�t�A���輻���x��a���j܎Դr��u87t�ʿrL�sX�d#!���=��	z}�6�]J�S�o&�m̴:\��ʌN�}��{ҁ��&T�Kԭv�ǉ6�[6�n(�����/��jz��g5�V�RfC՞��i��^�!�"5�"��g�d���䋉I��9����u�&i��f
�ќkWȉN�0iH��0CF)�di'|������yn�?
�����茋�YJ�4.�C������u��Ֆp��J�_AR�@�Q����UjU��8� ɺ&���N�����k�i^�A�U!��O�ҦKϙ�;Z�sW��`�U5�+�Za ���%�#��sK���c'2��/�=�1��������c�Lo}���=W���t�,y���^'h}�a��w�{�S����{�h��v�
�E�O�0�v^���W|W9�Kg��
�o!/�\5���I�	n����]�[u����n�����o��_�L=('3���&��(K����! ��R��t��꽯Men����ԛ�?XP�9y��Ʊ�2:�"�\�:������+v�e&�����z��ث�6+��וzs�N�b�1?_:�d*N��G+��Knh���SA���ħ���[w�G�Au�L�5㱮��v���s;M%\�Z.�;�>
�Gg줮�-F<Ք]�4g!k�w}��t�cb�f��Ӄ3���3��R�6;�ȒpĤ�!��qCj��"UD�jB�ɵ#�L\o5�~��e��;�Y<�6�P7�AA�u;��.�}x[$W֥7<S��hJ�ьڭh���q�+}����%'nZBO��N��es���^'��/;��'
������;[L��j����^;��Gܼ2RǢX6M*��']%�*�����c���c�hm7�\�B`��Ƅ�T��!�����<�.	�U�6� 1$���F	�eF�����M�2�d�?_�걜���<,s�]��!�_���U�\*?�F7.`��yO$���qIZ]0 �$90�"��jw`)�����ڿ���eϓ��[�6c2���@��C��
<�
�Kuq�ـʀ��:Ls�z�px�*�W��ɪAAn�0�Eڣ���������[#��ݜ���(���#IVˣ<T��?zנ�>$"�mv���4�kT�6����U���:`ؘU*L�t�~_;Ř�Uk��0���_1�r��:˞�����<�o����\Bj�E,�dѶ���P�1d��zjJ_@b�F6/I���
�9��Թ�֓����֦�	���K�'x�@�ȩ���0x�^����N'��{dK[.��b�*��WB�L\�u� ��!)h��!6�l	��n�s���7!ʔ8ә�ERc�'����4�N�vn��2��be1M��Z�)�r��h�Չ�,�����S��0�������}���dY�o�9R�M_���&��*�^{��:({�<Ltn��١����>�����|r��Ŋ�Nϐȍ�/.L�;E��9����d5�]װ�x`1�| ��^�U�A���^�n�4�7f+U���n���V��ӳ����F�Tᥪ��{*4S%tIi����߹:�*;�I�/)p���k�MwF�X.�(�!��8�CtV]k��͢�Z�h����}�"�/�&y���5�<l�3cx�[uKs�ю.�r�7�_"M��%��+3ٚ�L>�oo����·�R#��Dit�U��9l�7OK\�!YǷ �����o`ԏ.�t��⓲j�A
���f�&2̣}��\k�Hc0�m\>�8���y�O	[%���k���`�N3(	�L����F�]Ar���.X�|���!�"�~����Z��7�,����C�'M3�����d��v�ϝ�嵞���4��M�����T!��]7�06�/g�^]�rV���N�r�/1p���%� \dA�x�>�����̹7���+ܖ�oL�];w�����j:J�@Nn���mU�[���I�˭|�9;O%4�c9ʴ�{�܄T��_'��KO���;���شi<(��|$��@�c�R�����~�#8ӣ/����0�T�����Q�}ʹ��6r��o��\�QU��k������
{��$1�o}Z���n�}H8=H0+��[�m�p�.�d�6���̊F�31�&:�����-�3H��gKi
�V�!"������Zn5:���1Q�;4o��#]¬v]�&�iJ��JJ`wؽݢ2g�y}�@�5r�]`�,T��G�C���6wt/�X
g�:�!Ց9vsB���k��B?�z�A���z�Wk0�iz�3�k�{�o���.n���wK�\�[5�j�H<qH5���]X:_Ao[B�V'bx��4�.Ӏ�S�VF��*p�+�!��VJ�G6sDsˈN�h�S~���0E.������鬻�}�h�!�MNZq�<�r����U�-�~����h"+M�v�d�EYN:H�C:�K��}�Rm���<�|Z�R��u'����4�%9.�w�a���)�;��ޚ����WаaIl^*R��A�^ńn)#�ƅ�VÇx��],�Б�#�!J��\����k���wr�x�biI,t�AX�Ś�G�fesb�j�LZhd�ڎCC'Vp�z��;@B6�h��J��ɛ hLoL��;�Cb�nf�n�״t��3N�7Z:Q������,�tdp��t��.�-~��:B-�l�|�5�ي�+���|{��+XZ�N�c��Y�#fə�=H\V�t��6>U)]�\��q0�V��F�o7�zi�,�D~�B�����b &�`@~î�q�wm!y��D�}��ᶹ��{+TtYLJ�.
F��\@�cCo�o�`�c����@*<��BE&d��4ͨ-�(�G�Z��9K�%���˘c��CrDmCtE�9�T$]B	�h�����s�/.�U�p2Z(|�����òS��a7�#�ʰS�r�o�o�葞A�IY�]�O�P�.�%΋����B�������?er�a ڢ����J��}:�*�����]��}ڻm��	���Ep'��I����e�F&�R�֮C�O�)d��{\�p"u[��R[�� 訊P�:�;H������;U/+ֱ-�t�S���e|��<��m��dW!�W�\�	�,��v~Y=����ɱ����WJE��ldܻ�r�.r�*�!eeK
Y*t����&�|�]}�l�M"�`��F�h��	xU?L:m�TyqYGѬ�N�w�5{��u���Ԓǲ��9ֈ�ڨ�\�.�E �"�2�����<�br���Gt�9ڇ��dug��4�³A]EEȷ��ֹ@����+�n�B�@:SG��n�^�GF�W�g���i�Ks��b�<4D�ʝ�t����m��ʘzPϓ��SUQ:���4�X6kJ&1Pg#�L�<����w�1��c�j���%�N\gRq�`�CY�s[��ռ~n:�Bҁi��Q�K���0e|U@�T���K�zp�`x^�Us�x��ӿ�r��!��"��ty[�~Mt��ϡ\��ʝ4)q�����jMG�j�K��tal���.���Sd74�S�Y��e1p�1�u�mL��NG|A��X����ɯ���Z�x�v{�ή�q�Rӑ~ae���-Sntw|�$�L�& >�*e��j�v�r�w�8>ق��	�֭���!���Cju� R+~�l= %
���u;<��>b�859�n�G��U��Su����봎󑧬���Ge�;�f3��&�In6���0�QtDE�5�HSܷ~�S��Ƿ���i�7�Cyf�#�D؃���^_�y�dJi���{��G�dL�RVk�I���\Ȇ,˵[P�ƳW��_u9�3�a-�#���g�^�k���Qo�]�\#�A�6�7K�sTK[ݬs'�.iN�<�t���-*��&�⇟3���(܋���3t��'b�v�Z����R��e����ŷlnf��P����M�wd6�g���/*v���{L�-=�ea�*#��)�Q�]�ғ2ևps PB�g�*�^C(�u�=�:r�$�ՑvE�/��ni=9X�ȱ��њ^m��ou�>���[9uW�I�Rˣ�`�Ò�w���mCx>��5o�>1�}�0�N����n=�1+�/�0���2l�S�n�����C^�V'�q�\��=�p��I3Ze��t��+�ݓİސ��sÆ�0�:м�k^���VGZ�*h�-������z[b��k��w��s9��W��H���:t��gn����烈^�y���5�q���w@���NȠ�^�(+�X�邻�*�2�����벪�z�n�XU�v�ހ���(��d���Yo�f��z:���L��9�m^��}��gTT�RoN��b�4�I9b]oy�֓ۥ��ٶ/TnE�q�-ɇ+'ά�ҢK����W��L*k�Q-Ë"����f��{u�oOL�֥]���5�#�ݓ@VN�<%Z�+	{s/_Y�hm5�2;�W�-��/���WiH>K�]�;��U�n�,u����2�L����^�N���L�귁�nm��iv-5�\2s���r�6�n��4u*1$L����skq.��B�]S���¡�NWj�}��-F�,cQ�|���ڈE����+=S��,�yX��4%d#7�
�1�U�	�����o&d�t�G�g��ٕ/Vb|��{s��Q�r��%W\��ԇtʕ�Sv�nE�=�1��We���>$*Sަ$�
n��fv�p^eǔ{2v�trt��.PMqbd�u���PNQ��ᅳW�1�sz�{�yЉm6~���n\�[Z��1��&��U��.Qv�P�PfP�f��7���^���L�v��k�o��%�+ p���§Q��aŏ:j�Ef<���͕*��=KMq#k#��ʎ&
Q���,+�h�rյ�Q��� wHqL*��W�|���q�p��r�쒶�T,�]�HU�r 3�$�01I*��nVG����j
gm+�h��p�f3�[-�LҲl��L����5����r';�8�ܾQ|@!��*R��{DMZ0� d�9p�(b�T�NN
�E^Lk��bw�5�|b�z�F�h#��.v�9ۊ&r��aX����/4	mj�8��o�3b����
�f�N�,��&����U�K��Y\��5�����V�FV��W�>��3Z ������v���9���od��Ǎ��^�sj�$����J���dA-�Pɇ�_����ϔ�/��K�a�y�ss�!=��u�]r�sep�����Js�ttG2�w]uR��)L�F�vu��5��t�ӸNNb Y��9u�$�qE
�'5wD�3K�q��uf�qs����Țl"5�y.�;��:�xT�);�8�N�BjU�eEZ��:����* �!Pr[M�u�纺8TYS)Vd��^r�%�%*�N�ndY��y�99D@��Axt2(��z��䋎�98y�\�Y�ܯpp�< wR�NTS�I�C�E^Bd�Ⲫ㜼�d��y���=��H���9�+�<<�ۻ�Nn���r8t�5wk�����
�n\�*�.g�"��"��<��p��kBP�$�B��N�:QJYa)��ͬ2J��;�#ܽ�k(̸Rge8g����e��z�nz�'
f��9�"����$PW#w ��ju,����Ì6�t��D(�g�A������,���KS�z5��K//I�{��W�X��Z� k�K	t�F5$�gle�jn�e�#�} }#�b'�hraT���"����4F'}~��Q��v����<G���~F�!����S��7�����0�G�l�v�f. ��6��7=;s�.}�G�߮�]��w=Z*����R W߯}�ސ��ܝ���<;۵[�}���=!�4�'
o��ߜ{(�p)����!���������o)ɽ~pxw����������UߓCW;8�E�����8�?5���*���x��<�2�O�����<;�����xM�	ӵ���M�	ǀ������xC���8\>��;I����y���¸=x�����My���B�tuB6�N����8�?��{�}C�ޏ��x���UǠ��������}��o�rs�۟߭�'��?�������oHN�~[�շ'&�x�xL?nv��}�rԇ��>V.�S����=�z8S�v�f.�뷟�o��p>����ߐ�[���]�7��?����<�}q���<���C����Ǎ�P����z?v�|�'x����۷����s�������뿽�>:�̟%T\�ɮ�� A|x���90�G�
r�Ӵ��?��󷷝��O_=p}C��ۓ�G��c�np�٫�l����hoL�y�Ÿq�����Y˾���U�����ۖ0���[��C�>�я��i���yO	��!����9�'�ގ��Uߜx�}���&��Ǟ<�_����z��Rw��������P�;_��x��S~BO���7�o�s� qA�r��3��;���+Е���"!�w���xv�{Oi߿��xW�վ'��ר��~C��{C��q�0���ϓ���0���{C�o�$�����ߐ���oa�@���}EMZ��V`�0&lb7^���j3}I��xBC����~[~NMϣ���a�}v�O?v����!>,zw�;N<���<{���Wo'���]�&��������S{y�s���aw�{����ǡB"G�W��;�9ѧأ�ćx_�e>��9������1;�_x��v��o�{xw����7�~�ޓ
��k�z���a���z��w�i����O	������y��yۓ�=��&��80c�tF{*���t.�!��<�rwil�����9�:�Yĩ�����)��W���s&�tT���k��U�R��$u"�OQ�[F���Jk����WJYzk�օ1��N�d�V ��ln��j�lP@T�[S,�{��J��@�*:��[F����H�S��y�9���iv
�H�c�	��_�pyv��9w�x��aM���~�]����ߺt��r}M�9���`�����'��~���=&?��:��������I���"c~��/M%��~y�z����}�M���;��X=;)��������?�7�o_�{m?x��xq��{����P8������zw��aC㷱�s}��Dp�;�el�]��cs8�������hraO�P�zBC���F�99������N'1w��>xBO]���v���׿��)����?~�Ӿ;H��~�~t�nӽ|��؈��c��9�jO��LtW�G���fx94�/&������1;�{y���~O	��U)�9��&��?'�x:��pTbI��M��v��=��e�?[w���w��S�;^Oy7�=1�
15�B�PE�g��:�Z�^�� ���q�w�oI�?��<�����yM�	���ޏ�c�HO��X�~�'xw��<[s�<!�Ts�i7�r���P���<;���ޯ���rxG�!�W\ޟx:�	���4�G���������<!�0�����������v��	2�O���x�yw�k���뷔�Н'��<z�I�<|�	�F��2xv��ם$�t�&���:o�(�C5M���!~�)����G��<{�	�'��?�_��~����=���rraw�>~��˿;���~��|BM�	/��7�99���<�{IĞ��_��>xB��gn#�O(9@�ڹ"����oG�b!��|���V�O.�� y����y�:w�b�q9�<Y���gC2p���w�<��N������ǗxNL/������zqϔ9_q� (����G�y}�(�y���Q������!�G�)ۓ���������:���0�����P���ߟ�O�ޕ��ӽ���}O)����zO}�ؓ~B������aM�|�L�⤆ں<��,���p5���#�;��fB�䎭.!�}���O�����&����Pyw�k��{��ߓ�r}q潧����������S�ǎ?&��q�q�|����	2�O�=��Ǥ�;���>���ݼ&���+���H���MǉwW���-��r6`4�KI�wK[ᲛЯ$����b��ugf��3��..q:�|m�{cu���eτ�2j�ү��3��Ai	v����R�s���ܚ�׫�Fk ;�P+]� ��є�,��su��D��#O&)ﾐ������˃�y��=����N�?�?��.�i[�?'���É\yǸ97���=��]�1;���'���0���-��]���o�緅q����A��{/�?g�������>��h��"$�^vjp8.��I�8���N8�G�¿��'}?}�oHyL>/n�Sý�I��G��;s�zq���	��u��r�	7�yy]���1;뿹���|��.c��_��QR�W��H��X�H�#��;�����C���9]�P�ǯ����pU���{yw��n;rw�0���n����P��U>'��7���P��Nܮ��y��~O	���w�����K�>C;c�(}�>�F�����7�������w�b}�珮�ko�������˧i7����<eߝ�@�>���A���t{�������'�{;�o�Ʌ�������{C��w��� ��h�r%u�1����>�C�����I��}O=c�ĝ�[�ۓ}B}��<;_�������<�>���������N����߼yp�];O���������]�?~�xM�?1"!��c�O ���C�^9U^���������yC�raO߯�{w�xw�9ǯV9\HI������!�7q�����N����.<���oχk�a_����߾I�!&���~�������}^��[��ܹ�ۦl�/VujP{�
y��w�~���򛐾�'�וp)�;��8�{�N�~�O����;�Nq��O&vQO���~�*ǝ�����_�������^I�>�����h��w)7�t��2�}�"D|*�����o?ѽ�ɽ�����ܮ�q���P9$���������o)�!?��`�U����0s�ۓ�X><�ڭ�?�r}MΝ�$��~v�>�Ơ�@9��.֩Pv��!��k٩�8�a��ĸ`���%��O�|C�/���ɧ�hw���<te�O!��m��w�y?A�;�ro	�9��u8��
��� ����R����^���k��vw�E��s������|�\.�y����~Nq�į���I����<�~x7����￻yC����zC�����'��pǴ'w��F��O��<�>�DDP��oL�Ҷ��9�P�b���4 ʹ��5�0h����%��a�+��v�[q��Y(T��})s c�g�2i�I�������ϱ�{0�3�D��Q�&��0-�6]py��k뼚�lwh䙸�G�6
�:��]8̾�t����^�7X��(����Z��./eK��CC!��
z$�b	�~X�Q�<&�$#�ߝ�'�yv�[���y�:w���ɿ!~��߾xܮ7�y�>���7�/��=�������;�s�a��]�����{���x�@�����,���#� ���E�o�[���ÿ<���y
��aw�Ņ1!in8`�7)vc�8�B������چt. �ǝ��ܩ��">��# �W�X� }G&�;�sY���zrg�V�;^�8}�?}�S?P��[|~����N����眻��C����A��Auщ�S��{���K��7<��
q���0mC ��>#��B2;�0G��">q�_P�U<�X����vkp�.�m�L�E��roZ���s�k� y>��	�!8?����hyw�i4�O8\.��|��ߓ��|CήW��''���2�mp��;K��8�f|�y|���l��w�g��޹������>�������� �Hˆ�\0}!������������ˉğ�)���ǔ90��~��yM�	7��ӷ���I��JԇoΓ��ӷ��P�A~���ǽ�^���dybP���>�>�2c� �F?o����S|y�;�r{�>p����?���<�v��|x?'��pV;�!��c��C�qa.%�vX[����8x�wqN�`���6,��1�8��9{8{��>�@h����@������M�ރǞ��v������v��Po8�]�ڭ����x�����t�~����r��ҿO�����ǽ&�`]�ƻEɾ���"r{�Y�aEr��}!���H��z6~b4|yO!���+���ǯ}��0��C��>;rԟ'�\{v����܅�>��ӵ��z�S~Bp}=|�����>���F����@@އN�}�TmDϣrF[n�=�h��F���!��iwv�5���	pф08/-F�'��qهG|jM}�����j�s�v�>6:K�2gOW	�ń����l<�*_���r����he��N���es���X-��̥e�
�I' .W;,�>VV�#d�čl�;b�����lͱܱ�`�ܴ;��4Z��yyQEt�R�c�nb�N�%�!Y�u�{$u7&mq����u�v��5����������TәK;��k����W>ܾl���ر��S�§�G�+Q���1�9Z:��b~�'Z\KG��6q�Os9���F��B8\=�,�lНj���r|cD!�����m`���po�7��q��&��T�3ce��)�g����l���.+��#O\>���:j��V���T�j9QtD�&�(��S����F-��ý�5@�zEH�2quwM+�'�b�Z0�è;��ҥ<�7R�A�U�+z����i�7��8��<�%�t8<��b�&���*��!�#�`���=��#clbz�ӓ��n�@��q�MF_����7\σ� �q����S���;�ы�R5��3W!��WS&��Cm0�("�<�ŵR+�Y<ɣm��=�b�3���������MT�ȷ��!�6��������ey�CƤ��b�y�����/9{{F5��זCc���$�d(3�!�D����c�i�d��D���鍚��O���j�Uw�0rȽ��.
mG�.�9��[�Ϩ�e��]l��Z�����f�D6��U�o�����uӾ��9-��z�U�ib�Y����"e��1�Z_Ru� j����^tn��u7��1�t�샩�|��2���C��yS'k�Α�mPTc����OS�{{Rv�Hx�ϽW�ad�C�pJ^u��c���n�B�Vd�o#�3
�L��]�	VE�~�2�M܃h�{S!J�A��'r���k�j�v�'��H��;�d�F;���շ��Hɋu7 ��<�"atV��߻ĜZƍ�B9��Ɲ�}���r7*�@2��y����nxF�ם@��Z8OӨBt�������C��et���ʩ��˴�`�`2��Br�Y���+N<.j�Cy�nu�T�n���_�rATe� �TN�o;(�t�(�N�����̇0�[��0�J$E�@��]������F"F�Y'�@@�s i����t�p�r�~�n����˙l��Yݦ3&�����s��h�ըl��Jâ+�����&��f@�P´`u着ο���{4�Ї|�U=��ƀ�^o�u1u� p�C��{������C���t3�]Q�rDg�ƾ�N�9�s�8^Vq�U�R�g�f�-w*����z��Ġ�?�J��+�Eh*d�.�;�����t&���2���]ܨ��"���q�o�#����a�:ٱ@��쮁�zt6�� 0��'c��L�/S��dM�Y��ܧ���s1��U��,j}��,�T���S7<�kL�zt.��{��.\�:7b����c9�:=�pb˜d��X���̎ٗ3�a�ڲ��K�@�����X2va	Xaj���5:���2cc�vh�'1�3��΋�SX���H@8��2M"�q���]���]q�ꗆ�A���ڮ�B�'wA�S
h=wfmk\�Rx��1)썄8X��������ܠ��Iz�2���G��Ɓ�+�5��5�*��O/zxvL膵���t�^���y ��n�B���h�����R�[�͋��jF�HA�f�o���!�n~|SWT�Ӹ��D<<5(�f�m����184߻���ߌ�k�OX�R���w��o&�"�܎��e3��X;�(B�-�[�^����=�\2���'iYё��6] ��3EDr����}����I3{׋J�{��5�2i�pЄ!�A�.�҄����H,�.�,�.���������:�U=�=�٤?#���X���rE]������e�պ���A����L��ѼpD�{��q$Zs��7�1U�N���X�/�E5��t��]������1'C��غn���|D�G,�մ�p�i�ݼ�W�\.�95�r��KNnKn�u�Eq��y�M�ϖ���)��yպ�n87+L��:���r����D�C6�5O�}ϋy\\[j5mp��^���}���G ��|��8Pä�s�T�_V�E����_,�W׌�Ǝ�j��J.�i�5.��s��m��������ݠ�c����@W��ڰyy��G^(��]��^��a���m1ձ��%����1�q�"5�"��3Ă*f]�\nM]>rz:��X�_,�΃=�i�myÀV����=�S6wN1��j`��w�+Wf�-y
f�+;�w{��B�$�A��5�����_:cp)a�A|~ʈ���[VY�ΫO���6o��Y����r�tG��J��-����Eƻ�'�|<����Ʌ�����LnV;�8�k�֍���:t�@�5:� ���(��BӐ^Tdǭ��}�sb�m^8��������TD8���A55Ed+��\����&#����M���T��q�p[)q��3%R.+�2�Ԧ4TneG_ܝ��΀t� m���wT+Jɜ�0�1c��O��U^��)�oz1!���T̈́3�_�����j�0�pW�Ks۫�*�&����>��x{���N�I�I�H����7e�2�m4S�][A�5�1N���gmqV5u��8$
 7�A���9��u��ջy��<�jOU�ݵ��w�6;���=���0JA�����q���q���X]j�*Y�Z���3�	.�~��>ۻ
C��6:�a�+NR�h�B(<��g���Ԁ��k>t���8�치ˆz(�*����v��jb���*ﱕ\½/�����xk�U\�(`����6W��:~M{g�3�司�UC�rW��q���B���7�@wL�^H��7t0j��K���c�V�	��{�o��T�����ʦ�C.�q'KFx�+��JÎy���A�Wn�{!|���B�fF��ˬ՟�Yc�l�ĵLnNV��l���'\�H8d�f��~�5N ��������,�lК�j���!��"�Cw��K4�C������P��i���M(_�N��#86R?\b��e��1�}e�x��Z�L\(�q�L�mî7�A҇:��F�.�y��
tEDbu�FD���ٖ瓶e�X @xY��z����z��N`�߄�ф>��tZ:2`c�֔/F�C�S�*��ʎ�>�ֆD����jpJ�����4vH����}���c�j�<�6�,�w��Cp�k�`�@�gT&ކ���,��7T�w䭹J�j>��/V��AD1��<x�k�ph�η��*#��{���b��1�)��/�Lk����z����/�Z��wo�ڼU�HV�7�F��8cL:*�E[��٫�}_}���΅��Uy��kF��ry7\��4!CJ�5҉�b	��x��Me���hZk�y�+�w;��	��ڥq�O��mT��Y<ɣm��|��W�M��\n�L]��.���rYs��{~�GZ�y�Y�W���'����G{��[����ffZ�c�Of�����tP��v�
��(zk��b�ݔ���������O�A�,��'�Y�t����i��a�'�_y!�jʚ� H�#ԷN�VO>c6cC�:5���Y������?e?;A�\Nc����l�躈xFN��=��|y��D����1Z�x����N��z)��`xZ5,�>��딴^?*oC�[+=�Ұ�/UjDɸW1	��@+%�M}�S/����[����օOF?7!~y��ީ�끒M�����-J%�;B����̓+
e����JUW}���U�-�ڄ��l��$�,	�!
�'z�9�%�1@�t�ݮ!�STW�SY���TQ+�Yg\�J���o>)����Tw;(v���t�f����/���@�.s�!��@��}CbRh�c�d����7(�'�=46�!�m�K��ׁl�Ie̮rZɮL���ݛZ�ދ�T��Jre��qF3�g�]f.�i��C �⮭�.�֘�o�=���h@E��'n�j�.�57Jo�7i�)1g/:k�ό�5��@�����ct���r�:�hm��UZ�kT�<˝v� ͬ�)B�#q��-ޤ���wqˡ�"Ϫ�fq�m�+nS�QL�Q�o��]Z�1t��k��ë�Z*d���l�s�w��f�Q�����;�1��n����+�b�lɉ���F��0y�x��CX��rUv�и�<���t�TB��:S�ɛ�\�Z�Q�`.ڲ/D�B@P3��3�ꫵܤK��]�SL桮�ߙ�x��m��87j�-�S:��/�;]��CiQל�bW��ek�TRV����t�j�wW+aݱ���1n|2���:	�CD�mاnXB̓��y�b��\uQ�F�m�Ū�Elio^k�j�)N�m���"f�ؗX�ڛ���ٴlE��Z�6�p91г�����-D�j�Dɑ��q�;k%�5���f52�h�����u��	v�4BЖ!\v�0G�6�,�9&��W�N���P���R�"B٣�E�r�*�]gz�Q:�4�fŎ�U���)�r�s��ھ�j5
������q�:�	��`��N�tDT�������XS��=ޜ��5�'Ӆ޽x	�j���oc��]�5@�( r��Kll=�X��gɐP�W��5�G�<�[:�P���#q����[�7Ә09�����I^��Is��ʮ<48næ�ש%�j!ա�m+9s�![)�$u��\u�2�J ���C��~9^G"Y{	�x�N�R�k�>Ψ�\n�C����沨i''j�[�Sۭ�ݢ��>|-�{�uv�������"t�ɟF3~�u�ܒ�iR���/��ǩ]\����xx��\@�Gv��Z�^���Q��9��W�<��n#ۮ����3��W�3�6���K�ՖC5��c�4�Z����v"5�l�;}�u�Fք�gm��Իr�9]���`,� c�Y,V����B6b��>�p��Y��̹vV�m��f�C7W�r"�Di2y��M!���V�]��E�SrR�A3�O�ֲ��U���p��M.&=y.e�9�&��sw����l*}; ����2��r_n��Q���*֜!�n�#N�[�QΙy��RZԁ|��#�W�p]�42�̷H���_��L�!l�˝̰T����wX�-����૙yØ�vټnT���H��n邶Κ֙:���&f�t���8�dv��@R�A�$��-K!8��n����Ny����PN�T���(�J�9z"v�wwHr$�d���G#��s�\�M*.P�.cu"l��O:���"M���S$�X@�y9�bj2�uJ�ے�*��!!ɔ�r�z�D�N9�w
�*�qݣ�sΑ�u՚�wv��8��an�h��A�J�!S�����	���t��2��MrO5�=��;(\$�����]۹`�]�Dt�wI"Ɉy��㣞��9jD�ABE���^EFN�x��橔�.�;�$�s8�vQ�W'<�wGsU����+��R�4��%��P�$��
/	�s�%�Ԋ��F�s1c�y��ԓe����H�H�Z$H��8Y��QJ�E����x�u"Ӕ���\�WN5r���z��%)�)@��Z�y��w�؇P�uT��7�N�(�Wx���	����j��[?�����q�Fl�v�^@�߻��3��P(G	��=FP;��a"��t�;���ㅣ�߽g�d�b�mLS��#۞B�P�\�j��L��R�&���V2b�wfҕfʕ�����.���G.��݄�p�m.	֤us�8R�x}�^�X�H-�{q�r���\r�����_Zg���D3b!��-��*؃1�$�.�a
&�Kzz+S}�MYpL�X���h��
S7��&3�S�М�b��d�u����E��-�]'��c6��>Đ�T44��g1��/��p��4�i��CNxT����f�D�>��YY�yi�!�wC�j��`{���p�1����"��3J�� x+��P���cf<� �Ĳ&}�{�v]�}XpK_z�!����eC�:O	#o.��Rqq����6-��>�c�W�<�Qv0V&�>uLE�t��u��bD���D`D�X6��ڛ"Pd�z��":Qo�B��Q9X_Ʀ��en�[z�m����LN~����.�X8c6|�$\#��[�}Z����-���ѧP��귆p�vM�CB-���:���l*=����Ŕ߯��s��52a�k��t��* &j���>��A�t�]Nݮ��w����7c.l�z���n�G�Z�2X����M-�b�����Z{cp�W���OUc�]�2�E�j�xa��'��������T�d�Q�Go����ӚRh�b�{�@����m�Ȥb�q6m�Ό���ξ��gFT���@;�L�ȦX)�6xݗ���u�#n:)-�_V���Uq	�˚(8���k�bμ�a���TY�Յ�]|r�R�,ub$v���oi�/��{���w\����E��>?w����t�������������k��5I\���r��W�\�:�h��rn��1o���$�0��.�y0
�m�{���i^]w��z~��<<�f1=���{�#nWʁ�z�� �w[a�嚜򱳏������Ƣ�1U������c��sv���چ�fQ��ȻFon�[%(v�n�D8�#W��D�*�W�6S(F|�+qc�F��@���i�@��'�L$Vox�K�E	꛼2�f0�7>��s顴���e��*9u��'����5<|���*fa��j�2��ys@1���$gS�Q	�E�A�wH����f���Me'��{�j�����v	0��1���VP�u���o7������z��I{#��[�V���k�Y�4C]�SS;v��� �E���Հܷ3��y�T	�u�y%gWL�����%�1wMm��sD��խ56d�.���ѳ�\�_v#��>��F�R/��nH��gT���KL��ŀ19�"c�'j�����E}���s�"	��D���ľ�}��ؐ�z��=om�mUѿ�2��4�sC`;?	��OT���}�l�
z&SA��ΈW*�kC�Ք؍� ���uع���>��$a����biV�'X�};`��q�=����L�c:�q:wJe�vڿ�
�zPϡ:����К�E���+����L7Ս�/��Q�J���Ds� ��"�-/x����@V�X���1��.*�ڹ�q�hOU9��+~�ڬ�Wd��a	��_u�^��J�b�05춫d5��o���Q��L�
ڿ�ĺl����0��Lia�x�s+� �\�x�9�@���P�������!	���'������~<����heծ$�#���<.�T��o]dً7����Ѝ��	�b��[�#h<��5��ܿ��6b�cMΎ�l����sJ���wd�J�V�5�-��^ڨ�Q�BkZ�Ǚ�Cp��f�p]]~S�.��ú�c&��N!ժ��@� �k]e� E3,���́e�9��F�7�wA�sY�˓�N��6��S�����+o9f%O:�����Ӡq1;F��#��w��B�V�{3ei"+A� �z�p�oDe�\󊓜�wߩ�m������v���<��)a���8k�  (t�3ce#��ت��n~!����s��.z���J�A��癁��:>�UʸTt0��������@�=�mX*w��/�D�j4k|��k�{�'r۞������E�-|:����ўQ��Z�=��6��/�w8���'���4sj�_���jp
V�@�0�8$l�©���<{e�ϮMɪ.+%�ל��+�h�e�UMD&�x0�F��T��}҉�Zˠl}�)/.;�ͮ�k��\69�z�q�O���Ď�Y<ɣq��W�6Ww{��Gޟf.�7�=�����"_��ߩh|qF}g�ey�+˅�$�ь��O�Oc�&q$��	����e�����J�Zv�Q���I�*�������i�.u��
°o�x<Kr����{yOn(���7e��τߥ�c|�fa�s��Hk���ad��r(�9����-Z�����e�FS�f����9�?L[��w0��*p��t�ײ?e��M�hu�c���	L�y��ugܥ1!���xߚ�Z����d�����u��w:R�<e�9Z#z��M��$�T�u9t��H��\y:]t�Lcb̝A�nI��������:�����7��H��y}���>M*a��u����">��
������bǌ��+$� ��܅F%����sU�.:�E^�I��y�AY'
��kG'���� ��b�m�Wro�b:\���Y5�2�a���/�(+v��5�)�O�AjP^rG�OxK��S�I�0s�%��^]�.��X�|�9`�`2����eoc��T��T��b�4w��1\f����t!���k�J=�(�S�>�p�Yj�H�oS��@�T�N6`#��j��6�D�ᡒu@H=�d\�H�+�-�1��J�YmM��\t�en	zt`�rх�F���8T��J<>��e '�i9b�nHy�q�
C��J�n�:�B�������8YwO����&��R]2zU� !,��.I�Kf��бs�����b�PN�`��1q�����As�9�yXS`j�se��5r����Wj�����|Z� P����H��
S:8��{N�#!ͲY�ɮ�78�]�]C�7����3���ԐW�(�S�T#��:�B��(-1z�i�N�;�<*LF���������uMN��0�=\A��kTa�6��NPzn*�b��T�󷲸C���Cx��1������O]OUW��@���۷:̃f���3
(�^3�qk��,��6�m<���G3t�\n���P�`8�jv�%3�\��^�  f��mE��1uXQ�\yu� ��Q7�<Lt1}�<�b��[��o*���*+Rt�xD�Y���}c�7�ؾ>��U�l �*��h����B*��~��r5�W� �;�v.�q�g$�;CE���b�U1���Y@r���!�C�j:M �_8��w�,��e��T}%k�Y��:��!/:S;���=S-��]D����T�P�oâ�P��SP�� ��7%���J���4�4�s�yޛj�,�h��ڿ�M��4���b��_,g��r>q�E:��F�Dk�%�@��gF|iPjse��L�Q�S,��>��"��1��
��U%I�+�����(˚(8��Ƽ�ŝyda��kSn	�{Mž��o�Q�y�w����Y����r��u������2�Ś���QQ�z�^Xh܏���Z$��u�Ocd�{��⯗�*_���r���fDL[��
l:I��`W�(l�^b�}��U�g��;�q@z������Y�/O�Z��>�!��{D-/zdd���&|�Ic/:�UBcy�����ʦ�ˀk�'3M$m��)�Sz;2_hy7{O-;A^ X�k�j�fw�@�VjNa����H�����ؠ]3����(m�lngIh:�.촵�=θ�ڔ]qnu]������`P\� �m5p��gV�;����G�C=�TKK fϧ$	���CCE_ت���D��;��sv�����<'z26s��,��L��D�!Q.��J���L��_b����Jvٌ&��\�|�Ykufź��^�s��b����K�	����DϦ�GZ�cr��|~�g C�4&]ƩÝ�k:5�i!��欲R%s���˚���	T��0�#���=ƕD�er�i�J��x��P��4�]r��?kJ�-��֪0 ��#�'tHw0̒�T�n'l��H��&jr���Cf�n��Om�mUѸ����e���,�����y��:�*jK�Rތ��966[���ґl�S*7'u�'oL��X�Pc?e��v7�{.x�r��D;}9(*
�,��}B/��c�={uSy<4a����%��=��"�Sy|^�_QPy�k'���AF�
�1b}'���1�&�:���0�9��g%�.����pZ���R�i���lʏa�Y�kM�ƀ�eW+��r�J6m߯�dՀ�ֻ�R7��&EhN-��cq���6��c&;�'ޣ���-�)�=�yM��)����Lw�7b��Rn@p�����nE۵.�N�W8jd�s���ۏ��g�1�Á����t�Sg�q�W;��G�sH��}��ﾪ���m�28;=�[H�u�J�}��k���s����Ɣ;e������u[+!�W�LI�ڡ�ԗ�_P�*��}��EZ����򘎷U��5?dv�Hˈ�D�'/��a���i��^ͺhg1g3u�}.cI��Af�+�\�*#O�,���6b�Z�7>���̌����c�ᑋ&�	ܴ��"a���%��Ԁ���b�[0Y��Zվ9�2�ƈC��j���Ͳq�g�����e���<z a(	�t�3p6R?\b��e����#P��(��^.s��*L�N�0�����p��F�QG��!R5�Hg�d�|zN��R�v��z����9*� o17?Mƽ�o,�e��4S<qh�� w:���Jy�sU̢�=~az�8�z�Ď���;]A7�V�nQ0�XD��NJ����s��D��(��4h���*��Tq�ns6[�_iB���ri7\�,���&R�&[��6�2����'�2����Y��7���j�Ǔ���U)d�&��۠9�O@sؼ^�"B��t��59K��n�c�m�N[�7qG*��(�?"e5���G�0d���%�s�]&�KݸNK�%Ne-�@,ݖn�`�ՇvbRm!��x�r��×l{f�Ӷ�+�i��/ ��3x�,���X{��]32�IK"��*8�?�U}U��݃ֽ+h~��Y&~S���J_.��:��(��xW�z�CƧI�`�{��ܑz�t"��q{b3٭��\�e3+�A��tA��B��פ�K%��|��,NQ��C`���$�nݿ��v1��R��|v��P���N��c��� u�P�V_Rb�_��z5��H)� �St#,�2��0����|�>��d��DeN挞���{�͗:�M$��~syPř�D��m>y#>W0�,�k'c���tm�䘽D�V��5��_�d�"pg�K��+κ��wro�b7��d�ɨ�)����5�uܻb~�Y>��⫰��M�/d�=SSF�$Ԣxz�X9��ߒ��$+q:�^�L�eY����1.��zo�<Wp~�G��j�j��c�`����P>��^��>{,�\i��9��~��/��Qk�|�GR�s�������3�@�'�$�|e0s��$q�p�*�bԳ��)J*j
uݜ$\K�0XΥ�E_Cѹ��CV��`�Nò
� �5Y��;�=W'#�c������53�.sӑ���u\��O�z��%�<G���Y�{���:�r�ķ���E2j��m"i��[ڋ�5���-3C���~�*��՜���.ӻ�U��j�_�s`��ܲ���S�^��ҕK�6f���b.8����W�W���.y���ޔ�>�Ô6V�H�h��[�;�Z4���W���D�Ks����r�E�������|����� E��\k�NR*���/+����u�.������Ko���I|d�I���c����ocN��8H������8C9ewWK��tG`\ν97� U��$U�z�x>tċ�(-1z�i��C���`.�O3K�ؚLkf��0��]f��s��`] � {��|��x���Ҿ�7�Z�p�L�V�e�S�眠5��w����u��r]���ic�֐..'�"��a�'v_�Y���\�߷0-c�㺑����VK�X��B5��X:X�5�ȍ�YP�pD�M�b���tw]B3��cX��L�����z�n��7��N��ў35AjBC�!�y��PEvF���Qا��f�1Q�N�$�i��UI�L��s�C�:�L��"�\Ch֞rܶ���L�7�dW^����2���v]iPjt�A�굉/[V�23y�:Ăy�,�����ـFL��S2�RB-C��_Q7���h�{�u�due_�v�� vS=WNr�D7�ٺ9�,)�"5*+I��A�|�r:^tlӜ����m�������V�v��g�C�J�%:CV��7��m 3J���e��S�QcS���-n�j"t����}�М��n�&jH�ݷr0},���!�3��\ì��7Y@����Ҳ���6����k�t��l�X��ק�\u�;�C��^�kR�k4m서��+a�� ��!1.�ώ�8YJ�n<wn��2㕷Ir�T-�OvX��4���i(��t�.�¶�6s�-TG���YZ΍�\k�f��G����m[{	��c;L ��D���^���)N�S��.	QM�V�j��G��M1��pX�sc�\���ӛ» ��{�<�K8V�K_8�I�e;n����q��5��ſ
YR�0�X�鲝1��F-k:c�*R�o`�-���b����m�L˝L�f,fe��cH`�Um[/o�awK�@T����)�5��3�ol;�63�<=��wWyC�K�6"HWJ fm�:zGְ<�	�eپD��e���cR������@m�z���h����V�0�lQ�l��*��M������z��v@B}���\�k��%��<���V�]�̏^8�<��.̠D4�0�bj��M�s�Ch@�Y0�fή"�?�.|�[ɲ�_\t`��t��>(
%
꽠�XC8^�k�biMǝ�Wx�������Nƶ�_Ñ���M��{��8Fe��q�ӓ��u�2���0��+-W(�j�Ѧ�̙r�Pu�V2�rUp�΂����Ul
k�75 �[�.�L�U*8��"�M\q*��d��٨�8­�1	��#­8طمi�Z��}y"	b�	�=�_^q���@����iк}�;z�I��j�=[}n軄F��Xi:u��bA���ٱv�P��hF�ʃ��,P�R��u�c��7kL����t��
�v�39	u�k�T��X���p�Y�*fp�*Vm�nCZ�y!yW#�ۊýf�U�kr���WvY�a�{)LSSx��)-���\�{:�ޞ=��GMy|[�{X\�J��[�i����hf�w�mbF�ǲ뇻nV���,�x�,���e�뱋+�j�8�i��ܴ��k_Ig���L�`��_P�K7>w�VJF\YN	ӝ�L�Xl-����2�hbq�8pik�Q�j�Nn�疺朓h
�F���91�n�;@��=�{ݙ���V�@G�F�cU���z�,jԛET��N���r�Z�z@��p���8F�o���Խ�s��m��O���tgcW�uq�C���i<���H!��sn�ol��5j�"[��C��n�]�,F#[��ͥ��?e���4u\ċا[��WN5��u.5(�L��h�|qU���.�	�=�=�Ww9xa��WH�L��I2�Cu�)9̄R��uemB�P����^a�\s"�N�����.���諮�eR�ED��jJ�i��r:T%r����!FTbf�Ъ(���P��!$�l"'S�HK	'\;��s�,�ԫ̎�.Bd�"e�2ʦ��S=���U���BjB�J�^���<�JP�LR3�JNG)DR��9�""^�臫��A�adZY��:���y��D��ȣ*��s�C��[Cܮ��U�,��DTa\WOvr'	g4C-
�.GQMLZ��ȳ,1:�����ڑF��:*�=���]3#�"��4w#ڪ*�\EH�.�����ܜ���q�N膒�W�f*���eM"n�u#�������i�
'D�jê�f�CIZZ���99�JԜ�p��C�"@�~�"�l����+.����0ɰu@��u����ˋc�۰)�Ļ�Eպ��VRS38Ϋ��V�p���T��_�>�>�p��ʭ�ls�#�R; |5�H�7���lp�]y�B�҅�Em*�o��Q�N�ܵz
̽�|�t��z��C�"�l���=�TU�N�c\n������&���r�g�	S��m8��A���؅�[����C.!��ۿ��GGh8�b $��m���c�M����yc��C�M����u�K2��T����1Hז���{��g�h[�g�vR�)^м��Jq� ͚���`��"�����U�㔚����;��0�i��ݜ�;����幻�D'���H"-��ȋ�������YC�B�b�Oqd���|t��ԣj��q��7%�Պ�w�u��A�3���1��H�t��Sg@R��	B[�8v�ci��ΧO��j�amYg"	�D�u�*��%S�T�N��F�ey�G�����΅�R�1.#:�-j�0�ꟚR�i�`sϫ�9�"x�v�B�ƕ�61hY=pO9Z�KbEK��$i���mUѸ����Br���eX��z�����=���*J=r�'�ن�[�9]�X������ma��O  �q���gp�cUl�d�+Ul;�cy��9�4���eq*��7�֢���]G���o�����iU�Q9*S�Xd,�i�^:��R�A1�zQ�>|#}���i��ŷ�22LS��W���Tz;���44v����Z-���4TnN������@:S�Z#��P�R=U'�޹JNJ����γB��'�Q3a���\O�q�j��Uƨ�lmc*3Y���7�R�X��C`�`����Wh�~����M嚣���#��=.��b؋~vJIFl�h�� �|q�V7�s�v<�����*�*�xG��@��x3h;�Yg{�1�@B�p>��:�)t���]}�m\�ܩ�A�A��g63�oZ�S��v%Rj&�h�3%µ@%�qwc��;�R��ה�u�:�nDM���ܾt=R#�&̴���|@=����L��a;'�U�26�]f���Y���
%�cx��1Y*�v.�|��B�dĢ�'j&XT+��!��=�Bj5�|r9�e�<�$S[��L�c�]m�����02��F�� �������jUƂ�Ld�"��2�=�H�2J0;v�-ly�.�Kv���u�w̰y.6�yvy�ѐ�mH�M�M#�,ۗїf9���q��$ɛ�t>F�E&�)*��F%c�>5%�U�0�n_�V,r��@��s�"�N%sp�9̓���4�](fd;��C"�u$V���e�*O�X��d��%�B�f�t�+:�|�U}�}T��&��<�\wE�W��m\C��3���m����K?OUU�'�Ӱ�.���ݡno�Ӕ����a��b���pF��ա������ T�'!ӓ&rA��˻��r+[]�}6E��'�tn�Z=y��b��Q�	T94���L���.t.��"GD�s�W�e��1 6M�a�"�o-�v�Jd`Ӟg�U�M��Y<ɣg�zE���Vȷ��4�n�&��� �yP<���n-Ƈâ�Y�����x��Gc�@���e�B~y���Mf��S޹f��*����v�
��(zV��&�`�_�㾬~���J�U�A��E�9���xG(}�lX���&L+�*C]YLvN��ݎ�a��6�ɉ��b� ���4������;a=٦���'�H�(��5\�@�/�}
�EF�f�����/�2�+$� �O�H�W0�7���?MwOB�T�����@ldn[���5��N��n�˯;�m��U�t�q,�y��/�;>��u�+u�l�+:DZ�5�9�u���#�{Y*�[�g�$����ɣg�/�^�Vx��^�\�%���_ESF�쎜YZ�)�*�U}o�"T�K���;����+�,^Q�T�(�q�{��.���Mcؕ:�k�������ṛ6kw2< �*�pPY��ح���h���$�'G�%���ߒ��HVT�_+�.�"Y��Zʛ��5�-�q<E��e:u�q���D9���e4�pk\��1�4�<�_$^\��\��G:(�o_�T:C1�u�P���΃��Ę`�����Y�o8ڦ�y��E+*��j���v@��Lv��58���l��Y��P��#�����G
u�Վ��Eh�w@T�<���W؟\M�w,���v!:��������?`+T��^����- p��S��l�/H|zu}��D3b/��ްfdg�ڝS1�%��퍺�L���Ƨȁ \
^�q=)��dY�Egb�b�9���v�uuZ��1�X)�}Z��fs�8�I�44��O]	p]K� ����g.�Y+��=)��Q���lȧ�¤�G$�Ѵ�#]�
���Y���CW��Y�X�]h
0E1����̥�����kix���<݇\|%u�^^�>S��n.'�vӼ:/��}*3s�>4^!�<-��u�hhM�����+;7M�t�'���Bթ�L����wT�S�^ԉ��#���G V�%nl��t��c�V�k��Z��p�SM,�.T�%L�(N�٫J&�E�77��'q��ӹ���f4ؙÃFuv��?z&r�
��>_w[/ᕒ��*�"���c��t�^���v�;V�F[w��ox'\��7fD�[G(ƈ�Q�)���a}&C�3��|Ѷ��wr�����[!��mn�Ψ{�Ńf ���G����yw�>-O���J����&Y&z
���f�M-�G�ghb	fB���?2�߮�״���,�5�]�iPjs�a�Q�Q�y�����U��Kj3c8ܕł�[:��ݿ�gxl.�W
���i�t������]t��hbc�l#�J�#K���P�����d;�d�1P�*Q�� F�������M��W���ډJ����ONY��J�B�-ތ�q0�[�#�׼�������ұ7χ��~8�����D�f~�q@Um6V.��f���D���r���B�p��F�bz�Z��hRP��} F�w��c@;�˻NjJb,hH��Ucx�j�TL��n ��;MI� v���1Y�zi<�Y�s���/�Ⲣ@�]DC�!.��=�§ÆB�[8����n[��'j5��r.��h��X��e+�\/;�]9��}ռ�Uz���9�`�-��j�@ӵ�Hp��Dsnj̱:��j���Y#汒KGL��ء�՘�����)K�v��qVw�����'c��V�S�����4_du���]D;�7�ǠS�;`L5-0�I΋*kIODėμ5N"�}0y�z��N
��Ts�a ڢ�\O8u�*�
����z��K�'&7�{�2-�>��Mȩ.2�q��w�\�!���t�S��`s��N`��(��[��)��{���������g�aW��KXR4�Tj{ld6���@�@A2���eX�U�e���<c#��Զ���.p�@��6�a�i�V��z&R���4��ϗ:Ҝq8֨��b�F�/^�?w�;�q�f�+�3�e��I�	��I�*E�3_:��i���h���������l;�'��"�К�~[�mAF������"��+��������񫗃b���g	z��7�\ �Өb6�l?;2=����kM�3�B� XC̪������u�1�
  �PS�=�Bs�?�^�x����0�k̖����k뱻�j�Es����'�mAhԝ� 5�]�����"�Ԧ����pcr&�♐�*lÊNv�T��Z��h���C�gi�����q��{{�����J�9�(��ǖ�oR�g�d�j���s6�ƭq�{�Y�p��B� S��\ �U�<�U��gu�R�{k���z!�1�eq�"�%�qEYԹD˘m�l�t��ۂ	�f`)��6�����z�LY'
h9��ɢ�q;,<9ҫvdma��hYn}ˌw���L���B��V%���ѭ	�NWp�$�({0�u!\b��lК֭���B���/]H�NV�!g0����]vK� >=��0�DTO ���Lb�?9�sƈ|���~���E_�RfC�C�ߩ�� O�h3C��^U£�х�QGT|�"�I�]K�ۛ�c�f"���]:��DV7\4d��!��Нwp�A����* 
b$n"{F|X���{�/@��=@���F+�pF��MZ[�LXb�&�jp
�V�'�,R���9�ip�o�[(�AxnΣ,�;NMf�s��(T�����p/� ѥ;(�,�6nmN�3x�M *��4����L�?\\��{�6߂�T��s���L���,�w��U��W��ⷷIg�S|���lAL��T6�d�����T��>5�3�(W�
&���ݢ{z뙪_��w��|jW�}�wؐS>��7Xz�@yPj�XUYC��Fz����g��IN�p����$�б�r�|v��K��E0"0�j�����\��Q����_�K�0��ٺ�t�Y-:�����J�1IDq�扛�����n����3�����%!;�g%ٵ�t�x6�ܶ>omk��/cؚ�Y֢�T�9�����1����H�tc��c���<�Wez?��a��k�gI��΁'�\�`���:wt�1��G#d�����l_n:�.�u�뙆��ñ����\wv0���s���N<A5.EI�s�!H[�1��D�����$g��&��ضo��c"J�p�&=�J�ng�=�#Hi<Q�S�2YgL��ɀ;L�rw�'��S/q���9q���
yʶ������뮴/�&��"M*'G��/.��:��
u���.�����z�f����*%�A�4�)��:U��/��<k�ȃ��U�\-r׊s����q���_EM�]t�Zձ�Ƹt�d9���6�l��
Ã$�@��Q����gO-4y��U2Ʌ���Aw�p�Yb���h�>��m���*�b�8�#�����wmn\�wx3�I�a��>
���D��4R��N�q7�P�+/w�cͱ܏<��7����d���!�����n�"���s��.pCfn�\37NNQ���V���S�Je?��%r�BRj[��`8*rs=�O4x��Jϥ��l��k��f��5�ǯ@���ˍ9Zɩ�HV�����1m�GT�.�j�"*��v�{�U�xPp�WM	s���|ժ�h�X�+e���"Y�諭�����1y��׊u��G�?+W�"nHWb��{Ѭy V�̞r��|�������Ԥ'�i����d�82�d$`i�8鱙J��PZa7�����h���:�a;�Z:�d&�I�杚)��}
�	Y�0��߯��^�WA���'BY�.50f�V'��t��2{sgz��l�Q��dN ����~�kuI����e���^e�.k;���c�R��k�<��l;��l-LL��oBCd,�u��%}�\��a�5�_o9�]���3�oZ�]vc�ֱ�rZc�iҟ���Zf����Q����хD�>q�.w�����ƺ���^<}~�検����������o����Pvz�S}g$�t��œ)��ק�W4�r�t*��E���e���!ʫ
_&�Y��T���T4�y]�4�W[j�����q�\Rxg��{]q��N��`�-�l��J��)��xF���@����U��}��[H���¸3V�������1OQ�l�<��7������6��C�[�R����W���
��ȸ[�W%�u����"�6��qf�[˴�eE��C�y?������k�͓���~��Y���lv��8k���{poz���mM��[�7
��K������\�J�mRސ׊���F��'�c�̜�:�� �|�/�D�
[�C�����G��5%x�8���C�n*	Cw+2;�47���1�]�L\Ôx��pb������ ,��w�����P�SrZ�ѯ��i������R�v6�7�s�)T�����c���0��^�+�����|3���\Ն�;�V�B�c�������n�2v@�I{=G�{\XT��h�����i0�q��N�[<s@�|z{}���{��٫��g>��%�-sf�7V�jz�S=)��klGs_f�GK)��CY������?|�S�����o�
?(ߖ��f���nV��㞐�:�}��r��g�w�N��>u��=�٤��UE3R����v\�M'r����T��Ԃv�^>�oJ�ā�&�9P�)r�ͣ"zmǢ�:'9qA�Dͣ����r���T�z��T�L�W���+�X�qܒw��Wl_����!��5�jm�E�)�BY=�d��V����Uu���1ŸB�[�ΜX��2�a�5�UѺ*����7e�HV+�ܫ;�s�&���
��z,���CyV�	��[H�_ӴaN�$/9
EM�	�AРN�ҧ��t�
��l�+����
��2�@����y��n�3V��f�<m�j-�ً�X�gkp;v�Tm����z27�9�1�b6��v)q�j���#[F��^�A�S�*e�^���Q\�Xڕ�K;w�
\��^-]�n�
L�<{��2
��@��Ԛa.-8�Q��d6�NdWHv �x�c��C�^e��\Pg(��f)��v��_m�l���e.������e<,�.κ�(4�<K9J��ldK�C���wP喤7�Pa�[�Te�.X�d !x��\�9�:�����k�)X�>^�zl��z�-Nj�uR�YG;m��ȭ�l�;���,�w0a��s(��Y�\�ׯ�
��Bt�z�`�5�J_1���[��'�\��(|�^�;T�w$���d�N�wL�ž�yqYu�R�-Fu=�u:o�![K�����C��Ʃ���ΡF����ëc	��ԙҞ���;5{9�,�.[z�a�6Ad�۵�.�*����=dٴ�ˮ��hҜ��Arް�׍A+k�E���M���8|��8NN�!��� �]�Q�A���i�A�����JX�i΁��Y�����x2&��	�n�-�$c�>�A����UFh�YNۘ�֍�W�Qs��w���+��C�yԀ71B�m�h�.�氰��֡�[3c���'pI�t���&�a��Y[L<��e�+)y�(��(�чc�u�5����%�E��f���v<����uw�a��(����z����N�Ci�� �ofK*�%���ҥ�Do���:��`EV3Z⫫%�m>���r�=���1�ZǀɆ��ݢ�N	�[���u�O@,�hü�����]u<U�l	��N�f�Mؙ��b���e����R�F�u.��-�}1d�P
�f�L��f�yAR��0wv�5���ˠ��g2��O-�J�|d+j�/h���2���:,y���X�v�&��oP���޵a�����jn[\_��p.�\���f����clӀ�:���׍H�Ӊ���+ޏ��f���Id�Yyr��ᮮy����-D��]�u��WG�;3M��5b&��Ю��@k\���)��a��s\���Kw:�v�$����P��@/��Q�-����/"�gq��1'�X��W>̋M�^e�&ǔ"��D�9��݂Yb�'V��gs���nHT��e�u����XJ�لAQUPP�y�Y��]�4�CY�t&P��A*��{���Ha���y%�;�,��)��;�$Zar�MU��*�I2�5i�%g��^!��ջ��TI����'t��t,�ʓ-*۩���p�j�K��%s1�wAh.C�ZZ�:8�D�ԥ��Az��y���u(�ʰ���VDE!F\�ݘ���I�,�[���a�%�QR�0�P#�H�͛$�+$�V-M&����"����Y����DDA��3�WJ$1i�KR5L��-k%��P�*L��9f(\�it"4ws��Y�fIQ�F�(�-EYf%�)�K/LHBВ�C�'NU�E�t+#@�3,%��qB�ˢe�A�ZF��NK4ᴤ�a�i�2�"�U
�QQeU�S��f����U�%7D�/J�w7sQs��w	B�k3V�m�L�b{����u��V�T��w���.�5�Xz�J%b�L��ғG0뢮�9�y0n��#�\��yӭA�-Ĭ>VT��;��:5�<I��o*���G�o=.��ӫ��ǧu�':�C�;����!v��03�N��@�z^�"H�bs;�;�5�F�~�\����Kŭ��^m�9Q�fQF���H��i�,{�g����Y��G{|D�J𸟯�3p�6/�m���W��pR����.IY��T�� �:��m8KC��[i7�����t�����w97v�`�C��JN1Yʦ���_N�*x���+��c���\l�D�[�1��$�2�e7�kz������ԟ}����n�bnf��X�j�~�
%eQ�Q�����~򸶽�#@ɵW���|%
��7�RBl�B��m �Q�A�NR��ߣ�5ٮ3j.T"���||;��ē^�ێt����fwd+�O��iXw�q=�_6.a�3�r�Orõ
6����I���PfҚ�w�nB8�1q��Ҹ�p����B�,8����F��O�=鵵��帣Ym8^�`�j�3��K1�k�ߘ��ll2]X��GX;g3�WȩSd)	�����hP�됬3���Z�imk[�,����]�g1v�I��̢i�2��Ȭ6�Ne��v_:��uq�;�S�-Fd��v�8�諭����A��Y'��?|]��֬��k�W�:֎%�y7�������U�&1�	��ui1��2�d�G1���?\�����F�����S����s;f�&�F�6�\n._Cn5�,��vD�!�-nߌX�*����{U�@�����<� ���G7]k\9�{'i��W����f+\�)b:tr�椵;2e{k����ܛ{�_Z��c�;_e��;7Q���3)�o�1�Ѷ;�{��w��h�с/F^r�������r����ո#9['3���\�˔vR8�����S�[p%0�0��O�R�
b����"Ͼ�rޏ����n0��+(�;v\���:��k��U[��*��*�wZ>��4�U#�3�i{Z(���v�7 ꯧe���U�wQt$�2�D�@�fnG/��|�w�W����}���sD7��5Q�#Ӷ�e9�FZ���8a����+�Sn����k-IV�����#���k΄c�w��|����}�S���A�5�RFGU�VQ�\x��eKwxdٹ�%��Ҩ�5q�6GeC*vD�ޠ7a��]N�(��֢ٮ�sb.U��A�ΓeU�}�ܫ�*MP�gg(o�Z�Q���p�=9����U������i�&���)Ks���&���^*�����_<k��ͧ��]+!���+z���>�9�ك~�F�Y
������n7�:oHj���;��5����t9��0��P�1PR�P5s�G:�qڎM*��qZ�??w��iRk��&�5��1G:�)W�A�4�U��[��I�X[�[�.��Ox�m>7[�Ҝv���7��6�W�<���c���5)mN��Fcn;r6�C�/eK�R��[.����bk��kW��#�إ�H,\���bӺ�R����Qv/yi�/-�M�'�N�E��)̃��=]�׳�X@z;�w���5�}���闙}O��x�ܬ|�Վ뇶t�<�˪�c[�B��f�(���{�*޿��tS���G7�y/|��(x�s���+nc�#N��3/J� �M?[���JV���R��_	'
��٘_����o˩c�0gY$E$����M��Q�kL�N�Wn�c�����T�Op�X	�p��Ke�]���E��WT��:	f�B�����;C^�fUAckO9Rb�6�������y�{7;ћGk������̢�G�]�:p�y0��~zk*e����֔f����s��[p�޾͟��ʎc0s�v?���F���y������~�g0��N��د�&źonv��+齳��������[�c͡�=���$��4t�T�+�.����Qj�����s�5��g��ꬷ��+ĥd���a�}a=�1k7���W�����6uN���=u1ww�-���$S�0:`�?@|��RW��.��!�{���̭��y�)�yʯs����-D���A&(jJ�1Vu�J|ch�UV���td�c^�E5�=\���9��bܯ����KE�Md��Pu�RwG��݌���]�ҿ��K <�M�(�qॐ4vusM�qI�e��܊�]957+��>7����p��;��
rѪ����T��hb�aw��t�m2C\�8�$��������7�[u����	���[OCT�ۤ�Z/�N�����:��ּLw7
2���f�miQ7�vJ�!P΍���D��`�hIS,C'�Q�%僰�3ҕ$TM���ﾪ��ȣ���y�Squ�y����n5'���M4�w��k��y.�;2zk)��mKL�-�D8��/a�ܽ�ͮ{7�j#S�pک��\6��̓\_-�p�Y#T�m�/+��Y�j���\�~}�7嫷�q���{��c�h�e�#ޏ<:'�Iױ��!{A�=/��1��M�>��;{UH��ỹ�#��^Od��s}�z��4iR���ĽT��3�2\b�Ȥ��a3n��J'-�E6���f�LT�̺�ҹ��Q�uk��H��79�s�.&/�3p�6/�ީ�ɼV�dώ&\~�z��}[-��3��uѨ�P��+�b��I�ϝ�՗ٹjN5��_,	�n!)���L��~�D첯��
�)UZ��a���� �;�:�@؛獾��'��ި:y�T�I�b��u{غ;f�V�evP���#�{@�y��8�+�L�R묏K�y.�����GAc���v��]H�����Fİ�둦�h"�+��s�*����9|�gJK�i7X�)���Ŋ���F���
�R�w\�c�Iv���gw�r�h^���C�S�}U��|�W�1;�5��ɴT��ޅ�9gA���g�A���<�QeK�A�6��76e�ea~�=�4{όsƻ\^t6-���O����웅7K"p-�{d��FÂ�
[̀���O�ඕ�w�s��ECb��,��}��l[F�(�T;�j�C�)����Z��&���8t���-������xޜ���5Xe0��	����Kj�Ru�ʄ�̾!��Tg^�g�8�:mw� NZʱ=�l�Ȗ�~XT�s;��͊��x-�u�o�T�|����c�?k�&9������TF�n�M�=M내���K�9�7�5�/oC'����)�y`[�]=/��h������f��\d'�E�s9�j��M}����R��k�!��˞ti���H̕� ��V�y�q;V��z���1P��r�?��PO/9����3=�{)�#�Oqm�mliZB�����A��`��E1�	ĳ��m)d�vpc��#�v�ө*բ��g0��Ѥs+��<�ۺ�g��'bd���� �Ǹ�X����@]K��8�ջ�m8�_�_}�U-�땪y/	�� �d�Aw0*��ۈ�W����ڤ��M�7�m�-@*nVb7�Y{�Փ��VQDv�ݴ!Ϭ'���V��(z�D2��Fu�Qԯ\��f�n�{�;o�=�#���(�ݗk*��Z��g�[r�ڕݢb�'�Sњ��JZT�Jb��q��y�l�\�%��T*�2���ۺ��RQ*_�r�ˠ�%*5���p�\=k��ۃmWqw�#���p&n�Nr{�o�����)��4Zy����f�+��z�����t�ϷV[���Z4o5��YՉ�-�\|װ�f��.��_AW���p�{k�����P��`��-���1���kqŞ\/��BT;)�F>�Z)ί����H���P4
O�>�Ku��vӍ۹��s���@��i���9�m�v�1�h��a�^�9�>J�F-S����tT3\6��i����ڍ��Ϟm��M�37EJ�h�TJ�Cr�m�湺��fl�ē���wֶʩ�]r��{X]֞l�L�mK�����<}�H�y��G��[(���ٵamI��*`J�N�;���sf��U{��$�8�U�g���+b�N����Q�J�f�-��2����bjq��A�DO�Z�\���{�t�;��wz���=܉���^b���N�c�=	��Db{p�J����2�j�[����89�'����w<Q�XZ�λ97VvrU�sW�����/9� ��R9��g��WtY���y��9��v�[ҽ�0�ۘ�6Ǜ^��M�e?�~���=��3u�{Ôq(mk��U�o�9�D�8���Q/�k{�iѾ�c0*�w�!��ϙ%���_4�a�qz9^��-��I�n��=���~(�߶_��:���6{
	�ޕ}V�����_�]+�د�CYm�����:��Y�0c/��'2�J�EN���~����u�R��[ˌp�\=rf��F!�%�<�ƮN�o�@�܀���0(��I\-��[�_�rήaYU&v*đen��GAX�\˨�Ι�j�X`�3��e���1Q�::�Yljُ��!v�RU����kE�5��WM���9�pXW_\�\��Y��zJ�@Nf�!r�n'�+U%]\zk�i(l˵�D�ç�}�����ҕ�?������OLC��S��F��q�Gw|�J?@I���+�c�o�SuKo�^{�NfB=�M3W��N3i�sQ��:a}�0X%-�O��`�KChv2��3�z��m�Ұ�Rσ�й�(��$��S(�R�9ҋ;˦��+���O��(�v��F)F(D�6I�ri�K�q �P럮wT�e5��5�M�M4�wˍaB�ș��=]+�+ǊSޢ'�Øm@w7+wsk����O]3�<���$Rw�۳��vx�I�w)x��xE���ˏ_�moOL�=��K�8&�k5K���|���ا�~��4m�-v|3L��w%�f�����&��	���F�s���Ր��O��}���,��D���U-5���O1<�_ќ�r�;�)�q/�u�q��}��1�횲�ړ(uw`�kv{��U�F1�5��+N�a��Y[ڽi#��n�J�����K��>�!�57�Գ!��i��;�$aj��_9o1VRN��.�u5	ƚ+j�1k��!ܜ�0i�d�+��7�['Q啻���91<���6s�0` j���ӎ^�����nEE�ùF|��)��[{*���y�Sc�<��]^4�>�w�s�
n/hժ���W��Qi7��D�sQy'�5X��Uc��^��g�5�T�x���.oI�M�����Qo�����IJ7��嗍��t��ި�C��0Wϕ��C�f�~T{\��\g�)�V��VwQ֞w��zw��Kb�d�X�{*�T�\�F�j%Ib�u�:�K|h��|�����r����ҵ��q���{7��q����(kk2άO�6��nB{���|Ll�jc�{qj=L
��������h1��N�z����M+���%3O"��6tR�;گ'�fT8�L�0�%p44���H��)=��u-��+3�z_2�6(�f�K�\��v�
�L��l��@�_5ى��b�Դ�'Yq�0^�F��y�IY-x���؋
�[��:��<VA��ʗk6Cv�p���U�WF��E�Ղ�Pڰ@���]�:l�:���s���reX��Z���{�\\��POΒ/2/BD�k�=&�+(��y�UƮYN����v��hř):�R���Vc�����ޭׂ>�n>
���՞�������m��R�~o�0�}H���� �����@ �RN��p�ݣwh3��B̫�-,��K��:�F�h0h�QY(3Z�Dd��s�;Զ9�j<xe�F` J�/gz^�Ҭ�� ��R�?:��4�K^s\�Z޴�Bf
v���Z�re�����>ߑ����̡RCy��:�O6���ۛ0��k,�-�21�i�&���x8���0�*�{
�_��n�itbq,���6�`Ġ�t�P�=D��S�h�D�%s�9���{7��tj'f+0���e"1��vG�W�-�(��ȧ����� -��$��fR*�%:Νr��7ْm���%Psz�����C��֮*�b}����-��A��adue#��]��0w�%�	#�ٺ���.�L�"����0����\�-x�ն7���G�j�l@%��7���V_U��M��ғ��K@��@�-��Mᨓ5��<S6����OUC�"����RM�0=�%Z��*q��8��\a�s~�z5��+�̩�[�弩!�E�g�C���eKi#�P�הP����S��(��f ��*'�r��7#ങ��>��{$ z��(P�1�=K0�{�s�<6��çl#*M�1Ս�RTT��Y��z�%����h����3vB�Gn9x�ks�����3m�����!���m��X�>�����7���.g�ߥ�X�8��\�μ}���8�l��$�RC�������͛f�No[Ӻ��
��gb�F"�D�cG�ws�b�ϺЧ�x�nLΗ�*\�tѦ��XΫ:��Gi^���z�5�ԡD�gJ���Q�r�����V&j�WGK6��P>��V*���������ţn�
�p�ڷ&�ңAjM��n�xǜ�p�M`�p]Z���JQt�*a�7"�E��1��a�-A�t�+v�Nv�f��'�e�ٴ��u�
+�����]���������+�7�h�ܫ��R�s�)��ޘ2h��#�Y���RaQᘹ��n���ٗ]�(K{��:��Mj���}nT���NN�?+��gaV��e�3Y]й����=��k~��[
�u����l���
�*s��Y�\���$2qG�b��V���0��AR݄F�k�vn�&�bugq�Fڣ�M�y�fA&��� 9{�+��\����X��t6^��ɔ��GO"zweS�ܚ"L�C�& 6���#� `̐� ��c�EL7v3��+�P���+]Fc{�K���Kc��R�놘)��)�ap���!��̤-����5�$�%,,S2΅�L�2�EV�a[wC��Q� �Q@�AL��i*F����$�ͪ�LB�(�-��I$I.�I��N�DIJ�%K��
i�5J��
�%�$^�4���&!�4\���[D)u�d\�4�K6�Q(�亖F��mʹ�kq�(�Z�)��RЊMRJ�0��$H��QG%.�:������(E�5%��U*�YYE)�a�Cj����e���!A̱�'MK5A"4�%"U����PX�-*�%0HBR"�Q��TX�Vͪs���X�U��4�I)
GA�Hꊊj��Vj�H�	��H�	ĢΥ���dFӈ�t:J`�����.�X�,�LH.hbZQ�BI�PHV	r��Dj�� ��9���5�fr���j諠�͞Ί�!kΕ�OlE��q���� [����Ȧ��䀾�͚�#H��h(я�����}2B�x�W��M�i������n5��*~�vD�?[Aڕė�Ÿ�uO&{�ɓ<�w���u�j�V��Z�Ψ{'k�s��^ �b썮�%�NK�Rތ�|K���|;u5�X��R��k�Q��.p^d�*6J���o�c���$��'��Av	y�&2�;S/QO_;�ܺ�UU6�i�[�m�ߘJ{�VUA�r���C^r-��.���>�O��&��DVu�6�}^W���/_���.F�+(�;~�~����^ѫez�X�֩��������e���4��I�P�sٚ�/l�E���g5��ar��7��l�^���*Zn�M���'���=QHٴ��^(�]����<2��W����q]aT�F�7��ǡgCi覺:�����"E鳳�\��\���'��j�K�[�+q����&l���;�}@��gV��n��{#!��"c���I��oD��)��d��I����~��y��v�4$$��Qd��9mv%��ʵ+u��w��5`_m�']۬�\a��r\x�ͭ�+���4D�(�z���%�S:�t��Y�����"#��;�7m��[����ࢂZ+��g�gTb|C}�Y}y���F�6��i�o�y��zτ���*J��^ը��Ps�8�Џ5����U~��}˔:�ػ�'�H�G΄�. ��l�O�1�-zu��2z�R�$��n9�����l>YJ&y�y��,���h{5c�9%��Ja���"S��C}SP�`�&�]���!H������#h�"���M��)7s�[�Zi/-Sz=�;�1���,�ԧ\<�/Cy����D��QkpfuD�̸�\�w=�ܬ|��B[sh]�����x��v?r!mC�h�]/��uU�M��}bV���І]��!vwy[��%o#�:�N�8޵q�Tv�?^Lw���c2�����h4�B�q��ej<�)�
��k�"�
%�����q�6�����h��(���8 +�ݻ��z�R�X��XNڶ/�t"��fD��:�����ڧo�hkI֎3jeb�#�ey��~�&`��k�]�}�9k��H�/mb���;'B��
ע������+�9�+�3�qgj�/FAvw)�T�[����U}Ec�Sܞ���DNe;�*���F�G$طM��*���/(�;!�ٚ�Wx����.�Գ� �S�ƾ��	hr�6Z���o�s����VB+Y{^�I�+;T�ق������+�"���-��8k!9cq�A�\u$6iv%W���c{f��G\G 8(��Ir�,��u9��+}Y��7fQ�Q��I���+���S$�q�>�*b�jJr�:�g>�Rt��εu�!-����8�lV9Fc��_n���y��ж=�,�f�է�� cK2ί�wm�M+�;԰<�Ь�\T"{�k�1vh�����oWS]#�Wqa�nk��\�v����5�h;A[�B�����AΗ}�P�|�����Q�qr��JY=����h�����L:ך���/\
D[���4�U�]D9k�E��"K��,4�[Jyy��+�Ĵɣz�t�&�GѴ�]�0!`�N<�jApx ����=�jkeg��,��4ݽB����G���bD���u���.�o��Nі��9v��U#�c��J���+�Fc&a��8U�����EiO�}|%'N�ͅwڍ�D}	�=�)��ͭ�F�Mƻ�WS��:E��}[Ot���эOTǼqy�v#��U���?{Y��^�|�[��(A�~Vc���h�ܬ�e���k����.���O��m����2�*8=[�Pz��v�5���o��d����'-�R��r���\�x�>22���`�)}�z����:��Ĩj���|ͪM��������yG�tZ��/�u�g���U ��
��urr6�%���-������p)/R[�����g�����#T5e4F.D��g5�Ǯ�C��;������n���u/�έq��/5���)�ޡC��F�|�~�"��vX�f�C���C;9��AT�F�֞޸km�Z�q�7��x����ʗ�ϴ�Hȋ���ׅ�������ܷ�7ױ��q�ئV���m����MX�=\=NC�6c��ܷ�A�����s�����V�I�M�&Iײ]�"��/��3�F2�T��H�h��R���vWW:�-^������C��^U�΃H|�%��V\�z�����/=6K3��g;��@G�q�f�ٸ��_U=�2�קy�m|O�V-y�ςΨ�O��-�@w�q=�Z`].�c6jr̾��ya8S��>��4�=���\�>G.9�ɥ8h���r��<��*f�p?��J�����ěV�Pؽ���J��3��XŬ-;gc.������O�t�6�;�ƻ�pT�g������7+v]��Mt��vu��+�ٽ�.5-�o]�6�jsM��p����t�[C/2$hwjT\*�Qk�v����ļ��7����^�c��x�t ��^�������D����jc��y�K�^�u�X�9K녯�}'�I�&�]��T��<|�u�$���!'YO�����U�ڙz��ˊ��:-��R!m�j�s�5�-H���}�B�8bUy=p���P^Ҵ�zQ4�^1��;�՚������F��f�XQ�[/ݿr�'��̟���g���2�2�zۖaJ웮�9;Ӗ�k�^�kI)�Q5�ʵ����/,��v9o�h�X���A}E��Lٜ�;�~������_x��!=�ST�Lϊ7�p%L������޳�nei}O�0œ!�-��]3:��Q-���5��V� ���������Y�ތ*}�1Q�7����n<YZ;�]��?I��_b���I��ҧd���ǜbt�#Kb��5��}:Oljƈ}xq�1��Q^�+۱{^��u;<U�]a��ok��ޅ���Q9����]��5��ءs��*@�f���Q-騂���uO
"�p��x�^
��[/�P��邠��T�"������cs6q3���)GE�]��N��փ�����ڹ���w6���eԐ�ub4������}ͥa޷���1R3G8)dN]���nzE�oJ�]"��5���c�Ϝ�o��q�k!O!�����O�\JM��	�����B5�]�'R��oRڍL�o�ZL�b����5�4�F�Z��V�V|���r�<����Iym)����ީ���[br�ۊ��cRA�J�J�n��oC�7x�TG�e=3o�ѧ��c�D|=LF�:ҏe[�q�c(��-�c�H.w��JN��g;��pn��L>�ğ	���W΁f]L�:����k��A�<�(d��r}zd����Q�
 �U��}뎪�U��g��c�Ӿ���a������c[D�����J�[�uC�{Gti}�d��_�i_��]�k�;#`U�/�QlG�:֠θަ�
���7�[Tv����������֦��^Gu��_u;�/��&m��
���M���kz�;6~�g+�c3g$r���5���@��t�*���Q[�6-�{j�v��qd��c9x�W��{��r�)��ƾ�P��t�#b��e��<u�1��gl1ST���Wbr�ʪ`l�N~��Z�ͬ�ac��vy�[�SP*�k����zz������AN�ۗm�@zu���}��9A���[�q��Z��G�	�?9^��\[^�;fIYl�?��BL'Rw\]r��#��Cs�f�ķƠ��a��N/:>l\Ôg�".�K�"�0w�����Uε_F4K��M�U��{#<�ۓ��NZ����
�J������y1"%ªQ'�6_i�C��gGM��ܚ�G�/kS�W�Ca^��J���n*�P�:���nPǢ8��lS���ǲh��V��
T��M�N,a�M�HT@|�B��whM%ޥ��
h\�Fd�ܕ=q�t��;X���`��zW<�����9sPքôn�t$]Ԭ�+���9�糗W�a�]��CnnV����u&�֋o�hD�\��5�P6��unr���O�*7�N��-U�o�D�-~X~J*��%Vؾ]{}�Dsq&�Z�I�w[�U5)�MƻWS�Ȟc�Z�}[Ow��K�|\#U�֣��祿/-ܛ�Nu��Þ����GU��Z�R�x=�;;,C����Qg�vZ�÷SQ�\��Ր����g^^O2���{��`�V��wd7ퟆgs�'�ˈ�Q9o�)���F��������͓���ѥ�}E��]�Aw!�����������ڤ�X�v��]7�&^����_��|�+
#����AW ꯧ]��P��t��t$�o2����[p�pf���H�>ᶴ�WQ)�dv�9Q�@o]଴��Ja�ڶ�I�o{��?��C^�8��*J�N���V=�7nG�km�E.a<#e(�ĞF�/Ļ
�-]�&t4��W8�0�.P�#{�J���e��嶢���nJ���������\��l�m����w�<�'e�;V��EX�w�o�D'}��Jyc����]��t�p�V�u�Ct?U�nw���T���u�:����O:5�[oB�y�E%��SMe�yk��D�,|~�po��������ܷ�7׼���زt�oM=�[���i���q��� �|R�Qy��;��-�aޭ_r�V�ERC\cN*���9�WPGh�S�1nmԔ�C�ͬQ�t:1��v�E�Ȇo�+i�J1v1��\hT5q?B�g�r
UA�4��䲅^�Ó4�pG8��J�W�'�NTs�-��x�A �-eX�ڶp�B^�Y� ��;m��n{���R-S�ƽ鹵S'�{ޭ��]�V�Ȝ%��iR��y1@��q�U�[^�$~�Iy)�*�=��k�=p�Nӹw5Ҭs3S�=���oR��݌>V���h��'
7�s�h&�O��I�Q5[6a�J;ٽq��L�@��{�+QΦ��e���s/ӝ�N��5��\��c�ۨ���K�=Gu�T�qN��x�'Y.�u���,�o*�G�Ӗb���؛H�u��9�G!~�fsKّt��)���pyN�D����gË�T��}�Ç}U�.�]����P����
�{��c-�x:��8���qd���708��7�}5"����}�����Ƕxt��J�):�`^�NOu%^�o���޳^ވ�F�+>(�ڭ���XN�$���6��/?M�4Q����alW$޺oS��u��휯��/? �N7��{ᓀ�|����|]}�ҿ��*-�Yp�|�<�i�r(��V�e7WSR'2�oi48.ʧg�����%*:��p��Cе��^��7op�%ru3m�
<�ࢇs45%q������iざ���owc��91=����j�X�tH���*�P�k2 ,॥\՞n\
��v��ԦU�{z·۟7��Q���P�0�ﾋ{+T�۰�-U��	`�n�n�j�W�!Sk���B]����8x�4�\�4�i��q�o�R��6j���^�B�p��˙})f1L����q�mm4& "'�]�f�+n��.(�l�fՀڹg[��/S�*Q�O0ފ��C.$���c�%�(.����J�R��xҖ��NX�;�f��ѲByPm��E.�pNڕ8��N٦�ݽp�}ֹ�`P�up7u"�e�AVel�P|��*q���!.�u����m
�)�U�a��:��>q÷><7[�c��m+��f�o]����K7ʻ���C���5��\8�{�ΝV�kMT�-n.k�:zTީf�B)^i�VXv.z���|Mޙ��fjgYt��R���{B��I�D��wV���M�*ChC�G�a��x�J]pj�sn�ϕcwH_ȉ�cr�[��%�b��:�8X��h�kk�����R�{q��c^/�e�&E,�gF�k{����Zܼ�Hҋ��{��U�3�������[��Wu�\�+9�4�-���xD]�B���h��I���(��% ����DgEv#�iF�+o��'Xo��m=ע��o�饹�Jw����0�k:�a�i<��<�p�1ⓘ�3�7D����uk7��Ô��<�_cf��e(حv�ӹEȜ�U*�8��(>ށ�{Dǜ���\dAF� [�����S���ľ���t���+n�#O�m�tA�v�6J8��7�S:���Iv�.ˎ\ٜ�}g��.���б�lF�me����oiN-��6�!R�=<��]�IK&c�hY �^H%m�(%��P	����j}��5Q�w�9H���e�:��:2,�P�O=+�)Ͳk)ʘ�y�.^X��j�t�EY���ǉ2���Z&@KEB��x�]M����r�֟L���|�(���}�8��ҝwR�e"'(J��q�v�tba�[�؂mչ:K9S[|cƍ�� 5�"T:tRѼ+ �t;�fE+����������Bh����xݲ%�Y��+{���*��ȕ�=׈���h��a�8�y]}��;K�%g5]n��I�:�����0��-�C`]���/�n:N���Цp�Qg-�r���EC}��	}����BD)�-¨a�L�).���i�ú�/��'vڀ�9Ƕ�]���>�Æ�[B����w��-�]K�]@lJ��>�	��*��*��������&\��)pJk�*U�kC�Cߚ��E��Y,��W�z=(�;��WP�&!�
��Gc��.Gj�	4�;��T��ȱ�޶p>mQ�����}�୰��k��nc��0S�s"W��t���q��4�J;�Lj��c�ƀ���p���5Ы�ZS��M��z��P1;F�i��qS��N(e�� %��9�P�Jc3w5��7��yN������J��E�TP�el�-��	fR��PFHUXY��4*,M���6��AiK*�4٢��%�QQ��fQJΠ��UdV�Y�K4�D±S
�����̪�9b�V*t��-.�X�Ȏ��U)�Y�R��E�d�u2EiIGR2QH�J:��$%e�ET�I�Xf2�YhUY�A��Z�"�DQΡH�J����2Ԏ��� ���*�,(�*2� ���T�*�aeE4�LI*��:����2*��Ē�"�X�F��­f�[��"�#Q
�fDQ(E�F4�#K�"ev�%��\*�*�uZ%h�(�[TB���Ԣ��iJfY���j!�6m0ٕl8ZX�kZl*���U�5,�"�.��*���� DH �@��;�B̋���*��{%s�[�t{k�Gj����H]��]it3B0����S"s^Ex�W`l�*�Z�����eh�0�V&z�}�:����Ҹ��g05p�Z���+;v.�\ļu,�����nu\�[��I�>9\��o�b�Md�`dS������ٯ�����'m_]��;��Υ��m��\�&�Y8���24��+�{0+z��q�DL&Ŗ���*�#K�O-K��ކ�����VL���qw=���-���m�K�Gj�;!���A�_�M'�Ž��[��v���Y��)��}\�ߢ��^�c�����}f�gT.z�;i+���m=��&�뵋���!8�ξܮa��7�[Tv�8��{�%�����9|�"5��������������.��ļ[q�vk���~fnV�$��:U�<�=�w�2���N�����alW$ظ{�#5�cM�g{�O�3�㷊�mA'���R������geBX����P���?�%�dF,)��z��=�R-m7$�a��J�3lc7LP�	�Z/�=2=~�.y��ZSya'3YE�V�\�;L4ڻ���ֶY�eٹ�L�M��\t��v6��/�>i��@\4�5ɜ�\��`E���rU�!�9��d��z�s�e���F��<�|��Xp Ǳ��Y&�k�<����p�'����)D�U9��m|�{f�����|�F��(ȕ�j����t���r�	)�v�-<�b��m<㈥�
1�>�*�K�fo���s͑֔eȋ���:����o�÷ڜ^t6.a�3GaAi�Y1F�v+ky�}X(3i
�f�_F.�iXw�`y���k�T�n�̣1�v�
{�uqvCT'\h�<�j:�=Ȁ����+�5�e=o���P�qFV�,�������f9��y�۟�V�����oRz�{(Ly�.�;��5�׼y�*;��ԝ�1	��l�+h;��V���\�]�����f]�V�r�P+����MB�
Sq�T����g�-m�CY��9���ݏ��{~�NG��m.�e�k�����:�ޫ7�1ӓ�a*��"5�A^Z���0�2i0�{h>�^u�jܻ�sB�	�&����Z\K*��(�>���R���=���w)�
�X�w�JR�����,r�;��- ����LG`ړ����F�"V�s&к�Q�E�ߐ���#BR]h������'E�U���ƩIG_nW;�2�&u��������3��1��!���c�=���oJz�q��e�(�|��)�q/����(l]�'�uuc�Vs��®`>U=��T5x\M���-��gh�l�Ri�C:wΑ��MH�;%���9V�^ѿ-�%�Þʋ�u�]��(�^��h��'M�\��l�m����r)g���3�ж�d%�P�G_ղ:������f6��,f�����wH�7E\mOM��g�ύc��_ب:��ִ���[y\[^����2�����y �}y?w#P5%�m��Ơ��|񭕞��3}[�X9*M��߽�rn�PR�����Y�gV'�I��(m-�{�qRf�f����fx�U�����:��ymc.>L�i7�^�N�u�v���,RU(�BO7}��s�2f8��SDƘOtۂⷋ�w:���<cAi��i�����d���[�e|-�Qũ0���3S%�ټU6-��t���u��M!���z(��[Ndx���I�1ȉ���t,�G{��k��w|���\��@v�CW
Q����@�)k�Y�໒��G���*�5s��2o�9����9��a��j�D�r0
t���N�զn	�A	$�~��L5]��¢��S�ڙ���6�]�,��dI�-.A[�%^�]���B�}����n�|�'����޽��yg�2�J�C�LY��R��( �s �qU�����Oc�{��nV;�R�h#`}7��.���r��י���4��wS��w�I�S�:�q�+�(Xf/ArB
�q�,^y�xO/9^��Eh���mr��n>չ5�����3Y՞�<�)�
��o��=�ވ��,��vK�t!¹��箠��Fh]+"\��o\�Q��(J��U��_rM�C���v���h�f�D�1/&nkw(�Q�+�@���'g�}�ʨ�N���8}m6��'�.��L��x�WX�׃Ch�V,��E��_gY�Ȯ�җ:l�iɏ/xk�9�n����;hSz6��.Dz$*��ᦣ��۝[-uj\��n�I �)ٯv��VRf�ɒT=�*%�h�suӾ	��铕�!��/7a{Q�8�Ⱥ��m$�Yʦ� >U;<]�WXU)Q��7���@��еv&
��=��w��T�{n���Pb*��"����@Ԗ)��1[:��
��x-E�Qky��9v>��b���/�dZ(o5��9�u_(�\�[Em.�+�Wݥ�o���ky������BSߖ�,��m�gg�d��v���B��F:��J����s5�*���9��$wOMFd���rz�����7W<���Dc�Ϝ�;����2Vݬ�c����7���Ѯ�_�+\�e%�z��je�7�5�`����$�[��,�
�v�1p��^ �{����F宬S�R�t��)ϵ�Ma��I9��3�G+W��9zҜȜ=Wқݤ�#�l~�={YAL\��c0x�J�a^~�k��yk�3��y�uS�Aﮄ���Nx'q4��6�8ݐ=��: ]=i��A�\�4.f�{B�ope*on=�W�V׽@},����r�IŨ����rW���V>�=7j�^��yڷns��U��>�؛,Ԣ�t�{�gE9qq�&�t�&L�����iU���u,:
d��YWෆ�o.u����8��p��^Oy�c1cڼ~���INs�ޫ>z0��Kf0���|�Ԧ�ļ[p�޾�U�j���;#SN;)z�e|v��Q:�`�k��-W�[�a�x(���3Æ�e����[��n�
����P3��;,�҄����^�ݿ�ldT�>��I��O���W������y.�P��n,c���
i]_/�l:��\c�L�r�[9ՏOv^(k���i�ި�C��T�Os�G����6׻�os�GmQ>zjO/�5��-�y�*!JU(t��>���Ƞ�'��c�!�����w����O����۟'�ضQ��g-�HU�ؑǮKQ��j��� ��CSY�gb���s�;ԡ݁�^�������jJ�ݵ��8eʄ�CA<�j:�=ςn���+�4""�m��jyأ��l�He���b��U��J�5g�!��ᜯ��b��Y.�cQn�7#9�t.�yc�G+�ps����Yx`�6qj|)�1��6�7�듗b�q��'��9�P:�ئS�r�sl޸yZ�TO�j�$��k+F���R�O!�9��}r��JY=�QV*����=*�R�i:�2�:��L;���!brEDr ���.V�Ң�����^*��] +&{�"�S���5��Kn1��tC�c����1fc�JyStJt���׫�D����������{Y���f��^�iB�o�z�X=Wr(�e��4km|3Dͼ��\:�7S���q
e�L����̬���37w5S�){73�/S�]�,��'J)�ao�s�N[�p�6�݁3�	sr$�th�X/V��h�S凷��A�/�ޟ�9��Q��O~"Tc�����6P��~��Y���?Y�{��|�(�ղ��CV��^Ѕ��i�{�nm�����Tf�G�1i7���:�kr{2)��쌜ˤ�]�d��އ�M���J�sǥ���q���]���Ol��
sJ����h u�eϊ�/�O��$��5�h9���OL�z����4�+�k7Z�l�x[{|��o�D��3B�
�zA癋OxF�M��7ռ9��5�A�7�LA�cV���8�]ve!3�d���+*p��!��n���4G ��	��$!�ԓ����4~�Q:��!��F�Z{z�zt<庚�gZ�d��}����b��0�3��U�����Ao��5է��Յ5��Ȯ�Ԯ�C����)h���T-��Nϻ��3	[���'��e�Z�co{q=�_6.~r�� BQ�s�ߢus۪d2�P{o��-@bq���6��o���
��&#1�8	F��%i[ W-<�d��m7�{��o�ΫZ9Is���p�w��Q3�kI{Dx<�47�P�qc
D�wz��9<��+����mF���U4����c�V��ג�R�'��S��C�
~������qG�)ym)���b�{�$�$�����N�^�� gG� ��*��ti{2.�s;��y�(n��JEO9;;5˝[�7W5�>��s1���b�y�b���.�:�V�xѸ���X�|RY�Ŋ���Й���|_;��tt��n\��B��,��]^��g`���C2�9(��=�tZe���4��"�@t�S��{&eR)�i���M���Cγ�rsr�tQ�oN�v�B8}��w��% �Ť.�Q%�=Nީ(*����g�<���i�|Aߚ�T>L��N*7*D�#Q�ԕ�3n�aQ6�3j�aͬ�滺����E �+�k� N�&X�p�(1�Tj6�5z\*�����sٚ��oyK���4����K�<s�9ֱx�_X�+��ب�e�m���<j����P������+l����Wϑ�����JTj57�7B �m^����Z�=�0v?�On�P(t��
�;���+�A�-�����rqqG5�*�;ۜ��P�f��s
WP���}0T�s�,��m#l
t��rn��=���Q���t:}����r���,�COen��X�h���E��SA�T�@|�`YՋ�W&�:����
��R���_Jٱy,���	{PϨ�Y���c���|����q��t�@Y����kq���V�ƥ�� Q՝r���
�z�ƺ����+nW)�q�]>���E�G�&�s�-�M$�w��.�)�f���4i���u�O�r
s��za@����\��u��M�%�5d]�5L,����k�d�N<1��R:X�Ѣ��By�2@y���8Ja`<�u�\�sq�����mje�}R+��-W�D湞�h�f�7k5:����r�U����xF�b�Z��m�A��^�-��_w����&�l�y����<o�B�ו �l�}P����+��^���R�Y��	��b��\�h�}�/���߆B�W�ϟz��)�vTO\G��{�Dc��p�x~(].�~��$_��sƢ�#}[i�5/�㚥��Ҩ��\׸�:�=����'o�Y��͓(Y�W=㟆�������=<2жj�Ό4��9�,
�^Y����.+լ�G��9_�#՗:`_S�����4.���Q��Ԣ̌<Mܱ�zA�aא��p�+���i�z}^&�^ѽ��]�x��s��9�|xO��ǌ�(�pd~��^#��S]U�7�[�����/��s��]*9(Ō�wD�;��^Y�Có镎�ܥfOp�=��`u,��}jG1��=7����z^��*}�}I]ǐs�+}#��{�����^���X6J�,����_Cs�R��,H�3�q{w�xV�ƝOݳ��2��[�	�eۏ�o=y;�mˑs�3x�4@jK�d��2Gg{yEF�˘�v��+p����d[e���{ZCw]���鶳��'G"���1F�����u9�RA�j�l��v��
ڎ��8�Y{h\��A#�6��o+F����)kM��=u��U�_J˖��5
U ��.�2�����z���Rĩn��n��@�"�&+��b`i�$�ih�o����kM�ׯV������»!�xybcҜ>�\�e��V�z�ӹ޼��һS��4�l��\�(��u���p��s�)�U�ּ�ː^N�t�bu�N�Xι���&�G��H����Sz��>�Z�`��c��+y��b�t��c6�D{�d���o�m�!qA2���L���7�b\�����M��}n�-(�M�*�������Z5!�\a���M��5&I&��u��:�-�
���9�E;��wJ�q��F�s�&��jB�Ńk�7ͼ/�q��p��#�ڛ�ˊ()�ͭT����:{�ClJ*Ѷ��	ٛ�1��D"v�B��l>��+�f���Ӛ�.�TD����bѵi7T�:;��!�%���P��������R�L�ڃk��9y+�6錼<]b����{�ū�Ɖ!B�nZ�,�vK�p���H�lo�E\SJ��������u�Og8�c�YŶ�;ff�H\#���se�d��\y�8ܭY�r
6���ڑ���/��]�u.��f/T݄bu/��Gj�`3o��'�e�AbWg�!3�a�у&�iE`VqbQ�h�1J�Z�s�(�G0�-+9'A��t��;0� �d�ֲ��w�$8[p޵�L,��%T���2do�{O t����S�Օ��.Pa�J�\�kv�T�����w;Q�Q�o�,�B��s��]�-K�YMu�����iq+��ƅ]��V�=<�q��i0������F��$�sb���(l̲�bmɱ��VMۡz^�v���K�W;�X��1���I��w�uB�n�ǻM=�����1������(�� 
E5��	��&v^�; �-�����!ڳ������G4�Ȥ���i������;���In,�F����Ӫ륳�_&���%N��L�j����\qh;�U	`V �U�&\|-2`��E���8:G��m���ދ�6�؅]*B�5��uJ�V�Or�Z�t���GDIm�x`ʨ���V�]!0�*���6�MDѸ�:7�Mr��Y|_fN�J�C ޺� y3�^����Վ�G**t���*F�c^�Y(�t�[���/c�#ʱ�i[YH�/���5^u��pLwkTyʐ\�����
�s7�
9.�]���Ex�(rKr'8�ț������ -��v-n�k>���>i;�(�H�2�I:F�I�2�-5��5KT��Q�2�D\�E�5
ċH�AB�Zr���I,���˗(0���Y!Us�4�d�r�Z�4��Ȏ\��J�� J��:��$�ЖBd�$ʩ%8F\�Ia��S9Y���3��P�f���j'B��$�.�b	Hbj��A��.!��Z�Qi$��ڭ
քjERZ�LU��ZU��\���kS��\K�KL�2��5�b)��%�T� �ip�I��aEl�1�S���0�5)U�iB�]I�ж��bja$dVF�(��eJ��3*���j)�+6ʳ2T4�f���i+U=��XaQJ%]kR��22/:�E��åU���AjEİ@�m���E4D�U��y��S�Q9���*���F������Y�� bX�.K�Y���f+jn���#�a��tR�r��h,�Oz���T�����JbB�Fy)L�˘��h��GA]�����R8�,�%d��?Ee&P�u���{�q7>w�8�#��ȏt�z���mÚe�6
3ށۢ;�+�\��;��������:`�2��u����HM��֑���=k���=~�A�O�"O����yɼPķ|���L������-��pyי�t+�j��/�������xсS\�cl���5y^VO����s�@�Z�S؞&'�^�F��Gݿ^�*��윱su<	��T����]�<���.|,.����^9���)����l�y���q��d���%|�z-�s�L\?*�7����"<k��:�0�u ҖO K�}8�ߧ���زm��+��f�֏���Q�/J�~�g����=� ������C۱Q}�&��G*�d�e)#3jO��{ў�������^��>����S�=�����1���+>�e����Ѻ�և~��h�#�']��gO��ĸ��߆·qU�:9D������m��3���K��T&�R{����6/|{��p��xc�7J(�w ��vy�T+6V�9�k�`
��+�XÝ�{R����K"|36'�?P�t�һfus���Dm|҇̼�F['�iJ6�fXv� ����j9�	y�;=��At-�s�=��GQ9εyy�#m�&�g4���hoA7����x7���#�5�q�)���G�]ʼufTc�v��֭��Fn�F81���~�Z�}=���g����d�٘xh�T;��|pӠ<�ۏ��4F�,�3{�'��| �}�yd�E��g��ҫ���³�$�O�!�Pg�@�s�{'�=��CK�>��P9����W������o���+>���웮�0+?`�/R��^��w#�9����jc}ꮙC"�Q�n�<�����/����z�G�A�∊���+�{B_��[�>��H.�π�R,]swᑮ���{�bo��Æ}ޏS��,��ENnݙ��+/�fg6���b�G�<�Ӡ�X�)zdY�m�Dk������BEϼ�A�B��u��s���5�=��=�T4��T5�u
��F��>&&[�&�=+��9�D�D�J����y�N�RU�.���u9Ѥ��zH��z�iL�.��G���=D'a�C:	�~�>�g�Ϫ��q��n7��u�	��9}�@��\�{�:��g!K'�ٽ���N�	шAs�ɟ؎�i��~Oq�s��&z�}�_��y��mW��z|����P�����~I_��7ƿ3��?V��5��]�s=df޺}l��~E��Ԩ�T��lidۦ4'/c�ʕ����v��F\�)G�T���yO�ӷt+>i������ٻR��I�6�P2�䬎�^9�i�}��q�T��d�ۼ>
 tjwS{�^�ɚ�S���s�Y����X8�,em��/>�t��?uǳ�wtb����7��>��@71�>~�����������5��F}�}���գ��/�����w���]q�cפ���	�P(Y�ڝ�km��^�T'��
��zY>�0։�0�׺q[�
�<7���Vg��pUWda�y{�C���"���+�4'O�&�B�T���N�0�v�C3��=����}gّօ�F�oΉg��P�W�uU�s:�P��<�vGep��Ӓr԰t��2��0z5{ήu�����^��ʦ|jS%�'�:1�_��E�ɷs�{!y�%���}�9'F\�ƈq�x�����|��L��g�_���f.#��<珤����7	���Y��?�j�B��X�J|'cZ�E�c��֛��"tW���*���#u/�x޿U��}^_���1��>�`+g#j���S��WU��m1��ܥdI�OQ� R��ʟJ�����X��4F�my����_5��y������!���Ǹ�����B>$�a�	O��|z[.G�ͥ�hͱ7O��|6�KH��� [��V�D<޿�&�u��[�ݾъ�sJ�jw�Px�K�B�wECˎ:I��^�|k3u��5��G�:Yvb�TK��U�i����8�Qs`��ǌq����nVv���yHS�,�DL�EWR:]��K|��ӽ)EO���K�&�|��q{k̭�*#x�yIP�W�6T� ),�����Gceǭw��<��2�`�l�+v��n5�\M��֑�>��\v=��ޢ7�Y��2
/�w���L�͝���k]P���q�8�X�G8�֍F�'�l�g_�|Na=��h
+=���-�-��Zw(�\Q�Ko�I}>�S��#"mב���>=����+�����b�������گdqs��;�uj��}�Ϧd�#�z	��+VS���/M.t�_?\�ݏb��
�Ț�5���P�s�foޟ��z ��Ԃ�'�L>6}�M_q������a����n�d�P�r��=�+�c!{�to羠[��O�M
ו ��'�0>;�ݨPq5�ŧ�(�B��<�T̟R3��H��q��^��9�@z���bw��]
�NI��`�ͧ�a��/D�2g�����	���ï�o-���q<u���q�5�.N�Ox��;���՚w���S��V����\��!��ft�9:v�e���������>�J�T�l��� �t�~+լ�?D��Z�`~{\�,�Y�@^��hQz�7�)\p�m�kjZ��6���Q+�«r�I�:�(3��v!��,䜳�iL�{Vʫ�n'�jB���G@݃���̬)�,a�EN��uG�bx��wp�5��;'#Ou�&X��&���׏�H�£Z������W��O��5����Ҽ1�*N~w^@y��^G������я��0�!*�+LgM{��t��t�q�x�+;*t�d�q�xk�=LOL�N����qs9�bzr��]���;��F8�3���xyz�QueJ7Y'�I~4eT7���$1F�="��V��\��i�I�}}���������#}#��D{�����^���\d��,��i�w��Q��{n�[X�yh�Y\�z�,d>������O�{/H�|s�%��j�ni���|�W���}�3'6��]���}�3�~>�x��aF��G>��Bn}�H�g�q��{���EV����Sw�/�_�W����%���.��-��pyי�t+֭���۽,A��ۣ͌>uo����Q�9d�yE\�-0t�C��x�+Ҩ�+���C�g��2z3	��*k<b;��w���5lzQ>cӁ�9�K�rB�OW��^#�c#)���QtzX]>/'���ǯv1^�.���3�f|=��xdx׀�Z&���K'�%� G�LNΰ�F� )L�YJe�K��\2��<�k �/]v��s{����g� ��M̬w��*p�����Na�u����CWw�sP2u�t�Z5N�Ś�IK��=2'jo*ͳ�K�J��A������/��u�:��u`�P/&��X��#�����l���~���������{���H���@w�U�>ɓ�ލ�8�=Ys1Lw�L�K��>��C�l���]{�	�*�	O��m��ϓ��0��>��ۨ����d������f�>r}���p�,�P2|����g<po��"V}�Lz��G����������x�Uҗ�����r�׵�b�ʊ2�x��y���0�M���9��XM��cwuIu�y([>�Һ�>��9C�����B�J,Ξ&�L��>U���e�J�=�M�ye��y�>�i� ����FC�~����x{�;U������*���N4�#p>���N�\�2�'k��o�ޭ۹6�\�GO���W������z�=�ޮ�7�M�
]9'B�uo����䳑ڽ�+ę��P'��]T�XȵTY����ϣ���r7�<^�����g��{�Q��g�1��&�Tm{�=�6rg��A�3�&�,\W7~����W�V'���B����o;H��ں��`3"���T׌����e���)A��)zd-��S�ފ��	�^���yY�&�Օ�X��:���HGH��ڴd�}��6�]*`x���q�I޲Ԩ(❼m��!Q�V��Ө|�K�+<m�tJ׌�ɍ�4�nbXwXf��0:Tv'1�9�_;Oky,���d�Y�N]Y�mv��X8�R��N�Lo��q�
��Qk|���L���CO_��A�^�P��F���nx�=+���eW���Ʈ��K�����m_�}�ldes=��\8�������Q%K@�٨=$yǖN&'^x��Y����t}[>e���k7��j:���G�(�S`z�3P��������i12�*+9��X|vH����^g��s��q�f�o�������O�|}����r���WS�gE�\W*«��{3#�QR	��82}=ƆR�i�Ο�~�{Ϊ�'��h�ڑ�>��V6c
!tr�k�
�r�fI�"�Q�l	�.:�_	�+�������0L��>���*�{\�ż��ʇ�W�dN�G�
�yS�C'�f!;��W�t�H����-�>�o��u�A��{hb�W��}�^/cʬOܚء�n8��07���w��~hD�O��f!�䲉u��jy��[�ny_�:��9����uó���g�$�`�ؐ+�p!E��y��t{����{n����g#f}���~��Q^,��>g��F��}_���&��_xBi:��g�5�gW$%L=�RI�HL���w�h3djb;p��b��-�B}�
��`M�D����aɯ��<�U����V�o&*�T��x����G�%���9�X
��۝�1�H��IY�Z��\}��Q��w�Oeu;���t<�#�������t�}�c�>�[9�,C�����_V�9��x�FvT�rA�P�<X����&��K7��a��}^ ��e��ߐ��x����=n�� ��]�(ݖQ� R�EuR�M+�/]��z��5j�gy��bFouh�8�3��!���Ǹ���;�ĝL`px;��H��5���������̾ҽ��7^�\M�>w�9��י[�Do��H�2�߁��������\<�h�9y��+9����0o���}�F�{����"<oǴ����o�z�ڏM3>�S���1���z��l}
��$LK�p6:Z>��:јΈO�ٌ��:�㾙�7�^Uu����ǯr��W��ޙ
d�	�,DO�j�(\O*ZPA���#o��F������4�+S���U�'�"/IށA�(���'���*�g�O��sm��Y�:c����+�s5�����H���Wt.u�3p�>��;��z�AE����|G�c6����������bǫeדv��j�m���f��DHΦwd$��u�I����A�N�(�e�z7���p�Q�$����V���9�m�,�e�%>^2���n� R������6�┘I�Ǘ�.#W�N���+�ǋ�9��;�/E��Wr�j�aM�{���h��v��e1�ߪ���������6�hV���6Y>���� �/����20{ktI�~	\�]��)iv�߆B�W��ޠ=Jr=�Q=�ޜ����Ǎ�j�u�����>>�:�Ώ_�Y~GK�x�j��q�j��.k�\���{��G��N��
�w�N��[���Q���7�t���C��w5YgFU���X�/,�?_��	�⌕��n`���9�{��rw�o���N�G��ٖ2���w���t�i��ח�
�\�X}N�MFo��Z���ֽ�J��4�PMYJ,̞'�&Q@�S]U�/$dQ��:�^�������]؏di~�.1���~�s�]���"V>��i�$�'	~�s8b��(�Q�u웕M���}�JJϯ�pY���>�i��H�{��!�yׇd�pW�d����̿"k�s=��f��=`�>��L@j�]^�a�L���{�&��;���<^���_��r7����G}��R�R�{���Ӑ(>�Te�-ׁ���c"5�j9OԄ�O�i����3eެ�F����U(U��`q�Q�7 �}�>�Γ1�ILx�J�	��M��vW-��3a��3��U�ϕp��㩲����2�丢[I��ћ�M��V �3�}�&�R��2�X���SU�]��O�y6��Q�͝��f�6L�Y�Q^]Pr�S2*�F��*>�'�-��g�y�؀�B֩ ���"/��2���:�a5����"�'�t9r��:}!��x�D4o��-�u��W�V	�nOTX~�F����`{҉���˜�];�)O���C�3-t�o�)�͵����,M˺>���=Y��q�f�.=�WF��xdx׀��h~��o�,����m��@:$r���7��/n��/��{�L�������{����P��ޠ;���7�_�!SK}��⽹rԵKo��M�����uO������%>��YP�?]���^��S���ښ���#�_Y��0�H�Ǩ��'�~ળ�B�(�]�ǯ��G�OW���<�3{�MV�~�ս�=ʩx��׵�b������n��� �vy�R�4V�9������|w���t���A� 7��
S�QZo�w��a���Ԣ́����`u��C����+(����Ve����Շ�Tz%�;��C���/��x{�C�z&U{�,Gn׉���T�?1�)y��߰*u����_����o� }y̳�m���ti,���5n�kp�Yi(�>.��t��]��������q���Lق�*ж��)�TG�e>�:؃��8��%�z1�z"�[Y������8�}�8=	
�ZN-8".�f�~ytG"�jOQ�����}Y�^[D���\�r��z	"�߬:����
���<���
}�����&�t�p�'��[���:����)�N���h�Aqu���:��	��4���:�^u�9]M,ls�P��֭D�iqT:w����X:�.�v�i��䬺�}����գP�	�	���gC���=|Z�7�5I�4���#̹%������J�&v���CRly��+�6b�]�f�D;7	�Y�3�h�͙����h]O��
U',X�V�Sv]r��j+L=.[�6�.ұ�o��Ԃ�W�`C_q6v'x�3���C���$���� w|�N�:\"�J�;�,F���\Y0^��qٛ{��O1�-���7�k^b�&-A�[<@��5o�*�mQ�ݾ4t�ߛ�
��̆�]&��U�7�Qz�x7��CF�U����h7���8&��;c�9g�B�{GɵA��o����V�L�1���oA�	���v�	}X��8q�z��;2��ˮ��i7 v�P7z%�_�:�8��Ȍ��zh Jד2�����J��3!����k�,��{6uԠY[�o4�ojn� WV �o��W�B�}M,�F��!�P�v�oq�_��Mܶ��{V��t��o_|m�ՙQ���5fx���I)^Z.������X4o(��&�c�b��]L��};���U:=�����]	�����qE�*%急CWJe1V^�kSZu�a�q�ݴ�0���@�eA�*�ͮ|*}�%�u-R�\�)�f�GՈ��q��kt_0�;��J�}�eWM�Y�
o$r�7Z��i��`ɡW��nG/ml�C����j��5y�IҲ?���P�\_�[�>���r\?fR���iek��#u΂�ͪ���iJ��o	H&(P��$���W�64wei̘�YQe��8WA2&�e���ue����F,�	N	'L7
)�r���$�hVrk.3&hGӪ�F�V7X+��D�u�͝ʎ����\gw�0!��=v���{���;ؤ��%�/�D.���g2����:��;���.�l�E|V��ێn���Dmʜn�Т�����aq2��ȳ$����kD��Ůc*�ԡ.^f���>��ㄨ�$R����3zȥt�W�9ۧ[���H��ԣ�b�gVW)��r!�eAC���9�����4��bT��aQ�
�wh��Wܔ��K�)��[Cz����<F���Y��\�Zݼ���
��%��f7��6�9�����:��������AeJ7a4
/0�d���f�,�-�B1�B�V�Xin;V�F�;�s<�g�NDAͩ����14�E�#���i$��!�t�(:�L�4�6WU��br��<nЬai:�U�R�ILH����9!!̬���m[��xhA.�N�h&j���u,�T��'�e�D�Z�DE��ŉ����^"%t�r��-2̔�R�!�	T֥�E^녩��Ȍ�ktA���I
���$�,*�YR��8���,ۮx��YaZ^wf�5BEj�Y&��!Dt3Zs�D�{�Iy�#��%���Zi�Q�)�R'T��]�)LQN(�Tg�����=d�rĄ�P,���w12宂f���	J�2.�q�2�*	T���.9�r9ʓ	[���+6��G�ITKBUݮ�x!Я\�բ��Q�Fhr�+�=�)����T�!'���f�P �(��ES�nq�mv���z�FZ&ӤF�P���2uϓ��!�GS�*�j\��B%�AJc�G�@K�f��Hr��l���+���2lt��I޹p<�t��i�x��/�����z���}7\g��Z=���9^I��4t~��<�(<��z�o�^�>9�&������H�zs}>�HZu��k*=�C�)j��Jh�9�͢��Y�NH=FX�>E�����5�������~=]	�ʯ���*/����=��ﻤ��UC�m�QD�p���FX�)zd\���F���O	h��7'ut���W�H�J]z1=�2���=q�T5�u
��F��>&&%��iofP�tV���#�%J��+<F�{�+�}�L8��g���q7������ҙ*]�g5y�F�R�2����}�T��5�=/iѸ�J��o��k7Ѩ�O����|\A�S�ΰ
��2�k̎�>�m�����=d��A�zl�"f���Ϣ�y��������f�nW�7���}�������N�ց�뾛��x�Ϙ�L��>.ẖ�
pW�N���U�5�Ο���G���ż����v^]U<�י���F��{�r�+��+O���vHx�|�գ������G��se�~�]S���F�~U����{@v�4�5�����AԂ�Sf�7�l��c�H����焧�|����o9�q��GN؄�Q��5�iG�^h��u2q��ځ@�Mm�(�uʲh�{���#�"� ��JFME��Bs���K)��}sO-��)��1r��!�й��ϟz��VG��O\z�P��yS�C'�2a��;��U��=uh���@z;/E�n/^�_:�ǣ������K��M	ңrhW��R2�|G�?4{�=�k��ꏿJ#Ѧr�A�|N��^�+s����\���5>����\+=9'+��9o���B��{���9�Dܟ�C�-��4Ox�2*'�*1�ߤ�;���r+Ӭ�D/;�\���tL��h��}��t}�9'EڒΒ��<Euz�b��t<珤����O��{���m�
:�Z��9VS�+Ѷ�:g�q����H0��P�_�7������ռ�q>�759�[=���7cen[=����,3|b�eJ7e�x R�DWU)����gfK���w��EtT��%�$w��B���w#�D>���c�s��T;%GĕFa����&Wy+:�W�J�Iu����׽�s�~ӑ�^elyQ�ȑz�V�2��Ԋu^���֨�N������Ӓ�t��>�x���u�TJ�z�9Ӟ+���up7��-\q�W�����=A�P����J�M߽�s9�X��E�<� 59�G���AO� �gKV�] �����M#�ƪ�qŨ����ok��n'-ꆰd�w�{��M�4��MT+1]ŏ!��.��S��,XY����_(9|�t���9��T�k�K��N?���j���n��t�|7~��Q�֍F�~��dg_�Q����j=6�ʯ=Vs���wV�No�E|�Jsf���2&�yI������b�g]���~��7^���myQ�Do5e�����c���S&�d�	�^���1_e>�P�G��5���"��en����v.�-@�����!�~Wt<��̿�}� g�C��c��Dvc�AnW�կ�G25#��&j}h��S=Y�~/������� ���'O,����O�n���<��]rod�G�z=�4�s��R��;	O��v�߆}�^G!��R��eD�ǲ�)GI>��`�ht��s���^���_��~��O��Q�N����q���K���{���F<���ўarӮ%�?Vi��~3��zN��������j�΁**6e���� ىޅ17��ǣջ�����}[Z�d6�9b���ʝ7�>'t/ ��z��A�@yՑ"6<j���r{�)��jU�����>�|oåk��6�(��}x��F1�w��.�A��9���CW�)���A��%���߀���k��P��/�S���]�� ����F���d�c�ܧ7���؍�8�9}���n��nGڲ1�W&s��[��L:}=��C�X7�\��i�E����k{Wi�e,�G\ŗ�B2ws�G�Fڠ�.�C�>��q�|���xyg���웮��E�t������eueo��:}r���5�U)��F�w!W���G���\>7�����ۑsr%N�ﯽ+[%�6pg�|��@_մ�a�L�Ͻ0}�~ҼG���%����O��ֳ4���.�珯�lk�P@�,|�����|r)����zЉ^�Q���M{f�,�yY����v�G)z��ꃕ�b��F�������I���8;�w�|��IWF�zJ�.�<}�l?�|����M}�G�!�<Lt�WQ��P�'u�tw��Y��uEdl�{=�#/z�gޤO���'��4�>!x�-zp{#�y���I
q��Tr+ҙ�Ϲ�?�3�W��y��>����:�.���[���y��j��d�����s�Z:6�3�s\�7��q�y�Qx|{ޠ;�{��r_�P��܅�m�ZW�z>�d���r��@s�_]{����>�i��{p�?L�~.yL��S�
%�хQX�K��ҏ�)y�8)�Xg�X���:�gҚ/���,٨F�b�;�����t#��#.\�C��D�J�����9v��)��p���WܢX��6�FR.��:�]-�3m=���8Ԓ�M�٦�����c�Z�ޙJJ�<�74���G|�r�P��1FZ��&:�NqU^�ѐ��%wKSޓ�W&���y �N�é���vxk�V���j������0����07ɞ.Ȩ3u�8k�w�~�3{���\�/P/�޿ 7�������Y�顺v΋�̄�'2��<%ߥ�S캿K�=+�ԯ(��w��ۿ5,7�| ���쑐�_�'#�P���ʸv<��9'z�����qkQ�J�W��A4� ���y���Lx�}��i�x������u��WTgF�(u�Q���:����+�{\��I�c�&a��W�PȾ�(�j�Xy���y�/�2�zF��d���ǘW�o��7ƾF�F��Q���X��^�K=MՉ�ӓ}g���3��lZ�IE��CP����%���y\>�3�Ê%D*�,	/L���ە��署gN�>9�|u�3�~����������{\�;����0�Tu��ơ�T%,��W��(�cF���e-^�|vu��1����>��|οN�'������t��^�`��y9�ש�UyGjh���_=�����/t�
��r��䢸��$��m�˴�e	�5¥���ѽ�E�
�S;o�� ���Z{����$�2�Rh�*�kWD��4
��޹�*�:f��v�I;A߀����ຊ���R�ѷ�Ê�9����Y#ӎ������&1�kF��?[g �x{� �)�~u�{���/���ɮ�[t>[~|g� p�3:��F}6��^E*l��_��|�F�*��O�>2���/�פ��hw#�K���m`�3"���)W�B+�=�X;�yS���Oz��k�U�|kg�:vuD��ox�����l���p�%Ot@ɇ�'�b�k��ej�x��o\���D��W5��P=#���1��븷���{>~���*5�H�����}qwL,{���X<��Q����ܽfO�g�\�5������߂s>�z�G��N���4+��{,���\o�(.V�;�6�p�>��L*�� ���Ӛ���s��2U{����yK���6�6�B??{��E�֦(�95(�t�ls�7 Du@��3f����p6#��d:���r�:�C�p˸�~0,*���a��r�*��O�O��H	�
z}F6:�9ȍ�P����=^��7��U�i�U�ۖ�d;��YƟ�1�,�m��C�t��������2���ɿF	�_��v���Y7=ԝ�����ۻ�N'���)���7�y��,/;�m��R�#;z�)��xq�Q�_J5�vZ<�������gJԺ��CF5�B1�:�`�F�rn̔ݔ3m]���@w
4��s�F)��B��Q%�E�G/��}�*�"�ǩ��z��Sރ5�*;r���ez�Ǆ�|�����r�N�"��A�|���������}^yb.>��^��D{��{~����� �2�x����9co}jwV=�cѰ<k+�ץ���A�_W��q>w�9�����IJ��1̰�fw��e�,�G{kd�� ɨ��&t��+ŭu�����n'޴�A����N���x��}��{7|��C�9��L��G��0}$�A���|7C�F�Z��O�يܰ�? +vٍׅRw'7=0����>��6�������P�t��s�4.+�/߃�=li�^O ũT��Up��Qgޙ�K��F��9r�L�x���<e���>G�Ƃ���*3=
�c���,�t�Z�Ha����7^&��|{�a��A�R���|y����3s�f��öV�<�Es���Z}�>�����_j�������������憻��^g{(�lz��K��{��.#Lx��0�q�>�)����~�"�����{��{��a�5��@˟i�hk�(��M �MA�"�&=�C,,��^d�A��V��mT"ΔW����\gir�E�cO(p�v�k��dgJ��স�:�QA�n�́�4
`Ğ|Q���Τ�o]�����,{]_�}���}�j��6�rwMF�53u��M�t���X���*��.K�x�j��q��<Y�ic�{���}���g����͉��&���6x��F��?Tӡ�D�e�T�'��5�
Y9��<�MU���j3g� ��vϜ��9^�����^�da�n����?��n~w
��P�ofO�w��C?,�����z��M���}㮧��o$@��fO�`m�N<xmu���뒩5��D�R����>��{�B���~�s�]���7\+��RB���Ub�KV/Zk��h�$���� ꮕ]4��S�n��W���G�܈�\>7�:��a��gӆ&�:+��ld
&����$�	�{�u���ϟ]O��{�����r�x�>Y�P-�)��9ї5�~uy�eyo�6�Ӟ.�( yT`#�oᲑCUNx�~�&���EG��7�ppYO!ۋ�א����>��z�ꃞ�dV�(p.����{�����"d�ɪ��w�}�+���Z�8dO�팃����E�>�M��#\�>��w'�$SU`!u��#:��k��4u����X�;b���7����*jʊ^l���o���u����+��XM[R�i�;���NQ�K��6����c@~����3��g�Юو#��j�j��j��X2��:EN�K"�:�!��=b95�ǝ���^u�l�M2>��l���x�o��<��0_/z��>�"}�=8>B�rGJ'��q+2ez�N��N�{�y���;1ez�Gb��m\j�^7�3QP�W�����}��F��k��&��MKL�[+�E�%
�����>�>��ѵ+�h�|o�����W�����y��L��&�I���0�:߶�T2�dҘg�r��Nq�^��"+���i�w���u�<\�^䅖WwJ8�#��Q^���Pz��~�j��De ��!%�z<�+w/�ǲ^�D�>Z��Z���Wp��W�ߟ����*�={X"W���Ɩ#*~ڼ�*m\���x���c���
Շ�k�����<��z�7լ��wb�T�-��dU���W�LBC���lu��Gi�P��UǍKyk�
��쑎���s�P����+��#������˴�%7?M��Ȼ `�Nz�ܛ�nz�a`r���)�u0����P `y�{�����C��t��c��~�Ζ��.�\s�&;���
�,���z�]KB��	@7�5[�Q�mfL��V*�;Ͷ��J&08�/]�C���r��!t�%ĉ茥2�I���m-n�e���S�.��Y�g������ >�:t�oA]�u:�k��-��ŴejQ��}z�wqđr������߄�:�h5�#`�P��z��A�,\W*��tYO�/�����w|{'Z5�����hp���=����T-ф�\�jʣ�,	/L�\h9'c����#�JC�S�WPϽ\$tO��FB�י[�z�0,�:Up.O�D@���m�v�:nz���Ü֏�G��d�gؾ�Q��P�>�2���k�p�n=�#+�P{0J�=��f�碛}�eN�<�$��=-k��h�u�~��Ox�e0n��f(ǜb�g.������4�&��o�D�M���\�l��W��|�F�*�N��9y��u����f{*�#���l����,u�L9�3"�E�N�U��b���2�o��^UO?C*onG��<c�{��vM]o����_ɯYFG���9[���0N���v�#>����5F����x,�^|�ln's��o���Gz�C߮���������OzlHϵ�H������ճ}zPW�Q��c!��d��EV�ӎ�Y�ǅ��{~�W�}����:n=�Az�E������m�fd�
��D��� ��6�E�#�]�Q)b��P\��W��� �-�K�M�^�n�V�3�P������u�
�C �&X������ȵs]��IGqly�?,Ԣ��9u�R̛jřm�arX��7-�-��I�p�J^J�3�T�� N���37,]��\㳻������FҔI�y���!V��͛��\^���V�,�Rfuo}i�[-u���ḯc��y��aqPw�6�;�Ff��ϥ�~�*�h�Z���.�P�R�9��/~�s�[v8��B�0�LvWh �v�G��7��kf���w&�Z�X�)b*��r�͡Y����ӳ-]l��2��\�ʹ����{\[X��:)�_]�{��Ob��j�oc��m@��q��9H�`��t�p���s�i�Yw�#�AV�0�[�j�,�}m�D"�]r������}Af7��G�I�A�����1���L�8p��W�)⽀�<��;�z�(@�����oi�m��br�O�����j�J�GX�\Y�#�]:���X�u+�jaUz�de�+�v|i�jo;�z�9 �ЇJ8�k.ѥ�-)�D���] pҵrٸ \r�5F�,6-5�Ӵ���u%mB ���Y��U6m�v۽��^p��{{���5xq�f��%3���ً^��9ʵ<��6�eN�`C����-xI�Joy�{_a�vj5�{+!���SW:���
�hZhGÓ'����!p�g�4��j�	�]��wT���P�ez��R�ȱv��mǍ/YB�w��99��>ŇF�o^>���`�R���ސ�3�{ �/�S���akK"��f�� Նk"�@�����i��7ZΈC@]�=](]�����N��8�J���X&�ЋNn��%��0hh2�::��J�W�;u42,�\��O�T��V��7"�d���)J\��b����'x� �	���N��J�;��l0�[o"�CQ�Nj=sU�+�C�e^�����Ȋ#(���2�7e�lvѮ��h��ZA0��̄_��3�;��(�_غ�Ć��fܝ�ԅv�J�N����͐ڶM�Qs�9�m�nc��!Y�,��vh��t��:e���g��\���'�b��BvP'b��_XP�u%��lqb�u[����\^[��RzP�Y{Z�=��s���Dpm���"�&1��v�9��bf_."@����|��F��d��n�:�	���ml�tn�}�	ͱ|$ÑZ��ne%Yr��8���t���dq�[-��i3çS����[j5�P��]�ffV�P����ؠ�V(j�Q��hoEnI��E:�N]��V'�'�ܭc���Wp�t�Z��'��{��֚=sr�>@'�޶ʖ�7�=�}�Q��y|l̺"`�8�bQ��]]�{YG�M�L�t�<���_�R��iu �U�q�|�ͼq���=*-���-EsJwSӚ�#��Xd�BfZ�d��+Y�UΓ���9��Jyܽ$��E)CBwJp�Y�.y�n����k�\]ܯ*W\�$�W"�"tȮܴ%Z�Ĉ�j�)�r�'wKBI''v�j�z s�W�ܻ���#,�n��rD���;��a���Rr�q#̹I���43	B����VfJ��-���a�IB�9�������ă�uΕ8{�*(�M�]�Dz���8EE:"�HD�APQY�W:�4]�<��Ψ⊲���stY�y�wU=7(�����2�]�EF��bb%F��;���r9z������u���NZr,�1�uu��͋��F�EU�G"��GizlH��[�P�EkI�Wu��'B���ȏ �rp�\�]���r�� "J��̑w'rj�h���!%-�S/r��:��˛k,�%�ej���9*S�srL좞�.�ё\���0��B+ O5�#L�Or�a���޷�'�����Q9���5+�Ӛ����+��U^�2�1�R���6����{��zI����:��N�?�lT��sf叨�@�S8h��Q�\�~WᎥ������ϔ�R�UG��=�V����>�6N
��'�Ib�L�W��1qN���l��n�30||'s���U�����נ�;i�ឹ��c�u&W�q�Y1�7d��W��T>
%�I�ޠn������I��n�{>�����q�cr=����L{x�i�ۙ�I�N&0<�x.�	ܫ>Q��{Do'��S���P]�yb/��z2#}�w"=�C�z���raP�<m?Y�kG����������W��@K������Ͻ���~ӟB����IJ�2�V]��w>�%��o�W�g�&a�)�r�R�W�Q��Q��Q*'޴�A��㞨��@�:c����9�㠽��#i�35
dk�	>�&R������u�j�q3 1�X��w�]�^�IE������Y9��<�6��2)L��S��y��z���?)���,�x�A�
��0��*�
���}��z2���y"�w�F�Lf ӣ�)�ۊ]�]���^d4���������GO�k��Nr�����Q�
���t�����"�G�#�*�
YhZ|�˖D�=S�W�,Q鶱Yx���{��:�������^W�������OP�9r�CO����x�"l�r�j�eR;R֞�u�����ܭ3q��w��#���Wt.<�x��~���w�	����{E��r|uԟh|��ј|v�+��}�c�S=]�;���3��WF���t�^Q�.*{'Vk��zuW��zA�N���p{���U=��2�Gȴ��o�������8���K�I�����	qZ��Yu#��7Y>�9(z�·uY~
��<s�R�n;m\{��.���t���'�vW�({������xT|��g�#���~������>4��=�W~�szs�J|4�}�os� R�0|���W���UdW�"͌<Mܘϰ�yB7Ъ���U�'ɵC��Ҡ�4�F?W����T��]O�����;P�|O�X�zՊ���?L��\-M�����Lz'Μ�� y����C�>��x���C�xyg���쉺�3�7�O���h?�#�gc��!��R3ŕu����)��F�w�{N}�/r7���Xó=�nX���e�NLj!�VM� �d[=�����Z�YRd1>�4ھwê��zXZ�kT���`u�DOȓ�GU��iS�3^�YY#��r�s�k,��'R� gʺ�)��28]�ɂ�Xr���}�F[Ա�{�_)��"�n%�9�����J����� ��l�Q
X$�D�G�0.��>�����7�w�&������C��ʑ}[=��{���t�zޫ��gw�6
4���FX��-�1T珬H��3���M�;�̯`��Z0y=��v;�4�ǽPr��S0��rQ�p@J����!T�^�B^b>��,Ғ��;�C��޴8y�״���������W�&�����=��>ӛ��zp��[���d�.�����s������O����|�zp2n<� ��n�~���
��y�
S�[I��s� �Zo⤉��G)O��Ϲ�?���F�ͫ���R��^ o�Jr]J���Y>զ��1�S�f���+�3/���Q���Vԯ����|����������n5i���3[��h�){���Wdɯ�L2����=8��;���Yo? �9����xa���jᇹe�8�.wh�|��^��=�Bz�YF��Q�2,�>Gm�ڷ���z��q�`�����7P��y�^�_��Hz��G�Bu���R�{�V'�k
^ʜ7Y;��^��d��u� �'_�N,28��7�ݯc|4�u�7+tWw)��vp<2��W8�k^Q{T9�Y@S}'؊���;�U6j��:y] �۩&����֬��-��".{zȅ@����͒�N�K�e\7�����v��ݐ"����cB��h�Kd��零�8i����
�s��2z��~���uc����ʑ�<�X�8
��̱�q=�	z�zI���!za�ʭ"K�)ƚ���{$g����r=u�W���A9|��T'���Q^��6rN��r�cne�3�
�w&�\3�����}^&�9~>��=�v���l�-BSPk��o�<'�a����^�����`��(z��=3���/_�����i��&
S}Cױ�F� wdi�>�����[��\w�{�qnH=_`O��'��b�f��ly�A�E�-EO�>�J�Oy׆���1��,�Ǽ�=�ߌ>%GĔ ��-ӧ���͛H��Q�u2='Z��]A�׽�$\���g��^eoz�����p�:u
�\�fj�/g��~���"Zɫۜ��x��@�� r������1��&�}�dey�~�M��F����ފ㷰+�纽�}�̟J�f����끿�KG۬�j7Ѩ����p�s��m5)�p�;�<t_NJ�����wVP��e:j[7��"bm�м�T������5�=5�J|����Fl��6� �����WӱV�Ӫ��7�vYcCgVj�G��>�����/���ά�С������Ձ�.i���d8y�p@ozv��Zt�T󂠢�+������gm��*�tcVI�2��}y�;�V�ZS����r��b���j	�1��)HmyQ���K8};�}��	��9�3Ӱfaz�*�_e:�n�b�>p����ӷ��{_(�ul�^��wF���O���u�OO��4�'�d���0�psM���D�(��qv�3S^C�ʟ�Q��C߮�=�S�!��O_ʰP���H5��'���uM��T��|��f��+��r��ԯÅ��{~�W�}��~��<o�4N��-F�|��C׀��l=>�n����Q�M���;����uU�s:�P���� ����L*�ˎ�%�^��nrN\t�t헄x�fn����^%%�����;ɝ�"b�=��Ю�#�����y�Q��V�����߉Ú��:	A�N?�`�/�y��5���g��=��%�<�^�;GN��^���r=u��v�;��#�vT�����aO��uOE����CO�O�� ��.�<�O���q�c�^�^�C܌����R��d�м+�M�d>�;�IZ��A��3��}3Ҧ��)]\<���>g}�C��[㓓�6%����/@��'v53Ľ�]��������d��Yk]�*�n
�JS�x�����0����bc���ݹ�ҞީIb����y �yK|��c,J=]��{�rC��z�����=a�D�-+x̹��G&��:4�w(*�[u�ovdܑ@�q�"Tا���Y�N�us��]ǯ��B��D\O��NB�9�u��=W��y��{��f�^������������@�-ׁ��Ke溱�����&�޴��uI=��8�3��U���{�þ~�2���3P�AF�}�"b[��t�6�Y��۪譄��0N�����`~�N�0=}M����~u�2%zT�n�u2W�Ь���}s�h,���r��(/F�\�����1��V|p�q��=Q���d�� B�t[�3s]6Ye4����ew[��S٥�_y܏����7^'��>���/�R����κ�+��{	�@2;M�YQY]��w�S=]�J����]{�տ_�]������݌v,��z��̂�%{�~`�Y�k�[U�=�&~`�EX���1�V9�>���u�6��7��z�]�����PrXV6t;���U-�wK��Gvi����^�����)͟G{�S]��_����UD��Y�����|vv�g��i��j�Ί�P����wC��h�T��w�k}[��\g�үt"!��/��.�z�'X�^�%je_ymJ��E�!�ӈ�ԩ{:�� ���-[c7�zd3���)���gڻ�L��/c7mw'	4����ZgS�D6�K�;�η�L�c2"$�8�����]V+���<�w���X�k< �t�>s@/+��){̊�0
�(�:x��c��&#��-��.w��<�:���{W�i���^��!��x�x�C�C���'�FvT�^�(�;�u�q�M_I7@�Y�Tu�;�7�����#O�d\F9~���+��>��������oѹ7k�+�{^T����Ğ$?�2��I}��f�[������9��G���_�*��~t�8��y���K<�7�Ա���R,x�@��Sg�>}u>3�M	��W �o�M�b�/�E�r>jB/�G�K=~�p�e�`���X����6:[,��_DȩqW�ғ�}ǎ�}��S�}�Z3����w�#O_��A���L¸%p@J�>�r�'�$n*�O-n��JwC�
�5����;c>>ζ;_�������z�P%�.��P�U\�T���~/�'	���N��u�E��u�5������(�8�zp2n<� ��efH�N�G��9Mm-���D�G28�R��ER��^s�~=�f1��Q����@�yǣ�]�]��{������X9�ڻ��c���
b�݄�C�\^�n%W��M�tuM�T���aIBV
y�%ڥ�N���7{�9W�ISnή&�=C��DڗDT�G~T�+�9����k�6�]:7�����W�i,r��	��8Ȗ:-�YQե�_���.��f�S�xQ�~!���Vԯ����|���;g�ը���gT���6��}�-F��P���خ>ɓJa�#�Ӂ�J㣢+��ɼ��W���O����Or��x7ޙ�;<#���I�$yR(Y�1F߉�D�j�և7�k�.G=��s��k�f�4xz:�2VwW���۽�yg���x��V'�6�P^��9Y;�S�c�,�U��,�!�Q�:=��1�5����p;���+s���u�O��+>��#�xŻ2���F�H�kQ�K�7Х��;!��*[w�K�/#Mx���!;��I���k�3׳��������{����\��Mx�t����ۮu{��\uˁ�s�PG�ďO����ｗꬮhgz��ۨl����Ь��:/�$�%`���,d,��h�<�G|7�d�9m�������m��bl�q���ӏ����q���#�e�$��,	�|�s����F�����7�'������s��p��z�܈�Qg��y�{��xñrQ�GĔ���G�eNX�/N7�4�Y��m=��ν�s�k3:�s�@	VI��:�uu}.w�b+�-�盋�7�i�)7}*e�j)������:c3��X��6��ʎ+��\+	�nR���̷3(��Nf���n�,�x��֩.Ms��q!�������[��߽�$_�>~����V�z�����p�:u�����*	<}��Gt _�:�n ���F�q���n}�a�W��~�JRr`Q3���n�<�mM�y~!�W�צK�X 6h�H��끿�KG���"�Z5i��/תZ��u�k*���}���mh7ՀS�fiH�Il��&&߭�-�����lF/)�<�u�=^���~�����ȟ�'��X��3"�zj ����U��2�w�z���"�:��1p0�ތ����{�f�����G��Wtb�^~�F��}��:�&:}fIA��&{z�W&���М�R��b�u^�Wz�����u�`A/UP��Pu+�����B��H3��q=[N�R7��S)%��Oxzau�������W>G�b���ᐝW�ϟz�)d{��7��>��wiP��_�Q^��ܩjQ;@����ڇsY~G Ծ'N��\vڿuU�s*���>�G����Dg���o��}�u�����䜾�f���o�Ъg�tи��^��y޹���Jsj����w���TbZ�	�ȧ
vմ[�=o|ک�k�&{��z�n@���]u�`�,X���e%S�6''��5z�Ö�rO�u\#`K�VS�;B��P돣��	fr���m�P(����j��E�oLp_�������Z�A�Mz��%r�pULy��N���{��*�8=s:5zNt���tt��o�:\���������ע�x����l�ץׁ�N�����׼{���X�VvT鸲��2�7�!��*ڷ���FL�������(�>\�������!c�S��{�g���Ϡ��]�(�F�8�)cOzF�󇬓>3MA��.+����YP]�M�x��z3��O�܏u�����q�b0�cG��}}�;�m63��ᯣ�ĕFc���2��X�A�Q^�\M��ߴ�/H��ɱk¢z�X�w�\��yU爴}������W����5.@��x-��hb*)�\L\�������w=
�����ǧ8�>�8u{�FTzi�D��8(*��[�>/ō�m��!���F���x���ϣ��8��ه������wI�:�����J��A��㤇Q�������S����O��h{o����\o����x0�������%�ި��Ԁ�?DWF���nM��{���m���9tn�[5�0�kW!�n�E|ҦKϙ����ǥ���cm�f�o���o��� rln0l�������6m��`�1���o�6m��`�1����`���L6ߌ6у`���`�1��C����0l���`���L6����cm�����������PVI��\�'̀��6` �����������F�SX���l�D����)kScV�T+ee4�Z2H��e)J��
�j��i��)B%UH��JT�V�l�#EE4o�vd�4Qj��5��c�d@��5S��Q7Np��d�V6k[E�T�Z�kft��M�fj�16�Q��5�ɵk�I�F�T�+mCSU��>�)][��-���ڡ���b�i�f��f3[M�2�ص�뺦m�Q[6ֳR3&�l�Ui���V��+V�R�efR6���ة���wr�{�����E/�  ./}#[}�n�L��<��4�{��$���=�sЭ��ww�N�L��d:=kCM��F�q�[nk��z��]�w��T��ݭ���gR$�U=wnʍH�l�٤uLk�  y�:�����z�T�Y�g��&�#˻E�l�����  �E��ۍ�@Q��:w    (w���Q�E4z4g���t 4E�p�z P���C�ľ�u�ꎦ1�l�VN�  ���Q��D��.��V��u��ª�[����Z5�`uڔ���{��VmQx7	٫Y�����(�c�/+�����^���^�[�n��R�o'��j&��ݲio� �}��B�_w��uW�i���:��T�S]VէNv�mtڷw\�׳�Q��{a��������7Z�;�L�����۵���zz���m���۸�b$�S*��  �[wYv��k}��K�m�ogG(z��*�yy�޶�k\���S�s;�n{��PU��Ƿ){ܥۑM���鉪�:��w�k��r����lt��yj�v�Q׽^�lAe��ie   �|>���������:���S ���oz�ns�ٽs{���+�kO5Y���Z��瑝y���H�5��v�smޞ{�Ѷ:����P����z���L��ef͚�ͶZ5�  ��U�ѻgzOG�F��zKz�m��e�oo]� �[;ԯh:��W{һ��wMv�ە垷��]��O=䳑J ��^į/j�x��Y��+�������ͨ��,�WfE9�>  ���Q��U�����4*�׫��[��r���.ݔm�����w�m�+�M׽�h<�WY5^�A�T=��/ww�T�6�ۊ�yU�f��n�ݔ�]v"{UB�6J�뉞��)�   �=oo� P뷛���ثB��էQ7vz󤤎�g�ʃ��n��m���ִ��۶=<zSӺ�k��\�m[ݹ�k;Z�m�]�,�z��{nƀ�!^
fZ�V���JJ���  ��J���u��E��E��ջ^]���zY=�=��w`���׍�[v/O\=P�t[lE��m�!T���^���u��s�
����==�y�;��� �? �*���� �S�0���   �==4�U"O�`E?�SM�ɐ�S�&�*�M  $�T�1T�# ɦ�������_���?Aݟ����~Ϸw�4�1�/d=W_��������<�_{�脐�$�Ԅ��$�H@$$?�	!I�D$�	'�!$ IH@$$<�x?w_��5���t'��\&�B�E�/j�ͫ82��;���t�T��(�4m��4��;�,a���)RyM�I�"�&]dt�l�
�dmP��&X�n,��#FY˫s�`�XK) 4t��Ę�$�"A�I0���������3��gv���䲦Xd$�.�d���٨{4fU�����^���h&�(�kg7Zm�EZ5T���)aL���&��Z����\��U��$ysG|F��֜���<y�&,���.䲲�8$qe�:��J�饥$�\'��i���-Ǚv(��*!{4cSv��V�2lɴ�M�j�9���u;Z�B����b�@�++�,�i�F���PSec [��/8&-Lh�GG�vǝ��܍>S:�Pz�C�v�㽺19��������㳇v6/r'X�B�T��\�/i^S�H��[�r��SJ��m]:��H����.Ѻ_^��DѠ�YA�c6��Vow�q�١+3R����T��F�d��
B\F���s�i�D�b��%��2��4���yK1�@U����մ�q[ ���ʁ�
y���[f�[�J���b��"��n�,p�R,�X�j*��ؼ���D����.�5��hP˚�csp� 62�Zq�gKUr�`�(+�� nVKɢ�֎�x�8i�sXD�Mv[�Q�e^-�oZK\���B�������6vS��k�e����יP�*�$�qL�M�Y1��@K��)��"A��acn�2j� #n
o�7h̸��r���N��S�MJ�V�h�Saͭ�yAM�hl �W�]9��
���aF:�Pi��
��:�if8�P�$.#�2�x��m���P<F�Ûo�3CMj��b�S5pU���M:�D*�y(9�Z�su�1����#xy[I�l�VU�n́���Fv/Ai�e=�Z�	`�+It�����-��,���ۢm��5��lV-reT1姛6� t Ô��`��0����i�w��h��U�k_d� ��-�,�f�t��Fn��eTzq\��e���M���Cn����O�dM٠�r���4��tRX۬B��	��MZ/v��#�������4ܩv�0TN�;�r�K�7��&K9�XM)a��Kb�n=V�	ou�-dGUe]�
���쁰^@�#A+��ĭ咕c6Vb2Z�W����8�Vc�i5a����R��`�t^S)��'�v��7lM�&��*M�CS0�=��35j0&��TX[
[R�!�iis%B�xٸ]ڳE9���*B�fL� y۸a�A��zxodSf�@��"�=-L7�[7K�"]nb*��liʖU�b�!t��b��J[�*�B��aX�Hֵ�-��J=������ݩu�V-`ECM#V�"��Jǘ���+������r<�b˛t���x*n��b�ӌ
IV-���B��-�⬴Jm���Y4C�!t��R�l���2�B�G��$I�J�Jm�휻�2ލz�+fЛ6�W�X�M!ܭV��1�9�MpW�1T��z�lC Y�N���������6�`8u� �siլ������R�N %Cm��,Z�Ql�����Z7[1��R�����o�R�%�)ȴũSXP�pJe���i2q�8(��l�B�?�@D=9���j���zy�'�x&����5�����Q��I�0�%:#Vnс쬋HVѕbb�IG�+����pϲ����R�H.�Â�52��X���Ɇd���WH�k��H�qڰ@��+0ұ>XJ�XeT�m���e�!�y��A�q�S^����;1i�,�pr�^XFi�ҩ��z(�&�Ҵ�KrĹD�а�u�n��b�GXڌY�v��[gX,f���32t��F65jة�h|�9�r�V�ie�,�.G�ٷGF��8	��V���2ڲ+l�J�U	����³\H�㧆9�odl-̱��7e��Dv6̟id��=z�
����̺MH�;V�\32���5}{2�u�t��Ӗn��C�N��)���X���DST��7Rv�ףq:YU��)Z�s�[;�Nm��>jܔn��-K�v�2ּ
��Ŝ{�E�R�R�{j�r�6,
̖��wu�`պÇ%�Jfbp[x�-���m��͂mW7/4S��e�3n�70�7m�ܚ�^M@�P�����b@j�ҽN+w�� �@�5��"�l�X�i{�:��x.b��+1�Yz��d0G���幾�O4��q�if��$�$:�i��h(�������h���0��:�E���XosF5{SX8�SwCH�M�5&��s���������7��%�f=��.w1ȋш�7/p6�W
�Eb�`/ņXjM�J�ƚ�����ȴì�cM�3aR���w��',�j���7�LT.���N���r���s4h-��.bܬ�Sf�e��hd�����:C�f3�@X{=��&�o�t1]�gD��-h�!�CjP���ҔC�2Ruw>�l�KF��n��ʩ����Af�捜�[NR؞�b�+>&(�
5d
�v�X��S(So۱X`�lp]��J�8r"���y&3Ym�{�ʽ4d����a�3B����FF�C2ġM��j�˻l�`��*��q��8�6[�c-4sA�ҫZ��J�m��1/�V��+sP{�%�����x�U4�3e]�Ȇ�h�F	i̔�4]^Qy��A�J�P]�wbH��k��˸��F�.�\C n��wEK�(F-[ځ��A�(���51�ۺ���IY<�sS'4=щw�͘��i�,��-s��OX�Y�F],bjw7ER�P�1J�!��¦���@U<��K7!Ÿ/5l������7h:��Z��^?�WY>��t�oEX�(�f8QĨ����*���kL/^�3�)4�.���Jȵi�Y�&�wD�H<Ka��h$����>J��M�t��dm�sq	��ܠ��nG��t�ck�l�F����:O ΊJ�K�(V�YZ�9����w7F'�S0���^ ��"[i]8�K@�f��&k��F�kq�0I4�*��=�sB�2[Gv��Ј�)������j��fM��u�13�fV:��%=D}��i9��F�to"sf�ow�J�M4�e/�Y�qʖ�)��l���&��ؒ�F�Ԃp
�+��cN��/r��X܎U�T�iف[.�a�VP�V�!ٷ@<%=�r[[���,����՜�ǯ�.X	�ߟ5��/E�(2���IcQ@`�ͫא!-I�i���I���`� ��nD���u�+�R�)�Q���/*YY0wBS�*�v��5ݜ�P�Ւ�e��sV����+�l1�)y�\-
�E��u
��Ō�v�ƀ$�Jol-)�5R�X���-#����Pj�Ȕ�נ�%��(0��Lpn N���Ej���⻗ G�i�,@����۔J��hơ��"+)�9��f�V��1oq����DLDm@e��H���ҭ�(��ƝI�`j�sr�	mSxV�ɺf2��mՊQ���p���saq��w6��nX�;[�Wv�T4�p�F�6dAA#��ǁ���#+��gپ��z�AY�|��b�K�`}y��Uw�c��f6k4�h]6�5lhݪ�-iF�TX�e�9Pn� �E�ʚ�6�ݠ6��T��s)ݍ�1h@��]��?e^Pf�$��hE"4	��ef��	{�#[�34�;�Jv��)�5f[P�]c�.�h�굡y�L8�:*�@��a+sP�z����&����֗j(-B�Ճ�oS�Fq�B��f\DH2֧/����x�5�Kh\Y�kv��mⷔ�lue�#�B�cK�ybi�%;ݕ(� QJ���M틉����[YJ�V;���ÿ7*9M��������7Ӛ�p�\zt�]8R�R�ì,�����2�\k)u�(M��
Փm/)7�[��ܱ ���ȅ0m=e�N�y���L�f�2��E�����ɶ����*����r�)tN�����1kYV��r����U�i��V��{I�8\4>�Z"�E1��^ӧVH@�g&�ʄ��*U�2| ���J�eEI����0�[�p��kg
/h��u���G�޷�F�h���v�e,���dC&ax��v�+cu2ʁ�q�D�Q��Qf(#�1e��c���EVսBC�`_�]mE	���%�����貲�bZY�Ud�ZZ!�JJ�Ra�*��QK�Y�-��Gn�����xOґ7t�+f(�5���ImAD��[2��iַ�:ҳ]=,a7�1|�<0��5��P�Q$�i{������i��R4��f��9�N�/hP"��
_aɉ���YX�VPJ]%�@)cR��k�F��YYF���s�YV�.�7�x�a+HӺ��3%н�[�U%D6ԧ�Ў7�e�R�I�n�A������2� E,�p�i�w�n�u��f��jEjCp�n@�Sܗ{7m��t����Ӧ�E@�q`�)���K[�ixn=� ���)�� �Fjlç1m^���xX����dv�Y�"�!_K�rֱ�b��f-��A*����դ�N�t���i��(K$m����b�Z%�\h�vڻ
4�e���n0Y+5��-��1E���*�]�QL5��aͶi�I�͚^é����M�9 ��Y	������i 83NR�PK�jb���"�'p%��1\z2�:�5���[EQ�9V��E�P��~gZB+%���$ζ��i��C*�m��c�.�H�N�-Mke�[���u��&���%���j���X�iAm�Z���75ڣR��O�L�rE������L@�X���J�4�Ӕ� �Ϙ�' �j�ĵ�E;(�'�-��hKX�+P�����̶��n�Ce�Lћ)�#2�,�j�Z��5>9�Tiji� ��HlL[��2�T�n�t1�֔�FJcn����,�W�Ά6,�Zoq�wS��=n��N^��M9���Ħ�0+�-㻄TvekpX��T�����-���b��]�a���%��jKMB��ae^��҂+t���݊BF��3v��+$���*�*� ص.]�Rӽ��2S4`����1D��U�.��wh�ҭ�Tb,���x��KMy{X�8-�X� �Y�ֆ�hح�r�B���c2�Zڻ2����S��&�m����N�6( *�d<R�G#۬&��qf���4e8�)#��`Vh��7������2mM� m]L������D2��bv�3e���.)���و�5[�$;Rds@�`
�
�C.%j�l;V5Zr�9�.���E�ԣ�zr��t+vu7'�Oؚ��^EhLF�l!�<����.��8H��݂ZƵ���Y���6-�,���(:8�iE�p�'�5��ɦ�2�r�9r(�2*xFY�w�aub�͆�،w"�$�uڼ�o3T0Qg06*j;n�����[��+�K���70�����U�6	 vʓm݁7kN��[�8�YxN�-���D��N�Ӎm�������J5����@Pgb���Jhn+��X0 Śks'����
�R���6��0/��oJuw�j�
����#f7�KJ��T� ��U�BDbVBT��cN���ԝd�d�6�l:Yh!�Y��ˤ�Z��ojnc�6�D��/fL��S�4�͐P�yF^��1jWV~2�|���b�q��'<�=���کS1$Y��R�����v�!͡2@�f�詵��V��uN�?�F�av�ҁ]���n��6�^T%d���� �y�LQX���(�$�����Q܆YۻD^w�&V6.�#-Z�]4ň�Xʵuv1�2��ڕeL8i�Qyu��
#U�5�\�a�i�Nӫ�6�Yk2��SE!�х����[�5VZ��X9@�ZP闬]!�]��Vm-4�@̺WU&̤6@�0�H��6��vvܦrսe�+rfAiE�-K�i��Z8�ݔhaO,@-�;`T0�Z�i�v��u0�V�@�Y2K�dj� ��J��α���:ԁ%���VTq����:ĕ��8qT��.����mfb�$j"�B»	�q,VZ�ۅ}wAaC'F��U8nK&�k�B��5�����0ӣ�w	��F��6���+�Ov�%�Օ�3u��Ԁ�ۧJ�3-���͉¡��/a��Ju�q'j�f��X�մFs0��:�l�͓���5��2�`�F��v�Y�,�\�^=4��so�����&濒��9z�&����i�Å����`�.��V�N�@�w.V=���4����,Ԏ����H1��Ɂ�X���}��NfY���[I�|�nr�4-H�0�F�!��2��/ %`��!�[��(����." +Tp#�ܭ�4b1�aq��n["�FSR�(*!扎��`s%jC>2�D�%�B{J9(��]=�\�5R��s[Ӎ�-�1��-���bJ�MюVH����6���)<���0e��{jd�/$�5we&�jĊ:�pl8�"-l-����{l7����{�q�ڄ��{E��Ld�w��PALА��Ĉ�:l���ݐ5�Z�X`B��X���A���:ɰ�fV�ذ�Z��/QŴ�k�n�k�,PP��f����=�l�K��5��$}|S��wՔ5�aȮ�Ft�Ҭ�8"��&��1ap�mN��v�c!W��eS��uv��=}�Nk�b�0�}�z�c�r�����-�p���Pi�^�C�p�Cc/������Ir�ݸou��Kt%w(�1j��[g��S잓Z�3*��j����G(�}CMyE�|@;�w`[ըM�V��C�5WS�Ɛ�a��wf��b�1G�;\���$�o�Q�'�#�Z���F�r'&A���{(^�ڼ��Y �i�;k:(�%��y�]2¥�yD:�$Z7��Y�4�x�����]^�i5�q&9J�azC�0�VU)>��J5Ct��V�0�Q�;���=��G��<���l�&p����"�DbI��w�ܹ3Zm��`*�[��Gm����hw,��WZ��ʾ R�v�Kub���F�����1�b���C�����VS$�α�^�X�T����n�[����I<��W�b@�-L\bPʌT��#gfw�ձ����/M6ƍO4���y(6y���C���b����VN��ξ��V;@ �v����G}w�膋��Dg��ꋛD-N৪gF!�@�zP<F�����ُjZ������]�2���li��_��m������+, &�i�u�^M�5�תS��6\t��;������6&��*=K�vZF�d��u�RJ� ��Ea�==P=u9c�N�*A'�g1����պ���Om��:�Qd�z����	ڵ-�G��f�X{'F���+Θ�N�oy�ƪa:z!IPX ;�u��rE7�n�v�}X�ǝ���B��F�`�4��,����[9G�j��o��w�����f�<[���rrw�8/�U�Z�w;|���qE�W$t`vw�<Ц]5���s;Jy[ѕi|[��e�⟯\2��4�'���"�蜹��T�n�۽\�dn�\�J��s�;��H�����e�œF�w}
wԽ�$�8{u�{0Px�k<*p7=G;y(�I�Pp��(�J}�7�����q�}-W���7D;�`5ˋLcns��q�ط�{]�a,�r�N|�a��ش��f�T(��V��U��{���шm�[��6��×}N��������N�Mh��UZ��;����yk��ͷβ��檛�U`��̚'l6�=#+[�x���Җޕ�@��P��V��H����ӗ��=�׬�qo�b�Un-�p����Q�^k��þ.��{=ו��ng�\5�:��}�l*�ה��t����SК]k4�1�d�
�p�jS׶�U�¢��;�6�n�����O����E�ͽ��-#����G�ve�-����S(�����r>������[�sW[2��8��K�@b[��;������|��Sz޳���v�L��SB+2P�Uhbl/�	ɛ�g
��c�����u���%k�E}�mM�C�N̛�3������/[��K�T𤞵�K�:*�s�7=�y���bv���R����)�VRüΠGP�z�!��wmke)�}sN��X�w6�ܵRt�5�3{�KPx��^�λŔ��S����t��+��7�:	�߯\�yN"5��7'I�c�)���E�f'qK�o)��ܵy[�+�b�u�ep���W�B�wx>�����i���9�A�	�S�!'Q9�95g��
3����f��% h:���0�W�� ���m���:�j�5g^�]�.�U�X�f�R�:��̉[ӷ�-	��'�:��]Ko[|��[v�{� Y�FAq���\R��o��onB�u數�@��ު��lެ�O;0=�:���ou�43�*}�k,@�TX�GX�[ �;�y)l	��ba#m�Q��r�y��78>G{��C�$,�3���p/:��n���V�����)���]��	y���̩��������TP�J�}n�8)L����b��yy��|OS*�>u��y!�������o.)չ7HoȦ��x��h�b(2����a�[�;��|��434�;B��%�jE��b�k�ڼ�}ٌ_>���u9gx���(��t5���}{�vnx���A㖶.���e�^Ҿ�N�lO	}�x������(=�~��֋F3�]Mf��w��/�T���D���ɩI��ݬ�uĖ\ݷ3-Mx7���	�4��}��i����qs.�u�7;x��&h�C�9������/ss�,�V�ڱ��vҢ���h��h:a����n}���)��v�Qܱ-���T�8]E��݂�{���. �S�M�.�5iq����F���[8��k��q�?�g8�=�j��6�?�9Xթ3���	ý��� ���ε2ˢ�dTQ�/�:/��8����GΗ�.s��i����b�&@�M������C���v{f�t�9`�p�'#]4
���0JX�W����WC�X�^������7��8S�Ov#ll������yq�)��Q/�פ�ٳٹ�p:�*7t�P�Λ��2��d�Z��|5�?�^��=�;X�H����M��'���7١��"I��6��!u��;�T�<�J�Z��չy2f�}�"{����6����w$���G��h��4fE��|���'�vݼa����^6rE�iev�9Z:�[��L�-� �6rZ3�j\/3k�ve%��$�]3I��L����,(Mx��-X���w��Sc*J��^�^,�>;\�����\�\`��3`�(,�Ckuggi8�i˓�s���u%�[h7.@�:Śj�ǈv��ϙ��}�8��"���S�١H${7p�K6�7�թ��[6-#��Nt�[b���j?��}�iŃiݳ<��VP��]tM�a��u���t����f���p���OU�w�V�Q#����9/;ݸ�R��+����`Y��4t�E����Ƕ�������͝-l��������9Ш)��Z0�&��w�gue���W�᛾��.�!�p�-��O`j��p�7�9��QI����5��7���И�;7��t8�� fM�C�ȳ���q��/��۱H�|�)��8�vx�n�g:A���9����ُh��m��cu���t���
���$���uU�H�2�6L�C-���ow}��Ӯ�'�Ŕ�V�:�Y��1��.Oh�1�*}�����l�݆�B��>׮�X��gQZ1����/7�+�q��Z{t=�ǧq:�|�r�X:�b%pQd���xCyP,���g���s�g����!j!���/ްE�g��V$�ն�˟ˮ{��{o!그S80�;��N�.������� ����kf��%�'bİ�#��R�'
�`,`zѨ�[�+�v��ګ@M*�،��=K.�B�7�j����J�A�>:
C3}��J��{}xk�[`Fs�vBf��o��1�a_TZt�u�q����Xi^�m�N�3�t�+F�Q���p���$!�:�5޺���Z�-�sowPMIx����v����>�l��($c���p��8/1v�n��Z\&'���H7�8�� 4;��i+���k6�[�4sf��.ڍG���fo���8.�]/���Av���!�n�C-��s����sX#�^�Q�×ڏ�b�����+}P4tM\�+9 -���Uf5_7�q1ox��w"	�����=뽡�ɲ��Z&̺E���-2^��^�2���n�q�Wa\�IN��ʳ{tT?@��0F�t���bK�>����!f;�}h���W�f�2��o�hv2���:�;
��S�+
�(x��+��B&��L�Q�m�W/��j		���$5g����e̽>Fy��D_�A���{d9U�N��k��y�]-�f��j.��J	��h�72,��d���DJ��z"�m�6���*!��V�<[;�;4Vˬ�5�;�m�)��d����{}��	k�C8qGǲH��ˁ�|���X~�6��LK�tgQ.3���ͽ"%N����عE\�J�ޑǃ�"��l�H�5���<�C�cK�Mq��e�]��.���PnM�3��D�=���@�W�e�)�6P��ۈ��8�-��8�)V����7>x�#ы���h�7lVZts{�t�T�� ��6x�]�'6Y���M�v�j������Y����z[�I�g��j�І�����vo�b�XÒC�5)C,�M�4�r��&��M���L�N:{����ue�,�\��H�hW������R�v-�� ����L��9�Kv�;*NY� �2_k�(-;�/_os�x%��B��p{�7�AB�rק2�tr�	{|):�I�ܾ���Y��a��Q�!�hՔ:{۞�.�vם�t4��� �awn_��� �Ո�:��y�Q9t�ѷ]sb����^�u������˻�@��:��^'Xtpx�:��\����9��}:ɰ�^ӏqѝ��J��<7V5�7+G����x����s�m<i��-^��4	����z��pU��l' ���AmG�9P� f.��|�hc���H�v8-(�k`!����wΫ�\⢫�7RD
�^��0���:k�nvo��Ca����J%'n���V];h�
v�}��.U`��b-|�v�<s�鶙�6C����%�9;㖕;�{2 �'Ng�����q��Fm���K]��� �6��&e�>��Ry8v[��i�\{�&mJx�)�X�ñ�^��]�;ݸ#��ٳ�\�t�ATk���X6��h������)�ԟ-��[B$y�D�޻�M.81.�K�K�b���Ȧ7t;�iNX ��{6�W���E��J����q*(�K�ʋE�B�n9Ԇ
5����9a��z�Е��&��>�WkVqw�.�O�G�v��^�]�9\��`C�.�=�b�8�p�wJ�7>4D�mc�m���J���k�KJ6N��^Z��|�3	Ҏ��7g�����'xm�δݼm�"�8��F":��.���\��iWDq�Xh'�A �����X_�\x�A�\Ȭ��M^՛�=�U��ڜ3��[ʵ:ޥ�X4�GtJqb�YdƔ���^�`
5�����D���`�gt��	��+�wGu�V��̷s�z��lr��#+��s0��{ �89>M�
��C�7 ��M,�t�xD� ᠻ擑�q�}�\/���m�FY����e�*�p{��g�V���%��)�)b�b��|s�g:��#�\Սc)Y��Pи�*l�d�\���d9du@&�G��V��h��K�$/Mn�9H����wU��n�ݙ�P#�SG�g�30��.u�����f�g��M��3V�ϼ/��S��F����c)=����Nw�q�n��=����W6�)}�w^������7gv�'Ź�Z�s��g�����x'w�w^�u���,�I�͋peX��j��oEi+�w{�׺��렃M \�װ�#�e�u�Ղ-�n����">6��v�Z&����i}�쾴� ��+�Bi`�8)&�q��#XE�7�P�C�݅#k7�L�
V��7w�L�U�,.N���W�Ć���H�99X�td��XKA�QYݸ��������aMg���}1}���)�!}��=�Ķ�����u����|7�E�QZ���Qq�������+w��I���//4�P|iT��]�`@@�L�u����=�K��[��Qh��o�Yˏ�<�Ƿh�]��7oU�;+�N1����	n�,1L�Aąʢ偝}ZbV~&�L��Uoc��AP�2�=���d�;|��ǯ��$F�ǱZl͝.�U��y��1�W�2���H�}�q���'މ>�\UvUe
�p����º�m�F[�f��Wΰ��-��ua[�;�ƗK�ژ�3�q<ܛ����Z�)��@��j��&g�̜�70��L}NS���ʈHl<�j7��ɜ�溅u7jp ]ܐ�3Vy����%	&X<y�V�I�Z���ߒ�M�����PU��H�@�/t�׼U�N���)bTh�W±�����.��V�W����2��Xuv��B�'%�R�P�N�]|Rӱ�ޝO��-�y'&n]����D�I�[ �W�1k=�J��w�GhPԡ+.��Qvb�g�̔��n��9���)9QW�h��勝ڽ5�5�ϻ��ˋaHM���`����0�֮]���'r�v`8�	��5�Ѽsے�30�G��l�v�:��M� lÎ�Υ�� T�0Is�mb���:�d=ٌ[45]�[��E$^
;P�h�Ҟ���o ���w�8\�ʱv���VZ����G��Q�,=�]#��*rt(�k���4d߸,;����_L� ��/��Ո�&��&�Eh}�3x<��d��GR�W:ɱ}f;m������<�9�v���
�_U�ѻu%e��U��T�\��>�y�8n�t�0����6WW�v����Éf&EwN��٘T1�!��k�)9���Vq
��ă�ﮫ��{Zj��e��Ǵ9����A�t8sIRu}����]��Q3�ʝ�w�yn������k��5��hS�}[��!p�3�f;ߒ�|�̃��T����L���΋��&1�4�)��=ժ�zmc�䨷V4藟":/�E؊��̹Qq���X�M�XCY޵VöI�f���;�I՗�s��;)rK��O3xPK���X�S�\��uh��u���~�H��n��nv�p��v^��[;{����5��H@$$?�B����y���ǃ�"�l�7���F-��[���%�,ȧf��G;ӈ޳D ����W�R�Ӵ���gn����⊦�6	'6N��-��
�+�,�|����o��8:�����.��sA�4-;�#mVH}H�3{��ƃ�û�r3��<�e�|S
���sh�[ʳX6�h����8�ILW��ƵR��a;���y����[����Bk��{���,p��e���`+�T���8!�{M;����a��NzWս��ѯHϖ����܄fu���X��c�}NP���u�Z$]��sM��D�f��o�f#����E��'kM�K6�|�ڙ��ۓ#NGhm<��qX"���z��4���|xIBK:^���ղ�;���������u�
��]��'6�+U񑝳+7^l��I�[M#80�8i]�C���1W�m����껱-W�9���T/�Hm�ڬ�alm,�;�Vb�wq�pȷx1�2Ǜ�s��r�u�������vE�9=����<��kZ�.V(���e3�g�#Ws(���q�7v��{q��2'���R̧t��M]~<̹)y�rfܕ����Q�/�\ȏ8}�2�Nâ� <�H���v:��Q�=��y�SAu�o)�7��<�@����V=�.��y�x3j���Oxf#��	Ge˓�2n��êY�/N��}�G��'S��G�.	���2sͅ-s�xV��WAVճ�m�ˡ]�7�6�7#ѯ^�M�Bƻ�9b��P��]�l��A��� x���p�x-��|�a�����ZŚ/�N@�J��F5���Kz�
�� 2�4-A[���ڃ&��5�V�f�	o_�*����v�k{\v3���38c\�pp��
�d�^�-�ܦ��|$أ���uނ�Z� _R��y���]D���yH��i�� 6Ā�m��B7����kⱌ�ӈOyζ�W�B�Bv`�d�P]g�@ཉ1�1�R&V�Б�M^b��٣F^�7!��:2�G-{|��v׷qk.R�mԬ���h侧�VM(�H�`�W8x�黉u'"K'�JBt=��wݭ'e�u=��r���.�nd	'}��R��)9�H��VnvR4@��~��Gz�7����f쨖�>��xOV@�X%>3)0Ĺ�W7;��+�b�bV�P��6�og�ucyy�r��Bț1�@g=Z�U�~�.eNXGi�u}cZ��/���k�g�b�	`�Н�,u��Ӆ�qf�&��3�N�n����ZA�K��o�V"�ɒ���]Ը;�*��ʗ���@�%���ٝ/N�!��хgL�b��L���`+��p!��Cyf��r�mm�vu�S�d�[�rF�����S	
Kj�oJ�5�-�e/Zڂ�,0�Ysg,�q��E��[1f�ivd2!q���:�U{�+���,��Sh4
����3���Y���%Y�ԬI�������B���2vG���Bn���ɮ����v"�����%=���6�eja�R{&Ereq����k�F���;Pۻɔ�m���{��/�e��~Oϰ��;��z�%Nױ
Vn�,���T�c�`>�o�cLJ<���dtMr·#6���q�$B��wh���z7m̹�yܓ^��p/��'j�1��-F�o$���q��Py�^����'E�"l3�����it
�Y.�5��X-v$�%
Z�ǄuX������X�
��	���2��+=�r4m��x���2�r"�^�e]�Z��/d��a��Mq��l��e:���;�T��9�:u��փ�g�6�.�nm�BZhW�p�ݥI��8f^�V�����6u���v��]S^�jL�WJ�T�U;���m�x���v�[�^��� ��:���誠�Ҡ��=�X�9���7���u�Czh���kv*e!�g�S��'i�=C��5��up���ǽF-�T��kg�/o�X�Z�j"���AA����}9�b�\�u*N�1>�W@2����.��	�)�tGWR9��	�;���u،�+��l�yv�Oi�����DS]�,��.�#2˄'I��LЪ�)�ޚv�]�G��h���4]FV$;�yp��%p^��:u_ [0�<{��;�n���]�`����fi]:��=�@ ��dY���;�-�N�Dƴ�v,n�؋R!\vEZ�j�tOvhB<�W�J�	sVS�� �k���k�妻��M$i�{�PC�ʰ�Gg��J��Z�]��1z�t�F̫Mw��}�w�=4�b�����;�%sȌ��Wq%��k��x,7٠R�������VgN�f��&����<'ޙ9ޭ�3���|1i�վ��0gr]�u�72�,�Oj�ƄCkK�������3_݄���nD]P�K콄�q�
��w%�#5��G2�@�Q�{)��f7CWv�x\Bb�OÒv�q�ؽ��甙��_y6Z�Sq�sI�o@2��������V��n��|��c4���	c}}�J����;�u�+k%��z	��:�Y$f˫����O6���
D�\��ᭅu�r��#X�כ���_ 7t�us�
л%+r�̾�<*�%��g�僡R�:���oi��G:w����05�X�gs�,p���^�S�L�c]1��;��44�=4e"��=��u��6��ͼH����jwF�Z���@����-�W+�d1$z͂>0�'D2���պ3���h���>b%x����j���=��:�]D�R;�t�:v�/:έC�&��͓�'��|�h�NV�e�("�G'�7�y2+.Z=�M��dT'Af�j�#�����V�ۣ�su�lX�@we�*�/EN�y�ڟ]��Ύąd\�;�)m8^�d2�vC�Wv�;���`+��Ҿf��kv�Y�ʧB���[��wS{��H��$�B3��zk��"p$�o{nκ{=3�������bޮ1�0�{Hw}}sʵ}�f�V:���h��W;�UV�șh��p�(���s6t�ciSV��5�n��+���{���f��y'��5RI�{H��μ�������k�H��򥔃X	RhZ�k��]�s1,�J�8�c;��,�+�7�0htzK���i�Mf	3R�h��X��EK�)��yuvÜ�v�<N�ӕ.�ɼr��CG���w�rn������O�7�s��X�5�Nm]<�>N�IoZ���+Eo;��E��%ݻn�`��׽�=q�X{2�aK�l��ۖ�˙!��o�BB�U W�Y�w���6=eeg	s�ؔ@,�W�9��mh��u�$�[J�B���4���!u-j(}�%����ԫ`�;`&�
F^v	Ғ���|��*&�@�Q=�Gok�����(�譵ndso�'�q�s<� ̫��3��ػ6�5n�"�����=
���
�n�"��b�4��	�'^�e.��v-�5�
t0����_{����w���,��ZrvT�8֗O�t~\���7��d��؞�p�!�,K�>PpL���z��[�3Y5i!÷��8��i�g��n����ٸ٬��6L�iQ'4�]"�C�0Ӈ)� �ӥ�+8��֠ǋ)��וr��!�t��:6�.��獦]ڶ��AS"��;��Ll��٬��
��k5��/l]n�P�0�o@w)gD�g3@y��I�����zT%J����X
��s��'oMW	��qudӖJ�7�i�O]&�R�Sژ*L;|=���z`�p!�@��s�r�J�Ʀ+�{O)���%�S�w�L��ܻI�Ά6;t?)N�xV۳Ɔ�w����Xs�zn�촒�k�h���9n�ݝX�:�:�直3�h�Ρ��9=�"�T�%J%*i��F�B��0V�9�	��kaj�h�c:�֮g[&��ozVWQ�t��%�����m'�vm0��m��1��'y�<�ү��s4It�໨�Jx{F-�;F�:~�s��@������m���%�ͭ��<-�.���=�J��f+d5��<T	��V�M][�'er��n�8(hv�ղ���b�{�/����ч2f���F�JW\uT��N�i�����N�!ap��2(�=�:�N�N��r�0j�YGNJ��u��U�Ⓩ����>��z���)�j�l�5�0�Թ�ld �v+-f�3*��� _�	Q�������zƏ^��&S�hm�������gb�ٚixs�]e�!U5�1�r�d�G�,+�\��37Q�[�2����Zq=@R��9d6��/���\�dN��0���M�P�tj������*�bN��CS�9���r��ⲕ�]Vmr�u8�ù��`Ҧ*-sT�&�����,�NR���7�s�<)n��J
��[Jo
��QLq�8�ηhh��������H����/R;�:� ��)���peb�.�`�[�֥b��orM�X�*M§Z��z�GM��1��+�(!��e��poз'����2���i��-cP�1���VDR��^!�\��D�ɇV���,�ʇ�k.�쮳ʸi)��2����6�6�Q��f��ќ�[=���+LR���+`ڧI�.+k&(���]��ʋ�=4^�.wz��/��ժ�Лu��i�O��4�Q�Dv��Md��Fq�\X$��4��.������G�>���w�j��N"ZN��M�k�KP�ڣ�]<������4Y������6�{p2>΢��m�-��Og�}�����v$*����JF��C97K5^�3���s�Ԡ�ȁ6(��ݭ�4�ٮ�g&$����o4yN��Y6��r�)2��j�p�r��|��W�v�x)ry3����viVI�=끭�>�$��}�LN����/�n�!��O�){�a^����d�y���Wzh�ǖX�����	�J�>RV��2��,
�,�JC1�`+���I���-h�bIyw�mr�7������ao�(Q�O{F����c\����"t�]���C'vL���x��{2��B(�LHv�	��[f���G��ɽ3��![�m�]���v��з 쭧�g'��K�����zII�/�b;d�e\	m��`�Û��1���7���՚Ʋ��3��0��0�I���ҡ�ZuN`�}�9ݙ�{�V���7m�>B�CxC��dc2_<�%��ZՇ6θ�ڰ�n
��F�ϥn\����ޛJ7��t7,6	KbI�{�#n�_B{d�H�$w�������o�-<V+��+�r�t�i7�G�(㱀l\��=�9��AFE�a�c������.c${6�FHL�.7;�^f^�Kg��4�Fi�Iv00�YΌwU����<�A��m%.�p�89�-j
S����7�>yl�6����EIچ�LOg�.>�vd�Dj  E��{�C\��"�on`і����������F1�{�b�d�:!�f��=�,���*B�7�C}�L�Q�-)`�n͖�q3�_\.AiS�����8nB�<a��� K��i�#�}��dW��e��'G�kha�I�wY|aX�xm�lٸ8�Du%��`��=��D�l���O7�$o�%���	ԩ'�@ܭ'^f��`���[.*z��%��,AL�f&�6�	Ô��:K�ou�Ȕ��AJ��p��
T�3In�إ�M�������;[�B���qGXQ�+i�pT�jf�lblk2�+�!��)i�Hp���ĭ߮�]�Xm�7ĽsJ�0<ᝤ��&����s���!�:�h�R�ح�����KF�8s/��&�|B�;jx�]^+�x����H��S����z�~�$�^K\��	�;�T�"��}�8���1x;�~��\���P{��|W8ɫv��u���i��m�+7r�v��}����GC�Î�.�ag����ں�h�B݊�R9�~�+]�}�+�uo<��v>��%"�Q8�WSU�x���-����Fm�	uTꆊ��=j-�]��
�}�:�+��C���j�w�V���뇵7⑝T0pXlbB�����aزr�E�];K�.����5�l^9WmC*�°+��LR��*L>%SՊ�˃��A��R����\&��地��9���œ����$�Nl�i�.��O$䛑�@w���S�ZQx�L��"�����V/gP��v��Z]�'0���IV(���%��i��5t��tm_f��A�Y9����J�����0���h�6�.�����
���tt٥���E�DFI���=Ӝ��{Vƹy�C����1�c�M�l\n�oG���
�5��Ϊ6�Dv����)d�x0!Ê�m���1Zޑ8��� �,�7V��=ˑ�g�n�H�򢩝�x�9s)��#Z�غ孒�����wM���8�Kp�I�K���󣾷$��ѫP)v�־�Kw�ܡS�^��WC�M X���ٺ2q{��8G�m�(i�5�1l�b�bږ��а.�Ǯ��G�O8i�_B��`�>�D3��Lg!S	`�)C"���;���-��r������V���e�r����j$(��{������[N4�Fkh�H�j��T�%շ�ֆ>����tk��_*}�O6� �q�4{E���{��"�yRB�w/f`��n��5�ā���ѣ�[�ym����WnT�H�y�<�܅[���pr�>���ש_`#��.�6��䫓��������������Dg�gg[�oo�9�@��s����@^5l���Gu{ۈ�B�jU����
�Y�* >0�fr�|���ݓBʰQ݄XB�k�ػ��|��F�<���]{�wM�R�9n5���Z�C/��	KxuK���]9��ts*`)���+G%q+���g�짭�[l��fm�0��4��j
6}���݊�D;��{�Ѵ����O�dq��� Ms�|8��d��9yS:��^�FI�p��2��9��M~Qx��wi���A0��2-8&�}�n�N-��'qӕ7���Ǯ�`�E�wt�;�+FeX�b�₾�,t�j=M�����&�oC\�y�tr���.��f
��������Z�]�GP�*١��5��<�1�G��}�F�+ֺG�kt�U�{�x����ݪ�{ybb�����|�%`p9��p��r�ث�ʶ+w�����V�:�6��{9.zf�%-|�i�SK����/utG�5�������4���Q4������|XJ�܅��=fi��1o3�Ws�����[i]k	NxLцu�:>��8��Z�l[9f�DՑ{�n۷P:wx"��T1H�m]iǁ,�Gf�dۋw.�[��|�i��vp�q��7v=[�JX;B��\:gD6��k�;s�(k���S����X1K]A�{��նc�w���~���{/��c5lF
)��EDU�Ŭ����)�J����H��TƋR�cZ�2�U�+��ԬDb�-�Q1�PD\d��PT[il�����(��7)m��ƪ԰�PQE��mU�em�QTQej�m�Ա.\-,EVbT�Z�UU�kUKE�DƬX啩R��*
����kDT�ID��TUE�"R��YDW���U
�l���*�ֹIr��1���20UPU"���55�ihۍr�H��F#
�
*����+Ȩ��ŁYPEUQ��Z"6�DIR�J���%Jʋ.P�E"
e�jXT�r8����A���[eq*E2�q�J0���m��-U��V�bfU%
�V�E���E��	Ym����QIYU+Z�F��%e+U�VQTcimZ�
�3�_Q�3!o&���RF���Ė�F..B�f�SqܝZ���D����!k�O�=�di��j�W��u*q ��s��t���4�<����<�!�PUΕk���� ���K�]�l�(��^�K�4,��X	�������_Ev�l�-p8"�T�B[�j�l_w�$�e���k�e��fL��7�x������.�$8 }� d��"C9������z�M]y�t��O�F+u](v�n8���ȟJdf�+ב�9�VX6$4����೶�S�e�n硫�^X���Ȇ����xf��S9�/"��<C�P�\<ఴr��M
#�m�;���L���R��=T ����A~�W�����x{6���
��SWӁ>�g3�.�u�}_G�d�+P�;�V��w
�M<?n����V��LL�޳��{.ב^[��+�h��/�Dtv_��$�#�5�ey�|W���á�p�����5(�ٺl�!�9���LցN�nU�%���e�2��>ߣ���	�}�^W��5fs{g;qOv����F#^:���`��J��
��3��	��}�����T_�!�- ��J���5��Jd71�E�}�o� :iW��`���{��,	�!�u2q
�������Wj��O�MH�����_by���m��[arh޸K���g8���Bom�:GU�]����@�;G^�q{͠�+Z��ךa�<!B�4�J"���	�j%a��Ql�a�\�qn2��˶qi��elf-y�N������(����x�Ih����-k�P�<}�ou��[)�[����=tL:dſk=D����ו�ԋ�\\Hg��y��h�������F߬cB)�5i�^�xs��5����@4Ht��0�P]L�r��X�Ox?��7@��S ~�G�Sk:��E��rL�7������>@����_�I�\:b�ș���z������]�M�Xoefi��������Fߒ�0m��\��L
�H�.*�)^]�k�o�ȷ�)5�#��+"~���/�ר��������c]8}g�,5�`�0�zi,��b�"��\����g�O�}(�@-ȹ
�5���݇�I�r����&�`u��2��-S:��e�;c6d�K���`Yf����tό��<�Ն	%��y�a\�7%c^K~�<�{.�Ǵ�zhT7�X�:�A�h���_�V���� �c��tZ�ѻ�w��z�s��,=���gl7��;��n��b]Wj�r����'KT�:N�^��'*ڜN��^�G�.�Jċ�NXxn|�5�@�P^Z�[m_X�}���@��{��"��~UךZ����ڳ�)�+���y^Bu�>Nx�`k�I�o�q�^�Xx=G�����׍�9��:��\�bU|��8,2��<%o��Bz��G�:�e$`���F���{s�Z��g:�n�'��*�,ʖ<�Pdh�l<z(0e��kHqv�:o_f�^U~)��}�gh��ŉ���	��c>�xaV2�`g
�:�Q`q���~~�Sd�^W���1	FvDZ��i;��Y����g����KG�=���^ V��ŨZ�G�=vJV�/�f38��]��<ň�h;�ʂZ��+��Eqr�xoA�7���k����1k5)�䏘Bb�=H���4#VX�ܰL4:¢<I�"�l��4�mkfoUUc���ƮR�{����*j�ۄn�LF��_5�D��Nl�j�R>&WV�
���6��j��׮R�y ��0|�m
,V��;w<��N��U�"�w�Sz@�F�m\=��ݓ_�as�L7�4M�h���A�{x�y�=�c��=�U�w�ek�rj� � ���YY��/��K�[�}QмH�݆�RE�[P>,-=P6_]���\��<���1}{�7�����5Q<�C�m4+�WՎ�A�N����F緝�kϩ|��o�O���ţlO�C���mj�oqu�i:�w�<;|�j�S���<&
��FD�Z*�K�v�/�n�Xn|�tw'��,��J���_L��=����Q���~V�S6�T$�^�+���g�>}�A#��܃c;��������V��]�p9D�ښ�<�>�7�M^�f��V�#�v�g>���VgvR�z��T�����f4M�2M����Oo�x������f��=8)�
��cBge�+µu�2�z׌ڗ�'���~#��h�`�2pk��ۣ��'��L�=�Z/>��,I��כ��f}iڂ���x���Y�Ţ�ɛ��G��e��ac*)��w*�AGI�7l�	H⫶V2�Ã_f@w�L��;������碧�۴H�c�i��|�v���{Y>�pU��%c���q� v1�C�[��4�l�An����Rc��L����K���D�Yy�"�Q}�&�R�SL�ET��t�Wgtʦ[*J}|+�G5��,.�`�]v��}�����C^��bj�2�n\T=t�<��[Ô��+V�M�.LZ���{��Ov�U�V�	t�0c��(�����	e��M�O!�n���~�^g���xwe�w��z��s�T�A�x^������=����B�'��V�zjp>e��w�))��>`#�y#�/��F�2��3vY2}6ǚ�T�mh�)�����N~�a���z����'�0t%�BH��3g��Y兙��Ȑ���Y���@��o�[e/o��^�y��W�dq��D��J"t �c�փ�s'��hv�Z��/�H]^��/5I�4{��盋^�#.P�^3;��D����PL�g��Ѩ%xߔ��|���k �|\Z��iŜ�d��Q��b`��<���Ө]�C���z���L�V��9`�0m謶��;˅�Wl��BZ�r(E,P�ZHuZ���n�'�-`H�V�B˵�}[ռ�<�wL{�hȬ��EV�8$4�A��~��BB�o^i�}����g�	��ڬR�j�nH���ȟJdgt�'�'��OZJ��ǩ��3��R���&K�e ��<i�<R�δ�g:�o�x?�{8�5'��\A�9�u���f�m�z���u������'�
�z|���^�U�8:)����gb�%Vm�k.1k���t���G��ل5L5�ȏ�sρ�q�!ݮ�95NtW�e��b�TΞ����h���e���	˩{���M��]Y��c���'�At�n��-ޭy�͹���{ȕ�P]��s���s#��j���;���V�z��%qpP.��� k���+l����G�nnv+�]�C�]:]�ũ���+����Ϸ/�����~2J�7�]�P�r�Ɍ^.��-�WAI�pXJ?z�L�y��o���aUվ[�Q`�ڸ��{-���a�t�7�ڥ�q����x�Oͻ�KW�{vo�DB�	��4Ϊ��/�����,��bu9C����)!�h�W�n����	��:��.}y~3e����b[Ju*Eט����D���0�g���a�����Μ�x���QJq�;��<{��\mz�D2/U-�[N��pw����i:�=7=�.��[�GD�y�ǋK1���,2/�f�g�0�������WE�!�K��'��G�^+f�;�0.˚�׍����6����%���@�\�P����`��^
�n�F�[7
g��J`��G��*z���s<pE��FI����\ˠ�W�-?v�NN�sv��{8��A�X��K�r	��mĺ-��и��Vg�2��"�"�<;"�������<{m����`%��C�R����7�}6N�9�HG��B�Ci��d-aQW-�y���[[J�ߪ�0�g��0g�G[]�+���,�t�7�7�YFpW�<��k���>�:V�o3O4껡��!ܡ�t]O}�������S� Q��x\]~�����l������VD`ߐ���`��E4n#�F8/W���eم�H�őجRfR�&pޫ/}J+�QX�{�}�y�=��hIO��B�y�k��tɗp�ij��H�*��J�����e�5;����s���;�C�3�)%��
Ė7���y-��k;����e&(j��b ��Ѥ时o.���~]R���[z爾�Be'<�y �'��w�)�ye:y�e��;O�Mۖ�+��Yh���&�6̇}ׁ����O=MG�"���*�u�o}X_�Vn[�6������U�k3�<�*�#8U0|�W���]�:=z_ɓۖ8n�J[�Yh��#�{E����sJ��Uz��U�ʂ��A�~E��'��r�W�oE��	O�R�>��� 9����i;�a/���\����9��,Ꙗ�yiY'm���*X���E�Cc9Ӂ}��u;>x�|p*�&���뷩`Z��F��Yhn�k���O�C�Cz��s�\�6)�s]k=�v�������r��ޱ�M<�U%<�o�����9!&f��C+&0%���K�Lb�}�׸���J3p�{��F�X�a�d�I�o|�!�RUk���욭Y�-����}r�a�=�f��}QO�y�q??T�^�y�e��x`.�S!Ĝ���;��D��W�����㛣�g��	��o�}�S��-]��;}���}�x�G�#��=�m�1�=��:�I={K�E���������Y/�q���N�O�4>��gc�c�ؽ����/۽}4r�ΗӜ����9���%T��;%��U��=�|�6[��x_��
��y ɛ��3�WEm{�*�e7��� j1�ϋR�������m�C�la��]��7O1(�x���I��%�s�%�ks�_:��S�[���y�q���0wBk\��X��5����#ʗ�l����l�������)��^��z^��P{��z��GЏF�d�t�M��{+_�5�C���e=��S=���5�xʻ]��OG����{W"s˷b�hO#���E�<{z}��hᾒ�ְ�;;��t��w�zҐL��2N')�����t�-兵�,���	��e�1�:W�cO��:iXVݰ9$2��li�6�mQY�@��,3Y�(@t�Ԡ��V#�m�_*z�������W���so�����7=�F=�������\I7�w�mu�\���'����9v�UR��F��Ǭ}���f�W����X�*�^!@�/��,s(��ço���s������%H��U�t}*��CV௯���G99�>/�٬N�o���<��Ƭɒ4�����_għ�jP��lek�76	@L�sA���bj��q�-��l���W9O�V���a6=��0���k�H�Z� �\I{ۭ�7i��s$Ҏ�D{�|�9׳��Τچh�]�����-�(I�$5]�f@:O_�c�ϦI��uS��!��s�C�{2���ʜ�Wfs������ْ�y����ے�Y%Pï���l�׾����&��j��pY���,k�8�~ʧ�ݟ:��*�g�K�m|%�t~b���%��[v����XCP#F�iy�PHsS9Nw 5;(\����h"����g{��0:���^������-m�8�,6������mɳ�j^��.��P۫�eX��gg:�RgI6rƋ��	Z���:��(r�:I\Y$Ũh']���7���J��;R�!�>V|痔|ö�	&G�Cn�@�%��x5y���<�oL�=��w]�L��Ϲ����?oI�]��;;�0&M^�u�������k��No��g�җ�*}7��Ջ��.�^��ڑ��n��l�lX�_�t���v�ϖl��Ͱ3�݉#�~�P7S+ϣ��ٻ*yc�Wϔ��nSQ���������t�kv���E��;B�]w����+ŞK{s��,ٕ��q���-����G)��{�N%s<��}
�܇�0��]/8S���,'/rt~�~�g�E�8vzȷǯ�Ʒ�Y��5�S�8ߘ�� �bC{���tKn����kx��2��>�$i��ÁX���S���g84$=O۴xy�]�n�[ٰ0�oy���A�b[�
φ�3�}>zzZ�]��(n:�c��<��b�6Kz���K��k�G�=\�5倽&��=�w�sD�"�D����2�����;�ZƵ��{���-8v�!������Cw5O��6����)�%tͪ$G��F˸�Ш��S�N-&��9���i�|P3���H���]��*���\$	�f�v�Ή[�/n������&_jX;z�z�;u��`���W��௅^�J�C����L���bK3�^�0�,��1"�w�0o�eA�S��o9n@s��KË����+D�̗���qMP��xD�0Z�����j�"�p�=��+*a�9��wd��K�]ו"7� 'MՁ=�1�ĩ�JT��R�^���4oXCT<�@.eX����+W�V
K�I�fA}ȳ5��y�m�̝=�W>��X�h�]XF��s2r��AI7��i��-���rs�]X<��5�ʆ�5�	��!fm��3�S��J��08�9K����:�R�A�G��o�.�|8�=�C��q�v����fN��l�T�����:�����[�e�d]���׿J6�J�M!CLrH��,�k2rt{1�9Sb�ma\p�]f��m��59bk�'K�".A�]+2�,�|-1t.��hr똁�{����9.� ���P�^]Es�XB�|�ƆTvKڻ��)c1�k�d�W�4c�fCխiW,WK�r�n�H2Rr}-�X:-�ې��� �"���=S�ه�DT.��]�GD�����3^����j�M���`�䣠$�o�V�'�
T%���Bse�Cټ����X?+�p�$d��#��G��W��.�X�\jd?N�'�'�
�=׮��1�)� �b���J\��@���򢾔z�ICmJCh;R�|��YcK�uh9�;���	�����=5D�!3F��W*u��"����q���f���"��R+s�Vc��:�	3�i�f�/GB�N�
)*ݽ|x���1m$[碒CYK>�f��V�b�*
�U��}X�A,=�N@���m%):#��5k/z$�㯡=�5�d�Ϣ#�ro;~ m�	1�����Ya=L�X�pT�C���C���rb�˧�P#�
"DN�����$d�e;���Y���UC�G;��V�u+�e��=�ne@��n�1���5�nX�l��1\���H^{R��P�G�
�H���iG�+N�s��s�sE5r)��<΀��ݛPw<���U1'=1��=+H�g�e��hи݋���;�X����2��^��M��/)�h����UzBgSeݧoX��䨫Lh�h���-�Ŧ�Tt]���s�@�2�\:8��F��G2�mKd&�N��f.H�+C,����AA��,��ɬ����l	W�O_�Y���U�Z����[ٞ��Mn��j[mK!U�eDX�*-�ed*4�k.Z����D�m�c1Ĭr�Z"�QB��-bɒ�K��PE���f\���!�TX��S����V#"�[im��*����F�6�X�e)h��-DKJ�0(��J�Qmkm�j\iqqəLV9G3#mf1.d�1�n32Ȣ�dn`V9��k\�\cb�m�B��[V�JR����`�h4�B��5
�1���k���F��F"Ȉ�Yqhұ��Eb�s(�ha�-2��[U�j�[QUR�fV�(�����P�TF\�2�n9Z6elZ���iDp�L��m����"��r�"届e��1Z�R�3(�f#�,��PT2�&)�[1�V��U�V3+V��EfL�-�Ts-�ʅI�̕U2���,�V�jڂ�*Q���[ls)����)RDE}���Ǿ׋]u}�N� �ٖ����5���\�͘�:��Jl%�*ԏE�-�G7����E����K���2b]�Y��'�[I�Ž��n?yJ}��v���NV�v'��N���I-b�՘W=�y3�����]��S��#$]iOjy86����<�P?nn׸Lz�zb��u6��<�%�NS��s:�w�<��y�-��Ւ�
5�Y��i����:g���U/7�L�E�w�����ewz�1#���:��(6x�s�项�<l���evn�Q�.�ڃ%�'���رƪn6S�����k{��G�W۝5��O^��׻cov�v�|w'�Bk��ĖŇ+�O]��U��u��j�J�n�O)��z���w�[>�&���3���8Ė�����K�5���mK���}��v���^����5咼����~s�T�h{�ݞ����_{}��WQ'����W��ҳV���}^�~�r5璕�(�/5�D�F���r O#��wf��A`�=�$�lsU�������Bnn݉��2m�g�Θ��o��Y`�mY��)g���r�ky�C�� 2�����g�����E�B�8��ud�e ?����@5�T���[�V��L���ѷ�9�k^~~Ck��jXY.�zh]G����4����^tX~~�k%r|���ӌ�S�S������ض���+�����<i푯'9,�U��0���:v��JS��c�����\��պ�^��;Vb1�7�$62	_G:a}��bu�m�>�tɝ��p�iUYu�I�ۨ�#�Η���T{�hvM�T�~��Wt���sޣ��&s�Yq�}<�'PPA����/u-������\;���@tVk�鋢��q��x�X�uc���^η��נ)����N�<=�tԕ9�:i��&t�ϟU|�:vB��'M�]�e�<פ�ݯ=n�`yH���?IW����>r_^	*���m�7��וnV8U��ڜ�;�"�F:�ϤU���a���>�n3�9�AW��CSj��k�%�4�v�.���/>�g���̬s=�	#V��~��dc���r��LE�z��]���3~�<L�,ej�̯D
��S�f�:��u�����ٳ�h�t���+�iGME�®��
�X�s8�y�k�ݮ �!�f��P��&$�n�r�����˦�O2��\r?W�[����6�ynk9�1�i��C]��C��.׾�%��ⶊ�Q{���?I���z���1bB�t�1\ȨF�}�T�{�^�`^Fϵ��ڕQG��~<�g�zz^Rr�k}��=�\��r2<�|%7�ٜ�j��J���ktq��x���3����ۼ��d�+=�O)1�3�y9Kc�o�ꦒ�/ktI�ws�e��6�U8ۺ���愴u��ݮ�Ӵ�E�/��35�����at>�4���)�mه�x�L������T�ks��=�_J�����n
Η�7�g:��י��םM���@�m���/����r�Nt��=���M�vǟ�ƺ��ޖ�7�Y�O��]R������7��&����{���V�y��Ǹ����{v~��g����K�;	s�^��6|����y�F��WiDQ�]yt�zS�ӳ-K�o>q�I���j�{e�t1�w�.��\�.�V�ۼ=4��cU�^��X���̛~�a�R9B����}�9hBS%��]��u��)���aA<���;��s��V�w�Jއ���O]=���������v`�>�%�4E��|�·����R����d�W�������~{\��ɒe��T���>0��ݖ�'&,���}qo��-G<e��7�ӏ���ے�Y��Rçdq8�VVQ�����r���7oN{#�j\�]s�SѿK���Z�=Z����L����^���r�L�1�1Kϯ_�(����Ip�Rz?Cn�����n��K��'J_3�:��v�޺w�a.�	�=����=Ϧ`���u��������{��8�-Pt�/O�Mt�vw��y;��ǴR��­qUi��iײ�Z��i�G8br���T���M�͝�T}�L�cm^Z�y����WNO�Y�W�O�/���O��>�Aa=C\��q*S���'|ʇ2x���Rb5퇭d�'gs����&������9�/݄��'��X|�q>f�����Bjy�>f�8��u�m�u��a'�uw�:�d�3�y�Y8�	��s�d�ԟ�$�}�������x͗�Jvc3,��K���d+��XE�4q��#���ީ֯�ͫ���ۍ���D�mݞR��F�����w��rq���Pw�
X*A�A�HRE�h�����-�����)_
�k�4�0���~�ܽ\�������Y�G�(�����C�m�I����Ԭ�k�Ru	�7��8�ɩ��M��N�g���'u̝M2OY�w�Y8��k�~|�����g����u�8�t�$甝����I�Y���u��t��'�f���?2u+8�m�O�P�$٭�d�&��0�N��*k��N$�}�\�s�g���s���4�߾�����|÷�m���6���Ì'�<'�d�I>tf�J��C�hz���CYd=O̜Me1�|�S_���	S����N�`w����L��������s��"��eNü���?�v��a�^�x��O'�2I�l���I�iY*O�Z��q�Oж�u��R�O��ky�y��k8�>������{��!��I���=J���@�'=�߻�
���ԛd�O9́׉<d��	�m���+$�=�쒤�!��m
���{��߶{��g5����݁�8��;0�N$�?\�u4�1�o��}d<���$�<=�d�$緯4ɦM�� ��Oi󔑑g�e|�}�{]\�~�3�����מ��fy�IPP�ݝB�x��@�'m��RM��}��q����~I����'�����d���{�x���=w	�i�l?=׏�c������W׳*����n�o���D?}�e O�}���{�%ABd��J�Ĭ���m'm�0��d�?O��u�>@�<y�+�N��)�Iǈp��d���?n�z���_���f���t�go�
?}�}� �'�C4ɶ,��x���`,��~�J��Ô�
ɴ���Rq���MO��|�zԝd�吮�~`���{��]oO{������w�L%g�;���2Nxr����=@�l*��>��C�O�5��IĚߙ%J�u�
ɷH��'r�C�N!?k�<^�󟵜�\���{�]º�{���$�`��Ю(`SJ"��(J����U��<�^�T]T��n#�C.�����
��sͥ=�o:oe�����r\6�܃T�\V}�n�kU	���c~���4m��Y�5����҃)]-��f���B��_:	}U�'���.w~,ܓL���Y
�'�ϾβJ����a�a1;�?$�
C��P�'�,����'���$�M��ud�}��d�b��]���T�hn���6{�}�����̟݇2<�'�̞0�OO��6�2u7��$�X~����J��u'R�Oq��6��O}=�O�'��ҧ품�2�����t[߾�#�@�M>2z��̓O��y����d5�|�d�'X{>� |�2u��i'�u�Ϲ�PY%O��a�M�d5��xÌ��_�3���Nۺb��*���x�Υ���q��5��'5=�.�|�Ĭ'ϩ?3�(q���MC��0�	�y�>M2u'R{��'�'P|�k�'�u���:�d�!���޹�|��������ጞ%d:s���'��=&��L=���c'<��Y?2q5��=I�Vq�z�=��Xq���fC�N �k�䛺���߮�� zt�X8�D�ʉ������&��Sl��x�O��9�����q���~I�����9�IY:��yI�Y?0�����Ԭ�$�*}�� $}�P?�����~W�T��͋u��1'�(;܂��N�f�y�8��h�a�i��.��&�Rm����XO�2f��d�7���u���dĜg�|<~��Ќ��h^̯��J���gL���m��P�$d�V�9�Xu��Y�;���Y��'Xn^d�$����$봚�N0�f�k$�>do�-��g��y�>>��m+'�?3�Hm̞���$�C��~���I��o!�N%`k�ad���$+!��N{I�M2y�`x��'�,�o�>��/[���s��[�+$�:w�IXx�~��0�6���ZC�8�ԩXM��{���I&:���Y9�yCL�d����u�P����;d�&����C�r�1��(�þ���#�C=�zu�B'�2�<;i�g�݇k���+���U����}��*s`'j�MXs����VP�/8F�G�CZ�3D�A���<�Ч	�)9��
�F@���B;3X\�Yw�﷩�����7MW��t��?"�����~�����M��*
ٴ*N ��ɴ�d�jad�I����f�N3���d��N!����������k�����w��:��2|�vs����2i'5d�u�I4�����ÚȲN!��J��Öm
�Ԭ���m�6�a8����̆�q����~�?��~��~����^�C׉<C�d�$��<��4��	���d��<�rN��6�OP�C>���~��IR��r�%d�VO����&��߹�o�N�����_v��~����:s��N2q����+�M!����I��y;�$�$睸~d�����O�Y��'���5���I�ް������f}�y��\����������i%d��fR|��'���>`m��������C�s/4�_}��JʇygXu�s}�~d�
CG{��q'�,�)���9�ה�Yt�?w}{�����e���$�'{����~�$Y6�����I���y��q����_�<d��́��'�<7��IYP�=�N�d�?�d�
C>���37�e������߳�|��T=d�T;�!��~�X~a8��Y.�������$�j~��$��<���8�|y�3��0�O~� |�d�����
��o���y��}ϵ���޸y���}����a�a�N�Bk���N2|���t�Xz��{���u�[�:�����O�Y?'�Xq�x�5��<I�^{�ɦN��O;�w����z��..��Ͼ��y�8�䞠��I�a�|è,'����:�������Ԝd��'=d����Ę��&�i=k'Y:������F
_C��x��<ӝg폵~�'�������1��'g��i�M��y=��:��/����I��a��$�����8��k���N�|���y�z�z�~d���ǔ����';��sO�o���=�u@b�P1P뱔�WV�B���<=4�v*1�עf)r�N�3�5���a�!}i]u[ӕw�݉cƉ�Mz�K0
���>L]�#�[�w,ga�z�]�����L/�n���9F���|���������\Hr=[Ӳ�u�|�[rp_�����'�2��'S��1d��|`m��,�<��8�ԩ���N0�L�M0�`�βo�	��É&�Rx~�$�$�ݙ�3[������lָJɌ�C����me��?2|�e�a6�O��!�����2u*CG��):�ԩ�;��a�3�u�$���I�>���b~?��o�z���fK����ޱ�����N~�x�:�3XJ����z���?�k,����ї'�u4~�!�����q���y�Ru����{ܐO�~?MC���	����鲜8��QĞ�6ò� ��N$�>�)&ݲw��d�3�~�+����Y8����>C�8�e�i8���C��I�݇�?#������X��~��o���~���z��n� T'N��;d�&�<;��l�$�ń�m�]���3�d�XM}M�Y8����>C��Mag�3���cG��T��ק��w�c3ՙ��a8���Cl���yy��I����d����p�Ğ2i�����:��'�l&��'�k	XN!̲T&�M�o�]�����~Wt~9u��\����l���I���ߘk$�k�`N�I�s�d�x����i��[�z�ě@�]�:�d����;d:��O�~� ���5w���Ř�fg�����	��ĕ'��?@�'7���q��z}�Z�l'��$+�N���ԓ�s����Ny;r~d��<�r}�T}¨�_�O�k�	���^s�<�IӚ�XM�����I6�%I�VO�Rq��N���=@�C���<~d�'z��4��Y��Xnw�4�����v&��)J�inOv����<b���r�|��n���~���8�F��*V���M�`T�I<q��̇Y8�k��z�'��a�(?~}T[<q���L��op�P��t�m~V`��a�(�z�R.��&Z^U8�m�2CO�w��.��Մ:�K�mgvOA��2����x���L��-�ua5�9�v��S�	q3�.�CZ٨j<S�]r7�7۸�Y�����Ty��U~��o}�f���?}�!��r�#�~Q�4���܅C��%a��I�'�k̓�4o̒�2Nh�	;�'������[�4�}J��������~M���9���2�����I<I�� m4��<��u��
����PY%N{N�q��w���O�P��!Ԟ�~�^��u�[�$��>`s�2��N��}~�v��w�s��������;�?$�����p<a�G���4ɶI��S�'P]�xI�CP��u��}N�q*g}��N$��0<d���g�1�h�����j�=�_}����{�m߼��d��Ĭ&�Y?'L����6�~��N�4o��N1@��Y&��'P_>�z�P�,�~d����a�N%Bw���}�'s��-�J{�W޽�f�x>cg�">���>������'Z��&�A�C�q�I�,�$�+?��ԝBk���N �k��C��J�>��N��g2u4�=gw�����^��]��{��7~��ޘ���	Ӽ�i&����M�N�L�IY:��n�֤����P���N����&�T�k� �Ml��N��k��N��*o~g���ew��E���0������t'���a��d��M�z}�8�|����8�|�f�J��AC�VN����?2q5��I�L��XJ��z�����{{��r�|��3��i�Ĭ��I�N���9�'X~�0봜@�op�d�'��L�m�&��$�	��f�J��������R~��u�������y��;':�Y��6�߄?}� Y���6�d����m��X����w�v�(M�X|��l�I�Xx�L��t�N3l���|����J���/��_�M������X�y��Y�� ����<d�(�6�i��m4�1�f�8���C����$�<=�d�$�=μd�L�� ��Oi�I��MߠY^�<1��=��y|����"wt�v�o���v�M��g6LuƯvD9��c�m�w#����E���8a^��q����3���o]:Ώ�|��ٳh���8?'c��]�l�2`o�����Y�Y\8f�XT/'e��D�}���	=�����ky���!XO�	��J���!Y8����6��6�aI6���}�Cv�8�{C��}I�3�0��C�~��OXM�u�'�6�����n�~�^�h����������>���c�~��O̟����N!����0��J�Ԭ��P6��6�aa8��~�̇Z��3�y�+�N��)�Iǈl����n�F�v@��O��������C�ؓ�'9��4ɶ,��	�=d��$�sY%J�`r�aY6����N u�����q������:��;���_w�㇙���ߍw^{�
����p�	Y��u�s�1��<@�;܅C�'�,��!�=d��c$�O��T�'^0��t��Y8�w)}������=���7{�~�B�x��,��&�>C���
�&�kﳬ��a��ì:�bh;ܚI��;`��OPY����'�W�G�B>���-_}�6+�Q������w�ߺE�׉?'O�OXOSG��>d�!��rz���$���l�'P��󬒥a�=�Ad��;̝I���ܞ$�'�Xy�I�N������:�/�Cev�/�o��m�_u���,��j��P>|2������,8�<}Mo!�'y�'Y<I���@��d����'�u����PY%O9N�m+!����{�.E�R�?J�I���;�������Ba�P=@�����l�2/�d�V�ğ�P�	�:�<���0�<�&�:��>Փ�~d�����:Ü��f��o�s������M2M!��a�N�d5�p=a�O��{��y�����6�Ld�}�ǩ4��2OR���d:Ì&�ِ���(��<��j��?~3�z۟o����|�d�2z���~��'Pќì�I�w�u��XO;�d�'�{�2�'�5d��@��OZ�����!�?2u+8�=J��o/�8��d�|h��j�� }���r5N��D�SN����h�bQ��u���(b������ĳEJJ�X�FD>�&�f�8�^����֡�Q���c�m`E�2w�
�{��i&�{ń�.���/=uدR�� j��r��|n{]���;Z�U�}�Rٰ�$جɻ�3�������ރ]�0m��g<��J�Ԫ�7��p��h{��]$���z�2�h0�or�OV!΂5d����[-��}|�dգ�y|l>�gV��<pҴZ���#h��%�ݜ���_Fķ���*�P�b�}�!&M5'<��2�=�F�C�.��0Y���a�b�;�׷&����z�e��g���9n�}77�����/1�v��Z�����P�)���g*��:ˡ]d9E�~N�Z_n����3u����ctRn�ć5W �J�:Ne8�xne0:�7�PO��_f��]�E�W6��2s9�-AjZ���c�$�n�Dvۊ�L���,<J���o�Ҍ�m�������	5�ax��78gn�C"�n�UjBy'*�,�]F���paWL	�Me��b���U�����h�}p�EM�ݻ�E�������L�kXɖ�i�W\�-�[Ŗ���J��
��V��rB���7�q��ٔV^�Mh$�oy���
a��ר�r���^��y�i��.�X���R�Z"�;���ky�+����J�dz��<�RHV_z��@�#43�S!�0��wb��]Z�'�}*i�(��C+�?5��zW�Y��u9n��T�ל�)����J�/f��R��OժL��� �9(�	9�]�Sͤݚk����!oe(��9��WQg%Ⱦ�0E�v�zϏH��b��$�}�X:��j:��rgQZ����Q�{�sf��*K�c��ϭ\i'<�Evˏ���L�i�Y����fпA���g&
�hRw�_m�I��'���������w�>�=*�������]�쏛˝���;�5�v4��dP�#w��[�v��55����ҷL����ጬ��W�x��i�[��ly9�Y7�xg����6���.��ƌ��v� ��[R_i�%�t�ͦ󯾊=O]� b6�]	�h���D"X��u�)�X�q�j��(�.�[��ķb������gU'x�Pp��k�r���y0	��.�����9wb̓{�i�s�����N�qU����Y�џwWI�� {�x�M=�c  w��K|2��=VNd���v��:3?�w�ZL#FiN���d��!��iR���.�:��Ö�V'�ъ��\[�΍^ꋹC��^���- �#g����q��n{����cV�6�UK�T#�p�Q�Ӭ$T��J!{�S��]0m�hIL� ����胱�6�7�ݎv����j侳B�Q9�RA�P+=�1E��ݬ�9�����cǊ4������{x�7���/*K�!�A5A"�MJʢUbƶ��XPEEEkb2[PT�be��2�9JcQTQkj�V)\�*��&�q�*(�Yim���b�J,Qm�F���bPF6��"�[VZ�EAjTSk�F��9j���D[J"�LseDr�qܦ&EA�˂�*�-��&&1����*�3)Eme�m�X�i*�⥙KQJ�P��Ls)�J�2�663+kcZ�Z+���(Ŷ���#���9D+Q-�LG+���ZW2���P��µeV�e�DklːY��U��Q�F�Zƍh�Ъ�i2���F#%-�B�6�S�U�����ʫP�3e�VTR�m�UV�j�mģ�˕�
DA���aV��F,UŸ�51L*ڥTE�\S*���j���(��\l�c�)i\a\Tm+E��q.P\���Ŷ��TLJ�6!��UQ+S)TR?Q �Th	 ���v�k��+Wۻ�>|r����u��9d�븶��٭b��sw�������b�Vc�QL:��c��_}U�l���ϼ���AI?���|������d�Vk��N$��a�i��t�&�|ɾw:�|���̓���Y���u��t>J��'�w�:�}�3�����rC�m��V�N!�3t8��w[�2u+�R,:�Ԭ��A@���'wd�a��@��O�<���']���W�C���~�/�����&<�2w���q�㶇�Y<I�h�Ch~d�h�bI�f��`u4�1ћ�q��X=�a�N�����!Y9����l�d�(�?}��>�kT��{?~����W�}�0��sXJ�>O���%a�!�-:¤�֐��u52��m'A���I&:3y�s�!�y��':���w�UU�F_�!7�����R��}�	4���m�&�i;9a6�̟���d�����*
��'Ryl�I�N���M��~���4�q����N��� o�^z/=�xg_�{�l�����3	���q�ē��u�'��I�|�:�d�&��M��'?X�N!��d�	��6�d�VO����&�Raa� �uw����A�$�����VΞ�mo��[$�;��ϩ:��d�$��<��4��	���d����ܓ��M���v���;���q~�T����ވ�AG�}�����}15�PV�d>�=v>������^�a��n�DD.=�t���w�fC^Z�^�)7���% ��~��eH����v�T��cM���[�;wʦ�VqE{�QI�O���=w���k�b<��M����F��`2��Mf>������O�vx�:�VM�=(�T|^
@�E�5_\5��E��#x�h�-�,C��m����;��s�/���T8���K���!��e�5 z��|�3���ũt��;�����s�㮱��h���}U�R�����Ub���<�~wS���\�y��G�⟏*e�dRk3V����{��]�,{�	]��<�.�u��+�·2���cۛ�%�Wr����
�m&����=��E�j1�7Z[M+�Y��~����Mp�a�E��8�R��r���Zܯ%��[��z�c��s7�#5ĕiJm��rU�T,�)��mm�����U�F/;�9�r�	˘zv���ۇ,ao��i�\>H:�r��m�'y-'�q���W���c�����3�J]�>�S�����H;�?yY��;�u��%L�(^sc+]I�Re�a^˫]�z����T�H����W��+�����y�,�y�������ZN:��<%I��p]O.y炙��)����آ�:�	α�U����Խ�Ů����>��d��y{���}��jU�r�B��n��+�F$�=�i�7�i]Hfq`>ō�,�9���>�vnNg���H����L�^�����j�;��DA�����-W!�޻���9T��.����m�d�{2b͙���rKV]t�k_%\�^Y.��;���frޟ����>y�Ϧu'����w�=�ӏ�ގ_���R#\�j�Ui��׹�\�@g�4>����y��zX��ë}�Wzv��k��l���n�y�OqV��n.�,��̉;�䳂.������X��T/���t�v��P��2��(f���B���;�==���9�s�&�g�ΛN��a�c�=S��txA���X�p��Nk�q������d�rr���UI�}�v�o������as�a��򋥮��������iyd�}9L��n5ɺ���v�m��Z��5λ���*�s���wkT�yV�S[~�w�r��k�ޚٙS,�ln���c���ٚU����K�̏�)����[�Q��eL0�%����~��:tQ5����Ƙ�O:�!�Y��9�ݔ��w�]�K���s�{h�knVWSQ?Q5�]:;�I�riw
]�v�:�6wmY9c����J��UС�
�Vu����Up|�b�����[ڲ��;P��=��Ա�ں]�W4,�"�����%_���<���,w߾���؋�9�Io���6�:x8���~�ư�V4F4��L�Ԣ���Yz�#��txH���w���c ��q�9�A��o�Y�/���+��7���`n��62��ON=�o^�����>���1��hk�{�[��9�>#��Z��=��g���=��1va����;+K������p;2�D!!s�t�=�]�s�~Qoz��d	����l�d�i>�=�ޫ}^�U;���0���~�d>x5��J�W�;�{�	����O�?{5C��$�$ږ;%�NuX�v���ŏmo?o,���l�3�`>fXs#τT����wN�a(F{-��;��t��� mk�2�&rW^^^��<�J_G"���-��/��wM]�����2��_��ݮ[r���}Ew�/zS�2z��#��I�ܕ՞��,e+�oj}��������1��Y�'�xp[V���Sh��ŀй�'��hνMܧ>5��0�u����'X�|�y�W>KAtt�����;���L��!bl�e%H�c1 U��p��!V�3+���[��2gw�����Y�V�{��;z{��j��{J~>T��Q~r����@^]�|Gw�Ԛ�vj������'�ʷݴݡ�����1９��O��"��}�8.���.~\���S���ر7g��Oj����L��=5��t���co�����û$�Vz�I�X�Qs7#���v�����i�ڗ�7�c3E�]��*�f:�~�y��{��=����M㝮�	2�՝�{�|�g�u�c��|7��$7�A(G:a}��'�RC$��^����v�7ƍ���U�{jaϏ63]I��<{٨q�����}gq�p�"��:�ϫ�GË}%���{�X]���^^��껾�C�Dqtǝٜ���*pt�9����c�b��HL�Y�sr��7��ץ�9�u6�/>�&^N�v��{R�[�70��f�A�LJ���X��*�ʦq��$��m�R�}�f�E�	�%ge�����]�ԛeu&���v���
�4� �
�:RYݜe��P�L󰯻����k�R}�oZ;[�۰q�.���Y�=���^f.�y�*�����߼?k����~��x�����x%^���k$�L�o ��OmK���c�I�1��g�j�8�6}M�钮<,�j�Վ��K��]w�8����i{�J��=)k᝞���zB9)��ͽ\�{�-�����8}gX�I�����w��;R��v����x��_�C'��7�rtp_͗�`t��X��kG�Y���~=S���1��aG}*9�)9B��c$ևO-͝V�+p<���c� �%YO��ڗ�t�(����rAa�3su��wk�2iy=�r��;�|��RS=8>y�z�$=�c��H=NpN^����{�y�`�;��u]u����=Glz��Z�^V�/�1y��Ͻn*x��E̱\�_z�X>�h���+�+Ί̠;�;mC8�1B�8lbCc#��Tvm��59m?�笸Ǽ�g��1B �A4]�������AMW9V}�Z�yW%��v(���m�(B�?4����2�)�ͽ܁�cʄ�L��x���v�31��p�m�N;`'N��-��x,�-:�k1�����xV������W-�w��^[��L^�z�;iQ��h�>����T�R�sc�Zɹ=����B�ߵo7�R��H�?D��No�WvT���W���	��Q�D��n���=���j�ǌ������3������Ϩ:!{��Ջ��nxʪn�6�ۨ~��\.L��a����>>���]��giIl2�WDx��f�:)�|k��p~s���~�����v䘮h6v�aK�n%i����v=~��(m��CƂ��b���<�N��/#��W#-c����~|�;;|�c��`m	b:&�l�/Ҷ��ŗ�U:�X��>3�ӡ��[������7��b�/��oh;�}��vPO�F+�������]���{}y�����ծ3%�R�}�n�[���ϩO%^�]���4F�~�����z�����}�8��pc&���͏3���˸�̽K3����-]��r�oS]����R�����i���Ц=�po�"ܺ�:���[�)e���d��~�Ջ��s�_�����,��{�siǅ�̜�F[��U�9O�x�9t�/,�i��V����-j�8��SKbr/�}��}_=:��.t�Rܟ�OD(�����^���>�$�7�N�){�� ׵g�o�i��;�v����{/*݌�[�H0z�X�_�gt�Gr���ul�R�����_�^�:�;�4�/K���Rnp�/;�>�Bq�fu�H�8f�כ͸;����y���}-Y�;M;[R��__��C�8dT��QyR�b�h�H=�99�8��F���aV���k|���g,7���>�O���fƱ!��	Q�pN|Ǡ�-����%S�'Z����珏���m��vyڵ͛�^I���߷�q��S�ސ��Az�U�S��y�*X�(8G=�֭t{��f}���w�.���.�j��g?�s���Z�'b�N�|+���q=1o`�s��W�\��U�bo�&�q\�b�v�T�wO��Q���}��^�=A$^��_�Zo���)%�U�T��Վ�*JV8���BE����}�C9�����G-k񫸎lV�|����-;�����h�ht�~+S�܁ͣ)���Y��Ɂ
C�IxG׳F/etz�!c<'���DP4o��WB���Z��n�9j-���|y������>�| �Zu= �y��9�d��Ϛ��_�jXt���K�3ح��q*�j1:玵9܎_�|��rdx"��
���Ӱ;	}�,Nǥ?Eǝ���"��w����3>JG!��/���+���.=d��bǢ=�P�>����g��+�����M\w@/\�q�^�eq�,��S�C�����_mӱ�s^�/��lgc���G��OB����*�w�5��Q��bT~h{�n�5��Y[zZ��Ǟ�R2�W�6B�^}������O6es��MF3���o����o*�������9�M,�����lb�Վ��H0zܰ��Ǯy���fp�4��eS�]��y��5��o��b��b���-9s���������7J����H�T��S�x�_a�Y�)�*���Hld�����NU���e�[]��mM���yGS�ｕ|//=ɬ7�����OR��r��mE\�k�3�r��s*�l��ў�@�owMK��7=��y��vm��k�4�����w]q�A^^ �e?�t�mV�#�5V��"�3=�������=�Q��| ��[���p������:y����ژr�65Ԟꨄ�]h�Һ1��/r���ܔ���WvT����c�}%��;�֏G�/=�{���]ɾ�{���p��=��L����N��Q
qb�9az߽��t�om�u~���ͬ��]�����ے<��&\��a�vB| [\�t�z�}8���<z�Ʒo�d.��fN<�{�"����}r/K��]�W�'O"�g��.x.��f�90?o�x5��|�d��>S���<3����<//���}���s�UV�5�62Լ�Ӻ�yI��<ϒ�]G#mٿ�fvC��=��X#�xX����ez[]-��9w��������P}�Q����]��|��k��о���6{~h�~�(��K�M�J��^k�0�N�x�����?|�p����bO=�����`�����w%CSǅb@���`�d����Tǂ�b��0�"�;������]�>w���X���!�O�vu�9�n.J�����#q�{��Pش8L�0�S)a�j�ra@�vo���$됥ϡ:��j�
�t.=頋��������B)�ь�ql�[ӡ�r����u+/�U�����-�].�8�ǟ�q��-O+i;7�Z�5�����cPXK��w;���W���'4E�{dMl-a��f��oe�F���Q����6\ﮤ8��f��ʋyK��[]f�jhRuJ�e�?,��j�2�0փ�cm#l	ܫ1��*tq�֛.�a�y�4�<z�u�S�ly�oȷ�H4�$��	�R;[V��"`��,Q�
m����=��ҷ}���0'P;	��}4�ߞ��97�e�p����ˮeJ9��������w�K�W���Rue����MS�UXF��_����4�u���o�{f�Z�5k���&��u"�ʣѷ�]��Y4�Z.���ΛO�ǈ��7{����U��dv`���E�X�W��ҡGMR':k=���ӵvP�����D���f�˕�n��0�U�wp��E��TMvN�HwP+R�����It�l�޹&r/�s:�n�6�:����I%���
�,"J�0c;X��qŊ\�i�J��^Ρ]V���>�q�h6,�@s:�'��B�9}�k3W����
�]ϕ����
���k-0�����}���kΦ�:�P�G*��^!��6>��9k��n�˻�n:��1�ךf!WB
;�W<�H{Gf[�i^u�ב8�\��Ӽ�� ����3�9�,��:�����]^qt��d}��EA|�X}Vq��a�S�c�����������{�I^>�/�܍��RA݉��%S�8p��yKD�� u�۬;u�g����@�ʜ/q���I�V�bf󎮍:+�K����Ǻvw۬���d�7&��j�]ܧ2�7ⷧ�?X#(�ۙȕVS����~�=�~�ac7��εi�����˺u�J���\T<'��u�x1��դʄp�(�K��p+����_Z7�yp�r\C�����F[�x�9��f��w/�P&賂�RWy5�c��`��ǰ)�,�wS"�ԍmE�K����U��2�k/m���,`Q���2�|��+/k��_o�7��=��lt�#y]c S٠݊e��뮯����ڰP��]Rܠ`-����q4�Y�t���QRJ�OE�����ר��z�T2ﱊ��c��V�01'�i���_���Lԛy�m۽ s�Q����mVN�x�Czgq��H�d[zI���նά[h�5w^)\i��vgЬ��V���T?1\�r���P�����9<^���=.b6i���r��YmAݍN�"t�&�J�)m��}eʈ��mJ�Z�8��5����"+XV��̠�2�c1�r�TcU"��+p��m�QPms(��j��J��֢ZU��j���̊
��YF�b�Y��ж���V*�b�-%���-�ŕ�fS+F�bV6�)����j�W+�b��«��d�j��r�Q��˔��f�b����`�F��QK@�mV0���EiR��+��)�*�e1�nQh�J��*�+TV1��-"��ʒ���2�G�USb�YZ*�\
�q(.[�E�"��T.ek��R�Z��-2Ջ��b8��A-�s���j.%G0��S\-�����"�S
�[iiZ帴�VU�(��
����0�ȷ
�Um���Z���.����m�ru\�P�-�i�riX��oC˓��j\�T<�[ݔ��	���Y����w,5δ��.e���'�^������>�����RiuU�Z�����璊�Q�֣���M+Y����!�+tu�M�|#�\�?]��M]t���l`��[���:FlMq$�pi�p��>p7ZϤ����-�w�i��(��^w8s�[��-샥a*�eF�W����}���v���X�Ɲ�����|7�H`��vs�w(��5~��,�#%����s�����R���ÁX�|z�Q*eU�C�]E��I;�rU���R��Ԟ��Bs~R���`WN­�ckp����ӧ��Z{r��a�-~qj�\�瞩�� ~�,���b������d�/�Uz�[�1��4;�F��Y?G�y{���d�y:��ڈ�C�x��}y��ֈ��)9K�y���.k�����r3/���L��Y�&���)�Vn���vSvE��ө=���y�=�#J�N)o�q^?z� h!�"ǽ��>W%G4���)w5Z�b�;H��X0���o_q��ٓ2�t��ê{�ރ�!��Y;Cb�樭��KiZ,���t���ڜň�=}���p͓��ϼNA��W�18�������ܷھ���z	�� �s�?�5S����BX����?J�Z���z<c�DBz���u{\�)���9����*b�����t�v��ONw�ėf�m�O'����.<��O���N5�-��t����8���
]�����G�8J=��e�I����2N7���1&=>�t�Y���n��e��s=Awz�l�h���e=��̽���br�\`�]�c�4�l�9��df�k=�ޮ��d;�^NV�;������`�P�V~��վ�kѣ�s%tpؚ�{oyby�i���OM]Iy��ucr{��  )���Ʈb띇�E �q��留�Sж�|Buy%�}X��ڭn9ڷ�=�g	���Nt���ߩF���k(�WCD~^��0x��h��}��wT	O]H_8u�}�J9�h3���;�	o�?�3 ��_�[^%xf�܃>�v����GPڔV�s��W\y|�vڑ8fI��ey+��eB��[[D��kK��z�u�ltɱe滾!��p2�_tS������Ȋ	}��Z��|yw��r��Q����삵�&U��2w_~�������OO9	��h�X]�JeK#�_�[8�{=�q���U��WbZw'sU���������W�z<�㛪N[�`ڃ�o�X�}�qs��N�$�2��:/>tB�q�����^�.��<侹��N��;ݥ�>��%M��<�%�`�U����O>���{�L�|;�p�zOz,���t�C�����W���~Ϥ��$�A�Pl��Z^���A��)�j�}k��6¶���'����Y�-���Ӿ-=�3���g�>�~�#C�ό}yV��5K�Ġ
9}&:�)��-�w��� �^}��-��;Q��u����ҽ�)3���=v��g�*:���N���`7帜�oO�9臧,�[��l��^+~0���|�{���=��pm��"�z�ṽ�/��I�B�ݺ�׵q��3������c����\��M��9|o["P��J-��b�G׷�ж�T�Y4��<s;��[4��#����-�o&^ASD���7ǋHZ��[�(�g#�]Z�o#;���UK6VM��ĕO9�O��tR%ha�6Vd��-�|t؍Ί�hoT�8�~��������I�w�n8R�^3z��*��/SQ���-�����E��>������{�38�X:��O�.�V��r�r�#��<��^f��]��Q�/gD�Nd�3k<&-��䬭u���὎XN\�zv��<�ᾋ�n�fea���-�"�m;���)����󦹧��I?s���yX1wXbC��s��dau;�/;�KV�é3�Z�]�<�͚��O8\S��9��p�}A�����,%���u�'k�����싻ݺ�����}��qܿz�Gp����#̷l��=>�;�M�Q�\Χ5�S��L���������K�r�����>M�vL���h�}GI���=�f?d�8��W��K�%��We�/}U�}��p�,�^A����ϭ��l��vc������w~��f�B��s6�g�e�K��݇��|=)�����>{-ú�C���V
�u9�����9<u��
p�KFg����X�)��K�6EbB�(�'=Y��� %���:�f(9�w�Ψg,�gVLP�b��)tYn���]߾�������;h��xk��X}D�g��OҮ��b��n�g�@9+wK^C+�����i��\���Am��a�t�Y/��f�<[�^����'�f�d�;C2��|��^�nG!:�;bB���N�X�8�nK�l�,��]ck�;ۓ�W����7��ӧNP�����Z��u��j/����(�m����d垠���v{VI���W���#��MF2n�����l��鋡��gd�f�~��4%�_'����;��m�=n+7�g��UY��U[�Ia�^�fu�'� ���7T^���ub�������G�`�)�v�J���q݃g�������:~��ӷ3�8]V'W�u86�w�;ְ��y��f_N�Io�ၿB�Nǽ�z��������:c<�>���Wx�v^j��&ҿxПG�oS��eK����No�g�u��\�!c�B��]��%������w�ǜX��V)��=g���
�`I|�`nN�}�7$�U݄5����JWB�Tڤ]�U{�����Q��'��0�
�-S�!��z��^�Q:j�Q�s8�E���=�!����!9�3�. �rM�ݜ��z{�U}�����{~n5V��S�NZ<��nl��\�>2�WOe��g��q�h��%�"�>���+���'&��g����{\�.�1��������k�̡�B�B�|���:P�qw�7<�I�%i�Xp������]x�b�~��C1?Ulw���P��/���U��l<�k=4P��L��qU�������>�q��d���BX���g�~����[ekr�ǫa�K�OYR�}y�@��2OG�mԁ�/��e����O����KL�y��g)=����N�iE���jO]����lH^�}�]'«)v�2�G[��+��N�-�GW�!ZQ�)x�����x��k���TU�%��Y+�U�]�js��{��~f��W����m��T�?T��gz����]e��E~<�-\��٪��>��ϻv��M�-۴�X9������{�s�(�����R�-��]�YT9�T:�J	u�ޕˌ�Ŋ �4��t�u�y��p�����mm#�b��B'^^\��S|�l�kۭ=1�#��L�t�?���]���^�A�j��ڳ��M�q��M��{��r�$-ף���ީ5J���G_{������vI���g�nk5�ٹ�w�7����;^�a=6�K=�Z�w���o��ӭ�	;�ϽnXN^�tk�D�[Y���/�[ώ��%^�������R�Y�n��ΙT��
Ø�R��|\����ߔi���[]]�?+�·��r��a\.�}iк�pf��zTQ�sD�Ԯ_���R7����\�����O�]P��a8{���(�c>�����������.Μ,�����׎t�ht}_,P�XC��Z���v�*�h�h��ׯE���0�=����<�y����_;.���`�y��Ҁ�qsʂ����6bǕYx��ۚ�)�M�$y�.K����<��	��|��:�\��
˜w���Ze8������y����ԿI+äږ;$&�U(gEc{�:W��nmX�ni���fS�&I��P�^�ʵX��hr����K������MK��"�ѻ�L�t3l.�u:�w����KQ}s��,J
�Y��9���m��Č1�[����)�����&�#����f);���; S+��Gd�kX���k�)S(qv�{	�tG=��1e���������t򂮳�J����,��{�����f|��9}&?�5�>:.j"�Zu���_�O�����~0��u<�߷�'{uy��:�9�b0���~��|$�:8/�����6�X�9�l��m�c�����u5~�X�O5�WW�p@:zXps����Ĝ<�o�h5�9����4��e��x�R_i��E�5y�~�9��F2nķ���/7E��;Aɕu�F��f-�)��>�}y��z������O8�ܻS	\α���x����@}��X��z�i�~����XN\ϏN�t�i��uw�ڑ�Z�/�2�	u�\�����������������p�Ω����TyoT\񼣁]b�v��ծl��0U�QD�������J���q�'�����ݟL
݌CGR��2w��=c�*6���v�K܌��k�o���`��nV�e�ƫV��p]��^�����mv�g'��hx�-�^OAx��ظA�*������H_��t�ֲ> gZ�j��x|Ҹ��w��w�ig7�uW;$�;�!�ݘT��{B!�XV����g{�y�wꯪ���2�Sݞy�p�C�Xc����w�;��>�Gpu�,I0����mS�q��:�=���Ncj-�S��$~ɒfD[�w)��|Zw��e�	+��cw^��7���]�f_fw��~�^oT���sg�`��~(������;{�MG���=�����J�:��T=�ްy=t�Z��=K˅�叅X6n݋�r(����;B}�
����촐��Ԛ�/��Ez�y[۞��|NoPBqN1��A)�^|�[D䆟"D9���l}�J�u��g%5����Ʊ��9,X����4.��=�[9�Y��."���� (��~K:���4a�9A��n����7W�EP�sqݦ�ݩ��|s��L�Wm��N�H���ejz�4��\n�eﮱ�Q�����+.I��Ӏ�g. ��Z��9���{+�@`��`G++}T��'�Ej��&�%��߯r=�ޫ��1�80����MyX.��gO�4xn_��f`�vFӱ5	�*��#��G��*�Ø��ˎp��Ł������s����̬>גY����]��K����=���W�5�S��5�怩�]�bdסs�#�TTo���G�<S��"z�L��r�6hYN=�X6éQ�W;�ܾ���}�}U^���$�g�^�V+��x�����[��/v����7��.%,i�ٴ;�����0��v�g�8��¦!�;�*��ue�eT^�R��aJ��X#��(�5N�T��6-ދ�I��Z�m�eӹ�NX�^�a�<�y]#Ġ`���U+�)w^?�HOoz��w�j��q�
�]ɥz��=��	��OS�~
W43�P�ɘ���f���ۇC�<�����g��Y�K�G��-kl�,�S�}%�sy�Š��Y���u�AW�- k���˪pU����ċ
���	�c���T�5�L�j�ń1�~��hf���׏}��H�S�D�C�!��MrQ+��ϨS2���P�iԗ��歫e�Z���4�'�9�:1��7�T�f���(�ؾ$���}Y�vr�K�t�i�䟨�,J8�>ce�j�:Ñ]��Umq�"�F(w�L�aIt���F`���
u&;��j!	&�H�����x�%dA��]�pHj%C�uFM#;�#M�*b�|O�]�[k�m>@aGBt��.�)�Ŧ��[�`x����K�����k�)r2�gG>i.�ݻyqs����te�B|WnN���/����M��-1x�o���
�̧�4���SK.�hc{���o��+�o�ȱaᗶ]�-��z�w�v�$�	N�^�l�;���g�Z$�Y��s#��[ע�u�Cs���lB���(9n`�c���=��:��Z���Wo9���k흚�A�<+�=S��<��$��rJ.�4V����M2��,�V���7�y��l��Of�<�=�uo��E+�噽Ea��.`ՋK��̰���'^��������h����uOy��F�#f�C�⩏i|ń<m�|��L�]֨f�[Lq�s�w�A�$j�/,Ln�쓡^��FsY���x����;r��<L �:)��"�}2qo�+����X��tk����;��
���(�w`� �6�w�nLEgu�'fc=�
q��(rc+h�r��)m�L~����%B�ÂM��S���zN��B��ρwo.�*ۙz.���lPw6�KTޑ79��b��۩D���%r��dA�� ��۰d�B`�{�ԓ�n�s�\+-��2[����<��i �#$|F��Y\w�)����tn�LWKQp���w\ ǘ�#���,��g��h.�]����E㣒V��&�vZ�X3����g �l����,v��P2���;���V��P�K��}#��g+��A�4�	ww����|3Ͳ��q?z]�k�r\��F��o8[�u�F;Ho�+�V��[Ԅ�S.,�`*�,i��(������Q!�����S;
�1K��Z3S����mܫ��ş1ҬBw&e�i�ÿ)f{������ь{��SV�m�Tѓb.�.ue�7k��qK+1v�]Sw.�H9m�.�m�hv�P�ju>7��`�sI�U7�%�t>ަ�:U���\9��B����\��9�Tͽ�Cγ���!���"���Dք�3�e�I���GlY`[]CJo��z.��m1�����6��_L��!�P����°���hb~zf��ʰ����q����K�s0lxE3m���"/��ć0*��ax�z����Gȃ��tYn�kv�7�8��e�pEt�kn��z<z�}��3G.�v��,ǭ!��y�"ս�᫂*:h0o�{'�r�5Y��x������2��V��Z��"�e�s���2;��F����a2���b�K����@�l̻�ְr'��M:���b��}������43�L+�/TG촘�����G
"�+G<�5���Or�>Dou����љ�snV]L�Xu������yu���9a��!����Z�����oY��6fZ��n;��&N�R�oA�J�Eu�ˇN��u��#{X8>�G��H�ƹ��ˎb\�W.\̉e�K��
��" �ƪ(��(��iQ���Elr��-iJ�Z�j\�k�2V\̆5R���en*�-��ҕJ�\�(�-Q�1�U*�)kr��bZT�[J�-E1.&dS.8c�ZZ�)Z��PS31c*�cmZ��L�������aZ��QZ�fY�����1�����̦V���s%UK���ER��9J%�D�\E-���9b��3
�0��e
ۘ���c.,3�����q
�㊕+X-�e�*��8!��X
U��j
��Z��U�֢�1�W-��9�T�AAU-���S-r��B�a�	�ʸ�R�0X(����[s
"�UQLb�*V�*�*��0q��d�e��E1���j5+"��YR��D�)UQq��*�R��*�b�s�@T!���ц�΁�j����M�F�u�S�ׁ����x���r}e�{��M�]���pv�w:��f�i|�hN�����꯾���~mN��.ϰ+Xy�P�}��*����*Oy��Ie�>y��gz�Gv�./gP�j�\�!˺,m��E�i��_��Z�t�K�OX`�׾�ks̋�����K%��sm��>)�7Z�:>U.|�^9��V޹���R�e,q��.a9�a	w����wu��w�7�0��cC�,'�3�G0���$�������i��#u�'>]3�6��!=�p�C���K�����۰���O��*��a�˃�R�v1��w��UbD����8�,�c3;��w�дbwk�c=��\������)]�LK�k��ZXZS/�b���F(��$�\<�<��懞��c:5g2�-�����Ax�Ä�^S�U\^}0�x�ltL�lF.�qbT<�^G���~���k��vb�gU�q�Pvk�P���%\:R+GO���Y�;�#�&�u"u�����I>�%��:i�G�K���Z=<.�<s�&��
��S�G����Ɣ(SW��.�κ����$ŝ�v��i��7��}�W�B��P~��r��7"��S��	@�10����;�u��yF#���k,�Va���ZgQ���!vNq����Ts�m)�p�����4WYKoC-�W��y�\���G)���}��e&����i�ߏ���r'K�R2U ~� $�^`P��Nas��8ն������R\c�}�)�ؕcH�<��d��^�f�e��0�5%"N�7"�<�/�,N�{;�E�
���8������#�r�<�ب_�	*b�T>70/	���V����L�9�!��}UP��
�n��Mf.,���6`{�Wc��ih]C6��y�^y��|3���o��-Uw�fR��I��µ�c��h�6d��6��׈��V�����T��*�{A�Q#��'��]����3�P����M=�\��Mg[��|&M9��d�.<޼~~ާt��o<%Z��&Ě�>��o�׶#ԯ�/:����(�w�i��~"cX���u͢�hZ%{����po�q�9�X_��դmmthʅ�Wye��\��G��Vi�oS�ٹ�f�^R]i��=K�v������~� ����)Z�d����ta}v�d�����p�\|�%�7����A��aŔ�`�P�Ny�/�+~�|�t?��d�^��`���Φ�Y����u������7�$닩;����[ڱh��5m��`�0l�/f&��6=�B-���ǧ0�8�|��+9`��'N��F'�Ǆ��]��ۙ�8���d޻�֣�d	Q��۷��N�Lu(n���߾������P�w�ƛ#�Z��-4תW������"85�0��38S��p�~���F�������ޯ*�c��"���XE5b��y�*�t4�85��"{�}㜋9���c���$@5���]���1Q�*���Ƅ6GRh����K+�1�����qr��s�-���d�hD����&pI��_J��L�zĻG�������֎�t� l�����Nǯ��o�5���0�7��Vzx���:c}�|�7ё���
����X��dc�ߪ��L�e���#�sSu/��
eIn-�R�����<q����k�Щܑ�9L߾�R��D�f5�
@{8�x>�1ݳ�y~/APߑ���(fn��x�*<j���,�Ԡ����T�ZV)�=Y�w+����e���d���+î17��3���U�Ϛ���%-��Eb���e��|#5ړ\e�赬�P{<�v<�uG�z��+nS�6�^	V�2�!���lvA�*��Yc���1W��%צ�mz�uc,=j��3�!�&�](oBu�P<k�X�gT�͋s%��MKb�&N@XlT���_��C�}�+�+�W��{�7e�A�A�n�y����\�d�\�[Y�sz��C1X��/�<�.5r�tz�KD��C�g�O=�����}����
�;�/7��=3b�Jdf�+אlE����\��|�ц�4�����Z�;���re��}�q��y�xv�b��c��8,+�"Y�XG�u;�c������b�u�"ȼM+9e3�MXY��fC=�o~��/�౸�4����zy�rAN͞�3�=^�/a{��0+�C�-+r�3�W��v댈��ff��OiΜ�_:��Z�������D绊�ڰd�g���_��pSQ�VW�>��e\��sZD��b�g�< �Q7d��K������t;P������0VZ�'��i���*�&֑���J,�_����(��jPo
�,a�b��P����}i�yl�VZ<O��J�)�����7ֶ��uU|�}J�"����9��Y9Z�C�z+p��ҔG{�b>52Xb-yN�~�n��<����8�����bK�������#S�G��l	��b��3�eM�wm^��ڧHT���Wf��;!����A3;]ٜ*X��2���:o�!�*����A�ټ��aȓQ╚a�B�	�}%J����3�����LD�ͪ��_Q�V��w�Fw;�:�aɋ9�\@�`���Ruc�DqN뤶��hĤ:/�˚7q�E��7�^�SPCP��ݠ�9�-��|> |RS9���u�W�?	��n-#�Ph��R�\�J���Z	���iM�\#;�fj��=�'�~���s7M��y���rL�7�����A�+�ϰO	�w�c�c.>^T��2.�%�[RJM%���Y��U5��E|�	P�]�H��P�V�RK��б-��o�˴8M��8\&���D�"�Wl��<0J��&]�w�(Y�Y�ADi��ފ�N�!���80��c�PL���MIƀ�>ϯ�%Z��kJ���@׸����q:o�����X�ND���Ŝ;c7q������C�C��_%����}�*�23d���[hz�r�N���p*{gOM7Z�g�]K�a���>�޹�5:���JfO�����u��R�ݲ�����\�9���L��ӏ�Hg���{
��6�j+���r���U<X6��0k��=,w��Zk�n�9��-.�ٕf����{����i��L�j �Ƒc<.�ǚ��f3�kO�D���B5�yl��Xjj��"�u��b��G$��������;m�6���7@ct�Š&w�������Œ;��ҙKM��X3J�N����}�y���7�^��oo���}x����v��|��c�C��a0(]�+��k��	��CapNE�ﾪ��s'����,��?ԗ3��.%͂Ōb��:1E��+�d:�������z����Ύ�љ7�A�3W�ÁѴp�8�$�yo�*s�ۢd+ �F+NL�w�[�?$̮�_�3�Ꞔ�,6�m�T�%�0O���\[�fN�H����{m�D ���3��_�F�2�B5�>��d�C�#�>K�`�K�L+�Φ���apL���+��oW7�/��Sm���3�}=��a�7�iȝ.)4*P�^�����.��2�0:5��l-��pʕ����w9?T�{*ƑrG���d��^�L݉�L2�%ݘk{���γ-{#����g�qͰ��W��|f������Uz��"�~Y%L][��c�{Z���x2{���+����4�}�I�UB:����n��k1qeEI����4X�:��[}��C�5m�V4�f����c�l�rYO��|)5��Cךόw̒�,I�|:�xo��/��+��P���D�|���v��Z�2�������ϊ��u�c��`�:G�t��,�nw��Ļ��玱���۰��yE�^��a@��ǯ�#��-W!�:��ʚ�}�!�����u�i	�F��y,�g&ɣFo��/��k#������7��oq�Â�s �$A�a {.�'Oig��  	�q��*��n/�I-y�%XLƉ�)�|9C��V&�Z���Lx�g����ɷ��v{ȹ�7����Xȷ�^����;��k��䳫H����:-B�].R^r>͊�G�o�{#�7ْ�
�<(��׭3�D�^�P�,�T��O�%�w*�A�����	����ޤ��6�F����|�T�}�]�u�D�aŔ�`��P�-רtY��Saڋ�8��W�� ���Q��Ce��%a��\�Q��"9�Ʉ�l�b���(j����߱�>yw��z�'���u�F|_°R��F���+�5]A=���I#r5�.U��ft�:���Y"�9�&�]����*5�*���!��2�WYdO|0N�`��[I�z7�y[6%����"ڝ�$�j�I��oAM��H�˴x�ɚ��ܫ䢽3�Q��6��>H��[���;z�,,��L�o<rewmf��v��!�C&��6�������gH�Qf�C����A�v�y?T�>kA��/�#�ųj��w���f�Z;��AR�J�^��[	SI�*���lKX՞k�<$:|_gh��@/V��-���ۻ�z�*�SVX9���o{)S���}<�첞�n3f�c��m�_�k�F����w��zj�WR������ Hg���2����U���}� ;��:L��,c_�C{)RR�$�k�#�ƃ,�)�\g(%���V����ӕ���a��sT��!g������i�Ө]��=w�O5ظG���מx�qE�_-O���	yp�]������e���v�댼}�7�Z�W��c�ݬ�4�G���-r����mH-�=�5�)�w��yJ�iKͲ�{Eu�>+�]rU��v�x�ϛ�����f��q�t����
7�P�o�?%�yb�}�gR�pxt㮓إ�NB�nKL&s�|��^��E��� ��m���+�u�0G�5�e�a܆�9L1� �̘������;��v,Յ��̆vS����DpP����kޫ��f����0ZÞ&7j��Af�ŧR��U)֕ys�^6�ۮ2#p���mdYQ:S���r�ق��wca�gr�Zu�(��U���	����r��6'v����(�w���u�]L�T��B�`��i��=�|'�̏�W�#�֍k�d�WE)?g ���󀐍��"Ί�f�;W4�o��{�2��OH�Zz�jn�,=��� ���'�J�R�� p��FC��oOC�4�|��W����]ӻ�����C�~��t
��ׅ��im��>哮8�pE�7p�g��-�Η�����W�ǜʦ|9&|��_��kY��)��	r�yw��=���FF�k��汉زwWt�'R��AYi�Q�<�'>�v!�L=8�J�z
ӆ��T)"r&1���1�>.��u/#
��ʪfWU�Se08����-y��o3t�~/��KSs�}�-7�Ϻ��_��^�E�x��A3/������`S/ڏ,�҃���9��z{�9�4懷"�ZGR������V+����3��|$u����@&x�Z޴�����y����Gzf��ӟ�a�d��oD�hP!�A��e.����S��77�u���=�4_;D�1K,�It��Vd/b�k������}2Ɇ�6I��:_t��]��띏x+�}W~<o{{^r�Y���Fĕ��+�	C��}�m�.�|nw�P�y3�.�h�Q��H��T,v�#��W���sJǥ2ɘ������'*r��t�&@�w� ~'�/���%e�;y�����4��֡��|��P�p<W� ����-��e�y�5��̨
�`]K����U�-,W��̉�3*��E]"D���2�m{��^��4Nۺk)��f��޷)K_�5���Nlfٛ�%j��mӱ$�PX��i���ç5�N��R��{|��m�?�������e�d�\���T����(��1��T�Ξ�n��>U.|�^9�����n�g�)38sKZD���z�� ��oAL�6�{���x�~�m;w9�>���/=|?�'?5,C��z%Zٞ����3�ώk��'���~�ۢ��Lr
�b^§*��b�o���[�.&8���8�Q?f32��^;�蟖Ov��;֯�
Ho�����~�Է���z���cbX�ĸq3}J�u*�Qъ,q]9��.y8��Y���(+�p�yp]�"]Y�[J)�Ux�YU\et�U�����D�Vl�I�<nN��=w�xO^Jitx���%�^�Y�]P>TZ���B�qx/�a��D�^��Uc@�N�I�{��gK"��/p���ς�Z3��ؤ.��]��L�G��W�����E_�59q^{���Za{�V��"�~>o<Ӛ>��\�FX�hG���:����܆��m^�W(P~����z�r~;�ʱ�\�����/�����,�g�w�z�g��KZ��)��Z�]���Ӡ*+��W\-P�6�=0��x�����$���k��Q���\��p�_o�� ���o��ĭ��t��{��<�dǋ,�m�����	�8��9p�`��I��9}�B��e�Q%/�L��R�v������u��?�x��;Q�Ņ�NH���cH���P"�շ�ve�_^����(��Y��9�iY:�݃N���yu&>�ܶ�h}�;��м6�"�^�3//O�н$�q={Q��m}I�����ǖ�X�Y��k�.��aH��e�C��]��7���B#�/W7��,�f�ZT~s�3��"���X�x�u�4����P��X�ẉ��Tv��4E�Z3��'�ϐJj/'u��
Z�F�u���WN�X�J^ޮ��C ������ZD�F���G.��ٓ���J�3\�2�!��^��@�{|���1�v���,�v�d}Q�n+Hؔ^R��B'F=Bfb���j+�v���#��O�v��r��n��f����/'ۏ��0VHe���{��Q�!w��糙�O	#Z���`oPX4*�|��$��2��&��n���v5H���Z{�V�b�^o�o�[xx�l;(�NΒd,q�pg��bc��
;���ju�5}�C����2�i'����� p����'�-#�!�D���n�Q�9sb�;��~ƫ(�.���O�|I�S-i�;\�:��^�i�:�m<\�i+Wo^[z�1�ϣ,�S	��x��cR{#�2
�lL��3���.����}ۍ[%�7	����f���xd��:�b�X9���hx8;-ڜV����ks��%�8�o1R�{!({+��3u:�\@�6�gM*�wqPe����޽��A�WVM�Ê�:��+mjN�����'�%�JR1�5t�˃/���V�=}/�3�x��~^�-�Elt��26�QP���.&!��o&4���K�:��]n�N-��K��K	,�P�*�=�cޣ���ͦ�N���V2+�B�w�<N^� �*�`_(hK&4��TYw|^
�f�yx
�ze�!���e9Ҭ�B�5���w��n��\+[��SE�bݣ�k2��S\"����G��+��t���G�#�0M�Z���$�W}�9��Ǡ�.U��é���s
��h�:l5sJ����,��x�ۆ�U�K��#;�kz��0��xL�yw��P�B����)���Q�=:�K�t#}%X���eH_,n��d'mЛ�FPV`U�Ē枖�����P˜%%��6yЋ��T�(���Nvxb�:ٶ�Ӳ��{�X=��M�<���z�f�U\��ª��dͫ*�4[(k���7b����O�����׫WK��bJ�ք~�aK�sњ����������Z0���Z�����z���S��3����[��g����r�j
�%T���UDT
YU�F�Z,�2�Qh�E�+kZ+YR�����+iR�
c��5��AW��"��[dq�X8�*�QVUEPUd*U`����k&%E+B�,L-b���@D��11
5
¥AdQJ��X�l�e(�ʊ���T��r��´jfD�kQUDV ���1�\T**�+
�PX(bJ12�bEF)[l*���+"+��Ad��R�IQb��[b�Q$V�r�f[*Lfe"�,�Q�mAiK�r�`��5�5R,%T��QeIX���X,UX
�U��AaKlB�U�,��YkD��VBT�FaR�#�d+���*�V��("�ʕ��TU�DEm
ʕ��%T*�*��X����b`�^�{z����J)_;��Ò5��!�l���Po���HS����V�ꕮA���ݝdk����w���}��vm��WqD�s�I�G��P~W�����)���<�ب_�IS	�����A�N�L�Q�ez�gl�|�䠪�u+!����m�j�ˋ*�g���Ht�n�k�î���xnq�imZ By_�.�Ǵ��"�h�\F�j��_9����MF�� j��c���e��1�NX�g��k��G[�<�;������b=aݎ�%��ˡ�yyZ`/����Z*ǜ�U���I��<a��*�ϻmj�`<\�;۹�N�:�����wӊ���}�1��W�A�C�,y���a���]z*��ܦ=�6�M�R��3�T�����	��s�,��F�t&�i��=Z����YЩ���D�ừa��uO{�f���A,��a�nҵ�kW�U���p����5�"��qe9�=�7�-9u�ۀ6���땖���d��׎�+�Ce�����,�G�6���a&�a�牂�������"-���V�z�h9���	��t��8)
���Km<��`��to�%��H��63������J�fG瞴FzF�;�Y��+���g�0)�|�����g��#�*� Q�6����]Ih y���V]��egMM!Ku��_L�I�I��I��LSS��UvP�lP}}�+Gd�k+���{U���W�}��X�w�$�F�[�,tH��s�M.�W�TjZ�ue�B׍lԞ<9����̴�s�>�^�p\��GJ�W[��&�&pt��N��l�$r��p�W�|F�6�ƺ^���j�{�pU�En�O6JS�;p��q ��b̙]�X�[TM�,5EZLq����T�2Y�hoR��L�h!��ޮ�M��jV�i�jm�<�J�ʭ�㯩^s���n��	bZ�	�i��D����PP��6ϵGT�j�����8�Tե�m�Nr�.��g:����)j��A�yi*�-$�.��}ްy?t��tf�����jgǚ�^\/b�g�%-�4ȧb�{&��-�-|h�	��{8��<\��Z����Ά���=�h����Um�CO�ϐ�h:���M��t�;��
��ߒ]��Ep�n;L�g
?o�ٱxt�F`��yFX>h�u���B��T�k��(ఄ�l�z�!�:�5�i�i��E��?z{k��8,+~���v�a��N^!��]7�{��2��]S�m��RC�砖�H�w�����4�
8�`�	�%yf�Pk w�:_Pз�s�<�r����0$&f��{o�|(V۶^:M8�����ei�GE������
�p�I�v��L���U}U�>!M��t��&@��l*�g����(��*�����[o��z�V(a���b�U��^�h^���z�C�sڴ=�׌�^]�uK���?N0�G�bsr��=1�G�[�-nc>�0<�3*]����(d�ܽ�mx��QXӄ�H���#�Mj���4l(!N��;U��3�sW��3���4�[f�{��P��h��	���F,��zgN�#��r,��0_��%�X�b���y3�7��X}�<�y��]2�����L�\G ���v�}f�*�e��؆-S�A��[�T�hm��M*<\�������� ����k���I�`�2,������
�u�Vq�徒��Z�ݨEyb{䝼�骫Οb��qfH,2,K4=n�C�H����^a�KP�ǘ�J�9b����]�Otʠ�A�y�&܋qh#�Ph��ݠh5�D�WS-�w�t��y��:�Ό��ʤ�I|G�ڒ��^f�9Xx��$��{*Z��:�l�$�R������~
�a8�����> ��^���9z{�xrX��6ѣm��p��Q������R�"���6e�2֛1�3��k��b]c9�93��#���M4<�gٲ5��T{԰�_.�����$
]��>�/X������5��*ں�?��iy����a~���f ��d%¡,��2�ڗ�@��xh2+�s�*_�,�Vl��35z���ݴ5��������Ȝ��d��B����r�Y�w<��VD���8���.���;S����vN��=ue����e�G��aH����.;+5��s�W�L��P�鈌P�luϞ�V�A��Qr��uP��ij�:��p���3��x[�u�+h֯^�=��t�|��N�ҟ{���?X`ȱ�K���e﯈OJI�߇��5�����=�:�﨩���w��y�ٱ���@�bu'<�'�Y7��;�)���X~���d>���G�|u�1��MKl�����v�J�@��0s��� ��8����#�OK�֚{tY��7��p��d�f�^�������타����3���㧢~Y�O �(�j�R�nX���J׌h8�V`LlK��^K���O�ԫ��1E�T!�t�d:*��oFrZ����o��(��υ�dz�f�mm(�
�1�]�	}0��� �@�Qh���ˌt��Ez�W��?G�C�# 칀��`ɖrQ�=aJC`\;z�{�yB�,&M��ջ�')�:wԩc=���Ϟ�.^m�)%(v��^o�W�4�B��S���=��֑�e/l!v���a�*brN�Mgj:��Gk<�|>��}� �����E�y�R����vU�l�%����oGG��!��q	��SW������yA��$`y�g�B5��'��a�����Nq��ؖ�P������%^�%����c��y�7 �ߩI����39�r���H��]�F�����SݿV8;����I�Y(Pn�a䡰����v=�U�"�w��KƯe3dX]7�u���{�5�����<,�d�Dq|B�G����)b9����U^Z�+�R�>�'R��c�����ɉ��|o炡����$�Һ�GR�[�n��Mf|����Fu7�ݐ?�5CL��^����9��IP��z�T�"���ֶ�3,�3���X�x)$oe�o������\P�ɘ�Ϝ�G��SU�]���֦ppSWḙV}�*�v�K���)����ۂ�5�9���&cD��M�IϹC�ͯ�B��3���o{fN"ٳ6!�h�W�A�C�/�;��c\x�}��"��H�xx���W���]8n�t$fpř�����;�$3ZC/�a�Fv�{�ݲ�DGsǽ[F��4RBp�#y�lb/n���o�u�њ;�z�c$�u܇],we>	s�H�
e&�>I]�W[�wn΍^�p��M�ù�3�[�| �u��d]�A����Wyf
�zg�W�}v!~�x����襯��E�n��@�����AH/JA�A�t�3��V�
��2��%�*a@_�]2 �v<����L��Cq�ozn{�:�w�#=��;NK�Y>0W��l��+�.X�����"<s�<����1�;-�����'I3���e9x r��r�>k/��a�!V�e�P�y���亡��7�����|�#>�"X6Y"�s�@�b���*5-C-W�:P������G�j���S½�*���P�ti.��S;�֋��8Ѷ�}�X]���G�ޙ�1�,^緧���\�դ!>2����H���`�����7G�D����>9"�Eڔ��Y�Z��ޜ���|}E�JQ3	q{��A��"��1��.m׽�S�%n�2��;��/λؠ�L��C�x<˴���D����PP�����,�,t�UN[o��d��X_�w���T7�T�,�RՉ���������u����;bI^�n]�A0#��c���]z��u���<�5�C[���ә���3tgu��g�ih��Ff7A;�w��\S�����4�7wdB!�U�7�m�;�+��Y�C��Q��M��D�<2���c��Sg͙��=:.�(��}|�!�d~mz�΂_Uw8�ܱ�������=��zEv�JZ�L��ؠ�vZHTf�UX]y��Gs��b��̶�˽G��b|�~�/KEE/��h����p!�uD3��h�q͑��;����ۥ�HC[���g�(�n�糮��ƀ���b����ʐ[D�T����:��s�����t�G�=[�e�;�}�����Pr�E��� ��մCul�����ϴΘ�zL�����Ab��"���.�x���^I�쭷�����I���=���9S��3�.����j><�^������^�>KppV����w�pߕJ|�T��sQ�e���[1J�3@��(g��c�����=��%Q#�S�]k��x���L��u~��
��s�\\K>�[19vg�v�'cB}�%���~���vj�w�rr���^�);@�mx�E�u�1e-vsw;(����|�9<�%nM���9lc�>����Ƹ���ڈ��h�AaX�iX�F)��	�d�8��](��	x߮^�q��ʺM���qwA^N�T�];��Y��m>��M�N�%�h�BRP:�����^ʙ�r��u�)�z�sY�\*�'0_R�Glt˽gK�4t�6U��k�pR4�n
�4Z�4�`a�@�U�pܽ�֗U��tyzx��w���1_��eHzB0>ahg����Ip���b���(1�b6�������[�	���l�{��Sㇹf} �ȱ,�����5�X����PL����l����dzwU]w�0��c)�5i�l=�4��6�[�H�TD�Aݠh5�D���y{eV���3�����ɷ�j/��5�#�mIz^�/3N�a�$��z%KVl١B��wp�-�g�gO_WO,��Rz�x.���i8�h1�Xo@����7���!�wx�a���TBR�� ����U��˴\��!A�Qf}�0#IY{�|�Ԩ�2ņ7�t%M_0�$3�ew����/��/�ר�sg������ׇ��n�ϊ��3 8�&�c�|ލ�J�FϦ�*at8Ar��.���yr�'V��j���
��Z����A�
�0dX֥��yX�z�������Uxi�*����V6��-�^-�)�=�E����F�L���{�O ���i��|����+D�k6r�z�����Ӗ��[��0�j�"!K��xx�����=/�=b<��~�w�ӥ�v�ֆ�}�t�o;޵��4GbM>h��.�Dϕp��4���y�B��C�񚃼'�O����X}*��ߞwd`j{[�_�]H��]HN�����q��9�=�������L�p��Zg����5��R֛WSR��[w�]�F̜j�`��2/:���ׅ9��P�4o�I��<�(m����{��ߔ�`�'Ü���8�X���c��}��^L�R�b���F(�T!���o���釱)'�4�a㸄�Ǒ��4��)�Y��iD��\c�	V1�$����lܜ;M�ANyӥ%�Q>¤tbfrf3+�{�Xm`6���'R`��PtEh�ٻ܆�z������LR��_"D�=ʈ��"��/p���χ�J��&aQ4�$�܂_%��t�W�W�����j�
g�w1Q�r疅6���8���oVo<Ӛ%;V&R2�O��-oJY����B\]�b��ڻ��(tXy&}��s��N��U�"�w�Iy�,$�'������9�z֟*�Y0���h�R$�#��B����\[��)b9���<��ps��>y��O��;;|�j�Jx�k�x��Pؘiio�P���8曅�I��{��G��D.@�oe�OdXN�S�q��d�c_a�̈́?��rͿf�x�g����2Y����Em��iZ��w|��oQۺ̸^�BZF��1�0=d�v�K�<�[�'��v��G�q�U�41�ԏ+�qˠK��e���9	��e�}ɇ���Ls_��wZ�0����l�{I*R/R���}^�izn%Gs>n��z���7�[�����ZJˊ�&c�H�7�j���zϋ
�����գ"�BY�oW|�;�����q���m3�_+�;���咼��&S$�r�lnU��Ռ���"]�[tc淚��K5z
v7ٯ6!�o���C�,;��c\x�`�%w.Zk�&���|�ɕ=��+�*�먴tKp�Ip�KNx���d�g���{)C�f!o{^v�w�o�7�e6��WH!h�,g۶p�U]�9�L�+�.\:�T��d@g4����m���.y��W�eZ~�-�a��y��Xb�6���D�?�倿����Yǹ��+~m�u�٨�D��5�39x&��'�y;�c��E�x�j�m��"������*M=U?6n]��sH���H��H��`����)��e�Yk��P�"��Բ��zy�|(����7Q����d�upE;��I�9'[ս6�|8]!P:|ieOV]gb
mZ/��cQ��X��7x�!�b/7��Gm�܇Q3j���A�L.���(��k���}�zk�1�n��3ͯ'!��yx1,�V�_H�E]�$���D��R��5����;�����n�t�gٙca��Žd4ڮ�xYX��h}��9�G_k|;��Ņ�j�����g�d��M�\�ݼ0��{��냾n(�B���ۖ��&�Qm�D�t��k�x!=����Ih�1RԴ����G�ob��
�	���Oc9ήfu�5�X�'�x��"���d��)i��j�C��n���t�[z�o'��(��.��>֪6��t�n�j�2Q`#ћ�]�p�pO'C��	i��Z�O����f�ܺ���h��3�OSOL�Ųu֧�-[zi�s��e�sƤ�Y������P��C`|�\��jom>��.�����RI?#��W7�֍O]��,��	\�8<C�Gh(�Hy;�[j�;1f3�4�v�v��^�\����ْl�X�H��0P��g^����;du�\����b��"�> <��r
f��ݖ:�2�3��I�q�7�K�[��؃�f����8�72ѧ��r�6e�����e��hRw��1O��v/�BZ��q���)�A��{V.�������ݫ�&f�}��ri���I��ZY9��h��o��Ntz���, �\h�:��x���&���2�%�z�6�
B.��7T�6wgeH�� 8,���+����o\�?�n�%��Ns��f��M&�8�����C�	=�}]Ux��}�����)�nt�yf�+�ä��{���g�X�
n�O���>&z&&umظS��q�i�ms	=6������ڂ��a��`���(e��������'L�2�p�ap��q�e�T�sǡ�c�l��mz���Ɔe������4��bf�"$���ww+��c)�ś,񶥔�]N�v�0�[��u��kL�E���`�L_]�DgqX� �E<k��98��,)�ko�Z����w0��f�m�v���f��ь<�\�mQ������4�
�Wh)�������Hɏ�@�1��`�eݜm�t/���|S6�գ+!�8�[z@��N�.��1�)fŊ�����{t0Ŗq�v�ǎ�f��9ˮ��K���=��[�c�Ӗ	�{4^�D���r�ϳ� �fLF���-Yb5@h#]$����J��ܩ��=���%k�@��m�-�%.�뜹��_'�]�C�E��~��Y/���n��gjo,ʸ��FJ�{L�����^�"B��
F�z����a�_^R�ط�]���nu,҇o[�2��h]i�3t�|�N�
�4{�'���d.띊W:*�؝W�>�*�3�0�客��:��S8ծ�ݘ;2l;�C�^�ָ=vz�殧�$�������g�(�Ub �
�5�1e@��ե
�RڑPej(VT��X5)m��R��R��E�J�EX[dYZ���+ �b�b��A`�R��m+j�T(�h�X�-��E�
�Ub�QKl�J���
±���-�X�*Y�Qb��������E��Rڨ�R����(�,�`�)"�Y�²�X�%Z�Z�`Qa�QaX��AB���B�VTE�,h�,�ŋ"�j�`�b��XTY(ԩm���TUZ-�hT*TX�QV�mE�m�@���
5hVJ���jШ�RQV�����ʋ
���H)X���T�«����(����"ň֢�(�eaҵ�h�ee�l
ʒ��b�Q)J��m
�eJ��`-J�[
'�����}���ށ�}̈�%��W�G{�Q�-2Bf[�e7{8��gK��+U=Yy�Ӷ��t�C���F^��]_d�]S��䈀`;C�:+��EoO6AX+�?-	afn�L�	��Yq��A#�=��~�3W���)ǂֈ��a ���Da �/��u��;��/��*g
�m'Uggv�bi�^���.�w�Kj�
f�R�n�I&c^�&�]J0�2��#�:�������Iw��*�K�T7�ʘ��e/}0Pv��U�t�I5��DxT��.e���r�i��h�,3�`����=� �P�¯�*���I�H���<7�X��L�&g;n��U���A�7a��IL �K���$�:�A�r}��)�j�z������@����6S��3[����xWRn�<%���4��lE7�̬;2t��z=���+ZPJ�֬�f�#�;��3�w�>�m���y��'JKٵnڱ��^��y��5�doПPzXG�v@�ļ)�v{~J��_��/$��{U4��8Wԁ�o�+W��xr�E�p]o�jy���=�}:�g��
��T~���w�����^X���	����w�*[i��Y��v)�!I�ݾP�O����{�T-���,>�tBM2�/{k+��n#h8�'*������h6�x��)�;#��Ho���Yps\]_c�����gcB�XΒ����'���[w���ō#�����ܾ2#����R썎�(1<�>��l��G��H07ù?Z�a����q�}ul�\X<�.%��fe9�`hv!'W�U��T,wf�Y�R��}R"�pOL�f��Z]R�/���}�T1mg}N�(u9cy>���>�&��lz�����p��e��ϫ-'�C��N��)P�,
���4�]�b�<Vsqr��rV��G/�`R�C �;�L�|l;5��&���E�������	u6Tk~�{�g�vR��<l7i����/~�|B��rD��"����@���E�x��,˛�U�2	~k���r���l�*X�C���<׍��<ӓ*E��J�D�Aݠi�&K��V+\�篛(�.���n%3e�<Ғ��Wxg�9Xx��38ށ*Z~���=x���~j��F�bV)y���g�w�$���I��Pn�:Cx����%d�t��Yrv��K�ր���ky��|���ý��/)E��0#bJȃ��C����$�0�x-���h�9}w�Up�dˣ�dx�>��H�h��R��B�as�4�O1�W��;W!x�.|r&t��2,`U�<�_U��!�I��M��3���4o�3�C=�1�T{��$�՞�#�z�	|;�>}|aۤ�"�ю����gW;cW_.�9%9�i|5��>�Taצ�����P��Q�R�ш�k����anp����������BJ鐹ݰ}%&�`o��^֍�M@T��-˹�/zf�+Ӡ�ؽ5��fCk�{*h�5'� G�శP`��+�[�yX�z���վ��rܲ���l��A�鳬�so�>��� p�5�g�� VT�c@�)��01����������g�ZH�/�-u��~2��g�K��=W�ǃҨ�p!�E.�J��rWu��;W���6�����͆��}U�b�<�P�_�S�ǚ���N�/��� Dep�oY��YD�L��
W�ǂ��.�B����֦}UJ�t/�b�1E�Jo���oI��'�a���R���\�g{�k:Su±��xGǥ%��-����$2��A�[�E���K��$�(�B�k�����esO���1��g�t�'It2����t�N�L�V�{����}�.U�p�������FW̲�+��~����M��];m�]kб��ڲz�gH§rkq́f#��('i	�u�p���:�1v�Ә$��R�r��67���d��Ȧw	���\�.���B޸����ׯ��U0���{ܝ�J���c�kN�CB�%���{R����ِ����g�ż�'.q��:��B%�g[�G9s�Tۄn�I�s����ߥ�"úϖ����"��&HR]�~�K������2���lT�qP�$���GO_&�{k#��y�մ�G�L6&&���?q}�
�����z��,G06�p����_^����G�M9�^A��j�u1pߥC��
���HԔ�W�u+2�4�.v��ʞ�+O�%oe�2f�����⢿�ف��]�r��t���t=��}%"�`�\E>�q)�|��s;�yx{L3b�u&������5I����<��j��]����3������틱�_J�o��^�f�3R����o���,m>����h��m�xÄd��By�뽏e���p}6֯�*��`�c}��b��!/Z�&'���?�o${޸/�w���;��K�6��2��20MVg\�Y�ˡ5�L��L�(J�� Y�����ۜ��	Q��ŷ]Ut�H�,eV�,��	cI���'��ߨj�k�	�E�txof%y�\�o����{�����ue�L��a̖�ZÈ���nԜl�7��w\�:���T�O4��
���i��D�7EGfnǱ�Hom
��Z�z#W���M�"�3� �p2�5`�HJ�zW���=���s%�>Eӌ��9�v�5��;�貜��*��~�>���+�Ce�����)r�L� �ce�ufp��#q��ń����d�M����N^	��o��P��`�v<��_x��L��y�=Շ"�����Ϋ=��*��t 4�:&6Y"���h.�W��TjZ�yd�=��ZXO�6J�F��H|�R��'k&Re�`k��;�&��VrN��_o�>���i��'�gW��7E�ߔ5'���Ջ�f
ϫ�?-�,,���Mb����^��N����[:i�N�Y�L�6�]q�-�٢hGJ#e35����?S��!d�b/@�g�zot9]����yB|9Ǜ�f�#/>�:Շ����4�(��T�i�x�R�]�j����N3kugq9�lƶ^_����LB�E-X�(7t�l��g}T�u�����qΚYhf]��ްyL�h�,i��%���Ev�j��T3�X�ti�<[�����w׾[��NfwZH@���ș{�������%0������@���=Y0{�f�;2͆��Pꉱ�JǼ����<iѩ�㐲������(HL��ۺ�2�_h(�"kd�ae�o����Lo4�_
O�^^֫miܫZ�5�p�6��T�z��y����Qn���cn&5�cYW���})l�Ҭa Baf�G�n1�v������V�~�k��S����V�����VX�U��ս���.�+�^@Q3)���֯���;��U��08jy,�g��Vh�|�
���C�:��[֜��E����#�Ǔ�[���4�:�u�]��'�=g����&? ���Ԕ%��g�`��j�X����]�ܚ�{�=�}o��X���X'��w/:��c��4���>KrJŀ��� �uƧ��5�mm隼m��\\E��l������e�s/����Qhpb��=~�'��^+ݛ�&��:)�f駴�P�pj��X=���Nf���C��C�3�������tV�~�0?�B|e#�ӣ�Z],B�=�~&_
�,�����P�X�g;+<�< I'��,Hu`֛��g��<ux�3S�3�T8��(#�4��1O*���9�)�n>� ~�fңF.h1�(wd�F\���8�����O[Sܧ����n_�s�x������w�Na3y���8{�d��"��v��u"�ؗ�_Wz���rɗ�<�4T�Լ9^j���h�AA�,qI�����Ku]{�Ҹ���٧�����7]{ҏ�$&ϩ�A�z�D�A�WX��yB���v_h>��Cj���ײ�mͶ�0��w�j/��4*��k�'���ީ����W5wQ��h��^�
�S�;0����b�~�9�/%Y�&[kqi�$���w=����cX�⸶��}5�l�R�c��ҙ��ki��y��V;�fq��g�F������ڥ�Lj#�r����(א�I�b�c�\%�Բ�gI�ށ+2
��H���!���]�z��"T�e�� Q���9VZ3=Y�;��>�}�Ԟ4,�)u�QT&�o1V#���M5�C��`�C�(w�eه zik��T��W�Lެ6^�΁���I�YYE�܍���^��OQ')Jd+f0p	)5�>w��2��-^�������}K��\�tj���%/�Wz!xC�\@7v{�PA
�m��(����7�����7'��Σ��m4���^(��D�����U��h�BeRs�$� +����պG�tZ��c��l�<�����~��'��ӲM��8,.��\�w�	�.5�1VOT��G�y�^�OLâ�nX�7��ʮ�2��X�B7��v�Ϗj,�ٌĦt$jWg5Uyd��7�5��an"x�]�y���u+ӱ��6�N�ҚMf�{�yйS���qu�`[�xv]�^	}��m��wg���yЃ��k4���/}���ky+̩+TOz"X��l?���2{�2�Cޙ�!��5�b=�޾�[�:W�ެX`3��u�/-�8+C�*�KiN������aÕ�sgA��^�G{<��N��lR���2"�Ǚ���J��bv�/�Whc$�+|�Vm8�P�.F5WH���D��&���
͔b�rf?��i�&�9 |�%�0r�hH���t��^\}��0����/�[�	Sr�;:Ⱥ���qƄj���,�hv2��
�z����"[�<bQ,�k�(W�NͅV�Dv�܂�I�8��	�y���~�X��٫[�����/j�?28� �C����2���n�`���o�:ެ�]��tӗ�[�fIx���p,�lL4M	)h���(?+��|_�<����&�����z��y��	W�A�j��c�1p�P�0T2�G>��J�T#�X!��o�����Uz����ر��9g_R�s�ŕ�,>]�r��t����{I*�JE��8�v��u�|��ͼ�h�W-b�^+�mR�Ma��-%e�Xf0s�(��o���7]t@��-����Ky2���o9�J���:�ez�o�,�Fە�; !,�-DJ�8:��+�X�]�g�f��V���8q���|�J2q�G��BYG�7��<͍A>��c��ҭ[�V��Ul 0uvP
�Ҭ���5�������;�\���]�7���4!�m&S5�ұ5�n��?I��E��Rn0��S��^��
����R����^���Fz�e&iq^S�G�|�2=K�N����bϟ��o�=�U�;-�q��േȉL舜ZF�Ї@ѕ�U�Y�������v!�]j�YQt�7+;\S����Ea��({��O�Yr�����X�ݲ�O������Q���a�������I\D=vYNfE�7�����u��ࡲ���;ǥ>[��S�h�qӏ*��T��M�
�v!&�S39x&�-�?J�������6Ϩ.�޾�o@�pdz�=K`���H�R%�/���4��\ty���NL����T��}��8x�a�l!���.�L����x�iX�C=�N�&�&k{lcS}ĉ���u3����SjZG�.��h(	>!�D{��~���徜&8z�ǝ�o�[Sj�ə��f�B9��k�+���Z>6��5(����x���Z(��~3�����VV�]�y\wx����&��*ڗ�\QU���7���
�{��.���mp��k1�Q�l�Z[�Rib�h9�a7�*���
�xng��,���1\ywh͓�$	����NY�qb��4摍壻Ls:.�{}�dw���MZ��m���u�l����.H�qLP���:ռ�o甁��(�Lơ��Oݛ�_����~�_��<4��ݳ�y~9�Pߓ�Zz)j��A�y�]]�걻�ے[ ���0���ѹ�㡥��Fx���|g�q�u�9�v�K�
�|��jXw���s=����P�&ZHP�i�.30]�-圃<��ޢe�P��*���\=B>�v�+u�[���=��HW�@k�g�gs��[�
+�+���uѓ�@5'z�	�c�C���:q\� i���	��xXB�V�k��>G��.[�g�9�v	��?w��Wj>p���R9���9YG)��=Bia}���L,�'�\/ǎ�4�w�\�����HȆ�5�bv�	Cӭ
ʎV�<�x��_�V镹�i�q[s��V�ش�7=<��=���-��27/��,��L�[��0k�D��X/����/9{{~xsy�Sp���V|)x�<F�TφxT,��İ{-����ka�����:�c�v:]R�.��W:C�7s�}�������p�WMѐQۄ���]�������$�A��w+��";�'x���:ʳP.���N8�&��U�Ptf
��%Q���ռ�4�=:G���]�V��e����&��W��b
b=J��\�O�U�QV{e�F�6���V͑���Xj�Oٔ�;o��b+�kL썈2�UW{]+'�I�/�ݮ��������|�i�39J7��l���WK��7���gv�"�i�s�o0m[Ź'Z�5�o���sn�M,�\��@CM7�h�q�4��*`�kVf����"��*�E
�q ����(�s^t���p+"����Q��2�r�:���]��C_q�vo,�u����+c����r1ҊoH�^��v��a�I��s�(AìVa̶���u�A�~=�C�e�g�ئOvQ=�-ǉ�S���w�o�su\��ӹ�J<�b#����A�7|�	�{zf�%폘ܢ�0�ci=/V�}F�}u�W�5�m�&D:�zV�W��];Ͱ�\�]���u��=R���K����%�Z]�)�g�֘�/t��-�������bb�~�����o��L*a�-�ڹp~�E��5�̑z��]�/������˄�B=�0��u5�`(����q���X��xފ��Ώ��F��ox͑��,A=�¹����[µ�Ŝ��� ���gWf���X]tu7G���iI;.m��8ڜ�����ţ��en��m�C����ı�}����9��xmp���43��2�����.�oL�\_v�`��C�+֕���0���k틯�����l�|{P�>��w�.p�WZ�[��������q�{�톂�.:�Ϗ��{!��A_x����f�t��3�z+�=:B��߮�p:5ս�';FyN�ٙes���jR�}+�P<�UƐ��6�n��ȧ�v;}��N���.wf�1��3	�F��C�o��G-��x���mp������if��_��E{CR����MD�X���y�^-=���Gΰ��N���O��4n*58B�Y��7���٨��Cq��w@���R��ns����&��Z�|�b��VG]|��Ֆ��{���n��N�·�Γk��ڏ�4[�F����p��$vz�%+�bD�9��U%��+_�V�@��R���,�w�`Y�-y���Ǒ^p����Ӿ�±���d�eA�?-�h���,j���5'�+W��r��8ަ)j�fRwg�T 1|� �����cke�܅<+2�î��iN�LG��G9���<��pj3�G�kC�i��85�N��Eu
*���t����>�]lE�\��/��g[�o#+]']��ƀ6p�9e�P��:��t�]92[
�ʺ���jr�.�� ��r�j�e��l��R3��@L@L��	4�3�%-|ŋ	�ѵQ��V�DH�RѲ��ie�@PR)E��m�����U
�Z�*V(5�YK`�������)*��5�X[e�a�
��m�ڲ�kb���aAJ�[kE-��+R(VJ�ª
�X�	D*��*@Ym�T�PPR�(��Zŀ��IR�l�B��+Ea*,�bV��Q��m�*J�aQch6�(��Z�T���eT��KK���Ҩ�k�AT��B�������UT�YXتXʅV,X1��T��ʈ�*���"���""ūhJ��(���J�-����6��J[d(�b�DFB�Zؖ�kZ����ER��lU����m++hR*�ւ�[A*���Q��,X�1�[j��B���!D�TR*�-��~�^_����3�-7w�dn�8���SK}��u�:��!�iu��q6h�VG��T%�uJӌ�eO�j���X�R׽�m���wu��!�Ń����|n��i�U���m
Ok�b�������3r��[���/���Q�+Q��Gy��_���.�`V�a_�ܢ^�co�f�����>��R!>��A�n�/���L��a�6�&��W
������P�c�27���Ŋ3�x�Xjyo��lMw-a��f	�E�4=n�rE��T�������w�6�Yv�<w�ݘ��u1kKc�2����+�o$���q2��ù�w�V�>-,3����̿�m�6T#Zu+c��pD���FI����m�%�+y�c���!�A��J�.������q.�G�&����{+0wO�z���ej�k�Nx7;�JFs�f�D��!wR�V)tR��ś���G�Y��4�Ϡ�ɹ���t�#��8�߾j��CP�ϥC�vaxR:�֫�tyY��Es��{��R8"���~�7)Y�$�s �V$�B�&c$���^�~�>�Z���r=�.}%�ZB��X����T(���ԳQ���]YA�1f�k��_j|;vӗ����
�����uN�vc2�=�ۣg�����Q%���+W�ʚ4��˴a�:n��n�o��~\�.��b*��G�R.Q<
5�\q��"C�˖t�水���|����'�W]vs�Y7���%��Xג߹O+�P]�vc����;��K	�;�Q��Q��n
�B�jE��Ȏ�>2��M�I]=)F5Y�y�qvsw2�����zkC����'�ΰ:�=0h�`�o� ���B{�����ԝ�*j�w6���T�oֱ�$����Zh��,�E��T���ʰȱ�|=�Qm&Fe��*�x=�;��i�]o�枧^�~��@�ہ1�,g�/ ��ĽT2yq�T�9�[�0��|��d8��N\'�<^�hy��dz�ͅ����l�W�]�:�"׎��>~�}�n�Y0c�I�tL�g�(���fS=�z��b�*rڕ�uvi���ͮ�L~���i�J��}3`�r$s�JV}=H������W�Ê��צ;j��2e.]�n�î��x�	y&��\]�;TX�.yhSn���d՜φ�wWr1^�����w�����RӴ�I��`�Kܦ
:X��/]MMOXޭ��.ʣ���U�N�Ԓ�%$�:=(-�fuuw.�8o_B����mvfAdH��������5���.�/�:���
�(J����o6S���"C9�+oNV+�J���2j���+j�tPAoZQn�h|��lJ� v&�LX���oS=��Kj����u����!�9���Ưe3w2Ɇ��D�D��x���(tVׯe���LwHxv)]+��G9��� �*�ʘ�eC�XP�iih���]���A�1��6d�����ˬ��x1I��p]օ�0��r����?�"Ho<2�]O�X�g�N�Ydk2�Zy����7�>��<\P�T���Q#A�����[�}J�����P�t���ʾ�����f���Ko��!}�)� �,F@����S+��^^i�+��~$ȡ�ʰ��;��{+OR�xQ������G���f�^�u�8���5�ҽT
0G��6;	��-Wʋâ[�D�zr~5̨18����l��Y��>�h�J��h{/�q,c�֍	&��aj��dK�{�o&����&p����aP��u^k�D�.�`��P�s]ør^:�`�
���v]���y�]�y�c�k[.ԭ�U������85؄��L����9OW1(B͊�cw<]�ׅE���T�D�@��	�`��9;���: ��ᡰ^��վ/jq��Gh��	�(�on��(��"���j�Rܝ����E���^���[��z}zά(s뱴�t�i��k�|xӷ���,X�qt�ʃ]�d+�w�sI*G�)�J=WR� ڬC?ex����G5��,�G:��]v��E�~0ʛ<5ݬ�j_WE���(�Le
Vx�I�/@G�������Xpt��mL�J�۽N^B�}O��]�}2��T�(	>!�)q���eL�%��bm�y��G�RӧvG�!bo<pL��k�[�G�ݚ&4�:P��Cǯv�Y윩���ߥ����f(��%�w��/�8zm�H�a�Z���u������4r>$v���p�\�n��rq���]��2��<�����������RУ�E-K33��O���|§��7���sE��%uB�.�����R>�L�Y/.�]��tJ�E�)��g7Q��vBl�i!̮:�q���E{ռ�:��~�+g�������=dd5��"�������L����"8풇pb��g�L��nD3_�6/t�F��o^�N;}5lٽ��D�~`��á�h�0j�����k]U�Y���^yo����=d��~ST����/ށ~�oь�~�F�J�.����lx��彼WmD�[� ��1g�k�����'�0������G��'��H���R�3��S\[M(l�=ߏQ1��#t�3X�X��&�����>���������j�[�w 7��v汹�	+�},rY��o�!:��ӷ��/T	Y�{�x���������^���>�R�M�m�=B{V
u��jc%�jQZ��p�^�C�ž�^^���&��m/#��xJ���8���,IvF�wBy��!�d�=is*x�5���KU��R�����P�T��y�P�t�q&=��.f�io�J!�y̳ ��{MJ��p��-�J2<Q^-f��kЧ�T8/"��WT���_��Y�8@����g����yX���أ#C��bH��x��XJ��l��C�-��y�7��9V�a�2K�k� �+p��ה���H<*�#�!l_��7����\�qͺ��I���_�X3ߔ�D�s@����I��e<�x�ӳ�{_�jWO�[�Xv�l�}���<@�����^6ǚsD��3>����UcM[9������4hb�L�˩��P�e��iM�֔V}��pD������]hV��[	��w���)UpoJ�8"k�XHwX.�{A��\㨶��,AY�۷Y�y�k�m���N[��1���Hɉ�k�v������}v��{�\�p�!� m��!w�q�B�H���Jyu�)�giǩuZg�����dƽy���J�@�#��B���J�.��U3��q.�G�&����i{��7b�I�=9�ÍWE�K�����5>F�Q�]#�>q�75{�6/Et�2��h![&ۂ�o���m�ȃ��2�}*X.�/
GO޵T��S��������֣����"�X{�L��V$�B�$�`䔚�u��2�ij���r�+�{u�/���]�)���L��[��ѥf	]� ��e�)А�:J�Y�d��Vfs����� �-�y|��؅�Ԋ�y��)9�3]�Z�UnVҀ.�;�wUk+���ڣ�D����a�Q'�Pь�[������x3'��㬺�6<����z��/��2z��Ȭ*�m�Bc��V��ˉ�
uS)����\���F�is��������pX��=��+-�Ps�������X�υT$�b������{�j�CDpP�7�F(�T!�t�Ë��]�C��b��,�|{Z�R�z��ܶ�\��	Ĭ��}��(xj�X�F�u���c���Ѐȣ���4�*��7�U�VKCB�V�i�c���ʲ�v��|_d̴*�!�ř�u�MQ���Ͻ7o��$f���m:gD�f]�Wu����Ƕh��d�v�w����>@�f���_�Z�*�`�0�jm�d*�b�"�����gނ�r�|�U����솜�q�e���[ o~%�����k)܉D&)�?g߃��g�s�%f��۞|�m��U�3>�46¢4���q/5��ڢ�9s�̨Fl�+>ݧ[Y���S϶s�U痫�Ms4�N������`�Iq��t880��ȋ�}�W�g�l�=�&���}�E��=ѷ%Ưe3v&Y0ؘh�O�=��
sU�U��tKz����H^%�	��S{/<�=�*�T��C��Cs#RRi?c�sΛo�6/d�߉3�Z��"��5����&LDWc��mxc����hК{���-j{$�t���#��T�E]z�Z֞�Y�wKIX.(l.�9�H�r�����8{ݍ܍���tn�V[#�hy���W��%pr֭�߇#!�A�NxƉ����%��*��D�*x�z�L���,t��\���W���m��)1ή<�uȚ�T���7.�L���"=����@�н��'�dEӂ�һ5�gV�	\�yK��|:I���P���cf����"����yT64=�+_.*{ɓ2���1^�x�3
;�f�:y��+7V�ܽ�]�V������nw��w��pE��,���ʎ�Jʋç�nOd�<h)An[���8�~x�����f㚩_���u/��P������;��H!#���{�byU�bf��G��m�ˤ/#{I�-)�__�o]�s]2 �Pq'.��P�s^A���F
c�����:���ng;]�T	3�YN�VS�w8T���BM������~�s΅�uxu���ݱ�'�)�n��Yk��#�W+��Ϫ�f ��|)Ďu"Y���#��v3^]���O�;�Kg�����̐Sk&T6����g�%�*�~�Q�L�����ا:�[jL���������[kz
mKH���<l �4��=�V�X+�����S�Xc�LX��p6�p�\ϻB}���s,]��!�s|K���@�{�D���RU/��D�*_p���<�[6�*9U�Z��?�#A)��m؃ُ����:�jIq�PP_-���L�։y~8�7�IS��)kæw�W���Y�Cфmx"E����w �1�
�ˣ����A�r���8��ik��V!���%����[����;g5�n,�ŊR˦�n�S�۽�	����+�a���,Re�p�w:�8�(���c�M�r�(�5���9�r�z��G��L�7�N�w�]�����Τ}��K˅�Wl�Rr�ɋ���r���zƖqAC�i!\w�댼��W�[�3��|q�w�Q4�$<�N�z�	��y���U�N6i�9��U���C�
�3��[ҷ�W8W���:�&xR����m�������!F⅃bCO�M^�,!X5�}��,�?E*8����{c���郣��}+��t��e'+(�S�T�cO\��+b/���%��.���Ms��,�o�������}��ݷf���\pX��Y=^���V�wV�V?���r��ί�QrC�۵Z)aw�\�sW��v댈�ٕ$���0k�CQ�V��[�um���
f_ap���|]Cd�H�Ί�yyyU��h��/��b�As<�=y�{z7�A�k���Yg�-��"
��CW�x�"��ᏗU����2`�G�;��'U$4�yHL����\��*��#�B�pO}wbeY��S���پٮ�mΗg��z����hG/�&��ʝ������P!'R��ZF��w�)�{.봨xT�i�i-���$�zV�߯*v7���ǐbq��j��G���2j�"磟5~lW�^�J���<�t�C��3ޛ���v��A@��O��k�u"I�9�%�����-L�d�e�S���=�U�>�IX���8�s�k�5[��l��xg�wH��Gֳ��#�LF��r�{�`�Xd\�C�.���v�1���у�#��+�i���y�������iy:���m���la�S4��������Hsn�4"�2y2��L��͗�[�J���m��mT|��M�b~�Vu�
�������
�j�B��B�.���p��mĺ-�ғB���'�������A�5�`~�V`l�׏"�G%C�tH�hGu��>s�o��^����$1{]�{�f�_�ir�'Lؒ� �+�pHj�}.���|޴F.;گϟ��x��3-�.�����������`IH��I��Ϥ��5�	����}���ߦ��w�1���Q\@�G�x���ԧ�5U�]�}�0N
���ĕ�y'�c�F��[�����w��r^�8~�E�t;(��B+NԊ�ב����0���q�yF�o:�]����	���`�Kh�1'�����m?���RL��p�<�ڒ[סbYj��}�dRua�/F4Ѥ�{�z��;���^�܈�V$o0,�њFs섀��f��|j�%�Y�W*6)c��&�ʬBL��罔V!5�Y�$�` n�S���EF�q"�J���ܳV
:6���h�&M�#��.]
+����ݧQ�\�㵡��"��K�a6�{��(����-�Z*ctYM��۳��^�c��~�*��q_��Cʰ�4���0�m�8�r�y�!��W y�=�=J:�S���4]ef��W*>�`�_�������Mr�cљwqڬlU���)w��z�xo�T+�Itv"|�>�����Ӡ�W�^�}�P��=ι���6�Ih�`�]�ڶٙ�f%9�ѥ�Y!�m�XC����'X���z�QVk�ܱs���\��UkX����(ȵ�8m�0"�N���ѩ���=z��/@"u\]A�WNQs�b��vZ���|���m&�J��tM�t;b�j�j⦱өtӳ��XD�j�E>�1 ,j݆B����-v�Ϋ�^�mЍ�/$��]�lݧ�S�-�7�Un-�B7t��s5�ln�[�i�=�M�T(���ՔM�N���(�H�V�ǻ;(m��لav��ۚ�����e�	z�)��u#�DZ!Q�a��X�h����Pa���<  ���wM�v�s�n��e짳s������{��}��x�*���X�w9�3��jØ�nD���:^�׼R���A��S�z���z�SXw���g�83.�n1slO��s�����4�p�;;�S�g�4/5��Y}�EC�����u3Uyk�0(N����u���v,�����a>��Y�wn�u��ŎZN��l��V/!�{��M� V�h��]/���n����������B͗1�0y��=���@���7Ӊ�|��ʅ�fXU}���m9��
r�IQ4�VҲѽ�@Lejc����oo�������p�%��l��%�me&�����8�A��R�t��AlR�Ң���|3ud�j2���v��c�T%�La{�㛼{٣�W}�`�k;�����'��Y�w�^�G�	�Ë��6�Oo��������\��c�FAf[g�Ыa��@3�r��*�,"������f�I=<���w}�T���L�c=��0j��t+(�K>w1՟"'�^�����������uj)�y:�9�c,3��$�ED��6��tF����*��w��NO�P��a`����:����@L[�s
>���!l4�f5$�[F�/iTv���4|{�w�f�L�)F],
�N�La���&IKx���q�8uo�A�8On�ѻ��G�3֯����]�єN��u9���M`,#����[����^[������k��	.B$_@P&���
����J��
�b�"5�k++,@Z*@YF,R(��Y*6�#aF��m��H4��(�
,*)-�D��-���)F)�m���U��AQ��#*%kX6�)R�H���+"�+%�ab"�2,X�k"Ũ�b��*Ek
�+X%�Z�AjV"�+ؠ"���edkA��EEH�
�D�Q`�ƭ*+mkEAh�Ab"�5m
�����@�Kl��XԱV��¤�jQ**���dm%IQb��E*RV��*V���ȱ�T�,R�#l�YR5mH�@F���,�EDPV҈ŭ-�D��T+Ш��hШ�T-ԣ"ŀ��ŬP��J�,X�(+OɁ���,˘�X�(�+J���V`�J��*T[lZʅRՖ�UF� �� �~��D-k^�}��v���`r��o%�k���=�KGk{z�b�Ӟ�1�|�T��j�7����x��MW������S~v�K" W�����9�Lh{�"B��X�W���P���|�]z�.L];$�s�e�86ݚ������R@��cU�8]�Lt�/�^ue����k��{���7.j�-ڬ{BP���|����b�'�oS#gז0�xj��j�ʯZ��"n�{^��n���<�igO�8΢�YP�r��]-���C��*͊���6�d5�����y�W�ʦo�UT3 ��M�u	8�2�(�b)ə��g���q�m�n���m��T����^�f
U��K�^�r$s҄՟OR4?gonls*�j����� �E�ft���TF�K�p6���U�����Qϩ˞Z>Sn��~��o�u���h�9���3���%;V�E���`�^�C��ŗ�PŬdݷ���w���7�����s�JoҬi$�th�.5�)��D�,�}�D����J��w᳝Ԛ,no.�̿6�s�ٛ�e�07��<�ߢ�~X���J���0T2�D��^q���n�)�,L�H鰰�o�GV%Ani��6<�f���${vk|�������0�S�Sàفwp��~cY0��sD���Q]���<���2&���Wa�fUPö7� �"Ӽ����;��RF��e�`��5u}Ͻ{oo/v��2a?�K�J�Ɂ��r<_|t3ɓ��i�mx`t�fW�_���y��`��2e$��^%Khpֶ�b�a'(8`�3
���I'~�gj^9�߫�?�Ĉ��~�~˱�;mw�C�3U��L�f����W����a�L���Ʒ=���� a��Sk��>��:��f���y�:�>���R�]N1f{Bq�)�Zh{ӳx$�hipy����K�\��VXg����z툌�Y�9ݣ����C�NJ;㻗�Z�e1)zߌ�Ŕ����L[l%�H!uH�5����;Tc�@��w5�mZXZS.[9���]1R��8K�����Tאr*��)V�����]M-�L쒵s��3G�T	A�bՀ�� si{�J�u��.���M�~M���u�����,Ϫ���Yj+��M#��^3�P`��H�R%�/��P��C��lN�F�6���2��:<�F�	����-i���N�Ȫ�G���8q5e� ��O�x<��5eW���G��3B�W�j+
���$�ԛkr�J��X���n�����N����!��!,��^��_2�$���'b���h��\���)�ָ<u�ˌEŁa�jS��e���Og�5�6k��`�ٓ/)��Z0s�<,�J=C�򓍆�I���ym6��O��]�	��X�h� �I��+��z� �֔��N)ݜ�H��s��f��Ȑ��Ş�]�Z����# @��3��;	F������,S$�#�hLo'���/�8M�rG��f�#/>�:Շ�͏T��j�΋|�򜡴�ЕNY�r�g�G㸆W{��j��f5���p5�d�1
)����K�{Z��]�z�O�u1{��C$���d����u���,t2��u�$eڒj�[d��C�~Qr�7��S�b��(E|�P}t�#5��u�^]�+ޭ��t�U�J�,�;��S��d��Je������!�����@uQo�Z�K�r5�%�xқ�ꄔn�����ێi�nVf�>���wL	_��a���!�䳪Z�DP�6�XST�F�f);�շ�.��7jG��>�KȽ
�QK�L�NVQ�jz	��}]�!�2�׵ԈUsn�Y�)v�32ܞ]8'��FKL���O��-�z�U{�]k�V�5U�ǀ���S�n!��,a����:�м~rV'',^1n�H�+�v�ׯOp�e��[�����s�h;�w�����w���Ͱ�s�=��S���:e.���n�i����8 �M��Q%�`ΊVV�T�Lv.�duɰ!#'G&:��V^��ƭ�]>�V:��<��G�nmgbo1��dn_	Yz#wb��q>I�"�Tƻȕ��-m�4�<�g��ϟ��X5y+�."����WW"��*�i��79X�Ӈ,�\��/#�:o<�����~�ѯD�<!�"Mȑ�!�'C��^,|�~���񁸩G��n�]�0H+�Y�˧s�;�r�x��<A�[r�C��pBU�}c��S=��ߘb�7���WrD��µܚW��1E�f��S����(wK�xu_���+.�+�����Z����Q��&�;0Q=m��1�b;JL#��1h0������+w���{�PNo%A����]�V�,�Ŕ2��0�S��O.jߋk��w�*@���&akw��|Vl���W�U�
��6hT\��e�P�gm4���Jea�s���-�e�Ӝ�5����fq��. �!�t!�D��5�B��ۄ�<�s��}K8��]Jg�5*N��Wx{�����W���,�EE�܎���{�c�H0��W�ݪ�iu�ܺ���;K�sS�Kfw3�� g@͊mr��?*�H�9cr�]8�ǅ�3sE3E�++8���%t�^�elɻ<d��Y;�fZqq�o[���ݮd�Ŝshghw�y�И��>h�jg�Fs$8{�Wu�k����|c�܋@�I���lIYpմ{������YSق=E�j�W(�m^$�P󵂵�eg*��4b6g�֢��V$�B�39%&�c��
�!)_�����{{]�9kD��uw"E�xp�l�swׅ��:�9����0�u��7���Y�Do�_C����"�V��{KW���,'C7+�3`f��}�בC�j�3D�=j˜v9�yq*|�H���:.ͻHwb}��2R�$��3G�(QJ!�l�t�o�ӳA]��M�.y��G�YI4*�ܰǪ���yU�f
�<�Qs	u3�?j�CH�ҳ|8t2�K��.���z�Ӫ՚�y�N�_L%-G��n�̛��kt�%c�G���6�u��8�ʄ8��s2��'�C�.�#�ۓv�!W�@�z��s�^���E��RX,��/>��M�1����
���V ��W�j��^��/�Vt�g�����q�f��T0�l��>Z����}3'R$v&)=H����5Ua��[������F%z�7���@�˲��3��#�Az'{���f��{�ҷ�3����[l�;��+���::��ow�V�f�z�ț�1H������V*�^78��m�/rᚩt�ME�;��x@ߴ�k��!�h�f�m�\�b��̘�!���§�?R�2��tP��'��>�V��_B�w��myz_+cQ��*)8�6ʺ^�9���_5�f��sD�j��GΩ0��.j �;uC�1^\�Ëz�׭��6�
i�/����v=�i$�w����%3w2ɆYD�t�!��~��֭K-�F��#�Q�x�[S�K�w����W�A�T/� r�.͗��*[��>��eVl�=*���~��WU�u+2�!���Ma��Dļ�u�S�0��G�ň�f��'���o���.3�e$�9H�X*WK���b�S@n�Xs��i ⅄�5���*Q]���� s
�K��}��ϟ�k��[�C�3[����bk:�_C<q�y�1��CV��T�z�Y.~%Z��&���$���T&���/b�}���L�
+����[��G�ۚ��&W�=u�P}��x���%���+v��mE��%�gˏF����ݣo;�����>*
)�k�3�G�k�~�%��L[l$kF�GIb^g]�OO^��jM��vn%]mI��]]��7md[k{�����.�/���څ�C�-�Q���lS/�n*�������<�/�U�'9�=v2\y�r��O[���.��e���i��<X��~}q.�[1bU����iLNE���yc�S�A�1�K@z������e2 ����Nfl�ZV&���>�S�{>�]��g��5�6,#MZ��Uix��x�-�7�*Du�0��t�.^Tc��	nxUݕ{���YG�L��W�'�-Edq���QJ��N$pk"X��ڬ�>z����}u��甫��B'W�T���,�(]1�u'b�L�da��-���;���_>�)��Ĥ��g�>�e��<�:�[f�}K�Ͻ����A���O2�{�ñ�������S띘++�^6Y�ޙ7�8&Wvֆ�����4N���B��Na���ט�}aZ��k�#�j*�����C�������=��z�����azc��S^���y8����=� �H�D�f4�dp�q��35s�f4����4��F�YiY�t/�P�xuI���V4�X�B����x�hn�i]:��]��ްy<�h�Y=��������D�*\������P��@p��ZHSf�+�S�>q��uz�Mp��5���m^Qk��n��v�}x4)���^��rw���[��~8]T�&�`�{�$���h�`Ν�>�Q.m�<���3��g-q+*���n�)l��a�'�l_�U�#�^��X��t���"{8��fkѕ�Ma�7�{d1<��#[X��7�g�����b�o�{j|�f	Xax"�h����p δ�g;	��Ց�ֲLXB��*�O93�t��B=3b踋c�`K]ƨ���B���g�84�~��ml�&�z�Y'�����%�9�>M�^{8�5R{G%��
ߦ@p53���L?l�ak}O���~�P]:�Uf�f^?��,��y�̆xv�b�莸��ƿLd�V�q��6�ǒ�Z,��V�x��^g붝R�c�ܜ%Y���ge���:���a~����J;��ϓW�pVJ�Q9�����;����."�25Z�pTX,��ls�ֹ%-��Inq�� y~39�}�Ga��y���E�'�)f��`��7^��Um��ok���(~x(b`z�2��������G~/o-�WH�>*9�q�/1f xy�KYo�:�mZ(2%H,+sQ-h��L!ΧR�����vL�x���x���nQ��{ݑ�u�|U�"��'��v(�}�2�E<��J&���<Z1�V� ����mdL�(MC��V��g��]gk�ƖEf����\:��hbd;�U��R5bq�x��y��؝�
ٷ���A�5������/Z��ե��8^ij�f�GӵWRh톙�܁Y�gP�n!e�vsD�;�
��fnQe�n$z�k�M:�[�8c��t��/=�Մ�,�.,���;^a��a��ysN�(S�,6]ۙ���~i�h�������!���QrP���Ug_��Ҽ��O��m^1�0&hlCGO4������>�ϙ��!�z?{�m	N��l�� �l�J�s]��3Գ&�b��t���+�=����W�%&���Xoefi�j�.:dW��}be�͛$�t��x'���e��>�����]�4��E�JMf}���+"D9��^�T�Of�\�ܽi��"|4W�r��
�5lf�#���֢��W��W&c$��}���Y�������pp�WF�L�l�}�
�X���l�=����J���a'�DDOM]��fؽ��zK}��VjP�/��� �3�]�I���d#�j�{�=n����Vɼ���Y��+թE��м�ݍ�6�>�݊�a��L�����NYU�����<�>�줠��a�2ܷ8�;�tɽ����@ᱡU5��n�J����z���d�8�2�F��Ȝ��ݻ�:K�V9�݆�_�'�+��iG��+\{x4t7���#m�7�>Ns�w9,�j�w/1(���N��m�\�Q��
��ky{b3�6�o͊F�ř|$z���h��ze��(.� ��:��'fI��^�7����6��>.^&押�a��Gj�f
w1x��щ����h���9�x�z��J�Yχ:��iu-K��u��u�a�}pS�����-'Ί����ǽ)�a���i��V�/��U�`��M��T$�D�W�b�re^�[(_�����Hb��)�O��k��iP�xũ���*��@���%?VW�bh�l#z�qĝ�}y���^���`:d8ЍY~���L48�<q.G�:'<})��=}
r�P�Q�e�v�����k!��W�Rs�MW��9���N�̤}v�x���y�|z���߇���g���r~��%X�,I��.j����d�b`@^��u�����a���z��>��{�{xؚ��Nv�G^��*�ʘ�6\6tT.M�#����v7�LwavR3z�J�S#�Y�����k1qg��rÆ�i�����u~��f��y�U�:��P�+��v�Y%"�(��[L�Ǳz)��k}�-$~�Z�ǖi��\Y%�]��y��>�P�[�\=�2�%9�n[nۧ�[B���j"���]����V:{G��}M�� ��e�fj��?a�e(�J�9������ݳ��7mBy	q
`���"�cr���o��&��nƩH�kfc���{�&���cu�wz��͛���VZ�ͺ���f��#A��W%�z��I�(���(�ʋ��a&<�Lq�1�#�ۭv6w6 ��$]�:!�,�]�Ǵ_)q 3`�vq[1�=�b�v�����}�=E���sp�<�I�Fp��2ܥ��{<��o%�[�X��zT5_7=�Ao�J$��Ϻ�f��S��x�7ں���=�bJХ	������d�d���$g��|s��䦥ˣ���ㄩϬ�)�#YׁŐ�bç�]+�]�~�3��'��e�ٚ)o�[�֣C[����r��Y�[ס���,N^��9�(���-X�'������;�L�@��#줧>: �sD�\�(�8�:kR��2w�v�����
��U, +�`�N��c�y��� �%_k��x�<�6<<��>��X��A�՞k	�%��q%�2�to�"�1�܃3|/t�����Y�Yڂ&-qb޳��Xc�����3�8�2�C;I}c���ui�|�[)�ã�%��.PP�z����0.��S�àE� ��ۚ{�F�ncHF�U��tL��{")�>\v�g72��Ӛ�^��tƭY0N��,Qv��[�Ot=$���]]�d��������p�.�o�.��z�]��x���g}K�F�h��c�Cx��hUڈ��ݮ�v�c�d+V�`��f�!b�]�����ǹmC-�;%�͖�gxe^K&� ���`������w ���>U�;�V��{�1��(`���A�_A�zC�}"�������f���N�l���Q)�z�0-�6�1+r;([�;��:3=�,SEϙm۔-�D�)flXW���֌��^�P� 5M��F�ڜ1�0��ʜ}��K����F��pZ�)&���n3o�hӫ���9�s��0�7��Ehe��r�YS1�	]�%���:B���1N��Z�Gp��oT�����z�{767����ws񆕖��|�6���&���D2�lE֌oC�����'<靇�+i��!�7��A Z�M:�b��;��"3��O\WqΨ9V__l�5B���c�4<�2�����9�|�{�K��G^EB�yt^ӕ��.a!N=G.c.�'wN�<��O�Y�1ݞ�ɥ%�kN�n����eNX��>I������x��f:��I{��wFn��S�u�t g׍�}؋O��"�5�Y�k���4I���f�[C�-���M���
�L��������s��^Q��,�/d�LS7z���\�GT�M���y��~��>��o�<�n|'�4Z#��[D�͵��)�PR�j�U�F��V�U���(�mYiSd�J��-����̹kB�V[k
���"���ʬU��b�QJ���0+c ��ER6��DPУF�DA+Z*�X�X���C��f1V*�`�
����X�"�G�˕�1��Jʂ�X��R*�U��mFEPQIj؈���J�R�F��1q"�("
E�(��֊H���YP�eE-�B�X�Tĕ�(�`�b\�ATX
G(�*"�1��
*�h����I\f*"��0��5D���#,X&$ib�R�2�X�"���C2��VJ�8�*�%b�ج�H��PF�b1#�����e`�Z��*E��ERb%Hb-�FE����F��R�"��X"��͹�������?o���`L����c�N������,�/��N�=��~[o.����q���w=8�t%v҉����9r�3���w�tH�m���]��I&}�M^�ί%^J�,̋���:�2��(�f��^y-���V��U���!L��9C��ʱ0v���j�.X�h��-#�+TP{w3�k1�5����7�{��wF��x�E��,�Cor��uz�m-�_u��˗;���U�}����S�߬z,@t�o��7�r:��n�EP9��L'�����D�R��>���\����^�D�.�3�J������u}�[5QIS�Y��z�پ����-WS*���-��k� Ybz	嘙}\n�=ή|����1���g�e�X��e��8�j����
��b��DM"��cۑoa�w o+���X	��4��\w�1Q��P�}Yk���A����n����0��tʙ=��ҿ{�
0E��o���sly�uN����ɔ�_��6�j�)b�vu������#T���"'��nf
\���3�=2$.o<pL��
e��W-�ܦ ���48��إ�b�![RŰq�T�����*��*`�s��w�P���C7�It]�״�6#�V�[��ڣ��.��L�^��%ӈ�x9��d��g-���L�q���
�!į��+�Cvi��x4�8r�=�5�l9r���w ��ߪz��eqf�q���A�w2yhR�{V���Ǜ�b�]�@����)��;�]m�j<5� dJ%©��
	�C��)��4��y�Fw����ω�lK�y�<;�Է�}��!GR�������u�����`�x6��C܅x{�Y��ށ�jx2g�����BZ�r(D��ǖ�f�+댼�P�Ŋ��WY��;G&wo�kCd�\��ёY�����rCO���;A���A�ڽԥ��HZ[iu�U���O4�F�<��D�S#3��-w���t2Am�TpXc�����eX-�'=RN�-�p�%�ɭ�?&�l]Z��c�ϼభ�d>3S>Y�xe�A��nwR����Ƌ.��τ0�RP_��x^V`�/��V��`:#�"ǜ7N���d��?)M�sx-a�>n�<N�h,Wp��D��?n�k��Krp�Vp>"Uǣ�#a���(���A�牼�)v`��m�N'<��C�s��e�%��GE1¬�O�)n����i�q1R=*Q��M�U��3a,�U�^z���;�=;~K��f��f�T&�����/8�z5
����� )�A3�O�:�@��ˊq>:�@��w���=�|8ib�#a�ޓP�Z��x.�Y�(��P��_^<�@�ǆ�):�T6��ݾ��39�}�;�d�����0VZ0���VV��ɔ�׆Pcog߮�U�|*W�í��k^��N��'���է����e�Ů~�6*��6��[6����K�yxPQsQ-h��L6�N-
W43�AC��d�9��0z�
�}pc�x�XkM��\���ŕU�WU���+9��=(�y�ǉ=�)󺕹Kݞ��M�s��"���ו��X�����f_k�7��\���F�G@#�+�~��4�������$�!�R�%��S�ulL��1x���F� ��N�)L��إ7�wE=3�4Gs4uC�ᾓ3���X6t�Bl�J���w��R��u)8��*���<�R�5��XoD��<ʖ�xȯ��P��Y,����r�j��@��Vy��=�x+�r���椔���y�ȃ���[�ᄧ�{=,�����L���,�M#E��X��}�f�g���QfwL	+��
��`�q��L�E��b��-]����o"��q~8䷕�����H��Q���m�~����l�f'�w T��{&�����"Sz�q>�dQ�:r�I��{o�p��;e@+!��()M굝Ce��Vr��{F`\q����Ӵ�={5���K��6}v�0�:`컇 {KTϺ��p�l�swׅ��:�9�-%��Ǣ�;�۹~f>+�м�0g��5��\���,?!����vQF�!{E=�������z�Lnp��9�~������]�)=��R9���~V<d2��2R���-���rc������R�+�`|����}���n����CuH�k�,��5e��ϔѤON}�O��c�k(r�eX�3�S�==���w1x����y�#�����xYܢ:>����&�_��m���W�\/8P`�΢�YP�ә��=1���T�%lzX�w�W8=hָ�X�?�����>�`|g�-�} s�BM�d+�1w�x��:��fS��^���s6�jx�p��ύ�@��H�WU�����}3gȑ�29~�6���
ۛ½�ᘧ�)���8�B5g`^�a���rLIC=Uf�3{��wD����+�6>��3��3�}�^T#;�I���_5�cw��jZG���"���3�A剪֚[<�A緃�I'�T�~X̓��0m9f�y����l�d	�I��q`���[�ǯZ�\]�v��e.����-/1�o_�ׇK��E�خ�ˍ�|s��F;4������sq���:fz����*NIen��+:ڛ��vL��;i\���]�/ʕv5���n��N��U�"H�0̔�d�S7be������}+�Ӽ�w�&|:R$��x��(8������=�:v#��
����;���J�����r�����<��2�1�o�i�M+L��`�w!��.V�\Y�^L��{+����O<;|�i�J6�3�O+x)�yI*JE��R�����`�/E5�-aѷ���.��W�OT�ל���v�Ϝ�F�c榧uA�m���
j�|/�I��u߀32{�j;Z�O�C���^0�Ot�W9���3&���$�ܡ�j�쥈?-����r�t���r~����w�8�(�sh�L�#��g�Y�O%1��G��t4O)V��A^�	�\����N�v}Y��Y��|����S��~��(�~���<���w���Z��ܯ�ة�[@1!D�u��8z%�d�/%�������qg�Ë>�3��'��o=7�v�zT�.��%~�{��o�{�Z��Ze�N�VS�o����	7��s��L{��,i�m����e3��:���C"�Vtn�y��*���-۰Rwr�̰)	ؾT����%�-�#���u�t��xڙ�Ѫm g����/]4��V�@FΥ��V7�&�j^Q�Y��M�艝y�VQ9���nֻh�_���噾�i�|rS���-�B�.��L���VGMX����_`e�$�C���r������z75# �WD�l�E��`����G�������uB��O5}Eg�������^�p���x���k���m�f���������#��l��/�m뇦w�g�qiڰ/�0R�m.XY�߽2$,	��Y�����vvP��B�w��A����f�(��Wm8��u��K��+�Uo�W/v�&<�.V�	 D�>�j��C���-X�4͇t���D��������������1��5���[����u�Nr�2.k9h�S��KR�^Z��ZI�]��z�z�����^i���b�ͩ�p���W^\/b�g�	BZ�a�x},P�ZHSf�+��q�T��H��(f}b��8d��Z���w�'����FEf�U�NO�D�5��$+���(�)����K:���6�d�:+����ќ(���E�S#0wL	k��������Y�E�N��N�^�\�\�+Hv�$�����Q�8����>� U֘H��CYˀ�g^�Ơ>�Vh�{6B��zLL6t��M�b�X��4�^^]'A�� ���'j���5K��K�����Yjȕ���nFv#WH{�w�17��j-w�|��X�=�� ��Za3�r�~+��gF���K�
���$F����U��l���c�����&>�0�J����f�>�̆xv�b��u��,_n}鲋�]3���鬬�z�C��V�)�xϰ�5Ώ�m5�ǥ�8X�����'ZS��B;�93�3�#��]��Z�0j'3�x��n��,���gE1¬�2�w��fwom��ꮂ��85q�/]38S���#���O;�7�8�zR����^��s���jO���so��܄�e�S0W��XPB�S*����2����u��]5zy���9�K�Ori���p����Wk"���,+\�Jƺ1E�0�l:�Z���Z�a��uӫfy�|<9ə��+q>I�U�`��!]u�V|Yȧ��$��ޢF�S�{ړ����v�r��T�e1Y��t��s�ԋWPL��y��S����np��w�c�G���
�?h������A�C�����6��x(S0����ߗ{�#=�O:����/���A�J</hg�_Vݬ��j��x�Z:�:D`�W��P�oh�ݢ\ Ԓ,cy4:	6���9[wgT;��V1U僽=|�{Z֬������4�Dw�o���(ql�ȷ�p���|�f�����-ׄ����w]|^�eR]�#�mO^�ߝ���k�����B�àA�D�Sܻ6��ۋ3dh��9*���ې��iK,�|:K�w����L\D���	P��Y,�]2y�E�7��gs��
�%��G�u����[������� �+��Hj��Ef�d��|ݾ��V_]Q��H�dv$Y��w�����=֢��Jĕ_{�]y|�+�o#���Ukt���.��Z��FyX.͢����n|�T�����{�y�]"޷�I��tg���K�(���^̃�=��M��j4���X ��!<cE��ɼ�����E�yހw &_h.��V+��a����>�ӣ�fGt�9;Hl�3K�\"��}�Aal�מ�/D����e$`Ыsr��)�V`l�7w��̜"��.��g��<�*�"��l�E�aw0�A����<�����tX�ϣ���@lK�X�JK�	q��M�L�-E�qX�3!��_V/Q�s�"[1��k�����=k�Mh�T|����I�Tm���iBu#�9F�\�;�����I�i+2�ޭ�I'tb 5��k�X=ՙPv�Y�u�4֩�|�l������(j�.��>�t�?�1C1@+;0��_�#y|��\+.��G����\����LRTj�T�Zi����_L&��BM�tL�Y��/�S�۝���ˢ�]��b��+����ԤY�uYyJ���0�9Ҷj�W^o��~W��jF<~�9�Ѝa�A]�&j��O�gĨc;koIdz�]�j>��>B�oΦ�2�>����W5����l��'����
T-j�$�ړ����w�#A�$�nB�v+Z�ө�����*G��=�3%LX�����h߬��ی{��2a�u�I���B�������=�`v�G�J��@���'I�������6�d��68������Y���%&���GR�@nC~-�M[�qg���������wc�9gWc�9ѵ��~N�g@yI*�JE��Qh��c��Þ>-�I
����9w���=�|��t�����l��$h6��a��x;m$��SW�P���o8�[���4�ҵ�2�������&cD�d�0懕b`��}Tpst��j�`!^4�}�%�	.ܚ����A���ҷ�Y��8�]9�2ɋ�;�p�MU���	�ͩ�l�ԝr]\���4�ĭKm]G�X������q��MlT}�V'�	cr�|͵�gi�1�־����%e�7�L�Ĺ.dN��������a�״�zxT���ੜdy{=r����X�j?�t4O��
"���B��ɚ�]���kOAU�D�s~�͈`���Խo�V��)C�e�51�|�����^s�V�E����3JA쫤���xg۶a��H��*�� ��������e8e�������跻���8���lB_޾~��Uy�(l����9�倸� ������w��X�[#�3w���~>$�u�3�r�M��o�ϱp��+-E`�"��KmL/�`��}���Ѫ�\�Wa�b��;�H�L��s�����J3�)W�x�L&/�Vv���q��PR���[�
8Yixb��߽0�bm�5���߇AM�)�{�1���߽�%ĕ�d�B����.�'Ek�Eo�<���ޜL�0p�_�=	���t��m���]qr/�:�J<C�\-=E�(��A.�]h?<��閇iК�ߪ�� ��V]��I�5Ұ)���>�ک��l7��Vj]�[���޸}��;����`IO�!$ I?�!$ I?�BH@�RB���$��BH@�����$�$�	'�!$ I?䄐�$�bB��$�	'IJBH@�x�$�܄��$�B���IO�!$ I?�	!I��IOHIO�����)�ۢT[ z���),�������_���05ρUJRBAT�cgc!�klȚjd��҅)B@�"�t9r�ˍIV�,��u������r�D�FT%��h��J�j�Zkrl( ۖ�����6�m����U5���6f�XH�]�Ҧm#H�
�lIò:-kfض���j�68����l�٥dٛh6�����V��&�H�R��Wn�Qm�`%k%"j�hcfm��1-�       �4�J�4�hFj## �iS��$�J��р  �!�101��&E?�)C L& 	�`L�4d���`F�b0L�`�J$ L��h�&)���D�S�I�z���d�v@C��>�	 C�?�����@��OH�!���A��BH��]c���?�Ț���V�?ڞ���q�(݇� �@��)0 y�1�=u?c �$8����m!RB@!�!��}�<����pq�>�������ƿ7�d�����ВI$Rt�J�Jz� $!;`Bg9���ﾺ㮝$�H�����kK3��O�;7������xgܠ���	<�h=NC"DW����V�������xɊ�El��bеn,9Om�R�c�5�B�G/�)����2�	+��f#��f�Ā�e:��),�ְL�U2u��c�
��{[/�n��i;�b\�&(�`5{�rTBfRT�Z5#�&l͚�B03c�+fJRյ!R���;���S6����,<�`�h���4�S�N��1G vn�ݨ�J��$��eX36��E(Qi^DÎ�B��m-v��Y?[��9�
��f
�{����*��r�@oJ�{�����1aV���L�>�t���n�ck�^�N�۔��{M���in2���N��Ec";��{h�Wi�5���k4��X�"�Ǳl*�Xɲ�]��T�1'��@���.�㽩�Y���c(b֖ņΘħ���!$�8$�nᕻ+&��Ei�s@p<	�pc��Qn����Ӧ�)X��kV0���F��ȶ�%+��@��D~�YqD���,K��ж\)�W�VD���n�Y&�`<œј���W�TZ䧰�R��e
�iϙ_d�����C ?E3KZ�����.S#j�}y�5c����5�,3jLc��p�B���h��A=��D���nڗ�̸��7aإ���f��hEMi�d��:�6���Er�ख���̫̼�T)�XVZ�hF��{����Y�(Ԭ�pFjC&��%Gw\u���֚�B�헧c��K7v���voV�e�*4,���Q��~�B�6��R��z�H�Gi�ɏԆ6�̂l�P�UxB���u0�Ќh²�#�񜠛
������Xĥ�)mC2:EQ�Б9�fMkM&���4mJʕ���(�Ð�<�����5d4�'Wt���ފsjM�ld֯wt&�ѶI`� �u��)P�7$5:@4P����:>�)��3Tk-��:ELH�ۣ�n�ZH\���UM�x�J�X1�Z�3/���wR#]*��Ș��T�@�L0��h�Y� ?�r�l6�!�- ��2�/ ��n
����eh��B�ʊ�����u�^Uzj=@�W���������)��{t���4c)��ƚ�)��V�z.��B^��!"��j�+aW��$uX9�!��o@�W�A�1��]S��t�)�TCIQ��L�r�k)�:��5�]`�?O�O�+=�����=[��S� �Ozz�W�&=4�T��S��a��pf��{}6ppy]c;�<q�K�������8h�s��;#<wG>��u�{9�<�r!��g']]��/���r7X^��b_W!׶%wt!!�����x�x�2��61
�J�kd��a���ht���`8R�f��u��a��������޹�$���zo_3\����E�ӻsv��gJfa�>�݅s���/���S�(ǽ���!�}sO'C�g�4��Lx{���(�D��ػ��wl�i��6�/����	�{d�w�IQr�]".N�*vv����S���8pnvb�<�����t�!L�&�M�儙cBUQ�HH'��.��Vn��u��vj\�EF�$W-=����%��,� ��<��~�_7�Q�z��!�{ҸW�]oCg�W��t�8���U���J����'�as&0��qt1qr�::\����Wf�\���<T�/ z�p�SVWvsr���������e��вL��f��E\��8*�Z1��;�)Wr�C�[�2�>����3;�����Έf>�y:4�j%�^Լ�ں�qU�l]�M�b����K��ۧ2;v^}�79;4ܳ��^�X��9��s/�	�O��\r��1k[�XS�nsEm;2�!t7ϣ]R�,\&=�R��!y���͏ ̳��Y ŖE��X���q�N�b��<]��� ��M ����$Ǣ�'���rA)+RL�'w8Bj�Mq��y�Lf��8�W���2�j��cwYR�}�W­kR���q����xb��z��g�Cad!!X���S�p�ѻ|bc8چ��[����w���LP�W88nu9��nE;k��Xr9ɽOX�aV9	]�f����Yq�Y�a�%6��V�ۈ��B���0���+!��Aߥj,)�d���b�By*�
�"�Qv�k6"�B�8Q�}�1&�q��'t�!!���go�.������ˢ��K�޲m�L�Cz'�/��[w�-0�Y1��Kg'|�b:��Os ]R��צ�<|�w�����ξ�q��-�(8��Q�	\�G�<���;o��Z�v�v�um6�"����\6��ܧ����UZ���Y��n�z��� N}-��M�YD=�}xsD@�⺽S*����ڞ���u�F��{M�UÕ�]'ӗ��X�_P���ڊ6��}n>��v�7��O�������~f�=fo� �	����ֹ��������7��O�����}�:� @!�|�2�����߬�{������=h�$�� ��>n�D�ۭ�I����֊P��:󂹘Ʋq�o]��I�k��n���:Ni�k��r91�fT�V�بp�W*ِ����MZ][��7]s@�:\.�3�+�3@[�7l�K�M�i��n��$��$�4*����$7㒟�*����|T{&v�$���$��f��5����>:����wMJM����f��!&�.���yQ��\�L��ժءY(���/d���Tң�	`����!
\�&f�rM56ìK��(��J��^J�'���.���fZ�EBN�vV�g�6�L� ɇ������͙ɐ��@�X�H�I��uv�,7)a�f��CNJیMiV��mˊ3�(>IM�(��X�Pޠ�V�2��bs�V�'{W�v^��N���9�,�/�U�^�r���Zh�g#{����11�f:�>n�U�f��7��)j�ra����a5��q؆�[4�HصY��	��ݍ�6��P�1Y9Bra�ߎ��	t���k���՛���m
[m[����g�߷'��{���3����\�Q�܊�b ��ѷlc��X��c
tە}�*��y�V
r�\*ʥC�p`��M������T��n��^�A����r��e�[���ѩ���
��[~�;v^
�.������r�|ZDZ�p]E�:(!˲�t����|�i4&�s7��ˌ6G*
y4�S���S��Y��d�r�� ������F�O2m�Z�kk�`���oF��<)�3s�����J��	I[���"��/��[��[�m���]D�Ë:�sy#7�vNye8�&X��C#�IԼ!�W)GJt}a�o^����Z4�ݲӨh�"��COk01F�����YXt���Y�
aj;�nG
��L�,T�����AuYz.ﺑS5F �j
�S�AvЗZ۽�[YwHZ�Iڲlԩ V��ʵ_:mp�~�Ɇ=9��1�`٧t��T-��JN�i
�6�e:c!�`�fZg
X(f��1_:�*4��:��su#�،q�V+����Rm�s�]���:5]������ۊ�ځ ��/��p�]՝�#�^K�R�CI��w����[�5�u��y�o��'�@$21Ed'd(ys�><���'#�9_}S�Nz��N�]|h}�Ec��
��VB&-�ؼ5�cic������g>O�Meαni�ݝ֚1;Z���h�!d�^v�I��.��u^�P�4��V�}o�#Q����M�|���w��E�ۮ���O������V���Ms�UJ��j��\P��h
.F��m��r�s��F��\`��0K�(�,�9�q��*�a��EA�+X�q��iU�	\#��T���b�p���p�"#<�n��Z}�D\���&ͦ)ZË<͘�����ܮ/]�ȵU;�\�P�Vߺr��o��]�}F�S�z���:<��u͋�|���+<���}�{�*Z���B�kQ��a3ׄ͒�y�N�'B�ّ:���ś�Tn�5v��@�&�rJ����u��R�Rk�G���8�s�=ʰ�j�v��&���ՠ�؍��_fx'�θFx,ZS�2����srq��º�k,7�G�{�)V�|�ڞҨ�����T�.\�ڧ�T�R|5������E}{8iЮo��GF��Lv�y������Դ�+��v;ix�mD�B����ϻ��O�K~���}n�Y+�D���?+��U�) 3_럮D7���P0/?-�n#�xO�omv��^/��*a
Tn�H���k0J�GNu�+�*����oC��E3/�@�9��O
�nŶ���M��(����oc.O5�v`@]�X���t]�Nϣ{�r�Qp<O�E_dmZr�P��.�lt��j�l�b�)%r�v-�ۙ�Sx ��*�ٔ����H��
v�Ln���p�9���t��T��܍P�5�5�˫����\/��ōL�T�z��{GW��������䏺�vó}BHm��ޗ�=YytUgE�s�XeD�É�Nt�AHV��b�^D���x�^ݳ��֙oaG�RX>^�U;���V���к��7�U��$�y*�d����l��NT%�#�C ͡��7���Rm8t��%L��ɖe:Ꜽ&��t��x�gWF�"q�5��t�ҳ�8w�5�öm�q����L��.���J�oM}@PG�Y��A�R�6�V;g��Z��r㋥`)9qc��`�5p�=���9���� ]2xy��lA�c�{c�ю�=;��;?+��0�sN:�jn=�I��X��L�I�/l4�������8��[���Xa:rɍ����2�NY��	�v����0�t�3��0=&��2c=u���r���̳Y����YR�i�l�e)��a�l��N�;�[�{��j���
�#��u�j�������'žۜd�P?������]�Uf�VLSh���>b� ��%���8zyM$�T��7=٤��)���0�!�,�2�e�5��p���l��.h����]=kS�M������1��ZG��2�z!��X��9��؟���,��SI�{3�;�p2p�)Y�S��=-�f�ouS`o3]��mo�G��O��,���j��鈣�m�0��R�@�qd��[N�ϰ��J�{{&�1T���:�N�T<T..X���B7i>�c.�E�<>lWq��Kp�.#PӼ7��*�v�A��4�.�S~��P���Ŗ^	�[~�qd_�8�fѬ��H"}�/DDir��a��Ӄ%�����ܠ�էE���G�P[�u=;��z:±ru�BLHN�1���B�'�fw3br������2��M�h;�h}_�AOP��.\h�\4f�T�(�..�1J�WŪ
V#+�4�TÁ[iJ�K���E
$M"P
I) T�S���f�&ΐ���k�xƟ��/�8�c�Y[a��0��Cހ�7�Y�>�1��xX�P�E}@O��*�l5z���ESa����J�|&3��e'6�+4ͧ,Ω֬�44���
�2��7oC�]�G;``�y�z%�A��mx��ISL�)��0k�r�ũ��r!���3���)��:�M�M�۴C iC�%d�k�dBH���v;8�wh !�g���-�ˑ�Ã{CC[��3:i���p,�T8f7Lux��޴r�>��N(�q��x�i6�Ô��0�8��,�6v̳�I1W�Y���T������p停SƩ�hxM�z�ѥ<5ZNӤ�e�t��)]:O���Ӧ��Z������C�4���D�P��!��pC�3!�V5�d<o�z�8xn)��ql�0�a�wz2!b�
c�[&j#�ן����Y����0��s�C�{a�xL�f�H�T�68gI\0�5ަ���i���^s���	�k�5ݚgheznS���lB�[�˶�Cr��gnS�B����Y����I3gHIYĮǛ��'	�.^×��`�4���)ޯ���>b�3;���.��v�6��"t �*k��y�:x|j�dP�f�gx�����r��L0ЊWӻ�0����S�� g���˪a5�0]Y�o=�a�<&�����=�y���g��=�M��V�'��+�}D?0*�$��'hb����!�CҬ�&�a;y{��8k4�:C÷Z��^�s�Q��j�����X.�L��֏�+4�]g���8����Dk��ǎ�7���*=ٔ�w7�a�r��Op���'<c�ݡ��N�f��vu�������e�)6��9���a�g�o�����%�(by�un�5gHH�J�a�D?�`��x�pAΌ<����S�g	sv����i�e�{d�h�&��w��A�#�=�կ�M�'�
Up��ozƦ�4�'��2�81βa�M>;��e�x�ֶ�2��Ҡl�\o���4ì��d���K5�������ͯ1f2(�T�!�5v���+Z�̣�&8�]̷�����6���h�p�!��1��	�
ߞu�6�ib�<3N��Y�]���&�a��DXΆ6+�
���QQ�Hh�!�ڙ�
&�y�w�;�9�/N����]q��<�m�g4���&پi��xCML��x�Y6÷���4�ɞj���+��ƙ7+�賧�Ɵ/K}�G]ůp����<��ǋ��d=!�&XTۨ��^Mq��uN��k����@�[ce�o5���ڟ�����Zm��ۇ:�N��2���8�<'���z흦�d�(��]&]&�����^8�W�o\�P���Í�y���@#�N�=��c�*d_c��@z��]XQ��&l����p��7#�ޞS,����p����s�x�i1���A�{C6�T�[��pmcIs�=����i�������KY�%;3O|�(��0��D0o���P�>��H�i�߶c�gMm���T��qH5�<�����k)�~�K
z���L�u���l��Cޜ�~Ş,����|"��|v����
��ևm&zbٴ6C!����z+�H?�C���{i�kL�M�t��I���,Т8638t�m}�=�i����״�̻���Q�=ȍ�*i�R˜�7������b��m�j2k�W�����w(�WO$��2�@N�.��U��p~b1��"��O��g�i�26��#XξDd)v�wKl���p���G^*8�H�T���ݙ}F\/����tIb6�T� ��{���C��'�p�1{�S�TQS�ei�e�D$`Ұ1�*�o�}��a�-imqZ\%��1� �E���Æ.Z�+[J��3`�����ǚ��u��Y�X]*��
�tʟ= W�*��}�޹�x݈�x��{5�&�����lӴ�}{C�a	��y�8@:a�I�Z
�����;�N���Sl��!�!��J�$9ޮ	'd�L�+$2�C��B}����:ʌoƽ�uݶ�.q^��.s����gj��y�d"�I%@<b�t���A`M$��$+��I<2e��2�@0�RC	,4��;�@�a�	0��$;I
�i��Hm$u�Hot��	�I<0�He'�!0��o:�|u i�I2�2���$���z�RC��sd��!���I&Xe�9@�v�n㞞w �'�Hv���l�aᄚa���y�9��8d��	�0�9d�(v�6�����a<$�ô�G��4��;7Aƥ�t�cc�ń֔�_�6�K�E9 g�0]�5�bX��4�_�f�@�6�to�P����I��AP�e����E�K�c�L=���S��4�v�oϴ�>�|�4�����Lt��É%D�b��UA�\4X���5�Cg<�A�
�v�l��xe��]$jX��t�Ș�pQ�V���4r��K���)�b��,�{+v�_�;�mj�^u�@�)57#y�:>��-W�:�����j���1��z���&]�֪�] �45~n^_7z�$l{�E��$����)��_V��|ϟ>��։��u1*�Dm�a�C,��¡��n��Jt]2̜z�^>]}������4ie��$����X�y6=h,q+^�z}xA�΁�^�w|g�u��(���z:�m���f�S�6��R�%u��\����+g�� N��ʶ���=��TÊ�s��,�S9$#������U���ZгL}�m��35־��>y�ξ4�b��)�.�>7;f�KV;�i�~m�@��z�BVf�u���ܪ�G�n�S�_?~l�
���C,�>TH�`�vR��u�*�^pRV����Y�S'����/:k`���ģ*�2�6Q	x���u���(�:�{ɣY'��qg�x.�S>Z��2��u�b�4}�)(S���w��Ll���Z�������8\"�b_=ګ.�b_>��S����9#�4�mXԒ�nצ b�?j��0�}�G�s��vy���/2N;AM0D%*���2A�<�a�7���������$E^?�ӯ������#]zE���m��t�"y�i]�-Y��P��.�y�3���epT�;8Z�-*��43���'Yz�#u��Y�"@fw�m��-!]G�u	��Vډh�-l�Ȅ��+]���j�w)w'�T���yi�]ⷍ�K[c���j'n�4�DZP�q6��If�e7�)��V��ܜ���&R�u;9������o�E������Oh�k�$䑙;�J��ǜm�h��E;]�����gx�w������yy�oe�mkQ�R�QaKmb%�PeKj��[kKiYK[V����h�l���[k�\1hVҭiKh�J5���p��!�38k����f��	e�*���Y���k)L�8��-�:2�w�ǈ���1�_ ���φf"�f���
J�G�7�mٸ�_�z*>���ѩ/ܩt�-�GG32I�(�H���s`fR�:f*� w�>��csbጙ��^���h��^u�Fy��U ��;��avt��W�@4���<;*y�HXM���We�ْJ�vF*8�\ʗ,(2�����ۢ�E�����qM�Zp���^��[�f�7">���o��b[I���
��$,Z�۞`�����D:��{
����c��+��.>��Z�]B�%�Ǽ��1�Net��xqn�	��ÙR����N��85����h\S�Gֶ`��D��*�j�/�E�u{f��<�BZ�>E�ީ�wt��j����K&��u����q��@&*8z��V�S<��L���Ok�<�;ծ�e{}�H\�_B9�k����g��u����Eć�*�|�f��44�K-�"Z('w��ki�$K��t*rA}��/��xe�􎶽�����}&y��
�n{L��U���+�J�D=:u���C�oM�b:h����}��>��u��!]Ƅ�u/`p�5�o��.S�����6{S��Z+�0]�g�2��2fz����c�X�x�v��.ܾ7c�̋(Չ�����C�q�#TfD�ՙ�Y��%e��b�Ŀ#Y����]�j�mm����u%{�ﳋ*)J�G��r�O�Z��&�wqW�F��Ze�]+0�@J� ������]v|>�9P:��pє�Yu�r��fK+���p����/�7q󓽴�Kɋ����4�l�V��#s����*���{w �Ae�k��]+�/3��{�g�r��LU���a+ez��ď��*|�p��3�)��UU;`��O��'��=x��`�8��Eu�����-���T���1ۂF_bݣk�����-�Jr��Ѳ�UtO���n��x�4Նwq�hY/	�����tɆ��0$���aV�W̷��#c��}Q�����Z�M�f�ȧ�A�ܗ��/_]�`\�VV�9ڐrי.Sr����*O�Vc,魊r}Z<G(k�*�:3�c�K�r�WQ���p�K�7�w�?-7q�,��xΞ��q��x�us9;���S8��j�J�_8�;ӥH�h͘�FKu�5�l�-%%��g0��o	�\�S30n1դ1�s'O/���N���Xm͵���+EE�*� ����x5�c�;�YG.ε�9�~���[�����U�uP1Ͱ��#"L�<��D��{��p���}��u�wFS�����p�~9j`�!lj�����2*:.r.��B2DY�E��\��$�6��k,��͆9��3�L �����	��փ���W�+��yM�.�rF����6��R�<4`��m0�ֲ.%������wB�e͋�e�J�n`�ɲs	�رf/��k7P]�OՋ�r�rG�dT���%y���|�w;Z*�թ��y�O,�u��K^��m��V	����b����nn�w��,�^-��,��N&���9�;���ߐ�����#��ϳ��t]t{Idgg����ͮ=�s�e��s�}Qs�h�W�Z��L�XL���r�Ì"�;:$�v�{Y�y�X�{K1*9%"�J8��o7�k[��[��'��a��l�GU����Mr�B�=f{/1۫��V;�ki�+/Y�J�{V��3�qa}c���'~B�U��>�߹FZ���=��_3{���}��3�hH/0Aw�b�Ё����ڎc�����RW>r���';I/LR����m��I������������~�u�^�\Y��{(��I��"������ڢ�:8��X�� ��r*5�H��l/��md����*�Af?��U����J�v:�Q�j$j.SH�.�o"(��ύ��ѳȇBKe�&h�a%^_HI#��3{�M�[lU-�i?�w)Lf~��(jA�.�v 2�n���=�&>���8�Dm:�̇�kS� ���	��wK,d�/΁ɵ��״�I��gH�|�b��U}��e���l���q�����������9r�:/'k��H;�75e �*`�j� FAYW[0A�4��=���O�&7'��驵�3�T�X]$����x��]��A�f�Ӂ�2�H���2`��A�To\�qm�k#0�Jp����f���q�5m��i
]|�׸��Si� 8�J�ڱ��*��ꂒ��i�kb��-`{�i���gV*Ћ,u=��x��D	T(�F(�B�-"FJi��H;`!d'#�Fײ�U�L處��N�M�G[�}�Rr>�\ ��h�JCeĪ�~]�_�i�^��qQ�����5���X�}��t�}K���h\��z�7�O���@�wGW�%T����Íd*��[)�G�Nի�f�9/7��v��G���5��`���9z��áz�  �C�	5Cmm�-�KkEH�*���+mBڈ�k`�V���ҥ*��j����5�mQ���PYF�����9��全v����_��{�rtD��;�w�~��L�0v.�<�~�j	�ה��C
x:\'db�g;�{t�:���[��5yxL~9+k#�4��[��E�+ݫ(������y���^�u�j����撉�:f.�M;]�W�i�m���lE�T��g��ENʏr^����Wyw�X�ym���lS�g7&7~�{$�IdBH��fffrh�P�&т5\	lRџd��6Pڝ|3�g��T���rg�j?o�H��fC�M�i]�=X��H�~���]�^���� όl�Ci�����4�;�N����0u����u��Fm�v��k3LK��3\ၽҖn�b��[��𕸲��t<8]��^r^7݅�w��ᾡ<G�L+�jՍC�<��}p�m)&l�D�_7��n~/�]��\S
ynK�lYZ<�rr*B`�g�3/|���Z�w�z�liF����e���00>~�,�x�h��fj*��z��L��d���_y��z�V����}t-0j��+���8�b�j����8@���u͎�V�O=�+v�2/s��B��,yE��R�����`�'ވ"%����AB�*����F�/���7��g���`����7����GVt�qU�����ّu�+��D'lSu�R����S֍� �����K(cM
�2����֙)DtǪRW�*1��ȼ�)e�E,_{�oy��l���O<7L'��Y��/�6��
�A̙5�W������*-�ѩ�7Im��ѻ�ӌ<V9��2����R�;��_r�Rg.N8S�Ief/���f&��F��Q3��o^�v�Pٿ]���8fQ���I���~�s�1%�B/��u]�M��I/�T�2����eC�4�:�AUD�$��+�������Q�3�Ϙ���c��vV+�_HflE*����2�����aŇr�j�J�J��v|�g�ҏ�ZY�����9w�?��0}b��{��u!�%�oF�eJYDH�<�����F�P�,�Kާv�7�3�Y�pgj�ɗ]���[���z��0�%�����@cv���O
��އ��ˏ�VPe�]P���o�dO�	�H��}��;'�$��J����N�Œe��I@��h�w#n��v6�_gq
��E�$�
�(���FZ�{P�y�ow/j�]%�Ŋ͹/��q9�˳�g'p�IդΝ���&�����`���)v�ʹ���Rx��h��le��[J�kK+-����Z
,�DE-)m�d[-���(��UQKmKZUT��e�mh�*�Q-h�[Ub!mmiDh��EmZ"ֵ��Z�V��%T��-eJRҵ-���kl/|�f#�I;xc[G���30�9�@�W�o~�r)��&�6h��d��|�-I�����/�67o$�Ư3^?�b~7>�>�����#~p�-�=�v�E�V�����H�}�Y�X�����^f/�����~Oq1�"�޶6(U�dM;cׯOMV��h�T)^�nbr�-L�Kh� t�ۅe{�N��n%��
�q�$+܍B�{*�)V}��qs_s��I%���cU�|}ɍ�wU:2"�T�f]�;�o5B�9S���Ӻ}@���>��H��.o���F�&�(���NL��ӡ$8_S,P��d���h�Z��SZW����311u+x��� ,7�[�z��P�J	y����k�c�_z�z���$����{v��v遺hh�����*_7�e��"�i޲�DٴBD���f�mt�?�y�	�O�s��lWU�9��o�)"1\�C�B�F�0�,5�e�L�qUX�����*"�++ �����6�p���R�d�RŘ�fo17_NL<��.G8y�X��~_d2�;��˸E��,������p>/}�v��������Q$3���,;��U"a�.��45��L�O��qCrt��I%�p�����-m�y��//wo����+bf*/ٰ6i(��hU�f�K�H�gzRA�
(EV�lѽT����F��P̉�p�����G�{i}[+�F��A�M��Ҕ�/��ox���z�~�~�S�M#t\�H~��p���$
ϑ�"�ܯ��^��i�D?ų�q/Ү����vT�
f��6�X��x��<�Mp���쫇��:f��YR1Nf/��f���޾����:8d���̠�*)P�+꺔����'w�W�R��YkZ��[[b�'i�Ns��A��!�ۿn���D�̸�cg�^v
��r�|wp���$�LR4�/����[�����1�w/����>;=��A�b� S�^�n�$�������n9��K��r��"��,k�e�tD�N߻�d���f,�� ������򍣨:��=�y�LK������W�ᩱ^��tt7MQ�n�p�3���'��Pt�,8�{��2Lφ*U���;��(��5]�B+�N@'�"i�b=��D�B�k�>�/�`<�٠��JG��̵�/B.jjd�0W�e�բ�~M���?gxv��̎L"�h�Y9`��̽�;�+�r�%��-ul޾���M���7��ǹn�wo��r�,�CK݃^ҕ}�iU���� �(�h-�Z�-D��m�D���բʭ�Kkkb���V[j-���J*����*�JնE����U�EҊ������h-T������Zآ�ƥ*���h����*�*�?~��s3�fN�j<�I~<�fbh?�S3s���J��E��m�jу���Rei�*.T�u�����51��޺x�+����*b�g��^��gZYV�fqO��{}u�y~?/�����a�	��
��I6H�|�,�����Wq�S�b��lɗ/���Y��+�p��S�����/���q%jXn�+�ه��9v/�n ���R%��aɚ�r)������Ma*�r	�ߎo7y�ˇqG;[�(�J�%��Y�Y���$\P�*�ܨ��WwI�`�ϣ;
Zj���ˑ��n
ыz��^m顔��W'��?���m��]�N��-Wi��PL�5}$��T�Tq/��N��%�.9��\�_q�������Z���ʕ�m�6~���hQ<��q\yS؎�c=|��H�,�Ζ�2��AuyZ��XS4�.�泱2��{�^�<d��O��5Ͼ[�|;��R7!vORlC*M���ع��zIc�6w2�!��A�l���)�v1�`��#RSLv� ��oF��L�^�'�7n�"-�K�=�G�����'NK]z�ێ��\�K-��+�?�+|��}�y�k�k3��e�N��Cu�$����W�v%ąv�ZԊ�{u�joO?GZ?&��s=Gjf|�̻�^�iw5�D�[�NH!�;�,s�%����6gu�Dd��3I��ҙ�Ѿ��"=Z������=��Lq�����[�<����ãPXGY�xDP�L_�=�����i��6�E�ݭ�}O���n��P�%ר�~p��U%���ka��ʅg`���g1IX�	j��O�f�^��;����ٻ/ gg`~�X�cp�{�zXO�x�}�t���:�-�t�[�ީ�t�z��&e�+�i ���2��B�4�!Q��G�;��6Yn������x [�:ǡ�=�Pxr5A��]�!�z�zz�k�4�!�z���l-��):�H�d�l��J'k&âнv�鍘��w�ו�f�K�GRd��;�Q�a��J���� Z���'�Hy���~:�I@jZ�^�Dԍ����ή�\1�5�+jY7��A'�9cbe�:je��ի��։J���+zh�<���FnL�J����{0Q�G�Z��z$ް�H{��ᛮD��}�0�k#������]7.ja����nS�6�E��)'rbbH��Lxy��b�׊��VK�nu����N9;�&x�b��Jp�nb͢���ե��_&OwA+�j�f���|F{l��Õ��X����;	�:�EC��ή&W
"�Q�G�UX�(��8�`�LZ��Ĩ�l\`�Q-J�hءZ�ѸJ��n0TLP��m)FU+[�qYKh��m��c,���01�V��b8���cl���D��!�����q�>�e(�մr�G!M��܇���s��M �!)�s_����2�/���Ud�Q/[+tRC0�x�=�bO�����;|�mp�KW%���vlX�(y�w\5t�V+�rN��\q7Ի���w.�h�yr{:�/G�]ؽ�w���V�Ά�j���a3VR��yey��Ǖj������^*x�B/$�[�e@N�T��ծ/ן����!��ϵ�ש�'�rېyg��̡3��;��y̙R�е�Hכ�V�=
�M�۷��sb���k$�kke�T���Q��d����k��`����'�<�fCE ��d�+	�ذ��h����b���I�x�{�&n���|dyl��Э������aسp�)�g�׽!-����E-���
���*�e,M3b ݒ�w��8�8�窯�p����w��9���KS�{2��7�3ub�)U�R{M�S@Kw�hOu���V������t�a�9~Û��e�C�N��\T��ۻ��k���ϳ{�%�Z����%���`A8%��m�g��U���Ò_����l�٣���� �K4E7wr�@完"z���G����:�V[��3s s�ʽ��&��tS�X�|~�����>/8���ܴ��-e��z��Ja�K�'�E{{�����L�Ɲ��5�.E�=��K{��������Z3�ɪtյV�7FwTI���V���]�Y繣��yeܒ\���̄�[6;�.�:�U�C3%��!��ma�wμ��{j麻�恇��cU���v̖�b�c�KxU�ڇ�:k��wGݭ�K�����N����C>��G�y4����f��/���K�RGu�;�	�ϒ^.b2� �D��I/X�*a�����,~cѫz�+�N�a�m䑦��8�����Y�=�f�)]ǵ\u?&��vL�^���%����\7�9#��̌�9�%t�yo�\kJY����W�O��7���QB����y	��Y+7�KPޗ��s���gI����8G���Ӳ�=�k1!}ʀ��P�����$�(n]ˠ���s	�T��z�w�:�}����p�ɚs�X3x<��c�⎭>�q5�d;j#l[jͣ��2��/�G�27)�bod���MD]�D���x��@o���vr�uf�_�U�D��mݫ��P�j���!��}�|����ݲ�L��Z�W��g<dz�+��DU��0�
�q�ch���Bв���1Lb�"��*ն�\"%�G-��YmKT������p�ŵG
��h�c%-p��c#����3����Y8f�!$��v5Κ.���ث�~I}k�)A��ܞ�1���yKӠ�is7�DT��k�Ɯ���n��cݶM@ߛ8����"�͵j1MS@D�ӛ�f�VJ���J�wy�9�K\��b��9�-�*W��8ai�+z���r�f����{&W�����޲���\ZY��5=a��;H����7S�C)�CN]4�eD���;�f�R�g�TX���AG�wQ�,�hv�s{����S�dto�~�u��P��*���V��\}��܇ѿ/3t=��R/x<)�ȱ�����{��v�����o��� �����*R��Nպ��ד��,wZua��ކ��+���Y��`7�����ᗕ+#Z���,�-����*���S�IO��D�$�����M�Nz�m�4|��e����"j��o��]\k� �*��u�t$1��6K#������{�l�o�()wE���}·lT�ld씔�6Q	Z8��=�jZn�!z�vl�����8�8;gɠ��^)G}�ۖ��q����t���f�ͩ�Ь�N�����^Xu/\�+������nD��\�
$t���y44�mN^��T<��p`c�v���R�t��ߚ/W���dK�ZCx��j�>��J�����J 봟MVx��;�Oמ� Q��ܺ�X],��A�y��x��L��`�¢����U�?�,p�C0�$�[�.�VV���p���N��r{R��%���̑��[B�<���&	5����9w>�IS1a�83�%�Q�Yj����W���ږ5iK�;3�3�g�U�]]˒�i!7����,�Z<�P$����WMŸ�ƭ<����qR��'1�^��{&�����O'�$�QR����lV�j�o��ʳ�|����h���n��L*��Rr�]4����R�jU�Z�2���������[�Z
�~��j'��Z��W�����I$ ����Rw$��l?�`��x����Y�!��lrA�Gw􇡙�ъMl�of��&qB��-,�8b��[am���u� �y3	C;,� ��HE�Q�S6�*�J�e,V�H�ŋb�X�X
�a,��D�!|��A
"L�Qo�^)%&�d�[��c�@���Z���f����y�߾<f?ȅ�}���h<�K7&��ϸ����cE���>'�|Ö�s8Lh�̥�<���x8`�!H���h7�q�P�@���C��}�Sេ����$���=�@�C��'k�@d�a0O���=.� O��`�?�'��@�ƀ��?�������zϟ���>!���4�}�� C��I��p�����0F y>	�A��!�d���NhHs1	OW/�ht�#��`��?O��c'FX�4fKv`� ��g�����!���|�ɸ&�0����'��I  ���x�5ق�%~�;4$�Xj @ �:�.�9��H.�,Bd��NY�����3$=f�y�'�2y��H0,
���H*�T�m������������<��z�r}��j�3��E��{C�<����@�H@ԓՃ�q'�3�A�?l���m���C�g��"K4}rPш�_����!�H|~�����!O֞�߮��?nd2wd��>E>Ϥ��Ow��6Oq6|ć��^���=A�� �'���?@s��>2@�$�yL�~��D@H��=��D���z�GA��0"~Д?�$(2��i� �L�?�|��a��YrX���������h�����q��?x H6M��D<�p���rQ7XH!da4Y4Oǐ=�{OprI�8�Ǆg�6`�[H����'2I��!8JCPfY��d�J6��d�Nb�sa�:7$	R���,!�>����o�$]�ω'��!��>��C�����G���'�Y����4��������g�C!!�? |$�3@��"��4(Oy�8x>L>��=L$��!�R����= �?q��$|�{to�{_i"� ��l���~�A��$XO����s0�?���� �A��<�!�=�&B�}�vC���!���~��dpI��OO͐����< }g��y1�����:�h�}��=˿�������0vd�E}2�� H��O�ql��i�=(d=,���Їπ�?w�<�אOQ�)<��L`���l�����<�3��0x?�xH{FH�F��O����<wBC�'�>���N��'��$=�}��>�=�I�4��>?M��� �����q����c8���b}�,!���A~_3Вy}���w$S�	���