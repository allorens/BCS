BZh91AY&SY	��_�`q���#� ����  bB^�    }T }j��0hf�-h֤U�4IF�2�F��EJ�m�P��Z��ڛkV��l�Cc)�m��ֈ�i�CF�[5�FJV���i�I��Z��Q��#E�b�Zٵl�����
d�*ɚM��ٶ٫e�l�ʔJ
�[$�6V�QF,�jm[j��r�bkH�Ҷ��V�RTEJ��bd+V�L�,�ͥ*j�T�m��[m�ɕm2��Z�b�Ֆ�SX����6ũ���Kq3�a�T�[�P  �or����3��u��]���l)�4*��Z˝j�4�� ZŸ�;�7a�j�ӈ!��Q+e���㛹F��"�-�u!�+Y�  ��/�[�SM�yw��M5[[���w�����mq��R�K�O\�e�v�u���/xRm�+ݽ�sxz���M�j�-��z�5�����m��ey�w�Bm������V�f-Ul֒3eE�  [����&�>yYҕOV�6�޼�m�v�m�y�6�V�늓93�
^��\���u�m�;����ٽwU4����G��n��.�]�J��oK����Q���M&խe��`)�M�M�  8��顶���<{��V�IZ�ʷ{wqT�S�����}v�کu��[�R�]w*��=�um��Y�Q��W�eVl��ꊡ]=-}����}�2��	Ӑ��◽��ŵ�BBQ�j��J��  �d���֊��������Yw�_q��޹��N����O�%������U^�����&���j6׶����R��zU9O<9���Wm����S���M���t��-��}�\�cl�U[hͳkmVډl|   M������\���Ҩb���g�u���l���s�=�(m�����j�m7�a�^NvWl潝�4�Km���kЁGz�����v�t��^��s�m���J�-�٭[3lZ�f�   m<���}���WL�^��{]��d�Z���[����GЫv�Zp=��%M3gV�{�r�{v�^�g��)���=�E������ֵ+Ve��ֱ
�	6Q��   Mޡ��z;��4�D���cѺ�w����u{��7]�ޔP+=�{�f�c���Y��޵\�`�u�l�L�ȭ��l�mc)�  ��M�+��8�C�{��Z��=�=]��׏x�5��]�8覵F�a�:����C��[��
7�=�m�-��[l�"V�i#jھ  ���֦�/�8���G�tPG��נ;ʱ�GGN�<�z{a���@���t�A�w��A��竜�����  �  50T�Qi F�L	�A�)�4b��I�   h4 E=��*       ��$�J� �CF&4Ɉ���UT4�@     ��D&"��$̚��4�6G�~/����@�5�P9�V�~C3ӝ�K��yvOOvG��|������������Q w|y�_d?TW�"�
��p'��������S�� ���U"�
�L!*d����_�����~����d9��0?���d{�������>�	��#����d}0>�_L����}1�̯�G�����d}0>�L'��_L�0>�L����=2��C�#������`}0>�L��G�)������dL��"za`@<g�"��� zd@=0 �@�D���D�/7�C� �� �«� �� zeU�`�� za0(zd@=0"�a =0
�` =2*�` =0*�0*�dT�W�
��C�*�� �� zȏW�ȫ�d�0���>�� �dU�0�fC�� }�AL '�@�D}2���@S�*(x��	�P���z`D=2��UL�'�UC� 	�_�L �A�	���(za=2�s*��POL '�� 	��Ȁ�d>X=2(L��C� 	��ʂze=2(��~=0���@OL�'�"��P�����>�� }2�L�����L!���0���2'�@���_L!�>�TB�aL�=2������=2��U�ʇ�م�`=2{�>쏻���2��_L/�G��za}2��_L��������4�Ͽ���������g���P�^��S�Xplg�^����*�!w	���<ZK�N��۹[n	�W��P)�a-wQ �7���O�# f��F^�z#/sL�ʋ^'!�ݘ1�٠R+k-�[_���$���	d]�q���Ƴo�>�J�6�ͳ�4�}uRZ T�)���a�Z�䠫$Ì/�Y�-��z0Ի���٥f㛛f�:va�	9�.bh���B��VVmƃ2l�c�[j�[Vt�5�D<<��	O���
X�MT.n�����ͅ��!�Oa5u�)�gDJȔ�r���M)uulB���X�����(0�t
$3{X���[��)���VI��9Em ��]�5�Lƀk/M���tMq���$Ь[��ƴ�&�ZDт��=2�8D�M�����ٍ"��m�D�%��C��ɬڠ⬟��c��y�,��*�a�ս46hVk%lu�ֲN܈#����(��H`����yu�9���u*�6\�(�5���,�)Y �@z���3"��<�� ��[�ݤ�I+�`�42�
C3����ַ uj�u2���쵀㎣���K��Ķh5�jT݃�9��Zuª�t�*�^;���KF�,l��U�ݔ��X�K@�]e�4f4l��\���O�b��Z͕�����j�٢A�bX�P6���ԯ�����S��^�:ږt�h��7�Ve�X$wZ��[HT�\酬SV�AW)��BL�)��/,�/ub�fX��,���TU�$��Lt����y)�(��S�']Md�ݽ)Z[irĚ�p�a5)f��] �^`�q1x����630��u�y�����Y,"������;Lԧ���ːE��66�Nչ��M%fLƊ����ե�5ch����\l ����y�K��-��(p;ܗ�*���R�G�#��`�@[�i']�`�ܲ��n\D�0#�����v��7V���Tr��5�f���"�w p�ӻ��٣����]br�A�L7��T�x���l=7�Xz7���b�&�R�+u\+�Q�1;�L�����#ɔ��0����!�t����f�^"�i*�}ɰh_<�����f����v��"*#�ml���v4�^��M�0:'S4�>�n�ph��x�W3-��mԬ�r�n2����ݬ/r"Ty��&��*՗NUc�ycu������r^i*���5e�L3���a�f�b	X`�:�\�-�c*j�yc�zh`��3դ�;ᖗ&Յ��9�ٍ�۰�-�6Wz	؊���[�WM�#�5NH�;$�z��J�,f��m�eo�+�����v0��x���t���́a�ɷ����M浄X���Ӧ,�)�^�$�n��.� oV�T]cuL������-c=���U+̙
̹zd�,2]��E�5!�Km�3����ї�m��"�CN�.R�t핣I{YO7kRT�/\�v#���b�0�Ʀd���&`�`�5ٖ��ꋇ(b��o-���xH�a���y5ZWi��F��!Z�E�41��P�Z���2�T��b�찾�f @l��#)]M���IS/,:��f��&�ù��/A�U�O�LX�r��`t��l5��C���;�vy1A��l�$6�(.�
�fc�$�f���8z�(F�.��*bNa�	4��ƈTS���6YZ�����r7 m���XaV�i��Q���ݥ�6/��-Tw�a-�GF;h#v`oQo`yq�+t���`8I����n�oX<C!�e�W<
�`$r�������+HU��C�f<EAl:����r��D�׻��bS�\��Vn&n-Р��L E�&�/f��{yf�^cd�\�����:��m���k5�؏Ki��[��f����$�cUvE�ɫ����/P�ww�j�૭!ǚ(	 5�XqzԎR��ݸ��L��<�m��t�4k3&�O�~�BtMm��/�E�&a�aY�C5F� d�0e$�m̗�-��F�v��6bE^��,M�.����"S7~�A=q!�su7P��oufQ�
R|�'`ai"j*�����A�W��9vM8i�34��4F�ۻ�J�
�E�jY��cg[	��V����Q��HT%��5ݡ����������X�Tk1}�3�����h��5l2�����j�2F�k[b��R�~�9MMWـ��vVK@�֠�����ԓ7W���������:��]�.�3�j�;u�K��\�#��NA6��	���*_X1�]����k���l�z[;t���m3�L�U��(*V#GF���~�-k[�ՍQ%L�fLA���}C�f+@j�㨱h�Q�2�Ɋ�@@ඈ��;���ƞ�ʛ��!*VAga�y���Nҳ/$�ܩ.#Э��:Y�-�WR�
+L�����Z�:�N�Hn�W{��qC���p��M��l�������f��ֻ�A��!,K��N�9v��ڶ��Y-�6�au#v�յ�\��v�U̭
�[n��m�#E��]�Ifsd�C�ef#&����VӬf0m����R���E�졷n�Bj	2<�ɛZN��N�@:
��S�*Sh��/2�X�X����J���f�b�|�\�/���i���Q2��X�"R���j[Otn��Ӣ�_2��Im���J�×sI��FUܢ�{��E 9����7��8�гh7GT�	�1�X`8�#�����]Y�A��~��<SS̆��vԏ	��j�����ðT��4m:��5m�B	��[�Ѻ�X"Ցk(Ǧ�5�T�p8��Ӑ޼�e�N�C*l
D30�u�M7�!��n��zܖ�����B�2�v��i�4�)��"��黤�7�2���yCڵM��sb,���7[p2�m�{A����a�8��2<�{�A7.P�{�m]���ǱV�ӊ�᧑nPM��md��e]��E�^ր���,�+~ke��Abݨ~��Q9mf��Z̒�,�$SF������UV���AȉT�w1P����% E�8�Ī��I�^�k.�m1����iU��.�{��C�6��OUk�u��"�]���xr`�-�a��G77�262��v§������33j�v{���6l�F�H�-��K;��5(]�NX�,L�K�75��%�`u�j�Q��07n�����!��D!vƥ��i���e����3U��5��zȽ<�q\"X��ݰ�ZXX{(�Am�ɀd�U�����b4�����+.��+r��bY;3wv���p��ú~�/E�V��Z^�j:�XXc5��e��b��	�+T�G`�1�[� �NVXOP�%4�)3�T��2P�ަ�ҍ:��DX�IE�V+�J]k�Z���X�!u�e&��L��Z��,\�KV������b��3x3S����VY�%A%�N��Z,�ij��2uv��5{x,�_�<y���n�'PCR�����w!oH�iɊ�<��b���BB͛bn�+�I��ƴ��uh�����w{o2���9@SG@b �(
B1�3)
��a�!���8�ߞ<w�A�BA�
�HE��Y���4��;M�S��@%ZO|��6���XLl	�f�=P�C%Yr�[C��f����z����yo�{{�l���e�xi��)�/ hk�'Wm�4��&h��ٸ�RL�X��Y�����NCՒ�(뭊l$�SA8n��L���L�˟&U�u��*@�2��*L���Z�r�qo�����V�Xa��+�8(v�9ݜ�T�t���m�n&2������t��m�m1F�!����4-f6P�іj���ٗ6�&�g�k�uaM��U��1�@�6Z�n�U�C�U�YО歵/K�Z�nŠյ��*�@�9m�D�FG�%�
��X7��U��.�t<a	u7O�":���[�(�h�V	�Vd��į���;��֖h�e�\�{�8����4���,!�f_P����j�敀�L�{��8��L�f���;��Vuɲ×��V�0a��PZ�*�z�y��`�Y��^��cmn�Uݢ��H�?f��ՊrU�.���(�qB�����d�Ǥ�wv�l���D�Mk �F%RU�˚��eݸ�:��4.���6������F2��ON;�7P���l��'$��c���ętt����Dr�q]�+!-��Zm�+�f�϶�0���T^�^��HQb�4Q��3q� �����;���*�Qi�~[O�Sl<��x�n �2*�#S�H�4�e4���k�V,�l$���kQ�vNݽH��O��m�ͺ[Y2�Ж��m�˰D�Qۊ֕C]�yJ[h�6���nY��bX0V+4�&T��O��J�E;t�ܺ�n�{�oc���h�f^6Y��#р-;+�nn�P��T�:!9	Z�ЧM1�1,�!��:��;3i,Z�Zfe6�\yg6ų���p��SXʖ�S����ڨNPvJ�/YS5��E)j���#��m ��+��U$���K.=�R��eI��ȝ[��0�;a�y �"��c�A�ZM6+S�`6�jyeP#%'g%S��1�a�!,Z�xh&l������m� �˫�&����R?�к�%e7 ���7;��Е�Rƈ{�w[zti��Df�	�ui�%�y�kljQ������@PYE4i�܄�m%�c5����#)�u�ُ0�9��sѡB![N@H0���|�2R����+(3Fcq�Y�(��5B�m���m}�aUl�7�P�w��!�Rۏ �P���zqU���m���G��]F��j��۽��V/���1�k��VⲲ�H�`��ß��������&�ĸZ��Lن�Q��1�+j�ɼ��0���g7AOjE*�F씅Vv;���Y�C�In�B�5�ףM&C�)�	,n,�X	�Pǹ�ƙf����bރ��ܡq]a��gf��8�X�X��*hplh̆�㶦���Ӏ��hH+E��*e���i�u��bo,1���lZ�{53f	43*��2+5��@��e�ٸ��Ȑ��n�-;!��5������E��>0�)��H7i�s�Q�+Am�Zi^�}]eS�xYwy��1�E�3D�t�r���'K�M�4�W�b���5�Qc��3[��1L�m�mf*;�f;H�M����r�yIշ{C!>KBE���r6� a��ӎ���YWJ����	9mIA9x2�'Vq�9[0^()m�f'Om&�!I�嫭��mm�]X��hɥ=ܴP��	G)�1R����r�!���L�٬n"��X(�/DtU�n?�5Z�;:��ӭ�t�P�v�i"<ګw&�	�de���[��������66EY[S�&V� (.e�sK��E�;��N#�sr3���� c�p�����X�6F�W�n���jjc#�·f�a\.7T��5w�wD�������f� �)ͲR��z��.�6���ׇDr��eG�V�����Cm휸j�r�pE��5�FӨ!��Si` `g H�+,JԝJ4�f��t�%D�{5�Z6ӼʍL:�.��-���=�Ҷ���[�+r���	Lњ*ԤV��]c�3�RC�`���N�t)�@Zk$���A���w�ejO4�*�
�R�nc���bS��Mګ�7F�-���J�[�Ւ�L�;a�mƠK �vr��c����{H��xLz7ANi:�K�@�܋v9i�c`־��-ݴ��K�}�*P�ܼ{N*�&��,0��h�������Y�[5T۠ƣ6b�n���SM<Q��ݥ�����7]�������ֳ�BCz��`Q4�Ux`�X9�գ ��RTU�=l�D�j�R��st�3(U���]�v��Q���7�<$r�SX�����3.E��{�o:=��k5Q//J���}�5f�FfP���^|��5�X�pVP��r<�1*����#��Sm+������w{�wm�a��e��-�*�"�+55'����	����&n��R_<��{0�.�X�k�A,^cb�lYf�e&���ӕ�!٧���Xvet�#*b��z�OtK:,����z��gh�/�37Y��c(�I}��HL�l|7k`�b^X���7{.�kv8�����ȕ�61�l:%�ō���N!�2謤~����%��b���[�&����FEvU�Z"��vl\��\��+mIRLЮ�\��/pl��Rf( �X%$Y��(�V�a"c�l�[�i�iK�[x�zv��w����++ *T��GF�~Y���+��0V�ĵb��D�e�������֬Ļ�����4�7�l�B��r]��5>/�*]X�勐7��IK/j�� �n��(�L�*�ei4�O0�-D�g9uh��\C놌 .R�Y��Q�&`BX���J�d��[��	�7�o���̤���JF�X���͉q��P$�bÙUafKyz���g�,�5]����B��Uֱ��L"�6B���[�(�*,�Z�6�L�2���%J̙p�Y�,.\�b�U�
��(;�,��6�;�ԗ�������)YX)-�VKw�+�:6�/v,2�����U<�1��2�η�c����l�j�(	�<��׽��C��w�,s��</�aA�&� �1�P)�������ؾ�g��ϊ�<䖶�`|�xñ�	�-j�f�D�c��h�$��Y�&w�� L�e�Q�@'_cRn���Kj�V�D���1d�n����U|�c��o�p��b�z'�ƈšfqM%b�:�A�ëk�Cn5�u]�$u_0� ��q:�걃 �jV�p6��@S� U���t��@�{M2�2�өb����Ԗ-�F�D�ڍm�ȋPyg���@|1co� C@h��@��F�K{����>��jA���(^}o���]vI�
E�dD���i�lֹ�)�ua�2�:Z�GSO���T�-a�f���A�X��Y0s/5�]U76LKM�C38�`�|oE�:B7�����W]$���ufMʠ��hni�3M���)��1�8Ԙn��,���-�k	+�#4��.��J��~�g�sJ�-�8l�W~�[�s,��Y6|���2=�˸�{"�)��]�%�N<�\e3���7
(���BCV����ų�n�F�%�\k2q�V�[�M�%���v��(���|I1&�e[��ڕ�c?���c�g,��w[,E��_kv�NSl���#���Z��ŷ0�ޜ�-z�:u�8�(�������qs�=�ͨ����$�3[�}�ӭc��;ً�ʷǺT�&���n�btV�� �����j��cj��dz�5\��n^�	�;Ĭb�KIV�q�bX��Z��6�F���L(i=�����J��a��>Q�e���܋�B�q�gx�������q΋O��g0BC\���io/�7�ܸɕ�V,�K�p�[�B^T�z���#�I�队Wi�2�&�ZW�6�46�R���T���� }!���E���n<h`��C]9o��	у�=��I�ɑ��t���yuqj��F�81M�v�����C����f��܀��M�Rq«�䒭��p�^��;~���)���(�$�_o6�j��E��kv���5q�U&�۱��7K�m��S�5�	ǑXژ.�ǌ,��g;4;M�9�*f]G�tue#�]s�{d����{�NF�b5�]�,�W�kygx��
9Bn͑bJAn���kh����xh��-+�w��Sv��a�tv��dp���� �����5���Eʰ\Ӕ��Cw��c�FJl��gn�%fܓ��k��ֲ�):�0�×J��<�SqǕi��׵;͸��-�z�}Np�V$�ehU�3�z�i�=/��S�Ya�=}.-��^��#lɽ[L�`}*��䙕�Vh���K��^�B�}uq�8tVFF����ى���[����ӡ����
�7�l̈�R��-��i�W5���G����;�9�A�׶�ޢ�|業1�no!�6u�\k�#����<c� R�aFX����M�w��)�]��	����<���E�['Y��� �cx����i����ySY�b]�Y���.Z09޽V�n��]��X�^�tN>]��>�h���_N��Q��S"���v��j�ga!*�_�"DK��v9yW�IO.З��ϮK�S]����<�*S�KI&n���pnZztl�R݆u�7cC���ʲ�Ic��-"u���J,<�D70F��l��}Q�ˀ�Պ$ֈ���vʚ��%^��ާ���o�'��K+wo[����N�C�(�,{;iu����}��ӄ|T�@�7M����C泯r���U�l�lޮ��U3�Ƽ��8�q��FY�_��)��N�OѰS�7��407ܶ�w����%�&Xz͚e�a�������9���ws��pf�#n�~���������BW�s:\7wt�˱Բ��:�B�oF,��To��Q�ND��FF.�$YgB����Grr����|�`5/x����Bcʻ���Pn���=a��B�N&A]�.ج{CY{�{!�xn>X��/%�}v3��Ñ��h��q�;��@��=mg�y-�BYѕ}	b�����ǝ�e��&�=' 
n��5]�����V��Ó��4qu���}B\V5' �(��C��H�f�3
�/��J|̤j���zZ�?3k�ڈ��c�v���R4i�٦�g��.�ɵ�x�l��Շ+	��*(T�n�â�[X��t������7(�������ќ�a�Q����S��*B*��D��~�/����m��2�j���a��O�8٧�0N�Q����P�,�N����B*h�	�ՍL!�m��-r���v;�m8�De����	�[�,CZ��f^�'/y�#���ė�]ab�o�U#Fi]*Q�@�j�j�c�E�v�J��{{z_m�Lb�4G��{x�Ԭ��w�+�p,�\�$�ү+E_[�Ώ*=[�7�l����K�MQ�2��[z Q��yy��}�'dU��fۉ�J�Ӆ�֮
&Nu��n��Fv�*n��
p?��޳�ۼעZɮ��B8m�(.�
ZՕz�=G�-�)���|�x��pk+d�y1׼qk�����/��R�8���&9qK��J���X��[N.<z�Bff�!��ǌK%�]�/������P�ܒeYn�b՚E�ʲ6iK35��m�c�����ͮ#(.-��YHY���;�*ʂ�N�(��$�7����}(X��\�@�qj�xy���a�[Ǹ�VCg�hf;}�I40���[�*�;V�a6�h�5�.�u�j�ưc'�^�-��43!�f��7����$����ϒ��wQo���GpQ>���6��:#�{#�ܕ�%Y�m�
�F.�ں���k�f��9ׅ�d*Pɭ.�{��WZ{(Ê!ՠc��+R�v�gs)� �ι�:CXkw�.daw���v�DK8d]�X�z����m��c;����dNc)'F��w*��B�dX�`8�k�f���M�SÕې[�UԴ�&��Wv..T�����]���3���j�n�*:7��M8oe���G�����~LU��ՄoT�Gs@,�t��3��6,	z�"x4S4K��ï���<�u��em
n�M/�dK�$gX����5Y{��1�"���<�1�K-��Ы.7ι�Ş����YI���Za�1�T]F�u6y=ܚx��Y)��Y����aݧf�^C��v_�Ч�ڱ�IgM�jYn����Mǣ�2�h/
z|r�4n]��1w�w}4�"����Q�
��}�fd��'�*Y�ɛ�����j&�p-1.��[H���𳀽W�w7-<adit�i4Ӹ(�R��ڹ��c�3�#'mY����+e	���FH;���hQ	��Z�Ǧ�MÖn2Ƀ7q�����7�3Z��4�Ӗ�$/*��r�^���2��)�U�-�n�JС3m�Vղ��Zz�]۠�}���w���^�����l�����;f�c��2vs��&�.��˵O�]G��2`+h�*#�bY�ɸ%۠r�F.k�)
VG'�Hi<��N����=��E\�����?���2�ƨ�	�{yd���X#�����b�h�<�>xNurkUm�������W�;XI�k���=�Ұ'Rv�]��0���{���LmԞ�{k�������W<��fn��we��Ҳ�v�ŗ%���3�+;��0��[�ak�J!�w���, �[��s8��8�xٲM+޵6v�/;�j1��/�x��VYp��7�������r���}� L>�v�<�unn�}f�қ�i2s~<�5������\��U�G�Ȭ᫫��5r{Aak��ܭI<�2�7Ս���1��c��J������T)*��ux���:6Rͳ�s�k�)�8�?q֒�
�	�*=:ß��ۤ2b�@��$Q�cr���T�G(�K��O�g�XC�Za�d�Ye�v���k���ˀ�$ݒq]-u	Xnm��+�J����pwCOg#�����4���B\N�Ƒi��3��	�s\0d߮V_��,�����:���])ǻ\�S&�`\��;���.�,N�m \Gs:4�xOw~���[��i��4Y��[X���5�����=I�o�쥼���o�j�C�T�_5%���bF�i�����)7	oL��G�(������y�������u1q)D��C{}%m�Ȉ���j�t�w����{9��d�8�ʳ�6�̮Y1�&�r�\�W;N^�0-qS�!��Z�^�H�U�*C@@�w+�/�V�/�
0.q]��ۛvw�c�O��/�˴�����4���@t-VW]���䪅�w	7^�Ԭ��1ok{N�6ٲrW�[Yj?��n�,�E5IWn���e��2�K�Kt�P����c5wU�ZAȥ�c3BU�N�m٘�F��Y��Ԅf���
�b�V�&�ԗi�u�H��̽���wb��w��e��R�{�P�%cN.�9}6PY����Ļ^s�^
ʆ�k��oqMi���/y�0ͧ���Y��ӧ	��˘�é��Kg#ͥo��S�TY�&�o�s2�(k�AqIQ�e�M����]���ϙ�Z�vazM��E�ar���yF��%�:؋t��N�Y3Z�i�X֗r�u�Q��]� ���f_hӅ�d�ڄ���8�����jgZ|��r^�-�3�[j�]p�E�w����[�ޗ"XM�!�pS#Wwf�C}۷8%�:P����j�{�HeK�#���V�q!A�ݤ��<���� ��Vp�.�AWN��U/υ+�W]
�|��j{,N���K��C�)$76�(�t�Ӧ_u���Dp͵�i��v=�B����{E��ڃl�E]�n=�d�W{4ul�8*�zcS ��E�9�m��Y�b�1,�kq��S@=J��h����R��]-��)V����}%P,O%��j6�E���#`eB�k��*����R�X�����n�����,�S�\��ͫ�2��"�w��$�'+;�@��k�#m���b$��C �@��9�
�	C��!�R�s�}�Mu��i >����Lw�����tԥ��,r��y���;f�k��@�nՊ��=[�� sys
���B9����]WXp� �}]W.PS%��ָʀ��!�����q"4R��j��
��m�6^�d����Ȫ��LCۯ�m�ө�;����⡊�n���n�d�4�'t*tJf��%���}���Co9��BJt����gJ�3T�E�����K|	�yVm�'��wlw[��9�õ��)KG-��f�=v�Ax������%>"T�1����s���YI��w�OP�����6+�EZ7͚��	���'V�f3��J]���� k��ݧ���{�O.���r&8��^����
�E�v���Z�wX�Fv���Hu#rj:a��e�+��E�����!\���v\#t��}P�f���g���;A�q��^�4��4.�����A/�
Ɠ��N�(�m�O0�܌>n&�qS����;6c�u�Q�X$/9�t���{yWJ�ӓq��xW�s���V�ӏ7�ה�"@��F>�&��"�	���A}�fd�"s��ڽ�砵l��ܭ�n���Wfd�-2c�c����Y��rN�wZ�X��,����}�h=�w��;tx�4[8��3d5`���<��IN�t��U荞Jn��8��W����t�B*���[��1^�ħkg��.�/ �+Z'�DԽ��j�=�/��zUfݩ�6��Gc:IRd��t�}̌0<�j[X���M`G�[���.bT��Z�1��S����7S���ו��'jk-�6pd%=\E��S�3.�:�1k�rl�`��Ҽ�膼`���ʿ]\FGt�����7D@�v7q��p�D�B��81�f�㽃+Cme�ݐ��vT�|���C�N�/}�]�y��Œݧk��&en�췦Y�&�l�z�E���nt��8SI��;�1B�~�M�q�VL��xcy\TH��q]�GI"����,�y]8�ۻ{NP�KYne�h���x��#����n�;�)��i��s1}2M��cD�(ϝl�(��.v��[�q���h�4�{�j	W ٻ)��Ůa��W����mb�j1.1�|%��&
 �g��:{�#Pӛv�kgE�ȝ���N�)a묾���̆�l����h8�vtÙj�`�4ؖb��N7�c����wC���v8&nk�i��j1w{禋���ݘ
���n%���"0���+��3e;Lv�E�Ѧ�[�v������`�ʏ,ε�C;��+zpMl\�/�����z����C��[TI�.���7��M�O�[���J8RH�R��OR]�SeÝ77��vzlvE��CW�/�䲐E���'��j�q�5uf�_Q_�8έo�@���"����2�}�8������m* ;MԵ��02��i��o�wLڎ�w �d���Wl[4'`tV�5v8�
±3aW���4��^P]��\4�duY����KTJ�@��H�l/f�=���=gr	��t�]�3C�W�S����k	�蓀[y�>ReK�e>�sKb��e24�8�rj=��^.Z���l	�Y��ʷ&lz)��.)��wA�CbD�]X��s&�h��}�򛬗�ƞw���n��>�,�G�!|�%s������fm�����Ig�]_b��*K���W;�zf�r�h���v�5,�S���p�{O/�o�1��AL���z1Ǌ�J2�@��wơ��CT�e�ځխa�z��Յ���d�wv9������}Ѓ��in7�F��)���I�F�u�j���d����l��Hx2o���P�\��vP)
�%H��:�b��J�ļ$^\�r�����vcB���ǉj��)��/2�tС��	/w\�U62��Ь��X*-��}�kz>�� �J�r�9c25{�;�r99H/j��綰��+BA<MS}��7�b *I!�q��6@���h�ﶴo����颼�������^���_.�R{E�t����?R��+�H{�|I��com� Q ��������" ��R~$=���7A��t�籓�EE��O��<DA���������҂�������������}�������߷��ߕ��ől`XM�T��j�#@���]��tA�:�r�ְ�L�a�+A�t]�`:�rs}��u;N�]�b��|��m�9��v!�e��r�foU�W�����D7�������{�nk+J{[��s��go�wnK�0�}��m]t�v�V������٥��<<dWaea����%{�v`Yނ��ɾ��%�q��;��bk,�cΒ�B;h�8�څ�5&z�]9�Г}�px45�m�9�Ejn�Щ��˜��X;uLG��Ԟ��9�����d�d'�`�l^�b�n;�a�3l��芨,Վ�z��U=�K*��3&����v�u6�Ăt��+b
6��^�V�Z�Fytt1Y/:8�A���h,d'(��͆��LQ�
j\;C+�͏����;�KQ֝���k��)eX����S2�x����sKќ�������#STF��E�%�����^d����$�5 �Z94f���}���o�s�BL�F�tҤXs��!jZn�;��tI��5]�74�<���T�ʵ�Q���Y�����F�;e,4�WiUs)l��NB�LX�� ��f6�!�s^[�:��P�y��k'N�8���8R�upK��'�Aɹ�MoB.�(Y�Lpx�(�����}15���R摔/_
�0��t�(���mL�6�&Fc7��+U�>\A{%v���!Kv^�6su��<6��J���U�uy$(�yIm	YR5%�����c�%E��SGM�9���)�馷Cl�Z6���\�i�se�N����h���HW�ԓ6�ͻ�/)܇0��ku͑�K�`�\��Z�T˳u$�{Ӱ>��8��Lp���!�M��<]�cU'�I��A�����Z��M%!3��qU|��Q�8��Z�z������O\�v��7()Vf.�	��]�7���^*$��.8EX���d��I�K� �v���Jl:�ڷ;t/���B-<LnJtƄ`��Cp��^s#��Tz�r[]�M[�C����N��"�j.�v���yu��ӊ�u�Se:%]�UL�-|�f�N�Kv��a_�����vx��Nᳪ$������uc٪o���W��rm+�s-��1M���j��@��P�ݦ��X��7$��*(�}���@�0�3d�"XMLj��.l�Pփ}�>��%]��+-�mŏ�����3�²>�c8)��N�"e��z�R�պ=(|��΍� ��'>�d����^��T�	��2�e�J���-��N�K=V�)����M)�j	k�!���\�Ux���n��l��}�Dӟh6�c��NJ8��]�����TݠM*
h���4��L띓=��W��Χ\�7V�L.S&խ�3�Z�#�̬��	��V8��i1���/E��`F�Z!����'lwN��`�4�b��jՙ��]�k'ۘ�7 �	`hY�{�48#�qlQ@�(��kܹ+5vL�
Mö���r䇮�Ub�J4!���#�MvȎ�Xm����� НPQ���!T�&t�͖e�����Y��v�)wR��]����ʲ>���Lu��P�⎈�42уO���.=\�U�aӄ�c�>{�z��MR��R+7�M���Ax)Q��s��'uV��ś�j�'9C��)L��Ṩ�
��
r<Ɋ��,�X�p=K-���\hf�7y���r���L.?�Np�]�T����NP���$�[[����wr���]lpqۨ�U�h@�la��u�l�v jn����*�Ǹ�[�ċٖ�V����w�<�,���|���w:�����NY*�^l9��ow6_~�}��%�ð�sC�Y x[u��j�&d��fL�����Ӳ�=�����Y�b%�u�6���|�c��ݢc�,��0h�e�{C�%�i���tȢi�	2��pt�g�:S-��N�'JU�&K�T]�-9HNյ���.Sg�d����:�x2ɽ��l�Ks^:Lz�_Z�q�:=�A�?oP�c	/+Iu�1
��ew6U���T+���8�v��������L��!�fUޙ�@�t��;��/h(C�ڌ�	N��^�-��eŚ���{-���*i����B�ǀwV҅A&ez3��W25�f�,�&�WS�'��Y�L-��{6�{J�"�Q���]�ɛ*>�"�t�[D������ݶ����"O������e*�9,]���٧*����3�����p���ua�y���кH��Oc����]��Q�e�t�ki�|���c���s��V�	�E	w����妻rhsX�t8t��J����yTq����H�}��OO�G��������J��Zq��n��v/!&�t����L.��+��$Ia�m9�Yّ�m�m7J�X���OҨ���P̅.f��B}�BP�����6\�K��q�Л�9�_3�*�9�,Nq��L�Y��ǵ��MK5�}��ڌ223�����3�+Nۨi�C>��u��.�.�H�D�s�+���ʳ6.9S&�c�3�����-��e!�Z����N��\���H;���8EB�6i�4��`�&��9��jUa��MТ�ew��f�_T�w���{|j��!�1[\��H^�1�yrGu
y5sc1��|/�ԭ�P��D���I�41���c����ށҒ���w(�(ΗJ�N�&�*;��6�,�6�D�����R���0Y�gqQ���۝�Ẋ#6�i�O"��n�����\k"dŇ-��?h=]wG\G�:�
'Tu�V�V^Lu}d�z��b^�쑍s��#������+o�csD�kEwC[H�W�V�{]HmGK���i��hh�*]�qJ˒'XJ�Q1tY���*�3��O�؃^�ut�f�zK��h�z���H������jMU0LQ��\Ǻ/�ehc6xX��ɼ��
P�1�Cwfo3osz�#v�5^��1DÚ��W�:؁ia���V0��&��=�F^Ua�w)a5d^��^�u/N�gES�6������`�����x2��x�,�#�7�w9wZ�9��I����gn�5#[e.�����e�o ���l���2���9u�9x���v�3+���P��)Z���;��eKP+�n�-�5hs���q�t�B�	��<�ܮc�T�`m�C{j^�S�6�2AxU�툞�wl1hdp�ai���kw���N��)_1K:��k,.I��U�W��L��+����wt�1�5A{&�P���)�Y��C��h���=���n&����	�&;��Pc��I��)u3iN�����L0��x�!���@�@x�8������$�m84����vYLE1�XKb��7y�A�w)��2��j�Έ�f5���o�ϓһ���h�!��c3��T��6�pbU[��y�[At�xo�6QI#��YWzjº�X�V��9!P��7 Zh�e��ںi=;���B�|J��*v�y�N�Ar�k�K,r�&9{j��wã�9��zZ�Q�Y�r�@�m��t>�Y\S�j��uD�T��/VI��W���,�=�f��Oc�Z�����mM�]9� �!o#���Iv�9�YVHtD��%t�y+�d6�*<�<9�X^��[�ſ�G>a��+��uR�2}�s{�Q��L�%�"����g󓮇�%��0�R��V��뼲�=��zz)2ĝ����{Co\���v��.��e��s�޶���y�5]A�SIK��[��.�=3�LJsgۍ
��de���El.�?�]"�H»�d�܍E�4�����+q�Y��ܛ�6���yո*��8v!p>�4K�W���ؼh�f�v�4;TDd7G"���� #�Cz��FE[��f�$�#JB�N㎙)�'�4�N8�gyx {s�$;5I-�
��	�4����'g�Z��&J���/��O����tӨ�fm����i�3@$V���0���,�8�K�,��U�vJ�2��p�\֓8d
ح�S��P�� ��AV+3r��L�'m��~%����%s0A��B��7�J*���F8B�s��Wu�.ǣ �܌[�D��� U�Fu���sz��ڐ�E;jk�Y3+5�̛J�ёr���Ja�:^s�h�\�>�,����"a�R��%�7Zp33Xr�I���IS�G�q�"
�};2VN��z�3"f���$��0֩��F�_�U3�zc@U�n�Y3x>�GJ����`BCմ
��hR�v�e�ᳰ,�����F�"�],��O!��bL����ID{h��GPu4�">�Rv��ső���K��=��� ��)�à���ɧ��r�2%%�+�قwe���Y�j�Ӿ�3��[P��X��;!�te�H��|��7	���񃍬�i��5��B󖼩�8� �Xf!���Y5EP�Qâ'�|�ɸ��W��Z}��SSW�$���.�c5�ٴr����q�C*t�T�5��,����H�p�w�p2�^.ͧb�p垂p�mT_d��y��yΣ"���ǿ$��3���=�����S��/����Y�@���|)V�7��+ԩ�&�K�d�Ѝ�ꂚ��um��R�{;3"`k��Zl�����5]mٵ��=zV��á0\;N�z�G�|�s�O��]��"�]��Y,�ݶdf�Wr��òT��Aܠ"��t���MHr,ل�+v9M�	[��^��^�Q����3:��F�γ,U�Q>�9���n!�I�Kt�Vp;�o�dW��[�:��u���Ӓ�U��̛�>"����wOD��y��[y[���-n{����FM�z�l*�;� �j3�:VO�coo@�z��7oK���O:�5}[jA=���e#���"�&�]c�{��H�S�kyL=X�o�H]�W�$)[$���PƳ"��K(�X�sCX&�c6=�vu�鲗=}�s��R\�����"�^��7Ш�Ù,��h05mq�B*�\a�w{ϥf퍶��^�
u���jJM�n�:�ʗ�A���4v��R����Ɯ6���η���:��ǃq떈4aoY��=oA���\�/mU^IE��E
ț�{����e�K�j|�E�Dy[|���]|�Y,�V���X6'����a6�8��-Ŷ�6�]GB������-��FF�G��A�:�~em7�i�)m�ݣ��:�p�xZ��)h���zx�Ɵa}��f�9��
�������Y� �4!o���r�YzoE���#�)�a5l%ݧ��N�L(���[ǘ�Q�Zi���3Tej�a��EC΋��c`Ǉ�K�rTXdӨ]�FV����D��]F錱�	�V�%:ww�l-�։-M���_rY�¹��t���0��x�/�r�C*���Մ�z���!�%�V_E��w7�eu���dj�y]�S���ܲ�i��}|ksںoy7����B��y�t,˸�īEdE��I܈ ���wK[�VU_�B�7o7������G�P=P_os�*$E����87Y��`�v�떗�Vn��et�� V�|ys���|)�Ző�4��y_D�#�8;�pRb�7���e��;�ݪO��ŵ�[��=��]/l%1J�n�\2pս��ŗ���a(���D�@��'Jܥ�e�0�PZ���w6m:��g'o"OP)�L�
�}��pw*��Sd=�2��V�$N��/�������] �`m���nlwNqo��j�xq������a�</JƬSڔp��n�ָu@�mU����{,�Z��aw��Ҳ���oC[���5ޱ3�\��лmT��|�ӤF����	^uv�g7D�A���Vn��������:��n����
�WA�?]���y��ʜ�^	��W] ��=.X�gi�9��VXl��{�:}v�u��3�hX�quCv#
���h��E�Y]��:��V�֪f����<�nʨ��8��%���j��!�n��G�-��0�Ŭ���N��6x��ĖL�NmdHf����*�^I;�]9�t��3b���*��H��k�=Wu�V5�7�7Nv$�SqKݦ�����J�#iٰh�8��y܆t�Nk��RqO\�{j�����
3��rf�N�d�9��A�|qY�N{}ؠ�|�����b�d��gL�OC��=ͭ��U�wa�iщQ�W��I���Է�E��Z5�K��ćѭ�gw.U�׷W�(�pЈ�����p��Am[,.��r�M��&2��\����G�\��q��,�[��U�"vړ��9�ݗ�d��7&tl�EM�dY�i��ĩg^���V��8�|E��\{M���׉���f��ɺ=i�޻Q_�T{�2��{�Lp�ͭA��o5���S1ڤy���
:�$�	��[�pk7������n�Tq���7��^��ٍg]1&���:עdQGM0f�m��uV�Ԯ��]HQ�]3�/S(7�|q�݁}��`wč�k)��R݃�����˽�U�ޛ=�;B��8��8�Nt�N��;2����Nu<�7�&�Ŋ����G3w/:�u�lJi�s }B��Mm�o:W+qn*�Nm�]i�;x�Nᬑq�˓D��ԝ2s��U�nt�6�t�W��ݘ��5��o�۴hG+H����'q
��}-��YJ�Ֆ����BNԶ�E��2��owj=�x�ޒ�N7�/#�,t��a����ֳ���&X�ާ�)72�/�R�X��4jA���b^e&bs��B���3 V�v���ڭ�7z�/R6-V8����.�>e���=���n*B�r�N�`E�=��Z�*��儾�ԙ��vO9Qè����qr)�LΕ%c�>{ϟ?��4W�P_��?����E����Y�_�����||||1�_��fp�n�>��Gχ�|���E��v1�y�u�y�˭ā����ʟ�jFAE[@�PD�t�Q�M��)(���LS���K��]H��H���kܐC�?s��fn����0�Euu�������8i\5���z6"{�|�#�]�/��	eRL�a���kWl-C�`�gq��Y7�G�q��#���C���q��^[�Qܢ6�or� �eV�"�çL�D�cU0��U����n}`V�WN^Ә*<�7{�&�O����R{�ƛb�p�N.z��m����.�fe�> n��k+u��O��B�m7��.���es��/�d��h��dѧ�����I��
ʌ�`j^����r�l�7F�Ѱo@x	�Q��y�Vh悄�gUQҥ�M��̷�VlK'l<j�ކ��u% ���\��ɂp�OX���|�����WNr�ũ�e�(@���Y*�n��j���|/�h��Џ'�j�8Q�P���J�í�3O�f�nT��6<�N'0�V`��%�rpq ��ۙ9n�Y!h:�>�l�ؙ����=G�޾
�O���V�ػ^!������2����׼&1_���ju��)�{y"ȀU�)������V,���'
֨f��6��-ѡ݃C&h�rG��l��]��M�=�m�1Y(��G.��ѧ��X �U��,cr�8��]���/��I6!!���-��喞�$��Y�턨�8�mY���m��Hb8C�H���)�D#��K��3D&�B"��H
���L�D̂&�F1$((���n���˼j-�y��N�j��X����Gyxkx�w��kZ���D�l���D�9�HI"�"B1k�qy�����@^��t�΃mM�IM�����UN֮���4c��t:)
t(�@b��
��(���Hꔠ)6�h��l�CHh4=�X(5A݂�������]&�b����X���"4���.΂�x���-�i�F1�'mIAJ���
'��b��F�:t��5KIlb.�C�Eu��F�zuCv[�����M�S��R�͠��訨-tpUwa�t:��J��Q[j
(t��#�����۸4�Wv�	*JnΚ{a�h�Ѣ�gX��uѷpj�1OlPѢ�ѡ�����t�N#A��II�H6^�-�"&N���н���j��h��׳�1��ɻw[�ڽ�R
�B쿨��\�՜�'Ay���y/l���7�;���/���@}�1���b�: �Ek�*9��s���%[��-a��%�HGo*"�*�A�ίE ���$�4�f���n�����T�����8�X��!ɻ�>��f��^�/�<�����Ҟ��q����[W��({>��� �m�I=~恔������>�=����q�q�DcK�WU�vc���1�#���~�r�]z�~�)�������c�=�=lz����	�V9�����{���~�z�r����w{g�����0k������q{*>�B��܇6UF|�����d��U4��֏����������{������T����<h1��;�<Nm<�62�� w9Sf2'}��Av7\�6
��`WkG��`����ON�mW��}ؾt�}�.龹ЯHt�b���`Wq�9T�%��T��k܇��~\=3���>`zb4���;O+h��'�M:��̳��������?a�n����W�}�u|����_���\�i�G{�_h���0�����5Jɼ�ҷ՘h�E�9��th�3�7�����9�˛h���k���q��H3`��D��N�����qv�d�:.�Qs�)�A�5A�n�,�db�����e���QF��s؟HrGgu�UO��
��^����r�g�&��½���0�]����>�D���B�r�4!)���K]:����w���Ѷ���3'�xQn޽�9�l1Ώ�����������+�����5�j|��xD��z=��W��Ѽq]���+�'�Y������m�=�6�hgW�����|����!Y��6���k����,��c��˾ڳ�����c�W����z?ʽ���������T;�1�i�z�xڅ���s�Lr�=P޳T>�����E��zB�V�����o��ݢ�l1��y��U���l�O����͹�|�>�z*w�{9�uP�JC���ѭY��9��o:�Ɯ�fN���n7U���'2���w��������Nxk:�Ż�Y�o{���4t��7�;{Q�O�B���j�;Ȟ�F���ɖ��p�Z[2�b�뜇!���,9Xj+��ݚ]��QK-�J�{:m�գy�ǟ㜇`�&e�%g뻽	�l�"Mk4i�[[���Cg�)��]�����[�7������3�"�kP+���sڊ�IM^g�9��y����|��J�r�Ϻ����A��3ٗ�Ě�l�4�,5t��8g-k̬��G{�X�k���G�w}K��I��~~z"G-n<I�~��1�z��.Ɔ2R�WM���`E�l�N><���j{�����B����j}�Sr�Y�4��g�}p�?J�%��6oeC^�z=�9_�o���<k|�L��{|�O(u
�N���W��'��w��w<�u�#r�\�O�����{��gz���P"��E���̓v{�B�=��>�^��xל�������ܪ�L̵�[�܂L�q��5�vyV�Պ��me9�]�Usnu�n'o�n�{�ɏT�$���ɼ�r��y��p��5G���Δ��3z����3;�rn��x��U�qy7N����}-��| h��1:~����~�ߙ.�x����h<��s��Ҝص�G�z�P�6���.W�qY]��__7t�9�6t�VnϹ+o���p�Ո�wz���������g������J1ȑ��W�X�\�]�����*�Y*�,+fu�����ΰn5�L�{�����2�v}�2�8�h��o���� ��:�A�k{���<�j���$��=z��}NW����ⶭ�a�p�3~f����9��-��ֆ�,z�0�j ���X}���'*�����d�Frz/}V��qR�S��{��䝣�u������$73�{�nW{Q�}ܭ�I��=�ҽ��T��zq��L5�>���v�]o���<xc{^�Q��v�~��K�.[U����W�By��O~{���ӭ�<}�	3�b�;�ݫk��霯���5=�G���x��/�y�]�ndN���������t��m�^vA�]�Oq7��8��`n3���`Lj��)���گu���́%�fo]���PccGv�} �[3��̪
�2�0����β��ߑ~�3�i>��?I;������О?)���֜�-;v:�����;��n��,�̆p��X��/7�N���Mc��Żj�	�.xx�{@�P�<w�漖�>�mҚ�x��uvfGy�T���	S��V�)WP$%2\������ ��H������%g%C3{�*�ӗ��D�;����TM즞M\z~?T�!9Ń��-gL��|���^T�9�f{d��CŖ�L�M��Шj��<~�����eygչz�j��:�|��Oz7��˔N:���ߎ�>��A�޵@|�^º �%��뽸2a"v�轐��Z*��b�{��p��?/WV{�YZi��6|�����v0�}�-՘u�tia13��{��}�$��4��;nѦ��c�TW����Ν�d����%T��j@���z�d����^��MM��s=� �''R�]ݔͧ��=]�}���5�6m6�H��?v���A�0r�\�R���U��e���r���[�S��xu�VP����p�oZ����޳}ۦ��e羢Y��3��3Voo���:Eސ�g�.��4.���uwϻm�y��GŢ^OpN��W0����y{v{�o�{p5;��@_eW�v�y��,��<�4[�s�l�� �ye_}��\p��d�pc��Ldf�ΌݦB��̑�@6��c��v��N(��__���h�F�8M��S^f����ٻ��B�c;d}�p=�V��g*ٶ�C.0#Z��ʾ��`�,l�ڡ�)���m�gt��־��!>�K��uy�O������[��FW���0�/}�0tf\dN/ݩ�y�ǚ�x�LO?o���<����wn�c)e���v�E�αK�<OW��j���[�8�z]=�k܇�� ]T=&��yN���=~/|��>�T��v~�=����qh&[��pv.�����s:�mMR��߹����|����t�;)�?q�|](����o�<����s���OW��59�5��8hG�R~��]e{��@��]���]�0]�ݙ�����bOX�ʼ�@�#{?,{�>q��k�x�҂q�����}b���{k����,D���3G��-{l����[潘�E���oأ?a�x��^6�^o�I��W��� ��J������x�Y�܄W�'�սq;M"�c�ȭ�^A<1�|<y��F�\�W��-����nA2� ���^��k���9]|�Ы�K���k]��8c�k{�	��Tˇ�!����{��ŀ1��O7@�P!$��c�c�-j�z-v�luÃ����P2�Yw{s�G4�ټ#ё*ձ��w��},�P�˞�T8��yWa����te�E�;��{�N�u��yzǳ�za�:��YޑO@6�{M�j���i׽��z�����z���d�=��ay;g$w\n�������ץ�>����S ��{o69�\�MU=��x��r�w:#�j�ɋ����+��Қ�w��+��岻S����S����f��9��a�F���7m�A����o��'��{UV�<Vm��fo�ޞ�ڽ^�.�C��-�3ݦ>��"���)е������c��<�gۮp�=w�LTz*�~Ţ?i�W��{�k�m��Uv����χ�5��6�r����[=�F���O�ߪ���o�~دOޅ�{|�?&FP�?'g��g6Ѣ:n�4H9��LM��1���}���ǯ(Y������;H*����𪑏z�����:(o��G�!nfCh���0���|B�ʿ-V�)�*B���	����XR�qp���]s��#;]��	�0�h[�nh�Q��h�2<�<���d�w�*�4:l֕��T���e£��Ea�v\�w��&�b��zg>rڛQ�;��]oS�\�P8�Aw��f�+��WsƼ��NO�-�#�K��B��4G��Gt?-�>�L[�=��T�5�Ӛ��Oj�;2V�{�49���v��q����偊�m�x_B� �U�o׃u�|���#���npg��I�'��W�͹���cv��Fy���{��o�{�VU�kҼnWou#�/W��p�}� �:��h�����o��W�h����x����$eoO���^E9@���q�m��m!�|���v���{��Q�C���Ҭ�0����g}<��z<u��O=��v�#�y��=Ez��N��ό�����W���M����{�o{Ps"}��@d�^��>x�o�=��U�`����R���}gw��x}�)"O�^���o.>�]������9A���R�1�j��V��8^WװW��t}��`�����|��ęN�̍6k5�5�[�P�o�7Q�i���yK����KHM��{�Dj%m+:��җ{ɂ�)�(��S"�D��[��� 'Y�3�M{�&�5�L1W]2�+����*��(�*ל�y*�g}���n���{�?.�,�
��{`~��m��]8�[���y%��s�q�{�Ow�W��h�h����A4�]�J��qkُ�h����s�kɏ����{���ﭚ�9�r<oX[؞9�E��T*���k1I�E��̩��ш����P����>[Xsw(��mԀ��O���!g�a�elԞ�#N�t�oe7u���Iw�Q\�_�A���5L?:R����F����&{FW�L">�ٶ%u�;���kQl%�M&��yga��)��З��QY�Uu�ΰ�m�'t^5=3��7��.FH�,E�2i��a�σ�C_�U��M���&2�D���X�9�WVg2�t�����4��m� �@������*t������{d�RU�45j>;򦚝�3�^
�����zY��!�6ƃG3�"-�����6n��j[���e].�)LrF6\�,���tBj��j��lمE9��b��ݝ:��>�s�h0��-6-l�Y7U���`k��y���Zy�]����aO2;�[����3N�j�q�:�1��|��+G<�)�J;WZ�K5��J�J!D�}��^�Z���Z��h�}��w��FIr ��&b%���C��{��$�f��� �{��CV�*=늧Po�΀�,#���i�p9r[���V�w���9k�q��ڮ�i�
m�������@�^ל��e�ա�YԺ�<���y�k��Ǟ�'��
��a�޼Y�c�����[��ڞ:��Ü�ϯ<��-my�k��.�҅����T	�h~̭����Ϝ��ڞ>�g����ϺB6���m�\]+σ�ǴY�B��K =�xH�ݗQׯ͜��ؘ��=U��&+���f���a�#�珯<:�.�va��N��v�����9�5֜��w��umˎٲ���$�����x����g�Z5n]/N�}q���f}W新ǽ/��z�~�=��G�~���̡:��b����}�z�>oo����z}>�O�{<||�o?����_�p�������N�^����7Ya_Cw��[(�أ�gXUJ��к�l��Դ]Cܱp�.��j�s!̽z�ɛn�[.N��� t��1&�҃��PkN��S-��q����i�,�rK���09�i�q���6������q��������j�W�.n��6��V��z�H/����t�V.�I��˽��H�b���iX�*�nh��m�`�q��&ݚZE=d�M�II�J�C�Fa�c��E�"���R�0Z̥D�FA�ޡZ�
�AuY��mm�L��\�� �1`1��n�P.R��7^5[j��3%%4���Y�n���Pi�yCMU�^��ʛt����9�mr��ݻR��w�^�7��$������7|�ͻrV�� �Fi��άS�fK"���XO
y���{7z��`�����H�ᕸVo%�>ʹB�:�Q��1{��P\���Y�j�K�[jm��!�k����'��NJ(�Ib���c��~ �]��[Ձ� ��޼�)���4��U�S��.�u��"H�� 	�rwv<�1T3n�7�B�E�.�ơ3AR��Tϭ(eŕw�o4��SI��_G�]��.sH�6X�*t�$��[���G�N�󨻅i�q�ʹy�M%�e�M�y%�=�����J��\�%�}��2��Vo�\܂M]�p��i�3��2m/-�hRXm���_�و���~�@N�}e�{�0�-g���N��+(�U�Rk� �j!u���D{�+�g�����]u�<�Zŗ�+^�|r�i.�٦4���ԗ\k1�Ku2@�,�x������\�`֎U�/s>�i\�Wn�k�òչc3�3Д�J=L�Yc�+�ג�����+du��W�E%6��u�f_s'jcs���[�<��k:���jF�!��Mf�Y ��;L�==�4��4N�#��`�vS:r��8����h�)}Ց�*���:4h��;���u1X����� 4]�iC\�R_��q�^t3�p����z��T��S�CT.S�ǋ+��T�+u�6���r��%-���	�p]�0g[�(��}�Ȑ1n"#���V�1�ݿ��u> V�I���=��ª�嶨�#9�s]�u�zIz�q�IY\&��8�Θ8��|��g��uϬi�2��������x��^̵zz]�ے1��ǖ�7w9Ծ߭ζ-��Mw�"i�K�/Y8�UQ"�d��W��׫n��
%o���06X��Y�3��lU�8`{9���7x�z��P��˅m-g��L۩4���j+���\.�kق�Z�]����.L�Z��D<5Τ6��3��?r3%���c��#5�g5q���;�������h]��޻�Ʈ$*�:�\�.@�o{҆B6�r��}Zػ�B`89�4�6}E����d�g9�RA�9x�N�v��t٭X���pt��+�x�K}�Ө<\�-��+���z*C�4y�tT�tVm%]�'�<��|�.��.'���� ��T�6)zѼ爦'���4[m�� ѓ���b�Fg8�9;w��:#g˘���`��E-��Ctq^v�|(����mMv{��ǖ�<�l�^g�*<-�-7]n�y�U��(�>n�h1:��Β6�cy�^�]j+cF�AF�>Z:�ͬ�cd<���F���ׇ�M�wy�L�m���1��ֶ��o<�Pb;��=ƺ��.��<��z�m�/<�G3�^G^G�F�=�vǜ���v<��[��⷗Gy���yGw�v�4��.-QOZ�j��h�k�Umclհy��o+�k:�b��V�.�'DZ|��<�3D����y�;��1j:���馪���t'K�'��<Ƣک�9��TIK�ukZ1ظ�mc*��GZ�K��\Uּ�/ ������`����ST�3v,�v�[�;��U�	���~����#�Y���^�Ǘo�(�BV8��c,�H|OJ��6�����}���R���{����(gQ+w��x��� �H�d����+��a�,�Hs�&��n��IB{��v6�vι�^��ȿk�b$��ۆ�lG����G��M��z3u	��	>DA-P�|�{�I��t�2*E��+�:�pl��̪��ҩ�))A��K7��-�趃��p�����en��͌�~�ihD����~�?tuq6ë�Tת��7�C�ke��;l=x9:]K]��dՕ��")묙���M����.�J"�F;��c��ytxԾ�<��$�|����F�9�1e�] S#�:�e��Y�Z�ڧa��ã��@�@�v���Q��9k���
�hkr ��i�׽4�ϩ�>ځ,��Rc����}l�vN��g��:Y��R�۞�ܾ��K���|��7��(��2������{^�kP&=����j*�F�L�w���w@(A����3��y<gRV�7t/�0�(����� �s�/ə�k����?ӐǟkP1�"�/�4<Cꉁ�*���3�o�F������S�n#���|�9}�r ��Eٲ���c>���>-���v!"u��\�4=�d�e��s�5dΡ1�FdcN�/t��h#�}���!ɪ,OO��-b���~R�Ԭc6�w1;6���+0�*V���,��w�Y��J��#�þ���w}�|b��������.o)��z�ʦ4� ���{PhK��R�ԉ�_j�l@�z:��U2��V��V�Y�s}��¸���<y~�����1�?�>ZD~{���"�t1������9��� �30�\e6��q�0�g�е��^y��b#=��N���$j�������^���FR6��a0�b�ū��GP/Ɗq���"��~�&���\b��`�`��Tj�p���}��˥���{��t�
���k#ؕ��\�P������az ͗���o{d�F�bLE�y
)��wW��?���E�\��>����z�����;�.uުG\��c��[.�l�Z���߷nq�n��~�ߩ15@�dDʝo��Ͱ���|��Cv'�Λ�E/|��2��皚�0�}L7�����ﮑPw��.���jj���ʲ|̊�cmN�dR�gn��&j2��d�BP�3oB�e2�XN�l�oH��ܡ�A��20y�5�?_�*mvXRv\���(#V�=%b�/ns�����֏���Mf��c������yn�u�Oe�:�^�
K.D�`���n�Opg�dˢ�@�bX�fY�U�qD���:�7���,��7����7�9���/�a�jr������"\L��,�Gi�GrX�:jg3�-p�pL�u�m��˖��gM1C� }�s�>�����_ه��������	FLA�NI���K�G�[�O�0��	V�oEjj�<�3S��x�Z��k)ȇ������b7�+��q6�H���� �GU��.}�?>k���\<hn��'9t����r��|5#[s�~w�q f@����\�M�+Tz�9�T|���W�bF��R3#��Q�}A<S.~�"�{�Y�BL�LW?6Z��� k�ܪ/ܰ���ƽl4iS��ym58�p^��>��TǙ��0�y��|��|ϋH��`!|zR������d ��:��P��}��- _kH��&\p9j��F"��	l=��Z��B�������ܖ�elլ�m��� ��)�1�t�X,���6�ިN��q|�������"\��ϞXާ��^���>o�០��4y��O��9��e1�E�@����_O;`P��[�J�;c��k�v�_n��%��1��0b�<8g׏?�ym��D־�XʶLh	�\�`�냳5�1�N4"�`N�<�_\z�D5�yW�gK�X`��控���BP�7�	��\���>��̈�K�fy�jܥ�֋�Fb6��3/�j�'et�7���fQ*l�7�9A�g^V\�I�[��jwQZRR�P���h㦤t�4k*>�˭���=�wR��
yK ��@fҾ�nq���u�h权7xVC�Z<��݂@K�oT�Բ�R��dK��\γ��������>�������P��:|�~��a���eVti5Q�P��:�mç��~ݎN���!���c
�`��ĳ�N��4&#CޏB�D1O)�ʹhjȫ��X!l��5 Zȱ��s[@�hl��0�:�9	t
./e�ѫR(_ʼ=�E��z�Fy������K¨�J�S�g뱣>�ħ1���څ��#��uG��R��0�fÄ�7ɨ�D�lX�&9j!�y�d���M`��A���{N��܊f+u����e�Ƶ���Dൕ�o������魤C��t��i�<1�\��`h��dA��E����[�j�85M�U�X!G��T¼��T�}rFdT��x�B����z�V�yֆB�m�=D��19��Slv%V�V���jq����6*�Š�����?D׵{.�����@f��>�t��R��iIN�׏�F�a�>1����u���ԇ8�o��f@?k���>�i�ɠ���=#������K��Ԏ���W]η<>�*�c;x��s8C1�uu�4�4�W4��2-����cg,�u3{*YZ4�<Ǳɋ�m��@��{7j��j�����h����=�W\ܑ=\���%��\���@�ךne`�t4�`5Iwh�����x�����-̾rE��_� )�U�bk�B^9��Bm�m�{sU��m`��+����T[���xAn��XӝGG1�M��`���Z�@~}�B)��B+��aR}�,P�������/B�����{����SFXS�i&g��K�Q��3��@ց��!�7B4!��s�s+���>����.��q8�8D(��OF���/MUɯ��VG���/G�ca������י�iƣ;�e�1#�'��|sC	�	���O�|�D�OVE_��C���R�y�Fb�׼*�]�EŚV�a}F3�� b��;pCO/-�ci��B������J�ūbɽ9N�К���,s�ƚ'�1iᠹO���c�2}�̼���ov�JT�ylϢ{v$�Af8�.��g��ށP��>�`��U1`࿮Y0���)��E�X�O]/�E\��P�쭚�|��/z��R������;gH�W�dfCߕF_����DR�ߠ��V����h �hit����2j�m�Co�V����[&F��qh��oG��Q�g2���^���;��9Zې�\�����Yד�6���Բ�|�*�ltb}�������X�Y����b����q=p4����׈m��M������g<�j�2�v/���@*�+���g���q"��읶Q�11m>z{�5��F��c�y�xϬ�oJe��r��uj���7`���z�l=:��8#L�7#g�cR0n�/+��|j�R���_)�ХaI��ӓ��^ժ��N؂��U�#��㭇�#���������c�|�#F�~�!����7�d_�n7�^d"�è����S3#�t�U!D�n�m	�^�v�\��`y�v4F84%�sЗ p�&K|d���jD�b~wC�)���f���Q��?=�_*u���Q�1���#_l�ߧ����F'�^bs:��}[�����ۦ6� &���x=����N)��H������}�J���3��G����qq��T���U&x���е�� ��ja�G�}�F����8�[�O�=�(��\{)C:�nZ�.�c�yC�;���q>y�J��-t��j��Xh.R���}�[G^�� Pq�� ��p�c�w#�g��_n��`ӽ%�q ��/^J>}R�1�@�wt�l���yx���Ţ��F�9l��l'N��oW��:��=���q4fe]E����ն��~�8�8�!e(��M�\Xٖ����5�D9e!QE1P����Ps�ɬ�q�޻W�ZH{��P�0�Wb���5�q�ȸ��9�YcE���oi����Z� vb����1��f<.�EÝDu:�ϿZ�+��T���;�D%�!�E}�/�Лu���迕~�Zz�Tg�a?��?aι�C�6O.�l��4�]]�7��y�O���=,)8��Q��W%�����5�����ey�S��|v�b��7�՘��ƻ�J����B����ܸ�]E_>��k�\����?\ء�-_\�����D����ӷ�v�(�ܹ����Ԩ�ONG�L׋؆�BێkD �T��;�ʒ�Xwі�Ϲ\�����z��zh�������'���pOt���4��c����Κ8>�-��7F#_������L�x��P.��m�e�gc�3z*�T1kKS�K�T<O�fxU��I��:���|���S�l�k�L�:D�c/����0�/��P�o�s��m����˵q�"U\!I�f�mC>��u�<S.~�%>٤r����:��-W�����L��i;�q3��$V�&�����u��Cϴ����LS��)����B���ٻ���	���sϚ�B�y�c�x���B`\��Ϟ���.�o�&�V��o<l�\��ύ������(K�E׫Ϊ&k36�ű8w��g<�^�k���Gb�o$�ذf,�r\EICH맩+�4��>[\.S�V�7w��.��'J��;z<�u5��XI�S#b0�s�W�n��]�J�;���;l��M��H�>�2���a�q��jfކ_[��f�]��~<�}Q��֗[�t{�8��*T8�Y�	��w8��7^���Y��.p��z{5_���.<D:��lL� LAs�UT�>�(9��[�ڑ��Jz2,��L��V4�X㪠u��i}�C���</�^�s#dK�q�H���8ij�Ϫ�2�I���4�}5�����V�k�����[�F5���z�����D1΀ͥ���:2"};8^��>�x'[0h9�YM`��Dm�TZ��b�<��9.)��LאVG��rv��?��H��Xh�~�e?X�E�n
��_��bؤ����,��m�8�$6��r�hO]0��h�X���k���tA��vXuc�gP�9�}$��Sn���uP"�g��W�Ϡj�k^ɃQ=�����q�3���U�2>�Dg��[(�>x���֪(�j��孤4�s���Cr<�9Jb͏����>���$����*����%�"�VZ�L4��*��{��?x���-`�'�U�6ި5��>��(���P_O����_y�\]��2j���'0�wkknr�r����*#�M�\�i��� �D��A8Tjn�u^`o$���V���b֤{�؅)��ϣ�[���L!ike��#b�gT]ϒPݡXv�)���1H�a�(��+�����;7�ys��� �f����9���6���W%e�|�Em`�l톱��rS��j�Qr��:'W��K-��[��{c̜a �����.�)�������mN�U!?G�7�K!�[��6w@|Ƒ{�)�K���[eG[��l���m̥�5���\W����{���[����QN'�(�	��Ť<�E�yRS�W6n5�'��[��_�l��da��+'5ɛB�x���~u3<t/����d{/�܏�{آ(��ڈ%�]9-�������w�F�W]��́��|2�����h|��`�$�1�FxA%��UCkq��mHSQ��L>�*�uɓ�����9���
O��G|��Ev�Lh,����ʀ�s��'"�[�nj&|����5���Μ�Z�*I��ܵ#��0&�Z���.Ɓd>Hi�ށC��*Lf�z�~�onԙə���0��򕧙�����V��pȌ�I���hr�8;k�ۍk;j�0�z�DEOm���՛	
3^�����`����.�OP�PW�>V>n�dgM�&H2�Xw零��U����N�u�fO�x�3�=��L����3u��m{������Yk�;ZZ�Z��|>Q���wR1�H�u�s�xB��o�e���ݚ36wy�5��]�-]���
���j	=g>/`Z����O�0)։Ա���[�<:�sn.I�<l:"ky;N[��wW3�Kt��s�ꯨN�h���O?����ce��@yD��g 9��(kEz{�`Jzs/�e~�0����1�5*�����͛3]��ܽ�,�����j#�jY\Q:ј�4rae��)���L	*�dA��5�Ef��O�q���̦�Ҿ��C.5�"+���qDߍz1�ʑt#$SZ��[�/4��	��c��x�}�o��M"�KW�!��E�k��"�,�} ]��5�IWzn�]��7j]�q�閉�|4gٞ���9ҙl�ѯ�l�1#7���ߝVD��o�J�q;���'�2��p$�v�~���sN��0�K��ӓ�Uرe뀈j93Su�l.`[v���������3�~g��%��Z((��׀���_�{�lH���5�5	�1R�'��"� ������-[�%�C�'����񳿚����Q��{�\�L[ܸ��~�/6��?6��]��v+ѱ��	[`ߦ;�y�Xc2��t��z�i`z
�E�Vg;��=^jE5}=F^�Bh/�H��8ק�4[�Pܖwv��`���������_����z�����������a/����ĳ�2�f|ѯiN��^��S?��Y�嫙�3[æ�"ᙒ�e���*����p#;���-0�<L:�#n�ob|:"2��ȋ��%�V.ݫS(޾�G{�.N�P
A��{I�~v�k�2N1���Or�:��NRGLb�nJ.�؃�R�\��ࡑe!vff�Gq��1|�X�i�9 �Ē�3ZR�8��.��b�
��+w���Ô�)��$��䴏�w<�*�ϯه
Sq@v�d�X��1�R�!���uszl��hw:K[W%,�;bS��+Vd�������XD�f�ys,����G��+g��)(�/Q1'��9Tyn�� o�`��b�b"�c�$�e�=~�S^���P��o+��[�A��n�^v� �����31�w4tZ9�n7��vp��lw��)\ZX��#�SP�s�s:��ʽd��˚��7�Ha��,غV����	htB�kgV�/��^�W+��8����]�������=���s������K�Q�?k�A��pS+�VYa^�H[�/2��wv��J���:\틎��|��9�w����:�Wp��[�����(\�`������ƴU=�`\��O���І�K�(Jy��̷[��Zs{��m�9�E�M.�P��'���B�ms�=���&Y���h8�eNa�I���\,J�$��iUa��f�l�k�u�v&:e�0�Ds7���ף�㵉�Y��;����E�j�͗�MT��X�1r%{5���]��-d,�Od�w��\l)L�ٕ�M��{�[�\�>���.6��e[������ lO-���������Ѕ�j��u�Y��핫7o�v�p=���ؑ[D�����M^<}[	H�g����0�$�%��!$+��p��ކ���wG��tb=�|��8��M�X�J�u{�R� �-���Y�0�����nQs]�Z�+Z�Z��JY��]�Y��(_b�r��Ē�F�+BH.ͤv��іO;&^er�U"!��:f.KQ:6Pn��ӕ�p�Ķ�h�λv�[�t�v��cyM���NvTʰ�.��(����b��pOQT�W��{9!�S���%����Ʈ�QF�4iҖ�|f�!��mG� t����J��f�d��{eg`��gt[�2��4�� ���lču�4)A�u�rl1/��R������鯶��YmL�*��2X��/7��xh�^]v�L�1����^�L��6l��T���^1�+�;g��¹,��2�5���'*���q������!ɻC��3E$��Wk�Jܺ��%����,Z�'Z��0&��㐷��근���R���U+90Ҋn�E���~s
fc.j6��wCݵ�{��ʵ
ͳW���F,�N:���*(�os9a�D!w\����Cb�m��rsU��9�������w1]����^q� 5����Hb�@%%��-f��G��9��t�d�kZ�y|�o[03LFk��_���Uh몈��C�ݨ�
��uG=���[:H����j�(�.�6�v3��խ[N.�=jڵ���Cg�Ӊ�g�h��6hѪtDkWں��DTt��kX����ݎ���
鱳b��-%<��k5�:�5��.i�m�EJN���Gvi���4Wl���v�:+�XѶ+��xcq��1���`1Ӡ�1��Fj(�֊֌i��δFƓ1�;��E�u�F"�9΃�i�Th-���DN�����B�X֚4�ێ�H�KUl����S��4��j[�I�T�GlM�QWg�:g����"b�J�N�wv�[V��-Mڎ"�O]mmx>�%�n����(����+؟��}e����pW���9�.+�2Z��[��%"�7)�ײ�g>�|#r��n�lP�.Q&=�X靹��f�?�%DF�"�:�Y��y��{y�u�*���o,|�k��hVI�����\3���4.�J��lS����Ϟ�5�^;��\ ����57�v2���;�K.���K�!.;V='~�#�����lhcP��*MV����#+m�a���[y�-@�<H��H��O�E}E��#�X�`����m���B�d+�ۗ���������ˊ1Ba?4G��j`�a|�/���`�}�����v����w�(C7�ʱ��=��N�Ӟ%G:a��SQ�����1�3�:��2!>��"�ۓգ.�˒�;ܨ�m���`/=Y��@f�A��3k׹�b�]��\��~澓Zk�~�����v;����w�?qtW�X�a�^:T/O�9/~~~��t��若��5�����y���j�X�8��_�L?T%8�P�Z7&�\gz��Η�_n:�{�P���!��aF�[�0��
u���K�.-I��(��OŚ%]ϙ5�Wb����)��y���N�܉��˦��w��z��Un������C���޽6ӍR��$[�j�:Ŷ:@4[ޚڵ���Ŝ���W�=���m+A?��P�;V,pUec�'t��4��h���%��;y���:2ܴli[]���J2w3鼳�Y�2M��	-=%���a���9�z�,�ғ�e`�{���wi��rTg��fU��Cn[7����a�S"�:������o�]�~ ��v�����>D��b����$4�մTa�a
711�tp��3��ݠC���0P]�!�sՠ̳�V��>��N��L���m#t7|$�d�q�Q��_Ia����y�Tsx�oOT.������N��?g<�2�jS�.>th��(Z�aF�7��>Es�5���iw���]wo�n(�U0|{ư��O"��q^9j���d�Lc�r�{g�D ������6�}^ƈ,��&Ų�	��-Bd�cb�������R����3:� ���ǽ}�����b�]�[��7ʾD%��+�����	��u�l�:KzI�Vcv����騬�/Lԗi�����y�w�!ӟ����w� z����A���)��{>�Y�l��I���ϔ3b�{��59���k[��\^*�<k��Ϩs�c)�à'kՅ�n�?I�{Sl��Q�8m��Lަ�C�Rgu�XwY����� %t��1R��D����ȳ�l�N�{�kgm���Q����/�e>=ɮC�]��}伽�'�����{�d;�ti�����5?���l�P�2�#�'���|p�0��o1㵜_��h�BI��=����궶�u�-ݥ6mhӹ#�W_<�ư��H��:V�]�Y�;��a���oZٹf��[�{����N;�:�8�a�27B�̕U�8��@����,/�{�{��ǽ殓��>�w�߇��0���1R���<=CvCf�������;Q�*+��o#%�w,@&8���tUFwyq�0]������%Ih���`��<0��Wx�~�UM�xDB~���S��"�C��Jmz$k���P���LV��l$/��t����"�P��k���q�NU:�׃;�g;'�0�T\��_Sf�y��*d�d��<Na��e忾!�	��C�O\���/d0-��)n�Cu���Xs�eZUSs�(�~����|��c;�:��q��#��"�Y�!��cӃ`d_��
�i�ۘ�兀�Jn�E^1��u����0�eN���oJ���C^8��M/�G'��p�=|ZC�x�.,�E<:�'">���_��,ƪ�͙7��cWlu��T~��T����B���Q�i�������r�o&$F��\��g7.�ac87i޽��|�W���}88(��L�6F
�P�~��b7�ލ���x�d�2#lյ^a	F����̆t�䣛����?}��;@y�w�Lh/�3�)�|\<����x�	���Q�<�tnMD�?r��j��u�w͸�7���m��K,wݪa:��	ٔ�*��7eH��뜢�V���=�i��U�m�k���+�+��ɸ�$�Uyeɕf2�}0c�j��U�%�5\�]�㻫��dWY�,r������6G��_x�xxxmf"�*���u�m��Q�k���b�-B�z�Ɉ��-��h��O�Ɩz�d-��?zR�]7���}H~������*��ӽ�x%��X�&Ϧ�]�BO�#O�k��3U�q�
U����}L_3��+�Ks
�9�F��=C�21��t��z� Q}ŷk��ϺSś�Z�"�2Gr��?K'ҲKT�£u����mh�9N�c�����yj|�K�g�Vz�*!7k�Jq�W�z�O��D� ��|dK>gԧ�#���%��ڸ���l�e��{R3�Fc"_��]�,>F`�;Rʎ(�h�V��4�Q��I����߲~c���T�]�˛t"��w�fz<�e7�H��VӰ��."9�����1��T��k��1�]��3����j@L�������*ְ3�MV�Y6�+nۖEǞw)2+�09��5���],�â�zv꺎6&FAw�vj� �^)�5��t�_�)�^:�5D7Y��4}ǡ�y'n���걡�_ݲC�~;�Dؖ��82��=Х�Uw>%��i�
m�-�"�_pmɖ]z��Ķ`�{z�x��&݇�o%\�2�u�՗Idt���
�W�þ�'��|����yb��%KkpV㘈�Ӯq��(퓮��������6ܮ;�P����GC��tX3�ޛ+��KJ�lu��)�q	�A�.g�ȵ���}UU��W�_|$N���c!U�V1�����g�1�U�5�%��v=�����`��H��h^O_gRWۜ��<^��������9�P1P����� �Khu�YBO@��&pǔQ��E@�Qg~�ƾ�K�eP�4��>���8�!���PQ�t�^?r0��٠���`s�����[ Լw;͐ь�%L��:
b�-�UH��gz��⃎���r�䌖[��gб���1��f#C4`ލ��'�1M��L��/^�L���"������昍�<)��S�sQ�|g���P��߄E�~�Z�P��hm��!�MB\v�c�w�2;|_�>1��P�'�"�̃��q:_vw�/�]��x�x�M����O؍����ud���[C��]�?<�C8���T��5�˾�c]&�\Q�^Fs�����a��*�����NR�H���ffE4y��m\��M��
퀂��)|=7���P���^�BY\h����� Y��M#�⥿��X�\���>�޳!���z�?b�^Pϸ��e��F�' �n����k:���ĥ�����H�wj��/_��qd�}i��V�S"���e⨶�T�O[��Tq��d���=Q��X�NB�F�	�(5	����w�@_�轅@w]�}��8T5�hJ��N��ej��.�	�y�l���G���_�P�����'��c"����qmWp>�x�����������(Z�ՒM}ήL�:Gz/j2�L�׻OjL��}r��8���_�:ݽ>��a>¥k�΄AQnS;mⅵ��l��nL�Y<J��y������ڙ��[³�?����U|�eN�Sϑ0,���9،�t�Jj���xոL��r+	���Z�a��#^����VE�1c� _�Z��Ӟ�L\ɴ�������z���"0�/�ț�b��@fP�嵳���qm#"�JM�!�e���¶`l|�:�ٙ�ۆ��Xd2Ԇm=�3):��2���߫�e��=1�\r�&��B;�:�jy���zFuu�43��>���5�;Y�5�i0�jS�C����B��
8I"+��^cƬa�rX�V��{����4Zqy�����iGq^9j�����K�0Ϊ���l�ܶ��cҳ��u������`�G�*d}����~��]?{��5	G6���{�Y�2.�ځ���'�(]�Q��>O�"���>w�1	{S����yP����N�ӧW��m��w�b-İU_�U��ɣ���(����m�7M�l���=�C�a�L.��C�Y��a/z������'Vm�*�4*���vV�V�Jj}���5��⿦xT��ǽu9�,{� ������K�5��Cp�}˝�#�k��ľF]��(]������M釾$��o~O��R�b��-�2��^��`;��ҏz�Ɩ �л���m��\ea��4�����s��(1�O^&��^���>P6}_��'|�G��z���f��j�`�;�^�\QX���ck��-�=1��zb��T`*c=*���h>�!�nOM"�j�;�޺���ڃuH��љ�𭣨�����.�ϙ���H"|T��ѓϮ�D�[q&���H�����~ã�[Y)߱������g��Sr�j��@fސ��ϷG��ö����]29�s�SC+�|ͅ�m{�FU
�_N7v4=�����l�v�?؝ǟ��п��G�\�B�z�T%�ɯ��pQ6,TuaI�@�s�=W���W���7
K�/Kŗ�NV6�O��.�����]�Y�=S&������P��:ąP��tj�2}q��J~�p'��Q� L'��)��J��s��ۨZ��4 r�3�)�����-�[�z���{i�k�7s��!��Hw�+���NXXJ�����ۯi�d��y��8��,�2����hU\���Ճ�[��j�ǧ�� �p#��`�
���k��Fv��F%�t�f�c8��x^�J�_XQ�O��|;�mO=SQ��
���1[k��۟(d`i��2���{l�7cu�>`qN^DsK"���kH�� ���M����W����Ś�܈��Dt���z�����M���q`Ғ��E��;�{ɥ��s�j[P&N�5ɀ�=z�t����b"�P����xc�Ԯ'��KȈu ���B�f\\�����fL��|_�=X�{Gj�U9�2�cX���C̮#?6�;�*�mH�g�z(raL���c��~�en1�	��c���
-j�m���'���=�WT�˒;b��bز�u���u���	yd�6oz�t����W}_���Ui���}�{�O��:�T:܊���*����
���\�+�#�~��rCN�d=����+�b��^�q�hr�X���`��sE�1��jy�l�k��������y�G�o�:�.gXs1{.�OP��*F@��mxV��+�y�Z�kt"_�"����8?`��ˋ*1����>�;Nݸɫ1U��$��nvm4ҜB��$X��6\=���
8�: # _��0�N^O�Ʊs�ǧ�ye1�K�g'd4�N�T3~�@F
�������
'�'r!1g���Q�_G �ic�����0�Gm�[zi�J��If�[S$���d%4;�#���r�F�4R�K�+L�Gw����c���A�����Yb�L�nW<ySv����.���,c���q����jd.6�Aq7;f_ԉ#����? /��Mi�E��Gl����I�,�?z�:#�ϷҿR�1�����SyHeƽDEc����(�/B1�:�]��!�6���ؕ�hR��Mu0;^}sR{TJ^��4�Mi�f��Ho�V���L�8�'�@(LP{�0�_�-�4m3�:�Na�}1���{�):���#B۬�{�y9y�?;�����7��a�x/ݷ��SǀWU�#Wٵ�+������=M>4F�H�tLg��0X�vn<G{f+5l1���z@�VPw�a0SO��a�ꋞoyFk��27��G��H�vW�v�[!�R��_7�R<�RYClI���W`-���?�P����{��^��%z��<z��_`���*�Ձw]?:	�ڠ��7^�Gh����|�Z��j<X[9Q語"h��=����.(��R'�o��n�_�˔�^����p9�@x%�g	�;S�H1�x?o����l��
����C}/�Q�-��l�ށ9�yZaٱ͉�ֶ|�D�s)��]��s�n���� q�`zx��q�c3�I�GQ��\�'Q�m�N4wg������z��Y�r�-�*�T Ìl�tuq���Õt�C�­r_\Գ~�8��Yb�:u�Wqz{��'�<�:���Xv��N�.wl�0m���x���U�f<����Z�JVv)����.����U���*��f�xޝ�x�"��Y닎���?|&��^�_ʼ�<_�����Y���sY�;ܰ.ԣ���a�{�z��7H���V�\���y�=58\�����5���<���W+?�l@�>���T�Es�Ǔ�;o�WO���#y���������H
7t���ʎ4N���3��p��S��`ϩ�h�But_�S��8��3Y�fMH���~`a�u��胜�����>�ޮ|s-v�R�{�r���ت5��;u���kDޞ��;Ϡj��w7$�����K�w�'�9�����rd<Rx���:��&o�1��j���������~����ь�F������EFj� ˹��g>k �7*d��� N��~�=4JN|�eN��2����b3��;�x7�^&s	i�����܊��U��ޥ�B�P��X�N��`T|����(K��8]�w�!�����`}��NfQs�)�&�+�j�F��-���}w��nd��ԕ9RwL�T�ȏ%
�iއ�p5��E�uj��c(��!V^)��J=�)��$�n�\?3�～oG�����z�~�W��<|�|�?���޷���,z�4�{F؄�yE}(� b�w5���Dۖ�oH͡/0Y᛹&�����&�;pΠ��⣹��[ڱ7��;q0l���o�$o	oiJ
���\/]#���`�u�����q�8�.ӕ�,�f���2���7�$үa���Dr���!{�6��ڔ�B�^�L�*��qP�OR��k����Mi]��ҳ�:��m]g8�|i����׻݆��fZD.2����`��F�6��*����8��eiIμ���If���s\��z�d��{-�t&˳�%j��lh�o���NW��,�V�����C��wƏ[Gy��^)�l9��ڈ1wx��]x���f��-��\DU��:����Fq��J��Y%)j�p�F-��1�4��=4�qd�~ ���W]VF�}��Sm�U���ѼF�L̽�?��St��7���R;��g�U�_�/����^��酞�GUq��1ë9<�[�a�"��y���]��[��Nc�� �ݼ.$����H���17۫�M>3�[�B'$b�%L:X�͹�I�M=l��3�����<��Z� Ե{\B�����ܕ
+�Ւ(H����4�ֹFy6,�5I�߰K���;6�]F�ۼg~�[��3������%�H��e�\�H��U�t���]�lb��nD�M�ޑB����
�A�&����m�ff��~u��n�1��WrՑB�+P'Auc`D:"kc.�$,���B�ϬM*�v]��i[t�\�x�x�<{�ͮպi)x��,
�z;a=s����O��u���ri�
�;��:�v��#`-�ubNi���}��FAv�v�d ���o+!{t9�k�:�.W`2���YL�-�Vv;��Ԧ�x��,ޘ�!����iy�l�e8zX������#�Ѡ��^K�;��@��"��}�Ԝ{F��ƞ����"W���,Z��z����(��r{�)-�L�8˽�']����K�顂�KC�ku.�w7qw*jB�1�q���� U�?#�BU<�+k+y��tB_V�V(7o����ʻ"��drT�c��L.K{�$��7�X��ѧmY��ڜV�Ov�T���:I��c�9A*eLX2���H�G4����S���g��b\Ye��w5>`�b��W�4��`�W"o�q�wR�y8M�jv����Du4��&��3S�:h!�� δҲSy��|l�����8ګ�zᣉ͡M5Jξ�Q�"���<�������m�bT��qt���i�:������]�	��z���v�y=���b�}�`k} z��n]�l��]�3=�	=�0�{\q�ʶ\�/%�k~73���G��l[Q����G��9z��c4o䲸���.�˳�W�ϛ�4���`c%�]���=;�I�Ľzk,@~�"�e�C?�,�	��m��L��!�/Gm����j'�*��i۷EE;����ZѴcu���X�m`��涵j�Q�ێ�zFۼ熻 �fӊ`���Z:"Ekm�b������.ѱlQ]%q&'ct��j�v�q�]���s�6�!*�`�Ѯ�Y�$�5�I��u����(���էA��d�5Tv��F�l�z-�ݬLF�{��:|�SF�э�����-h:֩�s��Zz:����v��kwgwq�Z�4D���E�D��A���I��="&��4;ck�ph5[��EQlu��;1�.�c�%Qӱ��
횊j(�Q����vΩ棭=QN��X��Қ�&{���T�v��c�s�U�KY9��Q�>��}u�h��o�=܊�U�>w�.��~�0����2R��yZ�V����EEζ��j����&��"bO}��m����K�ay#���0��e0�kj���}N��Q�τ��;<���V��	%���gQFX��Lxw��\o����F�_��<���ɖ�*nP��8I^;�l���#�֬��ZA1�Q������9Q���B�Ê�7��e�.�|�!�K���蓙�%�_Kſ:��z,V�D�c~ ��x�����E2�8$%wb�w'�&�)��B
ޱ�
5��+|j���q�h/^.��϶$3��8!0~�ޜO�,��i�\��0��6%�$��otz�㊅���T'�x���~�	�(w;v���[��T}ⲻ���۰�Z���Y����g�Lf���j��\O�`�Ѡ�XPzu���[�p�j��b��\H��)��\nfK���.��܆��$`� �l9��p!]Bͻ^�ϰ�x�\���~n�E�������0e��ڦ�ۚ}~ ������Y90�R�j꾥���bS���$����ؙ�;♰}��*x��� �(��~Pm���Y�.h,��η5;�k49a8�뜩��h���E%����XeWlFr�eSį:ɖZn�N�����EwB�YC+tm�Ps��nΤ���7n���99��?�;Y#8;�~��4�m�ӷ9S��r뛬�ߒV�f�ے�^�m��� <>o�<m�X�-�Z�;b|'�o�C�bl����N$�6},�hu}T��\��t��4wIvױ��ͷr�O��Yj�X��+2��1�5��%�D�y��g�I����w|lG���'eF��l�<g�;�����A��5ՎQo^s�S���z�֕I~�!N�k7����tF)��y�6l=�;U�{�0��Jn��+�����v�(��i�m;��m|>B�Bݕ�:rp�1����
Ƿ�"�b��9WmIL���v�b���UK�/n��6���	�C;k�L��DD��x�=�4=Q}��}�ґ��E�kk�޸�"����Q�8H�z����x�4�B�H< ���9{�`��;�b�Sܩ>½�pA���Rɍ�
�n�Ae�P�m�x<�����e��L�=ro��1<�r)�/�}H.��"�>����V��*�y-�Cܻ0����<��O2j�1Ll�m~A�@y��QY�_�W�_1�9���� q�v3��{&h,��B5$_$�O����s��
�&Wy2�2%��v�L�y{ha�͕�a���z���g=-:>��R�`{�v��T��p���yl֐$ծ�6N�V����Ƿ�f��Fk�Z�Ek��Rɧ�=�J;}�OL�7i�w��w����,u�ayfKC�W��Y���U_}�W�_h~]��g�i$a�� �Z���6�'G/P��HQ��v�27�X ����0N�f�o�!��q��r%wF���q��x��t#RG;'�����4"�~[�׶=�W����3ȭ�y��tݧ�Q+�t�r�~����d`�����̳�I����̯�NggIꥌCܙ��Q渝PqV!�b���`S.ls�#��3��g��u�1Zh��V%��>��i���4��Bj=w^�X��\�ɐ�8�^J��y$E�ϫ�Ǭx._ Я#Z�n&W"�ѐj:P���>�U�}���K��fC�?bCm�Z,�8�bO���\dKή��I�Xᑉw����;�˄�f�3�G}�S/{��sl�����
 D�{tfݮ��z���&�(z�6�1≱>rF��|�.�O�5����-��F�C��(��z/ݜh^���5��ܙzc�t<c)��>��4����G��Rڜ����?����E�fQaDQ|�J��Khu�V�lKW�M�ɸ�p|�.z��{T������p`�ȍqy�����I<W�龗�nbQT�suL�h
�G�1����.8�ƨ�j�wL�]�Q8�лސ�"}�N�	u�9c72o�4]f�C��K!T	�3)�W{��)*Uk%c���xhF�U����_=���^��}�J����z���@�J��r���(�#:57���Lq&~Dh�ye��w�^}�H�3��ﱕ�% �=��\�ʝ�a�.r�4�K���g��Z�n��Q�\u�b�9��=#��;>����o����O�~.���}:h^�*m�n)��B6�~+����t��|���Zt=�d���GS	Y,�Ҡ+��Ј_)k����6��ӅƎ��Ѩ���,gq����H�3��Sv�zC�j���b�?5�pŧ����]�F�G�&�%�9��bW|��v�����B�};�cS�����w��.�^B���W�K}I���_0�z�wqm�;�7ѫˋs�M��2 ��Pͧdݻ�w�}�taw�,�|��
=2���8�;�f+OC�y��}W�-�J��_er�=%����Z���s��r{�s�4��q8���Ϊ��H�k��o*�Z�^a�i�<�vX��^��[P���=��_[�t����QB�%+8j���3Y&���k�%�MP�k�Q9����ߕ7D�C�d�z�ɡܼ=�t�O�N㷶�L&c���߅���s�����wH���z��9��S�t��5�^ڮne���#0e�����K��!~���꜖ӆ�{�F��N���҆L���Td�M��{k;��]˩7s��ӲR!�(��!$��ŵ��Y��	��a�[���
F��هE<W����;M\ ;�� ?��=�=�{����+*���Pf
�F\��+l_(���W1=P�����m�&z�K�>f���Z�5Y�c��e�4C���bZYgF��a�O׋(^߁U����ڈ���H|�a|"�}��_Q�2�n���׆\�lM���ۭOW����\�����x�^=k2�߇-�׬:LP�s�����Jкh+�WW���/��u�@���1کC߇L$���)�?bS�G,l��!��d�o����B�����<G�whO������I�jS��U)�����eߪy����K�U��{�NN�&��,~Dg�`��<��]Լ|�yk����O)d*��۹������}�YZk���Ha,���ޮ-�|�����l[��QRy[V���y�ݴ�5{$Ê\MBzY�2�RYy�>����#Whlh`� ��|��	�����tx��H]�q�y���7������W�G5���Mw��Cȃމ����,1�����{9���ak�y�!�#�{U�Q1z�Ʒ&y��dԖ�&�Ψ ���n�7�}u)^���\i��{���(�#M:�Ǵ�MQ#�#��"�h�o.�Eu_iɤ�o6��7g��e�j�AkI���.c��fn�����k݁d��	y��������)[W�j.��!�ʷ�QSK|ѩ��}����������7��f  'gT������l�,�xi�=C���\�CH�������%R����Dg5N��k��&�(ĳ�U�lΑ'�<�����ڎ��/)�Wy.T<߁�Ѵx䱷gc��Dss�8�:T��t_�ꉯ�]�?�5~����g|���&��{�3N�f���I���6%�p��Cb�$M�]Y}��H�l,de�>f���r�pG���뮣s.q_A{v}6�S�9�4^w���n��57jx&+~Ǌd���2�E�	���,q>�ѫ����'f;����y�U�	�3
ldw:���c�f�y�\]��Tɱ��9�7�=�[��vJy^ۮ�vY:4��_����hGD��	�pJ��s�k~�蛌G���~�YQ�wh\M9�6�VQ�lcq/S�oL��ȇ�ן[��,�A��*�{s��K�R[�u:x�N_�.c��7Wv�-k�����1�5�,�[���GN~�Ǩc���ƿK��z��6�i@��[�>W�๻:=ǆ��=<%��zaj�g�A%��F����L�ؓ{�"5ra�D�tmuzv�u���FF8˲���C���J�}����{7**ro�8�����\����cv�b˞�N3-.U���+C�nT�����GańT����'���� ,���{o�����A�O?�k����D��ǫ������轾O�����
#����f�Ж��{��'~M�i�������P��F�=��]zT;]5�r^Z�g�
�P�D��n��z�g��9�Ѕ:�w>+l�uS*Β���e5!|�ce���r%υ=Do��`;U��p�G7،���k���_5_&`����֐6w����S��Ih�S�i&�Gxe��${��AՆs֩H3x�� !Dņw���2��9�
f�;�p��V�~�>�g��#'�����r�ط<�����ϵP���#�F�H�z|"�_p�����;c�y�v��F�1��C\_a`��7��1#կh��Q��}W�^n�djH�`L�/j}�ő������	G!
���?�՜�]W�M]�RmA����������n�=yw֐�#(�"��>d��ݪ�I7��C�k�v*�~�wuR�w�dMǝl\��O��j���8�u���i�v�ӄY�}�.��꾙�@�9��3G�W��X�/]/���g�xu��2�^�#S39w�^Wq�
��	���BͿuU�N��z\�E�ʄ-T�3_]*��e��Η�nh1��CD}��Q�3} (�
Z��Z��+��+�N�x��4y�����R��y�zۓ5P�`�YM:�3Ձԙ �M��A�FV7�ª��]7�{Ȑ������ڽ��x��;����T6_{�c9�%��|k�mL��+Qo�{y�����__t~�(�RH��=�.�⍋\����<5�cю��!���3ȑi�17�TyG��)�>��Gl��ʩ�v��
b{���e͘�L]����Q�%G���l(����33�K�,����c�;f�m��U�ۄ��s�Qi�����U�5������e�g�a"
i���O�;u�x�)�L�����@u�5�ۛ�C��T9�㻁*���Ҳ����}^h����|�O�;w�ON�ˍw�����$`�D�h�[� ��α�Ϲz��f�+�rd3��[�F�Q�F[5�ã�H��ᣟ���~��B���<��M%�%���u�@�Y�M$(I�֋�}��w�(�<�v�}<"��=���h�5Y��0����Q���	g�3�B�;���|�8v^�x��Gy`C�˻bX?6�>OB\n��I�Gq�؞���M��-�gč�d..	�"�k�>T��z���A��$N?�������P/�x#:	26�a���ɬui�.����V=�-��ܻ�2Xe3e�{Lب/c|�'���������uۯ��Y�����_�r�;�Z���}�:�hX��W�je#x��:��̱~��h���'�z��{޽/LM���-�Әz�߻9��ǋ���ɉ��e�v]�ޘ���\�]�A7z��]��hh9l�;��{'_��r����������˾}���^}?�?y()V���d��v&j)+W/��ܲ��s��=�j]`��%Cބ�0}�ύ7E����VE�m��7'��>��
��[p8'O���g�W�~���67_x�C�?� �̀������u�%N�d���*`�(��~=�펚��|����)bj펂��Kн�a�%6���T��J�C\t��z�xCb���6�d<5�}uQ�mR*�,��Q�� ��a�B�*mwX��x��w6yV�l����u�(<�B�u�(o��MDr�!82��������?�$X����o~���Gǌر�x{K��z��n3�nJ�DKƏޢ���Yxth�b���#�� � "s�wя8x� ���৩���7!�/�y�i��Tm�մV�U�m��	9�z�j���綎�v�HA���f�ܥ�̢�<���;��F�dG����3�o{�fS��὘||2���਒��(��Ff�7ҡ�2�H&�7'�+�:l�]��C;R0]����~������
��Dŭa_����ʦ�����	vyz�� 0���}n���P��E��*����p����6������t��Z�L$��i��U�u��{�6)���*��f���d�eoԾ��Rk��5S�ň���Η���y9��O`�M�����O�)���Ԙ�+�iM���m��T�v��v2s8o<�H�����=�3  �330�f y�xx3�WE�fWU1��|��oA>��>֬�<u�!��~zy���I��ح�q����MA�����:�#�yY��ޝOAdw8�),$-k>��H�ޣ$t|  ��]�Y˙ה	{�)YY�o`�L�#=���J�rc��Ƒ�LdPY�ff[[��Ar�n2k��,�;�!&�S��#�LM}q,X�r�b�k�@�kz�5��$Ԗ�b������^Z8+�해���/�h�=�O�rd�iaY�/~�4��l`_3ׁ0-��^r)�^���7N7�����f��~��ɕ���0_�p�+´�>�;���Id����_��^� �w��w�����@�hc����3Ì�Bz0�xm���SQf���]-��f�$���R}Vc�!�z|��}W8��O�I�_s�"+�H�#42���8|���Ud�T��{+b�K�f��ч���t�}JAeA+�X��EBQ���D�&Ō��ss�yepu=�����%:�V�����1ݹ��b��w(d��M1�=���U�cm��?>����}�g��}�g��?f}9��������Z���!Ȅ��^�`�;xmK�z0-2˽zY�:�7���c�|����C;*�Ē�pgς'������u�X̂���9
�M�i}7��Ǟ�˅k��V �CG]����hv��W	;}�HŃ*�n�-蹛2����K�1�U�.X6���0�L��qgs�/��L� t����X�b�s��u�\��i�"q�%�mg]���@����8���L�3.��o>�ǯs�0�H��M��&�3x��Y�t����,xvW�ޫ6��e�T�����܏��j�q�]�X�Uv6gM�*�;؉"P�nd}.Fn�RrYo�(����N��`����¬��m��>�{Q�IӋ�c%�TS�w�nv,���'<=r����V���֧98����l��X�
bA��]��]S뤹���-��s�=������::v�Y��x�tM�gk)؃5�bc�6�N�o/��됫�gcѤ��f9EJX��T/c�����څ�:n�����ߓ�+-ࢩ�&�h;]7��<�U����mԱ�ْV�}g{.n�MZgr��
�9��K�!��:�ϖ��]O��F�dX���+7�5��#U��H(93*a�γ�+���ܻ�0N�Mn�b�t��*���˷>�]#V�j�AF.��
:�3*4�iy��o�au��2��%"��L�ڰv"D��C�̣�Zc���>�!WGy�4���Crm�1J���M���1t�3�����~�CG|��#�]x˼���w֍���42\����ٔ����D��zw&��1�����ѥ��(�E�M�ى;��%f�9�.X�Jݣɂ0Q��ZP�f��k�+K��;�N5\+:\!*��v�.�%Mݴ6�%�e3��g[�/P&�ysa�[[v`h�G�ڽW;��E��K��E2���(�AN�s�����ܺ�V���챙�����Q�U͓�n�2F���W��^�w�r����&]�Ԙkqd�
�v_,�|��/A$"O\��i%�.R�l�m���1�r����F�i�۬ub��gN���&ڀ����-t�q�mΝMEN���r�J=f��5�Rj�n1l���,+�h�[i<�E+����q+��V�V'�+iRƷV*m�rb��q�֥�V�����i���]udl蛡�c�ZJ��[�q�s��gt�%v�N�V4�kp=P���������{�m�c��d�#;ফ��0+w���Qc)"�$��+��Z�C�)f�Lg_:�ଓ)�9u��؇6�n��m�}Zײ�w���]%g,J����b��;�Z�4A[��.�/wk��Wp槎�WP���^�9���7�;&$ ���Q�ȸ��4R�lAq}��k��WW�l���@M.�>Y�$];SH�u;e��d itX��݀���l��ɩ��V��*�l|9�dF�k/%%ݽ�P���缭�珟A_$?AқcGlh�i����-iر�.�m��Ӣ��b�']D�]�F���F���G�j�cGl���"N�wdű���4th��:�����������ltT\svꠍ�q�4��b��vUE֩�u���EtU�Q���vm�h�PE���m'F���6"��Ww;`���V�,F�M�"b�[��q��d����n�[N.�ݎ�������fv�֪J��.�Ui(zz��w;w=�tj(��-��)���X�Z�UCMQ��ݳ;b
�����Rv�Tlh���X�[h��8��ӣX ��64M���Q��7n��%Q�U1DT��huv{���SV��]��1L�Nشb"�����**.�4豌�13E����"홪#�j"b�������P�7�{���V�!o�0�׼9���<:�W`�Ӹy�Ϲ���*�x�V�C^�4[�|��˶\a�ۮıq����<U�*�\{y��n�A?���ycu���#o:+��3U���JB4�@~ ������1ܺ�A� ��VZ��_(�e�����w��Ex�Ҙ~n�>=�uc�ٽV��)�
h&e�ٷ���T¼��N	���&|�1�h|z�،T��:~a�X���׌��pƇm��ݥ-������:�rMh�H���J�H�q]�,�bo�*�ﺹ��J8G��`�ta^�Yo�a��l�+��}<97OO�s�k�L-P�Ꙓ�N��F��8�nyhKE�<�lNXҀ�T����3b,x����;�V�;U~�� x��sI/`A�Υ��{�v�����EmwK������dg�����)T5,����Tsr��
HZ�.�F6�m�Т�~�ɜ��P��>�>a�y�M�-͞��V�J�/�Ih���5=�;��x��G����k�U�Ѹ;Jvġ�S�!�ƈE��<�J�)���t�[9����'���Fc,M�245���'&�>=R�髃��wf����!�
az��ls#�P�|�=CR����ss�kA�d�[Y��J��
'�~+�*���fH�_$1��9l�T{�����7����l�������#.R���Qu4V�[&<1SVf�ns���z�Ǯ����I����=6����rv��e`�Zq���:/�v{�lb�7�Η���|6h�s�M=��\�תngP�f7�r\X�_9G����.W��4�B%-	2L�`<0c��7+|)3o}�X����7Xc ���$X�T��7P����Z~&FT|d%C��� c�{"kv�O��/�ֽ���32�uv�ҩ�1�
����Q�Գ�-ux����Q>�?:�}hf:��
i����Sb�m�6Ez|/��x%If��-t5e;�P��T��| ���hW|�v_����Iw*k0�ǝE�ʄ-ELw��˨�����1le��I�=����j~PY۴������r���}5�l��x�G��`o�#t>��-l�Q�'��1��jex��\�����U�u�1I��M���{m["�����:J�=�Gk6p)�~G���ʯ�5Ɯ#�N?��8|`����F`�\��NNT/�Z�a�M���;˯3�0r�=���t�3e��>��k��c�d���!}���;�Qk "�����o�"��dۑm>�r��no�V�k_��wZ^��b���,Z����Y�q��E�e�a���BGly�g%���N��;{ϫ_�8����c�W�2��}�B�����Q��&^��\���6釲��7F��������X��s�]�d�X���ϡ�g[�Jo:���mڽ{����+}�އ#3�[e*��ޥ�]`���Y���\{���d,�&oI���g����[OWrU"�5:һ�ݹ.}��垾%<vBH�V[+����|@��)Kwڻ�\b����X
Ĉ�4z��=�/�������ϹϽ�;Z)�lvm؍c�L��/<轊ؾz�2*�<�0���k��ȣ��"�����Zv|�\f���a����_��#O���Qc�Ҿr�6{lqX���Y�E�����1���`��P��M]�@�/"�8��H�ϧ���t4�ש�=������%;��-nkhw��w�L��3e�x�0^�<��wIo�5W{L���5d���G�4?_�"E���3�T�(�Z��|PP3�n��%��;'7«�Y��3�旡A�7�?��� q�~]��_�F{H����g�>_�w��>��!�N��o�TF:�v�3����f����i��X#�k�g���W_f�D����%_�W���E9"Lf��hyu9�05��P���d��<��}~���L��f�ЃL>�K�UϜ�!�9𽼗�/�=�i�n�+5���Ǖ2f8A��n�1xw��6��+b�s�#j��K��ʉ��#�,>6�3���Q{���1w�܈Q�6-�D=�;��4/�_����PΆ�����&K����O���S!�wִ�K��v(��T`$�/xF�ϱkͫ:F�-�{͆�;3gVB����0G�o��l�B�����Eʁm>�ۜ8��i��%�b����O٪��{�K�=����>��P�@Ƿǯ^�y�n��+o��3���hƵ�\t�-a��/���`aX3�.�o+���Ik4�Q�(+�p__��a�Sܜ9z<y}�4�!�{����3(���/�럵)�v��d{f�a��ax}y����P�B<��>=ğ�q�=�Z�(=�P�y1�ySg3ԯf�g��%��6�t��t/Ǎ1���
\�j�Y_D�cu	�D��5���<�/�P������=HJ�ͭ&���2�殌���W�y��)�G ��ȝ i�O��W�D#sی�W��g�O<����z���M(q��Bz���|kJ	Z��\�;�1���������u�^v��7�j�u�v�^�U<˿������ĜT3�)1�a?3Ԛ��>6�Ǝ{�vކ�Ix�B��:��#v`��%��֛�p����ӌ���B��8���Z�Ԛ}ڳ��6/��ꨳ�o!CR�������fyTG�Oׅ��Ϧ���`;��/1�1�';r�a�>�Ǉ��wjq�k��
�����g=��B�d���A���_�#��'H��c'�sH�,^�o���Y�����P��3�憗.�k��^�GR k���JD��Iiv��zS�[Rr��J�!�RF>��f̒D~�z���r��ǰ.�.r�^�W1Y;���l�uH{h�}��}m�i��T���o �)�\�Q{7��ݽ�u��%���h �(�Yw��r>	$���w���]0��I����F��1BS�c����=�i/���.۹0�����SC/k�P��r:��V4��G4��p�+�g�l����Зu�E��4��D���S4���/��E16�<1�jە	E/�s��C�����Y�����7����)Ǧ���_x/�]`_w:��3L��*���+2�zπ���R��)ml��6�Չq�]����^&���p�h��d�-���S۷.{�y��n�dU�@g%���ᏽ�6nnc"�KR��4ܻe	��s�l�0􇞝V���F�����nl"�����B/j_�������K��`�>�_�f����4etK�&m��x�:������֮gn˂�Ws�1J�|���_�G7/��Ԣ�)�1]E?�-/_<�V�/t�.�ٜv�-�+��@w�؍�	p|�3p�}����v��ppQ�ę1�����U��,Oun�K�ޣ�����M�b�[g�qQkk��0�Q���ӱ����Z��Xz�'���^D��q��g>^�������ƅ������/▢�d�/z�A؎e�RHx��X�.7�b���;S\�/pНqS}�u*�*Yc:
�׺�v0��!R��'U�T��\QD�ۮbo_K�n�M4˾_kX�߼ 37��3�'~�^O*�O��1���@��w���ѳ�Hvskô���<��@���<p�N��]͒��W��T"4:�{�"��8)��{9A��rQ�27�w���s�4�f�t��ǥy�n�פ�Z5a��vМ��C��}�lt�0ڕk�H�"�]u� �֤a�˝�T;�C�,�t"m��|$U<�@EY�~JT��D���Pظ@k�%>���-C�˷W��2���"��f
ujY_gJ&����-A����w���'h�ޞ�.3��q��#ŷ3*��ۼi�((6�am�#���*,�)�k�dKIϹo^+�`,����������I�MG���l:��_/��A�^u�4����sG1��v�v[gꊻ���]|���m�+���Pp���(]��x�Ҩ�e���p�x^0i|�E�j�%���T�a-�k��Mi���;�7����D�~���kd%n�>O�_���6^:;덇�>���r���C[����:ѴsIn���J����~���%F~2˟Wh5n�g@�:�6���hn�{�զ���P��M'ƞaW������:Be��ͬ1�����][�ۧu9�?:�(PJ���co�����b}}�X���`�� �*���D�d�V[�rs<v>�>wķ)q0�/����u<�S7RК[���`=��y��{mU��i)ֆ?^N����\[�U��TZrsU�Sl5���ǲ��1����!�,8�-uɑ�'o���?��v΁��D[ͯfB*3"(�jR����Y"�F�8ĈGԊx{G�Ӌ�&p�D��r z��M#o�]�9L��r���ܺ#<ܬuE�m��k|�o9YW3����09��0X+�f��FH4��O=4`k�Q��F��ܦ�}�L�b�M���ٷ޳m����}e4��$����_>"?>���O?W�xм6��D�AO2#���E�-� �'��g�u�f���>3�}��_��h��@��|hD;<�w��#���sn�Gd󜷨�hrac�+�Sp9�2jz����v�"�8�+y#)�2�f,��cP�U*h���꽑���V9����1��z&y�9�.0�0^��.w�Uj���rak/�K����E�ɂ'��l��ϧG;�y�v�~=����&Gf�ҕ�i��{��gmv]�̝��=x�Oh��3�c����Z ɱ��A��2jE��x�,?|�1�[Y�ي�hc��Il�������"=���l ;㽮���i2p�w!�3�\d��������5�*o�5�Κ���q�����Ί`�mݡP��M!�E�Q���>GK"`��_:��u�X�,s�`]U:bD����uE���ލ���ɀ� o3U�pn�\q��\������}�n�G�TH��yyTk�k;lWg�3��o��+�%��]
:w��t; �U�D����~QP��:���z#�
�N�Y�/��@���U����o�]���*`����>���-�g[��͎kD �TɮRC�82���s~[�=����~��	K�S�N3�RGgc���{��^l{��+��G���f�*�Q��I�I��+E�����_pBZ�,V�Z|l>�E���/�G�q�lׯV�(i�,�L�Ԟ��,{�W�:\Zy!� �\;��\�]Y ���!�{�R���]XOϏ?\���1ȩ�%�����ۏ���ˍ��zt�_&�����P��ܧ�S�}%�>q���n�ٳ�S��֣������L{��Ώ:xaO�$�7g(�2�I�;�p���k�Et�+�n�����s���ڭa~D�d�9�a?w܄xWEjCIg��-\j�{�	\g)�����m;�j��_��80��F-�G0ŷ���z.���`Ɂ_g4�) �E���M�Ć���Z�>z�d�����2�Yh����slfa��]�T��6�i��W�'N\�5�ʬ���ֳ�i�{"�y�n+�L���J�q��W)kt@2r9y���Ԍ��`v���S�(��w��TUҕ�g�|G�Ā?{�0o{�ê���0n��mvfe��1���1s�b��O�z�z�I�cp��D����ScP��^`k���Xvq-�^{����@�;�/���F��G��'��F�0�8Ƶ=\�/�y.r�,6t�y��M��H��ꁳ�����O����k�)�aXVz_}Zk��h<�X�ǡ���_��u�P/zb����Z�sEj�_�A�L2��A͟3�F��������1H{�Twt;�����<N��ފ���k���f��N��h�[�Tw�6�8�F9���ze�\�8:�u!!tgW�Il��⢭C�Ƃ���D���PN]�P����0��x�s�����QӐ4+�����x���Hh���S�T1�w[�Xv"�����_`�7X6%���mz�g��d�pN��c�S1�ѓQ#�����C;��H>�k�G��kh�>/rj2w7V��/}�Tɫ8O��'0�ġb�O2m�!���5��»�S-�@�'�{M֢��:�8��-\�tSl���a@�̘/S*"N	�]��|pzE��A�%���$��t�no��;��:Cs ��:���+�`~g�+$�uò���>M�X��I:�����靚�T�W�;&��8��y�nW�tƖ�tS�K;�"����#��Yf
ӌ��f���K��8�2�ETǠuޅ5�W���0#���W��u��TAQ-0A?o�����2*�]�bu�	u�bt4�"��}�vn/ji����:k���=��'���J �C�1��BVb����༩���'ֵ���R���	P��?@��1��V�ܭ��){���;�w��HGK'��>�T����%O'!D�c�w���^\��l�`oN.�/N�z��\�φ~;�wߢ|w�Hw�x�Q~���s�sÞ�g�\��^�{.W��v��O�L�l}��{�D�c"����_�ι��}^�%�w2{��(��� �V�C��5-��ȏ��A����{�*�u��W��,�I�g�sDi��]�aL#��n�\\�n��<��N���BO��#O�QpXH��0 '���� �m�Ts����6��}�L���@�.gXs[���D��/ʼ�ȃ[G:�d�??{������t2��bW~A�kB���R���C6������;w3��>�$p��Ӈ���O�nom���˅���$y>��{��Y3��}y��jG�H�g��^{�ټ��cO��y����G����z�^�_��x����C�����l�wD���w�ȁ��ad�h͛FK�!7�^d���-7}�Zg4���Xiq�5��k�K+�7w�f��`U�e��ӥ(�闝��+����YQ���k��kf�[�DB<[X/5Į2���[��������P��cJ�zf��o_b&��>@�=�;#�;��E��p��K��������]�՟�L��(ôÂd�2��:���+� 	�B��c��c��zU �	�H��	�t%�R�(�+�^R����N_+�{m�E�ю�c�w��*��]j���F��Y˘1�y�ɚ�\�9ݻ�M����h��-�7�A�Vk��;k�=c��D�T:l���Zh���-n���6S;��^qߔd֪M�u�Xp�,#���򤂶�jӵغf���q9����7EQْ��X17Ҁ�J�Ac��"��
��e�ˎ��y����:5�U�r2ӫ땻VX��� �wk�}o���\�)F��|��l����a;�쭲̀p�@����`z��lR�4$P��&v;δoZkP3�d�P4���L9ۑ��+E�.�c9+����%H�/���Q<	�WE��z�N�$��j�yu�"�cs8���.0�) ��Q�k���w\�W+������Jl���cchh��Vl���G7u#T&#w�]��g[3c�6�XV�\�Ն^.#��KM�e�XA��&�އn���^��8v<�784H�XU��]����pKL ���%�Չ7>i1N�k���c���:ɢ�٭�zzn3y4��yQi7�s�ب�<�]�ג+q�w²��yl�S�����$��~����\dᥖ��G0 �2R96�L4TK�ŅQY
��.���m���w>�2�m���\�K�g_%�	m���4���$��m1��jѺ����/n�㩾�k�.�F�N����,����h�-ǋ2�`#-;��ng����E��0�����N�1%�jft���o�b��+o �tp��t���np�*S%�c(.<�Nu�,*�at��6+�(�3�U����R�n�l�N��:�v��B�n ��c�����s��F³�ȳa�N��˭U1!�gJF�n6G�c1V�de�ݑIo6vP��0�ُݍ}�2�U_V1�����PĔ/D\؏��di�ڛ��|�n��q�&ړM�}�p�XƁ�`mc� ���kr슙D(Ԗ��/j��vƽ��]^-(�B%���͞[�3Y�BNb�xL8�v �؋{��i���{�Ӌ����Z
��go�Ա�0p�B����9��Cw�[�W4�JbM�ތ�����Q�5��e��嵳s��'e�8΂K΀��;2�Ti�U�K���l�[6V�V�}���~uo���3X���EQ1u�cETTLF:��GcQ$EY��)���g�v�*�1h�m���Eэj�툩��Mf�jh�&��j���k����.����wbXc���3C=��M��h�b{h�b����"�)����4Tm��Fb���lUN"*��j��#���E5D�4D(�
(�F����h�'F"b��)�i��qUU]�K��t5��;b��b�������m�OZ���t���l�Hh�+��^�ff���1�����Si+Un��QpT�]�kG\]i"�j��kGA�:�QRm��(��"��"5�`�T1�3k4TlGGF6�DQm:f�1�;:�ƴ�Lv�h���"�����Z�SU�L�T:]DU3�Q�DQ;i����6��>�b^-�ŝy�H8�|�Ijt�^[��J�f�b�b�ηv��E�]�,o�UU�[�?����~ f��f`���{�,h���a?�zw�T����)��5r����+�q�O䧙���-jC�ݳ-�z=�!�O��l��Fa�����B&8�Ut���:�Oj��T���s��j��uCT}����eS����#�ݮ���񋘀�8��ŗ�x�t�^��ʍ����)9��E6����8���^IП�w�a��sS���'}Un��.p�Vȷ��L]�.o�QpΣ��Qi�f�֦�k99N��G����֫�w��9�n_O�W�.F��`M�"��n�2	��*\s��{�?eF��MH}�"MɎ2�;��˪Ӊ7��'<�2����p�C��w�!�)~,|�q�n���D�����K�vT��-ȓ��Hwv�\kd5Y]�E>]�&�}�hvzz.��¼ju�>l��BS۶�M:�L�Ϡ,��8IN@��W��W�k��β4�n��mnYt��9z���Qa���/�C���߼����~��:�����^0��{�#K�j�����7��>^�/dg'Bt�"�s=�u;m�yz�kJ�ם����k�KC��^2��E��Z��e��Z�x�g>���Sw��䇳X/xSK)�0$�->
a˅a�&oN�s]##�v��n�Y9wDx�
��(�����������`(���sׯ=}y���=�c�zO1��8��N3�Q��^Y�#(I�л�p'��@�H/Nd ����{�x���jaݛ.5��X��o�b`���cmށ3�1�Qq�1B`���M*:�L����1��j��0t��c�|�9b��|�F�O���7_��s�-a�(٭}�*OYǸ�3QNf�lE4b��ߩ15��O��?8����/ݙ�0�7c�8k��e�87g���rL�r���7�H�����ߜ����At��/X��t���B��֡U�q7���]״ƆP�A�<`CT��p�#��<K��|s^��ǘ�B"����I,"�C*6����u��ٶ;`�����96�3��*g��B�yS&����|'Z����)�˳5훾��~p\�)}��9'C��0w�f)3�	�lU�8��ab-C�aqR�[)ndK��*wӬ���Lyج
(�^J1�twQ�k�鄟m)�&�X�s��1���#&-�6�O������{lw�N ><1���/��i�R��s2�b>10ٹ�"ko�����y��N:ڲ��c���%����pa�@=����d-5�9U�����7��[sD��Nk,�Xc�#hd�])b[�3��YY�\�=�%:�Xk�"C�$�:�՝+��=s��gMu�\�b qI	���[Fi��Z��2�~���Y$	�$�ZO�o��_>|k��{�-�MR���!�7�-m�?���e�1|��ƹPm�|~�Qzr�ا����9�����wɘ�'��X+�X;�#ҩ����W�t��g�����7gE��,r��c�yN��r��mv��^�����׷SH��gQ�r�s�FK�W��l����qu�Z�����a���C���2�I�=>z��hWT�Ƒ�:����q���x.lj�]�q���2d2�S-
2�tR��ͮ�Й�.lTS)=E�I�C;��w����Hhԫ�`V� U�_�59uHz����Aޟ�S�@(v|��}Wc���w�p}+L(�O=S,t��fT.�"��ڃX���NԖ�&P��^aM}�ٞU�i��ߗ��ә.�h�ԍ���\:�:�vs��9æ/�����L(�T$����3��zbWҧ������]IPR�M�`�ͻ��f�[ �\!j-�rv/��H�$!)��%�>xt�몈���Xl�TM��3�tmˬ�՞���NFK�,��km�,��t7܄��]YG�]C	����b���������u�£o!k�^jӓ"�٧�N�M��Y��jӖmB�����;�v��z,�Ĳ�I��C���g�Y��6�]�xTY�υ���Gֵ&������H��m�#C�F^�N:�B�2Tbkɖ�ѤgvNc�N\��sU�� �0o �=�a����x�o	��3���V��9.YD��0�R�A��Z/}�'�5G�(Xn5�ES�S��ʹ�R�#�Ο^'2�aD�&Ł�P"��y�����x��>թ�k0���Q�y-�
v�A�\޽��0������s/V��Ml���� ���GD�3���u��������u�D�Z�TȹԦۈ̘D���1B񯭓������ܫ�p������d-�{��o���N��Ws�xNXpJ��v�z���I�&c �ީ��&Ķ$�C����f��46��?XTԁ,$&��y�Ob��Eֵ��QR���	P3ϟ�m�TS�n$�w0�����[��<S��q�/�;z{	�@�\�;��u#��э�{�!���Y��9��:�$�>8^nay!4�D6_����6W��n�s�����}I�{��T�ô�G������GA_�tyw� ��aQ����o^�u�����p�޵%�i���g�u�F|�05X�Z�۷̃��4z5���<�b�����w�#�V_���h�ϴD��|<|2��_Yn�b�=�+5n؛h��P���Z:�,u�$�o��PF�_#A��=\���#;vS���pToZ���lgnd��V�s:w�Z�'4��agb��຦G!�w6|��s��ϣ��������� �
 �h f���i>��7f!����?as>�g�z��q�h~b�ɈfМ��}�L�$���Q$Oh�UK6�Q�"������V�>̌mk�0��� �~%՛���� �8εf��0��4�eIn�T�$:�W��1��a=��$gq�v�c ��(�9�Ox����U�f�yL�a�#k�O"����&�����3wnᴘf��R�*��a���BVH%N��A�,[<7z䳺�T58/�T�Q���3�a�
ny�&��uq6�Aj��_d��Xu���������W����nZ�ƈ�T��T���|ǟ<��Q�L.qz��lM	\�����	ִǋ]�2���x�2m��!��բ�5�ɑQf�l\z�3&y|�S�����uйֳO�w?W��k;m�NWJe���)�_�����󭓡}�$4��"_�D��Xq�?U:&;�%t�uf������pGJ��`%��R+h)�Ĝ��he�y.^0,�j�ska;�����3W��<!&�?;���3@�N�Ӽ�����	�m����ydI�&x#)�:L��p{���]��!�a5�]"���U����P'N��K[/^�.�k��+�o�}QP;�Hw~V��Vt"���S�Z�«�z���([������L�����ͨ�y���$w|�(<k�P�8S�:p�h����>lq�f��}� ���3 �7�0f!M�i���l+����x4F8Pι�\�)��O�󢝨g)�&�@�\K���(-k=u=�����6�F|u�������@u�X�"ྞ_Wm��k��]��QQPr���]��&^<���J{,�<�}���kđ��X_>"?��6"���~ʘ[�K�[��d[N�R�w�<m���ጧ�_](��p^�8��F���b�������U�i7���S�J(c�y���_�3���F�5,��*�^�ňr��p����*��jA�,��]����וq�?�|��UٓM=������-�z鴴x�·0�_t��}{Ηܢ]Ԙ:��e�w�$:b�d�c}��/���;��z'�O4��J þ��&n�Q̼[����I�F�Ig�u>�D;=���1��Pʅ��-�鋨2�.���ׁ���0��D�j�<�I}���5&j��Й=�"�B�i����wf�BNt:wB&��:�2�����.��~���_\�9��3��E���*N���+���C�>��+��*��՝yhE�PޗԴ�����X�U� �lL�N���b���68��!a�GI��#մ��N��Z7J�Ղ���*��+uK�\pP2o��!|���8�nun;c�0�|������� ��g\ﯗ��oݲ+�)�&�Q��s�W):���A�=Z�O�X�m�Z!�OQ:]G��/�y{ �b�#zsRC��1�/��3���w*tr��0w�f�u������1eElt�F�3v�&�C.��y���3F4�d�"��)�s~�%��-|%O�*�bV���L	u��P��;�s(m�����jB���E��E�~��<�C4�)E�&ݹ����5�Ƚmu�H��/ɽ��T�i���3�1\��oB�gu$<*�w�4�$`��{�됎*9f�T��� �kXWL���9�'F�u×�*%Ή$a� � ���ҹ
����=S,_�)��u	}�רe�5�-���o`���I@�\x�%�3I�l��omm�_kڛ�����]�嗦as����ƅgJjޘNC��1�τt[��Lmxg\�5Y%[�ʃ��>�4���J'�"��c��W�-u���isb��Omu���WP�Jz.T{'��cg�J�0k3�|뷵������{�`�k��!��E�?(�k���i��.�u�Z�9z�S��3՞Ұ3��75��yshq�Nŧ�J�#z6*��R&ɑ��.b|K�%�"�{Au�i���ꔉ�YaIn˝J���42gi�T+�w��/"ѷ�����Y2��}���C&�����Y�Cq�>3.�9����]�~���,��������g���S�GS�@�fyT!�W�p?Ott��*X�T�mC���v�T{�3��zc���0�*����X��O�Y�F�?�xW�y�6�1gĥ�M���*js�e���fQ�<���}4w� },�;�E���Z�I��w�k���cgs���;[F��R�y7����gv�k�0�:�x��7K� ��v�B\M��z_R��]Yz2��ds��p�r(�_*�9{ZCE�w���*<57�3~���2p��5p����u2_N
�&Ŋ-Յc�6��y�15~L�"�����3l⩹�6�on.o��؁Y�.��j!���;�c�5�Ò�jK �N�ʬc��ճL���Uz�CzgYnx��E�j�n�k+�s ��W��no��b�&X�oq�"�X����Z��b�v�W��9n�~f��BmW�v6�r�^����8�ŴϚ"���bYq*�r�����G.S�2���zj9O!����b�q|�/��m*�2T��x쮘�k�y��YF��c|FL�Гsfe��d�t�(Gyb�G��55�nMZ)X�N3��cVv��:��ݽ�4�aǅ���V�}o5t}+�Ӳ��O���N�r��(��9�cɗ��jkoo��\��v��t-��f�
yz�t7��x�~ꉙg���|�&����G�8��	U��K��c������&XS�e��{������˻�q��?k�(�<"�fX޵T6����mR!���8��2�����0&o�l��`��:t1�7����l��~}�B)��H+��:y˰�ǁ�^�� �3ߖ���0��E*�5I�bZ����]ƅ�Phl�Dq�����D��s4�d󏙂��6~��/F�}�S�z9�2hI���hr����uជ���[��P��w�F^�{�U0�e���;^�C�������z�'�Ƈ���b(40��9�ޑ3��+~�f9ƻ������!	Z���r������&;�����09��"�7.5��t]�ʖ����u�<^�'�}��R�C4+���'����3&a�w�;AP�`�Wc����ӎ���>�`G�f����S⣊'[����Nч�����g������=V�l��鮭^�S�:���e�i��G{)�z��������DߎI�5�Qo;���z�t�g�0wW�-�/�1.b��4b�*�&�{ {	M�y�u�˓���]�c�kwp��4l���fQ�v��4�4B���u�#%�{1��YUi2�s��6�Wp�|���sL�V�s�Ę钝
�S���5�vuo1;%��l����a�������vŇ���P�CN��t�t�(��^7� ��kBQ��L�� �C�Q�����K�
cvO����w�@ף�V=����6�`��(����9ђj�J.����'�����s3�o#��΍wօ��ېC@�S�)�H�c
N?$g)B]z�*��+i�K��e��N���b{Gl�i�3�+��+ꈟHgU�1y�d�χ|}0��ǊgwAeF�q��7�,Hѧ���t}2�PdO�T^�����h���z�X�'�6�֧/�^N�#OɌy�@v��09��kj�A�/�	��j��W�s'b��1���u7�KI�7Z�o�c7���O��J'4�$n��	.xAg�r��+#�)w�Bk�gUԗ��νOI�q�\T�r6<�],��]y�5�k
�?pGW@�Wx��s{�%o��i�R����.�>
�<r�
f���xz���-?��-��:Dd�|��b�x��|<7oq�s��9����w�5[%���Ü�w?ܡ��S�d����<}�>�O����z�~C���y��>���w���X4�֚�	a��.�~s���el�����Ӕ��ǘ6wJ���Q�դ�qć6�3x���c�GX6M���(m�F���UeH2l�3\�1Y{��8���*�7�[/�8F��n���n�ɴJ���{�Z�Pv���􆞍0I�b�qGeBVc�1K�*f��Ő���$��؍�|���@p[�h��� ɫ�/i��KE�����#��mi�cm�����?=W1�C����קzAL]*��9��j��VZj5һ�r`�q�5�u8�.z��%wk���Yb�}��r�e�J8(i�9��[��-ډb���	p���j~��z ,�w�/·xCg�&�֭��(���=Lø�;sV|���m�ǭ�X�V�Gr�%m�Y}���3�)
�8槗f���[;���M]�9���lT�Bж�[8�g1���v��|j�QT�f��yɟ7�V�=�T�����Y�k-V_}�#,�V#���kN�����X�]!ih��Ȟ�WQ�A*]J�&�Qov��⇙��xoV�.I#� ƍ�}R��O�m�*�����52�,#g2t[���-���/�Oole��7EG$g+a��R9�;��C�4E�[�7;=ށT
����Jl�W��<��k&��H�b���T����zAѥ�����/��H���7-=6�&v�槽�m���ݬw"ܓdcn�1�j��?���ޅF�>�0�W��.�NB~���O	�u��*�FJ��ω��{������'�3O:Q�\��\0��G7��C� ��S�|�(�b�õ-%w��q��@cv�vO���(g)���"\˗�����fG0��rNsx/���@��Տ�
˷�]��jeiņк+ZvI޺��e)q�թ�*ۑ<�&#���j��4�eh�X���i:���21:Ӧ��:�)��l��#�_8^�ގw�Q�r�c�EnQk�Ƹ��X�@� �ʰKVUV�j�۔i%xD�r�1*qq�}r�����0��7B#��A��z[PЭ�įRk~�к�˜����"Ր-�Mӱ��57�|�@��A��A�{�N
;��So6���`��AWr�=gy��u�
�ʔ,�/�-�k�}�%dv:��Q"�,�z�֝�f������6�6��A��bE
79�U��L�(uY�f�銳a�lV� �|�rÁ����5d�u"B�҂�r�ús��c���2��&���f�9R
4��5�z��*��5+z ��7
C�J�������'s]1|+c��L[����-j���1��#ʵ�9m�9��{�.���a3����q"�"�4&p�kk��ݜ�Fڍcj��ƶe*ݮ���6 qu�sۄ�dNM��t�`��a��&��[p��sz���w7���:�Cۘs�U����!�+�__�����ĝ�U�բ�;��I(��f�CZ�"�m�^ݺ�:�6q�"�b�"KF��U55E%h������:�5mETSbCA[j�v�MMPSSAUu�ј�*c�1QѭF�k�E�QT�D�11TLUIULN1�ݸ�"
H����T�j���QF�H��AT[��֓MPDDE1Gc�M�0EEn�:�:4EU14LRWA��k�UV�Z��u����Z�]ET���R�05D�5MU���5Dlh�����D�T��WC��UAF�"����Fں5h�b��6�LDA�MSE5;`��T�T�5D�ILSI%5UUQTu�(&��MDQUE٢�*������֨h)��&`�()�٭SkK�()��TSm��0q��b���%�
^ÊH��
�&*""�)��X���h6t�M4퀫cTĔT��7ITQV�i)")��"��������_uy�����f�����ޒ�:�`ۖ���\�8r�M�����R�%f�<��[r���#'V~�+�wV��[02�J������]�˶wy��un��s��R��v�u�(�m6,%ig!�;��%�PLL/��Y�]��U{6�����wi�w콽���R��#�&�`��w[��CH�rZ�E4'�x���bj9��֐��x{�dh_��:��kD��	��s�[��{��^s�4��q8y� �s����5�Ě�F�Qj�������fR��<�:uf,>����۹7��=%��=�QB���&��W&GQ8|Oʟhu^^��
_�A��֭�'-L[�OY�R�\k����OE��{<�D�r�1�z���]L�SK����@��g�d?x�R�,p'G��z����R|��U��$�wK�f�ވǊ/B�Z���U���u���癧ٿg![�^C��h���hƆ)�p�+m^�l�h��),f�F�,���'���۫ќ�����]�����wm��-��C.�1�C1����l�,!6�vl�8�<F�I�Yc��ة��$�d�7Dc'�����&�lb#�bKb{5�Ӭ�[��<�gYa`�&)�EI�XOM���� d^��00p���˚�6�5絗��vD�DCF�F:l�p!�l�˾ �{o��ϙ�c�vB��:�}��d������:�b_��}u�LP�5���<Jm�J�d|M��Ve�e���Uͼ�(c�!n��g7*����n�[� Z�Q�cZXf��XY�G)Y&t�Y�N!:�����UC�ٗ��Ι�[��1Ƕ�z%�O��4e�x���x7G��9���\p�z���W��p��A��C�n���9l1�͊�tvq�w�R�~[�	�֣��%�l�\%u6i���F�n��&Q~"3���C������C�9��e=;E�D�V7�NM��,��5q1GWe>����zd���V_��@��.�j��ai�_E�yW5�ok�a+�O�W��R�w�u>���5�p����EH��� �����dD����)�M�%�Y�OݛmCr�I���p�21~�00��♰%t���C��}r����(�ұ&rRD9�M��qq���mq3%�}����P)�u�ܯ6�QL�M42����. ��WNt��s��u_g�k��.�|F��?�3��o�n�b�M>��� A����p��X����X�2Y�y�VO�dh�Rp�+�Vh<~����շRS-�W�Jh��l�cX��t��E�E�vkv������_Y��m��u3�} ����*���b�y��ZY��ht�i�K�,�n��ދ���UحCR	$˾�=��i���׼��ѵ,���ea����zZYω{�n����w0�H�Y�]��1���<Wg=���m
܎�����b�e�l�X�;�����8v�;���y��fn��Vp���@B��x�� ��iD���!��~
'8�@���}3���H6}���+x�B��s*a^4���K�\G:��x>�z�Q�j�X:ED:�n��h����/�s����-ݞ�߳���Aq:��4z�ħz���̚:[{^b��\����?7!�����/A��eR�O�ҙ�p�xw��<)�����>�	��jB�q�E[� ��� �ξ��1#���r%��og�	�^%W'N価W��T����Zy�EW=�\��%ŨyDj(�j�� ����U��B���<��K��|���ӗg9��f�G2;!AiZ�.�C�3oHx��
��W�k�$h��:y:��7;ו�YiS�� ]~��j��S�MV�'">��d>�����
~:��߲z�5B�Moz랓ϰ�P�숴�\g�
���(OJ�z�kƀ�y}M��Μ/�ѣ�ݤMS���ȇ'w�C�/@eC��)%̌mk���w�zE�eyW7@� �<khͿ��%?�
L�j�9������h�{y���ݛQg�R�j<����˝�����1̂�Ad
�+9��Z,�	�X1תX^���sth�>�CA^�s�I��w�*�mP|kSyz����?�}��۞y�i�b���0�2f�2<,ǔ�ɧ�_o�˷�o%�?�-B\aPK�a�����m��g�x��E���n�������6-�r�iv�Q-1&p�́<��O�$���+�;����&�F�{7�}�l���Nu����"�����±��/��|��ac`2?*����{r�}<TX����:�{�8��&�Ҽ��׬]/�`%}��~X��(�Ї�*�+c�bH1��S�C�C-��7�l�u@��K�r4�RsA����!��`X겍��iO�6�+TUK��ו8�2�ݺ���,�B:$��tTyB���)>�sQc�唼�Q8��@�����g�,�h�jv�@4y�QN���&]��84|g�7(E�9�G_<�Zrpj�|&�sJ8�3��׼z0,�vNKנ��)�D�6�>!��<��"㹵�g��I�z�Z�4�sn��<���F�����A��Gp��!�Ǡv3�80ι�K���-�H��h~��AF�,:�o��۹'vyK+7:]bx�#�Q��c�@�k�vQ�O���y���9�F�����-E��#uPɢ�z��5��A�.ձ�dS���wmv�9[���M�[�N^��U��D�4T���ewj�=���FaV���!`W)�ȷe*'2���܅���$���Ղ;p>���{a]�����Ɂ;����f�5b�V����p�_��"���&^�\��������zƊwŲ0�������T��P[۩�r�k�/0Ȝ>��Eq���(��5�m��ʷ>��m��p����~��4��{��u�t��OK�#N��g�����c����-8�b�k]�D��x��eՓ˒�1=�z�	��@��$9�vl0[$:�43g�hj��&m��� ���,��<�Q��_<�/���A~_Q-����/���]�`�}�����OW�o�"%�u��P��E�t�Q��M�1�hK9Ɖ�/��i�=��@��)]��Xv���S�n����^��W�Pq�	�={��f�Uӳ�)�u���!�^Cّs�f9셔�e��fm?q�Xa�?]�<�5#/g��ˁ�9�P���I��W&E}�������x�GU!K�Y^���p��W��B�KҮz�&�ƙ��(^��V�D��֋Xo_��M��͉�O6}�H~BpeD�~�.h��>d�� vD��;�O��g�}ڸ��U�@����a�_�U�2�4�VdU�F�9y�}�h�Wj�p�b�s^�S#*�Ė���2<�p]��C�:��gR���}2�N-w+)�3�8w]&���*wA�2V��^��t���`�U�/Z'Z%���#�U��X&Toՙ��=�S݈]l�/���/㾳0�{ℼ~&~����=L�0[ӛM��*�=����$�zY�������b�Q��V�_F&�s�tp�*>�yd"\J���܃8˭�N����j�纃T��	⛹�(�p�r�������oU&q��.y�탅[���E��T��t9�=���}�L$R���1R����s�0|tI,��׾��>c�[�4���'B��gI��߰���*�F\Q�U�-#%���y��[/l��i���,����=����ݞ��,��'�l�b9�DLv���l]��j\v�br��|i�б7fdؘ�3kn�v�V�z4\_*� �D�㡕�מ��=�z��]�[�N�Do�zI���[0u}�fV�11���H�mj��\�g;4�މ�46X�E�E��q됯��\�oc#p�f[x՘�6�����p��Ot#>�`��@����8&���75	'��i��͖=B�:Ks���#g`��ⵟ��,�Lf����hu��N�����
�矮:8iU�GL�.> mdhh�%M�[_����IՇ�|v/OM�K̹W�/�zNw�7d��5i{h�i�W��w^~.��ӈ�~�7ɥՄ��Xh�"�6o�v+l��������h��g!��$��}iqy��5u%��	i�|�Z���yBzI}�]^ʷ����3!�u���b}{�1q��X�_s�%��Ý�L�%���	����29���E}'�R�91�wf{�-��Z��%6�"�ӡ�o�w�,�{5���Z���Q�d���?��/Zdq���R��8{;�LI{e����$"�9����#_ٶ��J�m�y�\wr�χ~R��R�
S�>-��&����M2�XY.jq� r�@i�d}TSV��V7��̱x�6��%�+K�ԉ�;�x�߫���r7(�j3Ԇ�tL�1<¼;�S-��������-��f��2�KR�3��||�}��2�!�a�Ũψ�1c����_l�����o�%���}��������Ł.�N������9S��4;� :S˷7-�.h�-!�I�\XsJ�|u_��G7!�٩#��-�Q��ݜ󏃊ه$�ۀg�S2΅]#_�ٳLkئ���e��J���V�A���.�?g-2&���C+���v�< �=�ز�xB��cz�Pڽk���d�������;���5x�b�0B���n��b>���[�gZ�^7�M�e��J�a���6������Sʹ�b9��%��`P�I:��2����ʙ���,:��j��Or%V����ǲ��okl����1nV�̊wN&�ԙ}�vP��N������9T��W^��Y�:W�2X���-���;e���I�����y�#��.�+nZ|r����k���/m��M��?>�5�k�<�ũ��������,g�-OV�2�4f��u9|1��f�&�/cSߠ�˧�((�j{hxϟ���_~1p��v�W5x@���9'�/��͈�Zx6����u\̴c�Й�c5�0���C�:�C�vI�ٸ8Ub�;N6�q:�P~jªل��82��P�e�O����Tf��A)��_��6���o{�k�1w�.r�cծVz܇���t]�tg$_�}7�M_[�aHLǳ����'�Q!+���O��<��/wU	R���7|�Ef�d���Ŵ�ڊɣ̯)����%u�瘱�9�q[=�8��_�q��L.���5�30�5��
�pZ[����[~d�*�+��{����k�Sc��w��[�w+7y(�����ڵ�MD3�u���\=�!��c��+6ܧ��ذ��ѵ5Oo۴q�k������<uR��V���!q<�nc��P���(B�s7���;�k��������n������G[�Nc�,��jN=��ٚ�w�]��Ģ���_���oS[��\�2��E������1$m���L�k��۽dx����>H;�A�ܦ�����%���k���׹/��i�i��v��@14��oJ7�qҞ��>R^TO�z����>�T�#�'o���e���2�ߥ�z�����s�A�hm��ZdC�]E�m%EL�V��Ep ��f��6e�?��w�tb|e9�wVX~PƦ�p3l�ukd�����fT�g#Y(��B2Ԉ��S=��O��U�.e��Gh:��N�8Grq��B���T5������k%C���}�c���8�VfB�ڙ_eti;�ps(>χkX��x��"���\�k��������=�o���(�:Ű
�m���^�jK�s=���#o�"�T�q<\8�|���ð����n^cz��"�j7ʝOCi��-`�,>���t��*z`9_%>����|�^^�eXAn�<q4��F�4.AH2j\�IX4���L��F��#��n?��k,/���ۿb}�2���=�}�lnW�q��%e�i�eX��U*�ڹ���c4�%ܥ�C��Y�j�t�}��
V�m�NE�X�����[��6yU3F�u:�T��v9���J0M]���n�_kC��T��3��p.��T����V�Ze�6b�,��1ٷ��v���: ����z��wJY��A<�[�:d����k����3T���=�W���I����U���^E@�Η�WB7J]B�J���-��+��8g�iF�$�R�E_�S�Zv<�d�C&�qZ�Ȩ�fj�&A��5��1�{Q%{gbUnW,ț�5!���"[J��=�|�i��K�
j'���.V9�n�%m#z枷*{�n䬆v*�E�Ux�f�-^�u|�a����rf��H��y+���� +���QN�rv�.�Bä{jە��"�y�݊�l��U��IG��c�ա�^x1P���:w�^�"�ޯ��T�Fu��'Ś�������~�O�����������������59��5����>���K�C���Ŭ��T���2)(U8vr�B�R�F崵��ӗ�)V��z�or%���u�M�t�[��f�[��Y�Ǵ+ܶ)�ysyv;f�8_V�FSuWPP���U�Z�����[�x;hv4^.f�V�aB���n��L�%�A0\9�F+gn֭�d�æ��Y%:&d��>�N.���v�\����U��u�jծj������je+��k�5���;�y�䳶�ˎf�Mr�y0��q�yby{H����AA�͢�.D�j[�rm$]���;l��R&y�隈&9�!�¨��hX[�����{��|��͔�>��fg��\,�c�"�
�x�B������-���2� ���^�Y�wW٭����q�@C��mD%Z�]
�1�޵���@�WG��kIv��wݐ_��I;���q.]�)��M�ð�W���h�⽩���o�wM	�Kr(:�޶�ܘ^�~S	�5yF�v�JS�n�E��p�M��́AS������Â��i{�m��CΆN�(-ʽF��NKt�$�u��s.ҙ�Ph;�/H�WO�e���M�\D'�
󰉤g��J��4@���v�SV�j��[ޛ��7�GƮ�5�iY㙐*`uu7�M�xapj�}ϞU��,�ߍd.+!@�A��ɦW2n��6G����Ɨ�*P;��	�u��Yh&8�}+�����8�2��lj�׼'��c��G�ʾ��4Z/�E�/P<���_W��Q�?��M���ALn��'�Wbf�7M�v3M��0��*�`G{�ժ��3p��1m��Ep8���ԬͶ�`���h���ʥ2�6�@��!tw�Ċ�q6��F�ȯY;�5~J��t�&Q�랿&���V�c���:+��N�mGW�R��v]��{w����|�	w�9������aF�
5��1���]+sZ����m��U�(��Z0���6R�-���Z�m_+�]u�wm�}wb��"�o;��X���m6o�33l�r.�9��l�׬o
�o��I�rĪCN���gil�6u���e�e��DX4�e>�ʻ��t~/Ns�6�-�z]7Ե`��)�KOu�T�6��@z�=�du�uSI�ff�s�P�佧�r�m/�Ֆ�أX::��ЋiV8{;'%>�.�.��[ň�;�a�!�U5Jg�I�sk��Z�`Uڢ����g��b�).�dhe>ʺ�{�~\!1�X��ס
���u:Kf��s�ݮA�n��U�X�ۚH����U��+=�oWr��Ұ΋���2&����3Ԅ����|�Á��z^%B0�=�g�}o�5ԾE���\���1���F���D��t�+�_5Nͷ�K�
]}9�m�w}J	k�O0-q�ۗ��X�w��0 G-]٧��ʼ�q�Oq���p��q*i�����o#�q5U]Y�Ē�I�TA�����h�H&J�cZ(��d�5��)����ih���tP����d�)&b
"��5���(�6�U0I�(*����}]TE�k�SM-�CN��Z�*�� ����&��)�*��44RD��T�45Zj�E�1�:�����I*���kFآ��h`�SSDHRQ�����DRSJUUPQEh�q��h*��(�i-�D�h��Z�NŤ�i)���Z*�֐�1��(��(��IMMSLE3R�QSQ�4�C �S�[��I�������&�BDZĕE5@SLAT%S@�ZKE4Ѡ�Dl:(J���mZ��M%��I?�'� ~J՝�^���%�B�tm�N��6.i����Y+wo��JMǺ�KZ��Y�X'���7f^�/ps�)ӡX������������ �6<���[���B���X�[���}��oV����
?U)��i�J.,�@��8�ţ͉8��!�����S��v�nI���Q���c��I=q"���������)9��}��q2D*o6p�|���h'xHJ�x�Q�3��U�R:1_G]��F�t�����4Ӿ�q7Ɔ����Ż}>�,r��<��e�V�(B�z�Dt�][�;n0YWT�ٺ����3I�	 �����y_1�:&�r�|>ݷhާR:[���*����R)Mz��\�;��dM1O0oܪ˯t��Q�g7�FO�[M�q"l����nU!﩮�(k�Z�ڋ/v5�xs壍v��BU�RuE�ޯ<ŎɈ�PE��i�I�"b�S,����9sS�'ÈUfu=�UБJ.�ղ=F�W�S�)�mDh�m���8���p/s�8�[���EY�lx�t6(0����Z�-bGy��[����~:�X�3g���eJ����»�m�3��Մc���C��2���j��bppD���i���G�l������ɖ�k�<�Q�г.mV�����Yb�%�k=w�E���*Q�a*ɥxۡ�u&�i�6/��N��VO�ڠn~<���<��ox�H��q��v�(������
�e�#ѽ�gE0�#��j;�<��vk̶=6)��>��~�T�K�͠�֫"t"���c����⵼W3[a��3�1z�ƲL{׷DZaNV���W���۟&��[�[K\�M�#a��������]�j�{���x��T{cu�]�_��i_{Ś���ʟ'��_Z�K�Zv��f��7�5�L��cV���Y|z��s�$3�8�r�=f�N�E����9��|��c�)��l�فح��n�O�p��X�ڡ��7-߭v�� q�:��C�6{�]Lr*�0� �;N6�=rʫ2Z�\eƜڗ�S�T&��x��`�.;������*�;T��=�3^͕�U�wz�\��	����%+�vl�۔{%�*�j��O4�MLxb�S�tMKx�fm�fi�¯5K:�S�a�kLvOʼ<)�z�߽a���;�R���6sI��-��Y��c`Ы�[���w��p����� }ux���ɌPj5w#ɇ6��:ǳ��׌�}1]Ѱ!��Z������L($8�m�L������}�#�]wP0Q��N�u�\��)�ޖ4�f�YF�d��\�y	!��T�R��~�sʃ�ق@b5x?;/����Gp�� =����Q01%��E�[A+�)d�ڞ���ߍ�|Hݬ�5�ؚu�T���\�ַ�ϝ+/ږHd����p����H�f���Ve�k�0�n��-NSN��:��Q4G
���љ���!�s�]����j���U�֫��h{�?�|*�����X�~?�.��D��^42/�1��il����Q>|�K\�0L�t���t����ȼ�c���<x�\�7nO�8ŷ���w`U���A	��ۋC���ֱ�^g�E��פ����$�(X��#q�	yk��y��P��-�`��R �1�	���U���[Φ��ב����RK2ޟ.0[����Q^r1+��nW!�GQL��9aIk�%��㗻��mɪ��vp�5�5UE���_IH,E���b�����`��ɗ���ժ�r�p�Y\��]�;�ڙ��e�)���t�'5�VE��������=s	����v�[�(>|�P��r��{�;]�ySn�Հ��{0�܌uhoY�_�U��u}s�w��Ƒ�&1u��g9r~�lR�t�/itnV�N�P�V�M���~!�}��2�D�#���5��}�Ó�-xt�;�w�h �ɾuP����,����Ly�vb h��!q8�v]�Y�e�n��o��d�H��:�EjgY/"Ku#:�c:�q6K}��������M`G�N�6�ѿ~Z�\��&�{?d6Q/g�~K 7*��R#���;V��B��^;����S��B��!���vEfZ�0��N�3G�f;�'�'�oѻ.�f��iF�Rӣ��{���3KL��K6��ѧX�.���m,�6H����^�]>4��Уr��F/Vq�Z�H�u��J�@�w�V|�/��?X46Bx��
�̷���X�}�0�|0��F��$#�Rp��`�6���X\��r���[+M܌�[IQ1j���d���1����em�GbnI�mU�%���E���p��fڬ��&'m��u�u%|���q��Z%nN%��k3�t��y�/I�n|����F�On�%l�H���
���k��1���O�������6k�5f�TM"��un������o�+�^���ؽ�禗���>=8��#� GzE��W&�g�}�KU��(�̳�l�ƷsG6�_��Ʉ�u��F�0Hc�"c��u	��Fp�pC*�d�j�l��܃&r����`�4w8��$q	m�Fly�?�y�'m�}Q�Nif�ٵͲ�*���z�!�oh(�r�@g,���0]��1����c�I⡱�k����.��r���N����I{�3d?N��.4����,��j�묎�VF�8�e����=lp�=A*D�������}֍p2��C
~�w���Br����i�GI~��C^�&�i�c�%�#jm��LF�|���{���Sŗ+�¤�*��x��{z�T��	�;���O*į���
���� 󗱌�{nߚ�y=���u��|G�Q�ǈ�.��)��!���]�������n��;Vq#������r�JG�b��n���Z���� �3��9X���z�Iۮ��m(�p�I�,�5�9G�6��z�N�a�<`Q!���W6J��q��iü��}�[��s{^w^�c-��햣/v9My�M�vN�_a�D�^s�m�A����@�8���.��}o|���1�3�$,U�E�)�}q��q�$��)�8Ԇ�G�=��ЖPK=Ib�ц�P+2z�n/��M��;��;�Z��j�\v��q��u7A�e'�q����-f�u�	��mo/�.��u>g������@��v�H�Zo3o�����s��%��m�ړ�1���+�E�nS5q�:��b�k3i4/S�מ����V��t�vz��%���⳨�3��2�>�ޟD-�R��4���t�sv�dj���6�zm+<�a���k�c6���>�|C��Zҕ,��S�vM)����|�q�s>���#;>���][����- �m��n�� �p]t;W�gƲj��1���G����^?���sͱ�����Wa�ኄ�fº"όP�}�)%:<�<�w�(��2�6�W@+�&<���6S�R�p��2���Z�rg]��B�r��W�jl�3��L�SYoPtx�w"�g��bGsV� >x��G==~�r�|6p��Z�=Y�9�`��"�壷/��OU����C��e��zkф��}o�3�O#��Qv���3�g�[l���^��]#^C����2�U���e/gE��6�v�~m�ܕ���c�k�i�Ts�#�:�E���Q�|Kh���,��ˬ�)����E���K.�Ѭ�! FN��*v�ʝH��%����˂�/��^�T+��Wi�r��Yڧ����
#$%+m��x�KYj=��dî�޺���������_�8��|�5jV�J�(���yɈ�09�K�m{��lޘ5��E�FE=�O4�<��%#;�J;[�~�oq�Gte�W���l�s)+|V�h1q���
h��u>�z��2�f�75�v�h���Vk �Ky]�v�� 	��[��/{<mS���f�.�l��^f�g�AyD�妯was�Dd٭�v�;�J�mT�P���tȝ��V޳W�5��y�G�!�)��II��T{)��8���S��H��2��wr��햑�Y.���9\�-��su����k��͂oz���vc'y�lf��nH��e+v�؝��F%m�|��kl*�y[��N�m=�_z�W�U��6��ǼSo�w'��G�D�ʵ��h��`*�^gm�Mp��B�Dv���iUC���t�������Z�������q��3���=�j��(О��5ȫ@,�SGv�g��Y��x�B�n�r����O��|�>��;Q�����=ֳ��6�E��3w]�y�E-{Fgdq���i���h�b�
�E_$��mg�~;)�k9��g�m��k8j�nk(u�@��h6d��28aa��;����̵6�7Z5,�7�r+hW`��W�Ӎ��}���V��=��m���[/�4Ο�$��$������l^z�3�������r �:��qڢ_m���^�o^bm+����~������{�a.��J�^�%O�Ċz�zL��%W�iU=��2f;�{(�bij��X�Q� ̸�-�y$#-�x;g�,����k{O�Y�)�#)���כ�����݊%����ծ��HU܈=5�ml�e��Mu2�\"����Er�G�.�b�r;�������~գ_2^HmT򨞩�K[x�z���"0��Xs�ߺT��kܴ�;�k�����2�q���W^x�rP.:ڦ��{b[��k��K��e�����u�R���y v�U��K_f���S��.�l�R;)��4�r�v�$>��s�C�H߱7�@�R��OV[����/�3	O-�7�xm��}F�U4�0�^���MC�2]�g�R�(�?�jz	��J��j�����֭���f'�6���T����{^��oZ�$��:H^�I��Kх�g%��w91�z�WJy������/]����y"��ݜճ۳4�*|t�#�l���e�.ۃql�R��S��ج�w�s�@�c'1b'�֦�����u�[�"5\J��\ĳ�ͽO�<�F��\J�����W/�2F��4y������4\e(�d��b���kYy�{F�DM���Qw\�#@U��!�4B���c����#�I���WJ�VC�Ɓ���che�Rʙp0ç�';;��x�3�p}ՙ�4���,��Pʽ��x���/�/���Lt�ΤVv���(v^E��0V�t�ǌ�|�����~�4�~��l��ǄG���P�[��0��dc���3�v
1�Z`Im�|&D�.,Y4;r?Y���q��dK�����vU�v��R�m��� ��f�e��Z�f�񮮙Q+�nz���[�f���x#'#�����M#������+��]f���뻗��9��Gg���k&8�j7v��Qඝ�M:���!�!��˽�l<rxǥb�#��l[m�q]��]���Gk�-��˵.���e��)M��{f0O�U����.�$��竺^(�p�-�������C~�w`w�Vsva�ɒ*��[��Z.IqK7ƄtI�*G�\���1T!�2�v���t��5�Kf�S�V_}zZ5.��:�*]�8���R����'�e�����E�{�)��,�V��f����^�_�����}^�`�yy�ޟ��i����.�_3�q�ݠ��o��t-s_i�ޑ�i�/#�N�Y9�-�P�x�	W:n�D.} ��S�(��X�xX��-�^@�)�K�x�^�ųxX�ᜑ6;�GS��=�
�fw_7�H��:Y[�p��92+{9b�2oY�L��*�1]*��$�f�mJO6"S83�U�K7#�ӈ�GUDm���yI	�����_��su� �\p�#��t��܊U�K�!�y��q�+�Su��;�הO@�2M�6^'tr��P�al�Wcz8�/v«�nI��^�-,S;7&e>\��;��y^vNV­��c���`��U;��w7Yk �z9���yp��ڜ$=M���y�31ev,�A�A����
	���n�P*j�-�ʱ�s@��ӧi�s"9Y�mK����Wd&�6H����v����ǰV�K��gFT��
'INfQ[W�Z��]x�����V����P^÷$/7e��۶)�gAw2�S�z�r��$�3n���+&���E�-*�7+b�N�^-V��"��]d�@}�t�,�>6;�z��A3�OR&e�p\|��]Ï�x��44�ωחrWe�0�S���z�N]�1=����H�x�P���C��y��fnzF�*B5d��Jd�����7nl��O���k����+@���|���#��V��Q}�5+�]q�-���#� ��&oa{@�NU&������;[�+�7k;2�"�Amh[]	�vm��r��e��ذM�bVJ	����[v�������h��0(�Jd�N;1Q<F��r�ir�vn+rQSQ=�>W�I{��5tp<xB'lP�c�����=O�Jk��
�5���%@�Eo�7_zvl��Z�{z4��ƹ�+-`}f�����b���Hƅ^m�f�!��_�-��s���لe_�0�u�/&�˗LP��HYg��b:���e����
��2�E�s��R��&bLO��9%�C.�d
�Is��U�q���e�ɧ�X$pv����a� ���6f�Dݱ�K�Y�PX,藸2��a�2�7?&u�Z�]�=m|ҹA�42t���R��[{5}�gK�fư�(gC��#RGh�?^m�R;!���z�d��wKI#b�}v��eK�7��Tr��a���Y$��Ѫ�23tk&�ǣ6�"�I�v���A�766e�����������Bb��a(������jS���>:�G��蛛.�Ei/,EU�ޜ��U���_V�}O���d_e㺘��*�,����ޅ-�f[�5a|��O��7�r��Ys�U$V���R;����G{�5��oF�[N�s�;�ੋs.jf��.�ܲp�{��9�H��4r�W��6�/�j]%1�j`5v�:�Y��s���ީN�98�ua󙃻y:zQ�*���8�M�������DTZ]4RU:�I��ccC��kKBQQR�,TD�6��i��J#m�m�M-T�U��T���K�EX�F�Ѣ��ZR���f�����6Ml�F�ӠkL�!Қ�
)mh����#f��ڣK�m34RĔ���4F�E�AAET�U44�ĔQV�:uI��������
�"bh4Z�k[V!�AkU5CT���HET��Fض�l�Z���N��FقGN ����QHD�UE8�,HTMSkChtD�ECT�5%1%U4���N�1DPU"�S��hAF6h)j�F�b��$"	�
������A��U�	j���c�U8�!�Ö��,'u9L�A�&E��eM�B�B��軋��{u4�A�K��ݾ�*�j�j𣏕EGt����[c)U0Y%D	_�D"�i�0�_�	91���tk���$3z��u~1��c�t��uxB.g�ղ���ᮭ���~#��#�]r��~��U�{o�K�r��Ż+�O����p�O���|)߲�����VMU���H�1GfEi��Jy.匰!m-s��d>�0��"/���}�ªK�t��:�L��޾*�[�ɨ��-M{7���sīy��v��s��.�<�Z<ȩ��#��ߞ�?%��f�yE�O�8��z�E��6;�3����[�wLb2 ,7�wض>�޲�W7\�M���l�/u��h�����9@��o�Y�m�~(/�������D�d���8"d�+;O^Z��ѧ1"��H���a�K�C_;��M���DOM�s����p�ugQ��v����QF��BV��:��x<gP�F, Rƶ�ѵ;��t������R~��Q3\By�Dm� -�\���5�߈^�����\�u��;Rqp!%潴�R� i�!�w\�:�A �u���μ;���ʬ6��7�k��7:}3���3��y[���{����?��'h�/�n���eh�)׮�������|�f˽(�k�َH/\|�"�1����47������QR���V`��+���_>3ꬽzh����::.O�-߻�߰5�T9�$�=v��@r��$�3l�`��|ܧ���_*��9�^*r3%�e�D$ T{�ŝ#�b��{b�#Y�X��{Q��׸�4,�M[\�"N�KfG���BؙI���Y�87d�a��qu⧩Uv�w[$Uy����H�ՙ�
��<���E�f���Y#/U5zr9��q�{|�wJ�Y%̻qr<��͠�(u�6H#s&c��>3�ˁ��N��w���@Oxvn���q6���Q�����8ճ��������`�1A̑�+� �U�J^��u�x���X"^y�"�!��>����km���>mO��?=����$���(s[�O��Ŝ^��������F��o����q�����	�w�{�37����{�r��!�9���{��Dt^#f�fc�e�� J��m�P�ۍ��G[�����5oAG� \��%h��j�>�R��s|�廝���m�x.$�ju�cn�����ͼ�܌N��^֊�9Q���T�^ER+x�a�c��J����{����P.r��rZGv��A� ��3�y�?�'̝�xge-Q��m�����\gB�+9Oq���9�^2z�ZZ���u���.�����Uj����x�LM�{�`��-~���E$8���^z�e�fDs5~а�j�N�qX_��G��x������%�"F��.x�]m~1zn�"I�Q��U���O �Z�8
��/ѢbvG�%�CL<+MV��c��9=g��7��ڷ~�m��C�[��H�+γb�+a�I+��Ne�+k�j��W�UM��Sxˤ5�m,��㬎��-�]�oLdw���7�
��V{�e����J�.��ʶ$U��]8���Bp�wtz�Q�"�ۧ�wdYW���$g�av�Y�	�.�U��g2%ي&�vS�Y���6���v=^�H�*�~w��R���~O'xyOs�b�<i�b!��nipR���"гzFԘ�4F��u��!��-)-Y(퓭�m.F�cff^\S���@m<얳5U�]�E���J��G��ts�����V�ws��n`�T�G�N�B��*�arܑr薸wu��q�뇚���+�[�6�KG���c��ћ&@�Q|�0]�_�&f+Ζ��g�(?>q���[o���a�$[����u�oL��2�3�����\�n��˼x�z�D�x�x�����Ny�[��he���<�[��K��Z�z��mf�q�׉�7 +i�wNO���4}�[�ޭT[��[}����c{	�bf�]z`��ӫ��v�����d�o�����=���p���j����Ya� +Sr�g{c������'�>؎��O6-�A>�Jgr���z���c�x�;Ye��v$J���.Z�v���<nњ6ϱKe��O���+������=H]�-����+<ezl͊�Ѓ*}���]=�fqǾ��6���'��/dg���K�+�x��9�:m�c|�e���F��6z��W�5��ůŽ���T��X��v9o&���5���
��$k�h�5tqhG�V�/T��jW,:�X^F�Z�a�ihfQ�	_5���U��߸�;���{�
�f�� ���� �� �܂*#�Z�2�èS��ݤ��|{Qtn�ðq�쁉>�!�%Eoy������3X�������h)��"ڝ�E�W�HD�G�|��}�g�w ���x��.fջ���!���_�b�P`؜�M/>�\��԰���p��ҖZR��]��I;b�E�D0�8�<}��a�C�U�z�r~��_
�m�.^�2��L��M��U� �fH�r�f��x����t�Uw�.��f�Ců>��-�)�������U|�z��w�e�{�>�Iw��s-ղ�ȯ2�
y���]����{�x��l��n;8��+�m��n˞+:�����ڦ�9A�+�{�cD�=U;1z��4:ʂ�r��¶��f��z�%���Vp=�:3���nW�̩��~~$�x��e9�Jh�	�
��G07N/"^�NeI���v�y�[�":̋�R�vy�V_���Up�j�]� X3�[�5i��Rz���k��c���z�"���ZG�����W�5/(-.��2L+]gO.��X�}�v�F0�^��ɧ:���)8��(Zî�Tv���ǳ���k��ބ�hx��'^��JԞ�it���m��ǕrMF����{6)�z���ؽ�2%�YV�NVV�q��뎆�0���eǲ\ѐ^C�v��2���U�T�U+/&��h�}s�/^�dl��D��)���6)x�|ip�"|���m���[�����fd���x4��S��S�Ӿ���#"L��A/��#ټ���O��D��J�l'���Q@��
��-�M�SN<�_6�@9�.�ﮆ�J o���!���'K@�Ԁ5w�֝f��c�s��.Ub�9<��f\Vӹ�ǅݱ�n�'��ߜAC�~�k�q��L�N����c0�/��zʭ�Veo����b�i���L.���=
�s'��e���q7�o�ޤ{���@o+�9��� 9Mb9�����`m��<��p���U�x��%��[�����֣���_�xU#(�pˈ×w�z_/�A�͍�v�m��+��I���p�65r���ٿ�w��ņ�����y)]�/m�4�Z�f� �9kP
���
���b7<B�P�u���B���ǹ[�R��\aa�����5D�r��d������wz�����%�|�#����CW
|􏴤G9�����;c��e�;WE�vk�_q��&�"�U��qL?t����jUC�I�(���ɂ���m����,'��oU,���p�O���5�s\�dAF��m^��U�'e^���q�8������t�Z�g��t``C�]1؍���3zwG3�l@�=�q�3/N۠N��,��
gx�ǻ���k���=�Q׵�ٛ1o���f0t�/5�!֖-���5-݆��o��CӪ����$�f�;PW1$��j��^��n�l_G�VH�:�sa5��Y�h�-魢{<��W3����NR�y�_<W.��we�t��R r9BQ��c��}�17XN�`>�� =������m�+T����2�XK�[ww@�g�3Ǣc|��O�T����^�K	|��s��T�ɘ>3>��u��Z�b�M�C^���ngI����]�	��Éz���=�����"�-R=��+�ۻ�f>�E[�^+KFNY���p(��R�.��ާQX�MZ��<xu�?£���|����i��
]���z,I��uǝ���k,��������D�#�fP�'%zs[�pbm�g�����Sr��-p�������xѽLF��GUԗX�uW�UM�8�ot���8
J(]���\��ɚ0y���?�N��{�u�)x�d?�.�!Kj)��i�g{Ä���>W;��V�[�v'l��b�z�-#JF�F�On�<Wlfi�a.��B�Ή���
�'Ʀ<�Pq�ັu�h�o%@H��j�|�ݻN�l�˃y�7�dmT��A=$���^�b��Ɛ�ԡ��ea=c8�M<�=���x�@�%,#�~x��pfD��_I�<�7}��P��rp�Au(]�VJ�W�g��	�-�Ft �ͼF�JٖXv.�eTI��ʺ>��"#q�{�j�H�ʶ�ӓ��h��#��ck�[�<����*w�H���T�ٛ�J�k��8v���d�Q���{tz�3���<�M�>q���홀�ؾ�ų��Xc����3�����U��K�ω��p�aK���Zzr\�Kx��n��MPV��j�U�Z��0�K{[u�c����A�f�劧�S�0pc�O.��������P^wKOU�r��s��b�Q����͖�P�:X���T3���.�er��{t���@�B�ժ�e�KH\���(���4�$�S��D���3Yn����~�*l_n�r 7 Y��^N��ϭD[��s�q����m�{���t���sQ[�],5#����v��ع�bٗ��TRHl�B�˶�u��l3���q��5����&ﴈWR\ڮQ�Bz��U=�Az��t���=�
�Z�9�b��]1���O�N]E�q�����ARsx	�Z�+v�Xs"Ҭ�C��ɬ�r,��P*��t��%��c�{�,�).��k��a��6�n��o���Ic��3!��S�Y�������u�]�M������3h����H�J��%U�wfMx��=G����kVer"�i��:Xs��1K&��Gb��og!�m{۳��9.t7V�g�"�5;��['B���bdX^�b��_({p�yX`s�T��ܢV�C5kX����z������ȏ�X��J�׸G('�^�a��6��s"��+(�7��:�69>�p����5x �kC�ۛ{��k{b=R^(�E<��ܶ�*����*H��Xkn�/.ҝ���S95��gTn(�J<���� ��|}*%oZ��7*�ds�^�!�D�5�:i���T�EqN��h��m-}�{��/�Dl�A��(>�r|��jT&v=��U�	e��U8��x��A��L�8� �X��g�w v0m�i��Q�fE�g�]~��<�O�ܯ��1����5{:����z�pw����2�F#"�"�ؒ�rj�e���k�f�ͬ�?,���#�\���ɯD�06;5yt�c�/�gdKwF����=�{�E�G�N6�=�	 %JE�Z�|�u�!��V��.���g_Y�_I��fե�����- �2t��S���:��z��UNj㱺)��]��3Y������O������Dd�(���U,��Ƙy���Ye�D�~���V�|��6�E�M������2����q��q9T[T�S]��3�r�[�#����yz}>�O������{���Ƅ1��A����ޏn�]�,(���f�gQnWk����XX�*��A��54We��J�O�`�g�࡫�F�9�4��"�K��t>���'*�q��d)��M���k"�t�{�:u���@We��Oq=��:�{�{&I���TF��^���Y�[�
��iis\�2;�1Q��K{����}>�����n�e�U�bq�M�m)�icuء�����v��Wy+��=ۦ�RO<��0e�FG�/6�VH�W��G\��^��Ӻ����[u��GF؝"y�v�vK{B5��nL���ũ��;�Ƒ�ۘI7�l\�]q��\W�����;'-�/�b�����|e�G�m��#�в��̭[�=�6���:vNb���nL#�hėۻ�i��:���!pm��:��4n��,������kA~�!\��.^���B�m�ALr������ٵ��03	@�p�5�>������^�lt���~d�\�#�ت���"�zmd�H��7��mˬ�'˫P��7˸Ľ��:DQ˕����w���r4��i���Og� b�]W�i޽V|�T95b����,#&�׌X5��.s�|qu�5�#D�0}�K�<�����oጻ�Ѧ-:Y2�zs��,=�6���ӽţ��^6쥹E��t�V!�)�Џ�=�T.i�Vu�,�dO���w�A���e?�v�/n�P�f�-��;l&���h���4nJ�v*�5��Cc�m�P�3��uvEeDu��1��-M�^w��`�^�w����DG�^��K}Gz����.ew<�LUn���/Na�550T�e�i�B�����H=��L�*f^&i���b̗�Ld]������4tF�\��5/1�o������=}Xz��{E|_q��v.�vx}#��N�m:��Ӎ�v˖�ӹy����9��'�[ae�纑uc�Ŭ���2o(�t�P�uq(�q��DWd�����W�%��7�_9�*��6d�+�	�uv!�Y�^b�ݐ(:fE5 ������:�n�C����>ڳw�!�F)ҍ��iS=�ha�u.�ye�����]x��r��pf��̥���[y�gG��H����a$�
�	F�<�x�ڏ�q�۱FE�]8�87w3�y�O�Ҹ�=dƳl���.*�oh,k�wuy��E����6������#���_���V��+��d�=S{3XӏDdc4k�\}YNȰ�oGD[(�Ա���7������.��Ht�9����ݍ�ce���
t���,�vU��R[k*�v̔-*/��u�L�yIb�p�{�&�f7ݙ��Y���Sg����|WK�1]Y��.��n��-k,��ZR.���_M�6Tcvr�V�d���G(Z�'c���%a��w����E2��IȶouՕI�+{�k�N�]���ۖm�]�r�*G�o����
�I�����X�+lERP�4$Lm����I�R�l�u��8����+�)�AZh�i��l���L힍'CщN��"��������L�E�vM-����P�U-RD)�pk���t��Z4�݂�u�����:)��G�5Fڊ�n��n����h�;�������4���T!OI�#���h�((OA�b�x�/BUWݸ(�z ���A�v΍��MY�(*%��H[m�M=.�:@��ҝ!��N�D�j��E�WwwY�))�;6�JD�J+I�`��J(8�IAGlP�KCŤ4:]=��29�_���6����r�9���ʆ��Vq�E9�]�ݕ����=g22D]���;��fv���gn~7�U;v5�u�	&f_u��?���)����3�+5Ec��e��i�@��s�K)��Z�X��g��N[%��e�.�)wY��(���d���,&=�����KԻ��ڽ���c6���Y~O'v�������Q��`��������?+�oK������],Oۙ�t���o��nr�|�C��.y�|�#$�v�=C��y�[,�q�]"����S��Ān�6�S�-'�����Oy����V�-]�V1�p�F4���{62olR��f�6�'�s9j��s Qݺ�HZ�g���|�ď>=�����=��ٲk����x����[ٖ8�q�3<m�{�a��0P�˃Mí]�R\a5k�����N���g��~�@;�
A�=�c�,,�����{sLu
��D6'}J�Tz� ^��8�o`�B4P��TYy�������!�`m��zij��R�����^uanKo�W_��h0���J��nf�zm��2.fh\����ۣX��^�2�awT�ah��1>�.6�W�q^l�����C\�ƕ'�w���S��g)Q�����,�4���#����C��,���_+������7�t��]M�A��j~�&ݔ��졠�6���jl\�Y��M�5�^���1B�R�r�1W��h��pOv�QR[�T�5�w��b�|�O��YR��S	�y:�5|��s�JØ�o�'=y��OW����:[`5Ty�u<��бJmqL�׋��~����b�zv�椕(8���	]�z��*���m�Y*ۮ�nV��+��� @b3"��^�޹�/�P�|�1��N�R��V��Vт��^��fA��Z�96L�E��-#{!��S�Ӟ�A��$�m��j�W�O�*�=��/S0��+^B���f���͒�Gg�b,���_�x=�$�q�� �S	�>�i�et����?-��5�n�&�v�nڧ'w;�����a�q]ԑ(ߝwH[o�;Y��ġ���������|���`T����TC��^]l����lp�y4P2s(fwZ3Qࣲؒ�ŀ� q�86��C.��.��Խ=t.�Y�̼��\�\�7��FO^�]*�t÷]�J0cy�	�!7yY��I� "�v�ßknN<L
�θ��37v��㺵��嫉Â�
�V`�����eP(8�v����U�O��s>㺲�F<��٪���!�b\vE���%�t\��rᘘu�"3]����X�.zA[L���pWf�\�@٫���D�<_�H{c�49G�o��ڲƾ�<r[I�ݗ���B���/UȰ���F/�j�቏>ٟ@Vf��ų��z[_�������nm��c[��ܨi�|����d2/ B�",���sf(	�m�Spz�A�-�7���~{�i4�������+��W�Nԁ���~�4��TQ��p�31^E�&�Ӵ{M:���d<bOJ2������Rb��}��UB���T^���?jo+�mw|caF�UՓ^ཷ��� ���zG��&�T�3}Ҷ��	QĚX/A�SPS���jP��6�s�['7�ly��2����*��Ԗ�����_�	{���!�ڣ�!(�a6�ZF��=0�"'�-��	W�w���ۓ�K���sq4$�Z���=M���-��~\�����[{�v�����\w�y$�]V��tc�l�b�8gT¶Hxp�"��4�3)>t�Y�g�^�p�W�U�^��Ҟ�ɗ�֫�ڟ}�ƕ!��S��,�������

a�vu�
���V�@��Hq��a*ɥy�U�7R�lSS�Y'�!�ܾ^�#��4龕
�� �Mˍ �{�� ��P������^8�u�u=�e�n�����q�ig�w�=�6q��Vuf�����5����~�����_���oW�6+T֮}eAM�<����\���`"�e���^��O�C�=��F�S; nN�ﳒŚ�a^����;g7)h��>'q2w��}�7ũ��w��7����u�*<��nیf
��wA�������y� �i����]���wH�FD��S��q/�_o�v��:�������ډe�������s����p1ȼ=Ti\eT���w��P������4���V�>m]��E��(�쳯{f�S�A!��s�>�f���M�	�-J�G�}l�ʲ��Q��H���\����5�r�t��Q*�&"1��\�-�A7�͹y/��T���T':Y���;�����c��h�%"�CE���{����ƌ�^�g8�y5���v�ў�k�����4�+�^ �R�h�#�DIv3�W��%�;��^?h�<d ԪD_��5w��Oh�ϒ#n���0�9N�
wX��Fm�[�%u�|/⏮}o#�D�ĖM��iȷ���ۢ�m��oHa����jȥ.�523�Q�M��\��/� ٿn�j;�0�.y?Ee�;@Y��T�Wr|V<���p���_����S�BŌ��>��Va�ҏ0�_�=��5�(��n� ;��MJg�x�k�Z�߳����v2�Cvl����PnH��s5,�+��s��a�/��y���l˻d ��4�B�Ni�§���Y-\���={v<���yש�۶�^h���-75�}=ƽ���UG��<��t:��l��,���t�&��%�m�P�Y���� ����>���� �c!`I3uJr���D�X���F}�kv���B]ӯM����޻����D�n�&o�K�%��rV7���v�Wj�H����	]J7�n]D���茇{�b��|.1������`!����!�X������NQm߻�M�q�ͱ���&j�w�ϖ��@��H:��>���>m�p������;��B���t«��)���՜yY�6H3;<m�{�`8�+*�Utj���m/=�#�pG�_ɥ9Ǥ5��)��9Pl�y[�4l�c2�<:Gl�n��b���i�W� r��3t]�=�w'�@&��M��p�޼�t\A}�ͪ c������k/�7ʆ������'1���1ZtE���#��{z��mZ���/����E��]!)�ў{ǻ��YVb����I�.�nR��G<� 5��9�.�Y��/K������=��|6|��أ9�)���Uy�u��	��@	.�ȍlY�j�u-S�c�
/s`R���^�)W�^H*���:PFee�R��a��4�#NkV�� ���d�Z����]d�܀�[�ƙ���U5�us�>���Aެ��r�G�nh=�~����o&�����.�-��e�.<��J/9��kmG��ѷa_vtZ�b�th�K��E��7ؘ|6&��ft�u�T���*��0�\�j�ܴYS���v�=��?qX�io:�u�.aw�^o,ön"_6�H����V���q�V�C���rF��,3�Xk'�XG��S�S���޽>J{�I*`�zzm��ͭ��y���l��o/N�r]��X	��-ܐ9U����S?3,�ռ�v,�l<��[�_9�w|k/5�w��
�J�.���}�4;f���ԛ��y��+�e��ў�!���xM�'�J{s#{ue�akSl�f�c+	�Ȋzܡs9@�X-��7-��"!FEgu��^�.|V�~FpV�
F����]t��8��/��dXj����
�m4��G�������������==s��{�/O^�s;�E��@Vf��{qjf��Yuj���hOK�m��8���`/!���}/��ǡa����Sds���-Ơ�x]xo:�~���ʓO+u��p�����#�/��R�u�,��n�#w=t�+�͖]�9O�LB�>�)��i��J4:��$��j���H9���4��ܶ�A�;���Ti�W�Z}�׺E�kU�^v��|KE���g*��q�u	�����W:��&х<S�[�Զ�,�u}����Y1Y��ٝ�5�nR�]�f��¤�*����RC{��-�ji����-��1�ԣ��ln�ـ;f�U�V��HN}�s{J����ho+�,��n$m�<O�g	�x̷r2[T��x�\+%7z�uV��3��)�*3B��Yd�tNe�`r̪��;`y��U߃�kJ�a���]V��»A��g��ۼQ�E��&�Q{�$�<��j� <�M���"L��F�n��o�F�4pj�>n���<��]����X�us?���a{㾂����/s�<P��~�������m⎏7.4�k�.� oj:�ݶ�Gs��F)na�c���ݜ�HC�H�6?D�n�79C�+�������������L��Jg��~�fd6ٟC���L���}�,~�����������_Xr�#��;OvƖ296l���猁�Q/9�~�߫嘄�Iuf���Ʊ��
�w+���z7]Rr��A�]7����|������foT�$�&�t�R��Q�[b��n�2��9��S�kagyM7��knb/J�*�+{�Q�!�^�}��b��g:�e���N]`�d�E5�����ɺn�c�ɨ������ly� 6����R~W�x�� �'��ڱ��o�׮�>#ۀ�t������g���e�1��z6kؘ�SMeN�s��EW R�����op{�Y�S��C���9�a�c�[��S���f��	7�W�a���8ۭ�z�"� �)/.�F�wd�;]�����Ov`����w��4뾡~癒�H�Q>�b�ϒ�T	�j__3{;0���+��s��0k�;�r�
��_7=K���$��o%ł��##�x�t��eZ�v������o�*_���*���1q.4��P.K,w��h*�jV�QxVL�V��t��1��L���Bx�Y��m´�yg"k�1�{9+�JI��4�U�k��^σ�6��A=�����7n��5��/�I��XtL�����NE�YH��@�*ڳ��˙��E�BT���5��-�(q�:���Z_>�ފJauLRֆ��h.�y�q�9�=��5���y�̤����ݗ؅�N��]�v�cT��)6�C������8V�fFa���l4�	F���\J��2��T�i��u=�o��=M}���)x���
��7%���ݰ�C�&�e�y�X��#p��t���e�]\��ق4ϭ���3�}9�������Y��0[���+,�k�;�&׼����YOgD:�w�T:~���1FC8��T�o�^}��p=gI���;���@�*|�Cq�_�He Bޘ����x��m���ǧ[O1ٛ�z8����J̺]}>:��=��g��Z��;�-��ʤfl�R���dF�Ǻ�X��-sY���o�����
����MK�2,��@m,2��$�������b����7+G�?��1e���S݄ֆs�w\4�Q�� % P��\��n�~���Nff]��(*��;ʥzk-�7���������W�|��1�we��]�&��n)e�;��T���FH��46�k,�C��Ǣ�o�?[�����{ߦ����D U�� TQ����i�l���Ҋ�����q�������G
��2�0,2�0�� L�! *� L�0��*�2�D �  @@@P~��� !� !�|�E� C �C C  C C C C�|9 0 PPPa� �@@�T �A � �D � � � �D@�K�!�!�@!�!�@!�@!� !� !� !� ;Cª�( C*�� ���2�� C���ʰȰʰ��°�ȳ
����eXo%\0,0,2�2��C�a�eXeXeX`@��U�@"?������{ߛ��*(4� %(�*_�c���������������������*��!����r��ҏ�������������R �������
 ��?�� �@{���A� d��������� �
���7�˿q���`������P��>�w������ ��Ĩ�(�4 R�  H ��1  R�0���� J��( I @J��������  @��$As I  A  @B �  @ ��+*�+ B@ ��2�� ��@"�~����������*(��@�P*��?@o����� ��������>?��D U��0~�������y����'������c��<?7� ~���O����� W�!����E{�=�� ��g�L��a�80`��7��y?O��x����C����B ��<�C�(�����~A��������P�H|Q }�@�?�D U���{���I�W���?@,	�X?q�|�����|������ ��{�C��~��>��?�8=����?K�EE`���w��A�������{�����~�������e5���M%ԍ�!�?���}����#��/ >���������*B���*EB*J�E(T�JU*���D)*�
UB�R$�"!B�J�*�%�_v�f��UB�T�B���jJ�IhiR�U$(���$EU
"��*�ED�����R��j�Q*�R�E$J��RU*J��QEEJAJAMD�*PB�JIh�T��`�(R�!�*TJ�D��b��J���  69m���L��F!�ңki[T�*j���f�J��CI�Cm������Ec,*֭*U��SUFҦ�
���B@*i����i�  �: �B�
r�CB�
(u��СB�
 �' +�(��d�E�+[lk5[MK4��-���6�����U[Pf�-��ISYJEB*5��%%8  �m4Ԥ�km�hh�Y�̨6e�6�$�U��ղ����[-m�����#AV�m[V�kMm@�Z�ٶ���J�k%���"*JDE
�Q�  r�-eQZ)�T[5*4��4�2تjdj�ɚV�*�6�UTT2jـ-��0V5��ʙ#F�6�%EI(I
J&�#�  ���V`�jTd�T*6[V�@�Hi���ʵP%Z�jM�Ha�
��emV��T�(1D� �
T�F���  8t2�V��4��Q��0J��`(i�ű �
�J�� 
	��%��6�T-IR�������J("�  fp���5�@,�R�P5�A��M*�Sj��D)eL֨��J��H ��E ��Q*�BP%@�T�  N  :&V� � �` 4J 0kAE�` �`Ѧ�mL  5km�4 !��QDDU(IG  pt� mQ�4 m  Ah( "�f��, )�XX@��� MZ�  �I$��jT�cY%*ۀ n�B��S  ���� �چ֔ �X (	M`P Ѵ��  1�� �  L���;�E@
  �=�2���F�2h�` #@db)�IJ�Dɉ�&C�FL&���hU=�I�@m@4     ���R��1��10 �#L�&�L"�2M!�Dd�S'�bh��f�I��d�F��=4����C0	��%�n\�Ȇ6 sVn3Db)�y�K@2E���o��W��W�-�w��u�BB���r���,sw����(� �@ (�E>D(��'g����~�����0�:�a�(",�?r�h���	t"������mӕj\�ϗ\t�E�G��cu���f����~��u,��o����~o�mF��d�j`�����`-&�̊���N����v��j��.���ų]��$l�L$��{��E�x�r���fު��m�+@�U2�j��[�X��4���
CQ�bX����i�J�Ʊ[#XIGXʩ&�5�*f�B�	�VE����-ּ���h�W��n�-��*�!���$Ɂ�cH�y�i	Vu�qɹ��D �c���Q�Fҕ����j�Y�p�L�+�e-�k2aN���
)�F�mބ��Rr` Mm�ƣ�R�Ŧռ�b�YM��ur#F+qR��6���.C/,�N��P�SS�@�)�l��miN`AE�������LoE�{00°1�91�$1K�f�`�sC�Ÿj݄�n�n�[F���0*�2�-��+"�R� �Q���*��yR�Qɥ]�I
J��j&�ʼ����
q
qAU�ſ`zoA(� ��q٣@�MN^�v^Ò��b`6�0|^!����j��l���(:��X�v�uXA�QX�C)�ڊ�+���X�`�{`;ڹ��Bǡ���T07X�-�W��+-l�s ���v�8�%�աky�uR��fU�X�SlU:�4����`��q�&S�+Z�t�mo֛7l��ط�]���9M�`�V�7�m]�1_�^�����R�)f��"�Aϋ�:4�F�����b��ِ���pCt/bӒ6(Dnm#p�+�P�6+��\�`eͨ��v�"lr�n��HC�v�S)ؠ�[3��ӣ-L;=��(�˺'��bIKU]`��a)X���tm�YK�����0D���C�m��r��/0��Kq اY��J�gi >�o��nڭ�;)nPm�F�1�ܭ�KS�����%J�E�EF��ƣ�e�xs8�Ux��jHb��V��)���Ӧ��J��<�QJ�!Vfn@��Ae/.^jl����U��հ6��(VP�d�D,�'j��-�5bb� ���(�b���I�X9x�[M7��FJ�-�e�A�RJbeU���``�M̥ln唬�f�B�0�����h��2�ix��R�6ؽ15x����ĤG6m�%aQ+"/YN�eb�R�mVnK�M1";ge=��tZ��F��Wl0�7�H5��n��-)R�CR��%��yf�:�m*	llۤ(?��.���u6i�z�S��N�X�Qm����ǯ&-Z������3M)���P�/*=f=�eDs�kRˡ�˫�����-lY�' ȣ$�ʘ���T"�w�n^���"��ޠ���nR�����Ɂ��X����PƵ9�S�����{Z����4�r���o�W$D�i�p�D�H?l�Y�!�9��j��J;�;4����A���Y2������5��u-]��ց��3s;qR�9��� )J�a�T�Ё�2�GxYǶ+6Ճ7r��*m���F(�O�B�ljӧM<q�NX�p��Z����%����6�Q��ѫ&Gr�]ӌb��m�-3�.Ku�X{�]�,���,�ut�����FQ�eh��I/V�+P��ҀTY���v��͋3"��:�U[�z�ka)�S4�Ħnk9�2�)m����:��
��ڋnjW[!cjM	�V���m=~��J[6Z��k'�^�ּ5e`�H��W58��7B�;��:�E��E,R��l�'[ݣG+H���d8X�-��A�w/ND�z2���5AW���e
��
�N��t)��+[@���x�Kݤ��qw��zr�ji�ςȐʴ�X)�Ҳ�Z/-��j�p�H4a��2Rg#�cǛ��opfф���N�=��S7�!�NMA*�݌٦j4�]Ԕ4T����X�$,f,N٥W0��/Sŵh���t��0,��)��f�Z4����1 f-�n���Bl�Xj�)X��h*���q�X*p�����4j
��X6S���yfb_�@��ͭ����[��Q�u�K)�ek̶0�Ql�����2�t+�q�ԖƆ�'U�\���3wrV�8���Sb&+J��
��1�j=�LZY2a��fݶ����#��AE�Ghn��ۼ���"�≋?4Ӊ���NPI�4�d���2��*���M�I,�!�lֵZ��/R[����Ňkiag�)5x��Z���v���r�V6�[Cq���#,�����3�4�e<�L�);UN�Ek%KLM�`ԭL�j�*��H�7�1�f046
��q���F��t�D�@�w�)�5��Q��T� �IV��
r�T����
�,eKOe�,����ƍ`$��!C,M��$�c����y�m
Sm�%جcf�P��*�;y���Á),K�<�v�����?-�[x�8�6��rk���p8�v��e��T���-L(�f�T��3&խ4���T�j4���N:f�~�(:�z�U�w�ӊ�@�KE�**S�� 3w7w�,S�1�Wz�727��������7H!�䦶LWX�k17!��Wuu�Q��\:�a�,vUf^S׵	;̂\���9�����3V́�I��R3p
����zZ��6���1��ߎ��{�S�eB�ڤ���E�P[v�I�0����)7���J���'�/����Zx�)���˙�v��������?3��l
�����P6F���6Z��"��,����Z̘����V�v��WZ$���3D��"� �����X~��B��T�4����/eǷV�MM̆�w)hґ�e�k[�l��:C��q&�Y�� $����8�XXł����i��n^��T˅'oek��[B�Խ�P�6�Tx�4o���q�'�P)i��Ӷ��e�i!�t^*N���X�\zq ƚ9QM�k��
!,M�0��G�TkZ)^�2f�Or(5�R��Zp't�Toh�����(��=��!yV�wQZ��鲭�o*i��hz�f��4E���Өnd�y���iɬV,��h A��z�K��&��/�ZWMS�i�ԅe��͍Y�f�$\z�٩��U��{���"'Nle=���;�R̰��qk	S]-4��0��u��Y�R�M�Q��^Y��7�l8a�^�n��̽vFa0���t�-��4k~IŴ(��;��c�CB*��i�钊���B:f)3!����q٣F���r�����ܖ���d˴��h^��\��t7N���y��PR�(��Spѳ5eົ����,CKeX�X��Y�c��!y���`c����nުW�� ���Cn5AE47�)��1+�e�G��^n`6\4�۹`g�E���^�i��[E�5�a��t�
`4 ����lR�#DX���)YX5ʓ/*���$�vUv��y�jG��rou$�K1�/�u��qj� ޫWL^�yBܬ���j0hNΣ���j��-�r)�a]nCr��n��P[ 4�KH�f�e����2���u�ID<l����ɹin&i�Y��o^X�HRNZ0f�iи�h�p���b`IZ,(sEnхI�fVX�w�0kM���� ,�[b\t��b�H�,�W8�{�nق��b 2l����B�X� a��K��t��Y�n+gd��2��*��MXfh0ժI�4L��]L�X�������b�t�Bt�`�S{��CTP����0�c���Z�-V	,���t��{F��.�tM:'G&â#�+�X��3VM���ފAZ�b��� d�U�w�I54������	����D��@uT�B3�k5��j�׶����j�c+m:	!Enm���1�Z #B���Å�wԖ�Z��CnEA n���]:YW�(̲e;X�Ggm�Efյ�ۗH��D�6���*���L��`4�7�^�a`�70��n���,F�m�2��ٶ#-ꚋ��nJ�#��X���^��E�2S�#�Ĳ�)��naL
GX�Sn㙶LE�R�a�Mc��j�,�i,'Zx&�jLA�:��h�Ghb;�.�I������N���X�)�R���n��Ǵ����	�"��ޛ��M��Ӫ�!�2���u}^���-d��.�id�:52V
gP��J����)�:(]C�TM��η+5Ӭ�u���VV��.���1i�D,��J��t˺5��D��R�p�Z@;Q��ZjAV�4H7]��I�m�%�M�i��n���[N$�,��ӭi	Ֆ��+@PL��%Y�pU��+���(u��t_���3t�R-S)��B�A���4�M0Q(�A�7%X���l̼�K�������vi��ڛ����m��F�%��V�:���h��^�jL���ݚ��wOs�	)�L�+qZ.���nP0���hx>rY{AY��n= uz
�R�n�v�e ��̖tNu����Ӂ��hTf�ٮ�w^-��Z�|��i��Ǒh�O^�r�8��S���ݹb�"�5Qѡ���j��Z1]���u]�����@	�V��@��B��(�Y�v��\*��M���eM�D���u�o>�͈�OI�S����pX�-D�e��fMh�
�iՀ:*%���A�m�D\�l�hU�����a�� !$֬E���2�`Z����+�LF�YZ0R��+÷���T���N�����C�|�n�J]4�^���h�F�rb+~ӏ/K�OA��
~�����)Cp��X�%e2&�n��ϙ�� k�z�J{�����Xs]�@y&3z�Tra���-��B� n���9�-�зNk�P�Ҩ���!�JՖ�� ���� ��fd��ci�V����9(������(�ip7�i�pB�ʚNS���9�A�aa����J����rn(V"�*��b���;��ڇю�b��,�Sk@V�2T@k���T�z� T�T�, JK�ӖsC�@##9J�����f���-=��h���c�E�0X����X�p!z��Р�&�*Vht��EA�s"��@y�pm�u7,T�V�Im�2�ѵ���0 bʖU�������ЩV�O4���

bTh�݋�r���/�Cz�}�]��)��A��	W��0̱C3(��D!h�z�[��ٔG�Mͼf7x�e�"�!�ynTk[Ae������8�ǖ�	QD�M�K�h�����ն�*yw�Hn�����/@�٠�A.ҽB�ͺ;�'ʯcu�n�+*A�R�I�U���Ƭ1�I�c��:��bU6�+�H)	X��+f7�e��*ڈ���V1�SQ�݊ś��;@�Jilf��)aT"��=��a�k4����j}�ʊ[�e�D]e�J���F�xuM
kI�d�����3u[*%�-۔���ܽV��}h����zD��5#BFRˡwtB&��s@�w�55Nզk!��t��KL�X��#l(A�1�Tq2kq=�����K�ԗ5��ų7B��X(^T�]]�{f�[Sd��4X����뷛�ۑ��h�-�W$ܔ��Cf�F�Q����H;���hܻ1�R��%=.9���"��
]n�Ql����x.n;j�Q��>{VL�oN���B-8�֕��@2.`�Q]@�qӣg*����U�b������j,�IN���!�Z�za%�$fǆ����OH�B�r�[dX[H�,*8l�6�{N�S���I{Hd��RցQ�^��n��^��MV(��i�V�%��T��0D���oCR��Z�^�w^cd��+%9a��Lo-�Hƿ�;=f�m�Zs1RT�`b�'j'{{y���ZT���h����Zf�-���P��It�7r�l�e	LÔ�4m�"�w�V���k��\�����V���@�L�a�M*帴��P��h樵��
�g��P�]{W���@��IZi�L[@f���,Iª=kR���6F��ؾ&�k{A����T�k2�4u͗����e��CG�(�'�ki`����VA��p��VBn�V���.+�-��w6]c�X,��,N��Q�Е�5g�Ч��k��4�%��,�wo�L·� �|��Ya�c1��fըK�KH� ��oU��D�Zso�+h��mިV���.�Lв�1F*b�*^��5��	�7l�Sɻq��Z���[�����w)�0u�3,
m^��htܤ���\6�	��('�j����2VŹ�z"�mS9���,��G�6�,�����������jk���ʶpiT�gd�Ⱥѧni�NָKe�^+xqn� �
�Y�2f�M�54�B�֯�[óZ��KJD6��bP��P�:bįc1
�zKd]�k�m��0§��ֺXl���6�.��,4-҇i^�����"Y�`.�gʎ�n͇4�)z*X%<A�����I��+v��[�)/�;@$"U�i�<'q㺰�P�j�EB�^��j�uk�xX;D7�LLo�3��bi:k@�:�"�yV򝏧z����_���?���}��H���#�O��aѢ�4�]~o˭k^^�����V����W�P5�7�Q�)-�R������\k�,dv�u�����5�L�6�k��;lH;;�g��C�B�ݱx��A���ڬ�%u�B�	7�Gֶ�S���]�m�a�5W`�7����2��]�恆���P.���n'��ֻ&��c���^�ɒ'�e�e����9'K��_m I���"��m6bΕ�o�-=ۭ��QtN+��_���H��z@^� t�Ra�n;8y^���ɉ�J��TVa����&Ѥ*l�A�[ H���f͞4�r��I��x+��;/�YEounۺ/.8;B���-q��V�t HѤ�vY�J�;��Q������9ۻ��bԥ!-.ypY��6��C{���?d��4�op�"��9Ǭ`��Lv��S%�[��ks1em:�]BУ�Q�Ԯ��Ȁo�Ŕ���R��D��N��_9�I�&RYi7Yy+��ˡ��%�B�ʯ��/�w���oN��\�^� 3i�q�[�����w</��`�p��r2_Rt�����t�c�9�&ۖ����]W���3x�BjZE_=��y6bP���F���u������Fz���vہ=Q�P%�q�'H8�+�r�僤Q��>m��(��rkڡ�U�L�Ŕ��V^ϳ`� � odnd�Q$i��֥X�xUsn֪U����Yr$�:M�Q�6WZHk� �]�v�q�׳L]ڙ3/:��{zek�\�n��k�\lK����.u��Q�y��u���G սS���$������W�2��k/��vtTq�;�+f,˶�Y�L�.��C���K�b�	�2�`��&�y_v)�;.�`��}����Ժx]M�
��:��ޚt�J)�����;��+
g<˽ZbɕjMRm��Rm�3�Ӷ_=K��z�(M���d4pi��Jvd�|�=ݵ�����r�e
7��F�f�y=���:�5�rz�'u�śdB9-���dK϶��-�@�]5݉h�5��B�En����jW:jإVQ�V^�*owq:�r������L�l+�k��/foy�.ֻ�W�=�XF���-���in��p�	�C`m �������:�;��^e�[�Q�Af�[;X��wAC �:��ak(�F���䜝�T�&�]�X�TJ�&{��m�X�)��}����:m�yv���+��{�fM/�^(���,����ʖ���]�.���t_?���;ݫT]�q�0TL��[x�_������ʕ����8�C�zͮ�=o1�2�{3pN�q����$I�����C�9��]	Y}R��S������ohq��\v��:��S�s �r^c��#Z�C��^��4����-�0н��ݠ��c�*���W�3�%aH٭����0�p�Cl,��R�K;�Ui��Y�'i����w#�˳���-����P�, {�-�5㓛��6��/�r��UЛti$��N��u��!и�HV˛M�j�m�mdm�)vKclT2�����wr�(�Y��D���fW#b�:�zμ�]w�]�i����|;r��U�4����Y\�G���Ѹ��L�f�6T�ڻ�m@��@�ٶ���U�b�/)�q�Ƌg���u=f)�K� *�ő�d4�l�jD������V��TQwW��^�Bf�ˡ�:Uԝ*��ֺB����KE��va'y��zWLX�fꩡ��A����)��3;}�n��fUM�b:u���+��`���藙�/6�ӻ�:�O�����u���$ꚰ��u|�A�t�۩}ަ
3�{�K��S��{ .��_씟�>�1�/ N�W\㊴���e����	�<�s[�o�ޮ�l��,�s2�9.z�p7�J��h�#�֐ݾ�Ҟ�NKƻD)@��Ĭ��3�a劆k䳧>��}X��� z����-�G�p%�W�X`�
�.�������pP����ǎ��H���6JQL�]��o]�;�v�k��^�V��ͤz�^�|����<
��HWg;\���	vd{�u��7vs�ml$nt�x�mA\��T���B�m�p;F	V�����a�\&�ru���H����������4�$.������ޙC\A�VU��sTR(j��\ѬxvV�`�������yJ���u�J햒5�9�p6�`{�ҡǋ5v�˻��(P�r��%м��\a�B�ڍE��!g^�!W;�X�/(��B��Ѿj�������:^FTmpɈ�\6#��Θ�h?��9��.#1�4��U���y�̕��H�R�����C}�!jx,��Z�ޚ���(�ϓ�{Q�.�B=�Q��k;������a��lR�\w;�<�d䑮�ue&���ev:.���EW�$����?��R�(Ỻ�b�m2�յ*�gvSܫu�M������YL7LTiKS�(.�aѮ�]q�aC�K*s��hh'@!5�p�Йk+UCዌ��&��I�#�w�������� �e����h�����������Td��aL���P���s���轚.��焴�JS�W�|kCOэ=�|��y�y�<9W��+��{]�40�
�I�<�]h�i��g*���r��S��A;�n����NR����X5�Ѡ!��J�!�����Ю��y���/1&�]Ip�u 5���'.Rvެ#�Xs�:s������^��NZ&�k�f*�ܓ.v꫉��D�WLU���iYr�\�@�I�0G��1�f$�s��"���A�PX]�f�:�+DW��ee7ق�r�]�fJaw;T��L���'���b�{Z�V94w.�ke-6�p��CYվ�*��%�0�'S�U��×/�Q2l+ �_l�݋s�M�Q �i2��$�o����r� ��RLu���Gt�#���f��Oq��v'��� ��α�gel�CL0�|�N�t������@:*R'9v��ET��v�R�4��+�V�g+�w�4�jbWs�e�}��B��-خ��:Sd1ṕ M�85�S��]v���tX.���:־��*'���l�*�Y��S�q��V�����=
.�R}2Gk�ں$�G�]��$��Vb���v	�'V�����{{}\{'1V��P�}p�J�v"�1�N�P��ּ�"�k(n�b�2��Mv�E'����\�b���RC��Y���<��I�9l�ͧ�t��+��-ֶ�:�M�nH\��C�vQYR�a�k2�⡭�AB��]��/�����N�}���@�5>iH�;{%jmu��[ն��&'G}Ҹʗו�r.<Z�9訛�qN��v��J�D*M_[��:��΋���z'�_c]�,:T*�s�)��X��-dܑ��#��Q\+�=鮕
a�f����|�D��4k�ffXq�1H����v�i�M^�f	۔�i��d����s��+�e�#��ץɔ��{�2�LU�u�5�LWK[�0*�Vb��e'Sr�#o0��G�\��\9����N���z1��:5D1�����2�k(�z�[C��TW;r��z���3v�"���B���G�[�{τlF�T�w]����΁:�+.гM`�OZ|��;�)u��V�B�4.�<u4�]��Va�B�q&�j�~0�[v~9:Tv�e��_e��3[S�rS-�}#Պ
;�xB����9��If�>s`��7g�#N���U��
�ݫCj ����B��g+~u�[{���j��ҧ+���H�j�N��}Oe�t������kWX�/����#y�94�Y|���)mK��mæM]9�WR]b\~�7Y�qﲳ�c�3Rٔ p[���BT��G8�	����(���6n*�9v�FeKPՍցB�����X�;�&�j�Ӑ}��V�35�������=�{-�)��[���d�.3J�l�R=��ҳ�ٜ�T���i�غ��[K��C���\.>���������QR{�ba�.둵4dVq �/ ժ�5r�am<�-�y�O+Uuͺة�J�j3"���d�Ń�*LK%c�רu��kt͜"��z#���:�����_e���c�J�mb0��+Zv�2-�2����2v�-AӬ�vk�o�c�ע�5�&����nw-ͥ�ɞg7K�%'BJl�_A���.ٴ��ҩ<��9K-LfS�&�`�Z���6���ڂ�W�m�	e
Fн�&�*pX�K&vV^� -�JX'�VP����vĳmt�o�Vs�6�� yL�e�DV�0�.�{m�,l�jmӔ�[Ǧ�cC�Iw�]"D���դ&�G�{�|�N$�� ���N�{���;��m�<��
�Wv�X��v?�����(�K�0�6�g8f=���Js��{�
�w`�{���#��LF�B4��lީY���&�M�8JMt�_'�w�'c�����w���r�{-��<���c@�$�'W	F�:]�/����+LW�|�Vն��/�u����ƽ�>K#�����Q��W8�9ۼ8��Fn��7L�ѕ�ַ�	�c}o@t��Ne�,H]�5W��jof�9��B��4��/	ƀA��e�q\�ϯ4뿻!S7NY��M��� �>8�Z�����S�d�s(m�\CU�cJ���-4��ɔ���'��`���ލ�:��n���h�B�测�W>�tv�p(�\=J�R#�wh]v�]�rI�� ��2��%�q\�qt����'3X{y�g)z�U)	Wuj��x���x�oc��J���']�c����t�Ъn�n�S��P\���):J]pu(��K���d��٢�ⰴ���
���;G[Y��4�g;������o-�h�3@�xp&'ϧ[e��lM��v���&d������J>8��rI�ݪ��
��_wQ0.��S��������:+(��!�E�����Ȓ�a��7����-�����u��̢���D�tȱ���o
���B8�V����>��Vz!���&o�K]n� ����M�r�*Z����t���E�K�ڻ&Ն�՝Or���*��aa�+�S ���v7��CB4��@s�`�ub��@���R��Z Yn��:[���r�[��D'��,]w�u
y�h�q]:���qm�|{�*E˲7��A%v9��]�͋;	 ��@�d�l'7����x�9�j�y`;��ݫ}e5]�ep� c[�f���igUsT��/"�¨t��QA�6�Nd�D
�Rvn@a�K�`]B�2�^�6�
�����n��; �윯��}/V�ARG����)����:Q闕��۬�z��!+��t����\ߠf��]K)�8YqWF-�@�7xmh²vY7:�����ln�!��iD1�s���:Z��o6�$s+5��ZR��ҍ������9��j�*rRQ�i�e�3�0�D�Yf��K�q�cm.������T�^<�]�n�}!�V�D^wmkT(� J�z��S�U��lԀǅ!�T܁<����c!������]��h ";x̦]�9���~��S��J�!G���^ל@�Qy�j�g+�Ŏn��*Ɔ
��k�w��1vE�D:R�I.�EN̨,��[;���s �pIua;c�#��
,���֔��E6�ϳ��iɥ+�n���˛SX�{��:w��f,}9u�����z�Y�-p�:�Pv�:���H���5�R�����%�@�y���������G�E����e�=1�u�8�:80�|���2Sl�9I[�`���U���|���S�G�ms�v�W(13��Rٙ�NT4u��U2��h��,q�c^0�8��UǮ�zs�Be�WP0�Dp�U�SP-��0ѩ�Z�[�u8��u�H�Ǔ�w���z�O�=��'"�z!��LT5�a\lM_۲J��SE^�[���-�eK���o�xk$�pq�m�e�$[4:ou�	����%�tK+��4�a�(V92��4��3l��:���V�\S�p_H�ٕ/TNо�)ʼ�xwx���YJ��Kte��q3�aLh`	wdW3��Ě_��S��	H���6�y������9��6{F�%�(��/�ZܴLT���������Z��8���i�=}m�9�)^֪�̴FPt:��Ll����Jh�:���YԖqc�E��Q���q���(Snw�ε�;;��4QZ;I>�X�ӌ��W��YD��U�gJ{��Ie��%�[���M�gTc��mqg��]Ρ�u��o\o�����8n"u�^	0#�Vq�X�
5!Av�}�T�\6�Ԣ-��.G��ي	/��b�o:
p���Ktu띁J�slU��W�������:Ƹ����vB*Q�(-��(�� 7�U�}�U �k�2�z�ji1�E(��PU	�N�+{d)B�_n]��i\��� ���p���UjNe�gǇT���D&�-SPR��ԺXȚ��o����ec>n`ˡ'*�@:0:J�TG3c�bg&~��f��9x�{�읍cy\8d����0��a��N�~� ���K`����ļ��7b�N=���s��1��g���".�I5�ʨ����
"J`v�QUE�;�p5�gi]�m��]k���?�]���-Ooz=;��Zn�4�T��؉��w�����o�	%.�\��"M��Q������i��.��d��va��\�����u�Z"�"Y�m��K��ė��r�C�F�e���*V��X�)ފW��$"�`�D���ttx��+������rt_rMd�:���fP�jc�:�<�Ң��f�Y�v8�u��z��kc��e��y�^o)��R�����"iѮ���w�t_ky�v�ν�׺��`����3{�O!u:�*p�|�O�=�w,��w����B��en������vN�Mǔ�'Y�z7�(9�t:������[6�8���V'� ��O�A��hB��[�9��N�oi�3h
!�S2�s;@y�mcF�v��}���ڜ2��{p�nѳ�csG|'-죕i�/�h"��m�˨�tinoۆ(]t�V������"�K�&++eph�,h�H�ݧm[`և��6���vl����9��9O
��c��7�;�u63��Y��W�7�mNn�oVp&��Vroje���B3F=�U��"�o���1	{��I�`�	����
��jI4y�V�8f��v<]g�d�9����oGJUR�v뭓KWyI�w>S��y]�P�'4�a�<�vr�����+\Ɇ��2vZEY蒇����*]q�YR�	g`�Yy����ܘ���[��c���Η�\�i�k7c�iV���C��Sƻ�'>�+��9d����!�;r��h4VmҬ��)��E,S��M�,�@e�/�;!u�����l=�7C�f\��׹*cs&��m�n�ؾ�K(0IК�Y��gl�9Y�9��m`h�^��)4�"�ڢ���%.>ن�hZ����2�p���v��wMuӹ���*s1�"�|��1+њ�N��#��/�v���XA�����*�
��VJ�L����G�A08֞Ӗ9�jZ����7�ww�kJ��o����6_���y��Ny���UyW��D�:�b�Cx�ޙ�Y|��U���L��o���\4��kF�l)����B�1L8k2��֑D�.��oU�W��x��������]�����|~Yօ���X[	fn<]�T��[.`�P�*��نC�wb�Q]���l�|�kȏ�cc�r����G�}��ջ.��O��i�Y�\�ӗ���q-���'eh&A�t빒��h�W#�>��4�;L�e��J
l���`��l.��T�vr���R��떨�-kcqok�4�UI�U��`Rr�b�+��_k��v=�8
���/�7�9W��b^������IȺ�7Ӝ�:�5΂�D�ݫ�G�l�9�V,K��oh���%w;w�r�����v�S4�3&�:b L��g4�֎ @_."�n���໌p �w���a��|b5�{�g(�.���Ǝ֯��]�: VW�����X_u��v�-߻7n�V��<�b8��:fG�6�ݖ�g=�hR��.����uЬ�.����ʅd��9�v�cb���ü���ѥ�Ĭ��s�u,��ӻ&m�Fk�K�f�qL��9q����zj-��}��/l�u�Î��]��`���.ՠf����èԑܖn������l�n�
�@_�M)Y]�Y��=��,7ˎf�־����ƎyD�����߸G]��W
�v��4�w��R�%Rwn���V���t֛�������\���cT��݊���WL}��=�v%#)|�J�x��ĕ�6�!I[�����9������]�V�D�Z+\7�"6��Xf���[��lj��9PNVZ�5�����6��yE��p4K�
��J�%��/�ݬ���ڲ��:o�Z�e.��L�s�i'nΈo������P�A���[l�q^��.�S��EGy8b5ݙ[W�Uy�cڽM�G���Vs�{˶�*�����<"N��'�3�nk�S(+nW/�1�b�;�r���w��'���`GSFIu�ī,�v�gR�>�Yb9�u�Ww��E���e�s���c[�#m'*Z�:��[�t�I�-��B�9��K�Χ{���՘5,����8��Ȋ���=lK�6y��/*����A��p�wp8����n�CM5��c��iXj@�������'k��}ȵb�ā�n���Aٟ�d���+�oJ�� �G��׊�l��0uu�N��ܻt��ڢ|{)l4�p:m���VMp0R�F�#.��m��VD75f�B�c���os,�2ԭm�(����K39��z���]Ir��{M����;zӖ�⋆:�ȳe�*�H@e?�WEt��K��
���c�rv�-��U�(�5%���%�10k��Ϻ��mu���t�6�hW�{�1��aӒ���v�"��]iA�7�=�}S%��xE��Z��nQK3�(w�sͰ���Z��pHd���E�<�VWz+hWJ"�|@��m�ޗ�5�Vޮn�����143n��s�?M ��4\��[ա��gHE�V|�Z+�PDh��[8��͓G�D��s+
�7�97"�V8�'TO>V�R�)�^�r��x��"�+,��#�G�ѐ3j�#��}�me���[@d�n��b����Yy�2�:�kzr}�u�;FVp�;i�P[� ǝ[�����深�����3�a����{��*�D\[]�X�۵5"/�,�����2�-�_�wH�������$Œi�M��WA`[�o�.g�q�Y��۸e�hji�}�ۆigw��%:�X�Գk1�df|��U:�H�!�jƇSӹ���!]z,���˸�]�=�8�K���	j�4i�o74vW;�z��%ԝ
��.�뮴G0":��V�Iaݵf�Hܺ����B9�ھ�]�>z�����.��^&���u�݅�u����� �8<�Mv��]�h�4�1�X��ۍ�3�I0��^v����;�W�q��fp1횕s쁃��Y����D��s��ږ���p���QfJ�m,b8�.��G���=���wW��.�HI/0}�r�vtE�1Ďp���_ti��2�3�u�������8�wB�7Y��˵��P��Wl�B������g0K�n�˃�
�L�M7�$��ޮ<��1�㘞�7�Tc4���n�P�q��M��o�/w@x��%�V���%�S��{*,ⷆM{f�)1n���ܺN,��%���Ђw�����]ʒ�J�wp�k%�a� b���g.��j�w���Z�M����<�9Ǫu.��.A�b�/���"�6���.:�k�`����c?e���V#¶ٵt�|�9n����+�·!����Շ�8w���졚%��7�ޭ��A�uz��lZ;\�UB�wu�u�G6��skB�;���}t����x2���Ư�E��:sw��b%hu'�㛘_U�fuY�y%,�n�<ܫ��rP��wf�I�9���/�g8)���§���_n�6�͒��#�@���6�Sܒ��r��Y7�n!�.N���Z�n�s�J]�l8�u�c-gF̮j�Q��K����uګ%-�,���J��5��(�O��h�d��u&�Q{Y�E%Ckh��;v�_<ћm��OV����E�qB!���[Q�e��tct�=W���Q�����-':X�+��Yx����c.�l�q��ά�V�(�d=�)|iu]�%�݈讳��@5u5�tFLle��w���]�Y��,b��,��ST��W˒fHY3#�V�eJ�ڕ״:M!���Id�������D�Ի��3��S���������"�����JfV���V�'T���쥈*%ܰ����W,
�Xݽ�g�.o�1��5��]�ӋC+N
L*�1���r<�z��H�*�ևv��Ao���*�9����;k"B�M�:�6������W�Ʌ��޺d�
����ͽ�Iϧ>���Tl�n��\{(V���uu�řx2�Bje�Q��*}8�:ky�KP��5���"�ɏ���\ �#(�R�WK�U"�9���/m/�'��˷"+��<�۾8%h(Ц���ɲ�һ�n�r�c0ʔ�4)gF���/+��z0V,�ܰ9��>y{t� -�9m荫�D!��ձ����sa���:̊?��v�����R��|�W��i���t�hQf
*h��k��g/Hbxe������\��U��+=:�tb�Yav6��!��A\;j�V٣S���J�A�U���-ڭ�2�r�%f^V��#׳�;"f�*Α� x��;�JVf�qƱ聞��&k{��U`���&��uz�஖�:����������d�i���jzR�\�
�+�Y��S�2�� ��b��a�Rڨ�5�Ø�3z��@�����aC�'£Wqu�&Hy�lC�}��o�]u9�q����nv����:g�"�i���+�.\��sw�y�9$R���{P��ݍ�E���c�o]#7��y���h�R���y��<�(d�yЭVZ}��]�/�vk����v��}ɕf|�4.��`2Q�ݝ����Hk��,��6FB�V�L%(�n�<���R��š�����Ft79���oP��W���
o
����L7���$�C�"��JV���[ܭ;���R�:�`u��4	(���/���� oX�2G�V��#T��G[��]h�w�^Ts����@��\�Qa�_l�K���4&Ӽ�w��5���	�p�ڔn��[Q�d7RYX�z�sQ�V9��u�9�:��̬EܥEL�0Uu+R���sa�h�����AeҎ��F�]Ӓ�g^�s�:ϝ�X�9�q��Ω���gu ]�4����;����&U_$�5����z�F�7	Y�ǆ�L6��m�o��uٮQh��4s�]bΏ]�E���h����z]�t�l��i�����1cy�l�� 7��5�I�nS��Ȩ�a>�N�or��tH��m�2uJ�Zv�dy���i#˭2V֞k:�ať��E�ٴ����|�lۈ+ԁ7$��B�}��L0䧭 �3n�V1�k���'*�t�u+mX1j�BJ�qf�����r����쁕�]�l��opPb]9MJYc��G,��!�Z��: �xeJS�k��6�:��v�:TaQ_4{��`�V��?��]n��t��Q���Y����*̛.:݊���K�+9��@�R�N#���B'	:^�������L]���b���k�DRs����
��2P��]��ׇ��jm��`�AK]4�.^�����1%�>�M�l�n��9MC����1�a��&M\B���R����m^�Z��yU��ĵ��X&��W�0��W7,���W�N�FVgZn�S�p��|i�e���}��v��9T�]u9�]»lH�}|w�;�{2��\B�@��`'���>?]_Z��37_>���ZB����b�W�n����,@��ybk��%-��؞ܱtʼ��]L9l�a8����j�,[�}�_ժ[%Qd�w,]�S�&6n��mV��ʃM%W��9N�N����:n[��GYC�4��\ܕ���m!*m�Y&s��wS���޼�V���L&=�3${]&eҢv,�1�Ǡ�7-�J�O-f�7�+�O��J2��!��[C)d�r�7WFm�Zч6�R��Lm13 �����a��jDn,n��V{�:���ł�g�U�7��7@4ޮ���͠��;���r�n�V��]
;��{x�n�	��r�;R[�&���CM�\(Ùj�߃��bU�o�L�Ӽ�[Y�Nur��]:-�ғ�0�&J�Ƽ�r��5��@[�1�6�t��o^q.gq�zΣ�$�.Xq�{�����_ƔR�E�2*�f��x�iv�V���G���Me#M�ѦfH%�� ������%�sa�{��! ����e��g��y����-(����R���YZ�|MY��Mb���^\���]n�&���5*-�vJU���zr��=���C�t����H�Q�t�g�ɰ�͕�z��8���	ѝ,_N�o����>�[��a/���jm��,Q�Q�쟬���ۗ��5rU�v�o���[Mt�M;��՞42�89�;�����A�D������g;��b�t6��^���H'a�7+'>��\��}m8:{�!�o2X|-p�cf#ƨLy�h���wU���{��=��ٛ��qT�ٌ�R݅�U�G�a_ol٢�8�S��9V��v�*��Tj�d�����`C��������j�B�«f:��g�V����v�4C��b�>�3o���ab�Q��/3�'mc��mš�]�)�fa̜��u�kMu>ڧd��cC�`��"�7Fr����W�>���ĸR�h��V�[�K�Wq��Ć4*J]���O4C�CA��/)��Yw]8e�����gQOC�z�4u�(;���B�na��f�5�V6�-���ե��}�]!|�����՜�7F�Q:��K
H��z�n*�����r��u!��;�m� pK0 'Z��2��,�-�wv� ��:��! 7��xgE��ڴH�?��_�����$A��!�o�!�����z���p���YІ�\��;tG���;�w:p9��&n!=ޕβt�9oI�7����z�wX*Q��p�%����1�Œ4�	Pl4�p����Zm쎱ZL�Q��e�B��D�P�F�Oj+Y����,�/��˶[z��HG-�r���W1ҍ
x<_d�z�M�6�.}��y7mkp���X��h�1�(rՠ��V���Es{n�Q�/x.�����B��%�Ρ�1���h�1m)�1u��V� a��f��ol��T-�u��2۸�y�t�=���%u7��Ig���+
����O���S�]Ye%Ab6�����]���1�'ς����:)G�	�u����ٜ2��GW�&�t��O� m��[枒�@��+#��+ aV)������Psj��c��0���q-|��Y)�Ú�3�,J�N��{b���s4Y�(^��w���y�����kR�o���n��pƸ�!Z.�$�է�D�\/q$���T^;{�t���-3���8:�e3��<�j�Ok�,�O��ʝM�,ݼ�]{G�k?ʽ�&���S�Ӽ�RΘ�n�3�9���	yʺ��Y�]X�v���������ѧ���m<W�χh	]�Z���8�B�#%r+�#Ky�S�՜�Y��]�7�"�xQ�Wo�R�l�h�DE�Q%d�\���-�(�P\HT
¦3+$��E�
�`�+U"�aR,�a�
��-����)RJŊ,�AI*Kl��B�E���+@���X��1+`(�"1A(b�q��\�"��T+L�@P��q�C�I��H�,1
+X��YQHV+��ư+E��ffĕ��@��1�LB��Zԋ&$P*��f9�r��
,�%�C�cm!S33X�H6��#"��DV�*�T�+m�n%QDEP�P�iR嬈����eb�%h�aXJ �mJѪʂ��UA�j�ɈQ�Lb��*6�eOv~��1�Ô5���9Q���Hn��٣՘Ճ%�����l��GN��S�Σ�N���n�9�X�g8E�������.<]����篖?�����h(׆e�Z+78��<(o *]���my�l���Nw���Gh=���Ȋ
�׆=��V��X#Ǵ)^Aw]��7\���F
�F�Uܦ�z�.f~�0W���w/�V�[��TW�ᒣL��Oj�j^-�ë�/��
!��9�ׂs�p��":Ʌ�a�P�·Rx��N��3[wG�,��WT(1p)ۮ5�W�}�{*�W�/��p-帅?�^F
��칣��\�xۨ �:<,+.���U��4��u�,˫S�\?S���j���8��^��XƧ�����m�^f��K�.�S�!����Ό|�/�(p�9��u@ZT�U[ڎ�ذ�ܬ��Vˍ}tN�ip��}L���_�����7�[��$���P�z�����ǵ�;����i:oh�@[|���ҭ.?W�F��U4Nݥ���0`FZ��9��Ұ�N[)�[��P��e���G��K�b���Y�~���b���~�CN���E���?�-��f��Nn�x��"�U���a)Zm�"���̇Qd=�+�M���"&������sr>�{��Ce�������E�7�p���m�����.��;��ќW�Q}�+ܬ��{'Y9��H�$��t���d.Q�L�m�������q�)���X���@�:�F��;����s:)�j[�GB&�)��*';ͫ�X=�9Ȉ�N�s�~z��6����פ]>X=@�5[��W��K H�wc(.�V:P�N�.�X�/�����A3՜�(���k���C�6�0�� $dwME����`?8C�u�*Cd�V��ؒu�G�/<;��{�l��0N���A�G�xh�4xy����e��9���� ����e�#-�n����:/�X��h�w&�"�Ȉ�-6jTܘT�?r(r �%.Ƴ/���'���=_)�B�.jCg���n��$�9rV��7�5AuL=�K(Ȳ-�OwRaX�����C�$\({�RT/���6�$��u�7���#مtq�uhh�w�����OWʮsv2C�C\�����Î�J��@Z��t��2��[Z��s_�J.3�I�w����Ӵ}?U�q�g�qL��.r��N	���П>T�'-�RV�:�M�Ty�Cs�3��<��j��	����8Õʈ����=��J�겥Nݲ�*�M�{M��#����s�gb�ty(,u�Zj=.�o���n�Y{��u�m�s=V������)S�K+� �|�s�Y��C|sr,�k�-��cH2��҂��YI�w-�nX���4Y�KH:��,:؍�tO	�)Z�r��J�U������\k�H�ۍ!ĕC9��̰=W-@ڮߺߵ�g��V���iT�X!���:���'<�t��K�f�uTVk�9{C3��5n���q�dn�޾�g�-?1Y�W(O��1_U���&=�����K����U����n�צ[?$�^��\.5=�2��,��@������2��ѯ���gW�o�3�Dg�C��uCU���F}�.2/��-9zo�Y]
���|8쵰�f��1��f:� Y?8?JU��s+گ�7XyW�dz�֖z�}%"�o�vZZ\���a�U��G��;S�x4�������S��DH>�R4�J̍/z�&q|��S[ٕ�t���؜�yj�,&�!�����R����P�fs��"��~C����˨�ѻ�%�]n���:8'U8V;�*�I��B� �y��$�ҝ[SV�)�~|�k���V��X@��y�C�t�Ȉ��2䁼��������٧�R��}�oۣ���f=.h��zk�:S;
��p7r�jں~�7����h��瞥�c���WG�_0(:l��6�����\�Y2I�viP��.�4\�4�,M�ϳo��!��{D��p��tG����n��b���J���PWݩ�3��͈��]��|ɲ�o:�!���,d��,L�.��>���~�-Nɯ��v\\wQ�GI(6�!�u�}�ۦ{>��!�Z�c�E��N�_TnX�s��ok�{��,��ߧ$}v]醏�>��/�q�v;���k#�N��!FX�p�ܐ���Mó���}�G�gÉ�\	���^��*�	����r(���ZoO��f�C$\p�rT^d��������X��e2Ј�p�c��U-��7�VW4��=�0�Vlf�@q��4$��LpJ�M�����O�����{>Όd�|(�_5�*9��Ơ9��"Z�\VT��I�-�o��g�J�ƵL�i}��hb��'���N��o��m۹`�H�����l뵪��E�q.;L�Tr����AY�ɑ�����:��7�f���,��l�Þ�f�L�y��`�s��,��+8�w(�<���	�_3�tQ�]E�ut��ܣR����WU݌���k������S��.�ǬZ�^���R��"歋��].�4U�Pr8�+Xe)�g]^��킍oEMpR�J���B����4��Jv%���q��Ps���y`���Ҥ�\�;RHN�9�|�r��mI������(�҇ӴQY (�1��h#�E7�
wN��W�nL����1�c��;C�����# \7r�+g)�Q��~M�ɜJm���w"��J����;# o��uW	>��vϋ�Ѭ�Xok����yv��$pA�,�����s���F�=Q�4��fW�4ʇkz�8��jB������B��.mn�4z(���ky)�r����H����S�x��xfO����f�Z}VʵsE.��'�p*眮���U ���dPf�2��rع���o�s�j
W�=�����lt�q)X�f1��6o��ٿ�U}C��%{���Y\+�����g�o�l�Y���c��.n�$ov8̰�BN����AdPz�JyT|���#���Q�P�z^�2)�����*��h`8y����C�3�F}���8�9@rsh٨�knt��{IF�%�at"Y�y��7Թ�;�XV_��{-p����;U����*RVf;�V����8)�9گ��0 ֻ�B��p\[���8^_p�Qe��H"�O/{�Yh�"Ő���	�t>|H����#�Z��	�i�u�k�w�q\�oe$���+��ߧi�	|_SS݆`7��f0�����5٧8�mur��܏r�{~J�0j�r��!]q�=����c=�F��y�<8��Ac�Sʙw^�:�־r�ʞ���xY�)�_I�j�\>�P\�]y&��S�A�3��]�GZ��1R��z鱵�ηe��A�.���:�wz�ms����b]�DJ����E�i�^EgJ���l�5�F�w�.㈫�d�O�*!��*I��,� ���M��{FNG@��̸Vۿ���Z9!�;��r�ܬw��9@�BU�	��t�r���xLB�U1 ����<��J�u�1}ͼ�#�����0����^�*����+,u����,���}��.9]WQ�U��������
s�{����05�L�MZ��H���1@%Nl,a�?@	�b��xs�R;��O�$r�<�U1#{�6�s��ܲ�� ��B���u��
b�_�K�gcA+�؝�9��Z��e)"hq�O3���9zg��!�E�S���yPYU�l���hO]����ud�]��vWsK��[�.��[�%Ժ��]F��ۂ��+;�fE�ҹS���
��1��jk�W���
9DewΛ5�/�Vj5|�qI��u���.b�<{Jv| �W�KID��xʽOF["SVl{�Aj�϶��h�:a�=c{���t.�m�HQ��R5J�	hЫ:.�����q�8�0�(uE\���l���]t�������r�S�/���6n�����X�����C#���:!�A�¡�ú�J��UG3�Ѝ�����U������ud���;_*��!a3�g��DD���%�"#���O��xf�����{�֮�X�0������D��"�]fU�_�Z�;��fN :�]Ƃ�Fq��{�rT�z��k�$/|���b6i��x��Z�v�����i��-��ywf1.����t'�>> ���H����~�k<ӷH3�=�k
�����3��o�Ʋ�!2�=لF��X�9ڂ�R;��f������7R����j��6������My�������2�,���xe#�n^��tt��-��Y�2��/m�Y�'�ʅ+��afd�;���h�����*�WТ�L�ȼb^��q�$���2iT��)�\���.$iNa��ā���JU���y��6��I�u�+��2]áq?��Y��X� Q<%%��h��	��ʱ9��Qb�^mW{"w8f��`�I=�Wxa,B����� �[6Ĳ�;��BZ�u��i��#���n�7S�Sl0�eu��ܐa��Pdͻ@e�c#7+�:f7�1���]¯��P�>���",z�޹HO����r �D}��`ӕ���H�.�\��{<�<�fм��5�̸�pny}u�P�B";�B�����|B�ݹ{2��4���Tg{)ұ6��f�.F��;���dhg[|��h�F���~�:��F�x�7U���d��
2!�d�=�᫕�R^��ޒ���O/^��e;YD�G��q��ÿM��
͓iW��2�	�g��O�{P�*!��Η����P�lo-��86%{Evϭ���#�g�y:��cu��c�Hq/	R�פE�bqr���6�fl]+��T��b�	mX۞7���wJ�;���Ԩ�-��Q�4k��N'��auT�v>Ȕ��,�8|�Qd���
���������3���j�ΩFt��R�(gZ��9�(��8w�y���<+�\�u�ْ�z�w�D1�T���ˣ�^����z���8�aX]� 3����.��K�� W��qQO+�c(�ț��%*ü\�+3(��c�j��s]5��Nܧͼ8����^�5��u��#���&>$�9ڇ{1p��ͭ�{o{!4�¯R��fP����8`E��h��Z�L���u7�R��� �V�h�'egF2P�|(	�ϰ�v���C�=��rr��RkNv!��.��+%]���M��K�uj�E#�z^�ږĚF�n�����.Uя�=��CXg�{�<hIp�ؚ��AX#�U�Uf�R��[gr�zq,���3�o�Y�k�'��YYSN@- �$8|�9�][�¯$*�3,��[�.3K��a�r��0��\(y��L���p���3chd�+��n�m峨�:��C."�����څ�S���=b�y.��rU�:�/8[���,V�y�6zT�=��49��¤8�.:�W�c;	��+z`c�"*���i�^��Ea����ȑʾ�D�����%qb
��q���/�0�?n�p3�����Q�%˺#^-�1B̲B�&b���H�K�hސ�t�`�f�l'�;����ԧ��Wwf��DDTDv��iɁk�,�e�dk�爺�=���GE������LJ�Hr�-ɸ�Ϯ��j���"��ê>t�[oR�o����κaܛk�w	����aAګ�jR�u��Ѯ⮸�Ӏ>��|��Ï2U�i�	t��Rھ}i�#n�7��2��nQ� ;�n��
wk�����f����-�x�V��)�x8��$�*����V6ܘ���ÍLCE̯��L$���˪+�`a�-}���:�n^�hN㾖���H.+�E�'�é,��q��=�6۰�3�8n:GY�%q��5,��[u[�ofSJ���k,���ˁN�p6z����eP�!}�[�՟����@e����/{:����y[��w��XV]�`W�b��|@y��P���e��log�6 C��ŬKs�fdVC�;�d�-`���Ŋ��l������/�S�l�s'�r4�H�oy~�J7vW���qu]�_ΤGMĸY�)�w�|�����>���Y�����V�oVHO���4�%/
�.�ˆ���,�F��Aĸ�a'mD��4��ܷ;�{!
Q���k42�\v|O����([��t��T!�V�ZN+�m?IC���p{3{F���ъ���s=�6��l�c;Ǹ�E�*�}�i�Vm$�e�3��n�ū��x�TĂGF�A�en}��H��bb��X�'��"#8���@D}�G�B7���*?�_�0�5a�Tc�6o�*�Υ�����z��+C0��T��qn���Z�}sh �7��
�1w��� s�u@Ng7��P-ɍ��sz���W�A^�����%��� ��ӺHOi40"ȃ�qs��s=X-���4��-=�@�G�BV�̥/��R�Wf��Y2��.��G�b���f'{w;s6�ǽ|Ѿ�:խ��ݗ�,St�^gk(��7D��a+�7xC�#�I�`�QbiGU*V�����٬\��;�\��s� �t��ä]׵]WZw;�Ά
$�n�`[J�a�����%�NHmbce��w]��>I:L��x$�\%h���=GU�7�̢ոM���sV4,O:y��Vp�}���:�ݛ"��L�y�ܕ9][��.���4��ʯS�F4b�,�a��)gTwS)l�BM�N�����i�0��R{�V��kU[[;oC�u�:�6��U����S�em��uͅqW�w�OB���n�Ns�!�[y8rTKt"k�bP̫w�RY��[k�N�xaxs2��q!ˊ���{�a�4F��c[Jm۱lb�}�nF�$���U�����-�tԽ`��e@ѽPJ9e]AaƔ	Mᨮ�ӡ[\��8r��1	�y��:�v,Bc�}�(-�/woi���(}݁��,4����P�����̇n;��ec�ǵ����m�+5�[Uř]���EX�4%�غJh��2���0^R�<]>�l�U��T���z�zJ+"�fwu\��G���߷c�U^�{���,��t��w�����f�(�#��y�s;u����1+� /e� �kQg��ݾ���L\�|���^��;C������E��k�	�:-݃n�3�NfV���D��j����X�hz�gQ�(,���zս�s;Sw�O!�:��F���n�>�|�gZ&��MR�i�Co`U�}�vd����(�Z�<�.wrn���5+t�2�u>t(� �)\<n�M��7H6��)�3j�gF���E��P�ZQ�}k-X�]�X
C9]w0"xN9.�x4)*�:nP�� �[���椷4��_V�OU3�"�����LS��2�����,ᮥvT�j�]�4\���7}Q��m���������sU�Ī��[נ�K�`���>Αwpv*.�"��?^]*A��l���ۂ�t�A��}4:=1v�շY9F�����(�ԩe���.�A�N��Em�m���e�P|e)��4��G�A�e��.�Cy���u6�^*\$A�&�!����۽�z�,Z�c��WZUt:J	������Q�� ��,Z�����י�YQN/+i!��"�B����E��)*����1���oZLen�;�>ip��z`�0�f�&d9��]1���_]v��sHξX_c������r ����.��+^&��vFͲ0��_�*�fZ5-R��PR�
�)��ʬ�k(��ʭ���.\�8�I�ڥB��b�5������%B�Da��U��iI�H�8%E%d�������edFVE�aYib���ư�kYU�TD���e�*�U�IX�@��J*U-UX��X"(#R���F0�TJ�7011��*,r��h��EU#l+*Q��G,����ԩEF�0D���Z�Y�PZ���r��1)r�U�\U+feʈ��
«�0F�m[l���D
ZQ*��eQTF	l��!S���+B�B�*B�����*љ��D��R�*�7%`��T5��R��TW
R(V1Ƥ\m���� ��0
�LڰV�I�X(�j*��jz�����v�azO��}{ܜR�!}����ǰ���·1xt)x��=��tT�B*��+�)uJ�s�{�RΘ8��A����/yO1�>d|2��C�>�U:�DI��bJ�|`T8�O��6äĂ���>C��!�xe&*aS�;�<�� ��hu�0�Y���F�插v�8Ɉ}��ӏ�N'��_vhM����&�@��3"��+<d�:��3L��}֡󧴂�"¥C�b�{-`)8�Lu�a��gF^!�t��x���(c8��z��q �O�^���W�������K�f�*�����u,:H:��0��v�;���:I�1�O'>��z�ed��y� t�HV���5`b����d��3"ɉ8��β�aU��ɫ�+��l}1���lgH�[Xbs��$|q��8�L~>�@�>I�����(t�U���bO��s|�^P>LC�L1���'��%egIP��2�*K�Lf�� �O3�v��t����_r�9��f����{��n���'mb��q�`=�q{a�1�>�LC�+�oY:�bAgu�a�Ԛ{f�����I�c;��d�{@��'��3L11����i��iO��G�Ȉ�jJ�w�8�b����	��.>O���$�6��Yҳĕ���XI_SL��B��K���
��W�K�gWLC�.��L1�� �﹒i*�'S}��X
J���3��s���.����}���.>��W��
�a�x��z��q��z����
��:;�C��H/�4�Ͻ�b��4��*c�:�y*N!XV��? T�!S��2\|.)��� �����V�S�xV>���
��O��օ�2T�����:�Ұz͡�CԘ���P�0ۉ=N�ä��$���n��
�}��4��*O�|�!�==�;@|c��1�~q���ޞ^q�>�%B���w�t��%�����Ajzɇ�=I��O�Z��+����b�+'FSq
���c�X�W��<���v�Y�w�}IǶj>��L��mLN�!�UѺ�/M��G�@Iǌ���2� -C�����vϘbc'~fE�3hbz������ �aS����6�i���5
��%d��b��'l��'�$�ju�$��@>�>k���X�9J��Z�#+b�r�lS�%dO�w�14��|E}J-��A�9~�<'�(V��tʻ�}|;�f�:��'�j���0bRՠW�hf��4�D�3���M=/�������˦���}�bQQ�3�}ܶ����Q� t�"��=x� ��w�:J�3�{dĂ��7��a\@�Hz�Ԟ�<���Cl�;�}提� �w��iM���W��v�!7��6�s]���מ���M z��O�`q����N!�
��Оwq$���0��]�d�I��2C����y:�}�x}Z>��Z>��+�O߮�q������Ͻ�\�1�!���"���*���M�3i���ΐ8���S�d��LIP��tCi.�:�ސ� ��w����(q& t�ɼ1���J�>�A0}���ɝ�3q����Z��B�2}��ޏ9HT4��̓\��={�4��LĝL��I��u���SI��f�bbyI��>C9I��t�Xm���>C�;H/��;G.��^5�ms��}��؈� |b�"�Ci+�z���xv��z���CI>B�ٛ�Ru�aC�塌�8��JͲT�q��0*AC�M��z¸ã�gm1���ʯ"	^�7�ʾ��&`|">p�����t�P�=�S��'�OO�����I�{�Tĝ�S���댝��
ʝ��!�bI����y���& q+��n�H�L�&��"����>�σ�Y���g�}1�>-Rq���cߖ!�q�M�Ӥ��!�kZ��c��4��T�B�s�`q���8��y�4���y֧L��LIP��bI}��g�e標�bRE+ğ� l�B��=����Cb�_a�Y>k<d�s,8��l�8��I�+�{�>Nݰ+>I�Ξ2w�4�_9�h���L����uϹ��At�zם�����|���#w=���{`�	��>`{� 	f���gsW�:H,=NٟRb�|�8��t��Jμ��i�W����T;C���B���|��N��01��Ěea�뤟u���O7�w�~s�s��Y�J���u� �\�C����W٪M!��0�;5{N�8���y����S����iSHc��ǌ*�4�^Ӥ���ѽ���N�q
�}�[��}���gV��ǐ��;N:8��7�zN#�[2���|��\�%5���I�̪��_{�J��P�a�P^��w��0X�p��#S�m�7�u�5R1V�oQ���i�+mos)o><Ľ9Cz��]��Іs��"sgwSQ\{�OT��-z@�>���:aXW{�g5�!����H��T>�*�OY���(bM�}�x�̺{`T6���(z��I�{��פ�n�2m�Y=J�L��v��KW�'z.u��K����1>�xx�ô�a�)�i��$ĕ/��Y�K�w�;C���<7���!�J��8��&���tj�I�*m���f@Rq
�λ��t���8Qq�}q��s�yGd�!L���l�`}7q�d��ۦi;߸���k~a��;H/�<9�zCi�1�a����h�����ް=C
��ϼ�:M!����3�C^���@���̇���sT��x����7��~�Ğ�P�;C5kI�};�g/W�=�S���_�!���i�d�P��3z;T��C��$�6���ǈ��m1��皛N�4��'�&@�������1�GNf-�7�ޤ��i4�3�VL����׏sV
Ҥ�;LM>2bN!_(i�����qaXW�Xz{���%@�߷O*,���C[�x�Vp<��@�`��f�>X}w\���皳�����C�o]��q1 �~_WI9��Ud�*O_5f�(&m�@�Vx�L4�$��t��
�hty��t�$��s��}�?8�鏪c"��&g)˯	Q��%s���LE��Y�=���z�OY>5��X
NЯ\��I�����=�i���4��j�g/)8�;�� �&�z�Β�;2�5��q�~u���D|��@�!��޸��{v�2������
���=aS�x�$���0�g�s����z�����d�'�y3�h1:V���`i������Cԕ���Γ��3��*k�q�*AT�]�z��u�����w~�{���_�m;La�����LO����m;H,�<->f��q@�3�R|ʇ���ϴCMaPY�����;@�T����bO��Led����!��}ݞ������ﯵ�t��v��T�6�풢ʓ�I=B�a��~P1'���s&ُ�
��Ѿa��N'��QIǤ���'���Ud�+O��!�Axɟzv�������9*��T�:�m��Rc�$��m'�&X�/+�0jW���R:�P�Z^jx�W%��/�
Va�V���k�;v�;�w
�Cxg�|٤&�확��7uh���D�=�9��mfo8חňY��Tb漇����#��'�s�vޗ]�n.s�d7�|��z�6�^�c>�1 �=M{C\��@�)���&n��1��'H�|�v��&�|�M���|�S�`)1�ʻd�1��>�i�&r�`�u���ꏾ<G�,��U�-�D�١�_���i�g�}*AVE�މ��A}N�\Ci��S�V)��ͳ��t�CĂ����O��ed��Vv���Ĩ|í�:v�dğ!_}��:�����wߛ��>�uߝ_.�����!��%��O�������8����Ă�2T��5����P�v�����z�M`T8����|ʘ�Y�\��:C��a߶�>eC��;��Ax ��w��߮��{�*��_/���@1�>��p2}�$����V_:9����w��ϲ�_�/�uR�<�
ٔ���1J�<��Q�;G`\1�$*�s����7��ό���yˢ�V�c��9Տ�L�L�i���s�u_g��(�.4��(���3��G>B�O7�bZ�g�atBwC�-�^��\hi���U}s�P(R����7��p�� ���4-�\IW�ge�l��0���Oy.�!�q=����P^� ���^g,��N oE����M��B^t��g4�~�&K^[�j%��W��|G�i���k�y�5�	��tc�Q��w��0)YA'5�z���v��}�Ufu����\O�E/��F��>��0D�2�.��t�9Y��G����Dع�(M��%��(Y�� �a�D��zoVA�,���vPmM��ԃ̆��bk�6w����&�lK�*���x�j:P�kٲ�e�����1Qi��Ƥ�m=��R��J�vej$�I.\v�J��U\Љ��v�e��U�;�!�ap-��Q��&x��J����R�k b����W��,����cft�VF�����xm�l�t[���5U��C�Ϫ�M��GRl�}��]�<�c�*z�/ ���X<)��B����q��F,#�\<=);��#(��|Sa:Ƿϲc '���4�F���b@$ti.9���ҁ4�lLsj�Z�����j��6���u��_Z�`q���>H�h��zH�y�ßGC���{iؽQ�˷Ճ�a�u�l�'�9��z��o�cc�J9�6A�G�3n��u����{��R�Z��]쇋��X
Cf���<�dDw3����*:T8��L������m�b�-AH�%a�L���}N!�E���dx��r���c���Ij-k��뜀���Q�1e8�
���W$+�L܋g�ʓB}�*I<��P�}�B�=����7��$8�2`�
φ#����{�#�qGʽ�A�i����ֳW���$zt��_�>�ĴH۵�点lH��wh�X�$!�h�V4ZѺ`�(a� �C�)�x����%�kY�H�v���a�y��u����03�K��%�	.(�wʯ������
��<ۖ�Kb�c,4՗-����Iu��N�����c@��C��uQ]������X
j *����~�緛��L��9�r��]�r� u���y��.Ӓ�:�7�_mKY	����5��Hح�P�s��4�- 뼫F�(ٮx���DX{0![�g���:ѥ��I]v�\I���o�rq�*ZR��B3{]�o
�g�'���6S+W�6"�`��۠�wV�㻾q��s�yf�
�~�4��µ�|T����p�:"��yq��=o�X0x9��F��K��u�z�&�눲8�m3�׽v.&��g�nZ9�=} ��,�g�)��\*v;w��eή��?]+�u?��� \5�]F�;�v�O�\���?V����Zƹ�2��Ԩ��V_B�r��0�h����P+��2��f/���뀶ߵ%���[�Xq��Q��:�Ȑ��F����e�q��?�p?�W�4���J;X�O�C�zmND��)�q���F�؜�嫨���
�]����;z�KTk/��%�AH��H���+��Kzλ���RIO(�wfX�
��t��ĕ�S: �\�xhԺɎ����M��ϮɌ_wjX��lk��z+��o���k�ӭ�Xz٩�1%�^���;ə�f���J�qȺ��X\#�n���Bq:���['�Ba�nV�p6;�Jf�T$����t:`s;�`wF'�uJ�E�Q��_pN�
o���'X�*�u���/��@Tsy�C�%ҷ#7�o�R(��u6�)��=ݭ=�Ha�"x��JGb��u�^&�>�H:�^�X_Ep��:�N�.���}x6�g,�˗�Dp�����;I{O�u�k,���vxW�'����XC)mD�x��C��4?����M�	@�@/��4���Po���u���N�*G8d]�-�������/�o�{��T�f(�}�)��W��j�
��.d�������xZ2��k�����U�Ɨ�o�@��n�LΣĦ��7��O*p�H�U-(����9kfy�b���+\\���u�5��g�a�d�i�q���(M]�fom���"�#l�%@}r��'g��^|���ь��� �w>�Z��v�<A���b|��#�=K������Ʈ�H�/~J�ƵU�2�>�T�E���o=wkڱȨf�m�;�u�f3��MX�;��N�4e�}}9�4����R�}�������T s���b���ʇf5<����V��'�Ŕ(���obPR0�m�o-G�R�G�I|�ڪ�Vt�V� ��\'�Lގș�����s�+u9;-P{������-��o���-�����ܧ��K<���ǰ�9�u7�:VV��Ȥ
/;��ҡᱞ[�Z��,r��>\Ȭ����<�����޺Tq̑�o�5U�fG����aM�6��=���*3�i�b��fB;���tUX��xn!dɈ��!�P�
;�%=j��F1��6���̯�ݻ;{Xחvj��k2I�`�������y�À�.�K��P�7���%�y��6��펛qIk�k�c0� 7s�G\��"G:�D�g�ω�5r����Q��%�t�R�2���u]��G �ODs��`��,� 8\sD�B�_[�K�hސ�t<Ӫ&_f͝�/\�NU
X*ݙP��a������yq��FW�8ܣ?(��c�l��5��1��H�RXE2���FD��I�Y�TCG$�}=�I���=;�L���3Q$[BuV��U��n����34K�d�(z�ϗY��N��=��Lٌ�};b�NE|v���#�°�lIb}�gs��2t�-�"�駗
�:*Dc�'�b���{�m�w��~�1YJ� ����O7U)λ⡠�M�o>;:#K �yPM]|�Hk��b�gk�{W�+����wP�p�b���Zr;��]����U�o��k`DMIH�������Ȩ3��O��\����n��y�+�
�)H�O�ޞ��/o��(׽y0ϑ��[�a�(XV��0+���]�|.�]n���Z�j}��2���k3n|C�e�b}�a���u��
Z�s��5}wk���e�O�����'ݷ��^x���ˬ��#/���5����A�\�:\O�6�_'������D���XÂ*�e�N�}!�n}.��������I
:�8��]�������rq��q]�
�L����5����'��|�K)�tW��E���ޟ_�r��[��wm�V,���>k<C�,)Ĵt��>���0h�i�6��:�kL��9��|�W��r6�̳h��hZ0����6p�<�X������D|��z����]V��q����� �!+����<�a��젹nu�yӉNu�E�ͱ�a��k8�Pb�ɍ����ͅ�A�D�"��X+i�_]���QP�*�R�7{��[V3�%�v�%wS|/���: ��e˔�[s�*��L�kK��wb�r�w&��|�z���j����u�+��A�Z+2���;����T\.�\�\�0;6\�}]�.g\��K�^�[\�O�y7ڗ�> ?,��z�=|w��H�X$�ه��u�b W�2�RcJ��_T>:���\�0�����T|�壘 �wLC�����'����|�(�ݮ�@�ʀ��Q��.8t��.^y��eF��р_����X��Vh��u:��ύ*�!��w;*�{���/��<�g��0�`�>F�aJ�n�X�|1�p�B�<=�����X���:�18��+����|@��`,�Gt�X����KU�/<��A��+o��Q�Ӛ�n3�w݂�ZK��3ƈ"gag��g@�=�AzgҨ�W�ON ��!9��0ӫ�\�Qr}���]���:bCx��F����xO#޶;�����6'V�}�{�;�<ϳ�l�'��?!J����^�a��זӽ�pZB�n_/Ff�^��vX#ԍ�u�ҭc�E�/�mS��"��Vt�"�������V�e,�*�3��<��w_���~b�����S~}xpD����w��鎼2���n����#˦**��.o��Ο
n�,�[&n���π\2:Gg��F��v��������;uD�s��Ji�Ь����PP��s�-�/��0.�й��R�.YYh�w���`R�=���jWu%�5�cuu�{c�e��6n(3�O�ܴ�pl�u�\kr�1�� ��ʈ0�fṖ�Q6�������#ZӡpN��j�ne;���H ��[���b�t�Z��}���?�*�,N��k%f�����[&�F`yy� ^�:�X��X:�<��{�5N��V��̫��;�SeI:�_ ��$����o�����_p\���3s�`�AO���n�٦��y�,��u(��6�EBT�Ҷ�y��X.��<{OgĤ��\=ȼz�Ibn�}tJ��x�)5Sf]�w]1D줄ն���--��,�F�L�w�:^*1�Ǔ6GSZG���g3]d�1Q�K[�.	�*뻃�6�S��O�,ھt��������3��A��M� ��4:Q\v[`��Ѵe� ���.H"Ӳ^��B�dx*�J� �!T�jnj�����]@`�m{��t0�p�6�7�Z2�|����SĬ��`�qͩ�*��IF���ӶHfa�1��k����(ꭽQ��(�l�!u�X��F/�+������UY9��;Ҵ9btU���;H�<�@-��!��R��[m;��#������=V b ��_
��	6.��Wھ��;-p*�H6J�Y�,PT�ҭ ��9O��������zv��y烵+e�W!��]��wi� #z�J5*,Y�!�b�#ƙ�&��pQw�[��� t+r�n��j�:�����]��x��H����<� h�#���Е�k��.�Ѯ�]u74��r6���c��X�� U2�rʝ�|v�kc��p[���\B���:A���zj6NM�dz�t�t::^�u�aY�i�b���j��ԵN":���]_}b�Z�J�l�{�Gs�ۉ�1����.W.��K@��{[�<Q�_c��{0`z�]q+�p�;������V�K�N��L n����N`��T��\}WXj7�	^eL�368@�٢��d��.ҷ�jF����M��O�j��/T������>����˻��ldSgqѷz9u���WA:o����M\%
4���a��|2�3��k{�+���L�4�
�q6�]���*���u6�mfc5������JU�zFn���p94EɠA�ە+:T|!�y�XW;�\E�&RG�g(F��{�-к�O��Di4�:W��ѡ7� %�7�U���{ӵ�����.�}��rr%��qr���Ԓ�B��3��My��L�Ip�uڝ*��s�]!��eJ���Y��[r��s�w�����~!��[(��+X[T+
�EA��q
1A��˂L�YD[IP��*�R*��V)Z¸��J��ee[J�*E�Z\�ĩQU�*4E�[UT%Kkh�1��̭�Z�UĬ��0Ʊb2�(��m
�L�T�
%E`�mZ�AcXZ˔*�+m[em*�Q�ւ��ڨ��kQ[J
"�0��e�2�E�����Tb���֨�*+�\UAm���&2�(���l�S�b���
��Zc�m�V���Q�jLJ��kmJ�L�Z���`��E�Ur،\-�5[k�C�0q��[j`5F�噕c%`��r�Qb*"��l��cR�q�Q\���**�c�5+[h̴�U��cL��˙b�X��PQL��,2@��d�b`n����e��N�ݹ �ÝD W3�-�j��$c�)|VBh�[���ev9nH����B���$��������b]�]��X���2�m�?^:'��Lʈ�3��	Vk���o�~O�����V�Ԅ����F�GC�V��8���:2GH��L*������)W�̬l�'��!:�n��Z�������xˠ��Q�{az:�qk<z;����?�����Dd�=��{�ԝ��O"��hг�~�N�<�@�^NVE��ndL-b9ڥ\Bb1ƽ��k��W>я�1 <Ȱ 8�7y)����'a������#��9~/�N�Q����`Q���/h�1�8�D�w�c>�!�E�=�l�v�0��S�`9fU�")M���M��=CQ���F���|2:�"��\�}���$M.�1@b��pAB���p�*��k�(qf=�3�oe��#1�D0;�����z	>�yJ:�~�rO}�@s�I���ʚ\���vٜ.�#^ڀ��r�B
 ��8i�N��EA�7���?OM��۩�l)8>ǨL�E�!@2Hl���b�ম���jp���(�.�Uy�-��r�^��|�'h�����*L{Xu��C�M�:�TC����U��]=͡1�h}�f.ܽn���3����R��WP������WZZ�F�T܎MX�z�Ԁ��ƛr��/�����P��N���g:6y��Ծ�d崦��.� | {�r�M��q^�������KG���4v[���n��D��Q�ʻ�q ).c�u��ݚb���M!�8[�oʶ���پ"���]���q����dii�y���r����z�%��Y�'Hq�s�.�\���ZU��9��u�m�V��*3���2دT�]��G�)�8Q�;�	"�m}25EE���?t�o��K��Z�sp����
���io���N�l]s���^��Ajt��)?�������NdK���q۩�1��T9��}?wڥ��R#eʌ���ʌd�������߱�4�>-m�Ի�~
43��=��P��VD�i���t���
7M��:q�;Ey�z5U:�g��'[4�yo<؁0�LE助�����*"�Tu��Orv�-U��l��g��RH/z�|�y��^O���~S��k�y�ÅHqx\u-��*5��Sܥb�F�^��v��;9��&��$v�+���$s�t�����Zj��ʾ���l>��a��wAw�I�qM��v;�co! ����8�2��U�	������ӹ��1�p��f��O���]����J.V����Ƕ*�g�X�SG��h�ir7�7H�d
u�&	�s&�^���N�p�X�%߾ ϯ&^%8��Va���U����*
��"<X&*̲+�ϒ��K� �~�7ۜF��\�٩���z��٧	��(�QQ�<���@��g���Ќ{/�5鲦�~�y0o�T��e�7��?���X���m�� ��#�l�Sz{�,��t�Ν��0k��󨯊t2Ti��)���e�#�S��۰�����c�)�gev-�]�l�`F@at�i���ҍ]�TV����)�PQ��8֫�2k��Lcp3b���u��e�L/{r,5��5����puP�,+/��y� �ݰ�U�����GWi՝�E	U�ƺ�\��]���XY�R=g�t��Ab��y�:��%e�+��t�s"p��q���|�L/Ne�2�jx�i��I�9�h<5�_��11�{J%��ۻ����~����s6>�$e|7SƎ���v���÷�-���o�w��ye{����S~}S:WKK���.޸4=�-���dW�ײ2�31�.��|�ִE�;Y���>탷��MW��b�� �zC��t���=1j�kK�e$��LaUB,Q��!u�7��v	�;�D��.L���c�[z�+4K�["ȋ�c�N��v�7�c�ǃ��+X���3rM���������OY�w�������;:�;��a_�鈝5;1R^5�D84V}1�~��zU�0M>�{����tQzjd7��_hsng8�^_O��h�~�̺<�͍���K�ǚ�Ҡu'[È��֦ҝDg
���{��ap�ӹ������f��脦zH�:Xp���%�]P�)��Y�oP\�-��źt�ƥA�$ȥ]S�4A�D�#=�P��.���r\�^ɝ����@�7~�/�on�Qs�x������?�v��G".�p�U�;���,�5"�o,a�qq�G�ۃ��%a��������fJ���^�N��/Z��j6�x�}�W�����fE��M�@�ra@�?`�8����(t�!r�5#[��}� 9��Z�=J�F?��I4R�8$��3!ve�W.6H�@RC���I�Y���i�J��8M]���v��[��H��萺�{v�`�0��3�
Ⲽƿc�������m��2�z�tDu����bÑ�t�:���#��lڮ�{��:9[�)���V�;���1秭Xޗ�ҭͮ�"���-��sn���N]sA��X� s^)vY��r�C=����6��vd�"�k'E�)3��eC�IN7��KJ->��{�-[\o���J8�SW��Lo����a�=\�*���R��L�rĖ�}��}�y��ܞLT���Ө���v�D	f#)l.�pЅ��Qa��rp���u�4��X�����iN�7�ϖ�\�v⺣��T�`w;d�㙡�����}bm�@�"���qbG��/V����,V#��vzU��U+94�/��<�A�)�P/�vXF�������R��.Y��|�ݢ���쩸;`U(�!��_V�ĩ�+���TW^V���@�Lj��ڳ�Z������ܳ���!^ө.�}h�Q�Τnϕn
��6�|硵�;��"��-Y��Z���4%*�P"�H�S
�� k�������ڽ8�� �B��lLnlm}�M�Ⱥ
,c�u���=�(�%4	�E�G�6b7rg��jcH� ��en}�5g��@�]�����|kb�l'2&X̮SFR�s�z� �|h�ת�GWi�+�ٗ��{s����٠��:-98R�M�Cz��b��ng��o]�=Yϑ�ƴ[T�|��S�^!��5p���M>\����6 B�ذ�W(���9sA�u 2uak�2��6̛͓hn;�.��YA�د��,}��]�72$�'�G��ʅ6�V��-&GԔ[ҳ��9w�n�#�s�-+j��������^h��W�ջ�3X�ioi6�\%�w�����qV�r���.�}� *5�%Y^gI#��k��M/�k��|�3/�X1r�7֫�$��קb[�ⷥ�6*����t_nTL\C����f�̽:p�t?-l}����t��adZP�����Ⳍ������8��!��D>E!��@*�p�2YPo���u�i�[�J>�}�)�Y]�skנ)�f,9"Z�
���c�;���1�@#��k?mf�+���F�G��c�\�lޕ�lv���4��%7'�7��*�ljɫ�x�{id�xY#"��4[V�.U�+\^͞B��p������v�Ǵj�W�4�
���f:gg��y�B����Ȝ�:F���k�*�w��}iW����Όd������C�.7��]�1�^�٪�#.O=� ;��F��iWx֣��W��U����LD��/��{e����>�?ez�w��K�>�eW�`�X����'�y��a���]�B�L>[\����Lb*�r6:�_�4�xo�Ge:q�j��Dq̺\.��>��Q�	�;}�EAs3�3SI6W0����˄vmj�N)>B��ݭ�:'�;{b�SǓA�i�)�2X�;s���ϳk/�_5;���j�Y}��>�p�����w[�A}]n�d5(5��Xe�{`N�څ�Nm��K���7	[��T�eD,���[@Mg����A�� T�l��d(�8P$ӷ�y}ܭ��w�O�z�̢�x+�Q�=>mTuh�⡢8*:��5��Dg0����٩��.�!謧�rԠd1JTh�)*0����?$zM���D8�.:�W�^��u�I�'�F.y=�8rn�,t�F�0����#���]"EFÄ�R:�y��ޥB��o'�9!r]t(bZ��p������V�	�����5 ;����rT�FՏ4��?=�/��իgh�1R�(mK����y��G����ά�耾�"��̙[�G8�XVC9t������1�U�v�G`\wt�
�\�l���h�Ϊ����"�.�P�.���J��R/���U��A�꥿��~)�V�aI����2y������0,�`�f�v��V{5fP�@l-�L���j��0(b�he�NÊ���Uܩ:Ǚ:N/I9�sd��yhso'��'^F#Z-�u�a�Pv�^J�Ρ#��]�I�ꎱQ���w��;�ukY�;X�'R��ܨ}�J?)�I9��S:��Z4���=�sJlL]pT]�n2��${�&/9�d���G[�Ա�܂����<�2��\�nb����WK
V0i��+`�P��i�8�>C5�,P�OU�:����9������� ���v�o��Ƚ1���G#ˡ�^��5Y��pr��!]q㶬^�3ik������\j��Z{/���P6�u��e�~c>�M�Y<'�Y�ԩ֩�u6��oe�W���VFq�(G3b&H��9�e�7����:կL�ї#��g��Rh������|N%S~g:�Z\~LT8����x�6ܦR:-��
v�c1��2!b�=^��j�v�=h��@W:K�Mf��N�@�z���q��F�)�7����&{��(��_�T�?u��f�*�i���U1$��&�g�[�J��j���*�=�i��Z�&���#Q�Ȍ3�;Vq�k1!)�5΢]�t��Ew<,��-;���P޷C�ƉN�� �҃I��f����6�do�F��@�w��[w�%9�Ҭ���wr'�;�Ce�
��@��4�P�BѦѧ���7<6������uY��P�.h��ɍ����"���:�k�|�#� 5;d"}t���t�����|�/%�2=��h���D���wy�7}jf:�YlR���qقV����dl+*��{k���Ƿ��ѝ}�3��uR�Z���C�J89�}}��]�	 �ږ>��؊��K�  �L����=�#�$D"ʮ�s�
sȎf��ʪ�_�]��jd�<ޞV�����N`v�R�+�li��궥�
�ܼ�a�F�c�7]��Վu�"�/��W���[�k;4D��6M��'drSG3�#u0C� �̤wNJX���t�^���@U�Ȍ�Oމ;��}wn�\�� ��t>�LX�u���#�JK��X묊(�X���5�Gt+�v�=�	߽SUXuV{N,���s���n+�Ѳ���˜���L�9u���d�~�Q��v.�(u��/H΢�`�uZ�}����ۥQ����Y��6��R�"6��p��Q;=>��ʦv_
י�S��r�a����:���>|�.���X]�x���hK���Wxp��W�����ct�Å�>��>`�λ�t��o�.;�=�2�On|~�]о�:��%5�@��k/��%]�KqS������꧐������f���"�r�nV_B��$"6�©�^�P�^k�����̫zr���$^���kN����(�k�6�8I�ˇ ���dWVB�o�O3(�j����ӴܾZ%��'*"1���_ {G]�$���_�Gby����f,Ű.<��:|o�X�-Ч�o�v�@R��c5�K��KR������7K����\���ӫ��(�{A�E���%�j{��ex�z��`�����<�v<�:x��k�T�q�?���R����.���{���@Vq���?\����5t���3c^�U���MYHg�<Y���)��2��v2S5e%"nv�6��:+Z��w&���54��kT�9j4=��2��5��[���ׄT|�n��9�/�{.u�l�7+3�gp�d�^�`�JsU[ގ��]i��&��]}�Y"WH��\n�/��=��ή�T��Y�?8���x΀T�ٱ�_T�x�U%�9)G]��a��V6�����zn̾�"�,W+\ �V�/��pژ���C�DE��N�D�ntH������'x�JNخ��{\�y��`�	��-�|�T��q����qڜ"~���0BtjV�w/܅E�	�G�ܐ���q���ٽ�Q�� �vs\���``.��;{��p̄[��Z>��jχPe�V�]�+r/f��9��*#�u�@�k{�qU��d�g-���v]X��Y��3we���Ě���K�Ji�Z�R�KcVM�E��J)����9�u���k�'�hBcv��2�U�WD֎�*�i�N3K2��!��u-��[��t#�t弎I[��F��%�U�mu�ߙ�F���:��,B�R&�{u����̜����7}�D����Ϋ��/P�X�wl�R�����;;B��,5g��}�ȩ��ֺ��D��Rt+�c�=5�j��l�/�2H�]�[�^�a���]�E�Gs�E`�й�CR�ʨ\�5Q�YX�[�9v%��Q��46�٧���R�_b\5��J�F��%�&�.�e�U������ᮘ����ّ���a�uؽ���ׄP��Pǈ`J��Sw�{@P�(
YȚ:=�DMSks���D�'@�ܺ�K8+qj$��������p|�nt�Cn��Sx�:�ܬ�Su���j�d�i*iX���в6<�9�	���ł���Rh���II��o}ܔ�D7˾O����MQ��w���#��8d�]ːW��^��[T3(�1c�ա��(��62�u� �L����⾽W���U�2��s��q�}!U�2�Ll(t�2Z�L�v�6����WfƲ��E�.�o2�mXm�'��
/�F�x���NJ�7�f���5S|K������b�e����*feZ#���*�t�B�o����JZ{5��H�˧�,�`U�&����|j�5��2ƴ�xSȚi�m"ˤ�20 ���2!*Jm�>&	�h=�r�N�W
w��%�f��L3].���=�Z�^䙬wZB�Rm��t$���N����yX�� )�0 f�p����)�t�5��Q�ci��E�N��R$5�,��U��b���1]S�uY��1s�{v2��I�ڸY7W�[WH��]��VJ�Q�NbZ���RZ�� �gj:9�`�Y2�
c.�3Oh����;���v�h$-�=}PL[b���u7{1}�,���*���= �d�A�"i�b�(;��1RO;�@6��ڃe�nc�+�n�*�v�6���w�#�z��/�'5�]H�r̻'oo�I<���������K��;��-��M�Z��N3Iu�	� �5|�h���(!�.����Jz%�X����ĭ5�^����
��v.*�kW��D�@cx�t�x�:�-���#���E��V���W(�e,G�P����U�|Cr�撳 V`��֍�Lw<a�0�;�2��n����u!�,�x5V9}c�b�b������1�΋h��|��\�Ǆ�d����|j�ݓ:��lo�v�(N�:��pH�Vd��/u��]Pf����B�\m��زT�UZ�ƌnf5���\[��,�V*���b-E����Y�73
�r��0*�1��2X�V���V"*�,�V��T\�*��DKlb��0(�E�**�b�llQ��R13.1H�U.S#Rڲ�r�jUALq�R�9J���2��ˉET�Z1K�-��"[AV	s&��l��V��Y��*3-���fR���lmUT\J0EV*�(�f5\�b�F(�e���2ŨR�ʫmIW)(ō˄˂�ATPehF"��J��eE#����IYkJ�R�T`�̂��s0�UJ�#��n&E�+�b0Ƶ��¢%�J%QKjT*6�Xc1j�m���V���V,\s*�[ki�`�H���V��Uj\��Z��*���UıĨ�S�+Z�Q�Zܦ+��-lq�E"�hƉij�VD�Ԩ����[�� 	������m��e�X�07|���"nm����s�z��C���?q9\�p���T�^K�]2-n�PЅnި�K�������sos��X�I6@jo�*�T�+~�� /�{qW	
���ү|���$��|�{f0w=s-��mBmR�V���Tjw]ß\�/2%"`T�25�u�y�j�z��x�b��Ь|}X����s5g�<z��mV�}l�����w��q}N��G�����L=���z���=u҉��΍�w��J��>�-���K����`���'9�
��(���8�1<W�,��^��>S�T��Ӳ�!�_��a�E�g>���t��P݉���
���w��v	��cOO�� f�h#�`C*#���qؚ��<H��2���Ok&�Y�'�WQ����ddW��L�9*0���������<�a�C��|6���.k��9e�,�����0�Փ����t�9d	�+�$u�+�G:�f�~B�t��.p�1�n��T7�gAP�N�����_BY.
ϛ��c.��Ad	�=s1N�[��`�[g������C*4?�]:6��v�Hp'��iŧ�l�-�@��H����<������G_�Y��
�#3��X��t��mp���Z��4ЇF�``Zr&��wH�]��2��n���n��P��awN�/��q�q_3�R���$gR76;�$�}�J���s%A]0�-�˷�����@^&���xPð������� ����]_���}j6�5�)�&'<g�@^Q�nvN�z]�ȟ���I���LCfé��3�+;�7�/N΅��_d#ܵ`>b��ͩo�q_�uV�aI��Y���� ���*}EO[3{��眬\�y�C�r��:GY�+��6�z|j���V��qu���IM)7n��r�R����071�aBo[Vkj���$V�uJ�pT>��
�]׺v�� {��9H���n[�� ��S��h����dι�Ш6�L+/����/r�5ܲ�\�j�ilIG�^��o��|�o nZ��
��G�h?m<GM��g�x�=�D�3�_�02י���O�5|]T>��g�#W��2��@�/�F��rt�����ͅ/ۛ��iPe��~�����a(��F�C6��+�Xi�l�i��B.���J���5���H�z�LD�,@W�%�3�EŃE8������9W�3N8��eM�v�U۹���Ў���_�� �y]K�@�H�&�a/���I�N�zk��i۵p���N�]�(�t��R$5�fQ�Өi��%ܷz+fe���Ǿ�r���Y|���q��t�VH+$��X �e�x�>�-�b�D�:�<�5eo,��r�m�]Vz�dyqu.����m�����| [Z⫓���+gbc˛y�Y�9�Ȉ���vtu8��F"�%�S�)1�V�>�q�jէC�����P}BՎ�%:�8��$=&.5�Fb�N��B!�6:w��:�(�ҥ�ouk�;�Q��߉h��O�$r�6%Pl��y}h�"�3
zė���9�Q�1�jV�_�;��С����Ƃ�3�p��&k��>���sh�4�'�KU��ٳ�R�]�TG<[q�h��7>Q�<��kl�|o���S$.�u�
B�m�UM򴧺znCv~\l�X!�1�\�D���TX�	�ሿ�,̲���W��@�nM�����	�A�U���4���pi'��� a��HWf?`�2��F~#O`�׵PZ�vD�H��*���>ޗ��a�h'B�j�?f�<n��㽤���f��cT�߰{7�mt>��|�$>�}Y�@n_�N�\0�u4�����b�n���..r�u�ȂC�Zb�h����Ѵ�Q��S:����������UV�[��G)�9���W�;^M�&���r���eJ�A?z���a���&/����c��#�㻱�5�mY��,������չ��M��uw7{�苷�Ga7����E�٥���1a*�)?UUW�Wގ��޿o��c���k�D]���먝���yVq��}K޾���� ��{��mPJ�ѓ�_��J~��G����P�7^_E^!7�>�K���u�u�s"���VtTo��M��n��|FZ{sP�F��tО�����K{QW��n��'Ϝ���S�ߘ��|���MLիkjPr�&F�[�rKwY1��'q�.�Wg�����-�{��z#��t{y�'#&�SGC�ƍ����E.o/�]=iG>�b�d���h���4�l#N&������N�r���{C�֌N�q���6%����۸�9���ޛ��x/��t\���Sٲ�����&��e�9#�E��>Z^��˶
�k!ڇõsAD����<�X�k;�w-�>|�F���ºub�X�<�U�'N���{)�!;9��@�-��0f��<α�B7>��@b|�[��)&��G����t�6��j������FI�ǂB�ڂ�(E�k� �/��nJ��^�
�gt�T�:SI��I�{������R��Gf���M�j �u�qax7;
���bLȘ���悪���:Jl|�0����}���a�r��0����m��VH�?v���A�.bWD�ڼZNS�(�]T�{��~ehW�N��W�
��_f����|���	�)�Q��'lX�f�O;z��H���Ց՟^��:������l'9��b����"o���}�z����ngF��7O:��9X�:�q��R�g	��k'���s�R%+��~0s6�m��[۞��$S�m�V�}�歾��������m�޳Йǝw�g��&�s*�mo�<���ޑy�͟ugd���~œn��[��y!�쿓��c�N����2\0U�%.�9��}C�1t6����I�N%�ä������~��q��س��z�Ѫ���Bsv�Ϊ>}J�kR�ǣ�w�a_=�'��;�q�H$0gp�;�,��_l�=:#���3�
c�*���3�0UPE��o���N�Vq&�vIG+b�0��5����川2�_��C�Su�⃸��v�+�c۝cpD�ٙ�;A�hi��t��&�:��;���"@7t��f-[��mF�;���ͯ�}���޸5y��޼�v����9A�N��ˠ��;�v�C}��H���'k�UNUֻۤ֨��\��y��������}�X��B��u ��\��`9{���+p�e�9��B���u��A�3��Ϝi�/�9z�*L����X�o+9�\+��y�ML���6:�x4���G��k ���������~>��K�X�j��Urf�A��;5�2�M�'I7���/>���ןi3~�̌YF'?gu����M�:%I��Ȝ�of����=/+��F�NtRͷ��f$^ȉ�SFw�mbJP|���r�1IԞ��Q�uY�uoxoxk�N:�SN��&:{����uKn�R�d3����s���H�Q�7�c%�������]ڇ+\�V��C��į~�k�M�xͥ��y�p���wS��Y>.�$��\��7�u��R�N���j��B/H�Ǝ	b4M>��:���;']�-]ԑu-b�t��UF����Jj+v���r{���(pѽ�����ݾ��m�jډ"�Ά����}_W���_��a��y���n9�����sjM�[��'��\h<�f�T�Ԧ�sU�|��X}#���~���;4)�q�?!ܙ���2�j���&��Fh�\me���`=?�@.��iS������5�k9TK�ܞ{�s�|\�o�����l�@�S��Б��5���(��v-*�~i�Pk�������X��y�t����;����)�]FZ�ILqB]_v�x����h���\�N�(�r�uP"����R��ժAb��b7��л+�˸��kw�:�ĔU=��;-W'K-!�h�]xC3�g���	�^��ͧ���B�0L/"%k�ܼ�7e��,N6!^i�ڷNپO6��ɀ����\�W�f�����h6͉��P��_[W��T|ďs��+�S�)(�4ͦ���E��v��s<۷v%/]�b�5�~#e�Eg�H�ռp�Q�c�}�v��GvZ�i�'�wH��a�+h���A��Z����f�����@b�n�qs}7H!g]�{� ��o]�ZL�i��H�v]��9o��Z�1�@���[��ب�P=w�]�����[-���mIB�{)�j�Z�kg���Q�GTޱ�����u��Vj��ڕ����Q�Qg� ]��U��}�7y����;rV��To���-��mT}Y��j����{p�Z��RE������:�.��-���7�W�����k��v���:��88���.������v�6�Ͷ<����'��5���g]�W��>̊�^̋i���ϩ��U�U�6�+4О��TG��N�D����s�JV�Ҟ^>ݰ�����6;%m�U^��#DR4_b�U�[��Bk_P��|�M�Ҷe<��=����^�I�����0#�~ʷ]w�ڽ��7����K����������U�M�5y���Ⱥ�]��S:n���8�X�2��zX�tnM;� �����4(s�1��`��3�Y׫����w���"0���V�R��l�����gGڹ�4=Gi[NS-��u�"�ñ9�b;���؛���^}��,�<i�Z��:T�)V��	H�~��Q���<��6��g\���qM�V;=�����{����	HweY����z
�k�ۻ�7�hأ�o��o��/��;�N�h	��D�]��["�%3��_k71um��C�z^.ݸ�7Y{��pƃ�sb~G6v3��hV[B�c��T^�:�ک���XdZ�5���v��6��K�l��MVc��q[�M�n]�5	��Ih��i^�\�gԗ{\'�@��OK|9����giK�f�]��{��6�__����/E������T�t�z�x�d�U7h͹��Ѿg����)�ؗQ�ӄn�����'%z����(���4��q�?d9G�}�:X�+ۏӪ�䨯|�^�r����x�_���W�b����=w�}���'7�ǝ�d�,C���U����F�F.)�o^#P}�֔��=�6�G_f]kł�Z�Q}/h�27W�~�O�Y/���[��xQm,�����*�Ǒ��Z���odɟv�k%�O5�8<
 ��%C$i���+#
�|�,����� �)T�cj7��]��go�����I�����OHv��9q���6���pĽ�΂���χP�]�n2�����k�.����L	�ł���z]�Jd�Q�L��U|%	�S����j��:_�Z�&�2�C��2�o(��]�cw
GWmuf�[�=�o,����)�����cs�ޱ�O"�'IX��U�)��.�Ϯ�GXW�gjjG*��R�[zu���ͮ������������<g��{j#���n�o���վ��w���]�[�w�֞O0ȥ09�C!�ϐ��j�f�ʷ��]{r�'�g�̺\ռ�PSÒ���d��38KY�Җ�A�y(��{([���C/o����h��89��{n�oSX�������3�`����w֙�p{/�m�ޛ�HT7y;�܏8�u�R
�_G�cx=n����<�۴�\���l$7~��e����a;-Wx�[���W@�9W
�"M��t�X�h��W���-(��.��_3�6�^��4���
�=d���Y�����2�\|�^.�;�ov$�,|�n�h�U��3��iܽD�B��A�D���)dϕ��r�{��i�+�w1t.a��KiLc�#l�s{}+�)�]s33�v���w�����u���g]5�mK�d�IyOd���q��V�$��j�^h�w*��VX�F��D;�f���S��9�rp��S�%���x�'8������꽿���ӗ]�][-�*���ki0�<�nV/\��=O+3Cgq�h�Cnw\�:Ѵ�^<�̫�>}1Q���]q�}af��1wFNi����:�+���ܧ�V�v�(R�꽮�W(t�=�����ħ]���9(T�ӺqP�6w��5�(;鬽��
}i1t��S�>�u�[����)zk� �w."N�>	���MY�IDl�K4ҰUh�o�WK��%�Ƒ��<|{y��ss9�����:С�V[$��캾�v�ң��n+�()��p�7j�!NS��̥�
�,�ݛ�V�Kӊ�h���f��Mf�;�7N��	��6"in����z�k6_LM�aa4�ާ�v.
���Sc4]�=n��^� �����A,C�뺇+_M�f RX��M��y4s]	
�|H���;`��@7ժI'%J�T;`�j��w![�̼0��_S�
�l9�U�=|�k��[ǜ��:h]�PQ����R>�,���]��z�be9���Z��sS���;2(�\xX.���)p4O�E���k�1H;]�.]��%t�E�v_`T�c�:�h�Cm��0��W*��U�C���n��܀ݺݾ}��d ފ��yZL�V��Ko4,Q�cZ7�Pt���T�)�n)7
�y���W� �����h��90]�=���
d�S��m�C�.�O{Ocذ(��g�$�C&��.�v�j%�w`N�û�SC��u���j7Z��V��Y;W�1j�1�<�ա)� |e�ڨ��=�ĳ�"�y�NL�q�w�[��h7�l};%�X�Z�8�i	���PM���](�ÚuWgj���*�궧e��^��]�9�dWB��Z��W�*��{�ts|��%�9������"6r��A~mS�ok:�Vdi9� �#)��ǟ���ꍉܯOM�+�Q��i(�ꦖ�k��h��.��V���Yԧ7:�{����� ��5�R�ە�z�O��1yK�:�5\A�r�0H)�(�w%d���ְ�hu�c�5��������w���MΓ
˛ �tS���vs+�rVȸ��C� �\��Zrw*)���[��a����7������\W<�'���a��[3g}�γ��V�[e�-Z6����Q�e0�ʣEZ��̙cJ[E�eLJ�PP�TX�3��%������*c����U�a�R���+R�VұlG)����%�-��f8*孵2ى\���1��X�Ԩ5�&ckl����Q��jT�j�kJ�b����ib12�+[Pe6�J1iaj5Q`�-�T�e��pJ��iQ��FV�̫����r��(�*c\f	��)De�c���EE��.5m��-��KF��+�Sl���`��r�m,��L�e�ҍTEUE�*[kJT���S.aZ�mJ�m��0ɖ�U�2���m)�Ĭ)naQqml̪%�����մ�`�j��R�
գ*ҖZ1�*Rؖ�n8����Ĭm��m�X�Z�J��[Lɂ1�km�-E,[F��l2�U\s*�Pmh���f\c�V���*R��ʍ��iE���1�#���iZF�����[���2�2ʈcQ��ѭLj��UknP��1�ƣJ1D�k���H�j*���T(Q$ZWm�]yk�B�����蓏�zy�F��J�Dd�2��7�\2�]:q}�F����M�<�ザT8�r������:�������'k�䁇���<��!�
{JYZ|����oͺ��	Wgu�q��p#]&���c�I�9a��U�WݏTb�2'*��� ��)^V�Z�(�5�ʈ�N1[��O�\��h���Z�e�#}���[���=ߗ�v��M�\%4k�����B�f+C��.n�]o6�\vQwS˕?Q�_Z�M^rU�ķ/k���|�ж��	�\���K˙��CR:�.�O=�rr,xv��Իǵ,B���<6�[$�bw��53���EWz�P"w��[ݘ�L����ٝ\��v�iO/��M�*S�dvP:g�����e<�X�Y���lu����1u'���i��`cݠ�C��T�Z/��t8���U�<�>!cO�x�5��t�Ҋ}��}����r��S��57�M	qX9
��)��ق�>!*f�MH�C,�IY"�.�5����"pa*���1�=����A�u�S<��H �Ȋ���ָ�6�⭍�;(��[ �M��2�ɛ����MX�֟Wv�ڷi\&u��݄.zC�ri�_:���W�Rcr��7L-���D��dG'v!vW٩��z2���By���k�n0'�6reM��mP�4���C3�g��O2�+����R�Ω������巏���l)���yI�F��F�یv��y0J��ROf�km^��e˱��>�u�Ұ�=�eKj�:GoF���J��oV!2�j/���������.���F�ې#Gt�ҷ:_;���䱛{x�F��#-N��a��B�Ll�J�����^���<����w�a1�=Aq=���0ԧQoӔvzZ^�N����3O:i����Ĳ���Ss�{��.:qM>�������yFu,�, �Z�W�ۦ|��rH߫L���-�h����o�W�_����^Xޛ,�N!��;���T�W�sky��%���6މJy�Oy%N�����"_�����nY������Dt:$�'FS�3뜡Kh�B����e��u���I�,mK�KW�C>;Ì�
��lG��p�X�^���8k3#�Í�v�M�����M`�ma����ʤ�7ܧt�ۋ��qtw�o^
�;]�op�ܑ�$��� �TҬ\��g��i^5\i�S{@X��f�; ��r)o5�.���V�/{�t�k۳S����c���l�{�GƠW�����3��;�j�\P�����/���}�z���[��9L�3ܫ:U�*]���)���ԁ:A$F�E|����K�G'�X���Z���"e���1c���T�9V %0��C���bfFɼՓ���̝71?<S�ć�6��/��k��"3�vmN��yV����mSIe�-;r�Z�%<�;/��;诂v:�¬{)N�hs�s=d�u�p[�}������ov��Err�CA턫`�gbt�.=��wn�:��ͼr�ӷ,^�ޘ�M�}jeԛɨޖ���TI����o.0�ú �Ȕ��h�x�ZsNǦ_�kY���0S����I7����ɉ0��z���2-9ݾ��ĸ!��vP�K�[��h�Ĵ�$���G���}�	���قF�m�{��g\�tx�����ɷ'u��G� sQr�6�:���|��|��D7|���ޫ;���X�,rO9D����g��X=r�U����r�ɷ�޺7�Xņ������⼖q��[��?���N ��kGE�no��>�.�m_�橱���[�U�S��'�	�{��%�������N����r�}�#����RK��C8b��NVn�1,����v���gH5��oTc�|�����KS�|���|f�H]�\ϖM%N�k����x�u��h�vj.��U�#����WD������aW��8y[�u�*V\�������$Z��G̗���	O�����:���^
&�3�)���U�Ӥ�6�ݿ�Ka�}	 �ƍ�H����˝��R5Y�9���^$l9i[�;g)�9�[*�A+�;u�q���"�]T㸾�m
�V�rW`f�n�<�X�B���O����OX���^��wK��\�^�{���~��r�8����.�h�Q_<#�06����k�r�G�sk�7=i��eA��
�n�x/�Td�"���1��Aa����ܺ�܊�8��hƹ�já+�2�T3��`C��hj�ʻ��ZC��ڃ+��6��J�����6ާ=��e_��ف=��i\�}�+l'S�}���`�W\��$���oc��}y�@���2�1z�a\���O�����)�V�L����IΟ�U�޹z�ȳ}s|�V�U�u��M�tkh:��iWw`.�	głDl�Y]�l�W}V��Y��N[!�����5=�6oVǯy��)Ües�{�#Z�%X�W(���g�X���(�y�^�!]M�jxc��y%�>��_C1���$�|�g*�[=�g}JOmQX��/o�ug���r��tY��c~��Tm�K���6N$_�珼���3���{��}�y�K��;]����?%���f��U&5�n��5����u�6�Q�1����:�Y�K������ݮ��)O��q��+�hrź��X4�u�U�"�w��&ڜ��*v�n��Y��]jZ����`���m�P������o,���(u�P_c�q�
�dU�,����\#�H&����ὸ8�|���t�[#��pT��]�!�����"%��_E��S0�gA�v	K��|;o������W� b���ouUׇY`re���I��5���C�2�~���P{���x��r�|���)����N��_&���ZM�~�2�?s�#��S/=����gu��a�������ұ�-ָ�-1ǣ�!9M!.j������Ņ�(B[A�wc9*�q>��c!Ʒ¦�А�$�yZ�ŶU@� wN��rv]��.�Ek|���2����+-��Wʮ3�f��Y�r�W.�!�;��yb̸VH�j?RV6�=�f����G�$�߽'��N�[޹w��rt}c�#ϊ��p���5��6�\�Sh=���t�#��+��r��q����L��������9;��㏓c�>�0�#h;ۢD�沍�9�a\^n���Q�q��֭�9nw���5%
�=���Ҩڅ�4�[͚�"�b� ;E-�z�� �E�o�˿_�~���6�܎�:9��S�w�W��XA>��9��TQoi�G��f�@�fҾ3Wӥ���a�k�Č�0��G�0��t�djj�Cwp���7���z�j]�}_}�����7�5��ۢ�(�kj��YOAr�C��}K��|fy�#�����Z���o��]X�q]���[��-��9����#]�e��d���i�)h��|�7�`�
Ci^y���Ë��� �׻�SF6�f�aT�>O�zzr?x��+�G�-�3�1���{���y�i-�ĩ�w���K,6�l��x�k��ߍY���ʳ9U�=o_������k�:���{Ҟ�Y�'�4�z�<�T;]����Ջm�1j�8cK{����ۭ=w�-'���Rͭj��;L�N<��P�t�뺝B ���識��V���l^��Q���cS����^[����q��;r���Iq�j�v��Օ6�u`�j�Ib9��_��t��N-pyd+G���k����de�p�t��r雾���z&�v:�Uk?l�h$C�|�q���hQ\-K�������ܽkM�qp�<�v-��N�}�Xg+Z���bK{E�Vq.=�k؛[]˒-m.=@�VCg9�G/��2	G8�ݝ�ww����3�V�7J�wC�|���B�<;�������D�sww���{+m����-����v�Q�err�l)��	�b�����f-x�q��W�W�R�6�Ϋ�]�k�9o�M�;Xr�ق�4��r�b͘��ۣ۔�t/1P�r1dOz�:ꈠ��
U��5M4�o�����]t�,�����~��Z���&�kM���D{X�{˺S��aS�A��)�O+7Z�r�]�r�S�?L��F���dk�3�u���)�ud^��qj����>0o5s,��q���-��S���7��1]���1��9Cq(���7�띵��#.j�����VG1km�?g��i�]L�0�)�ϟz5�G�!9�E�M{Ԍ�7�{:N~��tu�$'ToTbC'��W��p���k@l�e� ,�)x@n��Ӫ�7گK��2� U��뉆9J]�(E
�E�xj`�+U׍�h�4ʝ;r��&�N�pq�̋��؊�=��޳ۀ�_9@lتr�ε�Wpَ�I\���0V�x��m�깎ۛq��(�k#�'��R���%X�ib�to�Qڵy���A��b�5�|j[;�L��m�;��	��]�|r	h��Cw���1��U�wIғs|]�W�i�;ɥz�m<���+��U�	�O}�l�/XקN�e��}~�i���ư��9�3{	����	��ڈQ�р��I���T��t��=��B�����Z�þ���-��yɅ�R�ά�1��Ϸ��r�)��(by��+�e���ӎ��ﲷ��;a���ά��M�\q�Pv�[��O,x�9�ͺ���V�%x���k�yK�������A����-3Q]]:<Lj�w7X�7��֭R�q�Z������B��#9�c���K]��_jcM1z�(22ؑ�m��J�1iԛ�rÔ5F��]��>�GV�0���;����;�M6���<����h�X�l���칷Q�Ss3�`�;*�����k��^�3��'9Ӱ�N��av��I�X�]�ܼtP�s�Y�i	^W^s�E]i<��UeZx��d� ��y�V9�u+���ӆ֭�n������T/1j����VH�Q����u�X�A������j��\�bt��%�q�@n�/sp���)y�Mw^�M����W�l]Z80X|���I���Q�Cqo�����(�3<�uf�J'3{%��[�';n�'c��G�?W����MI}-���_��o&z�]���5-7�=��B�q��m��o#�n�4V�sYB����}�����LN�w}���u�Pg��I���V�PV>}�e�Ά5�Mj���>7����]"��m$1��oc��R�A��K�Ub�k�b��,g1$�խs���\�6Ԭ���Li��q�*�m�j��=)�b���swbf'�����dh��)�1v�]W�F^�n�<�!\��4�;��<	���r�5�������D���r�)sxtJ�f�fǋ�� �S,�*��i*�QUY��7��!ԯ[���)�l�ұSIg�G���ǰX�t6��MV�R���5�J����a.���;�ŔT�9�h���vp=4b���IW6�\�%Ki,v��v��]<���.�ي�8��
zK��D��,j��k3i��{O$Z�j�M���5|"�igZ����<K;�c᪆��1+Zz�Ҽ��������;M�P}m]:�b�84� nM���ڳNs��}��&��r��m�Zybې�S�xr�:�儶>�̘����li\|��?Ii�Z\K�
f�u �=�4]o�A��VR��wf�����*��*�C6R��X6�jr�����O %���|���C{�n�0��J�Vso+v&�� �Z��ac���ܦ3�&d�-��
�wټ�c�.'�;�u}R�t���pz�u"Z��Ա�Y7��&3;%���V֚���X�u^:�Rͷ*�؈��}-��]ש�;�oe�k���-�#�Ыt5��GV#�)�M1��W���Y��dH^v����1J��"�k$��dX�|��##���C��uE��'���*�:@���W]��36#�p1.�6�M�3`U�����Ύ�9�[��l^�g��t��5N���F}�U�~\<h]��Q����R�ϖ��\>��%�Q"�.Ɛx�#3N�UϢ����u`����C%�?�y������������X��rYdB�^(��o� ����#{
­<�9y�u�*�Rd8{6P1��o1vkB��cY�if��U�+�K+�+��\��������Y	���LE��h)�)ۘ,JU���V�J�mt,���h����zog|����I�,�yf�yFVc��*����
l;\t�tV��/6R<(�&m�vA�`��j��+�O����>�a�-��p�S6r�(g���Nb�ܺ�8:2/��.��B�%sv��=X����!:�^�c�k-�Dr�W1Hv<u�l�L�Vkw+cy��t��;�0�z�:�Do�|q�}���V�u�<�u��&;x��ˋ̤�GJ+'}!"�u�tܻe��9�<`6�`�w<�c#�٠��q���u𮆥�7|1t3�t�*�Y�ŷ; �I4�6�v�b+�{�i�NR��X�P��uE�t�V�K�j��4���7���۰uwYI�[Z#�7"����.���e�aӈm�wٻ����pVR|r1M�7�`�ή<�������nh� ���3�^,�ʍ�d@�m�u°Ꮉ(z.F��e,��A4�s���yw�[�����Y�
Φ��'O%��N�\|�pӱ[���h�*K��d��E���vee��S���0u���v�v��˙P�U��QU`�Y�b�����beiU�����-jփZ+-3*G1�c��UZՔ�*[U-+Pˆ"�2��!ZQ�1��TeK[i�1���[���V�(�30c[m�Z��r�`�[bYQV6�W-TL��r���((�Acs1��1���+����帅b���J**$D[J��Y�cZ*�U�ʍ���L����������Aĳ)T�F�5�K�U����X�+����Ķ�����*��X�ĬJ�Q\�U�����W"cTs.GEX��jŬ*Ⱙ�ibĴmTDm��TX�%m�*�lj��,����Ƣ3(#\j��Dƫ��(�RZ%�q�+-�QTkX���*"2�����H�G*�1����RdAcE*�&R��`�V.+-��VE-J�QUm�PQg���{|�=����כ����ur4��bw���I�U���w�Ю�)]�`�Y�`}���Y�1ҩhĢ"i-�K� |�ryZr�?e���y�W3A�N򓎊+r���-�:(C�s���Ȯ����ąigc�s�E�s�6��Sa�f��g�Cܵ��~��8zK������uI�6��Zd�q>�).��5�h�_t�]�������W����9��^=�+bhcޖ��c;�:i5�an���jY|��,�(�_db��Y���MJϢ>���e�<2��Ft�X���7k)tSy%�����q!M�)������##Q�ݔ��##{B`s���o���,m.A�6��7�O*8�2rI�yܫ�7�W��͡��n�S�{˹����y-��[�&���8Faϳ�it�my��y��n��߈~�Y7E�%���b���z�Ӫ*���V���/��$�{�:�#�+rmQ���)����	�+��6FV	}׷33����uܨ�u�����sn��ޏ.{��@jn��K�y�h��Gb��cB����~��0��	��1n���D�Bi�=�h�
����JzF���)�)�X4�v��V���W���V2iDfY����hmo~��Q������⣶�&,c�<�	�u}}��O\"��uN���`�jo8L�[����)\S�h���w"�7����ټ�8B�k:�{��w�����Lv��z�'�U�)�����V��1�.�]�7�����[��nqůZy���~b8��_wf��"'Lr��0������aT0*���Y	������W�����r&����,�v���Z���;Q���u�D���y�w5ʱ�Ծ���Q�b��F�IK`��[��}+؈�߂y�/:E<3��s@j��=���^��D�]�t������L�1i����|v{j�\W��c>=��i�5:<g���:L��ti��~�ާ��/F����sP<�������9�elL1�[esF��|5�z�B�FH�q#���Q�_�G+b���<+=\a2�X��7�`���R��'y�/t��3��q�q� w��`�M�(ߖ:N�¸+�xv�7oA�^��.��Y�N���jt���C�<�`oM�T�T�V���l������[GKH������L���]s�n����Ӹ,�iVg .��Ӥ|�xK�';������}�����yԘ�o�^�Pã;X޴&�V;�s��K��F���u�{x{a���p�أ��]��k]׵�,噩�jq�V�S	�
���դm�72����������V=3�ܷ����f�U�m�b�nF�ys���˚��*��K#�b�6�!���I�,��Ҹ_^�l��*[y�-o�>����������ѯ�D�?Nn�v/`sG@}h[���n^��\c/�-5��������m�7:ə����C=Zr_��j���\��&���v�ȹN����U�Ic���N������ݞ�����뱚g�Mo�sz���HwF�&���jv�=֫+'\_s��Z��ve�y:M�~�pb���=�g��SFF����F;�4����sN��C̰!\��Z{�-تUQr-@���ً��[���Vd�p��I�nY��I+�:�v[ޚ;F�}@V�s(D��w`s��Wspr��� 0��ߠ��}�VL|�u����U�v7�/&�V�W�c:㺗���r:�J�M��y��yM���?Jq�@�ɝ��t�xg5��HnyPqbd��,T#�r��yM0���щ��;�
�[W]�fw�%D[7��w�n&J-'F%?wR��It�v��_#e�F�܌S�"ԧ5��O'�r�nMZ����m�7��lʮ�ѳ�O���uޥS}�ooI�I��z��t;F?iX�r����)�lZ���}]+:x�z�SZ��ϴ�g �m��~?����|�~�){~|��}�Չ��?'�<�"s��0���ӡ��ڎ�*�jyȹU�Z��~p*a�x�7˽���g���w�3O�M5%�����L�oX��t"ok3�;�����P=�ir>��w���x����A�~�伷�9pk�o��L��\���Қ?/To��>y��$�:���ۊ�k�䣍 ��]�z�3�ڥ
X�<tc�� 9W�K���� hb��j!�>�v�ܪx+)h�Npچ�0��������Fwwxoe��f��Z|����y�]λm.�KdaرO�������e�]���8�sjt�h_�+��[���|틗|�����"��|&�ا�e�]?W'�!4�1�(<gg�PS���EVŇ)o9{�fZ��������BI�i�wcOԻ���ά��o�L������f�K�R�r�D��"9��]�13��saw
�♾�9�7��N$�����������h�
�c"�{�b�����+�L��������#�i���Ya͎�򓎍+r�-ErE	�vr8��]�+�\��m=
����'T-�c�C�y�՘'�EV�V��Vo�5�@^c�Zde�8���<��G��{��y*���E��ũ3K�H�ۈwoN��}x��հwq���jOm��T����n�rk9D�㾦�r�ߙ����y�jS�'T�f�׸��gd�h�����|�X��*� �t+�������<M�0Kc�#a����we�	@ǥn���u���m�k��3�tq�.]./�u�7v,��@��ϋy˜��;a���_D����U(=ި�%�au:�E�Fdֶd;��9o���'�;��C)�q%˗��}�k����nm��b�V���]�m>,.!����o��Ooދ;���&�͒=�V6��)]�.êw^�.��W���o�jޓm��o/s˾���o
r$���r�g+�[�����J��/� odݖ78�8�{,-��ˬ�@��^�,_Ӯ~�u2�p��Ez7zzws�Y�1��?�V#�������	��/�~i� 3Y'��.C@�m��G�\o�)��m��
�ش��>䖄���M��U�/Y=ݹl'�M�޵���Jl��_t˄^�����R��rW1	��r�]Ƈ�k���u��byGʚ�iv����TK�ͼ|:��i����r��UM>蟓�Ԟ��)� ���ǹ�Y�Z���'����sϷ�3��]��E�Urt�A��q�f�"l�Z�RB����"ݙ�=�TK���#Nq�[B���P�%�uO:�I!]���~[�Sv���;v�j*�J��ػV`����&�s3{���UC��m�r��}����8�΄�M������#�E�]]�W�Z����׬�J��Vխ�Y�Xn��k�������}��V�b����׶%&z(��4�����2���oϒ�C3�ȧAYG�Yz��]W��\�4bB�@��\�-U�R�c�[Z��N���n�����zTD�{!;�c��Ҿ=qi�c�#���f���'�)1�Tb���A�Kk�F}��Z[C�:�_f�����D�R��/�U��Ǹ��!<�r,%�CU��$Gt�g0\�K^�ؙ{�j8����]�<�G���K���?�*\ᒷԯb���.�ȅQ���{S~!x��M%N�\����~��;��'�5{�v«�Ċ�_;��|�C�C^�Vd}*yg��Y/�s�0&�v
m���j�ᮾ���[��bQ���BU��>O���-�̴����v��[7�����ĕ7���pV�4n"�����;s����et��\!��ٮ��ti�z%có�7/-�Ȑ4��N�v]��Jk���7S]q� ��5��"�ɣ�\_��lu�C��hЬ�q�|�ȯ����;:oUmRJ�v�r���tPM]_l�-5ɥ`.au��r��L�)�2���"��{�{��dj��뿡s��"{t����yЭ�`8��f\LO�Y"D����ya�=_@s�+]�.̽)�˺D,oQ���7w�E�Z��ܼ�7���b32��F�lx)���_by�!]�.��;0{+[����W�����X���Sc���Rq�G.~3�n:]�v���_X�QG��T~������̷��
\�F9���v�5�n,��QS��q'gg_W{��3x۸>���XIt���@#f^�ml8��E��Aӵ;�L�e0{�̑V��'rП���]!lY	��*-OXZ���9��c=U޹^�A��	��=]���;����<�;�_Nq�o��AM�U��55�=�����u���GhY�W��T�=�-Z���(�K)U�U3c��x�:�<	̟a�{x�*����|Y�z�Q����c�/X۔�J�ꋪY�����M%�:sS��@e!�U��ش��`὾o�v#ŌC�(�.W�:�s8>n�)/l�{f|}چ�߇byQ���?%צ?%Lm{q�������|��ߏNio'��\��Ԍѵ(dtI����(�/u3�ϋ�*iǭ\������[�F��t*���u��
�Ro��j�?���,V����]:S�7m��ǭ��8ޮ�oi#e8�������tȍ�`���YcOԞ��V1��3���Րev9��wK�����Y�R/�|��<J�#��N�f ��ѹz�L�$;�mC^��)��T���wH홎n�B�s������/q��K8�Vq`�n�;���sHW�E�+��t�4=_����
�V�ve�r7��M]_<Là�>2�tP)e�W{���6�uP��}�O��2/�ۅr;������������P���"�jVv2���W2#���{����{α��})cT"Ǟ��f_��XE������-"[���s �o�,��:A���yh�e�\�t���;T���]���gK������V�;�tbu�F^,���$��'v��Vp�'��+ă������\��r�pZMt�մ�.=��������3�|5w��}�m���1�.��Kz�S̓{P���DkD�Ui=�y��c>G������}�OD\Ы�%k+�ݧ��|���rqG;�|}M`[�uv�XE��:jy˃�X�8m�K:md\𻒹�\HRB[�?ZFN�3z�k�P��^�G���-�O_6� �K~憿�Q<�������$�.�?�a�䢾X����u�^\a�4�N�Ә�w�ނmĔ��^?P���>��i�'���K/����M�%�r%遐6�H��Ӊ�����A��ܔ1��5e�j�)�3#"��ɛ�TE^�mk[ʩ<N6�g+�6�@�ᎄ�3�$V��}��TH�s��.�O�=���[��ܔ��JDh��܎�7OGxa�Wp�Ǝ�Ĥ9����-��b�)��5�.+���FJл�ͫz)gZ[2���d�Z�S.��v�Ik_S������L�f��2�m�-ܷ�^R��]zJP��
1X�]��+o�&T�J��+2��Y7jS�Y`���:���Q�T��ޡ*$N �Kb�b|�7y��'i�x�Z mG��r�K�]'EVÎ� ̾x�����J���+7hU-٠A�p�M7r�P�K��Ɠ��_.U��ٕҹk5� ����%:�L@.��z�K�����*vf�^:��5�'�僎w5�.�C��J�)�끮z޸��഼��V֌�ó�v�xm�N��ծ�� R��b��r�Wۤ_���q!�k���#K�U�[/"�=��75�"��x5,詼S^�Ŏ�f�j]�����܍�J�³��Q��Ƅoh�Wr�w�ԑ=3���ZR��l)��ӂ���8�sAړ��.X7���t��T4����/�mߨSy
��5��X��Α�"�tވf����u&�� W	#�Q8WwN��� '�euDe͊�H�r�S�&�0>�O �,��$��ok�\x&��/�u:e����m{�|�ը)��V��o~�S�ªtvp�ǩT��C�_*D�v�M �d^���|��V��Ǆ��)$��+}[�v��Hq�:�w2��ϭ���X�p��A���}P+�km7(�d�hh��y9�C���zP�4oNqC6���-S���`�N3*5V��t�O���wlh�1�Ml�wH,�0
���B�������v��6����ڋ����o�{9wC@""�S>���cf�)�P����\V�,�ŶVZL"��d���,k�A�rł-����TW�I�3u�-L�L]1vo�eN]���m��v'7BSC\%2�%85+E�Z��k�)6�a3��܃���q0n��`�xTuk0���8���k4�T�7l���z ��+6b�u���x�o����ngK��,Fs
��99�P(W���m!��*��m��9g�Ѻ�l]�-����XL"���D���{�'����>opgGU�-�v��o.ܲKy�D��L,���*p�]o&4�W��K9!\0�9@�!#\-�r_b�Q5սk2���BWM����[@�A����)�Xv��Lh�I �R��ٰ۫O4^��iY�PkʝN�T�2<[�ǈ�euݢ�n���ƐC8����]ǌ6��Z��4�vt��t��ow4�ώ2��%�!3M�>�[�r��X�X8%�!<SJvw�V֮�%��)���,��D�˻�k)N����k�(�r�X{��2� �����}38e+�\�p5;�!oՕA\]x�q�""rb��A�������l��F��u9��m(���hYK�o�*��t���-�<d}�T����O|�|�z"���l��l�i\��2�U&"��J��(�UA�-�`ũUU��*���TUX�\f*��G0bۘTUDq
�����a��DUH�˔���-J���+T��j,Eb*��PpJ	Z�%�\��$LlX�ch��"���`�PUQTm�`Ȫ�%�X
����j��DXT
֌QEF�"��R�����,U`�mF*�����H���(�Ūʈ��"��
�F,TDX*�������TF���*�TYh��"5�`��V
�UdU*�Q`��Qb *���eBҫm@EV-e��ƶ$��m�*�Ԩ��b"���X�U���Q�(�Q�5�PX�> (�����҅8�o<��4em[�6�Y�o`��w�Y��	)��:5�ǝs����`�a&Z�v��0��5�|r�}�V�B�PK��neC�O��lkOb��*O����K�;�[b�c�-�kS
����[�'"�q����Ԝb�Y��ʚ�"�۸��q���`(UղMt�Yb6�>vJڳ/+�*_U/�.����'�B��׹�Bܧ�&���F�*�'O��&����Y����-�ؐ���͞�/r�-���ȵ�kVR��w1��'J��Z�V^ޝ���gĹ���/}.vK�eғ�(�^�kX��52i��,wl�vIob�;�|p��,��&�>1��m񺙔��U���'�S�
�cq#-�޶�9�/X��a���F�H-΋� �@�L�l&���U"�:��-^��k��}]�Z����6s�P�z�>��U��ٍj�ut]��wg%۴-!�r���2wx��d��پ�-\71��n���}xj��B�%���n��,����9X8BX&��=�!��8�}��mf�'�]�pf]�4�ܝ(��=,s���4:]�[��y_35���o5�\���K�~[Y@J�Y�y��zYO{
���..��,M�w;��x�i�&�r�����i�\œN�Z���[�Y^����N潼)��Oo}��WD�ӏ�7��{���ʻ�I+�:�Ϊ�m.�o9M�]���F�<�P�v%�5�)��7-�$L�QZ�i��-_ØY�{�EBHr���U5�5��*��z��nI�/�(7�}��s�\�W�v�ȹ	�Y�w���Jǥ�-�5B��˽W=��3�s�!s�;��7\�Pnsab��Jm��c��;Zű�U�:]f���wbf�]�(p�&�r�gbr�޸��v�O0�0/{r�� S������"p��ܵ"/{�v��9{{)��i�t��V��8��?�n:6^�a���x#$��^��$$���w#�����m֥�4by���UKc0�W鰙�t������ϳf���ug��ؼ�uwv�|�,��omd�K��k�'M�\מ&*ݯ���ҟK�i9�lR6;QQ�799��i��\�7/��E��t�)�%lH���;k���c#y�}�t�G��穲��21����T�K��B6�r9M������Ћ^��^o�r߂�(��帜hH޶�B�Ŋ]�E����<�8���[]����<t�7���>��]e�oT>^�ry#v">�:�K��3(n�M����� �^"oԡ���Nr�/�I{��6xͥ��q_m�=>9�Չw����4F�-yk��S�0.��U��4��e,���˚�77�Re���7����ޱ���ܔuT�Y��:��܄����yG�Q���g�f��ѫ}�8�D)t�;|t\�[�@\�-W����7;v�{��b���3Z�=,9+���ݰ��ዦ����I�Oa�[ݒ�ء�z���!�n����~��$�մ�;�1q�UL�5�j���D��FBً]F�;(��t��vXB�@5ID�+��.rd9��˼2nhD�@q��#p&�f�Ë������P%��,��u8e��]bf�n�끗�#pM��9�R�=�m�����s=�t�ӱi5˺��;Wwwsܛ�]G�f������=��t�2�p��n�Ć����~��t�s��K�W.��q���í���S�2ʑ˲ة��w�@�\�a���!�ˇr7���S���3a����ݺ&�'�_5�l�*����i�߰���*���y�t�Ux������.�D���b�K��[Cy�c>aK��h���H;���y8D���=⻍?MZ����#��=�i<W�|�b>�a��E��޶��J�v>RP���;��j�z��@+�3�Q�iy^��/�ޞ�A�v8Z�WKYK����F���o���	3yOgV�>��.�/��{RN�1E;�q�\�چ�����f��K��n��o�/mc�g%ķs�{��w�����.�4�Yv.D�_L��+{!E3��z�zx=�+��~ڷ�դ+$�}�<�VU�/����x�{S
�g��V�ͼ}��竴$.Mvnq�ƾ��aŨ��8!{���
B�r��قT�-�ڴ^�`��b�6o�E�8'�D:�"S��.��F���n��Z�Y�B�c��_%���-4�^u�(�a�(�Ϫ���k6���	G�\�q�׳�E�t"����ͯg:[y��v�m�|��X�V�@��z�IYZ�V{ky��3�Mv�f59��`Ҷe<{_'��}ҕ��{���Ŏ��gĜ�fz��R��W�}��?r}͎��-��|�9V�-6�ܳn��U�7\�u���~�UB���R�1��u�̈́�3w)U_Q!�=[�2�w������5�ek��t#������w�;茉0qK���ک�Z1��3�)dr�Ҷiĭɴ�;�7YR��z��L�}HMdn�3�$+�9]W�� �sgc>-eKh^t��6�ʛ۾��aa��r�c�z�]�bE�m��o�!}�ao��w�sΏ0^4����Rω�e�p��tFa{�:f[��%f�n�Y�	�I5�1�<�+��d��;�n��'Z�^�����Z{Au�z��OC}F���S+#Q��]8m��-`�닆�}���Z�:��p��s�I��-Oy�ՙ���A���uR��It�2{Zu��jAl����ն�'ׇ
�Kd�g|��>Q�hN��':��6�'�Vm��!�ti���']�y����י�-��R�]Q���,��r���nm���ȥ?G����k"]E�|]���s�Ob��k��&�unL�2�M�24�M���g��&�73��'���6�蹕��rto7���O75w���zG���#�bL�
�P"q�e�k���x'ri��kcbg�{�d���ZK� ���]em�IѭY1�*4t�1$��xNweκ�|�qj��;2�8�v�q�TD��~�HzS�U�+p��{އK����K�в/�6̗"8���W=/��)U\z;���J{�Ds�!s�	��ع�K���=B����1��׌�=�t�KY}�f���MN�N�GA#�䓵���v�5��:�����Kٌ��F���H��~��>��6˜l����M�p���k��E��4��*k�����m)N>F��1�ZP���,�e�3'N�t�;{�,�U�W��eOh��Ds����w`B�˄��l�UVt5.�mnVs��4�����'�r�!K�ܱ[�~v_���y��Ƞ�M�m�T�l�[*����Sc�'�E'r�i��AY��.].6��6/r�+�b��x�j���cS�؍O8ɉ���0Ef�_��W8�F��ﴟmZF@Ődbs����h'/�В�]�����K�"�ۈuo���*��'؁ަ��ʘ���c��봷&���qT�܎��T����tv�9�b\U#*�6�;w~������N�H��3��cjr
m�}��;t���eg��O����%�i��9&��	Q��{�du�Sۅq��=��Ċ���� ec{I�:����j홺�U��2�m
�.o�M���d��75�g{�O*�K�z�T�]�I��B�9��V�xkB���8�1���/��E��	�pw90-��b:|	�$۹��=����R�F���Nq[c����k�I�ol�u�'ρ�.t��X�$�X�X2�u�p��E�Y}�ݔR�9�v�z�N_١M8����������\�yN����iL��u����W��3���9�W�&����<���Aם>.3���3|%q�f���z7�x�r��7Ҳǣ�¡���4ODw�k�Jx�B�x��~�������h3z϶�V��p�y�N��F����8�G`#y�w,eG|�X�h�3yK�4�d�̖�����΄����J�g�'b���/����A�Q$
�uTf(����{Ҷ�ˢ�ؖ�U�g=Ǵ���l��/��8}9ģ���<7'!���/�|Wi�/
���l�\�F����^-��G�qAq��C��J�#>>�^���������0�{�m-,v�ɲ}'|tԅە�Eq�9�\{�%�R�yE�騯��Q�I�X�=ui���!�x刊/Q`�;bn���g����r=;.=�Vi��/�!q�2NRԐ��)�������n��>�(�yĞ9L��!x��Pw�m{����3����H��9�B��*��Y�k�n��6�lۜ2�X�o�V�7Ֆ4��Ty[pu���q��oP#{o.�2�+mu>�\�k;�7]>�Jyr���C�pݨݦ�R��n�6��ǳ*Z��d³�+<����Jus���WY��Z�
=��Wя�wL�H�2�ؾzk"�9(�̸Zo��q�3������ع�WΫbK�t��l-�����c@Nu%�p���i�ΛF4�z<_w��ȫ�̍�1��g��yE�<_�}�c=:�����n���
n����=�\�s���r�=T|$�j��z2kK�3�67�D;��R�1�-T����:�{��P���f�ՒT�z���n�De��=�����T=ޗ2gY�G.�f��x�=9��|ĭ����T��v���}Vs֩GZ���ٲ7�ɉ�%��� ���N�ҭ�����N-�����1~��j��+��[Ӄ�B����b�D+�gY�(A؍�آ�)*x��1hX��1�x^��|����Sg�K=��v+����!d�-1��!{��^�׌�7����i6�?��e��X��l��uj(3g�n��K��fnf����sC7c{T��}�>��F�.:͕<�iq�-�Q%�x�������E�Ŕ��1n���kvr�3dk�& �wU ��V���bv7�Cc�v�Rݺ;Y���>5
�*`�$�5G�ku{��Fq�=y���U�s��+'&.�z���9��v�ojP��vo��kv�c���@n!M�41L���q�ö�Xꓦ�����F$dy�ؑ!z��D���W��t]�J�P�^Gсם垱����R7�����Zu����d�Gy�+��B3������]O�R��^30��ݰ���@�;9fo�L�׻�������Q�k"!��#�R��&}�f��X͠���l��D&�9�߭r�x�Q�����P��獎���R8�P���&�f#��������w�<F�{f<f��r���ާ4�4������3ƪ��/�'K����N�<��8�f��g����U\���z���	T���z]���Zo�s�5�N"�%����z��GG�y����z��賗U��=��4G���o�/�nv��ϴ����Ӭ�g�)�/�ӈ�O+���ҷ�*��^\��B����>K���~�蘿�lP����^vU���[B�wǵ�F��uj�47���^)F����SѺ�lw��F���/E�x��ͭg��{%u����<�}��#Z�|����뮻��~�{��+�����x�b�?QEi�+A��ˈ�&t��܊.}��wٝ�Df���2gV�Eݱ%@=s�:�H���qkT��4Z�R��'n�V����{`��khp�.s��Q��&Ӈ����|�Dd ����+�j����ﲆ7���.��e(N���qn^f�4S�u��ǡ.πxs9���k	�/2Dҭю�o=�Y����f�d��=��u���B,W�]EV{�*��\'G�!��; ��z����Vhݭ��K,�-Hں!fd���8�"2�w�Rt�����2��[Ɵvw�vX�����|�ُ&�.�^�vd�rmAyԣŘ
�|҈�ur��t�ݭՋ9�
U�*PUIq�z�Uш=}M>���ә�]���4F�hs-�ܜ󷯘mj��::��M��܎�캏:bT�Vdv��a�z�Í���q0�m͉aS�;1w+�"�He8^[�����z�,�:iv�k���wk���c7��mѷ�uv��xu�N[2���q=f��:r��O����z�����+��p/��r���7G�^S����Y/��Y�dj�q̴˚�J�m�N�=��7}6��r������s�n�Sn��J���q�B�ur��:׸()���7eh��������w���ު�R5�<��΅���E����Ҹ]aֺr/�]҄c.����Y��ΰ�t�bG7��ն9�ڈ!�6a.�M�����(�Y�T/1�┹���4�b�m;W
F@���JT�;���(Ju�S�F���66� +�Z��J�!�k��vd�%�
�5�
�b��]�Y�����!XV��T��o�k�TU=
��+d�c�'vR�������D88��,��I@����R�IrWv����e�s**{�3B8�Շ+��t{��m*AXŗ��f$jp=��%$�B���<sv�Cɫ�����Ӝ���{ n��ˀXb���+:�\h<ڴ��xCW$���.|Q�e9C:8�����@�{�r���Q�ݠ�]fӣ�YN����v���;�7A�wz>N�yi|�s���ՔR�f�׺�=�կrZs:'I�P �M�N˾�:��8�j�ܤmeNBV9�:����bI�����4��
���6�v�u)pޜ��J�Zn����91�fR1�7]r�/j}ٚ�4bx�u7W8>��{�{N���r���]�˜Ղ�W|1H����}���!7i!���R�6�ܵ+������}����a�@M�'�}�lD?^�{,�^�:�'����+ǌ� �T�.���ڙ������q�(V�!���%t��p�zU�R���#ڱ��w�"\�3t��K�p�	�!��KZ�N]}O\Gue�چwV��%���|;�Ӡ���j�i�|T3;ֳ�{���םg�}͡�0b��$XV�"�"%j�Q�V(���)YY��+YZ�Tb�
��DQ��UE`"(��([V�� U��(�B�J�DeB���V0h�Ȩ�@D���¢�Q�TQTD�X���"0X��B�X�EYPPQ`�iUX"���P�BT�FU�*�#X����j���#QQb"��	�[b�V��� ��#X,D�2,�%
��+("*�b�QV
ȤQPV(*ň��Y�T�#+UTDX�PT����TD��b1-���ڱb�T����AV�bȤPcB[KlR
�QdQA[BTw�<�a���yl�[M�5f����Pc�v.���7M0��M��G0���E�ʸ����K��%�I��[\��c����H��TQ�B�*��>��x�w�~����V-��z��O[�
^�B��D9쎥�k�<*�5."@���SЯ�֣��3�E炭ӏ���_�y�yd򗑛��G\D���㶜vϏ���q��S	H�6<},e(�^��8��fs8{�OE�c��kN{�/��x=�����@m�TD/J�����>C�
U�f-����[�w�K'�}�}�iAy���tP�]LP^�6A���&!x�jD����wpd�_)��r$澽��^�/U+��zx��D?nT�o��"8��8���~�
��|=�s���F�Q�����+=l�i�;�+r���U⏥Ǹ㬨�a�n"���Ro鑱��}�e�ώӚم�kRZ�_��ur��P׵���P	Y��:�܋�y�yΉ#�U$ܽ����ڧ˽��$o���Kv:Z����<����t�8mQ��yLN�z)��2`V%
y=n�:����M�OY�%q۝��c+t���i�s�3�N"7�z�ЈhI�ͧ�2u_G����_^#�EC7l�IKA��wt]0�}�����o�&鼺�_ў�����3��kf=Ӵ��L���\�by��3�*0��w09[���Ũ�����㶤�6����P��wL,��s�r���⍥W�e�pۜ��]����P5_�#�nь��ndL{3���Aw�b��~�\S�a߿�яW��9=����rޖ�#�㸋�(��A���Y��c]��`a��Z���n�W�^yf�.��*^�>z#zls�k�~&Ƕu�z�q�_P�7�s���:v,K���w�^�c�vmz�3�yF��ٜ;�gT��0�6:��6��wKuج<�G.�!�#��^��Nr��1.W�&��T���Eg�d�,��W���`�-������߫�s}Yރ�U��ן+�o��4L�R_7�S���y�yc*�;����U?f�m!>��u���x�oGU��q�%R�E��!�xé�ODw�h8�M�&���6�G;��u&���^tͤ�V߅�t�>�	q������h��?'D��;����*�F?�w���/t���XL��#8?RFϽQǙ�z'c�^���̹>�1 ��g}׽,ǥ���U�|r}�t,7�e���ұ6%����8�p�:]�r�L�1)�~�u;1~�Ф	�H��<�N�v���A'�#��R1%�y����{��34�	MƏ�K����#z?No�����Z�v�%�&\:���l�'��sx���Vn�����t;��Պ�
�Z�j�4jU�&�7�.l�o����a.��}Jy��>��pAxhw/[�ze�HC�W�o��؇��T����Z;��Ϳj���T�<O���v��>��'�j����}��K�JjK�	����C�e���(F�ޏW{�F�䛈�x刊�4��ϸ퉺�en����{K�꿺��3��$E�Ǟ�J�Yy����{ި�NLz4'Y6b�I�ʎ�5	��7h<���ZZ�dHQbo4K�뛟&��Q3�7��ٗ���T�ǺAÿ|��a�;S��(�	�I���Ȼ��r3�~g
:��hY��UZo�p�g����`^��D�)����X�j�'p�O�Nɞ�\v���מ�^�]te��ZU�����}1����\GX\�En�����o�X��Fp=^b&n�����{^�%��<7"V���>YU��ɭ.,d�����#]��w���a���W)��罂e�n{���F{�����]Z�˂��>�z�P~5�+�2gY���ʢ2�\��Q~�5�oz�g��W�W��K�Q����(Y��J���)�4Ew�=�L�#��Єq���4��1�ӯ�:�$��Nw6kOV��ZM6��
۵������.[C)u���ˏ{=���+{>����sη��K\�޻�6�)��VQ\��uoe�/��t�c'XY�՛ex�G;��9SXetV٩P[�Fs����r�:qK�fW����c܋�i`ql�`�_����8��Uz�s*�3�鿨��w���z4Qk.�+Kp&��,ޝ��5�`y�X� ����%�ҽ����=~����e���{�0F��wa��8��|�/DvL��9<��.<��˅Bھ���m��5��x��^�v���g�K�}=�-�u�|A��B����^+2�m�B���j$����EϭFL���צg"�k�y����g��|��Y����(�/��Q-l�Aq�	�G�z���(��������)_�Le��~^�tG��dh�^6"�X��|j�$
}[FƗ��~��ЈnF����^ŤeG��k���D{�)���c�ۈ��(�}����o������VW�u�V�r7�Q�x|�C�׮l߼�#��Ϊ��\�>gǧ	q�mew�;>�u۪��z���aX���6}���q��b������ޝF߶�{ڜ5BS�.0+s�{�k3;�l��}�;N?f�G��'b���?��n[��Y��9�b�9A+�az����ɧw>�۵�8m	��[Hy�ݳ�o(�V���|5\��AAAޫ�.��n&`�v.C5`��zA�6r�7ק4|k��ܾ�3ŝ��ϣ�no\��
TgT�}V[N��\���wl�Nu-ْ�&v�]Y��e��dO���H��L{������.,f�i�5�F���G�z�C��W������{�9-���~��r�����dN�%���*��C+h;��:�F:�o�8�toC�QcV�yf�����d�z_	w����z����)`��g�	��J�P���=U�>��׷^��|�zeϵ�AF�:�����9�T�Z�찑��סr��XɈ���p{�bf�}���|���D{�a�L�y3�7�ҫ��iT�����)��u���[r��
�H�n�Oߴ��Ηy�����b�7���e�BG$�}��c��U�v<XW���ȳ��P7n�ÿ`��s|���^uZG������r������+��}��W��}��n{�t=��
�!�R�+�z�m;�F)�nb:�RD/OY�\}~�{�aH����nu_��<��i��u�ߎ�r��z�=��g��řPc�h�����������+��ST���>�;����OK���쮂���؈v=�sn�ɋ
\.$C�M7A~��D�Ğ�����Tzl�ʷ�N��$ě��e��r��a-�M7��/��NY�'lw1����cЕt�\.T$�M�Y5�v�=`��Ķ�_B����zЗ���WH:C���n<�':vuŹn����t!�t{�'#�>�f��ϫ���>gs��;�>�\�hz���͟V��:�*!��u?S���ߤh[��>�ݪXH���8V1Q�W�+L�}�����A+4��znE�Σ�s�S�������!��X�2%Yw-�������.G���z���Ռ���'��k\���%�5G�
��U
/wn?.IW�j|�\<����pz��\t����!�ϴ�zz�师�X�tdB��]���za�w��R�tyuT��1��U��F�tڙh������j��*��
t�۱Xbﯻ�5�ǥe(��]�"03���Q��={�w��	�x���3�����w���ш�~v�J�D�ᗲ���*#\�>�[��>��{��z�Ez�	�eN��Ln�C��N?s]>��<�ת�=Y5��2gT��\�sc�j2Ƨn�P��A��A��nv�;�잴����>�d���+e7�w���ߎե��sav�l�`��^G���>{L鬡�^Ue���ק�V+�h�;<P��Tتq�O#q�M�צ�'���Ѫ�_�i ɚ��%����x��2&]b(ě�7���K/�����go�]R�Q5��k4�U��Q���B���z�8��Gq*�Vz�@�ջ�3xP�*�g]<�V]�wh��1W�Z{V۔6��,.�(i�#9��@dUqwH�峳C���g�t9�=��~)C�
z��é����4O��"la^/k�x��O#bK������|3�5��zR63�}���lP����UP˿��s�Ί3U�ž�!�/��l�����4��M�/֑��L#���蝏e:���U�/ �6}����b<�~��V{���(�٘�y��߆��M��W��ģo�t����~���yq��.��'�V���Q�����$/U�14�v0Jӹ�Wܽj=���+�>�^�u��EB�����wW���#�-�5���(�KGnn����"E5[F�ϸ�}�PZ�(�Ҳա�Ǚ�Ҫmm�#wׇ��f���W�؈��plL����ו�B��t�������o{q�DӞ�^�쎏�4���O��΢<�9��E�6Y����\7c���^Z���t����oj-��2f����wu����x��w�˱+����J9`L�ZO�N{��A�qG;��S^��E�oVÿ�v�v<����q�=���\�%G��hO{*P�T��oN�Lf��m�����5(��'\@�euӔ*�N*�C�#i��y1�E�l\�3Z%f����n�j�,Ǔ�z���+J�fX��kqf��q�����6t8p.{a�3�C�˳�����+L�#œ%����8�����}[�4v^��<].�wgg_�Kg���2,z.ZxJ��V��\��lOm8�����5�A����[^~�`��v<Q���'4�dN鿤��T�(d֗�;�`k��w��7�[&=ӓ�G"�V>v����=�;+��'���yu�E�Ȕ��.#�h?U.�~�S����y*S��T����Ő��+|w����=�>�P�{1C�������ߤ�jnh8�ް�z�Ϟag��	n�'͕��ïu��]{N��Wd�?S��藎z��\��7�MP7���Tz"�w����=��;W=��욅������/Sf�~T|Z;�z}ĿO��+7<=�~AM�.���+s�O��빣���&,Ҹ�r���	j�&���F}�
��q1�}�v�B�>��oM��wq��s�}�vÚd��
������@�f��S��t�\z/eV��gv���_y�Y���LƱ�C#�h+����D��D����8KGt�rΉ����i���ƥ��n�N��p��`~��w��pLW����Z�����$H�մ}}� ��%���?��E�휦o�)���? �<=&/i��B�ු.z݀�-ph;^�=H]���
���z�lN+$�wv���5����[ڒ���ᳮ��#.<r>���X��o�U��On��G;�!��ޛ�y�@*����dD+~ۈ��(���vٛ�^��>�0�{`���![1��NM>��7�頕���͛��Dy3#��9RMyω[}q�㔚u"��Y�o�ԧ��	��V3kc�u��fkK�e��5�u�D������<�GoϪl��弓�>������z?X��>ñ8tk��f�-�W,�G���,�w���9�DX[��x������v���'���9��^W���3�F���X������Q�Rd���S)y��K��j�;=t�b��[�ȝ�r^,A᯲������k��Z�OP܇�7���	��07�׉�S��'[�^�Qу�Ɣ^d�t�zf{�yՑܻ�s��W�KÔ�,���.�K���~�{��+�����s�:7�<���*�6;�5�2M��}�����Uz"o]�y2��'���W�X�߸珼_�|mV+����J��y�:�^ߦ�,>����������.-�VT�~��G�F|��o�����ǂ"�S�]w�*�fN�0>R���v�E�X�m%!��m�����heY�u�3;O��Gy�̗a�d��4P�~l>j����7�^D����=���P-��P:�p噢��a�Ig��Hϋ���+��QU�t�n:���8	���j.�Ҏ�kէ�V;Q�Y�K�b9mTĒ��}�ql�T7�D���c�i��{c6��:�����oޘ�����:u��0��'��J��W�a�Z>Ǿ��\�����RKW�^X��1O�$s����tP�[��~��󘈆���K����{<*��������	~;����4�J���R�҂�q�yQ�s.Lg�\>/"�eM5���~��Y+������~��ߧx����@�q�I�YQ
���F���M3[ޛ����Dv����&π27�MJ�ў���Zf+�s�=�L���u���nE�'�S���e�w�5���Kz�x#���,�a1�+��5y[���t��`�����C�>��SZz��w���߇�ꨞ��ǹ����`I\v�h/d������OA���Fʓ�4�ӗ�z��Dy{u�zf|a�����繑Q�-�ȡ�N���[:vC����z;�Q$E�����ݡ�=�T������R��|�=q	�GK�
�b�zkb��:v�ˌ�]���4v~�:d�f�UG�+&`͸ ��\%�L=Ȩ���l:�J��Y�ԗ�l��\�1�)д���=ov����4;�\)ͺ9&6u�m��-�:XJ���m�Q�[�4��tg(��F��0b���d8��ш���Gd}����NZD)��պ��m�m�y�$_T��g+P��q<���.̶���V�	�$�2�س�Ӂ��oq=8WU��VzT�����33'�emv�A��|'�M<�IAT#����@k���x^
[p��Tq�\���Z��or�yux�ٛї�Fu����{�Z�a��ŭ١�+D���m�+cxF=kkyuS}cR48e
kn�[Ҧ�������aTF<����'UX�����Ҵ�<��w�!�׼L��2��ԩ�c��]+/ͧD+�����y~���*�n�^�X��ɠL05d��6�4s�"�KZ;+��qʾ|R�=X�84��٣_Skww�W.�W�q��[˭��v�v��o*��>yL7�3_!j[�MAÛ�*��I��^��;�!�r|�@��!�r�]'�w�� 첢�ᕢ�שҩ���24�o_.̜��c<�4��܆ uI�n�F�Q&�P6���ۑ��vp���D�`�"���Uz����r��Ը��z=6�z;0����J]wGC���������G�{�p�ī�V�:���u��K+��^)H��q_݊�aJ�֚t�&�F��Y[Os����)��\Fm��$p;�-P��vg�P%�mWg�=�ޓ�dH�]	7|;8���(uY��CFQ��=XVHR�Q����>fS��(\i�T쬲���˺�n���0����J��1���W"����9�:BH��"��ܤ5o	�*�b��dB�v�E}�; ��aͼ�ŕ Κhi�	��d�T؋zS����	�z&�>��L�דk�օ���/��T��+����
�ͽ�ۢ��"�	1`� ��\����b::��ql��\���Pj�*V+�ݕm^��N��S_y!JX���l�Gfqo�f"n��{6&LW���#`%'����y�e�;�e�He���Ț�q*���и�;VomD觵��-V>��lc�zF����S����s5�����k����C�f���l�ȳ�<[Y�]=v*j ̸or����lWEY`��#c;o��N�$���v���Ӌ �sq໇\=C�Y=�C�Q�"#"��ϕؐP�)֕sU�J�Mq�"��Yyǝ�p�r#o���#��S���@��k��3�^�]u�*��"E��UTb��Aa��*DQ,FE�,�J�-*��"Ȉ���1-*����ePR�P*1
�0RT��(�T��E��h�DVҢ���U(��E�Ԩ�[DV,QQQeb� # �#b�kZT��X�*��`�
�a��,�V���Q��*�DYHT���X��UQX��UTQTUX��am�����$b0PMW(�,YR*�Y�X"�T@b(�Efe�LlE�5E�"�U�1
jʂ�d��R�D"���a�ccUm�Y
¢ň�jbLLB�9�<�~���E�yj'���'�%��i��!&�iy-�L�Ly���p�4{9�>�k�q�]��Ń�X�e`����ϧ=�f,��\~Q�=AY]S�K�7�}���W��\�O�-5C�����+3�2�>�
�y��^��Q𝜂�Utz�Miw�;��'+��jv��{M��[��e�{�|��+�ME�Fy\Y�����'����6-�|%��2�[#�g6:Ui��©1&��������>]겼;�>�:�T|GX�3Ƅ�2��D�� ?��=*ۭ�>�����"���[ɥ����q৕�o�Zu�^�	yJ#��o0�h���X�)�D��;��}Q{�c�yf��K���կy`�~�͍��{���|����;E�"��Csិsn��yn]Z���3���&;���)���hմ�I~�����}�r8e����Qs�n�O�����tm5.#Q� �Uʪ(-�a�/ƭ�bo�:M�(�~������J�ow�.[鈵*LG�-�"B�t��{�#A��;�\g/R�OW�Yεv�{�wDGA�����^r�fL��ȇ~{�mωD��ۛ���H��h��wdK��{-xj��\�Y�:��v�V2S��q�t��d���2���۲L������zx����X2�&|,c\��r����?j���k7O�%&�5N{�z�$X�
;Y{a���s��v�m��U��1,	�ӲʙsK��z
N�*�,��B�r��H�L���é��=+'C�Љ�-��������O�ϝǔ���w�*�E�PlL������0�~���Ww�'ʐʣ����ǫζ6+����53>=�:���5Q�f̘��x�̨�f�x�z�����>�ɵY������Z}��3@m�I�_�US�������F���J8���޹N��ɩ�ޝ�������q����������3Ӓ�Vr��x�,�<���_P���(r[S9��9�'2n�����6}�����"��\�OO����爿�w���J��={�3蚯_��ɥ��[�����z�爵�;�ė��e��5���8�F=U1��둄"������o>�c�'O�Q�o�[	�u�E����%�=b�?U.7&u�[��C18��eY����˯	^�'��n|7���=ޯ#�~�G_���m�~�P��RaƩ2G�h�[qx.��������8�ɑ������.��B���پ�B���8��e�V��׽3�]W���s��zbO�DOµ؊=�&�q����yG����Y�8=��������oߟv�)�'��6$K�m��
w��v0�y�wգ���~�Q��/2RI'՜z���~k�?6#v_Xu����x��'��E55K�v����Ӣ�F�]sU��v÷SLQW`wYĴ��v��[���Ds�'����ޚ�,7�7�gP��h*�˴��gsU8w�j�����u�8m�|��f뛺R4��.u��mWP^�:T�E�Z4!*�����.W�g�>�_[V�lQ�d��+t�\;��z��x.�E�t��~��1A�9��G�D��D�}>ä�wsu��x#1���^��Z�ǣ@�:�6<�AVϯbm�"���WKgo阇ƅ�$_�^x=�>�ϭn�/
���4��!a���z�׌yLG��k"!?eDm�QDؙ�v��� �z�����6�y�_��
���5������Vh;���>�� �_9��	�]��ԟ��Q�R������W�*���p�6��.4���\z���ڙ�HCܪx��f��?��EV����ł1d�o��N��^���v��z?^N����V�.�A�N"y_�z+�H��~�������w�=-Y�k�Wo��9����_�^���l֝f#=n6]�(K2r�N��c��(�nVq�������p�#זi��v~�x�5��~�[A�������_�Z+Q<�a4�k���+;���Q3�v�=z!�J����6r�'k�k���Jʚy[QtH�X�v������W��E�2w0_.�#����d��j�).cJj�'w^.�G+$�gf�[�t]�t���F��>�oLF�U7��2j����z�~��?f�밸d��,�����z�z"������(�(ۺ��3�o��c�ݍ�~�q��x��~��o�]�g{�Q\'JN�T�nf{�����Pz�S�����Xɔ�_�3�쩨\��|w��=�>�O�U^lOs�z&�2����Q~�?՟�������M�w�gBE}�*�޵�g��]��V�BK��Fw�R��}������%��%����'�JG���W���i�����bA��[��S��ǖ�F�)��t�����S�6�nx���*"��,=�\��Jt�����L���y��__�#1K�$p?m(/�F6=t꡿W���<扈l�MO�J�>�q��"��������4�O}/��8��
oױ�7kb���&7+c���� �{=Z�}^ؼ>
�B���Oi܂�wN�/M����Ux�7��*nb;�O��T�[���%}Ҟ�^���t�C�&��X�0���b��;��ZTh6�M�ޚ������������h�#"=����kV��}�����J�܎��N��rR��Qخ�S
� ��j����e�h7���#�����4�S�6��	���-���,�ӎ��9��I� �n���eGc�WH���n���{��x�����bU�3'$�o�r��N}%i�'����j�K����5�v��C�p����^8��!{(�xr��_�Lk�^��Xg*`Ǻ �������^���Hv3k�W�G�}5=q=��w7=�Ơς�Q_w�ߣ<�^#��/=��M��o��r����א�?[����~^��~��?�)��c�L1��v�/�`1`�ʶ=�]�y�ذIӾ�g���t����wy�>*��(�_�����Oi�F�o��9w�įl�=��XH��+���k�d����ċ���ZlO� ��8�����H������S��޴�D���%0}u1b�3�rѾ�>�V=���VQ)�NA������ig��KGJ���U�o{���܏y�w�J�>�4{o��%ڡ��u��D�4$�7T�&�����P���FG�n0�{�եkՙ^���(����{�R;o}~�}��h�ʝa�:�'b;�&��[%���[x�����.�ȟ:���hy~�_3�l�zu{����z��P�Jl*y4�1�ɬ���'�(�����S��Xs�g�R��G	��ּ��ÝYm9n�sU
Y��m⨟��j���)�=ynU���ߪ>Hs}ܑ丗�zv�����׍��s2p�����aXb���ˮm�2��yQc��G@n����ԕR���}1'Ĝ�Pl9h�pm�[J�؞~��x�:�"G���Y�{��Y�&���eb�r�N�A���_*��|���i�/�[J�ؗ���%��fٱ��T����c�<wڲ�+�N�E��G�D��Dȧ=㱇Ҵ�Aq�9z�x=�5Z�[�/-�#�er���r!��d
u�Q7%��7A���&���c\�;�v���Q�����Vu%�쎻����ί��G�s�Q9���2���>�&�>��!b���W�W��+U���g�O��걝~��U�UO������׾r��������ԗ��w�1���k[sl�6��c��%����}��m�I�_����H8t?"kʫ��B=1�&�X����i]�׋6K���	�q���=c'kfƗ震���^����<O�,�s���g�
�;^�bK��ܩ��Y=��ңnv�fһ�Ei���o��e�u��j�O�S�0|�t���6�,�y#�wgt꾡>�}�<E��;�ó��U8�3�Ɓ�;��c~��Q7hW+�|�F�gtV���$���jv|�y��7���b]�z�]���R�U��˵oekM3wj�A�)�Ѥ�Z��eGz�\�}|�uI�v�g��v�ku�2�Z���k����c��S���b���Įi-��}d����Q��ú�����|{\�u�j;�YD^dJDò{j����Uf�J��b�W�h873������4���N�w��u�~�G\���eG/�L�R\%6�?2h�������ȏ�a��ZT���]{N}���Z-�tXx��.�gT��R�u��3�G��=����r#:n���^�y��p��^��JF��|{�>�q�u�k�nFF���w�Oټ���/����_�Ѵ��O��3�\s��M��m�~�$��Q�P�v���=Ć���'M{-�y��. Cf���	^++�4�U�Y}�����o��v{brg���������Ҟ�	�\����- ��H� S���΢�UT��Φ�ӹ�������JGЄ�U���R����!߷pLU���X1��x��ٍ�y-�U��Q����D�aZ�5��)� |� �J"{�q-��&���"EL���v�����|�tu�яU��M>��7�餬�v�͛��Dy��P���lI��IGl��^~��\���w�5]�9�}�;��;n%��
i���^0�y�vl�(�wU�ݵ�L����m�����v)��p�u8D��;q�y�#w�ܮ�׋��6]��W01N��.>1ﯥI��}��ϡf�C��.4��������w^��`��Ȟ=���zp{ܰ+��۱>Rl��2��$��;>��2wO����z����q�U�"h�)ǖv�K�K|:;gz�x���K��x~��8������3�=�#J�����i�����=���=S�:�7�#���q����'�6V�b��z��+����?r�v��t����s�.I��KKBI��S�|5LF��m��d��:�{@N���{�(��(�ߞ㲵]���q��__�2�;�_K	�<0�7�S�������)����{���x��bFH����:��`�~�^����&�u�K��Z[�{J�iT������#G@���S#������b�q�V+���+LAG��#�U8���b���H�T�w�z�yE���I����}��*a�q��q�/�=h�B�ĺ5���uS	H�>���#.3�����Ѫ�����?�j&-���w�Zw�&1��~��8z(1��d6�R�7�B>��9o-�������
���w(2x����U���z�N}��̓WnaG��m4��l,����'[W\�C�'�FA�v�ku�[f��RJkډB�M���I�β%��������yY]�+�IwjIU�YY��U���%��>�c�%#���I��iAy���aE�m��3�O�"<��H�ʓpY�Kȉ�qx���ވZ|3f���{}�"C�˽bo�}~�ρ�WAX�{ە0������k��EV�ym_�Ly�G����W֨�Ӟӹ��b��^���U�~-�I���~��s��Kږ�#��-��gģ�C�&��g���r��k;�_u�+_���?U��1t����t�͘�J�p��T�K��+I�#�r�9kc�g����D���߮h���%b{�;ݕrTX�}�<�M/MG���DOa�������!���� �PNO����>l���>�;��#yg���3,���F5��c9魎d�_p�q��f+_�k����r���ڭ7��x����"��wa9�x�V��Fr�HY�JY2p�n�پ4i���_����>֯㵧�������n��,mUuC/<�Z�[�O�ݳ���I��b\��Q�3���3��c\�rf��}���ܣ�g���7�����Edx�5�r��m�7<~�tx��s������������;��xqp+���{'�yK!5eu�)f���v&���v:Eu��_��V�ZU��g=j�=�M/u�����H�u�G6��{]"�?�a��Q�vyz����p���%�A�G�\!�:�Я �J�Z���������T�+�%I��x��b�O�V�f�u���(ԟ"��S����B�=D����F�y�܄��^ڠ�a�{��/Ր��	\y�}����� �a��K�_z#��§q�NyFE�/S���_�2o
��솊�~X=����giGv�Q=���8�}O��t�3>�{��u��v#�6(�Cs�s�����hж���/֑�zag�'`�v��W>��L���ռ�z�=��Iw#�� �t�TP.|�p��}��k�iX�T�z����.�N�^��I(������Y8}���я�2��gȶz�H^���3N{�c�i܂�=>y�����U�eb���Fzv�Ԍ/)zg�pB��5���(��KGnn����"E5[Gf+�zo0�ņ�mߦ�y	�(���4�o]Y.,?Mx�O�ӟ/N�z�{,DW��%���q�t,�w��5U�{æT��^�Dg�ޥ&��>���lPJ�8jf|}�1�5Q�8h�8��4 E���޻�{V��]�k�t�=Ofvh�V�-�=�vŶ�S\+�D�E�҂������ ��ȹ��V���o�(�)�,���-�A��H[�iͫQβ����!��udh��m�L��|+-��j0��t
�2Y���e7d���bO�t�������u®�]�N�z� ���ʲ�`|�������L����%K6��b��k�	�U��S;��ݣ�ʨ�.�F��(��H�l���(����f"�t8a��eN�ps"�^��+�FE	u�<�6�\ީg3�-�J�=v�S�uk��Q�(��=���Ⱥ�h{*`���0�$+"z]��Nƌf�9���Z됦�������*,I㻾ң#S��t�=O*L���(eX��+�5�i*��ߵek�HMw�QxU�I38<heeu]��J�V(ވ,��%4����LaJE�-�>��`[�^��S�[$;�m�=
'����V���u����`H�X]�0R9ò�I�@�J)]���ȁ܋����Qѱ'�qkM|+~�nb#5���z��+b#g_w�L�V�orA�m�V"�]i<*�iB�s4�^n�|�mE�J:ݾ9c&�tȢX��v��*.]m�]��@���d{'_�L����V֎n�*�1�6˩y	��m˛ǁǿBk;�8�ɳ�fw'j������MP.�Yu��#��G
c��\�#�IԨ�Yzغk J�LeΪ0�A��ɚ���q��v'�~�Z�Y��9���CwS�1W�E��3n8��+��Vm�v\��x�o�lve+`woRb[�4�۬��5RD�m,����<3���x9���v�-�7���lյ�_r�xu�����E�hⓧ]DMz%濅.�M����^W,X��S��RY.b�#��ӵ���z���T�j��ˬ=�y��sр�l���-�����M3X��9�h�y��E[M1'ASJ6K���P?:��k�Qq�O],)
PT�=��f��*uH��O�Q��4k7VnJ�\%x�J�c6��SnӮOe�Њ�f����QT�{&��% %K�y���&�qeY��Y�ˠ��)��rdʍ��A�HB8)����ں�s�ʷ����R�l'�R��ˑ��[�q�@�,�.��i�2�D=Z�svA���eEZV%F�b�9�����7O�������;�Y\�)�9ȭ[���ƫ��d�eu�o'nt���zX���*�u�&��s��˃��]M#1�꾝X��uk�s:6/��*�")ZN1��]Y����tĵP�O�{����V_Q��O���윻�fg_<'"�:����'��c2]4��C�yqV_4�ۀ�c9m9Ac�����G���R��~I8o3W�l'0��%l���3F(�$�Ӫ�$�vz��Vs�2n�h���\��WV��W)j���,1*���X� ��!QAbZ,�DAH�̱I�G-E� �%QXP�V�`��V`(E��XVLB�U1�Җ�FAV0���\k�Dd���Zֵ�eTm#l�ED�J1�d�FL�F.R��
���
�mdY+TH��6�	P�R�*��P�R(�6�,YX�J���,��Bcb�PU�(��h�V�X�"��ED���V",U�e�(�@EdPX�k
�X%�l@�,�Y�E2رb�Hڠ�"±�,��a2�,X*�����¥C�h��f2V��AAIE1�����,+R�U���A�	 ��u=��h���5�Fh���P*��I)�"·/�2�� �ji#6sΫ7"��ޮ{ZmL�C��E���ws�3c}7��{�6��ok�l�=���}��,{����uS�6F#A��`���:(�ό�i��[JwG�='����1b�U�X�ީX|?j[��ps�=��̢^tWli0�����=�\���1�؛[s�����>*3D�8��&��>�Ӭ�zxvˈ�T}��k�I��o.\�x-w�z�RG���5�Zju��e#�?�/	��	����O��N�O{7kn�����C^���i��z���WG?](���(��)��T�����"�3_��}�[Þ���%O�xl�x�L���TF�ڝ�9�u�{C�\�O߲xh������Z��?B������N=�w���C�΃ђ�]�P^*_P{}���l����t[�V�KU����׽�ԕt�d?LD��sQ�E7B0\�*�jO�`^�͏t�Wܣ	L^���k7{^�>�ʅ�|Zb1�#�ɍ�+���q�wK���}� ������aǃc&���l��k�ݡW3��:k�n����.3�f�ң�U�ex�Ͻ�=3��f+cr�+�'V�wL>���[�2QW��WV�����k�9~�*\e���k�nѐ�:w�n�Χ�����Q�b׶0�af�
�2��<"�l�덎`r�K��tD�q��E��#�`��P�v�T;vu.���}��؊�D�Tw�v�M�<�x��d����a���"+��B8A��H��]Y3~�q~�D�wg#2�>%���J�PN�>��|��c�*
Oױۖ&6�x؋R����l�A������8���ؑ5�Vѽ+ǻHxi/�X~U~9��qZ�D'�Q��>�dǪ5Ff��vw���2��fnu��0��l����{��IY��\ٿ��QG6�VMM瞃v���g)��aʒk���V���˅�9�ͯD�ˍ35�Ǩ%�����f�r<��fʭK������3:gO�|�0{Dl���^�g8Nף���9����3~>����껽bN���KMDy�x`������Ǖq7�{s�s��zKGl	�,e{�����D��c';�&[GÜ�j�+�������{�\3��域��g������ʷ�=,���#��Z�1M�\��,>N��=G����X�ulGk�N|�u�u��w��g{�(�~��U>#�ë۞��{�F�3���c�֪�Y3���Beu;��9���=���~��}4�
�y��`_�r�Z6Ѹ���j�����*L�X�
�G���s�(��F�=�gIa����[˻j�D���s�]�v�4���ue�gXa[Kk{3�/yl�"0G����N��|� ��P^�W'P�p�W.��v��B�+Z�ۏs�V��T�
X�q}��L�"�L�;*jt���1��+��ܬ*�=ƍ#��FĥC/�d^>�@.'H�)� �kx�tw���q���K�k�\�y�-����v3XU�q�}�ļ��`Gh�;�F�LG+���JG��q����sy�K�}޵�}j:3�t�7�{N�~�B�~��9�Bh�.w��F���Z1u���S�<[��=���j��Fb���8����f:({-�E����j�D����h�ת\eO�&!�\���+��h�p�ƾI��\��q�<ߦ�"����)~���1�\�����t���Q�7 ��Tbi�i܂�wN��/��w�{}�����F��SP�����>�k*!ߞ�E[�$���q�3�a��2��翮/�z�De�܋�7Sr~]����z�d���%K�.�q�]�}�\��k!���t�6|ǣ�T��D�=}����#��|�aR�\�E���ŏy�OJ��3�0b��"{�\v����=��^��]Z���*~�[�Pyh�m�?�[vڱ$c�醐�{���č2&��/���3Ϩ��k7$	dh̚Γ}�[�,{��~�=/�3|{9V3���/L<Cϸ���*�r�6H�����׌܆�\����z�-����Pt���C����\�N�������:]t��Doܯ����T�ů+1���]�'ݡXo��{�bs��<-�?�`_�O�exK����Pv3j��?���"������v�Ax���C�#��eH�iQO'�~;���2�V�V2|�oK��M��^���^&��s��مI��P��LM�W����s�~**�X���0����Q��&��'}#��'7�5-���S~���6���0"�����A�[M�L�~�c�w��p��˜��T�&�\Xɝg���*��7���6��{ᵷp�zi��{��q�~�xؗ���z��+�m%����<��߀Y�K��lo]������G�9�eP�ni�q�t�^���S�z:��q�v��0�`��B'T�D���勽1<��V�d��W���h4jߺǱ�Sg�
�%�utlS�����N������t���1�|(�H)WA�h��hմ�I~�����k��pk`�������Q������U:/ �6k�Apڙ�.|�`��i�/�[J���j��2����8��F��a��M:7���|����Vڎ����̄����R��uve��j��8x3�2ve7Ļy�~��cüH�ļ�Xj�]`�G+�P��͢�5� epK��K[7�կy�f%+�=��v��{���g_a�Q���(?Px���<}�u�@<�tb,Z=r$/P�D�=�+g��o�ש����Ӡ�:}�Q�_ޞ�H�^W�3��9�?n	�u�Q6$�v���>$ha׼�Qb_��k�1!Y>t|7ң�O�(%W'�a?U���Σ�.M�{�t"��(73�;�R��x㫟\Պ���w����㮓�����ѱB��n3�����{��ǣ�)�F{}�R���7�b�3�7�,�7�`�/�A�m{����3[A����_�US��t��z��=��)/���/�߆�N��ܔr�}M�;.2�9�*�ޗ���\Ej���CE���p��3g�_�ű��&�>��0x~0s�tm�ӌ�:Wd�+M��I\^=�]z��=�o5�;V�M��-��C�+`k۞"�ȝ�Ix|�\^�����w��&��ԮW��B��[1�U1�;+̘�����<�
ǽ��ܤ���)����Ѩ����]�Ϻ���w���.�a:�}�#�cf����=,{�^G��z:���k�~�z�~���&��F�u�].��]RH�_��ݒ��uvwL�:�2'�Kۧ���8B�0U���z`__F������é�����p%\�Dd}�79�Ph��z{���*���Cfrqfo�gc�8r���Jj�?�)6L�A��#DP�A]]��s��{���g�v}'��nh8��W;���w�Ax�V�
Ϻ��Nx�_e�СfQ���[{��^�3U��xϪ+�kO��*��G9�E�H��E�EY�ZP���G�ٳ�$gTa�8��Vԣ�������������VԲ�A�l���ULH*Wg���T���p�pe�M�OO�6�N�]�����4�W��a����`z#e��X�	cWQ�U�[��G
΅q����׼��c9���п+Q7.��F�m"�>�I�w��S� �z�H^B�oΗ��J��Az�n{�峹���$}�k�)�ۂǦ��b~�^6#����$�P;�o�vlB��.>�D�][FƗ�ݟD����E�*�΢=��ȈK�VTv=��V�n|ɼ�k|��~�>&�ˎ���Î��F_�d�=>��gK�Q!�^��o\z(ɟ_��,�~��>�;ZL��y\K�x�Qxt������~)���.=�,�Ç�b��@�ԯf�o����H��S�߶�{>�N����	>gNϣ�������ZwS���^�؂2�e��05N�5��`�AN�\�a��md��6L���^���Aw%���e35�J_hW`t�(L�M'�dV0�������"�p�]v�5k!�e��L�Ŵ��w�Ĥ!��ˆw �ܺ�Y��+�u��t�:��6�+}�g�-���ǯG�~�����5�ʸ�Ont���L4sgh<�~�-}�#��M�s_���G��rxef�3ۏ�u��COiq8�tu�yj&/^�ص�;�z�����3o��O��e�om��v�����@��L��7\�\�P�;Q��O�W�z�f��[�X�yd��}3���0���+��d��la�&o�ݍ�����x����^Ʀ��*]��{�q��]�sٔy����(=2�:����NE��3{J����f3���*[oQ�}>�H���+犆�i\��f"Q<b;�*�D��1_\�$k�'FA1����}��﫝��}��^xz��/O�ؗ����5��ĺ1�#��U1S�l���3'��*�oU��QD�N��ס[�tL/yR��ǳ�F5��c��w����A99o�'7w'�w�W-s&T�����Z>��P��1�ש��T�yj�'s�hg�3�gs=��^φ�w�"!x�jj+����-�C�O�����a����rZ�Mծ�#J��UNp�p)������D�時N�~���3�d��6u/1���� �O%+[�	�4ãyV����4��aΣ��u.�j���_;��l�|v��v�7�Gyv�N�:�JT�ޝF�+9�D[=j��%��ź/;�2�ggN��� ��W�s��L"�i� ���1����Ϡ����/Mt^�=�}��<��T!��T�r#sׇ�Nq�6��C�ˈ�s�Y�ٺq��z�:+L�k���ñ71��AZq?-����f��?W��X��G��Χ#��T�K��+I�#�&�5������S��,��Z=���z���ɶz�mzSR\kn��0o�BS���5F{�Y�+����zc~9�Lg�-}��K=�T)��}��3Cr�Dr�W���b��ch?a7�jy�w<��0`G�~���Ѱ����6Kg<�����=y�ZoK���n"5[�����j��7_&D��6Y8嘞�^t�FW�{wkc�N�ٟFx�����
��R�z\F�o��:�z�J����D����わ/��?�XH��+���Y&7M˜��*�z�ɭ/	�H�a9w�!7�x���a�S7}˞����Z���6{���h7�x=�un)� �ˈ˞�q���c��}�g���Y��K>&z˪��g��g���=��^�]��m�	���*�/d�r8��o��n�.ΡQݚ�df�G4>4��k�^�|I�6"z�T]�_��8w����Y�W2���wϙQ������]kLv��8Ź��&+���{��H����=�;���;��DԸ����򾚺E;;�-C{s�F�����7��������>�~���)��w���ʇ�S��;�>}�g�>ȟP�B���<�zω،FGFRt�������h����=���;�\n��)����G�q�o.G����pc�b6!�ߨ�H)WA�KGۃU���T6���>���,<Xݿu���z8�o���mz�8zg�X���P�j�(��8!��|��̶��,y��q��v39oVc�8�#�9ģ�?I��ۗ0�eшЋG�D��Tc �=㱡U_��I����p��֣݇�8�.��ǴL��ʗ�s�9��pM��(��!7A���B��	#�'ܒ�Y!j�G�����%5%�~��σ�ȏ_�X����iA�_GPQ��}W9ެ��m���xM�ד�G���t�O����ѱA+4��Wu��b<�9��F̘�Ρ*�g'Z]�����6��l������ݠ�������f����/эUO�:�~���b4bzuh�%��4}o.�z2f���<n%�v���s��ǜV�`��� j�m�[�{��H\��?����{����(�tU���ۜ�z�P+�Y�;I��V!��:фռY:�:���i݄�S��ћ��d�0/e���۰Z��l���1��J�ks���M�5�N|6M����|L��R��T٘�_���M�?[�h`�:�:����;�/ˆE���[x:U�´����uDg��n{�Sp��̸�Z�F��g`�;��<V%�Q�;�;�����L��t<�3gӯ�i�O�J�'Q�1���6�i�a뗧Py]:�b��ur"�"R9]�Ǽ\1�c!u��ر�^��Y�N/��ld��{�k��_���~;���u�+-FǻE�s�ϯj����X�s����1=5��BSsC�]��J�_c��l*}a����po���^�
�@�e�cѧ޽�Z�z�cެV�K�7����c>|��A���i��u����RIYd�z;���e��wN}��5>�~�;E�lƘ�H
�� �\M��q�wP���7�jbn��^iy����O��l��
���'Me��gĸ�!�
�f�[N��r�W
�=I��Qx|
��ip��tK
���,�}�;�P1�z�ͅ�Aq�֒����fs~XH��������D�<����sL�.��'{O2����?I���|T��UU_��В!&2s�����. �".M�y�gȶ2����o���?v��5���	�" I ��A
(�A���z�^�A<�!D$�$�d$P��P5�V\!��]p�\�B�����ؤ(���Fq|1��;���e�L�sKܱ|�
�}�Pް��p�/���<���ý�����#с���y5��H��&�i�wt�c� ��x ���� ����bV�Y��������W����'�]0�h_C�W�7�IüE������u��F�&@J�h@Y��o�bڤ➲kH;�	��Yk�q��NlF�ܨ����w�b��",cX�v4��4�@	�D�
����tH�qҬ��%0�~k�%�;|�^��y��#�E��-N���F�����I���q��3��2�L�W��]��?���wR/�m�ɯ�!�T�����.��L��?s����b�=�l��GR����y�r-���"*�-@�^�f�Κ��[ǯ��7�NJ(".Ǩ��0���1���T��"�j�w�H�*""Պ<APD_[�w����Pn��T'� ���E�ce""`}CF�m������(��Bԑ�x����tM~��A�+R�?k���b���!&S�Ի
���EŠvo8�؋�7����w��с#c�`�<�~��dj����n�tJr���>L#C������!<�C�mJ|7k/���TPD^���v�F�1�2J����#�EE��[��_4�1�#�yx�M����w�RZ�y��I�����yg^��ݖ![rG�#���0�{��Ю}�uQAz���C��~�g<.,�w^A�= ��A��\��Zw`T.C�*/fA���`_!�j��{|�����@z�q�6���v��5�ep!
�NtyR�,��D�|	�Z��F��rE8P��4�