BZh91AY&SY��ftׄ_�`qg���#�*����b�      �                                    � ;�  �q�              �       (     P%@ P    3�D *E)"D�%"�$E*B"� ����(J��R���EP(�J� �*��
Q) ��$|   �HU*�*!D���@��& ��p��F@j,�0���T=�Jwc�C 8�*�����=x
 �  G��X= >�� q�\ ��== �0 �c���E*� �
���� 9u��'�4 �	  |�"�ETAB�(HM {8>�oa� �`��)���w��Jyox
R�t-���C��� r�����|�Ip mo���=�O� � qO�J<�w� 4�	R���a�}����� ݎ� =��K΀��`���A�{ <�v ^   7� ��T���TUEBE| ��X@;��f [�����u� w��{�����\y�' �9�;��
   �z=8����<��8�� �z���8 ;������R���l8����������{��X   � y�T��J������� �p��}���ͺ ��
��p [=y��y���@/=$�� zoXz r�    �  �|��z��^^=T��� �t� �d ��QN v�9 ��� �w`^ @ O�   |�R�A)AJ �.��=n d��@n���1n U�'ePA�[�Cv 8�UUG (�!��   |   ���n�.J� ��)�1 ��r"W -�@;�r �` �R@  ��)R� �2`�4`O�Ĕ�*C � �	� O�*�Bd�( d�     4�*@�F �&��Fd�	=RQ(B@       �=L����	��1#��12��G�|�����>��}�}�O�A�N�N�0�tT�þ�o�� ]���TV�T�P_��G�P� �� t	�������?��?��:>?��  �A��I$��� �
�'��&�!�"x@EPW��G����D�?1����S?~�m��8�N0�����8�N1�T�8�N0�T���D�
q��`�	�q��b'��xÌD�-��b'	�(q��`'��	���8�M0S��8�0S��� �#� �b�L� x�N1�]0��8�N0�D�1��b���"q�jB)�"q��`���*q���N1��8�t��8�1��8�L`'��"q�ǌT�8�0�P�8���q����x�0C�P�8�N0�D�`'�LN0��8�N0�T�8�M�S�H�0�T�8�N1�A�x�N1�8�b��*q�<b���*q�0��x�0��x�1CL1��x�N0�A� �<b�H@�x�N1�T�8�0�E� xČ�1�Q8��A�Ԅ Cl:b <`�6�Ex�Dx�y!A�A�A� �U�T�*rB*�lQS� 1UN1N0AN1QN0QN0N0QN0EN0PN10NH@U9!E� Q�� A� A� A�����G�^1A1 ^1A1P^HDx�x�x�x� 0�x�D8�N1S�T�8�N1S��8�N0HD�8�0S��8�N0S��8�N1	!�8�N0S��8�N1S�P���ңγc����\��k�N&K8���ـ�H �b.�ý��7C);l��^u�GP5B��ػ���A�ˇ�.<�p���-]I��-�/p�+�u2��[Y*˺��U��ye"��I{Gh�4��^{�����%NL�-�VB/pNp����p}�#�8���N2�RK����t����&�ڣ�I� �fs����1wQ��ȥ�;7{L��ۡ^C$$�>P����Ic�� �Rr��rZ���z����m��j�c �?\�[}d�hG;�Զh�{.�õ�7^�8Vm-K����E�:�8pGwr=�cʖ����/	�^�pM�'�W��{���"���d�KB�/ w^��0�� ���ŋh�݆e�ĭ:+pb���OsP�q�b	�0-��Ъbvj������pnҾC��\+��ՏU�N0���Ǆ��8ֹ�9����#vnP�b�q�Ď����Y��-
�u�q�T�7:�l��u�-[��ia<Y=0}��r���^l��Ӹ��)���s%,QL=r��}��o�s����S��-ז�����,s! ���H�<dَ��np_f�=���7 �ā���s�	��9z����q�������H�޺ ��}��]�.�^淣�>�r��'f��ڊ@f�˄tGw��2B.A��ţ,qS_�~@�����tqoL�g$�j.m�mA@����!Kb�$��m��=Y����on�(MXu=c��î�1Z9����\�6��X5p;����ǔohbe$#�3���2��l�{;X�跢�������c�SNM�]o����Qڱ�F�;��:'f�0�Ye�S
EG9��@r>8t=��i�d}�J��su72Y~��'&U��=�ծh��c;
�٪����߉�˦ H�0�%l+o.Õ;��>��1��Vţ����¹`,j�m+�@W��.����p�wLE�
ڛ��M�d��w� @��'\�͝Uz���[��r��M:&��u��y�R�Rʩ��K�9݀8�lqg�\�Q�\O��ql�LK����� �-:rmC�V�k�g��O�فb��3��ctv�=�w����{h�-Vw{C(eՀ���o&�n�C=�M�m�X,c�i4���t�$��"�{_Fj�oT�(��M-�qm��3E��H�r�ԘDК�=�G�r�T��n1�w�d�g���ΐr[޸W`��;N�:��A]��А�r3!|�Dd�����`�ns�o��Hbs㏘;}�rW	X�p`�&څ��:tu�voqٖ��s�z����j��:z�xW�F��|@��є^���,�~�z�^�m`��i.w5�r�@`P���DktRHg&`��ǁv)��y�Ǣ��T`9	�X(��yScuN�8��Ǌ�|�G#��.��3�Я
j��ܤK���B}�͝��#)�����&��g��,QC��=]A���q��.��Nr�8X��9�s��52���RR)�{5��W�<�6u�&Ǻr'�wWo>�nHY����Zu�Wd�7��	�z�u�QQ���${	�\3���@.\ܓ�D6�R��Ɨk���̫��C�et��f�-> X;���V��k�xsQ��'hS{oeĶ5.Qdǝ���<�K�bkT��o�p����f��;��Rk]��7wz�NnA�0�룧�X��p�5ԃq܌�z���Z�r�n�X:�&�wS�N3D
t�2��e��чp�Qϋؠh�r`�����%��]i���ġ6^U	Om׼�M`��nɹ:��Ba�/Z%%�����S�r�fY�vo.i�ˑշ�h�����8%Cvl�&��H`�M�ٽ�:X^؋�m��M<2�:2�Y�a�:�E�_����KF�.p����|���iK�����jc����|�K7F�^"x�[�^7��oa�VX�G[q)�I8%[�-ʦ�o��Z{�8CS��İh0͚���8:�)�l��Ƈ�Nuܼ� vN�v�N;�kw{F)۽���>�q<��W*�ى�V��ܘ�#���,u`�V�V�\��,�9�ġ�u�]�<�X�7��q�=���{F]:Cd�麌{���w�gwgs�a�V��(��:�����f\r��'i�wsL�{oAw{u��oqQ���K���Fn�t��a�Fv%�f2	1p��=Xu�:a�,�=E�a�Ch�N�OQ��鱡��߮٪-0[��5��ġ{kK���ڐH�
�G٧x��݈o!̈�L[��Nk�ci�a�q��99A!���]N���%ٯ���[����fq�/�G�$7�1G.R�I-#�xs���d"�w2S�R'n���v�jD3� YT��WxnT*)c���G>��q�NC؆�K�qL�U���}�(]�ϟ-|;NCܺ��n#FLܚ.���1�D�&چ�F��v
�ڻ�m�[����2�=&pJeY��S+��놕4ge�{0�Y�m=Yx���5Dl��M�U��vm���˶��� =˱����n�w�w5�ݑPb���z77��d�e�{qy��.ާxh�W�	����Y�k�uI
Ao۽O�)6�Og=�aswN�I�֚�,�\�N��4�DW�l8;�.��ذE%�,�u�B�>·L5#�x��:���6�ݧV_c���2>��]W�����5]WH��l�~!^��m�H֝�.�p��:���νǰ�ߣv��Ҭ"r�^쯶$)����pӨ�{�Ŋ>s	��ؕ���&tG�6�ƨ}l;�w:��=L�cn���ֽ����}�_��{�T�m���������_^}�Lt�3S�L�^�&�d��O�%\�ɇڞ\���[|�;N��ܦc�yg7�,���L���M�����I���ܶ_n���g����I$��nl��Ú:_�wN���Eۀ�����qʫ��%s�u��Z����o]�ܺwf��ND�-�SN�މ��4gVuh���P�u})�q�-�ռ#9�{j�Gdٽ�N���䖄!�׀����	��;F��:�ӺW�K%�i� �����Mː��i�t�˳����\��s��>���?u�7x�������x�E�6����\fvf-=T/��,��⥺wn���zl�	�6b���D8q�v�\H��ך�������Q�-�,�uV9A���d�A�ypS
��F2��m4iɎ^:�^S����p�f���MV�����{}��
Gn��j�%93u����ak�l�<���v6�浣~��M��ܚy,J�9�;8�fYR��nø^H}�[}�ŝ�NF�@�ʹH���2~/��E��̹�8w]yέ���]���Sǫ9��-�C,+-���8TI�*�7�>� ��;]���͙��{���w�ns#cK��h[�k�QgN�7��w����+ Ӝ�뗦�5����C� �4�u�7�N��*��S�UvZқ(rxPk��G�j��<�Gsr�{B�LX�3p���n�`�=W'o>ZXV��K�YOk�;q�l$]#ճ�-�8�]���{&?j�^
���WC,���&ֆ7��H��tu�����z<c��>�x5s���ݙ�9��↮�n&3�:�f��=�o*��-8u��[ʰYD΅ii��n��!�����D�7GM��0f��KI��4�7��{�eL��Ꝓ}hs�{5����pg^�(s�]��omŢ$�Z�j�����qw�x]9����ᦱ�t�ءmn9��u�*0���7���N8�#��np�j���C��E(x|b҂��e��X�݆�W1�f�E�5P�!ᯩ܍6�&!3PQ�hE���=ż�Q�d�tJ:k��r�Z�r�;��m�c�V�K��w�S�c�O8���^�s's�nrp��9��*��2�x�ӼE�6ܪ�%�̃������j8}��Biy-�_0K���5��"���k����bCt=��qV]�t�*W5#�ٳ"HH]G`/Rŝ�C�ޣ{���-�)���惸\��"M��Y�J2h�8��
�va5mZD5�^MLG���=ٴ흶�׷ѹs��y����,�y�;�}C���W!�!�)��z���7�;����� 3���Z�������vNzK�54BO�����x��
� �Z��.H���nK����b��$oG���.�s�u�2FEܰV��8��^� H�*(�q,���r\��i�$$FV�x��^�W��ù�#'z �՜+�cN��wDq�eĲ��sۚM;�1�����$*	p���g#��h�T�8�[�0����/��5[r���Y���W׽��}09�#�a뭚��J��2��%�˥�w������0,���w����eŧK$tUeCq5�P�bV�3�V�-j�Aɱ�\��륎S�[��hki�f��9j�W���0�}'��~��yâ����#�л䧎��g��`�8��P	��Q:s�_h��j݂f�v�7�ðE"ݲe��R�`�K�����.���\

m<(�	�wI�Wp��5o�=}(�W�sju�=�n�\�ݙ�oK�DFl�H�g^��2ԝ�]U=/F���G��Bc�y�P����Ӄ�ْ�Y79 �G���:F�j��B�]c�v� �!���}�88�E<�eM1��F���Ggp�n��Aj�4;8"Z�5�[�ݽ�����'��_=8WT�����(8I3&u.�㓲n�=��_۶B3� .���g^�UE�{��n-������1���Y�wBMdq��a�GW��O�g2�:����K����s���>Kn�H�i@5F����ћ�q�oR�R\����p��v�geUk�(}̳	�v�f+_c���t|~��d�����~ٝ�Z��9vri{�ةˮ��pgM��l�B�ة���bK�G1�g`'�]z�:n�ubt�c�nw"	������gmc�ÝP�];%;94T(V[oj�&�'��EQ���r�t��^��Q�J�q�7'j��]罷->\4"S�R��wn��7��������T����7H<� �m��AG����
8��3�Z&o�<�h���,�V�G�ra	Zpk0��	����WW�6��3^��B/$�]�� ���������PJ��3��֏�o^ష�_>K!���s�n-q��:U������~u�a
�U�V�!�t�Nv�"@D���ỎN�0��x�Z�p�)���\Eѽȝp&�[�����4!��/��vLAk��� ��q,��Ʃ����v�-iñQ����;�d�9��of��P*�L�|5�4�1�b���z'@9Vo!�KܕtIs�׈ϩ��M�u��)}+���F�y;�Y^�-\����:ۘqȷj{�A���x���wvc�w\���[�6>�R�ۇ)�2	�_@��ea�G̸i+##�t]� b����r��v���e�ױ,і���K�a�AS�Ţ]Z�`��@��kq�oA������ѡ����r���[#[3�rD����Q�$��.{��B;�,ֳ��{Q�e�b9VI[�Z�M����A���sRA�Gt�u����=�Ѻ��L�7 N�9B�n9ʬg ��,�`Ж,@��f��� ������J��.�M[fX�[��<�L:������T��i"���v����q����ڱk3�y���2Nr����'S�{z�pgx�>��U��¦)�.��!�ڦ�M9��b�N�SuY�a|�o�[�x_i.��.!-�"�-w��o1�����V9���݆�sd:�G;��ջ�'ڬ']�G,���^��״��vlJhH��a����3{RvvK�wP�� ���n����x��G��1�{�m7B͂i��Ʃ����(כv��}�N�� 1�ڪ�����d	�0���n+��;AӃh"�N&
[�d7uw0��09��E@�.bLv��q� #w�8!���Y�Jc$�p�e�S�I;�{��X��s�ĸ��m#npE�9-��@{���̆A����p�:vL.Gsqn�Ͳ����׫�m���>��C���d��Jt�A,�n���=t�';>�[��Y���hr�\8�O�={Z�s��1�Q�G>7	�������d��9>��T���Y��-�\d{xp����d3y�{ϟa�R���u�G����w�P����3��;��H��s�v,3�2�Ū��rnk�2��̱Ȁ�r���oA�:��n��ԓ��,�� �دR��K�wo.�݁vhgQٰ0w;���d��Y�z�^z��:��l=��׉�v<�d��gK����i޶͜�)?A�I$�t�N	D2�>f�<M$�;�[$��go��ߗ����/���m;��	����l���l�`�� �����/�_����%�>�h��!}�&�7I�Y0��n� ����e�����>_�pӺL'���^�u2!{j���(o��J�<K%�$��T'�vɇ����ɉ�Qg����dx��0i+ $�8�:J���wĢt��=�wI�Q0�O��|N���1+��B^-��F�O��|J:»aOаM"�6d<N�BI$�N���N��Ӵ7�Id�|d;����'I��Y��pFA/����Rga>$��Λ�z�u�|l:��),�K$�a:Jf�id쁈h�`M4���
����T^�}ߠ��j���'A��>:Q����Qjحj��EZ���UkF�bִm�QU�Z�j�[k����F�m�cmm����XՍZ�kU�j�V�6ڢ�V+l[E[��V6ֱ�X��Z�m����֋mU�b��U�U�Ţ��X�QU�5��F��j�V��h�U���*�*�V�-j�mm�Z�Zص�Z��[m�X���mcV*�cU�V-kXյF��j-�j�Z�j�6�mb��+j5�ѭlmm�Ѷ�V6�lj��UX�ZEY�BA �ObT]@*d�*���RG#����|��JP�D��A^��:"TN�]��/�33I��)�u�G�9�A5 u��^�E.�@r��*&]�Ts��= E��������������`���L>e���"�?�������W����>l����	�t�K}�fw�?yŻ��"y�}��>�ag$�I�-�9൝4k[ڼ� ��%�Yʷ���]�����ٚ|;" ���,��T3�"n�Q��t��ǯA�n�g�\���9���*�|�蚒����n�[�����(	�_M�V�K�4��eӖ������������ȏlȷѡt���D�
��:/n]|�x��dJ͡	�V�ӌQ����׻;�|�ޮ�>S����O�W�v�w���qD�}���酛�}14uM���!6����6�j훲=��Gs��=��2;�M�\U	����l{��為�G�������qϚ0N�{�� ��6[9��s]��E#��p�p㻥-�_m����,��|;�Bk���P��e#�#��;Қ������<� ���&4z�k}���{�V
<V>sJ�����S���dC,C�Б籣�\������d���ogP}���XS�	���;��}O���/t����K6#���x�����n��Ԯ��ؼ��w��t3׵����t�Y�Wc������y@d>�o��;q��{�˜ek���������<�� 6��w^�	ͱ�T�<���4悇���tݞY53�7E֓&��ǔ���'wA��#'C�j�I3پ�`b���͉�M�O_xSW�������|#8�˺��4��L���&=�L��Bl��v��Q�����v�2���F|;�5��ۓqb"�&A1�����䶌�a���U(��uc�g��ga(
w2��٪�r��?K'�M�Q��||1x�\���T�	�0s|�^����W���7|�?G�w`�/S�z�����Id�`<�|r$�E����������<l(ۯ���åA}A��;���?�/�*�WU��6����\����q!o��/�5��}L� ^�X���o�..��ʖ��ú�r����s�����_���=:
ʊ��%� $�r7.vZ�7N�X���~����^�ˑN8��"��ݓ��Ѣ�G�g�g�wv�Lx7�W���>�v.���9���u�R�lQ��]�b����ͷ�4]�C�Փͷ���\�pw�)D�hvj��l�H:~Ĝ�-Y�s���f=�F�5���X����m}������1��xx-`�Vù��w}8���w���]���ȍ߭��*UA��1�6n������no�����=�`��v���=.��ɗ`B%��!�ߩ�]�9�����Of���ӏ�&,V��XD������;͞�z�ٞ9c9��^�G�˯��u�л�sU]]�kO���/_b����qgZ��$xc�0v4�v�5*9Ɨ�I�rx��GV�^�Û��^��}�K�:z��ϧr?x#y���Ǝ�I;���y�ۮ� �=��܃�<���\Z;,�e8���h�4���wp����4iDJC���k뻡3=;o���j���u��B)��=�<[��/��u��5AW��ۀ��	��8�DM���i�5���y緆�{�i\��jX<����`rY��>�g��o���u�����4�A��.9�gp�Z�S���̗���Y�1z���i�:74%�×'�Jj�">����<��.ݴ���8K]�*y���s����|�7�o������^�H��
�Է�{�6��(��GB�k��Y`�^��$P�n嚍[��9k��{E�%6���Y�geɉ*�VQF��<�.9�{�W�i�gb�4�z����G�a'�6�:�t{��=�h0V�yDd��]D�L��V�.�T��=��Iy٣.��?%_�0{��˒�l�.|�G�Y�wm�U���89�7f}ڻ�c�r�t�Y�o��<w ��i彫��,�;�d��0�/<�}S}�/Ytg���r,[��W�/Z��{�����Vߵ�q��[��a���7�ɼ�I7ۍ��f��7�j{֙�G�%�8xi���ay�b*�����l:L��ǃ{ڴ����=�S��e8���'�(�C����1Ƒ�<D{�]:�j�r�#��� ��I������dž�f�yx���҅����c4{;i��ؓ�*{�w`�^��b��y�7�\v{&��bG�r���+�5A+���i��&���7q9�����>��h�3M�꒾�ON�3�:��|�{<^ȭä��[��!������n�",E�;��P#C��#ۘ3;%�,e.]�"v.�ܼ�LZy�����G%o�&�}Ǘ նjyN����ױ��M��x�Z.��$�p�nL��!�vDN�UܑOe�y-�!��;_�@}�rx`�$��Z���{K\=k�t��7��['�uc�����,��:n���NxQʯ��j�7q�[��3��V�6T_�$�{�3���޽����W�1�1!�Ђ}��;{<��qvF�x;��:���A���vN�=�5�7�ug]3�g�y��$�65��>��@�-~��Ho������j9���q�ңਥk���
pA�enh�=(��Ǣ�E�TA�����z�!�3��Ṡ{�����T�зt`]�׸,��G�^�|�C���]��W��,�m53�{{����h�}Fڲ
��{S%;�t>Z̬bNfd6X�(��]TM�-WD��8���0�����*���=��O�K��Z�V�#�j�l�ȫ�.��v���z��3-T�V���d�Dľ)+�gB�`;ۀg<����=�3��ȕ���n6|��׃;�c8;~:茭L:n�l�ճ�ͭ��|+~?o��޲Y�}���u���1�r�����:�gx�{��+�ۤk�A�:w��l1mPz�v�UϪ���ڮ��y�M���n��Tp1D>�jڦ�<��~Lg������UxS�w<�s��֫pW�i]��[F��8wY}!�OBQ�}��^y��&?>��$�k��>wc��'���n���^F��)�=����{���=����5�M��x��/9����4f��CPd]�x�_�����ؤ{Δ�8�<3��Oǳ��Hk�!G<)�G����9�_�ܛ��/?{]>߇���>��!�G�LƄ��}����c+q��K�恮-����邉E-)�ݹ���Bu���g��W���3�F2�{>)����>�i�ӆ�O����p��\�]5t�)F���8�?�z����!��e��5O�>�zYe�Nj�dwm఑���ҵb����x�i[�^y��yT�\���-��_eڗ�����3�{�sI��ޒ�����D�X�-]��w��wlr�W\�}l��I}�΅�������{{�����q
4^��H\P�2�s��װy��5�X%��K<"'�6=� "�j����V�g�T�e�%��$�^�����gM�*<[�#|ow�RԾ�")�$}���g�;���T>�,���ѵ;�*����A��ףڮ���s۾���OxC�����ᕤ�$rAKva��n�/h��{<ؓ'�~���=NrdF7�S��J4x璘�z�cs�HA[�B�E��yEH97��ۻ���q:�������~��|CA�z�YwR��Ƃ.o���V�g��{ӔɥM��H��&�����1��޼8��u�����N�����2?�U�/����xyi�{�,�T����o��w��oHv���p*o�r�|�O��ql�%�,~��v)��;W��A����9{���)�=.���'�fj�m�,�k��H���^�b�|T��/A~�3S^��HHO�XS�׉��J]{���Y�ٝ�w��m�ANF�?|��z8Ҡ@{=�A�����w��h;]���9�<�k����w�2��s��}���)ꦧ_y�p���z��?e�1�-�^��Y���������G�ٞw��<kӘ���ش԰���>���/��-���4��|���y�����>�2��儜�ˤ�>[�ݲ�.A��h�w�Ń�Ko/v�j�@�~m�j��G�PT�h�i'��=7������1i�e<<ƍn>��Om;n�ל�D篦��J��j^g[����i�9�^�<�/"!��	�:Oe���71���,܍���:C)�=��}{����ax�̙�X�t�➢���w0�P^΢���Px������<3��o(��ˆaM�D�ݼI�E�Yb%|��:^#��uu�%�vL�2�+�� ��[����]����X4��s��>>���'y` IM�\�k>��og���U�3L���|�t�`2Ww}o�s@9����f�A�G�i=A��)X�8,����o䅆�1l��<�B����1�˧����9�^b��*;��C]�;�֬qN${��S�������� ^X�/<ף�g<���G�#��0ڜa'xa�b��Yj�e�u}�P~^�/���N�7;���|�\����Ҟ=r?`��x��(te�x5N-��Ki��,��<�Ѿ��Ҋǥ.yPg�#�&��b�S��?O�2���2d�잋�$�=�����2�s�1�:�=g!D�[Ÿk��6vt��pL��m�۳��=�/LA�dx{�'�YɒaY�#����~�W|f��,��2rP��箒�Ú��E^�zɕ��� {��B�y��8G�ۖ����v{u��^<:.n���"<܂���,]���FhY� �[�{�x|�[����=U\����ds׺S˺���kƒ²d2��}v��4wP�0yu��}8�jJ�~ݞ�}�Wa$��G��rK��{�[5�w�nv޷��y������ܣ-=����Ƴ�/��HG�������u�`�<^?Xng-�QW�L�`^�d�ě���.C �s}�0؈�����.�x�ny=�O֎��:+��� ��KԚLܘЍ������A�x����#���1��<>kmL����;:y<��7T�"4M�Pi�|�yp��#��B^X����N��y�&Wa����g�";�o��'���6�{����..vIU��F����R�yPpr�9׫�K�z�h��y?{ɐ5� b��u8��>�'˚�������W���&ю�Ly��7��ֺ}�(�g1�+��V�KhY�7�ܠ��{��؇���Ө��r|��!�1��5�tYt����F���3e6�y0������8�iKMw��ɞS��g�@�Y�טfr����\|N����>#sT����ԥ�x��ok;�B�����{hk�^�1$?&Z�5��@��)���f��aF��\cg,���}��>�I!S�$�{�j��܆n�E�<�')������X��X�0Ae�\H�m�B���X,�[.�cXgb��N���}[ܫ_���pH�`hq��^�^5XNHl�j o��U�	�&�*���s��	�،�I��Z�Q&ѐzx��v�>���Z��}��@M?��6�82�ӳC�=Q.�"�NY��d�M�Sݽ~�r"�������=�}���lW�s:'�w���~o�/ws�;�9�ۈ��l~�}�=�����������M�[�s��Y��r�1�]�<C\�܈�v�_9�u���z�F���`��bd�v�lK��ϟf���Ý��l�_n�[5��%�8ǘ�7�i2����,�v�x���柷rxd�]8)n�rp_`�����
	K�X�r]��e�jo���C���������q�#��rj:UCT�{��^�ȜK2��L)j1��͌.d+�? 2�9��v��&;�[�`�'S�t����ߺ��Ov_f�^�5n�?!�8��=�;�؏�dȶ{7��z�R�z)!a>
Y��o�i���A�<��2�����D�g��=훥�Z��ZV��~m@�C#�'+���u�:��q�q�	E�C?�ϟy�6��=�"E3'��uS�;��xQ�۬WK_==wә�Nc!uZ�N�N�I���q��K|3Tˠ,$����X��r��+�z��S|��E�{�OG1jYG`#0b�K�s*G8i�}7,"���<ާ���3�3�W#���fh<x�Pe�d�fy��^{�`�)�,i����9� Z��b" �O��ȫ$�+�4�G��{7&٩����[�	nq�1��;	��h����}��j�b�@���ʿ��;�uo�)Q�X=�O+���yvӗ��0�ֳk��_{�UQ��� '܎Z�33~^�?qė�RXYS�v�l�Ȝ����o����zQ�}�洁jR�%��'�7[$�j`��x�q����6��W9��Ĝ#e�쫟��ݙW�gO%�����<� n�9����d���[t��M�.��'fU��d��{z�U��c�/n,=|;��AiZ�9�uw�qhilw�B��
d[V��?d�@��t������=�no4h�bG9/p��٬a�=	z�lK���{����%w�a|�'��ekj�{k,g�܇=�~��U=rOiŤ��73�lAt�6��~k��s���ٙ����N�[�h`����m�|pse�{�.�bk���U���}��<�{U�҇w�'�h��u�����\O�Ź����@�՝�s�m�-{׵�+�=I����,��x���eMk��A&Ǜ�dY�	�N�"��=�x�||t�!F�<�%�>�3Q�椯�{/mE��ӸiE�!ѷ���/er{���;�����|-Y�W�c
���{���~�t���3LX= a{uw��%}�^�� U����~����?_�_�U�G��o���������v;v�۷oOOOOONݿ�	��K_s�ߍ�&�9�%6����i��7h[Z�b��8UNb�6
o��f�k)_ًl��Ŗ�t�=���|��X�U�fq���q���WM0f3�{����U��Y�b�`���CAn+Y�aޠܥ��ѻ[n%�qC˱�@D�aWn��r�d:'V0�;�n��v�xKh��.�n��a�[�N8�qL�f�G�뷷�/Y�qDѵ�m�������w<E��s8q��Ӟ�M4�4��]���9u���.��n�v�v]�n�Mn�(]\y��n1����P{F�eM��n�َ�l����$:�Hh�Ÿ0t���l�ra̚����RbbX�*Qy�H�X�k*�\P��\���[Y�,�N�u�:ʇW�ZM���v��!�-�9V�z脫F�lZ�!�5U.���3f�LJ��=%�D�:n��(s�D�]�z1�guQ�@ȣ&��@�e��K �#Zb̺kW�`����9-�����o1\vY�:ɹ;d�v�G�c�atSl��Ql�Yl����],�M,Jl�1+�PɃz!j˳�-�k+��;��u��<x�����On��mۜpcSF1vN[Q�����������F�d�V���Ĕ��h��b��d�vwH/,Ǭ��&\U�*��x ���[]v���2��#�j���R����� NFҚme� �ivԷ9v4���*hv��ۻ1�]B�c�Օ��`���l�5�ɲ���(�m�ۮ��]!����X�Ki�,��F�E.%�]m����:���0��\��G5�3�ō�on��]��w[ф�v�˺��E�7J�4b�V����J�wE6�]��mF�Li1B^Ŗ��;�k�ѹ���U��P�I��0�!hɴи�se$�+-�@�ls�%{,�y���۞%�q#�Z'=8玙�k+�g��ﴉ���w�� ����۔^�:�V�Ү��RRUT�q7�f颎�7'eͮ��*�s���<��j�x��eG���|����ɱ�<�؜E��V�\a!eq��Gj�*�a1�Q� jI��w�sl��d�K��q�v�"��p]n !ߖ�ݠﺹv��>+v�>9̓�9���|�L	���.D�iXRLF8�[r�5�#x�Fr<�f��
_2��N��D��%m^K��ul�Z�kE�ڌw`��b����2�G��Q!.Um�B�:7��oh��۷��=1�x��;�8�u�n7]�Uɶm���1 ����[���SN��*�Sۈ�sv�v��Y�+���[*[���j�B:W�D�HẎ׷`�I�]��]S2i�nF�0��	2�q4�MnK�F�+FC'���7J]m��=ru��mƪu�	�F���$:��ϖ���Y�E�T�`���WK6���5[��PŲ�i��ٱӨ5��x�1;�����b6,�ᦍ�Z⛮��MnɇX�z��Bԍ�ť�bk��$�M[�XX /b�GhRSD�c0��G�<��yb�96q]�,v��Y�ݶ�������v�k���Ҟ�k�n<�v�)9D�o���wjS�{U4�홁�x�<��:���B��If.�1�V��Y\l�+#1��%�z˰�vf�	";Z�p����GX��8qϢ0Gn�y��[FNB��Zg�ixj�sΗZ ��4r��/[�#t͍4�ގc��Su�kLU������R���� |�%����:P6\ib�ns̽����gۅN[�7eZ�RWbXX�@�90��ŸJ�a\�-�9J[�	��dS���6�ŕ�T�˱Vm��τ�uI�L��>���C��-�;F�� �͑�M&#��.sv�'v	c$S��-�SZ�t62j.�Sv¬,K�qa���Gx�ni�7"	u��^��nx��Gq�v�f�	��]�V`����,���/�^^-�,���]�Ǉ9NI��i�vf�ꞃ��$n9�ݫ�eY�ش���]���B���tc�MN����&����Ft=�;N�' :̏m�ˬf���A#�B,�,XY��ϔ{q�'�[��0rҝը�<\m�A���I�ۮr=�Y:�I�'��FX7b$���^&2d��������b ��3L���4�.:�}r]���nm����UE0����f�m�-u�����q�\W����m�a�������X�+�srt��u��s�n7�V���g���ݩs;t���sfn���I���6J�b�	�6�6�h�5����u�.w/]q���C�H�t����0�`�F:�3K=�%��&�����GL�X]5�@��4�h��hK@�1��8Vf�Y��x'�d�+2丱��IY��u;�b&���`�ּ5�P�h��b��Fm�e%��f-"��F`�$ݣ�&�tQ���H/7.�7`�t\���\7os<�MM�����k��YU������6Y��Y���#��=<vշ6�]����`B�sY��A`5ӡ�m�(�a��9����[V�-��>�<�5۔f�]e����� �+
%	F,GS���{$č�s��5���k'��0�x�n.4Ȯ�]��y��r������z���uЕ�#2G��x��FLj�;M[�ZA��M,˚�f���c�n{p֔�%WQ#�΃hc"ʹ̚ljMXú�j.p��b8��p�$�G��b�eM��I�B��^Ӎ�1 �m�M�vsfefc5�oJP#
ZN�Fӭ�.�;�xq���v�u�F뇮�����8��>�=��n�$��f�n7�aר۴�+.*�,&�;m	]�MkLF���7V{-.�p��l�x�n�XJ��5��C0)mih�N�Ugη���p��ۈ�F#��������R�Ƌ������.1�7R�˼���=5�-]�WY1i��ʋv�x��vl�]Έ70mc0��2�)�$�q1
XX+��n+t��&������{�;����.�R��lx��3��GB�qv뀗w`�.�84��׷�˂b�Z2��f��0#B�[v.e�mz��;Sc(sq�����'�U�h.kc]�=G�v{t���3%�3�aʝA�:�N�i�)�<ĵ��lh^��o]�=��\q�@�y5��'�uݯD���U��8����W�	o��>O/�ؚ��:WLD����
�ۛ��z�kE�[��uÄ�ۭUq����K�su�63�έ��s�ăgr�q����}�=�St���(���ȰFR�l��C�9.	��<�{v����ۂ�اa����]N���w<���q���)iE&.�fq���ڪ��Fc�����4��܏ Ӵ\C�^Fa�ne��R�8���wY$�.��*���wl]���S����ڋ(��rs�E�T�x�L���,ьr��,v��F|/Y�&G�6;F�ݶ���z�2r�f:��RJ��7�#u�&���}i��<ϭ��h���wOylQ�K���â���v��Ǒ<+X�f���e���b��`�@��x���6m�.Inn77by����E�l`�Ѣ&�6�CE�)�W�SFмX�sKWm��X薹}1��jr��	��f��l4�b!�h�հ�a鴵�/N�Tsy���ώ�q:cR)m4ū�������37Q����z�cA�\�^�@�(�w#��2ۮ�����mp ޸�y!�]m!P���9Yf�`�l�9�g]�=�j�N�ƣcE<ٲ]u'=�:K/�_��|�{'�����xi����Ϙga���M�n�-��t��"񠵇]�=�������"\r�)r�Z�������윷k�o����d�q��u���=kd��Se#6�f`�:ȯh�rC�������L��hhk��xּ�]�.*hB��*8t�u�Q�o.T�*mkt!Z`����L��9�9�n�y��'%o����	d�t�HE��:�&�*0@4mՀ5�k���B=\��;k�A�&�:+t�bRY�������`�D�tA�n:�l��e��f�5�e.M���s�xqn�z64��UR;<��xSv�mxHR��9t)��&30
҃��mZ۵j�k"]qrM-��,^�A���l��dxl��Gb�Ď�1�CK��LAP[i���eV�rX��BnbҗN�]����=m�1�çס��v;��ELx�M�\�U��3����t���Z*�@���snp<T]GH�t�t<1I��{3ۣ9� X��@��K����cZ�5���c��ĬVā��01r�� �w,/n�*W�*�^�����솭�ķ�׬��N���44������q�m(�%��^���_o�w?FI�`�6���6�nӘqq��I�cq�\h8�78պ�้U**d�e���Ŭ�U�bu�<��yM��#����!v���K
��m'n��b
e6��b[��E�f�W�:Uk	M�谭Ҋ���	��\Xrm�pUy8�F෵P�UC��e�5�b7C�4����S���:t���[Jމ랸�;�Re�,\���<\�&�nɵѱ�C֐�;vX��b�nr�OQ�U��.�\Im��\�t�W�TF��!֦�. �6J��`l�e`ͺQP�F�v��,�x��6�����n�dê����v�m���0荫����n�h=��;:�"c \�lo!u;���=ft:%eB2`�YV����M�>7\\�`���om`�R�Qy���٫���\��=W�-��	p��7k�uS��{j�n:`��՚�6�3[5UU�P��˚�7��UUMSUUUU*�UUUGlݗW=�妪��ߺ�����Rߗ����H;�0�]�v�OX3sq�[L���u�����G�WJg�4z�1�օK����;s�5�-�rm�����*�`��U��I�O�|m�;���=��r���е��t4�Sć�3c��<l��jb�m2˙LCtB�<�ob���i/Z3)/�\2{���Dn\C4��]��\��$)&(l�.W,�;�♘wE�퀏��𥳐L�����	E0)b�*��62���v�F"�&c��u]wk�K�r�^�����&e1s�$L�v�+���H3Pd��(����G��L<�1�u�s])Ifwv(�,o��%�*/����0��|�ռ"O.���EGι1R\�f�Q��6�lbJMsr(����=ڻ�\�ce+��s]ݸX�s���^�Tl%��]����y!��#���*��W5��q�C3b���r��.�˛o7<��l�O׷�t'��31�KF}�5y�*+>;��2&Ő�P�+���^������	�pX-�h�v=��Uzs����72ض)(�aFiP�0�-��l�2ڂ�mp�=K�����|��F!F�ԣ
76+qvqt��������VP�!R�l⣭���ñ��\u��OY�f`�u�\k��W�3�l�v5�]����<�M�6-�<gm��>�1L�(�һEچb[4 M5t�끊�ͼ����eX�X�k�������ɬ
0��5˶n#���"��n��x��/hڴ<qUOv���E��]f��I�R�k��;7K!i�۟S��+<׭�!n�
�%���5���y�-�v�+�u�l��b�l�3v֛˴k���:�n�Іv�
sv\�<jk�n�5��Ռ���ں������LB�^cqR�\Q���+�;��Z�ێ�'-��n��>k��=6d���BX)���]�B�GV������f�'�(%���7-��08�����%�Q�m����8�R"��&ғ��c��v�f�F"Q\!���R5L�S�X�g�:��q`;1�ۊ�.|p��#]v{U�3��Xz����������<�fYpb�
ٔ��Y�� X�^�`�<m�����;��-��i��3��Nˋ���vݤ�s�k�u��xh��hb]i�s���,�3X3:�z�u�kMD%���u�mB�7*2gq0�un0[�:��u��l��v�jrV�(\ç�)�ܻ�m� �������)5֜�]4%/]���Jv����u�r�k�Un]��q]����,'��\�W�J˰�)��٫� �	��|��XY�d���rx����W�k�:4�����t^���1;p t�f��k�TIf���2�#:�p[���(½t��+gF���b�%Ͱa�,�a�6�k<��۳�R�����]V���܇�Yj��O���-��5T�4Ԫe�-���.�ĤA�<�m�nx�L�D	CGWq)l�Zi����>z魛�,IX<F��-���Ԋ��c@U�-Ql" Ԍx�RڔZF�m�԰�9X��I[,D��XӋ+H���YJ�J� u�Um���	eeh����R�Ҳ�ƌ��Qj^`�F�
��A-R�`��H�o)����Ae���͵
%���=K��?z�آ@r��B5[s4 ���M�B��g;�4Ks�f0��3@���� �% 7�I�{�¦"�"ҵ�)���W�,���k�-��Ֆ���VC���;��]���{���%�Ɗ�vK&�|�z�6��.�a���W�Z�M��I�d��	��q,.�.!���n�{����K�۹I��x�[��h��>���Lf^躥[�k-�h6�BoNT�K*r���%�������ʽ{͖詺ˌЦ��\��4^7�����jط��l��a����v�s���e�hD�EEԉpL��d� e��)O�#1�*�I �CT�x7�;<u�Y���կ��(fۀ��d������Z�02u��������·u]�^G�t�^�Yv�8f�x/A׊"ybw��덴x�7*�zT����Gh9��$>�3�2f�������-�e�-�ͽ�y+��վ��}�P3�m�No$&�<M��l#6���++iE�N�.P�r��x���&����Uu�K��[ $���S�lã60��7[Pފ������=�������e�|>߫�Ja��F�)��� �ne��[gA���ž���d���i�ke��1���xg8�&�+�5�5��-�3��#��œP�n��N����IB1��J|�xM9W��!5:�RTf���6���9x����P�6�UL�U陜��m���E�>n�>�x�F�_z�]��ﶵ|��/)���?Zrʳ-�?��;7�������h�:ۓ��O7�^ʷˆ��2_N�+�6T/&0�I���W����ۉ^�/�7��hJ	̫�n���UҲӘ��l����}r�׍䚼S'I���CmS���ZL�zh��̍�隖Z��4�7zD5�L���d�$�Г(|ͷ��'�;�-n/��t�lag�7[�R޺�I���������qL��YO��$Q��Z �."��4yl�88�e�ڦ�T>z�߼;�I?�`k+7\��ђ�9{-v�-����.�������I�`�8!I�.ג�ɤnj�#t:fK*ݔf�^6�y%Z���+�3����*�o%!&�n[U��ɷ��n��jS\�ag�2,�[�X|�0	6z���bz�����Lϟm��^m�6�7�fN^�J�7��	uS��;�M((0��󅁠�����3F>��d�����/AK��ڥHQv4��{^>����(��.��%Z�S��5�fj�����o%�5:��a6jj��4:fK*ݔf�/?��$���CnT����l�x�g�!�]��ź�#��ZB�5�A�F�Yef���e�?}��y&I�N�p<��z����n�����l��t�@��j�n2I)	8���1=��������71�C�Eފ���`��<T*۝êDK��$�&H������ߕ������W��2�Ṿ6��$���T}J�c٣�y 7����:��1��1mVycw����"[5��	gv������g��N[\}k3=��'��O73{�̋���Sǎ�5��wq����?G�����P�ڴj����ѽ���ۧ���6��_
��d���{���:O��=�{�6f8��u�F-N>AgB��k!]����4CD��ɾ}}bP�iMG]�*��kۅԡ����1@ƳM*��=ul��B�wAݸj2�öbJ�\Lu�J,���	�(�����͜<���c�=�T�g)�pa�Cr��b;ny��D�5�m�Q7B��@u�ku��'0p�h�S�#��<�T�Vw�<޺�F��m��[XL�U:�,vl6��J�f�+je�a2;oG���M�?5��b�#]��2��St5���D��(��Y�^�3)VDa�]h��y�x�-��i�&��ő�X�ٔa�*�;�<�۩�L�$����6��,�j��޵��pN���Z�ޘ��K0X�J��	^j��#Uf)�`�JG�����.�[/Vo.�b��ÃwO[�x�&	'����c,����$ޚ*o1�t)�j�(�fO�lѩ�/��bu�,�Ġ$�$�e	�7>�wEU����X����e��u��y!�����={�}�_��J�rc%�X4�i�l�Y�T��Cbat���Ubn�~<�������߮��������./Dȁw��ǋ"��-��w4��ne&eq�My��S�eB0�����;[�չ�M;������1���j;���x�tcw<}���aWù��4zB��n�O�E���S3�%����7"�B��sVZVna��m����Gf��ݎUi��e�4QE�]�m8�:�aN)8���[�s�-+���-k,��ש _T��g�}�5�lf�ǈ�Z �EވI�j�\�ʌ��ogS{ז�&�$��t�;e��`�j��<�v�V���E3e�Ֆq+7�-��$�$�i��Н�6����f �3�xh>�멣ճ��룭Uv��rK���rKM[	�Ґ6�C����u/�(�I��^jk�S�N;�6����*!Fk3'ۗ�z��W뻯z��>�޲֛/.�ޭ�����ي���*�9�w������{��hw�H�YՏN�kx�I:I ���;�݊���sn��{��E8,`)H'`�l[K4����F��w{��\_�����;|���STL��'�^���'� ޕFdS6[ʲҳ}��m�S�ΓzvM<ζ�Q��Ͷ�z�q���n����Ƿ6�l���t�I��r��o֯��q�D�3���}̖��_"�h���{P��/ gI'�8�ll�I�b�˜��[G�M�on!�u��`�M���&���\��>c/���m�JM���\kΆ˘V_*�0b�4ՙ�l�@�j��6����̏VEk&�(<ڣ[��-9��m�f�kih^������w��,Nw�=Xʻ���0��`�p��H�[捼�Ƚ@[��	�$�0s#/E*qx�0I8I���M��MЈ����*;7�{/:.�Y|���l�^�X^f2�5Q�
g!g�H��o�8���\����%��	A���!��d��A<�5�v�Q�4�t���X���Wn�X��vŭCA	�q���&I?�I��s�1��҅�+i1��wKfX#y`]υߧ)�sjڙ�{kƘ�>�ж���[@p�b��!3�/l�K�;Yrs�:i��wi��mCy�Pܐ��IOb�9���O��-����L��ݥ!&4�n�J�vQ���Ci��Q���ٙэu[�ތ���h�Jn�lr�\�� ���Z��2LW,���NDԱv��U�M���d;�ٖ�G�&�P�'�J��)�X�ob�I�dF�`�FM�fo�$�fڧ�>؝��o�I ����,���x%�
u%�v�����B�.�-���''�z˕x��h���m��w�;ǭ�A; ^�<���f���;TR7�z�N���۝A��-� A[�<#�l���n��g�G�n���.ㅋ��<��#��o���o����n��� ���ۦ+���&8U	�j�馲��bb�5C�d[�����X8����E�l�R��3k
v��{E`�B�K�(v�6��Iv��pm�]����/cLob���,��Mq��Q�'a�n���v&6��a$�1�H�1���S��{�0y�irL��ޗ�u�5��~��oNPi��P�9�Ů�ݸ�f��j`ٚjsC����	����s�X��0�I�#�{C�I�*_�_���b�4{�ί���\�>ᦻZ���8�a���th���7����f0	:�J�i�qw���'X$����нV#f�i�I�-���S7�n�|�ܶ��d��$�%/�J���hJk��I��[jW�vi�VC=-,7$�n8�o�	'I�� �I:{{�lP�KTQQ�v
�Z����
I����M���~��}�	HaD/����`�Ρ8�{�]ƺ6p�����u`#wVj�i���i��kV�/wx��oZm�w��l���j�z����XX�Y.L� �G�t뼫#^�o�5ע�ǷQ�_��
�����p���X��==H�/{?��V���jc�&ɹ������ϖM�:��x��\�c��Z٬��-�]��c5��KfX_���P��kN�1������$�J6DA���/li��9X�DU�fhI�}��	2I����A�Zgb��6�
��kxR3E�^-����!��}�����Ӈb-Z���o$�$��%W1>��k<��[ZҜ�(/I{ES�\$���jے�Ŵ�!�wg�h&���n��v�݉�A��;��fCl�6�kc�6�q���	=�`�q)0��l�l��V�*�37M�ǋ[�qz�͋�Jc�%&1���gù���u��j��YB�,�2��	(������Vg�^ ��� �]�l �����L|zq������v��<x��ӯG�������J�F�����T6�<[���nv�o��������L��j���.E�vf��B��>�v)Y��C݊Lv����� >N7��}�'&y�|�Χc�N��};Vz��)=�Z�����Y7�؅$��_�����a6$���B���y�����ۺ��	�<h�X��%�rcۃs�*���#~��{n1�����[�@5��o/Zq�u�B��G1�kc\vnl<�;�qwŒr[^U��&���V�w��M<�=:2���{�$/��#Nz�w�۞Ff���α��8��Y�yj��t��(�7���Ȉ��̲��3E��D⌃Y�Z�2T���n�`Y͛V�ù�.����Qc���b㺰�p�3)k���s��{��;��ǜ~G6�EH��OL�<ϻ@2g�r�K/�J��=���ٷ�$<�J�h��/p���{9?=�L�%7g��v�R������{����{.�|3~�;���W1q�d�c��	1{F2S\�# �Y6��p����d�F��ܽtk�q�z���d��d2�Y��oˮi9-.�:|���������	�Qϔx��Kk�7�L���d������!<��v���r1���)�!���V��}7�O�ܹx��tgp��:���w쓆���}���(���������yM��d{���޽��=#x�ƎMz�^zO�>^�yOoɋ��x#\g5�O��˰�r{G�_��Y��{R�Q�;����L�{�h�޸s�ڪ\}&&^����Mw��v���A�{�;�eWGD��� /]�p�K��-��6��%󝺈��׺�[~��$��I�2�;��ym���Eh�u��F�0�*���4�u�\�牃�#o��5	��F����|[�	H"�T�H�F�_\LE��5r|]���_Z�^W��bi(�Ԇǖ��B�5X�Ѣ"�h��ѓ|\��X�HF���A���{�����j1�K��(����"�=��[�u=�^y鴕�Nb��F���S��)\�b]�6���xY�������\��]	�/�<��zo"5�^oW˭�G������Y]-��z������/wv�wN��{M�^r9Q����m�������gwK�^{��K5�9�U�7�%���ݝ�c����ԙwo6��;�+���rL[�t�n��z�n�Wy�I�[}�\G����7��&��l�l�'1��6GT�=i���4A�p�]�z �[���i_:#�Â/: �-������ԲMuW�������*�ϳ2q�­�>wY� �ׂ,���v��]�xA�dT�y[EY=�y�8`R��,���͋������>/v���fD{˧��}ަ����_��l��Si�l�t�7h��ױc%-�F"�Ckq��m����>K-����� ݰ>7t�#8g)����+!��7��:ݱ�0�+�a@���#�����E��g���X��!�ٓ䂷��O�7���]m�[�l��"�!�ۍ�T������ �J�a��6F{[��t[7�-@۽oud f?�+-�H/sW�U*=v.t{/x@$n���Eݿ���]�����9��B���V-��t�G����r	������y�<2�h�,���0pE�j�ߚ��Nm=�4����O$f��QE�]w��jְ^dHյ07gj�n�j��ae��H�����f��4+։Nԩ�-�&�O��?@ ��rc�]�@/�ln��V}����n��g�@X�����n�����]&���M����J0Zs�*�W� �O�)aY�֝ې��.:�c�$�-kPyҧcf������9���e� v�"���W]��U*�v.{�{��K{2.:(d`yh"x8"��<A�`��]���!\�D���v�s=v�A �����<�9o=2�뼳�f�9oհ v��tY"�C�o���96�
ڽ��8".�@mଭ���|�F#p��F�B7��n7	�o�wX9�g|X�p&��>����i�x�V�@#��Eۇ�z���UA�]���^�F� ���#�����_������]��n������Ϛ6�p�x̳ۜ���X�/]�8�0+vx��Ȼa~>o>��2x��%�M7/ �`���m��9.����]�=�q��<��5og����j{���|��f{r9�ư��R]����0ˈ���Eb+v9q�v��gW;�Ŵ*�-s\�:�zG����7u��N#9��t��/c�c�,�X�YN;%A���L]���r�;'Goy��P�,�]x�ٌ�$-���&bK��Y�a�r���'V;xuZ�Gu��pm	�,���n�=q�n�tB��sZ��+`x�j:���q�<�mOi���crh<�\��f�=���o^	�����[��%�y�n�����qj����h��քt���R~����u����Â.�#޻`�o]�ۇ��4����n>I'5s;ܸ��l~w��M���7v�A�ۀ��`����T?z�la	3���(]��ީU��<<�{�#q�W�7�\?�����nls�e��S�Ӹ���l"_8�Ư��&.�kDkM�=BZ�,�PhdF�k2����l{�m@��E��x<��q��%"=��iV���y�� ݰ�VwTTvQ����ncp7��,�Ǜ
�Wѳ�w����{���}v��A���"���qy��*\߆��!V%{�*zY�ع�e�@ ������G��`�����Xd� �h����j��䤶��̪띬yB8��['���w,����z��s~]�F�O����A��<���aK<�ӽ�����#m@�^ ����/AL��������̼v��qO$�c�:���g��&^��s����vw�fG����2n�r ����p�*��3ZqL�A��w��A�s�Vw^�3���#y���=j� ��v���	Fn�h�[�����E��m^ �����a�9��Ԩ�kqb罗� ���|'���0�ɏsٌ=q�2�#���cu�M&@Z��ݻu������
��[��I��γ�������w�����]ۈ�l�]�.��o���ú�N�y���C%Eƴ7o#s���� ��pG�����ڻ]h�pPgXz;�r�`ieIi2�f��-�
2�4����^�88؃�WIc��{�V���W��D�����.�m�T��6�����G�B�n*b��O�=.��@퇮�A����ޣ�k�8��o��	���t��S:>Gyo?����5����Z��h9�%�x>�Ρ���F{=�Bݖ0��4i���^>^��#T��0*q�E���D �&�L��35t�q�vCƻ��ki�Ed]G6�%�A��ʻD:��U�E�n�\�Xۓ(m�Ƴb���{�znj���S��pG271�7n�Hsv�swo �6|"b1�qS7�kj�Wl;��A�`A���]�zx��zW<�p��yf����|��I-��A��8!O?����X>��������s�&�KaB�|��:+vtֿ�(9�o$��5��dy��
N�MM/ظ=�do�I�Ts,)���=��3Y�5a�Բ3�STٹ��$���L�}_���C��Y����=��r��]�����̎�a歝�ng+����2>X�}wo 6�`A�`��me,�)$Y`�h�pA
�?�]����q6�������A�>>���]�d�l죝k�gH��8 ��wky����Ä9�g$�Wn>m�������p�ʶ��	�Pr(p'{��L}[� ٲ��ݸr.�#Ç͡�vM�l߁�����K��.���&;ُ�f7M��y����13a�`���7�qtZe�Y���L	��^����f��ܗOW��<��[�0�qyX�l��4dF�[�����wtM峫��W[�j�
��>NC�y�WO<���,۰�]�p!��@6l�����o|�{�@��n�uO8�E����t�G�k�fdG����W�׎���v%�lq�d�\Յ��ϒ�1�p F٬�"6J����Nf" ���m �����?�l� ��xȹ;�¶8[���pt��q�8ܛ#90�Ay<Gk8 ������w�3���R�sU֐���{?��틙���F[��!��M�� ��k��k�7<��ac�W@8 �0.�< ��pE� :n%��9&�ꦽ��r�;T�dP��^oq��;\.�x���v�I��hƄ��s�V��� �3���b���Q��z��=m̢�%��75�U�æ�l3\�
"����Â.���v03�f��|�`m0B/z�f�B��#-�1�Aʷ��7m�����>�m�F�ѷ�hܸ<�γđ�jJ�i��]�10&��T@b�����<�-��9�)f\Bl��>f�&͛?x =���+���D�1�Opn�v��E�@<fn�r�E���D]vU����F�8�(�vy`㞶��,i�sŨ�n��0Ȕƅ%���m�&���A� ��\f:�w�����F��a�w�������,>��c4�5�:� L�-w0�%���	�+�����������2X�M�i�۔���IKa\.�٤"b0�����Q]�7��7�O�x���q�v��7a�bs�/E�`�3u169��x�{ԿkZ�c�9�< O�]�ˇ�y�q��OB罙��:�6�._3X �nG�_��v���9�x���]�21�!m��jX��x��9���p�AA��^���[l��e�ne���p��0Ƹ#9�Eۃ�.�x���qh����µ��C�(���\֢2߳{�U���n��ݼ]��=��^��o
 �W<B�pA�p���eG_N4E\�@,2����� !���J�|D�v�>�A���7m��ݰf.���7_����U�Z-�Pr7٬8���#V��.���7oựk�3C4�;-GX�'��!�����yj�m;�z��u{<������8wl����AM��[� ��A�o�m����r#�[dp�{����X5N��(�r7v�]���n�?�^>W"��&n8gG<L�ۘ��(��QV�u�wθBXx�?j��y�����V�;�"Z��3Y4a�y�h�k���yr�<�x7"���z+�A�8$ϛ:�rQ��a����^��A��g ���.���X���qK�q7�A�%�Ϸ��q���x�̲�&������e�`{�������)0�� |.�Ȼ`�]�z<m�,�v�������8�^�@�`�����OZ��DV?bo��|%���L�MiV��L[y�ŏ�͸`A�`��뻁͐h��!*��:�$������#Y=��8\{\8"����|;a+U�ᡛ},g��e��]0��hge�Zm��L��#4�ɺԖB8�	�>�f�+ʹ�H��87l��9���Ftgn����Nr{��oQ����F���� N�{N]�w^�M� 9�qj�[v���J=#[H|Kv�맭K�"+�7`�⷏�H�b��eVͱ��|0�x!0 �0r���6|�]����zcxmk-R����{�6�=r<ٽ�#6̀�S�=*ZԻd@��3�
Z�;��}�(�-����ܧ�X.i�=�3+[���R��P���^W���7�#Y;�q�Ӆ��`.�z͟]�� �|��r�9�v��-D8���7v�6�����]H�9<0�y�)7���1�W��<7�cF4_���E��	�e��7nwo�y���iy��W���7�wU��V�1�؛� ��$��s���1���3�[�l���D3�?�� r�Z;oZ�{n�=��yJz�Nv�Wk�h���r��o�"H�o��y�W+�o���w�{�;���7�巤.��0��V�r1dG�v��͘ހs1ǸJ��ױX���Z�|��p u�j{���]H�9=��)0pA��lUv�T�y���!o@>��p.��ݴ���z�$�r���q+��<�n��݉��j��A;�ݷ��x�n��,C(�{Oѕ᠎�qn3�n�8�z�&�;D���e끖�|'������Ĥ�)Pفw�ZC�
!�ܾ�f�ea:��� ���Bx�`������������9�����A�L6��	�h�N�M��{�����{�}w�7�87l����z�`�7l�h�{�v?��C�+�u�W���Nr�w�y�7l���.ڈ7o�]9O��{���l-��B\lS%ҋ��Z�nK\��æ�m�.�2ٔ�i��>m�il��9�������n�8����Pֻ��݉��-r���K�<���V3�Mݼ]�q�9��>�+ئ�ڬE�9�\Z���Y���M���^��F� �w8pEݿ�7y9�{������3����މ�(�l�圂n������|��A�=[����]P�9=��q�9[�gn�X�`�
�#����8��A���կ��`�䳫���ȷ�ov&�x��o �m�6��ذ�2[���^�����r���E� �:����F�p���Y����M�����7!=��!�kLg�Q�<q�M>;q����8���v��������Ǐ����y��d�x�^z���Ül�Oۥy��a6 q��ܻi��E8"����Kt����A�ǎ�o.����@=r'gg���ag����{Q�q�q$����i{q��l�A��,&�4��s ����G��!m�W�3Ů�h�d�'K=G�؏���L^N�w�G�J����A]��i\q/o/5�&�,��7#^�u^�A���7F�b�"�z�87.�n.p�޺��a���@�do���G��U�=�|gTX����ɫ����j�ޙ���sB�l��]����
9��oo�q;�(�����/���w7ޠ(\�T����@ge�{.�fګ[���g���ү`;�_yz'y�|���V�V��ճ��Ԥ����d�;�������{=���[��{�<�+�{_�wl=����H�{T�1E�i�|79��=ݳC��Y�P���[�po�x|�h��Sf��
Ku�x��d8|]���Y�}�;`����ً4+�Ma�<ݾg{R^~�{��g{�m�8�y�e��FXNZǂ"ȥOV%� sй����rf*<}����y��7�7��o��7s��V+��'�󌴓��.t�����[1.��� �>�{����Ϫ�A`f�i�?yU��c�N{V!�y��;^�-P��vф{4o����3jQ���^w�W�e�ܝ�^�B��nڹ��'y��;���F���z��ӽȁ����|�����n�|څQ���݇���Ϝu�^,,��zNis���Ou�Mrۻ]�n�}����]۝~��2�w[��gה��ߎW�]��k�sWv�K��M�s\ۺ��r�BKe��B�pz`��K�ж��Y�%N)�	͝ܮt�˻�j14#m&��3��{�r��=�A~7>8��[�М�HbH�yp͈��]�`��#FѨ$�7\�1ۡj"�F5y\�ŧ��1�%�ɤ�_W#mJ)*��6�)����K~wyn�@T��m��TQF)7�Q�&�|nDj �"��+��Q2h�%��H�Ľ�y���cB7��+�m�6*f�;�mi)�>72TW�]�h�]52�X#�f�w�_7矵ǻ�n*��&���X��q8���Ӱn4���N:y����KXl)q��,����b2���3hW��P[�L�9��>~��WgK�0����wn«�L��������v3�ItZ۲�l`��i���V�^6�!�.ٖ�,��ksc��V
#Y�s��v8ۓ���u�Y����M�m�Z}��nِ���8x�Ͳ��;-N
�F�V�;�ˬ�v�W��&�ÓXj���٭tg��0{1��q�<ι���l\K�m�ӎ����X�6�2��ʁ��;v4��rj��ӢZzJ�7&v�9��'o�����Bz�cÛ�5T��,�dt��`�X�#)e�r�V�%�nu���lv�0-� !��
��������Ee݀��gT�@f��m���bk к�M�p�J�4f��JL�憚��h��X�U.�L�j��j�۱cvx�]I��;I!ۨ{��8(㺙�v�ɹ,UǷ�z4Ϋ���;A�qL4ZSr�� ط�W/�lA�݄6Q�pC�È��
�<��6�u��S��Ɍ96��ȗ]=�8��F�l:���Հ��r�<b�75������L��tP++-�:�)X�1ѻ&���K�G����n}�q���釱�5֘]�.(�rW]�4]]A�H���9���9M���;V�Y�g���z�x9y��-#�&���F�z��f�N�|j��`Y�V/Og//u�����2d�\붅s֍	�O��|�@��+3�Ҍ��)^�6f�<�]4qnx�%�n�s��\C�@N�2����3Y�<�ғ�{W���[y�);�s�:�x�<�zQ�D5h��͖�K*l�	���g��	�N�X!{C5�i>{�.rM���|��cnx78yЅ�^;�G�'�����蹨�Ǝ�y�I�,TxgxM,�T�=r�U���j��T�Uėe�*m��6m�Y Z�n�ׂ�1�<��s�v���{�{CԎ\5eU����� ǋǢ*^�pTg����5ٝ����}��B�1��z7og^�F*@�L	8,�͢v��;�<ݴ��$wH`�7M�֤�Zq�1�s�ge�L6�L�������^�51u� ���\�ґ��Y�rJ� ����Lv\�b� ���:����3mc0�����1�.&�kqQ��L�C������Ah��qiZ?�⒪ՠ� ՇN���I�gV�n���򶮼�-"�g�5�����K~;�<Nk��l��n��2��]�ª/�0;ٽ��W"�;���f3=� ��.�?����H�a漃��Z���� x���j]��u�l-�Sw��[ǈ'u��ݰu����Ys�e����s�u��4C�*ȑ��ā�jm���UԵs���;y�[d�We�@$n;�{�?����.�8휀6���Tjd-�x����?�&���cVF��J��d߻ټ��v�|T^uF�R�〿F-a�05�/@aon ��s�}v��v��5n�Q^�v)g%�\��������A�o ���<n��ݸ�s�C=_^ձU�L$�4�;�I�7XJ�ԏ�Mgm�#��v�3)2M��DM����≯E�]���ꉻ���&�ٹ�G�Oe�1gk���	5��]�������y�Y�X�3��3��Kͬ�8�s$��r!�K�I䓹��o�>{������_�OǛ,z,��`�)��8��{��v��r�4&bڨ�#�{���/L>4�����/_^��E$��������L-q^]��n���<XɷD^��Al��.�8]�G�7m������=f�c+[cmk{��xw[���8#�v�]��m�ۮv=��a�nZ����L�fM�w��� n3��gI��Q�!E5���<A�`��v�A񻷃�`sٌ������rX2���XŸ�_	��{y�޽�p�U����؂Am�
��{��7��[~��U��G�R��5@S�Z�t#�\�g��B�Mf�m����^�ﱗ���.�?��j������:���7bn²v�r��O\Sivr��y�p|�/O�̨8 �`�>�w��h^�x��Es8 �8u��q9��φd�WxG�_8-���o+��0q�&X1��IL�-��d"L��Li�'�����u�+��Ƴ+�f�Ǽ�������o��=�ͱ��|���J���\�V�u��Uu��N��5u}k[5���(�|D>Q�m���')$^޷�~*`jp���y�p�����5������{3h �8��$���n��m��V0���/X{�����IY��r��!	�Ց�--���IL��vsA��s�'z�Y��������F[{u�$���$��{~�y������>5�~Yt�Vmb�Mv�H\b�[h��"K�����/g$�g[�og�,�x6V����fHnVv��I����xDU��a�N&��hǀ0��a���l<���eC2��]��`w޼��l�����w�+X>Ub��V��X���[�>8��|;����h;� �v!��� ���]���5�f��ӗ���E�s�10�� �	7����L��TwV�Oe�@ ���֐|�2C6�[��*������8�`�W��嶺�D�
~fJ7&�"*��d���z��V���v��o�f���;�H�ucb����sVsŌ���E;⸘��lN^zb"[��q��  ����!�)��̻#ʱ�R$�����>ߛ+�S����`�׊�:�)��[cv&�A8�� �����`�s��C	�9�"�t�bC�Ս�7I+v�xS^�e�9��r�z�����t�R����no�.�Yʲt�̴x��x��~h�3+����R�]!�F��!7�u8r9;���y&�A)3� �5���F���7�6���p��3{�2n�����y�<��Fˇ!&���yۑ�������a$,g���	;���ò4V��	�뮵��ӓ�-�����_�y�\!=���yW�E.�<i��M�yCm��on�r7�'^s����@Ǒ�]�]�������.US�6�u��eJ�s+���l53(�Ψ9���=���� ��f�}���uVZ/���)��ژL�BL+���ld���U=ܻ�AM�~+q��=���{BB\"����*FH�Zg��q�����]�T-3���a��i��-A�<����"���(ӭs�z��	��^+�2M�f�ˠ��v�(�=v-�n��l\}l`��B)��{I(����0�I�myd�@�vA���n�^���]617�D��9�J�#����[�ɽv�;�3�-�����&[���iSr��b-4�u���lҗ7p$U�k<���:�\i:Wn��b����{���Ѩ�m;j;{_V{���������!�V����Q ��9�f����l������9�ve�)6�}����y�l����߶<JLj�vV�K��ln�n>;nG:�Mf�[���pu7�x��%�(����u�;�=t~}�
:\�.���Y�{���1�fW{W�p�pF�$ާ֝E�B�!�U��x泐m��&�@)G�끡��&t�ok�M�"�zޢ����(��S��L�,�5���c*���t� �N��x�ȇʪ��еWDc�ln�nؙχ%=�O���Z���3��cY�>;���S��)0r
N� Vή��L�,W�Y������F�ѿ;����M� �s�[�mɑ�ߜ����>~�~	���z�Rgl#�m�j�!���:܍�o���i�lG<ԗm��N�%�Yg���O� �������̋�E��#��h�co%vi�>�p�l��a@���sfˑ�7��E�����.]�f�9��܈^�"����Z3�4�h�2㨠�[���C=�a�d�ϿM����8��AH�~��Uu��O��f�#�
���~��~�B~�i�l4D��s��Rmڒ�w	å�������$dPH�����n:�/��i}�-��-��q3�u���1�v�(y�v���#��|�G�s �'�f�୼�5936La ��xu[o�D���j�L{�Fk�"���E��¼@B8RУr�_f:]��A�C��g��L�z��{z2��h��7�0p@�o����-/ct@6d��k�!'�(��$���I��d�����y�#��۬�в��1Ŷ6�n֛ϭ�?�̓z
M�E�c w��I<!mߛ��h�q{���8����#�6Q.�LKչ���:���0&僖���ERN�co:�ރ&M�w�p\*�_��� �[a�&�e��-�=�u5�N��U�J������a�l�����g#׌�ނ����Y���gx���a
(�����n�>���@pA�9	8"��/7����|�XԻw?W!7߱������=/��]����朅�K,7�bhiD˽�k�0T������پ����(*�2 �(� ���i�����|3������ڱ�m7�kiI�Rg!�o�q��0��m;���aG�~�]��e��L���^:�8�=�t��)� ���q��A���!2!�*X���g�r�cYý׽��Y�3E�|��Sx?�#S�(����O
�vs�^���"�ر��3�<�3�f�LK�9�&��X�Y���+�t�h�t�)��Y���[����p�!2#j�fօ�|�-��cp��iݲٷo�-�(�8����L�!C��8>
�E#=8��~�'�#9�G7Z�q�@ɓw[�L86|���yZ���y>�5���u3�BdC��8 �� ���0�,��T}�!�b���E�&h���8 �058pBL�|���7�g����mD�g��t�f뀓V�f�[Wϒ���7x��87�����Z5o�TS߶��Vʖp���E�����Lp�z�9��I�� +-��ƚ`!�ۜ�e��6Ud�6�oPl�f�x{� j+Icm�ڪf���*�Z1�&���m�P
�)���N�*�'����y�Dv�Ȼ`�ȢƘ�rln�.n��5��&
��j��>�a>!'"�����g��L�i��f��wR;�;��1���n�q���D����<[��h��[�a�'���e���m�?�L��Rgw��#���E�&h�w�xc>6F���"�Ã�K�Rp�$�Gx�a�wK�n�X�Q:�]���_>S�|n�ow��F��$�N�;����v{V�����*��Y�����[���k��=�Іv�l�M��uz=����Ȼp�!2!�̙��>�;��OD�\si�s��G�g���q츫�����`A�`��T�S�R俤I\�@��C-_b���$��I�]�Ɩ��1*s�d��[����m�)�s����9l��9I��'��G���?z	�|�<w��B��3��O{Wlז�}�W���0~�p3�{8�8R>�v��,팟x������3a�*kz9�a�Bw��o@$�����T��&������*ٕ�f�b���kl�������?}�R��P7�[�kn�:�'/�r�5��H�-1�?Ϗ�MS��N̛Li��l�d��j��{u�d�� �7���\K��+���Z�v�v%������$.�@�c���0�#c
�K���+y)��L�csx�YvuY��WH9���Xݣf���<����n'��ا�sڣ/g��������������ܑ�
9�2�;tQHq�tp<X���7=ny�$�2���C9��>�a�5��Q�A	8H�j;���0T^�o��.�"S�M�.P#�����?�L�r�8 ���ʳ�>�[�kY��l��=��;E�Gx0 �0pF��(к�[�R��/�T�9��f7n��ȍ�г�Fދ�TEH ���dֽͶ]�Ns�ہ�g�ki�v�}v�E�8 �bͳ�Ӕ���a$R�����'���:۽r ��{m�i� F�+n��]~��V���&r	I�����I��Ev]�npc	��5���wf=%O��{�`M; �jp���	0�d5&ˡ]��ؚb�jڑ� )m:�ӎm��=u����7&�e&�͸��K�:��&�	��g��ou,���l�n�`���x�j�x�3w��f��'9A�]N��Z�	������[�6ȘGL�C*�$[���b��S�Is�^F=n����iT�S��h��#�Hqn�F?]��#�Kp͋���y�}�vK2[�s����/�	 A-Y���)X�Y5�#Y	E�BA�O9o����������n���o}�H�`��3\?�KwIh�+Vzs��c9�3�@I��)3�AI�;^�=�<������f=�M��/[�A4�9�#<�=v>�p�!'p��׻��A�p�V������|�';Z������R�DV`зa�����@R��&pBL� ��?�'R`�2�=)�ȅ�F�^��9������|����a^�'w�I�����]�����k��f�ɦ\/T��[�:�1On��Q�n.��<8����{�6� �o?���
LM.��߇v�c�U46pZ�xҴ{EآP�fAO��W�x2p�$�pJL�B�t�����8���yc�����s5��+`��,n�L� ���Rg��.���^8��U���tfYa3(�C2΁��N6��׏�nݻi۷l�}^�O���������8k���l�S͖{�y��k2�+9�
1��FC�@�C���L唬;��w'�q��~��vv՘��bv��_dԁ�Q+j:�D�\�`�=�'��BBoe�T���u� g�ܾ����:^��y��=۽~��@p���$�:�c�w�M��-���U�r�*�[xo�+N�����.�𔢚������p��C)1����(l�}O5�x�:��3���g��qp�SG,�̛<׷�d����Az���R���<Ӿ�u5��ﻃ~O������c
ym�7�;$�~��f�`�x�}���{P`�4�f]�̰D��["!�Mt'_{��4��T�ƾ�%��vA�ҹ���	�v�²N>!�[���>��|4d93v���UιǺP��l���\뭱X�2E�Ϯ��Z���P�{��Y�E:U�Fl2�}��޽�ޗ��z��M5�;V����-�z/]���S63�NAaQV ��Y\��;����}���wdx�_mS\�1�E��Ǹ]�|0(��'��谑��]ދ{���=��Nv���龃��A���(���H���&�Ll�Gs�6vw�s��č���"l`�����->>����wJ5ozk�7��z��ݿ���6/n��~��(�Y����w��[�=�.�*Gf��՜r��[�;�����Ə9	�S���cӎ�y3~'z��;:.���ݥ??L1�U�_k�Qs��;=����熁�Ş~�����]yW;߻���]��:��#$�I&��F;�,[�ih�͹��wQb����b�$���4m�sDҚ����ur���"Ɠ;� �놄�ˁIj	��v���R�h�}�����W1�Y�Cb�;�����-~-��QjR����-|�nQ�F1I�H`Ž�h�V��ԛa(����S
B�H�-$j���v|�p���ޱE�����b��P1"�T��D]��߁��&������6�J��̊ȡ"�gY��'�{�t]�y^z�ς�[#5���y�7�M$hhi������A�n�m^�l�������b��gl౸M0pB�����Nc ����-!3(�2�a�9=�˺q����H���ju�l�l���x�3��8)3�JM9Mu�c�ޏ,D� �I�{cRlB�e*�*8%�Η!�"֛��J�7i���~��;LE'
L��?���@���wkk�Ǳ�U�Ml>�Lsi�9nY�m�3-�fU�4S+�����6&&�zI��[;�+w����uUM�7 A�`��58r�Dc,3.���Lᬣ�˲M�F:h�e��l̷J`<�aDC��4�P�2u}d �Ս��L�n����o8d��4�9U�/��1t�` ���x�0r�7l#�u�^�x�wcw����r#���-�m��������G��x��z	��\>}�y'�;������)������{=ףS����}����݉�W��`��O���md�kf���TX��b�f��5F�U�V1P�:�Þ����n��� O-��.��d*�ȹ�&w�n�Ggvc̪hl౻�4�� �)0pA�e�O~����A$�4�5_�Ae��Kr�Ԁ�.鋬+e��p�:�tS�?>�Y~xD�X��BM�	?�(MvNa��}�Pl���Q�m���ɰ�t��r	I��y�R`;'|Z�87�3����P.�����/}���[�Vs�.����t�%�>��ˁ6�A�8 ��pRg>I��d�T�x��_L2y�YyoO(��p�%�u8x���� ���
45^<Fz��N�������(MvNa��}�Pl�v3p �t�E���fBU�.da����9�`|R`����$��l������p�rp��G7�3��!����m�pA���98rp� ��=^o+:�_;�QS1
�� צ'��eU� �y<��YHS��2�Ns��F(�M��y�d9hj�ɊPg*������4ND1���,�ZicU��cT������4ڊ�����?w�<����bV��l����y�^8�+�vM�6N�'��.7Xr82���z�H��i�u��[��VG��3��f[����ꎷ�kt/�P]���չ�Qf�mc-��8
\L�AM���&re�S�H@ܼ٫��lٝ�z������#г<�b[b���┵-�sr�����b�ױ��n'����1�^�k�vc����|��X����i��Q�*K5q�6-=w;͎qN6Nx���[�a����%���d�ξ���H�3���=����{�,�yٹ�ɶ!0m ���!'�׋ BvpC�e��;�� ���o�=ЭW��zf�!��7x��9�Rl��q%>؅�Eh �3�U�p|w�?�)8	4�<�&��Y-Bn'K<Xw[�X�8��m��2�����I�� ���L���]��3Y�XJw�w�<qߊ����������͘{�,���6�����M�E�F.�ϸ��	0rg �W�p�!)�}��x���D������rW=�vnWzCge7��5��"�Q�|������{���y�M�ʕ����(;w�㮭3�;ۘF�G��b�~�O}/�D���	3�I�ݎͷ/y���e����e�Rgk[=�s��zˇ������4�|Rg"���|��Ӯ�Z��e#%t\��r1�=:��g��"�>i��L�������˽5��WIdq�#�}xt(�mx
�,��|;����[*+MJ*�EJi`�Ad @��Q��Sec8�?}�l~]�S͖����8&���}�����1��\Ï4,ͮ��	���p�$��O����b�.����=Lm�=7+}!���� �n��u���� ���I��yn0����Ǘ��Y�.M�U0b�yp^�K3[�M�#H�W�&L�1����6����p ���.��Y���rUa��>BO�m�������-���F��L$��|��_���Y7�|m�hh�nb�H����ܡ��MS�Q.���]6��*3m��?o����F���BN�)?��)�X�r��1�)�=��U;y����g�3�g ��!6������3��Xh �����t�;9��m�ⱀ}�BSi�q���q��%�Nk81�ބ��U3�|a1�y�,�;k4���F.,��v�ó�܊��h֞�^�;t{�ԡKɜL}��l=��6n��ٞ�(���<yޮe��u�D�<�|�		dFA1B�[�xs{���Sw�+Y��L�jq�H ��9	0�S,Ϙ`r{�`0N�pFky���hj��q�t.�p7)��^k�s۬vmNwPl�2��cy&�|�� ��8)0���f�*jnZ��p���{Ѽ\������V��uÐ�y&��R뉹�mK��Z͓>�ڒj�`��g�0ͅ��lM�v�3 ��T�6�dw �DU���&���!?��� �����ѷ���q����Fveqhhg\��L���LL	0�9	�b�3:�bA�=a���6�qO��_r���8 �u��)2��؟D�����~�	fr<�8 ���L�qܢ�Ot�2D�5.�š�\�����8 �`�w\����Ħ�*���ĵjAYō�F��޳�
L���F�O?I��+���|i�8/�^�7��;s0%�8SeS��2w/NK�s0jelV�L&��	|�A� �5��w��}��Ư��'��<1/t_}�[���{��U*|��	a���q�4p����Q
]�\`���~����!z,V=m�OB�>;te0~�pF�!�n�ϒk僞��Q�g�v����-��5,qa�4XSi]l�M[��\i3������/�!�Q�1���ÔQp!'���7/t�9g9��l)�F/��(D�#q��2>I��Rg"mҽ��6y�b3�D�p �n��'WO?I̔V�7���#S�0Q��9�
pX�O��	��:\�p��y�""�W6tJ�Zޔ�xRM�|v����g �5��&�A)3�O��M00ѩgX�v��G�'ךj
��-�ٛ�⍗ �t��`Kfɪ<fm`�'[�}�HpRg ��8-��2!�Re���������rk����l��k�M�=h��y�Y2dm̳��k�i�i<ܥ��QV:�0&�����U蹜��Z\���++i�J�ّ���/�Z�Ow7?+������̔9�>=h�}2���� ���ﮖ��_�Ie#�a5�s��d�q;V��h�JM�hL�`;s�PH�tp��v�76��s7VT���=W�-�{2�tc�8�Y� fx�ͫx���a6�x�ov��=�<UAsb}���ܷf6]�)5�c1�%B�Tv&��ؖpՍ�飝s�.��F����n�m��e;SA��&mnր�ֺ]]˫��z4}*[�dq)�]����ԳV��nku�F<�5�70�r��{�<���2��v���W����������ud
[��[]a	�d,��[Lʲ2�#3(�zԱ\�ah���`�ξФ��c���a��g�3]x��ge�)��c�@cIk8 �M�2!�L��)�A���Yh]��~�S���݉l�D�p�|���`jp�Qr�p������p��q��0t����w�L�}�6���KOz1ۧ�'i��5��lO�����猲���f��&v��2谄3,�L��#b�������Wm�9+��g��m�p|[��`ߋf�r��dT.B ų�=�_}��`̻3]��s����3L�I�`�Е��QYf�k�6X�b�>O�%�Yg�><����L���V�����{� �p�oj�=�S1y�ҷ��Ek� �0p�`�'�`�G���6�ܿOE�b�;��3�J���z,�����X�p�Y_N'Z�&�?o$�*�*���/���W�r�ӹ� |D!I�O�q ���������|^�Yl�����n�n�L�n���MMWP��ʋH�b��g"���a
���q5�o-���C:��zot�w/����8&�|�<BN�7���P��6[�GT�[{b���?�%&|ˣ�{'���EpZ���L��%���`��ÑIÂ
LBN���0�Y�9�M�T*(�Z{С������95�I��	4��üm���A�<ޞv��*�����Q:̡n5Km�뭱@�'���q�q����0�Rp���!����w�󋳃8�ڱc�yÑI��7�|�m�{**k'rt��q3�w3��ὑ����q�-n�lFyl톮�p�~v��àĸr7��3~�p�(����z{i��e�Fܹ�͑�N�9��V��%�HO턣�8��y��$�L�;<��9.l�Ax}X7q��� ·����Q�VVU�~ z�i�+�7Kj"�ڛ�	�g 濜���0,��7�e8g��h	���}����j�A�w;{4E���a��p�|���M���]c�3�^�!̻a��3*�BfU����j�������*B�}���V<���)�p58r� �8x���-E��ц/39,S@�]4X�^Vm���빷���b�8�c]8 ŰXO�I����z6l5b37"Kp��G^���W.�2-{!� A�s�ʶpA&rg�n�G���vo�O�W5X4�0r�8{��b��3�����e�^݁ ��'�=�=y���w� ��=w��8j�x[bqY��^��Ʀ��s\���#S��I��|���0L����
{�s	 �Nsy&�*�jBF`;����jn ����G��>s_������
����h��Y�Y���b�w�a����9{h����܀ 3���w�i)�D��TT�"*Mam|���-������&r	ߛ�4�JLRp��"},�ޖ�K���h������LX��L� >g{o���`�n�	K���Q�����e�Z���ڝ�<b���5v�]6�!C�.���n�������1;!�L�9ܟ�Ro8&{C�8vA�4ӌ�5�kq�Go�O8y�x�98s��ρw����k��ɫ۶ꭼ`����qԃN&�9��PCv��-��h ���5.��bwxֆ9l��0��_Ł�`�n�9��$�	��$�b��̙��g�O4cF���b�m6����u�JC�����9���|}�(�9u��A&b�Gc��M���-oq�`1�M��qCh�Q9��$��Q
N�'.;v̴3�vy�!���+�N�\���0Cv��A�6��@;�ݳ�$�N�t����o��Nݻv۷oOOޙ��}��Z�kfh�4Lm�*����P����=�a�=����<ǎ{�b�J��T���A��a��<i�/�ś�fSq^�:�G�8^Ȱ������ZUO	`�WF��o�"k�{]��w�����L���4ov�:��Y)�	�}/{��xlɰ�s�T�s�'vG�}�/ST!��j�l�;|�Ca7Fz�[j.�����s0d#w7O�6�oD�1��Nax����;�;�q�7��z�o����m�=�fJfv���x�ᦿv0��{��w}�7��Q|�,A�T���9�o�[���?t�Z�X1_E�u�-Z��b�ѯރ
������^�}� G��%"�/3�;�9*��t3P3�%u� ��G;t��4�ص*�^Z;�+#oN"�̷���h>�=ssa��ٽ6�^�7X�P�8��m�=1��w�fn/K�<_����}����ۂ�"��O��Iܥ���t�{���٨�^��K���ǆ�/x�����i}�Ԗ�F%&��<��䝰�X��6@�R��\2{p�/&�̬��B�^6U����";�^��JH�O-��dB��]����O��'=ڧ[�G�/T�}Ͼ���w�9My숀%�=y��Տ��7�#�,fO_h�ֻwr�q�\I�3�za�^*�v�^�_$������_Z���XEn�mzulOw�/z�Lt?�{��{X�8cw������q^2e�c\��7X��&=�8�t�'�i��*~�`����2���\]r�S��I��w{�:�y<�^e�R� ��F!!6 �etۛs �j5��Tb*,lT2"��F11���n�wuF�.Y݊��\��n�<ԑw\W�2=�r�-�����Q�\Ż�s�4@[�y��t�"���ݪ�\$���\κ�5�r�yc��t*����^W�\��sInN���ߝ�~�]O��F����j��έ�掚�l닅���,]�U͌mr-k�-3�w�/�Ud���Y���f�eE�9�v�9o�}�}��6�K��E�b��ڬ"�Ti�r�Qю��"t��K�� ���`��tw ꑺ;u�x»������͞Խ����Rf�Ŷk�i�2V\ں[��ۊ�61̾3ծhi�%�#��;v�8z�%�M�N��f%7��vH�s�j�:C��m���W�ڔ`�`a	i��fe tv@�/j9���k�4�L�<ޱ����٘ʛ��c
�<��,i3��\���n�4k�H��c�D5`���n�m8@��C�)̻�f�8�2F�b��SCJ��Υ�룰Ů��5j���8�7�n�M�f�ix�ry�@a�]���m�/s�vp���ԕ�3�Z��8�On��>�{"���c���.!��j�bDjB3X��u�R�`�e��-+�VZqu��}�e�k�b� ����Bxxf�D�d��7��u�ۂ����n��jt[LD���=tspƋu�6ś����p]���tw-@��SxA���O.�������!�t�H�l;���N�ۍd8d��ޙ���ͮ���p�n�3F�Cp�܇E���z��٭\��jN���X����1= y}]$�/>��=qr����^G�ۧ������r�Gn/>X-[r�s��B���5W���7���c��w�3��k�n*�ixSWCiiv̂L��@5v�2c1nn�!u�&Ѷ�jNb�b�������P�)�t����A
3Q�sF[;���q���ذ��3��]���:�n�]���ł��.^4]����3	�\Z3��m�80q��kՁ�U��{Z����
	��U��@v�g0eńu�vS8/<�a; {B5¦���!���D�鎱�؛������zK#
�(�je�3������K�6㌷5�1�g";;����ຼ��B�K��fP���/�5KCVj�A��;1���*@\�t�-[���n�jۡ�B��p��=d'��P�F�Jؙ�
k��F8���<%��l[=vj�f� ���-�Q��"6���vQ�y�n�M۫rRhk�l��t��N�b�7`�m��P�я;mf���x�U�liۜ�e-�X7�,�TV�����@-�a�33K�1��A�����nS�'��x{��u��^Ѕ�ҧ��K!ms\A�p٨�u�a�o��?�[}K]
Ik���8F�t��vF�g*A۴n�����z7�>x��`���I��p�;�LX��N 6g{o�L��u�\2.�F���z����&�k��	�g>�hǧ��V��oQ��{c�::�����-����0���`.ة��ө���x7�8���w7nv��RaZ;�ҸM�.�"m�`=Cn���pA5��I�M�J"|�kZ��-�7Ⱦ(a> �N�I	0]��ŋ����^w���[8!�P�v�z�?�5l�� �� ���5�v<=��͙[t�}�гu��<'��95�ZÍ����g�'m�Lf�nm�Ź�.�;����e��p,u/,-*G0�1uS�Ut�i�KtC���pH�g �p�!&�>U�������`=Cv��:6ۜ�l	��> �����9������/?��$�g�֌��1�Q�X7N�-01���bX��bӝ��9޹5�s͔^����L4�4���w�N)���
d�E��<��<�>V����kōϹ@x�ם��c3��p���(&����O{��מֈ��\I3+L�̫l�-o���6�y���Q���f&��(�&wE��2ˆgm�˲�fYb�8��*uX�l ��9��%&.�4��Ü����ڛ��rEu;�y;�[yW�,��[	�a�[�j��[et�����T8Z[��;���y����e������ ���!+7=�ޝ���v��K��b��<v�l&�Aˎd��8j]�L���\B_�Ce뿈���8 ���n��t�|95�[�+xF�'��`� ��[y&��8$$�D�V{Nǟ��"8����T6p�?2�zv�M�����y���f
��������}	�\�H�]��x��p7n+����W�)*n��+iz�3�Z��6 }���W����\��׼��q�b��>�:`�=6�8�&�%�rLļ��T�|�W�a��R" Ͻ���F[?�;�@O���8)3�F�cM�6�a�N�ykO�>)6��k�E�|95�[�pAT�(���%�-n#m�u8w�]�pH�o?��p ��y�y#h�]p�_�lS�ٳ�������-��L�٭�A����m7t#Z�r�!�<���bC�u� ��q�H���l�[�:� v�7�P>��O��Dl��Âg$��������""��e��l��\>?�iN��[�'�X8#�����9I��Ro<�^F��a���u�row��ѾEw��p}⩀}N��3��e��zf7������\�!'I���&~��..�x���X���ۀ���9L�sX9I��Ri��T�fhN���ؖ"xFky�p�;^6��)��-�2����z2�W��b��㒤e��Q���@��u	$-�-�
v�����H�w��C3�0��Ú}nzt�<'v+t> B��
�������h1���g ��At� ��l��lfF�%���N���pu[p����Xޙ`;S��	�H $��?�56����4���D���jD��klU���"f
�&�%.��f,�Y�������i�~��0�B���%>���wj�s_�!�;P��D.��y0���O[k?� ��%.�L���滆�xyx����g �v8p�w[gw*�{/��p#5Â�;qՑ<�{�AP��i ��pA)0r�8 ���z��Xޡs�*�le^9����Y�3M����N�$�>I�J\[��VkaKG��n�����A�`��LUk66k�a�L�X�A9L�U$��5	+y���~�����n�9��[_U2�Ӵ;Rfrlh�p�d��<`�A����e󀱜�3�\?�I���H�����l��l��38.�u�^.r�{������f�f�ڴ��Ә����$��w@�l��V���F�]��z�F/o�y�����_�3.$+Dk����*�κ��[MƬV�W/�nz����4쐄��+��1�y9ê���9��x�KAS�GPCָ��b�D�!�ڜB�r�[q���8T������Hc��`��a�G��y.:$��׬��á��!AΖ4�Xό��\5ݍ��a#������}�=��k�N{�.p@�G�R-1D�lȲ�b�&�[3ep�����0����z���S�k��{��32ٟ/�i5�˹����,d�9""�͖�L���s�?��8 ���+3::c0mv�gz����o�4i�����0��1�!'I��8!#�Ssn&��O�k>=����s_�!�;v&��n�r�M�i��Uܯ_oɮ���ꚛ�δB{�	���W���̵Wg͛�.������_{#�ryf�ݗ��w'}Ӕs9�fʃ���cQ���r	I�o3w�7GVe㴱�2ۀ!�b�A'n��x�G�8���BNR`#�8���Oۜ�K}c��m�v����q7	�g�u����)56��c��%�����_e��ۆ��#l��v�f:jd��"��л�6.�D������Yn�#�Xv��n�8 ����v�ll���\�pF_y�]�l�e4�H����o8I��&AI�}oUsGר:1Ms�K�Ez�s�[��\��e ��AO�{'��~BjQ�N晾��}ϼSV�dN�0���M�z������m�[?�}9��D��W�X��e�57�a�Lj���060�.]�I��n���v��;�.�B�̾�ͤ3���Ӯ>�õ;�&�A9L����pRg ���7��>����A��I��n�\�er.��/��
�B�����3�����`i7���g�'󔛸>p|�Ň���5^�TOYy�,�L8bn �)��u8pR`����d�\Sˬz�M�7NvF�P�m��y��p�v��XZT�{)�D�,":[4j�*MU�!;�]2����s�=a��v��|iNِ3b��53�&�b�hp��`e��q��[��Z�pR�?�[�M��&q�X�'��0�w\=�v�gSmrN�{/�r�9�@�E�q���ķ���󂭜n��Rq�)3�AI������k/�fT�;��Pe�E�5���=��\�ˢ���?bn�/�n�-��5���q����ӻx�&�"'!�9�il2��bT["��� ����͍[w�%ھ�K���QG�0�w݋f�<��:}��9��2#���f�_A��}��')�pm�f6D	�#G4�@ ��r,��L��?�(�,�y�)�݈���p㻖�gSo$���[��BN�EPg�:4��Uʙ�=E�v3l��`��m�b,��l3�� ��ט8��-�m�nY�GO�i���u��T�]w�%�p��	�<�Q������G��[��5��5�yv[�U��(����V�����)�z��op�D?�-�=�FkM�K5;�&� g�� �iRh����7",͇9L�"�sX��|I���QE�)8��y�֩g�>Q�5���PM�{/�pA�D{v����2!�)3���|n�{~������m�I�Z�������Ĺ�w����SW���h���[L��Ц��&|����qS=�i¹3H#�.�����������6�0�l�n����V��mw�2G��y��qӾ �g8pBN��QE�BL�Jj��O�*w����'�{{���^�%���-�A�o8��L� �����=�=S� �ߡ���M��j�8֫�9;s��t7F�Hq�kp.������w�fX?�X��QE�A�N���݋�m��y���`t`���<d:��F[��dC���pRg[���=�W�x����t���Xշx�\֊;�	�����8>(���=߽7U]'�|ݥ�2�#2r\!�m32_�ȋ�9۶�J��mN�b��n2L�wՍ���t���C���r�y,*���m���~h`�5n����>�v����$D��_y����zO��V���-�A	;��Y�M"�ə�)��M�۔�R���x�7vN�<Վ]w1���QהXB�̙.�v�M��-g�����g$Rv���{6$c�0�����]�6V���{=p��z�YBm�Xf�^�|�W}1<kx�G��}�̯#�8Ό���C�A����/��3A�R8��Y`ɡn`�*+t!��k�H\�d��q�S���Av(������/�kl�1�HL���t]��ε��zH-���싥�/G�؍��%�#�CPQ��½.c��|A�(�tRT��� Fc+��<vuv�����;b~.��v�9���;c��Kx�Q�q1���m�R=��&�t�v��|��h���_<�7���~�\;Q�wj���pd����=�oG	�mVH�(�b	f����M���ɲ�u�rw�	?��
]��>l\t�����\�Zz��SY'���9	3�A�I��8�dm�Fj��X�� �'ٻ�'�� � ^o���8�9�5��������/i@���9��}V�AI�v�A7mjT�[�ݭ��C[یg�����u���W��7��9	0�x�dA])�vv0�[�#9���?��O}��/�dS>ַ|nYȨv��t�^��|sY��'�<�y�R�8	8r�U�����L�S�˻�'_� � ^w��?�0pA^́]������.�؞/{����y6!0&m@�̮%�:ۯb��:,���ۧ�m��ķl���������}�����Rg>I���o<�=]n׌�\+���[��b��`#Ҝ86�9')������n)��Q;8^�Q���l�)��*��7m��Ӳ�{�7���`.���&u��l+��'�����KT%�Ad,�U'�I��^�X�� x|�w����f�Ѹ|��h�H�v��A�o?�_�
M�O�oc��k;QF�W�����r��I�Qp�e�3(/2��nc/L���A�֢S�$D��F���`���	;�k��rwf3��� �W�m�9��%&}]�����v�gz�X��R`��=
��پ����ye�̼tT����6\31��n���o�a��';7j���h�M��,���?�>)34cY��͉�:{�m�@��g��L�,�T�l��&n�-���̡�v�r�ڳk������K-�H�?{#/�d�`Rp�{�{2�ܐg/;�|�a�ou�;�m��A�p�W;���7��Rg>I����w�>�^��p�9��طsN#����]�cG���?�=nٲټ����sʆ ���(�@fh��o��cӏN:{zv����۷n{=�O�����}��o����tBR�.�?v<�y\'�P�=Ʊ&������W�W��O�;7n����9Gh�4y���7��-5�BO`����/����n�e�#�^�Ҭ��D6�~�m�VH'�I�<�����*;��M��x�a��GuLt�ޘ��e�MGnN�E�֢�)�\�WU�IPvf8�⻲�;�ȓ'�4��S������5o|횏{|d�Nm=�M���zlUusr��ݹ;���9�ꟹ�hi��@ֳ����޼}=��ޘ7C�=�����sǸ��N}�=��M^X��#�qúFx���짹o�Gv�^�#�d�.�<�-Ș�Vo�p�����{ۧM���*��O[���|��gt�v�n���p�V��*\/<C[����p^�̓`��
>O�-��=9���i�׷8����m��KW��.k�I;�($y�,����:�,�>c������'�ʽ=�䏉����W����ž>G�ű��`|p�=���9w��OL�_,\�K�P�ڵtӦ����E^@yiH�g�yC�þj�u�:$`�ƾO�l~��[����4�f�o��������p�>r��6��d�,V�ώ��1�u��7��3;8֧=���=�YǾ����5���>�~Ʈ7̮�U��o�N�������R��/�|C����+ϰ��ܹ���6�Fz�ކ6�u�l��~Lw�����Nt�P���P�<<�z{�çE��\������)�������{'��'8�I��^񁞉��@�a�����z� ��YFϾ�3�DC�L`�TT����+�`	���o�|8\���X�!�2�� CM�"���oW4�3���$d��ܫ��~�����\��{�[����{��ʿg���毬I]΢Ʒ6��*��s���W-ҹy��͊��_�y�w�U����u��ו������/��yV�d��բ}=��)��,��o�b�wv�|�Qo��ƹy��ʋy�*��򋻍��wW5uݳ��_^[�I�N�p�nB�qI�TI�eW��Q\�����h��Ac�ؤ���W4c�ۛ���1����� *jʹ.ͫ��2)��7�nY�A�|� �/O�"�0i���zX�G��9���$��{V���H3���
.�/�Hb٢:��㭄8)3Ϙ1I�Fz^ȃv�,���'2���έۨO����]�E��L�ܠh���J���~��&��u�$�;v��u�\�*�^�87[���R.֤l��Q�9��i�t����K�u8r?�D>E�M�֦9̊h�M����P�/�n�6
l!��g ���E;I��9�-�C-���:_��7�c���s��]�qB�"ۜ(�v�r�5�f��z���;`o�p��i����2�&eo�v.4�w�ޭ��YS���a�E���L���ܣȣ�L	8pҙ�P�|��0hGU@�7]�m���RSE�-������	�g=���7�.�ױ��s4 ��k=?�w�q-�f@�^�H;9���>��f;�Ś����t��/P'����ʨ�㲦�cʴ����������'��NR`�$��(�%`�8�v\?�ܮ���$!�����}��o?���V��1��yZ�E�޶��F<ع��՛M�s�4�E�r�Ժ��bk���d�š�ڥ�>�oY�$��A�I�]�m�S����|�y�����C��M�sJV��L$F��ҋ�Rp�!&QG��6�*�DP����#-��5���BQ�������1խ���8n!�Rn�;��Þ5U��O|�L�T�fXfWL&e��7�7b��m�ud#P��]���A��E�y�n��7��n��k؆��Ͱ�p|�?��6�!���e�C<��y�)0r!������AM��ȥ>� BL��!8pBC}>�ښ@n�|��#w[��c�[�&圃���I��
L}>ot�97.��ĥ�@u�_.����٬����w,oR����;}�����.O_�O}��?�#e,#��Q�L߽�6h�J~��K���}�����Hk��{j�9�u8��9<pj�����؞8��P�4m`��D<�8M��,���ۍV�l[n�y�N���ݻp� \���q&��� W�� q�\��p��m�<d�i]]H\]�.�^!	��ؘ1L� �vbY��X�V8UN�ݔ�[d	a	��*����R�m�nl#�]i��ի�L��ߨ{O^�6�Cy�~��F��V�a�t^X��MX�ƚ���q-ݚA)��z��w�ᗯ�Dxi�I��}��6yt#j�w���\��{���-±�����&�M$�?�ۉ�/	兝�1�/3��:�-��[��i��90rl����-��:0�D[ �����IÀ��ݹ3�3�������Մ�3Z�D	�Uq�*�fU��̫�e�kZ�{��a��NU0���pF�9�@���Ǎ�Ό9Vs����#)���r��-� �=�A.���[[9��y�I���歓+nV	�gY�}�7/�l��=��������I��'
����H{�y���_�(�&`�n�b�5�-����_lK<wHu�u]thl[M���'�7Ӟ����߷��&#��:h�Z�\L1�����ܧ��䱘�W����i���pA)3���y�0��z�ض���3=��\��d�����@|0M\D�1�at�";�ȩ��t/(n*��~��]\��?�%���(>��q8�,^(���>��3��|��`�_W����F՜�]�pAL�v�r)B~����q�����g �&|R`��r�&0����kwec�]K�۾��oy�5l�X�$�A�N����nJ7nn���4��L�Rp��ݰ~��wN��jow�[8!�t��PEo0�jYϩ3�|޻�8>7lݾ�ǁlt4"aކc�Wn����3������on�	 �$�S�����3��Ƚ����kf��i��7���ѲtI�\7kJe�HM�uhp˶|~s�e<,���M&<X���ε͑�P��Oz��`��[¦a`�l�l��9	0pBL�T�s�S>Ǳ���1�� �XӘu�pp]ukw����'5��3%���!C���L�8�Zs-,e�/����w�X��>/�<���6�G�<�W�NB
p�mG����Is����F���;6�G�a��0���x��}4�>7=�4�o6��uy� ���i^���]*^�;��	L�#5��w��I����F}c�i�M��t�P#<�6k |n��7usgU�)�m���ZÁ���E��0�����˃��ݮ�JF�`l�����������/���i��e�4�iHr��V3��5��M$Rn�kp�'��0 9`杋A���&P:y�:7d�ՕJ]+b�ԛb��ɯ��,��H>�p�d�	8x۝�g��t�1m���B�cV�4X��8x�"\�Rf��?�^ ��l}nx���>��^`ǭ��wQ�ڶ�<V8j�Gy����EcT��n�;8�p�����:\����	8��q��Χ�\��P��yV2\�p]mkqͳ�s\w�v�>7l�������\�?q~ja>1O�@7l�	Å�۽�oo��W��F���O���y�q3��k�;��Of�S+g���t�C�ߞ[��V;+[`Up�w8ޟx-�H�K�NE+zi2��˨Fk�]� 3>�;��g�/�[9�L��?�M/�q�ξ��~�F!��ir9Ҵ%<N[൸A��υc)0r
N!�;�s�Ofd�Olu�&��v(�R+���I^p�h�9�أ�I��+��1����By�̦�-p��=��=�����{��p%��ڦ��{N[8�3����A&E�kK;Ƽ����W�-p�y[a�{���fm󼯜����p�!)�}�7[��r�&���;����BN��W\�M��D�umVN��Lc	\Ru����<�F�&�gE����^"9��v��S">�绊���@������-�Yf�m0���0�p޻`� ݸpQD�F�;z���	�L����"fZ�|��pNDx�s��Cψo&DO���ɦڗ�t�i۝�q+}�ww�u/7:�QC�p�����ǖ�+���ٻ3�ψ� 8�����N1rb�R�,�S�Ń���N�+p4���Á�����2�͋`�3��J� �|ͻnɝO��u��\C�$�1�h���PT����Ǯ�!�|�I�:���ێ�8�^��^Nۙ�/IrG�!,Ԭ��]y���9�[Iv�I��^Sإ�;9}M.�e�p�S7a#Z���S�,<��u�X�5���FTi.L
	^��Z���E�a	�{t���;��>`5qg�������Д���qte]t���;�����]����7Q���>I�?x�z��[i�M> ���74�Tuh��p؞w�du<�l�o
���L3<���9�%�>IÂ�Jp������U����<��	���4�C���n�8���duk ����|�L��V�Ʊgq��a�`M���EN'iv��#;��-��D̲��p���po"�@O�&�F=n��k �k>�i ���v��7gV�~'	�g9��y�.�T�r�Q�@�������QE�A�8!)��cfNg���x�3b�t���r;Sp ��r6���y�I�p]���������_����B�� �=\gmY� ��q=�'b
�|��a�a �.š��M����I�{N���)?�����}��Y2ם�|��;�w���
��"��탔��>�L�����I��$��M�ˬ�%�}0<���x�t������i���v7=ˡ�o��ڃQ��`I��1p�x!���s�<￟c=|W��  ~�Ӿ���?��?oٰ[������<0�հF'�(����w��*�.�e�<��72\&e��2�a���.�C��z�G.�	Ǟ��'!�jn ��r����r�9�2T��*��:���F�5��Ne�g3�u2Ǚ���+�ؘ8"�����M-��:�N��o9I��&p!'���֫'a��1{��ϙ[G�#�nֆ~'	�x�A���p��L�p[XP����}�}+���MSf����8�=�{�3d��n���k�Ih�$;@���ll�j`����! ?�oND_o;D�'"�n"b��+5��i��-�y��BfU�̫!&e+�S�Ɔ�n窘Yl]�Yݎ�e�S,����X�� ��BRD�v���Jy�]$�������͘������g ���������u򁖒y���D�^^�yQ7r�uS���[��vqJ���I��=2&�Q.��>���у1�؆��U71�ԨHh6��2Mo�bAKFY7J�3�8hO���`� �N�|�	!'2�*�4
�|�+�d�r3��ȇ�D_�rwE?'"��m� �����uתI�"A�g��e��"�0%&A	8r�0�H�t�B7\U�ޞ잣x�R�7��q���7\?�I��&Dn\�����A��l�Dr�!��D9�R��ͷ^Hz:�K�m�4�D�`R�HVgyo돠A�gSa�M>>I���i=�Z����g8
���0'\9Ç�p���wQ�G�s:i�'��"��M�=��`k��nr8�8
��7L��ޏ@)3'U�������[F��U��;��4��ynuGL#�<кT#�b܂Ă��vגk*��t�*�� �rk��	8$�pRg"7.A�J�e�*2q�����#��/�M����v��(G����+����H���'ߊ_���:s�Ϩw`���#��\�G!�sNv!ϰo��^�8�TŒ=����Ǹ��������ݱ�q����qP���i��E��p���8 �'I��ϟ_�_�e��މ\��6�=v:��	�g#��I���Rg�d3�l��`��	�k�Ō1�\�v=�y���u�=nLV�bf�-��;Z�>O������6Q�Â��$��u����X�uN��W�Ŷ�^ٴ��YeKԙom���j`7e�|���L��9
���_��C�`����
�p}��y�t7vֻ�ơ/��0o��9I��A���7�_G���\��,��um�3-����{�盚�zY���c99N4NI��A ܳ�@�O�M@�&�M$[��ړ�m� �2\8;����ˍ�ۜ&���f����-bS:'�� C^��G�[�++֕�Z�-"�t���DW�����=�G��L@�a$â3/�A��{q���۷��ݻv�ߣ����}>�o�����ӛ��ݸ�D�T������L�y�^^ąa�O����^���L��^]���<OӉ�rm"wt��%^��&�y�<�s_ߠ�ݽ���c<�؟�1�8�]S}v�9{}��l�Ȳ�Sv��y�qh����U���}�{�׹�<�O������	�ԮF-<�p����'|_
r�yO;�q�ty�v�ou��)pg��:�>�u�o�j��W��� ���x�{��.z=o^{�Q���a���t�� �=��Ǹ:���q��U��o����#�6�ᝑN�~������~��W-K_��Oa�f�|w�������j��G���K��u��bb����6Jʺ{	�r��ѻ�竲��S �lkrM+_Jf���6����O�y��|�-�[��E���י��ղ���;.zh�����^�hV��{ѡ�V�o��{�]Z����=8���p��3��Y���N�}ϩL>��E�\�Ns��G���(uyb��s��'��-M�V�߳r�xM�p���t��)���ƞ"M���;���d�t��:D;����9c��BӺ�f�����Q�����������]�!qQ����_�wok���{�݁�> ��]�7䛞��t�����%<�%1S���wy5s�P~�ʋ�_u���Ê���+�!��׼@XSU��yo�:�����|t�>+��7n�w�]h
��^��ޮ�N���ה�5\^ m5�g1��r3��I&���p��ǻ�n���-�M�'8c���#�r�`%o.)/��w\��5�8�;�H��܋�FɍF�."�t�t�r��*�u�ǑI=wR�/~u�bK>v܁ws��z\���#n��w	6�nAss��ѳ��+;�vZ��FɬZ���\,_���	���Pb������2 ��������Ow4��*��y`����� RYm��/Ym�R�e�����M�cD�}���a��7n�Ǐ�/ǻpSw]����Ͻ�D�E�a�j`����pie�Y��e��C�XYoT-�������q�y�zf�챧�~�}���!����]\�Bb�����˺���wf�9�\��ɷK\��3��1��O^���x_dae9��ݵ�EyCA����-�&nn���a:�5c��w^����utt��ގ:���>�+���9ɶ�%���ѻt�)�1�p����B�c��.8���@up�l)ê�M-��,6��R��,&v^�+B�����:�-5�e��fq`���ke�`�i�0�Wku���ی�!Nt���щs�5�&Ĺ�/]4[�d��n]�g<ʓ=smb��8�k6p�;uѹ���F8��.q;�ոZ�ӻc��Fq����.�Kt�oh���3��m�ӘȨLg7D+�[nɮ�bΛ�O+�ne��=�<r���<a=�9�����x!��Z�cm�f�-�^���X�F�;F�;-���d�mz��-g���N�n/:#��{�ɂ�f+`ش�f�Ŕ�u�mٻ��)��(C;��%��9�M��v�햧��4�+ј�����Z3cJ6��Ѯ2ԥ��v�8�3�jT�G1%��*[mP77ڶ�뎮�� -�ά�t1ɧx��Z�j4v��B(��CSZM����?xd Bג���]���<�Ek3���ƭH�m�qu$��ڝ��1�[V>��`��O;D��M��K��l�; Mu�oe|a�M��}�y,(qu�j$-�)��lK^+�n&�{�ε���d�pޚ�9��xZ�0iA�[��+��l��X��r�������U*��%�G��vӳ�@x���a�k��9%K*E)�t-��MA�i��ʖj'b�]]:�vGO������=��8�v�0�3aْ̎�A��ڜ꽶qq0i!Y�v�6�����l�`L�Z�UChipEcGj��d��2�mlI������b�GQ.�x���Mf��A���f�PҔ�f1ԓ
�q[�Cu��y[�T��UQ�����w���v׷�c�3X�������<���1�,�w'Ո�����;�m�I��Qv61��#0���t�m6.Q/ki�C��Y1.�b4ɘՌ�ĉ�
b��+i[��-*16�51� B"ioc<���ٍ�������G�v:��@����v�;�d�e�4��ӑ�n�㓬��d�&�n����p׷c�5�ph�z·\k�M;��l�8�i�%n�,�4V&�[�´���!GsN�11����ȑ� WQ��j#y�	v�q�pf���������Ð����[��&��q���q�)�Кy����h �p�cű��Rg�0L��`�#����EY��6���`����e���5�7T�;�|���Dn�q ����pa�%����̱�N&pBL&�	I��-ޅ�\�Kf*�ֆ|j�5����>K�%&AI�����{0K��Ю��8��!K��)7��L�����w�=�n ���m@#$���#=��3���C�ϡ0s�@IÂ���\f�e0D`݇�]+v�M7T�;՜��X�?�ٰ v��v���J�p���s�<�&Nmu����XRh�������B�\].x��P;��'?K��B��x/��������Otou�<>2�5��N]�<��v�ӌ,�����`� ���I�
L^o)��:�*R3]}#E��O�"&�F�XY-���A}�^@i�y�[ȻI�u�}��'hLƼ��"���������ft������ʃP�8+�?���ﶭ���hS�8�:��r�9��&锛,]<+[Q!��<|��L����	3�BN6b�����D���/0F&��u����bg�I���4��x|�Ë������L泐AI�fq~��}�h�O���V��{����Λ������<�Ð�����	0r:�XmȈ���:���ִt�
{�v��A���a*[��?Uo'����sjp���/f�X�i��`�Y[�İ��\�beqغ��ãw�_c�n�-�IIÏ$�1\�����bm�o�88��Б���{� �:��B�R`����L�ݖo�cu�x�ⵟ����ݲ��-�m/�����8%c78$ϓ�j���iѡ���k(��Y	�e�̲�L�4��]/��¯oj�6L}�W�Xr�t�S��Ű������s��iVD��'A��f�K������K��� �	�Փ��2*­���i��e4A�`�ݳ�A&p|��ļ�1�����*�9����p;�H!'�tgoi�M16�4g��8$b�<��s���z�©�9,��$�%&�Mn�q7J;8�����3�m/+"���p|j�9lI�RqCT�Z�Pu��ldL�l9���=�Xâ��A�wfx;u[[�'E*�볲��Ø���CD���8	0	0B�7.�bdj*�����S%;5�C�>������JM��޻p���93����{��c
��#5��=���f���ֳ�������z��BU�������k9�q�JL�� ��&zMs�w]�O&��l�k��������i���m��D&�8!'q0����ұ��/�
LnD�ٽ��%Uw�:����3���y��}���nn�i{Ms�p����m5h��]o�Og�r�ۦN��A�騲>x0�r�p, �{���{���;-�=!�G
�?-9�?R����R��Ә��|>��kݼ٩�Sc/>�677���x������F&r�!'���LoVԳ��+�[w���Y�FJTɬe[�=:���-b�`K�s���:�~Xuj��G�=���8�w��J�{��ɷ�MĬ�~��HκVۨS�tt���l�9�9�tC2�fU��ZW��ܺ� ���d=�e�Ǚ�%.�}�X����H�U�]�e��8���(h&��8���_�5ۇ͟]������͜S�/�X�3VikR��k;�8�����BNΙ8a�h<oRY�bnv�b��A����5��&qY}��ɻ��Ĭ�~w��l��u�m��|l���B��.>I�J�Y�96/�!���nn��Β�Y��[����	���|�=��ʎ�}漛�eо�+<l��謦z�hQ��Sl��Κ#�L�3y�6���&h�)\�MMQq�L��2ȹ8��(F#X���]c�g�a������< <h�.E2MX33��9��z#l���͂��a.)4�nd{7Om��-�N\6��u������g��(ۗ�='A�6�n 1Ӄ��n���pU����v�,4����r2Ɍ^JJFݞI�;��}����v�+�ǳvQK�A��j�H�]t���+Q��6�IKk�ɰ��Eڭ�7D�iyE3�Y��+q-�^s����p4i+wv�ǫ:������#����*Y�%�Q��	�b��N�4Ƴ�#��{g\���_��c ��[�͟=ێW<77���xi�����q	�:�:�E%-�s|�AN��tȇ)3�AI��j�Ρf{kl�9,��⭜r7��܌�I��˂Æ��y[ �����a�C��4xǈ��2_�]�ro8L�~�G2,D�]nv��N�Y�ڛ�䳂��� �&pB)��>38c�L�d0�c�6Qr	8~WZ77�5�v�����8p�//2Y8i����m>I��
L�"�r�=T;��ǈ�"��ų���;�6�Yx��<4��&��?�(�$�ވ���+nr��f�m)q]9�Jq�t]����(�dF�و�j:�`�A~��Y�o�������|���9{�1Z�u���M�"sk����fʮr��a��w��"Lʶ23(�w��z��N�j<5��));��n��Dd��_�^��i�K��}zo��ž�F���,Z�M���5��G��G�7~-�%M#)�j�"�~l�(���/�>]֏�~�4],�Fw��p� ��B@=�s�r:����o�� ��o:dC����Lw�kV=5<���&�П#,��\97���o���&Ka3�-!�~q�**�[�u��:� ���`Sy�"zg/q�53.�`�����A1-�}1�O~��봌m����7l=v��"�ÔQ�]Yq�7p+�e��5��{xs:d�4��9����u�JC��D,ڻ��ʎ�F6c�X����,�|���A0�!��n.{d^���I'a� ���*�6�4��[g��ϓ��,�m�8)3��L���ss&޲�9pxi�8o՛R.���Nt��I��8 ���&�����U������C�ђ����8lv���S{��>/��n�D�Y]��8��F�L��8�y�+�9]��FH�½#�����<�����{0<�eYDF�q�1��y���޽5c��3�
�7���:���n�yi8�o�xU�$'˖�0�ڔ4fR��`a�Jk���{�Y�+����y��O�XL��P��dC��9�}�d�=}m�-�9�g��L���s��w���\s�v��!֭����2t��������8>6l��Ð�{�!��_&o=��D?�L����u�8l~�n���A�������?O���'��)�?z-���af;A��r�n�
�lI��XaT6Y�L�f[�ã?O���ϛ�V0��"�x���˹��y�2�����4;u��Q4}������&&�En�8�;&�H�{�\�` �����FXL�jtM� �?�E�bk�]�c'�pES���r	8r?�L��m�3s�؈{�e9��Lg[�����7�)3��v��Q1kZZİ�����gғ�۹���y�&�����y=�#����U���������Ĺ�'��v�{�:�z�vL���nq���v5��N0�����>�N��Kk½r{�~�4r&ʶo�>EӇ�!�I��&p!2!�I�������Zϖ��n�����>t�7l��I�F]���+����z���ؗ��+S�����r���G�q;y�.ƺDw�{�b����n��_�z��s6�8!&�I��E�6F�+��������d/{���l	I��!�L�,����ʹɮsu[y:�e2��OK����[^�\�e�*��g�Fk �3l��oc�:�� ���8 �L����v"}�gЙ�+Sa�25��(��X���z����� ���fϠ]�{�n>EN�}�7��[�8	0q�3}����覰[:u����S?�0Ttht�-�����8 ���JC�R`� ���I��E]n���!0�̒�8��͙���]��/٬K���I��~?/�����	\f~����w��<��2\���"�%b��
ă錭}�D>�{���U?����� �*M��XR�5�͜�G$�BqcE6�H����nwYU�X��X'gn:��5։.�F<���n:����^�1-��tk���΄�{�֔�.+���9���6�ٽ�n5h=�:h]�n���\�a��Q`R��[eB�I�Kb��[��mW��7A�v��i���vp9Ã��]��^�UI�e��U�+�1	�P�l���7vB�B'n3�3���w���V�JL����8z���m��`�`��N��f��I�.�ɸ#����&�h1G����5����I�)5^�t��-��0o�XeN&�+��W0�Ӈ��� ��"�Ã��Ƃ�t󙩹�t"o9�`�s��c��Q]5nKgN�NSy�{X8)3�kim�Ђ3��.w�0rIÂo:N1�*���nr�;��y�̫$\�e��7�3�A�p����)0{�]��vy�����UG-9���W0sX�r�?�ww�C��l�ك��Í� ۬л[^��v�3ڶ9e�̲�C2�3,��f��8I�=[�=l-��v3�(��%�gc��>�g>�o$�o�I��j2�mɥ����YB��uh��lԴh<���=x��ζ��;YF��俻���>u��#�~1��g$�or[�y;�ȸy��V0�zHg�j���w��`9H�>��z<n���W�ӽa;Pɢ��.z���qd>@V�.�"�rך^��RՕ.d��Ȇ�D�n�}��y�Ic�5���������r��UR�C'����z�x{��������p+>�����j�����*�9��I��^&t6X@�7a�\����	;��Ra�uXn�l���_�Z��O=R�ʶ%��[�f��ky&�)0	H3�CU�+e���+Y�)8|��Oյ���.f2����3�E��cyDG�lH"����
L��
M�)0r�cf���c\�
�st�<�O',w�x8 �`�^�	4�Rp׻8�&��z���7��FJ}�V��AϨ:{7�Q�M-���0���@v0_;�t�pH�g!s�	7��=��]��T��%���߈Md���
Z�Y�|w���{��s���	7g7�j�2��㈢ �lrq��;�ūb�fo��8$f3�E� �Y{o��h��zx�p��/��1�Yߔ�3)̮�I�\m�ǧ<q��Nݻv�������ӷ���7�󜮼;��ú�Ŝ�s�
����FN��
��kK�3}����^��&ٸ�J˔NMg����7�ѩ�W����˹{��܊�'M��>�ݸ��n��5a��7��3��`Z��fz���z�ܞw�K��Z����7��''��9�{�_{��������Mޚ���YF���^"FE�~���渊��Qz�x�[y[��ٳF�pK숧s|8����G�}��>3��劧��A��fI�Z�[{�ؕ\:d�#^B�=����?ia;�0�<��`^/��y��=�t>�7��tk��_�4�����Oz��K!�}[����>^����%;�
o�p��$|�4m�h[�K��-�y�������IKN |vf���pA��7����(=ޫ�q��I}��^^�_����.�[�}��W	q�=�*�˷�>'D��B����V��� 6�=��7=����.�_����l�_�Dx�T��f��x�4Q���9\��|B.��q��~x�����>�j:&?�>�q<���`q����\Il'���r�ǓӲ���P��6C#�f�ˬ���YѦO�d�?1�`�f�8�_�=�)�q�g���#����ͽ�uo�]��o��gnw�3����a�H7��{|��2_=�w��e�p\nw���3�W�A��qw7�pP�x�o1rp�z2��^~�j���������vw�7d�-:wp*��/�����0��s���:��g$����^�r���7�
Ak̓?V�'.��p���w�\���IH����+ߝ�3�7;��0(������I��wu��0Y�a�wt�%2��\�Mێ�9���뫢˗i�rL����e�ęr�;�v�NnC��$��dR��1����_}��I�v��DE˅���.IΣ(�w[�!7w������Î�˴���wt�Is�EwW!�6r� !D�n3 �&h�+�u/��M>�ľ��m��w2��C ��˝s�&A�h $Ɉ��\��q�I�(��4R�&su ˝���˝ے\�'��r���s�!9��N�w+���#�'.��tNn�gK������dD��������i��7o�o���NX�n�������z��I��IÑ	�vM�ƙ��V6M0�v��7ll���}R�fܖ�V��n��MR�J�N�jXP;,���|���I���2w��f���@��V5���^b������3;�]�8\���BN� &D<��&�lk�2K6���1��
mq���j���śK,�LQ\�l�0�8�q�pF[y�L��:�����&��9c��zX!)���'�b�	��,��Be�gM��Y�2rn��ϑU��0�w��=��Z5��.��%��ۈ>7L��3_�Rg�W��|�Z���3,���A��`���&A�N:��P���tԁ�փs��pA�`�^���?�O�)3�"��R'(��ڼ���F0	5n����sSM���u�AX��E�<�MCq�c*\^�i束�d��E�̼eE�w�p[F����5�/;암�b��'�s|S�n_�i�ɤ�hE=�Qgk���}����.Ra ���A�3�Ki|s�h�B�~]�t���ŃX�O\E�-�i���9HpRg ��T�$�g��{��	Z��t��]LݩP�/l�8�^x'�;5Q�j���R��Y��/ߐ�]����TQpA	8|��t�8?s�S��󇮚�ە|d� ���*��BdC�Rg�?�w��!��n����pk87��wn�Wr�{w�W0pA��I�6r�7������]���x9	0>.
L K�ҙ����%�gn"���;-��8 �L�g>I�爻�
��Z�7J*癵�������g�'���/�;�R�����g"�{TC�`�"f��Ec�����)7����I�U(�lm��r�j�W��g�t�w���D+�9c;�K!=��ݖC2�3,��M�z���9EC�[o%�Q��b��I��zhs|2����F�ѕ�;O���Y �3R�}o�
�Y{����0A5�����\]�40g.Ţsu�e˘֛;�����+aquqZ���.�p`��d�XN��;kk]�&�sA,�)�#��lѸ�Ԡ�rs8��η4V:b,1��e�Y�9��b�5n��xu�[F�b73{�lpQ� �3,u�79E���Y��w\[� �/0��Y��T5a�ݍ��*�j�Rn�V�75�"��C���������,������E@M�42k����l[��Mj�ˑ�cݥ�;nLm��~�8���I�Ĥ���-_hf��t��:u�7�}��D�-��m�&i7���H	1z3�
���c^�k��Hm��gew�޸�`���nO<�n�w<&�oy$��'���1yK��{�Dk�:�������v�݋��L����%Qq147�T�����7[�N6��X�F򇷀��)`Ϯ�D�ĸ�{ow�-����o$��#]�ۻ澇���*�ۤ)|�������$��V��]�:b�l6\g��5Ў���.ķc�a���6M�ss���0@xx|~��
�nE�z�s���Ḧus',u�t��5d2�Uॆ޿�M��ۋ�x������"x�4�\�m��'J�����C�����z���A���g��9o@��R�r_�|5����c*�͊Y���4�\S8�fs�<۾�����_\�s4<}�Z��^�n�p���c�S�ө7��ww^w�ͼϹύ4s����#/�ع�\��M��JA���8[wJ���8�`�N�?^i��d厽��ػć��9��N��LN<�y&�y��]\v�4ߠKk��C�j3o2/B��v�!'�R�A�rŃ(��h�[�cu^��.3����M����2ɨseh9~��1��ޤ�y&���+�s��#�ػס7yso�&�`�t�� p�ȩ��.�^u��m��֛�u�8��B���+����v2H'���p=�yߘ	��v?�y	7�J=^^^���W��G�ܦ̆������P��<r'.a�e�;��m���*�;��4l]�z��mEī�04�m�����I�Kx�<mp���|3�O�����I�'q6����)Vd��;s\���ﰌ>gb��{Bq��;4��zἓ�&Rt���ih������4i̖�s%a���ñ�ݻy,G����Z�|����m.6��h��s^��	ÓHDuս�[�%�kŌK3��+����L�|e��wӈl�GWIk���[��"$ׄO+��O�g�I�3O�/;��T?�C����m��r�Cs�:1�����ی�4$&�-��eJ���lN���fOn�p$Jkf`�����l��sa��[��y$�7��n67��3,�ݞ�ns��w�qظ˼�t�\Ǿ
[����͂����9��7\�|L_2�4b1.��\U��/J-��pG[]��R^ȦxȊ�虽��Sߏ�.�x���0:����9�`#`�ٞ�',����2s�3��w�Vn�+����?E|�>	7�L������� �y�-�[�x�!�x��Iｸ��$�SC�g�6��Қ�k��4@�v���)b���hL�m����nQV*� ��0ΖC[�JL����*.�
�]���EL�L��v|����z��2LJ.��iw��U"�C���w��.�=�q������&��m�e���5����s�&I8H݈��j;���L����ҐlȇE��w�%��$�$ἓ�\�L�8l�qΚ�yE���4�7��v��흮�A�U/�^2LNI� ��9I���(w0@>(��e�:�3�����t� ��S^��w�#��կ�H��ޝǁ��Z���5��ۍ_�=��ợ"�ǯ۷�^��Hx�y	���}�=�.��=X-Zܜ����:}����_Q�垉��ʭ!��ݣ^{W&�Ju\�r!���t�E�;U/�'�c� n6�؍�\��x�ݭ�D���ze�	A����v:�X�[L띈�R�O��3�,�^I �2c�(P���X�Kq
����ok	�q��:ށ\��cx���O�� �j�m)*�C�m��kɟ��\�k[�j�f#P�h�v�v���m)���� �����K�mu����˓���B$��k��ha�g$C�"���e0	0I8	0̽Л�?lC��yڻm��Y4�{�4�l��k�t�� c��ڏ4C���^�;���}�-�sO9p�gw�����5Jg��v���%�����IG���(A}�RZ��EښhSo��g��CW��y��]�������w;m����	7����	7�wj-�#���^v���ӈ Jb���8-^�oNc���&�I8I��4F�`����\��n떩�wXk;�:�ñ�J��.������qI����u���Kѷ@���_W.��B��m�Jlko=y)��������M�������ڄ��뜜g��B�d�h� Gs�M�$��I�^oO�͙��82e��P�� fCX�������8�|��ܻ/'����Ctg��s������V{*�������W]�8xXٶE�? �}�������>�/6������n�W�N���=�yK˹¶jJ|�%dsD>@���zbh]㗩�wXk��[{�%>	0I���n�~d��E�xo0I9��흨S\���FK�X���`n��L�J}޻�G�������^�F��n}�mf��{���
1�7R�X����8!$�9E���3�@"�lQ�r���vzF��)�����n���|�����9���d�w)��ok�SX��oE2���nw��l� ��X^�I(�Iãk�P�Sm�2��o-�O��;N�*���9���,�?�uͯ��oS~��m��`�I�U���?s�;<T���uq��/�߿
�|KSwӉ9U�u$SNs`�G�j��93�6��f��\z
�].%�Z��iȡ12��om�ۮA߽�UM�y-��q���%��d���S�������@*���y&fwj��:��uf��í�4;fh=��e�<k���a����p�����:�NS�'��N3VK��8I%�/��0�,E0��0k,��4����T�c�1�b���*�*i\�w #XL�$���]��Ӯ��\�v�vAmLJ'4\E��z�y$�0	1q��g"c��Mc�`��*��v/
��[^wu���M�c�&��n�n�\�	k��0	7�J�w_nEΙ�^�g�SuL�w��{�P�m��&�HIk�Y�S]]/�C��W8I�76��zu�b����i��x�y���3��9�?!�i�����q��}�H���;w��}Uy�=���FjP�S�c�)�g[7��D\�Jب�U�b�h�g1�R�y�Gvv�J{��- �j�M���0뻀.�}q�4�2�R��b�ڢ�3�-ov7�O��sS�[y���h�;38��!ä���n\�9)'vw�۸�,�1���]lbY������=޿7��y$�:X�ݯQEH�6�r���jw�� ���5��q��0I8	0R!�M��D�����I�wgW;�N�@QyQ�|2��3_����5����$��&�J�GT�2�̼*��#*ڢ�3��[½��v��l���z復Yq�mV��I�,l��U!H�6�r�T0����f�S,#�[�	'#��I�L�ҭ��D���,�Ά��l����eK���Z<<wݻz|v�������v�۷������n{@JFn u�lk���P�.�&3?�k�X�=da!�{���;C9�l�w�}�9B��q�<�fT���vo,<X���ᆕ܈��wǭ�ӂg�l�F�M�G;����$�ޥ��ǽâ����	\�as��a�ǽO��e��'p�/�ӯ=�wM;�q���Ƙ���oo�;�C2�WA�}ܦw���7���b>�ᾌ���|3~�8W��v�{����k�� �ɲعa�ޫ,$�ޚ8Jcׯ��<|�л����:�\�wzI�OI<��7gw{��6ѹ�]ݣ�]��Ͱ�R��C�;�'����ud��	�����\D������G��7{._9�{0���hf�G�wq��qx�b�ӽѨg�s[F�=1������{��!�	Ʋ�.J�P(��wV��������\��ǻ�}�@^�Fy7�pж���� �.J�Q��[G���w��hI��b�^��'��>C7s|U�2>����`	Z��N�O[i|���({p�<�^�RO��w�/\/�u������oFq{��{�ݽ�^o�_i��G����M�/�����{'>�'3j\���WfzK����a�?x���d$�7du��ͳes�|w���}9��1���k�x�����,wOy>0y/k�x��)�#�=��:;*�鳽���{J^���7��C�#*}&���}3��K����􏶾��[��Ш�x�����v+�m
%��W�m7���m�cVD-gUU�//ZC�k$T���|�ݩ��.o�G���H%$R`�~6�s��ܒ��h���h�;��.L���];�������r���""�f���)1�䘌S i929��7|�{�L��\f��j76���/K�����޽8��L*���d���]�����2D�����۷�˗wN�����w[�%Κg�W��r��'t���k��b�u�6d����W.�wwu���w]��o�e�vƙ��u�f9�L�JD�5�ʼ�f�`��]���"O+���4E�wX��D���PwJ��fc�-�sr�"N\a���Q�L����We2�g9���q,K��>u���.cs>u�_��!���ȑ3:;�s�I6SFO������3M��1I\ۥ���@
*H9W9��.�\h������.ncHcII$3�����|�^��~��^���>�n&���\����N�,q6�Z���[�s�Jz�@ḑ��#�౩��؍iga+V�c�y�;�O(a7m�����L���XqAq�;�(�N�vO��v��N#giPz�ݭp#�ƹXTa�-¥��3u G@������0m����VcPDk��=af�2o<$��8�;0��,�i�U�vù�b�wO}��YI���v���[i��̺(�WH��F�!4[n���h�,� onZupQ�GUՑ�	%��Wmuҙ������1\.t��֐Յ�r�R���|�{s\�]���Ya՗�ӣ�N�u�<j�u�6�t��׸W�u�M1�]4F��B��c�gS��gm��כe�V����C��샺��n�4ti6Y�B)k�:�N�Jᖬ�&�h� M@�ZJ��KMΡ�֗A�JL:�L�Z[mb2�	�Lm&Ԁ��8c`Z٣�e�\T	��Vѐykgv�q�kxV,g[���ز��ٖ�ЃHL�.Y���d�v���z��cl�f��Y%�������U
�XB���-qhi�AbL�׶��c����Oժ9�5ۧ�ӷU��c�0n��9��9=�M��ny��9�<su�3����oE�h�2�҅�*��1��#��hm1 �˵�1u�Վ�M�7_vw�;�1�<�N��[��V�,Z����l��3qYy�#�u�׶4F݂��r�t1[l�̼;h���챇��ۍۡ�>���V6�틘x�) �Zu��A��7��[�� ǒ\����<tGQ�h�
�'%�E��nT�wF+č��L=�����z�<T���nn-�Z�L�.�z�0͈�����m�5Z�Y����n��e�x{g�λji���C����K��C��d=n���]����:.�`��������pv|��
F��}���o��\g�Z��i��2ݞ�X8�E��m�~N��7����|����A���a�]	f]ىwp�}�F>s��*��f��\��%Ĵ1��\F�<��Z�}����RwG��V���yɸ}���5<f���s�Zv��+��:�K�q�/bx��myzCn�9h�Utb Jlv�к����S�sN��ݓ�F���X�� �h��Au�$��iwm<��:88�Uk<v�I��l���p�z����8|�Y��TlO,]s����g>X[ �^����@0�q��R5��l��)��.�%ɠ���A�GQ��Q�ࡽ���&
Nv���D噋l��.לQsO�����:L� �q��G8"P̥� B���k�2Zݷ�����m���o�t��^Oq��Y�_w�Óy&I:Xlt��+#s�2�n�����NK�f�I�I:M�B3d�4�#TоL�\�$�&�R���D�3ם�kz/r�O�,�z����% ��z���N������k�=��b�#�m���=G�}w>w��ZY��#����������n���(6N7q��=�&��ѝ�d:�q=b-��RMWy;��{�(�������e�ou�/?��$�$�$����/^��ͦ�[�����9t�o��� =}�k�A��.<�⽞>$�ͯM��|p���pE�E��YI�e)+�p���7�7�N�]�_�g����k{��J���-]�����.XW7�y)I�Of��%�0��aZĜ����:M��JgD������\�F��pj������M�G?��>H* `�/�q��޵�o$��(	m��4̋�ż�ׯ�W��h�8��5�w����$�y+���������Hv,�>ir�BhSU��oA�'e���5ٸ��{g�䁍�>��y�tI8R�I�n��pL�R9sr�0ka�VD�#m�2��;�����r���z�2"=y��ޭ̞n{ރ���r���,���aw�q?C�(�:�UǂI)	>���6��TS����a���>_���b�#l�J
��.\��$��(V(�ي���f*��x�2�`�����*TM^�"�I��C��Aٺ{�Fw�g)��������I��y����&�l�n��xJM��x��&h���9����.q�2l��h������$�P{�����iw,V	�k͆�1y��Y.s�} ]�����g����?~�&,�6�#��c3x�x|S��=b��	�,���wBh�>G���N�������ާ%�v���5��S^w۹i٬�����p������M��#Ҩm���BJ�z���cf�KS*��9�C�Α����I�xt�~��� ��It�����[�og��ݝ���1y��d��wv�J������h��Ve�I�NK�m���5�NS^wz�z=��S��q�rG��k�(�-$;�z�6���@)��z{�r�~��۝2���[U5�5���r%õ�����z�|ޫ�=�J I:L���Fd���>8o��͌y�d��$���`2��o%\83��d�3���#CՅ�R�XQ�qmW��W���$�c�n�
�21�˻�/�;{-�M䓄�Wv���͌*b�;o�K0���+#'�����z���e����:܄�mSr��s�F"�����[ ��U��ͮ��C{�8�I@�>�2�d����Aɢ��9�*˲a%��)��\��&M�xj��I�]�6�_6�0������8��fk���L7u�M��y$�ig��L\��e�v��ʢ�z��ZJDy'O��P����~86/u�T�������{�s���EJѵ�s��y���̚AQ�W���Z!�0!���t?��6�_-�k�}���`�7��lBb��]���BA��S�M�w6�T��N�v�Ea�9�	��s^����խ���$�{Z�9�vֵ֏ ��m�ӡ��}I�|�`��ŭ��1�u���L�^г�L�/Wlx�A�x<9\�N5�Ҥ�t)1kc4��rWp&g:Ξ�@�r1cv�S���9{�,OZ��ö��yO���/����7n���X�V�#����L�m�;�
c���]*T�?��o����z���$��탏I��9�Q��P��!��&�L�q��V���#��<b���o`�|��s#��^K�9�N���w[sFwY���o$�<����5�`�9��Aj��S8��	d�]�3[�% $|�H�x=;|�܎��s{��I?��ݝ���]���ޓ��3]6Њެ-�Y$��L+ȰI<�w��+Dy֚Vz�^6�0������?��$�$��O������RS�y��
�#�jͲ(:�tmJM��a�"W�7�X��iy�9���֛o�]0��g�}�(���n��ʄ��9����:IG��w#���z���1��Qw�����O�a.[=��
kff���wO�S1^�����Uq�=ɶ�4�@���4���ZN�H�=��/��\r	�T��z0.	�  F(���u���:1�5A_q$�hໝ,�Ӎ�42:���[� Z�$�'	I螬�����ʻ���mlj/9s�|.1�3�$�$���6ͅƅ`^�dǈI��m�nz���(�m�U�Hؓ�\'u�z�7�O��GbM�n����J/D�&�+�s7¡wJLW7K��,�02�'40vp��7d�nx��e��㙋�x�C[-��^���ˏׯ=Z��$�R���C���M+#����Q��DBg΀/���S�[�=�O	�h۽�l�o�s���	F �{u�݊�M7ݣ��z�Q��8i@IG��Í˕���]TQ�͋S��ک[ؙ�W�`~��y��>t����8��<���u�!�B�BF�w��l���{?ǆ����ch�bjr��&�C-��#��I%#�V���B	�U��-���I�,�ˍY��M+#�npݧl&��D�����K]&�y%)0N*��nhuo��sƘuL����6�,��;���:�$���0e�~_�o��� J$�#V�7�I��I�n�U�[��f�{1��������&�z�I�I�nM�i�ti�oM��֡�5!��c鑑����'I��Aд���6����k�'��9�!��dv��.;R��q�k"P~�qz�v��I�L�ܰΟ��,Q�	`YS�e��V9e�W��{�|���]��ok��*��X=M�	Y�I�^�a�їM�	+40���c�O�l7;���*�D�:)�ww�{oN�N��(]Yb�Ǩ�"�D@�O	U���n,4����1a;��2,5c#
"آ ç��~�|[-d��� ���I�rS�	�E�p�ihY��2_9�o$����yk�/�}�]ZT��YB�lps�֍/7��&� D0aó�C�r��|�&�zj���뫄���_��~��+��̻��be�O��c��qv�$���tLƷ��xN����U�rvRПx`e�,<����-��s��4�A�]>���$��v1�˦8��A�`��q�-:v��q��y$�I�Ʒz�N�o?O�����0����uբ1��-}׭�xӛ��0)�3ؘ�W�N`��1����C�U���Mugp�y������1{��IGW�u0�m�4�{D�LĎ��3�Ƽ2����n��(s�����+O�5����mY�n���DͲ�ݜ��;׃67O���>�x�/�i��e .CR�4]6nɩ��CW"�`�!xi)0�����z�ㆄ�#��s�`�K]4� ������1�lY����PJb�/���f��f���&,�&ұ&2S�X���&���=��(�K�B����IN6ˀP���W=�ءݎ��X6�啡1�Eƭ`�n��n,s�6�n�:ၠ؛rj������ԣ��R�E_�O���BֳJ٨�rڰ֥e���A�wme�\�e�^ ��y �wމobo$�%]c�vu�3&Vt��Q�縩�o�w����oI�LS�Yț�z�͹�@�賕�գ)��-}����IR��8յ�A��M�[�d�$���h�\��F^O1i�99p�/y�L`�FQVz�#��&�/&�|�WX����s:v�2�f�ПW<�ػ^�=W��ov��Қ�87g�l0���o+F�l��g�k滷,�ӓ�lE�7��;�]ܕ䤠)U)J,�l�Ka�Af!ߤ>/<ˊ�I��N�"ֆly��	���o�t�V<��Ro$�$�I�z<�]�*�+�t�N��W[���!��Z�8�+�/{��r�F�I�LQȲ��[3a���e����Y�:�Dˣ��V�Tv�JjH�~Ɂ���a[c�a��a�0��o�}�K�3��o��;�l;���ݭ��I:L�أ�&"c6jnc��aR혂��^��k���~�������_w?�[�m䓀�d���N��'��DlN���c�,�I8I�LSs�K�1���Sx.Eټ�\�Ν���g0I�Z��׳o�e �Đ�iRҠM
�UK�bʸ�6���DK���ln=N��$�W�6�m�U�գ-�"-��~���l�0�w?�M����|��ʤ3����U��3f�_
}��xI8�L0��[��<�Q4s�k���j]>�i̳5���m����ӷ���x�v��g�����}>�O���˚�͏Pg�Cf	�?_Wӧ�p�Qx���������y�g�n�R|5�4k�ڶ��xwmk�V�F��u����{������TD��d<+�u���/ !y�qfC�o��������Ok?���8M�_������ٴLz{��u�C]�]O�%!�f@n�>��(�����n'&����K7C=��0���5��$kַq����{��]ȧ��{ׇ���fy{�γn^��z�|�v�>��$�5:OO����.�~�uW%��os�a�!�#v5��3��1Wk�/q\�S�ieᚦ��3���>\��Ň4�;J���ڕ)��|��FOL�#���Mzd����y���	�wp��f?v���H�n,Tnx���{��n�}���P���4��x���^��9F�7�{ô�X:�qI�N�O� *N�<��Mr����|N�辡w�w&p�Z������չܷ���i���A�^W���#}x��>nq��m�58l���~��iJ�R�m�_/���:Tk���v�Kaŀ�}Pc���6k����?�]5���Q��ˋO����~�lG;�����Y���.���ޚu�UӗC�3ށ]:;c�a��|=٪��{k���O�p��U�ɋÁ����^�<:[s}ۏ&���2��>퇢#�;��c?wu���'c2[�7��c���on{ޤl� �s�;-^雳	&o��L�z��o��k���ܞ}y��h���ǻdxr�`�(���˼eo�8��[����x�����o��v/L��Q>��d�G����_7�i=r��^;M��N�� `������H�'.DN��{�� ��Lk�75��^ZJ��%�]�Q���Q��d����]�/ws�����]"'wh�����~�*�t�\���wnBW.b��p�g;��spwt�{��6yш�i:ﾮnl��Hc4ɢ1S�����W5����tɲQ�ǜ+������t@ܺ�&��AF�M�d�:�ܹ��p1DL�˛%��Q����^��r��d�'��4�,�R	/�s�?nׯ;a4I}kp�II������d�.u�hD�`��J>u�B%/:0.�7^\���{�n�Q'8��T�L���n�����>.�/��K�]y]E�m$`�6�^k�ئ]�J0�vh��$����
1	r��`��ܭИk��+�܋
&s�W�u�cFT���R������)�d�$�j���|{~7�l�{9�2�l�oᘀ|��I��J`2�ׁ[L\z�nU��J*�f5��F[N=�;��o6��黨�pR�{۬d��&&�c�܄��?s�9x)�"��$��&^��	;`�)�&,�ͳsE���z����)R���jM
V])��t�f:���m�^�@�?��; ���	��IH	Z��;
�6e�.����*�4Q�<�o�y�cZh)'�&|E�5��C��҇���mYp�����a��*�e�8)U��s㗯v�&	*b�e(�@�b���M��	&��0���&	0IFV=�;���jDNy���
�ك:B�{Ʉ������e��7�L5?�3ٍ�d�1֎y��4d���y˶g�>��G���r�1�
��k&r[��7��r�S����b�2K�Z^FК��/��f)-��m0�~�v�]���w	&�\a�WQ[w3ѵ�-�.�Ӭ:����3w|��}�gvJ�z�\gdbKPGsIӚK47���(�t=�4���e�L�e��fB��oQ����5�����'�ooi�a�N--���`s�������LNo��yQL
v�	��������ƽ�a,c�d���g0	U�S�?L�y��z��i�~)�$�$�C,���d=LV�V����TVwxN��d��o$��":�q���$�20��ӳ��=Z�a�KE�Se�i�g[����N�	7�d�V����Z�h�3��l7�i���"X�^���n;Y&�IG���v/6�0�Đ�C^����S��N��0� v�yq]:k>�1��xIA���Ы���E|A���χ�#s`��ޣ7[�D�Ť�A��Q��K=X�2�7=�ײ5�v�T��.�;����5����8�lnK�:��\m�FL.�=,#d�Z�7\�j"�v6�h��X��T��u�x������\���.�4v�0�ܘPɤ��uz\\���P[F��ù=<	���?}��o)e��fcVW.�3�m@��p]M`�c��:�dbͬ���|��&�z��_�P�º��J<-�]	ZLH�9[�	��u�$v�Xa��;�����JBL�w5��գ-�.��,���-��zj�$�7�I8~U{٨*�۶�u�4�ާgו�-�o^�+{����(G ds���jL�pGS�l୾.�	z��3=,c�go����d��R��z��Ai��v0	0���S�գ-�d*9}�ӭ�ٽPZ/�;�+`�M䓄��P��kS]�J����cJՊ�����}�,l��a�k��!�j��;��`K�H���XL�ͬ�
�I�bkyB�.l��]�Z�cPv�W��~�oL�p��'��Y�wz�t��o���b��q�X��k�I:Log���B���\�ҝ�d6�1P�����ڙ$�����);l�]�= em&ڛ�r=ci�4b�I�w.������.�Bjt�c!�����{�ς�u�<���і�x��/�i�{��Qa�W6kߦ#b<�I(%�R��,srfo�4s�Yh&�}0ۜ���ʓ��|���j����i�$�q�ݷ7�������{��ȿ8�d��1��ӟZq�iY��U���;�0��mSJ���bk�������`3ݏwo�x�}zi�9��h`X�;�d���l���l���Ɛ�*ζ엱�As����h�2���0IV�պ�#�*�A3�2n�b%�o|�׬% �����w{#g��`.����AGh����}w�;��.4�!���tR�Ã�8�`/�$�&H�mE��s�/5��#;_���DN�i�al���b���_{xI�H���~�o�.�ћp�|o�z�ޯ�>uj�*[��Ղ%���mX15�E������Ҕ�&�n-b���j�L-0�Iq�Ӻ���6a���L5�'�]�~Yo8�e)�I��$���Ύȡ��"[����\Z+5��{3��d�y%8����{�Nuf'-��ݜqk͌&��E���cP3a�j�	� 4�m67$����`;u��y&--���Z15�E���ot�,3EkBрK�%>JG�'�-��%W�<r�2�uǤN��C�tه'+_�K7��Ҷ�y��WT�ߧ������I��p���;���M0�A��\Zkﯼ31�{�.�]���]vm;]��Z&��v��.�5-�ƴe5�E���u��x��Z��;�i�ti�Su/Xa� �g3����Dэz�h^��C�M�?i+w��S9��v��շi��h�#�Y�7G?��I���$�M�y�)�[ۉ�p'g6!��EÒV����J|�:���WG�!x��س�<%7d��A���c�ݻ2FJ�C����U�ۛ�������2±�IHW����Ztu���|ڣ.f{Y��ӌ�T��7�q:��Uo@���l��o��Y��h�k���׼�{��W�rQ/;���C7�'�ԥ*J��?�	)ңU㦱Q֡ۛdd99[��g:M��G�Qu��L��!�u>��x:ous�$�u��{�GHjY���/�}e�<��ۦ�ܳ2�ݮ`�y$�ۗv{"kz��o��:.Z�"�����[y$��}>�b��������O�=��	n�Xƴ��S��N�Gg����SM`�<>x��x��	ӫG�\`
4�����oWynw�禌���||z�*d�U�\��V�g^��kZ˘qF�����J6-���s�v.i��B�Y׮.{<���q]�:�>�jD���Ұ��(�0͈��9H�:��[��t�Km���&�klH+^I���Bmut7'N<Oyw�&�����a��^��ِE��NK�G��̻���3��%m�ٳ=l���,���sf������:�E����?�PC����:����^���h���f��f6&�$�쏽?V)�L<���p���1��6UI�k�����] $�'�y'mv�Z�����8�e��U�2'��4�_w�1���c��|usVw���`G�L]���+y4P�k�	�te���r�y3av��7��R>JC�M�sEowC�֮`O]��Yۺ$c�3��P��$r���ts���fy���
�]��Y����[�F��SW�����,
Y�������G���ֺ��D���Є�d,m#�P��������;m�b�b<��3��;�y�َL�$�7��W�t\����G^�I���\W� O7��\G�H�y�;�a�_i�1�g*%D����Ol�#r��<��.�a����M�p�
q�L���u��4�'���w�=��rBy�UN��o��z/�_˵���/�1�Z=P�vjV4LtSV�u8-ڷM�I��:��A��Z�dKWf����bR�}���p3��L��N��T�6�H[�r�W,}��t)kY3av���t�96��山��`�0$�L�{-O�..jg� ��?�S4
��z:$c�8���z�R�I1<���Cյ���y�sej�4!�A�ÖnBG�&��nF����nX��n�]0�o$�&]��˄�w3�k���@�,�k7g��+w�ww~�V9��c�E�B�^<�թ���
Z�d�]������$�cO;�ܚ�j���8I�o�y�h�C�mgM_4)-��nQwM�J`�m�yN_*�W����/h ��6r}�^�$r�x�uG�k;}\�j^���a&�ݚK�Q�>%�i ��j9��lHǐqh�C}�d��$�̞��ߡ�<X�p����\*3y�)f��ެ݀(�DZ`�=J_���10����'����#V&��)�X��e\n��T��&���z�lI����8<��i��A6tY�C����cP�BQ�z�%oYBYY���1����"\W2I%���Wi=1�\ɗ8ј߄�>[x$�}wp=v�86�0�y���N;����w�%,����̀3��E��Zm��͒ɘ������<�p�w����V弞&%�ř��r�2�S5����ku��O�������>�8M�X�ژ���h{��tN�qh�a^ow���xnۤ"��:�-��!+�ۓ���>y�3��g�`k��@����])/n�YHC��粛C ��V������N�/Mv��K�s�*�8���o�p�P��8�[�m#�0s7��e'�0��o/_}�=y���yS���#_>�o���L�f��L��0�稍e5�\�庹%)�As�\y�|��՘�I����*�:6�S5����Ӫ�b�qs�f��M��p.ל�I:j�|3h��-Q-9o��i7�����$eo�X_k��H�B7�T"�7<V��㵂L�%�F˙�=�z�M�����b!�e�C.��������I�N�z�$\di2�K�-�!+�93{Ѣ���d�]��ް�
�{g�뽋-��y�wn=v޻�L�k��xit׻�3�q�y˪�+����ӭQnsz3�s?���1�����H�� Z��*"/����� @슊�n��;l;�e�@"Q�ٖ�-�6�5fZ̵�k2�2�Y�3[3k2�e�f�f��l�Y���l�Y��-fZ̵���m��3[,��k3k2�f��lͬ�Y�ٖ��Y�Y�ٖ�-fZ��̵�k2�c6�6�5fZ̵�����k3Ve��k2�f�e��Y�ٖٚ�6�-e��-fZ̵�����[3[2�e��mfZ�ՙk3k2�e�e��Y��e��Y��5�5�5�5�-f�1�1ﮇB���1�1�1kf[fZ�ՙk3k2�Y��k2�f�e��Y�Y��-fZ�e��lͬͬ�Y��-fZ��̵�2�e�ͬ�Y�Y�i��6�-fZ���e��Y��-fZ�����ՙ��fZ̵���k3Ve�ʳ-fmfkfjf�ʳ-fZ̫3W��vm�m�Z��L�̫3���m3m3m3m2��Y��6�5�*�ڰ�
�F��J�� F"�F
�F���b"��QDZb����F�E�E1DX�cE�1DX�cE�@V5�E�1DX�cE�0X�cE��ب��"� �",`(��"�(��,b��"ƠP��-kfkl�Y��-fZ��(�(�7@�)L�G2�f�e��Y��6�-f�u�e��ٛY��-fXccc���Y�����"� (�F" B����?���A��}��P�S�{��T��Y���(��%ޕ��G��?�����F�1򟂠 ��C��O��T�$E ���#�O���4��⟞/���K���E _g���l'�{-"ס��L��0�Ȟh
��(}���$��
(�UA$ d@ ��5j�֪�[U,����Eb�"�bE��DX@Q`!E��E�E�Eb@T>Ԁ�:��J���[>����",���� �H 3��!��?7����@���a�v�g����* 
������5����(���!���0���:>�� vZ�>�[�S � ��  ���2����<4X��+��>Ѿ v�������z�aAA��:M�:.<ttY@t� 
��>����O���օ _�<8�Yt�~q��|�?7�}��z0�@�O�������
 
��7��?� U�t3�1�D��ؘY�Xx���>����=O<�)<�{D {��%^�F1�ô��4Ӑ,?���~M�~�QPW�0(>:�(�+S�z?f�;��!�'��PVI��`��r�:b` ���������                                      � �+                          �           }�@ATU)T��*B� �PP�)!@
�IAI)E%���TIPB�EP (�IB%*�*A@{�  :U%%
P� "�^ ` c�[��Ѡ{�TX9	\�u���ҍ۠ w{�@��J{�ҎZ${�    � �>��� x�;��z,s����AAGu�͠���t �`�S{��xn{���މ��=(� �T$��  (�  ;�Q�APQ�HJ�T=��{��݄��[�����zl�C��K�@�Ю��޻�UR�wT���6�Ҁ�RIV�@1I{=燠   �  _uwr�_;H����J��6� t	{�T�w�{U y��$�x�V筭���(Q���AT�����wmP    �  {꒥"�BEU)BJ�^��*��{�B�; '����k<)Uw*���Х*�o`
�{�J����ʅ���p9�    >   t�n�E9����H*�t��������]���P�� ���(���
9b��  �   ���*PII*���*�����©Yj�U��%
��)A�U
�IN��
�mT��������@�꨷n
���       >�O}�$���T��JKp3ۨ�Ozΐ�N{S�"�p:�*J+��\�%
�4��/{p�LC�J    �  TH����J�$��>�T��s����@�`&�: FrA��@���{� ���G:�*����UR��=�   �  n� ;nw >�Δ*�Τ(9�Ѝ��a��G{�{�p=(n �q
��0@rIA�����2*�   S���)*�i ��'��J���h0�6J��R�`  ��U)��   $�*m�T��h�O����o���c��	$�Y!fx~U<��Q㯇(�Q�����$M�?_��H$�������$O�@!$�䄐$�I���!$$?��������[�Y���Ĵ��vV�N�5Gq�+�r��tk��Pgt2��~9f��O��G�I���G]c��+H�PmȦͫLʆ�)���鯵��`��ŃX�ӷA�f^�@��v=�V�sʆ���m�8)��U醱b�30��{*������˚o�t��]��-ؘ�f��᭥2�aZu
��¨ElUmn��U�s2R܉Қ�%���&�)��p	��eV�@ۻn+����Sϱ�i��c���2"
���V�F�U�[�[KF��b�*�ں(�ejz��U<� `�Tj$W�w&oRۺ֦a7�m�m�Sm��J��3����+5�Т�Dn��6�%�Gf��n��L��0neTJ������n���4�.�	��p���U�R�+�4v���m��a�퍬u#pǻ�E�X�,��x^h�y-Y�&��F/�R��������+0I	�*`�:�]���X��,�gMk���Yej���7+,�3(Y��Я0�6��,lx��y)7���!Ƣ�70E��mL�Y��퓇$Ya
����v����I�D�Sn�ٱor��q�q�C=An)���v拓2ERjm�Y`�yP݊��u7�U��ܽ���te�U�IvqeҔV&�%f�"C����6�4���m(6��-6���6r�ڙl#���Cu)�^Z˒�1�F�k2�����xs��kfj�3�b��f-Ʋi��L�[cvӬ��j9�/ni��k̷$�JGJ�oq��^*ݲ�f��MSt�;��Ê�+��W�z��f��ÇkX���gn�U\Z���^��U�J�֝:^LFip�f�V&�6
��%9,o֣���̖*��kJ��U���m��P�Vu�VJ�����-'��K�R D#�N���{9{I1���[U�	R&��X�
7N�a��n0��U��T�!x�gD����V�4'`�"�<��	�ݽUb���f�4-��z�B����;���x<�e�g�U4b֝��t�ہ]-�U�6;���n�Ԗ�e<'05�mLa�z��p"�*Ȅ����(<�J���n��Xn7Kwr[j�2�Ed[{{�
*�M;NU�P�׷k-e]J�B���ے� AKC�HC��f��j���u�j[9Tj�XЪӷzB��� ��f���D�;U{�m�D]���dՓCsZVDp�/,�W�6�3&͙�ա0�5#cV������&Ɇ*�eKǶ�ZH�kP.8��l*V+7-����˺�C]d��Q�{Z�Lڛe ����:�vj�]-�:U�����R;�u��3X̲����Q�G��ʵK3
X���F�b�8�.�b=����`X\Ȅ���mm9+.b7X3rV�[o���5�O:f��X�2��&��o�)Bҫ��u[���
E�q��Z�,���k6�)�mnf����Tj�x��ԩU����Շ�~����4����3I��L����Ҧ��X�"�1�nS�f���e�r˔�����33r��.Mf���yj�`?DEl6�N5��h��h���:)R�z��0��:�2�k��i�/h��d<��i�ٵ��L���U���W����-J���fCcіrfn��Xh�V)��(k��,��k�����mT�74�ݿ�V���n��V%.�ZQLuN4����lWM�fZ{���",�5�؎��uD%�c^95��M�����y�RC.�e�Ȟh�7&ԥ.�(��0�F�t(��[t��֖��భ�1��Hǳ/r(���Rd����,�2�2U�^Ci�j^�7��18���̸^�޻��p�͋��.�^���r��eR9p�"�e<ۣiѬq���Te�4i�pg�s�b��"�8��9�:f6��VŽsFUd��e����F���R�ŸmJJ�������թ٬���x*3���Me�6F��^ǯ2�$�,�KI)�V�+&V�ݥ�M��ݍ1�R�P��#3�c��FЪ�e;��*㉻�d�x�]2�	G��v^��C�Kr�ӿ^(ΪlU�W(g���mf�Z�8�T�]�r�E(Ի�dZP�lR�"�'E���
�eFfķ��ZCʛ���VԱ��;U���F�h[��:�6����4*�
E�N�әY�b�9gd�v�E�0��Ѷ��Xͫ�N���,��oj;y{aM:��^��\�.�hWx��҂:�1B��ōw{l�+)��1ŭǶ˳�����P�Lt(�ؗ&UT�ٛ۷�9d�Q�z��{�])@H�5�y����5�6��歏��70d��̹�K�10LȮg�7�k�C��Qm�ӻ�T��^	Us�*�,f�]�������6Ń���1��
f��-M9���,W�z*�!K�0Ѻhf�W�����e��Y�w�5+:����2��R����t7E6����/X�o]�Mlco�X�W�!���Vm[�z�R�L��aQ�a�׋C7�_}�N�V��F���)�vj�X�L�1J�U�F���A�U�b�
�� B�:��MW̙��L����6hR�IzFшd��mb���I�zn�6.�h��6���uT!�2TJ��.�d��skj˕�7��*��q�yV�w2��klM��Lh���/s2E2Z�U�w(Ef�^��V�+p���6�Y��a��AEX�m�S�Y!�0�-+A�IV�¥��bJ;�� lI�]`B�6d�J͋�f�8+lI�۪�SJ�F��?��x�7�����X��Y���o$��^��ZZ)m�vV=��0m0��mխ֜ǐ��Ő��حػ\��S)-d��d͏.���j��û>OQn�=�q]T�Wn�CX�R�L��+p����سo1l״�Zi��O�L�1�k��Fno�T��Js2�
ɗ�q��i�"5R��U�)��8���lH^a�X[�͸$nebV]��2�flmMx�����uu�{b�j)^���GYDTRh�uR�Z9��2�5�+sf!(dU6YvL�{H�
h�U��Č��yg/
��F
���:�oe�7��ʆ�*�zh�*��V7��V:�T�"��^�P�F��ڹxV��I��X�a�f�k;�Rռ-��*���{����b*�ݤ嶡ͬh�����j�[�{y�!�mu�ss7��׶��Ge��iCU�]kѻ�YJ�UV��*�;&�nG��yR���fA�]�d�W�yT��Z����#ڴSnf$�f�9�3U-���I��:aWv4�x�(U<4���́S�j'�uuR��B�iͿ��T5���V�f�3p�[�A��гU��;�+U�R��A�U[̙J�mk4��X�^a�.�n^m���Uj�/�{hS�q�R��Rw�����X4eJ�F�5�t�UwUP�F���ɵ{v(�4q��2e-��u�/%mn�̲^nc(��A���Z�n���7E٬6�T�{�R�B%���]�:BX���LW����Vf�7�72���m��kc�4����;����pWڕn��X��J3p�)+q��
�4fil�w'[�H��b�M�W��!���U[��k)ڪϷfV��R���h4��j�n4r;?i����mF�sQ�6`5��0Ϩ]��]J&ޛ��������ze޵Woqn��;�ՒL�p��8f�A0c"�[��hm'���	CҕA��v1e�o*��	�o)ձY��*�^ꪇ�խа�.,:9�uH̖�Z�l��X��^)VX�q᥶��j���F`��+���Y�'�JY�JW��xv�,g&a�K�t��[�v���!L��r<��[�i=YlGT2�,��oU�y���L�7��bJ�+�ʱcq!�t��_�
8e�d�Jȣ����)��TܵGK�=��!��o-QD�ܤ�MyKMf^2���gѭ�:�̦����Mkn�UD�u�q[�s5=a=v-�����WR���kER�V3EƎ��lQ4��!�%*�DL{Q�N�y�ɓk]Q�W�`;H$��Z� �㌺����c	�]M¥Vm,��;�����s��<w��KNKߖ���
^��^�V"�U���U[Wuor�ad��KTö�n�;�T�,U��޻�	;k*�RB�ު��؈Ү�,Í���UTu�B��J�t���*����T��hۖ���{���c2��	]e��:UB�Fݭ�*�C�a�#7C؄�'Ӌ�$y�V�լ�/0�h}�-Z"deo^ݞt�\�,�#@�oa��k˳Ibf����P[I�S�^�b���|�9sNˑ�V�j�)*��-j_*���t�O4[�w�y��S�d�dF;.*Ћ�������U�$�q�jf�I�w���䣔f�&��웹�~��f(]�4�m
Q�����⯡E2���6ڣ�*�x0���W�DKǢ������W��&$���/b�%'���ne7�����┚�UxkCeVn���*�N���$����R�ZYY`�8�Ww2��UY�K�1u�ǃY
��:����ǹ��ZIV*�߬f����Yf�m��K7)��X�]X��h�㎮ި��&���,5}f�͗x,��vR�^@�0I	;tw!"��ҞCMԙ4��l`�*�$�+�m���*����yP���cp֪�cf�he�d�u�c�mX����*	���B�:w�X7aۆ�4�!�j�۽r��vV�����:
���<M�FfQ���ͪ.�P�Vsu��(ִ�A��I�tq�3��B���7w'�ӵ�mئ���(���p��r^2.Mf�yvF<�����ɍ�̇1�ڶ��B�ovcU��A�BF�T;%�u%!UF���Z���LE��ҒǈV<����!��CYY�7��M�r=��ʺ��X�����"�W)o�vd�וzEn[�h��b�z�r+�B��Z�{�f��嘤�͐�ir�nfhE*��r�߲BAx�'cnm^�r�8�ܳ��{F�ɖ�4�;��~ƥ鬪-��7�v�n��Ί�*'uX][��eM;T������k)��ّ�k�M՚n�0җ�x�Wr��#�Y�W*a�mm{2U�[W�*�ݱ���
B���m��ݶ���uW4�q0�S)ͼI+Vjڻ�1-[�#�%�e�h�+d�jc/yW�����w��V-֐F;�j5^�u�C8T[�/!C~A�B�
��h�Gw뒍"*ݬٕo1f�,�Y���0�A,ݨ��#On���K/V�b/�~Q��fFt^ӶLy��a�����6�Dn
�̮:.�iO�t�n��C�K �����vN�J�K�����Z[H�7q��v���<�\6���xpU��I���CUwB�J�p�	�b[WZ�U[W�dR'��n-:Q�) �����	�]��V�P�޴��Lڨ��j:U�dw��}���U޸vmk��Kw��{���B4iosM۩K���Y�-ZL���+iP��;+C�)��u!�*�^�T(=`<�FRD[��%��9%�U�E&d�ā˨�L�0�͛��=׸�7q;x���֒�lC,[�WbA++#�ZΥ2�Z!�YW$���yb�kk�����Y���Lz���
F궪u"8"�kfdڳ�l8�dU���T��N�k��t��m�]��)��v�zvf�A�j��e�Vf�mPV�V�JbU,ͩLa�Á���:Û�,-;ۏ�(���iӢf��	��Y��y�C��
�h�m5W��*5G�ɯk�n�4Ȭ:�KV3j�
�{n���.�'�5y�e��/2��0"e[?MҚ��ͬ"�{�|�Q㽣���ahB��yCt#�<�Ga*d����,d�ʽ����Vp�w�ռSM����4$�m�;�^�p�ӣx	�U�K��UYf5���u��.��j�aTGc��͇����L^�3*feRgl�,�Q:Ѣ�h�7�݉S�j��U�� �Z����T��wg��yr��E
&J0�[A�&���9����u�;�gV �n��.�n�iP0ިk/u��Y[zH����nS�{x�ݶ�R��J�osSË1%ʲ�~IK�q6I�I��F^���27�%iKf��e���A0�g4Q�̇
v��iPћ�6�,�SPe4���'�Æɛy���Um!fF٪g���B,���eI�[%h0@���&�M.n�-��HK]固�nn3
65!u�]�2;Q�k]K.�;%@�b!:��+0df�С�*�S܏fnD#4��)} �fl�۫"d�X����QKh�T��n?��ae���2^��wj�Z�aݔ̬H/�܎�ܒ���^���q}r��Qn��G�LjF����(�5U���ʖ����s5��Ow)ض]�����
]��i�mݹ�4̻٘b�Ǧ��n�Y��	�,��5�)@�U�V�+��1���Ԋ{Ks&hQ����bD�TY��]slE��E��U�Ce�7+0*ʁ�M�v�)LP͔%�cZf�#o����5$ʤu(��r��4)�p�t��d�Ϣ������\�T�o�������L
��R�u�ސol���m��d�J�V�P�
֢nW���u5�+F��]f��WL����r�sj�2��jEmB:s�M]�wu*mSK�F��*�t-E^�z3u8k�m��b��K!�/1�"��{l�u���!�K15�j�$���WT��Xb��m-����{����M�����(��v���Z�U{��hu�. eU�+6û�(�1�<��@r�I
�J(�ص�yWE!�r;��e��V+�[��'^�i�AE���B�W�UU��.�Ek�����(�~����n��������v�4�wv�Ȫ�nȣO%̸*��]�u�)+�ywyW3V�"ħ6�|r'"�`�Jղ�P�gM,��R�uc1En�̉�E2��S�7:/.�\66�^ܚ6��SS:Һ�Z°u���ߞW�t�~~���	'�"��TU]%UE]���wD�H�@"�H���P	$���$�@�a$ ��!(d��$$X@$��(BH�� �,$P���E$ E�	�X��,�E�a$�XB@$P����A@"��)$�) BH, H�H�!$�,$ X"�		HI"�(HB)��	!k���������+�.�B (��I"�! 
u�G]Q�u�EUE\@ ) E� �AB �"�,$�BB
H,�� 
�d�YI$Qd! ������*�����BHHH$��?��?�y_>o.���Hv	[�7��\�&�;ŵ��C�r�����[�}��a�k�Q;Te�Au��9���t��/"`��ۊ�\��oZ�Y��*^�\�V2ѻ�VRܝ�{�;�-�gm^�u|s�	�]Js����UȜ�]�P��$�Ssx��I6��>b�ox��B֮|��ڵ�_�7Hp^��P�/���.��wJ�`�HX;5N�ZCksJadCUp��]+C��b�(�CZ��[p:�E7�M�YQ��붳�7�����Q���eu��rWXi�5���uc#%e8���V3�gt�7�\��wI���Ʊx���3����/1t��Ϯ�\U�ruƟݱ�T���NɕҁY�hui��S�s���m�V��j���<ڗDW�{*{������W�a6rG�u����ar�>w�9��ȑ�,�UK�CϠY�\f۩�s�'�ņ�Y4+آT����!Tt�R�-���r�eh�6��U�z�;I�/n�X!�|̱W:�d��e��mP�\���E�Ţ�WΪ�^H�'%�)ќ����ōL�n��:�	�k��Gy\k��"�&fck:^vA���yx2N$�F�Y.Nɕ��+���`B�����U�JN�[�w�%y�+^�v���C+r�N���c?^�������d����J�͒���ʭ��/�7}��t_j,;��ݭ��|���q��+�L��ܻ0�xͫCs�3.��5n�t�Zd�������vU���V@v�2��x5Z7|c�"��zԽ�oi̺7��k�s�t�72V�އk2EͤOmT������+�G����
�R��L������e�*�-z?���^�x�Y�˼��r*�Rl"�a�����*&��\�{��:�j�&d�c���/y|����a���Sf�	"���hإ{]y��������hQ�ɢ����U��[K2�H�;vb�y���{	��Nn�x�VQ4�m�vP\��uVC�xȫ7�9��j�4�@j�!���Yk,�n�K�F��&M���]�0S�̊}U�T:��<�H�o]�c&�,��75���n�Ɋ͝K�n��ζ�����4���3hAm��x��Md�b��c����`���C����AL�u7}@ӭ|#�
��g��f�h�]y=���Xw�ڷη�bw��;�uUr��|�έx4u5�M�	SY,����yd�ܻ�$��8�uɯ�v��Ʈ�q[w`�M�B�^/�o��';vM�ݵk����ouick��l�ŝJ�$䢌��cw������t�M��v�*��s6헝��qd�>�l�R5���}�h�i5W��Dl��&vf��PGC�M@�3�$��q2�P���aN��q(7O�4l��ڝ���C�1>�-}He��OU��}�
����Jܳ��ݬ���Э��2�Vf���3Qѹ��+L	�i�z�݋��v(&r˔�I���z�j7vU ɐ��u�ZNؿ�P�y*����jV��KvCD�b����w��Lkin!�n��6t�h=ڏ���>�����o���]��N���Wy'�[3{;K�<��Z�Lyo5�ݳ8�8���Z�t�9YF�u�w��}s@SPwy)���a���EU0�7��A�e-ܗ�4�ݖ�R��{tu7	�2�e�[N��+B�n�ҭ�[�����R�y��k+o.��f'7ɵ��}�Kz����v�c��o�-�ss��5̘�}{|�� ����h�=���Fݞ;׃+�"gl�!�%U������}(�R�\�w_
y��u2:���.�]�vmUc�{�-��a�J���e��u�*�;�r�Ttqv�P�n����[Z4�v�)̋����|�D��(�׃���G���VV��5YK����x�7[��N��6�A�ܸI��]�:òuV�{�W7�D�=���r�-���}:�wV�E����|:�k��F����vl0��ǚ�q᭳���,����[��/��V��[����b��֚Z7��3����-���B�[�j�=,􀷺��w]��mlΏo�����M���!́�ҍf�޼��f<�z�}�#���底ب[|w�=� v�N���vP)�6��a�)��
Z��*�۽�γ*]^��]�nt�xl��^�&Kc��#6�WY�;
����LM���[�(X�xF�����d����	�E��w'^Sz&4�XҬ�{���%�̑��Q"^a0�6��Ud�1����+v���P���Nʢ�g���]K
պdf��1�j�	N��!)y�����;5lj����]�n���3Z���y�+1R�냖hK39\Һ�c]����t�2t��n�ʴr���g*�BH��rѤ��wU�F��֢{�F�͈vc�_wm�Z�yإ`Y3N���&�t��</�T6�gG�X�଺�������[�ΰ��`ԕ�U�uᭂ��G��:i�A"�835�U�5c���i��m-R�6v]���F
��ei9�k�Wь.h���+�����'c4�0���[�i�u��A*���?F)�܀���s�C_A��s:s�q�Д�ʮ����H��:�UE9�5\;}�T»mc=�C֡/�����\�+�Q�v�]>��<�դ����vL�X/���ٳf��)��v�.����o4�V�ڧڨ�k��2%J�:R�c�b��&��m){�l���]oen�Y�֐p�F���*Z�SG�.W*١���n�pt5�;n���q�GMoPʦ��Tʮܾ����[Z��ڬ��X��5��u3�e0�|h�e`K��p��ܘp�+�tK��wY[w�fjQ)r���v)KgMl�
���0�7 e�[�&�J�oD��ޢ�����ͪ�mf�������n2]V�������5`e�0�MT���}��<�ڬbYB�/�l�c>���+w:�S.�WVPYV�o��g$y����m�{h�]��W7�:�S:i���A�+�!��Jf!|�ūc8e�y���ۭu�����e������ovAV/t�A��]�<�����b�z����<�gs=�Ȓ�B�2���B�`ÌS�mZ�B��T��W���E�]F	w9�q<kn�6�Lr�Jf�fu�1�z~��oQ�D��bde��m�)�&�-�a�-�Kчp:9�Z��+"4u>�caui��n�4�v�y|V��hJ䬩s�Ḍ�bޭ�WT��\��B�n-��E�-�w�m�W�.e��X0�������nn���N%�T���w��;m��/���b�c�%�e�/>�Iv��MJZ���!Z��ͩڮ��ұgUq��h7�q��v� �A)خ�kx��ܚ�D%��:bU��R��eZ�Ov��*�nsӄ5����2f�tɉ�ҹv�0��Sz<�k7ilxp�]YX�TM87�rT��H�ܩI�Wگ9mTl��C\"F:�,�f��;.�M�Ixs�-=1�mY�}8�5x��/�mي\�̋ӷ�v,�'�o���8�f�j�e��w�[Tqd�UN�T�N��2C�KTkw%�6\u�Ċ�S�����v�����;|�F������xc*^oPqw
�ThB�h���z�wg:U��Zh��*��Ra�gpc�ܫ�h����Ѥ/f�W�;�As5���`9V�1�e�;�ъ�vf\+[�t���u�*�t�5�,Jnw7ʫʾ7��Jz�����a���x��z�i�,�ts���\��ܭ���zۼ�*�e�d;��0Q��=���+��]v*4��u�s�v��霥��j&����b��}1]�d�lج�ʕ����ʲ8�Ӫ��uG!TF��0ʊ�z�5�a˗��u*�+��䌕'b3�>�DVf=�GMº�&m�uw���g3'�Ϟ���Fq�Ѷ]�XKZn�ռ���`�!z��gu�{��9�ݻ��X��T�(wl(w�G�]د����¥(qd��짡��B���l8�;*Z}s1Ξye����z�C��ut�v���:���g����YE�)"Fͽ�D����B�]���{s�]o7v����9�(A���M�^O�����ɠ��m*�Ox1N��g^C9;��{�4V��Py'.'�j�Y�fUf��\�_f�ŗw�������,�JÛ��>�ËR�fG��:ly�3+�S�����zu�q=�뺣+J�V`�S��BK2��_P�X��ξ�z��f�n���rJٿR.�^�7�r���*ũ��ӰM�k�Y�uaJ国�Io�J�Jc��w�C{�mN�G%
r�^�:N�b�ܠ��Um.ʦM!��D3���}5ඐS�Y/s@�b����-��Jb0rʻ����_.Z�+�DV�J��*v�oU���k?T̾�f�u��W�7�K�j��hQ�x.�R޶�д˛gt�%T��]�wxm�ю�;WO������d��A��f���a������A5�Jݲw��p[n��}]6��u���rU��6�tO�m�qU�Cxae��BV����ڻ��٩�Xt)^���`�`�s����Z�'Y�9C=-�X@�d\��2� 5]Y�j���y[)ª�_v�wΌ���ʤ�8�k$#�w�}�'6����G~��u=�gc�o�꤬��;:,�!�x^�f��̻�˘C�۹���9�N��n�*Tb�yS��.iu�ޱ �m>��Yz�g釻OU�!}o��ͮr�K=�wK(�h���u��ݚv��bWc�]:�/qC��:�.�ke�J�����U��'��pZ&��2��3ƳH�}��_<�oe,���[\j���/r�m�W]�QUǹ�ķ��t��y�M������U���h�J�N�eZ���}�!ڨ����G%�>J�l3�3�����s���r����Cq�q�v�p�\�b�^�\4Y/�G���5��Y"��'7�2VC��rخ�&wh,_s�ˁ���u�yh��++lm�mQ��ʹ�ۯ�\������&Q�o�r2=�ct�ʴ���{�v�}�h]�ǵ�n�wb3��ɷ9Ȯ�8��n��Ӭv�ê��t����X�c�2G�G�|�iT6�s�=�,�Y�;�����[f76�%A�����ԏ]��xpU�-f'�MQ9q���r���9jwݵW!���o{6�-UU�}�2-z�-����z;���@�]���Θ6e`���٩��X��M��C�U�{���YB�VR�E��I��Lr���XNVoٶ,k[�(�@��%�CE�ʴ�]��sm^��6�B-�o<y�2t�]���ɲa?ew Β+����_#�y���C[��ab������������f���Xe
��w::GV���+X�Ι&��oJy��řyt�Ύygj���v�Β%o�C��R�%�w�����ʣ�S��y�Δ8&�ڨyW��&؝�+;o5MT+�:���E[�;o�PH:��nա���؞�R�U�S^((ˉN����.��x��ْ�*����c�c/F�Zf�k�{���v�#v�˵0�>kR�%A��U�MV	�_��Pv�J�UB���UA�B�;�m�G&��n��K��8R�ZlY�^�*9{4��/QH�v����x�n�2�݇��o2'�ð*�9c	��n�UT��6�\Q>�F.��Ҷ��w��ea�ȶ�'2P��^p{/i�ۃ����뾮��1��s3#������yۋ�}Ίᢔ��y�;Z&p͙�'a���UJ�9[yS),�����\���;v���`���GZ�4�������i����]��:���
��c���S�Av
�Y�Zu�&ӕHҗs���4ݹ����v�u��5�W]�V"�t��P��,G�%i�*Ɵ��?5Hr���7��&����w-�;��k^��h��#fHvȩ�zv7����:���b���z��G�S>���r�qQeR���3kJ�v�WB\�m���ct[5��X*r�d��D���:�Dd�(�f��ֳܰ�:~m��[�f�2��n�n����5Gq�[0ɕ�Ջ���7]��HKib�\�U���Ψ�k-��#hWS�v��Yv5��޾�G�����D(Ji2��=w���G���꾶n�9�|9g�>��.���6ݾ�=���c5U*��+�/�ij��4+�,fs/U띳�����.c��ufd�gAhϨ�&uCF���q�/`: �yk!Ϧ��4Ѣ.��Q-Zf%Uۚ���a;w^���6�wk��������;f\�2�89�AV�vͳo�s����ݹz��Y�s��}�˯���7��Y�)��i{4ǼdZ�u�$�5q
��yB*L;t�X�1�ϛ�X)��Ǽ��KKj����G��P�냙9�LΣ��Eݠ�h��ܫ�'�v5�p��Ļ�ڜ�젺L�;����TЯ������<��X��	�ٮ����XvS�u�I%\˖l����y{��^/FF.�۽M۬��B�w.jn]�$w���3+(����p�O4a���7�F������Y�uJz5���]Y\����:hUH���I�mn��T/oFZH�E5)�ȯ��(n1f�VޚN`��iu�����uU+:<��th���8^��XET˙���0b���F�y����{�X�=L^���-�U�ȍ�G�˥�n��4�N��^_^��N�v$����h,�_��!u�R�Y�+�������AXn�H�ob��l&�n��B��Ywbeft��ύ�'nu�u�Y��Χn%ق�⻭j�Wf?���+��F���$w:�iһ�҃����3���t��]��7��J����k{y�+{/��]�N72��o_v�{f¶��i$���k]��;��f����s}%���n��w!�cI!b\��L�J�=Y��n<�;�Y}/W���j�u��)�Y{�z歍e�Vʏ��z�U��9f�<��{�$B�l����	��M��c����]_Z����a�5Ӆ��8\Ps+��J��ø�N��U�b/v�8�v�����[Wk�0�{8���M2�zrqvsy[����� >ݤ�I��~�ӵ�vڽ�M
Z0=Q�d��j����l.2{Jv��CT`�[���#���Q�G�I�"3[�9m&��=r���Nb1j���d����6�p��=��3
r�%p���_(@2�.��@��v� _�w�e��/>��@n�5]d�v�7��ѽx9r�N��ٞ�vZŰE�r]W���qGa�aveJQ�ͅ�f�ұ����T��4sE�#���gt��`Uۧ��u��Cn��SN+�'�@T78Ƃ|�۞n��',c�����c�!9b��t������ã��*Z�f��]��Ϯ����^��uÈv�ۤ7A�Ƹ�m�ں��\S�j��nR�g������ֻZu�pn����ht�������7���R=�2���ad^�K1ٹr��bD�/:$tڄ�����m))kK�ka���칙�cש�n�S�z�Fs�[-Xx*��5��/R��Ѹ�:���❽]Y�sv���q�-m������i�vx���.�jz㷮��h�;&�MGe�f���&��,c,-p�����]˛��:b�b$�щ�@l�L���g�=[]�1`�vO����wl粒���m�nz*އ	i�]��clS��Rd���6e���kl�����J�"v�'E϶�β�;�8��iF��E��h�j�;�N�۴x����S���+
Ok+�b�u�l�Z���W&Y��B�F���h�N��u���q�6��.bMp�5����r]��b�FHl˚��s` �H�+v�y,%u/]�N.�Yfu�4,hH�F¤��ͽ��n%��<a���,���h�Cܝf�*;Mn̘�Vl��v��2]S`�9�+:��p��ў���q��ݞ:�{[r24mF�l=9��Z�F\c����犳����F�7����3R\ywj�s��l�È!v�0T]q�$2�4�-�f�M�� �Z��$Ѓ�@lʨnB7Yw��K�M�]����-���	)�.2v�G���Z��\�.n�.1�Մ��KC�p�p.�$�c�3��]���;.1QDO(㫈��Ҕ����SUH��čT�_�-c��h� ��pf�tFbhr\�p�d��7�,�ef�ݹ�Aݛ,�
��krXeC��A�sjں#���ͭ��s�J����	]ku<@?��?�c���k�7��c�YU�v��г<՛�[Vć����1�g���3ۖ�y����"���q�6ȀͤMNu��=�M��׵�`�t&�7\�ݰ�k&4��6�k��h�Qa�d��k���U{��Giۮ�g`�s;J\;x(6�K�������5:�s��b�Qv<���Bkn�V��Юn7&3[��Y.�C�u�y��ݺ�/ �2q�j��n�39�9�vn ��`�����^ɻ�3�������k-�vz���`1������ի��7���Up���2��q��so�6s�2�f��� 0)Z��_&�F4c)��,W���}/��\g���;=�[�	�z�)-q>t�n��6A�U��4���XK\�0�r2�+1Te���6\u���R$��X���jumQ���p�z��3lT�Q�1��JDҐ�J6�a�.L��ͭ�WSv�jE���g�ǰcm�ݱ��Zy�Ƿ����j��7��&]�����uW����e:��qu����`��V"z�ީ=c���[��������/=]�C]`t�/��lr��c �;L���`[�[l^����uNמ�n����Q.Av��vn�YG%��R9]�x ˍ�(��2٦��C��Zc��pny:Ӑ�r� bi��U(�4ۈ:K3PH�]v�"a�wf�7�$�F�;G\��k��&��-)3XE6.�l�.;e8�+Lhy6G[=6����_=�8���E��Ҭ�Z�G7���x�и��֡͘���#Cj6�18il��4m�����v��C9�nxc�5�F�v���y4v�;Ki�������#O<B�8ہ\n�S�n��e
a�keV(٩R�n9�v�S
O�9n��'d2���Ln\+�{hM<Ir��6�y�����d��+�ۜ6�{b-��{sne�;mtv-P�<g'җl�.�z��۠�:����Hj�4���=�Lт�yu����z�NE��m�sj��V�����O3n�����|f;�qv�,kb���bR�ڳb+����m�q��՝8�Pr���0� [b�8���,�0Xj8�*b����B���1w5pBH�fV�i�Ʊn��iT��f{j@Hkf��&X\���%t]��-��9���^ۭ.��RN���g�Ş�{]1�4ٮޭWWB.��ۮ�%e�lh2�˫�J�MfŨ�2��.ӹ���<�C�9���'<pu� d���\8�j#2XJZu�ؖݩ�!c��v9.q�e�	.�i9�5\�g��V��J�0<�K�=�9�."����ʎ�<�k��rSg;FK\�C@й�y�][ݗ��^�t�t@e.N-Q�c���х07E�vk�v�N�M�\����{n��������xȩZ=v�Ĩ�I�\�4���/RfnJ�MX��n��-�����L9ö�lvۢ$�%v�^[7i�-ԓ�˱�:�ikW�E�fut�ѯn+j�:����d s�tp�0xo�������k�u�--Ʀm�$o&��!��EKp[M�9\�/���]�.xl.��N� Ͳ�ף�h,�;�83Ca�85未�0Ƭ�(LM	,n�I�!ؚ7b�W'nx�m�y
�	��q�u����1�M5$u+D�T]���gJ�s馔,ʻ+lNf�6[vl2b��殖�k���aibSH8��E��[��Avd�!b:T�����ۉj��H�"� g�@�Q�|��p4�v�c7F6�m���K�)Q`�鲌�2�:��;���0�[>�z��}���M��n���5��͗u�	�İ�%,Wc�{F�u�ޡ���Մ{"7��aݍjkN�"���\�^��� )�x��Ȇ��,�M��̀�%{
��i��i/t���y�N�(t��5�P�[-��\�=�����_lUk�q�u�����h՗F��iAna��mU��V �1�;ڞ�ٸ,co�ؠ��[��Z涫:�@�і/%��ə����s���xv��"�;_WFz3ewǙ���̷�d��σ)�Q�dCj�^&HJ�M�X�:�ꫀ�����E0)�iS,s���e�k0GM*���q�Dr�d��mV�۟K�����m�pK��etr�eH��\[f�6�++Z�*���-t�⫳0]�w,[<w9��^A��{�pXS��&r�Ir�Q݆��۔+�k���K<��s�f�u�;$����n	�.+� �`śs<vڳJK������q�yB��7``��6]��W2�Z0��
Ŗ-�epS�)�����m0����k�Z2ꮂ6�*�g�F9��vԡpC,�S8��Į����/c�%mǝb�P)�ƉZ,�ܜh�h�]����Yw�}����}����	��ɝv�W&1�FkibX�B�M3���\�kd���\��������ƀ��DuMՖ��U6���F�gdPT��@�[���x\V��ꗣ�a�v��R��M��Ku��3�XvȺim�1��1:��8��Y�]u�Oi��l5�H��͂�R˄6"�j{:�����-]��`��%�Ξ��1���O$vVn�\n�7�;6V��m�S���c���q�f�[�FC�x�SD�ާ�ӵ��p �/a6�=�ٵU�8����������Ġ�3l�7"�ϓ��Zs�n, ���g�!>�Z����=��0n.r�����&�U�v�X꺓��O�6	�`�B(���t�ޓ��a޹�u���/]�.�jknl��b�����Ħ{%�'eSif�lK���5qΕ�!�Ln����m�{,�m������Vٟ'Fm��ͫ�.y��ϖt�6�%�جT�@���Ռ�.&g�=z��zf��I��l������n�3��ą GEc7iC#4��E0MK�+.w�HT���<C1�����<n.�j�����A�p۳�H�uFNycf���=�4*��.il��mϴumƎ@K�[�;����@�v�BGp3mGZ�F˕�S@-��2�����e��Ò6��`��xh�P۫��q�9��[�]�p�c`λq�u�u��κ�׵ �J�j�F7�NǹcD�c�"�CZ987]�У������j��o#�e�م���&׃i�t`5Qb�5����T��s��fŢ�XݑW�#�fźe�u��č�)n�lg�m�k�n�=�f�Ȇ.�5��/�8�s=rw�\b�u�S�gz��#�=xw��kBk�lЁ,e�JSYq5�,�H0�4YJE���*�'�;�uwoט-�C�4@�z�*]	�ز�1�̥�M��&�噵�Xbf5�+Z�ېQ쩏m\rv�@��:��ne�Չ���vY��p��l%=�c�|x�X[a����Qp���n���ԑv��eHK�»�]6Gil�����X������T#`fm���&��Dᜥj8�6�z�m�Ͱ��zD�c�Ԯ���	eXkW;f5&(4���=q1�m:i��j%��Y��,����C#2q��di��	n�6nU��ie�n+��{;R��Y��Y�5�\�{+[N�㫝۶�Ap��M`P�=m���N��S����s��`�C�����1ܿq��*5қ:��6fZ�u�����(��ʇ;b�4]�aP�O:.s�GN���9�EƖ���tr�s��S�l$��%N�1�X�RZ�(�n���\�V��	卶�
���x��*��Xɒ�i��u:i*�˼p�«36F �,�����8�$q�t�	�s��9��DI��8�\GDD�D#�I��P�9 TtNP�GGD�n���I�$@�D9 ���K�N��NE(��Nq)m��$�H�:'!9�Q������K1DBt�"�%A�D�!�Hs��	B�p�t�:��rAr@��DtP�B;�s�t�"��89:t�q�P8��:S�8� �Em�'�'r�;�p��t)��Y8:99'(���A�s����rN9��q
A�'��A''��8 :\��(9Jx������رƽ$�ZQ�q6�ǔ}c���m��vۡ�<�،�\A<&�K�X�<m,�����)�Ҭ�� �/Xݱ�F�.69튚����1��R�E^�y�$[��v�m�%��]j�;]��s��Av�{/!� ��'Z��s�\t�Kڱ]�vG��)�5�Հ	\j��c�`��*�e���`es�F���գ��[��Ԣ�h3Bm��K��X�mۉK�v��/4b��7�l��UH�,kZ��6�T�p�̓s�s��pv_��f@�H����7K�\�v��^9)5&5#��0Nk�[Y��)[�9���W
<�0V�C/+C��!��mae�je�݈�$�fJQRC��R������_ps�5m�iny{�������j^k�a,�xl�]3��Q�l=�ڌ<tn"��9�TV��)�m���a6�Q�^!�^��D���z ��ї��A��;]$�23m��H�F���aK6<[p�m��L�j�2�7g��K��1���<�8���%�c$[��`э�e�U�ݐy�/A��Rq�C��CoJvn�S��^SI�"����7sr��u;�6ND�G#���p״�RX�ڎ�#!8���:�t&��LT��,uń����1�xy3m��[x[��`Yy�P��.&nJ���n"u³��S��Z���7�N��8�qɒp��b��<{k�y��<;qqY9Ӻ���={nm�<�f�����9o\r�ΣnU�!�5�Ξ��7�s�ƺ.j<�u���`�f��v����*Ѷ!we]u�&�wc�`���ls}�����Ӯ��N����uT��l��塀�ո�!����2��]�W�͋�M�ȱօ�q�e�Tf�]�te�aoaa�5к��e�;cR�qr����m���$Fi�hu,K
��SZCf\bm+�-p��5�W��&5lt��neĹ�I$�]���E(P�x,)[l���`S���/XY�ݥ��J�V4�J��Ye�1)���B/[[
��^��r�,��ԱaH�V�R�D��bJ�W�)%Z�R#Z��i�l��`����ć,Z�:��EI+Q��޴��̵�F�m������,���O�������裋�K��j�A�`�g�Ĝ���t���9qaei`�����H���2����K\��k�֯s`�k��_��PBt�������l��?6��@�B*��o5���WȆ�7y��ճݰ):�*y��렁n���b�]�h ����W���~m|�-�Z��׽��%3��L�znp�민D��"4n� ��"H>��1��!2�9�=)|A���W��{_{\X�����>t�~��r=�冶���}�A [����mn�mK�X���z>��6;�m�'��҂�����D7CX���M�>�F�ī�(/��$:�8�q�1m�M�V��ic.�Y	���tS�d��7�D���_/�m2�y���#��r����B��%+�e�	�$���HA�!��@x�WO{p�dʺ��{�s�z�=�����U���OP����|{�t��Q����an���^�&�O�(?gxW��}R���Hg�_W��[��/�Ŏ��]�_'�#�x,,^��,O*��j��P��H��H��n�_�_o�u�ܯK�ʡs6oud�Ǧ�x�΂ ���-�!��A8�ugU}����6�Ǔ���<�}�]s+����g��˷{�qc���@����%��t-�J×^'��u��y\��y��IX���k���������6��:Ϥ��ߎ�H�7Uj���UMv��;Y���׶f���M�&9��ū6�̕o��YҾC���"	�v�wN�������"O3^�˼�I�֭L�d2�;���͠�-���U�~�(*�ތ���"~܁9~שn�x[b�ng�A�$����n�S�����0@#.��저?7A������;����0t������|Ȳ�N7٬^r��ӈBS�qq�}��e�����͡t�]��b�Į�(!tkw	�B�,�>�ur_v�%cO�}����_'�#�u���-�t`��m��AmY���H�n���ϸ��ZD���'7p�G�C�_ ���tźD�@��ޅ��7��ܹ	k֞k܏l,m��z4~%HY!|[�?�"��}�ŇhV����h��� �3dR�LX��	ǰs�uX�i���:�4��9� �vP@�Hh/����<��~�"|;�~C�R�kƭz��?{��mu�!�@�^�r�2߽T�h:��=�U%��Y��S����>� ��n�MDQ����>Ȃ?MHc�*�g9e���q�,�N�9��{�v��{4�p�;�Ǖ�AIHcA�u�t"��a�����tr�M����-���o�d�þ���<�\���;�m���a'u��^H�c"�XX)7}ou;�m���Md؏�b�ntp^[����Z�;v8�S)5j��طkRC�����n�_�|�h [�[����Q_g�]җ���J��r���:y�>�et�!�2��V){���7x4"����#�D�.h�:�2��E�E+���:ذ�j��Z<ǿ_��nm"�_�@/�m����~��h��#��׈�<����W�A!�^ �_ԁ����t����oH����H����t�No%�r��_������'וXrn�9 �ܤA#�|�A��&�U�Ny�~�o��.ǚGO A��� 젋t�-��ͤ;�n��2y�`��W����|~m�廚�}��8O+�A!dH?"7��=g��?�_7��n���[��uw��z�b�ȑ�5���U�'�מ_s��#�i|~m�(�V�z��x��ى֋���G�iϚ�}�5�:��ᮙ�wϞ@��f�}c����Uf�%Fs_Fl�"��m��:۬xK�r��mΝ-O:�R�=Z�Ő��ج,��]���&��ܳ�t�]n��q�4�����˨��ƺqIv�z��Vnq���P7^3eѮ(j! fU
\�f�س[���XQ-ͬc�<6�x�8C�'-��=��t�l��V�.Cmus��t��r�웲������ ��(�&Kt5s��h[�t�R?O�����%���i�S�6=n<n�sԽ�Eex\�3��vKp˦͔[]���oc,�?/���ײ{�C���eu�:W��z��X�Y�,A�_t� ���� An�?xT��\.��.��������s�������9>v���:D��L������Èۤ�AzW����dІ��L7ދM����������\/�}��y��� ��������׬�8��T�����F:DCt��:>��kYP��kd��E+��vȬ�)P��ޤ;��� �H����#7g��1G��}���v^�[��������H�� [���z�Xg��>G�y�%#��]\X		��dSs����U�s�ѻ� ;�e�җO�ǿ|#/~�F��"��J�=�����\/�}���c}�𶻎{c�M���r_7_7Y����-�W�#��{�W�Ӫ��w���nw�Z�3�>٨<5H_(��D�Ud��H�ض�ڧ�wU�{vs�����C�Ն�����:R�N���G���m�:y���쯛����.�G�����җ�7_�/��}�P�E���[�p��]=�H�H��K�	�!���b[�����A7( g�����������u+��x/���v3�/��g����>_7XA���k��ۛlm�f�"� "�ىn\+�wH��h:�	�	8����w��������
�ՂR$S�\s8�9�qq��I�Ͱi���4&,��[��_}��� C����� �����ʯ>�%��{^"�x�F6�A��=+���!��-�D7��X��J�H���_����ܞf��{�@�Α>A�t5/C�+��T'Ƕ� ���6�n�	�p,Z�y�������xhǽ��Q罵�uc��ẕ��lIR��B;×�[�}U�!"ӊ���T���)-�y�����u��\��U7���^0�wt�kd��A7+�����?6�_I����=�G�s�t�r����h'�����o������h �Ă3u�na�m*�^���n��6��"	n���ͮ�o��/�+�7��ܞf��{�Η���� �!�
�{�1�k��joX��
�f���q\�21�]�&vF��&��vv�h�sƺ�P%�I�����~�n���-5���û�C[�s�x��̣M3����{+�u����At�#�F�h�t�8�_�=v{�!7��v�&��6� �����{��"D�MG�/W�|��|u�@�_ ��o/}c�}}/wdn�=Ϊ.����	�H_ ������n��{�d���W8��������H��~��_9Z�{|GO O�F��r��_n�+E��p�9<+�P�0�� �c��xѫZ:bN]�T���s�֍k�O�s�+x���ٻxݙw�6��n��H|�G�i�n��G�י�~��V(O��c3���t%o������x�D#A�|A7Hpu���~	}��LYtҶ��a4ٱ��v)�(�|�j'l=Z���s1(�K�vX��h�G͢��)[C�K��sw���b�{�t(����-=�h � �ϒ���@�H�Ct���坩n�	y��>��z�>�䩥����̆���'�j��E��~�l)��ju�!��7���{�_��t����K�z( v�r��u��i A��t�������7BA�A)}��Q+���o7sÄ]}��y�#K���������W���mt�$7HCk��'P��^��>���"�'��{^:�F�S������?j�������B��+�K��p�7��Y�5R��Jn�e�uU��lb�V�9�^�������e��/{,F�X4�������3׋>�Y�ޚ7�/��<h�Ij4)��ǳ.���y���t;�:��w��=;�xwm���f���lBa�Y(����x�ck�p��1��r��/A9��h��&����:ڀ�Fk\��ښm�q�'	��u�jn1i��0��A�$EӸ^ӎ��w��ܜ�tnr.r�O�8�P�:f��3��%y�Xah[���6����~O9a���D_��]s�ͺ�nQp��3�E����ƬP��غ�r��й�i��c9˸�rϷ�y�Z��{�s�M׈���Z�k��ޡ���_�"H�t��-b��Z�l�>;ԁrrW��7����.�o�y��+��y����' ��DD��-���F���z�ޱ��Z�n�Q�i�j��k~�N�&�	�㎑6�?6�W��:�.U\A�9��_7Azt}�A�g�'<��xA
�A尃J�n.�C�ȑ�ۉ��E��n�|[�� ��"�Isi�F��T�6�{��o73��\'}����H���o���^d��\�i&� V讛��<A���8��j,��l���(�v�ð��z�d^����n���5��r�����~d5�H��+ʪ=�� �j������� �_?E�v����n;��x�yR�R�6ګ�η�D��"j��]>��b]��V���o$ˢ��6L=bo��V�F��nb�4<��Һ~�3�͑)5�T���K|��)F�A� �#A�6�&exI n�o @�t-�@�H@m몡������׏�������%p}�? '�/�;@��|�h"�/�sjPѣe}�Cr�@� ׳=������]78��}(!��<B�u:����?6��~m���v�������@I�mK]�֢ݸ�A[�A��n����⏆/t<=��}�����m]]
\���1�Pܬ\Z켾��5��ڍ�5f�Ri�'ο>2_�H����h!�<~�x�w�J��?+��ֽL碪����@��ŵ�u��n��ci�wvsY�@�"�ORjf{��M���]q<ޔ㲾n��6�7���@�~�H�"k��}���Oo
����[l.����A9q�][��zD&=wjV�ì�9�ݭ�\gfFXCJ�|��:D�9�C��Yu��;���P�a�;��gE;����ůV�M���H��{F��Y�Z��%}�gu���P5�G^n]��s&+'�"ڬ�� �q�[\�Q���Z���e��J[��)��G��.���Y�üT�+]���d]]k8f<�ӧ�0[]Ɓ,i�YQh3�^mlt3Vgݗ��]c�J�o��L��
�s�:�0)t���Ђ���b=Y���{AeT(Ҵ몕
�ˆ��]�p�뻺�u[��H=������t���)�:�\�lF}�-ߏe)�:�t2Rc]V8�YB�h�������ɻ|+�j��=�]u�컛X�o]�p�WR��4;{�vcmԻn������bf<��w�B��Z���S9m7e����gx3P��y�D;�z���u�y�����:�[������ȹfCSx@լ	�r��󶅼J�zF;�]h�lh{f���p���R�y6'+W^Y�7�Eѹ��Cs)��ۨ7vTn�A7��L�}�I�u[�-�Rƪ���3+�%�pyٺ�`2"*��b�˭��Tx������:��W�w�)ԛ�:\Uz8d�dڻA:��1�r�����L.��e�J�[[H�;�Tk��f!iVj/k�V�r��U��rӚoi�3�jX��S��ȊI�N[�{����{)��-����ӽkU^���"�Vmd�ͱ��(�r�-[t�IJ�۪�f�"�v뺵�����V��].��֚�'@�����ϟ[��9��#�D�,t�Q�D��	)�q��B�8JQJ����q8�2��d�mͬ�w "QP��0�\N$D��nt$p�%9ӝ �qrRkb(�!':8����q;4+7NrN�����(��@�8�9�I�
qm�-�' DG@*w $8���@#�:D	�'(�t9	ܐ�"BQ:��$Nr�D"�9�YB�6��9�������و�l����խkrrTAT���P�C�������{]��;�`~@�h��) ��J_;p-��XWv� �n�i<) �S)wn�bRAa�A�q �3������ׇzݢ��B�U���S)��P�`�I@��(G���mW�y>��z���=H+��|�
J��B�22� ��o\G������q~�
��2�)�6�i� n�i��YL����Ĕ�XPn�1 ����E����u�8�%FR�n�a��������y��+����I����q �*U�h������\�@��� Sڅ���
��Xe�k�?yW}����|��E���=s�8/l�v+W6�K���a�p�\��kC/-��|�W�X}�RTB�~��l��H(o�bA`cIwneRچ$;���~��(6��oֻ�<@`I@G����v����<;'�\CĔ�XW�\1 ���R'�)wn�`��Xn�- �0�v�H8Q
H-��WϽ3�ʿ9�a���
u�o�f��P�=��H,=��w���g�~�ώ���a�A_6���RP�0�jɑ��P9�- �1�����GO�����|s�����- �0)���
H)~��Z��
��H,1� n�i2!I��R��@��{�߾�~_���?nr��zm���$���
B����- ��������Xn�-��Iv�H,0aIwl1�$�s����|���-�q�6�l�I�>��
�끙D�>	G�_=ַ��(6��/ֻ�,���i �ᒗ��C��_���OS���F]�)�-\��{!,���o	�[[Yo��/4��D��'5sxz��3;+�ˮ�u̲e�U�����m��˼}DS�L/�c�_�G��
{E����N�P-���v�H)

�7h�������H)��v�lHO=�?��ߣ��|3�/�}��]����e�x@�~ t� �yA,a͸BМ�@�Br�+����/w�_����0�7]�]N�m�`�m����B%X���-Hk��X���u�@��i��I�)�j��) ��ݸbAa�� n�i1
H,��wj�ff�����>���o��RAa�h>�$�9��8new���^>��Qi���^�@���)���- �2!�F$��]��
Aa�P���P>��w�y�����7ºx�X�${P0�G������Qk�իy�҂���������O�) ���C��XWv��)v�I�^W~/|�ٞ_�q�~H,��sj�`��Xy�B�
C�m�rQ
H-n�H)��v�l�JH(T@����'�Z���>�'^�X��?��w�x�����ͨ�R�l������i��$v�ZAH9*�H.0)v�L@����~ߚ���������N>�@���Xg�pĂ�#
@��i �c)ݨ�U-{�s�o���y��>�5��I!���h����RAs��շ��{����Ă����j̌��P����aIݨ�Rb�v�l�2�
혐X4�]ځ�~�=ﯖv��� ��̨b|	�ɭ�ڥG�m�ݮ� �$�����ʌ��ځi ��ݸbAH(�ZO �$JN�@��2y���&
����U7츜G�Sp^�w�f������Ae�4��T:�͚�^�������V(�uN��.��5Z��x�4���|�:l��������,R�[A��@*�RfmEa2�	s+�Vj!�Q���ֽ�8x`�����%�d���G�����ݛ��1/��:�Q������ʌ*6��נ��s��;q�{�q$8d�Gt�g3ݣ����1��lj1�luiaz���v�̼�:��F��:���,��	�C)fm��xe]�';a�fű&H�d����Bc8���K�~?���]�CFm�msb˖��;!��(v��v�;1Ք�fYC�3����Ă�P<��H8Q
H-��H)��n�-�2RAB��bAa��{���~���<��m���A^m�ц$�������������|�ߎe���T-�FRA@��ى��I}��ZAH9PݨbAp`R���R
��C��X{οQ�=���l1 ��� o�ZLB�%2�������w;��XI{�D�'�>G���h���D) �\� ZAL
a�P�_��y��Wd� �h{�1 �����ZAH,=څ�h�H(�ZAH)wn�Q#�b>	G��|�ӛ�{;��8��������y�@�}����
A_;p-�) ���pĂ���E��) �S)wn�bRAa�A��AH{_em����}���@�h����Z�=��S
a�j���$ �	#�O¶k�y�Uww����z�W�a�H))
a�jɑ��P=Ӿ�~���LH,cI~��ZAH9*���� n�i�$Td�ݸ�R7n�XdaH�ZM�;Ɗ����w�B����KS�@U���s�o����w�{A��AHQT��i�RAjW=��S)��B�
AC7hĂ�߯�|���>yo�����{�?r��]hQ֘��:&u���sm��Yl�F����ӋSs��0M�7�FΖ�ߞ������
a�*Ƀ) �T��bA`di ����(��Xn�- �}�����^�i��~]�@`I@G����g�{�;%/9p-�) ����aH��I�RAH+�p-��H)
*�ݢ�>G���=���2�0�rF���ޏJ�΍#l$�~�t�mm��Q�k�R�A-@�����e!�2W؝�ة���{7N�߫��N�#��J�������@����R��ZAH(s�p(��?
���^o�U��9/|4��yہi'�
a�jɃ) �V��H,i �����xUe����/��¡�H.0)�Qi�$Td��n���v��0��-&!I��K�p,�#B����+�����o�8����,=�É!AT�Qi
!I��܁i0@��f2RA@ݢ�aIwl0a�#}|�=�ʽ慰�ꅲ~I���
���̢
A���PĂh=Z���^�iߒ�.� �$�I��K��
Aa���i�ʻ���������i:!I��R��@�) �ݠ�
A@ݢ�
AH.��- ��c����H�0C��Ă�'���{߷<���<�=��=H+��|0Ă��
a�j�R
��H) ����� �*�H/����;Q=[1Y�5�c[Il"ٹ�G3�n׫��cv��<��z��۫��<����OD
H,��K���
Aa�}�bAa�7h���$JK�p-37����]�dsGy��>�7`��>�m�߿/����~��?]�{D) �\�@���Xwj�) �Q�1 ����0Ă�Xn�- �_��r����U��|���I}��ZAH9PݨbA~�}�=>��﫻��w��� o�ZAH,�){p-RAaݨZAa�
@ݢ�_��Ow��KR���Z	I�6�H)
*��ZARAh+w ZAL@��H)�	@�>�=�:����5H�f|ޣ���Wp�2,��YX�b��҇j��E�:��eW���fV1;'q�Z��lFRW8Vw�}��*W������y��=��=H+���R{P���P3{f$4�Wv�`eRڅ�#�7h��
H,�������̸�������H,1� w�ZL�RAd�~�R��� �T������-y��>�A��AHT�勤���RA{��6�����݁i=)��T-�) �@�>�RA]�a� �ݨZAH(nى��Iwnx}�{�~�Ǿ_H)+��>G��o�&:v�s旕w�Y /h��@���){p-II�v�i �n�i<B�%2�u| u�Y�yl�CzH�R���h��v��	�2c'2Wh�\t5���j��uv��\��|�X{t8�R*�ݢ�
AH.W��H)��v�l�JH(G��Q~�]u��{�2s���"
�n����Ϻ����΅���['#) �Q�Y���$�neRڅ� n�i �ݸ�����}E���!��F���-&!I��K���@)uo�_p[o�=G�����$�@}��p��Z+��- � Sڅ����2�|�d� ��~��H,0aI�p��j�;�X�r�_��K�p��?��6u�.�s�/W�"��� [���7_7�-�~���ޮѻ���C~?9_t� �Ar\�9������Ϝ��J��W��Ś)_�롈�:=t��v���inb{QnӖH]�;t�Y̦l�̼Ɉ�"O��,�͓�=�:�LЖ����� ��>g���߬���E9ʲ"s�X�Ow*��Q�Y�0~���S��	ݼ+̆�� �� 렁n�Уz��gP����2[�8�[R�-�[�f�r]�Nóϴ4(�B��:ͫ~vI�K�Y~x��ϋ��2D��x��KNB�J�{o�e����%ՀFu}ΰHn��7A�":�{�sٝz3�7㞤G��ds�ٍ�I���9C���. �ͳc���jC}�U�c�q��X�9e��X�s�O�e�t<
u���}l'wh/2������"� Am������I;�]m@Fe��/�m�o�����\Β������Fu �������s�	�@��@��"	n���R�mW��� �����Now��7�#]�|�|zW�G�����'<;<Vz�1���e���}ث/Fl��|i�?n(�Ai^𾫫�M�65b�w�F�-[ �%q��E�R�����eJ��!$9~���Jj�(�Q��Q���
ݶ ��6��ے��a{����#3C	am���T��ϫp����cO#�zA�6tFG;��m��%x)�Y�ʎ��ۜۇUu�$c� lFZA����;1"����k�+�Czl��4jsֶ�݅,���|r,[�r��7����.0�kn0qqĚ�v]������Vv�#z��5n�v�s%�&�o�~~~<~XiK��8vyջn�Y�QXL6�3�J�R����貚�}�O~��t���-�;=۞�݂o���T^��3�A/(#�R�������[���{^Uy�g���}_-��_o�ĵ:D�oW�$gW˚��Z#\�X�R#�����n��0xY��_��~�����gdq�a9C�JD��_A�4�/N�}�~��g���#�R ��ا�ݹ���2>#��'e�ı�Ρ`�� � �͡���/��@��$_���c|~����1������%)���$g�|A�-� ��f=��mD�?���rFBD�JK���;�,�v�w��v��'��s�v�n��?~��}~$o��|�z��h!�S�����q�iߜ�����K�z;� �A���tn� ��������E�5���n���������:��X�Fb
�e5�bӳo�h�Jc�;�&v���5�*Ǻ>�#ɇ�B�ۓ���=`�������c� �3�fsew[���~�<���D���k����+;��̿x`�_����H�A�h/�͡e�!�D��ɫm�W7����SW�:�A�_7X@n�!���e��W:�r��A=��:���s1�b��c�x�ݛ��'I	�g|o>��W�/��"�"t�n�-�V��obBwI-�ޛ���.͂n���� �tn�M��#�lۣ��!#U�:��Zz�(ͥD�
[�R@ɘ�NY���s�������s�}���|������}���QL}_S��u��H�;P@�R �� m�t?Gy�%�t>޵F�X.R �Dܝ�G�돷��{���\�A���J�ߖ��:��"��t�$7U�Ϋ���x�ݻ6�Y�.��aங�ĬZ�(�Ӻ�Ξl��6㳭�52�+Q��Zr	�&}��̪��uHk�m�K+s�|>����ٽ�����&�P}�rP@���A�|�A�_!$=չ��x53kW���y�/�m�oo>��2Ҝ�k���_b}��b-���A
��դC� Ch/��-�@�X��gW���0o��V%&�zoM��}�~}���@������$g��{(�b��n�Vh��+5��
��-��-�X͌�bW%�B���:� ^R �E�@�Ct�~S���nz]�
��ǲ/۷���v��'�]��\����|~m|��˷�Z;Cj��`�~��'��͑.߭�3Op��W�4H����"�zR�g\�yH�ľn� ��"� !�4��r��泫M�]�齓�����w��HC� ~m/���n���8�����`���ۉ3"D���z��Oւ�p����@�z/N�޵_z�Ħ�v����o�k�3��mݎ���]��p�p�{{7�	I�pz8l38��3/+�m<}���R8)T=��g�W������_~���o>_7H���ݝU����{Y*�U�/�3_~*�̴����}�'�Dn� �� o`H�/�D��&\��B�tٙvV�.tE�5q�+lmnp�G*�V�Պ:�p1��W��|A��'k���3�s����N�Ct���F���8q=[�h ~ւ����Hn���~/l�vWf,w�$�\����W��h+�-�A�$�@����:;����?{@��� ��@��_7@�Y�$`�}�;7���-(7��}^'���t� ��Hu�&x��7c���y_w�-��'}m��3��8�#�N��%"<��Zx��y���ϗ�P@�A�7_7Xu�u��� ��@%�t���ﯳ`��BO9(��H[B��J����5�Tp��YOUp��r����7MT#�����\��b^Z��U�K=k,]<�1_<m)�e�g�+��m�{�yk[�*����wnu>�	O�o<�����ɼ3(���V���E����d��Kx\.��5T�͛l4jPU9N��	�&d�/�2���,�9܏�G�ꊕ*�)vh��R5�en^�ka�e�Us!���������=j�㮩}+T��-�z���{��GhŎ3��fvgf�.��Zr��k2����I�v� �Dgq�<1):-�]��[\̷�����K*My����{�gN�o�*z�*oS��`W��}
�������ꬪ�2X�HYs7`�����.k��d��OH�8(���U����m�X7;��G�]Θz����y��[ޭ���f��S�g��C�Eٴ��M��$S������^|��lj���j�B�JyΏfm�쉊�V�[���:�u�7&:��]�F�Н6�\x�[ �;1��l�hu�yjۖ)b죙���9��e��H>‶OW3]v�)�ޮ���,w��Z��6���,�]U�w��G�x[v�*�u
���Ȭ!p�+ �9a#�V�ڶ�&�_@:�����=*��ͻކ�Em�`Ӻu¡YR�V1d��pY}9�C5���SS�!u�&[͵���<lM�s4�Yk��f��]Ϊ�EC4b�v�R�ݽ���#vb�lI.��o{!Lei�Ί��	+����lKg5.L�/;3s�rh�j��>���1M���V^�Z{�+�f��7]lA�7(*�j�"�#��I�9��m�m�҄[c�vvFZ$�qHm�iв�R�(N�v��m��:J�Y��;�9ma6��vu�kIӹ �GvQ�3���im�f��8��#���b@�����᭶��Esf\չ�$�#��m�6ř�2m��qJrqN���.���$��m�';�)��gn,�8��:N�J:"8�wPuVvM������,�Nr �H:BH+m'r�gXɘ'�3r�*H�&�Y�,���H��i�Z�1E�N2q9�[e!+kY��m��8���s�6��I�y���	t�gLk��`�V����9�4<a��N�OQ`�b�!k��K�0ً��K�޵���vHk�B�%m�k���[��<z����{���8�����=�KS׆\�V�\�D�"m%�Z9��ɫgY�,�<�n3s���M\q^����Av����}�4��ZSg�-��t�Z2�ZToM��2FSGm.o��,�Z%�KB�V��te4�fA�#�m��Ɲ����u���&Dpԡo6���)h��r/���w��u�QV�-eض�er�%gf'"+q�e�Ar�p��Zl����Ŷ#Xm\c%��q�J�ݲ�3d�.�P�/m��>z��?3Q�`�,Y]��Me��$��g��94��\�[�Gu]l$;ӡ���oj�qq���K-j��H�;\I��co�N͓:Õ�\�؃�#ƫ��Y�s1��"�`pD��[c�^^����o3�Z����:ܬI��&�f�u��
�ue�\�y��뮍��g=��cm �+'D9�h�%�I+���a�����tV��t��I�ӨDa�����Jl����; ��$�R`V�����4�s�V�R5(��D`X�b��R��a�1(�6,3r��4� ı^a�wa���eC�d\k�IZ�״�%���<P���qt�RU���5�&���̱ڱb1�X%�Z�si��+\	�	�l�nr��%S��IUrj�*������M٩�uF5��R�「t��/��o9���F��,�3c��'sp:�ct��pGk�6޴��_\���LW1�h�p�j7�jmk2��`1+mQ����"M^]�(sݨݵBN��(�������� ��9���.XH뵪���x^����5���H�^q������#4B�s��Yz���vFZ��[��F�1Ѳ���k���\(��lYvXiln���rB	33i�Ml)�eM�	����n���m�S:�s0�5ΰ̡4k.%]�I�;���P��q�ۀv���{Y�$���X�m�W@k�Fr�i�,��Y[�+�Dp�}���ʛx�n�юrq,3��̸V`�� 5�j%6��];�f9�7UZ�m���l��;g��W9"[����Le���)���-a�H�yֺM0���oO"��ٶ����}�C�=t4��zZ7���C��m:��q!m��5��b^sj��l?O'��_�i��ml��01n�nfZ�ô̡˦5�\D	��GW���[����2�ϋ���6߭�5Op�!^cc�"h�ފ���W ���c�WNr�Nr��(��T,�2�ةN�έ Ȃ��>�yo<�7y�w�@�)|Aq�����_�-W����A���@~m[���7OF�1X��u���׽}���yJ�����H[_�7�gm���a�2�W�g �ͥ�t�f�z��̵0�	�����~��W?T�ΐ!�%��[��n��j���l�B������ys�6f�9��/��C������'�r�B�!oh�䮊�D����=�˷E�lV�:���,NU��9��3o3k����A� G��n����'{{��f�7z�O �����^۪�At�-��?7A [�����U�c��FX�~B]sr=��K�3o9����$]P�櫗�ײ��q���S�M�׭�9O�ḇ��z�`�ԯ��\l>ڵ��t��?��| ����	�t}^o��^Db���q��ԁz �-��1�A����)|Dt��%��K�͠�d*䊕>�TO����sy�����7�ϧx A��N/�x�?6�-���sۓ;�Ա�+�k_{����r�{{�3�f�7z�O/�PDb��ί��> ��������Ch ~o(���G�����sٲu���S�s�s}^ OW��[�׮���(w�t�]�����T^��k\��q��{pg0��K��kz�Y�]���1^�@��|u�E�_\�/�=�1����7�ϧy{���2��:�ń���n\ww&�x"��7�?_�2Ů��*�A8��^^{o[���z���&�� �(#$TS�nR������C����H�?H��D'£�,+�3�6�� w��-8�Qd���6���`5���QN+d[���Q�8�T��8fr��� >��v�L�w���c���[ j�R� %�D�����I�u��B�%c�`�>�=�̘����ٻ��Өx��`��U�z���
���w�9����ۿ��c�-^>�� �y2w���wKP�nKhm��?Q�Jl��R/O������<O���j��i��kK��J�.wiヴ*]�g��\iMvp���tո��te����<�I�)�IP�����t�c]�<ίz�S�*�^�A�ذgR �%"$�IA|B�$p�m����j�>�{�&?oyGo$��o��@�����/��
��^^Y���H�_-�,��|@����ř)$��vVĢ��zN���d���O�A|A/� �}bD�E������']ٕ������f~)*˻[2�������ibH�K; ��hË=a]�o������m7�J��-��jY�!��M�޻�t���pm3RHu,Uf�l�{�{6�pB�w��xF��7�� >���ݯ�7ڸ����E�]�.;�o�s٘�}�R��-��s6oy���7��Ӽ&?+9~�|�	%�Ktշe���������Ya��ꑳy'�qyK�s�l���p��˷6�Z������̎�Y(��J��֧�X��z���A�Z����а~�����%~�	�+��͡���2��F6u\��?]��V�
����յ���a��1Ɛđ�dP)B�cf~ps����'��i�7{E��Ԓ-I@�쭫�����h��>�M���ܑ�F����1�Yr�K�$�,��	��߷
��7�_ؒ		D�&m+�׭9�'��pZ+�p$�D߱�v�W�	��d��"}$W�H�������Q�ٻϐ��빳kkkc#<�a�c���Bؒ5�(�?%L�]��st���U��z�Z(V��f���ݮ��c��Z���?]�+}f<uT�{�K�3�sK�j�4�����Ԉ�������{��{���+����ѫ*���V��l����An����G���-���ay�0R \g�p3�����e�¾�&��o]��9س^b�i�cP�B�X`	��m5W���*�5W6�X�k-�
�a�����Y�����]�r�麷i�t�2�׬��i����W�|�A��F������)�3�N��$ ]���C���[��W�cΦZ�uݢ�����h���W[A2"�;j�K9:k�<$j	pԵ�˪0���`ǜ��.�Swo�f���׍������o��=�n����Y�_�@9����I,_�J�I_VsUJ)O�����_:US�=���uc���>��x�z�E��{e�f�V-]И�@��|'\VA�~��X��~�_��߃����u��#<�e�c�đ�dP)D�A���A	*��Q��X��L�C����r�A��u�o?=�ܛQ��yg��i��YCr���_wD4%/�$IK��ŀd��n�	;�z�W���t�76g_zuc���>��/�P� ���H��"��sk.�=����O��i+�vh!`�k�Մ5`ֹ�b�S4,�e���]\���u���'˾r�'PG��H���:�~�̼�ù���{sS�ϝ�1�d /]
 �A �)$�( C�ի��~w�t��;�++���u���Z����������S�Y�絵w�W)eĝAኸ���zc��_a�8��b�9�NȘ��|>�ߠq��.��潚�7.���>�N�@�=�@���>��=e��/<�>v�9ڴf��ݫJ����}I�x���s��w�9���;���|���\wv�Dݸn�7�j��&"۟��,��})*��m�[[�^p������'��,�ILk��r�~� ��H$�X2PDd���/cx��ݯk��#�My�̽��^���O~@�=�'P@�"_��8�,姭�������v֚�E��l�B����
�v�N�I���h6�6k!�8�}�e�|�s���7_O�BQ1���j�uŤ���mHS�K�C��w( �_����&2E�6O�v;``�|�_}b��}��k|wy���bH?n�
(d�y{�)c/o�|Gw����A��_I�"��?yz��=V��is�m��x�n�35�3mmq�xUQ*�,Χj�Y��1��~z��۟{qm\�����v�|>���L��7���ɱ��>	�s@���Q��J��I���z�z������X3Ծ �D�u��ګ�.�w�p=	�@"cX��I%�P���=��"��#��2��kد_W��b[��z���yÂy�G�o�[B�J>��1.�׃_������*���Y���g	�m �f1�p1�;��ٱ��cef*�tݷ�|���Y/߄e�(#$V?H��vn���=���F�N��c
�]W�N�O�ԉ?=��$�P2Wȉ),�w�xٿ7ʲ�z� ��'��y�~z]���/ ,z(� �_PFH�t�={N� �$	�yX"�I�|d�*�f�ˣ ���y��/y���j>�AN��I��K�t���w���4��&e�_X���ݓ���d{3{M�;���YP�����y�]��r�ke�u3��hqۛrbp��v}B:�}{|����U�f�`ƫ}׋���V{A��g(^5��޿������! ���9��f��(����T(���]L]P��GJ�c������{j:��� ��2EdIA,��0���k���R�yzsk<�nR.,���z�`�ٻ7:%t�td�)����#�	"�G�$�E�+w����6�|��f�ܫ���ޮc�^#�=ɽ�c��wr`���g��W�Yab������ ��ۛ'���d�3{M�{�	n+��' ��:΅_"��}�X��HA��D�ř)(��S�#ͷ~�Q�[���1�Ӟ˭�#�X'e����/����"�	Cef�O�_�c���/��I,_�oѻ���Þl�y��A�� ��CUu��׾������$�Y��d��2E�������绛=ͬ�M�3y��w���W�NA|~��� q4���/�݇f͞�0ō��gbv0�3�?!��k�����׷,�����0I	c7j����R�&zL�6�Oc�&hSP����|>  2{�*UVZ�-WN�8�6y:���7۴�:&Yn�՚6XkKHM�;M�4]a�,�ra�]gn=� �6.l�4q9b���s�pk�U�i%p��Î}�4�㋊!��h�k��hN�)���n�{�/O��)Fa:5��rT�����X�&�P4��2dҺM{n�x;7RIà��\+��M`�n���`�m��r�lrj�+<�,���h��u�q�%�9M���n�+R܌3`mamn��	w!y[_/+��`�H$�+_����F�Niѵc�{V�D���[�� ��_o��~�� �2E��gL����Sч�y|�>~�-�����<��j!�b�3bH#S�_��yEb���d{)�w�����2P@��D�!��������zsk1�ۗ��;�qY� ~��BIb̕�-��9�����UIL�;6Ń=HAR﷟�߇�����7�,���ֱd��3�m�x���\A��G���"�I����T���,W&����;]d�k;\� A?R �����_	*��k���^y߼��~�4�\b���Pvz��ٗ@Ia�k��+΀�+�WM�]?�,���[��d��H���y=���㗜�:��}�[�g���#Z�ޯ��h2R �D���Ӄ���t���P����d��k�ɚ7�nn$��7��m�j:��իK$��^��|�g��X�^u��F�VQ�I������� ��η�n��M�m��Ѫ�t�ڀ���	� "��H��pS[�1�4?kH謂$A|~��RK���|(�~��Z�.�<��K�q��/bAn*�(�!(�T(A��{i��g x�l|ӛ_w�f�sv��rK�>���qX"�������{�%��n;�,MڴMݡ@��v兺0��_�����K�Ӄj�?{ i�	))���}Y�#Y���w��}�b�Q�������Z�n"�2�lxqA���1��t���}r�{y����<�D��S}��^}X�w\�����Aֹ�y�;���mޤ?$���i��?Oa�d�d#+���P����Κ��m��䗼&};��n+ �A�b�r��nK��a��Ա7�h�����Dݮ 㷕��=;��E�U�n>uW{3�U^v5X_�t�7f��_^UGF*2�pou�W�9��<�{N��	�R+tc�j�$j�+Gn�?���S��L"����wx��Ds\4�X�{w[nӲqB���9�c��`Vd#����yuUQe.�\��*��pr�V`�ʷ����t�1Ԫ��Y��g�Uc�T}>�&5(r�J���)�ɺr��/n<<�Z�h�A�ܣ�:���V���k)W;�FU��R��2�����x�j�q�homn��/�ҁ.W|1�B���1}��b�vd�����*��][g������].γ{u��_KB����������?A�^���k+�^��9f��}����m3�m�fj�v��nn��C����O��B�Iݴ�]�KX����BڋU=Lʠx���fctU�Me-�q'h���;ӛ���RI]����4�<��+8S��Dq�B+\v��VE�<�T��31��7J�L�ԓ��-l���
� J�4*�?0�ݾyŒ���a[g6�r��aGi�K)|���v8���B%:�X����֗��VSi�ָ��u���#-O�;�����Z�U�[:wI���[u�6ލ�����*��UynF�m����G�3(n���t���y�N�kF�q6��ɻ��VŐy(��:�Rj� ���@���Z8�c��]�_�o�MY����Gi������U2�n�GvwtƧ�H)nԶ%�Դ�$�C��=��R�lp�f�r�V�]�[w���nK���f	��!�V�r��u��Ɩ��W�S�j��~���|��1�����
V�wmn��ݥEfېԛaFvHq�����`��8Q -�$l�e��;4��\Y�%5%���q%�����P;6؎����!G-�fI6�m���g[n��Z;l��͚[Y�ZE�k��nlf�u����nsa�;;�)9M�nd���!qdr��Ս�lq��vl���n�.92��f����N�hݗh3N�kv�lq65�np�\��f啘B�[\�ȵ���;(�$���ͭf�%�GYg��l��\eŜ�F�gE�m6i�e��F6�&�EZYiݣnj����P�K_BH~�<���}9��Ũ
�}@��Nl	%?RR$�������R^.���A|~�A}$B�)�����0�ᩇm��ؐB�|���ы����h2P@�%}$O�J��7�r	�l��{m�$��3��@��V}A���X�B�ey�u������}i�Z�����ƥL�֕F��C--�X�sXflm��*�U�S�V�w�7j�$%/)ݽʝ��Ũ
ފ$�.ɩO�c���@A7�<�X �G��H��4�C�L��1�|y���5�{;:�O��0��A{bH>rř(p��m�C�:� ��D{"_PD%d��"JW9�*��J���緯���L�u�_[�?H�_%�JDXKs�rg(.�����_R �BQ?^S��ʍ����oho /�����$���z�*A�T�t�}!���Wr�)�[�u�}�f���ٸ�o[�asUY��A,�G��{]�r=�^�*j�S��ȁ�}���ǐ8�j��܂?I_I�A�~�L�+m\�7&׽,�P���X�l�'�m��@�W�s�,�HH��[�uq�x�����ة������%��/'\�G3un��}�،k-��2f~+��|�����n��#$A�t��{z��l��oӼ���U��b5�|���wW�$������R �r���=j� ��K�	Ե߷}�Q{�-2�ڀ�误 I�6����"F���W�E�IA�A|D��G��ڟB�����&�Iw�K���{bA⯒���J>I]�[NJ��;�S� ������d���o����ٳ	�N��[��cj�?>��x����u��zX����R �,Y���컐d�~�v43"W�n�ʍ��.ͨ
��?t�W�E�ICh��V�h�yjⲷޙ�9�Ӂ�^v0Z�*�v����=zp��#ۑԺ#N�K�� ���"�{וf[�*���<�5���}�n�D+Y���б��[�+p��=�d2�E��z�Ÿ.��]n�[�w�u/^�6A�Rz.��%��}n1��G;�]�c�ɦ�3�F� �x�׷nAx���n�]��Ұ�����=-!-�\Þ�%���U� �j�1[�Ԗ�0ݤp��j� b+p��r�wX�b�gێ�j�Ƥ�*q��E�ֶ�SU��Ͽ���'"��ضVi��P�];��x�6v<<���Y�f�6��k�c�}����K?}#���3�IP���Mi��
K�r]�G�	[�z�^��ձ����V���i��0C%A�F�ݷ] ��Cy���rw�>~�w��f>~��%�����?IY�[�7���W�=�`�@}H�$�`�H���5)z�z,Z�n���.wV��{��]A��P@"�� �?H��/°g����yX ����g��IP��)�kLn�B]���h �{��=���l���ro�؈�ڸ���d��J�o�e���� �?o>���l�o�ߧ{��qX ��|$��X�݅7cy�������ٻD�V��⒐��1nYqi�1ڗlCV�.l#a� f��β�"�!�!`)	R�}s|���=;���&���c"��7���� Ȃ?H��E`�Y����x=}������/g.�/wTGuf�dH�U��5�=�[��5�ݳ�q�9ݩ�m�
��uW<��]Ŀ��������'��FO*y�5�R]��߈$^Đ~�/�+�Z�������pgR �6ł}@#%�YH��7�u��NS�g��g�'s�ߧP�-�d�#�}$_I[� �K��,��6�@��7Y�y����$���s�?�-��s\)��ڠ�9謃�� ��M A	H�~KdFҋ������Zcu��mƂ"�$~x�QJ$�P��;ݜ~�b��S�lU#tPUd�Q�Ż[<�Iw�la�XΔ@�iG��W@�4�,�|t �:��-�Az������nJw��8�m���%��/&�#�D����BJ����	W����y��.�B���� �-ҽ۔�4�N\���� #���)��<�ۿ1p:����ӕ�$�����H�����t�WY���hw�r�عJ�)h7(�;\�h���13���5�yptv�0s)z��'tx��˝Ѯm\�UC�����7�za�%�1.ێ��� ��P�%/� �+�&�a<�L����(4v�'�~_ICGT~nz����{����A�S��(ޭR�����b�
T� IH�����d���׵�g���3)7y��[�=;S���	n� ��_I�A!f�&
�ӂ�S�U��ś6��ie2�%�Vf�ȅ3�ا�ؑL��0���&~�],G;���e�7n\M�¶�����y�K���E�p�h���n�Fs��c�j��pM�ɂ��dOg�u�*����?k���y*^pw�p4�4A���%[�f*p8��Ǥ3�HAԁI,XJD	(ԙ���B�yϱVh-���d+z+�� ���dA�Hv�"���j�!�	 ���?$�P�MSZcu�A�F^' �؟�Uk�4f�ի�㖁�W��]��&�ٔ^��ˡ�U�f�xd�7�f�K.ˏ��=8�t]΄�x*fb7��q��f�?������w��D��I���%d����q�+2�>wA�=����y*^p{�w�%������J�}$�^���/��l���e��|����E)5�$�m%yu�����0ͬ9U���31(���4]�`���DM�\G��0�H?�<�׳핚o�W,�ohQz��kW� A\}�͐~JD�~Q L�}�Y
�3�8�����9��b���X�fwYrm�a�q�H�� ��P��F�6�lZ!LI�@�V��A2P_"�A�D<&����O[���@�w�J����C���A�/��%�	*R�"�wp�hlD�B�@�� ���r���O4�yz�
ފ�	29M㕬z���_<��r���"��X Ȃ?I똰��ٹ���,Z�g?oL���h�IƐH����T(�@R��^;����M�o++�Vp��1�x�Bf'"��C��-Y��m���`�]<wyJ�,�Hs�woa�{F�Պ��s����w�e~��Í��C�ϱp��b/CƼL�:�m����"ngdm�5u֮�q:���Evx�W�Ѵ�\u#�Z4ƃ���C��6�鶜���ٞQ+qv��Y�1&ݫ��.Ic�N:�=���C�]�r)�{���d�f/���m.炞ƽr���3��/��f��ْz[D��&���j���Ď���wP8�F��\��AfC<�e��RSf�u�<���K���N�]��U;���k�����ٸ�5.���U &����/4�߉���я6�wv��.tW�s�c�<�/:���vn7~ͬ�m���E��/��Y�� �%}m+�������Ȓ	�CU��=��An�;/���`�� ��}$Z=1>����пl�gl����!�e�v�3wrmz�g��9�����ٝa�4�0�q�A<ڸ��f;�h�ݫM�Ɇ�^{�ˡ�
�5B��}=���^���xe��RS^h���54G���ۦ��-�<�\y��ڱ7j�3wrnяk���1Bq#+Ӿ:�An���dN~.W���"�A���󱎧�����٪��o����Sm-�M�$�fmJ�;&��Τ�5fj��2�77M��1���e�~���y��%�����.�n�ei��&�5�7�F��y�8B�����fJD	)$�(f�ٿP����O�T0��V9��C���h�z��}��cG:�U� Ҭ+�;r}gY�3��{�]��㦻��Yk��SUt;n�����}�P�Ƭ�?r�՗���^�%���1�@NB�ڱ��O�y�`:�ޤAK��$IM��"���9���O_^vg�޿��� �W�E���/��$<�z��UFqo������<��$�ac��{2���h�ƣA��T85��5�O���C�@�"�FJ"]�-�J����C�����{ŧ�NJ�|7��/��`D�?H���%�3��{���ў�&x]-�qr��+�.r�v`䕃������@��'I�6l�o��N��/ޱ`�H�R��k>;�W]??y���6v��iD��P,�R�?��$���D�2E���뙴=�?\�?������f^�Kc�x�o�G� A��J���i��b�!���Ozł����d���+ Ⱦ�Xw�&
���d�ʍS{�{H�Qյ�.�Xiԕ�b�L_V	C�冈�ﱚ�D�������#�d�yN���� mbZ�N��Mc�} �x�9~�/�K���^���EL+E�a��C�>�BQ?��ê�ޗ6S�{���x�� �U)"��)�`35Y��IC�}%?Hu����w�mJ�C)m��̽�-�4m�Q����2W�%$��Q��v
�U[W�U��8�Iuчd�X�vh�m������-;ڮ]�]U�R�� �P_"�$��s1�xd��ID�17�+�ǓQ�eθ��sx�o,�����`�Ա7j�w�q2}�2 ����Ti��sk�oY�����8�~�Kp'�9�$���^l���۹�����?<K��_\�/��W�%CU-9b�6ۙ��Rئ��j4�FJDG�d�@���I,X{�˶�Yb��`���_I�dA�3��A�$�+��� ��4��k�;��J�e��d��;㷮]�q��"�ᵒ����%:�ð�(��k��93�F�m��y���Tĺ�xzk���c�ݲ'㯫����!b����1���������t�I�w�;ь�Ρݾ��u ��d��DV�n�������:i�D��*h!n�3�+u�%X�5�P�Lm��3^5�y��=�~{|����Q�$�-��}�_��/��}+�(:��w9�s�r����v��ݫ�n�`��D�Cբ���TV���Yb�U^�Q#��%R��<��_��#����ȏ^��y�<�\Mڸ��f;�`���<�+t���N���k�=�ޏ�r���h��y�������۳=���:c�t���u���r�$�;~��Iu�����Ҽ@�K�E^�cT�B�+��si!�@�%��W�Jd�����U��?�Z���w�,/�J�8O�yw��"r�I���Ə���g/�/�L����2����'�2'ݹW�.Aw�i�ͺ�U�TT�[U��v:��Zۣ[�q���&�z��ɤZ5]��YY�ףM�١���fk=2L<�	���v�XW�W�ǝ�8�V�ܦ�y�I�(��_VX����|��AT�e��r�RC��髮CFv�[K�q�.����}��i<��6]��:����2�����r��U�T-��yuF�g8�9ds��o�]O�|4Ӓm�i�,Ř����ld0�c/2��^nI�誶���$�+�o^:�A${��4sV�G�Q68�8�ۻ�+�UTNݕ��9WcU�%�V�'G��}+��[t��S6��h8�ME7EZ�2f�/�U��C5��xQXH�dK-`��U_��4J
�q�cI���*m�LB�fd����Х^Y�*�I�+���7�8z�;����47D+�i�d����I�}WJ��{�g^5�ޛ���}��J�I��v���Vw+:��-�RS3]�+�����W*D�x�K�Ŝ9�T	gn�}he�\�c��>�[���nڸ��*<
7f�fiLdγ�\҂�w֭S�!dl��ޝlvvʕԶ�MR�����!w� w���FX�5.������n�vPD�6ܼwM�{ ���výY�WٗT��W{+�>�}���uR����w*���2�ۛ!��l�u�-�^���ޮ��x���~���u^�9�h������;�sM�Ʒ"Ō��Ȅ�F|]�ڧ��	�/m�ʣYe�b��%V]V�
F��7�5=�5����_@EA~EQ��(�'-��[6γ���vQ0յ�Β��[Y-c0��6ݜ5�:�q͎JӬ��r��Z�a�GZ��ٕ�XY�XV�vfRE�nI�gٙ��R�:�&Yȵ�eő��l�K+;[i��f୵df]��dq��B��;��I�\ZvvF���+"̷.��vBv�6�Z��ٜ���,�M+	��bw6�[`VKj4���B��I��:�����gu�p�U��V��Z-��lwXee�)(L6���ڶ�nZvQg-e�if3e���:��gw-nl�-i�qg�6�;:136�`�"6�'e���4l��-��lз!��j�K�m��(�,ٸ�kK��)!w���i��A���`�t흒���nՌ^ĵ�2�Jd6�X�ĮYq�ۗ�Suq���8~����Q`(>�\�f�v��:�K�"�]]�����]�tv{cc��N�q�Ey��q��_;��|6�=rs�t��Y�h��J�Z,��l[[�.�ȍ����v1;���3N�F�[k��]favS��58�k<rV:��3p8WI�4���Or�)]:#��K.mV�*A��[(�VZ!������1H���|��)m��K�tu�pg@�����s���$�@�q�+���ڵ���U��,&Z�j��i��^��UIj���pfM/�\X�m�Pu�_dW�Ǘ�6
�����.��ٶ�H����Q����\�mt.u�%�b۔x0�X�S���ex�̚×k����=��\niz�s'j ����T�%q�vݶ�wc�1jp�[>R�{	t�qz�^4t&%�^+��`,A�����%4��x6f0�����W�ݒ�a�:Ma�6�7�\zF�{(F<;����S۴�'^Gρ�U�nV��4�q-���5 �pu\>cg[��2=n���G����K�1�i����뷝���ܝ���QI�m�me��enxR[+���\7�q�urz.z`5�n���|�l��G&�4���i����(]�&�屲��a��c ����t\���u�rQKn�T箎:7kee�V.�3C6�ii�:��ZV+��͸� �[ ��6n�\<�<'v8�!�j3�Ľ�tX;�|b3����	2k���7e��$)3X�ˆ���K�.�QAe�F;����f��K2�,���� �槎+uk�@��9s���v���0Zc����l���5�ǣ�G݄��P����]��4g�Dm�eyCs��������i����Kh���U�T-��n���5�f��r��`<���ӗ���\�˳(�9fxkEې��sG&i�p˘��O�fp}��I�a.mԔ����W�.`�h�z�<�ywb���pm�۝X�=x�x���'�]�˪�bEL�+�u�lc��;�L-r0��b�3�m&��6aq�	��+E�	I�v�!6���!�c�u��y�M���f�qی�����cE- ��G�_l� ��CBqٸܵu��Y�82�cd�3)aV��шk3i�f6�l��������\����/U�Zk.l�k�xdq�Z�m]���`���yU�F&�X"{�჻V���!���h�ӍR�t��P(�(1���@�������堉+�& A�+#�����@�K� ��/��Ŋ����.���]��_x���X�%]\�7� �t�#sn�/�d��2EdIC�c{2^�1c���,?H��>����V�9�D� I/�+H�[^��؆z��v�z��$��{5���]�_�;{@�p'�<l���+�^��4�Ƭ�������?I�F�N��z*E�oo5�ïFj�h��Q�~d�AI,Yr�$�������o�ꀾL��4#c��h�ѕ�q��q�IA;I4k��쭮�L�¥_���#�(�y�X���!(�5�^���\D�W�h��-�(��2����Kd��R���f4���m[I=[�Œ�u���c
�.���s;M�R���y�
��X^ʣ�TX׆��%����{8�7ơ�]Y�2-�3eX�� ^`���R����=�Ųk5M˦٪�� ����*E��͗��h�z�� N�V2 ��D�I,u��d��#6y��W�פ��s�J�:�D,+�D��"Iv<�����X�A謃"����?P�J�%��kD�mM��]�fzp��u��!�J_��K񒳪�vx���^�5x����������񞯤�H"D*�/h�x{�����f���,���J])�]�bޫ4���H74W50�S���t�veM�lG�������n����%��~s_��u��r�ϝ|�a�~G�&�@����uh �%"$�X2P@�l��'��n�|���y�37ۆ�ԽQM��[ �mMBr$�4,�҅�K����gΐ �'W�D4)H��=�EV׳ڐ/��>�ʊ�PZ����_�cskq���Q#�\Gm�,`��w�Z�^�5�Dp+=VH�{��Y��Bg[�M�g���N���c|����Hs�X?��g� d��+�$B��~��MPgmp �' ����I,_'5��R��B�yׁ���]�[r�z�;����R �R"IX&JA��H�ܿ�l�j�����ܨt/R�E6_�@�x��r$���$�=�8!cb���ؑ>ژ��R	�]���QLp�܎��g!���p���#�ǖ�����E��?z��d��"J󮼞�ߑ�}�T�>�0>�sxTv���( A ����D� ~�H�\TK�v0g��~?n�^�ݙ��.���y$yĂX�QJ1�F����W�y�ٓl��@#%d��"J����Y�-��������7�˵���<�o��D��E���,_��H�ǹ�[WJ���,��I^u�7݋�Z�U!Ӑ�9����d�Kyx=�_xDղغ>�׆.�[��f�۫_zt�ZZ�v���&�>T�OW�'�,��	���ϝa�s��g�㷓W�(xz���#��H��"�%m���{'��ʡ_j^�{3�[�-~YA#�$c�/�% A"Jnn����7xx�h�����\�i�zuن��q�V�L���+�U��=\J���eVU��Qq�����v�?g���f�u̾R������\�&�n��X ��_{�Ib�2R	+���~���9b���A#җ5��7��>��N_\��A3��H���6�k�.r��h��6�v�����^=}Zά����/��˙]�׾ gRG����)|D��N�ω��ې$�)1��[y�5��9P�kd�c�#Ce4�0�m����m��Z17j�;���~��m�<�<�ى�u�Ƿ^�Fo*�&COh�H%l�YD �%^��Kz���o���e_pŦ[r)k�[����[�ww�T�b���}���U�y����3��x:�֍��j��t����;��WS_Vc�B���bUE*�5e�٪+MP:����iM!�ٳKU�Y��Y5��"u�l�c&���Հk�8�[�k�-�Hy���g�����u�����D��%ay�f
�����M��'�2�,bZ��K��5��,�-Y4��c���Su��S����I��]�鸸C{
�@�L��J	u&B��mfD�c�#�	[��� �l�E���6�z�\�u�������ֱ���l8A��>vR�u�i�B[�uq�V�^.��9	�����#	?%3�JE4�o\�ɭn!�0���&�^�kuLoW��lY�� �$��K	����S��ܠ�1�|�V��>8�h^Ș��j�ȧq���ʇ�Z'�|��&��j^*M���Gb�ί�!��A%_%@J }(͈�<«۵�o.7K6�&�s�f�Dx���n��~dmw���9޾��k��5|���JE-^y�#D֧��?^F�A��E�m{��w��Y�� {Ԉ�X�A���2D%���	��e�u:�W�j�5��:P�kD�c�!�~Q/��X���T(eg��Ț�+�EX?�#�O;���ɂ-j�(-.s���R��J�]iv��� #ӯ�+H$IK�^k���նL���հE�O�әp(��ہ'}��ȾPό�_�ag����M��Ԣ��yj�:���x>�׻�Э��yj�z������8�;˙S�J����[�j��ؐv��|�(�i*Wׇn<j��<��*��ުN�\F����»5׈��X������-���[��=t����� �2P_"��
�7#D;:�⭺Wv���kU�t����َh�܂��%|��X�% E����.�c�^ ��b�� A!�^}{�{s<�[ǭ��#@.�c�FsLJC�Y,s���&2EdA�#c�U@̓�y"��y�#D�����~���ұX�%|$��\��8����J�H��b�������x.���8C��wf�c۷n �P��V��|� A �_I�$AJ{�w�Ƶ^�J��Fea���1�}�N�n��o�X�۸���Ո�n�J�R����>�D�ϯu�nf�����;��3h�A$P�`����v{�`�@�� L|���L|@�X�"��o��Gۣ)�i�b�8K���n�u����Kj����G��uj�-�^1k4�{q)��1Lz�0�ګ�3]W�ܭN'����H��fJ�I_I%�z�R��0�P`��{A|_r��iwzo�k�ݓ/�����V"V=�t�����{����p�ݫݤD�2R��e�0AԾ������7��e�d�i�J�'v���IH͖f��7�����$�YTj�V*��ы�vP��8&�N1aW�J���G,�����Y{��'��)�JE|���"�U Û�߈�c��wv�j� ��αfu|�R"Ib�2P��QGD�������6��ܶ��?*p���d������K�x�Ŵ6�����rŃ�K��D$�����+�޾�~}1fWe7�7^Z�^��j��`�i�U�^������(#��w-Y��S�޵��?s��$�P��f��1���0��4A�@����|��N�ń�樾ʙ�[���7/����ܻ�S��Ϋc�6]UN���=N���7�MIV��Ղ"��m�tv���s5�i�/�$t�D�ł� �+�"W���ڭ�����П�M;�v�Q�j�ʇ��s�@7"@?H��I,Y��9��>���\D�ԏ�!!:�ݐ���M��(��0z�ٙnh(L�̔�R�B�U@�C�fE�R <��d-��B�Wx�m��"uǘ���v>���)$��CYaoV�\C�>�r��'�v�x�P��~��)M��F�tr�\��}:��I7�.��񔫽W&���Mrϭ�_\���n!�$�$�߳s������y����_asۛ���`��R�c���8u�"�~��N�����������wU�R����۽S�׵˖{O7��q	+�#�j�?@sw����,�E;���b��Ip����36vd���z�Ae��`��WR�D]��V�s�7��)�;0��̖w����ߺ��|CU;��]��*mH�U�� F��
��e�D�)�֫[�K��6h��%ٗu=wn��"Ntz��Mtͳ�]-�cf�h���^��n�H킝\7��n]p=��Ӯ`;lt[�]t���t�n��ήF1�q���]pb��m�mk��Rf2�+��nC!���7i��u\�eӃ�c݋������t�f�v���߁���~E�M�1�������ծK[n��%]gPQ�ڭ�55sa����O��y��J>n�j���Fw-˥����]������:r�IP�.9Z}t%�{��W�?nO��[7zV]����ݑ$9�Y�Ts�q�R��t@IBH��vB��:�a�޽�܏�������fr�s�JD$�޴������y�O�}%l�Z�]�S;��҆�@�S����
�E�<Q򒀒 $�Ar��R��rp�{>�
�.��߅(7RW�S"2�a>�ϗ߹�}���vٹu���-f*�wl�7L��d�.S8-t�U�J�&�
6*��@/܀~�"E�v�r>[$����s���їk��wI0I�J��ayi]���CHO�1&��C��.��g�G��V�:_�TY]��Y��{�}z7f�0���\��z��Ċ��\����o�z@��r�R�Jfw-˥����-��^@QwP��wf�]�^=��R�|Bǐ�,o�d�{ꔞ��y��P~��~�J�#T����FVnc�7k���2Of�N��K�Gy�q:ܽ���盧܄�}%|$��$d&�������oz_l�����+��Ⱦ��"I$�^�Wv<��8��e
E#b��6hQ$�Tf���*쐣E%0k����6[���/��M�ǧ�Y%}$]r�k�w��I�����Ԟ|��ݾ���JD$�=Ʊ�/y���ix^�}��!�{4�u-�]�;���_t���{���Uz3�f�Π$�H���d^��3sޖ���{,V:<giٹ�d��Heu]�,����ڏ�OvUڵ�N��U��~�u��V&��N�͙��/g*Uy�ƹu�W����n]�Z�d�n�s]��i�"�b��
w�]��QDq�V$�\C��^�q���e2���b��h�\���JB���l�fQ�m��)��*j��ۻ޹]�]\�ە����@�U7�5�|z�]1�r�lU�2���lh�B�f���B��X��H����UZ��E��{.�B&빝sz����+{�}�l�1�*@��;�܉8��{Β	&n�3�X����iXٹ��Ue�������Tk�,�z��6avs(,���^�5+3D8á�!�Q_C\��r�#�痢�uT��}o�L�ٕ�M�\4���C��ғ���Y�F�p�]�g��7%�Y���Žڐ�޾����ٙ(<ު�:�ݳ"�R���e#��V�z(S���a�"����t�b�_{���Z!;=�Q
켅�9�H�Э��ʆ]�[��2gKZ�o_e-���喆l���#�3G]�0�6Z	S�M�"�3hE�b;��7�w�o�շ�u�iGpM.�V/����:㾥].7�\}��H=��}���隗�G�
Vaf���=��߫��f�9z�.o��Љk��r�]z*��kRVf�5���h*�}h�ʝx�mL�Q�ε��'�v�z�K~x��El�A��}�Ʒ}a���j�4Vs\��q:��d�w���>��&����©f����Y+&m2�d�_��c����1��0���]�ې6��]���؝��Ι�!�*ٶ�u�vڴ�9L�!�ekv���q�av`�v]�sc��G�mGgVi� �,�Y6��m�DYӗ-�3"D�ݻdf�H�X��6�Z�[,�gY6ә��n9m�d��vaY�Ga�M��a#2��ل���D�ZhB�I��g%����[[km۳p��a�C;kvgi�d����p���4%��e�sd
R�  KkI�G(fe�ۜ3;k"q� :��H��9ʹ�5��$qHe���gm�l��ve�m�0�v[��G!��K56Ԛ٘[��m�i��jt�ֳkhq9ft���ݱ�rb��@vi8�mfZpV����0�f��i���8��6��s�u�G(�,��mY`	ɷh8奺�IH��6�	UsJ=�ޑ%����w_��}$_	"�JCʺ��s�;w=x �N�$����r��3��x�}K0=�tuĿ5J�T���I$�12ݝُ[�g���.����!�/��$UY}B��*\�v�hһ8��]0�F�&C��ϕ�]� ݹ��/�Jү���u�I7�+�R��/u)�Վ](j�RY��ꤦ����))JI�wi
��8;����D:���<�O�Ym(��@�7d$�hPۏR'I�>ae�_k��JE��d�{2V�&�v��|+�I���o�^r����	"���$Ҋh}u����P6%��W�Lμs.���q{;{W��[�$њ���wG�S�v"���N����VW^*�a�5�vtO��M�r�����'�~�]a��u���0+��ض*�@iO�G�)(�����/mU�w����O�OzJ�s�\���$��&�<�^��u�'��������4��c4,0k�X9Z��A�wZ�`DХP�Ub���Q���j@�%!% u���Dn4��ż̓E�Ks��r,q�>h{��$�~�qM�kmn{��f
n~n�V�z�)�[��	�1H��g��ò�Ky���}@I_	%WZ��'΅�1V
�z���#-���߅*}�$_I_I���9~A�L�L�z ��%!�wc4�7�,u1癢��&MR��d���l�8����HJr��ql���w��S���s�|�_?P�/��;}�-�=�Yܣ���M:�g�y{�4�
v�,�[s�W4Dq*�u�6����>}Cp�ٗ���^u�p[�Ξ��\�|���y���Y�-o�����=y�.-t���6�h��������P7�묭�]�y����j�P�/�����۳�#��f��HNn�}���$��r�И 4���u[����,t�P���{E�J��]Bm),�/&� d�y'�N�qg˷f7<�݃fuMg��g�v��ތI��wgi[ �ˈ�z8�;�;��`��K>��SŽM��>-ڲA��60�����e�~�Z��R6d�XCT��l�&N����Gu8ۧ���d��a&խrM|�'����L^w�\~���O:]�K�1*��^��_9�I_I�.y����K�y�cϗ��5�Q��Z���>��9�$��g^�/N(!���?[��$RE𒜠�b;�zn�y��)Jy��;�q �RD �I�{UPwy�w���_I�}���~�Y����a.ݾ�t�G}�ې���R��4k6)�۩�ܘ�y���O�N��t~���C�RPA����x5R{�(��A^��l�]UGm�����)W]Y�r��6#h��vt�p�z1k�yg�~�ۏ�\����n'q�^�Q9�a1�+E;޼���7��@7(l�D$����㴅)g�w���H�Y�;.��z�<�v��/�NL=�q%q�s)ٮ�6�Pجu�Γ��hU�C5b�u��A�X��+�k����K�����5��g+�P��Hj�Qsm��bq8�+JJ~I:ي0�"��H�i��_�����5�^r>iJPI%Myj"���jɽ�$��~ޙ��%��N���#�e���"\� � $�J5�O]��I|']m����9cj�y@��IO�)��%��<���3龻7wwb���]�6��-f��K��396�C�qRd���1Č����_���6>IJJ]�y�a�cq��g���	��˩����_t�$BH����J(�\�wu/oLo�Z�f�s�Ⱦ~�;�ޕ�~�_vP~��H��$�%���`�����{�)���R�U�%R�ÉS���Z`�OVdr꺃�s	̒�v�U�-�S�ҥ�)Hu]�������TC�X��-w�sd������+}�$�	*9MPu=��(^�ݵ'/����w�v]o�tI_s��V/R����+/q	"W�I$���+՘��wy���n�#+�>��6D�BH��e�
~���u����	R�ZP�a(L�2L�4fؚ$v�RҲ��.�vl�CE_w��~}�����M1�[c5�1�5z���wT�́���/��$_}$�{�֏x��h_�oe���isuu��L�6���ͩ	b�Y���}:f{�wW�E$C���2�*���6����[�dep�����\A���	"W5%^�{�jN��w��*H���[c5�g~[��w����w��7ê�o�V�����+���3:\������T��yj^�ݵ�2�G��R;Y��Pu{�x6˳6K�R^�}{��~��3R^	)�$��O�i띙>N�=��b4��7��MSO~�㔡%qEv��v�2x�T��節]�*�Wi��P��4f��v/O-ے喐�%�8ݺ�S����z��x�<��+�w��?K~̌�}Oò��l�W�^W�g�+��$�$���Jb�,Ol�u���ٗ)��k����������[�p��+8��}O|��@I$�$�ǣ�9w��Lԭ�f^z-�7UM=�i�	P�)"�N��u�n�����߄��]�z(�y�<�?�!�H�:���/�{�BJH��I·�&t/j��/�g�����ݦ'L�(oy}$@Hr��:�jy���v�=����k2ݵVn��%H����M=޻̳}^՝��v���W��8���Vj����v�5�t;|��=W�6����V�))V����Q؛ٝP��ee&��1��G5�옧�i��s�tƝ�m�6n�<g�~��*���L��1^��o=#�t�Z���T�kF�-�Ɨ��R[��<�/:(���ײ��ng\�6�r��n�L�Vc���0ލ�m�]��6L�H'��٧Z��ZYs)�ie�jH9n�Wlm��́\K&&�)`��������G����z����듙\�N�%QE�Y������Ÿ���
�y���~�^�%#��O6a�d޷>����)gM5�R|39|���$RV��::��ӷl^���^�תuE��Zy�� �RBv�C��C�W6U���N�$�`CՍ��mX�׻�i�:	�v�LN��P��/��"Yyu�u��9�g���H��̜��u���X���|7��{���������)"�IRE$P�e/}�U���E���-�|����ɘs����Θ?mmKM��}fȿ�T�q&�3̆���ukT�mJ�m���C����k���������`� �}�sӠ����bu�f�W��N^����)*H��/����D&gx��˚b���om��Y����*���δumfʼ��i�'��g]Q��e�1�}�pҐ�=G����A��\s�6��7�ϗ^\��]vֿr˻��s_�}$C��ݜ�{�wT�|$��.���q]����;ݙ�pޒ���_�)"����;�˙��FkNP�/�[����ى��=�J���ڿ������yn쁎>	)	)JOh�Q7S{`�6�}뗱�R��_��]�� gr>@I_	%�y�V���<r��r�+l�B�y��f�c�[k��W��`�i��4�]
ifJ@����p>�RRQ�{��(����b��[�,8�J�K��mJJBPR>�N��^�\Dכ��"��cɡ�oӁ;�%����O/=s��b�h����? $�$BID�7�zR8��{*�ܭr�^�R�2�{���F,a�n��/���X�epַ����-�f��ֶ��fF��C�[;
�־�K.N�=����>�)"�/o{�5��l���BQ�{Y{�Q����ŵ��{�}��U��������/��x��g��^�>�ɪ����v�p'K~W[�I/����̗�/��vj��F��ݓC�!��`���q�ض-Qn��;��	[�rt����� =(I�r��w˒k_���}���{O��[���	"� $���n����w��H�l�={�Q�����p��q�Q��5r"�>�=̙��D$��J�ٻ�wz
ˇ��T�qX֖��r���M�����}%}$BЙN]h,A�nd��$����/˒վ�R�}���9e1���̪�D�H��r�{�^Kj���Sf5b��w{[����$��8ph%���5�2�_���f�~�J��!��k+���e��|�I4}%	"�g��s�0j�_y�{��WJ�gf��z:�l��JE$���p��'ϻ���ȓ������K��-&i����f[�WU�(]J�_XDت�E]���!��%It��Sk\ ���M�K��!��4�߇ۙ��Ix$��X�m�;�����<�}�0�a��ަf}X��m��4��يۍ.�������G��##Юn���z���v����߅�5$��JBQ�B���fos�K7�$��k��Mn9��yG���}7��R�e��J��4�/��%	%� }��Eڳ���I���+Ե^��}6ދn~X���v��w�~î��u�v�z�..��=�!�EWp;%۬)}��>��22F�������l7G�ܗ�A]jK�n��%Y;������pc0�(#��^�S�U�����0g�i�,��gTcLo}�r�JXy���v~��U�vJ��I��KH���؍୲�r�w����͛�0$_cM۱/7��ݮu�L�����]�:9����!Ջm�\���2�a8�k�p�Ү`Z��m�[�*����f��t�67�<�����Ņ����ޙ�*�H��:��[�`�����f�ɇ[��F�Yg����wt�"�ͩY�f�S��U5ds�VD�*p�A���ǜָ�δ�7^�mM9;;:�J�;r���s�Pc"����A�f�iک����x��R�ʆ�w��k��l#U��w��:�lm��t�		��Ve��Y]��kl�W�,��8�l�{hv�6�XH�pA�Q�ҧv�a۸yA}�YIDEi���ܩy�#�p^�H�܊[���R�5u�<���R<k,�{�g˦�8�R�pm��{/aE�U��tU+',n���h��M�\�}�^͢��c���]Y�4Z�<\4��l�e�����t)FK֒��^�*�6������u�t�#{;���|E�T}S^r�n�}ٕ��uUF�-�'�6�[t�0ovQY�e��ݓE��&7�g-4-|�h�U6��fJ�]6�˪��,S��^�����a7�Z�&j*��]�Cڮ2�a��6�~�pi���X�����}�z���s7P�0��+b�+�z�|^��$˶5�tַ���L��Lk* �(��δ٭����q���h�r\��A������(ᶂRq�[���.&�6v�N9��)���;+$-kNe�۴�GQgZ�	N�98GNٛNT�Ht�B\
�')܃���pqD��
�;l@�$C59�ts�"Ve�֬�nY�`��s�:3s���v[d㣧N�%)N��S[��s���!�2�v��N8�'
+-.#���M��֋0rvk��9�qw%�8q-S�ҳ6��$�G Nr��\���!��f ���Β;���G!�m�G,�ȡ96ܤS-(��9�9��6�\6ܹ܃���At�e�E��jED\E)�8��$M�kQ�%����K,�^���i�a�DŃq�C\�j��R�����	c��Қ��ɣ���u���29�Zl=d���Kz�B#v��"�l����7O,u�+6S\X$�s.V�^���g{l�	`�fDs�u�s�+왐�m�ׁ
cn,��E76G���^�L�/v��ǉ��h��	SUl�:�nIm����N��Ye��qږLǋ%h5e�8*�����*��.)�i7���Sw�cA�Yb�*\�4ݵ�]��������)�Vn=�:0�<�n����R�J�V��x��iaq�F�g��vٌWkN�x����-�&,�����ʃ�Nm�� �GJ9�6�Vm/^��Nx.��&��!��c���К0�YL�\��Zz4(��sY���K�K��tz�����ՃΚ���Zc�����h:���\��y�]e@��:&R�6�ض��ic��y��:5�tn�C	
��%&��`@ �┝<�z-�%�T4��Alc����Z��V	J:ת6�<�ո�v������r�g�ͺ�a�j;<'\@q��� y����\��y퐺6�6ꡫ�/F�Z:��+sd*hæ��vTĽ���Ql��bl󳛃 ���� ����u�2���I�C�-�c:��ݠ��ت���N�<��u�B�f�Vӗ9���Ah��*O��`��[E�;Is�iV�Y�u��n�ZK�H�1H�:LjXL�,{K��6P�҂Mpg(�
�>ŭkuh��û�lD�<�����r�Y>�}��춒]n%��ºP�`�m�ݓ��:�y�k <��h���d4m�1f+E3��Z�)��6�`Gc��	��d=�k'lh5����z0.�y��Ƿa�kT�(��6DsX8���n���f�'b��_h��r�������kif�����CkI�VB2�gy�����k=�ZM���m��0�[@���:���$nC��m��.n#<uv#��r���P�d{G�������붎<�ݚC���Mr�1%���6�W��C�[���ݰ8L���-`]�-��AX-W>���u[6�C��)���n2\]����ssòh���%��Gr�r���vհFn�`����k3jv72�z��{�ȣ��*2���num���Ԫ�jґ��ô؎��n�Eq�Mn��z��cs2c�p*��1u���%�iMa��?|����Mۿ<�z�ś�jM%u�϶׈n�:r�B��!�LMEG�&�{�Ԥ$��]�N�>�y�q��<�u��m�`y�H��I�$�5J���|�nM�w�)��0��7O~Y�z��b{��<��k�������PE�sҪ����s��pu-[��+{��� 'G0	"D]m�K�
���\���OopkS����n�[m*�^���~s�C���*H�E"�cڷ=�n�R��R�܇���׷� ��+�(j�R�j/c����3̪���|iB)D
�6�[mU��kN��J�kM:�]�ǟ߿�|����U�Lm�s7:�.}�ԟ�����y�ң�H�����m͞�+����z�ۨ[�N^
�n��I*�3�Bn��c{�Ϗ���H�a��$�x�r��$�vw^m[��*j�[z�)�P��j}��ɶ�N��s�� I:���X<�e� ���$RW�Nd�Rp�j��wJ�<�Rݡ-��E���D�>�pKA��\�~�vP���H�{/���%�g�r���sף8��q���^7�+I%�P�bܧ~��m�pOE�̛�N�ؼ1������'��~O�SOt=����A��Ǵ1T2��.��c�\�t ͘KM�ȋ���t�Ui�{�m �������{J���pݡ-�l��V��Oｭ�_I_I�KÁa���Ɲ�ϺE�ߩ��f��g�m��ӕ�~I4}�'��w�ؕv�{��%$RE"��x�u��ّbK��7I��R�̭��_.w7N���tVt�+k����ȋh�GXh2a�̻7��^^h7�Xk�2ڔ2������;2oq;�b���I�	"WOa��^�Rc��W�%�I���1�.��f���̨�^�o��+�"�H����˻���A�
�\Sf�*>�5�G��/��9	@	+�o�7�nI���#�]һ"ͥF��cv�`�5��kA���q�n�q������~�����S�O�i�֧��y6M��:�v�S?x�w������	(I5�O�����>Ʀ.���v�r\7��:�nn�KCݹ*��}�f��$�����A�?[�<Ĳ�Y=��;������I@I�Dn6P�W�;tN�'����k�<�վ��d�~S�{�t�m��t�8�z{�ާ�vh��n�*���ݐK�]�Fj�C���x���tp�J�6ɬ�/Ӄ���7���K�K�u�C`�[>^!��`E�H3��S����gҗ���s��L��h���	"taӤ�� ��Z5v�ut.�u���[�]��ևfrm1(�nˣ��Llj��Oc�Վ~j>X��9��p�3�D�5o~����[���c��@I$��t��MN/=@w.��h��~��8�ʞ�: =*Hk"��4�duQ��Ϸ+�ܾ	)	@I���HJ�m�n�޹PỜo�xm|��I�T��;b��*nL�˯�t5���E}��>����O��.�mHoJ�ۅb3��6R>JI$}�W6z�=���'4Oc�^I��>پ���I��R�Ǭ�Ō�_r����duf�я�֙���K�Gw����!�6�sY.GX��8#�5�.U��nmb���JѰ��*���72}��qI�x�X1��u���#]�Ys�:���V.�v
Dk�m�Ѹ��e�BI�1�ݲ5��F�ۻ$pi:C�n9t���j�7OB��Feݠ.�`X)���&����tYJ@�Β�� �]/WP^vNz�4�і&��I���3�p��=����=�0s��h}�vz�ܷB�k��m��沛��[gn����85�낎9��lG��>���T����	B�4˳w�'u�x�cė3p������j�v�o�����IBH����Or�-�f�{A�(U�N[�S_=��~I3�"�W�.��hr��{�C}����Eћ�N�^��}x�&�,���8�=���j�� IJJ@K|☯,�@���?x�I�;���ҩ�Gﳚ��/��J�'�^��o���� �I�Koi:֪��̼����X���W����J�/���$�%mLY��!������\j��X���>_	�&$cz���<<���?u �y��:[�u�ͦxJ�Q����n�90n8ت���)]]}H��y�E%�s��׺�EO�G�W��{G��[ƽ�IJPO6�n���[K�MT�]׃�]�ig#�I���]uo:�ڞȬ�n�a�W`k���՝��µ���9�XpH9�V��Thc�·w2��Cs=n�B��z��ze�Ns�s�{)��I5
Y@孩Cn 5����|$��׶�rV����91��u���c���I@I�w���X���{~v$��D�s�­��դ�E�b��r%���5e>���Bz!%|$��$@I�[�Ք�К��T����o�?+h����} ^�~�ɞ�VJ�0����X
'��1����[`���e0�4c�;Bhiv�	��آc��w��]	)IH�S݅���geǡ�̙�<�E,�Z��E$_I^s"-]�ӷ=�m�Z�Ct�밫k=;rs����7���Ijt՚���b�\������$�-�V���.��tў6g��88f�*�Ub>���Gn°#P�u$���8��m��l�|��;���� "q�b|�Q�m'��v)�u��v������/��$_Eh(���ѹZ��H�_���Yɑ*������x=��tM�����_I�W�D$��jmc���h�^y^�9�gc�f��Ҥ��&{5���z������W0{��vX\�h�8t�M(���3Bk�
\���z>}ר�RI����3Փ�k���ݝ���س<4>_	(ID<~:�}�9i^��7��|�ԝMK8�\.N���L�B�.���[��w��"�!%�5�<���f�]j<���]�����	)�%!)5����2��ݐ1В����������ˣ�-�Xu����kr��3���Z���n�fp��d�F��]L�����b�U�gDZL(�vy"�]��.�nw��]��~�/�����H��D$���/8ӹ"K>庼��K��ڂ_�.���NBJIM=
��}��T�]*�_U h�Z���(E��<�z��8^X�c���iw������t�d�����rמS�N���Tw:�vܩi��	���BH����1�?x��3�C�ݑKo_�ۏ*v��Yy�vP�rJxn����Ӟf��?/��g�E;�`�S�#}C7��U�q�A;&�[��M�J>IO�)�n>���Uz�_�ܥ��U[��z�1��߅�#lM��\�_�y}&}$_}$Re�f�4�TC9����w�q<�;7_�����$_I}����ތn�&�Y���}w*�Du�}��E}%
�\9�*�EBon#h�Ld��hm�����W�^���G���]K������0XJ�E!u����+�����s���1F%0ݎw���7���4��������r�wYWf�<���<�b�#n��f��V�iQV�豎B\s�v6/Tk`�=m�ZxQ���?<�m���!�Ż f�m[q��Iў�����pv�7k�����:�G�{v:���x��7ܽqh����K�`7m�Ìt'N�s��rK-���F�h��
�?g߽����c�g�w��4u:zw\��L��ݸ/3�f�����T�:����H��%}���\���>��X�:Nȇ�'D��.�~͏��IR����m�³��A�|��|��]�`�,O@��j���J�У��Ưh{�BI&}���9;e|o!�nM��6��vû�o�����)JH���5�oo�<�脑����<�=�'�b��ۼ��R6���f��}�|��}%	"�l�1n�?B�jꊯnf�Y�r�S�=��$��J�ڦ>;���,��4`Eg��ŕ�ôncF�ͥH�n���MDDE3U0/ ��[K�$�F?;��q�w�g;rx���2+v�"����$On�U���&��=�e9��α!H7��f�Y,m��x��Z���v�r�3UX��q�8��-l�?O_���_t�g���G�S�!�̾�����7)�حxr�/jҩn���"D����~����y���©���܍Q�J~I%�k;�+G�����U��R#7ί[����cv|��@ہ�ʒ=��?T�|$�}%	%�u�a&(�O޽b�2��ޔ��v�v��ȍ��o[�߽��IX�R뉍�k+��V�p���v�����xM^ Ҙ����?{:O�<|�H�)����/nd_���Ɠ���3V�*=�od �HJ>IH�-��h�U�l|/4ۧ^��4z�1�6�^���^��>X�Ȧ�k�ۈN��$BH�S�0w¤���xv��m՛�[0f�A\��ز���T��|�����p���t���Y�����7�v�u��&�ά�X7�U�
Ύ�.���f��&��ܭ��F��8Sx��a+���k{J�V����Y�ҬU�>s%nn�B1���w1Ġ���[�GRR��:�UM�2	q�k�6Q�,R�H��
�<��3K��n������"kb��+�^���xY�"(�<���oFՉ��a'��F���ۜ�^,#{�L��� �r�G�˶��g7�ecWZ�7J�q��W*��-�����`�z�a�fa�;su�{$�;%��T�Ėm��m*�Ys�gfVC)+4���$i��劣Ȗ��k��z,�YYv�;��^U�*ҵ��+��De.a�w��/7(�Z��&Q��c]�㒳 ݾ�$5a
PC{	6B�[�s���!�w���Bv1��9L"�U�2���
mط&��9�KN>�u�EG��c[�{�dV��7y��䕚/5:����Z�]�쪭PZ�a7M�Q�^�4��ތp�b��V0�λ|�K��]�u�����1�6�7=����oRUY:+wCn�q�fu��x��Y�Xoa��{�����۵לA���V��;wul-J��]��<���p1yZv�ݣE
��u6M�[;�fl�e��QBZ�pv�ea�k{�6��UYɭ�ki���ԡk�e	�<�f��뭕:�e��-6p�;U��u�5.�ѷ@�ݎ�i6�'�Z��6�˨lv3��*�?��e�#�Am����
NmiYݲ����%��r�vh�GE�ZRR%�s��t3BI�f6��NtDQr�և'$T99��'GI$�l�$�:t6�r�m�maÈH'9����	�qmn(�;�s�+;��+;9!�"∶���6��NY�Npm� ��N9�8�΂��B Dm� ]�۴�m��!BI�;qFv�NB'HI�Rp8!klmam`Q���.@s�Ds��Iܤ'���\rBJ$�G'E��8r"�m�rTEs��aDND�
tH�Gu���"I�ATmY8���p�* �8��8�(��EU
�AR����w�+�����R��� $�I ��:�/<�kc�mN�?%�S��^�ȿ-qm7� �<�;Qg�W�׵�fjӤϤ���)�!�!�±��a�o������iٷv�m��$�$2�6v5Tf_�Zl�����0X-ܖ�bܬ\��'��<Ia�Z}�f�Wf�+�>��6��BH�D�~���9�͖�L'���c3[q�� +6w`$�%?�ay\=�U�S�J_�yO۱2���^�ȿ-qm7�n~�$�NP����2�r ���^	+��b<ߞ��8��S��{����ݞ�{k�BH�T����|F��]����{>DK��Ʀ*[��[�͋�Ee1zZ�\F��ݛt�l� ��fY:bhFY;��F���ѹ�֧+���S��5PI���L��T�:���S��(7�$�I@I�H<�w��de(�����y��b-���ꏒR��Mv�}�����+}��ꥼst*��&���!fEft���K��T���Y��;��OϿ_<>H�{9o�<��әٻ<1d/�QUU�7��7�&IE�m]/Ó��Nf�|�`ı����a��H��)T��Ǿ���P����$���I�F���]K1�V�w�=�~����m7��܁��H���QܯnK2���{�}�d�`	)�oS��x�f��߶�R����ļ�=���LH��IZEx1�Uߌ�u*s�l�584ߌ7���ڑ�Q�H;.cBt�ϕ{m�g֪��6EE]k�G	ݷӠ�	�?r+j��i^�L�،�]�^��Yy���꾣k�-�՞�=`ͮ��s��-���������te�J�ʇhF��ۃ9n! \�x7ha6b-�W7]lr��ڀ��ei����kD �3z��,ѭcGlrq��j�[PW �8�ϯ�\��łݭQ��b�,!WC6]Q�1փ�İ�k����/c����V�>z$�=#Bv5�7Wm���b����Ps�iyш�)٭<��y�WT�c������X�֙�[vp�n��ET)*�(�h�]�*���t�}$_IIr�����G��sp�z��{\w���\����X�~��O͹Fl�8�1ӟwC���oP��>���EZi�k�5�
ȐF>�D6���������"M�M|A)����H-��	iϼ��#/��]}'�����;��H�A�uР[���t+�r-��/�B���Y@b��p'�}�y����|�>{A5?Tez��(����+c�Z�"D ("�Ń%[	ֿ��9B�-�׷gF�Q�6mp������	+�JG��{|陾S��{�/��������3�[Cӣ����W!��j�՞1���l�U]Y�2�\�����ˎ�X#�4"�����)LS�#�|$<�:|}+�ut#�_�ޤ2 $�,% Fu�
�b.��+��WT*ݏ/J����x���~yY�̲Fb���7#��L��80��p��g����l׽�.*Ӕ����2�F�vk�_��G�=�?U>y�λ�W�΋��AMM���@�Ϡ����@���:�	�HIH��I% ���/F�C�U>9��x�k���ǲ$�1�	)��R$�z���WxE��(_H���������3�R��#�} �^��/��Z3���}�_I@$B̔���"H:�U�z���Ȑ��Ɲw�<����c�%5?P�"JQ���ިJ��b[V}k4��=��a�,5b�-ѵ�,�Ů��3v�5�3V[I\6hↀlg��>�˿��߯y�d���w��opɧ�6�Z}CVg]C����	�:�� �H����JD�R���ԕ��y����oԇ��Eb�v���N�P�ܱ��$���P)Dz���j���(dȒ+\�9� BRE�Ȇw����h~��N���3�w�y�cN�<�����uv��זǏ:Uݷy���(����(Ѯ��^����g��w��~��|�f�w��X��Z�FVS��W:�c��S@��2R �$V��P�0�j�zPVm|�,��R$f�����c���w���P'�I�k�
�tu��}B�?{� d���H��$A%[���묳�0v��=���"w��K�8� n�J>J/z=æÎ��N�9�8�;�a���]�X���X�-���v��VԷ;�0[sj��9R�⻾�0}�X��l���ϒ� W{��S�<�xK�������߮����	�h���Ky���r���v/{����=�Vłl���w�^�<n�4Zr8Q ���"HIV�ջ��A|wi	���Ĉ d�~�%���|�WX��yd����MC�o	��$͡@�%���B+�r������F�C�B{B�?%"~�{^��<��K�c��?z�9Ȩ�O4��T�=3�4����n���e���G���c����]t��2�~W���m��Ux�U�7n�D``�5�"��n䘯�%��8��^��X���$$�P)GL�?���!���8^�<n�4Z�<�A��E���~&���rݸ���b����R���eT����^&.k����F�t�u؅��,�2�����}��ˎ�Z#��_
�����1;��MC�o	}WϸwM6*���P4Em�ܢ�J I_��(�7Q\���c��|�	�k���g�_	a��q�?V��(��S��^��y�	-��#�"~�$�T+�|���RUn�N���z}���\-oWܩ�"Iw�����Z�}���֓ ��$���������	�bx-��� ���x!�'�Ǿ+"H?nȐBJ�R� ��R$Z�/&������������h^]9������SD� d��?I~~�_o��)p����U�d�E�`�+K��YP�;#c'����םWw6���e��"4�Y���®�
X�]]��.}��}�P,����-*�߿�����ݛ�������� ��������s�X�w4��[s�Vl�K2���M����M{p�o<��+�u�7�޹�sň��ݭ�pv�-�v���"�Me�]���ͻq*X��{	�t�u�\�Jj���au��h�AMB�&,�����L����q�=Q�������6n�WU	\FZ	4C�3���֕�e,�qm&:��'����l�:��4j��\1�y��Ҙy�;W#c��VS@�ۗb��|�Y|���Ͽ�(�)H�n�p-��Q�v�+�����;�n����ʾ��JD��A�RSDx!b�����U��>��@;�hW{ow�"{�a�O�$���Я�Q�+Q[�})R��c~y"@"���;��P<IU|~JD���t���.��.N7�ynTK�c�'1�~�/��� ��D�:���}XL�� F�ȠuD�A�)|�����Ep���C�[�w�O{��#R��t	)G�
Jh�� �����	;[5�w���b'��P��[�������,)D�w��s���8af��(ݍ����رx��ƶ���=��%�6��3"�iA����y�/���u����{��a�����a�z�9�n���"�$_ A�� ��<Ϫء�o3��=�+�d���;C��`�t�_*�7���˷潪����fa�~Y�f��o��G��y���5���y]Q����~9q$R/���U�u(��4V�[�ǔI�$��.ʉ��D)ĐA��`dA%$U�ؼ���韞~�V�a6p��A��~ ��R����� ��}B����f;�ڣ�� n;��JD����>^�:�a�q��戨����Q�n����A��l�H�_IAd�,*Ҵtz�z����:����<+����Q qȟ�R/��K_oK���v'��ڣ��U��Μ�s2e�jx� ���	
n56�>�&v���P�:�8���D�D�R�����������8c��B��v{:�D�Ϯ�i��>�|�mCi[�Er�)̝la���p'���p�yu��C����9�A�"AJ*/z�N)�+�D�-�=׉�ܱ�ݠ���c�V��\|�};$�)�
F���/%<hh�ko��s�[-�j2efQ����u�Ӥ�z����^eU��=[��+]ޚ��b����O#��^�N�¸[ޠO(��O�$��	H��H#z�36`�׉��ܲ��H/`�ا���=]�M��N�	%46�ψ��	��`�D�� ��
�I	@�J��D?�)6�ć�����ꡇ��9�4>�#%|��+G6������'㡀.�a0�5�BK��-���:�tR���
U��k�؁���u�J@�"g��W���)�xW{"�{Z��8�c�p'�uW�)�J>�RSD\]go����
�'�.����{�xua�"8-�w`�"�J/+��>�f��,�喛ϰ���b3vˉ��0ݳ��c�(���7yN�3E�>�~�T�N�s��}�,wj�n����:�z�&���'�SY-�#�(W�z>�����qү��zS�����O(�C��g�۹c����m~9um�βW�^�L��*��Nn�u{�>�f�6V�X:�+Tحn^��>b�ڱ�˵���<���#�`����/dIJ$�����H)EM��1=��#}��͊�+]GQ���bc���Av�C͑E(�BR9vݕ�=Y�~�n���OޓDP�ֻ6:ƹ���1�]l1��1���M��H�q�Q�~s���O��p$��}_��3��P���.���%�q�s5l�oN���ڙ� ������2E"�/���w@޴�*g�Y�0�� ��H�]g�_w(��i�\-�P � �rI��E���>����?9���FJ@�$^v�3W�_VWb'8�1��bc�ޟ�`	6��I)�	)�Kug���ti���"A�_W�@��ר_i�[��w0�8�A9�5�$�����(�=�h�	(AIP�
Q�r7>��/dH�YeO^�(SnӢ�[ޯ�D�9BJ�|���یЊ����c����!m����U��<�}ڎ�5ي��K�\�uӎ&spwU�]�ai
�t�i�x9۹�ՠ�V�u�V�YF�J���ǨUQKA֌6��bŬ�u���p̻$6̧\�w.ɪ���aX���4��VC���s�{��Z��H㛹�����(sZ1WYܲ�Pn`޺�m��cE�*2U#;t��Vxr�mlWCtU��ͫ{�.��f��%Dj��S�R�˻�ֽTnS��̰�ݼ5ڢY�t�l�r0��r��N�r�,�uY&mmٵ�{`��ۧ�bʺ���e)]$CK���e����}J�޴77v�V7(�i�|]H+�ɕٗr�`Ǖ0�;7N�+�ViD����
�������r�דr��Hj�\;�si�Ұ�1�dU��t�:����ejCXq�/D})<n��X+�,��{1e���ʕ1�7W��;��T햱f#�g[j�!��s��(��YbkPQ�}��f���p������љٲCN��ZA[�pb[�����v8�D�"��1YQwU�M�����r^��e	��Mخ�=�ŕ�f�;m汆�E5ٖ���f�[�)�_bb���.��#�����2����]R�v���Qழe���4(�Y{�����n�=�R�2.ދ
⊮�:7.]V,W�Kgd��]�U�{d����es�z8����]Yx^<��g\ғ1$ۨVӡ�|�4���`wu��/����Yv�
����Ҩi�=��i���)���΂vLSfu\5�<;�UY�y�y���S�(����(�"��D:H�5Ht�I'C��%8YS4)�GqJQ� Q"\�i ��:	(�����(����D�J(�.t@�($�����̊q����$�H#��vA�$ĝs�Dq%'�E)@�D�%G�q�[YmY�rr\e�pw��E ��":N�"��8��"B�NC�S��(�	+��s���8�pq�Pp�(�)D���8T�B\"�.D��p�p�$�ptQ8T��E	�C��� !�tG �"�Ă'\�P�[a) �G>=x�?��j;>��n�:���一G�����ތ����k�;n�6��\u��t��˹l���{�:+b��.�n�C�a�[�/+��0��)V���Sy��g�\i�r�Ĵ���@R)Zj�0%�y��Jw2\ku�^�]F����n&�1۴{ҥ�at$��Afp��y�d�:)��VbX���v��5. �,�F���mrm(��3H޽�1ǝ�;�yR��MDI�.|�;=n��<l��l+��z����-���]3t1LRrn�+���qo�t
e���k���Z�����Ԋ8ヌ6^����m�s3T`����̫9�x-���7'<H�ܰ�Z:W���9n%/Kty�.<Zk�e��ۦ��s�+�ax�abкn-�j��uZ���q��Q��N���
X�U�e���;��i޺qڮnƣ�ܑ�w��/sUs��p@�s�1�LwC����ݢ��#��"�ˁ_
/8E�D����Z��{)u�OGh��ɀ8�%�ta�rU6�$�.ll�5�K�ƫ4�;5�F�^��x��o����8y��nR���[M�� �3T�W1���\���.qӀ�m���^r�r]r^ٛgJ.�eq�0�c�4m97Ѹa՜�ўw�=�۷1E����qVj��-�ڍ`�={k�s�y[! ���L���c�j��p�ۭ�V�<=�[WBgŒn�En��<'e��g�*L�ђ�bLsv���&�n6���P7n�	�.����.uƪ33�'I^��v�7]���!�5]�=�Gn�wZ��m�������'q�f�%B�r�JD2�
JLqr9��V.���4k3�^d�"�Z鲝1�;c��}j�:�h�<�qx2Q��5�P���]ia*F�t�6-)���J2s��]�!N���w��m2�q�ۭ�d6'v�]�C��U�nɚ@�==qOk��W�n�� z�=m2�<�]�A�`��%堡7>݈��F�{pi��Lt �ɗ<�.�d���Cb6�n��7U�e�uJ9v|���Va�ַ��y�ݳ�a�L��tJG0�6��v,��z�m6��	���kb�V ��ǋ��`y2N{{{s{���:���t�9Ҽ��υ�J'�Ih��s:��w�nň�^��T#GH����Φ�:�j�Nݛf�]��}���1��nl�r�����nM��:�tƮ�-���.uۮ���DT�U�.?@ ��&�]%������{��f�,zxf�W����P<5��V���X��J@�����P#b�\����g��)=|��>�Yn��>� �l�T�)B��eC�:������7ۖ0{�,D��0wj\�"���ǦU�:����R�v��߿L�j�9�.&��ݲ�V���v���U��ΐ~["A� ���{�sI���cd�xf�A�HK��=1�?[��:��A$�,%|�A|D���ݪ���	9t���D��fi����-ӹ���㙳@�5H��H �����Η�`�a��5h]�$hh��.Y���x���Xjݚ�����c�{��|#g�zE�H!)-S�ʷ;:�c�����:�*r#8h���� �r�u�P2R��$V���*����[�_J��.����W}�;4|�w�h���6����0Ǖ�Yw�Vg�qOeVqQx�y梶�}�|E��]]��GL�Mr�ʔ�}\8��?4��{�N�5��['��7����A�_%���CÿYi���7l�&��ݢ���5�֏�ں�!��1�d��q�͟�T�)D�JJk��"����T}�v�l���m
�I	@��WY�[��J����}�>��;�}6$���wH�R�?$��!)R��s�/l8��4}4�v����x���p��?s� ��"�Q�CG�k��M�'3��5航�&'�����&�W<w5��.����5��aL!�/m�Ap;B�o���H ��$$��JD>�{p�u��O=.�w�un��򶥐R�%�I����� G'��:o��T�c~�JR.gng]pM�9+E���Q$�$ܙ:�� Ȓ�S����`�@Η���dIA%|��-y+�Q����h�I�K��l�u&��Ҳ���8��]��Z�3��6��[O,-���C4�\UΤ�Q����c���ö��82�1g<�����bo=��9�����%�РR� ��I	)��K�*���2� �ޟ��b^�͸|:��7��]� �s�[��;$���{Cz$��?%%BJ� R��V;z(:�Ѣ�D���i��*�ݻpW{#�(�1��U_�����mGg��0�D/�I���X��D��7[m�j��{8e�В�d�zb�[��DC�g���.���/�o����������bؿp��u����W�wIj�x�ȣ�A�)%u�Q��N�^����w?P�"g���sò�c����J͚ � ��'�<�)�G�~����J���	H����w���W}9��o������$�1ȒT+┉)G��ү�;��=�4-��G�⒚ջ�7ǹ�e�Ng�f��p��jid����2�s+*��iͽ�����+��^�Eަ�]�ꕔ�X���u_�����3Z���f����f��OI��l�ܯ���H����%�@��H ���̭��ï�p*^r�}<;)�4�]v8��������(�W�+�������m��r޺d0�����c����0��-8q���j͆�i�6��/����F��Т�I%"@�Z/7g:W����Ez^h9�����Tx��[u_��+�H�W�����&;��=H�yɧ={�4^�9�l�p��� H6���m8�>��MȐF��?�I	*��R69��v���I{�ݹcr��NK����f�#\�(�� ���	H��Fk���A�Z�@�A	H�j��݌�����|1�}@�Q�*^= �OeRt�C�D��I�� �����	���&X�|=�A�S�>wø�8̦�Y�����H!�РR������7��Y�+���b�2.l�gk5�Џ�8U��68����,�܊\��ؙ���ѡ���S^�7��n�g9+�ӕvBR�}H!X*�5@�4h��� 08qS5!�� �l��h���3JF�ON�qU�&m��%�ƫ8�Ó��T[9��
��FͶ���u�%�{n�,�.�ղ��ɚ���`��T�ܝlz��ܷ<��<O�vig.t8=<�j�����l@ή�<-����ͳG�6����[�%���5��x�S�[�F.���w��?6"}Bk��F.�����-�Q�����u#4ec���)6��1p�AyA�����";��ۮ9�s��p"�rG��:#�)D��SD%2	J�k:���Fw��}�$�DڭG;c:s�^��|1�9� �9BJ"3��L����ߤN����|}9}%2R �$]~�2=�K7R��<q���Z��P;��A�РR����T(uj���o�?G���J$_H�u��H��u��}�ӗ-�0�G~/6h�ڌ��,j�}'���?%A%B�)C�\-lt{tX��J��q�gNpk�ۈ�z�=�$�I	*�2 W���ۛ����	��FR�J�(�bQ�ʒ���8Εк�j��R^�hQ��[�{���[����D��@?$��'۸�Gc�m�]?h��#ћ=���� M>�@�� ��H!%b�2R"~�%�K��x����#�6������Y��	�u�3	�[��p*:^��R7�5���oj}D�~��p[4��(���������5v�����_W�zD�뵯;��ƛ�u�#������$�����o�y���9���"A��@�R(�O��d�E���_��w�9��\c��W��#�{�P'�N���_%~(�=�ze�[��Q.D�Q�RS[��S��n�����=p$�^[�W��wF_
TH ��BJ��) D��I/a�z��6����
�w��{��9�×\�8�of� -�%(��JH�[�7۽�8_nP�2 �}5& ׷�ݡA��������>�ed���f{^�<#��JP$��O�W�(��"�4yiΜ�W��#���	>��>Uyy=)��ș�X��ّ��[�V�wv�;W���H?�tI���;�q���M�ן�j����B͡_�yy�\���h� ��_P#��>J�IP��R3��o���a��f�G�x~��C=j�����PA�nJ���j)[�ҫ�h:s'�d�Y����nG��[K4�W��v>߷�nӝ��ךܜ�e�;��y�q������'�R�?$��	O�-�F>1]�� O){c�xU��ӝ9̯SLG���'�7.�.ϫc�s��O�{�3#7l�ݫ�����.:�g��u��6L\S����������u�Z5w�	�?Vm
(�
R,U��~��7�u7�c�<B8 Z�G�v���W[vݼLT�^�eX�;C����������l�}`I]|BR&y�|�'ޫ�n9�p ����r�nw���t�Ώ���	L�
P�J8mL=�{�l|�l��Ml-9Ӝ�=M1ޠA��Ҝ�$����GӐB��>�� ~���%(���)^�>�>wV:���I~p������Vm
��AJD�R7��x�s� � ks���H��5��d��cM�wA-��"����s_L+��r��&s�Y�ۃ�����&�q��G1p]T���T��4�`��ˤ��.-y}��P3B��yU�{�L�
�A���JD��)@��!%B�J"�8_S�b��4���9�'������>Q ���%b�)H��g�IÂ	�3SP"�kn����ѳ]����7�%��=\n�t��[�$�� A5�h�������ח���r����᫄�ޣ�FU6��FvРZ�%HIW��Q �uj:���Ҽ7},Y�U��L>�z�vO�VI����S٢
r'�X�b��{��v$�8IH��I%"1,*�jۑ�vj�%��8�O��C{#����'�M���/��#;�9�!��Z`��D��H �������{G�ܧ�:y<5w�	�?���+}���'���!%B�)D�
R'�]q��>�?��D�_�OWg����&�mG~���'"AJ$�
J|>-�����Kwan]S��fc�)R��|j��΋ڵtj�bˌv~A��(z'���7��I�J��<l��ݸ����mV�G�{|��껵Q��^�?!=u���m�e�3GDaV-��2��2M�v�\�{MR��;�{���G�Ͳ����J�e���Ș�$pr\��9���c�?�}k �{�pr�n���˫R��[������W3$ƕs�ŶmCT��5ۇk�B��h�%�f�2j�m�k��$�l�����)���ڹ���^��Lڅ�����Y�|�C�?u���)���g��͢ـ�M�,��ݫ�Vk��3�J������b9�Z'��;�b!�e��-��9�3�m��=�C`�����vҍ���Gk�����}�Jk�5����o�;Ν��G���)��^jOk�S����'����@��+6��fq������]��9�_��I	*��JFG?h�����4��޿2���~-��A9�(�����H�^�Q�O����?5�(�� ��HX��V�t���l���}j$$-��1�:��+Wݰ$�H%%4!)R���`f����IoWT�Iշ��wǔ	 �u�Q�� �����������4ޟ�_-���x�P	�,�l�6��VV	(�h�oһ�`��V��)9�.g9cݫz�j����A�������mK���D������J�� �z��;�X�x��>�yKSos�֗�v:򦨌�����H�Ai~6�l����*���ٕO&�t��kh]43���Put=�Fk��'�}"R�.��9���c�n��j'���� fz���9����u����A+��&�ɶ�E�qS^Y�=)�um�'���O(D�b�����$��9!�_��nIU�P�U�	H�\�{WR�X�I�ڎ �g�+I2}qb{H�w��$HR�R,�ZȯzyW>����s��p[�8Q �H�U�|R�+�N���������U���_ز�+(�F��Mc8���k����B"�51�صڊkSK����_��O�5Ȑ
Q JJk�~j����ԧ6߲xj�!zEX~���� ����6/�
R$��_%Gy��;=R��Y�R�+�܉�6���]�^��<��%v� Cp$�wX�'p��*p��y�#7w��Znф��ۻ2��q���x�{�8 ]έDޙ5mv`N�}�u�@��cu B^�7�8b.�j��%f���3O1�u�!���q��"�g��"Z:�V�\ݷ���f��uppȑ��B�ӣw̼G�]�	�Fk��]n�U�ףs���F�N����h���y�b��cS=�N�4Ѻ����86B~���'/��]I:����^+��f���$�rՎ�$�uQ�Jjwr����ko0MB�=��z�����1���a�
VR+x`�KM<�Nffh�l;a�*��&�)k!�(�X,j�-�̭�JWm
k+���Z��f�ݯ���"���/.¬�ri���,@s���1WX�v!���j�'p��{�uS�U��M�*%n�}J��Y!�->�F�☮�"]�����w�>Q��sꠎi5շ��e<ζ�Ev]�Vc�R'%��ОHM�k&+�\�`K����9O����[ZMt��H{kQicuU���E>;�%EՃ*�/GSh_�0�7�J㽛�ɭ�Ɔd�6����P��՛٥�G!s��r��q$QĻp4ђ�f)U{C+IT�缢ٰR��%nl֖����ΛV��4̨J�{���Ն�:�[N���o�w�1�3��Uh���ۣ����q������5�,�C�P����n�N�V�o.�c�#e��T�'&U�ǺZ<�֌��U����ؕ�ձu���7�h^��+;�E��ͮh�Uj̵)�pVz�F��\%�e.�*|u��i��(*ڻ�)��������S{T��/b�PD���"�:��C�);��.p�!�.p�98�D����8���莜C�����N�:Nr.qΊ �JO}h��H��ۢ�)I.NN�N8� #��	 ��\�Nr�:;�r!%#��ΐ@8�):rH"'�RA:�N���:w;�.$ ' 	p������D#:��(�% $t�q8�9�� �˃�H#�G8�C�$����N��N:B����q$���N9%�ItBum����'9�	V""*Ň��3k�r����y�!�w�j$B��	*�P$)5��'�i�A��Ԉ&H��ޘ��yҔ��������ңg7,�5Cە��3%/�>��~�A���� BJ�WZˬ5�F��u$����갅��mGK�!�R� ���g����@��4J�_q��ˮ����E2J��hv,d5��,�g0܎�C������l���W�(�@JD⦺�_W:�?d1�n���j!�ܽ�uW��Q`������"~)D�~IM'��OdRt:&�D�����f�n�O}<�Jr��G\�y��?&�P)Fvܴa���s^H��{��x��W�%!��m�t��6m*��֛�O�`����A_M[�%(�A ���]�^�\}/���_b� ��H�O�-˞�~�+�c�{�	��64���n�s�_�EZ.����X<j�Ggi))��JF��,n�����l��뼽��Y�v���ɹVҝ�8���UI���ُ���CȾ����wj�1��ȉ�sv��x���}�6d��ON��%�sʒ�k���H?p����� ȇ9?�w:�N���V0��@����B��]��j1���"q+�jF��+2�oO~�2w�h���ws#7dLN�[ټ�3�-&;j>�D�[���Q��f�H:�H=� JJ~J�(�{89ϙ���h`���dZ���s���J�1���_b��t� ��d�]�J����txA�S�|��(�))Y�Z�b�j�;�T�CY���H+
(�(!%T'S!�ؾ�Ң�d�!����JD��ս���>�&�c���_M]9ѾP}�Nt���]?fl�
P$BJ��U\I8��wF�ȟ��w"��<��%Y�87�qD�~] $�
��#���H��c��Uyg댳<*�:��<m�6�Jޣ����SF��*�r�Up�i���ge��v��q��w�͜*��s��������T�����״���ۗu;
l��������B2�8����iM�V��E��1�,T*m,�2f�5l���4��4c��i�,�f�1xͲP�f,u�q��r��Ԛ�&���ܴm�u�����m��=��Ka�Epj����/d� ֻAj˒�K�]+5�:���ѻd�d�h��ed���ьЍ179�����>����F�t�f�FֻN^���FQ�͉�J�2����4�"crc��4Ag���RS��/�t�T�g��E��r�I��3o��b��A�D"Iv�JD%�O��My�����<���Wzc/ �Lv�}���-ȟ�P����$m�z���@���@!$����De���:�[p���9I��	���yt����W��IJ$�w��f�}?n�ώ�}%%41�X��G�&ee�<5�A�AK�.��f��q�q$>� ��
�JD�A|D�āu�Okݟ!m��s�za^A��ݨ� }4-ȟ�����{c;�O��'*�&ţ�(��3Y�Za���Cb��N�)�ۣW�y�m
 3[@ ��_%)H������_�R��{�+�J\g5�o(�0�V���_X�d�?"�އ%ӯۡ[�V�K��=���-�dxD;^��w�C�	�r��]�M�R��;��c3	1��K*a����r�o`�ίS�:�B���H �Κ�|�=��rl*�xxk��H+
)A޿h��A�R�}]"H�l|�S��O���;=V{�;|�]�y�c���_Mr�H��Y$2�?�;5t0�x���!(�,�e=J�{ةF1�^�(���GvVO)�zаGwU|�	 � ����%(�w|gjt�=�M%5���\�Ͻ�������H ���)D�A	HΝz&u��KD�-Z�aV��%ۘͮ�6u�a��0fk��.���ծ#Fc+=+�g��ڸ�{�-7v�|�	'mv��ޥ7�m&;j8��}�S�rz�Fy\�A2EdH��J����j4"J6<u�v�����Ww���b�cF���H�P�����k� ��n�|A	H�R����IL�B+���x�@��M�W:��0�.�rmݎ�ޥ��u�^É�ܚݨ*\�tD훵��ok���no����6eKz�/5�W���Y����h�?{E���p�ݫ���Zn�a�e`a>�b��D���E��|BR&'mv���Wu�m&;j>��� FB.�D-�݇���~mM BR$�P���E(�������E�0y�5�Շ�;��+�cF�������@IO�@k���99�b�Q����ߍ}�,��ܗo�0M��箅ʑ6嶙*��L۟��%�_��:K/~�"JQ$RSX�����W� ��磃|$\�u޿[� {��
�ؒ
RJ�|�H"fн{�칳	S�p����v���3�V���������IJ��z�~�w�^D��b�Qb3wp�(��?%"Uo*�G���nv��h���sI+�c����� ���%u�	H��U�O~��_�|����A�K�	�*�b�j��ʵ�'>yQ���$N��&S�7�aεr�=Q�M��Rk�J�����1�z��-�$ꚦj�bK~���g`�˪��f�ߩ:{i>���(�UW �D�� I]
Q ��N�h��2�=��y�=K��VU,Lv�8:�~����RS՚�J���*�pG�0���h\e�Ҩ�,5v�g�8��hE�ʝ<�(�˼�+�}�}�.���`���BP$Bε��{y�,W8�{�P��[���W���Fy���ۙ�e��b.� �k]z$s�g3) ~}�������Z�?<���	���A
(�yz�׽����H�E-����%"A	*�P8E�������K��ʥ���G~:�k�A���(�?$��J~���f�z�𝽁��Α_Q?R�0��pw��qV��1�^�����t�ڕ�(X##����d��2Ed�R���c��Ӌ_E�����]��9����H �������������?~*�W�o7�4��y�y���ug�m�R��j����g(��E����������5�v<���K���}v�c��YD�u�1~�ǆU����E�+b�x}�-��0��<�y��-��q�q��z7o�z�b�۷[�Q��z���q��A�0Jv(���qr�qm�lu�e8���c�e�v|X�=/T���wV��ɦ%v��CF���R�^h.�hݸ��%��,��7���7>G��+fe*�M�Z6�f�h��PŹ�ݯK�z����-��tv_hu�*�G������.�x���W��:�k�{mq��n���^%ܝ)�H�WtR���h�A�yC���"�^���W��*r�Lv�;�0u(ݐ�(,vwWl�=�$�	IO�G�@Dr���G��l���k�����W��<�@ ��$�����xԾ��{�A�wM A)
Q$��銸��[ى��T���~\���&x'�Oݰ'���W�(�R�$$��}Z�{�6��d���+��R'��{گ��*'Lv�;�A�B���ʟz��X���;q'�4	L�R�$�
)A��짫�¾͑"1m杼�s�V�q����$B�BJ����H��~����[g��4�Vl�1�9�Wa�����&� �Me�=�V�Q�r�-_�'�e��?;��}D��} ��U��v/�6�g�}!Q�udV�{�5Ӂ�A�B�tO��"����ֻ�J,U(r�c�p�ߡ�=�nX}O'W��W�0y�puO/=ƒQ١���c2n��n}�S#ޔ��]�W��H�o��ܾ�31��c����?PnD�R�H��~܃w��r	́ ���(�AJG�r#A]g�N^Z�9K.q��Wܣ�0$��q񒾰�Z�U�[�T���I݉��R�5l^+�7�3�����!���_���y<{H{�D$����AJ@Ib��C��r��6D��ص�_g�3��1�Q���4N>R��$]Y�~(~�~���
T���4��**lͮ�=YS�s�Rika�.+��e�cݵ�o��dk`O���QJ$��OЫ��3{�R˜c��!l��~��6�f��WH�u}_�H)D�JJh��^�1~~��B�+bH'7g�歋�|����t7�	�A玅�QS�+��<vg#C��!�v	������"�Ĉ{ߴ���A��z��5��^^u鬤R��5v>Wt���X�.x`�?Y��;z����B��+q���Qk�]2�=���k��j}�y�`�Mq���x�Lv�q�V��ND��H%%4BR$<�S"����� __����R�0�;�w���e�1�S�@��G���]�~�}���W�+�9ȟ�Q����)
Q��]4��ܗc��|��m�]7�qi�T�o��O8?<t(� ��]UX��1Sѯ.����d8��&*�*�+6Ӵq�<ݱ�Ͳ���[�m�U���J�y��?���'��"HIP��R=;Ow�;+���ݨ�"�&v}�e�� �Ȓ�I�%4BR�
P$��K˄}t=}ӣ��Ăl���E�gw�U�Xƍ��	�H[ $���z�z��^�="O�A �t��IJ>�RS�����VW�y�t^-�!��S�>�A�A�_�~ Ȃ �%�������X�2�>�/��m
���Oޮ������{10�j8�
�4Cy'=Px�5�s�J��8�5��uJ��H��mW�v|��v�ie�MLɪ{�'i��y�^�L
�I{Ϟm�Eĉ���]��p��� ��	IP�R����b~��1�����{�*��1�q�GҶD�U�|R��Ҍ������ys�����Y�7�3�ZA�̠G�T��ѡl`M��ł8�[��۷��������҃���(����*�~kؼ]x!'�S�>;V��՞��oʅؐAJD�BJE R�#PO��L{��^Я�@����nu�^&�G9�~j>J+�*�p���3����H?P$�>IP����?H���=;=�����MY��9/|�Ο�O��#7�.&��ɻsv�H���g�ò���L�c6D����	IM �{{^ťׂ~U<� �y������x���V{����I�d�"D!$�ѯ�b�h�z�p-e_>�M�2���P~�_��(��*�y�_�$�BI�!$O�H$��	 �PI �����I?�$�BI�$O�@!$�`�	'�H$����I?�I ��В	%�I<�$O�@!$�!$O�@!$��	'�	 ��I ���$O�����)��<9��4l�0(���1ύ���@P�@  �%
T (�  
!ATJ�P PJ��TP *��H�P &�  �IP�� U
P�U *�R@P��R� %T�� D QJ�B�E
@
�@���* ���R
IR!J(*�A*�B��D�P�ED�T$���U �P�U)((�%B�"�  h�P��@�T� O�C�
7`��`�� 5� E��:�����b n�T���r wc��@
�|  ��� c��� �n�u@��₢��  tx��Hp = ��B��P /{�t���((��s�@� { @�  =�"��)P�"�$�UE8 @ �h|� P�������V�:P\�[���RnܡB�Te��.�Q#��6�(q�J*�P ����}����J.p�L8Y4E7n����T�E�㔳T\����UUݺJ� 	REx �U"�T��@�UP�%{�+ �U�*�\�Ҝ���PGT�gJ�wa�K�J����;�H��;��)F6�R��O� ����zzf��ҊK:Uw*�4�j���7{�Cճ� q�U����wR w7��{�" �PU �  �R�@H�IQ%T| }n���Q�	F-P�M:\�P��w3�)Ww������i��4�)Q��1�@b�%QE>   7��ɠ"}��=��JJ���G; ��A �`�qJ���� �А��*���B�@�)�   �!RH Q*��A��� n�u@�@� :�ʂ� 6c��1���!�� 	s� ` �� ���B�JD�  �:�� r� q�	!� �� d v :70 uwRT. :�4 r@2 h7`����E)P  "�����   ��T�ES�0� ��R�A�F�z��S�4d��F�j"f��Oj��4<S�?G���z����$�$<<��s|�י<�<��HH@�\��$$ I5		�HH@�~���	'�$$ I@�HO��O������Z�?Ҍ��2;�%���&B��E)���г��w�RY8!�T�r�×��Y�m�-�mM�0����W�Lnf�V��Vд�Lm�̪�xi���񷄼��JJ;d�C�t��aJ�rl��h}���x�ܫ���e�v�ܒ+]l�����P�],:[:�9G^nMt�!k0i�ڄ#��X�C���!v�-X�֮&(�����F���5Z�SԲ���Ι���
�ۭ����N�!f������hȝ�-�)��ZU��qܳ��ݸAteDK�a
T�YpfF3P��2ȡ4Ԓ���Ú��.�cZhj���v��X�$۵Ke*Ѷ�X��6V��	�/YwG6��k,���Q�-m��gqUŲ��8�)z������È݊����Z��q̆΁t�)��m��!&���w7J�Su����ɚ�n��S('��P��Y�V\���5�[�-�'t+i�"�{���feh�� ��)����st�7@m�fY���ݺ�F��[A�Y.غ,A�ڒ��R�g�p �DҺ���7�ے��Y��mBrQH_� �߆K�p�S%ÛyJ"�d{B�:�Ц��5�:�R�e�!Ӑ�vjjZ(��ld�5�
��	��.+]V�Z�N�lam"�1LM/T�F$����Vl��{D��xȫ�u���廄�qz��w�W��.�"���b31ø@�/fU�YB�y���6�Y��@�ǳ.�Yffv�:��B��=����XZ,i�$����ę��F�y�r���R����EF�̬�&�w��ٸ�V	qC�y
-P8D�����d6[�&� �S�{Q4HM̎àP�V�R@BV�b#�6/[�Y�����RP�K/Mܽ�o��=�ߢ�*�Ռ������/��x�Ji@�e�Іɗ���Yi2(L����;i���ƛIK;�j� �2�i�G�R����1�# ��)׊TM��ͩ��Er�EQ�vpR���3a�N��y�6dP�6=A�ܬ2U��هYuC>0VK��f½l�6]�aб�9�?�J8�+ʗ�p9{3�gv��#m�̠�e�+I�	)b��ӳ��*ǎ�ʇl�Wd���a�{2%Bb ]ef'qe��3k$|�u�D�.��h�ɹY�/(���Z�^�B)]`s/$]�~us��3�!�EQ"�(Ԧ��4�Mʽr��Hen]��*��z7�键ڲ��G�T�0^"�"���)��,Z&��h�Z�r�;
7B�>��	;|��Gz���`�a��'�Ö1���rj.B��y�wQ�37Y.ܱ�6��1(�i�ha��7AV�̈��ժTH��ʽ^$��d��nX�ˡ��,��k�5}�mԣ�U�Z�q^��w*}lLZ�����b�t�̦wi��$i�na�� CIlfލ��l�ݵGY����RjܦFlR媻��;m<�Z�#�swN�V:�3sMb��J���0��$�{����8d�wm�Q"PӰ�)N��m���nlt�7���.���H���[����Fnna��q�ɀ���g"$�`s!��!L37�v`��V�K/�� �L\'p,D���N�y�:����$,��HwVE�N���+nV۠NY�hm��c��fnC�B��i8��\�y��3�&%CE�jǛ�&��	����À�j+ǵ.�q���X/4`��`\�0�^'���L`
��$wF���8�:z)��;��=����ݹ�ԩx��*W�{���uX]k�-����܀I(]f�fM�Y��zɫF���y��	�2�1<���bm����x歫���F���p��AK1��]B���q�M=���tJ�+Vڶ�I����x�i��B^�Lcۧ��1�����mǹ[��vΨn�Jy��������Yx��v�k��vC���ʏ�r�=̋��{����&�
�5�ư$ ڋY70�w�7I�z���V#�w�la����c����R��]�H��r^�[�TZ��x0�r�'	��.�ͤ���m�i�����������*�«'��&)�����e,���(^(152c�*Ľ�*������?]��Ag*汸�V��m]KܕiL��fT���)������k`��qZ��@���Q8���>W)a��mX[�eeC.��t+3H����U�Qh׎�!�+�w&�Ѩ�E��#U�댼 4lJ��ʣ��S7�����e���)�K���8�"�y9s�K�$J�M��uKE
\ۻsRSYe���I��*��x�9�ة���0\9
����	�7	�-�ے�&����lB�E�K�cg�	�Fd�hC/�TM�Hj2�E�qM[�p�FHd����̕�@xܗ9�P�Aؙ˨755�:��d!QA`X�.���u~!T�r��s(�Fn��m�9-&nX�U�����]�E��QS4��L<�7B���2�@�R����0��v��\ۋ6e�U(�/��r�r��6Q�%�Z�5r��������������U���t��:�Ao3ugVX̣c0��V�R�p��͡�H	J*�S\C�;�ɰ#�gsv�w���U�<ƞ]��
fiHe4���-�هFL��1@3i^+4�*�Y��Mį���.��f��xL ��p��b�m�-:���@ω�1�$�u%v���R����U4ƨ�)�X�֍�j�i��1Ũ�B�Cu-&�jp%2k��A���2�r�n�q�`���ҷX�d����5M'ie:�(Sk
��	dGc�x%t5ύ��	yi�'J;�W&�բ�k�p(�əvֳ&���%Ԣm��̚e^5�7	� ؒ�v]�iZ�*�¼%��һAL�i�(04�fB.�BS`ߛ�TY�\kZ�w36f���7km���Ac I�X`Zv�S�+^з�V���Gu���`��5,3���`2�Pnjs�$�毱�o^ͺӏf�"0��te]5�1W`��f:V��՛�#�9g	ϴQf�XxcK%���	$�6^/fe�cXãb%"%�6���4(���KFV;r��6Jv�خ����4������%fnjS]ݨJGL	���j��w@�*���aGp*�.7�,z�\�)���Y�eZ[Z H摫�KͭB�Ǭ��ۭ��fϙآi�n�Z4�LLvm^�Ȱ��M����MVR�ÌG�քbL�4`ye����j�s4��p2d�)e�묧Xkk�y�s,�֞�ƶ�e$f���n,�!:��L��O(�P�!ʔc���~��Vn�Mɸ���뱪�j�5&�WBӚ�u�L�6LVn��*QY�]�&�Җ=��c��F�ܺ��U�*J.Q�
4۵��d��Cd�0n	m�ӓ}��j��i���M/�Gt�G�;HC�*[�Y����ܔ�w0����t�a";���#�XL[%�uoE�$�E�n^��uv�^`{��#�Q��z�5���W�^�k�l=�k��"[9�B76R{�^�5fj�*Y�����&;��uҳ��.���1>�me9�l醷6[��RB�@��Sȹ.Y���MXLDMz�cj+/E y�O0���]3K.�V��sv���� `�"ם%)�Qǈ�Z��ܤ�$����9�oe�((���8P�4A�[؄2�R�3DJUf�k��ݵr����Ov�e�\�X��L���������R�ـ_�)[Ϧ��r����L^��Kd��
ųY�U�R ��Xd�f`r�*�̑'n^y�pha�vK&o��L���V,��veJ�L��K�06��Z�ʚ��;�cYq䣗�^���båtd�d6��j�ݐ�~u�f��'XNt�e�f����j���4q�g��(�˻���(nU9�%)P	3����'�F+����4�6�u���[6��L7���[ �n�D�a�Y��̻��L�n�b&4��xwww�K1�@����O��E�����s�(�!CJ	����kL�0^*ݔ��ϙ8�a�.[���[��՜0�.��F����5`�e��^m�+d�hF6f90Ebh��\��p9�!E9XV/c���s��@��h`���Ө�p-�.ع[�Qh-�ט��[!v^u��t�`�����6ҲU�`M�*��0V��XFV4�&�;%���c�Me�2&��^]^n�)��3S��-�w
B�sc"�8V��76�٩kb҉#
���n&�����T��Zum�T�mգK%�%��'%Lˠ���Q�.,�Ȧ��n��wRK3N;y��w�*ѵXkg%X�.�f��1^D.KH��(�Ïn��b���y
�)�mO-�-ڲ`9�ƪv�L���/
1a��յ�O�o9P���1�f��09��k,�7h 7�¡����n��|Mc��Y���.F�f�Tz`�&��XՓw;,l�6W����pdӧI�D�ɕ������øu]co��{&�6f�^nJ���kYK!��ZԎ-��>����*ڊҶfܻT�R��	���i*�]�oʱW�l���mf-Oj�q�@� �LǍ:��>�jۈf־�滞:̧��d��7��6b "h_�%Ey7�tf�"��O��ᴶ���*�S32�ޖ�mܸ����{��j�b��J6FҘ���,���7PE���\�yW�X�� �$�h��V#�LM���(2i��O1e!9)J�rf�F�����n�-)��K%,��]�b(S�O+�@x�p02}�.
2��a�}h��V�,�x6��n�]���e�@5���L��je]M�/32�7[�rV��(h�d�y[�z��Ӷ�KW�>ʕR70����*d�Uҽ�ּ��<���ȷ0'&��JfSQR�<����+pf�Q��L��,��k<[w�ඝm6�-E��E���a$]5^�r0�r�8�6R��u�R�d��rD�P�reؕ�7h�U[�P���<��wv}.�t.��?Ss�X�ו���vͻh�F&V��5�vb��LU�^��f�Qח�R�Y���a+�D#.���L��6U��Jܢ�k��ō�إ)���+�!�yM��4a��Vl����],*)AP~FbBE�]�u,��k!��-�"�.����ԫ���k
ٻ��i�G/�,y+ �f��M�nf{f�ͥNG��xqPj��5+��!n�x�k2�Cc9�&��l*F��k&Pmޜ ַ�M�h0 aR٫�@��*|�}2���4^k&��oj=��p$]�d�j1V�2o�7�,��\*�bZ��Eµ�i�cA�+A)6�b�nfi����΁��]��S��/l$nB���
���c0���e�62��HXQ���{
Ӫ�i7B\��D�V�ڱ1��$V���b���>�f���K+0��kmEL��Q���%lYk���$��fM�bRm�l������ۺ�-�؀��6Dr�귬�ۥzR��.�@D�&�vq!�]�Ǻ�큌�^�wJ���2��)D�!�7T�&nDʺ�����$���%��x[�&b�j7Y�n=o5D���[�"���i�Q�̂ɰ���%������V6^�ڵcY�6�feF���ܘM=1�Sl��	f���z�=��x%�{���b�ni �q���t]��)�^d3خ�{��[0�LKp՚%���z��1��h�E��Qb��B�ߥ�%*�+J���Ưl��n,-�vKY�n�&&�8��෗���j��>&�ȂsE4+2�dV^�tl��5/J@#��8�l$V��4�ڛڈ`�5���k6�9A�.
��۱�a�w�!b["��3�7�T�j���uw�f�c(A����4���ӻ0(��J�%$[���%b^�ӯ]�G�_�է�-V`�70����&f�J4j�j��h�f��2�*�m�w[H����`��ll�,�z���LU7r�^^䡆��2�
ǂ:ݵ%^f�C�Ȫ%���R�V�V<���X�HkpXu��Q�$ʠ2�/l���nh �
�(��"k^m��ř�X)hV�2�,����8�W[c"�XƛV�	r|j��)0i�E5u@��9�yII���`���yWI�ۓK2������$!V]/n�Al#Y�ݤ��sn�-̡��{@ۘ��!�7֞7JQK;x��� �dʇBX�xE���ǗKmd.2� B��4�`j.2Ki��cʚ$E����T�(¬34e]`QSR��U�� �bYĤlQ��+�ͧ��!)�wN��V%1�kM��q�au�?����B@Fd�F�8�"�hau���T�]'m��S�M�w�T�䣑5V(��Pǰ���V?����(Y�U<�&�;���fn(�ʯ��m���2���y1;t�V�	d���b 8j�h��Y1�zY9��g)�A�3,Ї�����A����3�����i	n���YW�7�dt��(	&��@*��V�ˠ^8�E{0�z� �a��
͉�e;�q�K�40Su�V���8XMld[����}@ZZwVf�����ܚ��H��sS�9�!��n�',YC#�mM�40E#�H�$�3@�W-�[Mjf)�3fc
�-5.� 3XY�]md�V�FZ����7e�e�����ov�{����#Mq�xE����0l��ڼn�^&���*^b
]�y��:���l�;��2bXJ�˧��B$�8�s73�[4�"���WwyWzM����d̆�G`����t���!��^^V/�b�D"���&|�2�dN4d����\ْDu��\��.�����@� , ���TZ*��Z������k[cj��j�j-��Z�5cm�j���֬U�ƪ5mڍ�Z��V5�QZ�j�j��kEmڊ�UTmlVգm�[[���h�Z6���ѵm�mլj�ōV�6�Z�mV,hڵEVūlm�X�����F�F��[m�[b��Tj��URZŵ�X�UcU���6�ZѪ�j�բ���F�ص��6ڋmEmj�m�V����ѭ��V*�cUF��-V�lcj�-�b�TV�6�V�5h��b֬m�_�mZ���ݶ��m�D�s�~�Q�̩�U�R�iѕw/wd��r�P�r7@đ �^����\�-P�&��sD����D�6�[�V�ugl�P
�pN����B*L���L� ���ֳEVL�u�N��;Wy"��%�G6e��k�Ʈ���~OР@j���'d;шD��'l�q�tTn(.�+P�G*Ur,�l7H_�5{'4iq��l�*V��Z�PƂ��G�7�'f՛�GE��Y�� �
�����fv�Y�Z��D)��=x���S,���ݒ���\��.͎ě�Eۿ�y(��lmE��[5���u'C'*B"%!);�vn���WK�q��d��Mi)�є0R��;2��d�c�ӹӸ/���5+^�uaј���]$��p�OA�gq�8�5aC�"����3QHM�Y��m��x��f
$�Jɜ�g���(��F��D�/��u�NN|8#v!
H����r���l̮;���*'�{1���|�ͧG[�X��ײ���a��bTd"tW�Cܘ�J���]hy(=1a�ݺYY�:ˌ*̣�m'���yB�*kE$]T����/��H*�݆fe���$:6�Y���'+Vs���R��H�T	�zy�]U��۲�z X��Z��j�k�`�A�Ӫ��YYK'$̖D�Y�ǮAk1J8zwtL�>�:�=vE�w]�9ٺ�`����=& ]����4:{�"sx����_]���Y5�)!���'�2�*t�%2u�cgv;� ԥ
*��u�5�Έr����kdS/��̦��İ�Đ��V�k)`/3M͢H�h<��/��5�e�J���ed55��-(�.R	���f�̮ۼԻi���[�*�Me i��n�e5�6/��-e���9]�X{�v	ZY}�f�2�I&nZ�W�F�\ؚ�vC�،��%�qoQJJ]�`J퍠m�6�k#
��ɴw{)�lQ��M���E�5M�:1�Y]e�f�7�+-��DX�3�^|6F�k���˻��������|�n����JXM�{� -�w}C���^;���l᙭�ٔs[k���IFd�ݹ��p�5z5�	-�]^@Ffb�VC��p�Ǡ�����;��*a�G���tl�
Ż��t<�f]��d֢W�;	}B2�J��^��r5�뎬[[������CO:1�MƇi�f&.2��PJ�81�b�n�[|:���wd/\�'ld��\z-e�]���e����؈�Vb���h�dU��*�u�{�15Ҟg[��[ݭ.�M,���/���{'V���4\k�[���2P��gƘ���V��ܑg�۫�4n�yN�Jܖ\�#l�U�0��J�z��L�wz��b��y�v�F6v��D)��^;�V+=��d�����vɷ}�Էb�h5���.`��>q��,p�
j�qQ�FX��2r�_'{�)���+[�I;�Bֆ{���p��r�����:|V�ᜍә�Y�����]�<��q98v�����)H[����Nω�H���㚎�E��A��]q�@$-v�d"��=��A�+e�2ýܡ%�谥��4;5��Jqb�9G/a��r)@�x���GQ�E��}W���˦���{�W�X&�F�kٳisi��Dwg}��VQ����Ȝ2��`篆,}���� dc0`��R�H��M>3��2�ȴV.3�)��2��S����ܫ��%,������,��v����E�X2�)��sk,7�)�1:v�-��E�6*��q�Aʵi�"T�i��P�VNi�W:J���;X<V�t�>b�w�eJ͝�d���a��Q�K뼽�k�s/�2RnV��]�RjdD̵��Wa{VvңRܟ�+�nq�%�b#1k"��e�2�`)�yR�f�ͥ��e�<�C ���fAmg!t�}
y�=���\�n��;~��BVV6}P�[q/,"�jS���)�p�IQJ�}��Y��b�`��k��2=E�M�e�r�X�t��RK]�Wu�`�w����]U�7�ȃP�mͬ�*�&��.�r���^3�m����v� N�V�y�a�ݍ��V#1й��*nPOi��Y+2�E}B��=�u,q�M������㙃tQK,JEȹ�Wǈ=�]�
�q��,F�WSR�gB�<
����ogP#��
��K�ϡ#�����`��`�#�$�ҹ�7h��]�α�q���X&A0�(�D���X�P�W`�ŭ���s�
�}ˢB�j8�3.���c�]�(�I�D�l��
��9�p��ga��N��εt�+ �����m-CQ�9O�/�}m�x��	���=��&9#���t�Ѿι�oP�{�i�hLz�y����l���%��H��$�^$�m�{���h�9��{9v66���ӫ ut�{�Vo�.�/#i���!��E���L�܉��"�F�����ʗt6R�l�y��&X��˹�z�H��Ll=��ǳ�PqW%(Ocg�#�xfͷ103a9V�1����˹0��J��Qp!L|�ʻc��V'�ݗ���N �&��/�NK�!r
y;㼣K� !�W]a��I.�@��u�����{*ũ��ub�v�p�@KH�e֍����u��\�����'+��%��۽����:ᦶ�W��`(��Zt�*�yeN���ͷ�M풥��/)93���&�7Q�}��z26�v+�Z�b���Ú݌�;˼ͧ����^w0h��(����K���n�8��.��v}�ؿ��B���m�J�3c��r�(�uzH4ξ�3BiQ��J�t PhI9��*/-��F�3xWw$�T�p�CC�6,)������V2���7�D7��;/���}��;��W��a�Qe�vZ�A�N󺵞|�`N�6����ž�-���)��r�g_>��*�j�Nhݮ]�㛈�uZH��O����R�eкX�'oshVc���;�-�l�
N��I�r6����ז����?*�t s��dF��s�+���%ΒwJT��=�hd�nv�j���൑k{��|W	^��!볚��P�v*�	:҂��8Y�D�YW[2�ؼ�s��k��^�S�c����ص�Ֆ�
�:��۠�D�V%���iT&^����ѹ�ǡӛ*�ñ�ÕV�ebV{,���E��Osn���ܨ�EP5/f�i�:l��"N��'wQ��%,�=:/��$�I��k�N	ww����+��ٛY��
�3v��8}��e�����V<�7���wJ7#��,df��}�i��漦�9��7!Q8KN}�9�#4��pΒ�5aI��n��:��q��ܵ��q����/�<�6���zn�{�20�����VUe#��:�_m�+M��٪^e\2�Qd��F��0|���9(�<�	��Z�r�ػe��t����֐�]Y��gWG\���)l/��C3lE�.a]+.��J��ʚS�:aE�fV�ְJ	U��7��ȸ�@l�6���rкahجX�Gx�7�øo[x2��]�*Ww���T:�ܗ}ur�$OH��SG.IR3ۇeХ46�<U�䫠7�Sg vh���đ&���λaQ'M6"��"Ҷ�.��P(M[�D���ٰ���-?���
4�=�+����v3����xU��nP����������n-e�I��m���л��f��K�8ln��J�ڸ�B��kK}ˆPy��&��݁��@�ӧ1v�x��Vk$.Z�uR��w>:6/�c��F�ئpI|^K�8h�Z��b��؍u��Z�y;��esC��
=��#ԙ C��q˵ϖXޫ�}9mV��w���7&�5.����A�-7ٖB�t��-t��3Vz��Ҙ��w�;7)�4b����2wVv��-И��c
���
S��S!���`�q��*(�����t(V��zN^�2q�'�mJub�����,#�qX��aD���v)��.�s�����+a��'P�X��<e��\� 4�v��r�,V�ͺ�c�W�:�s7�30�{.�o-у��ѓ��{��Jʙ�R� s�����-]���Cr����r�t���7t�|��*�Y�{i��&qyq-��5\e��\��ff�T�A9/npN֘ZۚUR/6�1N ��ᓈ)4q��2*��Ш)�h�Z�CK��R�$B�v�T��[��9�֑ҩ�Ķ�[�*NE���,ԑ"�FӪ�4�Lн�i0b�=wxz�%�FEV����W.q�ivm]D�2��(�����Kne8ϣ.noGo�)+���kQ��=FS͜���j���J�ge������vj2�,Vj�jĜ#e���m�7;�fƬVJZ���}�+K����P�w�d��jЫ����;(��f�ꚝ5�j���q�@m@"�j-`��������yV���,K�,�1�u�\��fZ�xv'�Q>e��5��Qj1��l0�X�e	�q^��0�����a�˗W\�n�
�q�ʡ�4�s�V �;��T��P��dɊRX+�R�1d�J�m��w�p����K+L�[8��#�9cYI���U�p�|�7F+��z�pm�7_>�ml���pKj��Pr͜
9�����\��cH(��jXY̻tfR�Տ�ق���e��_L��\����4�lcT�u�_!���cZ}�N�o`�l=v	3Jޚ^�MS���ͩSU,�����ֱ�e�.f��%EwwE�q1pE��(r�P�*) G-���^��Ύ=�y��l�-�_E�� ��f�ǚi�$7r����=D�
�#�D㮵SF���N�눝��B��fU���v�����hG]TK��wrnf�X�fi0�*Eش�E�x�L�l��L��sh+ȥ��"����ߓбFń
ݻ���.Ҹ����[��� ����� �Ro�Uk�����k�fa��݇F�kv�ٓh�5w1�[oJ0\�pkٽ��¥X��Y�G�y;]��
��h].I}s�-��
m�����љy��T�sL@a`�؞�y�)Q��Lz��3O`uisfPrm�J Wa��u����ѩ8���X�kj5�V*��$��ܮ'+Oۃ�M�A]f���3����f6���
H����)llP�	(Y�����ۤ�1�ɹy1�_8���f��Z
�"\ʢ�ٶ���e�{%R۩�E2�d�[V���؋5j�G�\��`�Y;�pǦR�+IߟQ(sBt�|2&	�*�a��7ZUd�X�.�;�	��nJ���'xξ�6��d��<9wUة�cm����e�z3�3#��3`�7��=���˘�F�6jm���dڢ5�Ik�@Ӻ�k32�t��n�lac�V��P���+c�T<� Ã�&ciX�Lj���+c �!�/�<���*��i��oxFDB�d�.��U��YB;82��ˇ��B�3+Rx��\F�>��sYyT���7�[ Tg&	$��P�tf�8!�Q�+5��̦v]lǔ�Z+�6�fvH�3��S6�1��
���YE4-�t��Z0)hp��npH���R�2��X�u������NPԯ&�&dVgf�͹�Gb]�pA�G��)�rn#Y�R�T/i�2q���]�w��;��x�U����_a�w��Y�����ܷ\��k-l�6e�	��cn]���\{�Kڂ,�tX4��@���zu��$P��S�j�{�e"vK�39����D�Ǌ,������"ɍc+N����C�l��3�2���S5c.�"ެ�L��>ʱ�IS�۰hvՌ\���`J��{�f��4P�2�Hʜ{���]�� ���|W	WI�J�S���J4�C��1z贲�H��E&��Ve[[wv=��Gv�^�Ȉq�zl� �C����Y��w����M+�v;h�	o<�/�Əlۻ9O9�ؐ${��2������*��3Iݨ�X�F��wF�x���ޣ;P*���ئu�z;��V�k�\�v�_d��^[��3�Mg���l)����	�K�ɀ��r-J�`/���ŋ(TL�Pf�;���8=�Q�u��j躦=憤ͼ�ف];�Ep�Z���)�3x���l��J5;��n%,uM�j^9FX�u����d�6��z��T�6[Q�(~�Łu�]�Z*5�`a�����(ܻX�n����Xۣ�
pÀ��b�J�y��#(&���ц��_5��5��n�6��Vh7��Yٓ�_n�<���5�4I�(t�l��\�mon��챼{����}[8��Y��ݮģ.�ɉ�x;�k�߰.�*'2� �U�T40���|����od�V.e����/&���|l��P�Xk�n��M�=�3���R���D4�R��Y������:eJ�݈�c)�l�Sa�rbY7Q�	;��'�.�@E��PHȲ����t����{��_�sK5X�Wz��w6���VY�I��pf,��D�Ca�{��Z}�i���2��	�]��W(��l���Q���
E���gK.�;b��X���*��M>�%g5�:�u6QI\ʉg��cS�Q��vF�!\a�5a�Ù/�gq�����
��0�]/`Ԉ,�̠jE�l�b+��7+�j�[����+��
U�(�6��خ�i{�<�R�ķ6�F.ٹw�/�P��o����'7�$)�j��ك�'6�B	�
,rW+z�D��V��Q�U�Y
7`C5OHt�2,t�v
��<�eCۜ�6s����K�k'ue��j�0⤢Ù&�.�d�M۽6��óJ��C����f��������k�8��2����i4��|�sw}�J�K)�`L���`�J�F������sYo�q��Is.e�v��=0�w�\y��meA��|ߕ�%x���z���w����$$ I4t�G;�j�S3!.+\)����1�S6ˢ3nã[Bl<C]��&,Z3�Fk.]
��l�ScS6�R�v�٠�r�ڢ<m,#f���nr��C��O-d�M\�3aî��e�7M���J�{Z�&4�� �����	��4��ZKUlIUt���L�5̽�ڡ�77j���f�����T�"�m�A\aL�(��4�i���ؙK9��R��hY�T�n52�`�L�a�Q�I�ٔ�uf�����r��ͤ���"D*�Y�[LَV_�K���.b�Z�P�\֭�f�F$�$c�ZX�JMÓ�р�-MF�h��d�1
���4�)�(M�հ�[.R9�QX���'��3*W,�4�p�B�P�kW��E�v�-�VX��s,��3�[(��n*��q���k��,&��(��Kk+`J���]WX::b�9�02�.�fnf��e�.*5�b��
̴���3*�l-��b�	1�.��ڤB��)i���2�f����)��nKġ�e�v@F�M-
Reڲj��6���S1u���@�b[����T�n4�m�Zb����H�r��&M�h�M�؄CZR�P��6\9nы%�R���0$�����ր6`�c6k�4E�ҰƎ�����, vζQ˚�[SL�*�)�&a +#(q�3R���S8�&Nn�e��]�Z.�"�M���v��k��WiB�T65�&�i�a�+��hd0Y��6��hS��)Y���-
sƊ\�aB�b���i�Td7�1���f�^Η0W] ���l�35c�F�b��%l�(@r�M] Z�T̥u���.�K6��R��t�n��,X,-t0�\7�U͒Ŕ�XZ�T�v)YL��\&��Pƹ]K@ɠ&��i��X�a���v�f-%k�e�V�$E+c��v.�`��XMd���v	x�,���x�P�+��pJ��s):�
������µ�Դ,��%�V�,h��T���Z[�����*�x�
�7z���	so0G�[p�u�-���I��r�f;CZk�)+�ːp4�SK�kB��mI6�H��g��-�;�`k<��|�<a�,�R	`����e�4��@ɠƻ��m!�e딀�3E�j�u�
%�F ��U�Z-����0��;��HB���3���l�SR]��2vʖ\�a�.B���Z�n�[Y��`��a�ˮ�$J.�2�ܮl,R[���n�nI�J���R�������Y�f�U�=eV	tH7M3"�ku�Lh���c�;Z����l
A��Y�X�-�B4�EH�$J��A�w!�5���	��B� BmHcF7L7JdҮ4�@�[�Yf4U���[AF��r�b��Y�dp8�����͢\���-KvY�F&���/j��Y`�1
`�,ؚF�[2�]��l]�٦��dE�UV%��ٰ� �p�� ���M1��Ʋ� �b7-״]m
�B���Ch]F4[w7b���]5$L��ijl4`-EKJ�Ի3j�E�df���ڒ�3)T�e,*G�^M��]H�Ж�;j	t��$���5�ۛ1-H���� l̤���:z���:��V�gX[���m�^ٕnΆ�#�M�)I�W[+���*��������2��%2�-�X����Z�\�6�LiY�8bZR����ҕ�4���lCf-1v�l��X��^-X�yһ����U2Cg!��K[BcV�&�V�<7��Tt6�s�D@�h�6:�U	��D���jA�a.��Q�k���m	kW[G+5�T&a0�(�����F=w0[�e�#�j�iu�1��i�M��D����鵁�v��i��%I�� �D� U�e�(^@��l�.5h�b�\U��ˬ�x
 �[*Bu��k�*;E��m��MK�سJ�6�L5f� �M ����#�V]-��Q�Jɡ�A@FMt]�(��!��n��ܫF=��[�»E������ƕ�� �9m9��ءvkr����7T�[,��
[`��4!kce���,�m���]f�1t��B�X��`�J� t�H�a��L��.뫱�%�&R���k,����"Ֆ\n��6ح!p��b��.��i�Zje��²�*ͮBa�M*�Fdװg 2�b�����<�x�)����q��:������tH���!v�m�;Q�靃��ˣ-m�*�Lg��ۅŶ@c3RiB�#l!I��K@�V��7T0p�@���M.�&
@/M��A�V]&�s�B�B)��r1�f$i���H��Rh�5W\`��r�-�+�P�TI��ٱ�K ��d-��Y��D�[��Yj�mi�6\հ�M5Ճ+x�ռj96�@��MI�5��xi%�뮕�D�%2��BX3;	�v�H�&�ؕ�V0h��{V��[`E��w4��j;e�孪�qrQ�� \)v�L�f�P��m��2�](԰֫,���465�C���,�K�GMp�����P�9�7X�"Q9�7�7WA�vb�ܻF�1�����ݵ�аFf��U΅�B� ѱ��d��#�(�X5���o�e����̵Wr��R�v�K �fƶk�:��Y�JQ��L���j��Q5����HB�A�6���I{m0�78��X[q�J�D���u��]@̰`Tl5l��!-�0r���5Ե3�ʀ���J��ŘZ��X�Chl����be��M����&y��!��n08���`#��J�6�v&��R1��u�!Ļ7E[k�XҒ��*Gg��)ذ��&�M�f�M��X��v v&��Y,%�n44X�]Qšh�!skbå��\���=jLL��Rc8�ֻ ��A4ٛ���m[��Z�Y�Ti1��v!��\��l&�i	����bRX-��9�F�,��R��CZ�rE��U�k1���5t!�@��ݘ$+n�6@n�÷%�v�8[�XJ�����JU�Y��]�li^y�]���ɊLb�t�L�u�,��ԕ�b5�s�������rŽYc-��)-�2�؍,��l�QeJ2锨3�1�c&�E�R&��Ҹ���\�8ͬ.�3CKx�����i-WAkn0f���
�WAlŵ�l�H4��u���KJځ]Ђm���Xݣ���cR9���6�fi�Jn�pgNmkG�rlG��	nŗ�+@!���EY�5�ڋ��;�I�mX��5F]q^u�@-]�me6�X�!�.�kl�[hF��b��.�rL�
X�˳u�@�5"f��d�(��B�T��!6U#p�+q�uIV4�������pm�(Z�Cl��6�%��Gz,O h\n�l �q��b�$�=v�6��0s@�]K��W&���F��j�jBf�8��4�+�L�W	.�-N4�כ���Ʋ��]�2,sqDK�m���]EM��kEU�b�c����u��1Fk���*��u�@Ȁ���ذ@"Kum\kpQ��θL�BF�A�B��su%L�Ie�Қ$J�۫���[��ɡ��!�K
v1��mCM`.��T"�WV�ʗR�iY��@����������t;�wl\Ў�Ō�-U��Zzw�|�K�r�X��4�3Ut�\�@��ط20/Q�Ђ���U4tԡ�����-u��(�ԙ���k���-�DH��J$��h�WM,Le�:�q��R�*�d�1�hV+��6%��f�y�#�A�-����`{:�R��ܥ�m҆K-֩A�E�Sݜ���٦nL��+qb�%%H�[.�.S]	Zb:!�-m�rݬ��琎��õ���:��n�;��k��&kY��YZ��q(̈��RR#�e��̕nu- 6�^R$.v��%�ص,-�h�4#f��6�N`�i�bݒ0�e�+�Q�*�d�Ьls,lG8�6`L��Ԅѻb�6ʰ�F��Z5�ڍ��B7A`��uA\\*�v�Ff�2�9��W���LKH��Yk64i-�t�U��d,�lm�����M�7�c��6*F����4f2$-Tz�1є��BdKP:�CG^��eY�]��\cQ�;3b�h� ,+Kc��h�49���u	���-R��5*�V���V�X��s���ZB$6���3;<]0@i6Ël��<�@�Y�6�&�Z��r��d�3
#́5zݻ2��X3iB�� ˻X%�8]�"2��'�Kn�kp!h�K e1����Rdl1�ι�]m-��%X6Tm�Y��]eҦڴ�A�Л4����[+��b��Q�n�<��A�@��DyTܙ���g�jT҃veF��d��a�u4p���qQDK�)
��ۢ��d�f�S���5F`��SM�--�4�Z9hCSV�5#X��̗M��e���+&֦��j�=a)WRڃͱ�f�R���n<B��X����բ������U6H;6[e��U��f�N�a�p2ѷZIa��`Čq�]5;F1��-P�El�u�X�b�B�Ykl[����.���b٦+.�+.ՙ�%ٳ4�-�fE�Ų��h�鄨IN@�h��-J��;�B�6��Y����[�fl40�A�#��n[[�@ؔЀ�ӎ��d��qm*]��b6��6cfaƆv�spJ
"̚[�a۪�mN5�d�c.kc�R���.*۱M4\$�Ѵe��Ҹ-b��dfÉ���+�Vkz�!kH,l��if�f����`��-�Td�4�[)3"��Xt��e�:.�4�X�ա�SKYZ<[�]H��4�%�n{�K��cj�[��$�u�+�\��u�M }:�ȶB�g��i[pIMnH]�`��r����u��5���)qwRͫ�.����(��ڦp2��X2٦���W-ٍ�faF:5��/��0J�ueF*.�kUˮK�(�\����*J�͖O��	��7 �TD�DDb�ۤHX��h�r�h����䟹�iE��;��+��$Q=��a1ϗ� TA�	�+Α���Ʌ2"|��EynX��H�`�»�s�Q,h2!HL��Re,RA4�n\������+�5�[�(�M	F�w+�N��7]��4QIH�r�˖��D�$ш�!���@��@)	$����1�H��]�&�LiM���Ɗ(�;���6�A�(���1�3(�%^�Q9\�t�
�@
"M|��N�4_v∓&De�&�(��h�+�� #A 4ɤ�";�B�c�eb	d�1��(9��j�ߋ���>A1�<&x,��\gX`h[��/9�֑B�$�mT�tt��T�k�`F	�-��+�]4��g�6i�/��]�^Ǆ����Y�]��D���e�a	�A��ua���v!���C1R���Q�P���7RY���$�f.,���](%h��fu��9)ƒ���3�ZB!]���T.�
udn����W(�ٚ�&�ˉKYKL�����Ё]#X�B�n�d�7�k*c�,����6��M6 aK��X�i��fQ�"�Q�� �M�l˥�� !�c4���fV�@�2�0:�3����2m1��-Ļ+�ڌl]�M����\�@s�	��ݙ���5�כ3j�2�=�JM&HY�`�GV�b�m͔�t�hJ�@d�є�����hK͔*L�%�#f�hn�RPn���ꡫpZӦ� �:��f�:XR�xG3դ&��uz�*�i�M�L�fڹcK�P"�5�m��<��*k5T�c��+���R��l*��F�1v����˞X�K5G6n�P�K��Ia�cCWDs��.�@v�fd-cFͥ�#IX�ر��G8F�!@�v�e��ҳ&U��ܥ����ʷ@砘,���*s��St�1�h�%pa�m�.�]2�G�(mX��:۠��Nf]���4�e��[E��R��3�֐����� �YJ�%m4]H�a1V� mSW9KX��M����i.���eP�e0�CkkDְ�M�E�$�hh�$�"Sv�F�ued��.�0W.�qR<d��Y��6���ja�T)h�LРh"U�f�!� ̳gX,c��k��i�����2����c�W&����3��-���#y��X͑-����ف�Is�$�Y�+0�$M����^X�˙x8a�
�1���$
�	�����V�v�25�9b�m�0�Ԋj�l��b�d��(��gI$k�M1�-��6�9h1�������`�DP�Z�
��KIIaac�VRڐc*m�$+֑���,-
aya+V"� ���� �j��У �6�5+o,*l�b�z�X�Zm��e�cVRQZ ���F�K��� 6��V�`�`	
V�D�m������]��* ��e�G6�pc�[sM�Ev�L���+�ͪeDȑ0����-ڐ!��d���S��Xd"�͉� �bT-F8�Q�C�"A�[^�A�D(������!�H�����b�m�rC�*|�) ��[�ͱ2d�͖��PFܯWX@���6כ� ����ó=�j�[���ٰfzA�˄AƼw>n-�^�EڇN&o-Lm�)�@�-�>��̍���9�3��
�qu@��*/'�,����Ȇ�[��myۤFߖ�ZB�w�}"�Hy�@gqH ��"� �-�:�ā���T� �9�n[�-�m&dL�	�9�C]��MQ� �,�k�z^�"vȐ[���^Cb���vK�,@��g�FbDW2�Qذ"�x^��p-�@Am�"�r0���d�.�j�P�)���F�0P��iA�ѫr�纏*}������ӟs�ŵ��uw���{-+�2��5i���7�g]-G� ��SW�36a验�3��
�w�TysvD�������{+�7�A�y��s>n��:��V)��\��iP8L�/K�n��j@!�ڽ��=u����n8��D��x���ث��+F�,@��OH��+$=u��ﲅ9ٟ
޺���-�$���S=q[�RQoZ��v�幇ƍd��'t*� NTy�P��Ck��������rf�١V:�Cuf������֧[���"D�k�CcQM��&�Z$�@�3������`_Nی��7�T#4��"o�\�7h#� ��Ԑ�@��sFN3�m�ɽ�
�%������WW�V������OH ���k��6��2Nday4ϠK^��@�^��� /�=��^��^�lN�P�j*���3LU$��NЯ@��Eԗ"��O+�۴�SN��v�A&�M$�ʚ˃(B��mܭ��s`�.:����<���ʾ��V���b'34j=�Z'{r��\ȩʎ�h�D]]F�;�������^�k9[\n4�&w�v��&��g,���3��󗛿 |q�Cm	-�).��=	�j�������8/���{6�H'.���s���~}l�����)<����;@�ff�s�1�E��iv),rl@`+*:[T�6�������?}����-�@�mU�\^�f�yryn��C)U�U捡[���uǓk�ۑ ��Q�6���<\��,=���#��7PQJ�N��[|nzT�) �A�FL��7c
mI��Ǩ�r$���׋�TkH�����Ee�l�3<$r�q������n@[�h�v�r�U)X^@^;� �ڑV��F��fT��-��r����:�F�73�@��E�Y׶���n��Ŷsa��=��~�+e�%�Ƭ�VWN�~��$K�`M��۔��cU6t��)�b�v
�$8�c�t"5�mȐKp�ͯ Cn�2���X��섂�J�R��U��* �gqO�>|��n͵��js&��Z]pJ�F�4U%E6�mK)j�2��HgeR\�T��T�F	�6:�����������Ʀo�����Ɂ�4�O�ɓ5���[�b���FZ�y�>-��n[j|F���ž���X3p �ڧ�j�jzFeH���P8�G�����.���ǒ����}����m�����x��܉=3M��;D!��@�Aw�ϐ^-�DmO�m&-��B:cv=~ �܉:�@my����"j���6h�9p��lZ�T6�֬�232D��k���|�S��7�î��^H��F�)z�qF��fT��-��{*<�"A�^mz0�5�-����hGI��e��p����n���w���-冥�u,lKg����G�t4����.R��7�w��o�޾�{����)IS4�ÉIL�+5̵-�ۡ ⛭�`�qX�vtˊ�X��4�%�%�pU-'����Č;a�e�SLBa���^nilˈ�bы�j�ËTvV-V����󢹥ٲ���h0P:�g�ܲia\�ZDv,V㔦�J�8au���d)��ɦ&p���b�+�2�,,�1�3�ji����/l(z�O�����KR�K+�6%���崊�a-���Z�5���?��_��ּ�m����UsEN눽3�CkJ��^C{sur�Ś�]��ڐCiq�}U�bsf�mX����z�n��؉���&l�3<'Ր�AƼ��/5S�H�����p(�m���Yn �ڮS��#��3�:���3��F�� |r��FnȒ� A�kȆ���ʮ1:���'�:� �������+kZ�َ��*L�RĈ1s6�僷Q>��,޵>!�Ÿ�C�7N��1*Ɗ��[=]{&h־�ؘ��A�����6���B�x����=z�}_���61-��X��t�v�J�B(�� �usP�܌n��?Y?�z�>~�� �55jw4Ɯ�*;Ѻ)r���n��C��f]�{H��'�\yח��A�@�ȍ�:b��X͚�U����D�p*���䮡�0�}k�78�ʜl]l�W��ub�K�u���tmI�fz���|�ӵ�'N��ok�E�L��h!sSFz�������Ҡq�;RA�/�r�|i�|���q�-�q���@��͜�]0�r*��1gg���F8������F��{;9{�Qk�r�� w` �j}Ws��s��F��@���I��C ;��AmyۙŸ@���!�������°s��؂���uX�/�8"v��Ay�#� � "�U�&�j�믵2d0�3�K���v\ۍِ�T�1"jڋ,�jaf�ڙ��e�uZ���f����A��uِ�!5���;8
�5�.&LFlz�W��߽>>mp���@ww�o�U�n۱�<�/|w���ơ�9�Tw�tR��9Q��-�1�ՑVS��#b�/�Bθ�myx��ψmIf���L����\.�ql��
KY�-\{]I�W=�uӴ;q�F��:�׶�ܴ__Y5�n�B��ۊ��������v�^�hD�iP;�9�@#�<�
��כ��&&��D3[�Q� ��^�!����:�9U���:�3= �k!x���+����������Am�� ��@� ��E�Y�m0�=�ƚ�s��F��ʏ"=� ��'ϛ������C��3OͮoQR�]�T�*�U%bG[a�@�P�\F�pm�٘�>z~��� ���CngŴ74g�Z��<;ZT �:�]�<���A�mI�/7w"����X���>^Cf��$L�oA�:�3= �N=��[���.'c}>��`��)cA�"-�[ֺbr�*Djw��/��F��	ʏ"=� ��ב�1eurSʯJZka�^����h�m��'�@;ZT<ԑW�;:R�N�+W��V�j|h>�F��dӱ2��4～�z �#�{N	H�Q�{8��Y�32�jٖ�}΂�������y�|Ch	n<��"Kq��� ����MՇ��Q��0�T��� Flyr'�͡���{�����y�Jۖ�9�2V���	[��j]��H����,�G!��0TK�X�:�|���_���	m����I�.0�"#tEr��7��TQ����'���۹�p���^�^J�ȋ�^́b*�v�Kg8�i� q�jH}�y�
�T���#���Z���� ��In ��V��&��B��t/���}�`�^ʎ ���Cmz|��qS�����z�����Ÿ�mH�����Ɨo��"�{*<����]�4�M�P;��Dk� Cnd�y6���5���c���o�D�EUR:�BW�bm��3�I� [���mlt��0*ʔGՠ7S%��{\��αC�����OG
UV�ƣ�N�=�n-hS)�W�3j-Nr�Sr��e%l�T���>z��Ֆ놴�Yq�@Ù�q	j�Ie]��Ĭ�k��\��Wa����.XW��lWV��!.̮�[������Ɔ�@,ëV�t����V.��9��A��lhA����cD���t��j�4��qUGVVmB�Q��`͸.�����%*�p���rW�lʉt`^3P�ל]f�n+4ֹ�2ʛ*;F�\��n�\3O>_�X#l-�b�۶nPt�R�\�(��v�r��#j5\Pc�}�g�<�{q	���0�[^@uUpm��{�qV
��J���5�kѷ3J:^@�͐'�͠�p/�T�DA=����>=����C���Q�
�r����dIn8�=5JVGV�r�XW������@����^�Њ�i�
eΛ��v�!+�16�P8|g9I�/�  �Ԑ�A@�U��Q� ��r$�Ǔk�v���T]�A�5X3= �p��%\#��y�H�����Ÿ6Ԑ[A�g{]�8�o�Hm]�ПⳔB;�W���^��q��׹�f�����j�\2`�!�	��̈́��@���v��^��kp)���Gd��ٖ�r�?s$NgG����|Ch!uH�`��`��Q�����p,I�/  ^�^ �ڐCpn<�16.Z��#���7�[���S/4O�X�W���#yv-�:��I��zsf4֓Y��iܦ!BAS����`�'�ͯ̀FtyJ���rU��I�5XQ<��@�5��qS&"�ٛʥ�r�6�"	�jA͠�n ���#�z7����1���f��s��]�r<�:�D��� CndB��J��$����^�s�AE�R��NM�6ڈA=\�5
R�sdւދ�<1�Ch An<�6��ĴƆ�N�lR��'\3����zNH�AD�eG}�y۟O�hSrjc��<5��
&T�*D�����c�!b�ͼ�[���
�q���ڂG.�q�j|Glp-�>�Uod��;\��;�W!3ѳ�5P�:9����t"mys�� EV��t51�:cֵ|�G2��ƃy��{bM�6ڈ�W)!�p+U���c|u)#�;��Cm	�D7�>�G��'�S͋h�tkeg޳�/�'y����1Ds��=�b�`��݀��P��	(�\ES[�Ta'��0A��%�aM�w�4�:���J��kKNށ�J�P�嗈�ס�*�>��̓N�ֻ;�A7Gff:?�;����ݜ\v���������Z�i��M���CwS�Cr�D�nB5��Ր
w��u�*��e�v��n\�u��;�|{;,h0]C
Ts��aO����멕�K�YYΤF���t�++��s�IaT7/{U9�l'�+}�i�*�*�8���0^'FuӺ&���G[��o*�f�X�{�D�ܼ3;59r2��m���6贓D(��r�[�3zU��9�+�<�ˆj�7�����_�R��6SڻN�����Hq:��ĀU�\E�,����)�˅�4A�g�}6�:'��a�i�pM�K��{6z�W[�b��`�Dѣ]�f��h��D�
k]�X��Ǣ�DK�2����&�t�t�WE�W*3�9���WV���xP�lcˋ�]�l�q%��XH����L�����c�<fl�s2�0v��~V��E� �[����uɜ�fj��b����o�p-�Ifs��۔�i��[	���79v���f�>�h�0�Eɪۖ� ��,M��\�}��"�Õ��-IQ��/9vQλ'-u`�M"�I�ׄ<vJ�,]9��+���6rg��5R(��r2��몌��Krݖ�n�3r�n�a٘�7ͼ�m��tV�i ��/�\L$�̓?[�m)3"h�	6"�0��(��B&+�ܣ��!�6%+���|�i��d21)1�$͌Ah�IR��	4TQ4|�a�Q�EI�Tb4b�cH�I�h6湓�ۘ��+р�1�1R��E$c)"���L`��I
Bkݺ���v�[�(�r�CA��1��)$cDAQ��d�7�ך��$��!%%i1X,��ѴF�%��5�F"�J3
���H�����7�Ԗ�rB���dm$BLR�0�H$��$�A>ܛ��䘻{S#U����:ב���"��۸����<����jŸAm����2��ms��
���<���&*�9kv��/#���m̂p�-�/}�+`1��#n�gV����0cm��&{����>-��li��2�A�rc�&ī��@�:J��ь��،�Қ8Q�mtk)O��@����7dO�p� �ה���{�0��fxz}HTutȾ�������!��p� �׎M�1���D��Od��)j��"wC�\�ĝ��=��|�H�q9p�zֱs�GnȐ|t"�k�۟O��h`�z��}s{3<�"m��w�>;\����"� �[jG�my
�b������Eǳ�}"A}[^U�]Ĵ�+ު��U	�� �i�"��z'��Dk��]��`��[���Ȩ�D�=�h���a��M�yw�p�oOvT��*d
r�Vb����x���ח�V׳`Yn<k���p+۴��ܠ�j��D��G$�L��r���3PG2 �1z7�Egb�yUr}�aAХ����L��Q��V���X�i��X�����r��dŇk$o�G5�CngŴ"U��4g'_D@��Q�8"۷�.syYu�  [jHm �xh��'Y����bA��r��%�.�z�T�	�B ���Co�UԎ��*=b�dA�R-�7��j�&w��}����2�����yq�-��ǐ!� H�Qȋ��G� ����[h/B��[����naP8�gyI���o;g���ha��� �r�A[�"��"An*l��I�ر`*^O����ީ��g��\"�W�n����;�f�,�\2�M�Vk�i,R3���*^noa�i�g�P]��lM��R���5��:m���#��<��8K�ѳU����OG���{G�XuN��-[v�@�g�H5N���]"<̛W���V����I�Wcr�Gb���KsK����A	RW6ŵ	HM����Z1���,١�ĭ�L��[
��7C���q�-�fRl�X�����c\WC`ڕ�b�e�$]u
,�
]�-`�*7�a���+��69�k��m&(fif��ю����3f0bXi��K��Y�nE�1\֔,��P+�e+�+0�E���� ���)�5.}�K/_>~u�����+��Sws}�:eJh��PJ�]c�q9�Ev� �B ��ב�	n"enqz�z�"��&�O�悅WW�QS��Dܲ�q�W)!�p!�1D�C�����uǐ܉-���j�!�m�͖
�kuRA�2�H>9p�5x6�|[A [���gk��L��ٰ(@-�v�vƩc��K�;X@��<��^y�8MP�{CZ�m܃��y6��m�o���x���x�B�����*��S���p�W��'�q��D�L7" LL�fR�b�q��c��YTĸbɵɤ,����ю�]^��$�k�OOh�M٥�� �H�Hho.�as��Ӹ��^Df�����E����k� gW�cK�!�P��Us�/p�̤�`�תq��Z�;	�)���Nw"G��+�Z�z�G��+Wf������=�xb���t�=�+���5:?mFK��X"��Q�v�-�to��W�Ů^DN�'�:�n<w��ml�sbp^�Gk.��,�;��ܢ�q�Z�A���  [j|Ck�S�hd�7p��ǯ��u�$��-�*ޭ��2����+�k!x�veZ�'�T�z��"}��Am� ��E��y�<r>I�z���<z�{��}c�J��@�q��dH-�������잂yhy��lK(�������%�6��wR"�.�$�*R��m`�@.��k^^!�"|F4�SW�
k=��ܢ�qIp�bq�NCI���z ��RCi�[� ���V3�mL��0��kӽ�b-唷���
WxO���^@����&�NP�~�d���x�{�I6��
�LI�=0�2�m+��*�;Qb ���D��|��QU�/���9�[���ͻF�t6m�q�zΠ6D�B�oO����,�a��i��꯾��'Y�]שU�Gf�E|��y�P��"kȇ��Ч���;[Q@�q�Fv�713A�1�㴓tT�\�T2��d�~;���jA�%��M�[�T���O/ �0\��.�I�B"W���9�Ȇ�ψm�.;�}؞�9�M��]	B�V9�9�h˅iU��4�6�m��.5�����>�|�!'� [��'R.�kN��ӊ�5lM؊�
��:99;��A6D��A��m�%�^#����Gl
~���>!�sV��Mv�cr����{T�Ǜ�G�����=w�������A��AHQU�]��`RAJ���6�Y�Ja�P�5RA`f]��WU�g�p�?L���[
7RKN��<	���6�Y)�ü�Z����H)���D��2�i5)��v�L��P߾<�M����)7����NoV��JH,3*�RhB��v�i��P))32���+/*��.�LeZձ7��O���$xR;v�L
H)\��+�7Z׼���J��F�}`�mB���J�ܐhfS��MҜ�Ӹ�V3j�����Tk�<y*B�n�S��=Zr�t�v��Wh��  ^����2S*�R
a���H,4
fe���AH,3*��) �(�֔���I32����9�*����^�s�
x$��<	����*s�$� [��g�%$(Ro�4��RAaF{p�AI�
`f]��e$	��@	>������5R�>��A$b}m�%6%�R�p�i)�*jh*U�[+�Q��꭫��]�� �ߴ�
B��}˵ ���;��i����2�hi%$*0�թ���ޜ�����������AJ�X|��%g{����o����P�JH,
�洤�I>���
Av�eCI5)��v�Q��
Rfe��6$���~7��_?y�w���'�S�Ԃ�R
{�X`p�߇޾���7yYZ��H,/��� �*U@�ݩ�����w>�H,��L3*���;��s�7����H,
�ڐXx
s��lCi��L3څ�i) �(�֔��R
gr��肐ZC2�����}�����{��x��ߏ;��������0*��|�I
Ro�XH)�{P����
`f]��e$
�3,07��:H)=��p���]� ����@m ���hr$��@��(��O�s���M9?_�%��,�R�Vm �S)�yP�D����};����7]Rq������� ��}�i ��03.Ԃ�P�JL̰4��RAa�P���B�̻Y<�眿��{͏�>� H D�� I�ݕ��߾�)8��>�Aa^P|:H)���R���������̓%0̨Z�) �3.Ԃ×|�}�����n{7n�PS���d�{:��=�^;����?�'�딯L����!��M���Lgp_k��b�J}�����$|�Os�`�1լ�5�DN��,���KW��a�V�cfGQ��j-���]Z/q 1��M�.�	lYv�j`/WXWfi������][�a�.�����s؁���\�8�T��\6Y�i�,Ӷm)�D��a+�6�WlRFf��l�t�).��IaB[\��rT%)��6X��	���p;e��̠c���nf�����^�h�!+�������[LKr�V�F����acͫ	�$	kln�%��M3͍���N�>�zH��wc)�ݨZ�������)���
fe��� �3*H)���9ϱ�Mwu\�>�]�ϙ) �ßk>��מ^k_k�Z_9`iĔ�XW�p�AI�)��]��e$
JL̰4���Aa�A��AHT*�f]���
xs��|��2�S΁�Ag�%0�T- �eڐXy����ekw��|�^e��� �^�>�m ��B�5����)������`k�{�:V���3�
A~�sʆ�
h@�>�R
ACQ%'��`i�) �̨ZAI�B��k&�RA@����Lw�|~�՟G�$���2��Ue'���<	���|:H)
����R�$���H,�d��H)��v���S3,2!�����ҭ��jw\����h�I�P�kJA`j4�S3,�)�ʆ�
h�oÜ��zk������0*��|�I
Ro�XCi) �ٮsw����k!�'�
`y˵�C) �P�����
Aa�A�I!R�eڐ]0) �ff��Af�)�eB�r����_=&�\�Rfg�yϫ{�>����.���*�a�!���C)�yP�	I�߮Ԃ��I32��肐ZC2����_�w��_I�,pG�Ĕ IDL)���,1mf�&�tZ,6E��e��ue�&�Q�In�H)$���l!�$��þ�- �Ѕ03.�M) �#�A��|̬q��ѵ	�ܛ���yP������k_7�6��N{�o��<�ڐ]F$���i�d�ʅ��%$)�f�H) �s,$��2�h����ANG�s�fd�l�ث�51Z�bqa	C���ke��݂�0!�F�ҳq�����{�i�u�H�Sb�u��pO����X��m=���=��@�<׿�A`~$�>�7� ���ꆒ
j��ǝ��]��U���<`Uݬ�2RAB�RwϬ!�%$�$��̻Y3�~���ҷ�M�
JMk�L��X{�GI!ET˵ ������6�Y�d��C@��
0�թ�{�k�s���V�y�UN�*�_xY��� RAd��a�j�������kJA`hi �fX�RB�$�03.�i��
����=�2���i���4��JH,+�p�AI�)��n�M2�
	I����5�q����U��>� ���>��
B��gnԂ�`RAJ/�w<�u�5����)���- �4��թ��RAL̰�H,�2�fT-II�Y�ҐXH)��0㕙������R�/U$�+~mϱ��]��W/π�Wv��d���	);����JH,(�ۆ�
M!L˵ �%&fX`_�b�]:��c���12AJ�!A	�]��q�ه,wPFmmw�`��h�B1�����z� �*U@�� �`RAN���62Sʅ����P��f�H,4}ߜ�M����Y���$�Շ�m �}W����kۿ��a�P���X�����I9߬��
Aiʆ�
A`f]� ����3,!�%$׵�x|}��y�!i&�)��.Ԃ�P5��@	>�e��O�~�:��ɿ��|-@>$�U@�nԂ�I(>�i�d��C��w߫/������>�V��) �s�Ci��)��T-BRA`PfkJA`hi �fX7D�ІeCH�$@�W�l�{V��H&����TW�`�)�+�/p��'n;�O�8(�T�U�HPC�d��N��i��g�L�i���h��R�<�ư��0���� Q�_ic����5_�π�v��d���$��XCi) ���ۆ�
MS2�H)II���H,3*�Rkg�{�k��s^���R�$�4�Y���{�B��$���0�թ�}|�:åZ:�*6uG�G�!)@}��
Aa�T-II�_y�w�e=�2�O1H,H)�2��AH.�;�$��̻Y�%$���`i���¦e�I&��e���O;n�����^䤂��RkY`i�P�����N䳹u���O�L�2D���nԂ�`RAO�큤�ͲSʅ��%$eڐX{\�w�}�yΕ���S�j��Li.��C���B��34Բ�a�U%Mj�h.�M%������ό��6�Y)��9P�%$�v���S3,$��ʆ�
'�.���&]|����	"}����P��o߾��ϵ��9�XC�II��ᤂ�X�����H(�3,064�XfPht�RU@̻R
AH)�����5���_f��<H)�<�ZAH(c
̻H,4����h�����xY����i��S2�i �4w��A`hi �fX�y:��^��o\�[C��i ��)��j١��
AOs�Hm%$�H)4�03*�42�
%&fX`V��{�缲�����c�-�6w�˯��|*`�I!ET�� �`RAO�큤�ͲSʅ����P��2��XhaI32��Ad鯾����O9<a����) �(���A`i���g��� �!�P�AM������w�D���<`Uճ�JH(P���}`i ����N�}��yG]��u��u̠�ްu
�B�2����
܏l�<�M�Qr�ʵt�Y�Fó����̝�7�u�$�Fi���x�B+_C䂓�
`y�[&�) ����L�$�$�J��i������`i �l��2�hj��>������WI������3��;�����n���.�a�H,�L<ʅ����~�$��S3,�
Aiʆ��$8ߒ�I�+c�p>��b)"�hR��t�I��GD�c,ɘ�U�݅���.�a�v��`y�l�2RAH)�y`i����>�ZAI�
`fU�j2�
��7u $�
�x����-;�_JAa�P|� �2�}�o=��j��n��n� �
H)^{���Af�%0̨ZII
���AH)32À��%2�fT-Q) �|�z����IΒ<	�`�G=@H)؇�T4�SA��v��}�tL�>�][>���R
wϬ$��~�p�AH,ʶL��k���;4�P=�����m$��C������ZAt0) ���6�Rʅ��%$eZA>~w�?df|~��ft]*��A[;Q���.�a�H,�L<ʅ����w��A`hi �fX��
Aiʆ�
h@�e[4��P��޵�ϵ�xO;���0II�sۆ�
MS>�H)Q)32��|���O�R��3�o�$j��� �*�{V�]
H)\θy�~�y�x�R�P�=II
}�i ����`i �pe0̨ZAH,�ZA`x�AL̰>���;�㾐R�7���
k���+�=�w߼�F_��FJH(TII�>�4��%${��I �3*�<����BRfe���ctex.3��?�U|��Ö-
�Z��ƙ�Iqj䭔$��eNԄ��w��CT�L�	�H�mC�[�,���ŷ�6��QD�Y�%����p~���srfn�s����hUp����s������0I�Cՠ�ev��ˬ��[�#�]|6nd)JB�ڹ��O�ޮ�V�F7wWw:�ļ�ˮ�}��݆���(��X3�\�avIZ�L��iu-+/n��l��ZG�q�Ah;���3 X�B:��E�F�
e�D86ԨsTs�w:�M����9�ٓf���r@u��J���Vj���hIݍ2�Y{�e��/��H�^��n�ww�v�r*h[���!Dt���.t�k��[>�w�Z�a�Zv0�ՑcO���r���	A�˳+(d>��wy��Y]3���V�5��T��K<a"EE�g��Tj^�w�ś3&�����+Ό��ƫ���6M�K�vT�;O�S;���Q�rL��v4���=��q�CNY�p����ʊ���`}��M�N��o�ɶZ`��w�=�Ւ2�.֦�ef�oib;mFŵZZ�jg��x��2�r��P�wT�y>U���N�l��Οfv�,ܬ�k*ٌ��۔KMa�M��;�v�䌂n�KfX)���2$���4��u+�؃D*��܍�N=W}ռd�ˈ��_+���k4��6^�{b�0d�w����}*i�n�[}�,<���ާF�}���ˊ]i�h�q^V&�i�G�d�r�e��]�H�-�����t_.��OsE�,�E�d�"����ٖL�P�J���ؠ@�E���fW.��p�d"ɢJ(�)(��RD��FE�4Io5�h�cg��Q�w�E����Eh4�H��50�J#bM�eF��L�đ��G.C���6�@�"l����S,lj"",��b�Ƣ5�E&�������5��,lF4`�(Ė)5��lj�`��n�F�F$�Ą� 8:���|�ԷZ�3����.�eɌ�)^��!`�*�˭����2]�4&���M1v����Y�L�m�6�hZ��&�kM��V˫DtwX\�5`�i]bBVXB�ͅ����1�fb�Jr��:�+i�aJ���fiLh��+sk�ݵ�ܲ���]
�h�ވ�,W��3�m!�5�D4���`3U��,�Y�`�b�6��`�kIQ��f�KK�,���������uSV\b��k%�F���ZJ�r0f�0Aݶ���S�1�v�[�J��,K.�i�Ѹ�t�42.
:n%ዲ������
�t#E����&�ԙ�a»&�j6Vm[���3f�`��]2�p��̵(0��
9�[6��X`��hm��Kz-&5)�1YQ� v�]�%!�GR�`bz�۵.٤�)�r����a)JM������Nlҵ`�h�[UC&&���Rˊ8���.��\UՎ��D�e�鳦4�m�E�v.��P�RjQCBP0�+!ucW�Z�a�P!,.�����`�-M�[SM�!�Ѱ��V���@�C�TJh���5�6P�a-�A.-N�Լ�qk�նd-L,*ۥYj�ְ�c$f��a�jP�GX�p�hS8�(bF� j�a&��DЅ6�M�tl���q��i��iSZ���� �T[u�p��GC8�l��y�c�4�v����
%׆e�Q����-Fh�F�M�V].�FQy3,j�.cZ11�۴Ĥ�FY�R �1���Xa��\]V,��xq6*muv3F��8x��.�l�+�޴��]�WY��%�&��eF	�lccYLSKl+��]���cEv�S���*��<�M�笻pB��
�t[���\@�(2�b,�-�Tu��AQ�����(�{[mm����f�teʪ&%�b���4�͡�,&��v�6H�U���͘��1n�t�M619@me��Fƚ�W:#��ݕ`��R�c�ٜ;2�m�[2F����k��X���'t��'�x'���)u�3�����^��2����K-:mUk�� �M�\�uW]���nC��:a��.�d�fIF�km�9�\HՆ� Ha�m(�K[U��9�T��P��+���֣M"KG�.�Q�a����n���a�l�ۨ���b��h�d����h����m�4d���A%�ŸVTf��\G4���	XϿ�?�[����-#���(YT�6��J�B�@�.r9��v]��Wz���þP~Β
A`y�ZAt
H)Fg�i�)�eB��II��V�Xy�~���}7���k5^�i.�a���&�|��ek~W'Xn��R;�����i �w,$��ʆ�
A`w*��%$)%&fXCbJH,/�w��3���~k�z�Ri
`}�l�I����`s������g���i��A�� �{V�]0) �����Af�Ja�P�/��/��^���Ĵ���ui���$��l6m �Te0�ꅠhJH,
̽$�I32��AH.�̨h�D�|�E�Rwe�_�}n	� ,�*����I
RwϬ$��=�ZAIȅ03*�5I �fX`m���2�N�
C���k�Z~��̫H) ���}�6�Y���{�B�В�
�2��Xk|���޷�����^W��AMkVm �P�a��Z����]~���<׶_q �<i �{�I �C=�i ��)��V�2RAB�Rw�`i���³.H)5�e['�<�~w�7�=�Ԃ�R����3����_}����f����ä����{V�]
H)Yߴ�6�L3*����2� �ߎ}�"�>|���~�.�.������5[%�6"� ���v���պ;!��H���=�O��'�D6�Y)����-Q) �+�ޒ
AH)���
Ax�eCI�om�O�pN��g�B�}������w]�{x��	��ݰ4�D��XQ�p�AI��0;�[&�RAH)����$�H)B�eZAH)=��8{�3���w�j��u4�m_n��� b#w{�\�l�r�`Lڻ�Ȧ�a(;�=���a�E�W{�W��j��7��B<�? �Ag��L;�B��II�ﴈ�'����sU:=�%��Dx!J�m �S)�r�i �;�ZA`x�AL̰<浖�y�}0��Z�w�$ЁL�d���S��`iĔ�XVe�I �3*�<����II���������>���g<���H,/�����X�ZAt����9�h���2�hpII��V�XhaI32�hm �}Y�����~��ٌ9�H)���/I ��r��肏|7c��H�x�b�E��8'T��
��|�I
Ro�4��RAaÅ�9�wW��k��߰�AI����l�e$
JO{큦�H,3*�R2� �F$�����͌��2�hW9[O��;��xKH(X�~֒���}����߾���e}��Ձ����e0�T-II�G}�$��S3,n�)�C2������o���<��˯H��YK�F�b;RP�W��Lt.v��M�M��IV]:�0>�[;) �I)<�,!���XW~�i ���e[&�I����L�s�������_u3���������$������[�{�2;V�^0) ��큤���Ja�P���P��2��XhaI32�q�J���@� �|���틀�zG��|��) �y���tAH-D3*H(��x�����DꟀ|(Dx<	�����q���L��9�s�y�����5p� ��� ����A��ui	��B0�h۸h��O�@��˱{�R���w������<č���#,\ẳ�y�֗"� �ݢ��sMՍ0�,n�~�4˪���  ��Ψ������� ��	���T%��w�[	���&��jl���������n�� ���u�;ڄ-����b�n�<��z{_z/u�Sy����ф�<�2s���b����̏fG�2g ���{����_<<��|�(:�Yʧ�}$�JK�KU����ǔp��,�+��,ҋ�`�\2�]�%�!HfkJ���C���	!u-�b�3 O]�+�6�`rZ�`A�ؤ�,=9>}۪�I2I~��>�>}y7k��_��|�U;ӱ�	s̻�Tc���
�C0i�q��ooyLּ�ffP��Vnh����ï5<PuH<��͌�$��^���u,YFW��Hj�5��
���=�j[c���Y�vy�$��T�t+W[z��f�����V�n�����CӇ��{���Z�.�xS܊�8���0܇zP{�� ����o��Ƥ?I.�?I�I�i������T��/��̻�U�eG�^�W��ZǞx��'���l�Ckoh)a6,
SE�е�5�Eа,ffX�^P�dvt�j�L����-2��Ӥ��(�%����Oۧ�H��?!���ɞs$~�5|�K�L����؃�.1���{
#Is�y�t{ӤR�{`��2�Ss1<�B=8
����'�D~���CR%�p��m{^�-1���ۚ�#���[��_4�1�A�,�UsV�	�n�ȉnC�IrB� ��˴�Hu�6%��7�|h�Uf��Iu'���`_u�n�9&V?^t�;�HY�Ժl�C���cќ[�r�k��6{�8s� �!ì��ˊ��5��[�W=w�xx�w���d�2�m�R�j�R��-ɦf�Z:L�s��Y��&ZY,�b:��`Pl�k��+�sk��Km� �ܠ��֙Az�G]���K�ݕ����e5��˺�aJ�_�>x�k��@��j�bcDҵ.V�n��:�N��Wq�@hVː�1�n�R�F5�:��X�:�ˀٍ�	�q5f��Z@V�D-�A�EtP��	�0Ʊ �ߟ�?�ݔ��Z�BcGA6a�\��y���:�W:�9�)W	6��0,FW��e/��ᙊjk��Hk��ؤO�ʺ��j��mj}�Iu!��&�6�^���^������%I=��@nd�\�g�.�f��{�ʒ]Hj��N����'(�]�u8�el��{3����v�ۋ�#�{5�!���^w�>d��nELG��=���.ڲf�z;ƶ�\��2A\+v�2��<u��r��w�dk��=�RVr�܌���
i?C��S�>��U}��[t̳:��un/�\�,����kf�c�M�y�߾����O^�p�? g�||K��4O�/y{��@��#^�_�9�RK�ם�5�n�_��@�{��{�U9�V�\u��T�m�tw]��e2�B�����W7�Zp�������«&8+�q�����y���=��MM}�;���_3�
�w�8�^����}�~����S��H�C�=D�v�RV�oN.��1�L����zCU$���Jl:��~2m�*����3�P3�T�>%�f�'����+e{B~�vd�fb�fI��M�9���x��"�܅"8S�Wj�dM�5Jh�{������ְ4׮n��Z���v4Z�����)$��$B�1F��p�31xfG�6�'E}'�
�P�ּ��#������jI"�C �2J��=�==Ƴ_Q��l��1s2�Dew�q����eGt�qQ??_�!��I(ol��je�=ie)u>�B"�.c�ܣ�!qӳ�2�o�Yh�Z����ٚ��Wmd�4(�&�Y�k�����7�᫅{�K�)'A��SDl�%�����z�]F�MdO3�
A���^��&Ｇ�W�F��yo�����y��tW��p��EP�Է����w�3��a�ia���?H~�I�Ժ��Vvy��p���4O�Y�i�Ic3=�2��Ģ��"%#2�LH:4� F���4kn�Վmf�p�Ă��͇��#����R����W{�0�s7�}|o�9%zg���ۚjCRKs�/s�hB��W�^���כk�b��{�(���u��={{��<P��üjIHjJ�
oؽO)��OA=^w��h�S���$��3��˚T�e���o�CU$Bjkc�����<=�7C���)��W�1�Jԇ6^��B�g��[P$hT��Ӱ��GU����먔!B�
��_Z�{w�78�qͦF��� �� x{�u�7��fṔ���GF%Pk�p�}o)�e.�Κ���@��72 ��;p3t������zJ!B^��ٹu
V�B`�f�[+��`�,������:\��fFdۆ�b�q��J�#�1��A�ev���_Hd?T��>Ǿ�;:�WPy������9�bʘ=��w&9�����Ԏ����}y/�}!�IrR��o����lW�'b=��P�{�C$��ԯ)������s��5����7��j���[�/y&�5� [�.;����5$��C%�7۵��vw�]����wA�\�,���pv܇���3�/:t�g��ݼ�/k(�ˡ���<�5�sfҍ�۹!�h0���������u�u���B�(������ϜF��@�0b'�\GL�uݫ5�9�sm.V�31��m���ز̋͛j�iRlU	�D��5v�#Ƀ3Cki���ѥ���1�Vqa[v�n����f����gDHݻ� �֦L��LbdImZ��n�#v6�����+��
��]a�����Y�]��K5� [�����!2K�v�.]Dtq6&�]pE�3l�pϿ����ꔙ��Cb��aL��F���Z�e�З$ML.��µ��F"���j��Iu!�oM�|��#�(;��f{o��}�ffe{26�y��������=�x�^p���R�#���^`耸�{�1�|*�d֤5!�$����m�}����B�����C�!���؟���z}zi�uR'��L�R{�=HW����X����~u��$�I$Rn]hQ;�n{C�x߈=^���H>�ƾ�?I.��I��s���s�g�.R��c���Y�f�Ar��hF T9!vc]�i6D�
T��Hí�{{2�1	��1�}�4߷��yea*�e�z!t�ۆB=��ّ�M�{�e�Ȫ=�V�[�ZζF
��%���;;��؂�M�p��uK���V��K��^��I��:��Qț��b	�u"*�C:���� =��]w��ל�s���ge� =Q���L�Sl���Z�&�7�����%�H~�]��eţ�\ծ�Z�9c�܀1��/T�fW{���O�z9�n�eT��gS=^�Q�~�X���	C]�&�|+9>�]$���I:���5^^{�&��`�R{v_R�R�M2���o�{�����oo����S�j1��e��&�X:6��LTe%��0�s����e�v��y�����{�2 �ØrkG��� �u=]�٣]���L{�������`n��������bͦz��GM�qb��(k��r.�oh��j��wW���3��,(�jx��==v�����X��3"��wb�JKz��M�H�گ0;w�}y���0�hw�)b�>/t{w�Շʰ%��օB�3��X%��2���
s\V2���6)���+���J�_f�f�޺z��g��(�9�{2�Q���V��m��li�f�]*��Ģ������2�ei��W3�I�e
�Dy�A8s{;Ŧ�Ȟ;O��F����:p��CZ#b���ݰٮ��8�ܙS��sY0��ʹ����l�vN�(�udҰ��i��Z�5aM��B�j�"3\ln�
>��{�r_%��70չ� bׁLg�E���t�j�
��,��[CH�_C��:죴,eb��)t����;V^�ēRv�P�b�B���+8��[�Vp��H�tK��Q�u��"�P��rۚ���pG��������^* sW-����v4,��R;�rj㙇G1�M4b���n���=d`Vu�4��t�u�����t&�����}|u�F����X�YD�����Up���s0���㥗p�rk�(�EQ�����`����vwF:�Sw�����{�/�v���7���G�]����V^�E`Z�(N��K7�휻{���ˮ�ˡ1�&JVk�a���q�V����#�S"+��\��,J9�G!�f�/�f�]\Ip���0�r���轰�N��
��H#R����@]�3һzuN7�/P�G�R ͛��{o�멂���$<��,�]J�X���#~_3gO�TR(c%*,�Ud�A"M��-���Ɗ��m$Y/�y�����1��EDZ7���-�nb�(�^k�&��KRQ��}�(�M���H�ݒ���r[y��cV
�h��^hڍ�ż�1ͮRU���-�Nd��5�swu�r�mo�<��+�wR�ܲh�sc]ݭ��������zh���-=�劍y��r�ו�����V�	�{{lt�gQ�����Vj�q����Hp�R?Em[�o�N���C[�8&<65+*���dN�힌U*��plڪ���I"�<��R������ۜ��ݢ.{T��+ V���)ҟ[������b��	��Y�1tn2�´W�Fj�M(tnl�g�����MY����ƫ�Ӓ�C�'���٫Σ;KE�G^�ֆH�������?}!�-��un�݆���8��~��ܶ�Դ�t5$Ǆ��t�����[�Hd5{j�.���I1�+[�sصOz�=�3({2 ��L�虧v��*l����{W�zn_a�t=�N������2�����J���3)Ȯ�F*�v�f���JS-o%�M�J2���<�a�$���7�s���yv���QTW'�i5W=�#� <=�q��YHjIuR~�,K�_�f�8�׈��[D�i��E_H=]Fm�:��y���������$i�t��8�,�2�jf��6&H�30$$g�m�vfNf*�tc�n�p��Z�'���.N:,������33���sٻ�j֩)o]N5�k�^�s=�V�h�{ٸ�p3.�2wkך�z;���q�\��7w����p��*.����@�z�x^���d�=�V[\�W3]Ƥ������t߷���z�7�%J��S��{ۦII&T�^��N�n&[�v�NV���-��`�����?T�I�ϻ�{�=�����oG4SNW�ٟ\�|���)�h����+{$��|����0��St:C�į5Dz�;S��G�!! �2���h- �f��Żq-v��[%,{(�W\�;d�xs"i��t �a�X,!�, ��\�A{-�Q����]
�Mx&�mE%�K��]�n�ͤ���DK���ـX�;��"JmS���m Ÿ��-��˵.�Sa�*��,uԼ�)s��1LR�	�$�����V:Xa��.B줬yh�),�\�0r���x|�}�����D�bk�6X��/8e�M��S`����ʐђ��.H	
s�}Q��^�̟>���w�f9l�T"9r��\�]چd{2=��0T���u�q�͚��0K\�-D�ޫ���f�»��Ϊ��231f\�<�9���x-􏜬�y��z����dʩ$����
�m���rc��ޅ_���'�FkS���#}QfW�u���j��!��x{t�b�Z�;[�@m���pp�Y����K�[+�ہ�L!)�į$�v�l��;����@�n��`vM�b
�ML�%���8���ڽ���h��V�1`�4]i��#\�� ����ِd�{mR��]���WF��@j8��銴*�w��a�J�g�F�	C'dQ���B��:#{�3{�%�:�d��D�燀�˪��}u�NFZ��R�v]b��B��������a���U�.��ԆI�S}y��_���S�������=�f��Ȥ2K�[<?��v���ۺ�+Ef�Q;립U�����6�}~�ݗ!�I.D�����⟺�Є������ge� O��WI"�NY=~�����_>�z��WaK�.�k��Z�qp�� J9���D��,`�,�̲E�>z�馤2K�븍��n�ĠxN�8Od���W��T���Ի��g�����|�6�iw��3��0=�}u��P�����b�T�Bʠfff����R�S�ST��NI4c{�[�����/�|�sm�+�6��ݾk��&4tɪ���T�d4%J�
��j�G���f�{�g��� O�����C����7�N��d?I/䵲}[�6��Cˡ�6u��|$��[�^�Ir�$�j#Fn�t7�2��%=K�fh���z.��vL�;};"ln�G{}@L�d��b�0���k����!unW3JW\]��l"h�H�sH32�����{z�5R��C=�m�N�4b;���m���}����dfbT��u~��H5�ڪ��F��Hk�`ܠx���̖�E�}Gu ��d�U"�T���e�q���[��Ń�M�ّ��Y��5��	�k뮆�;�-A=�m�g]b������j�ں���|�҇��з]�;��4R���ic��Y�	�1w�������\���Oo���s�T`�(����w~���>~}���E&�3>Cn�v��i-Gn��@����q�T�I�|�t~E���wV�fB��G�ьE6�vٖ$-À�X�l¡�s@�`���qzd�/���9���u�|v�|���|���ߺ��=��?T�E�HK�\fc{�]i���ޏwf*Ý��Z��Y�VC_>5$���w��f�4�_�����{O��4�����pg��5t=�e��H~��$��k`���ﭚ����w�k�v[X=7�2��V�E(��~�몐�~�\����/1y��GV��9fߞ�VO�!��I�:+(`ٗԗ��a���t���(�h:pf�(�Z�N��ua�>X
�aS��{���8�X�L���ws��K$�RwyN�6���?�I����`���\����[s5�, �5b���$Y�d��c�������ii���&6n%By)���h�])���\mC!�^�5�i+f����F���f�L�s4�R�-�T��nGfg`�@י�WMty��Ls��Xmx�USH6c�;R�!�YJ�cKnΌ#��1�!�5��&��d�K��1�XLM��4Vd�6����(���0���\cBne��L<�hU����tՕ�M�s��j�͇��N}���߿o{��4��"�I����*�Xv��ON0��dfb�́�����n���뫷��uW�=v[,��&�$�'��kޗOƫ��.�?}&Pԃ˻�O\;�9O���{�	�C��������bs]R����'�7�#3�پ%�Y�q���^;�wY�S�IHjC_I(3f�/P�L�ٌ�{Gz��m�E������fG�fH���Z0877��z�4��k�8 ��u�^�5�@�vf���$1Zi��9wF��Vq���?I��d������D����C#���j5K�E!�����_f�4xb��7�}��Ɓ��������,�� �ig��U_=�J7^�u�CW|�}�J�sZ#%m�u�F��ӎځ84!��xz��+`֦����;v&-�ˀ-��Q��o����7G�Ĭ����!�%�I�<��K(J�Y����ر`����zCRK�0���7GN{|���%��5��	�x���� ����ޕ���MQ_�I�I/����Ʋ�]�;���fQ��8��bb,�. x�d�÷RF2G)����{�~�� V�L!*�7V;fиY\�BquD0�]�7XI9�u��^"f�f��EU!�A�|F�y��|]:�h�Y��dگ���5$�}!��`���
:�ՆW����ut���;��O7G�d5T��>H��\oG�՚~���.C!�IF,3	��*�(ș�G#�d	��,B�Dk�e�-u�U�Gv*�@�^�μ�x󇞭s�/q�����^^wv��L���l�����1�d#۲��_{.Ɔd{$�|��rS�iCM�ԇ��O�7�/\7έ��|�]�Vy��r��aT㳮C_H~�]H�Y̷~ûK����\�������Vf�z��|d�R�d�}/�ʓ��l*��4'L��.�mT��l9̣KU�ښkI��0HIR���_�q��f)�����{vP��X�=�6���I^W�v*I"�������.q���|���
�p�����'�:)���U_!��x���h��K��E͍����/7#����r\��4k�a��v��Yѻ fb�wq�ᐏiGEº���.�[��QybfW���=��M��:3n9�Ӓ��4R���p�̜kN�+;2u��8n���'5�WaVe`�W�*�"�\�,���������C��$G1��Hh>��كw�^�B;�b;�Z��f@yv��Q�D���YA�`"`ĘHcV�̶�:#u�&l��F��D����ր�=��̯fG��A`�»�����tP�t�Yu�~On��+�"�����S��uWW��ݺ��n44�dI�!h����m�3-����nG������$��J
��iB��
�=R��έ��>w�d5RK��U��{�NCw�kא3 pۖ���HR扮r):+�յꞔ��W�jCRK��?T�QuZ��5�R���'�������I�%�Y����Ϳ�;�(�S�2��*Y���Sq�e��z��.�j�S�.�:3�v��#�*�%U��y���n�^�E1&�B2����ޮ9����k+�R��<#+!���*�<�x>�YI�"ƾכ�h��C)�e�t�35w0�/�1�VM�W�����oy4�EK���'Z�)B�e�5klm�_+����K����}�bR��Vl��G��ctgtf�`��tq��|�� �Y;�.ύ����)|��W�����pf�]wR"tۍ�N��s\����%�8p���|
��o&�C��Y��K�l��e����uc��L��`���nxm�+-V��-�w��'b�-��,\m�uG���'wV��6�W.�,�s*
��!�&�xÙ`��U��i���cA/�eV�ЌL���ܜ�X����2Z��²^��2�e�S�D|�m��mn���5�O�=��v��	����cvh��tkRtTAOj*�kX/#5ȋ�B��s����ed
X\���"'��K���[h�)<�ފ�{��{�:��}V��5V9k-�ަ31N�f���Tէm���]'Yٽ�c�o�ˌR%9���jT��!lNUgL=ϙo��h�m����V�[ݛ�l� 7�˵�Ak�Jy�}|,�T�	�T�ᖳ#ÉK]{C:��)i����ɨZ+Y� �E�C�"S��lZyEC���OGt!mƅ��T����^�2E��F��V����$��|
'�,����*�7�W�wh�ѵ��usE���\�Er�-ӑo{�Z����6����^��t%gv�:.Z}��/w\0nm�r
����+�n�ۇ4\��r(�v���5�.snwgv3��]<��z<�ɢ���0A�\�ywpnb�WK	Å��W5|�W��7)#[�ݸF�u��F�wr�g#�N�sr���"�wtS��7*-��u�H�˛`�N��^�I9v�k�wN������j����Ir�GH�Eʈ�ʮA9w�Я(�5N����������M�m@q�؛�����Kщ���4H����<�y,Pr���J��
͖�)��B-f�	]Y�ReԎ)���(�n
4��jZ�8��,�r�(ن�J<�Y�����^�S:��,v��#�3��cT4 ��E�hk��f�(��#�YC�v[�1�cK���X��j�ƛ��7b�փ�����Uv��C6\ �bԵI�Wg%��]�\��p�v-i���^�k�F�[��J�M��[��]ֺ"�a��p��.��a5�-qX1T��-�)�L�R�+L �b�5�j�&���mV��0���j=`Yt��^-��E�24,F)[��[M��jp�����K|�k�6235�P��ecP�XJiZ���AƘ�1]C#un��+e֋-m��t6��ɋ�Q���-�f6�U�a),�^��XJBӑ�%2�lۈ�voYvmY��e0��\��V�s���M�n̬f������	mƉ�`:�#n�k���!�tx�6��\�!B�(kfR�ѕؘ�1M�`���,�K�	1r���ŕdac�����R�D%p�Z⍬6���7.tH[e��"-��]mu��cj�	a)Z�T�3l����S=��D�^`��I�)�����n!�f�#r8�uPt1��T����h�4����j%	�����H�@��j�i�+35�e&D�D��h�D*��حv�X�[&��o��`Z��ɍ)u$5�5k-��jU\8�p:�`t�64�R.:��]�ɠ�]C�X�L�YX������voVQ\j��ĉ��ͳc�.Z�`��nF� lu0�����l5fz�k�l!P��m�����j35���%�m������0�H!1�&�be�J	l���4�K��F��C"Vٴ��a��[H�- 0�]
��[&{m]f����ˍ�k@���9Q�bS5��\4y�]TT
�`m�p[�!���M��a���tfF�)k����������.��x]b[��J�������<mŇjP�9��MnlݍMZ*���K5�e��m2�k�,���=����+p1˙m(M�J��R�lB�%��k�Y�5̨��Z:kQлX^`�٦&J�v����40Ee�%�R�۶�6&�Uh�^��Y� �h�bŬl#�F颖���&�-���k�D܊����6ѕIq��+U�~�??��� v�ɍi.�X�A�`)W0!,%.�����]4v�-�}$R�E�g���ҭ��©�Fz���@VǷ�3d����y��/�z�5]�vx�C՝�*�qR>��j���%g��y#�j��r�L�ݏs�4��}W����L�w
=L߾������I/�ޥ�o8^F�uԇ��l���g�3�Z��|k�/��v?T��}!���!��ۦ���@1�'�l�'���GeE������Ƙ������P7��&��Č�3[�K���bKP�4ճV7Q&ѱ�&E���刺>�=}����&�{��S4�\S7�{���'�/^鯤2K�]���K��`Ʒ����>�ӕ�UL0��bQ@V����8Y�2���8$��6�ؿI"k7�N��ʃ��a��[������t}}�����⏆ҏ��aP�Z�8���}����V#��ԒE�{=@]h�\0����LS�5�s��C2 �5�f�0�t�O$��q�Iyk�{���W{cE��\4�J,VHY(��7MI.��ԇ�;��ߖ����y8o�T�3:¡֯q������&�-�~~�=��<J����M�!h��ܳe�c��Z�:Z�َ� ��
=	z��$'W9�2�̀�� '��P;G�Lcx=��U���R��K�z�sG�ڰ·�4�V*�=�w�蹞�\xn5�G0�-�qz����m��<~��.�A�ZSc��y#/�Ok!��Vq���P�
;�'15��0��^��w�¶؝��&///4�L	��h7}��� ;{�A0�V�]G�v���1�ΰ�G��W�q!���!���
>�P4���^=�􆼽G)9G�=� �c�!���.�I3�ӶC���29>��
^���.��p��A�3�q�׳3+(��O��?����\�ԺgM�fu��Gp���Yq��Zě4�D�ʱ�`^#���g��2K���͖����g�gm[��� �NwIE�ə��H�C[�g#��V�����Vw�(�(�ǽ�9�)}YS�RG4�ؑ��<m\Ϟ��5!���7���dT�qz��Yٞ���/���/��vRXj�"�� ;����=&{L�
�w��}�$wXɛ&0����:��0�?\N���L�)��۵�f��[���X��n1���뫊��8�njԣ��gG��/�ǟ�_��ԒN�kM~��sꜫ)vm_`��9�#꬇�Ƥ����S�V�=�>��`�����ՆBơ�n�6�WB`�áJ٘4��ezb`�*o}{H�̏fb�����fLl�(;&M�ec�@fFf/d?gy��g�se�=W8��-����^o2g���lN¥{�nǳ1fG�,t�8�u�Xt�jcw�'nEGzr�fb́�)��h�Cjl{3�����=�ѽ��������.�ǫ��p�$^�d���NUO���q��Bz���U��.���́���/,Z�@��P��)]/�n�t����Vm���q��>ɸ�����jX�{�WzN�Wy!F��:��)�P#�{�Z71&$2�Ik���<<�C(�[k��eҺ������VҶ�TN5��K��R7Z��"�s]q+���L�l�J3���R�b]��4[�R��؅#�i��f��A�i0�*�&q���[�"J �p�#Jb�3Gl=n�dfP��f�uM�Ysv�2:�B���Ek�.���і��P-FMt*��)Rj�yJ�16�c˒�t����?ŭ��Ytr[T�eԳ.�#��vM��,ԛ����M�`��y�*�ӺE�=��q[=�ζ�����yr�I�3U7n����%�[�I��hV-���xj����j.{A�P!1�<@�y����w{Eg��;��R�I�J�նT��3j�B��+�}t��́��Y��2�J���h����~��C��`���?{�N�5'#�b���}W�����2G�1��{�
u��@���)�5��{������s��w�/-�;c��f\�6�	�\M���B�e�qK �0ۘ��î�$�>^�Zk��RK��)�꾮�.7:ˡ�=x<��w���$�T��y�	�i8��9�X+�0���.%��s�z� Ƒt�fe^2|H�Ϝ�u�=��ܴd�mi�Օ�ĭWe����U�EF,"�f�Aֿ i��Ϣw�.!����a�̣솟��r�\�.�d�2�3#2=��˹3wQ<b_G�4��m.Ɋֆdf@��*;@yW7ܷ��P̏:��9�h�װ�TX��R���{x���~S�!��K��	)V���a���<�6���a�����z�f/fF�1"�l�:H�B#&&�i�-��Õ+B!֣t�)u1��V4`ة��&bBFup�kݙ���	SLt�=���1���a1�`ϲuy�f@�ř ^vǢWFқ�K �hvm\M�pZ��Yx+h72^�u�'+��(s�} fb�~����7���z�����`��<J+�J�,��X3��pK��xL����$ٰ8�CNk:@��Z���i�ɤ#������f���|�N����{�5���d?S����_Hd;�_�P�gE��BjkG"봞�6�����Ь�����Ԓ�2�H�_��������)���^�n.�s�}�jC��æ� �J@�D,@�&J10�
V���<X���b;�Y��⮢�#e��]k��齝�߷߲H~�\�G������k�d{�����+ٙ�ᙈ^ΛYU.墮<rU;^#}П}���+��T�]H5��u/��:�嚪�Ƥ2I2�<���Z��e�r^�b����4̟fb����vW.��C�TS����k9�>����
57v+�����e�x��_�ú�=٭�Џo�V�tѬ���j�׻dv��**��;P]��|�c���rrƻbG������^O~����I/�%[rV�y1z�7�WzaCK�cm�f@��ɍ��<e���&ŋ5�+hꃛ�&���(K֗I�����f�vP�7Y�d~�����%UА�&Z��f�D���c����X�*�I��@N6(I]
�ج��+��-�Ȏ���]�
��P�;�&wL�r ��́t���ج�:�:��cȃ��2�9����u���d�.����
�<��^@���㘽���t�b��"3��g�\�_���HW�8������x�@�����*z��T��S,�ǖ��̯ Nd/s��̘۞�q�˹7X��U=�)3�KxP����i �@HsZԟR���[Nwj���X�Rڍ�[�v�DU�Y�u9�A��Uly�;O=6q��f���(�S8f�#ҴZ��*���^W{�������,�.l���X�ey�-��X2�:���� J�i�]h�҆Z�vՙI�W�4z���L˗7���4q2�c̋k5�X7%#l�.�+�L�И��QZ`�HZ\�	q6j�\��*�Ԃ�k��(��Pa-x:�.9����z�kM�n�mX�k�r1��Į^�C�a��@!����cD-��#�u%H���6�Yp��rg$ ͥ������c*9��k�K�Z���V4H��K6z�L��ˋMÀ����hC�옇��/��������k��2�"��B��f����!���1p�D�����i�}���a�E	}��ãd��01��8	��@��ّ/RGQ�dX��"i7��A�F�̏,�+��:;t���|�7&�{H[u�6����X���q���#�U�9e�k8��n�!&#u�"�"�{!x�20��c��-p3m
���Di0�L���ׄak�{r8p�A2<�b�'�l��h�.oN����`cQx@�h�p(�D20����foX�'�$�ջ%��v;e�ֶSL��lZ39�bF-¶2��dL�X6�=P�.8��Kِ��Y�kg��Fw<s��3]pP��Mn����
 ���ā2<2�Y"}7\����U�34e�q�[zd�/��m	HM�7j��UZ׽H��2�Q^�$�\������v�M��Y����WqQ��H0q� ���Uu����b10�Щ�9Q��k��ٳ�-��oq�����r� A����� �B���q[�^������01�� p4Y�d 9@̠�ܹs�dff�_��HDf��$��|�'����:R=B����Z��ۉ��d�@�l"3 /8B�� �D�Q����Q
۳�N>��)��6�O AʄA��K�1E�|_s�>�K<�_��lW6�&�4tvqX`��U� e�Էnt.f@�$��!h�_�} 
�T ����v��v���e�1����9ĕ9ƈ���@��a���ȯz��Z�6�IGr������Y/z��;�̞Ӑ�_/a�7َ4B���0F�@�<Bf@@�B� �J�ٽ��uP8Յ�n���.#e	Y
bO�qfj�πOk`8�鉚�]���R\ۼ�곹����9$Ǘ�t8�'h�u��j�,9w��f����2�b�1��APY�����L�w��LtU>��]mIa�b��m)�թ�\zL������\�zE�p��BdWL"�J	U���k�ҋ54���֫v�.���J��i�ζ�>G��nf.<��N
n�P���oq�FM_�1Fԗ���r�ʚ+P���HSn�eV�c�L���xW"*Vs�;.��kN|xK�+�7���h6�P%�0C�9�q�u�l���KS/��͇�˴2�;|!:*i\/5�VIՙ�.���[� $��������ޥeB�����8
��(:�bw�ZZ���غ�m�n��Á
Oi�)_Í����hVUdn6�z�XC1��*s̻�j]`ˌpuɊZ�Z�SOl�*�n�M��e�],�6��N/�'��^K�2�h��z�����h���6\Ђ!�.}l�Ҝ��V5�[EfRN��J^�<j)y]��:I���8�[+{��<���1m��쫴mh�}ji�5Q"���Ȉ��C�ʥLcL��Y
ʘg"�q�n�Nn�-̓��j^��8&F␔�����E#�t�Ԅ���o����Z�ja]oVԕ�4��K���� 9j�/#YY�� q�B%��Ӛ9:�\�;r��,_F8����w+�%�˺������%�Y�*�
��z�<�h�C�v^��;ĕ6nq�<�5c2�e57�s�B�Sz�0v�H�}����u��sW���s�Ą(�5y�F�,w.�7NQ�K�u��݃�w��'u�~=�]�N��XM��v��}�,h�����-wv�W*��C}�/79n|��myvY1���K������j;��7��h�\ѧv�wno��o.\�h�mو�,n��t����DW9��&�����ˤ�.�U�sWu���l�D�}结�L)��H��j1��Wu����r��ws ��lF��2�`��0��yQ�v6�F�$��4�*�����sN��ds�o�4�EEK"���ZJJC�w�=�'8�|���S�@��@�,��K�1{r�y1(�me�A �BF����+�Ld4��!��_,��]� �O�d .��WC�!�B*�T�\�;�:��v�z�
����78R��;�̞���y_ �_��}Ֆ���@:�Àj��\�\b�l��+�6�X���Vfe1M�0���8�E��A�^̏P�F�T����|���S�A��;���as��+�!gn��YcǍ����n��{�W��,�@�!�no����ra¼9z�m�6V1�*A(�C��¡C�
�!��K�^{R�t�T}���Xy�*V��
2x��"���dP#1!
����:�a�$n������ٽ�q������*x Aʄ����Ǔ�.��y3s`&��d�tF}���GN��q흷������	^�po�[���i�t�G�y�3�|�����O�����[Ǎ����1p��@���:�X�9��ӣg�ہL��1���/[A�^ �`��E��J�8@`+� ux3.�ƄL�YtBk�l�T:�6Ո�������2��!���b[91Vxnp���;���9��A8�A�j���2>�]
�Rf�����j|�~^au�l��;11�lT��T A���Fg��^k����N��� ��"�A�����=���%#ٸ�±�W(G5�����dyf/"3���<qݝQ> ��� ml��Y��*V��
���8\Vpܳ3a;A�n�Iw@H~�B���+�hf��Ո��'00x-��;aW �* �^Df%㘄m�HLFd�C��r�K�aN�����g�n�C(Q2�=�᱄�t�W-J���m$�M�z)�eu����fl8��m�q��-�6kb] lL�þ�=O�,��lm08W2馚�i0fً	5�R��,b�dM)W\�ֹ�p���%��H:�p�)tT��_<h7�*�6���K�łb�����R�p�6���
*��X�Z^�&rJ4si0g�ڷB�Jg=M����i��s v �)��if\�k*���3�4qJP�&ɣA����أP���9�W��3dU�Mw4P�����4n1��Xdf����� W$��F�j�͗.�Tq��f�
>z��@��Їߛ�4�}!�d����*֗r��]8odz���شb=$���@s���A��fÓT*99����N=l��_)����+/�:U�^F�P}~̀GNq��Ӿ��hs��{1d*>��:�qH���\�h����&���\��ѝ��Nr��9eǜ��ҔI�1n��J���Ѐ � �lA9���7U�����j�����y���$/2�b�B �ב�s!R��I�qG��kô>�6�dW�w:Ll��U�A7P��̀�}������3R�33)S2 $e�9�Z��L%�cj��h"l&:�֒᫭���Ss�!��yx��s#�1yWY�����`NQ�
��G\�N���R�#yx/����2=r�؅b��<�=��[���y�w�]ma��d�1\��;�����Ri�~��h��w+i�k`�;^K�t7'F��Ps�lA��>��>>��'��n�>El�]�T��8�ǐ ��2�:o���<�H |^���Fb^>�\��9Q��L^^�B�ٛ)a��6)��!�>��2��J����"F¸��Er��Q1y
vj�T1��I�;aW NT B�E���Ub�'������ �@Ddyf/f@U5je���н��t]Wr+���w7pj�ȃ�s!���:���]2&�
��	LJDBM-	s�"�n��.:�Un��y���@��Y��ϩ�{�<���K�و;��}'s���x&`qS��Q�"6�����ΐF���d/��'2<�D�Z�wag�G��>Ƽ�٫��|Q�2NQ�
� Aʄ"�y3)�Ω:v���K�p(�{b��K�CJ�!�-L���O=��*�:\=���SaH{�ݵ5V���SQ��Y�c^��N*ѡn�;�\�5	�_�G��Q[و�;]k���b�5q�8׳"���FbA����+�I��?O/ Fty�܍���g��)��f*!�fGc���Fw�`�@�������̈��j���ю=]�n�qE�e���^ʄA���#1/��S7e���f�
�-3t�%u7Bl����jٶ�2�4m�]���P�L���ۡծ��苞U��Y`�X��!�uY�-��H�sq��!W�w�����L��[�*Ӝ�`��/9V&�s6��ŗ� Ï"+�˹��t�m��3/� �B� ���#9$��������Nr��q,D�,���s���ޮx;n�u��q�<�{�Gl*���G���eyx� �(��1*�<w��Q��F8�ҼA9���uZ�-�\#K���c�8@>�w��:7"p$��{�=��2�����f�e[|�q�[��[�[6#rou��4a2�1;��9m˄,��m�m��uu�3_	�W�w���`�+Ӝ��*�g+�/��P�~���o���!�D��K���j�[(������ s"�\���ﾡ��eсD�+.�Ye����c�]�Av����Y���p`WF\?���n��LBz���9��>��S���#(�\ʎ�Y�À�P ���x��Ç��@���.+�wS���<Y���ڸ��cfv8F����c�&���E���((��5��7�.���<���Z��\ž�=g��(�Q���x���4}����#��o"�J��p8}4��}�T�nF���H�;aW Aʄ"�f9�z ����/�Ndy�do_B���c�(o�g��|�n»8p���AƂ2�@ʱ���n�!e��"eNywg��7n,�q��p+�zI� H��+�4�5u�rn�_	����v��\�V��;��wbԢN�R��}�ϥ��Y�bQ���5�
�v��ka�l���@�Q%�'�W��Z���K��V�ڕ�ط�-ؔ���������%�:[Fik�%�e3�f*�6lFk�U.�r�Y�t�Z��;jTeI�L$�[Ɗ��XLZ��Y�\7�4�MKh�����!-ݲ6��c80h��f�1m�s���qJ���Q��Ь�5�:3.������֟����2RjgF<kqi�3��EÙ��i�2���Jw�?�-�^�쌳ِ߳+nD�s�Z/��T�d)��SѨf�C�]�}��V���i�Qi�Qmo�i��'+�t��=5t�ל��3ޑ�v�L9P� ���fc��	W�B{���@fEN�@���fB ��$1$�VD,�0Ծ�֕vp������d/Nd͓̀[�v�{7c�f ����6�_ʨ�dD�eB>�4�&��"n>���$f@@����q�;G�P�s�-�x[�I�􌣴p@�r����ItǇ�u�9��yȡ�n�a�p]�K�1uh3����\.�h䘨4�.cG&b�B�{�ۏ!�Fd/Nd-���gR�x��)�$�Y�$�O�IL��
����@�dFb@��DwgK��l�f�_ֳ4�&�L���<j5���멠�D��xo#�Cޔ��}����j.�+��+)Yw�\﫸��3I�߼}P> �h/=A	�D����M��5����}9W�"3#!l,�}������!���f �dy��u
Z�D�Q�z[�I�􌣴*y{*װ��/�dQ�g`5��H>�^�Ɓ�Bj�o��S�l��x"8�Ä G%r�q�sQ�b�n��a���s!@@̉��8Nhn{]��\��{9�o��58�@WE�p�Ds!O�|>o�W���]��r)�m	p���[Y�ڂ˪������Z�W �cs��g��&��n���>��*�My֓=�GhT������D�msw�\��q�*Ӽ�|.�ݾ���>zoɜ駎g��{�%Dw� ����dj�VY"�P�tQ֐ �B� fR��C)!L�b<�V�D�/W`N�dm835�ҭ3�/�c�������Q�*!cw��[�p	����3v1bu�c��0�R^-W�b> e!]ٳ�'��S��G���D�8p�Ā�H���OR֫3�$�g#���#{YB�V鱍���z���08�BU�W"vl�����PBe//7�
 ��^#28`/ԋ���[�R�v�o��<�I샃0Dw�%�!h#����(�F�L��~�w�����5�sE��d�H�iWW�Kv�K@*K�^h6hŵ˼��Y�C��B���f!����S�Ӛ�^ãK� f�"�g��:&�tae/7� �Df$	̏"$\�aux���#<A�5��U�lf>�L�n�Щ�9Q��� Fbᙩn>q�4��x�s�Fb�@�_W��}닲&{�r�gi<��%�K��nx�B����*^n���d�R7#yy/P^9�-Tj��͑��PW45��C�f�"͞�MFQ^S)t������ʈ5�a�j���r��u�OY�춸�J&��x�%��H����ҩ���s�{�P���9Ё�/fG�f �̋��$%����637��M��<�^���@/f!LT3eB7d�L�(2�u���YTLR�M5R�m�Kv�&XS0�FjAD����}[��^9���2���/WT���0Dr�v������)j<@�n �1y���^Z7�cNy�����n��Q���G�5R�l�ӑ�|�2Q�$��s�\o�6���Y� s!0����*7��#;á�;Bg��B\i2���8W����J�7S��Z����x�s!m\N���;.�X2�G	gs��V2{U)�y�B#1 Ȁa�(36���mY��^�f���u��J��� ��D_@@8Q�E��1��㊥�28�ݡ�R��f���íg[w/�����E�V#-)��!�h��ԲsZy���0
���)�$�I�;4�f�1B�ޑ��<�k2acn�
��/�s�2�S{�w�z��t&�
qU����ܭ�	�샷pK��;�s������V�X�
�ޑ�
N���Dr�؁+iL��Z�U�y�v�=�i�!2�%U��P���ҦF�Kw3,ڹ�v�J�`b�S��W������dܫ��],GB�ͺ�����c�ʹk����޷٦�u���"�HV�ꓸ������]��;^(엙���I�1�:�-�7xY��&nY��d�ۂ��>Ό$�e�}ݲ�Z9�LW�sq��]W�9�c�&�>{�3�E�M��������Z�� ��l�NV��X������y :)֙��9�Vor��Jn�$�̼��B�;z�C3C�uѮS��ڲ��uq���Z�[�6w� ��,wK�*��j�n:��S��̕�l� 89Жs���
�Ddj.nF!8m�ٌQ-Jo��n�:���#���sb�|v��=6�A6�H��p�3�[��:FI۷;v���ȷ��õy�*�f���p\���=,@�Uױҽ��S%��}�Z��\;v7��7:��"��S"��it�`���bx���l�n���*hɻ��|�/q��U�ȾZoh9LC�����<Oz�),�[����]��8iV���G�R]� ʘ�鹺�ֽ)�K�D%t�S�}5�gl8	k-S|�Vw��/7r����+���5U�6R�"E�Ī%+'uЮb�s�48\��d�u�WR���1	�7u��M��ۧ:g7I�~���t��3s�ֹB#\�M��L6"��%1K]ݹs	`%L�-9�\�|�F�rSe��F�\�.t�|�"i����ۺ�LPh��c!5���m�!���6$4����N��:�X�ӻ�N�cb��yh��O���6e�':E�(��t�Q�b�"��#`�S�14/uq�wI]ݣaJLDg:&ja�����2���&!�.s@!c$)�r�3F$���wu�	�9t���z8�m2&Dn���7u���FGwe넄BS�H�o�ѓGM�+��\j�h�mq�� ���6̴ֱ֭]�o:�Z��n#+��6A�;J��j�p�1WZ��)s�&��s�6�C53�Jqɛ+6�:��RJV�˲B�X����e�u6iX�9�4��SiX+�ތ)���F3Z�{L��"vbK�]*��������^�49i�	�T�Y���s[
$,34lіVk����鶱%�ZBJh��2���5ֺY��F�Q�Rp���as�jX�̷Pt\�\�҅�3p�f��j�̈́b�2Y��G&Ч�X��Ƃi���Fc���,�#�b�m�%��3��ڕ���	a�kmÉMv�Jm�%��#��c�R'&�#�&���eԥYD�h��5lf��ITZ�`�΢�h�D���͜�p.(F����*�E�H*��6T�#��XlB��IhRZ8�a�)e�[�iX�ñiZ�71b��q���P�&@F��	F�[�$6ܙ�8���%�8�+t��ql�Sg����-����n���̆�7,�5\��� 1͛c���]��u�L�h��B��]��a�j��@ņ��ר���``���ˣL��R��Ԛ6���H��0�t�+�۫B=�vr�T�&�kJV��,1�uv��Yf���1�cf�lj�����`���iX@0-e66�&2��Uĵ"#�z�n��-�h�Gb��4��\g���+���<Rx�@�l�3mf!Q� �p1��
���1���tՄ�ҶU��XP�z�:lĦ�A�.�kl�ZJm`*�B��6A�e��a��A�v(gQ5�Q�V5u��c�у���6��(�`�`�Nȓ�n`q^-�g�u�D���\�nqX��G;���{W\vf��j�Š��u�1m ��-[�W0ɭ�@I�eK�&�ѭ�#X�/[X8닉��6L�@��2�
�B`�3�O<�h�:͝�1!g����X0���v����uaIn�������+m�t��4�..�7s<�`Q������٥�6�K0���$�+�fanRmf�іdF-Xf�j��"�S;TK3Z�K����-������/Z51t2jE1�mX(��S�[�e1��L���l1��䭄�c�%�Jr˔�%�LXgr�����c!���ID��c��`Cj��i)*���ቺݧ��c�at7\'euaa�@;9\�ljBf3���?��m�P�9w\.���fu�c��V<E�EJ��j2�t�tc����f�4t�F�s!r0�T�ؼ}mP�@ܝ�3�r�Y�t���QDŐ�����ÅĀݡ��;.Go�h�@�{�W���ά��X��,�|�dV��{:�2(���` d2]yo�r0��K�1
[�K��!���O5��ح٥Jق�NB_ �(Nd"3C�F&\Q*jL �)��[�>����6/[T8P6'hJ��9P�>t�0����L�#��K�o �ÅĀA1{n��q�D1�����s�o{'�'�\��^�����2�9F�`�#�ޒ FYHn��5V1�6���pJ��]bg��U�*i�ֆ���uڴN�Ӝ�s���0���;�zjX��"ǅ��}{;I��{�,x��Dyʱ9˱x�-4��8��S�M�%t����e[	+e�'i���j�E�۱��ݗ�r�E}m�1!ʁ=����U�d91f��q���rw�޽��6��>"����[T8P�3�%r�EƐ��A2,���y8svX��c;ʸ'9E�Ǎ���9�C��]����j�S�Ҧ����Ax��<F f@�^j���`�nG��8�{Ax� �lҽ���3ϖb���Vυd�K���X���J0��p��Hp����0/P6z�Z`�u�vc7��(\�� NT A��e/�V��x;!�8��I�4�M�����؉Hֳ��3DH��j�*��ΕL����@.�y��(Nd/m\f�~�P��0GD��`�a������G�q�� A��e	̄֮��Ӥ@�RBm��1��lҽ�����3Jق�	ʄA��p�t/9)�ù��,м�A��H@����F)��w��k����z.��T��s�l�\�}s�Χ+�]�^<㙄��f�=e����vܮ�T9�6�[���ew_n4�.�iV{����|�X8P�+h%���<Bf �Fb��X�px��4�CM�+���&g1=�<�=*`�����h���;U��'�.��da�̊�!x���^�����rC��y��wr�j�b
<�G��A8Ps#u����������=��G2�X�͡���\�J�7d-����F39�GM	�?>I�{=�B~��FF4����^,�hX����%���T�Na���_¤?Hi!Dy���DC����%�P>΄Y�g}�<�=*`���С�
��eՉ�p2�d��!Rl�v�@���da����A�	�"������ӕ�stN㩚�؂�x��}|�A9��FbZ�WL�)b��\y�?�S]�f1���&��[B�^"��ɢ%	�Z�`B������"�٥�'fR�Ӥ=m���X��V�YDHEB7(�D̜�R�S T�58o�N�=���w�X�\D|�Z'9s�"&��W.u*C� �c��wVu�F��9b#���"�G2 �/;9¬�u�n� }�(��)^�D@�)��E�\��]�Ņ�L��ˉv�恌�W/���zϗq�^^#1yx��9��3�N���d�B�.L�5y5�{�b〈'2�́c�T�4�g+˦�<���U�a�.Y��ݘ��̞�Bĭ��9P�"�y�.b���5����;x�"3  r�>�Ե�}�<|2znr��c(刎�@��<�"����^@����׉��M�/v8�� �^DkK�1�ns�gp�{S5�� �P�D9�����d�P(鲈'�"3�!b�E22ҕ��otI
����w]��PlR��r�x}q�"3#�1=�U���	U�mz�<\Մ�o{�Ed�S�j�=���]ӮhT�P�a��џV��򎴝|;��&�r��7�O>�����$��&�屺G��&4��᦭�E���e�Ij�t
�9#���YGA���њP�\+X��3j����k�F��v�Q��R,�7@���f[6(&I�1�m����a��[s03�iJ���� (�\�))l�\KVP��KC	o=P)i�a\b����tI��B+6,k��.L,�D�ڍ)�q��������~ۨ�fb�j.�2��sEQ�x�,і�s
���䔺��+����~�����d�BWɼ�+Xrr�D��v����&����>���9�����2��53�C���~�E4�4�����k6��'b
>�]B �/a���/A���#� ����@�B �8D¾p3��Y��ј��tЋA.@����q� Fb�1p�@�J�0:֜�V� A�4��2uz�gu�gaZ٘� ��"V��ވ��lq#@�āCb�0UI��k%q�{�n;�)����}&�n*�v ��\"r���a��Z�=������	t�f#�K�Mvv�R�cm��]cQT6r:�-]4p���� M v@���SR�"���Ωb�hB�*c*M��x"%��~ ���M��CW����[�z�����2ba~:J���w�Q��S�ҹ^��7�.z��'�x��pW��h��G�'oQ�Ȋ��͝�h��Q���"�ᇁ�u^��곰�ò��G K6@^x�2(x'.лۥ#K"@"�<�(���"3^9�T0��N5SĜ�a���vfrv �� �e� ����$6*K��iP��54cU*�A�/FF��=7��u!.6�.��@�y��lX��42�^9� pAb���
]X����b(�Y�����۾۪א�������9��P�B��[c]�]��VC�Ҁ�M�h�m�͡���K�met��ҙHm��]�Yy5X^��3��gDfG��Q�w9�s�����N�(��F;�v�N�͈�ܨ�'`#Ǌ����
.H�GFS��b���A#H�C�ՖgE�q�!w��* ��!�ow&���yDzN>DG�V"s�[Ǎ�r�����N�ad�V·��*�:�S��.7��e��vY��7�m�BS[s��q&tfd��^��;���HH�8�7rn ̪W��l㜹z��m�Y�ef�l�A�"�#@�ąoIі�2[u$� A���bWVd���,�� �e���]B����ܹĢ��}z�����Yb��X�9eǜ����{*p9&{��CrG�,.����p@��D�!3^#1�qn����|<���r�Z�l��HM��P)9ư��mA8՛l�խ]Z�]��m�љ�X#�e�(�d!�z��u�W2����uo{�w��"���/da�f$	�7B��#H�ش�	!U"��T4}�ߥr�w�ɖ�����;�6{8��f�<bs�bAIp�1��20���W6\�zd]�����\ ׶1�ڸ���Zs�\y�.<xؙ���@j�������<Ps#j��_u�ֲ��� �d CY�I��c|�Ox���81��bⴶ��~��l�N����,�xa쬵�zE��켼!�Iu�Ô5�O$m�:��{}���>9��9Bf?X��3��n�Q��;���Qz��J=�	��A� (A̋��5�Liy�֨��Z�\��*vm�6s���q.��L��)D����HKӖ���>�A��8B[Cb�1=��M�ȅ
ئ�Pڱ��gF�G����d�
�;�AՖ��F��.� [����=���2Q>��Bb��.������㫠�e<D������@���f%㘄zQ�x�osX��_l�h6��Px�B �9dA�̄�H1��Q��螏�A���b󫑳B؞��n#dD�@����]t�cz|��N/^�^��
�4���L�����F�i�ٱ>�i�ӗ/��$׆��]l��+�b���;������+ʣ"�����b�/s:V�g�r���X���3p<1�Czک�Eb[�f�I��l�}������:>��ݻ�A\�J�0i���$�A��e��e�R4�xqty��k�Q��]`�uMl5Q�̹Dt��R�Yn��3L�ʷ3g��
V7#��Ư���s�ֺ�Uqcn­���8�mi-��N�\�MYsa�%r[-���\ٕ�uN��ūF,Iv��c��ћMJ��mtq��e���,�[��m�B�K�hj
 X�4ҥ.s�)b�IIY�����>|!~@��i&�iB�2لk�Y`:tj<����K������D̰�=�>�^^#2<���k�3K��ۑZ��T!vw]Dp�q �A�>̄�As#���]9Y;�3�^�:Vzh[��Y����"{��^�^@����S�"��u���A6�x�b�NdA����F*f�8����*u[ ��/Fb����2�Җ�MmF*�ȍ����A[W����5���E@�A3���V���2R����7�ā9��A.���yI��������~�ܼT���x�ё�"y����fG��A#K$��w�9UQ�OBQ(���JI�
�1n³U�X����R�ӭ����Hl���;�׷�۽�
 ��Cj�ͽ����m�ٶ";�B���8�m@@�}x�3( Nd"W_fz��[+�I�x��(S
��+5[Pó/дn��.�����Ӽm[��W��A>GnSwă.��0C%d��^��+D���V�^��Jnu���q�x�^�ѳx�`��ȝ��Q�A3��9�ِ9e�T;�2��O�t��Ǒو s!x�3������j�N�x͋�26DO NT"��ey{29���#'/�����q���w`/A̅�z��;~�����?Z?{��J�*Vb��@�B ���Fb�̏Q�����r�����ݤ�_nD�7�J"A��9� s  A2�#Mu�����F{�bmD��
k	s,
��P�\�B4KV-�
���(n*���=>�$>��4��L{�@���s׊le��:*�'L�=��v[㋚*�-�#Z�f���A�	̄�YB��P��P�.v��W�vٮ[okU��@�f�ȋ��2):��U�Q[�)��j� ���=Ё1yx���d
���6��E]�NMpI���j�d��P]�d*�9W�%zg&V��tk�̼�<��_"�3����ʾ\�)�}VJ;��p':��Wc:Tƪv�2�8��nNe��[z!J��^�Ǫn�4Ë��_[!�kem,T;N����B����(0�Z�K��{�)T|�T�%�]o3�U�N��K_v�nQ���N���SJn5X��Y�
$�Q�$�L7
kJ5�6Ť*�%e8t���E0�6-N��f�i��k��=�̋�j��R�tUa26n�f+����=9p2���Σ��F�֧����M�*釴{z͚'4�<��j�f�6��j\g;A�(E�,᧰5��7oK���-w�����
h����ުɎ�pc���v�:����͋�}�*���!����]�����6�T�\�;����NM�P_��Ң�#��M�#j���].�*ׁ��̵F��yy�`��Gs��8��L���b�J�s��c9�S3�zC���LЉ!zл���*w*�#L�m����og��/���n�ٝ�/u�xm�ЁG�{poNe+?d㓥u^���
�b5�A˳X����X��P89p3VS��t:�6{�g�q��Mcŭ-vqt��'f]�kD�c��l�k�2���v&)T��M�2�WI2u��`�v���\���8�ta6{�N�����5��ۦ�;�T�D�y*���Ÿk��Cjژ�R���e��ņ4�K[{1E2������hv5��S�fIS���;7��y��v�p���]fv�W�ntL����gˣ{�E�;ݮ"�"�ݸ�1����u�(�2�H�@�$�1�'�4��̔�,�����K!2L��C"#A��]�b$AwtI�w}�2(O.o��Ι�BM	�.t����fE�$�$ �2$�0%b�u�\I���h˗(�]]4d|�_<�@�%fE)P>�ab��n�&bf!$$�9���G:A_.�]��(�$HY'w"J"r����P��D�$f�4��HR\�J0`�t�N��:N]H�2R��]g.ȉH2$1�F���2|��.������+����o4"3$H�т��m��X��D@�&v<��G2��*s�sݍ;|��L;���O<���#2<��oѬc�tM�N�yr�3�ɝ�}b2K�h"�y� dA�̄̀�d�bg�sv^��Z06o���ҹx�@C���������Bd Fdy$\^v���	$`*̢ B&ET��D�llf+�
���q��GE4.s&nҜ�� �� �i�Ľ�j�����.tڥx����uͥUZh�YM���X��!� ��Q���-��(6~��2٫�tV1�:&�'L�<'*p�Ff���W�l$��>�f@�+�s#U"�s���7�q��!^֫b#��� /[^̊#�#1!sC,�+vgDo�5@ݥ�3^�=l�c����o*�<}=���Q�OHΌ�JWMi�E� Z�n�<���ʦ��� '�+��^e���sk��D/�)Ǻn�Lr��c�(	�b���� ��CJ��j#-㳹��B��Ǌ�ᡮWS:d��Dф Fbِ#hA��[��Є��]3�3�c�X�@�cEΆ`L�͒ݒ��*DH��T���d����#�n�9��#��ʭV�G"�zd.mu�ȞeeK��%��(��i�����:$��+����.S���ݦ���P`����/8xB��x��b�)�	��Df/fG�#���������P�G�]L�g��T A��#1/�8p�1DZ�焋��KV�~�kG*�����|:x���b;l(�	��G�y�у����d AB�� |s!F3&�Vo��k�<|�	�ܶ/�WiY�+*�<'j
�5P��It���� &��Oe
��=��a�����
���c���>h�o]]^�Z���r+�v������#�eE�-�S�xB�Ѝ&�L�l������b�WYr�Z�5���@�l����������M��KHYt�m��hp�f����vȲ �5�
���Ղ�]Z��x�$΍ց�R\�Z�\`(Y�����#u˓+�8�����)N���
�rR�xwk.# �](��`.�!e���Zͥc�(�!̛ f5YU�K�3	�Yb�������\0у��&I�Y���˩M).f�m�Е��lhܥ���۟��=��~����w��^^�ۚ���j�L����w��� �Z�!���b�@@��s#�{qMgα^=����N�c9t8ÓQ��q���9�Q�N�q���^t �Ǘ���嘂յ�ž�ؓ��5m���QQ�$�xgs�@�x�@�����Q�����ӑ�U�dyf/ ��i7Q�>W5:d] ���:�Y3Ɵ���"}��/|mH �����w4�*}����r�q�&�i��\y A�D�� Amz���C�Ό�s,J�N�il�ֲ4p:��X7K�EN����(k� ��֙����a��v�G5�m������N2_.�DU�(��'5�sr����g�/�^/` A-�$6� �DA�I
��9Wx�'s��txj�1,�7�t�ぽ2s�yٛ��7_Y;`�Rkw�@_�E�;�{�ܖj�OhF��	;�>���Lp5��^@l��Ml�Z�蹩� ���.=�=@��r�w�f�>ꁦ��RAmy��m�/*�:��أq����=,�ԭa.@�ˏ A�D���yh7L�=o�r0b�#_/O�AzVէ]��:�iMW�v�
���{�?o��]@D�RCh |[�/@mȒ�oA��;�brW����U���x���Ut�r�漁���Bu����~��}'������s���U�..�ԗ	i�"�%��*`�9�%�m-�!�.�g�Bq�#5p ����ɛ{��u�+F���HȜZTe[�}Q�gb<�A�D�� ��������Q��1%xn����5+jӌ���V�uQ� ֤��Yfdm���c'm!>8�{n��N��܉��,��F���X�J��:�ni�pyͧ5�D��C�l��[
4�+a-W��7�Fk�޽���s��std7��˗S#kF̪<�A2�����ySΜ��2
��A˄A�C!ۑ>!��Q�}��A1�Z�;�#�J ��S��ʜ{�Ց��b���p2Y���tW&$�B:8�mȐKp����Z�|}( �kc�^�>��]TA��:ԐC��Y��ګ��3���DF�iv�f�.h����+�<�RR6)��ц,�z��$M���ś!F�ϛ�6���{:�XgW�Ŝ2���A�˼S.�P�/���>>mq��Vj�R2/)�౐�С�s��QoD���/J����<���D���-�Ӭgb7���Z�"��>}@6��mȟ��(�0᭵�i����u�YYuPLw��RA�x���Rn�̙��.O^�"|{ad 9]��V�buxLY�(Z�e���Q�>����k��, ����)�5��A�|�N�m�3u�͚U���h)$�ȩ��Kb�y����DokUrB�}y-tF��H��e�A-����e���w��w��j��������
w�@:��"�In�p'�ƙؿP�}��xOp;��KL���6)�]�cTra1�$0���;R;f��R4X^�>�`y���� 6���AN�އ��k+.�������n�k�:j�#� �+��[jA�p��rL��v{:�@Z��tm���rnt�*�}��28�CoP6�ÏnR�҈%�^n�Y@�[j<���8M�UW�WlpȌ
w�@�h�A���qd2�D6�}�������Q�"��uz|��M�b���6VUT�8���;nz�N�wF�����^n�%�� ��O�qU���J"W��M�.�n�9W:d] ��@��x6�	��i�靽�+��6$Kt�dp�"��{�55�9e�ya�vt"@�ug<�Z�3W���kj�}�:�
�	�j��j�*!�Ƞ]���'���pK�f�%3���$�!�
ݤB!��M[�et�R�:��$�I��;��h�$5��I�RiMU�ռi�i���.�C&n�\�t���J�5�����mEv�m�d�� �1�f"Ke����l3M��iRb�,m�Xlnݮ�keSɢKc�D�ցԚ���c5�%1�4h�J�f#EX��[nʳ9Nц���W*l,�=��~LlY�#���3[���m�6���ƴ�ҲRMPK6�p�X�={�d��{�!'�#� ��S{Y[�W|8dF#;�g��7drN<3ٹ"A{�ב����m]�s*'z�FnL��hN�7ݙ:��l���1�&^���"��WbA;z��/fǑ͹[���^�nx�f�}��^�������k�B�e������E��9=�L��S4�,.�G6��mO��k+v����1�%rQ�h���r�V���/Ck��6�A�^ �ב���X�^�Y���}�����\+ʨ1��j��A�#�ڞ��H댴�����h�F
��ݛL�UN�)���v��vJ
�e�3�w?/|�{�!��~{���|k�uM�tm�z8�ؐU ���bH�	��g/ C�����p�S�D���	k����f��1:[w�YZyT��,�57	�,�00��qQ�%o�,��*ˌxfoE�6\d��R�ʭ�0�&6����R,q���A8ژ��ٛ�21)[�Wy]G��"Kq=���*�!��W�Y2	�A�k�k�A(;�w����������U�PbNj��n ��Ԑ��|8�8��Z�V�q�w"Ä́!����GF�7�FZ��WO��
��n��%L� G_H����
���6� �lT��E����Du�uj��$�u�]�	u^y�$�[]��w����]ş�HhR,�Ф1+u��E0�2��I5��ަ�8�����g�O�-������ې'�6���=�}�������8 o�]*��3S�T0=� o�!B����?VΑ�w%�u���w/)雎[LJ��2�lH*��r�s��mX��ۑ�� s  �9H ��@�Am��e����p"��V�����i��ĕ���E5N��.�w`��m�y��P[���Ԣ��{y�����;�C���)wWzEB8k�G,���cC����� Au^y�'ŸD��6�B��s�o���/���v9��
v�ve�f��S�L@�&sT��o>�� �N1��@DwyI�^-Ǒ�$���1L�P3�yS;���}�e�ؐUw��Dg/"r'��ȑ6t�=Z��3��&J�&����c�l�
��:��Z���#�Y�3�*�3�O�yzs�@�  m���Y<4<IL�\�u���{H)Q� �������6П���s�����X����>�j�HǢ힦RȀ&�}9�H>|��zS� ��q��ε$_/ K��!����m{�b��
p$O`黨�/����bAU�	˄���s>>m[����=Ҫ#o��x�pŶ�.��d���)��	p��Q��W����uy<T�5�)z��Z�i��F��I���`��5e�b��nΓ���9.�ɝ�;�j����)�.��MΊ6eIȫ���@>^D6�H>-�7�f{��V�uV\�{4�wV��6��U9D���j��E�Am�;�x������G��R�	�8��m��WlF��t �n�i�M	�YFږ�s�&c�~n����:}���>8^ ���fM��*��W� ��8��̗A�Ȍ�3����x�[jH�&�{6��lW������]�l=�����R�t%�u^ ޹qy��2��K���}��������&n^��G������45�&u�g@E�KmO�m	�oOln^OG�D�ȟ�D��7Ӂܞb��\r��VP���<�p�߻;ؾ�[�>{x�Am� ��^-���5��"���j�*sǟed��T��� ��>n,Ck����OH�W��j9�s�����͸:�
���c��Z�͙f�ia�Ց:�V��Ʒ]\����1��
ͫ�mgk�Ѝ�N����_Zw�m�K3��s��{�\7@��	�ȓ��&xdhM>%�A[*U��г._7��s�z�
��zX�r�uP�fƓ�[8��Y>]��>QfƵ�X�ېe.� �١J��{gc��4�V�v_�h��|mh��hܡLmôI�����/h�:t���1���-9%"%�������r�h]fD�r"Ed-^s��n-��u��� � >9�ו�^�*�+;�pO;��|%��f)Ir�M�y�X+��`�_E{O�s��Ի"� WQ��)��n_R����b�9$�x먎�Չ�1ǯM	���Ƭ�Nd�[vH����c߷M���HY�j,��z���Af�"�7���5�J�N�(u��t�N�G:�j��I��	�B���T��56k��Qd�s[���8��eN(�C�ᩜ�w�(�5�K�Ɏ k
ljB�h�])���wQ�/��m�W��4h��j˨oeB��v� �jS֥�i��.Y����h�*rA��[B�Sq\� ���*��/b��;��Й����J�&[�x�ݑ�5��de�br��e_Z�3���tZ�Q=ͅ����"��+���!�qG�fe#��Toq��.гC�636>h����b��_g-������޲&��K���3%Xq��{���M͝��lL�5=��G.�0�v��_���1N����R����@�H  >����i4	�rf�b�'u�L3��I��؆�.rC
)���N�1;��I$IK���	$d���餐
F�t��"��8�IE 3$�*Wwb%&��1�&N�(�q(#%�I�n"h�E��a���yW"Pwm�=�cJP�7���)"��E�u'wf�뻴L�$���r���5���|� ����h%���/v��Dh��ĲN;0���H�D��LRm�J�ϻ���"DQ�n�
0��˻��\(٤ϻ�-�{���6+$�.sN�lPh�K����]�D�;��h)�	�scE&$54��'"�v��IcQF�l\ۉ���m��8͍��$��@���b�sS��(�'@�N���wϚ:i]+���(�
i\��2�[��c�#6�\㉇Fl�h!���qM���k;`��5imBe,��B�k	��eh2�&�2؉t��F�h�m�n W�\38b��wiT�S@��.*��[t�ح�����&�XJF�nSd��E�1�6.�uQR�m"76��x���G�n1����+K](r�,�2�N�@�3\��K&��TΆ���l��9������ff�lͪ-aUŚ�C,�[d�����p��1�퉄3٬L�ҵ�R�CM�����v��#hf�U�Y�� �P�.q�=�:Q �WC��Ԛ��!��1e�1l#6V4U���\J÷�m��,�C\��355��5���n���4fm�; m3��U�yܺD�(�]`� 0ڌMe�0�T���e�D\[�a��Q��y�УI�!e���a�����+W<�&!��$.�0��Ӱ�a\���#�U6����3y�6�P�Å&���B� �����ec֑%!-[k]�	K�V;a�X�Ky�R����lj9¶�.�&�.&��A��p�u,m6D�2�f�F�+V�3
f).����&�-�K1�	����B%��ś0�\�(�/���`u��ZS	Cikq	�`�^�f;��U��F��nD��p�l,��/mVm�-,+4t��)��Ѱ��(T�p�V��2����
R[���i�����3u�,��FQ�W$[@fA��%%�my�iqL�������@ݶ� �[-���"���3Ñ�58	�7��ǘ"�X�܎��sj:6�HA�A�Ye�1N�6���Ys�"LjF큔�kJ�Bi��)�Y�h��bk��2T�5n�u�Ök�Q��Z�&����cf�&5�ڢ��$Ԕ�Yh�X���ġ�m�y�8F��/��i����X��l�m���Rj�c��1��kUL��e�K3qX��m���aĲ�vi@eՑ���dt,�s�PF\ۆ��h.%^
3e���t	YV�ƶ8iu�+e!x���u�ۢ�snq.H��8t�a�����G-M^X�	u����u+���a��*Abl+K#�(D��]���6�׊�pQ�u�X�-, �[�eTt+f��ٴL��t[uvH���եu�0�gP�lwZ�dl,��ZvMXź<"Z�f1R��R��0V���{��w�ߨ�ƶۃ#e�]�l�h\�q�1ã6�a�sM`�ԅ�1v��׿�-��l��=>|����
�k���K��*�蘁�"t�*�*��S�9^�@�mH!���-Ǒ��<;b���������7Ӂ��W� ��\/Fr�!�''���\F�k��4ۀ�';��6���[j:-匡�z֜���¶2� K��_4$�|��6�&+ �q컶^��Ǫ����'�͠����d۾��6�����צ�-ڊ�Iڀ�jA�	n<�-�[�#��s�%��^@SR;�M����ؐjP�� ���Cn}>!��̶�7����1�(QA2�JQ�R^Uڛ��`2]Ll�,ҹC&%�ĵ�v#�ơ��v{ |��H ����W� �ԫ�ݍܬSË�1;�.BwL��ґ��ϣ��A�ӑ>:�myx�܉Ÿi3;��WނLa�s#�>R��1��Hx�涞�)z�<�9{sw�0��NwjO0�s�e֜S7�(=�]y/e����'�5鮮��;���9D�������n��UܳtY��u�"�-ǃƅ��y6�X��\S�R��p9�s��v$\$\/s��n��͠�p!��2ކ��̬R=h"� �����؊{q8��� AuDV^Ϡ���7��dwG�n��� ����qp��zȃ���Vt΢��d��S�rL@�8Ԃj� A-��Bw�:n�b"��%L�K5h���/[6�܎˫T	�lY���0�.H:��azkP'r<�f��^ ���:Gb�v����ؐUw�7�a(ڰdP�/"�o/ C�>��@� |�RBZq��oGE3�(��w�H�r����8
't%�]G��7�"@-��G�ݮ�� ]/"/�ds�ɵ�Cng��&�Dk��G��g����/Z�{�Y9����5+	�]�F�cgm��
!q6S7�T4���:��9�K�Fdw\���M����U^��#$����k�3` [�� ڒ^B38u:�sQ���H�{�Ck�cdv,Gw-!�Q;
�8�DD����t�b�|��"}�x�mI�@�YY�1�Ld���X9t�_���� K��͑%�@����������J�V�5a��1c�X�Մ�e�۪(���dZ H�1%p�LH'�5y۟O�j�/b>����t)�Y�y��43Qq�f�UV�氃�cA [��mI�	n<V��#�E-l"3��y��wr�5� ��O���^6��*&����^��+Ƿ���h/� A�m��u�Y㯮����*+t%��<���$��yr��}�]��v�U�$e�"7z@�Az�f��sג��Y$�Ʊ�!=9���j&�tYE�T�a�a�v�swt��y0���]
8�
9�@��X� �����+%ӻ�|!���j r`^	��%�u�Ƀa���� ��I��-Ǒ͹[���uT���-n����q؎�R\f*uH*��s�������+jDm�̩H��3fT���[����q6��"���8��̥R&f� �ƽ9�"�A-�Q�)��x�1Z�\5�i����r����n�}� 6��m�%�D]�;��?`"nפn��V�gIsג�.�I&O	�jH>�"��^�Lݮ�u+�Q�H�^@��� �ۑ �n<��W�3j)�EC��&�T����\{D6�O�m��(�:��u�yv��� �ҏ�j}P��z�x�1�@��D/Lr�E�\ #a��Cm	-ǙdQ�}�]U���׋����}�w$�'�g�栁e�|�Y�H�0��F�m��ۖi\��'V�<��3�w&\@��Fƅ\�*]gDp0P���w�vV:�G{0
��X�Y�� `^̪�'>��ek��!f,�5�)̹-��1�[apv�`]]4��\h*���E�s@��A��mҌ����j�I�.�Q��6�m*E�h��Q�n5C-B�h`���J�ťƊs�ci��Z
�5�.�0�h��@�˻��L�K�)�pia���ԅfMr�rۗb�d�^I]VJ �T��KL�eĮ�L�ΪA�_�翿m�jM�H��k-[+R�2�������0����.ΰ�'�,�Ǉ����qd2�S#�#4�T��juH*�HFe7�؈��^#^�������O��ޭ��"����f�'��)扜�]�����rh�A�s��lS��*ze�B#�� �A�!�^neN�T;u���3α=ˁ:�'�&[RA�Ax�ϑm�7h)���w"7g���!�D�ϛ�ᐄ���s�C���jW���NnLhq=j��JQp@꼟�̳D�S�Amy�Y;��
�[�U,Ё��#�y�)|6/�����G Af�@�ք���òeo����[=߯��&�TtƩ��TF�j�ms���uҋ���d��f��޽�a6 �kȆ��p.kg/�a�b}wu�3�!Ud�7�j&Ԑ@�A� �[k����y �z��Z�31��Ek߽M(w�y���B�a�l���9[�[Qe�]��J���u���'-�N�jk�I�Ϸi��S����4�����OA�����Uj�jxO��x����m�Î{U���[@,����@�� ��n[i�ӈ����+xҗâ�"\��
;���^���/Ck��r&r�y���ˊ���C�>>m5���c��u�;�L�� �j@>�ET'���+�\ ��Hmy[�ۑ%��)5�����X�ԽQ��형Ƣ�T�R�x����mȟ7`$sZ�N�$��Mh�B�	���chMܢ2Ź�n�� *��AZhL�t�o�>� �KmO�7闣c�@䝼
9�V�gn��b�=dujwc�ͯ Cnd�y�9;*Ә��<Ⱥ��7P^����e�bw�D�ɘ��-� ���-�Wr�����ZF�ϣ�������۝�Ⱥ����O�#�i)�l9�-�4���r�pv�xV��ݷ��{��o�۲�eDPioL�a�X�S���G^�^F����2��Mj�jx	��s^^!�"|Ch"�Fr��#g������6՞ö2�5�A9'o��ˏ/�Vϴ��W�Y���q� ��yۙŸD��6ª*�g��9�o�u�r�Iժ p �ε �3P@�6ӌ���n;`�6"j	��+��TvV��d��˖KF;X�$��Fń5�,2˓!V^��U���X��,D�sF���h���򕫢�)�T��U� ��5[����3c��yٳ>-��[�� �����F�E����q�ݪ�qz+\V��� d��
8 L��^�q1�E�𹛹i���V"w�,��Q۩�2B)[�Qm���5��X;:�:ԐFj�#�ڐCi1�b�U�=Q��"A}[^JzW+��\Q�Wk�PY���ثE�[���M���$�a*����i��������P�1m�"̫9Y�.���Z�J��DN�wx���̌[w#cj�;�p#{f|wP@�@-�$�Ÿ��E�z��<�����桙��
 w�����dH-� ��
Μf&uQ�
:�P�0��nZF٩���Q�YSv�%6��I���+	�!%D�Z2/$�C��!�"|[UuX���p��`�]dׅ6��ܡb���\F8�:��ԂAn<��N)�5.��yymJ鸜cb�
U:d��|r�y�"{;�gDGts�ׯ Q�^��@�x�[h���|��MZ���.�8;xr�G� ���@[^D6�}вT[�9�bk�!�A�^@�ޑ>nkg/���]��Z������,��u}!���>������|۟7$T��ZW8�T!����\;����Q��4*+�r��s^^!��>m޼�/jbÐ�3�kJ-�qU	y1YO��we��Ҳ<�2K��Ƿ�,m�ɹ?���2�l������E����Z��1XD��QmJP�@�13)҃M������ȡ.H�Zl�J�^�`��͖���M\C5�g)U&�8�h�aG5�͸

Q��qq�v��!B�&�9��a�Iuås�8iA��i��\�Ż�"6]�9��0�4Κ$�& ˦�7��ZAf.�%�B;WI���Hj�
��5���)S��J�&�^ά-5��kVn���=��I�߇cf$l��m���r�	Jj�r�evbi�6�5rW#Av���w�?�@���I�"� �[jE��ͅ:4]�N&v�(��]U\k��a�?k\�-ǐmy�BKp�9i�`��óo�Emȟ�!uӗ�u:�}ez� A��g@CŸ���.6��mR�Ej@��<��"Kq�^[�x���ʊњ/�E)ءQHw�\ys^D6���A [��;�)������qr�w�Gv��m]���L�b＜��
8 A��/��UQ���n>��0A����An�>my}h�Q2�qǋ���Ν�yo����8�<z��A�"��	m�޾���n���
�D��BD�h�jR�F�VXdb�x��`)P}O���x��=�_~�>��jSD��6P�̉��#�M�b5��}1u�ι�mp �������lQ6r�SD��&%޸+'�3�&�;(�b�}�w;˅f퍛˨���s��v��X��w�=��:hYlCɓ8p��j�5L��wއ3�f��sr'Ÿӛ��v���y�|��#�>-Ǔk�ۙ�m��G'{x��z)��nBح���A�j|A�Ax�Am�!�
&l�y5��Et{���I�Cq�Pjz�1�;*EL��Q\$�D6ݸ�|�T������|�pڒm[��j�ܩ3��ӹ�@�W���| ���w�>3q��k�7A�V�I���t�)l��M@Q�����h@t��T�\�s���Mc�Q���.-�!������ϏO��Az��i���r�lDx �U�&c35H2�@�-�$7���3��fv�O�\"�˥�������R�P��8���x6�v�*]�1txv���h/�"	x�F��>�'�,��٩�U��N��/,�e]Nc.D����Ʋ�;st�6�b�7}�.��@���9Xd�o�m�M3u^J�lR��@�%''gW��h�u���|�
���^�铵���.��I��X�n���
3���3����G� �B#�[4�1Ck/�V!Y/B�i#��jz������[�&�m�s�cZp6h!x��g��-�ݫ|��Wݘ*-"�O��L�R�ڹ���f�$kx�=�Fϻ^fo)6F%�FV�Ր��4%�8�g2��=k
��d�6�����YB�0ܭ�&=�%�E	n޶¬�2� B�!n�=,}��V���zH��:����w�fgZ(*k�X��b�'hR�tf���p�9�\K��T��k�J���-f[���u[)U����u�Y�]�@H9X�f����S�X�X�͌�s*�V��e�Yڵ����;�;˖N	7*��A�oT���X90�f�F��֪S�	�4���:ƚC�n�Ӑ�˼(ή���kf��⫌yW���H��]���x3��;((n�wڹ����.���ޗ�f:#��dY@rR�+�d�s��N����)�a9}yMv������#D,��5���:�Bz�=���X��T.�%)Iҥ�ڗ�vޒ�؝��4�mƯ�nwq��'�ք�uz�3
���c�)���N�+%�uh�+YR)�j����Y��|��em����7f���

��š�u�DT��|��z���I-�E����#	F"��!��2E˜�����Q���r�����#��!��HQFѣ����cr�`K3�6I���Q�F\�(���\�4w���A	�6�L��L����i1�D�6dVw9��wc�Ҋ���f�g:�ws\�t�(�a�!�4k�����QPl�\��7�-	R`0}� �]�/���C��rM0�c���r�Lđ�t���S!���&�JM�J.��G�LzEs�o���L<ݠ�"@�"*bc�	A����̑�v�E�n��v��!�s�m�66��[�Q!0�^q
�2M���s\u�&i!K�bRF��2�\����LQ�cP��Aj�Ecow�g/Z���z�Y�
9�y٫�ł���DF*c}5q��-� E��O�h/_eV|)�]�b�"|�S��pȒs�9W���9��݄	n<� ��In
A�R&׭��JU:�����cޯd�Y|U$�H'.9x6�	�q�7�����[)	��1�f�֑44�4me3�XDV��ĹB�]��"&L�e��Ϯ��F��|[j�+v�N�j�6���S���Nj��z�A{"A��^@�܁>n)��c��z=��ݙ��A�Û�a��[� p ��׳�X-������cjo��T��	�D6�H-����ۨ�i�8�.�ݜ�Ӓ*V�
��}�r�6��|[A����u+�i�=� �ڻ�|-N�f�6���9Q����b������6�F�@V��61ŰT)��&本#�V������ڪ�j���ϫk��"���Ja�%@��&���s��1z��fe:��4�^ ����p�-�/�h�Ng+�|��ΫN9��m���1�v�9����A-��C���
ݍ"*U�\Iل�]�1r�A�vm#.����L�Rkz��i��f��:�EA��|��܏"7�	-Ǔk�{aQ�����$T��I�a���,�[��zא����7�Ŷ��F����p�)�V�b��f�i;x@����ۛ"KqWu�ۦS�#D��yx���>�<A� Cng�6��"�o������ۄ�4���$��-�@�mH!���voB��ꊞ����q� �ݑ ��myt*5�Z��Ւ*V�	����h�����d*���㚼�
�RAmy�>�Ŝ.����U������=�L��Q�Tyw6D��ɵ���"��5�3i�el��mZ��i\������bԫ�7D�Ň���;D�k:4-��ԆL�;xB���k(Ï�d�z�L�jK��2ֵ��&�!L�	k1��D���cBXf�C"��<��t���˘B7&�ػ	v��,e���i����,�iw4� P6n#bT�Ye���66�hia*2��mvN��աz�h�\W�BX--��h�f)9-
�[el���v��^ƶ�ub���bb<%�4����i1j̓s0��Rdm51t˒��h~�����U�Q���[,��i	�+�E��Z�#�+�q7&J�bD�H�@�t��"3cȆ��|[B�&Fj9���P�f���!`�9UP�&g��E�j�N=�� ���v�-ǑIUќ5R��,p�!���Tz�na���FV�	���\"�^@��mN�s�ւ7�>�H>mpڸTtlB]�ET�����=��o����D9Q���Ȑp�!��CndT���/:ۉ��k�y�'�6���j=����Hy�@�|v��u�k�Vso�-�Yޓ]J�t��|u���q�m� �a�[3Dv�:�K�d-غ����b�+b��p�N\/�@���������Y�L%	���3����5�1�SYF����
���0&����"��s ����5[���mMڷ��zL�}D-�
90�c��glzA�["O8D�����An���eǣC����~5h!���3by�Fu�p�R���;����F���1��D�8�d��ԯ�6�uw\�9^\�i�B���F��U�n����'�9/f�b��_jډ4�Ai��9y��»�S����5�A�w��[s���!��}��w2�q�Uu�Q+b��!�.<�r�6��|Ch#���)9�ՒN�nG�`W� ګ�}�Ni4-�v�Lp@�9@�I���F:-�;��y>^@�܉��/�K,M$�8��hW'#W㻱�j�Ai��n�ړ'{"߾�.�``V#,-r��%���&��M�ev{	S3�X��PR�DH�z>5��/\����.�]j�['��\LlP��	�{3��`���s�:<�=d<s> 6��
 �[jO�]�tT������̀�'�T��o��zM�Qo���#�P�[�胱H�+k�^^"rА[�&ח�mȟ��a�F�2��W;����nf�����P�����髌���nC�tvU�"�Qt���k\�^��v���*r��ص�V�(�in'U�wN����@�	�jAg �[�m�!�����Q�����g���ބǗ�u��l��q1�@�t�.#u�����[s���7:g�y[��%����Ÿ��P%e&�1S�����Ԡm���dǆkC�p�6��S9�6r�m���3 �*J�� [U5�l�[
d�-q�� ء�6g2�!J���ߦo�l"��Cmz[A
ٛ�Z7��b���b�CТ�����^"���mH!�>��!��;��FUΆoa�<�®�v��.&6(�8�� ���m�]\�,��0��A�jA�-�@����iS�P�5k�{	�A����m��� Au^ ��[�7�h=�����-��Av�/6��ЭK2��{����@�3�I%�؉����Ɉ��h�q���33�#Y:��w15KJ�݋��[v�����s�P5g-���m�@Nq�+"�N��2�S�Ǜ^n���n<�>mȒ�	��o��*ח�]�M�ޙ�f6(��A˄9���s�B�g3�ֿ�od�Ϟ�Mbd�h�h�VR�LcCM3���f&b�Yu�`q�+���Tf�q�ϖO��ק�p-�7j�5'[�GR�[�T����X@���W�I݄!��CnD��@����1wP"��m��ZWL�Bѹτ8��Tx'��}�UvNN�]��~!��	� Amȟ�x��񩣙<�Q��f;�\]f{&\LlP3\�\ A�5�Cng�Ǜ�^"��9���U��j�>�^�@�[jEڮ�I���q=$V���]G�"��$�f/��j���B �7W��|�"my Cn7�N�����
�\��Z;3����};�A��/Am������g���44[WGog(���=����du��������jY�oM�zf��	�}|���d�둚o1�
�(Eֻ8V��\�H`4�X���^��̰l���a,î���q�I�t��\i�S�����c�"Ux� ǪC&j��!+�ͭ]�u�t8�F�&�-o��5��av�la[\������f��i��^V9�JIRLRB��bSLc�`Aء���L��*m.�b�9-c�VD�J��ͳ;�̢���z����j�-`iKRh�u�面��&s
2��~[����X+(�.s[��&���F�Mj��5.v&�mb�3�Ӝ ��/Fvϛ����1W�n���\LlP3]#�w),�wg`9qD����k�^nKmI�����>v[1�o  A/Z�v��a:�7nR�V���ΣȂ=�����@�6y>�x���y C��ͯ"s��p�D!IgT���sr(niP8��/K���
 �������5ָ�ۭ��W���Ȑsa[^]
��[�����Jؠf��."��LLq�*zYY=�U�'�o �pڒ�h"ٮȈ^|10�~��]qλ������Q����[�-�&5u(�g������z~ؾ�S�[�9kR[t� Un.X�I.ҳ+�	^P5�)����>�n��e��w��mt�����	���J���*���9��7k��6���א �^"�Tu�6>�'7�j���EX՜CBo MnN�HrƜjj��h3��T�]�]�#�]��y�fgr��F�z��Z��	&ɱ��q��A�^Cb���\D��k��Ƽ�mޖ����}���5 |�T���� �m(؜a���ùQJ�%����+�[��y]G�7dH-Ǜ�Q�+[t�:Lfd��i�G�Z�<�7
ّ��73�qA����:��l�z{33%�l
 ��^n�>-ǐ6כ�"��V�Fב��/-�ʽ�#5pu)j�f���1� Cn}>-��،�������L�R�K�i�Օ�M�!���5d�6�Қ#jVZ�3�L�:��v�f��[���j�^���6�J�#p\��]T�ܑ�����byȒ� Amy Cm	-ǖ�ySu���Q� O�`/V�9�s;�7iP gqH �A�Y�1}��n �v<�6�In��toZ�q��%��w���&�f�<j��69++^ M�N��4g���{L΀9���<y<��'��n�����&!�y4���Aǡ�%�`�t�r�5�۱>-��p;C���e��v׳`P �ڟ��͉u�n���#pT�� �� E�ױ\��h3y��������An<���!�ݲ�%�Έ�sT��̄z;�fv�٠�J��Ӹ��>A� �mF�@"8���I|�BB�&`Z�-nXav��.k3�m٘��p��ԋG�gcA��ձ�#�Ȑp�-�/t]�eÜ����%�`�t����.nr.,}�y�W�͠�[���jH�0�%�Y��bAʀ����ټؙzn-�L��O Au;dH-Ǝ��6�*yy6�@�A�ͯ Cng�6�"s/IUޠ��fv�l�y�@� ��C�Ÿ�[jA��WE�b����U��3�	�̈́-�!�w]�	�9���g��\"�_ݗW1;�]�B&����jM��u��̴�/�Ь}X2�<�4:�b(�8�7�s%U۹����QP�ѷ��׋���-�ڒ1�E�d���E���T�͛�S,m�R�w�B�y�ysvD��x����{jm��w^���٘�Bbb�8����71#)��]K���5�-�6�D���y��N�ykȆ��|F4$7h���.��T>b�}��Zsih �^�@�����@����u����2�X5����:*z��_p,El�3= ���1�"1�%n�2_�q��l@��mp ����*�r��{K�xm�R�o�EO � ��"5��� Amyr$Ue,\����C��Z�|���B���o^t�!��>3�������I";x��y�|Ch An<mȟ�<.�7�L%���]B�%�8��ftH>4hO9RӜ��}$$ I?�HH@�i$$ I?�HH@�T���$���$�̐��$��BB���$���!!I��BB�����	'�$$ I=�$�$$ I9$��	'�$$ I?�!!I�I	O�HH@�RBB��!!I�$�	'�����)��77�/�9,����������0��p     
@                 [�p�  �R�E  P P(PH ����J�  3QQQ(*��T�UQR�$$R(�R�D�P$AE$Q��Uo�h ��ETER�(�
>�Z(��K�Ӓ��%�2v�I�%p4�UU {�Jx��*��[�I�[`d��f�uh��Itj���
޽X�eRUEJ�QU�8
톟�6H�J�̟{rB)R)ﯟE^|����������I*I_3$�yeI'&IRJ�e�� ;�Tw�� h:� ��y�� �J� ���A݁��Y�F ����4{��=@ �� |��%*TJ���>� ����@�ԋ���A� ���N�2
P����=�h���� A�  l�0G@r�3��ʠ�� �EJ��U@T�W d>�݀ �wo@=Ǫ ��@4w`���G@2 I| >��t�xCGJ:.�Ӡ�S�LC�*�h�P <��R%P��BW�'�t:v[�;������hK9)�@
T�}��o� ��|�t�A�RM�K�Ӡn�*�d�     ��4
RJ��0� z�h h �0IJ�        4�j�0���       M���P       J"�EH     4  $ԀMJ�!�����Sj��6������ƾ_[j���%���t}x�w�Qe݌�� !´���J?�� ��D��D@�P(�	��� 	�m���_�_�X<���-A�P ��E�P O�� �J�M�B 2���j����?/�����I   ���[��}�b|�O�g��j����C��~����M����pۓ
D��9oY���9�>c��v��[E9%gK[y��κ�=;{�Y*��7�c}u�u�\����R�tq���E3v���<�r�N^��Ǻ�@H��/fss/oVy�+���і���hq+^{����rH��\��L#�P�>ʝ���ݛ�L5�K��xbı��	�h{�'F��^��>DsY�rz�t��ҹ��5Y�<FnmN�GHf-q<�(FIۛ�
;�pJGC��@�����Ly̵���pj�&՛�ϭ�!�Z�p0.�o[��Y*�)y-]�)�q=�+�[E�*���nD�@v��(O����mh���I�Z�lɲ�2�T�E�b��«�Yۏ�����[����;b�<Zb4��R�B�6&���ˋs�k�
�6>Z��<u������X[C�]q�gMɏLV�z�:�h������ֱd�\�ot�x�W'���8�5ˈ
}��(�:NȒٛ���B����J���f��V�э�͢��I�����s���� W��^K����c�Ȝ7�}�c�;4v]��I����Rv�zk�N�xucn]e�u��j���,�ۖ�0���D��Nc�g����]��a��66i���o-�.�o�W��&ڻPmޓm9��ܨw���&��F�ǎ�!�L��85��m�n��pŃ;z��C��ۓ_����d��;4skU��i��Y�sFiO#����{�c��k<k%.�ҩ�Te����Y�ڳ%,�á��G�h+Dl|��'Hᡎ�����cr���a�svoH��Y�2&��Ï'�c�c2rۭN��C�_6H�:EAҲ���<�.R9�ڙ��YV�/ڦ���T,e�v�BE���Q�q�R9�Vѱ��q���f����e����/5p�lҙ��&��p,��H�V�Z�ظ��u�g�Y�g$&��douL�4uGcx�C���mf�.�ǹE�j��Ǩ�/��O JZzs�5�l����$��j�!�cN�x����͆�5�a���o�j�;�As���d�ShJ.�0b9rq��>�9�6�fE�;����1�u,Cv��-����ݨeakw���U�Dd�*f�h�7wZ0�2� oϧtZz@)�
ң*�uD.$�T�m��#����Y���坸�h�f�F�kۇ��.��qκ�a�n;mx�UR���2�[��\K{��<�i)v,	���v��WMY��oa��z�OתF��vq(GP�pUkP���"��Ԗhy��V��@2�j�k��\�A $���h�@����7{�Fv������3���7�!���|�B	��uSN���#{5v��S������~=�ܩ���n�9u�n�{w�7STm�g������2�XWBqsyis.��ݯ��F�R�c�����w{Rf��{��q˽��١N�1M͋ �7�wB�a��Tqd��4��p�O���[�	[����
�[�-vji��ӣ��x�h[(T�i�Fr��p�N��y{'wws�(��Ë�i��Y�w�]�����t����5v�R6(� �2� �(:����띜��ion9X�W wᎡ8�6M�o]z�-�ĵ�^����Y�Z� D�-#Z�,�Mt�!�OȽzx{�|i#hLv�����3MRL��F�4�H�N���ڕVM���Ӏ ;@��BK���u�7]Ġ{���_	�f�������9֜�H3bPG��Co[�7qo>�_>��U�u>#8�\�nu�Ѳ�|��q�d�+����L�f�v-oc�%#��$�:���=�Ly`���Ov!�<�s�rt�� r�a8DA�r�!vA`����ES�(���t)T(�vrU&�w��v�W�?�y�˯�זr��5��|�產�q�p*�o��B���W��m ��O��`�>�r���h�*��j�e�R'��컼�������/��P`�j�nn���fW
��m�Ju�d��l�l��P3S��.8�&�Ul��5��r.F�1q�����]M�L�]�C�^���%�ʸ�j���ce*p��ݦ��r�yw	�k�k�S��B��.],r6���eG݃Is��c흓�R���n��377�nh�2�a=2p�G.3���X�n��Ҙ�wJᗇs��o\�.3�/���z��xv�r�*��G�����>���w[�3����Z=O7Cz�@ vv��!E���hĀ1�P���5.�0�	�s��c˅����V�n����7����f��;r(*7�80�̓!x_F�zmK��]��5�>U�9�/2[<`���F;��D�*W�3��"�������,�ӦGқ��re���ނ����.P,(g<smM�K6����+9dWYA���7Qd����x��p�u���{��g/�v4��η`�s:��ӻ��P�|1LT���X��r=;]�Nj�.&��Ɛ����e�C����Go[-�˅�)	�.ۇ��]�J���ŝ;!�����w\һ����9�ƨv��4���eE�7s��$���gB�Z�ܤ���M�:q!�Uۚ��z�� ��K�Ew�f��5�myMŹ&���w���ob�3�D ��7sf[�m�Ϋ��Nnwf��R����;���F����އ[C�a�ī��"�OY�E**�����2�NΜ��öwr@
���3j���6MX�;԰m�w$V���C�JnQ �N	�j��JxB�r~�P�
♬�LA1�}s�i�V��f�'�qɛ����N1Y}מ��,�Jj�kk'l�#K���Gl� �YQɈ�s�3�ހ�D��b;��1e�A��N�iWoG��'/�4�v ��;�sS�[�yks��ڦ�/q�uM���S��nl���ݒX���5+�ںX3d�{�>�-釈׋R�ܐ��������(�S��Ͷ)�p[PH�v�m�;�@e�kv^� 5cjr޿�Τ�{�f�q\{�N�S@{�+�<�3�f+,R����Z/v>���[��1h�K�y#���-�;��q�͌2u�kځb��aǗ�;�:^�Ԃ�ס,�K�j�W��b�v��Kv���#�R;�.:��C��W{׏��ۤeІ�<�������nnA��yI�u��[��	�zU,�x�Ip��޸�E�|�b^(��lXܳV��Z��h7�;�
�Q��']��*��4�;���{��QŃv%a#�`>�H�H1�t4�{��9���G���	ǖ���Q�}HY��L{</G���Ӹ�N�y�� ;��ܗl�k��[��t:�D1l���$��{9b�a��ʶ�����鋵$c�P��w��Ei}�J�eH�q±l������dķ�����.���j�K&����F[X����ɮ�P���X��S��G�4��v�i�����2v�y���oB��Rg����5|���otޚ���3�>6��s���O��vjtbk�옵i�s,ٴt
�̓*���Z�Z����p�X�7.��p�K ݃��.�B`*�����+J���{������w�d X۠W�9��r��:P[�)�;�� �j�0L�ǔeȺ2�9�w�p�� ����q	ٱQ�Z����3z�3z�!Z-{t�d�66�E˓5|��*�;J���rcZ���N�(�e���KGo]�p�{5�`�84\�7�11n�ZR5��L����\��*w�ss��#x8�야\��Q��V�p�)AN�qT7�u�P�9)��#�R-cO��&�Ō���I���ѕ,dA������܈�W��ũ�@�<*�X[jr�f<F�XC�'��7/v��J��}.�W^:ܽ�s�b#��ҳ��]��Óy��d��8��9�tl���u�\����I�r���P-Q�gcwV\��/�@��bz�c���'A�p���{��wg��4b��Z������[n���ya��[�ب��a<X[#��R�XNPN����+I�5܊��)�1-`�|�Y�I��}�܇��]�+Ǝ�R���X2�&�C�ӻ�/lӚ�ܝ�X:��ȕ�ħ���� 8���\��O��8v�7OZ�kou\�q�0T!<�'��F����ŅkѢ]Jo�$�^m�T`�W���_�לEd�Nq�sd�4�mێ5/�n����; �~�=d��ygf�)�g���b��惩I��==�Y�l�t|�W��x\�ypL�t��лe�&s�P8��e\cޜ'A���%Ԇޥ�li���r�F��)W�&.�<���\�'
�Yp��b���C��W�?��/���I�"}\��G����=� )��E)()Ai�PZV��V Z@���PT�UJE�E�Q�(�ZAR���Q�DB��i)��PhU��B�DV�P�V�)�R�P(Q
h �U���T�R��JU��V�F�F�P��)
U�P
%
B�A�Q�(P)B, d$|�}��=<����c��B@ !^A<ż������ɳ�,B �4i����q�j�խ��k{�4�f�e²��i4o�X���<���4q���zw�$,�-;������V�X3�5�7�w{ǻ��x���9�ӓ�U�ׄ�V��m'�__
ZF�JܒoMds��+p����o#��{�[��Q���M�P�A��j��������3�w�J{�ݻ�K���۷~���s�zUj�{�-���^}ݏ��֖v�}��.�k�6�B��M�jN<[M�n��0{��Օ�g����=��V���1�2e�t��G�Ğ׫����o�[޹��Y���y��]��٫ q�+�6�������yu�ằ�r9��j���ל�o����vMX���=�7�lyGDjc��>������wKU�Ś�6���7?`�@��o�]��껜�$�{`����`V��Wl�t�B����Ga�]�{n�G�+��i�M�kl���v��s7Ь:}�J�^��7�ge"�&��Mo�� ���rk�X�d���4�NM�]�d���X�<�K�j>�Υ�Cs�8��g��[N곩.�)��\�(7D�zTF�?8{ۑ����[���[%`���rY��n� .��W��1^s������V�زG��sC~=fv�R��<Rw�{�@�������ыq@�!�iEǡr�}Fn��:"қ�����=�3r��pȭeY�8rRC�$����U�guC�z����G�u:^�1]�g��R��OoOs�=���0��b��A��%��6]��VUN�*�s�T�c'_�����<3�5p��|�8�Þ^K�i���y��֮���'�L�8�="P"A[7���rL�:��3UNbI�]����z�Y�s��L���?j�4!/U���'&�P��$9���sdiFS3�ũ2�/h5;wL8�gY��5��Լ9{�T96d�^�V{A�ԧ4�� �U_L�\S��S��	lehSNV��Ɖ4�5���8nľ^�sE�0+����P^�3�( @|7٭���JxQ,׬Ξ�6���e�{��(�q���;�	��ll��GW��6�ێMx�#��2�o/�o���
�����H/Nžt'��v��yA��C�"���鼧��g�w>X«�}��׹�Y�Q�ܤ4���ϯZQ]��gn�&�T�s�ڸ1�3S�^ܚw=��]�Cc���k��\=^�u�g:0�>�n#�v}��%^���7��X������X�=.��Ҙ�:v')�{��yl�j�W����J�-dwk�`Yݼ8
��AM���	=���Te�ѷ9v?_d/&�v�@�$|en�7����nD��Rףr9�����(��򈛚��zj�/'��}��i�h�N5�z�QF�^Q��5�A�6��sJ{����!N��9��{�W ����:<d���^��e>�gL����ݪm����bܾf�m�l��<Y�Ͻ�(��{�e�@�n���7WM���iݘϟ��X~�y��:y�'��̀�K�[���L4�E�rf�oc^}���_]cT���i�)����'*��W�Y� ��׳����H==E	��d�b�,���Q�-���Z|y��Sk�C��I)��/�!<K��̚��Kf�*mm����)-=���wO)�^��a�>ڻN���G�r~H�O��v�M�_�+%�<hj�Xy�	��Z8���Э�B�����W�Y���]@��������������j����|dV�j,ag2���VxK��y_w�#W�xS��\Pa{|�=��:V��4:]�Y�
�[&S�wS'�@��[j}{��`�{ݻ�D��eK�ڞ0��4ӎ��Uw����tdDyx�_�k��_���/8�g����M��/�ܽ�	������عvs���� ���#ۛYY���L=W���@D�a�����u�=Tr5���/'Ke Zw��ۮ�G���5����t)�.q��B;�o�,.��q���£ʏ"҉�Ƕ,�|�­^�a�X�$����yd���tNj���]�Bۯ���'���W{{��v�>����ݝ�����7�'���Wy��W��*�vW�6g�j���=�ٱw�}ԋ��6��Oz���B���¼�ܳ��ę���ݞ�;��~��4S���$���'�Jf���Џ��y�ؕ�z���`�1�����I���oE�����,���<F>M���;ȳ�']3e�Q�5���ܳ���狾~��j��JG��{݇�;;˽y��i�7I���O�C��o��	NO
�}�;���B�q�#��H�H=ǭ���͛+Iy�Pc6i
mE	�Π��[-���:'�� [1��R��Sf���`T$�p�-�D��%.N�Ti�勘^O|��f쬸tw\���A��ꕞ�!x
/$�y@GY�Z�l��n�㯫�ԙ��4|��}�����)��w�^٦���̩qB��;!�گEi�[�h#܏d��O=�>/�a
!����3f���Y��9���-_+��ه��b��g��Y{qq�y��R؃�l�:V��V�"�y@[���<���VRB|
}<�|�3�e�y�v7�>Asg���7�/�%�V�w�����l2䜳���M�Pq���ۜ�9�Y���������td�v�&��Y�7��xh�(� ����HI�ltI����r��8��735C��u��Cf#�Qh��Q}���/�7�d��LO��Gt� �#0eZ�#v}Bkf��w:o��#!,�Ɉū[��#`!a��Х���rg���Pɳ��GU�:`���I����A^�Fm�S�cפ2UG7��Ҕ�� ��J�^�D���S�v�8p}3_�����Գ��:����{]��V�kn��A9Ι�T��ӳ���E�B���o��b�
�Q8wa�Hnď㈕JZ���e�)�n�s�[�n�^C�͋���O���_�0AH����w�����49���H�[�;\\3��!��\��o���qy�=s9UT�=�J7q�q�!�~�{�V�ܽ�n�{x�s�b�f�D�D��*1��|s|�Ƴ��OJYۇl��zsFM�Ƽ�aKv�lbV����j;�����Y�\:�S��Ip��&�f�����q3ݹ`�pם������;��#AU��,[S�N6ը��ڟR��wI�g�d3N��.U��k��b����쾻�z��u�wC�	�l�ϱ��]b?`<7֎Wf5�d���&)⽋@�l�u�úr��?<�r,�0���3�t����vt��W'�����)�t� ^��!۾��Ic�ֳ���4��YV�A��&*B�2�`܂�:��`3�
��ė����՘<�Y�{�"��4i�����^ދ�;���}먚�{iX�˧Jkk�e^�%�"�pRgK�
9����o0�Ye�[��
à[.�o�,Z��J+�Z{\x�B����ݏ���	�ي���/_`˃[�S^ik!犬�n1}�;�M���`#�hF�gNr:�=d)��u�{gC���vJG�3�D��y���ǯ"*C�}�۸�N�x��(ce��^m�M�C��:+�p?�ow-���w^׷;����j�:�l�羚k ����鋙��z���<��哆Gc�;�@k;���/r����{UD�N�kbJ�졀Đn��򡦲�V��.;Fm��.��`��tʙ������5��;�;<8-�4��{����W��;=%��>�.�M��9��]�i�_�;ݳujrmٛʿp7S��s�E87��wݜa����D&� }��Y]ڌx�\�8�C	�al�!(E�܆n.Z순��,��<���
�r,������A��ԉ����y��ܭ�����)ӏOs�~<��홷�bP�gn{������]�l�+�_k���C؜ �x�M6��F��c��I�3���ϒ����<,�x�;�۶N9�Z3��w���#s����������5�-�5#�S�u���o�-@������{�[�CC�=�ބO%��(`%��wT�Ǣ�s;;��BYwu���I�x}.������Y���9��M�x�/ױSD� �dU�8n9(�M�w�X��;��:>��{�?n����bW���?Mcɻ��o�ޞR��X<�۽��(����ln��<�{��K�כ�u�P�����=F��6π<��i6�>s��Ȇ4W�l]sG&��!C�Pr%%�-��	��<T������`�H���Q|6�u�.�f�V蘆f�w���w�G��^��oO%�a��Ʋb�Q?n�x�*�X��츒�u-%�"$��ι5A�y}raq��5}��x���S�b�^\A<�t��etƤ,Д�}2��:�h{�c}�Vo�2��䭽���Z��M:zs�{�W�M�q���#�hD,�g!�儨h���yx-���yF|�R�$����:���_;�=  Ad_�B[�`�j�ו��5��\j�-{^��"��(M��&�fF�WM��PX�h���B�hD�ٍҸbb2jL�/j�����l��{<��:[`fʱ�[�&f�t@��%���|���3`&F/h�MX���Gu."S6ݛ���R�VT�V�V�f�&q�g��,͎6��u���"gW���4qn����Zl�۞1peҰv6e@�7�f���U�y����m�1��.��.�3������i�*���6mGU�*�F�$3��)��P5-�c��d�5�]A(`YF�@�dqT��p�0;jv�u��n�ɉ@�P`)Mu�	ʷa(�PYek��[w)6�����aR˶�$3Q��cJhʸ!il�aE��-It��$���f�bJ$
h�B["�m٥n�Ʃ�Kت�Fm`�����MU29׌�i�]��-v��a�(GmpV�^�y��P��� �
�Kp�&)F��&.�ft2�0�[k�1���VjWK0l�)+�$*d&�m�3q�[B�
�X��n�f�h����Z,s�*�9���.ڍqM�F��(���	�ղ�+��́5my5�ɚ$�e��'�^�z�p�SZ��,-�	q�	\kr&mu�fRgS\8R)��T�Ŗ��9�f��J��)�����v���Q%��&#���R�Y��������Skn�i��tA�ack���0��7��4i��sˬF�4�ͱF	YlR!���0Q�V�,.�.��5�k3(C.bMu)�a���f3��-SAօ�Z�;�l�� ��$	@���c��M@������o�����bhyO%#J܆���b�MA3���kv!���,��m&�ӂUM��NCfb���^/`xi�Иc�&p� Y��T�����s�	un�)�!Z��˃R�R4�4Y������ա����R+�2��!LV�bR�`�e��h�@�HF��jL���#Վf�oGY�l���R�P�e���T��m�ID4s��J�m�6�^a2������bԪ��
ݚf�FM���8��e�،�̢kɛ��RS%�mC��4f�\B�40�c5H����RT�"��q�e��7�X�q�ң�
�	�Ť�Ku��م���Y[�WskuR��a-�M1��x�SD9Au)Պ1t^�[��7R���L-R˶��+Np�T.���� K�B�(Kuݲ�t!�u��BTf�-��1�L���Yd@�l��h̓2�P�!(�l��q%-c4|�����c_/o
y/ye����:ي*ݜ�B#h�T���Z��]�n���"��0��g&��ڙ���f�M��*�-!1��i��%�����p�"b�J8!T�T��Bl�SD�#R�	euF��U�nFִ)TC�rS��L7X��qy� �R¥�)K)MhƸ+�ٚ�jnZF����C2�	p�7]�V�Y�լ���� D� !��.��iy��l�f�V3,�; �#j*j�d��Qb��Blgmɬ�XQp���ff��B�y��v]\�t�n�U�͵�3m����� �t��@"�mv����0���Vݡ�XM��\KsT�Q���v��R�l6�)v��ceh�G92]cc����ź��6`JP��Af8�-�4l�l�����1�0��v��vt�e������U�F�{*E4Җz��i��Xq��-��T�SM�o5Uق�t�4!\��Tx���D��4ICGrm)]��*�R���Ľ�h��Xj5��#b�C����`�L��-��ň�D�e#�r�1�`�n�Ь;`֧,*GP4pe[�)娀"F�-XSJ5�C&�%�kX=-�h"L�+��-��c;e�֋\�W3XJ@qΘ(�
���j�b�6e+-͚Q�P��v��:�`n1m	��ҥ���ʣp5lG[j�5�����Aea� ����`�������`�Ll�
�-�m4�na��
�R;mJu`7#,`詬��LX�ԥ�lfb鉣��*��P�IJ�S�{Lʮ�8�L�a��܄��
�^Ը�.Q�Rip�Xv	qE!�L9\T���f���M��uk\��mtƫ��%�B�6;MÚJ`�3��jUk����H�[a��X��j974��-���lK6�Y��q�Y{Lq�`���ժj[GQj8Řj��n�-���2���{Ԩ�",1��Bd�t�T����\t0�l�F�]l���#��[m2�;P�K6cM��\��k�����&ȺkHZ�b)��0�t6����![q�B��*�]��I���ƅ�nA�v�զ�!	l���`]d�a+��,p�\T��#��a��8�eXQ]I�"�|t��"5
ĭ]�YZjX�)Ԕ��(ҳKf�u!��{*�L��:kb���+H`�H�&��:��J��P�k� e��1f,�N+�A��osrG!�JU��٣�� h�9�˺(�V�%��4�@������[�AmT(b���y1�R[�.#��%Y���ie�v6��m�P	Qr�h�c�\JW��b��P�i����	���1[�`j��o�����F��#��6ۚ�E4�����j괎[4+�+v���r�1HR1 ]+b#"e҅����ZKI���P���Z5l�b;]�V��L���c\6�6]�"����L�B$ŉ6��A,�CD��Qa��"_<v���0m��Si�q*1��WH4�c]R�A1"ġ-���f���2������j��\�
�vS�S`�6��:׭�+���7j��J��t�ee��3q��rM�h��3#�fAB�hҰl$h2�����;f�epn]i]CD���.��3���J��3PΉ��hV�q��v��.K*�n��9yyյˬK��]�f�5�%��TR\e0�ಽ���p�e��M�l��9�Y�2;�̤r�t��˫X���[tZ� ��\���R좳k���V�ҭZ1��ᔹ-y�4�����	�l��1j�l�*�R����+��mʪ����������eڳf0�e.P*�c*���R溙�і�CCL���:\��bj�G���\�a�5��]W!V�`lYcu�f�v�5iɶm��,h;8 ��عJ\�� �8`7ZǔĺңJ�CH�n�R63�k�*YFS,ٙ�nե�|i���y2Z���&f�&����3���[w���3p�s�B��T�ٔ֙ŕ���ܱX�Y����e�;eU�鳴�3�9r���O^ԓ�AI8��Jav�`S
T+�NW9�݂�(i��Phu��0�ƀ���ѶP�҇��^��C�έ��{'��w$�:˼Լ�М��:ΞTii"ywd�wf���()9r9{.��:�܃���"�t��9���"t<󼈯/.T�l��y/c��b��R7���u$���)<)M�h�Q���s��|�UAA��!�;�<�w&�(���rb��<�UG�i)����#䆴���=���P��9*48�#�d���ty`y!�lD�!�t4���II����f�yPh��ӥ��ݳGj4�#O6�4%'*S��@�.����8�䔘�i0m���jkMW�P��ܳU����篠kP#�ܸ�Ѭ�[��9��ݘ�l�Ԧ̚١BԆA�#k����`��v+B�lu��4�am���u�
.{Q�hPZŖ�6�En�˭�Mͺ�)¥.�ԙvvp8ȅå�M�k��ԥ��{S5)(a%��B��V�U�]�;U����F$"�X*�KI��:wK�[�CRƺ�n��"�)��f��6��1Eʷ*,��ɨ0�@i�V��[�u��c0X�P�6\M�"�K&E��8I�4e��lʄ�M,:��[kd�3:!F&���Wj�K��ŵ����5c+�)���"�4`)�f�ZMK��[2�9���4�+hbZIV��4)m%k-%��=L�L	�o�IK��ͭ�U��N��%`��e�,�ҫ۱3K�ef]�mt�4P3\�1e%�5SA]+�-a�M]�ڙ���Ѻ��95��%�7l˃)�7J�t��I1��1У�Uq6�S]rڔ�	��aV�Ylu[Y��(c	oiZ�lÈ�.f ���RѰ���L�[n�[�զl���6ʮ.G8f�n�:7j�-Z;���q��M���E�UUU�P����]�^ufҳYhזZ�U�J7��J�\�ƚ�Bݮ�2�0h��*+����.և^ZJK�-	V�^��� r����6YIQ+�)   �m�	X6��(cJ�l%��]4� !0�hRRl5�l�A�Bґ�B�^ml`��jU $U�_�z�k_�W8�c�����V�R�U�1�������e��Q���)���]˽��2Hrש�|�m�11z/&�x]��qS�{��'9�I�(w*�\�Qm��K>���m���1<��k��N1U��[Ffӡ{��5�g���͋>�^mx3����W*췰��͋؜��xm&@m.ڍ���`D�D�`HBaȕ�*	s�M]��Zm���x�yw��vѩs�b���#1��>m}[)Q�)�s�S��]t�ܱ݉϶�N�[lѪPO�q1O�7N8ӛg� ����	v�/;�3&��gy��6�ȇjm ۏ7ns'b;o�\G[ř�9�9[I��sH�0z׽�v�9�5���x[s�K����}�y�@m�}w�y0�8>�L��DfMg3��A�j�3uXB�bL��L�n%u��ƩX�74�JdF&g���e��{w��t_D�Q3��4ݮ��m����m�Ӳ=�w������焴�ޔv���nhC'�	m���7�v��h��u�NXanD/&[��75f7GvGwJ��wzb�m1Po*���:#��
�y�ux/p����N� d��̶���ᣕ�۝ꇏ�l^��y�p�N��)���!����a̼����|%�n%�IڧݭL^�G�vspčBm�	��"d(ID�	�Q3=�W��m-]d���Zw٘j-�bH6��%Q��6�6�+]������9�Pz�*���5�[M��1�z�q^�w�3����co�k[�6����z��`�vǛٷs��r�/�a�������iڙ��w=j�ຕ���c��=�16��nd����iQ���#���òލ�t��j���b�̇�t_D�9z�n���1	F�B�l��lep��l���kf&J&b ������L��y��w�|�)�,}� 6���a�Uڧ(Ոck�#�+.r��6���Q9(��*�y�5�y���w�}��9{!��}16b��Nm�*�le�{��_�}����hT<T�κ�c{��{5�Um�9����9}�w��<y���t�'F��8Fp�k\w�\��2����V?f����٣PF�؍�&mHn�BY�p�b��4,�kn�,$e�\�`�f�K�[I2���X�h�]B�ڝr2�wj����֙���a��͙�Sw�vByİ�m���D��E�SY��]jW�M�(ZS5y�g5��U��e�et��>��[�jU�c��=��0�1��6Q�"bJS*fw�sC���_\}5���9ݖjTD^�Ym��ɝf�'2^��ns$�V��}�״�qJ����MV�2�i��s��z�*H�:�m�̜͋���ۀ�Gv9��T:�;��}w;q�7�9������Byx�i�������������oYȇ���6��1�4��{E�-=�����(���i�[bʁaL	��ED̬�{!�؇�������ܱ9�nA6��^e��ʂ9w�e���,b'�M�迮�d��;��C-�c<n����i�=/j���W{�r�:�����y�9�^>�k�H�,>m�^Up��v���9�����q�wgH�d�tܣ�z~�|=���#�Ɉǃ`���-�@2�\���;�wv3���r�/3��VӺp�1�1q��.�1J2X.jV4u5�Ÿ��H#QJ*�]�e~�=��K�%�gnhfl+5.6/�N>>�F6����̻�;ͳ���� ��kNr���y|�C�F��W�p�J�}|���l��d~�L�9��`���@��x����y.EO�fId�t���ܲ6+^��ڜ��יX�m�rVlfR ��V���y�q�ɷ�߇�We�A�V��"�Z��u�.F#�6)M�+�2�7��ph<����y���vt�+�Ț�}�Q�k͸|6�N��է��k �u��}��7؊�+3#1�d᫦�2`��yy�ћ�w�H�nC�`m�mh������I�Ց�v��Np��o��9yQ�}8���gwwv����4��˔��4��1��/���)Ξ�ʭ��$��6�e�v�ꥂd�c7+ �u��}����}+/�SUj���"bb�2������c4���J����8�Ғ�j���a������Μ��ߔ��d6�x�xQ��z����������o��q��*��e�[{��cl��/�N���7�k" �[A��� �O����C��zi��m��"���G7�M�m��kj�ʛշ��z{nr#��Ǜ�����'��྘�&�&��������_L����&���Zza�a�*ߡ����Շtnh%|�����v�WDs�8�Ks�#�v������3fu���
9ڱ��f�ƍR�����5��IVl���t�U��0+����8�:�촊��KK��`�ҙ�F5%f�&`��s����M�������� 5«��[Mvs��,n�U�˶2����u�>b���Y];2�.��Z��z22�⬊�˯:@�=�1���.�H�oE(ET
k̶���F	Q��_��ݹ�ey�6܇ŰR�P��܇�W�v�����:Wãbj��W�\y�M��ͱt���ܯ3/����rk5����C�J+�E�!�ʖ�S�k$I�""`�)D���5���o�w�ܞ�ۜ�
�{C�:��R˛m��|����_���4�/���е+�)w9o#����w���x�k\���zb���w+=�X#w�dEw�k�|����Amϙ«r�(��w)쳱���2�O��h|�4�:�0�r����;wâ�7nw�QQH�qV�����z˚®�����y
�6����7������s��'��s �lTGv\Tt�X`�Z�g)Glz���!�bz���r�̾ճNr��؎[���6�ja�^x�rݴ7�}]�U��\�	��q��Ng;g/p��m�~�����b�G�x~A.���a�ϒ�"�	87�I�5�:(�\
�`��/f��H�k7����w�_�ս��n���z�u�,&�O�2'�K�k׸�@%5��5'�Ȋ�0�#^�+��~�j~�x3�G��͞�@�ּ���N�3����d��b�0f-����p��|��óu�LY����}�:�{���q�����6��M�9�թ�Ċ3�ܽѓq�m{����06-�e!�.�^�a[�S����s�k m��;����;��:f�+��Lk��n�㷰��a�T�3w��{Ƿ��C^�	��UA���������<X+�������{��vݞ�e��_�v�{�4_?{μ8|;�v,d��D���4��{�[�ۏŀ��y�����<�����av�v��T4[Q�q�W8t���ؘ��)0̾�g=����hoQ�������@�ͤf���wޫ��D�)�*{iz���Orf��ܜ��i��	�O+�#�Ϗ��{Q͇X/�:�	O�`�b�U��,��AJ`�I oLa�w~�bII"t�hw	˰v�8�{!�
��n�4>O9��r�`�O`ۜ9�sh�
�l�O�%	Ts���y�Hr|�O%)//JfYؚ�1)$�P逍��|�I�0^Yo;�(�!ʍ� �mݠ+����Hk%1I�v�)�ݤ
Nn�\���+b����vN�5�EګA��s�4��8�vƼ�/*��&�������4<�x��;'$��A\��v�$��"��v܃�QO t7lk���M!@v��s�(�t�9�r(���ʆ��j(";j�&���yi��d����	�C�)=t�}z���Q��y
�o��m3�"��Z+#ͣ�.緕������5M�A_V7*��HQ�c�3H��u[��l�N��n n����d�[��A@n"4G�A����%E��i�1\���=��M�<�����y�Nh����";��(���X�Z�teT��~��z��C<�Kb��u�L�$SS+�(�Ѩ�'o�/gzO�\�fP]�MA�a��j��(�w���(z�,�K8��},7壡�3�\�xU}����C�"�&�#Q�5�j���}eLI���Nf����������Yg�����`�%˿�&}>�J�������;7EV�s�lQ0;���<�Q"�?>�v�^�zA}��"d��=��j���y٘�y�B�3�66ozouz϶f$�Nu*��2�+��m��?�1$U:w]��IO�7����zc.w,�c٫L���'��}��l�������%������>D��TU�����C<��Rܹ��i�w|����I�����U�����Zd���W�>�!@E�I1�KK���1ZJC�%Τ
�\31����Yf��@KcKcf`^e5�6��er���!��:Z�XY��ݦ�nf��\vƨC(E��P1vQ�Ĥ�7f��f�1���X:�0�1U�[�`͠�)����^�k�� D�Bc[	\�	��t؅	Y�s��29�I�����+���9d��N�)�sD�;��GuN��6f�Y�۰��p�S3�$&��L�H��p�ۜ����!D\p���@��Ϧ�Tl����u���u��b��+���!+��%�%�7�PmB6�,��^�.פ�(��U�Qe��׿��*G�)̔��^v�+��QKH�%o��$�����;�:�\;j���)B�L�2z���Q��+rX�wY�vcQ�t7A63��	��[����?���ݡU�r�̿��fr��By,������>@��݋�0gi�y���zH�R@���Ȁ�5ؙ�9]{p��d.��n�Y�� 3��'�D�+f��؉��U���2�N���;��T����(
""`������_�91[��mL��}o�FL������t=��휥�ơ��P��޷�"��
.2��!w:�\&W�V�G�տ����8f$�%qŢ�����K��?4���N!�}u�VqI(�f"�-���	���������y�	:fP��dUB)L��7x7;a���1P5 �tϢG�1%�5������B�	�J�Ȏĺ��!w��	�5����\��	���ܨB�31TL��d	�$ɋ��Yܯ3/��Γ��1hL��]�9���P/h����w���2E̗g]���J�S�!��<��/���O�ķ�����Y��O��S�[ܳ3/��?(F���dN�H�2K���~V��C�1�х2s��V\���Cmő[��+?=�	"eL�P�(�[���b���$]�����k�x�,G3VjHj�8N'RhѶ�ۜ�Zm�W/���S1�ͻ˝��ȏws���]��ʓ3*�Y;uv_w+���$i����m2�*��)	�3>�]�˿�������!n��bZ�x�-��9��=m�ߏ�8�ؗ�������K 9�8��bJ�\��N�=��m�/�C�KW�N�I��6ej�푂2;z9P��o�S�g4��g0�^�1Z!�럂�u1(���:�e-׵�
��
BQҴ�C �-*i�+���5�����ؐ�A����kb\�Y�m��0�:��L8���뵺�J��e��P��6\��u.�2��1U8КQݦb���h�<W9j�m�3�|�O���ݪ
e�9�*�p���D!i ����C��{�����y/�\Zܷ1&'2�:���w]��O�p�ʰ� �o3���1$qb���o���Z��w�}'�D���#���j��"f��,�Y����:fBI�L���&d�I�c��\vr}X��&P�C�/8��A���>�=|��Z����(�1�6�k5Q%-��s��>�bG��*��7yW�z�}$L��{|R�8�ޯ^j�:���׺o�������փ0v 	Di�Τ򑓻:��T�K��]~_Y��\W���;9����Vb\	3(JQx�7o�4ud�u�?�j��m�ؒ)!���3���"����7yW�v�\c©z���ezd�K1ݬ�·�s�����gbw}	% Ԙ�eq-��u]0��s1��Å%��O����!��KW��V)=�K�Hi�31$J-v>J4ɽz}��Yk�߿]�)���@��P��7� �͇Ǐ�g�cer��8�دO8������5's�U�_�R��SA	u؆K�4�PW�I8{��«N�s�����A$�L�� ���?U��?�j��%����"e�j$��v����?>~����yWޓ�e21��O.�+D�AC9�Y_�bx�[�Wu��jRRLA�����ə������9���y��v�3(I#�j%sc�n��m�d�L����ۛ��J#}��8[^m5ã:��o:�~��z_ئ�m�~��,]��>mz��,���g3�duf��?��y�g��dk7��]@j��!d��tݶ�UG�6�T�I�V�$E�2)�����~���Z�*�����7>�ʷۆ���2�~��H��CP5ņ��Q��us��T�11�����>n^9�q��+ʽv{jg��`g56��w7|�"���1mU��s�����s{=�+�2��|��˰j"B\�f���u�2�Ze���F�����O���߻oK�#�uųn.�כdi[��׶����kf��b���>K/�]�h��&�R��P�	�"���{}�׹�>�N������ؒ����z�����)*=2����j���Rx��c����z���V����� ;3�<�<�є!#���74w���}���j>���Cov�����뛂�s�馇��lץ�GݱO��n�{��.�=�W[m�]ϼ�ʷ�kj"���L�NZn�]�5R�Z�
��<�3zn��xgvqF7O#Yx����:W3���x9�na���{���g�u�*-.�x�6�αS��yzBb��M;��˙O�T=���3˨����ѩ��Xtw)S��" ��+�l��-������d]��;u�pIwF/:tK��]�{�A��A;^��3���uS=rA}83\��:y��"��9�z�G{��I�;�����t�{�����q�8k �=s}<;�eM���z����A�س�E}���xzx��v�M���kAN��`ռ�*���(�C{��/%�_q�n{��^[�ɽCJ�N��!N,�T����	����@X�Jr�;������BR�Gȭv5����Q�켜�h,���I))�L@u�\u&���< �6BR�g�qm�XB-w"����5�v��P�guHV�BO���4�h<�;�K�4�����'�ЃɮBy]ƈ���F�G�"���s��r{	4�Bi�[j���;c�wC��;��P8���14��� �)��C�v��6ն5T5�AIݎ^n�F�
J���7"퐣l�2m�sh��4<���� ��α�n�����	�|�|z�
gJ��Z6ݰ�`�
�e�熖ykƀ�]��k4#0v��2�-�v�XL����֫�H	h�R�Z�&k�z�B�a
ٮ��@�,Wmj�b7]� �
dLQq5vWe�ذtB8d�Ͷt5�4�͡�6,ٴι,nh�h�n�;k�z]h��B��i�@M��aYm@�Q)6��,^���F4�C:Uֽ�)��^��W�+�K]�R+
7:�5��!V/��V+�������rQ�XL /]w���R0a9K��W� ꘥�y��b���%�ά�E�rxivݣ��{m�pS8j�V��Aa�X�+��;L��7bӚp�Ш�t�^��^�Č�[�2%�лM(�����meWEh��&"�K��v�`]yGM.uc.��`��V;a�&H�Љ)bɕ-���լ�e��Yc���V�D�P���k��i�\�v�F�V*�Qcu����p[T���Wb���긶��ľd��Rj!6n�K�ŷ��܎�����XW�)Jn6*���L쮶kQ�� � ^-�#n�&�l�ef�Q��mi�)�#.%2��U3y3j�Gi�Ic�)���A5��j���VM���Wl�U��9]�rB����;9sL�2��X�l�s���kEi5�A2,)t�65�5L�[��W�N���y㇀�,̈́QdpcK6��.�E�cWWd�ikwh@�"�;�&i�-��*�b\��Bl��fi��[`�L$�u�ՙ�Dm#���kAK��0�=�Ǝ��r������ҽjK3+�e�*�ȵ�S[��)�=���%aV���%u�u�Ҫ�s"13S����"�/~ſ}���D���VD��ڌ���m�d뵂r���S�2n��#7�^U���>o6���@�̼A���x3u�x����r{�16�!�&DAsKkͬ��]���n���%XCuk���)A��3��{.�mk��1��k#7�<��M-���v�y$���"��hͮe�`�Gg�*�����2����<��n��坭mn��sj:�v�+��k��4�vq��8��������^��˙���n��/�C�`>������޹��S�݉���xLW�K��o�߷�M�p*����qh{Mn�-�!�n�l���;���������s;j#v�6����U��Ҷ�x8�ݛ�m6ᲒVj���܍��w&Uۀ�ow��1��ؗ�$�Ũ$}�3RX�d�8b�"P�Gk��y�~��r�˱W�q�gr����NN%gԼ�d7#3����{��J��� �@�Ȯɮ��	��k�|$�[^g��L]Uw01,U�AȞ誥���W�s��o����b2��p {85�{��8��7��M�G�-� ��^m�EL�Z�����8@f)^�gVߞ������-��Q`�YygW��wD��������ߎ.y�
Aa�*H)�u�9����`x�:2RA�C��t%'߹9	BT�ɆRA@���0/�_ì�[�km�B��V�@�թ0���Uk�Xʭ�_�I�:~{�|J���%	BQ��Д%C9�Y�����I����y�y�z���a���@����sN7Ņ^�hJ����J���BP��=�'a(JC�O���C�(����Xsoy^s��9
A`i���P2��@��<�6kw�5�����A�� �2�AlHhJ7��J��rr��������͓���I��RAO�����?_2r��;��%	BQ���+�{�N�Q=;�J��]�Nwu���0<i����R{�(JO�rr��=����(=���%'����E!�q��~Z��@񤂐R
]��K�����t�BR����{�[�s��y��B���)�R��<	�BwB��B���L��5����*�V���2�������X��m\z�4ûѓ_� ��G�>�%`8s	BV�߹;	BR�BP�C��	BRp��B� ��2oZ��Si���0,gc�{�=t�w�$�[�P���Д%	G�BP�����zá(3&�hJO;�y���<}YK��<�
��YIt��X��x����_}):Ē��	I��N@|#BR}愡(��@����ZC9�] �z��w�+�9� ��d���km��1o6M&�Д%'�����J��mK��J�`4�Д����a���R�[
H(㹭��z��8�Rr�d��X�R�~sv�9��^C)0�P�AH,3���
A`\ݬ��H)�U������J�>d�% 4���%	BQ����JO}��J�iv���JF�`4��3�Ǉ/U��ֹ���w�$�B�!Hy�	_�	G�	Ot����t�BR�BRrM	G�Y$M�z��c3L9���
A`y�(J�����ܜ�)�=w�����Ng�m��RβRAB�Re��JH,;}_�y��8�[���(4��j^3�(>@hJ��pyv��=ڄ�HhJ0{��%<e�{�NA�w~};�8M$�����ֻ�w�x��א�%A� �%	I�9�4%!���	Hq�%�s�J��^G� ���GmC;ۜpUMT������e�.�k�
���n�}���0�p�B�����72e/�DD�K�dch�Z���
���ݥ����B�&x���%˒��#�./dpq�V-��G�l3J�i��4+�gG-�hq�����Y��!{�#5
������hf�mG���Z�e�h��-3�ja�׮�_�B}��U�tbE�1�<���s��v���������]	A�����p�BR{�'!({��j��(�09�/���;�XߖH,1ʅ�
C�����JAH)4j��AHR}���y��=ڄ�(J=����)=�' :�)�{��֔��R
a6�
Aa�T,�R���y޾W�9����K:�I�`4%	IϿ8�����f�d���8�H(JM�S�H��<�۰�&�v�+�����9	BR{�NA�����P��f��.O���s�Y���Hp��:O}��Ƅ�7�r��8Z�`8s	BR{�NBIt
`f�H)�:yra.�H�%'�����=�H}ڗ����@��kx��|��}����P�AHt���� ���5�9���] ��B� ���(���BQ����%'����RA`f�H) �P-�i�/~�d��B�T.�S�y~w��s�3�$?[S��BP�{������'!({��j��9=�������9�M�M�̄��j��Ü�l�G5Z�;}JO�`�v��>�BP�%����ܜ��t%��j ���y�yn��w|��AL!�,�Y9���7���B�JH,
լ�)Z�`9�%	X��rv��Cݩ�.��(�BP�|)a�&l���;9r�,D�j�n?R��T��(�Y��{����}Ӏ9�7~k\�[�s�k� @�;$������̤��S���w��y�F���BRw�NBP���P���ЊV�$X)�sP��wf���?��d�5	BP�|����Ӥ��NBP��Oy���d��@����Z�g5��^��6���sj�z�=l*���P�:=��r	I��NBP���P�%	G�C�Д�����C[\yF1�JAv�����Ȕ�I��' �:�I�5	P�[�������H)�:��%��B� �7��޷}�H)!G�Na(J�{���u���BP�%�h:á)1％�
A`f�d�W����SI ��)��c�3����ͷ�$�F�
��j��(���Ja��,���P��mJAa�s�/������L��ꮛb��[���ZL���u�W�O���'� �%.gI����Ƅ�=ڄ�9hJ=�Д%r}��J:gn��]���^g�m��RβRAC�k\ޗ�Y�	d�!t��XkU$z��?[P�%�4{�(JO}��v��=ڄ�2N���|���w�0�Yђ�oʅ�
A`yT��o~y���w��7�a �����)=�' :Ƅ�7�9$��
e�ŭ����4l����rr��Hy�<%Д�h8C�)=�'!(JC�K&��R
e��V�K���ɏ�snn�ު���V�w3a��ٛ�B2![�X�R�3�(�#[�Q	�*�I	�k'5���U�VH,1�M�
B��j�HhJ7�!)�O}��;��Ğ�P�%	FP���'��l����Z�d%$)}�(J����0�%`C9�] ��w����^k�m��R�R
AL RAH,/}��gU�Ch�?�!�j��(�HvД�����'vCݨJ���h$Y��g5!��ϘJΉ����R�X\��y~�����H)�?pr�N��rr��?6�(J�`4%	^��;	G��}=��g�{��<�#���s5e%�l�yïA sI�h�s��O�ͩ��BP�~@h8á)?_�9	C�4��R�	BQ�`s�ٞy�wV���r��t���X�;�����*���`RAJ�d�<�I��NBP���P��2hJ=�Д��'���HД����Vջ�8�H)��D���B�3Ǟw��1�k�6��g�BP�{�����ߜN����RɊ������Y�%�
A��!�Д��0t�	BRv�+��`4%<�I�9D��P��)�k�c�v���[[��o���0�StB���L3�� :F��?6�)Z�`9�%	Z}��J:�iv��2�
�q���M% RAH,-����)�R�:�ѣ�!o9������U�� ���H)���G�#���HB��+����&j:�q#(�!/��	5~�(���q��hV;�橾1{�sY��c� @ߠ0�Y�]'�|��J��|�(J�`�!)q:O}��Ƅ�3T���S(����z�%��ż����o_�v�H�,�FZ!3I����_>|��B���誑�͙���Ȳ�\�j����h��ͩ!�/v��N�wd��=�!F:&�_r�,��x��AdYDTH�;z�����!�	Ҳ.�uv�*��5�	g�uy�؅Z�"�F�A�"^-���<i����v�HYD�YP!�۽�Tk��O� sW����wN��d��'�+�}�,F��}V��`��An Y3wjb��y<����Ui,�u[Q��h��т����(jvk�b�nkmFTe�jfೳۖkq�mu�jwD�!��5�e� ��ʷچ�ڛ-�
���Hk,�]3�Z�![q��it��h:��6d�I�HR����2���f�ZfmLR�zm�Z�&xu�ɂ�𕙍�0�؏�ڃ	@�h\��݊i��Tlh!��i��XR��,b��%�3hWYc�}����t6�AN`[�uB0*-f�]��%�XC�@#�!����[�o_q۽#�ʒS;i(u�2v�f�� c�������Xէ��+ZE�!�}�;�ݒ�D���^�KȆ#�s�Q��F<Chd3��m-���Y[3�����-2�-�AdGa�T�W��"ϐn<���S��nƞ �P"(ѷ�wEL8��%a�h@a��[W��އ�!���ܗ�'�%�D"!���|����Ը��e�A�V��S<�X��7��K��>���D��8�/��:UE����+רؙ����m) ��d"��%��!W@�x�j��4J�Ȥ�CY�	����hXR%����.�tv�������� ��%/�ط����;w�p>g��Y�Z����0P#2 l�Z�Z��VL�֒+���N�K��ڂ//ח�p @�* _c�G NǴ� �V�wf��L8��<ϑ� ��k_�VGȆ����|�giʪ՞ڈ�wmT�i۽ w�>Wp �>d��
,Fk�L� #0�B*�Q��9#��e]��0f"d��=��L�ו�n�����$�ۅ�45����"��n@E�EDL������# >�Kws{#�\	} �|�:��ٺ+1V`�j�"��5�}$4�A{�;ӁA���������㦳���u9&������c��`�c>�wy��i�" �X����5Xs���/����9^�{e>,[h-��Wx��h��J��3�G'����ػsO��X��Y��M���^��"�ޞ�Z'�׎x�^l�ߝO��@~���u�z��o÷��D[���{پ"7�?7�;��KG�ў�kgl\����;ݓwV�l��>/����Z��7�.��v��]�,�B��I��/���o���ښ�ԦI�̹�3�&�f�=>��v��FF��|��Cغ� 63��{�7O��q�}�w_:�����}$�έ�ݜ��7�`��������ͳh����}��"������^��x��oW��� ���_{|%yp�^+���&�v�N��w��S��\���犦�U┖��6w{�|��8�η��_����>:���Y�3��*�l�-]l��L@HM�ٲ��E�}��;��c)�g��ih�PQ͸sp���"����I��Ӣ������Ic4:OnA݀�_6��[U��)i
R���4b
��y�̇�"��)J*�y��%5�4�jJ��
$*&�;h�b];c2�ڶh44Pl`��伐��Z�����伀�UEEHP���I��M �PX�#%!^�B@/�W;�����k��E�H�Z�g	L�I�X�gM@A
!���k�Wڲ���VH�[P�ƚh�xe��Y�Y�n<�utD�'��e_F̸��@%� F����q��|w��}V�z��*ۜ�.s퉗v�`R��&Tk38(�5��^-����z�N���ܛ��I�Ck�|d6�|����(uP$ݯ3��U}�rH�����CF�&}v� #EBd ��v*v�j7���ٗ"Z��� ��σhl����Y��8���������Vv���8�Y@�����u����̘�c��j�n�J������nD6�ɥQz�zV�`���� ���N�xʏZ��a)0�b��w��!F�Yq�ϲH���h"A����蚜����`�!cs�t��6X�KZ;\�@gAHdK+b�k{�L���@�q���P�A� ��6���(��6��{k��Eoq۽#��@���ș�y3��ht�>@���C^�)�����w"x Kj>��ix��Y��'"4#2���������.*�8|���*sŌ�(�Q��/6�σ���Ќ	��@����Y�6�H�	g�hH,�|�ȄZ�&�S�����m��Zdh���5m\31꓂l������6vT���y�v/{f��+�xx���P4)���s�1��)i�`2\�����.�4Y[1
X3�[��`��@z��`a44&��]�Eq��=�;y*,!/�
+	��Z�1X:��`ɺ@Q�7��
��mXb�F�9��%s�j#Z�M2�\�v4u����_�b�ٹ�aFQnt��s���TL��3���l�uy�$��V�����r'��7��e�PF�}���G̢�C&�������=�á����,�4�[V�,�u�Y�0��Mz�p�p0�>�*"{���'�K�GAe������� �)_(!�]E������������5�~�)�dI|������`�ޛ����T	hqg�Ax��ϭQoې� �aD1@�� ±�e��B֭f�]��� |v����������:��zG�v�Q�jp��(��<ϐ"}�����j͟)�M�ī����n��������iX|��� ��~�`$���=����ע����Y�������j�tz����:B ��D���3w�á�*ﱽ��@���>DAי�dO��C��|$��()ʸް��eV�Y��+�R��74!�6��σ"<[I�{�t,��oMf����t'��PF�"^>n<�z_������{1gˠl�Uչ��@�,�b�ol틕����}��� ���wx�7_����Wş#�w�Z�!�����w˲��ax���6;�U�p۽#��� ���o�}ۺ >5�Ԃ@5"����}G�HÀ�'�{I�e�F�30�����e�}q���3=y9�ʫ��3�R؊�{����������I�}����ḱ
��ܬg4���i|�.�����@���|�
�4shY�^����k��A�L-�л��u�6�HYD�Ym��uݓ�DϠ���p��A)P�a�u\�c�O�Y�N�;Ք�ˡ/Y�V�͞�wBH����13v���ȊAx�!3罰A�/���;�ܡ����"4�[UB�ؓ���	�PAyϐ��GtJ�J6��=�zG3�+ Ag��!�����䏯�A�A�r��]��殄���PB� ��P_E��Ƴ�&�W�:Q���1���o�w�-�iJFg����{���U���� ���#^9q�D�2�>nF֝�t�,�2��f����-zO���ͩ!�i�UEV�?g��l�(F3J)�\�]��Qk�q��>{���ˈyz��/���w���v4��\l_v�H I���@��Mej�n�3d!�Y�wuu�]	�/6�N��(�n|�"� �(�ЀC 3}�=9[��6����Aڀ|�Qы���Н^Ӥ",�y��#6���U��O��ɋ�}~dI�DK�@ �����ΛN�zU�i���5t'��PA��h/�	�q|*C��lE�U���/]�`?�%�-7S���D�O\r�)�9�7��8�����<>�Goa�mP6�l.^9��h6�Ҋ:g`%F,/S::Z�i��U]�� �,�.�d�%��M*���A�(�mq]M�Glh7]��(i�!q5g!+��Y�1R��Q,Ф�.�\ҵ9��F+��]�W*��ֶ��-}�>��
��.eVc[��m����@�I`T�r�'��!<�����!gU����N]@o���X�j��&�/�5��@���M�1��R���|�����ڭ>}��$N��w�>�d=�@>6|�-[^���M�l�i뚺G-z� CAx� n�5t�uwJ>���"||�tt�n�'.�6�ϗ��j�C�2}�5��^m@ ��5\c�}M5���n��ڭ#� ��dI�6���L�W1/�ɉ!kc��cK��8���(�D)�Hh6|4���漆�eh���N�O ZRX���)�� CAx�d A�aa���3�;0��r6	�5c������4�N&�#C�a�%���M{&�[�ewO�xxz�C8@G
};U��A�u��G�}�T���*e�>�F�� �|�g͡g��m'�g���o��q��n<�YD72���1j�C^^Ȯ���zꮄ�^�����ʯ�^d,��>M���h6m�4PΝ��ރ0�}gȌ>mzZ��
��N���AQ&$^�G�C0�hJ���9��]��%'��z9yϓp �5���OH�+�Ҵ��6,�&1E��P�V���أ�W�E]^���Ut'���F� n��.��� �D�AdY���&��ʭA���T��w�sF�G��Wx��Y�N�s����=%s�����N�^�׼=�J����1U��ς�mz^@�B�LL�Ȼ^�^}��W>��k8m;#�%��7rz��$+ G�>m>@���"�
����X,��nf��Ut$�Z��H!�&�g	�мQ<`��0"Q�QW*�l`�ΙvJɳ�.���4|x�FR�"O�Y�����LU@o�-Z��Dn^�"�j��dAmApxm�Q��U[ޙ���m�A,�dy�{T##�ذ�j��h"ڀC>�Pu1��OY�;�WByzZ�j�4�n�@��.��I�L8|���ۼ��Tפ�������;/����wU"{���l��&Q���vTȫ����]ֱ��C��^@�|��>d6y��ץ\{]��>w��m��g�ݐ �,���C�k��$p8r*,�kZfYT�6R�ar�������W����yu/75j캺�f%p���}�ȋEFc,8J��j%�6�[x�s)��J���ۼ��T��|�b����*��BZ��@���y��hs�������Ѯ�8m�#�%�^�%�e�+�R"ϙ׭� �}����v]]	���.`f�=sK�����e[� �%K��,aEMMm^o%1U_z<ϑ|ڐC>c�]�㮙f�8p��X����ɯ��v���%)���z�l<��H;��[ZLV(�%��:�p�)D�O��J��k<7%���U��N��b_=��R[ݑ���ҮEw��W
�+�X��\�ji{�S���p�m���K���V`l����m�s�������d쯘�%�d��_���1�N�݀�}zeo��flī��҇��փm��u�gx�O��z�+$�_bYƕ��y��'�{,�;�R��;�����s����i��\:���.yz�U�y��Ȫ7=�u� ���h�N^��n�����;o2���7=���_��{�)Pv�'gY��_'ۂ��a�;6����&�F���»F^�ђ!nX'�Ȼs��-�t�ب�7'*;r���Nr��[��������HE���t�o�˔�~#A��-Xc����ܳĭ>�[�Wq��j��Z=<�V�ϰlD�2L��x��S�T�Lw��z��2&!��x}%�]NŽ�n]�@�&^A���!*!�#��g�Q'#K��Ur֒"fms8�bߘ��R΄յݎm�ꪝQ�"��G#�0�K��4�TLhvأ�#N����F���"�֩H����]�Rw`��6�E%.�DT�kDQ^lPyj퀈��PSDT�T[���"*f"m�Z*�()��������#������X�݅�nˮ�a�5�\)h�S:�J��ĵ+�X�΁-�lm�J���K.�.X���"#,���3\�p-n�]6%Ηf�T�-[���
�Љ
K3J�5�\�ڎ�6�p�<�C��Z���T&����E�cD���]���wm3���6D�,aɡ��:fimݩ/&4Sc�etF`�61�VSZP���04��ssykk��63~���'�2�RX�2��^�M6뵪lD�G1�A�,hVh
5I.F*,�#S�h5�jR�e��hPl�#,��%v�� T�̻6�nN]@�m��ɡD�AԹ!X��]*it�t�#t�í���Z�[�K�Y�a�����J�,Km�&&qv��ɺ:�m��P�kVn 1�Lmm�!�A�͛�4�b��Z�TI���-�78.� �s�(���v�W]�
`��k��!�k��.�hnvt�أ�eS�Z�P��6�*M]0$6%�ݘgX�KH�F�h���3�G��Z�@к��,�����b���{�����D��`�جFԲ����-L��c�ԣhepM���..6�I�5f��D�kX��$�r=MpU����<��+r���U�W!Xʪ�c��[��/U�F�.��i&�ڃ���JƁ� �θ�h�¦6	�Hy�<�*����� Z͕�`�mJk����SEB#�H���.�(gKtYp�6���:��֠�iKa�kS8f�/Pd�c\\M�b% �g�g@.�#�l��cc�\!���!Q6��Ń�W*�7͍�mv������.�%��e�a�s�s��z��QJL�
� A�^���g͡>7���p�t@��jnaG�#��",���y�/�k���E�*>��5���v]]	�%�^D;ۙБ�zr=�	�Anx�>g�u,ۚ��Ԧ*�K�ş"0�[PAkȆ���={O�[�6�����n�k���p�tGK>����`=��4���BAg�y��j��e�>�9���lve]	���F� C>mD�Z��TɈ�!D�0�#��1lci�2���;\�#A>[Q�D�	f�>��*�K�C�-;>�/� ��i[^y(̋�����i���̈́�x��"�tmN���a��=	�Qۮ���	�C}����uz���okaw�5��#x��=����|%��k��ݻW��\��̫�$qmG�:��ЀYvI1g�w�����ϳy)���<���y�'2s�)�|ב Kj-y�-�!qyr�{2��dp �Q_tǇO�ؘ��Y�b�q�W)�5��3k�"&�SB�6S6�l���Ԑ϶�s�Nt�UОL�R�R8��myx�Ax�d	�F1�B�1��l�a�3e�n�1U_z�"/6�A���}DR@�Mz<׃�/���h�/�ә�܆�R�і���N��t ��v�=Szx���I���	�B�Ƚ�{��|�wr����K>�BAd",�ChC���T}$3��}����ΜʺG׵��՗f��� �,�n���t(A�����SP%�y� F6���snV��A�AQd�	���7��C��i�aqI]-"fHX�=K����4��}m}}�k����3�ݽ�Z����@�ϛ��>@�f�)�k�U=��:s*�O��NT�1k�p�:͋GIB.�Qw�'4�[}U�js&�9�U��Y��ͯ3�,/u����H ��Q�n z:�_vR᭲8�(��Vs5D�Uէ/�7�o�F��q��,���%X�NHR�1�o4gNKNDq�3�r��3�&북1�X\2�A��kh8Z�>�7u[�7�̬�$qmA|�gɸ�)��Rz�p&ѳ��fr�;&ڦB����b� �"
���#���A}d A,��}����@o�+�]38}DA���gͩ#8m@�{7��>�q�[{Qݔ�kl�̢3��t�V���>���� �-�3��uod^gW�̬�<%� ��Ȇ��Bd".��n�D/24K+b�gf��5P��>�Q��Lȿ��k���j-yݽ���n`A���[�K��τ�pΏ2��~�����iJ]b�6~/����<@�G&՗��ɷ��~[�Q� ��ށ�SQ�W�͗uœ����;	(��Ζ4kPm���B?�ǋ�O#b^&5���5	LVaU�1\h�K���+v������ŀGCK���]3�-��I@If���Hm���pۘ͹�ئ8�A��Y�.�`�C3M\�B��a�W9�PqD8X��ߟ@ߡ�%�� ԔT�^β�]eV��30�:|�B�mA�]S����"+87t�-x8^m,��(���Oj�d-7�4B���ml��U�8��A�-�¢5�]��'�$#T�yח�BG�CW�϶����ʭ��N""��Z].�DK��5�[����<�v�-y�}��{U�g�+�bm	�O�<&<�:�Ȓ,�p C�D�O��cͬ��j�6�'�O�W�5젻6�f =�P$Dʕ��Ǌ)�s���"�c�R�e}τ�k��5�CK��A���;}G����]��5E���D�3��<ϐ"�hu���țZ(�ܿF�>�ҏ�Y@��F������pvNh6�A�CE�mA���{���ڂ,����n<�a�������Y�uig�L{�	e[�2$�YQ��d��.�7$����y�"8���|�dA����@ �����B
�ܾW�xe6GK(��u�Oq2T�d"	���,�A�Κ}�*0^�n��w�wV���״�6�8�4%�2��iXu!��Vh$Z/7���-c),
���_D�>��$�,��y���*�| cwYz"�i>}�z�^@�B-�!1\�f��M��w�\����l� �QgG����p�3",�^mI5�����[�b�;fn��z���*+����=���NI�1ko�y�JiN�E�w�77I�W� Wk�ὓul?����j�4�Bd#M�V������s����U��|Y�#Ui�qp,Q�PAk�ϛR-y��j�(��ǌ�����*�%�A� ������ߟ>z�~Ma/�p8瘳T��ar��Dm�®.��>����Z��mz�TV_p�ɺ�䷯�Hy�|F ����,�F�'�& e^>e��svzaU@mzO��"�F�1ò������� �|�hU�Tq�f�Wi7Tτ�g! ��%��/w#��CA� �א�����7V�� Kj��gZ�qWO��3�D_���B����h��@�L,�y/4���*`�yb2pj��1p��<w��z�y�'̢p ��Ƀ�>�`�3[��c�b��<ϑ�@��Z�l��Lds��"B�0;�Yh?�<͏^l�d(,��TL�B�҂4�8^mx�﫮�����8�f�b���zt�=�e��>�Tf�O�T� ��ʚ���їV��ŵ������DG��>��"A�.i&��{����A��K>�E�׃�#�v��T�����)�m�V�n�� �Y^ �-R#ƈ@�h�Cp#��&��2g����$��1�gq軫byk�}$4�p4;ݞo8��V�E�kQz,k����<�NO����������Y"c{��'7hM����~�zk�%
JP����>�-cV�4@�[��k���b\3�Fkv�cf����
�C.Pnn�s��)1-#2�M�6�� �]�L�%����j
`nn�$�a���4W5�X�=\�Y���#3�r���Ͷ����_�i�Ļ�Ţ�!�K����[cfX2�%�ع_�O��>O�@,��d���ݍ����W���'�2�zڟZ�gͦ�5|��ix���u{U�u�-���Y�΁���$ p������6���:���FWv����$�e{��^-Ǚ����FF�w�o�s^�$��6.��v_�A��>\�'��P#��iy��t=Q���ޭ꾺�V� �G�A,�iEj��T��"D�d#ՙ�1m�iq�d�b�VDfbP�^����[^���EV^wr����wa��R���Ȍ^^m,��L����*������H_�z�u@�R2��N��%̅f��V6Ɲ=�BU �<���Z>�Dx�����5�R��K>@�!�E;ۚ�*݅kȈHf�Z�4�AM��|z�h�ɪ�˽n�>e��B �|���r��^�'� ��Z�Z�*����ut'�%� �N��Q^M��ϐ͏2'���An<ȋ��H�t����|R��|�:�ڒ�!N#����}����p��E6���@z��]Kq��>{���О�g�����]�ݾ�uWDqj��ú B�~ �@�σ0Cq ���!m�F��Z���ڢ�ŵ^@��Q�@�� �x��m�� ���z�5q۵u�ż�bv
5��@ɺ1��0�XJ����{Ǹ����]+h��C�$��9�On?�'�ݛ�ս���r�4����f��\,__"}Ǻ{<����k6E�n�o�^�Ez�7F�丹YK���Ո���^_L�@�x2�f��#��N��e�
H^�c#��;Y�!�r��+:o�~Y��.�����h��.����l�˄������C�%��²����4*N�+fk3u��v��������̇����o��X��r�o�����Jz���@��|&]�� �j���o�};������5�G��Y7�z|��w������HJgV��9��S�({0�7o�<���9�ݩi+ �)Զl������?S���eǑ%��a�K��j<��Q����E>X���si<���!+��$(>�1��*m\M�I�p�Cw�r���.�w=�^�;��\���'!�/wv���ά>ij�bEMel��6sl�I'�	'ēDE~�"���b7���5US%ITLMS]���r�LU;9f�j&���������
qECPAQLPPP�PDTCILU3%��UIITATTUUE%;j�f����U�*j�*��e�H��������9�Qh��!����51RUMUD\٥����("�(�ͨ������:޷�W���9����e	ġ�*C^����:��a�6�g^>ܾÕWD,��t��4�7�>}3p	gȂ��֓\ؐץn^���]�В;ŵ^�<�
�:��[�*�P$E��+I���(�̰4�2�I1 �B��� Y���Q�D��im]����U_q���Qͨ!� C>mIyg�� �� AN��v�a�WDw����t,�<G�j�,�*ЃG�Z��y:��7
�bv�z.n��#�j���^-��Y���U!e��A��(��쎞�]@�C�gȊ��篢����(D�ߚ��Зm�otK7`��v6<���γ;����������w9��_�^�%}�,�3��א!��S}V�0�|���Î���� ����D��5By���L�ع������\�`�`�*
�b&�3�o`g�r�k�ז�V��s������VO������B��p �,��ea�ќ�8B��ȫ=�=����� �|�B�6�h�����#P^�PgȆ��[�ګ��u��{��s�㫢82�FrY�������A�.���G)z<זEe�wu[���ep!F"�5](���e@��@�>M���u0A�^��ʖ7p�p*`M/I����^�'Z+DmDx��Iw{��dF-@���ri���<�L����&�| �f~PIHр�7��l�X���M,��/�cY���USnö����KiY�j�&�*�#�\ڦ3ؤc@5�ۛm�������y�`�����#q�T��åQM�J�)Ԯu��3n���gm��b��m������Q�s��0�ߚ�yIF�y�-t�Q3$/������CAx�kk����q��B�ux�gl��=�I�+�7�"%dGnH��@ ��������Uv���-�F���n�\ٌ�FD{p�p �,���nݝ�L	��>�A�ڒ^#I�X�* �^x�/k:�/�㻢PeX��26GX��#�+�7�|� ���j����pa���f��S꫹�@���j�!����k1�ZBT`���1&"A ı�e�VV�k�.��ت��0NA`Ad/�sb���L	heR��>�A��Q�k��ŵ�ێ�llW���w{���o�� �D��2Tr��b4��s��rW��N�dG�O��A{��)�oW�a�wDq��"���J#v{O� �m@ ���T�v��0�wW:��(��i�!��ЀY��c��c�U�֜����/� �|:D�wm����Y�PG|�`�|�k�w���_t�X���o�㻢8�Y^#9,�A,�,_v�� bȑbRA0$A"V�v#��-.�'����A�mA5��w��\�]�D�}Wb&�>��7g��%���m��P(�N�{5�8�p*`KC�>|�]}S1xA^(���7;s7�/v�~���pn՛��K�;y���&E�?wnud�8��מ �z��_ 7��]f�aǗD|A,�g@�Y�Y�h_u.�+h����w) ���Os7����+�����(M\�J��H/�dI�(��y�Ν�g��_��1}�Wv����>�q[Pg�v*_�Ϗh����=In��[�XA�-е3�'�V�ˈJ^��O+sko��e�E�}��zjvNc @8B>e� ���A{�*���ʲ��뉬���Wt+����|�g�0m�]T6�<�@��@�ϐn��ZP����Uuj�����K>bŵ�kȆE��]�����͠K��՗�r������#gb��ې�Z�:H�xN�`�sMf��E
�puh���s}�P %7���"��Gx�6�ϙ�j.6�n�	y�����uwB��W����hg8=�E��tq��+�M3gZ�e(�K`A��/�{;���{�D����ūw�S_G�n�wO��N/[^%��̽�^�- �MJ����wDq�(3��rttг��(I ��L���rN�8������\�mAW���[�2$������+�@��U�عf�*`KC�g�J����Դ,�a���E��|J�J�4	��]�ʻ��'��B "�=��y]r
\�)d��u�}�4>�禮s57`ک�[Ij��¾�-��&����G����T&���ݙn/��B�[Xf;C�E�m�i[,��Mb�&�cK��eۖF7:2�@v����QQ�����s[UT!6��u�kQ�\�J�Ɍ�ˤzC, XjM��tf��*��fn�"��ׯ�٬���k�F�wV�*�a�A`�t$���L؜C�g�{��^gܡ�vv�U]Т0�0¥02}K¡x����3ꠜ�c){�kq��T����|�B-�����)yk�j�Z�g�%�9V�fV�m輫�#��@ڄ�D���+N7�Z} �1�Ak؝wovҪ��\�׌QѫZ��#^>�  Y^!� C��ދ���.���EL
}��� ��^-�3�k7��x_aD��
Q13 �Q����8<��Obh�چZ:d���( ����x� ���ue𼻺#�c\��7gљ<YQ� ���#�;!�8�ű�G��͚d����������M07➫�쮿z'Y��� %�b�A��N��ﳨ�]Ю@�ͯi���Z��>alH@�t�7d	,��7��0[��ȩ�O�9y����m�6�P��>^#�n/���/��]���FբW3� �Nn ϑ�6�bC.���\:��}Kg6�6�U�
>�\F�"͡/�/��_s�J鉧�֋��hĨ0l&�`��-u�U��=�9P B>d�i��}ȩ�M����>�G��^g���j<GXj�ou�o��^;�"�����9�b���=� f����h�܁ 2��'̌x�+�����n�{DFk��yG�}ϰ��O�U<e����WvLɥX�� ��jҤh��1�����N�|>3h"Hgɸg��2xT���H1�� �PWVstgpJP�� ��˥1[�6�N L��,���W�25��Օ�s.�l�΁2"����h(�0�G� �4j�ڐ-��&\6���T���^-� ��^�����¦�r��m�Ӕ��2-/� ����Uj��g�pda�.vww9p��&��(��͡"�>�$���(>d CAx��H��OmNgm��Y̻{��Q�A�|��&,GI�,�^�RA�d.����|*n�W M�ES㺷��߱�gA�,�Sˣyo~	��w����4b���>ů��s�Öź���k�`�:&jTu����Fv�ג�W� %�ƻ/��"P���!�/נEq9�F-QfL�I���Kff빚�^F�*����z�gɸʬέ���v(�!�V����A��qe�@�-c��5�"}�5{�;¦�#���B!���[�� �@,�Ch@!�A,��7�*3w��(�&��D9y�$Y���5�')ҳ�!���7 ������9���xv��"E��@��!��^m.�Q"�0B�w������GM@>��y�«0��pC�4��Ȩ�pež��s��]X��ï*��} ����/�����������;r6�7N�E�Ǣr)�R�nKy����j#�xnݘ�����:�x�����iE]��@��8�5���f�M�����74�!�u�|V�o��	��ӡq`���^��cO?B{�F�&v]��)ذp���Um��v"w��.���̈;�+�����ɞ�>Pr��O�v��}(G�������!-�GܚZs����V^I��yu>�s�v��JwRS7�=�'&SUk���qA��v-��Uй{�F����x��fn�@�/�:��ۿ�����uv�կy}L�#R	�c�Ȳ����mH\)qE�x`��eUO{�GtF��U`��i����qbeo�E*���+�{@.s=��E��|0��&,�Hn��9�U�����9�swz]�
rT;�.'\��a�AV�u2!^��
q	��Х1��v�(�D�T�U5Q%5Ws��(�"
b�����cECl荴Ѫ5h�ETA��:$���F�)�lE��#Y���f&��ƝSEli(h�m���#���㦊�����&(��d�H�J�LD�Rh5ٞmE4S$�V�L\��*h���)���8M�UMi�UE!E[�UG`;r��t�0D4�RQEU�M-v�؂h�)����?=�\�8wN{*6q��3s�;2��3]�˖1�.�:l0eu�AĮ-��V����iNs3"il���c�eJn!���@Ea.a��4tі]��\�؃s��.����D���r=�(�)XF��KCl��9�%霣���1R�{@�+u��bc`�[6�hJ�f2��K�i��� �M��l��M���]���Eb�ַG��iB�"�.�X�(��3��bve���Bd3dtVb��^��-�f(�5R�Mqf(��h�+����f{ 5X�U�.ȸ���&����)M�љ)����&V�q1�Kli���L��գ��KbM+�h�%��Mֱ4GQx����3j�MnN�L�:�Zcumɨ4u���h����Y�[B�����p��h0W-V�3΍�]�Ĥ�[-ͳu�Zcjh�i ���93��қ�� ڰ&���W[�[RgV�-Yi)�9%�!6�Q�1J<�)�����4�W�i��p�[`����4g�����E5Vc[�uՌΎ��`�(%l֍fK��vz�ıv��͚-qsQ���p�K4!�ٝ4�4T(�b�L�U�o$+v�ָ����%STդ"]�qL�h�iZ�u1��\U��kL�\�ʰfa�UE[��Ff��ЎB��T.B�촡����anv&e1��c�aQ�jh���ߤ����C�����n�a�`�6�a5�<8�M!�G�Nb�K˦��Aƛ&!LGs��r蕁Zۦ��uȦ+Z`���"��Utttf�^%٦��hh�q�b���5HJ+4�ƺ�gs�EUs�
�j]�m���=��r�6��򚅬m�$�0r���\�� �4Q�<�Y:���b�P�C�:*j*ϸ�>�RAy�� C�0\� E!U ������y��GM#:<�]�l�)	ϐ �-���,Q�r���Sw�o5��b��i� ����^!�� 9�x�F;>�"`@HG̮�gw{W��@>4|�ѷ1ǖ+>�/6���!�D�M��z�!*�����y����>�BHeO��{�����U {���6#L,�J:&�e��t�3nr	������d A����F�w��9��b�!"bT	���ȣ���%��&4�@~/%X��Rۛ�s�ݹ5��`M�fYb���7���s:�%��S����:�hgZ��:���+­z/�,"e(B5y��^�Agً�Y�^m�W�,ީ'*�{����G� >�B|C(��n Z��QC�D��x� �-S����t����$�6#=�v@��� 3�,�A���f%é��R�=�شDI] �D5[P%�!����1��8��dvMn�c~�獌��6� \�>Io����/6�yt}Wv�
̬|�:�1���>m��,�T/��ڢ	�觹���E�G�A��q۷�7 G���p��� �W���H�]��9�c2���ױm7:l�g1a'j��K.��`�����k� X���\"$���(��j<����&c�j�&���b��;g�fV
=�}Exbc��(���@��h"�xv���g������������-�G���C>m\����ǮY�"#Rl���L�*4���X2��PT��	 Q� �R7{;��"m�����i�4�!�"@�׍�+�c#̌>Y�#�\]\f����#�A4QgG�n;��E�E�^��-[PAk�<�;3Y�=�\]1DqmAj�!�/6��@��ɩ��d��'Ŕ:����&��>Dt�|�T�2��ɖ���`L����o����x�e�{Ȝ�4S��;���r>�_���@���5��'LϮ�;є�ܝ�YDq�9��|�¡�����h>�67X�W�X���`���u������O���ͩ>d*�����.i�D!1ڐB)��(�PՂ�c-#3��kT��АE���;;Go��� a[X#.�{�}dA��r�@p��;ua�,�[�:+2�Q�}E}�e	g�ϠWESD�efנG*�ܝ�2�Dp��}u-�*��\!�A,�A���E�M���4n�I�7�"�P^-�Ade.�an�u�>��N�m��GZ���TU����Ǩ����Ġ����5�Kz���oC��O_��=;�fY��є��	(Sb!bK�DR�Skhe���]IV8�maIW2��Q�i�50�.%u�nȣ��\ٴ%J@�E"���ؖ�8�pR �ļ]
���H��b��ƛ:�Y��Z�4Ic\�*Vink�_ϟO�n���STJ�MZ�h��6��-�������,!�PD�ϛBB̚���³+"*%�}�$��T ̂,���d/=C���	�������.��MA��E�2�ʀ�B�P �>A�C>@��v	Mk��/lv�I�7�	B�"��@dc����J��,�E��[�k"�gd���G�>g����b���(@2$��E��u�dnd��N��]�t��NE�4�i���p.��73ٹ�\M��R�D\a��v(.�6j��e�]s�z=����曉�a�6��=�dM���f5�QD���@2$�B��1A[�X]��������L���*A��tr����Bbͭw��7r.���w�X8������������MZ��~�X(��3���Y[��4P#� B!��mG�%�]�*Vv���2꘣�+�:���̀��2z��>��!�P�b�4��I�7���N/����k��ŵ��ttEx�@;�ǻr8Vee8�@��#Ő�%�L܍.,6|���1r�4v�SW�Iu����ͷ9��Ͻ�z:���5�kˢ��9�uLW!�xq��Y���ļ|�y�$�!5V�П!2������tz��|ڣ���l@�j�����>k���h	Jg"rIPl���:�i��Ǫ޿�?�v�v���e�ͱzjtsNpN���_���e��#�,���@,��g�ϠI��{v|(^�R-{Uufk���G��-�t��ċ���P �Q��D��Dh]^�k{v�hJ�u��>m2���θ��0��e�#CEK?{�<�dq2�BI��!|�7K�=��p�p�o��ᗏ(�#x����6�B��D7	g�<0F樅��;�EZyy��p�4Qؼ�D�\��ئ߮.x���Ck̉ ��p�Ӻ0�2o�����y�qjס� CA���f��+ ���ix�����|�e��#�Q�.\w$��|-i�Ӵ��T�S����ppGH&��״?_L>,V�͇�YqJ�:�G�U��4|��>,�&�ڎﺨf�5�Vo>Z�T��	����ix��j*�a��
����K�mS�ɛX�9��u�]qU|���=�{�HO�x_y������T���Ȣƭ Ȓ�jH���I�j�h�f�x�Q�A,�A� �GP����F�C!�k�"�zՏ6����Q�J�A�>��}v A�g�HX"����+�x%dU �[ cy�굀��iy� �����e����\N�mvj�7����g@�D"^k=�c.�
y۽
��:jF���i�7�;������]&�}���y8�ʴc*�7����R;f���ߎ��1&�/V�G^����ZZ&�f�h�QL�[�3v���f��6�aYH$3 ���b�E�X��ܚl�)V���]n5�RQ��bT�"M+ĴFP"1څ3e����aP�@4��3M����\�Wk0�f
~|��b�����EJ1�(ܸ#�%n
�L�O��蟨C���W�J��u��5R+�dޭ�~#��n�}�;9�"��@ӽW�oo����D�/Ԫ[7(E����� ��n�N�w�.3�Wf�+�b�|YDg ��|��aO40� ��PA,��YY��q��Gj�ח���a{u!��D�@!�ݼɹ�K�ڎ�����*��B#H@����C����Ei�=�d1�WP���Ik���ZB��A	L)��da�PA4@p���'-foF*�b� �un:da�`�-�}%�n @8���v�Ŗ��̈�B"�젍�6`�ܶ*�����moQ��RqZ�cKYx{Ӄ�n���lW�����&�Ep@�m���u�N�b`@#�g͠IQ2��8��ݚ�*��E��j��@�uU��nV�^�Y /6�.��y�щ�X����E���,9�F#G�ȀA�!�6�����cK!���w��H�;��H�CAx�nr���tV��TǊ�K��ZL«)���k5@���u�Y��B�!>z�x$$</Ee�-����U�#��oz4q"@�/Ad�;j�����"Hļo B��7���U�<|ϳ��C%]-��W�(�Dk��@�כR|ȱ�_|�_����TcEگ^_�ͽ�șO�c�`S
[��Wix����%�}���k�g,�:�t�S�3��n�����5{�ۋ���0N^�H;�Ff���㏔����B>����9������S�Zy)�-F�����d��p՚Kz����z�8�s�XmJfxW��2���=��q��/+���U�/�>����*]�S���9��N��^�u�摩{� �M ���x���pT�n�$$��{C��Msv��i��mO=6��v!*�H?aָb~��D�m�J��nx{�^wR�I/m���,��<�5�{���:o��_1��VWx�c�屮w�ך��l��7��gOg`5a��Y�V�d�fq�3� m�FŸ��N����{o�{h����ؖ��O;>�77QZ N�
��"v���[n3(���4�C��F8�;+t���n���%����gn>��-�/�o^�L/ئ���	r ���{����y�ۋ�c#"/6��Ѵ��7�GAԈ$���np�15[���AM%W#CATwji�
��nmR�Ɗ
��(�֪J#��A3]�MD�1%)E'a�Oa�LEDLMRSQ1RTI�DM50S#ES��������b ����wprJ�h)("R�

K�(�Mh�!K��QBR�]·���i�nd��R�b(<�4PP '3�k�s;w9��E�U�x�-Q���C+�`���N���]@d�����=����(��n2yL	��b�	d CHڂ�d�P�a�>�-�;�G�����G�%�,�eK=_^�ߞ���B]�hL��Au#2Cl;\���nm�Ϩ���OD" �mABu���I��\�I��I���k�Q�>M����@��˪���3�p�Fޙ����] �D"�`������!)	�PA�d|�u;޵ۇ�3�"n�Q�A�fo�/�i1�X�狧x�](s2E]f�;�j�Qm�]+���M���#j)����c���[�+$�ɄBW(�sZ�RV��#�^���7_{��+�>#���5�|�l��u���Tع�{�+wޚ^����N	�I4p�Jz54��8�c�1�O<��	��H���$$����H=L�;���wF�����黺>욟�6��;��p����V��wYޓU\�����1������0�F�f3Sw�![��^�n|�SV��]��/2�5�Ƿ�vL]]����r/��6�h2�9����5�w��I�������;ǹ,�(��o���ʩ�㺮vx�蘶]�[��W7Z�-�Mm���C� ���`����yIq@��ZlLb����fSk��s��V�lP$�(� WL��-�ჇKF��l�$[��%:���ci��KH�;B�Ͳ9n�db�Ж���Dn�X'.��]6�c�Ib���e�*�ȥR5�l4S�����Lt��h�*b[�ƍq��+*�)�S

����Hx܆r����wAT�&�҆ET�dM���kO+y5&����u���w\���Fsw��0.כpt599W�gI���W��ۘ��[8����^deE���zZ�3���Buy�6�nP��פ�b�Y�ݘ�4wS����9ɷ�����DEL�Z7B`4�1oiB�+�و�A*a#�}��^mz�v�k[�]W{�gٱ�[���Ck͠l��5�����e:؄|�=t1bt������k����0��O��0��ơ��{�yj(wO�wAT���r�v�=S���z�n m_p��]�T���{�-��g~�oq����Y�<B��6�V��5�%�p�S�Q٦f;��6�!�ܧ�
�N,^���N�K^�A������x4��L	$IB"T�u�:lEu�6�"�'�W :�-�U}�{��E����uLH�<�je�]��\滻���[���p�U�\���A�VS�,��k�!�����5G�:n��d9��f]���m�s�o.��9e���6�q� KRwcvsw���g�-��dgj'����Kk�������:9�b��N�č-����g324������gx7U���������C�po� 悖5X�*!�Kq���.��[�QjZ��3'��N�m`��;�hڏy�n��=��}g�����K��_ ���_ueQ�޽�I�A����y������C�W���n��U���mX���
.��Po'GoN����W7/���UZ�����t�4;z�t��.�ܧ��7�\z?t���!�/��m�m>}4���$+�'��l[��3�\�h�	���ALLȕ$�2Sk�fй�AL���E��6���]�0����*��ֻ�u\
�-�z��6܆lZG���N,ʨ9�����|�lEDU�_�U/6�7�+Ur�5{F3��E���@my����C�#1y�9u����4�\��i��Q.����mǛC���]3��".����;������"����N6�n;s�f6a�z������I�ܨs[s-�=6�K��=~�~z�⍰u&@ �cq�:F�0M�*C[!�-�9i`�J�4�m� ˇ���8vY�f��1�1C.ƉL�3��l#����J���e�%�0��%�:�que��K�+�UEiq�Ҭ(�2����nf�։t޽�^�{�#���3j�}����O-MJ��d6��Ϸ�<��炝}�F�ֶ-�ЖS<3����n�$ЌO�l^v�N����y|mrU�'L��6܆U���K�<�=�
��6�������'xR�{���6�n�VGw_DS��F/��[nC!�0�=U`������\6�W\����<�+�Jk4CX�V�WM0�5iЂ%Ծ�GHE$������;�����T�-�7��Z�|����]��C���6�f�7��Z5�#��jtU�:�ʍˍX����:�būz��Uj����ws�����j�!M�۞���W�}4۪�r�>m6��W������%�iԭ�O7����y�'����p@6��AT3�Z������3|�@6���)DR��"�"<b6X����k�驖S!\��x����n�2w6yj�U�lQde�jgͷ>n�3<��������U7ͬ�t�VS.ޘ�I���o��1�7�'����d��G�yIsr˕x�~��xǷ*+���^�t̴t��<Bb�P�4n"E<Ƚ���Y�wͰϛB*�[Dc�Z�6h^f;��.��;[���Jm�>d6���`��Ĉ:�wK��o�ZCk͈�v�KR]�`H�e�
�֕����k��-+1�{�I�6��W����8"o[�:����{v�i��}�J�]��;�t]Uuʼq �;�����m>H���ޞ�����K��z����m׫��|V��/~_�}s��	�&�mɜJZ�b�TL4PJ&�����w'��p�M���&�%��,��L�)�ssOcqv�>��U]ks/k���W��pi�I���E-و������Z��L�[#m6���-׻�9�_�<�bl��w���Pg�������qN�������<��5�8��ݨ6�6sIͼ�{W�6r��x�ͷ*1�
&��we>׻�9�m�5���:�my���Gk�7
��@�i���qn���6�� {3&��5\N�Q-Y�\dTlBR��90FdD�'��{���ެ��vv��;����U���N���u�(L�v��5�<ɵ�S�o��Dl���Kp�Ev��y<}�'3E�^��}����U�Nc�{�P��q� ��]Zo%�f��*źI��0D@��Ld,6b2֫�Q�U��7f����E{[w�(�1{�9����{�ٸ�v�N�u���f�����"���0\2e[�f��u�B�x�$�0�/V�'�q��me#?'��e��O�j�SAj{~o^�E-yvq��_=������y�U���:��X_hx����cD����K��ԋ��:r�G�z_�����qg]����r_����'�Vq���v�����`i�� 9W�?kDgq�����B���]�U����p����#B6�f�Ȑ�VfXHx�W%qt�`I�� w�r�.ΞU��f	�]�7F��x����]P���*ƻ��x��h�%��q���z�Y;����*j�}E7���L\����C&�_��fQ������(B����,<�s:M-��`�-�p�y�@PvWG$���{'nɉ��M���d<��Hv��'��tHQs��y�A����@���AG$�^U�v4$@EI�m��(��a; �=��M�k	H�j!^N���˭�W2��%)
�m�r#v�li�a�]�)��i(9�k��ڪO%t� O;�~o��l 3^ά��m�YR��2r.�r��#4s�)̸���fk�#J7T��m��&��c��)
v�ط!lt��֗�
lG�# cF;Ŵ�0j�%Y�!M<��u�YZi���fQR-�
��l4�qI��%lG�f�4�0n�(,�ًv*D��0D�,e%a��-Z3,�
��5�ul��u�fe�f��.T)ss5�F�\�؍ڈ��VR�i�F�X�AVm��9 �Q�`�&ƍ�v�v��X&dF󋀼�x+kcj:m�(�s�W,���(���Kb���F�#�x�J�e�3�,Q�k���v�����B�dn!t�cC 6�RPM�mDs�E�rM*��BP���j��d�ޣqj6WM���gL,��lmH��V�h��.�<v��<9F�����9l���b%��Z��Au�(٬
�����m�DV
��@��	�$v�JZ@�Ƹ+�uGsM�)YqC���fjb��:���6�YbM*�Ě1�(k�kl�Òb�b��4�ǀ�L<�Nշ`�U�6WATV:m�]��arUM���rC����&�@��aC	m�F�Z������iv�Q�Pل@��Õ6]tW�ʪƊUU�F���Lr�[v��bj욶.)G��X�ͪ�w::Z4̹%ֹ�`#�"�f2֊���C#Wa5:ڌ`�v�;�̴�Mt��%�d֭����Mj6��q;HE�v����QXk�������cƘq�"�3v���K�.�2#K�6��f�m.7� .���t�nЄ�l�tQ�X�,cS鬿� �g�ܺ],��a]3�\(���L_���m�ve��5ӗU�Y�g+Uku��י[�5��չ8���)��)�����y�26���Ӹ�m��ӵg����ź����m�T��iDu�ec��Q�u\�'�9��u�6���V��)ݔ��3|%�a�i��
z�[�_���'�DI�:��ev�o��o<MH�͸5 P�g��^|�ѧG{��qn��6�r*��	��>m�q��x��܅�ܼ�[9���%�"��o�f�� :�?-�����9�W-����n�����ϲ�zTveW���F���F꼸m6��r��m�h��s�5L�xM\�����ɟF,>���lou�ź����!�ɚ����N��Z�ݻ�u����fUuʬp|���t[�N<�L@�b

�2b35�ۙ�L�k���=!�r�;��wG)�%��.T�-�n mTU�1���[�K���c�2/�zkoXN�ǧƼ�k����z��G-���mlNp��8�5��w�a���B���.6o�r�P�ܤ�5�Կw{�/wI�*��I�g�~��q�Ř����+�tr�����75Q���AѼN��^f�v�_Lc��}|�k�$;%(�S2dD�0�P�h��U�Ůz�ѦYL�s�3�jh6�n����וXFUҊ�t�y�i��aD�<���x/"�wG)��4���B"��M&�g���j�c6��{�3/�T㼞�ϛw*��)�@e��r�7y��ʮ('�2����� �û���wb��YOz/"U�P�Nem�����i���X�/�0�C*����?)�c{�ۿ��\]�CF3D�bSD#�cmb&H$f&L15�hm&ؗ�"��λy���o����>m�m��Fc������:�R��w�1�8�����m �l�P�/�gN��3\&���m5�3.\!�H�Z[FX̋��<��OZUPc���my��u��������ٛʩ���7�ye�pP�9)M���N��|z_v���-��h�w9G�a��*�;�ʝȉꗁ󔩎�&&��.�\6��B�\	ev�W�����c�Z�0e��.�LX��\��FXb��X�.B0��TXԺۀ�Vf�q	���S6G4�]�	�Kki���4���K6��ۚ+�؆���f�F0ЌUr��E����׿�|�ݜ:V�c.n�,B�]L�X�Q:
K�1�q����^/˼?jU��{(M:�o��l���t۹�9�l�E��<��s"�7�Ln�\�������w�!Dr|{*�7�zf��^&|�myt
:�]��u�oa��S5�i<��E�C1���y3�7�-�ݜ�gkgy����=0�&D	v!F��37V���2�kv�E" ��H�����c~W�?{��S*��8���qS�؇۟7j�UZɠa� 
���]蚃5�z�x�zz�a)�����yP��o&����S���u5������_�^3˽�u(W�y���I�$����(���9��n���y��6�p��T$5뺏6�f�WoOL��w����]Ѷn۟3��}���vE՝����Jf�{�[��\`Ln���g�67a�K���?���m�0etQm�~}����,���>�����=X�##�8�}���� �X�Jo0*CnVWoN���p�3��%Y��-��Bt��9ӳYr�c�z�Vԑ��U�d���z9�B&��Ť�
����d�R��ʫ��I��Y��a�S=W�Q�h�R���g���U���ӕQ�ޢM�[����53���Wok����P�psQ�z�<ǯ��扇�Gk��8���v�!�V��u�ډjIL��������J%�Q�e=�wi�@Y������M���gk�Ern��]���-�K��{S����Ѯ��5��M��@�����/3�F���o%�KM���oY-]7�Փ�B��ޓ��ܨ�ܫ��E�30��jNN�w����09\.ׯ>m��-�i��@��]��V<��>�A�֋�Lڙ�mY�̃T��f�.XF.:�%f*a#�^�7 6��.���*��<���ؖэ�{��w�p�/ӵ�o����SO��,��������Lu�ۏ6��;��ݮ�{�3�>�^m2�:���]�����ڬ̹���̩�+֣��3�Lb�S�m�Ch7��u���ߞ��f'���ϳ1�K^N���ѥ��	0Bq�+�z3=�'	���\��r����1����"��t�ll��1[�0���l�����b�ƅ6�L�%H������+Jn��:[�^��ni.��[`�Mp�Y�]:�2���J���1^ʥ��Fd[�Һ%
0�r큔��L1��l�h��b��Џ]6!A�}|z���h�;�7GC6v��J�� ٹ����y��m�t+mf��y�?k�nU��_k�ϛM�+�=����oF����p�y�k d,ki�����qf���f�4�K^�����D�m�z�b�]���X�'�^�uT���i�-�nv�n�C^����ʩ�9B�@o�I=�����_O�^K�ElI�B<�D@��D#�MRms����)Ίz��\2�^y��[A6u-��}9�p;3Nӌ��9�	�����q�s8�gL0f�R��]�7yk�/���F)Q]�ۜ�o
��g{��c��;���ɮ�(#p���i�ss5v3{�7w6w#*�c�X���79{��V��tU��Ji�b�=���t�n^se߲�=!ޝ�}5�2x��6���Aл���J��)���S��@M�GCk�Z�4����Z��m�mgt�FUO{5>�Y,�0��i�nS��6��h��W�z���K^����oai�j�i�7�|�G���A��U?F��ec��P{9�U�.���<{4]7�6��z]���^n�s��ѫկ#����I-��{�>�w5�}�lܛ�\do�p��Yn!�������{,Q��ci65��+���}V�7Ph*\��O��巆����9�н��E����k4V��%e��z�^�����i�B&"d��Wt{7�wo����v��p+�Z�6��V>�K��k�x�����G���]�.�Ϲ!���o��:��ɪ�y����F*�b1�*op��59�����F�Ӓn�v�w�Ş�ꇩ7g�N��I�@�֙��# �&�A��CpՃ�^ܽ;5�/����	5�ۗ=���o�3^��2棇'�s=�n7��"o��Or�<-2��)�����ܝ���o4Q�6�1k>�pW���s}�|\��xŝ��X�M�o����<cᯣ|C|g����3Z/:W{D�.κ�p��l���}�w����s��N!��x(vק[�:Q1D�5'B���-U	D��AZc��CF��MP�"Rh)
�j��y�NA�@��ZGaB�!�r��W���M��
���Ga��<�)yy�p�Qȣ�%;�Ҕ���X5�K̓Jv�)��#Z�vl�)��AN����tĞ^O 5�@�j�5��4iO k�K��'(�%U�S��vyw6 �Z��N/u��idl�R]�vNCʍr��ڞ@�;�;-�O"�O"�^��]ù��{h��)9�hІ��I�9�4ikEo.=�:O!�CI�u@]�v1E�����uH�Ab�*ݺU���iמc������&��N��A��iz���mo<�Ⱥ���X�;]1�l��W�@2�l0��Eأ졗\o�z���-g��6z���	!�	-[�ң���y�ۅceѹ
ݭU�'���Pg͢������k+3�s�W;�}i�n<ڹ�|�Y�S<:_r�s�;��.�{�k%����3�3���A�� f��ŝ;֦�xK�my�Ϝf>�qw����.�ݝ��Ǚ������C��YU��)�<�p�F�ԝ�g������f��C	Ϋ�i�+l�8����nhCn*�j'wpmUQ���ȷS�kgkol�ޘ�����f��A ��]�C�՘�j�z���?@��de���}���n;�Rn�mCh	���y=��(��^�����/��M�(���'v����zی���ug���;"�O9^�h6��E�ܱa@�{7/tM�*ݞW4�ͥu�8-��je�A��`Ի����ڇ�/��6�vY�d�*���z4����7LQB��f(!��u6=�v����R���R�l�:0
���廤�GPtrM�j����i��LŴ.�e�1����f�2L)	��X�������	k���l��b���y��-f�c�1Tiv���T*Ӭ؋5eÒ�l0.V+%Ʋ���uY�c0�Ur��q�����>�f5�Y�X��U�U�b�8�RS!bb\}���6�,���Ⱥ��J��Ȍ܃���Q>�\�:���mQ��Ֆ��u�#)ǳ��g����ڬ�ύ�x��3��^d6���f�bV �!���_v�vE��h��o��׃��d6��O;6�4���^����e�<c�^+2�OM\aL��F& ��36�*#��3�l���fz�!�2Eܪ�Y����ޚ&��J�A��������E�Ք吔��ˊ��[J@���w�����F���a��攝��V��Qo��9'��5�}���m�pr�c�z2�,B1nN���ڞo8�Pn#ٔ�'��|C�[^m3��~���Ыqgss�w��8�;���u�Qmx6�o���y�hU`�����Gx9B�y�e�m�}�z�*K��6�pA��nq���KV-�)AIr����g�P�s���o��8��1o;;���<p�FΡu�E�����m���g��7�חsLeM ���nE�0����HtL�p����N�ΥHohȨ�V#�g[ZAN.j�T�C�ӈ�1��c�O�:�rm��*�[^m�<I�**��r��ǻ�[��<(<WSk�����u�{TL�de��՛��M� ��my���o~�>�;D>#)�m��S+�T٦�7�Ņf�"A[�����w�e�~�{{xFu:�sL5*O�����qy9K%�N�IS���˝������6��倪H���A���-�@�#Q��o���M�w���[�-����Z^�ͯ<��{xd�:}r�]d��#n�3��^��3t{���}$*z��x긗�O�Eu��V�Xi�U���=������s��ﶂb뜌�����KC[m-]���
&����!B*D��M]��_���2��$T6��<:�Rdў�W�Ϲ�ɫ�k�e
�/2��)�b^�n�گ\!��'w��NӪ�r�Z|L���Y��M�]8��}�z99o��!���Z����묏��*�Y�����7r����!E�i��ۣ�E��H������tR~����`ќ��G~OρÇ���Q[���Z�s+ϒ�I+��>��Uk��F
���Ay7n�wI �3�F�)�j�:��0hYm��a�20Ҷ�v\�d]��� Q� �eۭ�V����!SvͻX��`Cvx��!6��аJЎ��5��%A��{�.��ŕ�vjPV�\�b����fr�s5#�խ}�������tcqY(�ܳj��`�S30��K�ۏe��^>ޔ��
�Ʒ��リ��!�m��H*e�@��FvUm��p�j��o �ɮ	._�6��Qmy���?�-��>ܼ�ꚮ�C-3�6��e�]���ۜ����9s��s\�B�L�6�mȎ��ћ������gs��W�d�^gѮ{9f��+331�6�����R[�wj�ЁS	��6���Z.��u'��P��}Y��e�6�A�#��S�7o �19	���o�~r�y�^Ɛ�uJj�����F��ʄ�i������:�1��N\����6���v�"7*&� ���ۏ62fmU�e��臓W��y�g͡Z�ژ��;q��u��s�����z���*d����N&�g���Tz�n��n<�i˞����ͯ66,=�����g5t�.���&�u&RR:jfu�Tv�߮��<���󊣻��n�W'ӝ)���2�m=p�$�Ӯ��{�\t:�R�',Jn+"�
�,�6܀�p>��PΥ�U(%m~ȶ2eTe���8���{J|߽����������P�w̙m�,y�I˞�kpO�k�Њ�kX��d��|�K}O��~;Ux��1=������w{V�w�r��\�6�6��>����[[����̦�s.�6�ٙбZ�˗le���=y�<3�s'�Rr�s�:�2�m@n�/B�͢��P3R���t'�W�{����b�5m�6�9���ޖ���V�W�ӀnA�U��yʺA��s�8�z��<%�gED(��;Vkq�gL�ݖ0����_k���*����xz�/�w?6~m�������3fj��t'�Y�d���q�W����|��sB�[G9�(�Ƭ�`�f\�v3k���~|���<���͸������5�%�p�mx2;Tf�Ȅ�����s�9��E�<��ͫ�9�Wc����!�7��FftE��s o7,�����S�wq]�w�s�t^��r���qc�a��d۰:�f)Bwc��3�r�}-{k����~���?��q"?��:�(���� 	����� 	��T� ���ȭX(-b�>�(����X�oeja�C�^��H 
E�B���IA�5ڒ\.%yA��jB �v���$��n��ӿ�'a�o����1�\l| !t7i5�7�k7����ur�$np;ቬh�� �����s���!A�	 ?�2rB ��Ұ�
���w��ϺM��~i,'����և��ϴ�|:d�G���  !���_����H*pKk�,���d2ZQ��{|$Ď��Ef��o`��-�ϻ�'���dT����`�a��I���R@ ;��ݫ�s�̓� ����/p*�s$��c�i�V��X4y�z�?��O�H S$�B��~�{�����?a%����gIi�����a��$�i��>��G��_������R@ }�������C��O�|~a�����56J�$�����)�I8C���>A�;��'������4{��� �|X����C����"oa�݇��?6dD@�!  B��C�$  �����$O�����T�E��įW�6bB{@�&}�$  C3'�ʣ �����F��t @d�I�B�L�`���&1M%D����d����a�T?N�������# @ !�`�~������ �G�!�������'�?w�~����D?���K�w�G��[�|�|;�ϟ_��C��[�}����$� �2��l�_����|>�@ }R~%� tX���O�s���M�Ԟ���}ړ��#a?<�\���_�����s?��������Tfo��1���@ |yi����W՜6�=JOg�C����yX��^�y�����C c �	 C��@�?�I?U�H>�| �_��^�_��B ��I�'�a��r�!�B�ؓ�O���zI>�'�� ���?�.�p�!D<�f