BZh91AY&SY�)����_�py����߰����  a^X                �DJ@$�%UJJPTEJ��J�Pg��J)@ I �DX��h��w� } P�X��Ӿ��������G�;zt��k����;�:����( �H�%_C**�����<�i��T	*���H�G���ϡ��Ж��m�!U�Ѣ��J 
�:�<�@�e*�EN�{җ���o;Q-j��ܫ]��F��j��x�n����=Z�2����vW8��n�vd=1졣G�

)  7��d]��g�]���zE�k��WZ�wqw=�K�vN���^�s�`Ͳ��*�^On�P�]�=�G9�U�J{b��vzq��pz
 ��������=1͇{�^�����a���g�v���<[ofݘ+�Pƍ;�s�.�:�e^��F��Ξ�E�*���ݧ�]s��$z (����>��wk�t��ϽJ���v�����{�^�6�����{�:�u���x{��n�'�+��Ǣ��ov�u��(�|vR�      m�@��P   
�� 
�     �~�jR�CCS40�LL2`�OЈ��RFh��	�� �y��h �� h@M"D�R�2`F!���d�bh�D�Lh��y12��eP���MM�SH)J�i��@h�M2i���@6턐��@�E�cq�(9�\S���26(*(����A �&� ���QEwIz�k�>_���� �#"���Eb�����TUI%W�ܪ(�x�	;L������ V ����C��u��ur��g�(��Γ��I*�
F@���_@0v���0cܑ�#S	�L��9RP����&#З��S���xD2)z�#$��uБc(��c({����g���¡�&,#�$G�&{@�3�PSJRd�sd*p���3y�f��Iiz�IM)|F�K� �e�q���p��_3v!|�JL�b!aC��ǝ	��
��%	E8V2���� 9�q�!h�����4��p�cJ����diIg�8�XjQ"fB�T3�ĘY�����K��$V����.p�a��.	*�$v��1��r�H�F:e�q���c8\3�%,�
Fi8�P�о��+�L���	����;��H�2��2M,���U�D, f���1��C0�1�3�K"/�H��&PݑF�a��&a��&md.#.�(b�8\h�6/�҉_P�L����1�B�p��]�0�[���r�L����=�0c}E�PƦ@�|��j�Fa�$��NBx����e8Bp�ƕ��S�P1�.�|�M(�8�o��f녃+�q@��\F����f���2�J�ac�c�"lJ͡��W�ar�c/�1�@�%�1�cL���!!�ez���!��&�bV�4�dk4��'��w�F�Z��D&A�:��\��6�r�c8�p��c*c���i`�N���Lfs������A�8\ar�c-�g̍#���[U	I2�@���)�!���PI	X0J`��|�q�@���ߣ!}#���7p�Y��±��.0�p���.0sP�#7Sk�R#
��<�Lc%�Kľc��>�L҇�,c��cci5Ьc&��ɚH�a1�������L%&h�;	��J����)�eU�e���f�ib�JGJJ��1�p���=P1��-,��8X!�֠��\&1�ՌΤ�DH�f��!��!�ќ7Qi�ڒ��hǫ�Y���@�ܢ4�X3�aiC93F�HǋFH���dbC�����e��3�9چ3	�#�5A#�C��#](c,���,�0g"��3��T�L������g9Q��h�P��j0�FK�RL�&k�eԬe�e!��(eYm$�c$i1���|���C���:Qc|�g���Q�z�c51���q�T2�3D�3�"�E��1��
0�)1�+�z��ư�ZC��A??�#4��fY��3��c�Q���Q�}MD��t�����G9Q�1�Q�H�T|��ڌ$���j���d�f!8dh�$ɸ�x��xҏV���ܸf�IV���<Lc��iCi�<P��mFQO���;P�,����p�ҋ�l�c�%8�5q_���8�Lq0�h���+%�(B��D�I���&>j�#L8۸L���ǩ�\D
���@��c_cM��\]�w�Qb"S���KHӄ�/��bL���)�4����c%�DRd����L�Ҏ0{��J�'�!8P�,���#�<P"@��5$��s��3�T�>�RK���|�5�>`�CK�)IC��!&Yb0f��,�:Y�),f�C4ќ�Gim%�$YNp����Q�r�⏟�T1��F;Lg6��֬���1��E�1��C�0�_�D8Lf�C1��F�c�͔�CT@�x��16�	n1��V1�|�LĤd��L����Q�T2:�8c�x+:�0���ҊnT1�|�Č�{�v�Y4�P�;�1�E�'12�mF�MD1��3F;��Iÿ�;�"�I�ڊj�;*�h�|6��˄I��c�ǩ��>Q$�B;�x�F�z�8��'��>���_��(��Ic�'"�j|��)�&�f��c�0��1�����RX�Lc0udP��|��(��c4��,�1�XD�G�G��Y$��?�0fK���j���!�5�+ ���$�!37и����3���Z�3K�D�Qc ��(e�alJz�����aN� �ިC3�k��L��<j(�$|�����P�H�(d	ڋ-�:(��I;�I2�wv2^�QC8��ID��iFDA	�(�P̱�1H�3r��M���G	�C���C,mY�,������C��،8婘M�q�J �����p�iG�m@���hB���'K넞&8؎�bwJ��.��	3���@�Уh͵�>PX��#���<J�_/��1����I�1����C8������G�$1�	�v��|��" 8Q��)�ƒ��֬��(����Q��i'?���6����&3\�e�Z��2�)҆3|�F>�P�2S1�ԡ�1���C�p��,��aCQ�!�0<P�,d�<(�_ɒX�v��3�Q�(c��hͥ�jI�LԤ�I���B?��|�mQ��.�2�8p����c+�3!1���1�	� v�ǩ��END��4�#2#���5P&%�M�߉�2FFR�(aO��}J(f���f�6����'�(t��c41��fϱ��ә��+�#�!P�E��.�V"�1�&p�Z��W�f`�2�3���,ʱ;��RI�2��I���p��K�P�VC[�>�Y$�
E�&Q�g3
̅��X���D��)ϴ2Fk�n��BcĹ*1(L�r�c���+%�iq�2��@�K�j����AJCK��9I���YL;\1�Ү� �H8�#)��H�(�YP���c8ı���-eι�B��T��W�4��T$��|���Zk&�W��^��?,no���w�:l���,�W�	=�X�'[ٳ����}�Ӻ���t~2��m�ww2}�i�Yǯ�q��b��=[^ڻ�a�3.�z|}���,tj3Oݟ��ג_ٷ�ּ)�:�kʨ^�Q=�Y����z���P��ڌUU�q�:���)�fFz����ܜ�j]Gvur��W�9�U_t⣞���g�>g�X�w�S{V~j6�Ws.m�ج4ݳ�U��:�����.G���8�+�w޸��k��O{�̹��<��"��Y�nl��tU�10��ɛK��KJ�0C���UI-t�O�g���#鷵V֋[͘^��v�ޣ{뻨��Z�ax2�w�v�ii�Uu�j��e�֧Ok� S�ճ�Mj���)!N��=��ȣ^e��/���p��}�E�w7$UF��x��3vl�5E�yB����w1�ӛ�33��ٮϮ~�޽/gEOm��H��'{V0ǻ������v|ɧý��2d��ze�i^��=<�;߳�~�����m�q�何e�����>R��/Z}�����h	̴�ڛ���6�\a�ٌW��uK�)TI{�yȼ��침B�2��R{��u�L���{�(>�{^'���&.�0����eӡ��X��I�����}���^�*7'��Nᛝw�/�wv*�s}[Q�i.�c��_������{���wiU�p�ǘ%jһ��6��n�m\Y)F�395ܫ7�䛚�2"䵻2Y��PU����]��Ƽ���Plj	�{r���=ʪ+�雟T��k�z�r78^�LV�Z����b�޺��mGfMdd���HË$��ӽ�v�g/s�چ�����OL�d��=z?b��d���v?<�̞��K��6��b��fL�y�rލkw�$����^z�f㣗G��}���d�;eط���������=��Y����ֺ��d��
�>�3�h{2�5�M��1���B�:gk�OWs� ��|�ϡιd��������K������l'��+ߎ�s>�O&�R}�߼[w��m{�Q�^��[���e���������Y��""d��g���'ʞ[e��M~̒u^���*"��Z�N��ۅӞ�O�{J��=	��&�z{�m�{3wI�Ϝ�O��Tv�Q��Q�J��K������.�靻��S>op��v\�FFd�)j��fu�yL�4��Oת�:����j�u-��Ȼϻ��]��\��\VL���{�!�.����-���>�K��u�=K3��2�n�����=����ِ�w�3��:B`V\on�٫�˙���v��<���Fܛ�UB�Ov�ś����:A�֥���ӯaÚ�\�ԩŗ�R�=�����W�ܥ�tD�n�U���|�'w>���rO_�ߎ���ۓ���(#�eZ�����~>�oÍ��y�߽駻&�M[���/}�Ǜ�=��=;O�;��r�M��6����v�vY=�{ޫd���g�{�S�t��C�[����l�x���>���>�S;��>)�%���z���݋y([Ź��OJ�se9��:��$�<��*�Q-x&L�J��GM�i��Krx~އ�c>���}'����3=/f��;Kަ�fg��*���O�m])�̟[Y5���wf��"BZ������ѳ��ۛ���;w8�w:}tp����M�u> ��U�WFϧQB����sf�2_�U������0�#پ�������~�{3Ǿ��r1��ٞ�{���Jw�g���-��'w��b�Vx�׌�?�C�ʲ���q�ޜ^��7$����T�o�{��{;���p���]������7f�%r�r��'�<�7 i�~�xѿO��y�cŏ��.��������j+&�Ͱ��r��{���ʵK��NKJ��PM��9;ܣ+V��Y}��eMn�Z>u�Mv>��|5���f��ď{2H}������i����A���u�كϦMZ�z{�s���*���S��f�)�����}�������!MF��:�m�1'Զ�R|��n类-�(����<:*�k��V���M�{f�:gMٷ�zq��i�۸�l�曻�Γ$�۝�F��D����ȋ��w���'��VϿ?��}�]�Z1� }��l����;0ڛ><�<w��s�6����Ϧ�}s�����s��������9�;� c��v���g�K�Vo�F'|��b��)Ɏ�[meV\w+J�7��Q�jT_�s^��<�m����̸���(�ا8�;�+���=RMN������`(���m͋^�~.�s�<1UM�"������j�U5��;we�Gֲ�w�s2ν����ݤy�޵.��{�(t����76o�����s*�g��ְ���9�Ͼ�rg��������+�WյW��l���m�a��gevuw-��ڛ����G9�\�D�/BS�Sh���b�6��\��l}�r�Ɉ&t��nvk�'�/S|B��_ݐ�;`}�)������z�n>J3;;wrfU�#k2s1�c�]�:�t�T͒�	����:Ց�A��f���jì�`o������d��Ga���B��%{ɭxU:wHK���v�_L����2��{���顏�2R&�<��2��<3�_~��V{���
ܡ�����oMMZ}�<к4��ϲJ2f˷UGk�K��&���}ř�&��E��r~�v���yĥ�����)(��GA�	���|�{s����N��9?Fv�p�xpp��˝��KUD�֮����m���x��9��3��i.�)���s��7����8��mc����=�z������y ��*����/��k���v=%��r[$YV�����}����9�d̏%�!�5��;��op�w����b����5��{���ݛ,�qkȫt�t=��nU�t��	�Y�f���۷�R#`���ڡ^�Qk���6"�����䴵���2s+z�k�32�]�ٵ\{�����M��+���������÷�ss�f��1����_����Q���Y�ݘ����ͻ=��f��c�0�jp��W2,���(�v�����U���$2�A��6m=�^�ng�����4}�����f�w��_�{����y$��~+���'��'��_�ﲝxV?u9$Gٺ�������2�6����i�,�Y�n���'J�?�.�����'ak�k۳=f�	ɶ���beۨ��A�ɼ�p/6m.-����Q�S�|�n�0�ack,�)�eq���m��m�i���n��6�il�J�+`)+	fq�66/-��/%�#��Ү%H]D�7��\Mi�oV��Ł�$�Jɋ��mZ][�1`=�o���OK*e�*N;��Aj3\�+£ �4܆,�׫4ԙ�-ڸ���v���po���T&܄���\�WT��q0����[ÄQՀ�Q�������5uK7�J��{/��%��3�,�C�_�,�W��J���v(,1l)�ut�46���ˆb�1��=�����ig索�?v�������c�r��KY4Y:�o=����;a!QYi�/gmf��+)
�n��3:�6�]e2˰+3�+\,��Wi�`	�xc�He*��fʦ��Ҍ6p]#X�ajS�]ڽtÉ�e���2�k����԰�c�4vts�i��.ZL���m�,��s��f ;f����dڔԱj.���FҤ��fݢ��m&X�s��Ѻ�f�����VY��#���o�����F��$)��Յ�l�u���6�A%	u��iO�Y�Z���/K�J�/5"4��_�p���EQ�u��CF�\;9ŉ�l���6�]M�at�f4T,6�6�X��oQu��"��9eu�X�i�Yʿd�[[��E�)cS<�<ͥo#x��)ҩcQ'�����ǡ7���Bm�؛rIk��27EkI������yڧ�'_�TH9#��'������\�@A2�G�0�����M�L�n��&�����g@�5H��;���`M<:��:��4���Qf��9���"ٝ5˜k�P��J��Wb��-Ԥ�MY*ǙƳ���������/��-�m����5�75�3[�Dt�vf`LT�&�(8n�0E���V;�����а���ʉ_��.�����v?��oES)Q_m����ҼE��By	(�g�mc\bj�F�mY،������ȝ����K�R�!.�[�ܲ>�YXv:��N7�j�N|&�p�^&vԧ��Zأ#j'6�}\�& "s�D}^�"�E��.l�aĴA.A��>��}ځ����4�@T�f�Uk�Q�}�&$;G����u����m��Ȩ$� H��wl�m���y�y�<��;��<�<ۖ�oM��|��m���m�m��m������-��ݶܶ�x�m��m6�v�t�r�m�m�m�������������(�R�R�"(P>�˚cm���m���m����6۶�6�o[M��|�m��i�����m���m������6�m�p�m�m�m�m�M�����<��U�,����2睮m�m�����m���o[��m�n[m�m�m�M���6�wtn�����m���o[��t�n�p�m�cm���m���m��6��>��Q�	|	!}� �{�>���m�m�m�޶�m�����o�m��6��xۖ�m�}��պ۶�6�o[M��|��m�n[n[m�m6�m�i��o��m����o>>��	�%���_`$ ,$D�Q@���E��#��p���< 9��?��iG���g�K8�3�2��2�(eaE��!��Ad�і1�QC4g1�p�q�8gќic4�Leь��cc�2$0c�C(��1�1�HÆ�&@� ��:�F�4��GN�u�Qպ2F1�1�t.0c���P��bc8�1�p�F3�qf�f�3�$ђ3�0��!�C�K�(��gX��!�" ���bb(c(�`{������~���ˍ��/z[ɩ��dm���fͬ�t��X������D=e��>m�e�ٝ����i�h���=�	_<*�u˼r��Rj4x��V�P��Zݣ�ju���nv�VT���h��R�ĥ�����	���"�-��[`0�T�9&%x�0��4�h�Z(��lԔH��-����&�-2M�]�bA�h�ҋa0\ËM��\��bP����4�*�І��H��vڐF��($��m�(�r�][6����H���%��k)k5R0%�wn��gm�u�X��Z��
�s	!V;{s3#HI�(jp��0�&�vڍH��,�Ͼ�q�|��51k-�Zl&���)e��Jn �����̦��P�H��u�]����x�Yf��L�i�V�v,	H�В٦��ƈ��`^!Ml�]�.�������ŕ&��� �[�� ���F5�&�Gm{EҒ�Ue��
��Ɩ}�,89�R��s�<n�k���|�R��k�l��{Ev*�)��V�em��t�\�,�v�e��u\�`"䵼�lfP�����RRA�#�fٲ���6�a�����9<����������9�<�UUS����{��9�s�z�UJ{����s��9�{�UQ^���{��9�s���UB�Uf�yǟ<�q�u�]a�����W��0~���ڶ�C���cX۩t�B�Zm(k/6�J@�훭��b��Z�N����݂��'��~J|�dv�f��m�cK6�[YL��M��i�U{A
k��Zg÷��/:m�o�i�I��
�Ou!E�-�@��XA�y�@�I꼣vB�&�j���$�����<W���~���ggD���a��4������V��	�|��%���02h~0�6�1�M��k��J����'O����zz
��*�ީ�d�s�J�u�ΰ�<c<p�������qŜ3˄�]���%��rj�5L,���m����IGޤ�&nm�a���];E1�o�r����l?����\�)���\��U�NDMD�K-�g!ʽ؝΍T�0�sȶ���v!֖K��"}DD���B�� g1�3�i�b�'Y�0r>%}
�(ã&B��n�Snm�wnf���!�'gE�N�<�Bk~��Y�q^J�N@hSҩ]�� ¼5���,8:>�Y�-9��*ѕ��$�m�J���D x�M�u�rR��昣,.��]F�F]�V�/�0ќ3��i�b�'Y�0��|G�
�`I'wAJE�@�)�ђ��K�ɉ���wk�ʐHԩv:�1�>C��!~�#�x���НJL����ц�
����ˏ�y��L;C�*_��y�3.9a�aA0�|��-��l��].���q�_:c4�1d���,�N��®�b{ۈ�[ŵ�]���ݿ�>���I\M�d��!zJ��S`��
�3j<i�@}ى��`3B�h[t.�#�m&�.q�f&�]�
�Xt��2��*JM6�4�y��i�Y[��a�����z0��=�U���eV1*~�&�>i�M!�"���U�L�o�^h���%����u��r���ޝ���{e�֍<�)ϟM^1���r��mR�lz���I�}�Q�Er��ʫKx*�E߆v`l�BQ�R�y,�N��Q��3`�1d���,�,l'L�&�nҡ&2�'�X��zY��u���Yq�|��/��e��qr�w�?'�����<�hY�#�b�ѽ�/��]"Ò�і����j�q*a�RF�)1�����>��K�dz8���Ҫ�l;�	@�R���6�����l�����m8��`��!���qŜ3׿�>֬Pv��-= M��Uz)�B���[m�|�Ħ�5��â�\_a�Οv_�R��e��J�ٻR��.`Ot��K$�"I:��v�V)�#��J���rIO�F��!g�;*G_I��JS�y�;|�ζ�h���'Y�0�^J�:"T!"Ek�oc���U���Y\N0�v�4c�~�>���h\��01Za���`v=�0_�jS���>�^|nTBRB��
�U����0�&�\�=���p���n'�ܐ�1g�B��E��(��~��O��bF	z���R�a��q��h�먾Qyyb��o.�Ő�&ԗ�I�T�!�C�j�
B���#�Ywyi�����Y��+Gwւ��R��9�����w;�jZ�����f]�� ��	蛄*F34�M��arV�qK��n�Rz!����<���q�1U��E��jTv�;O*�׫l��5Ƃ����:�R8H�p��%}TҚa���Tp�vq= �B�!�(oE��尘1TtD�q�b+B��,�b��eT��rH�,=;�FC�M��(D���0ӆ1�X��C#%��:��ޒ�WlcZ�VFN�G�n�lr��޾�+E�7��CFr	����}2a<��������7��U��v˞�^Y��0��
�b��M�Z��羫�ľ��vz��G�!�����v�n�����y�8��#�_�8e2�b�q���H��#�	x�+R�<�'�b��y�{����������������|�:�^_��������^8��<GF�0�6�H�M<�2�'�����y0�O2�<^^_��e�<��8�'��O�?1�L�������yk��<��-4M$M&�����y������)~a~b��y<���q�O/ɗ���1i�<O'��/痧���o3����α�?<�?/����m�>O2������:�O�[��y��mw>_�_�_���y{KO'��=��ƞc�>c/���vN/i�z�y�Ğeyau�����'���O�Y�<Y{�}���'�JO�}4fAtS�ܟ�vTOL��C�7�����x�Ux]��ws�cm��`�H5�V��*nޜے��g/&���'Оo�g[}���k+OL�M^y�wg0���j��s,�{`C��A},�djU	`��	��	����3u��1^|-����wwv��x�����{{����ᇽ�{���www{�>^���{������G�q��<��מ[�0�L��n��I$��WT���ũ�6FD� ���$� ���H�&��녌Y�
��j�@���_n���2]R��,JD"��R��*�RP|����m�j\���jr��fg9uy���r�4�$������_�PJ>�>ESmI:�D� ��x0/��5)���Ѓ���ypB e�"8�m����(�{)A:,����������4�4��,��$!P&�'Ɍ����.!����l�:�u	؂tJ�v�̧Ԕ��C*u~y��_��m�]y��4ˮ���;U]�I�EF"2��aF����S ��mICP�P��r��(����|h"=	~��sJj�� �'��������A�	�a+$޶�JzlQ���m)O%Q�%+[K�!�:2Q���9�6*>pYM/�R�^��(q(�����"��v0�FLC��C�'ף+���""l�VD�в�P�O���DG�)]n���
����KĦ�FЯT�.��"����O�ȶ@�`t�S�Ti|�κ�����<�,����4��.�A5%���WSIr6�
�Ɩ y ��Z�z���[a�Lo�b�!�[���$�UBk��M�׎2�G8��|�<Rw��޴���v9 $��B5���*�1)/�2�5nw�Y��n,�$ŕ�^jC�PMK,��2Գ�EL~UV"&�\ۃƊ�%3J��<B��zw�c�9<UC�!"!�d)�"���N�����z4b�	��	���W�Ȉ��*R*�S��f����U[DSiB�H��������$:�$�a<?SRC�h1:�	�N���3���f�<�'��Qa��!�%+�B�@��H����xš4L��s
"x0M6���!�d�#	��ϳ�A�X�&x&R���7mn[�g�b����`���Ia�,��N�D�a07��ꌥG��1\y�:����ac����<I����J��P���U���I9����0`~Ѱ����	#	c""$+!����1=Q��~��H
#���H���,9���C��Ȟ��hd��d�	FG���%	*R�"���H`�I�I�='��͓��'hAUR" ��T�GPb��J�p��DG�����w��qn�m����ݬ�Ήwkxi��Y=<�OK��HpaD��P����O`�v"'�IF�@�2;����E�*9'bN!F""@��R�!*r$�;�C	���c!؈�0�N�R]Sb��-*��N0�<��8���מ[�0�L�����؜p��`�����D��Q��$с�V!��B�|�S��7uj��
���Ħ��d(��� 	N�$=�cd>�{]+Q���#�D|�DbRE}H�e� {�Xq$K�82v%B>�y?Y�j։�������RC*�D�"�$qL���*��J�F=+h�b�l�d�~�ZĦd4�!��dI����" jO ��$�ȅ��!؛�h���`��{:>�%�3i�u&�(�'�d��M@��� ���v0:E7���
��i%@�M�i��I0K�z�E'�x��+��mo��??�������y�i�]mלl�U����Օr�t>��Dd�d?��SD!��-!:;�v��N�$șVh�`�S�4n�=�<OŰ�"Z}�����4,�͸�`���Jg�J&	'������cL%"U��}���*���;>OZרi� �����v `ñ�r2�'�J��Hu�I��j5)���H`����	|W"!�@�A�̅�qJ95V"�F*�Ep�!�'�)ZC,���0��E����H��ŲN�`E�>BX0�JT%U0=�!���������ag�(�ef񧕛�RH܎C1��<��eAK�x!���X,�;�a����ɈI��Jb��o���	)(�+Y�)r*f��==Կ4�4�KSZK ��l����p�)�M2��mS�e+�U�}I��ΰ[� 8%���o��
�'wLS4lp����e��$;��r���1n�]@�QĊ�AЋb�%D4�������²z!�	��NA��(��A�;�'E(�f�Q�Ɍ�hA�Ę2u1�0�4d>��}��<��g�r����7>��F����]��h�-C�KF�UZ��*<��#z����є1s��g�ry���g��T�����7P-��#��	�X��%��K�2L�dB{��D�8l��;??D�����q��[i��^[�2�:�n�vti$�}�UD�����|�0O��C`�	D��6h�4�Xp҈�RQ9�aĤ�_�'P���-��a�����%�hb'��6��aU����$}�$�R���W��:�"(f����C����ˍs)u�ML�3�i[m};6�ַ�OH����e;�Y$N�7�١�$��J ����N��"IvB�I'�6g�. �"w�>��\�26��V���ы�g���xpS�JS-8�_�?<������2��O�N�0'�.�c?MUU�)�-�_c�>��$�t��bL���R�r�4�n�Y�<�z�2e�����R�� �C��l�4��uD�r��,��bO��>}�|��bۍC5�:"�3J��9���4a���=�-L�k�:��)�Ԥ�"3��d��b��Eq�e��,P�ă�X��4��QL��(`�Q%8S�3�Kȥ,��OJAϐXS���vt�8�v���a�������κ�O���<�/0ˮ���1�����q�$�BA�S��1�6�=����}4N	'��)>24DM��	�	L;)(��v>�ۙ�L�j�l�pˆّ��a�����f�4�a�#���W0����Sߣ���+s1p���C��H�F�#�z�.aM�����b�&,��d��!R�a������~F�8h�UP����%k�.W��b��;N�OVi��5H���`�b-�[5�Z�co/��cϗ�_�:�y�y���M��y�'�h�K�k�K�+���<yz|�0�1��+����������[��y8����<C�G����'�F���|�lZyl��y���������Ǘ�W��e�<��m�|��y�^�_��<Ǔ�\�~'��/�/�.����p)�O���UW����~e��̱o������0���j���<��_����y��x�=ry=&�W������y~y�O'S���y����3�����&x�L-��<t%��<M�y�=s��6�<��O'���y4�y���ؓ�\������.��'^a�&�[̭o0����<Di>�#�o	u�0�n��zsj �7;{��Ǳ霃a�6�$'��)�lq��X���5��*x�SX���M���κN7�y_3������:-�*�A{ˀ06l�l�Tud�e��)�6:<��^��F0g�m+��U�p�Y�E��2*�������pq��H?����߁��C]P������	���>EyZP������]2>7�;T�vY�U��
9"O��mJ���mօc�B��j�B�W.eh�6ԧf�Λ��V����M���:j��L=��k4:�_WGE'c6Lke�����ǜ�"�ݻ�m��e��ӭΙ9pzn��G��5��;��;ݷ��	�����"=�)�+��˔u*�Hcq��*;�W�O�uH?^ES�g�?:�����T�[��K��\u����D�u��=im����fx�T�zW�N��S�˝����'\o0W�aEk�y]�?�{D1�Ht�cǑ}��A���?�7��� ����5ńվn�cf��b�If���8���ػ`�T"����Y%eQ���.����f䋨	�ؔ!���hhR���̷g\�3L�D�+�k*�Z]���ކZ���&�MuB�ֺk�R�vq-Fi���������kKb�8�]npl7�L�֌�hBa��ë���k�
ش.�֋��Z^�И���s����O���=�������m��{�����&�m��������m������z���m�u�[i��Q�e���L3�E�A>��*��"*���H6%��+o�_��!ba-��0f��	)�8��5֑��2͢�:�n8ֳss��oZ5bWF�b�t���Ҟ}x�Hh�rau#�-�j�G6:���E�c��l=��  ������F)v6��f��f�5n�:�ͮ�eV�s2\� ��}���~��O��ݝ�?f�ņa�a(o��ۡ��S�T��,�l��8�$��Ji��?[[LP�w�e�%<�z�Á��l?�,Kѧ�'�PB�
�ͅ�P���֮-��Ƹ=��(Q��k��L�C�h�a����7�>g�R�f�D�MSuݺ���a��6�??:�O���<�/0ˮ���:�����$�D0��z�V^�2ъ*߫���6����D��=��W��.H�E��h�<�y���?=$j��ORج+a��!�}[����O~�Q�V����3lJM�+4�%HBf2�iμ�FM?���ҟ6��:u$���T�~A�<:.�������0022?'���g�9���%����n�]j�Dˬ-���?�㭴����2���n��~��{��^*�!��O�M6}��-,������E�.WV�3MS�Z�]=O܄����?R>0�T��I��<����bJ��w*�3*[X��s�WϚ|�=W<��V�S�ӯ�wls*vs�y��vd2rH-"ٷ5%�G���z��-���G�٪y��Zk��C.Z7$�0ɏ~�WQݥ9Ižio�~q矝m��]G^y��u�[u�R�n�JD
$���=UU��a��:���~>��CJ�o���>V��U�q�lN�ϟ�2��1ͭ�77#�K�,����k*�������ҝN�3���u�^lߩ�UDȪtw��i|_���i�����8r�]�S�7=�����{��y�����4��Ҷ�;L��rRB��MS-?-X4�h�V����[/:�?:ag�x�G�c0g�/]���}_2���F_4�oi�g�eY�r��f#���"ʤ�MX�YL��EC����T�
��`���"��[����E3�YcԵ����jq�E1e]b��m�!/��M����4���<� Kp��q��%%�	�JU�
�X�c�!�"p���|jP���*���'-V���5�!��u/\y�F~��=Vg�/�I�p6�:E��O�m�7��y:�$����GA�`�=\(�4��)�2~�[ߒ?u'��m�A��gM�}��p-��;��a��v������7H�e���%Vڶ�io>|����,�c�(�C,f�b<�J6����$�V�N������=��������Mm�rW}j�}V�e��;�ţ��I���3�m�^���$�0����<É���Q�l���0C�����;���&i�y�p�R�c��+s3o.aj���N����N�����-�GI�_��ru4����?�I"-�,�������Ǐfp1�g�x��3zvv�DY4|��w�UTC�Juپ��_�.`��+��C���a18���/�i2Hy��w�G�Aʣ�I�Jwš�q��f�Z��O����g��Y,3,�׳Ԭ�,�[�*�қ�%��ݺ����sg�tA?%��`~����¡�s�8��#��j��|�;�p�v>�g�w3LdN3���ϙ�Yh�F2�fT�%n��̻��[D=MVY3[U�U����m��~u��uy�^e֝mם���y������d�� �mUTC�(s��U�����8D:��b�c����ba��1K	 N�:�V�GY�	m��}�ؤ}Q��`��_�'9[r��a��u$���p�hgk#&���K�L1\~n��O��G�ͬ�̾��n|~���������a;6��CQ�R����_��c�"���~m�sf�[O8����[i�c�Ǌ<P��<i^&!ʙ���߿F�q�QL��M(BpkDA�/�h�r��#C�{/7]5�i�q�F�m���-��e�Ҝ2�\F�8�F[�#6�` BM��Q$�4Jӫحh����w2�wm���,�O�d��X��l9��0D��G�`��g$�����n��5)�=)�@�j�<���-��d��7F�z�>�I������OB�;6v�����[b�qt��Y�ާ��~�f�a�bO߿�{�5���,9fca*�f��M�G��')�~��1��5H�k?0�~��b��(e�ï8�}�]��I$CL1U�u�����a��\>~�[h���ߧ���������_�d��]>C->a��=\u%�i��(qut�r��{���J��L6�R�jn�r`��NF���=^�SlF_�.��N?ÿT�#fQg�0_ௗǧ��m�
(���{�ի'P����} .z~G����}u��<��_Sϖ�y6�n�|�7ry������������ǗŶǞԖǓɆ��������2�"�J/x�<C<GƐ3����I��I(��/ܓ�<�|�6�-~eyy�-<O<�<�>����mbyyy�<���a�J�_��1�a�ǮW��&��G���O��K���_��/�/�/�������<���q~a�0�'�/��a<�X�m�|��<ǟ/���g���/��^#�����4��#��8�O�x�(�,�VY��޹S�\���~F�_�q��<����8�}r�\O�-�&L<�G����G��[�1�i��O�����|^��/��_4\�ev��̀�Y>x��y�Oɍ1�|a���r��J���!FT���zb���!VɄ��OA|Nڹ6n�i��r�W�.!UϜ���c�������E��U�c���!�ܼ����E���A��u�~7���@O������s%F��~�߻���;���{�Ͷ�o�����zm��www{��6�}������x�ƞ|��:�O�����/2�N���<��$�=��u�w����?�<�����;�~ɻ���������	ƥ��8�&i�;���~��؊)HZ7�9Jͺ1e����u)���	���&�N��&O���L�E���O��� I0DD?C��Xv�!�2BrB�3L�/�ṃ�k�&٣�!�_�b�W]~`�|˯8����|u�3Ǌ<Q�`�v[�!&R�$�HA� ��$�Q�12���*�u/8p���e����0�-���hL�ᥑ%,�`[>�u�i�}�N0���]i�J���������ܳ0��"0<)DC�SڸZ���C��Jfa�-0�Sn���ej���R�Y�z��\Mݮ�[���ǌi�8�+@:I��'c,����Y��!�<Q�ū��u1a�O��9�.[Lj9	�{y�e�-���1)&'_����1_	VL����������y��a��ѐ&5k~�����{zY�N+"�6:<num�O���޶_2vm���I|�>ٛb$�H[��eI����i�� ���՗V�0�B�Ɗ�6�j:H�� !(�B|�k��&TJ��t͛6�=��w7.Qp��DEV"�N�͆�i���_=8��"�M�G�!���pO��Fh~�g�M���&�(r�<��g1��q�}LW~i�3�?z�L����>��>�،�+�8����u��4|��&�Z��N�&,-���i- H�a��?7H��q�Y��өu�hĒa���Y��!�<Q�O��N�"��Uh�N����P�xa�������vw������WO�~a�����!^�_�,�Rr��[ul�E�R#l��u�����P��Uz}I��*�_��R�b�*3�WUE糊!	�<����w�M��&C !�L�$����g��U���:��ϟ�iî��<�̼�m���$���$�.d���=OS���I=Kmd�0Y�-��|m�ĭ��%,=���h'�g����-�(CL:��m+��@!=?e�+�ϣف�Nx#��~/f7����\u��v�۹x����ꏩ#�SGM�j��io��e��n$>�+(u�e�ӎ�UO8�|��m��x��1g�<Q�`�f�m����P*�қIX,���S�;^�neȥ^4�=��6�0�`vq?��-�ĕ��X������M��Yu�Ym��"��%3 ���P�d���dP�~�QF�Ȃ��%��<��*���'���]�-�|���L�4��J�F��h��I�p��~:B�$��?Ǎ,�c�x��f�{�R�_L(0�
n.M��L�M1��f����G����{E"��FҤM
B<�&�v;[MJ�[hJ�[�bM��(n�Yq/UP�8�� jO@�#�*����qB`��+�[{%�z8o�Q�Ç���կGЧ�*��\������`�z+}�b���� A�A�dyJS2���~��+���ڶi=7N6�WȨ�V��묧�U�7H�y�ߗ�����Om��8ا�*����*
E��,YF"�`,DF#b�`,��(+�`!��,S�hZ�YL�x�Db�ʵ|��-�[��֍�q�]eן:��K4�1�(�G�Y�<i2�|E��y8��!�?e���K�h�^�RM��j�tïw��!�Rݮ$������3M�+9��f�l�e.���V����XU��>�i���2���cW���*�!����8*�=,���<1��b�L�C�('%(�����cKl7�S��U���a��]~q���4��Q�Xy�^u��y��:���ܒI">���NCO&��C��Z�`��,D��A����h`�`Q>?#LD/��P2{�a�|�c��Z�-wsr��h��58����^��BP��}m�S4�7�K���j�[Tض_WnT�!�|�3Y�/��ѣ+`�G�L4�"T��Z͙a�ȫ����0�����������Nuu���^u�[y�����^n���I$��i��+(�IVqt�m����OatŔ�Ȯ�u�y��:��S�g>��1L&���~1N�w/L�+S���ӫ����a�!e��)��������$�'�(�K)�O���Y4�J�`�����2!�U�Q�}���6���~8�Y�?��FO�1y���&�͖��k�K���w&\O\y{[�q���ba�<��/�ᑇ�2�ĘK�$xg��ny'�^��b8��I�����yzy~y�y|G�_��2����O_��<���<�1�y�����u����<�-�-���Ǘ]hx���u���@�
|_�_�/�W��~a~a~O=s����y���Z�\e�J����y1��z��~oؗ�<�~y}v矟������'_���~'����K�x�5&G���xs7s���k�x��/��W���bq�7'�1��k�|�O�<��ʎ<�Z��Ki���V�$�/�Kq~|��?'�~����~�(��$jdOu����D}��y�����*W0�z�\�� s?mń͖�+��\N��^W����{���V!����fJ��ݹ�-����+�I!1v*��U���w�S �v�^jߗ�1�V�z�ν�f��e��������Rf�ף�2�qzK[6I�l�����Ǐf���P�e(�|���<q�bpݜ���0����[M�V
���1sqi!���֘�Zs�2�h��^v>L;����<�z�l46wK�Zm���L�lȘŎ�T԰�k�*��
���n�*�M�fe���Վ�s�WF���V�Gy�qb�Ji����6�.k��Lv�΅z�ܥv-��Ҏ)�<��#��͘�tX�^����/nʝ�m��=�Q��5�Q��k5�����u��5��:��ILDC9�C�.
U�P�M��Yk��&<}fŦ�Y[Lf�ͥ�T0��fWcT7�|��\��+������Xm %C��v��LP��m9G[��`X65!v�qu&�co��O-o���,t��	tXi�P͸]V��i�\�������)�	�v/l:��]�X;�����6�P�}�߼z���ww{��y��v�����z<�o�}������m������{�<x1�3K4�1�x�G�`�<o֙�P���l�
�Dr�Z��klqL�L'[.�@`�a)�Pm[Kl�*�$�Q���Kj�5�m����Yuԉlֵ�lq*�Җ���v�̘-�R�ƍ��h�/6:�4�i�qR�QZ45f6��?h Kj�V�8�F
QX�Zn�ri�2��):0���x��z��}�	�"���~�xO!a�N90B�������'(Q��h�h|i�!y���p}�?N�^~f]�|vs��`)�ދ}�������5O����K��m�F�e��ޱ�āsLÒ�j,�b�J�8é|}Lu0�u�򮙬��4�ϛ-��eǜ~|�8u�u�y��l����`q�0���j�
{Ҫ�,�'U����;�N�KJ��7��i��[g�ĩ�����r6���n�MS�3O�e�~]0糋�Ķ?4��$�[*���\�����l�_yݶ�e2ҫ�.n1z�0��Ae�)J�&���8�qx�R��;r�7Yy�$�W�,��RV�-��K~�ܗ�~{���e�\~~y��4��Q�X~y��m��q�����G%3裸H����Q��ӻqi.u�p����i��w�2`��J[�ڷ�?9\BS���T�S�p:����'(�Ga
�H�ݶ���D�hO�-Z�K���4�1����l�ϭ����2�J}��p��<0>��4F�)�><>��~��t�-�2�V��<�n�ےO���t�E�J��Q���8��M?qǍ,�c�H�xf��W��M<0 %SK�W�E?9��{.���ϩ�����\\���j�-D�J��$�bO�EM8���r�\�l���M�;����P��[���'����GV�3�?I�h��k����<��uO�E� ����'Ki��)��'Cߡ'6g��H��l�r��?3L>6-�[E����Y��!����<3b��������R7�]Rn/�i��qv�8�]�Ɏdĭ�6�����ޞ'�*�������}J��o�=�=�HM��&2x�K\[h v�m�В�c0�jj�y�]a�v� �6�f� 	W���&�,�UT�B&;�0��z��{�!.e5'AS4�6��J�DiOR߻�����qy���~K`�w��^]4�)��?o߱k������LS�cȎ�0��\�Z#Z[�$°z����Ƥ����Rхj�oVU>C��=�>SuiK�SLͺ۹��1�r\��C����o��M�"��(��"�EVwm$�f��#����w�Ï�ӭ����8�if��2F~(��g��:1��Γ
"m-U��UD���L�w-���l-�0>00CaO���?�e��h����i�ʵ�g����%I$��8�����?=S�ʪ�D�-ৎN�� �$������la��~���?9�����	�2�F^�\��xtP��ʫ?p�`w��\�8	����ᖝC��_~(?a&���q�4�A�C�^e�[u��ۜcr�^�I�*vo��'��w�nt2|~�3-Ěmڦ�h���H���ID�u�d>���P)Kκ��n�Wct��	�rGMQ�K��=�u
XP�I�0}|e�'�N�\1kF탌e�3M�L3L�8��}�J��w#��uͺu&��)�R���d���I>ե6�6��^q�ϟ�iî�����/:ۭ<���ԩY}⪢���
�|s���zCY��PTjpQ�&~����2jh.�6�*�:=П0ۆX#���S/2��'��[l�TQɐ��<<���Ncե���N��<Vz�d�{�d�A;(Q�;0��jVl>����C�?/mğ0h���e�\~u���h1�c$g�<3Y�vR*�з?������}
>�@F,K�}_wc�)|6�tK����;���$�wL�o�T�8'
�z��me���'�֦LFї_X'����eb9I
hхh�qEM�.�u+�j���%G�  ��1�E!��ȭ�Kà��=0��9�T�qT����O�;��=YaQ���A=JwE�>ޫ+xw>8P����F)t�$�-��8����a�Z�G�~�;-�ᖫdCKo0ǻ��O�dCÎ#�|f֙����+L֮�tt�^CmhYf�]���XS���	��3~-zq��Z�q��Y���?<YF�x�if�:��ï̼�n��uJ}Q^̒E�S�8wC` �|<pr����!��)��6��p��Ѫ�F˧�O�u�sU�J�o9��f�-v���2��xihNv��"�$����g䩳̗�c3JZ�:۳(ᙺ�fQʲ�"/����(��uʸ�d��0��ܻ��L���[j�St�?0��>��I,0Ê=R}tx���?Y���#8gf�2�X2�eH�,���d�2�"F`�h�,g2�I��4e�њ3`�(���2�1�1�qC$�H���2NC�2�1�@�Æ#�Z�:u�&Y~Z�<y�yo �A�@�1���cb2�0c$1�H�h�Y��ǆx�x�O��a�4g�,���$ef�&3�u��t�H�n�i0���#8e���Ȭ"rmO�]y�`.�pJ�qF��=�Z�։��n�o��Xv��������7Wuv`�b�{�D�Dt�v�о}�D��[ƻ<'=��ː�N��e���wNJ����h�w�]S�F��o̪�5�;[��G��k������,���éߏ�N����D�G�dw�K���M�[�j���y(�1zY��YW�ak��̹��{���������m�v������>m���ww{���ͷ�����z�Y�Ɣx��3K4u�u�y��m֞m+�$�H�[����O�&^ܗ��v��;Z�2}�.CH��_D7�̵�)Ѱ4B�I"'pt��gp��J �N��R�vq�HU��f�b�����DF�櫷-��G��k������a\ܙ|�I6Ɋ�1]��Ұ����b��WVѓ��+�"o�O:��J7VZ6��??2������4��Q�Xu�^u�Zy������G�UTC�Cd%4���fgA:���6M
S���?C	C�O�j�f`�V�Z�v���$?�>N?���ST|�d���d�j.<Xy7`����b�:��6x&��=���:󇻩s3[��7C�����uF�owɆM)���;-[e�D��gA��e0�_��~��5M��8�.����Y��!���(�����&>�-k���kk�=����ב�m��̘\�Y/	�;�	� �x���[�"�6w2�J��ۉ�I��M
8���-[��I�5?  ���ƃ}��ė�2Z�fJ�T�t��.1UJ'�O�x�F�
�7�7۞ �DTE���C�$Ǽ8�rJaL'��ɖ���Ϸ%aED>>QQl�dm�jv�Z�1UU��I��Σ�O��9�yZv|��z�Xy���F�S�&���TS>5��C��[�r�da�/�]^\�*k]m�+����.��0��~u�8�if�b�'���<_�-�v����̇��Np�e0>��On}v��.p�>��^e�8LQ�6�F�0DD:'���p����)�%9X3\Nc�0�9	"��D����'��Q3�����GMm����7ON��;;4�(o�|���Þa��~=���t��zl>�x���2)�~������-"�}Ei�<Y��8�if4�:���ζ���݄J�G�$��ؚ}M��/斆��뾗�i�	���GRT�S��DN'Ě]_���C�%$��ր���Y���.cm�J@'��>��
�̸�f���������ik�7M5��:����,�����.���)�<����ƌ|��^1MӋB�O���}MR�W�u��>hc��K0c�H�<xc4�[�����j��xP��Jtp���'�+���1��p��]�i�� ����^��KbZ6~�h�m�ǘ���3F��U����O�e9��9>���pM�'aO���pa�L/�}���e�b��YCA>F�l�irM�Je���Ӵ>�ƕo��Z.z�3M���m�D�Q�f���g4��22FH�f�7A����"Jd���J����zaޡ��u���ߣ'ϋ昊�=3C�%�3ޥ��3��3M��p$�$�R�$җuu#N.���͜#��(���c���s� �[Xl;�x�3s1�׀ёڄBD��P����
r��Z�Ju�g�{���W)E�Ku�ղ~ag��}�Q��'���;0��=)�W���NfdG��$��JtqL=?*˦\>옥�wT��UF)����ꚹ_n�ٛ����Ev�֬S�L���sG$���O���1$n~��%iŚxÏ�i�[�����<½�8����X}��0(u!��,;���ϯ^�A��2�}����J�ӳ�D�~2�VLx~2t�.��yk6~mt�;_at���/�淛�t��.�دIa���}?E(�!�J	�҉�va��|�2�����9M�$�õo~|O��~�:��>;��y���u�_?8Ӯ:�]a�y�\y)��ܒI"�����[G�|�:ܒ��wI�)��>����s6ۢ�?vBĢ~)��~6��9=)��ٺnh�뵍r��T�Tz{�ΟS� �<����	��vu}NfL>f�adq��.�֩�0�WБ�i��	�E��YW���O��0��8�ѐ1�2Fxc4���ݵ��� Ҫ����V6���=N�c����a������8J�WҕP�$FWJ�t���ۓ2e\>��"���6��e?	C��𔉰�O�`|XY���/qƜB+�%��^W��a��$�_+�-�r�L~��6q�K��SL��v�˦JS����IbDV�=�#�0�ǎ��3�3KC,C(e��!�!�J���, ff��i� g#ZZ2�h��0f���1�e���Y#$H���2L��Qc8gaa���ӭ2�<��yZ<��x��c��2�0aC1�2K(c�f�d�1���8��$�ƞp�8њ3��"K1��F2�0c8c4��@��!��,a#I�)2F3ǡ�:څqWj�!BV��Q
�+.�Z���ɭ2�݄z<��\p�92��+W�<�
�l~|�ݚtw��+�!ѻ�*x2��,fKnAc�/���0kq;c��;��P{�b+|��v Epc�P���`<I>h�[�f�;6��!�g`�zfbr;q2�P�&b-����,����D�&����ڴ	��LDt$�2����{ �^��xD�8�N���V'c�eƷ(�'b�]у񖯯�`cu��Z��C
`4�Ja�|W��S*u}Y�
oO
����pfZ��⹚��d�b�?��3���}��R�)��j����ׁ<g#���[˖�`��[w�ľ|���F�F2�b׶J8W�b�7�<�z���_k�md�.L�a>�k�����1���cǔWϹ&Λ�輱��9~[��4��n�9�j��M.�ݠ��.�m��m1��03/W�Z�� eۇ��m�mw`��m�iL7B�[���i�/��̔��V�Zד@�ۙ�]�scxSX�-�\�o��M/�q k�X�l��Q�^�J�t�N��6^�B�v���L���Ҋ��Ľ[�ѷS��� &.�E�9�0���h�al��1=����������{��6�wv����{ޯ6������{��y��ݾ��z� �8�<3�X�#$g�3O�ssT@�SEf)U��Y��h6%��]D��]�\X��MHk���R7�jF�r��blؔ�`ܭ{XA"�c:W�����6햔e��Pt��f:\l� 	6��4�M��C��[�36%;
�f`\̌�Rt~Fta�G|N���*������+�Ul�]��5��j�.��f)���i�ZY�"F��V���wd��GU[������C��d��Y�[y�ɐ�p9��޾��TM-��wTL7��P���'a��x�5��Wξ�!��v�6�#���p�q�Fh�ĜIǎ<i�o�1D�
�Y< �T@��X�$
�J	{N>�S0S2� �a��BIa�p�p�N���qL%��&12uQ2��ʺ|���%�n�$]�����);�q�]�Ŧ\}�Z$[g��0�e�-{1{=�j#4�����w���G���:��Y��[z7�R]�ӯ��9��\?w)s4�F%fcX�?6�f�����Zq��^Ǎ� gq'x񧋅{$��V�$�H�m�a��k`ݺ�X;HYt���iv����+d���,�����K��W����d��l��j5Ju6	����4����x���w t��^��!�&��S�L<�[��O}&i����q�_I+n��n�Lđ��8rԺa����m6���o?:���\u�0�i��������{�e��ٌRbX���D!�"$a�����X��i�C�	��?_�$;m�]�Zc�e�A6�F�K�]^]ؖ�c/Xe�1��3�'P�=
Pd;=�u9�-�D#M��S���$��W�!�-���3O2���`�6l[5�Y��̲r�LG+��1��n����БD·R5[2��a�`�3�3F2N$�4����;���K�ʥD�X��ͣhuv�V�4,�ڑ��Wȥ/L��$
#��l����m��[��XYK�4����SVZk�K[4I�����gL`�y���˷l�;@���+Q*qB��� BW�r6�$���\96�m��	7�/��*�lC�t0���i�91�0�rcG��q�+&�W�B�)���|YŔ�&���X:��M��(����s�E���;:���V��By��5Sӗ��1#��-��Ԙ���2�0���'��k����H��]��A�3L<xg��'qGx�����0I�**2)�W�{UX���x�D�����R�CD]�ʟ`��RH�Fǿ]r��|�,a�5�H�J#��o�á2@��5��O�P��Dq�X�T�U~�Dv����]O�u#u���V��q��{�K�&3�Y�Ј��})K�HR��~|���o�u��:㮰��̾q�yfb�)�Sy��WoJ��v�a�DN��wŖxD�����L�$�$Gc?D�9閭e�N�9)�rn'T�Gx�867ȯ?/����-B���'��Y�ﵥ�:��V�G)�~�x���G�:!���g��&?}���[t�1H�<��>q��81��0c$�N(�O4�!j\j����V"S�au��|tt'?N�XQ0O5��9qpU\�@EI��B3D~������<���)�h⪄G��P�!6׬+�7�6��	�p�2"�m�G%2N��|q�!}���/Yh��i"ѲSk��e`�t�~? ��*gD�iܱ�'*|�����e��>q�]yǛ�8��8�Ǎ<\���
n��\H�(�t��K�S�D꣸��Zeϖ����j�7�W�}�\Se�Yfõ���6z��)��X�a1�� �/� 8�f(�}X�F`e��[�k-9��DFm"�&:�O�#��0�=NU���/s��0amD~��{}��m4�0��l�t��g㢜�r����>%�U�x'�w�t�'B.~�[q��w;��pM�Uu�vQ ��|���q���Y(��Q��鰗@m��H)���b�`�:�SO��D��La�Z�H�.���I�q�>a��p��x��d�I�i�ƞ3 �����o��V"}�a�"'�<��C)�"tiМ��'G���.70��:�8�烙�4�Dq�a��� ��C��4��SN(���!1˒ԙ�s�F��i�ҥg��Wi���+��[B����UQ�n�h�a�*�Xa����9�/����Ǐ�8c?1�#�h�i`�@�D���f`�"���X�33Fp�i� g21-4f���+Y$b�1�1�2��d�@��!�C6&2�1��4L�((duh�N�h�(��<y�ydx��xG��1�ьc(C��1�2K(c��4b8c���8��4�3�q��ќh�0�FI�11�P�Y�gn6ۦ�Ӭ��GQ:�0�2�#��R���VDvM��i��Z�{$�qw4#J�|��}�1ݚs�O��J��X�6�|9� �-���~�B藅��hx�z�p����LkO�jl�N����B��U�f�7wǷ?w�}�)�����VjR��b���7.RCD	���RW�,�[%j�j��H�C^(�H��뺮��N
�
X�}�l�&����#;f��Es�����ϻ��{���������{���������{���m����wz�x����3ƞ0c$�N(�O4���$����^�}�':�q�Gȁ�3R4�4��g�)�u�\\Í�X6���9�����-�Lb�J���
D
�4A��� Z�sQm������3La2`�/o6�#H�F��K�4�µ�%�#NR"1��D�MJn�;$Jf�H����x�����~?1��<X�IĜQƼ�2�&��ʊ���J��<�r"-��"2��金�J�{��	�.��d�\�J��- ����֦�}�o?"���%��C&�q���T����4eU�u�)O����{7/�m�3K�h��sY��Ȣo�Тrz|w�ݵ߷� ��8�h��g�<X�IĜQƞ<i�5�#R�t]U]ZU�JKW�_b�F���32luq��&ĹV��)a+�T�����Z�W1�U��'��l��b4�6���W���S���72��֭�HUl$U )�Jޗᐘ��m�7K�����cBGU�i���ti�	��"���t��%r�e�r���+f��!���KlzNOǟ�]:���P���m����M�N������8S�'�O���Je�ngQ�Ӹ3��'�'���f����r�1��$��DԎB�JC��V&�#����7�h�A;���v�k�g�F�,�ǎ��O1�q/�|��8�T�W��R��UH�L2La�]b�׵U���������� �������4O;~[V)�|��k�2�6qiojOS�8Q��s�Ks�S5ҾG�;���U��h�*��O�m)h�>�F�~=��ѰG��x�ynY��5.&Z\4��vx~�8%�wȟ�5�é�:���D�����܇s�A�x��8��g�<X�IĜe�<�Ϫ���ܒIQ��+^�~a�eVqLS�)M�3Y0�5MS��\I;L>|«uXE�4��q;����`Ҡ�J
r";M3]F���+�a��7�n��i�a%M2�<����ݿ��2���R����[4��k>c�-4q�|#��ӌ(���p�x�ź�����<�3*LJ�RI%DX����ggLs����DNY��\�W�?R&�qN!XՓ�<��M5,�ۢU�C߿�{��&�����~i���'W/�Oֶ��?=L2��Fj���	(�oӸ���l?C݃C�&��l�/ٗ�ff�w���~�\���m����+���	MR92ˬ��矎�x����qGx��^ԶR�)���M����rB{ҳ>D�n�D�,ƨ8e�0��.4b!�%��B�ti���L���;�s��'� q	S8�C�e�s��T�ه6YU���T���z�A��N��~I�2"'G�v��Zal�~4�N� �'$�5KCh���K�^�4���Yu�O��b]��M�G��&	�<���8'�U�k��2�4�SH�s�.�=�Q�K�˸f��j:3��x�C��UUue�|��.._��V�->t��g�<X�H�8���O���Ub!��1(����J�"��0�a��~H�
��C��*����	�Ȫ�a�F�GߗV�HB����e��BZ�H�,�'�wr2;IL����D����ih�L0�M���2�n:�c<xgg�Oxd���8јx�go
��G4�ea���U��Q{��ᖩ�r���_��~�zI��"�QK^J"!��04J~<�W)U.f6��.��k҅�Ԗ�5����q{
�Í�i�r�rm���*�F�&)��橃(���ؑ�z��/�|u?Nx����v���8`����)NJ�Z���4㎼��^q���qG39��B���K䍣�z�w�d�SՆ��֘������ϧGc�� ��hmPe�g�%�cb��;����Yمϧ�Ò���z�+�]�T]l�qk�)l�=���Z�C��L�XDYT���r���;O��Ә��yà�ra�N	���'�Bڛn��kF��,��Vt��<��<3�g2M0e2P�Q�2F@!��I#�$3	���8њ2�h���X�"�@�1���d�#�H�� c(��fc4�O��n�:��0�֍e[G�<����u�]u�]8g�1�@�P�,����5���3�8��8�f�3�4f��L��1�iH�Qcf�1��д@��!�2�$c�$d�ejK��
EWj�[��#�ft���]��;����b�1Y�!�GI/�&'Oz�q����B}���o�$ʯ��T�{-��ty�����i�ů�|W�ɹ���C"��!�l�k2�frQ����〇TS��S��wt��byj�"g�#F<�bui"�r#F�"C���^7���O��w���Iܙ���-�ї��Sy�3�<o�����]}],RI֯#��!��~־���'������K+�Z�1�`wf��mS~�<â�izv�4��*�zK�۔|�Xh獋��M�2��q_{���>I�b�{�m��'�4R�8��]=�=�+lGN��{��F�S �ETT�q�Q�m�4c���.ܯ��!�Da��v����۱4l�v��UL�gf�7�}���ۑu��[[�XX�{Gi��/��=���g�"�Xe�V�4��ō�)i4�A�ID�YH�<<h�Kx-��+(^���'���Bի5�qUn�l�%��b[�QS]]T��:�ͷj��Y�6+��b��l\ap�{ks�)�\2�%W�OԾ��������������{�ǻ���~���{��ww}����{�ǻ�������<iǏ8c<i����qG3���w�؈2�A�Ʃk��Ze�ޔ���mmF�5��hե���2��
���uk�&��q�k��Z�WD�kH9�Θ)��V��]��h������� q	���|�]+tf����c,e��6	b���j�����%Є"M ֖�0��9���$�30(����YHjI�N	��/��b�66�-iI��l:�o�6�.��J������Dn�~�'��0}�����1Qq7.|p��̪~�]��0G��{~E�ֹ����<�g,��~<~?1�4�g�H�8��<:=3�h��X	檬Fxl�վԍ���"y�n��jgL��fT�����1��.�O��u�n�-��<21Q���oftpd�9OI����F��z�ejK2�]�rP�.�VXF�����%o�9R"'찔���0�t���Î�c�Oxd���8јx�}3�*�D�w�_���5����h��ʓ�����~m���P�ϻ�"g2��Eh�^171)4t�r��t-��~|��Io��|������UH�#�4�V�O�e���ɚ��g�Gb�ȣ/��T�����=��os�r��M���q�1�3��3�(��'q�����YG����U��L3�g!x���F�Ϻ_���Nd��W^K�z��b=0�/|��ĭ%;����ѺB�RV3Ȝ��Ncs+�	��~�n5�?)�����?���zC���U)�ϴiDAA>����r΃�?yNNЬ��Q/����8��4c<1��Ǌ<2FI�h�<n5iS0��ZQ�Y*x���k���O�Km}X��k�������Q�7��0��#A��.U��E�5p�YFZ�.#ַY���e�&�]���~_z+��/�6Ɨ���̈�'f` �6��Ͷ���Oj4_Fq�%��>��Í��9P���?����3y"'aC�u0���Z�Z���}�HĮ�q�Ѫ��.����+��n#Ov��J�U��\Y4��p�l�(�!J'��̭F�~Ԯ�]h �=��	Ra���-/&�?x?a���߀�.�E���{R��~�ьg�1�8�O:ì>|ӎ��+V�I��I$�Mg�d��ZhQ?zsƢ��3F�á?T��;<>��!ПQ��~�2̿E;:;("p�thw�Y���g�G(�W5+��Yt����u�kK�?�i��S�x�Ϧ�8
w;�:/~��Q+~���]�b�Ho�9N����y���x��#$�4f8�}��f4*X檬D���S�N��,UZ9�^�D]%0ΛG�7_P9���������ͯ..i�/��Ղ7���^u�6S�0DO�ɢa�
��ta�	�0�~�8�WԷ��H�[o0I�hO�䵫�gt��O��0��Z�-�?V��1O0�ξqǞy�]x��#$�4f0�*���b�QA��U��g����<;� �4�N@��gBh�_��扶[]��v&c�Q,�����g�5G�i��\_cK�wnSm��"9o��j�����S_9\��:q�0ۙ��h�-)4�L�D}H���ɤz�Ju��`)��xјqǏc<q���yyb��j��=����t����ڜ,-�=� j��,����Z�if��,�,�R����C2�HK��̰�X�)����ϴX1���Դ���&��aj����31 �],�����&�ml�� 8!]̍�3庺fgMn%f��l4]5�U�����^�����V��.�����b�Dql=KdO�gs��t���B`�)��~��Z_���G�WN-�����9c?�|��"����U�q�[i�7Yb}ϠY���#+�U*�5���+��i(��ag��NO��xQ�B��4��q�<1��Ǌ<x��qŚ3Y	+��A/���b%��bQ8u�{�y��U�b�V��mR�D�T��J�.8�#�4�ՄF)��"J���"�ߡЈz|v}Âo�]uv������aZ�ʣ��0p@;�������m��%���4�}��v-"��+FYW_��Q>���{���24d�q�1�p�(��`�CF�P�h�"��,d2�h���q�4g�KFh�7Ec,Ec�&1�e�C� "?��d�e1�f�f���@1���Ӧ]hѦ�h��ǫ�xG�<#Čc�1�2D0`�#2�IEc0cƌ�1��Ǎ8�ǎ<i�Op�,ј3�0f@�!�`�,c0�1�ach�!�c!�I�$d�1�1���_�TBWZ!H�"vO�D�^�d�@͜�W�st�z��oK���a )u�5L!,Rg>l��ܗ1�kLch�=j�r�`��e��k8�mD�E����Z��֭��Jy\L�j��U�����D���s%V��Ҭ2j�V93$���I+��^n���{����{��������{��������{����{wwww���x�ǎ<3ǆ1�x�G�2N8��a�|�$���S�xs�˘�(�dDI���pOO�CO޽l��8�Z��k`^3Cg�l<t^��,��~�ӣ����@�S�S���%��_��S�_�i���R^�i���1�&\�gB'�I���8&MZ{>᫯<���??8��κ�<��0�Y�0��TML{I/��4�蓮�#h�2��/�V�R>G���"�k[�	�2:'z3�YOM�f�U�ڽɂXr���֩�â`�1���a����F<���=I��)[Dx��0����	܆d;=�á<�4�O�1�pOfO�2��o>q��:��y��$d�qg���,ۤ�!0.<2Q�A�e�����tQU���6,{�[�,��h%"���_k�Kc�ݢՈ⹁b���˫IH�M��	�gM��GK3�Mr����mz��g� q3�5H��T�����nf�v�n3\���ӂy��R���Km�?3�9��Z=_�6�-�≰F�����s7�����E�����"S���:T��О��������a�m�M��Wb��x����'9�#�p֍̙*[n���5�2�jY��]t G��+�B�	2��ɉUZly����4��<3�i�Ğ<H�8����~��e3��0\�Z�ޕV"6t���H��Ҥ��˺{4�h�+ҔXH���R#%�QB�&�/\�ù����Z�'f	��6	SD��^5+E=�'�da����(��5��󪪎�ʣ�9e�۹&�zt'd�N�Ц��H�����}�>k��tJKqR�n�w��aמyǝy�θ��<����O�m���;�$��U~[�����;��)L�����
fc��l���^�؞~�?w;ò���E�Ҫ��B��BKÒ'%3mc�`�z~�
~?�D��'�_N�9B�QR�U_��b4�j�L\�j�(�$�q�u�ѾV����������y��q�-?8��ξuǞa�y�Ϛ|�o8W�Ķ�T!U���991��I��o��SO�l�	��V�9D}�u/�3�G^�,�c��,�q!!+ͨ��[(яv�wLӵո��N���%��W\]|�2�F�D!|2��)S4���<L���ҏА�uZG��=Y4��3ULu��]q�B�|����κ��\t�ǉ<x�Ĝqg�-[Λ%\Ii��=�=n���<���D�:��kmV�{Kem���{�#+�	I�3(���w{g��$&z�9�[UN�׹�����XA��H�!3[p�M�\�*n�%�ݶ���55�av���7�� q	g�������F���m&�ݝP�(��I����ҋ�-Uy�V�Z�u�R�J�zx'g��a�U����{�%����8��o>SE�"/�)���T]u��ZbHC�J�:�5�u.�ϛ6q���~���Z�]n�KX�5���wt=[:�;�w=>4<�tz؁(P�H�Ɣ3�8g�4��O<��>|��[}�$S7%Ԃ$�D��*,Xɏ��pS�t_�Z�gł�>�&d�Uq�� �2�RD~ϒ7^�7�Z>n�l�,���gGx��Q�h�fé>U�wW�9W��K���"��qD�w��ʍi����"��8!�j��"�L	o�i��L;�qCnh"y��$t���gB����<P�p�xc4f�<I�Ğa��<��Y���R^=�U)+���\�~o��X�4��������Jv�'��Y�3���ZT̻lv%hgo��ɧ��Ϙ����<�=V�LJ��H�m�V�ؗ.LS��k<����fSf
�"XP����$�e�.��<��<��0��4���Ȫ$IURTE�+7�����/�M��߲±N�t��8�����r~,Em�GT-��ḽ0�W�*0��.���+͘�5L}V+�K6�I)m��;�&*���O��%����H�&�R��$���;�7wt��I��&:&i`��{�8$�	�o�HI$�Eh��y��_A�q����rzŉfKE.�"ⰲq�w���"s�#��H��X�? ]T!	HEBQ�%!�*B����B*�AD?P�ȂA� �D� �!*����B�	UBRP�HEBQ��D��	` �JBRBR	HB��J!%!	HB��� Ȁ2 "�"B!*��P���"	H$%�� JB��A!	UB���D% ��%!)B�!JA*�R	
��R!"��*R)��"�(�!(�B���!*�@� ��� �D`�#" ��A�����A""H�$�#FD@F��dD� #H"DdD�DH�H����	���$��"�H$F$FDH#H����#AB"DdD�AdD�ȉ�FD��`#"$FDADF"DdDFDD`�$�"A"#��F�A� ��F"� �����#D�DD`���C�$�EF"�F0H �`���1�����0B1FD��#H�`�#`�A`$FDD`"#"0`"$��b$H0D� �##D`�#A��H$FDA� ����
$����F	FDA��� �2"#DdD�AdD��A""� �FD`#"$F�"2$#H�D��� �#A��2"�FD��ȉ�F�2"$F"Ȍb$FD`�H���dF����T�Ȍ��#H�"2"DdH2�A�Ȉ##a�F2"DdD�DH�� �"2"DdD�� ���F��"2"DdH$F #A�H0�0D�� ���A�FD@F�0`�$�!b"0DdH$� ## �@F��K"2����dD�" #D@F�2"Ȑ`��0�b$FD�ȉ�������0� �$AA�
H��@b""HJ���`��H�H+���H#�.(��*�
�PT�H�ĄD$`����D%R�B�|�V$�
�H� �)����cY��"���BT!	HD�RFF �0A(b2! �D �*BȀ�A�dA�� dA 1A���HP���!*�(�B!)T-��!)�%!J�!)Ab����%!*�)BRJ�B���!	HB���"��BQBUBUB@�dA��DH�A�DA�A��"�2 �2!D"�"�Ȃ �B*��"��*T!	U��!	U��"� �dA�	`�2%B���"��JB1��  Ȃ2 ��D!1�2!�(JB*���JB!$A` �A�@��%!	D!	UBR�D%B!)	D%!�B�T"��JB��BR���JB!*��*!%B!	HD!	D"�R���Qd�"�(�!	D"�)
�A)�JB!JB�T��!*�E!%!	UB�	HB�	UBUB!
��B!*P�BR
D%B�B*	UBRB�!D%T%��T%!	H���B��!*��P�������D%!JB!R�	U�!)��"����!��J�D%!%T"��
�%!�JBUBR!P��!BR��
�% ���!!%B�f3ad%!��!	HB��B!*�R��B	U
�D%!�� ��BR�	U	H!	HD%B%!J�B��%B�PB�*�RT"��"	HB��P���%!%!J!P��"�	D"�BT!
��!)	HJ�DdAda��H�!J�D%��B�! �"�H�� ��0AdAdA#` Ȃ ȃ" � ȄADDB��%T!
�BJ�JH�"	dA#"	dA"� �" �� Ȃ0dA"�!R���!*��"���BP�%!���!	P�)*�JBR�T%T%B ��A� �"� Ȃ 1A�`�" Ȃ2�	U	D*�B�$��D# �0A��!*P��)�D"���E!Q	HB��%B��!*�P�n�D%!���"��*R�D%AJ�BUB�	HD��J�B)�J�BR�T"��%B��D%B!)�����BR��"�"��J��"	HTBT!	HD%B*�T!	HD%B��BB`� � �A�	b�J� ��BR�$A��@A��0A"���т�E��r_Z���4�)�@g�' �`�(2
�!$�|��ho�^̰��c�O����?e�?(˨�7{�g�����tǬnczB�k�W��,,'���d��k=/�e�^�`�U���.2�;����5��o6w9�F�E�u��ry �y���{����!��E��@�
����?l���8��$0Ա(R������.�����>�!yϬ�j�bz�Ef�>��G�脐/J��a�7z�ѼJ�5f:b��LJJO:c��i�k�c���a<��&�-�t/��@�����{�l
wP� ;,Pr(��Dl@DjT9�Fؗx�(��a���U��oa��oZ/���7�:`
��"(���� B��
�����Pc�x0tr|��Z�����qpi��5��\
(?�e�h}�@���!��� �EN-�˱�߇�q}7��q"y�r�Pb!��d#�?w��p�y����'������[^�ŧT�1<��AQ�=3_gB�z��xN�M�\/^�6� �q8��"�<��X�,���뢭`8�/C3��crb^��`�R���m({z��!		�ؒS����Y�  ���Ł�l�z7�C+��)(��м0D�L��(�cb6�qe�b����E�O`�(�J���$'O~j3�zpAQ����ܛ����B��>�Vz�flO^�E�����T�=aŤ�<::���AO��%?W�}��`�%���;
@ԩ�X^�JH"�8�^N\O����(�[Y����&���<FK�$rI�HB������I.(([�j�����@::��P�l�C^w�c��R��^�Y�� �(��p�X�!*'2k�@v���܂��Xw@�o�d䜊e�Ey�HV8���:#ƙ
k�;��b�� ��q �����	��2hmK��������	�IÙ�8^��i]<iT!d��M5&?�����"�(HW��X 