BZh91AY&SY���D��_�pq���"� ����bA�               ��RJ�Rl�T%*�Rm��QR��)
�J���AIJ��U$���J���ED��4ڪM���R�J���J��F�)R�U(�B��J�Д�*�JJ�����(�*�� ���@�����T�$�AD�@ +���mH
'�6R'F�p���4�����]�MdW Z�%IJ,��L�!j�JRR��"H�A*Nڊ �O����EAV�`z"%)�x�k}C�t�N��wG:wt��]�qۻ�u�:�ƛ79S��wn-k��Jڭj���m��5��j�M�i�QNà�*�֚���ZA$�M�T�w�υ*%�^��@R�����q*R�[��oT�T���"�ƕK÷	
�ܜ�N�n��(�T+�g@*�m�v��4k�RUڦ�R*���@|�ZhTޱ|iJ�IwK� *%���Z@T�-��zގ�P+��o3��W1Ҕ$^��zP]׸5@����m����5'��wT�� ��()IU]�I ���JR�@{��悊TW�v���P��G'^��
����瞀^��n5�P�����n��B������UTy��ި
���z��
=]�h�U��	P�P)D��)%���JQJ{��� 	OwT{j�=:��=��T�������=((���=w��D���@䠣z;��ƪ�N⏽�*�H�ϸ�U[�R*���*�U�}򔔥 ;���� Q�pQUZ4n�燎���: �QJ�L 9\p(�`h�;\�: g��z �*�ꕩJ�6jM�>�Kl�| o� �q� ��0� Y$`4Z��@;���W���gP Q���]�� 'ZQJU[_|��*@w�� u;�` ��Y��t�
�]�� ev9 tv���P	;�8 4w�: ]sE �+�J�eB��P�B�A_}J�)@7�π���t4Ɓ@w��h�X��g`�@�@n� ���!�P��; �T7�R��@�{� m�@uɳ� �p�mv� �4��v��,�3]p f��@� �          ���)T�L��042"��Ĕ�H �    D�AIR� �     jxBi(��ꞣ@     $�JE3*��14�&Fѡ�i�*C��Q!OЍ����iF�4m	���O����~���*���Z�=���7����>���h9�m�:�����*�Y��R����EO�
(*��EU��'�����Պ��TD`���UϥAW���?�
( ��߷�O�p���8��c��q���c�q�c�q�|y�c3�8�1�c�3�N<1��1�c1�g��1�c8�3�c����1�c�c�n��zc�q�c1�blc�1�g�q�c�|lc��1���1��q��c�<c��q��xc1��3��8�18��1�g�q�Ƿ�1���1��8�1��Lc8�3�c8�1�c8ݱ�c=1���3�c8�c8�3�c�1���7�c<c�1�g�1�ǎ1��8�3����m��1�c8�1�c8�1�t���{c�q�g�1�ǎ1�c�3�c�1��c�c�3�c8�18��1�g�1�n��zc��8�1�c8�1�c8�lg�1��1�g�1�c�q�c�1���c�1�g�q�c�ǎ3��1���1�N<q�g�1�g�1���:c�c�1�i�g�1�g�q�g�8�3�8�1�c8�1��0c�3��cLc61�����8�3�c8�8�3��8�3�c8�0c8���8Ɍ����0��*x�>20�0tȘȸʘ�=��2�2�0�02�8�<`eaeaaL`a\a8���(� � ����8�8�8�8ǌ	��D��Q��A������A�A�A�A�T�A���^�CS�D�������R`q�q�q�q�q�1�q�1�q�q�q���� �*c�"c
c*c"c � �0�0�2�0�l#��)��������0��8��ʘ�8���8��8�a����T�q�q�1�q�q�<d1�x��8�8�8�8�8Ș��@��A�D�T�1�1�q�1�q����"c(��*cc"c � �/CS�D�T���D�P��������)����#�	3���.2�020�2&0�2�0�2���q�1�1�q�1�1�q�1�1�q�1�;a�D��1�1�q�eaLaLaL`N60�0�2�2��#�	������/�&0�GG�����q�q�1�1�1���� �
c"c�*c �(�0�ʘʘ�8�8�8�8��(c �
t�8�8ʘʘ�3�,�q�q�1�q�1�1�1�q�1�q�;a�A�T�dLad\aeddLa0ʘ�8�8�>2&0�0�0�2�n<��1�q�1�q�q�q�1�ddLd\d\a`\a`I��Q��T�Q�1�q�aC^�1�q�d�1�d:d\` �A�q�q�q�q�q�<e��(� �0!��c Ɍ�2�20�22.00�Q!28¸�8¸�8ȸ�8�8ʘ����(�
c �ȸ�8ȸ�8�<c�`0�0����)���� c/CWSWG����Q��q�q�zaLeaLd`WI�q�q��1�g�g8��c8�1���M���l�8�0c8�611�c8�3�c1�c61����c8�1�c3��0cόc8�1�c63�1�61��0x�3��g�|c1�g��3��3�c8�3�63�c8�1�c8�7M�c8�l��3��8��8�1����c8�lg�q��q�c�c�q�g�q�lfg�q�g�1�q�g�c1�g�ǎ1���3�c<xc8�4�1�8�3��8�3�cv�1�t�3�c���1��1��&0cLc&3��8�3�cq�g�1�1�g�q���1�c�3�c�Tc��{c1��c�q�1�c�q�c1�c�ǆ3��1��3�c<xc8��ǌ�8�=<q�g���3�c8�64���8�0c8�3�����1���1�g��pg�q�`�q�c1�n�1���1��q�lfg�q��q�`�q�c�1�g�q�c�q�cc�c�1��1�c�1�g�g�Ln��:g�8�3���x��3��3�c�1�1�c�1���3�c�63�1�c�q�c�lc��q���q�c�1�g�c�<g�q�c�c�c��c8�0cM�c8�3�c8Ɍq��g��q��;q�c9��9<��Ӽ2��g���Y���]���qG�"�]d�q�5.�un��y&��5�EՀ1R,���C��<z��j�WRkg����Ǭ���0�I�ih&���;@���h丵	�#+cmL���I���I�R�h�P�De2�,|�v4�Mx(
�m�Y�D�0n%WIc�y5�Yq�Y�]cUh�/�A�+�0*�:�O�vV��x�J�%�b�iPP�&��۽�`-�0ܚL�kA*���-]]���,ayI�0��RƶҶ�ѲT�{J���di��(�����Լ�&�&�ǷY"�R��c3]�d7m�L��2{��]��sRʷ���i�F�d���JUpE1ko�6�aB�u�HR�b TZv�$�yf�IM�2�J`�h�w�@�
�cŪ�"�f�b�0����)Gv.���HV��:N�T�Es]Ս;tU�f���ĩ��Kb�J��B���dn�7m��F+N�l�e���,�'X*Ԛ��^b��2��\�0�r�T�6�0�q�������Ѳ��MX֎5�VkT�Pm�"	�� lŲ���1�[�JZ���ĭ��,:��������e��lj����i�Y�|��4��^3�)�aҼ%h�/t����K9x��f�U�Z�v0����U�de���cl���5��J�z��R���&�M�K�t�
�,)�rALV*A�fNY������xr6+@�f%uw�w��-�6R����Z[r�1j<���wWw�dAe��e�C�w�X�ٺ#v1�!��Q�4���y�����.4�0Q�m���0�!�lku�-�c�k�a���]Ye����QN�����C`�g̵*����F`J �)����iv�&e-SX�p�ƽ�4ى�[N��E���-��qP�(м�W�w�Dr�Jt��%VhʑV0M��Ù�
-�BT�ؘ"�e[�Q�f����AQS[�,÷+d��2��cl֥��0?Az� R�t��&M]B��B���V ��y�0��SǙ�j��`��	����+&-ܐ��f��)��̩���w��ìӎ�S�i+�i&�`+.����Vlօ'��њ٤�6wefm!Es���fҔ@��>-	B���q\ɕy�Ub��cv��.΁Es֡+e����7Q�b�����K-2Y6m�e �X�k]�­d��G5����idA���B��B��̱(nb�+k�7H5�X�`�5X�*ܖ�Jdf�����*i�jȲ��ৡ<��+
��
����p����L�&5�n�#�
�����%)*�.��-�Ҋ��vdy�������6؈�t;�r����q@�H��Ԩ�UtȬ;�3\L�2�ڡ�QZ�z�d(4Y�աӤ�F�b�9����1ȫK�:gI�Al���w	NTi%7TR�[�Y�>K.R?+�y�Z;#��2��ZCi��ݸ�C��[U�f��V+�fU]��i#u.�TL2�ض�Rn�e'��h�9qJ1����ǹxsꎆ��*ڼj�5��ej�ˬ)6�֊��A��ʷ�U��gb�%��{Aj��)��2*�$wx!�o/#T+D�h��-� ��`J�u\$���kP�r�����˴�Q*�"+jlRmc��oE{bK2�XԬlXe�vsы��{�:��� ���5�5QFֳH
ӻRfk��l�2�'fi�e�;h]^S����)gE�{,e1WmD��A�6S����m��ݕ!W1�茌�#b=�1Vj\�&��P����ѩ���f쳕�>�D��+|r����)�Y5�^hA˖2R��KN��2
�ba�:�R�Bi�I���+8�R�V�.�R(�ARdhr)f��J�	Tv�J�'�]�l�:�S��T�v��V#@і͙���w%����	K9f!?>�˔�kM���fG˚.�n�&UAS���y���eG&�:h;���]�n���U�8�Pcc�N��2�&��k�*��M�FB�։j���v��&]^�3/��¥�����uvn�F��f�b@�@n�=%B�P޷tV��N:��p���B�J�E��)h�VuRf�Rǫ1�^��@����é7��Z���ӡ��V�'��$9g"��=�i�T��I��jb�Jff<� �KU���1"��Ka�1��.�:x�ݐ����
��r����ca����jɳ��.��l��9M�1+u�ۚp�,%�8E�PF��܂�L$۩�n���]�h��c�]�u+*��DόTe�9	���7Q8��o�.�u�i��?&/083n�͸��#�I�%��n`�5�yW�k©\�(��l��+ڗm�� ����Z�Z��ND�m�ƅ���mK@��(XFy�>cH,67�<�ʡ��e��V #�0�\0搁a�@��V�3w\��h�����j��z�ݪH�6����`ڑ�<�՜�*e�lͫ���w�]��u�X�P��"|s���Fl(i9*�]�F*u�:�U�RE����"�Ž�9W��%5^�50]�u�1��4���qMT�3f
��J���\M���Q5�IG�e=���]�f�3A��zj�T*M�*��x[SZ�R�h�Fטqd(*�Zv���l�M�Zos�CsB���!L.<F����m�V��Y���˫��Yf�%�F��ܥ�4?�m��;iaH�˵6%J`�1�*�Y��X^SX0�Y�v��06F�bJ������0d��h(l<�7B�a�ӥFЇ
���ī��.�^���V�S-n�f��m�D:��t�U�"
�Z0�tM�p-3�[Bf�*Q��z�	�G	2E��ѩh�����Ћ6"M+r��L8X�G�4Έw�7M�E�nl���%���1����*ʉ
oe;�P�n�8�&�ɩl5�`�*-�� ̅��G��b�m-�/A��(�'$M��ŀ�s2D���+�wI�N�W�m 7<e'D
4n������~QFPWb�q���^��Q�ؒ�*v��XQږ.��k�땗�3R &�AǤD)���	�Y[p��mn�%k�����b7xZ��؊ט��W5Ga�@�pme�ҩ�A*tE ���*�I[�9��m�&Ԛ�c)e�9y����&"]X�B�n1���Ӵ�f�h)��t(�9�Ǥ�YVv5`��}��	�����dB��J�Rme��&ռ��рD)m��Rm���6�I/M^�)�v���ߛkURk�ˠiL�*R�*�J�&�k2�Kǁ0F^��y���V8�Ri ����qn�#M��ndz,e�c�%�,��.Vi.�ONޑ[�*��5xu\�=�b���[�q�ły^��9n�))�/@�%�{�`Vc�j�sm�[�(ę��5���DR���"�M�
�^C�tˣ�{i<�X�V��ї�7.;�i�� ��%D�o՛�1vr��sqe�&��u#6d� wW1��(�)�[2�X��̀[L�[@� CK2�yr%���h�6�����Y�k�X:pE9mk���sn�ӊ6�a�IՕ�a�gp�,`�۵qfû�s4����+��������N�Ac�m�N��y(��tئ��nQ��w����rVf%Ѧ���2X��ڍM�u������l�B8������Mʺɉ%[��r�#SJylJ��r���	�VشOa[Ko,�lIt2P�y�z�`Nə�*uu�7�������'n<����2�m�*Nd�n�ahز�[	�L�S����������_\��X�;]��ѽ+r�LX�Q�/]�e�ܙ�+t��k%�Ȃ2f�f諩�s%�F��oVI��B�z�e�ob�zH����7�YlO�
�S���X�B�)y%� ̸�wu�j]��v�ԭ/,��4A	")��5)a۸e��[a��JX�ZW`�
V��{�U����
����-���d�J�,]�Nܳ�	�މ�-���� \L�QS4=MZܥ��&�)?uՔ6�N�ⷖݼ-����[},���ӗ�fB�E�{Kt;�35�u��R�)�*��C�<�M����*��cOrz�ƴ!#��wD帩ǘ�ӧ�n���.��-o�!�j;u<qE�iA���Y�*F�V�`P'F,�Dѳ$�bZ�n�����C���q7m�ܺU3N�B��Ҽ����H�)��Q^���,�pڵ5n���Х��6SnÅ�g,�ʁ�ز��2��w�Q�Z$�(�*VY���=���{";4���#p�۔��5u*fkr�S�q�-��#u��E�V$�� Ocܰoi�*��kul�S(�IV4�v#��d8P�Ira-Jә�[)֓n��J�3HHFm�3$Z��x�m1kxe�2`&���-*,'l��6��/IJ6�f$Yǰ2kp,�"�!S��W$�X��i��y�+��0���ɷe42˂,Pl	ON�9�����̊ �*�,����R���)�RM�-!�n#o)(���5�&�GeE���+]��Sc��s0�*�;�n��7���:��je�ǩV�dbڴ\��G]�m��PlwAK��Q�݇�lUD؁�V	�dRj�1��YH�!�u�V�����IY�m	���dywL��Z:��%�MO
��������B��Eĭ�k��;X�ж //.�LVȱS�f��N��8��`۟\�֞І�	��70P��d�pe�e4�&,�W�f$�¤L��PM�
���2��j�6���T�F���NQ�07te�/3BR�̢��.-A�)���TE��4���<�K�V�W�$	�^j5�k�<%��m;�w�������i�v2��h餶l�$kvh[JI.hY�:��u�G�wj�Q���a��9nKD� �b�B$j��i0n��h� ��l�9`ѳg��R�Ir��c'���攪Z�KF�[�a���Uy��%$�N6FTlʼN��Ȋ4\VŹl+��$��X�J�����wn�1��[@$�r���V�qM�w�m��L���Ϯ�V�hF���,V4�Zpn@�!i�7t���#`��	(��d�O��P�,Њڊ�	�J6�X���˦���k$3Z;�{HP�^�*PՕ3 �������]9wB��p��]IH�Ğ)�K��kD32�z�����ĕm�ܶb�������Y�F�^
���N���QxE+���D��%�I�i��M2���5�#�!ͦ�5�U���L���d���>;��d5�����P�)�y�R[��UҗP(��O�@x�(�h��$����iw����K�Z����FU��=)�b�qi���Q2�P�ᏹL5�����=���������N#�&J��f�/-U���ͽ�k��6��2��QlR(T�wۉnix���7�E���1+�@�
���&V��yj��'{�f��Ss�O�;���DI��%mjش�+��`�ب]��Ԧu�~{%A�i���[`Q��+ղƳZ�DO�E�E�����$�2��q���Cu^�}f��*G�.��J荽��Mø�tD3�f�xi��	�<�+ ����I�*Adt�X�F�kD�2\���-+ �Gt���U���RSm��yM.��y�ue��ZK{�vo!I�[/$�/�eQ'��0���9@b4f۫/2Ir"=M�::b��wy��GvgXFh*��s4̮����k3RCWi�oN�dl��{n���M�QС}�hڄ���#4Ҽ�Dv�t2wi:�{���(����><��<�u��=H�U�Qx�S�S����@��c϶Np.t���;��v 5�V+��Yr-�=�v�}nu���"�+�p�@۹\�ٰ�]nIK���f�e[Su@��c�����
+�"y�C3L\a�pe���.��淪0��;�c�mᾋ�N8���U�a� �k�;�O�Lw@�\j��1{���Q�4��(+g|�P�tjj˓Z��ȷ�.�X��]�y��#D5�V��b���7{�9kLX��
��W&��]�ե"s�(�K�7�٘=:;8��Ʊw �o���iλp�A�2;�l�4��:�`�ʛ��=�e�nDݓZ�Վ�h�T%Վ7��f�5�h�R��۾�ڤڳ�{zm��`p� 3[V).��\WY[�8�]��J<,�Me�ؕ��.ax�����n^Ч,cם��(GN�}����!I�#F����B27���Vs��={���Ģ�/6��Yf�&z�`�&(��.�ۧp��S��FGa�$�<�b�(s,��%���u��wAJ�Hk�[d���y����ti�yŔ,�vJ��7,�
7h�e��>�9�Gu�l�g� ������y45Y������q�m�{�+�cX�Ʊ��U��&BL,��((<���5^�w��K�4�a���a����R��هUf�f���D\�I�����o+x�
�ݥ�;��� �DܭtڮI���lf��yV(�M�/��qR���+�vIZ#��
vu�JBi36�lNH\y�N��mQ ��ρ\�>�E[�.0�6��	ɳh��qì�AI,����Lhg��6��B��7v��7�У��+@�n��Le�y<iXX.�q)̤�ak3$�r�K.��Ƕ�0�pճ	,�cV
���X�alP[�k���͎X��y��uZ⠇ﯡ�O%_](7�Le%��o�����T9������a$�{X8��*I��.�]fg�@�O+/PG��o�p�xŬt�-x#vn'6�\��Y'��U�o:;!!N�:S��'}S30ζ�I->�ʺ��U�^���D ���"f��n��#����3:I�oE���ə}3�tY�O"(|v��$�	"j���r�����)��&���=o9��@�/]�n�.�f��5qU�-Ǻ:A�9��gRˡ|	��J��-ď�-��z���� ��9���_�7�~C��|���
㝳	9;Κ�|�W2�f���,�z��tc����͎V��e����x�*8���<&��Ti�V��72��	'v��]�2q���Cj���ɔ�V{yu��;��X�y�wNQ���v�'��q��]�o�AD��zC����������U�fG�G���\�����G�n8�ٷ�4f'��Ccٓn3IZ5=��xA$��\��Nq�zZ�*�W��/pk*W	]g��wV�$��͹�r����3��&��u+~+8���Vu��g_��R���ZQI��G�t��k�L�ך�ʜ�WR��pֈ�GU�N�T�]Gbƒo��p�Y⾲�]�o:�tوV!��;T�W 8wy�J�#C�ެ�x��)Ѭ6�X�j�sO!�^Ế�̢�$���!�Y��P��t-��|q�b�&>��\�^:ճtyv{y��	�F�s�k&�n>}{2��.���h���\�*h;W+h$�n�O^vtJ�\��u�#]Gc��p�<��Y�W�m�V9�ݵ��+��캌Q"�"]�xJ�֜�N+��0�m`�vJw���z{p�E��ɰs���'y|�ZW�A*��_H	'C��3�U���ӑf�cqT�J(z��(��}�f�!Lu&^s�����ؔGsgu��yv��Y嚉�Q��czY�J.�gd�;�r�]C �7%�G�t�U�0�o���s���#eFe���p����v��+�6{�ԫ8���:历>���a���82��y�Q��3��[G4{���Z�o�e���6:�;�E^ �h�I���[��u��6����mtW���9�����}�E��B�A�w��S�rV:T�d�ƺ.�L�tyv�X�m�f�h�g6:*�]6Ɛ���ۨ����Y&�w�]��e,�k��l@����v[{ ,-����tQ��V�*<�M*���WEt�Yp_s���/R�XnMfHP�����TD�q��.��g��[�Pbd�*��D��Z1�q
r���uv��B��/Y���5�\��c^�^[�	�=��y���Kg�˓��]��\sd8�xJ`�ܱ�R���V�S<�k��o�'��&�s'�v�4��n��&�=�jIPe\3G_k-��#�M�S��5�2�1�ܒGN>�
+�D�/vG����1�Iu�)]䨥��e�u;o˝g:/\�b}Ww��X��ձ�2���)x�]�%�c�GrĘ�˗�� w7�^�E;Ʈ�ջ�˄NZ�����f�΁�"�Kw�d�톜��O{"�;ϜAQ}�w��z�g)���y��om�APȑ��2�Je.bL�	���N�ػ�n�`'�&�I���)>��/�Z�l�+�í"���gJ�ý�M�U�*�7����+E'��N�U7W>����s�Yl���YO.�[[Ͼ}�U讉]�n�U��o�����)E���7���vH�}�lM��y�xVs��L.odu�P��ؕp��vs:#���[%���PX5�汪�7�l�z��X��]�ʧ|�����8�U�Ba힧���>��+6M�f�M�I���풺�c�7�Amt2�v�����hgpr�]s8�CR�\fc+8�]w�3�7�v���*�:�Jq>�컦�	>�z�����	��)�K뵺�(�����>��%�I��b�29Y2�q;��l`AU��w�S��S�u]0��;81�v�Ћ�3-��P�$�[ s.�(�h�Utl��.�yON���k����uyt�Yν����b���7ݳ�Za�w]�'r�]F4rN���2���L��dpK_T}�:�Ρ��,���ݡ�<]g*Ǝ}���]|ЃZ�g�pيfv��6�י֝,�<�����K�Wr���g���Sn��l��ֶЎvQK��fsCb�1*�nfT)��pv�SQh��f
� �Ea-0�1���g��y�R�g��v +I�x�����&6�]�e.#�uiےB3U�͚��^��ʺ�e�x�DK�n�ǡ��KSM�eA��Z����k�7fS<!���j��D��>��h[�=ai�(�u��2�R���n:W���1��w��+jUˢ���3_/��;��a �&�]Q��N�B�Z
R}p�d�"�9W,��<%*b�ܲ�29�Gw=˺^e�n�l$�V�:�/(�z�#������vXy�x�}�2���q�wgdx�'U�8+��=�^6F훺!
yC� �y�^�!�[�Iށ�p��|�ϕ��7tm7�-c�,�脓��l����Z$�����5��X��W����F�4���R�r�`�E)�h�;5�����՗_\���9+<oA�4��d�֢ލ�༶d���I _R%"�c�ܦ�Ko4�a���%��;v�_IՐA��zJ��E&�`M�.�n��zִ�r��ڮ0|���]�W3
�R�ne������c�;D�]֤����)𘺙��mo-ݡ�do��ӔT�c��_r{�g[�w�gEE4s@���ꋊ���m�Б��c�ޯfίy���kD���� �͇�&��d�����O���l⛘<�^CaTx���ڮW={�7�������+��{�H_ey�R�iaR	����ܣ��ɩe�I��1A�\ƌ9�/z��ӱrum8�k�:3s1��uY�W�K��(�&���
뫾���b���P�E�e�(m�\�ʹpa9���:�{���M�80���<OL6+|��m��7��9�{K��y2+]\T�E�`��Sz�u�oYQ>��l��vu�؆��]�H:q�h;��mXj?1��4�r�z���KP�[�ĭ�w\�	���9��ɏ�.�N7�f>b��wWJ���9٠�|d�|�7�����G9�@o��K,4"B�t���*�St�����ԭ��^,�8��f��Su|@�v�ʷ+�R�(��@�]Έ䇲���U�]�'�eZ����~k|}��KKf������$��y[�r���)C�>#�w=f��ē�����Z��6aA����S�-M��.Q��ol`[��.��ͤVB��{)��]���m��)�W�s3�W�$��̗�X�H��7�������`�~�Ѥ��y��� �.�M2Hf���6�a��;
�WG���㭶g�7�i�wh�ފ���K�5����yP?L��+zn��S3���J����������u/�6'=vZT����u�w�vh
U3�bшd��J���vD�BM�v��Qާ�K�p;��m8|�8������L�$��&�\�u�^7W��f��oJ�3�Y��v�|jjx�d�(��d�gF��bp�5�oN�a�T���w �u�[u�_�9�\��VZ`4���j5v`�v�m�7:1{+�;�GsiV"�'{�y��rf�<��v'��C6������Y�` ��]�[���� ���P*�62oW1�´�ݔ��YzJW�֩w�b>�^
��dʲp�>ٹ�&�r	�	�oH��=v��Ӯ�GG3%�ڲ�=��-�U���1E�Z����u(i�4l��]�F��������廻p���P`˓%�ÝX�uM��Y��O�x)>B��t�U��\jB2�p�I�%!����dj�Q,R�23�]թ<e�JQ5�F����gY�ũ`L���P<���ʅ�H0��w9��e(��I��9�f(��3rh%c2��*�,(:gi������D�-X0���u����]Z&j�6���9e�R�ou�d�f�>G	�	�w�S��;uq�q���V@�����Ĺ��a�/=ϡ.�Zu��z����ێhxV:G�7��
���㆘�oMjP�c�IGɋ��&l��щu2X����g,�V�t��Z5c�B��"��m1{�RG��b�<ktk��ZF{���u	���j�����7`y�fۘgU[�;e�o�����sr�����T�ݛ�����0:�*�c;M*G;٬�^ý��C��Io/�%ϊ�
��p���*���ݙ�]2�4��b{!�w�G������:Z�Xφ�X�;	pE��D�>3j]վ]��G�n�d������fq�b��kjM��4��Y;������;>�eK=�#;ͦ��(v��n��.N�!�+U(����ڛ���Z�R{As;E�>ʘ�6��,��i�؅Y�A8�<GAr�ۼl��Yra�fv�8�t�yE��z;�Ln8p��Hk.M��<8݅W��[$��YZw9-���BM=۱�p�<�Q�q�qژ5v��م���R��V6�K.�&�'�v59�����,�/���L�j�m��t��Z81�W+��_�{����|~�&���)�qgI�Mɦ�Z/F�~d��9��qFﲻ���u�EC��6xd�͒gh��˥���@��zX+��/Ⱥ�7���\�R�*�ԥ�*��]3%�/G\Uv��J�xK]��|"F�|�r5�d����ͦJ�Z{Oe�`ݿE��$�����W�2����+tK��q���mT��u�D2���;
��\9u�EO����pׄW'���Z:�'�g�Lǋ���e��q���f�CN��T�N�XU-����2�qs�jp�?k��yֲ��E2K���P������j������fRMq�}Z̔R�}x�K��Z�i��^�e�K�rW�\�lOc�����tw��m�(M_P[��6�ٝ}�����,!J��z^jџ\Cp0s���PB;0�Eƍ)+�����4�u@���Ye-U��8թ�Qrm�xuIm01y$v��r�-r��d�r_��5��F��Y8�]����ǀ&K�m��{B�4ᭆ�2�\�1LC80r��]�MѼ���̠G]v��ܳ�5�cN6+h�J�3fX�pi4��v�_�S��m��L[l���(;d�d�#nͶ޸�^��DG�q�YKFG�Yr5+�3ď6�U�q�.y�̻R�x���2qΜ��&\����m���J��0������� �ڼ'jy�3����	ۙZ�wSz���b��;�`��;�zdr:'6W���N,[�.ս��Qw2`=�3x:QV�s�s��+Y�M#���ivNx2�����h֔�ͱj��w����R��SamMu�èugu�X"u}J��-����]G�X;' 4�:�k�\��:cF��Եh�.�v^j��_�u��[n������;:��Ƿy�D��f�uNc�o����f�����o�y�o���{�΢���-9}�����k��Vn�&��("�.�[>'؀m	��Ow�x��p�4ҕ%0c���JSi!n4= d$+;�C����'��!�t�s1\��X<I������8�{iu�GDLF�R(�B��+�w�j�˞rrB"�<�h2�����-�`� ��&�m��Sd���Jjp3��R�%�B��Z��BP>���>%PG$$�C��8�hi("�P�ה � �T�&��	�ˆy_}x�A���E�6�\@$ؑ�F(2X��.Bp�
���t-�����x�rf4O)�����@��l��"XA�����"�:�`��A�%T�4�K�{��=T4�*a.. E�m�����-��e�8�i��<'�'L(��6zh�)���d�(8\F;<V�vPf�-�`/=����XCKK� �ȫ1�mV�n�ؠd&�c�*��"!���4�(Kwt�j ��Ê$E2����`��N�LԲ��ڹ��P��L:%"B��0C	.�,9�j��
���*�Mʭ�X^j��CdE�  ��?�&���;��H��ܗ��I5�g`�-�#e��Cd	�P��,@ �GR���4��	��R0nP�'��,��q��<'�)L(��6Em�S7nm�M��E������8�V��	��P3	qq���N�]^P�C'!Q�������YYH�m�Z���D �!�cRA�V������.0^�Ɖ�5�iZ��mW!��*LA% �[}Y]U���A���&ď�#�iU�"�T�IxL�4�p��O�&K.��WK|J�#�I,ȉ��i2SA���V��L�X&�BS�&�%��	j��Ѳ"��c��4�c�Td�i�N:X�Z�����D+�/]C�(P4@��N6ˀ�R(��}@t�w
��xW[��a��A�E�U.>>Y-�.ae!!�Cwb����y7Mq��HTAq�E�쪦�(��+[�O&;g�0��J�%�!�%,�M&
E�|�/��pp*~������"�
s>~��K?�~ "�{��������A�\1��_��4��c*뛽Y��d8����B0oYݏ&T�ym�)2����6.�y�u�96Zɼ%:޹�o����7���ݹ�����M#�
�a&�U�{� U(^zBon�!�6r�*�X�]��s$�n���r�^]�8��l���[\9������Ҧ^�ݷU�sT��_�w���9�l*�kf�6��m%��u��a�w7�:�*>`>�ͽc4[$�ʷ�sJ���P��K}����գ�b�[�㷷:��2i��Y�<z�5�o�e��[d&��%ܤ�U���*��,��wD�TRV�T��n�5�䦤��dN�U�6sz�9���Q�������q�\�m� v�7t�u4�L���Ԏ�G7J;�ʆ�jb�f���B�ԁ��3e^-�#Yf	�խ�J�݌�Q˝��]J}�� �}��ƕ)1'ͧR��H�2��T��El+B�1t���0�k��Le*���g�8�u��=j�Q�Fd��Τ�Ia�qn����+qH�b=����w.n�\2�L�w[�~o(;~���q��u��]u��]u�\u�^:뮺��]g]u㮺��G㮺뮺뮎��OOON���]x뮺뮸뮽:뮺�㮺�ۮ��n�뮾:뮽:뮺뎎�뮺뮿]a�]u�]q�㮽�:뮺�뮺�뮺�뮿_��������~�뮸뮼u�]u�_��oooon�뮺�뮺��������r���-��6&�'-�u������/�0��V�]�ҙ��7���s����ޜ%�'sگ��'"�������D���%{z��)�h��Cz<,��*�ū�ُn�Q��X_>e��s]�O�"���1��G�&\u��;ڲ�N��baQ$�Q�ә���eV�Y�O��tZ6J6z(�r�B��;��]�Xq�=����^Bwfr*,Ie���Ңq��M��&����S�zT����8����vu�� ��K�
��EUݲ��m��L�ǘa��\��q��Ӝ�u�xU�Fm�U�U\T3�)S+8���4w���n�] ������)fƆ �m��X�C��֔�܅��������[���ü8�s�o��5��;J]��׾�q:�u�ux��4v���V$����eo]��ied~z��n��ު��8�|��(�F�;�b���T}EU�4�u���cbT]�֔C4n��w�tSr,\���W{ y��a퓏��Ǚ�s����u�!�ݷӠv�Z'+��P��H��P��7�=kY^����=���i4�{�-:��x
,�6�TfE�ܱ�u��o�����|q����^�u�]{u�]u��]u��]u�\u�]zu�]u�u׎�뮺��u�^����u�]~�κ뮺��]x뮺뮸뮽:뮺�:�N�뮺�뮺�뮼u�]u�_����뮺��Y�]u�]q�]zu׎��㮿_�o�����{~�뮾:뮽:뮺뎽��{{x뮺뮺�u׏ϝ�x+��Pݝ�����]�A��� y��խ��!4�7�h�7�ί/W QLY�z���(- 8��;����a#���[o�Ō@�HW#�	�ᩥa�@���z�iv����p�X�v����@�׏G�^�R{6GH�����K#�ǝZ��#�sF��ۑ�^��[0T��ݺ����Y�'c�dt�ZgJ�"��9��-��l�c�(�R��5����
�HO8D�m��UkUZ�Х����� �4QR���Ùڎvp��5_}W�^���#�e�)�y�Ӛ�Dp �Vm !�Hb!���������g8 ��, *�e�t��Sc�UHz����O� ��;�:M�a���`LvӲP��G��`�B�dF�b� c�V� a�V�y�U�a0�<�W��M)n�g�Q�gJzg�__J�G���ZVL&"��_����n�LW�ذ��17pd0	�̑Ԝ��]gّ��b�}*��(en*��k9��+$$6��M�R�������5xqv��Ybp��3F���Wv�W�{ٯy�Z8M&<�_V����D�[:>Q��-�u�����~�0S��k�1>��j��{a50�ԅ�L4����Ә�re���B��3&��4,';2����H�a�^��ʜNvt��j�z����U\�q2d1[��N�6Ϫ�N�y�qr�qr�͆M��\+F��[k }�Q��^<�T��b�c%��&v�ӷ�)k"ȅ<�u�Y���ǧ~��~���]u�]q�]zu�]u��]u׷]u�^�u�]|u�]zu�]u�u׎������뮺����]u�]u�]u�]u�]~�κ뮺��]x뮺뮸뮽:뮽:뮺뎡��뮺뮺:뮺뮿u㮺뮺������~�_��\u�ק]u�^�u�]|u�����u�]u�]u��;�Ͻ���κ�/J5�$��6p���w�O�B�r��q�E'�nhk7K��D���Z�L�.wZo�'�q��]�!z��-��E{x�8M��uO��V�#��b{L��SL�%�3L��q��Rs3q�w��4��ǲ1Pw�վڬw�A��R�V<o�n��y����S6� �_>q��z6͎qeh�benK̳��f��)� */�ɝ��.��;n�5�Ut
����k�@����G�/�ow���j�#W~�ŕ���<��a:�U.�e*֓�c2U��.A��w�4�<������ԼOqD����u0��݌�f]u��;�7��x7#��b�c7(tugZ���ȷ�3K�����q�x8�����a��k1�+	�x�=x�F�L�f��]��O�M
l�k[� 4Z�j �Z��m5���]��W�P̱��b! �P�v���y���{^Q�%���u)��N����iWR���owH���6tf�+��:���
���A.;�C\$���)X=lS�������ַ"�@�5����3�Ӱk�V
�N��h��'6��g�a<�`�YEZ�]�[�z�[z�ڶK��;�������뮿]g]u�]u�㮼u�]u�\u�^�u�]u�uק]u�]|u�]{u�]zzzx�뮺��]g]u�]u�룮�뮺뮺:뮺뮺룮�뮺���^:뮺�뮺�㣬뮺뮺�u�u�]u�]~�:뮺�����������u�㮼u�]u�\u�^�{����]u�]u�]tt�}g[�^o>NS�[۪��`If�Jk(���v�H
�����u�Z͹� ��F�W�������6T�άut����q��ʀ;�r��Yu�Y!Ԫ��{���"�Ϋ�}�����A�V���#6f����ʼ\ּ|+S1T�<����L)^���?�
#�M(��O��=jS��}�X[
!m���vu�u�p�,�e��{���qӈ�)��gt��h\�Ю��T�k.�U.��u��fN�#;�5�x���w/f�uM�F���%!��6�d�|�� V�*��N�;�a�C�{y: ��у6���=]H����X��h��w�n	PY,Z�W�]ѠCv��Powo�]�=/��l���%�S5Vw`�q��a\�,7n�*YmV��z�f.�����5i:%k/�a�W��N�� t)���f8�Z0����3=~w��#�AT�tK&̝*������qӻ}ʥr�"�drzw;��'X=�/\)����5W���+����^���c%^Th��$+x�&����X�P��מ�Eeլ[L��CY��"��[z;ek����]��$�N֘�<�,d�d������|g���������G]u�]u�_����뮺��Y�]u�]u��u�]u�uק]uק���^�u�]|u�]zu�]u�u׎�뮺���Y�]u�]u���뮾:뮺�u�u�]u�uקG]u��]u�\u�^:뮺��G]u�]u��~������~���Y�]u�]u�������뮼u�]u�_�}�tu����R�MZ%X�T&�A]�e�a*�E��ǟK�hQc)�y5J���vqɴX���/,�cM|nN���c�7{�vD����I2%m�[qma�vb��qs'�d:��̮onIa�\z��A����ȌI{�aa@���f�,����nҲ��h�m4EN��w�֢V`�zC]������X�J���F's(}��u���w\ˮÂus�O>�9:=d�^��v��[�� �k��am��ю)y�k����XqP�IK[��׼�K�k���k\E; l�W���R [���p<*�%�/"Ǔi
��E��g���:ޅ�={��M�Cj�.%W��
���t.����5����hƜ�Kov��rϵ��Q��:dج�6c/�������\����i�����ǅ.���wڷ���N��N��=���Yҋmu������_LU�wIx��f��z%Υ��%M����c��w��0���:��zg�7�o���7\e��6�N���e�٫Z���hu6wS��,�oMmss^.����}��Mb�e0v�S�|~/��﮺�u�u�]u�^�~�:�㮺뮺�뮺뮺뮎�뮺뮿]g]uק���]|u�]{u�]u��]u��]uק]u�]q�]u��]u�\u�^:뮺��G]u�^:��]x��u�]|u�]{u�]zu�]u�u׎�뮿\~�Y��~�_������]u�]u�]�����u�w�����{�ޞVn�b¹v�Ճu`�l�|�#��\�[��u�:z�H��uvV���>X�	K������H��ۮ��%�r��詵��V!�/*��DfHK����d��W{;�Z�rc����K����\"�乮�e�un����
��%�9Y!����D�=i3���k&�u.8�5��E��ɭ.J��u�n�u�Ś����s&@�#��r�CFaMc�����q�FiP��R��.��:�
�P��x��mq�=L����ʃ(n��%=�v�NG�Zf�۹+q;/"�ۢ��m��*�ڗ$'*l{Ű��ieim�|��;��tFԙ�xR��q"��`rX;��	J�f�.���D�Y3z�!N�}�o6$j���;J��Y��U:�ڛ��([����z�߃,�UUR�Er���=_�W}��Ƕ��vW���cл"{X��YeX��MY�F�T�<��J��5�Wn��؇b�e��7p�M����Eҵ�(c����I\���u.X���J}��\C^"h���}L����N�����u��Kdb�@�E1��N���t�/A�uv��#�gEZ;3��/z����I����V���q��\��v�<vN����usz�d�A�y������]�۽e�u���O�_8²t�H��5��m��j�`�{��G8�},�>�x���Ge+u)���^�V�*gu��x�0�ӬӼR>Z+���^��{��ָt�,'�+Dh��Z���C��$�?+���[�eA�og_@��q�Rnsl�fe�v�W���k2��1h·�L�x���(ӭpp�k"����ʲ���ѐp[!�����EҚ��»����ӝ��!��pf�5�B8�߯/��0[O5&&Җ��UkV��߁k���޾����j��0:[�%�λ,�IV�1��o3�m��B`9��q��g��nH��rJ(�&c;{w���Q�&�� "�UЅhz�2�s�xԳ9u!����V��C A�4D��nBI4��o;Q.^���G��t�>ٰ$I��
��6^�;�F^�X���|.Ϡ�v��y�i\�d�f&F�q�N�ƞF�t�x�CM���BOqU�8�{�n�Op�(�+�Kk"!�p��]W/�����T,���<���U�:�VN�Gi����Ӡ+��޶bZ�һp�*ސ��T���b�G��rںs+uh��*|qgk�6�3�]f��bȝڔ�[C��#�Ru��vT���tJ�C̣Q.�ŮU�E�ei���МŎ�(آ�q�Mt��Nmįc���^k�뽡���h�5[�.��ӓ�.�|����U���Mmǒ�t����ڧ�.�L��>9�h�7�o�����Tj�}�b ���������ݏ���rxA-�[��5�Z��-�<%��B��*`�-�S.�3�0���bC|�,��oL���������9i�g8��� ����㼳�^��]���\B�A3,ս3����.�`R֮�E��F��f]�����ڊI����!�L�b�%�5]�{�N�\��dտV�t5���U�M�u��-&v]#W2�3ݝF��8���u�K6λ�����_ �6+c�������{׻][�*{5W`�.35�<�:�lz�և#�)�0�����iLDm�`�x�-�K�8�����\j��諭��� �t�K�p�B�&*7ڮk�u׃��+)j� ���W&�
d�r��C~�8mq�����=wt�MW+q4Д�`5���tJ+�h�-��8u���n�Ϲfkr��3):�Ŵ~F�s��k�bs��:`l[�+Yu{�'(ٹ\���6j�AR���|���ϺTn��$0�ֻֽ�=j�t�1	|A�+��7:�#Ojt9�x�WI������H�n��>�r��
�ݭ��]e'ټ��n(���1Dme>Q�XZ��8�����c���]�֩+��b�;T�ŭ�����N�Hn��8nZz��pAQ�X��c�m,x{��cp̽O�$���wm$f$ņS�|���cw��B�e�ɱ�a��]`�[fi]�PY�����(i�p���:��0A|y'�3 ��/����xwk��siXɬ�f+*
�r<;�ȧ8MK9;�J�
i�+��m_Q��nRdu�hT�
shO>{�������uݡݗGsn��G9Bs�w_7y�{�7��?��H� �����?��/��/�o������@?����@�(�F"�h��RB��� ��i��aB��+v�#B$�A��PAV;4@J�*��(�|R���H�TJ���;�FIi� h����L,������
P�(v���o���j�ZX���k��kjv�����NB���c���!�R��iˠ�B���J5�Z��RGre��݉�����)��Y�	J�/.��[�A�PRY�r�q.��\�,���f�^�¯0[@D)�X�w`���a5�(`�gh�;�B/td�@��s("�oXX" [Jߊ����+��IXf5�wRΥjДRR���X�]%��W�sSXdZ��t�.9��M!��U˷����X�e�(
�w�p<G�7�Y�] �f,��+<�F0Ef��Atd�C/Bvr-���Zԇj6�X��]e�m�9��L��9d��r�s��;�\]YSi�<�T{�H�ܮ43�^o]j*.�X�[�uu�fM]|pvmӒ�>T�B�J�ɘs�����:z�$�f�3�R��-��[�%�K�n�Q[ly]�&'�_6��Φ�բ�i-u�(k�N��t�B�9��0nC�d�__Z&n�V*I��jKV�i�*�9MM�=\)�R+1Ҿڌ͢�7���cl�]܊M��Xt��4��q�t�hQEG�[F��
-q%I��cK&��e&bD@8�"]0�-�R&�)��0�T͖£e�d:�d���L#-��!\Q0OO��"���Xj	l�
 �e��rNH�\ ��-��\B4��	���CA�w\%�"q@�A�P!(�b7i�!��4d�DQq�RN���A#�I>!�ݷۮ9r$Ԗ}��w�9�9��t�OOO�>>>=����_s7[����V�n�ڄ\�-��]�ί&��Ԣ�����/�W�瑻�]�wl�*�^^m3jU P@1%�=��>8������?__Y��Ej�c�#�	E 4�rT:�^H P�HQ���<U˕���b5QE��Z��Z.sO^y��DE�幮V܌�d������.�kgu�*�J�70kwr�Cs��d��[�*��n͎��bA�9S��}|||{{~������>}�\��LX�w];�e��<�d����۵���淦�]p�;�R�-����돏��oo�믯���og����!�M�B��],������N@E�޳��������ۏ�������:�T�}�z��k�#D��F��[���������������u��<{`�e���
���l�܅5�nlm$o�\ץ��RREc�.���s����\�{]+��h(�1��p���*���Gh������4�����T�#@��H�>��e�s��8Ñ�ؗ4+3�Ln
��ʟ'��_},u�e�p�B�gPPt @%RF�H�PFD�����T�`��W8)Ҷ�c��˵I���<����y�i$�p5[�\�.���M�㱟g��0����RW��ɖm}羟x��Z��K�
���C��`T���V�%����7���W���*hW�};v�z����}��߷��q�؟:��}�{5B�I�Q�|]���(�}��o�x�B-~:,�����2�-��������Ό}V'�?v���S����{�E>c��W�y@����o8n�4!��j�f�56�;'O��BIn�����W�̝K5��,�!ڬ`�״��iR��(f��!j"���oN-^}k���RʀI�P����1�psMɼfmTh�Q���t2�CJA�3��j02��%eܥ�v�gW���n���m0��Z��;گ;��f��T�nM�5�'r���cy�N�7'�Ỽ,U�-^�M7�І�;{�U�̱����@�o�dɵ��`�y�ջ9b�g��m�<�z��\��1P]�m�ɺ!��+,�S�*�7/P����C[� �2�@�=�y�`�^n�fJľ{Z��3$��E�=ae�}�1v���iv���V�
�f\�h-����i8D�`�ߍAPh��
��4�;�����ujk7@��X����wR���Ti
H+�)u�;��7����%M��||�;�:�c�{���{3yȞ/>%����������5W�����N_J <u�֗P���`�O��U��},��|iw�mD<��)7�]v��k��7�AҔ��d*c{�7-�i�6l+����e�(N��	�t7���}���j�f��1�lܼR���Y���)\�e^bs�|�#�
���!i�Κ;�!�w��*8�ګb��^���𽋀�T����K�_V�۽�4^)�[G! �����I�l�Ǯ���W�;�"��,�1�����˞Зz���yx�8� �;�
��"�ey򃎱o��-���WA��'k�W3����[g��h�*���y�c5��$�uG�J���w��/+�vugn��fI#��ރ�{�lnImE��vvh��v�ɰ8W[��4� ����訌Q������|s��=�BY ;˥��r��v��e)��ʓZ�3�Ǡ>
<}�=3��8�E�#1j�|�yX�S���بk���t��@t�Bc׽�m��rw�^]ٗ��*}&n/s����M����>�PNuQ�Qlbƅ����}�zvJ:� �߹�6����`���zx꣙y�'�>���Wc0u�?�w���=�e&�H�-�����GTo��	���uT5�?��?\���/;���M
\�P����5HR�Z��M�?Wd��M���V����쑖͏�@�@�^b�,lpr�,�x��>:���X�{��=X�8�y�5�B�/7����� ��n�j�z+�k�@�|��M���B����hx�e�H�$�ޫ�f�[-���V���~qh����-ȽM,Uu��@��L˪>�kp�U�9�!�ab�9��u8����8��,r-o2�;�=�q��1g�<��h�a��������gt�f(������|�7>P�{��A��6�M���	��zJ�7Wh����7���Q>�TI���:>�����+5_�����RuEy�&��	����%�e_)nўj����m����7��3��8�� �9��s�6�
�=,i
����U�s��(GA}ܪn�ѭ�*Ja�UO��ڜ�
E[�xO�S��a/{e�N��ش����H�������y��[�G�=�ΤNs�v��FV�px>bʦ��n}�x%��R�Uu���.�Op{O77^�Z���Ƕ��(�[�BՄ$c���������}q��I��!�U�� ����:��L*�Ig����ݿ>���F綋wU�^��%Q�+��w�Nv�<�]y��Ƴ��5U�m	 V��W��q�ٛ��2Ö�k�p�[*;IP��}���v�U]����^�k�t }{:l�������Q����c�RQ7�b�r��Ĩ@�3gfW��<]������;��>
�tae[ T��� �*!U��AV�Eлz�r��<s��)&�X�ӳ�{0��E���9��	�(]s��Z=3z]a(2�8V�6j�"�j��dƋ xZN2A%:��@QV�M ��L���8H����!��N�q���0��Sa�XE>*���u��~�4�	�vT���z�9��e�+;#HEV�g��ay`��ӭu�x��sY��%�5��+7a���e:�ֈoIK�ݥZ���e]v����V�Wle�&".K�,#�7�����x渼�!��$;���6�aZ���,�؆� �n8�_�����u>��ݲ�X�@�[�ZQG���o��}�w�N ҿ���,��N���4��og<��J�;f�R|��5ݝ�&Ѽs�%�C��Tbm�G�����]˪��u�y��J�;�O��sF�k��/����{:������������®�>��?M�B�0܆2F;]��L���;��]�;��P =o��J|�[0nq�W�r_�[.q������r�W����-��,
�	X�P��0Ws���ce,����`MoH7E˴��3lE�MgU�hi�|iĩS����;YqW�ޙ]^��À�/Z>��-l�v����ƹ��k&��ُ�+K�G7M,����}9�XS�N
x{=�w[�ZA��P������^K��[ob��b��V�Y�"|�S{&onEtۺ�w�Ms��Vl����о��t�o>_]:���ϼ9���N����Ĳ�\T�l躛ĵ��9���<nl��^nnv
����s5�Zt���O-��;>��ewo��?}�D�ZW����ILN&�xLZw�u�z�6Q ��N���A���������j�K=tZ�:&��l�5�s���s}�?^�K_I�rWʐ�{��2�˘+������s�/�� �g�|�s֩C��CUZ��Z<�u�S�p���-�O��YX��!Kճb��m�ٸ9�w�>��L���Lv��P���'���s���;<��W�"�y���A��Q��Fƾ鄂4e$���MA ��	k��}��v�@��|�����lr91�j������3�7����)d�5�{�9�x؃8�ۆ�c75Z<;����iɜ�\��I*�rc9�ʝv(P��9-���-A�Ӹ���^�`�F�w�B��cr�%y�d<횽.>�Aw8M�p�U󪝝z�N�}�B����ɡpGག9���p����W�=�n�x����k�z����،ƍ���� y\�����߀ݡ/=��k[��Vj�<�#�5���!
J�'�'[�`j���y,3�y����3%�r��p�:$��4�{��]b?/<�xU��*��a?��{[2շ)�+*�jZE�:��=���i�RL�Z*��+�W>:.�|�j�����¯Y�j��o�-`��{�1;�&��L��5�T���VpW�'����֯ӘG�Oe������5��g}�^写�-��vu�x�%����f.���!( I�JR������j2�Y*�S���k���_� $�W>����}��N}���+�W`����{r�]@��/����}��t��I�	Bv���2��"�u���h��>�r��D8T䈿�X�9�(��Ũ��� K�7�B;u�J�q]f�~8,���.M����Õ+\G��)p�(�#�^^M��u+�չ������՜|020�k_,7�fu%֛���yO�u�QE*Z��p+7o+wI�242�
ޱ�E�2K+��]!�_��샒"b��H$>���hKE��ƉR�7�XO�2��J��@k��l'Y�K$�5�aE��N�%��a�!���]��d�"I� |��L�����7�3�U�K`���싡�CC��yH[G`
��rH��ZY鉩��Uz���6#f-��l ��(,��{����Y�Ŝ���Wko����e^�|�:(�,h�&L [0��Ɯ�Z�,�4��n}��z�$��a&���\�f���94W��s~��W���=:���7s���]�{�I+�J�^}��(�3g�^ ���QܚX��y��?fԹ)���]�y�u�^| �߄vWދ~_J�}���m��E�2el��2$Ӯ�=���gj��o���_��t���^��uw�)+6Dǲ�++)e>��F����8�sa�R<�j�*^�y��vGָZ�6V�\����X���]r:KDL h��DȘtZQ�D(� ��Y�p��4�  �T��]�a�-�a� s����4��0��[����
`�+���V*��8�oLG��/�
�У���JO��� ���c�SQ��1A�."
��!So�j��S`�[D����t� ���8G|�@+����v�۝]&��� 
�8f0L����I]mLm�K{%mk�����������V�����H�7�:?{~��4@�8��O��r������S�V��УQ�ݘ�[��Ŭ���xR��s�s�N�����}��������m]�eڟW��|��5���e�n�̖�Q�a��C^]����܂�s�^������pʞ�/vFLJ��R�ӕ�i\�3�
������5�*��|�5xH��@���h�挰�E�xUa�c��� �=뫭��p��z`3�lm�r��n�Z�;�yR�)�����;-���V6'Yշ��%D��U�`&�]�iQK0���Ŝ�_�m��P�OTW���7�G���6M�1�+���z��+S�r1�i[��N��si����;�TF�O+|��l��P����$zɾ|K�ǹt�X��ά�q�77-;��:�e^��m|�{\z�/�N�)���	� �=g��3Q�D�6+�(_Qd��i_to���ʽ���b�j�����@�qF ��m�wX��c�Ly,��os"M��|����\����\�P�h�|,�^X̽�ɧ%WZ�`B�^L̠)�x���Ϣ�ژ	7�k�Sȋ�2���u�b�i+�SU�Z�o����װ��{9��m�ǒ3������u=�]k��9�Ky�>w!l�
�}���/J�s���+
'\e� i���U��A0��wjR�!���2�ř	-{fk�H��0���L+w�Q�M[�4�(0� �?����ŭ�+ݬV�w	Ea�t�*��� 9�3�x;�7����Y&�)�YH2�#��-�F�!��2e��S�W��ڒ#
�ݣ�en�vqz?J������U:��[�Tyӗ�4���>����lR���l�I>]�C���C3X���І"gһ�<�}�뽾�r�c6#�:����ʽmfk�YI<��d��C�=�u�r����~�f�w�����S�>oztf�خ�$�t��+��>��^����uP��ߐg��m��)ԙ繯6yJ�T
�6�):x^ev���w��
�2�Y�R��u�5����IP���ݲ�,-�FY�:+i2f���Z�u ��b���Θ�n+���2'e|h9Y�n��m��r2�W@8A1�n��;�-��8�Fa�e�P�,�ǲ��ٳ��yk��M�e\W]w�ZVڙ�A�ُOY���)J��paν��HK	HU�	M�v�c�ٟJn��@WN�k:Z�6n���]�W�et��4�n������))e��lL;�oʦ#�����.�]Yre�T����!k+1m�ܖ������o8�v^.k#9�v{z��T��\����oQ�"Õ�������jn��"�q"��5ٕok�T��Ŧ)���0"JʘJ�e%��S��
l��|8��=�O1Ps\.1<ή��h]�ޙ�p�������rK��}��Pz�ѝe��v�����NF�5���"1k��wh.nt�q�]�2��]�u�F$���V	h�kw9��aN^k�:���7��h�V�8�黰�Ӂ��%��>:�1�
��M]#@���\�:�E��ZtbW(8�|M���R��ͣ��2� ������?.X��_����alT�LZ�-Hvk��텻#�l7ó�ooD���P�-�L�]��ƑU�p�n�R�}�s�]S\j������fv4�f;�x�V�ۭ��G���)��	|p��=��㷻�,8��.^.c(Y}�����1�6��U��S;J�f����Kp�0�`f$�"�[l�W�4h�*^$�ubo.]K�H����}�m��ph�N;�$��͡Iv���V�1��.A���>xQ�+�ڕ �#t�bM]���� L�j�[��ݐ�DP݆�n����M�.7Ӌ�I��Ӄ�y�qp���uۂ��-���Vt���v�tԩ�V��ˉ�KKB˼��%JS8�M�e�&tH�}����4�j��;fH��۾�ZJ�1RF�+��B��lbkV3�<��_ ��d�ف�SmT(��ő�r��v�`Ҏ���+�k�.�̾�0�0	*�k(6�+6<ǚ)�5>���S����zwz���B��ғC�"�7�Zѳ8X��d��� ��ޜX37^�V�h�B�� ۣH,y�T;���$ $l󋫛�x�R+|m�������׷����Ƿ�����<zgO/��?{��k_�������G$(��=������������ק�OL�;1.��V�H��i)�(�
z�Oo�o�����n��׌����ü�PU/"���Q����X�Pj��=>���>>>=����׌��gN��}m���TFţ���yu߾yxѨ�"�� ���ǧ�׷����Ƿ��u��Ǐ���Q}n.�_}^'���o�,E�H��b�)ݢ�7���o��z���������ǏY�o������׍;�>y��^�/�R��^��sh�n�ux�W�滺��W��5�ۦ�gty���b��@�1�O7+r�o;����u�^9x������b�;�cp�$צ��&��Tj�y�R�pW 2�6ܪ���^y�i����a�f��k�����{-�V�+rF	��c|u��;�����U7�0�3�s��z�����q�k��>�|�ל aF�H�q�q�z�3�k�x�* �B�y���e�m�wC��x1�0|&�.|'�5z.��7��Z<@F �����ib mc�R�U��8�{�G�{/U���<�>c��`'ӾsX�<���9��	�Yߗ0�o<��]���kxq�F�D���r`���k�ټO�pW~�w�d I �W:9l
��,���?|��[�O'�E��z�θu���>��昈36�{��{����Ba�a���Zh� D��Z����9d7�hyZ@_�����N����|���p�;.�|�ٗ����/���p���@F���Dv�� ��TxE�ȶ`�Q�	�p}��@B[�i>t�6�{�&�l��<{�_��g�
m:��}`z�	 )�s�{f e]�C���3Sq���+�o��2��e�x�����pJ��2Ut,b�qpE���{���@F1��Ǻko��j��L��q�!��sY�Ą��e^b��V��w�a�qܠz9 \z_���0wF,�>��h^�`��C�q̵�����6�#B?�=�ܑٻÇ����<#�C�7��j>���~@i�x��.i �,�������p*��JL�=� ۯ��Y.\�73�V���DF��n-˒�������N�)���L�*�f���G9^lr��×n��&��f\r[y��N3�g@h�
ųu�4�Jܤ�.�N�z�W]ut\��|�0�3�O�9��f��t�� ���h����T#y,�i��G�~+O9|jrs��s� �LW?��6{��%��g�VWp�rX)C�V�@�L�ʹ^�$��A �>7\0�z�#o��cX�����v{VC; ��<E$��tǄ�[�� <�^1ʛ��7�9a�9>o�H�	�@ǩʕϵP3�+�c"8x:�D#O����|O��5�[��ۑ�D	��Ԧ,���d|�����Goj��sxx ��`����D�m7x���H�(��^��ka�x�U�H�X:�ỳG7�'��;����ǃ�/�-�+V��O2�<ӅAN��|�|[�S o;�32tv�^U��O���dmx8@�if�@g^ i�ؠ ����v@�R)02=�m�4oC���c����;\�� =2&�c�@J ���H���@u�p5�#�-߿�è�Cw@K��4j��S�R�^���a��#�V^^�/If�(�<�k�l�����>�-��(�#�&�gF�f�d%�O࡮X�z>'��H~�.)Π4�۠m����Q���Xy�M%�>x>�O�M�<�r���A���粡����F=�x�2���w.��Բ�];y�k�x`���C_ �"b�������� �v�aDH�����e�q�>�����6���Y[{*+y}��q��8|��Wr%��s��󇡧�8<a=�νh]e��,2DR$�B�eFSe�2�R �
)��=��<#��p�����u.�H�=���w��v����
��L1�y���=�ce�I����^�O�R=[s�E�xQ��pu��;bo-ۯ�ߘ�ޢǵ�!+#��d��� W�_n6�G��;}��_|sP��|�������q�de�!'��s��1�����R�pxsg/�p{�8�{-�h4x;|@P�u��q��bj#cb��s����q�E�%���E#�4�V�*b����U�%#!��ᔾ tƀ�zg����w|�]wY��� �U #> d0s[n���ǫz Eo?S�;�is�T�����=�'��xq� ?P�ޝ�g �ozZ��SW���E��~�[P�{���U�� ���]TӋ�<*e��3���gs���n�Ը�e���m@�H�����&-�O�}>��a �k�~MQ@�[Uu-�QĀ��q��h�<ǁ�`�0 �C�i����W���`#ĩn}xO:
	��<���]r+7�Ah-q$�%�4>���9��������!Ő3�A�z�C�����0Ϛ�9��>�,�Ch՜�� ��a���kN��;��'�W?�<X�8���� �u���ȉ����"�+�a��7�߂N.@QI�ӦO�|�c���u�.*x��ƶ��eҖv/S����ն(L��Y��'�Wt݊>ۂ]�0�g�Q����E+iYF��2�u���w;���
����mVw)ن�]�yvveA���;GN]�CH���:�#���<�?Q�0�3�f��1�V��=�aD	�c8��#�]��4�]�� �
�i��g�	���0�����{gN�]�/̉>DvD�L��D
>��R��:'~c�����k���`<�md����{\���'y����ký^����m *w�,�7XC�����,X\��pO4x@i�,|;�|�w"9�ڥ5.�ջ��w���̠	<$��&0�kSOD
\�փ�u��� jm�#�O)�*�wh�C���]�3F���F'���QH#Ͻ}�ظ(��}a@�ϋ�p �b@f�MJr���[[ӄsު�`��0���ƏO>4�ځ*\\����$�#�Yz���˅å���w���T��d��;ʛ_\A��I��uo���>d8�Y��f�D��8٬�����Q�S��:��
\��۬iƄȉ�bQ C��� G��N3Q�s
1-FI�:)=tE^Ouc���#���b�a�a�����#S�`% �͐�J�h{��_W��W���U���mb[4b�Y�Z�7���fQ`b�a�a͇�z ��z+yM���dp��P3+`��E�GsEǍ8��!n֚{��	��W0�Đ�����X�x�K���ڭQ�}�J�K��4�>Y�+���awU��l��$��c��RG���{,�X��:��=к�(x��V�?�f�a�믜�����k�=���}��X�°����|��{ l�|�>�FIy�ݙ���a+�8�z�4>\���(�|�~a�L&��	�c��'|�|��^���y��6Vk��0��:H�׷3�Ѽ��7��~+i�a�[��7�����b���!8�K��n�s��m3�eZyn��3VǺ��y�����ؼ�����>�ckd�ڄ��A=W�@89���"�_Ga�,��z��i���BL��$���1����u���\�(�?b���=]����BkH>��b�Ѵ�6��k���{�W[Tqs"/b��R��:�c��7s�O���s��C�������۹m]��s������I��g�������A�/SP�S��	R�3S����7�BZI{88��=t�t��b��Ѳ)�8��H+�	�~N.H����	���O�>�x̨�;�w��\Kca�!�sǡ��{y1�C�
K1Pj�^�Q5v{i;1b(Yz�SO�Z8[�c�WOc���b�����	J�
]p!_E�9��\�}�++�{�ߑ�σ�M���K6�`���V"l���@�΋���M���<�V��rz��e�߇)���j~�*���|������e�7[I�7s�ח¶��i�t̓=C��{ƺvԎh%6%^�`�G]d�o'χ�.!� \C�4��j�h=CL��7p,`�����]7O8��E�UwE�1�ln�j�)�+��w�ji���y6�ikG�CQ�Df��^{���H��W���7�Hnqy���@cq�_�[�bX�L����ޣ�'ژD���''�9kI�t�ݜ��Cl��a��s%��[>�x
����!mÏ�S*��zK��I� �C�ab�&��'u�9a[��K�cv?M���:�n��ڞ=��cU��k���*}!ż�
�HӜ:v��	�G@����T��?;Oo��}M"0[0$ҷ���g�ql����:� ��ZW~�(�:y9�ڗ�8$T�Κ:�1f˭n����dgF���Y��<hÍ�%?�̅n��㵃Z	��K嶅+���ݺTع��Ųۋ����q���!��0��g�*�j�3�'�>M����/W�V����p��2�2ݰ�0d�-
j�ܯ�f6=(��Z�Ǜ|rWh�N6<V#�؃�,�W�z2�RI=�S���I㾦s��M�������8�Ğ��5'�/uN&"�5��yi��Z������3=x��Q���ڔُd��G!���������۠n�j����&��zcZ-	�:�kJo�^e�!L��(��㣔��z)W:��-�&��7JJ�H1J	!,A肜va&K4P1�*�Z�e�a�Q`�ƹ[�{��A��E�Yb䖟M�?s�q����
ꤳԘ�k6>9=0�Vw�ņ�r`IV�1��8�'3_��,(�%���G���	
Ȗe1�G�˴cCZ����5���@�g)��$OC��é�Ed1{dt��� ﱄ�'�	��(�ab�l�;�*�5:��$�S���}U�#���ƈKl����#˞�L� X��+T��g<_tB�"Ne;��h���w,�/"Ѹ��[�%�A��y��3�g�w����s�F�Cje;i�Pg��缎q���Wm�Ҁ��a��Y$Wޙ����X��l^��(;���!�|�K���+y��u��b�갼���?GI��ڑ8ӕP7i�ۮ�ry�o �D{D�8r�8�^Xi;B�sGd&����}�Y�����ce%�;�L��9�t5TC��,R��5�p��u�|�P�l_1ٵ��v�{�a)$P4�[A�{�}U�
��?t�VҖi�YsXίF�6�Gc�mam�6��5dN�N�3R�{��hv0�㎜+YÂ	ܥx�ͱ��O<�oG)����{�S��2^��~M������TaPO�~�?I�Jb7a����m��Z'S'��˿e	v�?Fϲ��˺a���io���P�(����l���r�>��X�y�d���6���y�֊S%��P+\�J�P��%nN�\�u]��F�JkU}�,���#�8B}�~�Չy���3ٴ�>b�b�q����k��O6���m��v�{�i�YI'�Q-���)
�=G�����g�$����|+�\7=[ �ۍp�z&.t�{<�E��F�9�J��Ww6D$gVB$�4�n��/ïx@Y��E���}�|��g�a�Em몌��f\����S�uk9�i�|2}�T�q�D��x�����>3��>�<�Df�U�7E��M*�
�_���@�P��r���!$y�_\�43!2�ւHN)X��C��V]�l���(n�[C�l�ߕ�F��@#B�~XI�t0�����E�Nö1��;�ذ�p(��y�ֆ�b	w~�E�������5�|�WڮL�l�"�8}�L�2A�c��UL��8moZ�[�y��2|��@����̐(�^��3����〃�DW��y�8�Yd����8�:��
��.����U�1КY��%k�b��2������;�24�Cy���%/>18��oI�a�P鼱v>�i4�O�n�v�6���� �p���>�����.wRm�҈�Ln3VY���R��$[g�l��\�m��r��b�[(���7{� �9dV��-\��]+U���]����[� ��+���L�
Y���QN�ե��qӜ�VeܳL��lG�a y��h٥�+�2��¼zӁǲ� ���e�DQ�+�q�O|�c<5y�#V��&����6���.kV��9cl�2y/9���rn�lf���ә� ���n�(�nk�A3���2ٸ�U	�����uG#ê���r�A��+�#+z;�j���#l�m<w ��Э���})�TB~콵1�ǝ���pa�vcy���%���j}E�����FsH��n��R�����
�#�2�?y�����φ���X�Vr��b'ë�{=��0Odi�rvf篺�7���9�y����p��7P�(�P�63���Kl\=T���4kqB����ڮ�*�.͞�����_�2����F�(�@�kF>8��6�Q��Sf�_a�)$�����*<��}��>��o�$~�d���OUoN�<)�w[l� 3�A:�o��w������C���+��G����bX���A�zŜ$�p>���7�ƽw����!����g��:�6o	�h��rl��,��y��|��16]ϮS����ާB�;a�s��y��y��tUz��e�����N�q���]�Nv��z���N��S�Y��&o�c�����ύ�F�g=w��)IfZ�p�����]��++�n���"�>[�I}��g2�=
צ��=��<�[�T!2��m�j`4�5�	&���|��4U�O�Jx}����b����=>>2�y�؎�~nI���:s�v�yV�{⃜�Jأ v���(3v��*��wq���W	��{I�Ip�I6X�X<=�nK8��K�Yg��y�ˑ�����k���!��>���jqv��ӗ�V�+m��=�do7�rEcɣ��(��(%s%Up��^4�XF9����Q,���_(��7���v���n�:���H-%��W��iܯ:Ɲd��A��ZƬß���Q��б�^�gb�����������n[[�:W�c��W
������Z�ŗ���R�]�-M|��w�n��g#J�zv�,q~4�7.���t�<�L��j�4�_�y�b�@#��w���1,'�5��g�I��}�B2���%e2<kߋܽ��?���.��<hN�1�w*��Xk����ܛc��w9���<2�͝�R1�c6z ��,�kqQ��ab�kۨ���x�x�}ۻv����_y��|���T27�6�X�uόw���/��|b �+ ��9�ʯW�M���ϣ�1K� �]�,��ĲE�^h���3�Q�z���6�#��C���1 ����@�w\.���j�;<5��aR�9[f��׆�=�Wès��:��yv����8d)w'�}ͫ(�SU͍VJ'�\�Xv��3����ۅk$'��۳�;݈��(�S�	�cD2t�}	���6����vf{��i`�0Խ��;N��-�AzL��ʵ_�yC�o����&A����#w)���"k]�r&�̰��{�
��ye�e��tC]gKn49��p�l��c�g-]�fe���҄I����Λ���n˵,��ݏ4gS2��yt���J�n�m���ww�F���X���y8������OT}!g�>��PH5j�wU ^�2M��t�i${&�]f���
ƍ6wZ�,u+�򱱎>��]�a�y&'�:�j�V���t�U���L��U�5�����cScN��9�pl�i�´��D��v���ul�02��&��^�O�)�α��)�W,^�m�^�玱A���u»Y[Ԧ�cɅ���Պ��[gr��nWP�������VC�ɯ���j����K�� �˙�$h����m�%;1Ra+=}g.@��D�ʐM�M�JBcQ�
wF7J�5��k*--�B�kϥb�,��M����0�{�Oq�
w���樊$+�
�Mɸfjc�*��bRGr�Ú�dV�ӵ:�B�tY*�!Эb�ۘ&3S�`=Onn��3r+�dx�l)-@ꢫl�D%J,R��g1��Y[�����_R潾leB¡�H�����議��on�t�+�6�
�k�A�a�V���q^�wF�q�%o$vж��"!(ƄRp5	c���"�i
&�)��5W�D����1����Xb�v�»�s���+c���VX:ʄܬ�Wưo4�4�(l���]��v.��5�%+4Ю�Y��<*��󒇲��ֻ�J�je@��"��ǵ4�r}}W�Q��K,Vs����t�s�0b}�:�E�:t1��
�c����J��gAϖT��{Q�5Qb�������H'�bƈ�l��/���.���.���3��]/�%ڮ�O��}hY�0���*��<���i�G����u����V�b[�;�'{yY�Sǃ�Ͳ�H�����%�z�O�N�^守yg���(�*m'�e������H����*z�0��r�]�J�YH��s�n.kVa�ܺQ�M�v�f��z�ü�8o��)�쓪�r;�ic47��s��B3�oC�%�&���3R��ez�sT�ս�[YK��Fh������N�y����*�BS`���7ݰ����u���y]ni�t���XiNCyQ�LXj&;X��q��y19�h�>���}��Нk3���Y��VsP�S�y���Y#��T�C�6�6�pzFQz�ʦ֔��B8�p5�%ѥI/4@j�JQ
�,��M��.Mȋk��*71'"����r&+p�m3�b��gd��eģ���� ��BJ��'�d@B,�Ԅ�QFa02�HQ��ENH�d��1'"�B`�J)#Q�.�b��m1\)Ԃ��WD�!0!,��H�ÍNB_���g�}q(��k�+��ܭ�׃����ы���==>:��8���?__^<x�΁�����J���-ʹ���wι�,UȒ�Gf��x�q�q�������Ǐ��}�9ǈ./!�C P<���|���{���s�BD�<�g�N8��q�q�>���x��w�l�4��s�7.Rvr����h-�_gӮ���������q��������Y���tp=�g��(�(=���E<�.o��y�3ǧ���\q�~��׏:�h����Q�I��_Ux2���x�h�<{|||~8�8�>����u���O����\ܶw]�}W�)|�~xj#��lT���Twr;�5wt9�]��>�lW��}k���ƍwtN���y�kŹ%�.�67K	�w��_W�;Isr�+��v����q.p8(u3o���UJ6[*I�K`B�J\�.��كV�WqS�WC����H�N:zB�2�	� �ھ�ċǺH�!��ZD�VT)��d�I��d�"$cM�)�"4�T��+�p���T8����X���mvx������j�y�s��~�J�.^�#�������}��[>�	9�S��1
p(�Ֆ�zJ�`�[�s�g�R�{�[6'�����|�E�-�#T��:�.'�����;[I^���! s[���|k�m �A_@�o�s\[�l�����u�3c���fq���4YW��u��\iT:ΐ�ޏx 	P�H��Ig�cx���]Y����<j	aM�������ω���,+���q���MxC׵���/��ȶ4�y�L>R�c;ZI>@�%�	��Af�+͋��֫�>��b���8�&�i3��{�ʶ�z�V�0�ռ� <�fL*Л�J�B�,j�^x�z�f��~�h�3���>Ҫ�k3ZQL�lki	�k'����h���;��e��_̘0������B�^�NY�T�;��a��"%�lY�̀G)���Q�c�� �<e�^Z����
4SM}�$tiL�WjR�m4np�6��,���t>y���Z@�b)x٘ښ �
EfO��a�(�JД���>��v�s%��dG�`���,�YM{P�|�K�Ӌx�Cx_���.ye�?v�c6k��p2S�W�:�R6��|�d렋]r�u�:ǨF�.����UD9��d�.�[�A��r�3,ls	�W9�'�"/����O�	��-]xytŠh��*es�:'�����#��y�����뻛����k��ͽ�J�+�Es\��r���Sc0��F�����ǳq@�����υ��ܭ��<p��y��#�1���L������u6qKջ��cR��j. ���>��z�s{{�J�Q(�U�X(Ǔp�����/!�=ͯ�����������g�O3�$�ϝ�w��?Cc�T�v����g� ��iFF����`����c��7'ͼu�梵�@��Q�j���ݙ�c`��t�&	b�@��u�}�|:e�ԗ�5r�9·�o��=�7��K��j5����4�4*��l�Hpݫ\v�a�>LN8N0Yoi+|�6A�~Z�&�Fdy�,��P�muo6����g/��z;��Rh��.x��㖂�����OC*c��|[|��4�Z�L��D%��Ϫ ������wcʣ�s3����>���3�c	���j�|5�!K���5�	,#c�*�'�i}\��k7'G#u�*f�(��q8K�3"/!�$(�NR�j�P�	^�N�B`G�s#�De�wl���V3�/{q�����պI��'���ѵ�6��Y�\�rߋy�hq�Q�(�`�� ��5����և�{iSa�/.�f�T�V�a��`�=�34�A[�U�(���il�o&̀���u��2�C�J��x�5�pW�0���d�_�Gg�)��5�oM�����ܜ�{�s���g��ay3��_>��{2��d���O��Vm,��iu��r���ʨo�"i-ؕ���|����
k"]�'����6O �lF����� ����7�39�v+�gKM��ŝ�¥����dS�/�v�+β�8-&�[_5�g� �+�$��A%1a�n�vx����{���z���L_z �ۦ��@��Yc ٲi=��M&������`���ξ�!r�~o'|bF�kq̔}�fX�����G��Q4	"�&7ƻ�W;��5:�}�t���� �D02��~��W� � ����W�[!��cj<�&�&j��;�I��G��:A�����<^���L%~������u��� GR�e*6�
���S��d����bSG��3S���z�D��=��7;��O0�[l��Cx����\qy�s����N��jp+S�s�Z�vidn�bEN�2V9���u��>��a!�1�V����L�xp�	��8�wnoOB>�X��<������܆)��;0/�4��7��j3�m�l<�t�* b�ł	_�r��D�k�_@�>��U�\���x�{�rב͎�� !~A�
�R�;����c���|�x�^�|���1 ���M����P%	�
�U;�ՑEmŢ���b ���v�f�hC��A(�W�]�O$ ������S/�S�n+���Lu�V���K0Yr-����/a�]v�퉚)b�ZEm�C�ps�s˜�� !�a��T�W:�c��굃���Y�f��蓷}m��{�:��&Q
�z���9�
�:H#_Y5�`kL�x�:��wnS_ykL_�=��wΫ�oX#��,~�]�|���[κO/wN�#�� v d��5կ���΄a������Aa\&�'�@������۞N&0{cPƌn�i��~5Liw�:��p�����3��s���.e��y���_vy��,�Q�|!�.^����b`95Y ��*�rf(�dO:g͚�wuwx�����wlQ�Q�id�tJ��+��/�����u��]�8en�7����I+�ٚ:������� ���Gy;�YJ�܋�0�ƻ�갭�:J�w�\ U�T!���X*�"D�_u���ú<��ndI�[�ދ���_!M�y*\f�}�G;�ˌ,�*�`�מ��X����
M�T�����I�-��ck#��m���#�qL�c�f�	k�ҙ��ox�O{��S7q�/����u��G��B���{��|+G_�a??��I�תiݶ���v�njԞY��׌��~b)�E�.�(#�; }Ϋ��bVU0ߖ3��G��6�7��a;�P�4�y�\����n�E[���A]\
�����E����ù�u:��UҰ|���$rsC؏�6�5� �e*&�x8�yU\��B � ��iE�y�Zq�H~�oX5¥��5&d�ky*�w��w(k
��X�UE��V�4�Nۨ��;�$�@����	9��+��]��J�J!��HHBhV�OH�ȡ�VD�Q!�X`RD�HPz;��ϻ����y7?��]N��"�������1'��$i�C=����7Lt�}� };�\��/{�]���w��s���Ǒ�#��������̿�[��
�9�n�z�	��ZR�D���ˣRx4V�4|�f�z�R��n<�[��'��t[��t@�|8}!r��K���F��k�3��i�n(u��
r�Zp�ϴ���5�$o��!�K�R�t�6�ڽ>�5��r1�xz�ùkr�҄l�h=�W�Oh#Dr�t��y:v�(�iW�AT;��2��=��7f�;�T?�S�;�d�]�s>��I�@E������0�9<�[O3bp����c��� I�H���i�7:����7ۈ'�9�J����.�78�"�z�@U��Ϡ�/��|�8 |���Xfw�E��%3�^�=[{���	'�Ú���ͻDQ$�s��Q�5�$�8��u`g�DG����2�l�ń�U���^��O�� ^�W<Q$_'>��Nu@(y�"��Xik��i��z��sXu=0�<jC�G9�����1K+_4����ͯ���R�5��ޜb+�|�Y7΅�\.�r@��e�l�8��}��������_�v���]�Pn��,/.���V�85� �{����ݯ��els����l�XEhk�;��,(UWx
�Q/G��ԟnZ�\��oW*���b�R��[|�4d�#��6H�����ޏ��Ds��?#��2(C"� ���| �������o����D4�;(��q�WC�k/)z�G�A��#�[�3?�)�h��A��<F�fZ�u�~�>�HQ=���69}a$�j�s�q0���'Լ�Dv=�x[ Xֿ����ۑ;�ϊĲ#�&��K� �i��#k=Mz�K�psT5�~�dCX���~5Lm��g ��Gt���k"�p����M��ˆ"i���{�g��vPk�&�p������g1{���hT�B�(e�R�]�c6@ �v���[z7;ԨW4��a.6�9K۶Ma�̖����ϹŮ�+�蹻m�+�F�{��x&_1�p��4k7��7>>$��?`��;~�k�(�aJ����P��\n��ݫ_@��2�,��o��J?pdM�tj��4%`��C�l�}�'�ǫ���:룱�%���l�n�~��N�yn��W���$��h�>a��_�SWK���X���,)�$,|)Pm�0�����;;o�j��;��	�s����t,�~�|��0����ϟ��g}�*qF&*�sl]iVz�j��2Z�K��/={�&���$��Ƌ�	�9���&wm�h9�4���ڜ��U�6MS7I�,_���1��A�KY�2��Rݩ��\��wˀ�{bR=}�qch�F�0^S쭵Ѝu��n�F�O�n���O-��Wq��nRf���l\�_o.������.���zG����ގW�P?#
2# dpdVQ�P^B�~9�~m������ ����(�����a���r�ߜy�m���¿H]�7H�`@���-Ok;B,z�]J�q��2[y�`ۯ�D66y4������K	�"���&cgnP3n�Eo�δ��Q�'��%}�|E�v�>�� PK�6f��� �'��6�&pR�<z/˹�>��\�}K�.�<��=3y��7�Fb%Z�,4�qN�4w� ��6�1���W0os�`b�g~�a~_. 9�J9\�����G��b�%<�v11w�)�ZQc�@��POԘ3�mp����4ѽ������S���XG lF	��t(k
��	 �Wi��������L۬���'�v��{�y��ϴ�>�`�e�┻�!�,�@�J#�ZVk[�+<�� 	���\��6� J��I<<f��E95��&��{>RM�v-t䳵_ӏ�f�`	�ަ���Ҫ�x����k�S]�]p y�CB`�=�����|�Uݎ��6�Vc���6|'�-s� ��8�f�w������z6�Sݝ����r�4يd��5>�N4k ��e���u3G�ެxW�2��4�kS��5�M�<0�B�o�k��4�̧�%�k�5#�V��&s&���2������I�3�G�F�֨�r�Fxmу��_G��)˫�e��*[]� �I,�����q0�ݻ»���$�1wŢ����W3��� ?�0'U`D�y"�`@x�xxMl�����	�s�[�(���E�o����#\c�/���-a��Q��&�f��׭�8���m�xzݤ�gG[#P�1p����O��x>9�3I08 <��������9"�81�"8�~u�O�C�d��3��,D�8pC�Z�->{����l����IgP�Pd�����d��,����i���Cm[r[��lӈ9�����{�N s��N��2�*���z��y�Ä���ݺ�%�j7�[F�i�
�4-9�����I�@Ty��0ǵ
��+\�2�';Vd��a���a��~f��Sh�A$�ȁ��c�>��,s�N��8�V��=ݩ8En܌Ӭ����T>�]3M��w��K���9۷�L{L�k*=}~�&=-DY����J���=����sR�V�O��rb��u�#�U�E��H]#�Zr!��[kN����<r9��j���^�Y���R��:_fz���:k��r�Vl 8P�򄩆���N�.]���>�κ�ḯ�{h&=�{�.�4h�&|x� �`S��X�G\C*�(�[��:�8	cjU%�2^�ؿ]�{�[�Yv�*4r+��7	��:�����v�y�#�M��<�A��.��|@��K��/��hy�C�5���ˬɺ;G�e�h��m&�G4v���k���R��ڜ�%&G)�4�
ջ��J�P>�EPS�AuM�b�A&�">F�/���yׅ�<�9˝=s���'�d\U�t0 �(��<�N�������=(�c���O�b	�D}�DF9�TtD�tH�/��2Wʉ8Q���,��|��^ �ZY�5��
;ՏȃM�{���|9�\��g�hf/���\�k�Y`|��f$bAP�L����싇x* �~爇������|�����0���a>���uz������-�Fm�vy�=��n��ݼ��*�.[������Ҳ��Se��b�,���e�[0d��N�xV5��C�=���^�*f:����5e[oL��L�f�l1�y٣����� ��ށ�x�]��M0sj�}T���;������[��[����V�E&�m�fy
�t��[h[:���f�K�!c���k;��v�׹���53��#�}�s"��e�i���}�؄�+}C,X��Īq$���s�>�y�ޔx	ְm)H���W?��:��>�~<w+ͼ�D�L�n_��fW?Ǩ�,~�����0�C����H��FF���'���഻cW���%���u,Z�Ɲ����Ξw��DD�v̮��2���Lo��'�\�7����X�j��[�au���F����3"c�-�pa�7����ּ2$�f\�+h��׌�\w��j��K3x0�O˻��c���꺜�b�l�C�ւýF�8�����ͭ�F�0��w�����I����t�����ʉ�0�# �ax2*C ��@��'���w[]ǅ��&���+6a�|��!�c:�5g���}ʁ�[T�N+�x�sl������ව}����zu �w�q�(M'����3h�2Ǜ����0K"{���r	^��v��\0�E�wD���&oe���hF�`\"b�_b����` ;���h�j���^���6��w�-ga�|�P��sL�t�����)ڣ\x��rXʪU�i��	/�`@y��s�V�I{�J�C/;��Ǐ�a�R�f`ؚ�'$�dq�ɮ;y��� ;�>NH>�ˏU�7��?1Q��0�ƃWs�:dci��/�'��e�3����;����.���Tӹ*x�vG�g3�mz$o
��V��R���P:�l^7�[�  J�v�V̎l���{�p���W���b$�'�4��D�+c�h�cǩJNXfm�~d����?��&�����.e��J��y���oƇ,�v�����y����EO�͇��Ӗ�{��;�<
Y 3
���2����sq޹Dx��wz��zvZ����<���\�K2���v����f�smي
�nEQ����ʁ�f�GZ��JY�sV�U�I���8h7/�LOVIvp���S����E.���e�e�%�M�R�qYUв�eY��L{:�gN�+i��W�L��;�d��ܩ��.%t��X��/���F��(X�w%�QU]ֱ+��8�.�v�,T�	q��Є��d��o*G�e��:�@J�]�.'Ӏ��ԫ�澻�_wx�t�dJ��Ѩ��:O>Qh��@wDK�p޺�ms��zZΖk.�ܜ���{��6�+�z��YI(����:f,����[4���|&N�H
t5�;f�v�;�a��Eǅɗm�������͒�(@��B���W/kK�:�g;V�rr+{�=��ٸk*w�Z��X��¬6���F�,^�����[��E0��mY]\��Q�;j�/j��wp���}�6k���.����,�QN���ƏVJ"�O{; ��gS�D��PU�S���ה\�r87�X�N�%��C����Ad�:��z�ioM)���ee@�"�}�*@-c�]���
Ȃ�I��3c;���l�@<X*S���tҩ�Txe� �L6$�>Ц,]�3"�%ˬ���B�{���f2�%���:�"�A����*@@�-m�M�tM�Z"P 	0+�UB&bK�S�Ɂ��G�o�ݩ�K�c���,�{�I{��Êb��J����f���u��۪�ڮ�]\{"�����Z��]u,�!��QF�9t�g>���R�2S5��e�B���5)j�n���*]vm<�6Y!�:�b�ϻ9d>;����3n�(�m�V��`�Ԩ�-mtΡV�r�ؤ7�;�R���p��w� �]��:[��:��nk�u������7��C���`z��tn�4�k.w�a��5453n*��:���C�5�M��rp���]
IJ�£��)�㬎c����W�[����Hpm��ȾKoT�V鬌;���2�P��ݠn}��=�?��v����)b�ؼ�eԚ��59܏�_x���
���h(OsgN��*�߱˚^�PL��QI7��ǴUu��}���[5Ծ�2��=�N����M5�y:�����!��Wգ��7�%���v���H�;oq��s�k��&*yϦ�:���_:^�u�ۏUf�/��ghQ�3�q�ܢp*@�N*x٢�݋r�V�BȲ8IOH�I4��s��]u��j����'x�|||.8�>�����o��}g��]�ݮb���n�湷#\�v��J�wQ|�<x�돎��8����񟙾�����sֳ�$�cr�wD	r�77wN�wt%O__�8㏣��>�g�;�m�Ɨ;A�h�����uѹ�I����8�w����v������8�����^3��}�伎s�/�\�(�s��D�wwSʽ�=\�S�G(�	��������8�>����~���Pnq^����}W>�cW�wPck��<{{}||~��>���g�����)+�H����;���.��x��W&�X��^���lE�v��E�w�㻶x�\���Nn�g�7������dstZ�.r�����m���p��vF���!ˣ~�Z���������wn�Ĵ���53��V{�G�c������ǺJ���ګ��K�K�;1�v����%]�)~�p|8@�  (0�
0�#�N�%� D��t�~48�/��2?�1o���;�q�t�l��b50r	�W<���n�}��ӕ�q�7��y��H|��������|��ُJ;�?5�`�Z�+nM���cdE]��dO���z<d_9`�)�a\���Q u��a�X+�E��`P�q�!��_lh���#����_3�����ӟc?��`��|M"!��i!��w�d�hC�H�B��>�7Y}ߓ�t3 ��A�$��A��-���Z�S��"�G�����0a�A^��	q�8c��|1Y9�@��.�n�ĠMW��S_��ŏ}�b��0:�q^��bI�:�G��pH��5�j�v�d��.�����k����"�� S��U�O�,�졚���|�f����'-�VzT��n;��Zٽ]l\6���������.�c�����	��,ϳ���2�>�� qr�B�}��8� `��׾Bo�ޏa�])� �&��6�N,���H<�S�7f��nr鑑���񟟏b�qû�����O�xۤ�'��-B��q�}��x�=��#S�SjIy��Z!��
�o�^Ё��#�m5@*7���	u)q!s��S��=f�C�L���:wo}<���Ψ�d|�3]��'ʺ�~���a�Da���"0�'@��=���~?H|>��; ��o�/������TJ��4���Ua��lu�`�'
�~`��=��s�K�q��PJ��.��� �ޛ0���%�[��E�P��<��_s�|��M�Q�$��|}#���}N4�ێ�ޣ�g��6�P�~�=�qg�=�7����#�{�}�8=���~�jS�����cHb�XJB��6cBdG/2b���e��=֫ۮ������:��Ӷ80gu��m�r�/��L�u5q�ϭU�-M�كs��Yxi<9d���M��8b����+���z@��,|��K�������1����w�qhO����Zy����oF��<#���
�U�����
���v�&���qFct������vw��tp���'�K_>���k7��s�9��x1�������<a��S����"M6�U�\������3�<�f�+�Y������L����P�.:��#:�:�)+��j�H�Ht?kO���i���2�P��f:�(k��-O�b<{����!W������뙔3���oS�U�=bRO����pVDa�Sj����|�giKai���'�ʒ$Iu���/]��a�e�iȁC;wI�[�O��XC\�h58s���_��A�3.�1�n¨�����N��h�y��2��Ò��JfL�#���ȁP��	.4ZO�@ԁ�!)�Q�gw\﻿�U?A�N� �!C�"$2 C*%x2��T�}ߞ�z��H�I���<�}=?�����`���(E<�c�~V_��_g�\��(�:������V�F�\��߄���]91~�L��0�H?d����U�Lֈ۟�xz��PZ����1@b�D������Nv[W�ی�q�<e�%��ؒ �UQ,0$0��&��@QY߾������Ǥs9D�a��aI"�{;=H	\� ӬH��F4y���$����Xy�E.��D���	��4J`<a��'�Ǭ��k���\�}[`cE��=���ۑQf�S�ז������$�َ�����o�D�l�@.���lɈ9c{$Kq�^�ࢯB�9ʔ_o)�h���Tj�|�7��*�ˎp�i�c���2���hL��a|����bs��y�<�I�q�df0�e:6<�0h������%臄���C%t�j��nA[��nm����z��G�ݚ�BϺ���#���o{�T��O��8��HmO�M=��:��<;�(�8�㩛��؎l��#� �T��
�;��"�TG���q��w`�#{�g��KF��jR��Q�6�ft�ؒ�6��o�|Hv5��v�f���xOo��k��p��sO���|���ެu�E�::�˦*PXl�7�I箊��1���Ul�&��]��A'�U��!�/��
��ʩ�
ҁJ�=�[n{{�����C"э�s��P d?kmw4�Ó���K��g�|(�J�z>�t��B�<=�ܵ�3a��W7�N>kNK��;��z�m�8V�noC� ������[0�퀸�|#��{S�43��/���C�ޗܿ8�{�x�=�j�\;�wg5��[�X��d�3��V�hC^Y�[�8���_e�j��>։����Cb�Q��Ş֓�����ý,4��$�8�`:�f��B����1��胰�u�Ğג$-uM �k|�{Ba�k�K�����>���|T	ݚ����A�G��f�j���:��D��H��`}�
�|����'����vڙ�5�����	.W�^��e�Q��"���k�����&,�4V4��ķ��0�C�#��=/��2�F-�Į�;��Y�,���^|]���跮+�#��ʸ"�B�r����W"r��b��E��cm�%LIqz�-�{�$���璩�4�<O���U$m�ʸd�R���>��-V��;���~t,��Lo���u%�>k#�U髰�%��%��T�XF;Y��dͫ�21��Lë���PU���2Ȯ�tڜ�717�0���O�gF3���R��s��>�/��0�j}�ݫ2%k���.��m9Շ�E��ʇPPdP�@e 9H3��,��������9�M�'�z�ûFKZ�Vl�X	� ���α���7/���5��<c��e)\�+�����"%�	�B��N��]���d.$�e�����O&��	�&��c���R%��5��.�u�m&�����k�q_9�Z�7��K�\��q���kĠy{���\�QV�\�ʬ��e�<d�{}�gI`� ���t���H�bp��	�d�23��@~O��
�����q��gͻL:�`[$��b��o�5uCo�C�b�S���(,3��UO�i)�Y=��8�ڸ6|����5�Ŵ��-B�����Bף�v<���Cz�Ũ�f �.l�����l�WK��f<��hU<������/w���(��n�����3t���09oW����rD�s9% �^�ܭ������χ�-  o��g���P��%#
M$i �N����k[+�,���>�|��o�@$
���l�����Z7��1,���w`cE�@���7��ʯ�����ls'z��:�=DA�-�U��u��JaH@&�68zh�xo,�I>��
�Z�k�o�������tlb��x�>j�JIn�q�x%��V��W^�Q�-�m`�p�װ(�����k�om�}�V3�;��g*��[�Dp~ 0�C#� ��¬0��a�1�I�6o�!�y��!���̟,#��ܝ ��_H���_���к8�;*�C5�\:�z���9L#�8 K�VU��X�#�	���
�?|����W;�|�\Kǹ��OB�.�.����������l��Q��Mc������jb�<�'Hg~B�u��(����;�-	G-���#�x���ac>��-�t����n�;�Gz3��/�\�|�>�l�@����Vx1�wC���^ w����.�@����L��alC?"�Q�K��
�J�mj� �W@n��؞	�7�m�R�Y��"g�w,���C���+��
�����Lk&`(���m���@E��e�N<y��ODM"kX_��]���ᱍ�FMP�ѫ�7U��xw����y�p�b���H(]��
X���z�uM^"G0�I;{X�T���}�V��ߝ��5����m��c/d���Un�z @�_�/L�|��e��qP!�y��Vs�ۇ4�i��>�YP�1�aE����c,�l*����h��wy��tZ�4_�[�+nG�����<�`(�=�W�w[t�(��v��tv�
��b��&I�P���z�`�V媓��dv�{S���p�}�`�Y!�s�gZ���8�T�G�ec3����;��a"�}��^�Y�����a|D��L3,�
�再9�;��^>u�\9� ?��`BG����pa@�`S�z�fd?�D�Կ}^�pt��+���R��A ��`{�6:@��֑����#u���x�i�;�ۍ��3�⅊��E�����1�ܮ��V>��m��i�{Ϡ:p�Y���M[o��A�U��γcc6��{�h���a�7�&o���-��@Tx���t���k܃��2�(5(�N��%FK
=}��Hi8�0�g�~�_�<_|oMyw)�o\4�ʼ���^V�x��1-�bm���#Y������x�Z����*�Qܛ0P����Σ�#����q�M6��Ɉ�Ҁ��ϘE�d�hD=򖉿�]Ht��""�Q۬���(.��a����}���Z<���%�$0` ��z�XDl)�J�G�*�]��D�9�NȜ?�-V�����Ab"x4�ߘ��FM��c�X>6�r�X�}J�,��x�AD"J%$��x��O�J�}8��Yӟ&%��ҢҖ"OL�9;gz�s����m���;i7���"�Q�;�a!.fM���B#�WmL��#�Ȧ��7�{1��߬�f]Oz:y�U�4��^ʋyc+��RT0_s�jWXy�N�h��ǦY� #���uW9��D�O-��ܺf��|�<�ENW�-�e�w@�CV��t���[�#�������}w��ww��զ�T?#"�ʇq��9*pdR�8�  9��λ���ݱl�`k}���y ���g[�����^'�{�����1�S�R�5�Ϯ��Z5?�0�A1T����;�񮯩�'��^ؿ���Q�["��r^�Nnz(di�~��?Sp�G�E)�+�ȿ$r��j��X-D8���3q�}T������e�?�(�#Fq��h滤�q�u+��
�ȍa8�k��H�zE�Ǫ��~�+L{��BP�+�^~��e��c���ٴ�n��p�χu:�#i�?^u���V8	b+���|�x`k�s6���Y�厮ꌗ��q���u���B�]�?9U��随ٝ������\�O�� Ú��l#��$��׏n�竟��䢅Z�G8�'��n!�u(K;(Ts��nsX��Gz�aV�,;Ƶ���9%�k_23�a|�_���<:b�*��t���ǞX»��(��䀌8)&gM�o�;0�i�JvcA�����d�sH�3�]���q��pFl��N�������5��Z�٫�{�{�R��
�=�MəruX���Yp]IBuM��/����Ewa�{�����)�QэF���b�Y�3W��R%.�����l{kr<n��99�,轺��KH>��{�gu��|�8a�Qq�d	:A����{��+��XeXd�!��>�@�6�_"���{� ��+bl�[��*=�2ޫ�.�ZN�2Fb�^��æz%� �s,��<4��������G@� �ߘ�����۲��ݝ�KY��t�_B�.̚�&��{��:�3�Fp���!�ɜ�0���g���n,\sh;�cP�����H%O��RS��![��q�a��"<�)8���`��$4�|��p;(�y*}w��&� zL6�[,�O+� d����tڜD7�O�%˼yC��O�����oFy��k�h�f�QlU?+�X�熢��e��DkBd|��!]L'���g� �����ܤ�}���b�)�X�IU=st�w$WD8��9�=1�[�z�n�#ͤtԉ�;�f�h{�F;W����t�؝=�;І��}깄
�R@�C�].-���bG��Zkf��?�L�j�V���CU���7n���ۿcxT�4\��4cY���~�5i��z\�e�����V
坼�7Y�n���bn<�K3���q �=�'կ�����s�n��K��M�Z����毘�͐���p4�z�&��'�������x�����M���K�Z�m���@m�������|�w�)�I��6��h��]��7��'��9��kY{��uqྫྷw��Z/��p#���p�a�a��+��!�a���@�� �vͥ���8;7�ٟQ�=xEoPvQ��2�<�l�y�0.�|� �̎[6�*�D�JfxbA�<��+�����Vy(�1f}�H�3���@I���廏��~�}���ɜ���ݧlK:�I(�&��k��>Ϗ$�R.��y�J�	H��I�A�o7ͻ�/ι�ZK<gK���e���s[y(���X���D�z��-��@�� nY�I
�����l��$1.����@�{�d����yka���Is)�i�H�����UL޸�Vrt�4� �2O=��2����4y�~A�{�}��qT⎀|���6N��X_7���=�X��(bz/�4�;d����m"��a��C�,�>k����+���'����x	��1KcBc6jAA�t���%�8�98Wƌ�ߒa��pxc�Ս��ε��u���s01#��}�1�x}TڞU8�HB�Ky筹���ť�j�"1i�e�̟G4LL�>�����.�=}����
��<��-��W\Ǟn�"�M�sQ�-��Ճ�Ѭ��1H���:E�9x���)�Su�z�f	�7�fG�L{�s�M�Kr��Nq��(��.���l7���	�y�ұ��/e+���HwPJ�!I�0Cٵi-���٩���-�3�u_�T�g5gR�1fgk.�K��+�=9z�>&�;5���O�/nֶ$�o鑊�4i[��,��9�:+Z�t��޼KOL�
`�*T�;:�rV]�݊��V�M���\��
q۝a��]q.n�Z��k�*�\����S��_U�S&���ֱhHr	ϣ}�0��ro���a���<*{~���Њ�*�n��7�WZ(�+��p�}1LO�(�Rc�L7&�*os�ppuwPV�Ι�P��]��JY*ƭ��,b|�Yۋ%�!d�b>�/�8(��c	�I���ėb�h`æV醩=�hD�Mv�{���^�����py$�86	���z�`�M�̻	���:�/R%�	F�	��v	}&q�ݦ����Y;Dt֗M�ukø)���z3�,o�Ʌ�)K5��wI�&��4�M/�p���Z"���jľo^w+]]E��^��f͢
�@F��r��+�V�1L6p�A�(���쾊V��Ht�{���u�B��J�h㍱I�J�$A]��3��`�;�<E2�`3��V����?Z��D����C4���4F+�ƴ�@���L��`�΍�Nk�*���$ɢ(���s��b�f�؁ѡI]�@U�L[�:�����*T���INJ��Kp��@P|�SuZr�ȸ9v#����ӓ��.�A;���֑�����d��H���w�"�P�ck���+��òT�+o���t]բg*F�A��t��ɗ�|���Fr]�L��hs�h��QQ�}rQ�|e�ϕ��=��T�z�䍛c�؁�ՂQ�kH�*�>�N<�$+�.;��C���N�x�>��Hΐ9VliT�����ݝo�-_<�KM���̐Σx%��4�WX۫*�Σ�J�u�Oou���9�r���n�v���Ưr�4�M����50+:�n�����Ω�04�!Jk6�Q�;����y�7����2j�Y]	��w�ɧ��Σ��R��b<�fM�Ҕ�m��-�;�5��U</(�I��I-ܓ��k(s��c�=u	�H�O5(�����A����h�3�JI�%a��rhy�Q#��x� 9��oz:���|�o��m��_CY�߈��3��[�ޣb3�P�WAQ��z"��g'����W/��Y��jm��Y*��p	t��RwoK͕��'cq��a��5�˄��$FQfL	b���CA	�4%�=Z�TJ�)�_����L�2y��X��%�"ԉ8Ą&ᆭ�H�M\0�AH[��E3�L�G$D	"2Ĳ)���)�L��JF�R鶙��I�.(D"�a;H�* ��PPe�h3J�	�Ģ�����J��)�$dĸ�tLi1a�a0"����$��Z%��#���x�Xs�(�I$�W&��{��Wg��||.8���Y�G�:zU_y�S�����A��/��^6�䈃.�y9�I�z|}|||~��>���>��7��$���o1D��dw�8�w�7C&=+�us��9}�D]
x������\q�G���~���}�>]�z�L��~��\���_]y�\�n�4`�9��x��㏏���q�~��o�������8\����;��$��]$����ɓ$��κD��^/���s��������\q���}f}����0D���'p&\�n�s�I7��3��p۝����zq������8�_Y�G�;���ɗu�$I�p�ߎy��t�Ē����d����뮅�'wr��Τe�I5���8nCӋ3������<n4w[��w]���n�B��� W���$�A�u�rL�������a��q&�a����
\饔ʐ�Ӷ���ⓠ�,G�`����r��D^�����v[T��������ނ��AC|R�$	G�F-"�H�!BB ������9�p�u�!�/�d9��a����B3�Ít{�ֱ(��I �&b�*<͘�<��q�����$}2q4ּ��Ո���٭5���7Q+�݄Kz�e�^v���q��Fy��q��#�&���o?j�Y�A���خ�	`&�zh�ˋ^h��ʬ6��k��tx�au�/�����\f]�v�2[�ǈh�z�\wB��B�/��rK���ـ��y�f�8k�h��׶��5ˣO�Ub���؝9D.*t�i�{3�"ӖgdTw�L��rG�5�:Vd�����vF���W@�TGdi�;���ٰ��aj���`Ldd�2Yszzp�]$��d�fa�߹�CBddC�$_�a�׃����Q{ �N��Ym.�VǪZ�[����pLO�	��%���?&�<�4�5�������=&�n�A�㝺�qVg}_w�c$6Ye%&���ó�eWk��Z+8������B!�Z�QX/�a����v�q���.:�,�ic���5oP��N�++����`���J�=���C�'cN��而�d�y��_������tc?^A��R��	y�Z&��ܔ��
t���!}�y,-#o�pڿjb{=$�j?g-u���Er!&hw,G��)3�9�;-pt�c����EWf�;���(��!����Vv�L�����|@7	@�ޞ�H2P��4o0}���{QyW�K�q!9���e��-�;.צ�;7�{�em]r�j� :ߠ��|ШF����A�u~t��L���r$��\�WLe�y�����A�ȗ�:��-�g�"8����QK�X3��Q�E^c:��y'���K����3�;���i2��T��u(;��(��_*�|��Z�t;�uz�벓m���w���"gr-�ΐq��� ;�K�Kb_1��Zҙ��!}cK�Q��:�j����7h�R+`y ��]�9�Z\O�m� �sS4c�A�A�����/<�$�7��e�-���F1f`K�Ł}Ą����j�@�JW��z�l�*�v����h��z����U)���Ѫ0��~$�H��S.�8F���f�s^ �?���:�!T
1��l��TB�h�V�����O�v�C�.#2���ͨ�j��sns��\��m�GȯR����}��a�F�=L� ��L�8�{0��s�O6G?�J}M#%���̔��{���=��w�h��M�q�]��ϵKx���JWV�Ԝ6�R��Z�(��J$�}�V��W��#!~��w��+9����;;Ԩ����Kb\u-�K���ft2��xe�{���7�8�� �J�eda!�9 ������������|�@�S�`�f�]����y���m��Z�B�U���C	�5���v$�m��Hmõ�1�����joa'�2�2��p��
ߖ�Ah	��*68�����U1��)��w>&�I�,7�E���OF�����ܶ&bo�;�?h������lA綾����ў:��4�ڣ��s~]Ҟ�΢s`O��$>���k����s�W�] �n0�-�9�s��U���ϰ|�}�����g�m�xJ:�=���M������|t��uz����8y�Do���]Q|c����Akm���t��K�񾍙�T)�گz1*8I�yc�6P���i<P*���O�UZk��ߞ������#L���ƚ�]
:�of��$ ���+�ء;Q5����8�y8�m���C��͊��][h�]p�E��{T\3՞��g}%rGݶ�A�}�ȇԹf��[ �=��Ǯ8��1�I�x�)2�ۑ��
�oٔ�a��b⏵-�Xţ���w �����hP�9��]��o�����|��i��$�s2�x�a���.��ݫ��.�_�5�w�ӲC��.�]Iw]R�a��y��6��f��,�hA��v����ÄG�."�2�$0������{�n�n�4����Q��V��I��ǒ�8�W5��P��>�R��_dt�	�UlÏ3���2��`/,�?'�e�����=�i?���9����j�{c��*�pu�`���tcD���sκ�4:��T~$��9�t��F�^���8��G5����i��kF�f.���<t�K���s;��@4�j;;|�ݜ��x�X���=5W��5��^�����fWm0"y��{#SI��[<�!�N���$����P��%�ѹ�6���'�����̹�}|^דP���xlu�:ۧ��_o�����6����Ο?���]�tv3y�p�4��LAǾ9��6�u�Zܞ?=������{*Q��QaK�8�#�3 n/@���ܹ`M&�s�o�p#�����o����x�{g���l#5�W�&0�@�M\^D��v��s�t+��}˞��s�Z�Z�Y�ty�2z֏+ҝsa8���])���՛9��p���p.�B�ph���Y]��:�����.TE����ݷ�*���+x7H�<�ز"
��B�<�^uk1�oާYJE�:��%����KhNs9E� N;�9!�F@P�u3��\�$�'��FJ�T&�	& ��Bl��% A����w������	;	�� 8x(WR�x�m���}���4!�Å���V�������}�J����Q&r}"��@����S���C�{7{�������5�ZA
�F���X��'q�܂�v��5ևX���T���n�7����]����|'.:��8ﻐNW�6�Ĭ��V?`VVT���JT�`0r�3<�����-Wng�N�|�z>H.���H�U���Uv[�;)bp�2��o4x20��."�d{���G.�A��1�����]ոn�{�H{�3����On����f�_�2�GAq
�>�U(kn�1�R��"c�ZI��si�O�\Y���ɢr��� ����ֺ��1�\�F�P�1jȊY�,z�Mb��u�;5�dc�.q��6���'��/��d�<�E���<ȉ'��ճ�����-D� *h=6�JI*���Si],�f4�{!f��^7�(nD���kJ�%����s��ܫ� Q���qw�h��EQQ���~a���Ƹ��L������?�K�`	VԈ�Ύn(w:3;�[����B`�}��9n�)�����z���|��pmn
{��8�G]����`������>�b�3uK���x9N*�T3��+�KVm"M��఑E�1�\����s������X`�!�j���c����(8	�s�����0Л��a���$�7��uoz}Q�=$u5���G%fv֠��{݂�2J��/�pCjz�?�P���,3��g ſ{�� dt�G0h��㲳cD^������kA�U����q'h+�a���Oq�Y��-��KY�mu�d�!��n{V��0�#طW��l�g���yC���L�g�<\ǣ�2��{:5��Xm�����`7v�������Fi���"dCkV433�_'_�69��Ǧ:g�ճ㖏?R���5c�~���ߏP�p�}��|������k���J�~�k��BЯ	'4Es�_�Q�ς��S�%��}&���l�8�D���k'�[���׽�t��ӿ1Y�N<�s�vp�"�Q+�;hBO��`֪��CV����y2��1x�������ީ����u�bL�@�4��ߘ����Uϻ�>3����w�vT�f*�g:��{�
����e4��s̴���7��74y�2_ڜw]��{��XR[`�n���d��z;b�`��'^/�Ս�Vt�䃰4����e�44�u��ݕ^4M��Vhm6���\n�s�ةۻ�c�97rbs�K��
�*Yc�}�-��R���/����H��k�[}"<e�8G?��bg�^Ju�߾}����� �*��
J�=��Outﱽ#�aR֬뻢j���E	B܍~@�7��[��3I��6�Xi��4�c����V�GJ�a�nSn�x2��2s1d-����� �x��C3F챛΍��eC_�͝���tD5N��4{3�	��rInf��gv�����?��Lyێ�����/��Z�m9/Ǐ�ka�g�,�Y�'{���w�AE[�ҁ�t�}����7CR�mX-5��dH/,���-e�r��ˡyF�X�����]U�G.!��i
��v0�ƭr�OX��YC�P>7��>=Md��͈�Y��9;s�@�����1k�;,-@Jp�OE&�b/�crѬ�s��r��.pØ ���
��ö !qz;�����m�)2��M0�B���=�M�E�2Y����+�ds�D
�O/�N�lo9����u�mƀ�Y�������Iѹ���E��ݸ��;Z�4���S��l�5�a�cD>�3Mxat�c�0?1��_u_��(ײ��8���Q��u.^A� k�|�0M��.��E�"1�
������F��7Y���6:��Q�UQNq�Ya�|�����)���qqSwG�k4�,�8V����2R��`6��O����p�!a�G���?�c��K���s�p�	mn��S�_1��g��&e�
7hk��T�y�#�O>M��������<�R[���ƱjA�h_O�@��=�8r����{�Q&3�؋�}�˝�^�[ҚD�L�H3�Y}�;W@�_�y/ҧ/�¥xn}��َ"4z5���+�&�6����;1�&P���㱬�L�"��2d�T����O]�Gy\z�pQ;��~���*O�)}1��P��;:f6��ye�|��AJI�`$w]���c�y�g�K�*v�&L\H���(w~�i����qs~{�����W4�ɬ[n���]	�[ڂ�ϸ~�s,v�w�e��v)Ĭ��CK�с̈��:|C�?2j�aO�'h슧�J��L�*2�@��ӱ�
�s���.�D��|d^��d#>[���nܕ:��"��w�����6&�ў�����S'��E�ps����ԛ\�l����{Z�}�T�`�T����Yt����H�)�XO2�k� vǝY�����!��t��s����t�*< 9d?�����b�e��Y߶>͵ɵ�������M�#[D퇈��SE]�zC�a$�N� ��'�Zm]!-r[\���2ɕ'��ڝŎ�`7�j��j�!u2
*����/qu���{�u�&%}��˺6��,$�(�e*I��hC(�
M�d��d�` �����Vn�*Yr�.u����������3>��IR	��Ϲ|>k���m���͎���@�k�}� �L%#$�w���¶X���h�V����/C�.ܠ4tDy�l�I��O>�gG�5[�I�����.L��X�����xJ��>�$��7���w�@��("?+"Z�����\H#k;��bjC�����wD�p��=�ak9�8�
�N��|wOz	4�煿�|��j��=|�h��m��Q�� �f$gd� TV��ƱLh8c��;�>���};σ�?c��{�p '�����jޑ�A�F��jr<�r�i'�x6�w�4U������t_1s�ޓZ��oD3������sx#4�⹤gq�uC�V�uf�!t^���C�y�I#H�|h��1l3��s��\�n����HJl�P�~'�(2�ZRܽ~��3��CM6��b����j@��J�N%Dߚ9�n21��t��S�D��U��gm��w��n	�����,.{^�*��4�j���bs͒�!��
����!�w�nG���5P�,Ƶ��R1�"QF�/�|'G5[޺�������,wN`�O�u�uw��{�0�!�"+{*G�}�1Nr��{�þ����U`#�t�g&��f�Vf:�&pԻWuH|���u���#0C��p`ĒI�M:�{��c�Й���O����QFݑ�ﭞ��Z��2^6VL��Y�l�Q��I6�m���ɤ&�l2��B�T�j�;�#(��R���v;~ϼ:���e��iG�:��i�r����ހ۾��dQ���cH���D���y��IS�����*�k{S��l��g� 鼡Ѿ�f��tpS��ϵ���ם8��/���Ќ1y�y;�!�@p������4	�5����0�7����k;�`�,�oQ�v�YĠ#�#�1x*{�	$ϛ#ׄG������p�l��f��h��ӈ�7�J���q�/��L"X�R��$����O���ajdy�^N��ā��Y:"��@qϾ����b0���e�&V�Wt����:B�G�R���d�����u����~a�S�YCcs���9xn��o4S]]�m�L0|B�13�}��mj��t�I�ƾkz��Ry]����)��"�y�"�m���{���0�8Iw�1� ����q����	ǖ샕twZ���Np��
����eREX�3��+�8�f�ш��tn����vC'��Գ� ޮG��j5��7Cv��Td�N�r�U�$��-@��r9���V,�=�MwS{| ����px\�O�L����b�d�!Tr���v�d��ù���� ��M��ej(���H
�KHbn_%1��}l�F�j��̭�������c�j�MQJU���k�7V-���>���N�ٸ�U��C����K�'T�*5.o�K��6�f%e^*/�Lt�O�aE�N�,��-���۶��|�2�cVn;'���_Q�O�Ӣ$\Wo]k]oU�̧�o�������wLVs^�c�і�_��;��n\O�����1R�z9ӧR%s4mY�p2,��L�;��\����:\]�#l틮o�O� ��G�}z���2%v����9(U��z$p%�Zj��Z�U�%-D��a_mՑll��m�M��{:V���en1(�IDs,[��K�����H�9�N{0k�kiu������-s��<�t:�_#���fGV1f����Z"���}�.����O�7�k{1�fp&�H���ɨ��/R�U���#��ꇤ���$"�p$`w �h���2C����u+M���7]Z�M��}MbT`�����0fX1��9�Ӟ�=�J8S5��e%E�}�hY{:5|_E�[r]�]5iq��5�Y2�퐴!&4�r!Ƞ�r%eHW$y�<٣,u/���ՙ|�T���93g�j]��ڲRV��<�`�h7���%���|�z*k�	6T�N'��#X7�a��ؽ�e����7ϳk5m5w]�-�KQ�p�����tD�KyQ�z�Wq�Ƌ��%|��{��r��S�|.v�+2]�D�]h�3��qP����3x�w��{4 ���?,z�qqg i�@a��l�Ĵ����1;��]�W�����c{u�\�7L��\���.�`l��geK��>˜��؜he[���5��o����ٻR<�i�H<Թ��!��[��&xp�/0T8[X�ڇyM^F�ە��ҍY�vts�p�1��_c�Ù��Ti�G-�^a���Npi�}��61�u ЧN+K]���t����1W����������:���'�O:)#tmQ���D7))֜,5�Le�U܂�Q�������>�N�ޠ�����5�y�v��=�Q7;�n�9�ka�ԁ��ʗ�<�2�����]��]�w�����;S8��RXnpi�p��4�k3t���hK�����T%C vZ2���՛N�z�� +��g��j^4��w�����8�����g�|||8���g��ϧ�M�r�.O#�I����΂aR�(����u�O__�8������?�������SÜdi$���v=u��|8Eo6:�**$��}q�����?��g����E�NX�s����qcr��*�c (����c�rܺ�&*�x��������?G_Y�\k|�|s
1��� �]�)���)$��آ���L���������q�������m�����gs���wWh��~x�����θ��"���3��������\q�~��o����B�����	R�B�@��H��I�9ƻ�Iwvr�H�w;�IQW97NLD|o�D!��v��!-'.c!Π$�_�O;�w]`��/��/�4!a�]%�����C!wnAQ�.�fƍ��ɾ�@#b�.^F��Aa�9j���iͷ��{-��+`���/�O���n^Z���ǿ��5��w�ye��2���6�f�~�tɴ��X=��O��S��צ�r�c�2}���$��+˾D���:i�϶�,�/�V�A�#!������H�_��G��8�A�/ihU9�<�3���pCu�Z�dlnv�$7g��*q�xmT��#�H� �o��Hw�ASύm�<�:�r�2���l'��y%u;�p-�-���jքʓ��wE�_5�94�~�� �l����H�#����t�y�P�	L�	���6U���2�D�z�8Z}ͧ��R�[;&,�w\۵=����g�9��b*�mŹ�aȎ��:+�SLQ4�Ό:�LH`Cw�k5z�`�X�q��r0�[>Z����VM>uȤ�����x�5��υ���z���g��c���e'�m�C:v���-�g���ȇ�@g��M�1�.A�:�4�Aʑ�!4W8��[ �So_,l�Mj;��?]]�k`f�4V��t��qC��K�$�T���0`�|ۭ��q�Z�"�$�w���nV��S��фI��ٶ��݌06݅7�c?��d[��u�5&�?W&g��ƚ�����Mg}���7����Z��f�W����:��+c�	�����kP��j��ya�j��JD��oia�����W�������M�Ӿ;���CX�!)W�[b�U�4&�9�U�{K��ժ��w3S��	I���p��\<H��#��1:yr���I<�/M�4sG��#�3�H�tv�ˮ$��H�4�t{�p�s�FBb�,�(^�;�����{L�rz���p���|T_@��3.�XCt��5��(�8�"0����]H��Ѣ]�;任�'	(�ő������떂8KV4T�_���' /\��\���h�^(D�V�[�\E�=6��P��'��hf�>ND0z��τ <>j�. *�/���R{�7I��x��4�@�m%��Tb�v���u@��c��	Ǉ����@Z�}����cl���Z��'�4 +����޽IW7e��`�k�o����@w��E�u�<LNv�P����i4�W�Y�@�����<'o���n�H��ȸ,"X-f��?{��[y�U�{���f}nS@��� �DY��v�O��[�/m؋���sһNv����n��x������ �8�Ԯqx��'/g���9�����'j����T�eW\v�"�븷`(�0�c" ����^��#�c��um7�k,��峜��ޢ�&�Dsp�_j�#"�y�,��3OQ]H;&U�%���6GB�BFm5Y�G�٤�C�]�[/.J
:����`�{�+��z��}����Mr*��:1=��m>�S��.��6C6e�e����wEJ��o l<;� iȷ��BDIi.# ��F0�`�B��!����/Ϡ�a��`��=���Ԯɵ��r�+�&M'�NRܿN{�^�pv���pBuF���!�.�f|ȼ�@n�o���v'�w�#����Dƞ�@\�[H�ܐ$�[xp��q
)53���!������9�R�ڹb�������	ٿt���Rr,���'�H2q݂9���ж/7g��V����n�!��y��ϸ�Es�dsJO��Y�N^V�M��(�m^�Fx��I%��&臮�=KI���=}�'}�̬�01iH���j��/҅�(#4�+��R&[�CH)���a��Ϯ$���n�	��0��<��B��Kw%l$O���8$U�f�|c�ᵩ3���9����ٚ��׶o�U�ld��e��<�Ϧ����L�
��s0fO:�v�b*�;r����g��q��cb���{�i���i��o~Y�|b[g5[�_K�H�I|�s�Л�l(��R����Yޏl�6�FĻ���ւ�;.p
`��h��������R�{���{��6��)a����(r��w(�m��1��*k�|�P�}�S��Up�}LPPd�Q�6�&��}�ܛ64�[�c���b�}�'
`�|�}�"�2�W���0���y��f����!��v�k|����Y�tZ��u�;��+Z�7&ٻW)�T=��P'��ۗ��&�o?t��:��P+qƕ���*�iˏt귚�g�\��<�ܘ^�
i��8�2���Mw:�2��ĭ��:�R��Y=��FtTZ}8/�� ��n�V����5��Y��7�t�]漵t\e7q�9drCO���_71ҨJ��#����}����c���عF2��ܧc�z���q��F���X�p �1�\1vffb�U8d!���<���0)ag^���ۻ�ֽ��c��k0G=_	[���u�A�ב�oB�b'�gQ���n91�oV��7278�F��q�g�c�7<���ѭ���;�=�1��5Wwy��l�p�O�%���v�e�1��yG]�*nr/M��e�i[�e�9����P4J��i���ɔ/F\�=��Y��a6����h�<�0�;<���P�k5����:s�����S��d��ץW���wj�Wӹ��ٻ�H�e�p�a6>�8m @�#�*��y�
\;�gن<�s���n΁b|E�m@�`I'��ɿ[�WR���]�5��~=���\���c��P/(w�nծ�=�`�z�q��t�=�-w�yPҼ��"dV�ڀ�G8�����/-��u��Ч`��^M!��q�=s�t�N�z�d����c7O\�O�^�c_�����}���*�H3֌������5CF
�[��3f=q�z_ѐn�t=�~���sr%8�����n$���.���< �}��͕/ל�^�/M}=^�(cw��\b�E��*�JW*Bۈ�,����\�����qy<�l�=�۪��P�+I����8�C�"��݉�#z<��]��������U<ol�R�&���i��p~O�<�U�X�Ood�uJ%�;��:n�xQn�v2�h/�J2��E���\������=��iw���ck8?e\�<��d���Lb�.�F��uI[����Ӎ*2�j9��KOT\��T�{w��n� �dA���I�g���t�ǀ����݂ܬ]��N�V�Js�.W��7��&�������R.����}�DA/���8A$T7}��^-�����v�b���I@�1T�b�@��oדuL���f��>���[d?4wm��|�R�lgk�<�U�2����d�J��Bm��<�M3�b0�%��)l�
��s�Y���x�R�Sj���S`ɏ>]f�oc�A%V��5j m���z|cˏk��|�&Z�4���l56uUر�k�~��|����/T�n2Ț�%��_�z� �,l�n)�:v��7����7�@��3��3`l<z�^=�s���1�t޲�CtIp�0��E����k��:�=�0>&j�ls��f{ʊX:�L���Κ� ���� ?UC��zs?��;�8֦���>��/���?����m�^����o~mE��i�ݰ�;Y�� ӯ7����y"��f�#�got��cӐ[l^�ɵ;�Z7{�;�RZ+5Fi���q�#.����������p
�{ ڟ��k�a��|�T���4h&��>�{�ن�rO�B.�}��wL����^;�ݻ�ró�W;r�VX\���������c�83i��*]'	!H�8���K��ȡaPG���(08x*�ӹ�ᷪ$�]����O/�:NO�~|���wg/�M������Q�M԰�v-�з�[���!�����єE+��]���몙[�]W�jSMj�[���-��TwNs{�Fk�N���O�uٙ�f�lU_��ʪ1iM�ȫ=��@���u��g�9n*���e�jŲ��>AC���o]⸖�g6��cx����Aϼ5�ت�" �<��s-0,��ח�6;����S�wM��,yRSh�
��l��f��T5%O�^W�\+m��(|>��ok\>��������������ĉ�㗚ε�l�i;9�ȡU�����eT��Y�l���̎����=E�Rw�"	vr��q^<��݀��>���e��N��GQ�Z��-�V��9� ɒ��U��4�+�	���5	۩�h��ڎx��&pns�ZHJS�!^ʷ����aM� Q�:�0�AR���xNP��v�$v�j^���&�C�MMw����αpKɔ-Nb�|-]���\�r_{�Quq�U\��|��O��L����V���x� H!N��i��}����$�֨DO� �s��Z�kz*��ّ��5��I�f��ZHon؊�Ŏ�"��`8�*����ʷL<��D���*��\�h����m��%���b��z[,�0n��4clvިי����8�������|���8�6f�7�����z/Y���3藀Ҁ�q�:bb\o5k�����ի�g��B�ɩ,o�K3�㾪("&<��jGtg�	�l��j���1�E�T�fy�j���!�$4���}��+�����|�j�eI$��T����7AV�i^>��{S���G�kg�.���6n�o�$��L6���|�{�Zm����U�	��}�I�]�%=꫎�5���2+r!�#;g)n>���0R}T��Z}�m���� ����=}]��v���֛��FU�%��g�6zW��L���.+��Gsv�<�H����ݓP�Xp�2վ[v�0�W�oG:t����9	�GX\�������R6�8��64������|���}%+����	�!��� x��j���.�w�t�b}�ѮܯWݬ~�`J���S�mA�v�ٶWK4:�''�׷�Hn�������':�[��u�l���matc=sY�3����Y��J�ZqAy蚠��s^1um�O��
!�?�ܷ�h��g�2�pq������O�"����d�}��f2�ta@��m�5�,ټ�����`D�;;�5���X[l�ۯ7y|;y��U�H
��7��oG�{ �^�ю/ۂ���/����o:���0LZ_�hW,��.���6|{p'F��]oC+����AS� _m�w�3/B�5R����>��>~�@wJ�ܱ���Ҷ�w�Ui����t��i�/FA�p��F$	��f�C���)�x���v�o;m>"h�����KO`J�̜ڸg#=����R��J\�#Bt�8�Rv8z���J��8+E��_����tm�*U �܊���:�oUZ|�y�;ߙף�hi�����HC�V=UPU�s_t���%ԝ�e>��͠�}��No���+{�̫Y}�vk�e��w�60��d~���yc�gw��J��rN$�-�U%���X���/��L��W�5�]��yֶy���Y
����u*��bg�}_�B����Dp�0� #�#7+o���C"�ĸ`�ݜ\9`z��f������Y=W�[��:m6�b�~zw���*kj��4םX�,��> �Leŭ>�~�e��B��Ǜ��y��q>Ktl�`��6p9c�lo3�ޘ=R&^*j�%+';թ�,i����Ʀ���nڑ��L��Mm/��Zby �{#o�s+�Ův*�����l�m�8�WS�<ꚲ��>�K>(M6��p&��n�7W�<��h���l�8�����Z+k<*q���O��r/b���Vl .j�����zz^Z�e�xRʽ{}���F����NΫ�pr^yD{2U�O���<i9���v���a~oT��7�e1}�el�]�o{98�v�ù�!¦�RV���L-�nm����4y6�bt���{�K,��u���z=��M�2S��k��z�����^�Im��xj�R6i�ӈj�oY�H�Znm+(�^��W0A�7f�v<��
�n6贬���ⴱ����.�,�ê����7��jOc혫-��ێ�`�v�Es8U���R���e�W����:�Fk���n��k2�Cs
^?F;��ʸ�ܢ��,���d��:��FϛB�ܺ}N,������R��]�$�0a�����^Nъ�=jT��|p.����*�iͺ�N��w^��-� �L ߞVL�T�J�K¬P�\q�j�pU��)󬉥A	�.y!�8!�1,#UoKY��Z�b(U\vZ`�����L�VW0z̖)�J�<a��BW n�y�D��E��<(u���G2z���Ty��f��*���o�����}�Up�:p��^���](ru<`�,
��`U�TH'�I,�߬��{�����o�J)֊���R5�������[��ep͛���#Č�W���N�PK���Y�97|֫H^@BI�#�m�eШ���L#/�)�Wb0io�df[��"�(��RDQ>��� �<2�/d�CV2��-�d٧k*�iV۩/�n��`,5��V� %�*���e4�6S�	�f�E��fz-V4�
��o�/%����&'1�k(�o#A�C+���r���xF6�@�B����(w�J�����sR���|yN[��k��Wg-�1t���O�e�'+�ak�Fؒ��7���"Gu�5�ɣ�u�]o5�
v_]¢]�4�WV��W{ӹw�W��n����8�B�株�h=�#RS�E�Σ 7�:�޻ڏ��_nN��0��1>�W|�[6�[�s������ʒ�LR:��n��6���p}ZE["���s+['Y(>�L���F��f	����q|cyE}�v9�AB�M�saqV�Ǔ�Y��7��D�\�\��c7r�!F�g]����joM�y��Eg^�l��<r�_o]J5�xj^%���|%sŽ�U�Z�M��Ce;��Z��L���N����js;NM� ���A����Φ\L�L�6JDK<�H-�o6�-{�:��..��љ���`��#����,N7֟u4zD<�a�z�;+VX-�|��K'iU�����Z����-���BkY��ټ�^�Zݵ����޳K$�y�Na�-��%.�gh{V.Ѻok��V�9NT j�R5�B
Rf5��Bh�Ӕ��BNRa��Q�Sc�(ڤ��=)�j��$
��bQV���hO� 7A�e4ɦP4���)H(��+P�Ah��d� ��N2(�B*�%S	�L��"q�P=��A��5	`�
�kv7,���u�!����@�q�MТ�ƪ�E�&�ba��T�I�H�ȧ���I�I ��6 	 1!BD�������u������������㎎��>>��D+��Q���1��λ��M�k��}{}||||~8�������:w�(����.��WM�ns1��'��8�����?����}���?]K` d$C)}o���~�YOj�H�)"1�=>������|}~����W=����,m�.J4��HI$���A����z��痑/9\�× ���ʾ����Ƿ����]}}f{wf*�M��}︨&����Br�S%9�G/Fz{}|{{{{{~?G��g���݆e�s�\���I�Ѳf��,�۫�9�5%�\��\����]'�u%�������r*Lb����z�F(Nk��G�ɤG�������'usE.v)��wq��L���!��on'w#Ji=~ywww}���E] �2��ܗz�����Hj����g�k�����tc��d�h娧ZO3�
��V�M��(8�.���ePE�@���Q+��d'���B	��r����C�mŹM��$Q�	P�!�I�?2�xw�\�k��0@uH����g�e�q�Ѵ�n��-�2�����9����kb�wT�dW���b7k�q���7Gh��n�<�U��1'��2���ŭ���2]3�.X�9�j�7N����V4�a*����kt���lnkEw�*\F�q������D�n�����=�-�:k�%��g�9O4s>�_V�e�hU��C<8��":�o���1$�A���|�6�k�x�=��݀j��N���\��n;�k ߯݈kا�݉ǡ�*�V�S=i�2f�����Oq��bH�|<g��8��= {� �Eωx��J�n�c4���H$�a�D���Ϙ{�guM�z��7=S�ϼ4U��;�X��R��;m�V�/��O7�cg���=��\3 ��b��C;)$��Y���j+ڳMXό�=�ېbג,0�|��4�e󬊹0(n�p�lk�!���ģ�==Ξ���#U"�6��KH�������D߸Ԗ�ɖ_�R��^�o(-�a;Y����P,�P��S���<Hďx��K3d���rz�q�'y/H=� N�����J��o�:��fy�`Z��ݎ\��1���W4�f���w�)Tk��O[TYV����ҽcIK�>��z<����׷h�4�ou���ԩf�E��^��)��uק���ă>�[�a��>V�F���//k{�
��]k��{��-���C����a���>t}�մ:�E0xz���*s�o����頺�fv�qޜ��Z��hG;�r`y�߯6�h�cb9�r(WUMo\N=����Ǳ�H$��r�7=0vr�d+��Fo���oKn�&H�|�����"z�Q�Yp[�9�Y��n{����=���!�(|�Kz=3��V�>��CCDL6g�g�-�]FV0�z���/���,�g�:=>�������l�6'M���vb@�n�Q�OPhs ���-��A9�������0�<��O��<>���05��S�$Jѫ�ن+*c��ҭ�`;U�������u�Y���8��@)Z���N��~�8<�!����s���w�9��F]�ߒ웓8��΂�������GlA�����P����=ޮUO�u��Ut�Y���qElj�V)��Fb�y۞lD���a}}wBbف��}�GoSw]/n��T�5ƭ��4�aM9�!	Q�������=>���\��b�Z)6���s�c'�z��H�����?x+��`�n<�s�~Ij�i�<�ҠkG������׬��G���z�M��p�1��|���p���e���Z�^|�W;��1{v�x�ݛ��R��wv����G���>9��G+�F��x|��3���)oM���ܕ��T	�ݺ�$@�[y����ɅkD��܊f����I2�(N�G�oy{&�5XQn�t�p� 5��'`�D�s����{�8��Z��t=p�oba\w{p@]���w}��;"*�b�X��ҩ�oo^�`MڤnRlY���~��x�{c�D8�R�K���\��;��%S,.D"gO�9����|J��q��kG�;���|��{Ƿ������g�J�鋘��;�Ǧ,��@��b<U6^js����K6�آ`� yv�Q����-�x%�;�>_(�K�BCc��c=����6z!qk���7�4'�D+��+�4��O�_���η��'��L�4<�s�ݰ7h�T����5��J���{k�
u�z��[�Q��A��8�$Ty*.f�����U�+�M�]��P�o�2=<���6�h�k/wLVDzx[fˌɀ2}�q
����4I�����vhǼ����Y�:��l����k<^�mQ�˺���E����Z�{[���{@�M�	r��][�4��o ՠG`vNT�m�M��5b�FY�=��6X���!��1�M>�=� \g_@�����Cs_n]��s`<R��P+�Q�y��b̲Ccy�2	��̯1���]���Ԩ�n�db	�ۙ@.��3�!r�����w��#=�zV��c�1�R9(bi^GeA�y]Ԩ�������r�������#~�淞 z�@�إWEJ���ڙ]��K�F���)�j[�t�<p�(�M:�<0^wu�U-m�m=njr'F�Z�I{�x4Ԗ��zX�H��j�C�m��&o�!Fe��2,#�2Jp��QD�2FL%����G?H�K�
9��^=�}�,�l�Bg����Ӹ��#�-{9#�����bE
b*�UIg�~���hȵ��>��4�{v�Ǉ��.���4�=Y��S�f.�ǝ'Mk��tE��y�
�:��<�_��_�˪N�T�������S�
A1�a�QD����y�#$E�qꝡZ�W[��oZ��,�BY��C���q[���<�W�)��U����������č�:fA�h�4;�^��'�>�ּ�Ȭ�k`y3��JC��^��S9w�!gZ�b�?�Ȟ��P��؁��G��)�Pʽ�#�Z����u.t�hm{z��p�I�^x�:��x��|XF�>��K��p5�[;u�jЪ� ��`>-�l��$�b�ff�<�����}�<D�m�R�l�I.�o7�C�Զ�q�z�D�Y��kl�@�q��{盅^�:�bՐ�����ڙ����bځ�d��Q%8�#weLD�M��jH���TC¶J�[��e�Y�;㙷��>�i��U�J\N7�*���!� ^��it�*^�-]��%]t���l!��:�ۆ�H
�nb-ۿ.�z�5/�0I��p< H���x�GWR��}��2�n��99�qr���0;��i���x�'���dSm浈94���I�����-U4zh�&	�W�n"�@�ks6�q\�+{)���������}�߷s�;Q�~�>?[�����?��[3�+[��5v+�دwH�۫���Ys�.#[ʚ�ܳ'��CX���_w1̳x�4+yF�_���r�E�������δ�0�[k:���a㫡�痟8�u���j�m�we��4�L�F��"�aG�I��a�Xc��V*�;<���{s���ǜdu�Df�s+�!��y�M�[�QNF��_��G�k`R��K�
�Ck��ݫX�ބ�z�E�f��f���-�s����Ĉ�T"��u�x����3�N���WJ�u���Dܖ�G�#�ϯs1�駣jɌぴ찿VSҴ�ͥ���'iԺzɺ�6Z4��Q�/�^ݵ-
�B�ǧ��g�6I�۷7*�v�E@�<� ����/�:�!�J��د�p/1�vt���C��3R˙_����^�$x�,<��j�r�m����G�|�$W]M.��C=���K�!���av�Ƨg�R�$���ډZ�ˢ�&�7n3��0-��.�^Wf��?!aV�q�w���f�U�����f��hqpY	iI��#Õ����N�د:�'aOt�b49s
wG�ɮ��*�/S]����eTc0�s-���#��n��y':�	�SA�o`n�)��2&���|{ 	jg��iz�Z�)���4���z���pSomT��{�S��9�RuF�ޫ=�!����GJS�7=޷#��5;�o�	)���>l+���h��Y�k-��l�~�6ٺ�4/<�Ks��ݙ���AI�b��+s���F�f �/��ܺpT�[�{����q[�Ț�}h�`������6�Z����O$Y��N71� ��+�?�����g���s/n��{������Я�A�iq���o��x�k�nS8�?W0 ����b&��C��A �5�����=�Vc������d�k+�h�]s&����;��g��Z왯�-Uf�	B�9W[{��I$y���k����ged1$�{��d
��#Ú�,D�9c�S��a�vOF^^�d]C��V���G���y�T�lWY�󟇚��U�Q���7\�ݑl���K�ÿZ;)(f�g�f!��CV'���o�]��r�EfǶ-�췶7�.���H<�6�=d�<=s�r	��+���ذ8�*�0�m>���cB�{3'`��hk�	x!��ac���X�ݢ�k�R�����B\���jL���[� =[�m�X	[y�O�`^�xuŧz�d�z/���#�:���B�A�r|���SY ���)�e��9I$����Cj�/�5Ѝ��d�%�;rZ��*���^*Z��fO��},�[�:vw���8�k�>�=�3@�ۘ����
�;
�o�a��fu�h�Cƍ�i��g�G�^�s��Z��@P�S��j�E��%z����;U�z���ҵD�v� ��4��{�wݨ�s�b�3ۣn��A�a\��]����ʻ#ʹh�8��F�4Q��X��
�l*U;��Ε�{Lͼ��gb!Sߞ�&M��s����^^�\�L��X�p=��e�j�U��!�b�-��L��b�(D�2#a!4&]!UVl9D���#�G8C���ğz��0r�u2�٥����ji�)�D}L�C��/��'t�/���g�A�bSC�H�w7 ����L+]�1�F�n�T�ިȩwpXʍ�<[Yh��٫`��;R�kU7lwT]{2�	��SR�V�����.�~��˰�f.x�o)J�;�%-m@���^���Fu��]5��ޤ��6ck.��aN�T��&Z���N�R��*�}1�~��ޟ6����X��H�}��ə�U������}ё���M�'���"���Yd?��}�5�ᙷ�i�6!꧹��QA��K�݀�I&����5���:�D�-P�TK�L�� 4Û�X�>y�_z�}���{Dt��q=uߡ�y)3x�Z��jw�`������=t���BD�l�)_(QoM2F�,r�X|�§'��Lm\=f͎�H[f�j��Ncّ���c�u����X�
�=��N-B��<t~��u#��6��ެ:�	��X�����듋1Z�Z������+e\'	p�:��H�Q[s�t�roW9WV��A-���ugj9kplSp��{�;2�Ups*�\
 )�F6\!���tnu���Iy��oL�����ha���R�{�\��-��D�ڭI�Nي��=S�ƞ3�M#�^|d�%�d洳MS=��fux7'�0��Dc�aXw�;�,o۶n�6���,�굟�ۺԳ[�V߲^%¥9ŷ�,�	�E��E�:G����LsV�FNfl쫲<�g8i����jsMl]	�pޞ2!D�tE7n^R��4��Ӝ�Z����������w���%����F���("�j$���=�}�#<��:��!.Q�W��Vt�s()��v9����='�5��G�f0����clh��2F��H~ �ý�T���f3���-��>>�οOS��Q���6���.o3%�7O�U�[��<-���Èa�u�}A�����\�}�ː�rTީ��g��y�uLhqa+>1��:��t�: 7aX҃k�T�x1%�\��Yխ�/|��wD]>f�.�Q���VEg�'՛��7�iB�"���Wp۰���R��c�]>���ܕ���f�;:�%�3.��"�RU���8՘Uc$w>f9��d��-�W�P.��Y�d�}�i�J�ɜ0Q܉@.G�ۙ�
���)�6�Չu�d]yƻ�nP��twNVT��+��qWH����\2U�ۮ�\��aZ��m���JGF�.wK�6y� ���e (ZN����Dg^�[�%|����jCO�xK5�n>����S��E�g3X*�Xy��36؍��3;����.��u����r�߅uҚI���T�ʬm��7���ޡX����rM;�f`ty�$-����S3�}yɍ�x��K8�'�r������u��,�Z3�ND,��Y�E�i-Ỡ�TJ{��ZgAڔ�;1
��S+����N���\`�G�Vj�;�\����\�tV:%�3U#��k�,qfe�p)b=k1�t���ϏԚ��n�NSr�`�45w�n���wo_!
�N���2 \��CL�R��)�v�nM�̓���B�cЉ��̂32�rً��݄��Q��̍ɠ�B�p�!�gד��2��o5Z�k/"7��U������h�۱�h�J\���;tsH�T4V�}.�:�K�С�v�&���f�4�j$��9`��r���Rwl������˔u��ٻl��uєV��#gQ�Vb���Ab�_��u��=ɬM����৶�M>�r��<��5�lΥo;*+��[w"�nml��נ������@h����d%��%m�;3����B�f�Q��9�Q+w�1���@�ٷ}�WJv���O�ݼ�!z�uG4�B�9���n�Z��qڬ�� �����\ٌ{��pS��9�ꉛ���)�I� {�������E3�o`Wյ���V�8�1�&�Imj%�O6��̰�l�WV9��1��}[ь��o)��4.�Wm�|F�R����Xr��Op�4+�pE���ǈ �d5�,�kn�p{�v����Tnp\T������2�������D��������5\2b��+Sɝd�����i�R|�Ο=zY8��M���ǯ������M����	�i�v�V�)���a`�g,����y�=Ŵljbf����9�g�˃i詾Qu�|7c)���q�C�^��;��ǒ�=��o�,)n53^�N
������uOH��sˢw�EeE�&����t��q:[L(e<g���$o��un��t�w#Nf>�ح)�l;�P�"E�I� �A\������W�]��ƪ
J���#�������������]}f{~�o9E���b�p�F�+�B��cx�6��x�G���;;��lݽo[���������>��=�:�Q�
�&r�[�/׈�Jb$�f������{ޞ����}}_Y���ݪ$���M	%��ʸW8c�M%;��L}�n�o��������~>����n�1QMD�T�!A�.}t�o�\�[�O����37o��x������~>���=��U��<��;���q��{[��>�q������fx���|{{{{~��:���� �x)c!E>89�Y�t}\e箫�I�n	k=;�*��&�;x���y�K�WA��&dDX4Q�`��ۉAd+�w��A�oM�}�e��G���E�E���L�]�P��ǝ���K�N�d��]P�mw#n>�t�V��ҏ^q�h�ސ��Ai�Ä8H���]�����R�_`��$K`ҨT_�:��$1�OKn��<��/��nh��諮�e=n��Mo�ٖ3H]ms��-���f�Ь�ޙ׿'�sw���I�yP�׌yW���~��9�{z�t]�d�n��n�V],�@9VI��}�1c����3�J��w8��s'o+����9!ڙ�8w~\l�f(��}��U�<�F�ޣL��niTؕ�s��mX�\�582����>on˯3���y��)�9�D>UL�1s�/�jIqJO`��3ۀz�6;�G�+�z3��'-���`�JS�{m��.3U3biKS� T�Y�m�S����<r�{
�������L����Iu=��,�;Tq���f�����5S���frk3��}؉�gS;�n:|S��L����f}wM���vK6^C�QC�ou9]��9Z�S�";o[�uL�3,�+���L[^����kͫ6�g�%����a��X �e����q�٣mfꝓ�E�� �eV��h.1Ԃ�zD�Ϙ/��,��;[�*����F^
˺�_�?H��eב���P��-�� f���S�X����|�t��SL�OH�̓v�\�[W?������bp%��݀o,]!�=��j�j��8��"	�D#���K���>�� ��D�t��[���p^�;M�,'�_�����M��y���Yw��rm%��d����5`��l2��OFҴDQ3��r�^%�o#�}������b��8�y�ߛa���=#C�mS���:[�w�� �_���U�T�ћp�!�K���ǵ�:r:Ħ=�P����ۛB��ҟ>�ˍ9��EY�7gD�d'R�	�%P<�دEk���]���vΏc��;�elk��
R����ǯ���4��*���0��47�:k��(tP��6�X�������j����,��jц�ډ�z���@���Ub��v����	�Wy��N�^�]&���#��0 ��I���Al� İ��z�~�؂_*�L��h�o	�u�PMC4{�>c+��#A�F�� (S `������D�@��Z���\Χ������z�q��N�O��d��6VQO&����Zs�̝���quM�hʝ� �w�P��-���,_�2	9-'#��!�9E�����m�d?8m ��f�	חgm���s�6�J����U�%F�E��j�жM�,�O�:���	�2=��y��JN�F�7����F慚Z�-4��c���5���Q�3{&nM2�I����|�����C� ��y�����,��s��	V��p����"en7���z�Yu�޸s �ě��q���L���RMd9�hɝ�n�׍Uެ�t�=�r*��u\V��HT��l����~�܊��]��=땽9��	�^9���6�ͳ�;h��N�r����M~�+]�j��o���;}�!wY�Ϟl[b=r۱-�� d�M���O�$]�pY����=��#�}>���TOo�,�f�m��}��e��N�7�^���o���[1�'����9S�n�v}�tWEݼ��p�Z�5�E޾@�[l����U���k����ZeFy��j�9�y;�u��$�-=� ٗn��流��&9]��n�vG8c���Y���̸sWVK��fL��=�¯7�%�	 �8�v�o}� ��7�w��(Ts�����RZ�����te_6���Gz�p����u������:�� �<	���݆w?le�K��>�k|A]�"*���ڠm���-�����I'/[áS=�E_%�ս^�`�7O(����0,�9�}��rki"���y8L��	���VǅA���Џ?RU�C/��u�-�Ֆ��ӱv�6��e!���3nթ�z*�ԙ�n�����M��ꢯ�����gg˂͔�G��L��_c��G~��������%�i��� ��{�� ӵj�F�n���>���̔�%�u��F�zTVq^tb�g
���u�(P����ϻ�I�0vY���L�M6*;��߭JʖRS:g��3&������#"-�b�d��v��hi��g���u]��YI^���ͫ�*���=?
����X����Z��՜����E�ӪP��ȳy�Ʊ��Ƒ�Q�x!d^�-z�q�����{�G8��Q�R���\���8�Hn�V����Ե�;O�����G�#ď<G᪺~��b;C��kߓ���S듩�[νe��K[Q��\C��+	>�%��������k66/�˷w˺��#S6�h�J9Z�=��3'"������9N7�^Ow����0����rn�_S{�`���k�ڍ��������>9�с����}٢��' m�!d�B<%p�{}}]������ؐ�a������a���I����OM]��U��`O�S��Fc���4�]ٳ}��[;c��_=l��Q���6����{܁���e.�:D]�W"�f��:��V��Ė.Ig���}yb�Fn��_;\�	�8XL��T��W����l�i��ͯ����늧�����Wᢴ�>�n��U�ͩ����	q���7@�82�<띞w����;*��+gz�xƝ����hX�-V��Ruq��c��Ñ,�%`�}��g�c<R��}���ȍ>���<��م{E溏>��f��6m�s�`٤�I��i�&�j��u.��y� ���f��{�kyn��0��A�Hf��	eF���� �䛙�SY��
�'w0��wH-SN3�4�����I��^��~��T�,Fod�M�m�~-���r�ݳ^B��j�q&vvw""1`D�����/\3{�d�]y��,�;\�z�(�#�4��N�i��0.��g0Z��#�a6B���[���]s���j�D��n̉��@:�O(�a冬��)�۳��/� є��Z����n�S�a`ey���oc�7'7����gn�y��i�T�fR���O�IJ����T53��dx�q��K]eY��7}���o�w�+�Hu���]wP-V��e�8ϿgOa��������Z���;�{�N�g�T��@��g~��;^��2���V�(׶l�'n�={��ӑ[����v��y�Z���4i����-���5�;ӱU����0�4wg2����*'\�T[5v��j�3�����!V!��Y�$J2�Ej��.I��hB ��pH�e���[�3����Hgx�v��tko�¤+0k`�˝LC[�u�S���Ȃ�Q�o{P���"�#Ŷhl6	�L6�!2F˄���8D���<O��y�F�""V��lar�/����&!m{]*�\u�c��{�W��ʋ���(��;.Z���u���C�Y�@yDumzRy�kT����������o�qN��T�)�y�dM���#�ݺ���I�<���|���6��B�Q�t���`�\B�����}�������ȇ��k�����Z.�U�j���,�u�8`}�����ۧx�E �H2{3уTc\��̃*��d��v�<G�Ǧv�����+U�H�������ѭ�[���j�̌� j ��w���c�{�<�q�gl݅�p�§w����[�MV��7b��q�1&}��E���Y�nPΖ�����\��̽�,�QE��� �y���U�����Լ;����k/�F9ds��^w�/�x���OӘع�Ȥ�dNʁ*��T�w�����һi����CB��}�#Kv�_&����6{��We�{�,��i����v�G6�F�Һ�\��wb:�`G�<�*@9���{��GpnMo�a���6r`������vۗ:]>�sx�u,�􂻐����շa��:ck7��x>$x�e���=Y��K7Un'�����Ӯ�T���t�[��8n�;nm9�$Z:���w�������@Kj��(+0��#���d�i6VǱ�ǥs���z�v{g3x�?���f�ʨqB�/��q�ko�l�Y�5O%��[��s�4uɷ�$�t�VƩͺ��XM���X�@΁[��l��#�V3�b���qT�4rC�_۹�'�c|��� �e����������S�t�r��t�I$b �czP*�(uQ��/���[�Cc�᮳��D$Z��L�{�>y���Q/�x�+�FoT�%���fJ���?�FVIΫ�I�m���dB�L���[��>p�9>l����gr"TM�n.�������xS����_���P�z�+�Z��B��er�񙚑�v -1��1	�c�'Wo�F��"t⽣M������,B;c�D�C����39t�FN|)�<�������0�Z�ǔ���x^bS������X�LHt=a�����;�<�N{���`�aV��ڕT��~(��<=�ss���;1�zϩ�w�j>B�z�f�7&dg`��j���ӵS}t�^*�9��z��	R��3�u����LB�>��'ޓ��B�e
��*1�@L���ӻ��[ܥOGuV�}����7ri�O�^#<�����=XՌ��Bц5�٘:�e<�a���MvةvN�7o���j7U[_Q4ϒ$�z����KvpJ~�H��lpr���.�問܂�̉L暫��c]��O/��XQc�@�g6O7�SOiia�����]Y�"%GL>���mT�P�o@�07�A�3��$�nU� W?;e��=P]����۴WT�!^��ja�7�u�;X?�7(�ͫ�̎��C�`�I p5��m��[��uUo�ۘq�C��\���<߻�O�܁u�ZC�-���2e�xl��K��[rl���I׈>G���ݳM,4 �����D(k�lh�,����s���R��Ou[���O
��9�h�rЗ�_��ƙy4b5mw����9�ס/��#��� ��rb�g�z�z~{'�Μ���S��ù#4��
:�v_@�I���w��RW���Xgr�3�8��V>e8!��\�fw��u�l��$"��!��.�x�^xo.B��T��pP��§p��ֻX�-*\�\��9�-Ng0�ف"=�`5R��zd��
_I��X�Z
��������;:3XL#/�^�܂�M�#+��6�n	$=���?��@�DTj�lr�ޘyu+��y��C��ѹ�[1w�keA�*]Tء�Υ{Q�놲%�3�5�S�ʼ�
_),-�[P�#�
����ˆ�`�ج��N���d����OR"r��v͵�,�pL� �w<�<HmY�1�\��oM��@�H���L�4j�Y���F�R�<tT쑊?�~����8�ǟ/�N�*��4�7ۅ=�X�r�Cs��7Ͱ�ҥ��X��\q�;�7�1�;�\λ�X]t��g":���à��l��JY��V6�Ɨ���9���K;�7A�3u�	������Qq��������9��ݡM�
��T�2{Tv]kP���sb�����y���ֵt"
, �.��Ut/U�p�S|&�.S��y�ι�*�\�dA�3�jG$��J�;�.��,�Sv�u�2F�+8TƤ����<j�f��%+[.)�&Ræ�фQ�ӿ%*�iV� ��Oi�	�6{]�O����q���)l�y@�^��
<ٚ`�ť����r ���>=��1]1���f%[NLc����\�k�޸x�+^�j������=���Ld�չ�1�$�p�b�f����Q�1�vD�e��YW�&��n��'<��W��5n_���2�6���O����ֵ;qL��"��]t�(��ԗ�������n��^���m�)��x�}v����i���ּ��bʝ�+-�V���y��mx��RO�s+�	/�1��ˮ�/Xa�b��Ӵ�s����hK����9��;��K��ޠF�[�n �=k`��M.�˺G��	�B�j/V��J�S'l�^3�1`Ҫ��N�:4���5M2�h0��D�Bk���X�;�b��'�J"`�XL�Q�DIJ�*�7E���`��I��Ze��Q%qS�K���I5kf�w3�C�=�B�ML��(�35B�I��D�4� ��]!D��L"�A&]J�X2*qY�pY��X����<E���(�T+��ʗ�Xw2MF��h_(�}r���M�ᮄVٻ�����Qwh 7����˫-ڷ����"���X��sv5��Ws��Qk�L�vfg:4�>���I]:.�!]��M��t0dk�Mz	�؟^�u��6��g���S�2���
�<آ[�m���-\U:R��Wb�`t��Q�	U�dUś;�L��V�����m=�fZSx��H�>�+��sWVX�w8_[�L�����00�u�.�+T�
��Vȸ ��#=�9��g�'jf�L���W(f��C��H�V�Y͔Ū&3�"�S��n��;�ւ�SLgr��/���u�t9{G�tx���N�X��U��WOqpu��[�nqf�7{/�9soj]d��;r���:���E���b�"R���Sch���1 
G_yS�*�tp}�Q���E�^�㭧��c$��4=������w�#�3/H(��J	�:?�p����g��\�Ǻ�3kg*ɧ����l;���I�n�m��u�wfX�N����������5	�#��u���h��X�:�W)Yc�PR�H�<2��9Nb��	m�:XZ�ؠ�
Ld�4�P1����Q�Z�ǃ�L��m��*EF�!TQ��IB%d4_a��*$��P2���-��M%��Ph&�\�5|E>j��"Tp�"J��!Q,�K��h�\+��	ea�Ӈ�Ht (�[q�IˊQ*�,��h"�
:d�)IR�Ơ~F�I�E�I�M��)! �@��s�`��Խs�����S�q�]x*1a�r�яZg�N>�=��������e���"���k�("3�Z�%F�Gy���o����oOoo��������w��p�GQ���sF�+���F��^��<�T���������Ƿ�������3Ӯ�Q5DDU���������C2�nE�D�z��OOo��oooo��:�����$cz��~��q�JX�..�w��F�k��$ӻ��K���<|}||{{{{}}~���=oϗ�h�bfǭ�p1����}�<�^����x�������������}}fzt6���o�r�o-~=~:��^��gy炒(�����b���zTWixۛ{[���痞z�zs�~i�xݞ�������^ڼY.��~y�dW�t���L����2P'5�%!�m�Ψ���-��~<�����VBt�S�Dl��fC�yu��u%h�I3�'s��2i,�t+v�!iWV �U�Y��L�8��˨:�9A²!�s�ͥ5��9RT�J�,�n&�`����$�"�PH!J��`��8A��Č��1v�V����3�ߝ Nt��\�kY������A���W��t7x�INOn���Ⱦm�oo^��p"o��ዹ��������H-{j��oS���ts���@e~͚��{C(�Fb-�ov�!�S���ުJ�[����ٓ{��A�������g��U:����)�p��G�_9K���{�U%��6�[��s"_s�D�N5îr��nl��;	OWU�K�əU��m?)��1�M=��{A�:$�����]��L̦F2|n�n�T^y&�&[�����g�]܊����>u �<��L�����:�YM�bس
j�L�|�~��s�n�P�N�-n��yZhRy�����w���&`mT�g���h�f� �`;E�z9X��{�C�U��^I���`'�5q�ҹ�N"�k��>M�j_j�w��L�,;�}/;�]�N��G�i� �)c��p�;�xwNV�M��W��%�̾|���f�Gϱ�`1ػ�<H� x�<DD޳��B���7qT���Q�o��n�R����k=(�ri�t��a9~Ial�9���Is�~:�=\����ѹT����\���7FC���x%w2�z��}���� �7�E<��'���jV�#\t��P�Y{s�k���Ҟ��ڢI�vٻ����=w�گϳ�S5�����ި�s��݉��j�5�y.~�W{Vd�iH� IR�K���Ȯ�M�}ї9Gv�.;*}��;���9[��<ӟ�E�,�mm�{��P)�d�C��w�����,6�u��}�6Gv�|wٛ�khl��dV�e��T��	�uxi�U��wl�.y>����ez�9�����v���j<����;�����e)���~	0���1Ձ��Άj��>���A.��g���J�co�&�%�Gk�.w�lv�|���Y��{�2��s���̠��d ��<���Rh�i+[�5/wy]����@�9H� ζ�+�v����ܴ��K�iLJ���D�
|��mC�8��v�h�CSwz,���'���_Y$x�=z�)�X��?{�s����)���;9�6tV��9�nZ�VEs�[+Fe�/���y(�S+���Kf������o�Mc�_-^��b��f�M7�26��]�7 ?�'����bP��	��Ιӳ�Q�^)�γx�x���eɞvj�If%��H�9����3bg�٘ֵp3t405d�r!��`_�}�d����~���;�5�b"0ww��m<�/�5�}�9�H6����{�.L���}e
(!w��ؗ�#�68�K+s6�t'��ġ\�	���0�JR���S*��P�pc�^毚5鰕&"j��J�f����Ϗ�}�OWT���S��T�B�k�Y��5��El)��6V�ނTn]	�[�~`�d�s�_B�py���2y�#��Y�y����u=�l"9ʲE�֝��{i��ד��m��#��8WQe^dU`c�R����cJa�ʧM1'��ϰLEoT����U?�iۯibK�WOo&^�|;,V��q	���1K�=�øK�z����UX5բp�t`�G?��$xօ��P���J�
J�̀I�[4�Q�!�`y��9���l�L���on�y��l���}�z�5�ߔ΂�-hR�H~�۝4	��g����1�n}����H&A���e��}��π�ܦ�w{�|'4e��pu��F}Qm������D�� Z����!L��7ז�#��.ߣ���&���(]�0��^��p�N:����d?.����*~_���%�x����G��	҇gv>f��㎻���G�b�,�Q��%].�u�'�x7��V9�o5@X�O�]�;l���_S�۷���j�昛2!m�l̝��]!��$E��d��u�zl��,3�����R�p�뼾=֤i]ޡ��,��	�2RV��"�;=/��目��7�[j������5���_݉��F�U3K�롦ʿQn%��w�ψ��*̷MI��"�i7�V�co�ۖx��Y�nY��Xy�%���TC�P]��i��P���۠�F��mMnL�eN���y��(�*��bƬ�w�1���B9�֥C��Z,��:��(!m
��i��&z��D�B��(�CD��5B�j���_ 8H��\��ɵ�tyN���]���O�~n�J�ٚ�O�(n8�U��ݲ�0[|��Y����̬�u��ix��|ە��������#k�ލ���/�g;v��w��~��ٛ��[�"x�q����G+�f��{J���V��2�=�S�4P��^P�m��XR�:7�8���d'ǻ\^+����9)=߷wT�Wһr���^g��i��[�[�������Z�1#�[����V��?b�y�{y_!�>�]j�#�+IcM�r6�$<�f�ћ[�V�ע���5	 g\�v�n��/���9�sLrg���V,>��5�4��z���gH	�n��֘���S��fD4��Y�K4��B}����(����5��z��$)��zB�����uq��/%F���51�\��a��]~������~��D���ȹ����b���N}o�sj`$���B�t�ݹ��4�eђ��  9��Gƾ����������p��;�����}���\ȆMUӦ�����֡Ҡ�p��۷kq�c�9�p��@�a02���u7�-?�i��6�zt��%W�R�d�7O{�k/X\�����!+��>�}:)%ᬬ��t�]���ׇ�")ne1V���YP#a3��z��d���X����w=�����s��wl�E�*�j����<��]��1 L�W��j�[�j��-�&8��l>q])]�B\����H>﫪�}�^���$�b�c�J��h���T3<nރ��R���r�o�2�xk<v�e�?�/��lm3���k�۸���{�&^iѹ�7�t�1ʏ4{�_����rɔ�����^ۋ��WW޵��~z��w���^魹��f>��]���4לVP�˭1oս���&PH4w�ً����<���';�N����O�n[	��"e����3�PU�. �::C���(��n��3{��ِ�Vf;�a�^��U�}F����d6��c�+�.E9�6�?y�ӯ!��}jo>پ޿D��l o)��n�U�t����K[[�k5������P�N�u�1%{�sM�*��0.�;Y��n�?��S<���u�Ӭn�GO�>�n��j��y���Ot���=�|*�Ͷ3��Mb�i?��}"����}G>�o�m�}�7���YY�i���)�"_۽=��f.��� �]{��]�Y�w�j,�f�Whۋ,���l��nw�bQ��L2�G�'��j��s�#����ݛ��H������c��Z�-u��կx��(�9�-�lA���{�Rl���7L'�.�c�[ܟS�@�j��7f�OsZ���L?gL���^���0�3�lfz���'��`�&�����h�	ۯ"�df�j��e��lc"�2�gDUmU6�	�V̙�Z�q�궫[.��7��k�ܶ�뚶m���*U%��UBkc=�p�<�+�Μ����$Pkzm�Im�K2�CK?#��;[xTTz{�Jx{�C�uYD�v���EW��/.���$��O���&�G0{�f�X��:�'��<��� 㧺W��ރ	ح���Vŭ:\풻Xˋ��i+�u�(��W[�^i۬ٗW�L�5�{@�����gT�X����z)���3~L�U_�UJ�<
�faF��s���[�[�r\iFoV���i��G����^��GE�U��oQ�c��8ެ�Ч�ޡl�X%m�BA.K88{Gzr�@M81����'Ύ�mWoWz��VL<a�������c�����Rg����nnjw�eK��Su(%�P;�Ժ,;.W�Π��]���;�j+݄ƞH5��K���f��*4��MƷ��5Ӑ+�qv��+��e�5���\�k@�<���8Q{�_of����$W�˗F�.̸~�x��;�z {؋]��kކy!>�_�U%�B;�V�.��Į1�3�|WGYbi�<��s{ʛϓ�b_�a�7�ݙ�o��ˇ�=�����a�R �Q��uA�����98ּ!��u2�Way���]���+�Q�R��f��s9�ҺLm��mI؁I��8��j���7�(mѡ���h�TEJ,M:A�F��PY�����oX�,���Y�;C�)���]�����8.�*��`��{ЗU�#sh �`ѶH�c��d$��!0���#	�e$�@�$�L5�c��� dp�8@�ulA��Y�#�dd`!�x��O�sP3��\v��f��W��*0UG��x�vwT�Z���V
���`xƬ�\ȏ>����C��7.f*�����H��Ւ��P&�����$l��;�9��^��ϊ�Y�ˈ��Y5��)l�Z�˦��5���Y�jq���&��f�(4��ӊZZN���j��פ�QV�-�~�n�2E%�^�v��׾�=K��f�6�m�w��$�1N�p."����p���j>.�K=~+2�H�ް�ќ��*�T^�4}ὓ���u0n����y��j��g����>ίm����TɃ���x�^Aoi۝�]�a!��y�n�$ؚ�t|)�H	�fET�����ՙ�}��{���'��� ���UU����!)O�Κ�1�X�9���L�'Ř*#��j���Ӭ�R��V9{��L�E�*{�;�v%��#�e�e猝��<����Þ�%�fg�J�t	^u��87�Ҫ�\��N��B&du6�kp��Տ:��]���������� �p��􆽱k�������m�kѱ\��7#��U<�U�}�ڪ{*�)�ţ�{����Y�����j���ڈ���MgB�@�����>k���BA��LE��-������{�^��;e�{�{9�
�]�fF��!F�{"�7k	�+�B��(����}����潈2�:꺙c�6�E�^���)����H�unpfS��n�1ws�v�x�K{�w=c}'�y�~�.�<~�B����%��$�}��T�d�a��t"��z�\̖��H�����`���)���{�����`uy��X�z)'U3�ə�f�Gy	����&!q޽��x��lڶՆ]�.�8ƶ��ǔؠ��D0��V�����g1Y<�d�ڄ6^�u�]��e��B��b��ׯr���=���Pq�lrv��b�m�c�[�**ً8����I��P��ۧ=a��ۊ���@��'���v9\,�d�[��I%Ӫ^F�i��)ۙ�Q]��f��WoTW��Lp#r��6�ҏ<�X�������o���u�c�pԱ��r����4�q _r�ڦ��[n��k
ۙ�e�7�S��l�ۼMJlQ�`���2�%��-�\�:�(��1aM=L��T�
l+3���*+�ّͫ�ۙ8�Ͷ����ľ��%�sU]Zږz>9��N�r����y�.W݊b��N�L�ӣ���v
U��v�&�0t�Ҩq�7v[�x��ҖV6�]a�ԎK��q��Ǔ-�����0�P�����c�d��X���4����]����H��*���\��+�5%2����T�Z�nfd�{ �9��Ke�z�oK�;��x�:_�T֪v�)�hp���M�i��__RSU�;�`��3�aY�2wiCr���nhf������0��ÜjRTnz�v�AvM]��.�R��K���2����Gx�'rcq�P�v�Nkse�j�t.}#��8��`�NU���w���|�Bnԗn�G:ñq��-��uX����Ap�+b���ɗ�o��Q�{$�x�5̂����e��X�b|�Hm�]9�YM�80�F���'z�'j���\%��A
4O�a
�EU*5�S�3`���W������Y�i!n`6���6(Y��P�<��$)#�NB��q�9��\�����RF5�n;���G�d��#)ۍ,�3k+)Tf��t�����E%\�
���������H_AgV2��N�T\��]=c���ii�%D�7dͭ�I��Y���zC��ݬ��*O���D�Qǝ��mr@��gN9�l��*يYsyV�&��5�x.¦V[szaueepi��Nu}z��@��+�wz�vz����ȹ�Zl��oh�.R���5:[�LK�U��ej�kU
�1����WR��,+�x�,0F�늽IV�ܣaR���΢���8�/�3eGw��
��P�۵%��B�GY�'�d8i���X����4^�5�N�W��X��S�2�uي��A-�W����P��y�<�ɣ���ݦ� �X�*
�a��4�K,�{u�٘iT
k:mb��W2ى��s����j-"��nW���=��ͱ]��K��^u�=�4ɝn�X�ΚrsC*����p �A���Wm\s�فZy���u-y���~`,����\���QVKjF��M��#��� "�$xA�s~6�o_�ժS�7;�y�IxۉDFO�ݻz�����������xΏ�n������k����+���܋&�<'���<x�����������x��}{tt��ƀ��4�}�>\�s��F�\��c�I��x�����������u��Ӯ�,6�㿍�*���t�6�W'.�F�\�ݝ��� �Y�ǧ���Ƿ����x�>�:)F�p���9���Cwƹ�W75�)o��7n�o����{{{}~3�������NG�rF�����^��뺘�<p�
�]0z���\|||{{}~��^�vR��(h�g���TckӘ-EPl�x�lQ�b��s��e�]���\�ս��0�ם]Er��9��sn����=ur,X�Q�_t�F�kD���\��W6AP��喲Z��S�*=�w�7km'���3�K�:�6	�1K��[:�;˗6��θ7���)���dpG�,��r@���U�s��B��]�^h��@FI�����B�v={[���Q��S�o\dr���F����cZ��mGSS�\����|�d�ț'#��B�z�]�@o�:�䨜l�E��+.���v^����l0�R�`�� �7L��c+���;2��BxŎ�F毓9>,�TЃv����nkp�;Tw/m-P6:��1��ު��Q�����n�ۛ�O��4�3g�ዷb�y_��j��;=ܻf�u�	�{w6��ٛ��~��q�X3X�����v\#�`��]ױ��.�N�`B��]dL	I�X�N�U��n`�5�.��G�.+��n2�90��)���/UZ��V66@���`���Mfb��a������`n�@�{�k�ps\�����"i�d�c�5�ȶj�p)NaW��{�8��퐭fQ�R��^>����%=�5��u�y�K�U���1ɋ�͘{��!����ุ�C�����
��}5��x�67�p�p< @�9U���e(� �����o�2��A �Q������K�y<[����Bt4�ޭg2q��'k.��5�p�~\�Jl=n<%S1��f�S��5�H%�Ph�[(~����i�U�`G6��rK�.fGY߄;�b�qcv�n�=�<�=�|��bV����2��kNZٜ�<��sZ�]�w����W6jճ��kӮ�=�նy�n�OQ����;���Ȯ���O��'��-������ޛ~��K0Yz�Y;O<ט���g��8�uHeO+�'dtr�fz��cz[�j�Tn0J�TXw�}X<-���5��`��ڤ���ј�r�}�5�䨣I��m�x������yOc�m�m;S���;f8|>�.UZ;�3���������ޠ�2�@�$����.5�q84}��%�A�}_�1b���S�3i_¦áW����9R�+m�I&�� f������[��a��g�� ��i��<V�I)cP��!��
Ap�ӧDF����[�2^=�gi��Nw�r�=�.�Z�qz�Ō��U���B�G [�m�Ͷ�R��i�P�η8���9@�3 �(TA�!E6��`�-�cP��х���i��4�w�o�o}��wfw,�#M�z;��i�b܏J] m�T�V��h�����d>=A͜���J������v/�����0�����p8uGJ�S��e�֣�O�d��í���c�6Ю[��˭�,YT˳�NW�C9���V��3�@l�i�J*��]�İf0o��&���q�Շ|Du��;�5����;tg�ǯk:$����B{%�Jm�PkԛW[O{@W�됡�k����V�2�� ��ل����!�{���~��+�"Y��k�d�)�`-�h`�-���m0����;#^kgΞk ?C����j�g�58ڣ�����ܛ킬AX�����Z�gĆ�b	���2�>�O+׾���]�j�٭�Z\��Nז����́M�%�X�84˖�'=,�Q��ā� �y�&w��<ĸ���L��~�9ZwSĢ�i�����5o����Z�oQԐ��m��(�X��|����w�AU�_�Y�y�.�y����rK��t�bŵ8�u��8��N�G���nj�-.�l��
P�ѣT$|9� �����S��~�S�1���/飽z.�j<�:磜4K��3�nfwD-��)螫��T<Ѫ����6��|����a���2}�9{��ը� _v������p�NK�g�#g���MY�����Y�҈������t
�9׷�v�۽]G�g�CV��(�Љ�[�bgF_x�ʼ���W0���ۓ�)�_b��pt��%�$�+� ���,�*�}�Nuz{/eb�!���zܧ/la�f%^Bm��M�	2�ai ~��>����n]�0�צ3��pو	��0Cl��DSU�t�3Ssɺb�>�>���_�E�}~7��q+V���z�o��R̅����I'>G���������L��fCz0����Ir�\�=��#9�۷�_Yۖ�4��c��ZM�hr����Mu��=8B��J����'l^������|[3S����~�}�E��|����n���\$��j �@�c����z�\[����f}o�5+��5�p͎QEN�w{��&�^�.I���*!��=dy<H-4V�fڭ-�8Zr�W/MQ�h�`r�3Ʒ��ۥ�<6Vs���Y���Z��IG�����U�C�,��&x8mm������,�Yj�ћE�b��:�l��g�71������U�K��M����W	�r��~ݫ�+
�>$,��8tL��s��˪	����&�=�ǆať3��ab�T%�U����������3Z��vU6.̦�5<��8�I�#8�l�쾞�Z¹\W@�j��\����DW�_fn.Ouj�����R������u`%�;6�\3��lhw��}H3U��'<O�G
wC6<�������v�M��\'���M�V�[�ܻ���y�R��qP_٦�?Zqb͟0>�q�>�n.�Xl����r�|㟾3�������hk�$/ϋ���k_
	��#l�۱�������o��f�c��|}6�s�J���^����L�}� R�H�x޲(��O��<7T�E������Bw��M3"�L�GN�Ƅ{��v}|ΥS�˂U&_vq���u
T�t���0��� @�#Ӆ��"!�^��i%�8'g��И6)����/�s�o���T�[6��JoQ"{��4�K�r�N�	e�U7Ɇ7���D2�!��=���=o����i��H��E�D�r�U=�(m��V��Z6#ϛ#��ֹm�~�ͫ��B3�ʔ8\�+_�m5�m�tNolw��zP�g&�L�r}��F���5����P���~�*�H��c.a-q�����E�FE������3�8�NϙwC��4���{���ݝ�xn�h��V�9�%�9�;tz����`�VB����:�k�͉|��Yj���`o�P9�]V�W�wy��Y]���0.��}���ı�$	�V��R��c��="`ɝ�7Ε�˻\A�s��K����mȁ��-����Ov�J����d�A�i�˞����ːt[~�w;L��Ʈn���-�ƵꥧG=��yL�ur?R�+d���	�D#�5�� C��7���m�3kUO�Z��K��;�I[m@[�����`�]8�p���`�����N��HA��-! h2�ER�DI�Ja@����q�8A�\t�⃳w�7��JO�".�u���VT�;���K�a�Rx�Po�͙���~R����r�v��w��zT ���:��=�>��}�8+�C��z9�%+k�f^�_w+�g�ػir��`�'ύch;S���d4Ҟ���s+ڳ�f�0����a_t��z�,T{W����Ă�����J"��;��o%"k$Y���ˠe�}IY�[໛����3!W�kc��Y�͙��������gd�-�wq��v���<�w��+����z>N�Ʒ��?���w�<���v/i��������
�#}��u(�׮���b���"�øgަ.�V��Cc��P�	4�1��_G�//.g���>y���/���Җ�åŬ��T���x��v�������;��v�n�S3%U�	Ou�����=&�"�K:�mu�t�Ŋ���)�4��e˭���
��yT��Y}B���/G��@xր�}6�{'V�{n��X&%��wN�,&���u&sf.�ց�+��jr]*���оT�૤�6s�ZE���#ď0�m�J�lO���gZa2g:D�������;��hָ�4Y,q;�7�j��L/���߶�V��r|՞��L������B�ڌ���П*����kD�n��}��i�t?P!�ܵ�=7dj)-�F�.�\ϲ��k��db�#�pR}�Y�mT�}Xn^,�M�Z�|/S<�w�V�@]Us��1���G���o0���o{�n�.'|���E�oOs�2V��u��)��j�5u�.j���c���Ҹ�Łb؇�[���^휵Z�S��T:}���V3,�\5��ڌN*4TnN�\�Q�'d!n�֠R��Fu�	�]>k���N��"��"EWw&��n?���w��Ӻ9��o�Ev��퀮�=ݹ6�Y�vJ[s1�w䗹<g���~s��q}��}�ʛ؋����m��78󞌱c<l��^w���������1�$�����{F�7\���t��b�K�Gcr��X��	%�)qn�v��%�;眞nk�����������N�}n/�^��DI[����.�e���U��%�u���9����X��Ǝ�\WeG�r��ŕ)֎�) ����f�ʶ/5� �}s<�}1���1#}w� �x�U�x>�}�Y�۹]9c{��VU�p���gR��@J�zpPK@>�=�{k(�=�j�.���3���e�7�Fa�nK�|s�6,V�h��ۏ���o�/��6bM:S<&�B��5)�8�ѕ�(s�����H;oL^�o���A���lr}oE4��D:_`�i�;�;CX�l\�eUV���N�Ne{���� �?�V��1SU4�~V��ɵ�i�З^�}�ƅ�{�*B�S��z�H���#I�r��CL.��p%��ѹ7뙝3�y��q�H��͘�ިW%��doO��M�hz����ou�8��i���,�SP�.���u���f'=��Eoe೻7\���7�,DO�+����)����]�0le1us�i���y����������[m�C�:Jx���V�ۆ�X��Άg\�=;#��oiG�yF�xG [C��P@QdK�Wgpcx�ì��Z��`j3 �5ֹ���j�	=�r챊�7�Ǔ��測�5�-�f�<H�{�#�8r֬�U�p�mBo^Qg{��kqck���t����9~��o7�F��۱<�S�i�O��0:Y��}1;Ǫ��U�-}b�&�k����VሿA��,5�×nr�隽W-A��n_�=����m<��c6��/��Ŵ�c�|(�3�-��\�Y�_@$n\w7��R��΂�v3T%>��t
��D����Ƿp
���e�����9�q��/.�m�Z�~��q��:���Cw��nt].���c���g*���ɭ^1J��'bs�����m�|�z���v���]�w���K�Hw����q�X�t�1�~��=���/�2�3���U�ۓ�~�<�u+���6.�,�6<Rjޑ72tyӤ2�޺����	�B<�����;�r�x�����u盟���C��޿9�PAW�������~����� ?�����ރ��<�A:�=�$��	�	E�	�E�E�E�E�	E�$:�Q�U�$V�XBQaE��D9�C���@�aP�T�!"�@� ! �@"!*@�(���8���$B�ʪ  �`BQ�	!E8�"$D�P`�A B�	AB%Q�P BP�U$A� BU@�BE@�	!�A@�! �@�"�
J(!�@� !ם �B�! �@���JJ,J,B,J�B,@/8�`BQ`B`BT`B`BQ`BT`B`BQ`Bz��E�	Q�	�	Q�E�	A�e�XB`BTy������#���#�] �B,J,H�B,H�@,B,H,@�J/����ϐp����*(�*�((�'��z����|�W����<����������_�����|���;��S���������Z� �������c�D_��ʈ��@��c�C�@�ڟ�/�����j�*"
���A�?y�/a�I�C��>��?�'�����A�C��+���*��
�%* "%-�@�P"D�J-"%�ċ2� ����
��,�4+0,+H��H���0-"�(���@��,J�2�
�(�)
Ҍ$$,��$#*�̋"J0H��$ ȴ��"ȴ�,@�
�(��,,�� �,�,²"�"�(ʄ,���,H��2!�"��ʄ�(̣"�$��	"Ȅ�$+0,Ȱ�(� C��,�,,�(@���H��$+,B�B���ċ*��@�
�� 0 @-"īH���+,��H� ��(�-",��P$�@�P����*P(�"Ҩ�,J
�" R"��H  :�!�����_�O�E(�DD(TT��@��������Po�~����?�? (��A����u����	����Ï�����ӳ���DAWC�!�I�=z�S�
�*��DAW����?���
 ����z��Q\���i��.��z�A���9��'�z<�^à;�DAV��/���QU���(���W�?pw���?��$������AW?P���TD@?>�v��������|O��?���A���ߡ'��� ��e?>�8����?o�:������W�AQ탁�|�A����N�|��C�~����d�Mf�20(	[f�A@��̟\���|�}P�����Q*�)� �JU$��(Wm@Q%I
QJ�$�kT Q@��T�*Q�$�D%J�h�EH5��m*(�J([2��2	#[k3ej�J�R�f�$��ٕDQ)���m�QAU�ER��Zj�I�-����#U�Z���*�PP6�E��VƄ�E�V֣U�  Ei�ZԊ�l*�QQ%)RҴֶT�j0���B�(i�l
$�(� q�|��ikl�YV�U5�騻,6�e�h����w5�mZ�� �j��6��ڊ�Z���as���Tֶ�N��խ+e��m��m*�EڶZT���X�R�b^ ����B�B�Ql!�{(P���Cܦ��i�Q��-���E��e�mf�&��ն�QM4R����J����KR��)r�T�۵��[kf��U#6�Zj��h5K� �<l�ZV�)f�աKm�i�mU��i����n��٪��L�UUQ�e۹�4��[)�F���Tڪ�i�s
�AAtm�`1"֐��  ��Ъ���mmlЌk���fm��ձ��k��8-��j�
�aVf�m�Y�F��e��F@�J��TH;d�6b�h�j5��A�  ���R �j)h)&UH�����#`ec;�̶���[+X���@�XE��j���GE]1UZ��N�isj��m��Z-����SZ�  ��UZжH�Qlj�P5$�XXQT�40 �d �h�T((�(�	� ��m�Pˬ�i��R����� �� ���&� ��� aݸ ��� ��aJ �, ,�[��  ��� �wb�@
�Yٶ4�ch���ʪ�x  ��  @۠ 8w ���  f�� P):0h"�v8 �Z�� J`�T�6+ A�ݛl%
�
����Z�+�  �΃@(��2�(
�F  Q�8�� ������4�  �hh4 �J� J�L  ��.�lmQ�V� �  �� i���i� �,� 2� i�]84 �  +��  �` hQk��  ׀"��M��) @��a%%*�4 �~�zO(� )� ��OH 4 �~D��d ��H���� 43R������0S
��$�Č �Q����C�
�A�8m�:���a���g�}�g�}��j�Z�{������ڶֶ���ֶ����mZ�[V��ٵkUm��~��������Z�aLâ�T��**���͊st%B9P%f����݉��j:���Z�F�+�nY0���kj�)�db��r��N�VTiM��em*T ���u�1�Q;X��B��eh�>�!Ki���Q�f%L�b�a��13�Gn���b����.���\UX08��D���Z&�弤㩍J��i�MGr����0�lJ�vZߙʹ4Z��e���ء�G�bfѹWi������ei�m�a�0�훺�%�����tHRQ�τ�Cok(fU�kV�1 �52L+�s?�pl2Ys*
qQ7374[m��ЩaQ�(R-쭏>X]*���Zgi]�{-��e=�R�icGeAAWi*v��%m���*�T0mXC��+	�#6`PI,(��s,�Ӹ��hȖ:r=ڹ)�"�j�,�H���8V	��`f���A�v]%N�(vǤ�Ff��:���Ӧ~�vC�B6肑5x�̸uw��NU�1崑�e[�u`YN=��NcȜ����nV�K5l ��۲��h���v�)�C5f�Ĵ<�BX�\�.��X��FFn�ى��ևmtP���8/n��)6�	�	��9l0�ӔFӭ!ٛ�%Ik���)<@e�Vִ�^c�¤�1m��S�fh�qS���L�ݫ.���镚܎�e)n�f}�Ɖ)`T�ư첫
ԫ	v�ǚ华X"����/r�)�_<�yQ�9�f��;&k���'�C�xf�j\"E��]fTz��T���26��B�unV��ML�ђYu�,�y�S��?Mє��
&.0�͙1Jf�:o���PX֜�@�d4���6��,�N�<�gb8���VeH���b�$B���db�5S��Ќ����\.Ga��'E�ƞ@&�˗i-�F}Y*�M�h�SCA鍹��3,46䂮�̠��/2��^��)ց��ً@,n�4,�$e��|-7�+(F�Y˹t1d�*���Y��j�Z���UM!R��EYY�ݼ2b�ݝA<��Z�"�VȰq+J�a�Rחj)�O5[ycf�G�"���/v��Ԗ�e�U��K�#z�
F;���LV"1!0Xbb�x����'D�f�e�3^�1�c"�-��L��%�nVe<�Hq�B�dQ�
��N����[W�,0��!0c�٤pb���(3Ue�Հ���+�%�l�n͙��V�wS,Y��-ZJ��z��+	�1VX!�ܤ.�1�sV2�Ev���-��)e��ve��LKq����	�n�%i;PTJ}��r�:%u"QQ�lcH�p��x,,��EKX�Jԟe�q�e`̔X���vnV�7R]�b�h���ݠ7��ˊ�*5�ʍ���w`g���D'N�*۔�cm pmÊ��@�h��dN[-�����K���S̨��li�]��7�6@�mj�4^ǟ�B�D����%�B�Á���2^7 yFR��Xr`��U����YB�"�4���٧h�)�l^�m�3dD2�R��v���Ȧ@T�Ĳ�Vn���MRY	kݐaɸ���A��̥�lY	�+��p�KاX�v��ùo ��
�Y�H݂��n�Ƕ�i�b��-��9P�l��ԮR4+#@�B�X,�ǥ[[I^�_ ^F�i&���ެ�܂��� �Y�,5�[j�n��r��"E�d�֊N����J��&�"����WJ���zX{R�ɕ�0��2D�N	0�Ӏ
� ��#ة6*��y���҇/eEX&�-�f�Q4�Ŕ��ȱ)A�����k^��W�cƯcYc6��	ؕ��\9[%4���U��S)���cR�/fX�C5�G&,���9(�i��!�4�Ɏ2��?
��}��שA�h�&�r��(ZI
�n�hcF۷EZ_5�Q[����P��n��N����5t(,"��[U�ܵb2)�ۤ�h�a�6^Q/	v�3]�ж���v��9��^=��U&��3*Tj=�3�T����n�A�E�D��%��"��;M�2ja�-v���lB����*�T����p����ȩ�M�sv���fHt��5U�OL�H���¬ЫY�͂U�;�Jː��75�{�7�պ���k���W��ME&U�y�����x�=�vd�H� )�l�yX�#[��n��t@gh\�a��01eXsL�n 1&�Գ���З�b��AAC�^�-ϴ��,�Ŵ+F��,��m��
W4fk�B�-����{�����׸Qhԡ(�:�Œ,k05�j�Ҩ4�w1Y���Un�g6�+-31��ї�ȣF��+iR�soL��X2kv�9B)�VY�B4�L(qjӵ�$!e���6ɪ�R�������Z�l�s4S`ңuq[`�_N1CaNP1��u�WӇ2D3-:шnds� ��&V���[)����e�2`c����`�Țn�A ���Kp`�S0�W{�e�$���مA�+�n�[�t�V����0?����و�f�;�Z��v$�fa�)���WS���|r��6d���h����3!��p�!���Q�lò͡s"��t���o�2]�RZF����JP�m��.��lR^�I6�r�A�su�e*l9�@���4��l��VXbՃ����p��D�D�L<�P�B�諦��ژ!h�/�K�ј�)�#rrf��z{�ҹ�m�	Vrܻ��	Qgu0���4�q�P�f��:4d.Y�4ڄG�����2����:X�	Ặ��&k���hC����+ܫoa��Ė��@⫩��H�c}>/>+
Fͽ�
��Cx[xL͛�����ws3/]�Q"0ɴଭP4g�!�@��;*�pn�G"���BX�۰�Ʀ����H�F[E�F�CT�V���t�;u0��]���(=�oj,��X�VV%dV�7�S��d�f�Sp�ï a�M��8eͷz MG�mm�Z�@8٨�l;�-�D�����mf끳��]�����l����i:+j�ٗ7.�dl`��hTFb���,���ո�I��Sˠ���n�Qɩ]�^\��Fnl�ح9&
5d^�[ԜX��.���Wt�xkZ"R߆���#�D#E�v��,�/rcwh�5�1�i��/,�e��(�r�[�L�xj8�M*z�����Z��h�t-�5�ܵ���1E�06ź,�X��qU�;�ZB��F�s]f�YN���j�L/G>��+��h+ز�N`��l��tӅ�{qXGq��2�C%�k��!����h�l�n�%B�F��P��U<�`2�U+s7m1����թ[���]a"�^ĮV�ˑ���{���|᭼��;�0R�cwjKD�i�voe�%��C�_H�T.'�T�2քԤ���;�X���c�db�͑�q��U�t�`6Qڵ���3b�#sV*����7)�֙�S�ER�j��yi3����!���˥R%��ad�+TV�LٮcZ�R0��V�0G��6�zb����l�`���6�V�ikv��B,K�LXKH�s�j,��¼��&���!Ln�FFk���Y��V��SA$Q*�JZmaI�l!U�J�3�y�*�kt7�iM��h+q[��vDŖn��C�x��ec0aTX!R�*<Uӆ�ꚅe=�N$�Oo��R�Q��$G	�Z�d������7'�kE���̬�3��,��R��b��l�3��ɹ�S��Ź��)���I�"�40�
sk6�h=|���F+B��-ٔ�*F��{eXmh��v�!K3J�YG6�����9}m��訫�،�j�|�Ibv
ڄ�ʶ�n��Vq�si
��`i�C��h'.]�`�<\!53!ʄ���m���$�̊�w�mR�Cu@�:��:,*Y�S����U1�Z��y�4��Y��]T34���T�\����{"��衪٠�Vf,�5<�ݍz�Ì6�Sh�ѱTgB�Z#�u{�����64��Mь,� ��Û��1�*|H�2���M6�7X(|YӁ[��l��� ��-;�
��e���������B�M�ʙ,;�Q̺Y2򵭏wud:FS�Xˤغ԰��ak��Y�mۏ6C��F(ee3���kr�!�u�HY�A͉��eqf۴ �3h]3&*U�I6�,�x�X��i��Q�À������GxTnT�,�E��N9h�ձ�!U�^������+�PL`j����
W�&HBG^e���e7�Pw�����ش��Ҁb�u{�H�h����m�D��,y�#{c�G$:�-���12�����ϑЉ�\q��<�&@P1������-�,�BTݏ�`���, �-B)�٫kF떅ʺI�j�hr�Y[��+�]I`82�nQ���3YV�
]`�,=D+���Tr��T�]Vʌ;Ő�E�YlK�u4හF�����{F��k)^R�S
����[����ͨU��C�t6�y`�PV́�k��e��]�4]��{I+�n�H�p�v�%虦�� ��S����:�4����90͒a�;�Btk7ښa�*���te��JSbVgH�Z���1��s^�k-U�k1]��")1[Hn�r��8��҈
׻B�5f͈iˣ��Y[&nШ�z􌂑�	�XR�fR��-��;i����B�����*��5�'�n+��$X&nͰ���Bb�c#I����˺�w5�	ӍjYYܵow@۴�ֻF���
)�"ڲeK��V�Y���@M������\�ST�U��2��v�gEBko2��[�>���#ؠ9K�
N��e�Ğ�)�I2����Ы�ǫ*k��IV�1��TįI�T����1���K7k2����T����L=Yh�Dk�k@� #����!)�J�� ��;�(�1�oU�&�3�q;�j��V���hj�wf�5�Tح�x֑�m�Ysi�؃4�,�0��[!'歆⍧� ��`��l����P��dS�+v��O���r��4X�:*0ˢ7���+��Ft���*^�u��r㔙T�x2�Q��n����7�*R��
��{,��XN\�2�AW���h ��)υG���Tz�R���b���*e+�1�S��Q$7�-:eэ�Uw��,X-��VՄ�N����Y ���U��S�2��$�U%�6m�N���:(���4!�\B�$�0�ًF�j�L�*Qi��W�`fIX���ض�^�9Z�
\&�;�S�f�WH���>/0V�,E%�E��
�H�V��&�+(��X^��`�ϊQ��me�ǹ�,�G�C"�����B�A�!`��+К�cT۬���3� g5ĊkT�V,�&V0*dF�n�с��n7y��c��Yf�uw��[��X��a�WD�ˍ���QSVy%�D	��%�AQ�����]X��gN1P22�-鬖�`�wNT�m����9+rWtn�5��XN0q'jn����*��"�TšKH��ӽ�]�b�j,R�y�@�Nl �k���iw%�&�T�1����C����֖f�[F��hd̦�[���K0m�gn���:v����a*t���CA�f
�������+�7S�(&70 �k�Q�:��m���g~[gY ��)+�����!"��#v�,.Ze<����V�$X&j��$����ûf fk!���R}`Q�-��L4���8ts0R�&��[�Kŷ+qh��O8r]��>פ5*ұv4�c����[��/U]���峊��ۥ�����(lM��~+*E��`4�y��� /�z��ԩ��:.��#E��b�)m!�N�#@Xٸ�PP(�Ocq�]��Գl\�y@U�Y���.ĭ���b�-(/�f���ADr�U�[f��3p�J����-�B�����zc���Ж^�-��ک�wR<�zU��	�A���O+w�X�pMV��zԂ��2Ģ
���c6�ҭ����.���,��-��h���躰I��4CO%/��%��I[I�v��,Y���A���w-���!Zxƍ�)5q�<L�eZ�J�ȵ#�ʚ��hʷLۃ��̧�*��J��.-+j[ۥo)* �m�u;c7@�U�XU)�&B[	ƆU���а+��*
m��%��3j���n�,6(���f��|���$���k�q��3R2�z:����.iN�o֓�W��m��2[�I̫Tsi�bI��n�Bq�-�nͅL(�y��f�tn��6��v��L,�Q?nL;
��+4��j�a=�rĬrh����Cm�2�]`-��]iW�n1yH�u@AG2$⽺. �4��N����{`ڠ卵����%]*���9*�SŮݙpeF�ڃ1�k��!Y�7IQ-�̤���ǩ֚[xRyU�n�p0�iP�ݗlڰZ�Ow��n����P��=�b�-��eiv�ۊ��2`�S ��2��X�Q� @��B����ZkU�5��"x�PZ,b�X�&C�tEK�{�B����t�cP�7h�*&�u�,(��:F��Տb�tv�dX�a�&c�2RR�n9|mn��X�o5h!7�6��!�t�|�#	�ǒ��W@$�h^��f=Y�n��寡���eژ��P�L�ֈ��u�&� f/+"8��e
Ve*ې
�L!�+�ܥ���cF䙄-�(�j׌=z�
50P���X�|l�2���Vk���n���CQٳݧP�s[�.weN4%餅wGsS��\�2ND�r�}d<���)��{EQ�dQ�ۍ3b��3N�>=H���.�n�+pwp�F���ԅҕ)ٔ*��ޞ1nm�SBt:PtJ_2�ۼp*=�q=h�V.֦�L��P�jÚs�sD��f�_!:e�5؅�m�Ng�༶���*o&�n�C�	��t�f���M�
�YwU$|�n'5vݮŀռ��'R���,��F��}��$䕨�WZ΢�غqR��(��jR�T�t�8��)v�E�U�u6eZp�9�;��L�����.�����g�s����JX��M��w��9Ē1��
+@��-��n�f�6a�J�78��jNO3Z���⦽�����OQe��[.�j�q��u�4D��hub��XdLnE�w�,�7�����,���B��Y@r��Վ�\rY\��	�=y�Y��;�gjErZ��@ݱs�-��=&cEܵba)�\�޹�����!S��\�������t�l�[v���O/2E�WY�� n��)�i�ۘ]�mF:�i5�&"� �]&��'fܮkjʿB���9�f���v8��368��,l5� ]�U��{QKqջ(�8�u�x�:�!���T������;FZ����J���h��*f��Ո���BŐ��Nh��/u��$К�*'L%ײN51+�K��Ԫ��k2�X�����w��/�.p��1S>ז�:�݋]��Y}5|r�wx�=}�7[��,�^�+u_qܔ��m��B(�At�ٕٹ/z93�r��)y+xH7�]d7�a�f���Fôhfޑ�ǣl� 1�X�J�������5�eoY��*P{f���=���Kh�-��R�$�l�CW�_tu�7�.�q���0�3��=H�໭�����IZ5MK�q�9_���f�ZEK�Ss3':L���k�/��v�X�O+��D+��o�+%�W�rv�:�N�t�5`�M�J-ޣlu�T�;�IQww�e���\�R�Z��eh"`�!|߾GZi���.���e �	�4,]XU���V;~D����:�^��o8%�������lƬVn��3����� N
ۙ����hR܆�or����,4�������v5�"�&U�֮�NR�U�S�E�j�0�ٚV��"�j(�N�|p�v��ڛ�o�o���(���I��[�O���K�ܩ�R�.��&$��uۮ.�N��
�T�4��0M�:bn��m_\�ں�wI5R�o��P��OmT޾T���v)���*sil�7>s0�f�z��l�2k���\S��Lv���W9Xa��H�˒�g(7��Ej4����%���вR�\WK�������:W�V�nt)���wK6��N])g����Y�i,��b�3�C�����v��p�wخV���%�ɒf֝ղh`��Q2tܔ���#�$��%��ز+W�|�w�u��Y�2X9��(v��&�)���R��"^W7,��m^}CPS�V=ھh���*役�
�m��э�ʵ����T������l���=%MS����gd2�#���Me�5a��C\�w)q�Ֆ�Jj��-1�$���}�T-����Iř��p/m�a
幧3MN�]��eue�n�w^��>E2�T���ǣ�U�K쀥�N6Ї-cFa��f�����6^l����1.�P�VЫ��ݕ����d�n�-��������:�Q<U���wJ>����!�����rޓ]�#,��JA��M�P.,`�+�q\�V	N�cw���3���Z�3N4&�,�b	mh���`��9D�Y�%�4u>�r�R���t{2�̷��G�f:�X�+��eYw�]�J�ee�Qh�jIP����2dv�
�Q՞yvN��oԀ�cdԴ�Yc�8�����K�����ɶ��I}צ;t�q�@-*�Ҭ���O�}J+����P���#�i�%�����N۩.�PX)�/3�h�}�2l(6�u��� �����)bޓ�f0�3�\�<�[�HVo�LP�ċ�+�U�$�q�6�^R&�Z�������Z��|�����堩Y�n��r��`K���ڹ:Q5iQ�@��鲰Ц�X�b���n.²�1f�x��q�p��-�`'YL��lU��i�)��,;����.���>�B^��)"�믱�I�t;�7��޳����2�C�� �%M2�sNIh����&�뫛�wK�pO�O�
w�ܖ�x�q��b檏��.�wJ��kZ�C�v�t!���ýo��ͪ)��4���NQ��w�f�浫�_jX�A:9�mn7��w��em`�i�WB�魱9�3;�b`�����5�+�s�cwM��Ku��Ek!���g��%޳���]���n^�n=|�9�"�ݐŮ�#n:[G��Fwv+�����E��B\�?�Fjv8��`;ª�:#��Fyv�α`�8�` ��U� 6o.�Z���DM���/�(�M�v�t �õ�I�/o8%jT�Gh�񱶗f�-�1*Y�޵yB�e�G:�8B�6��h�f��)^8g�l��R|�su�tgT �Fr�y�:�ƇulVC�`�Hӻ���	c˧�|MX�� 6���� d��/��]�&�+ဈ�rm�[�P���:�t@cp���]�b��U}��S��L���Z�4�fج��+�T���>����#O�}2�d�+i6k�dt����La9��'�������` I��T3��׀�J��Mɜ���p��XE�y�ᥦ���3.�g�L��I�R��u|���f�ݢ���4�]H]���*/Ob����h���ڼU�ܙ0�}�����$�W����u�<������cK���f+�;r��P�: �}׹jt3Wk����j�:�S�ݵ�^}�\=�<�ܵ.�MtKiG�B�LoN`
��6v�u0"�������z�s�,9KY�;h�zr�,=��N�A̵LtG�s��]���)������v�s
��#��
ɒ�-3��[��^Ӕ���"���.�AǦ�;�ko
�o3����&��1!�VN����@�:��O2#u�*�3��|�Y�Q��_F�:\��ws3�M��i[@�!�Ƹ�<m8e�~u3��r%7L}�nan�K7�e>��m�jl�O�6�/��e�tL얄1���ի�yY�t�Ck9�aeNG�_gvԭ���y>�������}�:g��K��8򦄘jT�Gd��+9	�;�����:�eؠ&�7
�3�B5E�%�YQ�ι}c���;#�-����K��!��7Hڵk����l����a���`�V����b#Zf�zf��`y&��/�8�ɏV|�n�m��#r�@w��r�*o��^%g�r��k��F����7�Q��(���v4������q����-Rںw6A�i:�DT�K_'I�$�$���S�]���0��YQ�m ?#�,Z$����w9ewNi8}�+�,:��WS�6���jIC�X��^�f��HR&V�,U�:y2�����軝[�\U����Qk���T�Y��0.9|����o�R)��4�`��n��k)EY-�ƍc"�8kb|%i���1L�-�a�9�2.6�]MHA2���w+��6�x̫�^���yN�Nw�J(���Ca���^�;�0-C"�g^�f�TOs]J��)m:��������9T}�!���=�"ӽ
Wځ�<ή�;"48U���˨�J륻�7��[J�.�ϱ��P��:Z�rS����Ӛ�jF!󦫳7o�3�wӱj�_�}����g�Ř��E��3�1ùj���=�]]E�*��am��Y&�ٿL9�ݧ��Z��$+E�m+g��Q�,�|�w�7*�C�'�t����*�Ĭ���n��%&j=ʊ��]�NZȔ��w��CE�%I�ɦ�h�̕
h��H�^��ɷ��D��oaN�n��9���6��3Ṗ�	���5+[�-�ә3���)��쌝N�qe��\��5t1- �κ\h�n�����eH{6ZI��\2
u3)�[�v_=��&�}�M	:n��N�����.�
�P8`X�̺=�6��t������%9��j��.<��W)��yJ;��el.���/��R��*��x:���Fo�@�M����<�u����}n�Y�ש%�q�|�}�(k.�m����w�hF��N�"�β�<���7;Ի�q[��t+e��!g����ȫ�4k���&y�� ���38ۦ��$�$�C�P�UM��]��=��Օ;�)�ϰ��;P��X�cO'�R��.��]C�۟b�,Fp�خ����w[3�q���w��,�|P�U1n���mG&�W���X�<�a]x�4�m�������&y�(��}�5��f��0*�Ջ�H�I9�Y�g�Ὅa�%/����fm��ȑdGk��[r��2֬�9�W��m�E���T�u(VhL5K%�3D<�b,�ѧP1�>��֠ 40b{|!Y��닡Á��4��ŉ�j������Ҟ��XI��`��0������bݗ�N��n�	���qb�j��g����K�����ճ�5��M���u�@g��ޱ�:�v������U�����.u�w�<r��rVj��ò�F�R\�sDEI͊
�t�Qne:��������@�����y�!�J}{���K�4
e��<�Q�ց/3u�Ȳw�q�4f��?�K`��v��I=��:>LM/��L�雓*�͞��ϩ�̻��*cbG.g'ɮ�*Xn�C��h+��������x��gqI�VK}Fݟ�o9^o-�,7ՊW}	�>'򒬍�dB����뛔�M�n2��4^�\��;`ꕢuo<��yo>�A���ֽ��Cu���Ӡ>T­��o:L��Pݣ�Y���ˁ��"i�N���ʰ,�ن��Q��k,�yI� a��W�^H(Ǭ^u�0Mk��Xջ����j�6�՝,Lrp�zo.��R�ٍ��P,�*`]�+�׀�4��$[W�&n���`R��#_>�.x���=����Ñ�}v�wSz�F�>f��.����\��Mm��4g%V��5Xo�nԹ�I�{h�;!��,���tw�}i����G�!u\�Qﱃ�n*3]��*�Z�Y��З�]�ΝǱ�j�ފ&�WS&IئU]fM֘��_Wwh�����S�=�n��K�~^�Sd}�M
�ڻ��BSٱ_.�q)s�E,��(:a/���x�u��Y�3�-�;U��n���+$�֌'@�[�Fa �4m���2��äw=�}wG,���E>����Wc�f��Al'3��5t�v<|C�B4u`ҏA�� ci�;���u��m����h��2�Q4��e��
=5�ξ�H@�v�iy�D1��b��{)�6p�Clg>h��c�����i��5�gfn�����.�Xnᄹ��!y��Ւ�IU�Wwm�\�Ǖ:���*;E>�o<�'�_+�9�z;�JQ<]��E]mJ������X�5-���<fq�6ZAXY��l�t�X���(t�7��W�����9�P�Ɓ3R�]C�J�481}�<�n^é3s�����c��y���$����;�ŷ�[BP�xM�Id�m���Oz�ox6�(rN�+�;̝^u�Ae* Qɾ����v �;i�u�8��R��nͮ�h2��'���|n^�a��\��%�&'Kp5�o+d�Sސ@��d��I#�.n�y0�Ç,E�C�O{fC�Vi����l�I� ��J��vsz뫁��P3X@=y����*��c59�)��Y��rRAW"	mn�]v��t�
˧�1����,�MZ�VmC�3G�QӲ19V��lѵ�z��
�'����K�cN��+a�^R���܅,�g^F��-���)��Ǉp�i��o,u��C;�ES��j�jS�-�#l]����m�5�0����(vi�G:b�r
o)��]�]���LS�w4����Q�>�z��:�ihP7���u��ݽ��W,��dv&�v�Պޤ��@�Z݃�F�/�����Xf��=��u�����J<��kGp7݊�V�:�G���.G�;�L���>�¤GN�ZƔ��s��*:5bSF�j��X{@���2a���|(C�Q�Z����y;{�W��]�Ӛ�NJ�f�Ұ�d�/��psօ]�8Zi8�1�z���`�
� ]f�.p���q�M��5V�w��+�`}�N��-^b婤u8y�n�'�(-9�\P�f�����&јqWl��:��\-�WIAT���V�۲l��3�s��X����V��T�@-Эo5�*H#]ێ�[]�X���ԖA|:]ڠ]���w��������f��G�w#�yүrSbt1� o+5kYy��8$�V.:���\@��	f�:b�Ǯ�4 p:���D>�y}Ƭ���>�ze^R��9�W>�f7Bй~&p-(ǆB��.���.���R�������<�K�<o�hS�^4[�=��	�ۢX���P�T�Px{W|�s�)N�jn>A��\{:I��z��V��j�0:��ʓ��I6m/l�\�0.
� �iv��Z۹h�3Du���εPV<H���;���ؾb�*���	wA����B�6�����SuޓPή�(���ao
��vr�%3������Of�X���j�}��%�h���/��i��d�%���S����3��Q����t���1f�n�/�s;b!��Q��<2�}n��(�`�v�geA)Byj
]Y=� #�9�n���3���Ή:{�rl��!�9z�Y���".z+y��j�ۋ��'�w���9L��gd�h7�����|Ռ�.L�}�w�Fi�؝]���/���ŮU�z�5+��呛}-�������}�fe���U������;��?�y�}}���������i�	Vٳ�i��5t�ѳ��E�N�����^w�,�'|Vp����N��p�܁zm�ڳ���XU�w^�8bzD�Õkrr�I�=����ҙ:u�-��زi����2<��;I.|2#L��6k{K㷵uX#��>f�ܥXsDd�8%KzN�7�)�-+h]�5M��yh�Ӧ/���v�jgV3ݲ�`��:`�o҃�Vu+2�l���Acy��� ��5�]���Io�eM��$t��a'��T{�[dn��:��J.,S�-t�K�ʳ�
к��Y�n]�O�M,�"�<R����dY/�ԉ�}19��\^��u:���z�S'����w�@���R���t͎Σ���osfJ&�;Ge��/��#�p�<�D[���-�
gm��2�4�9ݴ�}�M��ġwh->�r�����ЫknmИ���/�D�(�|�IQ����H�u��r���9+�SE��+���-!VŖ�::Llb���+3����ڲ4��k�oMr�c�K���ib�.W ���ᶥ���WZ(�����mfɽ��^#c�2+&��ήQ\#:�sa=�@9�����<XJ80��[�zI�{�?��769���,�Q���[cq��28��	vzY5~�k�'�E���j$�-�N�g:�44��k�ݓS�؝�&�k!d��Y:��sVm��'�j��*����}����a�ףmrnRW�(D�q��-
��I��ĭI�^�oB��=�a�p�C��c5l�7��v�J{Z<�2u #Yh�A]N]C1��C������}������9����2��[α�қ\EGt0`�j0��s�7� mm5�7I��TS���&����={��[�D�wv�,��8��pէp������eJ�ʊ�ٽ�1Gn-�	b׈ח��D�N�@�نk�����M;z��F�R:tW].w/B�]R�\��i�ǫ����2�H7Pгpv����U��g_r�Q9*��>#��vMh��)�ƾ"�q�U����d��fõ�{�ʈ�]ȕ�w(�.5}��^���!b�ޓ3��u6�H�lfܴː�P��up3��;�(���7��k��;%"�^KKa��@�@������K��imяV�mPS�`�J�T�.9�'K+M��Q�fZc��b1�IW��ĝ�����;�&�TtOR�v�Oa*� ��:.s7�jq�
l�@��f^�"��In���Ѭ����H ;�vDӳnc4�%.N���n�w��ǲ�5&rLeq�i�|;x�}2�1��t�:�q���9���g_-�sf�_u�^�K c����EEo���[E���L���e�mV��`�v�
�Z���&s�նp����k��S�\�E���@KH�#!��f:�NH�W�t���ټ�x��jQ؊���v�1�8� wX���&�݅C�N�� qfh�͠.�6-�8�e�)�O�ea�t��լME�8���M�G���Dګ�v�T����].�q�ٕ���N�FKJ�a'DG0�d�&}	w{^���ō�17�]N�Q_P�|�9.��r2.��Vr-6�xxg�')G]r�6�e�e�`��d�;Q벗'��:oJ�Ӏ��Sì��k��E�[���;�-�/�5èj*���4zǷH�y�>�-��6U^�ٍs �{��W�.ް�M�Nz���N�t'SbÍ<��c���nwl��];yZ!0k�p&�lrx�,W��=)��A�8K���O���R��.�7Wt�Z�Z���U�K��5���Ar�,��R|�Wf4D�.tt�_P`PQ7����5�t���g۱dpX\G�Ɛ��3(��9���%���u
[��kKNe��r!����b�J7i����8��x�e�eV���粹[ �eMӆ�G�A[��#J��2`4R��$ʻ����2v���*�Ό[Z�0�~]�g[*N�#G��آ2��x� ��`\��%��mյs�c�Lu�=�<=P�2%��6"���=�B�qg=۶v����Ne$�p
���f����r�]��N|UfK�%vJۇ�_|�wu�U�,���� e��Z�9���{ti5�!��HŗRJ�|�9ݺ�j�(h��ƫ�i�G_\��@ݺ<n��av7z�����\u���t���" ��kWL����<r�T��tά��
:����r���ק:�|�H��Y�
����r�-�Rwny��C�a�����P�L�I7|,�B+��ɏ�]֍��\h}7V䳘�p%I�B�R�t�/;x̗t��;YY�l:�3Ol,�}�eņ���
$�n�����Kn�S�y���q��n�
%U��[��.D��:�;�*�Lo@sb�ȣ!���*`�Y��e��.��ۙv�-jC[��w2�V��u-e2�T�Y��K�]y�uV<xR67+��'�A饽ס�t���w�˥�i!s��Y��T����v#g*��+>�F'��a|͈�n�:�n��,
�]�J��-	��z�pw��Lj
�tH̭0���g�ڢ���q̼���V�}:ZsY�:�B�fmi�s�_,�%Y�d���wbhK�E���Q˳b��o�{0t��N�u�rEvw���O;�>�`��uAr���jgt�1K�=�e�un�ɤ1v\K:>�,�l�J�0,.�g,}��v%�9C�s�Do#r�N�L�x�M2=��D���м�Q*�Eʮ���+�N��K��WATV^�MgN
�{�8dK�z%S3f:˗iu�x�B��/��c��4�P��,�"N�]����D��S��o	��)t9�f�L=�!��o���32���|w1yixw����ν0�ҏ�x���ӛ��|xV��Q��b�] �6�A�������<��n�<����a9�z��z9Bf��r��8٢�WÂ"�YE�eDb\	�J,��+��w�4u+۔�Q�*<=�Q�e:G��w��4�k�������v�1u;Щ�{ۡӘ�f�bv4�o2�v��^aHmd��Tr�\n��\���m�DM���
�ma���U3a�%ա�L3�Qe1��\�;��;!�!� ���;�ּ��	�oS%�����S&k���e�c�^�c�4.!K8{�%�I�=]�Л�n�bܙ\��r:3�P�ԝ'	pbn�vå7z�'��( V�Y¸� ���*L��n@l5nz�iE9E��O,�W�#����G�5����}F�YE�f�;����{{��H�q�i��T3h`��(����1NY�v�9B�4���]fS롓y�sx�1|&q�f�P�U������u3�!2�G+���4�Z�������W�υa	V�rR��B�G�mw�ISu3��˧�L�c+�[ĕkJrw��GFŷ�; 	�B�_b��N���v��M\��I���!�]�����)�Ӻ�j����<M별5�Ń��!]�)J$��K��w�ᦥ9W�vp���YP�iK�I ڇw�zw6�Վ��u��Αp2dպ���W}�iޅyy\���k4��p�A��(͊�+s���L�Bn���L�f�����1���]&�
�[�Q��<��2ص����s�5Pݸا���,9��3��w�_db��rM�Y�3,�`n��A�ju���t�N���ݵǩ5���3��5{��u�(2o���7.��7}uj\Ʀ]�.$)Z��5X��8�����|�י�2=֛~åR
�c�a͂�Z4^��.����M�"�>Z�1��e.�ŧ;!���t��M�=�a*/�J��S%���i�M
�s6�����W�bI���Q
�]mw_(u��/�9w���Xh�w5=	$$���J��Y�X�;P�\�V�F�P�z��miN�wԝ�ۼ��j�n�o!�oJ�Ȼ4Y�F�X[SWoq�B.`�Пٕ�E����&�;z�)�k:葤�V1U[�:����؀G{%<�7}��h�3�I�l�W�9bvX��u�����.�ˉv멹.o��/)0�*6�M@m_oW��.�s�q!�
���ޝި�ر�n�@�A�%y�j1�"6o����2�%0MṧEoohؾ�jJ�M�sm��C+A:2ͱx@�
s��M�����AN.�]
'�*}٣O	C�� �����e��*�f��i*G����ld�%�
���s7D���˦z��ek�]�����\���:����i�+o}��YYيeΥu9�q%J����lG�T�]�,�:k��,<�!ܢ�Q�l�n�*�'s���[+�5�3��8+���f���k-��
@'�i�o��N�Wr�1EE���[YI���+kӒ�u	C��������Z���J���iʝ<U�.S��d�=��f`�Ҧj8ri7�mL�Q�}���}��FZ1Vh±�)��pb��E�7Ws�^n
2�"��(Ț7>8��>Q
�����C���(�NN��6;p��@�	/:c�U�{Xa�Y�J����}d;?^P+�7�.X�h�l��̩-�--��+K�Q���V�IS�԰�:��t�r�K�S���Jnx��;N)Gy�?��Vx5Zu����7�u͌��L�h�M�Qݍ���q4�:ݢ�`�K5��"��a�����p�̛����m>�ھL�/�����]DuS��曏�4�͖Wm�&��ɺ�M(Su{(��+3��<ǟD�p����j\�q[��P�U�y���*/F^�J�wg(7�Ff��Qa�0���X��<�}r���J��P*�R�F�����8]�A����o&U��mÏ�m\����V!�uݳ��
ʘ�ͽB;�ӹyn�m.t�����]w#�L��Z�e�Ųa�w�N���us���C�x.�U�WRr���gZ�i��]h5{��9��c}��������JA��|��,��۟��v��/��W���i�ށ����Ɓ�72�U'�%:��khS���3iM�^f3Y�n�7�*���ɥ�u��;xm�f�
����K;���O�
[z�<"�DP������)}Ʀu����:��P�z���Ԛf4a�I�f�!�ߞa�t;P+����R�n�u��Өf=�ī8�{��.�.��B�G��>��{+��,���e]�M�v�S{��C�2] >:j�v�V��n&1�U�ٜ�WU�`���2�g[��c��f�`�7J�oZ:�⢨f8�����Ɵ��uf�ɝ:��R�5(��p&�ɽϱ_%�P9f�H�o)�-��
��:1҄���ھcwK�׽��
6m�\0��qd�W�oG(��x��d%���a�x��r�u�7-�x��o.t"9{�Z9+�"���ܥ����V�L���Xo�
��1M��S%
��b=���i-4xbM�K�}&.�&ݘg^'����޾��F�a�ϔ9�Ҧ�����2�wM�[�N��d31�����e|EM�Wz�j��E�m�)�:�qW'��f-�u���/����hOބYS�
�4iĕ���O�7��]����6�m��;]r��r��ƅr���=|R�ml�O�Ӣ
��[�RۭfŤ��Yj,t��	�$��V>S.��������v�]�N�
���ۅ/�4(�Oh����U��ou� ��*15N�z�����,�j�qәF��`���t�eL�F���L(��}jΧ�.݂"3Q`���ה̬=�4�-ݭIκ:#3:�l�т�V�Q7X�d�Q�]D��R<y����{�n�AK��n���	 ���#M�W%	�c�H.�W+�;v��~��at���Mvns=oz�Y]�NŰw���2A�ol9#�}z��Ө:�k�����ܣ�mF��<�O�����:�P�7/{�ܨYi���`8om�>�Q�Ņ/Av���}���J�!E84�����]���q�Q�[	����̬����1'��*�S ���z���KU��CfM[�`���|ʺ��ýoA��W�ծТ�e�Ru������Ӣ'V����6sN
�r�K��$Zt�����I����qRi3�9a�F�N*q&�-Bf�+��7�;:�.[ܓ�}�xh���nyh���r5� /+a� b�L�w%w�ڻ�b�HS�7����,O/9#{�-:���	��odߓ��YO���."*�h��'v��Y<�
\����j�32$w��'9F��˻�Z; ���7��Rj���t�u�[5�q���%��N4�+̄�k�|��%��QW���&�4��w%	)o:�-+��yj��3�Վ"�)�ʐ�
�����LoF[�wA�鏯������rd`�U�&�����Y}eW"r_U���$غ���7V:��k��$�WX.�F��9���UŖy8�����+�bH �!,��Z&��yB�=��DR�b�6#�N�h.��v�apݨI����[C	��j�B��]ˉ=A~��a	�
����-�kxd�Q}8L��t������F���
��<��H��g����b���]܆/���;2��5�ظ'LPg^6#�0���Χ��1eq\9*�KSu��>�f�|(\��5*�Y�XMnv���ʒ.ޢ�0Ef�K]�(�:�l�2��NZ�3Ht�t��PaH.�_m:p[S����, ��aHe������rTv�Pq��x�䙓���r������w����T78;*�B+���_p*27��)F�U�r�c� Tu��&��ڳ7�VU�5O�V�$�����)�Z5�1gl���K���pn�*f�m��8����e��2�o(e�J�f�U���M�n�G���W�}_W�|���a��D`55�(�9��m� ��t�r�sj�6�x1�k�f#��۷�r���S�Zw��`��kѰ�[N��	�A�7sRͥu��x�ѻ�t �'fg]�TwG���︈,���-�g�<�*n��0�6��l�R�7dyH)Z6�{ո{Dx�^Yw�YU��3b�#�6w!�x��#[���c���IVȷ�"��MӾ��kt��T6`�$�hL;�K��M-���5��u���T:J�+X���ቷ�3\�n�h�;r��d0ٜBkn�_b�B����L���dӼA\��B��/.��ع�t��!XN���r�3g�.���d,�>w#�_0pwaՂ<:`�r�\�j��Cy2�^�r����ϕ��F���HEǜ�\:��{�Ԧ$����[���X..k�����F��*�e���5��A��5V�]m;�=�]7(���Z]];��H���<%�� ?>k+ѡM�Mkch�h=��2 ����+{xU�y�g6����Ѳ����?[��(��++R��2E��M\P��>}�kNl�o(WnWF+���Q&��{�3��eu�7]؎t[ô��z+R�6&�5���J[ơ��HJL μ�J�+s�N��.�U��E*�rl��:�<+=
�K�	!�5`���K�L�}6����TTU{\�]�hMm�ɢ��.Qsnk�1�&Knn���ccX���s[�
+�Rlj�F��X�"#h�5;�-Ex��F�*Mnj
��F�o;��x�+$s�r��x�د.[��%x����c\���,[żn���d��b�F�]r�j������nZ���;�Ѣ�F�1��lE�5�K�VwTk��m�i��n�ʢ�1�5��ߗ緯�˫;��� em(�+��,Y�d�L-痐jܾ]E<�R�H��{����/����̼�r��r4:�v��{1�t��+�mL!�`����r(��/�3q�{;ō&
0��eQ�;V
2�=۷w�r 3�c��4�g�sj��w�_3�k�6��c�*���@�Q
�mԱ@0�أ����2@h�rz�U.L��g�<�\S���K�[��6����e=��w��W�\*���p(g����?�B��*�1�1xV��h&����4;�v�����Z
uo�UX�W��E�˔̌�<����khؑ0�㖈~<�cvg����s���L0zի�6�� ץ;4����ϒ�!��?n��]�;O�W��\;��e7���8C��M�����X+���8~u��
|.�N�ᓳ�T���)R�t{�ʻ7ӯ��s5+X=���׼�0׷]�3� �6�|��Vz��8x[��j�<�S���ާx���$m�G!9cE��'O��� @��~���r�,??����i�=B��c�0Md:���׷1��h婆+�f2ẀοH�W:(�kp^��B��e�U���e̦e�-��#�@��C�F�AK�8��P.V�'F5#1�W]I��N��U����0$�Y2�ƛ�L��^���l�X�_�����)R"�X��vu�o=���[�@����C��l�Y�-���p��z���zL�������k�䫆ϱ}�������'/Mė�~��~�b7K�V�X�d�6���̳��k�^Q~ 8�Q�R-�Z�4�c�g����>�~4���1���=Ak�;s6�x�6g>������HŉK{ �h9Qxv�u��x6Ӳ_��eڴ�ʲ�����2�i��xJن3ƥ
��O�D��Y�L�X����:��U�9=�;��gor�����;����E�IIRG)���a\d�d�M��Og0����h�x�܏;𬀔(Em|���
9-�'"\���#�*�@����&]޳ �:���^c ����'��br���&l�S }��#j\pP�Ӓ���htJ:�zT^Ъ,w�{�8���U^1������C�/L���l�Q_'!������ O�x��6��4ٻ�;��_�y����'�B��x��c_cja'���bɤEAA��!��F'wّZyV�m�;�8��R|}�L���X{]zɹo����Xug�qO��P^>�z��}�G˙��ķx}� ��6'L�:8�>�,�sm���?2^\��+���=6?t.�:�i�[��ҟV�4�UݑEu�}v�.ɝ�5kR3S��sm�\�vi�7��u���}R����ມx�(a �hT�S��$=b�[�	��ڑ��Q$��R�T�X#�X6L�{S��1^ \!���G��^_<z��Q�t�U�*� ���|�x����!�(Y���������De��0�`�$;���Ư���iP�:ǜ��N�a�>�M�S:{2�h�.��l�}�p�u��j���q�-�K3vgy��΂�!Ù�p�ҔF̈�}�SW��%k�~[��W{!���\��\I��+��~�{�J�\u{d�:�Yc*Ү�%�}c���4��j���/G��e�=�{+va[���6rPES՞e��W1.�Z��7h��R��g�N��}�R�*cީ�"�3O��j��HI5ۮ�<z|H���5��6�u�)��5����P��<������ۄu��҂7��!3x�pU�V�70B�� $eQ o�͊Q�pT�S�h�+�m�3;o%�q�&���^�v{��+G�g���d��`���[�@ʭ�aWn���rcǷ�Ϻ��٭
��O�<'��<�uN��������h�䧓�F���7�=���*���ƹ����~E�# 
fPۖ�N���%x��w]�M9�L)����nǎ;�������_���A�VG�R��hi���'/��˼�*Ц���Z�����s�7umԫ��2�B>���:'H��ޥJ9�9]L�r轪E��$U�C��(eb�3����}���a��F��i^'��l�}^}��q��Ū�e��4����Y�^X�Ak��xR�� 7�d�Z�~x��^g%3=|�e����=ǁ.C�`I��,N�W]f?"�Պ*�w���ͬ��m�c�Y�i�,�̀+���~}��}��g�}�?Y���:RnJ�o��,^��L��/Ү/Vmd��n:}j���?R��.{G���]o���w��Q�-�4e|��Ǐ�7��û��j��m���HX}]�f�U��\�Rc��V�s�vO#S�[B��������i����@����h�9x�>��a�u������ɯ���}g�͏y|��F�6�C�3)l�^�W���5V+g��/�B��%~2�����G	�Lmos��\�g�y5��&Ϋ�cl��ظ�6{����)H��e|�>��n��7��%�7��g&�7�{�,��6�O���^1n)ֆ/�y��{�dV�c��O��W�5`/N�P=���w��1��ֺ��'}o��� 2��������ﮓʼx�VW��ƺ{���ie�c��U�'���=��N��=�U�n�>0�'NŦ�P����QXȹ�9����8�����j[����]��m���Lk)�s�[Y���6�{
ѥ��@��:3�{��
m��/^�ݘai�X���=��(�yPA�zd�%��מm��x�'��f����ڜd:g�W�
�!�i�rP�LJF�*��X�u�}�ϨL���i ����!����>�b��o���%R{�mP�0�g�����;ƫ~��
o}�UE|&�vhU�YBp{n�F0O�+B�i���ۗ���e�͇ݾ�����;�8�Oo'�X�ܢ�˅R��=�Q�F{U�
��w�j�+֕
����b́)��0H^�{��+3x �1�J��e��.g�7j��O��۵�C�Ǡ@Q�WxVa�k���^��%��f�� &T�^� �5�U�=c���(���zZ�e���E�p��.F��7lfz�;�B����f'��K5UL<�l� ���Խ����h�s��N�o�����l�W+)������/�'��j���L��d/k˱��kh�nA��Rs�O<�)��K��,�ߊ`��R�<�����3��~Y*��d�gU�6��K/�Gu-f����X�<�µx�$�R����Gw�ͼ�bä}`�<An�~�+A9�������5��s-l1*��dV�0.����;��6�������E[���K�C�i�:��ꪗ���S�͹���O[J&���T��8o�̓ u���?g�z�
��{�p����,��s���yv9h�PDdIC$���+�&����U]��7���DFX��j٨ j7�!��6c�J�� 2�sCv�����0��L��Q}GM�z�B�1Z�o�����V��k�>3�w�ז�ٓT�t��Ux��K8��{yk2�c�	C�ʰOr�^ ��|(����m:@�d=̂�a*��Q�8΋ɘЯ��U�B�@m���r�ܼW���!n%�g���_�-�q9>���H� mV �T`���Fp�cb������y��e����^���@k��k��K���<+�eQ>��#"����AqxtYN��V{��/טy���~c���b�����˽��,
�s#�*f�g��4ꅏ��J�L\Y� >�oq���8P-f��k2�hٝ����K��:�b.I9.H���Q8*Xb,��j�}1 �]���l��yie�(.�T\c�}G&4Q)�&�S�6ἲ}�t@G@��G�5x��ʾ�ɝ11�O���a1��9��ٽc+FPN��\��������u�
ܺ7}��f?���Tf��*�vB��5��T[�G}+�����R�]�x�Z�ކ���	�)ee��+�Z�R�y5\Ŕ��sVQC+k� �/�|�2�Έv�8��q%�7��3�JÎC*6�B��])��~�j=�N�����@h�
���U��[�����K��qKk�P�w,V�m_�_���Z�<jt��q���^�:� M@�*�Z�1������a7!D7!)ܚ��Fĳ]-W��倧J�x*�ǃԊ"�
�77��f���:[F�x8(������1��5�Ս3�"���)�O� <%���5�>h;���#�av�mE �[^M�͌�ي�k�S�Gق��^�U�b�*��^b�x���R�+AZ��2�$���	�0�Z"��Tc�Bl�1�_5�G�s��W�سz�icjEe�ߞw�Ǧ3���+��0�����:PU���	�5��>�fO���gL�5b���P�,k=@5�^�W�ǰ�/}~u%|g֖���B��/��M��]�{Y����B �K��VϜ�hN�[��WP�qJ���u�}e�V�pD�o��}��U=�����(=�Y�'�S���z�&u�4�8�F��1=:# K������(F��T��ʣD���[13��Ul4��^7(��y톏�cj�)�����V��P�Y�+���I���V��eyK���{=Q5�^��C:�܂�@��j{pz�v�ܶ�]jH��H�#:r��9޼���r�gSڛ��L[�EF�ӬY,Yղ��M��j�ps��ͩ�v�Y6�hл���dj<��&�m�/�o�m�Ei %4�P�����眅^����?,���r��C�J[�t�o�i��/��4j-�௢��������@�9���8>��{�oW���Ne���M	G����v�KӨ�
���~�D�^T���ah�C��F���/Z�gcw��ۻ�ﹳ����5
��Yy�8�S���Ǖ��U���(������i�ݚk��+k�� �,��`���	֩	���($2����t�F�BCf�	�y���)}�ޑ�#���v�R���vO�R+E��^N���X\�
a]5^�ɈL��e�����H�5C�n�5KS\��ςLg�-�mf?"�X��Bf���0���G�nݙ� �fO� 0���^����к��51��UcƩbל`�P��?hv�r��hf8�b��p��@��R�e���yV.�U�V%x��ߞO���>�����9
�߫^Z	H�9�Xn3d{f��&UVS>ʲ���*�[S){���Ol�HS���h{���k���o�E�mm��_�]ԭ�>3������U��JT6�8��Au�W�/����;V9�Wy��,˥�=;�A����.AT�ݦ�g �H��+����.�)�s�"���â��Tÿ /����j�Wb�§�}����g���N#��w[I�}#,׏�8	�;�"LX�S0t��zJ�e_��.Ug����,F�x��Oԧ�<�NYݨ/Wt?K?{p={i�4Cw)z}]|�;�F�q/\��u�|SC��l���Ék|8���J1셴��^��#��UA����ޝ*�3yRb�ׅt5���w벻#U���G+�v�������G��������
a�k���c0O	]��iX�̎?odF���{*_���:Έ�ߣU�ղ�ph�
-�����#o9�����X��o��-��7�b�/>�`?/�}��s�^Ã|�9��ڳ��I�ޡ1���I��H}Ť>�
|例�N۳Y�Vl���5va�<6�/
c�����L�`:����Α#ۻ�k��P����Tk�ynH�S�Pc&.��a�a��0�g��=���c����7ҷi�o�w8}G
/Up]{� �~lK��y}�9y�=�2k
�zL;t��y(Kշ-пO�eN�^�j���3�G/4KM�����!�ggtHeт�SJ�A�x��`�0Q���J��L&ËoT��r�M��Pr�$��j�oe����ڏ�on�J���$!9���w���i�=�VQ����]\�J��]�^��!1�.�]����ĂYe�S=w�%��R�[���W���w�����p`>�?#�BMQ�[�O�bj�b3=~�۫��U�{3Q��{ˇ�x��P��La8%��*���т��z
��G���ճ��kt�~	��xb��~J���j�
u�X
uo�_V?J�"b/��Y�֪�JFIu�������u�s>V.�\'����b²��xQu��Ҹ����mVs�<�f1o��T�j]���mXF��K�<�}�{��B�|o�;�JKa���y���R�n���/6ho�i�9�����ٖ��(���xy����a:��&*��lZ��<r����Qs�빉p!~9��S��ю��a%5NP�=��O����+��`�L�g]��#� ��ر<S|"<~��o�L({�Լ_iz�h�Z�b�
�c-�����H�r���GZSɷ��e���J$��O�^NiB�f4;��W�\�B|[s�Px;���L+�t�$��
Q���]~��JsO@fkv��u`"�*�q�P��3{_�9{N_�b�����&��R�<XU	��xE�җڏR��z 33�6�a(�%��4���El�P�"��+��@��%׭.Ioq���}o{c:a�]Mȷ+f�n`����uc���W�/@����{E�+'wqPkyѸ
�ƟدSc�{O]ϛR�4��)5��9�Thˬ��}	+ �Ҳ��CcQ�6��y�"�⵵i��w#�8�Vá覜��<�*;�Y67=[����G��ᛠR���*P'V�Qgc0�Z��l�iy������nZ�)a7H<V5���X`틑x����d����U����ӥ�.�A�t�ySWӼ�#�D�t�ڔ�Pk� ;��S�m9�k((l�,Ŋ��;2�`Gl׆�OG����}4�3���>�Dud�np/U�G�J�ie��G_���tJٟG�3��X�3���.[N���C�Ho+�I=��N��ۧ�Mc3(E�FAxN�w�śu9r��oDn�r%B/0$R���P� 圧=괠th�`���bۅ�RB�JɁM��伻H���bԵ�E�0�uk'c���B�`q	cqv�3]��p��cOD�p�*���	��_V��ǝ���2V�ª#�*�.�X@��5Ҳ���{��եǓ"�.2nԺ��t���$�_P�۬��EOy��3�]^�MG"��.s8�꼃��i���<޻�pU�|��ܑ'M�O�d:��l��&}q� ��h���	%���o��_V�����Nh�#����Д�{D�ճ��c�-�X�==Xw����o�	���A�(��8���j���u��u�K��r����L�7eYu{a���d��eq�YdEul�c]J�`d�	wY��WM�v�����z,����ӱb���n3W�pۦE�MW�%ٮ4n*7X˻Vk��ua��j�D�6AB�cF�qM��[�-T�d�[,4q+�ѾY_>��-��3s{��Q��4��ל	�#U�6+0+�I�f'��(5	�˽�i"m�ԭ[9]�ۓ^�I��{^!�k U�q��5�z�0���[��Sw�o�Qa�����hg)�@���ۍ�6�,�lU���.��q��h�����g�� �yS����IL\�l����xq�pC2�JJh+\X.�<�8j�@��n_S)<��C�%��s��8�Jn�c-�e ��Fl����gm��k{z۔�U�wm�4~`�YaveѮ���V`.|�d�ڰ6g �>׊v�^n���-m^&�v8���/L4���Qks�M�F��W�S�2O��`ZIk�E^�n΂*T���t{��z��]�YJ$p1B��ǻw\�o#��3��Y$��3V�[Y�V7�wY��i�^��9#<�]>��l���t��.�/:��R5ò�d�D�(Vy�J��#"�l���xQ�m���xF�p*�hwr��8~8E����DV>n��N�%3�%�\��	�[J��MH�|��ܮ]�uF���������-XH{���)7��!];{�����lf�>�.��������ǿ������$EE�)��ͼS�(�nt�ّRm62QEx�����o�s\�TE��˚�r�V��cnl@QQj#b��/<�\ּ'9�]�1b�l[�\#n��sY�k/k��4cx��w:�r�x�^<b�ܮ\����y���snj�m�+���9�;�wk���n[��F�sE�r�μ��+K���T\����DQ���c˕�ܬ#� ����N`��d~:}#�1^��m��eHh������q�/:��78����s��]�gD���?{���;�_�{Z7�_K��o��l/kA{��͒����ow�<�O�G+��_w�חүk��������W�\�_��_J�+��[�wו�W��ݯ�}_}�o�|DD1E�l�����H����^�7~���b��o|�.���DX� Gܦ~-��o����ύ^��no�ǏkF�_ߞy�K��x*��~\5�/����j�髟K�~y�_��W��]��Ҿ����;��[�s��������sޯ/N\Y�dl\k��D`��#"�F�}��n/�W/k|�~y�����_>�U�o�{����^?�v��������W���������6����~v���y�j7������ֹ�ۿ]n��$��-(�8c�}(G�!���;W������~~y��/kA�r�^-��j�~z���U�x�oMx�����|^�ss>��}z��_k�}|���7�r�ޯ?��r��_��^�>y�����������OOJ���>��3��C�>�������>׋��S��忕����~#nWŹ������u�h��~�>vޟ�����jK~�7�����ޟ����~�ڮ\�������|oJ�W.��ΘW��X��Hz:7Q} �ƹ_/<���U������ﷱ���_�߯+�n~/M�^���r������;^-�\�m���׾��-��?}oms��h�_;o-��[�����{�?�
����'s�Ӟ�\�[��ή������V�U����Ϟ�+��_K�����|W�zW���^׵������������������|��W�ί��o�r��^1W��5�{���r�Q8�������
�~���DITX�;{�3=^W�E?���"F��Nb��6������v��F�~}zܯ~��=5������_�K~/�_?}_KF��������}�����_Kž��}�}^?���������j��6������_�+���{ǈ�H�� ��}?X��!n[�_߾ok+�/����^���k�x������o��������^צߏ߿=yz[�s�����z��W�~-ϵ�����xG��>������4E�.*����#�8aE���� }T(W�����?U��w�꽪�ͽw_�om�^*����گ��5������j�=+�ϟ~��ߋso{���kڼ[���=����}�ߝ���żW7�־��`f���fO�5@��yZ¼�j9�ou�o1&m�سB�_SSke�B�_�w��K��۰�Wn��~^P�z�*��t��P݉�������M��p6t�;<�G��{qډ��g3�)R�����[�ut���P�m���5���ξk:0*�uՋ����w�1��m$��}E��$DX��c׮����h�������~<���x�|k�����Z9W�~���~�������{��֮���_��_�?}W��Z6����_�����^��r���o��[�V;���7`��
ZO��>�G���}v�6�W�}��ko��kž�z����k�_����Ϋ����ߗ�Z��������{߾����k��z���[���翯|������hu[�*}}c�B">�:�6��o�r����s��񿗥����W�������߭��[�^�/���+�nk��zW��������^�志���_�^*7���K�~/K���œ�wT�Ï���e���}�1F�����߻��Z�{[�{�~z��ν����6��^-��������/��Q���/��_J�r���_oM������z^��W5��}_�[ڽ*�����<|k&���7;�����>� }�>#�������Ź�����|��.W���z���׵�+������o~yk�/���+���=*�o���7�n\����~��W�����^_��x�s^��W���k�(DE8{^�9\��sݝ��E_!O�ߊ�ޗϟ<����W����zW��W����o�r�����W��U������?�{U������^�*�W�u�\�?{W���żW⿗����m�}� EC�_|Uv�G�/�R�t��xC�k���_���s׾��~?��zWϾ�W���o�}^��{[��^5}w��-��^���������}���^�x�������{o祼U������������@�kտ�ߠA�ܛ����u���_������rܷ�������>��^��{_���7�vſ�ύz�:�^ߍ\��׮��m���KGֿ=y6�����+��[�D[��{���}-*����D�5;g;T�JU4�D!"$DA����͏M����^�zܽ��\���޻z[�ʾ�z�~+�Cz[���k�zWŹ����ץ_˕��{Ο:�-�\�~���׾�j��o��|#�����LM�/����ͮ�#�|Do��~�}z-�W�ϯZ�^/�������_��m�����i���_��|�����h��]������^5�����Q�+���گ��}��߾^��Ҫ�>WN���AR��cĳ�^<����=yI
ݰYoGL���`\�1R��	���RW[��{ڮ;=��~Tn�u�3}w���ԑ�Ơ�a��K2�SaG��R��Gu!��s����l�˺�2�i/nK�:aVۜ�pI*��}�����k��\�����zk��������W���+�/~}���snW��޽W��u����������j��^z{j��|k��~^��_k�}-���;_�k|^��������-�/��]}{��y���^y���*�#}@F���1���`��snnooռT��6��-����V��k|W>/����[{W��ޛ���zEF�׫�痶�o�������{��Qo���y���{}5r��ן���|�쎬�>���n��xtG����1C���������H�>���r�g���<lzM�w��3��5bx���u5\�S:�OO�tHJϾɮ�Ɩ+�
��?A�|�T���CqvyJ�[�R��0�z���� ߮���K@k>�h���΀���>Y��_ /�4=���qcW)~+C�}F��F�mg��>h]���<j|.��3�5V6y�6]q�PD�įe�v�̾�[�W��%cHW���EY�|w��۫��Xx:����>A�b���W_IL�r%�8Y��3�-��jyh����f=�J�`����z�=�ҹ>�]3V��U�i�d�R�N^s�y��z���>˷]�\��0���䈚V��t��"�.@YP׻�Z��3u]Xކ���)�R:"C~�W�b�V�ӑ�������#�Ȁ����(�S�H�3�3������kg;IN��y�ai����pCx�|�ҋf��O2��h�����+��p��!��U�poV>�X[�kH��!���+c���[I�V��;�E#�:󦒠#%�X�/
<뺩�Yڥ�ヰ�bo��t*I�W,`VO��*�>�b���u���������uo[h{�(<�|Bi
�L�A^Й�7G�e�.=� �k�|ϽwC�/+J-v����,��,^�}u}OD-��O���;8������}wD8W��Cܡ�F�U��*�w�n͓^p*�\�>��*��c��:-��Mx�İ��e�6�nr��n�X�����v��4F��+�_M�ώ�QG��*��&�U�k�<�/��|g����� �?"�=c��
9�����'�e^�~�|��[X���
O��\��i��L+qR��b��~\�W)�z*��m�<}����a�eS��+�jǅ<��S�� ��W��AU)���}�Lb����<�6�^���&دw���V�t�%xJ�ja�Pg
;��Z����?-��}5��5t٠���G�
��WF~xWs�g�__�8�=�ۯ^:�Ŭ������Xf������D=�lw~��7��S�m�4����p0��]�3��Ak϶��ද'��鼥�ow_� ���l�^2^Q����؄T��Ǖ�Q��X���g]�ŭ3�o���n9K�t��؉�F���/_ ��8zc�WN�V�w6�K�b���l;�o]5������L�Ђu�۬�1-U�n�� ����S0+ύ�D����j�����n��R�(1��r���'N�ݲ�pX;F�˼3r�rR�/[����C���^��󪆷y`#�W�
��yk7S�x:5U�7P�����PjB
r����j�Ț��h�Y��������fi�ZU����U�B�Dam���~5-��PFNUl�i�V_����%;)s>�>�wcj��wh��igp�y~��M���
Nyی,�d������]�Wx�]k����~�,�ue�X�{ �h9Qxvϲ����v-Ö��ӱ�vސ���)��' `�����f�g��b��zm�Ŝ��3�gr�z�୾�����DϚ6>�ݡP�6|\�>��YEE���É�Ǐ	Tp*��U�﷢ݩ�M� �g�������Ll:�<����A��PJeI�N�����+�Q Tw}��J<xeL��}���ݐS�bz��~s�x2��Xuγ_�U�ⵯP��@S�e�|�8�{ރ+s�˼��1��#��|�����8=&�Ǿ�bަOZ��w���}�uU�h�!	�c�!ZZ����om�}*&�A{�o�dH�o
X��w��V�fkW�`������Ҕ�;K�.�;a�x�ff����R�b�� ��g]־��L�pX�q������6U;��x�-��Z���S��
b�o�n�.��~��(�	h>�=�n���ĳ]>�^Üp�*���Pxn��`F�춵�3m�h�!�^%Z��9��_�h'�0ud�=��7K3'ҮՇV{�O��v,�uLx��S��:��:pW�36X,�B��,k�3��ق��2ϖ�^�n�dc�z��NZV�q�5�#�|6�6#ŋd)�!�pK>�0����:��a�7�z���s)��� �y��`�K1�Q��[�}�����ٖ��^]�����`��JS�D�Jg6S���A~WYBE�:��v��=��B��_V�����
�Y����l�*�s^ڄ��w���p��Ru'���x��8`�yJ~�����%�]d��OM�PV�T�]P�.v6i�G��<�m�n�C.�C�8ǯ��S���E]���.��ip����'~�)=Mt8e�y�u����=�n����C>9'K��d�7��ڟ����0:���^y�״'���w��R���	��ܯ��s�o
Ѹ���*C~s�Dt���3�@�81�1Kgx-�qx�����w	�n���Iq㮡M��*AQa�{η:�|�6�D�vw��#�{0a��F�_1�b��CQS�ȧ�Cďe��/���8<��楙D��SwA�)��Gb�3�KI��=W}�*�ݴ�ѭ�/�j-k�W-]�a�^=��AO��:��ڥ���L�U��6�ǯѐ��='��q�����')9��~����3p�ِ-�V����j�w��Ń���Y���w�WG��[���9پ���tk��=$������*��,?��T����2��n�1LnMin��o���7T��h�Vqy{�/���T/径��{<���Ԋѱ¼���S����Ku�8t]��@N�f�6p KR�P��A&3ز����kș�� ��W��}����~:�+QC��޸ �p��p�hz�_RXnja�Ǎz.zW5�{�O�Q�L�bgG��X���ﴫ���>3�خ���?Q���#kR�����+@Buc�~X�WY�Cw�3�i�7T�/O(V9�s
\hض�\�E�mdS�Ǫ�(5�� 7�FEg��޷0�]Vb�/�����k��,xT���V�;x���Ɋ��K{�s�za��:,�P]��g�j�l�tl�=
%~3��������KF���y�Ue7��Hwp�w�l<h��-���tW�`��P딟����;�n��K��֒08��Vo;�����1���J�3	e���+i���W+�N��#��wP�Q�}��;��/29��36�0�JKZ�q'�ZG����O.�s�8��{_��ݝ���k�C��pz6��>TCw*��Ժ�J`�׽�pJT�gv�yV���_yM
�s�Ǯ�>��f	u�`V�c����t�`+jb���d'��]\�s����^��ks~���R��0���r�TV��O��s�����}�O�ot�L^`kZ��)�=�gƘ����1�e����0�k%��A1~e8ͼwx���30+'�m��a�tg?�9��I�ݴ+�;ڞ�&[Y��u�<qc4S�Զ_����qV�BE�~�1>�>8����F0E�b �i��<��P�\�ͬ`�QY앪�k�؇���,�� ��3�"��M��#^�S����5�/��ZCX��;��b�7eI;�LĈH�5��*X�_l� mCy`��L���?y�g��ǎ��k+�/�$��Q�у�xz�|ʭ�\�=2���x�K����~Ed���:�۞;Z:�2ۛԵh�����e�Yk�J.��� ��hx��R>9�x{h{�^�~�{H��fΖ�^m����M�W�f-pv�Dn:}\�A����M�m�TyF��wÊ:�q�V���V�4k��z���IO/�RU�i������>	�e:�p�n�����j����>o�76p��Or=}\�I�J�]Y�*�.�|ĝ,��&oK��#վ��h\/��KV<)��[�ד�^�T�s��@F�xr�xkq^y���c&����%u�FME`����!�0𿅅e�/
/�\�O���	��Ww���k֘��B�����߻�U�s`���CC��׳�.v� �=������k^�@p�@��n�#(����Qq�	�aw�D�+Bg��AkϦ-�s�eq��4v�/����g 4l�W���
b6����I��$�
g�*�^��!����9 8m�E\dϏ�4k;2�b��˕;G�1�/����F�AwM�Ʈ��k�{Wu���R�zh�i0t}�KW�����G�/��!C"nw�!9zsi��ʻ#2j�=�ϟyW�c�u?C9k���۫ U��3�#h4oV�ř�yd���z��q�^�+��9@�U�yaЫ�W���O�{5�4e-�J��Aqxv����;��W>��֍�E|gr���0W��2*!�f�x�lj��މ��=�aih.eGG���o�Lt[��R�gp#|��9�1�`����A������A]C��N��d�d��zĉ:�:E�k|�,>K���Kpj�O#��Z���M���[xEcq�d�`�o�G�5k=Ǧ��-�K�Bޭ��r���<�@�pu�ɛm�w�8�V���������_���ɽ��u$0�#HgC��)����R�5�lvt�\���seZ_X=1�aY�=����2��S�6��"�UD�c7�E�<xee5�z��`������������9�^���j��W�?k5�. *ɛt��[��묓����@#hV��������ҭX�]<u����t�J�S�u��*���)�q
g�(ۨ"�jCD>Y����bY����^r�S�\<0���}�.��z��1��N&�s�����}*���G���a ���Y宽gVc?K�=ܫ��1o�����b��@'J�0��ͤ,P�9�s*+}Xj}^H��+�4,�mrv{λs���E��4����Õ/y�~b�A�z�������¸J��p)����Fa�E���Γp��ɫ>���H�Y�iL��hWS�I�ձ�ٗ���;y��T��hlV��K���gA�ǫƬVq�y۰vߠ��Bo�U��=u�
�X�>���_�p�M����c�.�xrC8e����4(�Ll�Yk }�kS��,%����	��я�p'+��v�st��4 �s�^U�.�u�+U�d}{�	��U�Du�o�1���,v�U��)�R��&Bآ<N]a7C��8> ��Z���'˴�N�x�Uѡio��Ʈ8Ϟ|���T<���^�ˮ%F�q��R�Wba��V��-��6�2�6�-���V$��\
�XiF�Y���4-Fs��йE�R�|��o\�^�"SG}d]�42����e�mc�������"<C9��6.ҶC!;z�0E+���/�,�4)�fu��T����}y���u�|��ګm�J����(K�d��Ӣ�ލ�w����Q��ߤȕ�����30���T<���`�ze!���}�
��1{��w-�t�"�g++����V�x~����Z�HkS�mث�te�]��K���A�j�O����^�GR�]o����ZUEzS"@��xa�77�.)n���Ӑ���&[�=Ë�NN�yn���[��a����]49�ݶ��#�Jg���n�N�{C4Ŷ���Όh8��+��,E��)��[���I⺰0-��\��c���V��X��,j�n�VS� ]˗�>G��Vڷ ��1���W��!f�Z���+���j� ��*��'�ze�V-�ee7�W�S�/\����!��\U��hy�ɸ��Z,�U�}ᩥ�\�&+pث�+F ñ�i#�G^1N��R�+:�`v��(����+���/0�Xc㯲�$h�����ʧ�m4TЎ��`�q�t_nB��h*6n�&,��U���m�t��$䛆����v9G�H����0T�)㻗�X�����;9D�^��t����h_jӖ2FV�\�k��K�ҍDH�ɫ&�r����U���ޫ��WEUɬ,�X��Q��&�0Ǜ��n���
|���Gϙ P�n�@���U�=W�w9���8���4�^ "�c1R7���1�8Vb|ܖ��I��7k_��۾6+�S�*�R6!E�F����7�V�O���qS�j��-Y̡��Fb���-��>��3�]9pb�m	��]R7с�@Z|��5�w����楐)�@;�+��Y��q��8�O��e�v����t7�9�t�h>O��!�����Á��[8��P�Z7pEW�IeT{ʙ�b�j�����������cF�P���r��.4)ŝ����Y��
��N����_#f_:���)zm�#�BS)��u:��uڤx�Eչ;��_s����[�޼A\�6YuvoN�/c"WKճ���(_]�u�0i�W��AӔ�{�i6OTA��^���2v%*�������vW�Aͷ�1��X/�HA�M�g@��09�z���E�����6 �`����@�y�Z]�TR�.� ��%yK��
5�Vn�q�.jZ���K�988�쐏�Up,[E�Wws](�6�\���6-�wv�u�oկ�s����Ʈ��G(�Wwr�sF9j�,wv�,s�]ss�u+s��S��7.��7K�-�\�G�^3���lG(܍&c�ۡN�\�y�kɹ܎](��(�wQΔh�-˛���K�E�\��f�󻻢�Ź�U,���fK���̜݉F���Lk�M�Rf��I�껻�a.[�A��cO;��LW��n�⁻�p�%�̺��$"���u�B@�yג]� �s�����d��\�O��vJ��\"�����7:���O���pCT�&[b^�0\�خݫx��%��0gv�3^���%�y�̐ib��1���|K��y�R{p���|)���>>�p�8��,]o��-*��%�}���Rz���ى2��1�zr=X=/�7�g���^�ƪ�^�/�#Uה�V@�o,�����[[1-�rϔ�����AyLh�X�7�����U�PEY %,��mO��=��//7))w�ł��9�"���s�y�l&%׼����}�n�����T+k=6�4��yuL@r/��s�PS�;��o7j�>��я�K$��Y��f��q�M̫^~˖��ʕpf���i�-���,�{f��p���G�[�g�d���m`5��0|<��@�cʬ��?a\�u.���m�aНs-� !{�4nhT��2�D�E�Vn<>���Dx����ϧ����Q&�{2��4b3��¼��.���ۤԉ'BtW�tE
�du���f�X��Q+���c=�);�]೑ԭ]�ϫ}�s��F;�9��!]t1e-;U,f̖h011	�0��X�����~g�����h��G<���|QnK����Kv�n��ݥ،푻Э[����Djm+MZ9q��x�\�{�f|pb繪1D��%�@�����ݝI1|�ͤ�W��bB���/��2̵�Y�=�sjK�r�45�6�d���C��rs̑d��5��G�}��t7%B���/��x�L����ut͢�E��d�I�^	�V]=��ʑo�oOqM���3ݜ�S�� <2,|.+�������C<��xJ��O*���(���R�H)���Nur��@�}^h���΀����He_ /������2���ANWcrn���Son�]�[�{U�S��Z1/N}&,F��:rVdU��8�����xf$=AuJ���rfߪwo�jU</!���=�:<�"vT	ۉw�Lu���0�[�!��"�B׎��&� 
g�i�P��)���1��CU��4�!= J��P@j���u�=����f���q�@�}q)9��
+��z���]�Ǭ�)B* �v�}>����QMѸ\��_W�� ���F2�W1�����q��Lj�~1�,��`�h�I��DR�)mj�\�sL������+y�4��0��������ó���>��'�xyt�a��`^�7Nb)�d¸�1-�>�o��`�B�-v���xy}�הU���iæp��1�������Od��w)v��~:�Μ��H>��q� M�]�w"n�n9���F�]ڊ��k�=�w�ht{wS[TD�Ɨ-����E��h�*���q����#[���	�X狣���jgQ�q<�mm�8K���6V��Dk�E�8:���t8#�ŏ��j�-��*"̣�N���q��(��&�����z�����6u�!�Lf�ૅ/�W��OL���L��E*u lL���|������b�����	
�Dlej3hve<���>�*���T*
��b���~B����5��c
C��E�x*]�GmUﲹ��-΋CFCWS�v�bP�wL�ۼ���T�)y��c)x<�����lf�<�׀��k��$8�Un�u�lu����8w��c\�l�۷P	����*�=�^(mw���+h�.=���k�K%֪��Z3�s�וv��Ȳ�7G�P�����|_�K�=��+lװ�k�k"+�]�¹��9k:/�g]Gٰ������$Ӹk�(fW%}ǖNX�{�9�ɒ{ެ�#���.9�B�#Ӎ1���O��u�f�X���B2;��-��C-�I�r��»�7'o<�D�R�tV�m���4ȨJxC��7���VP�"��[n�tp,���'�n��aF�)ʶ<ݺwj�ga㌪���r��u����v�&[&�����=:�KumB2��=��_G�G�}��M����lW-�w� u�k>���7��Y�5��7[O(E߯6�$-�^=���(.5�q��׽Y�1�z�>��[D�i�O}��DQt�n,z�U�&���-�??\?d�m谖����eG�j���W�Z�o�"W��w����r��W�_[���L�l+��u}����Z��s��l�{��n����+3F6�f�W�n����p��~�Y֞��.r�+��}��O.��^���~��G'k�1P�l�6p{D)�v�X�wG�J'���;�ߪ"�=V��'��+�+�9�q��Æ%���Fױ1�>�V:�?��xV�^�a�N��]�X���	��.MN,^ʵ��	w쇶�\�Bn�_({?/l���x���-�R:�w���B7NVW�G�X~nq�WF��8-F�9����œuv���u����x2�4>�]<���Ll=���.?s{9VOV�h���)Q��ĝi���B�F�A��re���6I�
�HW���ѻ�g�{��,�Gg�����yI��avzGt�݈��pxN�cWnţ.{YV鼫��J�-<�Uε��ﾪ�����+݇ޯ`���'�Pcҝxڊ�a����M�����=���\؊��k�Ԯ���Ib�Լ���?o��^^�9yr���;�L}}����B_r��������G�jb�x�P�K�s*�O�:����e�`�o�
�P�Q��ۛ�};j����G�Y�6�ԑ�>D�V��U�:���߆����2��ڜ��zy���<�^����T��k���2��4^�G��LJ���nNA�ף*(��~��%�n6;7��'�\;�^�mS�b~��iv�Ɯ
�-BTʅ��V%��u�>�P�٢��|��i=y[#9>~���*�He|�&<�Y.}AyZ��+�[^��l�)�u�J�Q�s�O��.���s}����+�Y�Q�*���kY����d�c�!�|0yz��Ɋo.�(�w�R��]�����q�'���t�چ���N8���fR���v�ĝ�7���Y���=��8\�E'͸7Vp���j埽.]}C$�e��GF4G�յxMY;TA|���q8�]�|��[�Mm\T]4����9՚U\���bn�	�V�п���U��^���ݬJN�-�oZ�4�D�=���by����Y���v�@g��k�	]^K�[R��eƧq*��;�g�2C��#zV�|^}�ڱpt�<�a^�g)���LƸ�[-�7�Vɩ�{P��'�V�Of�� nyG��X�O��Pe(�ecs�P]���E���_�:Q[�r���޶i�)�U���oᏙ�'���?b���4���0���$N؊�̝�]�,�^����Ebz�j��^D$���9X�ה��x�צD=�q+ؚ�����w���ot��{,���uqI�Ҕ��������
�˗Tr�����O���k�7ܯ��%p׶�u��fx=*}�-���0LRo���eeo��%'���>[V��!�}��y��4)Iյ��t�m�ī�fz����P�i�rzt=���ѯy�C^u���L�엹^�'(*H:��)ͫ}K2�
�e�^sM���<L�v�B�`�J�G4��mzԃ�	�s����<��ǽ������r�.Y��#+�xNNb+�`0))��+�V�9f�жr��'T�
Oӫ�<!�?��G��~�c�~3�^�P��3�����6��jtk�f�l�z���v{���A��<
z��'������'J�|_vuG�3�X��lX�㛾9�8��Ls�Ws~"��	\Ϸ��N�G�4�ٔ�����/r��QU����N��e��2�B1��Y����{v)n9��ڋ�1�A){g4�h+2��G���z�j�z
O�R�W��n�+��v�r.\u*N�v�?�ۻ����nN���	�P��O�Xk<T�Ɍ��ܶ���1���vOV:��S��W;�C�y*�V���{|X��\Φ��y�Doo��ݥ1�RP��x�2�g-����6B�!�'�2� ��V�w��˖�~�t���%���Q��n�e��G����}-�eT����d�j�a��j5�SYUv	����~D%�D���cձo\���^�T�ղK��#v��E�u���LŽ�[�2Sj����������uun:���6���N�N��f����8�G޴��0J%���l���e>J����_c�T4��r�����R�k�k�ulCaB��}{π$�&�)�k	��x]�\?U}�}_W�Ι(�PO�����1nѯ�˯��ˍt��]<�1��U�s��hI�WV��:1:.S�{Ӽ��Pt���k�K�M���m���L�`���~!M�J��]NO�b�>��Z�^�}4f ��]ч�K���ޯbWg,�����#Ӌ�/fS���v���xW'B�)xj�~�9�y۾�OʄB����������4���(xu㤝�Wy:��{۳Ij	^����A�* �/�x��3�{�:�v����ƺ>�;�;6�?�f���^'iޜ	B���Ԙh(�ۥ��'�������3y=G ����/Χ����W�ex�mW��9]wKW9�I/���1�+��G[�2��\���է?U����x6�P�?@���/�a/��������?\ч܀ݧ޹k���Y�ț�I���^~вmĤ�gq���m�����JKsT�;L�{�,�j��|��+�y<�w�Ć0��k�;o�N���;yX5m��M�Ke;r�Msn��w�Y��,F+w�ɨ�9FU��u�ȹ��^���[��y�)�Q��������K�y�OOM��_����:����+h�i�3Oy�z�|i?nM�6O%Ml�)SŠ=�����9�~�U������a��J%��ٯ������,\v�����zX��}]�Z���,��tD�5hw�W�΋���jǭ�|�{ɷ����E������*��&a�k��ϟ��^B���v61��J��y.��,[�r�R���ߠ=Z��Oӓ_7��@���z��}2Ǐ�5$�1�g����	8i,Z�KϩTά/��c�}��~��Ksv�*5�݊��߽~������9�ƒ{���m1�>�;|-Vt�y3w1E��@c���lj��W�ؕÝK*�q�!{h��;㘅��'�f�뛲o�W=?�v�{�=O�SL,��*צ�Χ��ϗѻ�}l�<�;}^�}�Sӣ\{��竳��>[]��[PuE�#�Q�����
���<.�EK�x?8�;k���}ңʧ��M���d���q���<��3Q�1,�4a��PN�^`m��o;�Y�P��3n�kb��Y���u����*U�c=Cf7��6�q�gL�gJ��b[�i��L����}}�x��T���c�;{_Y��)o�[x��8�շc�eDZaؿMց4�#�՚eC���ʴ���IG{*�oT|�Q���H� �|��,q�<9��KA��+�ڵ+��ۇC�k:�=J_��O;����ɖ:�=����G��^�*�E*edj`�K$��on�-��	��PD�ȇp~�u��������7
��	�R�T5T�yQ�v�n����%⍳^wEHZ�66~�N�@M�e��'�f�5��|�yP۳^X�^�;z�n��H����U�l�>bg\k��p��F�~j�5;r���"��E3\8���oRӼ��I���+K��B�!�'�"��DѢ���znTc��T��!�߽~�F?3�Ex���󱋨<n��Za�è����nV�~�驗�.�Voeŵ�~F�$�R�1����ӴƟ��.�M�V��E�q��n�sc�}/9�֏:Va���RԡZ��VӒ��+q��-�C���ȏ\`����)�gfs9+��	��D�n�l��Z�b��Ҥ֤�fF�kK��)�����s^��^��y]�[2��w��*��%����)����3��b�d��c�xq)P�F���r���(�b;�uѥ�άY]u�]1��VF�P�VR�9!p��X���D���Z�mV���:���:u���#{�vW��p��|ֳe�U��o/�!pe�|spr�;�s�pM��{N���')��oBmw�� �_)@��`�7[�kz䔔u�Z+9���B�편vVV�9A�VzΫaG�eY�ja�����h}��$HW�.]��֠�mkCz�_�E�X9�23��������gT�i��E\��&^G���(���,Ӯ2oK�va'��75�_zs�R����b�)n
�TY�WJ���2���N�!e��v��ϣ=æ4zU��n���cN�̈́2k�Y��[�^M���zwL�Y�e�/c>��Y�W�=���À�p�F�QΥ�s�EAkWh����BP�N���
���f�Ȋ�č�+�6�.P�î��G�G�v�:$N���(�Ӹ!R���$V�՘���(8:�o��=6�y��=�Ͳ9e�ґ,�K��u�yG�-��˛�C����#��J��-�[w��;s#����WY����;�$��apuu�:�}W�л�ە�Vr,�/��ƒ�������}��[2��n��)�u��o4[����e�����P
����wN�yy�2����;������ۙY�u�~~S������D���
�4�|JrS��&g=�C�d�P}��o�՚xb�`gw�x��E*���U�N�̖)��;ot��� �<"�@4w��ẍ��n�&�M݄,�֡M]�Cl�,�h
'�d&C�Ee �ki�ja�(Uݴ�At��c�u�����e�w�{� �ջ���Ӆ�[��'lE�ѩ�|�����t��v�KJ���.�[1MY���@����h��۬q��V��(����L��Z��׽�����:�	�P���Ub�}���Emn�f�8L&u頫�qcJi���� �1�YAѵx�-v�M�ˀվ�M|Z���cI��?X������-�n[���Vԡd5�����f���o�,�	�����K �Ӣҹ��Qm�ζ-L}ς�9m�
��b�!l�sM��B�x� ��G�.�&±Z�]����T%T7k��)���d�m���+�2b���%۝7�.��tW��&*�\h�Wa�Υf�=��{%��j�G:֋ƅ����G9 v�;٤;��|$�8ȻK ��$Ð]
勳rN�a��~*+���M�x���F}��?'�n�s��S��(H1�9)��(k��f"���NW\���ם監�s�D��uu�
�N�N\�����ws��7u��AEί:����b�x<���R��'w!���3�eΛ���]x�N;st/<nDM(�\���(��w`��Ƌ����]ܞ;x�㻮�wnQ�ѝ��w.��� f�"�7)O;ǖ����d�Irwr�WA������3�e�m�y���h�7g8�+�s	�;��7ws�»�����)��]&�(MЌ�䐅ݮE��;ݸwsp]v�;L��2�ww.wg\�됎hwB��K��\�7uu�v�S������%�mn��wR'�$�����<��՟ywg�hnd�Ġ���dA��.���YQ���c�����.���}�U_WD��6g�����U��ڥ<���^�ix^�S>X����R��oS��| �"��nt�:B>�qKbcҌ�z�]�����O�bW=�x��ш�Kg��]e��J��~�9k�
�ӆ�yq���k��߼��Įx﫦�-gi���z.��z����=��dI��s�*3ӻ2������z=Y
3ҤO���B^�aL�Y^<�h��Dt�{ݯ��2��Lz&v�E�T���-l$��70��{	\�4��ZL��=�h�joI{�V��JGN��y�t��s7�Q��=�{}ΐ��^^fn-��V�ހ��W$�9>�H���#ڤ�+�����������Ï�k���>�V3�� R����"W�{���cS��ۍP�Y�Ѧ2!�j�e�:�v���L��s��pV�{�F�ۻ
��΢N�h����J,��b���io ��Z9F#N��k���x ��[�gT$^QX9�G*Vq��p��*Z�.�u�H��7����Ez��t�R�j�K�)ث�~�J��ٲ:�l�*f�.e;J׮���F�����`�-�c�՞�3��7�4n�u�Wkl �t��V𤤃�v_G?D}�DDC��I�����u��z�&*���fO�EZ�*��Oվ]�Խ<��-G}s��-���k��{��)W�}c��<��\¾��'�z֡���ux:���)^�2��ȟ��KP��b���1����3��)4��ج�;�x���=� 4�uL�A<�U��^u�7�W��%��S�[[܆�>A�o+wgݔkV���%:���P��#�{��\[���rd���k��^�y|9{�,JQ��eF�1��iO�7{5�қcv0�z�Gv��:���W�ok�v��Z�ڎ��v�ǖ����}�����Ox\�q6�L���\�|w�{��>ĮQ�ے�]�G���z��S� ��c������9n�J��~o�Z��T��g&�R���uU����%�c�C[�{�nc&*�kъ)7r��ח�)'E޽z�T�B��ۥ��O�7�BvF+�*���6�����&��;����{�&*�"糗�#���љ�U������v�t�U����#��7U�4Q@,
kw9�gQ�Ճ}��JyD�B!jk�����r��MM���"]��ʻ�6���m<�o�9�;3:k(���R�nV),�v>�/7)�_��������c�	��|�gn�羷��.۫�f��q��d�Tn\+���D�u3�8D^1��{\gM,��{���^8���%p�2�BL�N.&�LRwa��{�W���O�cV�=�'����올ͣ��oBQ�U��y(�@R◨�������xS��j���z��D�����B+�[�u˂Z�?	�OH���_��[*gk���Kuiβ�ӽ�*�M��Lf&2Rў����kӺ�'N�{i¿���y�T�� ϖ9������dg�kt�g_c���2ש��q��e��,�:٪�T=�]�B��ڥ��ci�Ӵ����=�w���Ӏ��pםq�kִ�^��훵��G4w#��r ��<��L]G����ś���:�Qg�˶:�<�l^KlM���v>D$�Rū�{_P��uc��m)����ү.���V1	��jX��X�I�H���2�jJ�|QE����C��s�U�_���{w��l0OW��絑����X�Y�KҤ��f�_�fˈ-⋦d�'v��N)ܷ�h���~������m�S���I�G��xovǳ�E�ڡs�Z����{���o�}t�{�(��oP��{��y������,�k�ؕÝK9qͪ!{O�v�DX�珹#6Sl_�e���nU98oo���t>��?/^v�=p���U���7h�[s�]�a��҄r��#��Ν��Vv._s����ٝ]�vΙ����y��M����S:�0�);���_E�������F'��ߨ�l�
���Γ���Mmxz{qR��5���*�&xoǺmQ޸���o�S_��w~��<��,��{�*�����}��=��fs>�K�B4.��Z�E�1ZԿJ�O�9��YW�j0j�-ţ�D��J��	�SwU�_`2�R)[�3"�6�N�v*4��5�	��4O,'����}{�if{=�{"^���s�~ܝ��5.6�O"�3BWM��e���o]Z��M�ʞR�6�����$"�������?
�����|XTL}�[�Ȳ�VT�z(,XOT@W5��"�9i�}m �9�=���2���6gz+E�4	��Cz�u�[8��(*Mu:���C�Z�J�I5-��M�|^,���m����.�������'kYE�Tf��������#�H���7W�b�x�F,�\zB�13�k�h�>��a7,G���ւ����y��P)��U�w�g�����N~�
b4�1	�s�-��`{�]�i���W�6|�w;�n�����3����w����3�ǥ��H�SC��d防p��t�]h����xjr;�<�e�t����mR�0����	>��尒{�w��+��Rr�>^(mw���hײ��Ư�����.�1��Mj�^���R�UIK$���j�y��������y܈#sk=Qo���n 趮3[�lnJҊ��u��<Z~�:p����]��ף��y+��f�AF�M�̛�5��B�S�qU����J��b3Y[7	0�o2dKv�{�b�)ߒq��ن��t��{WpU��W��97�=��ݵ���;��ڨx|j9~ʵy�KV�*_�SLXy�L:�T/��Z�������ۖ��4���{���q�2���hO|��{z��8��j7�d�*�	¹u�E���.�-Ox���t��w`)%u)t�M
�i�xӒ���%�b�Y��4����tJ5�m=�WW0�%�sׯ.�h�V��pZ)M13{XsOkN�Ⱥu�}���W��I{��wя�ּ�����-�	0��g�:S���9��N��]^o���qk��o[�Ɋt�6���%_^��Ny�U|�2�'RA�]���طZ�WqO'^�C��%[�������5=�U�������W�r��紳��"j�.�+���}SP�3���Cx2V�S9]����wf�+�R�W�<�=����{͚�9U2��mU������o�Y���o?s��f�O@k9��%zm�|�y?E�\��O�#�ʺ��@.������@��Q�^<��-�|��5D���њ�G���Iy�ϝ�8O��{]����2��͸�=z�Lۅs��`���^��h$�
�<�{�.�}������򃲝F�qǊ��ߦ��O�Y9��j�=~Y&�����s#8g�M�RŵK�{_RϧP��V��>~��f1���zݗ�v�罝�J9����=~UK{��W��s�Qd�.����.݀!�V�r���K皊�WT�e6���ix�|���q���A����cT�z��f���{�ea�i����0z��y1�n�}YZ���Q��§L��N��tdr�gӺ��U_}UV�/$��b��9��P�Y^��8�E�G�ʌ�Z��M<�#���F�;9!hݣ�`��Hz�����q�eX�D�Ʌ���/W��G�y��¡���nm��Yr��
�e�ẽo�ZF�\J��VuTYZԨ�ȷ7{��:����w{����}���s��ۮ������nק��(⮽Nԅa�3Rn�"��RU�^O}C��m谖�	CP��dс�f���BSSng�.U�}�{����=&�����0��d�*��i(�Rp2�_�ot�nA��p��p�A�5���R��.{^�r�� �R/�r�~/<�샢hz��[j�2��o���މ/���M�Z�6�
h��B} eȓ���{2[�^��;\|iQ�t�]�ubs��;ِt�r�l��yd��o�y ��vr��u��oyVq>���6�>Kگ�D��J��.�_�"��pի#�j���^�L�Y����ͫF��|�����,+볉��up����B�r�|;^7Pd��/���`欰��u�J�(Hxb�<9�W!�!�������X��N��)��ׁB����>�.�=�O��o'��}!α2�k��n�$�d҇��)9ղ��}0��NI罥����Ec#���V��-8�nq�u^v	\�y�qTg�)���D�ベ�,�b`�ؠǥ��ٵ�s%I�����6o�.�=ݑ�x�������|�㠷�Ib�Խ�O�}3�)����ڜwh#���y��7}��cT@����>�*�Z�~���.��LyEaՌZ�v��e���ey{H�L��au���ܕ�}�\
-Z��l���|!L�^�XaKe����)S�կV��ݬbUz4�����8�
e�;7���^��<�n���<�w�o�&�)��F��n1�^�/7r��歿q��B�q�Gg2;�~{ݯz#ދ}�;�޹tH�do�+��t�.�zW�|:���bלkh�����Ϝo~S;);t|I�z�K7�t�p��Y�Fw����S�V�{6�^s/{8WN[���j�����D��L���M�:��	��Dkx�'���c*M(K����}*L�[8�Q�Pfҋ3��t\���?rJ��n��oy�孽t�Tq��l��3�����'gH[@뛓��`c��n��G�}�E\���N߲Ƀ�R�)���b��'���u�iu=����\e7�అn1J�N��z�^�M�2�����{���g帷��&�z$��$��
�s���y�g��a�q����Wڜ*�x"i!CT0y��#R�\)��k{nwv�Ɩ��]��g��n4�=�=\�҆v�V�uܖˑBi�X`A�M;���N����y�Tڙ��ϟ�����~��ꞃ����Dw�=��)�)��q�=�:�D��j�<sx�3�~ŀ�bs���]���"r��n�ߦ*Y�%˯3+j�犫.��D��#�r͈3�����q�ޯ?1���P�;����ּ��<�o��Y�ȿ{.-�?#Ag�Y���\����I�ugh3�ӵ�^����'��r�������k�o��3�.���}���^�|��K�����ӷ�gy�����r���ĮvHh[8�CŰ޾R�$�w�$]�a�sw�����|l�.�Pk�����̪X�e^���K��L�ˣ��mvq[^�R�BNn��+��x�	��]�ioWb���K����N'dgw@ɗ�Mj�fd�H���w2�v��]����j󷑑k������L�z�g��P���y�)�JT���'�_)Í$��^�O|5�D�д�Ub/0ш+G��� I��W�ϧ!��е�/U��^u:�l�M�r,�QkR�^*ɕU�Q��:�᳃��Ǎ/���t�{ݿ>ٜ(�ֵ�Ϳw���$�}��Sߏ�����'��sS�ڟQ3�OtT����Q>�E�U�J�wZ��/'���2~n��A-�0�|ʇ��vpyT�Kߥ�Z��+̌���h�ޞ�E�h�{9���d�N���t��-���J�5i˘ʹ`��c��8���\�j��a]���ƽ��%U�JQ��Y"5
�x8A��i���3�-���ț�$���2v�h��r����#uS9��Z�:+�ݢ���Ag�[�s�O�w��P����K��M5/{��0�/W�Wo����Z%zmX��x�DX�\��T����h���d�A�)qYtU!p�N�s���f��#�Եp53n�SIX����T.�ZN�]t}y:�8m���}6�J�
�U�vͷR0^�z��k;��h����-���U���tt�0t58�yÇQ�(�xk��3;:5}v�bу^󖘋*oE>|�k�/��ä�IVi��a�RjNe>4��$v�m��p�uN�8��i��ޫ�֞�ڵhaWRFpR�X;���x�`o�ǻ�$�X`�q�J�o���x�fqpCQ=����Y��6�5��}o���j�㶵�k���VR�u��Q�L9�K�L�&���t�ĎսG�ԥY�$�Du7�5�b�]G�S͙�%7N#]�8��9���Sa�s��E�����N����a��7��Ú.��Lu���oE��U s���]�c��N���*�*Ŏ��@w/vH�#G�/��QQ �Yx�G�N�Dxb�n��v6�� �O����fPJ�J�ݍ`�%���*v�3^�;y��\ֺ\��L��C������1숏�:�S�mۏ�o���_܏[ϫ�r�� i������a=�GF�%!إb�D��<q�%��]��y���ĄP�E��]kW8u��}��{y�yg
q��i\ӱ��7P�{M��^�� 9E��ܷ�fY��0;��<62�H�ٹ�M�{��=ɚ�A��u�*�(��_K6�ɷ���<B:ժU�޾w`�(6��Oڴ��DB�t��ۮ��[��1�gR�"�cz��)_g;��r�[5,m�sM.XK:�m\/�!��+F�[}�eH p�{Nrn:-���{��&�o=��;^��L�S��(�u�6c�CX�7%WSE���;�\.�'��2jS+�Ҷ]X�W҉�F�8O�o���t8��*�^�,��PW�f�ɫZ�}�,]��Us K#6�9``�<2ȏ�c4�)]T�'���v(E���%��� BP���^VVF��f|5���G��i3�Ʒ����}�w��>A�<��ϥ�%�c��AP��4z�Bu�[Dqr��
��vRɏ�eԕ�0y|uţJ4q���r뵌��e���}�p�֮��iී�%@{�4^������#�q(��a�=�ۋ]`zIB��T�Ѡ���M	ֶ��T�:�L~��i�_+���;�G:�]���ʴ5��h�)�����VU�eJסD��$��%��ow�ö��뻘	��=�����w�')�(�`�`���$TԮm���SVŜf�80�Ơ#��$���3��o���S!�#�u��Ed��VOgg�^��~ӄ�*�j�1�P{��`si���Bma��єƁW��wU�޵V�F[nk�݉(�sw為q:Z�ml��,��4�jVapWi?��dм���Z���Qkkt/oz.�S%`��V�N�a�}��7];�?3F�7�{B��@⩣�[3) �ml]�{8s�.���C�hi��r��p�:b�$Aˣ��.�n�\컷l��B&�����������_}�<p�'N�9q��r눨[�N�E��wD�	��<t�7����t���q�0wN蹺c�wN���.��.k���Ie����u�b��-ķwL�Wi��̑Lh�;C������\܍�s��e9����s\�\��xx���^<C΋��B��s��qv�u�.�]�]��""#'9�9��9](�����wʸ]u��&����;�9ǝ;�ήlW����wRdɱۘ��2]�:U�v�Ȣ��u�y׈�8�#��v5�s��^/ɐ���y�{��1�D�&o�ąY�!��wF���%��ӷE��v�owګg#O�<gY��j촷6�tF�Q.ckgg�T}��V���)U3�~�#'-B`7�h+�^���򵧚^w��t���\�y�FW�5�f�W��Z�L5	�;)�zW�m�,���w^��5-LY��]�zw�_}��q����Vҝ~�垧r׉˒ќ��5:g�e�΅���ܵ��X��^��}K)N��g�'z+�;�,?U�S�U���5��_�E��,�M�v���y^PcV���إ��|���8`���L�H�o%}��y�\�q�H���<ίV�^;V=�[�{7���O\��w;������k�DN�VO��y���^ț9�s����Ѫ��_�{_�+��C�d�f�*�f�?myecsf�rag*k������]-��ױ�ө�F�	_����0�$~���qq���E!�O����*ߎ��Ot�,��I�K����/�D^vp;l���;�)�w��+�^^�4wV�#X�����gv�@Wח/��� Ӛ��k�B�鋩���>�"� �Q��+}��wkv����d��8��t�i���=�*$;W`���Iu˺n�u��c'o9��m3w)�D��B�]D}�%�i��s0��n�tvis�S�5�b����G=/(��X3s��퐧�q�?W���<=�+ݵj������:�z$���|���̭��c%4�s��=ؿi�N>��*�v'�r涄������9�F3�m�a�в�Yu^t�TQ��4=;���q�R�
��0ݓ�����x�ޔ�Iy��׻���/l����!\k0�k���n�,�y���wT>F��-Q[���2<�ԉ���z�34�ذO"6�TN�u��:e:�	�Q����xa;ڦ�P�[|���F~��
^D�.����ǽ+L�u}�����5ʲ1�-�/���囙!�S��G���c�4~)bߗR����΢|��ku�>U1���ǁ�����]����{�q��{l�c�I���\Tw6y�[y���0�}�׫�
�7��y��x���[߹+��{�s��_D�t�<�a�0̞�k���t�$
m#����`՚���j]d���Ij����Wmh�j=����y����ڵl���G�K�����0�u[�8�yՊ�%]DR��e�bI��,+�}\,ҫ�ݶ۝�t=\��́��۴�=�nwV�zw��E�ꪪ�{��gb�'�?C��Y^u:�T���V-�ou,�L*�S8**6��H�ˊ�Nvn�U���s��Ŏ�}�=:5֘s��{Դz04t�"U��:m�P���Sf�ʲ�x֓;H��{��k�ޞ�m�����T���:�AL�5�qa=S��j�s�ɓi�߉���w���Z}���i�oP�=�yg��S���,����߰�T3ayɬ>Yv)i����'
��NY�>aFC���u��^ס(�sN�l��C�N^Ϥܖ������ޑ)y<�èhg��̦�m�ߪ����t>W�8R�u{��\�C�e��J]��s�+t=���B]�ϟ��M���5¿���^f��Bhݻ�����ajm�zi62�/:�U���̞���7�	�o����鼷o��}����[P�fK�<�}���NvB�� ���M��7�P���ͮ��ѨX����Z�]�K�Dpp �4�rv�h��<j�^x��e۫�5�h��o�n�:�{a�b��k�7�q����;f{
�[�Ϧ�ڌb�0Ka�3�����O��H�����9�9���PG7^~��缾8���3�����m�Ș_��P�r�>���w�7�a���f�ɢF�<�k�#�=7�R�[T����b͞E��x��ױ�	>5Ib�N���t��@y9�/l\n��؟+q���VT'��_�r/񤥕z�e�X��^�<�7��X�ף�2b3�'3I4�iec��K�
�3`�K��<����~m��o�z�z��.��ǖ��N���]�\��|[��5��jo�M�{���&�j���6�]�zs����Fzwe�������}�4�uV�C�?z_��VH7�:��<yV�3��:x��ћ�x��~�]��.��N磶q�_3޿n��bL�&xz|qӒ�C�����U7/�t�*[�����9Nk�	\�?|��W��*`Q~�F�W��s}�ev6<gB�J����^j�����nYX!*��o=yn����}45j�����8i���q�}�;�G�Q��H�Ҟ����yc�o�Ҏ��폐��V����C���6�z�����GRj�)�:,�;;�b�`]�m�WT�^�ya0����c�P�B�۬s�s�^�Ц���""1H5CT�=�Md��yv)nN'9�kC���CS�����*�>,��P�麅{��P�u���=����ГU|_��PY6��"����ۂ{��Ew��_���z��;]��=�b�u�eN��P�P���sd��.�w{)���*j���R��=��n��l=�|��/<�}���{U>obiV��)`�P���8A�ά�X�ul�}�%[]����o���MI;ʖ.�۹�ݏR��Sw��L:^u���vɘM��'V�^�_K�{�ro)����yo�5�-�^�7��u��W٨:��ɦ��a�x)Y�<��D	������`�W-~D�})�)��Ƨ�%��26��X���kJ�*�������r/�*m��Z�~!yuW�:�����2m+�_��'�d�ﳒ���~��䯸ױ+��Թv�m�ؤ6�g&����:8;�2����5J�݁5e�|����=��j�ו��?;�����۲w/V-�c����ʅeJ9�����o��i��[�{a�1"K�mYvG��X�/y��"-N��A
:4d���X���]��<���f�6��}�T󢕱���a�U&�];m�ru���^�X��>ē��L"֕��N�~dG�:��IyN[��e$��zp/[q*�J��o֥.�=���(�DW����̎���)���њ��{�x��P;���"����{u�UмpF�ɬ��Q{�h�D����<�"�F��Q�v��y�����Z�n߫��]Y��B�vJ�V�>D��y�Q��ވy>Ǧ�j�D�ߞ��*��H���0���-�h���[@F[v1���z���q�6=0ӅQn��+�1Pv���.iY¦)�>�S����پ��/l��߯�9op�8ֶ\mBy
��Q�{@ϖeh�b��o�S����R�����6|�"3h*��������@W���I�T0 J����[�xy�yp{�UI걞$"�<.�f19ڥQ�9��:�nqք���L�>�a5g?���~PA6���AX��J����j�`K�z��ud��?*�W��=�A]Q7L�չ9˩���0��xM��Y��f܈#j���aKM�g!��]�uѷ;e�gXy�[l�c��MK�WK��E�S�ދ�w(�z��)�����[����y$~�z�=+�:�~f�K�.��]B�{�����y7�������j���-���9Hz�k�����h�O�Ŵ����;(e0k�v��wm����~N>/ō�����}�T=�r�������A���8������vc'���}����$��SK�K&���Υe��]X���9'��KE\�gU^ƪ��Y�9�.ߡ�Z��q�V"�͙��3��jf�re�n%b�����ױ◔�^�K}��K�?,�7�k63M7��F�6.���B�};�1�qu��M��K�kщ���,V�$|V�y��Z!K.�m�����z�%-V�Jro����>)ע��bM����>^���7Ӣ�۾�r�Aٶw�Z�l6D�-�������>��+=�����P��y��Cʟ�~��X�vP����j��8ۢmM�m��m��
�V��*%�r��=t��W1�����3���c�.s��S�J6=gӚ}�Ч�*�x�2)���!��0*��߯gY�{�2^nk��i�F5+o�%��("�r�u˝j:�Gv���.v
��j�v�ާ���	������V]g��yv�]��f@N}�!�x<��Iÿ���"�/��{������I�����w3V�V*�}6�Q>Xk�K�/��D�_{���M���ǌXZ\]ө�,�)���m|9��y|�}�~�C��9}�	V���ϰڏ|���!�K���O�ʩ�`��J��,�~4�K���US/���5�-��oq@B_�Ly�wdL?�8mw����1�d"�R�ߝ�F�u|ڨ����pSq�d59��f��!�SZ����a��{o��m�]�:�hO������@^8�
W��ug��տ)������q����[s��u���;k���h<3Ԧ�4��]K�T�K)�N�7��W�=�)	��:T��E�~��{���ؕ�Wܵ搽���mSZ�B�NX� "cğfK�ޥ�@J�m���	M�f���,�!v����;��|�[��0�J�L<�;�:�y��5,�v�Ò�ivo�-IҽE�qnҌ���Ƈ�IK����wyiS�Ȓ�y2z�́���i�nq�n�7({7",�Ǉzw�L���3rḀܽ4dZ��]��f���݀\í��S�}��=/q�~|�r��^3����ͽ��%TB�H��:W�ު����W�.�zu*K�xp��}صE���s߄�ƠW���۵ë�����5��5���W�Z��o��W>	XHz��i��%}�����Ɇ��0�|ʇ�wy�ģQ�.q{��k�P��;��=�Rc����.Q�jQr����x�T[a�Ǯ�yI���IK}CE�O5n�z��&�9���G��z���D���I�X]z���lD����/^Td�yw�p�|r���c܆�2�꾞9�ӞfA4���b�C�v:{%��������4��V�C7��l�|h��Ƨ��뗝^���?}���7[1Ga��e�=��i�V� ������@��5�M���s���KvD��-C�_�i�O��T�ug3�}��,p� G�Q��:^������Za�s����O����
0?x(��:��n�f����A���|���nQ�W�Z�]�mŚ+y�csfG����
ή���Ъ�^n;�v�:�τ�7�3J���z��W	Zj��_�x��$�
վ��0�;�
k^�V�G��ٟe���_�/���Wԅz���)�Ч�O�_�3�d�}���yF��<^���މ����;�j�i����a�'��Y���뱃�Ғĺ��>��N���/� ��4}"s�F�_(���m�^���r�k͢�u.�<�h���G��C�:{�o+�x!�S�~?{����	kt�M�W5q$v�1EU�c���k*U?�~�����U�l�w]պ��ΏM�+�Rz'���Uh��o��3s�"�����'{ݯ�>>}��m||��U���;�ӞH�u�R��W�w����Udu��[���=�mG��y=��5�.�-B�Oj���KE��0�Uʅ�ڜ��_]&j--��Z׻��֛�up7���=���7۔L�]-�S9�`�����7'�n�R�y�2x�k�F������1����z�0��-ؤQ�C0�|0j��FSwY���U�i�Nx�a�t��7Y��̜d�+5�g��;q;af�Lv�q����-����ɏ�t�ܡx�m{W��t5+s&_;�K�aH
˶%����Qv>����u���L�9}L`AB��N�{b�<��E��\�d/���:���k.�*Z��jM��U��m�X������o�(��Y�L�j�;Yۢ8���;7��E.�$v�Uf��T|����cm%����m��iޖ����Zf}���i�Wwa���`�dR�JZ�V�OePjݫ/�<53	����޴%�y6�Nqu�Ž��I;��I���f��^�\���Q�	�Ҭ���b��=���va���7T��tx�KN�M���v������4�j�lYF���b%��Dc���OgM�lM���5e�Mo0�n9�9�Qnv�i�n�`8��X��:����а��{����WҢ�5]��]b.CS᫴�
J���Z橙�4����C8��W�E*���`R}�ྷ6���#�G�.	ޖpt�K9V�؁�)���ձ�>�O'���;���t���6_�[���Hf�c��dr�Y��}:��"��g�}�:���v�m���q�R�9m��e��8ܼ����eoR��dl1gk�C�W����\�y�7�Hx�� �e�Vo���w��|jf9C{&�N�NL�L��1��y�c���J=�
��~z�~��uGfI�r�����kxlL-�Rn�
u����7(�A�-͇�璯���Tq�fN��v�MFgh��
Y��^ik/j��Ctgd�.���}��_FY�۹nE�&��ǅ���l�+���t�M�n��_a���Ҧ?��:��4!!jj��ձո)ۙ�[v�.}&c4VF��Z:�%�M-������q}��kw��j���<�J��Yr��U3\,�y6dp����kw��
�yY
��cɋ��7}`%�Ci�(�V�ܞ�U��h�Ȫ�L�|57���L��jF�h��L�n��$�x+� E�<��fkR��X��uu�u}�Үr�87�m-�]���N�,�f�:鍜p����n�
b��8�u��ZøvE%�ḥ�d,����M��V��!��6e�%�c�CV́g���t�v��b�P�Y��9�uouڅ�����u��\�Kѫ�;CF�A%�����K9Md�6����
�yi΋���FtЦ�YsvT�GK���{9���% ��ˁQ�M,�å�9���5g���u���x�
*]�c��ͧ��A�����c��&��
��m蜛һ�L4�Jyۣ�i"��g���d�LB,|�YޥV.����=�j�U`���"6c����;�hՋNݳ��GX�捨6�Xw�r²�����u��q��= }��}V��~ �$`'	9��o�׊<snQ��鍎���*w��I��F�����&i�J.m�d�J9͢Ɗ)���u�1�E��f)�x��#@S�5�E���II%�IFETd���Ȥ�AEF�H�&A�
���h�k���D�h��E	d�cdfM������#��d�mDF��F��^5y��6fع\�Qh���6�X��ۻ�у�刍1�5���H���1����4Hk&�ͣ;����I��QIZɬi2M�w]� �0���0� ��L�2Ko�R�c���2���b}�w3��b�R��1\���}�c�2�^�#�i�3�Z:�9f����y�+�y
�x5&R����	�RND[��bN��5t�������ػ	��{��(Z�������a�ۓ�k��|�D��1Pv�؁#�f�w��J�G�OV�O��<s�zB��&i8�pKp����z�{ݾX.���<�x��V3���)3?b�q<ڥ_iӀ�nO�I^����S��{;q��n�����N��	.�j���W�~�^�S�Z�m'v;�l�ٻQ�~�tצ�w)�Xh�.-�?#�$�^NTb�tPK�Su�cޥ+MܻDm{��j=Xg��?���V���eN��^X*-^�8���(���Z��SoϨT�������>F��?nA�-Ӓ��Ң����e�����ʞ��-n��j7��5�����i��6e�J�"��������:|�t����"v����s�|�W�]g29�����v���߽����V:}�c�IeGb���r��^�����&��#��>��:�����8Zb����S�yuq�b�W�9]���p��73#o�z��$\��p}p]�uooA��,$լ���8v�iV|����E�����~�^���%W�v��c�5�8�w�t�{��Ob� �*Nꜞo�������5K��~��f�bלh��t{�g�0�+�ii���o�G̮���o�j��
�ڵ+�����p�}�a�S�s�̝[�h�zzo�<[��;I?S���(��0�@����o��/˞<x�|�s=A�M^�%]�M�н��m��v�|�7��l�!7o�ӽ]R��{����R�YD��j����a�{}S_&���y�EJ�#����h{��"�]{P��n*��U�~���e�?^]��]��=u��F�zz�玒�b���{���X��Vy?X�\�b�Y�k�-������"a����|���A8��@O#�Η�F����Po1��<���O�T�I� �ƻ�%c�\��Ơ�i�M�M}�.���}4�n3�d�y^�դV�긊t9�9�7��fS�E����S�ҝ�<���	v�F�o<#�e�bʭ�>�Dop	�Qò�N
����o�b�Ł�u�lO�co���uj�!R���7��b_"*!��k��HԠn�n���/����fWH��m�s��*�}G�%k�'�}X��y�y|8�����c_�}3�*���iM�����S����\[ݐʴ*�N���^���8����Խ�OԲ�P���;ˤ�c �=���+��'��-�3B����>ĮΥ��^^uK�v���25j+!F�ʏ=S.�f5y�fMSrߢ�Iƒ���y_J�5Ǟ*!v��YHzS�"j���/�7/mM/?=�V�[��=�
�Si�Șv�*�R�;�o�֢v���������n�N磌�3+��zW+��{�l�7l_�")�Rr���L8v������[�����Ɉn��A-�	K��1v<r�a������]P�R~�j��Jq��U=��g3�z�ڵ��{&)�%(ex��a;�V<��a�����"$�L��Y� �j}^�|U��;�}\͞���UE�,�B��o��Up=��Qj����C�����z�U�_�`<�a�^�ڎ4�����ߥ;\�WD]��-꥝��N��Oz��PငJ��X���c����u�n��
z}�x��+i�Y,��7�-ԡ��RB��.��)��Z�7؃���T|Vj6���=�q�1�1��*v���p���X;4Nú1�|���Ujq+�Y�O�zM��;�z�[��#�J�7���m����M�=�jz�9�/D��ˁ�M�z�	�{�z;,�hҦ=�.��jz�9@MG:�@�Q<�3>=w�=���W��_��b���x�KԵZ]#�{2Pu��yM¡H��.�U4;���虑̎��~���,��߳���
�7���:ש�
�ZURȿ���=o����=7����B�L#͟s��z,���o��H�䣝շ��2��=���f��`=<7�lyS��-���3�{:nq*<�l-�3�TB�u�#.;�*���`���T�o��o��\�>�܋������5՛�dt.���c3����E�~��o�߉��`�K1��1r<�Sh��)�ܨU����>�UvRs"��s�r��Q��Qҟ�Ķzrp�������!�7�e�ˁc����Fl>�Q�L`�g�gx�������F&��U%��o6�%�ș���8˙��HxFq*�x�<�����ή񡄦v#&X]�A��h8��h�9c��Z1O�����v�Pi�����JQ��N�5�S&~�iW�.�,��_��#@�Eu\��f�5&8%��Ax#�Xz���L����  m�B�69GqD��=Ӓ���6��fv�T6�a#�-�T�΃�6���dt��VmI
\�[�T꠳(EQ[�VW)���RexN�>�?�;?uO��=Q�=��YL�L��͹��6ݤX�gvpC]n���]h��J����wa�ρ�}2�nUu��_e��7����r��.��t7��J���s9f��=Y��Xu������Ϻ}]%�x���S>���]���Bp�'h淛����꧰�=6kw�wӵ�n
��Q`qj/�.ERX�By����]���~%�_F�"�8{k��D�aP<7�kG\L����s�f۞�Fvdy5�@�Q-����CrMB��':���y��`�#�{�\Ѹ�+N�b��xn�/�k��u<��\=ٓ7acjW�\{��`��vy�]�yo�XLuZ�I��꽦<��B�4i��MP�)x[������׹z�eJ��;�c���,��x�	1���n����/����^�]WIL"O{y9j�0>�����{|��g�g�۽��X[s"|��Izs�������W���2wŁ�T�7�]������O�jO��x@�j���j�+�*Ǿ��2c
�m�[5���mS����z�}U��x�͗m?��< Ș��ܮ�؆�[���C�S֌�W�W)֫�ֺa}Ab��q]�99�����4^������	��.S�/r��N�����K����EX��YO_0Ҽ�^�����h(����iT��B&�FSj�z�콱{�Ls�Ye�t/�/�
@-c��W��(h�R�/:`_�T��z��v\��E�}'�|�!ݑ�5M�%s����ъ�',��=R���#�{L �O	n{Ÿ]X=}���.�)i�K�6�6M�'���':�;���|���\dϙ�ΐ�ڐǷ��&e�G���!����	L�S3�o#�g�X�3��S}]^_���<{qV
f��{fXw��.���y�3^�u}������o�����9�VG���p�g>�>�d�'��,�9s	�D�Ӻ��-���穱â۟���"vc�g�~��B7�@�P� �;R/=J�6*;d)�����jzBV�uxչ��^��#�G�uuGV����.=1-����T���]�?H�Պ�=G�G{Z��z���>ђ�W����tl.�*_��}o"E�W���̜^��1��߯=�9
�����{�KF/q���?:պ|%.���>j��Fw���^��]��)_d��j.�Ǡ7#�z �H]��뉉�yu�"	|}�0��F��H���,m�0��c߭Vw[:���u_�$�G����]Cp�6��v���N���Ǭ�l�a���Tћ�/�p�h�Z:����KI��{���,dȶ�G$
:��csF�U:1!�(	���퓊U7�׳�l��M�Z<*ڮ1�����ĀՉ��s��
�޾h)�U���X�����B����;�
���6C��:0*�1����Fב
f�����^���zv���G��@o��W��\�L�:P���k>�w�Gxޙ����3/��g����ɮk=N�ﺄǪ=2T�.�<j5�p��� {�%���O��6��z���b{����ן��/�����7G)@�}�`Lm;��;�q�����W�Wb*7����,�$�Nz�^%um����{s��*���ޚ��O��`L)�@�����<������/�lK���uY�>��Q��4�~�; !~톱��_�{���յ�W��OM�#��+Q���8Ow��s��Ұ�1xyv�$���R*r�@�|�{�W�}���p73�׽@ʉR}>�O�{�^_e�+3�N�<�B�v�/IEG{�Cx]xx�V���"�2g�b�&y9���:���i3���TN�ZSC�e.�G�Y|j:�Gz;�x����"�Ȝ�ڻ@We?�L�����ٛt��9��⛞�8:!̦^}�a��b�}����'/M�/�Ȅ}E����6������c�f:O�	���%X+u���:�j�?��s��D)�C~���cz���Ec����9����]�yNY�}/!K��v���!���{5��3�-�)<5���X���1�p��jUq�k����z,�E��N���X'>t�e(�%F�n�e�丬��n�S�I�W�jGՙަ̻�β�2S3q��Wd��SR�I�2��Hm�u��MayV�����������@o��F�P��h�,������ 5����B-ۤ�P+�׽'���S��Hυ��!��>�5����f )��ɇ���C>�g�ac�Z��7��׳�P����#����$W;�Ō�0[;yt�_u�f@<�a�^Ř�3c�0��
[�}��{�I������"��WQ*�h��\}��@z��ߤ��qއ�e.;r�	y��>����6�GTl�)���M©�q��w���j#Pf�C���2�X�����w�!;J�_��}��;�ɿ���,W�GTS���M�� W;&�)�q'v��k�hq*;`k�5����vR�~���3|���~����k�OO���>>�Շhy��w줱��z����"{y�gr"v�������U�q�����upD��}�3����;9�����:A���F��`�����uQ��̋�w�r;=>�M�.��p1O}��$�1����Wea@�'׋s7�nn�Jqn���@�e��d�,���"�>rrh,��{�M�\�\�у[�_�3�֏=��A� �ޜ�wXK:Ҹ7%�.�r@��R��v���,���+�Ebx[�[�ѽ7�_�mg��:&�9\��F���BpydG]���Zj�Θ���	=�Ǒ�V�?L�-b��T�2�!+��]2=N{�s�}����Q���|Kg#���T��Q]�f�z�[b��ٞ�o�����htl�f�&R/6d=���X��T�ۺL��ő���c_�es�c6;���
�֝���;��h\d�f�&X]��a�q���l�}�n��P��ޟ®��^�k���һ�N=�7B��uK�U���`e�͒���6��)����s$�����3��oTg!��eh�s�,��-ʎ�`=��sC����@�O�w&S{��u�{�fc�zI��yp����P~���{��PW���Z��r{<d��)�lEuP��V/�����U������S5��\Y�^�w��7{IF��Oq��@�t�B�by����[`]�+C�����Oՙ����n�mV���_n֎��[s1q�<T�x�r�.��2'b['�Gk*����ᱏ��݇����]��Qy޹�q�,n�	c)O�����Ҥ�	�]]��#�G��A-�"|����5�m6�eL��g`x>@$��Jo\��7���Ų�[��L!JB���#Ն�����6�8�z����9��aR�|[��Z1�����9��3��ek���r�w	V����U�mb��-�U����
75w"�h�{�l��Ru�:�xF�X,�t=��(��]Y�"��XP���zz�t��5Q��Ey�&�J�x��>���~v��%~6�{��*��СT��/{��k��+�+�;uT��t8�&GY.����t��g��ơ]�ꮏj�ĳ�9�6�ڂ���@muW�`~��&D��/N}5��r}�������x��g������;,��w �2�����U{f�4�5�U����Wz/#��W���h�O��\Om��zsO[W���͢�2�"��R<�CЩ�
���qT��>�ʍ����1|�+t��g4Sf�w^g4�1���s��?��y�K�M� ��~57/�2�|�_	n{Ǵ���}�L+�dc{��|��I�]��?z�:ݤ���~F��;� 'mHc��V)5LM���酝e���9e�^{^��g��J
��i�é��Ȟ���2*��o&x.9�,;�]X��*'q{�z�R�=^��9����y�W�#��v��`Zȃ,�R�����@�i͂�����e������1����UП?Z�~+�ӝ��K���|�΀vn:] �UH�m;�'�>^;M~�N�]f��~W<����8굕Y�"DY��g,���,<X�B����)�����6Ò�����ʬ���2v1�"%i����煵d9���F��2ݴ˾�Xk�`<�B���IԷX��u�=�N� R��{a���^�!��C��F�Y����"�Alދ4�s��YE3�KVWT��0]����0V>�wϵ�o�cŔ��J$���֠��H�n�I�$�:7�����"Jk\��u�I���Io)r�����QƚD΂����v �{N�*�ʄx�-4ޫY���w�h�}�Z���..�[;圩ň���Ճ{��$����躲�&�S��ȹ�{�>��v|�P�}ןRR�$���c�O���.�Ó/L�'YsPr����p_5p|�w;s7Sfж����z�յv�cB4�Y�c�:��ܢE�R��a|H*
��:J#���!�彸��c�B�W��n�!D-�M��-f��`���Q�0CZ/�݂�A�I]�P׬Xž�79}���wdM0�G�=F�[*VF��70�`�3YR��]��!rfR�v�����f�3\&���R�c���W�m�Va�)��8�%Y.[7[��<]B����k�sX.`ٌ��������.��Zw��).��V*���b��ft/� ��i�=r�52��B�ZZ��
$.�qu�K�g<�m+�܌���ݝ�'����wg"�����Q��:_"�=��h:L�캽��v�
�2
yq Z�Lm���õt�]���[1:ǥ<�̧AAIf��{��g��l%|�g1,�p�=6>��u�<7Rf����9;q�+H���!	�,�ug4r�+��9!h��F|n�.)�-L䯷�Yw��[�h״D2:K�F.Ω��/��W-s��m��E��;��	���<�۹�L S块:�ħ�(�V�]�zB%��y\��U���Vȥ:��M1�;�7F� �e�:��Ѳ�\FK�i�p�Z_.�JsÔ@3b8�x�B����o1ʻ-�o7G"����rFG�f�Q�����Gr0�1���f���,i�� ��}ik���Q�DMkw%������C\��b�ś�J�p�`����ni����������g���8s/;����z�wok��Rڬ��oi�EWh{2�@���=�����gWZ0��eF5�}@�4�ޕr\�j�\��׼��QήKZ������EɜI5�N�C����8w�n���MR&�e�=8���+ʔѭT&�c��N�c�U&��=��O�R���9)Fk� �n��4��30cJ�U�ie�9��.�gyZ6�6���N0�lM�L��\7�;��"��DV���1�̬c���#�J�i����+�}������r�N���iU�8ֹ�u,�%k�tG՛-[;
y-���V)C]V�Q���Vn�99y�`�靵�/,uscT���� 
&��sD��n`�d�\��4��э�v.�,d�r�DX���I�vJ(���Ơ5��AA��4��s\ш�ns X��1�\�U�ư\��ؐ�A�x�(�Q�m�j",Q��EEs�"�	ݷMF��AX.��4lmʹ�QF������`�¹�(M�mt�CF�-�\5�*�A,Y#EE͹^+��׍\��wme�st�L��\�4��.[��TW.Ewv1i��6�κ���+�&�(�lI�W#DX�X/��\�x*��8l�t�99�z�|�eh$'a3�vn�ݏ/�������u��+y�u��s�W�É��F��1q[ON}�#ƣ����S��X�-������[�;���,{�_��*��1=����7��p�R����&{N��t�R�H��y.;����W5�.�lz��<䚨z�`�^ʩ:%w�D����,v��`��_ǧ��u�1�k�o��hNw�v��Н� 4�@[TZ���7�o.&6����ľ>�@�xkxO
^�Fi�K�|＇'^U��8���Ot׀
�O�<κ�UU�:l.;���̳&�K��9�3��;~�͏q��A���&OE���D��ʠ+�WI�R8��f�Y���ף��Ni��Gm!���M�� ����;��3ᵴ*$��>�<k]W��J�fC��gs蝇���(W�	{k\��S�\�8��\po�j�k�����061��>�����Eo kh�����]S^Xމ�/��]�<��y��g��V� ���.:��,���VI�R�݇��3Y�u)~����;�U�Cy������M�#�޽�~�Tv<�u�p���q�����qK:��a^��[�0�/�Sz��Q��iC�{9)ߟB���o���;}/v���v����voVѩ�B6�v ���RZ�nh={}��V%��»^.)�W3+�-Cm��A�w4:7�k�:->�u}� 5a��o�9�V�*5�#��HCʽ;|�u��x{bo=���h��st�7nk�9������ڮ`5�����-�������{&�9Uig�0��x�K�Ů0ˢ���?^{�~�F}l�/�t�EK��*a}�h�}�Q���������~�eӟZY�^t�;-�w��g{ݻU��.8�n�]ؤy9TrK�r�\z�;�qW�"��YH9ϕ߀�^�Vv�f���\�s��C6Ύɔ��ٰ��ݱ���/�������Y���j����v5Ed��C<�Y�R� �z�e3+%��2ls)�Ak�G{d�����&�/:��Tfx{c:�]�_F�q��x���J�x\���˖��d�j�޽����!9��Y~5A0�(v����}�J��c�D��5ۿ������O���s�hz�w��0�j}Y�Ƣ�jMg��[�n+'�`��(�g�*|���κ"�˒:X�>��������y§���:����������wz�ڭ��p&�S��]'�칒+d���#n��tZ.Nl�F��/B��f߳�M�s�XʅB���=Jb�H]7
��u��(
��@�Q<��g�ی����D��>����^�p�X���\!�ݱ�J�ưY��4�>Z �Ǡn�U2�����gr���
][���C�	%JX2YW������U��S��Z��n������N�����ޥ�z��������^s��q\=Q
h�1�z��@���ʀ7܏���ZY�����k���r�h�Ua��?������X���_��w\-L�Ec�'�P_G^�zE���)����o�zQ�87�$W���~{+��m��ou�ǿ	�=wo����{l����'����Y����o]����t�vV�?r����Q�ܤ�{��Z���fե���M{�y�8y��/�e�Ol膨�L��놳�s�;����F�Ρ*�/��"�מ�6������g����Oڌި�/&�z4�^�waK]2.�����eǶ9�L�a-��}zHɞ�����?"�S�6�Y�d�=2��ِ���X��1.�3��n<ߨ��:�{��p��H���<�G===9��Ge?2���av���63�Z>Qn����s�Ҕ�K�TL����Q��k�nrJ�U
�����)�ɖ;G�Q��&;ϫTk�z=;o�ޝ���}��﯆|��Yy�����XU�Ld��ˡ-O~JZ�{�!�޸r��_�_�\�<���A���z]�@��e�-��So�PvD�zu�B��<[�r��;�Ue�٤YN�� ;ёa�	�:Azh^�M<�Y(zrz��6�(Y�Xm��x�{�n��Sގ������vr�[`Ul���m)�b|��r��+i^�F��#жZ=�۳��N����t��@l����T�ʉ�ha�n0{�ף�}�z/(���ɱ=;��ިw��7{IFߤ�w��E��%0y���rt,n6�]5]�I��O�(��=v�0dA����r�v�u�3�S\��M��޸�y5�@�H/G�E�3�i�����^�z���r*�H������<7r���]'��GǤ.��ڞjx�g��+��3y3���5,��yw�S�9M����{��~&:�+�k���{LxT*�B�4z�nC&�^F���V}���s�z���z�������qWf�aȕ��y��]&�_���C�~��2;�/O�����VO�UGO�8�>����cz�ȟs���_f��qUcEߕ<z�J��V�>h~��ć��}��N��;Fs�}'��گ
��^���;�BP��m��^T���A�F`B%�V�ye�],�Dt�W���#�oO0�o \L�t������ۘ~�w�p����0�ս�3q>�`-�C\՟qf��"~��4��[�? 3��h~�^ w��.���VW�x�+�v��^�ԋ��BH�µG*�7��u߂��ý���ޭ<�ζ��c�vs ��һq�إ�Z��m��[���C�uG��h�����E�$�����X�0)��Ы2r��ܮ��5#�k�FTU�b���;���ݎ��s�D^bg�8��~�~w��q�S����?<�O��t���g�7��'����
�οQ_�Q�Np�a��Zġ�ފ�o�S��z� ���2*��f�g�㤰�0�נ:�묭hu�6����oJ�����V}��Y]���fQ�:�����7��|�6s*���u[αYr��]��x�@|W��ݵ���uȫ�V��r��d�"����:=��T�}���o=>��Y��:#�8�8Wf�q��L_�[ONDy�����r�K�l�J��꣱z�Jہ;}r��+���wC����(J�'�Y����Ӣ��iS��3ݝ�CxL_v��CѾ\�%S�]����b��|`��*�h��z�a�h�ށ,u};�����7�����I��3�W�9����e���=�7�*�q�⹛��!vϪe�˫;�/���o	�~7%���o����%uY�Z:s����@Ovd�{!�P'���*@銽�&���{Mǚ�'�f��2�:{,�C�0��d�ˤ��WPp�P�x��*P�5ZϽ]���Q'�G�%;�cB=�unG��tW)��t��y�WG�Z9��iu�,9�M��8;G	O�-S��f�Ͻ��i^���<����
�X�6��φMQ��qt�����2=�m�a�������n����~�F��˚��&��]�zM���J��ԥ��3������{�T*:��銇�'�F����ސ7�ͳ"��Ƌ;���0�`�Vש�����w�>��O��oN�5�`l�GR@�uǥ�3�]�����A��{os�Mm��S�r��h�_��톼�z��y�׍����i����ep�yS'���z�`���{��g��)����ޛZE���b�3y|�����T��c�� �7�F�%U�U��Y}7�vg��ҳ�Ճd�{�kCy'O�g�] z��r*�g�7.dA��n�7��Ҡ�o��CT��U,��9��m�v�G-��{�Ca�xx��	x�"�o������`�]l�@���)�s2�Ni���z�R<��.��ڸ�}ݶx�t�,�u�Ñ��{����Pw[aO�=_��� ~ί�"�q��-�h6�i�����Bn��x��;E�����������S7t���Ȋw�*#r�2��;��W�`�q�B�<��C�#ދC
��hGO���p7>�^����s>�G��Ρ�+��n#�T�U#�^X�-���|�A�?g��_�']W��?�M���"@�nТ�o-�M:��Ĕ�s�,5�(F?ږ�ʁ4�ܰo�6@�7��p-��B}D�֩�Z�YoU[�T�u�{���[�8��h�q�\�`��*|��ݳ��s���1��oU���,�ӥ�������j�W`Y����}r.;���ϼd77�B{=FFzw��0�j}Y�ǟ�s^c]\\�5�����f�#��I���v�u���]�uNH��C����简�_u�eo�0�p��ݖ[ +=�����R6K��ܾ��e�O*���TF���㸈,��MhU*��y`K3<�<���4.1�ӹ�<2�z�óҦ���<}��
�y]$
q�˦#ٔ� ���p��7�����:���8=%{�ê��z��,TB���B�RdwU�Q��X<�!��z���Y��o�Ѩ	�Q�����g�^c��V�h)�?��H�	Uݻ�>�,n�������>*��O2ޏTo�>�#������қ�b�ŏx�h��CuE��V��+��=��'��|�s�_��<o�+�n;�X9ٙӝ2F�N��e�z�#�rrR��s�D���l]bU+ꞄP���=�_&�⦧�7��z�C�#|o+�2��t��4�lS�h�ZK5�2�b���7dw�5�	R�L��s�s�������xt��_�����&��"���Jz~}v���/_��W����y.N���a�G��$�}d=���|6�^g.�ֆ�+�(V��H2���GQ�eZ%*�m�j�p���N�n����b�(vـuJ�O&8hc�r��Gv����atgF>���z�(ۺժ$ɩ�
�`z���y3�p�E��vxP�����Jf�t�r�<��{~�Q�-;��F��f��л��$[.w�@<������X�ﶬ6o�sb���h����/g�yy�oye�b�^_3���nGtU2��UǠTvvX�)�%���۞bB�k�ő�_yέ��n�oR{�����p�UYe��BsW�L��da֮�}3���W^9�p��v�U�_�{�Tu��$n<^�g=�>�nؾ��Z�6|'Yܮ�O7��ǘ u6�JS������7/M_�P���v����J7���������˒��خd}���~�ջ6x�2�(�����W�o��A�K����ݭO�Lx�㲙�gz��޴�p�W�c�X[���* t�O��ġ۞�¯�h�<=��R�'�|�4������۫�i������=�^��ue�s&j|�y3U��a1���������l��ШK�&tgNZ~�8ת
�G�3$�ST;�}}@R��7�qPL���)3^M�����W��Omo)��V'�V����e�7|ʃc���ȯ���u��j���_��u{z�@n$�ꊟ��8���S�Y�a�Π�*N��md��T�=�m�M��� �������"��1���4�R�f1�fM�7��>�Z�/�e�2=���]�)��Xn�3NO%��k���zG���GJ�������V&����}�$�'O���z�q}��b_�����Bc�w��qA�����:�Fq�<�O��
}޼sӳ�BP��^�*Nv1;�KT�g����fw�g����yS�z��nG�n4�&;�[=�0.<����:�6j3�'�u��}�5>:�U���uHA�Ux�k|����7��O�v�jn_�1�<��	�n�K�A)��;���(���_���t�`���,���)i�u>�)�A�]ɟq�ΐ�!�ޚ���3=n�t�A��t���N�J^Z:;v�]�%ʇS�������E\a���L�\EH;�fkg�gmo��t�Nz:s�C���N������ϣ���p�g>�>���@��S:�+�wҥ�d�2;����w�����Zs���7.��dB�Qgr<�g���Qy��\�F�F�.u<�^���*���Ke_��`h�Ӌ���f;��i�rx]�+�T����Njh�u��s��UH�N����t��O2��ͭ��Ӣ�t�So�Gg�vw`�eu)�g�C��x�r�Ѕ�UΆ��'��N�"4�F��V|ŕf�Nŋǝ�d�]4N:��|��MQ�(l�\�"��qt���r�Ȅ'e�	����^�y�L��Oq]Jf�'֥Nw9�燭2�s8N緸�M���s�����[}j��m�y��Q1��߽�:醗2<���������r����;N�`�OI���P!z&@�yO���$y��g�.J���t����C�l�H]����������W��:��X����Pe-��yGC(u���nO7����z����@!�����#n���2t�j7��s;J�g[��V#���������5z�<n!oPp;(��g�N�.�&}yݡ�R3&yv��j��6�_�O`·���G����L<�2zb�D�5�t<�=�w��Y�ط�~�tc@^c�CQ��A�6�&o����>�����v�������-*.�\z{�7�����8�"���2=��U�P��zm؎|�&ցg�:��_�����M�_���57�x���7�����Rvj�m����o����v�xӞ���	��g�b�3.G�Jϙ;��>=o���5xf.�J�o�nug���4{>Sa��-�6�<����lis裃�շ茙�Mx��Kq�ŝr�ߴ[���}�,y)кS3qN�y�}�м�A��Q�^du� �#�6(�y��z7�}�qT��-|r�d�8�NS�\��3M$��Q�wPP��}�%�"s�@�<�'s6�S�v�qq��;X�N����lӌ�n�Δ�x��m��|^h�h�FW��#����ڈ�֎ꄓr\�{�)cz��5X��(�x�Ɨ5��T�C4���^@�x��%&Yz :i7����Vv׋�扤�q� �1
��\(f������.�>�a���ӆ��ϑe���e"��alWc�)J\O<]6aʼ
m,��l*��"�P)����|��n��X�x���5T׹�>e�2�����(��	YN��Y;�";�N��œ���>tj�`��`,>|u�N��ܥ9n�h9���j��7Z1֡Cv�����s.
�y��c�/�S��}8H	�;�賏Fj�������u����)��ԥ�1ޡ��o[�Wg
d|#��t-��y��P�Pa��{��
�L�2�9֎1QZ��6>�s6�X��!��������ma�#�L��T�]��"�E�!R�W�>�N��}�	 ���9�-��,���M�g����h`ۻ�]Y����}���@v���!�/���%%t�E@�?���TE�֋�1*���ޛ�D(�5{򗲵iwC�oH����*���+�n���+��Ϯ�C�{U-�K[����:bJd�L���꠨b"�҄���X��]��-���l���kh�����%u
��ј5����	*B�h��sk�c5�Nt&��g��1nK��@*AGG��[��3�/4L�2(iwv�G��;(,6�)H�s�e�U���d3�TȠ�Sy�hbV�9���jh��P��)���6z�F��7�d��{dl�
���ʸ
����x*5�-]��Z�Џv/��S۫Ʋ��y�XƝ�]ٕ�;g7�41>p^ҭ�n�}F(Uk@��g�Q�8ia��.!Ӳ�%f�M�3A��7�Ӳx���8)C[��[ғ�T���*�	�����mU�[q�B�eZ�˯9z���ڂ����6#���n��L��>1�l�/��/o;6f��n�VHtο{QἫ�h-�V�}J;��]ھd��q򤝅�	/V�	�]�uqNlu�V�K|�N�H6� �u �uCT�'7r �=��|�<ɓ��^6��J;}��p=���s^��k�e:�)����]6�	7R���x�v���o�:+� äfg(��ަ�9��_bxP�^S��6�a�Y�4��fP��� ��8��}�j;g����Ƥ����h��x�-&��X+;�ʆ{��33*!x��6V�%�pu�O�4�r�:�nh;
��	�{E�C�b�k^�-��
�f�9ӳ���se8��5�!Vk/�}�{غ�¯h��nf␫Ɋ�r�@�4ˮ���(\#l��qͮ:Jba+u��d�{ ����-l腦���˅���:�L`}�`�&�Pj/��E�)m$r�E$h�s]˖���X�ѹr���6J�����t׍�^.&�Ě78Qb"Bۻ�5\�wi#cF4��"��\��6;�1cD � (ԑb��A`�+���A��ƌh"*�h���ĸh�ʊ"�8h������-�x�ыEA��"!��s]�EQgv�+cb�s�,Z-"7+�[Tj�lV�E��fZ-�*J*,��h���clTU&�.V�,&�M]��;�*�F�cdƋAW��4�slXب��܋t�IF�ؐ�ڊ��4IcF��R�cIF��C���B�P�e�C
��»�����m��͛OSՋ��E�ޤ��\��ɋ��&Cw�k�[��qY��ʜʥkO���B�������[��Rr��2ު�y9Tq�Ǻ�G��Tx��mȴOxj>�����u\�AO|��
���FE���h���X��1��N^��^+��Sc�ŝ=�<=�}��S7�cؕG�] �"��
��x@��\ge(ɱ��ɪB��#��_����<�z}�V5�<��!��U���Al��S��2E�N�`^\�f�����n�;����jf�x��ۑ����.����O����R=����ܨ>�������f&ڟT�e�oH�}��ș�
�M�;�Q�>��g����	��ge�*�2E}���c ��v�.���l����e�s��m�} �9�"	�5��q�l��ɹ}@.�=�ʮ�
�8�l.��=�1q����:���8ں�Ϲ]�w�4/;�F�,eB�P�6z����T����9��ls��y�i,�j���@�q-�3U���~��z|6MG�s��q����%�R:����Ec�3�{N��\]�%���j�u�]��
�dԆ��f�_�S�M��'������^�����7�׏Yli*�/c���'g92)����(�'5ׂ?�7Zn��'�)Y�q�驊�Z�}�	�ʫ^���� �������^���7�O�e��Ϯ6��������w���2����o-F��Y��W}M�����Fj����q�;���_��qF&o��y�9��������ߋ��,��b�����Q��x#��v�� ��*1W��r�F�z�s�3�6:����fE�;׹Y�9��Uj��힥�l5��x)��g��%t����>�	�ʟ�~��GH61F�P�A�q^����x�&�kƻ&|�/�)s���F��+��L���sp�޸y�l�}퀄1��q`�G\��WX��uz�
�v���S�C	�;3ȼ��vxP�j���t�[���g�?r���@J���#�&Yؗ8�����)�?2��X\�j�f�m�|=} vmz�_o��A�^���Hp�8��}F��:�܉W�]��YL�d����d��&����.iU4}ޤ�ƹ�=�Ƌ����Z����2�{8�hx�ˁ��=��!� �3=]�\����GL.S�nTr��������
���c �=qd��	l�g���e�kÔ�Ƭ���+��;����7=��酱>���i(��<]�_�:����N�t<�jMd^f,��̬��p�_G���8n4P EB���ꆕ�2���Qq}���׷����OK�S|߆e�ٝ"{��K�=x��ʏ&lw�^Hyˏ]^���[�:V����\��6\w:�z& ���}t��e㑜As�r�X�C�zd6�5Q��@�~�]��]~0ۥ���ݝr�nf.�E:���lӾ��^��-��3]L�;�y����<+���7��/�
x��Q�qֶ���vv��������K��oB~��gM�*G)�5Q���fW�׋���c�LS�����O����GP�ΓF�� yI�\����T��}d�C�ܿz����t��_����O`��k������Q�;U,d)��H�����V.#{H��C�ӑ5��_
���>���>���5W���ɜ=�����\u�#8��������U��9U��޳Gt��^d��?�2:��'i��wΕ�숟W�����^7��G�oK~T�F�gL򧿕���֥os�uu���7NfW��.)�8c��uI����Mi�}G�6�w�� ��KUUxO�M�ϝ��Nl�Du+���^F�J񿣝��\�^C�ˡ����gH	��R�>��:OY�^ŷ�V2�����v�p���s�cGo����B�۩��=Q�y��E`)���B�@^�Q�}
�D���D4��}�c}��rT�2�^_�!{6��p��̞�����
=�9�H���}P�#����ޯE+�_Qwi��C�@a�����xcvm���:��}�N�M�쮦��/u��7T�S�ٕ�X}}Wg^��t/:�M�S�,�Y}A�x;�V)t�VӦ88��~��A���
h��n�����>��=�G$��w^W;������!wNF��w�a��i���q.��#�Y�9��I�Ҹ�ڜ����������7���WC�z�d�,M�d�U�M�Z�t��R����ƻ��9jopM��O�e%)�ڭ�zN���'���`r�UHʉ�h��n����e\fևD�i�.�*}�� 6s4kE�3Q��y�cܳ\Ek�������1<��|%����s�����O�1��wK�Oo�����z%�q�ho[=O�w�s��=�*�3p/�sp}$.��\L{1�՟|K��S��n���Ւ���� ����8��(�<� -����<�+�TW����F����GJySR�yt(ӹ���<d�C+��Y�ʄí�4it���*�����WI��T8��a�
���p��=�}⽵ѕ��O�)z�,�=9�k���&�X�T*F����s�k����~�:g�дJ`������F8���w��N����y�ɭ��>���O��7�:�z�=Q��P1����^�MT!Q��tɟY�,���S�<!�эL�/Y�C&t*NLZ
�����-����2�� ��n�T��C�.��&���A�.:�q]��/=�Ys�ۻn�<Ov��nf���SR���ً���%�2�qm�dk{Gv AHt���5�=	�0E����Ѹu%_V�w�����3ޚ��<=;LSL���|��D��d"�<����O�0q����^��Y��!��U�p �{a�@�_����� ���~�!>w\쪸���s�,�{@�	�l�3p�v��lzN�������T��rG���܊�y��]��	EƋJĨ���8�O}��9�ٖ=q�@LDbt������rk��Q���������Y���͍Z&�����q�>sT�>5���<�_�Tg����Y�o�1����q~`�W��6z:��6q���xG�'b�e��6��c�1Uޛ�h^�,ɋ���η�`{Mtw]�8��_9Tr� �F�< ^d�3y-�q�c�MJ?- {����>H��f�=����s�=M�dp�S��G���p;ҪF:���-߲x5�cn��;]+��*�"�}��l�Z9��ﳲFC�j:��� ���Փ�J�Qx}���&��w'U�7wTj5{���W3g����vGq�dW�꜑�G����������j�=C���|�J� σ]�|��w3�t�]k�g4֚��%�pQ�_���Q����x�=E�ur+�N�"V��ۍ��rF�$6�m�'�$����=��=i]��Mkt̥�uرK���.�U�^qGf.ԖI��rV�	^�`�M��^����|}/����Q�wTF�::��VM���ap�-=*�<T�/b�ړB����^�Ba��=Jb�H]7����rL�7o��ǻ
rM��Q wӱ-3U���w��b����<�~z��L��!�ҙ������绐���vT����ۀ*!횑Ϥ�>؛��\�x�Ͻ��7�A�K�vgx��&��8{����u3�ap���d��uP��h{{H�rQ�D��w�}>�\?d��V���X��'cE�B�f�S��οO:�¥LZ��"����+�{�l{�zn��p,:�jFm`/wq�Bf^o���2�"�3��^7��=��?.��-:���l�4�3���z.@" ��?C��*j4�??β'��z�{tY�U��J�}�_�y�ƙ��u~[L�ȶ{�n?\n�=:�g���~J�-�[8O��w^ނ�lg���O�߲g�y�!��p�Q�j�yȜǞ���O�OT�Y���Ɯ�w�C�_\{;��0��U3K�e�u�O)�м�L�,.[V ��^�4%�=�7?v%#@��%�:eX�g����l�2f˂ԫg�cuA�)d]ּ�T����d�ׯ��C�*�nf"�ŹV����79�>z�Aw<�e�9Th+���i0��+f�D�N�%�bޛ�[Þ�~���{ã�Rg}݁��Hp�:���4��԰�Q�=���JfV/b�0Y��}�W�=C�z/r�yR5�<7|뇂����B�����L��D+���C�pE�>���>˞���o��\��r��˩#q���9���v�t�t��@l�ˌr�lLH��
���ʌ�Ѿ�ڡ�n�f@6�q�����
�����*����wL3���#\n�Pq��fw��莘�f�>����`z������t�}�X����>�0�T�,1���	#�i�/ٿ����y�]i��"�^��~۬��~ș�~�Ӱ�/WI�]y�4n�ͦjz�B�ǲ�Sq�	�� ��jˡ�A��y�XLr�������qWޑx��ȼ�y;,���:�{dѥ��ST;�C�PK��]ӡ�_�f�a�Y�ed����2��\���Oqh������p��U7ޠ7�wUh�j�To`�\�qzs�y�R�+��[$�1�;��?"��x��g�2j<X=Q��2Ǻ{���xU�vKUZ�_��F�~��D3B���`T8��J���Wj�%m`�_�c�����G7Xk�3�R6��m�x�$��/�a>0�)�İ�}pa8� M7ӮP���Q�ږU��VFo%�ty�0�#w��z8���%��k������1���7��r,��\��vy( ع�0x�������j}^�����9����/[����ĭ����<��]+鮯-zT�WE�Do{#���`��w/�H������o!����Z�W�aԮ�y{<�t�����7[�.���>0���
᫃�_?<�O��gH	�g�<��GT���^��=�U��J؜�����یp��(o�hR�l2���C�̊;M�D��능F�����{��wg�Ά�l��5Պ�ҙ[N���_�omVGmN��4�{"/l��Fǵ�D� Zwp;�Np_s���a��|Z>�����_W�U�Y^�绽>���Cʾ4�r������W�\d�<'eY��������y���ʾ�.��F�3��~�����>�K������1���0O�-����sK�pq�˭q�r/����j������Έ�ο�3��C�By���a���t4_�����A�h��X�񺓩�^��D%
y"�D�������]��t������'��鉚�{Iy�@ӳ�e���n}�$�W���-�z��
3-.��(oVՍ�+����kt��ܓA�̟u7딄כ�!�����b��X!��K��]W�,i4K�8a�MT�y]F�
����\���#��t�W+�%s���5.��^�N��+�M$���T=ه˄��Q�O
^�F˞n� �>��]���jC*��X\TX��^���^����j���/��ٓQ��V�:ϕ	�_oQ�P�@\T���Q�+����Z�� ��Yr�A�T�0�f�@�o�e���6�筌�~�m�{��1�I�Z�t��a;���2&���Xr�������,���<ns(��~Ӽt�`(���:�;8#xp1>��5���s�;�Z��w�WFy�٠������=pz�y���s�]���߲�R������g�� wvV��R{����ݪ�~Cc
�n��X����^k��=�7�z7�l-�^a/O�O��H���5�q:�-t����w�ho0@�~�v�g�ק)��=���N~V.z�r�}�Z��*f�fxz�z��NS3.xc;�^!��F�ޢJ��d��"�R�ɶ҉���Ю�
����|�62g���,����c��F�y/�īW/ު�@���>��6�f����]H��aΫ��/�h��ɖ�dl�n��b�cu�/o3L�N���ԙ�i��?Y*������N
v�7����D���q���m�ePĀ����=\�n&ՓW=��1r'/)j�՜{�iL�BЇN���i����m�"�R�NV�q�5��]�']��qq�~T���j-"�oN�����GQ���]fܺ�+�[��@�̕�o%��ެͿo.
��S��>T{^���uy��@ɇ��gѳ�;���A�p;eT�]�
2�5���X�]���NǦ����WG;C��.wM�	Ύy�G�E���/�����~>�5��\����@Ιa��t,��w�-�+ޜ��Bf�f���7�:
���tDӪrG)xe����1>Ug=����ʍ�B����\F쨂^��ڎ��R7�.M�/�qݖF�~���f>�����H���=@y��ڐ2��I���i��^�P�zT�|w��c+t�2�k:n窒�����뀡T���/"��_�����&i�x�j/<�~r6�z�M��4&*��+����:xݵj+n
�ْ;f�U4;��@�dԊ�r9N���w��<a���Wi�t�"Dw!���Z��V�/�wu�qUR���Ox��뱶q�ؚ�_EȻ�8��'��U�3^���=��FY���������O� 6T�Цs��*`�ܯQ��V熧O�:���?}���qQ0��,���M
wS*o't��.ث�밸��U3�:��2��[k�nf.T����.�/
}���޶������-�W�Ȱ��b:��p.�W�1��VC�b�3���9o*VV�]�v�גBp1v]��t%�F��M�e0mv���|{=���/�B��c���Lܖ��CZ���9X���̈́ѧG:v����6�klA�
�[(t�y�g��w���
]�L(c����
��7EE>{V�l��̵�^giZۡi�S��qf��qig<�8��YBv����w+]���7G���oYԯ��D�Rn"(S�=w��?Y�Z�
�x�e�>J�tɾ��>��P}���S��ڱ2��ڛS�&2
�B�ﳒ���\(��y�z�k�]%fա�M-�S�,*u^�"ʔڢ.Η�F��z���Y����y�(v<1[k��C���ǌskcAX�����"w�`+��ٵ���Л:�%�t�ׄ��VQ�+��{E�Xp�z�R'�.� :�8Fh":��;�^�:I��V-�W{Yy3K�lfuv$P-�xzJ-v>+x')�.��<n�eq�}/Snʷ���N>W]� �ʊ.U�D󾮵P�r-Y{2���-q����_ %�f����Z�U��'Oxmގ=��R�7���q]8�wZ�P��� �=��a��x�rΤ�Vo�bu�.�U�ۦ]]���-3�9�r���ĳc@��1��}E[���-jU�ZrYW���z�L�:x�.�Ok1w�,�T��z�����%J��k&a�V®u��|L}�BWS���eaR�qe�A_*
�nS�5��]o.�G�#�2��=� ݆�
����/�e�i=���m��U�h��4L���VC0��|S�%C��κ�A·7�Kcm���cc��^M�Z�r�֋N�*�� L,�,����#�.���Xa;=�E�I���,X���w���{oSs�rk����n�^�N`W�-t��M:)�7��H:��$��z�e^ncj�!݃��0p�z��Oi.S��:Tx��\:�B�u�c���>��k$N��kh�pt������̃���c qe��u�3�Qk&c�L�Ȩ��8�w�aV����m�X ї�e	l�
��h���"�/Un^p_d���Ϻ
�X���+{�{���*�luᇕ5n�4U�ڠ5ʎKy�D��xNjp
c�xok\��]�6�j�}���u�88�\UuwRTU�U�!i����{/����oDvz�
�}��,���d<�Q�l�Ѿq�;V��@���ң��M7�����:R��=;|b0==��]6}�j͆���]K,t׵������w�~~{���{�.X��r�b�j6����y���EE�	�h���lV�nZ�Q�p�4�d�F��eA�Tnsc\�0!&*�60d4V��&�d�$b�eΚ���x׍�h�lX�b�2Rm�j"�C�M���6Jō�\ADI��i,c��i�3F������jy�1i�4\�(4[�
�`�����c���Llh�4l1���F5F1\��V6�5Dh�����H/6ƒ�D���F�c��Q�\ܠڌTl���iwsh�[Qw�x
�D _�i�6.�΂<�e��<v�@���8� =[�	���.��w�
�$��J��qʖGZ�r��G3�ބ���˹utd����ǕyW��4Ǡ{��p=P�1��8����snX����/����ݝ���vߩb�B��Fpo~�����*��ʳ�_��C�J�J	K]2.)�y��o���bb���˩�!�U@�t_G=���O�l���+k�T?S�C	�;3Ƚ$?lmp�*�����]Wە�o�j�oxO|�Yf�b�֤�_}�f��6˛��@<�����Y2����g߱�dN�>���s��{�ړ?p|z��(pG��}F��Υ��������r<�so�1�t2�ӳJnK�<�X�snXw�#z���c�D�u�S9E���E�S9�n�B�0�ásu8�Ϲ	�/d�ɾ雌�mM�nT;�ԑ��zy��D�W�}n�Μ���(Ynr�z�}1�2�OJ����c=�������x3>�Bo%�za����J7�x�����ncH�� w:d�F��;���`m}}�� ۥ��@,u}�Z8�J�3c����UYV���_%^���y��{�~�5�ɮ�PZ;��n}�</T�����D	c#�cӜ�# �w��%��R��ﻨ�+#��!���T�����M0�":�e�� �uqRrQ���gV<i#�9��ֶ����i!,U�>'.F��Ďu�ճ1֍wG&L����w�v�I��3�Aea(������]u�Ķ��q���+w�3Y�����nQ-w踡QZ���e�E�4;�S^7ӑ'�U�@�@�J��o���v��c�����E�I����r��Ȏ/�7�P{1ھ�hO
�t�4�@\���:��B��2�qZ&hv�T��J�e��{ntڌq���^+��z��wL_�d����o�ގ�2=�*D�g�L�1U؎����N�E�魦7"'�~�''����p.=���� Tc�<{fpT.���ȟ0\�sINl*=5}��ɓ�{�J��[|=�>�i���W��ӱ��*�����2T���PL�K<�I��N~�-����b}�{ _���,�Y�~�o!�@��#��q�Ft��#�-�5�Ѿ�]⩝�?j�ёy��bW�����p|_��}�>����ю46g��ﱻ7�-Y�wT�Jhz*bo�u�=��l+9�%�"\���=Q�K��~3p*��]H��s5��س�{��W��q��e�6e�{��o�Z�P���R���^v��ʟ�}f�Og������Y=J|<y�/'��!������5��q���9�=��]���/xmWY����'���J�z�g�`��܇V񮼂��_��;�C�3�L����/7uЁ�v��a�[W\+2p�&���
\�%��GN�)9�5d�J^j&۾��^S�} d�g���G֨�xs�d��h��P��1{B0��;��7���m�=(��V�F���%�u8������v�Y[�:q�p�G*���.�{*�g�i����;-�q�Vp�t�A�Ϡq��bz/f��9�����`�������Ĵo����u�_Ӵ�pdt��O2�6�<��|���U�׊S�,�-zG?:<�OOx����(wO��"0��t<vU�}��mOk��������%o�vD��E78�[]'���n��w��p<�wMD�=�s��Ƈ;W�Q94}g�]�T�ٹ=L���p��5�'��|\�sjk�
�z��y�t�*�*g��+��{��67JK�=>7�ܻ��D`ڃ�~�|�_*�z��oP��B������/vg��${2��{U��3�ՒP��R��+��vG�4�zX񙨏:�
��=1��O��	�P:g*�۷�Ԫt|;�~��dz	����[����ǲ=>��oN�>�F�\p����b�c�g�#��9�^�9�Cj᫱����9'�������|�k������ �G�_�JƖ�FQ��eh�\O{��I��VY����~�3U톱��a�r5�W�[�Y��g��um:T�I��'m����Y�m$��X��+;��r��wr��t����j�"��o6��.G�`롛:~z����6�tݡl���v� 뤨��C��wB��:ړ�fp��7��r�6�c��E�os9u��?Wl�粀��@Js|e9��]��8�v�v���4�2ϭ��_�缩��Z)О�{�XO����g����~NS3.xc;��v�Gܶ�'�\UBS��t����F�g^b<C��W��}U`{���E^L��\FL�s�d7�T�s�\<�Ɠ��T�wV'�*G��v㕎*���[99(9�Wh�xG�'b���h�F͆��,������[ ��%��=�9zn%�x������o�.�{���nS��̕�n#%��EU碳��"�5j�t5�t�Ny�{;�������w#�Cs����UR,j��>��nq��Ҩs��zp�zP�y[��������h�}n�\wW��x�no��!=��>����^�5��]=�� W)��T>7�0�"}\����;�ò��uNH���\�q�=��$�p��%�|�ݽ=��U{��!>�k�k�y����>�����K7�v6��V�fyjT'́˩IdDuO��Dm��u�h{��ρc*
���L.�r_ę���ͅ��[����(X2Y���Z`��j��tSa�ݍ��fv�I��C6�7��B��O���{�e�m�^�Y}���Kixv\/���v���?Y�S��3�Ń2���r��c�v8��W�%�i' te���Eb�>��:0��U���Z�����>۱������'S�!~�����#�7��@*"σ��~�����d�yχU�mp���������Gw�^¥R�"X��=qC!��ʦ���*!��R+��S�Wq��>��{��}�y
��f�/w�}��Y��=�4Tm�1)��V:�z������b�{H�r
����w��e>��1�����^�s��&p���O� :���EL��X<r��O�XX�ӝ�;�R�e
7qq�z���o��?���s�6�<S�?���}���'@J�!9��Toeh�gx�b���z5xU��~�H���N,wde?U�ɟtǙ�t��k��^��dm�d��+�o�cFqn~���:3];�Y-���mu���vh{��73Ƚ$?w��Ǚ��:'��j��5�h﷕h��t�ND�W��(��	�\K�e�G]��ɔ�^t����;���Y]A�}V9���X/�Z>Ǜlq�&���뇑�%˒�oe\z��Jխ�^���ެ��`;/Od��F��w�#q�y��cE�g_S�,��܊�7��Df�2�گ˫�]�	�m��)��v!$��a��y>�N��ӫ���L��:�m�g ܉��-��zb��ܯe�ژ�Y�v��^VH�|T������]�jL��1�p�D����s�w-�e����sޢ��r���nM����}/��.2o�f�a�7�nT;]I���/b�v1�1Ǐ,�.�Վ�5e(Ř�;$�}�43�3�]T�V.2����7���'��n�%��*�UU�sz�*�ۥ����G<�*-Ut�3�'��]�������/zc�7kGѨ��}G$����tF�֗8zxΠ��*��S<)^�*��5onh�<=����/�aHiݗ�N�s�)�N�a�<zB�Rx�>�@�V�T
�C�ٚ������Lwj�+�fT�^e��[���{�<����<���d��uǕ]���=���﫺�*�Y�f�51���x�}%.��u��2��]���J��1�.�������kþ�H���㯪�;>�`϶3�fb��~�5����^��=�x����Cr'�~��W���c����;!�@������33�+�_?��Y���M��Dc�<�g��g�Ki�x�<3���M>W?J��F>$�yչ�K��^3�s���J}韪~[S��!G���~�>U�E��ίO��lߜ����}�^�f�q$3����]s:{CM�f���[pW].γxc<��ui�R_�r��lY[����\<2Y��:���x� ��z
Mp�P��f��M���tɀ_hr�Z���
.k�y��t�x�I�T*8����B�V�:� ��s��]��ob�6�5�^ݩ¯l���Ħ��3z:�u]1>�=���`{��p���OOuO�KUQ�5�.���Ħ]��F��ffg���w���Of��6�1��P��&��u�=��m�3�Z)��T��:��{�3=��21]u�P��9����2���aq�Xk]X�ҙ[�o �qث�yIgb��9�x��g:g8�����}]>���@��q9��!����ʆܪ;_ӝ��gx�Y��������`�&k�[��6@T{�Pr)]^Ӽ�2q���M���;H�]�W�����땾�����纬�.��P���!s�XQ�lߥPz�Fz'i��ύ�Bo�e1G�S3�p�S�26�U�ҫ�X�:T���O���������x��7����FD�z�_����
�=�iJ�G���	Ъ6wK>�f�����wgfA雁q�+���!v�O���ގ����v�U9����<GD�yﲰ����L<5��\/�Dk�;< ��vX�:��Q��\>U�Hp���W@Sc�w�m���Y����{NA/B�0������j���������^l�ga��T� �>�Q��p�/�YYX�m�ޅ~���w��-Xi�x=A��,t�u�T��U�]ݙ�\��= ݠ�h�q�{h��T��F���ej��9ܛ�.ݾ\p#J��mW���{f���mn꜓|�Tɒ��<%QM�e?�4~�W�a�W�_*T��ID�S
��n��Ƿ�v;t�'T�\%@?�2̏��>q5��i��Ã���zt��0"�^�o׳2������ۓ�9��@��i��pϾ]��S�D���83_���z�����X�U�A�V���0F�֏����+�zz 'Z \;���'�z�n�}���ko�}�'
��m����z��E,��x�y��ѯ%Q�9�����@Js|f����u`�>�3�����ތ˰YèIL�^w ��1��ވ��=��괳��Ǡ&ofxz��	�N�3'����k�޼��ʽ�Z��R6�M�	q�_]�+�~~ȫɟ9�'��d7q�v��Q�~�j̭�w���B^�9�U��J���?QgT{��f�^SUU���~#����G�6l6%gp��x�x���v�c÷y��w��=���]>���螣Qn����� �ۦ��+�����鉮��P�-�N��ٶ�!z���=O��:�*�P�<d77��P;q]���|�J���C�13(Ak�������/Z��ꆣ^���V��3r���v�+;��8rL��03|�Ox���w3��u�v\�[�X�q���a��mej#��$b�4ѵ��,��Ջx�W8����ɴM.��&^�,���3N�z�НCr��j�W�x������#8PiDen�.zwM�s��o\�����<j�-N�5�z��>h�!5)���Oz悹}��3s�ʇƢ���}\����;'dpw��F������Gg�v�s�mn���d���x_��S;�z�_u`�@7�}��^�mG\O������3����8�o+����g��<��M�� 4jg��� dջRhc=��Z�P�qX5j�'6:z�*��pMn��L!��:���r��y]$�Q<�����U�=���9��n,
�u�/d�����j�?�h�
􍨥�M�����Q�	�Ϥ���]Gz�W�a߹�����uk�'R^���<���(��Ǖ�pD�E��y��T=�ʱq���MG:O��|���ˍ�������Ga�y뇟{�^7��gge�<���&��G���:��k��X����-��#*�����v��y*�/�x�u��W�ڴ��5�e}���i���G��X�o��r�*��jqy-
̧b{�޹F���s�8<���-���֖~U3�g�҇앾�:����d	��f�EO�b�,)1�3�
RCx��h��.�Bh��N����'�Ϧy+�M妛�% ���Wf�h�M���_Iin���'6Z��XkiS�>�����{�q�αuz��ϒ��<2�����"\i�Kx��9R����p޲8H|�Ý�u����Oj��9�����Wo��G_�������z쬮�=Q����|���"��y=�}[�"Wzk7�w�B�{�^�0\%,M|���ұ\n|�l�=©�Ͳ�c��
yOƀM�〪���gL�vz�l�l�sb�3��;��\��2�;��|*��u,���	��oP�Y�4�e�L�o,���Xz^�W�9H�������S���FϨ��|���&f�U��m��s�l��3��}�4=s��>�ܘmM�nT;�u$o���r=�>�_��5߬��u.��j�º:��W���ٳ�:����C��N������d�)��ڇ������Yg�;&k���=]�˻o�_�&��zw�H��NN��qP|%��=Q}��"�^>��Z���G��
&�g�w�lq\��ϫ�zx��.���;��y5�@�Q-���ʠ0m����Y��1�Q�iu��V�z��	c+��)</�Q��@��xª o�j}.+�f��3ZZ�.�Uxu�1}+d׋�U���X�&K} .�ST;�9 zg]	��Zɩeć@E�BZڵ,rػyQ�e"��\��`N�X��񠃦W_j@�ɂ��-��n�<�(��;��C{L_-�(�6�v�/:�5%�Zy�ݬU�&|���1���G� ����bs\]\�m[�j���R��GW>~�9��e�h�vg%��� z��DӼ�w�3 ���K��Z[��^5������IVv\��j��ܕ��c��L�[/.�V�J��pfc��œH��S��}���I�ϻ�]�.4�T�ҹ;2���%IX�`e�I��]K(]!t63]��xVF��x�	]���W\�v@3e+� UQ�33`��ۆvv��� %'ev�me�t���5�ՙ�Y[��#����5���{꤫�C�E/r���;�'t+�� X\��((��,�+Vӝ��t��R3�!�-�1����}:�yi�wz一��5�5��
�b�ֻ�9�aiT5�E��n̄ .Fo��jҳ�c5::ML�Zݘ�5>�@��A`�+���p��Q)M�]Rr����� ��֜�"ωդu��˕M�Y���i�S K���,u�:�$ p���0�P����Hf��ԝ/�C�G�i]��S�+6[�7u�EQb� y�N�&w�3O�Jޖ��X8U��2�˵�z��������0`�]e�`�.�'VKK�JV]>�������h��ݾ���(>G�u�ܕ�����j���$�B�7~�K�|�	�>���{�'{m+l�B��o�".n�,�K���2Ջik<&�1A��"�P����b�����	�Nj'a��tj�,�k3Y11:^<1rg���ޮ�WǓ�Y��n����웬C]��is�w 5���:�Nt�Z��NWaq�w{j�[��J�]�6����ͬa8�q��c/8�݋U�W��(���4Z��e�3��u�A���x��;�����u2�oj	������Z�j�ܢ���/��eU�oVhӧ�:�h"�i��3:��P�C`/3ui���j�����+weG0�"��;_L�O�e����֗Q,\��C�_vJ��jM�T&�;��x�r�8\��.ߵrāpc���¸
ȴ�{v�єO818%�\��J,#��r�6�+��aq�!�o1!����V�۾I�|,V��D�7)��'m�Y�7�7��*���X���#��rSFJ2���`]̜��ı2��<v�z0��)UwH�Wć���b��q{qsv�"!��Z�:�rk�/W/&v�e�m}����yHX�y<qC��R���I�S��W����e���k�)uM��@��c�w1f�	���]�t}@A�w՚FV�)���J��� �8&^��TzۀeH��*�5�l7�jݓ���;Xg[�t�Fk��g��g#;.���w0�R�4��̋HZ����n#�0U�/:�����d�lS위Xpc�o�Uf���-�#��ߨ�����W(��ŊHѫr�Rh�a5��2+�����"�o�%�b)(-ssX�75t�ܹ�S��r��.�e�1RI�ܢ�L5���Ѣ���^*5͋�k�I�Q�+�\�h�Em�r��"��v�c�F�֋Qˑ�Q�(��m+\�\�mb-�h�K��[�(�msIh�F�sT[\����-F+Ţ�QJ��d�cX��`gv\�����I][i���wJ���W�TQ�G��ɚ;0�,���oA�7�M��#͡�V�Ό�΋ۢ���^�B2f�<��e~��f�?I�ʎ���ɯ�f�P���c5U>�q؇�w�b��N�}��	�JV��w�}�SQR+�B/�ϧ�؛��2r�n<X�3_x�'k�:��@\��s�V5UU�k��v�����z�­/^��3��GP�=qշ�������8}r=�i`TДY��23�'9��?;�:'��遑����F��������������謁2��W��G�;dj+:�;f���S9w^�=�b]�ղF�}
�a;����P��n���aC��=='0��w�iܟ*f`��K��})r�w�e3x��jC�갚�&^�x�Gr�dk�߻lZ�9��܊�q���4���Het�����X)��L�\sfXw��R�L��LpOb�
<^�t��F�^�W������w��{T�;�4�{9�)��2Nw��sna��v��x�+M������v�����ri�l9��@&��x��ɴxM�U�M�����^q^���˻QbҾC�{�1����9��Q�}q��WIc=1-�����UH�}��pdt��n�gz����bZjz'@�5^���cI��]{rJ5� �s�o��짋�>�+{U��qF6�T���F����d�i!F�L�KN�KHLO^2T!GtԼ��j"h���sz�y\�:w�oM�k�s���L贕�=����5ग2�;��V+!F�m�C%�����������3��\t�O�GWe���q�¡ߍ��ro컡�W�:�Rҏz��u��Uڹ~������l�.'�����;m� �3� ��L��C��o!�s{-3����W�n��1��3���g3D��Q�x/G�ps�g�
���ov󬙓�{w6F5U~t}�<U��Vߢ���2k��9�5
�í�4jH��!�(���;}��SG��G(
�{oȩ��? ��7��d����z)dx��D�Ԙ0�t��������dI��]��|= O~U,ȿ�tO�w"ko���C�����������D���Yo;'��`g��ˌ��Wث�M������tj~v6h?�l5��\����=ؗ�ճ��H��ݲ����L	�4����\yS'��X=&������{��Rp�{���9�{��X�������=������+7r��k�����-u�g��q�X=&��x֍�y
�K�ϫ�}j�׏o�W���w$z���"��t��ٞ��S���:��OsɮX<<�O���́��@�w��Y���v�l�^H�g	Yk(�����9�Z��h}�N�tfЙ�7��L������X�ju;�%�F�Jj���иs�Gd�uT�6��M��nu��to��ڬ�-Jhtv��9�j�*W��l�o�y\	]c���F߽D7�]xx�V���*�ɟ9�'��{��<`*#���<�;�///kg&��7)��J����x�t�,�yL9�w�vK�=���q�-Yz��M�!B��-���r�r��o�:B�%ԼT>��q=��Qf7�'���{n�q.�b�1w)w7s��^C�SÂ�r�HԞ�3�_q�V�5(W�λN��1__d1�
��Ah����fsU֪�W<�We�}�kܚ���v@%����FK^V�b����q	Ύy�dxU���}���娳�K�h_�]����s�f�R�=${�z����{0g��S�ϽP�����[}'��݈	��ϣ�^w��y�h� tgu�F�ō8'̬�]�����O�@vwݵ}2�o\�Vc��$�oR�E%3ԏ���ޠ��Cɞ�=����\w�����Y&���}Z7 1�s"�U��d��D%��6Uzb�:���zT�.�I �D�}������������u��xi�q��e���=\�G�f�b������Ҥ����p:&dg9�L�Gf߽^�rO�w��:�n��О����- ��·�����䷻�8�_�{�q�[ΚA�p��w���g�"������B3ox�,7�jH���381yMj����r��f���8d�7h�!E�c��w58��yֲ�y�Z�]�#IOf��;���{K����=��2��p�J�Z�,���I��Ch�56+_x]	����}f� ub��~�XN^T.���o��ٽ� S��"�q�L7ە�&�{�i�"���Y�����^���T�����^7��e��r;=>�O�:wK���	��|D�
\�.p���]��V�U�z'��s֎�ߠx=�o�c�\�K?*��C<��2;ݏ�?��,N]_�m\a���>�@���E���NC����-�������}Տ�����e�ig����IWV���O}�ꅷ���G_L������\��u<�TK�q���aW�.�ȓh������/��|�$�
��z4�>�Q���=2�yV7��Fv�G}��c�z�
|���4�b+�=�I8��Q�[��z��)ge�q�)�ɖ9s�딊��pk�Lx}\/�o|�\v�ɜ��z+bz/׸��G��:����(�ʍ������n2a�7��t�W�/O2:�?b�� EQ�¯߻5wnY1�G�v�nIk�@l����uP��N������Or��ݨz�n���pm�nἹ�J�/Y�uJXoT���ߤy��d�wnqU\���,fu�����Z}�*:L�}�tCS�i�ӛ��1@�X�f�.k^qv�\����.���^5tj{���}�]�h:�.U�̨z.2�$-�����\��:��2��TŌt}W��g���x�ٞ<��^꜔3�'��������9�t�b���S��BG�Q*%pU�G���!������'<���d���@��Q-���o����6�HrrB��[���{%���P��<2��<*����J��-��� �|j�US�5��ۿ���"���\e]t=�D*�
�+�j<_�U�1�P�K���f��MP�9
}@WD� s�|��7�J;uVg�D�WPeX����f��{��k�����C⪥�S'�F>���ɨ�Q�D��t��oo��J����~��4��3��M�z���J�oL�����Ł1�����ݾ�쮛5�Q�0��mo]�;��R��C=�w���Q��9�y��~�[���`����f���Y~�����)u����3�:w�}�`_�v��oeF��{���/��n��l�uDZ��W���=~��\{7��!�h��9�~ bﶤ/l��y��w]��>�٪�1O��>�x��'黿V^Me�}�l��=�.��L���1H�jC���_&����u�=���C#��A8�m���9Ӧacڨ���7.�ȫӐ��g��\�ts(��o>|�޿����i��F1���9�g!ؽ��;HͺkmKIe��ĪS��Iv�|��)v�f^؎Z�+8���;g�bs��Y�T8��Y�9��M���Urj_Q]�y��/#�����S��Q�{��"�͓�x���a���2����Ub�1�U��ļU�R�ϫx���%�9�s�R�]�2\�l�OF��w��c�{���9�L�^�2�?5���V{����K��
q��������m���O�o��*���o%��y���m>���`ά�t�-���b�:��Ogb����\�<.2lSG���wA\N���o��/O�L{:�e�U�%�go���g��ӥM�I]��(_uq�y1<��(?>f���Pл�������(tN�A����;��,?�����V��:��������Q^Klgv@�C���"x'=2���}Pc&.�r��/���a��<*�����o�5��>�7 ���xB�[�I�y��'h2��67��H�=�2k�/Ǵ�/|�L=�2|�M��	�����w�����݀��P�zL�R�$�$�s�]���#Ӛg���>�c�{���D�z�N\�T�V����|:�91�yĞ5�oUp�y z;�Գ"�tg��7�ܪƋ����$��1t8��Ҧ忴?�ظ=�]
�V.ֺ��N�|��ו����VS��<��U�d]ʍ��VP�N�^䙮��ѵ�:�(��b�ΎŌjj�J��X��@6+,)�H�2y����d9��fs-ÇY}�I�e��(��8u�]$^p%о�Q�z{�?;�����V�1p�u@�uǦ�}4=+��G����G$�>=���^Y׃�n�P�mN�hWK,w��iCӱ��O�i�7�x}�L��M���ެ�o�*�]x�WE�<�:��m���'������ޥg�@�ݮ z�]8�g�s�.����Y�ǃ�ڀ|z�_���V��;�ޢ�����is���?^�U�L����L�����a9L�UA��@�v�r�^{Q�"��n���m{�%��%ׇ�]U`<yqK&|�0��Ti��|}��LVn�n�u���ti���C��U�Tx���DS7�s�� ��)���'c+������3'�5��c׵k+��辬�X�7�׺|�{M�b���SA��螣�U �!]�<�i��:Ժ� mn�M޼��DvO#8W�ɱ��К�.5�#��G���G�>���򨧾���\*�07qE^zZ�y<�U�T�����.Z3q<�����;ԑ�gG;�Y����/�n<(\�;���`����ѽ���y?�g쟚V�������L�^�gOO��$�1>b��T,��ߪh�;viZD���D�����y��tP{pu(hbj��)9؝��[9X<���y+���5�+ǵa�5��[Z�.H��R�s������;hڄSo���O#�f9�w��H�;�w��S(]ΑN4]�cjsAl�T�W�X��#��_Z��"��������z�_u`�@7�}��%�{�Go���Y�՘�v7�k�B���;�Ro���tFCʮ�.] ѳ�K��HV�$�X��Z���ƞ[XA�'s(�Oz�}�&zv�Ş��mT���@sā�Q<�3>=�~��W{�쫏�;�G ������\m1�4O
�C�/:B�rduz�/���_s��v+=�T��~�@7߼��e�tftY���RӬ�3�����,��1���T=�ʰ#ў�^p�Ƕ����ye��к���{P���=q���U�q/���0�����s����l;>��y�^��[�-�R��R:�6:�N�g�TB�mH��^�w�gt���z���{�j��4,V�Ndl��ۛ޻#��Ѩ�oeh����7�?Q�����ʇ�5q39r��ꘖP�����=h��j�N��s#"�y�}�\r�^��wz����'W�u���١�Ǒ��4Q��=B�s��|��Ḟ�<(y5LM��}9�\nDwm�a{��*\�.^@6��g�(;��rų5KI���F�gr���;~8����)F�	ڋ�u`K&�a��޽9k����x��Gy۔�ә0s��Yi�܇7c{r4��^JJ�,epCyӳ`�u��=�t:#�v�{�����m�*�u0n��P|��S��4�Js=�^��s=�Fډ��;:�ƅ��f�&X]�V7��{�i������T���W�d8}�ϊ���٬�ϭ�~��s�g����k�MG�O�|����Xz}G���Ѯx-ϻm��{�r �wp^_ɂ�}���n�3~��Pe_�29��~�W4=���]��6a����t�eTv��Ew��UW�y�{��lV��w�� ���q�4g��L���x3�P���R����r����"�ﾨ�]5��]�����=��o�x����"��S��<���Jr=v������s�"y�]$�a}�(-���3�S\�ٿ���Fw�w�����_L�9%;jRe.��b)����v]���˴�	ǉ�gK��M��[�dV���V�����'��Y�(���A����W�c�2�&�_�V�=�,T.�F������{Ęł���]���ΟI�{�%?t�����<�^���x}����+�b�S'��r=+�y8�f�_��0��n��`^�Y��]G��gg��n�<7;>�|L���{<#�@�+�v3wj��R�����+vs�d�PǕ�Y��5��\��k:U���Y:�ds_��EJ��lL�c���{�V���'N�����
#,�y*�k���+�Aq��0������k3��<������IݙI.��;�����Ќ��m��9�>Qܯ��Z0F߶���j��/�����%�Q}g<ri�%Ylz硔¥p4�遊_�\oeFϻ.l�<��T�>N����+:�S��=/Br��vo�9��jGz�6�a;����_*�����F�K���-�>��N�,��j��L�UPp���.��w��;�jC����/�u��G=����*x*\��f�D�*��:;�R�����=Q�<wqJ>�(T[��l��]X�])�����U������r�Ｎ�:^u�ds�,����Ú`=��S�*;d��No���neCm9�V'ѼQ��4�G�x�9��Q*��ϣg�Q��P����DR���xG������ދ�߽��5YT�ƻ���Hƽ��Q��]��H���=1-��� �>��>)�΂��=��������T��ђ�W�Z��PK�6rpu�+����,���}�~K; h��O.�������V�ň��,]�{�&ǧ�(��As��Ҷ��#�j�Z��U������m�m��j�Z�v�mkm�5[k[o��m�m����Z��V����֭����5[k[o�Z�ֶ��j�Z�j�ֶݪ�Z�}mV����m[k[o�j�Z���mkm�֭�����m�m��U�����m�m��b��L��Rư\̿ � ���{ϻ ����>�UT��R!)@�DUi���(�J�A(����(J
H*H�H��%�wF*�f��Y�i�M�j���ܸfW  ]eT��-�Z��pv�e�t������wRY��3J�J�%(V��͢�UU��T�h��6Ĩ��		R�dqh�&R3Y[U����	8#We[*e`Ti�mSZԉG��L�QSY�[Zdd�����v�m�5��&�mZ�Am��� cT;d���Yhh6�*%p;����K[[fJ�h��    "�ѡ���       S�i�)JB� �i���Mc�bdɣ	�bi�L#0O��%A�44���@ 昙2h�`��` ���M$@�4ѣ$4'�dd1����>�O����?>O�|�]>�BHw�k�xHH|O�IHMBBB  �$?�d! I��������?�O��:�g�F0&�@�*�ZHIOL&APa��BHp�����}oz��������$	5I������3S�k>�p䲔E����۟��~�_��q�)��gM����H1��&˦�T�5j[/w0��Ƶub��e���k��=����P�vc��:���1��M�-��	z�(��f���5)k�p)qApԻgt�SeQu��n�6��4d�)IL�n}, r�t���(?���Go+v[���I�"��Ԇ�i����C��t5BHB�mܓ,�ϑŷ+P�D֑�4t�"�x���Hv�pd����B���u� �u6�B��)�{��fV�mQĘ,PX�U��/+q��VZ�ws
X���Ee���2�ԍ+մ�3W���YV֋)�))�d�7Oonz�
�j�(&��ѹi<��E ��fn��Ѡ2�B��d�s�Yd)x�jPF��5t��VjB ����d$n�)���٘���j �-�[��͖¬r���Z��([����M�$��B)��"MT�]� F�&��*\}Cl�S��n��z�Y�)�[��؆�6}�D6��;t�m-(0��(�E5���vK���u��;�y�^$gН�a�7$���,Q5��݋��2��@U��������l�.7|��(�y[�b��B0� �A�BܓR�a�j֦Y�I�U���4��dT"y�HӻT�5"Y{��J�6%x��b�Z���mml����Q͔Ȓh�<��q\�miV��@��i!3�L�#�,3a�����"^Ld�p�xݼ�ed�ݕ����F�&��Qf`�TT�	�W,�*Vр&�d�/3/X�Ū�n�w��H�5��!%[�r�z��i��-HԚmٽ���3k��(ܗd+�h
��3d�븮P�+q��Ha_
�j�k���o[Rac.V�w���\�D*����e"^�P�,H];�o
nIV6�72���Ui�Ŵ�)��ѲMKF�Jɧ[��$En�c��֧zN�"��he��9�53h������1�Ŏ�݀�2�=��!"u67om��"���(0��i�FT�)}4l��sX#��Ybڡ�ER�)�;��r-��Mf;8v�3eIp�IO/Y� e���W#@Va�n��{bWBaQ�Q���eÔcS^0̈�z	sj,B��f&��k;p=���b��r+�Bƛ�o/�0Lb+_-�ʷX��Xܣ��[�Pe�4�C��Y��0�`�ř�l��m�5�'2<��[�R�#�W`�(��Ġ���&�����kV,P�{��m��$�3��F�����0k���y�Z�M�%,L�d����XT��r�<�N��[��k@�*�H�T�]��e2����z�.�Z6D�{�Y&Q@ԛ��kt�z6��	�V �;M�Q��Dw�����3���H�h���ʹ��#�(L�u�liy�!zl����о90ۺ���`�d�1�a�[����?��*�P���]�Q��S�˨���n�Y#Iԕ�͢eA5i�b-��7M5A����SQ�������lD�����P�E5��H�Z%YH;�.7,�-��0������ø͆F�mEm�F�*'N��Yu`�N���J�ے���:v6ѭ�԰�mǦ�͈�A={��{��}g�O���	�/>�H��ߣ�Q=ƾ$����������N�xE�T�R��kuHoOnۻ�Z���Z]���Z��m>��lՊ�x�l��qaǺ2��"c�e�u�n�g���}��ނL3pU���C�\��T�:,���l4�P�f����n=#��[��@��Ӻ� ��bVG,������[�E�g'0�̭�;e�c�;�^�|������_��qN��D
mJ&�)�]�X��ݎ\�TR���*�FkT�X��)Lܾ�cvx־�]$�u�N�L��?��WHx����Q�,Q,�]�+Ⱥ��ж�͙�u=��Vzx��R���k:���;�_m��1�!�U�!�Es�*�-�/����{��ú��_l1<��R v����jd�s�v/��/v�ܡ���e�(Z~������E��ռJm�pʍ��26�=�x+��/��V8,O��L�R7�:2ﲦ�;�'hz�^T��/���W�N�кU)e�XP=���9K:f곛�G�}\9��l�*}_ۭ��ZWd/��Ϧ3g���Q�� ^^�Ēb֬�˂HVj��{�a޹�GhЊe�N��W�bJ��RѦ�7h�\���l3�]�G�6��2*��.C�����������3g��,I��-����x��VRu�Wt9/k3�-�l�+=ܼi��Ӄ*��H�&M7A��gb���H��
:7��2e����>K�lޝU�a,��~���x�Wa2]MG<���3*D��m�r.�]'���t~��V펕��սCt�I�(���s]k�������y���ĹW��Jr����/��nM�M�ᇬq��nNث�]p�Z�Y#kw]�,�<��M�6� a,8%�n�.�v�Va,�Nbofh�ػ��2l �c�-o;���QH��H��4ԪC�%E�v��c�(w`�+Wֵ[���;��rJ�l�X]�N*[]�k�Ah��<y�-�w���� B� �Wm��w5�����m�;T�U�6�ˈ!��r��7ث9�w�Γ�iP5cb<��o�ˮ��d3��@'DGN�D�%�pG�_5G�ѹE^wG:앮Q�$Egww'o�=f�u��mg��*���v�P�k>M�6T�6G�r�7{��w	K�f�������*}�o���av,��)i&Ev�]Ms}V��+K�2��ܷ�v����}�*��9{y&YW�}�����P���
� �Zj�f�k�],�ǜ����N��8�x�#��Yè5Qr�;��u��6^���	����q);P�*=�Xf�N����,��Oͦ���Jň�����Our���R��5�J�!�2��}�^Q�\q�փ�c���=W8��̚�t�V͎�[��[`H�^��G7�{n��]$�k5�SnJm��N�B7Ҟ��Η>����b�lYt�P����=��-ӂ�.���t�=\���!�Λ7!�������y|�b��ܛ�X��0�򧥐�9�������)0�9{}�-�P1�%�С��%}VP�=��Gp�ڋ+ť��5�X)�f
u7��M>���5�_ީ���Jl���lN �+�%Z�Օ����&T��KO;[]�2��)b@l�O��W:��f��z��W)���9��e�`���f��[!��뼬��?�����}��w�ؚ����$	5�z�v� �����
}�9$	O��C9;�=�E�~�����I�`�����θG�".�b�o	���N�����F	y]�#!S�{Jĥ�Z��/�d|�EX*�h�vrR-�3D�dC�լ:�	-j�i ���ޅ����v��oQG���v�/��i�����j�xEq���.��k�����ܕ*j�'r�]�[��,���b���C��GC�1e�i�9����P���s���������;)Fk�i��gJ9�δDo��e�m02��j�=�6�O j���%j8�ƗUЫ�2�vk�<}��(��r���_�r�����sֶ�t+E��8�h�*P�7H�����8xn��n�
�*t���ߑ�%�!ި�MNS���͝M����*���WBE��&�j^PCm�:ܕ0���G�A�OY+Q��x����3,#A�=9C��6�2��S�In�h��.dTd���U��'.s=ջׂi��;m��mŨ���i�lg(���ݖ1�Ӳ�*J�]Ư�	Ƃ�ܓ�j��b�H��MA�^: �o��7�N�%�(�����	Ye�8�*�w�nK���x���6����]��F�&	`^NWH���VR�G��_\�ZdP�H;���ts�u�WK(޴�}x�5E�ε�f�o�4�o�jA����S�0Lދ.݇�v����I;��1�n��1F� ky@ռ�"�ۤ�
��e��?���9��E�%H�j��p�y�̼I�ψ]�G�^K-�@o^��@��}*�L��^�k&��M|��9ײ���~4)��n�q�I�g��9T����f��ݣ�iAۛ�e�KOSc�C$�pt6�*]�	0�EW���/+6t=�*��s!�J���С�j���d^T9��,�o����Ґ�pi,�[��lk7�;�iQy�f%3���L�S�\e�:�u�hj�Q�Vu��k��W��� ��f4\85���u/bkM���[���i�v�[�N�U�Z��\��͢SsMJ	VD"�Q��n���W9�C�L���DQˢG�%���ݦ�	]g]�`֧����[3Y��+�&l��-Do/���v4�(��Ŭ�N�-GhV\lM�I�Z4�c iP*�(7��	wWq9;��e�N2z�D�P�.�B�b7a�n�4)5,��UlX�7�K m��ߠ�!�gQ��ҋj^���$�B�r�8��b��6��N[�b��E̘���*JTҺwW��pQ��Pt)	u�s_Zx�(D�g(7@��)w=v��0�j׽/y�iE&��b�a1̼���@ݭv��ڴx`����&I���GRe�́�
��[�qX�wc���!�s��7q�{�/���zά�upT�bá���hۻ��Rw���X��<��D����nZ�Y-��
�<�}�PU��ܰ(v4t0a�t�����Z�;Gl�;�+v;��S�;1�:�<���VN���k��q�ಳd�y���;v�\��]����ˋ(��wg8�e���fl�q&�P�L;�}�J{��O�%��~{.I�EX�顝�]�jD`q<k�܊���� ���3�z�ڣm�����4Q8��� Gg�Z���vB��`�4p��'���]��I�r���֣������u�&�z�����H�"�_聲d8@��e�{7DdL��}�������D��"�Q;V�-��&l̮}ݔ��k�kG���H.�/Z�K�]-�]�ܨ���K������P)�e�bDq��9��dz^iV]/eL�����!u�WtE+4!�4'"5S� .p6j��G;o/q��+��:�λP�����sDV�m�Cf�9�޲����oV��=t�N*,G^��3���+��z̓��?( >V��b���ch��KHV)3E��,CIzi��2�b�`�%Abł�V�ɍt�za�P�7j
�̨����M8&5Y����bJ�����劻��������'�s��aI�����a�Ļ�[�~���Z���F��:2k�퇻��_��b������0���>:�"�{I����͕�;%�t �`�Jn.2y;�8�Ņ�Zu�lĲ��&��wj��=2=�3�F���&g��$\*��/�wQ�]ףWr��FK���l�G1��=u�n����(+(�^��05��s2�[<���9_sƬ�l�Ww^C���2��稛�S�݇h��b3ܻ�h�!������X��섣{�ad��h�8�Mi�}3)^�F��b�.����;vc��c:� �|���r�Υ:s���,r�]�jꮧ�N�&q�	�X�n4Ӷ,˘|:��bЄ����@�\w;���%Tb:`9�TD��xF�n/y�ۯ{99xx�N�*�w"�v��4��sW����l�m^�tY7�t���s��G�o�;�;b��s���-66�~�!��6���>?���:�7�M7C8�$o&Ǒ�����V��4��v���<|r]r|%?uU�flJ���ܚё�>ʜ\��P�^���Jt���t0������ҕ�pd��.v�K�s���n=���kJ;<����S���mN�qi眕xg���S�ֺ���k����i69�x:��?v�{+~\�u0��A�ۏ�75����v��ȪP�yhV���D�곘�i�<�R���ȓ��Pʵ�f���mL���џ\{Tvy�d�^w}NÖ��Aq�ʽ|M���*�B6F�0����2�Eor�(fz�:��2I��!p�3�[��&��z�L��X�\�)9�8��n��Ԫ��B�QhɄg��8���P���ݕ�dpjy������ �y�v�I\�y�|`�G������z�wzP����Hd�1����6��y�!��+I,���..R�K-ɾ��ωhd_9���8�x�>3�G˶��Fp��".���%ubt��u��\��<:�%{r�D�7+k<X��*b�ptE�t9��m}Tv�(�F�&\���䓢��ht��m��v�2V�}��#};rg�ͷ�,�t+�c�]^(x�#�ϱ�L֊(�L�i-)�/yX����rL鏞
��cu��9i�.O�=��h���<e_Q�Wg%���R�&��~Z�T�C�1棵�L̸���r�I��,�k�\�V��n��QQ:q��,�/��Ko�}�ˈ�
��R��}���<^u�	�׳mϯ�ۊ��u�������c6c:�a�]J�����$��z�{ʝ�g�����_���߲)�U���q�-ݖnuv/���h]PoT{>k;���h���g�.���2@/v�^CN�E)=��S�;8s�y렂ݩ�F0�[�dԊ�ŷ�+Id�do
�I%����B_Vd�9��V���nP4r!�E�VuD;�S2�C����j'I�Յ����KX��|�FP̠v��R/5�P�7�XG���n�k�	6��GZ	QWL
�'Q����n�]J����-�v������LyM#_J�
�	�̸�Z�a
WN�'@"WN	>ud���ݻ^B��6hR6���P������]]�u�(U�ywJ�K� E\��Ő���MRq�5�ɔ�%V
v�K ��*�\��<���SIAKi�U�
��12��B�-jVE�&0֮���Аی��G-ֲ.e1u�k,��HEލ�P�4�"6щn`�-i>����?|2#�w���3m�1A������GǴgTjV��������F^g�M�!�mM��m,�%ٯ߱�����|��م>���U�1K��%ĩp=��Cl���F����V=��8xeZ#��x�l8���@n�S5f%ω����[e�V'���b{�I�3�4��Z+ףm;S��6�F�º+r�{k�LU�"��7��?,��q�ր�,\����L�l���nͩ��]W�x�h�<v�"Y1�4�K�B�AP�����G������W�ʸ�+1�Osh٭���-M%��4�����GN���K��wj��u@��j�N;��FvN��V$�@1��yC:@(�C�wy�!6�	�$:�!��dM �K�$+i&w�����tHC�Bzd��,�ၦ�2I&aǗ���HH�I�I$L4�'L!��]����Ǯ�<dXNY!
ʐ$�v�u��=��o��1�m��I�Hx��BQ�9BLHi	߭���a�5��3�!�!��	
�M�:�a�I6�4����$9f�����c$��7�^z}y��:�a1�Q�@]������~�u�����Js��5��{�������U|����|b@���4�g�!!���Y��p8I&��9Cl��Hc$9`��!ߜ�f�HC�O�B�����	� i�zz��]k�C֬��V���v�4�r�`Ld!�7��!�Hzd�$����b�i$�P�Lh�^tkӲ��$9��CoI!�����HOL����$'i!�$;`bI��8Hm���Cׯ]�a��r��$�Y �C�b�\����L��W���t�oՒ�
�}y�]��6�����S�4V��8�t+��G���K�m�W�VXkz�R[H����Rf�L-�x�����܄Y�����H�{���))�8.�&\#D͞��zsr�5�2u��A.+�d�]���>�Ws��[�O��,�e�n��`^�'��\fEޅ=_�Vv�L�=n(U*\�#��훟��)<��M��9�˺�d�3,�eZ4�i�Ɂ[6�pb������6��ؼ0�S��Z�ŭ*x�X���R��nݣ�
��]G�B�g�`[@����1��|�4e�5�k�5&骋�W�}#����Z�z��c}'�f���u��[�d���q�}�u*@��S�J�1.�S��s��������ʉK�z���"�n�����\[�-dYlZr��}��XV=/��^�.�:䉴�vv��.�I�j�˵�\���չ�����(��.�23	T|P^���b�����{Y=j	y��xo���
ƸD~>z��z�i{��:��qp#�lz�7=�lֹ*U㎻��h�}
��P��G��M�Bͽq�77�˸�:u,X{q%y����>[ q��OV�u^���a��]�ޕ�{<��۞8�X�}v�?t����Q��zt�~��x+®��tp"��+�k��VB|s��}�CQ���t�P�G�V�5"'�������}���$<u�\N���L�������"k����*^n���P]?䱩Y�M�C���_wd�Hq�6��f�+��)�@�4UZ+�H���j�[���3aW�����_}@.�ㆌ�������C�ʤ���*�,��ީ6�d�u��'6=��"s�'Y�л���O�S���Q��Z	�EQz��Q��\[��h��k�V�w�r������8�����pM�CޝԖ�r���̊.Rm��N�sp@:*���o�*ɇ-ʎ�S@���>bgz�����:�\�!rB�;��`�~
��W��r�*��a1�+3� ���v�Ď�"U�^o.���Y���wY"��(�1�-�s-�5tr�Ed��D�0wqSb�`�X�>�v`:!���L$MЉeKT��h�O�F]Is��� Y�8-.��˙q�xr�,�JR�Pȕ��)w�I�J���������@�Qs%�_T+"bX�
!]e���D��3���*�n0-u�&[-�F�ckl�)lj66��
8���j�U���J&YqZU��*(�lm���	]]b���2��Tƈ��.f]aQ5CHT4�M9h�@#D8�3����f��A�[�ӹI���:���P��Zyߪ�1���'��)�$�C׼���=����z�T�U#(����2�J�h.@��aV�9�h�-V=�f]J�V4l������W��E��X[c�������/g��q8�o}�M僝I:p���}�ʂ��C�*�CB���|g�LUr�yt\�x'b*~;�����L����O�s����	�B�:I�
����n���5ot[�k�y�
)�N��H8ŵ-a��Gh>�y���{���>Yj%-�r5f��:����R\o���Sm��ߐ>z^����|+�튋?Vy��,�W|�i�퍡���]s�;J�&�]�[�	��s+ͳ�i9M2�Jaqb�����Lx}
�(�����9�|�Z�鋶�f&��+�:�{�x�Z�'.ޙ��t�f3Hp&�^S����
c�f�
Ҳ��UXЁ���
���Z>B�	��}�䧽R���*��E[ߊ���ʩ��������D}�|���J�!���;q9৭k��k�|Rt�yt�N[�7�+�^�vx͡�T:M8���u�&��Iy�!�Rbr������=!y�']ӗ��,<q|+v��W�ۉ�e8�ޙ�f�³���,����8xNS���pc�yl�B���i��z�F�5v���9|t����@�G�ײ
b��>�4|E!T/�{q;ur���]C�L��Զ$�/�t��t���ֽ��_}��I$�p���c� ���!Ld�ܫ�LF���2�?+RG�	�����h�+I� ���8N�;M��x�98CGr�v��7iw�\��C�D\I�k,�)�;{8�����ѯ�B�B�*e�!K�A�v��\ph�0W�W�Ƙ��������T���GƠ�>oV��
����7�L}G_��긏���+WA���롯>5�����\uO�@�I�Nڌ6�b��#���ﾏ�uEOޝ�.m�[8f��n׎��<C��aS�K�W�V5��Y�ۥ1׶�^�C��Wi���j�ʚs�o6���n:f�o�r��.����ޘ+�b��D!b8V#Or>A�}B��ӭ5~6�!��r�yfsIP�:����������3#�1��ܽo^s���վ:M�ה2�yj������uPN5�� "�׋S�����i�T)����o�qn(Jd��$���ވ�")l���x@��	�_<��]^X9G�kV�t��R6~�``��~���W
�4��r*E��~5������Ҫ�U��I�ǅG}}�)
#�f���
���������?1V+��Z ���^w6�}xkE/OI�c�����{���xp��i5�^�uDa��s�O�`�C�HpB�V��p}�֏�������]�� �jZ*��_)�\�7D�~4�=�; S�nN�ˍ��e�
��W_�v)7�ud_����<�ۏ��v�eM�Xw�֚����t��i�i冓�.o�*p�qNf�4tS����b��%|F|0b�q�
�q�3�5���4�F�Y�Hi^<�n��Dx���p��֬�y|��|z�{��C��V
a
b#���T�G�]��x���ZdCM{M=���<��5:i���#�Ð�{����Ѡ�>�f�U���}b�us���
��{�P]��=��n���=o�N��3�����o���3�gL�Sz��6�������Vi�Ak������V֘#4�?!L1T���+¢��\/LݧI�qS�7����+�6���oo��-��㾳�:9�SǇk�8�ݾ=:j����m���� G�,(k�׃qk�R	9gN%E1j��^<�n��̼�~q���b�#�*�T���t<_���Dg�c��9>�N'0Y��N]�o~�����"n_�?x����]]Ѻ�{Ƣܬ��ø�,5b�S>��Ε^}[�C�A��8}�yO��xv�1Db5���1WƖ��ǵ�_`�^@����O��n�-r!��!HS`������[�4*�L�_ ���C�cG��q�r���,RGRq}�'Bڷ�QX(ߕA�>6 ����ɗZ,}�������W�a}_�O��:M���=Yx������Lд�=�aN<ۨT}��q�Զv�З�87�ʗVw3���:b�0nMKeew&���;�R�F+���1K(���x�K�qv(��Y\�J��X�f�I��8t��	�ƕI��-%)�@X[�
u��H�Ы	y)n��R��9Ҧ �@	��*Ӗι+���.���N���~Y��[/09B��Z����ko3��#��R�$:0��X��K�aX��+�,6�pc��X+�74 ���/Z(�Ǭ�uc)֭�
��D%��Y�̙Y�	(�kZ0k��@c�b/t��*�T�"�ѨwK5�2�.Tij�+R���6�aU**�,���ik���4[��ڤc"��*"��۫Y��-.�TUUq��M]cu�TQUU�R�R a
`� Q ��4+���I��4���.I;�\����UW�}�>���*�Z�����1pa��Ϗz�L9;�9eM����Vp@~xuG�U���c<�-�6�K��:��{�=<8���f����'[�Ol�/}ӗ\�;^n��������7��Y�<��^�2��iuf3v����.�z�,���&8��t����7}7�����V�c
�V�]����`�\Ub��A��Cs��gݥn���	V��3���P�qK��r��0rO,%�1���.��6�9�,��}�}N9vw�L�ߪp�v���0xo6:��
���5��Q�1YL4�Y}ٻ�g�{NYf�SW��O�����*gwL�v���%C�^=��s��1���ue�m
�N^���<��<ejx�a޸:��;+V��v*�C^��b��KB���:pt��T㞰�Oi�]��-CL6��^<�^��;�T�
×�Vc<X�:���Vt,۴��!U<5^�*��D�M�|u�2��L�T�5�I��&�q�4�㢬S�J�a��C�k�����/s��r����u֫��8za
�*��f�U�}��/���IQ��:N�=u�\t��KiӧBy�v�*�j�q�U`�Lp����)Y�����]����<N醞��Nxw�>�5F�l?5�Y���ī²�j늴2���ߔ�7n&e�;ߛ��;9�s����[�iٙ�������m{���\�ig%ﾏ��ņ���Q鋙Ꝼ}[��q�Zy{L⒡\C���5��/y����;q:B���kU��6��~tg:Ñ�t�7���*,�{�k������8}��?n^���
�b��C�,UW1UM4��	*�X����!*0S�PZ�]����)���ゕ���n�]f�*�|�
�����@�3[�g��V�V�A�Lp"�
�Xea_a"����6�<SX�&wq�a�ػ����������"�b�]{�^^�]u��c4�y��p�
����3�dS���+��(T�^i���zxv��g%Hx}�@0E�j��U�*�y�+T�m�T�
���NL���T9q����(��\��*�v:�*�GC,M�k���gL����w�4�wNY��|Ox�(h�����Qƴ<?T�=�]{MV#�4��1bi������ה�m��E����q���!ǽ�����+Wt���ǥ�朖�}K� Zμ�c��a�T�T�Lݹ���ޫ}>q��x��!۷N�ͥۿ0�v�gt�+�4��h��{gXS����g¥���t�s4������.�HxJ��<M;N;���\oZl�yi��&&'z�:�;4y|��p�[�r͡�Y�^1�on�}s�gi��r9�%J���{2�;uLR0|�>"��3I�s���
�a�X�#Z*�����������y{�wƞ���	�/��(x�����M��#��}���������+BX�]���%�5�^F��h�0���g{�&!S�1�8t�9��+��q�s��X>��>���=�x�>d��^�Eq�;��.�Ǐ<���|�ͦ�мq���۶,JZ��:a��W}ݧL�o�G�/����84>�kA��]�
hc2��X��@U��#�
t �{�Ϯ�jϦPVQeX��l��Y3;/�){�̝��	:뮼׆��i+ö������g��YߙU� �1\>��Vk͚*�Unz~!C����%]%|q����
�R U^�`�i�^\/����>�Q���ۻ��|�|�q��/T���ǮzǾ����l��1.�޷H��G��Z5��K(�AT�|2t�v�e��N^z�yC9�[J�������5KX�ǚv"�^)���&�)>☸Z�ۘ����
��s{�S��ߕ�}�nf�G��a��8� ���n�����i���q4έ8O8��e��GOՂ�������|i�n���?l�+�T��=�e1�t��b"f�^�
�����6O�S���\�(x��]�>L.Z0���i���]�����9i��j/��9�Y��~�s�(��n%yӟaty_:�.�������?��؆�+���45^�~3c�]�nf�>�m� k��8p����n�:��t�\.� ��O��F������c:r��b�j��>{y��;�����<���XS|�m�k���MY���^�v��c &�ݖ��e��Ab.�Ŵ���uO�1z:Z/c�9�dp�n4�v�}����%�E-�Dǵ�\t�8�A��N�]]ϯzV���/7
�v��QEK$8{w�����{Ո��ư� �Vڧ҉S�:
�T&��ͽ�͢Ub� ����+i[La/�+�Uͭ�wNa�k��w�;�����"�/u����\��͂���%m�kv��r*]ÊѣK9L�2QI�+7�Xc�iH騆���v�A�D��wV�@0����� v���/r�������h\�:8��-�sk��n��}ݝÒ.�&RL��\�Q���ݢ� i�U!B�-u�D�՚�(�%ab�CNa��N!�-�0�ETEZ�tY�s&pUr�KJ*��.�X��ֵ̪Ș�cp˚�j�(�4p���"
+P�]�:qJ�kt�1<�다���UU�t�� �nJ85貞��{C��Cu�[+��yn�8&�[��C�$��!w�.G*��d�9�`��H�H�%�+����X��^�^�4����(`Iu9�]a}�8���r.Yb��g����yMzk�:�p�Wڧ>J5�?}Ql=3[�<�Ż��_V����yǩ�X�Wo����rPEt��kn�J�4�w�#��9�T��Na�aґJ�*����,�?m�1���0p���k���\$�-�l�Ol�Sr<_���}:^n��t��?�}U�I&~�=�f+�٤�μ�m���YF������m_u�,6vn�}��d|W�À���{�qO2����L ���qh��������eNH�^��tKhd��D�rw�h
تj���Y�n7��ю�跫
���LgV;nwpeww���W��d�@VKB��Y<9 �U��@�suCը_5����P���s��f�f̷����gu���-N��������i�q9u�|��F����Kؒ��S�~G5S�����7/�Y�3M愫 �#y$��o�}_v?��`|+�}y~V�N����J���J~��j�5Ӫwn�Њ���&�:vu�vۮH�x��1e,RW����e�,
�*�Ʉ�	TY[�`yQN��3�:���L`9Z_b�%M]�x����c��6����Y6s�];TK��UI��S���n����)F�E+�B�V&M���\���,]WOD����d��M֎�C7'��CC���Z�d�)�5L������Uh.N���d�]������S��r
�#�����v��#�ze)��Ks�r��}��-�P}q6��k�:��N����1)%�]��}��8|���C}��+�2��+5�6j˪27LC���l�r	�;�����N�.Y�/���'o�V���v�o����O���w�نK�y��]1������8'u.0��;���7��4���<^!�i��o���Gk+��lx��3�\񌶸�4HEj���Af�C��T<J��=痾s;�]fsҰ/�ڤdX�b3|�݃4��s&��.��� ͶN�$�����ӎғ�t�ӻ�}�7���j��"z�OEG��Q��!�sO�)��ot�~7l!�ʌkk'c..�3�R�n��~A���k�Ïb�����e��4����#�u��3^{k��v�6�k�DX�MW(��;Z�0�v룝V^�;xt�t��_#����~gsU0�%�t��^��'W������L$X����g����X���z��1Uܴ�5�םo~>�)��W稨���abM�4i8�L�]�e�&�v�������n��=�zRr�Άg,����b�Py��⚫ⷆ����z�T��K��'j�7��{(�';�%���Z��l�f��u��H4�!�*Ճ

��M�d\��Vv�t�B��߻�?����J���`&
x���v؇.q�7�*s�\;h��i�՝�0]X�\ծB�b�w9.�ԻU(q4r��m�u��%�}�����M����ݨ�%��ȶG��:�^�U8��FjY�9d&�]��"���
\��+)�:Ri���-*�ͩ���z��2��7��;�^���i��x��z]::oUM�:�]��	�(V=F�T-� �:���=�+!O�`��Q�ޑ���'�yXA۬�ae>��S�A`���� �/U��˱�ܥR�+�**2��A(֪��,S�ess
dEDE\n+k)+.�Y
 ����U\h�J�S2���Ur�L�]]!����Z�٤���N��5�~��L�1]7���}_H翘G�~�c���J"~P�̾weա�s���UƂ��޲ע�;A�k%�¾̦|�R&��u������*. �
�V�V_�y5�)%|��Q�#蒯�Y.��۬��T����~pvy��v;�Kk�U���wؒo/s��}�W:T@�L��$��v�s���~H<��W�6�#�����RӓY,箺�E��\1�`���#p�'&�����pA`e��tFI���<+��9@r��FS�n{eS�B�WZ�Q��C��{�n��zDZ]�E/^`5}�uS��6��S���Bjw��Rq����vW�����?�дn���L��5"-��.�ƾ�RF�|�m�`϶Ō��U�G@>�f���-����g�z>Le�.� �9[�j��fǦ��oIwk8�Q>��Z�Z�U]�B�-+��굹����[���Mߪ/�r�rۚ��C�v�;�(�����`�=���b��D���bZ�� ��Y�l��Az�rHo.�*F�g��;�G�/�xv9�w���%��*�}!�ַȓ�{e����*U�*l�ֹխ��9���Ò�w>��Y_�b�'����>�ٷ��n���^Nٕ�V�[Lq��\}��1~��L�V7^�/\��M[OR]Dz�'��㞽�e%� 3q�K3Hmګ��p�Y:���f̛����N;^}�mn)�c'��ZVU�96���2�h��˔��+����`8w��t�[����]����>��*�Y�K �c��&r��f-M��d��P�Hpdk���ik�%'].��i�f��G5T�l�N��;������iTƛ,m��lŲn������b����^�ZJc�L�Ox��P�c�r�����$�S�(��팺��ע6�@"���R)�ͻ��7`��T�Bxg�p�&���*�f�GN���ɮ�`!��o7��u-ՂC7l��-�\��U6�@a�^qkn��}G*s(��4r\����H�Ɯ��9�^�5~�]�.�]¿��v���s��HnS�-)gi���)�Z:�d[����Wm��q[�z&�gMÜβ�� .vu�hEL�:�}�f�-��R
�S�0;�`t��(w�����f�g��W��	�tZh	t��H�v·2���"��t���f/���?��հ0�_��5⚒��n�ӌ�2�E����׻��=ܜ�Jǖ�t5��iXn=�r�0v9�'��ヱ(ꯔ��a��݆Dk4�ThܪЉ��}�uh^���[[��0��3U$�y���6{�-s��=���{�_�L���_��{�3	o�[�J0x�-� |6�x�Pa�~<@/�8���O9��p^%'�},L7X���fb[��ĎQ������s��Q��R�Ew�����\G�D�� 	G�m�fK��x�N6�.�-��N�w�kE��B�啕B((��ĨJKp\�\.+J]�]E���F-�sZ�'�6�smr_!���>�ES�W�����Q���֬������J����ԎV]e�rWg`��bM�Tg��C�z�d���|��\��z�:dwD�(���Sv7���i�g�-�.�U%�jH�È�����
9�h¨VnF0�� ��X�Dk�v�ok.4n�˫���R���� �FYhT��� (�����$c�� �[a����bRřX��,��!�V�<9����)�K�:�rۗ����Wz��^�	��#Z1�ۊ��Z�mJ�+m����
�L�rTĨk3��Y����*ۍFa�&���iF�R�Q--E���h��kkM�@
$�F���B���~����10��dJ8�.r�"��yݩp�9F~'�՝�s	�}U^�&���ag
Uشv���1�yR��5�[G>�=)Y�D�:���5�"�ɼw��5 ޑ`jԪ*�'l+�&a�F��P�SN08�^�|�o''�h��g�}�x��C��M+N���அ4��^N�+yULc��B�5��5v�{d�9@��kn�����Ԫ���=�nj�Vk�R�N�o� �3�v<�'��p������ǧ i@���ڋ��ꜗs�؎�O��i+�D�Z)Q��;��wz�L(�ǹy�8����ݽH�z>�n]z�L��ܱ>ߓ����w��.�����ֳ�)[��n�� #���<y���^^�4g��m�iP1y���wMSb^��&��k�1'`�����A�8�v�~��ݝZ�����]rh��8�Z�8�ﾩ#��]���N�X]�V�w�8��<D�O>7�����n���v�gnI%��O�Z���#;B���{3�@l&�*�<ǁ���s�
qw�}K�+��p�81���ˣy�L�@�����i�4M�Z)��~{Kz���{���n_j^��1��NɊ��˙��y?�Y�-SJ���c�Ju�!�R��6cs����vqH!��G�Nr�w��u��L��Nۍ
�8�Ɠ��bY{��š Č2�V���Z�K���bz�P�rP�+ϥS;��V�r9�=}퉽��_T�!|�f~�c���+��9�I��J��+��H�U��MP����=�n��{D�t�{��U��$i�KA����w�bUUЦ���Cy��ʭ�oT�/��p�5/T�����v6of�*����v�[�ӄ�w��t�Q�����-?���h�R����~���^4tG"������+����.'�Ɂ_H�ا�l>�rM��t�Tyl4��4�ν��%�o�w���I��������r>��v�x���Q)���}�{�w`��/W/DDDB�~�{�~�B#sE%�z=Qx�pi@/,>�0L�F�0Q;;�:w���@d�G�x;Ù��x�;����d@�n�ww�"zu�����b���^�ޫ	p`���hP�Zl�f�_����C�z����'K�������}_}$�8�?~������/��~��ʼ����P� 	�~�i��X��3(����̶m����B��|܉UT�LN�7�&���Ѣ�7�<P0�im�
l�!8��ޢ�u�ѭn=QS|׽CFr�Z����A���Y�w��x�r��\����د+�s��=FA��t�D߄-�'�����G��X����*z�xfR��uKY�����{N]�@ʕM�C�	���K\�S�+�w7���U����h������~GR��1)j��gj>�ɥ���۠���:f���_�Zhn\��q+;mk��:�]�k)l����WC��kIta�]�SA7������A�B�9]�d#b��6�d'NႅK�.:�H�%��j16ugk�.��F�쭘�p����������\�l<�)�b0�j��l8w��L��t]c�P9-H�̷��S#+���Su��R�+�V��4��� FnZ�T�e�4č8J2�.
�9�㖇�	˥W3����?#@� ����!��1;/�Q���2��X�^U��!��V�ק5��X���N=:� ��U��P7i&`��E� �@J*�8�>a�Q[Z�.��Q��6[\���իm̳-J*-4�M8�"�Fؖչ��֌�i\73��8ܮ4¦�5�����kh�U%2�ZYFb`)�r�R��nZ$ѪD�¯�1E
 �#�'���4��9N�{��UI�fw�Yz�;�t�j�\8r����4��-��x���S4Vn�5UZ:k}�� ��y��tx�9z��v=I5�9�z� �z�48���a�~����L�pΥ�[��!�
��!��4Y��N�8�"z�{�+�Z�/}.���!j�s~�)������t'�7�����Py�a}�4�	���0�>�!$o1xn�f���,��K������,�1h�a�q��=;�R������K#H1-f��ٛά��J�5��QN�yYS���S�i���b�;�X�{�I�/:F7Y�����r��I�;��-�sҌ'�ug\��,.煰�~;瀽\1�!t�_=��]{RR�ϋ�ݫV ���[�a��`����^�Ȳ��ؘ�{�J�ӮŸ�:Y��6����|��ʠ-��2=����K��ROr��i�\=��o)#-���x��^���b�<}����m�S2�3�[}%��-Vډn��>Z����eW��4�+�EtT9*�Wޣ�k��u�eF|��t!ܹ4�r<k\X/mj���2.@�97m�\w�I?2�J��uܕ�Q$Z�=���3˫o�:�~�%�4���-��WU��ԛ��kUSa�n�u��5���.KUl��X2܈ԯFC���К�2n���9q��)�L��탶-�#�D���m���g�g\���p�n�����b'�(�>��eU�X��&��ӈ^�w�R�`F2�Et�Boo@�x���)�5�un�t��W��X	��9�Z"5Ŋ~�bh(X��]gD��95V�[����t`�A��s�Û4?$�-��{Q��^\����Jn�˯��.{vm�bX����ߤ5�̬��&�Z�J�8�Νy���k;�F��?W�e�9��$�$SW�M�o#nEU�ܽQ�^yXj�"���硉D���s���u�b�$�7{zts��OmT��
ի�S�d��4Gs�_9�r^Zx��j��l3B��T��ƻӱ�0$}U�7����b�_,M�g/w�4��U�=�S�Y�j o �9�ׄM,����=��`��8^�/s[zk�{ۭ��ь<%�9/͢WP֗�O?n��e���A�3���y�K��Y��g�,�Є^�j.Y�	WXM�{��"�7��jj"bDd�Q���0visۼ���;�&�f��?5���%5��Y��H(;�jB�rn-ģ��;$�˳u�旝�_`wE	��~���o3+FB�Y�1�� �8pw.�x��Y5w��t#kx>���Ap`��6��
��&s��r��ҽ��:��u�WJ.��AT�-W�헤S����,������-νy.��$�'C���!r���3/^������m��h��"�:�{����]q[��V���4�f�:��GP,Zr��j |%Ȏ��*��� 9�94�up�ַu�́����vN�a�e�}�V����}�*%��.7�'��9�-g�D����0ةU�;��q�R+�|�����k�p�Z���s2s�����EZL5�Zԭ撯N-�[�{Y���⻤����Õs�Fܢ�\�o��ˌ�G���f�R�?�*)1�x��V��qf:�$䵊�dy2�#�2]2Ïe��B��3s�Q�Ɋe̢��"5�q����-��*�)h�j�h��,���k�R�ԭhV�xJ�����2ٙf���`�cDƕ��(��Ŗ�J�6�	mK1��S�j9�,�KihUD���`�J!�H����3(e���V�iV�ڷq
9E��ػ�0X��������9����u$].7"ܕ���{�ޝ�8װ�D,��c�[�P��YЬ�Ō�e;�q8���b����x*�+��ͥ���̹��:�_�őR��ԕ���ˋU�E΍��@*o��� �+��zgW�S�b'�+�������<��xD퐃�z�8G�������g������B��#����"[�p-���x5�o��2�!�ۖaC�Hw3.�ȕ��� ��.�m����!�`-����|��[.��3q۰��<�My#p�u�n��O2�pHf���=)F[�Z�#𿸬,��p�S0�Ll�w��\s�V�u�<�0�d��]W��x:�8Źx2ت{тxܵ�v�]��uJ�K�w>Eh�,6���ׄ��33q[�*�;-QG֒n�wBus���S���n�s���	�ī	����w"�k:1�<�`�W�_�[���{{��W�����շ�i�A0 ��sS&b�w��^r�:������k��@<3J�;���b"i+t�D�{��x��uc�ͬ<�s���wsJV����(���qB,��W�h�4���K'�uG�-(Y枬�&V�g<xNr^�W��b4�ku��ȝL��$~ �j�վ����:>k���ʱ�6�`w���R7�#��agNj�:��g8K�Vf�SN�uC[��^��Ik�%���r�T��k��yZ��O'�3�6F���琶�n[�bu��0�tE�Ok�@����1�7�*99�F�C�V=Ǘ�	:��.��\�Μ�)"�s�{�昝�\��D�u���0��uĿ$¥7+G��H��l��Le��䤻�����,�)sʁ�WG�N�_N��7����G[�Ŵ��a�ݾ�ǡX�66X�"�V� �X��ɗ�{=��
���>�r���㏹�]T����ӎvn�{�f�Lb�	�f�^�e�T}��U�����_kXXe��&�-;�3��'h��ұ��b�5+�P��I��"K�e���ӕ��3�#��z��>�^yP���ѵ�]��[�J]���~��+��D��z�2?V���	j����7��8U��V�"���]u�g���{@xTn��րRc�b��at�hK����uSg�L��Y3�W\��b���a��Ry��=;��W��j��Ŧ�j�Y��Gl�<�G݇�'vIϻ�Qo�vĮqu�5L�@S�0/vG��#>�%�`�$���OIr-0����$��9�����8�m�,��ȷ�n���S�zbt	F[�E�OnP�4~�C����G����Nori���0���)��)%�����cr�1O��8QF����Rw*�*;J�M�n}�����"�v�u�]X�h�F��P�j�*Π��o�=�[�����a�ԫU�21�i�\;��s3kLAP�lR�5WB�G;�S�.d{b������sMR!�]}ͱ{֍�re�=L�봈n�>�<9��+;�׮��#JY�4��NT��oEb��«��٨��t(�VV�D:��s6ݫ/C5[��!n�5�O7���%T&�u��X��N�\ݝkN�f�����gv�'�O>}]\�iB��K)��y�;n�g<�5q��� �"��b���kD`)�SI1�TJ����F���h�B��KZKs
����d�hֲ�ZJ���Ř"�*�U�`��-`,�RTU��R�ڱI���Յ@�(�֥y*ͬ�;�O;�]݉#J�̑n���̹<�٬Y+M���L�����*��:�O��9C�s�C[�u�x�}��WԎ/<�懣)�ׄ�ǵQ����Z�ׯ����&�G���$��S�a��)��Q�ӥ���bm��܅t��;n�t==G�ۨ�Hՠˮ>ɩ^q��!�����}o���x�7���X!�V���w��`��+8�N��Put��#�&cv�5��;D;��v,�O��  �s��4q�i��з���q2t�ۍN��<_ERo�}c���G�z^z)왡!�d�8��roY�4�δ�IP��o��o��5�9Sй�������y���[��+#��L����D �W�>5�F��q�9����'9�ūZ��
�/Ǫ	�	����鹅�G<����������uA�J�?J&e_�eU�с��K*YW�-�v:·�
�S�Y_3䒜w��[�ݩ�>ȉ��-�jБ)�����di��28�M�I�5�6�f������v����l�:\�]c���g�{�A�y��T!���*�r~`�Syݽ�豲�j�u[��uC�M�sC�u��G|�^�@	�~�t�wxo��+�1:=�Fv���&��qՕ�Ӌx�rV���*rҶv爓)��7KrU�W|{n��y�G�wݞ.\�u��Xa�g�ɣH��S�x�L�7["�>�Å�/s�T^Oq]C��߭�Ƣ��K=���K��r�^v�N�ZֲGvp���zv7I՞�q��\�}'��%�zT�P�,��1똲P�l;S�ў���Z���Z�&5`�=�5�t�d"��c�#��}x�e�8u�zHr��^��l��'�l��W���Bwס^{ܣ��=Cq���'_Nig��xx
П���
�:�S(%�2:Ub�f x��uW�t[������ٚ�����\9_v7�n���5�{�+�*)9X����C�rfm�ԟ�b��#5ϊ���/VY3[:�%�F���;�:Y��Ԛ�@܉fw���P5���l��Ȳ�Uy��KT�J�##��رi��ו*�׺�!��W�:u��'on��#���v���a�t�5�13�,��"��0�5�{rj�5�F�����oI��ۖ���CG�.��Z�7�nv��Z���)O���Ё�򝽃Z�ol ��Qp
���L���h,`$�p����빧��X}��\�������~��? ����ʕ�����Ё I�>����񅝄	G�u�����X˲���&m�����o�]�J��a �bI	���|�`��V�v�����g��߷!6�K�����@$	?X�}�(v�����ǻ�_���3���\�7������Y֡��q�Ex���qߥ�9��ف��s��5�a@��!��?���~��H��	O��BB@������a������ʇ�?�O����鲟��ο��������g� i�~!@�����O��b���g�:&7�L�}�����7�~��K�:�[�g�����~���O�_vO���\�����<$	����o�_�����@�'�p>�;��d:�����\���l�>&����G������#��	���5쟰�5
����4��C�v{~O�xk�y�d���?�<�3����@�d�����=�}P���}���xpj��=�|.O$�Y�O��߿��}d���>l�\�t�۞�y�������	Ot��1����$Y��i��:�nu���
y�?�:Oi!$	7�h@�$����'N�{���|0��|���G&='�8?�$	 I�p{�ğ�2`��?�tOk�	$	�e&�D��|���5��g�A�+R�?c�s�d8���þM��X?�� Hw0>ϑ���d�|�@���}`(�}����a���'��<��?��������>���X��D0~�'���o���� ~���?a�k��� I�|�o�|���-,����A�R Id�6}��a��?C����g�������	��?��8�9�&B��濾D2L~��{Ro�'��z�7��c?_��W����:Ù߁�7��'�r I��ϑ���~_(9�V�!П�!D�w=� <�B{�{)�ϋ���h����>�A�H0! I�1$������S�~G�s���`B@��O��C�8{8���oq�Y:�>��vf�!�B} �Ĥ�o�d'����]��BC� ��