BZh91AY&SY�x/�[߀`q���#� ?���bD���  _  J      
            @@�   (       D���((��P��P��TQPR����T�EP�
�TE@)	@�P�PQ$���� ��PD��@	
P H%B���A@� ��H�� �(UD��(( HRT�
 �`i P)'�  P�T�0��j@��j�@��%UU��QU�����CT-j�d�C����  !J���
8   -sMjM5e��0(V�2���c V�FV(�B�%���L*��PCd���(4TT *��
*��C�   CZ��΁@�N4�:� KT��P�@ �1`� &ƀ:(-S�U
 v��@ :*�4:UP��"�(�@H(�   &��P.'v�
 .K� 	��
���  tw:+�4�U
�� ��;�
3Z%F�P�U�EB�!Ax   mz���w5A�h��V�-Gp� (���@�N�U)љ3@ �i�n�(�$��� c+ 4*�( R�R �Tx   ��6+5�T)50 4��J
�j� ,Vhm `�(Q� ��  )eXV�� i��THP(� �E^   ���CiEm��m
� 6E��d*�1`Q��bb�@4` Q�b`
i@XV@j���%UF�T QA% 
$�  s�UU)����TєUU5����k�@�F j�3(���0(H�	Q��� P
$*J�8  ��TP,@U��U%(���TU��J��Z���J�U14����B�ԠmQI 
�
�UEU�  ��V�S@�a� U��P*Ԙ�m��*Ab��Pګ(�cI���Y,h��{�D�@�  �<	�T�P 4   h S���%Q�� �F���0	�2 	�`  D�AIIQ�1 0	�i�L�"P&B@�M���S#� ��S�)*z�SE22 dbhɠё�����t������"�~��a~�֒�p.���H{��q�)|�65y�[mt EEu��@U��
�J���cr*���商��>C�<����?�r!� "����$��U�H�1�>�������+�)�@� (DZJ�Ӯ�.�Ӫ���+�N��:�����.�N�Ӻ�N�.����:�Ӯ�;����:�Ӯ�:�Ӻ�*�;�ӻ�N��ӻ�N��:�K���J�Ӯ�.�J�K�Ӯ�;����+�J�ӻ��;��������.�J�һ���*�;����:�ӻN����K����亻�����:��N�듫��K���Ӯ�Ҫ�Ӫ�.��N���N������*�Ӫ�.����һ��J��ӫ��K��;���NN���ҫ���Ӯ��J��;����:��Ӯ��:����Ӻ�����*��N��껫K���+�Ү���;��봮�.�Ӥ��:�N����;����.���.�J�Ӻ�;����;�Ӯ�$��;���(Eb}�{_��!x�ն+\O_�I-t�Fv�P����tF`4�Ea�l\
ak@{<*�tt�ӗpb�F.�$��Ѽ�YmU���6�d��6�� �n�n�6�ٹR�u`�y�m�K�V[��Yb��43"f����ڷ9w�`M���ƭ]?ih(T���c�AR���!{��Q]9H��V�&�%���N��sj��ܹ��7�s6���H��$���w#5V�w,!f���lP�sK�oƚ�Y+a������Z�ڊņ�^�ڔ�(������K/P�ԉ�%����krH�S���ѩ
�sj�VL��S#�a�j#q]�[�nXO*�;n՛���ݷfb�pDXZc�଻x�e챘��{�U��R�+^�q@���S�N��r��t���5��悛�{W�ᣉ��,{d�s�Y����@I�N`ؙY������t�yy"�2�T��/n�#6�
 ����rL��'��[(�-]Q+4�J	[`����5��h�q�ͬERR�XՠCj�XG���N�QE��]�N�-5�k�n�4��	�ڔ&�	�QB�%��ި���P��-V�&�	�������	�%m7�4;�������BU�ʘ1�j�#x�T�a��Z@���[Y��EQ	l避b�T��̈́��z�K�e���QGRJ��J�!q��Ra�t쑥��;Y7/H�[y�Y�Ȕ�X��t�rY�yfM;N��QS����tw�;sB7����{]d��Kc71��{�Z�a�w�]↊�M�� ʺ�{�f��3�h+��fԻT���A���E�����^��݊����@n�巠�4)=!����c��,�������~����Ϋ�����<�g+\��򞑉L��!�z��B�eX �-�tb�Nʫ�R�8��$��&�'�����cr=dǗ�P:M�"��-�+.�t�ɔ���FfP����.��s2I
�Q��U��4��9�s4V�-�Ô@�n��C/5��n
&Ay��ٵ����&��T���,k+f�6�,$��oC����ٚelCr�̭�XsN��)����^���U�N�P6��Ud(�-Y����6�m%1ٙ�5��ۡx�v%�w.8�7����D����"�e-InȦe�ʷ��ovV�'��
ܬ�T�]�Nnk�7+J�F���[*k�P(ǂ�+M����:�����CI��l݈�͈-�Aq����H�v�f�:rXrn��͍��<z�V�h�I:���NI1i��t�2<��M���1�VQ��p:˼!7+f�
�Ғ��t ͣ��]h�4Fm 5k#R����5N�-��@[ ��^ݚ��JB���8���ƙ��h��6J"��%�̘�2.�,#;R��&Sg�*×�U�,,yx�棭�cǺ=�H$D���n�+Xa��2�[�#��
G`7�@F��&2�J�6I�M,���j�����^����[�c�Ea�:��g5��Y��7���,��� �6M�n��j���oX$�����z�-�.=N�m^�͠�i+)MD"��)�f���0=��i�F�����]ɵ �#��$8��ٻGseh��z֝)�R�6�������D*0���ksM�ȳYڗ�^�=1n혃
,H* ,[3M&^C�3(G��+Ǥ�U���T�Z���@�@�w*
>���`�v������{�����V��Na{K*�F:M��d�������4�N�)���l#��~�-d%�v�LR	�*	��CTe��1y�n��f�։�#N�[4���(�b&�c��TDQqSRFhM���d6��8R�S9{w�j��Z�l��z�OY�Q案Z&�'�b��R���h��;y��yW&9�2N�`�����뼱r��[���e(ҽ�d��L1spX�G���J��b��T�f�b��qT�;���#�[�����V;&%W�F�l*�QY�������zE��O͚`�7F͵-P7X��ɑd�t�x"�M'���Gm\���z���gP��;�
�O��	ǩn'VtE/JX�j��wc��6���ًNOE..�ҵ��;������&�rR���:��E��u4�s,ԚSw6�M�+�{�L����ջ;�vwXh
���{���¡
�R��f���┬ݨ*�n��w.+{Z��@/!�gs&嫢n�WJ��]f����Y�t�L����Vرy���ZZ�  X�3c��!,��K��$-�if��W!�N��̢�H[�qP�Y��b�Ƚ�[���^�B��G������]<�ց"w����f���]�y1��#N]���*�c�q��3a��Vc�p���7`TǵXc�2�+^�2�rջ�H�jefj76�������c�+G�w�w�k6�����A�6��+J��I�Tia��0��!��4����H+5�l ��Gn��6�˽�,�Mmʘ��B��.�2Ե�V�El�Xkle�<��J�*�mj7m��6���*�F�7l)�/ ;f�t5]+�c#�Qg6Rjd�2����Рإ�sh��^*тd�3f�B����Ô!�ܘ鶆�����B����u6ާU�*f7OTA)!�ݲ������,��^�:#蝙{Ym����t���b��ڊ�BX�M�uB���B4+$��J�;[iYVFލ��+����vV�.�#�	ne=�%�ݛ�:���3��f�S�]��A/7Ѕ�(;������`��ŅX;�bR���U�X��m�I7ux�+*Mkpz�cJ�h;��(&n�ݳ5Ķ�VR={�S]kY�M��SÄZN�[8��t�5���,FB�
��]�*�� ����V��lӶE-DU�+1���w�hYd���nL��Y⪕�����C�rs]Jʌ�4i�%�Cf;�®��Vl��9��IP��x��ӌ��E؛��"N@�ct���
�Z��@�yp�[]<���s%	o�!Gu/M[&�*,�sF�\C2�4�����#����X�%�̲h$)d0G��:��f�ޓI��n$����qiՐ�f��uk��2T)�����{���ݘ�%�⣎�S[ ̱a�r⬰�9Nͷf�J��Z�j�t�F��u
4,Y����w�+k��b��*a!�@ѶAGU�b�m��6Z4%-����5�3ٚ4���9���YSV��m��t�kj��WXe�)b�B��%�-`�:�kw�A�ENX���6�U�Tmn�쮐(n�S -^;���3q=�)j��{wf��!@�{qک�v������ۊ���-�i^;V�P���n��з{�$�0�O�S�sl�"x��]��)�!U��tiU���莥�"��74cT�73sC�ŌʘUr��!�y����^eZJ���<8V�O^<�V��lم�{GX�ָ�'VYv�Dfԉ�m�Uo5�f�h�,fQ����~4�b�U��kM��RƄkmn�V��i��ԣ�s
�����[�udmlefnL*�	Rj�v���մ$�h�r��
פZB�`�)��ꦦ�H�Gȯ1czX9wZ�[��{�p����eL��X:&�m�X��f�����{�m@�/Iq�t��r�(�5;!7������u��-5��b��E��×X��sqbu�����ؤ�aZ��"�͛�uJ�v��P�͕�NT��ĖTXf����o,*1P͓P��^��"k1l3+U����ɏ2�Ĵ��҅���ݭ�b�gF�3�܉RWyZ�]�E,��FC�E�e9ofT��
ҝ�ۤ���X�=�*��%�G�Ѡ�Xt�1�ca&U��aV%g!{�M�P�n,E)����X�f��%Mw�	
��;5k&ͳk`,����"x�Z��:������[�ց���Z���!�ĩ��dH%���lH6��&�Y[Y�	�'/<
�^MÕ�Gm0j9v�������ɢ��u�^޽ZU~Wu�W&I���-^��FigR:�����Tle�Q��og"6��8cn��­��`&�ȍ��ݛh�*ʒ�HVt�ZQ\Ӊ\u���e������R�e�om�Gr�T��YX-�b���:��D6�!IV37&��K9EU�a6sKT������.1�i�1e�ͩC+x�Y��$>ũ�-͡��v�E�Ѩ	tB��ܗ�f�=j�o)ӎ��+N�����5`_U�"�
�BI�i
�t�C�1xQy�!���R"@����4,y���A�\/#2�r�]�k2��h�Kvni4P{BP�wd!�E�`ih�OE�Z3.Ь�Zԉ,��E/eլˏʯYJ��{�挹��ѻ����r��Ɲ�sF�:f��X�HB�aӹ���%���!��K4n��kӫ.ܮEO(�1�weۓ��5���я2�M˔�N৷rZ�F�3(Zݻ����z��Y��{���V�[��n:
�R�VX�T��n��:B�rÃ�Ȯ�����҉[.�Ջhi{�Cv2��/mK���2�+ob��Ff/"��@B ��9m�kT����n�T�ն<P�^�M;�Cf��S׵��+ ʽ������U�e�Z�KՎ�;bSk:j��yvsDEU��X���,��3rm^=SSB��dS ��`��#�0����w�r�!F	�Y���7e\�TWG�}w���:v��Y2�k$Y�n����fE���j�� W-U�e_N7Gg�o��,V܀'������I����KeCHM�#�L�nz��%M��R��۔Ҷx���L��IA+pJ�)���E�!�qr���1�ncR�"vLH�o݀�Ǭ��Ӌ2�c+��vf��\ˡNf�h˖b��d*�մl7�-W�����m�;Bn�L�r6u���ڴ�&:��Mf9X���̎�o%X�J�;L䬡RRZ�^�"�F�M^g9�p��j��1H�
43.��D����d�������i��̽c��[{���v̔�ⱇ�H�c�a�<����hnƱ[%Kd,iJ���7�"i��E�bZ�{\5�*�s6�eB�y�f�f�(a����n����ܤ�zwe�U�0Qv��d��yc�y�#�t�z�rj��  tC�ͥ�U�MY�6���Ƕr�S.��
�$G�n��D�i �SR�փ��OL'C�/F�d�`f���f*�kF�&�]�TPw3����j��Ch ɒ�ڽWRP�S�"i[�� �Hf�����f;z����{#��e���ը՜jBJWk0�+F�6ojGkQKq�e䷕�m)F�Xt�i�M�u�q�q!�@hd"�ѳ)����Ʊۘ6ɧ�ѱ�����,��ԃ�)�P��zH6�V^H��QJ��)�ӠXm��:4��W��޼b=ӑ%�Ș{ԕ�a:#y���i�.��{tì�E���Z3���U3�P��)PV͊��
���P$d�Lb�CF�K�v��`k]��5"
�Ǹ�[�U�aV���
�h��tf�F��j�"��6�+��aa6���w0�"x�o�s0�'����� �:��X����)Y���a����V�[�,i��"e!�i5��n���a�#<�ZYMn�]`�tN���h0����ĕ�@[VQ�&��I�X˃M@�ye�yb%�uK�M�4�R����8��ղ�"MA�f���V�nܸF�;̳5i�=�7QN�<zeDb�ˍK���m����bzj�`�u��V٧�p�)�m�ˋ3�d��,��Z,eV-�KU�����'r��H�ڴ��0%0�t^e2��r�5�F=KkAȱ�S.5q��ɦV�pk8�mk�S(7�P��6^�M%��u�R]]@�D��H�ܡ���b�x�%�хVU�f���Mm]��U�(�%�J/��	vA�9eEW���4cn�U�h�����6��S�L�{��&��KY8%���J��n�l�
�U�ԇFrè�#a��%�V�wBsmM�È���x�kh/@�NF4e���ӫNI�$0&�YD2\j�u�!T�Ң�j�YR�[T���4D�;)ػ[�AQ�`k�q��ov�c��^�5�3V�h�қ�w��Y�J�]Օ�O4�+.�:��f#��n/[�/�.$r�V<!0�wc̀ԩ~h����1LL(�RFLZ����C�ov;�V$�ԽQǓ�_����Y(B�k�^���!��g.IY��+3�"#��=y*��M��R�+L���(
@Vn&#o1�i�nۓ���cˬ�]"���
X8����w{h�=�l�(,�dA��Kv�&@�5�n-��H��[Zu���M�I�U��[i1�ַv��Tu��t۬-���4�^D�lw7XC��B'gXt��dъ+*��2�)�.b��ґ�U`�&�KNS�v��T�\k6�A(ȍc�����&�56�j�U!��ubyn���F��;u,�r�$��Uޜ	��ј�����mk�f�L��9��VW���h�Þ��vP2����t�z�I��T
6q�^�[<(,"�Q�cqm�l���Ѹ�O�%�	ZٛknL���Q	-�{K(�x��c��e ����z7$lc��U��e2�Fދ�@F��Z�Yn��o[���6V1p1����ܱ�D^��r��[M�Y��V��j���cn�Z���Э�ej���<*�ր�+�:푍d%��K�b�D�DC&��I���D�)9/j�mI�m��.]�t�hQ4[v�'W�vb��A,y)��f�xB�{�d���wI!ݢ6V'k-�Ae*̫AT�Z��Df���]����|nҙĖ����t�!Z������V�t\i��Kq�Z��{cT�*��sq]bȬ�@�ُ�)�J�T�Ո�ZiB	%�c-��T�;�5����]�ٚD3��+h���v������^��T�����:���?��d�O�Fo���{��B�������ر�-gr�ݒ���@g((oomj��Ѯ݊�3�6�ĝ5*����(��/(^e�C�k�Xّ5gd��*6m�vXt ����4�8��4�dҽ��:�ܵ����X"�Z�̹m)N븪h�F�;{֔�N�
v��W��Y��P5|sz���:��{�,v����7X�)�ͱ�F��9�3q�KK���xq�Ykg=�`�kVK��	M�1ە}T�̉49wn�V�K��4D��5����l��~̇�Mީ�:�e���;�p4�A^�us5v�e�2��Dȕ�~vH�r���:$LJ.9����1��E�f���|�DsN�u��u����gP�� ��WݗG')���[�t%��;@��G��G���O����6]��ki��&FN�s�b(e
���ih����OJ[�H���c�7z�iD���M;���v��{V'w�#U���=%�O2J�<6�h�ȺnNR�P��@.p���mi�}��*�V�X��Vm����93R���Hd[L�^�]E��T{�ۭ���Z���8ll����
�+7��{�e�V�3�91N5չ��\�¦���;�wQ5�
�-�u{C�Ge���]ث19�̫(�̑n�hW%�YW~��C;r�������j�SV�]�1Y�׍dWQ�:y����U�ĳS2��-q+�bÁ<	2\�����o������uy�V����K"���;�,n�ݗV�%`B=�ӆ��ں�Rd�zƼ��e�S;z���5P=J�ZC���$�7�����Tke���NHp���X��N�\D��WQ�Z]�[8���N��~��!�I�X�p�S�����,a/
bܐ���d��9
���24� 	��Wh�t���RN,ц��{����{�g2���ý�d͖;����(a�2�qA��3��\���36Q�;&���C2@jk���eu-�+m�˾�@`��I�z�'zm�H�Y�7�F���y����B�+�wP"�q��E��h��praچ����bҌ��*J�	@T�Sp.�2�f�뵬wnh3��A�I���	h���v��n��5s�r��012�o4��,�Dt+P	ٽ���>��2뎼�|6]�zplz�5<�8<�j���z� �:��yV�F���J%s�:蹝���Z�ra�{��3��&��k4[9�TsV��]��Z�g;S�VjuLB�S��:R-,f�Y��.i'����D#'D�.�D������X�(\��8M���ꆷtX�l����	´��ijo5�@#���B��@V�,ebg�ֶ�5n��Ω�������)kv+��uw���z�ٴ�����$J](��z^n��L]ID�u^��]�Zy�+�:e��W���u1_�Î��`R�t�q�6b�¡.a�4EV�̅���ՅTj����RfW9/���2����FJ'e�ӕ&f�͚Mgc�hjA�Npk�p����m2d�����zs���5�ms�5� (z�nߧX�k;����6ӱ8��P��	}v��ܻ�XQ���P�X�Ⱥ�l+$������$�W�	{9P|ҍEVYF݊g���l�n��w'�=��J�gZ��f`�ŉX{hC\<|�-5�������37�����.fD�1��n>N�G.Z*�7% ���=W�MISE��u�4f�Ý����1;x�a�R���@jl-`�kz����V��������׋2�HoGf�k�ͭ�k���}�봑[�u����Y�o+bYO����KE�6ܱ$��^��b�[�d7CGng=�Q�A�oN|�30��zɄ
k�(
|��Q��1�r��0J�CcЯ�Z�
�:$��.�-�Q`��{v�q��IW�X���)�`:iR	���P���7m�7n�LGWc[t4��+��d���n֚Ip�P,�VC)�]ۈ��H�|/�5"��ݪ���J_*:!�Y�o�y�D����+39�MG�^\h��pm�뽹⦪,P�,3k)��*M±UBƧ8#oXf�=x����5���w��D9UW�5�掻o&����Y��nVPT�y	Ɓ])��'j0�NT���(pU�W`]F�)���[�0�K��*�ID�4�����]]�^z�Z��r;sV��tJ�B�@YP-b���6N�+a�(����N��U�.�Yw�0��d���F�ET� ��_�Yp2�'��ε���/�"u���am�ѩhDǕ�g�t�I�FU�j�;{���/�2X'�qٚ*�J��e;T�^�W9���-�x4#���vط����ei2hU�x/$��P�5@�X�ҸDHS�"%ƣ6P6Gٕ%W�D�O}	�,�0VF�6%���7I`lc�ڽ��qJ�����a�
P����ȕ6zj�t��A �錱��Q��%}���ڳ_Ӭ���8�&\�f�j�=�tʪ
,-�X��u�����h��􋦲���X��ٺ��b�hl�4���e(���HL٩QrZ���޼�����8Fl*��ܢ�L3�N�d8o�����++vU�2�=����B�3{o��c�}��D�t�u�Xh��8��jn�tz��a�<��t���Q�j���fB��S2Z�(Cf�2־V8�YE;�7����jđJ�ْ���J*����t�t;�i �9
�o-U�I��v��+�������@K��Lm:��t�n�Q\]E�)Xٻ�эM���^Tvkg.b.�����N��XƳ�	b&*^���֤�s�Qr�p��A��v'ssf0H9$���� �׮]<�ùͺB��K�3���l�v}��N��bⓗZ�u�{mn ��b�����F��O-$�"���AC� ��ܬ1z� �kL�3�i�w2mn*�U��Ζ�������dgN��Y�d�뽧|�]̈p��+����#.�Rwp�];7]���Kj��9b�ʍ��ffj�I�GK���w= Z��(C}z"�넒H|�����_7Iݎ8l�}�o��.�֡o	 S�-�'sQ!��f�{;1M�����nm��z��%Fm�Ƚ��9Fb���_W'���x�5f�UR`�"��� �w�
�E1O���z�Qܾt*s��y9��'������n��4�3w �3�n�^jK*��2��,��b�[ղ
��DB�Bߴ
ԃy.�i�YrFb�i�Yl�%@& [�Ԥ�5��n���fU��ef�-ǯ�.C�w^'�a۝��u�q�&zqf��@��v�}��~�MK띖,m9�X����r�
�/�t�a3=�R�c��E�\n��vV�x�;�Υ��Ыgrh�;��Sg i��#<_����Z��+,Q=jQ�3�� {㸨Ҏ��� �yBg
�uO���>[ +���T�M��\l�ֲK ��]��[O2���Uل,�P�[��_"�ˡ��ٽT�k	�Ц��3*�8n��ݞ�w�ړ�<��|VP5y�Z�G[6ʙW#N��1X��֝�ۡ,���Wi\,��N�i�3{F�a��+<����mHrtp]�-ǔ��9G�mJ�Gu9z�b�F�d�{:��c�	rZ�i�kj��kܬ��Ͷ��J@33�Vl��eFi�VJ�R����X�V 7W��,��G�RuC��c�_P�ǯnh����C�|x7H�zt��0�5K.&9�����ډ�h_1��Ioe˩5\�ٌw".����'�+"|Mvs�w�G+U�����9��-FZ�9��C͆�s���4�ۼ�yu~#���54۩:�z�:5����C\rt�wu��w�:t���i��#9��B�kn�ꨶ��DX��gN:.��=a�Uk���qwW���X3\�ئ�������ܢۙ�0���{���ԗ6�]���k5��']!u�og�駪fgh Q`����]�.N��D1�z�0��rU�o���I�fS���J�L��K��R[[�@R����/˻d�����[2�<]����\ٍ�d���K��suV��1t�����wQYCN���]
HS��9huzZ���L�����f��e24�-I��:��`�{[�������2Q-�ק(xu�azfu�R+p��/��j������e��z�Jfh"��*��U֌z�4:��'�+�����ECj˄l^�p6mU�7��V�<B���9h^D�ɣ,�v�2�k\�͊K����/�I7\�Є�[i��܆A}��I��[���}��/�I�<�
ٷB�гy��K�������.=��vt,z���q4Qq�r�DO�
�
�.�����Y�V`�0v6i���i).��`�W�wҺo^^Q���Hosv��h=����δ�L�N�D&\'GPfPu�yh�QZ+�{3�n��{/O@���<]��\ν��N2��A���m�oY�v:�#!����DBUmJ����Z��w'lG@���v>X#�q�~%��E��y��̺\M����,SqIKξ�H��߳bC�j��Z�C\o8�E�UŪ��X��j���Ş_��;T���Le�Ǒ�[Y�^j�����o1�bô��[l�F��n�s_�����ON�X�����&q�I��h {&��79J�o��y�w%�wcJΎ٬feL��)'��ͱI]�)��\��S����9+�bx�`�:��]�5��<ٴ��kzo6�2���B���\V�f�GP��Zz�w.�P��L���⹧/2�w<�L'A�[G��0 �,��ʖKu;Bᅤ��(���űy�p���;��b��	h�T�ݙ�nvQ��9�"$��X�H(�s��E��M��� R=d� +,���Zj�B6�ou�[�)s�we@�Э]h^;L�:�v)<{�ug�j���7�k�i#��[ǩ�M1bj��!�F�����&�w-�"�Հ�.��>�T�7;�	��`��V�y[�a��[$�����m�R��f�yɋ��Ef����-�kgj�C����ht�H�#�����C������7��W������G��-�B	�i�R	`�F(���J�։˝{+�t�%�#c	�cwJ��l�7
�7Z����E@�Dg�T�U5J�>�֙��)@.�\���I;��L�7��:-�b��(�k�X����;|�^��JP�A�b�`F��.�qaa߅<�o[��&:���/��"��>2�'SZ��&hc3c���yM�Ww�a�é�@.ܱW�͹#�{8���Y�,Zd�[��-��ˋ{p�����eܒ������|B����u���F�>��E	��Ȩv��3��u6��؄^M1�9�a���M��씒@Z׀t��E���H��o9gC-iXx	�g�YxP,�Qպ<�npν���,��HP�W���ɐEm�Y^C�h�)�ɣY)�Jb̑�$Ә6�b��ˊ�:&
�۫L(.��T�Kݰ�Ar���7#0���h�䡷��u(b횺�f��]P�uɌ��p��v3�\�Ü�#���q��y���/se���C�5�a#�u��[�����^gL�ã=�G. �M�:�y>��5�>|�-o3���7`��7��h�;i�'܄�oN��κ���\�<���qE��d٭�T��I�����t-���L\xmi��&VD���;��t"j[ƳPԥK����;�z���K�v����N�`L�!��?"N�YN��T��ҬQ�j��Ҧ�wa;Okr��G�w���o1�q�kV�N�*��y])��<$Gqd���쮨�3���ve�r���S"mq4(��]LwUf<e�)�u���Pt�-mpʽu,� Kh�B ��^���V��.�l�BV��7����]w'l�	��)-*��j�vm��������Ѐ'f��m�45y��:9LN��՚RWD����<
�t�n^�ytWl��u2�xn�\�W�Y�4����xowdͪ��6�7��l��7�3q��Ktߛx����Kг=��&PLj.Ω���4����7g2
����F^���dԽ��L���z���^�z`=Q��j�����!.�(�n�ö�)��r�Xл��:�kâ��s%U����^.�/�.
P��kc�B��+0����2�l� ��!PH;I��mN�N/tKa�h�ь���Y`Ҳ�4E#�CQ�^-X�Ј��i�{*�ޣ�r��G΅X�s��]���TB�uU{w}�Ɩ���H��	���z�rŸ
�h���H�v��^�4r�b���o*�T�ދ:�,ؑ��nA�i��k��x0==z��c��lV�J���<<�	��+b��cl��g��Oa����}��B�C�-$մ0m��cz吨�2:raV���e�_L����z�]�X�+�;m�{:d6�j��^�#�A�yMCUH�L�tgf�7"�K��%���S�H��4�7��E��̠�z2�(ȴ��pԑuR4F��@�Z%�e��d,��r��÷V����`"_-ck��fJ�C;�-ɮ�W�oasWp׻u{�1]��Y�R�I�P�T�û�B��FkQ�̨���o͘��e֪�� �X!Q5��oZ��q�J�b#T��s/�4[X`�M&
)'&p�X���v�Vnz�v6��ெJ���)�y�[ò�"'�-��f���%v-+j�� 1s���\6�y�#�v�^f�v�XE�ɓ��g6��µ�̀���
ʩ�"'4���Ĳ����e�m�'\���e�v��rț��}ˇwվCR��ө�A��׹�h��i�ö��7{1a�R���.74��]B�ZT^�Q5z�����\�4���f�v_s�l�;B��{T�����NVrj�q�t���/k��U�ݮ9�NK��
TeR���t����5ab��u�3X����E��R�Pˤ��L"�:�Ȣ�>,�5)@EsJ%Ν\hi�AR���J�F	N�����)hJX�7��0�J&�a�!<��r�e+Y�* �C��U  îzqq�i�8Q|?��>'O7W_���-N���;�3���(��q�Ύ±_P'9�r훏k7o��x��X�����j�-fQ�S������QcP���fFR�O����c�u˭�Wg�����}�ܣ�R�SƎu��F��c�yrꐆU�l��DʃDeYYb<�^m�9dI#*���+e��-�n&�F�������^f,�ܴ���VJ��'���3J)	G���/|���-)���'M�ǛS����=��� ���{�xQ��Šj����܋G*�f��Yt
�W
'^���TNjM�U�rR�Tw:RwUam�T��Ӣ�at�^ ]�C��&�㢈����B���n�:7tq��Ԟ<:N4�-�*�u"wME)����N[]��Ɣ]Շ4丒��b��t���-F��PhT6t $=GZ:k	�^�ػej��zI�_��r�
713ZJ��"�CS�Z�;M���*�c�ͼ����F�	gs���%ꈈ8M�v�Ʊ�V�@o�ܸV���iӹ��A��7��[�s�' ��������#�x�V9W�a�,��.T�r�1>QÃՀ/ט{�J�ĉ��X�1(ח5]۝��4
�<�}C�e�oh���I{�VՕ�v��s
!�2�Y�Fe�����ں�o�ݷD��w�Y֝����3j��C���n�`b�س���K�knn����kQ�$��A�D�a���	X#AAA � � � �(F4h���AG�H � � �#�WWVR���V9�Q=��3]���B��B3V�l��wui-�;p�"��gz���p�w�%tuuԞ\oNniv�8��<�ܙ�N=ԑ,֭̀l�ևj۔x:�:���d��w�,V肭\�㸲�-P`16�^���synE�e���c�GB���$��l:!]RZvIڷ��3xh#q0i�+�{*]����l�+�b���0d�/"4�j7*WL]A\=��a�*�l������ќ��lO���`1�H���0>V#Ӌw�L��I�h,p�b�V�a=˙()��9M�LՆ�f,�#0�u3�ֺ����Ę:R���	i۝ö�o`A�1W?]�fs�v�^��D�/!�^R�b�W�ه�v�7f�]ոq���(���ܒG�nі�_Y�f+�W�@3�}���*�mV曣��tm���f��q�c�D3��{
�c���eq;�R�=��3�A�y�G���֖p���͒�nf%](�B��N���8�P��H]�K��X�N]i��η��V��&Jיp]YMY�z���=������3A�-��.nV�i �� ��3۶�<on���PKF��׎��{��^5��mn_2�h��,m�M�����(�	�	ڴ��s��Z��o>4*a�3(lΜ"ἊT�X�������MЙ�GDL����Ǉ��2_f�	/�vS;� �؀ځg�0`���8@! ��AAG AF0`�A � �8AA �A��2��*Ѩ�T�6a�A���
ѐ�� 
#чD��p�8�t��#r�ͳ�̴�� ǵvl�r�^�4�+�,��� �s.��A���$ؤn��(kyԩ;u35U��	�b���5����U��Lb�Bj�3XCD�@s�ۼ��f��)h���z%����6�F�oT���5ia�N���hTp̓���ћx���It����έ<3��+��Z^i��yX���dV�b�Yt��]����٘��|�
S̝l��l}S^��#`G2z�}\ή͛g��۳k�n��zDy�#.^ŗPn�av�mʊ N�����o�k&!ȪN�Y.��������5�q���8�h�z ٌ���4un��T�f���m�p �x0�Bz��.������>�iM�`�d]�P�0w6�)�J�٢��U��ZM�rr�+��{W׼���D����&
oV�eu8OK'rѰ7�m��R�ؐ2��в�]�X)�b��z������gk2p���DS��a��ݤ�ʁU�Cf'�u�1fX�J��l�s�*�vn{k�e�4�hPsWt7�M��.�����s��4�WH�3���F0'(��nI��*R�Z��N�ߟn��'RC���c�>�lp��LNd@ol��2�
]rA���g�2jL��r�8��kF���/�̈���8�oVZ�.:�]囯 �n�H�9��v���}x�SY��u�rc��@r�p*a��ory�f!I���7t���`�v�@��V�N�۹<1_��2ŞYR�V<��)L�Sk���e`���E��d���YT��7�1.��@Z�FqhǕAٮ��φ�T�U�f�r�ڃD��y�Eu������n�L��:7��'uf��������<uyz��=GMqێE�@3z�<�D�BYFٽŨ���ƹ7���3[��ee
F���ɹ�4���!�	�f����4#��1��w�b޶Vf�\�n�k^�d��tZ�ozdW.�jd֮���[9�-�K��Ѣ�p��'b�N����V�$ 9H���.�<.F��Kh��VͽWF�T��k��7{��!���vM�d����˕f�[��;Vh$�h�L�f��z��:<���;���[7q˽A��m^lV0�U'MA�R�H-/n⚨��wRAF)U����7W:�T�	ܣ��o�M�4������sV�r4�Ut�V��V�y��Y�^Q�Jm!{����a�}��;������b�EV`nʹ�%�%�+9����R�e����L���J��tU!��ª[ߴ����m�&3 c"I)d�ӂ��f�[�)oJ��q���d`��n���k5�.�)A�"D4�v��&X�s%�yo2"�Y2.�ent/�xk��y ��)N��f�����b��ӣF��|]fLT��6�U�� �Z�h�O,�������Be�w`�s�Ѷk�t����YQ&��T�e��I�+[�l�ɻNC�V�QB��m҆�2�[�}y�R+0�<6�|��o}$Uڰ�E���&������6�����a�Ĭ��N�9�%�)��ޑ�˧�g块@��sH�dj��]Y�kZs%*�򘉊�J0Ü�fJ(J� <+ؘ�4U��Q�]7����˾NΠ/��[�.Lg����rQvR��Z�<��k��ݲ�O @��W[4]�0M��yt�"R�UJVL��;���J�G���w׬Hx�^9�g!�0dm���7Yj�3�E����C.	ų"�6D�k��A�^Ǚof����V�PlJ�;�r�U�G\�۲Y��9�ԛUe3A낌�@e�O,etr�Bӫʝ���4�h�8^*�FApR�hc7�:N]?������92�j]JZ�Ĭ7r/f�V<a�������%u�p�vɘn�/��ܬk|Ugo���E[4��e��Uy��l�[������BFҰx;!�x���Ii��ܬ�����*m�61�U@�㽴i�ѹ�-�=�ۄ1���[��%�iB3�(���:�87����ٗ(p����ˋ�$��Y�+�C�fl�X+�)�]�GS���%�l]v����('sw�1����s]���
�.ܙ�Z�뙏:!� 	q;\u�3:[�bu=�1��v�R�z`\���`h�)^V��`e<�S��Џnœ\��(��������ǫ��j,KP��X�<�'屫c	�n�D�2n,6eλ��Ob�S]�G�N�)�0�T��+�p�U��k��m>�`t�w�G���]p��{:��X��}�&�Ǽ�3g'e�7J�Σ��2%�헧\�P�ʊ��vL�#�����=̺wW����y�^jfWTBZO��h���GV���F���:��\|=��y˵@��mӕ������oq#b����f�Jp74�	�kF
��h������,N$݆�@�9�wfo�d��=j�\N�_9��;�>+C��xY�K�7-����NU���;B�@�w�s.�gRiְ�1膥�e�^d{j���w�Yf�yv5��V;h��!g�M�b�rً)��m�F�5�x17���n��͎��(����=��
��7����w��WU�r��lU1�j/�pf�o8���W��{3@3�zn;��4Y�^TT�J�jr~i���뭸�u����5���(
 �K.͎�-�;p��`|�X6��Y����6֭��aKl�x���^�P�,7z>�2�86��+u�����}�����6��x]ͳ�>��C�s�m��{���Q��5��x(�b��-��s��u6����2������ި&�ݶ*P�xw\��Z�T��1l�"�м��v�匥�ru�n��t�{@e�q�=8,:�f[f�X��:�Hb�Mb��ջk*d-��&�n�S�k�����-�2��t:�t�/��$�[&��uH�M>�ı�t��l�@��v��r�X�LtkW�^�4��5�y+���;�o#�6a=y�|Vm��/en�Aᦎ�ƶ!yB1	�1E[x,d�s�/i�2U����	׽F��G� P[]�5�/��#tR����t���
�]���TU��h�y�|.��kfP,�۫��:!��vkQ�N�M	Ll��X�nҩ���l�V�6�(-痷�:�p�Rn��5�BaA��F��<٥&t� V�m��*I ��m��W�H#S��m#.a��:ivd��(E}�B�v#���+^f�5�*~M�є�{a����o7���Q3���#ۺ�E-8(�L�Rn�/��(�+/o3 �S�޽$���'!6�H��s}�`�&� �G�<b�����!�N�N���!֭	�H��M�c:��4�q �&�9g,�Y�B=}N�ͭ�
��v\�ֵ<��&�4�w�V�ep��U���r�iѕ&�e.��-�:���f�L�`�ω�9aP�t,��r��N��C`�Inbz{A}����ov�x���6���,����r�b-V��B�\��7�s�'��:�s�:�)?
�Ivr	����H�n�P�C~�ט8]��R�f	��=)��V��b�lA����o\�Y6=���@�vj�ځ�[hꔛ�yVx]ΐ�����{��<}��3�Hx�U�ʣb�q��!h� X�;[Z��3ci��jv'�usuW����S�Ιx�-̚�*1.���̈́�Ŗ�gTػwL�X��(y�v_a�{�Mv2�o��ĉ�r�켭Z�� � ���d�9vV6񒚸��[y�t6A6��ڗGr��Yc��Ĳ��K�X"�M��X�������;���fZ1>���n�iH������ccb����Ԫ�-ڴ��M��l=�;!��ܩkQ��]l���@j�����)ť���`i�MǪ��I{JgR�/fm�U9u�V�S5�C8t��L'�*fҕ%��l'�0⻤�p�7�вDb3CP3#3%�_ym*�}����i����%��[��;4s�/xI��.n	Փ���ʩ���i<�v<\����xF�Pe�U�%�؝W�V���$7O"R�a�vJ�H#�\N��j�#r�A|V�x���xt������hQT���j�Eܤ�Ӫq��EwטeJ- ��#Um�l�Ͳ�����Zx_obzȫ�;/%ثFS!	�f�n��kr�
�!B,�d6���WX����t��Yi�Q��;�8�"�k,�Aڈ���DV�\{��;c��Rq�VH��՚�M����8��X�z�GOz�ro���r�ИU+Uє��q܏�a�[D���4b؋uN��dN|ma����bL�|䵨�Y�,��d�z˫�X�SNQS�K�f�8(.�5�8�hdF»�E�a-\8�OgYy�jEf�S�h�YQ�U�}��7�p�=��� fj�3��D�/!νi��J*h�[5ȃ�No���^d���k�Ww���`�����Zbfb�B�%�o���GS]���3��Mm�t;ar�g����c�P�=����k�nB(�������\q'r�9���ˇ���dS�)"��U�[{oVv�X���Xc0E�Ε;��̲��ʲnm��
�Q�^�K ��cv3�nTN�1N��u�Wd�����n��R:��:�5Q�x{wp�bB����Џ��E�IBW*(e#�v���ʴ^�F5���Ln�yq�����G���l�u�P2͎�B��*^��f�[�Ix��Me�0�ZȓF����*���s�v.��r�!-���Z
P载p�e9�7zqEJ=�Z�wveN�ݚ,8l"��EN�eݳ-�$=�.���9ϸ�����C�S&+�S��R-T[m�Qi�ϏV^�'R{�$n�x�Y�ړ,E�6,�7fZ:2�k�CV��+1��S��.$�R|�N���W4��"��u�����: nFe�̃�(�A,ٙ���/@�[�*��tkpl4DL?��(�9��^������x�֋wu)��[xN�r���E
#�LR� ]�,�>�Y���@n�T6 ���V�f��\�"�̊N��8�V��:��!*��u.b�]8�T��4V^C�m	h�uշ�#�w�0�y
ĳ�3tv�!�P�y�Ѐ�I��t��9k-��U��vE˅�ɺ��d|n7ZV�)M3�L��[�0�[�@�4�qK���Z2uַ���G��`����/]�����ڒ`l��x*�!��@��y�F����l�[�%��n��jW�.��n�p�b�rpW�_[��i��z�ع�8��ZR�mɍ���6U�:�<"�45vV3˛�}��:�B��vfwWd{���U�`E�$خ�]$�k3H�i�Î�B���,b�jӽ�V�	�fiS�.�̏j`�ۛ�����w�\���}�g6��`@��Dj�DY7���Ƞ:���^������IZY.���\�8%v`=j�;���t��4�N�[�/br��6���N��o5иw��+�����nNk�s�I��5���ڨ`�r*�ޱA������8F�
�na�PIQ9V0Tf)�-�e��]U�E�kW�v�����T�_����|�7�;���<"X;go��|��1J��α���}��Z���/m!�`C���7\3L��Vf�'e�UG��X�Nm�Y�"��j�y;Ms�d������chsz*�2@�Sl�ν��hAb﯆�w )&��=�5q\�)�݁��kr���i��5ّ>i��ץ�W�[
�jӚ$[�+�:pК{�(!�ۊӂ�tTTlC4%�1Ðެ��=��c)����%����f��Ȉ��\_��:�!F�hL7BP(^)b5:�bd\(���aHwK��0ˤ�4�0�
��M(���b�����c7\��{�A��m�
y[��;��7����N�G{5��7��w[�e�`��.�E�de�=�a��PR鵙�I��)��������f`N�m��h�r�7tA��8Z��u7����zN�D�jw
��Rv��j���HТ��9Q��`[��}7��㕈�e!��(k� �x�f�;�w7��
6hB$}8���h=�Gz�B�v�]���"�-�(e��wq�ع،��9)�d^L���6�f�3�:�el\�ж�N��u�ݻ
��2�9XY,�	��ch�J�lk�"�wM蠝��l���V)�	$g�xG;�ײw{b�N����t�է�fo$QF��c�Xۭx�u�rbcaM�Ga7�K3,ڢ�ю��Z܌��*2۫��Ird*��+���н�ʹ�{�G��n���P:@��	�N��Ͽ�9�'�9���}�z)&��m��㓜�e�n3E6�)ȵ�����~�?m�Ő��m���#4cn�6ݜ�˵�Zmj�u�m�J��p��~�_���~�ƭ�ֲ�A6L�ͧ`�Ltf�Rvg������I(M��:,�-�I���3ǛZ3�m�톡�hY�i�m�	I��K٤�s�j4�m�28F�d�;6�c�HGm7g6�����ȣ�f��##r��f��j9vڇ{[�'$�x�kmm�$���ٳ�$��(=4����I8e��mY�c���$�ͭ:8Pm��#l�.%,�֜��8�vd��(H������fgB��J� r��3!�IDy�G6�瑛nJI������f�ŵFwm��k_�_�����~��7�_�"����l�/�sX�>��5u��gcP���st��V�oP����--�y�n������mP���r�ؽ�PG�"���[8i��a�� �{yOMC�8:u塓t��s�D���n�g̚���=�wvD>5��|��4N��t9��\���3�ЗPI=�Ȥ7b�;H�1z���`p�+�%q)+���a�x�ɬE�;��<ځV�%�B�=�k�u$��4���W��vt�����N�w����:�'v�A�H�F�]���E+�Rbb(ٍJ�񹵚��8�K�{�=��M����kL������Y��Ww;1�k[����Z}�q�����)M�%�`1���W)�
�*�s
���owU͆怲s��c+�H3|�X�c{e�)���3����T#1�I�0y��\m��D����މ��A�+b=��㉮]��_%�6�1�&.M�L��K^��aOGt��.ψ[���r�[�0� Q�����y/m���H�Xs/e��e��jŬ.�lȩi[�7hXs���M�\�s��\MJ��[%�X���\���חz���5�8�kedU�n�<6�v"G{5	��nd���]���:��A�XR�e7���HUfvKܤ��f��c���Ж�ǂ��hM{NX]`{��j<``�[Zr`�{w���l{���ǟBؗp�z6�.⯴l�H�&�h�=��g���.ou����C��1�ճf�l����� 3�l�J��,�G^��r��,:.��!'RKC� �2|���R��o���蜘����kj� �e��f_gЅ�]�3����w18�1�R�wU�f]r%�n^��W�������U{�[�qvpRj��OO�xS|����bc0����9�j0"�EwA���Jz:��NbwȑIkt,���ݝ�Ϸh��g�6j��p�v|��2Խ*r�A�]`���J��WŎ��ߏc��۴B��rU�2Ĥ=)m�1^����IA9�B��ևQW��^s�qk!�� X��Q�V�>®���i�����[���� ����[�镶�ىԤ����06t��|ge3j-s�:>@u^���6�IU���rձVo�8�,���%���mըư�_�o���X~%<?��>�dl�}��b�	j��A��3.^�.j�i�����"zr8P��n��ʌ7��u7˩ \ʵ&�J���9�ܴ�q낄u@F�\��`ďP:��z��WW̌�m�*�� ���&�d��vL����0��ry1v�ǎ��+���{K[N���� ���c9mÁ��6~�
��<��<�'G*����mqǭ�<���|��k:F��%ό(�B4�Pco�O��D�����<��+�/$r��⤯D#�'�IN�t\e�7CU���]Ll-����r�����Ġb
�=4|0�VI�}��jp���]<-����J��|�X���+
n2#�tb�?�9���OK��v�F��ÓP!_@���s7����И��V+ ���v��Y���7��B����6y\�Ѱň�4NrW�ܱIc�������|���!5�Jm�z�\��)#���W0�X�T���m�CS�"�C�^ڹ�gY?(��Nӫ��7f��6Q���µ���sM�ַ&��#��G���4	���,VG��w���K��<��z���*�ze�ᑕ������n �����b����Ƿlm�Q�� ���E{]�]�	�&��U�B�E���ة���;���k#v��u�͉�M��4&����l����y���tOE��wv��)Z�M���C�%dp�4����5rpZ�� K��}��(:*��D�}��w6�cA۰�� 5J�e/�m}$.��A��VuM�J��Ev���"��-��s��.�s��g�ԥ\����,Y�s׃��h��;;����iF�%,�=��c���f��b�BE�s����d�.n��|�YyqY�Y�ޭK���;�>��.��~��9f+��`����y'^�d.�˕p���ܾ>X�R����{�R&�GX��@�2���|˹��9w}��.��a�g!L�7<���9��|���{���#o[��n6o0���&�1s��tۚ1���=J�Q
K1����^:�e�ӳ5s�g��s�3��@�,�S�}�nU���H�c�oO��r�0�QX�QT�,5
�/l��ط�e�%k��6�7�(�L�M|tm{:�*j�^]����Æ���B�*$p�A�t��p��o�Md�cq�΅�����.�/+�ՐvU���us�⯆��|�L��*�_�.�Z@�������NC�7�o*�f�����;�f�}7��Er�O�p��yQ�q��	����%�_"+=���o�q:�	)��h�\
�խ�c����>��ޣX ���G8�1�3*
yO"I�r��:]����J�ÊȮI
4:��Ǐ��^��Ag��j�ؾGu�c.�f�R�m�v�O(�Hm���|}��j��A,�^Y�I]N��U1�j��oR<��_S!]��"�ڔ�؊"��<;Mu$������+^�t�a�����ǝ��lJ$d��zE6����� ��R쌙�
��R����xw3��uܳ���|>U�>����n8GT��	#����=J��g7�T�ȉ���Y)4ŭ5y9�1��Ny'U�����LlNN�`ь$�V\����hQ��̓e�T(
;Q���t�%7r-�Q��]H�ba���`���f*NK���A�Ѡb��DR��PUj�m�;?^A0a��kˌbZ�f�LK&3/Ae���x�Ζ]f�*��7��o�P��&+��a8��3�b����I��z�;����z�6X:���9,���{0�F�T��v.G��qۀ�� )���˨�UÓ\������ �c'r�ID7)�̏W��:�H���gZ �D.�S�vc�j]���	���2��vq-��%�*юwVCߎG,&��WnɽB�j�/!��(�!�����x�%ڹ��u���^j�{M�)gv9����5o-c�:���$�Hp�L��YHT�t;6�U3&8�_"e�0�Fޢ�s<I+��ϻ�F.s7�{�,����y(�o�����X����Yg�����a#�1O��C"�m=2�=�����휼�De݂��c��	�{�Y���T6�H�՞��(0\�(wFȊC�U��Ҙ����7�kwYԬ6��Ȃ�����]�9��ɳq�"wS��"d�#�U���m��.�b䢯��bd�mX�'�A����3`�i�P�x<�႙�{��u]
��C)�����}m/�#��õ�h�oz#sk�4M}���_��@����k�q�q��6WC��<9|ז|������޸Z/"E�Ӂ݆�]Nh�$X|J�� �D�J4Rߔ�Y�H�����ܕc�	4�*�2D_s��8>\�*��|1�dGlud+{�}؟X�X�y$������VM�p��s�R�=ё_B�z����Ma]6N.[�l�2�bjq�b\�Zm
n������\#��,�[���8�����;�T���:m�G|��Y1P���	���ry�k�n��9�x�B���{Zu�4�e+\���gó d�7ꊇ
�'qP>�,�s�9[�����o3�颺:�G��c�v��,�V�ȡ��@��`�,�v�Z�F�W�K,.��Q��9���^�U\1X�"&�Of6��[�Y]R�ᱰY��ij��#U��
���T�Uǖn�J������\tp\Ӝ�S�̻=-�80!#������
��P2^3��W׎K�i���r	�!ݩ�Nn5e�T;C%F�	���p�f�a,�X/a˶�!Tm��efF�8dU±�*��L ��\6B�SGV_����`ޕX�!iGldsumF�Q�[��������n�2�H� �W4��{�{�wۺD��&3�t'�mǔ�q�]�.�2�OB;دid�Y��w���či�\�Sh��9z�:�и(�؜�G`��Y5�ň�d��=���z�r*0�$�ꮜ����`Ԃ�1Q��Ń�n�<�P���R�l;N��}_x:��HG��EX�]c������jQ�G�p�3٪øcl+W������=qG���"�j�),�%���U�@��:�i�Ҵh<��m�V���Q
��(�5���Z ��t��Ɍ�n���]wz���[X��#j�� ��tB��#�Ҏ)#:Ҥf{=*�pU�����[���u;���8�"���`WG*���%�3����q��7��*�+�P;���򀂜����s%�9�Vq���Rv�lþ��t�K�����jv�*c�N7�qTn/�JHY���t)L����f"�~7VᣝD�V����-�����g]��R�p6�q���"#Ld��5�t�"V���q�4^V�X��"Z���ǰ�Z,׾�ٯ���j��*�s �}1��FgpI��uo,�����	vv۰s�[0~�R�#Մ<Z.p +��'v�\Nw+}�6�T���]��H���b	�λ�ɮ�hӘ��j4���o���Xg"k�{�wE���3*pC66������6�&�>�ؕf��MA�������q0P3�v��Q#����y��Y�MUtB1�>[<js���`;����BPi���aX�o\v�״	I��-s�b7�e0bD;��5��`w`:(ND�kSy�t��c�}gPV�/�DP�b���uƃQc��aq6�F�,��#m�o1-vj�w⻓=��;�����;;y�q<����W<��k���t$���PO�6��v����gl_#���;՟eK͓z�Ӳ{صՅ�᭶�fTiӚ������n�H�'F܂¬��zo+O[�TE^��12,��6Euz7@Ϗlju�V�s8���U�p]�	�B���{�,�Sb��a�M�ֱ0��E:h����[<�i�Wmowf)��}Qɼ��젨������+�u���4����P�L�wCQ����ήkv� v	���.��Ϧ�v|���A������=��nAR�o�|�Gs쓫�7e���J��z���]V����2���x���@��[��{s�}ʱ�I�f&DLe}���vP�%
��y�%���:�r�e�ϵ�3�|�}˩du�W���[�Gvs�S	&d�a�����>9���y�,��|�]����5Iqv�)ڍ�CAe�MLKS�
����a��0��ǽ��������c{OB''�w�i�|P��d�c�aÚ����B��!ok���4�+}<�gokfʂGmt.��#l7�,8�k��*y��pcj މ2��u�7�~H���A�j������_W
5�}�T���U<p	��<C���،�lVcE:k.���% �fC(n��v���2v�&��ޏR�)\��5� f�9��uuB|:���b���Ee��-�p|��.�41]t跶v�|u�]\�C���XkU���S��W���A��������g6P�x�����J�+w�lfVcw�8 �6QY�P#�v�!2��r���3��a�\�Y��a��۵AX�v���F�F5�`��񕗜8�P��).ڲ�$�h�mJB]ҕLԽ?��H`�kYPjnk׈�B�;5�V{v�;�(=,�7�.�
�{]!�M���b��[ݖ���6�p�r��8�{�2�l�%�"������V&S���3�̶�#�2�v?f��lv�mh�7�Z�J�]z�����7Ϧ.���g;�(�U�Ar�Fk�ޝ{�Y�wNX��K%L�xsW��F���9L51�7�a�ZV(ʨ8�*�*�"���y�:��3ըI���4[�Vm��������+ʛG�泥�Hw���r#��𧛊�9�C8Y���I��.q7�Қ��n�s~wz�8�$F��B��U�6�u���=d�����b�6�����m�P�4��a��������x�F��P�F�^#S`Q��k,�o1,F�ѪDb�g1����Q����$Sa�.^,��B�d,����	.��6�k�#���N�o	ri�v��`Y��KF��ͪ��^Y۬����Y!�s�1��UZE��S̋�l��r�d3,ޱSmp�]�y٦1�i���u��������;��[�s)] �q�Z���h�����S�:�J�0�TV�JR�+7�u�{���,�]��]��J�wSK����]i� O]�NW�ّul����]Bpa� ��l�1�KY�P�r�`ȩ8n���w���J`.�����Zc.�B�r6AI,�y�0�ꗊ���t+)��/�ӻ���]k���{A$a<y
Wkݚ����U�j���n���e�m4�^��X2tY�js�Fl�h��ݚnm��T]e!4Yx b �N*�5r��j�b.c�6Wf'�ky�w�S+�6��][�����\m�hbi8u̡Eco�S��Y62-�M�՛wI�KT���i���=����L3��W�gu�`��-h ��Žob�%L�嫄]�8�f�:�r��E��������J�H{P������_f�
v���/fR�:]�j���A �0�27�*uĶ�5��uff�o)e��ڀPh�̳CnCP�t.�cY�_��WZ�I��}B��N�ͼ�� ~�,y���е��wiI��hR����*��I�S7B[��uud��P���f����uCx}�!��=�XN�
�`��;:����eFĲ�`"S���=ݩ��,Tn�/�|r��zKV��8��oh�)��
.�zwTW/��0��x�{��4�U�ók� -۬c���a���&C�9om~�F ����н�t����e�c��܀,��6f��d��,Ľw������g��m�l�j�yy�7��g3 V��p���$�6�{����X��/=��m������_����d嵝���������ڳ;����^�hr'��6�R6ѝ�w�n;������ڲ)<�2��9�Y���ۜw��H��vNgye�W�cmD^y8���ݒ3�:{#C[���ؽ��f\f�O4y�g�mآvٶs˴NC�ݳnQptY����Ӗ�n �fr$�2��ڱiV�n�� ��=�S�S����۴�m�I{i�km6�{�"�;�^���[fw��3Y"�ȱ�9/+9N�Ḩ[9m���t{Z+�5i�	f"vE�w�xG����>ݸ��|�;��B��n��e�+G	J:�h�i�˼��.M��_w�i.��}��7�����_�ϟ�������W��Y�Z�;�\��`�����2�3Ěp�iY�%mT�U!�S5ޏx��e���]N�S��/3������d�Ω'�X"���S�%M����K*/৆���UeI��O�͞���a��N(Z�3�����%ӕ�:�8��|	���p���.�ț׮c|���ʬ8kn{wz������B�]KC��_�
��T���Ϗ��02�Dv�[��w�
>u#���t�7K��W��հkE[�y3^6+D�>�W�D�[����V}W1���T�8�eiE����&|�ٽB3���vMh�}Z(�z=PD������8���st����߈���Wv.�����c�cup��M�C߭�q�UޟFq�,�_�6�=�'·�(~v��������+�qE��8j��sભ��v2j�d]�1�}[R����K���n봖>�. �ε�Gg�4c����iԄ8���ҫ��f�,oL9�C�G�}�s��{K(����W�����	1��dG����:;��5S�S����?9���=TiWl����z���~Vz��X���V]��6 W�;�!���@Ⱦ��ft� ��7B�������O�`w��s��xV؟k��]�v�7㷣�Et��R��)ձ6`�ړ;.��.u��\�r_A��2���Oo{B͙4ub���u]��W
� ֶ�m��B�26��I�:��#�:�gq�Z�e��$V��.���r�(5:���u��WW=�L�cnWIRǕtϠ�U�0����@�g�rW�9��,d Ĝ�F���\�=��5JZ���3��ɜ�fBWQ�J��� i�'�t3�w�����ɕW��C����U�*�}:7�v�U�1I�?Y�S��?p�0c��c�Iy�B�>���9I��<|�O[RCW��Ň؝b�d��:&DJ��z^���y�NA�y��LpS�b���h��ޓ���,q{m���07q,5J�`�B�-�t_�]��R��1��i\]P訹B�������b����Ȫ��X���O����cۤ�w�y�~��bnvT�	�2��+��k�NW�h;�KE3��-��o�L��J�ɉ����;m�~�H��H7\!F7�b1�~��P��<��s`�L��X��������RQ�����Q>��� ��Y���=��s��.f�ʏ�ў��Ј�á���3�'�yZ1������S�➝�7ΰ�1ӥV9z<�ځq�=��g*_a}�+ayOUL���"Q&.V*2+;��VA8��H�3"H��6!��D���Xf����%3�a"2��#��@��y��F�P��a��z�I$0]��(�����|�(sFZ㸄�D6�%��^�S8���*���S��P"�UQљ�J>�;���%s#�L���]q*Y��z�����"vj�70������E�nF���](����\�����lR�~��+<!���R��u�x}sE�+����?T'Iz��z���Xy���,]��4�=o�s�l�=B�W�a'���W*��.>ۙ��Cf�V�;��kލ�zm����4[�6;��7I�3bD�(1!��B	���WC3��{}�YL�<f���'�`홨������BϚ�󚙈���O��P�Gl�z[��8�WO�.�80Q�S���5��R�g�jߕZ�S�|��x���n����*�B�}�tM�F<���*9_���w��N�t]J�c�дy���(%�og~n���r��Z,����W�ި�)H�6�%�e��b�z6�	��}%�&6��gݗ�>=��\����K���Fr{P0��� ݽ>�!f��!�LwH��.±s$)�)����:�����A]�P
����B����=�S�^ɞU�wf\���+a�æ�h0�]�)�Sn}�(Ϲ	�]���Va�"�cf8X���LS���TAq��]�w�Zzƍ�x�*w�V�ˬϬ�7��m6�ַ����[ǹ(^���O���Z��Y�M��Sa�E��e�e�I�el�p]%�j�؜N��u/���3�����CQFin�!ll7Q3�!�^��Ǌ��T�&�%a!9�n�Z����d���,���v�R8L{�a�8���H�ۨ�8�u���>Uƽ�lMC^��~���}>�pM�Լ5�=�/���5|����{J����8�XW�f�<7lƽ�q���~�����?{ š�FD��~�2�
L�}K�ϳR�Ϫ|�u�4���v��"�ǹ�Cz/���|i�q�*Ç�з17�?m:����u�;v�i_t�/&�FN��0�b�E�^���>ϐ���b�|�a�z{.��:wÅ��+}��ǣ)��tW�ޞ�٧=�ϦhX��6*[신���AV����A��O{�y���]���~���ٚ�XX�d�i���t�>�=�{j�g^��":_����?yA;��x ��-�>�Si�r�hk-�~3Y>|���Q�Q�":hH��/��1�;�>~"}�����h����b�`ū�Ԍ�ON|�\�߂t�cy�?oިʊ�n�ƪ�ZM���Xw��@Jp+�_@���+�`�R���Q˗`������/4c�L�����Q�3c���`��i3lW*�K�ѣ����K���ک{�M�W]9��6���y�پ��f���s��:�[2P���}�7�eKX0XE>�ud��#�7�P�!΅{v#sQ�7sn�2�dL`23S��S 0�`�R��t�;�w%�*Nf�� R�O@ǽ�4��ɻލ��-�ȚT$1&����O]\s7j2�t�>�=۱C�hm�s����x���%�v�{j#� JAX���z)���^�u2�^	����j)|��kS��;�MOx��LB�����Ӆ]����B�Z"aXT"'�B�48SS1]>S}�x�c1@���~�\������Ae؈kԔ�!Wք�HP^�Ug�
�Q�0��W3A�P5Q�r��Y��=��r}U��k����uyiN��t���	wg�:�J���A�,�Q�'�U�'='�]����*���&N��y����u�yu����ޝ^㏌g��Ȋ��nol1�ڙ�na騨
�^ѳ�=ϲɦ}/�٨��n&��1qa�N,e�"���}雽�~�̡��>B�
]H��ɭ��z�2y��,���L�2��+�Br�X��?�8�y�*%�z��1^��ۡ��{!w#b��7 X\As�!�n���W��{ӛ9�Jpl�f�a���
�¨���΢�Z[}y;�Ή;;��b��RF�����=����Uw��c"\�'fl)q�3kz����8f��RfFK��g3K��}p�&�"�f�S[Ǧ�8��l�`�wV��Ъ`	�Mܤ"�\U\�Ȧi�Q�;b��B�^b��^<v��Ԉ�z"��9��7�R6��X�5L�N�T;��T�D!�,�ns�:��e>)��~���1ZT�u߽��'�!�ڕLE���Z�XB���&f���UX�����8��+�f2}[R���x*�W��i�q�7���B�"�j�����Є��Ԏ6�"Uc��g#{c�za��]n�-��I-x �sʓ?O����!����N;e���ъt.wQ�\��*�%�;Ⲽ*|�5�Ę��ŏzu��f�_�ؓ����L(u
��:X/%#�S�En���]���!~^��4��W8�eǦr|�&b�5�02�L�C����g�Юc�="�������k9��ݼ�n��9Q���̿���H���VH�
�����ԗ4$������VŸSp:ʇ+�^�� �*�}:����U�0):'�{R������55u������^2Lx̡71R��z��x$�]��[�5y���a�'X�>rFˌ��b�O�ϩw�<K"d;���½�
�]`�~�������6yc��Cw�a��q�ީ���L<w��M�N�/����^U���u���$���G�"���n_�_��|M�H왷EvT
3��(��c�N�`NO��d�#�a0�6�[������[�~�,�x�j�����Q�� �Ud隫(3���~�b~q�j'8wMp��b� ���Ó����Jg`ҳ�1�;��Wq�]�c�
�g��)d��÷:C�D�&*�X���}���h'�}s���ygL~~�A�+�����8f�igX�VWʩ�Ք�*jݏ��-С;Ⴢ�HF�铘������D��b7��0ڿD�� ��s`�L�؅c�����ex����cF�Ͷ�n��91��4���F|z�sѫ��8�B�6o�<��}�ʕ�"5��5A���ς~���>[���R�lea�����(υz��c���U�[�b��[Θ��#�N@M>�F�=W�>M&N6��ϛ�D���8���q�.��ϻ������|j�7:%U�{�o���H��a��o�ר�ΐ���/��ا��U�,_����"�]!z�� �]E�8��L�l8�� nU��Xe���,z3lb����-o�~Ϧ}�P/��0��&rO���]B�%�d��V�ˇ[�'����Y-��SmVCR��46\���7�F$��`BC3b�&{��tc�_���9��0�����1��P35[�W�M�'F}U��b�};"}���&��a��������V�������+��g�jߕZ��O�
��ه���3�PJ\��+��A��z����A,S]!s=��P=�JӀ�;�����wc��vOK�ޫ�C�A鸙�0��ӓvm�al8�C.�dfSR��+�‑gv�%��Vki+o�A��$	8n<Ⳬ�ʗYf�
̀����^�U��j)�-D�Ҷ�]H�����eDӝ�`��\��}�5��uYc�bXNA�\(��<9`�a�^����Fٝ�S��[��s�&S�w��/������ߧcD�gP$!_DHc�Ĉ��Q��P:�� �_��%�f�*T_��B�|��L��&|���ߺ�D�V.f�T&��NMWݲt��7/~'&Y�?{�cϽ�N<״�Uv(�&U��j �YWu��[�ȕ=2K�yM�۟@����'U&�n���^���<"W�3�_{ըM`&�Bq�Aj�<�'��\�:�/Q�Ke�"Ƣ'�{�G�q��wl*"�J,E+��j0/Sc~��j���@�q�9RЎ�P�!�kޥ�}��;}��;�lV@�D�"�~�k��F1!}�\^���1������uBu�C'a���C��$3����ˬ�yՑ5�B�z<*\}��B��s����.a�-Ǵa�����њ5�^��a��K����o�sӛ5U��Rꈐ� �>B,;1���q���*�纷�v��f5����v�8�M�����:{�Nsg�6 �ږ��]GG�����3�{bFd)Ȓ:s�,Bӭ��<p���5+j�닏j�y)��\�jv7:��f��|��+Py�N���_u�UN��.*T���/�;a��i�����%Jz��ڀM&�Mn�F�t�,c' �>�ƭi>	�zy���G��i��n_��B���'�L��wn��z&��z�V�k��x���p��0��$��j�{)o������li�r�kYmK�k!gϖTQ�Q�dGK��NŵϪ��~���7��Cc*!E�LS���>]��.�R3>��ԯN90��)_])EN�]v=,��<�Tߡ���3�$�
�P�.J�|;/��e�=F|�vҞ*�~�e篪¹��F�?29'K�|hoN;"h�"�`+�k�%��������a��t�ޛ�>�K�W~oGx����;2�t��N��Z�޸��V���@� К�*lT�K����N���e� \[�!�"�پ륱���_��(A��ʞ	_��®�g���,U�&�B�5�5�}��?y�L�u�H�>�vg2X�T99�b#��Ғ�HO$(/pߊ���d(â��W3�1�-��C��q��z+UE_X�[eIIX����@u8TؖĆ7P��?o��P9���u�j��|L��Y5D�T0��Ō��nt�oN�#�>1��Ȋ��p{a��*��z�B[}9�1�̎'�쨼l�l�:dR&V)�n�7��͉pR��[4.]1�LV�{���*6��W�i0L���L�;�"`]�7h�3���t/����ȄU�]�*�AC�n:3��[q�`����-��U��.�͒��շMNS�8b���z>�'K��;I�5Q^o�aV
��WZ)��\{/���Y�꬏2�Dr�
s�2)v�0v��@�����q%ul�K�'����6i᱓4<$l}B+�F�����S�⊪��cǸ꾜��:�z5�p���9�m_�g�;&�V���&����^Lx�R�7�jg§�X��8��{�Q��Aמ�j�r
���5W	�X�u�vzz5N��o'fT�`S�F�fc<�v�����spEӀO��}h� j��s�Un^�v2}�v�D�G� qI�dc���_�g[r��:�EQ�Dw].���/[��x�r�E.O8yw���D0�R#5ia�V׶`KTz"��K"b����
���DA �F)���5K�R���[K%r,�b�%ߧu���S�2�����
�lI���&&2;���9��3X6n�Vc\�=�h�����z��̡�nX*���Ϧv
�����D��@�f�L9*���WS^��f���PW)�����k=���*4���o�o��#%j�@רP��
�:"�ު��g{��]]���x�>�HE\���؍W>�7�]��U��x�:��wr���W1�ۭ��0���W������Z �R��2"f�Z�7��@�fA�i6Eo#\�kU�|<�]M͞хS���^�*]�Ճ�>;Ӻ�x-I��w���1�����9a��:�&)l-�60'R-4U^3��B�Q�'7Dx����*M7]�42�B�7@�d�kMԊ��fɹy.\�oU���2��z�
ٰ�uV�6�`�0B���U+�7��R
��r�M�[VcW��;E����l˻�3�4����0��v�vʝun�Н!]��ƹ]Y�5v�R,��+���SofJ<���X��X��3Ǜ�En�N�Q�γg�D�q,N%y��+��k����w�� ���M`+4J���R��l"���F&Wq�yǘW��4oYXi�e�W���7�m����j񥷳;�~#�{�a$���ި����r��.�i<me�vMX�Y$���z�j����.e�5}t�W�I�;fL�r��mv�yZ�]w���*��),d%���u�L�3���*0\1J�|�t��/�f�Λt��es
,S��s#M�Чy1��sU��ѬT�Pu/�p`�M��л�%�lB�w�6�X�n$f v���7��wc{����#�8=�����B��}T�O��WKr�A�L��-l8ov��RLc�Nb�7^��˳��{.oC����r��G��EN;{�D#B��U�2�{�|��X�e�.)��	�;���|!6�n�]��ք)'�w�����0�vt	��mkۻ���9u������Bm�:h鎮)vv��Z;L|m�f+ˉ�O�Ij�tU]9����\1ui�w�n^&��)mv4��5g.�;��N��N��Bj�{v
7l��������R�n��h(:5Ӥ��YKtj٧��V5ᇶ10�r�K{Q�����i�gp򕃷5�,�Y�V�#7e��&R�"0801�t����n�^˙�qf���n�k�Xemd�Ck&��dגڢ�u��>��5C���蓂8��Pq�뛌��5)IJCrF����br��z�T��e�R*����L��i��:N�!(�ÇK�Ř�e�Э��m�c{v.�@'������5�d:�3G-"��;�#���P�6M�8D������Li��ۖr*�f���eK9{�b�-W�MZfV�IU��3V���͘v���n��`�{YQ 5�ftH�ݨZ�rq��{�n�n����)ԛgz=�ks^�[d[u(ޥ�4�ߏ�q��C{�`�Tm\�M��������Wu��o;�t��P�GtAwM�I�*U$��cR0DL2�V�����NV��U�"�	�� �ճY2�aKܭ���c,���4V~���6�G:+�aTo[��)���ʉ˥3������s��{��N��/�)�egs�I��9�n� H����ǵ�S���>��ڊ�mQ�������~�9$����P�ml�q�D�b����v��!���s�kK�|�Z�~������<�)9!������㿙�.:';N$���:GAf qܳ9�{�A6�����or$���m��z�-�yy�ID�ݵ��O,���4���H�{זݨ��m�w�H�����#���x��J$'�'���оX��{F��prqYe����&�y4����[��=�N^`���[[�툍��k�X�ks��Q�J_kz�m��e��[ko����^�p�j��9ųn������Ӷ�s�0Ps�k�{��rI�ܭ"ӭӜ�c�z�������e��։��ydq���ﶇ>�^�ץ�n���7}��լ��s�o=�������n�|޲w��=���|���\t��n��X$^Y��(H�A���|�#ȶ�(���͐��6��Q�mnf!�X�8s�p>���nB�a�x:����ۍok�䶬�ܓqecF�;4eqR�=�]��j��
��$��fnT�KS�*�X5�unϡWC�ԍ���Z�1�):'�bf	mvm��z�8�y�������M)�q�9�eB�Ϗ,W[r���6,>NmGxP���Y�Y����\G�t���2���)��x*Qb���h���6 ��w�8�޹�������	{����`���l#*�4Ek��Kì\�1"���b�^[r������M�ُ�S���y�}P��(��
�����RU�0Ul!�s�ϣ\���N�,�3C�P�b�����S��*:��N�"�<��߳7{˘N���)�e�P�~�#j���~C�.mNL���=��剽�]��:q3�D{��2�ИgulwZ��#�i�=Ss�}c!=7�
���뜩J.;p�d^^߼������4�2����1���`�S2fX���X���{��P2<tt������~9\���G�z������~`]#����`���j�7;*��t������ok����r�^�=����kf�������+�t�C/�B|}sE��u;�nez��S�拪��+AټZP�6i���k;f ]�/��8Ntp^�D'Q:Y��X�%KS"x&9�_>?In�wMv���w��ĆA����Ztp�D���e�BH(����Y}yGs�a�P]@ej���a>����/_?����}������b�D�'rQ��ϠDD}�j�.��7�ǿ47���[*�2�϶jH��E��ٗ�A`��Y���;tpjm�/���&���Ḝ���5/�M�M������F$��`Hf_{_q ���=��}ЋS�6�4��~gϵ[3Q��m�o�څ�vT]LE�T�נ��Wr)�{�^����޸�a8��8fp�2�g�jߕZ��<P3��fh{�c�6)Na��j�s�Fnxԝy������"xI��8q���>9`�`<�k���H:#lΆ�)��|��xލ}Op�������/�	�}�vO�t��B|�`츇�{���*��(,N�w����{�^�vd��#9;�P�F�JtD�V.f�*_p����)�9S�W���b�.�͔�Ւ����'��@niLrW�s��-p�+I��4�>�&�i�BП)&�z�~5+���7��]�����ND
�ޭbk	����b,�Q��z7�٨Y򸙥�JZ�MzW/��f���`�f_��Ͼ̭��ߏS���M��ϗ��8��W�v�l��
�F��-��g�v����ym� �	�G7;i�	��u6�qvn=�r�NV:��4��,����D���������Z^h9�:&&��܇�`l	���]IF����;��Q2p�'{���!�ϩ*=yh��/��vH7Z��Yyz=�y��ض�^���#"BI-|��V��#3�;��D�`P�)H��~�j��nٍ[�ˍ�]�ӫ��o�bҹ"���;��	���|���{t�dր�(�_�ҋ�f9�Cu��F�����\�v������^��j��tcu�u�Qf?_�A�bU�+�V|i�G¤-�����>����CB�>�<=ٗ��A���<i@P鷃v�~���=��nwӳ4,H~��lO�oX؝���Q>,����w �1��qC�y������M\7/�����p0OV��T�xO��=����O�$]������xX���S�.�׭����.���j_�3Y�I�Q���tźX6�=�����,B�"z(�Q���XP�.�Zc�����/V�0��]ǌ6<s3SX�U���>:M=��aH��D���uTtX�+��ݗ�^���
3�˰n��*�y���X�Vj���O<��-)�c�8�^��p)�G�H�(�@��$K�8e�/�:v|�YY��ں�~N���Au���J]�-�S�<�Q���AZ+`R@+"t@1EM���qۜ1K�����`���ڤvD�u�V����g�u3��5��˽۝]b%�*�T�>{!W�:c7����B�THԞ�#6m%VrL�+ 3;�ڷ\H��,0�TJ�Aԅ8ӁQ�5��UX���C,��.*��b��R!�'��.l���P�����s.�g��P�@
�B}���DD G�/l�%:��Ң(ϑ���;x�l:9=�%_�����B�Z"aZ�$*�@���t2��Ϻu�f���KS�*�����:*�М	
�U�Z�Y
0詅[>��t�G�y�^��y2����DӭS������X!_vz���6%�!�ieAv��ǰ�|��%�:O<~���͚�dQ��=*=�]l7;��ޝ^�90O;����9����&�*�'���Z0}L`�JdK޽3�of��M���F., ��s��+A�7�U�f	��c��g+�5��(��ow�AJ�Bc]�����{��}�Lй�28h�������o�'��[��z��m�>����зJ���Z�-�����H�ٵ<==3@0hx�ʾW7F�{B�����V�]�8���f8�0�aUp��ɻ�{mc��V���Bk��� ����=�षʫ��[*��G�K����XB���8j��r�i�\�d,���6$�ݛB�l皿�'�vi��J��F~ߨ:�رI�G`�!�ˮ`;��E�8�6�<�:b�r����^ݯ�X�/9�X�%�ǻ�p�ז��L�Ky՜{x{�=�x����p=�Ip�C��kr[ܻ�5f�g����"�ݕyn�H�#�P�����u�֐��	��n]�b��"�X����F�z�")-��g;+�[�*�k�Hl���{�<(x�"#� G� |��x�d�o�X��f��ה��W��N���W�%
��(���ص)s��P���m]q�S7�����{;ޞ#7�,�T��֩k�9���2��o U��I��
�b�*P2/���{B���u	ϧ�^V�'��w�M�߼��:��σ�L�73tL
��A\	&H�^�9�k/ҧ��:���[�7�d��2+Y��m�Q�򵳚����.#�:�f#���;����{K<����pbs�b�&����cV��H~�|ڿ�����~�l���
g#�}����'C�ۘ�OD�*h=S�0����]��A���Ň��yU/	�����Da��m�fH�Q�tL� �D�p�11�NF��~��C��h��G�Z��{|A˕���ǫ5l�;Ɇ���*�k�j�3{4��\�$TP�b��ۖrĽ�yX���l
�{r����r�숬;fcw�b3���lz1ό��,�3C�P�'�#![�/�2�^�dyz�oY�2�f���Vz3Λ0hQLC�o��cj�ޡ�.l�[R���� �yy��ҋ���<��ǳ7�M��q�/+w<��o����G�Mf�-�u�cDk�=�z�8��!ʗ��n^S�Ő-��״4��ݹU�`e�+�����ov侉���9�&N��	N(*�����H5T(��w9\��Rي��Y��U_�
�
��P���> D����:�d׆���V�����`�����͌��0�B�a�?P�X9�8��}o��Ũj6����+=�{_T��������.;c+���q��fpT�%�lX���\'Y>�uh�y�0���c�c�����/6�B�8��+��R�Ǿ�\�������}�#��N�Z.�-�J��s�N0���@������}[�ߣ�O�j[:�~>��!W��.=㭒w�y�(�l�·�4'�lb�l�E���@��P���Aɱ|�L[�X�eY��^�ks��`2��p�,��9m��W�Կ4X}E��׆o �1&lH�A�`�z㗷�CK�O����u:!���R����~���������5;P�5�P-�L�KɅ=>�˷�gܡ_��.�Wǭʗ���?C�廙�� 9Xej�`աU���S���x���rf���,&wP׉����"�}�EWޑ�����
�,��z���V� ���>�?W�a����X�x�l��ZS�Y��bZ,+�*��+�:�]	󕝗���7�}�1����w��j�ɰ���
�S�XVf6�	� ]�ށVm��m�w��H�� �넱s-;��{N�CX9�B�a�y�h�o���ǷC:���@�NRi=4�M=��)ޫ�+<��ݦ�tWB�5ymV,����V�b� ^q�^���"��Bd@��X�x��˨���	�t	^n�7���Q��s�tD�V.d�"pp�&{d�ݾų9��q���*"��.����)�1�%qL�A���}+�X?���T����s��{G45�T�J�����ND
�jXM�����bU1��[�٨^�E3�;���~�+<I����C:`�~�y~�>��;z�N�lMF �L9ϛ��0��;#|�{�i���Ş�<�&6�jQ���*�D�"���٪_nٍU�Q���~����ّ��qaM�;~�4gƘ�e�2'8ߠX۬�}b�%�@���Qc�B�����}�kzi?���L�oG��A��9~�u����v����t�6j,d�L0�c\�B}�t��uJ�z�/I'gt����(f��D*�/G�ۀ�?{`��Ҕ*�["��c�?/j���B�yy���G�Z�6����P"��ϯ��r����bnf�'�L��t���\��������вQb���r���tX��/c����9p�j[k!c��/��Tȡ{���u��#���s2��m�Y�͢,�b��:	�D�b�j�����������b�ob��uYsZs�_��ɡ��Y�`}s6qn[X����;E�m�g�jSQ��iV,sB-S�ѻz������SzRq m�H�[i��ͳFfug��������_뺿�*���+����Q$�>>������5q�j=s&p
"�,8K�ť�u"�ڞ�ծ\�p\v��蘿,M6�a���g\��"�M�'�|~�D���^��f:Gݼ��"&|�8������x����{R�:�/7�x	��g���4P�Ę`���/�����s�1<�ezkWϗݬ��,;y�0�lηIN���j3��\A�[U�bH Кqo�=
z�o�pX�>ҩR9��T��M�T�.����Z�ㅢ�J���]�G*!r�,K��D]��*�X6z�I�I�g��,1Y鿪mϜ�ݕ	
ZM��`.�Rv}hJBB�*��\+!Fډs�O.�M�����x�0�ʹ�O@���"��n�N���K~	`�}������b�J�5���{"|�Gd׻��������YS����X�zT]NCr��ޝ^�pc>'�DQC^�ٗG^������;���~�AT�D�׮p˲��,t�0��~_�X���?>)��~�E
���'��A?)�&O�<����9�����E���62f�$lW�+�^�)�\�י��Ȝ��(2����_V�Pwg��>3$�yx������$w�t*׫�ů��U;��sf�Lݺ2�H⬩8�>�Q�wc���;�2�Aɍ�n�GUv�V�m�ζI�͖�ޅ�^u0�/����Utek�ܥ��8U�M*����@!Q�AX�|m�o���1{�LL����@oo�>��8�J؇��9�?�<+�Y�z��+�,�8����y�*SU}���\�-��\r.�"s�W��j�r0Hd���7ym�q�=��t�Wq�Y\�Z^��^D�ɗaӎ��1�](>>�X>�g��-ς��/���ϕ�>>����^Y��Q�f|�/Y��VԼ���z2�����\�k��G�x���ْ�q>��+=W�]�wXsc�Pk�r}_O_�l
1_W҅8�"	�lZ�fW�2���g�f��]%�.���<��	N\�87�*�7B(Ё^��rc@�@Ȱ�]�]/ɢOnv��ř}�y�?y�cS{���|�9�L��VL�����vK�2V]L�˚�_���]�t�S-���j���n�6ܨ�+[9�=��]D{~�٘�mtt��^�4S�O�ݖz�}����!-́S)ɹ�<|�caո*�}:7�u)��%���R^}���q��|'�*c��%	Q4�8Q1��>�s�,W[r�� 9�O�q��{^�/o?]Y����	%���
ݿ�5�l��v��T�
�����)rm-��W�b�*���̉��uF#6'6�n$��i��J�Ey�6�L��z��6Y�֘�ىx��Ӧ�)n
�z�HaMS�w>Y����_��h^�N�@E$G���3�7޵��C����0FJ�N��Fj&�DY����E�WOҴvX�oA8 �{�ѺEM��'�6qioӽ�^�a;�1�'��5�m+���쯧��%{�A{j��n\�����/3�˙9����1N�����{VDV6��u��p-\�ǣ���s��d��
�8���I�x�_.���-�jI���c3o�'��;ʛb(h}X!�?�N�݇�V� �lש5��@��@�*�a�C��Jo���`+��ھ��ϸ�z7��Ü~�p��tHY�G�ف�nũ]5y�m/r[��9ř�n����23�U�q�X�0��`�S3���~��=^�"�c|7M��J�4���)�C>�@�]��㕵+g�>)G�UDn��n�~G*\c9�r��&k�Ds�V�5�woK0v\������^�o��]~�V�<7�����Rؑc���H�Z	\x���e��^�o�_�����E�ŎT'�͌S���-�~S욁���Pa��y�ocL����{ǣ+n�
W�T��3���&�d�)�4=���꾛?U�<>�ٵ-���U43���>���'K��F_5�؝߯�>3��ڙ�R[[5��mu^��vq0o2�,�0 �1���b�n�������^ j8�\������Ε-��+�.~�EѮ5}Vm��[RBu���ق�!Ytr�e�`�.+8pnF��:�HPC����Qb�)^n�u$�tՔIt+�r�!�U�N�p}p��gGqg���:�aD�� �ܜRړ�F�P�pAfFE�61ݴ�5&S�B�T�Ή�������JU�[����Ȱ����G�ر�%5��O-�����pM�����n��k�����_k=���(=�Ģ��\dYڜ��6�J��]ҡEV��P�3�wS0�Q�9��^oa.C���kR�q��f��њ�S@��n�T�ó�D_��ErԲ$TWga�fB,j���e�N1͍��)T2T,z+'mB,�aw+��c�$p��K�W][��b�Д@�4����y�b˫�[�M�@��8=��i�B��wu��	\�.�j�S ��=+������3K�"��Y���j���E���x�]u�67�#��ѽ��S8�s\O3��� 5�9��O6
l�d����:�Ϊ����*k��u������V�����	L�B��i�U�7�v^>�<���Ol���7 ܰ��A�Ϻ�͉�%yoP�n���fl53e���DX`U��ECQ.�W�Nv�����kYޥ6gs՘�|tngjz���K��f:�;v��5镧w�l^,���nl
�\��X#���R<�N�C�V��R.�h�
��c\w�2�ݢ����Ck3�vͣ�s�4e��5񑨇+�(u��q�TY�)	��z�$	�Xe���1a%l�Y�k�S�z`�k�]}Z�a�47�B�j���g>->pބ�nV�Z���}�ש�8����JHYգ{^��.��&ot{M!H9}�y��-@�sEԎ�jݰ[�6:M�'+ac��6�\&���,l���q��S5U�gl)f��NUf�0�b�::6P���;trY<T��J��$���N�ƀ�t����ڷpHf�2�"͖;�.�_K���ӠF�lo�L���7Eq��Y�6�哭������{]|`�n��<�}{���y����o��!ѥn����epyϭ[|�YE�31u�v�[��������t�ỨR�/V��,����b���m�j�4��gl�v�9r*C�?39jBw��p�ò&z�LX1j��G�@v�R��pO���U-�*�|��4fp��6S��K��^�qZ�djɛ�]}��¨���m�-2���ոpX���n 	�[/�<ə�9�T6!�р�똺Y��H�+l�tĶ�)���o61E��C��]�9+�)�b��Bwrp�%F7�;u�V7/y]<usX[E���+t�x}�2��`L,�xi�Bu]�/FٗSFh�:��{Z&[�w��oo������o}�>%��Z���w�o�(�>o��6���9��В�ڄ<�gi(�ٲ��~�_����m^v�n�s:��;��H�֋�}�}˵�Rs7N�z�~�_������\	''p�g$�ԏk/�����'��""/� &Z�X+�%�����W�������l��m���t��<�ebH���_z�<�mg=n�q�k:'O;X	}��ͻ��Gw�C+FY5��A�|�u8#���B��q���#j�Q�!Ēs��o�{��q)<Ҳ�9�2���NIē���x�3�-A=�q�i!�I�qbJ>[��������4��2ΰ��7�ZOm}m�dj�G^Z��8��rDEC�C�݂��E����B!�Y���ւ�8���lAŦbIC�����,����2�����9�j-��x&&�����5�"\\��=o�ZW[6�]ZFT���8�'���Kq�/yк�t��.�ն&m: �$a �VAAK���Lo��C�� bF���#�T�r��\��V��`^�nsS���r�3Ĺt���3���/1�oʪgٷJ�%�����AAS�+�{cV�F��<S.��N�;�/^�p��2�7)�yHc�tO� ��]"1	�1b�� 9`�V1�V�A��{5U�����cS�1�7�}�Ve��9��n���5��`S�eZ�H��%��(O������7����b{R룱�y�����~6��7q��\(��9�:"U�bЪ��К�N�6"�$����]�98ǲ���n"��b����S	TB��Z3.3�½>���鹜�%Kh�����]P}ދ�o��X0����œa	�&�Bp�1Z��^����������=F�����u�OhDO�a
�#+޶��sӑޗ�]�ؚ�^��l�z�L�r*0�ԏ�N������g]mI�Y�.�nG_����Q�J�.60qvO�`�7�1�4��j���B<�^�&M+]"O�u�+VD����p�qc�������"3�����ޞ�(O�F+m�&G�m�҅;HU�8R����Wn��N�nup��qM�JI��Qۥz��2��I�^��RC.���=b{]�x�s*);f�]^�C���R��9��Э��r��3�&��&l[jf1]��5���.��d?� 䊁� *����;q��ی��5����kv7�b٨�{�Fҭ�Z*�6��ߣ�Nz�:(��-~���O�׷�QkϘ��?;1���h�V�N��6��V����4�6}3����ۨn���V��Ff1	�"�0g��A��{��r�����f��zciXu��U�횇�����!8�nmץ�Ę��q�N�ώR�tX����o�5�\����3Y	C{�9�QAF�:�/#}G��5����2#���'"�ATG��N�,]�����Ff����d�n�u���+I����h���	`>��u&�r&�P����t`�+��e▮�D�	�=a\���U�>|z���1�"�T��>��s@ǀ�~��{�;"k��$S`+�k�/���9���R�4�fv��9�6�y�0��:�%;��R��qN@��GD� ПtYno�R�җG�7/��q��>��U�p��tr{BW��p���D%8"ar�afs�G��]Hk1�&�"������N�T)9�u������;
��%!!o|Ug��J�q��]n��튌}su־��~�h��|ە3�M^Н�R�� ��>=���V^�x�������|dm��
�닲]��C�G�V�&v�֥U�M�kp���b�ʜa
Y!N�����KT�vF��CyY[ԋ#P�zp����?�����P����G��������8����*`�5s5��W	�V�T�e{��%��g�:���>�tc�ȋ�B�^J�sp�>``2������ꬩy긚�
QpǥG�˭��@9[ӫ�#�wt��RJ�����B5s�{\E%^�[~��jdM޻�geWK�߫��x���3����~��k{��}��_˥����2�Dv���<]����������3Tɺ�5a���_�lq��6��[�ݳ�l�������:[��g�8�n>�T�8C[�s���|�{ӛ9�Jn�sc��)Y�s���T��k� lxU�~�a�8���y���0�g�U�s�7y��/t��;�/}�]=�^�{;g#fv�R���1�]8�(!�Z3��[���U[����p�Wy�w�����klmw��>��Y�4D
�¨�E�ۈ��D5�0/[���wV�2#���w��1��<g���.�K~�͌Y>� ƀ�yNO���[�'�)�ge�}�����j���g<VE�i���.O%Z��.l�@�ؓb+��tcG�x�o��/�q蓷3航�P����i%��R�t��Tt=���!#aJ�P�;�����u���ݧ�!ڎ�j�EfN�����\L[i�@�9L�E�4��[�U�t��,��D�/Lj��Kd6�àࡕ,�U��>$!��2�v�'��{���W�T����w�%�[�ƅ��6��)�sג��v� �{��lʑޭt�F�K�ʘ3�0*\3!UTuG�S}���;��l'q��SY�`�/VX�Y򵞍�6ܨ����k���̸�.$Ի�Vs�����_L�c�*O	0(1-͊�數�T��{�p\*!�y#v����y�ٳU� ab�B�O�1�Ȫ�U14bz&�B����kң��8'��ؔ�B���RJ�x�u�x���?�g��(�䍗�f�hp�Th���Z;,t6��>[�f��'+��\4��B���������1��C��T�µN7�K:���bEE}�h�xl�b8͝���s'Ff��p�mrW�����+b�Ꝅ���`����Ѯp��X:�L�-�<���wg�^�`kV��,V��S�Ϳ�鬏Tؑ�����~�# ma��+����{�a�Nt2�hW�93@�C���%=S�9���h_Vl`�L9���Ü~�p�7:�"<-�k}u=>�:Z^�Lg�k�;f���t������җѕ�c >��^�g�b�-Ĥ?g�/�U�s�f� ���շ��-*���u�y07�9Ro7r�����j�&*���̓�)��%1�e,�A�݆؜ٵ$;�	r��دCa�v#;2s77��9�2�]Թ��IM�P��u��r���9��������*�׋�Zg}��k��ƭ9���z-⁑��~���mK϶�@X�9U��]71��s��joo��Е׬�����aL��SJS�7�^�o��]~�V�<�ߣ갅z,T�$n���/:\�^�Y�z �w0�X>wQqǎ��p��61N���Q�)�3횁��<�t�q�s�5~<uR����N�=�����Ti�n�G%{K�,�lv.�3z�g�#k3�׏3�/���%K�D�QM�R�8r�J�{%��Y�U�5�ۜН�R�ֺ���@��VWd����k��P�jf"�����'��@�F
�����2����M/H����5z��k����g�-F�;��;�z0�_t�?!=�OA�4���vX5�C�zdN�g���Px���Nѝn����IH�֋0���T H"�����1u�+�Pn}�h9T��~��Q���."������C7�b��w���f����tD�B�HR&��z6;[�g�����r�����RM�A�]���fJ�LbW�J���m+Or�?��Z�uoʊE���m��*F,	co.E�_�o5�	f���2��c�ӳ��u��Dƌ�O����6���&	��p�e��{V�T���5�ܿ�E�{���D�4f�b��i]8�dwR�oz�3���_5m�شL���:K��wjY�k��鑚_i��kL�tA� � ()����$'�{^L�_�d�)�lT۟@���4A9({ըMA!-�B9����\zMQ<���j��<��૒�&Dwa��"���n|3+zvK���M����aΪ�Bf�+L��;~7d�0G޴42�}6�eF|n��gƲ&����nE�'GW��c���Nɞ��&:��7Ц�v=�n��!�XQ�?{&�t��V+�mD~����/���k��L ߶|�O�mZ���[���u
�-Ƿ�U� ~x1΋g�n�}Ӟ�٨�����,�e*$_\n��坄���aP�#�>�ߐ���R�AM9L��q�Soϫv}�ޚs'�*�^
yz��wwb���7R��
�ßE,,�����M\7/�k!ckYɌ�9�m���E�_<��p�u�)NG�d��J3�)��qb�/c����9p5�����@ΗU����,�2s���`���&DtԉȠè�E����,8X��1h]��`�z�:�TN��<��x<����S�8eC҄�:���+�O8��::3�"�v^)h���]���W̷'Ӗv�^E!7�V����Wv*.��^���`!��}���HU��_t��K�fNm�&i�`�tډ��o#�	���03N�m�W]s7��U�<5��� N�q��)�1M��,�N@�[7F�e&N�{9��I��7������"�$EDR'�o�s4@/�.?&��-���`%U��3����Q�'A�+�(�_�'b�O�5=�Һ,5s���՘�a�v�aFٝ�S�:�B���#�r�b^��*3����f���{���:3�r��]Do�{��V���tv�u�b�]���2g�
��[}đ�-/b,|"cnDB�,1IL�t�O�eC��wX���ԝ�_Z�!A{����ޘ��"3٨��h���Q{.v��6���Ĩ#�DӬSò���V!.�3�����\��:U�&(<�aig��X�E����S�g�ꬩ8=W@1J./�=J/.��s�8��j�W��o#=�h�'<hϹ(�~l�E`~�!�o01��S"o���&+&�GM�֊1p×ǒ��@���C���b��w>�[�{ͼ����y���klO{��}�Lй�^S���O_R���ڏdՏ2�lz�g��'�_V}Ŋq��!�n���W��zW�;����;̟{���'�X�Ks�4t=~p�.�bp�������*��	���W��\�vMa��{�@�l�֪i4=�sh���&�o�2M��d����N}ʉ�=�'��T��xe��/	}���V=j;����&l�VP�n���@���T�q��:\jƔ�&��Нt�2��x�:������c7��-�MZ��y@NH*����4��c�f�3�sߗ~4gz�ӭ�T28���1�t�<�`��Fx�r�����7�4|�:Fղ��|���ky\\kxz}��Y����x}4Dl]7q�vY�Wd�f�	�0MP�
�6��U�5RZ�)r���f�,�@1�ה��W��N�����(S��O$��N�R-q>��s�����~<��ƪpjR�rZsa)�\�8��HВ'`/�G�r�̎��'��T�r/�up�������3U34�~���p'D�>��8d�Ra3���]Vw�c���0�m�>�0�0a���2+Y�����*5򵳚����x��ķu�˯���ܙ'�X���d~;S/�MGE9���Ii��ʃ<yX�][�rty˽v���걦lO��M�����v�`2tO�pT��jH�&&�B�(�:3�6!��ߢ��~�9͒ �����w��{r�������S�p}$l���&�q@�m./e~_T����b���D�iU��.?��mw�8�����!�5J�X\+T�٥��\�1"��abl^����k,^���y������6��^ *s�<�i���]YCH�7�\��	x�J�ߵ�`�I�=)��H�H��k_q���M�e�뛖\�j�9op��Q�Ԛ�l��\��s�Ė�L��M�Ν5�r�.���Vo�Ԧ��l3�@y"�B(8���?/`��ώn�~��,W�y��;foJa:�b8�s6z5Ɋɤ�T�4i��L.�]��{���t,�p6�o`������՞�)lH+��8ϛ��ڿD�-����Cs�\�-�&������XШz����]wN�~��辬��8�z7��Ô7-;���W���2�9t_�H]�g���lѝ�틯o��f����V��leb�Ϗ���}^�gO{�,Q}���ڴ����dA2�Vz<��x�dgϽ~� �mKͯD�)G�UDn��nc�����^���zwK�!��Ã2��2�ܽ�7�^�x܍ߪ�g�g�+b��G��Dv��RZb�LĊ�Y�=��n'�8�K�g����<p��p��61KeXSզb7&�����)鉙���c}݂�l`�����S�u��y�E�9m��	^�R�>S@žSc�*��)���\���vi�f��v'�ĉ��ڔ ��r��ߖ{-���U�5Bs�����ɇ1�eT�M#I��y����b(���r'��T����+�Y���V�F�މ]����"Y����Y�ڑ����tY�WV<J��)�8���goV�l�[�ldSݙ{km�!]%���
�Z"�92'+���guB�����0�Y�s��[��[�,��л�ק;%.M���cs��J6���_sү��Nq��z�ޯ�W��� �� �g>�/�����f�<��:���c$N��b�eFQ���R)q����T�D��6Ƌ�^Xuo��m���)��t����c��
=K�~�<�f��c(������B�98�.!���+���C7�/��Fv7�
03C�T`�^X�����r��.;3�k��b[�"e�]D#)|M�������!t�*���b{KGx�l�- ,G��}
k��YUn�tQ�����������Y6:*�a!8�"�����cV�D�M{�ۨ`𭇃��~�8:�D���[�G�	�z��BZ�%~�U�o4}~��K6u{;,CWY���A���G�v�8-	q��mK3q:<)@��[�c��f�|7m��Fֺ�����#+y�v�W�T�>vN���������]"O�۬�]7�1N=�t�CS#8�%>�5�ǶQ����0�;P�u��L[�o�Xp����T�n���W�,þ�,��F>��.w���Y��
"|��"0g�E��f8��u}-:p/���gջ/��X����̮�/,�v�n�N�&ب6���y������Y�vlQTB�>6�o��vQ�C���v@�70����&�n��:䀝P;	]��,ۨ�)b�̋�hdT4�Wj®�i68�Ay�/g*�y�%\��˲��7����J��-K��ѽ��p����[QT�H��c�� ��fZq�7\$-� 7CT�Mۻ�A�ru��w�S�'ȑ����W�����J��bCln�#3�pNҩ�Ǘ2	�n�f[23ۗ<�0&֎�6��v�*�cf��f&��Z��u�P����lv,�c��x*����R�1vtg��ql"�j@�z�t��[U�1+i@(m\���R/	V���ۛ�殽�]3B���ޒ;;_�n	����GQ�ٱ�9�a��AAZ���pۮ|)^7:(zռOu�.�EnL��#�VL�V����-��G&`B�ó*��v�b�w��q�ԩ���w�Y;coY]�9j��`�n�FRк.��n�bm�uu�h=���u�13{����e�/w�%;@n�V��4.h�0�i��H�;\�.�ǚ�{�Х�9����U��[�H#��vQ�ʬ1�{�N��Q9G&v�q�p�y�T���U�nt�O�D��([��,J����]ww�)���� $�7�r���Y�bk;��r�n����fޘ��tlš����1��[�
]_`%��u5z�j�D�J��mf����h���2L�/�ǜn�t�r��i+@g���t��ߞ����r�F����(���JK��`�=���9؎��a�cdޙ`Ω�\ե0*�U�D��X2�qsVA�eeR�Nk5eY��S�+��ʴ�n��bOO]�y��n��
`t����̾,{L���`[Lׇ4\4Wp>�Y[g�v.o .v�7k�;CF��8��ܧ9�@ՑD��O
���ej��=����)`<�Z�cW%�vd=�4-�,�ࠡN�
��;:���6�Z�
-X�r-�6S����i�v i��W5�hoP�QBv{yL�^7r�͠��RY@��ؙ-�BmhY�-v�t���-�5�Z��f�Y6Ҏq噕��+6��ok�����}����yA��|x�Î��{5�(�Ζ�]VzZ��t켷�*WL�������d�uXq�f�����V����F��#4���T��Α��T�c���3q��uʰ�d��C{��n�I2���e������]�EW��F�t-v��#�<'T��[3��>�Զk��mH�C�;9z�Ocy5R�v�[�X�`��a[D��1+k��2�ށ��b��_�X�8LE���'T�X���'��d�iB,[��+o@�j��q�n�(����>F���Nj�*q����QD��60�ݡ}�{��a��9G7h���tP�\��mIlSˁ�6㡹*g:�kkHp^��3:�{�����S��4�d�D�����{׽��;�����Ȥ�/cM�8�������i�a����+4�E�N��9��������"����7;���rA�i��$���������~�	#���r�_�����ӽ4����
;kE�3��8��2�3�(�;0�m~We�::;�k�;��u��G{o��8��2�����������j��Yy���|����Y�u��݁�6����g!�D]�e�p&�nGmbBu�s��]�Q!�F����r)�Z{Q��t�E��yg9�ݡ#�Nq�n���h������8�kt^k��+k�I(��P,�ܞ��� Btt]y�w��>�d�>מwY���2{�tu�y���:8���{ޛYo����ޗ�5mn� ����6��,���k)l��z�N�����Ӳ�W��ڳ���q��w��ýnݝ�QE��b?X6wя�E��d\�E�{5P�ax�V�{�r��g5���}�sH��&ʳ�\ܶ�l������0T��ӕ��mR�������닖��F6�}����UdTq�����D��>�Z�ϯ��r��n_�3Y����3�����:�u�`?���wn���=`�G��@fZ�bŋ���t͹p1\2*�"�udޝ�+=W�i{gTM�o�T�Q�Q�L��9��yZ�hYcа.�Y��]��=��{��}8If�[�58�Z�ƧJmԘ�"�M�'�@��@�D����2�P���g���ۅ,������f�ԷԔ��1�&q����;"OH���0;'�4�3bso2���hy�'6��Ec����#�1F����@*A��[��r^*P_�q �~�(c��ۭ��j)�R�j��X�1�&���0�E�^��Oq����p�C�F�W_V�vc�����t��r{5�'��&��,:\)���o��w���ϻ�Du�_�IߡWք�Q��S��]ʾ��9zz���U�X<+!F���\�%@�R&�b��t���	�od9��L;�}�q����=RT��6(1�U������YRs�q,J����R�˭��|�/�A��

��~��I����(r�q�A��m�d]E5N�iMɣ�X�*��!I���ݟh��{�LM��]�m ��HW��S�n�v�Z2.%N�T��b(��FI��f�i$Rf���*n�W�Z�፶��u�m�5y1��T�( (-1l���y�J���0�yX�n�߰1��S"w�����_�7_h���8���g��Ro�(I�a�'�;��Q�>���M�Gj�bٮ�� ��	���g6���W���<���ե/E�6$z+��7������t��ϸ�M�����0kw�tj���ښ����Q�k��ke��٥86}2���O�\싰؜�a�<0fXr8Wɟh�(���eW���֨�f<�Q���8#�`�g�������W�ʠ��_����}hϤj�_gj����1}�΢��{K�'�˫R��v2n�d]�1��ږg�#b黈��ȇ�t��7gj��>Ͻm��{�{�0*U!�x�����)��h�� �F�N�`�Բzhb��\w��m�?S�>,���d���D<�ъW:�#U858�r[����j�WlI�/��y���H�{�����*XrMCS�sאO;��<���~���p'D�9���������f� ]Ij���^!�#��b�����
���O�7SJ�s��e���Z�F�nT.��iA��Q�ٽ���h��>7ti)k��՗D�$�F�fXOOj�9�}�~}~w7��k�V�5�*��<�R�q��Ԟ��z�K������9�8-kv�/.�����&�-����͆�
"+���kb\�N-@�8Mj
���Y�%}I��=��W���T�������Xg�x���ݗ����^��1�%M��KS�*� y`סո<c-�wmD�1&���!���}e�����Z�0����pT��P"xI����
D�tyO�*��D2b���»�d�Ft�)��a��[`N�F|䍗�"��M}LW��xx?O6.�1׺4�q�r��kF\t���>�j-�����!���*�#�S��U���2��}:&�til��]t,��ŏK�Q�����r���M�^�������1�;�1����C]o�JgnFz���޿n��U���ɚ@л]�c#�OQ���^��>�z*68��>o��mkzdt�ٻ��Ng�i$�&s�4��b�f�y��\����V,��`?fv���ca�B��[s���/64����d�������{�2^��kz٬"�~����*��O��m���J�zM��k�&|)���7��^�e�5��Sޖ�ܷ�b��@�ϟz�VԽ�E�/��_dȬ��"}Yu���Y�xƚ�U0���t3T��Un^��k�m���u��V�<�)�Ze�~|tw�f)�+g&{5W.��-Ѫ=8����fڒ,l��֞��Ʀ&C��6�x1��2�v	�w�E6Ay;ot��ޖ�?R  �ߢ]�?v��B�u�fY�'MZ$�7�ٳٶGI�9\X���{n>�❃��}b5wt�Ȭ�ƫ�Slҕ���h�Q� ����w֬���	��bA�b���1��	�:���M	��lb���o�J�"Pf������z�d�Y5Hd1^�,9&� ���\<^yQ�鹾J����9h�a�Z�Q�<G��V�נ{�k�ʧf��>��1!��� ��r��W�-p]�j�f��	��=H��]۶L���֡�k���`s���P�T�nD�:�K�uA�S�+�g�j�;bVz��z�ե�˼��#E⁏��<׹�n	��3�&�DB:@��]NYF6s�
��5����p��k�4� ��3��S��[�!PưY�S�eX�P�D��Y�T���Wݓ�яfw"Ԗr�a�Pg˛��C7�/�7q��B��5�
tD��/e���c�y�Ƴ���{Xɖ�	"\�����e�'/I���֠w�*�0�D/O|U�\Έ��yԃ�P����Bkc�{��M*�YU�Ȭ+�n�����C^����V�5��HNeG��C"��̿;�;�Ɩ0Ci�E�|+`����� �V3>W���'W���T%���>K�jeK?+�b�`*c�(S����*~܆���%}�LQC�U}�0����h�X_����Fͣ���ᵗ�[�b��^c��L�eN�Bl�<N-k�U�J�W\++z֢*��:��M�;v�1r��Ҵ�f�	Iq���ޗ	^p9հ���Da��H@QN/s�[�7ⷙ��Q�� �{A���,mvˌ�j^YC
%����T��c+�@��Y�l�3t��B/�yq�����t.�!���b��ƶT�/MD��S����KQ�����%��A{mо�����}�3�L[�o��y�Ѯ}mvf�hNm\��=��Yb<�$Gz�MI��C��J/�_	�g��Δ�p�D*�/S��
m��������^�~'��x��3W9B��8U�>�}D��
pl�(v��Ǻ�)^
j�BJ}2�G����oz��k���1���:p��ۥ9�	�`Uv>�p�9_!E�y��:���ҥ���;�߷���vd�|��-��8�T<TrT`��BD�Pa�G�H��,8[��ױ�4�ؽ����q&s�ز�OH�n�J��='JmԘp*D�]Bz�WƠK��o7�Mu��O�j�.�!�{n��T��F|.��;U/g�V<x	��4�;"k��$U��I2�S�=O�]�VJ'ӽ� & e}_H���v^G#v�!��YF�N�IN���U�~ڈ.��9~s�i���v�$VjN����$�M���Eh�qN�Q�y!�U
���T�*C�Y���B����:���<�Z�c�f��d��RbK��֮U�Ԓ��5���]K��MN��t��N���V�1Y�n��]
��`2����XJ�FA*��B�b��-�NANH�B""Z��vָ��I/�'?}� D�4%�nw�c�ŏ]Dw�x��T��Q�������/t����\��G��DKK���DL5"# !P���M��N�T99�b#�[Rwmʏ9��������n��[���,s���xMtT¿�\��`�>R&�j�}�^�l9��/`OS�����Ǌ�׎T�j���-��"mO��uVT����ӓ��7�6�t�;�����	�qp���f,͆��ί3�`'�DR��p�>��'ndN��Ͼ3{5:n'hd:���g���e"G���G���z���Ð/�+�rv� ��Dv��!뭀�[>�(q��w{6d�Z	>����y���ey*�ñ�46(h���~����t�����Ÿ��lC��[�s���Lv,�y�۴j��1�ُD7d֊�V�I�?tu�H���a�8}�ϫ�`54ÑC�zP}�+}�����x���6�!�Vɳ�%�pN6�����|�������Ӏ��,!Ȫ�R�&{�W�fg%��U��0朵��`d,�q�=�c����ᯤPU�Sw�Ћo�}7�S����p�MF��,����#���9*�prխ2/�Xo�Vu˥�fT��	��*�R^������:��)K������MH���]%)�07��p�:���٭rؖ��+,��Pѥ���e�]NTm7� b��t 1,~}Gߑ0�@���]��8vs���:�`/���E�ǍϾ�X�?���P`ה��?-��b/_�)�wߏnu����Ĩ��dAϏ_��\�ƪpjR�rZl%89;7�*��������E^���Yǭ�L@��~sѢ��#�j���<��4�C�ܐ�$H�͞z3r�=����ɝ�Ss0ǩ������@�f�L9+`�/B���n��ە
���L���Y�}��w1�{(��%��ko���\G��fb;�`BL
BI
�\���>YP��s����ڦ\�b��e-�T|�I�{8T�����;mVϔ���pT��jp�hS�S��3�ΊY�� eo��ݯo����⤿�����܅�����a�sj0px,�K�O�ȥ(\�	10�6e�_A�c��'0s�`U�9ZX�/A8 ͮ�����1�7q���x¼��Y4���=n3-��;<xs�=�2e��PB�F��R��Gl�o���Ց�m)�	ߡ�-T�Q�{/J��f��ď5�߲Y�@�gadBr�ҟ�`�M[���%�N��S�~_�����8��}� ��"#c#衁�g�7ڳ�E}����mv)Rr��5��(9}��VΨ��hn*�{˓To[݃�%Ckj��V,�\�VD��A�҂�6�`��*ol![�)��M4>�ˆ���CS����xj-Ka���҃���Np��4���!�H@Av���/�Z�qmS^��?��9�A�s�X�����u�s}u�;�fvH��:�bYJU{^����a�Hݭ�GI��4C��.|��{��pL���z�P�~Uo�I����{0]��~��fY�+|����O����5HC��U�^�x1跊F޿F�.�(�\WO�,�y��U�G{����L[�.����B���1���s�U[����[��l�lc"�^ٖ�n>����fY�X�wc1����T�$Xt�<>�� �UG�x��)��3-O���}ޕ��^�v�Q`��W���\�(�
1^��A�ÖS�.�p�/<���-��	^�R�+��B���I�8x�p�����׆o*�I���Ćf�P�g>��������[�����r���;���F�����9�9�څ�vTsS1�>���.�`���2���8��{B����oV��5���pV���΁K��=gdM�$!=�	�12oơƽ��]+�`�2y���X��׮��B6��n���r��֋1����P���c���m �P�sd�?H�"`�}��HF���6e?��7\�6$��&T����a���m����N�_�M3����n����@N����xs�>�7k'�&3��
6YL�N����48q+Fq���1����B���1�[���bU�W�3iK�D9 � (��3���|mŦpmq��m�B[����`=�����5~�Cw��7�
1�s�+2�Ӻ<��b:��Y:�����:���D�l���q��1q�]�P
�S	TA����y����Yk��Ļ,��Ϛ��%V�@�zY+߫�Oh��*��
���qofbɱ�W^���6�'���	ǀh^��1~��I���r5{591~�T��R��:�2~�s�+�ac��=�2���<�Ϲ��R�MC~��~�� ZϢ��e�|n������W�%���1zU��4�v�Lnۍ{}����>���y�~�Z�#"p7�6�*V��ؗS�8�3�Ғ2gO���Ȯb�t�ԁ]1�r����.gƘ�*������t[=�w�o�}'ao�߶M�.�,�G��}�PÝ��:ط"؟`t��"���-��UnZt�8����[:�6��GkÇ�ƽ;�e���}Ӏ�zi��Lб!zlT�'�"� �>>�Y�Ϭq�nY�{�w�"�S���^7�������X��F��t�g����	谦#�.2NR��q��;]9yw�V��<TY�P��Z/f��{�Q``bA��G�)�-jz�?L�ZsT�ٝa�=q}�
���ԛU�QHߟo�ŉ|����I[��{v��ħن��Nᕐ�e'ݤ�G14�c���F6�^�-*c�1C6�!��O/���y#[C�l���u~�U~�}� ��d����3X�@ֲڗ�5���ʃ�*9*3�5"r+�è�E�DS�9�a�����}̛���~��Wb��٩+ծL'*f�I�Eȕ�'�|ek�fx5&(�	�,OG�Q��8j�ܮY~��.��;U)�����/dgJS�%�mUC����Xj��!�+`���%�����n�d6��@(��?7IN�������#zRg�Lq�k�׵�'���	�����^�u2�^	����xD���6W���[�����	b_��n�ʈJpD�J�D�	��ة��)�r}����ʮp�s�;g�9_���%1��B����V}±	�60UB3"����N��[�)��R�j������a�����?X���΅�ؖĆ7Pc�'�:�*Nz�&��	��@؀�Ǳ�U�q�?��,KT#�¡�y�B+�	/"+}N)��2&�׮p���)v97L��a��]{�~+=���%�N.,��f�_l��e�fs��ё97����x5ߠ8�ױ�� {�K'�ɺ��^R&bt�և\�WF%��,�T��{~�A�lK_u�k+QU��Oe���)c��%Hhi�k��{\�kͽ��a���o5U� IfP"�N���n�t2�m됎���le��"nt0�^��V�Rc(d��4�qS��{�P<i���Xo4io33hX��`��Z�o���ڞ���6���`�k�!1S<c��V���xtͣ���v�ӕ��s^�z�n.˔���	�:�Yr��HL��U*�y�4a�LJj
��Ό��pڱhi�g4�l��g4�dF(gEޮ����<]p�
ݮ��`+��F�_=���ܲD��9m��� -��di44'&a�W��+U��ŽV�I]Ckm���Ji�R�/7����s����{Ȑ��eK>�s��kJ鏯٧��ٝ�ONa��+�k�u��ӥl��(TѨ��U'H�;"c$��i��H��TU�,������f鳻�E&�^�-������t=k%d�v�3�1ٰs� «�v	gC��a�T��hx+/ɼ��[&�Kέ����D�`�a�rش��Y�7�K;c����9����&:B� ��AZ���Bn�ޚ��Rĭ�0�f"w�i؉��\�
ˋ�\�ͳCr��.X�Y@�c��Lhgz�brQ��Ajł�;hp��G���%^�[9x̺��M�9R7N��Z���N�id!gmf�݆![0�o��JYD��6��n���Jn��7*��08B�m��0.�Cj�]����J��^rU(���2�����	�<�����7���	J���?n���/K���S��KV1��(�׌��V�8V-ҷ.��d����q��2�L'YmO ��Au���ۙ���m�WORJ����"(�.|��7�8+Wv��DSt�f�Km���H2�WJ.k슐(k�+����i�AD*Q�YΪ��L��:�0L'L֋����6wE�6�O9�;:�`[D5�A�*n��T��<���Y5�B�Q���������An�������"Ƥ�[W��ŕ��oJ�:�鱯2�պ�S�A��6+1)��3���멳6�S�`�s��v�)�w՗�tw0�dvn켻6�M=�7Q�h0(��:��u�;���5|05|d��o&�Gn�o4
p�V��H�X�v���ثRep���L2��h����5��OzWZyF�rƔk:�,�x��}V� ���J��6�]�Y���3.2e�'^ERs0� ���n�8�ع������kt�̘�	j#qk��T�eѶ�
�|���N�]�B�k�)�b���� )R�	X��C�
���w�v�p��H����Y�l�J�+B��7	��+3

V��]u�c�i�ˑ��݁`������iΩ�N�gKic�ʝjh�nM�L��!����0����ŋ76.Q�s��Zu�z������)�q������3�0��1w�ef�PY��ځ�s&��6��8������3111!�mk�;�YGW��q�	Y_��<�㈑;���&iz�/���~��'?n�,����tVvG�f^ؙ��{u�'s��YٜY�i��[�.�����~�u�g~z�����yd[n����3s�8�8	̴,�)�#̞d=�//:{Zu�,���������/�|����+�Π9�����=�fwm[:;m����^jHW��}k�;δ�!_kGOk�4㲴���=,;m��孯;:专���I��,B�&ж���zm5��;=�������i+J��K;<�{jWv��&ٙI=�^sn���';�[W��e�-�f�Dwg[��<��m����cll��,���q��3K)�^���l�����6��ƷXPpv�5�ZC��:"Aa�������m��v�k-��lt��� �b���Kɋ�F��s�ѧ����&��7�H��I7T�@��B�t�)�Dm�m&�P��ŁM�t�L�#�,W4���:)�!l�8���5��Z�i���?�zU���k�9��ǏӪ��M�ށ}Y��,[�%LC����̙네Օ��n[<�{=�3�ɡ9�~���Y�y���~���+^�:x�t�ƻ|��5�YC�q�t&�!趱��Wz}2%��L�R��4�#T]8�?E�"��P�[�]r&wL0CNۜ5V���4�^���8���Y���O�������)@�FV]��ח���,��""�����
׭Ԏ6�"Uc��W�b}y�|�yN}>����������}������v�+��K��ݖ�=~�r��A�q�p%Z���.lwB��'�b^�go���&��O�����@���
����Ԡd_����sאw��o�55 '�恽��5Y�{��2I����&gc�Y3z&�:L9+�e�Yb�UZž�W�*�W^�[/;��b����ɆZ������r02W�Y k�B�������4���vT�.�_E�sb3m�+Y���8��[�C����7�v�U�1I�?0L��bi
p��)̫���7efu�u���₴=1$�j��r�9�7�8�����8i�*�ܕ��%^~�|��PQ���x��sZ
r��#ʹm��+�>h�W]��]r(�]n��z��V��rIp陖���qKgJ���j��V��
��E<�`�I��m��� �| � |>�����Lתً���P���J�nBP�,��6,2�ڎrC��&F�g�K�O�^����G�P��~���]�]?K��h'���^��\�u�T�B�8���|*�;�V|A�2t�����"��C��n����2�q�<��	�7��uOz��'}�~ɕ��Wd��yN�o:��:R=[Z]�ҵ�%e~T�~�����c�Ÿ���`�����P,�>��}����n��/[	؏C�Ȍ+�N{���Pؗ6���b��?,��Lx�����	�,�f���*Շ�뮜��}L���Ü�.�tN ��}=u�+�z�CF��W��Zr���wrC>��I�[�nz}W���S�:
�r�;ռP21��������=�v����<�e�_Q�Q`\�.��޹�,[�S��~�V��ɼ��7#v�����593r��~�$�ȭU���E�RБc����\�`+���8r���٬��f:f(,���N��3�v��^���~3욁�=TBW�a'�, �t�������e�6v[�%�Dx?��w�y͌�nF����9v��U�\�
�6���ڪ�Y�7ZW����o�h(n\��(v�XK|��1ĸ���)\�2��p�6��ؔr���\�E�KgR� sJ���d�o�=�.�ӵ�N&���bff O��� ��}6�uc������sAE��M�]Vf�U�6$O����B	�snW���F��{B!nt�gs�vp���m��~�np��B��e@����E�M���.�T<-����c�B�����ۅ��׶1���)⁁�ه����1ϼ'�쉠�!	�Rqݛ�8w�f�&_�1���\?�e8xr�uX5�uo��B6̷)NE9&B8+���2��:���Gu�����Q�@1_D�F}BZ��Q�ؠ���Z!�Η���g`o.z�
ۋtw��{���8�C�^Έ�}b�i�Bk�8��vУ�ۈn^�aw�@�UZ��ӫs���Rץ�
�y�\����Cb\��+*o�
��)��6��:��	ȁF�Iܝ2�iz!�b��Ʋho>�4ӱ�N�1Һ�¶����u���P�V���cs��3���2
8^�gs7y�ʂ�z_�Ԙ��^��~���轮�q��mK�k"k	7�~WG>�~y�q�/h�k$1׾�2��1�o�ȟA�A�H]LC�����������T��b�b�zl��4@��.�eT,igj�Ú3�u���wF��r���޷�n��K�i<�r�&�T�jҹ��x4���w�����2��+Z�90��)�a7��%�6V ޛˡ��ʅ �+N��N��G2X�0r;NS�R��W�b>� Ǽyqo{7��'��Q��]��t,�g;�oE�\�L[�h*Ç��lo�g��QO���(^�Z6M,�[9�P�v&+�GVHO�A�}!|��L[��[�㞗uI{�W���W5�n����� ���¤j�oMX��6*[신���A�H���b܈�a�{q�'k�q<�sW	�17�����2#2��p����#�.3�r��{=�x�j�&��q��(�^:����jY�p�|��ب�ɑ*���n=��'ގt'���+k_�+�w	�,8x{-�Ԍ�5<5+ӎL�B�ͺ�H��'���<�)�g.>�wz�/��9%�pz�̵����v)�ʥ|�D���8�i�0NʏL5o7=�;�8��K�$p��_T�}';/#���ӿ@+���$�m�z�Z\6)�s�|�ɕ�;%����	bJ�[s./�Qӝ�{B���N�(jn#��*<��O���_�DfL`��,
�DµB"~!P��MM��O���rUL:N{}[����݀�U�>o[��1�v���Ȯ�ѝrpR�	�k�E�!��ͶU�qsY)ݛp魰�@0�:�k5�g����,F-�ɣUL��1	��VS+e�JL1�m͚��R���Q�����z{V�$%]�LF6 ?��G� }��.������ߣW��2��]�/@�_Z�!A{ *��\+!F�����v"���H��*����r��pg�_W<�ey�IX����N%M����YQ`)����YRsូ������7�^�ܢv�?G��6�_�u���9[ӫ��迻��"�Z��7�`.��V|P��2Ϡa�uk�k�9�-�� �h�C�u|��ǖ~ʩ�U������'��'��Lt�ү��'����+Y�O��+����W:���V�Jl_��#E��辬���Ÿ���~!�+;K�N,�Ϯ$��x�ѝ�f5��>�͚S�l�f�t=~p�.�bO�����^Lw_����̾/a������Sw��[X�v��>�v%����
��թ�����Һ��û����'��~W �qa���5V幅4对��M�q�>��"}[R����j9ʣD]+���v!>�. íw�r؅�u�	u:��gcs�U�S�3c ����)��P��1��~zv��i}4��]�b��%Gu�{ձjR�uBll��9�U�%�6� u�r�r���P�U���<���#�B�t�C�P���M����m�� ���ohB��xޮu�p�.����S�B�s��C���̓V���]�-���
�J[����soMM1���e��ס��)V��|����q癨��4,�������@}���󴗝���7�F�BOӰ��J+��5:z������V����n�'�OG�7�c~�r٤��d
�f(ע`W�u@�f���%`0a����X�ۧANUG�/w����G<�au�*5򵳚����q�ɟ	���`!N��KS�x;d{��+�f��W��\T��`����������b��~�pT��P"xI�f�x��gh�i#���9N�
{,qv7!��2ذ�u�3�$l��D	 g�����گ-c��BR�B�����{)�M�CK���E��u:�L��Na�!ՙf��t�K�O��?u�T��{5�B�h!"���a������e
��}pH홴ﺤ3��$}4�r�B�G}����d�O���9)F��f�i�Xɟ"�1^�B�oa��������>�����I�UW'C�;=��Hm�Q��[��~�Ͻ��y���rgB��	n}S�N@r-R�d�C���|W��{�"ź͌�=��+h8X�ΉRvv<=��+>�9~����m�FO�բ���n�_V����^U���$e��sd%�$�́�|z�;���?S��Õ\4�C泱��dh���vfMz���x�#f�q�s
��F�N��/�R�f&\�/�v��`X!	����.��ê�c3&T_{�����=b����{3�>��Kdg���c>=}
2�Həb����|�]o��~�s�.��w:k�!uG�e�3�Dowc1,)G��Ӹ�Ϣ陌��sY��1��8ntJ�r�v3����f�R���l�׺Q(�	b�c��X�>�a��]JbGT��L!�u�x��M	�λ�v��}���O���qB�XM,E0����=�G�W��EԠ��9a8�y�G:�M����vf�&��A.��g��Oz�c���|��`���1&lH��bC鿪�!΃��Q>�"+�L["u<K�j�#�o���x�f}�ٚ�^�nq:P�ƅ~����7�G�G��\>y��?R��/���C7�s�ӆ�V:oF�V��@��fk����=gdO@��n\@Y���;���O��!?�NGE�A҂n��>V1��[�D#l΀�%;n���5��k'���n��}�~:�P��~�aɉ�(�ˈ|z��X/�f�)���Z�R�yG��zt�h���Pɡ�8�DK�����	�.MWl��\Cr��n ��b�|E���n"�����Y�/a^�M�!gtv@O蘉��-���mȑ4V�N�����6�1�q�-�ԕ"be�9�&o�Oa���}��]��F �;���n��TН�Ts"��$�`6�B�m}Ya�Hc���J�p.��c�]I:���b�����Ӭ��x.��sC��/N%wQ.���ؕ7�M��
���,�e�z�Ƭg��(��l�Vt��wWz�,��4�V��E����𭇀���,�<���H>�fzl��V�<H������,fV���ԺpwSbj��%�Xck>����*Y���ȟ�+���'}�o�k���␫޼Sw>�g��\l`E�}:������1ho�8�B�f�3�aDoS>'�o0{����n$��Q�ǅҋ�f9�Ck��1����
�����c�=�[3ѻMvu��k�v��W�t�6j/읉���[�Z�.�c�o�F|y��b�*�;0Øǣ&F<�5�t�x���ݸ0SO�_�8:{�Npl�f�H~�-���9>�z	Ō�P��Eb��q�z�8��Ϯ�Kq5�`�d,mc��z���;�Ns����Q�p��ц�>�w�3
�G3��<�ż>�Si�r�kYmK17�YPT��&DtБ9
R�8�R��)o���!�eO�L_�k�
���~]��fON��&7��B�mԘϜ��;9:*t�1\��"��]��}���=s��&�ˇ0`m���_Z����=�Q&+I����YqH��,�����4�ͫ5���/Rǆ�2�8��i�H"rɡ�
��U��#F�\/���Q���S6�n,SP謝sS�b�7{Y��
қ�Wǭ	N|h@���+�uթ|>Y~��>\��<U8��y��7�k�M[�2��O�Ǘ[lm�s�&��H�(�w ��$K�9�e�sӘ�a뷝>�yѹ�s��$��o�������{NbI��)L�t��4������0����7:~ɳ�"|q�'
�Oo�_���UٌGn!)��P�!H��ML�t�M׳�0�+wۭx������';���'D*�МHP^«>�²`24D³W3A�P��ݺ<Ʒ����RwC["j�7;����
���JRؖĄ7P?_�U�'ѩNw�f2�G�X9��b�]�^�E�rs���NM�t�(�����}j�m�C]�Ȟݮ"�[��'ew�'�����{5:n&�Q��*q���J������뽌��&{W[�g�Ѯ�j�5w�̟;���O�'=צpzsf�c&| lf�j}^���|-�o@o�k>���UϢ|����F�op}�vD8���9��`w�׽9��lҝ�L��i���9��EW�w[��e���>зm�j�Ĩ�ٟl�Zj�oZx5ЧC��P5���{�l�]�`r�"�"�f�b��֞˭W�1'͌�Z��Ղ)��r����������z5��ML�g�j�-�	VjX3@JV�H	���d��fι�6,���}�}�Ev��y%+Q�$)W΄��=�����O��K�;3B¡ᖣf�5�������֪b-�F���}h�|j��s�Un_:��8؞�1���mK�iG+��j�2X�����TG���� ���5�0�u"����ҫ��ؠ�옗�_gE���˖n\��z�+`QW�(S�ϻ/�9��3�jus��.9�%Z��W1&H9������ǽ/��>f��Bѡ9�V�W��,T�dX뫆gNz����EV�*���%W��iF�����s��g\���Us1F��c���7SJ7b̳�tȞWb�Lhۤ�/;+9��÷���U�*5򵳚��_�`d�d���
���Q��G�"��Ű���n{�Iص
o��*��{�pB��ө�;E��*���
�7񹉽�2o:q�^���&8�z=�g"�ǜ�eB������5W�ذ�u���f�r����s��dL�����z&)�N.���m�����e"�/��Էs.W�gՆ
�s��'b7���;��W_L�����I���W�<�蠘�y$�#��ur� ���M�t,[��.n��{�u܇`���ޅfk�-e�v/�܉�5:���zY�M�YG�ٷ�����^��gF��xB�������\�%�ݢz�˽��C�X%]�=��.��Pފ1�A{&$A����Vɱ�sHǃk	�)����ܮn܁�[�gK��m�����M��*4���l��N/k��f<4�Ұ�j�]З��M�ʹ�F�d-US�eL�.�^�pQ��N,v(=R�C�ۼ�U^����cʷm��3"xذm����
��ŝ����!d��Ÿs2��7yL�7ûC5�[��T������s_UoM�����".�U��N۳�ૠ1�DӮ7�����g+��G�5���K	[���`��P�Vmt��@��%B̶ A��!�JF��X6֌y�6���I��[]o�WKy%E�0�&���p���ڼ�i���&7`U=���J"�"�}���\��[�{oi����#�J�f��`X��ɣ���Q��kMh˭%^p�
ڳ�'2�=�+[�����y�x�ys��Nܜv�_nmm��:ʷ���7�h9a\a%f3�L�u��z��7Q�km�;��#6����ը�znÄ���b�m�Yu�Њ��˹��\p��h�!����ԥԻ�c�n��6�m��q9tV�y�ē륪����t�ZH�k{��D�(�����v�z���TP��3M�LdT���v3���,�.N�!L�X@m�\��K6����.ݝw=�z�|��Z�h���S�ۙY���­�X� �YA�Y\^.a�`s�/rc ��L� ҙmfc�.V�qj�QYR� P"�R|���w�gNb�)���:V3KTh:�E܊�R�iM�=���b4ich.�ńu�����
(�;ē�y&�7;�ɊÓ�8YZ՗q!(�G+1�����U����Nr\=s7Ij�+=6��hK黪�����֮gC���KtY�2
��K���tn��Ů��O�Ē�{�uDĲ�٥�^çb:�!+���0f��om��[<�.�P�g���[|v[�� �}��C��<%�+1|��I���N�e���Af�7�\�������͇�D��4@�e)^�+��ܸl��p1�zP&�K��j��R���&hD��ܴ �W*�qNF*WF�ٗc ��*m���tlvQ��.r
�ܻ��&�� oVZǮ�)ˉ3N޴6���m��'��U�.M,Nj��1O`z��LI��LV�B�K]I�����9.���E�[�U;���pJ��Mt�k�x�p�WX����s�VP\�=��v+^�I���TX-,l�kY��1S9��#Y&�)O�S�g��%
���t���Aw�H�Q�	9Fއ���<�m+y8Jː�˼9����Ó)+���q��ܠ+o�Ld���䒊}�&�hU��F�T( (���X喍mH胹�b��e�v�4ͷB��_쿫����rL���ss-���� 8.]���f㈓��nr�����~�_��3[Z\�6jö���q2��)&ւam�� ���B"ֳ�n-��Ӷȍ�$Ip�������Rf����6�m9�Y'D��m���sn�-�ɦF��n�H'.[޻�r)�)�m��ȥ ���$cl�謻:�msh̻M,��ˎf�ٳl�d6����:^���'qtm͹GCl��<:�k7q�P	�D��`ۚ[#۫Oi��iS�	$vٍ�i4��m�e�`HwM���ՙfd�쒰Ԓ��Mn����[9fQf��O�u��;0`�s;���uf�e�4[<f��ûX�p't%}�4���!V��a7	�,JB�ڛ&��ܤ�8��y5�%�e��B1Z��
�M�3LH��c~uA�v��v��9�#�f��W�߆^���d/a�]b8GSg�\��of�P��	
��; �u����3o�*9�3Z�k�MT�IvyQ�q}y�"C��~�#j��{����6%͙ɝ
G�%���=-�����wZ0�۶��@O1`o~���l`�L9�],9A����>l�D�;;~��W�"<�M�iM^x#����دb�jA5�+�Q��L��!�tX��|�c�j#%G��.����9�מo�L�m�7^����t�#r.�����`���j�70���Ռ]����5W�<�Mz���	�W�}[�ߣ���躖ċ�!���0���ں�q��fDm{���7�{��'��ŉ��/�[�m���@���(0�z4e�N��]B���>�����Y4j�������{	���Y~Sz�����4X|��b��8&LI��;ć#��P�e�zav_OZ�ɽ���J`�c�ؠf�[3Q���4'j|�ݕ���L��D�;QOáD�</*��m%=�^���y��ȷc���,bN�,���Հ��]yIƾ|>'�xV7��'iw�Q�2�r�PN8�Z�`[��eѝR�|2��}�F"vP����Ŗ������?�ޜ9ӛ�V�k:�_,���l�3؅w^����������+�Ձ(��C!�ϖV9Z��5j�]#t�@��هz���"��ڊg���踿}r��G�E��@���~�
$9P��;�^�V�A��!�Jv)�R+����8;`?s)���gDxO�P���+��迦k�B�(O����a�P�\����M�A�
TE�Nw��.�t�3�yqф��
tD�
���!P��NL���츆��7�/���z�l�
8����}ܩᢵ��3����U�E��V��hlJ/�Y+�|������pVm>+;u�O�6�	� {�<=�����6:*�����"�WQk¶�ɨ]"#���}��ݧ��/�`�r��F��F7l)�=+�{��5�L9oh1��轮�q��j]>Kӗm��g������D���"Q�~�{5ϳ+��~ˍ���WS��\�.�3���s��?�e��~P?�ʗ�q:��xT���fc;�oE�\ύ1n=��8}w��~��>#��s�W��{�`x�i�s��1�*ؿ��B|*Cc��>B,�ٍ�ͪ��~j�j�b���f>M���t,.�m%Q�,����,�%u�۶�7�j�a�}{n:l�ȾѢ��ô����PU��݊���e1��j��J۔n�����w�u\�ב�����ݾC����*GW_	���#�d)��1\wL��'i9�E����A~D3�e��,�1�����n�)��w������4�}UV ?L�bw�.�qw�����Q
��os;��L0C-��ꓖB�ܿ5��6���=Zdd�܊u�t����#�҃�7y��a��kȲ�}����>؇�b����3n\n���3Y>|���V��v*�%S�}h�,�;��D��H���A�)�p��{-�Ԍ��Ԑ�Z�ƧJ ͺ��l�*_N��y���XR%��Uj|��迩
�=unZ��/��`������I��fkȭ�K�Lt�ޗ�Czp�@�	I������N}�y��(�z������������{�̰]';�������v[M�"~��:*c����#�)�̫�DV^�맱���Xv�B�!س3��W��pvcۈX�j&�Z�%ñ6�S��UF!W��{|���fs%�*�����'~�_Z�!Ax����\+!F|xx]B����7&t��==4�t�����'�Eի�$x�3��%��g�:�J���A�ieE��ՑB��;�)>��\�j~X�;%M�. ���k$�(��FVb����ڼ���H��r13-�9��ʬQ<s�?P͎�޾g{�p��+a�h�%)r�j��ʱ�VV�u3y���8�qŬt�2���g�����l>�],����\.L��GO#d)S�V����"��/}y�W��j�\�ޫ�BLT!�qu9�\�
GE��������`G�W�ue�'l�R��"��M�j�����]���U��~�_���ǖ~��d��#��Ȏ�ܺ��ߜen�jk/�Q�����؎az� �$��p{�\�/&�����	�Z�����6�t�tɠ�sp.����w�+I��WӜ_�P�F�����5��:-��F�����V�mN�OL�a���
����$�A�B��S���4��!�kD��Ն'��q�a�T�<���l�F{��]�Fw�t&�XE������7���w�5�Y�Q^��}S+�N}NϏ��b�9�-�)�-s�����8��+�f�'�Ki��u����L����Pu�SW�e���^�R/�<n|��)�͌N5/�O�U�k��ݫk�0'��˭�W_�l
!_P�)�gݖD���1J�W;��WZG{�d�+����#����eߧuE2�Ml�@�ؓbz�ɍ�@Ⱦ��ft� �˞��[D�����G��=�aji��C�)�3�ϦA���b�z&1���f�a�U���^�S����-��.���љ�Y�2��2%�8W]�V���̔��4���#�;����7�"�#`̳�6�I���r2.�J׀�6��Ʃɽ�&Ѫp&�ZDƈ���ɬ��šp�\[�ɕ7C1"I��ى��hd��ӕ����ڝ��"�I'��ǒ�fP����>V�ѻ�ە�Z����A�\G�ul�G_T�$��n�QJ���\�=��b�2Z���B�<�c.��9
�N�o���b��~����rcP�T3n�Oq�f�N��dO	PaԸ����<yX�B�nBߡ���A�9�9"sjNe�>ޮC�Z:Td`��MD�B�LW��R�+��:�N3c��8+W�c֧҈��xF��Z�>x{@nY���*��Qc�^�ɚy�.f�bEEF,U�r���;e��Q��U�b��F8�A��h:f��_L�n�Aj�;g�\�٥��d�B�1^�W[{M�E�m�5f�ow��fn�/�0�g�<i1!zX���#C{~�*�^ұU���d�|j�L��ME���
��)���Xۥ���3�%]7��8�z4.��H�]�g:%I�����ڔ����[��Y������b���Y��u}1κN��@�1Ӡ��/C��x�dY�����>]��=�^��X��;��K����Z����@��9���FO���2� J�r�r���5}J�=;x"�qB8Bck���Jʆ�Ml���%fԒ�����U/ 3�	��&��S�`��2�z���F�y��Z�7%�q��;�Vb���t3,	��8t�
��iS���-��}��O{2��(U��S;OE`	]�7�����U���聗���\Zk��g���Xf0�Xf�3����fr*[/��HC��B,�]F���u]�q��c{Ns1��Pق,b��hߔ�϶j��_|��A���@Sڵ鎬���r%0�m�/������ӛЕ�5/�h��)�����9>b���'�A���!��WCb]O<�i{�]ЋR��V9z{- .�5S3PW�ۜߓ�>k��XsS1�>����p�����5k+�����9�Pp��9Xe��}�V���7AOY���w��LS��'|�,ֈ�b�IY�~���"xI�p%Ë8F��<�k�V�A�Fٝn���儼��Ew���A���vOP��Hi�}�.�O��Q�'�V�q�Z�`���	��L��I���{���vg��V�V\ϑ��8�V�\�
D�
p(MWl��\Cr�xJ�Ǯ�B�>����}TB~o��UvQWu��/CbiT���0�_	�K	�1���S��{8�fr��K�����Z��4~n�C�+��������,B#���;�Í���������M��k\W*ᓎ���'
�X�UB����o0�d��*�%c���"NLE9@[�韖5�\�B���k%p���.J��'l�Ϭ�8u�uu��Mܗ�,�keܘTܜlV	�i^B��UBÑ*�	ʏDY� �>��t��Q��'yэ�
��^4M{�W,J
Xo�ϋY�l�K��fEH��sq���=zH>fgjuMĿ����JE����T��]t�\lc.��к������[ٴ�C̿[������:�$Oul6�*{VD����R�G����u�Cj�.ab�y���}���c�p�Q�śgE���#}Ӏzsf��hl�_�*ذ�Z�������|�dС���yܻvg���/�k��-:p/���tW�ޜ=�9�Ϧl@~�-����*��TP�����]����wTP �_��ӗ�5pܿ����\��"7*��菀�\ǡ�["v�;���9�d���HE�E��ϕgWLo=�u��W��^B�j\�Ȓa�D�:�o,�[|K�z�=Ĩ>���`ū�Ԍ��Ԑ�Z�Ƅ�B��)C���w��d��ڝ��Y+��Q�B��J~�X:ls����x�P�u��S�S�dNl[G�y�99�RS���Nqz��Q�'G�LQ����������9�9�6t(P����1'aGo|+8k���ٻ�݋�(�0lN�=u9_V�tUb�i�6`���q�\g�y��w��=��r�BfK�v3,9�*��V�9�'�!��
�"P�m/��5�Nk0����@�$�2vg���.��T]��r��#|{ϼw�A��? ��e�Js%=�~ʈ� k`I�l@�A
*lT�K����|�׳Ɩ{����."���L;x�&��Wղ�Wf3�v��0�����B\m�2<�F*�w���}�03��oe�Օ
N}�b#�[Rw�U��)	x�Ϭ.����Etg��r�m_/rkɖ��/�_�n�N�W�[�K.��R��%��,4���������ӏ�Ǌ��T׶}�ۡ��j�Ź��A��[ɹΜG�pt_w�DVZ���AF9"fl睎�ޣ�9dƚcۙ��8�We���t�0����u<��t0E��]�.�x'���ؼ�9�-G,5���8��vD<�~��k�'����,�Һ�BVQ��G���<~�_���m;۪6�ʋ�m�>���R3�Ч���
3[�s���|�{ӛ9�Jv=3�t==��v�Ƥwoi���u���U��"O�����`��*���2�!���8��Uw�цv%�Y�,_�TU6�#{�L�ds��nb=�t�<��, }H��r��J�r�����6�����[V�`�rV���딸�v7/ROo�cEs�h^95lyef�2�M�.4��"�ۋ��UY��i�n�YQ1A$cN���؊e����[�
, `9(���:�.X�Xj���I��{��ڧ��uo�R�Ô��q��7W�^�.X�x{'�WX��_o�DlJu���Ȇ��[N�/����ҫ�}-�
d��s�v��vr1�ŋ�^(1����z��[�'�)�g�DGX�Y�S�s��6��mw���y�x�S�8e	�˛���lI��
�:1ub�2:������P�gf)*�|��a�q�7�7Κ�_?X�w8
v�賄�?�$/r�E~�5�(��?r�ʧ=�(h����wK�
o�ك�t.+Y���mʍ�򵳚��Py���ul�G_T�/�o/8d��-��w�':lTÔgT���,��`H��F�8;��,u��N�]���1�>��JԠ�=67�(�扄m�l>�����n��O�s�0��6Wp�lC�Q<S^�1g���7�:��y�<7��9�aw}��9�R�Z3r�c�aUt5�xC�w��U{�ۙhh�N3<�{�!�9����T
��ԣ�o�iZ��xr�M�p�v��J(�]�JS?c��v֋o��X�ۘ�n��L����eh��n���[�34vcxjrp����w�����˻��\����v�mru֏a��7z����v�l��{R���n�hn�Lk��l$�A�`X�����47��a{�2�-��{�w�e�7��8�Q�-�01�.�d�b�t
���a��W��i���w}6q�0�Ʃ�>�}�{};�p�hh��D_�~k �3,=¨[[��hi�˚	o�Wv+��5�;m4��7��6&�5�6��G�_oJm������������!�}Ϸ���v��;^,����u�@WQ���D��P�yze1�LT�:����2�xb���'��a��Oi��rR�#��7]bs�@�Ɔ�0��7�i�P��x|�7^�eh2;Sֺ�}*U�i�#�ֱT�I��J��"=�t/3v�+�9��y�S2��\%K�s�����R5O��v�SC�W@��z(���^����8���*a�u[~x���]��K�Yx(�p���,��q�	��G�����C������Wu��డ}ktT�ݬw<h�_e�oe�qvM�PH���T������Uf��h*i]�j�г��$�i���`�^k�kwjg&X]%�����zz���� 4�]��l����L	�66��K5�Q�N����-B�U�-����L|�5��9��nB��N����=eS��A*-�@�d�]����=yI]Ŝ��ㄗ�oϛ���g�_��z��(oof���,<�Ւ�\��9r����5�L��ɻ�����W����k�ۻ���M���[x�(��cVBk!u8LGfM*�Y��h���Tv��5�H9m��zIGv5�+3�g4lwզ��:���=�ov��ط�]�0��+6��{+�r��r�LTDu��*����:���o2����\Z6y��˴�]s� D��WZ�鵑N�6x��ap���w7]FS�a��ں(��1]��F��$�����v�)��ݒ4\-z�В/p��ܻ�ī����3Ƃ��/*��q�6�r�Zaz��ȯ5���1J
Y�uF�gV;Wb�v�8�vpD���,V�kN���Dfm�����6Fl0i�n���LJ�dx�`*��xvkŊ!N��6}�(Ռ��y�����!�_5t��<�2�˫��GZݺ�|���%ۻ�A'��jzVE>��j��K`�[D�]�X�������b�ΩWZ���:�f��aް��.F0���NN����W#b\�"e�݂�>-]\bFVA�����S(o Y`��b��g���G�t�.��w'>np���\5yW���k������]�差J�:�תkJ�Q�����@�hJ��E.��w������DF�����b�̧V���D.-��E�ϫa���0��ʆ��6w^T��ճ9;�K�����:Y�e�"fb=�����C�\��]v��,7vP��!
l�J�b���v����d�|�aL`W2��«���F��Ѧqv/;'�LIeZ�T<�if�3�q"�.A�}�k{���"�ydF��tq��ae�C3�'S@��d� #W|����׹�q�k�e�,1�Y�
F��ח��}V�qi�x0:�]�բ��]s�F-,�cM+�����F���u1y�����;
��#[ϰӽ��	&��-*[%#���KC@"���oC�lv�D,��5n%��fp�̬���,7��M��9����i�w�BՓ�o���(�W	�N��4hG66�ڶ��e���k�9	�����Aʲ�����Z*K>�����j]��v�)ӱk��J�
���笝�v�v��f���Щo��O�*sP΅���7�:P�团f�9���"4���:��%�`�f�dN7��K3!*�ƕĘ��7�.wc�)ޒ`�Û2�f�M�OK�-8��x䧆n�Y�)D�[���!ۡ�!�ڕYTT%�xe0�F����^]�}�+]7' .���2�<��:�e�ٝ�*j�
-�^��Io�����������H�33���u�6ٝ�Y��e�giAc6�Y}}��_��?n��W�zy)�A�Q�흕�ٸN$��
[vY�_������w�%ncLC+v쭶�	A,Ĭ��Z��m�nuea�i͢�������Y`�'m�/=���gkn.��ee���&�k9�g/k��"����s��B陵�gvgE�7l�.,賸����vw6���9�D%�VYܶ��̸���#�w�vt�ȶ�v�$]�u�m��6�m��leVe-���8A�ee�j��%�e�d6�qř����fÒ���8��+[M�K"��4�-m��E3q�`F�\�gMjm�\l�ƍ���F3'Gfl�\���:�ghGgem��@W��_R�o�T�\��eV��.�M�׏7^�E:�:��i��Fޮ��,����m�� �����n�La��6���%����'W�e���*?EpQ_1ƾ��_޿}^h�dyN<���L�|Hx��/q�K�;�,cv��߸D�T�8��A�A��9	xO��Uy��WZ��}��*д�Ҫ�3�
�W>��
��m�6�׻jj���d�}�Bl���lX)^��k�U<��g38KZI�Ƶı�`t�;���UW�'�˹�E/0�oX�{�F�_z��Њu.j���I�������:�tCBt=^�-~����6�~\�ګ����r�0=��5{���[��̗`uİ���T6��ϛB�Gӣ�s��f`�O��P�q���{=�~cy ~��Y��������o�.0h饢}��{w�����-�fk��k
M�߭�6��#&����v���>�^�y#ѽ�E(���
���SM��ͤS�=��nK>w����W6�[�],<����.��� ������ܱgv�C��[ܸ�gK�k�q���5qY�k
E�-�N�m��Y�O"��n�;e'��|�E�C}�uZ�'�V;3���2T�ӽ�Z��=�b�Z)QtT�F�[ۭ4�V���}@��N=+N��b�or���m�c!4}���E5�}�i=	���ͫ~3��A�=[�p���sOOR���d�z�����-`]�X�������+�=Ʀ�9�b�>���ҾN�.�t4 >�$Pヲ�ύ�|��ޫ�q��v��m"M8��K%���^}k�ֽ8���%��@�BC㐳�#p�٧g�%�@�a���>|_�K/Π��}����  Ą
�]��=;||�t�����>x��M���]oE�,h����g2/_f��0'�т⯇l��^��W��#���S��#Z�%j�;38I�k�'�rQ�� CΦ��{���ڝ`I��b��QZ6�6�s{�ɯ78äc�VO_��sL:�<�]-k~8��I2��������C�k9�������^ ���wՒ����:��Fҷ���n\t,��<*A�^�Y �GY�ꫮ9^�HR=���,�RRrq�S���NmX�/t�d;��j����]��33�ȉz:͗EoOT���V�&���7L���L���:�)h-��]0.��()^iN�Ш0K!��b��Z�Y������:v�66���-%�.�)��9A������ߓ^��c���}q�n��_���ٺ��z�{w1��i��W_�a��Z�|Ƕ9��6�4L{�c�!hI5/ßZk�^=S�i)��-��/#}�,'�[xv�|'ۻK*K{��u^�^�^��^N��ΐ�)'����o���}.��{{xRq9�����v��-I޿�rU��E6����Y�>����5�y�z(J����+�F��cY����)��Y!!�O}�1�J�u�lm����!��V@�Voj���n��;�{���rK�=�.�V���_@f����w���!%���uo|�gݿ2��|�#���'��^��>�W�q��jPy�!a��#���|��H�#�m��!R�g�W���~U�J�b��3�e|�B�y�ͩ��S��;6�w�<T�؞^]�ᾥ(��5�ͪ��퇰�g���|3Cf��f
ڵE㬼=7�h ���9|�;MfUb���QW��ZH��z;�������LX]�f.��N,̤T��M�ol�,�mfB(�F�W
q�;���]6�Bqnob�E�śL:4�Y��>��G���5�WygX}`�GZ�G#�{�6�u�vexi[:���[�]�͎����D�1 x5SOV}^\ޒ���Δ�#+�h�u��ds����\-�[1��T8i���?,�����s,��OF��ޅ޲GEb}��oA\���{]���dЎ��3��c{{XH�c����ƪ�g����a�ÿ��9��½Z�S��~�X�oP)T�c�'��[]��஬��X~���I��rGG�g�攫�I�h���!�$ v��{`EQ�����6��
��9ީ=�]"�iM��)�:/���6�>�5�i�E6<;�A�ѐ&5Ue��~�G��zY:��\�vȤ�g�}���˰}�{D�7��p*4K�q>�g�s�7��x���*)q��=m_͔r{M�ܕc��0��#8\"�z����۪����Ɲ>+�X��	"W�T�����W|2������9u'Z�{gD���&S�x�&حC�0����7�*���j�ٝǬl�-�i+kE���j�-ђ�,RP�986T-�@$Z��՚�����o�T8���
N]Qw�����"�Wu�:���۬�er	|���:8wP�.k�[�S4�q���x�e0���k W�p��������w�����݉��ի+n��b^�8��W��˽-�߆�o<f}ŗ��I�N�܃��^����oB1���~8=�z��8�mj�kZ�����nmoux����i�|�"���X!���c�	j�a������t�3��m����>DV�&��<��h�J�A
'���#��[K:���NY̵���`���ۏGtp�}u3�
��\�;r�h����Bw"�n��uO�u����A���Bl���SK��|^n>��:����X�@@�!���[�w�ÿϻ��-Ѓ[�}���>资��W�:�ud��CZ<#���wְV�_ϓ}��[Ȉ��F�*����c/�o�\�O��7�ĵ�J�K���|$�(����;W��-i�J�:����HQ�jPq8Ku�D���ԍ�*�&3�5Dٖ����^��>ͬ������yh�2*L��D��bOr�'� �QT�l�i�S�I)����K�-�ٜ����pY5��]�x�y{���ʻ�Cjh��Wr����8��=��^���y�3��.��m�͉-��hzԹ�n'�
Y���<�b��>XvbYE&�y�O�lw�^l)��b��ѧ����O��ph�����+���m�S_6���
K��|�o��������Y&nu.��!�%6s�+�N��5�i=k{��(�@�u�d���]{��i5�z���BHAP�_^���Z��sw����\�L��huϴ��;�zM{�>*�.M���]�@�_@}BH�}v�ԅ��)2.M���p'��[�L�w�s���f�rY���0$0���C��9�gvs#=�|��3��>��f���)5��З��=K0xۓ�~ ��]o<�q�����{0u!"Ӱ:����KD�ߑu�UGV �{h���O��5*j�����H�b�v� h�s/ 7\J�7�Z���:�5��/!f#�hSJ�f��zjQp����R�E#�[��W�K8�m�*�y�D��i����=�`i��&A��N)����0��l�V5i���Ǟ�|��7Pw�F��m�E9�)Vᜁ����8�ӑ�	�L�H�mp�!~�®�<��:a�s*��W�$��_f�TI	��٧�^��$��:��c16�zQ�[�if�0|, �Ox[ެ�����������5x&�FzE^���C�`��7C���$���/5�?1`�+7M�޸��0�]n⽪�yf0ׯ��o�V����s�:�e1���i�ע���m��Z^��{j,����ӫj���J�G�.�4�~ؓ�YH����m���}ѻ�K��Z�<Մ���n�_�vs�.��P}},'�[y�n�
ef�Q[�bt�J}�ir��g=�y�4;iRb)��B�*���.�����r
�C6�Y�ɟ]^�q~��fOi���r�(!�%���C��Nל�MT���y[2��>2F�x�v�
�[�f��g>V#ޞ���ch}(>��
�OpYV�G�p��yށ��-�m��f/��O�v�#��"��)֜Eo1��� �e"`O��g.��x��n��d�훻z�p&���e��i&7��A��p�f�֓����[�"A!?�����/5��L	;1���	�5Ce�F�e��gZ���е��|n���&�*|���q����#�<�>̐���x}1�����Ϣȧ�]�P2��?f,ͅ���z	�~�aTE3'���5s5�%�!#���;�|��a������=�K�=��AFߪ��Yݾ��r�I'�-}G�:7R9�6���X�*L��>ĉ�q˂��"���8d��/��pC��}�İ�J�v����zVq�y�DpR͊�J%������|�a��J�|1���5�ď�M=S�͌�]1��{0��{�7��
	���pO�SAp�f�zc��T8�o۴�O� ���v�����O���E%�_�����d����$ɘ,k�ƴ�՘��}�r��;�Y=�B?����,6v>�����z�r}�5������
��5�ጁ��u������՗��� ��N2�if`�;"dP��C/L܈'u��n)�k#�[Z���ul�6�����U"�� �:��.��W{/	(b�˗Թ���5���u-YLм����(�k�n>}G8A�{�u��ٽ�s���u��86�Ѳ�M䫼QOe��Φ��Le�B@`ͣ����/�Mی>>��C�G��}� yf	^ڧ���4d�����"�4��ش}g�A�����ڒ;ݙ�q-�ߡ�x�ǔ�%���/l��z��-�T)
qYuUx��g��<PE�>�Iq��ߌ�l�g�؍�W�@F�x�����>"}�G)�������k{׿s�>��˩g,fx���E����éi��j
��po�X&��X���7����w���'**|��_yE��͓�yx��d���{ y��%���^��GٜYy�:�i9Y1츼�'Wy��t��ݕ�1��!��#1О�'1��|�=���T/hW8`h�;�'Px�r
=��m�a��T�>���R;V7}��R��{�`��&�/�D��-�m/���"+lk���ϸD��ˎ��U���rg
�G��X�|)�܊����(����x5Xu[q[�(�T����"�yW'��x��!���u #���yH�f,b��x�����n]�nm�-C5	�m�7�:�m��A������(�D��}n+j/��T�A��ub,�HB-:;��步A��V�h_�[eT���|�Q�w~��c�ו�m����#%�4����4H;���RlXiLy��+�-M�^'8�Β~��_ed�����ƪ[���a߼>�lO-a]��W�ɓ`�,{���-�}���!��{ƉλՋ�=�n��U�]�s�W(D��os������U�]q 0�D��h����i�)ZW�Ivm�x��+2B�[y���L�g˽�y*�͉-ʪC�r3E'7��0��ƨX�pg|���l,4bZ�rӾB'Z5�s����ǡ���}ВZg�=�p&'�L3���i__m�����̈́�~�J>�x'ͦ�Y��{I��@���8����k��I�cM�xͭ���g|sY�`��_r2��lC��%�=RC��-.�\���81u4���A��mj��_e��)$_w(�����a��Z��î��A����u0�L�	��ȭ+Хu��7J������	G�cy> t≾�u���:����U��"N]�q��/4������c�6�y*}�g:2�]��v�E��cEg������X5r�9z�hO�KL�)U-d\�)�5J5!���Nc�k�FbY*A݊҉�g[ޭܲ����������� '�9Ɩi�Wyc�+�����YQf�V���^
H(f,��wԗ	��f�����s)�8P��5�W,�p\qqN^�*5b�3(�d�-i�ru^����I!�YK��V�k9�d���Y9�F�&����@�vXpQSA+��c�����er�b�����칕�k4@�/&pI�9�]����T��D�_0k��N��J�u[19�j�M�Q�J���&���l)�HF�3��6����A�|�k2'�h�ƍ[X%�N���j�*�-�����q���-��:���EX@��own��|eLË��s��S�
ve-�5�	�1SwF��|�Rջ��f; �vY7 �Y�sA�d�>f��T]�n����33E��5T�Ab,Ԥ��A����]+����K�Ç�����[��*����ln�D,��dd=�EՀ&-h�jɐ��s7$���(�18_MF�G���z�j�ջ
�e��'<ބ�Z���W<����c�|f�H������U�P0V�yW�. ��@r��v�ܬ�����n�wO���8`;�5��Iv{g;;���X!�����s�Z�SL�=��®��-
fn�p��ٺ�6l��q�-n�+�۴$�d�I$
�;���I�V:X��Ѥ���%��U�������=k�g"��t�;y����v�|�;l�CN����K+�(U�]'-��b��s���Ko�/ fiՋFԫ1�%��R���Q������ɴ�Y��WR։dg:B�J����{M�u��p8�ڏ�|�ŵy�|}ywn춃��r�rՊ���A+�K�FcBT��̋�.��w��,Pĉ Z�%$ڗ�k2wF���CJ�hjܻ�̱QoN��Ӆ쎏�Zm\�Y�6Nd���X�M���E���r�,��aQ�iX{4�{ύ���M��"[��]�5�Rv�+5`k0T�7)�<Cf�*GF�{F3\��T��b��gi�6�]�S���
W`��*�2u�X6��x��*,	�����-�U�Y��oL���'
���<'j����$���0��@p��&R�����3F.V�]���
㙀V��aᑞ��:��r���fgY��`^���*(�5����e�j��jb�xq9����U�ٚ�%سi&��ǗdѶ�!
����x"�f���ۂ�J�!�Dūڦ���t�A���]۶.�3��:5-��4�Є5k�҂�`�֖fS_x�zi����X�_wmR�c4"LJ��j�(�I0�I����b�����ie�f��YY�]�m=���)�kt�me�����_���󭛳��VvP�m���.�Cq�2�졵y�^e��.:�����~�_�Y��,*Ӵ�-)(#+
JY�mvE���3vv��i�+�΋,��e�8;�N,0����ݪ�$���Xfskm�eۍk,0��̺#�˲α'{zy�=��΢��+f�ˋ�2�$��f�Y[5Gq�Z*�2Ȳ��vQvu�vU�wYgl�E�V��qݚۺmq���ò�8���Ŷ���xyٔA]��;�n�,�+;������N[vI�Nq'֭�Q�km��i�JmƎ���tgql�NNBfrYۥ�v���kX�{9Ğڃ��&�gC,���M6������������� �Xd��y��K-��xb�F}����{��K�i�����QX��U�%ی��Z�@o��}glP���������t`�W��5=m+�6�ȯ�GW�4Ѐ�㣮�g��K��V��^%��s>a7م�/{��k�k��`�l@@��������sA�����zWE�[�]��k|�y�E�һ!�Wݻg��O��`W=1[��zae�$V��"��;��X��M���������:׉�%<�}�1��f'{=5
�%�Mv�����g����Z �� �]��W��J#d�Ӎ�6pA3%�Q/V��߉���)���b�z�{qp9���6#�B���V�o��[��q?0��[t��Y֪\U��]��㊯=�5ݨY>gKM��j"�n;��W�4��o}�Q��9� �計�.���}{�@�*���z��cx����ע���m��y��rM}�{&��1���/&��W_�$üi�{m{ȁs�\Mz���I�=�B�q ��f7�{~ڽ�0~���L^�Z�	�9���Tf+x9�Ń{-��{�jʫݻ�r����q����t෺��ٵjǷ�K��ի�k����hn\�*.Qv�c�X�O���8]l�o3�w8��]Kiv%+4��c&D#��T��üA=��_-� ��4S~�ذw������a<[y�n�[���2;g��o�q�I��Rwo�˼ؠ��6�gЁ�މh�H����RY�K�G����o0Oi���3��aP���D?Btl��)z�M�\N��x��yh�h�6W�'�|�G�=p6Cl �c�*6�Ͻ��q;y���(���hal�����y�Գ�Y��/��{{��W��;$�����N�ݢk(�>��,ͭ|�2K>��8���h������U\}p�cM\�j�]��mb�Kٜ[/�ݟ��MG2�]{��\]��&o.�y(>�ǲ�{�w����sZ���,jS&>쨋��)^�����#ė��f��N6 ���O��J�,���R��ݭ�g|Nm%�b�^��{����>N��o�:�x���	����Cyuh���f&1�x��/��yu������5{Y+b��+�VM&l����9���U�Իb�Ω��nH��{�1�L'�mmum��/S�Ɂ��h��@<�9(�0�0��7�J^�Z��o�c�絳H����a2���D�Rt����=��z��`FȲAVSK�+��J��'�m�L����0�^�CJ2u_@;�x�:+8�-�B��c���D�B�3;\u!�%�5�S�v��鼰�}��X�j��6|�ðޱ`6v	==tg�k�Cd�Z��[��=�쇓P#����d����R����g��s@�8'g��3��\d��>�`[}�;���K��CtJ��"��~j|�}�v&�������]��86P�������|����96��DE�h:Cl�Ƒ����x^3k���<N��).��"6��i%���]��^ϙ9��gv��:�F�D�#�(:�ep/��"�:���ii���6�(ǳ�\�8��K2�#��̍�vp�@!�jt� ������2�eh2��<:ۋˑV9{_�|���_I�sJ=�=�wmg���||�`���q�w����E׫����`�wx���M���GN���7�H§��j4��dFX���
cc]��n����]f0N�f��(MjUi;P�y��;��ܲ�x,��ŏ����{���\,{��rU���*��:$ķ1+�Ұ1)��l�����M����M���i76����\�C2o�*�9]?>�y��{�z���Z���d[��"}(_�{�����g��u��:�@��	��5!5ԏB��{&{P�gx��ڑ��q���.]�$N=Ҷ�b����� c�zF��6�r�܏<�VŃUt����Y�3~��Mq弸D��u˝�4w����"����{�-�O^XEg�è�J­H-��j�s`���oAm,@��[M�Wz6�A`A��m	��^����k�{P���1}m}<}�w�=�m׷�+�k�A��+�,��Y=�x5P��o~��c�ǖ%�ED�Y{S�*�"�c��5��j�/�%��k�Y,�`����_W��vm���{o/������t={�{�k��Ϣ��k���J��{�U������k�#Qy~δTG����7��F�X{Ŷ��o �w0���ʼ�������c����8�K+�;!���	��*u�H�kv#{��UѬ�ۛB���t�=�*��y
^]�o:��dUB�<�Q�^V�w+��ؖ���΋��	�:.�T���U�����7��ĎC��n�s9��}�^����y���k��U�#�Uy4�U�TP�Z�A5�������������a��4��ϩ��>�)�wL��G�8۬��_\{�W���v�ү�6�Ц�{�M��/��/���a\9ڶq{�S$mv|�\8�8��X��ZOk�JZU�8z�U���Ħͅ�<{��pj�ǰ
�k?v�r7����T�Pk�á���f��J[����L����GTw1�t�<�4��n���.n6��45neu�k���MM���^k��ק>Bb���C��>W�	�/3�A���RLv�X��K��U����Ｓ�ܒ�W�M]���ם�&�W��@A����G��X�_x�R�"_��~�Um7�6��o�E�1_#ܗ��� vh(n��8�����Do݁���u��B6��O6��(O^�G�ޞ���#N������a,<�d=[�_�����8�d�ى93l���P��]\i��g]��<�їE/f:��1<�R;�u,=����oN�eQu����¬ㆃY�V���g`t�ʌ�����t�Vgb��݉\���D�Jt/*�j��<���vS� `r2wT��i� �xh#�~��.��z=2|-��Y&�Pj�Z�lSN=�-̔3=�Wh�m��Đ� ����-D{��w�VJ�^
�v�=�����5��6kL.���������J({mz��a��J}��0Q]���A��wl���7������$ñ�Z�q�&e�g�էަ�Wu�4r�� Ge`���my؝}c���mi����:̘�_nl��Tg�v�H��}�|�U�ŋ	�}�C����|6w�l�&�^�P[�U"�m�w�{�3�����mKb������Ccڭ���W{��x�,�5�;M��_t�H��J�=��Xc|�\�j�Vh���K���0�(��Q:��ͺJ�i�S�!��ԋ�(N��>���T�P��KX��${����'�v��9��/��:۴�!�L�����N��ro��!k ҡ37�-�#h7��CHuq�U����27g\�!ʦ��X����ǲ�^m��xܳ��G�Z�Ŭ.��:ֺ)�c�ben�h�}�� f�]Y��[)JЊYNE�EK��z�l?�������cT�P�Ā�o�3M�\c3qb��K�q���z�?�9Ё���ʾ����X/f}ŷ����s����-`�#I}�4ϼ�ȃ���1�8�mo�ϻ��I��ҧ��#89.(�-{=|�<�b�-���JГ泯>LײLjz2��G��r}3���8.�����:Vc�pC��P�{��l�9�<��S�q���B���$�m"�_��5�����s��{I�Gُ�uw!�t-G���oT�W՚V�ܫ��&����ˢ���J��' ]uVg�q�|L�� ��#|.�R�w9�;����K�2��f���Ԩ�^]�5�����=�`�N�8��`f�\n�vڽ/���M���[����F�]���v�r��%��%f�>>�{@{$���ǲ(�OZ[z��R�I+Z�g<���5s��,#A�K�ىɾ�3��n]׷����)kڍJf��FK�eQ�O����X'N`_�6;�b��Č�'xn^TL>Z��X�=��W� Y{o��������z9AM�:�x���z�n�뻲�9 O�
÷�@e�n��1x�桲�nrQ��"���LK7  
rY�o����|uwCm�Si�D����K,�.gFS�z:�D=^s@�][��y�y�3�c��sS��So�?}'Q�^�%M]�v;����Y&n[t�C�l� |��^sXm��eo�-`<�*>��>�ZKƏQ�N#�� z@�rC^�!�My{q�>�����T.q������w���Z�/r��]�P$G�������U�f�_�w.�Ŝ��Ȼ�����`y�X-�[��9~�@�����3���#��n���F��M��[���B�o�^\�"m������B��1&��U�*2�y�2��Rwa_Tg��й�����3���`�o3ࢨe&���������M=9����z����h$x��_}���sR���8�6�|�T�����o�|֒��|	HW�h��.�\l�AL���3�oS�3`�gD5�3`�b�:N�L+�d����m�g�Ҧi.E>�u)C�yYV�����ݴ`�4��'N�`>ʱt���Q%#1���	0�ֻ����A��PZ�����a��v�H*�Nw�j��3��[�B)���`3��r�/Mɽ1(*�ƪ�����x�K/��1[{@m��{הA]�qv��|���~5�]Q?`%��z��[��ׂ(�שu�fn��3hy�B�<^��`�k����'�0\N@^��y��=>�r�׃�tJ}>,<I�x���dy��]��ޭ���g+n{�u#ݾ����o�Z;���e�|��&�SO�=.iTug�'��M�du}y��rP������_�m��)��EMK��8f�ͪ�VO�7hK��7��tHC!���!�C��\���̝��o%������K�^���C���A�D���q"���k�}�ԳWf�V��5�3�*ڃ4Zn�5�M����.��t9J���g�^�3����w���D�S�/��X<�?'�Y��K����Sk���-��������m=&�޾��H5"��oa��p�H@�����UR���.L!��2�GU%"䟝|'P�:V�Û�񀾱ԝ�(tc�CM��/SA�y��Q��Ü��DY�*�A��e��4Sܪ6p[Y�^�^�Yo ,��`,&��c�@���w��?:��gK/H
�h�љ&��Kε��{����Lo���?0�3�u����<�S�|�Ļ��[7��=��a��l�݂��*�~�a���C�����#1�Y�:�P7�OQۡ����pԽε�֕�+8"~��։��>��f����)+���/oRF<A_bO�l[a�d�4|1�VI��12Ù���s�� ����Ԉ��ݶl�z�>��B}�"ߘ��Vn>��ꋏ5�<��ɮ��2js	��2�3Ӽ
h_�XIc}�k�~�w�}+bxO���wZݱ�+�ֆ}>��~mW�����L;���x���Wig�^��m��X��ׂYX(�
dx�s��t��ޝ�>��3 zI���-�g1�o��g��e�͉�����}�!}�Q�u�t&���=@e�p ��p��w4;4�V���)�3��� va�1��; Yd�cw9�t[��ϛm:q�y1A�F17�x,;�Xq�@!�r�-�6�ֺ���7�oo�X���8&��;6U�Fve�'-/��V�%%s�*g	۷���ڳ[�)�xS��ꃭD�
QRl�g*�(^�V�.���Wgt�\ޫ24�/OyJ�����(+�G= ��fWKn��BF��Ή�$Cyf�N)���!^��K��B)�N�0+/+qnH���`!L�J��4	������8$e`�Z�������/!��ώ�̬Rc��6�VU؁u-k@n(�n).بc{�����E]� bst�f�y8���o���60�,q�nw��!�f��I%fgz\�hr�`+р:�u��%�O�N՚Z�e��	���[]w�G�F�M[{R��!2Ԯv9�AT�p�"7]6�\�u+�"�2�Y�Qp�0�Z�o^��.ںu���,��Oży-��۽,��^]����H���pe+�����0�x:޽yr*�w��0Rg1+1V�.M_���z��AF�P��������AE"���d�N�*7y,EJ(�p��7�q�����n\C�Y�[��/�p� 3	^�x�ÜOTKʷg"\�oi.w��M�m^��h��Ѻ��87u��C�-v�1ra���L{x�oI�!�6�G
{X�痶�/h;��Qr��:n����Oc��̍&�L��|K�m�RX�Pε
�������Z�r�{�Nی�,b�sy�yt��T3w	GH[����ouP�0k���vfu�.��i����^�7���%	��޶�n\]���b����_6���t�&3Jf�T��j�1�d��L�a2��n��cX��[�z��T��q�WE��C��Qu�{�O4i3��[�>Cr����БT+7n��6Z�N�t�\��q�E�#�m���Y����ʽ�;� �B�/�s8����%���Ջ�����1��N����W|N͡�'���MGp/IX��Ef��;��2�8+P;�A�J$��vuļƤ^c�&t��le�еyR����0���6�:�!�I'p���pV8N$Ne�6`P'[
�����aK��7w�n��(P��bh�@W2��w�	�h�$��6v�f�$�u�E���z�9b�V��v�ڹ7j3�;T8�)U��ͬ!Z�W�M���,ьu��\7)e��N�k�x�
��9����t�����\Wl�S�I'�K
��b�Δ/7{�s�0��s��ڎ��[vë��]��]���Sm��7�WR�R�*L5�js�*��ՄZ�V֓����-��u�=i�ӈ�Z��ꅫq�K�4$f.l�8ƌ �͹k3y����㽰-�IH��ٝ�t�6�8�f˕@;_e�N�=w�ȀKՍb��"��oo���z�wv_^�=�wg2��m�k#�Τ��v!�>���嵦�!F�љ������~��j� 6��Qmn&�
p�ѱY�gNRtLn�(�ͮ�ֵ��~�_���l�9��m��c�+����D�lٶ�rf�����9^^�D�e)e�ͻN9�9�V'ht'I˳�׶��r͔fXm{��^tm�)#���XݲӋ�פqm���xm�1�(��X�1�gY-�m��fX���`����;e��sVu�vz5��YbM�ٝ���Kn�n[�8�܉�[Y;�$A&Zm��M�tZQ�:�l��98�q������#����<�n6��l��e�쬰���&bpvimdƶ[m3Dw���n�۸�;[7lȽ����5����8�_�����������:Arb���c���'�SYY%�W��	;�n�z�LP�PL�oG�S�K���3�[����BZu��38��+�!RX
��o2{Nܽ��l6#������4l��g��/�CV���m��AegM�	Q��=鯸n139�/_�����6'�����Vw��K~�Kz�|�g�}n���}X��\H$�n&�_D��Q��{!fsߍ��\0��:ۼ	����3��:�}�<�������q�y�a�w��펾;���X��N��H/E���[�[�ql���\GBw�v�G�׵z�$����］Kܪ�4
�0�9��7�8:�'��hI�S7G���)��ZO*���'��){�HW���|��|����H�c�V��<B�i�;��<g�(�G�߉{O��/�AO��r����\o�kqMf�*I����#���H:��ZϺ�Z��_{ڄ�����{~Ѧjq��v��S\�5����G^���f�8� �S8g35
G��ظ8��\�&���"�&^k�#�#l}`��v�������0��s#y6�����v^�̇34����BV7p��lhS+v%k͉L��j\�wvF��o,�=F*p.���;���YOU7�g�qD�wq�޸��>��;����yD�����ZZ,z���Y8d��H_�����˳q#B����w�O���I}�i�J�V���<Fm�x�<���g���e]R��{_h��n13���f�g����!cL�����p���]K�b�z����O�#ZC��mlW�@�M��AQ}��q�BWi��0���6�%~��w�XY[u�_�oڥ/qDwwg�c:����^�io�[oLڰ*!�Q�۳�|yx�ni��BKC>#���l�	��/9�M�ʜ�د�$��T��Rs7RGd�qv��v�͈�,'�C8�ݜF=�g���b��x��Lӏi'�eyaX&��-�>�T��9���׾��ߝu.�N䖜�9���P���-�X{�`�	��j6��6�jQ_�y?m]-������{;�1���֮�T��D^�'d9$�J��K��<�E��so���0�l���]6�b�J)+�n�[��J�eM����F0�+����Y:���,�.�����7Ѯ4W*���}��]c�dD粽����A"�m��.xܽ�×>ϒ'�i_�`6B�b�Ru�=�Z�$�u�x8l_T���v����.m`�o؍o���qգ蘤��F�4ډ�dL9}�Z9�A0mk(�C�Anc]}}��
�-Iyq[�/;�cA����
M{x��d������m oу�6#��ń����7&Ƙ�S�xk|��SK$ߦm�B�FW��[ݞTg�|���l-J�KP�\g��k&�EL���a��ߩ+�H�n���^ݼ�����e��7ڹ�x�Xl�^�]���}pR���;����h��%->YB��|(�_W�x���}���gl.�3�0#;j�n�ߊ�� �����Ko���xKc��|̀e�c�5���{�^�U�Mr��'�$S�La~�-��٫�q��\Svv�;J�6�1ջWX"~ž���N,��݉�R���/�^� �S�*��ǹ�87fj����d�7��7)k5^`�׽�j���u�7��qR���a\���7D��ׄ?��aj��&u�hTﳎ\�oo�pv=�'��u%9妥��b��4�g{Ô�1R-n&3k����c�A�H��)����Z}��5��ҏMv��qgMg���מ��=3j�~=`����Xa�C�/�z�k�WgMe�R7����i3�5���'=4�2�S����85�\d�y����|��
���u�8y�g�5/|��y-zqlJ&�ߡ�j���8j���gT���W���wl��žm���#8�G7J:��V��I�#��tFq�R���
��P�xw�<
���]�)R:�}�{˻2��`%���b:��b�j���~���Q�}�b2�x������>9EN�$������'�T�G�����O1އ=��'�5y�ur�a����X�l[a�&h�c���~�����`98�欏3���1��g��;��wq	��)`o�X-E���VJ������>���MX�[nB��%�1�*�9	��������gm�f�+��Y��.�r�է>n�/j�4��tc��<:���kgXU�^f;��M
�X�䨵v�j4.oP�-��݅��B��n�ݗ�o��<>u]�3d��̗���(�í*��*:��up��g>>���6,�
�Z�j�ȵ�cʻ<FlN������e�G�fB����h.�^�-�[���e�,?g�0�����F�3�nO`�b��>���/F�0��E�>�hX;���}y~��*kkx���<9��|�7nY� ���%�6$PN��E4�wTʤ��R���I���<$���)g�i,<Xo0Om|w%��A����³�çͣ�(:����6z��M�ˋ6l$Y�|�G�.+�.���*^%�v"�K� }�>�`�9�X�2�9�~3���Rj�}�R�yiw�o���=<�磪�g%W�l��>>wx_M�m�93��(�/eNwI���Iӻ���0'�������[�|��oo�}gk<�~g�Ύv.��8ç�Լ��������=�=��BB�d<fx�i��!`�ڢ�̺�t�ؾ�c`�؃���r��0>r���#,�ћ���|霾�f�J��x�L�'itVP��,r�*l|����v5�u��e�?\�����^��.���KN�J��0��H�-��V��^0،�Y�(J�����L����{|�f�z}�R�r>ϒ'2�@��Yb]��}Q��ı��T	)oTt:���q�^�f��=a�>}ay��[m���Z���AST��������ۙ��F "V,�h��A{J<(�AVWU���Hb��\V�����f_e� ��Bi���5��O��O����?�2����<K=&���.}� ��68@��U9�py������m_~��p�^���¸�O��{�{!���T47Cջ��fqQu��kp�?M�b�ۭL��Gp�����1m�v��xX��~�Dng�I'i�F����<��E�\�{�����5k:�o���ڏ]p��!�"��B�_X�M����6�%~��l��,/M�l�m�f��V�Zc�`������Ze��ͯ}1Z�1�1������B��F��RjgG�B�ͳ�A���3u-�7�[@�U1Mh�qq��۵:��;(;��Ǫ�Iop޸gN��9���,�ض¾z��t������x�W�j31�ިw5Qf1����W6�k�瑛�93@ި�C=�2�`���N��t�ݫk}+ND�ײ�����3}h���m�u�MUе�����l�߉��0��0����[	�d�<y�ϸ�j[	6p���
D=�3Z���3`=��$��]�P��G|��y��^�����o��'P����������u��u��:�9{�%*l��3���q�{�8���&=�9���O+g�NG�s�	�~����,"R�v�"�EI��v�w䃉��	[!n�C}�����c��N��T�z�vz�4�}|G���7D� 0�G�CVװ����{�ݬ�*иڿ��V��;�9zx�H�{����e�5RU4�`��nV��2F�k����s�C��i�k���e6,4��^]7&��3L]W�j��o��{��񪬳�nf�e�}c�16֭-B�"�hv? kf��Ndr�ϥ��Cb��S{��G��M�ώ�����Ab���g�.ut"��8}�ȧS�s�lsܘw�p`�S�0�	Zn�k�^�X��ɷ���������\S��ȕ�էg����x����#Ϋ|.�u�.���5����b=�a ��dþ�lj����C]�!��ǋ���{�v6�T�ڃ��,�oV����{�0��݀m;#>���z�x��?{�޿8�1x,�$9M�j^Kv,��e���С�Azײ)��Bϙ�8|��g�m߯Q<����=�j��箚9������g�
��-_�M��Qh>꿸��������z����z̈́�q�}��BR����U����������9)��e=cO~3j�k:P���G���'x ��|��b�[tR��:��}6	��~M&\����tu�Yq��<��X���b�ïU7�u�9��م5/|��]��>�rY��_�U�O�MC�Í	�\t����4u`��σie��l��dB�(��6i�{�r7��}��^��PZ��޾�Ǌ�d�j�lਏM��RƬ���������sǇ8LoS}kp�P��5^�y��*��/0HC���}fe��F��7���b,m�ܛV��v��(e��@�kzn�;,�&��E}K.�TS��QH[F�>=9�y�r����r�d�2����ÿGu�yD�Nk�j:=��T!��ۚ�'�Y��ol�t��[��.5~��&����^*O���8"~�	ϼ�ğU9��e���>���[k�w��n�/��͇_L����f
9ꌮY�f��g���gk�/��U�(��ZH��&��/��Bn4b�\j�rU��YX�z<ᖡٯ{�q!4���ƴ]�8}[|��X�^zr�����[�vO��n�3�=�A����'�Ж���S��z�����S��,�h
Ӌ�٨�bl{y��6��yC�M w��OeU�13�/��vfqĥ<�on�S7k۷�e�͉����*��;=狠�nz�k�)y��m`i,<M�f{NܾX+I>��6/g�hO��&.��}
��:>P'�q��,��e"��?����t|P����~��]�r��Vl��s�;�z��Z2N������MUy�hTA\�z��/K���Q�k��S߻��+�Ř�τL���<��SH��	��$���ǩ1r�ءU�Q������r���	\+8B2cP�}G۷�wi��e�t�X�av��A�}J��5�۬	c/G�O��bō���﯊��}���V�P�u,�҇.�g�0c�}��ʟL¡r��9��Ү9�|3��)�g�_)�=��Ǻ�hK*��X�܌�}Ն+V.^<��r�O%���c�`���=��B8ȑ��_��p\��آ=�t�׻�:]���R�ϰ$Ne"l#����@������������cك�/5�"Uq��]��l2̯�͈s]�hH��Ni0�QܟD8PaĽt;��n �����9_&��C��y6��NY	�n�59�]�k���{�]d����!��$17k#o�ܳ��ۈƛrQ@s��5�����UcVO��Uퟻ������`���'ہ�����W�_˄�{jǖ�R��d���_/��������.�-('p*+Oz"�+���~�������i����r�wU)��T�]�JwWT���)�uR��T��uH�uw�]ԗZ��U���_JN��I.�N�몑;�wUV�wU)�UJ]UJ]��ȕUJ]UJwwww�W'I�Juʰ&"������*���*�����*��@�A�   @U`EUT뻻�ꪔ�����������R���R����)}�u�u��U�U�U�W����R���R���R��AUij�TU`EU`AU`DU`AU`EU`AU`AUa.�N붫w\��w)u�@���0����(" ����'ǻ����:���l~�Ɨ��~?aC�އ��rT�)C��}�Oǿ^'I� EErx������z�Q_�� �F����:=�� EE~�3�����A���{�/�W��<<_�Q� 
�+'+��λ���t���N���J��ܺ�ӻ�`�UX0UX�U�@ �U�AU`AUaU�U�  �EV �EYE@�D ���b��%���P;��=���AY R@�Dd��I����ϗ[d0>�����*+��Q�Oy��n�~�'p�Xa�Ac�����k�n�@DTW�TW�{c��� "��H�j���`�����q�
;Q�����c��H�٨�l ���C�;��;;@Q[8��w�&�GN���Ξ��X�p EE{�OH*+��Ր;G��
�(�#���el:܎}���*+p�I���{Q�(�\�Σ���� ������j�����'��<u]��������)���LW �[,�8(���1#��x��!�fJ�!(�i�j�kl��EATJ6�l�EI�[,$"��J�Z�CQ�ք6�@Q
�MKmi�64�b%��mT�on�U4a6mTЬ�b�eV��m�F�l5U�Ll5��(ֶm�2`�f�Q�SR�4�F�ж*�[6�ڴ�(հR�,ZcNwvfųKJɩ�,l[22Z�m�[V��,kUV�љm���6eiX-5�2�2���b��U�5kla[eD�kZk&��)�k(e2��]eN̨�e�/   ����u�={z�:�rٻr���{v��[oU����=�����ݮץ��u������zx
v���wo\��n���4z!���]=��u�ۮ��޺���w�;�v�]��Y疬�kmkfIC-��ck�   ���D�T�D����H�"�T�2O}|ۼB�J����BGZ]����P��iR�T���仫��ն��oi�������]m��{�ڵ^�t�y�O^ڻ��մ�S��{w��ޖ7)��Z�V��^�2ʹ�̳Q������L_   �}ݻ�.�_sw�����n��U��u7]{O^��]ޏ�v뛫׽u�3������Wv�ރ׽ʩw�޶��Z;ַ���׺{�m���Y�=��<�Խ{�G�owu�kn���ö���fR��"��UZ¾   �^��{��i�ƞ�J��޵C��r��=�wv�,����;{{[Z����uv��v��S���=�3�[���km^����ǵz���ޘ���u�{�۷�m��.�<�M�m�Z�dֶm[0E��g�  �z:>����*�w�=���^a��U��ڷ,ݺ�t�[�f��77�n �n���.��:�*�i&ݝ�������Z���5`�j�m+Sj�  n�F��n��}���C�M=p��@T���w:^ޝ�a�n�Nޱ�Cv�����m�4w��ښ��p�a@v��YW�z�J��Ҷ�ka3d���Mi�|  �Ƶ@}_p7u�і�Ԙ������{��TW�^��`W�]�ns�&��PΆ�]�w��^�m]^�[j��Ҁ����СozfٶkMa����Q�-!|  o>�� ���AJ g�å: 3:���5�)� ��� �� S��ٜꇢ�N��x����^��{�B���6-���ci�ZY%��   �����@t.��@���^��@˞�z�S�.x{�CTwE��^�7��=
��a@��^���������Ҁz�7�l)�L���#KK4���   }�{���A缮� Qq�u( w�p@w�� :���z:5@�k�ХP�6�� �:�� zn� uJ�|�{@�)T�HF�Oh���F�di�M���%*)�  O�JU5 h��T�S��  $�T&R ��G�����:�����ww�?��������Z'D#�먻^�VB*�7
�x{�x{޽��}����cm�`1�������o��6��ll� 6��������^<��4��J!��.��R��@MD�Y�D�K�tpʵv��t�"���t+�n��nTS*91JJX	�����f�����-c	U����m��.�WL㳌�ΧW.X����&�"��[l�*�F��Ԗ�"U���Ti��4�����n��b�RKY'�Т��1d���6%��.�3]ҡ��DٽA� �bv&����F��x�U���\a*���y��$u�rP�6K":E�mE���.���FITj2oS�A�e��ǆeaP�sv�a�2�M�Ob6���F�d���|Q�����x1�wv�J��.%��7ը��w�Y9�En������a}��!���cfQ��Xwb�d�t��ɋ*�͒�kن��+�n�KcN�b�K�egqMx���ǝ������&�$m�����4��6�)Yt3-# �r�4��YA`g�jU�W�
��M�t۹tR�*��X�M�]��1����n���DK�e�P�2�e����j�I ��"��܏)œV팩l��TՈN)A����(c�l!�"�ax���"Չ��)мy��t���q+&��6Z��e��)�&��k"��x�r��]!/��J�-1��op2��F)p�w�ұ�3@�C
.�X2�TVW7$1O/5�n�4B��ݛs>[h��x���ʂ3N�4V�r�]���C�Z�=�BDp��ok9z�Eв�Y	�1"�n��=Fd�0"���Q�ƨ�r��VL�a�eH��uS��j%f0��X0�^�f��i��3[�v�n�ҍ`[k$E��&�J���;�o#YHfXJeJ15pi���4U�4o���#)K%�cʽÒ�S:O��֌*)*C	Ph�0��heU�[�I3a�n"-@�,n����RwV�ջgqݤ���ҩ�\�Vmҝ��ek"�x��,��.��صn[OCHx$�P
l��T^T74�V۔�+4ST�)�Gl��Du�{�[��&�1.��v{{�W-G��u��%B�!�n���4͡	��`9Yo^�9DY ,�i���C7"���]ou�ڰ��X*�he7t~O/�w-�Xv���ܟ�)�4� .�m��I:h!�]G0�x�ʬw%�v&GM���,��UaWn47�^��2�:1�&5��3qf9�6���؁�i�.%M��5r���U&�?��`x�n�4�gk�GU5�mx(����*�A!{7�/2��	d�!	��Y�D�G^�?l7^J1��޵pK#�%�FfVU�
�m蕜#�Q��r�9�����p]�iNR�H+f�%����흵Z���,�3�[�7���&���n7��)��?m�BXĩn��C�J�6ъM��(47�Ӽ��q�&�7`U��jԭ�lY�ؔ�U���M:R#y51H:��<�&�ѥ]AB��"�c�U�ZE�"�F�QX�פb��|�k��;�N*�D^�xP�)Rl�R�֖�u蹊�wB�)-Ԇ�d�K����-��Gf֌���a|	%��'
R��[���b�-�¯�X;�;H"�-J�,7�iӦd�X���OUxpXU��g/m�ڬ�aJV��I��r%{���{���SP�+j��C,z����#��u�=�R�Aw�7L��!{sJ�!�M$1��������k/K�.��a$L"n�b-�)bZ
:M;�3U�[���RZ�=lZ�Qf�u�T��6���h.��چ���v�WR�HjT���]���#/s6�E�Mܼ�ɂa�@�77h�;R&�� R�&�LCG,��h�2r�7��!j^�iV��p��{��@�an��Ű��2j��5���sv�X��1ˆ�9�
��Q���$\j�؉AP4�ρ���`�½�/ݚ��C鷲-ɹFe���̈[_C�q�_�3�#5�n���f� �*b[(���[� 8d{�>+R�[�63;s�o5�%䵋w.1�XdU��50�X��Α�����n�;�� bGe�-�%a��m惂� ��h3fD�X.��P��ʛz� �MT�k�(R�#������)E�֍B�{��u���虲MS-�9e���QʫPY��e�e�c��vd��,�ۏ-8�Y*�Z��^ŔmZ�@:�
��%V.*�4:4�v(:n�^�W$� ��NX4���-�KD�Z�������%��۴o��OA[�smEG0ŀyb�
c��N�$�p;���u1C����m��yY��"���9�Z�>�X��E발UJjΡ�Z�E
&H�����H���E�B	+��clb�`�qX�r#{�N-��g�$�B�5/,���%�&n�0�VaW��0|�q,wwJ�V�);�o�i9�dٖ�RHTĀ�6nn�l[�˩[x������8:Uu��4 wCl�w���x[h�l����j1�-]\@�*��S>�z+#ckY�2���eղ��&'Hؘ�݈Sr�_���Qh���R�#W ��Q�R�o�4ޱ�cR�Ś��8� ���1c�uuq�Zs*3��2���Z�u�,Ƙ��3!����	;2�Qh7Q=�6b�h����&b��*��a�X�jjIw�p�q	���M	D�-
C���4�wN��.��ԧ.����XS�J�p�6�sd	�Vѭ%Ua3L十���%Rt�ȹ��[���v*<�Z�xJ�d�)[[�-�E`%R��nh#6��k%1pe&�:�o�B2�ۖ��A4j�7�@��%�W1�)��VJ�H][G&V��6/Q�$�Z0}�&���R�R�E�e2�:��l��N9#۩l�dd�\��QϯJj>;�-���v�`�`V���te��9v4������4�
��ӹ)�yJ�nBͭ�gmk�v �S�X[Ղ�87&�q]�6��tX�Z��	q�4����RMؒ�n����Z�Re�G2�v7M��M�wtŦsy��C�\�]HW찫31:6����V�m2����a���Q�֝)2��I��	mCr7Lm����\x�t������]H���K5(�(N&���)�4@ŨH�Q(��L��\��"HM���xT��/d1E�N��1�%͔��F��yGUk�)\[��{�lL
V��g��4�+�\�R��a�bz����t�����'/sp�궵���3cJ舄xB�CA�����x���J��u�mJV��ʆŜ�QO�5^��Y�9@��;3[��ٹ�ش�]XǄ�"{2���PU�J��S4-�g�WUq�N��N�m7h�\�
YN����وj��Ӕ�
��iMj1�ͣ*��w-�gڗy���Ue=Ņ�	���+��I�[�lf� ��7�1Y��Oe��o�]��7`0 -�=�U���l-�z���DRo\J�:�+�j��[Žww,���B���w:'�炵!�.٢Ffs)�x�E؈ږ������f�����f���4��͆óY�M@Em�
�h�MU��t��9[	�0Z˵/
[��(��r��J���E�U������FP܃Dَ}�o�7�S[C��[LOJ]E֌|��J8_4$a"�$b4`�d%�َ�]Z:�Y�]�4)�R��q�V��Z�H��]7�ɵ�ϛ#<)���}D_�\�>�"��[���ڵ�Ohk��!j�M�V�L��a�㥘���,��,��y���l��C5C�6] ��4b��rR���t��oDreh��m��*]f��kp2wt\��=�f	u��2���V�4�,V���#C��~6=�wY7h�N��qE���dZ@%Q�%��#ؐnM��-k��s��q�u T�a]�����m=���5=��Y)j���I���m��l���kB��zMK)���v Y Y,���.���s\kBu:	�lm�ea�&d��6ٖv7@n���;&/q0�i|�B1�o�J4�T+d-�@�0կ�?i!t57�nʹ��Yi0��K4Bxކ���GS��駴���6�
e�5e2�w1]% Su��e�2�N'�w�$飱7���ǌ��4�A�Z�=���u�ˡ��L՗&��Uf��#�'��D%�*�^V�H��6]�Ђ�ǴPG3�m<�ݧ-1X���e�M�suۗ��f�K�"m(�5�s60\"�ǈ���K�6H�(P�u*��eACQ�P���x��j�!�mQu�-����͕k$2˫�UlJ�c8D�2[�qˉHHSS��uxCm�!3���Y��c2�b�=̹AJ�� 76j�+�˔�-F�\����"�Z.�u�)�B��yOa�� ��`�N�Cbn�7�i�@äZ�K�Q�X�ģa����o�}uG�Ӻx��l�[�C1$�bn�f�����l�G㭡��TX�0bz�f�	Uu�j���	���Ɵ�hLZ�:p�Y/T*�S�6)��2)��.ܹd�孑n&��t�*8�[��Y+v��e�f,+Pb��&�Kxv!�k��;Sq��刚�I����g�_'��)4�t|CU.�Ȉ�♔�m�	�F�iC.�h��(ӭ���-�;��X��ӫۦں����vLd�9{"����yf�0a���L��X�N�GxXy�U��M�0�R��K;�1Ǳ��	 \�e�*P-�b}��W
�R?�s8\N�9ef���xfR&�����y�lF�j�*i�M� �/i�����47�!xb,�6M��*�F�n�^�Yz�r�6j�gV�I8�N�DS5(=5/K6��+*m�sTe�
e��V轭5��2D�������ROE�V#ĲQ{�r����i����s�!G�y@�#��-�H �9o̧��r=��Q�=���r����.Yĥ*���sv`av�H�+c��B`B���[X7;J��%Ǩ�ո���f��ceУ�q�*`�L��7�ӆ��dfʠC�񼩘�˻OGv�"�cF	qf!C%��6,t��V�I��)Â�Gl��	�mn�K�77A�ĥ����)t��{����R��#L�XG�DS��bo45/��jёR����!rf@t�~i[���=
Ę.��ʂc:�\������mc�H�Q)�/F�x|pY	e%d���
1\�53!TS��`c�u/\�/%]�ܒ���9gd�\�c��G��n�A���V\����+u���}�KçSˢn��F��^F�ǨͲ���svBu[z��k[�jT`ReVTр�"��坷��;�b�2�hQ�u�U��T�b�W%JK:�����5��nධ����b%�e���w�Q9,Tx���i��
Vޒ��J�kQ�e\�,�y���a��Q�)��sїf݀7@�2�y��8$0Y�������;����X�%���������W�U�T��n�z�]�b�TA����{�d�mc'Yt%b{.a�M8M�;C�o���p��w1���Q�
���,v4�&� B{X�:�Q��Z���(\R�U��l\Y2��k��4��+RJ�n�Y��#w  �ʶ��[Yu$�5����b��K��ȋע,c&���"l�d2��vEii%T��mnj��tFfV�ա�O*�Ѥ�	.���MQ�q͉m��%�K7�6��RiƄ��^���yZ�z�2��̽�xq���WV6�cɉk�[{6;�$3v\f�53N��NH6F�����f˚"2��H����ĩfF�o�$r�y���Ƥ	ɔ��2T,d��$����4�P�GlĚ��:7`F��6�黟@
����Pǖ�X��ژ�;[7lcYMH/�rKr|1i�)n��d�K�H��ph��Z�Դ�`���YD�c[����e	c.��D��P�������f�TmBN;�ݻ��6���g��#�##���˭hM�Z�
�nZ4%i;X2h��cp02Iopk�\�`"9�9O(ˉAY���.o^
or�[�C,%Sw"�%���e�"f���Y�.�=J�e�7�~=M�5�*mG�)N<a�f�T���%�t�T�Ձ6��۔%kKk&͵o+%�2�U�j���n�iD�,ɴ�e�`�{���H��� U�X����;M����M�-��"�2^	2Р�w�6���&��JKĂ�,8��T��-e(s&�wf�!�E���Ā���̲.��f��ϡB*/e?�����y�ֻeu� ]����f�VǓV���:Ħ���y�6`:��#A���:kmѢ����ٳ,���M�*#bUާn�P�f:��T��R�x�v
iI��������#��,FE����ӈ���EP<����q�GE����"�� vj�ջ���m`(L�b�T���1ͽ;rc��ĞVF5ղ��K3Xcwcv$`�x�C��P�fhM��T�^H��`��f�CvV�M żd`1��ڙW@��Hy5����W4\Fݔ���^��&����V�m�[q4��b��K8�mY�ia��.F ��WB�z�]}Y4K��4��A�J�Y陪<�D���Ik��]��q-�B�c��F�~�.�KC6�'4��2M�&ɐiט�t�AW����Ú�5D�@�)g�a�Ř^�Z�i�,�����\�̕���Tʏ��L.��n��w�Ecv:fIJb���/^��L:Ʊ�&�� � 1����K)[��U�ܓX7�64�L�����#X�i0�TeF��jJ髖/"�ښ>8���+:�KE�����~��N 5N���P�J6����Jl�e[/zm�,rq�kR`��0\cl-�:k)�%�w\�X�����mM�m���a��i0�.G{r���\I�ީO��A<�G;y9�����"u_U�o9W8r�ǻ˙�#-���F�1\T.<&�WwN�4C6�K @����{}Ž/���(��%:�g�.��e>���Ywj�vor��E�1>d����ʙZ�3;;aKn�K�G�֮��a�g�k`9}��j�vw\�(7��es��Ֆ�����k2L��y�ި�`�%N8��3��-�.ږ�3�ps�K s�2{hQ��^�g^F#%.���_V+��3�R4����
'p�d�B�jg?����)9�R��9q�%��Z�=�u�{t�vJ�1�P�ɸظ��J�ˁ����N���೒��N�c�D�פ+	�o[
Z��!ǧ\��)F�7���<|�9�J�����ѭe���u�	xc�E:�C5-�[#=Z�u�7�r�L9���#S%oY�[��kU=�$ǶzWdڤ7L����4�H%��sv�*F�X�Z����S�"8�b���Jmu�A�E�:�N�o�q,W]�t��b -L�� �w9>��Rv��2'�p\4^ı*`���"�Ab�����1e*���n�!�4;Ȁʭ���t�Y��MV񤻮��:��)p�Gk"/I7��5-�;|�ld�C�`N�մ9j=O��b˳y;��F����C7dLN]���]CV���}�]�GfN6��W|�Z��0>t����9���o':��u�q�p�������)�+����p#X�)Wt����@�s�;�[/R�:}\
Z8L��ε�:h�!d}p7�Y����K��UiQ(��ܲS�N�m]aU�-����;Y���٢���p����
m��C6���S���Q�3�3@j�ͨ�k�V$:���*��BWt/j:T�J/!��+@��Rӵk"s�u�����B�K
�FKǎ�Ԃ�����S�cjH�
�9r�|�o8Y6@卖�afL��iq15��ԮF�o2w�n��+U5$s&��,n'�M���B�y��Z��*��y��v\{��Y� #���ܗ�f��'ZX�oηR������L�ʸ޵��ê��c�k�V�c�H�Ǘ-͑�9+�Y��iƧL��t�8w%�w��2v�P���`}y���.b��.�<����t#B��WV4_"�M�=Y6Vf]�5en�(��0E���P���,�밹��+(bF)NcU�ee�u�H�����{E�ooi/�尩�����Ў��a̐����R���g,��
ѹZ�=�U�$��<W�G:��!�d	���:s7��D�t9h�6Y�7�S;��Ø��i;�*^dN�K���Էūa�Жe�e�}y�V���M������y,��ֹ� �.T��z��X{�5��-�X�V�C�`s��3d�W�鵜�2eۣx� �����-�T4�<Vqj`V'yw�>�)�\��N�Q��.`���
�,�s�(Z��n��2D|��*�J�F�	��:���ױ0r"p��uV�!�)�b�slPY�^�j��2�\�L��Ź^��ˊ�&Y:��m	�fTK�v�S��k��I�R�;�@ZyT�uw�Zb��h��b��SW�	��;,]�h]�Bu��ժ�U'M#�X|�֧�9���qضX��{�8�ֹ�"�NU����	 �83]/��Y����u�]dv�*m@�v��3I��]�� Hs��85���
Ů��SԶG|���T��e����)�u�G!�w)اx���CP&�Ư�n����=GW8ݞn�D�r�9:e��!@��VG�����ԭ��Oyť�[Y�D�+1�`*�x͛	�8�]:s ��#b��8gf����7%/�>�	o1Ft��(��x�l���9���V�iǇyM�ܝC�n�>��Z�K��v��gۑz�i��������X��`MwW;�	�^nYX�D�L��P�s,����j�2i�S�|]vV:%���J��jN{��u��[�@�����y�,ʲ!`��ي��	��5�U�)�j
6�P�^����N�iL�5T�/�r�s�*�B@�Pv9X3w���4�� �&�sTĮ�b�x��A#�.�u*�w2¦@÷k�p,_Z�/H��ζ�-ӝ4��x%s���An#S��wj\e8�Ku8�7eef�]KD©���5��d�z-���ܞvr��1Ç8L�M�j�P��{t�lIzKz�7�O��<S��0�c�7hq��bv��j�Vt��,�-V1ۋE�+��nXW�ê�x�g2�0ų8!lm"ܮ��Ʀb�lQ��l-\hƹ} �2���(�5(�W,�^��{#��V,��]~	�2�H��/�Qieq���f�Vf4��Ol1+M�N�R�R��q��֯��m���t�j���.ʽ����L�n�� �v񣳗TW�uv5uʰ7V���n�V�Udt�"�l�Ku�D�����3������>��C8���ƹ�#u�0�2}O�a�ڜ��0�&�g���GD8mt�7<NG�
���@6@��{լw-6"R.�MƴWv*/a�.ܲl�L���༁^���j$֞`P���,�f+zsf���V��љ:�f]�R��.���z��"���L&���Ϯ��P���n86����N��2��N'��ԭdLoyr�\�^�+	t-����(��V�x{YS��9��Kw����f�:˭�T�i�ZBgj��X�nfq����@��q�����	�&�X�vc)�4�e0�ȩ�*����jȭ�E\MB�,�<��Xx�(k�7��5+��Y@RW�fh�G�lB���&��,����k?"�q�#W��9@�e���xW^
��Ŷ�\38T��H�y3���Mz�S�oM,Mv.�����N@����,�Q!u�r�Z��U�����S�	�$�\�n��T��_JB��YQ�oV��mN�`��ʛ`����IS�$ʾK;'�:;��%���:*�l�M�Iy��r�UV�3�qQ�Ũ���.�wV�ެ���-�3`ik,NBn����5�1w+\����u-W74D��Se�o��&�K/24�P�[j�,X�Wƞ��C����%��/��L;ҎEַ*ɬE�r��i%j����Si��S���]8��R/&K N�i�}�؄3&Ыs�v��W�1��`/j��҉�	����*}���qD%.�Z�m��,\�Wt���W#ʢ2gHm�9]�V�.�pU�Oq+W�E�ɣ�3���Lv!�FTYGKX*��Ʀ��� ~�f�*��3��w�Z~T�hX���DJ�q�����X1�a����i�-�\b|m)�t$3*�Cf�O:���O
*L��+��%��p���vn�mͲy��l\��nº;��Nq�a��t@=��B�5���X/���tvG\/Ȁ�3�S_^Q-����Zs7lN�.v�� �A��\����'e!w)=�n ����[�t�����
��W;ǲ�֡0/�C2>�F�U,��,�.YQ9{7:f��J͝�Z�N ��T�ւ��iu�B��#WY������E�J��˭�QJ�t���u����D��F�m�g,�V����,*or���59��Z�G�+6,���F�ݠ��(��k�����x�hAq��{��4����k,�o.緔�q�ztEOcW���q��<7F�I�oWM�Cm�7���;��gV6v�����ԪN���A�m<�:y�c�.K@GlTH�{&v�\�;��C'���X�*�+1�Z�Rj3�Q}u�Xʍ�Ok���\nm����Z9BJ���Ր��2�Iz�=�����}Z�}��҂�NN^iZ�B/�b_��f�E�X�9�}[+i�j<u�����-){�hU��c��f��x\=x��Z����)��R�֮(i�YxD�l$����1�%km�2$��܉��A�:A��%���|2�ґuJ�y��Ǩ������w��8Zk:0֍�-*���V�n:��������M8�:�5Xk�sr�<��
k�a�@uIkv���1N��}�H	Dk�����
}*Q=�o�{w�#�m����Mf\�)#��at���"��.���;��)ub��Fd�� }��<r�+2����Ҟ :HdK��`��z"����s+���_ ��$P��R�vΕ{{4r�.����ۊ�)a�Y��v�������bOq�W~�3��lC(��vf���&m	�n�xC�S�9K�c���QB��v�+�\�F/��1X����{�f�[���@z�vO*���g��r��Ȧ�*ӽ�r�wm�nd���X�ɝ�K��G|Zq�K+kv�wLɰIՅ��m)y����`�ۈC�,W;e��T��<V��j�L3�q���]���:ū��f1GÓG���� �V�Og=�ˎ�U��q=/c��%.�,�(	i��G�U�ܮ���/xP�J�z�F'jq=\��9�^iL�i�H�ah20)�f������p��Ay�IH�b����h�@,/OWq��li��ظ�u��.�M��_r�ݎ�'%��ZN;P�`��[SU�2��S�˝�M��};Ȳ�����B�)�Ғy�5N�h��w�DŨWv�Z�#���+�C�OHQ�&LT���DU�k��ݙ"o�(fZ(�3�M��5�N���
WՍ�� `g9��z�^m	�(�Hfd@LI�JX:�'�=ǈ���ټ�#!;�IK�:���R��M��+��%��ܮޗ�p.��f��&K�I�u��
���5�2��ld=������3I+Ѣ����c��22����	�M�GH�
�*oQ�c'��$�K���2��\k�YSd��.����wZ��76���iFz���)neA�7]�K���]qb1�
ܡ�{eC��Q�DƝ#B����,<�:�\�[���C�<�y�]�vDr��g����Mr16]��>����Y�o1t���b"��׏2�ę�|�m����c�Q5���+��Qh�j:��S�y�
�Z�_R7��!G�N>���є=xo�[���A�4d)���rÔ
�ų�K*!�0�KO}��bZ�DO�ܭ��=�&��M�)�}[-	sNB76����(��f�hS,P�{1��U#m�a�r��àv㔺�c����S�9r��:�K�#���<t�����\/�Gz��b0┟1o;Y������Т,m4�c�}C��g\[�Kͦ��cm>�Os;�oh]bd�S�W(Tu.�˒e�v��}�M$�޵X2v+��@׹fT��!��CH����(�~2�0�"����%K9�B[o,�):q����n�RZM���vݶ0V�y�`�`Y[���$��_V'���:OU�P�K��Z�C}B���
���[&g'�RY�����)�D�:�p�I80�KV\�+��ӋuⰌZ��c� gf�a�� �c���fI�nث�!k:�����v����aI�*GOME3�m�m����*��Z¹]o�@w�q��]�j�"&��I��L�W3��®�&3�⥼N��nŖ���qaV�Y�JC��;�!ChXd�eur�����]�7i<��[� �,��k�HL�̷kp̜���i72�f�jٶs��X��JL�1�G/��.�kd�Ā�Y�X�g �����ir�R�����Gvm���⬤!*�`�1w^�j���,��vw����"��K)��&[��܅l;��Ʈ�]����nw0u)��d���ҥqV�H�m�W��s��::wEp���$�}x*:#hE��ۄS��Z��}�է�Дβޒ��:�Y�
�Vf��w�k��	۷WK�k25.� �'�r�\�0Q���!���<��|³��
JM��әA��s�`�	�KblE)��B�b�f�UH���S�G;�J��EGV��e���y�ýN7�m�Z��S�r$y�Ơ�Y-h�ԛɰ*�G��Ų��$g3[k嘗]�ٯ�5y�)�]�w�E�V靀
ҧ��D>·�ʽ�	3)�rY�Z�vAL\������ֲ���	�o2�(�2�/���,�r#�F�BB���knH��3�r��0QK.f�=i)�V�-���[/9e�nH˔e]]�nn�b
�gf��ITR��z�uV9Y;�0��p�w�2�e�W��O7��T�ԏ����f�b7�̳�[ǽ �Up�]��/�F������u�1�s������L�ן3����Z�vK��}|�<t�~u��2��49S\�H�J!�\ݮI]fX�W`��.�R:b���;� p��+��I�Z���iw*$fe�i�b�3�S�͹gi���wK�vEç�4"P��"�7�1N�]����5��ec�fk2�{��#Gr����_}4�J��K�I��3�mN�=��j*��9[m!��W�J�4w[}3a��i8��Y��X[:�gk�.�[4wYMҐ1],��Q�(p���"�;�f#��;gqHQ�Vr[0;�0�3cN�du���!���v_-�s�dA��Qj���f3��ਊY�d:�7�6��g��2�j����E1�p1�,��!}vF�����\�E|MvM8sz9{��	$���Jh���7�m�����DcF.V�<�����g7[��JT�;�=ph���@Ҷ5��T��
�w-���&B�Z���!��Cv5b��( Ӵ�}�������Y�t��'WF��f���%t�w���#��tD�[ ���y�Y�RK�✮��c@��,V%"�(���T���� {��� ��xxx�������2�6~L�®�fed�?RYȧ`�W���p�Z�io%H޶;�!&ŋ;,�fSvi}1�N_;Qh����{�bbp�]�p�/]����:� �2�M0�v;��9a�]7S�H���O�uʲ>�թ��[Q-���K��/���]uvM&��5�22AC�]
U�h;l5P�6ۢV����:XGPеm�T�F�e���d� ��9��73�Vg+C���\#3�Z3y�ZuM�kMG"�������&j6�\*n*"n���K	]���9Z����^b۬�V�4���u�����g�&3N���o���&��Rۀ@���ɭjG6s�3��\m4ɐȥ��w�v&�EDe(�Ec��]�xV�Qi�XI]T��
B5S�I9J�*���Sw&T+id㜢k�߆sܼk�����d1-]M|������kC���ޘ��U�v�n�]�kk�{) �h�����YEP�dW��Nk���{<�0f�Ň�Wt�\��8�M5�mC��{���IA�+�9�6��NuG-�^Q��5]�� GXir���vqJN�س��㸰���(Mըf8���iL`�Oot���Z����zb��"���#z	"l��^�+��

͸u�\����-'L0k+��G[�(ps��{o��;�����4���P�F�Q:�R�>U,S}�C�J��q?��*U���e�t�%r��m-������'"�U8�m�в�廵Ֆ�\���NEs�Ծ`�v�%n�H^�OnU���ٻ�(땮5�H�	��C��LJr���٘���C&�P�@��{w��뛁U����]� �n��YY�E^s�]��D�z,e5��s��t��awY{UgX�n��;�!�c��k���:]v_9����֕������s��T�l�U��}t�'������oVG\έsn�Sŷ4��%av�K;N���L����j)#8�/�Ԯ���8�O��&^�|�ZХԸ��4ѳ�$�s	�f��ӫ�/f��z�e�S�Vا2ȑKkkt\�WT�������Cw0�wcG�G�I��0�̊W�C�o[�R�=�w�COE]j���\�R�����v�yLwi2��?^����R����{�p5�!oFb@�F�+��:��D��fv�2���8��zN`2�����5�L�U�()P��J�(0-��e�_Mc�Z2���je�t�d*��t�ʺ���+3:�Q�]F�[]KRŎh���O Kԩ��IZ��{���U\n)��a�뛴̄+�o�+Q��w�qL���YA;�2��r���"�C�oo�@ݝ�] ���H�����+��R��} �dj�x�]\�P����Z����	�v�d�o5�t�y�8���Vet&S!t[*��f���9wF73
�c�[BX�]Fh�r��PR뗖� �j�B���vu��8�Uf5b�흙���5��ʳ��9\p�������	Zy��obw�٘��3����б���sc]�k��V���1�)v�
m\��\j� �q,ݝ�JT�+��0+5�e(:�1b��0L�Y��害AN5A(9���xX�8�"�܅1�k�7�(:M�L���B���g9u���ӥ��V����(Wq��ۙ���}2�BlSr��YPWS�7`� ��g����Ÿ9:�n�\t������u�K�M�GZ���b�%²rъ��R�Yf��b���1l�١J�K��I����'#����2|Vti\J	z5,��uHƓ��j�QC�"i��7Me]4D4V�-4hT��t�Ãz��p���gD;�V,3GQw�ӂ��`��;�y%���l������):Id	��kE��:wG{/p���t��Z�5T.���%I<��Ã������� ��b��*z�f�E�P��:�Q��ҝ5&�{�.�gb�wٜ71d�COf: `<�Y�5ї2�ԡ�K.�v�r@�jV�F��5���C�a3ӯ��\�qͬ���U1�L�BKV1u
�x����M�t�b�ѧ5շ(K��D�Oq��t���/k��ධ�����"a2;�-��j��1%*�P�G-;��^m�ː{;we5��iTq\E�<w��A��'
�H�*ɜD�r{9X���y5AJ�̝R�(s�*TZ-$��յ}���ˉ�mZ �ؒ�5ٺ'�I��o&�5]�C �Ǧ�����6���!��U�Ș�sR�մ��P ���WwQc��2ܖu��������R��4�<��tA��b�Ş��_Jz)�d�奜�	��G��X+�B�X�iv9Q�V��o�S��e���p�cvd��5���6��(_e�w�k�{{DB�n w)!��P�c�'f�~|��!�
�I�9r��^v�o7FWdx6�㹓R��/ga���h��̝�w�ZC)8X����[���uz]k'k��!�TI�)]Y����`;"B34�p�H������]#Pp��t�v�R�ƌ�U�.�0�bĚ�j�_o��o ұ��sU����h�[�5��w��@�f�y�!\vRV�4���FL=R��:`�h�a�Ծ�,_�wV�J��P�%t�\�v��Ɔu����ǵ��7��[:�&1yS9S`*�X�ڙ���d�����"�R+�=M�(dYmf�,ӱ�t�(P�ow'k+�Jb���<
�cx$��n��Bȕc^���3ds���",�=G�ܡ#�>�'9�����@=�	o9$�n�,tЍ\����WʞF�a�c�,��W{wE�)�3��Qc��NMul��jVi˜�=��4�R/��
��Q��ٮ�꿦��:���z�f���L����D"����Ͷ�XO`�Vd�PV	Y���1�D��Z�e]H��rVP�鿙[-�f*s*�t��f�S���(b��F�F&P��bϖ�X:#�	�R���V�<X�s�6nTW���2k'mʝNtY�:�;pr Bc����uu:�v�5�1���@�)H���Z�+�
7�r3kz�������h֡�c�'I��6iiyvl3�r��۫f��VP�b�B��V%�W���BL�gd���7r�8�c�R�����b��1*9#/Mc���>�~j��Vj�E�t����n$Y�Ƀ2�U�9k%n��>���tK�Ed����A�G���qs�h������J!S�k�˲p-�!��2��3@�3(�quJ[<KO1���G]����e���c���f���C(��S�X���#��n��ɘBV�A��-K�)6�v6�Z���Jъ�ɘ�:O�R�L�7Z�Λ�k
k�9�#��^��=t^iM�\7��A�];%r�r�-�"\�#��M@q])��ʖ��>�b�����1��%�ڸ�:��%f7��Lj<��9�̰2
aAis*�U���a��ڌR���+��<�޺���!Ӆ[����Yټ��N�Je�S���Q{v�����*�G��ܯ�-�����y���Āu�����l>�: �-��t���V2��5�|�W�X�S�F���W\ܣ�����.�
-T�9IR	�[{�ɷ|��>�"]��ˆ.bGF-�*o(u�Q�Wuz3��⧲��Kl�XG�Q������fR8��i��r����1Th���º�(�nQ���lV�j��.���Y�z�N�B�
�u�˩gN��]%��g���xq�5X'Z��v�[�2C�s��;��ri�ɲ��cF8ud���
�|I�]^���NZ�7��C�_T:�1��2uխ���/1B�n��Y5�2�4�ZO	��ZN<S>呬]�%��։�;����=�DN��7a6�]��4lԛ"WǷ㯙4��XwyDWm�_X�g@�0У�>6��N�z��4��q�&4����,<�+q`t, 3tC3���ɝ�qfv>U�ܔ��i_�����SN�w�'��s<��	=:/y�D+f�2^jr��](�K��{��_\:�}ΧI�T��r��j��޴!���z�|�ԃ}��wF���/��!̱����pɌ]�ڻO�8Ł%�jkfnh=1��C7�?	��d�ʒAYZ�P�3�C��:pu�n*���<-�iqP>�p@��}@� �F�s>���_EK�:�h�s�
��Y�u�7b�q�rl��Y�r���p7:�ѐ�����<Us3,��N��y4�����`�Z���V�t*���4�Յ�a���gJj�R�t'v��aB�+A^��s"�`�b�.�����3�r��3+�%�Wq�[|j�'e[�*K�5ɠAm���n�WsX�LP���LKU�m�Y������%�2��^����f����ξ3k���r���%�s R�F\,M!�������8j\feY�m�"���P���1�X_'��,�Rg^��+U+.�X0���%�	s����o)w%��>���XRud]J�5���K�ݙhgNk5�%�d�]ݚ�E���9�\�Ka����->�����&Вm��w����Y6�bu*p�r�y��9մ��"j.@�����p��L�)������������.�g#��Wn��J�)ѐ�tn"r�1u-�
�55�R��	�7|��V2s��dZO0m��\f�7�-�Wc��wSP �{:��t�4�ܺ����J�2l}xK�m2f�@<�R�˧v8_t,�%Sʍr��Y��ЮmC7:����J�xTh1HJ��jY�>f[�w��ա-oc�;�w���ku*�R���N���q��j�,r��KE���pB���s8�4�4���^���aq9�b�U�]=�O<p���1K���2)�Fs��Y����j�݃R;�*�Z�X91w9%ݳ����x(���8Ed%/���R���
�v�x�� ̽7l��7���1vU�)gZ��T�%n�Y�8Gn�H%��P6����mM̮��%�r#���' ,�lo*�M�:��QT�`7ï0�LSm��܆3n�Z���Z*XR.�-��s#����wt��4�)b�u�����SH[����' �+��	��'�e6��j�x[=Z�z�����W�:�Ľ����l���S�RI(���d(vʒq܂�_>?6�{�h��>��MǸ����e�w�m��1����U/�30%E�{�0�	h�d8�5�!����'/���̔#}>����	�$��4�ǵswX�:��m+�|H�hs��Ǫ�I���Δ2���3�!�g�Z5�g9ӡ��Ĕ���8�!Z摛�9��m].#0�ш��ΨV���C��v0�;�h�l�Qi-���>v;��3x� K� �a��O>S��HJ�uǰ=�bN}���t�i0�%�>��(5��b�M_e�|H�H���P��{�����Z6�pW�}i��
��|.�D����N����H�$�`q��vV9�4PyՐ�0����v���n����n$�!Q��f&����WWՀe�8� QV9���q�i�%!��Nʮ�ݭ���^�(;:��6��ܼ��Q�>ʄ��8�ĸܜ�R�b�]���Z��!�Q��+�.f<۩mqR�san�:�`���GKF�g��6��b0Wh���h
j�ZEcG��h8�n�$J���%�]�s���^�֮�����4��z�}]I�0~:�8��#
�|T��(��� �1;���]�vS\�Gl]��7h���GUq�+t��x�Z��_81�������Ln��F�,�����[�Lu:I^e�׹*��C��+�P��4z.�3yC�.�UȺ�a�.�y��@��u��˼�_'�W��yrO%�1IH�(8CA@����.���Q=�k�S��i�����n�I�@�NN���팲�V�,^pY�� ����(�p��B�� [;�Z	��-���^W25*�����f��)h6�C�'c�5����ҍҰzn"o���N�LC��_^*�J'>�W6w@�� ������M1G��[QKC`��]8#��[��f�I__VC>�E[X��n�+�لЖy�;���)X��]*��H����AX�1T߸�l�${W`YT*e"7 ��)n�f�"���;����f>��B �a&oN�TS;0����v^�`�vD��k��n` ^ �v��[r��iaFngD����n�k��������Q���7Ξ��k+>.P�Q�J�,���o�f4h���Хț1��9s2i�b�ꇛK �yI���s
2�;��ٯs��(8r_p�Ξ�����n.)B�)ԥ4j|H��D*��HP�D��uս��:֬ݻev6R�kke���Иv+���r5�BhNm�5�e���x�e��k��p�#w*q�&l�ΩqTN���އ;m��ێv��.sp�z�i��ĥ먒y�	�U5�X5k�BV��m��	Y6LyW6קr�̓����x�M�2�`w%�.:<�����V�-��jj�͙�[|�a�l'R*h�u��Pf0ͣ�p�cD�`�E��&���(N����.!�*�r
m��ex�o!��}�W	���sEj@�,V>�/0��f� �b�7.�j�oe��yJ�f�J^m�[\a�f-r����I'YT��)���p�F#t9<�]�\�z(G �J�3tf�w¶�P�l��''}|s��\�o�\"Ȍ�h�Rcd��)X�u|.�bT,�,1�=�pp�ѧ�ɺf����6;��njr�*����ƉV��t�wf��j�J�
:I���1k�1�9�{�����մ
ɥ�9!���x)�����q��z����T���ѿ%��u�pZ��mr�t�=Ք�R�	!�܍A[�Q+k�@�yǅ��ī�o������������m�\�������"ނ�Z�gÞm�����w��9��d�x�P��M|�̆�d����g��ȷ.�TJ���x��I�+$`4��\B��%z"��eV���t2�����sSm�s�6~�d��iZ@����YMW�޼G��vQ��V�b��捗y��!�TK3FwO`5��5�v�Pj��j{K�,�ͥ�-����� �7.�U3�̐Pb�լ�F}���u%!Ն���3�3��;Bh�-��]1�8���בA]��o��z�Ц��A��v]�K:mظ�%^J����ъ�;��e�+���i�mi�V�c��L�K�i���y/'8����)��u�s7c1їIx�{����W��s�Gb,��Fا�)u����ʌ������&F�p"sB7J�N��JĲ�<3�����u9��ӹWŇ/U��c"pk°tJ+۔U�C��P���%��0:C6�:�<��:ۘ�PI�"M^]�	Q��w2Cy�W��i��{P�b
t���;�S�����T㚤8�c�RU]9�7�¼o�V=���MH�0_1{1vs������S�R�|o���0u�5�L�&p����gd��đ�*^f�S�)�)ܺ��U��=g
�Kb�)��RC�ڿ��n������d���Ծ����\�N6wbq�g�ٔ{�]%Р>CA� .�?�̈]p�����*���z�lZu$�s�q�D8TT9��UH"�r%"rsvY�jaU��w����V��8��*9�DvWH�+@Z��UJ�D�LC��
/D9TQp��:�&˳S��-1ZQ�+ԓ""u.�PR����I���Es�wdE
���ˇ�듙z��1YNMʜ��9�.�$4��TT4��Gg��㧈I�)W�tB(����!��w=Ζs�̡-"+A�k�r�]vY]�ʬ@҉F�K�qP��r��+3s�u�*i��7G$�F��u�S��h�a%)�F�+)4Г��܊��܂�23����-+�Q%��d�Vb�#�«�#4�#T�LCL�tT�'3�am��"�U"�Y���I'Z�郻�	�����e)���4$®���M�Yi�NEҤOt��("��G�rL�J
�GS
�y� �R/:��r�e����i��ثNb�C�b=%�eܽ���N4�gA�`����FVЭ=Cs6ۙ�OU�@9��W#ط1>�_|
��=�35�DU�O���/㪕Q�RH�	n*�YY�>�V|@�2�@��=����z���@���D�g�Ǟ�X�!�P�6�#���g$�A]y\p�7�f�Lz�]zf��(�Gʬ;��s�\�_�R�H�L�눺q�w�_�_܍����N�:���(�O�sC(��XA�9�%;�%q]��%AF�
�z�K�U�u��W�����w!����>sD 7 ���ֲ�=!�^b�e����حB�DZ��pe{q�Lz)evo��=���Y�~R�4l�k��Pwë�x�s-��uO���D�R ��܅��H2�q�:u�j�L����"tW:���{|����i口w,�a��k���Q2��P���M��V�;�ƨ� "ќY\�u�W�느!}2u�A��5"-<(�㇛<W�V�\q�v��n-��҇�']R\z*��W���>X70��+x�ͭ������R��~��9OdqД��*��>Љf<��E<P�;ي[���P��2<����	�a@��vb($����h�:�uu!r�����Ψ��.Gw��5f'۵zu�a�q�}s��Y6����S���ݕӡӘ�丛�z�������Sgt�Z����"���w}�W��`J́�f���L��P���:�9�O�kM��sڱ�k�g�.��k�v�t���JG��Jw`�V
���ڦ�r��s�&v)������5����4��8��;�1�!v>�í+.a�c�V.ˡ ����r��K��� �3����M�$+Ś<�."k3w���]���ǵ �g��W�GL�y�u	����a�HԳ�7��ϒ�tb�٠�َD��2֝��>��˻V|�W��"��~ρ�!�v�~,Of�E�j�N�lep�˞�����Sb��n�2+�ZP�srN�wTt�IP���"�Y�ӕ;���RO��e�O�[�m�2�_,܅���B5���8��k�e,=J)n K�P;J�zģ�*v-���wr,��[Nu!W���K;���(*{��u�;9�kk��y�G�0 ���X��nא KV9��v�;�9S�jvX���������W�T]��B2h?z�#�e�rO�Г~�ۑ���9��I�W=w��6��s����VC�6:��le�����i*!ޝ�|����u�;1�ΡNH%҉F��B'�#҅�吥�2�#� Ӄ��鴝z��,8y�cK $�`ٱ�)�s��!�����2��6ntr¼�[�����v�m�8J�ֽ�5ks`�b�-�NUOx��>L�4Նrdn㋴�<�tz�S8��l�G����Tok���u�����"xd@�j,�qg����݋��JN�5��w^gZ�.����P��t$���)h�����U­?�j�8��1��,�C�>���A2Zv�����:��AGN�� �<�s�u�����۬�= ��cpԣp�f5�u֩�����0�M?&O,�}A�R�F���V�{����ʯ #�\H,�N�hb츇^t�L��͚�r����L�V�D�umR�7:w��}ݬ�����P_Ӕ�H>��G`.�Ĩu��1�;���Mg�i��Yb�\h�g��k������Gp��7�>H�p�����zU{v���� vi�vg&�c�^����iu���l�b^VHj�d��� �/�}@Uع��F�"��������Ӆ��自ڱKdg�s��3I�4���0D�D�(
 k��z�G��Km̃��	ʁ}����\2v%�f�BEؠẈ��Z�e�&I3����L�mU��/����u�SэE{��
��u{�#�M�k���d���bj�)�v]A��+��U�Nn{��6X'Ƣ^���Sp;ԋ�q�%�>�pu^�<�B�SJ����vk&��3R�"	�r!��c5kn9��[�5��R4�nG��2r���>�Fo�`���g����Ƈs��C�'�'Ü3F���a�9,}l<�C�H��]�ԍ�p7B�^)�R�mG��i�4��g
�s��l���m���k�]YB�0�� �v���q�6'���+��W]e���E�[:|�w�����oņ��i���O~��;YƿqW��p�#l�=[+"�s8l��d��ȓƟ-��Z���.!�oc��we���d�,�}^��A��>�
�Ј�%��� �>�@�gŵ�����b�����x�ȟoG4ʰO5��5��M4��`p�o�j�:A�E�4"^�S���:�E �&�)���'�q'��>��#�mgS���"ݞ�+��,����됻��\��8����ۏ����sb�9���zܓ�
o's�\�Ν��Է��ϦRj������'��}DznH#�2k<�!��7���&��ey���LQ��_ 7��3����LD �Dpk·Mw��caGhrh
�v݌�ZY~�h�a�tD����5K�V�ND��,�����4��21b���K�}��5{N�`�K�H�I�����rl�;�"�ƤŢ�5���b�L�� ���I���,�;I���Fr/0H/l)|.
���n�PZ�n�hCs�bq��}:Ug�3�@~;��8$d�n��q<��(�ղ#ȋ��_r3�U䧤F�|gr��Gb�8���͝;b9�hZU��-
#���y�${�G��Q�9�����+ �{˷��\�Ga�Sڅ9y��H��g�o�4��u9�^0N���|�K�J��5��F,�Z"�t��H��&Լe`�9,�}$���6���֡��l�&�;�9B��2APwuv��ѕ���F�;�l?rh���Ϩw1��s�{V@�a6���!�񭆖ϊ�b�qGr\�-�rA��Jْ�s)�A-Sdue
��%�9]<���Z�ٿz�ObYa!�Uv�n=����J]q�tʈ�Ժ�4n2����J���Y�|���s��ε���B6��o�rU)���8�����¨nY�wɱ�-��Y�.��i�u���g-��l9��
�^�cvj�iOExv�X���ֿ2���-��s��7�/�>L���b�=$�@�d�s�j�s�s-���>�Q�*ȥ={+1K�ƚ�����Ŏ%{pॉ�g
	���Ipm�}��M[ΧN�$�*wa�h(�w�ܲ��2f����eʘr6�n+�	9�wxa�$U�@�wX����tI)Dܭh��`޹�+��G{���vX�^1�"�8�$�7����9۞���~�c�!��#+���d��i+�[�� ���9�n\q��HkwKݺ���;�4w/�� �,L�-��^VX�j(M#�Ӣ|��G5.�g8l��Quw��^g���A�(9�g/�S�h�HF�),K���:���e2���*:��Z�^4`���VdĎ�OU���x��$S�h%<�+U���<M��������3z�ej�ܤ)�P�"]��ϢSkM���]�=�-�pϮ\#��<L�e�!;-I�3�ټ����<�Dv$k";�3(�'ݎt�� �!���[����$�F��Z�z�RE�ĜV�g`��U���m�@Q���z3K��gWmp����[�HD�����Z0ݾ��-Q��=qd˧Bd;�^�G4#�\�Qܶ{�̼��3x�Y�+D+��3LM-ҳr2���nC�����`/���T<O��b�|{^^�[���Ȃ���Z;t���3�ؘ�ܯS}"��5���q�wTt�$��W����;b��+O��n�m1�ASs�x�ֻ.�$��Y�� 	�^2,mg$�Ѵ2m%�i�E����,�[y@ �mTl$���:��F.:jntn`L�A����#�F�V��b�����+*�V#�2y"��l���sy�X�H�]�k�w���Fj��ol��������>
|p{�,܅�<�!���]�v;����P�	f�Q2"SĖ�O<�ozz���G^����ZM9���-<o/l��]N��߂���
��g�C	u�;P���AR
x�#tCP�t �
�ܮ$ϲ܆hP�59δ"��³S9\Y�YW�+���{_W�r�s0�)@�R�O�ѷ#�.2N
��N�ڻ0��ϵ�{<br- ���WR|�V��}z�l�>OYµԏͳ��{��ש��KU��R���"�m ɥ�7ѭ=�;�3��H̠�i�S
��"M"`󠖎fi"�����6�w�*wE�����L��ݣ�U �-;\�kx:u�'�!j�=�dfT�^UGV\ɰg�ޗ �>�TKZ�>��u�LNs�}XÞ7a2yg>��TS^ت�f%��r����$"ŬI\��`��kbr��R!�u�N��f�xk�|����u6[�.�>X���s�,Y���nG	K���G`.�ī�k���>�=�hMn����T�ЋQ5֎Mq�g�0s2�{�vnD�6�A���/��)ik��{��iy�ބ܇�w���ƏN�mٗ�U6�,c�8�=S��!��ۮ�:�����Wk4l�R2NZ���zjP�}23xEk�pY]�h�b��j�6u�Ƕ��=����yP�.$��@,�x.�¨b���"3T�{��kopO���U��Qz�`������:نՄ�l��ɞ�!G�!-j��r$@�ZDc�(�7]��yy��ش�jTiC$om9\����SI�Q<�$�q��QJ�����Wg����ڻ�#ٞ��t`Ȥ��(n��]�Qt�BIࡍ�G<W�5�S�@�
�=s2������P�\�|�B�Z�62\�Sc 3�1�{�w:�<Y=��זu*�{uz�
\}�/t������N3H�it�nг�C������m3�\L3�ze������&�VK��on��J��ة��q�Y�R������,OuB5{�Q�'�bj��d���'���eS�3v` p�8n�h5u��x}���j��4���?�uj7�E�@��[�kc���ΐA�tw C��{L�3�4�&�g>�f�b�I��#\+WB#������3љâ��O���t�ڞ��/"� 27�4������IL,R���@�~�{��`'��~����}�fѠօ8���l���YS')a�,�{Ul�����|�N�i85�ჼs��µ��o.�h��}2�`��)3�ص�ȃMq���&��]d�[y���8Mҏ�;�m��=�)�z\¦�j�Í%w._N{9S��At0ePh�='�_�9��19�3���@s��۷��u���x�3��I��F���5�h
ˣ�q�����Z�r�g���v����m�2D�VE*n��vu��&��_ݦ�Z%�FP��̯���=3}��Z�dS�x*�Q�@���+ٕk9�i���au=��u�}��J[>����2$bˢ_J�UqM=�^{�f�����9����L�w��2i�F�8�Q>肈��["��i9jl���u���_KB��1���Sٳ�lG:m	V'��p,�܅��n�e���6�]��w�Sz:�ͺ��Њ9�lm9��]8���x�o�5i
亼��N\��z�c�u�3�(�����%^��0�����]]���4���X%�},�}i+`=�$�&�x���	$��s�Oe���ڱ������!��z�F�֩�>��y�'LvUV=q[��&�0�O�p����sD9^5���}جqGr\�-ڎ��7�@����-1�ͤ�����፾������ؙ�/����ޏ�� J�du�&$H��[��C]��z��s)$��ĭS��4���R�k��s%gC}W��U�e�瓳RU�8A՜S��M�붑���vħWf��_��G Y��9��pQ���/}'��X�Is�2W�����"�!�3UJND�|�=������˛�f�,��#c�&3N,��	ݖCY�G"9L*���M4�^��l�J)��ީ�ʰg���(��^&n_�=Ҽ'�mz��s�]=�����,�����̬af�c��Z����"gv�C��
v,��+S�K"�' �u�A��u�Ne���)��KY������k�h�,�N�Up�g�=���_��Y�����|7͏��1���ڊt����%����s���K���᥯�m�1�$�ߩ�����P�,��T���z�b\ۊ�˫=�#m1�̻�tB���r�8v�T�UN��C��,�]^�x�{ck�ݑ��@Z�rfLO������a����u��J�΁`�� x)("E���O4�ݙ�8�qgˮ��x����f���r֍��ϩ���Hmě�t�qkj��a3e+�;QB8���Ⰾ�s�M���x��g9�bG���v�Z�v�bMVo����`L�D�984���>�o���*R?f�Dٌ֩�3}´U�0`Q��%�B� X-��8F
����̢����72�$D�"�k�+!�^�����1e��_�N2�^��� aT��QV�]>�}|ȓ�NT��5�����D���R�ge
�jZG�s��Aٵ%��8p� ���Ek�Y ��G%�8�^0�=�:V�Q�G/[���v�.#�]���Y��B��U�SQ&��ֽ�nԴBŋ���¹Ӛ�C��Zv��<�vb�������9��!

�V��yNS�8IT ����!�;g'5��6+�	�v�z�t��wP���$��F�a2�-�ˬR8xC7v�i�'�*>�ԵI|8�Ј�����u�=�L�J�pU�AwK/���V�D�e�>j���:��?f��C��1&���K�(��R�H�[³(�yM�ؔ�c��D��^m�Ә��3e���k��8M-t�a'��g9u �^_ʴeة�v�8�a��WX8��<�#�pfZVb�̣�6>Y�p��XuÒ��7�wuڊ�y����KJiR	�����`������T���<(L�Y���R���X]���9pLa�s�Y�okh���@����G���έ��
	��'�7�xU��>x��+�坮B!<Fi�)4�̛����&=譇���]�֤Q�CL:�ʺ�u�,w���S�!<��U�v�q����֏w]��2��v�w5c���]���*)'5+�r(v��\��9ڸuN�Y������`p���-����i�P����z��B�O��i�qL�o�%<��Q9��:�7J�%!�۸�:O^}�b�P8�J���Qw��L<Z�d�rvZ�'��ٙ7s�6!V�9j�^b+����l\)�O��!�rq��N�;�z�v�S��eU�{%K�Y0�-�[:��y ysvR��r���@�tQ@���&4<1Lz3x%Ʉv�3���V�Sx���p+},���mb��[�E�-����Hν�u���N$���x&�\�*�f,;����s�:��c�N2C:�!\�T�<:w�Xf��ݦ^꨸l�Hɧ��qfFY�1pz9mmJ��ƥ{���UFtu@u5T����w�\fQ�L�T��`5����K��jʩ��ojabA�R:=�g͇���r^L��}MX�١��5F.�if.���Sw4\t�����D��p�g��c���f��Ӊq�\ҍw=@6�&G�q�'��1x�2'�TM��+KѯZ�ϐ�뛝V�9�l�"�1����vԕzN}��|En�9αd	1�=���;���+鵫���\���!Sqe��ІEǴ��F����*m�]�c���ٌ�x��C��|nf�p��7�E�Τ��-H�Ν�ufmI��=���
�@
��sKUD�)$��Y�w�t"J�iRFwp\�X�R�l"JL$��0�*�0�P^QЊ"�DW\����%Ts��wp(�<D6�V��V;���e���Գ��K3��E�G�q1n^�f2�"Hs���"Jy�<��Ed�i&`�9��<�Tk�N�{��L$� �����ʌ�&��.Q	�vr���2��)[er���Uu�/=it���AAZ�EF%%q�Jk�
�BΡ�����@�U��Y^����S�ڒ.F������G=��DC��PGuBq��Г���(%��@�եI���N�p�­-b'UD�b�\(��#��SI3"(3
�:"Uʫ�w!]�����<ܜ��*�1"�TE��9.X����G��AE$T�N:�DT�d���h`QT�h��y;������`�}�*)�����iZޥ22��I1�����W�� D�Dݥ�[�Y��5��J:�>G/�J�Yyq��w^�gB�4�}�ȏ¼$��*��9$��?y��1;��%nܜ�^O���|��C�=q�*|v�F����a�����=x];H!C���3g��ȁ�ͷ�_]�+�y��wr���&��A${�<�����AA�}��Iz�@YdY�Rp���]���G+�M����ۺ1;׏�{q�?&��9�S�#H}�ő�I>��#N~ӌAS�c���tM�L����<��{��x����A���߻�yw�k��7��w�ߐ�;^����zBI�7�<�~���;�w�x@������&������
��0�E0�*@��^ԡ���f!(��㣇aAO���
"ݱ�$�����}��{C�aW�}����篽��o�rs�۟[����yq8����?X�}&����������G��aj��I��������W��
M|�8Mf�g���ϼ����\z�^��r�G�>��I�!y���w���u�(�}����>Y�'��E��}������1;��=o�y8}�"��P|�{�({F���?���!�V�Ug& �HG�Z��!�	#���z(��v�=��>;<��i=� d
<}�"	 ^lxId~>�����'~v�}��oϴ��]�>���o)���|ϳ�tD� H�j�����*�Q}��eV�|�yr��rF
"H��r���ߓ�r{C߮��U�\x��!ɇ�z<y��e��ݹF������]o�==�����k���#�D{��<�}$^q��3��¹�};�϶�W�@Y��O��I�]����w����q�\�z����P����<;��C��c��]��s'�}C�aWo8�C�ohI����ߐ���g��N'{����O£Ϧ/�����������6G���{n����D�7�ǉ>��6;�����Ą��ǧxw�iǧ���ù]�����]�&���z<X<;�o珪��"��'�}ԇ�Q�D>U=�޶F���7�R������x�HO�s���������n;rs��������~�������0�~v�G����I��{w��yW|v���i�=;xy��ט�P睹9S���7�'�7˽�{s}P7��F�Ȧ�2���m���?ch�7t:��mzi�{#�l�ܻ���#��^u�S�R�Ǒ�X�4ة\�y�n�"۱Q���eQ�#}8�Aؔ��z�хLu,줁�����V#KE�t
���4Vh�8�fem�op�럽du������;�ϛoϔ�_�c��˽�����S
o�����yw�k��t��r~M�9���`�����'���?!�0�����������I��۷#����}}���'�ۗ;������#�#�!��q���[���v��M���߯^6��MC� |=g8�� ��G��Y���� q�������@�+�m=��ݹ��t�^�}��}�#���H
 "=����7|��rs�=o�q8hq�=�=$Ft�K>�"���Y�������;HR�m�ӽ;#��z�������螊*d`���|/z���}����l�x#�#�a��.��S���='��C�y(?'�x����Q�'��7�۷'!�ww����7��}��S�;^G�P�,�HZs�5��eZ}W�v�����U�ݧ���zO)���������yM�	���ޏ��xM!?��Ǆ��1;ÿ���ŷ?S���Ν��Y����aC�>��˽�]����| ������Ull+����{P���#��i| ���@D
#��+��#�Y�hs��߻x��L���_�I�ޝ����o	�!:O��ǏQ�7'���<;s�#~C�<;r������NȏP��F>%G�+��̍.a�"�>'�&�O��&����v���r�� " �}�
���>���|��xM�	7�$�w�Ǩߐ���ly@�IĞ��_��>xB���s{H���r�u�ܷ?7ַ�޲��r���ߓ˿��'�|x��w�i�z��d����>�����3�0G�Ͼ�*��ɿwΜxw��������?'��C���~�x@QC�~}m����T��E�v��ޟoV����;�rcs�ۓ��������ǚ�C�aw�_#yC�~�|v��v��=��}O)������������^I�<���{�ER��}>�K�fH�<�ή*�머��Ϻ�J`i�>�#�Qr��;I�����Pyw�k���ÿ'8����_��0��|q�^8���90���8|0��:��Z�~#���@����\Ǩ��G� #��r�,z]��<�Ez��8���M���u>t\%���9��ݘ���>����O;f�F��F�s�mn�f�1Xz��iu\{���+�����s�b�Wڔ=yO{:�ڃ&�v<�f@ԝ�/	��K{�7gc뙚gc�AF�iEw%1L7Ԭ
c���΍�\����V���|3��(�}�b����]��@�����8]��CǸ���ˏ%q��M�99�k�F'|C�$����]��<��w�~w�}슏I'�H�ah����G(��guDnB�xt�� A۞>���#�Lτ��=�=$c��I�{̈���Y��2���D�a���C�$z��Ǔ�xM�����X$�]��.��8��>g�SF��f��t~�����~ޟ�>��s��s�8��㟈r~�|�vQC���|C���V��{yw��n;rq�1;��n��{���zL*���=F�� y
��ە��ד� >"H��a���.�SΆ}S���/w������n?¸�����v��1>�����ߟ��}���M���>'�y@�$�?�}���!��<��~q���������i�>��zA�#������SQ��e���t}Dyq�wୟpI��}O'X���'zq䣼[۷&������ۿS�w��������3���ü�H��xp�];O����ˏ�%w�ѹ7���LA���`�(���R�޿Ma*����1������yC�90������ÿ!�=�r���{g)��o�"��>�!^�
>G#�>�,�xZ��:r,�Y�Z�t}>�ƺ�w���I����g��x~�~֜h<��R�;}t��z����o���~�J�S~w��q����\yy�;�s��N�㓜s��z�U�E8��q>%�^ۏ
>e��,�Ϫ�O���@l۽?b�T=�;:o7��'"���!ɅS���6��7���>���G�nW{q���P$�뷷�G��>;yM�O�z>��<��M��>]�;�����ڭ�?�y<@s��Hx���'�yG�'��߄��y�_|�����_x���i�����H��K��G����bO�|C�=��
�ɧ�hw����($��=~��y@�����<y��nM�>�;�����,(t���SHD.w\m�v��Uz����{����i7���|�\.�y����|H>�"N8�#�G
zG���G�￻yC����ސ��w�}C������w�<�������~>�����G7�S�sc�J�+Mj��ek�p7)���۹�qB���+������\�ho6�fqq�ӏFU���%>}<"7vw��Υ��6�U���hf�<�{X�Uhr�f��v[t��ɲБ��2�Ҩ�Q+��)�:��bޗ���-��>�����㓟��χN��&�c�S�nB@�_]�'�yv����m�<�ߝ;�����~B�m����4�7�y���I�!}�I~�&��q����/��q| �o	���gs��v�}�L*��'�<>o�m�;����Aw'&~�c��#!Ʌ�x�=�_�xC������>;r�þ|��ԓ���>���v�~B}_�x��xW@��j�m��O�s~�;�3_@�gނ;շ�}���]������)�ޝ����]�ҡ��M���{C�V���Sێ�w�'���!��yOh{C�{�c�ߓO�	��<��I��K�QުJY?Y�+�'�� d#�mϽV�Gނ=k>� �y4����7�$������c�.��!������>[�o���>!�W�24�"�#�hx#�"�ہ���8��?}�*�O��3�k,���������L����hw���<+�hN�{���)������@�,����0>�E|&���{�zC�
���<����z�������Ҡ}Hv��'˷#̀������U�U=v���~��$�S7Gד|B����o����� �� ��||/j8�DxO��H�? �?���q��Ad|ׅD����=���7�9�������1/Y�i׺���իug���^�#��v�w��2���~C�o�ÿ��ߝ��缿�ޓ������9�����X��>g�I{��ϥ��x��fN]��W��M��������y����>�4RKf�=�{�R��$�#�D�����Ǆ���9߃�+��������$=/����R|�~q���k�}� )A�$�/���c����A�,^Ϧe�s�z)bdJ��E�X��;�!�k�
dW������G.�����W2�ė�1�;ǅ�1��*k��"��_F��Fs���_�T�7*`ܨ A}��X���nW�H�f����T$˃-o�A��ݧ�n�3�S�lB	��_m'��7u��P�@Iv���K4ug5I���X0i��o;&��nWG��uܺ*
�u��y˕B���5[a%�a[����%G6�X@I�׶�d���Q$k�m
�ٿ@��H�K�ڌ�������:C��c��^�mzY�S�h�HF�),�"8�YuP'g$�\�N�6Y#5���NY�S�v@M2��gu=Z�i��7=�4����a�塎2���x�O��)��I���`��+أ��vL�V�ϢSkM���g��Ŵ.�����Px��^c}\�z'��T��"q��j�H�Dk���H���N����E�C9��y!��o;��y��5'��Ab�k��48�� w0��Jy�nZ�=��qu�|r&zg-wK[��=t���J��&X]-!@�G�|��]B$!�8+��@YBB�v6R@�T��滮m��O*��X�de{�C�#��)�r�8k�����.&��1|�6��,��,*�wz�X���f�����'�����tkJnI�a�Q��RJ��xL;Ħ�����Q��=�%�J�Yo��LۛC��Y�Ry�F��|���s]�DLS2r�<d���i����8���7�ځ<)� �����Y�6�u!^��.�$�f�7���F��ځ�g�K�|xT�� {kz��6F��:�%.o�����ZoF�!���\M��)P��I��OU�hWyJ�]���	W���g������'t6��t�:oP�R�w�����p3&���Q5�*N���V���$�OG�L��]d��3i;Y�˜��~�ooi.������>C\�*�D��f���[�Ȯ�h`���]El��9�;�Ī�ٳ�
}s���9�3�����u�	����E�R��	>�Du�䗷'��2�K��wè�Aǯ�+_N�Cj0��\�I'���x�^^�}�se�:�,^�Xp��ΦQ�`YTZ{����x8�3)��X���@�T䮋uiS��gIV뚧+#��]A�PFv9�V',��d��sM��:u�'!��Y|�œ�_���b�>qx�\C3�;R����.� Ō�L���=}�]��VV��ve�7��T�>��'{SAx~�c�T<I��P2y!u��������B�� �zlZ��zZ�d�;F�͡9���L�
��ϧ(r�|�ę]ӉPk��{K�J�D� �7&����ʍN뼼1n��S)�C���M�yP���#��
_D��@J�E���"�*=(��̩�ڻ"3T��g�7��+	Őڿ'se_����*�D�-w| m�W��m��73D�_�nʗ1�g�\�hg�U��ί���+���������	�����xQƵV&RPg�3��-Gb��Y{��p�d�]�V�L�M+�K��)̂�]�]N�2��	�+7�7�P{W�x�Z�B͜���� #z�t���y@��4ȸY�gx�ld�Q�`�u\�u���@U��H�ND�z�����}'3C
 OW�M��i�b�;�Pݎ�]�Qu���I<2��`�!�Q��T�6�j���̾.�,�\:Lc������CGC�=��c���uR{.���]��s��m�{��l|������b����ҡ�ڽ���ͦp�t�ގ&�u������`��q�v�8-Ns�Eb���SY�ʣ�R̐�*�
�eG*�2�tѸގ���*���I:q9���`ELQ�pxxj�ԿJ���Z=�,y"�n��]+8�]V+
a��_�@�״��i��2o�W��{kb�H:B�M�F	V T��s��O\�N��%Ꭸ%��/3����/"�9�>ގi�`:�kL�nL�Avq�;��*�P�FHjH�7Jfh��Ƽf"}��yp�{�'>&�8dk�1����M�ە���� b��w,V�ېm���}<A������?s��]�ꆝ�{$���;U$�j��+���_9t6�3O롄m3F#W��ڳy�p�� �meƋduR�B���':	n@/�u&�y�޺LŒ����s����ɆκB��;��������lE)�"�i�QT�E @�ۅ��/X�駜&c����nI�μ�(XtJZ�W$�B�^�&}�i�%l��N�YW�Ԧjj�W���-r�_��he[�{z��9^�t�ɏ�������b�v��k^Q0�Xo��H6�Ȭ���# *�w4H��#t�yD��
"m�^>�t��MCҮ��+5W��
`�o�fΝ��M�~J�>W��Y�nB��3��J��ۚZS�O�oh���0s�5}�BFz&._:���=�ٵ:_��E�H�$@g�Ĵ���Y@��ys@:����J����i���"��H����R�\뜰���[��+��λ��07vZN�\2uߧ�W8�<�J�ag�R��Va��2Ǡ�"��݅��w�mcڊCǗ\m���F�'�x�}�y�����T݅loL���c����wx���(xt8���lq�deԎ���_�\��d�^S&}�mV��0稜�Q7n7xۍEZ�%ʯ���w �Ɠ�}����w�On��К�io!�'�K��Y�����o�ј	���R�a�L�۽�[�xl�X�����F�u.�-GD����R���1L����Tv��o��@����),oW��)���+��M�J"�o9����֤Y�$l��o��0�є��:Ro#M��f�_�|=�c����;����$.G�e����"�z�cSJ�rx��[�۞�Ƞơ����'{�Zu�J�����N���\
��	lO+�Yd�s�jGN��@��pQھ޷�ԓ�ܟY̐w�w�Эr���@=,��/���Z�/o��D8m|�����Ƣ�*���4�����p;�Fߛ��r�����eZ�N�'�Q\����s�l��Y�|�@�Aƻ���k^4:�9x��w@[��:�1g7�RB�),	�H��"��6�:�w6K䎯�d3؂kZfLNwS�z��_�{�O��5䧗��t��gN]��݌�Q��D�`E<U�ZWq�����x�글�3��W<Hqu<*Jc��K���ξ�s�C��s����$�"�I�Or�⠧���L�Vô��X�u����VU)O��n��F�{�<�{�Ć�;+e.�Ô���dmUN�ľlL�ؔ	��n�f���HQf�%!�Y=="-!��qH����&��\&+U�����+��%]��Yt�`�fj��ԒK�,djN�X�e6��c���טG
]d�d��$4��\��� ������E�һY����K�7T]4�d��GÍ��h�t�4
��RM:�t�ig��	����Kq��]?y�{���dgty�ҝ��p��@/��E8���;ı`i����<����Վs<�˿����lu���d�|��]҅@srN��#P���WDP~~�;��.XZ
��W,��u��/i����Κ���gP`=�8[O&Mv�3,�c��+N.%�=�,AN�4	�5��Hڳ@mt�B�y
^u\�­���j�Z��3 ��E�(�)ٛ��/)��v���~����,�p
�C�@x�.8U�ܮ$�k�����Νc%�^�T(�Z�T0��B�s6�K��>;�MS�V*��~yجΈ��c��-�����zE�bZ�KY{S��������7�(G}a�Iv����S��Y��Gn�1��WT �PX䞤�iO��Z{�w^giƑ�NF��*��̐O=����2M�3�^۠�GvnQ�f���9�ap���iڡ�]~t�ء1�D��Ǚ��̜��<(��� �0
qdd�Ե�Q�u@�3�3����ꅩ<��K��^+�}���&�w\i����^_m��8Ut�}HJ��tz��bے���^>R���_*��T��M¯5��'md����^$"� �����#��r�g�cĮ:�����j�N��rY&b�ut�Flq�F֙�r�\��ӭ`���:c��oh�}q�N��2�D�VeZ���s-��dkt]��Rf�2�]/+��m;��U�/|v�T�5��AU�Vc{�Z�ƥ[e72U��J�tʳ�Ec��MX2t'��dѼ����kE�Ԟ^�����ε*_i#��ԕ���i���]`�[^�i?�go�KY�ɖ�guYpL׈�=W
��qk�w��wZ���MOt��<����\ֲc�R�/nU�܋׷/�9׊FYҕ��_EF�]Q�|���u_R�0�콀Xt�3m.{4�k]k*���PN��l��LIqWa+��N�M��vay��Ve�Eob�9���DQ��l��7W�
ʸz���Kّ(�[t�
��F�.*�6��j���Ra��1�.����y���!���P�Ĩ3姸�yo���<ڠ�ph]3*r8����Ơ��<���x�q� ���ڲtϦ$���ԧd(7����E��.w���7����Y-9ND!��1X�yL�ؔ����u^KE���)�}��/�QJ�
Bf�^=�k�݀�1��.�Ѣ��(�����D��ʕ+d���㷄YLq��7_�Bj%�7x�n�rӚHV��Ҩ&]*�樤��8�|��ӟ=�]���e��*���jI^����q�f�j4\����f��=���ŕ��u+r���s��[פ����?x��Ub�],3<��kV��F�Q����+��S�S4mΐ��,���_N堹{�pރ�\��rS#���+��c�e�� ���L	>�W,�K?*�ɜ�%�m��R��!ε�c���JBE��H�v�7V{F1M�P���n`���r@�Z��+˪۾�"�Aap��S�]/�n�+<��>���%�;�8�A�F��������e��Y"�� ������}t��Z+��ǋ���mq$M�խ�`%7[�ZJ��(ehr=����L�֋w(�|�e�Y�G�^9� fZ�ط$%�����n|.È�[�ڎe�$�lf�D�2narr��Q��(.ПKNg]��3G���5�3;�1�ivۍ�t�5��;c�(G�'WQc{�����BP��g^�w(�X�"�0�5�%�_:��hޮ��S;K��(�4�m��_
Ǉf�¥�0=����R<���bQ`c�)%��n����'q�,w.Y��S�+�k������^)΅�I��t!�M��v�Y��r�M+�W�����#u�oN�����U�>��Y1��-�y�P�$f��k�y��\y��2�]�0M|�&9���W��cvR�����m�L'�>��իc.̩}05]dT�����������i�2�ڟU����V��ʋ$�ܫ����\���X��[�h�G��r�+�霹K-C�h��-Ŏ(�\�rDҳ*4Qa�j��-U�xB9��I&V=B=�A��9��W+� s��"#+*���E�L$9e��Ouܗ2�C*)u�w\D�� U�g�QQTEfC��(�I�dQΦŔVr�u�ADG=G\���X�f�y��n����T�5OqwS�-����RG\�"�7WZ2�G�eBG��t�f���ܣa:�'wvz\�<us���t]K3Ds"]�Ȑ��
�8��qn8�NV��Y�y&^����SΞI�5��4ڥ���EJڱs���3�*z�W:�e��Up�M���R�C/<qO]�)CN�.�U#,˗rO�̹ʔڛ��J�Y,����"��s[$4s5��rEbQ�t%��:Rzd�yŸ�sys(ϕع�$�� �in��.c�ǁl:ũWN}]>�L�.�����]�� ��}K[Z����ɒ7�Fr��|~a��C�L� d�B�Uܫ��C��ޙ=tlm�����z�����9}i�WAdw����f�5g�;�32�p2XY����m�ʎ����Qb�:�.r4�]R�g8Éw�yP���N�#��)P��I���6м+T^�%3�v��Ǡ���]&6��>��=�Ӌ!�i��T�yI
�!�Ի�¼�	==�oYrJ�;��"u1�GOq�ϧ��낎;	�$3�8����%�.�b*E��fv_c�39v���48�)WuEc)yW��	�� �\1b^C�7B.O
�8��8Z�����ݵ�U8ND��C�	i���H:A_l�9잗�qn�ϴʥ�j����n�w)��/�eU[t�}�����
�\rLZ�f/O�9�V��^ܺ�]j�/�x˩�x��o��y��hX�Mp�
��q{��O��i
�����h��k���
�ߛ5�x�V�0��E�r9���͂���|�P�\V���>&�9 QY��&޽���
�D�9�o�R�3�EIL~�]�g��Y�5R�n��"=�Hx�h��6��m�yM}���8����Z�p}��d�Y�t���+�R!��<��F�g�8(���n�8�º-v���P�.�QS����`�W��ﾫ:wq���h�5�Em�,
cy.W�
״ɿtδҰd�,���~f�:c��=X����*ǫ"8r҃�/���ti|ǹe^s�b�*�C�Lu�難+���`����o\�G�SM*��
�^ڨ��Q��0�2zO.��h�&�Ո�s������U��E��<�,�pӮ���4j���*������~X	J��oVj>����.��7�� 3unI�u犢cѨZ�j�J��ľ}�nh�k�tq�8���P�T��x�C������rOb�[�G*����,�� ����k���u���3ts=�V�P�/D2B���)5q@9�GP㖷�"ئ��8�Pl3{�N)W���y�w��*�Ș}H7JĆ����S��\.6d�� ��f.��y9��;�ԚGN�\+�*m�'�a{�$sе�I������4��r����rb��i�B�|�Yd�Ut��B�'N|9tA:�,	|cm	GG�wk��uR>Ͼ����g��_!2��zŻ=�ute��0s2��Zs(΅w�ݒ�g/5�׸h���g�"V�+NȒ�b��է�Q3/<�VL�n�s��2����ZN�f�`[MX��*Σ�-�OCY�b�/�Y=D���}����n�Y��8o�}_}Q�����Ʈ��S�I���l�铮���4���Q�V�Ș�%��*���e&ĥ
lGOS'!L_'����B�'��N'~�3�]/��Kd�ž��5�8�̈�x�]\H��	m��5��#��I�m��m��NmL��W>�\�U�ZYV6aA�WVB��}��T���r���0�|i��:8�c4�ϐ�9N��(��s=QE����	�9�툹��z��`�~�Ӹ�K�������c��\�'�W��.U��n��J� �;c3/��k���:�4j���<؞W <<  h����{~�Xq3cj�`9��tǮ�J���1��rO���	`���vBV�#G�^9���@�g��������OyM�?
�J���m�0�r ߰?
=��e��
���VbmFj���q�12XZ�����.��ms��\T���T�u�\(�y���J�bJ�; U)��S�Xr�Ü�dԆ��3���െ�-{M�vP�x6Wަ��j�P�Z9y������Bq�ǵ���cZ8y:3C���J�V���a��Ý��Y{��3ZuwqU������q\�*3f��Nb䗜�U�͖�y\�t�@�c���z��;Χ��˻���½Fʡ�]�.c�C���X?�"#��m�d�j��XA�#$!nʚ�Ԛ,Vp������x�글�3�V�Dt�Lt]x��$�w�jN�w����堓���0�v�jSܷk���ݾp@O��)�pTc��W9�S�8�f%���&��;@�Ai4�O8��U�|��~;kǋ���G2E.�f���T��_P�� (h�RE�#��AC���+!�b�kWmZ�h8�c�Xg(�oRϜ���@p��7:S�,���*'�:P���;���A��=��<3yXx||�G9�a	��C;����:A��%��̖��V�<' Ң���=t�lSv� EA3��u�[�s~GZ�le���|.9f�-��b����h�%y����)8/#Á�#�!Ws-�v�Pr��C��I�S/��e�ǄԮ�K���<BJy�|*�OW�?l���|�E�:�"�J�>*�Q�ĸh96w�ƓX/��{��-Mf��ݐ�)�j4s�hS蓘�.=Nb׶9,�k��r����E���L�8���GX��c9��֢N����}�MĐ��{gb�i��GI�fY�X�kM����U���d��಍G�+��=BFce/�.5gv��4^u_R2���8?�Cs�>X�J��.��F��P͏��{�.f�kk�5��Do%�`2Lz��6:�6�^����Z+Q��vk�|&�F�/�V[�Zr���IV�)�,�y����멒�a�eQa�{�98��w:�4��9SF��vjRH��cP�8���`�ш��*e�
��'�Ϻ�9eW�%�k�lʩV�F��xJ����p"Ⱦ8(��]d��\ؖ��+dW�Õ���>����Z��G�&�A�R�8t�Wݲ;�S@Ahji-�q4$�B]�cT����pe�r�lg�봘c�./���}�C��\�p�W�}T2]�ɈQ��r0]	��q!�iM�������f�Sye]27�aĘ� �qb�D.�$�.�ܧ�B�u���7��g�JC�\B�1�\,�>�������l�}6L�Q�&^���@�k���ι9f��}E��?\��o�r0�&2x��Rڧ���p4�h'�yJ��\e廮����p�}��H:�BR�u��5ʼvxM5��ᐋ�/!ћ��h����6;/jz�U�Cl�⡙��f2ƱQ�u�� *��5�Aֽl$\E�-�wwM���O=�b�Y{Ι5����8�5��z�.���a��G$�n�-AV�k�C�۹ډ��L���Q�oH��o)��i��.������F2������ꯨ��#����3mB�� ��I��BZ5r[ �{r���+�|�����B`^�k�=��[��82��w[b%��/ c��6PD�B95�>��t@�@SS���T��q�.�ݞ6X75���"���o�E�CB����P2u��ʛ��=����D���4unޘ�J���,�&�\�	��9��O�D]~^t�T	̒����Vzv���aN��JG ҺE�/M�b�1ܗ#��k�d�,06&�P쏓Y��3y�L���מ�+y����79��hܪs�U��K�=%�_�C=^9�;ѭ2���i�l�f�mĴ�?|5
H������+�{U��7��
υ*��q�3��IB��[ ���1g�����t�i��N��N���1ʽH2�bA�9�vm��1ֹ����kK�Q!{�n������b7Bܓ��|�$pl�Z0�Ğߊ��z|^��$�5Ń��V�#5��
g���z�)������.ՍpZBܓب[�G(tϺAH��,[;3<fY��a��^7�d�ݦ�b^�%��SְIEV���,mK6�ʰ���L�
e�ksj���˳ս�`�5:�H�V���	�M�/2�UKs~r�qVkf�X�.W.�&�E֎�kS�Sy��َe�u�:_(��]��=��ꯪ�TS�{��λ�����)]j �-6��{�BL�]��|���M�79gtN���wSZ�S|)���O	�J|gأ��,C5vli�ΛB�U��ʼ�Җ�#��b]ꓗY�wZ�P>��Pg����S���I����qL�:~чYR:�5�tJ���r�zX%������5˚�\N��U=t�F��|NF+�<��{"�k=۪Z{��^�z{�ZL4��ޟQ\�"4�K�e�v�/
0x���5�̙9J ʹ��3�B�9���}5*��Oi��f�MļM`t[�hQ���'���¬�I��NSA��Q��.af�����;�z�u2up){\Œ�R}�G/������J�^��o��o°9܈9h�F�q�ƛW�UC��;���^)%׋��Ԕ^�@ܬ^���M0YU����p�З:�J3���]nO9o�2�f!����L�޹zsAn�S���}�Ln�SM/���/�"�u��{OKbxe���Z�<Ph�_�%i�5^8U�R���V�"[aK^`�B���iywN:%۫�yk�|��V�ɥx��NTdngCK����zz���Ϧ}��<��E��,���o�Ś���((���ZaKqŠ��;��=��|�9�QD�����1���ܙ˄d�����s�f{Ü;�@�8�k�n H�z��]N���`W{QW������.��'�Zm#\����dm9�,��O���� ��$��o��S��O�˃�W_׷Ph,5!���!����.��Я9�g���mL����i�BE��^^��`�?\{^?3���	�Y�;��֋O�i���!�o���tNo)�XJmu UւOx���֢�Gr�{�g�:s�kM���K=�0?B���׹��~�A�����Ϝ#���@Љݐ���H�Z�i�(�oPa������N�u^^�u�����r���T-�z yh wg�i4�S�3���g�J�3��n}���1��H͠��8gy�q���B�4y)�Y3����g8�=�O)���j�y��{tK�.݌���l�uy�{�FP��O7:S��p�q���"�Վab�h�J�O}�:�刟�T�,��U��Ǹ�7R.��}�dCj�,
7s%�I��Ւ�n�檷#dSQk�jl hͰ�Hu�9��o�p���7ɱ��yO��)�/	����p����&Eyz�b���������9��E��$�g��,z^p�"s�BӼך�$��54���}�ā.�s&�(�
�|�n�P�M��G��m7ǱF! \�LL��N���m��������G��,܅�$���^!q/#iɊ���R�<���[-����MH^:����8(hw]�]A�סb}���Ne��K.�%׋'o�R0d���~�s�u��,�sFL�w1j�.K2�y�*�Q�4��B�ג�\g�r�4h9��2܆k�5�G8ƃ��1��u0j� 	S�w�)��}��j
��З�ayU9�6\�%&����5�]A�A�O��E������Z���W��k�DM��-qS����:���^4ω�Yʯ@V9'�$�Jw�Z{��y��8�3ʳ.+D�ړܓXS/(�Wp%�*�r#:BL���=YS.`l�A���^��π��<���u�&G�=;�t�M9g��Ҫat��:�P>��rߎ}S1�7֩��CڇR[IY���W'ϰ9f�2yd�}A��F���Ę��(I�TJ���&������z��w̙1#��fM�f�k�|��pme&t�R:zG	K�����:*���d�%��&f!�.�Κ�j3(9sC�e �T���s����������v��F�[����jt�o�{�j�<;Wj��:�u"8e)ӕb[�g,Q�Q����8��me��� igZ�uEj޻͒v�T��"��~���1|��k�'��%����f���E�ʺ|6rѤ���1��	��\b�ǎq���K����NsMٺ�\��S]��y�����>��>���XN,��uV>�%Y�yGA������fS郮��fp�ũ��*#�����]�c`4��g�Oe;�^a)����d�ٺ��u{;-Z�M���'� ��ҊU=t#��r�Y�4ԇ�Ξd{z;��;��w4�of ѭ��Q�{ʫ}|�Z�e��c���t��Ύ�b��/{
����n�{P���i��U&��>��A�c��7������[��0{�"��������G��]G��8hx��3[�,��rZ�p$�Y�wU1��5��W�t�"�YW*I.����|�)��Y���'e�n�!;���5���s�C��O��]>��1�E�t-����
��m	�p�o�*���.���_���o���	��hڃcv�eo^�wM�w�cb�����U<���.�	}��:0�cܳ�ëMxR��|�/B��^�JY{��nb��9��s7Az��)`��Qw'%wI�J�8�ܬ�i�W��ڜt#A������﫟-y���/�bk�P,ow�b��p��T�u�0Ã���S�0�/�r��).N��3yT��ѵk��Aȃ���:jTY0�b����m&y���=��L�g|��=l�Q[]��ŜڂóY�e(��&:��V�b�5tP�Wg�f+W����m�nU��j�ɪ]���x��}ʯw��L�W�>���	��|)����]�̩m�9�kW1ʰ��6�£�4Ʒ&�)��Q�}����8uǉ� ���"�\�l:�,���%��2���uZw+
N�c�s��rZ��y��A^�ZT��+�w�_(\�w�(�����`�D�
�-��+�x$�߻V�9X�ls+��Y�R�i;��ֽo��Uy��P��.h&������ػ�NrՈgH3��4+�7�Tf\���[Z�)���븩�[�g�sT���v���gM��ʻS_�@E���8�/rXܚ!�Z�8橌�����d�������Z���iiF��jY�e�����=2;��d�E����k��O2޹���	�K��M�J��K<m�b�Si�	�},�������y<��������#�O����O�W!��
�MN�q�k�g&�J�W]��Ev�+7�4�f���J�����qZ�m��V��uC5-�P����;U�0��Yh���KWzA ��S\�;�f:#�K�z�N�BC�l��e����N0Ua�s�d�c�7Z�fA����w�r���o\��;����!�X�����)�αɺ�<B8 �vne4q �]nN��u�bD�Xr������ϝFMH�����0vQ�)�S��P��'D7�/x���-0��s�7Lތ�mN̗-�i�bd�b[
�}�Qut��(ʺ;k}ow��ިk��*�46�e�W��_@��P�()����� ݧm�b<+���XR�hmS�;k��θ��SmK<4��#6�-��㋖Դ�P9�
r�r�U�t��Wu��fj�o]��6�ˌvTū���"7ΗL|J����e�z���u(@UCՇ�uu��!J褡܀��I��U���GGb���{Yx�R�Ӕ�8���T�:�6����!�
�{vV�{j��i�Ζ��b��zH��:K�34�Z��
���jK�c:㷏+m��� �+�S�$S:��d>�U���{�aC2�l�u�,��%�kxM�dS7�wl����\��т�)�JSB��v�B����ش��֡ھ�+)hRa����(�����XFY� |���-�Z\���^mi���9e���%�HE��\6���D�S�� ��ޔ-��mm�_	� i���|L]��Gq��ƛ��pcf^��)NK�xٕ$�Hچ[,�B�Ai{���i��3�,���ҡwn����s��+��z��0�%D�郆뺷\���BZNx{U��;�E�$U^�������4��u���k�W"���r�����!κ�m���<�OD�$��d��\�<����Vj��b$����8[��QDDNR��
i���j-%T�t���u�	�gK,�7=���܋,6瞗M+'3�=MݺT\�f�j�m�V^��g��JI���*<�Q��Wsr���4H"Vg9Tt�9�Q�;��%sna�ՙ�fvbV�T�u��Qw2��k���X�TQ�`j�EX���b��֑�B�q:�TE*u4����r!ʨ�,�VjT�Z(e�UHq2�3T2L��H�r9��F��i&�m)�v��R���U�+K���K������.����KI!BSTXGH�R"�Q �� i#�uۛb�q���V�ΰ�J��F8h�\�X�:�\���v�����cE֡X��W���2�Nl����UWթ���OSL:%��G}���k���V�(W
���0o
�|*b�8�rr��"+�*r���d�f�;s9�km��{~QZ�mDr�R����B�jsK�#����������u�q9�ٰ�H���8��8'm�<J�Ε��<���եS��2_�A�zV����S7�m��E1��%oAbX��S'C�lO*���E��Χ\r
�Jm���le��� �t��ʼ)֚�]�oV�y���wUytw�pH�JlY]��Wj��"�Np���H�_J"�s!.��u�w�
�5���	�I�b&X�x�3��Ii�}��&��-�
�CPy%��=�B0!k5rmT9�!ʊ���4d�yU��ޣ���n�2̈́�Rj�B�.�>��	T\N�	T���MD�	�����y�tp�؄1�,� ��h���\2u؟Q�"urY%A�Y=wV�9W���q��A̜<�W�a�C"s��6�Tm�x�8d�w�4C��`
�z��{$\�l�L�9�
����ta8T���s2�DE�kM1Ջ�K᛻F�6lTV��Ӻ��q�}Mj���g/�n*��������ם�3��H�,�GdlV����w}k.T��喦h8e����2.��4��Bt�ZV�QY�A��}��}�^"V��
 �X���;����3���	̥{K�&|S�#Qw2�V���R���nr�;��v��,���`*�;@�{�*��p�Ɠ�}�*�zʍ�&0��Ǭ�|�#�.�A8/2(�u�)�JqrB�8���(���1����L�R�n-R:�7P��Lh�.���/�ϻɍ�Z��U=�q�$�W�W���P�E��j-�gA|���w��gN�ֵ��׍2���f+ڮ]��� �g��߱��ݟI:�!
4�SX���s�Nn��S-�����Fk�[��r��gK9b*}r�Ь4�,I_u�y�䰒ϩ��>��P�W)�gU���Ň̺�0���[���P�hT
V�2ڰt���o�RC��\F� ���S�3@vT.!�75�[�~.��F���q�ܴ���{M�ΡƀJyu��S��%���֢�(�^�vL�N\z8N�,�N��.މ�&����O��mg�}s���	r���!9F!Č���ь��M7��G�K:΃�%���ex�&�.Z�n}�%�v�C��e��,(ݼi��."���)9T��ݡN14�h鵵w���V�'�݉�B�k%��n�Z���|�{�&�Q��Z�W)�+T�г��S�):��߼ ����LS��ME�#�̞:n9�z���r���V܅h&�܁�
'�,���یM�����ܞ�{���=^X�#:�h�F���a7<��Y��K�g�]B$!�:�m�@��u��>9����¡5�j�c>���7��|��7C�C�<��N˖I�\���,�DZ���w��~��Y��O��F����>ׁ�,u���Dd�>mTT�������ή���Y�|�N?��M��`�n��/�!��*Ʒ�k�C����%�3c̔Ío;mu�"����[O&Le9�S�]j-P�	p@�]�Y��f���
�u�����qt�UD��{W9.q�gcQv�5���m䠾�Ep�<Nc7��Hk��E��eTKM�3��tg)�ؘKOt7)�de�q
c��N�Щ���c˩�4��a����5�N꙾J�>��ʱEX�֗X��1Z���K�z�#_F�+��vl�.W4�_ᨭ���� �s꣢�u�Ï2��Нu2P0,�kO]O�� P����W�b��"(�M�㠪9�ٜ�E��,e�%&�s�d;�H���u�]�!�h_4�#k]&�r�'���[�ev[X��N:�l#4o�����ڏ�S��D�2u	��Ы�{�/�tfM�Tz������������������wv��"����/�U������K�`�	h�����Ur��O���>~D#*��y�ͳ�Y�j�@Zi��׏>ۣOJ�E]>DtW �
�F�eR��t7��s�����˻�0�y�����,�W��;QMzL��K$̢��2y *�����ɿ`�o`+��;xF��"��{f�V��61EK
3V���_v$K�A�'�w�-tΞ�N�ft��P#���q_h�_=�	�t.�z�9өU�܀�e����Q��c��<���js;��S}1Q*~���)��Lq���
v��'Cjӹ���S�9o�~���K,���+��l����@�x�Q�@'����
8�<+��t�J{��F�}LS�1\'��.O�A�q��R���fDt`�㶆n�b/5���,�hv�Ы��h�Ћ���C�1�4N'(��-��N��������6���望BuhE�_�*g$�q�w:�5�L���p���3��^.'�b���0*�K�-�{�giE�	��q�\���]}sC��H�LU��1��(�"J����q������̀�9]:Xw�$QHQ;t]Z;�K�N��Z��TQ���et؎R��"R�e`�bU��L#����P5�9d�WP�p2�0�X��7�P��_}�W��V+��Sûx>�kF��S�s�\L3�ze�C��jv܊+���tku*�J����j�W�GO1���]����k@�r���ǯ�|.ϧ��s��]E`xx'�յ}�,�~��n�k����̯�냝��gǾ:���K���|C��хң��k�Q�6�q���g�����h܊�6��L�XLt��,�y�!Z�::�\e�ǫ�E�=�()��b��
oP�TU� �!�jAQ����938�_5LI7��՛}P9�ݚ=x����Y9�kl:�/J�ClW��4`��A���qZ�=~��q�Ҏ,����5K�zz����M��C��w2�;��1W]''(�q��E$_-�p+�y�]�m�e���G�:� eO5�;j�5���I�pZ^�$�*�Q�I�wL�3���뎌މ�c)�r O'H�#ʼ)֚�=}��ß>k"���"P�'FÌz	�8��&p�=݇��i#�]#tO(�"��[!y���w?��+�xVq���(4ɛڤ^���(���:��8�x^�(���Z�\�[	����t��b�*=�J�`n�:����;��%����D��2��s $�'�i�+6������=kv�0Y���sϦ������Nݞ��L���Rn�p�1���`�`�WX�=�x =UV��{x�]�!�����	��$sr�s-A�t`S�9��5rmT9��<�60��H��*��6��d���<oɾ�Մ�r]^s�9�\N�	T��0ѓm��V�]��%I��9E��mK�V	s�}�%��v�N����8�<�C�w�x+���i��z@{qu����T)��Fs�g|�MJ�mǚd�{�y�<Vkj+3!��Ι���ť��0Ym}Z�[D��z��W�.�u9�H�]̻T�.�<!Wռ�]YB�ǭ!�ZW�5¸*�k��?v�g�.�������-~�w�.I/P�H�{���1D�~�M�U��5���%���P�V؅.�ke
��`cE&s2���v�"ڋ��;&^�;uڸs��;S�;���'��cMU�@� ��������8 �ᓈ}��O�8��٤�e�\�Z����x�s-���>�UP��ۈ���]77��Ǎ����=��}e�����3
FS�_X:ꏪ�`N [�Om��ݙs��"�m�c��Ѿh2T�p\H$�n�{��s쭿��b���?D[Z�?��|зR�8����%��SA]��5�!���x,�S��'+2�hY��K525��i�fn���S|p�.��!J��s,t���J9�5��#�,���y:�j�b��s�Ö�U"�_���꯾ü�qc�]���R 1PL_�}u��
�=�T:����~�˺����e����-���?8mH�T�����<U$4�Ie��$=��6��g�ֆ�����c#x�y%n�{
��v�/������{�>v��f��`��m:D� %��;�W�Gr�ɜh�E5t��r��c����=�|%���x�?AŴ�>����B'vBr�C���Bݎz���,��������1��N����@��g,s��n������q���e\R��oWb��p�+Շ��E;�����8g�ϫ����B�4y)�ɟuu>T���do��ne��������Ô�7��|�5�\:��!�r�8b�b+�W�}Z�nW(�r#aC��>���>���o�c�a4�)��٨�D�;-��KWkO]e����nf{��چ����1:8�}��kS�_Kfl��j��a�+K�xxt��J8s�U�=^p��ɓ@9�R1u��C%�5���g� ;Vr��O ��ti%Nhn�+�:c��O_)��T��	]����z�ҝ5q��A��Ħ,�x�b�L�ю�(77�߯�v�p|�ĭw�u��-��rY�4.H��1C����2�KۦӜ:Wiz�V����bWS�"'�{���36�^�:����C��g��h��(ok�#���d��2u�E+�.K0�=~�Z3}��[���Y:wB�/}��4�{�ĝ��܆hr����s�hW�D�C�g�G�r��+hY���2��O�r9�m��6nFD6�Y��0k�plu@m*=}�^�ӤTɕO'���e7�
V˂�hE�
w*��� �̰lD4�s+ a�eQa���q���L{��q�q.|��]ާ��/U���ȓH�<�%��m�5WR��]��FV��뺪Y���kW(��!��`��[Ν{�W�Z�zY!G�3\bZ׉}[A���oD~rܛ��,DDb�B?v�g�1�<n��9��
_H2v�t�5O;e4f{ʪ��j���A����;}W�I�Az�߹���3��+���3{>/��\�.�e7i'�}�L?�WM�Ij�'S"������M+>����x�Fn�Ko�~O����9*L��+�B?w@�N�9���@��y;��"�����N��j����v�с���������3{{��I��)����+$�i��I����(Qܦ��Q���7w!�=8��*��1�(�V��+\��]�O`L*�O�DZ9��5�6싍YU�\_MWe���� �m��2�Y��_;`̕�M%q= &jͣ�e7�:ce*���o;���{�f�S$�y/����9k*���9��ٴv5�=�n�:�L;g����Ի-kG�6j�.Cm�t:��(����5� U�"�̞�|����H�Τ��o>��x�'uk\*�M���Z�Mj���8Hu,u��ʳ�1��Y�/����T�.p��ϰu�<�C�Nt�n��s��b �ӵ��W����R�����5
��	��b�a᳑�]i�}�Z��O�Nf�n�~�����X�W��o���f2r�G�GԝY�g�}=z���v�?_u�eH�}n���҄�P�qGxv�F)v��x/�������s9n<f*\<��}aBu������S�x߳�������hnqCx~��8쾚�	�3���O(���j��Y+b<+K�qĸ�u��Kٳs̪Q.����4�g؟��[ QƧŊ�`�Y��QNﶵ+)��������A��rb�i�A����¹�ػ�v䡜�pN�a�V��\��V�x��ˠ�n!\�fMum�|��������5�'x,��w�j��n�,�`J�.�܍p��TS��Ƨc�X�Kpt�;��D�
�&�Z;�H������o�u�׮u˄�Ω�3is�XJ�ɷ
�\Mˣ�4$�8$�u��V�Kd��v&�Ƣh��E�;g*�-1����n!HJ�?A��%�q�5�qN�Pn4�M2��v5ct��eapo"%�>�]ٟlܸj#�u�)k��ҹ�`�u�!+����g�ǹ׶��Y-�y/���>T�QS�/"v��˛7U|�7��T�T�����l�`��] [�y�!���
=b^�;m�Bu�#T+��s��yu�z�uk\*��q�!���j�n�-q�C�[�i9U��'p��ϻ>�E�/w*�)�kI��~~�N��{}еu�=��s�y̵����U	8��&���}Kl,���/��)�#gڵi�F���{���-X1���os]�p��v�2� ��f�Q���@�$Aܨ��'E��R�4;�p�`Ŋ����7�S%�sJ��̥�0�	�̚�Y�Ȥ���ߣ�(lN����:�+����,��\�1�����{��yn��kW;"ea�t�ʷ(>��c_ީ�Y� �1�}�m��հ���>�-��NK�"�e:%s�f����;+��tޮ�6�n���g��а�U�P ��\���;�H�vt^f�Y5���9\���M���ѵ�*Ay$��1��h@m���/wtV�򦽳æ]3	G� t.�,�Sӽ�5]]#sJ)X�jn�'W)�%�MlTݚM_��~O�QV���^��K�Ih��g�����],�v(�I�a���W�+�'�@зo ��I���@��\o��)�=;x��f�[���W'�`U�u,3m�>�UfTo�=oC���*�
�i�h4�M$+[Ws$G���X��A�8�Z�٬�ԅL}lj��v���qe�p�;���V{3�.4��]�/iO`i��
�]"���nAj7F�;�)qz�e֘4d�Ye��!��e��9�|��@�x�;�,T�ot륐�8���L�R�+(�]{9ف�U��=PX�O@meK�S4���W�G�)��9er�,�}��igV9��6��V��Åa߁�IC17-+�m:�Uۀ�]���qc�%5*�u*��
��^��q�^�f���3Iu_J;�۴<�y�m���4=	����{�K}��nd�H�R�����u�v?� j�t`�S���ɛ�'jaw;���5����tF��E.:��D���/Z�^�t6k|���ީ��5}�� u��R���2��9$�=��Tq�/�΍��e2�-���׵tq<�ݨ^� X<�8�=�@^�rgH�ζcz��:��wju۫i[¥;
�Uw��^�>�H^���
���X��]N$��N�Ⱥ�����uLKWE�ݕסc�`uȥj���q2�<X[��Ӱ����6�S�Qm�}|la�l�Ƹ����ŀ97q�O�]t�F��ʷ9�I��]�+���"�̓7gB�EdY�O����xA�	�f�����U�e�i�D�ѵM�l�v��4��+���<�`#��,� �#�N��߯���u������K�44U�0r���f�7��&i�u{qɬ]����ٳf����@�Y�s+;�a$#����a����Ӻ�4���z��7{�<��j�;�6M��0��O�����]k�����6
g���CkVlvFtEs�ӻBb�O.q��<V΀٬�rեǞ�kU�{/�aZ��붆9��H�M��@B�z�#u�ݥ�ץ��Grg�cfa,u�;�����]8!A�E���X'Ū��s���+8�w��I����zf�Uքh�(Dr�,���%�Q�JJ���-E�a]SNfZ�+Q+�R�r"�PCY��%�Aq2��R*�wt�KԐ�"�X%mAZu,S(��ʺ�d�B�T�iȥH,S�%X���I�9�&Y�XdV(�V��ꤪ�e�E�:R�)R`�r5Q%2J��D�K2���J*�sH�:j�GB�db��2.p.hkIV�$K%�g2ډ��*���BI�4��!�f�L��ҳ"�*:,��h�26�č��	��B$�U+(��EfI�2Y�JB��aTIN��
YUHY�*�T#N�b"��a�����-*����"*)"Շ,�d)��4�֡��T��kD´()dPjW䦹�I�3*�ʑB*���G��Wﯿ~G�<G��\j�ns�()s�8�cS{���	n����F� �L�8�i�����k�v�5��RbjĽ��UU_Z�R�tҌ����-k6:�sj��Y�E���9Q�����9t��w��mQ��i��e���\�n��c��T�ʳ)8�TӍ�x/��#&��e���҆�u�be��e��m��:�1ִ{3h�za��?ks6�}�s�*U[u�K>�v�477������u��Nי|K+(�Wa������H*���6���G�>���;E㊞�yM�nSa�^Y�ܨݶ��NƲr (,����.���n���+�e�)�Ն�\b��}�\c+��sr`o��\�jqwwa��d��t]6ə���W3�V�w�o_���	tMʨ?A�Vv����˛�5���Rg���\���Y/9���8��:b��M�eL�8k��>*��ʙ�k:�]��+\g�i)l�ȗ�o�;�X&�����xD�=��+T[MT�P�]�!����s՛��[�3w����hw���xGJз/�[�6iT�Zs��BF�;n�:���u!�J�I�dU�F�.G�L��\I��M�"8�U�s�-���Y�2��
q�̊�[� x 9׻����_c=%s��W��%7�u�]\&̻���5�qH�_���K��k�2�NZʱ=�[9�����b�����3�>�VO���k�f�a�YL��[n9��v$Ӗ�ŵ~3~Z�?-�اi�o��U�6_-ntr9C�É;9����7��Tj���]D�7;��synAɶw��1xo�ʞ��^��ǅS9�ka�{�P^�9��;�f�vj1���9:�V.ɣӧ��^B�|�|������������Ę�v���ۀ�QF��rT������;�٥Az�v�V.��o'�)3��>g�E۾��!�L�%�O�x>�q��M��
�J���1�<@�Z�
.��1��iL��.�r��Wւ�M-��%T��U�h�8���ͽ�9��9r�����>+�F���n���̗�;GRZd��V������l�1;ɟmy����'��*�X���;�Q@�o���B������'2�p�@��M)ۗ�- MY<�2�s�����cag4363�WYn�!C}iȊ�H3���}���mdra�n���,��6\��9��c����<��yK��2w\ɘ��t}Mn�[�nC��^��.����I���q�x����"�+�X�i?8�7�i'[ƮV�������Z�C��A��9��g�>�ɼ.�˔�ӷ���2*m�V�2s�	TK�K�8"�P����4�nj{�4�qˎ�)�NUUOS �ٖ݉r�G�A���¼������C�o:����I/rmy��L��.�fZ�^9j�aR����NTΘ���	K.�f�p�M�\��[7V�r-��@�bh����Vd����ۄq�osG�mF}]���_r�T�T���ީ�=൜��hY��s
=��O9%�N�_�|m�w���ǟL�.p辱�-.�װ��ˆ�bes�SD���.u�M�a�5y���u����8Ѳ��WQ���brd�p���VǢ� �>�[�]I�J��;��If=2�]h���=�:�AOo��' u�.�y"�/`˛���.tet�6�Jd���3�6<����&'�S	n%xU�d �c� ѧ�3��z�L�ZE����[�3=g��G��G�R׆�V����5X���G�Z��EG���ʍ���X�O��OF�s4�g%��|Ŧ4U�����X�3�2��>#����Zk=�Z��롫�s�S�M83�\D�(�砢ܺOL-i�yE�[/�D:�pQޞ8�-�7��-uLچ�'���Cs�g��/�X1���=I��[㉹:�&m�5!���q�
իYC{���p��M>�
U=+�)
í�J�6�a.��{�FOwP���^D���!�CX4��^�_w�hm�+4���+��5�h(I�pIb�㐭��p�dv�{\��y�j-�����)�w��BQ���9��M`٢)������k�B&+��j3T'�7�+��M��:b��n&�����23}4�Q8��q�zY*�bZ�n�낋Y-�u��S��9����QR^�	�>���)m�< Ψ�ދGO#��Y+�t�W;�����A���&K�ږ:f����HY���&K�	�(C+v�-��@�r���햃�(��jۢZ�<-u=M-��pLf��g�.�RM9۽qr�;mI�)a�؝7���}��_m��e�<Uno�VT@ԫ)��%;惶�b{��@�1׺��Jz�e������3:"Qc� ��j<�]�μ���d�=m���¨��W|FNo^��W8Y�f:���Oy���1Wk�^H���9?-]�E��g�.�"�ø\����X;���F�)d��Fu*�,Of���S�g���K��R۫���Ɩ�%�Y:�,�sq��M)K�����/S�	n���*N�1x��4T��q��nW��#=��V�Y=֯"g���ز�,�w�^k����F\� a���#��Z�V[���}���g�8���#vY\�i��VUq})\�#�����	��k478�z�6^拔�ɋ�_b�ou�Y9b7���6�?�U�T�ytd�J�Ɔ����`��{��v���u�(�;O��|b��3�̬�I���e�&
x��K�+��k�'��qw�:�tt9�)��Bb;O$Cy+��.��۽�pf�_u��P���X�U1-�o���jVzA4a���� o�S*�r91wktI�gVq0�
��,�9H��i��)3�.W�+��f����pѪ�<�`��C�b������꯾��ݾ���ۺ��ܔG�+�w�s>q&�{l���P"I`�
��Zfi=g�ʅJv��7�S4~��܂���3N7;p�+��G�n�B�J&�z��
��. csz{�q�\�σiC�z��nu�hW�%4�g��rks:�{����"����q���Y-�y/��y���)�?�gOj#k�}&�G�t�@\�ͣՐJvʞ�����_Hx�i�����V���sn$���7�H
*z%87�v��Y}YJ�"��K��5([�6)2M�"���sW\�I��58����=��'H�}QZz�3��V�d^������?I�f��{�����s:z_�Y�M+��s�;�qzR�y�ou��ȯ���oAT�B�Z�lv�ϋ����8��ג��(�M*b���_rч��E|ZQ[��UO��L��_q3[�_,]ER�W�:t���:g�:���dn�+㵎�$���)nhP�
N{m�S;�z��]\�*s�)���Z�;�vJ˚Md�E�G�H��67�ge��	|��5��(��\V%�=�,ږ�1:I��;1A��&�ޛw�B�8}DG�m�%<�X�Gv�gv���U���	ʌq|���&j�0t��q-�^���A��UѶYY�Dt�s�� �܇y<W�1ݕ��iԯu_ejj�Ν��Ws�]^3�׵�k�U�o��g���j>X�贈����0��b�Z�;2v�&̊a��m�;O���~�3�)������E�Tt��Wz7J���*��M�s��#\.������ܔ�zfv)�<N�%Ud�`�_��]a۷�pz^5˜o_���3*�=���y_V*Ҫ��M�S��}@��zKX~C��A�
��7u��1�R��L���Ӛe�;q��BUDJ�Ȁ�M�z�Jޝ��@U�%ZJ<�v��ƞ�ݛM�\{|3�.:uZ��y�cI��`�3�l%̼�O*ֲzz�H��ٗ�/u��G%x��N�Ea�̼e�L�/U�VZ�޽fiUˤ;(�v���C+����j֐8P ��8�7+8�K����m@@���D��DyQ�g\r�=1���P��q���_'�'y�A��`y�V轸4�/��N���ޭ1�u�������	&���}X��|�c�Mu%��W"����Ow2���C�!�Q��Ù3��::6�W�5-�~�S��f��噼��^,����
�C_�r��7�������.{J��9�b�\�sM���}�V�
�qs�D��7W�<�lɊ�V14��ãz<�����wD0������=�k��~�4�7Nz�s�H^7W��8�E,j���������ݸ��=�`+y?T7xtv�oN/o����}}��ܯ���M�:��ۂ�v�,��r���(�����x[n1kSW���oLN�6Qnq�}��vB�Y�6��'Wِ�h��{iy���s_z�ě�nLվ�+�#����M��쾚� *w�2��aG��=Z��2����x�$MV�a�o�\N��ɶ����l��r�W�X���t\ɕ,����%��9^D������m:��kz�����Vv�(1{�"�ٙ�u�/�&��9���:-.W�ӗ���hAdp�)}4FE.�g)�����*ˋUD����s���GIc�+n�`i���%ר5m�
��g-�]�i[� ��8��;[����҃0q��c�G��Y/RE��7P���gn>T��ܚ?3A	I�JH��#m-l��(�դҩ�ח�=������q�q��ۤ2���o>��]r�G�H�9�1M�:��o�2�J^s[�e79�銈.=��N��S�!f.�݂)���c���~A���z�-dD�e���Jj��|jgT< �7��5���ۼ�t/}+*q��v�&���!�ue'/%�׮�d��^����{�t^|��}R\K��.�Ͳ����O[j�Fj�z�3�÷�P������%�؜]w��/$�?9T���6��(�3F���t�S}�%��E��?-��s ��-�N#N��oWe�Im��c�,�s;��5q�e�*��a:-k6:�sj��g	�g�Ꭶ��+o��ι�+:��W:;���g����H�����G�q���7/1�sr̒SV�X�/.�[��,Ks �¹�ܚ>R�������g(֘��G�oƓ#s\]	n�e������q��-s�B�e<�ыh��\"���HF�@I�s�nZ���M�)���V�/�S�������x�ox(�����U�o*��;~�����ȚP�D�L�aYnq�}�B��\��".��u�>D�������J7�yQ#������BY<�f����v3k%цlpkC�d��wٶ�p,��8߀�g�9�^P��E2:�{��5���/N�~{9M��cp>���9��9���'!p@�W֓��;Sz��{ْYt�bjj�?�����}���O�����7&����}P�YF6kr𓕫+B�Iuk?C�j�6w
֎�8޸��n%)?e�7(��p�ù�S���U	b�E{Q�%��\�σidD���	�N78eE�N�7�7�2�N��3|�	���K�Ϻ�}��%�w�)��-�{��s���a�ˤ�
z���y\8v�Ar�$%s��W���%;�T�JVfav[6�]L=�e�-�t:��{x���KT{q;sڽU"���e�r��3������*g���1�� ���ɱ�t�ۉ;;��5Ԯ�;�}�;���$�(s��V�� n���0(Ӏ�+1y�%��������y��P�ЅW�h�rm�ڹ�(�ىJ�:�r<��Յl[r+���Q�3]�X�����q}�����Ŏ�zF��[U��7�[F��f�QԂ���v��%A@[�	5WC�9�m�f�k���"v�����Lܾ��B�Y 6S�v�Ԧ3gi*��X*a���uHƎd��D/.]�V:�.��ɷ*hڂ,��(���oML=/G��䯱,��Ӹ�j�K���L��^��"T��7�& �<�Kt��7Tԩ)t�^o;:QB�#�(�|.��ܳ*�]�B8/�'��/2��8�ڙX�z(sept)9�8���4+Y�#�(��NY5��7Qv���B��X�"N��q�p�	M�RT0��f��i�P)�@�Xi����jҺy���oK�B��f(���J�����x��y���⺂�;�s�a��<%���URX�ֿ�4��� ��Sm�V	n��V�s@�X�޺ݝ���%�o�~�������H�_Ne9(5��n-Y�d���Y�ش*t֛���|IHW��`�4��R�9��*LYWƕ���Y�������-"U����Y�ܳY��6a/mPf�X��#ȳoN�h6$��m	q�ƺ�,��R�x�
�t��:�u;R-�-^T��:BR�0-Y]��S�'8�غ��Z����e=��a��\��s�}�Q��T'p��N��=����g#l�t�1�O)��R���.:�K�]ۭ���e �f����N���m����rBR�{ja��K�v*�"c�i��u��{�,�z��Jԃ�R�P�|�A��n��Ϙ���@:JR���z{�^�у�nlv��ew)Ã.���$���+�������q�X��s�̀5����n�0N$�1\�G4�C]�V�ȳ����lh"��}�@�R�Z��9��(C-w ��ݘVl�4��x��Lq#LP^k�$S9)�m�5�:ţ��<U2��R����W��p��Sf'A�]���g� �Z�V$ι�����V��k�V�:����RIf�G\��n-囤��u�^	PЈgl����L�5����W�_�%N����Y���%\�I��N��"L�,�}ă�Z��g��t��'E��R����*p����;-������|�� _N��ƻB>�Z�7!�����q����6���+����El��ܵuũZ8��U��j�Ò�q^Kr4��n�p�k`��r�T0���S��<�Km����bk\fT�ne��;�H�K5�vPH�E2��ۻ<�;��9�	jZ�DXf�E�-�R���̘8�W.6xl�Dk(�d�5w!���YsM��*B ��5@Q'0�@U����8Ykj#N�W.kId�����yVF�uZ��$Y2����R��)19���1V!��(m.j��hb�Id�)AJ���PŦCC��a�s�\P����DXE���t�Z�ʥQU*��й@R��,(��Ύ�P�j(R"�P��$��Wq���9Z�ĵi*ȮQ2/t��J�Ι�"ehQr�D*�E"��\�(��Q��',���T�\���� ��eVQ@Qp��D�h��҈�+2H�D')�f��V��4Y�"N��J���2���E
��*��8�AL�g.PPP\Ԛ����E|��_���/�O\��7u�y�6��LWsk��H7';k#���l&�������N(�m�[˚��C7���W�[�&�n;�����v�m]b.Bj5��M}�6��Cϐl]�O�ZJj�L��c��j�7�_ܯ$��˜:8��;�_}�Z�:��c�����!�xR�eZ��b��|m���}�x�g!s-3C��6���*_U���q׹: ��Ww)�xݹ
)� c���.��臍Ze�zp*���^�EV�W�c�82� �Ƿ���о��T'���|Jeg��g�����>�����ݽ���Ծ)��Dy�9��yZ�]^�@����H';{U��w\�[����;=���U��8��-pVu�j����تx�F��ݧ��Α��8o&�t��}P{��3טU=�!յ�g�i[��꽺4���U���p�(��!4��L��/t��5׬��n�=靠~%��	,]a�7��OKƹG8�p�2u�7�vFJw�XD��
�j:�l1�|o����TC�������� ����__P�Km�iН$��h؂{���僵������I"��/z�j���{�DO:��3��&t��������+��8�(���Y�q\B��<�>����n�3����7ݰ@��o�ku7�jd_�$Yx�'$�e�y,Go���ӻ/�nv�!P��	o�'�����Q�"M�л��(��k���5�K�E����<��M�[��=y%+4'�f&��5*z�-��N���E2��p�W���]\&̼��^,��AS� ��v�1�Jy]�.�f�-��Z}Y��\�l�ZIȶ�sW�şd�~{��S���S�/�iM�r�}�m�do.�V�wW�-p��c��fv��oQzs��؇pM|�����lS��6�;����<���O�����q��Ա�v��wP�s�i���.5N��wNFߵо�۝�}}�ުS|�Q9�*�Y#1�R�5��D5cn?f��As">wC��m�����6�͇��p�>�;�%Į��ˌ�E�u�S=�uF<��<�����*���4�c�e��Ru�8>��N"Ю����+�P��r~���+^@@�zS�2�VgS$�.���ӟ��+�p�Y%d�&vU�����L�\����؝C'T�vuZ��j72ޡO�k�#N��l/���w/5L���BT�$��Y��az������Z�Jc���|m�ɥdN�q���Qns�i�+=�Fv�u
3,�1��y�Y*�v��&㮕u(J5�Q���Pަ�'e���	^���B�E��Stz�!�k�X$�q`y�L�&L��a����V�].i�U5���R¡���Ѷ������'`d� � ^�����ݾ�Ksb�V�՗�.1yZɆ�#�p��1�ۅIEIȃ�4���������N�/z�;ȉ%Y���z�Jd��c=����s���BUA���9튩���[���=��u咥�����s��Y/9���6��a�2��l\�8�$�o�"U�k�T��Q�^�i���\ZȖ̼�^)X�(�3p�y]��4��8��VЇ�UHJ�{(>uq��VA)�4�f����y_b�w�o�k��K}L�`��-g�"�i�q��冻�_'��n�Ǥ�k�&&��T�ϟe�`8󚮲c=���"4����i�� R�h]�(,�g*��CޅS�������3:ᩮ��	��M�e�jt��)��q��R�N��yS�k�o����bZ�O�6.)os�VB�RC��;U�٥`P0ޣ�~�*��s���wqq��cT;�R��o��v��^H��?E=��Zԅ�o���>饚���E��3�B�SF���1�1�^,\읾I�ǲ��ۅeOf�}�Y�U>i�e3amW~Ѧ������o�\nN�zjL���EMׁ��t����C�[.+�;�1�c�r��K�=�'���3՚$T^B+h�����2!Yns�m�����b��o:�kS������,�g`ۋ�Ǣ�
m-����T������UƒPKQ�śU�t�je�)k�C��k��ε3�\I[A�G(.�V�ζ���ӻ���2]HLqLs�9{��NWǨ�=8yܙ�:z-ߒ����-�;�ZV���\rO��5ٮ\F2���I���z:��٘ua��nx��T��i[����^��.�y횿�gsⵣ�s����m�IT]���+��Lm����p˔󹣊��xze��� ��]�+⮰�Iv$	"���l��J��\���n�޲q^�;ygg;V,ct��1j.	�Q;�:/����9����rկJi{�,�s���SҘ�bG}c���2�vN�Cmk�T��DE±&�x����5H�����q�̜���j}Ӹ��Lj�����M�4E1(�D�U="}W�Z/��?.3�SJ��1f��:��S[d�L��U��M��S{~�&�Z�B/c����;܎��'�o��+����dG��%���-�t:����� �AڊvANz����_��R��K<�P�e�uq�9	��.��	���Q8��=���&a=�s�N����zm־���}|�$�p랁��yU�b%�tV�����*k�i�~��a��z��o'q�x�g8-k6:�� 6V�ʴ�o;0�������@*���p*�Q��u�� �z�5pd���z_&ǲv��G�	����+�;T�}�5����TX���1=W�2k�q�qG����:C4yj���r��������.�.�f�8��5&��Գ2��:v���U���T�O�"��|�\�hUp��$LR��w҂[�M& }}�TϠ���Ò��x�7R\κ�=���%�p�q��\iT�8v�J���[J�u�jt���`�*�������uJ,.��yմ�>�BO������Q�;��7`�����-��L����v�S=@�R֜�qJ�s��S����7J��j��;Y���p��m��i�@�=`��3]b2s��e��TL���0�evt���g7��>���O�)��R�Y\�7j�����ˠ�%������|,$�>���S*_t{MS�^�`����:��J���T~f�
��|[�q���؋1��I�e�ܥxc��] ]���ӕm|���ڽA�Ջ�n���؊�����==p�J�j%�ͦ�-�����mZ�{F3N��l�������f�*��e4��\]\Bl�ȗ�^} B�|T�*V�C�[m����g[Mp(fk���5*��z��֋�m����eHm�u�.����&�]ո���4_��(��V���9=��E�i�OnN�L;)�b�a�a�f�̧�ᝬ`�HB��O�y��> ?f�j�n�0s��j��7	uԨ @��a���oT�{&n�����w��L��N�/;�l8B�c�i���N�� �uv�Ϟ�7��f�����^�#��.G�~�*�;f6���5a��,��A��'bs\���]q;���r���_^D�Que�7�Ѷ�zfg1�@�龮��#3�;�"�N�=�r�o�����y��Z�t$�S�?C���]��Ʞ�2�j�߳h��.wl<���rbU�Ѥ��Ǫ�55������Z��r����9;��.wv����c����l��cIw��������&�5��η7��ʎ꾔:�܍$�j��VU�q})_�e}#��]:��	d�ܜP��&ٍ�]V���e5zIg
��Q��֏v˵�'�ÛKq��l�Xovi�i�bu�V����@Z������5�S&�(ʋ�Id.��a���}�Is�[wwO�ڷ!(k�5����A.��5���
��Թ�ޝvF�*���#|r![5p&��8ަ�`qˉ��ӻ2�-������w�KX���*��F�bQ��Gs�I��\~Օ�a��a�+W2V�y!�8�!�V�]G$XFp��75HV^��GANk۪ ��N��8��(JXr� ��&˷gU��q�LB��H�e�i������X����}�߸';�Obm��8��wfG6nC���eȮ�B���xJ����W�|5q�_j�>3��E���̼��Qy5;�3�u�\{P�}DEC�5!����_�h�d�4=�{گB�&��X��3���&�Y���s�cx�=�]@]�w�4^v
<\�Ϟ�M .��E�Sb�wU8Z�U�61׺�:F �tWe���F<ș��36�����J�O��[���m��+�r8ts��:�Ur���Ů�r�"�a"<���W_N�I�~���^юg��-x��=N�Z͎�����|--���}z�QӅ��U�ōu;��V^��S��Q_n2�U�]�)���D��λ�����V3v�iN텕ʺ;}�4�����c"��t�H��ΰ�.	]�3��jH���;ke��*K}��eH�g�eV� J����V�˽n��ү^�x�Cg�n7QM�[�m���� #����Z�f�*X=/]]\9ۚ,ս�I�F���������^4F��	��ʰT�
�&�iΞ;��N���w���b�ਰ���y�y����K
�˧ǔ��æ����f�(c����һ�!�1׷rA+W(�r�K]�9���{ҙ�]D����.��`J��d&��ɭ�u����>��kL�� _�8T�J���+kr��S���'n�-Yaۗ1#;�c����4���v'S4c�@ʉ&c�53�=BP�~A\�u���W��c\���79�&��E�N�-����U�U�EM����).���C���L�����u�1��zNHL�o>���sL���n0�Q�#��_WR/M@���{
�Es�GR1P,��wIKN%�����hA�HJ�zG�s�H�*.��]�,V&�p��k{�u��t�2���@T�����	���d]��V��{��px��������W"����$�Zn9���bJ�2�N9TM*ڝۜV�mr��Y�q/�R}��˭��w�'\�®Z��{����l��\��TW��\��1_���A�.��N��oҥ�!S}~�p2�VWu�j��y�C��E�luCՃ0ޘ�T���x't����͈�m�+�*9ǜȻ�va%��T��P�x6��C�h4��
��a����:n�Z�������bSs1wG]&����-�^��r�=�o'q�x�g!s��>�+xR����̱&E�:L h~�s>H����ETw�I��e��V�U���N��n����q�y���0y7�}5"�������ݰ�F����NWm1y��/t?���Yԕ��q{���e��w���6VGml�v�r�}��ɐu])�l�7]e�ݣF8�p�'[���}�9�i�Q��*#n��u���������
�s.�v9��3L7u�m���}���E��w�/7\�اfePP%q�F�A�
�Z��M�G8ks\.h��i��<U�媯��긛�_2k�}K�%��úo��{7���f�NWn�JӴn��|�z�ۈ���1�}�:����L�fq��O��:�]�x:�J�{S�ns����I�~�$W��[�{f.=Jٝ��H���n;�t��M]� Tӡ���r�Uܣ�X���f��C�EJ��Q]Yj�����B��g�U���r
��؝��-7���9�hDň&�XD�5۽n�q�s���	�p���p���]ԛS����"Y��i_7A��N�ͺ'�A�2v< �*�5U��
x'^��K�4ۮ�M�ڲ���̹,��r���S�e�����)�;@/�2��@��q��wM��%�����i+ۋ��[0�Bs]7jT3q�t	���׎]���U�rY�ע�.�Z�n�Lf&���ЗK{��(���`Ż� ˬ�N�	b�$��R<6�ٸ_�"Ϊ�Ohq���զ�-���Z4��l�	hyPpa�����MA�z��Х�Ȑ�����^�1>G"9\�Ucx��L�r�ő��M��]�G�y���|h�U���B��B�V�[Ʀ`����i��z�N����]k�����&j��W׼G>��>@�?^޼ǊU��i�fĆ�NrvF\ �//O��벣�����q�X�+�
�����Nޒb�xՅe\I0_Z˚��޼��{�ޕ�.Ηfv����W��luX�{��#r���N��^@,ͺ5w�v4�[B�����h�m�����k����yn��*ū�,�M����j0��oi��������X���,�8f�}�aD8��ޫw�:n����;z���Xd��"�R��Iu�3[���Ö�(��Gr���"V.���Ϣ�m�Jb��s� �Nd��I.�NFrt]�t圲��+�WI�b��u8~_]nJ�.AcG�;��H�7\�� ��F;��f�v:#�T���1��U���P�[>Ø�J�_F��x�7�/�8E��Zn�y�+��h���/V��z��I�r��;�vRM���ܨ�:�'"_U���A�o:SO�A��P���2��BS�E��A��)0��foq�N�qLΈ�ɀoS��2��É����9�C<�ґ���>�7}�=�$=�;��wD�gZ�����S+,�O��6����o��K�|	V��Y�+ ��`�^�Ͷ���Ob��qQ��,W�JdZ�&ULGu�Z�N��9Q�c�i9����9L|�s�g�s'i�Cb�c5,[�N��H�j��5�������xB��aX%���ƋRԾ��5�u2�������1ڬ�c}'��h�Nt������\�t��Ap�*b碍D���%h���}�A�����Wq���7�9�.�{��w����3�;kEp����잢����b�b��VgW�P��8�M;���	�df+�;ݬ�5��7�ﺃ2|0�D)Q��9�3�W�R-n���b֫_.��HȀk������XU������]ӝ�zЮ�#���j�]=;�p�o5(Y�Xvep�D�x�v?�9H���Ё*IIIYh�	SN��bBMPI9J�D����)�,�.Fl����.�4�TQt�$�f�%X�$fQFHR�pH�XX$�F��Ydf�4)���Y��+ZdlXG,�B(&�̢�J#!$$9BE"-8���,:BMR4��%8Q��$��dQ́je�F!&JѥUT���#Q)R��Aa���E6Pb�)��"K�$�Ւ�P�����B�U���S��!�!;�˕J�9�es+�Q9�k�P�;���ՒeUQ�j�BaT�I3:l�G8#�В#**�Vwt�.�T
���>��=��wNwd�4��DH��OVd���=F�kO�nB�y(�@�lr+���o\7�N�бB��t���ur����Xs]�O���>���p���Q/9�y�ɽ�Lo�J7I8��Ρ�˭�+�]�:�8��]�Cw��=]&̸v�8Y /gE#��1`���yv�"'�\�s��fڧl�d��r�7I' �n9��,��M>�<}�
�'�^gE���Yko�>���i�do.��x�u[����e�n���(}5��ʙ���P�WB/*�_��[S�lS�ύ���K�2+�x�GA��`�q�H���>��+���9Z��b��åZ]�'E��H%I��%�^B�zƦZ�j�߳k��0��߃ȳޟr챆y��֮��b��M7'>�QXYp�nTC�]��s㝎�������;U�k���ʮu8*$'}n� ����6M�w���y�F�Њ�V�Rv�o��2�RҮ��ݙ&�ʈ���a���z�6k�t/����Mp��2�J�y��(�o��MK�"'H7{��ڴ�	�=���u�ś)��3&�N��]N�mbH�W@���d㑍Σf+j���3/yȞ�j,o���K_=�TM�)oKn�J�S{��f�d�����jN�+{�O���k'"�t�s��b� y�}ښ45e4C���΁[����K��==ċ�n�/���÷\w��.��Y���4���HK��A��zu=}�^
<#A��{���������!^������O����@2v��.	���2\�ו�(�o_V�\�ϥc=���79ΐS+kw��r�1c9�f�haH�n84�P�k�2�K�y�l�ٴ��?3��[
�T��,�����r�e��f��h���|g��Y-�}:�c��C�u��ڡj��6�9RPT�H.�{+��R;]�����U+
���c����C�ˢط�,r�o����컸�p�Y&lOo��).Ǝ�=��Z�;��ں�Z�U���j�k<ȿ�|6�����q�����K�S%���p�G��__m�ϊvr8tq���\�eƩ{�v�@1j*g��F�s�=�_��5j֥�î�f_J� ,Nk+��!���#y�K��Aud`u���6���9� 5� ���Q,fa6��&��Q]r��ɤ8����]�!�ѹ֓�c�W���P��D��kZ�������:Ȗ6�Ut�T��$鳃8�2J����q��<4�t�'v�y
��Ls+�lu�k�x�h{Vf�{�u���N췳��V^�D�s���^B�-�þG��s!j�����Z�t����	v=����M(k'\Tbe�׳A�O�n�s>�(�$��K�o����5"���9�Y�2\Č��Gl�l�N@�R���y�^�aݝR��^6r��\v�tZ���H)�;�9��L�G��]�QJ�6�YC� ���k��Z|��' ����X�*��)�[<wJ݇�^�4�e�n���$�9�]��\c1�Gݻj_<h��oz�ݱ��vP0$�/�Iuk0횿�6t�k��i1��[�^gK�8�,�T��|鸎��8�.d��wb��m#�6�q�{�o���q˺o���1HJ7WReZ�A�f�������5}�C�[�wz}م{�,��9(t��R
���`-�eϺ����7���V��ID����7��!��@�B���{n�v��S;��l�5���.!�i[2��*VU��zg\
`�9;x'F��Z�5-�`Aۓ��eՌ�Ĵm��v�Qz�`����%�/>��nȨV��N��h���T(��Pb��y)���"�S֑ui�/"%�֮6 
�ؐ����������0F���V|K����Tq'!7���i�=��k�_n�}�:���q+�۴���y����bN�B��|��3��v�e�La�IE{�O��5�����VY��W��gLo'q�x�
�DOl،�QO�֊��\�X�ܪ��q�wl?Wt���Uy�jR���N���Y��fe[�3�T���ku��_c���Sݿr��<�MӇ�NN�{{�R;���WFX*�s��vAh�9՝�nԽ���'���-�:�Nk���UO�j�p��Ro��g!��v{;��doO@�هbf9����Pk*�kΥj�\�dpnn1�{��r������!�{�63U�n!�Ⱦ�*�7W��಼�b��WV�k�J9�w}Y��Bt���n��= 붱�8�[[�2V"�,Gs��O;e��*n��M�x;�M�4�b��%�����u0���Mڝ:�.�.!ZQ@�+u�hфŸ��"��m��Y�wgl�ԛ͎z�]���\sV��d��M������zuvN�ٮ�UcMB��{�Y��*E�ҹ�%̙_a}�$��4�
�U�>ۧ}�n����ؗ?����3�
�H2z7�`û{�����g2�a\q&f�U�(���4O6j�5�<��z�������e��`�)V���Nï�n��T�ı���q���Y/9�y���nد��nn3���ʪS�4U�jIU��%H�Y�{����(�1	�.�g呏�ԙ��t��:,�x�V������r�>ue�ՐJ��.�up�r)�ndd�KCI[oPY�f:�ĉ���1W���'�(�M2��]	[f��|��g+��z\*m�ރ���s��>�$�o�:����Wd�q)H9[��`��Ǧ���S9�:9���w̽�8b<�fv�.)�~�w�b�%��hBCs�$�[m<�7e*�Y'P;��y��Q�%*�p�LW	.���T����SҲ�w�	������5�;�m��e�c��j��#}��K�7�n��n3�R�\2u����ֺ�f\q���ls#��\%�>!�AVmԍ�چ-�7���*w><���e�zƦZj�z�!���z/��6G{Gĥr�R��{�üj�Kuҗ�_��L~��oDg�f�VtVk�ɸ�w}�:C��t*w��|����܇������m�:�s��>��x�+ u�5�p�k����|�+GvˏD5j���ղ�?Z���z��@'�q�[��3r.�K�4T�4�r����=�ҙ�L�*����9�+��t�>��r�'JqYYug_س����c�G>yJsd����yp,��P3��3PrK�J��$���uXI�v�Zq�ۅI\ܚ��4we��GG=<�!�8���к��j�����N3m���6�6��5��K��ZW��%o��e��n8&�a6��)���5��eJ��G��g6V����m�h���F暸��5f�}�6���ӧ�W� *���~������)�@o�4�"(fgf���^����(z�:G0;פ*CD:��v�b720��uZ�8Ě�ٜ�9ƹ􅇷�L��DD���^-ޥ�qo`N�jT�Zt��T�<s죥d���P���Fb�fwa��P�0�f�5x�#ií�L��Y�-�lB�(��]�=�s��v� ���q�5�<��� �M���r�%�o�_9F7�G��]G�e�n�,_U�t��)��]�_<W	��*��7���ė$�.T�o�Hɫz��j/[�(��m��֋;����x�u�s�G!���\�c'�s�'o*�]���*kֻ�ܕP�8����=�R�~?*����Z͎���U��x<�m���ȿWٌ�[�";��	9jQ����sx��r��P���s��2�+ �챖s��RȵY�E��t;y^Ŏ��m>��.�������w�Jy9�h-�t��Ь�����-��zS��,�+�M�qӻcv����b-���-b����E���Zʺ�������3V���*���v�ZȞos\7��2�=��V3��M��*���P�:�]	�`@�v&s�o��=�F�H��Jm-�����+)Z�p�쮦��u,�97���l�.��A���GձRNgaj5�QX�Յ�Z_a��G�1�k�ܾ%ry;Ph�z�,�.�)x�;�V'|�3�f9O���$��g����_ܓ��vk���ww�U~Y�_D���3R�^�ʟ7A���X���ȅ���V:V5�v���EA}�\^e��s����47��J�nUD��D�n8�N���.�J�먡Xc��s��Z�f�F�:�����LR�%��}W�Z/��<7]�4t���ms�X3��OOZM,�l��x�ᬊ�Z �R؞�)�[�hv��[xU:�v9S6WQ)�eO\$\Hޗ^-�}"���G��V:W�[v�g��I�@w�o�;6�����[Uאں�Iȴ�sWKїu7/�������D���w�QK��f�i���F���x�'es�I�1LGU�,�kE��}\���2�eھr7�ڻF:����=uq77���\��3�w��ڎ�ȧU8H��ꄜ�6��{�t�,'��~���&��D8��ލ@0��l<�j�[4|�Co��(Wt��I�\M��������=YEM�栕��n��vT�ˍ݌�ڹ*�w�Ҷ��M�Z�� �
��dͼ�/(M��
�؂&��+gw>(�����RG�\<�玩��&Z��Ԗ�|A�/�D9~sg
~Ū�H�Ҝ�KTf�4/8�*NGӮ+,*/�+��~���XQ�/�b�;��W����1���r�U[�ᬎ\N�7&�a�g������֌9��\S=�2���z�
ǐ�X��@�sՉ�Nf��w��j�vJe�%^�㌸�l���Tz���U�E�g�>i�7�QUEl��6O*�����j�.z�d��yJ_�+��.��]��*��6�9�^z$����tm�����˿E��y��0��gxg�	��r�$bq#�'�y7:Uϟ}.t�
U/ux͙�c�\3�~Y��bCC��Dw��l��z��U�W�C�Ku��cY9�+�7�T�*G7������(���(�ʚ�1	���s�=]�d?{:g��*g.{nz���*�%�xJ�������:h\��h��9��X$�k=b1����V�^}���:���-�#��KI��O��GRF��*��9�7���\��o �����&\�j;Y�k8GK�������R3*}��VJW��O�LP�9�;cR�����롂�^X7Z�U�yrG75���������]*!e��'.q5<��g�!3�vx���Ba��*��/a+rZ����yf\��_z�n��Y=w����S'�썚>˩��o�چFm�j�GvS�7�qɚ������.G_�$ͽSb���+���2���cc�A�1��S솗�
��Ȓ�_��z��=	�{*^e�*9�k����7^# �nzu;�!�Ϯg֫|v�D{r�Uo�c���e���,��.�����O^����~Ɔ��8j5��Ӌ#���=C��x?;���U���߲6g�V�����<�+	W�R���Uӷ>�?W�f�a���]C&}}�X��s�W�z�X��!.�߽��}�gߖa$����Z#���׆C��ߤQ
M����S>N'��+>��zD��~��8W��8�f�^�x���a{�̒*��n�dF�Pt��6Yو�V�$�~;�Q�~?E_P����>�_(�~�=�;_�����>���f�ۤ2# q��)\<9V�z�Ǽc�]�W�Y�gJ�QsU�=;2��p��O���s/�~w�"�OhR]>�e.��&O �q�F"��9�w���neܽ��Z�Ɗr!0�LySb5� =��ʰYN�n�Xf�)�M��Isiޑ�7��XDqb��C��c����4|�W)Y�eA�z��D�s��~�-؂V/L1���Xj��&V�w!���6��Y������!"�f��C��b�W0t0����n�ۧ*�ʆ�;A�i��)�����Ջ_)���*Y��M��zU�3����r��Q3ũ����{�/j���'--q�-bU�*gb�H�µNeV;'�N4�r�c�/�F�2�fl5g�
�NN4v]�
�L<��2��7L��'War-�W���7�N��T�8��1�D��g�T��]n�a}t����ӡ�?3])��7
Z�F��G(���՟e\䥖M�X(A�MViu�rQA�����<��S�L���Uݼ[�	�{c��5�偰A�vf8���^��b}�|�ݎ�����VT���}ѱ>�d�G�7�@Գ`T� �'7B�e	+�l���|y�������em�n$lͩ(k�&]L�pe*5}|/�S��v�&��u�v����4Q{����ԧ�7;I�Z�j�k��
�e�f�J˺i�[t+��,<7l���������[�Ź�Xu6r��館Y2�Y�|L[����.�S��㜫,�:��i�bl��x�`��e(Rڐ�K�m]pC.kÈ8�W<(tX�������nZЋ�U���(������U>ڭ�c�Y�J��"3�q6��pz��6��vŌ�-�������U0G�����t;�w,X.��j�;��#�5T����rӁgE�Es���E�Ůd�V���H�Ia�Z��f���ժ����o����m}��t2!�k�w^��M�%�v�
�ێ�ڬ����q���/WwZˆ`DE�O�j�˙s��V�]Z�,�>]r�if�_ ʊS�zC>Y·{2��jf>��/$�(������G;��,�T˨ۻ��S9
��e�y�f�>��+4��D��u��3��m��3gs�
�6�����B2�t�yqS�0���T���i>q���$l�o5v��;���K�����h��i���B_Z ٮ��,2�E�Wmj�)��-�����,�"Ն7|��C=�7��Xkv��4�Ff&�ddC�6�� d�f�6�涡X��Z��x��S{.=�nJ��f�V>��:UÀ%�v5e�d4�c�o�^kQIS�r0���9�D�9��,��G"��%��2����$����4f�+=���ˁX=�1��t��N89�"�Wn+:��铨.l��e��+~n�rOFMN�U�L�����zjW9l��q���X�2;&�Z�8���q�wr���g�V��NZ��(����z�;��q8�ҍ���"[g�F��3��7|�zG!��a�9J,��\�i4Ζ���K0'6]V\�L��U$�O8U\U��;����0��,�	�p�I�Ĩ�N��
�*1akCS��'��(��H����"�dUU�U+�VęL�;*&U�*������$�C"���T(�+���Yș��R�#��L&EAՉUPn���&�T\��J��5�	˖efTAr�T�! �X�UUGu
�x��쨂줨Ei!eu�D]�S*��B���iPQT�����\.˔QU\��ú�J!\)%�	ˑ�An��&U
��=�r�dQ	'(�ZU:�fr���H��<��^���g8PDd�Bt*��fPĨ"@�]�v���w0O�b��K���ǳl<�q�ŭױV(v�݀*�Z�������ռ�Z���w
S�(���lX;h�3Uޏ��,�Ýg.�3��yM�/	�|�ީ`�)�eQ\�2�(8>����c�nt���(d�O;2�Õ�9e���7��bB4=�"������rw�n��=��7��kP«�EO�U��>�BO�4$�^cW�Q��2�J��~x�G��t:P�o�)ot����E{�(0�n��� EE/Z��)���_��+��������V����{�׹�3�	_���O��N>4Nyˡϊ��*mȑo�27)�l��9^���'�g������x�/ӟ{���Bn�#����3=���� �����-2���pb]�����{+�n�����в��lo�i����=��̱�k�̺ީ��{�6G��\D*�:=^�w��w��Q�EZ���K���GO_����U�0�nC����k>�����}Y@ޟ��{�b���h�J�P��
09>���
����X� w���ű��w~;�~����zڕ�4쬬=�ԫ �M%X�z!-�ё0;�T?_�]��ը�}��]����~���?"W�Α�fH��?J��~^������9��.-ӛؗr���:A��%��Y�$6�Z}:D�����q'+���N����x����f9��͔�+��ݫ[,�W��y�E�6�$!m��!�͑�.�J��h;����@���;T{��v�^��?Q�>ޫ��Nћ�m���!��W�]�~�g�h�л��ee{��W6v��f}�i���e/z�ǲ�>#a�'^ٙ��\,�P���Bv�(�U;�3��ӧ2j�q�>��o�°�Qِ����k����{r=�j�<�,���m��t 5Cڬ�v��u��Β���D�\,�˵uq�1�˼��z��{�>�ޯx-�c���XBs�ꉱL,��W^��T��vl}%B��E9C$��{R��p=˯���ɼ��zL��z��z��G���S�;�ʔ�5u�U^zȽ�9C�x"_HP���{ۋ�N��}_W����>ԌQ�f&�ǯ���yVy��훫����w<F���z��Ȝ�š1)X��Sv@�T�w�\S��,�"�W�h����9�S^�N���g���� g��X��_�*�Pt�e��	�^�a����f;�)���^�S^d.sQ�{��Spr!?cc`{֤xo��nFy��۬b�U:�L��Z�&+BYR��xڮS�7��xO�)z�6n�`�^�ȏ'7�~���@��g���f�[���6�sYqk���g�V���3u�!����7�T��]����n�G�cб�Y��t�I�(R5��k�k�$�4��R4-a��:�6>�Q$u�=Jwxh�r�$N7b	-�magRۥ�Bjާ�Ulc�ᨲ���.X���7��Q+���$���s����-�X.SM�F筑iS࡯vG�=�b25�`��?W�O�nreP��*��/R)�;�y!�c�P�!����4Q����k����Nfl�o�r㽑+q>�>�aVv����>��6�ٓ8�b�M/���+����wn��_q�>�$��=��J�͇�1����&�ϮW��y^M��s~�`���̠�w�@Y����_�=1�"i�=~�c�yQ�� p�ͫ���Jww����N<�̝��g|2�j�#�5���\춡�CK��ir;�����{1�u� Ǝ�Dޯ,��|��ߡy�%���[C��x�]x!�v/_n,�,<��8?U9ۉ�s����.� ��5^���������� ��lL�T���~O(�W�/n�3	�z]�"�s�r��2;�u���^��H��7����?4ҁwq���/�9���=��p�°��Gn�ϣ��S���y[�uJ�En�SǏrng����٩��[f�Q����.��>f+���g"�ψ߫=p��AO�	@�q5+�5M��
�F�!I+�ڴ֏�h��HU+�ݶ����0v(�qbFM	�aQh�ꑺ[ٔ�s�����Η+�A�w�-�;��ɕ6,��-J��chB�4s״�8	"y�ض��K���nNͽӵ��e꥔�T��b�:�%N�>��F%Y���	~�����VR�{�����A����b{ۗ�#�33�B\�E��=�ǳ7�+}�O��D1K����pP�~Y��bCC��D?ut��`��U�W�CT̏Uz`k�}g��p�6�	�.Ԍ"���r9�j9��lF�i�xO�����=~�3R��]�c�z��u�� a���M��u�.r;D!Ϝx�s��z�?yX�9���:�N���P�vV>@W�"�p�!W&���}~:ПC��Uz��"��'!�`�M�;Q�cѾ�d����{v��>I_�V{��퇑�G�u"�0��C#��⚾�vS�7���V�V�Og+�;>�y��b��}�w����t�z+�����,�*��T���V;�
�{}���~X=+���v�_�Нߐg�3�4��n(�.n ����u9;˴�.O�qxƢ�yJ��U�y	��#O�4���ú�p�~����2+�Vp��G��<g^V��1����I|9�ŕ菍ρq��L�,6���,,�3��#ҝ�g�l{/�5'���R��9&�	5G���^�=Sz�+H[����k7��94{aDkCp����Ϙm}y��H4��rK;�Y�2���kq�����fT��<�٧M����&�&�|y�9���F�,�M/S�.��gHdեGܦ}}�˯N��|d���)7��Ի�M�·V�p�<v|)��H����N�|���O�~(�!�g��;8�>�y�0���9������Z�F��\^��ᑁ�傡迅s�.�`۩��p9:�{���ŀ�=%�^�g��z ����+��^��S�"��#�Hf "����{тi�>�{��h�Cq����E�=�O����v��ɖF?;����+$`
�T�T'�$��S��o�e<���3��p��ǧa������Y���6�|ީ`��`�b�}	����U�g�<7��ao�H��2M�S5-ߤdM�;�5�M���bB4=�"9������6/ ~s��>˾��<G���j�T�=TQ3)pv&��f��~c��2���T�?<s��Ѷ+���'��N캏����/��}Ab�>��D�	��0�h�K֬+r�/��V���&��o{ΗsSw�Տ	S◳ӣ޴��%�^��T�)�`�+�NTo����w���C��9�Lzןh�4=�_��Uv
n�#�>�L�{b����Hϕ0��i��OƑ�����t�����^��#K�)\d��lv��w�R�e���h�<8�������[\*Q��e�TT���(+|ӘE8��q��<ycN�v�5oT�J�|�Y܍	Z����hL��@��]���N�Xl!u��B�uj]&�U��1E�#(qʱ�3��d����vW����x�/ݑ���e���t2�s'��2l�mP6�0J�nF����P�G�*R�z�I�Dt��Y�8��{7!�'��#Y�_�-�܊&2�3��M��^o	�C؇�����v������U��t�t���s�ض=.�ݑ�Y���~�4��Ǖ�t�P��az��9׼"׶�E{SK2����������m33�����OuQ�̫��1���ў��/\��Yal?^I �2w�u�Kw�C�p<�E��#�[��޻��Κ�ܩI����^�ffo_���a�/z��/��6+2^Q�khv}L!�A�h�p͡�[ᆼ�f����|�ٖ����{�_��t�<{�nG��zN�Y��kht�׽׊=>�����Ӆz��� ,'�^�F�uq�0˫�������|=�{���w���Be̋޾ڞɎ�||݃�_��D܎f��q��Hh9Ö��y�]xg�דy�������$�U�z1<�G{{�=(w���tV1"r�8"~�
 �}obqa�N��}_W���b[��S�2�]<�Z�tR�]rQ�KMAL�;���}.U�Hw��M�Z�w]�����\�v��w��v|)�=z6p�xR"s��c Ԩ*b�[&C��m=
-3�r��-@�x��c�Z"�o��'R;�[j_g'ԥ��.P���k�ܾQ�KQ��}>���� ����{ p�[�y��BbR�^*������h�ⷧkl�3����s�xz/�?<s>�>��̐7ޡ:}~Ȧ u�!2ذhN{8=U���W��ܯq��c�+�<z�,d2���~���=�R<7��r2<�fo�X�_ʩ�zz^�ww���|�Rs�V�xJF�S~�����*~����6��1����߇�s=�w�!	��]>�798m�s����US�<X��q&�n�\��n+��[#�ǳ�Y�#!��g�z~������y�ώx,ʟ���M�~�	W�4�M�{@�ք�����U�q��$��%�=�U���N�˼��=�*��L}ﾆck�M�21������ʆ`wB�{����P�W[^"����Xa���Vnzw�;� Ϫ|���KAW~��y~'5ߊ�"�y�e����=<����t�b�̏��ᰍz{|�Ҿww�ꮇ��[��\vv_M�}[CPr4h�D���/f�歞����������n5yg�hC��a��%��H���8ߪ�����>�ȍU,���V|���T�c/��#�e�vF�֫gc�H��;$�^�u��lI�@�`HU۩HLj+�o݋P���Ρ����BiՐB�8����r����+�c��i]ٹٶ�	)��6&.f�7\�*n��[Wf�'8���N��@�LN���~���~��}�y�����a�s�\�(���FBv�=>��:����0�d��p����XUm�v��#�1�7d�����m�f���<}?+�������xMV+�k�k�#��@��O������}7����FU~�';�˵~��n�S:��Ѿ�6����S��˻���xk�\�9�����#��9
�C��#�3�Gޞ7=ޔ�N��}�E!�E���o=�W�����^��J9A̲�Ii$����_iRۗ����r]j�������#�y|��C;����bBX��?WIϷ��=��b�ʄl1�Hm��X,��iM|4#�p���Cs_��yS*��lC�Ӟc���z"+��*~�S�8�u՛����U_�VSn�b�<�rQ�L�'g�j����9C��L��]�����Z�&��ז���*��Q�.�T�A�n"j�z�L߬m���	�>;r��Sv�W�_{L�j�<%�&��Û�����9�x:c��*z[>�@_T��s�D�P�mH��̕yQ�U�׉T7[��)P�C&
lP!���w|�<3����
�N����vm#[�1�SuЫ4�
��%��IZ�ذ�&�;���Eаi�x�b��L3v�5�<�AW:�9)^m
SM����ث�B$Bmv��=N�p'	ԕ���~\c���r���Wa>�̻�~�L��*���H�LD�Obvhe��Gմ���8=���>)��:
�z�㠯_�ߙ�����튯_��ZY/Ն~Ζ���m(�V��U� �|t�'����s��8j4�4ڸ�^��0XL��n�4��O1�"���A�c�d��~���~5��GN�W��u9�^Y�G��\j��J��Ǡ���B(�x��G;�M_�}�X�ھK2��@����}5�$������[�~��>"�K�u�OH�H��V�z=���S�ڊ�˭��ァh������ǯ:}�x=/����F�l��d�D��0�8{�'>�^�����>[�S�;�e����/���=�|�ޙk/)�q���z�e[����^d=�=~�w�|=��F?;����̬��*�e2���W��\U��L�J�����3�^�TQn����>���R�����t�FNR�{����ڭ*��H�\8+�+�5�J�H��S�#�|��}����Wz�>ҿ *�]�k�tf�����U�Wp�d���{`�H�! Vs�m�k/[�5����-�CRƈ�;�v3rn��F��L0��L2T瓔=��(t˝M�C�mLڇPG�q�W����	����Lj��.�8R!��w��1��V+z�E��:���H�RV�NzP>����z�v
�V=bD�hI�a����}�T����=��;��\w�Ϳ�������?{ p������ȑ�M"����Ô����x}�s�����vU<���'�"�������V�<2f�Zȫ4��Ċ��C��s�C�I������P�ye&�5��0�������Bn�#��������� ���]ؖ�}w�x�?���Nw�g���z�o��}9�I����#�d{c�y�25ץ�~�L����P|���t��]MƮW�ʡ�%@���[+"_�3��N��盐��b��/��9����k�ZO5�,z5t=�ڋU����#���TL����#��W���~ ���_��ФTɟ�`�D����L>�9׳��X284�)@��B����V��VGd���c��w9���>qtzǲf}x��^�HO�XO�s��7�A���*��7	WW�����^��Dp*�#���[=~���~^ڗa{������fK�2t����i|c�C|���a|>��'�\��X�ݩ�#�7.�<7�o�.w���]!�@=O�+8(m�!%�Sq]��������o��O����p/~���C*H :%��Jf�t�dY}0��u�����H���<��0Ds"� į@�g��Ӻ�mL�U��9���,@�YT��� ��-��Ⱦ�oL�*>��P�i��hͧE�|�T�6���QQqwR.3�����*�MBΨi-W!z��p�R�y�R0l�0��;��6�{Oe�H���-D�:��������A"���A��������g�y��p���to�#�����ӵ'ky�#!�+�nJD��:F��p꒸�G,ɶz\��I�U9�����7�h<ͺ"�d�QK�X�ЕCk���r�
�h��2���h�+ �#��6�%*��ͤ�/�F
3v���';�Kq�N�m���h�7c����
�E���v2�v��z�Mu����͒s�o���*3�)�޹$@��0�ՀN�ԫ,�qk(I�����/�����Z�����g�`�1r�N[�0i�f����*tygP��x&#�ԇn;����#Wa�.۝+7 ��frw 0����J��q7����}ח�)�a�Z.��4�|Le���2�K�8i��2r��`���wOt�nj�GV�X��j��W�I\���STLJj���y�tW:0��0%Wd{�W)��Ӥ.1V�f��4�f%	W`#�+L/fcђ�5׵xvO��,	���f;@�(���ӻ��y���hrj�m&��y�kyvn���J;����Zn 21Dd�d\6���z�QU�aŪf��(�[:��׷CC�[y���ܺ4�.�W�5;�����d�[B1���%5B��Wv��U�w�W)X���[@̛V]2��=gZ-�B]ܡ"}���bd-r᮵�|8�I��y�t9� �=��Z-�#��2�{�fnj]��)I��\����A��{07B���vN��<o�����E4�ڻ8�X�Z��έbYB�l���v�'�	���{q�#0d��pt�1����:�P�KN�2#���s��aJŸT���+A�sB����\�]D�n��S����'m�
\�{!�p��η�Ӻ떑ݫ���"�J&�'z.��������=�+� 
���L=��d$v��)�DGP_5�r9���č�F��N6��G���,S���e��wj��U��YW�l�dMf�f���Ѻ׹Bk8C��(��ĝޛ=�"�K�U�bs�z�|4�4���I7@�tN����31�M����T4�t�xn"u��)e+&m�v�ȕM*E�K�N�M��P�[��ŸhB�[9�fb��*�#4V��i|1��q��q�WG5ҷ�^N�:�wV+�T��d�Uz��dUr�㪠+�<\̮�����/)>9�E#�߯md�GF.�n%*&6���cW����T�^wEq�oψ'�@PK��N\�	*�%��X'*0�E�,����C�C��D{��
4H�"�&\��r@�Ci�EQQQ�+�D���� �
�s��(���#��
",*�/'<�W:��㝥J����By�R*�y!�
(�J�L���<��*
.PR�ե28\�h�(�E^E�R'P��tNDDZ��wR
���]΄TE���\�Q]�s�l��R�#R�h\�n�:��WrKS���.I�D\�;�
<��UY܁<�6��+�;��$�i�W�Q=4Q�J-��"�r9��D\����^�Pnq&\s
�g��B9PD:�	2!��p�p��U�j;����rC�4��z����;�{�k)�TEy9�TW

aH�J����.ʪ�N	�s�zG�D��t��;��du4̊I*L��q �!$��@��Eq\��*����g�Vl z�Z�s�_B*�dnhC��\G��vn'�C��k����D�]-յ���'#������hP�p���XώW�|��>�y�_�ϡ:^=܏x/Z���*�������z�ܷ���F��I��p�	W筿�V�K�o��2=~��`~����b�=}'Z�������O�}�[�X���<A��n�����\�	�6����0��ߟ�6��P=L��tQ��L��U�}�����;�)���.Sȟ�@Pɏ��A��M��r�ɮw]{�LNŤ�>�u�{f�W�������7��ݫ����A��(��7:�'������B>���߳��1pPϙ�����2�����>�z��z�*����Hk�K���^3�w���yn�H�N}tP}���CSpq?cc`z���`{m��󽙸u�W%��S��^�`Z8�'����«��RV��[@���?5a5�������W���C�H3#9�Y��#����H?<�J���:\�ŋ�/��/a+d5�/yfX��#��n���,G]b�({U(���׳PG�P0��3�#k�gOZ�x[���JW�㍡�~��09��3����0�u��z�[T�mג[r�F�כ|��܂�F]���q��j�kD�$1 ��X�\��ns;� ����q�Ж�Y;��1�5o;����1u��q����ۥ0�x�m+;�
����vL����n���ʫg�ɅkT��ʟ$�!��]�C1���ٓ c��#K�H=��uD�;������Ϋ/���7[�=�������}s�j�{J^۩�����"���a��N{��=�A,�4�n��;�~Ɔ��8l#No��=:����\�p��|�㳲�o����3iGem�.9��]�U�#��U�5�z8�Bt8��瞗Axx���&c�t^�w��)_�G��=7��;*�;q��Y���4�|�}�^��=��N߇�}5r7m��W��=�j���g���"NWƯm,2�������m�f�_�����_)��V{�w�mđ�r�$Ol:3�������{L@��{n�ϰ ��G�|���r�_�6_P�}�����=~���E<�Ɍ������E{÷�������ڬE@�3T�i-(p4>5)����f�l�ᚮ�yϡe���_�r+"��p����S/��+��ܸ� ���4�{$��g^���L�Uz������"�~fࡑ��+"��Ho���"9��NF��'�����Cc��DȡA�ن�ːyz
45��R��fX��OLsH���[�1_��e\񧴤�ר�o[�����&�3&f��K�z�1����)�r���_��Gq��8�9x�I�/e.��$+*nL��.�T{���{]&K�;W��bZ��_�
�
�F�(lBBU�7����1E��ps�O�؍��9�%B���yWY,鄻�c�����
����>�u��;C�T�T|8�N}�+�o�� ��A�/D��.�=�I{��=V�w�È<ZZ�6И{?J�uG�b��n���=���/�x��*}�,�4۟����9� �Y��0T����E�e��>��ۋ�&���w��:=+���GO/e�-���>�̻�~�L����n9�ԋ���#*j.���RJ5~S�x:�n���VW���U�0�nFA^�!�Ϯg֫~�ۊ9�˛G�v�Dr��n�wy��� B��ō�KȞ��dU�zq]2C�zqd{]�����~���s��*�b���� �Ew�?^���+F!:6����]/*�pt��ϗS��^[����`�c��n�����8��9����Q�M��eW���+�!ND������A���mz�Y��R�}�L���5��e��-	����XX�?�*�������]�� n�Yi�Z�F)}t�D��ي��<ԝ��qo���0���y�MT�^�֛��0�h�v�٬�[&d�+�t�d*�%��L�[��eу�5��D�r�?u9�);l[��M���L��5�mc�����%P�p�������?,w2���d����`��^��~�O��1O��VY����� ��ä$����Y�ߟ	P��j��[p����P����ީ��o{!����'k,ʍ0�C=��Fo�a�X�)"x���ʞ�̀��>U��}"'��{�����X"����h�3�E_j^����3_
��bt
��R8"_H
1*�#�$���>�֦�+��1oe�畧�|I�ön����S����d���B|�ROq��M�#[�+�Q�s�,�]eP��"�3J/5VW�T���zl/�k��Wi?���8p#��5�
ɂ�6<�lw�1Y#��s�]^S*k̅ޏ�{�	�½�s�z�؉�l�.t��?�?�p�
o�?�v���������_����||��f�`�&��=�L��;ٚ�݉��z��h����P>\�[7H�N��`�4�/�q�y]�������>�V'mƁ��.=�w���ڡq�P��S���l�u�:zٿN���G<܇�	�1̢w[H���knXM�=������-����Tf�PT�3ԣj������������4n�q�B=I�p��^��\�ɉ��6�é�3}k���﫦��b2��܆�{���n[7$�X1u�-J���c��p��p���9�m����%�#��Rפ[V��-��Np|�e��
�R�_M/�p6A��ʫ�<�� �s�bO�������Q�ѓ�&���oּy^M�م몱���zp�����G��\���0�yQ������v�g�]߳�5��a��I���n�K3EC�u���~w�m�^9֮�X�2�ֽ���s�z�37���S�){�=uA^Vd�=�:FP�<+��w@�.�&�^�:}��P��Ǚ`�Q-��O��&��G�#�}�#��O�dL�:~�k(�W~�����"Li~t�jK�U���7�c�G�ӑ�hj)A�Tn�Z���r���rݏ!�B����9��3R<��t�Ү�p��M�P�L�J1s�}�::���^z��ǯӛ�9�\>Q��y9C�~�C$���m���U��S^��z3��s75^���79K�Ν�>�0���8��H6��H�5��D�||B�_ �O��L_,�_+oVQ>`{�uK����|�'�V�^W��?Y�F��'��pSu�h���Vq�Ӟ�Qwh��\t,�6b�JM���q��#7�ɟR�5�jq�ڷp�t*V1N�/kE, rWAwX੾�vJ��V��J#]��
�]0��sT2��".�\�:�;�Z�H!m7PnϢ���V����V�Ų�4���Wl��/�G���u�t1pPȆT�O�؟>�p=��dy�̷��n�p/v7ݭ.X��u�����*��MS��o[@�A�8�Sps��z�C�y�-"�z�%���q4�s����甜�b�UNB�#�&�B�sۊ�E��[#�ǵG��򺌆<��:����{lG�%�2=��;�:~�	w�4�|n�>�'ћ�����~�;-y����jS����N��e�-�3%��zc��|ch�2q�AV2^��D�p�}�RUv������gg��'�-�LV~X�0��+=&O^_�:��g�>�<sf�Ͻ�sp}�S��)��~�����U�w�j*��!��ǲ�s�M@�Q��{z]U{�T���yם�V��ΐ"��*��fZ�>�j�+W��!HѾ���kQS6�%�%��`����ߜ�xxX�:����Ny�ud�^�'��J�	�����W�������8���!w��k_�34�|�}�^��޿Hpc�[��S������#��i���Y�;�#NUp�,�S��C�9w��K6��h����a�� ��7���KOP'��3����͔��e^�ڹ�fX�ƀ�F9��x��d�",c8��>�%���M>�v]+��ӄ
��Żύ^����N�t����tᑎ�>��0JwTm�uk}�i�8,{�R�$u"vfN=V�'�����G��W��k�{���Z�Dt#�Hg� �
��p)[������1�;��Uv���Z�D=ۊ*��0��׳��E{û�2��Ծ��+'(!h0�n<v2sa��zv{٧��؟@�[����ߙ̊����EdSy��S�Gc�s,��:~wnY1�z�_F{��ݾ��V���PSP�HȂ)�٫�A[�Ȭ�{�x.	�����*�� �a��¤W��U|*�TSRyt�C�b�*�C�3����`�S�6!aO����qZp�e�7��Wp��dz�¦�Pj� ]Cy&ĉ^Us���W��}��{E���W>0����(�n\���,լ��ؚr�	��� ���1���{?J�r�G�l��ۻ^z\(S^iU�����'�}9�,˖�x?����y5�u!�,��㶳�&K�}�A3���E/[��=�ָ�x��������匇޹�y��zF���0�E`����C�i�i���w� ę(zV�Ë	r�����gǳr�~�CY����o��Q�9K=x)m.'.�.�N?���� x�!;�k�3�8_X�,C�Vvj�m��L0���Z�����=��+S���xқE�ҲT	�rY[Wni��_�\�f"���5��r�����_�w�+ώ���(��${x�b�ו�kb��v'WBԫ)�������V~�^�ō�+"z�^E^秶[@�i�diő�wW��RaF)���c6��^�+���~����������������w�:tZ��v�+�`�翷����`�#����6��S�6^9�`�U�wVp��ۮ0;�Cۉ� �>Yׄt:J��9W���O�(3�钽��36�ؼ*w����~a�$k�3q�n�d``yd
��9^�)�ȁK��<r��o^_��{2�,w3�'ٓx{�'X^�s��ߧ�~�b�Iڶ�.جeXy\���g���-��Y�^�$�
���9W�c�sL2��������v�����z�zz2�r]q��F��`{�Ϛ�t��T�M�އF@3�KW�6=/�����^M���	�|(�����P���۩G=�������Ӣ��R8"~�C&<z;�5Ci�g,�z�Jlp���4ى��}C=��egC�k�^z��w��tT�;�\1�!��-@�JǬMPlМ5Kκ��,������N3=�9S���������~�Ԫ����^�~��&��D��/�X����Z/������[zo'S���W!��׳F�`G4��5�P��rr��j�:nj��BQ��`��%��x���󩴐M�����}QcrL����\�wB�@�]��y��5t�U���h������h��t�=�0kיՐ����S����WG	*ꆳ���-�;�y]�����x��&q?<s�=�@{b}[,󭙷�"�`{۽}�/��3v��ߋS�W�w��'��݌�ezz�����1ps��z�|��R=�L��C���F{��nl����;Uk��^̀P�2{��Ϸ-x�2��yCW~������V�`����S��jIO�c��6���\*�N�'�ղ��#���M���\:��z����n�ϹO	pG�z-�[�����^ظ��V������CQ���W�l�t@�����0}�|��G�z�}�3gӾw�Ϩ�'W�G>�ٹ^ʬW�L�;�/sV��FF��≟�Ӌ���#�չ�#������Nû�
�~������g}�S�������*ǡ�a����ߣ�x/\<�=�D�^����3z���:�C}��j�)e|��ɘ6.��z}�Q�¦*	f�#Lyd���d�����-�[���9�`��3#����,*��z;}�-���wȓR\?:	A����mK�^�ɏJ��~��GZ�O$u#`�w��'jwcՠ��4�J�R�LM����I�)�>�"yӭ��ρ>�r��:���v�	����B.�'.v<\��wLkQ��+N`c���S��4lq�*汳�yZ�N����+��끀���%��_Czx���zh>�T���{��"�@�3	�S������Y~�n��i�5�x8-\.����{Yw~3~�'��,},�}��·�T����ˏ�.�9���U7]8�D��n�[�=�^�7
�﯍zˊX��f�")�gJ�ט=�Y���X�ː�ơ5ă�N�d����kԻ��C9���3>����y�jb࡟3�c�X�|ߐ=�d������U9��0�{��-���+%W�*�3�Kr����)���.
ʛ��'�lo�դ{Ç��G��1�xK�9".����:{P�gƱ
��Tc ]~c�5�jo>Ym'���*nBk=b�]��{y��w㇯-���@{Փ<��UM� ��P�?�r�U���A��iS�{Ir�h���痡V{U��/В̱	�X����I�Û&=��(J}ɥ��pя�	�����]݉Kw�K��*:h4�������\����O>��(?���F���
����v������'����I�z#��_��ה����I�=���N��3�>�ɮ��o�L���U;���G�Pݏy���J�S%�>�i�7ק�<�@�XGC,EK.�r�Uywَ�J��
�ܓQ����T�
��u�C)3�w8��Ğ�w\&؜\b�C��Vb ��9�Ȱkfbf�5���ՍU<ˏ:��[qD��	=ڊsM˖k{q�mr�伪k&�Nd��������(�܎��jgwǆ��vi���*q�*�
�d�V�v-v*P)�'Y6�~�g��S�2���n?f����Z �XR�/Aii�X�DgkesOvC�#�/=7x�K������lNcj(_7ݗ�k"�A�&��r-��&��r�6�C/E�@��ܢ��K��KJ9+a��pɔ�n���ק�*��r%�3����̷��0+u�¬k�]bR��%v
X̺޾��!ThZ�]���C ߢ,�Q�V�U��ױ�5�k�V�����f(�<"V�MY鑮�7%�x�I18����.s۾6)�B��(�0*�
έ+x]��'Q}xp1X�"ẏ�K\���f�g��UډqU')CkU�*�˻��"8'6�e�<���QU��	/�YQnC�~Ɯ�Rr�SU;Yv��u9^�����յ�J�������9q/B�
�'q�p�O	�,sF�sJd�b�[��j6�]I��#v�.�x�K����3��72+�#;�k���f��ۀZ�x��uΠ��u��S�:�<���M�'�u�Ҍ��h��u�|.\�'����ώhk����ʷ�n�S�>�d8��ڈs�-���ڭ�6c�	'�Ce��Y�MfTv��v}�MC7�n慊���9� ��Lkw�����~���������[�9H�ٺv����-�ݻ�2魊
;�7xÆs���J��k�!G�A��Mq�Mhlqi�}�#o7������bgb�[�B���gL�ֺk8;V�d�nMْ�%M][q�t�f�&���kJ��S'�b��],(ej�]g�(K�nkB���K��)l�m��bI�v����Z{��$�;u�����N`���!<ɮ�o�F*,�2��w��x�7b��p�ב���0����q�yt6�Z�8�.���)z���#�V��UY��xs ���PC��qւ��/y�s�+�!�gAT��oIu	���\�ҫ�k-3�S�8��n���,�ɔ��6��TTƍ=�ڡ���4۾z/Y�5������f�]��e¥��X�Z#��'u�|��-�5���ݴ�7æ���|z�1��{ɇ��#z4 ��3%4�a/-�;k+����CDŨ�e�5��E�Z�;S(�����v��ż-�1󭣲as����W��3:�2*_�z�"�t�u��2�!P�ɼ�M�7��'dG���7�
�Ymb�g˺�=;�N���"(������P�WUځ,9�W
t]J��y';/(��D�sts�W ���%I�E�n�V�DE��(��+H����p�%r�(#���/jDʈs����S���l9�J'"<�T��ҝ�)�'ZY!AZۺ�<�G �
�����:TAI��\Gfd�&9�A�j�X�b�c�:�E��v盭u�%(%W4J���.Y(����iu���"������"��<���N:X\'M����iҊ(���;�Qp㚴�+,��]����i%�j�U\�We23���)�u�̪��(�4����"ww&QȲNx��*2rp�Hʤ��%��"�eRN:���W#ͨ�Q�(��wR���s�(�z��Q��9�Q�-�.�NMeNsS&���t�\�:Ȋ�yZ�"$
+Ȃ	�p[��{�e���sj^Ǚ\^P���*q6���҇4�,!�c;�'�{P��.�Y�'^���Z�I��"���^=��Zf9�L�`� �xd�+m�E� p�i�gǱg�a�ߏ����y]El�WKںg˱/�!4~�H�L�F��~
�ټK|�#i�[��'��{��GI����]�����>2�;c=�-F��B�"�G�KE��t�Ꭸ%\���E���ZG�Q�m�Z��C/&+9�ý(�-]!�}�k����[�:�d����~�����nE�]��3_�k#�*���^���I�I7��}^�8���S�����>:+��v�� =�~^�w?��{r�g5]��|��ۭ��q^Ǐra��t���xv�z�Y�~�>#b+(���Nǳ6�����j�A�^�{�P�j���9o��w���YM�j�O��\�#7����{V?z{��z��{^��WW����K���$�ЏƀM��iM��{4Jo�"�+�Ć�[������]\����Ӟ��W�OxS�:�\(��9ݙC�s��(2�Iȩ}[��q���#�,<�u����:����d�]�T�U��ȓbD�*��X�~;�Ys%R�d~�f��e�E�ē��3G�I�t!(�cӠ�Z-x��qCf�BCKgeX̏�����!���J�R����ϩ+n����<ya�uҥ���Aي��# [��knebe����̲&^q���&����:Q�TD;(wJj4h�P�ܕ�~sބ�	9�k=.w��,=Z�w�<��>�ihHw�cm�~[�	R]�{�
�K��唙�֭ϼ�������%L���퇑�O�u"�0_xyo�=앛��M�J7�{g8x{n:��I�{r��Ӿ󼱏�s.��=2G���U�٥�0�G���*��Ԯ��#�\�$�ᒸ簐l4<C�����f�b�>��Z�����U�S��yw�{Ů��^�^{�7�j�����rT�t�[~��[@�?qdz=7�yS:�}{��������ݦ��W/׼�b�t!���U��:_}W{��E���5>(n���.�����ڼ�����F�;���g�z�X��y$�҄�\�*�&�e(���3����G�[/��b�܇�[�����'W�xT�<^�H��_���$�{Fo�;u�#ʱ�[�sg\��>Mo�]�@�q�S��Ck�%�~�!���ԍq�}����o��N�e�u;����Ĭ��B��9� `Jcc�J���ʿXz��i�]�5��p���S����d{ʬϲwދl��[(�G�Q8-i�U]��19ҵ;��ʵ_J�-�����4l�h��HA{{NзXP
1ۼ�;weK���"-ᆟn�"
̳���k�L+����"�]>�{tb��k�����s���YA�u5v>]fMZ�����Ŭgnt
�u��ۆ��ߥ��<X2��:>)-I�>�FԶ�6�׆G�דx[������y�v�+�Ѹfk�A�����SN�TW.����Nf�U/
�)��Y�>����c����J�}ח��.�=;����QŴ/�,��Z�5	����/��4&Sn/�'<p�!��B���5�GI\�ɐڵ2��y��#}��=~���(0�$L����&k���o�{�_����vQA�5�����;����V�<�f]�����A�E���Z%_��H��%�;�j°��0�C���.D6��1�֤{c���f{�v�F���E���Z}��;�x��ߨU��تlJ;�3}7�����䩑���=��<�=a.ӂ�y�ؖ����
ML�yw>��mP�P«NNO�e��D�8�zox߈�y�$Ez�^�Y5[�*�т��BK1�g�~����������V��Ѣ���j��:X��+��]v���E���n�/ �fϧ~N��5�Z�}�v�ׁ�]�ã��o�W~FV���F�~��b9.Vd�@o=�v�i.tDƒ���O|4�7c7�ꓶ�'E��ݔ��X2�c}�>PNQu�&X�y7uM�:P`J9D��.�҂V�@��]V�u@�`w�/�����X yc�1�Dsy�ds,^̗�kǦ�5�b���`<P��$���}ʜޝ��)~��cC`_�����37�垝�w�>�G�8�F��3�ʩ�7�쮊;:����%��x��Dv|<�=�k��u� �"z�3:���)�/z���_R�&�}�{�/%�1�����1u�[C���s�U����9��r�O���2�8z�ax{�<����r�������~�������|�#���$�Ip�D���[��8��}y,5����e��O/Q������,{$�`�L6���<dY�c� �
s5#�9�9k/#�>���ޯ��|�jj�Dy�^M���=&t�=nz��Iki��}�W�:�r�r�%��f�F�S.7ҧF�=�K�Z���ʨ�[��{>�{L���߳�a{��.>��r7֤p�v�D��m+^���y���l��^���
s3P9� ��z����3�y�W��N�{~@���d������B�Xp?\U_�rEt�U�S^�T6���ŇBj�� �h{S��7�66�H��;�����Jמ�k�Fo��B����� &8]62�!��ںht�B��x��7,���T3q��]�[��g�e3�> cR�25<�֚n_j�b*�%Cl�J�8�����s�,h'�ڐ�։�ޮ5�[Rj깮ML�,�s����R�F�w�,̚<N)Ǣ�|���|\�a`'���rm����G�h�\s�;I;�@[C�t�ެ*&��Y��ǒ��<6�|���:�UR��]��U�>*7�/'T��N�-�r߳��oR9~|��7v!$�P��^�>u�<k�(���M{D.�N͉��`����w�	�g�=~"���Nfl�o�w)��]�?W��B����R.:��1��3ތV�zSw���U�F�D�B}W������|VzL���I����>���sf��m\ҷ��zPx7;�=F��{
�=R����8w\{"�s�l@�d�4�2 �,��;���WC����@�F����w��*�
�Wy�zo�hnA�H������b���]/ ��:�MƯ,��ٷl�k�{ظ�(����]�w�~y	j�����h����۪K�J���Y�>-���5s]K�f����ʘ��^��Ou�Fy����[�:�d��P�9Uð0<�9ۈ�D9v|<�/ב����&��n��yc�AA�\�������������ҟt��	�C00�#���q ���=�^z�W[����[��QL�{�~C�Ν�E{÷�s,��9�YFU���	�!�ǻ� *�$A^�s�L��.0T	����s�2Gw&ÈQ����m
a8��0}y�4ROLiiҍր�Y��+��Pl�V�89�wnp�aX�;�%y;G3��de7��f�o��?0fM�OL���jq۴R��Q��I��:��U�P�L���L�Exe��"��o=�xO�s��̲�]	<O�ۥ��a*o<|�@�K��A%�H��y7?^����ICbߖEg��bCemmS�15��my�j���e�ǋ��wޱ;�LS�U!��@�׬MSvdg�S�s��4�x_]7�l��6����>��j��x{Ny���1����]�T�Ψ5Y��Bv(/*����Ǧ��]ᾪ��t�%2����)^�X$�&���}�c��U����X.A5��}����QٝIzA��{l@.���Ϫɥ/�y<�^�A�?%���|N�c΅���{yy�[��صr3l����J���މ<�D���^`��ß����w�1��e�?g�H��F=2���z�ϰ�Ǳ�U!�H��:�Q�Y�~9M!�Ux��ٹS�b}�QAz_��>XQH�5��2�NTWy�\�j�:��NVOWKȊ��Oj�h7�4�+��V����Ɵ^�D�Id��o�7V�9���׃�,ȣ��x9��`�<:�*�?��Km��	*쌱�G�_��t�]Ȳ�l��ű��Y|DN��òn��XA��k3Wb]�p������ɪ� �wW��h�����F[�QgO@�q�J�\�Ե��ZWH��"�_v�r�v^)�Rv1� سc�W1��t$ЬA.T��d�7jf��cӮ׳�7�|��~��w�zDo�����V�Yu��^��g՞���3EՑ4�e��s>�~��S�C���e���<�$���f�ӷ\)f�>��z��p��;��Q�%��P:Ԩ���uR�\����|=��/z��NY���S�.=�B�� ���d��y]���UK�@�=���9W�eT�y�����Gz���+�P�~w�����j�0�ol�W��;Y:z���|:>)-�D2`�C�6����]xd{=y7x<f�F1���ǯz�.1y��H�Gz���o�C2-�dd�-@'���QCT6�����EV=���ey����w,6��OJ{�d3�[^��P�e�Ĥ�Oq�V�.��B7=����n��$�J �[�(�ϙ�)S�^��;�s�z��27��3�늸b�	��^��{�3n����~���M0"���cW�g��/!��L�~x�G�ho���`dy�̨)���j�>�;Um8����R�ȀhMEx߬b�h�K!�a��~���֤z��G��_��Q����%H/;;du�_�m���+d���,@k�4yT�mz�'/Q"ai�.���/�@$%��$�y=��L��[�+{��4җt�SwM�Ga�a䎐Q��[o/�������1ç!���2W*`�Ը���p3�<�}ѧ���}�~V�U¦�O�P�ئo���xu��2��x�oOP����X���e[��ǡ*^�}�z�O��M�ڡp�Uciɏ��-gN5���rhLq����R�9��V�}�7!l7��!�Ez�q�w4r#ײ�؝��X�_O��}^98^ɰ�اc���oV�a�S~�2}����� �fϧS�-��}k��U�r�ٹ^ʬ,׺ ���s�&o�s�F�V��D��*�-Y�ڎ9���,���
�~�����Ih͵�מ���Vڽ�gѺ�-U��L��p�yk��O�=��L������<��P�e�3B���ɀ%���\޵��k��~���t��ݕ�=�OD�P������q>c~�2��Y���s�z�wݧ��<h{,>�܄�Ͽ_]I���<��w�I�.����w�ώ;�	[�^I��> �٩7��W�=��m��w>��^�[���x�� r�Qʩ�+eC&
��.t�����L��Z��:�V������tF,���A~�I������,s�}"؅蜠���I�/ߺ1�+�bb�`����X��b��N
��d�e���u�e+V����:������6u�)����:{^�e�� |- � �9:����Q[갯Wp�����'J�6�2R'|��n�:�]Uњ���A����D��'��L�o�N�;�]���U9U���r⽑����Ȧ��+�^`���x�Z��!۸z�(��y��_z��_����J�S����2R�}�C�|�/>�yj�y^C��� N<�݃ig+���ӧP�8j�k�z�*�Bg�O������"��.
��8���o�W���#ص�\��=�{3=��;[#�������U@/	�ؒ��3n[@��)�;�� yǶ��tV��f�O�y%����y�V�k���V�m\
�^�W�q��\��.9�}�ͬ	0�M/�#l���X�g��,FCo�(g��z$�]���
�`��Ш���_�Vu��Jex߯D{���M����q����4Yo�? ��.a��1��2q�A�ʗAz����ۼ��P� ��5�;�V��lB��]���9{7=:�ߐߙ�υ��͚#�^闽ٹl�c����vaT<�Ў�N��7�l�0w\<���.���O�#N,������o����{�Ȭ���;B��z9��v}۝6}[Cr6>+Rv��QS:�1�%���;��/.�qvs�w���l�[��!���0�������
8��Ƭ
�B*OXЍ�k'�����	M6�]�.enM��5�!f,hL��l�z����&S�Y��糠���	��ibYذt��G��w9]Ii�4��q&vq���^ɞ��({�es_�BJ����UӋ�8pr 2��`39��-ϽK�O�l�Qӻ�*��2�'�~�����]?P�d�;�"��������rW3�*޻�8��u�3{�n>��n·S��I�低�H���Ok���l{-O���".ۤ7��� g���y�t�:��=��#Ԥ�W�҅�qO!�ܘ{{�ӽ�xv��e���s�%L���Y-��t�`�W~��D�-� ��(�MmK=��G˄��Њ��j�O��t��'&�Og>���{��b����2ˠ
��GA'�y7>��E6���6-�dTf�C�o���u���a�k|�O�����)�SV8#˗Ѝnt������Pצ��#ەD�g�'<xԤ��!���ј���P�g�C�O����;"U糲l���wg��ח�\��hw����#�`���������լꌉ�v�Prk��͇~W��;�Z��|*�0�	}=*��>؛�t�>{ԋ4��=�-&d�@��=����{�xx{�cm���l����1����o�l����cm��c`���c6��66m���l����1��Sc`���1�cmc6޶1�cm�������66m����1��Sc`���6���6m����{����)���,% o�9,�������_���0���|���@T�P(T)ARU	*��!RR*���$�)(@"�*�*�%"��()A#wzx@
�
P�$�(&���J�PUB%(UQ@UQlh�*�R��)J�P�$���QH�D�J���R�RR�E@)J��(���U
��P
�U	�$�DE���$|  >�]�ea&��֓�ض�����5�[%R�aCV��g�uUB�T�B���@ {CV�J�C ci�O�� �N��N�@ .;� 
 �� (��: Pc��iB1
	(!Q
%x  y@zXm5�m�m�j�RP��X������lD�$6��c���YD"T�"�RT��P  ��
�S�А�0 -��h� �t(f��v!�br��w*�u�*��D)ZbUJ�U��   ���)J*��Ҩ"8]u]i@1ۡJ�D;qt�X�V�UZ��Uʌv:T�*5�
3�WcUU,�D$�R["� 7��WZ���j�V���1�J����U)Z#�����l�UXl�����k4UPj-
*��H�MD�!Q� ��Tz��6���UbiH���X�T�k-k@lLkRT�!���4
�؂��V��J�TJU)*P�)RN� r�A-�j��!�ڕ��[l�
��4B�*�jf���� �h��U�Z�`�*�SEU+mJ�T��Iy� 7{bkZ�VEe�kU
�EV�V��RJ�hƊ�Ci�Ti
�Zʴ ����-CdM�l-i��m5*H�#Y�H� nj�P m��SU�����P,0�5��-M�Ȓ�,�(��G�$
( @ 4�*ULL 0	� �h�)႔�T�U����4a4H���4'�1�=Q�A�l)�����R��#�4��h 2 0��UG�O�� h�     I %Q(��6� b02a�w���俿�����u����C�����O&p�מ8�"Hٍ�,�DIG�\H�@�A�D�#e���Uӧ$DD��%g����c�?¼���~�ٟ�����|Q���REU*�Bi	�)-Cy����!G�R�$j�HkJ�*��D �6T�^>��~����\�?��������~ԒI$��I$�I$����QP���.��.�@�H�It�*(+P���Ej"�TV�*�*((�DPJ�(���D@j+RH����.�".�I�J�-EIUj�T@**"$�	$�I!$�I$�BI$�I$�I$�I$$��?7�nҲ׷<�/���Y�]i��mt�*�=�{8�V��������ߍX^Yz힙c���,h�ޙG$f�B����p�qeo��P�C4����#K�C͒^���m]f)nF�w�䣆�Un�/y�|��8u`�]�p��(�+�c�x�����%�%%�;�eJG2ø&����m�ҡL�d�
���)�M�A�L�)��X�(UئQ�l���R<�	f��;��V^�@�W�Խ��l�;�:na���%<icww�4����f��K��*'jΝ�K>:h�����ɦ���ܒ�M��;5��K�mjK;si� 헛2���RJ���ޚ�,���a )���xּ}���0�벟�Ѷ���.�']k�������k:�ݹ7ad
Qt7�s)
�5p50����g�jl�ֵ���m���\[{tp-N�/�+8J�Pl<:Yֹ#J��*�W$ M��ˢY�U%Rb/��E��P����5z*��dv����霢�;�Z�j#Ku��Ax���u�h��,��ł������U�*��X%j8r����Cr�^I��E]�njFރ/I��Z5,ݳ��3F�TD;�\���"�ol˄岋��v�B���f����q՛���Rfd��e��uH�f�ïYIe!�9����1S-֬���M⊯Wn������9Djoe��o�P!�)�j�\ӕ0�a�1S4�p�*�;3%8�`�sCZ��*�aݨ)Ǌ�e&�5��v�"��[lUZ	b�w��%�,��˪-Ӣ2]�GⵆS���� w�#
���w�M��k���.wD�7kV-ح���jb��b�IX.�;��`��%%���b&���%2f��y������9�8�P�f�+Py$�B���lK��L��ta�CM�-U�,�osu�kM����5�5y��Z��e5�L����9��U�F%Weɴ�f�m^^�h�5u���O��k�YoR�ڰLX4�����^���N�I�V�Sg�n��j��fr��"�Ҩ���7����*U[�Ed$H������a�ut�])v30GE�՘%�em4�h���Ωolk���v-F존^g����K�Z8��ڍ�jw�U_9�]���^��,���M�����b�u[1���u�'e�7��x���z4iȧ��V/k�4�t�2q\��Vj��c���{�WW6V���ͫnB���V��k]|ԑ<,�j�Ր+�/3]L�ͅ�;r]8sL�h��k��mo��#~�C�"ي�յ�V��u2�T/q�������o��nv�u��$� E��s�h��^����8�`)e��6V��?Y�!47��0o���j
�s����8���t���4[�4��������_G�eiгaf�e���42�h�ٛ[�`��yz6*]��ׄRc]��٭�*�pGm^�;�];�cq�lK�'C.l!]��[����/��%�J���Y�f�TKE�F�2��Çv+*M@�TZ��)�bU6��Kʥ�U���
f�Z�F�SRF�Ķ�3N-�)�[M2��5H�����ҝ�NV�z0��T{x�]��I���+��tx|Cn���gp��/��l�x���e�ŵ���ȫd'0��n��5���8t`zj[ز:"��e ����Z��y�K��g�f�܈�˂��xs�"ܡ˳em�{2�,A�)���;U�]�+p�@,mhuY�l-Dͫ�V3�<��-vG�H����R:�Hg���vŰ��Gx���t��>Z��}cp�����e˱�b:N�݋��e
R,�ݺr�3F�787�"�71�-e�P$��Q k�i�.��������#u��WH팽�����J�P��Sw$�ެ��23m���������H�n�K�w8��g%r{w�l�[y��p�EX��h���N8��̺f�Y�$�2�n5A���2�]��"��ޢ1�u�o�coM�i�B�����OFY����S���qd����ʢ�a��D�0Y��,�1C��ЉՐ��h5y�ilR�F�uut$�:��賻/U�j!�(�u�	/s;>w�B��:�a5�֣�`�՜�,l����>*�*��E�^�S�ޫM��6��Ǧ��uZU.�X)t�O.��q�A�e��/N�j���ksr	/~&�{��ѻ�C+�����I��ڔ��M&�()X��A�'|y�K>f�wq���=hW^���J�C�Gcd����]�O����P�^^�]� �:�;�N�@�����:/i�m��wsM�$�!�mu�(hՙ�x�T��5љu�Z�u��;�)Y �k*ޒ2��|FӨlG�<6�Qb��Ĝ-n�zv�N���*�� wo4
<s(q�ܺR"2�*�t�ܙ�v�S�aM�-�%�f�`
�W[��&�w�ǆ�Z�Z�'���7`�ytq�"�)�;�r,o>�yWn�f��,G�^��ۡW�d<"��W�cdM�͢��wQ˹b��W�Ǳ�RF��?<�\C(:u����fh�#�+Iw��N�E�iC]�UF�)�6f5bML�(���6k�ϭ�tN�MuJ�&��b�j�P�BD6	�ob�)�S5������'Ϲ�XY�3�/,�x�_e]#LZ��j���T�0��c��9sV1���&��A۰�����
�[hX&�Ė�Z]s
�4�*�4v�#pOs,M�z�#�b����[Ɏ@�gv�V��y�*��5����,�'hU�_;�+Kr,܆	�N� �R�ӻ�P�0]��	��Q�h��#��BcU��+5ؾ߯���V>g,\�l�WrB�L5_;̽���ג�Q%�F��v2�n�M��Kl��hT�֑x�WJ]�6�:����iQt�;�YwPdۏk4Ķ"�V�YZy��B��M��/�B���^���օVc�R��V��o.�TQ�F˺d�b������'W(�ê�&R��T��K�y%A�cYX�%�2w�7���OAd�z��}�-'�^Tʉ�7X���Jgu�ݨ�+	�l��]���@� ����B7f��U��}�@c+�ޠcm�/�*�vf:����.���B�όwJ�i�q�1j�����F�F�U�R��^����ӵW��Lk�O 7�l��D�:��{�5H�Mo`ɴ�<6jX����=��sj��hS�pl
P���룴�2���*�n�x[���am=]�>�5waYc��;�ņ3㉷V���&1�k)��ND�7�5�)e��wqg��|G�{�x��t�<�V�$75�Y#4E�Wn��՞���4ސxP�oj�>+�G���w����U�+=���BYEaҨ:�>b��`7PI	�5r�&��Yf
���.�Rg^��(�n4�HkU�ݶjmj�8��Eb����5[*\svg�ly6�2.��*�8��m�%K������]:_|�f�'a�s,4r�
�K�0��1���0�cA5R�W�*��s.��d($�XM�]wn
u�Ŋ#gk�[	�@�ףsyy�=AST�#�n�X �|vެ��qbY���0��K(7�+����U�L�)���aD���õ�I��E�T�e�Y���L5�Ŋ�����G(�b���ot^b�n\ӌ�/�BE2��0UF�m#���͎�C�����vcY���!Aѫ���A��q#W�m�L���4qRm�Żv석o$O0�ݲ��+|��h�U��hz���l7�'�N7��yu�ұ�]��ǐ�9e#[-5�鹂�ʂ����f��;MpP��/V�dm2��y���w	ՙ�ٓЈG/fc�Wc9������+� �$�\t�vS���c�u+t���!�f��F(���6luyU���Wr]����n�V�9�{�Z���NY�D��c!v]k��uq�ƶ�u��5�lݣW34<��JAG7-�w*\�N�F-`��R�Bw�{FTK*�sD��\�5P�ЩR�L9Ts0�B)��[;�6��l�[<_v,X@�lqV��L�i�+[�b8��7j8�meMV��ȶ���*��5���f���M��j��#;�ud9ih����΄��@��2<���1)����Qʽ���Z�gh#k�K4]���`0�*QJkb�^(�[g7p�R��Fm�"�I�3���d��,����]���K���l�]�ӎ�U6���B�ea��In�[�klK]m5)��qn�kRO5�����ڠFl����dp�j�3�[	�S�u�����,C���-��z6��mR�QM�J���^^��o*��R�(��6��KŒ�Z�Gs,(q��;�ȼ-��.U�R�����%��N|p$�e�Ղ�u2�փMQ�΢0O�Xx��h�ޫW�]2,XЯ)K]ΈY�z��n�pV�4�fRI��pDwh�Va��+o������nb�B�1t/�k���#�Y�8�4��C�o����A��[�iMt�&e�cY���X�Vݫ�m¦Z��j�;z�D��!]bx,����f�ô7P�)�-�$&�c@��z_6��]�s��j1�m��Y�VU1R��x�e[�gQ���J=�	�kZ�.����m�v]�ˡ��k	�c��+�僵jV�I5CᚮŊ���E��$Uu�QҒ�<��ܱx��&��r�3�,�D0����F���5���rɋ)CS0�P�1��ڋV����c5-(�O)�n�eahe&c�yF��˂��HP�b:2շOVf�Z��x�����(�t�Z�:�1�� E-�X��nY��%����:�ga�7��ED�fL��
�¥c�DL��"����0-��g^ ���[{Y���u�:��2�oe�:m��(�x+6ƣ����l4�	���Z�[t^�-�V�!Y���36�^�bi&H��0c����7`�ފ��j~��E����,ǂ��mB�ވ����P��v��5�r
�� M��[D�X���M^��8�v��t��ʡ������
F���D^9�3bD�*�tX׆��n����;*��Z��Ċ��|�Õ�w]�\O&����ɂ��6�^�Wt+Z��'�q�n�V湗R�-�Z&�ٖtզ�-HmYz������tY�Q-+U�A�JQC.�@�)n�f�i�^���=�
&�X��yK@(�a�X���'`�j+m���5Ԑ�Ҙ�\0p�ػ4o�YB�����.a�������7m�+�
�(r�~B�J�ʲ!	JxA54�9�A�D ����8��~�������u:�+eƹ��w&ܥ�E1;h��ǖLp�r�)mF�4�������_˜��������R�n�� �F#��)�͚H���*/�ղ����<1Y�[rr�]��C6�:&L�|��V���K
���N����!���XvOF6�\��Hn^v���i�k�Ÿߛ���G�g��VD�4R�ܪ�c��6�f��^��ޫ�[�R=���y.ӂ��ss�Q.n]�OXe`ѭ���X����t���A�lzR���gT��h��ϝ����Gtf-��(�S;�b�qu�ۭ/��mf
{�}��47z���j�YY�����X����1��x�Kr����(���
���MZx&r�@�C��v�}[���[���qM��+b��vڢr�9&*W��>�7�s��>�ڰ�ʋ:ޱ8�!Xk+K��w&�6�$����!���YN��$����~ɶwUA�ü��5|�:���}�|��P����gk1���%G5I��q-�:M�v+W�A,���b5���]f�םcf�*_6�Y�F�U��J���ø-�dN�-�]*����1Bt��Y}����h�Z>[ݭ�t}�V��,����5�ڗ��/�G�h݀�1����Y#��*�H�S.-���
Hl�3z]ʻ��NK44.��&�u���h��ï�|��ws��ٸ��b�E��Z��:3��R�Yc�s��A�l��3��{1�f�d���(W'R�#a(�Ǡ:Ѭ���M���G�Y�7�V�fɝ��*�b���5�۶�v�� �C�؃���種��6�Vm+���E���|t�a�����9H�\��V�*Ŵ#��f4��O%�b�q�����L3o0
�fµ5wm�q䵸8���ld�j�����p�8WoCL:�FS�\j��f���,�W\& ��l��KA���^�Bo7�N�ݽ�ެ��h��}�3N��E^9+)��xHy>�s8�[u\]��>��]��j�+.�澙'y�Q��+X*K=qV0���T)����J��jnM�����7A����q_^�I�&V�;y5�l��ue�DQ�6��*Ȋ2��*���[�4i�w���'j�ʰT3U��S�E�[�uL4���������V�x0jG4�4�\�{;��r��3O�v���Q#k����w��S c�\ݓ&=���Թ �̷ܰ�dD�,<eM�&��f���ˈ��+8�(%�{�8.��!��Y�h��逹hMX�C-��:p���kj^��4�4q�c�]e���v^<c@�q'Z�vb����O�G�ݤ�L�n��xq����bzh��1=�Vn�S��-����vog������@I<�9B�,�e�e�$ͣ/.����sz��#	�6t0cT{u��f�#�c疞.��sX�b8��mZ�h�8D�h���%�P��GF���*��#nQlvqU�
�c�rc�����gjm�-O:�d��BZ�������
]R������_l+�� %fm�+λ4�E�|�*�/쌅,���ȢA�d�xxɜD̗{GB33�G-\&Y���O���w��L���(c�g�Ǡ�}����}�����Z�ӵ�Տ>榒ՋT�0K	�q��2�U�b�R��v��yh[�§T];/V=ǜeo(�K�Ւ�Ᏽ�&�w���7fJ��8#�=�
�"�����i]�λ+�w(�Il�i��Ս��pGB���oP�1��j�t�i��D�߳�E'��9tOe��`غ	\�2�a���tm��۠1����PZ��8�2�S1��ͻ�DХԬͲj�b{j6,ftv7{���f���벙��_m�5��P�2��h��Ƹ�L�:Ƚ�T��Q�e���DW[I0�mC���'q13�j���NU㽭��B�X}pUc�Lє��O\N����>af�e���h�֧v��I#��-���}�F,�r�+��+�岧>Ȼ�9ܹ�E82���;PV�ڏ��rA�N�Ru�"��7�$��������zt����]Z8�'�����6�6�k�J�����ʣE�.ޭ�28���w4�����4�y@n��%圬�������	[���+��n��)z6� 
ڸ0��ZC�bU�@"v�[vFn�&v��⣓�g9��3zJ�v{%��ׂ�}�O�ZXgWb�i���M��\��vʳ��.�mk���C�>�G���׽nm��-Zy6��t(W5g��T�0tv�����彇��[o*ùk����!�-�K��Δ���K7��#�]�������fB�5���D��Yg�L�T�#�C/r<|7M�*ƺ7�+fJFXl�ڹ_e�:�nk1oPp��wby{�r��$)�I��ڷ�,���.wL��8�;��uZ6�\�,�����͞4��"�������>�K�iJ�j�_k�-4�F
�,��%�� ����X��#�.��t�ϵq�׶�@���a���P3�P\�n�`N���m�Ib����=����[��"R�%+�`�������XW�y�*��+��S�h�o;�N���9�:���N+�w\5pu]��G/���[clp�@*��挆�"�^�LʊC����/w�@ ��m�V�9/	��!QeF�X�l�:�u�qv��n��/�.d�2e����X�4�U�Ь�l���ڀ���Y���TG+G~�,�4���\��gA
3hM��\�GUHʣ(nbP����,�<֦v�9)�c�fJ������CV�lt2�{VrB�ͬ��I��۽�W�$�Cq�@�eRU�I�̬���orN��2����6�:����k<r��pw�oYQ�v����nG�%�6闵��5�3�a妲W�˸��$1�;�8(9��y�{����bB��UV[`�7�E���E� ҳb��L�x�N�Lr�,���~��#�CP�2����;t�.\ �'��V$��wY�{�/�l�st�"���d���Jq��a�6�lv�2� J�Yc�dx�8il0�w�����:ۙ�L��)� {r���YAea��
�}������-i���qr�6j����u��Z���+��6˫��F(�B��z˼��۠X�)�LG��9 ��a����\Sk�,�a���n�3W �X�-<A`N�ax��P��avVu�����wk��$y����L�y�\Ga�dx���gn�s#�<s�>���Qy���Ž}W��ۡ�ѓ/�z�[{������g.��`e���d	/l"��W\�KC@
;�Ef��k.��;���O�]7H9|ͬ���b��~4٭QjF�m#��j�]&�K�ۭ8�R?hښ���{�o��Oq��kѐ1ide��Hzg.$F[�zZ�K �}v���(�,c�O�p����hb�書��#HI��^*��p��� ~%u'��U�\�ӱ]�Gw�֭�9�Tz���7[@�;�ػ4Vȅ��@��\�ޥ���pkWp��x@��X�t8n��r��fb�]k���Q/4�.H�!黓]
�Q`re��\s�&�֪�t(ع�f*�H	!����*�V�H���Bo^��Y��WfM����u�ǫ���<mVT���I����uvӰ����$�S�y҅6�A�]�{`Ka��⍞�,����T��Y����5�+�Ϙzܗ�,��n�r�BL��M��!l1+]NM�f��:)Iq����diMג�uW�)W,mi<GҞ�KK&�w��Q�X�$��\ukތѦ!t��ދm��j��|S��)6�C�d7&�H�$f<��Z��**�m[gd8&��{�Q��i��[x�����8>�t��{Ư��k���yob��w ���bf�Z����#����;�ޥ9k��7�K��I�VY&�Y�gK��Է6�t;\,INۦ�V�w�����1(�|�ھ\�w�\;�֨n�d��8+RKb����z��Q������"�ŝ0N�d��Za�ꔠ�)�t���7n�Қ�v�YG��e�=v�h,=
�&
��ڢ��<s]\*M�E��r�!����t��P���2Z�#�;�G}V먘$:����+u#�Ʈ+
�n���T_Z�
�12�oy�2;F'#me�O���V���Lʚ�:K����Զzc�tr����V{��_o5��xpW>D�0���!7-s�wǺ��"txK�b���l�-�-M;�F�7D�����
r{�˚N�a�w���g��Yr-5S/]�Wx�Ddeq{�V��`-���d�C�K��e
o,'v���
L_Z�+ڸ7��N,�9�Ԩz��F_�s��ߣ��.oc+QW(�	�V�Jom��K^��,���`Ҡ��E�M�{eS%K)�M�����0A����l�O=�$�U2��&3��]oT�N^��x�ifT�V�ݽ\p�9sd�O-C`����=ˑ�̚�ҶI\�(No���<�Q��,g����P�L}E�[=��.��Y�U�t�c۪�V���Rm��u_t�z.TUi�C]˱,���So���[�!�`��dp�s�㳣d����!F�ꎶ��X]���"�"��U����u�G=c�Ǖ�����f�o��� ��A��(�U<��-mm�1L�`KܽSc�;Vi耠�n�R�=3,����}b^s��K��	�14�R�"8��r���X{Ԩ�7�fE��в��(m���Cn�˴����u�b�
�}�)�����ԒX�,�U��׆��O+iv����XWr�V��*�m��$ʺ�V�o��PY�ئ"tWi!gG���pj��ʌ�{^u}�12�Q�TV�1o&mr���W��G@$��Bw:T��>����s��K��b5�`G�2Qn��5�9��K	l�5j���̟AQNp��4��AqE����T�§ ��J�v%�Z���
�Lh���hq��%.0�0��o��,Pm��'ow
���WQ��\/z�7�wB�q���Bh��|tc��K:{ft�ޭ3lWX{�ι4F��-�rև��m^��,�}X��f���43�gX��ݫM��5��	0�(�ľ��襫��{S��(b�tʡM1���n7~�:�UuO$v�����VȻ������ktsRN\u�l)���}��5�>�JN�N�:��Nu��=�*�K���qf���E�C\�kX�DVq�fi�����N�(D7>�)ɼ�چ�4�K��b�j��'RQ�]����;�Ϊ*[O/?��������{�mm�-8pk�?�H�|V5�V��ٮ!$�F��y�i�$��ۿz�S֍��$��kܩ��6m��+�]9�}�w�9즼��\��n�.��{e_mǙrٟ>���[xze����e�yӎ̦Li!�_R{��6���i�EP� ��|�*G�SãP��IU�����l\�T���E=�0�Y��5�X�^��F�̫��޹w%ǧp�w
��6�^���h3J>VH�[j0M
��嚢dh"�%���<�D+3;3������!+!5�o'0g����ʵ�/�V�&{f��00.hs	�p���r��e�~kcUj	]�cx�z)���,����Ƒ�ݮ����;he�����\�$���Wm�7ҙ���Uf����F�J�ˑd�29��Vܺ܋E
�V��؄�{��0�6FKا|N�yTԽ}[�� !�q�����c�Vre��1�p�й��ݷ�wMܺ���ӂ0��{r>C�dկkh3G�j{t�2�6�o7��E'��b���J��x|su���z�lFZ˴��xm��Yj�;�'Gµ��]�N��d����0*��J�d,ԣ��{�7�w��'��I*I$�I$�$�I$Rd�I$�I�-��Y�cz�� ���甏��%
�܆���]�Rܖ���FQ������K���[{��:�Gu���f�2��dC�{x\K���W+��oGd܆�Gl+�f��/��?�-���1Պ��(�q��P��:�_N<uo[���#���]a��,��1��%^��lown�T嘛�oO`[�o>Ht�nh��(%�6,Нŧwb�jщc����^j^���oH�{�H���7ٱ�ʝ��Xr�QE;��ric:�ud�ԹbJ�� �+���$�����|[�L���~�\�Kٛκ)���7���oUrȴ�g.�fWr��bkt��:;+e���ĩo2]r&r��Z`���N�r��/�O ӡ�@j�Υ� qv'w��nD!ƻ���SD�'��g&Q���e���D�Z{,o0`�����e��ڕp�D^�!qb����!&�E���Go�,]O6d�������U��L�U�h˗��$�z&v"��vst�{.в��ʹ6=R�Y6�ɳ�MZ�Fe���$��T�j����W�zI#�I$�\�H  IrI$�I$�I�I)|i&�Z�Y��}�n@a�����lQ�����GJ��pg%8+���}�-<+	��l�ݳ}R���+%v��Uj����R����lխ�36.�3z�1��QՎ��\R����� W^[�)�Y��J"L��ͪD��q�WC��A�n�^ÿ.�#�X�����C�/q�?<n���!,*C���jd��N��G�s,�x�vIՋ���;��s�b>G��8޶��\�3-&&��6��@�w�T	��Vں,�v��}����[:�嗊�9`4V��A}2oV�[��(��ޣn�f�\sv�|�K;����0�V��p�����@潷��eE�9ۢu���8^�L��U;����	���V�r�F''�*gJѷ�%�n���_��vKг;�*Iz�s9sP��ќ��w��*Z�}�ī
���fK�{�c�f��k�9�1�ԥwWh�;=��G�����eU)J�]�<�n�W\�U'{�s�
�A�r���<Z�-� T�WX�*�u�ō�A���ձ��G톦�2S����>-*�v�X�͑Mޜ\�"�YTx�{-�t���f��������H�GP��g/n'1��8%N<��ؼоy.譑����v�t�b�s�4%"Z�k�7�,�!�Mt�q�:�n7�p�x��O�&_��0�N����Tü����8�^��|,����d>�M�2_]����[Z�-�e��2C݆�q��{+����Z��6�>F�՝�Q�i]D�v�A�ۤ�p����5����M�0�,���K��; k��G�����d}n]�zj�*�7����k��t�gV�l�k%8�D��7X�x�z2D��T��x{�oQ�p؎�7�R�S�>{�0H��^I;�e�:]k��
�,�<����J�N�r.�BիH��Rb��Kγ̰^M��}m�B���sy�Q�_0%�ig%Y��/\�u҇s���Һ����U�p��+&)Z�s�]�Z����A�#��+)����a�5w��rAa�1qj����
�&��J�f�]|ぬ����xKīV8��J�W�j�Ws�}SwG\9I���u�#��凜�N���\hbL�H�(�_Q9��Y��Pw(�/^�<mke�3I!s��Xx��H��G������фK�oeZ���J3���MVGՠ�X,��t��1��Ź%"�:<�*^��܁�"�a蚳��r�R�!�nn��u�3�A��v[+���}��˼:��g��Շ�ZXr��.|�9psk:J�}7��$"�Fn"��R��.b�:6��he�i��`�v��H���.��ULN�K��CCZX�x*�!��!�v�^�qƃ�9Z�`X2_��+�RH]X�ё�-��ĭ��*��y�ͤ�:$���W���L]M���ja)�4���D�ۮڹM�U���a�����|{��r0������1�H����z�Da�)��Mk��r���4H�7�st3��ƲZ�7oGF*I�y���\B��Ćq�n̻�]D�xQ�B�c�̫lT#J�'�W;�5Pg#�.��)���;N��]a.͋�gS��<3��ھc�9*�;#IޡA��b�>m�Gi�_N�-Z��BJ����h%�_wX�\t���=6�-	�3�ԡ�58���#���5�w8��Y��˝��q�L�c��m�������:��������a2��.k��^P5�f������L��S"�8��U<�[�:�%S����2��gŘ�t-��b;SJʒ�D�Z�W��ɶoE*�G�v��ֵ�u
�Ri5��Xͧ*��f-y 9\zʳ��B�u�L7��roI�m}z:<.VPX<hcX���x�jz� �5Mq�m��ЗCy�����kM���}�f���nS�B�<�@��;�B�����L;�L9a�]��5
�Ѥ��b͉�(ӂ��Tl:���jc�+c�޺�7O��R�ñ*okoJeX=�E=�r�4����n$�PX\h�HJf��IJԾ�S1\�WG�֕`�׉\�B��]��s-�S&��iV��۽x6�]��)�E�!�#y��Ev����S��^;�1M��M���ʡ�fu��j��x"�20J�7���R�S՟�� 䝫�wZVb���]s��:��/���j�]nV�\کS�����:nX�NZ�W*@&;�U��V>�q�+S5T��Ω�v�N�:^���@*�	ܹ]]���x�c�wA�Nxi^�-6jaoi�7��It;�g4!�a전���J�XyY�uƴaJ��Z7�9텴�q��2��v7�B_M-��q���˺�DI��Td}��ݞ�w��Z2�e����\{:���fvp� �hֽg�^Ӣ���+R�YRZiB#!���u��B�Н��סj`ͩ��wCܼx4�����C4'z*q
�ͼ�[��b�!�;\z�����9���y������r<�m22'5]wlA(��\]�@Pڹg�/��wQ9vs�+�3��u+[�LZ�+�Pw�r�"��F�=�*r6�r�jZOT���ӈur(#mi{N�.8���8���in�VU�婍�Ⱦ����:�ጰ4e$Fc�[,c�3�v��J�W��C����# z���N!b͙w��l���m��s�&*;���S&@��{�DF�V��d�V�b���#J��5]sb�0"-q�.��V�)'i�RU�:v��	K�a���rWIy�Y)h@��/��r��im�!DpO!U�aPF�X���Q��D�IJ	��6L����@B���d[LM����G��l�%�t�*Wǎ�ꫫ�2p��z��/��-m�"��0�9��r��ˬ�'[�W�1�S�b���GUp+s��q��R,h���Q��'{�ʕ���ΰeM|�U��0#���1B�sxw"�����/\�q�Y�����9�s�
�+d�
;Ҵ��9��
�R���w�����*��c!O�m�w�#G���^��b�UYo&�	n�L��C15ҷ)菭}l=�"q�9yC!��i葋J�3 yZ�����*�4����t�g��ЇmJ�F����7W��#S�WD`���O��5ogo&��0�ؕЫZo��nNQ.���}��t#�q3ne�2�*"	��e*׋���E��{w��$�^=�����ˢ2�����*��T� =�E�� mʻT�d����庫��8N�L�ڹ뭙}c�s3j]�wW]b��w*�v�pL�0n�
�E*�;s�ށV1:�n��/�CCEp��2��P!Z�q���a���<D'���-�5��S;v��8�\��Y�v3b�.��jOC7	�#���1̳M��0�Gi����Uv�t`7Y�Bۃ:�����I��,t7��O�E\&3�S$�WXd`zd�
��Aq�M#��ʵ�Z����%<�5�+����ꏚ}N���"f���q��L���v8���QZe͉�h����1�v���s�6�݄:9/&�y�G���T��#���
q�q��d��A�/�����M�ut%G��#m�� �oo��t&r����h2{�fKȔ�q��xsZ���ff>9�鴊�IS�����A^��#���Ǯ�q�$ō��$�U�D���p�+U]�=����;$pM�CE����Y�]X!T
1�%�t2�&AK�X��
.�'fO��u�99F���{�=�̩ը�t�+S]��v,S��0��U��f����5��bW5�t���ݔW[R�fB���Mk���_7�z}`4�T��Vng^�T��Tt �sF��l���S��M��"sz,�6��NFͧ8��\��s0��hz���KH�A��e,�p���h/�u��Gn�+��]5f@vX��j�zV݃��5c ��gF૶���]rl��gc��.�Z*��5gNx�B���cҁ��0����ł��ue[R:��H
�v�I*Xͩبr�vS63�C�*��ӮE/n�Yy�@���#�5զ����2�H(,n��L9��-�d���JҐ�J��tK��0]��G�+��OU��s�e/U�<��버(U�[
��x�b�On彃���(�Y*R��l�S]��NpY7X���~E��
�0���h�[B$�','O����W<U���44��" ��nS�.
׮����*K\��$��n�܁G�He@ef�.��|fn���	�駮����n��/�����יն�X�ȋ��Դw�=�N��X�W��B��t�(ά�N�i�e�e&fc�{��<��l�N�{0�����u��W�^ym��k����e���lW8)MOT�je�u�#� n*��E[.X5���	�!=��̷NC%#�X9;���5ʭ�BT��9Yo��`�5vm�]�v_,�y�xoh��N���0!,�}���;*�{l�B�XHnn]JgH<V�\7�� ']M�,�U�L���X�N�s���G�2�����#n7����'7u�/�pJኬ�Z��ׁ� }P��Z��M���%%�����3p�^K-]�u�����l�c����/l�$��qϺ����`x0`�fzS�a���	���c]�ت��*A�G�Ɣ؁�3zDJWx+�Ds4��o�\����93Ӟu[0���Ҏ��B�Z&޴��y�f�7b�](Z�f�yG�r̺�yd˪��LF�UPh���bz�	�EF�A�j���������]�g��z��=#�J$�Z��k�/��{�|}O��P�
����D����zg�V��$�:�G�2���ƜB�v��$���y{$* ��k9G�T�s�Գ½V��QY���*/ƬH��*M=�"��d��3۔G�(�Ԩ獖�&yW�*�<��^Z	EDTJ�U�ˆ�)�YEJ���$�!yy^EE�//*�E$�PI�[m�7(����)��Vp�DP�Iu�)zw ���f3"�Ȩ��.�^Y��r��QRe��%��=�U�Z�E�;�~=�>�V�ȕ@T�s8�,�9VcԻ��k=P��QΝ�.Y4aXR�����}�xF ����������)/�� ju�V�N�q���@���X��V�̧���/��a�4l�N�{w�ڽ��܏G������r��8��2��7�'�\A2�
��㍈s�����£C֞���=�4�=�t`�YS�.�賶�8�Apl+9/���#z�l0�}�$e͌u�\��Y��𽒭�B܎��Ec����1Ԥs���^�=���cw�+�F�ʟ���4��!ގ�Q5��L�+�:b�8l#%��|H
�o���L�ѯ�>:�
0q���]_&���v.�O(oD��tݩ��;��b�����c�M�6{~������A뾋Jwj,�ۻ��ht�@��r�J��|�3]Ć���b���p�;����˫�f�ݎ���m���:8s���XǪ�j�+���ToN�Zg�r�c\��ݙQYn܎Q�%wjH,��r��� �
)9�*1�sӖ+�j��W6�n`Q���tzn_33�+hE�"0���7o�L�|%�|�S���b�_p�t\�sv-�� Җ�ѐf�;(�Î8&	�9իӾ���t��>2�m�<�������uA��}�B���cM}q]�fwl�8=%��qO�h2���v��o$���^���7:�2WuL�B��-n%�N+�!3_��-���֜YD�jv�1G!?�jL.b�@�J�꜕�
>>��ƽ�1d��
]���!ñ��u������Z��w�5�泋�i��x�F���s>�Q}c㻬F����&�~���v�+�����[1��@�/D� ^����Tlw[!=��M�,oV�e��3��$`�}�K��N�����L�-���_����SvgD��W��V;�JA۞ҵv��*�I�!�00AT��m[�D�Q�pŕ�?}�gU��}ᴋ��B|�By�ѓ'�����}ӌ��F�&-�Qzk��ޖ�v�M����6_Vn�pA�4��Ku�A�=z�ۡ�ĞS_ß�7�����;�_��w�R��	Y�^�b�����W�!��՝����ŵ�����{��$!g���1"�yo<�+˾�ɫn�T=��������vL�̖q���x��⑅(�ko��И¨�_�і��	]1�/���䱊��U3�����/��,�	l�-:����<�n��xv��e��@�2����Z�����FYٷ��O-��Ѱ�p���Ë�D�h��#�.i��n�oennT�ܢ:9R�f�J��\Sl��P�J�=4�٤�������J���S�oN2K�H3�Ծ�9����|_�{b�s�"��X+��,ĳY׹�o�jKw��E�	��S�ױOQ���겨v���q�Q��]P6���5-�N��r�Vf�q�O6��E���չ�17��2��V�a:�SVFҗ�H��:��d�"�Q�bk9+k_Mf�<�^Ŏ���ec.\�rz{`�t?��=��GiL�c���� �~�� ����D�ޡ�5����PH��iq� ���fn��{PB�+b�I��2O�����x]�*���㥕J97���{���2$]�UD�M���Ȭ�9�=��ޖ �:�̆�n	b�{�ԶZ�w����'�2�)Jm/]�����6�܎�I�ڰ�cu�d�����6wr�M�H`U5��{:�	�k��s
-�ӸV�4�Lx1u���Vm��&ZJ�<ji���76���XP
���5���0��u�����+��FA��E�R�]'������]2�*2���eQ¢ԟ瑲!��.܍��d��w�r�5�$��J<6O��*4ʍ�P]�A7!2E��5�K�׹��s2cʇn��]��D�'��X��ӷ��g�0Fz�eY���ڝX��Kj��h�yex���UMK�����^�����	���6�:�,oa'�6��mg�]�ۊb�OqBi>�.ކg���w��Q�����x�X�b"���n�Q�1P�S��Ǖ��,�/B�D�N�H~s����5l���B]�&��R�tu=��g�tH'DY]wY���KƇz��.\75b;��b3��Vߏ~��Vt=4H�T�n5� �Rެ���އZ$�JGsj=AG�9�f��R�4R�v�<ڧ��Bz�C�c�0h0VS��=�}�t�������[5��'�	.�q��V�m7��Y�|A�K��V��N���x��ɻz�h�sWSѲ{w�{'\5�D��.(kQ~��9�q#���ةrt�������y�i�ܔn��Q�������>�����J�V���9�1�P��z��M�C�fJ�ȋFu��yթ�����w?	��W�Pt ����8=Zo&c���S���v,ո�����ʵoAݷ>ᤋ��;�����&�ʜu���w;o.�Up[d.|�O�����Q�\8��NQ�Y����
ܷC*E'oekd,�9�H�p��Mc�U��^�����	�[�kv�K�\ܗp���;���ɕ4J���(f(i����4�y(q7��y%���)�݈w(���Yn�nd�n���[Sϯ);w�囯�����Z4#�'����.͚�q�#�ne�9�\�_�_t!Z�;x�wǓ՗�I�F^Ɯ5C��$(v)`�>oc���]�� `S,�ZB��Of��*��ι��')T!�b�ig���w3�<�7'��*�u��)�^��u�h'�t�u� �Uu�k����E"�}	�[���
�Kyp�x_?>zș����J�׳I�ѭ�yH�� ��>ܹ4�M��Y!��F'951�m�;��m�kr!��^��r�5��*;���X5kT۱G^"������,�������Z��iV8ڻ��4�S R����te�5jT#q[ ���,
��zYC)޽�N�k&վ�k=dQY�Fۣg�ۭ0D�Q33p�,�yu�rj́��(�ݛ�[&^gq���^�Ӧ�k����Z������9K4�P�7����.%S_d����Ĉ��^�㈮t�F�UF�1H�5K��A'�u<�µ���)>X*续�j�ϊ�,��w T���/S�I���r�؊�P:H��ٵ�z��yCU.�Ӻ�UPD!�=��(�qK���8�oCb� 5�#���T�+�`񸨎4��*�c;��cOFeu{>pm����\�{�ԅ�-f���w6�C�y��թ�17���2��Wt�'Ȣ�Os��ڸ'�r�j*(���J�V��m�}�ߩ�w���O㓠� ׶�C���$=�U����=�Z�.�I������9�!�:�9���2�Չv��%
���.����a��,u$[���q <�N�i�=[�3���ق������WfS� Rf,jf�b2�W��T'v�\l}�q�U�b� pp�Soy�@�~Φ�ޔ�ֽ�{PBfP�&O�����[�<ր�����e��&���`5N�(�fB��rU�S�1]�CS	��~�"��5�߬J6�(�Kކ�Fw����8�Ⱦg�B��ꥎU�3�:3u6彬�O28NIZ�Y�I����ñH�m�̷|[Qj/k�ɁS��"���am��%�-=�^��+v���x,�����z ��צ������/�Z�,�g��d��f�qD��lk�B,x���N��m��C����X=Y���x`�=X(���7ΤX�Z�P^J{�t��Ϻ�ë��F���S}�O%��Hݪ��T�zu
xx���Ǐ���V��TR������̵��p�2c�r�|e����q-]�]/pc������6{ܶ�A$���NC���Y��l��=t3�oc��L����5uRk -g2���%��#�L�`��'C�EY+l��S����TU�zZz�.�a��f�
�r[���QBSU��Y�ۚ�� C��$��ٲ�+bͫ�mD�m01��׌��eX��v��n1�cs�k�Wuk�>͝2F���{YW������}m;�&\-{�7�a�:��il�RJй����7�+�N�x�Wɵ�z��+$/��A�f�foQV���Yg�z��ߥ�T�7���;���8����u"�nO<��\Ũ	��f;n죱YB��Ė01��H0�' I\��+o��CG�iP;E����y7����k����k?f�gzzMܑ4��c��
� X�N��s�}���n��r�TW�/��깭!;Y�Ɏ���լ3�+I���K��5�7w1 ���=�d6��X�y���jM�W+��	�\[e%NC/�+ܕ��Z�fp3��5q�n)���c�y.��;�]�qŤb�����؁��*�N�]�m�����vU�96����"oOgX�|%ؕ���%q�2���1����Wܶ'C0Jdt��]UD�ż�|ʹԁ�(�'X7�Ŵ�7�n��u�w]�1ӎ����Z�YDY����yN��֝��M���N�]^��ֵx���n�f���B�c�N��[�S�'��JkYI�b�B�]�®]t�&����&$���IF�)�A:4��˥��^$M�)��u�\��"	zl1:�on��t�5���q�����VRHs�M���(������=v��A��Yy|���%��Zdl�é�ʻ�h��3�V�=]�и�2��٭�`����Ss���8�U�zK�Uw!Ӽ���>����Zd:j'��oo��W*�y��I��������/�����HG����K���vc�k�s�/2:��
��|v�	q��yb�ݑ
�z�d�-&��+eo�sp]&��h���N�x��5!������w��Y��5B�})�o�>$��]����TX�$��їՒ�:�i}.�F��s�õ}��
����T�.W:En;�3�bv�r�D
�A��kI���[J��탫��v U��K/^T�l�iT�7�I♐��i�=�]�\Uv�`q���.pn����w�!Ym�du�2�s�l��KÖ_8��n��f��Ӵ����+�'��ٸNw�n�Գ)���g7+C��6q�R�t�v�abÏ]E�X<�JÎ�*������)5t^���ž]y�Tt�mz�㸰eJ⍛2AO��6������&�\�xy����@��3�"��AH��Zn�W0;��l��S�݆�ked�GV�����X9�����\�SݣN,rΎ�/����nd��۳]W�)�h��WG�wڹ�/r�g���J�$��&DQ�!���o���h�Q�4��B����ZT"*���EE�m�QP^��h�2H�OD�#��x�)0(���DE^tm(򈼈��]%���+2(��!W�*.ФЫ������UUQ9y�-1"h.QUyPUsӐ�]t�9�tB֛�#�È%3f��M�*�����ʠ�UJ*�U\�T���B�L�+��bu��ȴ�j\QE]
�
����Q\3���^y�HS�f.�&��Q�M�@�vi�*�Tfv[DU��*�"���++UqUD�H�Xf����00�C�,�Jb��2Y��D�jQ�5�j�6�Qja�V����������Q~ V.ddY��)79�ӶM����S��$p�fx�B/L7��|TOUeu���zxk7�w�?�	O���
�VUZ�[��v�%�6�-c��}��#~_f�^W.�&�!�.oo�׹g/�G��nv�8EB�|���}?l>�t��Q.���`0e��˓���\�Dtt�#�P�9"-�5���żߨ1���K�s��	� ��&L��� ����paYӍm������9C-����nf������W�K?\�_��[�ic8�n���|���������FqGu����5��6�d���g5'��/+$�}X��]�ڼ���ϘK�a^c�����寧 ���ۊ[��V�i윷.��܆�^������U��ߑ�UxEE}��b����Zwr��"��KAy��ؔ���bݲ���:��І^���jƥ�\UpA���$����:��;�h�Z�&L�hp�I�(<���5�&��99M78�\6���~��0��x`�U2N�Fd��-��XP>ߜ\F�������;�d$}�DQ��*����U�oM�"�LԔ`�*�)��rx�3>ʽ��{S�q��-�O��������,�s��z����s�|S?�y���Xw֋�̻ME��|f�۪�~m9�Ւ����9�[�[�^���~_LlT�n����_���߀3>ӯ�����o!��`S=~���U%ˍ�_L|V�%�ܗ�l�Ww��n�m)�YU�/���TG� ��D�;+�V�}��<�aKNǚ�={ﳰ�w	+�8D!���Բ��gّVf�l��|�/�g�T��χ��Ζ61��v��g�ɮo�Jd�X�w}�e5�v�� �[�~5�~+tU�ǳ0�/OW�p����:)��q�?\�)Ԧ�xYc�����6r�m^3� ��ݠ�G�4"�s�Y��tL��8:j"��jl��s3w߫�`+~t3��U~��;wu1�u�C���.��kiL���ۈ���Y��?NkQ���l��\�Ǝ"�Ų
q�6��hX�d2�lZ���Я�'�)���/}8V�dH��4I���˺�5]7Bl�������}q��������q���������	r�,�e1Zu�*/_:�)��w<���,����"D�d�����e��-Q~Z��EW()��]�� �ʙ�Y�Þ��%	���8'�`֯	szX)t�z�m��b�%�F��Ŭ��~���2DB��(����X����[��{�*���q�}�""v0{���s_��;��1O`ΩM����]��c#}XIz���@��4
�j�f�4�Vv��Y��[ȞQS�u��3�dëz��$�n�0D袃�B���d)���a�{3U��B���[�Z!���t�;����9	O�BH��|W1�Z~�OZQ�}:�*2%?�gMF�O�zj�����z�i��{j�q�O_��j��O��˯�:�}����;��"�N�iWD����p������?l��Օw��]X��K��Fo����ΪyS�T��6O��Yw��V+� m%�6�����+���ee#�|������j��Q�%�GH����Oe�U��#'�^8�C�k�]����7���nom��0`��*xx=ʰ���.-��p^G��y]{�7>����O�&}
c���y3|�ncO5��{ǭGc� ��!�^/�c4.`v��� [y�ؾ�@q���A�j{@�l�ق�!�t2�r���}l��3m�zﻌW��-�Rb+�ߔ'`7�ch!�4��Ȼ�&й��=O�c�Qؽ�@w�YE֨r��������PC�j�ޞ>����E�� ~���jV(ͽ.����Ѽj8}�Y��|�ؓ�z�i��Ώ�wsI�P�l�tݡzo�!��5*J��>9-�\��)�P�6u��i�a��nnk;�LVw��}�f�b
{�<��9�C5Ob��F�hM�l^��wE�\��_Dި��GдW�h�_Ay}���/���_��cƢ�.�C�P�%�{�%�P�TVנqD/T�HY�`H����轁"�4 �5��w�1���k{����o<��^+���3�{�9�Z��/f�^ʖ�cP���S0�_C�p=@�	��;Ш���9����wη�s8��. �5AD�(���0n�C�[ㅕ��^E�WUk#�%ʠ�j Y�!���`���aob�/��z��������@̼E�*!�"��)ȍ���	w[���� b.�RH�acw�:�\�Yp$I�w�+r��g[�k�;�uZ��B���/��jE��h;�}����홨-��t'b;�m����ν1�3��0z>��~�T	�{����^��nX�w��M�yb��}3�Pv���v#��f�%n�q�ӕ��ܣ�ƻ�v�̿E�9�w6P�ކ�H9K"����;���^�Ҡ���R������j-Br#ʳ�w��ә��8>��G��GѬG��'��(@�^ނE}<Ŗ��9G"T^B���/b��^�"qI�Q��h��ܪ�����*�3���_� �������/�퐼\���S�1��A��j���J�ȅҩ{q}z0^�S���v������u���W��d(�tX+�7ơ��q���=���S��6�^�����(��S��5�V?���Ә�8Wl,q�W���f����E�7���f7�܁�����\�w٥$�Rؠ	D�i}Ω�@��O{d���<���Sh/ �7�-Ey.v�E����q~�Ncھ��o:����V�\Cؠy�m10n��}��V�Q3�=*gt�`H&��!躅D��qGqf��Wz����;;3W�(�z��=럝z=�����[�C�{�zDyq��K�o�5@�Z�qGb�#��~?}�#�Y�{�fץw�u� E�����.9K&"�9H�f! r z�	؍�ј^#�85@�.�K����ؗ=G�`\׫�֥g��3�w|�c/0�����z.�甆��-�c7�ʂ��#�脂���P��ٽ%���\�.`z�.�����L��~��������B"�̏��7�;qՎ��]�A�)Am��^�.⇒��Jb>�^��W0�z'��1�p�J�jo8�{v��@�@�f��^B�|�;�������rǢ�j#�z݂�.R�+�{^��!�2#��)��!���ts�������9�w\��o ^cx�"�o]����c4<�轅G�@���^D��d=3�ye{5�� �@�)�L����-}j�γ�s��¢7��B�/!{Qh/`n6�؁��Rr/aQ��OE�Of��_@�)����`57�
W�0o���w��N۹�9�{3ȝ��{���A�	�T'`n/���Z���/A��ɋRf.��"�/�`gT�`6oF�����[�;i��`ݩVt�ٷXY��O;<�v����F=+[��f�,te@�'@�����r�Z�2N�͸͌���ƳëLˏ}�^I������YR�8�]�ZҾ��7^���`nj�}d}E�i$WP�j \�>�P{A�R<��Q�^C8�q� �T��&
��P=����ψ��r��k�C�������Ǽ&v��F��H�7��P�`X��@w����f���^C.Yо�d�R��|L�v�{��k\�s�1-�q��O�;��c��;�^��M��-ܽ�A{�Ŗ��u�5Ш�-@r'b�+y�w��V��󞽯�u0�MUy�	&"��>��r@�j�ah'"�!h9�#��=�������5���%j����3�s��v�j-���.���#ȅ�Rf�9BI� �``�خo5b�{��Y*`��$DFO��-2��ϯ	�����GO���гa��FɺYsڇ�^���;�nb�0^��Spb���r�$(1���	��Mc�B��3{�W��}��J�����R�����,^"n��z �_L@6�K�B�NE-zN�y��1�o�� �n��4���<�?\�L��ށ1f�ϼ�ǽgP}p��9Bv&��X��ߘ��(��q3�7��=*��<��b��k�Ž���9{xA�	/���(�	 -���F���9�躋�����]�-��b�,��=@�f!z�����=U\�}���mn����Gax��n��PI�T!ؖ��⸎5�=���Sud=SPrz���/a{�^J���g�D\��.�*��۝��0�s6�����L��1�_j���`�4uF�3�O�%�G^]����{|��T�^}��W3jF5�n�٣7�B�Z?������G�̖�36tIo!d�g�^%��I�-���D~��s�O�b��R��"���P�ؾ��T�"v'!�Zg}���#�ޱ�.���)�������6Ƿ�{��ߑ�C�)dP/�-�S؁!m�z����v/�8�&��/�PƩD�NC��5�X�_f��K��~ݨ������o�V>W��~�.⽗-{
[t��@~�~ж��Ԩ��z��h<���B�5�w��9�1�w��o/ʭ^{5�k:���19�LU!؏�r�٘�9@���@�	"f�Br`�5*(v�'�x��Rr�Q�=�n�Ƶ����q�1����4`7�����������"����2����mQ��$K�	���bԮ�v>�5Rl��W���۷m!h�7X�0U`��������zn#h��,��5���1(d@���T	���
�؄��}uN���}��3C��1�x�|"��MF��� �.b�q}�RDL�ͩDm�X��Źe�;�-� �
�����#����'�^�v~e����S2�K �5��Ȼ�mH�/cw��q�S9��^MD�)��Y��{�^Cu��%Z�^;|c�oٝ�n���7{-B��u[�Pw�rԏb�Z]�#�%�A�/"]�	&b�qO"��������of��}�K^����s��	}�TE�	;�}Qo�Y�9zZ�A}E��Z��_KK�j����'���?OM��_��n�!�H�N��jnq��j9��sܨm�j��K���v�Ux��'d�'��uw���XO�/���C�º�#����2��u��o���K��eh�M�5�X�D�l�)_�9�w��޹��׿��TK@;�(�]@���%@�]E�(N��[�ŋ�{�����Ⱦ�!w��d����z4�>�W��b�o|�W' ��Hb�\1^��G H�B�wc�{D=��s��'��/C������ԼW�wau�>�/�n��g���|�S]MG١KC1��rn��/�1�0=��	2o6;Ш�Π��P3� �[f��Ǽ�"=�+2�����WN=3�>�l�D{5�9�|j��ף1��\��]��fh0;���1ި�^ ;{�!���-U�ۚ�1�c;�1:� ���)|P�TG����O���F�hM�mzKE�	�s�}z�w�.r�B�\Ƕ��-͕�b��9�s��t�\�}�X�^Eިtb�1-��_D.r����o@��^������[j��{E��}����*P�$��s���1�Gѕ
}��~�Ǣ�����r���/ ���쩨�@w�LB�}����/���Zu����;�9���׹�ۡȺ�D=���ơ�4!�����&���)^�Gp$]EyV�:�\�F��Hnb������+�q�s�ͺTV�1D�@��(7�����>���c4� 7��b�S[���� b.�RH�am���	������{[�VE�	�R����E{p�NB�^N��^@o���_f�=^�;հ
m�!w�2� �������tǮ ���+�C&��h�הe[��>AP�}���cY�8��.��gs9�[����\��/NR
��}Iq%�EG2��2!z6���D��.���|'HT�4QJF�_��O�3�������5���mY���ɚ��	�B������"t�I༬� ��6H���3ǲ�~��X��W��B��?��j�ɹ��K�{���}}�ۆ�2g)unj�y�ýv�)�ض�G���Hdr�6A�����J���Ӽ�)蹝/�O:�9������<Ɛ��-s>�U�s%�2�C�G:�B��{��g%�ٿ���)�m-���ڲa��U���QuxD�#���F�ᨷރ;F�[���a�%5^�t����9�9<x�|�׃��=��3�d�|ǧ�^`e��Ak��M^�G2/_�q�%��^׈Vg<-���>�?e}�UfU�C�g�d����̎.h;C�U�oSv0�k'�ސ�����c��P��Bz좙K�v��W�t�@���٥��n�**SK���X�[�$����CK-����w��Hqr{\M��C]�j�3r���$.������a��´n�Nʙ�Žy�����.D,���U3fZ��o�#X����a�,�v(m�p*$��Pe��Z�� T�z/u�K����ջt�������ww{3��.�E�2�]�˛N�w��C.�J�8�˾;�9G/i����}�y:F���1��q@�]���\�9]��{��pg�5W�ޜ���A���.	VsjE�s�r��C��AZ�&�Zu���X��\v�K�1���Z�������J2�FꝣF�&��zV���"�'���/z�)�o���.�->�*�N�;�t��|,��clc��]�+w���u�ŎĲ��L�:w��m��#n�S>�RJ����O=y,��ٺ���Ylo=� ��d43��:��sbz0��K�q�GAӧ
��f��"�8ٱ�is��+M<+[n��Z��\�E�/�jvZ2m\V~Tt�RIj_�㟴P)����������(���9�ԃ�;��3e��=Iu��ޙ�_pr�]ǲZrt�w�_ґ=�V�.���7f��3�u��ev�P�mG�N��DX3zY_v�;v�҇,X�T��Yʧ�U�����k��X:�}-�ap��q�/Q����9�.O"�>���l���Jq���/,#]���|8W���4�G����f�(5Pjg�][n1h��8*a�mX.]b�h��	R��R���,μ�.�ڻ�����#}#Hm�fq���N��3ڪ��V�y[ɰ���%�Pܹ�����N���[����փ`��.[f���<�Xp�������Io�GʝvueS��|L����0�T[ͮ1.S��gl�=�}�f��f-�0K��a�[*�ң��:B��C�3U�	� �b<lu��ԧG�:�N�2��9Pgk�Զ]��o�a��G�ޟ\ۆ@fw�:)ʺW
��ܗ��m"�ݒ_�@\au�͈��d91���û���x�Ut�y��P��3+C��Y�f=r��3�8��q����H�T(���H�V��~횇�tm�:�Ɯ�Ffy2��﷽痽K,��vM6�J��QA�ep��mJT�ۥ2a����ϐ[�>0K��T��H:r��!V!ַfz�W��K�ږ��==�]s����f�[l�7<B0�@�75��
ƱR�*#�%kb3*f�mvv���f�fj�3̌�R��j�3*����Ĥ�ɢѱ
(�]���TRLhL��"<�r:��y4d*q$*�ʪ�����
+�UyF��Qu
��*�hU�rerH��Q�#Ur��\ҙ�/� �jq�y$�n�[CR/*���vs����[Z�s	F��)��)J֤sӗ9-L�Q�^�fl�b��+�7������c��}n�Yt����|F�Ӛ�/��`�N��u���p����m�����uWu_}�G|�����[=��׽GO�~�����k��;-}}n^�i��[��{��&���/�x�܋�^
yOo�g�W
�T�}eȌ-^$������6t�:䭬��Dp���-L��:��js@���wV��js,o'�Q�D�)P"KQ��"�HeM}Bk̽[j߯+Ȟ��\���
5&l�bJWPo/�+F���ve8��9�������8D!�=�����kY|��"�k�5xh1��T/���Й��>��u�596oQoiL�JtD�E1gbe¶�6�2�,GR:T`,o���K���pc=��aM��!8���|�J۵Ƽ���uΧ�#������n���dd]{�,[�@ҝ�Ύ�9�h�N�����'�Q�!$pv#����q� ���D'[~�H;{P�&�37n�qH����O/�#���>��h;��߫.�@V��7���d3oЧ{_o��EE/
�)�� �6$�gR�Ӆ荶D����	��mY�h�@qǔ�E�J:˘ǋǄ>����Y���S��S_���A�yP0:�\j�B��6���=������f^e^w�f]
��`�o��iEVroq��+��N���-�[V����8�F* jw�\�i`���e��ɚ��^m���Gd��Us��9��t��k�\횹/wO1�����sG�n�?ll�{����o9�K���q��Lpz�O�J�,T��b�h�cN۳˛���iΫ��⽴�N���G�/!\��a�
u��5�.���!1�ok)VK}ڗ.�|ƯG�^�'��'=�݈�v�^�5�������r �����?��#,�>W \V���b��؉�e0[P�?�U��뺪���G��.w���Kl�|�+2(�f�tJ���(q6dU˽�z�����.܁o���nvX��^o�!&�C��g]�<�����L��uI�/�1�e�uWI�7��I�a�n�GhR`�z��]e�A�VB�ur�Nn���+f\�f�&����>�G�F�Ӯw<*(�]�-<�L��}�&���i�[�<0��%��{���H������O�W1�Ev'6���Y�\	���2�K���v��׻�D�4���]����%/%1\�D�m<+k3u��0_J�J��'��'{�����sm$Q�V;��7���_�![R��
/�򊁿(��w;~��O���+1��Z�-+g^;f�\ֶ��)a��M�/��v>�Y���0j2"�+u`2�rh�W4�ؤ�B������ٛ��{��� �U��gMD%f�.��]&�\�z"?O����ޠW/�ϳ2���L��z��ǨTnO��3�Y;�7��3�[�V"��}vH�������M�1f���ZRn2&WLO�.�*�TU�C�̌g/�yu�0�����L��%��\LdTO��-�,�b~� pUjr�����<����z�Q�E������sxgtQH,C�f��c����|nb��q酁ɶ��P@D����m�[��Kw�]�<
�6	�2��A��/�j�ٗ�Qx�Z'���G+ ���r�Ȳ��$ק�j��?
��l:������ㆨ�#��x�[Fi�˗�����K����񴫂�%[�q�=�n�z��3�P�.��nB��R��P�Ph�Jc-�*�)��NJy�L���ڲ@�L�}���3e�=�R[�U��Ǻ��0�X��Xn�RV��}����#ޙ��{�s��϶A�luͻީ"���2֘���� y�/M���u�x���ÙX���
*گd��H�$���^�=�Ci�;�x��̞|�'��f6�dY�d�G!Ů1���N��jB��y4��U��2]�Η���_���G���܆�]4���oB�:^���>@J�E@���c�)g�ph��۶������j�֬i�3�l|�|��	�<QE$7ڍ�j�0b�KWDE1��F�)b󮉉�žO��$N�Ψז�����j�k8�5_�^�B�v��)pҫ�LW)p�Iw]ޖ��d��J;b^�y���
�L˱��Zk��N�d��)9��/�h�ۮ>��mU�e6�d��p�v7���V�s�G�Y���:���LN�BU�A{slQ�R�UW�꾩��{�������ȿ�����	8+�5�+�8D.y�>�.��]��ꩩqO�p��`����N�m��,�T4��L���z:�\F��%�BɃW
��:M�W��"q���*�g;_�[1jg���$cMs��O��>r����sg~��a��FWd��̮x�7�W�����ǲ���xnlm�����w[�=~���iMhԸ�p����>PG��O4iǒ��j�oGh�0��]N'P��`wZ��΅�JSp��l�6�Ų�m�7g~�pX��:�cZi�z���j��q�$ݤ�Z}Y��F�:OE3S���K�����ڻ�2���Y�K��k�LfOxϮ����i��!M�/��]C��:i�~�\:��B����b��:�W���� �p�:���CX�.������J�9ɼ��w��_��U������w����cY���^�!�\�F纏�يs�1�3������PuS8�FJȉ)]R֋ 6IV,�8����C�0�]RP�Af�n�)Q�P���Ogo�.W�z��=�o���m,�{� Є]ك3���E���m�Z���\|�:F
9�lQ*����<�)�6�l�"Ac
S<��bx��U�Y�^��{��`�1���_��Տn�Wsٌ�l�s� ��oox��r�"� ����z�Y68dao�[ysƖ�{}:H�}޻�5pG܂�����$�@x�(c���o�T���NU�P^�ߧ��?��-s�.�^,�䪴�r�br�r<��X8`��Rv������Rγ��Er��<Fm#}���D�������su�2��V5$��nv��5������ޕ�e�<�\�	�3_S���QN_=��/�}U�}����聙����(Ώޅ�(Z�}݁\f �v')c�/X�{�WR��o���_�9fB�����Fb輌A�K�\0۽��o�f���Aڂ0z�H�p�n3�W9�#S�i؊�Y�@�ʷ	5~z�h"g�1p�I�Vm��O �Cn��ޗ̎'��o��(V�oEΚ�YGk%��"���_7V!�����:�ʼ'<MY�=�?{n_�d�̏#=�1����`���ɒ%^iEl�ڷ鍊�\�N��L�E�mvmU��a�-���ۅ�51Z�{��>���GD�u+��yL6�UamٴD�C��	@rr<O���4�*��K�<���\����x�M�J=鹨t[I/� �w؄�&B���_Q[�8E,���W�-���C�Vo8�Y�|����vl+��e�N$l�3���j^�lE��5wd�侈�����G��fu����Kv�̼�*�V����&E.���9�Ө�T^j.��=+�7;�/I\�Z]�sQow�ԓcj���"�B΅p���	���9��!��β��[=��ì��:^������J�+���CJ[8Q�T8�l���,�p�ƺ�"��g� ���!r-��
�����Ӈ2�gE��SYဈ͉�mz��w����_�B|�Bv��ח�x���p)�O@�*�F�8��\�ޖ�j}�ټ+ʡ:���ݾ��i
�N/���io:]t^n	�ȳ�wi�k$�b����3Û�޾:w�Om������W��0a��n5ұ2��o�f��IsN��
Aw'V�&B�'����;��2ǻ=�x���e��+h��W}.DvraN�2�/��谨&�Ǳ_j���w�K�\��#"���1�w��j���sU+6�,A�Q\��.wW�I[�.�^�w�Jq�\YN���ڂ;�/�R�Uu���j���L����3S�ꑞ���r���l@�Wle(�m���_�G`�%�#o}�TT���j��rj_y:Ʋ5�J�c��V�:��4�I]\$��9�h(�M.vW��ָ߇q������s�"s����s�j��{t/��w����b�>����y��V֊BP�=�# ����y���ǆV�� �P��8�[l�w+��X��:�,D��?��S�\'���6��ءc���dݝ�/��J��)Ÿ��5���Z㤺˞l2�w����ڲ��5UJ����]L�	�f��q�g%e��q�p�4軼a���D)�']�*V�i�f�هp`/ɵ�o���p��.��],�Ʉ�u��`RR֎����/.i�h,��Ż2���p��m,�T����ӏ܍���ke�.�.@[Oi�ԭnk�{G��oPu��tJ"̫�*��Õ�(�B�S퐃��g���H�S���5�qoM�\p��Ѣ�U������ A�uԹj�*7oC��^a?��,t��*���(şU�s)�9`{�'���%�[Y\�� wYrs�������k6��&���Ex�0B8zI�%d@Ay�V-��w�J꠴RJ�{D�@�����͐0��A���V�\oJ��z�>�sL���9X� we���|W[q�ȧ��oYz&� �����.	Y���*��d+l�<���'Qy�\]83kם1�Ӕwom����w��� ��qU�̧r�QS��X/Q��M�F�3�v��۔�L��c�"Ҿ�-��yT�+*�ڹ�N'kB���_e�i�\���cF9�<�P�Ť'ġےd�EV,����"}[U=�b�c�->���U��*�κ�M�<x8E�c�
�`�8om�s6cT����N��U�Фw�v�#��k���i��vhҶD|�5n����v<���0Ix6����(������b�sڬ9�L�RR��7�;{pp6��]\8��BE��"��\ܜ��Q�y]h؅�{&gL"�#Ƣ;��\b9���L�ewS�ߙB�ve�ȇ,v��v�*�p��۱����n�U;:I.��g]�x�$<��oP�d����|�mۭ����O}Z��Wh�7J}�:,�bîls��.dnS���Bƨ%�
�3Zm�wi-�ʪ�,�0�����F�=y�!%q�ٜ�-
��i3S:Aasv���{�q�����9*eu
���3�QN5}���ii� Վ�s=�
0[���iu�ulV���&S��Z���ř��Y��� R9�D�:�i@͍<3E
��E�N������i������5ք���n5������p\�΍��rV�MKn�����7����I;QMJ�"��$��f�$nc=��D*�iV����BHHT���[޾7��Y���^�S"*��ѕ{Fr��'-d��D%�X�Te�B��������R^T�M�bI������F��̨�SɄ��"b�6am�""*g&U�*��3�26M�Ե�N��T�6�S��S"����j���sP� H�ɌCS�DT���R!����S\���4H����
an���l	]���==Ջ;��Pu�<E�"�L�Ȫ"I�tݰ���Әnv�9$kh3Y�dX�ixj�DbQ̈-CTh�]�QE�Å2�m�B�	\T�(��۬%�kmP�(�T.gj5!I�l)Q<�il�+2��
�Z4Y`�j[jT��s*���{����O��OR��#���?�o�i�*��]qn�r��:yVe���b�s�� <j+�Q��Ż��7�kX�1��� ���Yַ�w������Y�:��<�Tv7�K_r�щe���;N~mI�\���}����b�JSp��ӭ+.'�\q�Cq�y7��ԫ�w;�X�.�~Ҋ����]u���٬���Y�0aP�'����qrLs��a��6�<���SQ���A.k�Nî5%��Bq��-���݃���W�/U���4�D�'%AK8������:�W�nr��R1��L�q\�Z�ڄ��C��|�Y��Bnv�����u?o,�'e���
�Q^��uLVl��0^�B����F�4�Z���W�^�}RR��d�#�B�Ɣv@���<ĥ�v�5�
�|!m݇���{��av�1ǿa��E��ܶ|�̬�fgkk���p�W��r^�\
޷k�OE��f�,M-ӛ1󗝚jťܷ,9�m&V�Q�dC��o:�z�y�������o���Ddֻ>�}[0v�yzVr�52 ����fn���3�m���͋~��Hʸ�Z�J�\�K�n1ɥ
n�~G�يu'�s�s�]7p'����e"��fF�i��&��6�F{�Mg%��.�k<Q���!�ͮ݉b��.���1��c�=�R������. �V<�u�D��"��#Q}*�hɯf��5��@�r�������W�j�IHǎ�̾����ݽO�n�D�bL�0��Ӻ�v�=����o1��X�Q�=�����l��j�
��q}����&o=;�ŘXy'q��v܌�.��/i#�{��M�ќ�"���yc۔�͚��n�JwȠ�ܽZ�#);�`j9;;��1���.b��+S4�ѣ�5v.��/�6�:(s�+x�aU��IpIq��U����G��>��G�������I�;:I�(�dZ21��5��yr�K�d�j'��r��G3շ<����gw��c3eн�����֔�cQ&�+ڥ@��"���6��댝�����^��n��D�����"c����T$���"���WfS���d�?��������d��}� s����m���?Qy5�e��<�C"�`�v櫭���𲶔˄�D�E�}��.Y�c�L��|n�j:��¬���
��JxUPQ�ř��RJYS1���,M����!��pVc����յL����ǳ�f;w;��۾����Z�rT`�q�upIB�D�6��&N��4�f�8�J�����D��ko�׆�t������X �����Vl�f� �p�i���I��2}�Ͳ�N8�u��/[�ud�%H�k���sJGF��>f3#�}�}_˪����G���O|+�\��vҾ����d�$�pٯ']��᧌�r�m��q�}�$��Ƣ�O:Z�����!U�*`GLޡ�����~L�Y��J"z�[Dio9���W�s��]�qEd��f����5X\߹7|f&Y���[x�v��f�3�>�v"kDM�:�Uʟ䖨�FЅfuHOE�������9i���R�9Lu��-�V�s���N8&U��~]#2�{x��ڷ�ݿP�f@�i5yq���}<��-���]TT�]w⨉���"���E���MB�u:^Z��+�3I����Ww��rk=R��Y�V�Aj眙�h��",]�:�KQ޺��o���ɕV�0����u�;�P�h���gF��RY\��ݜ�򴺀��.�j$�JV
�w70ЃC�b-�J��Uq���:�NP��C��9�x��7�O�U}���������{����w��b�7�\W	�&xIlR��e\+����[�y�e9A�Rv,�A �d�8v(�5@�T�F�u��T�V��P�e_	�z����{__���3y�s/,S��¯��^�Q�����s���`�؊�/u:����w���P}5�_��XY�W��K_,�]9�Ku�I��S��&���O���#��Ҕ�g`�I�[�����pt�V۩9#�ca�:P��7�8�W&��}�[[��T,	�f(o&��N��ڊǙYsy��ҝ��I������W:B����Z_C�����f�E�or79?�[��=>�k;�����(ԋA��d�<"X�˺��-������zh�n��̩��A`��������O}R�.�e��7
L�����B�Q�T{���rQ��#Eǐ�[h	MMBA���� 2(
�]޷�w�z�bM��m��u6����|ӉT�%|�轼Q�3���Zs�"J3�bȇ�$�̭;W��8�T�P���Ǿ�[��q��:/=!�e_;�������b��jjpVI&����\&.6�r�(9F�-��^8NU�\�m�[�R[�h��Z�A$�L�\���.,ڻ%�mnK	�uz��k�Jᑾ.gg���.�U�f�ګ�0*�^ۙ��h�2���X]���-�yN�[�����,wP�Yj+�Mn��̇�'w�\���x[�w�j�ϫ_`Yka�̗�r����i$p�Ck�:y;��W<XѺU�#9���"7GW�o�$v^��n	h���F1v5W��q�W�1�$g]�7�7 ��`�g<�)��L��T�����z^W��-�,`�k1�l�e��al�)pp.s��AdU��9m�|��kf��-�fmm��Y�`�����ܲh]�'�2P���jpP��ݽO�{0�SP-˔��Q��eތ�Ȱk��S����v�=tX�V8�98�i�BT�XWL�p��Ɍu�zo��0����o�m�뚱=:�mQw���g.0��o���mrhf~�e{����5�ZE�n���� 8ݬB��c�%X$���/�s�!����o��E&���~!��� *.��d:_M}u��y���z�K�t��Ջ�~:",�#��5���j��!����L�3���]�WP����������!|��}�4�Wp��h�^��0��T)���:k�J���Ί��7FM�8�5L'E��P�? �����BK��Y"�%�M7��ˬ=���ȭ�v.�Bn����W5��7�Z��s��(
��|[?l�p��;�Q�c�ۅmfхJө�O�g�<��|��}�)G�")`�÷fdN�tʎ�Mðw�\�	����p^c����$[Z
���go��q���yD?w��L*��nA�ؖ�����ǋ�=[]�g���}	��U��wt���"��S�Ed@�cQ�y�����8V9NĘ�[ښ�:ɚ�|%d���x�>�C�&>�Lxf������	���������>��� x�Ԋ|��{f���j�ge��mN�'����ssteԅr��Ο�h�?�c:���M����:Sz�ŹK'�+�Y����}��} �A�i.#�H�9~�	��F��׏V��M�B���A�]�U���T�JĠ;��;����sB���>�7�H��N<5h���_�Qu��|�Y��×��A�Q�<�yn�Ǝv񷗰Y��P�{�_�"2(����y��׵�W1�m_Sq�){��पf�aOg���Bj��uG�՝37�Ҡ��B�HR��D��B�3�s���2�}�����,#=l�e-����qTe���"�<�J|�-i�>�>�΃�G��I�Y�K�������炥:�uH1���7��h�X:s�
����&���)�K��Ӭ�a�b�`cI	�/���]���S��i{��F�ķ��tIdqѩ����b4թ�
�&	�z�Y���Q�9�w
�ܼ�ޞ�ma���%��-n�ش��"��S�NX��h�R�p�#:���O�U�0K�&/}^#�x���g����ͥx��M��f6L��4�:�ʢ��:���F�.k�C��<��UK���r����FM91���O��%Gְ��[�����e��H�W�:�Ѩ���.�zA�tohRu�	�j+4֥�5@jhs�̴��yvR�ϣU ���ub��FF��B�!&q�ä�u��������=ٍ�;B3��l�ffZL������o|�w�|�EADZ�g}���Y�{5�;]#�Û�UNo؀GH����T��5�}�G��گe{ݼ�%9|�4!mFCj��}u+�sp��a��k�5�lm�^�n��}ѭ�8k�փ)��͐�2r;�w��m�:y��f��h��EqIݝ�LЄ,��;=T.���h2��>�8�3~���"����х�]gJBVWS���4�m�27�T#�ԥ-.y隇b�������m=��\8�*O�Ȑ��U<`�HIР���@�U��vf4n���������>�E���@��^6�y�K�R��ə�̙�:�Պ�y��{������@��`����]�YN��zi_���k72_��j�L[8��{T�Z��ꄆ$�԰�@�,M����W�3X	i���d�_0j6����EÒ	�_5����Z8 �����S���.�ِyP�#t�y�i��['[�y��{֏aZ�a׬��7�4�e�܌]v%M ���5�b����BDX�o^�KYA�����*��$��Z���Q�o1VkwjW�Ԭ�@ȠHޡx�M�\�ogX��
�ЍE�F�pj�����#(�������6M9��V�`=�L�b�ْ��S̬��<2vZ�q�2�u��}t���(&U�}�WT�@�l�e��4�荜�����yٳ��������Q��ev�;���׷|����4�,�T����h�#�߳R�B����G(�ҽ��FL��U��c(vom���"�^�i��ޢ�HkS\o7��Vл�{�3u���q�6�@��n�m����z�c��.��g�����S9���3Z�����t��� t3[ޙEY�OE�e�cx#�40_!��rB.��ϔ�*z��k
6���Î���}�[�V8��Ӡ��˫��%T�2�k��{|��ƛB��b���3Aţh[��{[τ�	�4YR�ܛoN(��(	)r�T*X����Vd��{���l3#��K��-ߐ��N��?,�f��&Z�1BwU��X#�med�,LٖV�58a�,��R�"˽�`�B<��o.p��G	OUH8�M�����g�W��v����V:�Tv����@��<=
{�r�E�D���mf%��o��0^pǽ��WԹ��7Y��BG8{F���vk��u�1���ӥ���d>j���;�*o�2dݎu�,\$\�U\�}�o�E�d�}�*��.��
��_�-y�}��M�J�2�,�����3�0��74�U�)Z\�S�(�#��g��U�V�Ս,����ǭ�ٛ�J�5�4>��&f����#v�]��I��C��ڲ��J���ߟN�;��X��� �f�4r|�H��<��d�=�m�9�UO�ͬ���k�����\�9� 0�m�tU�
Ь�uWxGI ՚��D���D*�W>T��@[.�'p+"��:Q���t�y2���Ȋs�i��2۱�e[%����"Ӛ��]a����Rh0G���1��(/)p�L��B�X�|��ϗ��"�H��Q����A���D�EB��fDt���ݦ���42�Ͽ��=p��f+�51�I���$v��B��u�Kdˣ9��R�f�ذ���}��6�ԣQ����z�F$[�ѳO<���M�ūuЉ�)�Q�ԩUŤ�#�'���u\�gu�����.v����IU[\�g�����u$�;l�nyg+�싨�Lʋ�leL�<�=�&FG]�	�h!U��*�Y���+��Ԫ,�9-I"#�:x��WJV�(mm��/m/.���6��ӡѶ�p݌�ؐR�j��$��&�C!�]��i�v���t�ڇa�ݶК�-��WB��uuW%�λU�na���m�3N]�kV*��Х��F���W��8 s���w+xu]d�mv���w���=�|C�5�z�5�Z��Vy���7�9��E�U$P��?w�ߝ�_��kN� �렵q�����j%*�Z��Ȕ��|-���uÔ������o���U�%s%��
�'/���T��{��gR�,��x��j��'�q|b��nr�j�J����4(���˴�ŵ��kUl�l�;Q<p-���t��K+�znO^usy�lxvvz0n{ԏ�
����ooם"��S�������w39�Jۺ#Ѻ+��;5�Vt�?/ǿg��-���~3t����_�n�<��˃�"�����2�]q@��V������걦uy��=�v����#�|+Ж"�%Ňt�>#��cxj����3��n~Žj����H�҉���2������*��#q�Um��ƫ_�w��j�E���I�b�����ee1Nz�N{��}N_P��2��� ��g{-a�6ȐCT;$*42]ʔ]��7���+ξ���l��0�8��)ԕ�vM�2�(��L�����(�'V��t�GRظщa*R�f7���S� (�\�5��>�s�f�	�t�&o��;K9��`#�ia������t�I�v��ʗ�v�E1>��f�`��<z_½Zj�Pa�E���qf|���*��foKC
��,��09�B��1Ƽ�[+9ٵ��מ{I[��\lxw5�F�Ę#��BS���e��1&�Ny�s��wѳ�x�j����y���\�.;K�y���i�a�G��G������k`�U������ԛ`�_4E��� ܦ���J?1pk��R��{�;�����^�;Ez\P��o���5x��pdJ!��N��^0�h�#b�Is:��#N���uw^��tMH�k#!���#Ճ.�F�j%�A���p7]�gQn�'^�w'�L��yC�E���U�fO�,ٳDS�(Ȧ�����k��T��꘼b\yY%���Ao�:�x�-�b�t	�J��=g�].��M5�t�{����� U�wv��#S��c���X��ы��0�4,����80���,c�q_I��� ��*��*3��kӪNqG�v�;ݼ._w��T�S6�9���ľO�i�b�ʫ�;8h/�
��.s���<It���ppeE�M�����n�P��e�!_�ۘ@��j%G��Д��C3���Q���ų���ǐ����q��ڍ4���)M��E�#���Rx�T��{س�kә�5�9/�m��T]lX*eZ��M �x��9![󷙞�Kd���']������޷0"�)��4�)�Ĝ,t,{�89v����,��C�O�����->2����LМ�=�e���!�:x�WJRՊ��TjeJT�_'���Ri�XX��Hw�Mv2����QW;L�Np��1�43Z<�|�z�~;0K$�4�.AJ<�]u��]o����{ ���f���������C��6������g�5��ߨ:Ww�w����"u����9Һ�?L���>�%��z�kO�k�uW9ApI쵾�{Id���o6�8D�PH-���v՗��&kk���:��sL��)q�C�Z���N;��u�SF�Putt@��].��l/�'Y��BE��G�(����w�wٽ�h|^��&�����gģ\���}�O,�0b1Ay��Kв�j�+�5uS��S��c��5B��,g�^��GR�<pծv�����gr��P�>3�Ơ��H�:)Q�C&�%���Zu_dޥIҳ�ǆe\��?Ə��L%G��f�������S�u��Q�����8Zy��~���{=3����e.K�R�"�2`t��>�Et�[��^��tx���-�%�<�Pھ��^v��ʉr&ڵ�����=/7z�[���_\�NT��N62tі|.�vj=�f�����{.�w�<F�cH��a�>I���ս>3��ǒӕ��]tw�PR]�� ��m�vs]�o32�b"��+�q�*:ny�P�[V��Ϥz�uu��Z��`"��z��
��T֟W6l$2!�R�~@	�juM�j*dM�]ek9��=9���4���
��V�O��|�ww���� i��חO��vC�Q��)2��6J�*o$��W�6��g9,A�k��=JZ�I��s�|���k�(�AFDf]����i���ɥ�dZ�m��j�߫��QJ_F/(�\��W�h��F}����Z�H���'����2-]��H��1�1{�P�\�� 2�������;:KԸ��X]�����Ɓ�R֞7��,�7V4��;O����֣��xլ7�ڮ@x���rA�|lV�9:��`
�G���^����x���� ܂�q��LrkA��+�MmRy�(�[2$�9v��T�"f.X4a�o~b��~���D�x0�KW������!_�=���_R�c3�!���0n�c	�W���ᬷ9";zƦ���S����sj̖��\I�~V9Yb��#S*y�ڸ�c�h��܉�^%��5WJ������l���ݬU�F��Ft�.��WT�` q�S��j�L1�`"��[ðk�Vt������b8�Y�)�-͞ڧ
	�o�j��9�:�o��T�dhq��HG���,�'��b~�%�,S�C�7St]���VX�sn���k�����C�b��P��v���K�_#�8���KrRJ�<z��s*}d��u�w޽Zp��sJ%�����t��O�����zf?OZ5�wK��~6��#�දl{�V��k�]�ʃZ}^d�^$���g�z��V�����;���Q��B��B�J$�7' P2����j�z6��Y�yX��{����Xτ݂;�J����q��HɉES�:M�WJd1N�o3&����`�+]����[�^ �W-��v�0�fz[�\j�N���{�yw�e�3xCڌ�Sס���E$�n��F<puMՅ������I'�x֐���X��S���c��O�y�q���X����;9�\_&_OEk$@�(�[bL���,a4��Xt���;'�_w��kV�pd�qB�WNw�U~h�>ZC��&�c<��y!������*��v��N4*cbL��؅�p��G��D�!Z���R�<��|���E���Q��������>�鲺VAy|����T:�rB��z�M��� jsz�f��޼3�+U+8֡K*Gp۷g�2�]quoZ���(bT\�w2��Bt��ZĀ�������$���������b[5R��nU�c}�.���5x����2��6�'�\ĺ������Tt��C�"�C�[�Qwr
�~Y����4uK
�һ����ss�)v�L=�~!�rx��ΉLW���y*����eG�:��*�޳��֍�y��|��`�8Zlg��[�KZ�ó_e���ŀ���,�qjN*>1c���j����0��b���B��|��Y��E7�:��n��=c��'� i_5"�%G���X���P�܌8�k��$f�A���^/{˹y��_����"�w�f�{�\�B����V�R�Q�pl�0RU��3~���K�wC�z�.��^�"8��A��^�>��'�����~5��<�g�����]��[Fj
�ʗ��A|q!.~�_%���om3Bs��hX
���]�ѹ㌬V���l���l�����څ-_%huϩ��r�����R�j�GNr��yOF$�u��b����Cg�t5 ��^�A�(ֺށM�*C�DNފ�vd�o������o��/s{��]�^��k�czz*a|𡴇�0��J5��.1^�{6notp�[/8��jG�[������0J��a�}ݘa泫o&���A��1r'�L����/	���>�Ʈ���]3���y�=%i��G�O��<���#K�Ԉ�Q,w�Ԏ>C=��#����k��<:~���	����_b�\p��9�{;maڿf���6��T���/ˎ�*���63�	��W�ּq�tȃT{��)���C}���i���,Z��Xkʾ���jG�Ѷ��&r�N�C'��?����b�p߾ʹ�@b'��J���o��(ya��O}�^4g�^w���="A�=��7i����*�7�������㎧���l�TP���/P*��K����X���t�V"t��}�x��.^]��ۖ9��tP�]�ҭ2�AN��k_�6/xnf]���~���J�L���"U��2v���"Ĩ�YZ[�M䥺�F,�2�gM%��/(�r3����R���������� $���/��}yע'������)����,��͐�2r;�w�ܦ�d��N�[��҃�6r4Ɛ��t�N,�ڷ��|�[�Tg��=щ�j�vǥ+��,۴�ֵD���Hz�m����
��>�GM�禝�b�pmP���{3���T2׫��Ƅ)��1|��
��~V2>9B���2�eud��w�H�״�m���0�!�@4!� ]�K�X���.�)n/;F��Y��r{�f��R�F�_�=ޠ�N����0A���ʌ*Z�eK7��%bѝ~�j��W�Y�n��5~>8{�Z��P���F~���Y��]]پ��L���la�Z��FӮx���rA7K�cW%Z�z O={���q@O��E��&�jbS^|X�a$Ǽ��|Ael�^i-,y6ki4:zme�9�-.ș��0�v���W�U�%s%^����5(�w���8M-<=�](���iS�lQK��s-k�y��e��/�kc�;:���9piN�IoO���[`΂R�-Neh�M�G�>AE��(�FS� ��� ~BA�1��~�V����'7Zi,=K������/jqs���㇗��M��('�c��v���LL���H�w\�c��.\Z�����Qy���^�;����|^�9/�TvQ���l��g���N�zw��W������z�H�s���0���o�~�Ο���b1I�TZ���b�~�o�쳘Pfb�K�/�s�`���x{� �S*t��Yh����ٹ�G���#���$t�z��ę=$�d���r�5+��,�u�)�m!d{��PH1�م���OAԽ�R���d��_kEo�r��<�".ϰ��Z�]�l��8K5rXw��VZ�Wq���S��eش�d�t޷�*�Vc�����x�9���G���Uk�H��}��C*�s�#y�S��*]F�h�Q~6�F���wә/�G|;�_����� ��R�L*H�V~�v�X�W�+�΄�c-�_S�/ ���H6�C�j�(r	��Ȱ�w%��Cw�1ZާMD�Yu���A�Q݅]���Ef���#�8�j=��v�#���k_U��[9��LK.�G�V�*��+�߼v�G��):4O�k�-�9��9����`/�~�K�imPvC�o�0�̘��Pn��2��)�B�����yY�{f�j̲�Nfd�ށy����:�V��;�V��X�L��O��ɮڷ�eWQf�y�ϙ�܃^![�a�\�Y�*y��5F(u�Y��䫛���3�M��%���޺��2!N.�{l�K����ϰ@r��qNp�.���k�G9�rE-�4�+B�N��Ll��Q��DQc91Uܮ�w5>=><�N�4�$t�0���T���S���;i�v���%Ɵۍm���n,��zV�A�Z�Mix3]�3M1��D�m�S�S/)�
#su�"�f����O9�Tqf֊w�9�ړ���h�yN�)۝ڄ.�wj������>�����`Ss��hs�7���I{�+��;�@ϗ!��
~��V�*�V(�7e)���6��7�uŉ:�ᯣ�T7��Z*�:� ���9i����3+��5:�d3�Tω���݂e�KN����%����p��<�C�]��
�j4����ĩ/��[��^m��/�*����@`����Ԋ�}f�;
�038zs���͘�*���b�[�p�r��s^f��X��*q�o�̡�y�>�J�h��VpMk`��d���MN���G�*�"E^Kc�ݼ��岶���ђ��j����,��Iq�	�D����u��XQJ<ث���v��+n��ݹF�!�˔J]([����/;f��5�|��C��M<v�]ɮ�t3K*w�}w,9O*��(��M_K��n�s�f�7�FӲ��gG�;���y�t��X�!��mh�1Z�PPQ2�՗}Ȓ����8��H](�gv3��ͦ�R���0;8:]�걬�@�&�;�v��2��"�=Oo�wI��}â��e&�d�Ya�t,d��s�\��)�IU�W</5=_����>��g)*N]谔9���m<�l쐮H�&z��b�tO��x�kΰ�<�c6L�
:+8M5)99y�y2%Y��ȳĒe���5��:)�^�U�Ӟ��a�%I�kH�[\f���l�f�W��X��D�&��=*��W=&�'Q��\j�Mc\��ias&ei#m�Q�2Dm�W�<�)�*�aU�*2���L�1D��NNb��B�-���;����^0��%H���X��\�h�%6�9�Bg�G�G6�^QU���Z�^�v29�碅���t�drm/E
	(�>D��$��}���B����z��@�it�y�d�h���Y�+�����<w07�[�%�$�D��U.���A��o�﹚䴛�I��3z�E�K_�A�F��()��B��ae�mn�����^�:��}��B�o5�%�%DiBx��Tp��!{�ٓ��}�:��}�9�xe�;�!�\,
U�UdCb��􆐀�A�����̾��כy��Zb�����h>䈠pj��H6�mԙQ.�`1d)�
��EƼ����j��>��«c܉���N��,A�K�;)��і��9�4}��h���D<p����z
,]�P��gؕ|G��B�(�j-���ݽԝ�e�I�t����$���xO���񣗯�_����J
~���>��b��OL8��SӞj��ĸ#�!�FzAA�!���k�\N�o�0VM�
{i�'�J�T|b�eOz	��G-�YG�\���r�/��.-'o�eʞ�C�rx�@Қ�G�y� �+}��}�^b�FV˘
� �9���f��t/��>o�:G/=�E��8쮾RJ涙b��A��9���)^u��Lw��γoS��8�IY6��G6f�,����j����}�����������g���T~�a:���: �P{Q�KiB�3TMFVȹ�O�l���N)��#�m��lJ���e���[��Ő�a��C�U�!��	����N�~��6��%T�PH�X$O����������l�s|�{�-R��Hl��������:O��Ե$�h,h^��2�A�	KpVu𩒞���cb��/c@��^P%��S��=T*����t���o�ҥ�����A�2�3�!�6�/5��/K�4S��v�ʬ��{�d�|��"*���#�����H1�^��� �;�6��d˾�z�T}0��"u�8д�����&+�j��dȊ��3ƉHj��kN�5���<k��'0��	BqQ��d.�4��@}sא�/[{&zF��k�Q�)A�L���5��	��Ƨ�����-__gfU�1m@i�U�:}��tti*�P�/��-Z���t���n� �,�j�fD+R��:�O��=V�ESi��g"����Ɓ��e8y�,���ө��8�_�#ߧ�3��P�֋��M����o��E�f�B��/n�P��F�����g�7ʀ��M���ls�;���pb'��J�	Q����s���)$[���e�8��;�.4A	���iMB�;��mp�~6y/��H�x�<�s$� �t�J�N�L���ň{Q��>Ke~ߧu~�W��:ri��Gn:"$z�b`jv7��\�9ri���62w2ȋ�+�Kel��3Q��	6(A���/@���h2�>L �b��O\��"����{N��}�rdĩn����\ zk�]�əd�}�SИ(��ܗ�յ!D�p�EI�����:}��BHƆz��H7����5x��nS'�3PȦ���.֥鸮^@���{�����V���u�C䙤�����}�AН!�1�V��	�1У�u"X7�D��q���8u����ݼκ�q�U�n�C���-������׶_`V�T��CN>��B[�����R��OJ��d
9&��t�����Y�{��L{�1�D�i'����VQ�g>�eߘ�(]�~<h�-V�9:�#�۾Fn���z���G��jʁ�8䃋�>0r6�����.|rA�W�����z�N�٪��r�M��S¬R�+�(GPe>.������1�kj�����_�I���^Y_~8g�O�����"�\_�c���z�=��� S.Xa?���{��%��بu?D���0�B/0zVT=y<���å�V;��P4��]���:��X�t*�{p���"�UlS���O16�f�=sr�0T��4l�N�f�?�h��������`ٔ�3�����6+����R�q�\�>��f�Ef�x����������kq��r����j7�Xj�T�dCp2n3�(��їU�u���Ɖ���$kp-4���\;�0�]��$��u��>�2Y�%�;�bS�ب�j�#ku@fр�wl_Kw�xY+i�)-����EN�p:�'1�y�'8�P�T(t11҄�m��S�{�����VX�f2��X����Y5&nu���P;�W�G鈏L����<[�����j�f!�V��pc֨!$,��\�6,Jȷp�S`�8�����i�Nm�a�i�lX�	Z�4!l&l��''5z���5nuܞ�w�GƢ�����."`�����_q�YȔ5��ӢM����a�Tq;.�J��a�dS����F@J܌�}8�ԗ+��R���1�è�^"I����C���o��.�Sj��}�py�JL�t�k]�\lΠ��(Ws\�o�K�/�
�&)a�R�l���Y���+�n(���r;D-���M��UO�'�Hz�Eq�f\W��<�����ӆ�$�k��,5Qcd�k.T��QO*���MoEN�X��X�~���0�sI<��;�>��Nj�3�
}��B �i�7'Yw�Z���!p��?��!.��W����j�?��h�����حK?v�f� �r����>�V���"�b���-�(�ݗ���N�}���u#�N|�&L� �/���oJ���BT�S9�7��i�U�}(L�+���%��ӆO��/�E͵����7���/G��Y��t����O��HNV����{�\�ǻ,t�� �����F͛B������$_�,�=�dp�4�r���D\�dy6��v��id��G8��n���(h��X��A5{��o�G͝�P�m9پ���$�+9;�	��؇�:���񀁥5"�Q颲�mt����G���Mk(Q{=����g����^ł�Kma%�/M�%�u��˩��T�3�c#tp֮K��G�f�/iٱ�m��\@�}�'o���m$�$���[�z���!K��sԧJ��@�c1�I�转JSbeJQe�u10�=QQ�n�T�Vz�˛�!�}��r�b\uw4�5XϦ���e*��H�ב:{�0�O��%@�:wOw���PQ#�x��.��ɜa���֏�\�{>aɣ`B�����uf6�f5A7B��d(�ǌ�*�y�S��p�+�U�ݎݺnV!A�o5��z}Xdt�b�һSM[s��J��Н&*k?`$󬷤��B8��a;iݚ�J��E��]=
�#����͌k����13�T�Ld�
�o�F����4��a�����]��ic5��J�v���,T)��
�	���}f�`�qy�i�E����&ƃQ{�r|CT����9������F$����E>���g}�/�ų�$���c4��U+	K�M���yTU�	��]O�{�����_�\����v׎*���~0�!���r��=A���z����'ɬ����n�v���s�->�g2�x�"y���	Q��Gc�`Ÿ��;�w������F��ks�%5Xݧ�D+rUS���Q�����[�]�ɃO�q^l��\��R�����b�6���a]Ö��싶�_ow2#>�(�_�h!;��W�O�u�v��7;����N��z6��Qv��Q�5�'�4��kg�1�@�0Ο*\��ra>�3��1��O�s�Y�t�A0�d�K�i�������M����$�Y����򀕧oR��Gof{4yE~��1��\�)*R��ʜ��Kb�Z��TԘ]p,�E�a������PLI΅��s1�-��ݛQQ�������ꔶ����H����*8�������f_vs�˵�܆⃸0+^�w㲝T��d	Hcʬ.�EnkrR�1��őx�W�A�zQ�C"�B@�kR�8��M��[�{����wT�8�Xr,"��ޖ�?�����@��bbb�\e�'	�0��\�cjU1Oh�ɧmr^:)Yw�vRb�����6E-��ʑ�F:�0Jn+J�W��.���U���rA�ן�#i���~>#3�:�Eɖ-b�ɬ�Fu��sk$T�ƣZ|��T�yqϫ�I��ۺ-��	q%��W��ۉ�hR�����<hu�}5�!d3-ao�b�P*�]`�ļY��Q{S,�C�nM��VD�S��Φ�z��'�u)��Eu@M���X�Q&r�u����;C���w\�ƍ:c�Ž��c���=K:�1�ʆuE��Q7|5����j�a�\.[/����`�4[z22�3D�s,�a�U��j�s6�It@k�7�I��0 ���4���Q�㸋�n!���ڋ���g�M9�����vTg�����������JrU^><��L0�#�s��O�%�.����G�#z"�z[ó_��CW���'/3���{����0�~,C�i��Ê��\L�n_T(��2�ζ��]u��x�Wg8�υ<��c�H�ޑɱ.�9���_5�ҽ	�ě�jj���ݽ]j��Q��}hn�b�1ֆa!e�Κ�9U4�<���Ф�s��c~��M�-R����� 8{�V�fhB�f�Jg�nAy9)"N���P�`t��n�Ӥr����P�w�;jD��ѝ\�/h�^S2g�]������@/1�[�7۶,N��ݦ�V}�r��{�1i݌q�E�ƢIDa�!5��cg��_ac��	�Y-n
�Y�q�M�xӡ�jذ���gQa�5�%�%��x����O��}�{d���\{�WL
��`q-�9�ο
ʏ]]�C��,�ٚ-ݪ�����ᝧ���XE�V�����f�QI��4Hw���|ֻ\���'H�[Δ�f���B��aFR���~�\���`���C�S��<}���=k��c������|��`E�㲑�78�,ۻ�2^	ꌙu�����"(��lm����q�L��+s;�ҡ^���!���4S�@��܉���I��,u8*��?4F߳���[����A�O��iyN�!��bjwR��[/��NpC;���B�߽�`�CE="��->��!Xߎjg��~Pƈ�*��)������)/�;�Y�f��Tѿ,�$W����o�\�Noi������r0�Eћ��x�)hag�:���ōZsނA�U�;��Ъ��/Dt�����q|]��r��X�rx�@��h���6�V�;�ҞC~��=�/�����)���Ы�ظ���dm�,�ֶ�׽�g�C�T�(B��٥T��9{NYB6`r���� {O����wF�J�؅��~�1}���gc�(�v$�z�pN�k�*��Wϑ�,�|�ݮ�)�f n0lp�k.�����ѕ�%�k���j1S^��sU��X�ݨ%dԏ	�o�G5��|5J]r��:pd(�"�6V-0�\P��Q��t䜺dOL{W��a�L�8@��=m�]X����-r������*��Ɲɸ�W[��~$^�q�{�j�\�%�\.�1"n��]�	�{��ܜ���]���!�+r:2޺��nZd��[ʛu���4l�{&JkE�7AdXd��YsM��֒]��tr�{+�e�F�H_���P1+F���3#k�r���⬶��cr�DhS�I�Xݓ1�*Ι�)먵l��P�Y!I�ϸ��3#�B;��>�8r�:��2h���چ��bZ.D�k��{����;:��As���)�g4��vE�oW^�ȝ'�!R{�Ŕѵ�u��Wuj9�&MЧPtC���p��U-9�UŎ;���|-˥��n�L5�ih̘p����*[������P�tzo7m-�})�y�볕v��;�����)7/^f
ɋ��ܪ��خ�$��أv�y�TO�8t��>�,��J%3�ـ�b�5.��7�F��+��޼x�jI��Wɭ)�k���졊��T�J���_+U�$��kff�c5�U����L۹B����+3�kR�w͉�Vd�{:k�p��2�v�2,�7d��˖�f�].�4bwa��5�D�7�o��6���`��޻�r��sE��ٌ.U����F3��n��;�M?���jEs���sU�Or�z��`�Ŭ�j� ���3�s��T���Z�x��w�%�ѩ��ۣ�ۈ��6tq�%ܱ+�,�S+V��s7Y�W��g1N�GQ���μ��خ�!�
�"�����xk+	ڼ��T��dWզ=*�MJ�ηT	5��M�N�[���v�F������R�y�f
L�d�RU]�{[8f�#�
��s�Ej!�F��]h���PI �;b�J��;7h�N�nMb�:�ڛH�#3:�e+сA�%��K�,+m�4CP��nP��EPPك�{-ӳ��G�T���nZ|C��f���r]a�nn�&d����/p�w���(��$�(�$�R��Q��h��M��s�)%��!Q$
�UTh��L�P�U����QZ���{�$<�'�L�UJ�/�"��'"=*�
� �Wr� �2*
�(�2��*4��p���D����*�P��CI�rȠ��J�SK�I5OU�#��ܱ�J�*<J��J
'OO(��"\��J���L\QwL���(�]2�p�Eȏ �ȡ55�OMJ+]<�t�-���L���Ԫ#�*��/=2*�O)�(�$̓ʧ"	�0�e������}���p!�*�mV����r/�ûQ�=|�E-�CՋ��N�$��F��0Y��ɘ\ ��AX$������/<5����<C�॓��cq2�������L�(X�%�AqB�8�<��������"��B���r��5q�XiH6*$��S&R�"�C�A�}2߰�]؉7�z�-<`�}I���Y�w.�D*~��}*�c��Ǻ2��Iqʳ~�	A�a`�����k�0�>��kL�$*��</Vi�ݬ�o��G��凪���+>3�����N����Ŗ3��?]5a��>���u�!({�Q�=5�IS�y|�?�,l��Xe#/��#w��__����cL(��C�e+hJ^;�>>1��0L* o��u+}���О��6��^<p���a�Ce��z�`G�:�Oh�+R�U���Ԩ��0�V�%ʵ�K�ٍ�\GTʟvVEVKzOv:��6�j\�B��Rgl�
�	�Cj���kSH�9�S����6p�;��Eɞ���9�7���aR�k���}��E�3Uv��<���	:�rU�ג�u�(���_�����㺍������N�8C@��!)�Z��)�jÛ��x遗�+��q��x�X������ԥ��!�FCj��L=�P����Ven���}�Yb*���/�}<ho.�:�u�CO�h}q�`���������N;�����X�<���Li>92�y��\����=�̬�Yq�o��� �u��6=1[^D���6!�c���j*TWҺ4b[�s׹�^��<��ŝ���+։��2�T�u���t�o&��\UF���Y����t&M(�C"�Đ,Zڥ3�u�z�u2��@�YF_Dc�(��%�V��^�Pu:C`����GQ�L��������I6�VPoJ����+dF���h�T�42�w�Z�-͒�1o��s�jŒB�aH�cb��;�S�=�xC�1���[8��ڕ{�1](��x�Ɉi���u�R�؉����m�|��F�t$㋱�ܡ�@�J�Ŧ��C�����<SdK�Wd�{��F�E��������Ic�/��^7�Pq�E���:|�b
:�+Ϗ!��:���_Tp%N؄�1;)U:�A�K���R쉘X�?CLc�:VNL�n\=u���&�������+�8�?J�z��~6�VS�#�P���}�w4�{WQ��@��v|r�Ղ՟Oz��Iu�aW��.��[�S���z"L6v��\�{N}�Qy��Fhͥ��t�j�K����ݻ%#ļ��ѣ�f��2☍�cl�T�GI4�d��\ѭ��շټ�UL��d�.��^5�X���.$�x|!D�Q�BY��L"�F��_���gϧ��_���7�z|�����Re�;�˻��]t�vm��3"L�����6b~5���A!e��A�>�h[�L�ZĚe^�W84B��UU�8_S�����[LծC=�j�S��ݜ'��\	�{}Y��J�Q�Z�H23�0wf4!Eա��N�+�����t�odBNJ�H����]f�O���c:uL�H���L���x��gO�c����j�U��0�cv[7%�\>�t����rpP=�q��Z/��{��(�I<l����a����L�֩y���Fo�
K/0�C��z	�ծ��j^ν�ww3s=��
m�A�sڄ.�����ZG��S-�ٸh<�l:�z]�};�D��V�U�#��T/Q.[Y�9O�L�����; �^��c֧�O��i'�*T�0f�YS�f簥����s�SǢ�uH깯�͓��戰`�G[p{I���8ɦX�����U
�����]/��sZ+2��D�Wp\j^x��u,�/d�Ã���g�S.�cc�^)"v�n��Kw=��kپ���K���VZ'Oyx��"���Qn�=yL��+ZK�@NK���{2q�(ѱj��H���H_��Q4�vBT����E\M�w��Óqu޿#�M��b@Ԡ�f����tN�.�)hP
�Æ��nG*�i�k��6T�Y֧$���E�w��';Bvvf�yoyŶI𫒜����cB�V��7�b�?C�h��0,�d}�:D7pU������qec��I�|mc��U��X6��N�Y0��Tڗv-\O߳}=�Ϗ1��9<` i;N�Z�Es՛�:�v)�t��&�'Q�1��]^���Y�~���g�)d���Zi-:�Y��i���j�U����}�6�҇U�w������dn$�}�9��i�����đ���O��R����X�ţ]���fK�]ca��Nц7�y
H"��ƃ\�Xt�(B��܏�0�/��o�cof}fwP�V5q}y/"t�$�<�}ne�NsJ�7-Ą���׎��}I�s����Ѭ֏���M�r����{o�����~=)�Y&��Q�L�A���p�6/�eM��߯��tI���/��a��#i�X��m���}h���M�/���N��U�+���J��C݃	6�"���.��sO%nWI]]2S4�pO9S�x֦[ݲyG�]A�g��L�}�%�&d�Ѝ��U%�Yz���&Y���+-ډ(�� �{�����&����tWe\
R�)�,)s�hEQ38��Pl"Oz��E@����o2p����C`�}n�� ������5���+ߖo���<ۀ�A���:���������D��v&e&��N7�[䜍��NQ��|��=�����w+�ÿ{�sӝS(W�+lAR�\�.�q�~{}7���g9VG?����P��L�~C
�NwK�%�Ս�wT*�^ת'f2���e9�<��-0%��jA�W���)M���;�G��,���>@����O�z|�'r��t����[���Qf�GK�2w2�]�A���y4����P��z��k;�8�(ar��ٜ@�9\t�Fgj�ʖ�!� &;X�r!�e�J��F���+�a�R��5��=�;���Ud��#��Z{� 
����n�Ӽk�kqVb�C/`Vn�!k�
!pDT�l��&���;��of�&泚���p�w�tK��;jt
�u�2l�Boq,����A�8)ۄJ�P�{3F�Q�RՀ����vK��̩�W1u<�T
<�Q�b�1$@o��2g�;�q+>��a����Դ�m&i-4�?��@�t�P~���=��p��x`X�=�-�>�����������4���^�p:�Ɲ�������E�F�XR#���K���m]s�C���k����Mn��Q.��3�i��:�E��D��~���(�ö����.꾇�k	'����OC��,�~8`�]T5�[G�Y"�� n*��ݩ���j�T�hKD��+�{WHt]����QUw:-U+���%���S��C-�F�2w-�$A��*��~]6�)���k�/�T۳n���m��idSA�T��n�A�Agsވ�;7���,{� �s��a���3�~B�}sHq�$�+������\=�̕��p�uqG-����	芰/Y�S"�T��.���f�u���-�[$/%X���Ӗ��L��KT�!Id��âV�SJ���엞��)s�֟���.�bv.;�W�K�/�9�p5z��Y�ڋ8�'&�oPL�A�t:3p#�9m�yن �����y���d�,$����*�>�6O�V�:�� ���Q/��W]�u�w�S��y���l>��H�-�-;^�07�V�F�!s���$��~��-:|�4	;���������~\D�l'4&jȹ'j/�a��7��M�|�+�aD�KO���Tæ}^�-;k�(<��}de��A$�7�se﫧+mz��]�$�"�aq���>���{}�p��:��@ɬ���9����*s�k 9�Y{[���33��؅�~*��&�N�`xDm1Jώ������6+X�����4����5��ʥ�WgoU����0�ϐt����p5�sDX:a��IO�3��+oɏ[!������h���R��%�{g�VM]����A׹�9�w�s%����q��_S���}�L����DH�+F�,�\v_e�w�oA)�xke�ے���l�tQ~ͼ�u{�pWJ?1s�"��5��0P�7Q>�ė��e<������z�C��plJ!�����U���ix�P�zւ�*|��#����{��UJ�F�ZX��:��(��V���^#~�$��mb�E��6�s�"����=K>���Q�v����_�y@��,<f;����W�ke�\F�C�9�f��+Ps�G8}0%�e*�����g��Ƞ�AOf����n��a>y��1�K�ү���.�T9S�`�@9��.��I�#d���|��Ƽ�pk�X�tn�U7T�z�����_��7�q���:@����QV|��'���1�R����S���B6a��"goI���!ݍ��p����S����Q3(���W�O�����ḗ	�.V��b�K��42�9�L�V 5�Ai,�X���J���n��U�+=!���-rn��	���v����lU>F�4��,�}��V��;�LR���(�@�ly^�`���a�r����0a�a=؜[���&���]�4�Xp?Vl	����g��n���۽��	�����U��y/+	i�Or���.i=h��q~͚����]T^UO��?�tL���lvƏ�2�L*��n�,C��oJLuWT��	,&� %4L,�9F��4��`6x�F�+�&^�_����$��r��'��g��m:D��ƙ���v���m���fut4n�/�kdx̢Xz�@֟M|C�J�|�O �%w�W�R�����B	ap>�����!�1�ϭƄ���>0��jU{0�o��,��/�Ś7*��e�(iX�=+i�Qvv��L"j�i�n{3F�3�w������l�0��C>���wL�뭞�ͷ=3*��y�0SI��̯uS��=5�r�3U��j��$C�}������H���|O��m�<y���Uq�@�>8�w�\};�7�w���s,�W3�?�:TPg�E����J�Ф樞���lS�v54%j�W.��V�⬣�us0���ݽ����dJ�V�9�4�����ۣ��s��BO��B1�)wz:��:�����r�j���+ڝ��3!�R���7.+|�%�1�[m�Mƥ��� ��ya�g�eg327
��8�z��h��v��[HuJ(%��V�i��Iԇ�SxVj��#��k��\�{s�I���ZݠT3���5�Z���Ś:型Q㷁�k��P*���X][)�W�FX8s4�z;�^�%b�I��Yd])�o�k]��ʝoh8����mYoh`ԱW,�m3��ݹwI�C�z�^cǦٰ�63z[��v<�
�p�R*�s �0�FՃHE;VS��̈�̭�{A`b�i�rw%��ݻk�)s�Ϋ�'���[�r���[�k��{�3��7yQ�]c��8��au�P��#�KL�}��e1�z�J�k�nY���ˣY�x�ۯ��5)N�pnos4�]�$4{1� ���.�H��o0ʩ->���V�)nخ;��� �O���3�qѫb�H�ˏ1r�R�����L�h��v-}Z�o8�ا������e��K��,MC���2q�+e����ѣ)��W}�j�gf:�҃������#ub�MsK�������Ŗ�v�(tn�Ɖ�u��5��L��TD�%���R�%óB(�X�-�I��W�w�i��n�{�ɴ*�sR]��Rȹ��B�ܥs1ծӥ�A�u��L�4Bڴ�I��u����c��o1��a�0�H[�R�ʕ��4�0gb�R���`9d��)�Oچ�혺�K[���uڵ��Xss�:�%�j/l�]}���ʴ}up�3c���n�
7���t79�oX�X_)�>��M+�l|p*� Qu��u�U���z4x�.�L��i;�0�����3�J��C7����.6ɬ���Z����q�ڒ��#��(�	��`�E+�W]�q�8.��Pdl��ܚ�Ҙ��Ca
�N���L��O�#�/��+"W4�҂]�c'jt"��m��R�5a���3B�{Nr��s+��M<�d�Z�L�3�o-�Ûlfu��vK�m�?�����?	D���
�J�W\���R��g9�2ITT(�A��QCP�r��2�M�*=4"�!7��{ǄY^�Rg��hV��yAz�yR�eJ�����*	*�):��U^Y�f��d� ^I#�yd�A��!E�P[�ZK���{��$���	QX���%�{���Y����S��QzZ���$�B��$nEY�I�&b�$%%.Yy"Y�H���yX�g�y�YeH��IS���z�NG��BE�ae�R�'�jxXx������RB�E|�!!���i�I]^?#����ws�Ӹ�d�(�y\����L�h�:��3;<8���(����HW�߿,����>�q���qTGP4����5�Y�Yj_��g3`�F���ص���tk���zz9>cl��y�Ѧ4��u[7��n!, \e"��ǹ�+�$ϻ�<y-3��b��L[E�.>��^-��J���7��DRWEx�ԥ-3�M��w*���GEp�wh�j�e���X��Ԏ�t�$2 ugS�~ ,���X��(Ϲ���y�8v��l�»��9Q&UVˊ!J���.��ɺ�9`�({`����8�j�Soޝf^���!}abO��f;������ϲ�Y�O��nU@R��]�MQ��ܡ��n�He�B�k
GO�cL��յY���Щ=y�]u'ދ�t����lV�8�A��Qh�~��
3��z.�Ԋ9�;M�"ٵwf㟴a� ���^I��s^Y\�p�7�ԑ����u���:����(̕/��;ECK���C��V9J���u�P#$ʙ{�V wΦ��2��hT%�սk���]���{'>�+F1>ɼ]"ԢMn;&J��5'�$��],�X}&A�y�2X�'����Q����u�Uofd���%�V���,.bU?���)3;��	c,)��km��+ �U7��qOe)p�_����㶬/?��,�|��Â��g�7q�-�Kv.�F���Y�N*����^���]�6y���-K�C�\�~6���˱�Z���:�g9S~z�Ȼ�^��n�W�	q%�������FϷw�cbnvz�s�A��z׎�zޑ��;��yYgN�r�`%��]���p߅d&$Ћ�B�ڃ}A���Qp��ҘU(u}�]��bJ���J�A��w
�5U7��;���x���;8 6��F�_�}dP���$���GW���)�.4�~|EU��tp�_Mn0��.����Uw���q'R@�>#�a,>�1���53�����D$߻n���W�,�
�4 ����Z�9��Q�-�G������`�v�	N�]�o��(�<d����*[L�:�;Zٝgme%0*�,�q"X ��鳨7�����A��
J����hS�y���n��!�%�$���Rqbx����Fz1��[��[�rB3Ja���7������fu�:�w5�@�ؔ{�J\���g�s�k�.V���w��vOKt'#��{W������X|��r�=����+E�-xC�7�0��yH���wJ�3.�Zx.ma���y?I�����=��.k���>/R*�86�˱��2u��������avmdJ!��Ņ�J����/�!꼦�`��B�&�v��9'j��ƆY�'�Z'O_��r��BK�ݯ��/���Ⱥ�ڇ.rDv�uY��nL�֬٢0U4v}���B�)�}�	�_��9��Xӳ2���+�̢�Ot0z��9J����������y���T�|��Z���GG��%�KA�����2�OM�"8.���z+�G�2MyXo2��h���ȶ*ۜum.��ͺ������s��'u�]\�۰�g�f�fN���M�U�Ejn�B�\E��!�F��[��9ԝ|���^���స�!������۝�ق�Wf���M�>�;pzh��V˃]g'��w�R�^兦��Ex��i��nzn0�U~���^�3��0�z6�o�U#�oO�kG!��b�iqDio���z�h\~�������8�[��M��l)�bg�+]/#e$gW����F7U��?ޮH~Z��|�o����/��CWi����؞>����J�^a|��_���	J5��Zt��ԙ|����x]m���쓚�ki*���j��V ���K4t�$EQ��k�0�u��|�l��[�8��+֒�a��>���+<gÑ������C�����߳e߫��G�i}h���C#D���*i�����8א�;{-UI���V���Zi^��W�C�b-�[D:U������ey��ɣ����)ٵ��Og���%����0�>�Y��o!��֫�twYn�	]K���ړSG�t�	���֥��kr��Wz��q*�}#���m�F�܂�;:��jM�r4��d�ثU-CK�h��_��qx�B��Vͥb�(�M�{G'��ת o\< J���Ɂ���m�bC�{[;x�tم���$�}^�ңv�]&o��.F���dw�^P���fwm��,S��x]��v�G��R��������4=���b������jڵ˵&�fΨ~�m�lx�>8"��Z�#A�}<o�&�0�f_���;9ŦE�ήb�xk����l��͞E"�|�i���%j�h�`��	=E�R���s�7�P��A��z`V�`yq��d��ͤ!O��r�3}-��#}$�*�=JR�瞘5�>��
y ������{�Jͼ�fr8<
Ú����WH`HdB�<t�]bV���^ت�O�*�5^#�Y=��],KZ�� ���+��JzE�5 oK���=��F�%�[tA}x����ϻ�-��a��Ѭ.5���Xj靳��.>y����VG`��\��,�rє��("�..,��׷̃"�l�1�4�<�ܝ�{����o��_^����/�-I��zzS�^0R����K+p���������\�f����b�q�:�!��#1,*���$kˎ�|uUK����vizy���Ç( ���65q�Pq�R4~țZoѽ���g'�[M5��0��⨪�L@��ډȄ�S�ĭɜ��r��\&�Y�rOk-'H����1�r+�/���w�KT�*�=��M`���odЗ�*�bqy�T�T���A��Gg����vc���ǆ&�<��4�kdm�á���/?��E4�O�T{�'!�ݞCJҙqL����ˇ(�TVn��"�acg�~'�B��s���W$4�`A�ǀ�uVN�r��_{ֈ̌B�=3t�yX	q$�z�S�h����քlNI�U�l"��\S����w�wۢ���I������3Rfu!R/a6�FD��� �+r��F��cW����}�=GE�{�(���r��]��G�9����v���ܔx���wZټ�d�H��{�;��-���.�d���}?��ݬ��ėҪ׋ֆ�Nf�Y�GL}�O���[&�U�P4�;A�������Ҕ���ӽQ!�ۍ���R��@�f*8P��U3�"��<�')�S�Sz�xG���״�.����4^oA���mND�H�<GN �{*a�\�K�F�k}�#é��]��$�		 Ż3��9t,�7�Yw`A���u)ι��mݙ0�e�T�B8�)���
�����"���ѪkG>�ZW�8E5��X���b��\�o��3C�X����mK~}[���I-ԍˈiqÞ�m
'�.61���"�I�V`�X%i��A� Agn��ߔRڏ�\�����C�W4S��9�c9"��k�{W��{.�K=�rRC�O�1W��2!��=�T���c-�Z�6b35�mcd�YK�'j]�_IYx�8�*��i��{Ϟh�֢�((5�c3pp)�%#J�P�7n=d��U����K�pm��n���o��!������˺ξm�+��(���q��K��n��n	��@�]C��r:�R�˺뗞�nϾ��.�!�õo�h��㶇�Xp��H�喿#_�]n�o�3z[�ؿ
Ve���ܰ���Rٓ2����S��{��
߻b�k��
�)��#�ĝ����/|�.T��2�]Fv��u����%d�E�%�SR)��=j�!���J�[.���N�Kz���Jq���3�\}�D
��>!4�z��p�Z���~>�u�b�����v�fD,��NϯC�*�3�iY|	qDqo�Բ�x���P���+Q�C2}�U���v������9���Q�Y\x��+�<q�/pM��UԱ�2��G�2\/���ϧ?��)V����hj]�w���M5���ꯟ��P��3���:lZ�\js�L�L�T�֍��z}�#tң��0���R��՘��L|Y�P:C���EDq�g�x�鷆����Ajf�����f���!�c33EҘ�5qLtᧃv{f�bn�D��&�2h[�)��nU�����@��y/�`�FM�m[�;��7ܰV0B��-�W9��\S�!��B��(�F�n��3���¥��B����M򬌚q��#5؎!���F�d����kO�8�v��F�}-V����/4y���jb��kt��Z��
x�F����!���k_�*v�T��~������µ�(��O;�~�>�����g2��d3�w6Iۻ̿o�'���5ʆ ���]�����x!C+�����yj^�gyy�Y�ż��[�7�.L�vT��{�˘ᘬ�#j�`�dT˝�
��Q��<$4�=�!�"X�ߧ�(�����_J�i����>n���b� ����V�_W�P�����;���!~0R��.(����p>Dfnӓfg��ř]���o��\��%�2t�2�?��c�󸺃Li��i�ί:��5Y���[A��`��;_jc��mcet���[wC�`�Pt�p*Ԍ��'n+��\]b�ӗ��Q�Q&"8�x�Ո͞�.�`�Q��M���ټ�+֬�u������w- f��=�Vd�
3���^^S��}�竮��*K���þ���7�* G�҂��'�i�;V���o���79`��zK\DٙUS���i�2�خ�`r��/F�'�]���Oo
��q:MwY����IŮKA8��|})���1�t���
i'�s�(�e�%�
�困7���0�k�/$�Y�ZWD`uNo+e�;2`��[׷�� :�|h��0r񾌟B�iP
S�����/JEF�ŏ��ve)q��w��9x��$�_w�\o:���f#��^/Zщ߮�$����ղ�6`U�fԪq�EU6#�7n'��_WC��N���j`�S������Ϗ�5�.K�yW��I+�'{�^4�.j�t�cq�[���<���3�sµ�,.bU1�;~:hm�`�G��%p����Y��JL��.x�?��Y>�,!Lsq��ѭ�ż�nFy^�]��u}�����Ȩ��<,�,ٖ��V��R���ő�u*K��,u���j�y�{h�2� 4�_{udf,��y�t���aИ��`�>w�_h<9�,,
�)�=.R��w���)��0��%[�D#�H�w����C�1>S�5�y���i�%Ԙμ�1���vy�V�t�qƪ�+�&�7�R��%M�R�ɦe��on�l��s;L\�bT�#Xr��c���Bc;�FRuE���������M�$���k8(OY�l�T%R�(�ǵ]m�j\�dy�B2�����`�{[*\�B.ҹ�]�V�3+�g*j�6�CF�YC9���ڽ��]�T�44�k���ïj���˵����xf4����Vi/��+�,ǳ��#�ʹM��sV�\����=$��)&�L�~Ѣݻz�,������X�ۗ5q��&���5����&���>��Jw�c���q����z<q�0�Z	^�M�g��tec��v��5�.BsWz�s8u�߲��,=sOAn���`B��5"j22�%/��Ę�sG��Ƕy�[|f��o/ޙ»*�w�L4����x*��u9�bQ�=�Ξq3����9W �۵ᵓ��D�w���+r�{g\咲��y]h�BڼZk����/BΧ���e>k���0Iӱ�,��^G3{��d�2o2mW[KC޳��7��~U��W�;(�)n�Eq�-�Pv�+�u���R��WPޗ&Z�o�P���r��Ͱ,w�`"ewnP݋��BN�šHk.l��L��[j�T���3��Y7�X/�ׯ_mi8� ��2��eIw7z��|Y���Dڲ_&�WZ��G*�
���q��ǿ2y���̼�x�g^űtu�լ.Q�B'8m�QӤ�m��Q���eY��9U�j��ک��C����9{Ɠ���>�\y��)3�m%�z�Ы��ɳBf2��Jڪ�8&,��#gecKU��a釆�n;xp�\�s�s����y�jU��Ce��Ep���ۈ@&��:��/�qp�(�m���X���ܡY�eϐ �A�!T�
�HH@���D�*%2F����2B�YTQI(��*���I�h�o{�>���x�f�MN��Fn�P�Ih6�#u3#��+R��'.��ȷP���H�/4������r�HR�2�$���C-�ʈ��2�䲤��]Qu�1<�(,�D�/#�:�xTd��*J`�*�^.{��(������%^PUTg�k�3�h���yI�VII�0��yB�ɭ��,%�J$�<���u��8����HzI RA ���>�]�{�E��}U�λ�S��T@�YE�I�Ѥ���WSGk:5�;mЮy,��O/X�K�ڜ�d�2�Y_ϵY�lz��\g����k����j����=�=M{�n�c����c�%ԖK6R}�M�?c�,��Υ��{���w�~K�q���T0�ŭQ��_?Z#�F������*�<���q��y��Kj�%�Xs��j\���T8ݙ��S�1�0�]�5��㛷���z#1qd�9��%�~$�N���������,R�;�C�V���������*0_8z�OO�O\+��Tߵ[[*Q��[s����Z�s�;hz�b�cL�a"t��u|�t����
uҘ�䛮��F^�}Ω�	�Oݰh<v��M�h��������E��������e�������N�C��fpNZV�ڨr��A,�D�wWt�
�������sQ�0��!vPSj�(b���z�=E��|��sN�����)�J~�n���iۃ�K9���O[K${�N,��������u�ב���,f��l�GXc���et; *�T�˴fH��:��A��$�����"&e�0�e��t��6�噹����}t�O�ӌWF�;�1��}��P򅌬z���޴��A�
��I���8�Y��k6�ʼ��$�FÓ(k�*c��۞�����ܨ��՗\`�Z������.4h���s�=�7m�y��s������Nv�8&ST����Q�~~#>�qŗ�|�ì����=W�	~����CF׭F�eھt�4��V&Arj���4֦| �+�>�^�%��'��6vF�J��%*���}|7�o.�5���Su�x8G
C�}��U��d3}ic����8.b����)<�v}�R�N�<*c	��F����L��������H�ڷU�f������694�@�MH��eyh75�����%Y��#p]t�)tx�~|����z�k��y���W���98�ex�N�Lg�p8e=����dŇӥZ�k��t��r�cg��iߦl�{iv�p�r�sL}�& �jŜ���p��zq ��4W�5M8�D��:��nǚ�õ��=gG8Y@P­ԓ�r<����KR�3��$cb�X��\�Q�o�t]lX!��`V_o��	Ņ�^���ItE��Y�&�����[�9.S��cp�13�"!X�X�R��y˽�J�����,��/�m��X����mWM���]��KZ')��.1���|y�P%�ܨ�:|�z�!)@֗kyq�ϩ3[y=.<��O[F��lzuD�J�ǒ�ܦ	�"��峝���G�U�<�]��`*~tZj���Hn�ig�_J���Xn\�9+:���<��ٗ��+�&D���Z4�o[#N�P�r,i�jbL������_f�N�ݜ�����	>�(�qh0n�ثW�B���3�u��%���oU���KK�L�5�+���;�Y��\i{g�3��ͨ�4�}������ؕ7���w�:��\�"���et�]���*G�s ���>��E��s�yF��=~V./�+KvR=�T\8�7I�БyY^���5v9.m�<v��b#2���<�"�h8pa�<�]��Į�qN+A��q�15ݧS٪�3z{	n܎Q�_ p�s��M��r�C(��ǥ��1Y�F�����=[m�iH���Nzb��{��%��b��.[��c�'�X���d�΂S��N" �C|��:2��]���J⋘,!���o3Ν˞�<*�ؗ�U��R�9s�;�����`�&��(v;���fp7^���Jf�!P�s��B��e�|���P!�L���=�Zn�|������Y�w|y�Gcy�}�]-,	�t�շ��?{�y�4�~ľ�������l�N�t_�JS��F^ %pr�U��ׁ޸k�3y��N-e����'&��@@�-y.�O�0���`��Q�s���v��_v��ֹ��.%�=I��޾�H0G^�A���Ո-=��vj�\��E��Sđ{2��o�u[�~�~���T'�I�iT�v��9Nײ�V��4��I�Zm�/x|�m�D^vH	h��4��R@�uEu[�Q��z�|������ ���w�N���
�d��>�Z1�et��]}y���R 7����q�.�ӄҮ_i�+��hw���:1ǡH�)�{kk�s���Bi5��DuP�y:�O�a�y'C�S��Nvx�^���ˑD���gEJ�	��Ŧ����ʼ��$��	����g"�G��7�ͳ�{�Z�Rx�[׏܆��c�1�|��魷�G��3x��N&y�
f�Z�31mm��3F�1۬��㸰/?���%�H]���US<y��ga��6��������ݮU��}~�nȂ躗Q����[���"�ɁUq>���:M���h˗%�v#�Gb�w���	ruR�ٻ�T�j2Y���bkR������&����Jc�0���O#w�5i�7�n��G=N�0%��z5x��-����_�=hl��Z��#�ʻ��بX�B��HY&%�[�Ei잃�xrG/��Uk�0�'��ݯ��c�D+X��q�n��\ye3��+,�4m^֜Mp3�ʞUq��R��z�[*Y�.���Q�#��17P����:Z�1qXZ�������$�#��V8G}�*��=�'ա�aG�"t�\�ø#�\i���=J+3�۽���J#|-��N�}������6Dg��_�i�a��L��Ak��^vl�tE)`�ڗQݡL,���r�3���}%�$���<��ʲ����¯�1�YC���E�;)>#56=�ԝs��V�ۥF�|O`����~�%����1-#Z�8�F���yS�2�������H��r�/^����u�:�I���L���͞����ux�Wv�L�\N�W3�ؔ��؜5S�acd�k.$��֠~b�/�."I1�I�)-m� mM
�pD>��FC�3W���2��6���S��U��#{3���re��}���CC�E?��(��u
��J���˃��d��V��8��v�RRq�-/Q�u���a�ܮC��h���]v�s��f�0��$�gd��:��[�P(�{tN�D���Ѡz"����n�mIS���o+�Xŵ���z��I�7�R�����kv�wrq*=8u��p��Ll�Ư����'e>qp�����d�b���1���5�}�����r��k�,#��8���1̙�P�����].�����B�K7���,�[�N���1�����<�3;&WD.�FM$����f� Φ|t��k��VԊ�ʃ�A���v��磌6d�y��˾òn*��V��O��DV_B:�Lg�I����N��s�/[/<�˟,�1[�{���U�9zb�CH4�+�'���n�GW%z&b�5��8�����RU3E�
{<��HV# �'���s2���
Æ �:����:}}�@�(���=!+�ʽ�e��\���	�z��x�.aqM,t�����:��s%�(����Dy�=��&���9���ͨ�y�J|����v�'��ɢ�<v�a&���d����W�*cb�kW��ccI�^%�>�'�<C!?!_s3R�n��W	�ɶ�Xvs)J�!�d�ā�w#:}iT�����S
�S(�h]�2�#���NKt��Y�h���6��V+�e�N ��ݜ�J��f�Fi�	�˛���NRآ��*����ܹՔ�o�"v֍!��"4�%�GO�X~�����޹)��2q��|��cgE����/�V�8YG�j4�z�=��7���yX�sc(�Xp*,��9�v��
��"d({K������d#v�׹����;p�D=:6���*�;���Q9���Fv+uGMl%-�Ϛ6�*N�������Ʊ��L.v}�Nz�\�V�U;Y+E�� �򒯒��E�y�g�b�����g�������}�z�X]ӻ��F%��נ`�|ۻ�,Cڃ���"�>�2>���}7�q@��	?���.��׷��1�� �%��.�Z�q9spC���l��lX2����,w���J�e��S�բ��T9R�v
4kA�%3ns�7�=�Vd��T�8V#�������R�کqԥrIq�F�ԻJ�<v�����hj�W�}��]�{ad��ɩ�ܻ�\���
�.�û��8�l���Tkd���>���e�g8D<�@c����e��+h��U�{pm��yf�A��:�rp��Ms]}��)$<T��E�r*�|�)j�7�X�,��N�Q��	UPn�����Ϧ��7�u���4�@ݾ�Ͼ�(kh��K���Pa����Ҟ�D��J��=���k�DNNK�xz�;�ۣ70�11^�T W�2�<{�a��i�<ͻ�5J\et��ᝠ�¥.{��\�*s�uB|a���ZҔ�v}�ޚ'mm^������Ŋ���9N��Ǘ��������4)��A�/�c�˼��b~+����](���B ��7Q�ϫ�I{�P����漰;�c4�ȼe�snod�Y(���Rq�����H��jc��'�y
䒱�±B��>����W�H(��%�]juI�C��^�c"����4492r��zS�u���j��@V��Y	On �ju�c�.\Z�!�-\ς�w�4��ς����{r��~�b�F{F˶�6O7u&u�u)�ݽ�fMA0�uKg��G�K{[����݋tv�ѡ��-ނXϢ�Y*���D�4�f�J��Ƽ�V���.�����W�fj��a��j��,z�U�fV�ͫt/h���3�]NW\�KU��pcQ��_4�\�7�.N:<��u�F�Eyp��s_��CW�������8�+/T�_Z|�Е}���3Ԡ��<������d�_c��+]t�;V��m4B�p[WC7E��ܷ�I�%��ބ��Ě;��Z%�w�έ]W�f;陛ڮ�b�e� �e�t�2.NxP2����j�{P��t�e�}ĦP�o	ȸ�;�`>�栟P:ZD�$�����hG�q��y��ǏCC�� ��u��6�_�S�l�D޶��KO���Ɨ�Uy��̸0�団9 ���O�������� ��]���9���MK���8t��Y��(�;�zvOg'�}���(a����t+<}��Z�^)�����A˄��`�JV�s8+��73II��R7l�������1)]����iSF<e�Fܕ%������[;1e�v�Xi��]��捻���_Tk��D�H�I�ǮM��?��D����ލN]y�[�_��5�K���.�ڸu�(4�8����l5.+
�s�NJ�b˘���J��|خ�.��x�y��|���+�ٽN�_>�ss`��t�	��|�`��c*�aS0��y�;���C�b����&�S��,��u#�Ⱥ�f]9aI��u���A4b�x襱�Qղ���6��X��L	�=I�d�.W�iB�46���wO�����٢���N1�L�|in�;,s�����j��RQ���$��zT)YƮ��&#w�5^Ex��I� �}§	���&k�K�ӹs�#֬uh�R[A�=t��lc�%Wd��B�+sN�	�ԩ^�ӯq�'s��x���;\��n�?.&���Ȇ��x���.yW(�9ή�;]�f �?����d.�!���v�}�ƻGkqT�ۥ&q���$�0(t�:gp�'Z�O�LLs��iM�;D��[�Q1em����g^����T��I�
�o=\�;DwԻ���#{$"�[U�Q$���l��:ݭ�����W$Û0J/Gh��{����'Y`�h�Yk]֜l��Vt��M��T�sk-��M�7�����f�ҷH`�Wl�a�S�GJt�X�,�/Wm:Gu�3�l<��t����X���]X|)��*�x���-�9v�v��0T�k�/F��C!��n��C)*gq�fܸ��ڈ�M7���x�$���sW*d�j��Fn�93S`����"�s�;5�Ble�t�� C�0�7~�܅,��_-o�̃U��.jcݹ�w����_\��o8K��ʽ�y�M偏�hӂ+ Y��%����:�Ʈ��F;�,��[�)GHorÜ+������^�ۦqF|�
.\��_ht�H:!��ߣm�g��TKe7�����e\\�nTz*z���<��\3cFr�R�7�j�ed[*9@�Ғ�xk��	���v��XU�b4�œ�6�%}Ν�w�:��Q.�3�N�n���*[��ZB�k<,�/Vtm��r���ϰ�U74T��֢E�E�������W?_^��ϩ\�5�U�/�M�3�Ap��f�k��ϼ/����FcW��z� �M�T�����"�T��zy�<���"��+��ɞ��^�î����bM\j;"�
/HO0*�5�O<�/r��ܳr�0�*5Q<�+]T�Ih�"kn��e���hG��u("8��3�
�DXѰ1t1+r�&�*�R��5	!�����2!$��&B�Ꞅ��fF��qݜBT/fE�2mr&M�啓2.�/쿮���S���㑗��c���׸kE�ٺ�,����q&��,C�=�
��Q���@��7�ML�˛��؛Hk{Q:�=OພjnhC~Ņ��i�ަn�ٖb��dB2�n
Ь��z�HʕR�E�Uɮ)e�����{Q]^Quz+�h��1c�����׻6��i^WT x�Q}F�n/#������|����*���OCo�+)c�CM-�Qq��Ҕ�[+�Lm�8է՝�{� ��b��vv���S�ZLu���Ц�'S�,p�X��`��T,Gl�1^�Y0+T��X�+.^oI|������\���s���Ǥ�Ř��"3�ĸ�Vh����յb�2�צw�Y���NUҬ�.+A�}#�S܈�P4�+���(����/E�R�Gˁ��!n�=Z�����<�閮����,`�Wy�O,�c`,Cy���'[I���n'�8[�z�1�qM��jq�\�X��M�ջ�*�C�/{M�Ŗ�IpI4�'f#��r�ɫ�5g�˩�MP�Z��
��������kHKg	0�1�Tq3ՙW�6$d�/�5���N[E�
�a+���cw�Ȣ���r�2 a�|�j��Y׷�o�jKvѽ�+D+�S$�L�����C73�d+/���]��^�OvxҲ9f��l�ʎ4%*ͦ�i�{��iE�5���)�w���M���wO��'��蛇��n+�� ���-Eq��J�{"��Ȟ���V�Apo����h�ynb+��c-l7�ol�0����a(�����k�ú6�߶��Z��k�F�0���<�ejO�n�a��n<��xg���=E�Â��z�yӭ�ќ$'�Ukqy�_8o	
,;��È��+6��!�*�l�w��n�$�x^��^W��	��%�s��&\�`�\�-V�%{z���"J�x�ts�jB�H�0_��EN�E��nc�xx�}�roK��m� �(z�%3F+�`W�Ҽ����I��Hu'�����ۗ��bT�XS<�|PNE�3����TY��͔�s�_PV�s��P�f�2V�0n"����[���r��v|I�M��ʻ�H�&�� � ��K]����V���N54{$�խ���J��Y�r��+�OǜIs1U�T9�	ck�{!Q��P>�6l#�7-\k��״K����oR�V����)<&ʞ]��yL���^��ev�$Q�S��t���K �/E*�+��Vq�-����f�u�^Eb�U�0�,̵q�];�P��`:�H��T�M�+��\��.�2��q۷RS�쥤�Vհ	����0qr�bRu�F��N�Cn:2�U��DS��V���j����ᾂeiԚ��0�*�g8�rqC;��F�t0b�����S�>2������@D�8�4�n��;���㶤��� k70�gE8�3V����8����n6־�{1\tY}����m.�=a��_���{�w�p~����*%���n�zK}�3QW<�XꃳƥC�Z�g!1��0�y�0�I��i��g��V�Y�����\bs���u7�n)_38���Z��X]��F��(�J�Z����ǫj�ّ���*m��6���\:�A��s ���q�g�i �1Ŭ{�w�HY�P��:���G)����Y��9��"�c~����s�Q����Ĥg��Z�ʎs�]�+���
p���k,�2��z�+�2�����麒!X�u]��禛�����?n�c���j�=j�mԧ�V�jv�^�1�\�k:L5z���g326�f ��q�@Q+��驨H,BNh���3Y<*&:���V]��ty@\+�i/iL9/���<��6�%~]+c�|�-����2r*ŽEl�87��&��_�D]�s~��������uyxn��l%q���a�U����YhJ�gs׳��
����`�oݓ$(x"�;w�U(��Ku-'����=w��3g�O�OY�z�F��_�Vŝ�*Y$;�ͬݾc���sLN�[k��/tk������ɫ�:F9W�	���c��n3��Y�v�$b�z���W�Iy6xv=�CШ���h`0��1��	�qn?v��muf���vޚwe�bN���c!�s%/F;��Y��2���9:׺*E��b�f��r]�-�~�\�W�͛2�^e������:hp�|O8�(+��9�����^�YE�O&��M��$�}�,���|.�������"jo>՞�?C�BA�ȃ
��'e���W,K����U�#]"������Y��=�6�s]%ɻ���١h��ZW�ux�t!�g]�/U���\a�w�G�Tn;2u}�sg���:莺=#{������i=🾛�ZIo5�i�:z��*9",Z�[K��ﰫ��#3$q�������Ab,�|��fWS��u�>��!��:�wT�=Bs��"�2�9Y�|�����B}�<�l[�ڸ���6��Aó���v���{{<�%���W�~�x�r2��	��zU��-�������t��Q!�5�,c��L�du�������^kz��G����ɴU���!A��E�]��t�����V6f����a�7b��N��4K}����C��-%J�|b�z����Q��V���(1\����&�2@u�ۆ����Θ����_o���f�����U��*����Q���=��=��������}�뀜��������7֮���6�^���=p���;�M�b���mx��-�n�+�3�x;R���w!m��Hn�d�c}������ث��y�����{�L�Z�������.�
��_D�qx\��|N�7���u�Ff�����{%�3����L�q2q�ӱ��䨞�Ը�Ok!��kD��s7TU�"㽡�82#�f�X��Ʒ�XS�S+ψ��f��YLO=�{hxi[�����5��?Q��`�}�{�fPH\xP9�{��W�.�;+ `�3�ﺉ��L�g��H�A��pF�˓��]��,�f:w��
��9�SGx��G������.��o�m��Ú�b�v5"d�[���ün�lV��1���(�w9�hu_�ЙEyr��\�l簄0x�g�A��+�y�]Z�Phl�n�ۊ;�l6�;B��>�L�Y�׏��$v*|��C���<�d66:2$�A��ْ�m��2G�s& U�B؋�Md�S��lbӭ��W��k�y������ ��w���o+$^tT��.`	�$�a'��ȧ�6o]In��W��n6է�Ұo�,e���ϟ��x�V.���9�w&;O+�<��^?^T@��z6���[��n��z�����h��Лz�Np�^`,j/MszZ�-O�C��w��56�m����"�%�j�5��r��.{�o٢g�<;s�`,�?��3�3:I�Ib�4��Xͽ��=s���v�z��w�6N�:;-2"wk!�T��f���t�Gxs�qL�}SRc]@�A�)�s��۵8��bN0Ҿ�rF�v.�EM>��,F,f+���)�Y$�;����m�bÁ��h���X5}jZ�Qo�wJT�n�l,�Y�ts�����
���S��6-Ȉ�w�6OFX)��_{�3���̭/i9�i�PD����\�J�x�&�a�t���%��[˫AR��z���<p��S۬*��o�����Ƙ��9҃��2T�N��=O1m-]y�V�En�r"��=�m;j���ȧδ��T��ͦ61��N?���|��	T�9��6����(w��Ψ��a�>�왥�y������/n����Y�5"/��Ҷ�Ьp�_��eA�E��U���d�3A��gFQ�u�ҫ�'��D�f4�C8�'�e����\Z.:��S�j��v�%b��n�R�숭�v��P������{s:T&��7�f�@Ÿ��	�i�{�5�I��Ұ���>��s�걆Gq��2�&�{$3sb6�F�Ǚ>�F����gar��$u�a��&��f�;�1�l:]�ӌoT	�Pb5R��1�u�%�(�άv�%ͽd��ǳy���S�<{rq�=l{f<�"��~����|<aT@�"z�B1�+��F�6n�^������S�w�pK+�I�#�ݜޢ��n��lRs���e����m�D�q�oRkd�;:"I7HStzF'�k��W*T�K����%mds1�B4Ɂ�S�Qv�"O]�wx=��U�h��Swt�T�O-��h���5}�V�&Z�g��w�oc�������Ҟ��WJ�����b�$b��>ȐG�܋M� $��WYQJ�j[#�0ш�U��(Td�/�82��qi��/GK��r)b�TPE*�kHI��I0���]��]�BB]IK_�<d�!l��rd��2��!$	 �HHH��!L		0�$$$\�����!!H
(��(
�_�ٌ��wrj	_P�ЁA���%~=B��)j�R8~H��(DPT�T�J�UN�j�V���_-�p��X�p�FEə���
R�I�3�˭2�d�����?L��M�A�h,�h����;RB�j$��P��`���gΚ
�
H�h���7�ysv��U��ZMpw$@�?R�ԇUBB$�~��
�\L'x��e�M�g�'��H��ro�?Y����F���k���5�I�$�n�z$"H�r��H�����zU�C{7:FF�̩��F�{UFjF��\㮾g�B%�����O�����8^ у֯F��>����\j��,G��M%�U^O^�4ZH	"�t\�*3��Նt��e��,�	��
ڬYd1��"Ȫp-Y##+)s37���^����ך�H�{���f�e�$p"�4P�IJH�H��$QRQL:����p�'v��c���5��Č�x�L_�๰h�Gܨ�8H�t9H���p�V$���g�������W���4�-�ܔ�B$��X���u%�bt4w#�Gwb8>�hȷ�N	�M�6�v$`��H��ysx�N��Un�:�G���;�����8�q��j{OO��������#t�6q��(RV���iE�����fk0�?"X����T��Uӝ$�"H��9�B$��⟉�|jG].UZ9026<��C4�34�F�T`���y�S� �4M!ŊQU&�x-�i(�5��4���$\�5ɚy��'S�֓Pɫk�M£F�ݥ#�cĦ�$�M�����<Rb��@���r��$�n��pʊ$Qk�U��{#��7�u�Ӳ$^i^n��yI%��Ȏ�r�N�o�|�t��t�v*䓚p���9&\ё#��9��������
�u���z�nw�z��8�I��1e'�G���m����\$"H��N��ruWT�R�Ҋ�h<���6EO\$"H��ٍ�����A��w�q���8��r$Â=s٫j5h5Ԣ�HT�S���
T���Wk��"�5e�t<=[�*T�I��#fɛ���uZz��=ۙ���k.R��dw4��Is�4u�CL����S���.sj3*yj-J����,����Ro�.5�h�Sc4d��*y��V�+�7#�D��G�%A����F�H�)�σ�mm�;�$@�:��=��MI����֚�+B���5�ل{�mR:b�S�ˈ�W�(O_C�I��j��.�p� R�R