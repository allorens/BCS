BZh91AY&SYZ|4D�X_�`qc���"� ����bE��         ^B�J�
})�	V��5�hjT ��@(����*�P�a�U%J��S �ғ`%���-��*�6�#mm�:*�k[n}�
EJ*��UQFƽ�t�
%m�U��	RE[*�(��D�
ي�J�[�������UHQE��)�P�U�3t�ki�*�p���m"�8:t�,��ĥ���mH����Tk5��{r��6�*֐RUP�*Z"�z w%U*���     O#Y�GN�DkR!��EN��M1sV]�
��[n��M���,�;uE��}�uP�n�R��l�v���4�QKmD����   v���l�e@�N�
S��*���w�����}n��ZR�om��M�{e*��x_m
U�R�����������C���w==��Wg݊���=��_>��PET]jFfUUUm�   9�i�[Oo��oz7�>�u W�z�S�@R�_o�u�#j�{�쇠�>��{{|�ҡ�ҧ���QJUE��eR�z�Q�����J�̝5χ�����|�@����BSfH��   	��O��J�O�����R[��eld��]�z^�G�m�y���C�_*�=}��h��9�TUQR��@�O�������{�t=��J�����Z*�!B���  �4xWք�>�m���>�$(s�缩!}��|8:U(�n[�ŭ�Ԩ���uJ�//k�9J��{�oO6�{��wko��T*R;{��PU_m)W>�$"V�T��B�|   �;
�^�HB��qr�*���i�)Qn�n����JH��ks��=6ڪ7GJ�=:�=�Lr�+�j���������z��*�x��*T�aEUDkT�   9݇G�}�	�Z�t����\:
�n��� gs cv��t��:e��f���c�����@wN̡R�m�����|   ��4{�p�)�\p
�wG���=� z�{p��3�J 6uq�mGWp�ס��  l���I���"�A�  �=��@23�  �t����
:S�����q`�ڌ�{/k� Ѓq� �� �;jT���B�PUB�7�  �|�F� P�+� ��� � 
l� �� jV ���8��w�   P    �*R��0	�`� #	��{!�R��&&`i�&#��BR��� �    ��A
R�13Pɀ# ��&􀊪��     ��zTHL�2bG��0���1>/������8���1�4���ey�7��S����9����߾�۝��_�������ࢀ���P@U������ 
����O���������� ���UW�t U���HD/�P �����?�����'��S���k&�kkɬ�ɬɬ�ɬɬ2k&�k&�k&�k�k�1�������ɬɬ��8���ɬɬɬ����:Ɍ�ì:�k�k�ì�ɬìɬ:Ʊ2k��:ɬ�����3��ɬ����ɬ�ɬkƲk���k&���:ɬ�ɬ���:�:����2���k������k :��2��� � :�&����k*�������:��ɬ��"�����:��#��� :�� �0��*k:�&�)���*��$ì
k"���)�*k :Ȧ�)��k:�����Ȇ���*k(:�&���*k������kʦ��*k"������k*�ʦ���+�!�
c :ʦ����k
¦���*k
�&�3(ʦ����k�¦���k :�&�)�8�k"��&����k �����
k
L��
k �Ȧ��� �*�Ȏ���
:Ȧ0��2��k":������":�2� � :ʦ�)��k"�������
��k*� �"������
k*�������&�)2����(�*��&�� �� k8Ȏ��� �*:�����  �.�
k*�(k
�ȁ��2��*� ���k ��.������(k �ʎ��(� ��,�k(:�.�����":���� ��3 �Ȯ����� � k(��3
��!� ��	��������.����"���� k(� �®�+����+� �)0���D ®��k �®�0.�����(��������k*���2�&�k�k.��ˬ:ì:ˬì:�2k2�.��!�:�ì�2k.������ˌ�ˬ�0��&��k!��0����k3��&���k&��c:Ɍ�ɬ�ɬ�������ɣ&�k�k&��&����Lɬ�ɬ:ɬ:ɬ��Ɍ:ɬ:��:��:ɬ:���k&�k&�k�k���ɬɭ0k�k����&�k&�k��ì����ˬ�ì�Ɏ��ɬ���:��:ɬ���k3&�k�k&�k&�k��3k&�k���k��&����L��WA�q��^�����7؏�fX�L�Ge],�
h�If��o���Vw�b�dl���9��qlH�{�z��K97r��Ze��B�&ٗ$z�y���hn��x�Z�d�nm^HM���V8sL�^j��Ʒ�[f�,M,,�o^F��ǯ*֗ �h��)޽K�V�`�6�lSPŹjYh㌭����(6o��<ݢ�v	O"ET*��P���/J�Rg�{��j��͘��;�tp�z���˽���Ɛ�5*̈U�zbe�G[�xN�12�S]�h�]BZ���d�]������2��\YkAL�D�o�[�>un��w´V��Bgژ��+�S{C+.L� mm�
 4-'��׈��ۙR1r��VȈ�2N3��7����k��4�H��*ک��J!0h��&mb%<;���X�ɷ�m��Cr��)Xp�@��� fm���&B�*Z��YI��W��1�p�*`ɒm���dF'���;��T��b�`��X9o�R�n�/b{�,d�)EgS����W��%�$���l?�4j�	����˨�ݭ�mK�j���� a����6�&�XK�c3\���l
����-jC6�`��Q6�K����������;�6P� �h��۠aC�v4��'��-ٗ/�OX�(��Z2+�yK ;bɺͼ�u0tf�f�O0e����V��b�x3bB�Th��AJ-b�wN�<�oQ���Hvq�jݝ۵�س�~���m'�%�;��-�q�3R�Gn�Tӗ.ma8�]��v1m+�{�@	�{��L,XCڴ�p}�
I�jӽ�[���ZZ����)�-�!�sr���\��6��1�+YŚ�������vƸa��Ȧ�"��u��j�J�*8�����Y�ܚ
H��ha�+)�ܠl^��%:kp"tҢ3�����pi�uj�N�Q�gJ��R��(i
�@1�`�S��
Wtq�^H-ɖ�m�b��Q�"l�W;�Y�	��r��ɨ���f�A�Ca9�r�ຘ7b��ńed��f��[w�37��k���Q�ƛ�n�ݘ��{�h �X��"�T4fS;!hKMݜ�X��T�fk�q�ӡ�.��A�h���y(�I� -i#k!��b����ci�v�%Lˁ(���B���X�4���]�Om[�̅�V��l�26�hE2��3r�#�v.�f�Q�C˗,���y7��îO]�j1P�o�ˍiq�m��h�0��e�>I�w�����������	m��]�ug�%�mm;t�3�L��R�,��(?����IordW+Q�;piPͨۣf��ْ��2��;��U���.(���k���f�(˫;�����Q�r��7�(��P� �ep{\�.��N=
ܧf�>?q8�Ŵ�>�'.��17u�P�t^�� َ��:�R� �W-�S����C�V!!�2�g7�_CNX����Ֆr�<EkݩO"9!L�.j��.E{y��5�A�bB,Ao���ȡ�p�)e��Q�����RT�F�H,��ӉeMd�{��?��
�M��S���$�;2��z��^��qݲ-(��ړ͑H
!�9��bz���<��%u�9����V��Aő�oΆ7�1E�)�B��ڱp2��ޖ�MV��d���>�w�M�h��l �5���i�j%��:�ـ�Z�w��0���ޱ�2��Q�P-�,f�8��:&��3j-��nT�V��]�m��c2��$kP��zo"���b�Za�`/v@���hh�N���$^E��e9FQw�L2�5M�!E�-BiA���Y�{���Yha���',k�a���e73e��Ċa;̫��:r��V$c"*V��k��+�-IwB��[N���9W�[�UAgB��[�>L�e��Β�9�V�^e���H���u�\�7.��)Yy��2"�Ӕ
��ot��V�RI��əOZR�Q�ڰ�ؚ6�b��O%jJ�/��r�6E`������]l"^��ٌ��1�(b6��Jg�]#[�.K���8P�f�Ky�];x�f�s"&�Ƥ�("\&d�L)���K��R�����7��6A�/0�劆^Pڶ�.=_B��%�q;+v֤ݦ�n��m^�0+����u6M�!m�`��!��r:N�=8�j����������:{�9��+r΂����y��ت)CH]�#����,/h�!���O��Kirܽ���h�Cؕ$��b�mI�i�d-����0��;��&�j�X�"R�y�U��3���*�wy&	���M팗b�P9�:d�*鼚�H���oӐJ[>ddC�n�A�aZ��4怦����,�ַN6�>��v3�-��MӔm钘�f���l���f*Ô�iٌ�=G�K�r���Ú�]5��Э����ֳ���)�K��[�r��WbƓ���,�o�[��-^�̥{�D�:�l�v쑦Ȗ�f�a�w�%H�.	���D����M��Y�.��T͌[n=�Mӹ��D�@�Hnn�rn]\t�	3u���ٚtaDkIf�#���L+k�%���F��ST2��Hbǈ�٢�e��*˕{Yi���xk9�e *��q,�¶�raj�|���p��V�s�(iL�4�	�^,�s�2�z3>�6�h��+m����M��4�w!k����v��xj�,�v)l��j!z�t=	�n��tۨ^�剙n��6�6,�"f-��UYB��X&$��ۑ�w������GM��c�����>|��o!��`�X,�Zl�#-f!lnZ-�E��M(1Y��wE�jQ	m��2����֠�C �n�ȎV�gS��e�x��9c۰3��Ƅ�ǡ�}6J��S�B�d�6�ٸ�����n��ڠ��,��TnZ{G<	�����Ňl�fٻ�l�ң��;[آ5�Vo]e��3�b��t����_�<*���Ub�̖�J`��	�iB�3c7k���U�2KȲ�95f���m�\���(���d��C��7�1Kpd��mĒ�n
Ϭ-'Jr���4��F����'�12F��:��vO�2����Zv��gl�U�I��m�Yqe%��Սݥ,���[Pc�-ѳ���פn�
H�ӏ��(�m��Ð���t����0�NƬ�a�K�zu��hq��v}j�����i�x�L��k@gV�2i�cVa'h����Z�L���E	�K����.��z��>�)�$�/4 ��I�)ݨu��f̳'ЬH�uq��i�x/9in��m�X�fL5��4=JĽ�[ڍ`��HQЊl��Z¬�t@�=;�L����(3fhm��Rb��/m�[,����E�
U�H��Tؙ��/&R�yy�ڋk̓�,u.�5�Yb֤m^��/�&0yn���,�c2���˼����xq!����Ց�i$�v�P��e�����sai�+��SY�J��%��xn��ͳ���.�Ow��U�4(��)�uH7�&�91�ᣔ>&��9V]�Q�U7-f�n���܌�е{�S`�[Z�Ac�P��4����=�$�kI������V��o�ӉM�Ht��\x�o�X܁HNM�}/>Ca��y���%�m�_�m٠�bc�wh6�j�2-t�X���kX9��L���O2����-1�F���#o
�w2��T28�[pM�rhI���4Yӎ�E�̵*�����/21[� 5)PȨb�Z��K���6�a��^�o*�d 6��3�\q��_\���%U�1jMѦF�����qY&��"<�f[��+��Ql���	q�w�vMkk1�hd9���+m_�شЭ�0�*����#�1aL��wbΥ�⼨�X�6�m�*mnm�@�Y^�1�,��T����[DQ����r���[/p�'%����%m�%bFd�6�1�u$+��.��lRGo쭰�i��3+�u!J�Y(��ee�W�r1��e�;�&��f�0"fH�e�I�v�ma8�Zb��^�$�5鵕����Ke:���[Cl�ޗAw�V�cp��4� LA�j�w�������6(�i<�EĞ�n�Æ�$���FP�֩(N��y�_��1�̨/��h�{�!5�Acsf�)�x���'�d4�1�2d6�(b�f�B�n3���/�Sp�Ŗڦ7j��TVL T��d|����.z��8�c�u���ќ��H^�ÃX�Ŗo�H��yCz�qO��cr������n����,��4'����+@A��2ST�B1�k�(і��"�:MǢ�F��pX���lH"�m�v^R�1�Y��@i����3�mY��S)����P��GX2M����ҠJ���Z�4$r�v�8��ZM���h�k%ݪ��tLy���E�y�v�͹B�B&�L%��v˱+7*@��)���Ĺ WbŔ�bƈΤ� Oe���HRT�p��f��]i��^��Ѧ��~H�Y�2$Ә	��S�k"a���λ��j�e�h�2�㰖I�)�N��U�t~Wo&AX�k�,�t�x~�]<h���-���C$����
���n�X>���Y2U�Z5��pQoU�Ѷ/h�`f���'"8tB�U���b�ֳ��Z�i[:�3m�Ӧ�C����Tq5 k-4�$Xݭ	P���-i�xV
�n����$����zC��
��R[)���L=x�.��ISi�3g���G3ܩ�m)����c��Gf�+n�r�(O��
�ƨG����fYp��1-�����`R3,H�FH�x�xQ����`-,�b$�< �T0����&.m<����m�o%�ك3$�6:.̫ٙDj
����0�m��z�;QZ;DVh6]��h��o�w­'o����)���J��/���8��mo�*er"������
er������8:�va�(����j�f��#Ձ�j}����X4d��19aW�d�.�c*m�S�ZM�mFԦ�c/S[r�=R
ve��4�
�ٲ�mI��F�w��e j�^7�a���UG�76[#D�#��2�"�E����[�eA�cB-hd!�i��`�O�����"T�5�����f޻&�`)�'���eu���a����ن�j9�7�ܘ饄g*��A0�����H�V<O�6�
n]��'c�����YKV�&��f��@U�{F�-IN\����m�c��,�MVѸ�X���;E݈�A�X��]l*�E��YWlDn�a�,R�JU�ϝ�T7J�H���9��e����Ԉ���e�c����/���2��n�Ӥ��ր�Ime�Q6��<�O0P��jŊ��/H����b��w����Y�(0�õp�J�K2�3,cݡ/J��V��e`.T��������K!7AW�F�r���%��Èjb�,��A��$�b����'4��Gb�c��/)��1�h×�Cwܤ�IrHKB����sP�����ս�+n/�R�o
3@l��b��:qQ÷WL�:ʪ �}Udy�1�x�%k!H졎�8�6�\x��fTZ˪ɣF��ī0�Y33 Ӡؽ����M�G@,���v<�Bf�VX��%I
Q�;:�B�z���a�`���0����p�M�/B)��.�Hf��Z�)��u���&T�4=u���T+2�1�pU���֢*������KX$�coIpa�$u��A������B���:n�*a)��P��ח�wFN5��	+%�$Ɋ+ҫ&��%�x/L�o]�w���:ҵ��[e�`^j}�]&z�l�%W*#j��D`�ѻ2[e�;4�����Ce�x%�i���+MLݤ2�bJ�z��Z�;�h6��ڴ�G��|ͻ�4ڬu�rV̀a�fIM��y*�)�A^e�d!*�7�`���q�s1C���pԛ���S��[ZV-��d�Q���כt"�Nkp!l 	:.��[�rSVq,��XבZb���U�v�Z(1���5��Vk���h:O�ue�V�m�����m�����N�7A;A�mT�e �B�����VE��Gi������T(�v&�u��mPYa�Y�ڻT�n��Z�[��w��m#�+yS	�,Dm�U+D�q6��&�ԲH��w�'+�m*��IƊ���w�[W��wO  �HM@a���K:�t(vuBDY2[?ځ�{GP�:WI��,�"�
b{u�f����!�X�24��o0�gc
'�*u� rP�r*k=a8n�b���Q4Pl����Z&�(���������rF��p]YA@de^1�@	cPP���3�N��h���hD�D3�;�L�C���`Df�i`�.�U�8	h�ܝ*͠E��)'I�� U�C��d0
�`�	�ؽ�ؼ[�@�h굛Z�}�20�R��d<CS�`ƀ*^f�x$�"�[mщu[6Š���h�"��"^DH�r�0�f�D4Z�
����^��1����q-C�=<@Ւ�G����3��<E�|.�����H�m"���z��7=�x�p�!��i[��hO�	��A ��V׸_t��h��Ȁ�g�yБH���Ah(���ΐ��*���̇��M�GP�R���t��$7KHYʲ�$�h���*��Ն�Թƴ�9:�V�%��!�@�P��f�l���rl��t��cH�0�K�Y�$�Й捒t�*��QV���l��e3��fiV($.D�k$�i���v�鏕X��o�A``n��� h-	��0\���ITV �{k�pH�ӠeYc �qQ��WZ7DY�x�j�QL�d��g��@�m#i�AQlZ��Y,�]���.^��1�����;���� �_�O�G�{�	�7���_U�w���v���8��u&�[r[���m|� N^�ı�����yO+���CU�MWI�i�wZ��WS/n�{��]8���R-��9ʲ;΀ޙj�+���C2F�.���mqNМ���j�͍EĐ͹�^��S�6�]8���F���p؝	�-�+;ic��]���:��Z�M��e�#��b�{9����2"����f�m���Z���xE�{RՎ��ޙJ�8WoZ���=�S1}��ݼM��qs�&�1��L�U�
/*�\B�:x�[\�/�N���9�5��Ք�^tђ^B��[p��;<���dչ��
�t1m�)�97�tM�6l��h���lb�>x��=)8!�&�i�!$�,�90s�in, ���-�{��w�[����NQb��:{�h�Z�ֶ;���hxa���}�����&�W�;R۵y�l
XIahwU"/:��k���nY�a�L�s��X���]���m�ZSQbn�M
��no1��\o+��Czb��u�w�Q�o,c�L\�z���B���
�z��d5�  �yPe��*g��W�E���z��xѲ�n�=q�,����(h����Kvne����h����e����x����pwO�Uxض8�J�8�E��ef�~�:��Z�S���"�.�u��k4����CTm㥮1���O[,���9�+y��,o]+q�%X�C�=�Q]�ǻ�M��Vj#ݓ.��2�9!�����H�&�.�q̙7�<hV���;�WN�tՆ�h�����Lyr �T�Ì�n��j6n����ǹ���q���ӵwӈ4&�#��@M]7Դc��5YtX����3������K���I�˝���x��}��O)ⶒ�=�ve)Eu:Cd�)u�vFh�3:�v$@7��K6�{�a�>��솢���b��� ��0����wh6�J]�e�F���77]��Y��Pt��v������&�����,���ƮDᝢ��r��Q_�c;9����
�;�;þ�D�+�Pb�Y���ذ�;��V��I��#+i��}G����E�;w3p\{z2�*�r3e��8�&��d��&�;Y�;8�;�#�9F�ڊ�-��2�q�NgW0+��@��ͩu6����V��.�C��ԏn�׹��l6'+�A�Џ� �Ժ�f륱>����.�`�R�
εՊfb}�DS�T�˨����,����zoќ�ÌF�Y�S3ˢ�9+��+/��)gr�.��=G����R�f7E�mX�D0y�6m�2C6YO\d��u._.gY��R�三�A�ٝc�TZt<�A'��=Rʳ]Q�l�;���⅑��P�l\�c	f s����); �Y.���*M���j;7D����:-��'"!���3�^7��d[)I��ζ�u��R�$WWW�3��F���z��s�� �p����7�5�Gm�%���
�gf��8��Q����d��Y�8��4Gvм�
p�\�;�6�㻁�*��rJ=����N�QἭ�X_�bAJtޱ�9~:��1��n;˹�+�W�7M�qk�.�7c�e�x��a���譕/��
ڰ��I�}1\��y1���r��t�כ8=�XM�Yy�J7@���ݡ�bu�sp�{���l�6zw9ɴ�r�nL)�䩛�U)_M����*I�2�훖�A��a+kT���ݥSs�)�$����}�(���K�'r�:]A�9Iʼ�gR��渊xr�cb�	��⤀Yc�՝�2�܆�(i��"E�s*9Jt�_�ۍ���w��¸ݤ؅�����cv�S��1�J�����p�v�.���mLqN>���G/m�r��.����J4�w�^tUo^,v����1�S�~�����q*!��o1,�u�4m�{������`Q)B���BZ�0d|^W9{��ꏺ(2oXwCP[���=�/y��CT����ߌ�N��m�<��eK�]�bn:���ޙ
���R[UI�����^vo9x�V����;zEЖ�#71a����ޓ`���O]�]�k��4!0X̨�'kC��];��%�.��0ͧ�^J��M�������1*�֛\���Scf�-sq�T��:�Fe ��0ڻ�K���Ů��1�دWH%cG�d㽩O�M�AN��gE\��+2��(M���xwm̩��KIF�ԍ��r�
�v4+�`*�P>�浪i�9�:;���f�7__��W�ɺ.|n�']�����c�D��t}����7c�L�≸V��36 �!N�޽�����~�4�=���a���V���b35f�u^��F�üڠE#���.�-;�W!��!�Msd�)�5��jmp:�Ć+y���m҉�u������I�;��AXjŽǗ'n�u�e�{��"�znP{V����}�&F���F�Jc:u7��u��a�Wd�)D5N] �]X��z�or��Bț�Ã/z�[iLO(匛Z�����Y��y��s�y.�#"Q`h��{	�Horr�4���t���kEY��[�-u_��,�볔O�{!N/4�Qٻ�7�2mS�8�F��;u�`7���.�@�Sm1�oo�TZ��S׏.ݑ*5�F֋�!Y�ٵ�.��hwgU�8*����m� jp4���ھ��f���|�o������M�O!��msV�.ڰ(��8�z�l���кP��롙�w�\�Ш�Ɣse��H�bG�uQݨJ�A��݄ۧ�X��n����y%r���+�;1_]_b%�V�cz%}`���yqu2Fe���$��3�:r���_e�ƫH��r�}��7�]Ǳ_edM���v�);����͖�dr�=mG�;���D%7 �M��c�oX��뎐�F�汇����X/����!܆4�h� �;�f���R0��6s��N[���wu��+
��k��J��%��{���Sr�ԇ7\�%b��'� �1�v��y�w��G[�y;}y�ةH_����t�Sх�7����դ��[�:-��jTR�65=��.��ְ��h �NQ�ٛ�����*nmQF�+�£[�P�Y�^e)f]����A^�����e�ˊgu��^�O��yxּ]{b��*ݭ8��%�% �q:���8���\$�>z����)��C=r|�*D*��W��SiM��w*����b��s���Vu��5ǯ�M4Ca�ILuy��뭸ΛTQ��}K;6���i��/�,wݕ:�A��{�M���231��6()�L���Un�e��pk����s�ٖf[�+���i��o�Ι����.�Ӵ�Zn�Ҙv
U:��P�����N�ʇ,X�e/�y���}ʂ��r4��X�[�بQ<�}��#y�Ueӭ��	�8��butq*��[2eD�)iz_D��
�m����I4Y�4�{tjęa^���E�'� 
��2�Zr��h�2�a%�V4�+	JK���w�ѝu��G��ʰ:7]Qݛe�]s����W^��8Ix���V�Y�J!����	����*Zq�2r��rV�E���!��|�/;���\܆D��}}e�]���DPA����wBl����]�r����۷v`��K��Ikm	N질AYr\�YmX���Oq���k�{v���R����x]�x�e�&P׳���@jtT�;b�T���w�_bf��E%c�n�Z�V�|� PZ��&#G:��7v�����v���OC�V0�*f������͚��j�Џha�+i�Z�����-�핸�5�r��7�r�).���")ܵ;9�g�����*Wgsq�8�욑_n��Zcɵ�KIv�p����*��쳱e�ɐLSr^Fp]Kn}�$ݾV���).�f"�I	}��>t�6S�9\�L:����6�`Ѥ+ڷ�^-m���:������@+咝��&Jw�u��29oRb�������.��^.=XVB�Q�T#��Z���;m��u4@W�It�܍me.r�bq�'9Yw��!3���K˽ލ��u~��`��/�8}Օ�u9L ���N��1]�w�5ws40�a���W@�=�����N��f�����Vx�Ia�G �:5��=�ex�{{זCaK��W���fJbj΁�O�2�l��"��<��ݣ!��"	�p���M���]�t�����Ҩ:�x�^�J�0�{5�ei��3���ˆ!�.��P�6$�1G(ۮ��j������%n�}#{x�B�����;��tTT��4IX����bΛ��l|
���#��/%��AR�f���n%�m�ش���e@�@�o'�]�%+�%�C�K#��Cm�i�w��6����w)�]r�A��R	��;w+`�]ʥu�w��n�VYZTY��������#F��)��ǲoCf8ͼ{�)B��gu_P)�{���ox��m�n��X��Zc6�gV=7vPoy˭�t�Y���q���P�
�(��:3�Z�gkW�&|b��k(3v�h�C�M��=Ǖ2V���J�d2�|���(S}/Y��6[���fV��fc�ܬ�\�	�V��B�o6���hasJ�m���*zq@F��9��t�ڽ��y_]��\�Ef��o{���R��&ج�cSv��j�H��W�@� 蜘��=XTp��g+l*{I.���wDhz�Y�[:uضhef$h.J�D���L?`���"�k��/S�������MVy��uس�ԕeY�v��R�Br���J�i�
�<�(�3]�L�w��@��������+���t��Ĺ�Tt�w5�}db�3�/R���u*v�v>�*�qۗ�Lӻ��I�Z[�'�4�6��G��׳SBuΝn�WD�/;V�����5nS22�豰�[]t��;�{� ��H`΀@�^-��ood\ˑ��Mf��k�7W.g �$�BfYR��}�)z
�s Ʈk-H�̠�>�X,�'J��*���f^شծ� �
��ur��ٙ�`
Q�Ɖ[ �G$6u˥�π�\�-�'���L��ʋo(n�ASn�̵,9����rY�T2�7n�����*Y�-������>am�*R�WzL���p��\����4�����ol��Z�=\�㯍���w8�����:�t)49�r�*r ��#����5�]X�<����Q��]�t���g<�����j��m��T�����������FN��)m(q�fp�*���kǍ�B��B����C�	LZ�:�&���iT�_^Bf���Q��a���o���9�fё�ﬠ-S�ɢ��N�B���#��ve.WXt�m��\���cIӭRr=e���t��s��W�$�s�X�G�u��F]��অ
G�Y����\2�D��"5ɛKv��+uA�䕝J��_S㸺�����;w�|�
]2j4J�TV��o���[ܰ2��d�+�����ΰ�͛-K36�s�J+
��4CO7n�H;txS��H�������+��[��3��Nq���%U���M���;��i��u�x�j�=�{�PDˡ�v��<\��c�$��X$�o�rسy;!ʤ�a�2�0�(U��ַ��>��,��=��w$��2�jm�o�?M[^w�3�!��jȣ���P��Y"v�7�"oRM�Rv*�"�\���R�jCqIǕ��������{��[m�v��:����L3�����׫�w)k�Ċt��y}z�J�	{O��/���m�;����^���Z���V���./6�:>ʼq�n��T�
��뵢Y쫵թ�u� �f�AKt��v��f���h��-�ԃ�RM;�4T�N�$�9ԺK�^��3mu3������T��k��V.9��J�,��ѵV�7�T������y�V���*��;�1��{�c�Ê��S��G�@�k`�V�s����մQ#>7�z�5W��x:�B��ڤn�)t� 8i��w&�M-hA/T�o�Ls�bW�x9)
f�C�u-f�ѽ`,]�Q���	F���(\W�iv|½�p��#�-
�m[�b#�Q�ˎ�k\z�f����y�%Mo/�EZ~�-��FtF��7(�~�fhV7�nb9}i:�/`�,�c��5DWM�6���x������~�b��j˶�<�����3�n(����n�����CW^6I��ΒI#II$�I$�I$�I%}M�����;��!�`�����<����n�����.�g�j;s�t �}�%NEmw�!����`(}���6U=��>w��ߘu- y?}��O /pv����ɤ:��P�%6D�OL���䜞�{��_0��D���+�]�����E��.fu��? ^�e�b)I������?<� �rM�}��!Q����_��Q>�9��?W�?���8G�Q���?��?����q�?g쾚�D�~7z_+T8��*5��6-��S�
[B`��
QU´��ܣ%��˗l1a�5�dTr,�PS��y�NF���u�řV%i��*n�xs�ُZ*�C"���������\k�+j6n������UdΖ�f@�R�R6���&*�z�W3҅�"?d�P_t�ye;��y�Y/�����N/��;�j�Ǘvs%����ef+��CTP��V�_C��_2������d���GyP�ӻa9U+�������|�*�����Ԓu�!���l�`�(*�Z��m=�0�_p�\����nl5�*:\mnɁ*�J�kynۥ��Y�%��/�L���
ۥԵv��,�}Ժ�N�b�h�q�Q$(P�Mҩ�\=[�]��](���mZ5R����[�)Bgm]���T�{Nܾy�f-ú�Z�*�dj��;d��];z\{�s+N��-.,�|vD,�����gs�w��ZN������t��S@%��:����h��v9A_'�]������h�.��]X+[
��GRQӅR��Q��6^�pu�O��]׽5&)2���s�%	a3�:ɴ��!�ý�K�1+�m���#z�/*���d� ˵ݜ�8����WO7\|c���a��XRg�@��i�
��q�G�o�_]~?|~�x��ǏǏx��Ǐ�<x���ǃ�^<x���~>>>><x����<x��Ǐ<~�g�<x��Ǐ׌��Ǐ<x�x�Ǐ<x���Ǐx���^<x���ǃǏ<x���ǎ�x��<x�����Ǐzg����<x���<x��Ǐ�8������}>�/�����}>�O�:Z5�Q�S�n�gP<%m6�hu���N&�:�![L�y\ΤE��!�0���e�Fm�Y|��ךT9���A3����yRPL[��X��g{SV�7�:�/�u�p�n��[pei龱���q�0�B4���m\42�d��'�k�F^-ƛ���ϮS�1�	.�� KME)�ݭ������.f��Vy�{ST�B�U���x��}�ᐴF�{W+UW��򛊉&��nv�k��#�1d����0����a��r�pX9�8�y|t�p+a8�t2�a���T�dK.�%Ip+u�0r��0�b��d������ ��w�K7�q���7��T�V�#�u���(!��
�(�Fn��M5ͫn�`%޽�J^���jG4
�dRD�P���h�jͭ� �{p�n�ܫ3���E(*lۮc`�F�,��I����)sUO1Z�5���$�@���`�l�xyj��3s]NA���Ƣ��>�ŊZkx,�xQW��K2YS���$��� Z�n���;R[+{���j7O=���9�v���}f,"-�V������9v\eP	��7+
�VР���:Z\���m..śk�^E��>�f_�/6�7'0��=���B�ڕ�g9����ݟ�o�����qo�3��ǧ������Ǐ<x����Ǐ<x���<x��Ǐ���������Ǐ�3Ǐ<x�����x��Ǐ<~�x�<x��Ǐ׃Ǐ<x��Ǐ�<x���Ǐ�<g�<x��Ǐ�Ǐ<{x��ǧ��ǎ�=3��Ǐ<x�x<x��Ǐ<x��<x��Ǐ?^<g�<{y�s8|�0���`�i�@�d2eC�j�3o��v��E��wG�-��/^4����
N\}Ǉ4s*��!��L9s�˻x�t�U\[�����z��H9�+hd�*��7R�]Z�%n_��7�T�����c��%�׉b�e�0Q�wDB���+P��5{�en.��﷦��śu���#�� J�ד��X�32XD�f\��ʕܞR�[���x�$ђ�ݦ�>��QU�Йg� J�8dF#��tܕ�J%[;���AA-�q-�=�Nb��ދ�+�jRcQ����[�T�s�dԤ��ތ��t�@R�\Ӽ�3|7��~$0F�8���u�[]$m��7��Z�������b����`P��O�=��6�趃��5L�rqY��m��u��k�-�GE����o�9�X+Mc�,�{�N�ٽ��0�=l���;�.ӯ�A��5+�� "`�r�>��*W@qn�v��cr�����g��#h;�)��+�l�N�mp���q��4��m��}��]J����fd�Զo�Z6 ;�`#ohi�%�,襜���2N�U��8�Wue��/7bO�ט�ӌ�TB�Gi+��7κ��M��{����s������Ǐ<{x���^<x���Ǐ�Ǐ<~>>>>>><{x��ǧ�<x���Ǐ�<x��Ƿ�<zx��ǏO<x���Ǐx��Ǐ<g�<x�����<x�׏<x�����Ǐ<x�x�Ǐ8��ǧ����<x���Ǐ<zx��Ǐo<|x����>�O����}>�g����l��۪�uo�0E�WP\,t	���U����Y��RL��鼮-I�|���Y��)�E�e� k�hJbo�.�u�����b�L;6��Ӈe�Awʭ��p�`�9��81���Neni
Ҧ�n]�&�Y�i��MhR��Y7��b��;_V=��`�"����d�֫��j3;���ݫ���uS>�W�q&JX
��ɱ,�m�c��t'��nu���6�I�����Ԡ�e�[���[]�ƍ��3�)�8�^UL.��m93��śy�f:Χ�����
�:�B���
w�$��g�U7y-\u�4��MY�k�3V�( �/u�U����F��ۣ�k:�ؼ��e��8�I���o��'^�5u���C����ޭ�=e��ڱ��Jv��1Ռ���8&�y	R�n��I�5�XT����sg�cs��.nQ.�9���]�����m�_�9�6.�cP���ҐWȁ�9W
˻y;gs�y[������+�l�|����HY<xb�|gl���l��N��
8f`���%�SV$��]�I�WD�WW�2�ty���=���3}�H4 ��_rT�\��X;���I���o��hB�}T���l�%fzQ�r^$���lZP �Wu�ծ����s�x�TܬX�jR�\������R��{&�����bT��]/ \�{�vA�(��q�w�~@�'�ŶMW��ZN�d�y��is����5�W���,�K�q輔����Z36�T�6,�U����&�����%K���u!̒�[ܭ�/~�A����U9h	�D�5�\�p[v�hBFܬo���A�E���]'R�5T(��s"�7F����<���V�tἲ��M
���'p��WZ�f�5%�{��z���N}ͥ�ԕ�8�_u�7��$'gSb�Ƌ���ky��T2�����ۊ[j|��.\:�R�b��d�UWÕ"�7�J�ɣ\i�8D�yF���?��^w;�wZ�$�;w�h�"�ήlW�д�Y_ۖ�ķ�-�4�G3$�uv���d�5��N`�$��KZ�v��=�,����OܶM˭��Ϗ[�i�Q��־v��Q�RX�_q�B�*���W��h}�;�M�fp��֕v�uwI�(]�<~��S���iK��Dm�ōx�̳��/��#�d�X���+mZzN=�(�=��L+�l<x����!{Z���9R�4H����u�� Ó�͚����*�]�(�
��"��+��3�zB��Cr�ZKz^v�N��z�S���Fjƅ�]9U�
������/}\i��)jY���ıxB��7f[��[�#��ú�*�� n��1	d���>���#_U���$Vm�߯��X�-�u��`l�Cڨ��WM�ݿ���+md]"��˺���.��)��^*{YsU7;wr�'��$�}O��C�q��}�i�ˎ�H�h
����k91pwCXJL}+(V�����Kx�������N,�Q��X�/h�sr�+��k��ƺ�����r�!����S.�����>q�7i�N����Vwz�Z*ƚ�93I��-\سCSiWĻ�d�Z{kU�lna�5�ZVM�}lE��:����c:e0��4~��e�S#��p��#Ō�C���c"V#��9��TT���k��%Wo^������S��j�	��7>ue�wV��J�!�=����t��'��Iʥb�ŧn�yXcK��;Ϋf."��
�w-f5� �Б���X�%��2�6��й6���Q$m��K*�7����E�)>��5�S��s�s.�H�!2�
�V�K���b(ٹX�4>yS+��\#�T���:��)6�h,�e��3']�s�jœ�l����Um*JP�}_l�k��޼�m����l��1���vt��._:|s;CFk�b��*��nn����+���9Rl�}wB��̕eR�o�,/&
,sB�*e��yBR3�<33Nf�_)#X���E��a�V�Z5����z�+��_en4���X�n���{Wo�^ͤ^���8w�H�;/R�Fښ�؋	<��-�
�66�j�PE��qֽ��m��H�P�{�VB�@�md�Vf�]%�dk�(vDE\�Lu����O�T��]/j���w��Ƨk��1��'.��I	c�7⳺���E���3��7���i�ɒ��"��T`�e�ۼ=�	z�vΗW֯�r}�-=0{Ӷʬ-��J�2�Wq�;>��U�̐]�NdTA���4�P�U#$��|�sI�Q(Q��c.�&��*���iUm��)��<�b����2n�����b�+�.��t�g�\w�����Ü�ūuk��Mد���V���Y�l�qv�"J-���q��Jo�"%e�-�@S'_1R"e����ю4�:�s@�t�f7��C
�����B��k�ӗ,��V��6��^�`��'o��B,Ѵh.cb��d��7�7�҅U}*d�K��)p��klF�f.�M��p<�`p)�����A��9��m�meK��N��X��V��]��}5�	ur�0i��Cdb���܂Q��Fەuo�����n�����߾��
���j`Ql�qd�.iW�9��߬*��7����bG�X�1�#0-�V�de�
�p�ykF}��Y��2�׃��]!G��=���\��y4���z��A쨣룕�]>�V�ooF�76}5÷����r�w��b����;U.p�F�pbA�Z�4~�Y���M�����+�q�#�O���m�ኦ&�ݖD6��uN:Nݩ�F����/xq0)��C�b�����@t�e[M�Fu��{ǲ��ƹ�|��q㩵Cۨ���˽�t�up���5��=��蚕N��I|gtj�Yg.)mV�π�i��-h!0w��@�y��5hT�bQ�`W.�R֭���ޤ��΍D��Zr�Ѷ�]\��K]>Kv�]ꭇJ��t���6�]���y��Y6��ۘɳ��)N�pv�����\8#�O�
��0 "&�U�\%�w6l·VJ�wZ�Pݔ���Tv�o�l!���Jm�|�-ِح�X.��5��3a̴{svȬ�H�RewJx��Y����/ ��!g�3]��ŭv���GH���.�Hd�g�V<R׶kv6��,����	z��_^��Za��V�f�cM�ZW���=�u��M-�$�,G�*"��N'���&a�n��0`;�R�ȧ@]l�ձS��ݙ�h�ݷ{�786+,��u�Z���Y��E\��/�"�W�Lh4j��T��u�R�8�i�(Qt�����Sj栬z,�6h-k5�[��L�F��h����T.�.W���Re�!���`�/u��"���6��K�+���Vݸm�9u`�T|�9�<��t*�jA���Q����:}}99Ƕ>7�[ߪ�Aj���F�j�˚1���.�h<��^��nREb�=*��t�p�{ ͦ�e��;&�:����@4�j�"q^���n�X����f]vf��|r��wr��({\̴���/s��Gd���oR"�F��ZUW�F���2��Z�I;m�tMW�Y,R���b�D�!�n��x��R��C�2�˘p�[��n;�um�敪@���z�+:����ʖ�N�;���w|���B��ir�q췑2x���|���S��7�/�-�T������ܫ4#jnj�f#��*1B�8e�]XU�DM�E���Ǜgj�o6-SX�d������s�迵�n��;ᶋ�T;"���\?h�.���{0���`8�tG��2˧R3\J��z�Ig:��K&��i�kztJ=�c�ekF�]J�S�NJ����)�:�9|EIv35e�:+�osmI3��/�e��ot��[7�d��VK�Gj��%k�K�Fư6��ztᣝM`��QM[&�i��j���S�es2a���|�"Sd��O_<�����Zݵ'u)]NL����Z��oM��w�;z_\��*�Tzu�P�.o{1Hst����{L�D�i��#�n����s\�\6�[��l�L)Ή빹�v�����s�$E��x��C��Pؖ��j=�Dj���\��.����}ʹ,���xtq���ڄ�[�� ���Eh.Гf�̭k����uBova���P�pÓN^qs4[+��f�%jEQ���]��W�+��y��0��r��7Z�כʘ�%��N�Y1�Һ*�3]��q��r��Iͬ{�kp�u6����K�{*
˔F�}��J�W��U�GB�|E)���#V���We>�;3�D�r�A�[6B�'$�S��I#x�Z�1=܃t�MeoT�u�hA]�(�,�1E2���I�,���~jf�T�^��;���˗f����*���`yp���K���A�w{B]��)
��ۊL��J��@E+S��OA�T�\�� ܙ|=���G+<�ǐ���kJ��˗�\|8s�n�=w�a��v#��Bv����}_��J���ܺ�W�#W��q�)v�.���������3Ll�k�3.r�N�}�'Jt��疔;�y����__LvWK�rդ�Kw%l��jF���TK����8�ԣ����Ώn�6�(��Gn�{G�n��3�U�'��m�y�Iقf�9�,>�\�B�t��!uQ�� ���Qǜ���W��5\�Câ��Wv���?����7� ����J{�����w���W���O����u�;�?���i�a�/�"m�B���i��,�J@�(HZJ�l��,���D`%8����N ����m�i9�M¡���"�P�HjCe�E|���h��)$�m��D�(��.@QlD$H��(�dHH�m��H�p�����?(�E�# �>f7a�؄�	�M�t(��E@�Dڄ�e�g̈P�BI�J��/��J�����D�чwV���o��q��Fe�ߛ$rK}�ӝ�+�m�G����GcUIҸ�-��!��wai�;}�w�֋�<v:�s{���u;�J�9��9"n5�T��]�$�� �1��I�Kϻ���8u"WK4(�T���+YCn�v>�5 c.�����x��Ҡ��������������h�Z�WCqTJ�M��lF�����rac��#�jf+̵�z�Yt�mhC���R�e�B0��Yo'J�E�)FҎ�m1hF���v�����w ��X\N���ӳ3r��S ]�9wN�p�b6$wV������]��|��ӒK|$	mui]��f\	݌+���S]�����۴�i������R�\^�}P��ȹ�����˒i�O��T�f"

�V�V�S��B[ұ���3O��ӽO4��b�}*�ޮJh\Uc���} �/dY[q�Kˑ����1�*����N�LK���}�-u�y}cC�g�����x�IJ��K�W��ω&��]�[æ��B�.��%�N]�ea���o�a`���kʵm��0Pe�8]=�ׯa`�B��T�9�[����̲O,P ����Q�8'xM	 h� 	"!&g" .$�_(��"Ēɩ�
6�?D�%�Q���(B���i�BL(S���G�AL��9T�8E���c$R�F��B��� �9�O��"Z �)��*5Q��m��M&�B/�l2`N	!"�	�P��&JH����%� NRFH��̈6Q6%E6I
�	�)
�SL$���lF�!�ډ! I(�%F�("b �p�"!&�QHĈ�q�Q�5�`�\PEL�"�ԍ��M�)Pb@R*F�,��8�0�Tm��i'ɩ��"��N/�Ѡ
� ۆ!>�$�R6�L�[��A ��EI�$���"ܑG3��3�m�޾�"�2��p"�0�$���`ildQ��ff�e��U���Ƿ����������<x�w4�"f1���FJ�l[�dlV����n�f��OOޞ����<x�<x�'	3-������0727�L.��r(�sBcswcM����,3^<z{{{{{x�����\}}=��*�gjzzǫ����,̺ުè��]���w��;���h�fe	�]j��oX�tu��환f����]H�Da�Y[��ʑ�uuuD�f�%P�Y�#���U$H�gP�Ru�u�R�V���d��ud�ZA��.����e�f8�n�HfZ��ֻ�!��c��7P��η
	*0�� ��AD�E�����l�q����IA|�e �Ҋ�.�,2�/��������M�EZ!!E(���
.&�2�$��) ��������%D��_%D�XH��(�R!�I�D��:�-é޳:��gI�#(�2*���ڳ^�س(�+��#~f�m��gY�ldT�Vw��DN�L�Y�1�ae��5�Y���DfeFfs4��;��*(��黺���_��t/�I�������RJh�d����&�L��Ȟ��5����I3�Q\o�(Ȗ�1q�څ_XOM�����+c�v�{�wX�����n���?&Li�����4�)���e��$�,�d�i��q�b.(�b�p�aO�	')P�ݚ����z���3M>���b�@�Y �
I&I�M���W���߫�v{�Rm�}:��C�>^�Nq&og���6�;���t�{|�E��]R�;U���L���UP^��k$�}~��|x�CH�Ƿ+�Qed��Lp��2k�yH��s`ͯ^;�W;�-*�����ߞoޕ�bϼ���'��Z�R�\���=�ޟ?u���^�u\�;"�8�f�;A�t�`�|�2:1�׽��E	iz{��w������eQ��z��}*��b��;5z��Gg�e��֪�G�=�9�W7��~�H:tw��O�L-�>�4�]�u����щH������0����)�?o�y�a�[�f�+�_�/��=�o��zj�O���G�	�`"�P��FE_uP��#�χӖ�4��5;%�СK����>�˨T_r��l�W����3��vhG�?;�����;�$t��0JU�ؚO+o���i�gt=R�;F�
ǔ�jsQ����]enIw����36U���L�8�{��9��e�Z������U�.�z�y=�Vc�R��c5��ū]g��� F\���YZ,��u�b��ǩz�ܩ��|��6�2�>�}�q�S��;1���Tf=�:�ݴ!T�U���+���½9����=jE��Iv����C���^���@g\ڳT����Ͻ�Q�s���:C����f.���9�Oީr@�rʦ$�r��T�˃��U}���[���{;�߸y�0{��9Ӷ�x��)s�3�~~��'������#����KA{0	����u�P���Z�Iʼ:�L��\)����I��<�����m��]����e�y[ˆ]7uk����sb����8�[�_uW����1�������>�c�n����\�1g�֥v����^��y����uv��i��S���勽#��_�mg-�֦�'��3����4}����Wm�'(�%Y�Oks����y[�YER��k+Ǭ=�@0���*�+5�B4���Ч��kX��l]`�W[s&ɷ�>�Е��Ҥ���F�z�Xv���A��uDR+��b����^��o.�e����p�w�wF2���7-5$�̒t���XA�a���8ƝH��!��%�̰�nU�荒�tT�o�K4��Xz�h�u�{Ct���I�f�̼�k��Է`7n�{�-W,Mħ����g_�Ϥ��ߟ��"^'눨^���������,P�giCUt���S�gE!�����om�~�a��{��XJ��:;f\�'@`@�]�%��	5��g�����fɱnO}�ٮ$�,���^�7>�W�>�r�����G�X_;GU6��jc�#��>u�-�=<��|Ѕu|�Й��|��\-;��~|
�� `��OX1�^�Z�Ww�ySq9k�}>�rUdA��ڝ{�/���}횧ƣ�g��53_��1S�c�]t�մ�R�_u)�К�kqM����t����<�Q���b5@�����M��j�ܾ�{�����ؠ��#|pM>�h�k��k�d�_mo�g!��EF���߷Ȣ)zZ�???f����x����ֳ�Z��v(Z{y���གྷ��/l�A���b�;�F�c�^Q
��xn6|4M��Қ5Nd�T�*��8pi���m��,�ñ����ȇ�ճ1��]�	b�ڊ�U���?O�m?u�u�l3}/:����,�a�A��������ם^��ɂI��NLٷx�c��.j�we?{۷��܀dWpP���o�:=Q��j��;@Y��;^ٻ�9l
�~�T���Ds���J���3�2��J��}�����>�o+n��`�:;�=[|'>��$MW�Z5V��EC��:R��j��A�:��o����&򰆫f�%�Q��r��o�/��bSk��w5�����	�"�gv�X�d�dޱ��#���׀�6���;"��gm�HomW�,���f�����OI�w�3ޭY������yD'���E�@P�5s��p����ߙ����(��!o���yC^w�'�ڢ�����T�h�Wo�n9.����u{k2Z���]�{@��췼�k<*��\���`N^(�b�{��:pO����9���f��u|W��W��62fE�{S��u�6�5�I_K�_SMn�ͬޛ;"i]Y��.f�o`�����/3[����.�b����y�B�xqܛ�G:�G�)���[UU���� q7*���.���9����LHFd1�!HF
��!�Ao�bz_ǚ�RצD|��Q��MW	U�]�Y���e���s}�!�o;a�2���f��}}T�����3A��e'��9~�u�'	�~��&R����0�O*G���j�½�����RK�'Җ�R�������m{(j����1�p��['���#�=��*�z�T�{>^�^�g^X��v]����ReN�����bȹ���8��uV�&ex*��'���f���4���}'_x$l�	���\�~7��]�D���nS^ϯ�>\���0�eA�Z��<��{�n.�^Gﻲ�Q�&^�󖩭��R{���t����M#�MQJ�!$_�Cnb�U=��=��v}�g9~�>�}�<�ͧ��'3��'�zw�)��)'1{}9�����2>�xO�^�����i,[��8{�R�hke��渖�F]�vQ"UÏf;��,�ܣ;��H̬�Y1���q�Z�`QgY)h�K)�J��� C�:@2�#�i�9��	�5#w�N�9Ł�#9H��kq�*X�N��\������M����;}�����wU𢷍�>�u�y]���G:�g��/7���}s>���Bǭ�h?{V��bn��]Og~�C���矷�O>k��w����{����?@�����^���ji�R��zf���NC��������T-h���!c��9 ��w˫��*�g�gĿ �s�K�ϫ�����oQ� �-�9����#�w�'ɪa!�4�����As�,�+�G��h��=Ċ3\[��(�?9�?���W�E^��mz�;y�H;s��BյҤL��A��;��w>��'�����reͫ5^f׶�R�T/���n���#�����&��z*�lZ�]���'s�����*��t��?3i��Jn��>�z]�]xoI]m����î��&���T;���D�~�u3���m����j��8n"�����x���Sޥ�bX�񫙮������yL\i9���qf���� �\.�>Y����L�o�u��9��Թ�t�Wap�@Z��[�bŧ�;D�/[��
t�s3kW(�vE�1=}J�q�w�J�\j�:�(Me�yF���U��.��8��o����6���LD��5Mi�>s��3ʵZJc�彀��z�����9���`�����٩&���^���&�7�;z;[��y�9��mw���0*�~j�������7�]�
4�{������p5���ל���r@��z{��k������B忺����')��{�ml�����s��"�z�h����ٿ\�%�N�>~=~N��ru+;v�yB}�Ə)�*�}�Sz<k�*�I�
Oh��f-Ya�EW9�|$������:[S���>p�Ů>�|��7�N�9{<@T���������|/�gr�00c��H���3�4��3��zV���M�UNC�^�7=����>�b����\���Ԏ�iC3�X���}2�;X_(o'�O5�ސ���f;�c�N�Px�B�
�Dc�m=��n:+/l]�6 ��Nd���q�ͯd�Q@\�絙�a�7�y�t��T�����F�~>�֐��.w;�$��Z��p�p9��W^��)���\x���)���}`��Q�9�s�9&�5t덌g-����ډҒX�^f�ƽ�rڍ���yrb}���YP�ʃh5����zK^�A�-�R^��^�WWY�*O*����I
ob�:^IG�)k�֮�9;0f�<@����+^����WB�Q�+w�z���A��o�F�`;gt0z�:D��4��F[ꦨ�z|�)��b���+���8eՒ��T�s�y��i�g�k�
~��gM����X���db݄b�C�u����T�|���fV�)���~�W'��]�ʏ���8���E�c}��Hf�>u뛝�v��S}�=^l��͒8ܝ��~��!.5y��U{=��ޗ��g�V۱�q�'��C��E{q�|����0[���r�?^����m	^y�Jk��z+�>�GSޏ:*
I�� ��z12omQ{���y��Sy�U��Eb�˻�y��}Wukt���FQHR��C�mgo�Po�l���C�ĝ�]R�/��^�s;x�+J��zk9��G(&���l"�݊�K�{�^(L�ɲ�*V�3}r'wJ`ҫ7�w� ������g9��cNe�,��}C��	}��lY�%�DCm���L��T# !�gt�@��>����H!k�>��\[]�0܀	���W��l��;�b���a���'����y�����o����#���5gzF~7�^^m6��`���ٜ���5Lϓ�Kj&=��n��$�mY�;y��mu�`����a&{��^{���O���ss��l��Ɵb�����;�D�7�/��m��O���W�]/mP��O�>T俒�N�oXٵ�<�O)<�V/��Be:^?
U�2��Tk�i��'����&��̢U����fʋq�p��6�{fUA�<Ũ�U��w|�<^�@��E�	�ed��Q��<�^��k�����q�i�zF�a��������$a���y�i�"	w@|��rH�*K	�p~�a��<�=.Ϧ�>�6�dK�x�;$��<���:�j��:�S�b�53�ϳ-��`��p�Y{
7��ӂ��,��f]�� V�)�5�^��.�M�<%���c��k7��m���om0�eUG���1T��wo�{$�h�T󺴾w�����rjZ�N������)f�&��m���$��*��ti���V��ڇ"H*��o-��O��=U�h���ө��-]C.PGl�I:��8�^^fV:�b��MM9 󗺪�6����Y�Sn=�w�kї�Py��wtH�$������M۟e��kΫ�o������h��-c���[3s��ܿ{e1�w��o������M��US��𣾵���U��F���:`d�j�Z蝐��ß׫��=�����Z��D��@�2cZ�P��'�+<�����SkK;�k68'������#X���b�e)�'g���b�����o�9ѫy�|��=�އb��5�9Qo���}��X���i���=�ވ�K���Izy�.�?yd�W�'��c�U��ެ5���̩�d!nY��}鵔����v�FL�����=k՝/����lv�y֟yџ~�9�ϒ6zs��>��*������z�|M)&���Թ��\�ې�'B��N�j����U�޾�ъ�ѝ\�*2	n8Tu����1]�b�m
����,Z��]��ʮ�kjV�7O5)�XE�n��OG��fY���ޮ��M��-кF�p!��4��a�R
����AC8��U7�Ǯ�؋6we;FZJrŦ���Y�])5+����@��v6C�b��*�@�m����p�����@�*P��woI���U�w�
��.n��WR���֍�����M�"{�`j�9R����chR�.�_�Fi���X�U��Xu�I����nK������u�=��4�#W}��>���n�L/_U��g�\��:�s-P	WC������'�Tv_YP�H%�/���V.F�o4�����;Y[֬��!rlc�P��%3u�0I�é��c^3������B��s�i]Bc�&�qU��Vb(es�%��F�)!W����]��u@�ʽ�T]]a�M}���nf�X^�g�u�pV�
]Ύ�U�v],wDԝ�Z�%�1WJ���I�kZܾ�8�,��ak��kx1�o!q�c�55e�1Q�`ݙ/�}[����f���]��S��|~J��*��O���Z�5�
e]��\�#���WA����c!�V-��-L�C�Tf
��U]��(yǘ���C�+�K��;�lB�MEàҧ~����w�@?fc=�v+6���~��J�Q�z#s�S��Uպ����gFG��9r��퇛%��w��.��7!����_!��r���Ly/��%l�|��v�΍G+��Y��wNn����K�M�k9/�Āǣ��Y*3w7d��ƛ�{B��� qXV^ӗw��R��ɡ�z�<G]+"b��
�q>��70t�J��=�5&٭��+65{���[���ӥxΖ:�(p��J4iT!e�߬S�{ ;�����piJ.]X�7Ѷ�#��9����I��6�S��[�+X{�L��MQ�W��i��~��u����r���M���Cw}�PG�X� ������6�ouFzS\ބd��ӫ�ڹɡ2��p�M�p���$�*����؛6�ط����+j:ܫt]�:!X�G�(_]`y�V��Y�4*=��n�Le��	J����`-l@Mn�h����i�q��_Y�2Tn�����\%��5���2�h�@�X��*Ü�$��YY�:v��޳xs��X���(����k)����i�d��R��%�k��/��ت$V��wTn��faK�އ=y�2�����أ������B�1����ٶ*[A�e9&jۡn�G��Lҁ2Ħ��Q��(suu�ϞY�s6��6���3�*��
(��n�"�"�ʫ20�+7M-���6�w6ڣ|{~>>>>>=�^<}Y���{���eVNMQQ�F�w��EF�nc��9&``UTۛ�V:�������������<g�֓��0�
����з�+
���"72��ª��c(�(�,*(��Y�������������xϯ�i����Ys7R(*I˥Km'r�K7�l�#m���#s
�ҷ �ҍ�v374��!�p¢���2��/���]fELQdQT�a�dn��l�Kd�e�9c�DA�1a1Q�	��n㵖n���m�&a�YAF�M0EENYeVe5�Q4m��X�I3l�����s���")�0�7�*���w7�ݢ#p��'�n�YfY�ET�a�E��`N��fUCSY$Q�d��PPYc[��I1�1���,������	E ��$�$
��T`𫳢L�]�� ��^�j���)��Қ*g_���	bN�;���/4(q��0��30}Ng}��}��?'�Ϙ�vO>40׆�>Ly���� ��zg�ũ�Xgo	��z�[K;6��M�U���Ti�vo3��4���r�K>vp�_D3LW�ٱ�dfHv�ӕ�����O�	?��(o���߬�M�_�B��5�8�g=^�:�@Gh������I���r�{��\;Ge�kŝ��J�⥛��ޱ���[�a�%Nw�<�M�Y>�,����d�0�1k�.Q�/�+���n��[>���d��{��	��V�e�>�� �m��0��0k,���GdD_���5�uRY�@4b�}�`B*�ꖾ�~<�E�ۯ.��w�=���{ �����41j�3L���e��쮐/|���4�I+�|�Ĭ��#r2������ʭ~�%ei��шؼ�|�^:޻�����5E' ��"�k�Nc�vS��ٮ��h�{m;��U����pΐ��[��,�+������������6��J-98��/�֪�k M�ˣ�g���ʖ5}�ܽ�f���h�+�G����\��/���	��U-^���@b�^���JG7����38�&�I���o"��<'�%]xCH����F7��x\�%�`9��5wC���%��L��xx��r�x����[�\�(�]�R˂z#m3��pY�����Ŷ�������z9=��Q��剁) �9AX۔&�[�{g�w�-rv7�׋[��'9%p����K�6�tF��F���k+_i�����o�{ ��̼��T��|~?������o��Ԕ#+�a��d�m���Q�$��8@�{`�D��|"�\������P)����t1"�"�j�@zu�'����s p�y�6�,���cH��z^u�nu���]Lu,W�6L�4�ð�>�oK!r)v�o��	�lT�5� ��������z`Q,��-���S�rf��O?������o@Ӯ��1�{<\i��*K�B ����C�%ټͭr����jW�1͜�9����	<�*��F��4_8�ؗ{k�X�r�7��W���LsoQ���ʖ{{x�=o�z���W#��Ld�f���L`��vY�6�������y��]Rߘ3�i}��~�K��~5�Ͳ<�H�����e��Jo��>~�s�7��;<򱕿_�����1l���29��R�rD��m������`�t�7=��-�AWNΌSy�g��;�U+�@L�wʢ�Bʨw���Q�p�GJ�u�:<)��]��x�<��x�w��ho����-&@�K�"<7̀��)���Όݕ�ܷ��D kɏ
B��Ⱦ�a\�s���˞������9�m�%��S�3b�ֈ�l���{�'�-ڷ���7���"�씻��=�����E�ղ��Dݯ�W�bue��$F�Wz�P�X7D��B}���'��"�K���8!��zU�/��{�w2B&㲺+&�-�-�������w���F�pp�$w�ΐp�Cg���h���!�!��aę�Ǿt�I.h$� g�k��
�����}ɍh�P�E�|�Ι�yO��(^�J�P�b��������4;�G�m4E�M�ɢ��7�q�&q"ܳ+�K1`0^�W5�BO�
�.X��l&��B�P���Of�F�Gn5�;�8���
���>�1�p_%�uO��.o�֥�W��Y����24~�_t�� ,ԶO#�[	�[M{�x�?�O�}��O�.]��+�nQ���@�����	=R[��sR�~���R��z69��'f���>h��7oi쾋ງ�aƈ¼5[�O)�^t��2e�ҝ`�(�d��0�b��֯�g�;�f{��KU�t7!��8�-��p�zw<ң~�7kZ!�9��{��V�8c�Ul>y��/V���ZRXO��ζ�!�P�L"+��u�;�������|,�A3�{��̼ͩ��%���P�JOzrml��q�I�#Y�S����^$;ж���΀� �����K��C��F��!���N����녖�#C�ˉ"5Tj<ν�:�߆�+S�}<P6w~��T���}��lΪ��iXV}�z�~Nn��nƟ9���4�g+揞�s����.����y��j)���A}�3�؍,��'�=�vG:�f�φ�h=`g��Pk��Tf���#*�6��%�.u[:�z�vHq4�	ٲZ\�y���-m!�ƊS�y��߂�;��g��k�P�qe����ů�t��[>���CzU�����WM�p��p�@�`0ȈQ��Tv!��*�:7rt 1�x������=�	>��A��K[G��>��)׉��0�(��fvw.��d���Z�r�̄�-�Bj,�X��Y��� ,a�Ô �D���վ��^G)�]J�waQ�BO����.�w�ó�U�ɥ�Y�N�}!�xD&�m�L���Z���e�>��Ɋ�SS�;]�8��>�\���������m�u=ҀU�x���6պ����n�fi]��x2��V��I�ou��V���,3Ĳ.�	zx�;ҧ�K��x�dp嗏:���zs�>^��]�gxg��v�<�U)��2�z��m�j�RQ��U��g�s;P�)7��My��jb3{g&�R��h��9����K��M݅U��^�'�L�>5��	��mO�BOyv�n�=�_��|�h����{�q�^%a���ޣ<�1{bS�X����X��*7�e㩖��.���M7�T��dzXg���r�L79���:u���xЊ⫓�r]i�۵۶�%N�r8o��w)���nU�3�ܛ!�ר������/ @����\�U��L�Q�`t2������$��ӳ��7�H�V���e��
?BN4� ��{}�g_@��g�5wöVRu݋�@��� ���u���N�YNs�9���.���;�r��s!������������� <�
��k��(��:���0;̹��x,ܶ�T�m����Fv��3��oX�q��>F�J8ӯUW�F[�~~~=�LoP%��pƂy�*>|�e�x�P�Y�Q�u�Q�����%5��������Ȓ��@��Ӷ��a)Ɵo�唻��6A�������@u���<X_;x�v�zz9��ڐ�X۬O�9�Q01�F��0=���; �I�����*�Bn٫�}u
��ߚ�K�蚄N����t�ga�[�즱z��@���ٰ�8��28RUWA=�v�{2���-�+�T痶��w�����j��,���d�£�$�e�h@�C��>_N�L�6�O��ck�؛p���e�ӫ����fȗ���J8�3�N�y8���d��=us��.�y�Pm�K��7#��Y�̽�k��{ю�%��@t3�[�q�O��k~8�dB�{V�r�\�I�ۗ������ȱ���x����w�,�2�V�[�%e[n���M�į�@_�Q�CX#�w#^n�ZGn�6k/Ay}t
��u��F�M�N�|v��;}�V�����3q����S�k��X����ɗωC�
ͷ�8�ԆAks�K%�M*���8���K{.��ѣ)^����Du�`��6�K�VaѦ� �������a�˴5(n.��H��,Q��u�p�Z=�ZZ�N���9A�=��,�F%�{����w��u��_-������Lpq�L� G�� $W��|��H?ߘ�X���so��M�s樤��)�T]�%��6�е��O��ӄs��~�<)��\kc>(v�!�j5���(?I����~�P��j���͇�Md^���������<���j/w���V������drV��VF���k�M��:���X_,Ѷ|e.2Dd�z��^��n����ۦD��P/��,t��|dWt�_(-&�f[����Sz��> ���GF6W���n`s�zXcH�s�n�GS�B~4*D��W8�b�z6�<^��(U��B�����\������p.Ϙ����$u,�a�x��|��Ɠ���^�t�Xo��S�<Ʃ^�TXm���Bz���tMsH;l����gW(7d�ڱ��І�)r��o��1K:�>��T�X��輈�#y�
q��x��B��vM<�_P��%m{��\K���S�ff����맚��8潑�3��q�ف�^:����l.��ұC^���E��	��p�,Ls�yw�@;S�"޻��}Y	���d���a�b���m|uot�ٛ��-Z�����ֲ'L�`�˙cs�@�tmC�r��OV�qRފ�3�~�J;ORO��]߲]n9����5֧�ˆ��%��Ӫ��:0��j����r����9G9��{�2R��������	|�����s\dOǜ��33pΰ����o���r�b4,ϊM"�	!��1����� ���d�/�i/��'���ηe�P�oi15@��>2y�,8������{�$9��ݻʪݎ��̅���@�L��1,��Uӳϑ�wU�C3W��\<��ž��d�P
W,j|��oV���nzq�<	M<�3�؏>��xk�^4w�����3��Fm����G�!�̄%{��lz�Y��5?3�/�thw��2�c�b���YB�����Ko�G�����Ǚj%��~��%���2�A�iF'^Ɏc�/ٞ~�L��S������;4J�P^�Ŷs�z�M7�!JE�����A����78՞�)�cf�R�d��9��4�\�y���+R`鳜��wݡX�j��s�[`R� V���a�rvFy�m`3��[FE����C�2ԡ��N�#��1�e��T�����ۓ/�mKp�	ac;�^0�E��|[�w�]����]�f�ɣ��D4�H>�=q��vL+�q{sR����Ԕ�^5Էa�>����J���o�0F�n��T��I�KϢѡv8ɇn�kE�h�L������wg�u�2�zr�R�#@�Ꮓ
��h�Qԇ:ٜ.�2hd��K�Y/U����/u��n�w��GR�(n���6e6��W�>���jf���b}��o<�H�E������h�Tw�7��|�+˗�]�]o�wb�|U�bE��'�������cv1��<�� <��p<<c�v<i/f�6G5T�'�Hޝ��Gr�;[ǳ˨j��J�^7F�	IaY�3Z�97o[�6d1�6�o8�L�4y�iz1�̼��\���e�)��c���v�vʭ��6�:�Qh�6�<�П=�� ���D=��<u���M���Qg��~�E�띓E�C_Dē�l.���c]3���fg]�+�0N�"uu���:�菖�p�Hd[����i��T�@XZ�)Ɛb��灅��!�0�gU)��x��C��l�D9��`0 AJ[y�&�~|��Q�Щ�N��s���-�?pU�(�W�⭙��[B}ɇ�^G/S�Ѭ�e�|�K�m�I���~_y�W��n��[�X@�V@J�}=j���v��`�Z�å�LF�2��ߺz��aݳ<J+��Q�^�C���:=�T���	M`&��bʑV�#�N~O#�_����P��-�\T��|�= ���z��7�ͭ�Sl��,�X�7"���'vo���l}IM7u��^���ͱv1mD�Xn�drR����7�u�r��]�l���N�ޏW]!ʵg��{B��7V�K4e+�t���;�+�^�r�� ����o`���FS�b���.��B���v�n�mw\�D��j_'h��ބ�n+��!�8,���EZ6�NU�04qp7F��|�������|@�C��~{��]{����|�	g���p%T��`�Hְ�T� ���W�z�|������7��moDZᏼ�6ۖ!����y�+���K��Jn⦛iG[����z�۞�1cGl˫��kVi���Z�	̗bЄ�9�fh�,Lo�8n�;�^��~lO�O����]�zG_]���&;�[4�!0�A�[A�<����R�����,�Ԗ����V�{�'r_sǯ9�tL\J�Ǽ�3J��!Ѹ��|�~��z�k?��������R�>�ps=چ��n�X��D����������p{M���	�DƂ�߹�
��m2��r�즧�%��;��,/ҵo춽3� r�Ac���Ӟ&u�qk�cF4�_� k7Mй�R��p�K��,����ji2�s�'C��ȍ��n��Y5��<���s�\48�j�6N�q�������0�+B�0��R�C���eϣ���A�6�{��:c�c���@�.��3�YQ��q\\��\���;]�<1�q�'�t�3�z1��2�,n�hm��-��O��oek|鉡��O=��dy�����Y~�x�9�"������1>��F���F ��Tq  +����7��YR9D���@B�jԞ�ᡗƔx�0ڵN��\�#]���B
�r�L�70[������O��0���x����ۗʜ���_X�;_��i%�s�P���2}�wϛ5ͯR-
<�tu��9�ҭK0携�C�R��I󌰮�^R�I�D�l�C5w�9��2h�u���n�����yoL�	��B����Ifׯ%sM��]�,q��%�T�c�Ǿ��<����r�e�tbV���"��T!�)ى6�1�d�F%��e�D$�L�ۜ�oTd<7[�F���u��e>�EV��q1{���f�]�\R��.��A�>��>k�
��@��+f���%X��Өji	��c��&:cM�j����{��+֖�eۛ��6U��
	�8��5�i>�%�,�_N�v|r� nM��Ԩ�2��+'$��.]1����u�G�}jZ�5��=,�2��;���t�5�ڎs��A�m�7�m>r�"��hu��e�CV���K�1/^��nkgd�+�W��������1Q�dR�z�/�8���Eճ�;a��+lq���1��{hg�}���=��/�d������DK�Q�- ��u?K��/{^��?��C��$�� �x- ��x{��{q�hcU1�.�N�	�n�s:Ԯ��U��q��F}'i�I�xR��X���˲9N�wwIf����f3��WVZXM,N��s�C�0_%s�n�M��8��M�(���[\�}�)jk#���(&�5e:&.*�]e�{N�P�(_�Ms-aT���9I�H^����}���F��I�ZUa� n?Y�᫮W��K�sޠ@gQ�������}���h:w(������R��*͌��>8��c�b�.��ϕ�]6:�5Nd<ҫ�϶oh�����1�Gr���:K��2{EVhۼZ.�l�(�gM5����+_s8��Y�W���t�����_h\L�	�&`Ut�PڑTT�ګ{�n'3^�)b�:+�D�o�h�����7��:SWQ��:��]mww7[vۙmf�]�.I]��*�ʏ��RγH�&���K�*��S���Gi�y���-��3��E��aă��}A�s^�ыP�N�B�.쨶������u-YK-*qb��������(��:l�.�]<N�V��ǔ$_.�l&��)�WN�V��ʑ���a���W`��j#9��a����Okz��|�WK
�.�a�(�6.5�9�:z����oY��	��K�P^���❮>���n}΁�o2N������e���o9gϓ�W��[�������wM�ն��Jۍ]!F�+�$�x������}6��P�d�(�J-:j��y����^�Wj�t��J�Aƃ�ٷ�������ݵ�y�Q˧z
x�mI��WM)	v�'^�lyś�^�㮏���;W�i<W�ĳ�����ri��f�\��
�śZo�g2e���zBF�<m��8;A3˗�6��̼�j�L�l�v{p0�U
)�)s-��u��\��tta�ہ�%��Z)�CW�T���1%a�՜�M�kA�g#a�C�c{�l�A�Y�]�Ѭjn3"��YZ(��N�զ�w���ud�j��5����T��&�;#�-�-��K��Yt�'H
���;ӢfP�v���Y�(.�{����b���^F}�W��F��m�������i�G�Syy/�-{�c	�|�݁��\�'J ��;[���w�����A6���WN���<�6�x�.�ԐiPi�a�a5f]��n�����ĥi�#�ӉW��\z��U�H3T̤�6��]��rKԻ����u,$��*���ze]�<�R���n�9�����v��E^W��y*�%�T��P^���q9bVwU�=8i�,|���>K;�j�q!pT�GuL��s0��-Ó��x�b�
�we�ky�f̮���u��ͰrͩbP�Z��AҦ���)b�$����L�'���wS�x��h��:-ϻ��]�r��.�|�v��Xxr�f��@oa��;���5����6�;��9���u�UDԐTU�Q����cDu�%UN�`t�~���_G����VW�����QUM[FC�LTF�UPQ��>�����____�>��UG����W�ʊ*6Ȩ�2��ĉ�̈72�i�����3��(�*z}|z{~>>>>>����X}}FH�2(�g*����GS�Qu�QMMo��*7scs��E<̢H��0��\�(����2���6���
�7��p*�'")�1�371�*H���k�U�fM�ޚZV{���c]nm��m�UnE����EV`aS��6
J���g�L����eՕQ���DK���e����T�DfdE14�VNU3F��T�dцc�U$��5UC�TT�%4d�5YAE�Nn�MVfDDLU���MA��e�D54E��b���>u��r7���f�!8�(Bfn�	H1�R�P�JV�+m�˫��9ߕ�&��Ktɶ/%O��OfS�fdg��wkf��n��j�ar�Y,�6��ť�! $�
�b7�ad���4�I}
3�C�b0JD�.Eh5 (�H6�M�M��q��51��"Q�������Ȱ0�����-[HONW+�Lu��,�d��"8�p6	��k���Pά{�P��4�8�h�([1��1���:�k��1ԃI���(	fM����|O�;n='��#k�����l���wg�o=��Hs�g�P�7��?2�J�k�Q	Ċ�g�0u�Ƚ��?���uHI��=c�n(��,����|OzD��:>�1�a�Y��P�:��y�d��߲�럷�j���}����q���n�q��Z�W<�;��f��T��[����$;A:�֬G����#�7c�f<�����g�m���z�v���8�0���q��T�=��ۺ�:<�����*����gW��&�����b�B������V?֫�����Xf�=G�(�vQgn�b�Tϝ���d��&>�z����3B��oL#Ô+z�cCpͧ�
�NW*��2�B���y|�`�P��F���^��ޅ�5�9�r��o/HQ�����<����.{���n��w�ןn�2 }��w8�j�C�[�.���v��=7�78�]�B]%צ�\|3���h����:x�&�<9/�{a>���Y�W��n�l�ޓ&����cG6|��u۬W��0:;h���)�T>�n�X�ξ`A���et�5h���y�[�¬�f��4^�ڣ8C�����1敽R�{�VtnR���Y>A���|߇�Q�a�������=��Q�z�G_[�x���kl^�Z����[[/]�#�ŵx>@��N5�~�d��eٽM���(�!�*v^�}RSͱR��o��ls�ڦ��5�Y�mI�u�.{���(��meʈċ+��U�h.��Cȵ)��wT����29��k|\⊷
9��ё\��ގ�r%���s��]��Z�7����M����d󃔧�qFK$�9�;5����Y�QՆ�i�7��ql��O�]D'MS*q���/M
�7����q���_�K�(��h���Oɧ{�8M(`�5�j	�6�x�} ��ޠ+��v(}�=�?M�s�h%��~��[|�}��^�gāeCh��	�����w_z�i�U��A�p����`P~"0��*�?�!f�`�Ns�����}裃��u��Y ��y���1��^F9�^�Ԗ/"!�@f�����=;��]jEl�)�zsZ�[����:c9�Z�����<,丶l]�b���g�5�9;�"��4���¶X�"*8S@d��X�j��(5E��έ6'A����},��3m	�x>3��&�u-�#K�hf��ż��;vA܋9�]$�߅���k�ގQ��yx�c��3ǳ=��HW����ܶ�f�	{��.f��vz��J����J,�R���F�k2�|�iU��P���WA������:,{�a�6���S6⹘l�8/�|>~���aVdh����_?~=sٞV��'?��#��%;�;�����w�X��S�A��i_ib9[Wo�]�C.���<V�^��"'ñ�r��!H���|���3T���QmD:l����.�rsS6u��z�aT��v�V=��1�햠`h �0�8p+�A�<�F�q�i����M9|�����rp���Ō��1~�.%�P���J}x��d��X{G{�������SmA�޶�oWVj�o��;Z�խ��0g�����W�XI�,��UL�{�cW�X�8�Ŭy���S�y�_5�W+*�vw�������/�|t���]0�w�I��� c~�8�Rfۥ��lwvS�C��6�����l�sT���C &�&CΙ\����,3i��ܠ�l�ڨ*������
��BToCd(7���Z}���7�mIoM��O'����=0�J}�v=��q޼�_% �A�[ׇ�����F��{P��C��� ��RZ��+�T�����Y�nqi^-̽�GEܶ0PZV���0�����_�~*x>uB��`'�n�����u��b/]6`�Pn�A��l4�sk�<,=�:umf�v�����\�:V�7����T5�ܹ��p���$1,�0�5 #�b�Wٹ�s[����n��պ�V���x�j.�بyd��l��^�)��� � ��#�0��	
��{����X*��M
4ϟ�+�ڗi�݁t������T�/��\�u`��D@֏?T��Hf	�Ip��:��xkA����,Ҷ��:��}���e{��C�`!�\�	�Ǝ~g�-2q�W<�@��)p�|��k:��	��pl9�-��� ���"Kء�o5�Ӓ5f���ps�
#��9���0N��l0���v�wh;@�YCo�m�pNC���D�l��1�!5�Cw��=��AU�� �
��_�|�Jx{�����}��0�>��F�Yw�����/�}4�u��#��n��K}�15@��E�n��^X�+�'Ι�H����	Q�kٮ����1tU�6j�v�8�A�w���lm~�D��p���E5ߺ���q���O=�x�1j/�Kn۰,��\<50nQwX�5�t�'�3Z{;���2���t�.��ls�נLRsι�=q�S?�����t��W;DЕ�����^�h���[Ȧ��J]�������aTq^~�K\��ªCֲ�50Vvg^�~3u�P3&0zR6{���ooZA{c���X����;^7b=��N��-�XHh�ݥǒ��
o���5�A,�^;@�<6ڏ;�Cs����t[ɃO�6%opjZ�8]�jM4��'sƷ�5ǉ��)��W�Cv�WF�-@���v����0�w	$*!@��� �8��ys�H��p|�;3�)�� ����C�}����Y>�k;�`&��"w��a��-��r�8Q��*���y{�w�9z�0z�s�Y^q�4	zX��\��y�p��u�p��\
�1i���WuY��,w�l�)�N��ju�.�Q�F/�ѭ����5 ����lH3}���d;6�@9yZt�4��T������H�ш�s�������Xǀб��+������p��مQ�S��&�!^�/)���z+��i�j�ܫ�m���	��>��	^��3y�������q��g*vv�^n*�sGJU��-p������9�{�M��dm{::�qڌ�i��`W|&���8����oT��s��x��A�I9L�=��=)-�9���Z�Gq�+��3
Yw��n�xX����1� �n�#9�r���ge��a�+D��(�e9��<���c�������]�ߤm�b({�8�v��%C���>�>��v_�K{��-g`rza�ӑ,����^�.�ORC)m���U50�O��������5�w���ؠ��r8Q��w�q��;�/�P��f^�9N�3�I�u �Lr�R�׸��,��K�I��^��W�t��{#����ו;�>��pvZ���L�]���L[;��*�mBi�-���T�,e�=����v����ڹ�Ώ�gϥ�_���PD2 �=���9�����7�����?e�"����?���o����-!�������ˆ�+>^��*]�l}��VB&{��Թj�"�綨^A���&ҪD�	v�3E�<�3o��e3�"φ�#j��r���_���CPy���swe3�)xޯ7��;���ZL�2�H��f��߽�H�Ď�S���_	��ۢ�yt�ju���s��9�1���8�����d��ϗ[b���z�W9/m��[=��
`�5�52�U1gi3�\j�;q�U/	��h��קٞOd�2��*}Ҭݍ��.��D/���{�����G�ƽ���̱��K��^����2�H=R��c0�{ڤn��c�����w�l�=d��36�߳��l\��X�}�с�8���ӂmI`B&K%�������J64�f�.畭m�QL$0�Շ�-C$��\�L}���@o*0�sfy���E0<��U:w=1�=B���{�ni��w��ƆW%������������G�
�;'g�eڷ�LXw����R�v���O	᦭�W�� �+J�ԇEkG�8�Ȩ"�P��Ćh��ZG%	x�vj.�]��R����&�햱�Q*��wh��tU|o�Lސ�yڤ}�쓮�-��j��]���0�oʱ�A�w���5��*��  ���>��aP��%S޿|����<�.9�*Lb��|��(�֞1m�Ř6��4�����l��2�9�=峕�6fҶ`�L�heN5>��	�j��y�����#<�0N�"uP^�Þ��Jtw��nKھ�/�}�/����³�/�س�P��s�a<�N��Z��X�x��j�ky�%۳S��o�p����C�L`w�	�Z&�:�t�rtA�;�d�+Ca{���'�\���h2�G�{�4�y ��m��{�7���,�_��E܇m�,a� �4md������=��?W6�3!��I���" ��s��'���1�D�U�<�!�T�,BUL;j�L^�f�<����mj�hz�V+�}�	���j*J�	Y�y�F�א�FR���b'�ӹ~ղ��ԼYk��a���-�~*���U��dmQ �j�Wj%FϹ�Z��.�~�z�%tˬ��ಭ��<;�S-Jd���{]�9�!��\��A��x]yJ���5�g*e�����
��6�� Բ�����1�L5+�ݸU[uZ��>����t�2��]����9����i�$�"ؕxR;X^o/��s��Ϋ\|�j[&酮�QԞ�K�ϖѦ�i�r:�]`G���t��b��x������|/�di���1,��*�>x,�����>�:�G	�μ{�Ƨ�����������o =�`��ZG$�D�����+�'�ȿbje��DG_tO��k΀���FCMʂ���>�T�۷TJ�0�!�F7X�m�A��,R��_��"��+h���җ���gT��=��\oW#";�œɶ��s<�6440g~Y���3̮�2����;:hs�$�e{o���0wt�pT�v)�����ZV=-�HKsC/+�aEQ��c!_�'i��d�XF�BcAk�~|��n�ϊ������l�}�,��?�M������ҽ�#���zn#/����`��;��9{��<�]R��NyV*�XÌ��ް���u����dKM��W}�{�'7jw�����&/*}"���?�az�>1�Sa���u�5����Ǥm�zl�NE&<�pV�����?E�r �H��6U�}��C�����Uz=��CqT�b�D�Nb<2���"�/�P��w	\\$�V
μ4.�~��nV2}<��|u_EbT���u3,9��[��o(f�
X��:~fkM�%߬8��[�{��%�a��ѐ��v��;��{��>[�\k��b�U�^��|�;�h��&����it����-�) E��Ae�^�R�#y5ܫ���L����l�{n�1J,K��j������9m�t��"S,s�{�\�����aAհe�AQ� >�8A�$�ȏ�m���o	Pm�C�K�"DF	�	 ߾�|o
�x�ެ�b�C��mzD�P�t�${���I
�(�x�u^S��<��^�HJr)�x�^��T��b�,���}r��	ў��;�s��=)i�}\�͆�*���e�%�|oL����1�K`vxX�;�2�Z�{�Um��n҃%5�欺=��u������n��1��F�>�#-p^xFyp��4q�������]�Y�o\j���FGM)k��++��Û����VC���>[�K���o��W|����Ǌ�x[>��=3:�����n��s@
��˞����/������new�����[�1��➆���+v	�S�^��X �˞|K��}�@4��,��^,�.�l�ڦk���������P���P%��:_��2d2Y&1�"�+c���cɼ��_�r=�'pI13����p��[	�l$�%�'�O��Ȫ��e�f�7'Y�=ZL�G$�)ޛ��E�^��sxt�a_{����,0A����3z������)��H�Ƶ�J^�)6���F��'y0��t��7k�r��䬿z�ɚ�(�^2oj��)��oj��gjdy�5vC!��S�[��N�;�N��wq΄�*^�V�v�c�Q���ص��R�jnb7�k-2�k{�@F��N������*�*�Ȣ�iϟ��ǿ�����W���|�S$8'[�0�CBc�m�r����_��;����E�G-�5��u�+����S9n�����}D��&���*�x� u��9a��G%��2f��S^a+qW��=�r`XbU�b�M	���85��ȁ���lMf�gsT���'����/NqX���H���7ˤ⃝����wZ�lP�;��H��=����Yў@>�e@Pa�Kո��w �C5��~N����o�������1^��x��r#3�_����.Z|�i��Ԛ`�"J(��OZ������ux����(��\���ve�g��p���F��\���Pv�;
�p�y}5��-��9@�3ܑm�#32�)���m�H��g@�.snF�Se��-�v�_�1�[F7��-���Yħ,�w}�`ڄ���e�ȁY&M�b
s�O��+�\�哒��|w�n(g)�9�B1�t�{��\�}*ڤ�!�z�d3M^� O@�S-s�O�Y���5�Qb5> '����r?�W��~	��R�ܖ�)��Hs'EG�������[L��N͎�Ϥދ)�`
Y�/7r57E�	�(�]�8U�/EνF��N��"hT�,��ܪv;�\��F��5֬1m�KƁǔ`9.BU�Scr�{���M��&�l���r��F������{�%3��*��
�i�qR|�;��-:�W	b����]՚5.�Y�:}e3Ҳ7h�/ �+.��N`S%G$����WW}�����A�j���[+y�ђ���	�N<��m��������Ի�d�&���}��E�OEw~]�f�z�\�N�H��oj��ٝ�љ2X����]�ɠ�{��V�߶��Y/:�MJ�9�Wu�4�r��
v�$K��e&.�[����x����xR����,BJ��)�/��{��Z�QA�^�"�ꐫ�e�έ�B�t�e�t�)ѭ����kB�C�^�V@�;����8m;՝4-��I-�)�����h^j�u	u*7�ӸS3��L3�R��,��"F��՘�U2���M穗�)�;��V�e�Z���[�-��;�f��)Z(vT�x�	),勶�M��-�N��-��;l��:v���O�·�Xc�Zk4`���z�%i�ڇ�s�z0Zں�I�-�,]��&e�u���ݜ�\p�z^��vg&�!1a]�AD�5.��sOy`j���Wk%�F�uw.��˸eeu{Dv��LhkN�:j��"BI�T]�K�3�T��xq��C�e*�-�*�^���z�ޣ�@�MS<�QݷR���f�RiGi}��w/Zթ��|y>�!��,ԖwRs�A���}�P�w�jB��;��C.Q��8�n��.g��ف`}�0���2��X.�5�A��)DKj��I-��n<��(�����牎���F�Ϧ��L��LȾ�wږ�T����FM^�#<�KB�	�.@w�?b$�}�\�����{j��)�u�!w��bv��Ԉ��"�uq U���=my�����Z�j'\Azu+��K��Z������8Z!�4bۆ.3`��3J��_
֦�QS4�}S]*J��^!�mh���3t�9�v���R
L�\5����j�k�|:�iKT��j����亳��NNc��ziˆ��e�D�c��h���3$������f��k�]�鈋\��1#5h��c�]'�ȋ
�;�U��H@��Y�Og���{t�s��Ř���0)�s���6�8�0�P�=��i��G���m����S��`0��DP�x�-<ՠ�X�fh�}N�@0�7t�+V\����m 9F���+��$T�wMҕ�E�x�vӷ�.ۀt�4h��y5kӊ�Z�0�+nӵ��� �&A'�~?�50e�QDKIK�eEDe�dRL�E3��������>>>>�}}~���ϰdPTe�o���Am�JAD5KT�EL�M5�dld�X�������|||}}}}~0������T�d�Q1U&YS�aFTAEY�T��f�lZdTU:�������|||}}}}~0���a�DMLQCW�f`dS�cM���ݢ��.���J&��� ��*��	�	�
V&��*/q�>�Tt�YZQ�3u`QT�Q��ZFM)�aUA�[�6f)Ud�U�Y8QQMPV����Sr�"J"� �"����h�2J�����(hb��
6\*�)h#q{��ʷ3�ɓwGj��ª�������SQm�PU1-daU�dgX�a�D���U314�1QQ[��SU5UTӓ�D�cDPDPufe�nl��733/��Q%W��TfaD�X�y ���OĀt��w2�si��M�O�E��8�ʓk�SmV��B�Wt�{Ԩ�%�%�bTY/w�RW��n�X�y��o����w�|���P��0�XB�%�@
��b��������=z_��^��@�d<�lϝ�at������VC8���+F��LSH7<직�;�YCC(0c��V!�[a�m��yO"ё#�q`Ҟj���.����&�D^��&k����e�g�ߠ�k�6ߩr���Z3�-��RaÇ�gD�9X2�����_�Š��Z�=��ٺ��D3�fO���1��uʹ��ԓ9���d��R��!�����F��F���R�i��^��`7��<�04Ba��N��
��Tw�S��C���G��vs�_��k��y�^�ﮅ{���4`3w<ö�T1Ynh[��t���R�X6}��5�g+S«�c	�tϰvbZ1+|�O�A��kt�M�-g��">�'�:�Ρ ���X� ��,f>�i�D��$`97�&�1���{��|��Y�-�}ۀYX��Չ3�Ad���a�^�dw�]ĉ�"��Q��S��e��� �.9`kCjF.�w`#t�$��|�9�B&w��_D8d���;b.՛�>Ç�S�7l_��v���L�4Bտ�.�s���t�[��&��ڭ�7�K+�'�� ��2ķ�y�>Zi�7�f��Z��[(�f�Ӈq��Ż�����.��/����WW�r{�[�~g���v|77��?A(P�L�rP���0d2D�i 3xx͵j��kx~8'Z(q5^d݁\�ǬG�37�,X�E'�|i�64���q-W���c��kuY��B�S�Ѱf��ڡ���D��V������m6��O��Wk�9Om�����=��Äb�C�ߣ/� kE-����fe�h	U2/alSm���Owc�F�6a�i��a(C� �����,��k���ݑ;�	0��]0��Mݞ*��nch��Ք��D.b�N6K�8���=�zQ�a1�m\�/�CϵJ��g������	�Qז<��SH?���6e�����Z_PF�W�O��ߖ��gT��ϩO7�V�v�;b�m�,�P���$M�G2���IF75�x�42�&Q$���G�������Z�T�\�5v_]��G�C/ީn�p*9���o����2��9�&4�����4;�Q�]�ؽȷ�k�M\,��a�%���i���K+��>&u��-r�<�T����A�Bd0�t%���s����={�֗���� 3;���]�P�����*�+��kk�΃ܲiJX� ��v"�F���b��v�Z���=����y,��l��ú(H�[.�t�Qm܄lኽY���������%b���]��s���������hiD�Kx��
�tζ�ۑ��\�X��
���?@�~���	��@�* �@4���e�	=���zo�j�d����%&I���4[���1i�&��|�<`>�Y޿	�|c#5V��� ckP�.ucU�_-Lus=CT�8\�����`� ���PL�A{'����S9�v=3�<*����՜u[�)Ǻ�^V�;�v�����]w���g!W�̉P�D�E�&�K̗S�L=��:��d�Z ����ˠ�#���⭤:5.���{�15�GgO�_ew�w��R�y��MG�j��*�jk�f�W�Jfע�q���t�?bv���>���'�]��%�}��� �y(�d�h&;�qO?Z�^��g����}�)�W�)��=w�5O�0=>���>�u������\Vx�L�_H=�
�:e�K"��7 ]O
0qڵ*Flsi!��k��3��x�f�`Y쭟!�F��6-p^xFys�:��o+��|�u�~Ә؇�Hv��ۖ�Aj��y6�Zy\��_Ӂ��@|��>��3]�<'ޞ�56�7��-dY<���9�O��*��g(m�7BFwHɯF0ts��g���^x6��>���}�4�k�Սy�-�ɿ�y�̥����Y�4����@l!J�r,k
��]���U3�9并"6�i�=�=�F�=w�Y��<�@B�䗧n��2I���z�B�{1[��̾��-�U�յtVƈz��{�0���LS% ŕ�
�����1(!��	�M_K��R'��s�c��}lҎX�q���-��+�ͼ�6��J�_�u�Pϼ�]7*"y�8�������	����%�=D<�Х��S�/2g��~i#��^�<�]�}h�EP�TXm�/�Y�e��u��vO� q�ZD�̷[���A�C�VP�p#��&��hή4H欵�*-��ݷ�.���^~r�9�u��Ϲ�mp�QKH�`��F�R&[�\y$�{,\'n�c�hW��ޟ��%N��~e��
�ӄ�"9�Ȝ�S�"�^��!��핵���Y�m�R Ko��7�<�����>{��v�0��2,4�rZ�����9��M���C��j�ݤ�;�!;8�ľ��Q�v|��g��%���hF3IWA���&вm���:��=�q�uG����_��j퍎�H�i�59��Ƽ	�-�Zg1�B��&�j-�,��6��r�?�2�v�'�+�K���j�oB�_EvEdT6� A�L���ߵ�&F��ͬ��G[Z��J��fȹt�(��\�vA)e����1�h}�|	*�k%߭���w��s��Պ�R��$qTP�m���t2��P�i�S�WHamޞu*V(�o{�����{�>sz;��~T������!ApIZ�P��}7�s�{�
��gw.��n�g�ۍ�D��+k������&���{��zsd�nz����osz�ֲֶ\��Xt9yO����K����v�cGܠ]���N��?qo�;Aw���8������)ٸűd6:D���L��|��h��>[b����߱���'�d��<�g��^oM!�P����`3Eb�/[1������T�ʵw�*o&3)[���VT���~�r ��my+ ���ʄ\��:k&ޙL$wT����7j�m�ܾ�U��[�K<��A�hi���㝜�Äٯm�b5j`�(�TXwf����{�s͸mӯ�CZƫJ'�N�Ǟ�8���3�[��X4q%�0�׻b�H���{be�Z��)�&.NZ0� Q�/EGs����Z�[�{[� h���	>[�r=�⛟b{�8;����B��QX;T���D��8ŗ��Aޞt`��R@��}l'��ɾ���@>�\������v��GM��kݎN(�ƺ�<�p^�&�q��}�����Ym��͠���,Ǌ�IU���5���Y�[��d0�S��sJ,f�D�~4�]������ܼ�R�2�^EL��YuD�U��v(Q��8zٻY{B;�%8�s��r�V]�5���\;/L{�����V{VP�9�{�z�����NA?�U��'��ݣ��#�3�P�+w�a3���cL��������+�?��&V-K�y����0|!@w�yc�ʦ�<Y�1�:��pJ��a�����3���]
I��E.�]}��WVsCQu��8z��D~�ƚf{�q�k��kȼ��:��N���u�Q���4�ZA{�� _I�3zB��%X���K�d��{3�}�`�%~��'�r���Y�SG(	�J��z��<���q�L�J�/�.�W�ew�}��\�H;B�gצ��_����5w)d��/Ԡ§��ʮ�f-���[�jv��͎���*.�lNW����Z����k�	�)��	U2.����,�aO��+Pte����l���b�T@Y�酑o� O4��לr=g��}�=?D�L,%R���Kh���{�������R�_ܞ�kZhu2fo�!p/�c���1�^ыYH|����z�]{�	��a�<�I���3k��Y�Q�æ�8��v��ˆ�?i���3l>���aPB�?�,淞����Y�u8�k�o�g�Ɖ�q�i9%���oBse�'@�K�6�9;�$�����V<���2?m��5I� �����vaAm���ݥ�������{�|�g��<��a�#�C�02�� �#J��#+"_=�DZ��ѹ0y�;o=��3R2�QB!�� (�Ab�����H��s ����'d�����x�6�6;����u�	x����T��5Ay��]�cf�[g*�n��𖑶���(Q�⤱]��=���`�ؘ�L�`K����յD(Ⱦz����/-�1�4���(�����C�_#S;��4�<d˾O�>�.���{|�K�����gP{e	=K��z�='�Fl�e�ғ儧��Kdd�w�6�C������劥��Qu0'<|"5�� �ά8{��(�7t�`-��k�&�ޥ�y��M:[�7�ά��DMm�|�8ϘE�\ᨂ*(c�e6�Ν�V�[f�/+��cp����<�ў����ʾ�i�6���5�P��Lc0��\�"s���Y����8e-vc��N���N��m�L�i[HyF���;6��N��u� �k����:�����)���}�Ŀ�^Xm�Jk՝�9@	�9Ne�j�D@=�i�+2�S��9�U�Fo��)�����U;��Ќo�L?�0�;����t۬Ĳm����K�-�ٰg���Z�7d��\�Y&�d�oҎi��4��ZKr��NY94���������{�6;�E����0�Ƈğ@��~���3�/SN����p�*<��5iV�/�q�2��в������W5��y�>}��{|��{��B��$qF�7�����}�{���?~s{����n�{k�]���e�.�&�
[#��Qm����.��5%�Gp�����(��:`K^�zs��]���W�<����gI�G��y��k��HP�b|}�{��O7���8AD��|&q[=����XØ���X����F���z��vX��kIި����˔�h�kymCV��b�����J���+졷�I�����ь:�����Rw�!ש�ץ�>t��p!�����^��ak����#�נ���ww��c�*l �Sf��k�����qє'�Db�M]����r��a5%�cә��+�&_��bי'�Ɗ{�I�3W��,%��������O/u_ԺX��P��Ӥe�ץyl�5@��H�K��a�9{�o.�4cY�\Lc?�/��[1�V�W�>}�f����(���k1�fj�ˆVɰTv�=���ؤ��
41��gM4����ѯ�¼����|V�ԉ�10�k�'}�����f��g�H%C5�а�%�_8�a��3E�z���d�͌Ƨ��e���}ɑ�MD����w����gsp>w�4�|nx���������v��\�"	��с0v��{r-V-�$��H����b�Ð���s{gg+���e�����lN���أ��VP	Lۏws�L�Ɍ8$ѷ� ~���%)�!��J�H�2<�%VjN��W�������ڲ�}�q����d`i*��hOC�^=���Ԥ53��ͭلe��O{" �o蘶)���N�9q�^��7="1�AK,00y�gp��]z�me�K��R��#	��e�s�=P��#d��h����6Ma��-=�����U��ᾖ��o���K��_؁����K�<���Sګoe�),�nokm;^0������&��,k��
�Sl%�=�� �4X�
�s����5<��Ezi�mx�o(ڹ�zNNQ^	�Ƶ�n�2�1I����*o]�{�S/�u��oF�[6��C�P ����Vm�f3�� �3Ed�0~muk�Rm�*���O���W�d�[�0���۞��!;D�++4��^�Y<��t�Ւk.�z���'�b�s�e�=T2��*U�6V@Y{�����cT����|�?Y��5������Im�>u+���6\¯�k=��#O�k�{gq
��$dlZ�69~;Q�⡅N����9���W��/�n,���^'P�#]l���C��HW��+?����약e�U�WX��$��a縲خ�QH��+�b�H�b����&}Oݍ ���.��1��
�N`�i})�^.��0n|�&�e�Ü]J6���r��9a��1Y��� �P��P(C������w����4^D��Ռ>q�d���'آ�i��jr8n��PhԒN�l#=�)����������&�+M�qy����e�zt��74��D�"c~<3�
)y�Wq�&3?I���:q8v=�9Լ�{�z�z}�#cR�֠5H�֑�-�Lf�7���ո�0��܊�m���Mp�H��й�����jq��b_Oa�ܬ���q���Ӿ�]]����y�ȼ4�˽�?<�d�aa?�u�X�:"�xY�3]�
��{C��U���i�O��)A��L^K����O<�|�����2s���ƮK"GZ������"�4�-	f"WM�3��W�F���L�6�~��c�}�x��&[��۫����{^�s9���ׇZ���{�񡳙- ��n��9�	Ó�hσ��%t*�Y۸S����6Ȳj��m}S,/�&�[�*+(V+�3�=�S���J͙6.����g�f��2o����rj��̓�+ɫ΢�uCѽ�L��K{'�Y�v��m� 0EA��\���]�I��[D�x3�e�DH(sgW'B���L6�iݯ����}V2`x[}FV�1N�delݪZ�5��a8Vc���,Q��G��OT�^�e�1��I�2�KIw�=2���]5Y�4�t�_!m�ty��^�K�\ْή���������5�h�J஽�Kn�mrt���;7��4�<YEJ���k8�Q�8m��PǷ����bB�LH^#a&b��7%�j�WJ�)��qj�:��ޗ�M]�O��Z�=������,S���yob��·���cz<Z����s���Q�A}C�����u1�4ls�9��Șm�K�l;��W�%�i�s�Y��jp��(Q4��G��[�IZ�ytt@嘏<9F��+Qإ�z8�N�R�_PK!U�Ƹ�,�X6�x3ԡBWIq�R8d�1���w8e�qe�E������{��M��V^�yi�۝
�̵"UIK!�|]	7��5������6Ѯuh�NJ�gNT�H��C��Ou�9d�1������sK�eY�т��� ��&vX���4ݕt��Hs��R�恷xtmj�-(��곓9ڃ��5v���O&Ϭ����202�;��#�m�+rV�8b�z�ܫ�}(�`^���Y����6��m�o���5�M��2��o�\�C��`-̮�N\�tVNշ����F[�.L@۰���ŊB�WŒ���VC��?q�62%�Ukw �<���$h�L '#���}.�kz>�7}cH�9[ѽv{P�FbfBqmP{u>�u�g��θw׺����E��y�lu����P�k��ˬ|�6bYb�jl�&�	m�r�����s��p��_bO�fFr�N[��Z��8��,݁U\J�4Kڳ���c�\;W>��Rg�[�X�=뭲�6N�9;�Mʆ���R��v!���u�om��M�%���hX���ʺx8fJ�N�vLr.�����l\K��U�WU��´2[�:�u.��{��p���щV��m_u������\�2�d�:E��c���
5ˋ%�̗�4Y�
�k+�=/J��a��4�dn-zU6�����v^]e�[Q�\Gu�v���m�Y/B�v����	�j�]��Ǎiv�eg���o��wI��~�f��eKn��2���ءEMQ^�:=���ᤒ� ��S�]O���}�yi0�4�!�P��n�`�2��/�����ד5�*�1ve��ˮ�z�2��C��B̏J�kr�M����#:�&v�����ݮ�>Kj�����3%#:?�t��g��������ھ�8��j�[���ij��^G�ZN��̾2X�Z��R��3٠�cR�tVwq^�QM�GpLb���2].쩶�XS���|�]M0��![�< �~@�'R&����ED�s�M�)(i�(h���a�ݑAC����|z{{�����_�>��O�K��EIf9-ffa�[9U��LAA��6�rd�"��lu��������������Ϭ�DL���os32�2�@ʲ2-�v��
(
j(���Ȩ��36֦�z�+�__^���ߏ��������ϡ�P\����C�Ȫ��,�*,����hL��#p�H�0�06؉:��������	�a"�,*�Ĩ����&� �$�(�2(i)*�kw��"�(���6J
:�Ƣ��-�`�6:�.�	�J+,�
�)�0�&C$�#HȪi(�-�*�k3&�s2̢�'%���Ȣ�"J���2������(�-����y���&E,SE3��-15E5M7V-Rfc�&KU��PS�a�E�����A�Md6�4n`Dll%�U4m�F��F�$�d0��� a6XD����aJE)m6�P4����ys���ɷ.a�3�$���h��,�=�F=����o2QE�]`H���	����s��8y��y�N�"b��RO��F�D�p� �)�� p��@��%#@�Ʌ�_�7$�Q��8C&A���w�޿@>��0BCF  �13�8LP��;e+���0�JFE�aH�d�����$�߻�-�(�f|�x���<]_��o�~��̊U�\�.�nml��;W�G���>*`��ȁx��q��]z &Z��v�khU�<��x;�L�.ևQ�;n���-�/T3�-k��M�Y�m�Ƶ���8jL >��)����lx�8� �c��[w���ѷ���ؼ���1�Ԕ��zh�a��YL��@񎳚�C�����7�OJZ�[)�WܨG<��F�v�";���g���������3����6u֔Nwl�Ur�DF27S-�`CXk�[���Tsr��B��f{�3lNk�wVP�ֹ)�8� ᚶ����B^z@�y��m��8�0�&�[<Щeyڧ{4����>\������%�D>�$e�::��^���KU�1�}����	�[2�q��ӝW׳���w�L�Y��U&S�ߥJ��kNuf�e�a��!F�|c8�j+6���nY�ѝ���,Y��z��6�35�K��D@5�s���9�PF���d{�x��8&I��Wdv��3����׼8<�c��C�=¶�!�.��m�ِJx^]�=���(�pp���?Db�d�ok)��ζ�r].�,��wD��e59^��PŨ?�C�h�r���ѽm����뾱n���S#S�i�C�2�#�I@� ���^�t$35�3�_P�g	�{�f���/��;�W����9
�'z�̏A��vZaz~��`��o�E�ُ��s�\;@��Nܺ�>� E�ƒ��:5.�9ٵhi�MG��oRt#]y�3�|P=3�`z�y�gC��Rf�@3��v�M��p݆Θ�mGCo'��{�H]��S��3�P�p�l�t�ܘ�+z�� ŧ�,�2k��n�N���)��z�	��,�1�[^��ȕ���,���<J�Eە�W)�c�ז���<B�t{4��fa�\�gb��h�%�\��}XdSe ����Ő�V�˱��^����茵�PΤ%w#��까���+��8����a�G���:ЮN�j��am���kW�d��Pka�4y=ь�E�N�9U��zص&�����c�s�5L�6��c��'�n���1�Y�F���|7c<ݰ�q��,��x���Ϊx-3�+�q�/���9r��1�LX�m��X�]��}Kv�ț�r�N���C���C3��+��^�.���^ӈk}=/C��2`-#$�8�2�效��Xr�ҙc
k�'#4��ǽ^��k|���SW��ɛnS��wrwq�<�{�Vtf-�k���l�ر��U}thV��,�-�9T�u�ӛ�/�跱oQ�����V�NG3gT۵��dGS���e�F�|w�g�˾��Ϛw���u���?#=�2��d��D�)���~7��>���'g�����:?�#��l^DK��������
~h��wn��c�%_0;3�G>B!��R��|=�y�8�э���"#X��s˞T!�ףP�ʹV�ذRw)�)�+sc8^�L��e��thv�L�]���"H�es�l��wNU�i��v�U��ǽ_{׽���?�K�?�`�P^�/`�3�w���mr.��xs�R��E����iD��=�t���%g�y����g,j٠u+����:k�e�;�_���/��o�k�;iz�xlN�"|�ΫE��B�˜�B��N(9����m�1����T�U.kIk������>uCo9�:Q}��V���	���b������������OOތ܌Wk����kK��!޽&m�O��k��{�.��u�r)J��{WZ�����p�vt��E��g<��0;_w�B��VF�{#j�h�*��{a�������̻N��*唫3y�l�;����L���sг�l�IM�u�H��u�������K��K�Oo\|�pS�;�ԗ�^:Цu��<�QK��U������Ro?a��Zk/!���}i�)ɇ�]K�vMY���������U��G'+�t2*�K5S���u�\��x�֫���Sn+H	�I.�h5��_]}u���O�37��^%�kLӬ�w����q#���R�`5��1�ze'ң�x��3^φ�Т�L�
);gM+-s�r�c�,��j3������,�f�b��ޯX�����&)�?g��wm�Ke����|ZYD�N��燤w���8�!�=$�^�pe�6送|d>�&�R[���ʂZ����阌ZֽK��X*vr�]�����T�����h���:���E~�ʁ�*W]Vo]�E��������:��(t�V��I�2��:��B�n��A��n`޷��D��P4��Ը��1��!�Q���9a�-k�j.ͽp�O*�'����0�:��W~��HL���Cu���ӚJ���I��8i�hcOA����0m�X��&���7�Ϻ7��-���&!���B�'�X�[����;4���ƞ������O���=S��������	Y�����`Z��G��
�/�kb�iB�Wy;�f�♜8+�y	�>���g������V/%�X=�OG��8��1A��fDP�]����7�䩪���X�I9�[�f�F-7�n�c��Z�9�Y��޻2�D)�nɡ�/'$M]];���Wb�,˞zOE�u����28�N�Q�3F�n���������^j�۔��ކ���.��|?� ��C ~*J���=ڳ2��f�>��ODm�h�d�	�ec6�==!�5������|�����Q&ro�HtT
��Yȩ2��1��3S9M/�І�}e q��-#$j�w(�e�
�j׆��:jb�Zʎ���ff�]�M;����T����B%o��~R�d;M���y�=`��p��ʁ�HS�bk����I��-5���}�`Y]Do�OSǹ���CuK��,��Uk{J��Dr��ק����?v����_�l )�	r�ht�^}N65�N��c�Ʃ��['��-`��o�kZ��z���1�{��:H-�At����</��S&cf,5r�����Kz������T��9���]�`�f���h5;=L���w@�<s֮yX��U�M��ȋ��1�r�.��>7�@�X�7<�/������`m�i��l��;�]oY�q�/�.������xj�]:޵�F�qU���sJ�s#u�{nm�/��#`kzk0E�y�M�J�xyW��ی���Љ��㾿�C����$:G����{��`@cT�;�.�5�ԉE��1��:���*.��h��]D�I�{@�u^�"�\�w+A���ZLp�GH=4��q����������{�Q�|�_Vن$��y�H�f�Z��8pF*y�F���ںΔ˕��*#��.Ky�9ל��w�7����fG .s����̏�葁�>\�����5xK�k>tK]�V: ���}0�wFҹza'[�.�B�Os��R˥����<��0���)���S5ŝSy@�`v���$�L�:��J������a� �a+(	�_O��\5�p2�'!��p�C�0*B�/X��^m�Q;T���y�g�>l
kd6"ӣ�3A���*�|
dq$w�&�����̜=�1�N�$���ۆ�
����P��`U�{V1���Nw���K��rO79�K��A����y�9w~���N���""bۍ��4�v��Ɲ�ܡ>�̻i)c�sP���Ә4ȵ�����u�W|�cU�j�Oꂝ��s��3�q����k�p�|M���Nfg+*�oey+���p ��]v��)�<X�B�;��J�q;���f�gB������,mن[�t��\�zZ���c��5�v�< f���|B��1���l��G;��]�nR�i۶[/���C������w�Ncݥ8��yˆ��v�D�����w]�Uj�^����L�F��H�2:���k@��e�\�M��:�UaV��-Ύ�^���%R'�P��[�JW#�k/S�DI m�A?aG뫻�-(N�Q�]�=;qnK	K�����.����OeL�g*W��A����۝}[W���&�ב��@�&�q��3�����-+��s�0n��1��q��F�dAP����{jv�0>���|n��ٖ:���fC;{$-{v���]��S/!_�\w;d@f�*u�>��bØ����ef�n�܋e�8���f;,��=���\���1��4��m�wT�s�c��Qͳy}�[���7�Y�E�7���� �\#L�]���;C �S�����Ȩs.&LT����]YC�������m�
aU��@&� ߷�*��WA�u�đ ����#��&_W������R��o{Jt8�� ^yS��y4�^*KAz�͟]w������G���F�GW���v;PM���AˁK�p裰�(�Wt�-.�mAgH٠j��1m��ff���� ��η;�V8l�U�Iz���AG����ff�'�T5���ؿo\c�mA�.+��	�~fm:�jc֌���#�#�{��\C��$�$9`�\3ZsY^�nE�Gl��jd����;���I}��c�=D찛�N�" ��,�M2��_o�Ii����G������IY�}�(޻�hW:	Z q�5���=��wa%�V�^��&bHu�7C���Ǚ
�8)�vSE�S����w3-a�7���w�M(��Kץt�)v�T�e�ꜚ�*5���z�t�4��:�ze�_2	��K�*�9��������|��3�������ĺy҄F��,�WA�͗���w��P,��3�PU�a�Cm�2���Ȗ����	�G�������KK�r����,��&8�<\��-R���'�,��u�VW��Dumǹ���,cu��82���AWB��ՄQ�3�S�S��7>+�_gg*��-Z]i��Ȟ�X�|`O"��t��7a1�1I�n{(>�7�.�ݧa����F�6��W:��]3=>7�G�p8\隔csg�:D�ze'�	O�[	B������5�3��u�6���H�����$f�a���+ �.��W��A�͘��LS.~5;�C7(L�oa�+Җb��L[�s��;�@�,��	~��4��@�aZ!��Cɝ	z��V�=�k�A�]svyG7%�b����j��H9A���cǝT)�Ѥ��sTNZ ���;ѳv���!U�/�L�KQ��-��'�g�q������=�6��T	)������=�o���Y�)7)0��t��7\e�d������:�\��n�:���}z�ϥ+��n��u�W5��������i^�#E����T�5�ژ��y%�\�y>F�*��H�� '�+��t]=Huؗ>�������.���e��s+CI��e�S�����v��x��^i��۳��O��>?~C��% bG���n�e�s��۝|��yӷ�zh�A%Ɗ�2����f>���A?�'<�W�qg��=����7��ny)1�^�R$#C[��Av^< �1`���׸y��_�X]�
||��`龻�b�Ɨ�TXX&1����xgv��~W3�Y���Z�L7W�)�)���GP�@/�u����`��y�݈�Dw7h��^x��<���gAl&{�]4n��������{��^��#\���lxg�3h�3t4]t�a��S2�q��bo!�Fm�s�:u��#b%��>���<Ȩ���G7;.^vn�yTWQ[�+�ѹ	�=r�h�3|� �=�/2c�F�t�w�FŌ�}�&�2�zT��E��,���T��4���~/��<w��%��a�{n&�~�[�8f���{�N�>�K?3+�1�}s�h
�;��e�׎D��V��sE��U�3��w��$l0F�y����'�y+�Tl��U�<v��v��}"��[8�6�'��ٵ�H����d�7E�%��x�I�C�jEעe��a���Z�&��ml��')�r��įp��_Mܗe�f�()������I�����ݤ�W�q��D+m<"f�皂��H7�/2]H;�nބ����u�Λ������
�η~��I��c+���dkg���4I��SF�u�:ޓ
�i֛}��:�c���&���F��d�W����>?<���Qg�Q̥9+���SE���I�L{��v}^�r�90�]"��U��4s㓂um�X���3�w
u�K%�C�ݞ��g��yO�S������)P��[M� 8��BWMi��؅N�Y{����<6юo]�4"�\�è�[a̍פ���?z��j�eX�������+8�+蟈�6�w���E��7��T�p�Eܶ2xn4n�b;(ũ��b��9��X'|P�h7�4(-��uP�y�T����D���R��Ah'u�ʍ��i�2��������� ��`D:���6�?W�O ׾�s
�6\���0mm��wl1I{��Q��%�}���8��)���H�_������/X�t&]�Z���
����#$2����E��H�34]�z,40��&a���d�a��M�f,�7O|]�'�����+�>�fP��8-��g��e�0����������Jŕ�ܣ�t�Ϧ�՞v�ϋ~�Js��hr�Q�alU4U�F2�lv�KTee�(��XXO�Lr	{��q����{ʶ[�S�வS�O�[W���+8����.[��۳I'9l�mʂ�3Ud�7�W�Fi���ݨ�'pFpќy<��7
�V(��Y�_2�>�&ϡ+ �9� �Q�2�%��'�LdA֞K E[�b�8��JGu��K���3�#���W�*:X8�Ҽ��I�F�I�7]�*T�,f�9��I�e·6���7��u+jon^��h���/uEYo��̚��r��|���:��,˻	��1�v5�]�u�V�k�����tDY�$�@qB�wfgX}���e�,Cu���ku ����Mՙ`�[�����[��4B����\�8rv��g;4�5�v�5��V�!�r��rHA�nE C�}�{ͨ��R��t.�չYǨH��ic.���r�\�N�0n��g)���Я.b��guJ3���x���!�G:@�Y��4AVB��ъb��<���r���N`�Gi'���������}^�L^;i�Y��g�X����;��oIv�nS!&l+���u�%d�\��o�[m�+�w�Zr�H�Cv�d��)�	5�wx��E�Bɮ�R{/x��'j�f:<\7��n�V� A�_�����멣�������W��-�k��M�zMnt�[N��X���c�|�s�s��*�«ʇ��'O]�,�qT��f�Ap��iś�d���,V��:�z��Z�#��t�����&^u
 �K&i�rAw�P�<�3�C�#;�վ���s�z�	h��.m�+���vg3�-�Fe�U���p8^`[{6^cP���U�5�@է��ng;�#]����Mh ���p��2����#�P��[��($��i���xyD=��Z���.��r�e����6jt���S�V��YC�,�ї��7L���D�-:�ӷ* �4���d���6Kұg[�ZX�U�\+�M�bb}���,D4��Q�)p5��I�A�֊S�_Q{:Ǝ���X���	�I`)T�ں���g1
�2I�C��kw�ɱ�0��o\������S�&^m*bR ^��2��y�W��[t�/i�$=$��6h��9�fv���`̩]iB�[U����IX���e" �����k@e�v������ux��qݱ� ΒT:��ʡX��<i��'R�yi�[/㥫�*Yj������.��ע��V�����1\.��W7��n��E7����O-���Dn!9H�U�k{g��wt�s��ҼU��l[!w"f)�ʰf�C���7��A�4$u�1���TހU7#�<�*ͭW���X�����¾!b���0�E5�|���Zj�t�JM�h �c,�qr
�i���ǧ�����������Y�� ʃ*�"[���Z߸mAKDT�[��U��s��c��oooooo�����׶}}q�ʲC �2$
()�1(�e@E��Y%0Q)T�hz��������|~���>����g�eKE5[���f�Q%9���"&(�*L�\�j���7r�"�L�����p�sb�����2�1�r�c3'+32L��*����7Qu�啓�nA�nePVY�de$�LEm��g�[u,����0#�r��3,ZKp�p�!�����(�0����0��Ʃz��>A�+w�d��`R��LE��|�W(�s3"������0�q"ʪ%0��&�vM�b�(�b����:�h����2��0�"(���cs
j-���H6l�ɦ�͝�Ҥ��R����ʀ�����2L�*v�(� �w��;��v%G6⠳f�]�`�}�Q�5&�%3έqt��
�����K�����2��0�@�y���:��4����D�����EZ�ՂSg�HS�����#^���/4)L��;���z�M�Y6ڼ�W���a����<9�i����$l��`�lCV#�=���,�y��J�4�~�(>n"{�j���~�n�YB�aK�f��g�e�H��\��̾���[&J�
·tW-ڥ��x�^g�y��=��I��H��IV��{gm�h��.uѳ0�ݾ��jvc���^�sJ`�A��0��^usH�,�{�0�JOa(M�����Ul5�yml��������-�XJ�1�3/.�y��M��C�m}oP�L�/�3e%:�^qˠ���W)ܬ����f�<�4��ۋ�ԡ|B���	��*����i��9W�P��\��ǖ��E��-������a�5,�v�l`��,!81�B��"������y� �����#a�S�����]3��^YD<Ӯke�JK%�g��B)��1�������S��W�.����a�A���y��	CW0�[<О��g�L7�[�j��B8�d�_�=G˧��U������e~��J5�o��|8�}��长p��:�FqwJʼ���:��w0����0?a��[�����ȏ+O$F�T���CY�i}le�i�}br?iM"��l1ԾJM�>�Z�B.�[�ƚ�Vhu\��͇�?|?� ���������_��������zm��9\rq���s�>�����4�]�i$NI70��wY�7�Y.��;��H�4*�hX�B�ܧi�v���|���9����b��9X{�O�9����4Q���������z��p�d���>���'�J�{�9�Lv�\���x*P��o�s����P�o�&;�>[ o�S����F��h���p��I���. En�.�c5�Q����A��ͻ��G�Tt<��|2'ѐ�S�[�SP��{��|���<61n��{�2���m�(7X0!�F����ݗ6;���|Ħ��{�Y�ӯMp��k�뫧Pb�H`�н�����������dC�=���)���7+��Ԧ�P�v�3z2,(��}�j������k�kj݄Ǯa�Oַ(iJo��l�����{�f�'���m?Z����h-�񨶘s���5�S�Z�l�
脟,%;#�����]5��%�M2�\ZvPθ�zkw��=8��vGà���	g�uR�9�KgO�l��Lcw�LH�RM~���"����Ok���RÖV���wYoC�b�8���^jy��sk�	1����u��Hu��!��-	��?l�rp�����V��U�o��Q�|r^훃|adt[�wי˽��lm^d8�8Uj���hu�s^e�W��|H��_��P( [��+ݿ#��/4�E*�	��&��N����
�ȃϿ�]�~�����ܱ�޷��jˋ�ڙ�>��ϯ����a��P)��72wz�)s������M��S����(�<��E����ʰ�~<�#w��,۷.���lQ�x��4�zSO�����&\P&�s�p�r�G0��)��6�;�f�O�k\�9�*�nE�������>!S��H�hVg*0�����Tw8�	Ia"ֲֺ���p���20Ÿ����`,����-z��o=	yc1������ԌŹ�>��^F��Q�.T6�MM��.Av�>Li.��{�<9�(�=4�\N	}j�v��Ѷ5^LMR�F{�be��T����Ì�S���/���lM�=��g���yF�V����$5�?0M]\�s-b��Fk�q��9U�9� �S+i�����_J��Y���W$�0亙wG_�E���~�_O�X�OM��O͇�2�������`ܢ��ع�p�ѭ��,��.�k�v�m>z�1�7�sj� ���T9��/�	�=�N'!år�/׵.А�� ��vؿٱGK��Y�oc��v�΁���ó%Ŧ6���\DB���Rrs�ˢ���U�
�g��/��o��̫
��z�;7��rLP�)����0�@��RH���vg9��X<�g\=$���1ƹ���r�׮������H9]���=Y'�����>y��B!�%:>�2�9�"Uq��h%t*}�cV�����<&x��N���Mz�%�%f��:6І��q�s�eP��ƨb�Ĳ�1B�H�Qn�uWϔ��Hr��w�qZ�����50���)l�@s�aǤri��M��f.��7tKn�Tĺ=��U9.�E�@��up�+MH�p�k���UfsWdr�g؅c�*�|�k�]�8���&��l�*���M�q�l��05�}m	4;��g�b��FiR�/(��ɤFt�C��)��^܁�Z�Tsu�c�\��z޵���M�K��z���S �=�x6�a��x��y>��K5�4#��NC��[ndn���tj�9w-�Y��O(w^�g��� B�����<�*C�_��m���ѱʀ�AO�֣2i.���w����<��1��y�s���� ~|�?p��P�Y���x���0Wy�w�t��Ó�c�H$֚�D|H:y�����t_say��'�\�ʨ���}
gDʫנL?αc"�>�|E�^��8#�T��QWs��8���hVn'��`���h�:�ug�H����;�z^��KY��:-�FU�$��+n|f��..9:�L&�����l�w��C[Ť�J��~>?����K�,I�!h��8��	�����>�؇FO�� Zg\�u�{�ST��#��eE�4�1���3���������e��&x9��]>�o-��`�+HU��&������/��n��͢C�e]<d%�]��tfW�ۧ(m��5�u�BF	M��0���2el�\�ѓ9;ЩjT}�L�+�L���vy�p���w��(A�0�-��cY���5�+>�D]qY��z^c�ܓLzf�%��4i��()�_ӕ�g��gK�)�T�����Uk��2zɥ�k�����D�]���T���m~*�ߣ&�d8��u��&�H��ݝ����n:�)����2m��U_�~��=-�pq�qw��,%�qC����.f��Yu����v�P9x6��	���I��)ؔ]�%�;���� �Y�
$�z����}��kߴ���|��kAW^ ���B�'�kߒ�����-U���qr�ɦ��%�̮ȡԲ��m�Z��|a�O�����6�ؔk6����)�J�3�c�#���k�����k���yb��3��v[�������l���w��h���V�Wf�[��5������%�D_zQ������b����GT�F�![s�r��\{
b��>����K͜&�-j�����-[��+��+�_$�>�:qR�]������>9�/H���g�){_�x@��M5�.�|�wL.s!I�.�E�s����������_��a���vM`Ǯg�/i�y�Պ�#s�q:f���>����MY[��|d[	��)��@����l�ῼL�I�{@�"�3����<�5�	g����^Sg����]i���eK/qR*���,;��r{���g�|r�]��ī�b��L���+��L��~{36�V�,z��4;���uj�ΑJ�[��9l�8u<�1�.D��Z˷�k��h�$_ɒI����N{ξKj��s7�ڐ�!�LC�8"�cbE�>�ē9¹l
%зf݉���#;�`��>�M�K�W�w��g[���e��m�0]��V��D�Y�k[���s]�}����u�'��vܞ�?����e��C֥@[��ux����^��a5�e�t���9�Ʀ���3�)��Sn���?[+:5
���8˴VF���r�A0f��w��۸�/�^�G�&�t�ؠÓ�9�Wo6mbW����:i&�D�,D[���v��+R�<��]F���ur�x:�}��~޿|k��]`	�������Ջ�SQ�R}y���b����+��|{�og��R��^���j{&�\�T���g0ֵ�c��?.�u6SK��%?{��w֗b�Ɓ?�eFjA0�̉O����)��)S�tm�^Aa���Uț���\S>,��)�YY��{�G�̖|&a�/i��k�@x�^�I��>c�魳�Ѭy�R~[r3ASx�ߚ�n�d��D�ݎ�~Dz���W�f���u ��='�S[�@���2��Q�ǻ9�5���h#�sA�ᔽڸ=�v�H�5gڭ!��<4��v,�FH!��h�]t#�B܌�=�����y�=���c��G������̎��ґ� O[Gڨ�qY��^���]�7�0�Ϊ���7����T��	����7iR[�P�ç憮+S��I�8�^|�;e���n��Ow��y�̅5[��� ^��Re�j���H�d���j)��|���i�<�g�M��[i�G�g�3��4P�O�j��͓B��ʺQ�ٔ��*z�bPX,j�ju�;œ��o/{s��0�QD,�A�[��6�fN����1��	ye"/+�ڭ*�%&.(^��3.WF��kaW8˫z�x3�y�S���Z�`P���J�w����~xN��P]�J��ۜ}_�+����|��U�u�������S��u���.˓�q����=՘'rj���b)�3r����˾�|��M^�!��́�v1�+���)�^|�W�Fm� ʎ���؉���{-��Mӕ�t�ՌT����.�v_ ��-���<����شS=Z��ų����� q�0�^��^c!Ϻ)ґ>��B]���{du�Cwe��f&;�*��'�{�p��s�]�Չ�)A���|�����^���z���\�\���*&��KVb��V�;'w�3 �ֱ��s��As����֨L����Az���7.f�؇����(Jy�<Ai��ό4��S�~��b�o����`��[qk�l븏y&y�/p����'ϊ�Fo�L�b�w͑b��x�u�߻�X��
%��s�t{��ZbT}�Vl���f�B��}s��%�ۊX�Y�vbZ�]Ke������� FF�l�w�>)��~�{ז/=p��x���	vjxdwJ�y7�Kg|ǭh�y�L�L�tM�v�e��2[�8�2��)���`���
�uP]��B &Z댤��B�X�Kl����7 �F��C�AtÔ�m�
�n�Sl��f_�ᾡ�B��b�>_��/�Mi�=���\h���.q#�Η�ޗ�>����s~d���eZK�:k�K���-'���3���5�"��i<W
Mhcp��}�h��col�J� �Η��h�3/�>]�mD�_�T+]��G�F�[��Μ+���9�����X���X�gG�Nt���r��U'��������|�y|�3�T������'M^��>��S�k���FDH�K���Y�Ù�R)wS�?twK�`1����tu��L��~;����>6uzI�!��u�\2$v���^��(�^��o�����]^��({�7�ު�j�;�	�6�V��c�b���Z�j�`1y���]|�A�M3�7�@p�la;��� �K�ayM���W,rڳ2�2zzb�^ɏKOd�'����w��-�<ƻz���O�r+;���t��8�*7����-�#Z�����9�1_����v!��&6��Wq�k�Õ��3p��d�Y���*+�(����t7��l�q3|�⦱�@��})+���Ύb}t)��=���b���Z\[��m��h���N�9B�3R�خ���bz]t������m!�6�ˁ\D�bj�[`v��R��:#g�>���5��T���x��O:�^�(o���v��T��P���V1F�q�y�]���]jhg��D���_5���+�/V#�� ^��c��B�wM�����y���*яlb�h۳L�t9����������*�:�(�N�y+��6�J-��ٽ!K�>�ui�Vغ��Q���w�����
_s�a\"��a�я�܄߇�@�vn&&iGB�t���ɭ<2lВm�v}�_�4́���H7��DE�zQ�]����Ġ`����=�	�:�����Ĕ�{�O�*]e'�uW!u�P.d��.�yy���P��M���Q�$1���}���g�d�0���vE��{��2߳W.�zE�_�);?3}>���m}%�}!�0�֯>��`�����n�i��6�it`����!�	d,����a>�}A�G��\�.CsH��M>��v�_)awB]P&��T��3պ]~��e�b�O���{�b�hjM�"�^�9_D��Qx��O	�+b[g:q�zqWV���L�ʒU��2��j�]<�c��{�m��wmw��}�0���n�����6_��U�wv���GyУ�-9�"��Qa�vy�=[?]|;��>�5k�8Ű7��ȭ�˳��γ�̓��-{uM�л1�Ɔ�AN6ť�M��<`G�m�L�E;�j�a�w�z�W$��&�@w�;��wf]�s�����Cu߰˶�o@q��w��m2l����gC�N��t`� �x�y����ӷ���WWjFآ��nm��AU�N*�'J}�+r�������r�+tJ7R{�ٵ�fޘ�,)\H�r�-U)���*%wԘ�;�c��Z�u}�^�S�Zy��.�wF1�<�j.qrO%�͇Y���ʙ-f�%)I����i]Ǥt�|*#W�[c�\�w �@�dvSԧB����-Gq�N�Gj�����D�꽓��V��c3��rvt����h�`!W}�I�qv��%����{F���$:���X��_P����&�Ͱw\ł����ٴk�B�Q7�s�X�-γ��m���1F��"�ڸ����{h�{����;`j��4��~�zz��]�cA��m>�v�"��󺶅�1��Qt���G�	�u`� �U��1x�q�����p���5��W3y���xN�GnM�I�/\��n�����U��7s�Z_]gp���M��t�o��b5z+���� ��.b�:"����4��b^0�Vh�ݗ�Ⳏ8��i�V��#>T3j>��^(�4E��J5���-��T%Y�
�j�A���%j��α(��ւ�%�������<.���G%G��ى�$�J��D�qk�df�G��5�Mu�s��ޥ�j�T��w]Gd��\��)O5���6��~G%�{\t�����ėB�n����[�HA}�J��P��|�kL">(�@d`8�) �]
�+)�!	��-�e{���Y�妬�9ԯX�[.4��3��(p�]�P�Oeܩ���N�.��y�暽���b.�i���Jt&��e[3r��.ۨ��;�ru�[��YȒR����ͬ�<�H�[s�R��-y�T���d�A�(��
�u��c]ܺ���f��j�y�O������a�x��骵�[Ձ�]��P�и���7�]�o��bAu��c�܁�I�\���;A�y�"�iYk�ǆ�FY��W�>cN�=f:�]4��{��� w�0�떱Gv
jC�Fl�"�}��1�wj9u5W���uVP���[6�o���EL̜E5}��H����u!�uA\�Cy�.ȖqC9*�TlN]�j�n��u-דXx���\��[׶D�XM2��9sf�dB	NPa]�zhr�[�S�:��3��WE�OB�NvK.���U�i�Y��=�2�iH;f�s�07y��z�K�M1y��N��6�wrЦǁ�sd��[[��p�6�`�Uok�x�8�|Z�3i��.d���pxp�ǈ��X�kdet��'�_.��"I�:�����z�@�O6r"���qi-��N��ի�!�[�$m+#�3yw.ThՕ7(K��E�|���jV�0K�9�f��&���reuX��D�:gF�u�[�hQU��>F��JRTCE%4�����:�M���Cm� �2�)�c"u����������?__^�__Y�2�NY']f�d��NF�K�ܠbz� ���n]E�3��ǧ���������������=��������3%��r2��3a�*�L��r����$�26�q��ק��������믯����d^��AM��J�cNN�;K�����FNKT4��X�UR4�4ӕ��dҘI&>��5�V9�n.Y!��bR4�Y�EU��AM-D����ST�4���d�ٰ�e�Dd���F[l�m���L唁)�e��T��1��������3�$(��B��L�*	�s
ZM�$6�f�hlȂ�k"�m��l�3*w���,���t���b�r)(2r6����*�+b�i=���&�����i�6
6v�5��,�[3a�$�ȃ���f��Ό��!�2���(��~l%B`j� �.0���H,t�ծLoV�1�֖\ĕ��z�(Wk6�p���mU�����s����љ��F��g�j܎�\J6���4�LE�!YA�P�	|ZL�!q' .HڒH�E�JH��R6����	¤�5u#�Hb�$�Д�n|A/37cz΋�m�h�7M�H��?2�X�
Aw���la���B���p2R$�Ʉ&߻�!���W�D�����ט�B�}%�X�x����l�mO��z��4og��С����8Y�u]c��ܹ�C��~U���Liaa$����g�V1|O��ﺐ��T�Ӫ��f&k/v�1�2c�|f�U�if��?�Tl<�Ϟ̉�d�hVf��4gyD����ali�+��ld������g���T�j
;��r���fϺY��wz.)����
[j_�>���Y2��;;��`+�7�m���ɘx�'e�J� ����w����4��Y�}㆓���R82ik�����)?X[�6��47�g��k�5-��NӰ�wn�h��mE���z-�m������Х1��t�w}n�D�ʞx]�Xe�W��.�z�|��i�Y��"Ȭ�(o�~�x���0}`��A[��y��]�Nf߯���kG<A/��9��"��bL�LP������Y2׆��_eL�B����9����1ހ�Wms
��^��j��|<��&���'�hM㶠a�OS�O�ٔ?Y\uH�� ��;��zۄ�(vdak}O�vt��R�~�Y��!�����q"gKw��M��ZdF��"3xkn����%��h��o��?���?z^��&Z�1)�t�(E���c��#�\���WL��t�{�1P�u�olɱ�!�{'v�L	�ް��~0j��ˎ��N�>��H�)�y�eH�v)2�6���
0Y_TH�y<����y�V�2�GNl�ߎ��N�O���u5�>B�r_��زhU{yQ�6!?�2�RXC����A�o��u��`-kc3aA�%(y�	C�s���>�@�p�����p{ӯ�3�7��.wNr��G�ev>��ꮢ�Ɠΰ���7�(���=2׌�n:}�[�k���^ڐ�<ϯBMH�q�7{F[P�CG���+H/:��,"��]�]��m���k�ޘg�r��/���a3�v���n��jeb�7�3���񾪜�V_^������Y�D�}��#�E�;Fdr}k�GIn�R0H*m��	t��6a%{�����1���3���㯄#����}�c��+���$��Oc���jFN��p�G�~sy3��&<��DxTh�Rp�+�����)���ސ�·�����Eɷ�#EFڵ>��$��.���4��먗�|f4h�祚�����������s4p��y�D<����z7�<fLV������P�Iw���Z�ʉݭ3��xv��L	dq�1MJ ��
��}BM::�꺛�,nWm�27 4�Γu��iڻ?LTF}/�q@5'��"i�m�:�3a� f�����B��\�3��l�Q-�|��@�r���1�"ݙs˽�˽5���{�(	���_��VY*��]Z��ӭ�����2O~[�UM���;��}x׭�H-�P!s.2y<���w����qd[T�	�h�dN�\������a�u)���+�9�m�b����s�nF�3��.׭�˓�]ðP�km\���{L�|}&h���[iQ���c�,�c�;�����Q�8*<�0&"Q�6Uu�㽲��7�MO3�L�R�o_#"4qU�.�!�A�v�W��<��s��y�/(n86{Փ1�J 0�˵��O �CҽS�'8���/�x��8V�s�@6l��ᖲ�b#R��f��c
�\�ݮ�x�H��6ws�\�O(��-M���߲y�F6��2z�]{���l�������r	ۑG�$t��̡:o�H�]?42���Z�JH�ġ��� ,3sfV;n����p׏ax��Z�zW�o��+��[��.�+����7�#�3�r�R�X�T�!4|F��̔�*��ۀѝ�z+�t�
<Ý�Uz���Tn��^E�oxA&��f6a;���QAeK.
W�6K\���iJ۷>�bX��\�\
w��V��l���f�xυ.�T�jٶ�a���s�C��U��fm��Q���pѬʪ���{���ڥs��>_=����>}�$�DEW$���dL�k\Es_q����!�>���P>^�Z=������'�aQ&��x����1-�~��ٹû�e���{����6���w6�
����vcj=#����a�ȩ=..{��d>�+)���d^,��J0`�f�kn�:����gE�S��+��:�ԳA�;]�{j�R�.l[��ý�.슞��i���U˞j�Ro�wo��,�%~[�ֵC==d�=�<�3��<��2�cc�MpBؾ�ў����k+|MT�6�����e�D���c��(GR���lt�`�2.Ws&fz泻��X)�zf��KVǍ����#}�Q��<����ͧr��W1-����!�]��^EZ��fQ�C��+��8NN���kI�@�����3)��pg�a�/[O-�49��Eb�0��ZƫW��C]:�Op	�t�M��c#[K#ص[
8i��W���\��	Q�F_&��s�%�}� |{�(�Q(����n���X��2Z*�a�"�(Z���)����'�ޓg��>Kvx�+B@�0?���^��f�A�D)�W�ݪ*�(��ީ׬鑺ym��SKe������Ɯ��ڔ�"�BP��be�a׮�[��mo*�φ<3����%��k�`)�e���]������=��k��b�Ḵ6ur;�[�r����;4;�iv7j/7�\r��P.���#!����=�r�$�v�H�����S��̷l�5w[���g�s�.���,�Vf&�n��y�ƺȊ������S8Xy��Y"t�hq>�>
Ղ;i��m2ƟK�TC�r���5}�{����f�Ī�+�Y��/>ԆOr��M^|F�Ca���p-��]�^�`2�l�~�3�3���>؟(Ҷ*Nu)��g	�=!�4a��s5�;�5��J�O-L	M~���ҫ����~�G�"ݕ9r�O5�Y�N����md���*�c;���BսH�\Nq_��(���x2�
�@+ŀ�)PJ $�3$.�8�����L�2:����7�>�q{1�G�q��㵵�xn�q�����S��j�C/��]@�������r;CT��Uu^��@^7p�ݫn���޿�ׂ�;:��V���z���\x��WW>�W�5!���Y :[6E�ڬ�m���&u��s�i2�+4k���n�ԍk���p먿u����weCGE�c�䟊�&����i=�x�a*{��2���vQ6�s���&��6�zKvu_SR�Η�4����Ou-E�1݊v��^�L<���=�h��g�:�؇V#���ʄ�f�ћ����"����R<y��2�����ӽ·Ҏ�Z�$gyFv���>��<Y�<���<�ÛQK�'pe�\�E�!�<�W�D��R���>n���Z[R�@�3r�;�\���+ v)7��`��>�:���־��i���-�C�ϟl�8���C��Ѹ��d��Y�h���=�y>׮���,h5k�>��^O����X������~����г�^[��ѕ��û�)\,�,%��I��;��z��V�9kYUy����(��v�M����-�ԽakɇVd:w����&�%8_T]�Iy|CiC���_5N�\��\䂏����uu�vݼC2����7�Zԭ��]d�,���.��8�s��oɬ0kMƟ����"�Sޮ�ʇ�=w�G���T�H�M��}T�2���W�!�K[�[�V"��ؼ��I��R���<u�x���q�R*���	�
��}�(L�|<�.t�6,�x�j2�r����U�gr��ꌷ�U16�w���x��ܖhSJG4�^J�bT=��\�7��� Ӟ�B����ocdkY5�1�Ot��B�����޼V��$^2����s!�p§-f^��z�W�zc�=�#I1vw�d�5��L�XC���/�[в�VKy3h�잊�����5���@R�Ws�(�gaЮ��،��S��z��<�J���^<�
��<%wM�/#�\�V����O��[����h���V�� h�~^4C�_����]y�AnOUJ6U�є���1�6���ժ!�*6��("oo��b�oFz��5�'7R�T2�i���>X��֢~˩KO]#��]�n<~��3v�b��r擏싗Z�N�vV��4��mq�rTm�Vӵa[� S7k�2�v�l�;�k)����P�;[�&J7�����+����M�/��l\f#R��9*]�g-ֳ���I�j�z�U��D���-��9�p�P;��!�9�mv���y'���c�4{���v#A~Y�~^�پv��̡:|��&�t,�8��ފR��a��v,�I�)�c]�~k0Ot������с]UQ;�|�_�PܗK~����C"�Y���y��ᩎ�g�����)���{����k9��o���?�B�гѹ��2���y�|Kt4�64׉g�-� F�O�P2K
3P��O78�IB�oE���l�M{��=Y�>��!�T^��n|���q��.�����O,w���d�� �����-�5��<���%\w�[�jm]���}�K��[N���g��F-oH�W>�Kk�$�*��Y�X:��Jg�'���M�o�/���;w6���ǩ�>�)i�����sr��:�h�ǵ�k�O�gon����&8H?2�_"yE9�
��6�U�����͓/�Q�<��O3������p�	�=f�l��տ:x�G]ͼ�
�V]>+ۆ����������O.���3�_`�f'm���M2��C	cMRY�ճ����A7��)��w�o&3<���K��ٕ`�/NP��<x>NIiu#��wfC[�*�=S0b��A,i;"nl��f��z�נ���s��=WQ�jhf|�
��oM��Q�͖��=R�����bq��9�R]��AF��&�̳���z�1^;z�VCs�=�w�o�N�T5�D��$��	˽�;�{<a�rV��}�%�4Ĥ"���	����vR�<�Veg�t�XC30B����n�ŕ��߫���z�29ҡ�F=� �Y�	����L6��}:c�0i�>~m�o�h�g�Y���3!OMt�CG��ཥ�x̞	�"��n�3�l�kʑT���""��k�)<���<�͡C�_d��#:3�[[�oLK��,��+9���4��V���OCi�>��b Vs'u��4�%E��Z�7"���#���T5��팩:ɵB�k�-�z3�v��I5�(�ˡ��� ���!���`��1�֝CDm�:�f�k&��=���f�h�bf��鍺�0�p�\���4]��/fg7�m!�>9xN𣒝����=Se�����q �i�V56�}�ٯ6 �,(�<g��ٯ�=�u�W7t��M��5!�r��V̌�O-tͳ��騹����8Zx��-և��G��&t�Wy�<џ,�q9Z�»^�z17tvZ��V�i���Y��5!OՎ�0���u�׫�m���=W��^�ƍm�^�Uǜ���zXu��:]mG[=����ڏ���Ϲw��(l�*��5[���Y.��u~�+B s�}��y�IS �~�lU����\BO8��|WM#{B��T@j��sU9�\�s�T��}�bԉ��S�'x��Rz�M�\�o�Z'�T��'J���3�g=3P����a]��z(t�T
�*�wl@�e��f>)�Whv��g�u��y�.����~��r1>��D d�F�imqf��wZ۲n�a)��L�ߝ(��J݈�}ι�ll�����bUۖj_@�[�ͷȆ�٫��|���W|_m���%��
���:W3"3j�&�dfm�H$Tr����(�Q'7/����w�LSJ���a����pR�#f7�d��DF���_��p�n:���nd�����J�K���;�[5^��뫪��a�xy��r:�9v����>}�պ@�{g��[0c�	e�WZ��d�K.�l*j�i4m��\nj��R������F��J�_`B�"V-���������X-����F���b-���ue�����=@�"N�s�/{6	V�:C}��\6���#�C7%ܳ���oQ��f�:��i9�Hf/�zzR�;+�D��k��;uoJͻ�v�ʏ�r�{�]�Um����Q8,��b��
,�0GI�33�d��&���ǹT����&�<b�ܺj����8��������C*i�͆_Vء�{�6;��&=!W�Yɘ��������ntةO����	�)kB��9zk*�Z�4&�٩��ਠ7�zI�Y���,փ�����Tk+�w!�0�(�]�6�*V���CN�3J�+a�U�J�VO\�ڽ\�8��2��7���\68*�Pw�wz�mg62N��ʕu�u��X�(K�u1�����[�4l�v!},��y��<�77�+nS�bU��8�D���6igO�a`������d��[�h'�e�
�ؼ��E��7iVM*��4�4V����H����|%f���c���.G� @�ԷY�^Ǐֆ�٘���6W_E�tn#��#��p	XrE� %�Bu��l�x�ɉ˺}���LU0]v��G�ŗ��Y|l�G�o
��O��
]s�Ru�38��\y9!���)j�8z�{�5�W
����6����vﯚ�Q\:���?������2���ݽ�h{�R��ג�uK��'Ex(�7���!�8x�I�ɉ�Q�(�Z��2��۸�c9ٮͪ��eb�.�,�C!6/vN�b��C�;�Z��v2�v�4��]ƚS�
��1��{� �Xj���;r��+�w.�1q�Xz�i��ϵAܫ�eۦ�z��B=A�CE�uڛg��zT�ж� i�xRa>�j��A���(V_G��7���8�jp^9���W)V0��e[�����X��'�P���i^%�MС�&�ʳ@���8uMY����d��|$%"S%�%�n�Y�,>yj�'��v*՗�.ٶQEN]Z�p�2X�\�T]�{-�����XDRN�t�y�%}�4�s���lR��8\7�>��6���HY��K��zU6GK��v�}αC3J�OM`�K�w<���h{R��-�hA7���,3A<w$t���|�)�ӌq�Y��������&������F���DUYy�V�C�aBD�����������}}u����*����2��"�02)�3u�����)k$�ĳ )j������׷��������믯��{.la��f��dl;eXAIf9yuFGS$m��V>�>�=���>�_^>����{e[d�Yf��9m��C�Bl��R%��ZT�&f4�DNMe�d���d�V�Q��&I�;���+j�̲:�p�t¡۫#a���mu�me�e�yl]]mRS�[m�fd��ә��lEnFFy�kU]K�Q�Yl��5��Ze���9�n�mf-Q0ѵ9	���A�Q�TfU��dd�[��n�\޵���ʄ��(�s��76�-���Ў���h:܈�� �7w'g+3,2f22K2��6�2���623�*L����܌��e��,�� ���P�aYQ��fP��~ �O�a4P��5��\�fZ���[�2��!�v�h��̫|)WL��m_7���]�Z�<�p������^��w����Fۦw���Q�f��@��4T]�X�P��ti��'~��jH�����1D7�[+�#U����}7�K v��Yp�� uE�i��� 9�c���ʑǱ�KצF��[KѮ��fȗg[5���4���뉴�Z������WF�p�ʌ��g�/��������3y��aܑҙV�80eH6�����z��m��g��9�"���5�f޻�(|Ǣv�cg�hj|4ͱ��ͣ�����$Ŏ�Z�D���x�J	@�^;����;{
�p�@�Lײ��[��!�Ǟ�?tڻ3��m_m4ìٚ�Ϙ6e�i�9ywZ�윩VЁ�}SWs绀ܪ@{���:�SJ����7��J/Q^s3B�FP�kh�ʬX�Am��P�WպZ4�ە$���:��k0�����R���'$r�T+�l�KS]�]�f��h�i[��_�>��d�ѩD>�"�Z>'��̕ǋ�2��2��o��)=1X��Q����$�!lևz�"�̿�>'��Ct	�oD�*��$�,��\cՊm[4�G]7��Q�zlV2u�]�Kͤ�,�E#L���dV��{�����^�R�H�~>M^	R�T�Ҭ��5ٕUPA��;d�3����-]�F&�9&�E�4:���ҭ@��aͭ6��"��rgv���N䙟��4^�o�5FS:<s��?xy���:���{�8��Q>���������~|N�s��`
���f*W`��W�lm���
�Un���`
��͐��!�����C��Pӷ�:M%3�������u&�ԓ�ũ��y�3��ZC�e�T���۵��\g�C�$}����O��g6J%�xª�z���)������gw|��f��^C�fn�Z�m��棼{3�n-a=2�k_A�"�KeR��Hq���$��|���P��`]����.=�蓇��,�ɰ�R��S��ګν]>mO6���3'��Ш�2+�n]	r���0��r�<�j���[ne
�ܭ��iށ���6�^w���aV����]/��*�$׽^0�:���Nf66>��)��]-8O��'���aߛ��nd])��Vv�HΨv�r�����a�g.���c\�(�}������d��;^��8���� �#
?�Q��l ������87���*ڼ򍲑�T��^�umA����|���4��
:'82�;�me� _���\�2�#l�:Ż�S�27nT���/[�d>*�v�|R��Zj̭��r�Rڡ�ճdO	sm/�^�1���F����M�咵�0a>�Q�����Tژ��	z̽�owϔ����i��-�P8�K�h�%_H��<��u�y���X����:�W��_�-�����[�8�B�(�"]0&,�����!�<l2�i'Rݷ��Ԣ{�����B[>�4�Á�l;[vP��ؓ��+v����۔.X����G%����u�:����=�O9���GnX��S��g���(����)%�Źh�d�'U�,�M�l��Ѯoo��[�~�"8���su7�q�u-I���G�5�ɭ��?J;�a̭2R��b�8���ܻ� �p���ww�FmI���k^�Z�V�SE�t<Ӓ�u�d��<��0��9��L��*Nds��㹋��vs�q�r�����R�F��w�Wu���zy�G���m������_vk+��N�%�v�g�܍d��7�U�:���@;)
��S�<=�y䋭��/\��V�����t�#�L�~v"��Y���7e�28�0���f�tP`�@�0�p�<E�3��
��3/ѹm����;�R�[��Ӹ'�)7ή��5��%�ʹD��h���s�=��׼��9U>͚�	W+{��(ؑ��=�����YHD�������3��<R��3H��<3R5!�)��l�^-�&�MZ٪���.۰�q �Q֤�pǱq���/�jKtJG+[4hyfk�?���M'o;��v��U���y4�&��e���f%G�2��sR8��<�g��Yӻ��5x�5ME�n�M�.����p��"n]�X����!�?�)0�=���b{���6��U���W�lc1�Ǣa�s><�i�9�bΉ��0���ϹӡKԘ�F�!e���;B�:a�]u8�<]w�岍�O@� ����)V�W��y����1�������'G������C;��;����%��cHJW2b��B�.N]�_����-f�fI�x��B�c��w{������恉l���n�-�U{B�q=����7]���Yzk]�\�[�=��wQ=lem{�maW;��o�r��;r�f��K3/+7c�z�z@�P)�D��Z��Q4���E�����_![NgRv���R�4f	nΘ}�t����1c�ʺfm�m�ii=�|t��	�;df�	�o0COy�tB��U��3��Q~�+) �;a:1t�9�g+��~a�!�ۋCcy+���zXlxz�2�d�k��d�|����^&�G�"ƙ�4��q��M�Da��B������|��{R\���F��P׾����4R�	p��v٩#8�d�mpu���t���v�o1�8�}�i�#�x�Z���y��Q})�\yݏA*bl���e�1#��;�!m\޶09C�v#��1�X�i#�E��̅��{x͔�	EXYZ��[�!���<�Rݭ�ܘ�帨�<~U�Wi,U6�L�#��,fuM�3�_srպ�����t�F4�<���A'�����(Fݍ%$� ��ǩ������e-I\��D��UR�i�Q�/�ve�r5-��MV�S>�Q�=� ܪC���K�>��L�wo��LN=�gvw�<�k�O�SFW@myT1c�G����]�!]Y�l�c��Z#./��\S���@��5ЖPJ=))��4���/X�5�N��>���7q��8s������Gd6�%~	R�Un,���q��.�׵Q��N��B-�ej��)��1�9,-�lg-�y�����ݩ%�Bx���ĺ��i�5�[и�F�� ����^��z�6$������)m��:�����zb�4�*�j6��I�w�+��u��+�ՆN���l���of1����G<u�:�]S눬K�<՛t�J�x�A��!���,��̣������k�hf��JӚIH*O����t������� ~X������l��(���L�߯�3�ή�w�9Ofͱ��ܜ��<F���<hT�.ŋ�
�IϷ32㽷j�FI$��u�^^j��Kji˦osL�g��@�m2Z� ��/��9�bya����Rr !p�3�� �L7r�u��Y",�n��'�Wt���c1��C(u[���y�:��~ah4�Cqً%�Â���K�ܷ�jRl;�����ɖ�ךdr����qb_�77�Τd1h���Ȫ� E�D��1R��%�s�����f L��H*�Ƌ۩�me����ƨ��~<[I��?f�#��7w3�As7�"N�8���-��+�*���fQ���@����k��9v�ux�w�*���X�y���}9���m�:Z�C_5ޚ������rh��wb�C��T�04b��SR+0q�4�pQY5.ۓ�n��F�A��sI��U�	�O2y+��ΪGj[Vd�Y�������xt^��:ConD@�*;��M�l��W!�h�{�ʾ�b�l��㽳Q��{8و5�x}��W��ɣKy]�����O���/�����S�є�t[v�zl��_.c��U�",�f��0��vɾ[z��v��R�'�V;��}�)�-`R�ԨnRT듪�Q$�L����{Q�\E�;mk��^g5��e�s\oP6��Quz�+��:\��;�v�j5��K��m���~���o5��񉰽��y�� ��ӈN���b@[}!��-�B~���ˣYU��BJg4��7���m��|���C�������'o3��vԞ��eC����YqԌX��뤒��a�����M�����꫚�fM~��+�&DAF��^�\��k��n����+�>��\�$EG-H��=�?����ײT>��*��L�"�GD�+�s����G{Z�8U�+�Y��͛�f*�s�wF��g�@m�^C��#��7�6q�?p���;$�����Tp������V��m��M/�Kܴ2+�ͮ~�E�i��^Z����eס�<�T�������:&_�s,��-�ק'�H3�X��i�G#2��S�l`G}��"�{��
6>R��G7��w����/:���S����4�9�C~�Q&)>=*����r�C<�9.�p�ʤ����KB���p�j�ҳ��Go�WG��)�9��=ʞJV�R����l�Zt ���K+�o)��Y��{�X�wKkh:�p��]ͽ�U-�N>Es�-��st�n��ܑ�����q�k�Q� v�3z}�W��y�Ԉ鉜H���197122�)"CT��r�����^�������RQ뎷�4=(��M��o��ṕo�>�]ݙP���/U֭������/xО�x�R�4���M���[�#\��qIqml�U|i�i�`k+v=3�@ye������p�ë$#�uyN^J�g���'p6�*{;�<�ǥu�9��l�^���h�m�ƨ�Щ*��UD�s�h���طS�=:�9��߷]+�OE�.����rY�Aݑ�� ��9��3ұ+|�N����sk�7�R�\Y�giI��7XG���w(�m#�5l"��(-}<����n��y�zJݬ$�i��3`�g���.2"9)R�B�s5]S8&���;;o8�Z�����Җ=�7�����`ho�C5� ��r���v��؂6ͻ����ٳ˫�牸�ꮺ��{C_.A�m��d��L(6�%5�A'6�9�3����hV��Y�U��i���*>�=v�:2����{v�����5}�m���}['�)s۶V���^���5k�IˑǛ'�f4�}��[�����V��=�����:��_��1�����}#�pO#l��U̹��_U�w�g�ve�ő/�<p�Uؾ�j�Ӽ�\���j���pvOl{�I�i���g�j�tV{ �×�T�i]Ӿ�?D������,od-Z6@�����e��s���k�z;�7�E�]�+{�;'��^�oy����s�:��g���!��+�ud�����)[����J�`U�s@N�,������V�-�EBd�w(���ym:Ƕ�j�aσ,���4�޿�J���ZW쌂��V��ܔ��3E��������U"]��W!��D�pQz��tk�[�w_4M��J�ӃC�2k9�k���\z���ȺSC�YZ�}��!������'I�`w4�rR��r�K{�%	�^�mRJ���E�
����i�4ﶴ��%\9L�Y5�α{qjU�z��gRuX�ƹQ΋�?����뻮�\�urݭ4�W��/��(�ۏ�@�v������ᛧ��5.���J4�(��<N�EԶg����)ف�]���[ݭ�*b/����w��ok{8���-'��j�
S�A
r$�s����d�[�jbٷtq`�M�m��*K�pb.�C��wfvڸ88'��
�<�mz�ZO3k6Y2ҳ�d���-����B��.���{Ϭtܦ-1��٠��BݼK6�e�|�UcI��Q��;��9�ڔv�0��lRaI٩{���s����i5p �Z��.�*%�'2�˹QV�ӊ-���2gX��!��"�^mT!�֥M�S yJm^�I�8�.7��)v���U�Pf\���]6����v�xml�gZg���wџ�wb��v�w�]0��y��l&a�2P��}�S�j�1L���6�˵g5sE�Aӱ�ҙ��I�ӧ]\溤B̸���/$�֒m\xA�q7�Xٓ����-�:�c�v�o��5�v�K b���9�D�U�K�w,V�ʕM��w��ø|�*t.�޲�k�r	[Fl��|��%A�M�׹*�L/1�e��|��T��\e��wWu�2qɱk�lUޚ�(/�P�WW]5��e����Sm+���ޱV�^�R:D�ʆ E�v�BI�n�&��wM�ɋ.��ڤ5�j�@��+KŹ�p�[����нV�n�f҃w!oo7.�u7A�}Nv9�.������d��Y�[�ztp�����"�V�E��5�����ш�5�h�����%�+9G��'u��/��<�buۻ8թ�o$��Kh�
.�ji1�v��Z�E�sH�4w�ީZ�!zi��Ʈ��{0�B���l'^��l�"#���m���uԶP�- � ����1�Q/s>xy��j��3�8/7���w4_^Dβau#���sr�F�"BT*�h����4�v]Y�M�H�.i�]�������e����i�iK�M������j<�[
�Z7�������g/��Ӿ��u�ѫ-��kjY��ۉ�DjL��Zڈù#��af��I�˓nA��u%���e��	6�k6�Wf�O�rP�tx�ҝ�d�|1yj*T��ɇ�R���V[�	}h�{��k�03c�[��]YR[kOi|��#y2�7JB��,�TtQ�۝DfR�/�����of��,���;�%.����&��W6.�����]���E�(>T7T=�nI�;E i�Ku����;Ir�-츖휉�!ۖ野�gmڛ���;�ϲ%����e�\�]|?s�_$	��(�HD(/3:����R,���α+7�*30�H���;z~�=���?_��?��___Y���((2ɠ'��2bt�ȶ�(7ܳ*222��������Jݰڳ1�2km���_^���ޟ__���>���9dPd��C�=��z�Ͷ3o4莬���� �00���&��^������_^>������fXV94��l�|�t��1�ɪ�"�r���0̘����ɋv���r32#J����M�3
rvȥ307p7s*2
���چ�,�
]�
�X�-ܴ2�̬7M��l��3��m���'��Sa73f�(�s76�m�����0�ͭ�bi�����u�c�y��FNw�n�rrں���7*�v�݊�L,�ksws6s7���6��Ȯ�.��(q��2i���2ɸ �a��0�I;'����i����fd幎YY�NA���&M%.��15M��VfV��h��FEn?n���z!�p��6���������H�q)F0�9�!$�/���>�"dA�%��:�i��R��c��P7مQ�i4t���ܵ[);��J����y۲��9�]��i�x$
�fß&$A��e��)#��H�E(��˂D�rP��'�AH�p��h1!���.H��iT������P�@�Q���L@�-��l�$�PI F�/���Nؐ��˯�d�1��RΨE��dKa�u� ��r���ü�|/����I&&(ɽ.��?b�׊����p��avދ�#-�hӫ�꽇ɷ9Gbv҅Ew,�N;�Yow��Ch�<�ƻ�W����ۍ�P�&����&c�1���ԯ��u>V^����Sc҇��5瞫�� !ggV뵚:�`�]d5�@d���7	���F��v	ꣶ���[k6�T�p�+U�
��#�0o]F#>��Ȱ,Ŭ�}ӽ/w1kh�^�<�����7z^:�=S��d8>���+�9� ��3rnƠo2K�i�'i�ܑg-{5�f�!��8:�zk9��o��ze���s>#�4�+���6����$�I.T�}���Lg<X���'�[22��G��Ƙi�|�j��,n�MR�E�x��V�_�9��/�g�f���YZV��{L���U���*���Q�J�Zr�~��N��>Y;�u<��2��O��Yj�];��t	T����{�2�XL��x���^u>�L�Ѯ͐�7���7#T�u���Uӳ�nV��=��ǰ-�Eʜ��f����=���vy>;^L�*�����p�^�>-`���W$�ڼ1��r.�shӵ�m;�����3*���]���0��YeazP��r�ӻ�M��9��<Uu�T+i̧R��(Hg��� [�R� ��]�+$��슅�='��[��{+�+&�-��2$������-v,z��>躉�q�tݙ��������-8ꮬ�θU����.=�-�|����h� \d
����eo[qHߺun�}ȃ#��ٵ��g�8E�"=��8�a����g�6%26��G]-�H�Ps�y)��K�<�i�q�3�e��gk�U�����3;VW����� �:��-n�Fl��雨u4u,j��{6 |�+��vG6���NZo�ٱ�xv��M�uor�o�:��Sv������p�?]r����Ā
>�ڸ��������R�v&9�GC�	1��֝�V۠Q�w`��S�e3y��wS7{��7�Ӱ�z4������4Ӗ����>b�Yum.�LU�͇`��j���g{�7�9aa�l]
|���o*�}_q�T{`���M�]f�\��Ӵ �-����>�^�4���Q2�2����l�2��s��
7Z�t��h���������'m&�a馞�|�ڹ��SN���D���mHۙ�CW�sՂ|U�K�UT�m�c�����٥�:����z�T���]�-6Kޤ2^�K��o�m�vt���v��ۼ�:)��7�K��*��Ԉ��IO�z��<��Rs��b�:s'MN;0lcJtX��~��29v��EU�泂�w_v�GJ����t1r�0���
����op��c��skp�޺����X���:$sC0h�~sз,R&�]}W7�lM[I��Z6��m�-l��"+6C�ٲ+�V#�c��Y�o�3.C*�w1E洲��Y��7���LA�^˦�+�����l�wW����m�5��ՂٌG}��B�0�?o��:/8�xm(*(�����`ά�V>�1�u���;z�+h!�h��W:N��֊׫kp3xӻX�ݸԙ\��n��Z[0S�\3g>�jI�����`�x����t7�R���##�꺾|�$�g��^�m?7�֯GK���j��8)�gi�u3=�ژ�,v����p���e��A�l�,�m�r�;Z�+���_�m.���!��93���=�/�Zղ͇����N�k�Ǜ\6������w����ʯi+(%�sK<|�@�� �����d��ȧ[��8�V�1�k��|<��9���[^���~�
��G����Ӳ�mZi��݄f]OH�-}!fz/fo�����R籪�u�U���[(4k2�e�虽2#1LX���a�.wS�g��X�$	ݾo�S�1��1�M��+�g���Wt�IO�n�n�:;�d�6����ݜn��y{�f�lg��RH�yG�d9��O�х\�k9�RհmSő���v�]�9F,R
�o�T^j���m�ji�[��.5��1��������g)r�1��J��,��6�)��� ����$��3U[tO#��c�SAm�Y x�/����GݮR`���0ҝ׊�-l�7��hԱn������ɠ-�������}��� ��9����Ӷ���ww`�<>�_$�TZ�ή�\�x�
���f�n�6in;�mMVz���f�����Q��8�]~W�>�n�E���6�m��[?G-$6�Up��i<�;�ᅆǍ���^�W^X�[E�޽�є�y�H����y{�ؑ��Z�J[>�K����oC���M{�s���jOW�5��5eI�r~���?���,�Y}͒��
��ۥ�3��n�6f��6��.�,��"�=[.�|��A5��8�EX�[���q$�}��+�[f��8��7�ݲӆĪO{�1�=5��{d��BB#��2�č�P��w,��կ=f�f������v�YO�����c�yO����L���P�������{����سn.x<��2&��8�-��w����"�� GY�M��=�����q	��&긹�����d��*=�A����XG�F"�a�#mc��;\��W �����}h_3F���iwKG-x�[�r<ajpsvi��d���¥Lt��u}a���4��vJ|�Z�໙��wl �@3���)t���i�z��M$�t]����2��k*�Żw����U��r��y��6x����v�Y�Pd���c�x�if3��7��nȅ�<`f�`�z��4��*Rө�l�*83��CI^��*Η����TU�����ܐ��d�l��RM�{=�z�NCɬ��Ƚ"�y?E>.�D�Ϫ����!p�v)e8�:�"69�V�yȴ���.2Yȩk�zv͙�ҫ�YR�%Uhq�2�z+n����D�*[�KD��gZ��3��"N0F@k��*�1���=K{9��RΥa�Ǧ�b0��jU߬i$bɛ��L�P�U���ZVӭ��3X��\ ֳ�ʹ��[,��c�t�TWuz�
�	-����imr̉v�5�W���ř�t;5nj�fq����&��r|عen�	l]x�*0wv_�V���Bu'��V�dNQ5�.�}j�\����#��xqK�F״�u�y��?6�X�[�#lq�+{PE��s+,��>��S�#���JF�k��YC��R�Y�Y/{Y[e����-����e[�Ģ�̇C��gm�	�7a�.L���(�8�9ȁR��T86!��p�7\�k��{λ��(�+;���gm1����a9���:���`RS7��	j[��M=N��|�����ߌA���}¾����a�n}�����#ìQ{����ܔ4��=�ݭ\�^��V#�q�/����;�>��k�#B'��������X�If���G/H��;Ǯ�N��s�eN���{��Z��������60��#Sd�q��ﯱ˽u�ۆ��N��� ѐ^C��n��om�m�m����e�3j��
T���9촂lGj��V�q�c�ŗ\(S�rw�k���^�����b�Z�oۀ+����q6��գ��>��E�'��T��%�2�9�p(���u�6 ��g�W*yh��8<Vء}:�4$��]L؍4{��!�~?&c�'j����Ӥ!.���Sbګ�c� �{G<��q��4�}�1��Z*��<|�ťĄ�I�^Ic�y!����P�F!]kc��W����mur��i�����Te�;SE�bSB��A�8r��$����˽����_1��*�A(l�[�v+�iYwJ�����9r,���x���yxD�'�L^�3�Fr0l�2���ﾬK'�ynS��~��Iu�;��-��[��*�V[����ٌ��22A�����I��Ov͹����[���v� ��[9��*���6�=�q9�M�/F�h����� ��5���A=�!śh��-�ʏJݿq(ܼ�ֆׁ6@�I吏�sxB��SP�n�@�ffc�>��4��<[D	�Cm���e�ٙgn��J��r���C�@wY"5oP�4�(.���3#�Wd�t�����ʁŞ%-�&}�Y$��`�X:D>�w+��(��]���,�fss��]�kԻ�ɽu ��ua#[^z�4q�8]��:{/�q/�Ú�Ȉ�����}�J�H��8:�7���}�����MU��ef3�u�P�^qfmr�)oY��9D��5�5Eu��`f�s�߸s`x�׉ƿ��y�̈
��E]����tu�=S�`ch��9F.�c�.�c�c�3`�D2�:N�w��R��k_m
�-��Qwk-�I�Ϻ�t�H���>Ж�/���ug��Gյy��"�N��Z�wN���BR���؞I��Q��sb�����Nf������A|ڄ�M������N�/�!(��	&"�3cp��4r�� :Mo�0��*l_E�=z-M�}�'�YzkM���8�i�u��l�\y��	������hi�0�!�3׽`�3v.PR��qS4 z�O�@l2�OV�}��A����i�u\B5>F4�ՠ����QӇ}�'m� RՍRz㹭�S����	�T���jU}`����('عM\�;@�E`-[jp�_6�<;���Q��*��*oL{:W�� �H>�VY�lC��8x6\�(��\���G�Zda����{h��d����K��̊ ]�:ww�+/�_����>���5쩀�3pW���y�]�Y'|��I�b�^�& 0�]=��M�J���.o�� �hoY���qM��'��ٛ.�eEjh|_�oZF�t�*��P`ى-=��^��%�>;Yڦ�m�-pk���sa]���OQ�\��jZM�&�ָ�@�X�p;��e-���%�kf�q�,	�v���m�7�]����Vpō	t�S�4�˺��ww*$�Am�u�J�	5-��q���^�����[���v�x���<���q����^�`���W�P�/O{w�k�z̰Z:��6����Y�@4J{#�y.�w�g`>t�mҳ�����m7*�+�y�E9SO�u�m�Mc�AF�l�+|8���Vb*�����}�a�;���i��[$9�C����X�#�#Qp�e�&뢃6����|Kf���Q���O=A��a��� ����S2�!aޝθW6��ہ��(k߸�x��<U!���a�K��3R�^����/����m�ϱ���p�[�i@�g��܏�������d��w2ݐ|������:�S����1�M^lE�O��
Ȭ�^y!�� �1yyb��4�ta���g�I+g0��6����A�U��%u��ڧ�#qn�c��L�c����cU�D�\��ϳ��mE6�9�w��M��+�[��ވ��>]��jp�al}M��G�:��\¦.�֢� @]�Lk�d4A�d�Ƭ]Z�PD�Ȩ)����H2�k��X�Il�.��o8KDp�ްF�KЛ\NŘr�\���U>�{��e�1�k���n��/1\^�z8�K�x������RFݹi<,�v���.�MB$�y��K���g�\�Vj���WOr�kJ���;.ȝw6�u]c�����i+��Ş��(l���3�e��ճ)e�_��P*�3�v�{�8�9@�d�n���}J���A-H��L��wvt6�V�u T��z	�஺>�I̽�
���/�����VR��e�IK,;y[�%��GQ�l9�M��˼�Ɔn��{x3 ��]ZeZ���və�I/����+��@�:-J�������wF�Ils	"A�ܻ'1Zp.[����L2r��w�������Use�;�-����0��n��ȹ�AQh|Mnq�!�P+�pԝb�38��j��øwV���%�Z*ͤ���e�l���rǋ�n;�*	0Ōc�yՙ���t��o**�����:� ��U�&���K������E=T�2�����b5W+L��G�7JfP��N��F�N���+4W4]%Xm�>4�jfLˠ��j�章����%YyQқ������Ap���P������b�[fژ6�D��nn�0u�2�7;-����/�Q+�V�%�@G��n��L{=4!��p��Ȉ2ym�.��\�~��u0��KUj)�Y홒�]sV�ipY-<䫋�v��]��1�n����d��88���}ݡW�u/����;b�aǹ�J���I����ҍgY�X�K��/k��z���.Z��A�'�o:��Ef���R�1V��ur�_n�:����V$.U��w�"�kVYݥ�M��gh]qf��0��Z?;ŵ�B�5��ڃQ.|�a��H�{&������pǑZw��͋>��{�nЩb�boB��a��{ /�U��#��k48�T�#S�w���O����ɣ�$R껲ԥ4:hŹQ���r��ڄW-z�3m�j�Ǵ�w[��YpYt[������[]�,e�f̚�jtu�I�lnN����X�eCn�a�pR����j��]bVdԻ{����,�\�iWL�z�FV�Pd�t��H��V]=��sj��0�1!��Ҋ�+����f��d�*t*nU�d,�{��Zצ�u�SӺ�����7Q��㹏��n�I�[r.j�͐ ʰGC ��
�稬W�u�7�2%���m�N�
�LK���%�C+1^
tf�Qx�lۦ;[�x�Ku����F5��V��rN�v@���Q<Wz!�u�e�آ�Z�6�V�+�r������j�'	�~����h�o�e[ގǐduiV��VfnfᙕM:��zz{{{{~?_���__\�0����q2
rh�"� �-�,�!�31hLs6L�����׷���������돯��bg���Ɍ�ldf��mfl陎de�VY.���==�������}g���¤��wp�\#w9=��d�'[���iddlV�{��ԙ���EY���`a;4�XbP�Vn�a���a�Q�%������t�lǸwL(6k-��ʈ�����$��$��,̧s�-3h��2>�=E�D�gV��<ӭ;��<�"*��':�w��&-2�����l2�sZ1 �c4�0�����
"6�rL���+,�+1p"hgK337M+6�-�3L<76�32̳�M�w��� ���w7t�*�2c3(��
�,�L1ª`��
"��R�f��7j���=�y6`�䓩�u�y����ǰ�����4���3n�?DZ��6o*,Lۧ�h�逇�D�fS<[U}�v��{��G�b�������U��p����4����ۈ�~굷�{y��j0�O�ି���+&�.�[�|�wfC^�ޛ����i�+_z/����=7���	�k���W��K�F��Gn۴1�MC)��Y��A��ɑ5H�U��w�]ohn2�Ί�^~����	+�Of#���P��� �bc�E�c�0�Fyq���Y;}Ѡu�Qi�����i�}�ˍ�wz�.TZ�����U�!oH�(��^T���C�[0��2�9J���Gv��Iƺ�f�|��j;Q��e�r�����޾�#�q�L;��k���؟)�i�G{���a���xعԤ�kL��%�6�ě�:�=�x�S����|�P�@����*�w����������
�X����yc�=��6 r��}mن�ݵ��,��w�wy�`"��t�7��9�
0��wFթ�jNu�lU�k�RtK��=n��yt�:p��k������i�7��*�ٝ.|�i����l�}h@�&Tw�Ή���ʾ�߮wO?;_c}�ME�#�u��gy>�X7�|��.�~�R��0b���{�� �2S�i�ˉ���{��OڛS>kY�QeTM��]�ޱ8"�,���z��mY[���;�J{`�lЍ4k2p4�jc������ ��p�4^V$�6�O�dr���j�n�^'�-�.�.块��fK64S����i�x�x;�r��-���&��Q�9s�*>�g�e���M��i����s/��oC�f2�R�u��5ҲR�V�ȥW�����q�4�O\T���C?�3VHr�E��ŧ�g�>=+L=�g�2e��4�M�_x�J�V��W�aAD9�d�u�ţ9%5e2r�t�֫�������s�ux�� ���ވ�����dƭ�����4�LwGmψ'f����D�cT��qV��p��!�j����w�F��ww���WdM��goJ`�L�]q���;���Qs���39��{q�Pz0�4��h��f�XᏫ-+;������˂{M镡
y��n���jٻ1��h���i@�[�:���wd�Π�	����
׊�ˡ���.z�a�l�.n��7I�?Ed6W��A��ιg�_v�9��֎;�/�Zղ��3	������̛���۾m[��μ�fbO��gt��������=�Rr8��.�i>�-=�kv�77�e���n��!���ra��>"l�ǭ�MOmB��j�{�Q�aS�C�&ծ5ؘ}�"�6/�Z�m�)��x�C'Dt�\�fh}RJ�]DE�̿dy�x�^�S���ѱʋ�M�t��&�O�-�V��zlG�M<mԁ�� 3� ��0��0PN��#�������D��3�b���� b�h=L�7��/�Z���a��|ˢ���z6�f�%d'�7�Ҫ/P��ye3��D��=��"������� ���Ƥ=�H<����WC1�7�]|qt��J�V����]3���r���x���>{��M\��r��"��gzR�n��{��ӗ��Z�8�w�ʏ�Z��5]m��^9wK���P�(��gd��5V��1$��fL���X��N�������\�#� �l�C�Z���><�2��=�r]!l#�d(e]�4�Vh׊Wf7��r-=.�]@���+R�O:S�_���Ϸ�/X��y�IV�ƕ.����-�Kj)�KS���n�M����t�!�v���U��&�'��r��Y��:�A��~����S�_�J�%�w�F�ޠ�*Մ���,�u�.L���v}�0C��|�]� ����h����g"�W)e�h?fqW~�0ד�3���6t�an[6ݟ�b`�P��/C)lm��K�e�J纁�2cuα;��n[,�M�C�vZǋ��&��y�CR�x�1�ov�.k�D�b����Ԯ�ij�^@��Co0=��f�6�j�QU�T""<:��������xº�����ToP}��?�[�=1�Ϡ,!��^c���e÷s�����o$d]m'�8bL��s#a���d�]��U�k���r9��ߣ;��߬f�m\�}9G�����>�ȗ���\:�25/�Ǜ^�U@�[[D;��K�P���e��,{Gl���ڻ���㗶�6Lbzȷ2b��!�M��f����e��0�6	�@������N^�D�q{!��:w+a����+��wNW��RW�sƟͿ5�ǣ=gR�OncW�H\�2­��uA�ǒ�1*n;����٭MwS�f&�EV£���rC-�m��E�"�0����m��*{e�޶z�gV(M]5s�*O�)U��q�u�ٛ�6���IS��%d�V�;��de��1��2!yn�%�72��+�*ӻ0�2�s��;fhUm�)*k�exIkZ�؆�"X[���a�R!y�H8�Y�v����K7��H���9fAݗ��)�L�1~�-�u�3o.���x�:�|��ť������[������0r��Y��p���i�ٵ��Ӄ��كryQꍁ[� V��u��7�v���pP����|7�Lù>�����G�(��2���,�S#o�9��dHw���|~��4S�/R)_��B�F�3��e{>�7���zg��j�:\\i_�s������^`e�R��%�{��ii2���sIYP�ōE�����Kj���۳�H�rjW�y��e�4�l�8-n������:�f`/(V^prT���.�Փ�;(\��TVv.�&����*r���E���/;ρ� ��_��E-ۯ#��Z������hv(�Z�ǫ+�i�Uf/)�}Q��e��YK9�T�q���~l2m��гW]z���;���i�mgh���,������3�r�e��������a�fJ�q���DMM��ohL�8�I����+��$m��9��/���ٻQk�Vox5Fuq�����l�Mϸx+�.*�����}l�?Uq��Sݡ�E�bЁ����S>�k0���t���9�z�y��{���"�j��Y����k��6�:�܆*�\1��d�7,�OP�ǟr��N��v���{1�(��q���j�-�x~a/�i�V(��R��Gέ�b�����<ܥ!�>�cY�m5��^�)R��$�������Gn�Xν�1S
I�i��8��yN{d,�X�_�n�Y~%"l-�ge� �F�N�l�ӵp�G���s�[����}r�Xp���ʆm�&i`��|�����=$��E��t���[�h����5D��{VCDn-�t<3�Jڹm���|���в`�;/�i�f\���G!kk�a���^lgc���I������/��������` �,�g;��pp��?��&�"F!��� H���wuO�Ϫ_g�e�rah��lr�L�cWt캺�0�ď� ���O�7����i�_����i��m7n��QSW����b�Q��� �WV��N���p7S���x��SDI-Λ��๮� ���~:��w$u���l�Yl��ʵP�x�����t�̊�!��T�|j��j�i��,*�-�fյd6�ҧ[���Wx�֚J���w5��Ee%�sHLyv/6e��0��3�6u=�3ܡ��$����^7�m \�����D���P���	��l�S�c��c�H�����εڼ��٘
�ؾ�j��X��B7�x4��j-�C�wfdÊ�R	��) �m�k-�}��쫤�c%to�4<E�?\)$��/9ms��/�&�N�gK=�J�*}1?:�Ե�=���j��ﷻ�.�F|�<b�:��4Ď�[�^�_1W>�WV�8�(�Y�&(��XhCpd� ���s�����zt��1�OYS��*p��iW����7hIj�[��S��]���4�^��˚�5r�� �]J�n�b�/��T��=�jj��Yu{TӖ���� lz���f��S��^4F�awo��:�_��>�0���Ъf�O6B}��P�mz�����a�;9d�K_vpq��}F�U=�$�W5Ǖ_ZuRۀj�,7�Ց�O�&����Z45�*E^Uf�(vǚ�u7�cM�H��@��Mfme���1�pˮ�>;=��3���PJ��׌��|/S�W�8��v�\s�0v�b6�M6��^!,��V�~J�qJ���=�[jl5��0��J�(��9[1���%\|[yv{\��V��$�k�y�w\��I��p�L=3w��Y�W�)\�t�	C`[���ȼ�\�̳_�l>dqW��F�����n�[���λ6؝��DAީ���3�[���y.�N��aa��5��{��N�L��9ش y��^������|��J�f<E�ʬ�q�cd�x�3�=l�r�wZ�r*�s�g^�*v�p}՜X�ʛ�ofjj��m�f8Wv|���쿱�K	:�f܆�e�c-�zq\���K��6U�Q������s�ӓib41�Y�
�bk��S���{d��ӼHz�W��yv�&��w�!�!��<���"�Vnq�I�xܷ�#�3���Q�8�}ӑ�����-����nq������~��g�_d6�ٶ9����^;�C���aa��4{uNȌ���	�f��!JFĊ���W���~���/���K�%��T<�J��f��_0�RD�����|`�&�랾�4f���B�x+E��͛<�s�9���f>7Mk�i�6�/��D�H��G#�y���&-�>����	fyM�H;L��B��9�V�>�#"�������[���2�[�w����	�|�b�(�T-^3��K'kVL�ջƦ]!���j�o�^�C[l���<2�> ��̓t5,�Q�hYU�]�z-��֡�WyѦ�'��^��޹��\z�i�_y���=iws:EIq���I���2�1���Z[g5��\�OL�����gywb����c/:N�I�^�����t6��<ۑ���Ց��6�_r�����WV,[ ����n�ɷ��ֱ7~n��]�ݻ}\�N�VT#�o�ٳ�3�2c��x0�	�Ū�����&�w����S���<�Y���p�/�nF����q5���gˬ7J�J�=��=��Ν;�����x�>�J8�d;�I[1^#:ǫ�W"���_²G����Q1����a�>b
N�r2�v�.�u��\�#���ά�1r����绤��vx�hNX�fv��e{>���33��l^] �9ϼ��(7twP8Ւ/��sվ�{Ff�jV��tl��׾�ڣ
�ױz���ƞ]��O,YϜ�Ɛb��w��[���*�6��[�H[���k憳6�i ����7^=u�<}͛螶m畁��4�S�d��l�#�4h�>|f>�B��i�����U���]&o[����<(���K��I����Ի��3������㌳��HUnܯ����a��W� ��6+���82{��hl1���Ϟ�W����o�������h� ��� �*?��i��@ +�*��١�� �O�Y�� ����
HH$���@����J$��4ʤ�@0L*HB����10! 0�
�'l���J0�*H�����@ �!  B(c��
�B�! �
+�(!  B�!*�B�!( B(H�� �H��
�膊�f(b(�j�b�*�n膢�f(`�!����!���H���@���H �
J ! �B(! �B�!�B!
�B�@ !�B!*!H�! ��#�!�	B! �� @�(B!C� B�@²��! ��!(��
HH$��H@$�
CL�M
HB$��HJ$� �)!"�)! ��1�CL�HB$����}����0�������"(��

$T��3����g���� o����w���=���P��?��� >��@�Z$��?�������0W��?�������U�^$�������?�)�;����؇�  
����A����3�_���6?���OC��C���t�N�����a_��AAp�@�*K �
� �B�0)J�"L�D�L
HJ$�A*�H$�"@H��$��#�@2°H0�0,��� @0�� ����,���2��,	 �0,! �,�(��0���	�# �H� ̋"0H2�,B1(�H*RL"
��RU� ��A �A �A�!ZZTJ �I�
Q&""(T��D�D���Q"(�p��X?��_����UTEF� J(�AV�����:���?g�����pt�������C�ߟ� U��x��?�~����������?ؘ��������~��  
���C����;��䈀*��W�~�����J��/_��ÿBD@~����J`ס9��Ӡ���Xg����ϯA���� U��C�Y��_�������x�?pW�?�:��h��������R ������`�@~���ρ����=C�R}OX~�5��,'�?����>��=O�BO���  
����g�?��)���O�x\������8����������AT_������<�AE��nG??��������1?�1AY&SY�y��_�rY��=�ݐ?���a�}BH�J�H�"�%D�J��)H(��$��H"R�Q	%J�*	DR
E�*%m�IB��B�*��)RR����� J*/�"HTJ��%B�J@��B�hҢ�
�o3��*PID!R��(���T��(��������R
�*�R���@��IU"�{�$�I!`  {����f��UU�EZV��[hC-AE[ZEb��@FfUm����*-��+�*�e"[j�S&�n���Q�ʒ$Un  �:(�B�P�pX
(P
P����5*r�[Ui�؊UF�Z��Xՙ�E6�j���ZX�V���0
j�f��U�$IH�  ˪	R��h�*k���*�2��FR��h��Z�eZB�M���5P4Jl�J�D���%  8�*�갤*Z�` [mD
*�i�)KTi$ �k+Z@41�j��-QR�*D�BB$U�  -�(a�@ؐ�R�Be�IEl��Fʕ�f��� ��"* �SR�V*AUUD�P� �   ۀ2��XB²�k4�F�&P6Db�mj��Xh
��*؆̖0T �R�H��T  8�s)��B��T�k  �� j0  �` �6K
 �� f hYU!(IJU*�*�� �  �  C  �d�  L�  U�  V  K� `��V  ��iUUB��RR�� C� � ��  Y� 	�  � 4c-C@���m ���@������)*K� � 
	�  ֶ�  Vh �` (@�  F� Z�  �0  ��� ;� J  �~@e)QP@ɦ0�	�� !��$�%I�4��2  "��m��G�h�   #A�JU$ �h 2b`  Ed& C#)�F�5=G����<ԂL�A1T���0Lh@4�d�p�8��
�$��k50�b+&��iBB����'������o>��c 7����c�<�� ;��En PC�@@����� �!���~a���K� �ê aP�����`�|�o�����)��� 6����ʵ.�����L�n*��c�qs%�A2n�q���$_�}m���
uw?߿����t?��z�����`Z����YӶ��c2S�67����m�@�{0*��"�,,��<f���hVL#F�mVڤ�p��t&��,2���aф]�;AL�t�v�C1��7C2�2����W�|6���30��v�\�i�P�k#V��R�+%����Gh�O.�Ub�QP�[����2S�iLC3Eږ<K&ӵ���nV�# !�BA� v�B:o�T�$m�22������*�Eh
���+1t�3(ZZ�O/��^�*��k�����Li^�[r1�#{���b
�0�V��v��A"@Ƕ�V�jލ8I:ǹ� Z��`�fP% �6C+i��U���M&���sq�!���d�kE�ʺ)�uyd-�ȺyS2Hۤ2#�1DU`�rTך����/3dC4�Ê�����/r
����I�f�"��.�u�fc*�hƆ�*7����C�aػG'w)s�mc�	�gK�Y�t�9(��ӽ�q2�:P���*��� VJe��T�Ǵ>ka i��u2��V+pZ��	��ۥ���ʶ��41M52�Ǎ�iͼ�d��ƣ�ڧA^X��
ə@A+Ubܰ��bì̠��QըR�� �/,�B�W,i0�f'$Y�9\7Ib��.���0!�:7]�7N��M���n�'K����b2q�ǁ��N^k0���A���ګ��Ѵ�ZQ����B��3C���aS�T�ź�&)�3�4��kj��	\���D�x�n|�X2-:F��y��a(D"h݈�`��h7v�S�n5kb-�F�St�*A,r��Gihј�^�5�IUǫ+Qxƌ/Y��e��B��-���*{�dhn�ܸ���oqIz�,_@-�'�53܋,�� ����.T����%��cI%6�o1�6B	PS@Њ� t�gtd`[!U���.�����Z]bܶ*9*<��2"*��.��I��l�Q��[2�mc�R�A�l��$�|v1n�8��;yt���ԙۚ�y��R�����yt�����M
ݗX���y�&���B?
q]�b��-�IX�c5TUt�	fBP}fҔ��(��-��4V=�f:^ S�QA`��٭c"z]��u�nV�QeLf�7%&��[�^֙aH0]��VF���CB;I���yt��Qڃ[��ڳ�H�zZF� ����[�������]K@WӧR������Ud0e���6�^H7o(5��3Y5u�V5�441L[�P�r��2\t"�X�w�'�L�.�����f�#�n�J9�0��0(���� *�0S�i��7L�<,��U��=Ӵ�<T�{ �܍B��w�q�X���͵�����E^TTrM�(ƱP92š�?��)��[[�Ť���
a�]��6�����%Y!:�h�U-�Td�	�o2ѭ+4op�QڛO@�h�fصf�SȢ�u��!&+l�6�r�ִ	7L��73F'Cq8>w7[���@��NR�E|f<���AܑaU��{%^:�QU�U�n�Db�1#Y�*�e`���4,�V�"��2G.F
E��]=մ�&T��&/0U�=Z��-�RU��48
�]�1�q�ɼx���d��M������'[���V5�
]jIԋC.;D:č�va����y�1�I�
X�T�n	�m�H�or��b�[B�v��+�m�)Kԉ�AO����tʘ$��d��f��襹��ժ�����kZde��Ð["��m$�47/m}li2*�m���� i��ңkhb�$�6A�EY�j��5��Tf�T��FɈ�i�^����
Z+AFhA��!���2��i�b���R��P2C{u�G��M߷�6��>����[f���(�r����Q9Ce^Zw��V�#kp �bI^Њ�ʌ^'�Ɉ�kł�vԨ��,�f4��V��n�2�;;�4�T�Qe=��vmRW{Yf��8"fTu��-�n9C�!��v2�:�*/ojL�H0�����,��,��M4ۧ�D�{)�sF��4�9��t�uf�{Ve�U��lܤX�RV+T��2�%iIf��(��Ϡ��m;��ڥWX,M�+ �v^�	1F�2�E��afhԑ�,XZ +,��e:jU�.�GR�M��d�Yl�4���7�1b���ze�$&��51X�3U0���[��R-:˷zB\x��"΢i���>�
��@>Vi�wH��.�����8m�
q
ko):(�0�yxvXo
)�*�m�D�bY��Uj�ɒƭO1�U�Ӓ/��;X�ڢ�C�#�-�q��ÖF�yj�e�hW���� V�tK/�P�7�1�Æ3��졏fG�n�0"Q���$�\D�3j�1���7$�^���ɋh�d�z�]!p[�{&��1F@M0(U�u��k*[����dbʽN��(�wq[v�(A�����6���˳��	1�)
84��^dB�$9N����Go&�N�ܻ���[��lLb��匙�y�Dn��juc��Ʈ�P���2��ܫ ���^̠4������(�MH_jV�A��q��7���ݨ��ۻ�k
��ʔ�l�Ԫe)Z��Aj�M�[eJf��٠�2J�D����Qͤ�v-��d5$O�iT�6K�Gdj'D���2n��q����U�������a膥�J郂T��X��|�J�J��ڑ�Q$������ �ʷ)`�w-�f�@EM�@K�!��t�f!�&+��Z�%�jV���
��(���1�.kbn�ZK�0�ݔ���[ �VC)���ɨ�p�A��Ƴq�N-��V�#&�.��bY�3��a^��g�ww����2�-A����A
E�y�em(\�Z�wn�cn�6�O&�)�Ѻū�ԣ�� n�Ц�!JQ�jȤ
1��xQxn�[����l���cs0�E�3]�j�m&�ō��5��Ek����]�sF��r� <��%E����]��8#8��˖E�L���*�Ř�位�6qôç�մ؊E�$�k�ڼR�mJڻJ��^��AJM� �f�ê$�;7�t��+N�b�]�!����Ҏ�N��h�5�hU�o�����*;r�N�:���-�,R����'ڨ��gd�� ���Xf&(�Z���U��&��X����M�;x��Df�W�����APP@^`Wr�V-9Xrͻ��z歫aT*���utkDZ�W��sV�z%�J��;4�X۱��tVm�F(Y95t��jX˛4��t�3%K�ڵ���@<�R�m���d�S7&JJ��5qf��������7r�f��ET��\���j�]*Vk6�8��7)t����(e�/�v�F�ŅU��ZK��!��t��@ �d�fҀ���OI��.^���CD�5I�B@@����ۂl�1h[��nXB���KD�hc�%kDӄ-�n�TiL����77> ��f�4�>ѣu�ől6�ͽD�n�V_���,���P'hm��'YRV�:Z�,�n��:hI-A�#p˫չV�ӇsY��Lk^P��2�����*��!z�L]izv�i��������e�����&�6ͥ���'����j��1�f#�A7KAZ&`�e촷tU(%�$�3oi�z���j�c#K]5�um�"����J3��`cѷ����%��ֱ��)����H�N�r麐�h�G�$��ұ�Z�V���n�qL�d˦l7u�E���r0�1@d�vݢ�mmmE��RH۲�A���3n�tTx��.��N�P*L�+F�q6�7��w-��Iϭ�HCt�H�Ҵ�
V�``E�t\���o-n�d� �1m�mcbb��ޒ^���ŗ@Dt��-�-�SAh9�v�[�{2��ET���#�u��u����kb��5�B'��cQV6��L�M�fl���ed�Ii=��������)� Ǖ4S02�yJ� \ݍ�x���,y��(�vf�MƦȍ�q-�ز�l�nJ(��5BV3x�)�oN���Sz*@�h5�I�P�J��r�5P�+�Q�n��>̭)b�H�);����j�-E�7d;$I�X9���*��+ƅ�kXV��6�E�I*7��:7wCL���v)��Y�fB�[u���V5cF!���ЬRDͥ�J�ki�����6�xN��*�ǚ��e[�Bm5���7�o\�F^�GIfQv
��n��T�^r�*e+'�ݳn>�a�i�fZ����>�^_ȸ@{���3l���73R�*QE�$1ye^����I�򡫶�x��:(�� ��?�
\�5�yvt�)VX�N��4G�-�6�d�GC 9uuI�p��m�fS� U�i3�)*�F�̬yR�j���X#�`1.�9-��3l�'%A�*�t\��^У(-P��#BZ�mf����9�6�@3H5�X0�jQ�c 	L�v+`��K*�`�r���4�L� �n�k�wF��&��
�IN�o�i@eYKՖSwl��"Z��C4�m8���V�n�i`ɟ.ć�t2��jW�2)��V�2��(�e�Ц]n�L��f�x������V���{s	-k��VC��5���Gk�;������f�Ĕ�Rw.�j* ��t�F����4�յ{��xvL}t�Po.��C9Q-��e��22f�QRf��X��YtY���j<R���髡�Rd��Q@�*�R3v��C!}��i檺0��Nn��4U�,P� �[6흔�R‌�&F��Ҭ'��K�:��%P*R�h3j�oV�Uf�Tf�76�(2j��40)����nnm	���i�BSZ܊ m���<Ր
��뽚��k>ӭ�p�қt!k�bn���f:Xr}&�l��Zr�f-7RbbA&^��w	��� ��GB�̧@|�lĨЇI���S�� `Uwvx%B7�m}�2�I�y���l�����t^�th�gn���&K�Y����է�,�]���yK��R�܍��Y.��l���j�6�T��7ND�Oi�osd��<Z6іn��m%/-dV�1�$J[��	��`�>�� ��į���@٩=N���9r�J���������­M;�n�*����� 7 �V��>�N��B�+n{�[.���{h��J��
uf�+ �K_�`,IZ��7��d��ば�$�㭇jť� P[ݦc�4i[ l�	�ug$�"�5x#5Sdݻ��R[6�	�{Wh|ooV �A;M%�����2����ssh����n��i�4�d�w�w���כ7H�w�[�y���v���P�z��w�ֳZ��	�j�=�b��CSTv�4���Q,���*�iՙsVEuOj&Z1�S8��e�w��l�@��N���v�4���]+�E*��@�[;��Z	bx���'S���f���t�2�SX1EMc\�e�:�5^�̧�̔�H暷�l�($��ub݃ee'�*zF�ʻƱI�VRTv�-�o,�B��!'��Vp[
}�F�>�����dc�!�9z�ڹ���۳I��C�D�.!�2=7"ܑ�VJ(�Aec�.�6�E��%V���,�Z0!�Uhf�cbBK�*Ѵj"��&jrXQ�R'Z0��w"�J���%ؔp:[�rU훺�[��{J�B�ғ�f�%N�
�lKF!WX�dm�JtB��o�֚1��Y�+l[�5R�z�]�y�L�%OA�m��\��j�?6J�؀�ab/���������'￉�7���p$��=��G��tw�����'�;�_�D�ǲ�h	vO�����+)+'Wjl1�M�9s��o)���{�hz�^:�]X�����cX�|�c�\�B7n��6n��{-�x�ȱv��z�P�bQT�1:Է�.�����6^a�k#����WO�0��zq	�C/gɽA�]C��w-:�Q6A4��F83� t��XD��쏠γ{K`�zl�fu[��gܻ^ �+t�?tb��
�G�C��Q��y��e����5����`�Nsd�{E�k�����:�e!�,�]i���T�,2�Vv�;�u��d��Yp�9n��h�\�s;�Or����D��{B��k������Z��T�q�ˉAu��cD��k�}Z{΅�7W�{�uy�roiԒ��8.�Z�c����VŻ���y;����s��Gب�Ź�G��˕�K��ї6	ss%�4>{Ъ�B�̻���#B£#�7�pQ�Nzgf��_\�NGw��˺��2�ԧ����,w�#.�Κ"�Ɉ�����{\�Q���/2���왩4�uZ��x���;Q͹@v,zlt���{����X1����� n��1��|y}�[�ˬ�WjQ��ַ5����o�Y(��}��g��hZ���U'+f������A�go�H��+}�,d�%čڗ�)j�쬐IP��K3���2���+	Q���6������`�k�{�(�La��tco��`�Zn�S97�j�$��թt����ۤ����4e1�2����u�ں��\Q������:������{[Ӭ@���%��%[��A;Bu���=��
�'{���.Ԥ��^��=f��`3�Q@NםN�z }�l9O/ˀ��z3ʔ�x�a'(2�]e南�o<51h��#��es���^n�96��˛�_,��	|�]8���)��	����,�=w
��Ȅ�1�
��ϫC��Ҿޢ�i�z��a��}��Wsvs��JwM�ƴ-��d3V�EW k����ƥ��L�Ffr̖r y�\�H�S�T��L��v�*R[0k掅c
w���t�Jh�����~[��qS�t�@CBb7g��zMra*�ݹ~\��=-/c�읺�Q)�ص�:���Uuu�EV��nYة9����˻y����r]��^΁8G'�]+����OFr��5��oS�7n�@�n�U�L�.�Z��`�<2��i�t��/���R��Y��Lb��^qzQ#����$z�Sμ�0�,��Z�Z��0�̥%�B�y3/��\j�du#P�t�u�ggE�f�"���]6�v��I\DWG����Yz��vy@�]��v��Y��\e5��Q�Z�����L�ԉ���)R�8�Y�էz.�f��[jq��b�>#Fә����Qq��s�^r���h'�ay��	Q�|���ݟ��@!t5 �����V��K6�ݴ�Nft�X�vu�.�4��G4|hB��yN��1�E��l���OD�u�H=�wG�����j�J���ur���D��@���Y�s�(�G�B�'EPK6���w$T�W��<�;WJ[�Ŕ�-Ĩ�|h��u���N�،g���U.;ɿJD�ve��!^Z��7��д�P�h�ju)&i*�J���D��o x³���vu��6���t�HH��G7��iɰ%����b(T:�i8�<�շfK룙��p}�΋�Z!h�S�;�w�:�r��mI�^-]l�-�٦u��Jf�@N��e*|(�7YA>��n\S9��sFP�mu�_mͨ5�vw���9��D7��Ǯ7.�SNJ��Q�ۨ6���xϯ;��,l��/���v��їi���olr���$���8����jNs(��-�WbA9����&��M�$sOg}G愻���7��r�ޫ�����B��o�T͹W.��9�1�]-��wkHnt����avP����D�A��Q��W]W���u�[c4��|9֋�m�w���u;5��\�-!N4l�e�ܖ�p�,�tL*�q�룖'D�êH'^�fVtK2��@��"���8^��ɖs �ǥvu4o;iˮ*'��t��W[٣��+C�՞}4a�:]��n+\A̝�,�cVb��vѡ1�ɷ��`�R�UJ���_-�1��i�E�4ã�=]��_ ���rv�;�j�Nd���:X�w������v`Ǒ�ҽ���IJ-��M+F�%]�����j��w�+��v��,�-��}��P\iG�nn�6냹�:�;�R�A����o�7���'W]u��N	X���s%��ۼ�4�0;��A�z�4�C��NZ��A>ù������N+5�Ұ�+��%9����������ٚZ���\���������t�gT:�2ڙq��ń�V��_	�u6,@)���L��)]�A 1����\��T�v;���&�lie��N��]�;5H떂��C!�\h˚�� 8��k��}�j՚��a����.��.�lD�P���f.�7	�>�^�h�w��P�`u��ahT��Տ#��C��+f+���\�iv�c�us��Z��t�6�#u1O>��������ٽ�K�L}Hĥa7e��OE�S���e���.���V[�]3b��ݺ��K��[���E�n�}������i�(��3�ǝ�����aj�P���` "��")]���Ԓ�����N�5B�,�Mo�q(�dm�M��3-��Ƨ,��-+U�8k��O�IQ�i���V���:�d�!M�[=���(L�-��p��w�W^�sw��mjW����d��P���u��Dc���z7�W�%�]�U���Mn�\�ԙ������w���aU�[$��O��vs�y�ME�9;�� _'ݨ��öf��YPۖ�h*���hl�{y�ik't��nhs�:��R�e^���HUcHl����r������|�e�Etu���;��,P�U��N
s{�|rKmp%^��������+�;�[�:����c�c��
l�8�
���7��I��:��g�P3X�Ҡ��e(+�;��6!٩e�9�5E �����j(���l�6rV�ư��כ-�JfI>�R8m4i�죸{����L3w�R�۰�����,.���E��y�b]b�SE��Pw�՝�)�߳:��.f]�Y�����-Sh]kġ,ዮE9u�Ub��ܭ�A쮕���Vz���M����lu)�gA�G�$	��e������hB�һ킹�zjNyE�IiwE�f��������,9϶f
{���3�ah�XR��jh�c�R�2�������p�4�,�i��5��j:�-�2�u$�=���u��ц�l����ۑq3�mH��{�����]����T�u�\�˚�3)��i��ͼ=��boX�zWv�>mo�����J��66��e��bV�ְZ�s
���3���'��νٗ�_q@]�"���B�9^�qh�Ր*�f��`��:�@�T+n�;\�Vٵ��{0�Ƶ���`�,>@K�N���U���^WJܛ�����(�ʇ��0I��I,�*\��������c��B&����tyA�o�Z���D�k�V��j�-�]��u��3��l;ĵ����y�O�M�����q���+���ڋ�V�e��gK�k_6�^X�svU���*U�-�X�֌�ue<�QuDn6�Jٵ����=��hT|gc1#��׹�"��^Ni2"xx�\A�CC3@Jgf��ɶ+j�/��;sy��C4�*��yxLx��vG8�{Z���Y�R���`<O.{���k���cu��>�C[�,q� ��׻�p��H�
|38E�"���D�Q����z#9���bSW�p�i��i�}�i�U�)m��j8m|�Vut,4���핐u	���DR�)��%�}���d��$ �ᦪ���v�Cjw5�ȵ��b�_mӶ\�8�wPWZ'�R��ڠޑH�y�����;r�{�t�wV������rWsvWT��=�2�y]5#u�R�N����\K�*Ta�B�X��x�1ǻ����en�v*�{r�@V7��v���Y�d��n����h)v��mu�%���V;�h�����_f���m��SX+	�B��Y�Q<3z�ۋ�jԷ80�-��c��d*��y���]}��+讧E����ͼ!��Z�J�ي�8Z�k��PKO��wk��{+��,9o�׋Ft�F�Њ����N�ԩ"1�������U��l��� �w�vz!˒�'6�y�����2;�����s�+���So�r�-R�:�yp�A�u�g*�-����q�Kxfbٳ�I|/�U����,NU�����k�q�3�/�ԉ��u���L:;�.�K'v�A�&#����+�Z��S�v�ʡ\�� ۭ��%Y���.�n�}���|��W"��T��Ӿ`��'���-��ĩW�v�ѕuԻ���/+0w�(��:�9��ݵ��$�������*Vaw7Wq��`gni�X�����✵�6՞Q�ьK����'\+6J8�|{ȗ7h���Xg���ٷ§�&���Ag`�t{oU��Z���E*է}�p�����em�nR����Y��S�Ötn@����܆�sh�aP���V.����[�ƹ�wX8�*{�5k6��7t���ǚj��wJ���j{�H�h�o^�[j鋳x�dC�ݙӬa���P4&Qa:�6�I��{��yN�ҭ��*��,˦Dk5x�k;O��찆�X���W&0���;S���&|.�9���iq����^ķ_����)ך���'����:��0h��ھ�N��9ptݼ�T���1h��XE���a\�|��Ȩم�[���/�}��뭫��Su�y�ٕ
�x��2^#d`��_J�;(�ɄNX�q���5����e��]M8�ы�$�h^d�d�n��:R(k/C����y��V'����<'��	8�LN'v����(�ύ�΍�P� ���D�]OpV9-�1W(��iGF��-.@�t � ���K����/5�d���U�p�}F�
� �k�^�-d(e���w�����z��/:���h�^4Nk���w@qP��Tw�4��|w��
�{���A�|��n�E��՛���m����e RF�X2�	��m�7w.�J���:�B}5˫Uo�w��!b������Y����X�t�f��gM�S)7�!q���{Sf�%p�D�5�������U��O�;n����� fU��8�B�E��']��Ӷ��wv�]�	�]p�E�!�T�N6�f,N�])Q,e	��[�����"ZYaF�ɖ
�犄{��|4���Q�s��S��#�n�"[}��ΐ��땳����m��Ѯ�mV��Ky�ɋfp���s�HR�����%���Ql������yܨL#@�*��MR+n��R�����*�eJ(,��zH]<K��ӕ���l�r��/��L�7b�X�<�t����ڰS9T��>l��Ds�+ye�t����sV*�ݰ�| )���g�j!ά��V
��gv9��oo�=܍i*���.^�AK-D���G{C�B��}��۱W�b�d<�ѯ��M�ɽ�}�+�d�]b�5u�Ń@�`��V��0���Ĳ�/۬�o����y!���oK�I�HV�p.���]�����#��AF�:
�'���65����X��n�H�:�	����Z�\�,���9֔�V�ղ����WS�Z.<�}���Y�����[�a仯��-;.S�̾�4����җ]s��gvet��H���ڸųVD��F��;o�.�*8�/����_��������?/Ӥ��  #�$�Ui�D-Z
�J�A��UEUPzN�E��g������i�To2�?�4��i7����/d�& .q�X��.7ǳjobx��=�]��7���cy��Nk���v�3.��"s��H<��V�V�v3�K��x9�7S2�,�Q���N����mv�1��o_+�s}z�G'��7�l����`�t��fґE<�%��/�������_1p�u�u��^�*�� ��Z����0���9���.�(�ʶ�,B�:�҇����L�A�R���m�e��u��j匾�b�rwÀ�#F�'�J#o+���x�N��є�t@=��/m�з�zo��X�uv�3�V]�k��F�jQN����u�p�q��ڛ��^Z.�]�$�(&�����KM7˸��V��n��.c���K����r�(��BC���lZ8l��K1Bn]N�ٙ)l�>J��ـ��1�������Tի+'Q�ޜҌ��(��T��w&����暛n�t�%�[W�u�"]٬E����+L�r�uu�ǻj�ddc�!Rn)Y��]>��}�M�c��T�1��|�)[�c�Vt�ީm�&Ȃ+/���8͢��oy]��\+;�&��=E���%��ۧ�(]��d2��v*%�zUm���o**�p�YI���C����;g��an��$٨q�V�|��e�<&
w�x���@�;��y�����J��(�j�(���L
�mF���ec���+3j��p��	@�6w�t���9��XL����i���o���yՊ�����Ʌ��Cݴ�9��5��0 �Z���j�%M9:hr�Ö��<�Gr��}��C�m�7V��{1G9Ӗ�������%����6���sn�fD��k_n�/,�pw�_%��j� �Yt�Y�ȗA�'��ͥ[v�u�6��Xn��ln1��Dm�L����q�a��q�iF�/��a=�vm㘜�;�!G�c��f�u;�����!�@��;���3�v�wKx-�\X���Ǵ��J5��J�*j�ۓcW��s�|��XغƗ����'F�%17�nڨr�wU�ռ�msH��>8�-��hT7�0檽������#�Sx��n�!+L7G7l7�1[�3�d�x4dO,j E�÷5�6���7��c?N��Kul��Ӌ9L���{�I��]RW��O&��p�����XM_�i�8��ɡ�pG��{ֈ3륵H��>����T鯳��wGQLmn�P�G���or����ʺ�d"�5\�a^ӧ�X<�"�,�]yR+Ƿd���e�5V;�m� ۇ����}PP�����la�
��u�%[Y7��l�; g�{��m�Kk�l����,�T����&�J�űX\��1ɻ��9��jKx�0B�\����A˧M�էp����66Gf��:��q�ko���}hr�F�=)��؇@ y�]p�����ܡb�n��g#��։�����ݭ&��+6I|+y�{�/�;v�Q�E���KOD��V��t���"tlf�L��1��T#;�����(u��y�-�]Jz�n_$w�Mg>��3u|�1��ۑV��)����wz�pD�7���O�Ncq�Z��ީ��@V�%u�*62��OkyR��p�se_X�-o�i y�����cRʷ:1�R�U����9[z��W����CbE׸l�]okq���,�)�jSwIF,���2T�ڻ>	�]K�fW��k��C����0���*�gt���Gx㣉���xb�Ï��U��
�"/.t�f��>�h�w�:P�=��K��72�o 
6��j�_3�G���k��W������9�c�1�tV��ygt��&�V�+ŝ}ԩ�9�FZ�,+ǗĻ��
W��)�y�l����M�ε��FU�Y�w+Q����M�V������
�yr��Ý �al�+��yR�`P�g�P�{Y�-*�G>��¨|��K��䄵+2���$U>2��	5��6�ښJ�ݭ�{\�$�#������Yv� �e�'V�C3+��B�rT�TT�4���s�W��Δ�Pu�EH�Uo�a��ᘍ�L@��T����DTh��#�a���\�o];f�F�� �JݧW��ꫴ�/{k+]���� �����WV۽�s��~�J��-��n
���Zd9�7�ԗh<��j�m�]R�.��}!���1R��o&.#���2�bS�I<-h�+)�SSٴ[?=��Up�XQH#.wSK����;'Kǒ��,��%rGH��\@�u+�������N�9�w*k/��u�t| �d�nv�.o-ƍ��۳tr!�ʺU����uOw���9s���h͚�����Է,�ԑ�͚�]�}7+u`B+�)-&nv��I�q���:���*K�̜F���,;֫�̢��S���^��K.p2��[kكu�%1�s�M����.W/:֢Nb5��/m��8M�n"9kr7A�jZ����P��1��b�>���%-�H$�i'�e��s�S&�m^��5W�K�����;A].�aa�J�ⷥ�}�⬒�C/6t	�3gu��列�N�z�ƈ�D��2�1$�^�J�˾}ˉ�`8RoE�[X���L�.��H��m�Yj���U�Q3�07��
�s/0iA�4���M�k��n!-$�*��j��a�k�1�d�
��cG w/i�s�<��Q̹�&\UIj�T��{j�����ޠ�m:N�uR.�)�DR�'��٫gR��q���1:҅n聩��z��Δg�t}[G�m�����Q�Up��U��١�nJ-�"�C��wv�x���a���Qj�'Y�W��j(��ye����CWZ(�( �]��`�3�tSD�wR��IN<��vuep�#G�gP�#�\@�V����.�N\���L�BZF�o�n��0�ɫ��r��6���e���zi�Mr�<�fT��1iF�k�*Zn=P��Om�ж�ڼ��Loe>=78R1�M���2a��;����q܋�jзS�e��nҭ5�-��R���!FX�ܻ$��.�
n��}W|�L87��Π�{r�q�\%ե�k���!T�(�f�m��Ã����������=���Ċ��s3�gJ��;�(r��)ȏp=�u����Gu(֚F��(�/2��a�i��^�i(
kɜ�w]�L;ֹl��n��:�Ѣ�������˻B}9�F�7V�L�O�ݠfVoc109��v�6�Yaw�k�ae�͠��8�n���_],钤5TG���X �D�P�̡L�K��2��W���fG&7�׽�7
��@̺�q�[��\h��%�:��u!�G�4�[gQj����f�j�k	�e��[� "�tZk_=y�'���\��Ϻ�n�]۹X��n��>qw=N���p���ފ�ik��bQ+�3/��K�&�a�9�;�A	��`T8w.����t8�d+@Nm�����^���W�q�Af�.�0�ۘ���E��v1čJ��
����Tn���ބ�L�CQr�6��z���k�t�:5\���X��K`��OU��+Cn-�v䢕��;����][���%�Ѹ3i�h$�t�ԛ�MH.�uq��j�V�s{i5o�0����hØ���pR׏�����ï8a�����:���@�r��0O�l.���)U9��m�C��� ]dZ�n	s`�����vm��[�C(�8�c�=�I�Α�"�
ʮ�!��K��ɜ Z�l@u=ᤉ.߅�p;]�{�͈Rwz�ur�:���R�RPn��xIĨ���$ �n�L[��L�\����$eD��]D]Όn�LfZ\�*y����L4�Qe�φ�.�S��1�b�� �u�g����8�ڶ("��x �뢙�Y�R��RY���JG[]��lja��Uܮ]����ԙV~�{ٿ
g��l[ Dٺ6p�[n�s+_9Pϝ��9t<����	\�Y�Bk�P�}�tN�t�Y�rU�Pl�rdб�i�����:���K�]{�v�������r����ѩ\'�}\U�h6H�5ˆغ�V]rrOڲ�a�z1ɀ�r��,��/;��'#�Yxq@��c��Z�z�t�R�(��6�s�>����Ys����\i>t��޶�ԇ���h
k��>��`�w*�	A�C�P�����q��e��.�*���#V<��(��v������/M
�}��&9S�A����f��|,��#u�X���mS�/z;��l&�l���n�7)>�)o[��I��+6�x8w[�����]pC\U�F7����u��3�Qvȫ]֤��Ջ�r�Ш����w7�MN�ƒ�Ы�c+�G����I��"�hq��n"jg�i�.��9l�s�^]5՗����d^i�b0����I�n:��:�����z�w���v�=�S�,*���j�U3��3:�igSt�`�Ԃ�g������L�]��m�J�]N��-�lU��6�v#q�{X^��;��ٍ������|�%�m2n:����!�,���K��d�!�������/2$�����κ*�ĺ�hWv� ��뼊'��4�
�F���N�����;��p��̓w��`Q�4˙Y���|���LV\�\����寪m��T�/���:�n���2k������+��zܼe*j����;����Ӱ+/oR�S��F)A�+9�m��jΝ���N��|%�3,�N�m*�:t��f!Ǣ̈_dWH^�����{J�ͻgpee��7�zȬ��H�K��4A���L� ����7���`�iMՇM���ҘSkAT܂u������3.=W�Fh������s�Ӻ�MZ���e�=�Jp�8԰��:�K�+�|�M�G;r�뜂�z%�+$�^��ߌ�k$�r�x�*u��8��Z뀻8��Q�h�G<ɝu;�w2���%Yl]�w���s�|6��/ks#ke(>�Eg�1�ӲgW]x�l��e������+HڇTĪwt�=W�2���ev�!ܴ���w�9]i��֪�b}n��˪ŚDֵ��{�A5Wb��Q�3��[�ѫT�v�MY.uJG*_<H��PLa�*��8�2����]�����}��S#�:��2EG�5h�WlS]s�@�~���M�r���ذ�˯WcTĦ��c�nV�1�����Q�AԳ�����k�[��P������;��J֣l��ÒM�u�Q]��C�Z�>����wn�n�m)k����7J�Zj���ر*9�t�6��=�{z�F�:T��R��;����oP��8v�\��-<K(�n�`�����ʉL1G�<�J؈�붻7���d���b����a�P��*I�c�z
��@��Y�E����;qt/C�AoC��'�ݼ�9�^9�v�c@d��t��#�@	��yS*���ϵmp��gi^�̑�	��I`�
!�����,Ѻw��80>
�@�8u�@��R+n��۷�:��J�f�0�cc���]Y��M��*M��u�戩�_
�N���Š9�Efά�VX�ذ�h��v�z
}���K8I�K]H����.��cwg��6N8��ᶙ{:��S8�7�i�wrE��e�%�����Mb+�k	mp�ۊ�,��[�s�`��wZy�,�\済��o4}�z�����z��,��`+;��$��B(y���Z�"�%\;|�����]옂t�tʇ�>�o�GI�j�;xbv���]�gq��j�)���F�*��x����q�� e�9����ɕ��c�o*7�^B���m�����;��F�@�����V,x//�������n�1ւ���A�G��p���|�6��ϯ~���y�/�T����ҡ�v�AS�?������"fQu{M|�]�'�h=@:��p�Ye1j'B������M�,��-ܢ�)b��i�L�̧�,��d9�|Žq AW%�V.n���(EK�E�:�,[�{$wZ{&�(��y�/}�o"���,_���E_KR���L�竜obv_5|J_> ��d'L�9OD����eiGAI܈�Ќ���p���el��-Z�/+�=��!���^,��Mk����8��!WY����#��㛫h��� l�K�B>�e�CZռ�����p>*�c�M��b�"9�����[��Hfڈ�x5f�K��eڥ�ʢo����:S�������T���L1�d��'��ۥm���fՊKo0 Q�ň{���$�byJ�Ca}ܽ���uq�qZ�X�kGp�9Z*�c|:��8��v;.%���I�������QۖPY��c���gE�Ԝ�j���%����=��8�����i�Vb�	�V��9��w���vCX:����:oV<���������.s�=��7��[۩�o:~� �4($�v�G����
�N	^�y�s@�*�ҍ*�9T�YN�eQz&�H�q�9z�I�N�r�x	h�s�)�'#!�r7B�N�u(�9E'����.���ۻ�:ЏP'[�����*��x�g='w"$�=�$	P�'F�"Ȏ�ZPD���rS&DE���	0�+������b�DVZmڅ(3r����Ov��#�/Yc�TN�9���듳%��/9G��D���EGp��r]�J�CCR<�R�Z�^d�J�����B�'j��JIqл�N�8JF�Њ�t"�%g��r=�ss�w]�g�wt��K���3^�s��t�I��#U׬������})�ǟ��oc�"D`��l7��M�gR������vWT�/��{��֊�T�v/fD+�W�z�%�pU_�\����a�.���O��^J
�T�
��p*&�W؟m��Q����{�&x �T�ֺ�(�X��7U�O���{��b�]�=/7F�:Փth�\1����@|g��C�{���[����5Y�����JfG�`j r�rU�y�G���`i��؟�y����YB �P��%��q�u{��Smgʪбl�3YL	��p��A�8�К�YlC@��p��I��]��n�f08è����=(�@�yL�U�~�1��ؑX��OUFR�I�Ѹ36�V�z���L�Z�C>���*��@Lq�Z6>�X�Z�{����T�H�yf��޶t��x0�xc�o��OP�Əg�=�E�+u����W2�*#����Je�'�#�
�h v�z��̿�Ey�@J��Z$!��x��k�ڼ�ੂ���ơHԛW�y��p��]Y<k4��U��_�U��J�+-��T2CR9���^	T,V���w���Z�t�����6]]�ZV�1��΃+);�-��m�8!s�V��G^�Z�O_d,:{%hzH\����Ƨp7�b��*�
6��@��Vl���Դ��cВ�uk�Q`�c|r�q�;\�g��yJ%Q���7�D�+�P[V�KU�%�s �-��4X�ܟ�/e#��@n��lO�s��ҳ�2��y�O�D�v�]�O�k:��GV4:\����HaeN�vrv;�5�o�Yt��p���E}5����|%Q;����2��s5�o;��UϚEbH�t�?DE�G�|Ϗh�F�|uA�G0�=���@���U���U����A�]���^@k���T�T@���ie��KG�'��¦"|P��-ň/X��t*Dt�1H���T��(�\�(Ǝ30�ɔV�(�������h��Z���SƕY������:u�@R�U�qS g�<)�c^6F��▷�w,�~�7F6�,8�=O��a�&��[s"0�)�����]���H~�gNJX�����LH{�Ǡ,Ƴ,f��1 �B��nPݵ�� `��9���L�:�2�|�237CXeh�����\�c�g�Ƈ3K������4�'b�6ݓǏpOa1��@j��M�]D�\es�U���w�e�E�(��Ի:ż�z�JcV(��r	�y�3x�}Ba!�4F�s$n��2��%Ѭ1˳�.\Z�6�4���ƿD�绋\��5Z/�Nt��j��De����	T��vzU��_j�}�w�7e{�}��?H�҂�YǄ�SJ�_*�ڳ>�V)�6�[��I�)&��U�7V�;a��}V����A}v�>utps��x��Q��܏�dLp�����;�&�3����5�i�U��U���4<5�T;f+���mU�(;��P:��}ȜЦ7��a�D�dk�P+u��r�`ϝ�fS�&u�5�[wV�;&���o{r�3�YP %:J D�O�Oq�5<ʼ��.��,Q�*r]�5�W#+8ΣaŻW�A
�I	�ͩ�$���8Ռɞ�Ӯ��ry�K}���[���O*,�+��vɋPa�0amu{��[��ob�'~���1B89J�2qj�<�K�*�u�\��'�@��� ;�`׼r��x�L��G�k`��o#`���Iz�2��Y�v2�8u���f��e��y�r�ZW"-����3z��-���"!U��T9���Lڝ:�<�1=;�i�U�N�rx��?����Hf�zETk¸*�'�A�@���0�����e��WM�#:���ǜe�o�Q�h��^^�|,=a|�1' s�=���O��֛3k����p1�@�e��l<7۵
�i�� ل��J���jݼ�-B4SUQ5��~�3
����^�����J&���S���3�;��ja8�9�	܏���Q�o�{Q&�u�t��qxGG6��N.����Y֔�����7X
bit���'��J4>� ]$�Θ�a����)���(�N摊�b�����h{'���¦�1�[��ne�0Zzc�������`�pM1Z�J�Ōg��J�ʳ�\���l��on�/W���������`�&%��}B��C��D���߮e�b_��3�������Y9�I!L�Kw���ވ���y��|V���<j����n���s_��u3�9sr_Qpv뿞9���8�$�L��HҮ�lh�D�4r�G\�9CEO>�F���-�ƥy[3��Sb�[)���k&f��ע�γ9�z����f��}Is��m��gu����c�8��$o�qz; jLuǷܹ�T��ԳX2�:"aO;c��Ea"8(= v\UHeJ �U8SˮT1a�Bv4Ce�1�N��1�҂���-���rP
E}�V���	��cqf��<K������W_mh訆�OM�:w3pԢc�n�uR��������\�e�Fc���������UonDW�X��X�h���uK��.J� ?��9��S�@�/�En:~5�$���.�^�̀�6�r�{���b��������DS�� �����X���Ѻ��>MXʝ�+I�9����6͛�H	�k�aWyx��l~HRƾۋ�+��%O�n��m���L˲�����0��G*���BZ��/��ë��3��=X��E�"��(�����c ���\�@�Ʋ؋���p����7��;pe6�DX��4W�V�,`�5P���4��)�p������:����kA5¬���إB�Y�7kl������1����6��ѺV[�Jgu4��������t�h�)n�6��*���<�g=�چMSr�4�N�Md,;S&wWi����A��e⌥��p�3�t�SX)��r0�?H�B;-�ٱ�u�F��t�,==Nz�V'�n��x��W�X�R��W������a�uL��V�ɚ�/�z�i���ҷ�;gh�X�6a�g�E��jʞ7d+�hp;t�3λ*�>;�(jd��Ǿ�N�|d*�8�x�uL!�pō�:�϶@\Z:+]%�r�v�~괭\������ĳT�+�|�;�.phwb}�w�f�p��b��}�v�)s) �.�ZU�j� ����S*U応8;�qv�yw+��7[8����h!|/�=>�r��Dp��t���t5��ՍӰΆ�¡nF�B�
��T�t�ǨG����b"��jS(#�|%Q;��?p�ڮ;�M�{pu������s+�Y�1��˒t�X�0b`���N	;zY��8�h�����GB��O��d��-�&�:���6� ~Zxԡ@��@bK�Ҏd�׻w�N:�U�����}�J��m�������a�V;ӗ�)��9�3/�z�G:˥�
BU�F�P/D��]���Υ:����v)9�΀�\ ��K��tj���ђ����_$�貭��y�ҹ�?8n{N�����
�:]C�gcz��x�}@T|�\���1�Ӈ������ZՋ�;\eF_\��hE�0 ��%
��2gڦp�`U٘U����o�t_��'�T��*�{�X�O�ha�针E�ͫ�Q�]�\y�ާ2�C����b��o�l�BÌ��s*"�gf�k�Y�������3t��}�X�H�sSR4�CH��l�V�Vʵ�_�j���]��늀��{V+����b��b��?h��n��j�lD]��r��#�:����.���'d�gRWqW�P�����PU�<xASOq�T�ՙ��Vq����n��<���FW4�tS���®g8�+�Q�x�����w��s���)l�r�g����z�;���֝]!�O��� ��4�pq*�J����٫�Z;'P��a�f���)�-�Xky�@���@���[�*�����檰ӗ�GV.�w��7a�y��5.�PU�|.|���:�ݺRH��m��789�VS�5�@�Z@W��޽
g��.X�f���F��8�Ĳ�Y��N�sW*�՗ҭ��ݠ��8*�1����9N��J�<�@V����)J���3�,K��&q&i�Vk���r����@��L� R�>�	^nOB�%��������+�D�f�x�Ȼq8-�To��A
0���Gd�d��㯦��G;�`��9��v�\�1L��ȖWc�"���#R��Wh�J;ՋF.��f/m�������f���懰��L�?>�����*r~D
ϗ���ƣŇ=��vYd�s�HeeD���b�����r9��$0�*9�ѹ@V��ݫ��� ,B`8�O���.nMDqB�c�ߠk0����*�s���X��q��lh�SR�\A��څ�,v���&C�0�j��5�3��ka�oV�t�G��'U
�vS�🲗��]}���쫯n܇���y�M]�hD8��q��s%�{?O���J�d� `��R�]�1������vzٻ��xV�:F��‘Sk��	��^�'j�j�9�+޶���A�71{7���Ӊ��)��@��;��ۭ�{��G���;CP��bN��Z��+��Ir?�3���q�וoXu"��󡎸��3۽١mΌ-��vPZ���B�`�{��vi�MU���ɯ�
��0��w[zܮ�Y54
2JmY��(Q1B2��������l1	J��������½���ȹY���j�]W�xk�gϢ�(#�~��1�H�6KΏ����m.�<x-#�[�\=���B+� ߊ�3T�x�Q�f���ʕ�u�`ִ��q�] ��5��:_C^�Z+�y�<�[]Wb"�3���jcr+�g	���9����E��dF��1ou ������K������ˀ�Z��M�甸W��E9� $x~}sW?h�����Qqf�D�� �v�$�=e��O@���.��/U}#Oi���x*�;�(���#*���y=��g4�;r�sB#�.;�����b��F���3*����O�w[�WE�(F� ��<�*�z �@���@j�����>pi�l?\���U�a��k��^U�n<��{-N��<�ݒ��@��x,879åJ�CW=���.3k�R���zV����͞�z�lh[��*41�v���Tk˵ʤ���r�v;f���c�|t�Y�i�l���L�3�j:���3��d�v�Hz��S<�7	Hʒ�ld	jY9u���$Em�ݢ�j)Ol�֤��m�jt#3���U���'��ʩ�'�������P��SJӗ�.�P��"��q�,��@NӸa��r��.�#6-:�6C~������AV�u��Ѣ��XP���4�����bT�^�rdr�wF�!6�{��p��,�?!)�+g�3� _�W�]g *3t7AM�@HWu����n�,�]�>�H�@�v�&-mf|kE�:�����x�7�m_w�����l�+G�/�K��Z0O������,h9�L������s���s��4cN4paV��N�����W>�t8��0�����b��F�'���At��w����y�ߝ�����¨9��ϊt�O8[=�w����	�������Lx ����kE1§�yo�1w�� /h������Ǐ�����e�	����߫�y��pX
����(�95��F�>���ʖq�s/�q7B�8���q�˶��X1��oU�
p��j��COl�!]]�m��\��0�9�9b������}���lu��uf��e��L������Z8M|�l�V�2�]��t����W.n�mv]��m�E��Ă̪�45w�K��G�v1�51F�ݵ����A�<	��"Y\�D�wt�J���6��g0s�ʽ�VoH�;��D���><��^Qnjw��M\�ȧ`��gc*A�A�n���W.��2�Y�V*�y��"]%�9 �����^�u,N=wWv������ ����t=�LtEL0r�R��r��'ݔW��a��Vi��e���f��a;�"�:`�ܕ�:᫴�ẁ3�n�	��3-�M�N����N���o0���"�O��t+���J�37��l�7AxQ뤕i }��˫5ڠ��WgìlD-�G��M���|�Y׽�W�4(>f�XT�ޘ:���Nk��+3]a�i\ڹ��l`/*�a$P�+X��U��P����d��L�t�]w�X�c�Vr?\�����ufV��tqS�Ej��;z�(�xE���L����p^�}�tq�fih��5Q,��g�������>陃4�F�9�錋 Oǣ�4�+����F�6�bk�p���m%��{)�ʇ��L_g>�j�����3T���,�݁+��wut]رdl0񸶸����y�2���C8Vq�j��O��;���u�E����rJ]�����y{��"ק�ZqW�D7~��!�IM�#���'~�g.�7���5^IƔ�8=/6�ku�8D7,�#���n��t��j	L��C:���"1S��vU1��X�PX3"4��L틇\���J��Z��h9Ҋ����Z��^pr݌�N|gtj���U� ỵ���\y�Dp�|z�^%�{:�>gx�d��Ih���G�+\��t�^kQ�=��M�Y�N�O�qY��n-�����vA�:ヰ��:8̓-�w\�cw�+���r�|��	��&B�Kp��e�Eh�6-ݧRVkz���m.�������.
u��j�:��(B����F�Jh��b�Ѵ�Gvtdک6 n�`��7��8�W.�]gj����!��^��XN)�̶5Ϋr^�^lV];A�+�xH�>��Z�T�4�%2��=��V2�o��[�A���S��QH�����϶�Vkvٓk�e��>����]L$�[bv�VE�K#NZ��9K�?h� @ �҂4��5UP��Yyr���\1.�)���$�E�)Q*KԌ�<Ȋ���-ww/'L<���9��vE�����R�U�˧.��y\��s��6��Jmi$Z9��+κ��L�OEWP�Ty�ԗt�I'�DQ�����K\�DTQ��K�*�-uĜ��
4�
'Bs²����xz�%t\+.�拺;���9;��z��\�B��qw6Vd��L�Hz��w�����ܨ�+es̫Ԩ�Y�8��T�`��S�ˑ���9*r(�s��$�3&��UW-wM\wr�.#��C����Y�N�NȪ�E�wq۫���%h�\�S����:w�}��������<:�����t��OWIv��7���b���Eqp�R����/���Ͼ�����0�ۏ)���|l��aT�z��}~;�y:}�,�����1��N����)�>�r���M��=pxL?,!��yW{M |B"����!���in���iy��)��r�����_ݤސ���y�����xv����>1���aw��v<';J����q�<��כ>���P>��Bw�>;�ǫ�
�c��ru.�lg���B%ﾡ",G��ǈ�����nv�u�<&����&�|�ޓ�;J�����yM�N<�|x�?|X9	�~~��C�s��z�˷&V��ʸ��<z�O�k��߽�u�q����%~�>�#��$zO�7�oo;���ߐ�UǑ=�&��࿮��9���m�<;N���~�^�0�~��+�4�w��9L/����.M���A˻�:��Ȭ�ў������:v��e<�zy\������㏨s�����������0��?#��o.���������-�����������ﾼyw�xC�� ��7��好�6�"�>�"?�_�zO_-�]�4���O^8>�������=&��v97�'󷟑���C�k���ˉ��L.�~�䝥M���
�_�<�~���tTd��w%Ĉ� #������C��7;�]ɼ�&M�<�����_��9߽�r�����s�r�\~q}�� I�!'��8���!?/~�������������˾}���99�����]��L>~���Ǖp.�|�!��ǟ�x<��><��=?��]�7��n?!Ʌ]��I�7�$ސ��?!�{|!�A|G�B�R�����7�yy_����
[���SI���ݼ���y`��@��x?�}��ߝ�\I;<��߼q�7!>ݾ'=���}M>��ݏ?��0������˹���C��y#6��JO�R��>�#�7?��>�Cߓ���$���;˿!�?nL*��<=�~C�a|!�w�^1��i�o?~w��&���v�a��������ۓ}Bw����[n*��V(��'V��� �:-�[��tk.�ە�:{4NN��1��ǜ)Z�V�jt�:�rֈl�;��ZOV&�v�����R��w%m4O`�DV��q��e�˻�6�qD�J�M����:�o��C\q�MNn�5wظ,���C�Dz��xL/��?;xI�Wx�mɅ��׸��S <��?' }I��݁w�>;�����av��܇'�9��?���Ă���nD��~�����z���{�����~7�M?�Ƀ��l|M����M�������?��[���oQ��8=����x�?�|v��{vޓz��i�c�7�o�y���}C��?|Ro�H)�÷�s���{<��ԝ�x����7&�z�����q��90���������ļ�q����F��}����v����Z�j�V��>&��v����~OcSO��{���0���9۝&��90������)����q�>'�<�I!�z������;z�nL.?�^=��0�w��?]Vx�k��R���H�#�>�G�����~'�g��=&?�_�y�c�o�N�>x��o=��rS�w�����I����}`���w����90��(s�8�����y���_�z����������������C۹?~��ov��{Ohs�����q ���7z=���{BO'�޼}v��]�=~�����y����8��l�SH!��#�,���}����ܩ�8�{��k�>��NSxB��O���xC��!�?��<&|C�x���o�N'�=���	<���xy��s�_��< rN߾����_	�0����Ӽ!�4�#��������M���@���Ǆ�Ǿ<"����g�ݼ<��M���q�}����pN	�n߾G����8�����;��~�� G�{�~�@"#��\>����^�3^��xM�HI�ݴ����X����x�o	�$���|Cۏ*�]����?&�I�?�Ǆ�$F$�P�G�~v�����Nӿ8��|&���b��N^��K�#�>��#�n�������9<�w�����'o!ׄ�]�N��0�����xC�xC�y?X��������$�P9ʠ#����h�W����2L�����%�-#{�|������õʷ׌��31�Y�Yz�v�S+2���?bx�{����b��������Ԓ�G[�՚K;�[�E��o�Uz�~o~�|����<���&��q8���x�ĘP�����n��<:v���7Q�\~�&���`�\�pNL�O�=���]��{�������i }��">����i��~��\�c��E����c��́\~B�uP�eE(?T��$G
�U���Y=j��Ϋ��x"kLA��P��2��K,D_*�-��~�@�cnM�Y�`t]��$�wE8��
�P�89Ѐ��/eۘ��[����4�wK@�K�J�$�FX���o�Zi�SƸe��1ױ� �"�L#Cfȅ������v��X��5���D�ҭ��3��υkąG/�o�d�ݙ��M�w/:?z�[�@��	؇r����_QW�[	>⊦�)��M{�\[�ފ��֣��k�+����}
��Hp���r�&������Z����d�T���4�[��|!�p���"ݖ�E��/�-F;Iȗu�U�!GFB��a��(E����P��f24W:�#��K
���7C��Y}r����V�n��X���f{*�շ����B!���.�ġH`�v���_�U�9�9��\�I�j<�m}���s}����ۼ1�8��{��K&���l�v�����hK�qgP�q��_Ͼ���w�u�����O�[��D�~��CWt��i�6x\}4VQp�=��ia�pP�|���P�Gt��%(��8&s,Ch���E2[��O�8�N���J�e�*�g��P� _VQ��-ʊ�a�1��xU�9���q�Mh�|� ��y\�]~hE
�����pc���b��+:�ҡ\tm����ÝUB�����X��NOKD��U9|�������g�&1��i�t���0���)��ULU�����
��F*���mw���&��ר��ԅU3
�<
�u�Ҽ'%T��� �:{.r�����ՈO@��V)G^����@�u
�J���f�5+�o�nα�3���o:�!:�2��B�^Cϒ���s͊��U�X~P��:U��y+S4d%!Y��߶�-5U۴�ţ��Ϗ�(�:�u�I㞩�r�m*������劻�7��,��_v�t����W�J���F�՚�)�S����+~��~����os:�>��C]�r�C��@�Ƴ�;����P�Kx�W�xS}�1{z��l�����I�*o�
�.��,5ß/���P]�k�@hd���n���FpV��{t�k��O&G���s`���k�X�hx]�������Q��؇�=5k��gWE/%�*jA�H=h
�Y�Ϩ�{Uk�@�8ooWԑ����qܜ�|��G8���Q�.Su��h��pR��W������et�1��������S�96����UC��tNP��C���t���2��CSJ�qU��\%	Q�E4>[D1�����d���sTdx\�_4�l��:�%����B8bs`��b*-� :<8��><0Ѩ��jr	ϛ�헚��z9����������xQ)�+�N��on+�wP@�����_=�\{oxGz�g�φX5g��{����Ipy@w��ں�N*��M5��*�5�ɯE���Y��(����)9?�y��T>P};J�dJ��>%��z�"���F�u.&��⩱WW�r�׊�H�@�B�ru���k�.2�$�Jnlt�v^����J���P֒zk��oDVޫ��9�KR�P3�f�X-�n���U_W��w�+h��W��p�49���Dtݚ�j����G�	-xp�d{u旊�2M��Ϫb�vUrB��}=�{�FE�����p�>��K*�o�8?r�ͤ�@� �1?c��8�g  �.:e�[ق��e>f��`'){�/f�K�R��F"��p27�	���7'�&3|�c���3f���<��{ܫE!���fx��ٌ�X�S����a
����w�S���ո]���;��qb�x����b���%|e�i�Z�X���� �B:��Y�Y�a.d�1��G��}룡
�%RZj������t��lp�}��x@��T�Ս�+��_J�EA�r���G	��~�� ?,�W��V��>ٱ��or߰�޸�(��yp��ƙ�����q�;�@�d�Oh�eb��֎q�	��S�m��42�qCyPB��BF�'��45�xW���H��e��%�+��=�w�iZ�NX�	]Qִ��6�ƬFE�n�X��qtS+h�m�ܾm8x���I5��1D���Pr�����Ǽ�D�v���/�`W�L�����kf"  �}}�ٙ��I���6"4!�<&�*6���cG*m�u$6ꜘV��^3E�7g�����4i��Ey}��9F*j3΀1�ƕ,�Nb9�vp�*;x�Y{���ك$ ڄ�l��v@���W�K�b����㮏�=����sK�^^�F��Qξ����� ��+]Q\�/ǅy����w��)��2�%�2D�#D��+�����M�%�&KE�s*:��F�N+8���ټoA����xdt�F�C��*��Cm�������h�?`u��H_cK�b��l�ٲ�ޖ:".6]C��� s%�f �*�.I&
�zon�F��^6��,S�U_\���
�xV��‘S�˘�K��%����n�7�ͧ���V�:���#17�MY�F���Cڎ� A���;Q����s����p��c��g���4ź��x�hUM)�c¶��53�'I��F+�H|{@�(�S7���7���;F�}\��k)�]2�|�A,ۙզ;j��Z4��1B/`j���@�uk�h�7+.���ݺP�R��xP�:�ۑ>G�)����N�s�/"2�kq�x?UUU|<Y����_����^&�y��}��؇r����Wԯʶ葡eZ��Eα�����^��-��8^�ִp��J]�
�y ����R��2��֞ān�<�EdC���6 �&�ƺ�uh�o�բ�w9�dOL�|���}��
���_`M��i�ETlҮ�^��b�Y�!��Ä��עeT?f'�@�l����&� ��:*�H"sƟ���8��8��k��~7�V*R�E�^���Ԏ���G2��؆bxT86��|��N�Gd��j索X5p{�kr�ȇ�@�����y�EY�T����D�P���?�!�-$�+Jz����(������F�B)� �]딜�B "���� j�o�1f�]���MIp�g���,LGA�?f����̨�Hb%l�0��jzX��P��]�M�I��"�Օ���N&�J�U}1�1)ı�e���E҇j*�틽���{�Z�l��N/;o����*t��+w���KF��pL!��D� ��U��};��Z���Z6�XChu޷�N:촧(N�ݦr�ѹReD�X��F����t��;���h���ʬ�}�}�F1;��bph@=��@b�رB�|X3sFm��0����r�M�|�V����v]1¤<+j:����Pd<+αh
�i���F��كit������=��}��R�1y9)/�pֿ$+@�u3��>YݓB�r�l�7�w)���W��;��L����o��/��)��t�K7�[E��*^)��0¯�>0wiq�`ǗhrÜ;�uЈ�z�n��k�j��w\n>Ȋ(j7�D��#LV���3]}��j\�tz�b����B4�N����&a��r�G
�!�j;���Ǵ��	ӻ�~��Ǽ�¯z�m��/�� LQ�lh��˟��v�֪g������<�����C��?Q����(����u���ʍ��XC�U��5�꫹�6΄)d��9S�3p�l�#z'L���hY�1!\�(z��W�e��)���n���Sh(��GP���մRW�u��5_%abV��D�)����v3vU�ܳ�Tث*!���M����V�U̽3�z1�]�Vh�M�[bN�@.��g�O�c�"=Q]�P��V![�����*�z�`���q��<ʅs0��s���+�"���˒��P`�>�&v>����]�2!�M��P�7�4���x �#S�5�{qn�ځ[�(��{����g�g��� t~��~;�؟���].�!�3�R�H�̣�,�mTbz�����d�K��	�W�
jX�4"�����bcXu�ql��ӜtZo�u�w^�g>Pߑ�)���pO���³lb�k���Ơ��j~}P��C͡c	<^)D�H��v�������a�]g*��N(=���y�h�	+��]΀'��O��48��i��4�"2�V�.�����a���\k�ꡂ"���n�K<>b:�ĥu���;�����١si��C�:.�kY�s��a��}(?��B���%���#��߷�1i��,G��ɘTa�M���+������@o���.��N|c��2�%���ŋ]Z\���>��u�R�w�2bI�|��ʳ�g2��=����7]3ݴ���8mJ��e��̴;�7:=�!]Ƅ�8�+�!��z��֬p�Q�m��9�i6oI�&�|�^^>����W>��l�C�u�J�^����C���dub�2�wW�cM�	˭�y�4q\^��Ԗ] ���m���gi�ck_m�j�SC�b��J�����&Ō��C�t��m��=w��֜� �t�R�=��t���:����Y Ҽq-��:I�A��Vo��֖1X��X�*B�_Fp��.�Y�x8�al}GU�|���;�N��|Nk{WN���Tz���^3`<��``��ɵ1ϕ�Pe�Œ<y÷�O�5y�T�\��HG�^�x=�\1N��F�y�0uJ�� vU���2��N�r�`{���uq&���X�.Q�g�O*Ǻ����,f"�PF���.h��.�U�h]��-��)Q��_1c0K�۾,�y�y���SX;����#8`�5�2�
�6���e63��7չQ�>�{;&����|�ocY�i�d��U�w��W���]�]�
���;�z륢4f��O�<�z�u�y:�u�1�l��ۨ�]fR)\�d`�U�4�-���}�x3����-d�����O���uc� �3v���k5�Z��Qk�ʻYp)y݉oL���r�-�f�'w����ǍE�����pݕ�攱�yB-}3��.���\�{�<�K��f��Gkn�z!�7K�Nֶ%oM�~tX�ɛ�j�`l�9mI
��/�df<}[�gk���;���J��3�����"��>"�bo�_Vns���D�I��3�z�ZKu�R��\�`9W���v�6��;Sjrl7Yki:���ٜ����,�}n�eZ�}r�h �p7���b�w��{�naח���t֞�� �7�_+-ȷyM�੫dee�u��\���Ab�0H>'/�wD��s�+��G}}B*u_g��5aܗ|�c���$I�4C����R�9�{tІ�֡wA�گ�-��9���c�7��xd����W%@�����!j���L��2���&��N��mǜN
J�upaܹ��)�7WNhZ`�Ć���{�˫;\(u��Z�V�I�l
��,���h��%�\�.Nw\��b���^═�/�&̖n��Z��q=-3��=v �ON�m��t�����mvԷCX|� �-'�w�X/���U�����ˑY�*�3�y%�ȫS��Qr6��]���՜�Z�Ȣ�"����w�죦���
I���e�5s��Ю|Gu���>)Ȯ��B��\�xw;OxdQU�<t�u��'0��P�GB3gL.bӤ�E4�]��ʢ�����Q�@p�J���=7%؅DTG�AY
��QQr�[��UDE¢�8�fQ(��Zz�2����E�s�S��3�tJ��Y5Շ�5��*�c0H�eTDE���W*��AgNйdQ��%\�D\�\�QAR� ,��H���V˶r�V�F�����8_���>L~��z�*v��w��h�mK�er�����]��z��dH�9w<��3� oJ�z�x��S�?}��D}&���6�h�kf2όS�U��Ĵ��~U��p���*���&�{ec�Ɍ��-��Uވ�
U���5Y/��X�T�����0��䝖���!d��1����|�Ɗ�鐎�)�'@��[S{$Ļf�&�oa����a�?N�N}��!O2�\:��`�ђG#W�|�cX$��}9�z�3:m���P�0*��%ݺȹ�u�V+�G��FB�ۖϲ�#7�w���f\=F�zr�K��l�@�
b۹1��T����ա1w1n��Ϻ=��iS�Hx��~��EnTW�KÐ"����w[���xЭM@�UD[0G ��&�n�=Z(�[&��K�E��)\�ѿvl�u�4(t&&3)9�BUp�� ���"���TCEneG'jrg�q��մ��cڮ��1���s�B��K5�o7]ۧ����ζ�g~'G�o���+��2���l�u�ik�M�ʴ���a����u�pF�q*�b���7�O��о͆72GW{��ކ��g-VdU�|b#��%�Y��[�A�ӻ��n�>cl�ws��g7A'���UUUSڼ�gw���Y�ٸҙ#DE캇qe +�,X����<#���L���pK�&��!�����|7���)��r�Y��o�-��Σdۼ�|W��#�W��εNn�=Όu�'Ta�u�T �b��
~�o��-V�a�n��:���f���9�BN�f���F���
�}<���$�o*GV/Eg�.���/s�Ո���S
z(�>����>s�;>��9F��=#v�j��oj�Ĩ�J�TY���u�L�����6�{���=ʇ�˛�|�HXÍʉ������Z�_^�P�^�']����[��۔a8P��+�ʽ���eI��gp�:���mt�y�n�S�5�J�E�c�ޣg��ܮF+�v�a�^Ez�[�o�T'f��!��9/z�,o��Ѩu����ݝ:o_���6XtNFrۛf�Ҩ���R��q�h�x���X-�&a�F�os�-�ӄ��*S[e�Ρ����=5���wy�*�ﾯ�����͘�^�u����)H��}5�>;b�Gui�U�
�$�\]?�s���ξR�ɊV�WN�@���|�ɓ�^hݾ��]Y�b�)LϞ\����1��U��/d��:+^�S��oQ���&�Kq|�����bs�J���8s��޹<�N��[O#��~��N��ɺ�O���_l��FC�;�ť^�B���-ҧ��صY���5J��A��l\�=�I�*��wb��Kbc���8Յ�f�u1Sj��ɝ�/�53:8�z�����%�T�	�ɫ*��3B��W�*%���FT���]��;�E��/��ux�a��t����O��
Xs���qwA�E�I,��(�W��S��{6k2qc�0L�7<���N����k��j ���;{qN�S��]�@vw;7�]�+p��B�Y��I(���]�g�e{�7j��U�5Ր���p۱���ޒ�Y]J�nL�4�w�����vs��3�`-�{Z\�V�K��_W�}U�5N6����}�ܨ���O��eɷ���ՙ���
gTҌ���o�w�VϺ�����{$�Z�5��rPHy���.]q�얆�gwm��n���c��wW�b��\�u�W5M�f�&H��j���8�{���VC�(�;`B0##���j;����t�o�`7Y�+��fuA�-�ڈ��E��9�4M����u�g�w�s���%��g]w��{>��N:a�{���v����e)u�qr�tڃtW7�(��)�3�0�ޖ�k!mB��F�>�*둗fz٘�s�&�8��r=q�YΞX��ѭ�;�������g׎~�Xn�GF�XS[hN.�p�6�وH4���t�k�Z�hl��ٸ�U��+uD�ˎu2�X��A_`��թ�3��lF+1&^��'}�3xmf��ҝF��L�n3u��&!;n5p?�/rO��5�V�=�GG;5���C}3�O:�yu�v	ީr��w5=���X�z�T���}���{�ΩVvh�{�;QЮ�o�ԫ�*~R3~�1[ۡ�7�P���Jѧ�1Aލr��3�j��AZ�h����T�V���v�\J���&)�ήhx��OݟMk��rw�3���$23��8C*%��qվU���^�3�'�y�{I��>�v�<B�A�Z$�N;���}gS������1�����erm;;$�|o���2�3���ռ��&��+��X��zL�&9���e{��㍅P�%P:.��s���w�Z2&��.�ܘ�?c̯�j�Z2�ʘo�[R�]ۊD��T)y�_(B�rLS����b��u,��;���M;�J� �	P�|-��wc��ط��#����)a�0*�~?kN�_����ʰ�H�����β���:�էl��s��%j�1�تzV�%\�YVZ#A�:�t��1H��f��S6�0����/�7h}8��a\��\X��;SG��G�}�����a��>��V�R"/X]_W�G�Zww�Wa�Xmw�&[����P��S[�~����C��Cr����+��jO�j�bLw����4��9
~�&y�:���U1u��{�P��T������fiL6w�;iT	s\P������q�6��tO��1%ȃ�l����&��F6�(;-�qQ)�0��yʅ<��0����n�"o_�K�S���󒨬[K����ue����'�)i��VHճ�����3����z[F��YW�~�3O���R����o1K9�Y���uyiʉW0�e�C���d�����1��Qs۵��+\6.�j���%���uزr�Wv}A�{�[^�Ӻ��IEoF�rb�k���eG2c�1���:uf����E^��V	�j�mX�Ό��gg��VE����O��y�$�:��� �ո&,%�`�T���e��Ǹ��6�Y:��$��Q3L�Y��訹�D�5Ԙ���ع5s��\RN��Z��c
�}_U}_|KE�=��Wꬎ�d�*>x\.t]V��^�U���NW��۞���T�̥�kU���o
M-����3�E^o�n^^{�;�~�nm���B-[�s�c�J+���t��ФJWc��%�2����˦{��v�D�9��v�u�&�oIQ��[��b��UA�P�o'��x"~��s}9�Ӛ�(�j�I�K^�kt��a��:I���	�Q���l��c#�u9�{3q��<�3T;Yu�3��
��q�g�qΣ�à�-���j�k��ջM�݁w�r��u}��[3��HSC�N��H�i�7m%m��ȟ�0->��c���͈ՠ㽖�*,�(N�����F��F��|�4;(�kb�n�=?�3߯��wV��r`��D~��U΋���h�[��Ø��e�̩�m����֙�2�N�CL"����P�V��Ι�dowZT�]�B����k+���b=vr�6R9)���2�}W���9�Kɤ�hN��4��UW�_G��1�[{�=��5��GC1I�������kj��B�k7W�Xg�M���ɞ����K>r��eMY�5�!o���)��1��Z�9;����p��l��9��(S��b���ھWЯF#0d!
�aJ��m���T9Κ��,⯬�Z2ۘ��]\����޵l�J[Զ'w��zS�U�~��c���oΗ�)�a��9�v:�"��m�sr���[p�fU[�D�%?��kE=�(��"x�/�SپWvWֲ~n���a,����c���NP�l9��"�+y-��c�m|�dӥPݲ�\#�c2e�]��ow���������Tb/�PԺ�JO� .l�T����p]8w1�Ρ�U��޽9=	����j��T�d�����;���qW�1U�#:�M�M��/kk�y���Pf���%�:�Ҳ/�
 *m_�WF��V�h}A�fdT�yǷu��ƶ&WX��^ �Nu�f�5����-v�+/�Q���ꈈ���z�;��<��G��i칯�y����ٞFV������pj^g?S"���J�0�3Z����fb9c�W'-}e��潞p+$;����J�e�|�+�[=�Y�d��J3N�f��Z�\m�mWE-�è�)	y�6[�8���~Q�N^m;}�O�"�=/˨<���ڊ�F)AޥK��ھ0{]Epn1O&�y#-�ULEf:�9�-⎎Pw��g��Ũ��˛B��^���/����8����K�s�������
5�@׫�[Q�{�\�ݵ�d��H^/�i��̀���u�愚o�u��Y�9���C�IyC���!Ε�ħ�	%����>��F�3�d	�s���:��v�8
>���6�|����B�O�%4'<�zF�H���	tW�^�)햻�{��[t���;ds4��i���F]Y����j��QmǽPv��y����`Z�P���������'���b��{A�Cf�m����}Dd磞�^�U��\7�>r���4�|���Ц��&�f�
�:,���r���=��J;��kdT���G��+9����˂3��+b�9o��9�n4g8�������n� ��ގ��U�.�Y<D��׏����e	���V@��B�V+��w����Y�rwsT�_\�+v%����+��=�;��‌_�D�&�)oOd����K����b��q��WZ���e2���7�c>���z��9��&y�:�n�+������K��&̃����{��ݶv1`3��\ش�:EGn�����RFfդ��j�orۃ�ʋ̚����(;-�qQ)�)�kh>Ê@���ى����}�-��j>sJŴ�{i�
��*���ʼ���(�����F��m�";)����Y�fl� �p�4�B�ٚ3�8�&��9�V2hn�N��3Y:����Tu�x��k:��lu;�蹋����Ɠq���Eh�8��[�;XǏɔ'v���[�f�����R�3p���	��дb����$�*U̮J �\(�w1�V��� �b��N�mr�Bt�A�dΡu���$m�jA[�n"��9=Zg��񡽼r��VS�t0l��{4�vs&��m����%�kCb!q��j��Zʲj'Yy�C2�u^��Օ7}��g�u[�!�2�փ�13{�+�q�����s]ùv�4�nL���96��ɚ�FK�z���^?R,��Uy��&�9�	��i'��ˬ����yaN���|(�к�1}���)6��{n�U����#Y�gh�)<�-�TwK"�����A��(��L��c���Køj=�|��=qX{�R��v՛r�|ҕ����b����w�L��9\4�+y���.���f+����c�֫�"$,�Ok��n�����W�a�����e0� �{C�h>hRg����+2<��S��*�gb���4�ω&�� �u�|z��$�mTTy�\7.Y�����ݸ�E���F�b�J��)v�q��H]�*Γ3 g_!V%esOix��2����)5��ٙ[����������Q��?�q��\�p�'��M@�F,���՝D1\cH��2�s�pAj��C6�z�Y�ȯs�S�`gb��wi�=�zhm�"��ݜ_z�0�R�)�ȥ�ɭ\�������w�m�
t�'wK0B9�4Z4�cY�}��,�
�7�/�r�இ&�[�n���B�r7ٴ���3.k
�m4���'5+��7 ����HQu�"�X��i⥙�83j��H��� ~t�-�Y��S1�����(�ٳ#��yʈV��Hi�fή�a�Cp��K�w|�A���Kdc���c��4��l̆�!pv�^]!�[�
C�%޾�ޅtR�V�[v�ӳ��=�y�i��9f7�7�2�})�xq��9#\4N�6���ep��Kb��u4�U�r���'�b႙��ד�wY��[�f�ܸ��8�Y��n[1��k�'����sI��{+;"j�����m,Σ�����KA�������@��	8R�*�.G*�*�"�t�(�ʂ�e(*��NG�y9����fbP�Eɗ�ʻ�G9Qd��Fe'�J�W-lL�U&G�-H�KXs��p�P�5:@�����ƭР����ҎNIq�E�@E]�Es�AA�S*����)��\����E��2N��U��\�t��	Zp�LԸI҈����(��©:p�U�REӑ\���Q+�Er���D9�(wBsѹ��i,�:�\9U$!�\�E\�GÔ�z�9��qݬ(�H�D栓�{��UPU��O\���"9p����jE��}}����߇�m�I߿]�
�0��E��`�Ծ�$�;�3�՞*�B݊�G_R�v����?G��D@��bm����f�5�0Ռ�E^�7��o��sr�N�7���\�,�u�,َ�?,���r��&��N�9��v�l���7�/�ĭH��wk)pi͚f��1�78Ԝ6[��ʹW��%<����$7�|~A�r1���dWҙ����r��^����۹K=T9 ��9YU��o���s/���Kr�� �"GY��}�`�c2�
�lvW�̥�U��E,�R�c�`.	:�]�t��R�8�71Ô�P܊�nm��pS��>1������{��sB��)�T+5��԰9��#Pܲ�#t�]8w��ʦ�B:K��7w�@Ϲ,���㝍\��5hq��連r�ժfvZ��8��U��Z�M_�w��M	�����i[1<̗ndh��,���U��j���Z�C��Cu�W�J�f#�V��޴�v�]O��3�%�]:qf�im���t,���άl�![���m.���um�6�絶j��|�K�:@�v����S{@e>�sf��DD}��k�B��'k�t9Fc�=�\B��U�R�c�D$�wg('��U�d+�jD�ܾ����s�_Rܜ6��ά��Q]�6�,�� +���j�=����kϗ��Y#'�����4�l_r��/�q][Uf�L^�љ7,�>��I^.��.u[��f��ߺ��Z3�����8����}��,x�>]E9B�t�7��K��rn�3�2��w���3�b�G��uv|����7���7��R,��y��C2O���+�f�mDJ1Z�Y�a���b���p����g�{��6W��ƽ���P��%cwO�Y�Q����)�*�]�����R1��o�B��|l-�������zOtO�����0p��9o�]
����EǬ�ն97+����Y8Q�hs�Z��ι8���.���پ5áб���5[��Jr��ܖ��y��f�E�%��-f�vٌȅ�1zk������{i���}b�����8 xF��Y6UU�ˍ~��#�ۍ��h����v��m�,�鹾�J��	F�Y/w��Ys|���{�d5kj-�u��}���)���cGW�D\lf�Z�����䟇l�*��5��Cף�[Un��%e�b�8���+�3�G0$��EAX�UP�޽9=	�E.���u�����z�3Ы�8�R�q]�]{.i��
���FFtUl�a�2kZ;��ꩩc��oR�uk1�}BU�r�f��b\�Q:aM��a=��ɗh�:ل��Dt�vD���K��Ő溲95����H���5��z�6����C��>���-n������$��57�)�k�<��<]D��z���y���F	�L���z��m����ڋx�G(�.:��Ԍ7mM��pv;ˇX6�ǐ���TQm_p9k�־�r��S�b����ה�K!����;rS3=�����$�N�zx���im�l=;v�J�i\`�����U}as�0��t�i+�֡(�~�r��Ϸ���R���-O���z��p����?_g��wj�#j#q����^����>�ǐ�Y��$��%�w�5S[���[�~T�Unr�ڲ	Њ�8�DqcHT�R�Idl���(3���lMձ[{]ՓGTB,�'HV�a�x�"��-��2�U����qz:PUl�MT��g��7���P7�����:��%��ZحɊ���S`ʌ�k��h��-B�X�K��w�\Fj�-Uxbn�%�Ld�yweկ�}9�z1�Hh��<�U��X�m�rm�5�ws���Wt*����rC�8S�
v*�[�ʃ�@�SUG����f�.��u�ϋ�n�}J��=�:p:xX��=��ɛ���^�v&���q'^�ޫ��y���Y]Yu�G�f��^i� �u+ot�د0����Q�XΤl���QW�j���e�������;3�C��!ġ� �vĲ�'	@r�dR�{����%��IwW�,�����Wr��M��~�>���gC֗<د}W�wƫ���X����K+b�d\P�yջ+9��T�M���E�3������pr���T���dԊ�K�&^�i�gAח�5��V(?l�Q�B�fTJ�]�N$hc��B��]`�to���E��b�O�
$�/x�-��S��קkў���g�>��nYqyQ�UF�>���]ӂ�h��m����9��^����2��v���i嗜$9MC��I(��Dwi���^4��3ݱs6�r��X�P٩�Ł��#Ds��?E$�ˠ�m �{���'�-�}�^�.�r�>�Nr'8.mD��݅�ލ�|�˛{?^��s��<���l�*=���9����
���"Y��kZ���_¸ř����3i���N����Uo6�YҚ��}b�S@�[��N�t!��D��[Д�� �4*S�o	���I�v��͈��J.uu�z��e����p��kh�uЬu+�i�"���U_W��������v�rᬷ�ǇTѱ�FR֤��v6��ɽ���1��S©��+|�9r�4�<1��κ�-�f�s=nW,�ZwI�O�y\�b��7P��5V�M)F9���_*�^ڜ���ع�kr��s	�퓉�?)q��xu�h���;u����0�Z�]u� ���*��
u��z:��Ew�K���B�p��bb>�����Ϋzf2٘��=wʹ[[YSm�o��7�%>���S�@T�o���uګǵ�A���qِ��Λ�\�6m֑�)-����>��
���t����qI�0����G�N��^}������!`J�m�'3D���{e^&%��%�G-ź��T�MMp٠��S�-�m��s��XӋE�o'���iH�"��g{)�����}�8�)6�����)��K��әs�Ҕަ��|F�5u�kP*�A�ռڮ�ø퀢�����)E�u���m��ϑ/R���+���w��g+~���瑱���]�k��D���>�8�#,����r�[y�uDB\��F�������L(��Ͷ��~�!v�G�`�ͷ���i�a�ٵ2�Ζ�9�Ƭf���5�k��r�u�v:1�D�R8�ѫUOKĥ�Sw�FF��voi|������2������Z�+w�h^[=Ֆ���Α�ڝ�r�n����J��Q�A���iP�n�v�b9R����.�ퟫ��c����S�0˶y�ӱq���&�o�R�+�$wGgW.����Q�4��(�Sj��/#q<�J� �K�]�@��T2��������?SN&�Y��Nu+��j�w�R,�����E|{.j{�&�[�Yɭ��օH�^OP��_t���%�f>�����g��h}3�d������zy�qjqq��8�MЎ���/7zT�O��z�w¢��E=�/Z$J�Md�v J�:1Q���N�R�*{0K\�����P=1,�bW�p�ʊ�~�������s~~��=6�H���u2݅�)���>����ή2\f�.Cs��oN<b۟��W�2�i��� ڋ[c.�K�&��[�kE��F6'��M���J,�9�k��������6��LSΫs��(Ǫ���7��y�^�B�kVzv�����,�E3Y	������m1�wH���+�b�6�~y}P�,ѻك�P�ʶz������Ϩ���8ui��1o�V������yjo��e.e�Tz�%������M�`������?r�gmwi��׽Y�uf�J2]iv��u���Վ�7�!�ttϧ-ڑ��4�X��f�-e�\ɾ	Ʊ��GeVgú��ݭ-��mGŵ۞��<� �\�M�g�w7�P9�i���Q ggQ�j-��ޕ��KWڄ8q:8f��� �+][��UԉSo6ĸ�ú�0�a���tx�ݚ����T��V���π�ٓ�ڵ)4�[��G��G�e��%���M�EE��r�*�Aj�ɫۯ'aTs�=3����'�A��\�jx�5P!\�V*��wS9*B����m�uڥ�فz�66�98U�D�K�.�
�bn��֍�Ε�.��Ω��>��|��.>�R�Y��JF1����*n��i
��qp����OF��Ʊ<���_qJ��z����-�7���W��ڬ��F���g��BZ�ښsqa���D��5�9O�7?G�[ͬ胯*/2�ב���(1��Ÿ�Vk{V�z3���s����ۨ6���^NWر��Gn,�����沸m�׽��M�w{�5@��ܭ�;*3��6���~�\}Y��)��P��o�-�!��&����T����⻹i�pf�ݱ~9	���* �[Mdčv��[�s���]F������5��B��<����"o_Gk��W�s��q����k�	�����60�;t��$�m�.X˷vچn��� ���""#���W7�Y��ي7�Ѳ0W��q�]"ڝ̡b����������_OA��N����\a�Ƨ�@��Z����r>�Ng�Ҥ�u��ſgP�+7Ӷ��<.��94��vFS\[��ռq۵P0u�
wࣲ�Y]��������{Q���ǹ�N��K{--�wlu�c��Ơ���"ﮄ��ގhJ�m��Y���x��NQ�r镟�7���S����QS�uO<sE����覦b��7A����[�1JQ�Țյ}K�����V���?l*����1�잨��4S��Es�̎;�a��s�����=����9F_7��Yh0aX�OW�`���ꀮ&`s�*�73��zg-��M������ob{X�U�{���䥧�R��*8��m��Ǘ{���I�,��6ݑ������@�|N������N��.
o��ۖ�䙺�XkXKU��-ۥw I��2��$VV�Q��"j�դ���X��"�u�S�)����H��1dZ��jM��:��&%�ǐ;9&���1���>�8���sەz�U�

���[2G#D.$^�t�ʰsu���s3�^�m��fټ����P�ܝ�T���,���n�Rsd7f�lqn��^�kk/v��)��U�!�,�\��'}3�fnPlZˊ��pf�7��`��FLU1���,�hb#DO���b滁^ق����D��t^�d����[��>q�����u�
ܗ�ЛJ��w�)OM����N���fӴ)�A�h܊��٦n��u�YH�}�yeh��&j넭0����w��k8��Xmc%����ܘ�����(0or���U���N̬IPT�;$fX������:��=�w �\�v��pøU����g��ew�-8rk��A�9������[,��7x!�
xH�۾��ACeK^�hv\�5���*��O������	Ws���-���e�N#���5e�F
5%�G�J�,�9bn��9J�:k�.��r���Y��*�������5��XzjﱌjԵ�'1Z���t㖉���Y�G[����
������n�����R਋�\�Cx�ᔲ6J��t��OK2��Ty�hB����ǋF���w*�)]EBߦ�.�[�*�T㼮mvv�-�`�J\V�+~}:���m�f���K���5�<�K���q^X�>D�c���A
v���`�����V,Y(�CR�y�mY*9�+;�bw&����WB��������7I�mU�Z�;��]8�.����z��ӫ��mŀK��sU��a:mQ�V6�;�C8!Zlޒ��DҔ�r��<=��x��p�J��[z��Y[g�J�Ԯ�@B̠w�E�;�Ir��\���� �,뜖�)#/��w.��ټ��ݥN�B��C�B�v�u'aw<��e��N��o��7&�A�\���R�z���l�m������Il���0jZ�"��n�k(8;��_u�8�b�QGj����{q[���+jr��չ5�4s.p������ͫ�|�9���$�卖O\�m�r�������T;��ô�ZJGsT�c]/�R*͊]�S���,y��*��jG��Z=�{x	��� �s4�0:N��������B�vCy�:q
;����
�@�d�K��KD(*�*�Eʢ!Q��<��ts<g1re�W�TDS+�teW;"��3uʹ]�Aʂ��*�U]�J���GUhWr��"�U�.ʮ*&r#�Q��%�UG9AE�a�^'&\��C�E"&F(�8ܐ��E��"�w5wbL.Res�(tNGn�s�$����Y!\����qʑ�M��
 �I��DQS��r��w��.UW�&�˄�'3���rL��2�TU9�P�ۜL��(���]��Ey�5�
��S*�(��T쌄(���u*.��sΧ]hҙ"�a�z�7S!ersB#��r��.P\T�Gs�p�7=��t�?�gw�_=�����޽��NEV���ҟB�9�rP��}(-qWN�"����O��fs��\���^���>��L��m8��0�����e���h	�����U��b�n�Δk��,��?l����	�-��x�������V�|�E��N���ﾢ���[�c�N�q]-1���Q����0�N�աt;i��S6��}�7z3�F��p��`sϬ��0nc�wa\3˰-�W�������P�u�F�LX�SP���:�bv���j�[y�z�ݍ�f+Z���Ծ��oh'�q���Ć(ӄ�G���jV3~Y��MOA��4�M�8�1Z��;\�����ՍW]v�_B��7�i��u=�_���>J{a�s�x�dF�n�%���>N��]xc��VK�n���܍�I"%��WD�n��~��Y��[�q�N���
:!�#v��/̹C����_M��J#���9���-#�3�[y��x�.���(8�nf��s;f���a�}͛}݌f�6+����ԧ��l�����õ8i�p�<�*E��{Z�j����Df�7W���7߄rʒCS���8�#�½<�V�b{����5�gp#c9Ś��2�j�u���Pʪ�ע�n;n�r�1|'Z��oҖc�GW�*���y)����T��~���׼��B�s
S��0Bl��֤JʍG+!h��4���i�����50�s��e�"a����(wI��1p�ѥ�s���S��Qx�6��R�.e�2�nh�0nַώ�w����V�������e��M����+�U�ʸs��=�W�7��1��fڧׯ��n�R���S�;N�
�o>�/̼�Wa^�[(WwKiSW�V���=(��׫7�ա����x���7ީ�*O-�fۯ��m$.R�S����C�>�kI�AD��b�_nm�(�PΖ���{�O��Z������7Mc�κ_vD6S��y2�H㲱�좖��Q�S�ǫ���tc�^�,�![v��U�3���6G����f����
c�%�
��f"H]C`l	��g~��ﾢ���fW�S�ޕ�ʨ�vro�s���~�}X;DR���B�^�(F�y�Qe��:�4<�.���ٳ~|o�u��=�gOp�,�̯�bz*%�U�u�*�U����fG��Ϧ����~t9���~�u���Q�}٭fɏ��M�7ռ�6f9���?s���W|0%C�TI1Z��U�X�[a��_ew���3_��t��T���.;>�B�s=}j\B����f=�Ҙ*�X͗�0-�&7c��V�M)�tw\X�yC�ْ�>���᪽[U5�v�a�ݓ��|���p���Z�d�mMɬ�Q1V�q�Y�Җ
��ȕg�=�}�V;���s��Ӭ�cFU�j5��2j!MS�[u��ŀ�zV�������TyQ��`��#�J�(�ǀ��&M.�s��6�u�M����D�=�7���݈�r��;Υ?S�8�g�;]^��Q���wS%�b�;�6H�IO���x�a��9M^u���]R/��ɺ�Q�L�R���2~۞��_�:��mh�{y�~���g1
���OI՝���[�I2/��| ��t'�J+��R�j��y�뭬ò�#K��n+�e[3���Xܲ�򠪣�T��2����O��X��;��U�=��m?
�c7k�����A�(�����r�SC���ǩ�`��U4�D5}�F��WG*l<m���.�J��j�ʠ�n�j�{�s��5��}�R[}��}��ץ�گ*ɴ:!����E�1oE�j�;�8Y��i��{-�����C���U���Y�R��iO;J���t[�����oF�C��c~rU��p`��lnz{�s�jl[��ngT�OW��t�Crʸ:��u�b�yhߚ��B02
��^Y8C�V�f��ز��������l��n���^�s�W��)N!3��n��k&���M����Z潦B�rL���G��1M����B_G��j_.���hsK��UW�]�X�w�(5��,�^����n�s�֚��~�O[K��)Sϭ�}ʌ{�y����w��<���=PE`�0�w)�\�������]*f3�t����i�{@W�'1�tc"�5S�v���-U4�/���pfA���D�ܾ�zg�{�<��f
�2�c�R��A���Sҕ�ȟ����F6��茦��7s�j�>NyԪ���1��G�S~�꣕:�0��YL�<s��+4���z������:g�r��1��t<�Lr����%F�b���~�y�u��,��(t��|z��u,���:�^'���Yx�I3Tu�r�"��o��(�����؇�U�&�)�y���ou���4���ʆ�^P����iWZ�E�Ue�]�N�u�:��GS̈�ë:,�r�����q���M8�fd��kٛ�n�7��n��S�Kj %�$:����ӕ9�0gX7P�oqF�72���r��-y�;����>�T�����W��6W<�����D}m`ŉ��󼕑����t��r���%�ad�X��+ٴa��z$���A.?R��W�N�͜`7�����coo���ˍ����.�&��ֲze8ڝ�>{^�{~�_vǸaf�Tt�S��B����
q1\�}}�}+2a�7�/�����n^A\[�=�j��WO��v���K]�ՋLO����>��}�]��}JQ��a��U��[lg.����=;W=�ߵ�?��MD.��n�R�b�WTS�e��C"�o��[p�*��Za�=�s�!��j���<���oU�����o`qL�v)��gl�t�k��7�\L5���2�.����w�H�!F�����ͨ�S�,m9ڥ�<�0���C�м�����ܱ�JRZ(�aun��֣wx�x_NuK�o4	��kg7GUŃ��lVf,��IRʻH)]�cr�Aƃ�&��9���w^�mYn:�+cI��gq�ݜ�L�qM�������UU��o�B����:-���V-�޼]A罴�.�9B;� �uM޽��P�B�x�u�GeAʚy���-�Խ�����p��bx�>�/�uw��>����N�������[2�_��թ�c��]�:�q̨�q?6~�ޣގ�:^K�P�-��>a˃�὿O���e*��Q����f�ܿ�a�N�:���/R��d4c���h�|d��������nE���:Yj�d�iw��hwO/�Jê!�?d���]1A��ER
�V�h��7���n�s�ͅKT:;*K�)D�55�5ܱ��F�mJRJo�W��ʇ)TC��{ G)�I05�Z��v��%v�I�1T�Q	�ꅁ�S�!�k�\���uÆt��6d���S��5lJ��ʂo���5����Eg�ίM��uD���[�)�F��lk=Vs/ާ��}���}�&/����R�z�v	����h�UjTF��O�<3�j�}W�3%�BR���CqD�Aeo���"ԽZ�=w����9�ݑo�cw���e�5���.���]�1S���Ģb����Ԯ��S{'�>u.:�ȭ �^&��@�U�|����;��Dl#.̵��\�HS�L�8�b������Ǜ��
c��+V�����}m�ŀ�F'?GJ�U��;
3�V�]��`[J]�_�_6������^��0���2�k��ۨ��ӭ0�,a9�+t���A�uox*co���۬�U�gk��Q:��G2���n�j���ja��[�G+j�kbV[��׻;�F���:[�UnyqV��U�4�R�ǯK������nnHG�z��|��M3��:�^�̭w�L�R�C���|kF�Z�YT���5w��٪���3Y��cDXOjv�U��]�����$��*��=;�}�r�"�]6	�Aj�h��	�)�jL��\�y3F\\Y�\�o/�=� �vj)�c���/+%*�W=�c3W	)?�""&��y���pC��Kj�W��:��"�άr����VX�s���e��[.�v��%�Q�J���aU@�쯥�J8�SjN��m&���p�Wf��%���t��P,wW�c�m;�Xw#^��j�P.�/9�n��ꇻ,��P���nQo�W�kWZ��l�R�&ıvED�C�b+���_n���ɫ��U�7wX��Y�Z�����J�VĞ��UX:����m�ݷU�L�v�*h-��v.�,���U�u�r�>oo��ڮ�2r�B�<�[	WK�A�5,�}BU�f*�ޒt��q��C�[c�q����P�+\:��n��T���}_U2�@�ub~s��osxfu8{ۯA߱�[�d&�r�[�7�!�딒ݬefN%�L���f�9�wk�(��nVJB�v&����p���ŗW��XP+��`(����U��k�O��nN��4��`�F��.}�v}��5x�����.c��jAӢ6:omF���DD<���,h.�Vݧ�sv���\����+S*2T��t���}�ܗg��u�/���q^�䢋x����1Λ��O[�E7��n��u���6��C����W�s���P�����P�&�O�z+�s�{�v��������kUqFN��ړ�C��վ�F�9���kX{��*ɣS���8��|���7~����|��ߟ˦(�/����*��W��hYP�J�ֹS.�q�_���c�YҶO?�k�q��:<W��lm�sv񜫾k�7�d!���������2���S`r�EY��W��l�?��T"����rDTʆ޹��޺�0^!� 5p��{�1���0�[�H��>P!\V(ɜ��^�}W+޳=�K�֨RN��Y�B� J�}\�n�_q�6S�Mu�VT��fSUN۳ܪn��l_]O��U2���\[zop薝f��U��$�m�dF����5�
.��Id��a���!�ϒ
�W>#�5g��Z��}�Ɉ�kz�L#6���-i5cYsC
�G�V7a}%vz)�������䏴jR���5�� ��po��l�[��2���)N���l��op�.���a���4�V�7��#v&�˻:y�u�F��KFmj�-�H�s�6ʚ�;d���n��H�Ԛ���{D:0�<z�[��Z�r�m��}f�@'M�}6P|8h�Ӄ��[�-0kBKspSz�D:�@53�;�*�<��w-_mpY.�<��N�4�t�R&��(�^�y+����>M?�����}�\�˱�����m������ٗX�'��K��[�	km�yN�+n}�2�pH�NM�98e%��D��I�0	"57�w/�����niyolQ�wi�����N���]�/�0lqCJ�sT�ccYbu	MQU�^�[ϸZ�bM�ζ��O��V�/8m"L�����p,��gv���+���5�5Ge*��kkpV+�cc9�n�zu�λ�zT]b�1d����5� ���7aۧ�E7�v�"�z��T��������D_9]8N���P�3�3��/o�QG8�'�����6,;ELh9��I�X�ݷRb&�F,�c��iͣm�`��yp�����&�l�\�U��2����n�����QY��?�
���͂�͓� �&i6����{@���@��wV\��E>Ŝ[�19�jua������YzP;Ť��譽�Ux6�
M8�0-��[�ma�E˷���6����W�f�`�z�����\�+z��dǱ�T���&+��RNu̳P樂��x��+�$�V���|�Qw*}��T��ˌ���D�7�����j��d}bhZsu0266XJ��ާ:[ܓȲ��F�k�%��hc�Wsph�t�E���C��J۩[n��?*���8��	X��totx���$˝\�K/�l ��YE�2e�籍DW*�2��lv�i<;9��ֈv��L��cq��ޑ�(�ͣ�.�eNCYM�"0q�S�}�V�|�.��+�]�j�
(��J�k��[�^���!S���uO�̥�H[G�؞����廙]�t���-���r	حI���Wǒ���eNqnR���&�(U�*���)�uԀYg*��ȧ3���ۜW)�$INZ��Y$�@�+��p�:�:IS* ���q�Y	��"4-֕U���H�#ԢHJ*rL�� �Ѥ*\���"�҈YAs2��E�Q8�-������N^��{�ܛ�!\I�"�w0�S�A=wi�Ö��Gwr�'%NU^q�r�6�3�#�*�*��T��T�kNGe�A9%��'�*
"M&�ng��$TP\��8Ei�D*S((�t��rr(����.E���	$;��9����DQ*�p��Iʪ�kw�"�&����Su�\unBUu�^����3��.\��\���ɬ�P"R�e�S�y�+�r ��J��H�:D��\�<�s�Cʷ'aG8�I��9����
N?�>��{�ޯ{��l�9����I�)r�4��+i�CI9:¸E��mN�-v�m�z��F�z�,��]��G����%�N1b���J�ؘ�㩼4��!v@W1�jOj]����/)&��ږ�݉��Y�q�q0�D�L�}v�e���˵;Yہ���c��i�՜Ek[�`7��fUjv�>R��f�D���ux�1`6�DmR�&Ɐ�觅g;�s9L]�@V|�eYn�Y����-��;�a)j��(��Пf�8��ntc�>�h��߂����Z���p���E�k3�t�׫��*/eT^x�M�Oe��VE�;�w2J�@�L�N���7��N9Ҏ�S�=��嫈{Q+�W�hN�,kr����*u���ʴ��s���?g>�'��D6w���`{�#��K/%گb��7��ϔ�.�+T���]���G<E{պ���][{1������ֶ���"XEܛq�:�n	[�Z�;��N�h�e�[�xC���YN�K/0�LK�bZ���C2˦t�K�p}�"�yc�6[���cgZn��i'߾���/m���O�Λ߻՝��[Y�+%��m��.��親R�l�ۆ��u�=�<�G
�*�tv�MV��]GPjB�v�����ݖ�z�j������W@��|9a�ֳ��%�Ԣ�9]:_Е��3Vs�e�넃��V���� BY�7+4Z��]�������׻���8��iH��Z�9QF����/5��LB���	��
�c{j_4������]N��ks�|DJD֚]
�_��֡�<Ӂd>h�XUV=|9��6s�;�i����*�6�-����8ڮ7ݦ���8٧�l��)�v���������e^e_��GF���9�U���W��ce�	�������^ёѝ=�93}��)�_!w�)ח�٪���E��*7"�.��k��HHjV2��)��iN̫-���m�qs޷s���KD�tܱ�@+H�v��Y��m�������\��Q꺗�Ry{�����҉F^g�#���3<������)�C��&uf�q].~\�ǟ6��yg)����ʁ1���M�O�1Sn���:1ּ��A���o��k{CT����t��K�77cjZ��S��^TF��Ɇ�@SO[��{Ǵt��c_w�⫻����PR%�D�@���Nd����{���"�W���vБnuc�����'`�T+!����d{�eQ�e�wc�O��U��|9��Vۥ���W*��Ɖ��
���G�7Kh��y�ʯ:n��c��v��"�G,������Z�$·��e�ά�wu�Yoi�<�áO����O&߶o�g�9
΍7ʇl�)����u��T8*�#�{�:��kS���1�sP��}�9]�R�{�HB��(wa���f���=.-؇�u3跷Ϗ,�T4��<s���]��ϣH]�h-��<zM&e�/s���w$+�Qu���+�س�{��o����g+�e=.���K\4���:nF� )8�p���Y�O'B�tbV�Һ�+��r������e�?���KĂ��-mbҎu�˅�[L`��;KK�����COY�ɘD(^'!O��1����&��o�le�*�t�x�2����mj�q_�-��aۘneu1�u�űFS�g���.h���'7��qG��aVm^�?U�ׯ
�fg���owUr5!�;U�t�nh\v�)�ٟ��]K)�CŻ�e0CWٳ�8��`��K���+l�g,��Vq�b�R��Qɮ���c��o �o55�	dڣ��7�ݍ�F+Zp�.���*�F���(��h�W�ӽ��}C����,�5�F�����?l6��OW
�V��=�D>�^�r��'of�0����y�3���'G�q{7�a�KxmM�0��e[�w�;��u��k��<����yöP[�6���ݞ�x�y}� c#:��MvtS�R��RJ�Zt����ēf-���0A͗f�Xwp�w8$���3R���R���5[���ǟ.��6gE�����=ϛw�&pvR��Z�w�V�s�}�.K�7�pN�(bZ�=㋏���o�7L���/�^I0��gU�"���!�&;/f-��іo�!�����p��.q:�QX��$ά������1x�����1<�uCx&��!uv;
�A������U��+5�l���ٮz��拇�Л�?=��,��_<��9ֱs�������*��<s_j��ô�GL��=wS�gK�7��L���T�7�*����ŀ�ZsT�8��zMŪv-
�$lcהط��:a����ʷ�����Ũ��@GOi�܅�[�j)pV�o??h��tm�~�uS��R7���:8<�%zbW����Q�T�P-�-3���Jג�2���#�kU��Ʀʏ��ӒU��'b�x��S����{s�%��pp�坠�dR��Wu�)�\�N����G���P!��]��]վ��o��N�IZ�\wq�o�P���հ�*/<r���H����PX�:�Ζ��Z�}���^�<�����w��F+;]�86���IlohX�s���ƹŪV1�[墯�I(ջ�/$:�5���*�g'(�4�z�p
8�sh�OqN5h;��7R��s���
�3�;m��::�T��Ľ곮�OUr�_��4j�w�d춒���pc�ٸ͹N��rQ��������]�l9�r�.�*��?_c��1�SnXT0%CVT��J�]�b��RW�����g�w�=�oGR��)Ж���V���o�Sb+9-��a����r�f�4�َN[����0)Z���֕lʚ��CT#���d�N�d&a�|����T&%�j3��heC��;�d���>��������A+�ْ��R�ʒ�bQ$�J:R����J���*x�ӆ����ك`��-�r�}/,8��e����&ؗA�Y��-h_ϡ�n��5��H�m��
|%��fJ���#c_�dM*f(����V�K�mg�gM�{6���Lw��i�?ep�����i��O�UN��[fcSwg�v��'w����jP"ۀ�a�
���-�;���pV�8-�ۼ͵�.uJ��Aq�J}�GF�u�D�o���;�"������S��ɱ8&��R�����x�T���sV�*dn�8����Z.b�rv՗���M�b>uQ���y9�$�1�zLô���y���'�lsetl��o(�3<�uf����|�xSg7%����yz2�Un_��l>����HOȕ��(�N�׎��{|"����Şq�eI�E�7�|�%���w���O4�mt��R�����a�k�����cn)��*.Y��/ej6�AZɭ��N���U�҄쬞�&I�Օ�(njkNT��G!��O�[���j����q�kkv�����[���et�R�i�_1a����g�9r����gZ�F|ܮZj_2k��i��[/WQ�
�Za����Y��cu��E>�ލ�ξ��5���0���.P!L(�!8��-U��Y�En����B�����UzyJ�+�7�8��_Q��ܮO1o���
�#�BQ�&^.�ڜ��EU��B�R���7��6u�mʱ3͜��U՝p#_)q�	�*f3�u|)]t�d0H�%&�t�����r�����9�T�{.|��n����~��8��1;c�������4�#���)��p�5Kp�1�+��K���O���|�r�ꟺ�j�n��F�uB��ϛ�;��
NZ�@��݉��f�s�vQ��{��9���kO�g��y�O~��BP����7K!�ۧ#r�+����mT��I�������=�Vs��V̿-O���=�o�W�_'��Q����5�S��ڷ��N�cUlvX���y�W��u�Ơ��t&�Fq��,u7 �xy�WRb�8
�޼;��)��s$�;�L8yN�*���������WF�Yǭ2`���k�ڎ\p��U��U
�w��J� �{�wuwPa��ct��DV�n-���Ly��l�4ƾ��Մڨ�h۵��� 4�['��5�'mE�����;�=CG��F��3���R������z{j�k�q���8��8r�֝OR
L��͛\�W(��%l�3Q2Q����{p��UL��<��א����Sv������Ι�k�j���ֲнi�����b)!��U�o�S��b��@��6��'?%��m��'~|�f+�w��7��;��8�;j�n�\k
~�s�s��%��{*.�bb-#)j�����:W�Ȳ|w~�qn�tW�:���W
o�֜u�ήw����+����G�G��"i��VW�N������+���-v
,�NzP������Й��]��4��s��P�>�	۬V;��B0����5���0�>��f<7.{�k��	#�N�1
�noא�N�2�/f��G�˵�т�Vpݰ��z�;Jޜ��y��u,�Qx�6��R�����㫷XK�L����o����(��v���bk��U&�w\%/R�0�'��΅O~�p���Dn\죕?S�\b��ʸ���9T��jeN��Fv������g�m���;P��9~<��֤��}������֢�<�-}C��e8f�k�iI�F�{�yF�/B���m���0��Y�_[�Q��#��JS�΁Q_V����-���x�ꇱ(N����}�Yި�>�p��^����K�XyA9�DOW��\B1��P�%�ߪ|��\�̫��R��Sܻ]�P���6��P��t���:���<Uz�P���Jˎ�-EݢV�3$��|�g��1��jk�t�/:k�)� ������<�.mC, �^N�
�W�|O��#�nȺx��+Oep��V��|�i�VdLV���;Kt0b%^��W���s�YÕov�b9�xvı�-�wc��&����I���:*��0����:�����iC�>�`�z����v&iĦ�+��y(VD.!nk�imt�O�c�d�yc����"]J�u,�w�X�>�qiY��K��v�ѭ���(�e����;���b�&��l��Xr������֥��*iX��o9DӦ����&p�����kI
�W��I�%9��Tʮ��r�O��g$�[`٫n`�����ڡ��T7�$��ٳ��%	��;��G�;%XYE����G�����y|���������;ϴVS�Ֆ�o��!�Y6�I	zFr�W:���->{ל/��pN��-r���X��r���J��B^pR�0�屉�}|UԻB�ʙ�6P�V��"��43Gj�;õu7x6^7��]���B��Z�ϛ��dr��>C��;!��ת\��l���̅�)��kn�Y�R���s�z����l<��J����K��O�b���a�����l�2��۔/�5�0MG][Db�bti�K���g��<�o1�p�U�	����> ���wkWLz���*�
��e^Ԙ�4�N�.�9ff[�q�����e0�7�'��>�:�K�;oRMh�a<�67���RV�&���:�Ik����m!}�ʰ��IJ�N9�Lj�j92��hIΫ���|v��3�$�5	�;��Y���%c]ԫg �k�`�R둕�)
���.�{���Yjv�ډ��dm�0R�Vl��%Ǿ����E-��z����An���3�6J@�_X���
�&g	t��r"��tC��;�q�e ��$�l_EJ
�Z���r���۹W5T��E+[:��n|�U�W����TDoà�Y���jZ��Y���G+>��[��7|��M��˅Ǚ
7[��[��y;�1u-qMj-�˝ٔ@���V�̘x�����p)�:걺ű�TVc�v�eM+��������]{��V�E�,�� ��U�<w,C��<m�p�z���A��{VV?5�e�V	+�R��V���+�*.1�k�Lav�`�f����Gd�����V�s��7ݝD��]t�ɵ}\:KY5C%̽޴��童�m[{Ӹ���rgC�@P4QC��C湪��"¤�<�*��VG�PPs���i�"T�N�uay��H�S�DF��� ��C�x�^dNl(�E�^d8t��Iap��R(�y;�z	2���U���ӹ�rs��&�F��I%�N\�i�i.z�u���+R���N�q�
nI:��D�.R�)<��P=w4��J�SZy;��d2q݇��^�듒pwOwwD��U�r8�E\����+S	�rs��QM�9�t�]�t7ti�(��c��g��]!:FlwY����gr����:M8��p�ܦX�Y�A�����ww�;.�hvP�DVE��Eܝ���I�#�ⅺu���9n.5�ِf�a���oX��F7Shm��|#䖙g���6,��2��<���5��5n�gj���n�d�+�%09*3�bw�[��:��T����&�C[�ގ��4�4Q훫����lm<V��G޺YG}WM-��R;j�r{��Bcw��i�6	}����o3hBߟ��uW1�d�ӻ�X�}��Q���@M��蒚��H�糐�#�DҦ`v�=U���Y���GRF��&b�;�d�qx&��][��Zb�:�Wªcn��2���yV+R���{Ǯ8�?'�)n�,��+^�����2:����^�Mn���/c��늄����o����h�']�rEӃ�v�՛�o:_R�.9�g�v�XCu�+�mzb�׺��C|����j����gE�ד��1�ގ.(K2��:ldti���F��JUx�\o�;���X)�|n��m�.��$ b+��{ś�i��5�Pea�e��o�o@�/	{����+&͕&��e>P-ާb�u=��q-���1�[���y��
�fq��jU񒌋���d�gN7�Öz+��&���tm���c�,S�����ۤ��Kt�\M&�{W`�Y	T�*V�a�Tb汒T9��s��S1�Ⓔo�u��ŵ�Cy�;�[�{�Vگ"����>�S�]������ �W4�6롾�K��c:VV�v��x&����s-�w/x����U�}}ܐ��1S�V�=���Ld�7�xK E��"川s4�g2E8ۥ��(�7�긒~����z�k���2�n��{�^�i�/��m[�(���"�t���ʫv��r�ck�iY=�!��<��i�g�8W��[&5(+.6.�J��Y�t�;U��-��c��W�g�s��E����o�RJ=��	�!DSא+�R*X�)ϥ�'w�U��T�n�!7[�}��#\���5����:p�"|��K��靫Gd�ʀ��k�w�K����aGk��G�y_7�nB3{�kY�Ұ���p|34����}E���3�xb�d��8�+\>����!�
���#��ǉ�H盽PO]����j�g�o�Q��wo-��P����"��s�h�UJr��1V[Uf��OMF�qjwk~����}��l��0��6�r������:��ͨ���/��K�z�m-��q �u7�/*���<Bފ�=�CY��ߖk�̩�~�*�<V���sjB:��k�'��u㋁�{i��%��a8�V!/mg���{"���yr��d�P�ɝF���h�$la����]&o�W���)"�m���n���G�m���"������p��tmx!Z��´�R�[�蹺w.;>��p�.cf7��(����a@Ϣ��/�x�\k\��=�7��zi1Y{�N��V��?_��!NQe��-��(5dz�+�_\�y0��i����cJ���]������rG.7�����>���WB;RR����;����܎ Cg	<~�ut����1t[��y�N�许��u��@�}��`����u��Z��[̙�)�����U�B�B�"�^��g�j�x�/�gp�J���%z���3�H�'���vږn�gp��[9�׻P�v�<=��L���Yn�ɋ^�o�_�[�y5U�B��yډ���:8 ��|�~��giLYs�k�μ�m��E��I��S�M-�{�ǮϾ&W�@A�V�Q�z|;�L\�W�b��G�^���)���������7�UU��@'-���u�D����_9�VI�^�U�1���P����J-V�����l����ȏd��y�_/W��C�r�C�������ʇ�}zv��YQ1^���B�ί`�*�f�_�a�+���I^uM��y���'kg�X�>��C/����%��>�Y��@��zO�g��w������P�vb��F���>���6oݧ��9�c�G�w����uw���c*1���	�>~�K�IL�c��&�8�U�+��jw����G�㩀%R���b�8�d�D�ݸ�#��*��Ï��U�\G�lI�u-=�0����S�S��LlGY��]�P���unT�]v,�?]>w�U�Ո�]�
�V7�V�@�L+�y����A��do�3h��\��m.Pr���N=�[4K/R�+޽����W~���Z)��n�٘����t�����a�N��Fo��qu �?E'F��=9�z՟Gz5��C�9G�*��6���0&��
��#��/�,�{���}�ɗ�sFO� ��w\�:�q�䳽�L��,
S�}�M> BZs�����V�G�fD�(/�y�H�:�]
�WV�� &h��T�TK/�a�}sZ��=��z�_\�m��z��^��/�p���G�W��4�Ԇ<��wa�U�<��"\��DUH�[(\O\d��Nٖ�O)��4��W<�������{~U�%��LO�n=�U�{L\��AA�ޞ��ߋ���S�a���wf$e�ыr��Ш�Ѳ@xj����L</��\��ݪ�UB���sU���Da���`�@���7 _L)B} )�u�k�����r��2{7��T}��W��4[ /U>���9�9j���U۱֟㳕��W�ukpQ�ф�6,5��5�e���ǙbVN�J�Řĩ*"���z���Ι��P�,lb�^�a�Nա3�][��yq�������!,�����*������1�ޗ���X���j�u�2�{s�Wk_+x�)�;%���9���}xyL��S'��|ik�����=QQ��,[�?��o�t�2��=9˶Z�p�l���8��T����O�<s���}�"S���A��o�rEJV�Ը���ݓ�Lz�)qB�6kM�c}��ߔ� W��jc�W�,M�~5/]Z�*�H��̯�OE�$]�٘vj�*����z���G��;7�������z�Y퓌��|����ح��G��g�h��*��9��j&��r[2��IM[���uC����1ҭ�Z)��wl z⩁}ꇝEt��y��s�<f�����a���i�����F+�S��u^�n|��e{�	eIAm92�I��t3${�_��Pw�~���X�a�O��x!��v���x���q�(��Pr�d��vM{{�CX}���Tzj}�Y����!vΊ���.�0��z \����r ���HR�F�Ƀ,���'`-�#��Lu����u�P,���������}Mh�߲�]mFý-nc=J��N���M z�k��6&fΔ������5��8"�i��un��@G)�48W^�;�����7�����$�1�NŻ�'d��n�!c]�]OGW��Bn�ȸ�z�ni(�,�Y^� \v,�gXGӓ�r=%)���~�3��,�������<�ȫuNH^�������R�8w��3j�y)�|N�~��Bڤl���ۯP
߶��Ϥ�UP�X��~>������-Y�EY��ݔ�@b�m��g�baw�O�=ty�zLz/�X
�[+'�x�(6�Ϡ����V���c��i�涘�)�X��#��#ƣ�����1�]��ǷW��ɟ@Zد��#dúU�a�ϴ�s�vc�":�^	L� �F�mx�Pv�}�q�{,�{T#B����n�V�ϯʺZPݟx� W��g�]����;��]z<�q�p�3�Q�W��o�TGi��c/+n�O����e�=�u.�;�F��XW�s��N�c��)d��m�	]S��o�;ӑY��+ܢ�i�l�s�x�#ך�����"ً�U8w���y���^fn�r��r�i*e#�m�� 4κz-�U� ���*���NE�͗8�*�[�++�0�]7���^6к��ռ�h�,J���f��e��]Ob�3�� ȵ9���Ǜ�b]ں�b�ݎP��o�
w���;wy�%]��/x�O��w�	�-}�"p�xWf�%3��vB�.�Hފ[^����:���n*��H��S�x�_�3��{�k�
�R�DaZr��Mu��ɗ����>��5Z�ޜ��HmQ:��:�	�0O˿f�K��ʗõ�t��$��x�zO������W*<�^�,��	��#_I���R�W�ɏ���Y�}�O����!�G�9��n��Wx�o�tU������Z$6l��vI�=���~��h��P�y�̘�NׅG���<��`���̹1_/	�2�zj�_����w�g(�q�r�rP�pNٻ�x:���x��1�ω�����pv��8�����^P�o{$��>f�&R� ���6��wA�Ο�w�����/"�S�o��>����~ˀ+�{�&�#�x���U�VI�^�U�S*	���ԙ�z+}�����>�/��̇�H
#�@�^�@6=���C��𯴽&^����̫c+�ᾴȞ�ɚJXg��	���]�n�Y��ͫB�^�W�[��Y\�A����y~c³5��U����^�Ѷ�\�5U�Ю�Ǘ%N)H2["��D�ӈ��Jז������w��
�w�������x"Oe��O�P�������ZnvXی�hk7v���0�ֻ�.��͔4q8�w��8��|k���N�Ç�͎�P���v8���S�>���Z�%ފ��:����؍���s���j�<mz`ͽ��<<bo5����,,��Rp�Ȫc*2kL_��� c}R=�, ���)�ɻ����nT\Qb�vvKCj}!{�ܹ�tR U�U	�κB�g|o�}$E�o�������H��޽}�>��=uQ瘇�m �H�*$�F��0+}P�Edς�W�W�<%���ݎ�ў׷���쵖�
�\s�,�{�;2�[7E�1J�W��q�n��]���r_���7��Z�2�gp�%+����ᐧ(����EH}Pe�ؑ��|�i�ޡ^�n�0�۞�,.������",Ͻn���9NO�t���
��������g��n̐E��烼�����-��O7d�j�JӜ�VO��o��kO��1���rb�\]�V�nRfxE��xc�Z��%���@m����6v�W���\��8�.a`�]�a�!�ѺO�1ϔ���!�S3��rW%G���Q#�v�j��)k곰0p�웰���W�����*��A����W��X�W́(:���=��'geכ �a\��eyQ��?G�����[�$��A����_�f|&�A��;~u���U`�l� pM��G��=?D�[�
$�@r��h����C��y��IGo�O}��k�f��rqw��k���=�3�z�ׂ�Vwbs\�O�Q���;~B�Ԅ�φ�����3}1��'Ɠ���|�W��,���z�Y
������W�>�9�t���;p{M��|�3���;�g�鯻ޫ>�^r�n���ƾ��**�r�r���W���g�c}���SL�Q�����"��(?Fj�?��/�D�������]�� ��+�Y\��}�o��m~��S�g�����$h�=5��Ӂ�bc�z:�G:&xa�(<���\�zB�xC�׽��_�����/TL#Ȼ��F#7��V5A���3c�눪`(��7'ɂ�e*��^O��r���m+��'��]O'.����Pm�\����M���ۗEs��29-��jLv��ݍ������ԷK3�3�Wl���+�آ�M��&у���i�<� �9#�%S�|l�u'�Kmru{n�	C����U�>kr�9JN叠��@���6�[▼\�nΧj*��Ν٩Z��S�T��������YB�_�L���c��lR6��G�991��[\5;�q=�����g!WM �Sܾ�]J�u�&��:ér�s*wwY�J�B���s5;���h�*X�JK�\8����B�9�i�VS��ΨgN��%aT^ęǁQ��lu�8�ٲ�.T�(>}\��3v=�_:��cJŧ���2�	�&]��ƻ�\�+y�P�,j�ts6�Cz��K��E]0�ȩVp�K/FЊ��.��	)�{�gq)*���8a�����u]��r�|J])��!�A�����\�=Jm��@MJ���tx��� �s��t4�F&��i�Su靕�^��JF1�����F�Ԑ�[\n����X{ٴ���V���(�U��>ׯf\��fY��{��ni.�R�����g��1u]H*.�R�ΚZk�["[|�V����R��`��W�����5�G�9Ll��vmc:y�ǒ��m�������
K�%����3}�V���C0�c���#�ka�nΤ2����E�W��3���B�JZ�xЭ4K�&�+o���.ɂ|2���hSPfl��HM�LbT�2+xE<���<D|E���j->D��<�ˮ�GoR孑]|n���H��	��zK�|��K5)�^>%i�+��9�Pwۨw�ĳ7�&_n-���|L�a�9NS6���jG"�X�4\r�kp�v��L��h������zq����d�y�ܗ�0�6F�����P��_o�N�>)GJ�����z�҃�c�r,G8����J�3siX8`F�˧W��m�գ]�T�O\52N'��+�t�f7���z�ms\�[vm@n�S7[�Z̭j��G�F�TrE��],��ff�ݔ||q�x�`�5�ē.��Z@{8�y���oXk#��lb�޽WY�0�b�*���w�6��)k���-���h*�5s��N�K��
{��S�).���&b�c]v7���E���t7Q�F�"��� ��Q4�rsf�<�Ǎ̋��8�T�/�L�t<H��v��|u'�kx��"2��y����[�×�����(B����:w3����$�"ir��2�'=̺NBȺ{�9s����8�V�����*Լ�I��I7t�:Bf��)9!�N��͖P�N\k��v�P�)\s���Z8M�Gu�,��KD����nK����=�']�")̉"�(���+��2�J�"L��#�S)�s�y᝜����%OR(.�eI\��w[���s���	�G��	1,"�ѧ�N���&�T.�%u!�s5E�*u�$�s	�hsws����]s��y;��P�N���tӑ�u�H�Nr���4���T��\��,�E���̋	�I�9�t�*��,�v���גb5�_'�R�����=S+�_%v���͠L�)�	f4��U9D�8�y��]1���67��Ϩ��[�Y(�E��zs�2;\����%��u�gЕz��"w=E'61�Z�5芮b�"*.R>L{c'ë�V']�>n_uuk�(W�<}w��+�/|��9�,���f�m�G��@�=���X�ܜ
3��Ӻ��f2�v�>�o����=��p�	'�%uR�����]s�Py�{���np����G�ϙc�ol�
����~�x�<��Q W9d�c ��Rĥ��[3�:��{�g���{�������w�G��{l�V���� EwHUv�)���~[;D׸/�9�	�ncԶ��%��7�@+~ۊ�y^�/�U\�%����ؕ�X��^��� �I�2)?W�`,e*�}F*ר/ND�@�* �A�v�������0t��YkoC���Q�����D)�X�#��<K��w��^��3��{C�ۀ �ϗ���1�U�a�f׸�s�k�🺽^����\�Чr��2��&�v�y�+����0l��h��k&p���>ՉG�Y��؇"�i�ea�F�E��a��lfR.�7wU�y��Ú(ĸ����a'��|���`�zv�xc�o���7�=�D�N�FǪ|*<���Ί;s�x��ʬ7_�Oy���Y����n�<� �m��Ǎ���ſQ��~r8�Ǫ��7��d�B���t�w>��_Џ�Λ��_r�&�񿙌�K}Q5�.t��x��S�P�v�j�gФސn�^o�'�t�;��1z�3��^���;�Á��s
��Ι�&O6�&�Vz�鷤��f�S1���|.#&u�ɟ"�D����<��Ow�y���ߧ�[؝�B�yX��*��7���y����n#&c�{^l�c6z\����*ޞ�������ʔ<9Np��@�6�j	���*�+����"�ǒ�ӹ{�
���vRf����w+�z�~
r�/�n@@Y ���;�\�]���x6���^��F�&<���L�>����tU��q�.O��`�uM�tB��������[5��le|������j�;LW���)����D8�T����gW]:��>���9b�
�i�pf&���=����z�IKj�w;]�R�z��VkS#4���8F�%t���p�t��#�S^�=A5���nv�9-���XW��+4�{�[˱���-�t×8�+6�':Da�{�J��P�1�~X8J'l�g}���U�3ω���5�ZyʏMVlyv��=���8<��:�������>�b�����G�J��y��Ȩ�+�Ъt
��\_yߍ���^DI�x��5��5�/O�����#/1���r=z���z�O�5@p�G�o�O���@����ǰ�ݨw�mx(�w����a��ϊ��f��B��.�f���O�P�,� H��Ρi:X�+ݾ�Wt4���g�;�agL���'���_�g ��^����s$��_{�Y�h�z�ɠ+�/�.��땧�,V��#}7��P'���js�o�'���6}7�򤩜�G��^�جSÊ���ʯ����|o\����{o��&����&q�N�_�\�l?D���|�m���D�'#u�.�>���Y�;ҵ�W��@ҹ���Wkt�]�w���z<��G����;�3���P�7l"0.+}p�0�"_��xz��/el�x���ܨ���T�2�;wLc��:HpɓV�7�O�*`�m�"ۍm�.��څ�E)��8�Nz�S[�λ[���m��Eԩ"Vm�p�`�������cYz���g'��on��/g#���B���#����A�uj�n9�g�ߘЭ�F|���bV�t@7���^�1[�����!���aTF���)�Z}5�cЧ(�p�Hl���Uo��ѕ��V����#}�W1����E����]L=;��޷p�Y��Ź+��%�^�����f�A������g}YX8���zx��[�59b(��{���D��^]�	�7��F
f~/e�%vN`(:��w�%�K̫쬿n�eS>9(r�xf�Ƌr&Gz�Sd��҃V�W����j������nS�hvzG�ᠳ�����^ +��E�Y�UGW��B�d]�}��Z�9��~</�¤�zL�^�����w (������C�Y�����u8��E�`����ke�2t1�UP�Q����9�I�x{ځ��Ǘ���ڥ��P?x�c�r��d�~y���aߵ��ge��^��R�|��ҧ��������fy�¹x�>� ͣ{@>���=���͝��n��;����MI����	PF9g@n�s{E^jF����G���ѹ��>[a�&)�elR��ط'bb#-ٶ6u�ӥf�`�lGB�7�;K�����`_���"�L	���.'*^W���g3�:�������c�f|��W��=��k%�>x+��O�a�aѩ��~��Ѫ@�T��hx���z���衞���Oc�P��"���p��G�&pa鸢�����o�gG7�������n����}3�ި�SȾ��G��V�r��<�������~ȵQ���(^�=�\,%عu��#�}LR<�T*�f��n7�,��&�v/׹��uT��>����p<���"��Lǰ�v�UpBӞ�q��G��6���I����f��y����K�G��*��-�,w����b��Z�k�2�K>����>�W�n����ǂ6&:,��D��R<
��DY|^\^%r��T}����6=9<�������~��j=c$�@K&A��`G�^rǞ�5aZ�~��=>�c4׷j���N�֝ǃ����\���GŁ*i�%��w޽�kb�FR�A��H�=�n��<�5����5Vm�cel�� ��5^%0&��Rt4cr��|�77+�ګ�W�k���&��T��{��>5���#N�Õ���E[�����'6v�gb���S���sA>�O���H��~.K�H}�Q5�ȇ�D_������}G�jX� ��d/���L:���^��7��Un(N���gz�-w�(0E��ux���>F�L{.:�K����5�����B�%��H�F��Ͷ,ߴ�;}qY��k<4�=�V���	Ax�#ԕfy��=灚�j<�Й��bK���fװi%�,�_{�B*��!$e}�E���xn3��f���I��F�R���ü��'��H=^����x��0<fߨ�O+���PGrf�i��e����
��=3Y�ew�a��E��UB��3�ip6��+�~6�g�o�'��ߚ�#���c���&��~
zװj�ў�2kJ���L^��i��uz{ņ-���q>C�n(LӮ[�wޚ>ㄮ>������cc&u����/:d`��������fU��}�'�N�P�i�۫�["��Ii!�����[�ө�&o&c�q����r��B��wtgה�J*	K��k�5��U<���;�*]�&�O��F���3�������to+ij=\�&*�����ܰ�9�[��\�C��vc�������ʜ�J�\�UӞJ�����s^V=��ޱ�=����#��t���ޡD��(IP��W�+��������'�ݾ��D�����\z{�b��W=��xW*�˿��nn	�0��d{�=y4�����h�z�Nx��L{�Y�1��������'E��F��ezK�$6w��s���X����oyx碦D��@���2W���/N׃�x�O��tGn���1��o�������z�ǣ�O�l��e: ˝�j��p�;*`3�}3��|�Vߝ�]��k�lϐ�.��פ�*Ѳa�*J��>g�w�.�|K�{���Nv����IH9>E�?{�p�x��u�o�50��U��d��Wn�x���O����
�Bb{�x�r����@� R�z�
��&W)�����r�S;�f�>�������Ҫ���+�1;�����ϗ��>y�**}�ݔ������rr}�x�ZX��p6������߇D)�����L{�4�t��]:����xj�|��q�]r��e�W.�sb�9������ġ�.��{P\*�3�}I���ݻOf^�t{�4	�����VQB3n!�31fs[e�Y���k8����3DP�L,asW4�/����|}�%����+J�
Ӭ����X��������;0������W��	.��ٗ>~a\3�h�ζ�[��ө埌�\���G����\��b�x\�ǳ�_�M���6��g�Z����f��3�7�a�M3��|�z+g���L�g���
�}H{*a�'���x%ohR�(3�a�[ꄰ��T�t����~�>s:<!b��s�� �Z��rY���
wPfs��>��67i��az@�����7�G#�0�L+�L���9|o�^��UYe�o'��~�m�׹@�d�UHU.�\ǃ���r����q��]L[�#"'��^���DL�@�H����B�вd��u�,��b3.lmD�GEB�������{��~S!~��q�ܳP��'�ق�ٟ��c�\s0JO__���=�ճ)(T�Lx����(���;�=�U��%��@xT�Ok��ՙ~�Gt*=/5���N��$�;�B��u��CP-�Jօa�+g�[�يT���(X�,S�CF��!]�6)F��MӖ��& s:���4傦Ζ���u�b�t�5�v���M-��5�����Ln��>�i<�Mx �����{&�c�>B��S�"���W+���ͭ�QǴ�|^�P�u�4iz@^7
����Q�>'#�g�����C��ݬ�j7�X��sQ�X6�S3��3;���B���>��~�>5	�x{�(O�0�� \(�����:�z����5g�:��g���W�<sf�y�1~1ܠ�r��ޙ���؋�cȞ7��2}��5�����`Fͭ�>�W���^=��)�n���	��(��]�'�0�0���Uq_�:�%u����:�ǯg�ٓz<W�F�^�2�3c�τ[�8B[Eȉ�zn���&be���nw�=`�> w��w�#Ȼ�u��x�����^���k�br/��ŗbA^�`M�p��}�p���Ñ��T�7�m^�k����jK�,ҽ����SR�蒂ٟ'�s�X�c�>����U5�wPV�?]�Z+Kh���*�ME⊁W��Y��#��d�-Vm��i���K԰�+A��yﮬ�e>`mb@9|�Z�u��ls��t�X�����:R�1ًsT�.�cˮ/;� �_E�U�&zˤ8P��\]���sr'�g��;7Hfc�[ u��w(uFe1	G��5]�b'�4�/9�����\y�/�޿dxdt�������lET�
�ꊲ���g���+�]�3�s��_���6Ώ+{dxW��w \{�4�v	VMёt���f����-o�x�f�/{��%��M�zxc���?S�rE����nm����:0t�A{�r���cў��������aY~1�ɞ,����:� ��n�mV/
>�7&��|�o<�=�Q�lܡ��v̊����`,e-�p��LL.��v'ʛ��f�R��~�n����0Q�50���[����=���i�#$�]��Zs�n��X�Ei|��~�n � ���z|����Y��׸�9�fz:��,�/��X�G��VW�s2�����޻p�|)��#n�:va����L��.��
��vk:�W�O���G��� �N���Nx�S�bߨ�O+���q���Dv��#�'�����{��jw�(�gJѡv�yV:mi�gu���nXb6�eЛ�X�h�b�:�*�$���;�b��b��ONGoc�݌��p��2�30n7�1�[[ĺPh}tЬlRi�p��uq�gu�j�E�8d�r�ZVL��U��_f�X�,��r	{g�oZ3���bF�&�Anz�u�]0��o�p��B޷����Me�td�28��{Y��#8��h���'SP������")p��gN窧AN��c3��^P"��:����u憱�V<��׾9#�ƈJ صy��&X���z��ΡYR���=]Ώ]>�����om��X�����B��S]pvX�GYc�4)66N��L�5�_H��5t]\���j���:E��]:P�{��� 4����5>ՙ��wse۱Z���AK	x�S���5�T�EZ�$��j4���1u-*$Dw%#S�^��U�]�t��u�9cl����h&�(e��K��K�*���ɹR�wH:���W�^7�P�%�Ұ�:Ȼi�����ƲU�ŋ�4/(�7nM��J��"���禭�m�ڟTΉu�1�d�ݡ1�Ue�5�g��1%�`�ra�Ų��8����4u�)Ήq����wƬ�ϯfp���pcl����;;��u�-56����1Y­f3��M.wb4�Q݃��6`sU�p�V��f�5%
n4�r������9����㴺������~�s��˫w[�۬k�%t5#��rӪXy�r�'y���	�\PC�bY1��Eذ�g-!+�p��q�����ã��ƣ�su(S+��)�u�é����-��+[��S6�r�U[������f��k������m�]ïJ���lc��(Ұ54�bi-/�u�눀x�*t�1���}jP�`��,3�%��%���T�!��3�]�����N�t��M�
)��J��̯��>�l�ĺ�����7^���淕�7z�d.�Dʹȩpl7|+X�b �+2���[Zя92��+s��m���O��N�>�t�����m�e�Iމ]b+��V��i�2q=٣UbqZ+9���K(�����)����Dr����ȯR�;�fz�gW}ó�<���i�S+��ov��(N|�W=}��|/�ϥ��:9vRO�u"P ��F�L��$N㻧���3�u)�Uc�r7q<�L�w2�	:Z����sú�ʕ&\.H�;LOw+�uJtZ���*rr�*�吐*!isP��Y&�K�u�)����9J.���[�U��VX���R�Y�2��Վt�h+(�
P����#��^%��(�UbiWnF�YFf���DDē�L�IE+�.VL�	)+w	�Z��	�/q�ꊸ���w74�S�ҵ#���Z�7q
r�;��(��W1�E��*-0wYwQ!ɮ�@��k��*�^m�)2D�J5(3	�-k���9�.��:m���%i���*��J)���}��^��'��.+��T��J�=��B��u�zfj�6#�ՐD�[���i��:�X���i�zN����{�׏�.�F@���o)"��o�ƣq즻����0�B+�=�x�k���!�"*�ʌ��댙�Lk!��#�q��Lt���32iQ��\���f�c3>�j�t���=�NN�U���c	�{��/#�Fn��$�=��z���\���[�DUﮛ�>Fq�)�S[����䙸ɘ�_u:�C
M{1��9u�,{�d�=�.�ͺ�A��8�g�B��v\MB�?RT�)��a����W���OG�$kT¯�Wq��,.��q�ޯW�}*��/`���"��ǰV�<� ���/}��9��y���0�}[���\}���u�W��Bb���������S��C��0^���J
�ʽڅq;LTx�I�q	��hl;��d��r�7��D�|��2 C�T�:�'l���O�������59�N\�;n����5ǀ~~܃Qnk�@�BZ7��T���o�|;�LZ�;=�Jz����*==�JW'De[��XUta^��.�'h�ճ�c����6���i�ۯ�j=�S����#�<�Z��r^n�r�� 8���s�1�]������qk7g/'7��U��@s����3X
dW#�5��I6=ٮ6s�'9'�O��\^w�p
�#Ʀ_ʾu��=+��3<m�ڕϣ��޺5Y,`�1?r��?H֦�{����@����W�6=��i�y5x��^���^}��eG�k��S'ƙ�>5}w"O��$-�mou緄M��V�>\�>��Q�~�Z=q���z|<MD �oz���B���L�7]�d.��wb��V�޾�$���t'���E��>Ү2|+N�3��Ł0�@����`Bvr!粟��{�4ϣ_TM}���ʄ흇Rp�eR�t�E���r�������T�S�>�B� �԰��Y�tR�7d��U	��7&w��c�#'����V�ut��^�)t���C�U�(�{"T��c�D�r	����W�r��7�U��l��;��/H]9x�.R��yE���OյC}�9S�S_��ή?�	���
��	���U�7��atj��)�ÉJ�~���?��%�U���Qi�v�_!ߟ���-;�z� ��wCT��]�X�sv��|ixo�V�R'-Ӭ��\ܽa�e�fb=VY��c]M�]�'�=�'V�PsXʔ��5kT����lc�����R୸�}�A#	��N �u�5�AR۪���]0,ǃ��;��A3�b��a\Uhة`�z����u��t��t�,\A�-�X{uR&	�,�����͎�|'�'xM.���S�,y�鿞��UA�L�/>e|`����/i�%q̆x�J���緔g��{��Q{JO����˂�^�\!��@zzn����L�w��H�q�g��A�Yl�i<�� 9����� j���=g��Ud��ٮ=~cF{�=^����O����	�]�4j5z��G��������kڹɢ/O���[���%eN71k&�ܟx�F�ft1�U}1��'Ű�ұ�0�w\�H���v�R�'���?����6�'t՜��k���F�c���o�U�@����O�y:r���/g��Ȩ�6�\�Cˌ�qC4�g����Q���~�������޹��'��"�<���]�>�H÷3�}u�y�� N�ڑ�롥��\-;�.P6 !Q�Z2�� nf����Pe���/۾��fң@�����igVꥼu'�J��ɼ��DGT�]R�^���-r�.>������������1׏���]~q���g���<0��tnG.�:�V��p�^%S�J�K=Cx�Կ���.;������_�(�g�Ij;�ro�� o�j���wU�_:�o�2�W�s>�9duo��9Ru��Ѿ�nn�o��z��A�����<��L	����ϑc	�ld�ud�CԸ}�ӼX\a͏tˑs~�>�/������n�1��)���b�=E�}g�]�J~���.����sB=�T��������5�_�<1N
�c$�6O@[2G�^�{=){pEfmw�ߟ�1�Qu�|�q�Wl�
��n�_��x�8�Q�$Y3�?o�����/W����#B+۵��Ǐ�A���������uNH�HPwpf/H���'�c�\�H�s�X>g0�+F{��Q߉~.M���O�z+����Z�թ̍���uP��7,e�b$����ǲc*
���a�
���A>Nr@Rx�k3_����:���8�׽��p�ڴIO]�k��Y�B���͸;
���0��V�<zV+p�2�o���D��TZg���g{3��#�����Ʃ39�Z9�z�i�HwI�X��4c5����CȶA��.�mB�0��I�WOI��<�<�}&6T��S.n��ä����c�J�Up}{l�V�?Fz�������9�`[P��B�������0�3k�FVoS�˶q���k;���4OW�Idk���ު�O��	#+Ί:va���Nz%�v}�/q�9�;��XoG�� 61[���P�A��N;���6�v��q�W-�Bψ�>�\������]���M�p6�P��ߍ�ơo�%ex33]Y�m3��N������w��3�{�;鋍r��#�z��mw���3j��>���5Z�6}�w�l�;�'����z�=?\��3��L��� ��B3����t��p��<԰�=t�T�TbyR#SتD��ӱT���1^)����q��}��/Ѵ�B��Si��J�nj��>u��H�$��5
Ti9q>vʫ���c�[�7#�Ǹ���Qʻ���Z=�c{����9E��6KsR=�.�t��xȊ���Ilve^�3��������Q�9�X�yW�_�&�q�ö��
��9l1��&���r���z�!���8�e_��N�MJ��QOiy�uoU�C��J"�)��YjQ���x�U#��#�º�z._��&�0��������@����Ș��n�#�{���q:��I�@�#Y�3��L�'�����aL�׻P�'i����Ɨ����R�//��>���ތYd[�RcaxO��0a�C���œ�n�����^���;ʋ~]�S���FN�%��������U̐/���ʀ������ݝ��"�d^"s_�s�>s���d2�©����\j<�*S�w�S:~j��q���w]��=��g}r}��U�!�H1̟~��!u]�x��̀��ëQ<��ty�/+�˻�M�gmG�#6�4=&v2���T��d���|u��+�y9R��v!mvzr�!{�ʅ����Z���ǉ���<��2������}u߳D����=��n�Zч;�����Ug�����&�*�h(z^�=3�ờ�>.��T���Q]D�{/�j�n$��敖�3�2���5�֏�W����1��Z>㹶��ك4Zb�}�z��|��Fu�$�>��"��M3�B��L$���o+"���Q�c�����)}%�ѽ��U��p��wӁa�;(q{��t�P�ó����ts���S]w�F�a,�<��s�t�E#C���o��g�Z��@5[��T�ް�i�ߗ�G-/-��p���Y�#�������iA�wP�9��щ�C�d��i��̉�W\��� ^�G��[7�>Ǆ.�T�B:�n%�C���>��=�+�k��~����Z�?�x���A���,�����t�L��s.��Dr��]VU_�wo���NdixHH��d�g��Q1����(%λ�T��';�������w�픮s�wgнn�����,dٸ%�$\�,_�\�w1�;eǯ�{��m;�s��x�xO��n��~�n�2 px�1/i�۱ T�g�����9���{�l�#eρ��;��=�U��%�Ā��=m<I��xov��q襕�Y��1�5�¼/L�G������{�`T[�\��lj��yJ��u��j�{�]�+�-6\ܞ�i�/
�a�z�^���������<}�R�_,���q���slE�
r���G�[ڿY��+�8xAD���sUG W]Z��C��kv�Y�Ű�������Z���� m�h��;v�SJ�T3!d��ޤn.�.��MxG�|N_���F*㲰+���5�ƙ�{UT>S'�"�����P�3�:�#էж��_�D���Y�p�O�x��ѓ�l`��c\�k��FK��C\�wz�z0yK�Ys_{�Bi<�� &'�O90�c+�P�٭'`y�H�~�k;#�}�~#�� �gU�����Q�{^���v'p��F��Vqtlj���C)w��z;:UF�}}Q��:a��ÜK��+�vkE��Q�P(f#�1Ѩ�p�ܔ�z,��2�-���J�)V}Cx�K�ɿ�+�}mT�M=XǢ��T1�:X����X���H�͆]S��~ɖb��9�2;},!�ǵ{�Kk5��s5�޻�>ھ��~�,��uL��ͪ`MO"*.|��1ꌟ�˧!GQs�5��x�	r�����%{ޜ��=����H���Զ@��/W{w�4\^�м��;�1�'�:}�Ϥ��z���8�&@�)M�;i���n��<������#p�����u�kN�>��ŷOGf4r�s���ox�}�LM��Mѕ�U����:��7v����jF�뺝��l��'Ȋ�8(�%xzeoj�Ġi����%����z��wǣ�����]g��R��6����V�a��_�O�C�%�j_G�u[�����+�d�\ �ȣƽ��gg�=Ӡ���ǃ��m��.�0"b��u\ϫ�ԑ�h��Y�*@1���n��+{�[2����>T���m���8�`j��[ys$Z�hѩcQ ��#c�}���T*��9VX��[�pk��;R=�j����=��O���*|���!V�x|:Oi��1����^fx�23�zh�GLd7#Ǚ��p{py�6)z|*�]|�0�8TĿ9���]���y��%(�ڏ	�u�q
d�*!ω�G�T"����FTy�Gr��wK��7��k�ۇGٳQyU�����@	U��Nx�����$'�����d�� ]"�{ۖ/��&��JևRr���3e �DaP2��	���6�g�J]�r�E�`�g�^���͟R�.��q���9.pjȊ�2�kK�w��3Q�G�]@"`�'�O��N�0��@�܌��(�}Ys�L�����葯hڍZ��y��u���Ӿ�Κs��P��w:�]ʅK���q�����SU_Ƨ_o5��������rg<�ȅX%i�[�)Gn�v���7$�]oYu������|�3�7�~�'�6lت�7=����L��-/{�o�s�{ټ꽡��G���B�^7�}q��H�yIiu%�[[�ԫ�Q_+?c�7�s��H!Q�¾´�R�P��1Nq��L�'����97�1�������E����0��׾�W�)�5����Q�ޯW��NQG��F�3c��ڳ'��x���0�I��%��T\�^\z�)�[��Wx�o�tOJ���:�J�=�'��d��l��Dg6�D�>�ʽڅ���EW�sF]��_�������h�=9������T���xO�Dw��2�CNٻ�x8��2�v�-��閜*�H�L�zb�D�s�
��5�$	\��D׭���vΛy�-�/O�yEP��	��>'�Y�jz���S�+�������vL<��9��۾y����d��iu�� ��������{� ��<�DMHQ�wNM�׏F���A��C�5a���d�>��ܮ�w��rZ�	7oK�z��q֝}����f1Y��Rd�҈ʂś�\k���"�f1�p�Szo{_@�ՔE)�\��V.�Uˮ�M�H�Z�F�$�ϵ��
�%[݈��T��A6�#�b�oV[�ώ���9ՠ�i6z`�r�s��̨����\v�-_ r�����Z�;�e�wEC�)��\�ZK����7C
��{ޟe인�[[.Pĥ�N��)��K�6��ֳ�s7(���$"ѐa��w��^�ۊ�� ����+n�֫�#�RT4��k��Y�Q�����!SML�t��ff�:a��Z� ��)�=soUL-�ΥՊ봿�/3,4Ϧu�[hGC���EP��t�0��ccL�R��u��m�nMW�oy�����;)t
dU��_a$�S9±|~�{-2ݶ������)���U�-�i[��˩���ltwCA��,.�,��Ũ�V�N������`[7�2-��:y�;�4J��]��������l:�Z-///k�Շ������k���0@����8����T�M�'6P�h��E+R����e�v�ey<m�8#�?F�7��b�ec�[٫�Eߥ{d���H�`��w:�?L�5�$�-q��i`U'؎oZ쿱�x^ӕ�2��Ϫ�y$,/��W`6�Ζu��b�:8��l�1�Tۘ�Y�F���Rd��p��u����Wب�\�m1�j��{��6���+'g V�u�Q8�R�	��N��U1m��I%]�Bͨܝ9!�y;��5i�s#QR$ԇ~�?�-?;>�#^s�����!+�wGy�Ly�Ԋ��3#R*��:�έwb���J7�8�7���/nRڋ�z�;GG[�iNsQ}Y��+��tl�\���
�N��T:��V�8�>4Fa{v؋5v{97!���v�_R:'�8���H<g�a�4������le;��L�b��M��Y�}x4�y��{%���4L]�t5!�W�K����26g7�����l#*wK�)��+1�p/��:�of�)s����ԏe�������<2��0�������x0���*���XC���l���>�XE�j�ԕ&����$Bj���J3����o�R���⮷K�f�'js�/�����Ҷ�4�u�>�`d+^��B�� �^��'5M�t��v�bhk���ljڹ�o�f�Qv�X�p![�����9o'�.m�՜�	��/8���Ӭ�������6�A&��Rn�������#���w�_��}��{�]-f�ID\YZ�*�*�|{���#"�B��Q��NZ�w9Qz�L�*�*�OS�(�+R�����,��BYb܋�/K�Y��r"u��t2-����# ��;�"��iS�Ny3-R��L�̺D���6\,��.^e��B*D���ɮˮxr�#nBꢵ2�:vkSl֖DK��8Fe2(��QPE��Q�$.��]�Һ��*�*��q ��"��ȧ:d��%\�2��e�B��T( Ԋ�u0Ud�H����"��:�PJ"�Y�D�F-&�:t�9V,EY�-@�ʼ��Hu.W�{�7����zʵ���A�6nt���!=�tn"�.Y�>���;���쾢]��z�P�/O8�6�kq�j��opG�A(P�?�n�u����3YP�z�X�2|c��}��qS���Bvk��5���W�wp�3�aᯧ%����vrzp1�V��z���q��<D3��9���i�>�ف1�]��I��F)ڋ��iW>����M�`Gnc��2+2��ީ�9J`'8�#ز��*�\�g����3�)��k /�t�#7�c��݃�wt���x0���M��J�5����E Q;�U	�{8�.��W�7�=�-��(/t����q�.���3愠�Х2�$�ϭ(5�1��^
>3�Kn��ɖ�GZ��GQ�Ŗ�iTau������]�;��/G����;g�
�����YC�yW<�K�S;�-���=��6J�+�u��ni��@l�R)�=�K���{s�j�}���B�����Pu��琐��jT���8}�u��+�X�:%�pJn�D��,Ys���u#��3kj�+�$��n��]~>�����xs|�i�"��/_ ���D ,n������n�RU3&q�ڴz�:�G�ŷ�8�K��we��I�b���@nV$ep�P�:U��PY�v�9Fw5����9U}���{k��|���J��G��wy�P��'̈o�__�����yFG�$�^�o��9�2
�=�*O��.|'^���nD�����;��A۾����Nzc�f�;*!�O�-�Da�^Q| Oʀ��ˏ���8�VW&⳯����@�¸���Y&�^�ʐa���h��OZN����;ػ!�^�������u������
�=^[,i��,z�T;����z�w��Ǿ�t�uLyD��~���O�x��g0б�3��6�c���Ş�[�ў�����\�鯼�מ_�_��'�\�C���-�"H�����:�S�>eW^T� W��p�<�|$d'��~x+���F�9ʂ����練�P�G�N�\b��z�}1�΀�S~>�c�����hf��Ϝ+���]�V��gN���$<&[u����}g�7��K���TL#Ȼ�u�W�c��H�9U�{�~��E����%�V)_^�g����f�k����z�ۢ�;���b��O�� 2��Ns�N�v�S���(�G3��tqp#&�/��5ֻZ.�+�����T
YPk鬋���MR6iVu�)��c��ږ}�ћ�߀_M�+�����W�73��� �w5]�5��*�����ݨ�{(������HAf�0(�#"�ȱy3ob⑵�V���H�yʯ!l��k�p����sS�IF1/
vl�l�zKd	������oH���%�=�KQ�HGiѿE�Sg��1_��xLz�X���P�NmE��z*�{=q,F�b��򢾳��Ʌ�u�P��Oq�����J�{ޯ��j��$�֣�w�_�|H2n(�JJ�Qf5��j������:�x3�g�M��]��璂���<B,q�?t�~�8���9�5�ǩmR!�1�<�m>�}�T���}
���w^�.T4E/!HNّ^^��ŷ��yKgoW{d8�9&<ڠ\�>����e�n��b��>�f�\=��|:N-��ڽu}�cw|�v��#+ê>SD�JC��~��\懽���`��n	�]�S_���y��&�OJ�݉)?[#hX�싨���u�WU��0�_$����r��9�������*�S��[<�*�T1���.uC�wO[�h�S/�STv�>�;h٫ٕu��q�g`�&��P�e�����q���.7�zx��bc����,��^'ֽT"�t�?1$e �,��z&�y��i�g�l?��U�Զ�Ϭ��uj�W?Ξ�s�#Ɵ���t��s[أG&��)���gHg.Q������ۅd���v4�Qʀ�^��n�@��N�;J��}�Q/����B�<t_�>�	eSY5��;�d3��[D�zi��{¹Pˁ'���f��2��Λ���y�f�튨ss�,a:���xN�ג��νS��~�7�2'���U<˅Wұ�zZ���H�:�7�t�,�&��X�,j+{<x�Y�>�&c�q���X�+NZT��Wh1�
p;����Q.�z=������,�4����1K�}jW��\k\¨�]���T�]1c����Ö�b�[�g/�ܻ��x���ޛ%����JW��x��&�
u����+$��K���OK�g,���^[���%��7)��� x8h]�Jf�v�S�����q��!{p�x�PTJIh?B�R�k[��������d�ؓk�M�2��ym��i0(|�B��u4���Z�Э���սյ2�<���L)��Y������zK��:-oV&�T��]2����;M�G6<�:ܶdq�V[�ôr��ӈ�o����jpo�ꜘ���>f��������F��wn����78������u�e�TO����+�� �[�*Ѹ&t�^1ל�X�9�]�;���1\Q,(�M"<B��>�� j��������9���X�,��?/}^��Ǵ����
���z����z��x���yp�=ܽ���k�/oWp�a��Q�ͯ
��/I�ʇ�_u�0�>;��}}\�D��ŝ[�L��2�9�E�Lv��~��*��ic�֖�}~��|dG��nly_�H���1��~RI�7��nv���iW>�Y����Q��m��봷�e@��遟B�񥾨�Ǘ�>7�`)>�޵�5���'�~���j��|ԁ���f�S J�������W���<ab�A7d�x�黷=�s�u�(^����]!y3�������
](;�u��w�FBzi�^�~�1���2�s�q˻���m>ZZ��۩pV�(5QS��]q-����6�ʲX�pI����Y�0�d�x�}(Z�Ω6wv�l�\�nt8�ޭx�-�H��gG�w>\�����=�Yoy`z�P�k�f�����o���w����#d��/�0���lX�{/�^_�����K{�g7�>�Egސ%ў)C�]>t?�xʲ��3<��s�o��_ �v��&�ߧq�r�q�U��3�9E�{$6o��R=Q.��\ǃ��}����ˉ��s���V��1�u���+޿\{�.O��Z=���I=��Μ;��"���C܄�h~��OՕ��D����*S�#������nG�O�x+�窞��:C�k�U{�R��d��� �:��|��>�u�Ǖ��{�.
�Wt�d�x�����b�.� B�^�S>��τ��O�|)l�6O���� �n+�/fL߮����껮���Y��GTA���@T�$�<>
8�4�L:�Q�UW���������N�a� ǉ[
�������+����*4������N�n�"Lj�Т�g�xIُD.�(�/Ux{>j*=�K8-����OW�����y�i�>�;>�MtU���q����g��,��8�>z����a�/��׺�0c>n�>��n�qئ��2:�Ax�ߟ4� �hƬn�7�M'Y�k1�<���$uη*�����������ۓ���LR����c?~�g�b�P)Ϗ��2'���y�1�����yz;���/{2vokG>��o����8ppǲ��(�����W��O+����]���ݠ\,��3�Uy����z�}u��=G�T�������@L#^>�����uxGG�&r<刪\:gw{�x���[E��U�J���3.g=8Etφ�z�Q�\���W�)������v��h꾭��ԣ�!��l z������=-/u�7��3}��ѧM��������LǺ���d�rJ�+"=�2B7�DQ�,K�����,���<�^�ӍK�n����j�f�Hn*��8?#4���9���q>\@����|:�|"~��ќ[:����_�<1N
�����v��Yw�S��0��G�1�}��0���J�RF4y'�G�_�\�u���^Ê�;i�z�z��cIGā�&�� /K .=a3�ه�;^���{މ{-�wb�vEN	��'U��km"��)> �{�	\�]Q4N_j|�ֹw.��)�����.�٦�Fd!Z��!��Gc��.1v����dpn(E�T`�k�l��b�c᝟@Ԭo-&/G_��F�p^��"��9"�z��U� ʜ
��aY�zc�x��(�}���T�DN32y�{�qV�$9�h�,ZR��dW��ǎ݆��ܲS^G=T}��WO��d/J�����@�μLWҧ���y}[�び�Pǝn{�\�}����X����SD�_r���H�Nhz�u���b����hȮ�@��R�z�"�pǳe��S��mC>�S%�ω��2!G�]xg��V� ���>�����uv�j=���;ɛ9_�M�R b�Tg���J����uU �T�;Y*�ߔI�n�xZ#M�:�7��;(e�m��L����M�p7��j��ǤG�d&.r�����Q�1�V����\�kh��Y��e�Q�Z^����!������d�{T��o,��V�#���u�j����'�6lڨss�,Y���^��<:��g�Ϝ�e�#p��]����ʚڌI�B�W���CӫK���?~N�T�T�������2ka�#�r�V���N+s�;���"/c�N���=�[�s�u�ae�"�(�x����1t�֯��ײ q,��3{��e�\̙���ut*8�36�O����.Uz�bruw�\��|͓�ׂ��Ҹ�}��w�/δ{#�=��f�9|��V6��5P<0�����t	�n���J�0����r�㨰�F��0�B19W�<�P[�Ez#j�F�܁�Y �)J�T\���
c]n�;�lԉ����{������yEp�^��IQd�����S `��^Jf��^��{�gS�*�\zgA�_�r����L�~�!۪rbׄ��������{�-||]a��ѯ���3��>'a9��˃�~�\�@h�l�|��'W�c��(+X��m���=,�*#�4��H^��S�=�>������M>=7D׻�nϾ�S��N�MB>�꾦4R�1=�>5��p��{�xS��X9��L�}�.���_��xV���ͯ
����ʇ�Q�tũ���-��΍��1x�Aӷ3�{)���IK�I���zp:����Č� ex-�W1ڄlTZ�����λc:�)�rx��q����9��,��or��x�(�k��Y��]�{�*�!X&=�Lr@����K�f����/os����j����֒�Wӻ_P&q�Ʒw����������������$���F��~�
���7���X�W�:=�X��F��0/�ߦ񥾨�w_5BQ��qn���{�������~�w������l������#�}L ���M��J�7��[��V����G�g{���J�Ts5���&w���wR#+7����;�z��`r�L�)מcӝ�j����n�)�6��]�xTE��^9���{)Ė�K^���+W���h�U�ſe{#ޠ)��Y;XJ�LT���#�z6�B�e쩞�#[~�C�x��έ߆t�n=�Cd"ͪ���F<�O�m���ͮ͝����1�#����j��zM��z�ï�,�����w�T&^k�Ԧ��h�({��a�߫+\*��/J.Fs0GC�3q�|=�B�ϨD�������G��u_�� >7z&��0�T�w�}_���^I�9���c�������O��IPUW��2"���$��UP|;ЗU!�_Hb,>D�������h��q�q����}���m��>x<{88<b0�{@61��0`�?�ϧ�>w���҈�+8�{�BRUT�#8� �6F�+�~�}�w0r�>�B�Z﹊с��8\��[��Nx�~_�{�D���~�y~}���m�?5{�f9������:UT�a ?��@�V�/��|�������J�����9���$I��UPp��?b���"ʣO(�^=����)����kH���g��B�7<�{����4.9��r ȱAU1�i2���M��ª�냍�r""��b"��%	��|#4��ҥṪdK���U6�hw��ֻ��پ�� \��������%n��h���]�<�脇��N҄���I3�eEUA�[.���C�4�?�;_ڍ���k�٣�IF�g��ȷGX�"*�*�#� ��L��[Ǐy�7�J�"P@6<ǣèb��hT0�"�$�d;�xH���Py��>���A�{D�������~��7���`?py!c��T �X�H!���B>Fi��0�Ԕ*^@��xX<������~�}t�a?��6<�;�Q��CB �Lo+R�(���UU�׼�;�ܛ�UT����`X��k|�{�_�#V�0>&�p�Z�B�.;�;���t��pG�./fQ	����ħ�q�x~>�PUT������V#�	�Pyw{��P���+�T-�1�C�臡�܏�yx�Z�A��v�jB�R�ȔI�Ü�`h%#����z�r�+n@b@�|7Dxz��
���t�*"����Czx�~��ОL;oI ׈�OD俪ӻ�r$������*��?�
@��D�O��5����UUA�Cq��`�;/OL���b�+�V�s�ʔ�`4 � ��"�f�[[��.�p� }ް