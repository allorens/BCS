BZh91AY&SY9��S��_�pyc����߰����  a����  $    D ( �� �B�� EP��          o���}jP  zf}�PP �@PP	  PP�Rs���OOGM4gw`.n��ۖ�����'Zu�**�#�N��u@��Ӻ�;j�f���ݝ/o�I;2�ӳU٢RI:�� }b� ��Z�����!��m�.S&E���R�;����4�#s��5U�4fI��Gm��T�GT���U��� ǀ؁y���U��n:Z���u�%;p'@�(w(lw`w&���{7����8;I�ݝr2hXP _  =�{oC��v:i��9;iu�k�q)M�u�u�gA�;�w}<��c���m� �q˜1
� u La�
 �=�͢l��p;�n��5��ہt:k�p�M���].����Um��v�p�:�k:ܻ��@       
              
�JU<C=J�TF10 h�d�  ��
J� �&&�  L���*�SjaM1 �hh�ё�)��J�B �P4�   SU"d&@�#&��4����F��==&��*(!��Rz�j4фaɂ0����=8qr���7,{���rrw�m�&�_7�������"y	� ͳy3�?ܸ�����66͛�ݹ��_����p��י����i*��#s�l٦rC���9ˎqJ����6͛�l��L�UUU6}��-��u��c������O�������U~�ɧ���{xl���~?_��M�=�%<s�Ĉ���@����p�;�c<GxA�	Y��=;���:���E�Y�}$_�x�3;p��ӆ���E�[k�����y�ׄ$�>BʨJ9G�蓲 ��Ē'(�ʙ�(G�Bt��L@�?$�3"{�Ǆ�N\'��l�H�A��&/�0�'9s0���L,c��:�	�H����r"�^LYÂdza<#ۘL�)�t����x}3�tr��Y������ē�%(��3	�ar�x�F#��vbDG�1�,s&�rc�1�O0�3Ae	1�:#VO�Vb��9��Ǉ�B	eē"t����'��	᫘�,D��f0,�V�|�fbDF{0��9ً�	L���i4%��"`�&G>��&(�b����"$�<'�:p{��Y<<e	���QӒ��H&!/�(�	����.�?C��<�f ��N�J�t�$�,����KJ(��~������P�q�	y3I�&$I���zaF!��R���ID~��0����8rS��c�B#�LYe��2&�a,�x�N��f30s����vc/�Q��H7��N�;�:t��R˥�A��5��t��E�`�-h��hG�0�Cq1����Q�DBx�ra�D��}�*�! ��"=��I�@������"53	,@�\�	�r"����0�#��Qg�B"ac�Nw�,j�q�>��ǹ@��,D��Ĉ��� DN����>�D[����Rb�� F����"#ؒ���M�aI���H�"�͖s���B"�	��� �(s"d����,�.�<t�<�JP�=��}1��AD@�$<�D~K{�e\P�Y��ds��<�J`�ȁ<tj�~Bk��@���$�q��D���1�M	��r'�	D,O�(���ġbx�(��8 ��IxO+"Sŝ:�BxDj�pI�Ĉ �pD���y�H�GýbdDn:"G�&�����<�8t��H<A,Ģ#ȁ0I1�OJ	�"Cq(�ǉ-���I}1?!_?G��b!8'���"{��Y�y�?!�q��E��JQ�<�2`���P���������2@�}�ĔN�O��C]�O�ƞ,�\ƚnGH�g�P�#�L�7�qə8K��(IX��8q��u�JX�r%��%��'Ǆ�c�Od��}33S	�L#>'�_��Of$���<O�8"v�m�Oc3�8w	0s���O�dDtb.jf�a���.�=�$Ϭ�Z��c��G��)�,� b>~}2z!fi�,�fj:%=���$��"Q8[�&������N�[��u�&	Ӣ=ԕӼ`��'H<FF:#ے�u��ڿ��uV���]:����t6u2�d-���N���N�ř��+&'�5<y�τ�<b��g�����D��2&Q<:5蟟��DȎce�"bħI-�K�'��Lb#�Ȓ�M��NBp�}@�"Nv%~Dr�l�B �$L}�$,O����f%3��~��=BQL%��&D����w�3��:a�xHy�}��BaB`��S�w�OJ��
�DNng�x�b��"'b"�:`��R��py1< G���2"x��;'6ýQ�?��i�;�aݽ>��zI�	"7:#�f�8fA	�	5؜�OD��g�e,�ӣ�!8a�����`��	���B"X��$~ܒx�J'~�K�I�����'����&\��`��ȝ(K�"<�	(���:'i��G;n>A-��:Q"TBP��0�rc8&D&�L�c�	�$���(O�Jx�$�z����IN�{D�u���$��#Ϣ�s"xp|������y3k����rU��΄�dN�_Y/����G��	M�ф�Jp��~�(�T�"s��fk�Y�"S���L�I��Ʉ�0���$��;��{�3��te�c�k��N�oN^�>�d���i���C32	#52�3�6%�A+����� L��f�Q$�A	���	�c	;�	��������0�E�D9�X�(k&R��Bx:'�$y�|�7	G&?"7Q??9�?D�2`�"#��ϡD"=�Eȟ�똞�pD�"-��ȔF���O��8@��c���-��	����0��Q<�J#�G=0�/bOB%���cț�2'�xx��NK�PI�~n%$I�':t��t�{�&,N	�~����K�,}t�����J���K�"Ĝ(~��9	#�`�"/bOD���=0���.c�l�ޝ3��L���}F�質�w%a�5��'O��:n�O��n��=_=�N��}	�;��K�ĥ���}?x��'�"#�$GH��O=�#0���n!<I6t�p�O&�5����Mo᳥�����[:k�I8{�@�L:= �c�p����"Z#�����tLN��rc��}&�J8��c�LY�	��;���r,��'�ē��$�D�����añ�6j����F�Ӽaӽ��)��D#qe	�����N$D�Q��>���H��0����`�$D�0��8@��$ߦ��,I�N(�Ʉ�����<-�D�bDFc�`�����H|MQ܄E�~�BI%�"�G��8"�Ɖ�1��Y�[19َ�t�$>&Ix�QĈ�aGXOI��8x�9|�D��	�a�3D�'"��j>Anf0�q���I��%	C��Ex���c�D�#����Frc�M+�&NLĜ�õ�t;Ǧ��߿������A��{�'7l�o�|\:Ϭ��v畝�ޮN{T��
��L�{'���ˌ��7;����C�&�&ٳ��[�: y���94�����݉r>�����,�yevxc)��;��V���|t�nL�uX]����|�g9�e)���Ʉ��h���\-(]�Ͷh�3?�e�}<�=�.����$�d� C�Fg�����������3ӝ�*xx��\>t~4�X��u<�C`�N�}0������_@���=9kZ�u�y�w#�G�V��i�ftKc
NzB�3��3��C���"F9$��|�&rJ���1̘w=<a�M���T���p���L͘ag�C�ه��J�������~�~4.M!�@�:~�ã�?1��Ϟ����ޚ���tip�3د�:t�ᐦr��P����x��!ñ=>X3H3��|8|��
:n����'� !ӧNO�8���+����4Y��W�{g���p�������ӯ����~�z������h�ǌ~~0�Cz6k��>Z����ٳ��.�����O.�5�R��m�OHxeUl�S�8i8x��&���8`��<S�xK�6ж���m���vЫ�Ǭh��]�LY�s*��� 0f�Ha�͐�<C�qq����)㧎�{���hK�0�Ja��O��SB�����������N�?��ܐTL�S!�g��Ɍ
04�`_N �L�3��<'���iNjxp�����~�8B������;��1.�|4d?S����&t��f�3{<C�Ӧ��;�L8�CL!�:y�ERA�<p���O�O7Ҟ�\�x���x����;5 sģ��x��;� �K����i�W���4�Hp�8|���di3 �����AtA�� �|gt��3'O���ӄ0���e�C0�?I�:|��2vp���4�|>� }�H7&�>Aæ�?M<��w���0Ä�C�JC�<x��O�`3)}e>P��<0={9֗NxÅ�AAp�0�Φ�a�M�:S�L<ol�>/�0o�y�k�ʘB��x���ϗN�:~4���-8q^�����>Ɏ??<|Ǫ�cG�2�?�(ϕ0=����(f�|��)�M�<a�S��p �OLںi|8p�c)��<~(��;���D0��:@)�u��&��7S��<p����;��0ẞh�����N�����#<P4Ґ��m���Ӧ���1�9��I>�dӀaw�*���m*n�a��o�:R�I$��' �Y��{9ќ��L0��}��k��ኸx�N�L )�M7�\��2tvI�2�ܳ}&��g�tK��}0-��`�W�������<}���@��Hi�?Й)�6N��F��Ha�� y�1YF�a7����܎`A��7�zp��g;��gM �&�G�Ή���l��̌gJw��7��}�3;9��g��Fv�3'vC{��rrm���q�4�δů��(k�h싯���HB��S��)��N�`~���r�c�&����K$:\��	g������N`�0#���3r?s����\ɵ;=7���{�޳9�7�>ç6GS�ㆴ�0��'N��9~ZW��)�M�z�gfa�s&����hFg��Ã���ˡ�\��o8��s�&��IL�F�x{�m�w��^j���$�җ��΍�,��L��p���0�NN��o��<� ���w�����Y��w�a�yy:|��x�˗�˽��>�L����-�
�z���N��i���:r�+�'91!&�6{�C��=�ӽܺ��3��<g=0��R���'����N�M�\�o{���s*��X�u��n[�Ǧ����(lӹ/�®�3�͝�<���X��/�2��t�9˙��w�3�:�6L��w2p��}�xI-�bۓi*D���W͇�V���vZMQ�nM�Ƙ���p��ɯ���Ky�����zl��Y�8�vt�L�@��t �\�o!�#���k=��Y��J�ays��Ï��q�H��y����~ٔ=�ӓ{�×��3f�ۡ��9k��S��{�v��e��y�\�K=���wl���׶\�r ����P�6��|:{�r��l�I�	^:Y�+83� �B��`V��(��?d;����#��n;�Nr���ỗq�zC�hr���|`�qNcrvI�8e�y�n�|��X�G�x�9�U��9d��ڔ��sr���9vr(N����e=$^']1�h�s�����5q�]��I���%�G��Yݡ���N�ݘS����f�����ǳ33��s&�J�zf�K��zn.�}S��N���Yo&��,�+=χH2�>]�sxĳ���8��~���8fW�oN�4��uwswL^9�G���I�̟&��5��3�Owl=�g��?Kß����3F���&��w)s�܍��,-��I��V�`3����4�ʝ�|��fn�NfN{��fw��&�2p���ҩ=�Ҍ���PN�D�95y��d���&c��8|��7�ä(�?8C�4�G;���&�k��1y�<�~/K{ɇ���:2�rv����L������<����z	����/�Y��N�`-)�Ř���f}#�8�3�:e�Ɵ�L�ܟHi��`Ɲ4��N�8E���6�<A��Қx�9;:3��O��Kǎվ�s%{={8S_'4�9οi�4!�H\�?ML�Lj^��;vz�`��
u�Oq?+�
SU{�ݝ�1u�Ǌ�����i��1���ɓ�i��Q,�Ҙ�{��<�4ḟ_`v&���N��'�?z[�(��ݒrx�Ȕog h��8i�\�-7���@�Kܤ�0�������*a��}{W�W������?������(�l��_����ǿw�{-��u�7o�<ݻ�v<�~*��	5���n�'�����ǋ�g.�s��������v�X/�J�	j��|�����j�n7G{�۝�;;��1r�j�J�H��Q��K�u��P�������i�(:�4U�F5���o�� �sI�?���;J��D����l�]�d�Q�\k�M
�u����Qg7dj���/���J��u�%J9��Y��8�Ʃ:C���ZX�
�zm��
k$F��R�!�/�r)��e���ɛ�AVO��u}}ʬ��<�yR֞�)�<�IUǨ�ꨖDKb_}#�4�0uz�UB�V& N]�����8�#r"?�6�����P`����s���"��(�ϵ���64A��۹1���pJ�E�ڀB�>�)?�T��i�-Q�ˡrB�J�D��-&5A���Z��Z��>ɤ6 X��"QmMr`Ћ��
Z�	V��U�pt8�wy���'f)p���7���[��*���V� �EELI �1KO�JR�$R�DFJ�E1 ���b D�	FSv��KLTP�J�\��-)�]kR��v*~����_ l+	Y"�!\���D1T��b�M@�i�R� SVT�SP���q�y�U��$*T�es�gQ�W��B��R�T�%'۔V�Cl�;V5K��4�J�E�Z���DA�!�_b��Z����&|��ەD&bX�D0A���F�z�ci�ZcܔkP5�{0}%Q�$�'�e�$G�^��c��_@�=ti����KG$ġj��"T���1��ᚇR��GmH�h��B�mU[�d��]��*5_!n��Ui�Ғ��>�r������=�ůD��:flxx��Ux޾�0�g�n޽�qn���z:�����������������oo��ϧ�OO��������������U\a[Y[YU^��U��U���߫ʯ�^*�U�U�եꭢ������ʪ�����iUz��\�����>���>�#�����>�>�
yo|�V�W�
������������Y^��wwwk�iU_+J��ZUx��aUWUUQEUTUUq�U[YW�|}���� ��">��l�-�H�d9�s_y�s��9�qx�J��eU[VUU�UUTUU�����TUUq�UWUW�ҭ*��UqV�W�ʪ���Uz��������v>� >4�7wy��u�-eU_+J��^*Ҫ�YUVՕU̻���\VUU�UUTUUq�U�^*�U^��U��eU�=�/9�݅�H�D["�-��//6��l٢�kD~���/���m���rp�y��nos��朞�c����H<H��pN�"X�%`�'DÅ�F	ӂX�'�K<Qӄ���$��'��$$J AJ8"@��'��&�W�8q�F�Uh�j��	���DN���$�D�8"<��:&	babX�a�aB`�abX�Y��t�L8"tO��:"A �x�	HI<H�p��'���X��`�	�C��UV���}���J����-K�.��N�wn<�쩎ۍ^c���X�+cV+�(HX�$�5�V��b�!	Z�A�/n���s�u�lk;�pd�+�[#���ӛ�y�P���cˍ9eU� GTr��Ƕ�66�ѷ:��qa�����=�8�7Q��ݒ���ۖzC����sŚ.x�K�y��v7�m����1D����e����`��a�1�#v�9S��GK.�i��)�����:�s�;kc6[.r:g������.��������ش��[,��b5��쫤ڶY.(ٲ�%�7=�b�p�N�x�.�˜��hS�1�ֵ��`]���O�ɍ��m��u]r��Rc��:t��:��m�v'�:Ƕ�P��u���6�7F�/<�Cɝ�PyZ4�G�^3�Xw+��Ӫ"b��Ȫ�+yU�f}n�'̵�f7��&�ݮIPV�At3��ޮ�%�F3������	l�'���:��#�c\����n��b�y�-�|�-(��"nA9�P1Uju�H0��ڢ��6ɸovZ�yM�痶nN�M768���K��z�-õ;��������s���al���>ۓ���6��gm�����ujю��u��:8�mp��X��m�q�x$8K�$"q����X��G�$�{{{r��l^��=s��q����)��h�1��tF�9�T<� qj�iE�\�\����r��=cp�c��\�q��J=����P����"����17m'�Q�;�Q�W�A\�V�e��8a�D@Ў�1P5�nӬFC�[$�"I��֮y���wQ�ᴈ �o^����W�ɺw$�qGq��m�Y����]��u�eZ;]N��bvn|#�Gz���;Qmv����[M��Yc)c'�T�a	�b�_b�5�f�E K�J	֚g�i�)�w���ܯ.���%r`�Qn�e�]lf�W[�N�n.7��s^�e�;+���v�k��L���An�����.r<�9uv�q�8���h�v�<�u"�ٵ.���π��ǵ�/��	A��4�1���rHN[��֋�M���� �m\:]h����#�䛝��m�u����,�b�tv��L�b�����mڴ%�;b��k�f79 9�
���W��m����v�/O
%E�wyY]ݶ6,�Z܅b�3�t�+��9��u�J�1.\탗���m���ltu^��V��O�p��ej�ܒZ�����u8����Gi�N�6{��ۉ+�̊�����㣲/n���,a�i��Ǯx�#ͽ����5�{mmқ`�0��0(X���2���!�7��$Q�M����=r����:��_��t�.�#�7Ӷ�rt�n�5s8m����G\�x���F��k�N�6LR�]��D�¦��AI:�g�Ж�top�Ѳ7�01ݜ�=lv�-c�D��s��ܹ�=�,[��]�{�����:u��c�����؏
]��I�\sΫ]��d�x�x����;tp��hݎ���7%�̹C�N�[K⊢�{>^Km�w/\�'�h���7��U�6zݢ˹����8�R6Ұm����4��X����V20��ctVѴ>����\�{�-����á���}����wwwnÿ��������n���]������II0��^�돝z���e�
�0�xC�y�^����~���8�kۓ:��t��r�`*���ظڇ��6�������P��ݎ��LܙK<�=�j����	�c�d�=�z끍���s6z���cq����za�ffC"r���7p�/B!6	� �&FF�es⨋���2lV�Sס\�a؜QҨ�D�m�>���"��tx��k�Z�u�ͽ�Ƥ����m�2b��ͻ�&�q���mΈ��z]�n^�,��81�c�c���t���ѓ��G;��=��gr�V07k9��2p=uGvĎ�)dm���[Y�wt�-"�n�LoUR�o��G��&�8r�7�N.,�>�S��U�.%�(� ��hO{6�	����S�������>��x;��$��>5U�ꎯj0{V!�8h���/��)9Ub7\���|����4�㋦�e���Ǿ��}�U�.��C�J�$�~sV��[X[mԛ�uVWK���uf|ѳ��h��X�tJ(J0æ	��7Yw!C �!�2��CGh���2�k
�ƾ�.�GQ��P��vG���Q��N�*!����­!E���K_�\u��e�3&a��vڳ������ڿt�,��a>E��0���|V��0�bX�bY�(D�(��'�68�� �E
Ua�E~���Z���F���1�%}K�T5Gh@�F�UQ*�]G�~>X.7$u��Y�ɐ4�"����y.K�W
�tF�[3z���"�y�K�!�����U�QZoǥ��j��ӿ'"6-�%�ރ[@w�,�k>)��M��Y�X�pJ(J0æ	�����_@'#�����<��䧮=9�d�lG#�E߭+R�9E�o��X?��(�'*����Dtx�F�cU�]:5�	e�ڮ/ā�Z��I���'���Q
0艂%�e	B%	FtæΆ�:u鎜~Yw��Hi�$�QQB�EMV����d��L��fS/ͺ+��m+m3��S�r�lݤ����3���m��]�\$Z�g�.��6n�l�����Mz�e�ox�X��˃ߣ�j�v���s��yc^�1<X����U�k{�y�S�⺷Si�8䲪�W�.�G�|�#Q��B�������(d{j�5M��f{=bcgӬ�|��eޭ�퓛]ߝ�>��z�qz���~]K�\DK�]�>��dm�)'ޣ9���:`g��%s����kZ�W/g�-����8�=q�$���:`������L��o��[��_G��&�#��9��}lU>�mU�e����;V��c��n��ǉT��,A'�V�.�p"�#��,����L>��k�cO]�G�4fF%�v�4v��I�A���x�-0�v2RLL|W�7�ģ�%��%�%�%a�����0�}AQ�0Ҁܕ��� _~ղ�l�G�C�A�Dn���9f,�w3��s�f�IG��2JH!+�����̞�D���uZ�V2��G���}i��GH�e��lG{Z����+50��1��>�qy=y�̮���|��_6㮸�K(J(J0æ	���t�����3p��(�7���hCT\)�P�:*=��fZ���7�-&��7�ކ���w�z�
�4�����6l��UmJ����!�VY��K,���[���VQ���UY7:K9�����O$�I�[m�Z�7���OZu�׎����J�0�xC��qۙ���@��ݛ��]���.ሶ|��d���$��
�8�i)�G�Y�ԖE�꫌n�ٙ��^�u��ۤ.\oq�k8eLY���x�>�rm5p�^��f�D�jȮB.�D��b�>��X�eY�Z����{b�.w��g�Z�t9�:��5��r�_4}Bt�hAϹ�ѝ�R��f�vr��QM<�����oc���x�#3sV_z֭���q����#Q��-YUQ� �2�!�PV�	��̳�D�l�ɭ[�G�V�4!�4}�S�j�8x���D���:a�gCcV.u�P9FRl��!��>X�r��Uv��=���!��RQ�0l����d�+�at�,�Q�,9T�ՍQ��﫢4�bZR��~௢�U,���������_��aЏ8Y�a�4J�Pq��Ұ���4��"�f3��̃�>46j/T^&~X`���/e��>GĆ�/ǉ�ƌ��l�<|N��h��IH��h���RF�I��a�ؓdix�:L��i�釭����xO8x��Oa-�N���V�'HN�i�N�Nia4x'��Г��	��xRɠt)��$
>����Y<Y'�h�x���Ɖ�����<O&,�>���~���~?G��_��~�~4�?��`�Ji8F�&I�i�p�4��t��4���t�tI��f��c����ֿ��	ӑ�<>;F���#��/�d'�,�,�<JG�d8_���I4�r&Ĕ�S�dI�	�#���(��ƞN�Ƶi#�&��p�r͙ rl�b/����ݤ�G�����O�L���i��x�ɱY#��)� �^h�g"�j\Ƹ}��r&�g87�]~���Z���f7>cQ�^}�֣k�Vk�,WQȩU�dAEWjs��V�Ȣ�<����^ǁL�18�1C��	�ɍ�������]��Ř�\��񮝸��y�����ˆ93FLz���>��\ͻ����������ܻ����7��������ln���]��A��,馉��Y���ˮ��u��m�ڪ��q�$U�U?�G�a�rXudҪ�����X�Q�*O�8%@D��5#�%�7!�H-**!ٗ1��,�A� �&'j������,�0���TS���C�M��щ�u/5�!o�7����ɖ����^,=�N&$bJ71RmOqn��g���+9ԑ��IJJ�g���2|�MY؎i�:��hH�N֙�ىI�� ����SeF\[+edU�0�º�K&=���פ�I=+������<��I�#qD�*ę��\u����x㮰묺�N8��[u�J�I�b��ݫl�%Y�?a�A��$�n����SUG�X�&Q*>�7G�,G+�@��Pp���#P��?|f�˥����H��IJ��&E�l&1�[�I�F	���`�����2�ߞ������{^(�Y4����S��֘z���!UTX�2Sk,K�ٓ����yV���bU�	���lE�md?,L�'�K�h�Y*��$�$���K&�4���L���~��'YLE��O3�^ukbG��j=fM���������"ɉ(r*idx�1�$�/~q����O��i&�Q�N�K4�2]�����i���lEI1&�D�2H
��>��jQ"��@0�C�� bѽM1;��M25p$��s�ْ�J�z B���;��gל�^TQ�������~[�r��^���Q�������)����z�&�fO�j"⦨�����d˼��������s�����5�Z�{�B�l���u7�����I�L�pǘ�F��V��[')�bFcoŹF�A ���Q�
�V�z�s�䕅W�a9.m��_55fM�?[��{�����ҫ��G糖�ͩ숱1,��ec[��h����W�A�;�e�`!cU�	CAi�nY;��݌�duUē=V�Ri�c�Jº�L*��f������br������j��䶋%�Ɩ�Ŋ+*�Mdj�J�Y�J+�A��b'��~de�x��%7,�	ѯ����4�1&kLHm�U~a0�1�G�������ʬUi%��?2ᅉ��~<t�M4�M(ӧO	����s��:\�K�UDDJ�j������"�.`�H��'���*�+߇��.���vb���r��b�⴦l�U�&#��V��V$W���fq"֖?,L*�f�&
}>j��0��J�VIa�X�����|ԝW�S�&1'�S�id�Q���^�#���U^FثO"q�g{�����ɫb[q��zH�
k�餴V۰�4p=���؟E�s,,c��ZL*��Z�e�W���bK'�0�Y'VXj*UWq$�O`��3O0Zx��&dx�4�i�U��k���Z�nE��f&E��k'�F2㭺���pM$�J4���if�>�&ff	��,>#�����lj��~
�����B�F�e�h���I�ڻWc�&U_�L��TMō�[�ۖ[i$��r��K7'8_-�RW��"�T�͵l��@�T�Qk�X������`V�FS*��{b�Y�J_U�
DO~6h�.[�����2\�]�5Tq� �W~������U^a�	�w1���)�Y��TvY%��*���UK�$�R�e#K&�$mM�,EUpa&lN>��c4���~Wk-��,8��]��$�y�u##*G%�5bOY�`��8m\65I�DJDF�����{͓��$��a�Tş��������<mÏΰ묺�N8��^��q{��[E*�T�\�⿆]W�U$�nkoV4�:u^GL��y'���Z2aUT��E�a-AjTXZ�YFQ��w	T��׈��8W*&M]"]��yR-�Y`�l"g�%EY2�ʲ�Y,�~�.?4nǊ0Y�IY0��F$6V�b7,���1�2�XV�Fi�a�{��ch�-{���|6�<Ë%�̳���^�\c&\�u��j��yy�c�!\e�JaSa�ZR�П	,�T2�2A(H)��� �痗_B��td�'�F$����0ڞ�x�L�ǧOŚ~?�Oƒi�t���<p���c�I&
����6^��4�����r\��+l{j�1�|3�9�xۑ�$UGJ���ٝ !o�����nv��>���tk��-���]q�Nq��k;��fp��&o9��������ۓ���r�r͓�LB��n�$A޾U����~���<ֲ��7U�CŐ����T�I�:��1%Q_�<�0e����S$�U�X�,���0��j�&����X��56ħ�_��'�`��?	3YTА�H��id)*	P2�L�VW���bG�U�S|/ܬ�c���d�
Yab�1��ɨLA8��VU9��_�8�i�0�S4j��s�fK��j.��PA��Q���\6�����}>e�O��o�:������8�:�-:pD�Y��9%�|��Z���MWj}����߂���r�G���j��
�!�qe���c	���k�e�}��ˮ0������)�M�*V%id|�*�8C[j�`������>4l�����S�SFVD��[�5KM3���v���������s݋mչ>?��&�+.���;Le��7��Yh0�.p���1�ţeqTԧ��i�-ƻF�2�J������W�Oc9L���~x�뮿<tA?I��iӂ'���<p�
����-UPD��>�e�GfDё`~IG�����O��	�OU9LF_>b���M�>��bV�=FC���>6R&U=J�M(��Xb+��p������(�%	X^�jD)$G�\M��[j��*�TI4��L�J��x�5��_��KX�<L�0e쉁�7�)�M�5�XV*!?dd>jF���ϪD
��M��~ڽV1����E�=�4vaȦ��3�x�"�����bq�2�)����]z�������8�x��xчN�:x��d�%�I�UPMT*~����4&:�����na��	�L�yL~\51^��D5ϾW��\5U 9���X.dO����ôC|��֋�>0�qF����;ſ��nm�w#JO�	�0�a=S��I��nz��׺����<%n��UV��H��l4��2���R�������?���د��g��}�f?RfO����)ְ�]����6Ɵ���H~ �'��x�!4Y��>4O������OG���xz>	�$�J)#D�0�8aZY)��x�4B�������x����<h�Z|a,�pI�BO�<_�<_ǉ��<l��G�<'�œŒ��� ��M
h��">|��'�>.��&O�'�ƣ�y|O���ŗ����=���?G�v�?��?����|t�x��N�&�a��i6��4'Fb0�R0�>/IÑم���������'���觏G���xp�deOc��'�'�����~��i4~&����J𓥐iFN��	�i��Q�'��Vg"?<{>���;5L�gr��xUӖ2�wӄY�wr��� �Ӽ7f�<����s�q�v����C���7������s�o_Ӯ틜�LD��{s��t�pٰ�Q�'xE�������2g$��Ly��r�G�	��֮.W2V�δժ>���7��V�X�$N�uD�g8�f��r�P�,���j��z�
bm��s�V������36R��׳V�>ψVq��9s�5nNla� ��F�nTx�ɵ]b��P��myZ|;��uHU�I�ȫȵ����,[�-�����o�V(�c�J�s�G1�c��)SDB	_�L���u�g�ȡ�秞��U�����������U(�1�ֱ]������s��73.��~U������Uw3333twwwws3333wc�'���DM$�J4���if�r=�ctm�@X�1U�YO�^�|��85��1k�b��8���N���L��L�nx;9tr�p&�1��X�Ṵ��h ��=n,��s۶p����;��;[���X��v)���%�١��c2�Uׄ������m�퍳��������G�%r-��X�8�����\ѓrql���·Dn.UN��ۙ�>[��ހ�s�t�D�<�\n�q�Ս�q���b�/Kշ��9�����G�у�+�����8�t�g':��-��' ��{���Y��7g�xIlz���;�`FB�����\>�p֒����8�w����'���c����ʢw���{�)=8�W��5o1g&;w"y���۲r,�eּ,��/y�����fn�'3˓��O�����s2~�=�rop��L���|t��sF��W(�pFCF�N�@o��U�Y�m��g�=N7<fƟ3��x��!��S��d�<>��C����6BF���:�i�O�������~~�u�����>�$��T>�eeV����}~�~]J�x�m8�<[v�2�~�	z��.�]ݬn�ƨP?�Y�>�B��r;j;|�\�z��n<~~~~q�	��i�t���4�N�=<�m�iUi�O�v���y0/�k��h��Ո}��A"��WM���4�����'�~���;F3+���?yn�Ux{4��`�?<O'��qT�R7	��+AW�Y��(�U϶�ǌxۑ��v�ػm�3�佛i�;��c���}�x��c��'��K������	�m�����x速�$�J4���if�R5	�e���#K^�Ui�?ia�~y��/;V�o��62�1�0�:6|T8�\'g?~C(�տ/��,i��+*��S���K�{���˫��ܝ��d�S��|l���~b�H4�+�LE�Eu�V�l2Wz�F��}�1p��0��#3��>e��̞�6�ܫq��g���4j1��Y�1���Ǌ�c{竊��Ҽ�ѕz�oq�_�<t�D�M4�<&�ig=�D4O��K�Ȏ���{���/�?Wȇ�}��ʬ� ��2Iwc�xպ�*[�n�E�94�����ݾ�>��8r�f${���6��,������4l�*�o��Q�?V�ta��⦅��o�WO�z`�u(���-���{G�ǋ<��V31��!�x�v1'����j_&�Sn1��ʱ��a��_8��<m�"A��pҎ�K4��d��� P��g�F����X�&5J��5q����W~����,#xӭ���چZ���7+dM�Z�����s�<e�?JM����%ٙ�\�DkH�ן�'�w����M�]�6c(�Σ5���N��퍒�ۍv�}�{m�j��[�
���!�	�}���.�ίhDD��gύ�[U�
��`�������d�
��y�~U���wg��_eI'���ɖt�g٧��/dԞs��Rnxnd�&#6����Էn����j��.�����к��1m�>8fY'c1���0m���F��5n�c���Z�)OXW�5P����ҿ[cO��G����ed���w���t�Nw���l�/��mf&�Yٷ��'�Ye�}�'��x����#��m���??8��W�Ox��6t���h�fHK�#��ui�SV��%
0@�5��Yx����X�]���n��ߦ�Ǿۧc���1�zR��n;3f�䵔���7�ޣG�3n`'.�>�U�{��������IM�@�3*?}q:*�T[��������T~O��M��
Y�Gc-o_[��6�c�]i��2��c^��cl<)Yc1���z��~q�o�8���0��gO<pռ�4Y�TB����2�/T��٘fz�p9��믐��5G�,?mw�]_��˳gL����D.ϩ	��&V��z&��4A��D+��\��8e��.dVNa$:�O�9V~?pagVBôUf����-�.U�CT%̸ֽ�g��Fg�4l�[i����3�;�ۭ��	�!uճ�wr۵����Ǽ_�D��,٪�վLGp=�l�<~~|��|q�t��aӦΞ8z�c�\���q*!cFglKUU�>1�?Gc���Sg�Ko~��Yͭ�ǣ���}P�B[+h�C�O��m]�G��b|�r]�љ(t�z�;[9Ifsgm.�w��<}<.7�q��վI��a�����U90�X~ͻm�����G
�^6���a�/�>~u��6���M8iGO	��]��y9?w�4w�6K"������h�P#��n�rc�)g  BY�Hg+ꟹ���UkG��\�o��'�ط�Q���&y��^�5����c_>��,��.n
�����s{���)Q�Y��,�V��v��m�˙|����t�F5�~�~q��.��y9��'���&cQ�#��)^����ӏc��&{1���F�X�����2~�Ct�ѯ�����48t������Ɵx�㌜�2f6�y7�{��M6��؟2�K1�i5%C1�V��WZ�/�hh�|p�aa��+��X�T�0�q�_:��?8��4ӆ�'D�Y�Tip�ǭ��UQ	�e�<B�?V�щ;v25��>�����le�v�D���l�����0=G��]Q�@�z�v�7φ~���'ۣe!(�;P wܘ~�ȍ��1�iq��b�Np�_��Q��Ð��5=x�:����d�:�{��`su�$�e�h)���F��t��4L?Œ�#�x�|>!4{�>4x�	����}��	��zFF�8i)4��p�>'��/����l�D�~!���=��p�<x�4O�ap|a �<K|Ox��=o�����l�>=|'�x�x��׉�GKR.�4AxS��	����:Bx�C�O�ǣ���|>��d��|'��c��_����9������:5mBN���#$�IH�$��>/�I���l~<M�'NE��th����vx�<N�������!�����.">Ő�d<60<A<O�����ᇏţ��~�����ц��iI��$�i�����������nO��$��n�w�7s�̫7>�k��x�=˽)ޚ�1������m�ղ���gV�j���d#kZ
�y����#���-���Qy��`�c�nק����:8���ڱ�ԭI�u��"�N
�>c��o{�^�g)d�������]������8D��;�;�5�����۰��nfffn�*��������������������,�4�<t�D�M4�	�6t����D���5��*�N��v��;�_-Ʀ�^W�ͫm�79�1����n2�Z���飍�,��R��~�р�%q�FF܊,3��Fc��|���S�e�Ұ~$�q��O���&�Y���*�jO�Ca�;4�V~~���n>�2n2̲�Y��a����Ow��<m��x�n�z���獾8��<Y�GM�<p����H��aUUD�ӆ��|���>J��ϝG�(�TM-�:��H�)��h�vo5��*�f�or��Fz����4�P�YG�!�t�b(���^FޫF�UXm�]~�a�O�|@CgR� �%�;\6ڝ�i]i��cL�+]�O��;F��VC�7�WU}S��3�a�/x�󏟞6��뮴��:l�㇈ގH|�q�-t�-Z����-�k,!��m�w�s0hyQ%�E\m���d�� ��h$��bvE1BG�bnG���!Q�ɋ�;_E���4�oE�Ž#Vs+Q�-�z<�S[q�LM�c�y�7�_u�1�y��/���/�.9���z��&��ӡ�i#4z�H����稅��&��V�"@��B�D?�7~��2������k3,�|�U�F�V�l�&�ޅ����pe]��e�a?Q����{������q'��5%�~>�Ĥ8PR����5��n��ұ�ט�-q�2\��R�-��������<Sgf����S�䕆�m�~0��LH4�NQ�D�Y�H�Q��UD9P!��Y�C��QZ<a��ڔ]%A &uB�|��ʻ~�I�3;b~n>�,�2�e��u4>�eJ�V}6O(���M�~�ψ��r|%���?�9��2֮-������I�����jw�=)b��v8�K#�L'x���o��Ɲq�_:�����i�NtO	���ԒLCWvmUQ	�Q�����Z�Z~������6�<V+���*���r�NL;��K�vpk�x՘��v�5U�0��h7���FI�٫�B���MQ���5_�l?��Tl����=��l<ԣf�>��˔ҫ�,�e'�Տ�p�t��-��z�`�~����z��s�͹�[O]z˯μu�����q]<x��:l����QO�#B�D��*�!u���{[�M^�ʲ�/U��Z�+t���6eH%א���~>�z��SFf@Fe�#X�LO�J��#]�ns�o�(h,>�Qw@А���Y�/"����9:�Z�M�6��V�U?G�O�O�SF#笴�/�m���97��G����̰����ǎ��'�Np�<xM-~O���c�s��nQ�+��Y+����7r����'H��_�� !/n*���Ų`�$B�L_�y'6M��xc�b,��l�Q~1���e�p$E�W9��r^]7\�7Y.?�s i�B4�c�sd�}�G�MC3Qx�%7Y��(��S���t9KD�T]_x���) �]!���e�XbX���5��|y+��dn�`�����ѰC�Ra�E��6ɥ?8��57�|V~U����곇�ȩ)J��m�ڬOc�d2]C��>�>b}�mS�[y�	T$���k�����/-X|�\�[4"^�x�Մb~6U��0�ǎ��&�pӆ��gO<^Љe(�!�%J�b��֒Ѝ0�p��ZZi�⪢��U�(�OQ��WW^�#��X�0���4fm�r�]F���0r�4YYBCG�}F�_T���Q��#��O�z�e��)��q�a�TA���)5�~˽"L��%��P�(�_p�Q���<p�K��9�W��z<x�}��ٶT��93U:{�f��V�í6���x���ǎ��&�pӆ���if�� �UQ���Qx4X��i~=_v�|���QH��\�f�Y���G6�ȹ	 ��a�\��y����FMG��䞫^*���F�V[b?��]5�R�p������=I�@�\�Q��w��k��zv+gz��_�]�ر��C����4!���$�a�,�����+3�����q��_??���zq�q�:ӭ:�ǎ:�׹ыh�+���⪢Re��E�	��5�%x����}g���ԙw��3&AR]�.����񀆪U2�9���Ͷa��e�M;��ʼl5Wc���Ki��4Jp�f}�K���b�o1��Z��&~;}��8_(�,2��~9I�Y�!��z9�.�!�D?:&&�ć�$�'�a~���O/���������`�:aZ$��xҰ�L&�&�0�#�t�N����:������z�^��N�sW�Xu�=u�v�m�z�u��M�>��"l��x�x��'�h
0�40H:��œ���d<Y<Y�����<O�ǣʋ=����l�p�_�g���l����?�ӱ��������]����:>�'����_�G����վ;o	���|���x|a�{�=o����<>����!�'�O��E��c<A<A=<L=ΐ����x�M��ß�������wH�qB�����wI�C�[|}ϣg�:���P�y[�nzy��(+�w�64 U�F�����~�@���zǼ���&�I6�dN$y�U�,���rV~[�:_<�����}י��G��۞�h�b��=X��Z��_�n}�ٙ�ݶ(���
�Ϋ-���՟W�)7�-.�'|m��v�SCd��=�{��0��B�i3^����f��)V�`�?=��k�ȥǂ�/������l}�sM���S�\����s�u��m	�8+�T�u��-`���=����	-i�E$��O�l�6 �nAB[�s$��u�;�2L�Y$drH�@#�:�_��w������ۻ*����������������*��{�����(񥈘'���&�pӆ���if������wm�lU�]9���5N��d-�7s%�S�1.�={#�x����81]���b[\��mЖ���g�������[<у����ݚ{�['�\魑T�^*�Ͱ��k�$
�\fU�>5��g�<U�1��^�K��{t�B=��������F�LO���E����]��������m1Q8�S]Y0�&�~6��Qi�6:1�;mմ��Szlr ��yw-LMgC�`�v��]���v�yت��b��m����S������ �V�knۛn�gsv�M룎ڝ�|S��1N��1;�qۺ�x�s��s��[<>W+�BŞ��\�Ym����!���.C�6�l�r��&\j�8����=w��Tb[�QdlS]���#�[����#ܤ��F�yŕC����FX��^dn���?�5G�B�K��?��pn��&�ѡT���D¼f��Z2�����F�����h��)�x�<-p�	����`%m�QϹ�����l� ��h𛦰D6��:cS������(Lt2�>����[k�M���ݕ-�SUijZ�ě��?F�S=cm�n<��M:���:x�`�&�4�t�Y���1�[��4e�*�!ҡ�=���i`�䚒2����0��{�Ҷ�������h ��.��	a��u��;�$�a�@��7VB�5VA�H|}�lm!��yw+�M^�,%�5F��R��v<e�|�ɼ�̶���V9XK�s�Y�tA�������n��ă�Y�:Y�a����"i�N:l���>��	d��6����$=8l�<4J���q_���ŷN�����əƣL֝-X�o�����]�Q�r�EM}k�H����3��Z	�\!�wy���z�P�P4���t��:����������w6�&		ų��>!�K�Q�7D�Q�*��W�^��d�l]}�%�#����'�wU�@Ī��kTA���&���t�D�L<a�Μ<p�Wx��eJ2���mUQ@���΅ѿc���~���ڲ�e�&��n�tl6g�B�r��ϓ-��|q[V��Ó2�u��--*�_��FO/�kݯYxj��j2�����L8�5��qƟ����s?4�^2�����y�qɨ��oZeMGL��͹Wt�����V1,Y�&uxu��m����=m��(�i�D�4�Ow�N8G�`b�5�R#1����j�*�T��ED�nEZ1��iUjX���R��� ���k,aZ�'�|�ɱ;dj�4"�P���,�qJ��R����xcM�8��b�6J��fAӃ��4�33�QS���&��gO�!g�!tpK(���(��[w$�tp�ㆈ~���?=q��L)_�,�p�f#�V��?,��Ђ"'M����*��������q�IZ4$T t�G�˪NQW�#)���Y��浌�f�&I�d!突�%�j��t� �֌��K�Rձ���]���A��J8hgIQZ;��<Y����Ζ�"Q��4O	����%�J��J<Y�LO��.T�J���1P~a�X1G�PlМ�P�|�Xܼ����Y9�+
S���yų����<v�!���0���v�J���<) Q�~Y�替e��kz܆�1�b���:n��Y������?	��V}� ���atquד1�x�u�L�l�SQ�t������~4��gKH(�i�D�<p�1����dVo�UD8P����U]�������~�٪9�L��3.�j�W�6��q����<�J����R��LXfXTYՓ;o3,�{u�m���Qc�={�a�U�Q����K����u��9���=�,�h�R�����{4ԡC�l�P����H���ڍF|��޾|��^���㌺�N��ǎ�u�X�U��*�-�UTA>,��m������E�D���<o�{��y��ɉR�����M���E�{W��g[y'/��<��J��9W��7H�?�tH�u��� ������_���L,Wb�ߝ�z�i�30a��fS���aJ�ܷ(���NM0�Y��J4�6t�㇎]��H��N�5����(�s�XԒb.A8�rd3�r8�E���uE,�ʛV(��� !/vwWi�1�/J�`�?�哹�wlh�%��j7�9�W&���4�;j����bx(XB���;t�h�0r�IZb������oh9����Y,]:޴gI��ڡ.�����}{�l��>��>�tn�5>V�oL������?}n�Å�[9c�F�9Op�RU��oB�$�Ls穪�]��V櫂4~��#��6���7YU��U�Q��h3��L`����Nq9�8����5������h��t�������tiE�aګ�F�"��~�fS�pæ���,�`�%	��<q�^��I�-�[/X��1bv�[V�⪢'���t���f�bJ۱���<�[k,;r�6��N�n���8g9r=)�4�6д���Ѳ��r��Tp�B��h�*�}���˕�6���Xe��vx�_Ls�M��3���N�\Y���Y���+�g��coL�=O>]�_"�W�_�4�ۭ0�m8´ A0�
�N'��,L<&tL����,�%�ǎ�p��'DD�"%�I" �X��"""Yepˊ�
�Í4�L+G8�H�a"H�$���'D�4�f�Y��i�"%	�YӢX�&%�f'�,J:pA�8��Y%�"Y�x�H8IBQA"p����ӂY"xK:`������bk�Vd��.#��vX�a�!���j#�a��v*%����/��S�j;��8����K�jֹ����8���b1f6^y�q�;꯽ݜ6�[�:�`ϣhi��70|{◓cvD�|m9�wܳp�b����G�8_�[�9�Z,m���o�w�nffn��*����������f�ff��ҫ�������<p�����$�&�4O	�K4�q&�Wb"a�^W��&e�\�>����~\,}9�4��gK�<,�U��o�\nq�����$ğI�h����]]~2�|]�PӖ��Z<6yR�a�V�N�/�fl�f)�W��飍��w��0V"�4�'�YH�=6��g��m�1�[+&���ÏmZ��6���\|���H(M8h���i�""
�鸵;]�U�E�[Yf����WR�D�4���kFù�Z2F�Ѻ!�X~�(��Ѫ��{��x%��Ӑe�HtTh0C���Y��[a$Ê�)�+c��i��$��0��y\�e�Ϊ���-I�U2�\���i�6ݑ�²�X�~�Q�[�V�8�����rO>Ϳ7�_#��=x��ϟ�?=m�D���p�<'M,�k=�ҫ�TLE�Ƴ�2X�(�{��\��"����&���^� ��Q��j�^���[����лk�n*�H����]�����\y�k\�}~�W0�m�>wk7�y����cn��_����;ۭd�`�����V9��'8h�W*�t�L	�������"���F$�W.܏2ז�J��z��&MJKd覍�s�q�6=��]����F]��`�hC���]D63ڿ�&e�<`��P�^�.��E�o����Y\eS��G�c��$T�(�ӆ�!��,��9DI'�K��X�igK+�2�:��u�j��Čن���UD�'kJ#��ʭ�mF�I�3�N�3��Vf�Fr�f��������=m���[��~�pf#����3�}�l�X���C�������ν�yz5�4��ԃ�v5+�9o���ݩ�6e���� 4Q~�2}U�Ç�Q��>�W�,�}$N�l�b}&������|��筽�W�4�xM<Y�i������9�MI�ڪ���R	*���]�N�~[��qWL�7kփa�@�(�]�����y�Oޫ�e�r�"�0�v��H���q.|�&t�qJ�Bl<H"p��y�!.�6�,���OҪ�_��2a���,��T�u&���m>Y�y[�#�����\�r1����|����筽"@�Bi�DK4�f��>��DB��х���+��v���TTGp�����k��iiAq��ژ��5�|A��s��U>`WXV(�Ų<X�Zxǋz�+���ӑ����G_>Q6p�u䆨�U�4�t�4xNb�DNU���0���������mOۦ_2�Ϟ�8����~i׮a���`�"P�p��,�L��x"9�h6��$���{�Fi����J�j�0Ѫ���BZeƷ� !-J}��)ǖs�Jd|���>:���c�"��8⏼e1���
��	�T>�%�ώ9�k�^@�\]u�r\�s�]�a3��WS�7��U<hBL	S��U��]9=��ڊ�~<S�l©�#��QZ8e6�$�h|%lފ��q�}�ʻ��d��/&'��aM����e�32z��W�%�N yCT]h<Glf�V����L�o/#5����9Bh��J{��p��ٙ�?e��	��,�$��t�a�N8p�ϝ����tеE˶��UDR���P��/H����m^?8~0�J�gK��D�tg6��6��a�f�ẳ=Z��F�d���G����O~d�z��q[�EBE��dt�'��P1��@�|�}F�X!h��������.����Zv~�0�[G��$NT2�,�~><i�a���`�"P�i�%�Y��_^�xb�l�KG4���b5�c؇��;a^���<�?Fi�cl1VL`m������%�L�o<����B���Xl U��a����Y(8�!�P7����n���o�eg�q�ɪ���Ϥ�?t�ݏ߄�4�~0K:%�"%	F�"Y��4�>�El��Ypa�J��z�>�I=W�'�|lk���t�B�Ը+a�����~����S��u��-z���^&(�j�Ή���%��-z�Tea��]Y��c�Z���r��7f���K��z�����ՕT_nmvM
~K	(ٴ�T���V��D���n2���^>m��<|�^?A��&���H�"p�<"Ib`�`'�Kb,LĲĳ�G�(��H
0D� D�IA8$�bpJ<tDD�<W�0�¸p�F�0�
�A���$D�<"%��A:"P�'�i��i��&"&Δ%��abX�`�x�Ģĳ�JDD��xN�B`���,< �$�$H AOLGD���:x�<%��0L:`�%��������9��8'9��E�0�����=��.�֎�A.���{6󜫝��܌8��v��#+Gsk��fv��7��C'CwWG�&)9
�G�Y{�H�d�T��8�|7���-�9��i���������;��}$�S�-����5b�1Tϩ��̽˂
��{��vdh�:�I�bmo@�!@{ǭG"�Lf��N��3��g\Z��s;�"�]�3�D˕߷q���9t!�h�2FI�����	�ښ�SFE²�2�28��R�m3[��ۏ`�q�Ca�L��u���������7���@���6\[�ގW�9�d��YI�P6Jܮ��v��7��]깹��fn黼U��������*�fnff���s3733w��xӥ�&	gD�$D�(�DK4�Ɯ�Cz��Dԉ֪	�,+v�����j�q���u�t�s��u�W�[̆����pud^����:��&�,5\�q��Ǟ�6\�c�ng��=�wF�s㸖˽N:����+���g��44�䷁㧟r�Xxy�v�daNVX��#
ܘ�|�e��6s�y-<OjMp�a�3�s�.eԝA�>��@���d�8-��Mu�v��p�T�v�[��tG�q���V�kU���g�������n��9y�ATt�B��>ݡ��c��=�����n��=�|�m��ط�����i�=gq�3�<�L�乊�m�+='��UD;Z�s�uP�\�M6�cR6�]Rw5�����NQoV^�m��Lۣէƺ����l�9&�W��ml%nة����������������f�!�	WG(�?��<;��	��ô�G�&�ތ4�xd��s��S�,�}G5���Sf���.�p�0���~�^�����Fp�"�cZ����8�>��y����E��������[���|����ɳ����/��o�	4�t���	bX�&aFa��p�Gu�B�U$��"��2Z,�P�(�c
����UTA����h �����wd%�����Ts�����[�e۠�C��������˯ߖ�v���i��gV��P���(��r�,��6l?k�}?2��&-�<]z�rσ�(�`۾ƛy&�����f�ǫ6�6A��t���X�$��Q��ig�6}o!�9'ڋs�UTC��%]5�=m3ђU|h3Z���4��Ǐ^�=r=5�4�{S���'��Y��K ��K܍�X�dх�rs2��͜���v�?'���բ+�(�~0��pd,���6|n�CU���,��^�RFA�V0B�'d�0ӇDO���J0�~><p����y��$���%�UQ�Ã�m%�hCB'�zQ*Q��?ȑ�:Z�8C-!�+Y�O�\0HB��ߦ80����'�@�u���aTw�����_���0둨�Oѭ�G_O�ӆ�4h8!�il�IL^{��r�r��e0���V�zeOϣ��O̲����a��,D�
0ᆘif�j��T�7xdtf$��I��e��^�~y��;+�Al��H��UY�  ��{�����բuX�Wj��i�B����>{^�"�[��ϻ��^���뭡��cܟ9Dݵ13L��z]ȭQQ�b�n�Zڷ���d�;+{�;�p}�VUnTRId�eC�%ԯ�0�WA�g�8oa��2����ѺЉ(�]��E�|O�4����T�����?/ed�+���珔���^|��_Oc|�i<B�,���-= �Kl�w� ��/G��Y�wF�s�w�X��s�3�(�å�"a��b%e�O�|��^�뫷oncq�[%�����h�J>�ڰ����]���Ӗ����mbߟG���x꟤N�����c�2_���?mx��a���UhD�Y��ej�FC>�$�����K�m�Y��Q��at״J;B\�p���K`ᰅW*l�4ez�Xz���%�X~���T#�0L<"a����ı�(Æi�<qג��d�ͭ�ꪢ�R����]j��j��a[�����VQf~?*yzlؕίu�~f���D�J�"}�Z�cŖnn�5��x_�9��Θ@j�l��fR��L��|�q��,t�Ȭ�W^��x������ET�Q��c�~8x(�?�<Y�a��,D��_4�뮽u�6�YĨf�Wx����<f�]P� O�,�/��	�<�O��%ǋ�3�K��G/z��x�r���g��a`!?&��r]���H�[5_@�!��W����(�}�	\;�bv���F���ik3�;4�~��ݯY+��y���f�JN�@hL�G����ŉb%Q�,�K4��(y!���i��T�sט�jɛ��^2�aTAc��m���̔DU)F�������� ���՜���?��~���+=��^�s����[�C��d\�M�S��ZMBswI�3w���w���yd��i�$������g�^�*�(�rm��&�M���n~��	];�.Ue4޼m�ޙ5$��-�f1��mNGe��M��i�i�^aVX���7����^Lɵ8�%��'x��SqM�g=���d��L��᝶e�i�5��0��������-��V[>m�����~u�_�|��Ǯ8��ό>8x����+@9>I�*�5^Ő=F�|b��7��a�cV�6�o�UҴʕ��~}L)i_IԘ�p!Tt�j�4a��
hjWQ�A	����B�z�O�h���ל�b�.�'9ň�_��������)f�xe߭���ɠ��(��ú�:�t|�w��wvZ�n?G�����_��~m�Zi�$��ҍ$M(�J4Ӆ����,�$�,L��bY�<t�D��$DB""&�B@�Q""@��p舉bx�>p�+�+�4h�L��G	IaH�"%�b'��"@��pN�4�M0�MM0Ot�,Lı,OX�X�x�C�B"pD�0��L,��0D�IN$ �x��pD�<'���&	� �,�9}���]c'ގp�"{����x�^�0��^a�вU�<T�ve�s>�oܨ��'�U����6D���_�Z���z���1Ȼ�dH�U�{O&��]�s��C$���; Q<^3w����wP�_��cF|>s2ws������Д�)p��y�c�YD	��%A����q�&<~�B����I�_=����0r�ns�՚h������g8.wow��{��37wwx���{������s33s3wwwz�ffnfn�首i�4�K��gş|p�㇎�*�!ߍAc������|r���-�l���0�a����2���|�~�q�O�~h�?K��21�����U��G.�k��?N0�Od����FOXm�n�BX}Hr��گtSj��7y,m�m)ǥ����?w�4�Uƣ
�
�4ӭ�~u����"Q�p��4�K4���D}tEED�֒�j/U�Q��=�B��a��Y�lC_��\�~,��,^��a����]ϵb��]W�5W�_U(�l��!� ����S	e
r�4���(9#(����[��K�V�L4@����Yå�߷E���M,����ug㥗A�=y��1�D4|J�	��?h�X�"Q�p��4�K4���K�s�}�Hݕ�f��@�*�C4EM�2��9�NT�'k�w���T��NL̍�3'��ɛ,ŏ�i��m?w���ؽ̜�t��"1y���ѓ����}�9�oS�����_��ȗ���!
!bj�٦�����x�����̛V���wFH'�x�G�u�w������.��
ۛ����G�U�6�u�Z�l�?Q�|�F���(���?m�R�d��[U�����~��$,���`�,I$���DOŋ�e�/�|��^����l��Z��,������svu��'nS��VÅ�G�#�4�y_+�}��E���q���=�fUZ�p�*��U���yd�V�ZY��0���������<�Ѳ���rbȀBo��s��Zִ2��g��+U�	4��&�ٙ��#M��
��o0�Fՙ[�]Ɉ���i�W�Y'�:x�4�N��_2���]u�]s�j��ȵz�Z��V�=�tF�f��a8�>%eW��0Nו�G�����E�4~0 ��o���2e����_�9&�^]�ʺ�>MK����:];[9��תT�ѕcN�ʝVś�~e��Kq�'�m�+n��1��/���L�Ͱ��D�'�4�N��%p��4�K466�j�H���!�l��X�ݖ&5��U�s~0�w�B]��U��Z�X��g�:�O����=_������~��f++$a��9����̄J�%�ǜ�|5GM�{]�mZa-�q���1o��<W�����z��Y:V�\�>�x�ݽ~z��N�h���4�BQ�,�K4�K���\V�}��\�PăSv:��IƓQ�:vQq���d�.Ϊ�"s��nsol$�y�M:qfiY�W�����y�GW9�r-��\�}�uG՝�U���>�v��q�<G3�����{�Qܖ:J�Ӽ�	�ٜ���Z�}8�Q�,7���v���~{�켼��8Iw��J�:|h�=I��ÚMj�Q��hG��il��A5�)L.��!���20,ؚ��(��� ��!f�|I���(�YQ�e�Q���%w?}�%�ZJ~vŎSx�r-\ſv$�kU������pm�L=Vt��ƍ0DOŚtD�(Æi��Y����R�B]ͪ�"n�I^�r3�c->m����|�m���M�����}�*��}u�'�
�>�k�]��Ӕ��3_������E��P����j�:�r'?�'%Q]���r})��q#��
��b����o����+���Xx�'NLG_����'�Y�0�D��:"P�a�4��,��ED&���|���ϖ�a� ���K��G�#�Fj�B$Ц�����Y+�6&�ݒR7q�����O���9z�9����e&Q��a�Y\0ª�n=�Mi0��~��ix���Ǫ��\a֣j�=S���,�2Î���q׮���Ζ|a��ǎ8x�|�T�*�"v��8:�t�6{���B]'+�珨������iLf`�~�/1�c��TF6n������	�IF�5-�ܒ~�z�ٖ=]ib��W&c�� �~2�WۘU��bJ��,�a����p�Z��$x���˳/��\jn��Ej7�1�q���G�N�(��(�� ��K(A(D�f�Y��Q�h�i���,K��0�(�D��"@��0�D �"p��"X� C HHA8(�N�@�aH�B"P��'D�D��	�;�<&�a��	��i�a`�,L�bX�%�1	%��I DN��"IfxNA ���H�A�$�H�	�'���<"a�0J<$=��������x�;�!����=���:߸������kqo
�����C|����}|p��e����6�%8�qE���=��b����7���_Q����j��w�>E����ծ�/��t̹#O�ԭ�������2&�$3a�M�|�vf����|���<�;,0t�œ5��Mr�L1��ٽ,�ީ�Ǒly�v5|�f~u�N��dW�������}̵�;y�Ȭ�t�V!\�QL��ww�ӼSrn�ǌm�y�x������9�S�rk"v��[S�W�;d"�VH: RD4��h�4m�s{Sl���w�5S��J"X���ݏn)��YdN6&���'�K�N;g�/�o�-������www�ww{v����V���������n����w��4�MK4�BQ�,�K4�O�Y��Fתb�d����=v��Np������s�;D=�N�#��m�Z�8�i���n[�<�Lu�v�)I����d�KH�E�dk��&+>�1�\c�9y�[��gq�.�j�cttpvF�\��8W<h��Wk��'7O��-�}�ݓ�����[��\���6�c�����0]#��M�k���!>7&��ù���V��.�v��Uc�t�z��FI��R��]���7X�Y�hU�r���iQm�?a�p�%�+��q���_4�QV����q����{qp����yy����l�p���e�[�Rj�^^�wA��k!���l����O��}��� ��r/��
����ř���N�w9>mk�����NH��X�G�ɘԐP�C��+�쯾.�8NY���C����њ5I��{��sv�u7"AdE:a�%ѳƄ�V�T���7E��J�8&�i��]�2�nQ#I�Z�A 4�V�!`ga(�0K�����h;F�hHw3l��ִj�ڊjBu��{j:՛3{�dּ=?��2��L��h��>�o�e�]�I�:����>q��4�BQ�,�K4�O?|D(�����Q���%��J�VXX�t�ݪ·.�|�X��v=��+J�d��0�UV�b<e@D��j�5�.��F�kLn�
EFc1%p��gll�>8����b=�����l}P��VAb��s7�L�Q��4��8a��h�Y�DJ�8abif�i?\m������8����_,��1��LG��t�l+��Gv2��lNJ8_��]�N��T^Z�t����V2�I~�a1e�\�e���Rn����4p�!�H{w��70��*�|�6�Ua8�r7/�_8���a���^>���Rx��"xDOƈ�Y�M��:x�㇏�� �t�7�UZF�n��W��9G��F	ϓj�{�1�8��F�ř��^nj3>��p)|lI[������	��g�FQ�^UA>3ԭV}	��ti�hXF�'�AhK�ZÑ�F���va�nx�ڵg�c���0����d�i�m?>u뎸��[4J�0�bx�K4c�ܘ�j����X��	4&�Ҹ�"TL
H�劊B
��8�� �+-�����"�S�'��ɹ�+qs3�cŎg�.��V�uw�X\o����Jբy����{�ޭ<��n1�@a��^x�M|[��չ���=�_���^��n���N�f�
*Xb��L�ٶUw���ɥy�؋窵�ϋ8M��'�hD�D:>����3cX�+G����j㳕�I�eP���^���ȜBӚ�7�����^���������4WG�<a��'�O�if�4J�0�bx�㇎�m��Lڪ�%�R���|u�Y8]}^9G�_Q�uFe6v���].�'��K �SE�bY��&�Y�7R��N��]�{�.���f�1�+�MI���Tj�r~�E����[k��pĴ���_���+���vx�G���j�֝0�a�i��4J�0�bx�K4�R&�]��9��� y(�QZ�c3��H��,�Q��+��hh�1�>__zzҵ�����rm����(����8'�勵J�1��Zl�8m�ak(fK�\Mb�Dг�(��^hM��|f�م��]O��~�y<a�d�1�.�mn[Vc���fp��DD�:h�%a�Λ<x����K$>�D;�V�,��UZDs_���� ��4	�%}񔉡9�ղ�컶�=�0fY��d�ar���ؒ���p����j���Qm�ѩ�N�l骺0L!��d��h2�^���s&��7]����6�z���2Z����0��ɗ7n�W]���}GH(N�f��i��4J�0�bl�㇏>��$��9��F��b�,�k(�i̬%Eª+n�^�,�5�r`��Nw���)���;�Ko���ș��?�v�hL�]E������Vd8�4��sH�<Ǎ�Z����"�j�m��#G�w�k��z<�y��ߴ"�$�cw6�g8(�<�����U��<��,�?��Wdb=beT�ͱ��n�|�'��k���*�k���߭^ܵ���C�H&|�=M�g�C���6o�,e�wt$ �P�H`�|���ww%0nTjHl���D؍&�������	:t�i�O�~0ӆ�BQ�,Ox��$��U�M�e����`�(�||X����ؙGo�p��$����k��٧�`f����.W�^.���7T��,�=��n��^~'[Ǒֲѹ� '�2�3�1�,�'+��A<!���Sf��tQF���N�Wp���H2"�ި��G����	�>T��h��~zu�柚VZq�~8q�x�$H8"Q�<"YB`�a��i�4�N�X��H�GN"#Q""xD�8$��D?$$���K8"X� A�$�����
$� ��E�$��""pD�8% �$�&N��M4D�4�M,L,ŉ�a�,Kı0(��Q�DH�'D���a�H �$�H�@�	�H�	btO	��X��`�	�xK��aĥ2E��������f˙�"e���q1-��s��k�ˡ�Dc�WHq����{;0�E����1��J���㢙�k���g:��l碗�﨟h@A���]�Z��� Q���kY��+i��2���T�r�������6\�b]k0�vr=j�T�s{�s��?^�����������������ۻ����wwww���M,�MDM0ӆ�BS�ͽq㮽u3m�ʬƣ/���g#2�u�H$����]*z�V��V	��a��'�D��ps]�)E�}&dr�����]K��~_ˬ��<~�-�l����~�y&ZW���X�nT���z��tp0F�;D?O��շn͉�i��F�<a�Ǐ�%�i�D�(��'�4�N�91I)�^�V��2�FU`�SG�4}���S3��>1�27#B{�5wzn�:V�V��L�n��')0��c1��?f}Ʌy�n�U~:~v_~T{�ψ'~%|��[6'*���|z�w�9R�����V:�\>b>�įU��#%i�:��ֈ�f�p�J�0�x�K7�T�}2�n��F�ϣ0��M*q�l�9j1�$�J�js��V6�Tn";�pZ)4Y��+ʵ~ �"��X��{#�����2��
>(�,�E?Lş{����(y���k�\8�����Y�-rLb-�u<�����9�t^ʢ:�=Z�xՙv��;u�����^��U4��)8@eZX���2ڶ�ek��-��,~!�=o��VL�aym�ΐ� a�	��J�_�VeP�F��S�L���9:�}���̰�4�y��rpS�S�hƨ�\�1�,Z���O��fX�����x�OiǍ�zi�%�i�M(J0æ	�M,����\д�fKڪ�'�L>�j�5Z>W�K/գ�r�](�'��3E֫��Y�OQgD�� r��6���K޳�nX�[��L'�q(�"h���I����1�Is�������Q�d��u��\n3�嗢e!<0�!�_n���ߧ�>���J�]Va��[q׏]q�Y��4҄�:`�4��<r�!�mUi�X5��:%�Oѕ9k��1���vL2��ڳ�W"����$I�:l	B'�Cd2�����rߎq�}.S1��[�&Y�Z������g�w���~�����ZV��1?O��/��0lÔ~0i,DH���#2����4�`�51�Ϟ:��\qǮ�ᦔ%a��i=�~&��"��qUiTJ!���=Blj�_�4��v6�}��* �"ع3�l�d�lM�Z��2|'�U^���J�#MŏU�g���_�;*iZ�&c���9���u�cҰ��œ_[u^���v2ʶ�,3$����j���^���<a�&i�4�(��'�4�>.Sd�k!|F+~�EZd����T}�'�(���B�IF)kj�\+���}�!�Β�W"l]���6u�����|8�9���wv��߻��c���NϮ��ů=���P��,X��2<�w��v�aǪff�5ֵ������St���(�hM�tj�V�FT���k�#��w����Y�4B��5Z�(�s헓.d4�hk�eح�J�0�1�,brfI�;�Ƣ5ے[.�Vӵ�&Y����kA\OV��d����%讒�4K:i���Y��4ҍ(��'�8}��H�O^-��U�ﶶlŶ��5MI�L��>G�q�V��M�|���������C�!���)�A�X�W��@��|ԒZ|���˓sO������!̯��ɘ�T��V:�?fbL֘�f��ƘA��X�Y��%�iF�Q�a��<u׭��yX��&��#5iy��hT:|�f�����C�hjS�H�M�NΒeo�35Bf)��Wϊ\xf��������2YP���tv���lٰ�ʿ2m��3����b2�keaL� %�x4��xM,D�,�J4ҍ(��'�4���#�-�ydbŶ�\�#j��j1�-H���K�uw߬u��IRy<1̙�.K�Ƈ����.V�+,��r2����w^�q�r{�yl�g��[q�i�_6�i�m1%X��v9n�k��ѝ;w������{r�R�􊬪�4lٳp�������ם�y�u��������;�8u�BF���ciw����2��f\��cR�<�eK�X�"E��DH�",��#���dX�!DAmD�m
$DY�"�5D�h��--Ѧ�"����h�[F�,��D�"�#[E���4YDE��-�h���4DYD���4Z",D"�4Yl��h�,E�H�$kh�-�"�B-�m#X���&�mȶ��h��mȶ���h�"E�b[I���m2ibD�F�HK$%�&�I-,K$�I,�4��m$�D�D�ȖKid���%�q6�,�-"Y$��ɒBId�ȉh֑-&�I,�H�ibY$�,�Y�%�%�K"�&Y$K$��D��2�%�%�ı"ZdHHK4��IbD�i��X��I2ș$�M-�%�#�ی�-�%�l�[H��$i$��%��Im2%��ZD�D��dȓ$�H�Ki%��-�Ki�M-"Y"e�ĲM,�-��Ki�K$KiK$�d���%�%�id�[I�[I"ZM,�D�$�-"Id�%�H�nm$�D��$Ki�,�Kid�X�$Ki��I��%��F��4�i��D�-�im2ĉd���i�M-�M-�%�[I���,�&Y!,�Kd�&���&Ki4��$��M,�&D�M,���Ē%�-�%��[I��Kidq6����M#HKil���,Kd�����m!-��d%��B[Kd��D�e��X�,�$�I�X��KibM,Ki4�2Ą�)dQg,�8ɚF��4��2f�pFւ&œi$2ɉY3Dmi��8�$�����Y&��i$ą�h�k&�M�#k&�D�-6�6�f�5��L�ő�Z3�!���TUI,Y�s7���q��s�pDZ",�E����"E�-B�����!h��;9p9E�dM�mY�ی��h��E���Dp�DDh���h�"�-��.$[D�h�,��"X�g"E�DX��"ۗ(rE��!"E�u��e��p�h�mDE�H�������"�$Y-�"ȶ�g8Ȉ���DE�H�H�6�"E�M��""��,��Ȉ�2"-�#Yh�dH�MȚ5�����m�m"�4YE�4[E�&�"E�4k"m"E�2&E�h�"E�DZ$[DE��-,��D�,݈q��--�B#DY"-E�m�"h�E�,D�l�4Y�"h���h��h�D�dM"�D[D�dMD�dMD��MD�dH�$DYF�&�h�,��h���4H��E�dDkh�m",��""�2�,��,BE��,��"ȑm	�"�",�E�Z"DBdD,��""ȑ��"�QmB�hYЈ�"5�4YDE�!�,�BE�"ȑ����dH�DYg�в",��Ј�4B�h-4!"ȑmD"#Y""�H��E��X�m-�mDE�H�"Ȉ�"-�DȲ"5�m�h���#[DE�Y�d[E�Dkh�mDE�l��"#Y�m�dH�FM"�&�h�D�m"h�"�DX��mD�-�M�mD�"#YDE�dY�h�,��"�",�h��4�"E�E��D�h�dDZ",�D�mD�dX�h���"-�"�$YDF�DZ",��h���Y,E�mȶ��E���E�h��dDYDв$kE��2$Z$Y�"E�H�$Y-E�ȑh�h�h��YE�E�E�E�Y��D�DBѢ9�h�DY-Ȳ-D�DE�#-�"E�!mh�E�Z",�h����-�d["�&E�kb,��b&�4X��b4"�""Ț-"m��E�D[E�&E��[DF�E���2,E�-�b&F����dDYD�E�,E�dDk!dH�&�"E�w���o���ûY�պrgf��f�7�?��n���Zٍ���R��g9y�����v������ٞG������G3����~}ǣ����sI�ݝ����9oA9�����6���OW�:x^��ߏ�g>�~����N}������p��f�6_���[;�Vp�~��{��{�6lٿ�<~�a��ߴ��ɷ����7�#�m���f�y���kpo��vos~k���=o{�N��l���6��?�u�rm�y�����Zv>�|�ω��1�6h�<�g���$����;vܛ���3ӯ�p۰��yvrʌ������~��3�����9�8���N�]����{�׎�<~ǳ�ݙ�vi�KEo��|Ώ��s��`7���pDmD@�����i�P�A��^�c��a��M��r�12k������D���}OW�v7�X�-c0n��q6H�(�����l�C6�`�������ow��w��n���y���E�-׫��{w�P���uÙ������׾��}_��r�oOnB͛6n3��urZ��o�����~�ݞ���T>�W��՝����;��[��o��|iǆ~��~�so��߹�N�=�o�y�z����x|�������6l޼|V����|[D��S������Ws}�>��՜l��oN�m��4�>3f��Os~��m�/���i��˖��d�:��`�Dԓ�<0�a|�#�~f�<1�n�ٛ�DVZ���*��M$��ft���&$))��O���a�?�)OS��)qK�C	?�y"y!�n�1?�*efi�I�l�&�*��[�|���$H�lt7w���W���{��n�n3f��r���ߥ6��g���x�\1�?���gwx��}�y�Y�&r�~L�r��g�p=�|}��}F�dm�ל�|��o�ߵ��Y��f���S3�&��}���lٺ���|���f�c��6�O^x�G��g���n���i��>��˷����i'����n�`�sZspp�6�[�܎29}�>?��������w4O��ї�L�~F�/	�����F͚oμ�y6���'g�=o#y7�\7 �x6�.M�ݝ���S�wgo�h�����6��o������x�^9�a30o�kg-�|���gWo=����\���s3�������N6��t�upoc�u�`��;���V�Vpp7<�x<X������w$S�	�ص0