BZh91AY&SY����_�`q���"� ����b�    `                                      +@ 7ϊ��   P  @   �J      �          
    ���(E@P*��U((T�U%��T�H)T��D� �T*��D��TT�@R��  ����Q)R!
�T{��rPwwT��9W6C�tU��P*�v:$7g@q%ptY��n���   ���� 4��j��;� �8UU�� ���w`���g��� @e�<��� y�  w�h  ��Q
�TE!J�% �� n�:��Cv: O��� �p� ��� r�y ��)	x a� ����P 
�  ��� |�� ��� � �=+���y;� �G��R� -�`������A�c� �    s� (/������T*�E(J�R� ���݀>��� 8�94 :���TU��M���  ���9����PVt ��W��k���F�  ����w� ���"\ :���� {���z�� =�
S�n� ���=8��A�� '�   �| ��P�
JH�TEEE���� ����=� 7H �B�8� �X��{: �/0 c<�J� w0��z��    ]� �7� ��  np��p��{!f����� 6�(��wwB����(  {�  Z��IE"��UB��W�`��� w`w nP����A݀r-� u�����@;����  |  �@<�}�;�
p��C7wC Y�Q, � �� ݀�[��      ��*T 4    )�&��� A� @ �ʩ(��ԡ� d  �i�T�
��ɦ�2d �M4�&&�S�)%P��L&L L @���IS�!���=M4z������1�|~�c�@��N��z>e�&.{:�=u� *�e��@xU S܂�*��ȁ X�'�������ڧ�� 
��
���U ]�h4`_�HA���}��#�2�{#���o��`t��X�_Ł�#�#�Gm�Sl.��;`v��� m���L��;`v����Sl��#�Sl���;`v�m���Go��M�8e6���)�l��;n��;er���m��T8aU�W� l �T��`U����D* Gl"�d@6�Ql��d 7D �aU�.�Ev�	2��@l�`� .�Qvʣ�]���l�;`RdP� .�Qv��� l��aU�
.�vȋ�T]��0�$U���v� m�Wl(�@� `6���	��*�ACl�����` :aM� �d6�(m��D�
)�QBdS�;dD6�m��
	�l(��M��m�l���*dD6��m�P�	�z�EM��aA6��m�P��*!�@l�e� �	�UCl
&�EM��2(�����<e|`l�����d��d��a��X6�a���l	�
m��2��<���<2;`v����^Xv��� m������bs�{ ^��%�(x��"!����ܖ4Z�"���{���!�	W�v;X��vGO}���� ƕF��3"�p;���xMäU�w5�:T}�v�z��R{7h�Ϗp`��rLP��<s���:�rW���%�>���u��{Rt�K��gf���3n�3jnvI�x�����
����,��](L���uC'j��QN�:��6��O9�7M��[f�+}3�����w�5��H���K��7�B�q�7���\��$�t|� yBvPV�������Z��f�v}3B�$oT�g&�0��8��V��܎�{���`�Se�0$�mwgu�%oA�8�ͻ.(�"0F��-���j��������΢��;��Ť�Sr���!�ꮹ����PK3~�4�y��%�����{��cb7/|����� � k/zc\�:�؞t����-��p�.�.�f�޳l-��ɌK��Cz5p�!�7&��7�pW�uBqй����/�w�٘ݬ�8�C*�0m��[y�FD��-8�5y�-�p��(n��3��K��+�˸5�{~z�;����9&bȠL������e��]W�⺞t��W��f�g�d��Wφ�`�Ζi�k��g�7w+�c6Jxp�.�+�]�$�u�o9w-Q���h(o�jէ4���`�cp��2�@���6�p�X"t�����Kދ��{�w78sR�����ot��R5���=ޜ��4�.��t�yno_c8�n�;IMn�!��^ϵw:m�5�\B��,��S�y޹��>8TŌz8v7��{M�㗏`2����C5�ƹ�o�o,�x��m��էYgr�5nOoM�a&����A�ҹx�$ޙ��p���෮sb�u����&���Z%�z��p�̃��%Է�rn3���T�F�cmas�E��q.:�� �t�rH�4h�Q'�����[��^:�C�X����&�w4H�Z��
�/��؞��X���w@�v�s�]1�CA�'uZ�qSw)���7��w]�Z���0��JX��9cSs ����wtg۝8-�۝�&M���PĻ;V��F�\V��ŕ��X�:��'2���䀍=���t�w�)qpΒ����'�J֊ma{Ǖ�3�s:مorȆg?�kv.�uҝN����f��o�XqS����w.`Fn����muǛ��Zk�&sk�b@�K��5"��|����'f*�8��͝�!|yn��=�D�K��k�~+)�'�T����\%�;+sFD�0���+��ױe�x�n��'.R<�K#���!���A�[^S]�<G_.cZ1�.��.���N|�/0��d�`�F0B��/=w�>i�D�����>�׵ח#D�-Q�7Kz��m�ΎY ��[����3TP��j�!�����Q��-����NI�Ⱦۨ��/mA�*�]x��p��b��;ۀ����蜗��m�9����(F卬<�@wc�,]s{4-��F�q�1�FC/eb��Y0�泰P�n�d,œ��nX�􈌝�q��w��
�|9A�p�T�)Y;�_T����29�Y,}�ESY�O��L�n�B0�OJ�&��@G�56�׊�]q:�.����ɓyA�GWP���Ӎ�xp�w���e�{r:�긜eu�u�����2��nH76�Q��Sw+�_1�p�Gz����ҷsN���ː��6)�i�a��h����)��<�Z��˚`8yꜹb��rL�f�y��믩�؞��O�`�*�50��6���=�w���Mk��V��6��S���g�Y�gjM��vof�iw�;�{.m'��t���Z�/�] �Б�8�#�N�����ڝ�blp��N�M����z>{�WR��0/�a���۸�4ֆ}��wy��K�Aq��̵Ɖ���ιǷ�0�T�zx�D�uu�+;P�=�n)t��Y7&��P����74�gC��������ᖭ��}��hǇf�.F���w���ע!@h|�oO�����������.�q��ϖn�C s���K�s]\H �1��Û�ʶǷxs-*�������K�xy�w�bn<9�_�#�OS���U��th`����hc�I8�Γs�OI�i����P�2�cj� K��N�1��;�yG�0���qOԨ3�9���Xocɍ�o@�7X�5��]̨��.�l�s��j��罰�h&�)�i���Y
V:#��,��<���<�\�9� >�C4�m�Or��*�^��w3��ww�[�����[�^�^T͸�ڦ-VojE�z8�q��γJkZ-�9����e�ܹy-�i�3H�����޹p�x+s�/0�t�����?.=o�.��6V;��Rc�$$3�qj�0��8s�2l��n��'-[��'Gl��z���j��Z��;dV;AL&p��f��t6 �
����h��qF.��`����sw�Ӻ5�{F�1�"�ԞƦ��k��˨�>�ם&��9�;�����i�Q;p��lǲ�"�͉��f�U�s��4ov�7��s���@7���J�N�D������[H��i�fI���&���݃,=�v��G�����4�w�v]BoM���z;qU�7Cyq
��U������ȑ{��~�s�݋t����w�F�"U����n����!5�c��\^�B�Ν7A!�{	�ε�U`�Yc��'{��AG������΃����Z�gn�p1��
�N�5L2�뗵�P���nR2�gE�^�>�5α5����X��m\ݲQ���\� �H Κ/,��S9�������
��*Rr�P�xpx�!&��z8�:j�ǆv��ұ�&��s�H<�^Ó�s�r�����B0�m���f��^˷yIxc�S4r�Ύك��'3�3è���uw�O�G%$n
��{�u�t�A�כۑ@�]�[3N�L�uU�I���������@�0�KE�V����J���q������&^cD��_ork�nCSwn�ֻF�:s��8�pԨ�=���A/�5�G�����i\����nKCw��Wo>}K��Ǆ���K	ar[	ȵ���-i"���Y��!�֍;�k�����Dx,#�+��d �{vh���1+���uV\8������nԢ���|���Uv�Ԧ�v	ٷ�h�*,��Wgc��T>^����;��Q�;���oNjg5j}���S�_��k{�'����i�Z��//vn뷳�����J��&Z�m��Z �U!�Rra����bE��-����f>V�n19���ʃ�l���
ggvߓ#	k\2��ޘ;f�+�K����p�{;��95r+��iwH �	'�_v��h5�$�'�w���˜�5��D�ȁV߬����]�."xFs٧.��Ne-�6$�ws�o�AIZ;�a���.Y�h�ۿu<1`k�\GQ��l�aswsr��f�z���ش��!���zf�G@�/m�ϸ����'9��ݻ�ك���*���Դ�}���w�p���6���2��Ow�Q=�[�4�}ԍ���e+lh�	�x����ڵ��jǕZD�VC�{5c��3�����B�l�8���]��D�K	WnAD������$�!]Kk*8���
ӹ7/W&�i�}ǆ�,n"����GG!��x$����
�p��fhq�ޝ�W��6��k�Ë��hP4��Zj���|�v�\�ܬ���lFNOݸ��|w����fd�ٝ: &�7���p�edD�Ϋk�.T�L/����템�[��?6f�ӧ�b�~�D=�u@Ot��p $���������x�w�nI1�Z�zι�|~<F�ɔu�4-[J�����c�:Bze/�l۪1K;��yq�8�%ϻ7��q�bѺfp��왺��%X�sX�Y�֦s�#"d���|m#���nX����������!���ٻ5���^�"���Z��ws|�X�3�F�����ɧB��0W{�w�Cy��o���m]Q:%��Â\�/	��(��b���4C�H7r%��$���X&vE�n�Z�;��nѶ�d|�n;��Y���6�^v�a������Ñ�S�҇7#�g)>�Uݐ�e�-cF��Qі��F�j³aۍ�f��Hۏ�nR��X�ts�qqcBݮ��I�ܐ*�iE��
�K�:��$�qE0��w1(;����R	'P����V��>/.jɈ^�{���dC��Fk]Vh"i�<���ڱ,Q�a+��2��4����}1��.0j]ۢm�xN}3h�l���R���	�Γd;�Ri/����� �Z���!Wa�7��"ܦ�w6f����K4�W��J[Ǳ���MU`\�ʏ�<��D[�@���ܰ��/�vth����9�Jӹ�P]ǌ?i���ŏ�I4h}���V�X^Fx���j�N�c�y�8�MWB��I�w՘s�lZ�;-
u0]v.�<�#�&��?�ΰsY�S�l����鸫/zIŃ�@T�̓Ԉ��)�ښw�5�6�YzVF�Ը���[U�C�.h4�8uq ��-L�[��Vu��L�p�����(��%��ޜ�b���Rg^;�n�Ks�e+7�A��\��T��9����]G�>beD�V=<ҝ�6�C�n��:�T5rP�t�� ���+����.����0c�1�Z㇔��`��Nč�9��v���f�������ʳz�ǹ]i\��I��V���N@�D�i:�ۆW�'=&,2�rc�S�Z�E�V��n+j�ί��ܘ��7:׆�ү=ۜ�� x��jz�op0�3@]��pǂ��S�:!�v�gK�M��2ȱ�p�A�yw�z$BL�^iX���U��8L���Dv-�UF������r��h�4��:�`�����B[1���Gm�{�*-E�ئɪ3��u�⻝+��ʝr���k���x�J�����׍*��W:�Y�gk���{Uyڒl��ۣ��	
��j�籂Y���9{N|�l������{�F���Lq��88�87a�˲�r��z�q����'f��S���޹�P�jkX�o����Z��4�)��U�&����ԑ��Ʉv�`ӂǕ��i�f��6�����N>I<��4��D8��ą�[v��>ߌ�����9`А{����9E��CV��=Սo0�[�nF�.�͸���z=N8vL����B��ѕ����~pj�
n��qo M��Fi���:C�F�x�&�r���9����^K���N@N����{�YW�E��f��X7	���ȧ @���t��r�z���x��*�I�'��8v^�N��lHf��3S�<bsd�cq�tb��:b�ʼ�*rޖ�Q���bl4I-ʆN<�.��G�����=F�|� ���@�i��z�����Y.-ou�un�{�H�Dא�����dЪ���X~(�\��o7/.�:�ɜLdts†$;E�܃N��@�b`��1�T��9n�D�����T�Qs���.,gd��+��w�l=��л"vqV���w89
}5St���5�M�~y��zq��|!�J(��P)9�b��=�'-O�}�V�FUî�9�W�
���Hظ��6�b��'3���N�#7�S�K��<�Xp�����/9�ܐ.2�����&ser�u��FM7�o��#�!��8��D�f��r�K���9��n�3�-L�cT���<����&�U1���Gc�N7��T�n��+[�k������wY�Q��5�+��A����|����O@����Dأ=����!�4��$���u���]Ȥ�Įڴ�:%�k�ǈ�}�H��ӝ�J}T�l1s0{Uh�>�!�*���`!�}�Hg4�2&���4���ę�|�;��k��i����t��wc{���og>���h�A���A�M|Ƙ�!��n�v%l[�҃��B5h�W[�g7�r`�R���k �����k�<��c��|Z��s��lD��#yl�#�y�q�l�3�콬ɍpQw�}������D�.��z��N�f�c�ðn���v�Z��6�����,�[����E[J�xIn>�c�m��"���V��W+xUָ�����r���nӂ�0��S�8l�r�r�h�P <���uI�\�֢�Q`f���C��b���u�켔�d�a����ݍ�:�岐��nNCK������z5���4���ڌ#FV�kX�����9��g�����p4̂I�.!�����i^*��_��n'\Ⱥ������DM��&�;y.�N#̝y۸��2�4+�j۳�sW1mQ�/Vns]Po����<W�qu�ϱ�9�e����ܰ����x���ň1�L_��;���<N��~;pa����Ge{'w�y�t�ȂB��2pKa��\.qɤ���y05�.�ݞ��	{��CmS���o�����>�B>��G�o��F�z^gY>|yʜ��1�ڌ>bs>�f��O�K�.�z�ޮK��jZ��[������NB{j9�L���gV}�$J����v�b�^M'kY�H��,x�����H`�S�j�U:͢�.�j�F��ȃ�8��qV_��>�	%oHɟ���_��S�����>y��<�;�s���!Q(��U(� �)@hR��DV��J������+��� �H�B!J��)J(�@�҂� )H!J�(��J!J��BR�P�� P4RЪ������*P� �4��J�BB
��P�J�BP�� 4( -4�"�(P �(��"Ъ��(%(%�"P"RR(҈%
�"!J�4�*�("�(�4�� ���*�H�@���%"	@� R ҅ �BPP-�R�
��H�B �@"*(���`��$Ɍ�q$x@0b��L�][�ۂ�a�OD�P�W��.�<*�Vk1�(|��o��n�i�ptQ֑yV����|�F�@�Q�:��댝v���:��sd�)����b<q�^�	łck����{F�>�q�宠Q2��q5Z:0�V?ϝ��x~s��s�Z1c�7'�_����@D�׾1�>r	�_S`
�/��?��a�w���|�X���9>?L�w�����g9�R����{��>����5�a�=��/��R���q�5�px��{����B�숾���<+m���T�C��_Ȋ;�U��[�q�{A�qy���T���i�kI�玭���n��~�f�N�A��8�h��Ўz�� �F�%�}����]N����丣8�>���br���B2��`/!�ٔe�b�霫��q�ޯ8M��6�����W��Iņ՚E�vzo��bw���h���0�IG*��!�dۙ{:�B�.T��0{�=U�{��՗w����`�ׁ`�/o��k�1(0blŰ�A�#�v	�2du\�NY�k�2xm�4P�i����7��4z:�+t<�6�g����r���Ԙ�GE���Wg��>�c�ͬ��K�V踈�w]ך*��t��;�l�+�����W�f����*{�w��d]�f�'���z�2��.ݡ���뻀{���_\�=�|=Fz��`�Cxq9�r��o.�謞<��ѝ�¯}p9����`mr��Tv	��=���04]}B���x�����V�f��i��>y��Q���W�^��o>ջ㣄d^�^� xD�L�ViX[���t�ờ_��.�e,�:��K�|��<�X&_ь�Gq{����/I��L/���ۺ�^8�{)S=�so���y]�6���gaA!����3���,����`�"]����*�g2ﱂw�`�������3��w����F�{�e�������N�
Y0ۭ��wf����\��W���I���%��Y/o9wܷ�֪�� ��}༫��r
l����gK��7=���na�ǹޝ�=���>�x������!�����|V�?{Y��W4���{-�;9ѣ8���D0�y��ʮ��u{g�g|1�1\�E�a�64x���,�os��"FUd����{/w��*�Y|[���ǽ�|[I{|���&�[M�,��wE�t�b#z+R�9��-���{�}�����Z���g�=�1j��罹��[��{r���,�Q��v�o�ww�<�='�Y��=��vm�|�J�a�$rH7{O}����Z���XiQ�?�Ϋ{(�z�ݱ�\g��LB�1�������o�Զ��1RtF�P�5���4���O�˞t�(<V?d �3�H<ΰ��C9�����ZKR|<�a�^,�7�R���o?l�Uݬ����M؎#�W�t�C�er�4<
+Q�p��c���7��npx�8��3��0�$]�~�a��vY=o<9�����l��1TFx�ӯQ��<�k��^�Ĭ]��N�~�^��Ov���kFZ���[
����pE}`'|g���|��uȷ�ܞ�Ԩ�/85�zf�����9�Zz��d�^��U��໣�F/���^��tt`o1�E�l$�b��z��8���U������3؏��^�����/��s�.7��Y9�=��|��3Ft�a���(	-T�7�ܘ.��r�����.�T]�����2��o�}>�����E1d*��
.�au�3��&\��0�b�d�`�a9����=�/!���ፃs���1>�hD���E:@\Z�s�E���d7�i*y.�(|�t�ç=n��3p���+P��q����,�/���jg�xt���{�����vo��4g���(z�k�G���op[{�������3�����p���]�=��#���Ow_�pv{t�E)�|9�A7ⷂX �k�_=J�nL�������Sg���?z��7�w���ʝ�g�{o�S���.a(1�p��Ӹ����ܩp%�<��\�O:��Jѿ-��#^��c�6��� �(�����C���e�hO��̓Fn=�P���/g�7S�I� ��Rj��v����� `Gw/���K����K�f�x���;�����=�uI��qp��.%g�l�)������+u����������Hk�W��5&��:��L�n��Ie��8ǰ�+wo�3fF�������_@d�ww)��ᆥ �U�I�f!�M������o����Z���� 0�7�i&>�e9��ooš �N�����jh�w�\w��Hdc��^8��w�Z%KN����!�ۛ�f�S����l��Km<��<��ڥ��4���?<�v�y��yvTB�$^�#�K���o/� 8�s\�7��iɹ��н�1���9ݴQ��䷺�ws���}n�Z�03}i���㍿M�z��Q��^Y��8>���-])p�ʸ��T���e�ԁG�W�O}ڤ�xNd)ܽ��H\�mͻ��5o�Ly�2�Ñ=��7��;9M�胏	��X63x�Tՙ��c�RZ�W��cCJg�������{�2cbv��s��{�=~u��{��a��#��.��Ɉ�>����ȮD^���1����g��Ya��)K��w�=�_0���N���	�C��X�K��}g4p0jo�2�wz�/L��'yzc7�h{���I ��P�W��%�61��sve����y��C�=���'{S�t��4��۳۞�:����e���*1<Ϭ]�e�Y��
[&�T��S-� ����]3=��KQo����j�}@�J��6�����1������z��{{��WG1z��'5�7���b�Ł�C�����M�W���e�ѩ*ͷ"��L��-�6o&��˷'�n����o��W�Ŭ�����O
�[�K�_����f���E����|�o����_>��>|��3��o���H�-��n�#�c<@;�vx�u��0G�?9Ќ�P���s��:d~�n��vv���7&��<�z��ٽ��5�#8/N�/	��>�Y�-���;�����Eo��W�]ң�'��{#�����KC�^y���s�b�%�F��y��h��G���|qG�4���-�K4w�r�;y5�8�y�ݲU�����i������c�k�ykW}�ȫ��Qw�O�|�*	�Q>����<�!�:L�>�=��ض{6�Ox}�'�ZDq pb���$Ѿ�=����=a�s�j���{��Nw/�)1za!��Wi�"�K�xOr����ǹ�~�O�[U�W�g����x��AZo���^\�zf����x;�^�X��HB�P+�속���	6!A�=���:5xC{��
��"�<j.ygI�w!����'1N��gu���M�w�[��)0F_h�PT�CH���b�` �}�	x�=[���^��/�\�L����Mev{ܧf���]9ۻv\�X�z\/��B���g��N�e󻚽� G��bez��3���{�%&(M8h�	v�{
Ƴ��R{sg�!>���*9���w�&1�Ͷ��h�k܁zޙ툌�-��)�r�!��Noo�,A���x��oh�ɗE��b/9��L�+R}d��/۞�t3xq�bf�i)��IY���3a_�������+ӽ�m}|w�䜖N��]q�{�w�����;O����������wnp=\8}��.��ֵj�1f�FQ�~��7 ���Ǉ�����[�����1��\�t�kF��ol�#�Z�IR�G�tP2�Y�N��wA��.�]f����B�~ó���X&d����w�?"�{ҋ��E7��,�����Bh�~��*;��v�~�⨒-�Z�^N����}9S�47`�ZO��0�61P�Nc�/k�?v����s;/����m��e<9�跍�R���5�{w; �z�5���9�����dG�{�	����{�g��թc���}���Pb�,a�z-·�(��X^�P	(�N�`���n|�L���稿b�HU�T�{.�����~ɤ=F���E_^��"U�a�A��M�e����׻YB!�k츢���U�__1hqhƿL����G_m��eU����M�>\1�m!�zd�"J���f"�͛������=�����/�Q�ͤ`��Z�I^C�9��#�=�A�k��·X����|]��AL��Գ��}�݅�CE�H۞}�'���_N~w��d�:��{m\��c9�ӛ�x4��a�K�7q�8q۵�tys�4���*m��
�SDqb�{�k��}�N�ge=6go/���N��{�F|�����,ja?�,��|��u�"<�w�)q+u�'4+���K�n�K�@T;��/�z���3�yz����JK��w�(���>X)�ۡ�cN�K� �<b��x�-��&�8,N=�a�b����Qd��P�*h>��ڼp����h�}�_��6o)��}�Es���Q���&�g����o�ґۖ�r�������y��ZM��sY�.�>��ن��gA��
v��w�����/����t��!��Mhg�ޟ>==�x��>o�Ȋ�ǌ�Hw� �=���y�ٿO!v���,�}�o��>�B�L�7�n�-�Ӓ/{:��c���1`�X{&��$@y��_ˎ�Y��|0���2���c�:=�{}m�9z狫,�}�-����P
��܀ V������=��v@#�g����=��)��=��&,ݯ;"�Þ�ݾ� �L���e��Opک�Ȝ�������&���k6���?/YK��sc*y���ޯ���u�^UB����]���k=�,3��M�5,��c�wt힂� �>�����ߗ�扌�{�F�%�G�c�&��=���B��nk��l��';�ɧc��o��o���.posɳ���5n����ۥ�gT���ή�IJ��$���Q@I��r��t��/����Or�|��-������76q��I�������J�C}�뽩>j"�`C1��/ld�:�������̺���n˱p&]��>�g� A�˻�����dE�۷���{V���#��wǸߚ�7@D���7������(���v�c�ݼ�2{����\
��B�f4�{�%�tm�4�5p���s��&�{HYW:g�.�:6D��GA��oQ��6��y�� x���i�T/5�G�i۫6x�OC���od�-[>xC��v��}����{'��K�!��~:c���G�p�K��ʱ�(���-}w����&���	-y�G/�,�V�ܠ��2t���ͧ9v;�u' րx8:�5��n�N��;D���^Ӏ���;����v�o��E�w7|���-Q��6��gi�MzQ����w�sFl\�u�\%���{����r��y�uw����ZW�ޞ{8�>���.ii.������Ƭ��W��כּS�Z6{�W�ǝ�}�`�ہn��j�&�vh���<p��-���q�x��qCo����sE3J�b�؀�t�f@�t�_+�j�S�?Z;)P{��_�ãG�3��*�s�3-
(7}��O{+@~ر�0&�kU���:zl^��u�<~Uc�_y����wn<�|��'V�7<��uzdK�rD�(��4��}�,�4��۲;yx]#���n>"f���y�ƍ><�s;�l~��21?{�����~xU���w"h�h}��0���7o���}�����y{ی���؉^�E�ֵv <�6N��}�{�=��߸`��{}v�+ނ⛄n��q7�aཌྷY�^�^[���b뽇7U�٧��'���@�}4z�aW��.;�O���ٛc���j����r��K[;��t���;۞�O��yyB���p�g&���� �:n}�O��g��w�3ǳ��{g�m}��'tm���!�]���c�Q��lǇV~�f�(n3��*���F�5��M���'',0�j<�Hp/�a^J-aK�|'���cc��m�=ㇵt볆�4�I��G��%S����Pf��7٦&�в��8��@�]A�3lG�ٚ����u�fs�{����6�v��LC��d�N��.��ɟeѻ"��ߦ�J�Ͼ�s�r"�>�q��==���~g��'��ʎU��Tj�:���Ʊ��Y�Y��}�  f�7g�����lK���o��F�꧂��;�m�	�&�5�v_>^x"��n#�ǁҗ^��/�Uɭ�ڭg���z(���i�ýڈ� ��}��E��1��t8u,x��'����_:�Rw.��w��v�]o9/|���>߼��Nd�C��nL` ���{�,za��d=��X��W��C�b
�Մ�(��>�|n��`aj��y{����<�_L{���Їx�\�^��M� P�޻�n+���`!�eߞ��]O}��alCfM�ʗM=��n���e[������tsu<GJ�pyԾ+�ɻ���������Iq�h��|��n��a= �xw�u<'o&���5�t��r���\��Z�/g�߉܉�G�f�sD�HC���K���_ oy��3�W�6���s]I�{�'��腸��g��o�WZ���ڃ�U�NS'Nw�a����ݏzy��gon j4{���|��q�7���\x�U����i�޷�*�w�q���[��7O����/xx���$�<�գs}/��or�G|��!��&{�C���=VW�*в.�Q^]��m�у���{��b�7v�W:��3�y��
�"�7��'�w����o��U���<ST=u�!��k8��GMv�ۅ�ُ�-��{�f�8#=��ǳݻZ���<ͣ=��3��� kl��cZ/������K���#~6�O�̓�V��??Ot|q�o�ػ�U�k�(Hk��Fi��2�s��R�=4tݻq�*�h䉜.��_�d�T�k�|������O��3�[V��J����|�nW9a z�4���wwx�l���I8��>����� 
�:�?��~���ؾ� >��~��~ח�����?k��8g��=��w��J� Ϫ������v�O&��u���Y��60�g]S��.:�0��]^�p�9ǭ������Yz�MP6m��u[I�h0���:��Mj�m��Ϙ���/A�qø�v�s�aCgI�ŋ�U�@�n3��Cu^�O��N�ԧnr�Qq�C�S�9[�⧋��%bn��$�;�s�3ڻ$1�b�=t��s<=&�̠���շ]]�<�uwX���N������GWlZ*��k�y��mn����KuϞ����[�;&M	S7��nCbY����,ۈz]�<�&9��z�5��T���sP�7@�J�@K�UcR�B���M7X�ac��W[��I�F��FͻJ�H�)��v���)�E��MR�H]4�lp�W3����=��v���~d����	�����U�t�n]v[����^����`.aS��w;a��t�GC�n����UƯ���zK�툍�N��f�k��f�v�pHb�:ˣ�^�[��iH�K0�9۠:Ղ�g�����d��68x|��CT�� k���|���e�ǱupZw�j�V����ƞhh����n�4��
��b������c: =��iʹLʛY����
���4\��vb�aܑ�l�/��i��gY��tk�a\p3���gr�����fNf�1T-�T���EB�5���z�����[n2�R��!"J�mWmfz�1qqF���z7V�R�`e�zȋtN�=�϶������u�hر�ͷ1�R����T��3�� ͵��p�eA��Ș.�%.��siO�a��[��t7i�G�7Cn������@�팧b��oY݌逻c�v�ۀ��v�%60��v�=�;0'�*u�5/cWZ���P���s��7;�!�!���Fj��ݎ�pu�<��|#�-�y�H�%Bd�W4�oZ��:u���M`�Bm{���5yt1�Xf�7�=�8v��=6����K��C�J�7\ݴ�u�ـJYz�v%�O�@[�^n
姷c�����F�cU��3Mzy�Zk�RG�#c��묁묖��kWB�n���lbe�e;,M�:�\v:䅩4��KCmX��sm&#�t<pO���&��v�c��ۡ؍�����nT:жXgӘ�j��<m����zVݲ��ACi��[$�E�/gJL�u`bR �n�:A�q�pې��9	BպibZ]u��Y�)c��ų��J(��-+�l�]��/OgQ�����£�R���@�6�4eSY��l�!-Ye�.�Jj\F���0�oc�5� ʫ���yz�Fĕ�@�!{غǅ�0�pWS�6r��jF�Z��JK3l�"u��t�b;��;M�;\���K��Z�k�Xh�Im�sd&�.,�A�V�ic�1�W���;��ĀRf2�k�����OC��jp�k/�w�o�Bۂ�,kNqη��ѹ������p��!p'tٛ�)�7BZ5����W�7�&�#��c����`��;����&�ٖǮV][c	�
j���5�tm�oW:MH��Mtݦ�\�Zg��<�m�(y9!F�v+E1�n�=m֚6֌Nt��tGc��t��m���N��'�v��-�]=6�W7Ak.��LZ��tc�iij�jk�%�0\S��l�ͷTgb�W<G'"�n<]e�'�m�`1��M�VIlt3��I{mװ�,&x�
[�|�Gm�=���u֘�mn��s;�}��)\�=v�P�B�L�@���>��6Mt��l����.n����A�嗜lp�!W���4�ꑱ�b�[)�����ؑ��{	�Zh�5Lχ�M<�m�R��Pv��Z�X[����!(6�{v��C���q�0:�Ǣ� D�n��u�nP;]T$�ɝWb�q��>�>�;&��NRmє�v��d8N�d���� 8tB�M�f{8�ڳ��$�׌�YA^�Ӻ����s�[���Sa��{7�㶵�wϐ�7�P�'���)�|����87jN�"n�:!50ʲ��(m4�쥩�k���NCu�!&�p�P��nǠ���֮�ON#���f8���3{]�n��J[�e��kak�A6�j@A#��`���e���v����%�T����[7e	��ܚN�h��64�@�vZ�ű���'��9����;��`�	y�-��o,�a�k��没�q����-�ݪ�+\T���Z}��î�7n��v"������]��W�`X�KJMM4� �K�����n��F+�A�yz{.m��%,1l�;g(;,�e��3Ɵ\��X!��Z{j���R�W�͘���<�KGrp��[nlt�upk�(��O�g0 U�2�pGn�$�6ۙ�b�����נ�q���4��Qxzx�E�Oa�����qOmp���B�qq/1(��֔��3��)��zҜ�=Mry0/"��w�	ۂ�c�'�m�¸-m����cn����x�Gӳ"*fv�������'0sN�a�-G`Sv�e�7f�x��06 lsϡ�ܹㅎdՎoWC@#�.�j��,)��\Ya�iq-y�!v�ny��<΅����բ���1���i�����wVQݞ�K��Yz��\�s������\.`�L��XJ�����=oQ�vsk/@<��X�d�Q��c\j� ���y�L�ǷZ��p�W�LFb.Ê�iN�l��Ck%l��B񬵄�ĢH\ea֌��&��-"��+A�h��#F�	l�@丁4+�MwuT�Y`b�]�kx�k��jKi��氅�F��6��q��v�/�`0�E9ͣ���7<Tc�,fg��:k�c�"�Э�֮)��`��6`����-���D��l�m��ۉ�=�.�!,����Bmtuh���
��Ը��� D����l=e!����l�%�С�,,q,��{j@�	�@�e���6b�Z�LRѕ���M6<�<!	l���k��4&��\�L%��]3FPa-v�m��&���n���e�.;���*�-��ݹ��i�+X̏\�I��n�m��ݦ��7O����<�ΨE5G��ҁcF��������[d]��۝�r*���&�Ϣ��FM��@�mpY��cR�#�8�;ss�-�1�֍E�[���\���S��F�Η_0����������&�4�\;�D0�-] ��ד��lk������"��f�A�q�k�o[��I{!gGmt�H��s�͑g0�4qa���a��Nn�㮸��c��q��r�Dv^���/�=;�ܖ�m��:�OY����6�iph��{\aǲ��F�梌��\�km�� :ӭR�옆�%Ԃ�_	�/�ҭ�
�Ҍ��d�'�8i�"�ܥvݧX�l8}R�Wf��M��s�#�Tr�q4���J�1��f���Eh�Y�͛��Hu�F�2�;�[R���+CYA�3ru��?��
�1GX��б��w[k�r��ȚA��Y���0h�����ґ��l�.�(:��MA�I21�\UM���3���#f�n�WP���vz;5�v��b�r���fx��t�AWYܧX��<`�HM.�2�[Al�#,����VG�Ӹbs�:�If��Y��r+"����@��ڐ6�Ɇ�)ú��2�:�V�`ظ�� ie�/4ѓ�l�؍͌���tϵ���f�K(l8�p��/��۬_8�n�t)���x۵�v��n��0��Sq�����n(u�L>�^��]n���<���S�Xf�/1�p�Q�S�(u0�na8fx��7O!�$Ǝػs���9��<�����n�Z�`��9����j���3�]���ήg�=��������-�v趖�����'^�q������ax�<�Brv����V�3͗��H��װ�l��a�N-��z���r�7U���� �6;uW[�m��]<�� ^F�c1K�=m�M��fXR��f.��u������<:��f�-��uzc7pz���H\�/#�@͓KC�n8�m�K��0�=/�sZ^Nj�n.S���5X�Z�U��a�`��;��ͨ�;������v�i�&�z�э����y�l��O,�F�����mIx�W��w\^M �\��甘��'[�{t	�u�T�Dz4��
,��ti������(�Ї�I=����S�њi����Z��X͌b�4GY�5�ղ�o.i ��-��[d0�a�Q��V�\�m�c�n;z����-��.�KA�*�4%f	X��9��x�Min�r�3n6#WY#��I��<6Q�/��ѣ�Y�t"�ۜ�,��iY�[G�����/H��m��N��,�ڜpI7:���mMB&�{R�+E��1i�慦3B��s ���B�z�3���&8�)U�1N훈�x�#����p�e�^M�� ̦�Ӯx��xg�9ɩ5�B�v]���{9�Z�f��U�-��U���]�9��V��oU�hǨ���K�[��6��`��\�J����lw	
S��=<8!V;pz�=���q�N���u�[%YtM1�>Vc���̣c�p��8N2�zz��m�NN���Bx��0�X;�<��F}F��ݹ=q�yM�&�k��f2��<�<���5���d���N�����.�t�!�qoMR{M�뇫f�JI��+�[-��G����i�SPsuWSx��mUUUUU\\UU��	&�<�f�d�L�ˇ��+����ϺM<�ZV�"�ylbU͛u#�������ȒNO�w�9(@����ma9�vv���y�^j�mi9���/��>݊pHw8r�q@�F�slHsm��C�B|��i}��ŝ�j�@NE�m�f�{Y��R���ZvL{�zK{xα8��9E)"E)�hJG�YQk�޵�"C����&��vg9	�B<ܛb��;k�<�6�۳��}���i@�@��g���p��W��W2ʒYhBGRsۼ� �2�pf�-��=��#�϶ 요fG��/D[b��':JI'%%����6�m�we������҃;;k'̗�e3G��I�IĔ�8�q��l�H;-�v�G=��s����[c?+���ǹ$���|����bۥ���XS,&���b]yks�y`�hֹ���B��5�Eܶ:�XZ���s�\h2��=�ѹ7j�9g�vΦ}��5',1�uۯiLZ�6�Ve�� <�4��>��ysa�V��`�l��	���=��#h�ݬ�r��^;v�1�W;��ǜ��\R�bd�6�t�sȝppDw<�A�M��<�e�ڜ��8�=;Y�)ر-���L�5�05[5U�%�˦<ac�q���#Q��	 qml㵞�j��K�5K��xa�zՄ��2��n"�6���i0�he��uI��1�Y0c���Hѡs
�f�c�+�M���Su������XӤ��I�]!`-n��E��bʛqɈ�J�qڙ�%�۸�VŎ��1��rkWb�E��Hjcָ=�]���ۧ��g[�s��Gj��!��ڴm�s�ulv��}$u0��-��,.2�-���V��u�*�,��d�����ю��^ׯ�� �s�XA�Z��fсm��R5��E e��)��6��ͣɐ:�e��^2a��&W�SS�P�%Ғ0��spj���bn�j�k���㒎[P��X�׵>5����r����!�n�s�m1�1ٌ�퀰�5c�˙R�IK-W^@,t8sc5D�6v���VM�ׯnzȍ�Bm�h+n�7L�Ǡh���>�P��豗uv�k�ےL�uE��X 9L\��gk�+�S�q5�����g%�Zս�M��q�l��a�=mp"¤R[+a��LL-���e�5�n<ur&c�.!�Qꡎ%dҦ�X�Ĵ+j��-��r#��v�es��dU��<��n���n�08ؗ�V�:e�#�{	�K�Sph��q���d�ZՇ�ǹ��3b)Ɲe��r��j�"��[��Fp��·&}��Xs�Fȭ��:����ib��H��J_"A�i�/1����G}f�O<7�vF�%�F)["�R�"֒%�($��6����iW��1)kV(1��m!�ض*��F�Nh��R� V��1RҼ�YV�^�I-D�a[Z%"�R�"�!ZV4�Ye#BZƀD��XA���"5�e��)�O��[��!�!�:4�ˌ�M��4�I���-�d4:֨�ks�˟����jϭ^���|Ƀ���^?Lm�)���2�R$�$�P&r6٫2��q��۳{Y���y���������R��t�I[�S8rZa��_ғ���0�Jmm��ݣsw�(NdZ}�h���7�Ὣ\��&	'W���!1z]L�F��I>m�c�Z��,�qd�o��ךݒwg��[h��{o��C���d`���ey�e�7�kVi�����¢-;;�-�U��䓏%*�S�=Ie���O\?�כ%"��������]�;@	k�m�>`������ ����F>�P/�v�fn5)���wʬY�7q��Tʑ�Xϫ1���=wpۏ�Mot�91ڲ��G�nd��$l��fnQ�s��W�N���B]j�v/��v�G+�s���f�CEK�R�D٩k͎S`l�)Ƿ=影���w��d�hW[�wt�sd�V������Zs-[��lO#�~+Vh�i���|)5c�L�<�W���a)T,aZ��I�Mm���{��Y�ࡅ ��1���w;/V·�v�^#��~>�awo�m(n��ˆ�˶��{�m�:�������$�֦-,����|�{�<�����֜�3U;Z�^���W+�Xu�8�� S`����q9[g�i��p�9�u�C�����=��O*�X�澙iZ���:�gЩ<���vo{߇Y��Ƌ��Y�����G�S����<��vٙ�ז��Z��5�l+��1�������q�ܗ�>ouw��x����1$�׵j���U���ʌ�8OXj��:��͚}���������q^��=��y�ޗ߲�_o���J���m�1*𶸹�UnO�om�g��ݽw��|{�R�8��wW��Y�V�[S�=��y$O�	MŰi�;�Afέ�;xpc��,���p� ��ݪ���Д�Wl�����-��Y��c��s�[-׵ROq�	����~lk ��/.ngwf]���J���z�J,�S��U� �p�{�0BM�A�حї����s�x.�A��|)5cy%z��-��[h,	.=Y��I�I�S/uT$3ʫ��s7�tc�I̬��Ka5���$����z�w݉�>�܄�Fd]�S��K����Y�
m�Nk��,��U�з�/�����/�%�-s 	<���/�uq��T}��L��i��-�W�j�X�0|Tj�gَ#d��]�3����~�喢`4kG���DL��k���F<ʃy>jU��t�^���#�*hϯ�K�w���3]�K�qsd7&+�]CZ���%��p KǄ��}��3}k�j�����74�Ȍ��Y��|d��Qcv�f�]�?���oJV�cJ����w9O�.�k3"�m��d�+�L�����+[�'&�N3��W�T5]DS=Fn��*�*��Ecy)	:S��5�79��`��I�+�����7��M��W���n���?��-�,��_f����A�_�,{۝j�هq���y�
r���x�~���ã���͖1�a���o ���@��x�[��#|\�+����_�C�z�'wK��n��z�^�>����f�9��'��0 q|&C2�Ó�k5ul���c���a���|]������ۭ۵�eq�������H.�p�+��S�G]�W<�1��ȅ��l�:�;�$�>�l�`��1���m;!���[���4�[M���8���ʱK6l�e�
�U��X�:�
�X�7!s�n����xm��qgE���H�o=]#U���dk���8Z��{~:���E֔�Mj������V�<��13�JEl�(χ��;��O�D���F�rsA})�u�67L�sb]���a��po$�'�lLTԾ蓶�z�6M+�g���
�Vf��W�St��������3X�I8J�0S=��Ƹc��t�[�]�+3"�G�[y�[�)I�����T�?�5����e#{99���Ѓ:���j
�3e��N>O����f	0	e��"[Uõ�V�^)�Hլ�lͦǅ62�7�^��v�]�F�1u;/�'�|��Í��v%����9�v\��k���fF�ci|�+�����[Ve�~]{V��M;��x&&v�6-�Sq{���p�x$���/6��T�$���ϭપ�ǿ����$�Q�oyv��C�_1'N]�X�uo�g��bM��ņa9�W��*�5�I�U�{���;S��7�5cRF�j��V�@H�]\H	2M��
T&���p��Om��2��"7¯o�u�v������Oq-
��f�Dش�V�$ޝuw��:-C<�f=��B��&����u9{���W֟����w�4�#=�����nT)�u��8�)?���vB���ǐD��X�X��Vs4��B��{n:���Qi��Ë0b��6��f+ߧ���RX"Hd�j���{��)f�3�ѭ�?�k$�<��L$E介��m���i��0lh���{�ך![�U��a�Q���Z�-��{1�$��P�Ɗ��±����z��7�;^����w�G778e��$t����3`{�זh�nz/v���c��*O���v�Q��0;̋�9�&^�T�i�Q�L=X��o$�b�fpӵ�,��<�u�P�Xy�A�`ۆ����=Z�����k���`� �x$��-zHt�_D��645Xy��e��6�U�M��ìIYzQ��:��!���^���=^�Ŧ���BڳL̤j���1,�3n|�'�w���$�ʳ��;�a�Ie9�/*��d�Ž���˯#"��y$�F��]�B���W�-�=d�e�6�b�E�#fb�oU5e+;{r�9���g���j����{�&B����_)���&����㊶	0���IX��N��j�XL��a��;��杗�z�гBM#�fVm�y�6�h�>�&<>���5'	�'}��r�^7H���(�稛��j�`����#�}�P$&�P՘�U7����և��1j� �E<�f�ˁv��X���J$X�w�c{���+����t�\Xǻ�0³\��*;n�IW*a��Z����T*j�Lf7,t��h� lf�t�w�+���؃<����6{n�x���2�Eҹ|ݣ��\��Y�;�6�u�2�w�k~����S��i̴��FsSy9xj]o�[e#�y9�Zeڤ�,ԛ±�K3��l��i[խ;�� �x$�q'%���'mK���hy���w�a�+5�I��$��5[�)�i�io)a;�<�R��ݭidne��\�����.!��'��l[���7�K�
�ئ�r`���e:a��7tycP]Nh	0��p��ԁe�{�^��e�Vㅬ$ԙ"�6��>���ݩq��U��ZBS�e6�
��0,4N �+Otc`�����6�ָY��C�?�#��Wx��-�п.6�S3VI-�ق;se��;a�lvT�6��pn�շ=�0�+b����,�B����-�h1�����P�����m��*m4���I�6��\P��ll�l�e+���/��ͱ���{ ���F�bL`�$Ћi+6�s`W�����.wM�s�&��b����
3l��K�tɵ�=q�ݘ�n�+��Q�p!�kma�k�����Hb�n��v5�W�,PLM	��Qĺ7B�˦��6C�)� -d��-fkJ1N�C<��ǵ��V�m�Ʃ��҄��$�l�l��n����[�yw;���Ź̼|���8�[%A1��v[�8������d��$t^��p���l˼LV�:�E ������mYm�4�^Eo(�Wq얼o���{���հ])��kCͣCq�h�a��뻋�l�IV
p�P�3�a�d���V�F�����^8mI%�'��f��n>]�D ����ǉ�,t ĺf�ݝ��*X�X#�L�Mel��\�6��o:a��;����3��r�jF�,���pv=~�{�&��I�
�=�����n��r����3�s��X�8�!���t�o�\���ǻ��5��4UoG�/m��2����hʀZ�s7��^Z�:��ڛ��L7�f����E��u�{[[B5��:Ld���9��4
'�Z��mh��/N^B���8�`�y$|��j�P��Zde֬�7S�m���0�/3X���.�4R`�M�l�l��T[�-h�&�>*�&�I�w��Y�2����ml,[E�M�z��\
L*OVcCl�d
�CoVA{�q×;6�T�Ł3`��2E�ڥ��9��k�hpI����X!0Z���їs��Z%4ә���݃m��vo�&�o$��$�.ruT��l�v�þ�^^�y�A�Vh♽��Yb��/V0e��]�K�jC�N^��z}����^]��N�8q��� ��ܼ�v�"��f9p���i��|��=;�TT/N�d�</ǎiS���Yi�����o_i���u�]j��eG<�m5��O��m��o��|�x�빾���<`X�δ�m�Yߛ���d��AK�kS	�z;���vP��`�=�u�ȗg��t���Mc�ƹ���w�=��2d��~��������ݛ�Q�����7˒'�n�ϙ'ޙ��FuS;�2�C�-�<B�}�_��=���K��{�}����~<�wv���gkL���z"w�<��r#[a���O���}��}qhʼ��C}y�q��6tqMЛ�_�t�K�2q|���p�܄:/�'��5�G<�c��p����Q��v����ʣӦ�Z��˹�ێ�����iok��A��<NwG�9�큁�(}�_m�6�����1-,��vm�k�=;�>��G���>zs=�����&󕇻�8q�])<R��TQ��C��컫��3�Ж��d�y����Ors7�v�����3�8{�yN�\�����>�ٳ����z�u��<�h
���𐩏D~���vP��i�i�&�d�f��{!1>�����������K;H�~��G���P��L�|Z,I�m���:�w�Ω��GG���~уΫ�|��VȾ>��뜎�7��t�}<��L4.Ľ���z�u���֠fG=�*����G�xp���<�kNu���]�{|�d*ÓT�}���.|;�{�w��=&ABp���>[_z{��{qZz���y���_;�W���gk_�R�N`�]t�2eC�������z�2٥!a��m���Y�X[m�HK,�fkcs-�{�����ֶ���b���[z��]�!-re~��-ΰ������w�6m��_����ؾݿ.���� _Om��y�yZ�޼H���l|�/���������ޜ�����γ��$��{����Va1�`88=�ܑ��W�=&ȫ�{�Ŷ��,�zy�uzw��l�<2���^|�����=Z;K���إ푂�g=�k��� 4���!DF}���/,��j��μ��U�u���pۭ�ee�:򎏝��-�'��o޳��8�J���E�YYߝ����T�|��-	�z��W�Ӓ����h�����-��Y�n��E�gy�%6�y�� ��p$���7�8�s���9�i�&�z�g�^J=�"�����<΃�Xt�y��me�ם�aCl�;�Wm��+�ǽ��}��{W���|�VQ�U%���Q�������	O�à��b�K7��%����_�V+Ȼۦ�ScF�W�� J`�vzv��A���9w �YY��|l�a �'��{�.��6�)�z�)i�͙�۬<.���yѺ�u �,��\w�����/}㠞�������8�� :q{3z�������4���]� �޵�<�����!]���v��k�%�[�(����6�p��3�gr��gV�å��� �a�u�59e��m,�H�.n�e?{�޲˙O���n��ݼ6�ͻ|�˧�����m�x,��Nw����o2����7o��"��탂 Y���-���/=�UQ��}Y�]�ȩi��x�ۭ���\��k����T܆����z�s�}Qe5�9"�oB7����I;� �*P郍]pf"Wf��a�}7� Wz���7���}��w�\���X2��}�R�B��w@��>��Yρ76�D�e��,������m��a��������=scD0n���5��H�2������>��ؚ��)SfU#af1B�c��v�k�P)�e���>��M��{�Ӭ���z���z�&zpw�xxH��X]�pEݷ�DތZ�,���=W�yӢ��kk���^3�@V��I��R`�~{<>O�r�/��}o�Ow��	�W#���!϶�S&e�j�7��/-h3 ꓾���gw=,W� v��� ]��gf!�/x��Y��{�<!����q�`+�Kn	��v����'��f�+�v��7�ێ��SuV1�m���԰p|[� ݷ��r-�-��µO��	�`����E��]��#^��~�TӞd�2�T5Y�||����x����7l�>���|.��5�2��cS�-G���r�q�c�^^�1a��p_D&��Vy��z��D��x�8��]���7p��a�7m�Y9�G6�����q���j��M�D0�AY� v�υ�>�s��{f�
��lOM*�(ɩ���e�Mm�H�;5:,NT6TR��XC'����\�!����C�n�~s���m�fm��f׺���[tk:�jO�v�e�l��������Da�L-%�-c�	�kaV��X���33A�K��,y��Xٺ��]�31x��RI{C������T�b;c��E���we��rmcG��]:\���uۥT�v��/[���>l84k��GFXɖ
���-����6��Q��!�v�j�/z�),֖�@�c7Yu���=���u��I�R�q�%{؆M��翷���b�֝=4�;Ύ�1��F��qIc�u�Jfn�ͷ��~3��>�
�E���]��-�+���j��||���jYo�6��O=E����o��苶s^,��&;��cGh�[ ���cj-�3x���.��)k����Z��Eݿ�c�E<�g;o�1��g"O+x>]?���wn��۝�b!���뾦Ⱥ��/���A ̰B́ �rn�?y�fH�S�����nn�7��U�[�#�l<���|[܌�J���;5�Ng<�`����)�;�p9M�s���oz���������FET�Y���㿃�`깗��%D[�?z�{�	V�-o	>w B�n���!U��ߒ��~�<�C;�����l!b���A�ܖ;����Y�3t�.Ai���;Ի��M������s� �cǙŚ��S�sUxc�57��[�b�m��P :�υ�"��G��ޯH���`�C����톻��!�Բ��i#�ч���0h��7Q�ܦ-p��}�A��~|C�}C�6�j�q�ޛ3Ƶ� ��s{IT�,￾��9c����[v���������A3�z3_�n۞{��O�uS��;����9�տ���ݰrۇ�2'v�.]�%)�����x~�^��V�<B���
�]7���Y&[��1[��k�AN<鍷����9����講���573,�7AW��OFu�[��G��8������M�<sG����W�t]ȳ�/-�^�EV>�up�h[������u�� 濟��Mݽف8^�{�������&�k���i�Ck�����{u��W`/)L6k@ծ���*|��w�2�;���۰pE�������P����q�m�Y�[��A�Ñ�m�<E����v�A1v�-���?^5Ĭ���0\gk^w5B��X���	�`��ۂc�ݰ��y��bP�aDW\Ex��`-����.�z�|�%�^1Ɲ子b)鹮���2ݗ��
]�Pxew	�OJ����y?	<��\+!Eإf]&��f�b�-����=ӫ�Ms�>�o� ��3[�n�� ��Ǘ�[7��0��Ucy���8��7nE�
����X��&[��x@ �C�֮���nl�6���3�n��zG�]ǜv�
�fk��`��x��;�y��
�Ȏ�w�3,��`@7ln�ufOuQ}1+�R�����X��ֶOQm�k���.�6�SH�gR�k�Mm�����8��Gcwu>�W]�r��_o-��o[��[#4f6?c�A���>y����1܂c �Z+8� �̘s�4�0r3�>g`�3�3���Te�ֵ�I���p����ٯ����;�M��a �sH>�שc����y�>�fa	s���w�1K),�ѩ�L�pA[� v�� ݸ���deT��ə�wX/z\?���;�1��[���c�缸gνn ��� ����v��ʚx�g��=�aR�����x�Z��r��Y���`�����4�|�c��׈�3�O8޸�z>{��5���A20���௽�)3��^�g>�`���]�u�dr�kc�h���뫅�����/SB��W� �lx�������o�{�n����'��Ã3a�=�acu��u��y1	���Ŗ��]3�iM6�p[�[�)���]��A񻷍���ם��+�O�Sq���@S���3�!��A��D]��v�:��E��=� ���;��+�����kˆ|���A����`���9�֧�۶!�}���p I�.`� ��z�.�M�,;2�#y	�i�[���7zoz*�?��wq7o�������L�J�����{�����xIŹ��NU�LC#���Rv�5���`�n0r.���AnW{;��/e��'�T���v^�]5k�kY�8�>=Z��k�$v�swo�s{#�?�w�w��Q���|p��̺��r�q=U�ɖ����^�مv�@���g��t���d��m {!�e�2�oɹ�g���xxk�f}*�6h�d�Af��p��bh�۲-z���"Px�R\�&�v�/C�N�3����,�!pa�z�p݃ۜ�J8�v^�v���船N�toͼ�>�;v��lti�M՘���s�Zg�C�7Zqm��F'��]����l�o8�(��Y�0��R@e���2ֻ���g��m�˅⮨踵7n���01��L�lQ)ٰۮM��ߓ����e٥���*#7�'c0fq�V�Hnl4�������߀A%��j���`�{����)��{���:;K�v�0�'�m�O��f?����x"��Z��þ�U��A�ǅ�$���iYYUm�Sp>�`� ��]�h�z�$�p�r�X�p�J�8@k��.�W�0k���{ �J�]�aD�F��d�C��7��}�F;���?�&�� "휄-�-ő�XݶA��
��ۇ���ֽ�1h'�J���U�8�]]v>��#n��z�]��7w��.��d��qB�r!�ڊ���v9�NeU�������n�8$��/�^f�КV��ty�9g�1�Ӳ5]�̍S+�H���}�f˧�wK!�z�����0r�p�"��x��8y��sp�e�e��yS��".�|�>�֒7v��.�� ݰp@���7wfa��\"�29����&�.7�Oe�|�wO}8�=0h��9�r_a�X��"�b�{�-4VS�����.�Q� ����|~�������b��;���,�w�oz*�n�]ڼV�eV�u�o]?��M-x��o�����z}��3ۦ[��/F�,ɫnM���EvD�����G�7N���&n���p�|�,$2��bFlDxݿ�U�>&��Ý�\��f7����g�a��6����g>�׏v�A���.�v��u��;x*�g��|'�����GzV����9-����v�>|/���K$�|��vԠ۫�hm5Cs��3$ѩ4�36����y��\�o��|%�z��/�89�� �����6�s��y5m�i���;g6)k0}� �`�]�q<H.32�g9���Ms�&�4Y�x������&��'��a���׈����n��9U��|�����X������ln�,�ޛfs���o;���Ml�5���zR��F�uj��og�z�C7w�1��f��g���Zb�i������O�9���U��Ϯ+��rq���xx{5H��ooZ�,���[��B�x2v��y�LǞy�y�-�x�F����_W�R`2A�ݼe���>�����~M�2�����f�:���s
��y�ݸ��A�E��\I����O���SN�Ϗw0��f7uk��� ݷ�����ﶢ.��' U�����qv�,�n��jd�]�Z1���n��%�]�3������A��a@�.�?����3�|��f��+x@Lb;E�-�������A�[��&����o�7l�n������cz}=ip�wm�m���ϣ�)�*㽴��	�`���v@�v�y3'z�,�,n�v����`�p�]�G��sn���m�<������.s���׀A�8����v�B�fr2�^E�b���v8Ӷ�}��ۇ;��N4��54Y��J��l\�'6�����ҁI��A�PۼF�L!u�FS۞���kP���>�y�f:r�3h+5F=B���k�k�z��ME��2p���R�� {����;�����n������v�pn؍?|)��/X�x��ҝ݂�����w�&%��������.���
��K�}��B���aa=>����n�v�6�6`d�n��&�3d�bkv�$a��a��~�o��6�g�p�����o��|�����V�oYۍ��SFִ�����O�ɼ�5�����g ��� �#G�L�s&���V0r�p㯰`��}�榋*{ҵ��9n.�N��߫�/�����gōn��m��ݳ�7v��ν���)NgK>�uu�u��bX8"�G��`� �dfd@����5f0r�p�"�Dxݿ�ou���G#�b^�v�w�����i�;��
�A����U0x�+�.��n��v�]N?r�4R�2n_v��E��ӭo�qw��k̇}���<i��zxt�����������3�1�:5�}�X���+N~�0���G��Q�ۻ�MiKLʤ�'gg>�#�$v�ǜ��L��ͷN�ޘ��1��ѹ�w����q>OX���+l؛=�:�^<d���.X�<��zjۥ]]�Ú�i:�m�;]Ti�c��w�i²����i��Ap�X�x����F�X�ݴ�>߼�/.)��)>��x�j��Q:{|�!���l�p������I���g�:�fŰk���wӜ&�����|1��u?	ϓz�cpv�,�ރ�=�j��D���_-�s�ׇ����n��/g-I.��+�}m��5C{J*���%�y~?��nk�e�4q��@��=t�����<`�,�㛛�N����ͻC˔�;�Bj{=��~W�"���m�{v��Յ�c������zY������|�Ei�z<�
��ܸ<T�禼�A^�������Xx�8��ns�XF�ʭ��j	�i��B�v����7�q�/�uXj]��7�1�ߊ=}���6���3� F\>�r�*a;iq��n��|m'�+���`��ҡY��W/o��ky均P�����.�.�#�bA��G�\k�Kd-{D�}�/N�'S5�ƽ�7��sGtM[K�.�����=�f΋�_�ZbM`��}4�Nv!1j-q�a��؎�-�}�y���obv���q��^����L�#a͉�Xf��{�D�W�3���x��>b�2�=.O/t@�v�>}78�C;�#�k.2'&?�<=sFn?'� 0���G�Ӎ�.KM(k����L�/oJ��h\4��@�n�^�eN��u?=um���ßü����,����Nt��8⼽�=�G%p�:�:�Z�^��P�[׋˻��̎:�.+3��^[�þu�j��
8�k	��9>n�}n��9μ���sl��:I�'��#��:F��[�+��pQ_;H�["��^ru�w��W�!J��giO�μ����׶�N�՟�b�r�Ǳ]�6��6՗��^^w�w)T ���G^btqtgfVwmlmE�rqgvuu�{�Yd�qu嗦\w%���;;+.;��Q���7o+8�������8�+..��ܝKָ��-�uI�I��vqyv�{vDG)�qv�-�Nt���TTwE}�gb���'�ge�ӒuA��s����y	��G3C����@R��8��n^�G<GA��G�\��B��ѧ��Om�4�
V���1�t��L�����۰�e�tY�I]	Z�'���|�n;��-k�))n��&���z��5�BK�ʹJhi�MW�2aqG�Raƺ�I.�^���7 �*�ku�O��<��w�Q3�uַH�v�p^5k���´L�,I��op� �dS�����vk��5Փ[K`S��)[�0,t7�m�J8��1ۃX���264,зG87j1��8��h๭���>���kˋm�h��;L�i�B��¡íѵ��q=]q�ۮb&�.�O)�ݨ՘�Ȧof�K�]b&�����a�sn�v��u��H�LG��f�,��Y6CP�+���W���;;��/��M��W�ѻMf!�P�]Yl5M��˻;g2��%�܉8ѻ-�fc���;�бa�  �n�c��^K8�D�/���QΘ�v�`&E�A��wnPes2Y�o/o��I�M�ۇ����4kmss=��!K�A��]ml]*���)�;�1D��++vc[�j���X0�l�M�Ъ� �n�VVlkoV-A4�B�k�z����u������O�1�tH[���-���Ie���"��	�Yl�`���Jr�!5�z�v���K����^���2-ڣ���k���p���s�;����u5��x����.�ŗf�Bs��qY���=H�cIG�P���a�.,���2����\V�[tn������M�ۦ�=]؇xŹ� 6��9��qg�������<��DkG v��d��d��{{^k����MƬ�v��M�|��g�Ct�415ا�b��g������imrɳ9�j/4=�;���u��h'5F����)u��E�\>ηm��7:�I4�ˤl6;v�$n�Sۍ���9v:������5��=�-OQiLڪ���F��s)���t��o���EͲõ�7c�y��R=m�hp�F:��^�K�{<g�c���.*�Gڮ]���zm�B�����@�Zf��r�4P�&Y�ˣ�`�ͪ�q��g�<�o<Q8�:��R+�m+w%m�7;�cvmZ�LL�=ہe�)TY���y�Pb`c�]C�e*�f(]��=yݺ�0<�� ^D�q�.ָ�������/��j*)D칼�glQX��!�i���n�f\�,��
���O<�Y}�y����7v�KJlS�ɟ�%uuµ��,�-���"6�@;��	�w��L���o4�.ȏ����ƾ�M�Uy٭��s�����󛶹RՅFd㈐Ccy�V��A���v����q���	�4�bjn{q�(ڞ�[�.AX��w<@��=v��è���K���A�D8+��wo��O��ɟ�U�]p��2�f��ӱ��#�1Vz�#�Ñwp= �6_�����zƊ���N7�Q��񯧇�a�^vkq�x �ci�8>���Xޏ�|����f�}�=,۫��`ҥ=q��/l��3q�p�>��"�l��8؟'���K��������fϮ�^���i��8ЊU¼J�"�/5�!�i�7m�47���E���������V����b�g���P�Sc�9�!�k���o�+y�uŰ]��D��N+b�0��{�تʲ#3ŴԦ%
�\�
�ȡ0>��}�|V3�M�<z����7��~Wuuµ��fX8 �dx@7l:���.3���l�=z�=ۇ]�z<n����s&Z�~�{n�XJ]Lʯ;5�Ƕ���7l�wo]���9��2�����	��|�����e�n\?_`훝��.T��R��[�Yb{\��1�w�H���[v�oŋ]���`3��av���T��˞����7���5]ծ�C�퀱d0�0��k΀j��v9��ٙ�3fqC=l[�Tj�Xn�WJ�j���m�-f��8z�7��p�]��.�����l���e��y٭���ԶCnQ���'W���A1v�V�&탑�Q����\_o�X;?��B��~�^���� ���|{�Fs�#wm�4Z�nlŀ�>� ����,x![y��9�z� ���uO<D;<Ċ,C�8�z	�^�rB�8�!��%�c9�gY���ہ��~��]ܴã��#Q8�#!�ܐ������x{�xɆ���S�`�Uk��	�`�"�@7l�]�p����LMQӧ��ۘi�Â/6#��ǫw"�w�:��nkp>���1����p=�7��BL�Qc�J�;b�U�N���u卅��c�%]�[�����0�ÀE�����o?�{����yG��e��Ui��ؙ|��fݰ�'u�8`�/�V�����Z?_�ߩ����-p.�M�<��c����vq-֙U���{6�)n�xq��,�6�[ �n��q ݰr37p�_X�Sʚ����Sq>�Vv>Et��m7���po��n����_��1��f���Aqv�A���AŐ ���ݰ4\Yi�cO������4d��kѐ�w�o��#ێ�̏G�c���oN-Q���Ų��Ms� �8m �����u9KC��Uk�kqצ�xVE��j2W9ށ��ۏ���>AZ��!Qz����?Ӡ+��$�3���g������~c���48q�9|������LAy���*/�%=�t�����ف��� Ϸ G����M�v�Ȼ�Go��{_�Ϊ��fN�"x\�v�Z��v���r	���-���S�n"s�T�ĝk���.��[��6j37cF��
�hBY��C8���a�S#�8�n��ׅ����2���qm�93n�v(�ma�]8�=��y��ٙ�&���������b��,�)X>���\�r6����UkEk{��`� �l/�a3�;'����X�����,s�� ]�r*�=7o�������yFp�7����[� ���sv�W��o붠|:v��t4>��a~3*x������	�;��!�Wz�z�`�'��F�(X!n��e�m Mݼ{�]���hڛR��_�{��z�����i��h�nfX9ܶ=v�/��2�QW��FEÛK �O�Ol+����owm��ι���X+����ɻøB\�����|{�Y���:�9�{5�
�������q�.ͱq�q�['��6F�a��ъ�	tH��{i�h�$�(�I�f��V)2$!v\���#hѵD�wU�^p^�g<��=ȥJ��Z���ی��@ӎ�����@��=��
���G���-�펹K=�-��v���m�e�R.������5H�l�S�����1aaƹ�X�6߾~!`_���b�a�x������,��,m��G6&㰇����Kn�9��`op#����]����dp��qyۭ�\ee��=��_^�v?�x�3�A���o9�`��t�w�
�5�d�\�we�`������7Q�Ӄ��Uo����[�"��En�-O��˽�����pA��Ó�v��}]����UN;V���S�첍U�
��Ae��k��A�p�]�@�}q��1�$�W�� �8p���v�q��dvr28D�ȼvkq����!Цq�a�� ճy��^:�%�cH ��D́�t���;d1����<^c6Y�ֱ�_&q*΁��n��G��ۙ�����aM�n�|H#/��qI�BF����э��.�S7RZZ��T�O����ү���~ ��x�/_��gwo�6����]FmW
��F�t����F�nk ��
�A�Â.� l����؛ˬ�DQ��/2a��K�&ʜJt����n�Mkt��qH}
�hC+����O�٧�m[��t>淳��K�\Abʭ�p~��� �q��0�#���g�>���O���n>���G�0���ƩZ]E^V��S��7��.�6\�v���G=��m��kzj�l��aWyV?���&���k!����i>
m+V���҆֌xj!��8n��J�]�n�'�����԰hӹa�
� �8�wn�G�v��W|�F=�Fp�m�&��ȧ���'�O9���n �X�A�6��ݳ��H����߼V�9����t��6�9�݌̝	�Y㋁vJ�g���y&'�0)n�ܶ��}�5�	�`�K\A�e� ���έnt�Z�9�d®��� c�;}��4�e�8A�p�u�� ��W�����o �l`Ӌ8���#@1Ln;(5��9
g�ڭw���R��<�xٲ�4�[e�f�m,O��8�H,[��.�`�"��<m��l�#���p�(;�˒O;��y�g{�N�zJN�u�e�ѿ�aӞ̊��_�In��y�>��c61'U7q4�#m���Z3qj����r�����yc��Hsv�&���l��@�;5��0r���p����^�:l��nxl�Uޚ��l����9�p�"5Dx�k���y����m���owr��-`�}p =I�^��p75���GN��6_��ۉ�����0o��Q8"�+	`)��s�6ē�&N���rvKv�tF,iGkil������|�Y���y����E���hwF�7�O9���5��1��.�n>���-��ݼx�6}v�Hl���p[6^����fːo\?nks��Z���
��Y�(�p*�8"��-�1���mC-bk}�ȇ)3��qc�k>�i ����s6��Z0Hޢ�x����x#�q�`�#�����ۈ�v�e��b:���"��g�3o�1�-�#�]���ǣr��1��9y٭� �X�� j�zt.�Ϯ�zTb�`��|ƚ�-��#6n(W�$^����YO�-~��J��ߚf��v�"�"��<U)���I9���,@����q�_e��2}�e�uw�Ľ�p �U��`���*E`�a^�n���Ů����UޚΏ]�r�k�� sq�oR[�ŷ=C����!�6�l=���@�z�=�9kZ��Mj�gu�z'�9��=2���G=75:���p�ψ&��<�%k��\�Y*+���F�B�^S><��v��w�v�yf�l����o�>�އ��M�nyʼ���rǏ��pnۘ�fN��p
�x"m�AX�����p.�p�����YM�x�c�<6<��Mg@&탂I�p�"��G����>k��E�К��2u���Zm��i>�o��k�v#���ൽ�2�޸Fl3�6;���L������-�`n�8 ݸ�C�P`���*��=B)��v�\>g2n��U�n� }�;��7m������EL��Vu�S�a�W��tQq��"��Κ���ǀ��'.�Z���F�b/�O�ƮEa���|7��H:q����Sݶ9�)�#�<1λ�n9�g�X)�#� �k��C�K<�n[�!����G<5���K����v.x�%Fh��E��;Xe���҉!	� 9Z�&�;U���Q�GL�v�C�uL����
su��������F�8���A�%�GK=����^j��m��^��z�^n�v8N9����8X�p����^L"Z�;p�0��eM<%�h D��Ě�]�����~B~�5'�m!� 2�Pin����g�8�"�Щ�vǇe�C@���A�`�#7A�`��v�����B׮�c���� 'ݲxc�+�� A�p�"��;Ǽ\n���ƌ����7Y��g��k��n|ۦQ���4V��S ��Z}�&�{b_�+���s�9W�0;�x�"�8"��<E������YާMQЭ�]�r�;u���x �[Hy�]�@76�E�0�1�q3�Q~1�r�Y�zǋ�E����������*��V��l�r��{a���"tp"n�<u���|n���md8�#�3�����'�=�km̦Q��ӴWw�����-� ٲ� ����n���Nl�@3�b��h\�f��m�&�lB͡Wk�����96Ct���n��z�C;7�����n�r2�= ca:ֿlg:n�����ob:Y�hKy�[a�wo@�6C����@���NKut`A�_��d\<<�1eT�w���.��&�Z��5�������� ���ɾz'�\��h�^����gǽ�{�������swٍ�:ŵQ�!�o�s�<E� ��E]٭��roh�/���gǈ&����wo$E<e��<ҰҌ�k�g���6�8���>qv�]�z<�[��\���p�a�ݘ��C��>?c�1��W�����x�G5�n�Y$O����}k[�Y�`M� ��� ٲ�7k��u\���6��۪��+�3� fϕ��wp#��ȬՋ<�� �z�e�⍦��m� �[��@�f[�ħkl��qE�³���.�;3�n�o`=���E�>�i �wo2��n5(ަ�������|���yb�awp#�� ݸpE����.x�>r2�nۉ�ka33�_�u4w�i��n���u�� ݶ���cTL!��<�a�C��Ȼ��Hn�G}�8\3��ӧ����������gכ�������l��c
t�V��f�cOh���&�o�)k�3��P~�3�n]�t�{��;���ɏ�5ۋxr�M>RN��_D�N̈́���=�]�[�.���d�4L�T���cQH�A����^�G�i�����y��Nmh��}�-����>�z�l֫�{��>Ӻ`�O��-8�Z4sۗ�trO�Ah����>9Ԅ��m�c����܋V/�h��B-S#�l�K�=ȣ��n�������X�T����?3D�����g�{�/;�ݽ��gQ3|F��F���Vmar��4r((Be\YVM�Y���ˆLEEc��9C�����������qg7}��t��=]=�=�=,>�>9X�#u�p�)�@zդ������vD�{��"���*�m-�~w~��S�?]>\��g����ٻ�1ڄ���o��u��bC��ȿ�Iޫ��>sL.�CISi쫉�ϱ�z���ٛ#�޼W7�*�j4}��Dȭ�y��{�g�a�L��a��狁S.��P�ұ�q�d/��ރ6y�~��O��f��V,A�.�t/iaW}��o$&���ЕZ�Xřsǎ_wu׼z��ڎ�j�s�'f��w�w��tz�����y^�7_���C5�k}Ʌ���rF��Y� �ww���$����o��{skZ^���B�`u��+/)60�p`|�7W5� ̓�Q�{|�Y��R>Qݼ����<��l!{Y�[<��UI�+��׳�{׼!W���5�g��@BM�������tZ /�X.��`����������׎����j8�vd)�`sfC�k����q��\�� ۨ���u�`��8�Έ� 6��Agv�Y���u���\q�vY^���m�gS�GSk��J�J�:����D�򼼭�v��^�u�%�О]�G^X��E�ye3tDIg[�QW�Y�A�w��ٝ��ړ����.��):����:)*)N�$-�,��+"�G\E�G�GG'=�:::���Tsl�.�vQPqG^u��gvw�wwygG�\]�Qt�TE{j;�m�ڂΰ���^OV�8�ӝ.+��죪��� �.����;;���E�unYեe�]{h'�u�wvXGqI^آN�8�ʷ�՗q�n���Drq���yA�A��Y��j��2��fY�$4�%���
<]��o�w5�*WP"�>�A����v��v�G������5�h�._AQoY���jS�Ϸ;q}R�!�B9�������&*g4�%Y�2w�m�r8%\�z�Ñw\��ԋ�أ����C���k�kV���M2����A5��u��&&��'��hywޛ,�z��?��K�`�v,.r��b�^��Pd^+�8{fj��f��g��|�	e�H�/��2�(��p�����6���B�Ns���٢��8![��	��v�c�]�����(��9�gڙ�W��:��K؇��f��06?�FngE[����y���o#� BLR��&DE<2�<x�<�U��4�:����Z�q���4�	I�NK���q�L�5��t��p����q�q]S�(�Nw��d� z�'�w~ק�|��#A�D^d6i~r{)I��3�|�~���r9��^��>wt��A���ٗ�����`Q"1�c;�,mwvr}���_��p�8�C���|!2!�I�5�Jy�A�g
+���Τ�*ӳEpG�0+9E ��(_b��\Ý��$b��Y[WE�F�C���nK��g����lp�vr���"<����#��=nM�QJ�/ûY�3N�:�/{m�IMLn9��ZHpV���������퀛��I7j6(8�Y� �8p;7[��6۝C(�Qޜ���ْ��L���ܗ�h��[An����?�!2>I�%&z�ܰ����5je;k��j^��sU�p5�Qr'�8�D'��QY1;�p� �p�,w�L�q+t��n{n3N�:��b������Z!��uh�5��x�E8`JL�(��r�'ǭ�|�'D&Y�ח��ΝFU�zr}ހM�.��%/�Q ,��ݹv��#*�S;ӳ�s��V���h�Y��7�����ww1�{Gk�4G��"�<�̽�*�ˋ{7t�223����3�X7���gt��[���͈��[q��6�ЗC%�5҅�暎cr8�n�q��d��x�R�d�f�;Lu!����Iz�՗���[��	�Ɋ�yѹ�;$�]R���v/��s�9zή���<����6����/n�c�٘���4o]ŋ�:��[��0�b�Hݛ��D�Ѓ�LC�M�X�g��]��1˷t0]l�G[�S�:�=�|��~�Z7b�Z;:���j��K�����k�kB��� ��c��Y.�2���b
M�&q5u��9�wkA���w�<M���T�$��������9	;���[�mt�,���w�M�8V?�V�ݍΛLӫ��n� �ֳ���r�l\�Dt]d����H�0�h ���E�)0pA	8�Վ����å�U����b��W�5n����z(Y3P#lYkE�1�L=M�l�󂱜��qKsQέ�YF��౸�n�?��;.�Cvߖ����	0�����0K+���0ӽ�|������흍ΛL�+��n ��g ���� ���[7��-cNI,���Xw�r˶D�u�C]�Xq6!H<����qmD�|����]��u���t�>�o:�ݵ�"�K���8�����.��`H����A�gW�G�Fk�g_x�5Y-�f�&$6ǽ��`��y����=�(_����,Eٿþd��h��T����)����B��Ӡ����80;L�v�aJ9TS@t�� x���|S?�'~i����b�X���c � �p��nniS8ab"�R�Ȫ8 �`��9	8$�S;�H�;�]='�M��W�����A�k��RoW�̝��H!��]wM��'�60����� �8u����N���^��\�b"_q��ȶ���v�@#������I�AI�����I���\.:sٌ���o[�J�FB౸��5� �]��!'[����%��C[�]
O�% ���Y�lF���8<k�^mָk���d�ձ,�B���cL2�՜"���i��}���I���z+Zz�)�p2��^7�N��FY�Ex�9r���X�kb�KZ��7�3�cj�g��D��0r�p���nY�O����Ӝ��fK�V��	,�ݔ��^m��:�6��7{ëQ�kX6�%�x]y��xgr�KGt���N� �eG)��x�'nN���դz2���ؗ[�k~��q����m�]~Y��{\������^��{�v�U�x�-�N�"����� ��^db����(��L=����M�E�"����+t�?lS��U+�����9��(���ֈ�U3�	���N�0�9E�_�Ӟ�zSb��8��j��}��wt��9z� ���I��C�Q���u�-�|��(Kh�\���&��3�sҋc�Z�M�E�ع�тf��޲ߞ�?Y޽p>I�Moe���J{Ȯ��g���3�{�$���� �'I����9�|��2c�lV�W?��'r����~ا��W�x�[ō�9ٯ��I����UVѕ���zL���ù��aDR`�)0�t�v����YVF=��;�Q�ޜ�nX9
�?����I��8"�\
�!ڂ�d9O�c9�&���^�m*Sؘ6EpV����@��|&3�v�Yu��h�����ʚM�p88�9�gvlz�3�ӫ��P��61-}on���nó*k�z��]Z��k<<g���^��(�Bs�.���oz���!kX2��Y2Ƶkx���KO�W�oN��ы~m�݊���R������rk��L����E��b�{���[-�˦���t.��[���/'j�n��Ok95�rT�9�y>��������Km��8r�!&}����u�����n��8�y̓�#�^��>�p�p­��?���][Iݳ��X�*:�s4���=l�������Jo�Ȯ
ہ�`�>� AI�	vOL��tb��~|p������]�pBN�'�=�n���3�)�e
2�'J�o[��x�f�����M~�m�W�f�1�/��(W?���BL׻�My�Zۙ�T�w�8����N �7у��C_/���L�0Z~p"�!����H}��2e��K2v�%7dWo�y[� �?���/�	8�rC9�1��MMZ3�=�����s��3s۾X�&�؂��Q>��r{�=<)Ć��*�X}����:���o�K�<Q*��[+;���9`,߾����_�u=WtE�z��m�8�Tr2���z��%���
7v	�u�q�V�q,���BhW+K�q��`�6�J�4Y�n̶�3
�Ś�Ghe�A��6u�vCX������c��<;��՚Y������r;��sf2�pqI�fss@+4�빖�mx܊�\����,%�b(j��q�Z���,ѲQ��ѡA�mc��eN'�SBh+��P���U�R��~�,�H�9)�ek��t���c=�=n�	ڪ�9\��H�0C��w�~p|Q��N���S"efsttf�������n=�b79�����A������3�$��L<�'�CX*��bgf�q�ء�8m�s�]N7zs�.[�.�?�	m���,;���w���`�1M�@-����5�?� ݲؤ��
]��=W����*����w���&���ǈ)8{�87.7ZVfP�ҖKf�L�}����$����7\�WQ�Q������r!�ӷG7�AƵ�o%p|T�<��!&̸ۈ���Hc ��L6o1Cn�У���q�Ӝ�\���Âp�%&V��O�\���<�L\�ř�v]s��U�<�[^�+��"�P�f��av����Yϱ0pRg�/.�c�k�z2!o��pױ}��.��8}��g� ��r�����3U{B�?W\;���J=�Uw=���P�>�}�>�']�n��	�h.k�a��i �3�o<-mF�كކ��ҁN�=���ߚ�=�=E 4
����׶�XNw��=��EuF��n7�r	Z��I�z�x=�����g���fps� �'�g$ê�A���y�=5���c]��q�Ӽ�\��v�$ޒ�y&�3����q�q��� �I�MD����t��b��FD-�{)���C2OӰ̀t�A1Âp�$�AI�z]��ax;�����r�D�W���x���+[��M�)4#QG�~o>�}�)���FZ	c�(U�@-iT<瞤ٻ5�n�F��ljkjWL������������%'�؍�p�g��Ԝ�V��r��!��f�[]�?�dC���Ro<�9�,0S5��v�ƅ����+V0��Z.ۈ')�qX�I�^e6�0�6�Ñ��I��BNR�!'����K?0��"*�y<ɛ�wg"�44��z���Z��
��;��};�
�!�j�\L��D�f\,�T-�e5���7|�ٓ���Q�z�(iV�ym���ڍ���^v�{�n���o?�L��8!&�ZU��m-�FN����q��)8|��r{Mh�vk�9ޭa��`�#2�n���v�����E����vރv�>�8)6�M�Ayc�c<u3�w�ﵦ��bhk�୸Poba ��܋� $��)N�7uZ��ĳ�0$i�L	����m�TuI�O;&�>:�d���u���6�����"�ÑI��'��_�9Qé[٫��n!8���ͺ��^,t�m�\��]�	ֱ�5�f&ְf8�8�ە���0���w��5��ٮ��V�~�l �39p/#,��x��]��5�%�X�Au�v��yr]���n�r�t�sa[N��U���G��
ۈ')��*�9I�����0)Ç���u۲��_Y�@ ��V�?�I����Gzr��U�٫��nv�G�=?bE��o���P�enWؒ�f�rm�Ȗ�1x~ؠ��Ua���~�~߱ǝ����]�[�Npz�h<V#������Z��+�)B�)B'\e�o]�$M��2Ƶ�������＇7l4Ə�46���(�lV$���֎E��Np��r��"������<?��H�A�����%���.��Au���Xm�5�Jl�ۜgbb���X�/|���zAI�I�Eh���-�\_m�!q�Mne4�{�B�sX?���N�Bw��ȉ�fD^y��3�@��u^��ʨ��v�U�n�AV�u�M��}���"��9�Â� ��]���Ѻ!���\�gSX�f^�s���Lݸrp�)?���m ��j׈nȕ�����֐|�Ep�[���[���x�pr�9�ވ���մ�A�z���F��y�L �`�������*n��f��o���.�P]�O����k��op&r]�ֱ�:�%�:p�����������v�O��z�}��Z�c6MI�Z�F�*��-s�ûWx��q���h{��|\���zeNL9�E��#'����Shg��Z=�Y5�������9v��pH�H\{@�L
0aD �Ӱy{�1��=�=��{Ga�7.q�,�_t@<��9%ǽ��M[��5*v���������]9��߹?o�kk݁�w�{c�V,�}���u/1��D���/o:y/[����-7{��(�!��[w��Ü�P�(r�l���ϦLg_;&�W�����$}��`�9Y���14�^/��Xfq����S8�7i9�����>�H(���T6נ@�-c�t��5���k��\�m}r^9�/k�2̤uJֽ�j�+��jK|���{*:��^L�8\�3�=��â��/܅C����J/l�/^<�xM;�G��� 6\�]c�v���Ҟ��Ўs5u��b�}�o�o�GE������잝0`�����=�Uo�nL��p��oӵo�q��W���̽7��F����[V%<x�0�K=1r�|���l.��vi�ﯜ��/���mY����,yv{�q�X�xt�Ԗ\�_g��@x;S��;Y��T*�3��Bʠ���h�v�_=�V�N.��B�۳(ޏ�d��=)�(ӝ��{�_�l�ͣ_{G�kl]"�����~���w�=Y髬��6{Oφ����u�#pi�=���{=����Q�X§�M3������G.Pd����,�ɂ���V����!ۘ�/����B1�X
V��c��<�_<Ӽ�޲�'E_Ñm��.���.B��.�m�QpYY�u�M�*K���G��]�9Q�W�续8�˼���;�(�B�
.θ�.���������3^����.���:$��;��8�:������ɭ�n쳣����ʣ����Eegt]�Q�hË{^�]�����w�g��vw�t�_��[�{wU��|����.�s�#��e����p��.::�W��^uiyݥIwD%�lH�do^�9�icf���5�K��貰�'8��;��mGGˊ����+�D�|�:��믙�q�|��Q{ۃ�o�YyZw̻�nQ���gQ�gNRIal,,�:�{��3�U��-��sa���� !r
m�W\_����X��X�vv[ v,Iy�T�X��,��,"F��3��z�=k�������q��r�vX���x]���WWY�F��(
Spc��[�=�q��o9�V�m��-�ƌ�D&zKvB��+����낲�hFZI^J]�ZhTYI�����KbZ	+,{+a��k�4�EZ[!y��T*6Oanx�ψ���@q����nx��:�F�;=������5�d}P��|�RU�N���Q 2��B�P�ƴn���9�
te�8��\��m�RN��i�����n��[ۃ��vM���V���U���x�K �����gA2�H���A"�v��c���n�F{+��Ǌ`��DYص�G2�-[p5��X
�c��X:��V"�qz���Gf����}qq��A��]K�xw�u�cBR�fTKm�ɠC5���!�F�\,����w���Wa{Y���s������M�s�,{pV�F5�Ɓ\둙�ɜ���-��E�4f�k�����C���xf�a�ح㨔fv,�15hQѫT��m��Hn8�,v[s�O�lq�C��gt��g��wh.pn��R�e�nֲ�Z�c�j:��ӱ[(E�iI�v	�7j[v#�`��Cn6]�]����`��,��g�k.�"ڛ.��86���k���NZ��=��q\;p�x���5��C���(.ҷ�VD�#��-�X�����xyfi�f.��g6�1�܏��Y��2��sʥ����:&8Q���Wp�������Ws�N��ƌ�5��0t�DK@6LK����#�����PV1ۘ�Qw=�8����91�`��6�$G�q,�56rYz��ǐ�q�Ge5����x�eYY�ݸ��Nc��n�9�+�P[n��ѭ�����D�jq�SV�3�9`���^�K,��l�e�[:[#�?�v��Mq�l�5��2ն.%ᵂ%�1�v��J���5�CL�1̺:�6v��4�qݳ��Wh���ܧ<vjE����q�]�A5v�n����:镶6&����E�� l5��,�N�N�x�m��<�F�T*m�SxR��y��\�]b�6�qC)���˨V.��.�<n��[���KTh�İ)�v��ү�߻�/�&=v�ʋkD��N�^��<U�3x:�p��cV�������Yn�z륞����E����ƞ�m����w�����|9_�-�EӇ#m��?x�7l�n��Oс����B�����fx���zW=e���୸��`��V��I�c�.���j|������9	8�����2tP�UOî��7���A)3�ǋy7)oH)3�N(�&n��L t�K�L$��on;qcGm7p*m��;�|E�8"[I��۲�16"����`�&pA&&Rj�眼�����l���Ӽ랲����`|n�M�Q^ �$�r1��5��Az}��_pD��jX��r��m���\�5Ժ ��`&l�K�v�Or��o?}1�=zc�$�q�s�wU?�S�v�x������#Yx�����g>I�e��@6�G��8 	���ZZ�7��'������L)�̳(�re�2Yws�EVV.�ܗ)7����~Y���hŠ�s��WA�1x�F1�)�*�U4�w�x� O� A� �x� �q�`n�~���g�Mwm�s���	X��9n�$�%V<�C�+J7<C�����a���BO�)3�!3L*��g5{ט�a�,ku�YpaE�`*Xw�>���I��Rp����8��U5��p�P�Z���,����)?���v�꧂�R�^v�p �\��]ۣ\L��o}�쳐A�g"�9�L��8)0�{k�k��t��;�dsu�h�m3��V0r��8$��S":
��{vܽf�MP`�rŘD��^��H��@X�7[6�v�\.m�Tf��WD0�^��=J	�g$��pRg�h8;�r��Ǳ
/�8A�n��=�\n_'X����`����.Eɜ~��f����^�:C����S��])T��n�ճ����sI�]�4ﵓ�B;��*C�Z�?�"��AI���̻Q5����E ���rP����K�sW�D>�$n�ҧ̧-*e3��Q�X⨪�362���׽S/Vm��wĨ\�n��l��o:��8��m^��%I����H��Z׳̸<ٶ������,g!c!'�y&��=����46��@=,�p|�?�֎Ŝܟ���:��,oE0�3���f�=;'�^��D+���!&pE&B]d��v<s�	�ʋ���<�U�s[� �ճ���X-9���ߙ�Mw�?v"�Qc��Q�Is0��jݮ�Vv.���삁�A͘�X�x���cX?�+9E:Nov�l��\Eى���8���յO;Xl�����ȇ�);�	I�^n����s�q5��f�s�Se�����u��Ӱq8pBM����m2�N�L���LI���_��K��F�dk��w\��'B�J�^vkw�&���W7�i��8>I�޺j� ��A�p����'�&��e�dݘ��m��5�/�^>��f����0x;;�.#���`g^���۝���W�^�>P<ӣ���iY���5gzd�d�w'�ޚ�Q�Y����Wv���`�3TT�N|�k�e�w��
L�NL�?Mnu3�o�\��m�gP�C��_�U��|3�i0����8!&�4n��:�Glo�?ʼǺ��T�uO\�8]�V�G�)Ŏ�چ&ٸlk�c�p��y�O��U����J�I@����*�:�����g��w�:�xq��Ӄ}c,����v�oMc�����F^����X>�u���n�2n�Nw������E��	<�P�����g?��U���m�	�g��nM> ��_+13u>���獤&�]�^�e7��j��'R`� �8!'q�ɱ�^�=�L;���ǉ6���y�Ҳ��O��J�n��Ǎ�~�j�i����g��pBL��
LRp��kd�l�0�у�4��^ݲ�綘6�Nw����8\�/9	;�D��y��}���ube��M�Em)hyY;������j���%�KBJ���������~}ؼ
�MU��Ȉw��R�H���ء�3B�o��ҧvߞ�����73��.�K��W���0�6��Kگf��rT�3sx��:�J����`�Rv�v�[c��z���&m���e�%�cE�9���N�r�GgC�k���=m��Q�au"]�hKo(�Ṋnp���/nKv�W3��O]����֐Y���`��[3q��d���X�n����h\g��[5���]R�]/���S�n�֌�չ֌Ұ��a���}ϒ�����	Q��������I�v��V�b�D�4��1�R����߂	1��#�9I�$�&�N!ӻ=9#E�G9��Nv�<L�T�Ja��0kw�x�pA	8rw�(�����P��-�����ͤ>J�[�<�L���n��pA����}���3�N�<�Ǭdb/5��u��mkbֲt��LͲ�'1ޒ��M0R17�[�հr��o��T��av��4�5�Dc��Z�A&qU�r����/��p ��z}Cx��,XME�3�������L
o�Tb�"������K�ք��5&̡����[��H ��n�Ř3����!���C�hww�H#�(WL�2�A�Ơ뇛3�ez�fՀl}���,���5��&�
Nf_[e�o5���s�[��7˶�G�����9��x��p��\6��bmk`-q�Ft^���1��Y��G]�uk����q������*�6�0�����+��):����6�Ŵ-�	���)T�83q6���xx
��>[?� ���W�qX��g�/�#��`V�r�9=�[�/�]#'�Ѯ�d��׮3F��H���f5��o&Dc"�U�4/UŚnu5sh�8������&�?�s"�� ��E?�4�1#po���8v���l���r��.{y��E�����p���o[�~e��q�L��7N;����YRe1B�����f�Cf������0=N�9��AZ��(��N'9Oޞդ~k�0)����I�����V�o<���^�Qɦ٦!�˵��v���{}u%�������y�:##��zy���3w[��q��Ntة�e����$�E;y&Fb]����<h��O��Ák:�.���Ћ
';ս�8_�^8rۛ�w��MD9�gی���$���ޫ��p�M9*%�V�ѠJ˕YW}�m��(�"��C��5���ƴ��K���7T�ǻ�fy�Ǽt�l��f�%��-�������찳Q�߲[��s�� �`-p�\�p�"���&ƛ��h�"������L�d���w)n��R|��n �j�� W�Li��<!�'�EX�>+����"� ݸr�)�q�&]���N_Vn��o&t"����c��A�p����	��%�F]Rmש����g������i6��9v�;b��F�5`{qՁr.��6���^���/���K��� ��V�Ukl�L1�S��pa{�(B}%:��`6�Ã��
N|�&��!�N�9��JFc�?��:rj�7�TBRi>gf��l��ȇ ������z⯨p�Z���,C��`��9�>����x�Z�=��D���SQ��:���g{o�p���)���D?�L�"���<�DLM�6�@����������zv{&������@F-��_|���x�`�t�s��*w8�Q�vh����P�^{���R�j��k�C9	ᚻ/�j[=��3�=�*Sa��m��Q�܍�T������MZ�f#�y3�\��Vl�5��!%��@�-�����8��Ξ�zT��3�[� �g��:ȇ)3�	IݺY���'�����Tk%k���}�փ�est76�E	]B�6�UE��q=�8�w6�:�w��z;�ۂ��R.��-�VB�k.e�vE�w&u����9<�,�f��(���:�?�L�����Ra>=���RF��r��*�x�W�Ɇ�5:,�y�7l�@�Q��.ڛ��o1I���Ⱥp��e�>IÀBM�L�Q��(��llU=�����U;���nV7�Z��ϡ��#�,������U,��E ����{"붹�d3B��m�pN.F�K=��}{a��4���dC���%&s^,9Rhq�56OUa��g�;-����	�&���1�@9l����E8	8�&��fy~_���݃9���9�/g�����>�pO�i�㯧�ɛ��@=З/�������)�픖&���X����������y/훵�Sq��l3�:���0��0 6o�}Y���7�@6���Ck��g��.���#ۧ��/=$�>'8���n�'[��E��D�2=r��˽#���8��C��'��h�sѱ��.4uWܲu:7ju�ٻ���!D�z��T}r'ۻM�<�J6kmt�M2ؑ��(�t$K�&YB���0ʾoG\ŵ��W 5�Kz_�O���UO�^�I�-��ѕ�X�]����L
�԰�f�h�̡eO���L�.�*A��$�?�o>��fd��M	S�����FiޜW��� ��η�V8
�||�X2���i�q��*�wb����`����]�}=��C4Ug{m��A1Â;Y}��u�;��[K�c���8�*��>��{�~��m��T�S����`����L��=����%�X9�5�����:�<A\�R�?�I��99o�]Н�Q�y٭�x�F98NV��Pr�`�g���0L�r�$��RǷa���V�
�V�s��wY�U�=�Á�`�^8	K��'򫗣i��r���n�1b��K�1�i���w ���$����!���R��1��c�m���� ���9�9`�Tj�^7݊b�=�&6���+p��`'��;�
L�P/��	���MW�T���i>凸)iWΖg� R����S����mC�ږ5�z�׺��`�Ӷ7�i�w��2m�3���y��'����)7�C��������;�o��}R�T+��n ��r�9I�&�Fv����vȍg>���AIÂ� ��%�^(9�Um�n�\�<Mf�m�vÈ"����y�dC��8!�ܦd��et'P�A��Ek��L�S��c�o�Ŋ��g80>+8wY5λJ�=��FK����	;��Q���J��!��p֩���q�wu�<m�#rjn�s[�c?�:�C���x ���W��P�WY��ZX�D3ـ�0Ę���	��k)�ڒ����0iWMy���L�W\!m�k��;��r���QGΓ��M���������}���O��xαs�L,x�?�L�r�9���j�ͦ���buϩ1������ŭǮ�	`6*k��/�-0�ۇ�gCn(�E��p-HpN�."ֲ�&X�5����yyyyyzzp{}�>>�����倱���3wI2���6�fn�C�9�vÞ�H�xr3���NH��5f����R�������lQkY��NB�$'A�Ir�����n\�0D��9g�ax�Ї9mT��[���G��9y.<M��z<�w��y3��g���C7l��t�G�����Rg��;�Xk�Lܹ3}���=���;�.p\u�g��	��/��=ʎ�nú��3�g��8�q7���o ��^g_���m8=,�G�{���0v-Pަ�{6r��zd�C��5�[0YO���^�|���HRN�:zKsǻ�gN+�v���}<��u0�g�ΰ�Lѡtw����(�<���gmU6Pz'{c�/��������k��޺_�fkVrTǚ�y��}y�.�\@#4z�;���� �%��ދx`�#ɂab�~��u3���%2h�F6Xq��U6��ښղC'�h����c8�Bvxy����N�j�P����`���z�����fd�~7zp�O�ߟ^S���E$d�9��� �9t���Ec��_5oe���t[{�웧<�S�i�7%j6bL�H--A�~�׽���=�>��'6� ��o��J�-�r����� Ӻ��W\E�N��3{����Q�����V����?=U���U2s�{����p�����4����;^�xn"��+�d�o�m����[�{R�C�s���˳o*'"�@���Y��qR�-Z�.^E]nOu�q�������ѝ�Zν�:C9�E7�A�ErL���ǱwR���Jw��m{�gG���4�ӓ�8��S�u�(���cce�ăm�;A�E�}�ܔ��\pVw��eY{���w_�o>�d]�츤{gP�kN+��}���ù�ut�vwgt9�o{ٯ�����/k�����Yw����3���̮ӊ�<N�㒂9#�#������G�z�kΎ�+����^TY��w��ҧ�Y���m�w�����+ ��Ύ;.�-�z��;��+�u|��r�ʂ�{ۊ�2��:���jK-�w�wZve���89��"�O��+H�;�&�W�y'vTeo��]�y�vVt\fD��YqY�OX\N"��=�{1E�������5bi+��o� �z�}m>I��	5��6�%�:Ů*���es����̐@I��%�=�2�]��yoy����:��:y�?h�2�?�G�4�|Rg����[OV�u��X0�3�l��|����b��Y�`N[ �k�(��$�3���z���Ǳ�Ib8Mb ���q�v�{�5sՠf��5-fȥ�9����z���e�����|��\�(��=a�W�����1�b�oq�����	I�ü�͑�����C��9�ӂ�/���>J����b�w��޽�������^0w[<�4h����[��5�ĳ�@���)�O��N��X����X���K`k��p`A�`-p�Q󀓇$�2�2���,h���6�ǊdC��Q�]�'�.�%yۭ���y[߿����bw�VI���n��'?A�v�zw����Wd�\S���}���sU0�b�/1�`�"*n�Cc�7]E����ڹ��9�g���;���{1�-3S<�G�w팱7��:pV�`�ְd��Ȣ�h��"c,X��e1߻�F)OS4�ל���׌$���S".�L���5��xM��)<����a�j�.����9Bx�랢84���et����6��c���r(��?�>)3�X�V����Y�a��d�v�z;o�'��3�	8���>��H��h��q��5�wsKt͇J�[����8�C����Qr�lϛY+U�Z���8`AX�:N�\Rp̚r���p�-�Jݍ�+�ѕI��.�g�&�"������!�)3������;-6����?�[?�%&K����z�&��W8}i��+1����*6���F Y��|Y[�]�pA�g��9	&��ΊR�W�-�<*��7���a��������qRg�BM�e�q�9�q��v�#ϖ��yye2s�gn����t��J����vtW$��^�"�_�A�sV.(!m��Fa38)��Q�bhh6����<	�5(QU���6�c<X�\Y�e��lc��^�9�^̎����95�wsS�iǞ�s&^��ոsR�ـ���	fm���䁥B�
ShT��2�`;�u�:,�K��0ͦ�ȯ���8I��'<ĳ,����e�b�L���f�[+@�j�կ;2�[nwC��ѭ˨����n0nlQ������k���&�W�P�C��!�rVl �yo����[�c���GjXM��sY]�XF]�����E#��t���C�޾�'���l�p�`���2����պ������I�e��^/H��ڜ8$�w�&Rg� ���E�֦۩���^��b��o=npi�E��0>9m�8n���!���ED�5�����NO�<[Ɗ/�R�%*<��m��A���n����ۉ�ٰ�v�q�r0�
L��Rg!�u,��]���l(�+\9ӥ�!'.m��f�ȫuSK���4p��j�O������Ȓ�9��2!�L�cF7ZX&���{a[�w=_pi녜#�[ �FH!'�3gsGV@!�TY��.�ɀ���h5]tlG,*M���#�J���:��CЎ����{����`��Â.�?����=�v{8�?NYYٍ��q�K,��Xi�>ۋ�c��1kX���]kH�Zי�́6�vnl؀�"��E�JĬ��V�9o<�I�#��ӑ)g�^�|��Q��^�޽��a�&���5R�*UB8վ�o�����6w�D�3�M���っ�pAZ��m������{1�'�$��\�km��lo��V3�JL���$��)5�6	���:c��j����֋9�7�q���ݼ\����,p�"����%��'GgQʎG�:X9
���ȇ�����9�p2���oq�oJ�3�K�j�$Ƴ�m��DH)5x� ���Q�~���Se�f~qu��7�3�u5�Fc��A�p�]�ȎOW����̕AA`���~���mm��v�[�6��q��p�=�Ge�sb[�w���,�~e��ݏ_^��
L�R�c{��u����aqQ�.�dwL8	�Vޔ�8!&BL�uVT#cf+Y������M��Ok����Mӌo1vcq��9�0pRia��tr{��B8��s �IÔQr
N �ΜީOۏ��*�%��Y.�bڔ,i�L��'ި]E`������d�-���Z`���h�Kն�l�h!�������H�t&͹���UN���>�a ����!�Rg-�J�K�0��l5�� ޳�AI�R�#{��u���w�s?��o����8i�e�!c��	;�� 9')����h����55���DS���[�����n!�)7��/v��[����/�Ҋ�U���<g��a�K�49�&.W�͈v�ƺm�U����w������0pA�ȣ JN:��2w�b�Q���F_8z����:p|7�?��?�dC��� ��y�۳��"��o?��q)pW��W���=pÝ���0z`�n6_fop��k���tH9�z�9&�����L��e�k�3�Z�c&*�cʳ��1��o1vcp ��r����A�I�N��J�ۅ0@�%8���)8qVd�p��W��F_8 �6�hz�e��A�����4�Wwo6�W���lh�TQ��4k�
��'�W��f�]U�0�7�O��,�T	0��TD��]�A���~����&*b�[�u�g���=>&r���l����nٍQ���5�oo�/�1������A�ۇ�I��a^�Ԅ��-d*x�.4�wa��Ձ��չ�g�=wbk�[���C�#��<�߭����o�p����|���NK���O>1̺����ܺ��û�Z�4�ϡ�X��v�%&ѓLX
�C�����7nE�;�;�}FU�����Á�`�-`���	�ݫ������b�Ζ ��pA�9��MS*�L7��Fj��M��Q�L=5p�n���mÔQr'I����g7z��ѳ�q^���>��D�:�箘��9�]z�*n ��ֶm�oT��@�g��g!��3&�IÐ�s�����l_x�Ç�bWv��W1�F_ ��6�AZ��	;��� +���A��Y�ޏM~9eѨ�5o���QӬ߯��~Ç����}����� �)���5"xg'Z��Ǌ��������ہ�.e*o�-퐴�z��`����3�/u�>y���:Yq���r�r���^c��'nne�0���툽��W/fیtS��:�6�.�in @�a�d���J��skak�f����l�ݳ�9tg�<�g�r�㔮�zF����ف�]��������AՓZ�,���g���i;q�Be��Ik�-�Ҳ5��*�on��W	�g����{V��U�=v-h�Tt󵮔~���%g�����f)��v��c%�ۚw5N��q�3�TlZ�˘��[������@GHpn��>)4�ml�f��Y4�գNy�:8;���b.� �8s���:��8\�O�=�ѳ��F�"]�S"&1��StD�c�]�����pF!�I���"�"K�O�`��1� �`�!&��eİ�aqg�����
�z=����K+���#/�V��yk����o8)3��UN�ٲ��B��|Rg���W{���5�5p���x��\I��t�`��滛h"񃐓���?�p�$NECu������{i���OlK�K6,��n�����y�&�K������#��~ޘ
("���!g�.�b�<w=.����m�(�v�T�qX:�_��}�	�`�\9I��@IÀ�$�gu��{y��#/=����=�����6��X��BO�$�I��S9 MF_[Pn��$��h3/��k�"���/{O'����/=�ނxg{H+_.c�=7�[.�ȵ�yU�7Y�2e>*{��"�Pz��_k���9�����Ă'��=l���Җ˽��y��MZ7[�@�`�����L&!=P��fH����m�pNk�07n�zE��cr��>wD����\�Ȗ�3���1�J�pA�9I�AI�Dq,K_�j<`��C^k�[
�����a����d�gu�ʛ��1�F_8 ���6��Z���SY3�v� ݳ�E����3��:��9�=��'�yݯsz���i�`|o���d�p���-��V���ص>fwx^��#��;l�^{�ca�80T�]�4SX�5�����|:_��I��2!�LWE�~G��(�����Q�,g͋��Ca
�r�L��;�I��54Cn��L�����޽���Q��/�E�rZ�%�5�cs����Wސo9���;l��)3��Ri���mM���St��W{o�����d=���Yg_	�wE�.b+�����'���R�c�y��&M�v cX�^`bFo� �|�wk��w�v9F�۬+�[� n8m ���BS�;,E��bu���X��R`�&+"�Kw#�cevcqƩ�C`�͵>�fߘ�;�3:�L���:�LƵ���y~�(g�8YR{;���ܨ��##?�+\8$�pa��u�	�;@D/���.Ψ� �h�M(u�����L@�&&��K�H��}����e�_�����Yx��Ը�vi�8��(��w��ޫb���r�؝E�iv�����Rp��(L��۝���b�P"%�� �`�&)��Kmp�1W]���	�`�y���S�\�$�|aF,A�g>�p��`�"ӈe�`���9���:�W�T<4��Iv�H�����2x8$bg-p��&�v�G\c�R�k]��n���0pk���<�.,ك��C����a���3+��`�eIY���Ub��a�{��n�k���o���a��<�<o�&�f�Y.���p�k�5��e���C(���H�y/T�(�RL��>�Ӂ���÷�%		3��8��~no�'+����o�����2K�pܩ{���`&[��0��A)65�V��Y�Q1�h6U̢�)�	��K��T7�d��vn���,q�Z��x;n���#�d��2i8S/wVu��k���O>EC֞���&3F�z9����kz[��&pG5F2艚n�n���oD���{�
l�=��
�f���s9m�i��B�l!�T�pH�g�8;�vޏ�22�?m�N����]C�vcw� �3�A�`�)3��)�3��m��~h||n�ؔ$����x��Ȥ�!'
���cu�L���o��w��g�;�R�����o9����v�}v�&�~wDe{!�Ȥ��wxχ^��Ӓ-y�1o���kbk'��������������fx}.�볞;޼�-���1�pL;129G�3�F[q����
�gg�0��v<:�G^�q�E�����:��S6�R{/�q��s�yL�0��s��5��|���kW��$�w.��w�3<jg�;���&�<�µN+���ۻ�=�����O
;w�`��ˌ�ý��
b��(�j��(�f�#�O���/1 �p��JGs7��q�%�ž]r���3�/N%N������|Gч�$�!`˂��a9�0TB��Ny�!rX���r�}�??�����z�t�|UM�~����}��_v�z��j��G�����z��6�[+Z�!�}5��囊��y�i�V[>b�iݧ���G;|��ɽ�wo��\1��{z�{9zC͝}C�E�t�2��n�����J�Ndf��f���ɽ$��o����=�;��+��t��qc���Í�[����{�����w/�ִ�0����^��r�|M��w������o�'/wi�r�oy�h����>	΋p�;�[���o�ĄrJ���"B��<�����Pqw��]�gb�^O=�v��Wj���z�hޝ��F�[,��(�z��徴�M���?-�f���#�ݞ��1�~��o��ާ��+=�uXw�}U�BGع�N�og�����e���'��I��]����:z�k�3�,�g��vO!�U�~{Z]�C���-���=��x\@�f���w�[���vyqbn�(���Q����Ռ@�NL�D���\���<�¸/G��w�=XøW�{n�I|i\A��vd8�w e�!՞����&!>��;�n��V�����"�me�����e����B���sl���+*�ח̾y^TT\twq�\Q������{�wq�,�ݝ6��:.���z�����DtwQwλ�k
.��sj�u�z_J�ׯ��y�i*˻(�:�筮JϝgE���y^W{���|�֫�TWfe�Y��������:�Ϲ^w����y�y�g�YM��wg@�E�I٥oj��EE�|Ҷ�[�k�������ʼ���]�{n�㢳Jҿ+�,0���$M:�Ȩ�>�$q�Y}�V`ͮk�خ�o�z 9��َ��'l�$H�0Ene bE��i�ehv��l��f��CZ��n�ўd�'7d�O���+�Dso
��/Z5�)`*�l�eD�!a�=�⒝��5m� 붶��Oa`Y��:�7W(��N�'�ݻ�gf�/n7�<���،�'�!��,��YY��X�aS�t����X��=4۶��sh�n1�Љh��ˌ���t�q��N����q�W2��Y}<f�X�\1�(�%��j��� 4#�vSع趟;�	� ���8Mc�а�Ԍ٬ƌՙ�&-t:^���	�����L4�.KM.�V��s؛ԭ�(3mx�<���\E�+f�%��Φ��,od35rh�#`�f����[GjF�]��mCM,t����]���n�����[�� �f�)���Ŗ�#ͥLcr���zw���c�n�-��%+V�SCL���\ES1�n&4Mh���#���\�u�º�<�{�:�֧�`��l�`�vϭ�sҵ���Q`��n&��γ�ʴ=��%�##�e�r�>ޕ���Jn�5=;���٬�q,a(�]3��ZX�a����eu�+1T�����B��Nc��m���A���շGi���m�"�}���=��O�#jU(���;ef�%:�J�	f��]lH]�ֻl��F5Ѯn��;Vp��,f�Dc]I�n��EhX�|�.�g\'d����	��jc�,͐iJ�A�cb� �`荍�kq�\�L��W�=L�x�L�I�W&Ś���s��٣72�ˮ�0�aE�2i�:k!��� d�Ƀ�+��
�1�vܞ����H�՗���ɛ�Ɗ;k������b3'U&c+�g!�ՂF�Eiv�[�n���po;RL<N.^���Qol$�z��j��ܩ��@؏噻�O<�e���.5�*��t�����k%��.��UY��X��N�v�l��~��>}�����jN�x�ڽ]uv�u`�a&���K�R̓\<DS:���K/et�jba���F[ڭp6��bq/Qu��WOk�g�Q�%�
6����pZ���!���A��r3U�n��ŰX��E������٬h�BM�/��ܗf�K����ٷn��0U0K �ef�-��7vb�`�,�<U��u]�Tv�V������~CCc*6�k�k�m�v%���v��&Q��!�����׿)G���u���s���`<U4嶆�å4�����6�u4s�p~����L]��ͮ��bƱ��k����GT��9ǯ�[s��'9�~��71��J�y����W?�0pAZ��K��P��7�}"y���3�v���?���A)2ݚ��-���5��k��Ǚ��n�x����a%&A	8����sۃw!�xF[���Γ��U4ݱ��mКsvc{��9�=����^�}��o9�g�0V��n�?�7o�L�	��U��q���\�Z6�����{+��j�n���������C����Q�Re��m�U���fL�.�SRa���X���퐋��G_o����췜O�&��&q3�E�sOpǉ��f�x���W6C�M�0�A�X��;�i8p�..�8 ݲ���ЬλmG�#�o�d�S��g��{I���3��'��{@�r�^�号�w�SI���ߠ��N����C.k���	O���?���Y85st&��]��Ai����&zW�x��7�_��r3�A�`�!&�L��l�&Hy"�6�������UFV�+����	$V����'� ����Mr���A�'�ށV�|�?���3�swx��+�/[�A��2>
V:����5���ט&`��8 ��9	><높�dFU����p"y�l������`"[�v?���>&�}`t�dfͫ"��y����v~��r�i�独q��ʙԲ���jt&���9����CkaŰo�AV����]S��Z����2��lT����ȗW��� ���o8	?��M�)3��U��n�9�=M�=�������[x�D��\7�A[�����Z%e�1�b._����� �$�G�&��t��?��l�����Y>�dT?E��%�� �Ηa׺V�p��=%�O��ӑ�Il��5b�������Z8	6����*��}���1� ��q��$�A)7�i����x����,,�l��?�p�V���;Kө馌��� ���0r3w*���g?�뀓O��g ���I�+,�2kE�.Q�g�������(W��1k`m�����)8�uK�Pn��iy��fBLy���`b1�f� �GMq-H:���f�\P��b�p�׌�h}�؟@7,}��%!�|T�A���{���1��4Ʋ�t�f�AX�pv��
L�!&r�L�z8dl��j�s�8 �8+X�oy�&#���+��������+\?�I�o_U
�+��.��S8 ��g ��{k��	�m��-�5��R�1Z���9�Z/[�
�A�[�)0r`�l�\]ϜU��b:q�,f���w�	?�
�7vy/|#0Of7M3� ��kD���{iޕ�V�������sTi��g���/���Nɞ���w��]Ƶ��z^ǜ����N�;��]�t�E�u�t��߆ �ox�>o8pj�
�82kY3j�.h�jR"�vi֍�Ӈ���s�ff:�"��|��e�"�Â�Dx�ȅ�7�C���wB�큳�3��xc�ыS���qA8��x���-�%� ��tſ_G�e����r�9�&}���;OdANhO��!`و�k��P�|A�p���I��BO��?�I��#5[昮���R�q����v�u�q���wq�A�g �8	1z��|����š�X�A� ���L�'�q�����ɝ��3�M��F�8&m��Z��BN�&���3Й��C�Y��0���CL4x���8�����;Oc�NhO�� �`���G���C�άJ������'BN�
L����%�9n=��C��g�H�vp\�������wq���4��vG��휂�{�P7b5���Ï�S�gw��'��;g��j�Z��Y>�w՞����n�=g���7ӽ�p_k8���7	�����81�0�Vx�#�ni��1��|���ٳz��=��n%7m�>%<W�Y��^�Y��ّ��p���5�:0p��1�Ѷ����*��k<]�Eu�3��T=��w�~`�w���ϋ;kֺT���݊�,�v��EV�ǋ��mv:čc��QM���Ԩ<#ͺc�e�ƣQ�6�T)�aV�m@��n
��f���6��L�@�4u�6�6�翳���Ѝ�c@1v��@Ж�aQB�$�#���]�P�ƛ�ﯭ��;L�'
L�$��ʻ���=t��$j�<goOg8�0{V<0�X�.��)?�����u4�MHه����s��9��gwg��c��4'��p �����2�9I���*a��f�g�G�8�g� z�9$��I���������S��	��(a�z��{�=O=c,O�2嵬9��d4ൌ�s���ݳ�3�_8pw9�8we�W:5��Ӷtǘj��e�&[t������'k������5��&|Rg�0o[Y��-�NҊ�u���,�n���7G>���pV���/;ɖի,������?g�B�t���DM'��He�3{ܶ�́�u�Y�v���%r�A�^�.������3�_�8&M �p�$���2dC�h+��Pâ�=��n��V�����:e�����%&q�,�0 �&w��������6]��~'����S�$׼��$Þo�2c�m�6vMh���ȩz���z�@�ӈ�}�W�O�Xlx^fܼc�o�G�p�pA����r�{�^_�r_:H��~,�/�A�����7���Sko���q^cL��u�S#�@>I���3�+����"���1٨N�;��A�[��E�	0ra��8�"r��fA� ��B��D=Zv٨��xg�[� ��pC�3���]5�K9L�!&&�av޻aKW'�z�pv�A�����(��Śy\���೼�����}X��I��z�u4c2}Wl3_ߩ�ľ��9��+���9�mӷ'��3Y��"�V�1Tu�}���K,�}?{9���> ��&�m��D_f�c�9z�����LwE���˵���p�5��BN���&FFI��v���m��V�ȉ��ۭ����7�Rc1a��.
g���G��:�'��p�� ���	0��<�fa�|�w�������5�����z����M���^���ך����@�lAvsż����l��|2�\�=����0�"rMak��Q�~�[��9I>�l��BN�' �H"rΡ�nٜ:�:�JL�wx��������nG�5��|8Q�#x����8���y�$kYrE�`2kY;c]�z��b����c+[uʻE����s�������h ��m�l̇z�j����%&وU؎�]���RlO����`�/�Z;0�0�F��3��=��7l���t�:�s��9=:npp��Ƣ�Mv��7�X:b��,u�r��\����Z�2������ci����n7��8 �L�q�[�Zl�h�/BtY�	T�����c��`�F�aQc@\����<g�$�%/�"� *�%��@���ɫ�[]��A���1��)3��I��Qs�U�nÑ�5��A�p�6Q�`{񁯆kc`n��9=$e��Q�� ����T�MJ-EC��1%��Xk�D��ȷ�V�a❦�Ffm��¤�[����(ƿY��������7PE	�(?K�Qˠu��l>��Tf'(5%?l�>"m�����pRo9I�S"��e��"��r[pљ��c�S=
�g87x��`� �8sf˂
N�/�8���4�>�@�X
{35���)It!6��K�X�	�ZI�k���}{��A�ۇ!'���Bն�3&��%�v�{��O��/y��G!ٗ4	I�N���8#l;u;TKB�8p��8qy�krqƆ�JOQ|���e�"�Ð�@��;o��m!��9���L���wż�`e�Y�c�sB����1񩞅h�������nQe(�!C��$,KO�\8n���2!����n�L��s6=��T���c�Ί;%+�"Z�Am��"�C�&C	 ��>��f��n�z�،�����6OQ|l� �8�y�d@8�����ncvs��vKl�O���q��I��(ޙ�T9��LŽ�{D:;�{��O�������SM:y ����k_��P/;�w�sp�qs%���%��'��	5�jYH�	T�suip@�:�km�:Gn�[�|���Ŭ����[��h��F޻������ښЀ�6����9��Q��e|1�2���qˎ8�%N�V]�+��m�\�گ/UQd8��tT����ƷJE`�E�E�D���.�Z��mt�O(��M�l�#)�#@�V��N�H��/j�o~��>�X��l�u�cmg@z�6,\t�q�;a�u��uvn-�������w���:��6�/:_s�a��5��s�$�J�M�7���0��Ӈ��BN�E ��ͳ��l�9��H~T-��U;��_n��|Rg �aI�櫠�2r��܏0 �`��9E�V��h�헴���r���)C������6\k8$�&G�4��6�8���M=P�zڈ#Z�s|�A)3��}ۼ��p����d���m�1=I2�����*�9	0L�4k�E�Ͷ�DT6gdd\�h!�Sb�^hJ5S?>5��p ���#[HpRg�3�������d���,��2���3��b������s����U�6F��ŗp������o]�rۇ|�I��7ҋ���FOQ|����f��J>��p ����ȇ����p�����=u��L��r�{�\'΁��S�W��l�������{ӧ/Fw�|3��&��$��!�z�O?Le��!�s�r��%0p�}�G�C{�e���3�W��n����U�Y��L�v��(��Y��k�_�g�^pg��j͐�kHֲ嵍G��n��I��\V���UC�E�n7x����>��Ɠ?�%&�*|���Q:��CNk�A�<\�����jQyC\�=(��#/��G��{H�[�y�hJ�7]�Bk!�L�>I�/0fdC��M�tU��y�A�g��1}��.�P���s㉃���v����$�9��헬�ݸ�|��[%}������-�8��>�N֐:��t�1��۳���� Mkt�����>��W�z�k�$�ǈ��d�W��b�T�����nM�_+SEūhj!��g>I��"|R`�#Z�"�f6,�E�Վ34R���ڝgA}���V�%c%����9��6��1M�8 ��aֱ��b^��<<<<<;t�}>���|߭���D�w�ӕլc뽻ޕ!}���dȱ�^����L"xѷ��;Wę�D���'a����iY�j���t�8�N��uJ{�w��qL�~�R|-wNI1_k��Y鞓6��vP��<R��l&���QJWƉ���㇛�oϵi��o�̻��v�!nuٝww�｝P|��x{:�'\��
�8�`�&�V`�wrv�.��{}}��GT�ӱz�v/��H�װ
����v���\��bg������<9���٪�g��2o8�z���5�{�����NǕo>@$���뽻|�y}����j�4�y�ao�ՋǹL!������f�C���{yg�ݹ����&�y(�E�M�vW�nh\}�����4��5���Y�#�!��]�ӾY��]��<����4��@���:�N�����n�5�4��v���y@|m�M��.��}ϔS��
y0�k:8�<]�VO�=��]��={7Q{�[���㙹��wxB��wXz�`}1��ss��9��ž��)�sՇ��s��x�"�;M�֭�{�hi����l��%���C��a��o�9�Be�5���4Ìm:�e䛬�޾���ۋ�ݺ�xF�y`�ɠ��R*uI�v'��Ǖ��5o�O��g�6��ޣ��ס�ao�>��*�n��=�{VL3���;T����Naa%n7ޝ/l�y����2v��7�"����#��\y��w��s���l�����I���9�����;���qQ�xz��l���f������oV��-�@� ��Ϋⷽ늏#�y�ˎ���Υ�dgDu��gtwzdw>�au���&ZtYe�y��:8mgw����۶�e�޷A�����Xm�������η�g���U�qZ_;;���/M-m[��s�쬾]��%�9�Y[�^�q�y��՛kmu�������d/{ݕ���$�*��#�{F��m�Fu�Ko/C���ΞZ�^u��mDۻij/��N'ppY�~�����8�lY���R]�i�G��.n���2:,�8�ˎ����痔v��G�����l��֎T\��k�׹;8���[n�{V\�����pb�V�L��CWz��8�8]�ro8I�����q�� �q�����Ƚw�&2Q��|�nU�r=�����2��TK�����_0���0	0�� �&pA	4���{���MF��<���9����b2��	
��BN� ���2N��0��l��6�茺.��c��j�l8��S��u�[�/GJ�G_'�����e�}����m��0�VvD��S���L�z�11<��o�����o?�p�8	3�;*�so0��6��x�7�F:�jٺ�V�7q��
�pA�C��KAZ�/}��tY�g�� �Ӳ�����ȣ$$�Y�VQ���7�7���/�|�����U�pBM�L�r�9O��m���Q�;���4�v�� ��>�܃����3O\/�r�9 ED�F��kU!���?/�"3~bypk,��xq��2�	�l)�;-e5����������}����'��c}���{{+e��9�},���#s$�US|  F}��?��.��탐n�8>	T�}��?!Y�:����+�U)�n��m��[y���r�y�LXeHYFY��f���Hv�v�p�É�9��؎�S���L�=��}r��BZ�r;�a��?��	�`��/\9I��@I�vp�Q;�/�r^�2�8���ӄ�[�/�	��1���o���z�m�0wɂ-���j��mvA����x��O\/�'-��.�?�L�A��1��abi�?�D��0�7�`���O��0ź��\��]��eR���;��&��w_�
L�l5�Il����w��b���5N�&�
N2��\)ݗ�ʨ�$e����Sn/�
�����S�<Rj������	6i�ڙ���M��T�nv<L�'��� ��-����L�plm�D���'F)A����S��{2��[4��Z�nE���*�'S6���0.�&�=��.��/�����������|��������-�������@�!���N�y�n���j�pt����A$ˋwc���늝��s�e�ϊ=���^�Q��C�i�ɹ}
��WB;���k��Mmr���0n�:\�c�I�]��)�v�'lWOf�����1Gņ�{�cfܜ�/J֖R�&�-�]�b �7i%%+%,�Ť5��L�e�%��s:�k�Nұ��q՞-��v�����s,w��I���͉�����
���V�\s�X�8�T�m�(�mbjtѳiOs�������e�pBN<�)?�Ѧe�>�ԫ�'�ۼC�3v҈c�[�U���?��u���v��g ��8"��3�W6ύX����!c�7B���ꈈʨ�$e��4��=�>p��.f�sea�ׇ���3<:<Gk{�̹����[Y�l;��9ݴuT�Gn�T3���
Uf�4��)�����v�AI������	���B��-}q�s����a���dC��7�uϳ4���9���ޚn ��D�̝ve�x]y����L�5j8mkX�X2��F�U���p���o���ꈈʧ�$e��M)8pI���ȆW����={���}��Ը���\�̎��n��YU�R06�(l��bRS�3e���[������l�X�^�AI����U�{4<­w�CJ��;�wU0@��x�$$¼D'�Q��fR1Y��8�)*
J�Έx�Pu�������決�n�k��M_S\�	&Fw��F�E�����BY�:���^Yp U�ˢ�5O ��q��iu�uϳ%*����٦���4*އI˰���O�J�^���5w3�J14��]�2��gDӈ���^p
N��^�pΡ?�'G)�mׅ�`nm�Suڹ���e[�����g+p�ʋ��V2LO��F���J&�K8�v��\�0mT��71�4��;q�R�:���_�����͆I�_�"�)��+����o
d M�8̮���p��	�g$�����$��2�چ]�{0�4��s��}�#����L;@d���5U�eȆ�M���"�e�2��sʺ���y[��2^�'R|����	�t���7�L=:�TC�4����x9d>�zH�Ox��y��E�~�ޠ�y�^��㋚���<�7{M�;<|�1�H�y�s^or��A��Ms�:M��JQ��64�9S�K{V��M�}���ra�ri��{�+z�D]��"��po$�$�$�O���0ڭ{y&���2%�u�z���mY��H���k�$	��?&��	�1I��'�.+;Y��c��OD��oLu�5�������Z�V2M��F;,�[�*l����8�+�R u'I��J@I������7V�p-2͞���ܘj��|��D���Lv�;k�*��3�DNܸV��$���rt�fj���T&�19�0���Z�2I�	3�'��Q��+�7�3<���I8�vY�a����71:8y��5E�t�?;8Zݽ��16*�C��Ź���'~�ʝ���2�y�|E��D|�<�Gw��zO����C7�|/������I�Dm������i��۱��Q�;}�"q�&
��m�,�:�n��?�=�ta���At�1���%�ôWJ�H���n.n3Rk���&��6!mb6{�w��(|Wu��Y4��K^[��?�qJ^�=o�Cv������q쟱s��ũ��nw�i�;q�I�6��j�+�,:1��&��$���T�0�F�Gd�n�Ad����8D�)%�wp.�ݶ��s�ڥ���I���[��nǆ�]{��of�%�s6�ú㧜{��I�$� �c����mY���쾖j~��~��Sg�����y���!�u���\��D8�k'�Y�Y�{]�3е�[Dx��2ow�3w��!� D��?	�g�������Ϫ�O�>�t���Y��GNfsk�e`�t��7Z(i��Oh���i�Bxy�tu�����%n�0��u�PQl%v�BSc�=ٕa讍�ܥ�F���N �C��GF�ͮ9�T9���b4�g�n�W���<a����	eMٷ\
�)6֖(�l��K1H9�c����pAG=<Y����g�Siˎ.A���eB,ٷ=��p\�>���Q#Q�\GKf���:��Ǧ9�[/]!d�/7e�n�`������/�&[׍I8	0Y͵�����Z������~����6Vڏ$��a���ϙ���©�X���V#��ݏ����kyc$��u�;L˛$���}��O�`Y��l��n�z��|W���	8��s��M�gc��	2I���ڜ�s͒jhƁ1�Ғ��=ռpŋUV��|=;O�]���;���g�t7�x	0I�"�&%�����< C����6�[#z�	J���RS����f�{�l�w�O���2�:`ILV�Q+O^��]��Ha]�4?2q��x������㖟�ڱ�nq�}�Og���q���&v���5�LI�g�W'�;�+h�8:L��T��U��j�l��v�8`k��A���Θ���d4k��Y�ꖦ�$焚���i����Ѕ��9��NӊL�1;M�&[����9��zLA��wH<����V�YF�ڕJ����k���$ד�Q�1ꗕ�;����d����p�t;m�{=F��3:Z�KsEv���/�wl�I�m͹��f=f	�S�7YՕt�>�NӊLo$�BS�F�<���g�z�d;�fa]#�$��rq��z��c�'�Ax��q��, ��N^�V��9��6��x-5�ʈK:6������a���$�+���̡Q�o�N�lW<ji�;�!��=�SZ�� M7�:�]ss��I� n�n���]ۯ�,y��O��-?~�*�}�_��<�dÞ���������d�{�n���$��S 	rw���_YB��r_d�`nx5�#vD#*ى����qիyCgo�x�u�R`�y%޻�̩��L�o�_�^���[y,�ȶ���i���2Y�3[��Y,~�8o?��Ԙ���R>�1�R�΄k��Mr�r^mK�55���{�ڔ��^��}<N�}��~k(�:�wl˶�U�d�V6��d`�mۅ�2~H�p�e�0� ��������~��߈L���U�0�Sv�V�)N`��a�bn�<�{��ݶ����v���f�vt�raۗt�՘n��c����Z��`��	��������`���2�-j�OGZ���<FZ��jlZS{;R�;�]��w�2te�X�t[$3mxE��ԧֆoB����wmHu-�3��ʳ�62�6B]-7x���L�r�o�7����?�Oۤٵ����	��4$�H�ؚ�I�L��"�5�uˊzs��ܗ*�a���nZ��o�SkK*�)��7�W����>b��3q:�u�J�������f�v���07���L�1�7��ROvq�gK��'e<�
Fk�f�����y���?�z���y�k���yصu�)�L2�����z�o�)�@!r�n��Ǯ�Օ��C�Y0ʭוW��?�k{�ol+�m/	[RG�Z3�I"�ރ�U�>�nO�7�N��^7���l���i�!*��)���ൖ5$�$�$�����[�Z�w}�Ö8v��h�����Q�@�7	��z��o_�ٙ#1��d���8�E�f��8�m�|��u��[Rw�Ο?�&�Yr��[��9{{t��������;}7���Vv��9�V)v���*�����t�n�v�IyY̳ۍ���i͌�b�\~bC|zh�r���3�OaԬ��r�@2�A�]C�a6�Z���~\bY��}ݞ<">�a}7����D�����h7|�G����]C��(9<��p��cůi�|�oO,�lgϲ6�7x�Gw�����?����
�O`�Y[��C�Ƽ�z'���e{q.s��q!�eI]��w�c�FS^��l[��>�b��|��K�PU��Z��r31�hX�0��;�g	��M����K{�QP�zz՚yE=J�������駅ڛ/6nos�E���f��Š5wf�g'�t>8����R�U�}��z��v��֐��I�v���K�f���_����vO��}�r漴��L�l3WX�{=|�Q!��1z{����aؤ�������W4��m�� J6g����r�����-��[���M��c�ƶno�>}�N�����B9cWר�am����y�;{�S�]�u���k���'��=��|:#�D5�o����Xc�/_\��hZ�_Y��4�e�+��� t����|��+.�(��,��ٍ�>aā�4_�7���.��۷>N^�<ӌŏ:�Gl�q�\`?���A�3=�nV�%
��)æ��g�{u�t=���=�W�Y�۞С���������۾�}bn��\=��D�7���FGݥ0����,J�޻�u���<zͮ��d����x�</��_��d0���{oX�>�c�4�8��[���"�3�d���Tt��e���y'�%�)���Y����㣛Y���gح�g�R�N��3��У��켻7neh��.���b�+�tj+�4ۍ��L�鹸JK(�zۺ�𸭲�rv[�}}`q$�a�/�<���(ⰰ'���탁�I�Y�,�(������q$�)RO-�nm�]6q$Is����y��n[dp��'H^�9$[~�nr��Z6��"�,6՜�&��{��y�L�{X�$��v����'=���% Qy���C�Zۙ���{���i(Nrmͤ�ZH9�c"t������V�Gm�#cm�sm�ok��9ͭ���HN��s��_5k��'H�-,?��O�>Q�3n)�@�s��Q��tdⵑc� �X�4P�ݒkZى���Z.�9L��<Bs�"J2�XƁe:�L�j��H~w��M���-��b�;F�.*h���Z��t�h���7k� �����>���[s����WYSV�NeiB˘5 &aKqs�`f�Ю�rpOV`n�u4a&���i��ݤ����I˦�5��VM����CMB[��Ʉ�R9/[��c��j���㣑ʣ�{G�N��n�X�i�`���:x�f��Л.{S�.���q�z�E�ALXݨ�^�b����g�۴�p�B�0�'c���nWؖ´Y�aiP�x��W�6�e�	�	@K�+��H���6�@����|z��nc��`8�TBgQ#kV���$��L�k �(YkZ�&��5&�s�- �Xj���՛�,"K�<�kNwI��CTcY��ٍ�!t�R4�َ�&�J��)55���-��0��ܛs�4��8#9�����Nݩ��A�
u�tԎ��1�j\�v�Ҧɬ<W,�4r1��uC�A<`�t�>��|�]��gku��f�7(ż�۷+�thG�z�#QpXF�u(b�i�Y�4u��D��=���Ŵ���i@�J���'A�ݼiq͹�K6�v�������1�x;Gl=� ��ٳf��j6�2��0=nm�����9uZ2��aj�k.�SX�S�`�e�1h�h�ނ�9��d=r����x�b�8���z�Xө][��`ȴDpOt���R�ΐ(�5�A��!����b����#ؕ�u�4���u�	n8��w<�t]]�cH�tn�OQ��%��D���k��7Q�9*���%���)]jK,�!�Z3{m��:�n��V6ō�n��{#�m7V�n�3ֺ6�#���l�<X���Jg������5�ִ�8֬�b&%�:nXlcB�ɉn�:7se�
�#���n��祆��YX�K6�)2;iBˠ�T��R5fa��˨LcZ��a��A��Y�8foZM�;[��9I��M�l��s��ۉޝ�zO�u����rXح<�<ۅuׁ�ヮ�N��r�C���Zٹ�/+B�tksM6�tZ�{u�����F�M�U"t��_����X\�0�kp����O���Z̤uF̀sWEu�ng������~N� �v����ʔri�����WK�f�mz��bS�p��7������o���wh�U�4j^�Y�7m�W���]v[�3�}r�ok�:���y���'��v����y!�[eK�hr��PBa��t�k���:�:g\z���-�]�wM�N���������7�B�Ww[2�EѮ�gyk���(o�x���f0I��$�J݆�p�6�a�[XlVc&ۺ�eAL{/���{]&�2~-ջ�Yfv\������8�Z#v��z�pm.��0�3����l&-!�3Ӎ���I)�6�k`�Umu��)hy%�N�����RN`d=�B����}\�	*a���ȫP��|��F���2iƲt�3��X����v�.��d�F�/�#�̼
�u�/��	��0=7y��l뻸}ɗ�YG��r�X�^2H��.�5��ީ$�v�>I�7�OU���)"�5���k��ǔ���ݎ`�$Җ�w�$qj�� $�x[���p�zǅ��;�g_�uq��/��E7��n	�M��^��+��y���7qMeþAOJ��v���,of7��p4�������F< 5� P�`��k��f2t�r�R�uH�1�[\M��S����x�����I=N��'Vv!�AV^�r��	Ƕp��/q�m��8#��yl[:,�}�k9��ڗǅ��8D�I�WՍ�kT<C���5�����JBT=�.�;���!�z��~Ӫ�b��V�#8��yt�ѷ����w�?�A?����0Tbi�?�`h��v�����lęwW��"޲���w�0�o$��&	7�H�.��8��p����M�\i����Ȫ��J�8�ˁ{�V=�����]t`�JBL I�P6��c�K�(���X[)�j�x��&��$+���@�Ni��]�%gk$����u]��0�Sh���q	E#��K��3�xg$�g�0[��8�ote��~�Yo/�=�]��"ީ�uO���{��0�]�����,ٍ1j�U��^�n�lhYz�����9R�K;�:��_=�ݴ.�$�y+""�!���mǑ�6��oi�:��s���M��x$�y�Pyu�ֶ;�B|��o$�{-Y���u��������uWJd�߸�ʐX*O�*��3�ڤ�����I�U�@�Ot�K�4�^����cRM��^�T0��T%��[��o$�U$����U�H��y�82��<u��@�����������,�bl��o-�Z8�aX�i<`�����b��1��֞I5:�&p��Q�$v�-��w�~������(�M����擓�1����3�9Bj�uX.h۝k�	'���������.c���a�۹�̾���w��v���ᖒ��Z�V��m�A��w�����O�I����6.���o���]�c@������途��(O�}x��8*�с0³�6�-Շ������xF[�4V��Pƚ2���L<� �J����7�юga �*�t��x��w���X�$�8��r%��_m��ǥV�T��0��<�{���X*pD�
���ǹ�cW���i�ѳB��OT�[#��|�,r0d@cf�Q�
 ���X.,��z�D�e���q�2B�6���ӱ��n�֭��G�zsI<��.*ݨ��G"�9e��T3���4������*%Iݱ&��{a�ͼ�[-
�խƇ^@<)���b;y��7$�:�cr�{=��{%�c:zv��mn��\�b��ؼu=anP:���Y��*n:�a�6�<"�Vn�Ns��0�ظI�m��G7#A�v#J$����4�j]�s��,�T�Lޢb��-�ղІu��r;�hr]��?�>��K�Z�I�I8�Ʊצ�#���^�@�Y	��ږߦ9Ʀ$��$�-�:��٣�U>ˁ�ܸ���*s���z��y���-F���L�}��䓤�	C̻4흾�w��
xCī���Wp��
ĒI&�m��SG���7�z��S��ݼ�kze�:�q�Meꦼ�˴��K^�VVy��o]���I�I�4��O�M|�S�WAi��9�++����EہI(�IG�����V3%tѻ3,�eӮ��oalu���.�lk7��Mq�h�3�g���bw�ﬞ�%����D<*�=�Y�w`~Ƚ���2�),�I��n.���<��j�q�x܁vn ��Ќ=�\&{z�\��^��L�<�ʦ�ޔu��/.Y��W��c���o������"�Wq3����2j��&(�]�v�o_�����:�ƭ�~����&� �T���I�������V�I�Iґ��9>��� ���ײ�GT���zn�$�$�	0Srg�˕���q8�y�ܬ7<"�$�Ig���C�衫���zV�?�o���v��K�l�C/�ҳ�o�ߣ���	���S{o�$�����(�ֽ� ���{�E#J����Lg:%v�hh�Y8�c]u�f�Q՞�s8����hi}��,;$�A6--՘ry�tR���x�Ru��s�����`�t�$�فe�u��v|�����Xny�E�Q�g���x±�Iu@��W��<)��w�>d�%�go^o>U�Z=Ǯp���^���vay���재w�m� 	��gIŝ��!���矎.cM&!����[�֖��f6�2!�����k3�S{{�7�`�p�f�����ė������nD�c)�W���[���gt3�5�o$�$�M�	�u��Y��&��G'��Ue�fz�����$N玽��j�`��e�;��ah4��)��������ގX��cuv峗1 ���/���W����8���_���d	��,3��t�r�����I��&JE�m��A��Qh�q\�{p7)�ۑ�X�U�onw��ś�������zs�ʩCy$�2D6tQ���̛��Lbem�����i�I8I���./7�<yWp	7k ��zɝ�wn&�Y�4Ç�v��񡪥���
�k����Y15FP�������g�_<迤���;W���DK���ۄx�܁��L�����Y�cS3-������%Xb�1��}T�l-[�&��%/����sm���y��b�]n���zɅҮ����&	$��i�a�g���`�</��4K�l&�o-VJ6C��S:�n��eMi��uup�O��{�;�_W�L�ܬ7/��o �g���F{�0��f��^lv޻oy$z/�n�BW�;���/1��g�O�*�8U7��ϒ�M��L6=�ӻl.��'�	S���@�
QL^�Ż�EFB�Wy�U��I�oI@I�3͞n��5�����	6vU�i��7���Oo^3�=֙y�����f%$�o��zJ;wv�u�W n���[�n����#�����S�{Ra�7n<<��vz-Ğ2�{���{r��]w���#ZSRlpf�n��(lc�.��[?sۑ��W�R�Ѕ|��-e5��+ecޘj�T���6bb��˧��3����Uk���\Z�X�	(��t��.��%�J�N�����X5c��t��ѷ'I�Y�g��+�['G9�}+d��0��7]�gO����C��b�Ay`�]�y'��q�Ѭl�f��γ��;��SKфI
:�����;н:p5�E�De�sջ��a�6C87��Օ�ʗK�*�_~�{��#٢�6�]v�Uz.{5ױզ�;��C�xɺ= qx������	���v��zY��!?+��n�6�nc�íN���	'	$�6Ӽ,٭��m����f�tL��9l�����ޝ,��ŋ����DG�VÈL)7�Kww^�\6�_`�V,)�ء>���X���M0�����]��ECI���۠e��p���9Y��}1�ty^g{mmO�21��BZ�z��]���]ۤ�q�����y��R�I@_M�Ɯ9Y�[ �gp�kI)*��byÑ��Steӻ��Z�y�m�"@T��� ��L��00gd�=rq�I�:�k��m�c����ȿϮGܽ�^��7~��m�I�'�I�����\��0�I��ig�w���^c����9��/^�Ur^5rZ;���
0���n?t����gũ��N�Zt"�kνW8�[Üs7�GN5��{������$�N�\�
����t�.���f�Bqk��6Q�����;��ZeI��P�y�H�ZZ�ձ#ԙ[x$��#pf;e�~̱Q��i�������O�[S$��I�I�CK˖�O3�O�w���'.O]�pڷ�'��%3ݝ=L��[2۾z�y=�ю�\ݝU��$��j��ᮮۣ6��=�S�5&�g_���ɗ���9�?�e�;�ojÍ�2��a� ����lY�>��8��I�M䓍��pt؊��i�ַ�j�c��.s٘*38M6���������QݳโLI��������}o/ݳ���˓Zۭ��qyƫ^vD���?����f�n��oXlL=3`	=9Ç-{껱w��|�>Y4{�"��׾�����-=�v�GC�^N�
�`𝯓^��07G/s�Y�v`�؎�k�S���=�ftm(�u�]��ew�fX7|=}���6��s����F����/c'i��vq��h��{�HDy��r�!���Q�U��+,�.�D{ <'v1O�BxT_ho~���^D�gs��wR7�~�!�l=Ԟg�Q���>�{���q�_OxY'�¢m{޷{{!�ᴓ{�}�����6W/]��<>�4�2Nc�6����3��i���Yѱ��1�{޹���_vs�z����1/w����R�i8*҆�ޞz�?�%�	H����<^h'5�/�����v�#��ɡ�{��᫯��AZ�<��_���I[�	6jm����a�x��7`{w�v�Xh^}�,����X1v9j;��Ӈ�'����z�����q\I�8�Ѹ"�.Ԯ4�K&`�~�Qפ�a�
{�8����u�.�;g�7��L�oo'��h^Q�^�k�OJ�b�BW�~G�?4�����>z�NCݽ=#�������ď��K�7�o0��x�x&���7��Y`���}֑��>���ow���H���[ᛠB� k�ݫ�Ȝ"�Bצ�-I���x9o���}�h�o�[+��{YG��p.�J��C��
!�'�p��4����G���'�J�g�`ýB}1�ޱ�y!��t����ƃ�"qH��揷�k�H"�� w�c��g��c�/+gX��ȭ������nݷ�zw�n��Y�9$�N�H?,!��0vtk-E��!%ű�H(�Y�g�כ�}�(I/2���$�>��,�)f��u���<����	z͏��yy��{d��t8I�[��p.H'���g-�Ds��%rAy�dw��1mm��6�f��ۯO���t���u�b=�s�ZL���B��G6ݝ�-�D�̭��:b՛�.��1y�k�g���ny�G~�{p�v��4~o-Ε�dI�I��K޷���>�??~�m�_���o��������%�Yԉ�YŶ?N��4�i"�PE.p�fla��SVv:��w����0�pv�3�տ�7�o������2N�&wcѲ��M�8n����q��j����e���3-��y&	'&J%�e��i�[�[d���0��6f�S��o%.OD<wI����j��ݙN�n�8�f�^���	˓����]Yݬ�/\�luh�3�gl[W��������9�_t��y�3Z;7:�k=s��8�`�p�LM�Y���2�Xts��s^���3��m�	����k��IVƝ|�{v�ya>�z�\�&	"�Otb�����DgBd�w�^���%0w�&&$�+�H��U�mz�c�&�8���rlG]�p����Φkk×�3!�~~ǃ�.�G����G<��Z���{�� /y���M#�s[�N��T^�A������CVUe�ʼQ���i)��Ͱ^�ޙob�	0I����'�-�qbh��h0��a������װ�&wz���7v�@��߸��E����"b
a�	H��q5�g�$��4�Z�v듭�4`��iKJ�A�&ҟ����O��bLy�{��|%�_`M�INW��v�8��/���I����&�t;*���'��:2����y��������J,S�Qw���Ş{�qv޻��n�#Yl2k�U}Qa�L.޽oRd�Ri��Qw���y��,o$�e�̇��-
���⩣f��,[�L��Y��
��$�	2IVLm�.���{r��l���'u��]'�$������K[T�\���֨���H8��{��Jc��o����<�;;�]K?i���������{������(��0����1"���\Y�Օ���5ţj�n94q@ͷ[��u#f �۩ttЦ�;B6Bif �t� ���y�P��IfM�b�f�6eDu֌E�	�5�F�js	�Q��Yp󦫠��if���X�d��g���z��i�n޹f�#q�\��u���x�>�����&�c��v��q�NT���׬ޭ��\�t9j3Z��Y��e];׿����ͻX��VD��'k�Z���xv,��s�ܰ�Hi��HI�	6������Ua�L�o s��șW,7��'��a>I�t�^���Yߘ�x�Qeu�W�8boo'K��5�MwL�]����t��RE"^�u����*�諾�0Fڼ�e'����� �9�Ƶ7{�7E�^��d�7.��r����g;xz������0|��$�$��$C�6�5:7g-6+���CB��t�orS��	w��i����`��]��V�
נ�}ɹǑ�72`�0ws�gg0H$�Fd߽���.��v�n����3���2Z��mhV�߼�"2uכ�N��`'�$|��z����=S�K?��.�w������L��ĸ����*��q���s�ow�v��Lz�U�1Q�b��F��1՜��29W6Y�*]Qk�h����Ds�`6������6.�[�v���I�Zurk�=4aB�=�XOs��&��Mgv��UCj�r��C]�3�7��%>	6���ai�ǣ���،b�r؅�I�/t���3���Z��u�i7ر6�=2)X�m�$���o/Y���;o����𭭴ې�ũc;L�oz��)L��3��������_4����3�[j�Q!�6�2�
b]-K�@���h���>���������^�O�r�z]�3b��̓u������$�� �)����E� ����v�5gly7��^w�V<��`�f-�f��f;�˨v5ݥ#��|Αy�s������L�"睧O����tݳ�#5T�p�������$�8�s���<����c���W_�M�R��i���5I�kaD�̺ʗ�	U��g��{�Z�J|��AWU;��MZ��u�[���x���{Wf�g$��MS����m�I?�oW�L�-i�%o��s�ۡ`ї�����]^w���o���;�𻱕�r�4Y�w͇����f�][�k���#�l�L���ݟW[�kՎњ�V$�8�H�ً��{��O��s��኱ҳS}eާ;z�l0�k�gK��`{q�ȫ�� �q�3g��hk�`7m�Ҿ�󱙮*낼�0c}ΐ���Z��X�S人1�kMdIC^^C��Xz��.��0I��JUGO�Z&2eغ�ǻ`ol^�]��u�������6���;dIr�4!�ĵqI�)���Q6b/���F�gk];�:{|����=j*;��as�'НkSz�����s%��Bw�����&�I:I:w �����]��h��vkSU�fh�oyw:LM�춻�l���v5���.��<�(����n7�^���V٣P�[�Z��~�_������ݣ�`��؇s+
��[;#\k�>[hU7�[�$�}I�t���	�xa��W�+��u����R��5����2JgA�9�����z{_�I�o�Dc�J�41Ӯt���yW���h]����o]rS������;c�#+�1^ �?ry�
��u׻�ea]W��y����ߕX��I��`I��f�z���i�>��&�Veꉌ��CEV_p����Q�J��f�W9��tv��ٽ�݁2[��E�eL]S���]H�Y�"v?@�H�xs��v[�~����C�i֪�tҕ�{�/tE1�ʑ'-a���������܁�4bK��q�s�U���7��d6-�RC����'����y��l�YHLq�t�қh��ˬ�%���R45�S!�[bM� dJb�R�
�e���Ib[��i4��x2�8�i�-f�b)�۷k<��",Z�̻�Fbi�3e ��\h��X�sԠ�v��Zv�Vz��N��[8��ϡ��6<�:�u�QsGV6���;FS�*����>��*�lZ�*�ذ�t����=lu��x;yu�W~>��>��o���T�:1�:5�\�"�4C+X[$U���y&���k�4��!v�|��Ѹ0oglC���u^p�����h+�j-ػ[��M��I%>�V.Clf�Ag��rVS��Z�v�K/���V�'��d�k�uD2&Li�O����I���?V�����U��S3�ث����c=������?�L.���yu71nn1�X�F�t�(fcn�A����8�qI�M�T`�ii�;���qᚂ��/4�Mic*�K�M	���+t�/mϒ��-썊�۩Hy��;-y�.�$�l^��7}r�W#/�)ɬ�0v�P��U뀓7�$���n�(���iy��_I��4=�˃vf��H�vцw���M .��y�V!É�AR�6ƣ/1g�s)�Ѕ3�!����a��*���>����Ĕ+��[�0%��D{_���(��^tu�l�p�3ɻn�U��6*���56OU�z�������v�&�}:N��2�7����lM�b�n��r��b,��c pμ�\�˧r�kġ$��{�Wu��:�47VVG2��J�t޽�^�~o�������U۴0��2�ˮ/�]
J��R\#��i���,� 6�~������V`�{�ޜ����i�3��eRDvvys+a~"���m�]ǟ�=����sEX^]*�����T�{.Z`����aX�I
�]xK@�+w����}���I�I"<�Q?ǆԳ\�~��=��Qt��Z�2�k������y[#m��Ϣ����y�}������t�����7��R`�X%�*-���5Mb�y�*o_s��7��vԱn�K��v�k�p�_[k`��׭y��Ϋˋ��״�G{:X{{�$ޏ���O���Ww�1m�nV�嚓U��Vµ�NJ5��]]����wo�;��~��g.�rmI�[�9�J4K�r�/�G�u��f�������]k$�$�UV�Kk֮��j�J�FR���޳/�����S5���y�v����!���ml�N�4�LgU�{'2<���V_��h�q�)���$�&�G_�m���h��靻Z�rʣ3��*���u�Nd�a�x��|ę$�5����]s�R����z�C���c,�*c����ؙ�Z�C�鼺+����(S����<_�͆{����u{"�s3p���c1�|�]ax,������$��$�-smϫ���=.��v�}tے�MS�W�N8�	0	'��c�0��� `�.�Sx�a"�,d�v0H�&s.9�w/��rB[��4l�Q���A���$�.m�f�>Y�����@�t{�������wty&��$�l�_m0����ш
�qSWxg�9E�D�RY�~9-�޻z��$�F��U��U�	0I?�Q�y5˥���ͩl̗y�����I�L$�u�[m�y���W����k$�vkyU���5t�>_w��g�8�x�s���5���w2M䓀�X t�>�C;��wao^���|������\0��I��������?�]c�� \h(������p���L~Y�.�!��g(��A�,0++# C"�
�#!̋22,³!!"rȁ�Xaa�E�EXaQa�=G�a�E��EE���(���@W#��������E�¢�+%¨�ʢ�"�*,0���
�
���0��
��*�*+��2�����(���0�ʊ�
� �*�0
�� Ȫ�
�"�2��ʢ�*�s
���E�XeQa�E�DXeQa�E��E�EDX`"�"��#0�0�#�#� C ��
���0�0,2�2,2,0�#��:��`֠�����(Ҁ�)2��0~����������;����?Ǯ?��>�����CG��>������>|�k���� 
��~_��������vȀ�*������D��'�/���~�?p  ��� ����^0��}��4������ c�����X�8Qe@E
EE�QiE`fQaQ`�E�EUEQQTE�Xad�&E�(�)"� H��B�ʐ������
,� �) +�,���� ������?��� ��� �
Ѐ-� ������=�A���� ��;����  ��~8��q��;8�Oϔ�f�צ?w�N�� |d>�������� ��@ U�~H|a�Ј�+�x}=�� *�?/ژׅ�r6��C�Ow�$��}<�@� Y�����|A _�v�Z�Ϡ~?�q�����O��C��C�@W���� U���p|�C���/4���i?L�|�����6��s�� U�?ajjg�Ϣa�����?��t����e�*"����0�PA��������/�0��?�b��L��xRDl{� � ���{ϻ ����o~�AD� P  @@   
   @ 	 
    X }�    	( � �(@	PU� 
� 

*�� +<T�*QU�T�%*���(T�B(���H�UU HB�JH��*��P � @3uR��J�$���P�}*�vp�ݜSw}�NgNRW�gU���J�wR����J��RRn*�t�9b&Z��!J��R� � �  כ}� (O7����� [�� O.�*Y��K�TT�A�{0�h�;;��L��QS��R� N��@��%HB)TQ���))��S6���=5֋g!�R�T��{J��%U3�*�`2���%É7*/g��z�<�U   | =�����D��������!a�W6"������V�)n��tFmTSl�`i[���)UO| �*"�
��*���f�F��٠�CE_w�B�
wgT��-`�
��'�n(-�U �O�G��W�����n �6b����Uݝw��Sv��2��IK�  :H�� �$B��$���R�<&��[�uE�T�wp)n�F�Y%6j)ZЊ�(.षkSvt�P � ��̈́���>��U�����2 �f  k�dd�B�� ( ` ( }� �)@UT���(%=P��%��P��4U��0 ���i�@i�U2n�J�G%�t�  �^�
 {��4}�@+�`uN�:�[����J�����)�:n�@S���ݺ��:=@    T�@%*Q���dƐh�F	����J��       ?L���*i@�   F i�T��"�� h  M  	OԤ����i�M1�h� &�҈��hɒM���12MM�'�����?]_��'�@����D��;7F����wF2�d�$�Mя��!gА	 ��J!0IB�@$�	r�a �,��g�?����G�h�<A���	�I! )�� BH� b"��IH��ժ�b��?��>o�d�B@&����%z1��i�c��n�w� A?��}��������	:7+�,Qa�6e���r��f��Ӑ�QKI�<WX��7o�!9�U�7]�i�a�f��A˽d��h#���U��\wY��$��z���w�ֹo6�*[YGJ�)A��q���q�؂ܥ�#�)X��X��u����ͽ�BQդ��Usl����wi��*X;���5�]^�r�w)�z�6��d�F�d᧔M`��*����ن�-�j`�7j�e�p��x�1�#R��^�Ҽ{MA��k7$lx-_�e���3Oc�¨��܉��ȼjD�Dc�B�ۍ$�n�@�^f[Q���Y2jwU���[m�ٻ��C>��KoM�
1�#��S��XkU���~C%�Xd�e9��V�Û�Y��B�c����e᫁],Ӌr@���DFƇ+t����ˎ���KI�Z4�h�4�e�b�Sr��&�&U�,H��Ƭ�xqn*- �)�l�9i�L�.�T�r���V��n��T\za;#��n'�����RCX���C1���:�Pbg]%F���B�k�s���,�V�/1�Lz�	�:�P���xr�Ѭ�BzF���ޢ����[�Z���:�-`�����)�CŎY`؏/�7Q�X�V�k3
��b�//.�e�N�h����ڛUv�B����]a�kI��G��J�m��.��R��.i��-�H�LP_7a�t-�s71*�@4�mZ�aC8c>%;�q.>�#���P8l�%fnQ��Xnj&�bm'������7Wt��K�Ǣ5%U:�6�55s�����5Zu6���zq(��Yqԥ���=.QR<�:U-ݭ���sq�Ę�0�PBJRl���5Q��2�Յ�
�N��a��Y���![F�MY�����S5���÷R��6��e��9yF+2���^�"u��U�,��7�]�Xq<�/�DB�M73�����ۧ����w�Q�t����zAI��eED`�HE
R��\���ۼ�-��*56��0*8�p�/5[���S�V%YYN��ݭ6$�tɖ*'[u�mc��w(ɶ�qx�j��.�m��HcN*;8��r�NZ�ȲG��͡�xj��W�4c�q]}��>��\�4�dЄ1�fG"&^C�K��ǯ�v�\ja6j�9`ʧ�S2~�,���W0f�ub��dE�T�f�qƩM����ݰ�Zc�AW�ܺ�V����+t7�2�i�1��G��/*��2����UGri��M�˼�M�ҍe ��������?4X7�2J�uv��9�l���9V��6e;	i�+�.��cY��������`�(�NR�Q�UV�E�Yʁ�Y�Q�6��2��J��h���jKͱ���RUM��ڱl��&�aQ��*20e�Z�j���8X�J�O����Ӷn�֦^7��a5.�ɦG"<�s�h텔���b�j��7q��˻��q.W�N���H���&Q��1fPan�'p2sor�V��b���s6RTl���75��uV}G&*YI믫.`QÖ��*�֜��6&��m��{������,B*,��*1�Z�&�ā�8��ڍ���%�Zp���3r�e��yx��Բ��Q���i�Є�v�iyU�iQ�hK��uusE�J�,+��H��{�V�-eЕ.T{� ��kW�]f�R`.��F&��KnS̻��l4�n�*��l�yy`�{�jVܖ���-�Hٛ.�QB����k�3v��ie��9�rL��I�*�qH\òg�1CS�TB��T7,��͙��B��.�cm�N�5*�9��ȵ�'peݼ9@��HN�xa3Eafm��1ݝX�$���0�wr��	z�NUj�F*�C�
�gG^DDV ����1K����.��;b����r�Q�5{�0�U�1캐]�JJV��K
V�
��u	�Yy�]曆]�O�zWr��*�*��ʔǹx�4`�umm=�,ٽ4`����̿�,u�"��Y�]—-=�FD6��*E�������'K��J�]����ތ�4�C6�e�As�4#SP-e��q#����T�
u
a��;.�0�_ek,��kr���b��S0o�-r��^���ݘ�eT���j�]�9��̗eE�Gr�Q+	X�����j�֤����n���h2Y@����J�+�vĪ6���/![E�&�WA�X��"�r��W�zouJ��ۅ��F�1ɔ��8Aj	t ԅ��d'b��4��lM�#s����ǿi�V7X�%���K/b5`��a��1�YX[�Ecm��l���RF���j�����5U��W�e�;75M�]6md���.�nfh�j�Q�D�a2УoojB��S��\ۙf�:�T��d�[(���յ���f
�y��o"st�zhUj�zZ�Ԧ��+	����U6V<��R�YQ9&��
�+:7b����A��oM�ǔꮱ.f�6�*��)��pf�C�cF���δMӏq�i��°\X�Z�3��q����-��Tr�֋0�Ʀ`5����5��Q�eBj5����[)�ׂ�q=+˵��TЧ�U��V�V�x��ܣz	��G�Q�U���mq�Q��^8��!Z�d������G�r�e:�u:��f`�.�(]��;7/5�z���v�*�n��j��A��Tx�Tki&��d��ş7�K���Z.�(2�6�^m�v����2L��5��3/M�b^d��rI��kD�f����І��M�4X��YT��A���p=ڙ�k������!h�tج�Ku-[wE�N�R���4��f!U�:R�O�/�z(e�+{WT6G+$�*e�7��:��s���Τ�=��mF�
f6����J,YMٯw�L����*z�,��]���R�c�<x"j��H��Of!6��M�-�U�P�6	y���x��4D�FQ�y�h�"]B�s"ByR� f��R��Ȁ�`v�=�z��;u�`�Z�B�r�ֶ�Mf��-�1}J�<ۛq��ѥ�-�3l�f���,�p-�K�a]�����kv=z���w,1[�Mݑ�R����f7���.�bz6��lm��0�ڗ�n�1��4踴��MT�Ӵ$��t�p�"�V!���D�nDV�K�x���W�0U��Ӕ^;��e��+5�;g1�r�ǔ����lYT"Uac�2]bL�^Y��6ʭ��.����6�UMT-ùd�5I츯Ud���
2:�m�R�l�KU����(#a��+i��/�5nhosb�Ř���B��L/p���֨t۽wu��;��N�c�)�"5����������Qn�|sc,�L��X��u��S��]�SŒ�;۫�����U�)]�x,��5�U�R��ɘwr^�k��f�l���Y��4�5w���.�]�
�/�bF�%4ꖵ�Yeҁ��H��fp��h5ote��J��em��M�&�w��mU`i�
�t��b�;ktDr�m�f�#���bULjr�]m����5QxvӘ&h(-^����up�����M�0��S��DZL�-ʼǸ���U�؅*��l���<�ݷ���!���`��aEd�D��ҍ�ԳY�M�B;ʰmU"d��e�1�4��Mư���%^����Ǹ�c�k��*T�m�c��9�����Onۻ�&-ɲ$��m�ʕ��Q	��dW�/r�^*�B�ڼDh����8�Vz�G3r��80�n�b�5E<�(,ъ``��ˊ\g㚩�R���x�n��CM=:��j���0��|�S��B�Y�%˪O)kF{��r
L��Y��u�S�Yy�[�;��U9�!�3-���idLCe�M�P�XXRә��U^��ۚ��.�˺"���S	꭭��P0^���ݬC���fݍŸ�V�W�`�j\R�sn7VkR:�ǐ^�C��T2dt�J[�{GuLV.�ئ5D�`��4�^e�n�h�����v�K���۬���Yv�^Y��V5�/I�l(��9Z��tWb���$Z�UUP�h�9u�j�����S�e�5�p����92�bf�ܻ�x��ו�-9���b��n�h,M�p��5�n(G������C�"dA6�Nf�[��ȣ��TL�9�"D�bm���f��3�Yb�X;�D���Ywi]��N	uTʤ�M��W�+�ތ�푕U��UK���6ko^L:��a�c��IW������n��fbl��hmnl�eG�z3D��4޳
ݧtBڨ��
n&��Uy1��m?���>v��"9̓���%��W�.X� !G"���H�[���I;��m/�Ӱi;[� ���uBQ��p`�v��rc&H٪R�9��:�ڠ^����ڃa����e*[G-٭qMw�ld9�����1��t����e��=��f��.ڱ�MZ@�Y�BՐ�f=7�srfJ.��Wv[�Z��ɸ��T�B�f&V\��^o��'VF��Jn�5��Z&����ɰ�aꭧ��7-UK�l�X��+�)fkA�c:#[ZN)�^	���,��md��]�Ӊ���&���Ԇ�'�g��0���Rr2�2%:���"�Y�^`)���Ce�+&�����v^�Ԏ]�H-Z�z݇�C2���D7�y{�j9���Y̽�����^欨ⷂ����&�֩�Mi���45�une8v�1Z2��u�A���+p��bVAt2�	{+k0^,;R�̭���^ʗj�hV�b]P�D��Z�q;�o/eҼx1�nܳY��$M/3/3m#2��,n�/#�uv���NhR�D�Uts0�[z���FՆf�8c��۱R����5�.�Û��,���!w�B������%V��{��gH���r��pU\�y�
�n�eei��j��,=�ICl]S[.)�eE�#�y�+"B�Ͷ�-S��!eUb��m�řfT��ڻ�1!�����ݦ�6�eRr�1�����wx�b��nd�+1^�ȡ0V�Ul�ڒ裌��˭��Y��rث�%I,os���V�'���Uv0F!�����2���U�̚"m�{{u2Y�3tL7H���n��ï%ʻћEɳk$����37�� 78����]ؖ�k-٤e-gV�������#��WԨ*�.�D����U�e֬�GQ���P8�v� ��5U0kU���^�e��H��m�BP�vV�q,�)�M�s�wQ�@�Th�䭷�ۭo��3u��E(�W��Y�����[��,Z1�w�gv�W�#��-b�U�v(�oD&�ь0���{����ȩ����t]KyE-Z3�Ŗ�7%X��i�Su�@������i�zE�Y�GkY�3�-A�nU���Z�A{�ܻ�XPֱj`���j��ڹThйoN(���Vd�;�<�{���i�R�:�Uj96\������(̣�{6�Gpd��lkYI**�.�ي���!�,���U��S�[͵a(b���vl��`6B��U��bɢ�a���:(�v��RE=���U���ǚS0�*����/Y�Y�R�P`0*���:u�±��q�)�F�U���8��4����ȨZ+H�	LŌe꫈���*�$��um���k�8�!VQ��"�p��NЖ��)�{[��X��P�J�݄��
ڎ&k]S�[U�����֌�������{�I�"Q���H���,�OS�P{�$�� X)$Y
BH)
H)@B�!@Ad�"�� R �P)!,	"�a Y$�!$�dP� �$�I�,�,�(YH��		$�a	�E$�P�"�
"��)!$RBIH��� (HABI Y,H�� 
I�P� �E�U��E]q�wQU]� H) �HE�) Y! P��H) !d�d!"��R@U $"���:����.�㻪8)���}O�������W��� �+�N�{�$�'��� �Cg�݀��������o�Ð����Q���2*�db����]���Ⱥ�I��]ghfi�5X=���>�fc���ff<����U��rT�;�J��USJ.|��j�:%���~+�Zƻ�������=x�j��J_74��7YTD����f����n��i�uB�<��o]�Qn��ʮ�2��<�OiG�[���&V��+��_V�.̃��,�U�Nc!.����8M��v6f�k'�UR�s.�u�}�$��S;�~λ���=:��U��y�����]��̎�N��'tnո��3%^�"3k�Z�(�8�V���� ���˧�NS�ɋ��ӳ���+(d:��s��[$��ٜ�s��.��@��^�	ăC]��v��dW2���1q��6޽P�W�6�=<���{\�%��W&���!��J;Y4A�PB��31�;�>NZ嚩ʵ��Hi��Iw7sĞ��Ce��w�w��-wz��ݙRm_���T�e���m<��2���S�������ޫxi��|��׋�vs�g`�.�]���Q]*c��<ݘ��׹�!�>��4c���<}�=�g8���Y���69��/����*�.���i�.��M���T���Q�sZ��xv�TyoU(���Jݳo�y����v:T�����v�J�+e�9N霼j�f^�e��S7l]�$Rt(��5چ;޷�w[��dx��Ջǂ�fÛ�����H�]O�v;kA8�c_;��>�o�Kgj�AYL$~�ݍѨ���v��6E���������WA�����9]�bv���h;j��r�fF]V��}�uL�e��/2;�N���VV(��ق�4z�-�a�S�U�!�&�Л��:h��d㻆Ķ�b�$��Q�����IA�R#n\V=ݼn��D���`�؀���EE�y�T�"ވ°<벟>��P�2���Q��=T�ի��3#�X�O�J���C[ڥfV˛�#,u��!]�T�%��)�YwOb�dZ���k�X�o�>ɐXe���U��
�.�a���ˤ��n�A����d��q萇p�4��3NR���WcB��<�
���uo�Q�ۮ��6mil,v_tW]u8Ԯ�Y�+��dj�%ղ{�5ʼ{`�`î�R��rј]eV�j��Ǟ9��=k{6�PJI�z���we3W�P�퓬�2���D� 2{#��yL���e�ʶ ���T�sV��J>�Z���×�F.�[7GK��E0�僩SW!������n�-�ؖ7�]���e���wu�qZھXr^�&l��C+7��NNt;7M�w:�fl��W�^І���w�D�It�]r�:�u�-�,�Yu\���嚤he��9�S+u��tܻ��f�Kݕ��]�i��,��B3F�cWkF)�)2f�^�������s$�B�7������{s����U lPUX�غC�2ph綻 Ն�ñ]�L��Gn��M\ܢ��&HN-�QQ�={�jkq�j���_�ֶ^�6�k8n�*`��݉��#uK����:��lU�B�p�}���Y�ֻx.2�%���W�F��5���oQG�Ɋ�蔙S0�7]��u͔]6"u8k)�sL�N�mf܀�dU-�o-u��kq�������jUY4F�'K��]R������]Ü�ͫ�����t�����l����f��Y{���>���UF��b򷎙N�Zv�����ΫVu�-�.�F x�YUn��7�eU� XO`疹�ī�Ua*�8+�S�p%�{Zk4�*65��b4���N�[/]\�;���Z�0�&���x�����a7�y-�
�+j��\�8&�u6��[:��s##w�i�vf%���D�[���՘wslڽټR�c��Yys�ݵ�vfuk�8ݱS=�����cv�
}4m7E�](UV�������h�V�;�y�c˥8�HUj.%�=�9u�q��Vwi\��ΥnkȂ:�,�w�d���֩g1d�v��p�~����Ϩ:��s���^=���r
�D.��C8ˍ9�K'vff�D��Ӱ2g6Z�U&���[Y�I��%:�WYT��x*ɊAZܛ}W�t�3{��
�W(��̒���6��vf1K��2�3��\:�r��F΄�Ό��dVުy�-�aVZ\��ۛ%�Z��t�N���_;�67eK�dʗ٢��P�z��v��9�/d1.��ƚ���z7�-�Xs5^>��O���B�CiS����l���w�ֶ�)���W����Q��[��i���(A����"�m�J�'2M��8'uҬ�/1[���J�����l����ux��e.�_m��&
�'.�cF_K�4�ɾ����v���WF�*�[f��8��5�:�]K��;[]ɍ9Ge��Ʌ:�*e`C��w:��o��ܦ:;�B���^�I�.Zou�+�2����p��"����yy�����/jŎf�Bb4�v&��� �ݖY��JJ���{t��n�Tq�(l�q_�O6�j�aɢ:;u\�j�z�;v�.��බ�U6�%�M<ԙ��1��D�'oX�g"E�� �Բ���T�ەFm��	��M<u�)��TN+c0QÏ�lD��! \.�lL�cLpݳR����qK%��t2�P���j�}Z��jLAk�7+0^al=�u:��t�Y7�yæ[�w�Z�f<9y���^���Q�����^��>�9rfU�m:#�m�ͭ���0os(ެי����i��Ƥ8c$\�jֶSc%���,�ӫ^Tt]Ҕ�X�sm��'eM�EԴ��f�dٍ���r�S\���(-bg��|�'�4�ȍ���e���+����*[ƪ�з4-85��]%��ʽ�����N�+5(��KrҶ��R���A�̙�C1�b��b}�s������݂�hm�Hg%F��tv�,���c��NEd���I�&VȘ������gZ��m�C����٪b�I%�w�ߍI��ֆ�-hD\�u��ꋲ���v��\#-��A�v�P�mp�ʪ������B;����v�!Ű-��@X��:�̖�m��N�%ݽ�8|Mc����3�n+<��t�u{��C�������-�U�cP��*�1Y9�N�b��𱖠�y�U�м��9�G@�u�vn�R��>B�k9��w-����S�c뽮�Ue5���O��#PnC�ͤ���kjWc{����X^U8���c�=� u��6�fX�9%���V�9����2*Ɨi:�<w�-�wB�?hKOwǴu�V8�Kun����%Ō��Y�jk��++.�!�P7���EJ�[Q�n�J�w�V�r���'I��6�JS��Mc��;���=�cϨ7����V4d��y��:#�ZWً�V�n��PR�Ϻ��>V��椶�o�$�����RD�Y5P3��:\�(�b�vNCy��.=4U���ȖuqP�w{�����v���O�q4Y��2Xv��tjDht��\;���ѽX�<W&X��$;�'6wr����@��B��+�擽kr�jڎ��}j�E�+�#�g>	������&�d��.���r�����[�������H�]�t-iJ�z��]�:��e�pWY�,}2f�2Yy�JympF�Ʋ����e�tט�ܳ�'t�#v(�����}`6ږ����ܖ'sK��'f��T�HuL�#ۻrᬕV#fb���/�Zl4�A���Uфޱ�]�	]ު�E{��1�U�7/���_#��8.�x�t]����~�!�v�y�Vʑ*�S�}��q;;*�n�Ibk���5{aA,=[�vsܱ�ұD��`��꓃�q^!'X�9��Ty	���3m�h+�Vؙ�[�_kǛq�U-��n<:|iX]�Uܞ��O$��˞��;nh��:V�c68�ں�7���+-����*�d��<�.��o=�]�.��n������5���%��E�c�����jC�
ٗSo�I$�]�9<����45[���K{�֫l�iXj덩��˷]�c���6ƺ���S��fZ�7]�_|d�ܤ��U뱌�)�G	�Xs��@ӽ�Rn�v�̜Q�$wؘ�lιhm�7���w�e<��cY[rb���l�pl�c.Q��3�ټ	�guC`��8�W�{�!V�`���)]X\��9�U�4<�R��쯭���H���=ט�aZ��p1���~��[r����EF����Vm����!���٘�r����l��lwՠ��Z˶�e	�q�]8L�́�j)ލ��Zw9/�6�C��!\���׀��z��٬U嬧W�u�MTx���u}}��|j���?J����_qo��R�2�s�����$���f�Н-�N�Xr����M��.ŵ���Nvq�4ۺ��ޤ�
��ܹ�,�-��G���1iYy6B�dΑ�F�N��J	6[�u;���]]����hm�f
�\�G\f�X��ݞ"�x㹴��mUr��\5�ñ�wݛ�k�F�U�r�}��3.�^��;�@֙ڻ��J �M�&���f��sOUڭ. Sn�����z��r������&"^l�Fn��KϤ�6���ļ�Y�5��Ae(��qS�q�
k����#2o/�"X��UNa��az��+F�H�u�ou�f�=��5#�Q�%7JU��3�+V�b�;Y�(ք	L�AX��۹݄_w>��7��]u�{u��,�*��F9�,F�m�˪�X�7�j��'E,W1���5,�NlWs'�z������6�C�N��,L�Ub}�*��9R_uX�cw��3Y��#p����0Y`�c�L��=�����fsa��Bا|�5Yh��uf�Kp�=ժ�0Y&Y���	{��cY���	2������8񾘕mnm.X�W:��mAy�(�����U��{�Zfe��%n��eZ����T0��c�2���n�+�'3w���-�ڮ1u�!��rmN�34�̬�̪B�L�⦷�mJ��?���@�*��q�ƞ�ڝ�x�5w�ۑ`b٘�{����f=|6u�o&թ��5 ��=���2��JP늷;m�1�E<]�S+t5��U�r��8��;2����zI�0LiMt������7�r�;t�+
q�DXXn���e���7�]�*�ޔ02x�g�V��U�smi��Y�:��̓��^��`\*ȫ��Ƙ�h*f�Uy�ڥ�7�[c;!{XU�)7˳���l��,��K�tq8�u��𧁫jFu��'Pڝ����n�7P�����Ѵn���j�r���f8w�&�'"=�4&T�.a�:5��R/P!��m[x��*�ιD�|�A�=Y+vT�a+7�u�7�!9��T/�B�TǏs%v�"���h��꠾ˎ,�.��hu�otu�l�ٖ�=MQ�*��T�t�^K��fS&a=�Vi�p{�²�b��:b��I-�i�C>Z-�l��]Ҭ����Ť���`���U�ō[AX�vi�w�2�C�I^Jx�n�s�t:�,���V�ձ,9Q�]�E��|]#���lUuuv63lntLw�q�Ν��֙M\92v�,��!Y���uX{�-��f,�UV<j��ܳR���lu�K A�����dV�jQ�\�Se�Lɥh�L9J�S�]8:��N��0�n����\�!2���sCC��T���ޘ�8�aP;�����9BEB����j���ct6�p��� �+�isù��;�뾵Z�7ߡ=��B@"�_��k�,*�\;���������K��m�J#v�	+�`��t���^�֎&�s���u�`��\C��W7TrZ�\���N�ִp� z����]�s\y��ήX!���Λ�tl,�Sk��ј1`��K3�Ȏ.5�$�e�i�+�:�&�Йn�R^���䝹䎓��e��x�s]8���-"7����>K�4�H�Bb[kels����	���&���+v-zG%�ñ���9�vx��nK��w"m�F�6.�Y:4�07Z��p��^0�� s��]U����Ya%�XV�bkFn��Z�t�s�;�W�]Y�`��+)`٭�͊��"S�Ꭱsn�E\���<;8��nK������;Ԫc]�F-IB�b��0�@��,����ø������l�qi��v$�����T�n��^��a�6�u��ٶ;^xvhY���ʞΎ{�I���N������X�p�K��e.��IK^��f�܅�\y�e9�����Ʒ�b�K�b5��W�<��
���śh5-�Zd�0�4Q�%�jh&�����n��6;i�j7��u�Ό��cG��۝]]k#�ېSquƖj��λ]+�̐V��(mBmlB�V4�B�4�t�\�-v��Y��Bɳ�b`*i��l6Y�����B��H8�:��f˶�*���/F2]vM���zḖ��b�KYb�ZI�mYm�ϳ��qs��7eF��b�-;	uծ6@<c��ʜ�u%��1��e�j�]���;�\�٧&&�WK4�����ŭâG���:�����V6c���k�ȄI�'i�p�vb���v�J��4`Ыd�)0�k��l����5+�+s��ۉ��uWg6����'[;�W���0u��w�{Sѻg�-F�a����jɰF��m�퉈�`�,���.����]��u:��<�E�m��@44��n�7U`�lՈ���ф��m41�ZJ�髬��|;.1uہ����g"�p�g j�t&oQ����
s����K�9�Q��B[X��o^q�n����2i�xt�)1C��Eq%.����\1Ǎ�� ��!RvD�r	p�m*үי�r[�@�����a�M�)��ݗ=���6��G�������*\��N=m�2Just�Qv��˸�&��1m�P���:�,-��.�b����Y�lɨn����G�ar��.���)��C'��,k��̠T{e�{y#�4��9�uS�Y�w�q�[Ba0�ū��sa���J����G q�7	�nk=�&�NA�Vⓜj���rq'��\����U�s�Gqg$��s���=l����:��y�{'LؙS�i׌�=Ոz�=\됻5ۭ�gpl�aV�ac1���<�M	���g�㰢��b9-�]q]��V���}�$Q6c�X��J�m!�k�i�#�zۏV�=<X<��9��\U��ܡ Kd��n1��^j��Mo)w�h�]�]�%&�I�NLݲƺz@q���V%jW�v�om�S[��8�k�E��r�%�=���#;��룢�z�;Dܷ':1u�o6`�{0��\���4������=u�S�M�!�5ת�ۀ����h3c3��q���W$�3Ü�Μ>�J��1����Fn#���2X�1�V�	m4j�;\�2�YcNoH!�@Ջ�	;����tʖ�Ǯ�gL���K���A��[=u����Y�8�.�,/CVM�[sp'++�	n1-�{!��;�jH|���ݸ+���*-3�����yLU�����[Vq��6�Lcs���s�ctg�溵��٦/<v빠ǒ8�p����M/.�f6�(�ql��ma�SX��3u��j����y�f�a��:ll�f{gG!�C(C�lK`�"�+-�УTJ�46�j��S,��^j�eq5.a��k�vZ�K�6�l;���JG@��l=��ͻe�l�e��#��畤�r�$�Ԕ5ݩ&@;K��)���x�kZ:r��KP��9wݐ9z^ܩ�-qV����k
ͫ���on�n�� �D�b��m3]����������ˁ�a�e��,8����m�v��:�o/]�G�������=�$űɴ�a�孃B���n��m9�`�΄O+��e�+Xf����rVbxFԄ���Y�9coTw �<[$=/jܦ�x�����q�u�{pټ���ĺDĹ3,�|�T�͡-��:�0W[=v�v�f�	l�M�P���Inc0I[.ݲ����)�9�Wj=S��x�-լ���=m�8���k���:�vx�d�g�ṣ��F0v.��)jl�L`
P��G:��-�%�![�����hzz9�Iu���M��`�-��p��`5-�^d�V�q�u�n����`����P�q�7���v�tL2�V!���#����J��H15���e�3����A��<�,��ѳ�q�b}˷�)�V�+a.,\Y��\b��b�)ӞL���ͺ�5����yeomC���j�xy����U
�s��b!t�.��5��0eqs�*+�� �ucgS� �6!I{=�i�N�=rd1�<��i�0�`��	J�ān��m�����4��VƘ�7,��,%�b�%(�nf'�Ν��p�+@fū��0D�6�|]�y�GN��si�ױ�8j�@\��훱��8��/��q�kn3��������kB���]��EI���r��,.)x4�U+w]Q(6��"y��x�K�����Z����P{����kst��n]���溱v�wI:ܕEg.�V�k^vx������ۯ1�.�qx�m����f�G+Ըu��<�v�T/ksr�x���[���v�^8��d�
݌�r��!�kJzݺ��yBՅ��V�u�s��k讱��O5��]�3ٸє��8Cq)s�=�e4�v�u[ <��x�`h���	Kۃ���yC�ez{�x�[����xCuN7;���[�n���ʛ9{zM��u���Ӌ��f���(%ڳ)N�+f��+��K�2��$WϏ|1��be[�b� 7;Jq��(�nòΎ���3B7�˩��ݝ��B��b7	l��uS��[���݃FF������N�.6��u������u��]�!&Uݍ��6M)5��K'.�s���qn�쎗;s�;V,ۚ���U��燹(u��n�e�K��!FP�M�Жk��.�9�mB�n�Gیg�v5n��f�[��a۸���Ʈ;Y0Q���ιz ^��6�1�p�GL�aJ���]C���'Wb]sq6:����c�.�&�f53qS0������[�^^v�F� �نt�K��Xp���)�c����������w��\�7a���F�� @-���mN4��ܛ�:�ˢ.a��6�<d������^�#�[����n��_T�!�ۥ��by�t7=�gP9�/.Lۚ8Kf�A����N��C�V�����Yae{7c�p��q�z0�`Kq.�=�֞dy��;����[�{t�!�61Ƅ8�v�R\ �����}f�6g��x�[�a5�hF�5tp��е���-��]�l�b�e3We����5�fGn���G$�a��@U�!Z��q��A6�̮��чS�+��-�Kq��w1�@�t^:�Ƹ�|����ɢJ��?;�7]l1�Ϸp���ɬ���!�oc��QՎׯa���˷9�].��4�tvNJ�blJr�D����qX[va`���sn9���j�C�Ն�:Q-�"%s�HVw��<�v�{v��n����rb�+���W3m�:��P9k�Z�*ݤ�M5UUUUUUUT��S�UUUCn[j�����Qe�)�z�\7g�.��]X�v���7;m�u��G�K��0���mWZ��[f;M��<��藌������8m��j�sl�ے�"h&��^�U�#�mn�C��IV���Ϗ��x�]��,�3T	�*� �|�PK��ۃ�x�C�.��$����"V��NNM��v[�;�jIH	�VCm'.?��G�r���沒��p���RMQs{֜�Vr$�h�	��R8�#�8Yns�����HG%8N�鶥<�)�H��_lC�����%|���L�@�rp�6qO��ځ")��	Yn��g^[j(�R��mB�|K[�$������{���|�[u|��j� ���y��Jmzw�����G�o-�[g{g��{i��g�������׵�{�������˯���;;Fv��#k:��+�#���Z�m��]�_(���-��C��� b�۩hXș��A0���T��R��a!:>x�kJG�J �����Iunښ[�&w����������p�h�施p��+�HbȺ�qa�<��yýV4N
�AK���-źW��3�.z,�ۭ�k�8��#z!�\e����Z�ZY�M+i�|�Ir�i ���5�d���&�r����f����l:C�*f���b�M���f���30�T��q�Y8�`���-��$s10����KbZnE([�/�븷KV����Xq���ΰg��d�>|�U9�X=�ڹ�6��^�3j+�u�t��;^N�HP�ŝ�okn�k�kx�zCn�+WK�G�۞܉��z��g��&&����[��*�n8��l�v��F�<Ѯ��̚�`ƽ�8�@��5��.���/��i�H���B��$���v9�W"���D�&��yp-�Pt$��sWYh���� ]LM6�`V�]�LԵ�m�6�;�և'!�^�1�s����n�u��ϳ�ᎇq��{r>S��@pV�pAogn����=��6��	ў��S`�+8��1�&�cL��B&���K�	bI{k�Ca�m�=�zꛜf�Tq��tk)v�=��{nD3�\�ܤ5���XA�P3Rͦ�bKڶӰ�([EM��G$��];\D�;p�\=�\�a�p����	�K�l��`.�B쮊�͑.\�[$V��"�B�.���ˌ�\�mͮ��q��Y0`�1���ܫ��ۉk�P�턺�٪����U:cr�ݖ�3sgC3n�\/���s�Gv����{m���*oA%�@H��<�R�R� R�Ж�z��Z� ��b�
P#[oU;Oh�a{F��$�����:؊@���^m������������-1H% ���,<�JL�ʱ�ª�h?'��? 9�r�]��h���Jٛ����n�����r�|A��/���e�f̪��x(�F�?p5�'�e��A�B�!�͡E�dD��e�;պ(� 4����K^��t��% �|�RԊ�8q�u�X���	�T�G�_�
���D�D�C���Q;�eZ�"J"�j�~m�����T<���9L:X�W=��t푧� �&F�ԃ �{�!�i@��
8�K &�QmQ��/��-�F���x]�ab��|Ah��-���j
���QB��V����&/.�\t�v��X�GCL�X?s_vYw����C(���f׫o���vB���.+�IsL )+�� f0(�hQ����V�z=�����7:�Up���4.��H�x�rq�T`���\�d	[��d��˕��F��dG�gS ��(�\���v��� f�m�G`H�pq꿢�����"n�m`!Mϻ�w=~\�,��C?"���0�'^\_�_(�
#�?6�fzt�]��U��E��!|Dј*�.����B!��hP ��@���n��+cQ�9�p�<'l�<~r�cq��@S����y��n�ڪ��F2�`�m���u��"];Sx*�\�%ai���R��;�c�ٽ��H���͓�����A��-ТDڢ.��n��:~�C3�a�}]}9�?2wP�[YCr�{/�6B���@���C_ [TCh^:��O,�|��wx�k�������K��<1T��۞����|���ٺ&Uɒm�D�f)�Z�푧� �L{hQ��[_!y�a�ef )�(�&�B�zW3���ڐ��?�%g	w�;���B�eKk�n��
�5ѣ�����67����Z�kfʕ�!|A�?�R`���|�F��qk�����
�hY\�n����])�$�,�%M��Co&���9�|���A�����Z��Ns#���.n���j�_Tz�f�e��V#�"c4m�;4Y�_3DVoB�vn�xW<Ոx��|[W�-����l0A=ɐj�dQ@�j�Dm�\��ݜ5ge�{��eJ�	��a��� �!*��2󨥘2�	� �T���-r���9������-����<\��:�^�n���ED�\*�Đ��["E/��)������:y��x0n�O�eW8�o�8�(��a�T��,�m|�3[mU�����#���¹�Y�m ��j����o�ן� �ris�`SM��3������ �[�2�P.l���68� ���H0E~"��=^�����ݬ�*Ws{jD�+�gu\F:CZ�sZ��\�9�wz����h��(�f�-�+���4��0�cu�F�J��g ��_<��_0�5O���!K�>g�圣����s��h
��VChP搻����ˇ���}T��t1���[��EJ������y���b�/Hҁ��hQB����].��Aڿ
�3����?ab�u�E~?U1�K�˸\&PrX�.E�ySv\K��O�8��3��-o�>���69���}�#��U:������Y �MЂ!�'<p�Sv3�H��ʹ���8{��6�oE�#�Z;�s�	F�T�5!\�aX����.P\�0F5�[ �2]l������:��n5�ttb� �Ns� fQf4`K2�v���+�^�.X��ں�^�n"���L[1=���x�Fݓ��C�r_�}�������(�]���a�
��Grb�����n#b�@���R�M�_i\6:�p[R��WP��k�3�c����������0<�!�a�(d����Y4T� �D"��SE��+�@�ϫ��@6���O�$��s��!�w�t�#A�L~�`Q�~!�[T���ij� �k����{=�+��h�}��|]����+�C(����0�p�]%^y��3]jر�z�g&������5I���[Q)	�E�����Bi��Z��qUAwe�B	�3�\0`��E�}�L�� ��|j�"�
.�Ugo�窩�<C���FrVV�!ue��Mj�j��)2wǽ�z����/[��V�fq���[Ү��C9�K�¡Uj��L��8ZT���T9��u�-V8ƦA<Eӫ��t����
x���ڵs�=�٭�1Т0�A=ʈ!����n�b�ngKU�+3{�X���4T�� o!e�@�Y��I�6�UvڳV�d(	� �*�`�`V�q=�������Dc&jz�wk:?�5I�~� �B�mv�z�ײ����L[9%;;�p{T�`����|j� �112"�}}�|pO=ğq��T��9�j7���b8A��6�ûk�교�E�A�W���o��Ь������z��ʕ��5(ʗP��zn3:W�V|A��k��`����[ט�7����V�Nq9�j�a�	�LwXh��?�N0�bg�!S�*Y�Һ�ǰz��7�/�.��
d-�bVR��
�<Ȏ�� �'�>�{lW��Y/:�y�;j��Z﫤*��5n�\�0F����h)�1(?�?5��D�7`3�X�y}an����"�?�%nۦzw����HD1�8T>�A|��Y���B�-|�t�~�9���R���n��s��@����`���Q�
��{��������[qڵ�rC�qd\�kۍ����=�}���� _n0�R`�D*]�B���Of��03���͡�2�ͪ��O3��9P���c����=�/vg
��� o! ����;Y��m��@�� 琯�-|�-� �B�������Ŋk��{6�F��'�n��"�U0�R�Q����v�{A�0����@Q%w���LF�hq�A�Gjϩ�ʕ1L�0�T�c��Yy�W��P�ͬ;pu)��^�LS6�Y�]�'I�Z)��Ҙ�����#��E �&AЯ�e#�d^x����X����S��B�&H@���L��u�����,��l()`mDP��%	����bZ���-PC:�Wp_�P'<�hՐ[������9��H���C�L��Ф��[��n��	d"+u�����A��Gol���
�bPdQ�C�8��7:��`��|���hN����G�����]��N��%�&Ho0��_3D"*�L���H>e
��d6�(��������j���v,9��!�~m
-� �B���}T��ؚ0(!}�p]��b6h(��b���[��*��%�Ҽbջ�h�&��k7�̖�|d(��`���ecW�c���.8��녒�^������U��ʹ��*$���$^6Ɇ��M�	rMm��76��ZT@3�y8g��'h �7k��uvƫݤ�X��x�nx����Ϣ��h{�f�-( �5֩ac6��MSPЦv���o@k���줹�&%e ��0��m��a�&���k�8{t�92$��!�tt/(�۵읦���~}���,�O][ۘ���6�~�/�9ݴ���h$�B0س���2S�(�T��z���X�5�P���ݸ7zB ԡG���̀��͡_����O�v��0�q�\!Z���c�ۡ��wXc5��3���ܤ��"S����K`�PKO���ﱅk���گ�!�e��{e�6���� ES�{��gV������d�E^R���2��@����"���C :N;;Ds�'�f,��٤�·C��wXD*�цQ<ZF3�k�4���hcmE��`˰Ъ��03:$5!�v�ogݔ�u5I�MF��O�y�٠�	�5�O_�SD��F�'+ ��W�3�-�#�ǻ�}q��'�/�Oz̖��n,X�����X�]�Z�v�
��s��H���NL��B ��B`��$�J����-8��y
���"��T�l��S����@���jE/�5I�j�{×S��a9��Ȯ��'d�:x�b���(�?6�m`#�N�������0A4B�x�.�ގ�4pD�@�!���ݳ�X;|Aݡ@� �ڠChP!���cڳ}����B��-���QӸ�.��d�A�a�j��6bN�٨j�T�6~��m���C�GF呣�Y�-��d�\K���+�{�}o��d�8���`�T��f����1.����cR9�~i���
#����XA��o��/R�g)3���-�����K�7�
k�[DL�c$�DY"�:Ֆ�i���i�z���W����=6+g�<���*�0$"F���C����/*X�wx�D\@����|�t�>��o�)��.���9*���ڹ�x�0N]���3�=;U�f��� Y[�(���9|����U�T.���� �f����Y��JsRs+E��L\�Nn#X���W]ȉ;;�������fK��I�ӆ��7˲ �F��`�a,�����n���Z5)�x�ec�U�� �6����ռ���Z�>�,��\�pk�[
nW]RKU��5�k{��3-��TN6��u�/��]GI�3�z�OjO���F���ja��/6*`�tͳ*_t�Sfm�ˇ��_K��NpSnaԹS��<�srw5g�k�Ub�`�{WKXR���\�_$ξ�J�ku5T;r@�����Z����[�Q����#,p��ı�,��p�t��SZ�U�$�[7�J᷵��]��;�nUՋ�Ӽ"��%�+9�A)���o^��N��w6��b#0�܏9��s�ڭ�W*��]Sb�t�rK84B��*9:�딕�Wcxڻ���Q�����D �/�����UX�P�����	}Y�6=y9��Z���DZ	Dv�nsܕՇ%�*�b�T�##���(G	���Jd�����|hGWb�WTX(�����:�������vt{�ow��Sn�9���	0�M��"N��K�B�}�����)eHll���Ye�	�\�K1�\��[��+Y����8���skR�-�ȏm^����~Y���˽8��ƒ�(�m�-S��Շh�|�����������۰��v^x3#�׵�WK���\��%�[m��sc`��ҽ��rt���94r���:>dsj�l�n����;m:�J^�!K-�إ!3��g)�����lw\g��_������g{`�=���|�n�����m!�)yj{VFQ�Q=�:����]���,-�$���ˈ�V��޵����(���q������:]gfbskE��9�3��Rw���o��V<�/8.[U�~�:!����V�R};�;�$����
H)�T�) ��ʅ�R�E���$Je;���ZRAa��`p�R��cΰy���h���R֮�) ��fFJH(R�H,0V�]^�w����!�AyTAH)<B�g5d��H(�ƫ��\�� �;H/UP.���h�k���� otZ`@���]�@P�%$7��0��I��8u�^y�밤����n����u�^w��=�<8�XcT8H)
*�Ψ���!I���R
Aa��-����P7�- �����t����`Ba�P��PS�a���֘�2��iHqR�c���H.j��
H))
a��Ɂ��P+�Y���R��
AH9*�C	Ś�z���r��]u}y(�-<��Yߘ���}I���(i%$s��0��I�
H,�2��@P-) ���1$�@otZA�D) �����s���p�� Sr�i ��9�0�X;㚽ߝ����9�C���<aI%!L3���a��P(�,�A`a���/9�s��u�d����$
@�-0�I �U@P���XV�p�Aa�� otZLRAd�S��
�s|��\�5�1�z�7�/7�3�Ă��ZAHy*�Ψ����RAh�� ��B٘�I{��0���,RAIX�%k~w�}l9������z�	 ���� ��n���1�t��<˟f,��I 9A���I ��������]���n��R#�c�s�Wݙ�U�e�����%l��:9��'h�n���M��ۙWG��\\L^k�|<G����DuE���Y)��H%$�$����iB��$��{�[!�WM������[�]Uxk9��;C� �b�X�}�!hM$Z���4�}_k���d�Ԙɝͳ8̨��k���E!�7`�}{�����D
H,�d��$���;�a ��H)�C)��/~��}�y�؟#�O�-�|	�^�oz�f�Vv[��E���u�
Z0�UH)ota ��RAv��������B�02�
5�v�漽�vm ���ˢ
Aa�H.:���8y�5�:��P/4ZAH,�d�L
B�RAaG^\0�Xa� otZK������Ad��H��i �u�- �RAh�@����L7�����
�E�Nz���z/=~M�]h=���|4��<@�?H))
a��-����A���A``i �`]� ����\F otZAH,�9�F��U��z�L�`R�) ��up�Aa�������R� d�]��|Ǟr���y��Aa{���AHUP��pQ
H.�5GR髼@�AH,1�BٶJH(TC]Q���R�$���B�0�H(��XH.���]_R��[ ��B��;g�һ�S���|���~C%:`R$��ÿ*�R
�E�Ѕ$��H��}�ڸ��;
�~x������yY9SP�ro1Õt�<��0��/����t�����щ���L�2D��'�
J # �$\�9v*ґ	J�a+B���U�m�]ml���vs*�>&Q���A�Tؚ�[q(��ie[�\0ѽf3�!�q�`n8�6ǳ�mvCa��geT�����D4��8,�Rxk�f��̬��^�;��Ɂ�։���j�Ú]��~[?S�B�ؤ��[�E�{u��;\GAƽQ�*��z�$�����P5��qD) ���
AH,7���,��P�7�0�X;�5w�w�/�:��!�AyT0����Y���Wn6y�+�l3���e��P(�Va ����Rj�C	����H)�d�uP,II����ߞg9��7�- ��I�
H,�2��@P,�<ϖ��<�y����Ă��A�� �*��H) �7wH)q�oug���~VoRm �c�ZAa�
H/*���RR�\�ZAH(��R
AwUr����?��d|	�ĶW���)9��^qO��o�@��i�$S%:�������ᄂ�P7�-&����L�uP��XouH)��������/4ZAH)��� ��ý�- �1���Aa�[�Uw�s�>^�u�;H/*�) ��*�R
{:��.��W�����i ���r���jT9�C	��7�- �a���@R
Aaf�p�Aa����i=o����tH,�N��,�<�-�󏙺�>H,/t8H):��(�$uP�� S�l�%$)�$�B'�3���Ar�M��l�e�I����fs˫��V��[�4�-&K�}5�-�	=ޅ�-�Y)�z�[&RA@��ل���I�T� ��B���k�u�~gw��^t��@��i ��tW^s�/I�ʨ
AH,0��	 �w�-&����L�uP��Xot�
A@�贃�!I�.��cΫ�NH��Y�n���)Lf�-��̌�*�GKF�Xcx3Z�4gZ�4;+v�>�Q���"�u�\y:�)� m��H)�5P�z2RAB��Ta �w�j�x����<�f�� �� 
J��B�0�H(�Y���R��W^u���<�8AH,3�B���7�-0�I�)�����·��0��I�) �Te;���cV��c|��|��][���5޼8�X^�<$�@gTZAH)�Wp��Xoufc%$(C{�	�RAwT
Myۯ9��ud茤��G9fI��R�d|	Cg�[��sS^�}�@Pd|	Y��N��) ��5�]�ݼ޼��CĂ�l)�xg�{�����MR1�`�ynB����M�fޒ��,x�B��(�����d0��"xp�=��蛀��n6��	�K��7\e�9��X/h1���W��	�O0��L~4B���{z���ς~�o�U���Չ���� !�~�Lܮ�_��3�H�����ͪ�f�<s�5k�!w��hN�K�2�j7�����i|�5I�j�[/��c���&J�6�s���F�'ؤ��4${���x�ٖ�m�s�-Jt��Zu�5�#�=������y�U-��J���i� ���#u�F��}T���5&�����ͿQ�y�ς~E ����\��Q�ؘ"�EA5I�AL?��ju��}���t�^���s�/�l���(���#{*��N�����c~�w늌n�5���5������5e�����6E�}q��nPb���5L3w%����\��O|Dv}K���#H
��i� ��d�OB�+��q�_P0��5�ޣ�emhT��~_��|9N�憂8�A;�D6����`3V2��v�=��<0������[TA,����v#��Wk�j(� ���r� ���;	�f��8+xA�L�����C����^��Q	=�e���C6J�gUc��
MF�ʌ��ˏj���a��=��D����P�W���m}E��m
-��)�pߘG�����g|qs���o�D? [T!�swb����E���j��'	���k�9�
l���Abiub�в�� W/��0����:k_/v�Q|$��gOKE�^�2��k@ �D"�@�РEvL�\���������u����
Ɛ\A�a�EC�5�N�ܟsC��� B�WŵDY�^�ffX����ϻ
��5�Z3�-��Q�%H��d�_O�����0x��]��
.�A���?
,rvE��(0 wW�!�P ��h
�U�ݴxF�ћ�3�!c����CO��m�E~�CJ���3�����q��P�}��죠�fZ��7��-L����	/*��\/0<�����.�,/}�� *�k%��d���(�=:�ݜ��:��r��<Wa�Զxl�x�`|h��b�ͫ���xÎX��I�ũzxT#�.�;q��p��s�3N���![M��-�5�1."Mx�/)���"�n��Q����9X��F�R:f{$@�'Zݎ�m��c[��&骁I���ߞT��N���6M�Ý[��=[ev*����h��E��^�!���0A4B��ou��Zs�ygz�a��b-�_ _��ТD[_@��{l�T4�%�`�y֟ncN�\ �4"u˚�o\u�g��Jj'z���ag�Ղn��v��9�vN�O7���o�#��}��_�Wŵ_��_{)�����`�&$Q@Wlr7����hU��J�7.��2^�G�9��z�"� �j� �T�Q|g�~������ݫ���. �3��J~ �!�$}�׿��u����*f�ka+5J:iuU�A��ĢIr�j��ݠNrAhՐ�<�Ru�����̑�y�/�1p ���?S_6��,�x�º�g�kΛ9��-��9{ΫB��x��
a�ӟpdj�K�J�k��P�U�s�.m�Yv�嬔< �}��9I�8B��r7�����hR�� �K�R�s��n��u}M
#
���|�C 6�M{��ߟ>��ל�w,����\A0B �?���K 6�۾��ԩ�� ��Wܢ��G�3��Ɵ��Q�ޓ�n�mi5}�����e��Z1�R:�ʤP<�mu �
��y����
{�1(
 U/����t��妸+�N�w� ���c!*�G]]GEpO:��%��Y��p
n�K�l�zW�H
 P�`�|:�n+����\DV��鋞�4e��3ɐM�"���5H0A|�n3 F/�^0���藺��cO��k�a�f��W����َ�x����-�ͬY>b���˿�@h�;�74Ъ{��n�����-��a<�5���<�.�~-5�qI�8M��ܒ���xn6|>����3sA��=��օ>`�bP`�K�j���T���F���j�@��d:�dYG�T���o�U�T�%���""����U�Ӽ��t���@�РAk��mY�N�F��ē1�c�1s¨a����$�+��Lm�nƷ�����p`��;pn�-�����\;�\ڀ�c5}߭�{�w|����O2�o���}���[6}C֞�2��U��Xi��u��J�K���k�00�(�܃I�}�����-q�Dg ��F��R���6�m��@���؀��_�[���{~1�^i�ĽܷM��li�ݪ����t(��YT68oZ o��3|�� V>�n�Oa���g��M�����+6�Ǘ2�_M�j����WA�6sʻ�.H�tt�dI��ա���Y��mfAȬu7X�Db�YO�| |#��9I�E��?6���
3��ҫ����>��Օ�Ik�&g0�Rg� ��Ԫ������_+
"
*D5�	��;<�����q����
�A���X'e�r���"��-�F�����
��������Y����u
2��7B�j��4Gt%nl����,��?i����i�;Z!�%R����`*ڈ��W��� �0(�?Tľ��3�j���$���w��k�wCﮬ;ө���;��!���3�²8S{�1�F�t���y@�F�ۨQm ȲB�j�|��g�C�V�=3Od)�У��"�K�<��ަ�I�7�<��}W&�	�)��u�omU�y�K���xjB�4S7N#m�wlBUۆD)ں��u�sp�� �YZu*�]�+�]���ڏ]�`�������%�R�4�Q����y�/,13�Z[cCV�Ûr�wr��G4�]�)μ����X��݋�fәFvU�.��5}p�{�w��=��s�7�����Yb������]����UD&��4��y[�h2HJ�������>�Y��d뷘8>�86�ىǉvIwT�v�C>陵;V�+��k(�k�_{˻B��h��o6LТ���`��ظa=y��
�ϵ�1�Ǻm����i����%�fz� b �=�p��U4�K�
����	�2P}��WV.�Ԥ�%M�x4s�����*�B�u�ַ�+�h�Vj�OI4+�s/v,�P�MરU�yi���Y�yL�]�ܘ���E��E�9���M�7()0��l�S��V��^J����h��w.����G&vi,���SQk
yv��&�ĭa�c�qV��E�K{�^�pD;юr"�C��ͤǤ��ʅ�g7J�Z�Ǆn��A��TwC�}�g�*�T��V/�����G��g"�ķѶb�e	i�F^����[���,���!e��*��!�ؖ^�h1:�f��v_nזG��:��h�ݖw�\�|�ڛGH��j�^�\Cۭ<�5��Q�TS�׷7�{�B����;�Y{[4��m^G���/z��[Q�~w˼�A�:����;"��m|�8�vyVw=����:��X��]�� �ډ8ɖ�dYHRDL�9���]�����㼸���C�+��8�˽�]�y~���h�mݝ6�{X�~��h�ו����#��䈹;̾u��vۭ�w�}�����kQTI��,;�Iȫ������E''yX�O۬����vd��H�v]�P�r�˲��O�u�k*$���mi�QU����I�߷�)o�q��4]�t���U�,X�i�=;�B�ݞO.�[ "k����Ye��X"[�)�tHJe��e�tv5�4cll�9�t�����y�hF񌋺��զ]i�s�� �β��V�u��f���J�i40/նm�fF$��k�A��R�ź�ƣ�kS�lFQ:`��vvUMv��1�s��774�M19ώ�۰�1���	N��xP̊��c�����4 �5k6@�&)oM�۝�3�(��Nʌ����*��m� ��˳C�`䉶f���+��[�^����;��ZIwoGS�x��E��c�˙�>玢٧�ַ��3��7o&��vk6n�ݻ@a���+���Ih[��;[4�E�v���,�蘔�	��|�2ٮs��s���b�a�
��h̅����X���1���Ǝ2I6}�25�l`�v�zhz3���N�^6��^�;XyQ��cK,��jX�I���cbS����sۊ�Yy���<�_b��n@7k^N��c�V��.uf�[!�7mfd4��:�������4�w����f-�cغ�B��=�U��8}$[\9P�����%�]��j��f9����h�6�]�ƞ��<���nv's���`�%ñp�ᛷ��'��+N�K�%I�2K���6.(�@��˜|e���a�2G �\��/Q����k%6ؓU�ty%Ν�����7v2�`��زhC�cF!4ذM�6ҩh��E���Gm����e���г$���:��"��jM���X8�7F<��D�h]��m�\��Q�oiIR����Ep�MR�j���
#�muknC]C��[�����86F�l+��ͮ͠��l��:�f8�s5s�kt5��B�����ŉ�:5ջg�"���Z����'r��Q;b�g���[��X�]��	�͌Lf1�u/�'MWI���Gǁ��Z\�t$8�w���8]��6Ƃ��]:�xw�x�@����e5�Q��Ycl���'�����Ʈ��ݜV��,�I�B�����0<O2MV���� ��Ƚ@Q�BAhXY�Y��iȟ6����2���3H��_l_`,��[B�}#U�߰j�3�x��2{p�0��!|�XdQ� ;ɯ��`� 4�6���D�e��OEG��ۉ�a_��M�AhՐCt?XC�z=;��NYKc�F���Q��0��R�wn���T\ ol<[zKx�� �~:B!�(Я�?5�-�D�������%p�#LBd���U1��̎ڨ��Pl�Ȓ��=i�X��)�����Y�[66�����I����r�5DY	;'�?n:�¯P�t�氼�|��������e�k�wN�f���z�)˽�뼛G�S~�z�Gb�̱��۹&q���+D���D"Ɲ�[[��,�����/G�>��GX|~����6]�{u_MӠZ�	���]3�gWlPM1P�`د����A�����? R`��Sm���x�@�Ƃ��l��� �b ���QG���Y�=5�-X{yOY���ְM��4;�]�Oj�|&%�"b٭|s7;�gb�Jg�[_6� C&�6-�5l��^�ı��n�ɛ�/�!|A�a���4E)g&kw3�����8
ͩT�4&�]c6i���6��	4J�&���� 6��xA�^�]�i��$^W-7!g���`�+��L3T��DL^O!��������K��ɷ�A5�8��/�5HK�r+��Gx�2�,�A>j��ۡ�x-����l�����gF�	��Y�����L׿Y�+1��V(�sd�֏$� ɽ�U�:��9އU�)����5I�AQ@�������ں/��_��g�"�6lk�.���9no�n��j�@?I�n��2Q%|Fb��N��|C<����%Σ��of�}�����AU0�3Ru�'f�ԋ0�	�	��J�Rf?���-�x�-����L!o�㲟�<��K�Tǐ�<�۝93t/�`<�U�3����E�P%�(�sF�YS�7�T �PgE���{c���~�@����A�~��U`�Ǘ��t\w�Z)�H�j�u��&���uA��:�t{r���O��)~d"����G�}��wO�-0FR����z�˽}��*.�%� �G��������ꋛS;�kr�ì��hdI�&[Ǹ�"h�ȇ7����[mV�k����K.���!с����Āoy=n�CѠMj���An��j�;,�����E`���ck�w>�����r�&A�?��~ULv�z"�ox${����s�`���rk���=�������R��_����?)�5I�ƈ_Wth�약�Of�|�7�#�
����&?U0�~_������9#H��ۈ?���{�tݸ�Z�A��s��I���������P!�Vmx=��w �ӧW/^[��4�L��wP�������Σ��xi��"H�A����U�Ү;%oe�ٰ�0LRΪ�<��/��Dk@3��[U��C:5��������a�g�^'��]�|A��@�D����7�����c��{��L`7�ı}���T[��lr�+b+XyTڮ�9910� >}�۾NS����5��V�;�Ùxj�L^��p�ޯ7��v���2��i3)H������O.t%��I�Aj�����r��K��K֜�S���]�7nx#.�ݟX�[=v0�qn:M����3� .����[��Uq�	�Im-Iu�A�:G[�Ss�����ߛ߉4�ЃgG98�v�C�u�GM"Yc��=���{��Q�Ց�
	�^��VJ�#O�zϮ̕��0�,��C5�-֪�M'|��n;k�H1I�H⫳edtb�˗�aW�^!@��@���z���]
� �&5L3������R0�E�7=t�9δ�6���9�?�R`�h�Ct>���2=�,�-|�b�_xO���9ͽda���_p�Q��bH��Р[T%��!�j-�95z� ���VF��{6_L!��?#T�U �n��І%
D3��,�8�v�uѢ��2�>���Q3џ�����x��������-�����q�A5����T@by�wS���o�#��;��㪹�+�����DߟJ��%�WHu��{O���9s�Ry��^����m��`��F6���|>��@�_�#���/�+1~���=Da� �&#5�E���ϬJ�E�@�Y��|��ddS���u��ѽ+���̈́�?�P`�H
j�m
��P�h�R�"���t�zs���6�&���U�G.��,�/��w@�РC? []X}l��[q�� �23����wOQxA�O�k� *�:Z����^�\��v��,�6�u�,qפ���h]c!ۍ�7��� Gj[U� �Bs�߷:���8z��u-�{��v��j�|u����t6A�Do��R;��dqca�'+\p|:̈́�|~����G���{�W����i@��G�Qb3U*:��5O�ˎ4�ŷP<�E3����~���/U���J]!瘝sռ��]�/C�t�����"�VS�NETX�� >��1f��b:�|A;	�sXd2�����X�+֣�@�YB�֙���\u־���a>`��s�6�gu}C] ��[TAn��l7�n#DL@
ᇬ������6\A��|�5I�A�&n`�w:tC$��
#�f���P,����s���%r]�һ�o_l���I�dm|ۯ�Oj͗�^���|���^��|��#v��`�Ct(��Ad"')8h�oM�@��O}~R���=�s�W�񸀠�ȶ����p��Ӥ�Q�@�Q���
���~�샚�y�K�d D�[T~d�ǉ��+j��ڿ�m}�NY[:ץ�ZC����hӈ���v��_��#ED<J*N��M[!�J��ܹ`�44��1'����iڹ�D�]o��*��u�k�@! u�D�Lz��j�3ID��QS^s��:�ad!�1�nW<���^�~7��?6�,�}���}�;.p�W�N�o⬺y\�!��\&���%�<l��_=��QG�9�r�'��K�T�h0�_�QրdY�E�F�����ߗ��_1|�:./���U�:�xN�d���5RY�yč�}:�i0A8B �0��L�����1���|�Vxl��}@�1
 ��mY�D3���О�tk��
 �Q��-"�$�=��	�".���̬ę�vL�������5�-���̗��B�X`���k�MWF�(a�A;���a�E|~5Li��j�ͫ��s�"�6ȭ��O��;��8h�{��`;Z�c1��.�G�^̖�.�.�6P�n�d����� >�|�?�=�g� �,�b�.�❅�֮6v����'�3�Kٰ��ԯSm�;��Q����f�-�sO8_G���u�̌�5��0Z.��ڝl�p6��a�N�j���ڝ�*�.A���	���rY`�r�"�q����BH���Wm�-t(t��H�����:37������連Y[�2��f�Ʒ�,4Zjٶa�p�(���#*W� ��:��RA����l��Y᳤<({���Ճ���1� ��
2�%��n�s��w�U]"����)H��<��3�Ck���
z�|[I���<��0�Gm
�~@�/��c���nV�u�&$�>S��@Ƹ�7XE�S��H���\=���!����Hh�W��O>��:@��	���~5-��"��jX��Y��4�1֪�֬�4�=U����}���U��Y�3�Bk�$A�_0��_
7#\-��{��8nh�{YЏ=��̥����D̲Ԩ����{ׄl�^?U(��T�*�ټx:�:��r�؏Y5���C[���Z��֪�"i�~|�o���ɤ\e�Q� N(O��;#V�P�q"o�Tn
я���rq.:�^�����v,d�E�e��9+i��;�?������z�~=����5��?՛w�K/r<oPY�����+W�Hg���t�?R_T�荋Յv��/���v��ׁ�(g����C(�PX��.���������ڃ�{�0P���Z�����;�<��k��Ad"�Тڞ��=�'!N��_���E����N�Ak�j��9��_uf'�uq�������R644uts;>,�u=����12ٌ2(������ʼ����Z@U�r���2B �0�bdD"*��HH"�b�].�}G�|��a��ͫ̃��l1��㰾c5�E������ӟɯ�\A:B6�mg��F�I��|v��Ix{/�/���t�*�>"/yuc�g��q�4��ҲiL���.rCu������1V���̈��nr����G�Å�E	աP��x1.���6Ӻp���Y�/7��Y�����3���;AF/4Ve�&��gE��1[���dsW�ޕ�nwZJ��n"{�
z�'fX|��ټ�������w��Ou�ء���'7Dfk�<}�nWV�ՠ�v�^&U���ܳ�^��U�˛z]����J�v��ݥԕ}����,דf��'����F]Uބ1NW�h�P�i��7(^�p�{�;47\o6��=W���f^ec�=�za��7�>��fT���k��a���Lemdd֚U����=����p�4iPb�t�J��s�ŷ��z�;���^�}�k%=�<����]tp�;�4����Pv�U5�캕�nv��v5
�T���3���$�w̌��5}�������4��y�^�к��F�|u2�;�Uj��n�kju���:�\�\�mI�R�=շlYsa΢*eu7ECLX��(��<�O����b�7s�����"�CL_h��7-�GF
�6���Y{o+���c�貹odTi�Q���+71[�7�]�]Y�ՠ�9۹��L�{������胼������N.<�"*���:(K�۬��s>yͰ:%�(������۲㸊���GgA���Gol����F�̼�+�:���ymk~�[n��;��۵+;~n�3���8��∋��{:�+̸�m�!GGw�]�򳿋þ7�ݝWά���y���U��e�ؾe�\D۫m���u�����6�����#�!m�]B�����"�������㓯㴸��
;+�*
+����:��mv���˴�)���O��vvt���k�:γ�����gy�Q�ۋ�;�{�qq�`��H��T���U������I��ZW��A�	ҵF���)��@�$�{�}��<��ƫz�b�Z�~k�[TChQ�<���]�TGZ�HP�ʾ����Z\A�DnK�٥�`�ު �x�},X&D(�FIY|������	�f�̞�b>��T>�����bّ��z�w���}�&��Uٷ4vE�hD�8�'�r��qζ�b�s�*��|4� ��dT$B��ew���U�cp��0䩤:�t�;Y�����(��I_T�'�V��C>?3�oljEOs����\/��Qg@���}HCt�t �#O�w1�����U���w�G+�T֝M�]�����@�_eY���_I+���EV,P#uг�Qݗ^�l������~��3�0EB��ŜцJNL�__�����(K��k[��A�̳�Y�1��ļ0I*r\�N�B�r��b��5�$ T�sW�=we�uS{�����CUU􁻰#�mS�^�u�К�$Y�}��,Ⱦ�?wyg����Z04 X5]"j7m
[-�Q�g���;mLnY.뾾~}\�~�$���%
	{L��/�s�tX���=����$������!G�$�,ݦ~�k�b�<�|g��!]Y/�gz�]N�t��@Q��7v�{�mY9e���#�n�&�E����x4�u��IU*��`K]�	� �"_G�i�L!$�,Ip��*vN�bA���8��"�2m�n�Y�cO���U��`��vץ|;��M�`Ȩ�D(�%}"�-��}��T�^�gzfS��6���� ~�#$����KW�lf�L�e�
��\*��*2�v��m0��R�qDU2���Uj|��F�B�c�R��x����iG�D�2g�L�N{E�c�C�m�bX�
Ƕ��l-X����ޞ79���u\A)��<7Y���s�I�{[L�Y�`Q M6pm��R.���л�Cc��˴\SE%�:@Iu�xyR����sb9c�l�TM�޺9}�k��ـ0:xN�F���~����;�
7���z�M�������ݺ���kya��}~�n���/|������� �^?^�u�К�)7�d�k����#�Z� Y���@&��!�<������m
nZ��=W9�p?���K����^�|[b����0�D��� ~�J���b���k{��/gtY_\@z/��U��(�[������� ���Y]�	j�{�W3�kBk� �"	��ñ��1ǵ|�0��X	�
 ��%U�w�[W�$`T����W9�p1g�5����(
��$�������g�&GO���^{:��^���'=&5��L�<;�j���׎<~��#�`Gƭ26B�̕���jcv�9��g�wܧx�����q��__�P�D? d�d!��!�u�ޘ��+0�k���w�n�RW�Ku3r�2��^�9�j��rw"pswl��cL:�  �|�<=���0�3�kCk�&D2�v�r��G^F��ȼ�$��r�"� d�d�wlx�&2��v�˺��Yj|A�5�E��X����"��d5��ZDh#�j�%��_�-���y��K��b�-ꕘ�}�/k�B�����D�/�ڄkH��fذ�-ǹ��]v�6��l��zŃ"�0�Vz���ͺ��������;���m�*ݐK2I��Ty�s>�>}z��ȅ�J�$�@�ͭ�o�M��B��1��F�נ��#��b>7i�A��A�;��3��	�M��y�~N��~�9�`�(�{J���8�(�ڲ$B�������dɂ��]uՕ���b�_(n�����gf2!LS�����r�qlSރ��M�Y1���|>1�q���k�ނ׈?!F�Y�P �a�1�N�z�q|��V$B�uf�/ٓ}��~b�fw���w�D$_I*L��M�{ίʽ��w������m|�	%}$��u{�k-��X�pf��8�%�˱n�fLWvn��'=s��n�n�/v��	%z��n�*^�q�T�w#@;�=@H��"XNAW왵-�_zn�ɫ���i�g�e}���W4���u��o $�$��9_qҳ.�+$�嗝���|����H��z:>���Ϭ]؍Y�j�)]t���!	��D��dNFԹX�+VuK��'��{4K�Ne���u�ީ̷���q̗���rބ%�Q��9 ���d��D�X�� �9���ж��/��wl]��������˅�3Ɨ������sw�b��̯���I3���7s�v�y�(0���&����\uP��e��}C�N�)8}Q�w�j��R���.ggv����{��_wu	$�AGrF�yA� �J7�]4�b�k��.Л�,^�����{���L�eo�d�}�Z��{��7_�,�l��y	J���=��Y΀|���3��ogxVggu?|�/:���k��{���I$� ��rI��6�m<t;8�앭��!λ���m�l��K���SS�����m��&	y����K���R'��W��h�mj�d���Y:�f�d���6�3� �biڐ�5�d�Z�:,f���ϵ�K�u"(:�*��&����or�)Ʈ��9�۠��9���)���D�ֈE�81�mv����e �J[&�!ȡ-����g@qΎ�q�����ɰfc%v�3k����f&����� ��c6�8�ғ4�)5����	����O���V�]�C��B��{�g4�0R�>�!(����U�]��u�NJ�3���%��ɉ�'�7����e��<�bIBE��d[����y��%}�W9vF�#3���J�V�������;�r�]���Wh}wr�鞌���=�U��S�%�| /9�v��_]��a����ݒ/n�n)�=/}�.��I�sڇ�8��V���	�	%}'=�\m����Sk��7�Y��S�<_}�I$5�>G޼~.=w��f]71�4U���kt� ^>S��F0.�U�i3��z2���v����{�y�O��UX��o��I%}"�j�3'bZ��x���ͩ�����7)����ݩ�UC��E��-]�͇���y2*��3ݹ_*﫥��]�� |�j�������7�z�?q˼��e}�R:7&^}��#���耒T�I/�ث�/�n��x5���z���J�K���*v;�_6�W�IE���Wܫ�5�| ��5�K��Wo�"�	�v4+������NĽ=ܯ/<�$RD/�[�ں����^�v�@��B��"]c6�Q�6b�(�CqQ�]!������w���U����vH�)ڰ�cb�(I%�%}�T��.�����(=��z��O���g;�[XL��+_�m	JI���:^PyV�߻z	�������п@�v�K�:HMe�I�v�g"���;.�q�B5�]\�}��ݜ'=]=ڮ^~{�� �W�!���[���r}"��/�k�4��u?|�w�4^����f{k�6K�I_H�����M۔��4�Sz�+OWC�i��]�{��x;��vT!�4 ��,�!\P]�5�23k�iU�WW����L�D����g{�j����R�iZL?-��$�@OR>ݫ�_=BK�~���Ҿ}����,9���u���Xm$���<&�>��vi�g�ɫ�@N�H�)%N]=2���d��������mM;��W/=$��<��9�s#�\�`ꆲQ�]U�EN�!߷�[	�5V�f�Np�4�ȉKB�с�Q,]|wo�Ri����Z�� �g�ݯ�л��C�#tؗ_�s��WϺ���D$���U��Y�/����lPE�(�8j5��u��p�u铲u�D�E}_�=CzK@�u��=�}\�_��rW�6��fn�}��I!�S����򚭹�$s�`=]��n'����f;o���pu�gޒL/�ʽ^���Lnf����2��ug�x�D$��H����w���։��P3�e��Ջ�x]ݻ3Lͫ���oI2E��N@�
ǎ����X^|o���o�<��R/������V����D��}�k4e��b�lܾ�����Wټm��o�XPl�^}}H0�]����١hR8�gY[Gr�ȉ���Dk1+Y8�.[s��B^�#.y��;�>��eL�{װr�Ę�a����j˫��W,���C.ś[t��^<�4�Yf�C��:�d!�]��XH૕�;AКs�,���]�,հ�$
���.�j}�ޮSN����̥fhZ���T,S��C�20�m���n
�⊡<n�Q��܋ƥ	�8E*���6�karD��p�F]��Е�^&&�B��D�]��=8K��P�+K�IrB<�]Ƙ�ޮ�ܩ���#4i�;���.;�#�3��J�Q��)vc/�J��"���*�Czu
so1������\ج�gq�cwC{������̷Nah�$fۑ�S���x/�:�ym�q��;���g��7��r���˭��v�yH�i�̺�݂�ڱ�O2���2����"�T�u1�7]��������y����f�|�6f�:U�&�-���ۣs(L���#�u6w��v�s"�ٱo]��;b�Y�U��NS�Ω��ڱB�>A�"TL�Uf��o9ڜAWLq��"��@N�.�*������wM�]��-ˈ:6��ٛ1�Ʒ�������%5T[)
�Qk{Q��u�w G��qAܖ[n����]�]�rwk��������$�󣲟�$Grw���?��������QE�튂*��$�֖w��w|���E?���O������.���iŗXS�q����ם�=��/{H��;���}��.W�y�Y��w�&e�u�ۯ�R^W� ��ʷ:;�m�I�˷�u�m�7޸���츎/��T�Y���W���B��΅�o>�zuěJ�����h���\Z"�[�5��$��egX����4^xTz�<S�z��on��WJ�F��� F`E�6I����v72z�q�部%�j���(�o�F�l�Zi�.��ɧ����\�3'��c6ټl�m]��6,���}�m�b"±��+�q��,b;{�qeM��h���]�p]�n\��R$Ĩ�V��e@V��We��[�v��-S)�w��]�p�mr��=�K؉�����]]7Oc�[�찍4�Yc0��.�b$l�|�K{g��.K)+�X��8���/V�X6�O<�n7VSk8Ύ�7F��v��1�d68�sv-�:�4.G�������eըM��ZM�taQ���tV�6�jV�#����a�]5b�[؆�]B�fkl��԰���%���fiٱ����䋗�Ü�]� αu�ǵ���ָ�Ȑ���H�B���UŻ�7<<*q��<l�Y��!�+)�Y�[˓AqwF��v�;�wY\E`z7�`c�7e<WK�,��y�3�q�Nݍ�����SN���+2f:�&���k��d�"U�ۭ�S�&���/q.�s�M��뵘w��-a������]����fd1+��g=��Kq�y.�K�9����{ K-�eRX�3���1�ɦ�Ǝ�ErP���suP �60�Mi��aI+���βz��v@�;�^C��l,�c��v�ic�������Z퍄<Q��CH�û�	��B��xm��^8ݫ%�>ݘJ��V�uVj��x׮2f�=�ّ���Q2k��{���|����D����^^�q�jG�böU���)3,��P2�����������^�����&6�
����v;Cے��7[���hЃZ�`�F�GmpqI�*F��b�`�q�9��⥺���wZ��x� ;�au[n�Mu ۷�k�^�������1/���A������<Ѽ�m��З7\5��:e�a�����P����gm	$r�����2��ug��(��� �]Ҥ�Ē���;���ʺ������x]�7�$�v�b��j���$RJ�wɪS{=B���÷���o�G���K�I�ob����'/�z���*��Vx<_Q�}��G]��}$�	�<��ױP��R趮R�7��a���7�d�x�!F7�X��F-�& C.�O�Pf�@���hLgK��(����mX�n���â�P�|��f���S%�|ԡ�{�v���A��	�IB�]�MF�f0�g8�
��25�.�z�5��\�V��'*�#�u��t��pT���y����ۣ�i�P�}����~��Uq��q�ou�
�6Ԓ��"nZ:�l��v��	�G���ݩʛ3ϟq�Nxl��!}y��v�ݶo�Y��
���W�9;�`��y<���yC���WL��wcڀ�&�k��C�:�ꬼ��|����X�6�PxX�������g�<�M�ilU��&�ku�߹���nP7\C��=�o�	�:�R�S~1���<5��n�t�6����m|���-
������7<7Go�s�o��=�7�=h{.n�%
���i��u��g��V=~�.����~�םg{��|ɡ�����{)c܏lj���w��D�uҫN(+�� ��]���IF�����i
�)���fcJ�N�g����'Z�۞>O+Ñ�ڮ�~x���@cM��h�f��My�d��k;������y-��Ψ
�=�b���u�C������V�u��㡉z��gf�U������4���S��^��J�wW�?Y���w�o��m|�[C�����n-���;(��:�D/�*�U���g�:����x��56�_6�yO)���6eyׁ��=8w<��^��i��4-ɔ;�j�ӺXo׮�_�������V����ut+���g��a��i9cg��ė`�x��5�뗭�j���uj�sSq��[{D�V�C�|>��o�RUP*�bߌ�ȝ�;��{{I��3�pjjm ��a�e_d�uD���@����I�b���sM�T���V	Wj�IR�"���ɶ�m6����ݙ-�4|�5'Բ�#y;���m6�{[���=��s���w��𾝵��7=C��c��7��5�_�k��[yO�mDL�|�n3!�u']:���D /m|M���9nsYW��6�o�y��ud���ܥ9��Nߟ&�m|�o��3qj�����g���|����C�����7:;S�ڋ�҈�U���*M���7Y5#��/sB�y�XC�V�v�	�oR��S��c��o��DdiF��� ky6��ixqn0`��0��s^��&�YHddk���m�y�n��mu�F	5�6�6�˦�͠Î�m\�)]�A�y���nJNi�E�u���n-�B;�u���kLJݷ�v�X�ݳ6�yYN��ؓ��{5p�89ָ��1�:�;v��D�5k��>����u�=`s�Q�^c5I�H�JݬMw\��LDǾ�]��
��^F��ڨ��GB��#;u����g/�_6�@�:1�q��olf㿛z���xwVK~���&�dZ70�o�u|A���!������̽ɇ�vn�S\�m|�vit~���3���ky}U���ڗ<���
r��t�fq�su���m������ݾ~`�o�;��|�ܛA�q��t�����c��V�b�vv�j��g�8l�`�XP�����A��ͬ~�6fo���M�����v����ޖ���\4j{���Esy͜D�\�@Ĵ��iVL��;Cnx�1^S�U��h�er}}�#+�� :}R���t>u��]3��<"u]Z�*e�u�开m��7��9p��F�^��Y.{��܃h6݄�G�f�:��hc�>�y��zl�}Oڴ�"�;L���φ�6�mۺ��W��D*�S��}��<����h������>�����h�4;Q�a0cNAݗ,%���.���-u�w���@kn�m��9��Ւ�?!)�����cA�A�j�Z�j̚�=��+���|�|6�����:�r�/�m���y�򔲁�$Z�֜��� ���L-��8�[Ց2� X*A�5�{/xGnAEr�Yvk�BOZ�����u�[��=G����7a�A�s5A>���1d_6���WxwV;�m|R]J��Y���m���#ۭf)�p����kæ��sA��Y�Y�U�nU��(�&�Jl"YMCP�4�E��׋��"۵�5���o�u��RH�Q�r�ODs<������Sd{����=a��7���}�Ǫ����So<ٝ�ú���ͯ����z�����A�Ѝ ���ڱ��|
�g��^n��t�^�T@sM��h6��0�z��ο�hG��Gg�]��r>h`��p+�d����^�F��y̺��Ɠ��8a�:���\�;�Z{,oL솘�r�_]�-�T��� }���}������͖��|qZݙ𹼿q�ɓ��ܛA���ȃ��=���M�����/I���ل���W\&0��D0���V��UHU)���q9�U���Á{؈�i�g�ۑT�m6�B��N_�pБs�}Gg�]߰�>�-h�z_Vt�Ǻ�9�R�/� �v���Ai!���A�3ܻ�^<�m���f��p�s��X��׵�o����+�V��M����A���j/׋;<�FN�w~����1��T�rf��0_dZ깛����U#�`�*v��W9��m��L(lihݵ+�V��������cO�}���\�{���)�9�n�\��X�p]D��F��u2�g����:m�H��l͍ō�J����5�˩g�C��U�rC�U�9�ų�ϷI2(�VqeD�e���vI,%ע��]����W[��q�"waSѶ�d���Z�2�>v�,����$'�j��eo����߻�5F��%�ѤLؼ\�l&�J��G8�Η��&���|�7`6۸����Ǟ<�}�2^�A���m6�mex����r�6b����%+���ի�zv��v���q�/=a�m�9��,�=��Oً���4����JY79�z����a���^����<���nC1RN���:�\�_6����'u{ݑ-m�㻉��Vm��TUقο'������7�܊��qe�kmv�["���>W��ҝ����}x���]G���]tJ�lȭR��
�5۰Bю>L�qs�u��l<�Ӟ�$��Wz��\�ݖ鳣��R����9��@���Е,���F���J����7oj���}+�w��.��32�`軐�M�'9z��=�*K������@sM�a������r7�v��~�]/+��;�}�*�����56�h6ط^��rfU^�+;�=W�ؽǱ�����Ъ���i794wx3	��pb�N

d}�����i���n.�5j�R��w圛C���6��wx��6W���&�*�>�C�}�i�&��w�]�s�u�����g.��:��}4����<F�?3M�����r�zl=�W��s�m�C�aj�C��T�HF��#��(�ӳ���!ڙ����g\���n~�!eA9��y���6�rd�T�NKק٣��mh�xK7�ha��y�],�9;q�*�ve��1��4M�Ͳ2ʷT��2	�%oD��gbu���U_*�w�|�X���2��ƹJ���|(t��v[�*"�H��[���.��{T�A��W�{��s�Z�����.��iR������0��(�)�חr��+�qur�d��Zޕ,�NU��B�j��t���	%_����A�_Eo�k1Ab��Ħ��q:��o3����6�ԥ���ݏ�U׎YE8���������r�D��ko�5?S��s*����N6�8Cښ�1��a��n���nj�]%%N��4�K�m��u����5[��iy{�1���u{��
����djw�	���-�f��lWV�k�t�}Y��n�]� �yS+	�n�8���ʶ^TY���J�,�4�a,2��ܣ���t�t��.��Y�z���7U�5�ۯ��kj�c�2��:r���޴ޞ���r$�ݎ�!�_aݕ �k&#*2DuB7�x��^=Yv�t!�C�r6LNL�ٙ�G����_�������:=�qݞ��Y�6�����-�(C<n�,%-U-�!�vt8�ה^^m�**�{]�zft��Q֝E�^U�q\����:���J�Q�͓^ה��m�����+8��ۺ�+$�6n�.�k�:��Φ�%��vu��h��<�[����n��,ˉ�W���u>��e�ۯ/3o{��rqQM�w�ue���ekn���e�gF`�Ge������f�������|�-��N��.˰Ȣ�d�,O�� �3�����f���m�������O���O�7Shd���w�Y����l\��"���Ś�i�m��}�t���ר﷫�.����>�UUP����R�xW$�IB��Q�uhd5�q�V���eQ�B�7D��`�e��<�m�����f���:tby��OB�an�UU�+������x�ȳ��Z�{�J����ի�i�w��}�2ݯ� ����x_foS*ŵ��a{�޻�y�|,i�mٿv�.v������8���^��T��K���s1��V]�,�
�Sǜ��fܽn�`� �y�پ�e�|�3՘�ِ��2F�.����y�}�ݿ� ��m ��������ܴ���bޝ�1�9����HUU�=Q1��8e.$T��|�Z�;v����o.�!��v��@�r\����g�����#>��{�޹�y�|�2�6����۰A�@l�k�6dk����m^�4�����x��ooj��8;�u�݀�R���\ce������7����+WÚmۿ�﷈r͋`wd�_g��v�u��N��d�2���7�ᖅR�_��ܞ�鼖�Fꗲ���֗i��e�ܛA�;���\��:P)����N�2D�7�kp1�d�5Na��Ι��,Ԏ7�s�ٚR�u�/hϞ���wO^~R��AbS���ˠ�Qc��6u+��{ry�Q�Q�W�x@�IƬvw�v3�y�(>���Fϓ�7`����ݎ�Cb��;;p��z�<q�I�/!�W�`wn�S�n�g�̒k�AvS��0�1Z-�s����J�#<k�	۶�G\�|����uǪn3m�p��MT:������~'�mɨ��ηf5��bb=��-��\�l��'2�_ｋ�|����Q{����sk����0\��������k����n������ݾ���Σ�,��f����E��ɴ_7��>]ٙ���+��k�!������m�GJ��ϧ{��m�ٷ����Κ�-h�{6WJ�7��v��m6�v�����tˠ�o����1�)6�����FM$�V�t-p�2�&����ɮ���K:�����TB��wVE�w\_���:sn�w�SÞu{��{�*1C���:�m6�m}В6L�'$ޫ�zȨ岕�yr{�O�+������L�vF!���!
Dscmp����Kv��z*�{�q�k���s��T_m��`o�+�:��i��{]cTr�v̖wg�k+��<C"m|������u˫Ɖz=�vݿUun�Z��w�ŕv^�v����·��ה���۞w�۝�s�=^�i��~8]U��!d{iP�*o\�Yܙ� j�q�8�n6��eX��o[�߄�__QT�
y��l�5*T�lU�{9�ҽ_۰��A�K7R/�7Oj�O|�v�/�{S|+�{7��Ve�g/�P��oD[p��:�:�U.�;�����כ�Yq�O�'��~s5�\�<�R�t�*��	'��6��fu�'	!�N�w+}��s�=_�WÛvn�4ŧK����kC��/}���>���v�p�6�_6�yjg9,��c���mV��
����x<_{Pm7ݕ�o����Fd״��b��6�M����*z�M�c.������/��_6�k�5ܮ��3����d{��u�V}��`6�lor�8���wp��%gOq�u�{�ڪ�_��S����D_6ݶ�Ι�ˬs�W�zZ�<Cڱ��m���~�[ݔ�j���Ҟ�޼�|�{�H]
��D��äT�V��Sd,ih
�3�[�v.�n�(�����D����0i�N,�;�]~�m�����������IWv�<+ݝ�wSp��Km����}}�c.Lb�5Lb0��:\gno\���n�	���5�oS�9�~g��{��{�ۋm�H��m�m]a���ww��sYْ�tf�d:����H	�*�(��dkLN��A�Mӛ�G�B�^��7������Xm۱#�KN�=3FgK���{ZU�/�ً��"L�>��k��i�SFM&�z9����/��˩�W��������L��ז��zo桜v=��ÇP�;r�R�B�k�٨���;r�v�P�:Jz/E�̫jv�]��4R�e��E��B��H�[G0��n�Me��0̈́jv��7 6�2��V��K�ⲙ��q��ۂ�S�;��t���9��Z�1Y����&�l��p��hB&�!�6&ji���4�R;-=CEj��t�w\�s��M�дR�zZً��z���Kۦݯd�5P�Q�������]���R@�.���A���y<�ʫ�E�8��r�;��|�K�T�S�����0�䞖LF�;���g-�i�>mV��*/�����:��4��;o��f!�A�����g;�O�ͦ�o�hf���	؝w�r�s�褐9��ͷ{)e7�s;�������'��w�{��4]��Gز��Y˵6�m�n�����޿����+w�b���~{Sk�ܼ�������/�����v�6�L�){H�tk���K1�-��S]ӟn/�����ѭ�V��\�z��Ug�yk�Y�yF�h6��M��B��e
��7-��:I˵F�Tߙ�]
g��I��w���/4ࣗwJ��C�0uE<���\꽷UlO�:�=k�V��/�I<��m���J�UR0"����7P�a�{��(7��R���X��;�w��	��h6�so��[��{�k=᭮���\�{��'�t�7o|9cA��i��m�m �'��[ғ��);�=�R�n�T�ǐ�1�G��~�t�`�0��g���ԫz�/C+�ͫ��,�K��ח���h7����^ÝֹN�]Χ��{=��_6�^�!�8�ֳ��yoOd���k�o;�\~�����@6�n�l��{/,Оu�I�<0:������f��T�)�|)�f��G�y�k�v�=��	���k�@�c�u"4�q/c������Ow���D��T��U&�����TG����m��>�����[�(	L�ĕ��wX�@U*��R�R�Zr�~���.��K�z���F�i�۫��cW9�
���
@,�Ӵ�E�u1 ܦ��,3�l8h�b.+e}ت�Kl�m5ѽ�(�3�{7�nI���l������=:!dF���Tԩ�ۊ���ze�ߝeb������b�j��k�ܺ�g5�]�c^[��.���b�m �c^��;s���؀�B��N�Q�9���J)����O����\A��R"�����"g5+*7Ȋ�uvf{Wso
�n�+1�n��Oϯk�� N{�Ÿ��B��>�0�������=:s1B�b]���1|=��������va6�yr��wV:z7M��Q�^���c��#-m`&���o�z'�݀���_�~����Cr�o�={����6ݏ�Cf/��It�>CY�����s���hdM�>�̩Wٿs� ��ܻ�c��+|��O���wb]���f!�M�m�^bQ���hgi�_�C]��V�h�7�N�|�h6�M�����ffm��^��\<&N��f����ν�s��ꄤ-2]�f�n�D��;`q�ڕ���Oz�-��;+(�m0��o,ǀ���D�����ڮ
��U^vB~�96��a�ov��B�3Z��eLB��Xwd�h��/O�&
B�(v
B�k;�z�[��b��ܥ��K[Ђ��Mgr{Zu��WV�jYM�.`�Ы��!|u>�Ӹ$=qY�j��dq�h1�NQ�l�c�̫�2�_j�h��O2�]vQ���lx�ۢ�we��t�;4Pe���6c5mL�E��n�M��$�Z�w��˱R��w&8��*6�N�:�Ҝ�qT�C.��FtY�XS���6�a����L=�t"�*w�u��y�u��YP%�wh;��Jw0C����Tr���t슎雨���h�gy�{NIa�j��)��A¸�T�Tt�tƾ ��վ®�����3j�0��n�}�&	jh_vыW1���ڔ���;�<=.��u�wHr�h:0���1n�5x����݁�F�_Ұ�Y5�e�[�Ȏ����zi�-�9��y]�<nIͬX�2��v����t� �vD6�kvpnr5�=�s��Vf���i������	�2���Y�f]j;՝����ҟc�[ۯ�P�v6\l=�&���=3.=Sn����%]^m��ڛ�r�
��+2�!/+$c��$z���"���B�*9�� ��6�˯{Qtw^v��#�3���W����"�������6쐸��F���Y�[t]���{��u�ͺ"��;�-;�aA�dی��:˰����|�û}���$�݇zi%��蛵s�I��^�u�V��t��;ڼ�����v�k���N�=+���ί+��U��e�[����L�9��|��8�$�iH����q�g%�vkn9�[v����+:�V�oX�/����z��#eպ���g\ylh^���&'���&G����+��Kof���c��R�p�fל�l�m��ͪ-a�au:#�:|Bq�vxΪ���v�ힵё��T�Z��f�#t��;�N�gjX�á��-vͧ����UyY|V	��8��Z��q��Vxڳ�"q�u���.,W	]uXR��:�nz}��8i�N���<��]{t���m2�]���"C*˳G
ƑI�]2�k�o.��5]q ct\ Q�ef���۴\���9�ݍ������!�[u�$Z�ݙ�z�y��rp۴㛵ǆ��%a��Y�)2�Ɗ��܁���	��¾4���Z;R��ɺwGV\����N�N:���j�r�V�H����Ƴu��%�b^��΁���1�]8�sG����wۦI^N�����胚�F.��=[v|q��\=ڠ���^�9�7^%��.�仵����I<`k4Km��4iWb[#*鴦��嘂������R�Mx�i0�qԚ2�.Ћ���k=vܼ/`�)�$yx�m��thu���L��{������h֍�YD�t�Ձ�Z@#����H�7W��#B
��:f8ݙ�7��f7f��k�h0]]>��7�u��:�l�s�J����Q�Ķ���4���\�[g 9�q��I����3YU{9��B2�^7A����f���v�n\�&�LM�-A��f
l`Kqf����,����a�vY��O XU�ntv1<�h�G����4�eێg�Ѻgp�a��t�����KUZi���d�2�	]��M32�h��y�!�YcO M��/4���PS]�J��l	P�&6�.Y7���������\m)�Y[l��E����]Xͨ��F���ə��)vS�[�����E��dp��h�w]�u�Cn=���n5e~��yrS��6Ӎm�l�C!�ȃ"����[Zgm�J�~}��� 4���J0�u]ɥrVZ
K�
L&L`6�6I�Q�:v����3�3�8�w#_}�!��Ne����UUT����3{:l�R�o�	�3�E�����lW��&��7/6�����m����Y^�`���ڧ���1�^,��m�����u]R�fn�mfc;���Q��2�O#��%��Sm�����K&�t�b��_>�bk�1w��mT�����z�dV0؀�5�[0D���.�
1��'��S��a6�Y!n����UER�9����2vw�lu���~S����{�l�)ب���D�3x���C�Lf^�A=5�**����.���{�w�g�#,��Չy�ʞ�"{�#�슱������D��^�>�]���G}�U�m�p�]hNA�M�uJg��w��������V�|�n�^.�:�Uv}-�Z־m|<��k�K��d�>��A�ή�b�{[gw�9��6�i�2�w��[�
d���;2�M��}2��B���DW�/߹�4�1�� �R�m��]ku��ˍ[<��2��?�V��m���Ǟ.��.�^�����}�v�m ����CA�:�ἔ��#C��o�j�3�3����S}�/��)��~�w���ͯ�C�'��pOX��1�����N�ơ
�.#�t�þ�w�u��=���Y�0w-�kP�]�ѹ숿}�,d��2����o����
�[����oe���<]�b]z��Z5:�a���υ����a�ڧ3E%�6 :;�4ם�	�S�8�J�7����\aB�C���([����z�k����̅&�`Bj!�h�B�U!T��A�7�k+�]�{���ԃg*򶇼���m|����lJ48�[��9���[�8lb�74�Ū��sW�����M�����^�I�z�s��:�h�g�p��K辶�۫ߞ�����|�a�v{Oo���u��Ǣ���oʆ{2$�1��=Zd���v���sNK�Ni�����S�z��S��d:ԣ�����>_�zXm|A�����V��J�=	�����u���hsn�od�9��[�ed�����Z2��S�ŝζ+�G3
b�b�l�]���xO^ϯ���o��q�ֳ���WcDh�>z�q6�m|�VEd�!��bDb��{������w�����1ɇ^�5j�M�7�:�`���Y���|���htA�i�vUz�ދ=�Z��{�>�z��:��^�#Չg���F���ͦη�<�O��<C0U��ή���w��9U *�pZ�ޡG6�L�θ�O���9��r�Si߾��|�Q���unB���nR��l+�t��y�zE�~��9 ��oO�aR��M~�\k�V�ԷCHl5�e�����4�p�q�wM�E2H�8�)��ZQ���ECOh��;��`]��t3`�qrs[1�g��lz�V��bJ��wc�ݠ}�{ku�#��『��V�[,�ieр$��+���X��flv�Qu�k�ɺj�y�����}��sv���v�v�/3vZ���ݶ��D(����ӫ�>�SفPܕ�O|�7\���"Kދڛn�mxɓ�M�P6�ѧ7����O�'8W����p �{{r����c�ت��'P��_f�q�)���;W�K�Ub7;�}Qs=�w�n?h�ا�����U�[ԻJY�撙�*�©}T�Q�y��v{0�=�Σ�8S�PW&Wv��to%�����1j-��̜�/f��s�������d=@.ӂ~�5m*�UP}vԸ΢����:�#�<�r��_6�q����Z��W��I���{h��ݮR�\r���&��'\�Ș�@�A�:#K�}��O�v���+�9j�}�6�WQ��jP�]ɶ�6�W�9��i�{�i�x�|*��M��m�r�yR���Z�q��aHY��X꧂�q�OwL��L�2��T�^cq�b��*�h�7����&��]��6�����Ǩw#B����j� d�^��l��u���-d�B��p�B�F���'�R�u�볮��к�5��r�r�h6�m ��^[��:׶�z���v[������9
�_���-��Cq=M�7�E^-!R����6���Ä�W�:�䉛tì�4ni*&Y� ���~���镽�d]����q���X��:r�7�G�����<�Z��۪�M��f����r�;����~�9�*�ٓ�
b���Ս|���ِ���� ʵ�}�:g�l�\��[�D��Pm߹���_r�1��.V�n��:����,��tO�ӱT-�Z�Wu�g;�ڏ�6���+^k��a���8���wUERH_ǘ�֯�>�琞_n��λ��sQ�Z�M�;�o�p��'!ھm��C񰼍�Ɵ�m̙�O�/��h�id��ҳ.�*}v����=�n��Z�Z}z)gT`]������V�p��b�`ԉ5���d��)�3M�3c�KP)�X��
�l�8pEXꑕ2'�}���D���m�� �3vO9U��ί�'9��¬���S��ڣ�5��0��'[�����2t�s��MDB"m�~��B�ߺo"�
�*�fw�Ϸ&\����Mz�Uu����vޗ���Lą�9��ѷ���+�z�Zr��No9��6 M��.6aJA�H�űn*�i�p3���l6�UC&�R������|O���W�nJ���x[B��f��/Y�SBjm�_6�n��^m�V���[�{|+�ux]��D�Ô��7��~ѻ~����~�J�YԮ.}5#�#�T1uc*�M�@�y��!�"����`�D?���n���;>$m�Ֆ��R�=�ptgYfp�@�7��g�4t������g�A�E&�.9:��t�n��2nJl[�α�g�e��ob��ң�8�-�ۄ�-�{j.N���-X�i��fA�������Z��ά��IE�=�vݳU���:�����Ɩ�8��Bƍ�&v�_6�O�s�?.��̃��-&���8��<S[���#�@�d�1��r*����Q��g�������7G�U��_g�h6��]����)��n��/;�o�s�>��y��Fr����_�Sh6�gz�{c�V;x��xA���:���kM��{D0�m.;�N��=د�3���_
�Z^2ψ�7;�-�/�M��ĉ�����;hEV���7�F����RI6������$3pI0�P\5g�\����f�dZ�0���(��Tjy
�W^wC4vp[����l를�=�����m|�����ŗ�����A��j*z�jd�us�.�^���t�\m���s��sL����yC��hG˔�z�����Q�7�1u�ң�3��Ƈ�®��Vn��_������#v�������raћ�d��/[����ɶ�7z�n+�8��^ug8vpY7��B.����W�dn�_6�������v?<J���
��*ܶ�c4�5��x�*�ј9���p��Kֽs�r����S%�����	��m7��~3��s�_{�P�tyr�^~�#A����W�ugpP��i�[�8<���D/��V�mwf2�S�:W�K����,���=��M�8:B��J��D��Ԏ���w�ݻ5lU�.F���".ЭOr%��gv��
-C�I��KW\�k���B�\q��[��uJ�M�tw>�:��+��˛	n��	XM�]1[��P��IF��Q�ך����;$� �`R�������<Wu�jx*�q�Ki��hWl܆���X�Ų�u�e^��=��;��������2���͆L ���Swƹ2�}���@ic��C�v���w�W�������c��nܢ�,u�0=��8:�:ȷa���W��ܻv���Z�^\�n����o�:B��T��;�v	sz�ˢo��(������ȯr��+Gz�jڳ�٨d��PL�Y��\i��.��t5jʾ�,�ee��6���[$�%�n���J8�7��)	rmc�j�w/+���0;[Gx�jPm�d	����,b�n�m��!�i#y�V\Ζ��}��Q�n��P�U�
�nؙ6WEzT[I
g��;U_u��F��Ҭ�uʬ�U���[w��vFwn�{����FS�뵸j�f�[[�V����SuyMވw�-��2�ǭX��V�ޜ�Pc�8ȕ�Ic���Bݝ�:�v_i�i�uK("�1�huS5�/2�[�tl��qΜ���Ȳ��n�ar�Y�~I}�Gd��Q�K��kZ��\Q�n!�6�ֲ�Yh�{���ww������V=����W��#L,��_-����{n�;B���^��mM�+�ݽ�̾[ֲ����g�y��Ze�e��vvڳ���[��&��ّ�������YM���+�n͸�lێ����&v����M��l�ٵo�zֶ����Έ��hwm�+2���n�mnD��i���6��@���l��V�۬��<Ž�zؽ����(*�%9��<	&��7N;�w�����!�Z�_U/���S ۾�I��nr�����N�����}7l�y7ȃk��m|��j�j�u�=F�!��['W��_���v2��!�O��h�r��&�1��z�h74�~q�_�)�-�ڱ?���u*��WV=
'ӛ%Ƴي��3��4/�M����_�ՊW�rp}��Dᗲx_g�רE�q��̓�W>�����h~��f��'�0l��kc���i�v_6�v)'A_
�vkk#B��͎��Y�""��j)�L>q��w��봱�k��۪�i添���ń�E���h�&Y�����eѩ�(̪���٠DdZ��� }�zW�g��6�m6=כ�r���No}���z�G�Y�Z;7���{@O��e� ������;\�I�`p��N�U�.�iw/@�-h6�m��[��Æ��պ�ɓ�Uk�֤_6�A��{���{kCg����޿a��^�_oo77�^�G��؄��6��f�[U���{d±�ο|3P~M��m+���������Z�{��sc��A�2�4f>|�m�k������U��οnf���
��i��7^g�*�A��.+�yU^۾��/Q2\��x�72^��6$�Z�VYp��Z�A=巵��їw����e��~!�_�2���]2�]@���٬	�E���ς�6;'�;�5�Fѩݢ��n��p�8+U;F6��;]U�*�&ڶ��7�1�q�nyz48�Z��==�e��mk\B1���Z�21��A�2VЫ��v��g���[����8�3�26i,���5��;�P�~߷�}��Xq�t���:�I;:�^+���p����5��R�n�uu���/�Lo�;z^���:|�K��ͮ�%�]�����uV�>�+����v��o�_�qfV�/�!�6�A������C�`U����7�k�h��M�d�y�}��:R���}������	��姯����m��M��m�/og���Rv���ޏ���UK調�0{�DCj���p��Gv*1���σ]UgN�Q,�F��n�Fסּؾ�A��ƾs���7��/���%�c%�d@kM��ͯ���S��4���B�g����!������s�ݼ�E�q�]�M������c~��I�j�:'"h�EG���U������g����ׇ���z�xA�_1~]�:%��_RF�z�wl3v��v���XodKSJ��qj�۞���LGc�_���v��zB ��F��mO���6�'���1���0LJ�{�X�bʈ/�QUdTA�JOh�Iy{�����;+�_a7��z�:�}㶘 ߘf�3�ک���xrx�О`;��l�9Nutk�]�6�h��Q���Wos{���	�l0n���wږ�x�yFmσ�1����b��)��V�����O���2�=1k6Ή3I��m_�x7��A�����������z�7]�
=�4_ :�0~;��n�d]��7lv1�n�^~6]�}<o���󓭪� U&�����Bs�Y�����t�q݋P���آ)2e�-슻�rCM��U��Y��F���y���K��_?�ԐM�d]�����+����C~w�g�?�"튾�S���zsn8tx0@3)�D���l�k�(�}Bz��aȨ~����#�؜�3^��F�g�07���N��u��1(0 ^?�Ԃ.Й�ڇ�{޸��Ǝ�4�-Z��[\�#�p��q����5���C�i2���?����q�ؼ�^�zy}�Ș�zr9Y�?��g�Ȼln�dl_<�*���#ˇ�;i�c��T�<O��6߇G�`����A�wǬ��R��|·�yI���.��k��Vj>h����h7}7�����J�/�k�,��wx�k�w>_G���H����6�;��ν������?��U-�����c[���x9����20ML���Lg��p+0ƭ��|��л݇w`���bH��U�޼2&'k�W��� �؟�]���A�A�]����S.L+'Xy��Ks��'ٶ�:<��L���H��(%�I2��fa��"�@�$�[����1�I�0*h~���xk�lv]�6n~og��_�,�_�`ݯ��O������=�ډ���:{�d�<\�r�`ݦ�A�E�]�G�͉�ލ���=����͸��v9[���^�����ڽ��Gѫ�`�����}T���4�<=v��;�oã���q��_]�&�0Eqf��+iIh3����;ݞ�:���"��1H0B�g֌A�y�$�h3v�h2.�u�G����a��o'������G/|A�0A��$n��n{�展R�7>��֭bм(d���$�;c�K��/Dh��.����
AOoo5ennt���=�UBfr[�a�7�fr�]Z�uhljG�b�\�K���f+l7\�4[.�m`��q����
���;�s�v8|e#�;P�]i�nur�
�ݣ�����)��޷����y�?�.���l\��=���m��QY+�S�Щر�o[[��w�{���+l�ݦ������74��6�I�:�j���oS����~r�3
&o]6�x�r��{F��\;�Q	�T�u ���ڐAl1^��x/	�m��:�B��6�_��X���n��ݦF��_r>�P�|�h ������oݾ�"���׃��n�z�Ir+u�!�s ݰ�"�|��ck�+5��0�wLl��aم�����񚾞_8��"�$��1u����ψ7lW�E*��7�ã���dgdo8�E��}Cv����!FE�Nw��f}�Vz47��gb��O��r���� ݱ�Z냞�[u��ķ9�B"��8��J��nˎ&�������_�����v��Vd�ϻ��磗���Bּ֬~�a��� �n�"�����0���c�O���m�բ�����3&�'#l����4�k�:u�"��SSfgkT��W�y�����vj�r�`^�2/�?�ߴR��^���^xį��a�w[T_���^��&�i�E�ݦA7h�q˒��������s�&-X��v�b�w?15��f�/�5��/�)������1������s"3�N��z=����	�&E����[�~���B~�.���k�G�̦Fj�~v��K�'���O�?l&��f��rṣ`�K6���H��fm �E��W��Ԙ ���ڒ	�N�ޢ����Q��(@��\(�kuՎz������_6����ee1>#�U|ow��G���e�{�xNb��0��q����q�y}~BMZ����O��lf>��x�����t�؏JOldv9Ril;w�����w1y��&+��4W]����2�IƵ��������`����A�.��7k�ӛ"kY�V��0A�զ/;���������9��nPd���15�r�Grv� ��`]���ʚ�r�-��c�z���^�t� ~�O����O�뵣z[⽽;FYD��b  �X�i�X��\�h��c
W���Kp��Dh�x?��`z���7l<��n��O��m�=�`�ʦ}���b��l2=��$���k�m�o��}ܾϏr���?O��Ncw�J�ܠ[�v�F�?z���|Ey�	�� ��ܿ��aGA�w_G�]�R�1���+��o��O��3��d]��Ȏ���.�C� {�� ݰ�nmý�S�ۏ�`���ɋ��G��A�c�s��FE��s��X*8��rnfA,���\$�Ͳ��G(�=OS%@���jX���m/�y�n�?]���ݫ��WY��iT���������a��C�Z����R"����U.���!6�	#	*<r��Q�]��ma�n���DC%#	z#�w�u2��.��E��ޏ?d�z������P�)�N���, �|�92��0E[����}^W��F����"��Fí��;���fS�~��}_w!��2=��E���ݬf��q�}1���{�
<��@e�&�0�A�v�����c-R�GS\�wlS��/_���\��>^��o���2�d��}�"����|{�"�n�]���^�����;N�\�۫�Yૼwn8=C�̯�����lP��꿽��@(Z�i3X�o��/օC�l[Yz[Y�#�v�n�9f�;s//N�t���Z�j�K��$p�z�[�#�m`�l�{[U����&�l��vb��}�l[���3���+.,��ԧt<v�vUk���>#I��;-����ck��8t}�1c��e	Ъ;�6٩�38�h';,��S�m�����d�Wmۗr���;��d=p��2t���Z�f�YŇ+�)n�=m����v��`0�hVZ}��w���ʳ�q���q$WL�}�_^n�:�雗��^��+�A�!�%�:v,�s�K#J�e;\��J=o1���-D#y�i[2���B��hu}1u83*1dϰY�n���.�γ�8�u�V�b��\LS���[4ZS�NE����$D`͆�CY�j�=*We�V����V�g���ddGg]rZ=�
�em�pD+g7A̓�ok{�c���u���vX��Q�y�t��7{�����,���-�䝉�*޼�X^��ʪ����Ur�.���Z�����}A�.����W�j�]��]J=U"n���Xl�&��Cf4�Κ�������B�{������0��r�c�Զ�����{���[�t��'}Is��y��i��(��7)��"�p]���(���u@�-�ͯ�_i�3�2�&-�P��ʜr6(Kou�F�/qz��P^,��6�eiR跽�O<�; m��{����.���;k=����{[j��H^ݗ��u�_��m)�������%X��3��A)��;�[F:&k'�ޢ�{"qÜ﵃�-�����[8�h'� f\tNR�\�'!պ3�o���"X�̢eh�����۞�
�i��ZJ���mDu�d�+@��-<�����Ͷ�6���f�D(D\"�������;#6��F�"��Zy��.��[,�� ,G�w��׭4�v�W�;#�t��;Hj��f�#P�&^mRT�^)��ɃJ1���4�l��.˺j3�κ�e.;Ȗ�6C�.y����gv�M��A�8$��`�R�\	���\a�>�+�.[����8s7��n.dVGc��h�U@K��
������`�Q��DZBϣ4
�%��:���`:��7q���Sw I��n���2���\��W-k.� Օ�ۙ���=���4���4�sm��s�o$k<��:M��W�pq�q�W��3M��9��䗊v��C��C���s����;���7�V�J�v�҆-��Vq^�oC2
v:�K�]�"��#� y�vvv�7d.27�n���ۭ��.nL�6bA���\�k��J�&1շ<��L>� ���RF�����nc��v�X��U==�u���F�&o+jX#-M�F棴�������l��<K�>eH��gV�u�@��,[v� �Z�P�D�A��'�쁱��=��Iv��u���I=n!�p#�c�͛ 
\��-l\puִc��:��<��\̒ۮX�X�{M��;XͦB�1pD����/��6B�����n��m�
%�[�t� 9�6�X����J����B�7vK	e�H�B2�si�L<j5˃E)�u�^�c�P�������љ4��H�:�l`2�����Zb�f�ÍqCR`%�$e�݈�{NSWn9�!��nɦ��N+�I!���l���N��-r];�g^%��[��0�y�㌝Ec5ST�Z���*:ɜY�!��1θ�s�.O]<Z��6��f���RSl��
�����Z��>��瞺���k�Z�F�V4Սŋ=G8�4�Q�dtq��<��oh��`��ۖ�b=O7Qtlr�V���G��	s��1c6�HM&5�ie�ؘH����5f��.h��>c)�F�Fv�s{gFf�7���'�� �iV�ZX���%TZh��|��=��q�pl�����,�=ϯ�7פ�?]�����#������Q���uOr�ս^@d!'��"�E�`���*�O�V�bc0	�^ �/:����3����Az�<��u�͂�կ�C�	hH7k�.؉���{��)����x�* ��E�}%}"�7i�a������LM�b�z�#����kw�G���"�:��b�A�L��s���7i��l2.ڎ4Fw�7���jm�F�=&#w<�x�Z`�/�`ݦ~�V�M�7���ῇ$~o��X
�Z7n�Z<�H�w]FcR.��D��(x�����_1v�y�®�O�7n8ly�Ǔ��M�RA����~�a�v��j�De��ԧ��}|�����-��<.]�u���^[�:Nug;X�=}{�U��.���w];��*���W&�֕~��&A�;��؏u/_���`�bPdv�7j��f�)"D(�@�g¾�
����_��^DxFmg�/A�_;��_0n��h/E�\^l޼@H�a���"�=ћ
��>�ݸ�z���L�R+�7�#\xO[�?�kݯ���2.�`ݬ��O�gg݊'�ݑ�^��;�
P�3(0A�n� ��
:zro�SU%�F�7 �[#���ݜIO)�Kh�M��
��PC|=8�u2��.�?�Ы�[G��1�sk;�x��㽭p-dK��
/ʾ �"�$�ȅ|�%�W�o��>�`����=ӛ�ʺ<7n|���#uE�����㗿p�0��O�5�Ȼ_]�.��׮<aU���I57�H�Xm�K
b8���sRR�ۚ6���;VF�)�P�$x�.o���;��o^#U��˴Z��K�?�+�"���
IT5����m?��������]�-�(�L����>^��6�c$oi��dh�}��A�/���A�A�]�`�����_N��w�ǆ�߃�0L�`�3Xv�wl!��<_Ͽ^�nfն�&W4�6���y�A��q��uvE�"3�w�����A���&�1y��~���w�W��G��;}#���{gq2�l0E���v�2��pN�#�|����-��ޙ�9�|�x�f� �|�7iq�Ԭ`1���$����7i�A�`�~�����Y�[|���L�3Xd]���ݯ�l"��7���'�����p���6�w�&%�����9;�ř�qBr6�݃YB�ڡV.�ھ�k�L��Q��}�a���)kQb1(U�2h�`,�k8��_1^a�v�7k��blVLF!���Xb�p��~�F-�����I�؃7k�n׻M����~cT���Q�xS�&��M�=ds�+�z���4X�_G!�:�f�2��'cѝ�1����FAHq�.j�` �0Ȭ_?���2*7�P�<��{�=��Z������M�"�ڙ�W�&7���,?�� ��k�v�w���^��{ev��bگ>^4���"�AE_$Aw��ʬ��9�(�/��a��N�t�Z�����RdG}]q���<���"�	�W�H��ݩ�v�[��V��Ƨ�=�m��S��bP`����c(E��(8�a᫑�3��٭13Z�8EVe]�s�L;�Ϻ�Xӵs!��H�͝ˊb��R5ec��(e&��0Od�"�{b ���}a;�A����͕Sp���1j9�gh6X�8w[���<�y�y�qZ�''T�q]�/+v��n{%�%Ǝ	M�:谽1�4�$��um�v=����&�k�g��!���w=1�=Q��z�`�;Қ��Z�7�����<��qֱ��wO]+r����X,D�!#�_�`�����.�?�п<���L�1mW>^b���ѩ.�iG���m3����~`�v�#��yh/����&#�c�#c�s�O�n��R�o Ȼ��)�ҸF�gg�|��L��ݠ.��Fx{=_R��k5�{�x0LJ�v�7i�v�]�*bT�z����Z�@]���{8=~��G�cڏ>^��4�Q}�L�QX4֦A1}w,n�.��iV�yڏw�+j�7g=K��pZ��Z~�`]��툯jZq��hե�
��P
��&e�A��;�>|�ǉ୹�J!�~�\A;i�?Zݧ�ݯ_a�?��W�=�Ў0�K̞�����5ɐn�d]���L�Շ���Qk;kz�����|�x��41��d}b%=++I��JU��/o��Z"Lvi���j�U�l/ھ{�^<����[�|�x�f�{`ݣ75��3=����ʟ� � � ]���E���dN���J2�*}��af��1i�܅$���B��|��ηִ{�W��A�ݦ:�a�{�����&-��o��3�w����
"E����~��o޼a�G�X��^ȷ����G��L�ڸ�����b��&�1Ṋ���C��� ݥ��!�@���LDh����@:��LE�v��ޝ��ʌ��z�z{�m_�65��
"m
��+��EDG�q\x�أ��R2�ڽ�^�^����@;�7h�~������\�'y2.�k�R&5���<�)L����l��,%z��j�y:t�n'��)�A<��)�9�]T�wm]�\�Zk��Zu�l��xZ��coN�[�~|���'� �X�ڒ.��ۓnM�C�?�Z`nد{egVx��Fnp{�	�O�7:��z}q�O��~�0��`��O��l?����s0�=�bbk/�{�k£w�W� Š�h3v�wlv���{R5}��do֠���G4umuq˷!sL]��8"!A�d�ΦA�9�E����1�x�"�����eF_�2�}��E��C���?I�hW���a��r��B~��5����1�᰾v�#���l��7����0gW���a�v� ��������.�'��g��?|��A�E[����a�W�}�/�ݲ���_��/�G{��)�?>^�R`�������+���͵sR5�(��8`������d뺭�aM���Md5���ȋ�<fL��Ju��Vf<�? ^������dB��}"��[�� ȱ0�WV�����1�ᰇ��L�;�r��B+ڳ|z�A�h���q��-��y��&;y�1=Bcx7)ת3����}����8����3��y}��[�>v�<)�1j�ʍ���s�W0�9����.��v��{qGj�|F���z�c�#g���{Qϗ� �/���X]�cƾ2��7WۈIB��W����0w��s?n��2n�#v�>�`����a�.����2ңY<+Ū>"u}������xgF߬��nxS�Ġ���dLǯ��{�m�v��BAc���+�����0�g���wd�ڏ>^f��<��3�ځ��o2��%�v�Ы++�2�{�AZ��l��e7����/�g2�vD^����)F�$�F�ɨ%����c(�c7e���5��m��J�])���X[&%�By�k����("TB�u�m�u�oulF�����RiGb�s�U�)�Z��C�����[���==t�-+��,漸��5!lj<]ea�+O�VM<S�F�"�)�\$���lG���;k����T�{� 8���ji���{i�]b�]5�B4��q�q�#�R�9փ7k����i���y�w</�-uG\x��)"�F[�7i�7i�,{ӕ�/�A�L�kgw��]z�z��^bPd���k�Ƽ��t&pZ@wO������n�c_�}�*d@��>�d�ڏ>^��<��2	�L.��]������a�y2.пg}y�ɨ�����L�����O�x�|G����a�����|��f�g��ߦ���H5Ɏ���ݪ�7>��&%?]����ݹgt��O=z>��M@���-
Ռ�2��ZrՖ��������?�8�����Hz���z�NTk<��ę{�z��E0�;��A7i�v� ݠ�Z'��F�s#��d�E
������X��u�j�.�Ѽo~ٚ��qy=u��4�w�zw����vF��%���u���ژ ����_�9y���1��k���Ix��f[����?�?IB��W��N�`X/Y������.Ueڭ���A��a����E�a@~휮wy|��3`���a�ٕAF��_�N�����Ȍ�ޅ}��.�q��~�L���ݠ�"��>��
����B��c�7|����|��J����]��c$����;�e�.�O�(Ma%�s���a��ஔY�Ǟ����]-.����ߟ��r�`�v���{1uW���nx)�����ͫA��G��D0$B��d]:��gpHk�w7�bٕB��k�'j��}��dg��j&�}��%=w��P �B��
2/�B�����f/��~x)�E�珹�ܢ�LA%�k2.|&���]]W��j��9s!,�ei7u��拘q�p>�r�v��k���*	n�E-u�E����O&�v�Q���~+�P�ȭ4��G[
ܳ�t7��|FKT�ڦ�7:�(3}k�ȫ1���f������b7u:�������\s���Փ:,d3�]�s��f�n�nt��ǂ�WW.��Əji�e7�wһ5���򝻗�έ�%�Y��tEb�뒫9_d�:��V#�NAZr�(��j_sͣ"x����A��>�[����D&s3Voh[�\WW7&�����t�nr}�횾����s�cت�X��
�1�8ގ�7s��Yv��3݌9�-l�e��U[��k��P�r��^�f�Y՜xC�E���K{�۴%m���۝|�c`���&Z��Ŋ���].X+��I��=o{l��v�[�g�r,nH�[��'\���Nm�zŘ�W�ǂ�裳cw�fhOz�gm�Z���N��0��a[�Ǭs}]u�I��UVqS;j㬳K�����,�{�ꙃSSvT�WCr���������V�D��kc����^�t���`�Z��[���|������B�����I���[�9�i���'`D�N���e���wmm�6�޲��'[-��&	��$���G:���o�d�[s͛m�t�/c�$R���ЈND� ��#[�����.��f��mp~i�����"I9$_�;���`��JR��)�z��N��{����9����|N�������Ylb�[zmY�~��ه
~h�ᘎ������U�3m�PDG�~����8Y��qN\綧�$���S�۸p��gz�lw���{Z��p|�$�� ��B�؄E٦n���ʄ}���ﶿ4r��sn���JEe���8�ӤG�m����:'�Y�tskm�H�e{�vs�P	 �b1UAw�tgX�]�m�{��3�B�/�C�P#yfC|E�B���a���ݧ{���=�w��|��HL��1�Ϟ� ���n��"�va�8*��f�����h�w�xxd�מ/�g�ݧ�v�$��=�R-�8���`�nv�m&�8�4i��J)�LDp��	� �W0��_]�y�3�3|�s��y�����T9�?��?����n��������k>��>�W��fODz�_�焴<bPdm���~츴~yy����>���$_P���]h��^��1�4Fl�<^��~��3����@aτ�YM!`����R"�����F��m9���x��^ N�a�k���W�x��_��-�����;�B��Y�tudv��ܽZ�nJ����\`���;g��U����v��v����8���ϺYW��؏
�������@?���������L����z�v�{e�5���g7�1&,ɣ�� ���\�X>����Ծ`f�Ȼa�n�c/*�l�w�Lf�y��ݴ���JA�c��I�Ȼl�����>�<x��
�|��0+��=�/2�7<9���0A�2.�g�U��ٿ-A�j��TD�P2* �nץ��	^�d��G�������bP�I�_1v�"�7^�����v�du���v����ٞ{��^x��^ �׉U�������_3�L.����A�7o봳�]����y�3/z4{�ENnxs��nW�v��"���E���F�A�n�bXW�α�Z��v���ٛvpb}-S��)�Ř5.���u�Q���i#�����F	���(8M1" �`��AQ�ƭ�F�;p��灆�,�n��;L�i��cf�.���e�� �X��I6wQ�3��]��*<��lnR�%m:�l��6s�7'G�XW���zMh��⇂W
q�oirq��h�Ѩ�v�M��f{v:K��!���pjk��޽�=���-�6���Ѱ��s;k�]2���٢� �b=R�~�_1�]��ݧy����	����V�fyZ�^�����2���7i�=9��{v�ތ#%���l1Y�Cby��n�z1x�W�_�f�n8��^����}Ծ�C�7l3v�"��wZ���o�Yzv���AS����7)�;P/�J��բ�_*����������<&��s��0LJ���te8��Q�(QP�A�QI@H:�=
���a�]P��}�;�^�^���7��_0n����j��ԑI4�|�+'W���q���4.�KG0��ss�������/��g�7զ"틾՞��$�78.��F��wqՄ��?��a���ݦY�{���M�9�^���ӣk���NS�=�r�rbl�"I�SW�rd�����3G�i��Z��{�빎�	������Jw�Q�J��U�E����+��$�_#]�qB�R�>q��Pتy�%n�z1xL��ߘ����"�3yx�=S�HX �"Xg12.�b�ڳ�|{�)���`�r���Pw�]�T���0���2P�"��z{Ќ�ww9�q�Ǆ��m�+_8C����v� ݱ~�~>o�?��=�B��n]��Cf�C������=p��;>(CF���Rփ"�|����G��}�	[�^�_T��}�1W�)_��=�3z�ݧ�m��A��qe�塃\��u����<�.�J3s�w��)�G��$n�S����,��r�D�P2*?H������u�C���ocXlb���l��[;����v�,]73_}0P�Bݘ8���N�G]��9�!��ٻ�0���a�}*<Ᏼ��+_8C�n���dv��v�c�S��Ư8��d���v�ц�}��kroы���de�JQJ� �C���b�5k�`��k�|�{��Ǽ���{˞w�y�����0A�L���]��?]���y�p���& ��A
 e�Z۲YX� iF���
xxG�A��J8f#c� �\����?��i�����>�Ż�����j�}�r�| IB�U}"�5엾�b���<�c��)�*�3��&�&��A3��~�0��Ls�Vx���1ÌZd~�+���|A�J�QIB��'��v/%;���Q�~�����"�РdT�ףoe��F�\_P2*��ݱS�>�[�
���@��EA��pW���H3n�v��f����S!��y�Mg����Sd�W)��]/+R�iK=�t�}�J��������?�~���6bD�g[�J��9��n�oы��gS ߟ�jH&�nU���_w_��lro�Fнu��$�w�Z�{p�g��v��Ճ6W�(�a��ȻB��gy�W;|x1����V���Dy�������L�v��s�;�{�Uþ>��?��;�ݱS�J���^`�� ��7ja{��	�m
9T	�U�JD�ꑊ���6m�ħ�k٭:پ�^���7�7k�n�"�%׬UĿq���=������v�����y��W;~��9+�[����v]�����O�	�Ln�f�*<��u�5I�����;�W��������3Xf�|����_�
�s%%삌���L��9ǧ~X��D�*em�vZ����n�G(eZ�'*�q���.i��% �DS�]F׳�K2�@u�rI�4cLuՏ.5�Υ`BG��{]Yc��:��:g1,����q�ۤ���k{nK�S]f���[pa��4viy�q�<�8z]�l��H��)�Ԙ��=ʃ������2��W]HYbM7U��u�k�s
����&j*�+~�]���~n�\O;V波���{C!�-[ X)���_���_g��E����)d�v�ބ�f�1}k�zyn[TE��Z� �v�����G���5����p�2���ë����y�s�����J`{X`��]����H0cS ���]��ԐMڪ�L{��^��:���F�^�bPFkݯ��a�v�>�g�бz�b����/��a��+wU{ޔ�&����_ћq�`1w]�� �^�"J��B�I_H�p^�y��Dszϭ��w����k���"��a:������~�����L7����<���u�� [��ZW|����,�>����2ݦA�1y�{�c_z�dn�*�S�u1��B�������`�y9����S%y/F�Z���j6�s��\O���u����!6r�؈�e�̂�ZJqM;�Y�oc#/n8x���>���^�U�zS���b�������n��������2&��փ�7i�nخ�	,��W�~��\m�s��?v�.��v�7k庆���:r��~�U���n��{�s��c#w��0LJ�1Ց�贄?-jd�a�D�P2* �B�"HS^i�>�B���+݋��5�~�^ ����_]���v�m�\������-2 �១B	�F�n4ݡX��;�톡���
#�m�3�2���L�.�U�x�ܼ�߇?|��G�09����
��ݿ���A7i��g���;�3��`�&/7��1��;�
��1(z�Dv��+�B�#e}@��!��+����,S�xֲ�~�:��5^5��F'������9b�M�b��ʶ�{��5aa�QVwj2�얜ki��z��5�r~�_����
2/�Ȩ��K3�HU��h2;���QJi�x�ڼ��~��rSyt׆��륂H�o�7�`���i�n��i������(�*��z�3�^���R�� ��7i�E�������"�)�D8�'lI]y��$96�B=��A�m�/u&K��ן|�/��������7l:��}~�{Y7���:Ƭ����(Q�T Ȩ�+�ȅ%�F�������Y�Lwu~5����+����	�_?�X`���=٫����%xO��b�n�j�'˛����L{&�dN�4<JZ��RE�v��ܾ�iiy�Y??�Э�^ط�g�ܹ��^ ���"��o�7%�8mI^O�Z��kǵ��)���u]�ndPӽ�w��7�GK�X�2��5YB]t�p�;��}�ҰA��]�7h0A�a��}wq{am�W�+�{��j��s��&A�0E�v��q��1ú�E���h�9y�ie)?��gʹa.�n�7��B	�_zАn���v����tv��dN�
~c��ׂ��Td�� ��dv��BM�`���KG���/�vì���O��7noы�M���0���tܽ{����P. $C��!�����^��֫oß���}�2.����L��p��W�x�@�?���7i��z�>��~���A�sv�Y[V+�9�;��{�Ď�V#7�,M�P�:z��Ϩy�e϶=�(̊�k� �Z�D;��Z�]j��>�����*|(��UW�Q$��	mO�I$$~?�*w	$$y1G苩�Q���n�:(Ɵ�ك����H0! B��ٍ��1��F� HH��F窞��}n!�RW(?y=�P�B@'�$_D6���{�׳^8x�{�w?J�s���𑗊�b��k��z�:�k��߸*G%��37��o�I! �!��~=�c��G���>D �?�jH�	����XT�}���q���'�t�钏��������ϡ����8G��$�:��~U�.}_c'�%�ӢXC?)b�t�_��{R��?qY����
������Ϣ���O�>w>�D�_�I�?�E�I	 �yx�;������2�Jd! !�HB���Y  Hw*�w�Qegֶ�W��ɰ�������x}�B@'��i!__H{�}�Ǥ���	�Pg�S�`=�c���$��~S�i(����ۿ�k�����(�HH��*r�r{�󇮾P�������,ъ?z{5������쯧��k��g�\��&@���OgA�=o�����?�=��HH�O�����E���=3���X��!G5�gƉ�	 1��I	 ��hD���a�QMI�c���:6d(!�~�G�XH@&�G��F$��r��@�#�z�BHFL�L�Oy�I�ϲ��:�i*	��39��Q��-�T;ٜ����I	 ����}���'�I! ��}�8�}����a��П���q��8{����{�a���LT���>��'���>��?�=�����6���T$��	�I�ϴ�>�U$�������I! ��2�cԳ�?H~�~��?��{!�=�,�����63D�
?��-�W��&|��;��c?_�������uf�|q�_�z�HH�>'��w��7�_,�B}�
������'�g����P~�d���=��@'�ē�"{`O{�O��ɿ��Ԁ@'Ğ��l�c�A��tML�:�'C;��ϝ�MC�E	���>�=!<�M����"�(H=�Tǀ