BZh91AY&SYgU�܁_�`q���"� ����b"     �                                    TI`} �����   �                 
          P   f�=
�"�%(�RU
EU*�����AE(TR��QI%T�(���J�UB��QPR�H|   6EI ��ATJ�Ϡ�6�Pw7DE]��U*wgc�%Ϊ����9:�R�*�T*;�D(�ݹDP�gW�
PQ@(7� ���.}%W��H�_F<�t.ڔ��<�ު[klIe�o.Q)*�$�ld x�� =�UU� m������y 9� �  G��  �I!T*H�H�����(� 3c�� {��S <�{ ���Q\ ^�)�0��=�:<�{ ������y�<�^� ( _  `>@=)��zS�䐥������ �� n���'��`=��|�T� �|����`=���� ��   <� ��JB���
��$�0*�� �= ���v ;�T�p �h � r;� 9��S�1��p   | ��C ��+� �q� �1u�9�w*�� c�s�;�����  �  {�)"�RB��PH�J@�� �@��9�tg`��I!`l wX�� q���K�S��@�x   |  ����;��ડ�!�P��Rs � �%� �� ��7` -�O
  �>   �
��Q* P�UQEE =��s�;��àG "8�7`r С� r�W a�v�   <   >���<�F�u)J8 d r f�$2 wDE0kP j���� x     >� �� �)Q�!� �&LЊ~	���P �    z5RLJ��`     LA��T�%* �    I꒑	(� �1  B�IP4���=G�=#C4�����>����/����A�7�#�y��l6g�<-��ι��PEx�o�E�TO� E���PEp��������'��O��OU?� E��r��i� �+�0x��PA^{?��~?��ŕT�L(��dE7`U?T�T@���UN @Q���L���0*�`�L���AM2�:`4�Ȣi�T�*	�M0&�M2&�L)��(r��a0&�CL���
i�:a�i�4����L	��(i�4�r�e0��CL�� i�4�`2��Ni�4Țe2�,	��"i�4��#�D�i�4Ț`M2L���4Ⱥd2.�WL��U�/L��A��� �"�q�L��
i�tº`0�0:`2�̃�P� �t�:d0��:e2��SL���4�:gfP�(�4�:dM0��L��GSL��D�i�4�e��i�4��eCL	�D�"i�vWL���i�4Ț`N�CL���*i�4�:dM0&�L���0�Ț`M0��L��� i�4��ɦ@� l�a2��L��D�i�� �"i�4����SL�T�i��L���i�f@�(r�:aM2��Sf�*i�{d0��4Ȟ2:d�فtʺe]0��.��dL i�;dCL��_v@� �*i��
��PGL�*:et�� � L
� �M2�L�aAt� �T� )�EL�&�@M0�a4�"i�D�Ƞi��*�TC�x?�2|��q�ך<�7��r�ݙl.gḦҡ�X�jxj�J�᫜�m�!1�ݹI&	0Uۗ��wX�3GM������߻S��
��^ސ�#��3��9���&�=���;5j��a�f͸�c���'��@M��r�N|��1������R�,SYǱ��ۉ&�gsK���r���Z�C�������g���)�Q��z��o]@�s��N�h�J#	�@�������P7�Mh��	&k�g1�i���i�}����:�Ɏ�"֋њ󰫆����j�f=�Źe1�vbZ�t�ˣ��[�l�@L�G�'�K0��N�m/w�Q�fJͲv��+�2
�1��~�25!���j�zj�_Za��H�
bDU٩ҁ�;��4s���-7!�e�X�;�\VΆRSjk_.�un]=�ڦ�u�gYʙ�<�IϨiY~۝�S"���*�x躦+�ʇZ�ڳ�����M�`C�AݷK��`����+����:�	�q\��MֶRYݰgw'$G-�ʨ����;��üB��%�-�1b�6���
�ֵ�:�#�ƌ���;�/��́��Q�秾
=G�e�a�VU��!��śs�ͼ�Ą�h;�ͻ�f��ac��j[�=<4=ݷ�����8��G
ԧV���nW �#De�jw���4)��j����jzY�kܗN0/A�ݐ�\ppn��Y
J���ѐQr��8qP�+t���-%���D����S��f�C9nM1q�vnj��z�2c�HPM��1|��M�o2�6k�? �u����]6�M���1NʩY0��G�C/1�ע� D�0L�b��hu���7���XG�$|��xr��աp�n�X��j�s����)��J[��ncF��JT[�����u'ױ3�X�z �P�yq�3�`�h���.v�h�2EormZk�OO^����\�ء�t�%�<c��.=!�i�ݐ^��db�ߩ��d��Z �&�5��|(o��w���ݯ9ь.rMM����.M�8�L�<���&����X�ȁ�ݫ�>�A�7_mS�x4|_$N�v8�����#��o�n��a=R�fLu�ib��Ӳ;��L�^�p�u}�����N�j�ݎ��`�n(��s�YQ��@�F��PwH�"�Dk�xm�Y��no.���2w|ۄ���g��7ި�&r��͸9�ӨLw��C�$wI'r�os�����Hw�P�/	;�x�W\�+S���p �`d&�P�[���(�N�5V+-��ѸB�=#y�ܒ#��[�*�����JA<�SG����[ݡ�ui�4�ā�h1�U��3iK�\�Z�f��q4o'���쩁���x�����[��2�W������Ў�-�\R�pn#C{c�q��ri�׺f�����f��b��Fu��b(CjZ��.�.��r��ɴ�LCa9�wwb�>H>�!ݹ4�;�.^�ˇ�歕5�_>��t±����mT��P�p�,ņ��t����-�u[)IZbX����gip�C.�(����23��� $G��l*V�� N����$tވiKy�͓,=��I�����zE�@�%����8�򳴾X���J�^Q�����h��K^�x=!�T�v�־��IĦ����y� �t��z��<r��=X�����lWq�^�ghy��9aQ���-�R,��Z�Ҕ���F���׋���h��hkud��&Ԑru�C������ea��,��]ε������:w����1WͶv��({8�h��sn�ٛ��\� r�F�ۏr�8D[��j��P�<���+�M��pg:�bMe����}��4\���[�GW�%���ܰ��1�\d��y���ٝ;S��e��vH5;�;��ŦY��)��4N�VQik:-HG�h]�=q�ӹ���r#H�y�6�coi�3�|̃/1�v��Og����8�WPѸup^M��?��47`'�j��I&αn��\�>�3rvD�̥��� 6}�5��6��TZz}Eװ����+NY�L۫�5��7�{�R�<v��j�W^�:�;Nm-���O`o����ol�)��u7�9�Ȁ�W��u���@*�(��罗�@�j��S3�I���V����ֆ˹*�l�,���K�Yd�6�ϩ���MLn%�~D�k&���"�#�͗]�f���u�뫩[ݒ��yh<V�s��2|w���w!��v�Aїgf�.\C8u��e���ϖҦ�De0�Ȇ����zu�YO*�2�$j���+��E��g��!�9��w�����۞߽.�{�i��쉍�šxĖך�uA����Dww<��_
R�[779�>EP ��ۢ��4`F�I�3����3FL�� &6#u�ý9[�P�pAڱd�'��C%��;^�Gn1طc�����p�� �f�ՀBn�k���õ2O^��w5l.I�R\�D̈�cD��,��d�n$>ƛu9p4{l�Yƙ���x�s�a���.��P��Ѹ�md� ��WC��n��J;���M=�PH�g>ۇWK����wS	b�B͑N{���������u��幷���̑�˹���˰�q; �f��ze�f:������l���Y����X���>{��^Q�sf϶�݋NR:��y:�i%>��G}˷ M�8ę��2���"���V��˗<�:�g�n��z�t�*^0nO���0�CskGs�y���Yvs�̲����&乲w'�	��s�Zf�	�M��EqÐC �3v�,,W>-p��N:�ɔ�9��Y��ݎ���L�aޙâ��V��,e�-.�������M�K�Yza�E�}�u��;�`1A����pw��7zV�!�p�}kR��K#�(�p�c�5e ���`f��ܥ,#A]B�f�L9&�Z4�7�.n�R�岼h���\����d��V! ����II��G�nIx��wJUa�a
�^�4m�[CNsK���}j͕�h�gA�vNc�H1L:�f������
ۻb´��l�G�}�>�1��f��of��7�P�fÜ����,�dͧ�9`�Ժcn�,cv�x3����Dԭ���6o�v����ݲ��ݒ1yu��|{g���������'�h��~���.�g�nA�Z�"�o+y�r�طh�[�{��Nǰ�#��{���oQm\�p؝�x��iW/�O9�f{�����s}�@g�ǚ��9��iYhk
��\#���U������[�F�e��wht���s�F��%z�0�J�=<4�uYPYjsF��G���z(�{u�P���8Nzļ��6e��凲r����&�p��͊��ĺ����oW.���fkv��uR�i����]�{��ʎ|Ƀ���,f���q!��J�c�:	;)[�x%��ߘ
�Mߨ�m'h״w��{�q��T�G�AU���cJ���mK4��3�;j¢�3�:o"�k�bw�IK�ŷ���;�d8
�Y��vp�u����+�+��Y�����$�F�j�!�۴E�M��g^ʝ�̕d���c͘��������1oaU��
���.2����P�D]��˻����ݯ�<���;G+N*{���]�������nM��n,Rf�;��v�uY͚;��`�IwXi�rb���v�/5����t�Vmv)o$����#�[�f	�,�G��9��sr\B�"������ѝ�*��S��F��Mq������D�g�;�h����[�|��gc�w���7���a�Ф�Ǎ���T���槒�Sb�i�C5$kDlLy����&�m� �ƙi�I�ÒO-�&՚��VvƩ�;��3���8&��7��ݧv���e��H��q"�;��2c�l���3Q��p-�-�վ�#A��ګ=Q�78�k��F���B��#k��w;�pη��N\"�A��zz��S�uʕcur|A �����//kG-H�ޫ}��\-����P�q:W�U��%ˍE��tn]x�s��l|Lcv�Z�a]{��v�/L]e��2��u�a�r��ƀ�����t�K9�w�s�9a���h�L>�*]F�61�e_��4L��$"����~�����s�r/5J����]���3^ֱ(#3;5�������^ɦ��	�sO�>O�e L?G]8�*QN��[��ު��MfkM��;�f��9�KH<x�$��y��-7�Dy�:�_j:��L�إ�tf�m���L<av���G��{r�Q&�/���]�E7w��Zֵ� ���Ʃ����H|��{��1ݘ��s$�T������h����o��"ĴD�p��p.��s_=�:78*ˑYĭ���^�~�"g��gʦ�X� }W���,h��3fL��B���	�V�t��D�{�iS���}�Z;��R��c�f�]W/lަA�tnW�Č\hո�.C�篚໢�������ui�R=(U��G
WM�^Cz|�t[ʜǈ��ԶUݫ�wf�ۂ^K������,�v�nv[�ƴ���*
��:v������ü�R;,��L�$�Œm��;w7�����P<�'.|�l��!�
&.+6��>}E��˛���[|���ܗ =z%f�!�\��^3ˏ,p���I��J�5E�w�Ș���v�u���=N����wN�����V�d}`���΍��_�u�,Q�J:�v=`���/5^Ն�&2"������ܽ�I��J�C{w������.�=�[F���a�*�{��)��\8���9�Tâ|�I�4a�p�z�k�F9b�;;x��9�]!D�>�W��I3sw"0��)���7[ �;g��"��^�qf�^�vwLx9�{�eX���֋�+�K��s!�;��cm���:U���C�<���M� �w6��y)%tQ3� G+i��p`�ˣ�ʥ�S�X���}U�wsN,�yhˌ}�\���Ý���z�L,]�1�wq������L����Ҟ�ڭ���{j�����]ÃN��;��!�!�r�uL��U��xd�����m��M�����_�f�[��r���V%X�Ď�7s�X�Z� ���k@D�Z���J��3�ͥ\N�-�V��qVu%�O]�n�8+�3k���ޑ��1�'k��q�������y�t:Br�z���Tk���ٚ{y<�w\IJ��8hY����;-�5�ZЀ^��u�)��k{�DwNȒ�F<���;����=;�v�g����N�x$�&nh�g#;P�ݿS�&�;��&g&�
s�qZm��;Q|�� 3�ld�^�o^��Fe�u�[�f����s����7:��D����;c=Z�ch�~]e���cAaqǍs�����0L���B����77A���ܳ\[Ǚ�&��{G<�����K}�������Me��^kD܂�c39J�D$��Jރ�3�{@�X�U��s/~�v�bM\�X�?kE��h#�C�N��v;�E�;6<Cwb�Y�8R�Jk���y����1�kz��.�pnW�e�P�8���]h{*��xAG��s�O�tt�:�II㸷��e�&��)���n���(B(��+�+ ޳�.�Hy,̵��&c�Ӻ�.h�;qm'��x� ��=Ԗ��4r���6��L�wfC�E��NۋN���>`X�Z{�,2���*B�l�;5�{���*�I�f��&k4r�-ں�H X]�{nَ��A�>�E�Ɗ��5���ӈY3t�"ep������~2a%���UXp}��wt�Y�=%���ѽ6�5l'�)��t��;3{2�f_�#m�gvh!��Y��8;�.o�y�W���;�Zѐu��]z��^��󺂩�Ȳ�)KQ�޶.d��<��-n�'h�ځ��s
*���"m+ya��.dv���a9�H}t��W�'c8|����74�".ǚ��s���s���:�@)�m�{An]��(� �S�m��������7뽬a�N��_H��T�>ǽ�w,�lX� ���x�.�z���.	�0-��;`�P7��ay�*x�zb�q.=��1���T��Awx�g3̱
f�Z�@���R���D��P�A/g<�
p��!ڈŪh����@.�| Ǒ��[��^����E��2�����'�5����:C��H�{�:���8�C���N2��t%�ovU���E1Oc����
;6ͥ��¯weg��`m��w�Y8}<>�^�,c�(K��n漢�<�����"�)���l��ZM��t�G�L�����=�����Q8D�v{���%���iN`u����K�J���b��4a�f��x{{�
w�Ȼ|Y>���ʲ����(�ni=SUe��J�r�)٘�iz���r��$��yŢ7�A?�	�d��1�g&1C��oj�N����-4��v�}K��,"ݥi��wt��!;���ްFZa1�1��Zl�؝�m*�OH֗�P�`�l�@$�$���QN[z�����KZ��?q6C<l\�������x��U�a�)�\�(v�/�!�BR��)��C��t.[?�:?=��:��O_H�����~S�#��T�P2EZi�T�
C%@)P(22%W!�%D�C!2@ � 2!EJTF��$iL��T���J�Z6�mQ��*��l�(- 
�(�B R�4� �JP�B�*�H	B�B+��R �H�B�+B"���eJ� )BP�*P+@��*�H���B�(Ј�*��@�J-����J�4��*� 4� ���BR��4"�
�H� �*���"�(d ��*Ђ��4� %
U�o�C3�Ô
v�@��:�y|
̵�K���]N<<.���Cβ��e[��-K[	���B�9ė5�����!��W��@���#+|�v�Q�ع��w��y�R�Ӕ`դ?��>�q$Cʼ�;��:�)�Ld�fe��BSK��݀p�Vo�M�������}�°�04���$5��Z�p��WK(�jZj�G���6{��t�;��������Cwr��|��o���:��i�( �����/������?K�?[��K�Zl+;Ϫ��Q���"WJ� ���Y�uѸ�t��w �lBnR� WF��՝��Y�d�}��t�|�ĝ3��U�Vެ>�Y�z��G*�  �wd`�Ǿ9�3D�G���*P{sY� <;=���Xj���e��n!٨�������庇��0w���أ����i[�O{D}Q ��"g�����n��P��_lL����j�?g�ݧg��}�X�����+5�m#uOk���{
hՓ�Z��zFӼ�y8�5�ŕ�[\ӷ��޽��o7Gg��c<��;ۯ]�{�.��{9?�d�D�zq���;?;���<x4p���=�i�=ܻ�KI��VO��/-^ނ�$�_wc�	��{�}�珍��7��=��wR�Af�#�Dd�����t|����r'��u{Ɂ��8%�A��D�k(��q�������j=
tA�G���xꛋ\�^�a���n�4�Kv��@��>�С'`�v���Wv�-��w�a1��B�hi�5�-�2��|�A��!ʋ��zNY	�~yĹ���O[Oy��<�LM!��rv]�8�WX�m7��sG8�;��K(��N�B���+яf��q����+���_���w�o7o���3��1ۡ����R{GZ���7/��a�쨀D�-�ᘼ� ���ٶwv�F�y�K��ntB-�t����vɣ٧��ic�R�u��]QF<LY�g67$���/z��а��ﵾ���ҸF�<\��k��z_}�K)�~Z�&A="�/oW�G��gv�H��+�n��(����{�T՚�WY�J�]�Gʁ{�+� �y�Z��=��z�^�BQlg���2��ƬYo��!�Ŋ�I�^�&�c���
�X��6́��y�-���B9��ja�*�i��Y���۪�-#���߄���g�'�].u~e�k��|r�5d���f�<�xgy���r���o?j=�*��Hs��W	�;NY|��� �{�=�z9q��'~m�h�{��F]���)�4��9��l���x����O����o����n�/���g��D9��Y�#O�J���.��.���V��wfėu�#��W��y����� Ys^��汤v����;���Jc�E���0�?j��/���9 +f�E�'�����\D�����y���e�{~�wY*z7����I�}�/h1���м���Vk"W�=�xMㅶ�ީ�{_sݝ��v�۱�l�FA�� 4�����
�{ݐ
o��?Z��������
�t�W��)#�G<:{(�!�������w#�ۇ�k��d�l�7˲�v�yc��GԢ��Y��r _R�n����XA�b��7.{����};g2A,��/���5�$R��t̓�q}|�:�u󃟇{������n�ǻ잓�o�ћ����u���o��~�o�oK�|��v�ү
��۾\#�~�d����x��i��`�b5��T#���
����$ɼb�+�Q컓��"���=�<A�#6"x��ǈg��ܱ�����?V���f���l���b�xgm͞b�%�@��3��V�����u눬"�v��.�g��B������Ou*��Z6�O�nz񚵉���r�ف��b�^;�k���W�e�;���3[SƏc�3j��콚��0��7,�7��l�w��MH��÷dkǗ=����}�A{|�����-��xe��;H^���/���b�F��8�bC
��{���s�>��f���a����|׵��=��2���e��W�����e��ƯjU���ۂ-؂C9a.���=����sO�r�Ӓ�a'��n����f��v1��s�krS�ӷ��XL�{ϠU�������dx�����s�,W{>Nnw/z�?>��oFn�_4����n���4&j�e\
&nn�w>!x�CG�����pr!����~Ʒ�si��O�M�y���\xo��87F�d����	.�����B�����t�>з���Ǔ:]����ŝ��+|:��y��̜������gS�WzhV�<��:{7�V{=|���#t`� �u�����牸����Ǜ�E���+�Y��wƌ�]A��ۯ�I+���}Cw�j��f��8y��s���]�^Ƀ�ڴ�ݔ��� ��s�?�קh���^\�<�oWny�uNA2�Ϗ35g7���Լ��L��r��aoc��몍�9qb)Y���a���S�Ed������"�p�v�@���o��v���-������/�k��ww�w���z_���;�kSȃ����7�u��ļz��=��i��|�gI��,7-7:}jU�w���p�J��s�Q)������ ,��K�v�Ά[�g�>ʻk�Q� �w_z�w��o�o���������M{}�J�����^�˚�0��G�!�y��5���O�գ�L`sJ��%�Nn{��=�ܔZ� wi=���o��8i��j�
��y�F����k�4m]q��M'�nL�� �z܁^��{f��ؼ���<)g�Y�Z Q�,�y��Uc�r���/\����9�n��vUb�&)v��u<=<Ώ�o�������r6s�i���؛9�� ��J�x�v^���s�+���<��\.�2�������:�5|]0tEe a����$` ���{��9���x[y��o �����]���ݷ�5]�;W��G�v��ҝ�����Z�{��nq���V�_�f��2I�P�i>�Y����̦w���i��� �uv���`/�>u�f��,���;֯M�Eo�͠ԙՔU�^�A����i�r{M��ٌ��9�<z><�*y|��0����`�W���p�3\�=��FF�{�V��D����i�|�G�S��:}�/{����{�2�k�z<��ƙ�կ<A~�H�{ӽ���Ǔu-re��ݫ��:�	��ٰ�G��U�S����9M<�/�nx���[�Z�!��|7�F&�'t����6n]�����ҽ��M���^�ɕ{������.�v{�^���TY���X��d]�Ü�ޥo��Vx��gv�=ݜ���1ד�o���UE�n,�.c�p�o�n[����ͳ���K�:=����]޾����-���Jŝ�'�=��vU�g��ۅg[��{sg�*�����;��mA ��@�]c5<݇�	����W>,��5���j�}뮲v_A�."�}��sV��|s��j�2���	Ȗ��ӫ�%��]�f��p��j�*�͆M����g4<b���g�^>��J��p��n�v{�kE�{���ڣ���� ����^��c���-+��ާӲL����{zx��3\�� � cΈ��ڽcz|&v����p�]��c-�݀B�M"0��Ӗ�Tަ{g��đf��}��?���bw�(}�G�^t�N���P,}�˰/j.1�:gy�V�{&#���jg�C���1a�[�=z�H�2���g�|~ a�~Ù���5�d�x��d�QK��Iq�N�ʢ�����/ �XA�߼�eya>���=��}�M؟�%#�:���L��l�����]�*{�]�X+y�QG.��e~�QO��|��У+�������7*���gϠ=����b���<�<��h^�nG��g;��̾����揭�z��.�n;��R�݁����g���T),���Fo|�ǒG�����S��Fé]>�w4K,��6����5��PqV���j��w��(�>�
p�qB8g>�y��^��kHAQ����ŉ}v�칹�Ѹt�L�l���}�wM�	_xo?+��y�ò��ڲ��ΰ8��p��Z���o4�w���s�:���Ӭ:9�,5���xQFn����A,�	{��O�9�`�0Jíq�{|h�U�b'��=/�-���[����+//{n�p�;�x,�Λ�=���Ǔ��;�n�m^��X{�y�ޗ�b���	�x	�{q��j]�/X����5=�o��l�þU��(��R?C�<��|rh��w��}�*rߧ�7�OqQga���[�y�R��_T�ťe�5��%��α�a��
��*B��&\ͷ˖L�9���W�fÔ!�7�).�x-��␸�=���6����o��������.՞|��צ��=O��_`#|{'�x8�;����ݮ]yg�Z�q�Oxh1���M$�Mi#�
羄�w���'�ª�^8�����N=<eٚ�V�k�=�7�9SD[��{2on�O���|t\c(8������e&�S��\�d��r9��I�/U�a�Lo�=G�t�v�z�
�,k�x{f���#?d���N��6�nG��}�m����;����=�Цͺ)��n���υ/����Y����<&�n���3X����w��s��U�9��ׯ�g�|F8��o����>c9�޷؃�y���=�G[q�
K��g�pvv��J�������B4JQdcNo8uy,>�=�-ͪ��z%�{���lb�(��{� %����9Ԫ��w�yf����W۩��� �^�p�pl_ogG�	f�}����P�{qҀ�wt��y<��6��r��LW�=�$���b�j��l���[�{w}V�w�>�{Lܙ�z6i3�dp�uM��>���`��x�9�-�t�Jgݳ����z�ڷ��!�=��/�}�<��R��`�Jo�>~��߈~��]�$�<+��Y޹���y{˷�1^Yg��b	�}9g�}}�W;�k߽;��.��y1l�3�¿{K�O�8���A�2m/7�z<;{��;p{}�����N�!f!�*ӓ���wuxu<,�o�g-��mz%W�ϗ���|���h`�C؈U��e������xp�w�њ2k\1���2iìs���<7ܺW0�<����7�w��8vh��nyJ{���@{�<�1������],�b�=�ӹz�.+����Di�a�e<DG���={���xOe\���������v���K���+�JA�{����6M��gy��d��w�SfmG3VŲb���V���s~��e�doq1��*��/�i}���������4-�޾+h85x"~y���Y+���#�$<�|�W"uN�86�}6u�Y�M��V@����_�/�����:��M��{�1���K��w��^1�����{Dc͔ƚ	�o����_�����g�'��Ij����Ȳ�˻}��v��F�to	pK��׺S����9ub8�|AI�W�_U�io�o=���iw�ލ@xo,�nt?'w�zQ�|��1�۳}�Q1�O��=��p����\��1�����o`���Y!�T~�Ի��G�3r5��v)�7���y	D�p�uL��Y_�Sw|E�g���a�7Z�����m�ٽ7$��C��X��2=����(Ό��u�l{ ��w'={.f�k����*�[�I��ce��˰�i�ss�R�u�
�������B�4)+�N�<uFc��O,�{�"�HY�~#�3|���������yÝ�.�dB*�3��Y~F{(��'�l���,�Jj3ڗybbwk�6�:�<�]�װ�x��5�� ?g�ň1;�ͩq����Ҏx�g�]Z�.���� {U/9����ٷE��s��^���r��W?k#����.v��9e��ฏP	��H.��Iwʉ�{�|qn�����[3��dy7~{�����,�=i�^���~CU���d`�=s�z	����nh�=j#��k9��2E���/bj�b!{M��/���"�oZ��ʄm�-c�+�n%A#=0S�.}����{�(3��g0r�hn�^�(��^��?I9|�������GqӚ���ܻ��v@}�-��4.�h�Ƙ���� ɷs��WcOL@�!'ۃ��}�ݣ�+�}���G~��(���F�}��c�2R'{� �������g�c���q�$C@�q >>� �I�ŧ`��{v����}���8p�v�tL�{W�x]�Ѳ�%�p[������ϼ��%�,���>�ً<{}�c*�ƈ^�Bib��o�0`5�x:g��������ڀ٢��V���H��g�t��j?�J��V�cg�uV�x���#�+O�(�ɮ�l��j}���7�w�5���J��p�@�q��ҵ�T5��#�=U��@	n�,'<�����8q��Y#K����/v�����4�W������U<|��q�N䟏�|��>�|�,/�v��9�$��B���f���x1�G��{���'���bRxz�Ojl��<Ykt��9���}��] 7��M�^�x�V�F�o���w=���3Q��}Q��I��o'v�sI�q��&�|�̛�}Woz�f��Y�;�f�ǖj��.;�,7خ���ƙg.�~>���8��MY�^Sû~�c��x�\T��
���7�Π��k��3�&���^^^�����{��ɵ2Q̇�g�a������Y ��|��0W��������HS��n*jXq'm�<3�y��s�5�sc��[q�6���콷	����W�Gyo0�!yÖe���#&�uw�z;��-��\3�;�y�Z#�Ig�8��QU�}�<��|������9��ܳ��;y�u>��U��`�Ge�9��c���9�e���.����S��^z�<�n�0�Xq7��ݽ��O䯏5���M5�(�<�G�%�<��u�[9��=ph��������cG���������~�?K�?k�?k���?��><>>3�������g�����_�|0��X�3��&$�����О8�̙�����k⪪���*����5�svA1��2 �M�F�%m)�*=h����SR��\��ݖƲ�T�8�����,�2hr�b�gGMu���2�\�G�f,li���\l�P���$��JQ���i
Ź�f�ͦ�]4�52kPBb-�(��W�36�Il�wZ�)�.������t���u�1H��[e��D%�i,V$4sZ���\���̰���B�K�n4pgT���b�F��A�ݥ��:�qIIk3,]��=t�tLX��e������Q���H���i����3.�bʘ
+]�I`8�y��ie�f��M6�!C�X�\�u���z3bF2�]�G1C�����2۬�������v�i�V]�j�X!	Ch�-Am-1, �SWb�5jqe!�u	�bb�va%��-�l�sb�)v�g&`K���,4
��3#�[eط5"0���ٳr�Df�#S�J�l�h�A#:��n�0B��1�g:(4H���@�le�X�2�\6�ݱe@֐s&��QD�:��LƦmkE��1Gd �[��5F��;h�ݥ�tɣ	c��/�֤�v��R�	P�j� ؑ��C^�vM���sM�0՚i�6핊���[�6��%��l�4rK\9ͻ(�K�����H-�w;#)U�E��5�)ۭ��6�P�n�ʚ�	�M�5�l)˥�3��J�Lʼ:sChiMn%��6��6�ǎe�6�5�c[IeSRcZ&�^jv(�.r�4��E������6�f�+%�р�)k.�3B�B5�6,n��0Mf��Yl���c�]�P�F��n�12h���I�,4�ٴ�m�N3	A��1p��� ;A�L��+*��pf�ƎŹ�3��JQՄCUNB ��l�&p2:�\��mu	[4eɜ����:�D�6n�ce�R�(���!�P��)Nn:�n��1+Mr.�M�V�v*��Rg��X�@�YM]t5�Ceh]T`rbˠ�aWD��K��p�4m%�0,q���F��������c]�ʎ�ݠ�m)-�un��C����A��ڀh7�5�x�����l㛖ᅑ�L���V\g[4�d5��`����`��;�t�[��S-�XXKu�dLL��3BW\��i5Zb:1��Mf�fB�e� ��Za�6m��٨6�#͸l�N�aVT�clՎt�!�ؼ�]����%�bekk�nec���)�dB��̻v3�0�N��\g)%��Pڥ�`���l��T�gS[TbV8lҥ�5K�ph�Z����,�DD�,Ұf�8���K���K���f�X��H3ipq�fPh�SK[�`9,kL�e&�Xh��#z�4�A�f����&V]q�!�LFhE�:iH�\�BR��Xlm��s`ܹ�����L��B�MKH4Ԓ�l�5m��4z�2��K�#��,),j7���5-7C��Sip]��&Fm���W05�KU	�&�n�Lۛ\����Ke]�8nK`6Q2��7�R���V�G[�"V6ٔ��A5�ha�j�&�vD��P�P��c&�6�iev3J$n���؅���.k.�Й�偊P���.��Z�NЦL�c!D�f�r�����+(FJւ�2ZFʹhڜ�-Cb�JZ�n�):UX�G	\�\FCn�m��-�
��U���+p��lP�b�]z�45�CXM��4���c,���9SR8(]�ׇ8%�L�sj����K/%l�ص�Q��U���[#c����f�ڀY���s�c(mq@٣���io$�f�aTҋ��֗����U�q�Z*����KeMD4å\���m��ױ ��[�,�i�a�0Ձ�ڹ��p�í%5�gj���N���̦��*;k��G\��f5n55��Ά��uR�Z��n��H�`-�`j1:�FU��˩m���ft6��G9�,�+��E�Y@ؗMF�͈@������K6����Ջk:��-�G)��1�\��D�5���]j�ō֝��`�!���� �@��աc(���aZ[e�)�R7k@ڮ&�ljd��喨c0	c*�T�J4Զ�%�b0R�k0���3[+�l�If��s)M
�3S:R `qneJ֕��hcF��Ơ$٠-����K1n�f-r�Ze4�,Z����F�LMVa���î{f4�Bj4����[����e�6YE׬����fl���\�؍��dÄ́��I�)Kts���"6͇:� ���豲P�6���"�%J���jkk�i�e!)P,��ܽZ��aJ�-(�h��5v�	i���쉖l���������2�]�%G.�Im�1��1�Yz�X�S+j��I��Q�.����+����%uV35��GG����s�vY�� ۞h1��K��^ջ�،X�k�m��J����L`����&)�5��[/Y��k�Q���̴B�� ��t�,٭���pv�hΤ	\��r�Ƴ@��D(u	�5X^l�YFP�eq5�)�Jk�=�1t�bKJ.�$-a�]S9�tj� �tWL�����gj�F��ҳ��.[ٻb
^ݵ��;Y�����꫉K�0�p[�V�p��1ك���1WP3�c���]).W��Ye�K�#0�xCp�e�v�h��+�k�pc#�m,�I�c�n�)�!�t"vn-�"��٬afa��� D6�A+IK����B͍YD��ƥ�-*� �����7�6�Q�h.���&���6�D䥕En�U��H��LPK�T����*G��P%��[]
M�6nk.�W�Q5F
5�Pr�d�XZKb@��r%;f�&�!S3��Z.qa��52�07J���f�T���ic�`����Y���`��`˴�MK+��fSF4c��S�FPlY[u��X�Cj7i��ѷRn�tЀ����q��k��r��l�6�fev"Z����$.;4,�`���kI�)a,�55�l-�n�Z��fk�9Z;�#cJ��3���z�x˪�]V(�^-u]u����54tV4��]�C0���ݙD�5��4�[�����R�3��%��4;f��6mΦ�ˁ	bW$�j\F�u�B�f�r�3]��m�݀,*YeE�
�2��q[�\\�����z�Yj֑�E\j�������\˞\�e��+��mәnsV6k�a.�L0cY�«�jY��\�+u���HY��i���0�Ij�bh`�@-F:� �um\b��*sЮD[0�dZi���QІ����ivp�F 6��b��쥰b���!�jƬ��]�[�XE�%+1���כ{@$4aln�Aq4�{Rlh�"�(�,cIc	��t��M�\-b��F8��.!5��e��Hʺ��p��]��.l�X=��b��׶W�&��\2�8V�Z�Y�l�j�M�n�D�55/4���(��.����+	f`mjM�R	�p�I��F�-�3d�S&�Gp�v��-��cc3;���˫׈�6-&Ԇ��m2($qn��e���QL$h�R�V�����as&ap�+�F���"���V��6b&�s���b�`�c�8)ͺgea8�b$pڹ�-�L�j��F̹5�6E��6��.F�e���ε�����SF�KCk�B[
�pF1s1�e�ٓ��R�Յ�q �ri�Q�d����6�lbFk
͑RV�*��B�X����+p�(-�3]���C��j��F�sX�u���0,�R�M�t5���*�l]�3m��-��kl����Rlfn6!K�ɵ� d�Si�frkVږa��lc����u�(:9�.��CD��ػ ԃBV���gMm���*XM�D�)4^&6-�l"�k���DQ\R؛Q�(ܲ�#�����K�bU(���:�3�d��
͛xhh�taˠ-�f�����8�c,P�6jb�c���Mضh�4�bi\�Y�W����I�H�K(�[��K�7:�i.10+��\�j�v�[��K����nCb�����jT/`U���47]�@�$���ۅ�΍Z�)
F����c�5��65p��:�X6:0�nmK�@l*p;m�]l�)1���N�[��v�1�p3�$�<&.%�r��R���$x��i��D��[��Ģ��Z��f�Ɣ˃u*�ǉl;&U�MM�����m.��26F0)�qs��&�kU<�q�A:���KY�����KC��W�Tݑ��2g�Y�x�Ҏ���q�m&��r�E.t]e��,����,�5��M���,��b:4��WY�&`���u6�V��e��bVKL���ͭ�ű+�EW �W9#c���lL�Z�lfS-{2�њ���.�d��f�$+-���[Y���"��YP�����L�&]��L�X2�����@l�ˠGm�5�J05u��A�X�0Қ�M-kŻED0M�LX��m.�Fl�gcL�D]��q�l	b��4rP�.n&�Ҹ�'cB��)c�LM���k2�;�Єm(��3j�ܱ�"�X����܁���\�&�iP�ɵ�Tvն-`b�հ*��!m78��cd�"0��Ͱ`�1����i�fo[Z��Xm��f�*쪪�ݳڬ�i���۞�����,�3t���.a(�Fg&��\1��s��:3(����mL�fPsJ����Q�UUUUUU[��L��d\�U*K���x���b���r�o�y�-���M���|�y��єf�0�In�Б%�u�wu���\��r\�)!�Ŋ�6@��]�f0.�8I.p	'9��H4����w�˅�uFX�I�]dD(I���S�ܨL�J#��ӻn@�ň�u�����;��I�o����
���r43G��$d��b���Lb��cAnt-c�A&�$X�b���:��m�v�9��9rƊ0d�j)7wPS4b�,`CD����$���+�B�rdIRF7.�H B!,h�ns����6#h��1�{4h�X�W��鯝]AI��B���;��IDQ��j$�2g��2�b1�y^<�Y-����I>�ߓb�:{L�lC5��!����CFdn`���01`�bYu�f5]5ػG��jeev���X6it[vdуE������.�-l�b!�8�d��lC^r7W��%���b�v�P+1f��a�[��4&9�p�5fkSUђ���"�m���mj[l�k�2���,v�ǲl髚��[e!����J��Yl�k�؍�f��R��,Z��<Į���֨U�3XS��+^�Vu��d��9�oJ�MQ.�B���^��V���h�DfxR�Z����U9K��6�JD�-%+�MR)�*���롎�Qqi115�HK`T���Rm�c,�U�V<�B���SWJab��f�����;Teְ�5�,������3�%�P���u�ysm�MVXR� �$.���l�� ���8� ��irUΫ�v�79�ld���h�^ݜ�+�2�SFj�#Q&pMu���^r�X=��l���b9*�Tn-�1��˸��]�-U��D���s[2�&�T���4���v8��u�+u�.1cڄcq]�d�7x���F8�[�L�Y��hb��k--�P,���
���͵�KQ.q.�l���Г��U1���-�xR�]ms�л�s���-���\JPn%@G[�!ۥm� �"M6��w-0Ŕ��k����ݜ$�ƬR&�щto6L��mb\[IP�p����g2k�C�4�a�4���˒��eЌҔK����%��i�$�`��֋a��kͅ�%�WKfQ��H��+ke���G�C�
G�(m���vK��!)(�j���Nځ�u�o3pe-�5i��������Ҩ��#�R�A�b��a���ڌ��Gi��6�Se���X�a��m�L�ker�� ��Zc8��5��ʨ[.��v]�.vs����Kx�$�$�|Nf<RR�Z("ҥh��!lbB��Ԋl�����IѭY,�%F1���hU�V�-��6���Zǭ�V�խh�m"��B�(��Q���ձ�"�Jp�Kc�G����[�ʠ�F��[l���,F$ ��@��h�ט���U���]�e�B�lB$H�R�c%XX��ƫ2�[ ��Hf�r��d�鷛Q�K��6@%,��"�>6���S
f{Q�@$���2oyT,6��$�%?�|�����ܗ�:�.�b�	�N�I k6ڂM�����>��� ��qዧt�0IЃ�s�A�U��Qrq���|��$�Yu�>���箃3���x��ӫr×�Ɍ�͸�A��r��r�~Y���WG�C!-��A��yA�v��A�O��=UC&�ikR��x�$M��A;L�����B�K`A�G�6k��Y���
���rɒ\݈\��݅��`@��l&��x#�l�	X�߃����e��� �3�+]���k�
{�&��/	�l���x��/�˸�0f?�n-m֮��sYg���3"�U����	�U+jzٱ@�Cf�׋@�ǪYM�Z�<`�����jj4���DPm�e�Y,����a��c|QMM���}B�z#waW��Ł���Wl\�N��fzz�p�T�P�Hu-{�Z���i����� �S�g���.T�b�&t$�T�;����c��0D��ƌPH� ��
Ȑ�f�E�:�8�g|	*w�e��݃y�<zZqo�-�`�"b��d�il+�®bL�F�=�$�6q�S�lYl��(Gצ4)�)c��;uٶ��N���$%�ڦ�6���`�X�8M����>ݾ̕hϰ���|�@^����7g"Úd�����z"	��}� E�q$K;�������� C6������ȀI�܈�>%�޵�׈v�8	��5ӹN�'�D�I�I�ج� ��^�5����%� ��"��6~x��5��^��I4��^���~�\}����F��^�ᦃ�sG�=��;��s�b��t��@��/1di#-�LNF�Ǣ�m�r�;��3̃;m/jThFKF@76�` O��������h�A:H��`��d&Kń���n� �^��-W6������ A���@$���~�ħϑ��9�毉�,$���et�(����S�p�!a3�.-�t��D�}��n�gvv�{��/dA"|�o'�'��:��)�V�ڎ�9�H���0g��)���m��g��Ё��y��b��h7�I���|�$n��<tIpکR�^�9W�ECΊo.���[�`��O� o��/9C܋%���$^���u�x����`�w,؂D�F��t(�)�X���O����ź�g�}}0H����^Ȥ�_'60��ޒc�v/�~�������~�+�����g�yu E�:w�4S�3���b�L7!\T���CF�͗9w!_�o�	L�#�ߴ�
-�N�ѷ��@�m�Lө���'TcT��CeD@$�K[��
�}0w�{jڿFA#��	�XM�ójf�K�ZɁ�f\i�j�.4Kl�R�̺ⓓy��K:,�8`��4�lH6�� � H'ծ�c��i�5mcguƃMm� ���q�M&�1��ޯ�8\��}�|��;=�� `���2 �� y�����	�u�/נ�Q�-�����h"H5��˘f�1�*s4ӼD_��i� �o���_�h�X�SAٝzm�2�������\�L�A ���f<C�-�ǈ�V�����	��ǉ�8b�6:fY�p� �k��`����k�f�f�
���9���rw" p���K�D�#k��k���oe���z̏=�77�\Ȝ���N>�������{����w�A����s�ûp����-�f�!�xc���p��������:�Yj/V�V��\�f�la�xˑ�D�.�;G��Y�����mV6�y�L�J@֭�[�Z�f���h� Ӱ���ی�	]��Xb�@���M3U�����ds�X�BV�ff4�6ʅ�G�36��V�6��U�&�(�h��d(R=uq,�":�,�Z˸��v�
�˸�
��,cԺ�GlU�p3F�4&GGm�t�Yc�.΁JM���ƚ&-� �#��E�@�y�SK�xs�:��� ���]���O����p����-��S�Z�5�� �'�f�|VD�L��L���̙/�U(��*�����7-�!x�����rr���*�����O$�k��wi�'��3{�N�E�Nt�מ&�π�3ܟ��~��$�
�Ke��1㰣�ӭK�ªB<H�$�DO��q]����m2��r@�m�0��ex M�JA3��{} ����n<Ҡ^����ƴ|Cz*�} ���f����^�{��3�E����V�׭˜M
�s�G%�ęò�1�l�C(����,�(�[)�9�5�]^�枲%��E�����t�Ēb�`ATom:��� ��d��	���j/~n?΍�Q�q+j�x��fRy���2v�"�C��`;�-��Mfo@����;���zr5q�e��S��|�M[�$�v�P	)¨W9%fNRܶ�Dzv50�v,�0d�H񘍏A�u�	E�/i�-�J��J�i ���	#S�4y��mjt��8Ŏ�^�ܸ$7�7�X���@4OZ�A�����jɉ{��"]�b��ͫ\�3O!����|>�7����5Mn2�ة�����DO��:��x�kZ�ˍ��� ���[�&�x�J��������ay��Ա{ef5��6k[t"�J�Z�����p�"ά>\���&2��'ě�ׂ۩��H��{q	4�q�3�c���H��'~�W> �1�\�e�#�
ͭ�	�b�ƀI�� ��܉~�}/A��q �h)=�2of��D���$�#ϫC��;�<6���0��^rڨ�s���S��C1��3��ٗ;ދ�;8�ӆ�>=�Hz��b�P�oc/XhW�x-V���>����I�|�|�;�������!7�,)�-�V�,�{�Dy//yψ ޽�A9�uT���V�6�zLM5�<h�d���X�p7�A����k�.~���}���}y�	5[�#/"�J�������H"[��X�sf�b�b&�jgXE����
 m�`�1Ɵ=O����36�ÍL=����� *sb^Y�͜r���V��M�l ����	>g�4���2d��O�N�A������\��a$�� $�f��qD��i�6�j�ߥ8PoB34���̍��H����ۧ�|.kb$���'T�}P�Y�`'Ĝ�ǀH$�؃�aW����8Rs-��*�0����ߜ�3 ��؀A!��f͖47��`���������m*���Q��_��8��7ٲ蟕%��9<9\V?*���Q�w��Q=|��!���#�ˉ`��ǌ�GÖ��?_8�|T	���G��d/B� eY��o-��MCeĖl��A>1�o�]�$!OUHA�}z?<����Su�8u%����gR]�4L�j���qt4�M�eI���p{�6�d���y��	�{́�[�4Ta���c_)��>���}뛥�e�m�� �����qU;pn�[�}�}$����f�P��{X�߼߾v�5�<x	9��`A�,���I����u�2�	���<u��~x�c�,Y8JAںr�ܾm^x�@8�� ��)���^(�>�D���.�".�%��=&�س Zh)9��N8u��m�?ߓ8��f�"	��ϣ�1��ۆhl�%yG�����Lq$q�����җ�@��)����~��hV�aU�}�3Ƴ�˳�v{��l�g��Z��4����g�}��q�
���T]e�X�Ѕ��Bi��]�j
�I�*��GGb����XK�gM���q5��ڕȩq�3u�2f��e6��:3m��"A`t!����B�3��ٰ`�^Ά�L<�)
�iR8�[Yn6l&�^��8G�Mf��j�G23km�DK0�K���8����F0�i�ta.i4�uR��G]�KMn���8ʶ�˔�Ե�UJ�-��A��[�-�e8�V����]7GA�.����;\�,��.f �N�6G�$�}p��bm�4�O�2M�d�8]'`�X���5����ݪ�]���h��I��� o�"����xˬ:ZU��"$����;��߯������[cd�T�:��x$�[Y�	�-���g8$����sb7K䶂��b<H;���I5O��/���e��5���c�͔A���Wސ� ��@��x��	���i�ǉ��<x�#7�[C�\Qb�H�M�ڲS;�)��)GV��Ie���c�:�g	��,�'gb�fx��yP$X����>����3��Z�=�Ժ�ޗ����0 0w�� �tJ���g&ٙ�� �>�1 ؽ���k�y�K���bo�7�wqQ����y�uj��~A�'��N�"n<�Wz���r����qE��.�;���z�z��>�{SN�@>�}x�A�܈�����3F�dN\A�HY�&��I�; ^dy�H1[����9�� ע�)H;���@��� ��>�=`�$cM���̬3.�D(��m�$�i��!�f�c_b $�f�GF^�p�1Z��KT�S��;�Y�'3&#6A�[p�7l��w{m�Z�'[5��H/��D{Yn(!�~[�������HF�r֪�sqТY�m���n�e�������gi�eT�Ϟρ~��1f@����]<E�o��w%��,�x���ֻ�1BЍm�� ��Ǉ;�Ɏ�����ذ��B9��?d��A"'v ��TxߐW�-�	H���~�e�I<E��ɂ�ݐ|3�7�Q t�q������������㏏�{=��o�����@7w3��21�0�F�_-&����k{]w��p鈌�P��b���7��bv#���)��a^�gb}��ܷ��oڏ���|�ك'�Ɩj�TH�;+��=��˹L	Y6�ځ9s&�XhQx�a2�$�����?\��zb΍��Q��ܕ~�c���i�Su�[���͌d#8�qyፚYA)qrD���/�����b�/����f&�O���O&�^��6{���p�ds n[�$�۽�`�G 9�b��o�ע��Y�WJy��O�Ӱ_���#%B��P����֩ہ��6����ߧ��6�(5S,mL[\�yvUrF�Eq�<�}��M���UD��,����hjڋ~��� 8{8A�;������;��`�������;�����j�E��;
J�'p��mS��a84��D1`��=2�!����9�0p>�\r��P	�������;�}d`G�ܒ��8c5��z?zJ�oLݕ�}�x7u����y�L��=���w�9���tw���@	������wQ�&Q�����7˻�&��c�<�����p�������ĺ��������'}7f%O@5eS����K7�!����%�>	�����1X����C���n�/�r���ֻ�%�u�*����{/�����sП_L�cۄ䞡��xpHR7�˽�����gN�
�<�ۋ=�=��^7�z{yvz�1�>@���M�߬��m��p���F<h�������F��qA�B����]�^��Cy;�4��b
2f$���Dl�)�4�(����/q�����#r�E�.u��BD��Ȕ{�1��(0.r`�c0���^t�[�M󺄟�f�.\̐$�`�K�M��=݂wr�#'w1��oLQ"��v����)����y1d�(c�|���7No<6�ي>wl��$ܮn\���:�wzjg��P�ve^��F�<������H���s\����t~�����w�^#���ή�wp�#twR�z�ۯJ�Nd2�����RS��lk�WW]�wnWf蝜߷t����f2r�r��.!�v�|��i�;C��t/���tz������pw4���9;��w-�I�̽�5��uH�(��Ţ�@���HH�����X����;�Qv��$����)U���E�v��wr��{�;v��s;�f�T��Ի��8�S���[� 'CY!@l�Q��8ۭo���)B�Ƶ��rs�VBe�￺�v�d2&��
;վfnY���$��=G�{���������?�w=�dK�����<��>6�lC�g�o��Ghzd�z$�L���3G�TF�E���" c�|"&*� �#ì�s�Yb���t��$델��巔��0���5�0� �uӶ�s��$I��&� xI��>�S'�}��h9e�1� �sZ����@P�`f�#��NC#N�\�*f;`��;�*��g����8�똱�?_ͥ��If,����"gqǄ{�� �:�o|�v�䌄�l��L�%]T&7̱�������9�+L���ָ�����|β�{-��l��P�9`3�|�'�'�L�+]��9��Ȍɷ��I�#��I�7��r;C̙0m&Н�l�������"�D��!�h���^"H�B�<o�:LS��H�=YR��6���R��0O3�=�x�
R�d2M��~��w�}��buHd�NG��Ǽ!�rK��2��ms��t�N�OϿ=m㙜�[ry8'|:"/��V�Mצg�#������ #�/d�|�8��(N_6���w���LJ>�I�Ǆ >�5KK�k�I�b]�l{�Z|����|5=M��Ƿ��CH5,��#!��*02��Ӓ� �Y��8�h�����܋��#�|Q�������D��B-�O�������C�M������2r%�\�;���Iy� ��Ӯ�=����%s�>p��O^o�pN b���������O�~p�������jR#p([����6L�E���*L�B9�m�v���=|�I�Ѧf����B{d�����Ҕ��y�ߋ���	�x׾p'1�l�zd�MdIL�X��K�#�B��.�c>s�2sI��:έo�o�Y��or=C�I��ε�rI̸O-�'��s��c����Mw����HvFG�]��{�<s	�d�2l�Jfaǿ<�D�^�%~,@���v��7�p�����������U����k:{�����/Ĺu�[���s+x���"<�%�����T���>�6�hO|���K�@d��ǿk�'�IT
�N�$��
�4G�x��<�P |���'������߈9�,���C#����9$��!�X��;�}�܈�њ��o��}�G�ټ�|$<��}���fw%�˥��C�&G��t�$�R�2O�ѱ��@�H�;���1�B#�}S��rY#�JQ�>|�N%)J��<l1�� ��n�Y��w���-{��������W_Z6�頍���p��?qqa[R������f2��s��-��,����]���+Tux�y�0q ����@��4��e<���	���ٛ�kpa�j3a��ͦҬ�.�Ya�TQך`�&��݂86��6�ąm����A��	hbd.���hF
!e6Ֆ����KIc�H���\]-�k�,a)����VW�.qoiWEXZ���K�M3+I��X�b!Bf���D��%�%B�B��L�$�)
�vYM ��s-Lfb�Ѭh)��P\c\ځ]�A��!���n��b2�5�ZT��HgT�[`�l�Yk�b �K�n��(',�0x�Gw��D���6�m8@d��Ʒ�JNa���;#�G��� �W[	����
>�����#v]��<��w�9�u�HHK��gg`�H�|�6<$[�P���9�rt%�<�%+�#	��u���28�Y�1�w�`y�G�>�'�k5��ک�av�r�����N�G���=�M�MS�މ߇JMuַNd�\�$�A����:��w�@�|#������^�6�����L�;�w�qJ�L� ׻���؞��R^���~}GcFo]"OD��p�{[8K��cƳ�}�H���s��<�Pd�&�w�p;C�&C�d�>���'>��s����b��<�����2:��w�9��\��I�v`�O4G���SeG����$=�C��C� �@���S���5!���q�s�)F���:�rYrR�}��=�y9!���&��V��V^�����rSS��v�Ȋ�ֳB�RcU�e6]��R��Usf6�mB뵵���اs�ďp>����|s.0d�˒u���JC��� 9�:\�	(�y"�Dx:C��Ǆ(Z�X��:�r:����m���K+�fO:O���m���ޡ;N&;@ ������vuh6�����V0�'Y�i��-�b�5[���4_>U5���Ѫ+�ز���<�q�y����W0�DWN�Balvq_��Dv�?�e�R�rN��x��2$�K����@d��\GEy��;����I���d$-�I2w`�-��d����rS��S3��qĥr�)I�gY��vk���JR�#���� �%�2\�ָ��%(7L��MJ�L��X39��#�|ծ �o�b��v��Y�Pj�/H����aB�m�7��^��g�JCx�K}���!$d<��A���=amu�YÞ�%�G�(�5q�<�� �^�+��m��͸:C���w�8�`2R�	r8��n<��˿�����[{��'p���q�#��&C��.3�k�x�^H2�J8��7�9���;�5��������M1��,�t"B�&���+m��ӱql3f��Q��߹���p�,Љ�����T��o�	ʹ&ͱ��m��y���R�'�]�i�}��9�嶇~��9�@Co�hϴ�1�<�}�@G�D���>G��C3)����o���r4<ɑ�>��s'2�	���t��g�-7�i𼇘���>�c$ٓm���y���L�S<���q����Un�n�5�����G �C�ɯ��t��x	"Y��q��@d�1��G>��a9�@���"<����pXu���i�L�dd�#��Ǭ��$�ųPk+lV>b�v|�p-�\.���Je��_"�^ZV�6L��e���F�]���@Lx�=�r��d�9�Ϝ�ļ�d�vE����du�η��5�V�+!!nRA���G��Q��� ��}KA��������|G�Hx:��s29a	���F���9���>��}��zkG׼O�	��7U��=HN�C������M���'�މߜI�ϝkp񺓩p�%�\��v�\2���&F�v���5�aπ`B#�i�#�ADx"���wt���L�s�d����uAe���(��A�$e��o)�%uyҳS6��Fj��\,�٥1�;J�l����q]��)�0p���7J^I WlH2�Iy%�ђğ/>>��3$UT��)��K˧�D�^��\F�d�����<��|�	�0�r�[��6�6ʎ��ր	6���l�&B(͎譶� o%��B��/�[#��7z��2w.��w2e(ͨ!$����"@���[3��Ѝ{l���It�H�(ǒo]9.L�7a>���N��9��&h�h�
�hؓ8���Is�Ăd�	*W/>J���Φ����'s[ydD���y����nkվA(x��؉	ׯ^)����a=��O��	��s]��nr��8��XV��	��W{.U�='���� �F�IE}R$J^_) �.RA��+LG� BI/%�얙G�1���,�Đ̌�2'�C��3�ǖu4�>���9+a	s|Q"�2w9Iܩt�W�Ѵλ��f����u�\�hEkX�Z_��g�1u ����73���H�/��`���t��HN��[D8{�9�%�L'ܗ��A	f�H����.n�i��G�g��̂�aW��_�L���Z��^R^@$<����QA &�$H�n�v���'�dΙ�E�� ��d$�Q�ƾ��V��Dvjt��ׂ�$�X_�BI#��*D�Yꀝ�3��ŝ̙J/� �%���n���t��T9���	v>J�"Al����+X�=��m($���Q�|�HY���;si��ԉI%��Nl>��a������ĸ�d92;m�i	OOl	��x�Eim�[��)���?��$�al�I�!�f�)��n�WnN�>����Sk�$�Y�U(<�_�Fc������	��aY�[YNma�{��~�����5F��%��附l]5X 9�-��+�.�j�v�YuB�[YU�C1V�R�C��cr[ı�mַF3e�M飅�d�mhmf(�PFۇjE�Ѷ�ݶZf��2-�\����x�o)FYm�3�#`jRaU� %����[�Ҭ�:�Zcuj��M�`�T�)I���2i�Lն��i�C�t!s�0q��M(vL�g2��D+R�5��H�;M�Ym8ձ�ʮ��mn�nsG8���>�������&v ���S� BA"z�%L�I-��!#�{u�*���ԭ闔��K�m�T�I�$�
5��D3suit�@�	R#�X��S�~���	.��S)$���D	'׻m���J͗נC��-�q�A; �LH[�X�R�32W]1>2�H$}RN�5c���>�k�a$��%��@��{dH�549-�;;���'�UaQι�.�]��g5�H�n�K�Y�^	!��"I&@�����F�Bp��Y���փ#p�@t3��ŝ̀e(���e$����"����4���F�^I��HI$��d��PIr~�yH��ܜ�����	���)[Kx�wt�ى�mZ �C7�5#�]��f��ܔls.����l>}��r�ț�'i�n�|�)y,��!$Z��^|��h
�s������QI/-��g=�ʈ(Ӕ�d���0���}}�[�&���*�ウ�i��TH6�p;C����&�s��bi�V�=Y�f�I�����x{WNϯSXkg&��_�����y�hD:�E�A������})����]�*�Ii?�/) ���A�9����0��Z�E_;�L��g5D�OFA%䨾�9$�%r��.�D���/���#s�	������B ����0N�8S7V4y�{g9�M`H��葀S$^�:^R'|�ϱ1�>����i��H�v@�#"t�D3���I2z�Ro�f �X�9�	G�ѝ����p��&@I��?l� �K�[#�e8�q�;4�rA�X�	&vO�(������]�1)-uR��+�Ţ�1�VN�Gw��
d6Bl�&_Y�4�^fe��"a �+�'�ew���P�) �;dH�IC��K� �la!"��s@&h�iS�#��B��0�̎��%x$�'͗��(-l�i�I �ǂŅ�lAٴ � :(2g`��t�zW��2=Տ2�I"<}U9xcٻ*�e�7Wa�1�J6��R-7b�پ�}��d�d}�Ϻ�������2c�"��7<������g���H�5�����3��k���>B��#�&J
>��>��q?y"P��t��J	vO�2�}"k]�	�ȳ��K��=��s+j�lP
��q���H$�I^�<�I$�����ŖJ��I{�m˒�2щ�0vb.���r�D��IEvę>�wB�}���ݒ`B}�y	 �	Vμ�F|�{dH�Y��f�2��	 a�E �)_�a-��,ŮA�P��ؒ�;;r�ChRj����q$��ܤ�<o)7=3��G.y�R	��dL����-(C��I�w�q���$N��̤Y����d��w2e+���d�|��'^���.:l�L_�%�Iy8�>�I �4�m
�H�z���T&����{�H���		NS��Sλ��a��J{:$%y ��u������ECl�ϒI/%�:�(��Qݲ ���P�Q��]�����̀��6-�	S�SNbI#��I�$�]��L��IO�.||}ox���:��j����ת�J��{����bc���\ZD�+�Hd2���[]�{�B.�_.!��]0�S1*�����#ޣ�xxQ2U\�F�R�B��
�J$��>ff|۟=ۙH�i|��O�L�]�QՑ �I���!uVg/�A�o������H���dA2����>��FF�])L�(���0)��kZ1t�B4���,�Qe΅kYP�	v��[���
��R~��>�v��b��m�l��!$���H2JH���C�H���d�<%��۶���J ��Q{�&V���ӳ��I2y�RnzfH	�}`˘�l�*�mR�B.�D�H�5>t��$�����{��8���8�%/��ӤY×�d�q�/�$��>�H��K� �3<w�^�U�M�v��I$���$L��Ij|�y	/���h�$Y9Nb�O<��]ց[(���z��3y-�ȓ)"t��<��I����ӎ���&����L��BB*�D�:"|��L�0�@%˧D�架3D���M��p���2�Ib}�ru����v��P Zgggǧ��Ǘ���g�����z��v�V��P��a+���]-v�m#{�k~�0�:@ģ�{��dF�m�=']Ԥ�b�ϔT͏d"?f�9�s��<7<�p��~��nD׎nsW�����AAcQ>y�G��c�E�K�L��wX��-�������K�YՁNv�_h[��y$Nޯ��K��� Z��wt�����\�le��7Ր���;�=�3��3��D]E[���0�Ns	����G$��n���Vv��3;S�Sn�^N�Wg�۸>it��1��7�^Ŕjl̇��e���%���Wp�4f�%si{J���Џ_k�VB����<��N�^T�6]�:�K�ѵ!Y/��&�޽�-��C�ļ���O}���������byў�>~��Ԍc�`��r�n����W�۶��4��zf�S�}���WaaDZ��٬�{9t�Q ���NU�cp��U�g|�24�w:u�<Y���R�=��; -^��c�c��x��P�yn{�9�-�僃h�*���#�,o���w<J�ekuyB�{N��yuwi����D�1�M5b
=�/|�;�=�N�
'�9��*��s>�Λ4���ު�^yq�מOz	�NU7�ެ�.�Jg����zjA��}[��8Rʆ)���,������V�=�8:J����S$�>��x[�n�{�z�3=�>��wi\p�zoh���0�,�P��}�c@˒�,��}�Y�D6�˵�#(2l�[JG�s$5����1���O��f�g��=ݰM�z����3��pj�������#H?|�,g�y�*M��T!�Z��VE�ev �R�n���\��z�SB�$�����������<��ӌ���,a����u��1��90^�e�uۺ�r�np�t���7+˛|yy�uݓ����l������{�	4�W	-��t@��V��9-;%_��/v�c����!Awa΀��� A�7^�̡�n	� �7-�{�����wW#F�p�BP�ro��M�{����������e�<�;�;2@ab�3�r4�pI��5<�ûy{�w"�H��nWu�7.��nr�������`�sv4�r�(���ו�|[���h1!�t;�$�{��.k�Ƥ�Gu�t���B:�1��31�=۳&u��e=�$�iW��� �r��2F-� ���g�wr�+���͵�����˅+��J�=FՖ�Ci�M�3R0�M2�A�.Liu�SL�lk��-��`�Fd�4x�"iv�2���g�LE4�Y[6�3Y�m�[�hb^F[(�h��YLT�m�mm�U�ZXq3���.��j�M��I�-k6�����B���6�d�ew:Y`0{MK�.K�Y�2͐��;T��3�8��UX&s{1İ�������ly��кmK���r:����&�ԅ�!v��b^^8�M���Kfe���fe�Ja�(L�^J�\�Z9KcK���2�]���ka��ܐ��6�H˛t6�u��
�i+Jjf5ixs+z�l٭wQ�S�` 4�2�h�ذ��$љ�<��^����[Q�ׂ�v�Ի:Yw)[u@��\�:�"����l%ͦVF����u"�Ķ�d�G)�s��W5-�"`����DP�W��5��
�(�H� �3�f�Ǝ`0B�vvl��(�Rb喪[�[bGB��6���V3"��������Vh�U4Ų�Rֺ)i���(FnKS�]���6�
��q�͵#/i.8u����[	6�-��;�q���6h�t�Ո�C\��\h�j]e"�RԂ�kZs;,ݔ�[�3iL:���n-�B�#5ƍ4Γf�0Q�����KR&	n�z��T����ݝC+T�Tl-�[-�auG7Ts{��tX��2�����1T`J�ni0���e����N�8�lL�����M5i)��j�w$e��Z��,��W�+jJ���Pw&1f�� �K-v�̓��Y�b8�66u�8Xh�.Y�лbe]�-����kr����d�s[6�@�l��@�����%�\�ȓJSF�*-���^ݴIzҋ���B�Y��4�P��j�Ñ����P�n�c�6J�.1�K�Qn��]H��Wl6��֦�̈́ٵ�ʹW8ty�C�y���1�����wN���$�$�HJ R
��5��9�o�e��ĩ���ʭ&�B�Fh��)�Њ�P�H2���\�j�4o$&����Čڹ%i����]��bbʠ8���W�aL��Ա�Ʋ�J��F���m�YE3m^0h�,��qJ�YU�1\9�q��,[��>hyK|����c�n�h �Ki�	��h�[�f�
˨�[��m�������a{Qa5f��*�+W.�4�+�ړf�vRSU��J\Ŏ��}��YCD�d���3�չ&RD�|�s)/$��y�B@C�{W>d��efȂ@������" v����
bW7e��GȟJc �y#�F^�do���IR~�rd$����(�$sS��L�9����+���t���ܤ�<�)7�3��[G)��$���NCdG=I4�le�"P��\�� �^9H�Va��tܹA���U$�U -���t���e���}	����z�I���wl�V�)����
	!+j���/&�>+Fy"�:s U�����W=�&O��Z�w��`?W��.;3)o5H�A%��"}(�qu�֟d����"��4���0�&#�\!T�D�3h�Y�B�=�c�~�,�)~G*�O����H#�����1O�$�]=�"|��s淸����*^BI$c�)Rq�kY�2)���ڨ���@'���Q�ݝ���}�+���ӧ�?L�_
��&0I�� �B�khU �ɫ��x*��Q���Wf;��p
���.=��}��8\k��s�s���� P�"� (�$��o�>�$�	/^<re$^]?l��RGۗg�,�m��zJ<�Rt��
 �6R�J� 	uFęA$��q9�"2#k�!�^�A$sΩ�P	/��"e'�un"���wr�2{�
NOMH�D��|���y���)���Z�>bJ�ݑ5�fA$-Ft�B���;+�Ӏ$id�H���>vAܳ��ɐ��TO���'ܟr$B�-3��vtd�0Ih�i&BIVWH�E$��Η�����6��}O�?cP_���s�[���2��`�I�SWi�v)c�ҡ,��z�و�_�������FD���s��^��D�%�]�A%�O�/)C^�$y���j[��D��I^VșWw�PEHv!"�B�f��Q30���;1��B���.�n���@%�["HBHr|�y	?�3d��s��k�%*rA�Ư���I����3ꬉ �I���9��T >^>=ֆ2t��8�AY..����W3�7`�TZ�fq���w.�n;1��*���T�����TQ��O����1�t�,������=��>� � ��i�"R���2�ə/����P��u$��9���7F��.ZJ�ĒQ�� �I�'ܗ$�\�<� �gR�ð5�.:��G�^����A$)n�,��0�q./���2�	~�v�>I{�rD�	 T�r^BI$��y�V��[nHm�oY�
b�Kt#*#5]u�T�+K�WR��&�&�D��g��j�=�����;�.��<�ڃ��2��	i{ؘH��^���K0��Θ�7~WSr �f��KϒI�O�1�0LIgh�	�k� 2�zrj�bN�����L� ���=P�I�͓��xvb:S����)�BB*C�	p��\g�f	$�峍/�f	 ��u3��ٺb�6	�k2	/j��yHI�f���Ja�vٝ�/��]�h%�]�FGA�*�A)3� H��D�m�i��I-����3�GCv��u$���U��L��Y��A��N7��S���wF�;���&�w��͑��ڃ=<�)�0߿;�l�����;��;߯.�߯67�{}�������QZR� hEZTNr������x����rI9vr)�s}X�d$�>��\F=n�ճjo?F�$��e��$��:�e���D�H4�c���MU+�b���P���Ƶ6�W%Va�ٌ.l�9���2]|K�'I��d��ܤ��Ȅ�^�3b��� $�IwWH�K�F=2�`����e;R���H�Φ�%*�n�2!؆r�ɐ�ʉ2��E(<��T��D��۔���H�V��J)&=������[[/��/C�\�<�0d�h&h�i���J��O��!c�����I%M{Mϒ^[=�&R���.��3�O؇�|��Q�y$�[�"Q($�Ol���$5=���7�v���f�$�ݴ�L8�[3�)?�A��N�Mp�M���9���c_����Im�m�Pd�H+��L�����$||}]�Y�$�*�C�x˱<≟q�4�c��謵{�Y��Ɉ97k�oX�۳�����Q|;��T>�t���ͼxca�f�|F"Jc�}:w�:w[ӺN����_�Wj�3�f���L����l�f��En��pM�t�,����%Զ��v+�r����7�6ᙲ�[B�7�f�ff$��.l�`.bmH37b�����r�M+E��q)0��Wl���сH<�b#YJ�XLLl�6v�R�+��o����`�j�j���F�]Mu�A��	 n��r�r\.sv(��r����-�v6	m�+FR.3ͷ]�ˋ3����aW�Տ-A�٦���l���ԭtF-��5�4�^�32]Q�&RK�%���%�w���e�{'|��a�QA$پ�	��7�ۚK�;"��f{�
NNL�@*�;F�N�H����t4I�́��K��K�Iy+F95�;Z�/����݌�Kr�$�	 ����BD�<EGu(w��H���>��M�K̟�^RM���e�`���Uy3G[m���5ϙa�6��$���L��^����^H�Ζ}�ѳW|�w����O��$��Ԉ8�La��3�I�-qyّ	y%�nKO�Gl�U��՘/Y�4^��U[�"U��a��%�"R�Ζ��Y4�1O��U<�}�B��然��4���Żes4��7$��	���Yj�P����c �'�d�������>�Q7�&PI��dL$^KVt�HIE	�ӑ�Fz��Zb6|$	O��2B��K�y���9%s"�ك�
^@\�X�$�����>�K��A{x�2�&�0�K��LZ���^i���(�-�oW��$:f�����*�x9��7�zz����U��t,k>��z�qysB������ZF��[޼��>5���q�yIy ���i�W�O��3�
�������-�l2��~�Ə���	$W��)�E2�V�N���Z�	,Y/)��Ζ�JB��u��Er��'�f"v�����*[	�p��@9|���o"�K[��e$K��Bl{7[��c{���͝��s�y�$��nZ4u��H$�U=�&Q����i���.��I:��y$K��ZD�'g���o?|������!`�Pt.%��L��saغ���[aQ�(.YP�=H\�����~J~��'t�<t��t$Ib얙I"W�{$I9��ۍ����gEԼ�I�}->��ZL��f��Қ��.���Z���b�	-�7�!��- J�32Aw\ȟJ)%$b*��8���rp7�9@![�݃�
��ٶ��fI���[�,�J|��|F�U�=��/�(���"㋗��Ȟ��r��K}�W�⳥9���qfnj���<��f���6�YI&�z�Ĺt�YP�q�Sm��=Z�m��@�B)B�4"�#J�дҪR�Ї|��o�H,n�i���߮4̥�]���w|)�I�L�t-���?��wi��I89M�A&R^��$�Ij~�q����lqT�u٭>�	$��:���d�;��a+�z1!%丽�93��c�j�<�[MKI$��~8% PIr~�y�VOQB���;�Z��!e$2l撱�k[n3��FaJ�C
�y�X	�(6�������u�V�.�3G[H�JJ���JI%��%�-}��Έ=��;>SA2If=r�)
�A��ǰ�A�o��vt$�rE����1��I ��z�3��;@���&�e�s5�� Ֆ)��R�$ӧ4�pC?�v����)�%�$�����P	��E"�&�������2A$�����	.O�/!$ވ� �f%;�. ��mc�3YO���2Bk�N�,����+Ԟ�^BI$�_KǏ��K�eA�t���F��?|�U5{D��'�ot{c�rmG�������&���{�������@�����[�&/	=Ǯ�4�>ܧ�`�,@Ы@� ��ȭ �*YW�=��zۋ���ߖ����ػ�=ݨ9�M¯$I��� =��`͹�i%���>I�����I �_K�A����b�'^�v�9wt�4�-��!�euqf+�� M�Հ�L�
�Տg4�����.�2v�x�H��LJI%��à�'���M>z��6	�kc�sy*}��e$)td����=����P��Mo�c����Gfy㼒Ib��y�K� �_K����	��n�/;�"����ok�/O�U�
�gbJw�T��l��H���^}-�i��M�m��~����y�$�KVF�ϫ�ē���){i�)���A���$zkE�lԉ
���G�3�����IK���BH$���uj��nʀ�d�e�2��NS�G3�ك�
\����)g��$o�f%��ʨ�sػ���$5W\���A+̗�H(��Kz��J ��b�&�,@�L${2�w����L���n��ڝ�N�nt��qP��˖(3�ʞlض{v�5a�g��.���3/��&�G��P�su��$�桘�o&$� ��� ��H� � �
1;�Iz�_���~\���M��yM�6LK��uX�Bd��l����L�I����ƒ�HL�rև:�K6�n#1�Ћ�5�.�bI�{6ԍ�e�,�e[1.a�i��\�i����X2��hM&��1�Fm45��f���]	���
m�eT�t����-�u1�.M4%�3K\�f�XFP�wB�c,\�0�s�n�����5&�ХC&��)y��lEi��Mf	YlF�]��F�ԍ\�_?~����\�.����x�}���$������2,As�<�O�C3d��^��yI � ����W_�rɝ8ws&R1Ӓ"W�{<�L�O��|�5s!/$J
���RA%件�	����N�Mp'�������㍈�`Y��U$���(���=}sI"�-M3��n���K�%�QA"{��}){���XT�;S9$�7�U9|,�f,Gwn��Fq�R$���HI��(엛�4��2Itv<�j�g3��gj�	���J^�IQ~ȟBj-QM�&cb.g��7RKb��RH�ok}(J��^|��Nqh"�1�F�$�� �cv��aub՗;��kZ2�k\f���C:wtf�'K1,���\���?zR3kk^	���v��Z�/�vޒ�y�F ~'���w���x�i6Sݿ;���$���zB�j;,�����Ҷ��P����0
�塏��p3�+����K����ޓuo��̻ۮ�!AbEJE)T�E��E��.�������<�O'<�̗�Q���I���>��j��~����#}�v.�ó�$������0fA&/{	�J0�V&��9ɡ��	 ����yG��%�z���ӑ��v`Y��I+�]{�TRx���32Gf�DI �������$%ϒ�j'ky��r�IA$��x3>��°����Y�Q���T���IFW^��Wh$��n�s���30u2�D���-�I��O>�y���ZU�4��X1�Qs�M�t�)2��ō̭��R]�e��J\��O���O�ŝ��#3�1$����I��t��	��8#���?��y�	-O�/)<Q`y�f,霆
W4�4o36���W�к�M�F�l�%�I
O�/�JI$�zQIB�]-�;�O��i8�������SM����ǿ������Z�e�JI ��y�ޟ?����z}���g����g����Ƿ�O��Z�;���Rٞ�{[�8�dx�Үm{�S�����{f@Ύ�4����zn�/x����Sm�wz�⟎J4ٹ���=�T7	2��o��^�R��3ޣ��vM;�.��_`���G�Ν�k���9�{N=��4�ڣ}�kG<�u�����į���W����3�ޕo��5��/������;lK�o�{<�!~o�=�gb��t�ڪ�=�s�.J�:�m:e:�QA�;� ����]�aec����ε^���/�m	\=��Y�^��e�c�݌CP}_;��Ԩ��;}w���AX�����t���� �����Ϯ{|6���=�r^Z>�[�t��~T{����O{=�h:Z�o�T�^[||�)v��?ypv�>��Z��x��;U��o����龛y�;�c<�����uP��x=|��iZ�ddx�k�'�ۤD��;������K�C���LkE<��v���uS�A���}��s�N�dӲ6v�U�##`��B��X��K5�f�*���ݏ��3���i���Y>�$�{�p?"��3��QRZ�������)��W���v�m�wh��rjY��})�=ܡ��>Eb�:e��ƶ�Ee�5�����I{Ȋq��d���=�nL�������(��`�DDr$���TWq{'e�K�v�=����Z��7��G��Rd��1d��K5ɇ<X�9N�����ۤT}	<0c��{O_w,��
 �.x��;��}�Μ��,���yƀ�_��5�_&��;`�>c�3�!�?}G�9�ș����DA�%�!��U�Q�^�=:]�o��F���wy�5�Q�E�lF��D��X�2nnb�r#	����W��\?���E�7�u���5\�%\���Y-HD�}v�)6��[�~}�%;�͌~;�b+�5�$�cEL�(�.c%}Mv���V�L�-p��b�u�w��]W���,h�-r��c_�s��=�60E3�[�h���n�A˗7��k���h�ݮo*.mͷ5˳b�p��"mr���W ��n\��}|���Tc��nm�K��o�PlRŒ�&,��X���d�����WH6�PRHt�? )B� �(���JA"I�x�#��-y/?y"W�O�/)$�����JYb�{d�]Ӈg0��9�/�:l1��3$�Zr�&I��I�O��O��ͅ�XyY���9���{ ����ub�3t�L�J��/:�	���ۗ�g�J�K�I$����QI$��^D�����ĸ�Ͷ,�9%2%~���5�4�+p�X)��K�4�E���EBfrJ`��bdf,c���K3�I�
�GL�I%lk�j�Hy$~�y��0�c�T��{7�W{/!"PVے��+��Iܐ�ŋ;L�b;��aܔZt=D����I$5���RI-�=�M$��S>&���/���>y%^�� ��S�r*z�Ƒ)�/׳JI�kr=I�jz}{H���%�J$����y�������SM����,w������	�I)w[H�J����My$��>>>l�:��r$`�]n�swQ(KmKEt{�=��������i�V��n�R=u�l���'+*p��h���};Qq9p"]C)XS��LT�8��F����Z�Q�` R`������fu��kny��o��q;t����F��bPH���Ùlܧ��#���\cD���A �^�B����L9.�[�c�*|	�%2jggJ�&�3Y�)���)(�����r��\fSR#Q�L;N�m�� Y��O͓MR$�v�I$���%�k��0�װ��s�����Q@$�{�y�t�c�pK3�I�'ˋ�́	$ߣ�nq�)��Iy$��I�$���%��/%'K�͞�FS�Nx�4��f�-��6�������U��
��#յ��ڪݬ$�Z�#�IВ�.����)�(jdRvv<�����t�(�Ou�"M��Ĥ�C��J�)��Q�T���-
��%�������x�gE��v�,~����^	g6J�4zm�]�L�]��^欦�I�+�����Io>ʙG��͂���?3�aδE_����e�EU�#�.[�<����u6z��z� �{Z4��j���Ĉ�T4�(ef+��Dȶ�z�b���98Q�H����Z)�I�H�BBC�t��$8����R������;���InE,H�kI] ��[`h���f� �eڷ�� �4�A�pD1.Э�[P���:�%�C��j���(+��pˠG[V]6΄\�,����к\]0DԵ�dI�΀�Gl�ٶ\��U�:��f�at5p�c5M�R�:���]-��%K.$밳�3���$DP�Յ�ՙ�{;mj�;5�1�X]Sf�B�Չ�nVfiI�Y�TF��:��mu&mwT����߶���wN��'U��<������JI��S)CiA=z32T�ݴ�($�dd�4=�x�ld���uB�7<ґ)^f�ФJg^��V�E��HR��^y�Io>ҟ	E�[���t�w9�M�����UN� �,��0W��������JۺZ��@*�l\�I=j���	&�=�rH$�7l��S�"�'p]2��]ߒu=�ȷb���:Kys&�;��3��D��I�KZ;oJ1c��'�(%6�a��D[�P�dRN�R��v6JU�f�\�u�.1�U��Ԕ�N�H	�5��Q^H����J�֔��9����ĭ�\̭ٱ�h`��Rk.�:Ħ��c�&���B�P��}������l�����ѩ�d:^H�[��e$K[�I���:˭и!�^ܼ���F���^oX�|L���d�Ӛ4�)ʟ<�$����n�,���Źƶ�9M�(Ҡ�I֓�y�m��(�{Z�1�����=�C������SN�"i������"$�hvf@���2�8 �(&-B��>m<0�C]��$�?���bڊ�f�Y�&�Z$iR��<��������;�_9�y��0$�_7Ӎ2�4���c&9�o?y$9�-�����.�U-g�i��RT�vC�	%�vr��LC.���В��>G2Ze:�q�J^�4a�&A�X3�H�ţa j�m��j��ω:�/$˲�Fi�X���-5nʦ4c�Q<�Y��)	�Ƒfӻ��Eݮ�'[]!�$M���|�r�rc�F��ϖ�L��,�h&R�ѐ�e�/slCtܧ4��L].t#��X]`@�l������viLuc\hėd�ݚ�ZY�����}�k�i�Ir���yI�.���$�v��R^Q��(1��%4��|��I�;���	&gv,�T��Tϡݧ��#�Y��|���	,k�i��Hr��y	 ��bݍL�Y30׻��x3�E�0K��.�9� %�v�<��H���ÙI$��'VZ5��w��	[Z�%>h��v.b�!���c��������%�c��Tz����.���Z�"K�[<��s���o�V� �"�BeH�(RJO:��w�Y���m���O��/�%�$l!�ago31%�
�%�仺ۇ�x*,װ3/%
;�<����KGC�>I ���������	%-��2�݄T5d�p��Z^vdI"O_K̦�9��ĵx���|�X��!"P����� 	���%:�_5���5v��/�p���&�E��#�.�):��F�ĳ"�vZ�46(�Z�.�g����o͑��]���'S��!�y$��0�� �I��-2��^'�eo-6eGCh����̗�C���\Y����*i�i�J�)��P���'r��c�	$^����䗒@p[�Z	���;������3��s��hb��K������I,W��)$�˛���a}�Oy$9=����Ak_KH��AӁ�ӗN�ɕ�njۏ&�����a	�ꎙI�����D�A%䐦얙	$����<}�߯���YnlN�d��<-�l�T�A�+��j����M����b��yt�0���'5̌��ڋ��
sAs�s�fa�o7��@����$x�詛�T�ib�-��@.n��$�{�Pⴳ��d��~L�j! �JW���z�oHu7�I �%�$�F�brI��֐%Jy��ڿ[��m�-*��M��Ż@��1��V�q�mm�C1����ZO_���}����)��%��؜�I$�7N����S�1��Ol�Ĥ�/,l���~�m�ɊE��Iu���&�i�)o��E�`��I,l���K�kGkL���v�l�'�ܤ�^� �J�\�GY3f���QK[�@��I)QY/+�$��ub��
73pM��9@�IK�;Z})G�ȴ>D&�J�O����?p����n��R�S�`_����Z� $�G�zb�����nJ%9oS��P�,场d�M���S���:/��j����{.[I�� �IOLa�D�>�Ĥ||}��f˶)����wR֠C�{���MR����Z�ڣa_��5D.��\3���H^��>^@�����1��8��ۍ����v�6�ڣ>/�Vd��U%e*��(К��>��w�\��&�$e��Y��u�3jK�s`�e(Gl�#1,�.�W��n0���iMt�r(*�/Z5c�ݶ�W���Һ�( SL�+��C1m.�9���]3*K�aR�pQ��(�!1�l$6:�L&*)���^K[LI�e���̩��ذ��6��*��!�QZR��P�1�2@�Lع��Ɍet���bե2"�,cK�+��L��j��ˑY+x��LJ�|���Ҹ���b���f�P!���J_O��	$��j��P9L<�K����B���W�fR��4�t�bfBQ�#Ґ	X高�#%�\)հ�%OLY��H$|u��%)�3 �#c��^'�Ng��=DۺdE��Q��i�@R�K�g��lЗ�3$�T�� Nr�I �K�D�y��%%��A3PA�̙�3rK@�����ȔOF��9��Jzd)K�� wff	$�O5򆲹�e�9ޛym��H���yJY^$;�g2v!�L�5���e �	b�Q�Zxu���r�ɨ�3��/#�	�����P!S��E��<+�w�(Q.��&dK�i�\�:�`��u��[MX�"�K��s,1�g��z���3�L���Jq޹JI$;#�E���%�ڢSb���?b��
c���@�5���|�aVY���s"q3t���G��٥�N�ύ���<���X�_n��1X�Ǹ:�׊Y�N�?o� 	(٣�I� ���p��0{�U����Eg���x�5%D�Hĥ���~��fV7~F�W��7��(�	'|N�v����9�(��('r��!O[3)��z��	\�3��	�J��y%䗏\t����|��3�s�~�i�:	�&N�6�U>��v˪�Y:u���516)��/$��TL���j�v|�yU
���%(�A�b�39tKC��Q
��%]/3�-wm�h]t=cn�Hؙ�H�x�����Kz#OŲ�b��`1�A%��,P,��15Lj�F,�ͅ�D�Km��U�բ)4��<�~��|��ԦwE�8�ۘ�	I"qv'0��KzHHUZ�=��sOv����e%�M����E��L��>�WM�J���M�W��Ϯ:���%$�J۱Dy%�[�d	]�S�w��0���Ի!)r	f!�Ț������I"���R�IMM��U�w�~v�uNy�D;��-q�_��~?Ұ`"{7��IB��u�ٯ�^��P׶�fv�w����c3:�տ���y��;����C׈#��G�����GܠB)%���dJB��!�9)�X���=t�n�g4��S|I)W�%�ʇ�������<Cݤ�w�\�*=
�}��V9v	�&N�V����x$:�"}+rpE8�r�Y�U�|�آ I${!�ϥ @I#�1)N�=�.-���^N�M�Xi�(<5�.r�Z°e�&Kr��Ƀ(7;�dQ:������%��+i��A,�|�)A"QΎ�����	+�+,n��	?`�����%��q�Y�����|���^I{Θ�I�\$�	 '�0̅�dt��I'4����}Ζ��� ;�N]2s&R鷩
P	$�ttH��"�.C5�����m�I����H�GLJS��'K3�hU�n���/n; �	 �D��RJI��H��b>/7m�zh�v�xioK;��"n\Ld�VTǚ�[���Z�4*����x�nǄ4:5]��*���^\Q��x/��l��x�x|@ ��| ��Kw�H*{�0~�?R݁H���A���e���r͛u,�l�����2<�I�0L�$����ێ�����ג~�CJ��m7ip�V���(C]��Q�6�b$m�aGk�-���{��6b�L�����b�I
�șD�^I��@I�6�q&f������H�ىJ`"yg��39tKCϗ4�	 ��H�=��cSKĩA%���2`�AI$7b�E%/u#o%��l��� ޗL�A��v�#�&0JA%�v(���(����� �˃D� o�f%$����آ�;a!��r铙$�[���n��H�ӷ%��aoz�^H��0ȍ�ŷY����R@��LJHuNq��$�O��g835ʁ�<��?��7y�-���<�3I[� �IK�#H%bL����������돏�����z�~�h��R��G�>u뽜Q77��/�6�����Ε\�����x�I�'��:�zL�^�3\�+w�M̑�I�I�AT>dzzD��aŗh4�j��{��ު�,��.�uG����~O��s5��ɨe��g���_b�Oi���7��~^��ޚ��g;���E��{�6��	y���mg�S��L�vw��0:�b��z8|���=�WK�~{�Bݾt��ۊ�y�_����8
t`,��y�&�/�&����{Gjo��D�Q�����C;�ޓ`tu�oDϟ� :>o�D�Vo�>�{�8�b,������[�~�o�gQ�w��<{���1���w=_Ξ�4�پ��9��}�lD�� �����Jg�{��&��=��}v�l�}�Ϭ˞�W����vh���;�2]�v���\�y���f=��2O�������Q����K�����~ǧ��x�DbQ�N���Nwtx�d�3��b��=����*����sx�'S�}��vOy�߆-Q���Ԟ�����R�|��
vUA��
J��yx���/��Z��z��<���m]׶��;\��I�!��G��W���j���z�-U��7�,�Y����������{��c�������lԠ�Xw��6b�\#�
K��kTj��J�P�:'�t�-w�G������P�ކ�e��wޛ���ȸ�s�\�P����yڮ�/�.ƌ3������[�����5q�U�ս�7^'w�xf�qr.8u�c]� �r`�2�&���H�L��
C�|�I���z�aI���Sb�^���Sֲ��K����F6ŢŢ��Fw[����E�����o���g�p�F�ﮤ�cY4i#�XƱ�m�!M���r�1%��bM�m���"KFŽ�nr(�F&k�0����h�ל�E_;��j�巗M�ۙ��QQ��tہ���ӱ�ؤ�4	��l[��o5\���nA�6���s���4o��,�o�nQU�)�#Q��m�I���r#hɺw��Kp�c}.xWw6�of�>��k���b��p��f!�MY�Bak��\n�\L%�9�ͭ�K+j�N�M�\�e	Q���.�Z�;KkW1�N��\,)j8��CM��E�iV����sĲgEM)1�7m�5b5&�\��؃tJ�\�b����.&lm,���2�����1J�@�iU+�(1�ia�-��D!�����*jJ�&.���"Q���&��a�vBk�9j��5c
���Q�&�U6�VYM�[aU[�S#IJc����,^�[/!����0��={��Cl0Y�����[�P�g��)Ja �,��ZW��e.r͕��`�#5���L��rv�к��1E��q5f�J��<m�֬!y3�%�%�f�faD�����aa����1�l��%6rU��!����a��wam����ͩe��,ل���w��\�l�mh=��k���L-Q��,ȓU,�������L�ąn�ȁ�f&f��L�Ilб&as�΁4r�A+Ib�ZR]X#�ݘ��+��*,���Y]�	յ�fB�W��֦<<�����%,Fd�'c9��iq�i��Z��4�SV�e+,�:cV�r���!q]c�bh]�m����ip�#1�l��є-�{g�v�;����ڻA��lT�ke�1az�l	L�F	ma����6c.��Ku�=`X)���dc*]6�\�Ha(i]H��42�l���s�+%��A�e,[l�A\��)�Xn���@3��k��H�wf%�Mq*P���ue�bh�a!h3s+40��� ͘	���3	tQ����Иhٹ�9�]�����tvB��	�ڷ�&iu�9� @�ʹ�asͲ�"��*��Zch�m�A�	\���IBe�Њ"]Kh4����p��]�n�YQ�k3� �B���:�
;B��JG�%���B�a"�S� h�F�yY�UW�i����o<u�.UW��]��{���ߕ��_/<�C�5�f��V�KkH�k[0��hƃ4\T���QԛvL����<���\1VݬB���vm!���L�� :]t��\P�:���Ya ���Y��ƃM��+Hn\�PdŎ�^��Vf�0��X풭#�鮚�a�C�G���X���R:,�%Ѳk31dU���%*�����.�pG9�M�T�^Q���U������IUV5�c�K��{K�)-��u����3�"h�m,m����?o�3� ���@\CM�~�RH�Y�! A%��e*꽡��95�8��}ꈴ�^T��<!?����w`��3�M_����JH_�?��ѭ�a�tG	D����QH����D��`n���ܘL���\	5A���fb��-@?.i��f	e�̀���3
�&:�C���w��"W�6�r`$���4̠���r�"�݋�Uyɩ�s�"�5Q�뤒�ܜ�Iy$;"4̄��^8��3N1�i��I�4��,`;:.�2s&@K&ތHU�fA��$J������:J�~Q	 J.cL(�<���i͔	�y2���A�,�Jvt���,v�M�Β�P�<Ss�l�tÂ��R#V�f~�?��c3�xo&h��I�%�T�%��1>I`�	��٬�;Ai�M<��(�ژ�"R����N����uU��D���ې:�p�UN5��!ˎ�H�Ag��Lm˴1�6N���׽|�����8��.w�?�]�mB14���YT͠�t���3N��| B���I$^��3)$�����_���^�-�o���\$3�Q6̙�2b�n�}��	�p���}��y%�p�Nޑ�U$$	 �f0�2�8���!���fb��-/+�i^BP"9�R�l���3��0Iy$s����	 ���J6����2I����Ro\a�; �b��������ʯ0fIb~Nh��5�'��<�踲��I$ddĀ�	%�|����d�(b����66�B:��m5�J�e,�F��-%Q����m�������1��?N�J��HIy!Y�I$����0��՜�DN�̘� J$�w1)/o�����,��sb�&h�ޏC$�"���8�l�WF�ϔ��� ��LHI$�־O�(��s��\mVK6Y���}NXd��Pp�+� �s3)��帣ЉA?�x��Vv�؃�G�(l���T�s��y-b�uM�,������g���B����E�ݞ/$���ԡ�2�:�q""�+e��� ��z;a%䑾��%"K��Q�
��Lɝ�LS;<������f��S���3
h��J��\��הy�̟ʺ�)�*��&�pJH
�s���0v$�
�˩d$�@*�|1ro�xM���>V�^��)%mڜ�`.�3*�zVE��I%�B�5v�0�<`���"]�"��讠�rՃz�[�P��~-�V��,���!=�?#��RX�B^�K�/wDa�q��K�gn{y��v"�A$���zݓ�HP�'�2s&BQ\�>R� �8ٛ�2����9�c=(�7�ֻS�[�E����4�>U�Q�԰�����sщ/_i�u0f�
!�܃v�R�I#�
����Ie���	�0��.1 I.m�I~|2��p7(�_��I��XŨ]���@B{P'�̓y&���2����ޞ�>>>|m2^��1�h�(Bg��ǳ��/�.�}���E|	�D�|0�AM��Л�|/�M%�@�Gג33�Ô���kHښUI��>x�K�P!!��gP��S:I�d�w~Jޟ��H}��2�m�^(M��z��@,g�Iz|3(��lt�#[9�)���V��A��t�֘���GLKn��5`�:��a@.p�����Y��%��kM��H%/ϒ���::b|��s�~Q���{�Q�i�^I.|�3)z�"���`��T�˘2[W:��GSܮ���	 ��?��H��LJK�kD�y1ۦ�VO0��o��j8t铘A���D�5�� �I��$ar�;T}�:�=U]$�|�+�{_�L�B+3X"�(Q]slf�ݺ�G��#��#ȓ�n�6d�Gu�Y���uV�������E�A�:��["A ���ɻL���[���f	&o#fA$���Ơ�כ�#S/�N9K�jƍu�~��&�������秎�ޚX}�����ᣐ�;�,�/���7O�.#���\��8w�Zͭ��������m�dM�d�Y�Y�_
Rb���A�h�u�E����h�Չe�*�e��:CMA�Z\ib��GYMVՋ��*j��G�z�fsf5��9�ca��qIv̆�Q��TÂ��5��\M��e�i��@7g2��p�.J�l���1���k��Ю2U%hƐ��^�&2�a�"MiT��,̳8"�й��j�s6�n�T�t���$�>I�[Ċ�Skx�.I�Tƺ�Z.��X�h8�ʵ\]K����>
A�m�m��"��dH ���؂bF5��3ou�τG���O�LQ�LJf,�ؒ�%�v_�swȇ73c��Ak�jgĒ޼���B��e&�"��YefvE.��U��>$�{o G���Fnb"���WC?Y���x=�`�k�Az}d�l����Cp��';������Xl*��'wtk:z$ �s�" �-����xmk��&.�f|H6
G� B.�}�a��皹�<�v�PX�Q��Zx�ȟ	 �^�WsY��r�֎�޸�K���Ղ��,�0�kα�����DҦ���n�0�\�:L2E�xE�Ppη��.d�@=w� ����`˔�,:s06��d�Aξ�N=�ę$�ɘ3'x^-\��x�*������Pe��!b��g1x��`3Ӆ/�ll	����2^.�5r�Ӓ͛���3��xn�^rk0Z+��۽ ����>+�k1�O�y�N��͗���f`S1fĖ�$���I]M��	�y;�˴����A>��=+���*n����]�;D�Vu��>�;�GB�桪��O\ļKM���}]�2���Ի*)f��I��g�~~����çfNc�t�B$���@v�����a/y�Y����|O�"�dd�&�9S�4(��Z�ϙ'o�)��er��
��J�p���Gk[4��4i[��}�J̴��;�nz$8�H3��me�'2=��^����]t@ �|�`�5���'�A�:�v�'�ghSI6Gv3{M[��^%���@'�[�2I�.�ř��/�-Ku ��v���ܦ,��gSV���Y�1 �H��TRw��LF�q�)�1��ˉ�a��l�*$���o/p$�����)kNn֓N�����oLh-����{�ص1�����bC�N)�u&T�R��O�d)����� 6��gĽLifA&b��-#�:um��;x�K�� ��M����Ao?fl�Cs8��b��ǁ"��l��A��i����A ��oB|�v-#=�pKv� `	[� IǺ�"뮋�m0�>>Z�q���[H��b�0�k�X��75�=M-�������
�pW]5Wq��ע���mL&�8�j���혒I�$;�" 0#�FBv��w����ǉ;:bA6IC* �;�
�-�D�><:,+�Y�x�H�Ι�A�n����|k��y��c���4�[$k�g��d� �@�;$zA쾈�I��֝L�]�e��$y�32	�����µ);�Lɋ�ϏS�Ž5�\�h�3)͋9ћ3�&�� �N�+��fx.�w£K�?/o�ڽ�`����I���G��M�-/�(i�� J\�j����G���n%��b�M�FSg��"��dH<�W!�f.�Y�h`���5������tێ	�1Y2>97� Gs�����ǳ��ք���,�#ec��f�MA�ZU�uՌ1ײ��n\�ֺ݌E�s~|��/�&G�w��rd	 FvD����9{77�tΡ/q��!O���^��F��A݋�fs@P�ڡ���6jZ��Y�͋�$���#��ȀSC�����B��s���@���P�w�]7�y������6k�c:�H$�����h_Xr�2	��p΢�~�ʶ�k�� ��@�H*��~A��2�՜��Հ�~��{'�r���̃;̂�W@c�|w�&�vW��ue����x�$�+n� ��t̂��tF�����}~z/�,��ka1
l���ŗKP�:Ӗ.F��lTÙ�VFe4χ�ݎ�\�ر��v���ȶ�����w^��ɉF��
I�C�ML�i��ࢄ,����K��y��܃ -͹�N���!�k*��bA�.�V0���]�ד8�sj�n��U��(Ƒڛ��W��e���J�ب��t-�����V���X\gM!]�i2�#�	���CkD �6°�0�����ù�E��hc$]���b�Ѧ ���&G�F��eK3���@��M�tm	�xn�VG,�0.�^Z[��e��Ֆ����8�`5u�vq�·sK�ȳg,Ķ�1�� ��nCO�7�d�`���Z�h���ĩj����H�2��݋��މɒK0����ة�0���]��7��4H/��CfVFGt�G?�Rr�]�3��P���A ר�L	%yv�	wa5d��[$	\�� � ��~�)��F�T�w$n�^mY����#řD�bI�/���	��ʆ�Y��f���N(�� _�b�$;w\�|@��=�2�;9��S�b��d̓�L�tz���7~�8!�����l�]Lu�L䙕��f���c��0�f�(GX�]������n�������mUp�	�ܘ�AOw@���컬gx��˩G��
��c�nj4�,1wr������@���m��ӾB,�esܟ��?�(�7ֆRh}����3ҳ��w�u��q�h�#�������KB�Z>1���4��]?\)��=��<�23�kz"�����g���ZH��H�~/�,읦F��H�^5�� ��E��\T���*Y��	+6`I>3��NI7l[�˱wfg7f�uL
.NR=Ϲ�K�D�Y���� ��d��ؾ[O���'��QU�>�\���L���(P6�P ���M�Fn�/�]��KVUț�@����ـJ���'���DdJ��y5�j�lh&�beꬲ��l�Zhf4�kV�..j�I%���N{���̒H3�� ���f�8��6��z����]Th ��f��e��\���3&.�F[�`"f�vl>6����vol�3���D	�� �����z�|��ub��7	����fd��0-���QpA kl� A��������˧ON�\||||||x||}�}�w�̇�{�ͥy�[�jGk]��#7�/xew��{97��Υa=��/*�����x2����rX�y�}�>7ݽ^X�d��'Tܻ�2<=}gQ�?`�5�U���q0f�M�K��P��ފ7���v�;���7h��ݍ�6�h���Y_����]'M���Grǧ0J[=��1����~͗9 <����|C�\]7�h�����ȱk���Aϼލ�7і�U����V�}=��{|��wD�=�#�������~^kv�m�<Ff�@�cC���l�����g��;ܴ�x᫜��������kQ���'i����/���s���7�I��w��}����m�z��������F.V{~���_h0q����?3����ӔI�������/�ـo�zLN�`}���xj�p�y(��^��DKf�h�ދ����ﯺ{���;{G��]�	�d��G��u/7���P7�[��p��8n/t�F�卑~zB9����1����֎<�Oi�u	v �|=����o��1�}�]�����i�Gg�q����"K���aC9�3^q�ᯆ^���G8���
B��m�ӻ���0��F����g������y؎��=�$�4�8Z=�r��9x��,�sm��Y�)��9l�P������h��'o]�>Pyo`�g����Ϸ�6�|0p.��&j��ޗ~o�����tSٵ�O,Y���Zp��ف�����w0�@�mi�y�gx�&�gG�]��!�C�U����A�ȥ�<Ť��9\��F
>9�wr�Q;�W+�ӗwX�w�:�W{�yd��W�v�r�ݽ;�=�b�s\�MȻݼ�u����6**6�u�scss���*(����{6�&�X��b3����W9˥���c%�sgq����sF��.k�_;��ۥ&+��71�ᢈ��ms����e9��4�WJ,��[����-�iݵͯ5�wW4#;��p���X��aݍ=�k�k	�Z��k�ݢ��ѷ���X�����涪���'+v ��Y��@��?���v�n���3�4��׉=q ���V��`�k;�#�P|I��{����p�ػ�3��M]=@]�5����r�%[(nyv:ل��$�mo�	�5��2i=�L��t� �X*��Hb]MP雃�ٶF9v��i�v�\+M#�ԃ�N��5`"��ˀ>N��*= H[�`|O�ot���eŚ��=@��<��"��n�I!�\��[��/ă"2�VRK��&���D�-�Ј$��{�w~!�j軦1*{p[���I2p��3�I���� �w;&$E�7�T6��l��	$��D����ss����'w)�j�L�x�b����i �n��$��əv�����:�࡝а�)ay.YJ���MM�E���y��x^w�=C�s���rӖ�"��]�ں���&ky;8r�M1���M�%��b����Ǣ"�� Wy��Y�;N7F@�	9]�!S+��q�b����S���/snD�z��5����V5>��Q\��aL��Bg[t��&I��
�;��3݆�ųש���\]s���?;��-F =�nDē�A=]� �#����p�>�׳ �U�0���Y�x��H��� ���[����=�2�H�^F̀O� �w@�ڈn;<)L��{�C$D��r���>�l�$�U�A$�]5�Y՜x�G˲:dA �wDrAy�\K���L��}aO6�uH�~T:�v��{q!���7[����Kі�j��bFvoL�}�S����'w)�i�D�A$����[�Abn�G=�2�Y3�A>7ב��`���2x[������o/II".h�e\�Ȍ������nf���)��@�R�ݷ�lỷo��հ�S���R�~}*���)�_5g���#k�Q8�-6�n���q��9c]�&0ݕvf�V��yf��i-���i�����J�&��J�<�+nN3T�E�8lR�]�K��� �l���"��wmuʌf�ؙK)I�f���&kz��-��c��`b�v�A�Z��C�QZ
�R�vu���a^�R-�����c��[]�]F�)��B:�8Ɓ�Y6
�Y�vb�HV���Dtil1rE�Uʹ6!a��tKu�Pҭ�&�1��2ЫH��'A]��r��ڽ��cb�I ��Ȃ	�+y�����1���j/���|H>���gݹ���4�I3oÿ���|����ǸiZp�l�WEx�N�����`o��F�"Dm��>�h:̯Ė.�D��0 �T�l"	-�rx[�6s�=�y����؀@$.��m�L�i�I�L���y3�:�I[}�SM�O�S ۽S)��!
�z�<4�^��
ͥ��	������J�m"<gd���1�Dј^$oFD|H��� �g��X��v�{�v)w~���B�%���i�q<n�X	E��ː1S,,��w)�B�3V��l�}}���b�;�N
�;���M�$������~/i� EI��� ����D ޸�h%�O�,읪��vgĀ@�eve�����߽�?���~��/�I;؋'��۶�ʀ�;�pZG�X�&	��x�J�9���w�O�/�q�5��YN�*f�\�_C#�\��H��c�	��s���DI8=��h�쁺iN�;�LΦAۦ��^$쉉��U�[�p����읂-���/���D���p:̳Ėt�Ex����R��,f<��� �����7�y���ٙ�$��_Z�7��7����CyJv� km�L�i$I�7�c��dZD�k�4`��-~�@%C�]v̉ ��{2t>�+�y��<�I�"��ѝ��0,�Vj[5v6�b��k��"���ן����qTŝ���mیٹ1$��'�בP��()a�O�z�d�����0L�8J'Ǣv �����26�T�!x�f̉$�^?�[�[0x�x8k�<[hS���坒x�ל��u�A�$��YkY��~i(���5��9cd����a��q���Ǿ�vʙí��2F�cS�-ը���+���۔��ji���-CY�X[ө�f\�є}�o �ןu�I5����&��%Ӡ��ٙڇF4ɘP�XI�~��I'���o�\��S��mƴD�A�Θ�H�d8��߉,��
�U�	&y�`-������O���g�{/b�'���`޻�*�0߄���|-�R�Kt����A!Ũ�m�v�k�%-�ѣ`����V���n��ٟ�s$�^\�b	$��{!n=���m��"|	 �����Vz��E�w�3���e��uei�����*=���~�'ŀއ�> �l+ۡ��D��f�a#*�@w���R��b	'����5̨n��՘O�=�� �N����-�9gd�dg<��N�S�w3^�ޞ�$U�ـ	��L����/�����yBa��
c��-8*}p��p�M�n��.)|F�Ey?m�˵�z��!��]`�9��y"��v�u�m,�nW�Z�ڮk�3p��i�x��t����vgi��mP����YY<0��i�[?����� ��{1��7��虑��bm�Rh8�Ly�D�%��+oD&`C�Q1sJ�bZ�`fMs9!��ܤi�M/ߒ���~���t���*�� �ga��Wtt�+�]�n����������D�u�,Hj�	�/C��E���Wy�x����t6 �k�2d�{�n��>��W����A�r�fvx�4��G�n�dI ��O%�=��>@'��;��B@ޞ�8w3�p�;�N�Q=^�㨍��O	���{�2�|{�6줔�V�0��|�`�f�%�ˠ읙<�6L`��y C��Y�VH��� �H���I;׎��d8@�v�)�����<�MQ|6����s�'T���g�?>�{���vno�f>o���'{<�J�G@{�I:��������I�͡-�P�\,�4;:�Ke��$fZ��̺S&�($�#	���y����Kn&ۍ����r��p9�ua\�ڰ����"ؓGѭE�6���͓h�h���d�fj�&$k��q�iʶ� v��`#���B	��]�tΘTٷ#{j��"�bb�T�X��ɋp�l16,��ց@m�x���;�H�KI��j�鶚��ASM���!Msh4\�.`MJ���+�÷f��Tc��_>߂WQE�߿��֨�A��ؒA$�^Dx���A��O�Odt��A,�BH��$m���8`r܁�}ǡ��|�&k�bA����7��_k��*��dX������s�����5װ �L3����C�h���7�vD�Mu�S�� ��:�;�H3��q�o��f���Q$��Ou�Ay�q�V�w�/���$w���p�;�N1� ��;a/ԍ?t���yh���{f�fA���@'��L&bS�L�'4�A-~f!��+X:X�V��ɊA�X�:�S:��;itɜ�(�5&�>{lŸ;�'b�Ҷ�;��x�	�w� ��c�n<�"�I�-�]{>�u@��ȗr���3��mQ�M���}�ئG&���o�X㭥�7Vi[����ˉ�������	nn=�n��9X4�le�e�:��8�*��fe���b�8A������#Ǻ(]��U��ڱ�������@�m��'��$��|���=��)1S}�H�؀I��� m�Y�,d'Ha/�=[H.���P.���� �;�+�:'��܅Q>3�X�*ˇp�ggy�e������ؒ�:��Nu�sR��l@ۋ�$9���$;�� du�	�xx}XO���3Ӟm�1�	��,���w30�4D*���+��v�b���ߟNX�,�i�-��k��m��$�]q� �1��%Z	���}v�#[_LZS8!"����3̌n��wL��V�謸ޘ�y}�1�Is�fI;R���,h_u��{c��	�(�v$�vgi��MP�$���x������N�і5B��PY�,������}@S�����z'Oik����n��_{�I���@r�:M�k�U�Sc�!�ϑ���9��0O��}3$�9�K��gN$Hv�g+0�1�K��$��D2�fD���ܖl�=N�ݾ=�w���>�~��C!A:A�B_��H9��Ȉ�Ǟ����7���	�~>�ވ�A�ȇ�U������ǆ�Z����Zc���S2�jk�Ⱥ�n�X�;RMa[-8)��|�_ы3�?p2��?� ����$��{�w�����M���a��9Y�2	��E�;���:3 �N�����w�_Zu�KV�	�nL� ���ΑV�e^5��;��c�(2v,����H:� ��]��w�nI�$c�k�������A eH;E�tC�wfv��-"��xY�����ؐ	YY>[�Ͻ>��vv��\���?lV'I~�zI��or�CU�f5����?��g~e�oU����6����z�}F.�i*i)A�ڪ�ø���'�Au� Y�̉�|e����~���ʛ�Iͮ� ��^������-���?f'�n�����	�1������,�.�U�86�P��h��5C��s�b[>������H#2� �<��B	�w���芙�Nes¡���p�,��&�a�q#N����h�H�%�qH�n{0yy��i�����K{n�ϝ��gp��c�+`A#�� I5�1c��2_W>�$�s+\A#����L����3<�k�J����κo$]�#�A����v��xU9��t����w;�=>�k�gb�ػ�;UWMP� �ltH&�5*62�஻x �n{0�ö>w�^�͡�����ח�O�o������{=��g�����F��2ő�H�.��	F��D��*��K��B2�^f[0,�ѧ|��{���_.�+�՛����=���K��Ƿ���A�V�ͷW�A��_�];�����8���FL`b�.o%��ȅ8X:b����xK��ڝӝ�����@�n�7 �Ǐ��wO*��3|��
|��?��.�4�V������Gq˞��i>kޝ�]�Y�]��>�Y��M�������/א�������S��V��41��<�z����-��+�霞���@�������6��X������r�^��R����zN�7*Ze�0Z��웯���;�=g�Z�7��.�#�z�r�wR���{�*��W�ո'�œrM���xq*���wQ8�2�ݎ]O���\���ӳ�����a�1�P�}�B��p��c��t��d�㹯7Ŏ4��F::z�<��{^��ځ^4��y�|�־,��'ySb��\:���p Ng�������pU�E����}�mwwx����;| �e�>��/}�'`޻7gL�7^���W�λs��=��T�a#�J� `���?_kkoC������n���P�or�pmg*�{ʥ=��o|��-�nQ�\�l�>އ��uD2�]�)R�~<�t	�g���gu�yt�i���U>����œȮ������TL����M|}�e�V��A����W�L�A���O�W\����D9�U}	F��o���٬��>z���n�]\�����뻆$r��|^I�b�vif�E6Ko�۽�>/7.k�\���Q����-���.|lnr�j�.���F=�7��g:�.nwv�V���*wڝ��+�*�~}�"3۷H��9&:Y��\�F�DQd������r�'t�ƹn\��D�Q\�����AwS�㻮���v&q9�6/�E�W1gt��cnݻcg8�"�(��t�.\"%ݣ�1w\���ֹ\�f�1�wwcs���t�b9�\5�W�����~5��;�e	���FƏ9���.rh)"
"����渶�n�s3 T-#dB۝���5��5��cJ�-e��L&�V���ցB�f�b�*Sif�!ف�UI�8�jA��i�ݲ.F�:[0)�]�ZÎ-�uE;WR͕�iK)Ua#\۳��^H��Hc�6�Y��v�.�bQaZ��M�h.!��F4�c��5�b����D̶FV�۴���"�2� [�c��f �ʙ��vYaM&��ư�8-�c����8H�XQ�Zf�]�����,������f�n�g3 �!��n4,ZfQ#�K��� !R&ˁ�L�뇛%Ŕru��������K`\�f[u����`��F�5s*%v%�n�kc�2�����h[\37��܄�U�rsz�F!m堲��1�1k���F�
1�۞�n�I�m,�,،4esi�7X4[�� L�p��L��XśBlMq�J�j�Ρ�mViQ#v�(�Ѫ,뮌ΣD�ͥ궭�,)4�\vK��l\ę+�5�����6�R�T �F�0�f�.)��%�t�s���P�@ڭm5m�.�-і�����.��CX�� �nVقԀ�J	-�]�Du)B�&9�f��[u�-�)j,.F�^��R��\B����q���+�33-�ǇM�]�B���
dq�hL^"[��1l��fYV¶�SDl��Q�Z&V��m��t֤X�U�0��80�!c�j�uU�Q�9�9,<By��O�2�Ka�3g���	�J#ukZK��b�H�4�"WRԕZ66l�XC6i7kZnH�M7�u��!`��l����0�)�n�4:�K2:�kQ�զĲ��4%���Jm�Ќ���x4]����\ݴ�[� ����� هj)�A�P��ZZ�/gb�p�qB�Pm]���+3,kN�R�dt��+�R�F��ۚ9W���ֈ��S@�"�GB�.W�f��f,UW0�ɶ6vv���|�W�g���˄��va�u&a�en%L,G6L�-"i� Pxf�"����K��f��c;��v�y��B�S;3!��-���P3UZ�v��v.�X0a�2��ii� q-��k�#�O1f�9�pǁ�*�%�28M��tm�K3��kfBnE@�2�u4���F�0��J�i\]Fc6�
ی[NiL��[�� `�B�hf�2�Ύ��k�(��r�L�3�\����S`	ó����GAv��"Yݏ�YqA �si�A>���뽸�ӯ��� @>'Z�L)�[1	I)��L�GWL��z+�n�~���Ȭ��H��D���$�Sзu�%1�X�W~��ݥ[�p�.�����$ی��Kf��kyg�&-ͺ	������wc�H�̡�3��:0#�G��+p�׺ăݭ��A ��� �Ou�R�����&�q�	#�$Y�9A��fy�3r&d���{h��i_h$l�O�U>� ���$��؄���j+��ˑ�i��Ey�i��i�ii�g0�ib6d#��GX.옄��+��&.��3��=��A3O�>�{�^<bT���3���O��6�� ��� �hp�,��D���y����*�Ȕ�#�eD��馸ǻkT���<�x��Ú]$�B8��H0�W{
e'c��3k���a���~D���tI$����Ʒ7�%�WmMr7O�����%D�"��i��$����&b����7%SF;yH ��̙�����7��}֕8v�b��A��Qʠ��"�&��$��{>��$�������m�mGN`�y��#*E�E��wp��� �56�i�7�$�g�+;`O�'v��5���;��gT���;^���^"׬*�P�ܫ���6үlcE���S���ݔw`�; �V5&M�B�2g��"I;�� �N�>�+���'Y�I"�� �P����1p��;H떓`��L�ǭ�\+�z����� I�����n���f�^��j�p0�%3�@�y�"	���O�>�Ɨ�n�����a |w�쥯F9��>��������3Ӱ���cpa9�G�z^�g���4n���§/\�U3te�J';�$}}�ss�m�وJIvD;1�Q��[����1�I���$�M6>�$�:x�	11�
}GQLY�ݞd��q��|s��H׼
7Jn���1�k6�	$[S�@3��vĘ�km�� �z����+3tڎr*�+�b��t-i�u��n�)1V2��������G"Ɵx}dz�Ʀ�D3��2����a�
Ȩ��@'���c��h�̙w��ɞ';"dH=��n�'�o|�;�5[i��{��l�Z�tkC'-.��A��f�i�xS)��w�Q>�l���� ��ї�m�m�wQ�I>���H�~�K���AH��S;5
�b�Dfvky @l��y-��� �{�\yy�˛~md$��׬\�RI����L���.dŎ�M,ј,][m����#sn/�{�S�K7
�}��z�<<<��K����<����o|�>f!*%���]Fto���؆��v�y��Ջ���7� ����Gu뫵�t�
���r�?��~@�B;v6F��R��JP.t����Q��a�V:�(-�G:��O_l�o��Z��g~��z���^K�bbI#���요Z��uM���{0	�>��/���,;�vp�̂�]|\(�Zkd����ܽ���%���vD�I;װ �v�h�T�����Ȝ��-�0N̙�Y�x�㢼��lߥ	i��Q�ã1�E�F̖�^=װ �����ً�Ι�k���-�t�e�^��-S}�A �ޭ���5���n�R�%��_���8�q%�$�U���_�d��ʯЅ};�}�ל^���މ�����	�7>>���N�0ѳR�
لP\d�RМ�ȥj�$3[��8��A��=�]����8��N{xŎ�n�{��c�����;�+v��T�N��o1���*aܗ`�2��LPr�f�t�µ۶)��&q��!�D��[� �4\A��ڃ�m52���[6�ن�MJ�ʓ5Z�j�s��[Y��ݥs�d�.�\�\٪&�,s�Le�ȜU�5U�q�҅jV
֗�e��,�� J�� \Q#dif���l���(54�#&�ƴ�F�5)B&M��pf\Ƭe�t ��݅��!R͊g�I�c������]�6�{�/���,�=���fA�]�A�'[�L [7�P���y�'ă�x���K-�� �;���=�]�sz&�7�/ć�[fk���>�s���k�Y�[-��7d��ҬE�p���ãr+�	&[�a�F�49���D���}�(���<K>����r��9�*��9� ����	O6�ϒ��ޖy��φ�b$�M=��vb��',�Ӟ��
���|c`B[{���~����]�|J�}0O���@w��ycX����y�ZK�GYl�qU�5,4 �+�v��M�5�ġ��1b��Q6(aCt��$��p�WdD	+i�$�<��.��tD���;u� B�|0M7e���)�˴�L� �s���ץ�v*�� ���d)0�Sf"�-��M<�ҩS�H�} �?���=r�:����%ҩ+k�Mx���#��=����%�Ce�$���o%��d��c���3kfC�y�%��ıd��Ag��D�缉� �l���P�˳<O�Uφ>&u��K�V'�8tds�i�Xpg�-�'�4�w5x�Rg� ���n�D��{F�H��`��$�&<���fz޷��I��7�&lՙzy]�H�w�$'�2dג��"��e�ds��z`XYm
Oŕ�7� ��Vꖊ�+�[\̺0�le���2�ƙWs�׿��b�:)�;w�MP�$�� �@$o_@��Vύ�⺟�x�N��H�a�6A.N�ZD�ͱL�.�[ZfY���>'2�%zB ��}�^sr�:���2_�LU��L&���g�ח� ��@���y�J�t���*�%E�-�,���i�|Yl�9�����K(;fm���x�:v�&��I��c��{g��44��a���Wă���> ���� ǧ�`,�`�� ��TY�ld�@w�2= �_<W.�q�ף#Ld�]��dm�ݭ�w�:0*�a���!x�q[�D�g����ݙ�$ח�nC�A>�n�$Q�r��gZ���{f,X�����4n4t��íZ�Z��M�����i�T�j1Ri���z𥥎�Ȃ�Y����f|g���y$�ݪf-U=��+�j𻪹�	� ��<e���ȳ�p����u�M� {�f��3�l�]I'2���L�׳a����h�E3�����8.
N����ͯpI2���H=��u��n�kɌ���H��q ��φ	ۑ�ҙ0.�C0�v��HӦ�^x��'ǚ�	���=�"�]&hz�Q�jӶ$x����<�{����ܾ����Yvj�������+�%A�j{9^ed��9?b[����<��z���7��_.����=qB�_+�̬����$���3͉cS&d�0wg����N}q� �6�G<�R%K�w��Oo� �Uttϋsd���-6��%J�K(��n؋+4R�f����+�Y��,73,����eia=�?~?#M����ן��jl���$g:zdy�W) ��mV�3�|Dskُ/Ӵ���Ȃ�S=P�}��M;k1�;a�A�� ��׃�D��L��H��~¥���P}v:��2,�3�gh@�[\"I�^d�	���?q��L�� ��i�B.	N\�<�ӑ:��;���m0�'Č��� ��ќ2!��1B�x��y0	؎��d;�<�w���@�dD&��(3d�O�	�w����q� �N���O��Y���H��1Q�Hyo!��8�N�]�}�Op]��|���B���4�E�YϸuM��Q�eȉ-�'(&
*=Q6tFn\ڵs�eX[��Є�5��h���a<��1f_2G*4��V��0���"j�l�K{��)n�(��1�ь%{i�*�&��.�\%�$2�[(g9&`36-���v)1�����nŎc��-6�Z�C-��i*��G����-�a��gMPKW8ujMr0f��Jm	T�e��5��A���$��2٢���в��klrhT��m�Bڗ�[4iݘ��H;3v)
����pVQҥ.�9#��a���F�B�����D���\��2,X;���.��D��ιȒF�"y�"2{!�9�x~x0 ��2d�Wn�$��:`�̀_�b5�\��k��g�=��ډ ����'�#z�=�-o�7���l��IKC2D��g����L�<H=w�*�Qw����ct��%]�1'�ױ�8*(jd��;�gi��MK��h~�P�a�vr�'��A�$���f##^�^��,����H��F5���->�pA&[�`�H�fW{���^�I;�� 	��`��jڠ�s��V��d�NW�M�p��B��e&&��\Z"L���+��9�G[��5�z����H���A���u���n� ��{0n���M�5N�֜��ě��^mX�I&E�9wy����=խJ����+��YE�<��6�W3X��T�w�ORumM�ʸ{���E���h��]��iq+{nᙩ��8�.Y�n�Bb�Y.h�_���:�|I?u�<O�������M�I��]x3�]e�1)ød�љ������@'�z�kvN�����F�'Āw�`D��w���$F�HZZŊ%ܳ<�s�Ocfj+Kӛ�����X�'Į�����ə�=Ӷ;�Kf�����sc�&w,ᝃ;���D@3]�^��d9y�/V	;� �O������
5��&��;�Y�B��IN���v�̮��i���Taq�ʠm)�X;Dm����g�8[� �r��}��^$�m�|H5��t;��/=@�nDO����&�7Aӳw!�m����W#�o;j�a�W��%�KY�O�{�gĕf�v^��{�c��Ō֒d�3�w�.��  #z�b|I � �|}~�O��������������������33c��K_�t�j�qJ0��3���3���#٤\�z�;v\=���X���%{��Tթ{��@���fxk6�� �M�nD3A���b�1�ۮ���:�{f͹%�ǪK��ꛖ��/hQ�c��wnw�*��yN�����e�xn\%����g�?^�=���G�5Bp�NҬS�y�v2��y+�ޣּ�w�^�1�e�䷣o�냽6�7�߄M���dc���P�w&s��}��lͻ�����l8�O#��wiBn�:4�7PP5��]��8�w-�t�G�{;���ɖ*����a�����^��,o�\�� � ���в�_����AĎ�
�}|�x�7o����3w��՚@�����"7���O��������
�;�=(��u˩��"ƈ~r�!��D��M۸�U�(~�O��Y�=�������d��.BQo
}���\��PYn���Ϲ�H�z�?zO��F��q�f�pv�!<�n=�����f��ݔe�q�\�C�Þ���|ʪO]o���bC�y�i��x��
Gu�H/Q��p�h����:�w���{u�W�|�p�iE������CB�>��;�i�-[=^r���'�g�K�t����=��V��jy���9�y٫	��y�,_���� ���h\wF_x��X	y�7y9�v/���D��|�=>&��BzmԭԻ�N]n.G����k�hf6`W�!�[iY���@D��ؕ�"�(AJ�đ�|R��g��1��,C�U�4}%��e3Vq��Z�����M�(1;������]��5�捻�h�Pc\��������������))��s`$חH�Rn�O�]��cy��t�M%��%"bCwn��껺�݉��(�Myt.����ܻ��J��Li0���)ܗ$dh�
l�r"&Y���,5��a����\�$#h�!b2;�ԧ;wtL�N��;�/{����4�t�&����iGt�5�����MΜ
0��͉A���p�w>�{�S�>=�9�H��wv�gu���R3dɢ2QI��lgqN�R]ݾ���-D�;VRP�,� N��8>�ml0 �;�L�Bz�[1g��d�Vڜ��.�9'X��l�|	$�� ��n	��N�s6��*���"$�D�7�(3�g��92H��Ȃ�t�����$U��I�Ι�'�{� B�6uWN�c#h$
�E�J���A�>֍l�Bᆖ\��R`{@�k!��r�v����K�|>L�ܳ�v��� �ى��ȀpD��f����~1�I�����Hh�<Z� �rϩ�o�5�l�>�w���~-��ǉ�y L�wlO�i�Ĳ��)+ݙ���GA�@��Hwf`���>wι�H_^�|n�s�Ka�N�>�9#w6f|O��� ��:�Ԓf,Y˻���/���d�Ԑ԰�'j�bA$�}�y^H��a�m}ƻ)�#ӱaI(�F,6��Z�RۛJȑ�	����+�_N�DyQ�m��E���R�͉O��
�7�-���	���{�+� ���2���W� ��=�O�Ɲ�pٖo$��R$yz��>'�����;�nY[I"����B&��2ܴ�a����5kX����Һ3�b�3�]�I
|Ř�d���~��I=w��>$�τ?�,�2U�:kw��c@'ĝ�؂0\P����8g`��:�� ��*ӣEϯ^�{��C� 76�����j���;�	w3S.K� ��:�/ęnm��'j*-��n%Uۚ0m�@$�s�m������WL���j��<#�Z�H�;��OX�Y�z閺'�'�O�զ�S1E�����~D�s�6$��̧��Y��D�>�s��A|+��?ޟ�<��O12c���g��[=��eε�P�9���OK���3�|l��tV����8�B�b��Y��wqШ}�������<����e_������3:	1]e7�4O%&Y�$�]4^3m���sIIb)���.��f��h\a�&e��$*ph�l�n��#B鶶�c�Qm�f8��m�G@�Vj.�qYD��rM�0Zf����\0\�q�����l҆T��G��:- Y�����F�Z��[`8�me��lƗhH�]4��׊B
Rf�h�4vf@��2>lUƅ�nh����)\F+hjUƖ]��0�ZӍ�E��rlf��?��ܰf�������jl0$�Ύ��Y��d2<�*�����A2��`Dt���w�Y��O��\�s>$��ջC�^NV�w��A �	���#��]��'Ǟ�:�5����/C��wL��w��=t�`����$���.�����۲+�x�ѯ�=��!y/W�8�kvLC�p�zo��ы��`˪^�$�j�"I���Gv�]�7K�=1�IZ_����u�A�L?WFI��BXbx��r^m��'��
���Aّگ��XEk�!`���?�غ0hK������3B˚i��	�.u���Q�SR��O��Yvv�����=�;	�ȃ��˲I���)׃ �H��ɟ�E�kN��0wd��W^�v6:�w�.+�w�:ܒt�����ĥ5�RSe��F��8��z?������N8��$�c	=�0yƼ{l�[�w[&����~�>$���fA$��́ ��F�ds�����9��$��QY��OU��s���܀ �g����L���0��n�v�t�$��ǎ�I�3��gL�+}÷����݉ ��!�>��MՑ#Ă/��t6�큇T��X��^�|	���NɈp�/"O<l ��Cl'mv��eU2�b.�b�z$I�� H���^4�c��w�P7�+m<2�f�@��hl��edf����ڷ ����so���{�3u�����&�+�+���Ot>���k�x�dE�̂A �fDO�*t���3�w��~��B U�gnL	 ��@���<g�ݿ�l_�����Y�?���abX����wz�����mx�e�kOE2's^�W���{�Y�_v����o���훻�K�r#�<��)�f�}�u��0n��j�,�%��@%����.��O�'�܈g�}/��$����1�1�9d��q��3��0r��#��	��A"s����ofRni�
Zr��� ��p;��wt��̜�j/�kg�M�d޽����~�I��cĒ:�:g�fK�{�����1>��,hX\Z��D4]tÂ���kj��h]l�ˍ��t��S�}�~��1b%�q猈��D	}2�1�۬9�����|L�>h�1e�2�\�[GWL�Dh�5����	>'ِ�}:�z�"��7��]�~�d��f���6�'Ȃ:�6$�I��}ъ�+�)�� �C��I#+g�e�K��ɱ;;�	��5��,�c�}'���'y�>;Z�$�̍��$��e���d�Po��ޏ㡃�u���Л�[�5����پ|�j6Lk77��p-^��2�sv�������^�������+ԘI� Dd�|=��޿����lG2��gd�OÀ���A ������c�^x��z0y#ٳ3 �	���|~YCn]d9��@i�E�3�s�]�dŋ;0l�m\��F�`V�\�V��9���q�ԟ~�>��Vt��~��j����؟@'��q ���S���g�$u��$``zu�r;�KϹ�, ��i;�:������ρ�]��'�om���W�0هI�+A��.Ab�'`]y#}��''0�g!2�j�8I#��'=^G؆�d�������&`�ӽX��v�]�'�'ǩ��H>&�,�#ĂG7>̆eW��VI#��&|M� P�lvgr�w�뷂O=5�kl�v��$
i��>�ۈ��φ�<�<Y/�J�g�j�k����Q8�tc��r����N)�fX]��Q2�q�ɳh���J(`�"�[<��j�1̾^=�M1��W�p_	���}o�O5�r�j�it���e5���@A��a��biM���/i�� �Ε]�^�R�enC�ġs����Ұf��ͅ�u͌Req��rK�Bd�X͢ۊ���]�2����Q2���d�v�ZS6���Ц��YaZ�رb�6@v\V�����n�¥-!*`��k��R�^��K� ����-#�.�s]k=���R�.k���sr溡	��Dtn# :9�ѭ妹�8N�,�ǻ:x�b���"�}\�s$��׹H>އ��0����B)�dI#�������M&�X�?����}�����ݸj}�W{��@�I�̈/��/�e[��yE�m��]v:	8 R���C�p�z�3Ձ���̬d�C�m�흯Z$��>G��wC�yH���R�����2��s�7]���ӀI��$u�<H'�[;��8��>K�����x���S왘:�2c���ۍ�R6�r�5��� �|:�� ���2*z��xx����q��T�-�3���9L�-�ͣ2�hM���k3+�������?0�t#��b��	 �C\x!�)Wt̝��O�O^�ۼ�I���T�mi.ɋ��E����� d }>�X+'�
�wd��<��a�N��w���չig[�x#wq��G�r�<�ļ��i�y=�b�Şh-�yT�T5���9�k���� '����� �bj��$��7�bzr�ج��;�0.�.�V5�� ��LH �G!�1�����Cq�I�ޙ�p<%���%�I猠�C�w�O� ̻J�>$���[f��T3Η�d����W;Ƀa�v��X�x���I���D�\�@]�B�x���0��Fq����8(��`I��8dW��2�GX�:�Z�,�TLcp�J�d�&��~�w���.�t���K\ Ovl��	Փ� ����
�7�4�căy��	�A�b�Ħ`b�[g,Fx�q�s\��Uw4�H�I}�"=(��fG�h��}
���]J'00vL��-5�'ă׷�@^��l)��;�3�t�<྆��_���I�ҁ6y7�,�JB�b����ͮj�Om<���,���2�2���_ �>��#<��uT�@'���x�z�$�ɝ��2zm��2s�d��JvA�7H$�޸�|Ot=���<k]�	:jF�t��gK�D�{��`�|g��m�Mʮ	�*ɦ�����G�'�^�ב_#�]k�%@�<�e,HZJ��ƘX��e�TԳ[�Ca��P���b�pAg�x칒A�o��dza�U��zk���2$��s�4ɭd]&bg�1���w�w~����ȍ�$�����@�cf�nc!Ξ�KN�σs���lN�� ����w A� ��\"O�~�syu�_�S�	#/nO����$KU#��郻�E��eFJ|��|�2�p �Oͥ��F�uHą�7��<E
�m�We����A�e�L�ful���A25�&!�C�J��`�g8�ጇ�����S�j�1�5&��ٟAW���H7S��z�$�Y���?z��mp wLIMۻ���uGD���$��6�"j��@$���jع%�7L��ui)�t&�F�\DL���\�,4�gw
�ZC��&�1/�<m��2��O�=[2a�SS[�n��u����@�׺�a�J�����މ��A$֧���]۝����$�{}0	����|q�Z��Lle[w9�nf.�1�3���sioG�>=�;I5�����I櫧xy�^��2 ������ S���;���;�2[�j�ۤ��N�v�H/�|���H'�y3�Iն���\$��(��a�jebJ���"Zdv�L�$]lGN[t�t�?V�a��� ��<璪׽k}��gg��_]=���{=��g����{=~�_�4S�al|/�)N��f��d��ʪ-�Xl��p�6u�]]r�n���{ž�B>�W$��@p՞����~
������I��c�c}`o�M���9K�7�Ӕ0�~����z|���-G��+��������4�K��lX�&<<Mڂ5z%3�S�{�_��StZ�jF�=��'z�j�7���R�?�G�g_x�?��ot��N���LK���]Ի�RgnAGOt�0�s�}62�{G����佧ݏga�����Yp��f���o�{ʜ���j#������9�X�3h9.)^�o�����7X���'��!�(ph���t���\�Nŭ������_x�y�zj1]۸{n֓�/�(w_Qk]��<6�àc���yT�=���sY���x�I�sօ��;n�#��^8h^�"��l�!��]|&lO��M�ϻ�p�a!��7�L��Ƹ�a�����\����"C0�ic��b*D޶z���(� x����0y<�jsgʜ������x?{g�,���+�5c���{1�v�;�=仧��[/;�ŵ�"�wώ��3��`�F/w�V�_���|6��c���6Q��9L]�б�h����B�La�Z�^ʩ�f����1�^Tq���\ۼ3���Y�*o�s��
1�Ri��g{uU�j^|�/��G�p��+,wf�ٸΙ����U������Gt��[�;�ˬ�/;����M��>�w��x$���B$���e}��ã;7�<e���֎_b��%p��<7ܙ#a���Jx��c:pb%�\Z(���s�`�?)	Kĳ��Yo��N�2A�N�fk�IxS����/W&��;�QYa��|�f��+��������`�m�߃���?I 8=�8 ca�r�s\�"?s])��	Db��7.�w�&8��ԒnWC�t0�spf4!� �9���R��w"(�����u�D�77d�h�I��2b�#���q��M��rM$�&�1�2"+��W72'.ƤR�2�[���ɓ�D�WYf��\��i��~=wˮYA���r���q��3�D�ۓ!����D\�9w-؝���'wSA%�4�HA1��c
iw]#��4S1���
Xo1Ȓ��8�Msu� .��Ӻ��w1D�"hW�pR���IMI���8���Ewq�$ic `7u���.��N\��$������=,\��i�k{\�wS&wjE��l(��[�C]-�D$�Y�Q[nи�qZLZ1�5h&��X�Z���p\sh��йm��R�r�jD�qi��n��IL�^�;6�Ź3��[N�	B<�B���
f�3J0�$!�����uՍa�g��F�E؋��^��e�
�.�.�--��3h ���g���V6Lcl��U �R֥e��D�2!��fw���a�*��h�U��Vc5�a�m��A�\��Q��aTb��*f�ٰk2��n���l[���<���AbƮJ\B�lZmSE
�6��\kS]��&�ڳgkƌ[�lţ�Ҡ�� ����k��*�-�nƎh�JD����.�T*+\�l�ГK�U�u�cXh�X�a��,�h,��@���4F�Q�L�ơ��4s�Ib��LYm����#u�ٮ��R�rq(gPah��eն���"����v#��ҭ��a��k��fu@p��1Ln7L�&C�ጭ�h�bk��,%cf��XKԥ�ȕ�Y1���IrX:f�;���u��Q��Je4�"0
�hi���՚V�5�͝�Ε��t�"��)�3�l�(ݣ�o�j�&3���&a�mR5�(h��V�76ۇBۥ!Q(me���]B̬ԆU�!.H;�mƄ"uẘsEFK�,`3v�oa\�4�7f�g.��%�u�r$����.JXH�-��b<��1��2�6�W�l�IM (�WV��3bYD	Qv,��f��pU������X�%�b͵#���-��Ўt��Sj�j"P���6�Xf�a[Z�t�4�D��)v��eЁ���<��jhh�s��� l�4�r�[�n������a
 ���e4`����JiW��Ƅ� ���a��b�˰Hb`j����Mn�ZLb�taf��K��Qî&J�&��kC`S�h�Zܪ��Jmq!�ҟc|�y�
����8�-��#_�� ��#6A[Y�t�q
YqeP.�Y��Sm���X�1��+���]th���7fbؔ4��N�%6��"L��p9�̓@�Gn�*Xb�-�V��7;:D�J��[�D#]�5���Y�Ȁ� �sbƤSl��-��0��˘�f]�%oP�E.���i��u�	Y[x�,(˜�)a�KU����[�ڙ���\1	�)k��c�fjQ�sO�>���L���x~�k�"A �{�b 0�\ᬱ��tS=�|�F��̍��#:\Sh.0b^}͑pA�w���x�mV�>'��fI�>=կ�2grĽk��z��Dǹ�V��b\Y��s>$��\/@�8v���S���I��L� �ݶ������)��A��;�k�aڔX���D�H5�o��:��q���A��"&b��S�2M[�:w%w
W��d$�e�>�>ff��\�����	ne��:9�ǎ���ּ���po���p��$��,�5����ۦ�\J#�i�빦)vd[*䏟�`|e���b[�%�8�7r�	 ���d=OVt Z�^�{[z�A>$޸���UIe�����z�z�Ϥ�M�׫�;i�7\9ԑ�Xr��"g˷s�r�����~���F�B�ƻo��o)��^;Թ�E�fа��\D�H�9SX���|���H�����D O�����$�<H�kc��� ǰL�`��p��(�����L�6��A�\�-'Ku?f�>$��Ǆx�c�� O��猬Aܱ.	,�Qw-8��Uq�VLi�A7<�`�EWt�O�Ln��抹� �u��#|�<��v.Pt�&#�H�O�s�ěWر-�Uqp ��|0A��2N]e�Z[���ߟ�}��6�YL����F��a -�*��r2�	���
�@%�kj8??g�|�Z*�7��~m�T��D��� E��h95vz:�G�#2^�#�2�%�	v阖�Ψ٘H�dE�4[j���^	�ޙ^�&Zh_�B���|�
G�'gN�g�'��-�F '�kzbH�����]W;�=���	�����:�'"��\���YW�ӤMN��Qlr�'Ĺ��3�[[�<�C`CO���zh(���(�O���� 6>�x�'{���X�\S	ذd�Ƞkbl>^��!��ο"9��� �}{3$���x�i���F� ��x0H�6iZ�pIg��2	'��=��s���&ଶ���왒	���R��0�!��!��P��?��i�hkW��^L��A؋	��Z�Y]m+j�;Po��ϙ×��|vi�<�3۳	�>$ugD�&�[6�W6r�`�Fu��K���3�gN��M����o'�����Y��ې�d�O�sfd�N��wi�٭Ƴ-w볞')�Z�)�L
��mFH�W�U뿏f��5%����}]��	��ܘ����IP�Y�;:t<��ٝ��K���_������My/�׀H<ʭ^wsD-䌏��GW���=S+	�v/��U��v��=��'<=}�W��v�<�=ˣ�o�6F�;��)=��;�M�k���7K߃�'�;�2O�{��)��;�z��D��@�*��F4�-����E�b'�bdI&�� )��P
��"h�N���w�_`����R&�ib��5ٳ�df�1dC�3��D�@m[Y�����LC?������o/`A� ��֠w�(�fWYn�Wf�Ϗ��`A�ǧ×��d�)��fU�E;�c��ƂI$v_Cx��u�1����:;/Y�	M��	6�-�����A�0���{@틾q*�N>nx�u��DׯɁ1�<�q �U�KP%9`]�-�bǬ�UrC�ͳ	+�����6�Jh�z����k��A�Ĥid�]�2�d�m�L4��f�WuǪ�>x����Dg{�d�>x\8tu��M�^�b�h����9���������o=8���^Q<x��"��}���-��u���9��ٞ�D�GY�0���v�| EԚ^�cY-/���VX��݌lґ���i�)Ç��7��a���b�-�qj��5m�	
Ɔ�����*;�-� ���5��@�G�;�غ�B$���f��f,��uiWKdl�cR��`4س��2JࡶW. �
B��桝�i�=�F��l`�*I��e4,�u���K����j�e�t� -�&�]��,6if�cakԛ&i�s�����]Xֆ��<S�v,$���ݓ|B�k">��2y���ѻ��Ond��O?����Aܱ.H,�O�+�&�j�:�wuMۯ �SY�O�{�D��_.����A�W3�೤<ϋ�5B>#;6�I#c�e3�ut;M�wobk���_L���!a�n�س3�:g2y�2{�D��ۣ��ss�$~G�{8�>J��Jv����O�G�^�2�	NX`�d{y�$I ������)�Jyr�!��o;�d�N�s�gb.oNo�^���e(yX��v-͔Fݍ-ц�- ���qV�s�\���i�Mp�ts�����`f����&q�A�ݨ�A>=�� �����؆2^��5p �G���A"����NŁd�D�ݓ A����VwY���2:��O�=�_�]H�{�����F����\��6�7､�{7�A��g���e�Dםrw���3�_�懇� O�;�d�}���� ��+��o[�6Gyz[P�d˗@��6�s$�}|H�D�l��38Mۂ�9���b���I$��<
v�8r�t���/���UJ�	�y��@s�Ex� �gG�O\��㢚�/�pc�+g.dO���ˆL�3��<�� ����94k��9��$�ۛ�or|d��}U״�f�Aߞ(��5��i\��[��h̅����c�=�%�V�1s�څ�4��`�Q!9`]�.�k��I�� ��@�ݑw����]�3�A ��D��g�wt�y�]5O�{��T�c��|I'���J���������l��G_;��0t�pS�`K'�%�j �|T�<A>+��뺢�0�d��p�N�ﴍ/����%�Լ�"����`[���?3�l����=������#d~J�o��_`�ݸ�с���*���Aܿ�%}@�O�E�,�� �g��GWN�ʋ��A��p�z��	*w�@"{g�{����jՁ�c�A�ܨ�	�gH:y����A�;J욡=�Lֲ|J��H%U��$���O��jʹT'����-�ɴ)vF��029ژ�lηheP&�����+S8%��69hw�ᜳ��
i�A%e[�$Ύ�9tZ��g������D��5���$WUs�H��v�q��h.�\#���T���C^t'�����G-��ef�2�t�V˶l ..m<X�	���Z�������0f�t����[�=EG�ql�q �MwFL�M��p��X��H-�P�z�3\9��*"^  �}������7��6�s�zk�Za�X���U&f��6�2I��/��ݝ�8
~o���_�4L�}�6��Z[N�k�ˁ��`��)����B3�r|�Xȏ���Y�@�[����X��t�%�j"w�	�>�u��*	w�q$7��~�A�������?��r6T��N���:kQ�YbL����U�Ř�B�MG6R����k����\���t�	���>�$	�f�x���x��	�fd� ���'�����;;��dy��-����
s֭��ćA	�Θ��F������U
�n�͝������9f$��S��Q��O]�G�b�8Wm��P�sMS���&����'��d��`���A3Ę���ц��z���*j�I��3��Z�9��[ Y9Y�"E3�d�ذ%�Ȑ>�>'Ǜm��<WXurѝ�.��d��\I�/"w_����tz�����s�fM/��X�e�.���Zsuo��#ۄ��j��p��4嘗	���w��W�}��*�r!3����%�N�=i����p�>-�v��j��4�Ú��[��s<!/�8���.5j�q�҆D�W`��[��d��Nk5kJ�:�sHv�0,\�����D�4�a���{V�Ld�P�X-��mբ�������-s��)�2�����/����R[i1��
�ؘm�3i�f��ڧU���vX�K�V)il���R�S].���=�����궐��;�#a4i2��X֩�ճX鸄Ų�9M^
�M��iX]��\�[�\��V2�d�Nv����p�%�=���GL�|O���@ ���<g��*s����Z�"|I>9w�H�Rm���3�,�::_���O>:QQ��H'Č��㭼�	 ���wYQ�[�:6����'w;�x^1=#|���x$������3M
'��v�O7t �6#X5�]رE�2�}0�1�*��w��z�>��Sot��e�C+~�I-��� F�N�ܧwt�g�+i��e��$�2�����OL@$-��G����tӊy�lD;n��i�$�$��:A��RN���c3�t�u�B����
�TM,0�fYt�9`�������t��K?�֜q �D��̜�R:��n�w��ہ �mVl1N�(�y��ޙ$�>��gs���
/΂$��H59��U ��=�Ei���Ѭ4�����}`�M���������e��g5v���-��vR����������^BW�}2I��5��^����GB���'3�,�E�y��	 �nlI#��g&T�S%��h�O���@	��wL��bA��`�NS3�]ܽ�j�����׵�݀�ƽ}I��bI$]{WN�.��0����<�����]�)�ױr$��؂��<%7`�MM@�I���A>=ׯ DhS��#B�D����ԭ� Xm�ױ��� �(d�փ���Sd�Z63;�7��;���L���c�>'�Z��J���F��G����8��kg�ݰ �i�zd�n�S�vI�,�D���<
��b{ǼȾ�|H'�dH'Ǻ�����.xr��Ѥ���C$��w��͋G��������z�޿G����{�����{=��g�������P��!����h��=�O���3�L�3O��<�,�ݽ|6����E��P������28�X�/U+��ȩ�tCS8�]�==/��-pb//�u���
�wf���blbrzn��a�ؖ��v�ܽ���Z0��a�6�UD�o�nyc��i��q)��#���{#o�t]}�`�}�&��k�������;fx��.<1e��G=F��q�Y��{��`J�%���C۾�{��_{" 3��?ks��j�{p��))�|���َ��1�~�p��7�Ŀ���+�$��W�x�7a��ʽ��z�%��L�_��i��!|�[}�p�����k����o{'�K�y5�� �/Hm���]�噭e���7®�77�W�� ,�F�Q�'��i]�5gc�����E{�=�l�����6q%w���Կ��^�F�=���c�Q�Yt�l37�����{��u�|e�v��s�r��\(�����wuÂ~΂nd����x�Ǵ8 �뇅�Hd�{�������wK�txLG=9�Ftf�w:S��#s��ڼ����`ۏ��R��]�I�ƺ诂ɧӊYD�:N��2�-S����<º<���U7r�"����x��z�>͏��{�����1V�M�=�J]��x�v%�!��^���Z�+�h8����������v��8��|�����r��$���H[:m�KH��l��w��Zs��Ol�C�:Q���$�@��xx�I���,w�FH�Fa��2��\�	���c3@��h$��g���.��Q�wt#�Q��M��%-�:H����s����H��^늑�DwWc #$����iw�I�n�e9\�5���	�<��<Ѿ.R|WH�e0�#I3d��$N�i�������]��]9�ȗf䨈�n�����CM$Y3�rAI���wD˗	�l����
#&��]D�d$h�Il�(��H$9��0���HQ�s�'uĒ��5�vP�"�(�e0���܊e��QRN��fM3&��0M�4����M�rR��Nn��\1�6III�75ԙ�,Qb�"&*������|H��������i�>��D�~���=c�
�Y���=P1oZ�F9��ח�<L������ ���5t0l�{ǰ��g�A""��1fg��y��<�H+����-m�������7�9ٱ!ut눻��P'϶�����lX��,���L4�q�˓m5����lk��K�\Mg�߿t�����{��.dC�޸�$�Cot ��ާ�z��5�T̐}~G/��xv��w)�� ��uS�<���ŏS����}x��wO��u+��0����מ�$v�6�d���I�ڀ �J��I �M���A�'hǒ&���|��=Wք��ݒ$ �3��URe�_�y�؀#��< �AU��<D�o@��X�MjZ%D�^f�޶v�p_0�*�m�����/9�p�z�Om��;#���)Y��K��:�<b�w�<7������UF����Y�Y˗y��ߊ��lH%�(��ХX]� 	]�Kgt�k��Q��oJ����t�Q^Zō�Kb��W2۷X��\�E�4a�]��X$�QJ�Ϟϐ�.6�
ͻ���}��8��q �-��&+���<�/�[� ��q荞A���t�f}��@�v�OѱPAu\y���t�٫Cr�6��߻��'�?�	�Jm��=߅��f O���D�_�e|\��xAY}���3�o^u��d���I�ڶ�nf1�j�L�\ˋ2H����R$�����6�Ͳ�)�i8�p ��A{�VId��w����I���je��UyS��*����3��gĀH;�� 7�D׷�Gw�����{�{�'�\s/_p�&�y�����n-�g֌ݙ�*�W�g�g��=���x�~�o��콝g��f�-���lr�-�隘�H,�[s����Y�RmFc1T�6�X����36��2�������U����[�F�d�)�s���G�$ۂ���M։�L��3XZ���e�%f���Q������j���X3nJ��L��j�(�H�.%�c�5oa�+��]4��cR5�@�MubLZq��Jу�e��՘�ٕ6J��J���R�Ư��.i{l7$�Q�KG	2����R��źО����fA3�.�|b+� �}ؐ�^C�� �#��i]�Ǆ䈪~ɒDy���fg�wp�@��&�_e7�s4A`�׹��M?dI䷯`@ �W7=�	Z��]�l`$=F��A�:p�3�}s �:�b$��.�zo$�작$�ݙ�vz���Iݜ1L�&�˽p��(���x�w�G����� O��ۈ�~�G�{�×�'�յ2H�vt���d���Q�x��1׸x3�0�'u��{��I'��= ��?d��h�m�D�	 �p�2H|��Hn�4zݓ3a�2��.eѽ@ˉEhL�w���+2�i%���w�ٚɟ�/����@��Ϸ�qt:22d�	��"F���f`�˗x��:�C��=�8��PK�q= ٱ�1�[]�r����.��|3�]j^�	��K�L_1��ʢ3�_����~!�{��Sy�����Dn�p'��>�ۈ$~��|�1�\%��27��TY�a,��.��ź�=����q �b����0�T���Σ�)�[��z2'�I��c��pŝ8f�W�y�Rj�;�i ���2k#�A :�`A �q���cb����< �Q�rΝ'vp�3ȯG){��=q�%fK]�v�M�O�v� #���Aݸ�]Y�F/@KX�D���fp�RČM(�ط@љ���5�],�.x��4�-C�￟�7	���8|��e>���-�!�g�K�<m���-��ڈ���.�4IwgL�;̼ut� n^W6n6��C��	�� ����$�w�lWn�Ϭ�KFP�4Ys+	vf	��w�/� �H=�'�U��B�c���W�����x�X�?%�>�nC�����\����7T����8��㾳��C��ޛ�'9�}i�f������o��'���d�x�!�;:	��@��~������b�4�h$��<	'�c&A���m[0�:l����{��#��i����>��2#��@�����Ǝn���c׆v����t�$�:�'����弋KbH ��.5J��l����4����vie�Z֍]�c�e6���w�	�e�������A��؟�+zv �w���Fc�\$w��$�����vb����I��x��9z�离�$�&�2d}��t�� �����/���=Z`���̉	����k�A ���A&�z2����ex3������$oN���`gd�3�.�@�v�i�Fy����$�]�I��s�$�Ʋ<'�DGӡ��z�*]��Voў {�����&-�bVj�nӝ��S����U�W}#Ļw�KW��#��gU5��HOE��L�o���>$K��H�d��w2[��AsU�x�dZ��Z�����'*:d��};�A:ݑ寺�/Y�~�ed�X���m���ʴ0�\YV]p
�-t��2�"��f����~��;�,��7j����v��q �m󥸥�b�	�ޙ� ���}(��;n]ӗw/�L�^=�O� �D�kXS'շ��ޟ$��x�9�c��i5K7X�zk��֌�v\��3�I�E<�6� <W���y�>#�c���h�[��x���^��A:ݐ _��I,��Ȑ���n�����uH�bAi�� �n�O����ηB�s���uS+՞�+BwL9r�4�[�ǻ#`&��]h�6�lrWWDx_��p$}�����l42��#dLzC�eؼx�"n�,�oeyrm�AIC�Pa�c[�
��x:L:{tb���Oyu�D��.���T�i��	fbJ(!/��������5����00J˛Rkk6����k5U(��p�xͲ�We�g�6U�Mc��{�Ǝ1555��U��0RնU�R�K,YhP�cq̤ts644��jh�x%ZC�CJe靆�]L
��:\3���e�M�^���CD+�B
�)�Цn3��e��F6]�P�i�`;�Y�4.�e��Q`�EJ�����7#WiVVŗ*H��n*��+0%�Q�:�+T��!�������2wd;���b��|�{����	�����ݭ7�1 �����Ⱦΰ�pŝ8f���|��
��.<zt��l KvǠṱ���S��.�dH�}ܚ�+Ϝ7��.�_̙�e��$*�:$�K����̶\��ȋn��mO�<H=�	�gm������Рr:y��^\����g���+�/�fA>$�v�-s��r§�Q/�cč�^�K;;2$'/T6�dg�@�g@�h���o��z�1���}�� �I��<��z=>����!�'��ُl�ʆS�h�.��"��6�s�B�bZcf8��{�ÂwL��;�wƮ썉$�DwtA�M��Mj�'��펙 �z�i Y;���HO�b $�gkչ�����\��͛�nu�	\��y���c��Ɖ5-D*�M*��c��m�3����#K~��Q��>"��sQ���z�1�Y���H��ɒi#���3��V�ㆆZ�VY��J���L9�I�1gN�]�>�ȏ$H:ױ�y_bk~Zj� I�͘�g�ȃ��DU�.�˻��&y��53�+�h���}�����3�$H�f��H����TF>=�$���'��T��wp�y쩈$��M�4�H��*ܘ�ۑ �����J�s���zku��`�~&�-6�ն<R�s�2���6]�knX�˃M��wj���ݙ���=N�|I�͏A�F�>�]�/�ػ.�j�D�әv��KwL��3̃�-��A��cvt7
c<O����H5�9� �m�&�-���{g=Q݌����w4Z+c��[���4�}:˞�C]�Ap��J��;"7ѮT!���3{G���2�Ra�,�2:vM��H��s;b(=jw+=�@�۫{�X��s���v0dj����MN������'��L,0N��NL��\�8D�ӽ9�Cv��>$sS�w�q�� �ք���`AăYõ˺r�����vg1�ǉ �tlI|���9�V�>'Ď˸�I������-z�h�
rfD���L�ww�@�B�8t��Me��$�r�[y���1�;5��b��_߻��wp�	?�و �y����[Q������{2 �|H��c�f6;�3��	�z,��@ˮ�輸jz�o�y*�7:�h�@���@��
��.�r%.�Y�;�g�&[�"I�ؑ�A�Sw�N����4�8\"/��I�l�k�ձ� �/�l�,��0d�Tϯˢ�c*��j{h�b�$��6�2}>=ռ#���+^��;a�^��C����-wS}��rn��Bc(u��8e�>'V��CXl�s���b�r���"F�,��^�3�=��i�� H�n������`���ND�F\��+�؂���p�Y�����<H5WO�'z�%OO��ͩ�$�H��]L;K+�5�E����J]+u"�Tu5c4����Hm��]��w/�fxƭuG��.�2$��=ձ����6����G�B��I�R9vwI��B�~�qLѝ����L�t1'Ď̍�>$�؀w�Gn�,>EJl�[�Tײ�gwfbC�y�ѕ� �H=�� �rVڢ�2&k�Qs�f|{�"
��|�	 �I�g,���'�УN^�l{ǣy���|ss�'��I��tYv-�3��'MΒEN�L�e��r���Q �NסzB e��M�Uo#��@ڋ��!�؀IY��z?I�?w��.��~�W?�@PE���_�m�?�J �/���a��n8�&ٸ 8���
,��0���*,ʋ2�̨�,��� �2�̨�
,��2���
,10"̨�
,ȋ2��(�*,�2�̢�"�(�,ʋ0�̈�
,�2�̨��,ʋ2�̪̬�́2�0�32�)2�)2�+03+!)0�+2�+2�+2�+2��0�0303+03L���,��,�̬����30�032�0�+2�����3+0�2������,303�0� C"2��C�*`�C�� �0"�(C	��0��C �
0"`��È�C*�6B�`� C
��� C�(�"�;ˊ�
c&����ʋ��`쨰ʋ��ȋ(��2�̠�*,ʋA��0���*,0
�(�(,ʋ2�탴쨳 ���0�̨�,0
̠�
,98��,ʋ0���
,�+0"�(�"/�\�񃎠Û���UfD@� fO��f�������C�;�?��~����������������:76�-�?Rf?���~�����~@(��~a������p

�~$"�������O�/�����~�?� �+��Ӈ�~��Sd�=��:������~�? ��+�g�ࠠ� 2�(!J�,H L��(
�ȕ&�R�U5������@ HȀ@��� 	
(ʀJ���#
+ �		� �  �J��?�H��a�,��?��?�"("�"-@+B�~���������B��������:�Q\ׁ������~�n����>�7�x������~ ��և�O��;7���E� E��}�>�w�N�ͅ@A^>���oDE|�����^`�� ��g�s��d��6p7 Eo��}H�o� E�����:���w����po߁������@�q E��<#�~@(������'ܻ�	����~x������N�	:�x ExNi�:z>�����u���.�S�/Њ
���ǎN@A]������~�}����e5���9�h%� ?�s2}p"��@zѣKF)�)lR�R�(&` [�T	h jؠ 5@� ���հ@��  ��
	ς����( R��
	HP��T�P  (�P� ( H PP ((�
P�P�i��               ��    �P             �        �7�nwt��:�3��6rn����mu�*m����ӗv6��
E� �k�9WMn��% P� �   �=��܃Iq@:$n��ӻ�5��� ��w�  9�� /@�.`�X�P6(=�t��{Ճ�`�w���[|   o�        � f�{�@^`:x���c�4y�� �� �Z ̓���]����h� ���4
�� p =��lw�@)B�[�  ���Y��=<���E� ݚ;:^�]��c�����Xqp ;��M��{���r�j�ezI��<4\ҔPP |   �     zP  ���\�_o@�j�ku��Mnw:�L7 �A��Ӆ�f�Zղ����kn���Ӏ�]�m9�ࢗ\��P)!@P|  6鷙���m���m-� ��V�sj��u�f0ӛv֛+Nή�Y� ]]���Yq�[ks��-6�hԫ���6�(R�U �  ��      z��b�6U�]�Y�m�\�U��6�iV ��^�/0:�)t�ͦ�k�*��K���ڸ �m�n��6�ks��0�Ed �   w�����U����[M� ��ڶۭ��n����]r�m��[�l� ��΂kl�ݵ��ܳ��ks��[l��I( S|   ^         ]y6�s�T25�ˍl�7,1V�mY� �v�V�8�kj�YJ��nYv�ƴ���jTp ;���\�Vf�l 5@
}�  ��|����wi1�p ; :�c��9:�QM�ti�n`�M�k��\��Rw7Wm5�;R�ʹ������EJ�z @��b%)P  "~�U)��@ ��~�M)( ��R�B   �M�)IP���?��?�?�u�/�������_V���f/���B�P,����%I@$$HB��$�	/�$ I0��%�H@����������f���_�-�1����U��b��Ti�C��6Rɔ���*�l��(�.H�����l�F�.���.ܞ��$0^ՋM4��mGq�*�ݬЃ&�{�&^���A�51��O2���FU���R���h���4��kvq{u�Mk������k�.�dm&��.���u�Η������fE
J��\��׹To
��8�lop�w��h=�F�;v�2�,��լ���L"MSr��hzCu&c=qT��e�%1�,��Q)��⼑�t@�Z��JF�TQ�'���p�R+ODP� N����l#�\��7{B��͒�D��-�[P�F�Zֈ���Ӛ,VcI�W ����/
�6�;Ӡ;P���Rږ����[�b'�������nl���.m��Y�͚74l�4�M��-�v�Y�n^2�-T�vS"�X��.U���<�*c�<���,3�C���N@1��C��H0�!B�n�Lw��-�:��7���2桰���S�7X8V��x�;z�nL�#n�I:t���a���5��ÛӦ���u�&L��h�ԩJ�K	+* &`��M�V2;8.dO1�Vmf�z6�����0�S3kC-�F�-�n�:O,#V&��d�W�.��O�� �sF{0!L]�L8u);�X!�4 ^0� ��W�^݀.�"�xĭ���"�hS�%��r�Q�R�5r�+���ɤ��*&J��͏ON�8����&�W�6��]ٓ��U����DX`��KTs�6FZy�b#��B	Sd~;D�U'S��"ˉe`R_�Z�^O%�k������tq�x�;X3FZ���n=6Fc�ފ	h��qQ��ň���[z�xv<����Tos)#z=����)d�b�2�����3mt��k�B�f7t��2f�8�vp�evNP�]=��9(��w4J٘�2Ws����!�q��e�ع�r�ږ.��Zjˊ��B�ۖ���k�5[#��E���h��������L�M1X�I�t��ܘ��M*���^bKv�sJ�n���Pf0�˧a]�9�	�7�,-��x�,��{5�n��[��=;6����~�@�HF�߂�(	��;H�on���&K���`�beD����򏋑;q��䜘���>v��*�2�.Xǰ�YZKq�7i���=�J�AN��Yֈ�f�Ҝ̪�����)n'IG�NV=��O3N�PWe;��D��d�d^1u�)���F8�&�ce���kb/`d�@V�!l�
���-f�`���nT@�����f�	aI�V,V5�%z��'n��;��@�S�&zȖ
�D�ybP�i�ۉV����*a��m�v&͛kDŕ#sLT��"Y�4b�R��ܙL�`�e0yT��zx���a��Je��gD���NG[dTx^g�b���d�S!��n��e9�իH�����;(�i���ӴN�j���tŃQo-�k&��rL ��1�ɑf,٢ 77U�U��Le�/����v�*R6�=-^i+�'��#�P��1���+.�3r��elP:Q�3��;�>4�ʷ�z$&X��lܱWZ2�8Bw,�/X�W6�a$Lx��
}��{s3�i
��]�Kx��ˏC�80�H�{g\a�z6��J�I��L���@��EC(ܪ�1-k"�c��Ҋ�I��nM�Cn�p�qQBנ�b�Zm]zx�S,eE�!�	-j�f��s0U�`r��ݩZ�;�ϰƙ;l��è[:� ��x����)�k1����%���p�lrXͼ�����q�Of'Wy�^�aS-��`^4kt�����ф������7����鸲��^�{�Y�)^%GYM�q;��ay��D%�]&�p��.�1�D�]���	���r�ݵ��b�ka��u����뚳S[�B��M�e�ܼCi��.Y3���_�ӹsA���R;VsT+ Øm��jY�R\�L���+9K�h�TCD�m.d�+��Պ�{d���:365�S)FHU�+2S����ߦ�A��Y�jn��U�� �,Z�
Cl�WRm]���᠌2�C�/���1p%��m
w���]��R�J��A��.[��4����x�,r�l��Ԇ���[Y�ӏ��Sc[�� ��	.\Ԭ�,ܬ��6�`!��!����,��em�iQ�kwbWG#XnD�r�גϳn�9]y\��=(J�Z����+I� ����kya1+��V^2l�5 ݵaM���)��`,���[yg2}��Tw��v,�̬I��� t�@��WN�[�!a-ג�J��Рܥ��"\�e�wZ��Ӯ������ek��j�5S6M9[M��reMܤ.�k+�+.hsi]mj9D�̣S"oF|��tEط$CPC+-�j�{r�a��u��V�8�$d�.�˼��Z�� 2^���Yp,��gl=/o3�M�&��.�VRc�5_����K�M'��"7����ͷT˨���l�Ȇ���1ݷ�k]M/,`ۣ�^%ciҨ(���ͳ,:�h1�B{6�b�����h�8����*,�skt��0�vH�_Y�M
��'*��׻�����b��z�������o )Z��X�}���ʃu���)�I���u%¨{��A��/��*T���ƃ��ǔ�$�e=���2��nL�
��%+"�1%�EP_A�ګL�Z���p]YR���`#��X�P+3r�eA�;l��/v�dh[a}�!J�$�2���tL��P�07��W��6B�9[�r/<"?�[�	�悶����u�A2Z�1�ֵ�T�6�n�J ��ʼ��C�fI"���ypbʽ,��yn��23o6Y$�q;7��l�����7�m��^Rwv4m��i�ysl��ChL���{4G�n��2�h�k�ڋ78�h3j�U�Z��)��
%lYmn��Y�XVdsf�V���g������Ȕ�8�a7&Y���U��C�رrR��9�U�	VeQ�1�{�T7�N�֕�����j�VI��ni���q6ٕLMV�3U�mF%�T�@�`Z���5c �*,ܡ�ws,`�su��Zʹ�*K9H�1̪̅�ѵ�ϳ^c�1�#u�F���S6�d�̛����Q���`d�*�cw�Ӓu��<)���E��n��RSec5$��� �ͻU�����x����$Umc!�n�,�XZ�zs1(�4m��p�Q�S�7pջ*^���)nZ��me\͑��y���ɚ��� ��Y+tq�(VXg*jٻ2��ܶ�����ј���an�;r�kR��)m:�b�M�9Yr8����60�;��B���'����6�J�3Yd�(븕ԭ��JkXua����Ө��@����	�ݺW�l��W���3�1�����^�U�\T�N����^Z6�����p+�ɘeĈ���� +z��ǭ�X�ڶ�M��2H�K��DyV�U2�i�7��*k�4��ł�aP�ݩ��(,[Yu��$t��a#N��4�E���ދ',��TF͆��ҹ&]MK(;�^:�Ȉ���AMћVڪ˖)̫%���L�(ǁ����F$���X�C�N�	4ar	����-퉇��B%��<�p�{J��1�2���j���6ne�*[ 5q ˣSH6�:W�����^X0&��q����b�_;��m<4�^��m^À��B��˃w)���Y�nFM̒�5���LN�V�n<O���,m:F��0���qZ�͌�)P]�&�$h�����#jP���[⎬���ʺ�5�kq5���55�f��BH?�us�*��G�1`�(_�f@�݉���Ci˨7��l;�i)�*� L��u꼸1��f/�����IV�giG��S?Xյ��Kj�L��*=�ݼ[N���h�Z����x�j���U�Ol4�kp�R��G�@]���Tt���k4X�ܗV�M!�w)꣛c�,äȩ,��*֒��z��*ܢo@�`\I3�ꔅC����RR��7���t��h��d��5v%-�3�spZ��Yiy*�!PTr������ⱉ�d��FB�&�;mЃe��Z%�2��'Wm�c@��Ǥǰ�r;�Kv�mGF��V%e�vj[X1e5���#X�4�P|��Ůn+
kZ3)'�;�)L�Zr��7U��^����s.<ѹ��f(s."3,��w�6��j��I�DdƁP-�zN�c+	���9�m����oc;���[A�I���N����7r�Hسj��v�%��o�5f!t/v-0ݘ�OE��t𖉥HU�Ī8*�M�#�شV�2���j�E��MYSv8ڈH2�2t��ת�^=�<�r�U�V��K�x�<�ә&"8⻌�҅J�q��z"2�
95R�P^+,RA�є�:YÒ��*}�d#3R\�O��R%�
�Oh�ur�P��T�"��bv�wq�Y����w��%�{Z�Ź7akY�3*EE�մj�,Ӭ	�����[���6M���!���J��C�v�]���T������r1;3�N[�
�v��i�v�9�yB�u�1�v��m�Nl��%۫Xov��v%�6��0�����ʥ�U�ܘNf���(1�iP[���	�΍N�Rb��/F37o'2�Su��D�2�+ ��v�0��˚��M�2�#��=�7%���k6��L�X�e�HV�� ����՟
5^���2��ψVk�}�����qJ���0^/Z�!rW���Ͱm�vu��U���`Z@nT�t^��=6��Y7 mm�R�~����Ի� R#�����3�����B���[㸬��!x�f70�S1-Q�ދ`���\9e���l���<u�REG�6��5m���&%�w��˽���L�ձ^���
���`5�DLX-�;�AB�f��t��{"���M�V���e`�Ɉ�n^�x�+B��`�,&%�ܑ}Q +R��)�Z3Qom]]�6��T�͋����y,��TdO���DJ�KjT�V�9y1s���L��P���8ޙ�:��njo؊IVU��V��V�(ږh���[O�*���eՌ��o��P�K�Sm�Y�d^�)��w(:V�SW�/NJזU�ۦ����v����H�ɕt��lKN����M�TXP]���X1{�;�U����_n�����*��يAb%�Oi!F1{�շ��kBk(��ʼ[�j��M�nTL) �D}����
Yiޒu�"YVa�w�QJ��E�I��rķ��U����*���$�@mUV��b�Q!�>�m�ڳx-m��fñ��i�Ph)<�j�#CBY��u ̒���Zoq��E���޻y4�e���ػ���[;�j���K��t�4�-��/�ֳmnR���hQX�ɲΨD�CP%ԇt6ao	D2�q�HG�EJ���"�Z~R��&K
 MDw.�',+B��VZQ�V��i�hV�.!���L���(���t���n�.۴���u��n*�:��Ù��2��#�w6�X�%`2�^2�C.��F�)޻�-)���XM]��C�s-�8Ԧ��b`��U�Sܫj��(�͔���Gd�Y����(;˥�o!�W��V����jsIƯ4�!�[.d�f,�F�i���4%����3 �%�&3�mǉ���/�pc�0�k��Q6�錧w��w�	[�ڙ��^���QͿ�Q7�>�6�M��bly�lL�e<�bʔ�J�R7X��
j��i뺹#�7�p5�n6� G��P���M�����J��
ՙ�r�	5��N�75�f�֬��� oE#�%��J�2���%����S+FKɄ��{-���*GN�4�R�Z� ӈ�k7fYյr�`�ܼ��.�  ��j�F8.�fl���2�ɸ���҅����i��X,9�ot
˼�t=2����f`P�쁦r�bz5Y�opR^���;�[���ݚ�e�f��d�5/9o!j�bdƜ�M�	ۭ%k��C2��C�˭[B(����V��٪\sz�^&M��w�S)"--�P�Ʋl��gpn�)h�GS�t�	,�VEL�;_'�Gtn�ʬq����T���WO�X��� ��\If�f�j�j�"=VR�Հ=a��$z��ْ@w�*V�kkE
�{$�X�㸝�r=;���~	cj���y[X�^"bq]3veL�.��庛�sp���4�bx�K�u�qbR�H�#$3@<�����wc���+0U�����<�dҍ��T��6�EfneԆ��lW���7u%Z�*	e`�P��
�*V��O��a�e�r|p��ʕ����0ퟲaLݛ%IY��.+�D!����=��m+d��z�v�	�v�af��6�L��A�smRxi�7`��dWPd��`a���x�X�x�L^��^��DX�[���~q���yQ0-�T%+��+�d%ܒ�73k*�c��E���ph��g>�E�a�Wy���F�e[�V�A�N�v%�o]�w7)f��̂����;�h@���i���(�a�gg�3o,���f,��(Q�[�-��G�#**Y����i��)�$a�Ǳֹ�3nS.a�WZ��
�(ȳm[�1+jٰ�i���yo0@�HfR&�D�Nm�4k5�j-I��h̸��bw2��
�ƞssk^m��&��+YV	2� l�K5E��Z(� ���B��Y�P)�.,��G �g�Á����=�^T�U0���1$��B`!�$i	&� I!b��6	$�BAu��u���]\u�utuUGUuUwg]���u�WQtu�\wwgwewU�gu�Q��Y��wW\uwt]tUTu]�]�u��u�Di	F��6�H�!��WUY�u�wq��gWvw]u�w]�e��gu�W\U�u��wTwwq��t]wwq����WuE]�]�EQ]�Www]�e]�wU]�u�q�]�ww�teWg]vu�\UU�]wVu\wYwv]]Q�	`�$�i%����.�����������:�������.����:���;����  � A���HH� �$���w��c� �
y�iU�R�
8ث��e-�������W�iL�wG3�WK�wGr.��j�m��������uԬ_�3:vpm�RD������V�߯��H��@֓�ۯDĪ�l]���2��<}A	�[l��Y!#z"u�O	�Y�nbҸfL3z�Və�Sv�7F�*J��ۊՁQcZ7Fٖ���WSq߰�
8E]<�l�,��jwpL�t��e�)����SW�9��x��"�
=Ǎ�tr��3Fm�^>:_U��3�l�x��/<������^=
�m���Șt�Z�2�EƝ�?f����s�ch탙�e�FL�R&r�W�E� ���]��Y�U��"���mw'��2�B~U��\a�g��O7�Va�]���CV��kۺ�ҨH���j�zn�M����h3��h9�:�;y�K�X��;��9澨���Y�f�w[|�t�0+�[�V�zsɃ��x�F�]�e�:���7�sњ�N&0��ĭ�=�Vm��,��F���d]�u�`ʼ��ȭ��gk��LՕ�9]�iuݮ��ݜ���h[Fn�/ZX��V��6w�A,m�,�'�k�ͮ�i瘱բ.�S',�N���	�;["Vq��6Hc|�uj���*d���.�w�"t��;;@=�\u��Y����ݷ.�M^P�Y�W�U:�V�SA�������!vV�n�p�j����>��t���K͝X�_���X�X]�֝�s�ٔ0g-���v�t�Ɔu��Y��Z��kFv>N��%��[YQ+�Xa�*Me�I]n�l�O͕e�tk��4�w�6˵o�N�pP�hC>�2��;���Y;/G͡���Eun��j��H"*6���;T�}����(p��^�6��1m:��&��6���KX�޻���S���d���������Rb&@z�<���D՝�n	d�+N;���<Gw*��7;S=�NC*�$�mgv�2c����Ymd�
�+&˗��8��:w0�ܝ4�ht�cd��ok�2�q-��Z)˸k���|la�u�r�عe�D�XX�a��͘�\r��O51B�zV]E*�v ��T�sN��|6�겴l���ES%�v`/Gq�R�����ذ�5��/q�WK/LZ`"q)팬�uc��f�e����31��K*g�G��n���VI��c.S�6�][b���ٻ�..k{�{�6š���~DW^U��uq�
��×J�e��g�cw�p"�k)�a+Nٰ�o�]��JmP�T'F�-�y������+zr�RhTڜ�4^��smLَ��Ǯ���_Bv\��u&�UC��:��,�YqE�y�5�1uvI�����yl�f�:k�bU�՝��N�J��n�����c���K̓M�)k�J���F�9�4�e��؄"V:ͻ�)���|3��v�vRiZD�1s+	]Y� �j�O^�����ٵ
�{�te;+u��2���s�̔R�g!{&rS�n�]�ՍЛ��PU�ˎ]�R�K��jY�	���ِ�9�a�)�\kz��<���D�wr(H9Ӹ�F۬�N��KM5Y)C:���[x���Ճ>�=]e�l�9͆q�eĲ�Wu��8=�ܻ^rX�G��3=`ĺ��� �lgvi����YCN��;��WiŶl���KrB���U���gJ]Csv�d3/e&X��.�o4ɦ���w����+aO%�a����vb��I<�v�o��λ)�lbO�v�e۱=�4#������X�ɯksn�Cbj�+��\��'c���5��cB�h�Q�D��!��V�v�Iu^'���#�����Y����ӕ�*f�h���N�f��BG0���ښ���V�j'y#�|�Mn=��M��maA���y�Q���Y$�]^K �1r9�;�:Ƅ-G� 현�6{��P����F��
����Ǜ�����8�j��h���'yy��J�7����j����x���8J�{�h�&s_ۭiY�l�
�*�P�[�G�Q�r]��56�˩3)��YZ��
N�YS��#��W
۴y��.�@���9Zv��K��<Σ���l��oDww�/�W{�\��Wu+�r��9".�Y��$�w:��u61�\�ݛY7����۹��ˮ��p�ۖ�kv����b;�ҷ���MEV
ٖ�륯;6����u���;R����V�������U����	6���f��
�`���^W5s�<j�H/6o�xM(���Fh��CZk5o[��e�Z�[�����>O�`�s��jB�)RL��C�wT���]!^�35jT�X&oYR!����=�) ��)���ҝ��M�� 'L�޼�@��d-����*�j��am3�ޭ�V����w+�9�h�7�����;{�zmdyȝ��B0`����m5�57}r�t,͚�!���gz�vl��[��Sj�/P�B�6�b�� }}�����|>7z7$�a�9ڰ�,uƒr�T29�Mх���Wt:�s�&js��l�K��Guo7J��e`�}��I��е|��SY���nfY���RB��N�3#��J�MZ(>x(m���;,�ev%zr�%��\�ފ{�m�2L�ĥ���L_NTsxu#ػ^�@��޳�����@Ớ���`��/ӇDt���4��(��ѷ�k>�z�,�]�x{`�x�)�;�m�)ՐTؕ�w1��q�HU�%�������ʹe�{|��EB�>��L���)a��M� N۬�]G��rK���K�__V�b���L�C�aU�7�z���k���#�>z���^�\�-���(��Ӱ������ҏSv9:��^˰���Q�Kvg>��]A��VH(Q��%Ϛ�%ͷ��9L^NU�_Q�ɬ&��GR��Mgy����O�����;eX���q6��N���n�ͫ�E[��ee����id��Mf7>��U2g2����__#�hZ��Zy$��n̯+�@��z�`�,X#%��*���n�O�v�BT�W��Gɜ��L�.H�w.�s�Cm�꛲��k�Y�^��+s�\�n�1���Κ�ы6L円+.fL4�k�K��bZ[� ����oͥC3�z%r�ɖ�G�j,���������lۜ��.��U%p����X�:]�9V@9*����(7�u�V����wC�D9e�⣜H��ۙ�9��]6R�lm�˽��#��ތ$�J�q�e´u$.�l��P���Eer�m�@ԔsMe(�D爦��,%JYw�r�+Xv@��c�:��v;8�^���˳��Gc��˫�o����fm����zU�m%7��}-�ǫNA}YcnN��-k3���7��6C�Z�+�d�`����dJ���;���:�rWh�2��#��.�M,����Yv.]�"���־* �.�;x�ٚb��T��%�I^P�g�ˋZ���B��*�܅𽘺�Y��@Z]���Q�m/
�}v)����	�z���ݸ�� �mit��/E_b�E�io=����mR_5��*ݵ75�q�^ldP ��^�U8��v�9^�f�z�J����]�g�5{�m������e���
�Ј�P�e����/��Wwk,�V�LA�*-ή�e�����4�F�CYْ�m6%�d���&*��4^G�c�v�\����1i,
 B��OK+9�������i�(XB �}��^ ���z
׉�(�dK��[�ɂ�>�J�o��I�n;�ή��x�?:K/:<|�pW.�#���ͭ6����xF�p	����������e��V��mL�xCm��&�pP���2�*I���n��pMX(�Ȧ��8A��c�V^`��^v��LҮ�3(��/:��(u���e!��,݊�Jki[�#o�����y�ZVǈ}}3E_�6�HGg9��;W�N�\$���W&ܺAӴrg�Ki�䩾%�[��ɜ����n��9K+���Z-��ne%�2�+J���bi4v-�C�N��E[�>j��޵��;��>������&^b��� �kT�N�3�[�B9Bؕ�_J���j�4�#��ս�qv^���g[x�
Z��aP틃�t�j�CO���tn�*[�a�|*2f;ۋ�E�h5��K���'	F����aF�7F\�2OUUݬ�}^�d5���5i�����k�}�R��M��{hl��Z��A*.�umZ7[�
�ݘ����L��\�5q��K�Z�cJ}�f?���n��[ٚV�N����y�}���y��k�]�]����m�Z&�"K�����M�	[s^s����LK�kv��^uM��^n�ɘb�۸��ⲛU9WMgGPU��>�ܴ�=��v7�0t�7��eI�:53�la
��5����oyV�W�
��]pEW@T���4e�,'��j�Y6�V�^�v��<s�	G;��d�g�+��X&Sio��u��V⹻N�zh6��%�j(M�ɵ6����^Ӳz��<O,�pPr����K:��1+�vV�i���}��u�#;z�\�V���5ϴ�����h�;�0�!���8���/�zv�r�1�J,�9������,�����/���B��T�͊�̶�6q��a m���F���f˓��	����I��5�Ф�D�[Z�C�G�Y��.u���n��/dt=�,UV�\���ze���]2�XgJ�z]�+dȆ��)`8s/v.�ܼ�3 ��Go�M�Z����<��N.��ZWPU��cU�o�5�!�v�>�ޠ�[���� y���r)������Mswr��8gZ-f�"�y�(n^�q�Va�C%j�4V�Q',�Nv�T�4v�SM-�� 	����U���#W@D�5<�P�4evN��w��& -�|6�x��2�Qtf=���K����+fAt�b��<�v&����nt��C��[$$�#YOE92$�M}��en;���He�zF�� �8m��S�g^`h�=�윇U��0��IIbx^q{�vK*X{&u�7�;^R�u�kF��ٕs}�t�a7Vj�a�w>�*ͼ��ls�U}�QOna����m�d�!h��sul�0�*��L	�4./�U�;zT�<�t��e^�}� �ح�W�����&���^k'h�!pRw��Yݕ!�Ƞi+��E���y�`e��Lf'�X5^}n���e'4�U]��f����m��v�v��+V�4�q����"!y�EX���jݹOc����o;ͫ[w�+��,��������9�t&�	��mM]:��
�\h��XwL��Ar>�q�vm�S@�ۗē�E��Z�v�兇��EӪ������I�}��F��j���	a�|;+�B�7|.�#�P����gҜT�m٨�	�hLHew*[��v���C�nDWl*�9s��gzV7W\1=�SqvgK��A��yI2���pv�� �.u����oi7V�ƗP��y���U���bkr�2,�)�un���ö�̱pO\��=�./KZ�����5�)���j�U���Es`3�5ҳh�x����������$ع�,J6c-v�iN����w��v�Ǌ���M��E^����s��uz���]�o;[ƥ�x��W}Vf���Y�u��0��gZ�gڷv����"]�Ox���|�1h��[�ۧ���Xa��t���|�κ'3�Cmd��
{[ę3��ˀ�̹������:��6VQ'(��U\�w*G�����bQ�̒���x���q�5��"��F(�e꧚!o��"��fw^�Z�^�|�{�v�j�#E��Ffe�e,���j;rR�/c�ֳ#��Ӽv]b���t<(��Y�����(5�0Z��scj���cXz���Wn���5�D4y����\�ё���Ѭ�5��s�B�ZX���:#9���EB��i鉉�AKk�F�Um�7��S6���Ie�U��;�긮���B�C+d��Gc���ԗ;&ir���'��#��ׯ�s2��]�@�j�f��&g-�՜����c�d#s�\
�6F�̸{2���7N	�V�2�S*�L�pR�L�6Gp�0�o2����="�8|��Cv���e����X���霵�7q�13
0��t���}�X�uKɮ��Y���l:���m�N�[��fu������&�%P��٪OG���*Z�ݡ�\��q�1�]��c�s!����u�e��B녫4�C[C��a��Zso��u�����E���jd`n���'I��iۃez�h�v⻷��cp�^��&�����J���د�^���`�]{*s��. ��XZ�Ӎ�fstu�Z�(!V�XT�uk9�&lu�Q�V�5W{��xɽ���u���qc�^�ߐ�2�j����Ŗ	�V7����>N֞�<�X��B����.��2���+0��e��4-�d�m�����}����d�ąh��7�ݽY��c������ܾ5z�0�րz�<`��b�6�=��3�p�jfjx�\-u �l��\�&�_p��,�o�n�u��MٲI΢����ĸ'u1���zk(o&i��n�kxd�|�cE����r���>���&�h�n�yԂVI�ޏk.�VE���V�*b��q�@�)WZ�Βuc��F,uP�@����gi+Z�����n���r�-ݷ����5��-r�#|��yԉ5w�(�X���#oRvx�C>�xeD�e��\��ǝ���b�r�J�{�W�w[�Ed�1�j�`����ӻ�짻|�Q���+��B�D���_fT�}Ւ[�ٛ:�vѼS,�o�����r��ˮ��Z�X�Q�gFd��ˉ]Ͳa��8z��Z���h�j9:��ֆi�A�j��Wor���ź��M� ��_�P$�	&$����km��i�CONi�@pb�gKr7=n�Vݛ<�Ou�ٺ-٠�m'	�k�3���	�<��;q�6"�۞�s�R1v�;�ڍ�7�srإ��$�q�Y5�7n4q�k��pz�!cMg5�ֆ�Dv��5��;x�m����[���o)ܕ�MA�#�k�*�lp�Zk�R�A�8j�Ǵ���]�8<v^N;�(z
��Z��=�9չj���ݸ��XG��݌=�]+ڄ<㛝�-�f�,\�=`Ĉۅ�c�#��vN3���:3y�2s�͏7������;�2w]v�ָ+
ó&�;��n�[nw&;c�qb�2�[�i���C�nմ.潹�ֻ2 �X�N<�������$�ٹ9m�i�İ�Xg=f:���#���5̡��%i�v����^R۱tr�vMڧv|&���;A-٦k;��\I�`�Պ�˨��;{Qn�g]��h{u��h6����݀�<�[B�[���nk<'L7l��u�ayr���ю����Q��8�4���b� 7#gE�E�-6b�(p�]W���ໄw\]�����n�g�I�=	�+�R��vl��Xy�2���=
�rI�jlx�۞}t��@��f���]����Zxn9�˴cn4���.�lY ����uu���ѹSF�zn�gn{5��N��-����v6��7j�4uw]�,:���*��Dݱ�ۗv2���/�����n�V�=�Dc�lk���Ypr�u�$�\A�x�v֗#m�u"WE�lp$ɞ���/��7\�!D��<v3�w<]eV�72�T��}�kgͩ�Z����V���3bݥ�.
De�xݹ뚍�����f�û������n���g�EԽ�x����IƳ�������0�T=Y�]�]�� ˛�[r��OY�{<;%�v7;�l�'��.�Wמ�m"[;=��������9���ts����CՋ��^޸���ǎݶml�+�C%���d���[R����Gk������^��S�X梮�ڞ^��$�6���Ǟ2u��0vv�.v�k���k���W�d�<j��[1u���8�f�૖�.��ˈJW��;�:�l�x�ݗ�j�����=R�q�yY�nn9�ݞ���H�y�I�����z%�''����ŸD��^:�ჂNCnyν]g!Ճ���%:��v˶��BM��W[#C�v3\��2�����R���spQ�'-���Q$����:7�rQ�����u]�v�z�D���g�1�v6#N�U ;u�ڞ�}5\��8v��Y1��񣇸.���ly���\��E�Dv�w ְ[�y�=+�4���1�7Cq�Ԕ�7-qŻe뇈S�c��z�j:HܛN2l�"���];�a�li�#���[���^]Wcn;j�;5�;��	ۍ�g�[��'A�w]�l�=�s�nS�esт��an�Qݖ�1:N�b����m�:��Q��ti���f8{�CMGX��x�)�ըF-mOns^�Of��1F3�M����ݎ�o8�Mt�غ7ܽg����FBwmz6j�yl�Cr���l).zMu�f��'^b����_;�;n.�3kv�ƃvg�YZ�Ѐ�Wg��ѫ�&��0+���:��Ra�=�Ձ;o$��x�nt��V steӉ�gv��㛭�������v���-:���=<��Gj'����ݷ3q��k��Nۏ6��ۭ�r#�]8�c��yQ�f���On��י�k�W�]�oY9Kv�s��;�v�v��pS�y\v�'�;o>.p�G��q�8�F����i�݌�܊�ϵή{"q;�ZL�on�B�<a��ڃ#�Zn/m��[�����W7�8i�//�vJ&E���k��s�w!'1�ۍӣl=)��ZdۨQ�]��(y_\�sS�w><�Ր��g���bKSu����<,&��N�����I�<��<��ܻO�^w,d쇑�l���q�g��ۍ��a���{h6tG�+�s���7h�n̢��3Gm�Ÿ�彫*㒗h�uE<te��u
��Ȼ	��W�� �2��@�1	�1:�BP�ug���}�1��W�H�f��6��\��Gn�rq<�n��;�"c�՘�d�6��4�,wm�W`6����9�39�8}u�]v���ݫ]�u�<�Gm�R��Z�{t��X�v�.�\ez���������;����sv�/	]96���\�n��sd�v.ٻ������ͥON�r�E���A��,$�:�
�Y1`�guۦ�n6۝�nk�5���\���ٓ��h�	vՄ�����ned�7�o],�r㭳�-؋��<l��������oE����l���u����E���q��
ku;q"n���ø�5����ҋ���\��t��9q��WG���Ss+�Ӥ��sa.�N�ϵl���1�#�Ԫs�E�^��/��{q�v�>^:�]�k��L�۬뢻��^��m�ܽ�,�W�9qӷNǣ:;���`̗:�[�rj�;��6�=pN�]�' �qzy�9ɷn��#���yN���g,�L���̽�u���E\89+�����MI� p� �\�8�2dz{�ajyc`$ ��ݤ�8U.�e��k��v�ss����ܾ�wkZ�֌�v��+���λ>}0w��F��ۛ	��y"�F�ݺ���^�f5��ܴ<;k�vH���K��A�'�ԗ�ɋl<m��G����ˮ(�Ml�kv��ޙMծsN�s�v�5��w��]����Pqݘ�\��nv3�ë���z���Vʳ���Y���[�=����wL�"��Ʒ=gn{Ā:��f�<n$n��+�sm=�`�f��[V���}�;s�8��k����=�Ųnz��v��Z�un7\N�9��E��F�T
&4�	wm�:�f�s/n�����`Fn�h3'�x3X�x��b�iOa��cv�eMlFy���<�u����;�r���c\fm0m�N��c��vM��2W�s��E*��B>�'@HR��Q�B�@~b{Ggʬl�̱v�Ɯ�[��A�؞�wW1��#n�:�\sԼ6�nps����V�y֜����=�g)xx�w+O�;[^�m�9�vN�\X���{��@���J��<�˥�r]���1y�.��i��uԽW
G[�(�8� 6�ۗ�I��E3��j����^h�m��u�d{g�W���`c����h�q�;n̚yv�Ʒ@4'=�.y�����쁻%۝Wck��n��u�>�D�p�t�Үם�sŃs���[y:筻n3�N�m��X�pk�e�Z��f�%x��%��������3���Щ���&.�ոXoO�����sn%�.g��Ty��.��qc�U�F/Yvݶ2�qpm���9�nR�ot����۴q��=u�.��T���j-��{2Y�H��<ӣ g���J������{lq��smV��n�7�Ɯ۳m��h1��&�km��e9i�3����#������8;y��z�:�u�'�'&��ӛ��X��{F�M9:��6�͞n �8C�Y�n=��8#<W���/� n �.�9m1��Kd�n_N�ks�Yw��K�=�c�;�K��
1�n����x94�$��	�&سk�U��;nٝ�#pf�ֻv:�l���op�m˷��6�.� �&��GY��/3v��Byp�ݹ0��h9�.L�h�3�.6�r0�\�������.�v�y2�O�^u�^M,[qa�5�u�1�v�n� RD\�y\n�m�����ۃp����G�NKF�w!ջ&z��n�Ʈ]�5UZ����;�o6Ĝ���Wfs��vu�x��.���	��Os�tl\�����n;.�u��.$�y��ɺ�z�����j.R�c�y;R�&��S���0㛟=�Mk�r%���=�uKr,�uH����g�'O.��2�=8��ǯp�q�,<�G^�,mXA䬖a�uNG���wG#���nnyS��R�H��㔁��x��X7%��'S�����.=gq���^�{pY����n��v��=N�6�IM���Kc�������v��.Uܶ9������$[z|7Z8��ݝ�0;�Ev�C�t�E�	v[l��k��h��U�x<]-�6��IY���;r�������J��:9��{F1��q�5�v��[^SL�vB�X�7rLᵂ�D㊁���7m�tv,v��x�lqk�=n�t�ǜ�OG]��tx�6�������Ȇ2���+�T����2��hBAۮ��nܛ�[b4��F-�v� ��
�\��x�����j:7��3ڛ=�h�p<��wi���6{)Y�r��7��y��;7%�>���N�uݞ�n�c-��8�z�ӫt��.]����9����s^�d4���m�����b�EÃy;�;�d��e����a�^�8�شxY-�Nλp�Mݻ6�Okr���ōZ9����
�Js��\���u��������۞�[n���܆g��g�P%�w�P �΄�uh���FY"���qW�=̘����{5Ɂ�[qı�uٷ�A�ӟm�[�v���c��2� ^�-�pN�îy���n�Lch�][R]y�}۳�۫+��oN��y:+�x����N	���{��#8vM���7>q�+���:N\�RnF^�b[�����s۷m��v[p�{j)(wdsV���t�I�%��v�q�F��F;��1���!��k��"�O�}�m���5�]k\y����3y��u��ٰwn�%��ǎvB���]�-X�}@��Aϝm���=��ng��7T�8�f�;W ���z�Ě�P<5�h�jS�+i�=>{��>[|���K�G(���YvZ��e�-M�!���	�`�$Q� �m���`� ��f�8�[`q I�!���r"e�ZwmZ8��6�r9�6Î��'	�� Q\��A��$�$�.S��RH���9fHYl�����Fd���N���ٸ���IӉ�fH��'%KN�*v�):!�"s�#5)��%X��Bs����'Yi��V��N[vm�H�H쬶�t"�r�R�[k��2�$B�ȡ�Ds�f[qZ,I��sgM��!Ci��)��e%Ë;86��&�D�Kn�$QGe������u�����}{�|�{p������;�7y�,��i6�Ol�w���ë����ƻ�A`�핧��y��^wnܑ�,M[��<v�/����n[n��wqH�9[%�y�x�r`:�K[\�θ�<�nN�����fٸۗ�1�vp��ݍ�lgi�.�|�`�UZ.皫�6�w\-���F;s����ct��͝��6]6y��.O:�^��]LzqǌOlG:{;\*��6ڻk\�כ��pqq�hD������l�N����{nOZ�h������A1�;&��q;��;)���گBT4��9��Wc��a���8��<����f���j�Ӷ���Fϑuv�;q�>|��z5�l�L��F޷�ɳ�gS�e���]�m�����i��T]�۴ˇ���"���,��=�jv�����R��m�^�-y�:�`|��ѹpgl�B�y���r[{|'{�����|�x��ӹ\��K�ì�k�ɷ��v�M쁷��6����V��<b��zzE��N��n���u��%[�=�"����8�<��c�׆��T�����BC�[�7lJ�[��㝸�0��=�"��V8*D"�c���k�(�g�y�6�99�c���{X
�]�ok��ΠJy�X�笶�j�η�}�m�n�E����kx���e��m˻7j[-��[�=���v�窶�t'��)\c���W' C��9�i_��eq�	��8�Vv�s=�8ɦpMq�6�v�2�a[*�����Bzp뮂��v���Uvŭ�lp�6N�ortjk�t��"��E������*�ЈB���McU`{2ǜ�-��ۮ��=3E�.���ut��7b!Cm��9�Z�bv��ذ��5�6d4լٺ��-�V	��"l[��qv�8S�l]b��t<��m���wf����j��Ź��۫r��:�9�@��1�(�^{^���e�k����۱��ǘ��ݵ�%������f�����6X@�>;&�c	���|8nW<ako^C��ǚx���{L�Ӷ�L9�{݃�?��u!��>��{^lk�{�,�M{6���d\&��Oq��s�yCǎ�A�c�<�ۅwd��L�3�sʜS��m�a�Q�x�pUC��G�d��A�s�S�� ���g��S��8��n���l瓟a���7l��ld�݃!��w�?�����'��k��I���w���8����l�'��P&������{�y�O�ƞ�a
�#tE�������Zk�2/^�k?~��͓� �</�#m*�
�o�`cx�_�����~	8i�	\�=�����c$3{y�	$�+�m\�HҵF�X�uc�u��j��[~D���y�~�NP�?>�GA��xbܖ=�[��'�p/hH�B�([>�^��N�n��6��>��8
\�lP-�����<UVkח�um��6��Ƈ+�JA��1*r�N沽�R`4�O9..^�_�>��Ң�����y��<i���ka]-��~v�ڟ/?y��~U�Wu�j��XWl�<׹�X�zw~\���K������=�\۸ܗ;��뢼��+ �v�S�����wUТ���`|o��N:��\��c��rd7R��9��C/ �Μ�x
��Z�P}��ޯ'w쵅��X����6FX�C��}��խ��kggf�V�^��'��|tӔ=�$���'�v�`��X��o��4)I�U��+o	�ᓫē&�7���w�nٴ��ʼ���UYמ�M��F�X5uc��^�����`�޻�y�Tc佾�	��`�H;y���ɬ�w�]MeVupD���c���[n۵����>�����J�&�����A�<����o��Ț4�*([o'Y���M�������6<D,�!��m�|C�"pmt�T����y�6G�^]&�1��|�I�c`�#�o7� �y��x���ɿ(���G�k�I\�����X�9���H$|n�V ���������v�#�a2��.9�y#�{�Vt��!��f�H�n���&�/�u_,�j Sy�|~����C����4X(P%R7D_���)��~$�ǭ�L�;��A��-*�rbꬡס�H�=��p��W��������@A9Ks�Rȋ��w�<�$�7�0� 흊��s7�J(�az!@Ѽ��7d��f���뱷iP��v�v�Qpp���
_]��Tj��$����X�=6w�dʩ��윕�����	���%��@���#�w]�zt{���u�nz���0A"M���*V�W��0͋ٚ����
����=u�덶�{6�Iɓ�t���a�q̙ ��{[$�y7���\~���,��KnbN��jl=�D.��O�����N�L��K͞��^�s��#���n�5��顴�B&����y�k�86�@�wetF�W)[��`�{�L'�����&׻}����v�qO�EcWI�vm�{d����)Va�:���H$ʕ��	�s�6X�^̐⧲���D�j�d�)�v���M Iu�\�nj�F��=^;q�wk�]��t�j=`��X���l���9]Y�@$|O۝1��=��V+{��@$�J�{o4r��[rʴ��ow���9��b}�;3�x����u�������)�|>-+��S���ɴk�-T���ߺ��A��a��)sd{����$�ɽ|'�~߳�������AX��
�ü�_,����a��A�6	����hXX�h!ڶ�3�z�]٫��j�� �ݍ�Nov�����Z�'6��
��S �o��uү\R������x.�n�G��WJ\����^�]���|V#�#�،
	d�� �Ե�x2���+���GLg��X2��57V��A�����R5��U9��ظ;��h�g�^���/v�1�ל�/cn;-��N�<�wgXNø�2��1�Ѫ;<�u���jT�n�����n���ܼ6z�{ެ���vݜ�[���B���=s��n��9��^��jڻ�`8�=���ʊv�J�I����6���s p������x��(��I}��Km��]�Һ1���R�og��yx{O=U�۱z�[h���1���M���� �f=���>l��X�T��?�lzt�&T�{�	zH_՞�}:9���	�!}t~���~ޑ�A��\Ǔ�����H�l����`�>��Y{q=ƪ�̈�����a&�xZ��M���I���m+3�ʕ;;� H$fs��H���z�+�yYvA�Ux{z ��Hwg�yQ������ݹ͂ILu�A^L)5}����SQ�PV d��׵��ci�����y��kN��7�<��9���v��sFs4� l�Ɯ�������h�v�5֧l�bia]V|�8�U��(�V�w�V�]�Wx�g��wgy�~$�U%�<�R���"�u��kt({ޞl!��]_���b��dU�nE�?R�>u�iwfW�bn������\ �'3^X���-J��]X�u?f�9�X�S��yGeI^1w��B���A$�zy���e^v��u�^Xڋ�ݠ>~�'`���6H�.��= ���=��A�E��F�Ă@�~$Ṟ��o4r�K[vʵ���w��9��u�{��4 �/�qΖ��׫�v�K��P�FN������U��EY�6}�}��׫cv���,��y�Tꀡ���X �l��y�i��K�?!�-<���v��� !�B�Wm����8�4��7��y}�h[�н�b`�u���s�O��4,���'�^�w�ka?
w��$�a��d?C��+F��뻶�[�� �;�i��q57=��I8�]x�	ގ6	/3����s�8I�ā�_���O>�O���$�F�6��
ler��*�L�7�j�{Y���Uנ���n[�;}�[�Z��^:pr�g��˽F�V���|�Q��{+��d̕���;y��������}�Н��(�����K�J�� ّ��$�ݮ7�?���>���1?g6	��ե3��
刖����^��������`���o�r�<'�T�x�'9�>$�oO0	�����t�E���uWj��+�<:����|<>we�����(G����:�������f���uEY��Ϻz��8�`����L�X�>_z�?q��5,��y��ȏ>)�1A�^�{���u[ɛ׺�Е%g���d������~��퍅�P�����*����n������'7�x2OQ	���+⶧�+A �7\lA#�tb+��6+�U\:e���U{�֮�0}��I�7�6'����D�B�F��f����v�T1����6��e�ӟp�M�;"��q����.��OVA`C:ƚ�sy=�GQ�"�V��IM�yF���ѫ^�{���=����Ha�{Ҕխr�$c{�0H���� �p���{���u���f��ّ�2Aq_�
|���O�<�'�;\�Nۖu= �h�n�����6�{4U��7��d���$H�S+����gb垔���$�s�a��*���t0.�B�]ڕ�,^s`vw{9zA����ᩞ��̾�������/���N���QVAB�����͂Aks���&����uW����;;9��$53��~��J��wuJ����=y�.;*ڙ�|���� ���Z� =�z����f%(��� ��PY�A�_TM�~:r���}�6L�!s|�<}��H��e +��]C�԰�W�i����b�����]�Z�b�t5��mi��ye��㫶r����z��8{�$��	�U���Y�.Ɠ��i�;��* ̿8RUV8 C�S�Je����v��p�I6��k�v�n��ݞ�V�Ύ�,uψ�z�r��M74&�g<�\d���۷kg�=b���٭��J��H���up���ډ�6$1��S��ۇ�}�
s;��p[Z�s��<o5�[]<��r���tyȽ]s�y�<��3Ƹݨ���K=�n$8^�3��k����m�v#�sϳ��.̙�`x.x��+Ρ���ˍǌs��"���K�}T�g;��P��ҡ��{��K�`���xO����6�<��P���{}�����
��ӒC�ˣy���_վ���+�/&u�26gn����c��Gg�u����B5V{.B\^F
	XWH�-�/۾$����Z}��΃�%dw龄�GV�	?oG̈��,LQ3I{3���ŝ�n���ل�B���$3�l�'������5���v*��={wvs2��ט���v�c��O&/�����T���~��9r��=9�`����M��sKδ֟�X�[Dj�\�U�cAȔ����/V��
d�ۋ�ߟ_����|
��#v��$���'�zt���2���$tͱ�~y�6H���v__�a����2��$u�(_���O�fj^���	��^+]�.�5�d�JDWU���s7���K=�����g���V6:#�i_uL*�Э.�뷥��{5��y��	9��#gNl���_\�3�t��Ԅ�R�b���`�e*�\�({zw��_�wu6��m�I������=�]T��*,^���zЍ%����G����0A=:sd2�:U���ų޿oR�t,��sl���]�@��9@�.� W_EK�oĊ1\D|	��k`�gt��2���Ǭ���}�˽����jg�8��Z_�[cf�x�s��{T��� �F|)Ug����-��w��9�G�;�y�H'�Aʎǟ�c�������@'7;��:��Y� j�����y�j��ic�U���I9��n�Kԗ�� _�6z�m����佡�G������=��P�|�  �y4���/uC�*���(�0�+3����^ӵT��YY��Ζ�9�
�8�S3ewN���&嗬t9k[����Il̲pT��an_�U���#Um��a���y�vrk>�T1ҭ���H���YH�<m�s{{�pav*���H�J��%d����x~m��ǘ���C>B�R�a�Ȟce�7��g(]{�P�h��i+�K4�wdUs̐8K��ܚqƦ�W�i���-��^�g^�k�D�<(`�q���7wtj �<}v���B�l�=�Lxss��ʴ0�5XA������|"k[����J��ܤK^*���kҞˢ�G3oh�t6i�U�ۄ��K�]��Y0*�۴� 0�X�8nr�"����7P=�$�Bun���m�KYۅ+�,R�Sa����z��v�K*�'k.� ��_-!ԫivZk6� e�$�XŎ��Ц���z�Q�;�l�=[F��|�ҧ��x�V�	�.�qִ�|�2�b��M笖�_g.�2�i��wY{_-�٢�k��K�]�]np��&b�	Ţfn�����]]�&E֎�UaK"�A���%����R�q�P�=�
�
���Wx1'�Ϫ�U5����\���Wja�*Է�S���H!tiwI8���Zޕ�,����nn*��gT^��#��`D��I]����J�`F��IJ��A���5�Λ4���K�aE;�p����a�-1R����w�%@ﴋ-��9��ԅo��bz�8W���"��vϐ�w��RE5a�?/����a��,�4
#��8�)��,�I#�):E���n�.N�"J9Î��gGL����Jm�p�i�&�t��rH���Iħ2ę�h��A�9"r�	m�6�#-(��"(��\\)�ܖb����p�u�H�N�`�!�9�9�$��8DY�e�8f( rP�f�P�r�RPQ�s���:���喝m���r
D$q�BA�\�:�mn%$����ِ9�N rD�s�%$��.)K7�I�E�$�rP�tN��h��I���ҁN$�:8�\C�9��H�-�qqG�IG�K0BD�pӥ#�e�^��N�� T�I	�VY��7� ��J��wmrJ�}yt���C�� ����_���۹��l�tT����*�d_�{��{5�������T�/t�$����;9�0s�U�_���߼��.F��<��mղp����<m�5�"vV
FGTREu@8V�l���{ �:���N�s�vJy��'�uuH�0L���>�&�a���7T=kMm����( �,@��3oD�[vV��_yz��H�h[�
 �W������~.s�2I����b��1�I��I��6>����XxEe��zO=��3��BXB��HQ ��q��'{;���i��X0x�MXʙW*��ڷ��^ú�LS��	��:��D��Z ^�[ށz���J.}+���S��w���W�Ь���:�׾h�=���iU!,D���N��,C���It
o��|)����t��'�@׻�dVf]�W��$H0'�h��q٢M���mu`�u&g�=���.IH7Pv�B���*Һ�Ue��{^�x�N��l�7���J~������k��26i�����Y5D�%xw��`�}�<�� ��?�I��#`����d'z̅Ӿ����ר��+Wj���v�;�u���� A�C�Q:sֵ\��+vdl�	���� A�-gƅ j��������T����^��$rs 2O�L���U5'��8��,_oT��/6%���G�������� 
��C{�K��3`�a�\��	3y�O{��o��Rʢ�y�8��`z��:��&(Ї��[>����P�6���eJ�͆鏰�Рܕ��3
�{z��ܲ����7�n)���W��H3n�-%���>|�m�y9���Ͼ|>N�q��%ɵ\[�7�1����,>�U`'C���#���mqA`��0� �@oB�/;v��=4fA����#�(���j:[��aN7��$��y�T�ln�-�8;\��;�Zj�Xz6pZ�l��n�e�e�8��r�O8�x����<�<f��&�5����vT����ڎ7U�W:��6k�-�CNN���T�G
�i� ��r�܎�|�򐫠��*��7���	=���	��H.z�]\
�O/o����0ɛ�͓�.��8N]��� �U`^v�е����@$���l�I�sްOK=\�����{%I��4��h��]�T
�k����'�~:n{�~$he4�d7�����}���3R�D�'a�����y�����½�XLF���`U�{��g8ݞ��~�9�H�vcl���(TM�^����}d�9����d?e�P^"#���� 7��A;��e5���ǜ�b[h�Ɯp���mb��f.�n��!��f9����68"��D*�{��eb"iբ,W�ٙ��D7��I����!uPs0wn��a��������U���*����kd��4v�n�ØU�}��2����"�{��YR_����4R��΅H�ֆkx=�.��A�ߕ/!�K�H��W�N��8�� |W� '��a�ud�(nq��0шe]!Ue��~=��d�M9UU�%v1�3<��p�I��x�s��Y�+E����N�旵�s+�N��}��-?=]�*~$��q�H�������$�)�}�"�	5X)�%M�pf�ϯ-������AΛ�6_.�k7���+�^���0�=ӹ��of�+���b�Wt[m��yy4<P����TB�Q[��Չ�:5�X�*��EB�5D���闕�D�q��$�����/z�w���<��h�x���Og8�~��YAP բ,W�}�� ݌�w/>�]��Ad�sy�����͟�)*h���]�X=�R"��Ѽ�UY��|$���$���|���o3���Z�=[O�Gi�^
�N����[K:�a!�Kl�U������-�����k1^�� ^��zT��� o>��	���g���#F`h��uDUYl��d�Η��/��	9���$�77y�Inxz�d�.O{����;����"v'5�繘�'�y�+���o���[�@���`�H�����F!��Q�W.��S��l���_}��Ŷ�ӻ8^�g��xc�&��0�6�;f�HvvÀ겧GD�~o���Wi�K?.0<24g���[A��DR������$�#�7�r��c1�����Y:k��8���r��biF�J0�9�w�cLQ�p���/�����h���7[������F���s�s���+��E���`FF9�w�cF�8�7��] �� ��5Q�3��k����/���P���4}h1�1^{ܣ��4��&�t[J�A�0��4j3�_wR�}��Q�#DM���ر�iD�iD�{���V�LV�Ͼ�'�ZS�Q��#G/������[f9�|�[�DR�wݢ��A��G=�j��l���Fo��)�+��z�J�ug�:����Ϳ�����<n�߮Z�ѯu��M_}|��*����w�h�*ܒγ����F�N����Zz�_��~K�Ҍ#�F0��4O�n䟡��z�3��э����������?w|��i}Z�[$�����[l�N4}���PC�Dh߽�R-�7w��^n�Z���CG�k��O�R؊�ܻt�`��6�r��7^'YTR�SuS悍�w�N�G4C�4�1o��ь�j(�iG�ʺ-�L"b�Ch���F4bh���g��2}���u�eVn�b��iA�ҍG��A����o�I��O�����&F�o;�x�G���{�[��{�@֯{��AAƂ8��v�L���Cj3���H�!��(�������W�޺_k�q�m��K�>_���Z4�7���m�F(#F���McJF!�=��ۓZ�}�5=������#AƂ���t�ʂ �Gy���9w���?�>������bb���F3}�{���f湾�@��iF�iG�{�,iS1F�D9�o��bF���}E�On���{�ΝbK����RV2���.3�	����V|��dh�v�H�!�H����=������j�#ύ{���e��0#Q��7�F5�(�Q�{=�Q�3�>G����"u]���Զͩ?Tq{�9�>�_Fu؛J�h�I�F�1A�s�n04^*̫|�d�S�B��ܬ�w��m�r�?�%��{��nD祕S�b��.�2n�9��Mv�鶦�X�9l2b<�Y0g�����٭��W�F�n���]��r7�;�>|6S��`�gn��<�0��cډ�َ�_l��v�A�Ό�M�WY�0vsg;��%�M��/g��ɮS@/'6�-˰:�ڱ��Ԙ�^c��#ˣ�QЏ�;��:}��;k��6��}cwiTqqojf��Û��d���'��2�mnܞ7h(G����1gq��DW�}�𬎑�+��\/����~�J�[�F��s��icQ�l	������s��k��m��;���U9H�����F<淣>�zoZ!��ևh4�b�s~���(Խ��fh�=s�K�s�xV�Q�(�=��-р�"h�Pg����b��Q�-���}^����.����\�%�o˟�Wi�B�cIm4?���wA���I ���QxA�n4�5����{������AL�����L߻��cXҌCa{~����D\>�9���JѦ!���(:}U8_\|�s�s�+���#a7�w�`�4��b-�����F�8� Q����&WR����eA�)�?~��E���w>5�g���>���;�Q����A��J>Mw(��0��=���e੄b�+7�F1�Db����Q�X�4��iF���2��ǈ����I�?|d��گ~~�&�%.��������a��@Aw%�n����h�8}[D�u�}�O�|O������̍��i�c�C`w|屮 �"84���e����y�g�{���)�� �Pg/���kQ�l û�F0��4w��9|}��>�N�m�#�}���b�*���u��?~;�DV��()��7r�w���� �=����o�;�1�<)K}q�c�G]�Qw. q	3NP>�n����?Ho_w����$�ඍ~���cJ5��o߿Y�dh �A{��R�!�"v��ǭo�eb'N���gu����!��[��e�R'jv�L�/w{��`F!�Q�k�E���(�Q��|��z�O���6���4A�1A��}�1�F��(?���z��Mi��c}\�v�ZԳ��ў���J��{-�ƃc�DR���E�$"8�G���A�!��~�n�m}�����u�e��O%ƺҌ#k~���4E��c�/�ϛҴi�ƈ�5��Zh�(0�Ch�=�Q�X�����a��_]���FYg��[F!�q�r��YPCb�߽�R1�h#��w��Y�js_>�:�)�^�9�l��TvZ�8G��3����Ϫ��ߗ���s�Un~�.��5�o��F3��ҍA�'k(�iS؆����э4F���~�ٹ^��7s^��s��1��9�o�c#�Q��;���I_U�7\��P�ҭ%ƣG/��1�s����_s[��e�D�Db��e �-�5�{|�cX�Q�l8sW�{�{k~�a�(��N|k��}�i�1��;���[E1�&�=��k��D" �w�[��K����~�,�����������M��twQbWO��E�����<���ܺ�\�i��W�v�����?�UW�}U�=߫@�#Ah#������lC�#���[{$2��V2�)�<�*�=��Ql�~��Ͽ>z��{�������cJ�A�1�{��-щ�1���ޢع5[�o��icQ����򒱔��)��g�=j|kL�_Y�dh��yA��A�����QlC���/^���?o�6�h#��oփL�bP��|�cXҍA�A���z�a�h�d.vs�~��9����i��on��`�{vg��뛱i;;�w\��,V��Qċ�795>&��{�N9��jO���i�ɢ>�wt4Sa����|��iA��6o�������^��7���~߳[��A���AeA�qDs��)�/���>L�h�R`U�ۢ��j&�k��_�|�_��o�J�J�)����DG���э�#أ3���,L#J5[���$�^���~��V�����tR�Z�C�k��˵��1����}E�$h#�ƹ﷾�ӏ�|uY�g�d�����#�ҍF�a�w����!n���جNW+ϖ��o�=�(}�}������q1u0�PF��s(Ʊ�Q�F{������	�Q�|����Ŏ�mge�̾OzQ�>���2F�ef#��X�VT��_��-��xD��V�
?*9<h�Ë�.�n���ط�k�7w���ꯐ�~�Dh�}�R-��G5��߈���>�v�L������b`F!��r���0�9��ju��LCh���e��р��3���,F�MF��s�t�����{�Ǯ?�{1z��`���RF�t�7���N�:۶'c��b�	�GU��}o���R+Z�~^`y��9���b7�z�b("1ɾU�
b/��N�����-�~��H�!���D�;���a�Q���6d��d�J���h��[��E�A�b��}��=z��g�h���GF���203����24q��7�U�
b��s[�r��v���)��G2�s>���M�h1�ř�r�f�M(�iF�ں-�l 1F�F��ݽԮ{잩��<��4D��3���!��m�Z�-4�~��.c��'U���Ic#Go�����V��4�") ̢߽���CqN���S-���L罾R1��9�_v��6����a�oޣ`�!��7��ѯ��N2i�1�Dn�����b�#F��w�15�-{|~t���g>�y�i�L������Ch �}�] �!��9�o��x���מ־�MN?�g;��t�q�����������Y;���ZHH]!�o*a/hY�=����	TG���������3�!���f��(ZX��x汗R^P]�1f������0�֪���QG.U��SqΨ-uK���lf-��]�m
���e�Ki@K��G�nD��,�^�a��t����t�bڽŐ�gjS�y�O��/*B*��M�]���2j2��n�y��L72��C�K���hur�a��M�_I;j�#W/�>�K����Ε}X�i9a.5�#ܝ=��G�<�U�a�@�"X�څ���;uwx|�m={�H0�H/}ne���,B辥t���XI���c��2:ُ�R��ww��%kd���P�j�X���}�[���h��j��_b�����oWj�5U�9˯���	���+��:�yh^�ۭ�6��<�����s�LvrN���e���飻p�˻�9�]#ר'{�Bu�iF����	.8'	����˼��rIn�]�NY}[��ց��e-[ا,#5%�v[W��,"��
;����oB��(�J65�	gt��xT���+h����`!8=�G���run������=�nӳl���&\�/6��:���U�������_�i%�d�l�O��fVrmMn=����k��f9����l<��Ż�_���n���Ð6oP�&�9B�N�I�Kp-g�^b�i(�S]�j��c1ە�A�{�W��A=�t��n�g
����C�1�[���3����RjL��B� 	�!:��nE�am�N�,㍛��$����m�9�
r(��ȉ"�" �J�H:3��XqfIs��'q'�H�I�[ZR���$���%�		�Q)I˔���tm�m��9�I"�r%$���8���)9:�Ӈ8�9�'Rs��#���
B2,�.
q		�p�!m�#��:	H�f��BQĄ!G%�۔�Q� I��!:����p:q��mb�Q�,�S�t� S�B�P"B!�GH��'8�D�v� �':��p�GNtK;�+-����,���t$�]n����l��^�؇�*H�"���o�
�Y@�B�낉nbU�D2� �T�F�D�.n\i6���s#x�=06���g��=�皖�{��zq�Z�A�/��u�5����Z|���(;Xhk��H�q{`�X;c��M]���U����M=sʌ��sn�tG;��v�嬉��1ۢ�xK�כ�,6l����{Uĺ�%sBvB�m��cVt�Y�/k��H �q&y�U��vB���v�a9�c��h9���5��Sq���9rr��U�%k�#��۳�֭�-�V�qG9�mlu��5q{\{u��K�˭�OGl��P��a�v����n�>N�؂׶�<85�W.��Ś����vgr�0v�z���.ׯ!���9g��g]O3g��n�ygan�r�.x�E�^���6��9���n��W�X��15�[k0=t9�����ٹc�ۛk�śsrc��"\�v<m���`���<�fM��)��I�wZz�F�D'\3 �s�1���b��gl�I�Bq�\�<ˬ�KX�u���PK��r���m��C���'ԗ3�ۍ�#n�ʈ����gs�rv5���6瀁31�aWa��6g]�{n㱭M�1��1�r�� ��q����B^��<X�
v��m�v��\��Lv�[gn��Nd;y���n�:�^M�uŮ��v2[=�ǣ��ɹo��e�;r�x���kS�p���^�\���cn�K(���:x�U�'/o]��{l���I��7
����������t���v�[�+�p8�N^�-��yi���Ibꎕ��n9��[=oo�wC��E�='j��K3=�'�G[g[�B�\�D㵹��5�۷!��+�;��mQ�%HGk�v�Ts�k��� &�;K�l�.�"u[�nwg�����om�M�p�U[�3�<S�����p�ۘx���פ9vڞ������Y�|u�a�ڞz��F�Aʱ�j�Eۚ�l鵤ݛ���{�f{&�>K�y�Z�y�a�۝�����[j��=���E&��S�����G�;�z�ہ�\����<ٞ�'����Ɛכ�ѻ���x���tmncb�Ƣ�6nR��݀�ʎ�}%�3�]e��)���%�0���l��v��muuG%4�9.zqEq�f�z8oa2�5곝�c7=ֱ��ы�T����F\����5��w�n�s�Sj���v�&�E�u�m�ثn���Lm�fyɓ������9+		(����%���K��I���A��*豥l#ah���F4cDh��*���G��|��}�o�c�X5Q5�*�+lr����i���3�}f01��=��<h �_)=\�d���X�����ƾOh_!�ro�v����6�3���HƱ���o��7��w���1��O��2|A�����h�E�F���Ƌb��F����"؆��F땻�Ok��u�x��#A��=WH-9I�{|�c���|=�6�|1��i��3g��1���{�[�Uk�6�4�Q���豥lCah���F4`� ��w�[��u�u52���M,j4��o��RV2��G��־�j8�՚`X������48�I �w����%^[��O�݈��A���AL�d��{��#���(������`�/Z�s��ui��������do9��
�q�X�#G^�[d5�vu��)k�$��(���rv�����m��&��w;H)���#Fw���4�5����1�������Q������Aۂ ����F<I���ǲ~M�PI$���X����~��c5J5����oҾ�ʾ����q���Wq5����w��
�(f��(�l�CW)���R�����:幪��k2����o�� H�/����AL?1F�4M���hƌh�h�Pf{�}F1`�1���~��W�뽮7���^L�P�98M?�>5�}���24wy�R-�lF{�E����G	Z�u\����S0`FFh���R-�Q�4����z�a�#�i~on!7!$�gʿ�?�߯9���\��y��1�lCh�\�XҍFC#��z�`bdbA�󕔂�ۿw�f�8A��)�]���m��c�Q鿭3g}�1���F�j&�o����V�y�9|��߾�
0�b�����hƈ�6(���}F1c҉�ҍF���ALV��ҮONOU�M��V��RX�_� �l�����І�k��T�n�%�@����w�~t�uw��LCh�swA�b=����"H"8ro���������o��]�t5��z��F1�Q�a��}F0��3
���|޴FM:E�`���h-4[a����}���Y�e_CM��Q��4��`FFo����F�1��YpC������s�<�?߾����>? ���NWf�I��ﵧh4�b�w�Q����A����YH)�l-1F���sק�?ǟ���)��J)�I�LgP�"�v�)�Ky�����L6n�m�{]/��y��I;C�7�j��X,��4j����~���$�W��_��Dh�D`g���E�`�4��iA���n���K;��x�+���K1m����3پ�v���jq֝5�4�6#D�o|ߨ��$�#���.z��[-�h�}�R-�w�rs�j�}��Zi���P��Ѷ�9$�P�b��z
i1��w{�]�Xs]6s��C`g}���C#A�|�f�Z�!�"H�w��#������sُ����N�9듎[g�8�pq]�=]�7�V�)|%���'.
�J���w�m�nQ���ƿ5�����f�Q�o���i�l 1F�4s��)�6��\�y�LF1A�]�Q�X�4�Q���r�����ߜ4��Y6.�F��!�?ݞ4�#�f�~��쭁���E��lC}�֐S:&d��w��#ƔbSֹ��`{��Q�Chڼ}���|޴FM;F4cDu��H)�lV�4g��R-��Q�F������g5�����l�1���|��
b��?�~�u�Ƿ�C$�{�M��rB׈4�����c/��{�}��@�Q��J>o��
acah���F4bh�#;�z�b��>�;��ʝݗ���ݟ�g[�@@
��KZ(����#Po_AN<���]�~�۩���c�ܫ�����s�� _��_��҃Q�^�IZe0;C���}����>������y��`�1@/���/7�����k�;����׹h4�L�6��w��#�iF�iF����(��c&g݆��g�|{�����!s��sƞ�3���u�Wn�����؂U��_��P!%�~�i��4G�e��F(�4s}�(Ʊ��C`f��Ql�2�������h6���e �PCbDF������|=|��ڏM�h1�ŝ߹F3��(�9����_Newz�}���z��iS���;�o��hƈ�#f��Q�X#JF��Z�=�z�5����Q�z��2��ן����oG�j�bG���<b$7����"H"1�YV����̜���U�gd��{��#�iF�Ҍ �7�z�a�Q�V>��sG��z>ӴcF4GS��	���5�7{Db��1D0���R-�l���[�q��=�V�����r{=�u�؇��}�F<CA��3�s��}&���i�����f5Q�o���-�L;�U�ݝ��]�l41F��~߭уDb��}F1`�4�Q����n������ɻ�y�7��-\�S�ڙ�r����v��є�d����<�ц��Y]/c�[�������2�֐c{��7r��}C�S9�I�7]>�ܘ�w���@�߲�����ΑE���<;c�\�n;%]uqz�"�s���z��ku�j��U֞��OL����9�)��-��vCkB%˓�f��FzU�wUٸ�3��8���"s��ܚ'ő�1v��5v��wZ�bw4v�6�n9j-W��=�F�vN�7�� �5�*cw'J5��q�Kջl��T;^.�Z��`I0Nu6j|�a����.ͧ��:�YnNvs=�ݛ�K<]���]k�XDV����Ю����_Ě������؈��E�"8�%o��!�!d/��t�� ��L�w��cXҍF�`g;�Ql0b��_��P!,�ϖ��7�sZK��!�Vd��aK�Ε�m�x<�_ez�Ɣ�20&o�����F�'��9[��lC�њ�N򶏽�U"�F�8e��_1����ZfY���c10#Q4�Q(�;[�ƕ0�Q�m:o�ׇ���k���4Fw��ŃҍF��s��J�L�۲��ִ=hq��)�c#Go��o��;X||�w��6#d�^���؇�Dph#����A�Z`FD��A����F5}�[=���ͥ��F�ߨ�Q������5�������0h��s��)�&�m��(��iJ�n���Mv�{ˌ��c48�=[�PC�D�#��r��Cg;��s�=����Ϥ>"pv"�	�6�pp7c�,F���K7S���]�s�е�i��* Z�|�k�_w}紶��(�iG��� ����D9��-уDh�f�w�}\���_3����b��i@j4�j7�V�+l�P�:�H��4�MY�Ch�w7A�x�A�#��_k_zj��~�Z:��k�#��������r�)v?2�%^��{z�Z�y���YTˆ�U����^���ϯr��^%wZ��_���5����(��Db�S�kv��������)�J5Q��x���j�Six��iq�ƾ˫Q�o�b����H�E��kwAcE�F�0��{�cX�6펧uu��O^{5�Ì��G�kt��pC���{��x�Gg����j=7���cw~�����]z,�~���:�6�4�^�E�����!��rэ4F����߽�1���?_7_\x<��[�(5��J�lW�e�[S��\Zk�����������!1�� O������N����q�����MqM���S�l�g��r��cJ1�L3}���1F�Z�ݹ�ԟ�_mV���
A����
���;���<���=3�4�yA/�����Z���~��G�#~����F(�4g��Q�c�����E�0dh>���W�����P�u��ALC�A"#9�r��CxV�9�$���>�Mi�2�.{{��6�iF��{�����bT��g(�4��b� �"߷�Z1���6{��ŃҍF���S�߾�������_}Ԛƒ�&����*WEK��ѝ��A��lD��}�/ �">��?�^�F�����OH1���{�	,��+�{�{���r���T~�oۉ#Է��"���U�^��5�[[�;�gp�a�^8�K'���Y���>�UU�� �~`F!��w}�#��6�?s�����D:V��>�9T����g�����>�)�~ճيf��Cb��h�WyH��5d`g��Ql8�A����A���Ͼ�����?���~�n�lCy���_1����ZfY��(�c5Q�ҍ���XҶ�J��>���^��u�m��)ѱ�4D��{�-�҃Q�������[���۽k�u��?ܩ�&CrO�����!*l ��n�ױ����{HvgZ4 �$��������k��l7��!�r��Py�A� �;�-�x�"84��VZ
e�f���9&��^�?�kn��R1�iF�Ҍ"a����ch�����֟��3Zv�hƈ�o;Ahh�(0�]�q�kU�>����}�6�4��b�=�1�m1��X\�'���O{�����u����>&�8W49�$��oӴe�{�ߨ�!��(�6���-�l �D�����3w*���:�6�����Q�X0�Cb}�e%i����o�{�k��SP�՘�6��st�ϧ}O��4�"�e�bA�nOv��S�l�L�w�R1�o�{^}�u�>��i�@�	�Ya.���e.y�D��� =6������ȴ��#݂V7���x��u�����}�M��I�m�ɤ4�~���X�ɿ��#_�A�0�-|����T-�0�Q0��~�cKZ���Q������X���;�Ql��A����ALCb�o��R1�o�f��j}Un�_x~z�|M	�Zƙ�Ʒm�����m�۰�{=��b�Mb�@�fs��C��m�����A�xb���F3j4�Q4�|��+a(�Q��o֌bE_{�齣�/�]{{���iA�҉��;yIX�`B��Ya%e��)qi�����k�K?�b7zƷ���{{�h�AA�4�s����l����{H����(Æ=�ߜ�+]ϟ\׻G�y�4L��o�?�Z#5�h�!�Ogi���6���GF��������^�/�=��q����6!�N^R�!Ⱦ@|�����7���(��2׈4�L^���1����sz8��6�&�j(�w;E�*aah����[�,h�Q����c��񼏲����4��(�Nw��������jZ�����24g{��h"q���o;�QyM�~������4�7�g�h4�`FFh�g4�j�Q�4�ù�z�a�h��o�_H�5����&�e�MQG�i���d_�#�5Rjs�z�q��|@�xPz�k���ap.U˹n�1�����g8/{���/�_%�f�Ca�
�Cꁧ�YBp.V�cV�fƋ���E�vܒ�Lo;���k�"�]2�suջ�4\ݳ��<U���n���ŷ=[���Wj�����X���k���CK���3/U����r���ξ��M�<	ìm��2m��T��m���-��mb9�ą�gd ��=��6Jx{y�`q����<���gtf5�ֺ�!s��T�N��X"���u7p�3�W��"v�uN�a�Tם��.�I�]�7?_��w���p��������4#��n�i��F(0��wE�m(F���[F�/�o͓ۜ[���k)���H�3y�"ݍs��f���c�SP�Zf�}�1���A���o܇������v�i�X��&w=H��#أ=��h�,aPj4�Ϸ�W���C�瓚�K�����Yz�O�$ѡ��YLdh��t;h"q���{7��xA�n4�����9�C���|A�!��4oy�"���6�{7�ьCh�3�p�|���q�ӴcF4GS����xN����Q�.��Q�h�U豫iD�b���!�8�D���e ݚ��js5z��bP�C�O���i��s��R�#rפfؽ���c1������+(��0�������\�p\a��4^��E4[Dh����E�cҍF�MC�w��|�#� �X��Ε�jt���%#O+���gl�vwn۶��˸7e��c�c���;۷#�Vs|�����QR�^k���9�ߖ��D$y�v��IG竽��,�@�����Y⶜?���F���)�&�j4�0�oݣ`1F�S�3���sZ�_�4[D~���1X�1zΞ�a�z��޷F��[̩m7��Q;������FV����Tv��N^�{�!Դ�u~z�i�b�-�[���������h�G�+p]U!$~h�z�~M[J5d`Ngz�`bdh#�q����T؇��w~��|F]sH�!�_o=;4޾sSP�Zf1^{ܣ��6���k(�Ҧ�0�h�v��rk����LCbFw;�Q�X0�(�i@j?N�RV�L�_��,�ꩊZ�g���������Pm8��=��PO?'ԍ.ʩo�G{s$y�\�B�D]�(��|,���yxH�WH��1�&���$�[��s_x%�}�'���:($�6�5�Ǣ@�gN��r�E0�v�ehp�����m�R(�r�=�7��6��ۡ�s__�A�Q�cw�����đ��j�6��Q;JV\Ϟ{��ZL��C�ӓ�~[�����	�� =�Ch���z���FY�8:E
&�ɺ�x�J�| ��t�vg@��\����e�{;�t�ƉX/m�0ڋn]��e��(M��̍e�K3��j#ҵĂYD^�4jW�b�x��=۲U�h܊�&�-뵝/��";� ������Ռ��f����1]G�������M��}ӝ�C���s��vh\:���O�of�y�b�9�ǫ�3��yt_
��)��kkv���3*+�'vr�=����'b0UV�3�8P�Y���̔6��HLC(�ZO����xoJ�#�Y��m� *��Nuʷ+��j��صj��u F3��j��бl6��0�D;�Avź��e��Cd:h���A�t���Ǭ�J���ԡ�\�9�.ܟE����g�~��v{f�[�X7�%���v1����5� �bಔ����b�Զ��|R�X�I�(w2Ł]�����u��J�9�w�L��c;V!���壌�N�& �u��IL�+0�a�\�/�SEYzmCWK�wR�[��۔.�T��s:΋�ܺ�ɚ0,s�t̬U�s73GM�w���a�5�m�+y�7��I%qU��$˨C+V�9��Y��Y�{kl����[�h��ans+��8�[��r�np�1\W����q�)�F9��Q�͎�v7�����Z����K�ejWPQJQ[���;lS8,�*1��W��2w�N�n��9�C&jK�)�9�� �62>�n��X��k���?��*�n����_����[XB`;4$D$�.8�BP˷R���p���6��ېSm�$D�N�#�9� ��Bۑ�J�@!&dAˎ8T��D�Y��p��m�l*v���&a����	#�� ���� C����,!À��!"#��$rC�"r(�:D�:��9�de�e!B�wNt��s��;��M��S��&�)�Nt�tB9����$�@�NE%�6�I(��9$���J��S�mhB��)�$�8�s��"!(s�N�m�:q�\�m����Lc�������ڋ��Oߢ�W6^�C�p�-��{]vp���w'�W��Mf�$���g����{�²���y+�S�&+U�ʖY�Y�f .�1|9rHPI���Ͷ������>���@ztT���&=�u�?y	{�7�Р��w��+RE#���IBq�޹nn��g �h2I�8���g���j׿�V (>|�
'�:�]/�1�A��@v�%�h��8Hʺ��寕h ���U�\��[XO������fv�IU���/��OT߬��g�Fe�]o���!@|'Ort ��O��is5�Ui 3^��>=����R6�n�݊i?9�����̹�z�g�=~$��� ������~��m/uqHZ��.��w��z�[� ƝZ��.�9���*�_JsC��r)����b�f�e$�?%��)%�Bo�	 \<߫~�o���>�z�i�MA�w]�F�$C�����^�,`�14w?\���	'�~#��𺳞��ǣ�˽���MB�C��M���R���Ys ��u��n�ګr;��l�n��R�;����;�?��9K��-�X+L�c1�{ē��6	��i0���"�l��X��٘��I��@�{ɏ�7"��C��zr�ۻ��s8��WaA��ۯ=��cò*��u�bU�ye��(�5�A����C�`(X7wwB���fo����I�m H;���� ��W��6vz���n�����0H�4�kEѫw�fU����g{��d�U�+��l'���`���������Vi���K��u�ۃ����)�A��_!U���,�!����u*�َZqX���s��h��C�Ġ��u�Mw{V�����I}�vAtvJ�9���b{Q��b�z\uێ��f���nՃ��[s&Cx��Z�܅ƫX������XR-�O[��qݷn9�������oe�&�����'A��q��apO�y�����&�ۋzz���:�	�K�p:a4�㳛m<�<s�l��z\�u�ݹ-�(9�!$�p6:�!1��9����q�g�Wf�q��ѫ�5g���MF۷[���gW�mۋ`�z��B�u)�tr��\��v��^lR�ܺ���~*ՠk߾ג?�0��Y Sފ��ׁE���u~�sW�Z�<jQ5kv��k��{ZZ9�yx�^�q]<�2I$j�+�gv_�$����L���E�E��к(ٴ��Ϭ|)��!Q�������|��U� ����!?+t��B�V��=�5�drmu�<0m���<e�Y ��t��?�{��z��@�x��fx}d}B�!(X7WwB��sۄl��OT�ec ��{�B�oD��������n��YJ7������|���ݽ<�.���ODZ0�p^��c�#on"�
ZY*�߅߽�U-B�7g��Ή ��'Bk�9�¸��Y�ÒU� ��D���]ee��8@��v6	���K����W�d��*�֚�V�!ĝ�53)�8BX�ڑ�;����V�֙؆1�>�v��;o�������ƴy���y,o��> }���:�﹔Pڿg�v6���y��oYG��I[3eR�Zݭ8������o�?�����V*�N�?7f{Ă�����E���t��^`�װv�7GN��K�o���=��#L�^3��w��W����-k���N�iI+TUX�-���@��f�Õ:��� }�� (����s�κ���l�԰[)%ԩ ��3ŭ����v��������n6z��r�����P�р��%Y&���U���}��'��O�( +�smP�]�A���ۥ�_�Tk���1�]��8�eR�i���i�ga�Y+�O����|I;�kd�A�.xX ���':yog����B��?n�޼�a�L;s�� ����(Qf�n�u�y�9�S�VZb�.X��O%k*�����Ev;���h悖�6_ڻ���{|ͼ�u��n���{w3�}|���s���m�7���lg��z�Y�4���ZqK4��kw�<��ּՊ���:
��o��N�Q�;����'�����+�lR6m6oS��Oϒ�����KD����'@Ct�_]Fk�x��k�+�/�+�ѠP_W��Z����v�v�]΢yk��˷W]V����0s߿pn��Ȥ,]uw�ɱ�Iuzz� ��_{�n�u}�\��'�A�<(�C<q��岊�����Z�,�ߞ��]��'�:�C�oJ�������û�!5u��	���.�q��eVV׃�q������rD]�ypC��Ut �5���L]B°H!]�z�����7�J����}�D�L�=�I/:s͠xP���}��S9��ˍ��[T��.x�V�J�f�u��}F��w��kh	f�R�j������[�����y���ryI�����ַ�Gڌ֛�
W���?��(T����ϴkWS�ec^$~�}�?�v��9S�}ڹ�������(�%��w��J���[$�9ܫ�q���O�겨XJ�V7���X��u����3��s�a�A2v�V7/.��{�j��|\}�?_���Y������v�$�]w~���\���D�L���I"N�l�v���F�7�����x��J�M]աv��ݽ�I����=�zuz�&��5��H��	&I��"G��6�,��ޓ�/r�֯C{�m|O����dHޛ�?��I}/�.�z�_z�}͂WH���,*� �y��I �O
�C՜zm�h_M}��E	��0 㺯�y�D�MrY�k��L+�T�e\`j��͂�:�U�wuҙ�=wt��u�҄Zt �]/��$C�r��n9�J�?�� >���۵&�<m9s<�X��<�O\���&���v�,�v���ۯN�7'>�3�Z�{tM�h�t�������6]�糺ǯv2>�r�}���=��Iv�t���zxxWiݶ�����w	�Eλv�'>Za�͙��tqc����o��^_��#���x��p(X[��C��A���/W���;��j�K���C��y�E�5v���m d��9�ݺ<���j�v.����'@I�䓊�{�~��C��Z���w4�{��L  �^�UBy��D7�w<�}9�۵�h$ER:���ޝ؇ʻ�K�Sb��o`d�N��� �ڤ�7ے�p��g5{�g� �gNg�k+.��߾�wF$�S=��i:�vs��r�����Iǽ��H�S<(�$Kj��F�Y�l������u�fq[+� �q|���aT�Ws�6�����6րÛ�������"���5d�J�Q=s���r���	[ӛ�D�1�=�����7��y��r����~�rR�ӷ��8�f��GnaNh����m6�n�~~��\� hڴ�n{� �5L��?v��g�5�\����l�7��
?���XP����M;۞�l��ǭ���k[w>2���o���(�K6���c��[!`]��V8�	aF�}y:�q�#u�D�֧p���՗eH�X�/���A��s���^���M����]��q�~�&k�lo�s�E*��U&�7�qx�=s����;sj�'Ğ�7�~�s�ǗS�Tb��Kn������no�{�� D^������ �s��J�[��`�^���Ė�Uh݋�M�y�k��H<�g��������U���Āz>�2~$G;�K��~��w빹���
�I�VM���N��FU����P]P`ժ�o݉�ͨ�m��p.w�H|��2Ds���ޘw=]�xo�Wq���x����O³NuY(P�+�[켍�n���g�{��� �������7�����*�~o�]�Q��t�V+F��*�x�������	��A�K��X�7�߶ǈ�wF���a��ms�"���o�]q.���w��m�W�R�d� z�Vr�U�����^�]��	"]k'��7�����7{�ݺ���H�R:��$�N����{l��G��q�?2A'�L���c}�4[����b�[���Uj%�Z�;���}�UY_�[��x:�ͲI��������9�)<��QE���X�*�W]b���nڋ����v��ı��Ѕ �2��"i�>��_�ȭ�Uh՛�Z3ۛ̒9�̒I���/���uTE�d����m�~1�f��G��Q��%�s7)��w�;�m�k$k�~`�Ojs�P&��E}���S�ult��'^v �xX�[��Hj��ݞ��+/n�b��	�kl	=�g��.��+DҴj��
��ƪ��l�g}@��L  �^w?r�er���n���k�dR��6귖�Z�Q�\����M���8oyԾἏ�j�
|NM7|�Sb�����,�M��H9��^z���ԟ}��і0n�x�_X�������@]�4��K[�ӱU�+����)=�O@{��w�Yъ"6ZR�kr)�ʙZ�&�c��h�Ÿ��ˉ�'.���g=~~��?���5vk�����'�OE3$��[���C�s=��������瀣C�J�!U�f�=�� ��5�P�n��� ���^��Gk�o�~n��{ʫ}Sh�L][�����Y(���Q�����ϙ�=��2�g^)�f+�&s�a��:��B��i]�ݏ���+|�}\^_Ă�vxQ �׽�� ��5�o�滾�dq���ٯ�j���p��D�_P^�F�	��:j�o	}|���+�[E ��o� �zsn��Vݞ>�b�����+�Qo���c�4��[�5b�Wܶ�aVe�`뮧R�ec��hw��U����ا{��p=j|��k��6���]��4q��h���{lЯ@J�6q�'</i}䝃1kT.�&]1��]��ᗂ����7*]���3�F!�"NxU�L��]�
S�u'���7kg���� �mM$3�`AK(��s.�ҙ��nE474�����ûrъ��Z����y4Iyt�ҙ^��.ލՏ�D�v��h�*G��sm �i`F��|�>���fgɀ�<�`��eD4�����ޱ�k���}��]�O I�c.P�M��K��t�ˊs�{r�Ư>��v^!ݜ��q�t��8�}|Њu���H�ZI_&_¤�'*�]{L�ih��%ќ��÷��7s0PX����r�^��,���<K6P�g���`�wT�/N�H�w[䵞w�R�4��L��I��im��.�4�{I��V���Z�wY�25�I��2@��]Mz���2��m�SX�n��G,�u�h�ba����3`�^v���-�K�z�t��]uk��Ō�s.yW��u^����5������/˱�b���6�u���3x���4�a���h�y�^�'xp��ZF�RZ�\���gq�(]�#ʐժ1R���y�ѥp!ٕ���7��Q�(���ʜ���51�~����|�W���P�ҋU�����`�̫��R�F��DM��B��р|���Y���e񾴮�[���)�+GT�:�t�G�Z��m�W�v��{��gt�᭓��R�mC%
 �!'Qp��98S�D�t���p�q�G'(D�Q���W%9Ӌ�[�	Þd�p���@���N�J':@ �N8<��:p�����$p�$m��Ml�QI!G��IH����M�
rG���,���\q�DQA{h�:.:�$�7#����������
(��脤萸�;p�Ns���,8)	8��R���(�;1:"���8�Zr9A9ː��qs��C����� D��:"����8)'8��I��rr!fe�Y��9����N���9�'$� �ҒTp(�%%"��QDw�>O����>+���|hz�۸|��N�XM��<�����s3�
�9:��:����Ӹn�#�.���[�n6���͹��<��6��x,�9��s�1�qc$S֦�.�u��X�m�l���ֵ����=ێ$������p�n�z��;��n���{<rl%�=kQO�H/k{/X�˦������Dg�sշ�ݤ�n#X�x�ʱ�Om���_�F-ڍ��]��-�ع��O5�/h�;�9�&�Sfٶ��٭�Z����9x�Σ+c�\_���o�l����t�r���M����:��"��p���a�"���\mcl�$=��v���{Cî�Յ��b��wj9���ɸ�C2M�	���,m³��]kL�β%�9ax�w��N�[�����'j+q�9:���Z�nݎ�r�E�8.��^�J�<v��P�ڜX�Z�Vy%룙x�gp�{co�{���������n����q����w����,pg�,��]����z,�GW0Gm魖�����a��#�r�n�m�����[�6+�|���/Ͷ��)ݝ��hԷ�]ۃwY�l�î�����G7.��ENL7�0��t����Vֶ�#=��k���:�^w�%����k���������mn�k�������pq黱��p�&���v7;<R�ӌr����^�Ӷ�f��z��9m1q���ɹ��x{�[v�m�v��=�W��������wHϳ�LDG;P�f������zQ�
±���!J�"�b���8N۷L.�wa֎�v�hzC���ƮDl��:���u ��pD��	ܸ8De7��w]�����^�{#�y�m��b�d܁y�d�]̦ӫ>b���$;�sOa��h���ݘǃ���znr�Lk�m�]����v�i����mr�"�E0q�=���(؉9{[�C�uɻv��l��n,aMأ^Ӯ�{;cw'q�Q����n<�K��Mf����9��w�ݘ#����n�j�!�6z���:2m�����v�=�:۶�v�mκj�m�C�q��z`�ژ�t�i� Ҧ��Np��%�v���U����l#��"���Mq����1�!�;#\:��d<��ck�tM�r;On�;=`�,��Uɨ�ԋ�h��H]����r�8!Ľ�t�8"Ls�Ƿξ��L�D�x��;KWs[��n{r�ױv�a��!�d�۪����;\�wf�l����;�T�b��7���׵���� �H��m����i
C<u� ���M�o9�X��n�Ydp�9l���3���U��w�3]["�q]���2=��'�=&٫��`���=�\:��n�
�p]�=��ދ�S,��W�X�L�f�� ��u�H����e��Ȉ�l�Q�������{���~]��Uy�22g��A �ۆ߂�s�<'�{['�vQ���	ZWD��=�	$��ՙz�[�2�r�������y�G�P���[}�Z��a]������l���56m�X�5͊��H�����\�}���',^U�7�����T'����O-�^9u~&ɽ˯۽�f�w_6�'w=�?�c6�*&��-�g^ׁ�����y��{�ޭ�1�p�DU3ɈH�]UKoUnX�뾶�����b�� ��^k�Z�$�X�iU�~���oNu�y���䐯�ʾ��o������v�r�����הMn^_OwĊ<���)#-��ֽ��ci�>^j���}@�l���d�i?�v{���A�=g��siU|iR�e1׹ޭ��1/��]O?2I'�ܯ H'����ΔH��� K=+�Wj��c�?q��������*�aL�lA?����>��57�ت�k�?�ߣ� �Y���&+�!�X'���щ�ֲ��� ��o�Z�C}�甩��
7�w[�f2H"u��k�}f=w1��ךZ���)��Q2S_=r�y���:��uU3�	���$����$�"$|fx���a�l���YX�
��  ���`�OG;���fn,�{��޺
��h��	�|ۿ<��'�lZ��yv
zk=����W�h-���#Lw\й%��U�ˮذz��*O�UU~���߷i4��o�so/+)U*��Zj���2�[�@C�NIP�>q���+}���|��V�V�(�Z�
5".�_*�WVS�� �{����1[��Ovi]1 ��By���(W��\�	�j�U>�8�b�Ov}�J��V������]�Q��k�nb���l���~���w����� Wj���Nz�$�u�$���٨6J�[����'c��5�g%aU���}n{��;ULcީ�&����K�����H���$e�3���o_��b�ʣd��毷������u���}�w25�v���9��� �Z�Y��ER6.��~�;����u^.��>�a�'Oo�#�緼4׼�yv�{ڷ�;ʆ�VM���J�JS��R�*9�Z���R����x+����A�����ޞ1��9I��}�bUc�ݽ�|�X�'����5T�+���Il��^�?7T��6+^J��O/s֌� ����	�:Okd�s�ت�}�&6.����km\�0�l���'g�=tKpg�^6��إq��\[o}h<�B[Y�;�NlP���N�� >��^����zT����*��Y�n��×xB��o<,�j�ScO�_tm�o�6Hqخ������&1�j�~��/(�m1�sz֟ AΜ�� l�kh֞���d�%�H!ޜ�KI�9��=�H�c�F�M>�糝�3S.�meߐ{��, l���̘��o6^_*���|�C:sm!���j�U%b�J�L�0��,��l��ӻ��x�Mǭ =�6� �N��������^{�v�p�ģMR���{z��!���;��J�eY�z�H<����f>���Ă<����k�%�ɼއ���5�l�ELrq�^xv�:���������^����c���Pll�ݵi܅����]��㮱뫥�)ƻh$8�2\x�� eZ���:�c��۩{;n���Ѱ�vӊ,�C�`\��7�[���7	���;Ax�r�d^��M��=������z[���)��z8쐸T�92cÍ`ݎ:�v	��ʀ�/2�s6t�u����sNmry���)庞C��]t��&��Ps����W]T�-�ܟ��w3σ�7���I$�S�zID�)�b4z�x�Ϫ�o��g�1 w��1*D���H!-�����l�O;V�TV�UA<��4�H ��ɟ �[����h �ڽ�a����\ϰ>��w���evJa��o��@y��6�6_]�l���}7p�x������﹙�oo��d���cf5��|��{���k���э�?Q$��=�%h�j�sF�- *oϷw}m�����]9����*���>k�$&��o$&:lVz�0��|��I'�=��I&�w4!F6�rN_��]2�l���w�[�n�6W���^9�������rY
�_�QGz���rE#-`����1�씖v�x1/�@$�f��HPMd%~�w��s�緶���v�j���Kr59����R�U�e������]/�׵�]���ˡ�����v|�
佫����L�4���)v۵,�t��W7K̮]������E�Ͼ����$�}߷�BM����5�)��B�<޳kA�#P�L���5�ݝ٘�H$/;|�K��I����mʔ�/�D��ݹ��D����5��.��),�IMw|=�7�ﵯP>'��&�$�hd�4����o�#�3�l"L�{ ���3���� ��Bg7�KJjm�dS'�׽6��]��$����	y7�4P	/�D�`Z������7�B����Bo�%L7Gs����u��ݯE���,q1GcB���V���Ѽ+�y��!$�Qo��$���n�Wʚ�߇��L�33�I|�{���+��T(]��B��ҽSvK;ڷ�f�	vwG!4I�M��d�$tM��E��e������u!A�YF��[d��.o]�� �̢��>����V��%�@�3&�����GOs���7«"�N�V��<m�3��o��&�"��z��C|�������6�X�4[�(�ܒ{�I$����@G�o23L|�Rd%��Ӿ�w&�������D��~�$�Y?Q,$��ݹ��Vw�4K�ВB�9���垳XE-��SS|̠;�{�����a�K�P7���I|��m�h��ݭ��v��d˻�y�5d�o�
�ѥ��ܻm�AB܌�iNM�-�ۖ�N�H��|��hZ��H�Eo �[�a"f�l;TH�����V�Zq��C\���R=�y�C�;1X�_�%3w���d�t���n�D��I��x���I�OoN���	nnp�yv���\�N�����uUB�U]�(Xm+���d��g<ĉ?��Hn��[D��G���V���٘F�zYF�XUwWV�&{_8p�*3�@Ꮮ �w{� KW.����?:�X9em($��u:�P�jb���|��͕t�<���0�¹v��W,{��`]@Z�W2�9�^ɮ`iUOkl�33�\����3f�0����HI S�����}�}�����D���vf�H9���5��X��U�m6�T�k>"�UmH�[��.�9����!�G*�Q?�m�������U-��V�)L���Y�9�$I/���ĵ�+D৊���[�IM���}Z8/TW�v�o�>����p��ދ"�ô�(N���$H ���E>���r)�Z�����q��@�%��V�Z����K�G�m$�L�.�;.�vN}S��f��xI$2=m��"�9]Uk��e�p��" 9�<�П�4MN~I�H����%�fC�y۶�}��f�:�'��[e�&ع��?I���ք�Y5�i�o� jt��d��G�To� `�ܱLM���_7��U1=�\��s�Bv�������Z �"i�k1�{��ڬ��Wi�2�v9,=����]ѡ`1��^7:�7[].v��oi�����U�vݢ5�$!i9��v��l�v�T��=ev��-��^�q��\La�u��ma�`x;m.޻N����̶�X�T=bM����6��Ƭ��a�k�]])9}vѶ6�L�Oj����{�ѹ|�.���=$�0cW[���x�Ȝv�|tn8��֗.��牜�t�L�{0�����ݰ�����d#p��cU�v�ɉ۱ظ�2/c�
G~{߅�9��d$�;���;��ka$�5=9?�4I$��Gn���WL�X�(~����	$�0zst��}2�	8�%�Ɉ=Ns� �n��w�^��1�oأ�	$�I�g<d�$�iQ����VG<z�Xʵ������Z�bv��bF?w3� ���$/9����1k�I?9�h�D�oƷ��ճؠ�TJf#��okS�z�-]�m��i��$�~��Q�%$������
W(���:?n�;�$������ڊ�J誫M��ά�Y����J�D�G�������S[�D���6-f�sy�_z�$�]{�/���m�r�k����&�S����۷\{F�olˉ�'�j�b	"�������ݞ6��l$Ig/cv�I!7��0%�=�VՓ�+91�,$�����i}~� ]d�9	-�|k�����7C9��R�F��zB�����j�*�W��tC3������*ʿf� �V<�[U݀�EI�R8U��H՜W�7fw���NsQ�	9yI�N���I;�{�J$�O���~W�M`~Oԏ#�r��e���j7�s|��}�y��� G��Z�%w��I&x���A�N��I>&gP�"0Y��U�X��Kn����P( $;���>��6��Xގ"-��+�쭸_��n��� �%��SXk���'ĒX�i�=��|bR��e�;tI$�N���$��Ϳ�'*^S�qU}Y��ꩡ�q:ڍZ5ma���x�f��Uī�5��W,���2�|�u�X��o8%z�[��;3y�$% �����gM�u��r¨���i-���H���4���j�]Gw3�����Xzo=$��=P$�[ټ�$�H|��m��~���u�k�}��Ho��.~]��9Z�L���bIc����$�%W�}+�/���S��X�f�+r�%���G�����o)���kwC�D	4�ɵ��@�l^���P���L���������Ζ� ��.�;/mf����R��3P��#*�b���z'�U0����ѥ
����A=.�p]m��&�Lɝuwy�Pƕ[Ά��%�J�t���,�wS�}��޽���w���J���p��w�U����Ө��lw��Wd�7� ]�{��#�ΥB�C����9V*ko��Y׉Z������(f7mHˢ������"Y���_Vw�VF��-\՚����1��ٕ�Ǿ��Ӭk{��[�����&m\XB�j�x�gu�Mb���u-�1�#�vPy�f{�9�Ts5��qc�����B�S7�
ΝY�7�����f�+f*���&��\��U�j�Yۼv��A[�GmmCt�e���Տ�����-*��v��Wۅl�2�Lq�f=#9P0��lQ}��
�yr39�JJ�W+�Wg]�3z���
P�Lmu��u�ۏv;=8)^\�Z>e��{�Z�������w�*�-��mR�4/�1�i�5��-��-t7֕՚
[j�NK�<rv����n�"��D�4�^�Ԇ*j����R�E�3�w>�ɻ���x{�����Bݹ�Rswp[�B4����Ŏ�
�����͍S�:�Uw2-��4Y�{�i��ϜOCc�I�w|����/�]�L�x'gu�S�6�$v��U���G�&tȇ9xI �ʃ�*�j�4ML	Xf�m��������%��e�K=���㰦j-�%�D!!Gq҇Gcd��Â�����yݧ�q�AI��p��k���,��E-�9C��Y�s�kY�Yg�\�=����9�$���9��$�N�����ۭVZ\�t�l�v�ynO72ݙ$cjJ�S,S5ge��(�.s���+u搊�kۡ��:�0���C���P�6�9�mγ�&��+�:sf�O.˅�s���96�v�ٴ�:�"fⳖ�Y���<�8�k9s����痬ˈ��wYEd�	hy^���֓��� #O=\I-��o$�5��)j�a�Õ�o8���wYH�$�2>K� A��o7��0�s.|���'4��N�{F��nQ-mR"���кϭ=��� ��+����������I�3���AtO�W�rs}5�}�O�堙!e��dli��b뭫Z�չg�v���݃�%c��-��;�~��ҙ�V�/w9��D����I$C�<t�[�^��]S����$�K圵�-!�S�"��
���;̭�l���pç��.Ǎ�I��+[�H�B�xA�%eGt6n��c��=�I
��n-��,�b9�ٙA �ŕ��$�Ҙ��&��3� F�wy�`�f�>��O����FITְ׻��������s��ԐI����	$�η�$�'��ޒ���ն��@��Tj���VnT�+��k~A���[�O�4��*����wu.G.�Q۴6k�-&ʕ.�
w��ߠ�r�9��$��Y��7b��U*���.L��1e;gy��v'*�ٹtI��M�$�O��lZ)$����׳6�����TO���.źI���!t�Z-�����:0�q�N�Lm���eP��|]*L�/�O�]�?	�'=L$L��o J�'e�u^ui���J�����fP�T�썒�Qx[�<���Bh��I�SX�躰�MQ>��X�Ot�H&z���(�K;�]�v=��F|V�B�=x/M�PH%�;�bA%�Nyo����\�I�̣ ���}�����gKm�V�W�z�o/#�w=�g�$�-���K{7�ϒA$Ÿ�x�V߆�读Ϳ���A\�~^�O�%S5��w�$ '��'X}a{+�kl�}�R��a$K&of`I|�S�v�v�K=�~mS�\^���wʊ�	���N����]�g:����35oB��3~W�ԩw��)��X+4�n4��z-W�����"=T⃑���+7g���r��m�v0��T�NJ�]F���=�F����cs�7.9�Ɉ9s��hz���*vZ��K�PT�{[+h�6���.�7��R�9��;��.\�{��P����x��)<�q�\�2���.���r������r[F�z�[n=`0����Y ,"]���q�2�amfF^+��'VF�z��;�q�}��P:-ݽ�1�&e�϶���+�n�����Ⱥ�I����;��ϖQ ���ǰs+q�Kr�f�/�a7�>[��)%����`,�O���dp�L�{f��A=g�Kt�Z����kv{� ���6������e��՘�϶Ũ�Q2_����k�߷�h���ڥ����iz��˗��H$���a$��s]����7����
��^���{����u=(�-�s��Mk���I$��N9UF���,��Iޙ�^��ٝP;-�����f}C�>����W�{��a<왘�H�-�;E��N:&{]	霽+�c�
�R�a�^f�ڎ�gϬ��l�ݚɟs�M�Vku��"������DIT޼��;��a�$��Qa$��GL%�U��Ʃ�g%k�����^���\�Y��:�-&�yI�a-��N�];���Vl�#ը�o����d�p�}�d�U����,h����bK�^s���k<���b��G+;��G�����pPʸ���|�I|���4�H.��n�&o9��a'溇��G> س�[e�So�K�SW��h$�Ӛ�;�;ֻ#2�ou ~W��d${���52���n����uEr����EMyz� �S�ɢ@3mGn���'�=�9x�Y�wg̛����d�}�+��֪;+6�&�=�;I�7�Rt%��Q�%�����*1{�{3a{3���w�����n
�K%�%#���r˅�u�i�i3�i�$��kj>n�j,����0���f�ߎ�|ݒI��⣧�� �o�$)�KU�aM#�l�� ��cbՑ� ��_%AUX�y��������>�^���N�t��_$J�%{4�C�wo{_ ��=�N{:��z�H��KU.Lt�1,�@��{1����ȵ&M׻���K�0c�%`�ّfWm.��+��)��>V�n<�w)m
�����ܜI*��ÃK�j��!�[%=��Dl����C��M��I���h���vwfg�'����UW�6|�y�TK�{d1 �K�o7h$�_wN��	$����n{����^�OQ�"�̡����%��+Ǯ�o1ė�8��Z輫{)P�A0��S�D�&o7�$�	��ם�]�%AH0�珞�$\Mn���'n�r|��ٹ�`�m�6pe�n��}m��TQݭ��^��Gb�t{�Ѿ?��I.�y��	���t�:/�.�����R/���^���O��P��9-j�g�4k��P@��ܕ����,p;%%:o7�$�N/k�ZG6
�����0��~�i��NXI*����ϪH�yXtI'� ����ۜ�������	�]�T9���
;$�R��~�w��Mq�-w�!�7��6q"PW��I|_({����x:Ϋ{Y��<y�z8w&�}pN��5��־N� ��/��j�vɓGe�D�s�jAt���/T'����ū{�W�9�δ-��{�MM�$|�������~��㙙A ���,ֹ��ޔ;'9gĚ��� ��W;�N�(�9ޱЃ	��b���A����.����v��:��Ͷ�h�Tu��
@�1+A;Y���tP�2XӒ�y����3���U I(��������Nsu��$���^��mE|��]E��`u�}Ś$j���{^�c�'s=�Wݏ1 �	=+��$�h����?��C1W��{���Kf�&)K�%Ɉ�k_@HK5?R�$���˻egN��݋Mm��� ��f*1|���B	�qN�I,�a��=�Һ����y��� g�N��I$J�餾I�ݙj��=�{���$/�Ga�컫�B�˻��q���\f�d�go��^�*"y��zLuz:%�����h������}3{֡�z�[�nh�<�/j�l��G���.ۻ���`.��^]�RZ8����q���m�Op�=rjL�+��no������}�ձ�2Gj�)�I뵊���������UPa�<tBk�#����w	ɻ�'��? �{\v��l�-s6�m�p�m<=nF�FyKq	#�+���B�m�7b��f01�qҵ�^��+���8^.ʇ.�:�;�y8�vs���-ێ]��VE��� �m���VピJ�۹�9�Mb�m�m8��tX㲻�rH�s��m�r��t;��
#����]��nM7�����9^�b8R�*֔%_�����_�B���Ν��A{��I�ݳ�3vFO?j�P1��ݜ�s�1 {��3�kJ��di�_�U�oo��L[���m���Y���I}D��q�d�'ݾ�r�?|���&v$��z�7��\Q^�|Z2��Q�tw��_�t��%�I"n:"
�75�4�w��1Q������Kf��H(K���l�+��Gw�]�Lw����ۧ��Mjv�����%�\��t�|h��w�ͽ#)�̠�k[S�D�\����ВM�W����;޺Y�$�՘����� /}[��)	31��>���UV4H�9Z���6wE̽���&�!.
�T��Q[���T��ʋ����f�d��t�y���H=��D�*����|�-m�E|��{3H8����!,jf�L�P���qNڽa���jֱ�^K;n��T�s�oVu.{|\�¦����-�~�����9�����|w�������1��v��=O`�����K���$���h�RG�[���^e�3���M�-h�@�9�gƽ�s{[�5۬��NGoŕwz�Y�6r�D�O{{�B[�q��j+�ϋFX�J<ă�;Ų�뛃�Q'D��G�b%��w�tI$o�jǒ��d��b��A�$�lٽ��٣�$��	r>[ۮg���즑��Z>�D����!&��^�c$W�%9co�h�Vs|�˶Nj2�����v�c���'n��^뱷�\�؀�g s�8��x����#-w�{�7���ă=�]b���d��[�7m����ID�C�؝up�70 F�9G?�^3U�%g#�϶<���J��#� �I|���Ii%9clZ$�vwK۹��~�d�q�������wHSi�x�'����$�(;���ɫ�v��n���-� 6a��1�r��5���K�͇���l�lY�A"*'��^�\6�I�i��Cζ�v���2�𽋕օ^/ar�s9$A=�spg���y�����~��9��]�Lj��.�&|��V�INX�D�[��3M7�WW����zV4X�B�O��J�(ݒ��w��� ��.�y��Xo=Cd�j�W�K���M$�b�شW�!�;�1&x����d�WDt%H���;4�i؋���H�`Wv7t�Rc�gu�y5���_ql|�d�B_�.瑽j{3�����I$�gvf|�;OǱ��3��ӹ�@#�7���k��0#�4�����!1O
�{}/�K���JK�Ս�,$�gvf$N��z��m#�밓i��%".V��>� >���$@$bv3g����}H�Ǳ��%�;�ϒN2}���⒫6�6�Jo#)��=bq��	Q��[	/�U]��I>�I$�W��w�t�ǱC�1����m�����~ʽ�
�F�osq��n�2����mr�zx|�q��0=�e����#>5�a��Q%q܎�=g5PU�W��\��ϑ$�W��f�9�Z�({�c�O�L��l�I|�}Z����r�xz�}"�����r[gn���V�O�8h�{0�Ț���uǱGV���j
&R�~A׭�>� �l�l�K���N��v�+Jn7��|���om��`���"��B\������z%������%%�5�����o�ܢI$�+��	)=�:I�=�:�"��,z�$����tW�}%B~ �~5�b��<>�xp�<s����RN���K"����'���XD�U�
ݴ�zM��;,�"o����ݭ�@�ms�I$�Q���� h�f�o`o�ߖ /�	]�H��� |5F��,�2Z^Un ��=$$�"q^���I ��c`y1p�1��k&S�i3���
�C�4d����p��Y��碖@�y[tkb��Թ�jV���N�*�̕�}3�ŨP����mLά9w=��7)�W���:s|��7�)ekȫR[L'%�F��U�%�Bɝ{V�p 
7�0[W�SXa0bUy��Nәy���)}3�B�m�.�6������wu��!��]r���r����c�n�ߕ^rRU�̫��������z���n�p9W��T�B*�N��_rY��^�����9|��x���SK�Ôh���Sn���';[�^�ي��l���ר^�'�Z�ǶGf崥o�S��r�tL�j�K��p���n�O+,ze�	�P�c�|R�)�w#�2蕠�	�8��x�$�Cn��p�Y�Y��u�W����(����|s/���4*BU��)�vJ�=���X������%=��ƪ�
���:�n݌93�6���Wg����2�L��@�sSp=�r�)߈̯矅�M�ڻ��w�we��D�m�L^f{m�a�2�\��S�x/�QA�,�2�3��Pq=y{h����H��}���F���s+.a�ن�Q�Hg5v6���I%B�+:�-�#P�k6l��
��O!E�G�.́��Y����؍�7+�F���_Z_�n����Vv��F���}��.\�WNn�����ƻ�ݵk��Z���V�Vie
��)��h锇c7Jե}���Q��=�t���&����c�S+i�qfp7À���,+(u:2�2�7���5��25ؚasn�[XvX�#�4�Lb��iY��V[b�г[f�����,�㭦��5��f�,"*ʙ�ô�vէ۰��+b�mm��m�Zٵ��[`�D[6w6��e۝�ىm�[%[���Y��gMֳ�����ΖX�3��2-�shζj-��9E����f�+mc&цܷQ��6�Y�Yٶɱ�gqۤP�KDݳv�����lu�l�v���-��:����2�m��v[(m�Y3q�a�t]��������6k8�m�w-�,���&Ӷɶth�� L�2:v�jX�6�,N�d�m���6֙�N!fA��[�,�m��xÏ�g�:8�P��'ղ'�5�'�o[����ֈ=�cm�Eo.�q\�q�����-�iI�|�+�Ux:�nv����b�Ķ����0�|��<A����ˮ�ն�K��Gn�mO�/]�7F��.9��<�7�x�*V��2d�OJ�v�^�7mͮ\��TWGn��F�=�ۗm�5�L]�X(F²�DՅ��#L"G��b�3n�X@��˹�T���3m<�q�ڸ�Ɨ;ni�ގr������u��3=%���rm�l["���͗��=^s& ����c��h��$	!���ZAod;$�N�H:ݻ��G;p��0r<���v��n\��l� V�>��IӺ��v��p��l���J��yG�6���ۘ5��+�ڽ��c��lun�s�l;�n!�nk���u���:]��OX.cۛ�n���j�|n��/T��ـ{IGsr�܋�k��ގ�����p�uk�=��uۑ�c!ϝ�n�D�S�A���n{m$�v��[I웩��l����l[Ș���1lv��W5r�M���dۘm�L���U뎮0:1��cv��.��l����'O��󵽵�;�ᚺ�5�z�ͻRs-Ш�����>�EbӺ&ۋ[��;c�=�h�;��]<tM�^���˜k�˾ϗsj�I�Z���
���g��7	ѣ&z���c�/\q���e�;{�,v�6���Qۆ���=���\E�N���ؕ���n:ۖ�� �G9&���n�0sG���5�0=��Ԭ�Sv�s�w]��&}��"�]7*���n7<�t������[���s�������+�.G��ܷGe�O=��X�nۇ�w�ㅆ|l��݌��n9��*mX{dͮr6���8v�͠嶮�xB�J.T��	��d�d�\�G&ӎ��\ąӊ�,��m=i�0�0��:�lvd��;�S3���������m�Mq�:�ե5������{q\���=6㎽���k�դ"�5�"�8�u۴�q�&��k��Dn�ŕ�twq�;��n�&ֺ{>�pvݱϗ����x:�)ᣎ�c���cq�N�l��N��х����FVE�]h��7k��i��/m�痶��; �Y�s����%x�v.[��[�=�Bn^�vΰ���wn�9�q�/I�Ϣ�y6�;urq��9�Ng�|=��7n�{����qv�9��7X��V*ޑH;&��9N�AN����5���EږM�X��y��}�O��b_����=��7�� �wYF�>��G��Bҗ�]��'��o~$�W7XM�_�>����v<σ�[�f��{�/z�Y�9���~$�4�V�I���6�&�]�~x��}/���>�UT)U���sF��� ���f��H=�o�y�!kJ$Fi^o4I���7�$V|����v2��L�v�B9��>#w�y���t{�����O6��͑��E��֗���V
(���A[����ߐI|����b~��=ӈGI����,�
�6<��$�ݙ�/zl֎k���l:Т'�Y$�5Qdk�����;Z��Y�R�2})��*������ld����ә�� �y�[�ϐ�N��$�땯kN&=Y���E�ZuF�5*���WD/>9yLr^�j� {g����^����7�������x*v,[�բg��V�9�F�)�.���b��gв����qP�qqzsxg/a$�~��2I&��ޒ~'�+�u�����wAyZ��Ԋ�����;�>~% �t�y�$�;+i_z�찲�y뚠I|�Xg���ISgvf|��h�Y�/ЗS9�N����x��H6^c� ��%$����I�խ}��^sX�W����hUi�Ԫ�)^:+ݾ��?h��~N�����5��EH1Q::E�2N���J�M&����9��}��F튱G+MYk�R|���:�i�)��k+���92�	ϡkV:KU�[8����B�oo��~I ���x1J�'�Z`�>�ΆVR_	�n� ���I>&to�H���J讱㙑�{O{���]Qݚ��K������	 �"��h�Uf¸AW�������s_xQ�_�^Rg����'�@�W+�_�V{�d�>����[M�����ON�wGh�$80#��x��[���Z�������T�k�{2
[�I�]��hǻ�N����Nn�$L��oI������6�TtT�ǘz�g�ny���wt�w�I%]��>�K�u{]0���jyŹ~���ױN�Q5���6BFK��R�\Tl?kx�^�T�E�c6�I�;33�G9{|�ߵ�f�zt�[�Ǉ910�Q)
i��!f��Nn�Fm��S�N2�s\���6T�[^|�*�P��]�������⼬:$�j(��yy���]['~�n�@!"x�N��\n�VY42�ˡ�^=#��n�>��>�9�~ǃ($�m�v� �<�h�;՗_�t��� ����H1��+�^�ֹ 5E��D�����r��as�}D�~��g�`ߵ�ϴ[�^dNr�[�c��dm�Ur䜙�~;	4L�ާi$�CT�;%����ن�hL�ك���r��9KmT��40xwc$��kw��6�^Q�H�V�gT���-��c{��\�5�l�^��<E�|�G����C���&�Tt��׬�o��~%��y�����~s"K;��$�Ӹݒҝ���Us-�:���9q��gt[R�Ї�����g���i��.����d�x�Rl"^���ɒ���|�kS����"a�m�$�IM���K^�[�����v��o����ϴ}�;J�#���+ӽ'К$���0�]��ȍ��H�ߚK��{{3I/s�9Wg��4�U6��E����w�k ���y�"RNi8��d�~�\��
[�rK��N���HM���	,��+\q��\z�&�w�2�絤��	���K��ٻٙ�H$���k�3|�3	���`|��qy������l��l��@����?t�2߷�����=��Ě$�o��O�$�9_7�Y�7�s1j�;�x��̋w<�X�4K�YJG��12��� }����<����n\DCװn�˨/q7���:�\5N�gY���ۗ&���uee��z�ںQ5���\�Ț��n����<e�r/d�'D�����'�����LOJ��W��\�h�v�(����r�D�/n��˓\7<�k��,��yz݃��㖷:��c;�3��u�,7��Y��V�E��la�{vn���λ���m�p�q���_-��q�^�{s�k��[��� ����ݳ�6oK�0<X-�Cp^(�z�۞���`>.W�ǬJ=�����Ka��k�-��?{��,Ê�(�Hv��E�$���s���Hg+\�b��~zw�8��6($�M��ė��19#RK�K�\����NH��{~����a����������w2�#�U�8i�N�|j->v�DFFZ���f�2I/���Z%%ʂ��wY�`L]��$���6�D�?�����L;V�i���;̨�5��w�@]{��I$ε�n�$��cc�/L����������v�VWH�+������:$��c5�;,{�e�0�qOI*�$��⹼ �I��o�@�/{����FڌL��E��I>V>�-:���8ǭ����S�vGC������ߊ�oi�Z��BI?4�'��I�Ѭd�qN�d�������@!"q^O�;��xa7Y�fc0&Oڱ�>]��<<�静�+U��C2�C xśwo��/.U�z�cqr�.���e��\i���}�-�Br�0�;F�2^�+��U��ʾ[fiG,�t���
(t�ُ�$D��k����O�F� �>�zy�+�34^s��V1����[���@ ���3@=e��E�~��w�����s(ρ��y��@�oO��Pp [6�����
c���m�($�Kb��K��Hݴ�I7��<e{����z
�|\33>����U���@���/�ߐ	���}�v��[�n��˖�i$���($������}�A��3F�<�X��
1�nϟ�/̉��6z�r-r��d1��,��$j��%�*���T�db+��|�Mk�>���3� >@}�v�f$ꮦ��i;w�����l
E$���vp:>UIPF��uc�|��Lg�~��7;RO_)Ud�$����2�����>Y���.nq�z�����z�z�1,�A�w��{��#kyw^x���^�"Z���I�ں�}y:t{�U�]PY�b�� ���OWJj�����]�;��U��Y�;�O������'X���\D�H�������{����I~e�1"��t����"I:<��I$����G�}+]"�VƮk�&�A$=�ly �z��
�]ɟ����� �2y:��%w��/�<R׌����"@��2wC�{��j��ۯ���6!�w��ջ.���s<\��fbKf��g��γj+u������AU޼}�s4 ];��"PIlw�0�ŝbx[�j���7��Y�ݘN}���eQAVh�b=��̃}]�ޏ�ҫ%�� �M��%��=Q�H�����c�yPm]/�(����Ϗg���-�9̝O�&�"��v��>�W���I����� ���2w1@���Z:�N�Gko�k���LW���.�4M�\�IH$�Gz�I�����}�@ѡ�֢�XB��S۾g1�Tt	�]yIz��R{SLt;b�s�懃ǡc����Ox�Z�=�.�b%��`��5�'fg�"�.�MR!U_Ʈ�0�h��		��ݎ��ߝH񬝪�I}�����M��ݐh�jyF�o G��������8�mTl��>W���63��=^�.�v� �=���we�q���}}���2)��Q{=����~Nɪ$
�Q&M^���z�ȱ�oBH�Y�\ؤ�x��j�&�R�m��=�0��#�����wM����71$�H�i��A�ck2s������w��	���d��^�K~�I�Tm�I9�H�0�Q�-�I$�L�o�E ��c�`�~�ҡF��ua��3�0�n�ی9��~��K��; �H��O�@5��zM7�ɬ��|���d'��'���v�:�ϛA$�N�y���W/]k���ܠ%}��b@$ ��o4� ;����ɴ���
��V�؇2ǳy%}0�y��wzا[�pe��~]���T/�om��6�w%�wgu��'kF��^�뮴h]׬M}K3rf���F�5@���^WX�K�rvi:y,�i'�/���B8��h5�[��yqt[��t]�� \p�s�S痙8#66��88���t�v�SN�lk���G�¯ �+����I<9,i�l�l�碚|�{)����ۮ�NMnJ�zg�Qتz��\����cX�Y���Ϗ�I��9׌'�Ywen��s�
cm�4�g@Y��2:�v�귄���Ν��S�s����z��8�l���z(;a"����e%�2�����ِ_����	 ���ل�]�gl�����iuY�]��ɡ`k>̣�,]��1�^~�c�o`N�*y
��/cv�:�(���KI}7��	$f��D��+��gW#�B�u��Z���f Oo��!?Ix�J���#�s��@{�D�&�vf��:��EREVml'���ZLv�]R�I!�#6�I.���ĒH,��oL�sy�۲��i�{;�4�a6�*4�Q�]Xmnt�+�O�I�f��ɣ�o[���I8F|���İ���٘�I,��d�����x�σ�q�B �*Q4�u�TEI�<h��v���[Fw;U�&TT(�Y��$�uZ���׿|Mr�t�$�L����MQ ��d��K��B���D����$���B�Ze��s]���;�}�;v{;s�]]��iV�R�0�6��s��a駳O��t���ԝx�Ǳ꼺�Y=���J�ub�m����<]�]瞶=�9�I!;��1"R�ܶ�(%7d\6g�ݺ�����J��r2�r`O��3�I$�we��JK�mNǖd���|I�Oo{�O�4I3�c]��(Z�5d߮��%E7�ow�I%���BI$��  *y�oVy�2�tI��w{ois��b 1��+�g�ۙ�v����w=�pA�ΔI�M��|�)gn[i>I!���WD쏟�j� >����/6:In�z�ϔ6g^���͢�a7���Z�mF�o����'ޮ��h�R�y��'П�on&I$BzF�� ǯ���s�31$���~%����l]�WF��o��cm � U���V_vc������y�	���3��=�)��{YԀO)�n�B֙nLSۖ�i$���%%ݤ��k����o�����P��AQ��Ux[�pznu�e�C�����R��G�T�;P\5���9�t���zL�����dv�sfoX�gc�.�vO���\�;�ތ���+�SYx������%_�2�E�y܈�5�ַ�oŦ^� t������5m��(}���oq�h)b��%���qNMg9!Ѻp��Ԭ"�gW��\���� ��n��.�v����Ԙ���U�Ŏ�a��4s��y�2>nb�S. U��D�Θr%�hWV\�������޵��M��2D}�������w�uv��IVr���L�s��B�E����&܄�X��V��j�9���ԼQ�w�ʾ)9�²M�z�I��^��3眺jai���$����o�oƽ찶��0��ԭ�$f:��r�e�႔����8Q���T�Zy���R�X���9H��=�+KTa
�m#˰�kel�7�X�C-���C�ܦǕ�^�uVk�X�V�^�C%�i�z�z����NWvbk���un�	5����S�c0�o�:g.�W-�Ͷ����o{�1�p��λq��C5>�s�!LQY��Y�QW@�v��޳�u��ܮ@�z��n%dg&-�ֻG`�T�p����^e������:'�P���8�6�\��Y�[���Q���m�Qf��ɜ��c	[f�vv�gX�CMMe�QB�=�#}����)�;M�ɑZ��z:K��˩z*�c0������dI���Q�����;�Z���O���h�H���� �#��X��i��Y���Ve�gfgm�+#l͑���l5f�ۭ�Yp���Z�r;kV�m�m�e�m�l�fV��A��6�#�8�u��i���ҙ�"S�ZpvY��[��2�ٵ�n�����90SV�iY�Y6kfs��h��[l���f�L�q�-l���\m�[�2�m٢\l�ka�;2FY�����0�m�e��n��L�0��7m���kN�ѷe�q��[[2ɳKq��cd��c "�Z���Ĕ�ȃe�,t"�j��m	�۳�d5�q����[Gh�M��M���+,m����Jpqs��H(NY��!!��gee�l�Z�m�7B�K&�%���;m���:I!6ݦ�M�����ێِ&KV��ݚA�JkE���k@��f�kMbe��PIkZ4�q�6�m%�6���XF՛!�7�Mw�H�y��T۰-�{�X	��eDN9k�����U-���۩��PY_%������$�2f?0�IN����v��^y$Lv����Y *ȥne�]�3����{�+�rwܕ�	+�~d��Df�����Sw��	{݄-���?G�=�+4hRZ���.�j��s�͝��A�zM�nݖ��)֣;�r;���t���^@؁{���Bv�f`K*��0�B�K�'RHI1����,*B��Xo幝�BI�s;���w��(�Hݱ'D�$����%Q `�������~�Z�V�b�QV	�-�7�l�s���ĒA"�ǩ�^M^f�w�I	�i�.w�����yN�n5b���ܘ^v[�7x��'�A�~��"zwsy�I%�ٵ3�+-Uq�i�f3ԛ@�Wv��\��h�7�:R�S���ŋ�n��`�����f����U/���Pչq���p�Ǆ�%Z�+Q�s��ԫ�՛7�y3TtI��� 1X%�Q�@�ܘk�総` �=9���Y	���I�[��$�����	/�Aw�����\���׫��l���U��ks�����$�S�;������nM�K.������J��"����oس w���l �Hlۍ0��j�V��1��IC;�����9���>�l���쳺� �v�&�"s����$�&�{�$�M;z�/{o�+��S62.�� �8���b�}�)������I n��vI$��>�U�۷�$�ݽ����K�j7I|]n2yZ�*nט��]�9�t��z^����';9�$A$�q�%Lti�癄L������ݙ�!��zBn5j���ܘ�y��Ϡ >?lt���W�����5:w��I$�{v[$��P��Ǖny��w|W���7ſ)��w��ޥM�BF�8#yŮ�Sb�t��Wp��k]�����nm�U�d��7�oL�t֔Q0Lq���on��-��v�/mn�c�ݫ�9�E�k�"�6|ㄗ�l,uZs��ogn�i�;��㵲=�&2#N���IXw��urt��n��-�Ք7���o;[L�e"ѣ9�:Æ'7=��*l�#a3�����ucZ���mAч�����gu��`���GR7[���o`��ۓZ5���FZܨ]v7u������s���g����/]t��Y�!�,H�q�+���'z�<�>��}��F�-ws��{��{���� � �{�˟���j�K%��s����ӥ��%�[�R_X�7F����da�Dٗ��Ey�,�����h�D������$������]2�{����^U��$w��dy�e�8�b=wۙ�}��D�iS9�q?:yW�e�턚).��	0��yfL�T*���9I��z))a�M�RP �x�TI��x�����)����ד��m=�x���G��\πF���Uj���^b��Q3��6r��o�Ҩ�����	$�$l4PI;w�3䛭Z�A�Q{�\�6��	FۖPpP�񓴙F�3�W7L-Ӯ��Z�A�K���}	<5j�����
�6�	$�HM���$�If�����Kl���o��9��n�5D��{��f�z�c�-w&����`��I���<�~x�=aӗ��6�S��"�3���l+|/�F�7!}�n�zߥ׻�ya�n7�4��볗���W/}��$���HL��7(�D׸�hxsě5�����'7�i�HL��izs��4Oow��I &��ud\��������y��_%�7���{��/�4J�th[au�f�J�	��J�ɏ�C;s�$�K�wfg�$��|�z�3d�	>$ѥ;���([M
�D+�Տ~|ـ$L����b��J+��H�����/��vf|�(-;��Z#{�/5���S�hV����Y����8и�պ���s�cM�*(�`�� ���h�#��=	<�R�ʛ��۽��l���o`��;��iw\��=]��=�����S�}����$��B�պ�$W��1hS��A�2�
w#i$�t�oI/�Ÿݢ�[3R��g�릴���J�"� Z�L5�������=�b���%�|{¶���!���a��D�t�0�,��'g3.�$p`�����5��^j�[X��&x��o�{ڪ�\�v�Q�1�z3+���z�$ר��&��ޒ ����i9��@+NJ92���=��;����ۮ�H�nǘ�I$����I$��n�����q_X���RHod���%3�B���E+6*���(۠�@���fR�U��]������{S�f|�	$�>tI-	���,���I�����Gц6ȣ`|[�$Q��g��ƽWG]��=���k>�W�	\����YR���x����Ľ/��4I$�7�4��v�-�L�{6F��I$�/���[�nz:�U��k���Y�AϞ���y;��9�y�|�IJ|�_!;��E�34fu�.�3�H�%%��WV�~jyg:/��!;����/�ypRS_@:�4V����k|�Bƒ
��69�u8�w~����n�9�߀�w��I$d�?0�(>����{2�����F���]=qK��@���r�Q��;6���G7,j�l_�J~�E�F�mBn����+����Ȉ믶�����T���7�Oi3=a�ݵ�j�VvF�I$�w�b����)ә�HWV�O�AC=��"�A��fg�?wVkӛkI���Gg��h�(;�$����֭m���pX"�H�"	V{�P���a]R����o�I$����~_$�H۽�>'r�C��<�*���$xy4�r��x"��%��Xk;�oil>woT=�WY��g�%�$�I��Sx�ϻ� {��nE��=�����<䜮�]w@���\}���J�'ӹ��$�� ����ω$��ɼ�~~��V�0�D]��ʼHFW/oh���o���	�y��4N��7(�D�)�F%Oit(�$Ѱ�7�'$۔@"����t�IP�h��~N�ΎJ��Xo(׺�P��2I&�ozHI�$%�ȋ�����[!�U���-[$�h��2��3W�,N��t�� ��B;�.I�ݲƝ�T�fej�bϭ�2ެ��ٽ����瘀�J�mr��
nT�.��W-%mÞ��J�������p�^���ES<��8��ӫ���w/Y9|��<uR�˘�����Na��շqua2ㇲȁ�r$Hρ� W�H�ȡ�J7`؝؎l'c���y�J���s��[3���[Y�-3@^(��9�-���/3֊ӎޛ\���!jMRui�{v��$�ul����݀:��mOi��ƺ���=M���-6�/;�s�k=__A�����]�����vz� �'��B%k�I�񻭾�!��=�E$�7{3Hw4y+Q��
�#=ə�@H7�����bZ�����ogpl�P��f|�	 �kD��0�,vo���p4=�R����U����������� |Z���o��h$ǽ�!&�4W2w3�͹'���KV��W��f�:붼@�>�9�Ē_$����D5�Q�k�y�p�xej���!(��Nj��X�V��S�\�%���Q�7�wOf[���7����D�IZW�$�o����4HON���w؈L��{F l���+��%1ֳ�g�����ƞ��Ä �QUS~߁���l�e��{�߻�	$���ȇ�'�kܢL�]Dg�o��)3sS���D���?��*/�]�t	����m!ޑ��	h��{b�"k����q\�;ⳬv_�#�j���-}����2
幬f��ȵ^��M��V�˳0`�V��N�*�dj�^�R�4�ga��oВ@Z�ȲMh׹F� H�oG�Ff/lıw%�{��B���})�I$H��0%����:����o�'_/s�lA����y�mA��D/ҭg�=��a���%5%�^�S�I$�Q�I���{�z@/MI�P�h�W�>�LےzP���կ1��s0�t�瘻�L5��;Me�/+q.�V�4�I&�h�@n��f|��K_�.]Y��{L����#��?�cj�k$k ��ǆB^�q�͹�{Z��)H+����2Zʪ�zyrw^��I|���6�I�۹���$��Z1�خ������:�Y�&�(�u� :SL#�����ϰ{�V���[9=�@	$��{���H�۹���$�������\��S^���yHB��j,ˈ-ԙ&��;�}	�@�[�޻`�8�dt/e{9
2��j�+VN�
}� �lMB������ʱ	�{}f�l��=m����o{�G1ȏ�%����a-��oH�\(1f�)
�H[i���������i$�濛 �3������&}N4qolQ"�=M�b�^&��ٻ9�XN����QN:�:C|	jaٱ괇9��	$��3�������b�U�I9yn���-�0v�q+�u�v�[��<�壗��h�*�N�c]F�8���$���R��^��+��`��Z�sg���|�K�*�����ۯİ��7�	� 8
UtUo�j��ՒNǙ�g�GS�W�k��Ic����K���[�K�)�G�H�>�\�y�ߨ���$P�̏��s;���k�=�J )7�kSYg�L�.sy�s�^���K�<)�T�!f�UӶ���{BH$���1$�@{]�D��Hv��W^ҷ��u<hє��0����a+:�A�c��˼�]�ͦM,��E+_'{ح�Ś���r/x�^#�6�;��"��&�{��r��*�)\ǯrk\P�h�����N�F�M�tI���zI� ��뛤PI!��l��`��[�1���~������.�$n���mG\�إf.�={y��7d����~�Zf=���㐿X��Y��J�J�|��I$�r�?�X;�Y�%�iĤ�H�M����w~�9b�`�Y�i5�r@Z����=����7�� ����s��f�9.7�%u����$��J5tUo�)��o�H��cm$ODG?}�ݕ���ۘ�\���x�'ݦ� �vi���r�������$�{��MI5P�&�?zo�&!��k���=� >D�ys ��JgT�*��ث�d��? �	fN�^��a}��âMQ$���A�Oޛ�H�����د	�����I9f��0��١��	Y��ah)�UWD���Gk��>U�^uٙ��s�j��|qL]�	�3�uۻy]��9N�w��c�]i�4E�o��L�x[�r�r=W*��$�;��>jI�&�����i�*n۩�95��������e'Z.pe��;����O+e�P��x�2�����R������S{���uC�G��_Y�M�������NІCU+�fYN͙m�H�Hx`�Ev{p +���z�&7��V��pA�n��1K���ќ&];���¸n���>��^WS�t�Jt&T	�uX��mMm�;wF�ۯ69���6ܿU��H�*�K೮�A���Ȯ� ���l;���]F�&�-Ͷ+@8�'�[����8ϴN�"�FM }��ܲ�F
tV�﯂�kr*u��%���@���ޙ���o_�����{j��-��>���׮�)}k/�T��,pS�n��{�,�U)�IS�Ɛ�?��sI"���e��x��v��݁����fc�YT%�k8U�3�	�e�R�H�vGz\��U�Ӯ-"cG�K�+n�����T��&�*Y��i�Iu��6�u���Rw�#m�.q��ǑWN�5�$��
����a;�[:V�]�gxAZ/E�+M�ݢT���ۭd��i|�e��Gx�Iz<��!��C�1z;s6�D5c��pv������2��X����]B�)� F�_$�/(Z�d��lV�--��7��3&���tBi&��qrm������ݖKm���Kkkwn�Y��27(rk[���3i��m�u��:t����ݸ�C��̥�l��mQÝ�em��igf�38�n���vkk Em�̦F�E)��ݓS7饁�v�"ͥn��wfvZN۳,�Z:3:���v�n�Ζ[m9ä�6�.$�9mX[Y"$�i��mfY����Im��2���I9m�m�k,v�,�;�!K���;7m�Mۖ���d�a���-2gvӚͻU�(L�;L�;	�+l,�6ôt���8�њ1��H�����Ju�m�i����H� �m�̣�gF�	�Y�f��3�� r[ZR�n���\AE�l�pqA'gGrmiGGn�gZH�ëK�>�*�P���(�u���c�tm�A��<P8ԋՇ�v����=����Wv�J�݇f{��V.,��g=��
�ڹ`����9�jC�Þo;ɻ5s���[��kk�Q��C%�f�{C��A��s5��{s���n$x9k�:�]z�����I�;�;-=�k�E;35�>���X����64�Cv��,�m]��0=��[����u��q�0���A���ݳ�ؽ�U�,��ctY���ڜ7�P��uf�0�q���ܦ���v�+�X�n[���5��w���o&Kv	�9K�^���ѷb�;WH�@�K����˄�Yy69�^�7=*��ۋF�0�f�;�25�v����*���S��-rW4�v�X�����b6��pvvR�q���z�.�a�����tZvCPp�k�qv�{BF�l��ݮ��r�&����IN�q��ڌ]��h�#7�َ���]�sg��kI�{L+v}{d�3�t[�:zm�,.7e4v֒J�n��b�zK�vaۃrٵ�cz`N�O�ۊ��3��/Y��8��\.�;\�'�K��(�s��m;���m�ns.@(F�܀2=�������c˶8�9z���^LW �1��ɑn�m	�74W^�q��;�v�p�n;�	�E��)rk�<ݷ�\�n���R�v_nQƍ��|�a���tD��Mi�=��N�9G7n71Gm��UPX�ck��/{<��1�;xMb�cFvݣ��23�O�8��=[�W���\�G�<�����S4���ۣ������k��H��g�t�wny�b.���׈�7a-��ԤG�Lc֣v��&�[/�-�xX�v�����\�3n�u��y_h^q;��+��z�.G:�v�-F8�_ c��n6�u��ü�X9�/h:xc�����(W��W��u�6����,�.U1]C��	���i��\�W��n�T�#q�b�w=۶�Z-ˎ�=�p��r<�ks+D��<�k��+8�ZplӍNDNu֊�8{vv'����;c�GX��;��1%�M�m�3@O�Q�mۆE�svݞ�n��l���غ�@-�ᱭ�oe�Bo;P�����1�އ&����[��lW6��n��F�l�� ���{^Mƶ�G=�T���i���mg��Avnz�5D�w4�����t����&��<�.9���g�ͺݹV8:� ��q�Ϯ��s�yݶ͵��v3�nzz�,\S�&��X����:�q�)]׾���.`6ߟ5��4I��}� ����ðz���� m�[��ot?���c�u�s��U6�!���A$_E��m$��٘&`���)~�;+.pI|��zR�+Zj׍���>��{��{�T����aw�� G_�y�Ϸސ
�P�D^X7YW�o�.�j�2�_i�ʓQ$�^�~%�{7�0$�9��6��xޢ���@"?sy�AF�4���H��2b9�w��� �w�~%:�{tW/yt����&�_\��s�@%wLl���{`���ٍ�x���6rd8�z��m;K�mŞ�X�s�o9��l��huu{�R�ϭR��|�34|�w� BJD��[��������͏"�I���'�\)�f�I
�����ی�>�3��.�>̜�����mw"��ʻ���;VtFzm���_՛](��[>�օ�_m,��PN�[(KS-th�qf�ś�Ϸ�ߚ �vo�$�I'�;�6H$�gްf����ل�[d���n�I=�{@���g� f��Ht3�\�H�]�;��h������$���W
�	�>
s���y���m���S�Bh�I����I�<=#ad�f)y&yh{}�I�&�P�
�E�u�v��
s��K�J���9nH�Á%Y�ޒ|I$�gs���?��E2��MK�����B�W��r�v����Ӛ�ZG<���@�J:�>�U+�5ѧ�6�"eYl����*I&w�'TI��I��2|s6$1�w��C���BM�x�k���R�ϭR̸�W�sh
��:����&���sI$����_�$���͢�J���){Su��d���S�I�h[i��4Ia!��l��7����ӈ�۳�o=IT�hf7J����qX�4]��<�C���ї\��uO��_
9��,�t������$b���eܦ/�Z�2>I|�Y�M�����,7�נ�8�~��׸aOL$��\D �#��L��&t�̝�����é���Jm��;)HZR�mz�u� o��kd8_j>�&z��H����f@{gvf�w���#W�H��)U�x�x�+���K�f�e�MXX�����E��k�{�2���B�[�)�ؤ�D��m$�Hn���	J�[��_ʳ)�)��f�>���>|��eVa����bPW�Ҵs�>񙖔�'�M~��I��w��h�^��V�6�����!�Q�R�ϭV�V��7���o}�y��$���kd���A�z'�I$���+�����s^.ɺ�QB�Z�	��:�y��(���~I S�{3 H�����S��}\":.{���
�����<�q���������x��-��e�������ݤ�S#�\ �QS������Ϭ۪ȃĚN�o�%��ItH(Q
��Y���̢M���Vz_eJؕ����I�q�$���ل��ͦ������:�˝w��+[7[�l��hbvMT����+�lV4WS��k���Ea[#���9!�ZܶR��H<��@}��s�I ���TM�|$�G;������������$D]4
7tj���槶�E�0�+%{m�G�w��$�ݽ��$�A9�ۤW�Vy28!����({;s�D��)
�	U�gƻ��{Ka�7�٬��}�:ۼ�Eb_�<I����zI�$�`�m�6���!,���lˈ+�9N={�Z��TH˹ʄ� �m2@y�+�V�L�Utx�n����f ��8�1a]�bж��h��?����T��.:�O���$�I&�N�m�I4ty�Ѱrz�Kݘ�G��6���X
S�]���U�k1P��wm�av	���u�Q��ܝ%��'��Fe2�Z�VD��z�'@�p��5�j&�6��U6�q���j�i�8�/J�x�(�[]��*Ca2��7]�n'7a���� <�G\�ZlA�x�½h�@��W�Ƭ��w�dwev� h6.d�{nN�.0t�v�F۷<�QY�K*p�Oa��� �8�K�q,�h��-�oasr�I!v���]lS��v������t���N7���ͺ=�S�����w��qm˚�������m�Z�6�x=u�k1�����	#u���
�����i��W�#��^I�� ��!�����IE��]Q�	3~~۽���q$�n��N�ܐ�l�R�b�o��@G�b�g�%�� ���d��<�cȠ��{G�/���I�e'@ѻ�v2���m2~$���,�J�շ�Z^�́%�I�߉a$��7���O�<� �U�b5��������{�	��h�CW<vKI	�ݘex`�Nwg�ygfM�B��f`n�3�BYb�wV����I�i$�'s�]�2vA%Gy�N� A�'�"	'��I(��;W}�Źɭ���x�r��Tm��/nS�v��n�$�Z�w��ea#-�nF�L�s:yuTX�
�E{�s ��ޮ$�%����	j��cG{�����!'G�Ij��-$5� �D+��mngL�H$1�n�v�D�=g��=(][�1e%��f�I�+.�U�;˰��oj̫[Ʊ�łe�q]�%Um1����cN�]Rn��,v�.?
�y�1�"��I'�q�$�I���I(�L�EϽ�y�׹��\���m�nW�z���~&Ow��$���I���J랷=�$�Zc����L���	x����D���.���w��V���a�t �۬?�Inwvf|��$D��W���V]{gA�=g2�Ti�7�pR	�Xѹ��qH��ͮ�[��<���pj���	!ٽ٘�I!&���殚��k�����u��4��'��mv9U�k��v4`�Ԯvت&�*�c���c
&�^O��X(ڻ5���݌? '�w<�	 ��_�L����:ӻ����E�d����<��$m�A]bB���ϰ��]�+�אޝ���I	�{3K�km���a��S�e��%�?-$5��h�A������ 9��` �L9}
ޭ�������Ͳ��v���������L%/��)��A�%xA��7{I5�v�������ֺ)l2)�q��ܡ�V�[!�\L���]z?rH$�wvf�HI����ܞ���l�r�`+����^���߼x$�O������Ht���#��v����hD���$$�4�a��7�n�U�N������=H���`/�.������ϴ1 ��g30Z�_�l����ۏ����+�.�.<�F�V����v�q��WB#q�"�*�oX��o���&UgO|Wv�O�$�'�|�D +�z�'���7-ě����I���m�=�;s,�e�:Z���1f76��5��צ��g��߱ �Ir�ݰI$;�m��H�ߧ����-��Y����O�Cy��Hڂ�A\�y�\�Z >��30@�44�o�fnj7��y�I|�C9�Z�����y ^��b�K���{e粴qs�X !~�"I$����L�o��#]b׃c�
��<
�`���
���G4���y\j���l���H�~�z�n)��ǵEZ�W�L
�S���7���a��ԌM��!}��+3�ǿsX�S^d�Q�d��_o�T�$�3Ӽ��a���`X�!$�F��Z�I��������ۥ1k�z�͞�+���˘�'�i�'�M;YS�7L,��,Ҵݮ
뫇��-$v;�:��m�]�z� �'z{�B^R�tj�� 5�k�İ(��vA@L��1���*N�8V���`�/D�?I?�G��I$&���	 �MǄ�=E�F��{K�O��qB؊���s���s��r�?I�"�2^�����}�I����F�$�ޝ��!��0h��E!v,�7G�kw���L Fg%�I�$����I$�P�k�͍;9W�MI!��m%̔9�$�DU�H���&`�	�'&�������i��'�|���&�_n���I���[O�gww�/p5�/b���ו�rdА��k��W]t��.���νq*��d��-]�Jqn��+�6P�꽨�e������dbk��ZwZt㵲��4��F-�ln5sDu��e����LmB{m�{jWsGͷn|=^��/n���;9^+�ȇ�v䣺r\s�+��d��n�n�=n9*�Za�w>�bcu\��:��������=�7%�k<�ź��Wl*ms���WF���ck=]�����jCI��l�V�8�Гu���cII�s6�yٸ޶������gf8r�+<i�ї{\�&Gcg�]	�u�dk]���h�������0��l�bA$J+�v���&�c|�6����If���	/�(�Tݚ�tm����<�Jv{v���v�U�Z%����$��;3_$�75��PI�����^��ί����Gʬ�t�I�$�<5y`d�$�^��jnD��d��O���BI$�����vX5�؊���s��W0�s~�\��l %]��>Ē_�Os��I!�ъ��,/m��vz2MV6�$�9��B��H]�B��F�H$�C7ѷ����d]f*�|�s��q$�lyPC���g�s\�]�3�E�G~����K\���Ψa���Suۃ�9�
��%> -�[�V׾q1p����jx��$���&����H>KĽ�:8�.o�4I��W7�&�o�l��� ܯ3���u�A���h���v����Tf�/�hє|��!P���RWr�ݎ1�i��M�eW��	f"tt&�ԏv�B/3��jֈ��]uɍ�	 ����;i$�z7�RK�Ύ�T1�!/K�{H4<���Z��ʮi׮w\�A���sh@����U��s�t$x��?"�Aa�F��Q����L���w���\�{�w.�$����$�|9j�I$��zDU�<��(Ě,)�MW:VVs.���6�I����_%���}��Sk>kV=�PI/sv�A$�Il��{�wm�E�˥�T�-II	c�Y:���@c:ړ�ʢr���PZ�#�*��k{�qHڂ�A]>>oZ��|�1,�	$�N����]}|����j;��z��7d�֙���K��(k�T~���g;�=�Oļ�J�,o�Ȱ	0�kƒ�%ӷ�1$�ܚ��܏|�_{\��Gm�nW�z�s�B =��ٽ�D������d���Y�Ľ�гR�Q]<��ӖկZ�5�3�!�z^r@l�鷑�r*+[4g\���+�Z���5�%����̾����xd�:Ӻ��ro8+��{6Ós'^)�O��f�kcR��]j��l���i��S���_V���lC��f3z�o;4��5`a3��u�ap�{t��xa����Ѳ����Wێ���R�+3/�W��L�7����\G��4�'q�XJ�Id�����
HMY�p9+�v�N���%V-���}{�cůu,Zq�ՂĎ����O�f�\wEu���9tQ�MdT�G����G=��Q��J�a�4� �˪����3n�`v�U�5������[n�ǳ�i��1���+K�����1R������b�E��x�,f:��_�[ɨޜ������T�j�άgCp�W���-���-!�2�u�9{��mEa<,��k4�Օh��w�Ro:<���kC��K���U_GQ�`���mB��|�3��n�er�!��Z���U�	f-]nRG���YX�>�g(1�=��9���Z}��MئЈ㔂�׷\e�����'�U]L�����V�5��5'T{�j<-��)>VG'��L���8J��W����{�����c�[���"G6iM���h�1��u��F�mں�]�:��Ԉ��	�����2�ݗ6�M�:Jw��w�w]�¹�ѡ;������d�w����r�t�/�MS����7��{��6�omʗ�1�5���U|ѱ���7�E#��p���۲NN�H�B�6�J"C�,�u�8]�tI��vhL�ՙns�N6�e��vdαm��)���,�h;kP�:8gk�;-m�h��bv[� �mj(���v����8%�V���c��h@HI;;'(.6�۳�a	6�8�Nl�ps�!���Ȝ�l���E'E��)m[��8��5�&c�a�D��E�Dr6Ԣ�9-�IVu�!�ȉ!���'frum�ݭ�Pᵓ�t��s�!Ӄ�8Dr����fNqv�ۢ:'!8[ZN�H��k\"C��I;��H�n�$��Ȓr���8��,�'}��������k~/��b��=�w���lZ5���VU�:���y,_��_|I%���<$��H���I8��\ƻKu����/�L�G�*4��p�c*��g}�ؒA.7����<�z�ډ)���I$�v�f$�ICy��,��������~۽�Wv�WkWn5��L�黳ɺ'�lY���ra3���Z�;����-��Z�O|�8{��������> ������t�sZ~5 Nף`Z($��{0�wĊ`U�̫5�xH���$�R-�� >g��x~$]�ޒ|I$�9�A%��^S��mb�(�OAB:$�G꿩׻���H�o7�y/�'��v�4l��a$>I}��ل�	 ����@{ݬ�,R�Pr�o���s��W��Cj��0M��K/�<ľH�Y��	��N53=��ݏ��Op�����Z,I��ZդP��2f��Hx��Ӳ�R쎟���d��5P�cyi)/�;�O�[�%a�V�7��+2��4��m	;����]����Q��7���(�I��sm�����eN�a�&�K����>���nZ�T�n���a�z�wDFk�mN64/*���}zN�_��\}��v0+MpQ���H$���ǒ	$�u8�Z�>򢤘���� ����P�U�b+-w���S���.��;,Ò��N�bA%�K�q�I$s����'��7�wd��vǻ��R6��PWXy�]�� �3���H=�����/�7BK䒇;��H,���x
�U���[�/od¥oe9�)����Jbt�$�k�޻I5��zL�|�xNJ��kS�Y����a�E�l�Fs���O���!�Z[ݛ��Τ��ֱ ;�9��� ]���BT�=G9��̅K6k$G.�X�5B�B�r�>#�N���h���y��U�U�����l��Ҙ�EEޞ��VI�2d�&��ΊWj��j��GF��݋��Z,v��g���= 8�m6{x�݌��	P�n�;e���rЗ �Gg���A���tt���[i��f�Oum��[z�L�ҙ�9�u�ۑ�=�Qs�t��۵��m��x�q3��S�qG�p�uO.�@�0(�d�q�l�u�o;�՗��葸���,���'aWs�:ˬk�_7ncv����`�׵��\a���u�n�֭/g����-�H��}���P[%��Es^B�7�ϰ9�\̤������KW��Sq�#�߼O$��^��B��H�J�t�]���%�No����������]����I$�wof`I|�}ۗ1A�M�~���2z�Wh+*��D�����Yݼ�bI�y�'ys�>�ug{��I)�b�A%�wN����9��ؤH�.�!m�;#{�i��wa)+���_$�oN���	/���ư��x_y�w{İ�Ssv���
�U���Y���̢O�ֵ��/����
�'Ě�|ݲI�wt��#�~O^�{Z�o;�Gvp'p�r{����Uu�̘1��K�]�����6�+Eu����~B���������鳼�?A �~&�V�k*�{�	=�;�z�J���B�ȸ�� ��ξ���fª`���F�1~����Q���0��)�jWO놃�ۖe+Q�&)��xʒ^[�U~�]���1�9�n�l�A���9�n�ͬ�{�9{ěPi�=� ��K�{͂���H��=n�=�;̒H�=~��36�Wh!j��f������]M� �{g�Ē	���z50-�X����
�w�*�f�*�gܥ��_o����.9���,>�c��xx@ޞ��h�����HuT�
TQ��;v1��u훩�"��Zn=�N���X�v������D��*��뙙��H#��~$��=$nu��C.���a���x�ΐ�E-�j�s��qcO�ز��5v�����$�r��	�ѲA$�e_���;��LE�d�؈����;�����ܵӠ��b|}�+b�M�zݣ^����O=�>5A�R�>�l�ü��r���0�s����:�֨������ר�o!�}J���v;�xP!8&nt�	�NxX$��=��D����h���;bϜ��pv�$��)@Mծ��O.O/%j��g�Ü�*9��WiwWU��̌�O�7����ʻf��n���w����;�g�ƾ|����]�TNEF�@5>W���e��ƒ	a�89�&0��,�d���ަ�3HU�B���P�}��2I��<�h[.E�fO}`��}���P�EP���T��[����kٌsS ۓ�����`�/#��ׂ�S������
��i��]���:oO0A�,���Շjm@A�7�$Ӻ6	�-q�Z"����潯j�j������'x
�Nl���<�$�pۛ���;�t�y��KU�v���w�ݬp㊏ۆ� �k��kLǹX���)�� �qypak3��-��Re�Y�7}��3�6OԈ8��($��G���7@P�NU�~�d��YU2�%�5��?d 7��^`or!�RI�Ǟ��+`������V�cN�V��8�.�s��*�:Ń8��q3� ����߿��Ѹf՜nl0A��`�I���"�1�w5|)�0�U��|H'�Ѱg��ت�.��3=� �b����Α�����~;;��?p۞	�;0f��q־ ��'�%�"��)7���6H$��, |5x��~��Z;-/N 
���?�w9�{8�[p�r��Z���wӎ��+�Һ�C�lL (
㏮��{ڵ���l���t�{{�S��N���ywf��ж͟M��go����c��~_{��`�����X ����v�ݲ{3>�zx{gn���fL�+�8Z�ۧw]��-�:YdaX��J��N^�^3�ulnI��4��U�E�~5��=��F��D�䄲4굷QTX';�B�6g��M�j��mສ��Z7��f�bH�l��.��gBޗ6��<��󷇣�_��b�w)W�[���]����`wW�M�:ϲp�vxGc˝p읹+��;g���^Z����mۛ��*G)é�<s��;�h7[k���n��,yؽ��g���0��]uGu���9��9��^���䳽�j�����廝���!���g��D��m'W?��!X�Yָ~O�pPh*�nkd�t��Y��=�4��aM/w����o�gusK���	U)KL{&꥚�X��v-6��A@m��P ��=��c:!���'V� ��w���ۂ�ƪ�̻�6�{��cI��]W�P���}[�	 ����#�z0��O���!PdRl{zG��KA����N�`�7�����eU�����u���t��#��դ罾�}�w~�&;���K���@P����o���{Y�k��n��nI��$���h�u/�s�e띥윁�m��u��.֯�����o�	R��Q�y�g���n�6I$l��1XBU��^��5y�_�9���h�V�ZUIvR��9͂�*��hY�j�C�����U���͚��z�^f��{����pߴ��z��%7�f�����tq;�ܲ�}Qz�Eݦc:�	$����zvs��[���o�[\n��_�]*�*�i�j��u��w���>�B��%��ӻց ��o�I��ٞ9\	���j���p�9�jٝ��- e��t �<�@.i��d3��Y�{����@�@]�I�Ϥl�0�o��x.�ݴ	���� �����5��)�,��6>�Xr5$nF0-hek�V0
����aՍ�;aFonC����������jŊJ�p2�5��n�y��'�~�Y+��W�����Ff�`P�t� ��V��+7T��m�>�� [�1My���	���W{��� ��YB�;jGF��Op��ԛ��m>}I#k	�s��`��|,�^���Ìk�}�>�G)`��ý|��A�z�8݊[u\�4�j�w/��[U	���s7�]g�8e�M��F�*�&w�9��k'����NKT�-,��{|�o��[��2�=�G�Ӽ$�ʳk��H1.L_jt�q�0�|�q�>�.i�l .����<�(
��.\��R���l��#`�a�����l���nQ����X�īsϬ<q�c+���Zw�n��M�s>�kB�>���<�{UDJ���k��3$p��� �OO0C�]�B�g��.��z�>i����ʵ�x�6�qʪ�h�={��w�� =����a �i�7��`�g���rE��uu��E��N1](����|�u���v�ttpwQI�h`�9�`�@��O�Y"�;Xz��-���^�s��VIf{}`���� �ӳ��<�p�zA��F�c��<i!<�e���?Jj�}0���>3̋��5EG���_I�f����Z�-�H07F=���wdF�V׬w�����*�U�V���[uB�n�� N���n*L�{�H����ĀH;y��<aV�>� ��8�;��2���O0Q��4:��Ζ:^�slz�n<�ܩ�7UG���Dm�cWϯ�׾�O���G�$�~��̓�Y�v֊"�Y�+糽�éشV�4����}�Ҙ��\Gk��'�z7�$���� K7����,���^x�MY�V,R������� ���0H��O��Z�����:��H���$����.�/@�"�X4P����Q���mq֯΅/oy��P�;����[У��^�W���o����,P�:�5d����_w�y�H$4���:�o�he����7��cc1�{�yH@���	!K�P	!K��$�	(H@�� $�	/�$ I�	!K� �$���$ I�	!K�$�	/�$ It��% IV�I_�H@��B��@�$����%�$�	/���%�$�	/�����)��M���,�0(���1�0   @       
  B�T �    P �P 4 (     il|  [�$��"�*����  ��	
 �
� mb� ��� 
H)T QE((�P ��                                       �      *�����\��*�\ƥ�Ԫr�m*U+� ��Jͫ��R�hqj�6B�C���N7 �TS-R�����U *�  ʼ�QW�\�
��t*���F�siT��l���\�"K� uR��#���l���#�*�y��B�)k�ki��          7�J��'m*\Mتsk���seJ��p 6J�Y���K�R�Z�rk��(�� NJT�3�=���)Ax� �  �, �� .�  �`n�� ��4�� <� 
^�R�P ^� $(�f�`4.a�N r�)�{w��
�E�4Z  �      @ �P�EX9��@.`s0Qr��'�@h {�� <`GB� h@ � #A��t ɡ)Iu�"��   A�@d 4� � 2 d �# ݸ  �ݽ@� zw��B�4             8 P� ��C ,  H�C 7��@ �  H��0P �W�   � ��d� @C  �2�G 4T� �F �2 ��� 0(	]x  �         	@24 2 �` `!���G��C- +  $2 �(U$P<  z� �hL a�ԇ6Tv��Uū��*�� ��I�/6��.�j��R�� 5O�&*J�L��4�S�M0 �j�T�=OdP(D�*�IST  ��T��jb�T�@h2d0�I�J�4 GN�����vƜ;�����וm����E�x�L�b�(h�y�T%	*"�BP�BP�(`R*=�UJU˧N��<n߶�i����㝦���NE�������]J�C��N�I�=};�-�r�l:N�h�E{Y���T��i�N��nW3z7�;��&P(y1�ve,�~uIA	v=����F�3�����D܃w`�:YC�g<[+ې�dZټ�s�:�����fG�a�Q��C��"@��0R��{X���Y�����6��9׺\����ZL�:r�I״ `����,��.��A5�E��d��]�L��QᗟWZ�!���B�Nv�$"�vsMGӐwAHh��p��������&:y��@����:f��:��l�om�A�U����Օ_�dZ�3���Į�H�f�{�>E���М-���[͗<��=�,�;�����d�,�NkI>��ɇV=�v����6K;�3l�Lnw#^Ү�m{k}�\k��s'7�����[.4{I�'���cp`���-��>��Iݱ�,�c����A�ez�<T��uec���L�L1�v>pr!����Ŝy�Q������3�7���y��wKA7c��wS�%c�� r��FK"��v�k�5�*���8\�QS*Q/LG���r�Oo̵���k%��R����db�D��V�5��J�餝Z��^<� ���i��~$��	9Z�򗦣n��eyؠ�d��XU�:��\�Q�}��Q��_V��e�FЍ��m�GE�v��=�k����SRVJv�R!�(��c�q^B�/hyeK����V�Eݬ�SX86v86>�\{�v�{�����X@9�^O4U@�M�Z�n����Ids.��AcX@��ó�5|wN�]9u����:Z�� w���&Sm��:�A�.��4�g'јS�ˈ����F��>͎��+W?��4�{Szy>�[�2�ň�mڥe��K����ӆ�{$�Ei����	e�
;�Cr)K�6�=$��nm|�>��彻�s9/�q��f��ֻG�4Oh��ĵ�n�0$EG]׻��9�����G)l
�W�h\�f��df�b��� o>�y8�v��;YK���(�W-g!(nLm�@�nW�z�%��{��ta]�͉IN�q����ҹM<jC�����`v?���JIo��y���� 7�6zU�&f��Ҕ׀g2nb�HrK��H��j�:%���X�uZ��c۝��<����Aۼ{X�]΋��gV����+0v]B�����9l͐��o��Z�s���!�(�3jg�YŽ�L%�Ƽ_^�_IԘ X�
�'k�Wp�kP�����od�6h�;q9�
w^ższ���9ڰ5�k+s^@�崾8䋹��nv���p˱�ؖGd��H�0����rv՗��nUVTRn{׮�O]���˲�Y��0̆��ׇ~"`�@�;_u!�R�"G����w.Yf�(�/n�����@����@�E�k�9U��w�J��q��Y�<�zkq=�f�[�=��z�׺79V�k;A�)��Lm�ɛ.,��^���ڵ��[��{j�>�fņ��qk��^�"]2���F{x.rއ5[��Vt��i���Ռ6=b�S�"�S��Â��1ќ.�o]nm�7��qW^�e�gf��w�d�n�e�l�g]]�oVm37ۍt��Y�����a�@ː`'U�����~JG*��K*ݮ��γB��r��J�I/x����t'������Ī5J����F�c��v���e�`r���6M΃{�OP/1ډ��A����db�����+M�ϒغ��<(r`��d8�a�D��͖��n��eB�3y�4� ��b��a��򝻈{a����IT��v���{e�Q4_<�!�4}��}����5x�v`X�q��{��Yђs� �m���5�b�w <9\ү7>�������4Mg9�1-��C�.�c�{��R(8�� �{�ܛ3M��M\��'{�&��	jp�r��q�5���1��'
G;̴/::�D�5�j}YE��n�s��%<��5VR79��h��E��`���ˬ(B׭�9Z�0-c�#��IO#0PY]s�XqqP�A��^G0G��<�rSl�qwc�^��X+`�p��=C�zK���6ݡ@���Ɏd��e�5#4�d듮�ƒ�L:�FN�y8�qn#L�&��CWGC:��Oc�3�=�m����� ��&��&��s�ɝ�ȂMtĺ�&�!�{�^��.��vqȮ@x �!���F5�u�� ���"�՚֏�4U�:�eL�	�ٴ��dY�nK�Ŏ�Oh����:�8�����o��V���p�49���nCWod��D����$ �
ǫ`��G�	������[��D��������Z�ƛw��������<�U��-˻�v�k�A;^u��b��t�ocN';܎����l��S��	wMs���'Tvv��r�e�ؐ���9��9k�[�*)܂"������=�	#���g�O}aͮ���%|3S�#3/n�TG�#�rh�x������{D��Jkf�l���F����谐3FUA��Q�_!�[�����\g��i�ɭc����r陮������A�ڋ�8���uAq��)e�-�.u��2�ZP�yźV�f�>!Pq,W �AqKwq��u������2��N�/uU���$�8՜��-���I�+IH�݅���	��@��x�'��	�2Z�Ga[�Z�q��N,3eaG�d�|���]x���Q�3qv\>^z�U�8�IE �m�Y�f�� ���]�-X�i�n�ň��v���tR���[ǂΧ���D�(ޙ$qu�@ݝ��\37���vy�ෲv�����Su4����p+�˚��<��	T9�|2ٸ�	�\������X.v4*V��oI��;���,�/��:�{�r�c���g&�۔V:�X�G{w�]c�X�v���ᓙ�DRP���!9�O2q��;�����'ܩ�@ξ�e7��Q�n��%Qܷ�J�d-+Q�ˣ�wi���~\����MЌ�Y�
�T�f'H/0��� G!�ay�$xˀ�.�Qۖ�K]�gE�n���1*]f��Ul�H
�O\Z�O�GH�:�v���%��0R����ä�J� o:��r�_r���q5�ь���FI=p�Z���Gr��f�\�U���{{v���|;��%	���d����Y�`��8�ζ�V�T����J���N�k�&���m�s��\���{Ob�����\g�kgRx��:�����9zt<3Q�x������`���&��i���^��MY��k���p�Рy��ǡ��Ap�rv������I�"�-�a0P�w����{�P�4j�F�	.i��ٳ����ݢ\��2��1��}�9d��fp�v���b�����"p�r���.�����#��>��jt4(D�W������e�z��NەC\����ݺ��{꛰0�bf�u�VD�>:B��;��כ�0*@�]��W<�_H5s�;ӌ�H�z�(�R�}���K�f�\��ƻ�Ɖ�LK�57��:%g�<Z�v����[���t>7���a�\�ɻg 3�\��{��7�V�u�9�i�$ZX5�]p)3��i�{�:#SHSp��,7�h�=�,���OӧNP�X���v��(�ɡ��q ]v�� umCA�#5��T�YIh�-�b���Ywn#��k��G����o�W0���D\�h�y�M]սv��+W�8�Ӈ��t�͇(�:��a�3��T�p�,5�� u�#��sh'���K �Ί�Je[�!�ynS�#������{v���N(s�a;�ͽ{��펙��z�<�V]�����m:��:��s� Kf$�&�u几mY��6�u��p��Ҹ�bF^�PlDMJ;��0'��EU��tj��_�a� ���6�S�yvh�[N�����`�׊�d�˲�D�9� pǋM� x�L\�&�F�y�iW9��$�#
�rg5i�*�u�ۚ�	�� {Y�j�&$x�k7U�]�qؾ�f�za��`-\U�6Fs<�9�􏳩9���iY�pJ7��9\���@	-��k?2���Vj�{���9�-��E��=�x4�m�>�"�D��y>Üdb&w
�Ql|�Z��M�m���[9HK���&UTt���^����//��?��@�Af�ޑݜ���"u%#l��mv+���0F��hW8�&w��n��	P:fݼ�Y�8m��q	�pG��A��Q'U=`���6�ʾ=�Hڌ��v�"
�Gu�$�Y���\��E�H��W��1��*8$���F	Ru/5\�<0���yS���v��#�W�M1�B�
�59q�����s�Hڰ1V�U�}kV;Oku҃�ȳ�܅��=٤�\����{C�#6��9�։�X�m�ܽ�q��@�C�����[�{:� �$Լ>1���7#�n	_%ϔח��6:��ٳ8׳;�7(܋oFB ˱�5��wB܏W=;��J�q%� �'��#m%M3�:����m�<9T[�Ɓ�0ݏp�+��	uq}�xz �E�Y�|�h�3����y�d�rظ��Ǣ�;�gL	�Ę�=9w�lKK4�^*F����nK���6���P�,yw�����hD�ɍC�k/h�\�1�4������Oj�A�0�����"n�7uJ:;N�YǷ%��L��m�v��_��WY0ܸ�ʄ$|xd�m�Q�7�t��Q��x���˻p���6� ^��X����J|
P-�vo0���u�-��;^d1����r�[������yh-}rދ�����4�dś7H��08d��6���R��t,�+9�u�t�;n�'� ӌВ�vQ� 
4dR�A���פ�gnQ���4�˶Vh�7$�M3�I���ԻUq�&��߲�V����]h�n�:Dm�9��.�}-,���s�\Ѽw
쵡S�X�JA�Fi�n1����[�䄯���t�j�l�r&����^�qN�19�g2h��`G�i�C3j�1Qg�cyg4;��)�&NUŸWZ�j�6>w�ތUuFm��&w�=�����!��"���*Qa|',MA�u�O�X&�[v���^���:����6�����or�@gn�؎��v������8vS�^�¸]@E��:h��9q�[�
�Ğ�8]3oZ�\B�e7s��4iW%[�A�1��o,n��8Lv���i��P]�ݨ�rF.*хW�ܪ}h
���!c����v�-Z*N�b��V1ɸD#b8:_���.��ڐ����@�
�$!���sN�ze��S����(ǹ��`���������4��Dt�ؗF�3����J�S��V�Fo1�\w7�d�S��}^s�.���}�Gn'�я�6��^ܭ���9��sk{l��q��x]���yzs��>���N?mكSzy��/��,`�F0n��75`%ܦ�ը����t?��Z3Eݝ�l��[�Ud�)Λ�¨�t8�Í�l\��υ}>J0ވ����7qC˦"
{��S�BA(#Y7�@����eӚ,enǴ܇����dpM�p�ɮQ�'���ʕ���o��3#[��̰�}Љ%6
�=��Q��B7ܾ݅G�q݃����"�%����wU�:�8M�L�C���痻�s��6�B��W��[�*�OcW^��>�OK-�c\����+	�k�A!ҧҘq�$	�z�/N���_����:Z��fMc��d�@]�EO��U�3`3S�(qr�V�*nsZ&u��>.@��1����v���od��M/��`��%��=>�-�)�R�4�ç&�m�P�:��E�5�rr�h}��T��wa�zgw|�BV����iE��t���ସ�qC���`o�^�@#~w�D#+K,L*WR���{�P��@�3��;�/f�-�hDRM� Ӊ�g=絼�IV!�â�L��'6c�W�Sv߇i\9$-�4��y�EU�VN&�i��\q3��he�c�eP�͛�v�Ɇrv�wp���Tl�ޢ�E�a/r-zs@צ��6�0Ay8Cb���t�i�N�Юp�N1�s�u]}ۃ�Y�eUt��zh�	cyk����w�,%3A,p�]X��:n���)���i���{�6Io1��յ��[gS��Ն�E�lܯ����'����j�;���.p�pWۯ6�P �I[��Jf�m�6���	 f�Mb�ǁ�B�㍸¨�Q;!ܧau��'�
=�pւ�q��oT�˯�����UA� /j�8pα�{������e�G�}� "J�Ӄ2)R�!�@��4dרL���]@\�"���5� 3Dx(8��byC�����FWÍ�fN�d���\�N*���Pf�]���R߉��\6�>�	�?� J�	$P�(@� P��(�H�$����
�"�� �T�R%BH��BE *�*BI��$,�HX�AIa$�H�"��	"�	�@$�P�-BHd�d�B�I X ) ��HHVB���d��BJ�d �$+$ R"�I`@�HT�� 
���E$�BHAa XH
E$�HBHAd��@�$�`�VHB�	�Y$��Y$��@�$�)$Y*+ �!`E�"@�a!%HB��H )!*a
�d�, B ) �HIY�!����'��g�}�A������4_�L���C����X{6}����#�pMm�l+1ӏ��^�n�əV�cӛ��5b�;��}�ؗ�2Y�P��`�k�#CG�պ
P��]��i	 ���q���Y�!�nչ�:f�Dp�H{<v�;dOz���S\�����/M�������%{{!��xE�������wy�I�2t(��p.HE�2f�m��>�)��w[pM���ú�|�*����90���ڃn�Tz3B�u�BTP�z��{�����whӾ�G��r�O���_-f���嬋�8�o'����O��������k`�H��q9xS�@�	ں\�M���>����9f�6�����s��	�b�}t�0ZX}A���ٶ�<7A�]���K�〽��GX2�����!��\K�Oఉ؞Y�(;�F�=1����1y�o�LIB��<ϡ��np�犟c���^�XWec�w�!�E���Z&P�vy#�U��9�	'=��y�v_dW�\�K��}��!��䑮�7���f��w°[��-���~�g�C�g�¤��5ӌ�-�� ��c ��%xCV�H.x
�O^:��m�ެ�w�i8�>A!���*f����o�m[�؞t�@�T���O���f/xt���ޛ�y�cߖ1�o�� c����oo�)�a\��f���q<k�;��;/�����1Zϧ����k��M��-�L|�j��z����<�}�k�v�Aa9����8t�A�1�}��G�vo �^�}�\j"wZ�755U틦���E�t͐�x�y�����Z�]�Զe�įM��HI(��{C��FhDH�M��m^�|j�C�ӔZ��B8����v<޹6Km�W�ϮF����<�篮z"@����_��ܒ�>�-�6_�@��y��g��X� E����� �{~��+���H����Y`�kZP���J�b��Z7���Zv�μ���n�ƍ���V�U�q�&��n���V-�B�c-�bt:歖v�
)4+c�N�zI:�{nj4*"nj��bqW�~uf�w[,n�nߨjSAL7�ϭ�lF(��jl ����+��~Mz1V��b�w���|�ڪ�U�[*�HD��b����VL*g-��8��h�@��׺�9lSG��t؝b�=n��]�{����=|Ϩ��h��gnK�G��yڪM[�U��<�I�����%a���m� e�Z&P�{�I3��BM���:n��Q��f��mLj�Bu���s1̸�J�T�_�f����R�B`$Vֈ+>S}gM检�� �Q`+^���r�����r���RR��M����r��h�h�����:����pz-���DD��U��0ƻ�(��h�yK܈^�&��z�����a�x}�4���Ph�������E�<|<|���
���Z��x6�Ny/d�N_4;D�}�Hh����g�j�Y,�Xe��P@C���m�E�Z^�=�f���Y�[*=����ߣ�i�۔��2��۽�
��%�����;����i���)^� ��"tȚ;����V��|R�� ޢ���5�rj�}V�)�v%�ٺA�H���z6#~����Kx׷ůn���0��{C��&P��.Q��P�q��Fg�/H/|�b����a���Oz��
m�=�7.w�{�ޕ�/�C��3�����~��~g]A������mI�*����W
����K�З�Δ��y�.��ɒE��H�be�>�t���K��o'�}�-��Eqo�30t����=�s�y�P0d�6v�|�[use�ksY(�u���Cܬ���u�'��bKۊ���5���qי"���,ݛ#l�2sY9���T�{6/�T��>-�,k���*��k^������};�����ѳ��t�=n�*ެ�[��L�Yu�vwIUi�(�v�T�m�*3<��7_�ט��Ͷ�U2� 4XV���y,�U�^��<��n���qH�vn���G+Y�u�l�-��s�vD�zb��tI,C�s)hR��԰��]�V�nס�b~��}���A{��xv�=�ѕ��{�?��y���p�����{�=o���;�"|(Y�s_�b��E��̆�~"�{x�ؔ��ܰ��;�	)�{��w�������ס��NPH��v���ǹv�@R�̥c�}0���[���S~�2	r���;�)�hv=�by�x�[�/=��SV�B�o5���n'���n�O��]��΀e�����1�R��t������o�=��Lx ����
��7�����|ت?�ǒ�^���=���h��O�&rl��ʩ���|&ǂ��'���˹�ễHn����8rO&�Pey����{��C�u���ۈ ��O`,_}ֳ��{��������ž�'�Ly���l���:}B@��1 ���qx�C5��.��u*��FW΂;r����M9���gFs����gR����X���;n�`ܳo�3ROP���������r�)y��UX�|�$&��6����dĭz�ؓ_�x����v���wI��w��07�.T��ԱS�u5�y�=�{@.Û=�a��T";��s�>�E��;);��l�2����w%�|�W&CtCՒL�X)��mx<U�� ܙjX�P^?T�˯:���FbaR�}��Z��Ll��A���0�b
x�G�׵�jIG7�>��/b��3��Hc�u�a9G�)��Q���:>9���O�}~ORF�E�\��zn�~��Hb�ǁ⾝���\u�g��׶aC�+��p�>�C��#7K6(W��N�ĩ�Ӿ�	ɩ�������#��v}U�^�ݭ�C���:<X/Z����3#��� ʇ2|t�L�;!؟#�a� ߃��n��.���Hհ뛇�~}ƣ2<�6o�ۉe��w�Ս��fe����ü�O1h&>�h�i�	z�C;�8g���ӭ����3{=��P��)�鋹IFT�z�įj�-��i�cك�*��O9�������o^��S�__a�$
��[v6��a	�s�Xəu"wC;�d(���_%���_{.�0ǧ��YwV�ve��=�YG��~�;�§t��2Q�8}ּ,�<=��ZnK��4�+��Ց�z ���s;V�	��%����cm.+c��k4a��!-�{&��3�OAίEC��&�r�&�/@n�ݜi�������Fu�<A�uz�`=V??h�y�jyEO�᪎��%Z���z�/>���o_^Ѻ�1L��� �X�ǲ�}bZ=m�Ӛ�1����1���@Ͳ�>��'�K'v�ëqeQ8[��ͷ�e�؍�^�hQ��B��l�E�����7J�:�M�V���K4d��]����ޜ׭{B���y���C�Ǖ�»7c���W}�x����4�CK=Q~(G�Ŕ�^�CN���sT�ڞqk��b�����엵�C��qQj�^�����2��:Y��g�zk�����Ma���ٝ���*��B�0s3lA�꟤<��l�\�v˼C#|����7�(~�6m�vz�3i����0�����k�\|o�y�Z�}��>���7H /!x_a�PY���ש�aW�����z��w{�u7���� ��FR{�şd�ͷ"���Y4ּ��1^�������+�9�j�/��ޱ��k��N�>Lgt����|]���q���+����;�r<�e+�}�!ݴa/��wC;��47L�I�=���O����\W{Fn�^%��\�x !ޏ�/Y��|�	����ʝM�������yv4�^�h�dy&��3�v�����H]�v�=�ёz����2��h��;��[���y�=�P�f�o�Ke��v���d�{T�K@��}wv���i;��$����O2�-P����s��y{��z����<���pˑ�t�=���������+��æ%����o�=V)���$���5���䞗�5i��B��j���ڞ��Hn�q�wW��^  [���>���Q�O��~�w�Z'�����Gw&��Av�T��׽��+-�h��+�׬��ޞe��+E{�~&c��X��'��>��"�/'��k%���|��<�u��[K��Y�W�����r��/5�*á~�����2���\]F�:����2a�r{�.�3W��ɶ�]�>�����{����xv�睶�]�*|4�}B�]6v �^{5Ե��w��c�.~uoO!5�����1^��e��p-nu����n�B��ٹ����{��*��tỖ�����c	N��x9��f�����K�� 
��ec}Wb�� x|@v�ڟefd���Y�{�vɅr�݊f��۔�g���Ɨ�z��厼;�Ը�w�^�h�˫$�5d��ϱ�Cm9�9;��3��LOL��{o@�n_%��jl�n"5H�n]��.��}2�j`q�i����ǽ����H�,u�l5�&O,�v�'�w7�͗u�=sk`z����\��j5˷A&�܋��ޙ,Qp�%�w��J_��*�4ۯ*X��C`���q�l�?v-��0�Sw:����vh�zU��G_�ܡѡ^U�w��mc{����Zp��y<w�v������� 6N84t%���p���c�^��b^/]NY��`�Lw��H&�5]�|��]�^,���k/!�7�����'��3ϯ����x�
������(s	:�5�Ν��ξ	=��ý�b�<����4{$�G����ڔ��h	6��9u�y���҂1��ǽ8�'�?�g7[a��+Y�wt_M�jK��z�7ڷ�t������yF�7ړ�G��s&t�� �|Z�r	�Dk��\�[ڑ�����{�捀��]�ex�w��m�f]���$�^�	��i�(�,ͻ�ty`�^�Kiҏr}<sk1Z���Y�eoA;JX�εq�3�@���{`�������7��AT=��	�<�/���<�m�	XǛd�+����|��=u��﨏7x����Is�$Y��Wg���y�f���q���U#����si6h9,��;7�.ͣ��FvT��ˇ�,L�1���w��{�� �w{W�}�۹_��=^��8(�y[�K̚��D�d�����L~G��� %��
O1Փ�n$&v����0���+ϵ�l)�fxg��g��ph�|�T{j��v����<�:�_����Y��5�޺���"U�m{{�ܝF��{��d1;�<foo=��SP����-x,���H��ڄ%{�iP��g�p@�{B�(����x:q��^j���b��TPªЭ�Y-\�F�M�������o;~���{_N��_d��{�EPj-l���Z��L����ч[�ױ���&���xD�7Y�6ƌ^�r1wv��>��zFm����cB�X�>Z����"����D����#��x/ik����vu��>������M�]�Ϻ;��uc���]L�x<���Nұ�]�����B��sN0Vo��a����ࢳ�e�Y�hשv/)�\�m���hޜ�p슇�7���^(��6a'4� }�.=��A�je������}[��'�������r�;���zJ��{oqT��,' ��[[O�n^���9��i���x3�7h�𞊤�zOo�>��g�
�wZ=�x%�@�߫D�6�&�G^��[œ7�S��1X�����I~~� �]��E>%p��a�`��E��r������<9-�l'w��?nmZnsb�kV�AdSyf��5�ؼ5i>0J8n����(�3<�zo����Ho�F���sw,�%;��5N��I���M��i�������$��h���(��%��,�q,0K*xV�6j��Ą�A�c�"պ�t��=��[�ZY�.
d�x_?C�"/��N�t�R�F/�w1�z<���!(���D��Y͒����ؠͷ�W`�y�oB�g��3c�����3o��@�б�X��i�x���<1�w�W��� �ݗ��Z�U�	�;��];��m�)��!�F�yK�/U0�x��]�3��^
�A(K�Ɲb�K�L�U=0��\�����g��_RP\���rt$鳒SW�uާھ�[�*]�z
�o}x���L��,g{����UKٰ�,{��[��L�p��p]��j�S��E2�W�LY8]�����=�;da:�┽W�W�7؋��f�S��{�f���L�٨��k��q��)�^ήe���)��.N��ӛ��6K��ޕ3��%3��Q$�tJ�ܿM�]�2m��G��74���Y�ԛi��9{�j��~8�~�y{�T�;��p}�7�J����ڞ\$ܫ�]�H�1��ؗu�y6,��sFiS�F��9��k���T��f��e�;���#|`�	~�/��vd=�Ru½���%�;�7��y���uz�j\��������꭫W=s��ыθ=<8�};F��8������w��?�صw� ł%�8.��*$n�z�p���Z��t����5Ō���|*S1�Ԇr�����ڀ�~��7lᴾ�b��h8)� ��<�{��DڦY�u�m �%��#T��9%��x�;Trz��|�����;���b{B������	N呑��uN'�y��@s����V8N�7�x�j�OZ$�����xt+V����o�vs�>��6��{!����i����{Q�nOyH����IU�2��5���8�ڭ�����X�*��7�=/xq�^�����s{�1��Uŝ����Ú������$ I)$���Ύ\��m�냧�]:Ƈ�jx�9a�\��Qڇjsܻ�g<���r#Ū�sFl���uX��!����f��t����s���:;����SN��e�OX�X��<[�}W�a� :��x��v���cy�9Ay4����ݰ����x����pnc��[u�����Ш�[�nz��.���{Dݫq�-�ρD�Uv��Ѱuv��u�B����͒��q�������U�ു.�6��6�x^Z�wH���x��4m�b�)�ͺ�t���zAS��t=���b\�|�R�\l�gl��]��ݧ��.��-{v��Z��tvb�V�+a�Gt9�=�틎8��Nâ;S��m��h�@�J��n��Z�8��E�h8�bO�����&�l��y���N콮pv�uM���+��v���g���bv������v�5�.-�&(utAz4�����N�,��OF��	�n�ħ�)$�y[VN[���8��=D��VK�cz��Zٛt��m$�&�R�L��m���W<�v��Ńs]����2=�܏2n���J�;l�ӷ;�s�1l��,�e6�Q�ݶN���LF��۠�齷�=9,��r�3� �7q�����9D�tY��m�q�q ��Vuۓ	�m��gW[�8�]��G[�>\��M;7!�=8s:^�EE��Vܛ�)�t	���v��٬ϰ�)Ծ�v��p������e�]��y($7Onʜ��u �ő��`��V���1��jr�j�z$n�-�x���Erm
=�Mu�`�N�Ӂ�K�nւ{n�N�g���o&t����덷&�u��8�qf���Zm��6Z�S�l�Sڢ��N2GQ�^ƭ�O[JE{s�玀��ݫ�V�R�7i6rJ{�y�k����sVz9�,���16����vlûa��[�F��v����ms�9�����7$=>t����g��և�N�����Ǯ^wgr��&h��l.�e��\��kۋ��Ig��9�U���Ƀn��#�tk�s���$��ܽ]e��;��������|=�]�k����VWpf�So\f�n;h�F�%b[GG:-�v��V�vp4��7k���l�	��`�"���j��;����l��nxk\���8����V��F-;��1��ʯq׬�Y�nwk9�9ٹ�"��[�����l62�+��������4���\�(�z��l�xO�i�Sv�v��g�ce�%�ڣF�7X���{�㗷4�u�L����c��nj�=����ri������ޣg&���u.j4r���n��&x�Z��q�ۚ�uN���4�n1����7s�q�����r��כ3�^��ە�m��\�i�w59O.ԧ9�����nS���.���̷On�A��I�\;`�^x�h�������ۇj��Ӭ��$lJ�c�D��v]�=�����^p�׭��!�[n�ܜ�����CS\;g���uWnI��ݖ�ͻkgjۍ� 9�瓫��8�:x8|c��\����h�۲�gͽ�`��1��Ҹ�X����:���좘�ۖ������;7Z�/�r8�9+I�#�z��v�ո�h�΁%�c�77��'-�t�u������T
����{��\؁fWz��r�w�ȧv5<�n�n3���8I��89�z����u�;�O> �Q۞Ĝ�dꨣb�<W=�+!��ծkkn�MƕH�Y㱀�<N��l�cn��b�S�3Z뫨�s�;��N�ɲ�r�r!�Oe,�!�V�N-ӱwd���^܆���лt�<ud��W�뤍v�7oe���s����p�k�K����k��n���q�r�k��ɲ�����]�k.1�w:x\�5v񣰵��\mŹ��ѡ����a�x��#V!\��6&�l�6���s^�1�JX�n�N7�^�ju"]�Y���]���`ىܖ�w2��S�rn�:����6����A�猒`&͞ϱ�W��6�\v�w<�`#��㩼j��v�t]=h���:m׶n;&�1�n�x9�<9^ָ�4=� �kx�絸��F�J��c��v�0Y��I�e{:�nKq�[�g��,:"�n{0M��v76��ڷ3�O's���PC�1����Ǟ(in;��t������wm�c�{mS˳�6�6�[��(�&;t��<��!�j�맓�^�!�֞�Mݍ��ޗ�!q����e#��O���L�N���.��w`z����ن�W���Y��v.9˫��Ź]=��o�s<1k�λ'r9�o9�G���⩧����c�;O�W/k\l�㣁S����G:�V�8t�a͞����y�6�۞-n	��ӷ>�]r���g]�����\<��b��&�,=�[])m��iݫ��\ȇ�n'��3���<I������!�ڟl��n\OV�8��nc�o��\N�8yH�4V}�a���gj�;HTWm�\oY^u�׻{D��`�ad�FZ�t�q�-k�l;m�N�.a.E�ո�S�W\�9��u�Þ]Y�h�k�3��
�$z�<=[���ld#m�{!����cix&;4ݳbyй���!�������:p 3���� 5ӝA��l[paG��7Nˡ7LDy��&����X�α�í�o ��	��v�n��r�	���ʡ�tq��$Sm��������F�u�/�8n�+�ݐ�h��]<����j�G��'[ې,������cj۷M�gz�h�6�y�u��G/ih:.�]��癎y��m�-�e����^��L�{n���-24�%�T��64w%���/;���M�]OC��yG\q�ឰ�\!ZA���@�Q˶:5�::v2k�5��Zϲi�ݷO)�J�^����%!���^��V�Z��Ѹ�⓮��%5s�7�L�E���
C�Gl�w;H9�֛w]�{q�u]��N6�g�Dw[px
�f��m�ֽ���[D���#�r;�k�ι+JF���z��nب�v�g��Qn�c>��scU�`������3�)�8�l-���/l���;�ͺ�.�kU�6P�b<�ka]���$g��h�W=��si�B�q�v�e��<�{���wm!s�v�lY(B����f��<���4�]a����5��#[��v����oA�&jMmF�p]ks�#`�+O<;eŹ�:�v�����]����9�q�3�-���dƃ�����:ѻ;�v乊^-�p�O>[�zL�]�t��5�2����GRL���n7۱����ccE�k�%�����z���n��0�m�ܥ���Ok�7������^��ۇv��jbn�W8�2�{�e�jsm���s�E���F<�=s�vx���e�8����{���j\�vQ�wd�{�,o=O/=m�c��Q����m�&�g������;y��{m�ӊ������x��C;��
W�n�� sv�;��OdW��u��n�t�k9׃�.�u�qӷ��d���-��nbC����j�������Ƶ=�����֧lh�l�nyS9�=��;=��g��8tl��l�y�!��vݛ�b��]���<��\m��(.��^5"����ݱ���۫5�4{h�.[���^.ޞ�\%�;۷z��Q�s�ޗ�].x�=���.�sw �ܦ�-�E���v����n�S�"�\�܇&�V���vz��\n�۹ꃐ�bw0g�C�:�|-Ö�U���K�[��k+�]3l��U�m㇟1���sbS'����f����mwc�7�4j�7:�6�	��%9+�w���2�GQ�y���nMÍ؈T���7n�f��ێ���=��nyKV���Z:{aK��`�e�y:뎟b�x�f1��������yC�tm��9w4-W8��[r��B[�ښ�9���9;]�]�+u۶�luv�⣕�,t��9��s�����p�K�]bQ�+]<p�����w6��н���X���Ɲ͎�&\7i^��<�ۃY���!\�hޏ�c�)�1�k��d�>��q����g�������\����{<ٷW>x�e�#zp㔻�0�1��X6�b��/�-�5����E�vT3��S��V�.�2�r.5WH�r��h6�u�V�{�sB��;����m�����Ɠhz��붑�]2y�Ǟ���Z�`ۺ����y�Y�Z��=�l^�/�<���6h�N��n�tvvwZ:��p��ziv��au�s��l�l���jR(wa(�Q��9��.ؗ���n�Q��dzQ�����YH�5����M�����Q����I�wa��u��z��X���xÎg��rKb��.��6z��ɡ��C�볭X6w^���6;x����=�s<=��\��:���nM�t��j]s����r��F�+6L�<�Ȼ���n7�.k����Tw6��F^�����v3`<Inܯ�i��g<���:z[���l�N8v6{&�P�����6]�����D���N��|`�q�5\�rH���=q�v�&=����Y"ׅ�s���:i�$[i��
`+�T��<=��v��k�5b�-̧i9�s���뎣qb��8��|q�y�![w�݆�q���F�:8M�m�� �睻�C9P�`L���y�����OY^�9�+s�3�����z�܊o3�W�C��ă'c�X�u҃�8��e�F��ˮeK���[�o&.ט#�r4�R�ol7n��v6����-�Ƽh��@;����47�:�����$���c�bM�'7�m]l���>����4�]vN+��܏;vy���sIO[�f1�]��T��ڹ�����5��lF+��������.�.�aont��z����cUS�;a�;f�Z�`�\�h
��e��v���0{���{��Ԩ�[H ��UD�Tj�l*,Yj��mm`[T1Ad�Q�
���)
�Hm�E�ZՂ�J��Q-�U
��aUX��EYX,Z�ej�FDVT���ʐmR�kmU��maR)R��Q�"�AE�PTh �V�c*(�YcE�YX��J�X�m�IX�
[m(�mQ-X���jQkD[iX�T-��PX,
�X��Z����T*�R�����+
֨�X�[jVUm������,`�����dP�eiXT�+Z1UQ��Tb�##iPm�*�XV�,��Uam`��
�U��,�l�Q���ҭAH���j�%IX��Y*�d����V)Ҥ[KZ�Q�"

����I+ �����(���P*"d�I��337�B�����mɲ ���r>yH`]q�-�2���.���-�C�#1�ٴg�������>WTu���5����p.+:T�]Nn��"�MvN6tl�N�庻���l��/��lq���ٴh�c��]�v��9����눷7OXy�絽�tKtv����[��a�ǎӲ�%�����ȝ�~2nlG#�.��\F�7e��_^^[�%�#c���A�vy��E-� �vy���V��;F��t�e��xؼa:��\o
���'[��k�����k�]z�����O'�ά��\n�n�Y�m����.c#��\sg#����j^ ���À��m����Pn��ۍs5�h%:��4�'n�	�;{\޻5���ٛK�]�H��$89�X��x"��������p�Z9��ܤve�m�B�gv��iy̓sù`^�n'z��k�4p�m6tz�ux�c�]�����X��r�\REq8�,c�O˶kG;0]�m���v �z��Y8Ɨ�z�s�{v��Mm���\�t��0z�8y��<{;k];�>,��GDm��7��p^eۮ#ɽ�]Q�ٝ�^u���lujzɺݎ��i��ژݰq��i�SSG?3��|�v1�������vݻ)7��*��{�ĺ(s����f��x':۠��[v�w�瓭�!�|�crmm^7����iƣ5�������v���,>#]xM��Ҵ���ܒz����!�8dB�8��-�öz����Œ[��� ��B�]�9-�9�s�yۚ�痂��WR�-0�ܝ��m<^lp�qb�nt�n�.���q��\�{;s����^;���o%g����ې읞p[G#�%չ9�� ��7L	�;�@\8˃KӁ��!���:n���s\�.�-���d���E�c�u�u�c6yy\�И[�X�����	7b^�jw�A��FCv�n.����:uMI$��t�T���1���3�w<�7gx�;�/.�,ȫ�ዎ%�s2�Ul�.#��ce�x�Q�6���C*����r=���یn2��&܂����9�x��{!�/"��񳃰���v��dw�M�.�0�gv@��\��%LJ�TW�����v��۰���a��;�;p��m����=�<�+�Ĺ��m��0m�)�����U1D̪�&
�d��z4��N�\XA��E�yV'��"����Eev���H'��(ج�eF�)�N+<f�Ϩ���
�wF7:���@��{lY$�)�4��]���y\��w�yQ�/2��B(�
Bڒ�%�εo���W� � �o;��p����?��qYjm���i��.X]s1qW�o^.��z���"!�Yjm �O_O�n���ʃ�I9�t=��<���Gn?�2[��B�% ���wk���'�L{��/�8��_Z� �����/�=Ʀ)�4" �@���(
�#;���c�F�
�r)��\�3���wMۧ���~����a%���$N����$9��v&j�5aM���l���U`mW��G
e��eCv���v�H���n�۴'n��#>���}�L7xE]��m'��d��a3�%��8೷����HGx�a��zxz�𸦉3J�uwy`ݏ?[y} >���V�@#�������D�������|��+� �Q*%R$��ŏmZV ��ܖ� �S~��6�ߗ0F�Z��A�s��+͡�!��!mIv�v�<��n�h��>>�Wd@�5�-�=��ٞ��db��\4��;޵V��?���p\���:$�I�uY���{n#���H�j� �G����!$���j�Uה�Ⱛ&0eБB��e�:y6�jz�7X�9��39v�O���'fݪ1���p֢��'͙5��	ޡ_R%|��l @|���o�J���jdј&��$�΍�5�r#U8iS�p�y}ӣw�����Rj������ ��\C�*h[�NW�����0�hE*��wM� '���b�aQo�[�1n]����08���a�y����v�|�̯j�^�(��^��8�����S���!�C1i��/A�yc�;��)[��Ţ�A=αFx��Te�ف4�!״�>5o=�1�H%�nM� ��Zm ����Z���i�w���z�6��ݥ������!mIv���mC ����&��q��V�5\�����"}�i�@�iU��~*&k=�%d:�V�r����$��SāJr';�'c�t���_/kĢ� ��{�;�T���W��GN{%�� ����ն�!x鈟f����ٗ��`�o4�qg-2	r}������U%�Umi��x�՚�7�L�Ng4� ��-U��.���zMDW��o��~Z-!C�+q�"R0�o�w�͠��$:l)���RWϧ�?����i�� �BP	!�{���a�L�n��/��e���e�_z����Q�֪"�G��&b�J�(짧���yZd�`���&k�؍o�[�ó���a<���Q�Py��'�Կd�q���R4��0Ǟ�v w ?f�#����a���iÀ����T�D�;���޾�ݢ��=��[j� �;��i���9e,��#vg�w��]��̅�/F��/r�-��k-�;���j�#lBӭ-�0BT�������mHSR_�s�� �ڜ�V��|6o��S��geآo�>�L��Pxh�[A�,�._�WL�F�J�t¾)��`� z�b�,����?K��z8矪T��֐�KG��>��l��qQ��M��d@�S�w����O }U�Q�W�I�Ϣq��SQ�rK7�N�՘޾>���]�*?EDDGt�� mv���/�O>oTG �&�A$=:�,FBʆ�l�������Wu���Q�ꭸt�QwYi C�^�2 ���Wy�m^C�pW	��}yWOF���O+���+6M����׼50����so�\�����7�e|�1Js��}�ؐ�������v���z~F��B25���#�m�2��;p]�@^-�>��o̝Mk���{kt�k]�;l�Qb¸��\L�G[����ٷr�n�t�j�7R�%�y�%��FX����\2���Yܵf��i}]ϱ-Xס��]q�82n�mس`�u��܊��낻Z�
��o�����6ۋ0�m���훷nv��'�@�4a�zv�D�FnF�LoXꝬ�a���i��]�x���Mֹv�	�:�<���ߟ�r���
����V�� �:o����z���pbi�����w(�H��땋J��>
' ,�TR]����`�	t��7��?n�zr9Y ��� ޽i�Pxv����Ѭ��ڵ-%�94	N˒�{���H$Num
��L����ʽ؎�w�� �������ŋK�V�ir([������~�-yue����o#��A�f�`[��6��b�����z��3i���/]�W���dH�
Id��u����SU
[y�۽ܬ6(�wv[A��l��0�X�ƞ�<r��/��& �P d���ٷm�yF�i��ck�K��aw��8��������s`�"�H��HTg��i0@ ��B���=S&�J,̬�������-@�ͦ������*f�T7�զ�$�L{���V���?W�]Z�,�u)����~7�j��V�"���7>dһ.�{���j�}�]g����F���H�Ʉ�����靄�����o%`�wX� ��Zq9Ȩ�Az{}�3gw��kj�S��bN&��E%����mC �r.��:��O����z��� =��4�G:ȫ@R�e�S����iu�Lr���)Rπ�'w֭�>�뢬��;�j$s���h����v�򋸆�9_MES�*�z/� >}{M����n�v���`�����>��l�v���}}�?2�H�	�ʈ������yۛۀ�;\bz����cL�߻��S<UV� �{n@�*��`�����qTm�e����ћ�W���L�Bk�	���eF�a�`����}},X ����R�붣��n_%�U�ب���4�.�&�+mT(�x�_�kkkޑI(Q3JB�B{[`�A��� z��J��w��u�Ѩ�8���\ZO�Ѿ�Ǔ�Rd��o�a^�;����"SI��<�3��w��k�Y���{.{�`��J��7�X��@(���� Do_U�r�1yPLm	
�K���������a^�$�[��� =��m ���[���;l�d'@輦L�X\)8
jK��/2n��u�e��sVWb��'��ӱV��^M�4;��L+}���G �!�2��FM�#P��
D�[v���kj�pA�Γ6�ئn�g2�����5�QU��,��TZ ��� ��2y^g%��[�e�0�I,~�wi
��\���$��_P�Wa���w�˕T�j��:�m����O��vמ���#�u�S_>�pL�*E*�(l����D�u��� �S:�l�ɞ���> ���2�'w���P��4Zh�iXB�i�����Q������4�d��A����&�HNxf��]��^P��1B�n�6s�~�2��C�9������� ೵�Y�{�<��*3��O$��:�V\~U�5����I*y~wj����ßHSRU����I!5�����}�NG=nɴ��m��$Nxe%+70���=���"Q�*@L,((��[\������6��D��$�LơD�J�M	0`�'��L@M($�s�/�Z`�	��j"Q�0�sξ96�-G��s��v�	�����(��.Tp���!�2, N��C|��}8�@���q�����A�t���u۽��{gX^���15$�%��*��A$���݀�;����{r}Q[��� 	��(�	#:a��I|��e6� `������}=���Ȟ߹N�� ��[�C ��p� �w_U�Ǯ3U�<gs��($e�X��:_�,�HR4���	�iv	Dv�SL�ȗX[� ���7�D
*}�X�k��:l��ߺ��C߻[���3���3y�G�Brq-���~W�����H
a����:�W�Ъ�~�E����ǀ�,�f7�<��Q��JO�@�ݷ$[��m�IY[����k[`<��\#�Ю%ݞ^-�Z���&L��.�vS�ʕ�8�7l�����	��	Eσa�Sכ�1vxT�lô뵙�J�kι����8x��K�w%�]m�wr����F*'��cN^q��9m�c<�%�e���=�����f۲��%��9�e�)׊�9��c�f��Lv��u���v�q\��VÄ��Ƶ�L���[)�G�����=��eϠ��0��ep6�I!⯩�G��m6�~t�Y1�Yd��M2���P	*6M2Rp㖭.�d�a�+�˼ˡ�E���w�b�>����A��Wv��_���_�j�����#0�%;yוRI P붚`���ױ��y�� ��P�i.����8����$@�(�I��	5�ܖa#h^Q1!����H��Ol�$�ٽC�誵��G�K���.]��2�h�IR�	��i���Vo�v�*�z�z�����)A"R^��v�(.��(�AG��9�R>��x�э؋�xL��>���^���sv���
�$�������!�B��#�r�" >��i�����N�ϫ���w�Is6]��>ϔn|�Rj�A��o��+ay@f�����dfP��c���u�ٽ��fq��
��5�f�*�&�
����θ�N�L���ց���w}z9�A��ܗi ;7�Q$�R�U�C���ڄ��h���r9K[����J	dΦ���j�M]<���h��6���PI�z��@>gx"�))1In��+ͮ޾q���I$_e��$��i���(���i���|��`Z�WpFӒ d�l$����)%GiQ�wT�7wҀwSa#�9�� @EOiW�������ϊ"f�ش<���8s=�ns�Ǝ]^r�u��q�Ez:�GW6{ٜSd����'Y�����W�Iv�A-۷����$��J$�^��i}c��e�"(�.����T�{(�w��ˬ����`�@osi�4��Ҭ^Y)�W����X	�b
�_
���û6հY�]��$�ݏ"sȫƧA/,�ܻ���)܋��;�ك����{o�w^�l���j�U�Xo�I蚅%m����x<�����yyh�io�k���
�َ3rS���DF?G����g���z�b������=�M},����tl���U���W�%��&Ak��Omi$�݉���ۚn��^��UC�����7p�ivM��K������xYO��� ��+X|���������\0�G�X��l�p����R]���1����l񄜜���
t{���7(r������)�{Y��vL��`bӮ:��ӓ�'����kU��v�g����^��.��C����զx��1������{j���/
Z���!�_�8^V%��*�!.>��Zg�L��ռ�+\}p�V��&��A�rѸ�Ck�Z���Z�{`�Xe ��w\����S��]Y�{4�}�v��VY��❞ǩ����o���97.��/��y�UY쁨o�ӳ�p���k����H�r���E7��ށ�<��-W��f��x_v�/�8_�э����g���F� ��ފ/-�Y���|o\����5b~��yf�ٵ]��`/�W����UW{�}�|(��Sݚ���x�A��#�o���Od�ux$W��w5��ü�+��+=XչE�
�_l�{~͗�zvJ��Dc#���b�m^j���՗P����u��AS��g�ksoy��5+�z#!H�h�U�F*#��fc��t�|���D�-�#��2%�^XS��w���y��S�d*E��U�AJȱ�F$��F�����ʋ��B�J���YP��R�T�b0�cmV*ƖJ"���m
+hUAEmQ�F
)V�V(�ʁA�JJ��H���H�XUJ�Z���(�X)k	E��2��("EVѶ
��J�,`���-+hJ�6�P�E%eV
4k�,"���)��(PYR�eaQ`)*�,ekR������őjE��EEP���X��*��b��XQ�AB�jV�F2�,k�*��T�,��V�E"(V��J±�*��c-��m���*!-iX���`�,QU�TQJ�FAEX#Q��"��A`��E�,Y%J�"��Z�ʊ[EXJ�TATR-�ֶ��/�~�r��j��%n4����9H��zWu����s�_G���-[ ;�D_���(�ܭ�q�;ʹ�e���IP��p�%;C*x�$A#}[.�uq�n�5���BP��6 ]Yi�Kz�]�A�:"Pkߒ<���R=����N�F�(�x;8\vT�Pv
N�g����;��4�&'��Y�A!2v/�  ;�)��=S����Gv�O�E$&=2�I|�V�4�����'����	�s6�ۏd������� �ɆRH$�[Ւ�%c��u{G���u��kS]Ls1%AD�4�B}[��v�S��@ ��Ys�ގ�')dG�����H������*|�Q�d�{�
������WA��"Cr��ܾ�`OwZ��$ţ�F�X�ll��
��v*��72M"+�܄�NX;+��[����=6O*/�G���>�qH�z�5|T��`���}��tY����$;2�H
�^�L��p*i�6���| Nvۇ����#r��mҚ@ g�mY�ʹ��2�{s����;�2!l�Tr A<�8������n��SJcn-�۠4�[U�������f �2F\��uO��D���v�I ��{y�����eg�̷j�긨�@�n�ҜX�pHӒ d�m*��Ce?fj�M{�Z.�qv 2�i�=�i�@��U���:�=�+�)��"bTԄR�%Kh&��� �u�i y�{55Qޞ���c+�H���Ţ�/��_֐��k̖Ԑ�����;�1:���o��Gk�6J{�b�"R]['��'���׎K��6~���T�BUM���W�#oj՗��y��Gw���'s�l� �ګ	����f�*�ȅ�z��Ry�ڹ�S��y� ۯ)n_%�Ȁ�搙�^����%^�'��z�I2�1*xݧU�>�@ד��7x{�˻p���;��ϲuM��5��ݳ��6�xd�s��1	�V�ư�	�b��;��z�����f��#�gb��c�9}��u���v�i�<��nr�9,r�kCc�n`,�ƦyM��Z��^�g�<��(���gu>ރ�kz��ۢ0�j�ӎg�xH�	�m{�N�ɼtF헇;[�2ᱳm$�!�^ԷD�j�z��͎-��i��q�¾�:�������t�vv�{p�
�;^�	�@3	��,����#�D��ZI$�3�� H{Ua]��]����˯E|�O۶/�H��2⁶d��-��E�FI�C��>�sp�{�m$�A���$�\�c��H�{�&��|+��lϭO8;24�%	T����@ �/j� G-�5V� ��i�PI|���I ��Ñ `���]��~T��ڢ��#PW7n@�Hɾ��I�wD�Ⱥ]�ׄ8>��(��ׁQIJ"�q^̉$�H�܍2��Ǚj��"<�}�6�#�ڛ@J	t�pUa�Ja� �D��$�r�oj�ȓ
���9�p�KuoH/#E��Q�|P�I/�K����H������ 7�����w��[�Q�/���I'���)ą�Q_5
G)X	ug��H$s�jo>�y�2�ܫ�;�5(����}x&�1��c,aJ{��Lk]蠎��@[ŏ->�vm�Og���e����-�~\�����᯷��6�$�UђI=�l�-d'Y!U������b���e�lIN[���ޔH�H��eH���tނ�4[M�G\��;�i����+ّ�$@�,�I��y)zRA$=n��Rוm|�ο�|`6\�	,.��$맂�"@�Q�8�k ����)��Zs՛�7h#�n� �{�)���sO���9R"�>�`ln��:9�.^ޡ���BU!�1�:��i��]����BL7#�`���H
�'pA����@ ���l���V·_f�'�����U�D��],ZA
�xEI�B9$�K�����,���1T��6gh��@|{/)�:��i� ������o���_iE|�)�`+���a�2��[ +���S�f�׫�Bq��N�4�λ]�2��j%���^�1�u%��t��zx?���;�Ve"��R}#�X�6�b}�{�1 [�/Em�������z�'�H�����RG���b��լ�mEN[��O�i�.����p$�G��Q�'�u
`|�=[$��\�y�J3����c�fF���a'W�`��"b�Κ��j:+�G���v>��D�Itδ� Ɬ��eE5>kj����F�7�jŎѷ���=���ٰt[p��rq�uА�q]��%B�(� j<�륋��Wu�AT�l�͗�A�~Q!�4� FV�M�l�?"����pQ�Ϛ8^y��/����IɽB�
����H}�#Y��eN�׾a������rIV��m
��J-z�H�ସ�k�vNF:��� ]�4�%}Mh����P?H�
G-X	Ow����<y�Ay�����OV�hI"zv��2r=,\�̯Y�+/3�<*&��#���P\�74{׽���������'Z�׀��@zcTj�b���wC�|>�O�_�v����"&�p�S�,/:~u�H$I�=����=j"9l�t��4�D
�+d��>�ڢs`F_�vpI$A#QD\�'8{J����s�i���Iܖ5��&ԛ��.������#Q�
s_|��ڰm��Eϝ4�@$�N�d��=�s�z;Ք(�xG�Z����i(d�Gw�N�jᇶ�/�cٜ{�{} (��"- �N�D�K�|ǲ�!��8ˏ�/�K�	�q��m�w�W��H$znƓ��}ϯo�����>�u�_� ���&�J>���S5UM�v�׼�;����� zzmI| �6�6H�]gv��Y]��"�X�ST���#��!p��/ҍ�Ne��{�[�u��;Y%� u쫈�i��4�k��EO&������-Q>����O�q"S誫�L���RA�w<�������?~"W~���!�,;a��w�߄z�7������{�������^�vnd���/a/h*!C�k�7SK��H�u�c���w�?��C��x�����F8��=�эSۉ��C���v:g6{\lv�p%<�v)�9}����&�v���۲�δ�t����e�4Ywo1e�n2��Ձ��Kv����[���8����;���1�Ѻ�D	1�L�ݦ���j�]:�ۡ;;] ݞ9&�L:�vh|ű�m��ܛ�u�)m��s�<=[v(�-�2w�����
'e9�_���A"K��v�H�쮱d��{�F7��OM�&%A$�D�e6m�F)j*���N�K}m(i'ճ�`��_���ޮ�/�Ҭ$|6��2 ���j�R�n�AS4�J��Q�1���H���)�AQ�N�m�g#njry��а"_��́ ���>k��PIB��[��[|���/�vw��D���Z$�2��l���k����ҀH3ݔ�`�o#�>���S3UM���9Mꯚ����Rnu��6��e�D���O��u\p�V#�z������>�n��u�n����ݨ=�����vL<���(���P�d,�~Q�Ē$.#��|����u�Au�pX^�yu�N����m�����L� Ow4�`�����AD�l�.��#��N�K����v�����{�X��ˣ��+�HWWӯ	�%������Yy�W��)�+1aX��˸�j"��5Y�X���I/�Is�>��� �N��V�H���&�V�}==i�N���T �t����P�\���A ��T��ǽSռ@��4� ]7]%��(��U�J�T��뺃޸��ˠ�������8��- A=�D;���N�6�[P�EA1B*6�,�|���I$_n˴�n�����,�֛��� �w��e���U��0�$�a�"#S���T����6����-�nM�/hr;h
�-�w󿿟O�v�xL�VD=̾Pπ
ɝ.@ ���	Z��ĩ
DxʗC-T���5�h,,�A7��D���}i%Yfl��6��È �����D;�M2 �r���������F}i�����E"��i�eL��A /���:����]c�Py��-����͊Kݻ�^H��zٓV�7�����,��%���eE���Y��F�x"W�Y��Χ�m��Yǅ>��޿/��o�k�Uh$�~�F�S'E�D�(�N\&T�1;ƱNe�E��.AA�>Φ�sy�J^9j0v�_�/uW��鈡�O�%�ϭ �	=�7Aﻻ&��%�'$I4}�,Z$��zŁkq����(�R:LNQ��عz�̹�=��m'��� .�q�ۮuGm�,�~��Ӌ�-��Q���^�ʚA%�E��l No4�A�W�Q�V�uof޵Ω��;��M�
 ��7$�}����J�V�r�1���/|�� ��e8�=�i�A�G����ª��D��X+�"�1�j�K�~��� 9�nA�?p��P�[�� @��X�%����w�����i��_.�"�ٕAQ{��4 ��i� 
����<Spw��<��g�j��G���e	��+���\�^:���2t��Gu�S�{�t+p��9�	�-�/lG��#�sN��������;��$ 7�����k����/�4.�iհM; ��� �+�������r�~�����y*�D��vػD���5*�!�8��|	��J��C-���Xj,�g��	�ٗ�U��d�r�W���w��߿�OH$�Q�*{gI%��>��	
��^��<��u{ ��S�� >�i���z*	�2UCc�.A���1� 	eo4�D�Z�Aꪘ���m��{����d�#rK����I�7�� �+7�/;�i�v4 GWu�� �jT��0��%�[����v_�����s��A<�j� e�hDDZF�k"}���7c�ڷi��J��QER��i���T��]��q�]��^��i�?���- NۻL|�F8�ke �N����IP=s{,�_��oC��JDՅፁ�{̆�~喰��6�S�0�؂)�G�:U��;R��{�_�|v�No ��q	�|��62xz_hG��t�_�Ol-�%���bm�k���ܐ�{�;��Ԣ�a&ד���'�>b�^ڱ�K��/jFG�EF���	�Ӈ^FYX�N�MZ�Yϧ!��̢1�z�t��	���5x�9r�@�C]�wjE�{������G\����x�#�
�S$��M�y���u��^��${黧��b�Df�Um�$>��Ĩ]��x��{$��}z��`��5�9��ۛ����i'�ݹ�J��'�;ҍ�_I��	�ɑ"�^{����9�|�]����kq��Pp���c^�}��@[���d K�-��&�)��}vi�n51���]�q�^�ł�<��f$�+�C��g�>��-����|��#�;��X�g��h���h��p�}�E�g�sR��,��K���xK���`�<;��Ho��<���Ū,�P�;��ɋsM�:�w��x4V���M+�>�}�k���vP�ώЛ�x\��f�-�{A=׵E��M���M��n<k��Y^��a�и0�a�v��������L�+~�J�үV�׃v��ǔk&rMB�b�el�Wr����Mn�W
�z�G76x�G�'� �~K�4j�J�Ŀy��n��j��Mq���P�E���������Q��C�LQ�d�7��=�������aܲ�3�B6u�r��H���U�0X��R)��g� �X���eI(�Xŀ��P��b��Y%`U[J�Ņ�""ED(�"ł�@���
�V1�
Qkd��#"�%V[jAE��D�ʕ�(��1k
�1���+F�P�*�U"�*�"�(�)+
��(�P!RV�*�A��`*��YP�(,YR�-
5��
ł�`,m�,AAb�V �m+"�a*�`��1�դ���)h�TX�J(�FJ���YPDX[d"*��#X�T$P��V(��ŀ�b
��9onbf�m�mm1�$���1�n�p1�<�6��9��%Q�����4ums]��7��Odܜ��!���Q�����8��m�HR6-�k=W=�I��lzx��nN���s����;q�������!������g�n3Sֻ!��|'+��Z�v�TA�g<e1��wdL����p�ݴ�t[I�[C$Y��#5�m\�mZ�'��i^�y�Y�ƪ
p�ק�8�m�\�۹��l�; ;��zۘ��P���r��6e�1���S]X��sۗ��6��ǀ�^����ڎ��rz7e��60=rQn5��g�cc۬���܎�n0��Տt�M��Z�n,d�q��j�ЊOcw9�ź��y��*�W=0p�i��As�OT>Zg��O�����f����ՌΎx�5�wd\Wu�W����n��OcCv�q��������r���v�݌O��X��9^7�kZwg�=�f�/R�q�8�ۭ84�X]�!��.� �����8�pn.^����R�yǱ�D�t n8n�F�'V���̊ڀ�1�WTD�xz������;���k�,���h,�7]p�e�[m�x�uϭ�i�G&�!g{1*�أu���$�s�x�R�oF���3u���j��Z�n�n�,p9'Sv�(�(#��:���e��{1��q�܀��=c���e�ۛol����]wr�Y�u�O��F87�i�����R�k��1q�=�nF��ڐ݋���rs��i�Ƀc�s���Z�:Ӗ4�h��;�5k�S�XK\�uZ�nj;<[��t�P���9��X�:$rs�ce+b@�w]\Ǩ�^<۪]��n;[fAᮣ�r�t�����sn��2a�gjźs3^�lX:y<�a��e燆��l�XhD-���=��n�=���0<��[ɥ�϶n3$r�[���\v�M�[9�v:��ֺnSH��g��s��m�[��T�jŖú[���%e�c:��$��D�i�8��6��g�����������{O/Bk@�#:�uf{y;rp�g]l��y4��ݣgpBGj�����m��ح����8��Gr�ܝ��l�=g(90��n��v��n;'��Y8�8Ӻ���,g؝�97V��ms�����N}��õD�Ӷ7<=�u�n�/�fbк��W�����Sۢ��������ϖ�����n'{5ф�[
V�jx;\Nnۋ9 �]q�
oQ�����T����1���W��dG
p�3�������Ne��[��v.@ :�[h=��/_����&�}��&�i��^.�&Зý�h��wi�m�$�~&���`�S�6 ]���u���D���z2��^16cID�T8�/LT ��r� r;:c��-G��&��@ mv��V�g~�$���U��fu_��a���'@�2a1`�Wsm�Wk[k�WP�]�yM	U�W�)��ϑ-�(�i���~m���{m(~����3�Fo�G���A�[�� �֚b3=0��5.������؊&���d"���E���_`��ۮj���z�����6����� QH)͜�}�B�	 ��ڻD���i��>YW�{ϫz-EͲ�/�W��u��)UD�������0"7�r�������P����u���ݛ�r��	���:XZ���2�XzN����>���t���[������s�ݾ��b�kn]��4��.�I$$����>�>�_�7����֛""�Ř�O��N���[�����n6�&��L�>��j k�0�׏8��� ��m� >;�Zi��Vb��҉�ZsH;zש�*���m��e�` "z�*�W�ԣ�~I�ޫ�B��߉�|P��.�]Y�f�H����ZUl�}Ay�;���ۈ�h�^�� =[aX�qn|�o�~�~V�P���aM�\����{. y�$���+�W�ѺUf���w����ߏӵ�f�I5��v?6� g^ۆ �c�bl�b���(�O{��#r������(����Ƨ�4��+�:�^^�ͻ��@,������_ ���"�2��K�b9��U"4��[Pς"`�.�_,���_4��O�NS��n�����������y��3��O�����/Hiy�c��xΚ�f�\����W�y��"~��ж���G�O>�|�K亹�~�@��ߚi�$��l���ҩ�����n;�S��
>>�l���K�=j� ���l=��|�ݖNyزM 렠`W
��4e��-*�"{*��Ɠ��]x�\���
L����kl�/{����;��]Xv\�����4��u�A�rt��u�ڰ��ŏi��$��$�_���f�_������kl2і��~1�v.�A$�N.�J���b
�������7�w7r��뿻$"Kkx�>���m�`	=]`N�]�D^m⌔���w��i}�]C)e9r׍ע���l @^?u����m{> 	ɭ�� "{���u�F�D�h ��i�U_�mT,����@%\��� 	����|=�k�E�S~p�d�S�bj�W�L������l�蒸�J�0`���rz��<Y�x흭�ҎbQS�}��UU������%x�≯�%������n;h����0>	��o�a���&�ޭW]y��5�/�> ��w�D����k�*{��]b(�&G	#i�Ci';����^��lk�F���'i.�.iw}����;�W:��E�v9)	��l wy�Яk���l�8mAx�A"Rw�6�:�$�$�K���vP��*�o�gEK~��v�G�> ��h"wy�&����]h��ue�e���A@CpDLӦ���� s:տ�5��]z�72N��y �6�����{z��k��:a0�)ʇ�;)�n^{";��B+�>���0}�j��9�)�z�v�vQ>W��v��2z��AA�եR��a)�鯚u3,i'Ԁ�6���}��L�
魂������~�z6f1�傇�(G�3F�98�>x��~)�ݾ^�#[f�>o�ժ��_j�ݧ]�sFw�y�{�vcE����vT�&��dp6M�	۫�.g���w9�C���]�k�9n�y2��ON��0��m�=u��m7a;����.H���v���ݢw,9�]���:�b�l�7�l�Z�9WN��d����X�5��<��62������]��W���Ã1bt�o3�k�6�V;K�m��z��D��f��;M����\G[q��ܻ��nS]��)9m�b}-;��0��u��l=�nم�.1��[ff?���O۵�U(�3S�����`�=�j��W9�P	{�wM�}�"�]o֊I �fأt���'��Ew�SM�J�9{�#�C�˸� ��6�+��, ���a���
���U_@�I%���V�i$���������1�N�#���W�t��h5�hE�J����~�
�Rb���	�޷�8���Y��6��x�Y
3}fÔ<g� �slQ��`�D��r��z��\� w]�dx����-���i��
٬��D	]ͦ��^�]�y��?;`��B[Q�1��LF66]�6�۳�������v��M9&�����~��8�ko�At������'bԇ��}v�]s�,z���bŢJ�s�Q47���`NBPP7��Ղ�H�C&�����,=;���ik��C],#2��$#���%��{N�˻O�wŏ���M#g�z�^���<�P锋��m������;��� >���� G��Ͳ���9��Sqt����i��^x8C�$QY��IĻk*�  �5�f9D�dZ�y磽J��t��h�|�`�L7�D�(�UUT��=�Y�
�ϓ�y� ���
����I'�\nN�.?B�_Ts
�� �*d��U:g^y���NesHu�,�U�^vo�-�ӂ�Y��v��"�g4�sOO:=��Az���u�����+��9-���]�a�͸����i���&a���H�j@QRzr�Sƾi �y{m� ���]�W:u=~YZ���� �����]}*$B&���m�4�['���^�髝%�)���m� ��踆w�N��W�y��Y^I�7pp�Զ��ͦ ���1 ��c�z�ݙYt�ڇ�z[�Ǵ���y1��f��ۊrAp�\Ǭ�ܬjK�}v�??,v������w�%���V�A�$��,��L��jяo������O��V������0_57�G�(UJ��(�®SN�z\;�F�u�&���̈�2����
�k`\W�35߫ɤ���7�m{D0�Al��w:{B�PJjzh5Y�ײ>�B40��$�vv6������" ��k��d�噳�Z(_�p(�P��1�#-B�B�ך㜉�b،m��y��d�I@�"B�o%,�3T�7m����eesC> 
鮂"'����}|�g���� �VWCL>�7�G"%�EIrע�(�K|T;����� [[� *鮂��������X�9��Q����!N�	�\�$
�z.C�N(]���OzOe��z�� �
鮂�C�%���%qݪ��R��;zŹ�ؿMh=t��� ��dM� {�x���Y�+:�t`iu��x.���~I�r�<}s��u�m�Ո���ǜ������<:�;a�u���d�~ٛ���=�/���?�	%Uu�صaW ��bA�(�£��I<���m_z���:�[z�L�R��p���Y8�I��ڻLpǙX=����W��1�uĳ��û	;q�F(鶎��b݆��K����AQ�p�F}�sC���R�	vmc�
���� >��n#�����vr�jԯV��I�_%��ץ6M@K���W{��<�	v��ޙn'ý�=����VD��|;ۯ�!%�]�ߨ�uG�ZX5�(�� (�.Z�Ś	�۷��I �ѓv��q��	���f�A$�}۷g�r�<�AP�A9u$�罒Ԯ�Gg�;�=���� '���yDu�3�6��Ί��y%�G<U��Cw�6 D��vfN��$�WK�����p�[�1l���≤��οy@._�t�	������0��̏w-�����%�eS���8�@����5���=Gw*�'�����2�ⶒ����W�K�~�}���f~���B&aٳb�Z�����x]����&d(�Ճ�c9�;n��Nb���X0�gNw`�9�^9��%Ә2h���r��тCy�h�zO`��������ø45�����O	'#Gn�s�.����+�k.�ۛ��{3['�9�,����qve��tΔ�NQwhw��s�q��o\F��U:�b��O]ۍ�k7&;`ޮ�y�t��aѴpN�����^���Xj�ך�ݒX���o�ېH 2E~
�N5�I$��ο$'�����nh�o�7��, �Y���>n/�ʡTT����Տ�3}����W��; ���۲I�]]Vh�.I��|���=��hIVN��Qj\�-Ow��I�����	��<��JҮ�ރ� �;;��Ȓ�]]Vh���'h�
)˖��'�F�19U�ҢI+��_�� >Y}n@]U�0�ې{�	+P��=��K�X��T2N]XDۯ?� WL�r_����Ocu����~�"�m�L�]U��ʯGz��v{*.e<���q��0CA$�Gvlא���D�{@θ�@���ӝ];���~�v�	q��S|c��{�@}M�HuV���u���������@�G^ۆ��Mh�p� 2Eڮ��|�K�k��"�N��Z�|s�L��;���^86dK/�%}|�]������t7��[h7� �����Ɵk��[�����_|�O6��~@��� W���W��ݜ�� �����;\EB�AU$��s�"�+ft� ��!Mrr����<u�8i� uV�a�F3'������r�u�C��%"g�~��9��:�vm怏�����+*k�w��Y�:�f2VV��}��8�1���`e=����?ky��_}����d�,�LeN}�~��N�bg����3%�QN_��Q,�6�eE�c&32Ɍ�,��o�}�Y:ʴ|��{��s�K�>��xϓ�1�������N��fD1��N}��ٌ�9��23�d��������<f0��>9��}���)�h��uj:�E��n+i�cvv����y*9�N�f{��*��'8i����q���w�a��L�f2VV��{�8i������ɉ�������p��#/���t�������~��o��Y�J��$�c�s����f'�O|����s3F.���4�2T����������@g�@��Z��>�n��?Q�k�<f3�c1��YXa�7��1���3dq�ɆS�������r�d�_u/+�_ؼ������_���:s�����֍���c'S�0����18��Y1��LO��������c�1��03�!��w���󟪢���YY���x���9�"���Y淦���8U���H�2.S�ρ�nG��wB�l.�r���.�)�#9U$�xc��	����N���TJ}��s�!�+���|��Q���y�`�,	a,��[����G����ǝ�7���,����V���'�nw�^������|4b����*�1�ua;�R�YzCjy^��c4����9��m�l�q^ƻm�DzD� �H����D�0ѝ��������j��|({�5f�e0����N��k�;��9���= �^������H�8::��Č���m-�nK^��6{V�8+�70n���UB*�;�r�sF�\�Ҏ�!i��7���V�HV{��3i��DG@�/�r��~����Ƹ��E�h8�Lk��۞�����J�����S�g���w.R�wܵ6�-t��ö��gD����[0���<=
 �,�&?p���^��M��5кz�-�s�Ym�ɱy�8��b��z��^��o2�f�;.����'ҷq1��,�<ʄC����㾒�/g#:��q�{��~��}�< ά�����^|�����HN��|u�}�k����c_LJzQ`�t��1��s�w��ߞ�>��Lg��wa�������9������OP/�m��g3�+{=��Ӎh6]�͍{,����#]�Ť��N�4�ߴ�RD���j��#��n�s�Խ�'�HT|s�j�}���'�1�{s�?*N�%,X�U��"!�E��(,X-����A`)�X�(���,PU���A`*��* �F*��1QTQAEE
�X��"�+dR(�TX�����������T*�,�,���(�����UE���f ,P1*)�H�����"�$Q� �Y2�9`QPA`�.P�D��PQJ��P1
�Z�
��"��Z�"DAV
e�"EV
��Q%jV�.%`*�QE1*��H�E�����ũF�X�Ym��*""�DH��b����*
)1�`�����{���³��c1�����߻1��c1��b�O���񓬬<�ݽ��bJC��#�~d~�մ{�<u�{��u{��~g̜2�d̳w�kݙ�4ɎD�LpLd������<d�<q��LeO����V{�����o�x��$�c�����f'�L�8�~�s1��u�C��u�&��Ϸ�'YY�!��0f3�{���C|Ϸ�|���:�i��w�߼1���3c��J�o��Y<<�.Y���LO��;�W���̏�C�t�G
�⻛a�m�܆9�ΐ}q˺z�[��\qܭ7[q�l�� (��Y�V��(*2�s���?~�L����Y�,���S������I�1�&3�L��;�Vu;c1�=�u�5|��߃��[��ٌ�Jʇ#1��S�������Vy����X�R�5ì�N��Mw��a��J�����3ڽ���u��p�L���Ɏ&2b}�>�}d�x8ɉ�2c3)���w
��Ɍ�$�c�'~/�����3+*x{��3�h˚1u��CL�ta��y�����Vx�3�c1>���γ�0f3++{�{�so9��=���~�ƙ�88�I���J����Y:��YY+�b}�y�³��8o������kW[�N'��k��f�{��ݷX����2x��&32ɉ��{�}|x�q&3c1?{��p��u�3��3��k��f��k�ӟf����_�=-M^9q�yz�x����o,�7c�̉)�P,��O�yc�dY�N����"X�x�{˭w��x��$��8�P���b�O���������4�zg����N���:���������tq�dɖc&L�_{�vo��2c�{��6��߻��'���>7��>猞'�����&3	���y�³�l�����g�߻6�dG�Au˔����;��&�����B�9��8�F�3��i��q]s�Gx,Qf��t���ߦg��1��u����d����w�|���J��YS�{����gP�c1�&3_��vm����ě��/�.{���[����c&�S�y�w�'YY/�c&8&߽~��>x��!�gWz$�l��)��&�X\����y2c+%c���_7�z�O������'��Jʘ0�bg����+:�a��J����{�l�Jʇ#1������>3���ٴ�{��d�+'��m��ź���gv8�Mw��a��L�1����;��i��^D�LpLd��s\׾��r��������q�Y+3)���w
���1�Ę�r!���vi��YS���3�u�3F�Yu�i�d��7��4k��~ֻ��+%ed������>f3�c1���0�]��4�d��8�1�����w�My�y���ݛd����b}����^��LL:s��-sWZ4��\�:�a���vi��Y̲c�k�_��x�a���+�<K���_�ʞF�L������u�3��fD�]��4�C��c%ed��������a���������Q�ߓ�ѣ^��V8y�N����}�]����E��.x{�Yꬡ�z�y�u
���Uc�����  ���j!(� ��Q.,�2v����`��v�829�1���^��k�j���C��:�F�M��=])�\�s�R�7��l�cN�m���\f
|�j:�㍞��L\pӶѹ�ǫ��9�CJ7d�y4�c�� N.�]q�y��`�V+yq���r��˝E�{7wGBz�q���^K���G7Cn�)ۨu���ݜ�7%u�䴾U5��zf�'�^��N�n����8j��.8��{���G�����N���L�O�8�O������J��YX_{�vo��L��c&8�ɉ������VJ��3}�{�ߚd�e;��p��l�����!����6�Nf&g����х�tV�\�Y��a��>�����̈c1�����׾����˟O��׽߻>�1�Cc1�	��g���6�I��bLq�əO�����O<�.K1�{�{�x^�'��<�+�N�by_���R����M����]ٶc%g�d�a�LO��﯂O�$�c%eL?z^�kϪ�y�Vx�a��b�a|�ٶbf3�f3��O�����	�1�y��_cn�!9c��#�|Y��=�� ��jzV��3��VM�f2a�c�u����2c�c&8�ɉ������OY*x2c*}�w�³�{����o���OYY++�3��У�"��3�#2c~�S�"���q:������!�1��3���O�����1�C�Mw7�}����hϧ��"c1�f�ߜ6�I��1���fS���������p�1����s��g*g���S�sU�_���%�	�"Y"P�sLv�/:��<x���gv"�y�����������b�5s�2q>a�~��4�tɌ��&32ɉ�~�}|�<f9��d����>�y
βVV}铽���ݺ|̬�w_��f��q��Cc1bw{��a��c�v���V�[�:��L�%eO�}�6�βVVK	�~��{�������g?:���+�8�2(�Vg���?݁L�f>��pJ=ì�'^z���5u�^���s��}����?���_�d�VJ�c&&O��������Led���ϻ�q��\c1�����\M%~������#�"���S4ar���!�m�����o����1���b{�{��:βVV��=Ӷ[�ww���~d}ş�2��əO��߷�'�Y��1�S�}�C�S���W��:[��ƹ��6���ֻ�H���>��q��뙛��C�ZB�������
��R
P���8�@������څC����~�^���������b��~��x�3g�i�~��k��5ì�N��Ms�h:=gY0�1�&Y�7�k��Y�L}�=�.aҲx��S�����x��x�&&��ʟ��u3��&2�VVϵ��3�fu��߭ҟ�ZS쯈%�H�LA�!����n$��0^�{f��ṇ��ѫvbc�������֭�\����?2T�����!�1�D1��3��>��3�0Lf0�z�~��1'f$��u��;����Ι�������ٔ���{�<��d�f2c�LOy�u�N�b`t�}�֮�b�5s�d�v8Ú�_l�p2c02Ɍ�����u]o<�~����\����O���0a���ϻ�q�N�1��C�7�kݚf!�f3�c1��m�q��ϴ��?a���{ߚrD�	kN9�L�N�3��~�u�:əf2fY�7����ri������S��m�����&����_��2�C��֙���U�`�Z��6,�;8�k�{?eV����8*�{37�C����M�m�Q^n�ֺw5� I�<���̞�󌘘�&3����w�;d�W"Lf8����vi��YS��w�Mh�r��kp�8�����>ߌ�����浚z<g�C�df3�;�6tY�0f3`��a�������8�1���`e>����<�y�y�K���^�ߟ��d�c&8&'?s����&&y��~��-�5��:ɴ�a淯6i8�1�e��Y1>��}�_x�w�^s��1��N3�%eO���q:���1��M���ٌ�Jʇ��1����}ߌ<�c���:�l����l����'�{w6�cce�n�\�e�i�$��M�v�B 䅨�}���� �����$�8�Ms��a��u�2�d̳o�kݙ��2c�1�12{��{�<O13��������Y+<�~�{�,�l���Y\C�kl��Jʜ>���j�֑�]rgS�O��=ߌ�C�c2!��)�~ߞ�_'��k����+:�YX`��a��^��N8�I�3*}��{��u����W_��3��w;�߼��}�7�p_����t�~�[u����Y�2u:0��l��l��2Ɍ�,�����﯉<f8����3�a�K����y�:��1���c0Ng���Y�Jʇ��0f'����񓬬4�֤�i��p2�C�����̏߻n�;v�����d̳2f0��_�Vi��1�Ld�Ϸ��s�O�1���?"?~�]|	�n�ߡ�����ݏ�w�kE���������we���E���yw�(��=�w�ᛊ,�o���������v_��$��'�W�$�2�}[A���~Dw��`QAj2��8�'��~}��~3�C�c0C��������?x�e�΢g3�g�~l�����}�8Vi'f$��c&L��������c%�1�LO��{�/D��̌�ߦ&���u��>�M@�f�u�����0��x�K�t;�]�\��c�?7�/�i3H�?a��#�gካ(",2c3,���S��~�}d�+�Lf&0�bd>��� ��ц3�����ׅ�_��~K�w�ef��1���b3���񓬬<��~��C�(�5ì�N�����l:gY++#w�����2߳[�����u�e�g1�1�Ld��7���'�㌘��Y�O��{�,�%ed��~7���p/��{+6���bg������*)~���F�{��� x�fc1f3��l�+:��cLf0�����g���<󾕛I�Ę�1�2�o��o�O'�c%�1������&'Nw��Z�ы�5��N'\`������w}����9�y�'��Led��y߷�Ğ3+*cf&~߽� ��������%���ef��Ƿ�:�>nvx�!��f!�17����a�x�a��z_�k2�KsF9�L�N�3��~�ãY�J�əf0}�l��%\�����/7|ߧ�8�	���s��猞'�2c+%eOw�y�,�%ed��b�oݕ�Nf'��s��<����[��g^j�V#�ـ�ɦ|�r�{sÚy��)������[�1�m'��SQ�8�k�^��ڸ|��o�ť�PĪ�*�ۘ����|>���|��,�d*l���dq���8n3�®����z�û�r�$wc+����5��l�#�iq˓�f��={
F6���u���q�Sr��:��mۈ��H���˸ܼὶ��E�l�4<؃�ٹ���ۆ���;,es�^J��\\�]���δZU�q�;����M7h�m���q���6�՞�k{L�'�qʂ�n��ͦ������պ�u��;'�H[;����3�c��4w������֗2��k�g*k�}�}g�3�c1f3���l��βVVJ��'���³I88�I����˼�ۤ�r���d�Oy�����,�J��\����ޯ�>x��!���]�)��M9~d�u��o͕8��,���ם9��y�O��~�Y:��I����3w�{�,�u�3�f3�9�vVi�������?�v�O�[Jo�G�v��H��?�Z\_�14A�~�'\f&��9�,�'L�3,�^k헒Ͳc+%p1?k��ܿ}�|�y��N��2b`�&32����pY��1�ȓ�!�s~��q�3�<�tֳ4R�������#��#��:��������?{u�C�8�YP�1����9����d��2&3y|�핚d��8�1�2������G~��{�^j���c%ed����g��O�~��v}�D�p�`��2u���z�eO��&32ɌɖLO���w�Ğ3�;���������"Χ��L9��� ����d����<��+4�YP��f!���~�~0�O�=�����~���%qH���$��is��'9�lô�k(;mʍ�w������Anh��4�̕�<����|�u�2�d�,��5�e�d�VJ�c&&}��{�<ed����~��w�?,����w��Ν�c+�1�����Y��f�K�Q		mFBRW���G�?Eg�ۿ:��YP�~���u�����p������>����mE�1.�w����T��b>��]�bJ:�-�tw��T�SE����;N�^�W��J��j��;����1�N{������d��0Lf0���o��f�r8�I��c&O���������rY�������[�O�����N�by_[��:i��n\��ɤ�5}ߛ*q�&3&Y1���������I�1�&3�K�]㝾k��w_���2VVz�3}|׻+4� �f2VT0f'�����<f0Ͽ.���u�s	�|�}�J�f�	�{��1�}ٖc&f0����^m��Lq1�!����<d�<q�#���2���{�,��<|�{�s�1��$�c�g��~�X��̇��~9n0TR��d���߷�N���C�df3߹�l��Ρ���J��?	���}�xVi'f$��c%M{��o��O,�K��Ɍ���w���N�b~��~�޼�߽���4F|�De@B���DwM�hȜ𝣱/\�yT6��]���q�������~o��M�ѭg���>a����Y�J�L�c2e�_�����I�1�&3+*g���u�������u��|�����=�핚d��q��Cbk���~0�<c?
y��8�h���d}��̏߻y�,�'I�c&���ӧ�����L������;}�6_6Ɍ����LL5��}猞'�q�Y+3)���w��K#�~g}V*��r�)�����3�#�_b�8.2��~�<~���~ߌ�C�c1f!�1�����gFVu��cLf0�|���<�B��0�{0�������b�	��_cξ=S}�Sw��}��|<9n�Z�E����d=ڳ�c�x�rk���B_5��Vi'�Ę�1�&S^���~2y<�.c&2����7��LL���x}�M2깗5βi:�_��ʞk���1�~�c'Y+92ɉ���}|"O�	1�����߹��:�c1�c1�'�����Hv��s��\�nm����C��f!�1=���o�x�a�����n]j��L�p�8���bk���2w,�L�1�׺�e�d��:��>}�}�Y4�1�5���<d�<d��1�>���ೌ��������~�Y�3�"�g�ƶ��u��l[�4� �=�fLX�p�pu�m-k�S�g�FT1���̸�8�qO�~�?�N~�o�x���J��YS��n8�Y����a���Y��f$���￿o��s~�_}�m���sϷ�O��c%�1�S���7�d����籺ְ֫�Z�c'S�0����T�tɌ�������e�Wo�8���{��u��&3c12}���Y����Ȇ3��u��Vb��Jʃ���s�7^~�k^o�߸��������~3�i�6�)8�i�I��b{�����Y�L�Y��e����l�,�&9�Lq1��}���=��N�W߇�A���a���|p�߻��;;d�Wc1ȇ����Y���9��^���9�L��!�q:1<��}�����zi���<C�df3���l�+:�YXbc1�}�o���YRpf2T׿{��ɛ�]�s��Yߤ2oޠ#�0z��֞>����Q���z������Y�.vC���sQ��Bn[�ǲ�g��/��ն�+��.�g�?�����Ɏ	��>����'Y12_ǯ��V�hˎk�d�ta�پ���&3�c+%M~�������wk�}�����?&�c12~ߟw�Y��f3�c2'����Y�q��C��1����}ߌ<��.����_K������l��.�N��'	h�7a[S�9�{��u���a.�8����o����r��ğ3]��l;βa�c&e���s^켖i�����c&&���w�}�3���2U���6���o�3�?|�����;�,��&2�c1�=��ef3�~DW�e� Q��W���?G�_���<���b{�}���n˯'Y��}�=Y�0f3bc1�N{���Y���'f2a��{��d�+%ed��?��}�ӿ�����y�/D�&%x{�c��GL����Y�W:��tɌ���e�������$��YS�K�׼n������y��,����c0C�Ȝ�[�����f!��b3�����1���o�N�-re~�>�g�G�ݷ@r���^ps(�2VVL�1�;��e�d�VJ��S����x��x2c+%fS���?sZ�G������`��!��oݕ��c10��^���Mk)�Z�:�'A�&��Ϸ�<C�c0�c%eO}�y�,�	����}��q��c1�Ow���f$�ęf2T��~�}d�<�++%q1>����N�bY�/=3�]~�>�?�����r��)L�ule�E�3�7�Z�X�㱏{�>A��6{-;��������W��v��;|�fG�i���sC�/Q��ڹ��㥝�=$TN顜�w^b�Vz�cܢ\����_e�����^ۖz��̨�ga�z䠵龳ؽ%rW�� ��y�~��T
��=�h��gT2�&ɱ���*ڬ8B��Z5Yt��zlz�9�Q<j΃����T2���F{׈�=�>�j��C�}����Q�Ǒ�aU^�O��˩b��-F��to��{�S��sT�ힼ+%���6������Hu�s����kN�S�8�4 �g�e3A��x�ϱ��7Ho{)Wgǯ*�,=U��}�Ӿ۲��!q=4�+<��j�c����)�nEn��C���,X�u��Br����>���4cp���{�z�(Y������r�d�yv�$.�tw��6�o�܆MD4C�i�ޤC^���C1b�b���F=ۄY稄�W��������vr�sױ���p���lU�������{�W���{���]b��
=�w���z�xD�zRО2���轝��<�.�a�7�)%?{�)�e[�w}E�Q��+5Y�X���cŁ��ʹ����g���,����<�wsƽ�4�yc^������hF篡 ���o)��|�| ;�xm�G�����L��5��f��Azg���l��.I3�`�o����D�=8c���n�
�J!�  d��b�"��Ŋ�DQH1UDV2�8�IP1��J�EFH�"�$��bȢ�T�UH�ɘ�`��(��E�UX��J��T�S��V�c&$�J�*��5H,�L�̈��*�Af1��Ո*��Z5�*�DYAedEA`�PUPX"�EQX�Ĳ#"��T@Qb�ȫ1��m�%d��dD�AU�Q(U��R��1�
1�E�EZUf!X(�QTUUH��q+U����%��V"��X"�c+&$U"�EE��X����U@��E�����AeJ����PUb�"�lH��X��j��H�UTQb��Qb�$U"�B�H*��2�&0�DV(b�
ȱf5� �*5,ATb
)�[�� ��#@�PZ �!����-�oQ��y�:ƶ	`�����n7+��]n*wkz�o���=h �{�f���v�S�yy�x���҂n��Q�۬6�z�m��D8}��73��m�%�%�:��f��]ΰ����]��wNi�y�c��#�6�T.ۦ<���^�t^���nƈ�t;��iն�N]�Qqg��v��v1Ji�(nC�u�z����FP 09��C�Q�\�x�g۬y܊q�����\�K�����\�`��#���=��a�U�g�v봽�>��v(�M�|�=k�)\���d�&+��������m��M�㞱�ZM$=�u9v�#ɻv�C��v�����͌�걍���s�\�����E�`�<���ggv6���N,q+��G�;��m\�cM�ئ�*��:�/Yj�.܁��7���x� ��^?��m|�{ �L�Ngc�u�m�Gg\���'crT2�3۷�n=�vۇI���J	Fg��wnvy;;�������W��.닶�t.`�.U�6�m��cEky����[Y:���L$��ckθ�� ���v�9�gdSBc���Y��k�|[p��lݝ�e1�s��c]8�Z��q�{�:��Ş�;��\���u�Zִx|�nSYT��׮쥣x\���n�xNy��u�O@�ؒ�Z���m���[wh.n#=�۫\�*�W\��n<��Y�.,�"��mֺ�[���cQv�v;q��L�7����,�/	��sI��׭�f��k+�g�;uk�#�δ&R�чpJ�&7V6�:��
	�Z�{s�=e���]�+�˲F�Q�fr����<�qt��`��g�8�v&�c�"�:{aq���sFs��;>��^8�^�q׊\槫�b�n{�Зn��ʒ��ܲ����)������km�cLj��N.�*簇Bgt�"X8�h��ݺ��i��ms�A<��9���67n4y�Ci��p��s�7gT5���ۅumӢ��A��m.T��7=v�7���s��;�x��ͼ6��f�N�vt>����ؒ�ۭ'f�mѰ]�d8㉎�Z��^�y+j7��w.y1�����y�k�;��b�n<]f�ml�x��9M֌�;'m��H�6n����H�u�F���M��L�0��.�7�;8gXZ��u�0���;f�5vwm�N�]��ꎺ�v�4��9,j�[.�t�I��A;�"m��[�]�.M���s��;.5���
bq,����K��\�~�� Y�~�]�S��&3&Y1�����������c�I��Jʟ}��pY��f3�;���߿k�s�C���k하�YP�3�3�#k;��x���?i1~�ԉ6A�gv8�Mw�spY�N�f2}�~<��nw����}8����v_B�2c+%q1�7��s�O��&&8Ɍ�)���w�;d�W��w��=���s<�하F�?2ս~fI M�K�C���'�翷�<�x�fc1��������!�c1�&3s�{�g�/��������Y�>q��YY*w~}������d���Ș�}��pY�J����^���fD`��?}�<Y�W�_�"�w�{b����2Ɍ̲bw�����I�1ȓ��f&{ϻ�AgS��3�f3��߻+1~��g�\����1��Fc1��"��k���?����CH��p�:�YS��y��g=�1�&Y�7�k����L���[����<ed����猞'����8Ɍ�)�>�w��Y++��[�ef'c17�>�K�ϼV~/�*$�����h8� ѭ�뭹��4�{;���l%��a(��a6 dp�Ĵ3bk)�Z�����&��Ϸ�<��C�df3�{�l�2��c1��"c1����ef�q�bO3w�s���~y�VN�9���~2y��p,�Lr&'������LG��s5��sF\s[�&����]J,ь!��|N��~���=�f�u(��jxN�9Yۛ�)�{zw��9M��og�ˉM���n^�W���G��ۛ2�BVj����Z������B�BI��~�u��BL�O���{���D�3c10a���y�{�,�%egD1��y��vVi3�c1����^x��y�!J����7�0����gcjD�$����:8�Ms�saѬ�&e�əf0��_l��%ed�1=����=��~�������9�~d񕒧�2c0�~��೽�c+�&3Cy���Y��a��u��5$p�����!��x��}��}��^8k��{�+6�YP��bs�~�β�����	���7�
�2VT�q�ɆS�����z9�{��9s��K�1�LNw�{�/S���w�}N�f�u��ֳ������w�ʜ�c0�&32ɉ�~�}d�+��N�ȳI��L���y�N�1��C��K����͡���C��J�o��Xx�1���u� �B��B�/��50�ɫ3�7ryԁ�ҝ��a�:Vn;�������K]i�^�gR}f'�����gY2e�ɆY����+6�YY+�1�>��{�<O1<�{�_�~S>�Ͼ�ɦt�w������Ɍ����.��핛N0�bgǺ���:5�k.��u�N��&��Ϸ�'YY��C]�﹚����'�~�͞2��c1��YX;���+6���Ę8�ḑ���w�'YY/�f�g���K�ƅA_��~��V��:�%�{��s�q�s��e`��seO2c3,��S_~�ݞ$�%H�	�b���Cd��ʉ�W��um�=�f���%����ɤ���HN�*a��7��r���Ua��8i��eIl�SEa��/������?����ID*K��oݕ����ed��?������W���i������Z�z��_�]�k\3�q!������_l��+c���݁��J�Xk�y��c���<-޾옆$�TmWPG�g���mu9$Q&�	|"AO�����!Ԃ�YXk�y��ed��^~�����9�Y�}�xV#R
B��k�}�;H6�h�����	���"+���y�mrB$��0��V�	�gA�%�
[>#�B��1�؂�$�{4��8Cq�d�G�G�[_�",ed�?k��l!ԕ�aX]}�9�,80�7ϛ��=�}������@��vVO���FT���߽�:'P.�[�!�42e�~�G��ݕ@X*�@�_����]�g��>�������߫�HV�
�R�מ��:�@��&}�9�,�d�T��y�\�Ѱ����:0�)��=��:]fj�-ֹ��>��bIP����~����ʐP(%@׿s�wo5����Ͽ �<���k���$��j��������S�0K��\�"�{�W�"3��m��w�:�Y��S��s�:$�%ac
�?}��0�*%M{���?}�Y���"�8*�s���/��ۘ��fZ�'P���{"1�;�𻢽�[�u^ō�F��/e�C��?y5���D���������}���?}�T��~�:�@��_ﻭk4�3[8��Xo_����R�3����R��p��������������bK+*g�����2T*J�Ͼ߻++߸���wsx*9��]DӚ2n�J��!�M�T���5�ϐ�� :m����~��ߟ�Z֋�]Qѭg���T����Ԃ�Xg��{9Y(ʁD����e`p�`y�|�?}�3�_�H)�y߶N�
Aj�=��,��}SY���kk8S�M}����++%e�{����n���I�~���l!���=��aRT*K=�~쬜����ڳ��3���6�� ��-��2ֺӎ�i������aƤ-����l����`T�s�g�����ǝ���=O �R,L�Ϲ�)$�Q������
���z���nf�)n��q�A�My��l���;�u �m��{������YR
���V�(ԅ��kϾ��w�������?r���{�y��x���������љ�k`bq&w��eN�2T��k��l�N��k_^��Ý&0�
���}� ��¤�T���l��Y(ʐS�y��'bu���|u�����^~��p�w��;_�������'Qц��Wc^�����y���� ��Q�<��z�pA��&���I|>��"�cl�r����������unzC�Lc"�pv�����k�(N�n�=��t^��4l�bz����p��F��n�V��x�(/M�wv��Q.��+��v���mP�CϹ\]Z穱�:瞮�ѓ�k�
������Gnʏ'���=Fs�a&�*��#�r�[��ö�U����n�[��l�މ��^�]H�vζ�͵q��;v�r�nS7�{b1�w[�.ܩOb�0Eۄó���戛���o������w���7���w��R
B����vT��Z0*_u��p�P*jW���w�y����~�;��H(q%@�_k핇V��Yp&Z�$w���`����@x��>����-yy���$�?M4	�?wX����\�������T&�8Dq�dwt���$�{�w����t4��z�����o�	�{���<bH��j1{[=�hmm��,�U��|O�y�w� ����.;��<mx�o��~�h0m�K��� ��e���,��YY>�#�����6-[ӟ	<��b� .��EH/"h�[<��i|����Q3N��m�IÞtv��3G8�=k������p]��]0�/���@c�e��=,�@��m�$|WVA@�� �1�
Xd�_|I?{����㍒Kr���<��?��gT`'k9��gK��_�K˷�s�.h�*儞��n�v��]�E��0��5��[�����K�?�s������ĒN<��d��VAD�ݾ=��tW}v{�O��6b	�M��� ��ن�ZJ��+��\�ο�WVP�~��#�7fGw�����S���dvn�ŐI]YO��i�Q�7Ofa������B�i�F/+�~$�G����������złB�m
��F��k��^5Vj�~��֤�ڴv��Z�e��g��nr�q�:�p����E(!Bߊ\!E9	9anm��H++%A?wI��7�|;�}��_�+`�H|�(La�L��.��+�j�����ŐI+k�P'��GH4ױ��{�<mT��^���p�P�[�f<�@�Gd|EJ��/Υ;�-��>��G�[��EI݇5M�����
�<�cfT{(����U�q*/�EmS�uT!�'�j�y��9����د�����?,��(I��M5�'�z��l�و$n���U2͋6�mgU�@�;�i�~$��v4����"綅EP��DF#N(�盛$��=�}�EvUx�9��}_��� �y�������
���̢��bB�R���v	�t�[�#Eֶ�(;mʏM�������k��#��7ג�$��9����â��J��>��O���Q?�G��!E99w�~��;2��緬��Cמ�8�I�H�N�w]�L~�~��� K���(YP4ˊ��Y�����A�ns���ʕ�I9���?�����͹#qH�9V��2���U�k��'�G?g]����U��9{�=[y	O:;w�=��S]=-��O37�ﶛ7������w��J��;�E_ǿ\���/��/(�1��o�?),�?*�5��I�F��w�d�WWJ�ɞ�k��X&{�_5���`�WV�_�N�
��������C�������;W�Gs�0�t�y���9fw'"N�����P�k8=�Ɓ�������@͵����[�o����4	�}�v⧌�`M��G�]+�I��s����/ώ�H$�>��κ��X ��מ�@�z������S�`�we��u����O��-b��)p�wIvh�~>y�b� ���W���@�eFS**����%+�J$�۲ β��H]�K��U$A ������'v�9 _D��V\�OĀW�r�������0M�w�X'u
 �B�ګ�=a/{J��kK��_<�!�B��Z-m��5�y�9졷|��%K+�B�Q�t�?�m}�2��� �{�ޭ��
B�Ab�<�p�$	���Qvvb��7SܺM��kn�rۭ�ѭ(�,���9^��HZV6��w�tf+&6��[hc�Լ��9Nx�6 ��ۑ-�{����m�TnG�9ǝ���n˟b��m"����4�-ɨh��p��>k|�x3�;��6X���WRӶ��Y3�6nN��E�6ۇ'Y��T�������۬%�<[W)\��xg���<T�Qm�	œ�ح�9!Q�{\e�Zw���˔I�A#cҫ?y�J~'�ϵP?+�������@���E\��~u�(�f��!#
5V��t	�����7�t�l(�[5[~` ?V,	K�]( ����௪�Yr��L1J�D��	�{q��%�\�ݹ� 1�P�H(�k�xe�K 1��9w�~��Uc2#���*�Q$���@�����^~4Կ��#=��K���
�*BB�fӟ�:}�Ӫ}yq�Pk�j�P$��9��u���Dq�߅�Q�b���-EQ7��n58yF����
�u��E�ƪ�G_�ݿ?jy��Cg�.
��}���$��m��}H�~��]n��F���D�J]�`�-yD��O�6:Un�I���s��hK��|��D���=+
� ��	5�W*J?]=�l�s�6{G��̏`�
���{i&�˻$z�ږ����Sg��y�$��ݶ���w���c�]�d(�b0�U�M�@�H8��ŐI�gؙαm��-�jV_�ł~$5���$|I��۷)��a��T
'���3|���{`��������7�� �}t��IxʤW�ߝ���, �"h$���V��Ǘ+⻚A:��^E�)U�I~��O>������e�ys^�����l$H��M&���[F��tu����]�jh(�����w��"�]�.��H����#�\�a����L�S����3��x��B�}��jW��f+2/�38��  f�n���.�~:�z�{,go;%?��0O�7@�]�dA�(��7�gd��{d��啶����d몕Vj�(�Gu=B%�n?<�V
�m��b����W(�ww_w�����w��]�m�wL �{�oLu-�2ۡ��M�ž� ��/���X�*��O����z�+������M�{w�֤L�zy��qW��w<��%�@a+u}������Ui��FJ�r�6���3xA�T���s�5�%Ӯ�l�m9Ϸ��;��/v�eA��+ t��(T'6�:>6��]�ץ�e�%|�F�5�.��z��������C�L��k8c��X�=�ܓ�Mt��]��/|z7vz�sҷ�S��t�\^�O�ۉ�oS�SדC�і�o��Ѹ�Ҥl녩�9F���L����Ul��Tj�{�Vy�Y|1N��1M�^�c�j齔�H#/!�<(L��ۂ籭�{=J�a����
�����,�^���eX��LJ�}�s_���ih���Ѽ���ܗ��{�|�K��,*syw�n���S�/{Ӊ�]&{��kg�^�����zC蝍��Y{N�H5`t�Ul�llL�H����ܢ�J��QC�A���/5n��h�+L�v��Z�h�"����z�t��HUOA�kږ��f��gn��Z5o���BjHח��r��A׎�0!V炽�y�FJ׈���Mm�bc��:��6����m�$�8%�c9�wovlvB<����Ş/����x��P�w�֮#��j~�<z�7~�C~��z���̓���,ʩ�X��@�UDPEE�"����QU��B�+�Ҫ(�Ɗ!��H���adnf*��rʩ(,�TD��XDJ%��U#D�+YU#)1
�`�	iDR��\A@�Em��X�#mb��V��TQ�*֭J�J��PTUdYZ���2�Jōn!QTPƲ�A@U�6���������آ��J*�"��AX�T@��XԢb"�Alm�m�[kZ(�IEq"�*Z��(���n%ڪѪV�E�r�A9IXĶ�$�mUk+�¡T��Ej(Q�\�e����ikTRV��R��PZ�ҴF+V���h6� �fWKZ���+HѨ�q�H�R���h��D
���Q��2⢸��"����U�Qc�Uc������km��m�Z������mkU1�W-Z-*(��P�F2��5�Y�_s�߹9}�6l_�
�Q"��8�1݀��}^E�[�?ٻvA �e�_	ok5�y�x�{B��\�ρ�"�P8�tv\�H$�ێ���y=����'�}wb�=���&���+޵�ٝS��epMȔ4ۛ��޴-��>�|�/gru���w�%�W�wX�����s8�om�g�A�K�	��~�ݮ�	8��uR�ٗB�d�(�y�0!P�ڊ����|Fby�_��:<��� ��.�|H�]��o4����˪s�~���=�{nD#���NXjd�$�b�&���n{�4Ol�OĊ[��4�<�A>=�ġ�7�=����I�j��0�W��~:��Oh����cWf���k2�Ѻ�l��v���=���6>�}1R�����j�����y��s;;�*��o�=�֬p�x�iU=��΋�-��5���=�x�����[Y5�$q�mݶ��.����$wgP�~&����~�=�a]���c���K�.:5�f���_o<��ͶȆִ� q;�Ѯ��7f�ᠣ`�N>;�r�$�h�c�I$��ݷ`�喪^m_}b�o���}�p��JE9Z_��œ�v�h'h��O� �^��$�?v݂�{1*�{n%X|(�(ZmE@b{n�$�~ͱg�A̘6�����L��?��@�H:��`Y��r!�/�r��d�\���"^t�I�y�b�#z]	�����K�� �w��L�K�A>������#zT����b��F��(u�v��IΗB�.R����]B*�o���m��j���R��^+��d�rsy9`��W������{��i>��<���f�F�.��� ~�um�㦚-�	�.��DT&	���=r豅}�p����׮�2�b�h��ɻvt�et[li��Qq�{qQu���rz�ôGe����;q�릟CsM`.��s�",�A��1�nنۥz)��l�{x�o;���l����|��_A��=�����:����4+�5�Bv���NNy�6�^�˱����j�:�!;pd��Hݭ�vp��ɳc��;Qյ�n��:�����\�1��:P�����~��<L.2J���q�m� HΗB��>~�K9�-&�ꤸ�g'�U����)�ʃ
\f�Iez�����ݶ/�~�B��Y���Y���leiK>F2�(�*�~�ڲA̗(�.Wf���]�*�q�ҁ$[��@$w]P��/3�#J�1P>}qf]�\���� �����A#�uB�$���{:ܧ�7�� �~�~���P��r쩗(H"vt�w=�f߮�{F>ct������+�@$ݲ�R�A��\𯵒	-�B"_8ː��0O^Л��v��ݟ!�h�7m��������l^��j7��w�d�wn��$�7�Qv��E����ؽG�v�X �캡@��e�@�	�AR���t�A�Y��]��ޞQ[�s32��1!TG�e�5��1Ϗ�g�p��Yz��}ٿ�u��;{˾�)x׳.
8��P��*|�|�a�3՛����꾠D��D��pt�̪�۽�TkBE��P8�u���vJ�~&��n�s{_��	��W�	3{e�ե,�ˌ�������}���ة�&�rP$���_	:��yC=��fh�Ѐ�w:����,�"4�M�o}(�'��i��z��aq��G��W�{�0��<��b�{��h�_��+��d�:�p�n �\��v���c��0�ь�P�
��L9Q��	�o�RW�9�UV��C��D	�_�n�X)�rw�c�<H$�ܔ	
p>��f����|z��������Az���	 ��J�����o�{�}�%�i�{+�h'�T|�H,�DqT�/'@1ov�'e��=�m��T��̚�جx���7�NPd:�@��.y�[{Tς�s˷\��a�/Ѝ"����)�^�vi��vW��� m�`�v��"�a(N1��/ƶ��${�(�G��n�<��T�pJ�sN�t;}����JY�1�E9v_��������z�;(�"��I'�X�I���z����g|�2�I�$� �u$�y�nx��m���h�#LBgȨ����E�Ł�Ɣ)�b���$�~ͻ �9��ݰ��ȃO�P$���v����n�PH��9V
��(|{G��+$b�~��w�4	��ݷ`�Ϯ}F��t����=*x��jU��\"'��w�d�y��?lj2U@{���t���I���`�Gt�H��/K("Dp"T����&�:�f��vD�� �Uwg�ޗB�$�٩b��^hU!��2�B�y��Q<�w=�|#�o����w����.ϔ+<4���2�(��f��Iy��6�;��i�㆙ �����Z,&
��%ܩ@�~�샓�2��U�%]ݒ�A��(�X�"��=~&��&��\{t��Q�㫰��{.\n��ްu��׾a��.�3��dj2�r��{j�'2T����H�{]c%s�EAF\Or���e�$��T(����ϒ�f/v�	��s�1$=4wwq��˲A����v�@�urə�J5X�ՖOkw�D��ʲ�zW�a��	�<�rKnw������T"-�b��_ID"q�3���=6C+��$�o� H$o5�$�Wvl�Y���iH��B�3ƅ� ��%K���t	,���k��s'�^�?R��_I���ۺ��'�[Cc�\
�*�E��=#^�QP�V���o{��1���s#���Q�:�^�����T�|	�WcWP��,�E��{���#0=�$,Ǹ�jNƺ�pͻq�Ƹ��n�������k����e��]�f���}��r��y�tr��I����U�݃l��|�����n뭭=������u�.���.9�M�^��t9�mƮ&�b�0+�6�����3�*{;<v��PsT9P�mUn�':x��p2�;eA�w] mp�{�yVSj��ܐf���`��be��y���nt��O�r��q-n���u4�L>������|H"��:�����۳Z�<~�w��hP'�iv�@�X7	e�����ӻn�"W#Y�3�=̩Mo1@���B�"�{M�U�[�IX��TF�1a�o��J�ͱd{��7�g�c�+�g��~���(Wvm��'�;�C"_D����Z�]W��p��(��ggX�N����R�ՒfV4	��Ή�{�}P%�ƨ�}`YoJ�jn��۾1L����$�
�ޱ`�7�W۵Wu;L<��{��Ț��(�dO�%nܼ���r�V�qp9����[l0�(��,�G4��8)�4��IY��,�~$�T(�s�ێw�+��������p/Zi0�J}#���\�O�G�������Wf�������u�U��>%���_�������FY��S���P�	����|�wu���rMO�۞��w</O��4�=��������y�/�u��Q�31�=�4��G
�	�$.2�r��om�$�}���G�R��]��q��]��4H^�X�IҨWą�����0i'�P���.�%�߼�Ι��G� �T(�H5�ҙӋ��O�w�Y��r��2%�N]��r�$�E{�W�+̹O��%t�ݓ�?vUP�	��]�(Va���b�1�q���v��bw<�Z��G$�9nװ��j�߿�{}�DD#q� ̫��zI�A&��Q��h�a�������UB�$O,�O�p"S����(��8��s���y��`�~ͪ����wt�L_U��� �����R��V �����e)�:��VJ$�̂����.�d�B�r9���^���U^�����i�ݸ�fB�U��J��m��P髿P�^���B*���~��l�ҳ�u���U���f�Ͻ�=����}�PWĒwt�z��t(Ђ8�)˳�ݵ����o&t��juJ$����
!onҮs2%��E���Y�C�^� �""�j�mzP ��3l_v{<��^�.N��T(I5�t� ��w���ر؟]��d���]� ����K�
����U�ֺ��d֠j�G_�y.]�Ĉ���\	W�e|H��n�7�]
��N�����Q$��䯁+�@��IqB܊�꽿��h.Qݛt�M2��.o��H$׽҉���v	A�0O�L���~��H!1��R���|I%goP���E��w�}����8�;��30�۩#���d���x�r嬐D��DB��n���J�ò�e}ݟ]`�*{%��:�+ǌqY�\_\�R�k���u�dn������g0�#ؽ�DC$��=��n���K;��[�W|I������<b	"(�(y��@�A̕(�|G����h����Wwm�ǺU
>�t3T��D�S�"��ˍ����*�)�<k��캭��w\8�R�(��f��}��H�����J��gm�$�Ϫ�����3z��OdB�o]���%�ЉH���z�P#ʫ�g[�n�sFg���vu�'�H��P�������T�����W�}�6$MȨ�޻?Ϫ
_�[�z��^=}8�I]���}U�}^W4���D�o?�s����?�Rq�?�5/� wJS��_:��=n�H��w�?�A�)O�q���(����,�+����S�(ݝ��U
$��W�>�b\���W���ɨ
�e�H�=�J��*w�~�zǮ�U=�[50!s6{��+�����6I�a�{�i�s���'gt���<��y�ö1x˹�C�x1-�ytb�9�{T�t���%��i�'���/=7��Y�'Yb��8�}��+B�ڟ����xO	�Y������,��q����P��%Zn�>
�%z�8)��_�f�=�|�Y���;�͘�ӻ7.Q,�;�{|9������ĐҢ��'�ɾ�Y�p�$o�|�؃��7�?2�a&�dޚ��y���p'�;�^��׾���f�!4b�b�d�m�ʹA.���l��L��r�����{��׳lܞ���nNk8N[�����Gw�,��wI������� ����{n�qPF��/E��=T�j�7ZS�{���~��x������B�s��.����O��^�޽�^��	W�f����G��m�L[�ǠL冎ȕw����Ú}ӴÕ�8��p��sk�à:x扃��P�5xyG2q�A�=�wڄ�W��o�O�Bn���6iO��/��ό�N�}�x�C����:�p�{�'L���>�KO���$jO?E��{�\�Ca�����rC�)��/��lJO����D�n��+wF·��h�7wY���=�ꇺs�VL�s�T7���p�r�m���*��P>9]��%��]�~�<㣓���.eئ��Q�����C/BG�S�����ѥL7��d�����G�gF堜���`7�j�3`�7)�۝1z���
/�G-m��U-UTU��ferڕTT[E5�++*T���EmJ����-��[մ��J�ԭA�
1�4����3+J���P�JU��X�V��mm�@JҌ�J������Ũ���i+(5��b-�Ғ���FХj�Ԫ$QJ��*E�����������Q�)X����KYR��,(�R���e�QQ6P���b��J�1-��"�� �lU*4�RVU�J��JQEDXQ)e�F�-��J�Q�Z�1V�-Z��J�Ym�� �aEEJQ�-cF��
�JV�����X�ƴkJ%+jYE�b�E[jZ[m�Bڶ�F���-�ѵ���-"�UE�A�X�+E��[j��Х�E��YR�KJʕ���֣F�[E���j��ED�����6-[V�)A�j�(����ĭcmU�ЬD��-�D�_n타������ri^�<xςD��ݸ��[��TnC�<n�M�G�,^��>wϘ�;/b��^��SGg19�ve����3�g�T-�z�cp�r��f��p��ձ��u�ɲ���4����#�K�r�nz�̡4�r]��Dx��z�Ol'f�cg��{���+a��ɓ:��ϡ8GX��#�x��>|~>Kl^˽��]��ȁv!�z�۞�c �dիk���W]�oM���P�k\scNp�쁻m��tӬ�PH�4�Pe:���v��&���}��1n�܎�{�s�1���T@vv�q�]sU���)[l�yv�w�=����v���������68+��oj�{W:#
��1/q�7�n��7N�L"v��q`S���9{y���1�x�=C%�t�l\�B���
r���ļG ���va�8��ֺ�b6;4�m����ӌ']r[�2y��&��7%���$�n�ʞ=8\/e��:���Wckl�;��ѯΦ��v�A�G8�nx3N�;q\��W;ہ���w;|J��[X^]I���Uӯg���sw4�̛-v��븚�<�z���7Ϲ#Y�;��z�wI�{gc�\��l��n�����ĉ���;�����N�i��e�S�Ӱ�����+{>k���+]�k�ݸSc���h�kn/W\��݇�ݞ�}�����z�8nM��v�<�S�/<[�g[��P��v�bp�{�-�xsF;uӇ��]_6��[{nL�Ծ.�R�cag�����h��`�ݫ�F�gF򀩰�����q���R�:�y����Җ��ֲ�<��z��xyp�k���.k��v�tKvR[�]�\�O�d��$z��gv��麃�kF�ٽh�.�OL���ݵ�ٲA���ؤ=�ӻ&�Nݱ���i!�k[M\��ϳ�;e�u�V�׈��YX�}��H�m����nc"��m���ntvu���e�B�5Ɩ����x��fy{Jv����?2>�7M<��=A#������u
3�6�W2�l=���`9�������>j��^���_�v|^���&�6"���nݷ)�z��7E��3w4�-=q�ku�\pf]�v.�׷i�V��`pѫ��s;����un��gg�����@ϥ�a����`�q��>T�����r�wmb� {V8�:���eڶ���(�d+q�˖N^��M�u����-��K�������,���C[��K�C�nN\��}���?��A$E� };:��O�T�I?^�A�8v��>>wޡ`�yT(�&���"�hq��^�I~��.�y�۹��A$�ʡ_�{�L${}\����ng�GY¸�#���A�I�҉��[���]�$�=���G>�	$���`3����q��:�Ŵ���w�L/?��_A$���(|I�5��bװ_Ď��
��\"�h!1��R�[�	���`]�Y����W�!��ċ���͔	���k�9"j�v�=��i��͇LRE	�����Cڬ��=��H�)��	�
iS�=�Ï(�L�>���'t�$t̕����l{����g�/���Q$��ҁ#�ב�c��	E9v�g]�|�a~x�A5Wj[��>��JR�(���΃S���Gr/^l������A�V���wq(/=�J���>��<*w]��4�
`��ʦ��&�I>��Wĕ��b���fx�3����4���z�D�bI���<I ���A?��j�E�f�ψ �܂�wf���<���8�9w�^��*u�V\�I���O����w����SZ|���pW��C��_�k����q�@ͮ��'��jQ�Y���U ��J$�W�z�H�B�S�[��P���N8�{=m��n:C����SǤ%1�5��ӡ����@�(D���[Ŕ &8*W SΕ� ���Y��j�!�I�<��N���zi$.�۲'�QyF��:�䯉 �+�g��F�����~$��ڲ��P?���߳43�U�]]-GA��%��>��v	̕+�A �Z��jT�e��x�7轜�Gv���M^���uy�=�qNtQ�۫���Z�	v�b,���p��h(�h��۷�w�\8#�ȶ�p�]���� vJ�D�>Q�1R�&dU�}��Iu���$������wJ�@�޾��z�z� �;��_׶p��H�HD�X*z�|A#�����uw*$��`=ҫ����D�"O6#^*�_T$��b.�==�u ]�㍻c��#�z����nϐ���1��&����q4R8x�V����PQ��(��B܊�];1 k��X ��T+�k�+��.��:P'�9+�Y�R��Yn��� �*�����@�3~�ݵ�,����h џH㯁�A#��+�I�Q����uOo� �l�I�`]^Ii1�d��������T�/Q�����	�I��(�f�7�_��S��cO� NS��w��Ww��X3��7M5��+V��$u���=���.R���73s#���kѶ�^S�r)��Z�uy|NC��&
��̊���J�I盷~�ovL��o�G��B� �g�e��m�����kzIk�" S�2	M^�q'���E�5Ҫ�̛���+�Ͽ�}]����D���N�_	�ݬQ ���~�r��R������|J젫�����G�o�Y5�l�✫ef�`$D��T	s��{u*�=�ז0�z�	�
�m��_N>λ�-��}�^���{�|A:�6���W(4g�8��Ӳ*T��{y�*�#�T	$���m��}PA0���s}{�������Tf_$���2BQRU��Ϋ �<�_�)URr��s�� �����#�U}�:˝%�w���l6�n<�}�ݱ;U��H��؟
���������W{�\��"�����`�<CE	Y�g�sC�P{ex�J41���z��P�ԙ����N�t�Kxi �\b������t	�a������7n���,s���e_7X㵭�c��v���1g��PG:������<�i^�^f�l�Wk^��;v�N'r��M�l�v�r��ܺ��K���⺑GE�lv ;<��r�c��Y�q>���֖M�v-Nٳ��_t[a1=�<l��Y�7�F{"֧mtٛi��H��Ft�*n���	kP��p�������;��0�m&d]x�ʾ ��7n�'�yΡ@��;���~�yP$m��u�݅r��+�G��J��y"�gE1Q N>ͻ���9��=ެ�+E�6s|�W��q!\�L������G%o�X �O��ֳ�Q]��O�wn����:
�S�WP���@�v��^+�yΙz�}�}L��{u`��9�Q$�}�����F3B���v,ű�(4g�8��Ol�Ar�TA^��k��Y U_����2
 ���*1�>�����>��d�QR8��=[�ڻ(��'�n
s�@Z��{�������LpE!,�/�=7:���d�� ��*2�꒤@�޻9�P'�(^�P��fEWμ�y�={j��h��q��3&�e�}�	Ɏ�n��Ob�A������+��q��<��谐B���i�Y;�P3����E<��f^�1��X �s�P$���ܨ�o/�|ƺ��z��#�t�~��#(D��z�P ��܅���^>�W=�N9�(��w*l�1A�#��/�}s�_�;i{9�X�o=+�A$�{����������C;깹B�50*�0�-%����:�,a�~����eU}D���Q}�^=��-g_������tA���Kclc��蜮�pE���=3ќl�A�%n',6����/�rk����D��\�~�G>ͻ��}[�w�(�$� ��UfߊZb��1).�~��I�];m[�Lޞ��IZ��� �y�m����^�;��`�����BΉa�S2*�u�_OǞnزH=���:��nz�UU��!V6��ܧ�m�ܣ[�����77�@�y���ͣ�u@�ޅ�H���C<�����g������ft�^�b��}s�4��o*���lY��x��"&"(D��*7ڽ�`������՟�|2�� ����A�t����Ǎ9��${^b�@[2�f&�H8�p��%w����<���������'��N?f݃�?s�_^$�j�ޞ~o�@�ʀ�Ɇ4�y�cvvgݎM�X�Q��M���۫�QT�[(�w�����bFT���$�WA'g_�~ ��u
Ւ�˕�3�ܫ�A ��۸��ną��%��@�
��E�W@�,�;�@'�n�'��	�%�_��zpn=�ņu�H=��1)(/o�E����$��u[�~Y��\b��夓�۷`��u
kɐ���2��՘�5"����W�V���M��ꬿ�A�hCVE��sÄ�o��Κ��Y#�F�<F�Ba�wq�������~�߶n��Y���ȩ3���zC��,#"��Ğ�}w�8N�"6LD�Y^��I �.�_���}�����f�m�lʡD���Qb�}��Y�������`�q���CY���<<�qh�lV��8A���(�>�a��R6PqH��rU��t�Q#��TF�������wX?�M���i�(R��r�M�Ov���Wm`'�FM��'��T	D��ぶk�v_��&?�E!	��1�9�L$A�	>�U��'��/4�}�$��@�F�ڨ�]~+X�8�Ĥ�/���kK���SC7P$�%��G�TI?}��]�J��7��|r����hB�2'�2��n)k��G<ͣ^�D���X	���=�D�5���[�W�(X��>�X9lT�2���y.���yViR����3��Ճ/L4�[FV�n���P���������Y��Oo��;|�N{���M�V�y�ٶ���:8�5m�n×�˃�9���`�9��85��q�/X�ɞ�����>�a;r�걬]��
�܌j���jR��WB��sӈ�knb�#�Ǩ�f��4;@p��k�D��P�	��y���8��4/7�2 9��v=�XI�}�v�iv�BX�'<����Nԙ7=�;�k�Okd��.hJx�@森�۪ye�`�v��-���G��˜=m�ծ�Q�dI��	�l!�LD���8�E���OĂ~�۷f�K��r�oo^�9��@��1����R8h�{Y9�'z���s6�X?7ث�A �����i�w�ؠHu`���� ")v}ʁ q�uX'�k��v�muW���#[���u�m_��1�aL�a�J=7'�z��>�V�mxn,�@$���u��{PyE�{�3A w��P5��sGb���αd��*z���լ^W�T�q��(�y�6�O=���$'�\~#�*C��E$���[c��9����f�=�l,�rgu�@��`��=Z���};�{��L�d]�������ڰ	����P�k�=�-����{뷜�O�^v��E��o�	�`P�.��z|ގ�[�� ��UY Z���أG�ͬ�p��!��Ljf@^U��f(�����{�a��Z>�����������}��M�^�6c���1�Y���~$y���$�T���)�ߥvgE�~+�kcn(q8�%o��jWĂ{�+Q�A;�NQZ}��$u�z���M�U`5�!*8�Հ��]�]����i��I�ʠ+��Gk�.`���{��X����0�b0�%�rP?tY�x!Bv]����r�6��O�U
$���Q�}�Ʈ�i:�\"K�>�"�� �Q��ֻ\6J�ˎF����{B�rv"�w�����^��z�g=ݶ,�F̩@���W�}�wK��6W�����N�o��R9���S2.�-x������,��H�ʂ�����$�2?N;fٿ���7�E.��فB��z�|G��T	$�ZFM+5��Pt��y��.H����'���+ԱyZ�,��d��x�'�U>>�[�ٰ�d�߽e�V��F���%������ł2���(L�<�<�rT��^[�Q����;��đ�=�|�[ց��s�+9I��+�o�>�|e��� �nnv��� 88��dJ/%M��	<��k�$�<׺G�^���h��N����!�_|���t��~���1�������{�/F�sʵ<R�r�R���oPqR�����Q�7}��ވ|�\��k��S�whsA�*�}<���z������|��6i�j�Ȋ���� ;��S��H;Nq��~��C~>�������lM3�xB��e�h�S%��	�y=�`�,|`��5q�#������}�d���i�}���؏je�ϐYU������ּG}���>%��HGP@g��;q{�O���ۓ����nIC+�3w��8H��y=��<||��|��[��ם�^�^6V�j,V~�.�����_vL��-�5�x�ܩ�I�ߖO3�x�כ_?up	��^>ڰ;�d�1�:y���|t�z��ң#Wj��ZEC����T�zf�wS$);X�,mYFﺃ�E�O����'�oN>��� Ю�Ιtk�(�Tt��{=��oS���Ej?��4���n{'�Cdj-�����T��󽺚�h��z6�x�W;�Q���X�8�8bE�f��^<W6�.�cR�p��?�����
��h[U��iKh�F��ZJ5�Uk[Z(6Z�+XQ*��յj�A�*��-QkkYFڭ�m@F�+JԶ"�Z�-��V,�+Pj���Q���Z��Um�F��(�ҥ�E�J�mZ5E�ARѶ�k*Q�F��*�mQmQmlj�[KF�(�E��JV����[j1UE��j4�")Z�V,J!eh�Tj%jZ0�Eb�*��*Ҋ�A�JRűEJR�R������Em�jV�h�[`V����hT�U
�m�+X�QF��K
�mF�l���[V�m)k�Z�Rت5����*+m�Ң[B�PeJV�*�E��VVXԣ-l��KD���
UQ(եX��-�V�kh�
��+m���m�J�U�-j�X�օ��[Z[mm�ֵZ��[j�b�PD��߱T�_���?l}�P)�k#n(�9!%m]��o@gA����b���Ϸw�uI{���O�u�HU`�D�D��BGv��U� �>�a���b�96O��
$����A]۶.n?D���?{�c�?�an�C����fk����v�v����0�n�y�"&b.''�](�z�⯉�v��7��|�Ac�L�잠+맼�
�í��1Q˰}]�v~(߬�G�����+͹�I$�=�@��+�6��v���;y-���h���Hi�̊��u�D�O�vfز	�}�}���	OyQ��m�g�ᢗB�l��N]�T��ffD:�z�����r�I���I�����,����ۨ�I�gO�.�4��hy��yz��"ύ��b�m�F��`{�1�'_�p�o+sѡ�U�V�U�'i�/����P1"rC�f]��?=�F��&�E^��X�|A+�z�~]�B��ߣ�3o�9��p�J�x��X�;Z��q��-��tV���%ٓ;s���@��BGI�j�����vA��yo�FM�z=H�iv%�5',�P�)���F�nWě��E�q
u;G_�<X	�Hٝw�$��n� E�$Z"��Wo�.$Ug����G���߼���>X A�yMv���e���_�D}J�Bz��h�e3"��y@��Mur�+Q�߻�d���
��܎��������p�K�a6�P�.��ʔOğR�Tw�L�����{�d����A;O��@�矮�P�P���d���y�У����j\p����/NNs�W��{|[C���k+g�9؞d��{.���� ��h�o�i�Y���!BP0�� ��.���sùѮ]j�5�������9z+/M�"u�9�q�\�4��O�v~d8NW���N`a��n�{Xp��q����2k�=8wL��{,�p.C��ָwg&�luu�+�z�J����/0��vcv�gn5�c7-�۵n�n�����ۛ����krv��;'���n����1�jrR��7M�]���m�nR-�,�Ѧ� �`ێ��6'�%u�ϐ���ۦ4�e����˃\ɐ1rC��]�l�I$��ܫ���]�'���^ʺ��T��-���H�Ï�P'��|�R��S���,�&Т~'m�*!Oo���^Y�ym��0`qI(��J�Z�TH?:*ճ�l�����>��WĞ�ܨ�Wb�"q0ق(�N���XW��++�|O��O���
��v2�fy�$Ou
x,D
�A2��P�u�D�B�αs�J>���O]�'��B���N[�TH'ⷻ���p����� {���P"6�IBaE	)�^����1+�e5�#ۢ�/C�W?��߇�+��+nN��~>�ڨI[��ܸ�9
�������?z߱Q	���d��7"��꾱d�*@xP�-����c��w����*�KR7ǉ[�$���TN��{�����i��hdp8_��
�0G��Ի�`�o[#��=y)��$I��g$�V�u�$�sy�_Z������xD�(E;���4�$��۰H��������Q?���Wwu�"���e�`��Qy��t�xN��s�|��ĂJ�ޫ'��t%%^�5@��d�F�ݍH�L6`�9C�{6���6}��?l��g���ҍI+;v�^N�@��
�
K ������W�W�-5�ĝ�����*3t��SQ����d�r��A�WBi����Sƾ ��� ����(��b^*����0�����dW�FKn"".]�}�_	�<�M^��g?$I]۷`��:�W�66��aꇭOd��?Z���dF��P3*���O��T�A0�����G*��]�F����g@W��Y�S�%ɗWUY~*����ɔ<oYЮqW�����?���b��_T�.���<	�y�b�%�U
����K@�����T}y�ˇ�f��w�W`Y<ꂉ�����뾝�}��ܰUne�����a�Ka��W��d�=5��i�f@�y��_U�~/z��A�ӈ�(jKٔA�M�҈��5��2�X�A�}y�Ah�� (O�/��?0�<�����1$l0��9cfnP�ܩ@�H'gN4>)^�;}#�ڏ���KΨ(�|<%l ��A��#�}�}�{ց��{T,���B�$��Ɖ(Uz=��f�`�i@�qr����Iӟ+}3����ZS�3�_��
:q�H��"�G&�T�W�Q�
�\�F�l�	�G�M?Q[ݫf�8�=����྇��b�܋���v��J��m��no���.w��*���:��W���6��c�������e���
���@�P �l����l_I�j���R�'��ˡ@�FL�k�H]ݴ��HVQ�z�����v���K��*S����D�5���(;������n��5rb6�a��p/�%��4I ���l)y�˙�����(Q?�|O������Â8��>���|\�:��b���`�I92q��!wn��	S��qu�1_�ϯ��@���(9|7*x�Ăfm���\�z���s	��zd�_J�ݻ"�mM@�f}4ll��~MF�3׳�O~?�  3}�۲A#������ܨ���H��MYz�O�H�7"�2��Y��R��ߟ�2J��-fK4	.�ۿ�mAC���Y���_�Ȳ�	��?e�w�ޮo��j�F�&�
���z�U���D~y�$+ȷ餜��s��J��	�\����H_v�	�&wQ9�"�ӛ��^��M;l���RR'h�YĮ-]Y��$渃��c�����t�#�"�KB���n�pU5۲t�q�l��vW��vy��˺�J�b�U�Lx�\�xNy�t�y9p��rIv:D�{ql�O��U�t�֦�A�G&�$یIȝ���c]�6t�i�i	Ny�05����>��g���볷�ې��[��v�8[h`]�=�È��ÍC��]��8��t@�tWK��n��Es�`��I�{�V�>� lǊc���~+;���	�ڡ@�j���XY]�K�h�H+wz��yZb6�a��WǦ�M�^l鵙�S��> ���W�'��ܮ��5}�"F��g�ݷd�veJ$P�fi�p��4	'����T+�oE�	[,�Xr:�<|j���Y�;pQ���A2��@=9�1	�f� }]�b�޾T�3m��E��S�}9��Y�"���}*��,�̪OĎ�8��;o�w*�q����&$�m	�tU���w2g�;sX̜m=����L�������$H��p3*���zuJ$���Ɓ���>~!�ޮrn�ǧU
��ğA P6c��������>���#����nJ��<=�b�G� O�>ѹ�omË6���#�/g�G�����!��v���w.�����_���HQ?7�q�A�v��wE��O/l�t�Zb"�A��P=7%�����`qU���}ӳ���B�$�:�D�vxD��$*G.�{��ϰ��D{.ை#�u�����i3�����=w�4s�B�?gY1Ђ�e�#��<��9�ml!ۯ���W��A>ʚh�y���wM%�����-���i����]�{\m��Zٺ:\�p�^��Y)l�4����}�3f}r��z� A�OMA$��۳�}�.Ⱦ{r/T ��q���W�eRf��Ő]r�E��f{�(O��~��Q�v���s�ona�Na��`%{G���@�l�k)��A ���e��t=�7�\W�4�#b�J#�+�;ٴ����B����u�6���Y����5��q���ç�O��=sH1���o���2�=�&�ej��︟��8����n�S�i�i3��@�܃٣39s����V�I�S�D�I<���~�@��o�]pE?N4ks<"F�%"���[� �+�}�P�_�u?
ܒ�6�vł	�����F9|r�y�~���'���ȥ�\)pn\���[�����=eλx��s�SD�kA�����YL��}���ƾ �~ΰ,β}֑e����T�_�?~�g��3b}r�ys��_{f��wo�|H$�-���� �A���~#[s�x�a{�O[F(a�E@�]��d�ζQ$�t����~�����͡`�u��};G���@�l�v\�&�7૯A?�W�Y�ζ��{��t����s�j,w��wܔ���'�)����܇0�����z��ߧo���	?x􈺞&���,'��Ɵi�W���?�wT64�G�n�$f^��'�2^X�*<Vف6�0H���:` ��ƌ�NL������~O���yb��zh��x��>M�e��JH6Mu�6�k��MTէmXǕ�	T����J{�����n�h1"R)�g����I�Y~'zM5�z^D]^݂O:����Id$��a�맧�����J��o� �H'�u}@��4�$��~������P��R&'�*�Y^��'�}��IY��i�����`'je}D�7��_a{�O
a�D:Uo��4.�$���I$��4�$Aם�����]yR���.������1$
�wo�i��=���Aȧ@����I��#�vػT=�;�z�=_&9��993j������қ�����P�G�������ËYgV����L�<Ox�s>_,N�Q��ۜ�x<��(��ӥ��wb���:^
T��w]Y^�z	�툑�.�'�}��.~}��{�^t9��ږ��[��2c��R��v����cڀ�t��Yވ�|pgT���օ�*v)��Ӯ��@ξ��콧x�[���@�-Y�6�ʗ��Yt���N��N�}��*`j�{8.�����oo��3\2۹��¨��.�6=�Y�_���5�O$������/vGé��%{���d~�y�X���h���T�ԥ`�П�V�[�*S�K���WK���:�j���VOo��t,�MOy%����h:*�o�N���2I=6o�$+���  w�z��ƹn�4O�����AU�g����n��O/�y��T�]��C�jyr�2c�;��{�����d���2�ɜ��v>��{'��d�?{�z�Z�ui]ٲ��H������?q��/0eL�'��{�y���7�d@��Sћ��FۑL��N���#�y�wu��ucѳ�
���ƽ��@it���PO,��н´������DX���Ou�1W"gݾ�oko�5����[�]�لԮ?,�w���!#S����յ=t�!��q�@7|m|V�3���R��ISn˻�l���oH�J�Є�_vrWQ�j��Y<ɽ��4��kr�^�}1��L��{<���vL��D����J� �{�m���M���ZҖֈ�V֢[EDe�
��k*1��ʒ�����%�[m[m��U-�RԴ�J��*6��TUQ*Qj�KkR������Q%V��,��ҵ��ʢX�(�h�lh�R�J�AV
�ڨ��Z�kiER�XZ�YT��5�*ը��QU+(��h����R���5�aRڡR�ڥD�*��-��TYZ�E(�ڭ�-JԬ��m-E*4�+,b����Kh�--FU+V-�bUT�VX�1X��DF��PkTj,��Z�(�X*���eKJ�UF�KJ*
��J#([Kj�"*ZUTm�iQb�[F�m�-��P�QDJ�҉F�V�ЩmF�m�j(-b����ԥF����"[V��UA��R����cl,�EY[S�<���5�>��|
k�׷9`�컇wV���q���i��E���n�v5�"�v��6�	�`���*�!�틳���b�tv;_���+U姃w�A�]<d��WQ�xq�ݸW��QF(9�=���c��w>�dvG�5N|[���[`-����=P��\��z�˵�b�(%��+����^`��/�w1���k�Z��;m�e��� �an�����E�n�=Ȝl�\���]�}���Y�ˎ��cE�7#u�P��n�=�`�@���6jqb^���z; ��N�3����w`P,��vT�����˷�<"콁���g�L]�p�0v�V���v1Bq��\<�7\��y�Ɲ�6�<�SJ�5�w���/N�sh�2��p:�[�F�)�t<bc=�v��j{ :�c5�/i�ײ�m��k�ڵ����[��u���&^à7 �����ڃ�<���9�C��q��l�`x�q��{xX�K�>ط��z4�T��Uo���O���#��FKR�k��q6�3�B�M���y���uү�)��\]��'Z��q�O[�8���]�N�ug&����z�u����k��/��XϢrs�͖S�iΗ��D�m���[\q�O5�Ü/�]���]tm��k
X��y�4��#��l�٫�pq͉�������jt��ϝ�w;�[
��^���t���A��S��d��ɋqu�8��u��Ps��୨�q[\v��)����ۇpVm�m��^�vm�G���j��ݐ{��w��݋��mN�����;u�uݯ<�[1���>$�+c�F	�oL��F,��n�>s]��2�v6;N�zڭs������8u˹r�ʅ��t�%�q9	ܮ�u!�l������0�.;m�s\���Uf�iw���om5�k:�Ң�n�Ѻ�]f�v�7\l� �f*��;ի�k��`���/8�s�!�nwL�n˞�ϳ���un�#ѡ�v��9� QϮ�;U�d8�W9୹C��]�p콶ڧ��z�Ny��6�r�&�4��뱛hT�;q�mɫh�	�n�v:���w;j��8�*8z㵧�c�d3�l�&��9C�OV��K]��F�kW����C|zl�,w�T�1=�:z��	���L�����r�v�[���ti�� ���c��U���׋���������x�2��g�b �v:6�Z�� ��ю�}��~�܎u?��W��O��S�@��<��u!l���]
 ��S�f�$F�H��]����gӢ�,u�{��O��O��8� �����&�ǻG㊽v,���¹��e4Ñ�ܞ"�$��m� �Yzڌ��Gy,���O�S�H+����=ޠ������E�.���h�XycͿUA���_�%gvՂ~'ﺲ�]
�8�����N�h��|��b1"Ȩ̻۲	=[R�6Gy�ɛ$IS�I����'�*�y���G����ߖn^����A��d��HR��g�{����v�k��F7`,�Ս<ѝ������ڝ\@َ���4	��Vom�$��uB�>�u�~�*q�I���ڿ��v��S���tmd�A8;A��gv�Y7r��\�P�T�K/���a~�4�y�n�srg��٤�f��6�	����+���w��z��^����g�O�����q��H+=�W��PP$׷�g�I�7�tӷ���A�b�:�}[�X ˩D�M�w�h�4��㤒
��n�'�˪O׿:d��SL9ʞ6j��~G�"���`�Ge�
��OWN!�5X��O�#���}ޠW�	�	���$�������$L;�^���uB�$���h�AL��7���`����d�^[Ge�;\c��s�:0l������qm�V2�L�y�>m�fI�ȸ̻۲?�u(�	���֦e�Y��$zge�|O��נ���Rb:S��@�]��SȸS1o���` }<�
;]4�$�V��&\>]3�����ۄ��N"�q�;��Q'�^$Y2K�z:5!�<�=0B'��2x���Cv������ua���7t:����&*{�w�/0���顪��C6�A����ݳ*�a��l6�=� �.����&��`0��b�N��=����{�R�����=$�l�'k'$�;]��� '�����8�E4Ñ�ݕ<hH<��]KJ�e��̽� ��z�A#kf$��;lX���TI��7�4�"'L2��+��9�9��9��C���E�6�6�����n�EנNh5�8�O���$�u�m�|�3��A���(P$W>5�%��6�2\�F⯏U�زӧ�`�Ѷ��>r�a�I����	���o(����I{x�.% P&#�1��Hc�۲	>%MW��v�F?z�a�� �}�Y���	����ۗ�|��ǢO\�����IǙ�`��*F6��z�j>ں'Ej�OH�V��*�.�K[<w��@6�^���mzwh���z�c���f�=Խ�j�>�k�6��V�oāUS�+N灄6C�"w��`�J�r%�7FC遙���$�~�,�*
�/wv�+�K�*�Ͷd��l��	.���v��ӝr`y�\u���Pb6��������덄SL9��<��6łOݒ�P8��TOʎ
����@��^w]�ٔO@\��>��vUߥA�S�TpW]�:I?os�������:�e{<o�c!7�r��U__�I�T����=�=7d/���ګ������۰A=��P'��|�P��1��s�]}L5�ҕ�M{�(Y#�U
$~�4�^|�1׉�U��%e���K�!!?�3�Twr� ���}�Z��J��=������>�T(��޹��;�I�%޵��>
��8��q�/k�7�e�b;���)!�d�9��ow�m��}�;�4�����l
ε�ѱ�-�{q�~\X� �p��:x�dܜR\�wV�ak�&�g6�X�,+�8�]��Z���ങ�V��n���������u�W:������M^���ή���z{���O��c�q���ֺ5��{n����J�=<�������0l�����8��g�`^���u�V���Lm����u�7��۲d��V3č��M�����:��i�v��H�n�N�)lQ�}u�I�v����r�Q5EU �@��0����b	��-H��v�]��;���$��h�(��
����;o���ʯ�,��F�)���d���v����wg��ΕB����sMA�j7���j�М��#�}r�w�D�z��;ї�R���Y��U�~�4�V��A� ����W�KJ�9��߉��~$v��D�y��J �'՞�M������>m(\�@���>���$�q�m/$�1<�Q=Y�(	�������l\u��=�j����&B��z�8,��e��@�L4�5��@�ոXm�?���ۯl���|{+%H췄Q?Ϸn��z�^�|����2��(�}�8���Ɉ'��"u�{�,}d飋�X\�W��c*���Z���;��<�������e%��:��\c���{ �9�o��{:?�D��4�LK���]hY���o���~$gT�D�N�ݡg�3c�h� p�ʿ�D	m0�u��7��60��G�8�=?bQ�`�:�@�� ����&�$pO�.P>��z+�N�����SI<�6�A#�U�gP7��n��wJ�3��%Hn*���X=5�|�{Dks�;�d�H�w��$��shX'�(�\�۬���p�ʈ��Q�rSy�v�S�q��y��q��Ԃ>l��Y����͏�,�,)���@��8��Œ��쮉j���- �H>{�W)��'͂Z�=���G��ɩ�I�O۾��I?��,�<"�:���o�T/7�h�=�& ��Bԉ݃=����	/c��Iɴ�ю�:�e;�e���)x"���C&h�~��[f^���QЫ����}U��/+��,p�e�;.����Ec��xՎ�s�$q�m�`�_I��:<Z^�d ��	��z�&/���ʭ���u=�d�G�d�(��5-��uw���ޒq�������	�e˳�� �)��#��l��xb�Jy^�!✨H�sYUv)�Co��q��JG	0Zp�P�QlqNG;7m�-����ӜF�z�;����0�ñ@#qp9*�ş��S$�H�s��:�;�,y���@'�r�C��*�P�#H���\�U|H7��mp}����'�e� �	���U� ��1WĂ׽��t˯|,�T�l��-O�qP9��`��1
'�.enN���z��	�s󘨐+g�0���"w`���o*�o�o4z��	>�1WĂ~;�u{Bl~埨K�S赴S�q<x�E�:�$�����o�V�����Ճ�� ��voL�����1��]0pFs���eg���8{�E��ٵ���79
4�l���SL7k~�� �L����{pՂu��ē�sU OĞ�`^Zk=��=x�^��V��@[�L
x���m�Ꮁ$�<�;8Z��M��4�[4�~}��߮"�	�e�qX�ʉ7�jH$oM���׹�g������׸��~=�_����%HN=*���S��d����5�����5Q ��b�9X��V��=��=Af�*�P�#H��h\�9Ӷ��B��S����h$�zEu��2��2K��*=��qp�}_�Έ�>� �s]�(�ut|�_<�~�h��D�B4�R��w��$��L����եB_�9���׹�`��b>�1�Z��eCW�&��W��+����#�|�=�!P�.�Oi\3��y�[��N^y�]��)t/x[��)^����E&�p�̀s��l��9���Ƙ;bg��������c�J\a����k��qq^�Ӧ�Nu�[��m�m�n�J�\�!�F��}�E�X��Z�Ȗ��q�x�z��WK���:��)٘�k˼ɇWgm>+i����<�i�69��pݍ����{6�N�|�.�7�çj���3��9՝<v�nyP�'=���V�r;l�/2q	7Ms����ۂ�np����nv:���k������s}�)�����ƾ$�y�b� ��b�}�hNƷz��W�����vy�s����|�r����@�%o�ok�_	 �<ݻ �:9�P'tND:��w��V}�)Ou�Q*@p�9*�łz)�� W��c��
�{��F�͡d���T	�-[.$i��q[6����&���Y=�D�7��7����W��Wv�|I[~���R���XEϜ�QȽ�'�<4Uȯt�5,�yV$�9�� ��4������ �"��q(�ɧڸ۪x��eV�
wT��9ý����A9��p`!�E��7�� �S���fǦ�����N��=|ϸ�^���~=�G����/>%��q�������}SG�ޡ�����k:��{�E�������Z��){�\w���]�|\ո�b����6{�h��йd�7Y=W�<�D�s�RGUVg 	���U�?�ޓM�]z�o�dۙ�b�Ǿ�j��6\�+ʽA�M�|k�H�����x!�B�.VH��!D�I�W�MDc�Ĕ� ���k%f{s�Ҷ�Q?�L�I"�'$���;ZEv'��\���w�V���E�.�\�D���o�n;9�~��מTH'��9
$������>sm��;N�sg4ۜ0iX2[dy荖��؋��c�lf.-�W���/����CE>rE��[���S�$���n��U������	�� Ma�D�ADdR�Wv]�q{�/r��V0�Wr�����[9�Ewn݃�N�>��wHh�)���ȶ�n=���@�	���۲v��53�r�B��Q��:��y�gv�:<p8����=�Ue����Ҝc���,�z�ˠ8M˞}��R�*��A��z���~��f�����n�gs�c�n�뷡�/)�l��˗�I�Ln�{�M���A@�T��6�C.�J(��GO�k͇��d܊�2Xl�!�\S:�=t��������D=���(�9��ԡ�V��8��c�_N�u��o�v�յ��B�����2w������w�pk�'�(���n�LQP����l9=�n��+��A��S��2D{�����M���[��^/(U��W���g3d��;'i���|��}���L��/͂qx�C��� 7u�#Э���^��L[c؛�Y�������&n�vE"�@��>�[�^-�G�mמ~n8��˯8ENz����ǀq�A+۞"t?<׋dza�O?c����}/[���N��n����A^���]5#Wఋ���b	�>v �K�@$�^�x�tJ���n�6����#�:_6s����n�ûW���y�i�&\))óF᨝���p��Ͷ������<|�}�.��?y>�yƠ�k�)����_]�9��z���t�K�s:md����<n�}��tܑ�pF�;��U90sгK���		�^�e��5��Vv{��$x����{�Я&E��z{����$)nAy0�߇M��h��S� D8 �w�b�7�6n%��օ�	���80nLidy�:�N�AL žw굾r�i}�i���$�m��������UB�V�P�m+-,VֶҒ�YD��hŒ��,��[V���Ukkb0��m`�mKD��,DP�� �ڌ
ƥ`��j�,P�-�@Qcm��IYb�-e[KZF2����U*������PYiE,XVB���Q@QPX� T��F�(�jJ����Z�2�X��+(ł�R�E�K(�++QE��,���R�,�iX(,�["�[J��*��Q�UAT�Y�T*5���VE�V(�X�X��P���"$���#*�
�VV�aZ��U�B�+QV(6��l�a���)b�h"�B��
(�B�[`�e-"��b�2Q�EU+(ԇ��/$����&:$���ݻ#���P�����+ʽ��/����'��N���n��Ē:9��t/E+����=����A)���J8�jAEl��g�:����R���G�{�7���h��LB�����B�Lр�#ND���mlv�y�� \{:x�u�zs`�`�mby�۸���M��,)]�K/�A ���'���|-���7�k��Iw�lY��x�h���H���L��0���Y���q�$����A=�(�|��鄑.Wn�'���D�ADdR������ئPg�G.=��J����lb�xH����`�OG1Q?h�F�ߔL��u�'�3�����n�H��*$˧<�jCy�t/s雍�����7&�z`�-�u�b���F^ʈ~`�p
ʦ�X{U���U����D�{I@v��|J'���W� �V��:�8�r)�e��_� �l��C�5{.!Oo���{�w�?�������ӝ���C~ʤ
 ����9�27�C� qۏ6�9;	�A鶽Rq�Y:���$���Q�Q(���|S��@#b�O�9w~(0{Ԫ���� >�Ǯ�p��q�XR�.wʁ%��/�_�zgz� �Sռ�*$��rg��@��W�X5��	'>rEE��S�)��$��2ﷸ[�ۭ!뜨H�r�O޽8<I�|��ȥ���}���>�Q{�`痽_2I7��P$
���V���Ů� \uj��C�����CS�:��vݒ�^�L��T	�~�@�9X�~+w���4�}�@�oJ^S�k���=G�/@FQw:;���Ξ��C�_�ǰT�m&����,m�����TJ�,�fʒy#/�^�d��x}��C�|��"~%���lc�=�Bݶ5�Or8��M�vD~v۶�t���۷���<�v�0�d�n\�Z�q�!=�
�.뇲v1�&�����q��[��ۓ�T6Gx�=�/7A�j{F�ш�mn˒ެ`�GG ��%v������I�u��h�lf��\:x]��
Í�S�:�c��me.73�@z���u��&�]%[-��-n��In��v8��uїg�+��Ϟ��s���tN�e�����Y��O�˛�~vhl�k�	�	]��`�=���%g��_�k�rx����Օ�PJj:�*%_4ᯊu�bɆ^�je3�W�[V怈$�tOĂ�{n��Z�v��N�g^]��q6�l��Z�z�HwvݐA>�=��!�%��ъ�x\(J���ڇS� &|䊾/��U�6�Ewh��r�T~Wٵ	�Q�y*��=��3�Ey�*'o�b�$a2)c���	;X��5��ݛ{���{J���	�u�&�_t�@�^���!$�5qV���8��v�����\�sùݮ�]��B���ܽ���77w�<!j��Q0)�u�]f0@�m� ��Qh.8�z�^ϔ�C��� �wy��qk�jhEML�LM9d��j�3|g�����{w�Q�vb\6���\Sw< A�޽!<&8�l^w���L�.{�rzo(�cl����o�)�+	;v��ͳ�` �֛�":�iE���	sX�S��֝],���8�*%_4�+�'7�f��f�E��3��炇SN�` OgX�l$�L�|����P�nE
��K�:���fCz�%ﲰ�	/�C�v� #���cͨ!�$���+��l>���z�bH	�����2ʹE��.5�\�����M�>*v�`$��_3��{�Qt�w��?��v��9Ւ�GGl]s�5�����f���|]D�c3����#P����P��)_�@ ��������Gm{��6��4��r�ij�U!;@�#H9.Z�3�'&P��I���
��>Ꜵ_� �W�dD'sO���\Ju�Уڨv�"f9ɗ-�O��(4JK��U	-��(<Q��:+�/n��!˽Gé�<��v��w&�S�4a��;��vQW��j*\�51WvY6���'� �6�a�z6>#&�*
�>�i��/eڝ�>Z�戋A��W$@ɼ-��D�u�5�ޥ^�6��t�g��TD�ĸdl�l�u��RO����g7}�5�թ^����- ��� 	�暵i�9�����(C��ۍ���;<��1Ӟ�+��&���g�h��dm���?>��%Ҙ����l�W$@�x\4 ���z�ՀVZ��Z-��|6c�#�E}�����{�-[A�o�(�MF[�n��� t�� ��i����w[n63���Df�b��B2���|�ʎ�	<Ϋ��),��6.�����F��#roK� N�4Ů0n�#b9ɗ)��?/P��������s�̈N�� .��[��M��ֻ�>�����j�9�k��[������_>�cpd�˧���zΝKF���c���#���Ղ�Y�����{+}e��ru̸r?\-B�椳$��Y�Iu-��M���w޲/՘*�
��-�@Of��PI9�_%�������H^pD�r��.�ݹ�{]�5��y�����;OjC/��:hm����24�26T9�d�W�I$���1 �R- ��ѩǷ;f5�s�3�E|/ٴ,ZB���,$�fH��ON��C��sCQ`=�ض�H�v��
�r@$��3➝ϧ��澽]k/">1#	C1������(b �'"�� R��w���ySg��δ��鬂�J�"(4�،�$�aWL�UT��W�9�*�`/��p�l��`|wU�^kNn.��>$�u�b��0�p�"���M9h���ޛ�EL{SudJje=�i�VMd� �|6`���z�tf�8K��UE<$�E�e������m��pC������������k*�U��.�둯|q~�n|���sïu��ۥfw4]:1�ʣn����Na��ch��m#�����qnHX}��n�t�v�y���۶��ܼ���7"��9�3\;K��8����0n=�WW[��h�t.�n68�y-�A[�gF�Np
��5��ڠ^z܆���]<v3�G4mF�8��i��/a���#�iL.�.틫`�L8M�z7]\.�&2q!EY��q�u�]&��V+���A�on1mKCne��-�g|����G�I��N^՛I$�'ƚ$����@k��or2�9���֛ ���4�hk�XB	n*��I|�*9�cε���_zմ�
�=���d�����kk3���V�Ÿ	Q$J����º�gM���
�v�
Uwb��@)魂� �+��������fJ'�}L���w9���i�2������.ڼH���;�'�b������C5�*�K��&2��d�,]3�K�	�m����"=T��[�=�x?� ��i�8e�ڕZ�Y����v9�Ƽ���;j&����9�b�;YeNt�Uvic�	!j4%_��p�"���sϖE=XDg���h��i���ŕu��'�231WMd �����B\��1��RQ����Y��ZR�E�j�8��� ���g�����E��G^�#Ԉ�:���w��N?��=��[쿍Ŵ���]��d��9 ڼ	��,Z$��yq2ɞ�+B^S��7��Z�/U�i�O;�ͤ��f���ڛ�X�"M�Wh����j^�,�h�2EV�4���Ɛț���0 �3�m�z�Ȯ�ݜ�b έѤ�ͥ>(!WҪ����>�C;3�[�I�7�n��^���@ 9���� ꩉW�{����!���% II�V!b��%65�zm�h��2�G��5��I��λ���q�Е��$��*�خ�$�ݫ6JI�bT����J��J�D�a?vػ\oK�$�7͗)�O��P$���h&�#�8�� �sM�t�&��L���xY�ol�<��X-Y�i�m���E%	=�P�	$�7�	}g��m5�(ݎ�Rk�w�����[�7c0ʑ"&j��Z���V��c}茟�����O�m�{;jzo��_n1���ym���Y�D����_։+�bD��3��$-�\l�l�uȏ6�e��}����	f�U�h$`[UX� 7�����Ǜ9Q_ o6ՋR�Ga(�)8!r*��*��RY�]=�=?w铩>�����~��@$I�u��w��{=3�Sh��_0a⽸�y�䋫��R�)��u&���m��1�݁�&B��	��B�$���@ ;��l4����ˌ���6|uki�@��UpX
�qD0��"j�2���$��̼p:�]�P��uUh_�|�W�L���]{���	컱���kX��6\�a?G�_4I=�Z��	 >�wG%y��t���jg�� �x68�[m���H�	>�Q��u��"���K5�T�$��eb�	�~Y�}d[���6�����k��v{�����~Xf�̨�6٣�����<�_?]S5��:g=��\=�����S�G|U]�`��3��$-�\l�n��/U	 �M�W���[��=�{&� vU��H-��(��{��n��"�ୃb0۫��[���\�_`�z N�8��q�w��4�0���ATg|m�Qh �.��Zl�L=�����;��A4��W*7���0�d
jK��=��-Ug1z��B�:�ig� 7j�o���i� ��{*�_qu,�g���������(�r\��fb���ev�P��^��ܺȜ[T�Γ��D�^�� ��i��qf�JpF���%�
yz���^S�o�D�<e� �V�N!�Ꜵ_����^�r$��+�-*\�;���H��)���HFҹ+���Ш���<�䶖��{�a��=��ߠIOu	C��J�	C%	C҄��BP��J�%j���P�=�%*��BP�BP�(J%J��	Cʄ��BP�BP�BP�����)��ͼ��]G��9,����������0�?�L   �       �  ��   � .���( P�h�  Cl�(�����J(Ѡs�H)UP(H��
B�A@�TQ  $i�AJ��P@��X�7Z�3����d��A�6z��dyj���N��E�{oX������lTR\}�!=i���˹U�*�U�^�ڃ��P{j]4"��\*�P��O��Q*�Q*|�X�G���5��OA�'���=�LW�8��=|��:�Ӡ'�gAE����@�)I=��ђJ �>�>�CCZ+��/{��d z��_a�: �:\t������E� �	�A9�s��o�3�t���hzz=q�(��^
QT� ��DQ%IB�}ꠊ:�zeٻ2:��g����� �jzu�Q���zӋ�$���>�ȕT��]�M���mQseg���N��m�bW�׻���-����$�*T�T|��`�:s����;�:��睪�:bt`�=+��iu�)l/��ϭW�*���=�:eS����=�W�=t{j%��+�*�      5<@))J �d� 14�2a4"��	)T��       ?&�� �@a M  i�H�I5@      S�L��*UG�ɓ!��L&��4��&� )#Bi�!�=���S�ި�=M4���G��/���>ϳ������q���$������P��B ��%�@�>�H Hk����2B 䃟=������?��:��w�� ��`a @ aD�� �!�`�$�� H $>��žk?4����������P�  u�I8����\����h�H>Rd�9��T�?��o<������J����?�$�S5qs2�L�Fe�jZ�w)E�IyR��M	�f�t�+ �K4�`�u��҈�-���㌐�;��̼GK�<�rv���ᢩ�毹��<�6v]�Z��x�o��&c�n��lIl�e=�[H7�F��m�/J�1�+J��hB
���\�nke�m��:����օE:�w\��'�>[�7�����I�Ć�tIf��۳*"�/q=��U��y�Xn;���l��Z��wp.���g�qx0@W���.Е�\E�{���m��6�`�2��{�o(��W�]]�y;����;�ݱo���0W��ż3���ΰiلt�V�*�wv���qi�ӧ�*��2�0�Ƈ^Ͱ�tT�ˮ��N�rjW>�mc]�8�΀.ێm�O�;��C���vb�]u�M}�e������Gl��kJ��D�q�&���wLX9�v5x�����ۥ��m���z��o7�X��9�|N����;\��h��t��Vo' �e����-�Dz7x�=�;�Y���-=��;��Ax՝�s�|���v2���t%����Hu��������$	ܵe�T
Z��,^��Q\�-G��%����w�E��vRd���`ż����tbא���[�vL|��\�a,�x��Iw;)L9fô�����%�u���,FA�!އ�ɪ�̳���`BX�.j4g_��]�4�|4߸s�"&�=yѫ��;�'� ��N��:�Mb����P]�T%[ >(���N�-|��nfF�MŰ�o�����u鶾׻D�s*=ٹ1E��当4G�`�e���׼&�_�0 ���tBݫ/S�,9�VA]�x���)������%�N�ΐ-DI��_-�	k��P�#��qwN	�B�&�����vsج<�{1�p3��<��+K����Ö ��ל%�ʎݐ+V:�n2m���'7^�Cm׸؊P(��w���ġ�]��.��_Y;��S�K����/��,d
���UUچsV���	M���7MU��te�5�)��xt��/v�� �M���w�ߐXȇbi�t��q�t�v�.ר�(4�N.��{@�~ߢ멩a�^�5�`'�r���G)�W<(�[�q�=���Jfe,4�X����wqH�;��[���ED�)�M8���6)o/��9Z�%�@`���]�z�r�	��Xh�IN4�����wqq
�*�ɭݵ��-'[���}xj�F0u=�5����%h�;�-Ӷsah'��лwxt?ndexw&�f���O8��0��d:����Q�!D���s�ˑj�Um��Ν�8��5�ڮ�kہ��9����n;OW�8/מh@s�F�79eq�.��t���I�xv�F�p�$Ij睠�\����5����
9��V�:#0�>6���(n�y��U�nt������5ۗ��-� ��N�NL�/��䃎��VZFp<��;�Yz�wrWC���.\TTӳ{j��@!j(B�B��;#79wq��޳�0�rݚ
�Ǻm�z��u��{lR<����3���΀�k-��<�#�C$q�q=�(��nL�gHN�rXƒ4��t�nj��X�d緤�d�4k���;��:|�<�_TS��i=ʅ{XG�+J���N碓z�뱾4� e��sz�咅��=^k^��
�G��� q�JKi��N�d�9v ��k	�������{���W	&�Aۇ%��rZ�����֞H�d����$�Y4�����v�D��	�I�]X�]�t�?J89�v-8�I�����n"7���9_(��i;z��v��l#�K�����T��jh�,+�53�lKL��f8wr�b�n���5�ݸn�}P�"-�Ǹ��Ԡ|v|N�Q���)��a3R����k���БѠ���g"�e������)*���h��;fܝklN;d�JM�g��ǩ���n��;.0�v�A����.m����nl�cN������%��q͓Fjmٯ�wV(yb�Mj��q��6S��qQ��tu�`��ŧFr(5�PW�βH�g{Jc��;a9��=�ҵ��<v��j)��>Nt�m��Y3z�9D�M�&�b�Z��q)vǤ�齓s[���;/2�r�Fq��:LX8�{��7T�Ǩ���~���N����GXr��[ßN����{w�nuC���q����p� }z�����(�2���T���\yAٹՁ%����C�y>P��7��7waB�Ƚx𓥸Q艏	+��y+ZMBv�'u�f��7�?䛗��ʙ���	���uk�7��r���H4�"Ž�@g3��B���Bwy����lǫq̅�Oj�v�AΜ�������磩(��L�'�%��K�;�:Ocy�"顥R�\{�t�\�Fw!��@X�x?{ާ���d��}��b#,�2��wj�٠�r��^�{٫nWb�HE.����Ihڏwd�EةFex\]��2�13�v�[xt��枛�l)^w�6S��N��bݺw�؜Fc�^]��zM�O.���S��fVC��w9��q9�&`K] -
n�{��z���4!y#L<�[�����IP���:v%�*vN�	hn�{�J��ٰ�F�Zt _\]܍�q �����}��Hծ���U/	������� �T��aҮ8]ѩ���=�r�Rm�����1'���;Bw���LE�7q�;v@�lN�v�fg0�*����k ��FuQ�ip��2��1{���a�wW�Jª�E�V��٣55ܡ���UQ�/�Bs
x��FD��r�Wgh���}�F�]�f���.D($�oƜܮ$37Q!	i��̭q��D��$l�q�r�Q���\�7t��.���� �w/�`jn�:������:�P�)v��ru�����8{Aw}���{5n1pM�8���u�8��)���������FP������6EF,�C���v��.AVn40��㔗5c;{���˚��p���������q}%�%�:W_�^%�ȳ�	�{ݜc��Cz����NC�l<VC�^�5wwZ#�q�:-�8�tۻ��U\׋`]��9�Aℛ�m���h��P<�o[���m͕0���]d�n���k,���a\���L=y���Cť�C*���a����72ky�seW #T�Z�*S�^X��#�pta.,Z��MI]v!5�o2{7al����Vv��,wvQ�{P�Qj{w:�I�f�ı��S$oDUCDo���i����m�돨����E����gns��̽c��n��ȝ�ѐ&_Q��'�����!	h�ٽܤd��#�S,!���6����K+]�8ճ�5���n-�����20ڑ���0v�x�=Ģ�͝��M�N�	,�6ѽFWp��óK;Á���3sV���9�S�U'7�4�A��t1�D�]�״���8�֦x�c��/9�N�C����	Y�}�)�_�:�N`�̟jI��f|x�A9�W<Ӎ�G���'�ts;BC�aOڐ
� �H
AI I"² �VH"���XH$�T�A` )d�(I�	Y T�P!"��"�II!��"� �I*HJ� $d�P�@�$XBP� �$"��d �I)$� J�$ Aa
�B����
B�$�T!R�� �B�}_��~����}7���|��#�$! ���͒H |��!	>�;�V�O�R  ~c����Ϸ/����S5�7�eӺ�Q���`W������HboT�S��;�U��J"�����΢)���zq�}��
��� �>z���T�&N��Үk���˕l쮚��ރ�c��M�����H듞�{{LC{GoH��6d���
�+�X�H-����C�6XH�%��7�"�Nb֪�՗��ǈ]e��R س!Y���F ���xGA�w��qG�*=�ۉ]"I�{�<�E�:�x�i:g�`�Z۾#�rz�w$Ŭ���ad��+82��wm, �7�őˀΛ����v�.�\2٩����f|�F;@Ci
�y%EK&�)aS^�º����E:v���d�fW������x�-�X�p���m{������ۗrk�'��*��9���?w��J�c~�������z���p� ֹ���d���n{/sGF�Vr�s_{|�;�R�g����x��[���mz2q� �,{����z��Ջ|�����)�t�s3E��IDndV�{�u�kL����0�hC�Y�:�����.G�����ɼ�Ol�h�9��?iLkwR�y��a�08y�U�.����g�μG��]}ش���k�o�&��c�0��`}�7���_<w��o����o�"�Z�$�/�s�p8�A�f����PV{H2u��,;��ul�EՕ��Y�������[���v�'o������G�9{�.��V;�e��q��(�v��(�g���ڟot"m�~.�
\Y��2ώ9}������9Lw��3t�q�^��V�
e���hT���R��Q��oi��R��&A�_8��g�LWg9^���OgV�[��6��������gz��{��4z{\,c��\B�O7��u�E��d�A��n��#h�9����*��q���|sGf�&�=U`_M��>�q�t�@�Er�k��:�	�.��Y�ă�3������Gw{�#TX�T5K���k-�8�T�:�z��[�[QQ�4�wڞ똁�q<Z����m'tv��fXw���So��JZ��O�ؽ6���+N*y����R2�/T�ŎgZ�G{�R{�D��U��^s�*Ɗ�`jW2��g[��~ʇjslD	Tm�u$�u$���N��]��>`C$�]&S۽��t��=a:R�G����j��l���O���7@���W妐����U��:��x51�…���6�(՚�Y0I�F���eU��� �O�(dL╗{xd��h0r�3����	`�,��A��STsRk �J��FlV~��s>�q�;w���W)���f�b�^���y��=���-4��{V�\X�W�����sۑtі^��'�ӊ���|=���o!�o�Y�t�N� �X��bY�{��`�s���G����ܳd�p�:�zw�y=�??:1��c���h�Nm���䕝ў�{�E��,.��a��ށ�vx�otf�Wvh��y���4�Ax>}�,/�0W�1�����{ވߜ�)�S���*��&{��^����v]Ts�޲��f�-�S{�/x���໔qo+��Sf#!��os1�v������g����ҍ�%��땀^�}�3ڲ���Q�5_v�=�\�RΛ�W�V��w��瞽���s��3.w�xa����u�Z��sA�=m�s���u�#��}���pS%nn�A鎽ݺ���h����gw�<£/f��}zѫN\�PK�j!�||'!�f�̞�>rA��TE�>��A��;V8K�봱���䛞��f��c�d�!Ы�c�4�5y���&�=뒅��j��ˋn!�k;%R�W������ה#������Z�ŸM��~�s�S��o�U㫇��ks"׾7��]+�A��h�ވb�ș�ϖAiy�V�n�I��ų�j�=�Pߍ�����Ng���M�	�/{���KF�U���~L�q���=�E���Ay馷yݛ�}�1������������.jg�>�Ć�'[��N��9/K���K�w�(e��wn:�=�[ͱ�Wo���4f�nv^�	��Ds�Z���|�`�b�i�}���T>٪��g�>���d�կ�}^s��4�����Q�'u�Oz"�{�;t���e��/�#��چ̎�`�Ɯ�>zYޒ1�İ� �}�Oi�FL���_slz缹Y��]9�8�#��VI�)�g*+)��S�Q�u��>T���h��,�8>�pɾ.dȈ>�_���1Q������t�s�l�_k�܌mz�/=o��.��6�}����l9f�Þ<`!d�F���e�C !1��b)6��.`lƦFI]I�.���U�d� OՆ�E��igv�?@k�0��g��ޞߚ��֬�-	GH�T�;����"l���}��{��g/U4`]���'�sN����Y�ҧ�/S�a�d;w�s��zG�;�p|���z(ܚ�c�z�S���^�Ί�q��Z�)�Ȭ�{�4�6b�����͞��.
�.�3rn�4@��	�L�}H�{&�;����t��H�8�)����ד\�]�a�x盝�4��o,��{�6�i���{��\���4R�\�Dڞ�o���4c^���v�T;��-j�
������Uk�M��^���.��+~��0$��6�[W,}���s��XBA��Ǿټ`���i�29�<F��L��b�;{5��2A�����Ȟ�Z4��s:�����������}����B��z@p�ɷ}�z�zؚkk]O�����ۋ�=�#5������N˿C�#M�+�L[���r涶N/,��2��6^4jp��<�����?v����+�w}s�"�8��&�n�y���}.t�&w#R���*d��uGUz�j�V�ۛy���A�d��:�R��ᨹ٨,���;ٶ.=nr����N�;|����2�)��/6p�ׯ!�{����ZYU��'2�t涵�9L�ؘ��~j��[�=z�!�r6���1�\��B��Ȱ�dAx�E�;�Nkʇ/��ygv�͵��J�x��.��h�Y[s�HK�����4�i�+M�Z��d�8�x����Bv�ۛ���i�`w�����*@���ZV4�M͓�E՚�w���'����ھ5�fq�nC|�{MC������!�{��;c�yo�;��A�?��}|�I��}��1��M�cxtl��ys�&nѹ8bj<�HC�ﵬ�c ���z��t�1I&�[��kS��=���k���F�Rnwa6��y���ăRe�&�6����0�B���x���zu4���._nn��B��c���Os��׻���V��k5 ���N:ӻ$�盹�鹹\eY`˾���]OǤ9b`{���yf�����Vk����^,���ǃ>}�~�/f�P_X��4S�w>�v��|���0uȪV��6u}.i�$��}M�Ot����x�̰�2A/7���5�=�o�c��8W���x��.BO �U#O��I�5^-�0��."�wM&�JHֈ��=�����{�Z��8�/%��>�z���gp(\��|vM�9����˽���3|ߐ���]_jW7��.꺭��~�p���r������5��]>E�>|�u�&t�k(����wN�U��φ�#<����ƹ9���m�n�x��>A @ A���@�tA`Q����{;0�9������nB�af�����I��p<X�s#[��%��4�a�a�<J�Q�ձ�!q�u�1'i�n�9qjyN�U:`���&�i�% �+s�D=j�Vwo3�v�ue��`5 /OO;��ض����9A�Z��܍�j$F��f�AJ�����웴��[i����x�F�m'mҺ�^�\�̺�CJ�f��Z��S
ku��U4slMUXb�3e4V���p���-M��鲞j]u����w�mn��`%�P,`e8UZ�ҁ�<�e|f�^@��A����.ی��R�Fv��Aڼͳz��.�s���Ʀ��D#[n����x41��0iFJͳی[��.0�P��]��4U���nGYt4���s]A%�l`��6�#���5����$�q�u+xp����xnӸ�9��omtܔ�]�
ɆX8� Q�,E��)�D��1GO�c,V2�z=��v��NB�	[]	�rm�sc�mw3������Iw6�.���ظ�%�>A�V���ͺIڍc���Ĳ�K�b��m�QyI�Ll�H�<�ivf��ʐ!t�Yy��ڭ���Z<�]�I���9��<7�;kɺ���{�f·0�:9+OE��a����mt<�\ö3pf:\�b���fA��냬Z��\��W>�lu]���`������䱙R3h뵆
�xR������R�4�6�۟.8�j#�Z�1��J�[��fi�h�=�(�k�q��B��nL�f6d��mf�5�h, c<�^Es�h����o<�XT��0̺V˶�Z���	QĚupÆ[�Ѧ���0J�5ܡ�0�.��n-%Y��X�\]e�h��X�9TѰ�.���kn�RY{6�B�̗(Ʈc�p�w&��f�.GW��v.oF�;v��E˴$�]b^�ְC0�M�`�ݪ��t�qM��8��6G��m� ;G%΅̨�ƙ��;y�#���W�3�sY5�݆r]t�[�oq�Ȳ���uώIy�=�;m�ݠИ�wJ����Z�S�;/=�hz��`�Z�Q��m�t>C��3�}d��bE�8�u4f�D��[�qf�1�
;qn��J����7W61���X�h�d���Ӗ#@����q���:�t)��>G;ݭq-�ƶ�� �]����r@�Y���h'/+V��X�An�8�2��n͌���Z2�$������Ú�}V�����8��p�]�ML6Հ�+� b��c�v;(r7\v��섣9ɹ��U�ě���#Ú�z�m�U���Iڻ<�;��ύ�n^�э{�<�M��z�{u��e��m[ʸ���15>;�x��^.���x�Us���Q��گSֺ7%�VJku/	ڭ&v��Dt;Xacd��X�&���H����kTk�yl�z�9��œFyjh���(�4��+�i�2�M`�Bgf��Euz��<�Ig�[6ݮ��[�P�.���8�1t�z�Ըw���۔-j����ܽ��%�aWO<�'X���
On���5�#�iL��OY��˥8t�l�M�<kX��J���t+�N�Z��7H�w6��N�Ax�M����sI�k�����rŀ�d��U��n$��ͭR5�.�qu�s6Zk��tu�#zm�WA.Z��B�y!!v���#4�z����:�L����Iny�]�ˡb�b�X+������][�]�$a�Z�;t{tl7Y���Ø���I��6Ɯ���!�]�i�=�3���e���\�t��j��Vk#^����5s����]�bӫ\�H���ؐ��VY�INT�`RE_R<�z:�E�9ڼ�Az���m�g�Sb��.]n���8T��Ϋ��Y�WV-%"��iwj���͸�<]+�.�H��/L=k)�\R��j�eM[���ģ�3M��r�s���:S�X�"�;Uۜ���{3��^/t6�nw��ZnxN-ʢ.��6���m�R.2��櫛V��@t&ڵ�m����VwN��+-ڹm�k��r1q�U�7r��0�rJ͗ia)��0�&n�Z]���\P�h��%֍�L���9�%h�c&�,+��G%ݭ�ی�D�	��#�9��
e�t��1��T�Ls.��ű���r.��M�5�ve�M��4ͯ5\���Z�/0p�cef�+f`֛9��ۙs�����aYn�lN0ݮr�h�eS	^�ĺ�7�����{
\<u�FW��^b�/gu�i�۝�����ٮ-�^x+�ALqku�$� ��`���`�0�l��q1�B��&��W���<*.�ދ�����mm�=+&�z�˩�\N����h�u�z�pζ�lWg�]7j��V�v����t]n:��qPuW�K��nmt�Rx��=���79�<Pgn�k�5v�Ū��������m�����[]�����UV�ԷD�T�V�\P^���2v�nGx^�u�UqU���9�I4�{�`pP�qj�hD����\lW��/4�nv��hJ�!��[	��L�96%mA�D�B��C�gk�׉�{��=���a�[W]�06^�n�GN}�f�]�z�5�����͹�ګ�j�)[��ͻ��+RlP��_����QJ�>2�{�-X*���TƳ�Y�cP��J(Ȧ%�T�����i��8L�+%H��.��@rbD @�"D�0����Lqej���
ř�k
�v�M+*R�%r�E84�$�蜒�x-%��2�Xu�u9$�����8:o�㨜-[-���6JI����J-IZ�ud�QmHf]1B�ˋ���FҥDb�[z^đ u8��C�RNcf�r^lA��;!���<3���5�n��tZ;Y{�{@��rYm�>tv��v����#�h��b3M32�d��LT��[�
gUv����/=T��{v�'��Y�v��x�3�ݮ3��������cX�y/c�̇v�x0-��nޝ�2�n;��y�Kنꭷ��[�Q�u<� ��Z�im�"���y�7eZ�rvw�u��ا����8� k�xnU�L�`��:�U�.�+�&�.���1vkg��F������qc,ks���U�\ݲS�#�����4z�tћ�X�#��Z�M�ɮe�8�)�ձ��#zah�
��	�k45$���f}��̍�t��7qr\��Y�Ԍl���`�����<���FZڙ�L물�ɦ�S4�s�)�v�D�D_WS�1ls�S\�&f����9[�Y|3gl%�+I���i�m�k	\�Ď%�^�~'�/7�F�;���0�&�v�ԩM�k�ϯ\끮�ta�1U��mU��΂�Ul����v��K�j[�;Sɍٵ�9a��.3�:CirYPU`	e-^cQN) Ee
E��l"��F�m/^V��+XKT���kly�[H6�c[h"W�eycy�(��)R5�4����T"��ce��-�.e�k���x{��;ֵ�[�kT��4��ou��J�eX�<���EfUK�Ov@̿`���%h`�����ڸ֫���X�!��3� 'ֹu��ڹ��#�cH>��3mWc*Z��S���e�|vz=ڙ�\`b0����Wj�6��=���x��7ǋՇ����widG��j��v7WC��(:�tHGl�F�`�v������'�/U����Q ��Vg\ � De@�8b"�5�?��3�B�|&TV@5CEj�]c�
wF]�,�ٻ�8�؞�k&c��ہ52��������(#�yR`�}8"�w��P��f֘5^x��3M��x�����kLQ;<��W�)�qWFT� g�$q�/�Vf�/���$�?;\Y����}W��n���I��k2�Z�IG��Gf�.x�s�e2E�,�]^�����A�L=�lCgS�8l����ۀL�dZX#�r��c���JZ�4<4 j�]x��Y�������pO�7a�w�j�Ǚ�p���sFm���
�r7ݚ�x�j��oa���]&�կo!$���9y��RV0��j��ßr�L�oK���+������f�*�s��گ����ԬsJj��e��)/nQj﵁h�iE��~�d2^�	��V$b]��4��Uj������?b�3n�V@����l.N��a֙"�����Ϳ��\>f�I嗄�:�������,�I;=	�uz�rl�3�3'h����.9�vo���\�׬H:��nM-��1o�	2���6��K}���O�0�3��ʴa�������T�Q0c��\�0�$c��$�M�X�����,��_��<Q��A쐤\4���&	;;�uݘq ��}�؂���sN�<����C�=蠀�6�����ʿi���l���Al�u�I�k&,�bd���<�g�Č��ǐxeY��j�_CE�������@����{Z`��h�Md�M�N�{f� |J�*�JD�F�7ʗ�}��q�>�܊s�0/e���(�����*�jS=�����4��m#��H�M���v��n=����,�FRz���'&�΃��ʾ6��ٹ�q��H\��u=����9j�Q��[S:��Pq����/����� eSdR7T���3oY8�[�Ƙ�>�`�_n�7�ug#X_i�\��A����[s��;��ya��7�o��N�s2r���x����_k�=�bIM�yq~8t%"�����G�~����+�b���j��gȜ=b1>x��Q��R��v�V	���for�\8�j�	M���Q2��Ω�6V�Ͽ��~j����H+�S��� �VEٸ�f&�͸"*�8|�l-Y��*k���jaH����"�)�DX����5O�p �� ���A�ۖ��B�0��)\X
��胲q�m_ݕ�@��3ܣ�		i�ɾ�Տ���� 7�p���A5�Y��f"���Gb9;kH��P���G��;N�w.<�չ�*=(�eMK��'�nl�{�U��/�!wi����pA�yĻͬ|r:��ѵ�T � �i�ī_Iѷ���y���$���d$hVk��΍�al��(��N�j���B�(�7qg]�̢^�����;"�c5XEZ��CE~�Wo9�[�H��q��.�3W����rAe�h8��2��ӟ!d���51����!Ox�z�=~J��=��ԍ��1L��n��-v������bo�R��)��xd[�w���̈/)��=`-�hr�9oq�H�~ÄI�S7R�^M�u�R�X��F �U����]���]6	$j�*˲��Q#b��(0��=�L;Z0�v̨P����˺��~����ߓ��,�3ym<s"~��N��
����#�޸�~�6�%kPKV��W��!�]�"j�ߦ�>�~��p��Gj�U�uq���(3��v�&����c;o�}���:N��i�a�����r�������,��I�H#���^����<0@gvD��ܷ���t���$� ��pO����T�H#T�3q�����Y�pL����÷b�0[Z2t�7��q=���j�u�a���/����=�SN	D����'6�1L�
�7w���f
����+J��9t6�T$�R�M4ܱ�Ō�s����㒱n���<�+�u���Z29)Ƅ�\��+I�Ճ�gda\Ŏ{F\2u�x�G�����M]n�qa��dcn&��j�ДӺ���ͮL�:��4�)Sm�`M]"���E�sE+��	j��/�ad����{-HG�9��K�3.�u)vMlF�Z���|)ˑ�o,�K�x߃*�W�Hp���n6a9=���, �Ơn6X� �����p���c\( +_��Ν�]�x��(p�)��4es�V���	��fU���=7��}��}9L��	��>qٌ��G*���S���ߣ����}�l@�����D(�@'�H���p�WI];�#��"������z5E�US��*j����(W���0�p�hG�I�ow���Ρ�-<� ��&N[8c�%�#�ֿ0-qbД�f"�ۭ=�D�d��H�EF� ��[Ft�7�'4��9���cF��AZfE$�j���=�w�쪈�UM2i���6�DvʫjWz��Q+��Ў|ѝ��b{����LYo!������7���O�\Y ��H�)w�nm�>��WV���;z������^���*����_�U�VV$-�3�n���<l{��Ƈ��n�;s�kl�y�B��V-�n���U:
��N���F��/|p��^ڇ/�C����{�����}Ӽ�ý��&������t�� ���u_�u�ω���Da-)�`�!�2��?j��r��w���a���gj�|��O-9�`�!�d��"�A<���.m����i!����(؅�eP;��Ɣ�x��yboq�^�5�ֺ̈́�B�G�}��\��O�>�]2}笽ѧ���'�'r�<)Y����έ����6�C�1�z�^��z"���Y�h����>=ܗȖ؋��~��+��:��o�M��D�~�^龙�R��s���Ʀce�иr��rF�^Ud�
"�*2�꼏p�{�^5h�ш�mm�Q�±dƪ,�q�J8�0�IE���"����;��pe�N����U�7��M%i�H�D1�)S�BMl��7�k�$�Q�p԰��	@��:��
�� -���R�B�!)�q�����u�����i"�V��R�UYJ��-�1X����Tm*�qiE�-nB�G.��*��+�"�Ea��h�(�p	�(Y[H�R�(6��UEaYEU���Z�n�TX��eU�m�E�Z�*J%���%�/A�X�KK-'��9l�Kz w��3+m�.X�1
�2Շ S��$���I���}J�"�EQ�����}F�A����W���=�THk��[�U
"������@���I�؄�g��]���[y�Ԃ�E8�E]1�;Pٰ�.���������D	�~��6��ZX$��Q��(��z4ϋq����C>��\�f����U0�
�L��Z�}����&�\���U�(������$R;��Pt��=V� �C�{��H�VlBma=JT���(CČQ�Ω᤺���*��{C��Ə�Ę�q�J�h8A��]��k��cũvvA�)ח,�Ԏ��v�H�
m�Ӕ��:dM�^�u~}�����5�}� �m�Ѡ���[���Q��P��2N�!�F&�*,�[�z�z�H�lz�1P��v�.�U�(������z�}�[��������R��us��W�8 h��xnUV�9��(���H��2+5��l��liis^�e�mz�����+5T����TLҊ:tx����t$l����[9�����ֶ��D8%�EF͘ͨ�a5T�:�Q�Ͳ�]�+up$�3V�\v�Վ�:���D+/b���l�ra	4�X�24���펜��̧8��.�-��Ӻ�l5E:�s��P3�H��ղ��Η6R=�ctܽ��<�S�����4=݊>>R�P�uQV��Qg�7`Auؕ��Kb���l�`������vpޛ�&�D�: ���𪥒_v.�ݮ^c��K�v&�hJȓ�B�\�Δ��Ά��Y1פ�qzS�M�ʦ̓+Hdl�oS:zn�O?��˘]SqWmq�V��SQ���T�me#uUJ��_u���W)}ò���UQwJ��8��dw#��+D!T6bn3�KjMklN�>�uWK�mܯa��B�fǕ� a!D��,��>��$�&FTO�R�m~s�NC�5�/cbSU��Nnǣ�5�rz��1U���k��U{��������Ɋ'�51Y
��(����� �o��W�"�� [Z&��r���hƈ�mG	��|���@t��6�)�Y��d�q>א��O+"v�gE(�~"e�-���
�s��A��ٓ��{3<�)t�=Zj�4�t���]+��:�����{��/6y��A=�����ˉA���1��RU��{��χ�zߟ�œ�_.�N �9?��+[����bG��blj��Ż���K���AiJ9q���e�r�'qnT��+nӊ:�`�#���emJ%x��.0 ^�FgE�ۙ���mX�^���H姽ả���=0����I;͂f�a&xĠ�1a(W+$���gq��;ͼ߀��?����U��|OU��4�G��l�v�����C�f)��
���@#Y��e�M>Pg_Sxiu�g�QoD���{��?����0�"�A
��N�D0	�23�ԟ�T�1�O
��b�J2�2$��zg;jw�yRoh�� �b/[2��i�O^�捨P�*!?cr�5��8I&�0E�&Z����r8'��I�}�A&��E�Q��4�����	��>����ˑ Ʀ	e20�d� �+f����Npj�2(=��R`�N�,��-`�Ѻ�.��:�E4�Z��/b�U<#3b������ݠ|b~Gg6f���l�l��X@���t�w��-��,ƭe�YaR���maT[�˻���f�S۶e���}�
.���s�,uɷO���lf,di���mm���S���j�*U�(��-�\��ƋW~�����]��o�`��Vxh���_�?��h=�qRo�K����̻��7[M���
D���T#
A|�'��	�:��f?�Vt���G.�7�����j��$���o�Z��mz%_�@H��..V�U�����@���ו�s���d�7AC��@ԊD�8��*#�ܛ}�U�D�o<��#!/u�8n����+<��:���{n����B�ٖ��{n��%K�_��v̷lr*>��q�5������E����_�� ��2F�>`���މ�~^'v_]��CyC�8t�� �UW�|̛>�l�щZ�^HfG|@t��!��.��]o�����V�y�I�8�/v����K&�32�7hD�˂8.�1lĆ��f3��V�1Z���z�OՇ�	G����M�|¯��0l�7S��*��l�*S�Յ���$���>�ś{K��h���E9�cM��$(�p�O5����r4<����Е�v+��l�i[���9V�y�"�}� Z}���Ϲ���iݢ�L�s,�����>ńҸB�W��9J�(F*̔���{�����{i�3i�N����L�1��%%T�(ЪJ��)��%I.��I�r��͂��LwP�B|H�cH��(:E����iX-��ӣB�����.멜��U�(v���F�4�>+����K��6������tS�O*v?�������=���ud�P�#\ش��]�&��J͋Sd7gʜ+0�-l����g�N6oƐ-�.>��+Z���A5-�,�F[���{�z?N�%(t�0Õ��^H�r�mJ�w����ă'K ����T�˘뀁J��a:�$�ql��E��� �e}J?]�w���-�H媩P��|^����Tkt��a���}�V��U>X��c����uLlB�r)GNSS-1�2�#)�.�N ɍo��~6랴�#�xc� �@^d���u�s��|j�Jz�/f��V)�P^����׎9����ɴ�%rg����u�5q�g	�MW�m���t�WjK�;| w���p�e���So��TR��X��Q�^~7u��c_,^~�.��o��^������H�~����Z*	s�1|�D_b�x�׷"sKm+YWQ)
ImK�
�X�3�������:߼�ɔ����8/�3��`���=۾ܶꙥ��G��Q����<����t��'�t �B�sŕ�m�D�d�vM�gsĝ#x1�,
���+���ߐ��KM�V��z�z��p�>�A�xx^���L群5�`�E��e� A���]<`�3�N�;���x��7�{�i[�����ތ��� S�����~`lIS�i��D��5���<�b�e��*�ƒ.�άz�}8��?�'��؊(�^pR���XZ��� YzT��'R � ?o���x�+X�NNj��ȇ��q�&R�J�V��(���9K��-�1ƅ-R�E�ԥ�![�@ܔ��^�-aIR�Rrޢt�%�[pD@:R@�qo+Km� �M�5 ��0��%�D�6��(�$aBD���V�H�I�;�t��7�E�$�cաZ��� HR�� �s�fS̠V�ش!$D�8�m��!o��}V~m�����iF]>�X�YG���轵�,n@��Ѣ�V[�7=A�{sx�;���1����Z�hb�
�^����4���ۤ�.��n�]�3V�	��2��nX̬X�m�.٬��u�jX �l�x���6�rV�N�X��ۀ�@����{�椂/���.y݁ޮyF����EՃf&"�f�iID�\!l�`v�T4[m�Za��T�p3�4`9�U��v#���̣Cp�U6���]����;\i���:��n��:b�������a\�/a{9��f�z� Xh��꥘�ҥbv��sQΖ�O����αX�X��s��볡�#�u��A\j���
�[lf�<�e�l68����ע[�u��W�	���.x�-RGm$v�(���S�9����'`m������g�.n{c�	];ZM�.�玝u�� T��En��
�:��$#�:�ڪ��.�u�ĵկoF�g7[�MUUMV�l�+r�A���n�:��*JX�"�jEu�#�Z���,�	�$� �� �k�h������@��׮�c1g�x�P��7[��V�Q�es�2zޝɛqZ�Ox�P��N���ps'�ͭ���òh1r�H!�ݵ�.ۗ[.�Ӷ��֫�����c[Qƭ�3`85[Y��m"7����"�L��}����;7��Q���	?kg^fT#oC�Ëڝ�g� ��h��-���{,a���H��=I��q4�D!��grCH��)��B�d��~�����T ��eho �4\�G��`�Է-�9_I��!m`�I��)�q��M]��*Bݣ��e��M]���~����� 72A������Y�����	����"댟}��;��������fg�r"fl0��dMl���L&�n����x�^�e\@$��H`��&�O�ea)�+��?��ω�߶�	��uig�0�<p�h���L��N���G,~�#���@��f9��<#����v���|��Da	t$�8�暐;Rm��Q	�E��=��Q��2󽻌_!"�����LZ�~���:E8��^��ws
sb��n���WǛ]��$��7:�	���p��������� Ͱ�7��!�hŇ�Y�gT���o�� <����׼�!jͦ�N����9���f�չw�ݐ��ڤ[��z'/{:�����u�.u�P�����w��4\Z]`�T6�Ӝ!��'��=�(�wh�ku�Վ.ois��
Yy{�Tz�ܘ��<���N@2��&�{���"ro��g�bd�ݢ�v��[)P��Y��o�W��m����2VK/�6�LFvc�
5[ܩUOD�l�����s�b~\�1��w�W-n91��1孝�Q�#DQ6������7��&�;+����>_��1�z'��jK�����O܇ v�Q"c�z)����u��cf��l	�KGD(e��a�[������c��I'>ڜ΄�s�oݛ+an�� c�dC�$��}7�䣅ԇ�\�s�6m�qw	�<9S!	XY꼟Yd�*sr���d��UtN�k!U���ύE�h9Q�i�wN�'����3�����moV�р[e��J-U��L�"豫.6-i+J�cKf2[@wG�WWN4ì� ��c�sH��7it�ъ+�[��\�����Z�Ӧ�9��.�wnW�m��t�+�����7��h�����@�|���`n���O���g^�>�.��u)S��=մ��sQ�m�b�EU=�ܰ/����aʍ�����;�+z9҅�ζ�I'=Kû,c�7V�,��Srn뫖A�Pn�#��n�i��3)�/�i�ӈe���V*����"r���N�;�WAF��DotTĂ��,r�����H�%��V�3y���b��*?�xg��e����LyG$~�֧����z�.6+ш��1��Q~s�r�V�ׄn���8�C�5��΄�=���ݏ�eOi�/�@ts��r�C�<r�A"M�RF`5�B�lQ޽}��|����n���2�a��Iz7_X��N�}�qު:z�����5&0U,�D�:M��a��o��^?�w"������s�N��ޑ��?/o_�e^�<ۍc�j���H>SG����	�~ϵ���O�:ueU�8X�1�v���#]�(j,�
2��U��2��{��[�L�aמ����R�+�:��vڹ�h�W���t7� ��f0/���l�����)f�q�;�ŝ}�;��i�PV�� ���ۜ�B�0;bF�f-F�;P�N�g�)W����.ܸCgx�
��X`�t�"|LV]�
�#˹����x]�q_4�E���Dj�x'"&ji����� D��J!4[���pFH��lǚ,4�b��8�Z��=
J���c�u�R����=�3���p�z���
Y�\FM{�������M/_s� �옝�ft�Qᗬ�����ՏQ��'���ڝ�74��GrF.�]P�,���7a0��W�Kƫ�Q4(�l.;�qE����ӿ[����$��W��}k�#7Ex�Sl[�lI��ºС�
JŠ�Fh��-��0��Km��Km�l9z<1AήB�7AY�N)����9��.�Ӱb�a���u�ݲm��J�Nu�W�m�r�v꺏G[����mISW����>�w��{��)h�x����P�Is����{�b�3S��%������!��fc��C4���mm�)�P��3�)(�P�lv��JzLf�ίH�4s((��wln��ƔB�o���S9�#A��6�e4�]\�����07������󊶞A���Kyݲ��2�.s��e��=�s��\
޼1BDC��b�I��˸�^י&�����7��5��)}vk��aJ%α��(�9b����w7/E@�C1�E�v��!���ה�ui��H�0�d)f�q�ۓ��y�[�e
��Z�f<}���6fX!���f]r͏l�V���NS�c�uNH}���[��*W#���b}�^�2�s�r^3���97==�/Z{ ���u�~��0"��
�#Gn�FN;��c��`y�l��4���+�9vyg�m�J���L9�Ξ��������l��W�W�j�t֗��e׬���!.���y��1��^�X�5/�{��?�+gy=C�h�&Uø�_g$�}^�6h}��h~Q�ݝ�^F� �4{�RB��#�����9�O<������ޚE�5�����G���;���,?z8mi���ͭ���Ǟ����2=���T�}�\�F�d[��ϴ�ݶ�J�y����Ns�"'||��O�#}��^��i�m%��'���s�'F�����'�?Dk���q�I�{��E��Ί$�a`�v�p�61�Y�����B�5R5��i[l�DĴ4ܬ��qf[�06N?f�oM�4Q����k� ���Z&$[���2�mF�FdDX�������O��f*.5�[�h�V	l�*/l�f�,��]�"��t�[UE�����c�	��-�1C-$Td�eAb�
�"(�W[�C-R#j�8�"+ �k"���M�V"��
"�X#X(QkE�eUQU"0M�����(*�EDPX�b
�(�FF"�j�&5Pb"0APQ�b�X�(�J��EPQ�c�f�TĢ,b/�I |{�|!�ϟ�aAW��K�����c3'�X�ZEH�C1����*�=�~\�K�=痆���	���C���T��IR�EG!�U�D�%�Q����}����n��;�o�*)�'7m䛪�،�31�v�dɝ���h@��3����v�޺�{��O �H[u����X�ʒ ��
���Z�ϋ$�A,f,�	yW��K�+3T�(�����{� z2X�e�R�{^�LR��l�̐E�*a��)ba�6`�Bh��N�&��������������c����h�MM�&�0�2�6l�6��*��f/q�խ�rl	'���Xѹ�U�׽6�V���k�S�$�u��{k��r&K��Aq+�O8.�9v���ۘ��6��T��s<��#<��1�����<���#�;'��UH�u������_�Aw%�b;�r��#d�d�n\5v7'd��J଱�Y��n���PF�e�c�S��y#<�+y��j	1��)����u��fvu���.�b��8��(�ˮ:����UX1�[mN�鞒��e4D@0�^�P]�(�c��]��oe����\�W	#D9
y� �W��9�o1T��
�:�q�9K���+��쌤=������cv������v0;����I�O��=Uވ�:��Owl���7�o�!횚,v/��^w]Ar�7UM6�7��?�q����J��1k�
���B5�MAp�hׄ�g�+���S��n���1�`#]5$�����٥q�P^�� � G}��S�n�_f���T(C1t�<0m��������r��;R�����s{�����~݃!$�̫���N3�z#�������[����	1	0`C�&װ�kj¹v��{�_����V��*,�ރ�7�l^�g"!���Y�����r"����ܕ���{Cmg���U��&*��l�E�[��Έ��Yε)�e��9���1��c5��{����9o��$��4�2�*�>�����t�tU�,�5�\	M*$t�g[��{w��b�^�۪ޮ�n���"����*T�A����pbp�m�_i��zLvu��^�MU\n���y[�`D��a�ee���J��.�N�ͩ����D7*'�W7�.��qaAu���%��$�F�/����ؿ	�m.���{�E���W�JڳYB�I�E���1�_�<�ׯa��\J�v3kTDU���!y�=���=��
��XgX
�{ b�!6���l�ۉ��\wJ�ݶ_LA�d�c0�.ɊͶ�҂��k�4�fMQ������#7a�Uk_�u�ֱy�t�9ą�Y��d���/eT��3����R�y^�@e�@��Ī`n�������ە3T)_@s��N���sz�E�USIbş���F-"���{�t�IߛB�}�j��uŏ).k.��ne���Lţ%͕�"v��拰F3Γ��a�ꍦ�s�0�S��ʩu��.�]DBR� �#09�0����b�[�-B]3J挎�m2�&�Q�ś���un�&�j�"��?gȥ�ĸ1���?�N�ݡ���BiPq�bl��zn6��Oى^�����=ta=�<�c���XWɾ9{�
)��ݎ�T�P:�J���9��l]z�"HX��ѻ�.�I�P��@^u��}z�s�n�?�Ym��QA�'�@H�)��E��U�A}�J!��hf����s=0���h�:K�S�&����a}�d����3����d��9r�3�6wbvD禎p��N�/�����;{���7,#��)�a��e�EFZObp^c\E�lč�i�B%����c�������	��s$�l�[��gp��"�d��ȡT�"�
�\vgLɵ%V�������ѽ�c{��V*.6����aJ!�R��Ҽ;���8����q�u���ɵ�1Ȭ�p!E�{l+�e�v�l����+�8m~�	���U��R�/m��J7?� �w��?�JM�'f\���ߦ��v[\���Qe�19��=��DC�7i����MuG�B-��ՇkJ';S"�mw�����u1�xUs�⺆L���VS���V�˴�.����:i�[��aAg�=1��k����ٻ����D��T����]��K�݈�{����ξvuW��̸�TVU)��N~�������H�G�qQ�����v�Rm`q=+�W����!7��q��]�W��~yGM�9e��[���:ǲ�)��DDw��|�wM����`c���[����ۨiF��R%f����g�b�wjwwG
�8B�c�}w��ث��;(.��H��̷��k�t���+w_Q˫s�8�J�%A�6��
	D�_���w1�ν�����@��ز�G���8~^�o�;E��q�ec��z��uǏsZض#ws��&{��K��86#�c�/�G2���0{w���d��J�7�ϔ�J4�.��o�����9�4r��Z}�v�b�Ol���1�C9�x/:8Lk\�m��Vꌽ=��{�Ujnf�Ա���`ZuuSAy_�d��:B��_Z/�U�" �f�kV���b%�{զ��t4dN���Z\.r\uN"��݋"o5�Xїu���D���/ad-��w{Z�hT�s�!m=g�xN>��K��<��~��>¹���T�>�՚��qL��~O,�C�2�[�MݹܙS�RV�2�d�N�9�H��nZ������3���y�ozZ�
�^x*�����v�����>$�	>�|\����5X�3{9���;JWh�R�i.��$,��1U`��Ơ����EYdm*(�b���**��*��6�`�UUX�c�Q-�

�*�����A�i*��*(�U�"�,��Ue3�U���(��]�;�*m�
I[O-�#��F��o- r���	�!�r����!$�,�#p�R�7�	��Uu�V��C�U����`p�~�������з8��߹N�@�Kh��t�0���`���^C�xٍ��s�;��A���;t�����h[�u�Ѯ%J�-i
hc4���
��l^Tv��j�G[�tM������H"�܇�*j�8�� K�#����r���n4�K���gW*��0���aAP��b-��ދ��<�ӝ��ۑ*�j%�+1�+� �嵲iol�֚S+T�eѥ��j�-�	]��@,M�!t7T�f˳C�rDЊTзj�Q��ݱ=�r��˂g��r�A��k�S.�C�Þ7;K���Fn,9l��@=��]K�.�2ͳ]���xy<I[�,�ԛR���Q�M��]��5ۘ|kvU�GL�O#���M���VIf8vt�r�u��v��X�u�3��X�v֍�Sr��"�OIpֺ	ټW>�mly�'\s��am�A��v[��'4N�������� ыuZ��<���Hz��X��.b��U������G&�{��]�XրǺ�w[qv������l�f\JbU�?�t�K�-<�X��D��N�3tԘ��k��n���݌c�y��Q�9r����WZs��yv�\���v�\�IB%�ю���R��y��;��WQZ��Z�ޜ�.kNGWNu�N����v�6^�i�S���C�,"!N#;��6�����Ck�n]��������bvu��:�ӿGk��f���6�/a��_�m�^�w$L���{��l�ᨕ��IR�����/Yv�x�e����m��ϳ��^^	�~�eV%XV+��
����,�!?Z�m�|�"<�l����%G,��~�W�51k_�m�>RM�+�C{��y��DD�����p�3�-���i��oJ%jsq$C������1��g��.�KL�1=�����C�*�y�{{'��n�5���<lX���:���ْzC3G1�5�h^^�F�r}�w����ܨ�M8�6���MF�	4D@0�m�Aw��9���ׯ��;y��P#+IQJy�9�.�+��}��7)V�s)"���4m�	/���Qxͫ�'xg�\��$\���J��SPs�N�UJ�����{��GMb�{� �bYi�b��p�˿�b�+�$؟�&���n�Z@�wXc����J*�Jg�\���MBezN޾�[��h� ��l6Z17��mUߓ������Hp"�A�ȃ8�3WhV�ȝA벂�	EW�N�pH���߉�A�75�p��r�`СpyD�3�8��n1+�z�wPdn�F�RA;$m\v��b��I�g= ���W�������L�� FOM��d����Pg'A�Ok6۝��������&	�ؘ-��C}V �k�ţ;�b�J~>ٶ �6��X���8�
p�bP�&��&4Ʌ�¹v�z�}��"x�&}5�����V��Xp��ou��B7)V��O>N�J���@�ͯ���f�%&��hJ$9�dv ə�c[���,����L�'a%F�bW_Iȱ�.�	&�3��vz"����(�h�^�����=����a��^6 �����蚳anX�u�#��6Μ~�k�=1U�q�0/�{h�u-
u�d����oe�z�r�skb4p�H�f��&��X6Us��f�)\S5<��譺�V��]��Ak��QY�dѮ�1 ���l�	u܌b���ճcx�rk��cj띵��g���$��W[/fR"\"혺���~O�Ee��[����� wZ�ia���ݦ���K����?� ��P�P�#/X�&Щ+
°�H)4�d��wL�eH(]���5�'	θ�lM�/�\�fk�H,3���
A`s�Ă�R
$:5�}��{�# Ă'>����t���n���&����wo��Y1�����i �Q+��i �45 �}w�y��MrAH,=��
u�7��u�*t�ǷL�%H)=��Hg&����rN�j0�8��
Ad�oۦM2�VR D">Ϙ��'�T}�s�
����F�Ρ��h],��l#�#s]u�Mnv:��a�T4� �-�<�㡁R
AN}� �l@����Rc��
$�Q��]0�
tq�3Ѯ!���q�����:�ۇR2w2C��E_`��U�+�c5�d��ە���s|�d�G� ��|>�?A "�`[�����R��0$��o�}���t��6k���u���9d�s��2T��S�:�4��V�a�<y�o���'�C����+��M� ����i���������$�;ֽ9�G��R�y�1���R�T��p&�++%e�,4�~y�{'	��Ăóz�9��qR
k�p:Ci����i�@י�Ϟy��;J�z�1����-8�I���C�,4�R���������T5����]���ִ֔ۚ����u�����z�YFJ�T��!���aXu�$�&q��yϧ��6	}�1�L��eH)߾�`o���[����k:���B�A�wߝ�031�Z0*X�S�9�4�@��}�bA#��:�Nex_sg�<|���Am�����p!S�}��Cl�����9���$x���ۡ�iT� �LE��;77t�ѿ��M]c�3��g)J���r�N��=���π�
>G�HU���X�|{a�ЁS��kyΫ���r�|�1�gCƤ�(�P�J�q����l+�$� �;�d��󩴂��S�<�m6���u����kya� �|�H/�z�Z��
�q���ed�<��
IX^f$����wѿ��K�Z�
Xٺ���SvW����y��{
u�p=Ci����@�T
%`>w���Xy�����=��
Av���i �����u�+߹� ��<��pJ�[�4��V+
w�CI&���34��Ǿ�͜'s��6�����u�,Z�ިi�AH,޳0+X �����\��w*AeO:��IR���'����#�@DWsj~����� ���3I�`>���<	��0?��#�W/�B�(Y��ीOᰇ<�KO{#�8��'w�������8���ЁS�]��}]l�KǙ���R
AOy������޹&�m�a�l1&�*J!Y(��s&�P*T�p07��}����)E�B붚M���GSfݐv���������N��
t߫:H)���bAH)5Ͼ��^��=�s'L�k�$4$��si�a��m���kp�'(T���6!�J���}󞸜�����$��y�1 �4ԅ-;�{��}��{�p�xQ@�:A�������s��R
AN}� �AH,<3����ֳ|Ä��HV�y� �����}�V�c�9`r�sC��<y��ΒZA`9�bAt��P*u�8�
Af�y冐㣭�zz&�
a|�1��V{ٽ��ӗ\CI7�!���Xs�43H����_c��"V�3
AH)�|����+D:��I0�\{���v��AK�2bk���Y}���+��N����f��S�=��HUǡ�\'4�I��WCWmz�U�y?�����t-=��6}6�Dp۹����^��q�+,c�Q%JRZ����Y�u�BN���a��Ѵ=n0�ۓ]7Z]��r��1P5�cL��8��c�CH�ƙ���nkΏ��﫯�'�d�{��2VVJ�T���!�� ��H):��yهY�t2v�}�$�����c�$�îN8P��Q��@A�<[Hs5��.��`7�Ă�R
w�=���+(�Xy݆!���RT;�R�xLsdx�<R�.+����'|���6�FT����i�@�X�{��߽bAH)5�{��a��*]t�=��� T���c;����|I���S�8�4�	+
°�I�
�X~f2s����p�R
w�X���N+s����C�I
ZB���Ă������R����؁YFJ���4���N���鎔��z��.�%~�r�67l�6�L�Je��gZ�ޟnfw���bAM���OYY++|��4�P*V�y���>q��*AMg�{���|��i���u���\�s/�$i��߾����g�jTx��R�8��H[�ҥ��yF�K`IŊ�� x~�>�`$+�,1&�*J!Y*_>3&�P7�bw�xNSlO9��j�5�H,3��H[HR���$Q�R�
��]�tvy��� ���
A`=�����a�z��[њ�8H)��y�s���9�8d�T��:��i�P*V׹����i�0y���m��:<	� m/#���^��������}�1�d�
$�Ϟ�C��獓�܆�
M!X��2heH(J����|���~�N�����7S_�� �&��'���S�c��|:��#�H{l��
AM T�u��Af��}����Nٸ��a�4���s�Ӯ�kK��1 ��� �Ad���z}��0�XbҠT��sk�H)�`� �`W�u�6���
�tn��vk`p�����
AH)�=`C���VP>��}�&&j�ז�Š�ཛྷ�z��2n�_G�<��`������&�8_iV��''s�uZ>�s7����W���	�nH'�8a��@/�(~�|����hɣO�}���d�]�PWk�]�riO���ڹ{�{��N�*C
�}���GN����T�ei�qKl�뜹{w7[�?=���u�-�@Os�l{�+4g���z���}E�����3��.J�^��r)�_�>x���GE�/N�{O�ٷ���g�{B��4;����;]��L{H��%Č�;�Ηؽ�
f�V�Qt2oVU'��x�b�3�#V��<=y��?sɥ�ec�����Ü�S�w�Ǘy����NM�v�]��1Hǰ���Hg2�`9!�����Z��!0�A����h�
:qƥUZ%Q�He�Z�UE��#mA��m�(��.�1�V&YV0X#�`V+[V"e�ĩ����F ��*�҂5h*�j-lƊ���h��X�*������h������ ̥b,USMU�X֊��Z�A*��EF�
�Uթ���TR�F"%���U�Q�� ��i*���"��0�X�n��|�7�^P� ��!Y(���Y42�Q*|�]�`l��˼�Z��q��^P�㣣��9�- ��c�H)P*s�X�q��VT��!w����;5�1IX�f0�
��{�ٚ���!S�z�؆�
Aa�v���u{�����xޱ �4ԅ��0��Fh��Xi4�S�ۯ�_�ķ�2-#�x�M�kl�ML�1���z���^�X\f3ђ�(��=���m ��rH)/�����}�8d�.��H,�P(�7�M���Ê��u�x�Ă�u�}����`:�c�k�@�N9�@m6 T�ʞya�4���� m���*G>����'¾����kpĜ�S�}�؆�
Aaϖ�R�o{�q ���;�{��+P�&�*^�7[y:5��,��3珛�rp��R
o�0!�� ���I�*J�`>w���\q���Q�Z��U���Ƭ�wQ�Wx�v5ќ�6�^(�j'��>���H�	=��	��`S�:��u����Xg�GIil�s��o�\��7� ��� �AH,�9��I ���l�|0^U�����6�0T3����)s�-4V��-|�}���۵�C���S�z�4ɶVJ�þ�3HJ�R�-��bA`w�Z�o:HtZu�x�H-`V��6M T�������
�FK�9���YY*{�6J�����á�a|�!���B�����M2�VT�{��^S�=�4��|7��[� ����H[H[`<���]0*AN����� r� T�ʞ�a����T(���c)�C�)RPɈ�G�"{���0�x��YXqņ hJ�D��3CR
s�xs��� �
؆�a���7���ٮ ���Ă�R
y�8v�hq�<u�<�a�
��XbMD*J�d�w�bAH(J�y�z|D�q't/���\�n�4bn�ɚ�?lX���w���]������F�����O�.�nmU(W��p��� ��.� ܵ�&[�t�]] ���(\�.��5�[�®-%s�wc����E:4c�ܼ�<q�3F�V{n;)`Mq]2�]rf�4�Z��k��ԩL�5���i�孶��>_��j�5��sC��AHR�|�$��@��~`H,���5&�{�'� Q#��7�R�8�~�>�ji��A$W ����j�ݠ��+J�C���T�����yׂI1(2A��C��\e<D�6�n��� ��P���A����E\�J1
A��V�Ц�'q2A&3�yת��z�0�Rm)f�Xd��cE&TXS�ɝ]��թ��穀#o�	�8��X5�?n����F���%�H�J��9�sڧ=Gcv��(�*2�X��W�gT,��"����6Pz�����'�F�]4�pJ����b<o�d��1N�A����+��C�
PFʙ}K:��ψ"m�	=���w�Y��^�O8�V_����r�%��e���K<)�^�:
��O���R��fWk��_~_��6�|�@>3�� 7)�{�]�n�nS蔒�a���)�TT���{mH7���ZHD\s�]۰b��	�C�eX$���t�M��{we�v��Gc���G�7�&=%���ݮ�ܹ���u�a���9u�.G��@w!.�%��qTv�!�{9Y ���"�I5<��I;��TuK�
�p��@�{�:��\F��&��sd�YkT�7\RR#��l���c�i��|��>�zW��"� ��z�W��{*TQҞ�`u��)7-��M�1Gg_:�zĤ���ΦIWI7t��bH�@Vc}�:p���a�ɢ��B�I3���n�\"����w�^����X.�5WK�n���;�)<��z����E��!����(uU�$�/�͖l�_&A3����.W&�@[U\j��1�t�^��S��l���@VcN�dt4�rI���D�����;�U��0ZC� ��	�~�B�V�K�2�^T�d��#w7
��S7	Q>#{_����%$�XuFuu�g+��TۀA���;㘀�ؤ���u)V�Ԙ*�:���LH=�VtL]�#�u�@U#S�ӈ	�KS���E�ꝩ �)�]U?t}*�8i��)6b�G&�.ͰM+eв���>�9�=Y�"Lu��W:ˁe.���:�3F�-�%r<f��t�rug����֖Ff�ε��K2	���.����Y�u���w�4U<���uQ����q�pK���2���12I7�F�5G�kX���#!�/�%N���}6���M�d���$F�仝������Q�L�+�d�"��r;�0����RwnT�8hF�t.���L�{�ݻF��L�d��	%�����6�r��=<�p�$W ;��\��\R@)jb�֎dlA���UW����|�5-\	#)y�]�
���e�����:�,%��8�=uAf�K��e]ø���lQ˛]�=_c��g��ӻ�[CQ/]W���|I'�� #��@���b�C+CJ��w:$�ݸw�M����"��	�>�,��ѽT҈G�W�>�؂I�p�.�R�5��A=�=�� ����6(q�1�;S�Q#u��7;)����$��e�qa��Ԗn�u�5Z�vPԒ���C�=V���j�꼎Z����Ģ�&�Iz��A��D��mtv��]G��G.�|����3�k�}�)�{s�?�j�߹�X;nn����|�^��;��s��H����T8����#�d�( f4�̭��W�x���?��\Yݗ�0�i-�rc�{'��M�I�{�x��)��t���{#5�lg'��^EE#� 7��B7)��͕R3v H�l�	I*���F���S� �sS$���8�eT�(�O�(7�CZ�H�L��8oO��	�A��G�"9jo2�)7�x'�hA{M |o8_hS»:�M�W�o2��5F�Ք�8��S�N�
��gޡ���f�*��J�TH#����-(�XV�&�� ��b�lR��b��e?}#�(�EI.d���kr������}����7���$V&�n���Gr�N�㟙�LwR��#'��"F�iC��"�"8z���
�H�����<�m\G�Ou�n���>�^g�GbPnP���X�]�#Z~ �5q��9���:��S�G_Q�6��;���R��eT{12�X�}/;zc�� �W/�����%=Үᜐ��B�MF{�,��\�@��ߓ�:}쾄>\�>=����{��3<{%�ײ?<]�Զ_�����q� ��&�H�L��=��	��N�B�Dy;��} ��o�����u�T�mE�G6�:��R���7�*&w���U�	4���!^+���a�Fu=�[�פQ����<u�S�)g�e�aF:r%��\,�Q��{JV�,n�^�g��WNDÖ��u϶�z����Z|�x�2Ֆ�܍sS�I�y���������7��T�Of,��
�E�Ȫ����a!\7ޥ�)�73�������AX���y���
��Pk��eΛ{fe32/ٺ'<��t�4���o���_����~�ԟ�07�}|��|����l��"��R���[3;ź.��qm��/!_"�U�%T()���iJ6�T�QEb�NEb"+�*V�R"*�Tb���T��\ZP-��kV1Ke�e�Z���cb*1L���QTq���`�G-iElcm*[mea��1U���X��j�L��QX�kQ�+\��E�Eێ*+"�.�ES��1�UE��B�R�D��`���cmjcLjM����V,����TUm(�hQ�� �*�ˍ��
���Ł	����Et��U4�3��0��R��������2��`��E��'K��ol#22m(�(Yo)��Me��퇐��2�ɳ���;PY<n�k���B�:9�]�	��bv�e|���m��[fѱ�hƻ�����fA�
ـ���|����BfR0���R��P˵���;�H�������2Yێ���Mvo4��2Z��e�N�x�9��͌��E���&��J�6�?����'|ͺ:�+N���]�9ᝎ�=�kf����7��F{�}����ی�0��i��t15�0Ic3��T��c"�6��ۖa��j7�{aq���x�:�.{E;�u�G/a�u�����iz�2�nMMV��fǦ�s���1�H�K��P�g�ݣY\�*Bņ�DY���j=]�̵���!�ë^7Sô3m�ۋ���qS%<C��s���������-ݛ�R�n����
�Qs��������b�n��1�͵�b�UT�mV��s ۺ��[���yw���^-�ű�*Z+��i-ְΟ�A<��4v�յ�ll��P@)X6Xc����F��zb��q\��%�s��̐��v���Z᭽�#���s^K�S�%Ɠ�ӘV뫷]qه���Nm�܍�Q��u�i�Dbg�٠l)e��e8���CJ��)2|H5����L�F�SL������c����f���R�	9�d�*�q�v�F��6)�؃z�^�pޜU��vV��b��J��6ꩉ�.�$��'� �ifQy���Pށ��>�ڍv�,t�^�h֨=v;��h#2�}���T����R	U�NTQ�n��TG9z�?"9����6 wi��d�1����ꍨ#eQ�E��BI}��UE�5V�0��6����*j��s��I�������2M���Y~����]e՗���q����W^��H;��wi�ﶦX*6d�R�,Yv�2I'�H;�.=8��!�
I+ўL'��ʋ�B��Ϣ�>�ȇ*+FH��r]s�5 �c���w+�ӶT�n8fj�P��6A��O�6=��Uk��� �ݤ�vǰ"�y�B"��2	$�?݈�O[�ZJ��j���"�����p �b�3$�O��I�A�T`��3b��l�g��t ���>Ϫo�Ѐ܉�D��fĂ#S ��k�A�W\-פ;L����G;�[֟|��<��t��d��l�{w�����|�48H(��)J����ƊL���]������>�ɾY��#o�}�R���T�t��Ƞ��J]c�\=bso���_���� ͒���PH��q�0�̻$�"�aor�7/��A����Ť���U6�c�Y�j�r�A�؄fRV�����
b�T���qV����5 �"Ķ�gt��s%��g��M������3��?OM3��L�nS�zwo���ER�R|6*H�φj=nٕ�[����Ϭ.���Ͽ]���$�!S�����r�x�lR�a͙�W��J���#Ʃ�Iu2�;��vԊ�Ŭu)yҴ-�`���9�{[B�0��5�#���9��pF�����`�wTWNߥk[K�J����&�b'r¤��*�$rS$�����\.���k]�@�����^��5��oOvv��6z�)%�D\���.��Pp\CI��i��"�w�n5�=I����aGڥ��rei���Qأ��րsq�m��$�u�Z��Jl�e�]K�u�=�zF����k�[t�d��f���7`�t�l�`ٓ�P[+I4��դ#�#\vo�� 7_�sd�'S ��ps��1�F�f���TL�ݸ&eɎ�L�i��SB��gg{����p����ݜ�`�� �v�7b�dXl��$P!�~ ��p�WOn}gmr<�H{/�z��G:�_����S��Ss�ݽ�EM�$F.}\j���B���~��5�R�9x�H�l��]��yJ�H$��{��"r:���)�]�6�0�q3���O��7u�e?��~�.��*�>�pF�d���L�<�"7bX*&d�k�uH�ő� �X�F�fzUZ����N���ې@s)�r� nq���\Pk{��R��m��v,�Y��D]��ܥ�dZ�#C�I䦂��:�� jX�(��1�Vp??�'��	�LI�B`\q�R�E���eY�>u�}T��d ˦ �WӇ����{&oՖ��ŗ���`�$fu�w97���y
���ڪR����M	YNª'�ɛ������﫛�&~�ŦFΥ�~��2S ��ϳ5�eǖ ��R�A͙��&v�B1h3]�s*ɈoĂN�d���1Vr{�w��ў�ʌ5{^��n�GQ��I��v��^�������y��Z��\B���l�c���6�x���h\3d���ϧ-�$,R���Ů���j�K�>=~�@��z#
K���Ff8��P����'b�$*A�N��o�Z�S���n��'=���󪕃7��s�����g��"�e8��π�Ai��t�\L��� ���_TzA�L�n��K�����/g[����0�Z�;6�N:𢖎Dj�:�= �@�oǅ�7x���/���'h���֚�4��!X��L�D����-픦�- ץ��Ч.�s�Dn6|gD{In�ǈ�l�"�����Fc�"A{� .�03*�s�G���R�x���dO&rems�s�A�lF�`��rZwe��1&�v����۬�Gv]cG'�h�EE�WUzA�n7s�o��I��>�]jir@[B���[���t���M��ny11����#E��ݱ�zn��v��b�n1ә֧����M����5�0�=l��;nv�\q;�u�u��w���.�m΋hv�is����Fk�cYku��Ͽ>�8�1Nc_��|��c(��enϢu��	�XU^3ɂA~�/m� ζ״�Q��7��+��X�$�I�H=��r��N��k��&Ń� �6)V�]2��"i�7�NnzhrSB�;�:l�= �b��3{���A�ܙ��C-Q̮�����*� �����<��j���y�� �q�a�8��v� ������XO�L׀�Z��(b]�H���~hJ�/�\n���vD�ެ�[����0c�y.������t�$W&}����/�M��U"��W�.�G�� L6_kgS���P��FJ��%{�`/e4�8��^oh��m.<G�B��=7 A"�sĒu�A;��z��l�}������&����aK��S���s7Ui�5�W�f�/e��ٱz^&}��=�P3�t'm�SR��gE²	#v�	;��'�0�qar�Hj8"7���$￦k9z{�}�'ڜb��w6��(:�d���kh�ʥ��32o4Fɺ���v5��"�+�� =��s}�d����z�j�KMի����Id�<2nK8,b��UfV*�h�\l���p}�P�u;,��+J����A�j���%�e���;l��;�S团/{��;�b�;tj<��E��o�qW��I؀����6�u��3�@��%&�x��FoaU�4����zb�n�>�{�u3�Yh��GR�3S��/�3oIInR��5:�6
�դ�������7߻��>} g��<\ը}P7��7����,>�}��sOެ�r;�^{����{�ژ�ڬ���_wva�aR��3l��=X^3�%������";��	o���]�A�=0>���y�p��?VM�u��D]ȥ{5?0��|}��}�O*.2�jt�U�QTH1r�m-�P�*;Lt�Ş��yEE3V��<�t2�"��YWe��DA�(�Y�
��D�*�ZT�EU��k�F1iM4Tq�+�&��E-��UE ��լX,M6�ST���1Qv�j��* �[Kr��&҈�-�j�ֈe��"D��m�cT%� �Ro/�� hS	&:'��Y ���-�1)�BMy�>��h_�n={�F�rY�>]�J�I[,G��d�x��7�E�ݎ:��a�R��%�Q��{� e�!�Ê,\�>НS�FJp�Y.�i��m�h��=|��`�Ǧ؏�����=$����L�L+9�Cey���>��D�`�7SA�S��c���7��qlC�E�`!si���l�eX�2�=�K�8)����32	;���KR�
.��U¾�*��+^��܈�Rr�v�Xu��d�#	�>����^�C�R%b����'K�ME5��W�����ܝ���uQD�	��:M����4��Bm��I�������+�(Gכ!�Xv�9k����`)���+r�o�f�=m+��I�A�7v y6��9��`��^6���b{b�F栘�P$�yЄ#��;�;ۃ�ꔘ�pY���k7�bg9L3�UW\U �c践�ػȀۦ�̉O�f6
͞�&�r\wH �Եsuvi6O�b��ʪ�0C>�?LN{�\0���������f��uU�5]J�l�m�k�]���v�<�'�:}���5%�O�)�m]j�&X\�˦�RKc����^��!X퉒�H���52#��5����^Z��ѹ�
v��iL�f�tk�F�ƊL���]��>�_��}�\�$��p	7�>�uy%ۺ�$tFJ鱵�c�.J`!sv@�����6�B�4����鸂E�`���;�+�9�'��6l��Q9\6���r����!{�0;���7x�9�M���\��,:���ǹ=x��;P�:�{�R�����s4����P��5Jꋆ����϶��BAM�@Y֘}�L���n�Ò��l��)Bª5�0b.+{�V��M� a�s����쏐�}���SKb��Po���>�|w��� �ܟ��\�����}��M�2WJ`-�hA�6�ϟn� �i��EnA�Ų�wX�ZEr�z��ٹôw<>m�e������G���^n2�$������%��%�U���n�G)���	-Ԏ���(����v}��	�	��H�؂��k�[���r�=�*����k�;r���[�`��q��
0��L|L��hSF��t#�YT"��w^�u�z�덉�bsD��<w	���uj&���2tF.tg���1����ۼ>�@v�7�Z0�);f�ԟY�A����w]����n�$�+ރs���w[��Ӗ��L ��)�{9ۢ��x�EM�$#�8褤�DJi�E>�M�^�z��r����w"<w��X;�2�b`�o�#�P�]���֟�WprZw'�ڳ��usE�UU�$��P{h��z���d@�1���U��w�ҍ��$(�dG�S~$8s/"wB�M^9̤V/��2����C�m�{o���`"�Yk�M�c��饢��cQ.����24υ��{�R۳�n��&Z3[Q&��* . ��H�A6�idI �7D"�N>�k�7.+�|�6!X4��}\��O���d4�p��L�,h�)\k�A��p�#grQ��=(Jkr:��A�E�yu��n�<��id��d+�b�;�w�r*�Zߎ�!�ks�蔺����]���р�}�g�P��LlP���%D�=�,�Bm����Y�5�V��,�ԎT�VtAl8��Dl�˗�b����U.q5XE�A����*��t'8�Y�v1�g�s�u�v�ӯ�tڤx�8�;�$�;��gV�FP�]h�q笙E��516�.��V�"�ѣr���V���d���4���O$�k�sV����#%x~o*�Y�B��6�ٻ\4a�Q^}M�[-�;or04L݊ ��V��z�\u\�Q9P�	�pF�\qfL߳VȻ�{(Jj�sGo��G!�Gg1l��|��]g(��!�s�p����W��ZC ����3k�һƼKșI����T{c�G:-U[]��>R��c��e��:�ǈ;����4L��w=��FJ���oĻ�Ҷ����#Ϻ��R#�w���7�w��vH�1�/WG3L��	"wcۈQ�^CX
特�H�uυ����.��h ���ā�#����+[��}�����l��M�R{ k݃](g�uGn�<X�?N��y�@;���D;��W�z���.=..]L�h��71��-:j�ԩ;�F��
s���gM��ޖ|T�m����i�±M׳ӯ�+	:p��w�/N�c��*���0��O�I��|Ύ��X1i�亥��""���Z���95X�Y��i/#ڳ'<��`t�>��[]M�[.��m��u�^gu�c5f_�)E0��J�2��Nl��FsdZ4}��L��{��^;� �uEQER2냭�o%���~��>����n��,`!_�C�on��;�PkF櫈}D��h���7L�u�!���1�gL��K�g�*�Z��g@ob����;�A+���<��22W���D+4��s_ٵ�9��������]��!T*��"�ԝ܇���6W8�aZ�֦��&v(q���֓���`�3��9�^\�_����@����c{c��-��˔��!�2��7ɞwu���YD�2��ݺ3�K[}L;ܧ��� m��4��R��a���G;D����}M�(��o�-޶����wB*�]R��⩑S�{{>;m��)���YϹ���+S+���G.sm�.�]�__�v�f$i(�N�H����&�F���Zw
k��)�/��R;-�fN�������F�o�/O�s|8�E{g�O'��e燃6R"	�dEE�o��c�˶�ǒ�ˣ�Q$y����ׂ	T�k�6��n��ܻ�ʥ��pS��&ݟ���o: |{�ܧ���3�A�{�9Kf�^�[ܫ�UN�sZ6�%�Gf_X/oh�c7ӏ{]�\Q�\x������K͛[x�'&��X�^�^�;�y���f���Yn9[�gjO�Rw�mr�sN!�p��2<���{�=H��A���.����r3�P5!ټ���k3Uͷ�7ƵfN���{٨a�Z>�+���aH���`~�y���N1���'���^7��w��N�vV�=Ƕ��m+�W��f�e�����0����޳�ڑ�;Zw�;. ���V E�I�+�
�x�9��#���_�8 �d�$YBʬ��eS��j�kq��j�ܬ��YIǖc @�@!��L��U��oWP�"���Ki���p�A���oX�a�kF��yc��lSmE��*�R��,A!F����� �"R���J'[��JYIR�h����j�j#5s-e��f�pAYl�J"��V1'$�o�P�Bм�ZF��R[;��%8�������up�.�,B�{=]Y�:�/�v��xY:�l��t�2��L>��[�k��p�SW@��hu������\ʢ�h�·M�[���,�۝�uY(X7��3��]	Pٮ�����0�OFy'��t�^�76�[]�*h�i\.+U�G� �2�c����T۬��kGZ�6��Q랷m�f�M,v.c
���Թts�1�+n�X�>�L\�>�s�孏b�6X����1�`l�(D�,m7a��]oeh��K��uv���<O]����ë��X��n�Z�y��,��.�[� ��H؎e����v�+����;e,���)q�YQ[�ׂ���vL�t"��]�D3��mH�\��xM�Xn�e;��\�ƣ�Wn�]���*����Q�X��b}�cF��g�Y�X74�X&�V�M�*	��	b��0�46�����wdo�ͺ�]�xジ&\��4������t]����b8�sIj{5�UU[QU���v��O����${��v���іY�{[��Y�����0�w;���2�g�ӳ�/c�ň-��p#�� �#�P\�ƹ89N.�E�nr��@.�l�ف��h�����<��nͺ�Y�vV'Ô�V�u�6���Vuca���n�r{=�`������29��Vדs���� ��m����"��[�k��VTU*|U�;� ���6p��*f�E���0�.��}����s��D��h6�O5��QÛ�\�������������g���Q0
��*�*!�v��c�G%]	R��r��2	"�ʨ_{��9���ؓ�1�Tn�>�Jm�U:�/˫<��K���4�V�
ޝjpt�͞,���׏M�������d�.�F�{�o<�W��	̃.������[ghm��TC"� @&,VS�O���Z��H�d2L��{�9t(����I4��A �s��FSF�O)�����߅����/o��D4�F��pQÝ֡��ߞc��`��MG3�v���{p�����8^��f&}��X�ݝ�����EyyNi���}pG|�f�u�jT /vC�V�22WF���w��@	���I�L��nn2�t��G� `X�7g��|� ��"�#�B���a���{�( |���։���'ܹ�1]���[��F6��PW9Zk��x*�(��m���=�kQ~�+�p�.���x����.V� <� �\_�d][�����]2��tn+ 
]��e+�,��oY����{� ̯�i���{�g�uOG��l��dB�Ur�F嶪Lj� ;��ma���z��n+O)y՘��F����L�b�#<<�S�,�Qٹ�3�YR�>���`�k0S��������j���6f��	��⊷YMev�2�M61��b��T�,�g9��ڨ����1ɑfK$���M�q�����Sp�m��do\��^yE���=���oS/�0ZX���G���nm�y��� �9�p"�����jn�Ο�eh�#s$A��n���DWWT�8u ���Y�V��]F����+S+�z_�8�KK���A��w!ζ��t�`\�7G��|w�ʱ�`-݊ ;���=��ܫG\��9"ߣ0�G��
��(�47v������)y����0�.��'��l����K��R�9A+Riv�y�ъ��k����q�s�@2\&��[km�tg&��3�ƃ�YV�ff�JB[�)��9��.�Nm���h,��W1�[t�����h��S���v��z�.��Uz�QT�i��rDu�����u��f>�*��T�۬7pl�pS5�n��߱rr�0^�T���÷�!�ie�ۢm���{�O�u�����]��:>��o��{�m�@Xu<�fN�vd��Q��m���	��9*�^Ϲu`��4�m{"�:��y<<3c<�Ksl5h��1�c�|���.�A��Ӆ��ԫ�ǯ#�w1�%��
�id@���GD� 漱�l�<s���=�ˬ��D��W_V�C������H�F�-��w�*������ ��twla�L��w�!!�0̃��CʮX���etLW�R�{}��1�L�`��T|���U��=H0Ok�b����;���Q��4I>�̦-pJ�Y]��}�g��d�_�S ���X��:#������j����,���ʅR�mh�#sZ�<�s5`�$�Z��H��	��G�۷���Bɶ�l�X,q�)^l�R7�.�en�Y;7�!�]#��8��'N	$�k����lD��-w껻�f3�o��f�T���LNkT���1g7�wi���]��c���|n5,�T���:�F���T|㉺m�鹾Ej� �)C�������������b!kin���O��� f6´ݯ��X��'R��b����y]�gs.��9.X�(Q�F��Ȱj��3[$��:���MC�&`�*���5��0�D��4�c�<����2�;��n�7x����7��#n�8��WK=ǂͯ�cL�36�z�S����5�LZbC Ym�b��s���,�����w���4;�1M^b"=�5e3p�k�K���X�r���f4����_h��9�P�TdAr�D��#�ә9;��f�A�a�q�톢�����t�wY����sV���uZ�"k������^�a�I;\һJ��	z�$�N0�Ƽ*�|eLn�ɣ{�a�H8%C�E�g�.������~d�4��RK4�mm����4:T(Y����pfs:�7&w����9sV�3��@·4�j�`B������sp�D���7���xSS��ǵ�s��X��)+��2�1GMGV�4ud^u�΍u����E	TT�rI����W��ۯ��^@�Wl�[T#�By�{`��������en���j[$�.߆�ЀK��Y�Ԡ�CC�Oê߱n	��H=�?A���i��� ���g���7 �u\�����`�	��*ބ����w�L�H`�wm�7��:���:;�4���."!6���!��<���(��ߒ�'�}H�^u�&�,� ��"�����;m��s��k"S�%�lv������y�u�Ɲ̙�w+.�#��$������h�d.�8	,!!�0̙�~�TI��\s�<p�����n6wIH�]O�p~�a�ȏ�� �ZF�*<� �R1�P��o�x��P.E�+n6� `�{�������t���#P��P��mK�_�������{�@�I�`��{=����֠]�`�@Zq@P�Ҹ��/�G\A;m��Hfjw:)0�Cι
Z\�P�B�<h�����r�_t�v��K˻q"���fZ�ߴOMB����F�t��;�DA��ࣔN�1�yמ��|s��;�,�v��>��
Pj$:qa׉������Z�J�/��<��X�sy}�8�H�S�A�vEW��5L�r2Yf/�#W�j���LV����K��T��\���mu򷒍Z'h�|�{'oZF޷�ʧ�׮�T������\<�2��d�೉9��}�C5�CW�7�g���9�����ә�����΄�nY���'61�=ˊ�ކOE��\E����[�{6V%o�[��-{�֨�9��.t-���m�RU�[yj�0L����p��`Vm^Q��?{�D�4���'���K�
Uh���D �d�!��m��VM�;%5SyU�F]
}��^BJ��V[\h9aQq��1XT6�E2����7t��ۥh* ��0�^nil�PDPDm�L����K\B�&5���Ȱ�,�1S-1�T-�ib&!r�̦ �Ȓ�;���D���#l-A� p���^�ZC�Jt�t��;����xH�@;�(D�l��p;�N������mjcr��eq��QE�5��D� Ł ��� f��%���um)���F
fW,S�����"H7��a	�[ܑ �Ę�k%��þ8�q��W���T��Q��WJt>�B�>�rx%�+S�@�V� m[����{|.��$b�'�T�㰟jjn��u�	���wl�j]�r�WZ=�P��o�t�[�A�㖅̀z�0��UR��k2�����u�ϙ���������J�2��|I���ޯ.�E��+F 7u�b�ꭘ�;u�њ �2Y���A=������o��Vo��`ż>��H3ٗUk���������','XBS�F)�>�;��Vs���p`.^5>�֮ns�ث-��*'�I$R�GLC$��F�����H�Z�4�8�v�#Ǳ���<x�"�_R1�R�?6|r���v��@F�\@nS�T6ga.L��QCb�	'q�l����k��wd@w[0���ʕ�V���PwpFdǠ�I�~ӄ��w#�8�������d�x�g�i`ɍѰ6&�A m��I���޲�v�mt٘�O�vqfj�vl\d;��J5�zJ�P5륧�Q�f�O�����*Җj#V�s����:�6����	�wd�Jq44�3m�\�0��WYe�K)`M.f�eK� ;WNj]uv�׶X�8�]�!(qf+g�n+`�=�&yݬ��\X3l�����E�..hwq���܎t�99��bz������Lv�eaȭ�\Ş�7@��0�'Tvk��~~���Pwf17[��[��![J�4n�U	�-�lZh��WO]T��a���4Ѓk}}�ق`z�*�8E^;R����=�ڭ�w+�#ag �w�e���c��5�cf��շ]�%�Z������N�m0�� ����8�}N6���K���9�Ew�g{,7[���┨Ⱦ�;�)m�ÓS-7wiRQ'O�ۤ`����9J���E֌���Vg&�5�|JEj���Q~>긂I�&:XC�X�ǋ>��t��8�J��kڎwj�- ��O��Rt$VH@�L�Dفi�J*����I�l(��b�t�F�?^�uS�Ҳ���j�V��1�t�۬���I8����2�p����f� �w���sM /vAo�����Z���ˌ�|x�g���3]�y���288fL�@�	;��������T][�[0��ԡ\,���DC��M���K6�ژ�8�njp�$��� ��þ2�T,:�$�S���կ�ʈ<��h�U�������qB�$���w�c!�A��j�����Ke�IP�g��l�f����c6�|�|���(�Q_����ulC��l1�50��2�O�i��+�*:4Ќ��z�����hФ�<��b��n�4����������̦��<�UG���yp�Wh��.�-��l��m^��7q]nx�a��]H
Lb(R�jL�y�v�ϸ.bGAX��յb`m��6��T�B� wrNP��پ������
">pL%0��\�K+�������u�>�&�+�����&Ƙmh�t����J���M�\��H���F�R��R��X13\r}�n�~����ئ{���]T����⳸4h>	��f��D
'�z�(H��3���N.;_U���d�v�Gs������ww-^áI	�:�w5��Di�-$.1/[�*cW�;0�0\_�^6���ƷV�c���H����ħ7�f&ѐ�:���]Mݕ��Hhb9F-��e�SF���t�j�nB5*�ݬ�nv���ص���z���W:i��)�fJ]��~`{�]���u04�gK���o��߄+>�������!wi{!�>�\u��m���a$��u):��B�� ��C2����(gp�S����y������b��#y�\� ۓ��e5^22�CBտ�v`��$5iw\����r�)R�ަ<X���_7����f�`����|�5S�܊HU0l�&8�%��,h������dF_G�`�|��	f9���u�vNQ1a��w�;.�1]E�Fй��
I�Zl۝��,�y�I��}�~�z�DԌ"�_x�D�d�������o��P�w�GR��9�L�e��5�2��/���O�(��I(}r%ף��A�~�ŋR;�?jaqv҅���{���9��A%DX@���@�칾�>����#�.t���4�a���$��OwUb�ʝSi{�@�wX�]w��PA���J�hDA�=�~��Q�_#j�� /u�Rwu�}t� �,:���WB	%V6�9�z���e��"n����q���9��]���X|`MNl���a7;5�* l��~�RR�c�����ԥ�;r�4b����vm�|4*�0�=�O��]��ȃ��P/�w�ˈ~#gX�{P�����/��%���V�y�ӶʎFTy��N'p.k[P�Ұ��9��س����݀���w��5<^�<9N����3u��_^��ަ��EDb�v��=�����+�:P|wޑ /��;$�7��p����ISq�kS$��'j�����ۅhك��m���nlw��$�ڧS�t��>�$ɘ1�y�s�߶O(Z�0�ԥ������ݎE�\'9�.,P��Z��i�9�F��Î4��ӥk]8G=�QY��ݓ��0A��B�V����7[A��y�X�
ʿ-��Ղ{�����۵w�;� ��R6QB:��!��I�e�z&�H�Lqi~'kUWZ�6�mz���Б���u�u�ضgo�3X��5D�Xd� ��اj�{���F}K���������?��>�V���� i�t$ ���Rw	 �Շ���C�4Ì���5�O��h��M�k�<��Ĭ�l͈k7ɽ(;���$	$,d���^(RO�����O���3\J��Cd�,����J�� �	���v�ϭ���}�!����?�DL��a��C'�H�4XtjC����NiC�&|u
Rp����̖�!��s�f�� ��Ry����<��� 	'0�� �BH@ ����XY0�������|>�����x	��?����_�'��~p�C��4��턁 ���������C��� g�?JhHs0%8�w�!�=��1����[��H�O�~>�y9~?i��?ON%1~�'�찐  'GѲ�#&�ˆ�ݮO�D��.B@�`� �V@�Y��ȧL�����?�\�!��='�넁 �'*�O��?PM�g�k�'�~'����c��M�ɰ������~���p�����?Q�?/�~&<��q���}�e � ��!�>��#���P�w����ph)�4���0�����/�����C��ܟ07	�P���t��gē�~!�~��C��>�  } }�#���~b ����>7'GP�:?�
��>ޤ(�Bk�$�� �2� ��O���v�h-!�C]��J$��tl�|��? �,�H@ �8��A`�Od��i"��O�^H@ �d�@�9�Q��l��.�4�A�Z�����̄󀌆I8�Y��$����@��L��^��pI ���a����H}r`H ���0d������?��?��||ς̞�����!���!�I�j��g�D0~g�$�އ�<�~�~�	��>�?��_���� �?	���|ߜ/퐴������!�� '�6~�=L?�?��a�C�P�?�}���C���|��:s 3 ���.�#�����ϐ����`����C���$<~'��b�~?��!�;<����D>\� >ߴ'��k�'?_��?t'��(�@w����a�0�����_��d5 P��nH~�I��� ?��~S'�C �~��	�?������c���! ��?D�82pM�pO���8��!I:�� ~�͜�Ab �q������	��s?�rE8P����\