BZh91AY&SY\���߀`q���#� ����b<��    >{ᵨ��5�Ҫ�SU��m�5����2PJ"����(*&��Rڙ��4�
�lԦ���١RSX�ԉE�h�o��)�٥TM�h�MP[1����Ll�%*��Tl֫-��-�%(f��l�ɶ�͵J�k`ke2��UY��6�2Dx��f��µVգM���UVf��,�f�,�*P����l ���j6��m�l&�@�b�m-m��Z�Jً+m�XԙY�+Z�w�!m���́� ����ҟvr�G�Ov�ךU��� �ٶ�V������0t��u&�R�q'f��{Ӂ+n�2�`ƯvE֬��N����m֦�I���E��hjx  ��f�(+���q馕t�iq���
��U�g)��G��yim��*�C���֝�;sx�ԻeI�Su�R��ڛz����^��7Bݥb�+[mU+*���i�@�5[p  ;����d���R�����z^���u*\�}��ol.�;�U���;y�J��[q��|J}�����ϺU��M�|��J��V�z����֗m}�٩�ښ-j	���  D}�S���v���O�T������.��)�<��_m�s����>}򮚄�k|wϾ���{{T�L������}��j��{�	R�F�Wt�jP�n+p�W�����)H|�H(E���1v�  �����*:��Lz=�U٪�w��{m=�)�ewx�.�Rh�[yz�尳)V��ox%Am��,*�{i)�W�v���;-M�/w���n�^]�Ueӻu��
��֦��m�2�3#� ��J[�O^z^��)k�����������]������ޝTB��^���6��S�z3�T�o=��ٻ��T�ǝ��Y�zr��i.���_3Z��d�Kf��4�4ٯ� ���%)k+�Is�J�hu�W���.�k*��Wt�ҕ4�q��R���{h�U�]�:Skf�;�������oou�N�{��{�U���C UuT·��IA�B�D��jm�����*�T���P�z�1޺=����Pѯ#����h/+�UQ*������sɺց����� ���D������2*kcS6�f�$�Zo� ��x����=�@��Wy��zPνs���c���֥�����z�PY�l�����hz����]�އk�(��U�UE@�$�=m�� ׾����<��;���Q{���E֔ކ֝Ux��颯t���^�w���^��n<��T���+p�֗�       ��R� &LL� �&L�"��b���2i� �� 4�M4ɉ��JT� ��  a���J�(� C&`LhOIJzmSC@ �h � =R i�� �SOP4��<��_o��}�y�8w����V
�Ţb�����߿-�^:���{�﷟1 Wy���A@{� ��
 
�s���@ ~��#�����G�ҧ�� 
������ 
��T��EA�����������V�?&���voɑ?K"{`O���`N0��D�(q�8��1��q�8��d2'�
q�8Ȝe��"q�8aN22q�=0�e�
q�8�e0��P�"q�8�e2�C�	��q�8��d2'���&�"q�8aN2'�)�D� {a�
fD�
q�8ʜ`^0��8ʜ`2�fT�*q�xȜa�q�xʼ`2�	�C� @2�<`x��fT��@2"�dU8�
q������"��g
�� G��0��dTxȠ�dPx� d̈<`PxȪq�T�)�T��N2��N2��`U8�2 <a xȪq�T� �AS�(_L(�T0�<n�Q2(<`xȠ�A�
��@W��/�@� 3�����^0�`2��C�#�̩�D�
q�8��aN0���8dN��	�D�q�8`�aN0�S��݅8ȜdN2'�wa0'S���@�����O~{���<`��{�Ǜ�>0�ݽ�����2���ld��۔�,,���2���g&V���̈PtQz�N�a�oB�N�If�^����RJ�+p��%ԏ6��[��#P$�p�2��b{tm�`�W��"��n�J¤le���$ݸ���y,�'��Vh8cn\���)C�����L� Ʌm�S��5ZD�f[�l���ie�X�c^Ēݡ�A�q�vƙ���YcH�F�Z{iC��aK2�cnL��傅6���4M�vɴC�1K��B�U)�ٗb#��[qjr�)
Ûv�� �#����\�ZkU똝Qä��:�̲6�k���6$�`�T�/��ÇP�B�U�48n��WKI�B�H��0�T(vp<��u���ǚ�۷����g�5*�m��3c`Œ�YYO�p'�)ٲ���Z�5�w칔�nT�P�6�C �C�s%%��N[G^S�dz��E�@���'W�aEX��f�r;�Ps����5��k � �X���avh�5h�]\��hϙ�ř$
G��Ͱ&�m�Y�&j����YlJu%6�G�
�//�ݚ;��ޅP���v\:�	�at�Z�U�v�{z���HkE���d�%�����q���/?{��#�7-"yf]u��֛����m3* M�9yy��kvh^cF�Ƅ��Fm�YY���b9��������AA�܃e�������JISY��b�a�	s<�[5���>H,X���W���ךYڛ���2��ػ�)[̗q�"�6
{�Ń(�H�QnfX���D�J����h2��P�)*��oD��ƨ��cdf�KƎj���5����6f��lǑ��vrA��#F�aY1AIdT�[:���F!�ݲ���3�iCG����y����Z#ĥ�lz2�jg�{�"���$�xт-;����Qle]bB��2�U�*�Gi]n�'D�NV族$1Ԍeָ�̬-�����1|l�snԔ���K9�E�т=�ڍb��0S@�+,��n�Շ�PL����������},.uK�����A��R*�1<*�gi
�Ly�-[Ӻ��㮈�֐�M�G7�\�F�<t���^��l�ߙ��ƍJ���?nͼ�V�v�hʏunj`H�m�d�rQ"�Rۆ��fn�7S.2�6�)��٫q2���(���-��c4��4m�ʰ7R#b;�l�#�ov�,Dc%Ey��2QP��J�M�`O-��8A+;c5���b����R��L�*(�ٗ0P��2�ˏ>��c���x�@�X�{̠��;э�Kw�qf�m��2�D],�K,�J�/v-���Q��B�cEz`���E`�TK\��-��n:v�ڤ���1:ợz*P��3d�;
�7"7!�m�
�bSY)T�e��1%�(mfհ%�ɛj�R�b�AϚ��[�1l��u�'Gx[<�J�	4�mf��;�wQ�K(P�Rҋ#UD,�k�R���Z�D�${�^�hfֽ����a1Ǐt��L�Ո�6ab�Z��B(Ƀ��h�'ΦX̖�2�g�k*���[ó(2���H��nZ&�Uxtmk�&;�[� ��Vc[A��K�f[�!ON43ha�R�ll+�*�FU�p�6��0���]ʞ�:�Ű�}݇*��S���I����-�3(3���e�������6�
�,L�.M��I����5�)�L�mٴwR�ٕ�u)���A��f9�J�u��4�SC��"AT�Qd����ܻ�4���&c�f�BwJ�#��Պ�[w��{��0��cL�a�'ܼSqa�Э\��:н�K�+C4i ���NT6�L��:P!�st\����H!�Yָ��FV��[��mO*f�8�}rá���n�qA��ػɢ�M�r�8���Rz��&l�g�!�%:�.��������02�4G~�#�v���%��*R���N���`a��j�U�N�f�������tɚR�3��;v����4��z��ˬP�7$Y��ne��Q>2�b�#+$�Y��z�@�J:��� w$un�;�G�ڹ�Qh녚��p�G�lBo2��� 6��U�f�zvƧ/,K���әf�.b��Y�F�V5�=١qi̈́v�\#zI�i�w)
G.U*�e��՗[�ZFm��Ǡn��/�vٴl�U���M�Z���^���L���* �
����m���0觅 Q;2��t�SB��Y*�R�����y6���{Q`ǣ>l���[.�^�5yˎ�e�6�]�anR�5�(��q�ܢ�:���YeȖ�\8 hVM-�9Pݰ~%n��l;6�GSt�7���x��u��<��f˱o ��hn3�C;�	�4��Y�s[m+o"�fa�U�r�H�K��4un@�3�4mDVVU�r�ʺf�a�W�p�):�q�j�LH���&�D2�Ɖ�j���\1�qF"��f2�b�|��8hےmI&�nV�%�%iP�9Dk���o
ˁV��ַI��3X�6�j��hPQi{z�@ј��y�VY��Q��6����^fnV�S��6���(Ћ$Wr�2ʏ �!��0�Z����u�LҴ^Ѳ�=�h��V�v�������f���e+ض��D\�����6+ur�Cf�L��LY���1�Ȋ�����7��*(k���d��~����M��2�-��q�`ֶj©��7s1Z0�Y�� ��z��4�����I�n�F��$�h
f��f�����bF�(�Q,T5pYݱL#%�ʱ¨��Ǉ�p��W[[.��r�Zsai���yVv���o吶+[l&�K��S~;���ĩ���Ri���c[R�O�g`�����vͺ�O����|(Џf��RYu�bTf���j�5U3nT�E��E�Y��h3L�#�be���خ*��|yֲή*�.�d��*լ������rԅ�FR:|��k��0PGnՅ�x��r�]vf���G6*� �Kk5Zp*��-ߚm��)��;�r�Y��_]�sZ�L�����5��J~7a(5'�Nm\���z��`׏@�igF3� Y�`�qi
$��G2;�4m\E^�z&�8$�6 �jeMj�5�4ޝ�Ԕ�o����I�
��w�ʼ%k�cd;n�<��f����XtEDc�%���k�U(:7��ff��Y@���Qsb�&d¶R���r��0ḥ �/5��,4O�3d�zMT�[�Q�K҆��#1n�Tm�v4�%P`�7G%f@K�f#�g714uD�̤�kŐ��ysZFk[��e�;X�$���u��5M�QV�����*=oS�7��b�A��qԶ�	W�
4Um�YdV�Ck*�������,*�UScFC3\f�n]�Mhb�b�YZA��(U0 �83v����s,[�CE���Dl+tr��7.��͛����3	�.�T��1�ఞJ��):�H�7P#NcǠ�S���+7Cs&��ѐV�PVЛV�Mn����[&�d�wlCz�5�C$d�ݒ׍<q����na�QglV�dC'���i�Q3�U�j:�3A�)�Ũ�,�XYtq@E�&mnG(��K����V+�M;��G	�k� %l�x^1�&�`Ǹ�@-\�kw�����y���l��ie�|�@Q�j�ѽ�d!mлj%%�l�M�idp]��1᧖���A��gj�JR�H��4V�a�XT���c��L;�LL�R��-;հfl�����B2]�Z����J�uywks2�b�ɴ	ѐ��Uu�3]��:T��ֽ{na;S/fhke���)�,�?��C�tp�M�Ӧ�S���~��˻hmK�̸ݸ�i왦BI�/S�i���J�eP��TO�ͳ�d
�L	��݁��m賮��e<�"��D�ͼf'�^�����St��³��j��`3h�����{�`s�W�']�o ���*�l�
�hV�%�X	��IqKL�m�E* u��ѝ�n��Z���y���Bwb}wlD�ub��n�Q=t}Q��[u��f�'Sf�A�n���܆SV�d,ǡ´鵇S�Y@Ь*ؔ71��Z�T�W)��2�[(U�x��T�
R�Y��h<A��.�����IP��&D�R齢��BJ�A,��q�&��h6���U�s1��̆��wqCE���W����u�b͎���Rʎn�P[��,;���V����lb �[��(˹�ܤ�F�E7-�*���R�kp����'�qB�+�D�0P`���[�E�-dL�t��FT�t��E�F�h��)�[��6���YPlFa�b���,��h��L�Иk2-����k.-*B�[kB-�w��٦	��F�-��m��{�a�rn���а'�M�*f�%ipm�sM�k`B�Ըs0���~؃�4,���b&�N�©бZ�ɹ���`�6���g�'�{*���F^�e�}���c�þ�z�"�.�k{P�(!����`�۴oNJ��s�AṮR��YH(�"�.ed62����5�]B�3l�E-qj�An*�X֓�Ec�#�j��m��+/�\Hh9�����L������4M�I��%n��Kg�X��{��1yx�����ܽ�+�+X�X�l�«wszֱki�J�/m�VE��27���+�uu��r�0�0���elp��1�$ll��A�MÁ����A���[6$wJ�`�w��{�r��q��y�����@��^fi��쓤\����6f���"[K�x�j���5g#��fRl�((.�S��'u��t.j��y�Z�:NM���-�ύ�Z�5�C��m�X�4� �Ҷ�1F$�u�o�eh�s.�X� y>:�e�ʹx=jj�JY:m"]OF��e��j1{N��p��ފu���3u��ג`���Ξn�+4�If�ꉧQV��5�K0�2�p�������Y��u��mřl{L��l�/Zhg^p͏X�Wf`:�S��+b���m7En�;��g��JJhR��^�n��r+ 9r཰�6
�6˻u�~�h`&���!��X�֧Y���[F�x�>��2�3>�"�E�����X�v�RJ�[_E��@*z��@SI�b)��Y���MU(��qR��e^4P�d�d)X�]`��S6T��
���g֎L��Z�����t""�}�o��K~e��DA�$�e+�35%�V��df�݅3Y���4���z�BŬ��N\��6�{���<���۰����D����uoB�3���5�V���B�/��H���J��B�(4ݴI��W"!X��^<g���Q��&
a�n�k*,G!��F̱�X���&�����F����xŕc/!3l�����czc:���[̕.�fM�sS�;s//a��D9�ɣj�Xs�!Xzܭa�2]Z���{�%a��nԪ1PQA�"���S��6en4f<�F=�c;H��N�3���-
�i%b&E�B�Śݨ�!��7��5��Ɣu��:�%��G�ru���]�Ξ[�Ż�2�T6/j%0����Q��H-�[[���~�s5�a��{��X�`�[}�1f�h.��>��@�2[�+�v��";h<b2�H��L��y[�*9��n����2�i���i�֌�Fɭ�9��g[�{xSo���ch�z�"��'�֧hk!�3WJڼ��¾��ۛ���2�sb2"�P�/11cE�r��M<�϶��F�i�7k[��+� !b]�c1X�GRwxF��P0�!MbUI��Gv��]��0B.�V-֒?�#[e��]�x���l����`���C�����n��&̖PչvjSJP[@�s\�t,�eܡWX�b��ȽH-��×�laӵraQ�i��5Z��SsijƄE�n~�X���eʳ��e8/�[��䙪�`'>�Nnm 5sQ�Z�SQˌ��NZ���1�Zwt�mi��NAB����K,H��/E�l�i�W+M����<�˕��e��h���jӳ�ݚ�{o��Y��X�Q�sF�UP�ӼfD��`YI�5w)6��Q̦�.�
��Y����46�P�����˄�P�T��~�<H(?�q!Gm�t�;ic%��fȚ�n�+X�MS��b�Ӎ�d����u\�A��M"nUm����K���M
X�;
Ww��`��3F���R'�Zvw4Z,D�I�(J^є�$!�Ӛ�A!Z��І���E��6�,���:�c+��Z�b�%f6h�R�A�Z���]ə�i�Ō��7.��v<��'I:4�b��K�2��ܢ�T�t�3�U]H/wf�c�@(ؚ!^T܆�2�	dZ�WH��ܻq���LD�K�7�B�85cf`�XʵQЭ��b5�cUrM	�4醤�c/�R��5͔p`C1�Ҷk�oS4)3�wY��p���u���j�qVau��S5$�c�,����F��s�k��Zs�a�KT7
�W��d����ak�QM�,%�����Ʀ��2J"���R�ܬ��oi���g7q�&�[W�l��,�˖o!�PR���4�;J-۔�\0�li���T���ު�;`Y�o
��;�����Յ]��V������3m-�;���H���b1�;�9>Z�e�gh&Z8���Kč�K�Y�M�C�ufPD�;����.�HbI\;����&��e�ad�^1�6M	!�/�sɡ���~��	�{NÆ7A�jP�+�P��Nժ�Ʉ���o7Wg�-=;{E���X�JB8�u��|�����pzCU[$� �&�o��8uC�,�_Ҩr)���ܽ�
���N�x�P)��si��ǫ"jyh0vfb'$ل�oT���Rn�L�3X���-�xO����v�MY�*���~{��j��� �ޟ�{�	���>�����ju�h�`�F&�XW��ʁ3Y��H(�]�Q�}���wx�h�!��"���ZE.�FV&47��٧�C&WLY&3e��%lڂ��c&DcQw*u{Xok�W|[�i�~x�r�uj�m⵽��\:���]ì��F���r��x��L���,��h���&6����.BP�u����������n6�\�Bk�[R�#h��q��!����EQ��o;�v0����/�Ѽ�Rn�`΢��Y��Z��GM��'�A�k���jJ3X��Q�F�+>�QKk�Vf��J�4��]I�9���3j�\�8s9�d�4�N
\t�Sɼ��5���f]�&M�#J�-؆�1�u+Mn�M�����w+��awaȪ�pW(M�ɼ?G��Q�9��o���\�[Ǹ	��I��&�v�A���n�c⧷}m�l��|o��-�p������!�j^�Ar�m��Y�L�7��:�	�[.��R4Vm��"�F�=�;���Jb.-b��Y���c �{¸0�;��Ww]OqP0^Cl�S��%���%���k.������ؖ��@YM�K��Y�peoi����Wŭ�<̳����Y
V�#�,�K{p ai9�U�������=���l�*K4z��zɣր�q�9��g��S}�	XH�0Ղ5Cu���c��F��P��Xʽz�L}�3&+�e�m���/p[��ධ��Y����4VKj_jZ��M����6��=���j��Ц�t��9�STl�Z���F��;nI	�b�-5:F-��q�J�Y�{�a�9]o2m������l���8U�-��[-WKt� RtU��E��U��8%�bNR]��k����7i�fA�p�x�f�M<hV�����q�,-Wp��x��fw�I��r-�1H�0�N� Zp֊���=/1��0]]�oQ��"z����p�m�9c��j��wa��8��X�t����ڴ)=B��y�٦��y#Sf�t��n�c��WY�g�5����>8�@�K"t%N��E�Wѳ�4��:Fd�nN��5���TR��O�Ν�����\w;���{��E��R���+C���]�p��T#�q�n]t��P��H�f��][4&e�j�Y!iE���I0���e�C�5�m�^ң�ћE���j���]jn]e^�=Hp�%�{�d}l'��{mf����ت\�)t�8�4�9����*G�%f��7�]ǅ8��1Vc�dvz';��y���N<ti�Z����}xK9;��!�ȣ�K�8P�0����'"է�S[B���խ	�;-I0�1.�6�z�����^�t1y����i������}i�e���ҝ,"�U�"Sy��Ӵ�ݏ��ܬ�&Z�����L��}�)���e�{�A60.d����^٥���'���A'fa�f��œ7Aͳ̻B�f�NV٣{ظ$l2z�Z��;t���Ç3��*�5�<�W�f��mi��0ޑݵ�lש���ǁ�e1�w��;.:��ZK/ENp��8�����mnsڈ�����a�=V�9��)��tJ;��}2��o��O�
}^�b���W�X���H�h;=��!/Oh0b��X�]xի�%=��b;��j�.J�i���9OFf�:���fZ�7�+�^�;B��v�)[xj�'{,i<�X���e'G(d�bm��JWR7�Ԣ;ǔ7��Ц��r���;�hސ�Z/���GpV[׫���*Ӷ#�w�hem�A��(�\ُ"T�&p���pEôД����J��l���M���w~Z�M	�@ӝ�6�뫄f�j�x(bcf��)����d9�w.����Æ��q[2e���*��Z����>sj�:����Gz�ގ�\.�nQ�y�����N�mN)�41Cg*Jx�YDN��V���elV�K�ONBW�Е���"���1W)�Q��HdMZZ�v~{7I�W��f��ĸ�[�\/�j�v�`�CY�-�)�rP��o'
�g�xdÊ4
jn�-V\{�����+6T{������͋M^tmr�}:J)~�G�]\���Kz�kgO͝�s��
��-Ř����Lb�n��C��bQ㈲#j���ΡHM̝��m9dӭcE�h�3Zݙ�u�Q	[�5%�̫�v��}�9;�FW~�@A�^��Y�SR1eE�=�`��p|*)KE����[�r^\xT��\���:i�hP �jW� YBD�<�dI|n��� 3���mI�2�ot��[3�T�X(�]���9V� 7�\cu���j�vu�ɵ/mc��:#ٜ�g�w�,�H�n99I����p�W�f`f����k�al��^�Ʒ3���ƞP̓�={"H�}r�eՂ6Έ �u�t�nTt�'����g�ۗ��f���Bw^rm��@���-:�R�m�v	+T�nV>�մ�Ew�8G�����y\��s����t�ٟi���:jK7[!W]��4T��u��X,�f���V8Vm�$}B>7N�{�]��˗Y�/fq�v��,-�ud��A����n�vf�^k�|6�����GB�i��'/���6���)�mCV(u��a<�9���U���ۇ*�kU+�t��l�V�74��W>R�����ܴ�����s�w�DLm]�J۰��RW*�'��֯-�x�3r���P�i�T���%����.����Җ�	���U�ƣ%iޮ,�����a�%NF[<�a�v���� ��B�찱�wS/��*�6����t����.5��/����+D����F�&a��{�Q-S�,�Γz�5SX��9f>�|���Vp �$���.]�%s�[��:�JR.�����!O����J�b{4�O0H��|�Q�V���8�&�M]�.h���7���ፅ3�4���I�<��ep��i'gI�f��*^�R~�7Wٔ�2tm��i��bT\&����qtm�e�y=`�b��݃Ϧu�d����0���\�L���c�����F���s�K,�MUô������a	R���p��l2�d]��u�(4��-p�uݚ�K�����}Z��G�ؽ��LDo5�.I�"��M95�8�z�RM�Wƍ.}�%ʚ��2x+�q��y�}�2�����,�����Wܖ��c�]���k.�켺Q�j��R��O(ӷZ��y��J�����Ô`��o3w��vf��qR�e���Y���-ėppo� jM�cO:��7|��Gq��b%/nu���T��F�ֈw�L�WhC�A��wf��Y[���F����{���t����|��~�뽬f��
Ր�������f�7�ޅ͚�b_,��o:S]�v^�6mK3@N�U�xͭ��L-�����6�[��-l�R�[a���N�a���z�䦖�Z�����.VΡ�mp���Yg4���
��4���xr�]é�A1�&�EY��9�Z�o��j��X4o<���z���R�ug=�F9�'[��EO��.�שR�<��`ޫ���-w�o����i�zk2��9at`�t���U�r=�Y�y[ua����m�+
C��"�<�������V���1�ȩ#ev�
T���z���0��Ԇg<�tz���
�r��[8*F9�F,�:�t�k&=��o읔Ec�"� �v�UĚ��:w3tQ���%̦1o`�S-I�d���#f��T�fC��U�G�(j��^�'��M����^�7��ujX�����_�lX}�L�
�,�,�U0�s��vL�0HY�'l&�Ѩ�)��w]s��syh�U]8�"vA,Yv-f��CT�c�'ad�������}Uze�ݻ���jnW.�/2�����ڣ���,�� ��V��8�Br��fZ��\]]K����bvn�G	����K�A/"&y����/�����N�9�2fLEsC#�l��juڑ/��|�X������mb ɝ�Z��%C��V�I��Z��c��aҏTm��E�2!�HZ֥1X���R����tiή�?����z'�� �Wwhn��61��Ʒ9V��cl�NP��NW; :+��sT4�t`B�KÉ��ћ��&ʻ�7{\��q�WDl�5�����v��b@Τy+�nsy���_f$%�f�͙Ў3Uin�#1ê�,��:�z�����ԫ�34�mq��ńt��.v�g�㏭�Z��.횻�����B�&2U��n�+/��x����bt�J}�+#������w_6fhe�U�.��C6R�wU;qq��0���k����\ݸa40K�Wn�3�=]a�eNl"�1V��E�U��{�d2��l���Ǆ��|����0ic����u2/pP�D������=�x�I׎[���S���':��UAB`s�ʹ�Z`(��gr5;s-v�+.|�,��ԧ�z��y��N�B�j��F�F�+b�v�X�֊�s.�!AfP"��8�-oP*�AZ	S�I�[keN�l(������[����hB)z
�sb�����U��_`c�m9ʞ�����n%m���ufvj.�@5��6F*�J�0.3��/cޫ��[�~��!���<4*���C����T�aׅY��h�UW���Ӂ��H��V��f�J�Q3���w���0'slj�`��N˗�TF�[gA�5���e���fP����ח�9v"�M���h�c(�YcsU��Ԅ*۬՘P�F� ����h8 ��r���R��S�g9�5��K	�%
�d3��+�����Ʋ;��6�庴�Zr����ͣ�GB�X2=�є~QK(�ۗ�W+��K��zYw�σ׼N�{s�1�Eֆ^��Q.Թ7ԝ�\��ZC��Q��LG�V+���,�����H��Y]�Lk�̄m��k��U;�]^V��տd��E��6[�n�i3���i<��pY:�Cw/�s��.X�t�ӝ�.i�U��V�n.m�.*�b���`t4��@��׹��Sq�8�Gy�4%�4G9�#�V�'v��Êv�BŐ��F�ʫ�;��ụi7HrmWW^p���u���nw�K����o$|�1[��ENH[ٸ�X�þ��;o�8U�؍�uR�C�7�.��V���J[C%����v�O�n�zl(.[MWV62�4:U�KbWdƮƜ�)�P��p�ܓ-���$��!��
��bB���ک_�`�N�,�\��St���0�c5�!�@�U�7i��Jڦ:�:uk�N�.�˧��K�)fD��c��rZ�]#���xv��G>�6,��TU���Si�7�_U!F�:r�<�[�û�4u��"����C\�:r���z
�{���&��
�
vfQ������KXJ�h�/7F��Ő��?P��m�V<�y������"޺�6��H�cb"�E�:)�/����D[}%ݳ]��nvj�hI���b@���U|u'f��{��a;�b�ɯ�)��Z�^�����Px�\�4RK������-���� Sc2tҶ��oW�l�ݾ��zz�m�p���w)���tN�]�F�'�'x(������*�eа�/�댙��%c{:� �1Sh�J��0��LD�nAcz��#����}7�W%�� ��g�]lȵ]tΰD�)���SX�2�����ᨐ�}�/������ٙ����V�ᣪ�6�s��8�7�>'Lj�*:��� 6w�N��a�����2�o�d�-��{�3{����ŏ]uЁ�JV8�.X*	\1n c���܌
����u�; �$�| .��{]sT�n��8^N*ܥ�=@N[��W��lB�7ǻr����2h4�V�M��y��s{�g��ڷ)gSD�c]�ݼ&d��;�s���0ܧ8dn��Z�	�f.lt�
>WڙvB��*�^[hs��ʵ���
�1Z�K��jY;p��:��Du�������[-1���+p^`�eU[;d;)W;�G9��!�s���y���L��֝&�����7x�՞�y�/_���p嚜hp�ڬ�f����t� �1V���&�����qΦ��c��S��6�e������ޣs^��[�h�
n�v�)�q�Iz������6�i�ڣ[���s�ĝ^ַn&V���Ė��!�yc��}o�H-٨����>�1�J�v��v�V������d��u����q����a����>��ߵ<�c��Ŧ�*�uGP�i�����iM7,W��
V�p|L�b/T���[bݛs�{��i��as[$��eYƞ�m40s���ꝵA��qE����MP��8;v�:�\ȧ��m�
X��
Ы�%R�\�� j�ztU��^I��oa�{g6�渱*�l�^r(��	�*+Xe���f�ʽޮ��V��X�m"�tζs;�r�/��:hW���L9�'.��{h.+n�b���Q��+}X��z�:t)a���M<�ݗ���:Wh� ֫x�|cs6�3�t�����;�O{rFMA�ܐ��-�8tn�� ��w*ӑ�DE��p�@A�N�Nm�
{���l��2y�\�q�ǰ tI��ǣ&nؾD��B ΋���!��/l�x�bx+9j)-3\�#�t3�9&K�2w�/c���s`o�n4�n��ؔәɀ�@8Н�`}���Of\��߿}��R���C������'~���;���/~��l��f��;ܻ�v��^��|˺�h���:��>e;�b�7cBu�AԞ���y�piz�:lg��45���z���y���h���:�K�|I�(
������;*"��}�}�/��O���"�������O����������8��Ŗ���h%8��l��T`Y4 �Y��X��t�[��z��P�����FZ�\bܭ���u�H;Vr��@�{Vt.c�W`u=s���>�A�aӍ�����v��Ґ�R�	�kZ���ռ���wnaQ�ؔy}�u�۫q77N�WN�Z�֮�l� x�	Y0^jT�\��,.u�=����{����{� ,�gC��"��\koI��ߝ��]��\�rV���ka�ޕ־�=J��e��%m������R�X�;'R-%�4���vҙ��)n�������'�&p+g5m��F�%���5ʇs��:����Pi��ꬁiB������%�ؓv��/ =��0�S�G4�V���N�S��vVE��(gIl��)�t��Yӵf����aYjK�B+������ۀj���{��*���f��+�<S�� �
z��2�Xw��K7z��=ʔ����۶[��4���&�ʎ,w<�>�_iXt*�\��c-��8Q	��c���0s�0���GuAqkf�`�
4�Q�H�T��g6$�)Y����"�A_��,|�����3(��bhoH+R*�7�o�Ql_X]mX��g2�ݪ�����kRt%asl��y{Iv"�ԡܜy;�]	���5��7�����$��mf͖].��:��}1Mvm��6D�VZ�T-h����ս�k�D�!��\W�Y�T�xN�k�a��NjF�x&���f����-R��Y�tʡ�9'(sEm�Gt.���`hq��)l�<�z�Ս�FwAB��1�r����>+3��F�\�I��ݕ|�Ez��r��Oj5�(�X2͖,���U�W�jh6�!@��(o������Le^!]����K��6zk/Y�������qŦ�犱&���!υ��[G0B���G+��P\Nݼ��Sմ��[���[&��q�s�Ŏ���v;e�v�ݘ�RDl��5	#��i+W`c!m� �0�ua]o�nl]�J	�]�ݏ�'���3%�e�Rۤ�T�g)7�j��CZ�jwJ�2u����\8GԧN�A4;�����Y�ހ���P�U|��ܡ��]9kx 
��k�����Yf����sq��(VԚ�왢��|���<ޕ��=U��܋3�d3;�DZ�EN��^���<Z�AW���+���mi��si�Z1�ՠ>�Oq�}�dJ�疢���t����+��D�vw��Q�z�u�7�S�1m
�̞�H%,�T�{�n�]͛��tMqI�<n�M]9b��h�uwpm��%��Y����iu��w�N�Y����/�$�u��-���ݜ�8X�T^�;Y5�ۭ;Φ���%]^e���GwPԃ%����ˬʐј`��syu��t��p܆����9�S���1��S��@��. ˠ�u;�9���ϳ��7�0� ;q���=��j�a�S0_,|�f�mo�
	�h珌U��1A��5�WuG�3tT]�#����p3��l�=����*	ǹ�D卥�v�2 ��ݴ���r���7����
\o/goO�\ܻ� �1���wlZ�N�QI�$ԚV��9s%ZVħy��s�hv��3���8�lZE�I}�[��.eWc����GI�٭�S&��[��8
4;39�s{ۓRlX�ю�U�+N�v�ĝ��e[4����T�璳Sy&�r�t�"8o�-�|CJ����Q�2����˷��MN%���UkE*]ZC�m"��op1�1\2�8-��W��|¨x�:�F�Fb�2��n��S���^m�����]<�KYܤ����������3��Ȝ�*���V�+�/i�X|1>�K��,�1>ׂ��uS\9j��O^Ҝ���*q��G�=8_m5S{9)ڧ`�S�c�qW��d�Ĩ�,����b-+Z��ˇ�P�0�pe�r��8ԌR5��X�S:����2���B��#�Yrl9xvG�>�RSz�rR�l� ��~�Y |:mqO!��J�����gvgo�C�}5��y�PԆ^n腭���c��FYM8�]���@�:��;{�kƇcq��𣀝2��,�J�&e~(��l��n�{�Qжwf�s�S��۫I���Y������E���Gu�����d�V�����\��r���oU�T)8��NA�.�peE��)+V��ٝ65r��b�t+ ����g�un:N��e�O_���F�(r���cY���eq���'�#q���!�k��F�YFɮ��)��:ݔS�w�k|d^s�ys3	><Ӓi��>w��t�Nt����� 6ﶬg_l1�ISRW[��Rz��ZG[X��F��q=��[���م�@f�Ls��_L�e�������ʺ�;{��<?βR/�|yE$7/�vP�z��\M�ju�\�����
�h���׳�������N� ��||9-tb�NW����[�8xYB���^P�A[�]�\�tv�^�lZ'�R� Fvd�]8��<ĺ��m\;nT�v�iN��-e���9t����Ye )pH4��sY�7��]6��N�=v��oAh7[6�b�q<���F̬f'�m�\���ZZ-�;�[/���M�:4��TF��Mk�{���66�ѭ���ۙ��N>�:tXY[$��Me��t������u��O�p�{!ۥ��"K��6���%�r���᫈=afhE#E�m�6r�+#4Wsz�p�,��>�C��=� T5Z������z���.�pY����y@Zl�Pr�nت���i�'^Nƻ�4l�׵�$ƿ��#9|��Tm@��|m%m�qΒ��Hi��q�hw+
̷u39�n����Cԩ���Y+�玦Wa��n>�/�\�M���WK�q����[Ė��qsd�4���fb4�Ev�ov�t8#� f���Z��Kb��wm��H��%X���;Ik�|�1�ϴ��z�#�Ȋ�ڨ�q���I���ŊU����,������k
TC�I���O%�v�-�ǒ=�<�gf· ��ܣ\R]o*t�%��0 ;�'a)��`�F��2�æ�޷J>4��i+Ӌr�p�`�-���>�k�J._uV����C�G����n���l#M�3�����S�έm>���B�m�7���IP�C/L��I��ʷ5��'�-���	��� )��P��!3r���!(�m[�,ݵ���n�b�6��AV�������0���8KUw��\�c�������>��sd�@R��պzu,[]Jwm�SjCr�q��H�'�[��>:�f$:ME��w�m�x2����{��>�}��^��S%�,U�3��AL�42U�Y��v�1�7v�a�� �#G,�D�y]�P9��[5�=�c���;��U+�/�	�9���!]�& ʣ�|�K%S��;�^g$��lfdPum��JM�S���Z�]� �k�w�ʻ�c�&:�+1%�~3]���j룏U���m2�}%ݹW{ؘa��b�X����Q� nZb�}˗%���,M�=�����R�h��O���A���h1�J���^�/�b�Τ`�9��tR�k^v�ot��]�|��l �(Џ��xF���F���0��t�tV¯����QVԕ"|�nj�ؘ�[9��6�;rֳ۔��Rp�(��؟0S�mcǭ4�7,FƄ���̺*އ9_J`��ˣ�$U:��%P�1t�ҹgwA���Y���,unJ�YW�Kt��o���3c.X��S��"۹��ɶ��T�T���8�[W�;& @ۍ�����I�rkpݜ�髠�W[B����7{r���V�X����q���on��͑O%u�K"Q]ȷYЇz(Z��EV6055b�j����шfw7i�u��� �{�,���jä�b��5��#�:�M���5�:��R�c�}���#ٚRgq����t�Lz��㈢�qbf�W�{2l�i 5���ĺ�sn6]�yx"^�u�{tu��V�7eqr9�q,P	O�V@X=�	��x�bs�s�.��E�<8]�ӊ���8'���CU���6�KV�7[1�v2�q���҈�}HMk�α�$�"�h�c�n"��X��D)[n�Wp���ۢq��46uKI�`z��\ f�qƐ�O$F�-�Q/�"����d��S'�oQ�a�v�u�0�Ʋ���9]�?YB������˸�r�#�od�Ų����L<Ҿ�0���#�H�����'�ח��yd\Ap̾z�Ls�k�&b��bk,�q�v.�e#�e���,��j��f"p�J5�����H�C*I��f�e#ի@��Y�Y�%�mlxqRަ�8�Sp���A���^V�h�t�=wΥw�]��xj���T�݆S�Ro�,	���=�E*Q���[�p�}�i��æ�m��9)u'W+�}C�fi�v�#������a�p�.;��W�0�X�e�$I�~�X0]�ֆ�A�P�j�p�nݔ��撱)��]���*į\}��E\%>�k{O<��*�o���."p�[�^l�٥�'}�kE��5>�'դp`m�ҧ0�tv�F�9��;�;Zr1S[b���ˡ�bo��.[46�t$�W9��.��d�b���Tk��!��Q�+�vR�.D�Ɣݤc̻Y}�����ga��։�<a͛D�P3.&��ol�v/~ʇ^���6�l:#�0F�r\��w[1�OXz��	��Y�7[Β(�� ��u��y�8$�<�8�w
%�̮�b��Y}#����#e�Gr�OU�gi�{�⁫�N�=ɓN��(c��B�r���G���UĕoXz��vʹJ��Y��&�Uu��Qԧө`�s���7��X��^6v�p���D�f�qcX˵s��xTTˋ�u���-Cb���r�F�$?��>k7�����]�LS�:����0"�WDћۓ3�ٙV�լ���ZH,F�<�4A�l]GR�h�T�Ӌ0����׺���6s9ɋ��-߯�*.�@����2QhgS¿�+�͒(�][h<�32�T���]�t�VI�Lҹmguv2Vʗp�C��h���;o�2���?B��q�L���C-�9g�6�S3g9r�70c@V�t
��,�7*P�G>����yՙ6��X��b�R4���4-GL���� �x��9�ue5Zs��K�n�Go$Y�O�W%�ZY������L�x�A�<8�h�Ɖaf^�PV�R��WZ�k��ֹ@^.�*�^�����)��ƭ�]�µ�JR�Z��6��V����j�|OS�!��v�M�޼��Q�T��PP���G���G$�;O��݊m�4W;VC�=WA����4F��@�� �1X#R���k��아����2h��Tlm���u�d��\d|r3�oD�J�/���X�Λ�Մ�Q��$���\�O&o�YWp�����5�*b$����k���B0�|ݥ���o��>�`�J�����Sj�Ő�k��d�gʠ���#y��7��k՜�̋gQg{�j�Z��O+E�2�:U�Y��4�sl#��Wf��i�d�yN���4�(,���wcy9�y��5t7(e��ՄYK��ha��4K�+E�p]j;Fќ�i��
��R��Nu���r[{P���2�[Y�)�q_+��9e����)pUԣ�d\�^�z4���M�_
݃r�2,�J��IO���.��9z$F�e�U�7n�ʱ�����'+c�n�[���ФR���M1~fh��`[L�:�'���"�І�I�ç]�wn�w//!�9�pFtu��[�����t%*U�М�/i��6�A�M��L�)�E�
 ��4�v��)��6�ͱWy9�%�^��!G�t--w�f1	�3.tsu��&��U�c��w[�
(�GN����X�`�R#�l@�(ñ�p3��v�Ut���
��p,���x��	\tW{�t]����*�GF�>���9H�g�<����M�[(��	'\�#V��!����b�Ի�KCG-ɔ_2s)+}Bp���5��PUҎoL�X{�lŦu֮�L�\Y�Q�6u��B;�t�'8Y�+�Zp���`�YXm��eM��QmV�32��ܠ�`R����Y�S|g!0����ne�5�Ol�ՒP^:��SA�zvee&bWY�{nS���{As7�lή�+���m,Wԅ,�#+N�w�[�/-�āx�ha2�`]�A7�͕:�r��^��B����#)ð�o��(�M��Ъ�5z2�7�b�������9����QǷ�!X�+*)0б�#��4j��Nö�?�y�p%��\�<I�V���m�+����h�35դv(F��G{@'�n�n�zf�V+�o�ºֹn��*�:ú��o]0���*�����D��8�a�|d�F�]�5��]oY��h�]L=FWW,�1u^�L�Z~�V3��s��B�1@�#J-7k�ָ��xe��j�_*ФՋ!6�����^A�S���:E�۫���[׹]W�v9C�\Փ�ݓ�j^��r�X�[|z���R�'���@yLQ��uҐq�q��w�-�vF,��LǼS�8+�^��&\O\ս�%qM�pc��ܝ�-y	��a�'�	}B����
J���q�#טoѣI��9�β^���o�))��sE*�QLteM�ڗ���a.E���M���asb���4L}S)�Ja�[�T_\���{�=	U����&����1g,tn�$:��Lܝ�=V�b�+6DZS)"
v�JhX{�}���333 ��4~�������?�_�������~���_O���}�=��g���o/ٽ�zX*ww	�b1bS����cA6L�*���LHY3�jː9����)�Q���ҕE���%���\j����'ev����*V3��w��`���V�9��
�Q����Q T3��!���U���-\}��m�Y��]
vu�3�]+��2U�C�m�&�W���ݫ�{�	9�v0��T�����Ou�$��ɻ�}�{/OƖ�fQ��ҳ����F����cP��v9v��n�o��834����+]��qRK�VЅth>��ay�(��i"���;pk�㎞(�;�h<�pIn*�c@�p"�.�7�QI�%����@��Bkj�j���Gb$Z�f��O%]d��ሳ�>��ʎj�}��=�i��zuu�.�uS��	qk&N�]����!	[�Q,��A {U��c�iǵ��a2wD8o��;�o_n��ԑ��J\3A`4�G2�Y��wϜ���o2ᜍ5E靔T&�^gYf#bV��3��F�,f�C�Йcm;���R�'H�]p{��940m]�[��vM���|4H��Cyؔ�6I�,[�TR�S8�s����wz���(��Ns�N�&�G6�j�ma�K)�Fg%����g���X)��*d�YX�'����B�-،�%��I"��SD��:�$N��s�)��1���h�*l5���J���u�#�Yφݹ!�E����39v�\��4�B��(U���E�4(�@���iA_���ۑG?D%"�$� 	-�B0BS��! �l��,4�N$	g�I�Ql�(8�`�D�_���M8a"!?�2�d�!	~j �PH�	&�i����ib0�	 ��xf	��"(Z)(�*(������F���"���hZ(��t�T��R,DCLHSCT�AR��LE��!M �D��L�H�D�C�D$AIKIQ���,E4Д��,M1-�i���)���(��������������JX�
J)���j��"��*	���
Z"�Z"�(������f*���QE-T1(RU��!��������j��"
�h�����j��j��A%!ESUT1USUP�%RQM5]�>Y���m��y�]�ڷ��5e)n��9�Rtn�{�pܝ����:ӥ-�����e��^\���1<Î����[��=���2���
a�Xe$�A��_��~��ܱ�P��	��\��o������S�sӱ�	��^ǒ�08�K�����N��;�5T�st̩�^'��ȵ�zZS�\�*��Fbl��p#U�هb���qJ���ݿ/W�j�<�����j;�E`�9��ՉK�_��v�럟�n��2�L�c�ӗ���=W<�GKռ]21�N���Xb��Q���2�ɜ���yҍkpT:g�]��g����ɟ wOޮ�ײ��_�n�����a���v���νfweZ��լ�"�߸���g����|�ʞ�{W�E�x���D�w�pv�j��}ZԩS���_����A��,�I���ӽz߰5�`W:��u�J� �v�3zI/z��4���$���9q��;�,9�E6k���Q{"�深�˙����ݗ��z����4���������>�%'��ܜ��*奉��9Y�}2f,�/C;k=�)K^�|~�[B�;6�3�,E�h?em
��S��Js;&��f"����Z��.v'����-�:�[.�+���޲�d}YnR��A���;��q�U��Q�ia����|�&�sxM�t2���Bc�Zy�O��L�j�"��|0�k��辺}�*-^�o|���kՈy49d�R�nv�c��39ͣ'˟ƕz�g�W@k��{�õ�y�e�~����cY��_��4�{�e��c5��8�y�A��͜jZ�u�r�m6�#�a�2��yP�����ꗧ��+G�D�b9��̍���v�>�����O6DOz���uK��w,�/���$�
���P��n���6�vgE⪖�^]½���d����d7u���'��m%Z�|������q�W5���#�G��j�g���)Ǵ�l�v-�77����� �yt����J��X�mi��d�GV�.�9�p������&�g��x{�L�<�;�������-�*��a�\@j�=l�n���cl��
�~�a�W�_����xܾ��s�LՎ�sXֆ:MZ�3.dd���4Z�uDl�[���4��5�!����u�a�4�̗|�햧8M�!��D9��+v�V"�dD �Id�\A��*K;���U��G�o�S.���{oL��R�U�2�=��ə������1��*P7k�*�Q��8X�
!���4o��x��$�7� є8��ᵰ�v��:;@��1eY���;�嬎��NS��߇��Դ�qBB�ک��n�7�$Ξ���KW�u�5�9�i��l��<e�2��Fc��&fg�y��Y�2���{X^ޟ��uH�իy���Q�Uٓ�n�;�S�M^��z��L�!�[_D4]S����Q\��6���ݦ�|�Ɗk�40L�br���g���&��kv���wu���`s��\Û�O+��MG������ߣW/&|��y,(w��<�{zc�������N�������74)%�6��_����Oܲ����eg�V9eQ�c��������;��N�WLY���'C���(ܯVcjk�����|ѝ�EF��r����[�|���|�SOe�.�k/�3z�8'�=�[Uy�n��F�Uzp�Y�w�8�L�1��ȯ�Z��<�zq�B�b��b�3�[[Vb�k�-�}���XAHU��+�:utn�\���R��]w��c#�"�X�s��n�W}�:�A����h�yU稗����� �}}��k\s}Ǜ��Ůخڗ�������ۇ��I����i�9L�6G�ww�nWz�R��'�����l�|p�������v���&���dȳr��[Nc=yҷ�_��/?\��T
���c�_�G<��N�5�j���/^����Y��}�z�H���=^�|o��#t�^cM���8^x�1��;�{����9��-ت���Tz��.�.�)��-��[gT�;ϗ���������[y�ye2/�e�*ϙ�ٯY��h�6#��s�������I�B�w��hT:��yVS��=��1�.%��oՌ���Oy�t�1쯷����<Ƈ>PusZ����8�C����~����?/�#.I;���C�^���^u-�������h�#c{ZP��K56@��s��ѹ��@RD4Z�}W�n��er�Y���Ϛ�o��ޭ�<N��w��)\�h����ҩ�s[�"aH�l�N�n�ɼ��zw���,�+c�d#E0	O+[Mx=/a�4�b���u�)�}�踳cT#{��'E@�.�h��ӭ��_Ɩ��ܑߚ�K��C��jFS�C��;��w/58�Jk�U�V|�K�H���^W�5������q��;Qm��4W�����IG���hibTۃ���3-�*sk���j�͍7D���}�66v<��7O���֡������@�3|o���q��g��N�W�� E �w�9ir���yOz�o�����@��u�!����o1��n��ᑪ8�<缱�_ux����{��ȧ���[j�ާ�Uף�Êu������t�ix6O.�m߻u?W�|��o�+�q���@��If{��\����5�:�^�7�sK��_���C��s�����W��X��}��wd�u�ϑ�mi�Gg���WV��Q��ڌ`�;���v�tO!����^&Ni3���L�ۙt+���J�~짾�:�L��~]��n�-��p���1��¸����`S�b�pH�CAK��=�)�-s6�:�X6-�r[�<���횉/��6�,�&��F��{���ѝ�{�����-إu����"k!n�kV7�ܥy����^U�K:�uc�|t�:�����]9�6��d[^m�{��u*����{;>�g=ٚ����P=7o�����w4Ǹ�}��K��Vk9�x�z�Cru޼��-[4z��hn�ݛ3g��a14q��;�-�|�8���$��lpÚ(^>x��9�]���S����/A�K]3�{�G�E���zMg��gg��eO���+Y��A[;"�;����4�+ȧ����zB��Ned̷6�(��J�3�g�^�8�:0��_�5�Ғ���I�����[G�&$�n���v���y�z�V��1.���J{{�ܵu�����m ���bʐu\��g���*��`�����۳���P*��F�D٨�k�?bN��u�?T^��,'�n�e������{郞W���׎��h��+x�Č�8�.Xi��nr1�Y,к��3h�+���л� ,�H�V���ə��o�05�;9n��,؅����@��`�Wv�XU �=���\��Ʒ�w�v	h��p�ݗO���u�TM�Ɣ�Z;���9]���Д�X��):r����SX�U�/��Y��5�������u/`���l��RS�v���mhmD����So���[���&�k��n���/�x{���g�=~��uOPPC4�����Nՙ���q̉���Ξ��ߩ���R�� da�a�|B��z��з��c�3�y�z}�z�&.�
�RjSӑ]�װ��^����Օ��26��������<y;���so���~P�Ҋ���(��׀�ʰc2�֟_�m����?Y~��s�ǅ����3�#c�,1��~�Ƅ��mn�߷��j��ڰ�=�Iv��FI6`�=l� ��g��ۢ6�@
M^�Go����c���I�����y�ʐ�]��{�;7�{|�*~Ǖ�o��Q	��h���`�E�d�mi�y>��/y�������g�g�gd�g;��ݣ��= ��' �1��E�Ce�c��B���n���q�C	Z������O�zO��6�L㎗����	�T�?��Xą�h�4Ύ�c�����T���ȞR��u�(�t2�N��5��l�8$D'|q�M��҆t�s� QpV�<�/�B��L%��U݋+[������u��wKk�	���$�eK���z�r�=�5��d��^{�s�Gw��"83}�R{:�]4��M�:�o\�;Z4�߬�z�Ȭ��&��1�c�mԮ>�7�r�HC���S�c���r�	/{a����WUɤo!��p������{�p�7���C���3��������p����ߴ����6��j�oR�R���N����E�.�=����Cs��g��&�(o�*�Ko�M�q�9q�O�dܸo㝣2���o4��fNP�u��)n��(.°㠟k^�[�n��nx���Eo���M�������g�q��9��;�]޼��نe���F��z���G����yvV��yv���c��0�^����f�M��o�9�s>���;���m� g뀏>�u�c�Z�X�|��^{�f,�w�Q�t<�Q�2��/�qՎ{������{�~�����G�t�%l�-4���9����gt[�![��e����$<���bT)�̂Y��l�@ڀf.Zs�{y�"�!vstҪP�@[s��T������0����#�O&��}�z����(yV|���>��t~�J���ތ��W{�'o�׽$�Be�E�������̹Jb�������� |bH�OW���M�Vu�����7�u��Uw��Q����9�7Wd�/yگ\�����}�ΒO)�;|�/�b�����SOwm���|��^�����w�ޕ"��:�hU��[*Z~��3��ю���hz��*�����K��|-^�iyw����,H;��о2GHc�����(Iʘ��WA�En�6�~��5;�����'�A�><� q�O�}��d<d��\ws�*�rf����3�S��I��F���H��>�l�4��k��sbj�X�{޿z}��j�,+gx��oW���O�1[A׏�͵��Pa � 4ꊸ�v_V�p��3�PD��ǝ4�N�&>}RQ�U��{|�)�!2e�%jKm�Xs����U�(ٛ�`gB�e$����>�'��}��S�y���x�[Yx�6N���G��@��dTe�;{=�%��ʂ�M)��}X��b�`{�V��BCy����- _8��7cH;4d���������5�<�����vk�������5k�=�WP��(�z��i��2ut�sI�'OV������+ϗ�="ry������j�K�˝ ���z�b���K.����χ<��ٶ	��(�m븑�!�|�[�;��L5�^��',E8���9�G�ӵ���>o}�9�<H�c_(�Pt�r��O,~gԜ�`l�ϪL�[e��:e����ݟ��h��TJ���Qnq�ʶ� �P������������S��+uCmY�Q�vT�V�4�l0)=o����գ�U��e/����ƨ����5�5��}�z��%".��zh��/k���,9^�e��>��>�9e࿂�4�/�<��v�W^9뾨Z�,f�AA|��'m�u������c���[�p���x��^�g��������}����}��o�� b,��7N"j��C���B����t�)ζ�)[ʋ��r��q������m>�x#��;W��l±��|��;��z�#��(c�-�X$��9�k8����M�ssO>�w��!�y��6 s_W<��t[��x��l���kps��i�8�q��ڽ}��$�u�sqfg�7���	w�ά5(������`'�4���a�+��jr��M�2'wë2���Ft<�:[V�Ec��Y������n,�L# �3.U�R����n�y�l�pr��"D(���ƾ�4@�Ǆ�F�'J��m  ތW���ˤ��k�������uպy�Z�*��9%&k��V]q�%��vSa鲥�}{�m(������(eMғ Vq�ݰ#Q��2�]��^slJ���X�n�!�9fu�M�2����V��V�Y*���c$ND�G�ۓO�wsj��LK�ʺ� ث4���9G�.\f��u��EZχDV��	�]���Xxw,�r��C�n��j�9\x^��/�	��fUT��u�,)�qxe��� �ۡ�4���6ޝ^��@!pt#��ݫm���m]`۫*A���T"f!�FE=J��/�|�z�J���5]v�T��4=�x�Np�`�����-ǳ����q=YHh��j�����K]Ύo[#Ue�
8*n����9$�f49WU�4f��o�f��������m�Ҏ�X��s(i2��Gq��E)�P�Up�G�Q2*;ۍ�1��Zؕ0�m��Ǉ�P���ב�C���	@���6���cØ���R��N-<.������Y
Qc����KeN�O6W��a�����}���r���<zX֒�ծ����X_=Q��N�.�Ӡ�	�5�ѓC�+U�w	7T�j�ڻ�+Y	Ws^�ïs*dj�@�s{k�Yw�]|��X�1���h��e��S���r�VB�ٍ��9�X�l��+h%O��E����DE��k�+�F�� 5؆s�e���T���)�KTt�DT�xs�j8�#p�yF8T|K��c<hT�ҵu��I
'�S�O7^�o+,tC��d���l�2�,�p��dA�j7l�@�.̈́Wi=l�e9u�$A��#��V�HP� ��
�.;�A�5�{�ݼ��fH�xgm�9l��n!���1�J�
���W\�	�@��$���Q/�sf��أ�5�t�J�}X@�bt/�Υ��������I/�����N���ϮrVl�$�%v_��Ozٛ5���	�;v$����+�h��Lػ$�VQ�4��v�k����Y�ę8���V]��Q�r�<�En��f�#�[���.�W
����:���dk/:���V�m7[{���n:�y�+�:�=v	pDv�����l�4�̾�s�S��a�Zn�ک����(�P�mJ��55Li��;͈�윏I׎).�$�m�s')_��5�-%D�QK���5EDRQS$�,UMAKDL�1%4UP���CMEQQE�P3-ET4D�$EUUE1P�QU�D-UEUU#N��@EJ�UMT�QAA%3%1]F��m�JQELTM%CN�5iqAD�U�Rh�gE�:�������4j���A������$�UY�F�Q�h���M�D��*�tf����j�F���Q:6�ƪu[&�4h��նvZ��#Df#a�,U�ZH�FtV�M���d���u�1�Zb�����Z���ch���;�U�b�@F�5:"k[;E�M�X�V�����ϮWֱ��-��U��)�r؛ �xfD	PSw-�s �KRZsw[�I)r�ӁO��(�V0=�����=]�b�}`�~:hux�����F�z(��Jj8G�)`�Y$VQL�P��滼�Z���L�2���?d�B�/z�"�}��>�;N�Y�f��/�(x����d�BpX���ڨ�Yyڹ�ų&�YS����E(?���gfu�zP���!��v����,�	Ţ�]N	b������AA69�W?�*1��^O�g�$��e+8�>Ȃ�6Orv�y�5�=��l8�eo+"���9O�K2������<�)�ǫ��g�j�����L�#C����D�W� ���R{�ZY$�8�<opg|�q��̆�dܪ!���`(�S��?���NL�m��L�A"G��Vsd��?��ϵZ3{�v�-9���[�I�>j�O�1H���S��`��}j�l;*���*�J�y�+)]͎�f��@J�v�r=|g�P~R��%Q��%��T/�,�oj���b����teR��l>���+C:���i��|�X�̾�A��p����� �QB�kl�۸��M�
$���=����7�z�r�����*�D�j��i��R�\eK��~@���<0�Ĥ��䘫���D�{��w��o�4�jO��	h�!�diǭ]9�#�]�$�B����m�t��F�gWfL��V7:�wH���#V�ZM���VL���m�YNh���/��h�vp��9���n�BNո��t�
��&%��s�������a->>׸AI��~+(���w�ό9���5/�R򟍊�<󝪅��{!Z	ܫ�
���~��=}},����ۯ��0�H�Ƙ��?��ǆ�p �T
+-�A�Շ��&�@)ܡi)L0��:z���\W��sP;l��(����p�/F�>�E�ދ�޷���%锸�cu��>��e8;�[ j�Pt�g���0n`7T��4�T��㨖�#��$?����bʹv){��9���f���ގ�0����S��)�٣��q���h
-ָ�^)��㩈H�a�zڜ
��ˈ�ެwhx%ݽ`��ש�`�e��6��&��9�F�i������@4�v{���/�f'D�}�H�`��XjjY�-��\�,�R�;��f9��l^����v3��z}�����Dz�F#k����7����#��9L���Sߓ�،c����{�QA����d�)����x;ED�7�fm��G�^o#���P��1��A��1E�+�#o*��z x{Ǩt<�uƻA٣������ml����T�����'2Wݓء0N�~7�Y*�ԝN��s�zkC�1C�L��=�>��ޯHR�H]V�r^���[�i��gN�(�y����ب�M�]����ć��v�uo��w�����e���rW��k��D�e'_�pX=�qR�Dj�4���S�,W�֠-E'�Ô/l%[��m�]..�ab�o�aɢD�ޮDu�#ɯd=5	pgřu�1gܒs���S��<jy��׌vVt�m^K�u�әA(9S�6[�m�2�
�׆!��6�2��"�X���P[�R{�-�fKÐ��9����P%W�Y�Rf�Ta�RA4'���0�u�a�/�ތ�щ�Q��;Me��n���:�*�
	T��#�p��c��#���B���d����ƙY����*G8�֝�~�o����s^EP�4e��\��FK%��q>f��\��S	$���IZ��9�!�	�}9�:Tt$wN�B�&��~`�J\n.�N'�qh��\�넋0u�ّ���zOE�8��_C"�gn��C ��mb(ޝ������^>�J6;�1qB�s\?��w;��u�.�gK���u�٪��C�b�Y٥� �	��־�sL�ׇR�j濅>ڸK9��wي��36������u�}�Y�����^�DYE{����L9l3�����Q���0�f�F�Kc�)������)������?��W�y���Ǣ
�]ijb��Գ�I=��<�{N��5KB�%�l��~�K�N�����V��U��Bt�cZ�N�ۚٗ�a�k:��Q65G�����L��F]������d�*h���#��5h9�W����ވ�r\��Eʳ��ڵ2��>kk��	�O�R�K`�X���h
�J�ˉ�a���S�=�0�m"�,H*m�r�hNC�:�N,z�[Du�������ZcZ�&�e�l�����E��)��ڦ��t�~B��BD�j�w<���5e�unr�U6n���w�7���+�f�?�TC�Sq��һmn!�Exڠ��J�V8x���f���X�s��L�����D9iwƲdH��P�Z ����I���1��(M�8�׈m)�=�@ꊶ�쳵f���z�%����/&��$Uj&QC�ψ�v�	�+�6�t��`��6�3�&�ad[a�R�u�����_)��Ow0*��F�|h�r�0.p0��4���մ�����VU���b%9`��l�J���ޣ�rjr�05��yv*�^I=z/G`�N�|�D�V��j���j&)ϝE���<��Z�Мg����foT�&ɷst̅Hg� "!>�]��@��T�Cz{	�D����%���
(w8����q��Z��$�63t�B�n.O�
V-�u����i���w���v5�BEv�R�d�7�;jP6�6��Z�f;��֔�d41gP�3�et(�cy�6uI*�n�� ���n�s��Ij�<5�N�a�C������%�j^�3������sק	5�=�V�]�&�pgl9X����^�-m���YP5�Qi�v�)k��-=43q�X���V�kK�zX�)���^c�Ly���\X[�D�i��y�ϐ�>ƹ�4)��r�<Jg���T~���2@Z��P��ʴ:��� lT+����F�_�V��W.�Y�C\��Ƕ��{-��Q�l�p���"λ$5��G�[U=�cmK}�o�)?b���Dz���{s�d>�dc.{ �aw��xh�����M����,cɊ����m�\�|Y�>�5ϼ�b$�W���Hq�v��x�^<�0HM���f߳��'\ח��o����\�J���%AOSQ�s#�ۙyw-cx˶�R�h�,�T�nfU�l�K�!�6���^���x<� ?��'�*Y�~��Ta��Jh{eIu2������s���m5��fW{y�9�/�-�3��JI��3���7�F3*v���>��Śf"�>BY�C=�鹝���BID�|N�&6�Y6�uD�޸�3|���I��"�d�� ZE�EQS�a�E�ed������@�]�����QR���*E�-Ӽڧ�it�ܾ�Z9Pni�[�鼮�!�ږt�8��C�lj���E,{�����7�&�&C|j2n��Y��6�GTݹ��[[)�Lo�Dݼ*� �L�4,��c�b��$�
+	�Õumo�&��+�77��p��x_�Y����b�
m���=��/x�.�׸{Y/ihD�h�e�#=�n��4��q�6_���(�����J-?�_W�ʠ��n7n{ė|�{1��y���X1������� �+!�;�F��TQI�_ܢM�2(�����]9­^�Oß\dp�+~�C̯�3�xd��;\�r�Y��N���d��:f�4A�����[�@�ceqY`ؘ�0V�����0��E���
�r�P9y,��>v>°�ЦC��/^�s�q��}u���
&��C5�V�q���Q��Ŝ��b-9�i��u��<�^�Ў2)�@�0��<Ξ�غ��,Y��k�����' t��壃+;�3ô�kMf!f2Xu����ur��mi�%��q�F�1�d>�z�Q���0!l6U�ڳ����0� ���&�8潑�3��X	w܆�wx�w�%�����A�Ʀ�]q����rD������G��K}�0u �U���.���P��]ǟ3^������&�2��/$��|ZT�*���Wr~�W��^�r�{������{cr͞Ʊ3��rƎ���X���L���K���U#� (UK؃�3�+�U�;>:�mM=�r���H�XNi6��|NŪ�'��:����#ݛ��Hɔ���WL?��[r����x{ư�!T[F��Ȧٲ�!�)�6"��{"�2\�5�u#8Ϛ)������e��-�;���<+3G;[�N�r�,����e۴- yۺ]b��(��~E칳"�	�)�0E�Û
x̴�m9���w8��rA��Uc��_��h#"[!��I/�����d�#� pk�����uV%}�,�e��05�W�4���e}J(�J�Nh�*��n��l�V�t'U^DEi<�rrg���0ڷ���XӅp�W��a�W(��Ŕ/_�T��PyҒ���ٙe?�,ۄ���H��B���,���M�C�m��2Z�J���ۑl;�UI�&V1����Z�[�b�ԍ��ke�]�f@�*M�a�I��ek��f�]kO�Y9}��	3b�N�)m���u��7s�;�cl	�~��-��_�T^� ��I"�t�=�ظ���b���c�9�7Cϖq����b���C��y)Z�\�ڋ,��*<���uz�����l�]K\8�<�S�a��q�'�7j�4���6���G)� ��H,��|���4=�(�	��G"CE-
.)�Lё�iQJ�8h���w9��Q���-��[�#���PU���Oo1_-X��ʌ�WۼȢ �Z�B�[Z���Ѷz�u{,��ɖ:���b^�	�9��ƪ������9���ݛO]w�*�� �6�H:��%����S]5L��2����0 (q�ki�����ZS���Y��\J���<pY N�=d0�r��80t��59�TS.��-�,*��d �%�[&�6:��^�"@�J��k�!q���Ȝ��4-pgd���z^��\�Zn�M=/���'17dD).3���Ǜu�+1�}a�U���:_ȋ�D���D�jp�%�>���b!B:4�^�����w*���?YxY�����7�e�oՉ�Gm�xSjd<������m(�S����z�6E�UT��wAN��Ρ�E�X�T���m�=t���ܨ^
+'�"�1i��̥�'�X�N ����G3�C<)�RޣB2=wv�Z5����)�_E�x�\)Z�`��r-�2'��i��&9�[�3�d����Y���"iAR�?o�U7�D����	���O{����`gF�Y?"��O�����P��mNT���1q�j�L��"|�/#�U[ kEN�<�Wa��Aԛ���[���{W��>j넋��'��b��JDu��ӵ��@���f_��.��Q��V�=�[�嵏J��i�'T�[/B����g'G��������4�xhV���馊�9r�e���كu����5�q.;0�u�5y�fن�u���ۜ�b���۾���L-�Gk*8­��ti�2vS�/g��}��~�\�.�#3���
%0�2�n%T݇i��(mJ����q�xMZ/*	��e�c{Jm�*6oa�..Q����SM��0�gt��H�F1I텭WI��n�R��k�sL�Y�J�oo��B١�Q�0��2�.ɫ҄&��	�v��ib���6_Y76�*N>�	���h�*[��&���p�g@�ѐ��s�K���6�W�%��;U�z��X�	mr{�:s��_3DbV��(�i��PA��[�)dV^����F����!�'�F��z�e�F���ԪX8S&�̢��f).�����s�D�b�9nZ�m�	ޟ��?�y2�|s)��H�����=9}��&Q`�����Z6���>k�ƄFkj0i-`f�-g��I�*��X'�(��+�gl^�
/�AOH��3���]��A�":���H���C>ʻ��=.���Fc���
�(|��Rbz�ls=ܬ`k"��
w(���J�[�a����5\>���ˎ�򣈪�b���/�� ռ�7�w,C�V�-�6��	�����R>�Y��*�����ѭ�S��`���|ͱ�[�ه�g�H>��������{t�6|������D�d�ly-�ݏ^]�άxL�@`}����2��F:�P�v6-B�4��>s�+�Y�:]��ٚ���6�2�l0r���F hu�������}�7�=����y�����ܢZ`	3���f	�a��Pږ��`v�wA��6HCˢ�M;����0B�펪ʅm�z��҅)fg����]?�r���	���Q�;y�MG��\M�%��1z��g���#xa.���F[�+�Ifע�i��մ�@3�m�1+�F�|�py>��c��Ԅ�R���S��:����ic�a���v��r��&o��A��O�
I�6G&���3��*����y���A"a�5��9p�A�5x��q��	��-���{0�)��iU	�3�S0܁5}�{�]!����"�Ⱥ8͗ث�Xu�/
I~J-?S����[����@۬z76�İ;!�u��9����*�;,��vZ��J��d�"=8=�E��.0���l�b���GiMJ1��"��H�KlCM��83%vs�0H#��C1�J�p�6��:wC���U~u�����[6c($����$�ZF�`��r��˼�O|��݃%VsI�"�����վx� ��v>Q�����~/�Թ$�5�������l�}�^>�O���x�}��o������p�����VqT���䷞Y4�mr�>֫��9�!��S��ƴ������2^�w&u�H�br)�X#.�=�(���,b#�f�]�0dU���s��=�Y:Jy�3fO竼|ڿy�ݹoؑ���7r��T�2Rs��}0��F��g5E.�K&�œ��/(�urFR|�!n��m�̮2N����0�"zZ|�"�qVe�Q�<YaD� �-Q�S*�:n��6K��Q�;�Ed랽�s�dT����۟h����;�f��]p}$=+Z��)��S���\���1�n$�L��jj��i�4D�aWqJ�t)V&�#ܼ=@^�m<��4Ջ�;��'%��K�N��{MV�� �n�2�T����}���u���%�,��~dp�k�+2Ŋ7��������D��goh��'���b"�\��8�+V8��(&o�;&!zo����%�E2�n�H�B��Szb�On�꺝����/p����=5�����Q=�s�l�N;��'�j��
�#�Э���5���[E��#��J7�U.��`�O�D�Q�Y�:G��r2��1A,���u�U��A`����Knqzoy����M��4Q�[�X��=3���/H��O4u���x�ٶ5���KSn�u�KU��y��)W`N��/-�go.	L�*���'(X}�ڸ\�e���r�}H
�F���)YÜ�Н�z�]�ޱլ�����s캀Z�'�ņA����}y���ƕ:7v/�1�K0A�����l�d��g��'np��N�!0ryn�@KK�5�C�o#�Pe\������� �0�\�(���\��ȒfM�7���6�@����ua�`�L4��2ۆ�ܧ�;���d��Q���y.6�P�'i�>�gPe3�<�u滳d,Mڃ쬦���k��Nܠ�:�"%md�ϯ�<�6�B!�)���:�뷿-K+R7ڜ�&�=J�ݫ.����w�͠�����^aJ%��y:�aI&��u̒���� 7zm��C��3�f�Be!}�p�CR���5g-�|���+hZ�����p�75d6{)�5�9��
l<:�^���Q塉�d�ȧL8�m!ә����N��,Id}ݓgAy�ED��FP��c�
�8Y��R����eL�2ݓ&�aiŢ�3גs׆�����H�[R�0&�D��8^bD�ƻ��.��l�UY�3x�,O�_	�\eSRWa��tkge6؍�	e4�LWN�4ic_˟+c7�����/��W9pǁ�.���oA>�k;��lp�z=$�f��V�GIiT��+,��1�_׿mE���VP�b�!E���:��5]r�e)��oy^��Zfʵi�qF�M�[4b難-�p^�]��ux 5&�m��bZX7ҷ-���K�s,h���
�<�Qa�}�J8�I{��wP!7����{�]7=�Y�SEn֜�Z'B��
I7���#���0�7WB�}�~ERH�
 ���փ:���Qbs�u�f�Y��i�#lbV�&KmQU1I�EkQFm[d�� �Y"�g-�URb6�(���&$����b�lv�G]:*�j!��(�����SFڪ������I$METPUDlb4�"���h���&��v�ITR�PDb�����֤��v2�6�Q%D�PutLE� �����1QT��*"&)��*h�%D�V ��������"�*J����%���b��j*	�b)�h�������������*j�Z���")��h����
�(����M�DԅZ�S0�D�UU]�E5Ո��*"��jb����j�
`������"
���i(�b�mLQ�-���{�Q��v:�d I���t��y^����&��T�͙-f")D-TH:֩�ftĳ�qؕ꬛�0�i0���f�n��\�FvR! āD�ۄFB1ȈM(.G�@߇�����n��m[C�Йv	�s���\?���_�yԔ	T�g�T�:r��=�&k�����?�����HM��-2j���D�����d��,�]5	p��{�y��C���N5#"ۭt��Us���a�q�ч��8���XH<F�)���s�N?���V9��ͱş)ݽ9/��kL��c��n����XZٛN+ã=����˿()�ň6g;�N|�����Ǵ�(��H��̧��NSv��&�Ȧ�/�R���&�<S=�#S)�s�ge����؉=��e׺�ݛ�u����^8���%	P����f����yM��ؼ/��/e�λH�Z}��64A�}ܤ����]��/V�ڽw�ٝ5[�A�*���� �77�i)�Ki���:=}:Af�J'T[���V���^�܊�"6�K�|��a'T�{�K�(���\���S ����2�3�Pj��ҏz��ƅ0�>�:���m[Ļ]���W	׋�a�/Ƈ�����+2�V��g�=�������qw����H��2=7��2��I�i�](C���~��sug=L�M��W攑R(5�M D��C^�xĿ��A�;��D�	Y��W����c�׼�Fٺ5����:̻���x�u�s�������ok/��f�ܶ.�&M�6,����ʺ�3	\�C��f�/�WZi+}�o/��0�r�̅��&��wG�x}�<���*T�/�{�������е�Coܶ�^���SO��F/�B\��� ��9��m­�C�̭����3.<�C�L$��(�\��{ed�V���F&<R��G�af֗�c3cP<'I��ɧtSɄ����_������
Ԧ)�L&\C���-q!r��_V����y'ܜ�֫�fP҄�c*���r��<��^:��U�-#%���'53�`G���v�c�g"�^��/�A�%�;��:Xu��&S��@��b�R��m@oƟ�_�t�6-���Z�;m?�'VO т��C��Ml�x�0Ϣ��Tt���	%`���>��'{�O�(���Z��ˁ�{�3����S6�y��y��}��'@���&yT��;�m�q�c�[Κ�傌N� ��T�;�P�	�(���/��l���.�m��o��wc���-o,A��B�������Ş��3H*�3�O�R�|Oζ9��矝j~��tӈ��Z�
i��	Z��K��-}[���A�H�%M�nQM	�\�ؽSlgs���5�(�@��ʸ�ӧ@��6��"�W^۹ڮQ�+aX����c���UN���xF�.��|�HH�70k��^f�}+,5���Y�����I��bk�\�bk3����dR�Iԧ7���V{�BX�o^!}�1�J�������97=�g�p���5�����ǤF��0�[�1���7f[���X��N�d��$���]�\kQ�d�����־��h�==0�?:"��'@_|��x�j�j��Ϸ~��v	��l7nD�x	h��/���֣��ЬV<y ��ma�~�F ���4'u�<���8�A�_}nW`o�²4� ��[���I����œ�_G�@n��r��!����[�#u��	�#!Tb�BcvUSs�����ŕ����ofcF�����B���_;ҧ�����l���B�R����b%9aa*��ܕ[q�8}�L�%q5=K"Z9K)����k ���ݹ�-�쀛����iR����4+���ɨ�1-��d 9��X[<k��>��#���T���҇�ouP�Ur~��j"k ��\�ƪ-���g�|z��-��%0���Ym�X	�M�u2�#qQkc6���p�������1ʙj���A(�层���]��xy�)���1ؿ��iv��5�nv�]fo�.e���S-�����G0l�Iv��3P���es6U�)�Eu�m�31ͬ����jj��m[��0emaRiGI���xŘ�����Iofnj):V�T����[�o�zi���vF����#y+�w����{�ׯ~|�����B"� ����q�Aᖴ��N�[$��i�%�����%�5��6h�#cPa�Ii��9��EXތ��2�Ή�ol���g"N���t�4���>Y���l��0�z�~�녮b��m�̛���kN���5T3J�5��&�u�I�/���p=C�����LF~�h�fh�!��ɡ�v�M����a��椈��(
^� ��!�/~��}�}'QU�%�>�����X^�g��Cf�.�v��vB��e��M�Áb�B����0�
�ԵG��������=���wnOn��k,�!t����p��Hv/�0��ro��3�Y�2��S�dQ��B,���&2z�N��0�2yU�҆O��d�������ݎTۿ(�Q{�/=�p�/��yƚl���Y|�1B`b{�����7
��8G���=�s#+��DW="���z��k'�a����q���a���>��^0f �so��k�y/�b�M��ǵ�c�&�'(�vA&oa�cL���XPb��JR���ef5�y�J.,�R��¢���G��W�{�Tfp2Ǽt��Zg4��I�瓖�٘E�z��p����Z�w�ebS�c}�*ʻlN,&Y]͋%��*vqk�ŷ��ލ����2�WA��b1�͓���Ίju�8�ٙq��#W�rݍ0�W��h1����6�]hjT�%��{��7���*r#1��4U� ��P�Ｒ��5�c�v=�^g�a0SO��a����i�XU�5x�n�B�D��m�s���М&\��T=Khu�VP��@����Լ.z�75�8Z�n�8�f5�laƖLF�{���%r���(�#��@���wx���M��Va7w�	�v��#%꟧����{9�)������О�A,���H(��TI�J����c&jݺ{�u7��i�P�EF�/%�yi�Ξ4.�J��o�:z���=׉�栄���)(.�cN�4�U:�$�THM/HDS46{'��s�wl��fq�<�t��z"㑁,E-�a��/��*6�sS_<�;���zZ�Y�P���F��߲���G��f����q�r炪�)��ܝ�0Vѻ�uZ��0�Mc��b�Β~�����"�_+�|}�2r/U��t�D�=59;�O{h�7�T�1��?��oS��jRm.M��e�k�w���y}�����g�U���p{X�ETJg4}��Q���m��<�Ջ��0N�z�.8'���;r�
�]�W�Z{��6mqÔ�0���dS���=��6�!k�WLѭ�J�.�I��-��U��h��� ��Z�ќ�gq3�����5��e�w�/�PwJ�>��,��[����������W+%S$F�=;�^��qmB�Ә���r81��6�FD�V��w|�P�'Gl�y�j*���c®2s��4�1�'�WJk�W%��}�~�9k�)z��턲�l�w�k4��Z~��;.���j�r9�^����0�1�S�ɍn~xMm�z.t��0d�n�[����_|w��/����&u�[��H�k�B<繋H��9P�S��c&�;2��\�
8�؇}E��|^J|���^���-fP���^���SO��H��ˢJPp�ǅu7�ry�jN�ȇA�Q�ȣ(����N��S~�%>�O��V�^Xp�xàNY�mɬ��s�׺����ؚ���̰�1E���+����I� MJb�T�G<�����>��[oY߅�Ͼ������R�a����νo<���D�Ӧ�\�<ü���`1<�&�Ǜ����;��wMl���p��KP~�(�Vp$w����Y�'	T���.�O�+�Ҙܦ��P���R��C>�N"m�F-T<�;�1����Y�xa���م���=^t�ź:_禇��eY�.�rܲ5֞�k��4��:�������Ԡ�����\�6T�\-;GrM�k91ѻ�����@���Ŋ`�G.р�kl�7���4N
F�/;r�9Ȏ��1�.��ݵ76@���k9h�c��(&��:�w�=� W� !JR(��_X�����W͕�L��O,a� X�f�Li3\�Fjc-pg�cbr�G��)��hV�X�����i����f[�A0Z����}��W�X�c^�Kϡ�^ tdA����eͭ��m�9�['��I���c#n��^$�`��MZzs]�m�z\��N�Z�]��!u=��1���К�DH�QqBk%��lȆ����'¯5�����d�C�!��J.2�6j��O6�4r?7�?Ͼa�~��W�۲B�~����P�nK]�P��[�/{J8�q[���q�w:n���T�j��m����A�9l��2=[2,W����Ĉ$�L[�ͭB���-j�[k�Ьy�����	M  C���z�[ �w�E�c������Գ\�0e�˔����*Y?X�4�l�omyb�bڈy���`���&��ڦ~q/�q.y�;ҋw� �YXb��9ఞ3)�璪e�pj�n�k+QQ�0/�=��yr�8���.zִm؄�Ly�!����G*E��"S��M��J���I���~=�2f	��_���MWm�֖��V�r-�h��L�jY�7!�m����VC�UH3V����w�> +�w3a�mV.���$��+J��E)X�a˝����K��|=�KɐY�`��3"eηk�<y�@ � D*�BP��{���JֺJ�)�cL��[T���}0�xAn���������8�JJ{u����2d�iM�3|��>��'�'b�<��G����o妧3��cq������ٺ]�����qc؀<w�.���J	fy^�l\����=Ff�e%�`�Wڇ�D����z6v
�ޑ[�w⫾�0�t
���<rj<�w��^?���iQ��`���X]�'a�4��f�lܖ����[MV�k�.�.5�����y4)�k���z:<_;����f�p��v���`���"K�kaJpÑƸ��폎��p�3{�������4��3dz�d⦘Q����\r`�mk�Q���!��&�mWf��:�C�3�9��.�8��V-��# �誵�+�����津����-�w62���Դ;9i�T ��۹��v]�M�C��ӎ��3(kZ8�0Aޗ��G��Q-0$�B��3����Q�n�}<�ue���4vr��������;$�ӴW��k��y�5�Z�׍I�ɭ�1�h%ژ��s��x�Y�������ngl���3�S 1P�q����t!�4�Y%mC+泑M������7��f晻��o�/��sO�v+��Ǫ�q���zg]���3�C�$���5��u��qC5��M����w��M�����}� ��
B�ZJ�( JA$�A���{Ͼs�Ǫ޻�޽|g1���A�U������FA�t���g����G���T�����\RK#�Zm��	��bl콱u���|�-޵���R{�Iױ�2j�Y6�K*�l��2��h��C)7���RX�:�=�(���'@����'�h��ۋ�k��=�)?_�#BۅCuv9[�o.����lA��]Onc�h��>�^�&B�D]����1G0�����D�Z�q�T&�Jʝ���[/�!Tt����+�FUհ�����ע��A���;-C�ǥ`s������ZW���xP#N��˚�����M��� ��H��I��@��c{-��v�9���n"yd�'$,�k�������8��"��5w\��%���Σ:#�裔8nv�3�`$[ ��u��fD�皁����AA��C��v�2)�~��hN���9�����TI6��kh�~|��57;�uT�Z%������_<4s��[��`N?Za�5�ߕ�g�u�J�ś�ofy��Mҩ�(�Ɓ�0s������tC��1X�����ԡWS���g�z#��%�C�@���G-̨��֌��ݛ(�t�o2���+X|
�ꞩ2���
/<�Kh���M�lV�ׯ��qn�����z�O��u$����F9�p�8n����R΋ґ�3�T0a�i�:r��]A|�ŕ�c=O1n�뫱���Ϗ=�4 �J@J(D"$ȢR"RD����(ЀP������������~�����(F��i0"@�� W-�p���o�ӝ��h��]o#[]��)��%��=��w���/�P����Jadqb���v<7�1X���3O�o��
�˪�<�����ml��V����}�?�����T9D��T=U]���ud��S9�5�k�7'R+�)����%�m��n�������7�ty�F͵�M#�_c���r���5��4
w�{~�h��� ��m�R4)��� [��C���D��虫�QR�(u�2n/K_&�c�4�G[���G�ʥ���P�)E#�竚�A�J�99�W1���Z���
�NQ�$nPT)���NLG-��5SOXi�l��5şr��ޛ�sf��;+n�\T�~͹�M���nXV=2�`�yz�CЇ;����*eT�t#�5���{���BL��DM@��N�)��kQuߒ�}����A�X��^���������w�qS��.�:���2W�A�����I�/,q�%=�4�X��ѭً��o��z}>�_��������{��O������Hz�����eN���b�J�>������=��዗_�oe��
�i�n�G�=ǝ׍ҏ�U�Ld�hL_��Y�vi� ��_n�h��-�$�	��[D�4eI�Uj1�=���9��\d]ౚ�X�˳+����K��/i�j0��o	�Z�R�g
͢B�su�A�7�u�WV:��Z��[}�	|6�q5R�0�tq������&����s7oJ��Q�c�Y^m��h�������V��aa��v��"LG�fn��Jj�p��t�|��o���G:}���b�Nd��T�^�&�+0��"n��^�Y3hgD�wm�������ac�h��a�W��\�m�g7��f�]%!��X�q�3�wV3��!0��!نW(��fd3N��b��4��Y����q�D0u��,��� ��Y ɺzv�8����؟ћ�(�y�KPB����������!�WpN�T�le���~�!�u�Erɖ@[��X�1=��-�cUt�΁�:���P�zGL�j�u6������Sr�(���W�T�:U��f����8�I4�me���X���5�d"�D���|VK�{�S�,jK�M��y�V�E���͔&k�����薲��9���A�0�)mjv�;�6�j)�LXzn��3����x*䃙�����Q�;/��i|�-J��5}��v;(J���m8��@q$�tήup��{P���֓p?o>XpS�o��>��a��3Nb:W�[3�:��'S�?����]�
��7Զ��G:u�o��U#��b�=������ �u-�I8�u�GcI�wur�b���qj��w]��̓eP��H9ѱ<�V;��P��g'�)qL`\�l<���l��AuK�Y�0.�u|��(��;&���
DF̳�fr�V��Y�Y�l�ڄ�36�+���6̊˹Ko�j�j
d�Y���R�}d�j�q�Ⱥ��T�V�̗o�-��MN�.q#w��<z��P�ߝ���:J�������9����u۫a��(��R���J>{NSɇfѶ:U�;Z�m�U���>�ܴ�!�y�T�sH�;s9ܾz������y����F���]=�3��b��.{Χ4��ٓg12v2Y#5�{bA�Wa�:`���y���JM�%Z�}��F��1W���y�kr�E=N�m�����j������bweE��;�i��wznS<T�Z��Ԃ[nf���!�k���nናg���p�@k�0�3�$zu�v����p���e��OW54-έ�]ۉ�o]C���K��T�7�����sY�֫׋fB2�1�����X�\_6&6ro9��#��$�r�{����DSSUELUED�MQM0xɤ����� �
""*j�"(�b"��DA�[b"��� ��f�4EDQTD�UUTE�����"�j�*�"�
)��(�	")� �m�!LMM�TSDDQRQE1MEM[��TURS;8������d�4b*i��	
J(��&���J
� �!�`��"Z&(�Ѣ*hh&�J��i�&�T:*�f���"(����b
����Z���Ӣj�����ib("�h"����*X�(�**����b����$��Ѫ*�f(&�h�j$�*�**`��ӂb�*���h����
�����M�E^_n��{��]�mOp0Et�ˑu�k��蝾�y�2]��u���Q�N�Ƕ�ca>U+�Y��\��y��
nrˈB���v��]0G� P�D$�#2�@#U �P+J"L�(�@>�{�ǿ}]�w��{����a����ӓ�1������(�E�����*V�d-�����3]�Z�"��OQD��:3�h�4l�.�φ�82��w����\⡡O���s�l�h?8n��0�� ��g�`@a���I̿�g`�J\o���$�Ua�/'*[S�I@�Ġ�X�ьAv�\A-|��~����N��@����0\�-/M5��%�4;yԷ�=���F�_ϊ���:k��*D�[K��T4Ba����N-	���۫��s^2֛^SM͵�F������cZܙ�}5RD{T���X�@�=��w��<\"�j��e|�s�:^�w�Yx����x�Y�xy�=�ěl�)�A����Dp�c�������{&��nTl^e��}}Q��g�y�?�[Z�/ǩ��ZKl��C(�m�q,p�/�9���R�3�X��s�Tc�9Iſ�-���d�vUQ��ȷ���M����ќ���q���ө{��߆d(wՉz�:4sԜ�Hg)�FT��.9�EL���k��a�ٍ���g�3- q���Y�Z0{ݰ\u�-B�yP�ꃸ�[�=�8u9X:9�yhc��a�I�-'O��f������d�n�IN�@�H��V�h��;VQ/�L[3kL[R�^�+���*[^�)^�� ��^��~�b��hTb�JT`�
T��
DiA�% f(P���N�;��;�䃭kbH�h�ܦS�o��u7�"F����T�h{�Ȯv%);�K7B'n]����:��!�^֐`�5�,�M׊i���of�U勿bڈy���Ty��h+%�"��UvC�q���/u�84M��WXW�̦[�%T˜橶굕�(�̘5����̐�7�',�V��5�%w��	��ȨgM�p՝a;p�(t9�:aIT��Ī۰�uR֧��5�;���?=
sZD12jv���	��@M��<��H��b�����~�S*��7�q�t�9���~-˨�\[P"�l }��49�9����U�z��n�T��v ��7!��B�TS߃�%��R;��F71nv|}��A�-��+x^n\㖹�d�Y�����u��oB3u��NZח>6���ʏ.�b\��mL�^Mm~2���]0YuJ���|rl:�t%��5��M^�馯_q����,r�W��@&�Z��K�.����c��K!^=Ua	d�Rk�5�#�i�1��!��Q��_�=D�mr��E|����gl?���?0n�.���α+�:��T��.�י|���x֊�n��OP��q�W��K�y�I��h�{B���oqGĪ�i�
���wy��N,���:&Uh�0��=��>�ٽ	����C��D[S���dPe�ۜSb__-�p9�6����(o���ߝ���'Ȃ�JD(R%��I JEh �	��Z!T�)�i ""�]��h�E����Ko��X�A�*�@ǁ81�Ä�_^�3�u����V���UI?uz�i�<K��;z��k�!�]܈�ˈ~B�٪M^��N���m�(^� ��O��o*rEm�.�ƾ��f��MMww�6p���v�ǁ͉[�3�<��)�����83��x�26^��c����=)Uȓޡ����e%l�~P�d�R�3��������o�TX��>����u��I]z��K��^�c�b}��2|�#%�]*��M}nC?���:��V��@�)�F�Q\�j�4��a�˞ni�#��vis�0t5'�-�#�M��ֵ��cOM���6��q�i��Ek,6��2%�ˌ�iݮ��M� ȋ3]���S�{�������>�x8)��@�!�9�b[��j,O�����ɁL��E�,a9˘`~R��������L�t3���[�˔Y~8Q���i���re��{.�<`c������`a��(e��3���pΡ��%*M`�T[�����^�im�r!������{ _�͜E؇iy��6�}�sô� ��gh��慿\b��u�m�̋�c��c�z�o[7�&VBç�8@�PA��]$78��gie���q�t�z�U�*yF��N�W[�4�6w-�I��A�x���ɕ�L��Y�Q�_Ͼ���|>U)�j�i�h�@�R��J)�=x�s�o�;v������M#����{	�j�7(��Q�F,tzw�z�y��.ij�z���#�Lʣ�3U3�*^1=	y.M��<������v�;��u�ju���SÈ/|+��;��"���/�|ya|�/T�>خ�4.�TXm��:z�|� Eޔ�p��#����������Խe��GS�?����]�ő|�Z�`k�Oa��i��Koo�(�>�*O�/b��h�m��ߢ"��'���x�)xHܴS9�;�]��4.�ѱ-\3��5��`�����0��-��a�.M�1L,�<�����ީ�]�m��ОM�p�v���K�1[���ODܶ*�]�5Ȗ���#R��ǲ|�6��r��eo����B����-rg�e����#p�SuQDC],�Z3��g���ŞG�u��Uȩ����m��^k0���v́V'%sЗ�qm@]�y��֛�~ma�2���l2�p:��穭�$��yEn�h�>��JETE���*:�}s�V�Z��2�o7����=�Y��<`E�7_�ʘBi���w���|)�3��"�i�ʧ�m��U�ghB��pl��[�O��NZNqhAw��n?�u	�YӸm2��Ay��=��˗�:���U��T������z���R��Gi�U.�w�>W7�s�6�B���Q���ߟ~����v�|�JR�X���e�H%�@�F�h)��H'Ⱥ�g>}�K�_`S�%�T����d�S�;'��c��[��w�V�5x¸	[��p��l8�ر�te��)>�,�{`��qw�jH��e��cײ�3��[:�TU�I�<�f��9 0R�˪��B�����_p>\qP�}�/���dx�bԄ0y��Y��л]����͠�apͽ�T9鄝X�N%�����4�Xۓ9��%�Ų';+2�d�!�G�Z�a�tc�y�ay=��
Ԧ)�ΪS#��pf9��ˎʯL���5InZ�"]�(�	���t�3L5����0�>j��-ڞ���=s �J���a����r~�h�6!�����c9�%�Z�ʜ��O��Ұd�*���1�n�Z�1�n���ї�j�Oi��_������U"5tlh`� ���M��{^w�
_ ��	1m�"Xm��S�U��qjGj��j9�+�j[Z�8Ŵ�]�q����ށ*��<=�>?^������d8ic�\����nĽ�&1�ɞh��6!�F�gCk t燷�/��d��wIU��V���EK�C1a缱��u�;�I��3P��2�u��.0��/�@�=���ݻ������TU&X=��]
b���6k��o9��t�)�#��y[�٦`�)S��SM�m��sqwNo�N h9��j%��l_%�!�V��)�F�a�a����z�J�浹��|�"n���G��8<�'��r�� g�����01�J�Lݎ�]1=��VQ��WV%�<	޴�ٸK֘V�'g׭,���YխKHbx�G����$�����]�t�C�C-���E�Q5�觏�D��Ɲ&g�������n��:*xO*�ŕ7S�Z�PCm$�'+ګw�L�:4s��!^�Y������q��J�1��-���� �:����$%4W�HM���~Խ�B��b/��B���B�Z�]H�mE�7a�j�aN!6����>֐zMcX�Y?^)�9֤z���R�-]p�1y4M�٨H6���w�m;h�G#�Dƻk�=t�:$��q�L�UL��j�n�Z��Mo�a��x;�s���#��7z��mXv����ԝ`��w`x���=�?>��x�P���ܻț��;���l��(�����;-�"�>2�2h�/!����\3����-Q��W3�R�D����4ؾ8/7����~M�c�����kx��,�zS��#-��p�GW�XK���x��|g
�oQ�w8� ��m�Κ59тU_>�=���IS[y�re�r��鴪n^���0�[�͙E9ˋ7/%@m�R�X������z�/���������8�{���C3]e���wZo��qw�%t��^�]����Ǿ�;���r�����"@7��<�7�̝=��k����1U�n1Kz=�a�G�EW'�PK�ʤv�凌���8P+�C�"|G��}4�%�i��藵Q�Iΰ��1b��@���q����X3�R���b\���^3�����,ΎYk��ݭф�t i�*�yxЊ:���;����~�+-O��=�j��ql��ھot��㧸�N�> �F�lYj��yP���-G���e�g���h2��e<���sw�:�7)�MnN8��i�NJ��b,�� -0ա���jhgnU����ݸa�4뵌рV
'�VD�4D<a��d��P���7`�5$s�~L���Ř"�-R�
�v��f����w��ਖt�\t۱�3��$��$����5T�ǰ�6�B����o����*2v�)��0���n\�H)�h�U^�n��B�	�a�#U���9]Bz�-��WV�ũR,fy{+��ϼ��H���s+Q&�z�S�m������JS2zJ�5d�[����3�JbL�`ڜ���La�w�M��á��\Ԏ�JXSk�l ɪ�K&�K*�_����;a�3�Q�
���#\�$����C1����_ ;H\��MK5&k`S�,�0�˕����{�5e�+79�W�� <&B����c9�̫=��ً���S[�Zej��4�T��vr�dU䥙u�[�Puֱ�W����<��ff�y�}��\�	�V�>�D�{k���dz���wk�4{1<�C�=��sо�G���.���������e�k��SiQv��V���͇�T���T"<���,`��9�5��|k�V���j|�QN���..Q*�>�-?�_PYV�Z�79/Gc�t�9M��0��ť�n���O�u�;1UC;H+Uy45���)>�%@���Gc�B����+'�+-�ՠ_�!Ɗl��qom~س�
Xp������PE�$,���p5�#��Ev���;��7<��9�P�ۊ���ջT9W��|��M?F)��<�7)�9&,F'��yY�]�O0x�eV5Y�1��"�I3ؤ�4�a�vZ�Ji��\�ƅ�u)�Z�gN���.�κj��C�s_<bq=��h�>v�d	�j@���|�K����L�����bd��J7�nx3���d[Q���V�qT�i�!�b@��Vi d-�v=Gr��K��eb�M�j �5.64���v��EӾ L��\a��gE;��6D�ǐq�oRJ�d�,yn<M.�cq��u5B�e[�s�����K6;jS6qj �|l�ׂJݝj��bM�^��U��ٗ��	m
�*��2L7��J�8I/������goF;n^^������i��<伥�8Q�������b��ȡ��{����?��O� 
�<Rs������2��5`{#{����'��&3\�`���甅�ٴ�9SxMXK��	�����f��B��|�3��Hd�Gi�c�ǪPE���yha�B�;�a�1��O|h���7=
��N��
��`)^5V߂��R����ȏ],a�a��0�a �X�
��x"�c��h����yErh�y/J��v�ga4��7�Q�-��*P�����㞺��U�_�����2ἴ1�Kb������uӔ]���S�Z����0��SɆ�|�5Bjc���c
$�2N��t/mE'�Ķ�vyN�:�eK5:�G��CЂ�����)��VBj��b���J4�η5z:M��2�6�S���Z���n��ke����L.#�;�6YW��Sa
z����~���l�m���I�]�_�S�Rj�:j���m����=��ɚ��7S��pT�)PvGF�s�����_.�C������Jn/��J�Qx��O�N��ϐz�+��ɲ1�`�C<2�7�Ǝ|�O"�v2�<��>���e$[�m�5���<޽��q�s�"H��h녝�OV*��W��1{sT��C�PE��^�cs����1�n��Uv�U���o`��B�̟)O8	+�eu�w�"�P��L��Wm�0�=��HcY�u�bGw�ܴe���1��W�t���i�N�[�����'�J�zg�l�����c!�+8;�n-��� ٰ�g�=!A�u��W�@<��ٛ��[+�x��x��偻�K�1�0�r����^<�u���K�;�ļ�[ϣiG.���n�&�z�'U�¤�E��z�1�i��ޑ�P,,�7v�&k^s�4u�n�H:k�a>��P���5�j�6��ۧǰ��lC��,�x�,^k�ƕ�yO�0O0�{l��8����۶��k�����(��M@8z;��)��~q�h���r�W8V�%�l� �L�+'�W�֡9��og��:<�gE�eFL��ʭt�Q��H���A�{e�`�J/�]�ġr)hgdk�43�-F�c_V���i#�ڙ�E��6���E�h�r�i�9CUc�~U0�:a�y�[$�dC*[&�9��(���yl%��'wAM6O��ݶ7 �T܀J颌�Xv��t�eyJ(92$]�
Z�l�l�r�E�լ�¦{� ��My5�6���,�Xʭ�͛ol��ػ�ne�������~>߇������}��o���]�`9vjy��*����<�T���a��yx�c�@"݋a�):�v�fV~k��R�u�C�;����=Oyۀ�B�M����-1��Z��l3���z�ƨ��M���O�uK��i<��)^�N�h��ϹA�tD�G{^�4��LF;��}���.��6hdN�rȟ^�*Ţn����E��ȫ<�[�k�Ai��صEbKY���p#�9RjL�s�#xp.��w���I�]NՙVQ&b�H�,�����e՞`b�".l��aɼpMٜ;gD�;��c��RyE���AS0־���'M6�����bT��d����y+G:S��i۶	��t�>�u^����$�I$ p���2�N�ZP&����SV��Ce�sv�<�{���DvJ�q�/D��}]
����g�9���K�]�o�����m�ZjV�{� �7���I��]�bK����R��������D�x��p�շt��!���jf��ۋ�}�NS`�J X��-��MICdE+tXq�\�Zp�;q�a�RG���G��xu��:�n�6���B0�˳'%��bem�Ƒɭ���@3P<������]���w��������qZ�3y�+Y�X�\�6���u�G,�@��&�H�!J�ٹ��W]b�h����)��PjN��p�8#P�<���B��ݨ*W|6��W:|u	]G�˚� �S\5e[���E�ɷ/���c�3wTAM
��+$̽L-R;�vA��2x�K�iڟ1��ܹ����z�y��2�^��d�n��͓Fuj�.���B�b�bk��%��E��Xu��[��nt�z�<���z���౰�}:�n�Ma�RH��11#�e9��$��k��Dڝ
Pi�Q˸Y�y�[���G�o����ڸ�q3%��Q{Ǳm�-�*oN�Y�|k(ۛSD�uH�g�ٗb�'bK�/yjx2���d{�ʱ�3z�3�j���c-�kyB,�)]>�l;`�εao<68�
ɂ��[��sr�&�J�U+Nc#5�r�n����.��hĨ��oM��ɻ����X��Mb���{�>�:Yʆ�4�,f2$m[Ͷ�,�=�<�X#�nb�ZA6�!*�C�;v��XF��*�޺n��-"~��/-G�W6��jܷ�E�;��ECzT�.���q�-i��n�� ���:�if��u���m��J�,��v5ٝ������єN�%��{�&jX����I���	�o?$�5�ĎEN>����.3[D�훽�v��#v,͜l�;Ƨ;=y(�߶P�E��CL�k�&H�շ����4�c>�u�c;)*V�8����M�.-w)��r修9��g�s�Is���)�a��ohi4cc]��[5�9�؟��4m��ci^���/��6oJ����e���%T��;����5@��AG���Z��
��n���|ć]�U䜧#kE7��A�T�yک�������U5QQK@E4ADE5CM�PP�3M45E�@P13,CDE!K�����E�!DM5T�@�J&)��J�&���&���b�	����"�)����<�k��bH���6+Ri�DU%5EB�hĴ�2��S3AIAEASEUD�E%4�QAD�TL-�%m���)bh��6�DQPDED�4̔DQCMQAlb����4���QD�E!Ei4U6�h&�H��(����*%�%")SI��(h�"5��)�	BP�PRPR�Z4�P�)MR��"���?߿���W-��0�!�dwk4�r&���U��W-�&�z:�MJ���u{�c���|�]G���y��p�0S1p�.�0��v���ͳ����a�8cC��CM��(l���	/����K�=��>��0������ 6@�������寁7��{�g�8̦ՉU2�9�m�7�̕~Y�Tȴ��������������MY.EC���b��M9[��|������g��J詣�:�+[Q���X��葑��8�^EA�E���^[�E�xe��pM����h���c�B�al���T�{����ڣ����}�&����l������8�I��Нn��;G33�����)sB�CzD�w)e;Ϝcǖa��iv�1ؤ`�$���E�h��m�ls:��f�\`;��ߪe����Z��S,m@�QEG7-����Z��h�{h���_t���0I�[�<���r����D���������Z�3Q3:�q7[��sbj���T틭���q�mA�6����7��ip�kLz�qv��k���{u��	�03!�>��.����c2��͜���G��A.��u���F�<�kM�G]��#�И��OB�T䄦��4!�l�#5މ�+�f��1��"�*[�Z~����N��&،�3b�@��c.sOj�I穙�""v��df�z3���w�~�u�\
N�놝ճ�8�7J���KeW��)��!i��ԋ*-�ևQܽ4�/�mn�wK'R��=�NlwJTX�Ǵ��6Vb��iISnlR[�Y�]��ٌ�> �Ȩ����4w˕�i�G3u�^m�ZF���1S	������V���[��p]�z�tS���T�Ay��C���A.Y��ݰ���E�EH7X'ӌ6���u�<���'-.��J�0�lB��!�k��]�N����SQ�U�q6���7�Y<P�3q�(E5�A/j\���˞y�a�R�T��G1bߠ� �u2�������8CO'(��V6�I%�-oa�frơ}y��Kr�ֵ�FC�h�'&d��v�q�>�����ab}�́*�F���Wl̑�Ź�\b����yꌎ�(�M":a��Y�I���C��P��A��~'˿Oz�8��0�+P���{	E�'P���l5�s��v=���爲Tj.�Z�R�ҧ�àw��#3��cjM��O(㛁%a'��du �E���]Qi�k�;4U�:Z;�U�C�p������zv���Z��E�Q�F/�6��`v�.gj#t���e��T��ɕ��o�����|��,�yw��Ϡ�]����P�S�H��G���Q�*�KNg�����9��^�
�S�����~�6��4��8�+�+:�+/�
f$�.p�2̹��.� ��,P�J���z��yY(�w2�pw�mb�;�)�8B/4Pޚ���M�Q�䳵�of�I�	�n��ҟvj�2�JjJwr> q]v���*����~~bh�z����Z.|Dϼ�E9<���*w�z��*��ȧ���,����̮��B�2�`Zy���f��3m�@���E�vJ�G_
��ƀ�vy��_-q�}�Z �P��[����C��t�Ԍ�b-t��.�k٪�-0�C�)x�C���)�E;j��î����w��XOhǑ���������/����0�fˊ.��v��_��ΥO[~�O�A֧���̀�!|�t�~�|w�eR8}C�~��Dݵb{�e�P�и0���=�}K""I=Z�O�Y锿=�t�Fi����T�D5վ���Q� .��m.�uO��A�X0�����@Ψj�?�yƦ�����&f!EU1��+^,KQ�d��A�v{_1�q��y�ݜTw<�sT"��NK�v���z�E�QCj�I�վ�dY������!�!v:N�z����,�[|�XSP��H��e��cb�������<���i����*&)��_Z'�u:�7:e�i�>Y��Nc�^�[r�[)�zsؚ7��웜L�JHR�\l)L�S[�**-SwC��0كO����&�kי@%*J�&��)���¬]�ʔo{5I��.L��2�ָ�[9�j��Q�-��e�,,Cn�A�-�4�^A7.r�d��4�����-35u�p;��������,^�$*[��������u�o���-��ʷ��S���o6s�e���e��S�M�3F4:��nj�c�,���F_����@!���f��(��*��W�E�����}��a�����.[�����;��HH��}�<����橅���(�=�6�A����I�LS�a:y2�׉T��V��L��ѝ˨��X/�j��J�C��!�7�Aa���]����zZ#tM[�����˄;-W0��g��Z�;Š�0�A�
f��@"�e����L���=K���W՚��=�B�J���].�ڎoscZPXHZ�/�E�6�8�^g��r���G����Q��g#ǳ2'�K�|�;��W�� ����%�s<�U66���}�7W��oZ9_.���4BN�05�,&���b�Y��oX<g��3��1�*2�wgzH&n&��C��	�L� Y��d�޴ˑ��?����2Z��d�� _Ct����	��Uk�o�2�4ZK�r�g���
�d��8\P��)�k���̗g W���*&t�GM`>஻�RZDRt��{+�,��8�Q��z:#B�hL:n�굂�����Y`6�w@�Z���:����B�x9ݛ���;ONA�;���=׈U���Eay�oX�ޙ�Y�.���HP��\�7�M�*���W�2܏=<�wx�Ӈ?�Ir��X\{������!��<�1ѳġr ���@�����w�GC�9�3s����G���J�^��^�P�*�"D�z�(�9��6"F�Bm��2#�4�
��ty���.�q�N��}�PT�v�wU6��)��O�m��X�~ˁ:1eD?4��e�e�ѫY�J�i�-id�-�q<�tdn�x��6�ܥ���eֶ���U� 
;0�6��m�8��^����ډ
,:P��*���V�KEնl@������J#uU4l����4�_^�Ph��I��H�(bh-7.�S2硛6��ةC��zIt'�tn�u�Ȏ�x`�*�m�4�@����בO�S��KBO9!�p�-�2�[��w��I�4�D�xt��.)QN��6'��
���� �>1�Ӑ��Q'��̢�<_�C�)T��b�S�%��޹oP�v�Q*�;':{5�;ff�R0Ci�J���R#v�g��qZ��y��}C�W�'�@�H]�>�]�������6/i87��!���Pq�:��݋��Ʈ��Y���A�.]bzU��Z'%��|�V�K1�ka���TZ�B�ٷm�*���f�ëe,�8Jh�xv���[����ZqD���rp��	�֨�>�m,��u���af���ǓDe�tk-���{α��>����ެP�1������<�\|Y���Ňk{ȑ5��<7������9��WT5��'3)s��(��A�t���L`Z�0�F�F8�v#0�|qr�x�Gk���p�&%��N�i�w�<�l�p��l��:М���`T�^��!,5K�ײ�2H����$d&,�=���M홢�ڔ�A��+hrЃ��>�����ϴ+�vW[e"5�����W��ڇ-�l�h�����8�Z��z�A(?��8���8Y��7M;ܠ�������L3¡�4�������΂{z=�峜���h��s�,h���c���}s�noEl��&s�g���S@u+����]\M���5�2��M�L��j	d�&$�ÍS���r��ݙ��{;��"�m))G%Y�����jzM]�6iLԎ�P�ZǻaM��bl�k-����m��:E���;�&Z��K��ȗ.�	>'�p����+�M2=�I��� ���w(�j�G�L⭻��|��sط0�h���}$���C��d��:��]8z���|���okB�ƔQ�2rSe�&O���P�X�u��_a9b:;���J�R����]v� 렖��z�S"xu��0�]4��hє��뒴�	�����'�vn��n5]�:}�zڣR4uw41��t����^J}��
�@L/aho�H{���ϔq���À.�}Ae[j&�1��{*�<c�'U��5����}Ͷ�"]����O��=���=�Qk1E'�Ĩ�im�,�l�1�ges�bdf�i[��T�2ZZ��.��h(p\�r�Y����]`e�c�G6�7d������zc`�h�Md���kzݵ�P\s^��[�r9@��+�R��䴧u6�j�X�Kɾ��Ɗ�����b��]�vBrf)`�3Y6�i��)�f����e�Ƽ��r�&���"�,ܬ��$�Q��l��t�����n�`�&A�{�8�P������"�v(�/>�%v��f��BytTv��2��2���zF��c5S�4� Rf��ݳ6�u������~򭔇��ػb���mމ�a�fl��&�<��l��UY�i�����O�[�#�2���K�ñ��W\�����9�NW��&I�T1^+%2�ơ �6ge�]��rOYrn��$V�W��t`h�uCh�Sbj�xB��h-ˀ��˝���=���a�}�!��6�5b���x�-ynx��B��'�����to�dut�wC 0�
n��׻�>�p��Z�v-E�Jh������+��)�v�Q�Dԫ깧��3�x�c�B���jM��Lw�#�^):�������׽Զ~�~��t�,�w�|w���4�,^� �T�U!�U��"�^[=|_�z~͌.��W��g,ap���*�A&�9�������������]>��#��;������;��i��`��'��� ��(�}���y�a�WJH�d"; w���=O��
}˶��t�s�+]�����ژcC�cPބ˞�(��x��킫tT��Y�S��hu���(�^�O!�=�r�9�b��:��E��cD����q)��c�c6s�,�Q-P�`���9tjTJ"5��q�Z �՜��s�;����f��*��IՆQLy�C96v�y+��\������puN>8x�Y�7��~�_�^�V)�3΁��~��Aݤ���I�VĬ`#hn��o������-���"_�b���C D�=Q��yP�#]��m.����}f��T�q!]���FK%�����.�eq�ص�C	g秨F�q��}��E�L��+���;��~U�
���T�Ű���n��FK	�.@}za�?H�`���0`WR6QT*(����K
�b嫍M��� 4�8����y0_k���A#�.�e�.���eg/�B6�鴉�{��;�/Ne�}�M�dE{��L�/L�d3+0G(*��9�l�"��ݝH���3"�wy�{Cp'X0."m�r�]�����c$�X^��X@�~�Z�F�v��P6zz�z�:�n%�+֣��U6�q�h)z���*Un���K>ߪ����S๙���LpUG�^���z��XX&5����z-�d��3��N�[ưLv�,�\V; t�Yru���[ߟԋXD�������6=�p��U���U��A3HV�����̖�7,�፝�d�hV�~Vͥ���x͑�"�z獱�$-�������%��n�rN:�6�"�Jm�`-�<��몎�g�兀�T��d�t�umR�c��ձ�@�7H�T��/a1��T �C��9�m�X|��th�'tW�ό����ճ͗�=l`��V�L3���6+����8�MjBmJ�M��hز�߉����~�u-{�^��y~�2��֫O<�mA�S=�RD���
��u)d��%���V7�U��I羧�g�U9cku����..�h��Q�
ds���l��z8�
fb����z����N=��J�<���n�WE�x�̘h��Q����\��t�;	j:sr���#�����n�}�V�Zb�{��!���z�W�M�.��z�KZ��J��oݼO^�9L�a�F d�V��7t��(��3	���2�T譐N�e7��N�@�ҙtF�{���W��d����:ʐ�Dn��4n��Zz��52��w�/rmbn���O�����_����TKo+������d�aFX-ف�莚�ǟ���Yt§]��H��;-(��L9qF)W�uG��Co?Q�/Ɏ�v8�.<
�ʖ������!�D��dc�rsC��2s����{��zD���A.�;7b��4�'(��,H�r��Exk ��z�j^	[{*e�@�%���5+�-E��Gr��j�- ���j�]U0&���o�π�	ޟ��C��L�_(t�ޔ@����o��^�5�W>�D>�z��{�?N�P���tj0i4��F{(��w�x�;��s*F���lZ�W�s��̵�zvݍ��ǟٱ��D��:H�yhgdn�2n5���`Ǹ��u�V�����ߗ��^/���Ǜ�%��0h����W��YkdNG��xrЇ=�Yl���q�~���3o�Ŋ����7`9���QO��}g��k������,a�����I��z���j�VQ�o/<�����c'��T�E�k���Ϭ.3���1>�x���}~�//w�����{���w���XS�����W�f��+�d�N�$,Т5��k�F����+,:YVI��6�M�⬝�Qֶ+�ydL�č`G;8��Ǧ_e����QU��T	�uXKg����g&)@�RZ�0v_q�۩��w@�m��l�����H�ob[v_s�>�;>:kV��Y{{g$K.��q�<��v
X�UN�Qǡ�8�H�Qb�a�o6�b�����+h�ԇ�g�xh��ݮ�Jw�*�pظSB�a귰-k#�]��3-�A0#qc�z����k�X�h�]Z�e�gxIq�+���U�o&���B�o|��<	cq�L+76��#���+bYV�HG�����A�T�(y׸:��=0Z�ە�9�c�6ঝ�Pb�X����ż/3��Jٖ�Q?��k8Zs�*6�*���4�@��謫�4���b.o*�D)O�F˫��^�J'�vKՎa�Z�t�K�xŔ:�[�tL���-`�ΰ�y��u���q=�VQd�ֵDE/pJ��ԖCso'un}��֟>!�LX���]Y���GUA)�j�'�[�Y���.�XX��r�P�������ۮcOj&��
�:مC�6��m�8�o�6%\��=
��7ܖ�
� �v�C����]��v� �������Ks�b$��E�-@e������/�8S͸��?:�6�镵�VAL}�u�����r��r�z�p����mc�r���mu��P��1��������z��0H��o���
`�&�Pi�����Սu�2���à���;J�E�X���T�3x�ǯDL�RY�4��!�]�ι���ׄ�U,�V�6LF���zI���)�� [y�]I���=_i֗3�U��b����ظ�.��{�h!t"��*�mo}k�aM!
60M;�KL�Ā�4X�b��t��w]����T������[݁���\%-Cᴨ�mkMc�t�9-����]�xuйzn��Ua7� e���A'���\�!��~1Y���Ww�
9���@p`���TrڡoEc^�!vz�&ӒD��o�Y�0�ձ,�g�^P��ּ��̫�HŶ(�ȑ�2�w�Fs����Y`�삻1�QT6��te���z34�7J�\ى�#B��K�
��*v����{��d�9���.���,u�9<�y�:bY�]���\$���1t)�;wZ^��� �,�qφ!����y�6�.9sj���\�_vG��:� �n*Y��	�����V:��Y�9���Hk���6��X�`�Y@P���fV��[ݼ������i�s�k/�cy�򇴛�K)�E-��}��s�R+�ĝ�l�2�U8rwKJ�ʜ��#"��������c�)�
<�'-�	#i��6�b��{ÔRj��#��<�i
�()��(
��)Z)JF��"�*%i����J��ݦ���F�������6ȕE 4�PP-%5AE%P4�DM4'Q�J���h�����"��(���i(X!"d1��)����*�(�h��"J�iJc%-QIDPQ!C���D�U@�EM�T�%44�P%SKK�h�R��T�Q�IQSHSHD%#@�R�AK@R4��r�H�д����������rB��V7�,�ok
}�N����V��ՖX9����r����`����X=�}��玒��3�M��w���H�K�lv����f��o.��xX�8�O�Ʒ1*�Aw�}�w���i�1+�cY�/}��)��Y5 �:�\#�;g���HP�՚�ea�.*i�ns-�\���U��KW�R�f��j���wk��&�� ��n7R˾���mw�
�%�'��#�Ms����5M��#4H蠽�`�_k�p[����ō�&�K'mW2�����(���(�������/�,�a�[�QpeZ�=J�Xݐ*y��6���a�@^�Z����S]d C�Wt�c�L�E'��m*�z���p��yS�';C/&����C��4���G���u���8;5�!�:`O�i��w��G7v*@�3Z�[��%>��kXNX7��H�zB>����S�޺�j���s+_\���m�Kg>�Պ~���C��Z6�ͩ����rj-Q$Y6���ιf�r�x�S��+�)�%�+�}]�e!H�E��)�t�kg�t	�棰����Yf�T��l�ڇ��޷���a�y�n�3p�Y��!��HX*n���׬�ڈm�z��fI,3ڶ���A9T�|�U�I�ӯuϪ`��ҷ�F��-�8䊉8���Ӈ4����!���>��L`�nP���˂�WG����'��{NW��]ᱺ�s��ٸA=s�i��\Χ�$hcU���@�ֵ1������
�|�6ۣ�MM�ͪ�2�	$s�ƀ�h���V9��ͱ����Ls�fl��&����w'g��Ǳ�ܰT��)��Ԃb���F�S�C]��=vz��O<��G����^Z��}or/�	�g�sR���C�e�s���@v�.�X����hn��A���P�c��tɲK��OT��f��f�zG�ڷ���!a�T�*�q�sE5���C`�h_E�{�g~u�w-a����������k�P�&�ג����	N�jRf�`-��Z"�H�͋a�x�X«��о�C�yO�\��΋���/�Gcq[�:��Q�bM��⏻Ǔ�֮�ӫ�?
kЙs�p%>w�e�%_s��`��*7u�d�1�5q=�z�B�NsAg�Z����Y�����r���D�+��Sђb�[���m�f�4F��kb�ص!F+c;�b���� �,vzC4�)E��&Ru> �:_��aU�E�'��c�/n]q|��>0�J�r��37�7��۔\-,���G�t��J�u�������CI��]Eo��6 ��[*A��M�Q�՚��l�	�qL�C�%Ь&�*�Dq���J�v���{���[�@]��maɄe�����2���z=��[r�,�1,g,�1��ܨE�{�S�n��\j���YU-j@�g�/�S��M�~���.�ֹ`D�/FJT2<�p�	��z��h�&[Z&����\,�:ӯ"�b�.R�`WG7^y��+a�Z�����@�`�[�i)ƛ�.*���LwVSo[2�{h������yP�4*�ҭS������j;�e�%��ӭE�6����k������h_n藹�`��X�ô��z0�̼��t��uX�(��s��כw����䵯��"`��}e���Aށ0u| u�Dai��x6=�=7�4�U�h�Z$�qC*5�j���=)�ШӺ���RΆ�b`/��GS�@��3ʄD���\.�o�I�9E����y���j�K> 9D��{	�32����;��Ϯt�h�+ҧ�Y%;"�o����y6�׽�5'�	(�8ab�܆�"T��П9ѳġs�KCng�Cb����|�Ɍ���M�
n��ҡ�V�(]f=���ǳ���=}Kl��9B��눯u�!�ߧ�#�IV,�U��W�y~�l.��%�/�f�藶��9�xX3��ڙ��B���`�9tM\;���.c�<���Y7ɘۋ�����`ӧ|7�h�:�M��+�'=\�ʝ4�W.h�8�t��/�:xup�0�edxY_����t�Q|)5b��9�X���MϜ�u�]�V�Z�xԏY�d?��!y���"� �1�SO�|Z;����ܡ��Z�e�c4V'"���W�[��_��~�o��Ÿ���sh���3��M�-�7�d�P��6�t�^F��T�6б�i�nӕ��3��C>�t�D�+bh^�"�nfF���
���)�����!V� �b�f���	*���M6�Σ�rT�E��X.�H��=G�u����}�5�	���<�EŘ�E>y�V�|�do?Q�/ɵ0��O,�0�$Yp�f�8g^�"#5&���c#�T7����J�O`:�]��9�mͥ�҃8�a��T���	�� ��b��S 6H��[Je��]Ew,\������m��@��)Z<�4��G�@��&4tyw��/�DE��ņȑ9�������x/�n������B=�)���`�I�&9���[.��i��i�{�\�8�|�HV=�Xb��{��>��
�"��Ց/�"䭊��v�1*n���Ѧ���[$����I�����'����[=e5��%�nf�F\ل[W-��~3��"�{bS��7/�[ی>0���t6��89�	е*�x��ecobi��-�=gM)�=�<��p��f�x��˄pkgo�k��hb.�6��}���Y��ZX���~��y}_��v�Ӯ�,O�*�cٹm��EjR��HQU=�o�8�|���%�Ac�b�Cp����@^��Q'��:��m�0ISi�׌�Bu3�Y6KN��ׯkw$x�g�f��ϵCBSE��P1���6n�T6i2�
�W)fϋ�b0�e-9[�m��g�e��{4�Oq�o#�3��M ��6��1)�w���S^�|e�ã�"�=Q&箭��OEe>�����vz�l�R!���91�}���^��au���2��{,�a0�򙘬ٴ�1��v���~a�}��.�o��&Y���A�%�b"]�˵g��A"Z��ի�Ǟ-Z}�j�a��W{uƹx4�7���|����R)��S��Td>6��vT�sz�,Xz����Ҟ)s���]�lۆ9�y�T�q�*V�OI�P��,�aעrn^D��A�k�T<��X�R+|�����C���7B㙣s��{���b*J{�	P%�ޟVӮ�"<r���DC�Z`C���+��8L�����Y�ۢ��v��Ĭ��L�.�a���,�7n�.�fDv�=峰|����'h`�ӧ7gM�-��YŎR�%�[:��sb-�C���ݍT���H��l��:;]�S��YvS��)8ŕ���N}fWRAp���d��\��V� -��`��K��?2i��zv���Z�7(�{�elx���gsrb�������Γmr��09���@:����^S�<�̠KVZg_��Z��#�[��k�ۗ��{�h��O���TI�J�8,�����[�tⴥr܉���v])ܡv�i�f�6��Z�����O������o.���=s2_Q/L�.,�cI|�8؋&u8��F�5Z����^��r�4��8��L�;�j��F���H��!������Oh�RvSߪ�'\�)��3�%~������r��g�PU��B��b�D�d+S�0�(	�7s��d�iRͩO�<|���Aݙ��Jϵ���4z���.vW,�o킒� �}0��Ƙ{.���|�o\�-�Y��M�]�t�,ǳ��z`���(�����_����-�"�B����r����;�S�拼wG��0�a��0v��Q|�Iv�yE	�E�^��;>]i��Jb}*y4\�ʞ��2l��C&>�.���S��/�~��z�ө���=�E� �9D\�d����Uʣ�e�^���i?Lyb�Z+�2��Ѭ�]%	����%r5t��O Ü��>��nSL�@�v�o��`r�^YAv8Î��d0�M��Y�9Po71L%#'^��2������K/bɈy��D�]��6�8p�4rm�v˰.�=G��c�ػK��X�X��	o@�L�9�Q�囮���Y�/l)	ʘ����0�;Z�bDu����f�Pv����Q�D2�4Z���R/�T���{���B����e�Z$v4�á���	�Ƕ�q��p�|z�!�d;�n��Y�s����>q�����~��,�3o?����R�,��N�
�	�,��`k�!q}r��jX3�k��u䋤7H'��3���LS��,��c��6-q"pD��A42��ᛑ'�~�#5�a��i��ƛs�%�uȪ�4e��S�8JF�wYX7R0A�%�x[[KfDʚ�f�������ң��n�r�0���b��K��b�t�-Gs�����K�9�z���j�^GS�d�����KCp4�U�;�ӳ
e�F�^�d5Ϸ�L��X%l�ϓ�Vi�n��]A�z�PVp�֝��s]��R����}W4ɍ�\�`�k��{ T����݅�����຅�0�c��U��9�S��"�c���d�ƚ7x%�,=s�<:>���hL�z�z�I m-$���M߼�#�I����)Y�B�V�֬����#m>�;}�j\�$p�+(n%�����~�.�$$����wo��|Ep�t]�!��A��wMu���:�)+sgw��/l����=���,�",�����Ly��if���呲e��(�����6�KB�CT���q�Yg%�f�jMv��C5�����z�
�d��Z[/�%>��;���׼B�z`�>�Ϊ��f�Y����w�����d�K/�@tkW�2�P��a�78�?H��|:���_��n�f��E��t��۶������*eC��+~�G'���o�ٸ�~Z�[�";�����*6?�P�q�n��U7�D���&�J�V9��-�0��n��ib<���H�&��2$?��<�dd/�M��oч�
��r�CB �#�ٕ��&�Y��#՛3h�넋�gʑ�2�ݗb`HvGp����GS�����T�T[��5]܇u�	�-�L�m��y=QA��˦�'�Y4��&\���q����K�Hn�K��S��fD�޵`��,(%R[�Um��u����O�R�3��iA܋]w����|/�h�N��A�j�	��Pz�E���������t�'Z�)���cu
��ۢ��Ns���6��Z�U\˹):�g���=B\��7�Wj5���q�+��G���1Z;3KQ�;֨�	go ńc�ӻ�Z���Z�O��ͥ�NǔŁƻ���7N�'c���AM�\�`˧&���:�����{�����$�؇�,�5'������Kȉ����	tqD��c�9�S�ڋ�;:C�Iᩩ�����r�3��\/&Ż[�N��;�pj<��0l�؆&5��e��u��\�`}�.���+��A@w0����/WŖt�x�9zF4���k��N ��{;�p3��2"�v�r6<ڃ�XLs_<0��PkLnp��؜<�M*ym��@��U���Uў�d���kZ��c�p��]����W�x���4m����4��i�����/��c�:���05���.�8�fh��5��;CMJD*g���0��im�[�o����� �z��Z��TQ�c.X��d�Jnm�ZF	Ud�{�[2����Zs'����ͅɰ�ӂ��4�a�.�J�Ե?��_�w�{2�Q����l���uUN��M�P����d���ނ�̱�����"
�ٍ]�5����d�`�Gv8���J�g>�g:���b�~�+�x?���h�
��4�]�~���}�HT?�D_���]s�����s�Y���gm��w'1�c�/���k��z[�-�� �لd2�eJ�{
��Fɩ����m��}�T�K�qT)vf�K���r��#�o���|O��j����t�4e�R��'Gm�ot!�0X+Y�s���k����爝�����Ё@#���d#��Ƌ�����"+��BC�DȖ�MK+U����a�����:r�uz:$���RuσyM�:�4"��	�hǪу�r�5�֚+n&�sC�a�E#����8²��4��--���Z��N'+@���c,xFQ�p�n�Z��Mnz-L���t�?&�XM�q���&�����=�7f��j�a���UvU�%�2o"Лtwmrr����gP?I�z�Z������ ��#s�KF�)ت<�V�d#1�zXNp���S��s��n:l$�a�9�pj^;��/)�߫hW<�A\9��+w�3�ޙ~�ul̅2�T��eAlOa"�:��_PNME�$�vJ�&<�3�Y�.�j��}�Z�3��.�/����>m�J��lb�gOkc�ZL�5��O�P�w/̵g�+���?�X塂�1�l�y�jq�]C�@|33�Ì`h/�6�dOP"��Ydou��:���3/�HCׁ�h�?��U��gv�Yx�w�%��>������x�}��o��������ww�}o��V��ڞ��U����9k���
�$M�G(�iZ�e����H;i�Dѭ�ץb�N%�q-Z�U���({#2��,>$�b�S'�pd���.���/#U�hq��۪�m�/�����2C�f�0uˇe,�g=9oJǵ��I�AE��"ڸ����z���ˀ��=2^rӂ�tiVӥ��>��X[���o����V���F�ʮ�A��nAG�J�Z�Ճ���i�sa�r��4a˒��7�p���ەw��,�͐�Ge��w�Vq�Nv#i�Hn��mO]cL�����ɽ7z�WQ�37!�J2��8��}�m�����k8�kd���R�:;Ul^P�O<B뙷r�)��5��d���p�w�kZ+�.�1�䰁�Ncw�we2_)�ȭI��6����q�(��ɤ
�˔�Fӫ��>3�e��h��E"\�+l�S�ƕ��Iwi��V����g�ʼ!��Y��쎠Ԯ�a��1��䱪�&SO��;�U�E��#a㦲��R޷t�y$�{�M}��c��#��0���s�j��=�X�=ۄQ����jO�`��,�d�p+���V�"��S�}Z����5����g1�נ)Q��w��J���5�i��Ҭ7�O�«Z�|�W�.���Jg. ��o�Rsӕ���E
u��!9خ����aV��B76ž,R�Y�I��'����U�AG��:L�j]�]�O��/t��6��ʾz��K���ע�N���13"���\#����TM�vOFܹ�'������Xx#�����9��
��<��J0�X�-`Ўrb	V�t�޶�i��U��.����mTuf�.*����r^�k��u}�5*T@w-�#=�s�gr
z�&�\���&�%�E,�Iq[|ҕ�܃��gZR���΋��j�W^�=R6d1r8'��^u����i�{��n���gEеc���|r�Ѩ�(�1R�kT(Ex�7�Ma�Z�P�.N�KZ�:�_��m���:��f�Ix4�+���T�ZA�:��^�DK:�x�%}N��隖b�Mf�t
nY�� �)0N��8M:�۽&�V�dOgwV�3��O��%�n��Cd��k�*���i��"�L�z�=�̝�fܸ�����oi!m��n��v��oH]�Nkd����:+7�"����Y,'��uՙ[�Gǵ�QP�q�q�o��*����e�L��/�3}0|�V�b;�0�Tr�J`<!����C�&��O�+�û|з:���U���ͻy|�K�,+T��lx��`ű۝�������tNU>W����dM����Z�����|�Ҙ�[k�����{p͇[��-��mb�1�i���s.���w�mt�{4_]p�z���[��y�v�,ʰW+ k+�/�w�[J'It���^��r� A]l�]����i��kk���6e�Q>�WJ���!&�*�>����

�
"iB��!��(�b��JR��h
@���i ��(h���hZR��hi�"U����)
B�JP�(Z �
O��Zh)iR��
R����J(�(h��B���b����V��J�JT���%b)R�((F����{@�(b
Z%��Z�
"�)h�(*��()j�P���S5Fˈ6[6�<{���қ�*6����{$�)��WY�s�o�%���ia��N�j���ЇqVr���;I!��H�I���a�Uz��\���[1G��_V���,�5�&�=�Y^:��fpϝ���pE����͋'#���M��׌���3�~m\�O6˔t�[6_@� ���+��L�Eje/�a��Ԍ�>�>|>����
z�&f��e�.��6'b_5�.�Y�v�@?��.��(�6/�轙fE���p�#-�7,]�:�̌�Å�>"ػ�K nNeuܽ��AP�(�vqQ|�I|�P|�h�%�h���6j��"����q��@b9��+�MS��zj�XÓ�?�A�=^�����N�⫺�ܝ�#��S�-����R�N�<�V9��>s�Ɉռ]�j�K"�[V�&I�R}��B�[wGYpgc.��_NZ��ng�Dv1�齐�!��[�������J�cD�\�8��d�^m��V9��^�Ū��׬�P��;{N���@g��E�~� �,vzPط�jkc*����"��<B����(d�u��w?�;f�^��a�Rc�*p�(k�=��^��S;�j�����a֍�<^��e��0������n�n���-���mJ.�����{�=�������b�ŏ���Os�����"��fv���&�}��� n��Y�
;�Iػh��d��M��:�괖7{�ŃPZ�פX����n��<v8�uN`�% �J�����%yV��]��|��e�6�����=w�9p�2�dV-��7O U�㝼�gV��7�����r[w�B�τ��E�S͔�+�ɗ㖫�ZFK$^��pN�ϭ#�]�F4jo���)�bg	���p�b�y-t�3
��G�=���,�*\a�����?s�����*!S��c�nr-<��;x팲3���7���\v*}�Ӫ��R_ �rf��\V�B�z���$�'��w9��P\c�C�o��9���Z�Θ؜�x62:0/Xq[�k�?w�D��&zՐ�n>5:�\ѯBM>���gCa�0������2�5��a(��F�B�wf�5���'n;Ӭ�@���,��}#��]&�7,��*Ə2~��3mT���S���$>�����{h�3�=�"�*�r��q8A�!��
��>�6О�a��TuO^_� ׫�
ۦCt��J�:7ؚ<�M�wM��f����g���%�9آ�Ѱ�wwV�f�1�5"DW❁�2!?�������9��O=~ECÑ��j86�l��7���1z����l���	�`��Р�w�Dy4�e�[�>-�
m���~kL�SP����dOcP�Qy�s�|���/�=�0\�Z�<T�d��o3p��l�	�oCs\�8у>��r�@�!�3;\
V�pt,�/�õ�nM��>�&e]��o��%Y�C��X�l��tYx�9	k�G��u��G�������w����Mx���C��wMUv���ʢ{17eؘ��0�Sk���P���ƛbʬ=WD�3/k���aj!2�	U2Nw��OTPh�o*�Mi�zTAz�\��t��*��7L+�/��[uJ�.���]���4�و���*��؊�cyϸvYԍF�1m�j��s���	��Wsy���9�����mj�&���ݺb��E��\_�'ֿ.�n*?5�а0鸮��k����؁Y�
��6�����������g���T*�=��_RP�C׺-ޒ;6հ�M<�R4G��!y���Y[��\���߆mL��V����β*T�9P�vY���2�A�
��ld(2�ֹs���'x���]�(~}�B)���:uٱ������q�l�z�w�LI���7�A�i���݈�����`�d��9��Ů�n"��g��UB�ڕ�Q�(8p�5���yS��7`���^&}��VL�z��,۲������������t:�۫��:�B�,B�
o P��ײ��ڵrl�Ӯ�,e��'=��l��x�ĥ�i��_V�a�N&;eյR�/�Z�y��lFc=թ����ʛ�oLr�tS<,��9���u�!l���Ŵg��d�F3(�2]�S~o��*�)�1����3j湖Tm�����R��wZ�{e�(�x'Q<��m��<_5�S�e?�	��w)�����{%�芟�(B�ϋ��l?g-[�>[d/o��~�<���^���!o��cч�ނ�uicJI����J�t�/�x�<*J��&%�Ef�)ݸen������g>�����	}޷�}�Y�WVu�&RK.�L</dIP�mĉ&�c������0��EI�y��<
M}pC=r���gLy��y��T�j��ӎ�.�dKWe�h:ꁒN�}d1�ű�lЖֵ�gL��Zy'� ��d�B�N�5]��kY:����tyb}�-x��a�QI���h[u��z�
�n�5to:ݑ��?UP׈˕B}�!�G��RM}2�Ց��s~R��%R���Z~+�V�Oѯ�KP���U�����^�s��6l�����#?@>F��)�.�qv�ܕ.�/P��g��5ϋ�F��R�|Ū�/V���W"@���י��(k�(pv���:f����h9�����E�Q�F/�5��^�a�;� Ϭ1�������G����������:�gUEG;I���ڃ/�+4F��W;QǝwYVP]0��pr��ӌ�
ywۆ�ctn=o+�i����U��Z�2+�Y�C�㾬����Qmb���޽薋�y׆�h��$*y�uty�C)���U"Z�nW��c�D�J���a>�����j�g��|��[�)�݊T��������=zW�PNMG�
 [���8��as�ЪE^�@��<󗒋�='��"�ĪL7s:skg�t	�捴h^��Y�Z2�;[�&S�v��� w�R�ZH�¼�S�yOYپ.gS���������m)x�o^2 Dק��U��=,��XLgȶK:.�/�ր��g�kUb��W���M��W�s�;(c��;�� ��R,1��B�؏ʀ�ߊQ�q�L��ӁC^�\{��7��u�"�Z��Y�MX3D�s�Lz_�Rl.K�/ɉ�,�9>�Dq���ɝ����mEOoi� N��k�t���3q��,^��oT_y����|��{"u
��Qӫ�`�i�$���e��u/X�ڻd��Q0�/c�(zB���l�7�]�B��Fl�:����9�wɾL���"l���L��TRj�]��a(c��J����^K(Q�8�[m�����C���1��w O$y�p�
prO��rb��4le2��$O��-\�������N�%�IjZ�// d�(]K2��h8H�, ;Z�Y�����J͇���O
jSw���71�ޙ"������;t���=\�A�	���rdф���	��v)��5G�F�Z�|e��+2
|�4����b��o ����7_�3�+��vW�Y����*�L����H���#ɯd=7�-SK@�V5���C7�%=n��S�c��"Y|@r�oج^�Y�6��ke�]�4���K���'� Ǜ6���s*u�o�}�.�f\T���):�QC��y�����-kT˪�$B|��������������C8���L'��b���%��M���&Z���!���hue*f��@��>U�}��TCR�	�X�Ǝ|��&�}�L� �\��FK%�'�H[L�� �0�r�&��E\ў��)��<KH'B�~r�q��GggJ�N;7��׭Gs�=v�mJ�3���h�buİP���:p��S[&塀Y�#�u�Yw�s����"��\l��E����H���+�� %/�@�־Q��L0+��S]�_�F��G��.��&<��U����\U�֧KCw*��\^����C΄g���P������/��R�I�2�*�U
�7��C!�cc_��H�an�r=�4�9��
ވ�;.	��c�(�z���~���!>��^$�/K˫�󾈌��OR���f�T�$��T�#?_Y<Z��W�e���`�ڲ��0�5ArS�._�v���Jslh��⫮��˾O6ƭ��GN��vݟ���Y����\GS�҉�ӭ��VJ�i�fe	��q���>9T�6��߄�;7�"r>�]��U"'�k4�2ul��d����!���F�w�B���N�\��gy'="���Jw�w�@7v��B�����?X����y�ꝲۖ<�b��I�X���i�D+���Sj�hP�(74�f��R�mk�q�+�U"\�m��ϻ:��^�'/��0U�Sjr��"D��N�0���oQ^�oo:T.uU[�-��`�q�JX��SL��VG��z*Ze���"�h��eQ/�E]�s�t'�牦�U�#�q��)P�K
f%1�*��9�j�n�k+QQ������PM�N?v�I+_�nM[\��#~�Y��~�����������N_�e����и�"A��/�.�	5}�qT�A��Z���9���Jn+K�ΓH��b���(����nD��kR�R��8L��zd��ls�iE�&�`}��.6g.��lW<�Nn�e��zg3�Pۅ��wu�n�����.��b�Z�/$��0@��=O�IO����m~���H�[ ��j�WB/�Z�^�3�
J�g_7���"b�Z�D�T�.q������(�{�Kݢ4� ٠.�޽H#F�p3[�]�i��A����9X�#���݂�'Oy���0T������Sk��kNI6U�ۖ3�qYu%Y�t*��1�G�^���4�9�~P�b�����Ib�4C���4r�k��cAk������Ee�)�Q���qϳ{����,�������.�`1���%�]�Fn`I^�x��-w�R{��js���Y��aU��ܨ�{k���ݍg�4��M�2{ME��%�&�g�1�f�ݗ���\���#P����K{`_G�e��{}^��h���[�9�#�S�zF�����y�f`�T0a�ٍ�hrw�9]&�� Sڧ�uP�#\ӱ�օs��*q8S2��O;3�5T��:!��DS���*�eC�	����Yȣ�$qe����S����b��_)&�œ=B;���i|��U����O�L�X��I������~��~{�Ul*]w]u��t�v_+(N(˚���P*����ɠ
̪�߽6��i��7+Q��|{5��j1�C�x�\�Z[���gJ[xd�*��Y�zz,�d��뮷2L����{��������l�Hh��1m*���
��l���p�φ�0�z��=�h6f�˕�g�S�m1�	�p	@U��6h7�U�l���e���n�P+�ӌs4\ʙ��VY(�ƪt:س�)Ϗ��=�^Mb=O<�;05_�꯫��ó�'����E��'O�2]|���}{]oG��n����Ԟ�0�P*�v�w3dѸ���ݻ�F�̞��I#Ox�Pl�*��\Z��BWq�~����H/�yf=����7��Y�8�n���]yFN(��e�fz<7�}�҄�%��M�]��g�Wt��ܹ��ݐQ�����rYi�ݮNS�p��eʨJ�a9*w������91 �u �՗ТЖɽ�;���a�Ӯ�^"ok���gHEY��LGX��U�ȫ��ɟ���c������^�b��A�C!���:W���e��~^śt�ܲy]z�k岒b��r�������u;��a�7̳�����L@Vf��t�7�Pi���gp���ܗ�ͬ|2um6KHs�����5���m��EM��Q����*^�:r�Sf���n���>%�w*{�+u=�_e����y��s���#����%$���u�Z�q.
�Qw�ݲV<��(C���aY��}ŕ_����܀?(-�j��S�S$��_\�����Kgv��c2�9�x���NEJQfM�vD�*���+rV��8���;z ���U�A��{�5�ۜr9��˹@��32^F�&��Z�)f^���mR��ŵqee��+v}��3-�WWjb��Vp/ r#$�>�����;���]�ؗ�����ٽ�j�c^��ӯ�R1UϤ�T�7�����7�vvoY�����ț�� R���w���s�߷|�fC�j�e[�6��3�R�玴!�J���O��u��fn�Ş��ی�U�)wm�}��/E�9��=z0_`V������D��ܸ:R+zv��9�7�h]aL�������?���%+�9�'�~
�:�M^\�z|b6�f���#�^�p��.]���=�yʽ�U5r0Sr��,��(֝�w��4��RV��o#��s�G3��	��{*E�n�#2��ӝ�K�oz[mT�f���-�(�s�W�l���3�Z�#)Z� ���0ë�yp��"0{;8��eZ�$��O�����=�>�w����y{���0~؇�9Dk��z���v����V�t↗v+������!��Y�o3�\')�L�ݮ�7O� '�N���������,���򤼷JW L�:lKy�]QV�#D(9�����Az_T��Ù��-7{3���9��{�F˵6TշXK��@�9K�^s���A���vwga�0`!�]��ut�nݣ2���N���5�\R���Y�a�,f��dZ�j|ĭ�;���W#{�Nn2�e����� gV��jt���-O� pL��=,�M�Ӹ݊��[�*�1e���2��5�6�#[�p�X�֯�*+�cU���+�9�O���{���ƒDD���&'�v��-u��ս��<� )E%��ڛ}\p���-�j�V�z����m���8�p�j�]�o�bQ���7jV�Xs;�q�q�}� R5v���FL����zk�j�C�ip��n�l�\�p����jSp��Z�0V*�dȋ�Vk���:���k����h#�"�K:B"yU��՛�lX�uq��jT0g�y���Y��Ԁ�5��JT\��\9��f���ť3���Ҋ;V;��9���=�5/A���ĕ�'��"'�i���U�>*������o��=��)ւ�&�\U��jܵ�
̶�Ђ�yZ��极>:*MZ�-Kn�k�CuC���p�����O=��6�i�D),���f��,Ԯ˗��sC[n���j$U��:�P�H�����S�Ʉd�	lȐ�����Ҟ��ڟ�Q��+��Q\���~��}0U�䏒p��o�݈H��ຶ�<��t�8J���u�0�V��r��37�ĄC-�,������wN	gF�6�擙ڼ��#������Z�B�zϻ�J"�|�v������7g[#�zV
�_צ��r�'}%�>ҢUrٶ�� ��m�\���<L��m�p�q��s��NT��.uԑ2�J0�.]��f5�e�l�T�c�S�,�=)�fi�'٘�:���m�2�v�Z[��[�r�͚}�t�yk,M�[q�34W*�K�fʊ��q�HBޱ�7Z�t�9���|ĤK��d�;����P�F�QMWs��c��(}�i[��x8Fte��{N��JN���T}C����+��W�珴/&m�bt�/u[���STV!�ԙ�$���udP�߭pL�)lWj�i��X��9*Q��4����"����P���,;ܩ���rA9�i�%t�DC�V�U��o�N�a<�y638Z��0��Kd��u�a�n��Y��oFX!����8�Yk2]o+6�N���݂֨�qⴽi̱�7;��[C*E9��[k��tp>�K�㴱��D�Ϸ-�kr���H�O:u;���&��O7f��w`T+&�-�J�����[�K�z>t�5�x����iD��2+=:�B���̛���#Y�I�E�Glq�o��r��7�8=�`�Oǰ�Z�X��i��(�(�)�H�(i"�*����ZB���j�ZX�iJR�i����J�)V�hB��j��!���)
(��J��)R��#CI�
D��iv�	�)A��֨�)(Z�R�M	��5����
 z��4�-IB��o{���!���cN���"J�����EݔJU5Hv)4ѵ��1r�\,�2�t��u�o��ƽz�Jl����Wc'�3�;���n�����/�B�{�u�^�6�Ҿ��]+���v�wmtk���m4�^#t����R:g7����0k����d�^���)5n��������/d;ŎZ'%�=�"�����vE�j]L���f��n'�g;c���[�5��q�$x�R�e#������%��t1�� ܹ��ZF#16���'��n�i����3�3��w��e�%F�v�L:�'$���T���c��7W}��3I�)��Oƶ6�l��dy3J�$���W9YUK٩�R͝ON�X��[�vy۲2�I���9�.�Qr5[L�G!;'�v3+�:�r��5uC*�E
��^�bgY����y�Z��if�U]D����exdN��n�p��#RF:�a�gk��/-��f�6�#�ERR�^*�5K,ɯ>[�7�=�0!���=|���{�&���n�X�����?ѻ|��{b�(�R����n��S4&�8soG���Wu��6��9|ZF���'@Ys6��%�|`f����Td͖r�`�p��5�9��v!y�2�S���#�:�t��U�暬���,�߽�q杋K���JN*���Xr�6�kVEbZ\�y��x��~��E�<��vo���e�xtm�J��T��5�D�?�/4ow:�y<	η���[B8oO�{�9�%�s���-R�ɹ����|Ƿ���ݠUt�fp��,3�"з��u��K~ѻ��t���z���s�x�H���rD�Xu�[,jm��WgC�)���ʧ�8FC�ms�:S9 (Ϊ�:��k�)�}�vx�1���te��4���[�uNv�oEHf)�El�̋���[^��XOm�Y��gdl1}!��.�0.V�qˈ֔�������&̋c��[��{��i��/���&�vn�1��ǉk��p�|}�A�;a�9<�VfX�����l�7fϛ9���DV����n.���4ZLS��@x�k�t���3���\�8^�Ӧ�)�{V2��{z�~�ËIp�����k�[&z�#Kz����=���&�ޏ�o7.זk�-�ulN�`*��
�ܧ8ޜ|��8��F��ĹWg�n6��kf�i;|�E��d�*�r�\��ܮ�,�N�`˶���e��D��F�x�u��B%nVS��n�s�H�S�W�G+u>#-7����:La�	�P�P�9|.�b����ւ��HE�#�u@ջ��s���>�Wai�Mno�sz�U��o�*������K(^�U�9�\�){k��؆�٢�\����}&v��F�7dڏ6�J喷�:�,�Q�hYU��,��$����y"jN���Y���徣q�o��Yo�a���&�r�
e���v{B�l�5�3Cƶ�� 9Ms-�|�8E��F�UO7����\;�֗+e+v�[�ו��Q#��C>G�-r4��tV�/7��1�9�ͷboOt<����d�r��"�2Ν]A�`<3}}�ܥ��D��Y���"�L��3B�)	n�~�QhKf�6����)K3׹�p��і�괣
��MO>ޚ��V�,��s����K�j�ݞ�t$��G~��c.N�}��#����/7?d`�)����q��{�!��j;�w���:i�N������0v^�*�燢�.m�у�La�ʹ|�Zh�Ur�`�m�ܾ<�b�*=��%f��t�j���Z.T��Sv��y}utS9ȥ3Y�A H��`�kw��?�_liN;g��WD��̇?��FU��+�{��pF�]��ai[��Ŭ��٢[S
��_���Z������7�k6��j�%��N���{q�q>ɣ#�����0`I�2��SH��/8��C_���{������xG)2ܭ����,�^��M�ֺ/,C��y������ߟ���
C5%b}���gZ��k��a�Q��ew^;��r[%��J��o��K�5�E��)�TͰҷ%�,%��/��5MVZ��o�֘fC����C;ܬK2|BsH�͛�,��8�[D[]�wd����Ϫ��[�e&$�I�� ��W���k��\�P����,X��s�8#���;KmW3��!f�v����g�o�ha�A�u1''��Y�훭:����x�8J[֧$�/r����19�f�3���?�rF���E..��M�;����S��n�]>���-�`�
�uk�]W�
��$K��6�C�a�y��Զ�	��15D�+)n�`V�XՈSdج��{m�p��fʿ�����ΙB)J�J�+e��Σc�µ,6Z -cbR�y�>�����zI7�4�(�t����%o
G6��>(���u%�RV�;j.4�=5���Av��*�H�e')n��8���F�<���߯0�>;.$|��}��\*��l�H�D�~��"k�n���(�<���R�����9#E�`����m�;��'�7��
M�x�`��S1D�i�(3~$�Yi�)�A��[y�̆���$�!��u�\�w\sj������E����t��,���<d�n-iv��j�.�mxϝ]�b�w�}̑������K��h?N��.�m�B%��W=;�8��"����mO��1�Ų9���8�	*���betM���fw�j���%�>��<����9
E����a����e9[O�p�kw�����i�[����9+M���ws��ݒc}>�a-�άOldTy�fjɻ�Mvﵚ�2v�F8���F�gC;9r�S3���<@8׽7���	�I��Ic� ��N�a���f�^�k��^ӽQŘy���Ù�$X���|x8��z㛷�ڰ��S"����P�.��5�kG5�x��ۊ�f*�e0�~誊&؝�[�ֳ{�{6�~|��䣒
�45cE�w�j-T9KTڳQ�u��B����30�b5d0n�;���z�M���*�c�
P�\�Q��t>�qRkq��o�.��ؤ>l񾄲��8���S��,+2fl�Ls$xW"&�#!�U�i���X���<d7-�g<�%Kz�U�mH��#&��a�*�kE��A���pWޭP7w���3�u�Q��Ow�F61�~�#�%������E�����!�˲��`S�)?��\&7Z��$�yț����:ދ����ڏb�|ޜ����:�ѼvK��,ù��Ud�7�ͥk��{��2p���*������4��qLz��A9/����/z�qW4O��|(��Q�ZZ�͑��{z�p	�`�3G.Oa{�W-{v�_Y�B������*G{.mј���G<�W\�I�޺b7�^z�'��Q�3�����-뿐Dջ���+�o����gs�fU�5�h�CZ��C4N���Ԩ������T�ˌ����	���'u�bCWǝ�oun9P����Un��M��k�A������Y�������i;Xl�i����ӮF�+uJ-�L�L8k[��%La3�@Xn�m�y�;��eZp4��N���N���J���c��������e��U�ǲ+�"�wfh�3o�o�Dw6u�A&|
� �:�6���5�T�\��c�kYkOn�/j�L�osC�L������FO��Q�[��T�o�(,��m���]����Y��v���U�f�wYK��I[���l��[�kN�}��;yMo�����/[^;P���{X��TZ�U�U�;A+�*��$*2_\EF���̗�ǚD	Z�m8�	��mA׷;��ޫ�㋢��y��h�0����юo6m�=�2PG �e���k� �����)gP}D�M��s�����F?�ם���+$�����ӆ̅	���-�\��I�%��{~uY��L.a?��ɳ�L����U�i_6��\��:�	�&�n[E����hn[�CU@��5�$[��C#����d���i�h;�M�ܩ����c�F�,͔�fk�}���AXb	]�O�N�<���zۀ�w��r��s]�V�cx������M7$�P�4#�;W1�������=�\o��ƛ��oi��	Ҥ^�G��wB� �y�+���v�����?s����r��p�#����u�����&�*���e�����Sa���2�A.��s�eX��5˳g�oly�n��Ee�c�wn�q���%�0 kk�Ы��1���S)>����t�j5�����o��&{m�+/n7�a�-\� ���>4}�����]w|�%���(�����n"0��}C�Z3q*l����g\`I�/�ff"C�>M�/�g�J���#�u'�{P�+_��~������s�}�6�t��򞤧����Q5چ��O�y7��"� B�=5BKJȌɊ�/��6re�
�b������5w}�^k�EDl�T�z=v(��~ �|%ۀ
���e�ɇ�%�a]r����[�J��[��Oy7�Ib�c_[+��6l���W	
����af�Z����օ.��=��w2A��'�h�8���-�SSV�h;�Ƨ\�32�Dsu�#,(�z˼A�|F�M�M9�n��\smT��K$5�	�Fƭ�����7�E���^�Xq�᳃U]c�*QV���u/o����C�C3�R=x�V��¦�����]��ɂ�+�� �B+�S�1�x���n��9�eqIm*��oulc��E��=*��s�.��f��e{~�:��/	P]���o(�97r�D�7���z�d�& �3�:��wL[�K��%#�.7��}�>�z����I�.'^���Y%_�z	v��p7W��Ljޠ2WJ~�Ѡt��8@=һGUX�l�/Ղ�Z�I�Ua��s]��i�ǯ#i����|�j�Ԙz��-[uM:�j2�=�[`�ń��6ψ�l���8a�&9VE4�5�<�*ɶn���_�ZI-¹�R���;� ֟1�<O��Gu����U�� ��%��:���複Spv;�n��&��"Y/��c #hv�l�iy+�c	��q�ΦxH�qM��b���LD�2��,�f
{��#3���f��I�m����sG�G�E���G���Ջ��h�'�7�-�p�f.=R��I̱�:���K�}s�:;$k�`��'���2���[{Q��qvv������d��V-��s����i�	%[�~��QF3�_Z�7w��$9���XAD�QV/��]���u��u
N����O�+Z�/k�7ݠ���3������r�u|����W�Ɗ��i�qU/AUA��i��Z4�W���˭���(��.��?t�x-� �4z�N�k3L�lD���R�	uE��OA+��5��Ж�D��8v:�fud(�efr�q�Gt,�w ���id�V+���C�cE�Iߍ�V�*��ϙ_HtEɯ�ڣO�Ƹ�[t�@���&yMf�$�r&��pr�]dm��l�d�m��f�t�L"�8-�Ի�έ*���KCkoQ-y�ӝog���jl�^˞���s!��9M�d�Z�s��y#�{||}��o�����{���w���������,����鴵*>�K����M��R"m�,��sw[�@�2:H�P�(;|�{���w*�uu�+2n���l�Q쬕��w�=5��g_$�T��#�.m�1�O�g���8fF�F���qk����m���.>ӓ}����`2%j�cn�*cQװw3�\l��|/Os��`�׎�ˁ�1��R�c+�tMո	�����c�s�nU����BV�9��Pcy�����6ܾ�,z�om8�v���ub��o�r4	[Ɇ�k�����8���"ڼ�:�)Ɲ�:�4�d�n1��x��V�rhրs���]�I3tp6����bIlҌ�θ�8�h�ca�^��N�`�K�Y��(¦�#�f�F�k]L���U3i�
N
���q��F������]��ˇ��Dz ��8u�tXُ�z�]��O|�J��̬@о��٭j��,r�w7W05��Iw1�gkL�I�����{�����zm�R�̽b�5*��#�U�2��}Ջ2���V��*-<�J�����J��f�Ƥ4��f�4	@k��fF�n�w�r�:��J�H�|6])ݲ�œy��y����C�X�(���KQ���f�!�x�,�	��X6wV�S� ��Ԉ��s��y【��݋��DU�s�"hN3U;���+T����]�;�nQ����u�Fu>q2�N=�[�.+;��/�ή{�6��(�F蠻�K\+xԛ�29�����K9yy�ٷm��*bCe���b�\"V���%F7:�f*�j��3*)�l�s���je[��Gb��z���k�*q��KX�9���*�掜.0���GL�Vӗ�au�T;ռ�X�ʵ&�]��SVo@cs0Ptp1º��溳�[15��cN m��s�0l���T��zQF-���M����.ݠ�S���Y��� �u��)H!���4>Jcݥ��*���_p6p�Ll��4V ��C�V3H]��opr#t�41�&�;lm'H�/s/e�0�:�2�[8Q��<�=7��b[���\��6��7�������743rt ��n��Vn�X�{Z�;w�����¦7ܝ%����-�5a&d�4 �h�.����)ݞLU�R�ط�v����8�#��\���r���oщ�يfK��'�7+m��P)��Z������.v�U�P�2��x�e��o#��Dn�
��R	[��]�upV�;:b�%㶦�D�>&D�u[��{[��"�^�u{ٺl��-�!F�!��|*'���&�M��X�ew<vM��mdͮ�8�J2��2�>
V
���BvB���(s��wH�sr�<U٬���Ϯ.e�C��;�.�6h���}��9fH��⮋���On�w��׾��㿣ƭ���T��M
4#T��t��@�BD	CN�)��`q)B톖��ST)�=H���Hu �	Hh�i:�@�=U�о$4��=��dM�@��i�R��'Pu�!�
z�N*���GJu�և�t���J=u�:�t�E�]N��GQOR�Rh�:��:������z����(�4��J4Rui�n�!�1%�Cԩ��记�ء����+��)���Y���m�����ǭ���-�� �0���N�C0�1�4����ox(^΄c8��w{�ӡ'm)̕\J��
��]����pN!ڦ�D9�N�:�7����,��ȍ4�,)l/Ȣ���d1�q�"@#��s�o��s�:wx���B.e��|�faֿ�W�*��|�[y�E�6�	y�=�K,%ź�>+/�Ǚ����i��N�f6�E���3<�z�*{	�o�n��In�y'Iw+>t����&͗�ȴ�v��Wȗ���<ֻ�������]�J�Q�3\��q��-MN�ԥ�����n���
2J��t�;��j��gT�n�ez�k������kt�h�.��������wt�0�g�?�6�f/�F�k��e����讐9�:�ގ<�ᥟΨȇ�ҰT0��'v�-������2�9z�̻4��R-.�l
��T��K�l�s/���nY���͎��R��X�	�VBV����_���嫭��~�ؓ��� �_������بj�z�Q���z���O�����'�����2�6C�.�����9S�~��fT�1h2I�\�3r��hvz�k/1p�ޑ�|u=+I}�I͚�*�t��KP>�c�����n���sC�z4of^�îq�^P�؄sV�\�S×�����L0\���N�����\�l	�;w�[�P�{���uA����m�
���KM<�,�h��Wc-�
��s�c��:Aߟܧ�kz�{�tR&�i��u�$Q=/0�*��fO������|t�]HWxW��wg0̘%傧��eL��W.��x���Nk$ݭ���'�@����!m;f�-�E>cl۽ԝ�����&���IS)XR͕ו��꽽o.&oCA�;f��2����vpN���־��Ƚ˺b�7��A�:��0�}���D�Os5u�tSM<�c��}͘V�R�vn�������9BO�Z7a\mWD����p+�y�=�z�d	���T;�[`b�J؇�f��`Z��*���"���;S��ݭmS�އ��͡�}�Lv�O�hntf�8��h̪<ҕ�����-sl�3��ߧ���Kh�	�P>�WWN�R#r)��.�0�9V)xU��ڭ+-P!��({
��-��`��M����TYN�r��t�`ގT��go\�čc���3c�J�v��
��I[B켾�N�|��@鶆�T����jͤ���M�*�}�]��,�^(��|�o��e�\F$V�o	�
1�!:�=p�;�i�3fK�s��2O�fqi�뇤���q�}�)���2�H�[��-@�~Re�[��ҚCz)�J���ӕ�vhq6��6S�u���e�w�qI�͈P��3��`f:�x�������
�*�	�iX5�Sw�y�_�2y�kG;iowa���i�l:�\��L�;R�9�UK�u��=��u�� s��z!>�����'MM�Ê�b�x-���ܺC��"���:���s���9�Ǚ�����).�	r���UuVq���Uo��_7C*�%��z��yid��u}�@?A�oB8J[֊�qwqʶ&�����ݙ!L�`ʜ��s\�ci�`�����j�$g��q�W��WH�N����71MI��D��8�UyJ[0���cۗXڰzx��
�;�_�>e'��WlB����ckt>�4nn�L��
or��L�2�e�M�9�r��l��[�f�R�s�j�s�m�Lb�6��א��o���f\���P�oLn��u��aj}�n�%��#�� 2عս�6�]r�6�w_D��2�7ܚ��pO������`��ar;tܻ8k��Nػu:{m��\Ow%Ҷ�g���f�e�>���ز��*eШ�����$ d�yk�m�8�H�!M��l��Xe�%�f&U#e���wq~�1�5X�(�k�(�����9����0��uzg�/Z�4H�e�ݱB)�k�>��O�z6N��6��ǚ�F�����he����M5�a3{-8�|�Ո�E�_L����N�h����a�K�ܳ�6�[@�o;�!�l"qُRa�i߯]Urf��=.����<%����f�{cҲc��R�d�k�G
��v�0R6|�sv�S���L�n����͏cj�.�Z/�n�(�P(��*�,��H�n���d<dN�gV�
e���ʫN�����=Hs6��5B�W<RԪ/��y��ۈ�
�;��s��wI4�VWꚫ3*-�7X�����}�����~�(vZ��q�G ��(�ʷ�@��d���4������e[R�E�&�P+K��q���RW�dU�3��8*<�0��c+�*�i�J�=��b��	�.s�e������(���wZ�#$�>��;��n�7z�`ű�"V]��>���ڣ���Y]�)�(���fL�V�i�����r�����͇�,�%���{�,4c�q��ҕ�jrM<��ƻ<^;�A�l� �N�hrzd���_
�F���uR�1���V#S|7+�w۲0��Q��&�$�܇{��4?��յ�#��B���҃�֑��/5��֓���V�RΨE̱���6T�	��Jt,�K�z��i���W3�s��䓼�\��١ϙ#�����nG�d)�~�5���c���I~�J;cι]��k�k�t�r��¶��M�-�;�*�7l�{��nBm��M(n;�J��dFg.�'ln�T͚�Q����/�q������ۇ{z ~��d�R7g2Vy���'����M��:C�;Ձn9���cQ�� ��R{]���F`,3vcqm�}o�!��\�f�n�s�|iQb��3v��һ�P�O�"�<��n���R��*^ӼI�w��Vcq�ٵ{�*z�s�g`͈��*�M+�q$���B���t�B�}�m�܂pK�(h��&,�*hۼ<ҷNb��pY�h8��a�f�WTS��=��i��� 󮃐�l��b����e��k��F�E�Z:7�5�O�_�\�;Ű@*�����7�T���G��������݁mn��7��FfKϷO�4���m�BV� r�\1&~�kep���Á�k>�j�;c��"��i�;p�4P�	GN~��LrIfm�OW�LS��ٶ�Q6O��CLKҫ�:�=R�*���T-IȤ������G-���5StM�£�1�_�-�1vri�����֒���Ϸ�2{����8��ʶ�̪c��n6���
3����#
x뻷l��������w|P)��+��c�Gz��I�[\�"N�Hl�S[�˕	�d(��oy�Mo����zCrH�3|���u���㷶YOfle��z\�>lni�0AR.�>y�s��L��1I�����Q���B
F��	���$�j;���ǽF�`�\,E�W��{��fl���[@=��9j��(�Z˵[�8�]�"�r��N�i���Z�C��C6l*�X;@O��*�pA8T�mц=�2�yݱ5tz�>��}�Nٔƻ��%���j��X4D�Q�o�Ʒttr����"5��羀C���������٤���-�0�;9<3�:�/�WK�f�\q{q��h�S���5�ٮw���4�ޛ�r+	�/Yn�D���N^�6�*�r��jm��7F{|WTv#^�]���y͜-8����{G�����T�ϣ��������a�Xb4�{��8"�=-w�[����#�rt�5�]4��;Fl�/Á|��ngU[۹:�HrE�uW"��0j��Y=�[�����O�[����t���X�_�3��B\�Y�Oʨ��yX����;�CQj$�-1y����3�� �S�X�[�0k+�{�-�G�q��9~�ך;H���Ys��m������I�7轃�JW=��n�Y�|���Y4ފ���!�(�#�}E�952/)��㥶M4[�t�w��-2q��`^���F	Z��$��b�.�,L�ͫzݚx3�E7gS�7���X;E�}\Y9+vd��c���2���'��<!iW��W����m���#�>���b����w�q"��
ʔݺ�>�S��+J�)ou=��O��67�����ݎ\uf����N������g^2�k�Z9Cs#�a����z��_��T��ބr�K�~��������m^ێ"8g���D�������h��!�o���$���c��҄ȍ�k�ik
�L�Cmi�m��A��50�P%���oTY��䷍"��FL��G�`�LpΪj��8v;vz�	��98T2����>��)cOP9�Qۗ���]����ب��S�B�4�zL�:�ّ���e��O��F�r.�ik�0e��z�ܖ��;�vդg��B�g�oC��@g��;+���Y�t��.��1D4L�Fb: ��]�p(�ށhLtfo,�@��"��;˴�D�[o��^R�5KCW)�l�e^��}�t��q�2�����c�8��P���h��f��q6����j�6,�v�������w���fn�o͌�V��]$3KuT(e|sԦ�M��:v�a��wlog��<�"�\��j��$ ��tW[jV����8$�b�H�7N;����r�3a}vnt��"Nv|½W�%����B/#S*Vr�6�MQk�:������G\�Jǹ}����ux�2�|]�O[f����f|����Xd��[5�n�tf\
�+6�>i�l6���i4�S�����a"&��M��Z����[]}�]�2��)(�R r�Y�˭�l,�A�`��ʕ�u�Om:�B�k׶D�!=�ʣ�a��f��)j/+A�*�]�}�d��첥��c�� ��x\a��Y@w �9���+2�.3S�]�>NYp*��H�v�%�˅ǚ��of�����)Eq����6-��+�Z���߽8����e �-S����]k�2]q��ѽ�יO:La����g�)�
��{�&���z�)���d��`�n�ˤr0U��e�[�-���0ct~��1M��mW��OyM[�\d[�3�UJ����d�4����9�A�9�b��~�-2�^���t�ō��>��9��`W)s�͂g�8ۖ�ǑÚV�U�\����F��޵����4��eX�>�z^������|��Ǜ�=��W]8�J��߈�a�C�ğM%g>|sogc�z�U���N�\z�oY��){c����e���zV�ɯ3�v���2�S<jb;���}�1;p�x�If@��Y���4S=S�ز�yS3���O�mA5�u�b5*;�ު��Y�2T�`;�1��4Ћ�s ���4߆��ls�(�m�*=��kß�`"�r�Rl�Ր�U�2�^=Ͳfv|M�2{_�-�w>#>�!a�3{x����n�qvH��+Z֯rO���d�m#�1��ΐ�h
����/f��5��5�j���(Y�ڱ��9;C�`��O�ө�lR�6Ӑ�*��ƛ�O	^F8��Ce�U�1G�ֺfKϷy4�FI�Y)[�r�SN�{���G:N6V[�獀�M����7�=�B�I�E��A$9����퐀����%78�v;�n)�k��N
�Z���@��������ɥ.3u��}3u�gs6��J��fW��W,����>�/w�����{���w�������hAݏu�Ϧf����ٷ|��f� �\J��9�h1�1,��ȩ�i�ܭ'6�@��{��;�D	�fwo;�N�������_H�3_�YbAkf-�M��@������Ymh͠�Mӻ{e�N�a :����H��%�$i�1b�/Qu�$_*4s�u�+nP,1��Hv�����t6��a)�H-e��Gs���o]���k �{fS�ft�U󹜥ou飪����(�@���t�7j=c�i�45�Ō�u��v�j�`��6��6��F)8�#+Rc��S�ʚZ�����k�@HA�s��j�S���e��i^g*m]	����m�E��!�G|�9͎�K[����<Y-���îsOAR�14[t�.�k�[���M�f"��]�+n!�;ov��f��V�t[I@��Tö��"�� 4+M�L�0�ɍ�u��� $��
�cuSIe�Y�S����)RYl����lꫩ��;���$딷3
�
$���'m��^ 4��@���Xd�ok�*�J��q@FB�
+��H���,�i�Wg����d�]�R���i�����D]�����n�;���3�syN\���m�u;�tdR�t�u��㑧�w{/'h�-�d,��<�.n?�@ �].�w�˴�sYYj�J�U��f�����3�ʖ��O2ӿ���"�����V/�=%X�A�:WX��| u��J�r� Z,j�i��8����Ni��я�r��S�̹����;���g�������},TN�����/y�����t+[IB�	�����3w5"�1f��5ݼ�gA��җI���ŕ-X���\4��ǺSS���`|�+텚�ma�c;�_+*I�Ч��/��*୦v��I��97tS��Y5�^/5��V�;w��ꀶ�ޤDz�Y�|�&����8n���> RK��c��9nrS*Q�8���J,w{�ZwB�z��ݑ�]��:�W��.ld�Cz�emƺ*Ĝ��L�!���vU;����bn�2f�PЬc,�����z��˶�/�GS�]�ρ��Lxhe�(�����>�IvĐe�n�ƖEXM�қI^��p鹒[ZT�6tA�JTF�6��e��.ܼ͙4p��%;9�����D7��]^v�/1}�7t��貰�Ži��b�E��p��Є|w��ʳ����N[�e�i� k6R��}o���},b���I��CY(��4w�vA��c�÷�橉�2$��<��������-ݹt� 1.�b���N����1|t`1e�[���y�.�Mо8��ɽ�����SOLr�:��<"ݙ�fISNa����]%�{o]1�q�m�wD�4hȬ1��ͽ��:]w0�N1U�X�4yX�'V�"jE��K�6+ɋ3�"�q�Ej��[�v�ުSEٝM��52Cw��{��߯6��ώޫ���A�P:R�4&���P��t��t/Ph�.�K��KԦ���
�MU��@�#�=M���:�z��@u��������ҁ��N��)���M���	Q�@�C��B�C��4���{B�)ZT���!TU-&�4&�ЄJ/RQ��M%#�(��D	E	@h4�&�IAM&��CM-�t4�
�
H�*��T�AHĄCHL�5T�CIC�AAESM%U4�TSP�!B�S�E!�)��'�r�s�j1 �{{W�}�"�U�����V[�fgR�&�i��Қ�@����z�x���;qb�����XUp�R���/��D=��n|/M��vAVj�X�"G[�m�	�[�㑕�§�i��*�$�6O<F�ͮt��d�#�,޳Y>�ky[��2ٗ���|�3:�V��f;�ࡣ�K�NP[ Y���]M�%�T�l%���u������NNF{f�/Y��� �3�=��j����������q$�F�5Wf����F۸�;4Au���l,�=0�Ϯ6�U]�ď��fK_�}S�G�Ln�!�"������������l�BޑQ�����kwtL�0�����]�WƖ�o�Z�dw��ρ��1]1ڋ^��OZ	`ֳ��Eݦ��ZG8��� N�<���y���:*s�{��~���Z���)˰"K�͑��V���	ިn�<Lْ���J���+se�d�ߠ���"�O����p��8�@��B�I�/c��y�7� �ڹ���<��PF�����7�H�B�`,=�Q�6on�O�Cei�f��2.�]j���ջ����j�Q�|X��۳����bN��6(5Q�Ws{,�;Tl��[�y���5�q�v_p����y�S��9u4����fw[� �Y���a��,�;���fbo������w��e��9dGvl�j�!�^P�}O������e��`��ѓVx���O;]u��f<Әd�w0���/)�[9S�_H
�
�j�v�R�jDt�TԔ���wu6��6��ö�֐OG�5=C*�n���j�ˬ�h���-}B�c��4� �U���u֤�R��^JUuf.��u�[��B��ƛ�֭O�/]��>�FM��kM�@s�8J\�m*�ٹ]b�:�v��}7{����YT��rlr����ǻ6Ό�';4��z,+h�ji�w�&��u������igq/�d��7O�.�3y,��i���L���]�Y]����5�h������r L$J�i�d�~��Jμ���PÝ�:������y��'}��<�uPH�s����}����@Czo_���d\�͛*��8�����0��&�O^����MF�[�o��6`=�w�WBjJS;�uI�=�&x�A}DT喛I�UĻ���*m��}*"�nf��]��v�4q�W=�����o����V�E���dB�9�y=����*���<1&�4�l��Q�(mL����um
0c���~�R��,c<wVZF1
m#7<��5�me��(��5[;����	�	���6E�o���&;�'yd�9�JȌ׾�]Շkd��L��L����}W%����Ն�N�H'�:�D��|�tݲ��dq��ɵk�p��\+9b�qn{���`�:.���؟!%�Z]�]l'a$g`&Jp愻�}/�z�,3T���2��%ߝڶ��!q��e�����]��I�r�\��b��B)��[v�!`=C�[�-}�$=�n�3 H�rCdr-������n+_�UT��&6�Vc'��a�˻������FZ�y%-�%s�����j��t��Q+;QU���Q�����{���3�#�6ʟm��(����mj�����䗫��۴�3<Y��x�vUW~}Ms�ޏ&��|�P�)kz���JBL%�Ɉ�`4�3&H�®��	��l��p�*ה��0�N|)��-J���'��ۜ�kz�ɼ&�b�o'6��<�s���}	���n��R��F��D�厷�p�l�7�-t'ݛ'!ƭ2��Qe`�ۺ�\y�8��b�n�Q=���ə�?W���ߦ)����q�;�+�_�S�~��\��f8�	��#^�J���[>Wy=�)�6a��w�����!T�4�ʼ��Z��u݌�!��2�5e���uƘɴ�7��Y��O��g��qY�U�&c1m\�"�}[��m)����,��M�U۶�Nnye�%���D�C�k�� ν&DԖa�,��C�Ms�sدތ�=���3����	tI6��T	�g��,�MM�����<dDjU3���_%S|����R�I�E�N�{Nmݚ�O�NH���;٭�A��+�=�FJ��x}u1��)���G1�w�o�'pZٜ�z�t�k����F"}BB�ҫ0K�(���q����s{c&��I2b��:��+z���j��(\�8�熓/��(���=^u��=y���:�M��`%[�4�/e�g��`��3�V�rЕ��]�����m��6�!N�T��x�N�_c�O;Oc�-��9�i3'mJ�z!"��6�ͻ'��;,j{0n�*}`��0^8�v��Ep�\��ckju�§Q)�e��WrIo,@�������.�*Tŷ���x�0�G����̗�-�+��:�
�j~���/x��taW��nn�ˠZ��x�jU>�FDMѯn0|��J���
A9h�L������1��/Rݡ���h����륝X��SWMߧMT0�j[�Z��KC�ֈ�8`w���r�R��!7L��v�0�CaAݻ:�kF�D�ܲ����1�^:NكtT��Y�Ecǲ�N����KDl�}�㛴 j�P�M ^ĎoY��6��,Ȑ�Z�lȷ=���b�^2Ӑ_������l�Ё��7R�nI �fj�L��Tty)�4`e=�Vm���q|��rC����jlT(|�|��7�����ucN�Sd�7[̬q�)��uSh�''����}���66Ү�cq�� �c�L�%�;�^W�n.�d*n�����6����9F9��~E�2��4n���	����ݘj*X�˗�q�-LܫCl����5�B��O,Ʉ&��V�Ī[���G�\���N���0 �׎^�e`��Z�����JLn4�l��Z�[ZN�:Np2��c�y�g�% �.m�(9:�ҙ�c;��4��9}/M�x����c�������� [�z�x�lXoeu(�?9ױ.���;��"��A���Ֆ	��m�3��ߧ���	FVb��|R��z��±�m�pj��)=k������M=�v�f�iX�YP�'&�7��U8���ͫ9P��fb4;�/Ÿ�k��L��1�[�nfI2LcOA��/��a<RVd��X1�ݗ���W������[a�d��k;Į�A�<Y�Ou�K�o�T����iH���v{��VTZ���~ᱽ�ь}d��x�T�V̓�<��v;HoC���m�]?QǆF�5T/6�[��\x���y�#�MM�:,w���U�F�넉m��ZH������F����;�+/�R�Ԥ��
����~u�YbH}� �hƧ��3&B����@��#�����׃��F�ĥ��U�W�����
�n�54Y�g;i�}��&g�L�Ď<���R�ׅ}qS�.���_dnB՛ON�\AM�\��s���>�X�&����,����n&��[�w�Y�ޓ��&�{�][�U�&%�s�t*G0v2�7�É�q���|3�u���Pѐ�:�}�1d�9���n�J��f�W��*���!��͖!+�"�x��θc6�n����.�XL)Q���G �s;��Ǎ�ڃ{������t��.��{�`�ML���t3�z��VI�n��k��a���=n�:���mԫ%����E�+��Z����/\uO��I7wym>ϸhv��z\���]9Pw{k�-�����4�w�Жxu�We'�%[{ue�q	m�!��Z5y�!v>p����45�1g�
Egw,W��k�Bn�L[��P(���������i�>�$�q��.TlZi��r�d�)�{�opw{ػ�}!��_�ɞ�u�N�"z������7��z��_n��.��t�f�M�k�i.�%R�4�_H~�d]��F�y-��ϰ��{�$�4x�#���x���-����:�^�jP>�ݯm�ne�C�W���[w���W�K{���A"�����X�z�{���ֺټ|#XI}�p��=5Yk�3�s���[s(�'��r���;��q��/�d���y$M�b�cr�\�j�9���t��#O�V)��1vS���0��k�KSPl�����&�w*�k�l�˟�ޮ�˻��������ǱS4{M:���v ���I�E����x�4�~W���j)���+HO>��U�W�c\�|���e�����E�����Qu Y;n'�ؤ�<�א�����=
��\)AǡW ����2�Ulte]���9fVm���j�n���ܛ(Jx���c��@�s7y�Ⳳ"4h�z�#��ً�	�TVd^2� 1�"��ݧ!���}���d M���sߤ���7�����guG�o�r�� �)�^���	I�1�������E�gSGqF�:�^l4qg�tx�z��!hlr��B�`�wg���@���az����I�E�'~+��t�>d*��N;���`����r;��(Nk����}��U^��\S�AwZ�sF������3pbV�w�w����k�D_u<��5]�e�z�]KM��9�b�����<���/e��S�"[�xP9C3�z�l��z�'  �yt�}��n֍��ܟwSq��>�(�$X������#d��4�[�+��;�U�aN��/^���P#VWB9p<O�ۗ�Ds��9�m����̤�UM�9Y�	E��o�xC���pq-��*�]xV7�ٖN�Tuv���бQ6�[��j*;V��٣�LF�A�w��[�]����~��7�%E�f�c�f�s��.~�z�|,O^��Á�����F&>�H���j�{����ԈD�c{vF�m�=��)��)� ����,�Q5[�_"`܂Mp5��H�x�r¬��C߷IQ �,�Z�;W�4�u�RDc�ƚҩxGC��O5�}A(�'�S:�FT�&���옃}4bƉ>7:i��6�-e��}�]M��z;�D0qߛ�?y�� G*�'��+&V[<{S.��pl6�� �uI�����l7+�ܔk_n��K$Q�jʭ��*�X�*�l�6m3�U�N�^U��*���Ehɭš�2^V���r$���vP���5J�y��]�8�6Җ7^��"ҧԱ4��X����s@���-�@{GI��rm>L፜ߵ���d�S]u�����J�c�.[�jT[�+�oA�c_r}�+ޝ2�lQ�B��j���1��Z��=�n�����8ڌ�)�rr���I��2�b�������ە�����K��$o�[�wR��ኞ�L�����{� j�G.mn�pi1޷�ֽv������:�u�p�$٦��^a��Z��xD{���u�wmQ�D�c�)�щ�ٵ*�{�����H+ҸY㻻�!�:OI�ТЙ��{q�`��u��Dmfٶ�M!��g��>�˪�$��̢Ve����jm��vg�o���U�wys���7��*=�s���݋,�YB�6�3;>n#��I�z��5�Jn�+,#}QWL��4K
�:�i��G��Üu��j�=�ɉ��g�w�ԕ�?9{"0ѹv�Ղ�38�/�%��t�ۙ�34ΈE�Oo'�hx=�i�T��&[U�WCi��e�B�17ʰc��r &�#U�e+ٸ8ѵ7����"����6���;lQ�Ca���s�7�������9� *�ި��{���
��H"���}GG���>�t0³̋2�ʳ�2�ȳ(�
̫2�ȳ�+2,ȳ
��2,��*̣0�ʳ(̋2�2,³"�2���"̀L�0,2���� L2��3
̫2�0,ȳ̫00,ȳ�0,2,³"�2��ȳ �+0�2��� (vd3 ̃0,� �0�3̃2�3"�0��3 � �#0,�3 �2��3 �#�=w�'�ΘFe�f�d�f�dXd�E���.e 	� &  �@d@	�@&@@��a	�&U@�Aa	�& �Pz`A3  L ���v�U̪�� 
�0�ʪ�0 ʪ̪��P �UY�U�UY� &D �UY�U�UY�U��g�Uf  �@d 	�U� eUf	�f��VdY�fU�FdY�fQ���=(�0,��*̋0,ʳΜ00,��̋0�2��� ����������4��ʠ(�����G��><��>�����?��O�y������>^�����wc����������>/�  *�s�?_���tQW��  b�~���� w?Z~i��|ߵ�  *����s�?�㤀���S�~O��'��o��P�s��}�PeP!P b )UY� !�U��  	 �U�	@@!Ue P�U�!Ud%U`� "  "@�H��=��	����t~	�D@TZA� � ���������~aA����`}������  ���`�}{�������Nބ���>��v?w��}��  U�r�?1�ڞd@W�  *��?G���!QW��?��H��� 3�����{/�<`�v?�o���������� ��O�}�_���  *��}��y��~?0~����}���I�ߘ?�<�@ |~!����� ����v?(w
O�;�S����~����.��	��I���  *�O�|��d��������8�'��E~�������wEEz��'�˻��d>����e5�g@?Ř ?�s2}p#���$�
��P��((PUU!$�
���!)%QRU
@R�H�B�
!H��IB�@�U��Q!%P
�UJ���H��
PEUTDE�T��IIJ@TT�D��	
D�H!AUR�T�:5(B�	�*�HH��R��"�	PT�PT�T�P��J��TIH�"J�A"��*�RA U(�)R:0�IW   ����kkI��P­�P5��Ih@�%[ a��)�*�R�������3%�iL�M,��Z�ڥ#F�a6���T�f��(DA*����   m0�С��CCB��, ��
�B�'�
�
(L�C�B�
]�ͭ�Ҕ��ڪ�SBʶԴ���2��HYl�V�T6�5[4-�[km��ʶ�UD"�%PT�	
Ep  �sCmZ�06ښ�)L���֕S-ZSZjkE6�JZ������cm�c@k%X���RڔC6�6�Ȇ6ZʹP-"J�P�����p  3WJ��P�i�*�JJj�ڴ�ڡm��e����ej�,)[H��V��j�j�f�*�ڴYM�h@�U-[j�)U
 RBUT�� gR$�l�Ҫ m%����$jUU�U�� �1�5@�He�(h3I� iIU"��QQT�% 8Ơ�`5@-b��3T�ѡHѴ4USjV4cE�֪� �Ơ5���ʊ��iT)$AB�$*)*(p lu�Z�C�aUTбEE�ʭ�a`6#jգ@ �L� m��   e
U
 �Q"IDI. M�  ��� !�  �`  Z��  � 1` (*4�  h�@  ��T�TQUDTUp mp  �� �Ƭ  �  4,��F��S ( Z� !a� 4�����  �R[h�
�B*�R� :���� �`  -)� р�` �j���*� )K�  a�)��Oh��R�  E=�	)*Hd 21���a4��M0O��)   T�i�  $�R"f�T���l�NRACD��AL�ig�+�E�0Gr��ϭ�����׵��;t�}}�����Z�խ��]y�?�mZ�{�ֶ���=[j�����խ����V�����[_���߼���n��?�n�26�٬�jˢU\r�4f��ڈ�Obj��#;hmdlY�Q=U�$r��j���j��Yқ��B�3i�W��kC2�ڨ����["�-�u������J��yVӊJi�3W{u�RxT�x#P;+2�t �F5n�f��:��mK&U���J��*�n��0t$
��ӁMc!��D�����nD�`;����(G�U��o.��fpe #6�m���ƺ�VAgs6��(��3i� �B���HҨ�+i��!ʙ[���kr�hL����.9Bʶ��6l��v��:.+�]�h-����q�4��F5��P��ID��7ʛ:FU彬�:hQ��Ą��n���ؗF�,1��Azn�H��#fQ�y����+Ţ�TE�30Qy�����n�Z��0�
�i�>m"h�t�Y����7J�7EnTd��يh��V��6��{�x�β�ԔLT,�h⦞�)�0��D�X��Q&�A���XF�ј��W��ŕ�j�ҜOvck@�73s6�����5
d���U���WXi]�nV�\ʹ�,&mޗV��V,iok^h�!T�E,{�XV�K�[H�ˤ��kD�)a;�g�>��pJ�h������N���0P��V�:Tln��O���M�X�r��(@������׭-H5�L�Z��Be��t�-�=O%,
�X�z�圬7��\X^%6�)h���+kj8�����kFf�T�h�����y��ʰ�Xj��ܵ��tbʲ��cT�M��.�eH�V�l����L�w�g�W1�ct���X�;F�	�Aӏf����/b
��SY�V�F�RY%��yz��5mMN�a������ށ�Kd˭FAQ��b����,�@21,Q�Ve��L�]�La����mr21��^P��)WNf�!� )֘�lt�ܰ���kV�lQ1Y42���^휕ȱ�Sn惊'@,�P�Rf�Jha�Vf���i��,����I��p=m��T�(K�f\ҵ�2UӋ0o�T���
0�t�I��Y�չNk�6�j�U�Y"i`(&hJ�)zC�n�ɧ۸ou����,���ڦ�;���1���úL�pnӹ-®�YJ���B�׷R��֤"�[��Zi\��5
nHۨ��^���a≝M�ݩf
�Y(�P�lMn�^��f՚����{)�7rݞۚ�KDL��2$��"�*�0^R�3a� +YM�ǰ�W��2���Z�/0��ǔ޽f橗L��tWIm*f��$ˎ�w&H�B� u[,Ö�X�Y�T6 �:��P1�4U����&��V3[vcifTh�G&c�E�j��0^�Q{omK�0�ldhGt'*'j�kvh4ݵxi!b �u�٥�Y���b�%�EɎZ��D�[�dWjܷ(������̖U`���y5!{uE�MS˔%��e��Mu��7�ƯN�E���*n!Re^H�V3RJ�VE��70����%d��/T -뢃p*;B��(*xŇh�"`Yz-������x�9���Sc�R�r[5�f٠,=�a������#�\2�ay 3��J����ۈ���0s(K4��+m�%�Wt�U�*r���D��1�!��n�4�ZQ�ǣqV���H@tӏt<F赸�Aj\QVf�f���0F�Ŕ&t�H��fi�k 2���ج5wM	/TQ�/1n�kv���^V�U�m�{�klQݕ�ee]��'/4̃r��`�e�����Nhf�n-�ZB��4�%<�m�6�&���h�śgY.��-*��ؘ�a���Me\B��`,ˢ^i����[�� DaT�ݛTP�Iʗ����+(��LV�2'�C0�P�4��RA���K���	�g@yY�!D9xؔ�m�VU�:�q�L� (�Ku�@�۸l�
	i�$f��usG֨�3`l�w6��9oi[�0�wAZwM+��J��-��3X,P`m���b���
i�%[B�9�a�Z��e�f]�$Ԡ�f۱R�>kV�.
Y�R7��F�ɱ�X��-��[D=Ѹ.�q�$YM�t2��Z�����m�����z�N��r*]�2�$���(]�n����]k9g j���;��F�w2Z{W�kmAxhF�7lʱ��j�����J��M�;���l���w*����Q�èP�%�*4�Z^�M
�QQTmܚ���[e}��E�R2BuEq�����Z��H�[�_ٖ�D%=2#4Ј�x/�Ε��X�^��Z�ؚ��iAi��M�����r@�(��F�PB &�Z{(+I����&֛�����b�Yk!��Z��T�]�[�7J�$��rm��@�v#@����f�ǘ�b8%�T�R��Y���R��y��v�,F�"�-GU[���n�Wi��e`"���ZAQG&dU��5�Ȩ�k�]0���y����5�{���Z24�IeE�2V��<[CNnD�kXk7w��vv�j���k0 -���,����&��LN�������6^H2���ԋc��ij�^tꔳ�9�}Bi�Ld�cK7*ݡŦ�ә`[z��u�oS%;��[ g~�N���L��ʊ�*!3n�r�K3N��mQ"��j��WQ
z�f^�T�&���Q����]�lщa%&�!.´�!��GoE%u�e�0�U�t�2q��i\�"k1v)P�V�����8Y����5�sm�r�F�p�F?�]�;�آ�H�v�C��olm9�2��)�.R�( �馳k"6%m�-�6Ŭ(�D�t���3)�Q��U�����hS/�N�ܸ��"��嘩
X��WpƵ�P�S+^ù��#oN�9n&:JTj ,l�-�8��Q�N�F�|i�JU
��ڰ�8e��������ɹ��V����Yl�mҼ)��or�mV*4(�Z�0��n&tf	.�������
�X Ս��E��d�w[Xj�]�[H��h/saN�:,�Tv�Ku�� 5[[W�d��d��(����+j2Ï7j�&b�o�oFb�)U��b���t�`����n*��׹���Q�N�c��	���C�v'&ujx��a]e�Xi�esx�m<%9[�6�n�aX�Y7��`���<��#�>�c �f7�an��6����.7�Tn�ǹ���
J��;�
-j�03�j��Y� =�Cc�����vڲV�r��4T����լyr�R}ȃO+-��ȉI��W��bѤ�%�b�����N��
̤�#���M�Z�)�6��T�yv�,e��x@�(�[�֪0��f�YZ��c��;u�47YZ�a��lmޙI�VyB���;ڛ�R�7-�*;�N�.�b�˼H ����ܦ̓j<
:�YV*΅�@�e`��u,ڴ�t���mĭ���6�`�)뵖��xj
��.:��߀��A�+��8r:�Z�D��#r\/tnQ�#EJ�.�U�9> �f�#WEC��M�[R�t�G6@*��]���Y-
�${j�-<�4�X,��v􋠲1��Z�1��H�Pim���ȉ��:�ٲ�,B�嬥�Z���fc����	
gmZ;�Yp:>��T��\w�j?�Y�`ܑ�*K�fm�.�qR�/4�c�iSsu���:�$͆]v{nL{l��)�w�D�e�
m��5�@c��+���U�A�V��顸����[�[I��VDL��߅�b�,�&	qaK2�N�	���v���E�BީkH�-<(R�ŌVT�)m2��r�c�(�hf�i��Sb������hL�F�t�:��R�2�(���tc�դ|�%����^��+�20�0^U��U��a��H��B�,aT/)
s�*'u�S�^ūH(��Z�!�.zجh�r��Ǧ"�T���B�z~I*����ɧG^i)Ū�IKW7��rZz� ��czIce��A�L�1�F+9O��'H��e�@=6�*̓U��A�f�Y����	��c7J!�r��.�b���Z�{ì��Pɫ��1Jb ��̷�i-1�oF��[�Su�����7[�YNb8,��%I��R.�SS�[U��P��:q�jg�l�tK��W]�Mi�Ե�@O�8I�,�-��S3l���-�ܒm�n��ʽ5hK@:���
���OX�F8���AɌ'z�ol�F�=б�j�K�0��"n�p�[��e\l�6m<�n�6�)��t�V���:�82�6��%�"l�6�{>6RO��M0J�.��7Z[+
��NKҤ���2�{���hc�,�kľ�.T�m�#�Q����*:��wAbBJL�*�`1h
��y	��*[����T���Z��n��@�
��ڌ� ��J�, ��M�o�m���� �%EVb9�;Lj���Ow
�)kXCA��,?�ҧ��f�3i���*��<����N��������Wx@`Ӓ�	eVnV��I��CIZ�������K��� �B;�y�������ҥ�U�Q�m����5�05�͝N� 6���l�
�(�vm�Ѡ����P�j��U���ei:v��V�m=1����D�ae7L��x¬�5�JB���x���L��[Z$eX��R7@}�K��)7w'Ҧ�����F�&���Q�Z���b��۳%�F�X	U�vE&Z���C�a�ޫ����0���-R�^jW2�����@�c�ԕGs����A��B�w�y��X!��J��h�bY���[*������0���;���`��òd�1�ͭ�0j�5g1\Уˏ(D�;A�+5[�Z�aHQ��xwR�f3N�ċ?�U�-�*�A!�R�4��STf��֩�Ђ��2^czj�m���bm�qnŒ�sK��v�]5E�6�c���&*���b�'l���*��(��T^`���j�Te�j�S�t��L��PIS$��6�\����j�,���b��[��)�;�L�V�:nWI��N��ven]�Ά�(�dR�����O"�&b�9J[IF�h�B��7��ϭ��� p�!P�d�b&�V����y��fԵ�RK4&�'))�O!4ȞQY��v���$�Zz�Ѐ�w`���u�EKJ��J*- ǰ,R�SW�D׬P��\ [�1}�V�����j�v��" @,Z�P!/Eܼ�V#Gi7P�V�e�
ʐf��JVZ�n�-$"��r�'~�n��w��i�V-n�3N���Z^ed����TC��K�ѷ@��YҲMP�ӑ�Fc�enѬ��Q`e�+30dN�J�\�+1�YE��Y�O�n�7��L��:f�M��4˨P�e��U �4漎U��Ru%���V����L7&�6�ٳ�KU��a�G^�Ql����Mb�&輿�=����z+:,�o{F�!�J�͏VS�q������2S�F������rVE�v��4���f�+v4�B��kc'E��6�K_C[����z��}
3bN��
���id�D��"Ж�M˔��'�+-;��&Ve��`V&�Y%�T���Ml�������w��YkPs^�E��%"��aRM�9*[�'`�J@���լ�/(�����3�+�0U�|�e�h����ɣ�B�f�X�/F�P(�+U����"���	�F­�¡��Ơf6v�YX��Jʼ�Y7�;a�T{ud�m��m[G*�ܠ��X,��3���i���`��0lІ��aY,^��$�@����g��7(�"%���� �2>X�a�
%m1�1˷j����:�3PǸoYY�iI��g�"BZ����+�X�������F�TṂ��	������K3 ̚���E?�+X� �LL��[�����^e��VAZ۷1B�ۙ�MLY�i�R�U��CP�É棡di;�Q6�wr)5˵j�;h��@d��b�]�t�Mx���2��j�A��Ҏ�+X
5v^���+T��K[v؀� �nL�M8�!.P��¦�i������<5��K�^Q�ˀ�N�Z"ۊ�YR�4����ni����߄e�cl�LO=��4jR��c�od�N�j��J�H�
�z�t�XDI�&�KɒR��R�0�Ɇ����xu�n�Cl[I�*"�&ܫ�kZ�!�SW���l)�r�V�#��%m��NA���N`�/Y��bO5��,ҔJv(��v3��5=j�cP�)��ܻ�*
�����F)5���)�X�i�tt�e� �5y hÎ�̢L�Xr�y��a_C�`m�Qb�0I%�SY ���Ū��t-Q6��\NTݥ�Iu�2�֢M;���uƚYZe�ֱyKD�٭f6���T��Գ7�t����3_�X��tc�9�e�B�	]����N�HXg1�l�#�P��`mip8P��W�4od�z��y+#���l����X�V�k
;ѮQx�b�ݭ�(��Za�v�/�r���؃V8��JJf�4t��*^U�t�QM�R(�&��(��V��:�i�k)\F�Z嫥w�+J���6���ue��[M]���(K���jm��S:�n�i�(kM��AQ�^�1x�	"��[������!jEukp:
1&�e�5��jJ�)���fӨU�r�vӹOw�5�uf��aU��"��G7gCc-d�W�E*���,��\R�3���xm��N��̌hs3F�k����B���%Ե��V)��.�B^2�Z�n���ԧ��N����v��>�,PJ��
[k쉛��M�re+���_�5t���k�{�}xr�qc�9^wpm]��y�.c7��i�0Y��y�-Vr���y�iM�%k�X�IdG;��8��h��:|����{�vé��Sr��<��,��
7b�[�Y��H��,-]�/lt��)����p�!�C���m���;���<��ʇ	/\l��	�n����X��W��ɯ�/r�r�M�b�v��]���p�4�<��k�X�d���u�Sr��U�m�]γd[4���U&�Ưe��":vMtg�J��aHm:Pރ�X���MO�Fq:nڵuj�qk^�P�A�]�Q��%6��VF&��n:z��$�g�b����v� �͢���������ӝLe��3��b����>�z:�����-T"�M��yݏ����7A�N�w�����^p�k��al��ة:Biē���7��`�/h�/�+Ѵ6�\N�#��q֗bfeEh̛�7��]̒򓛠+��UwA����ñ��;^pІ	L;��V��Vɤ*�g_�Q�zX;:S8��.�11z�&S��-�U��6�ZL+V����\~s��vY��n>�q_�@�!�5�-��[׽D9�h�9
aN(�3]������4:"��e�뭶r>��T�	879�e�]Y�:�ǹz����,d��%]� �X:;e]�HMo3k��]�W�)l9%�ɽ9�V�i_[�]��X��o	$e0*���+����?��v��=����=?8��N��n��Čp�[	�y��.[��8Ӛ!��K��|�*�e��e�k�;�G)/��w\��bG\����X��yv�*���b�3:q���Eт��jH� @�p`ie-���-���.��쫁�Y�y���^�(]�0b�da��l)TB�Ig$�u��r�/��gsjӾ�f�7�mM�׭���Qξ]�B&Anl�8�p��ɲ�N�>�U����zYt�{m`I>��0�{]c�}���������Pr~���Jok1i��n(�_n5�sN��G����r��#Ṧ�t:su�G�)�6�A��)n:�V�jd�0��!v�%os9��տfe �x�w&�x�p�7*�kF���E��!���:�J嘴�f�2�鴾FR�Z�sc�l�hsZ��SB����fб��Ӏ>����wh�Q������
�֪h�Rb��w$������B8�4x�+o��Y'�6�Fq�M�ܰ	v�f9ji]V�G��չ�K�b#d�i��h�U�o����۾a����q���(b�1a��F �Ge,�]�Y�tZ�ce�w��Bw+�3����:��.�R�e*U�T���u��� V+
��]��؛9���r�}�ү�yQ�r�!t�b�t�\�;�P3����BP��v�W;O8_E��}���t�ra�k#�Ղ�p�!�ݮz5���괼}�j���>E�T�1�%���˷�ğ3�#Sa=�8n�1��9-8�0�T��t��k��m,έY�Ò�u�ޠ�\�೬$momsǘ�@J���{R𬃢G��bs�Qe���/Qt�$u�� ��"�([�׬7��V�}�JF�e7�7����:�r��}�(j�n*_+}b��Ɇj��e���f]:ag��nz\}�JZ,	���e��k�l���5/�?V!�	˦��`��̕�N�����ڔ;(K�� :��}r����|�f�I��t{�"��j������>�K����dw: �ncي6��7̙Y��,f1�AXD�K޾f̫�=��ڶ�*#�:Flc9��ٵ\T���԰�l�1RPp������n,9)���N��k��Z/w�LDgk�bR��߲�6���,�*DB=���.f��cx�į�ԧWR�ͤ:�]̸�����������ZS�	�}n��=�upf��cۏj&��:_D%��r_Z(�ذ���ά�o9>|�m���r��[0��d�C������ʵq�4��{V5��;nQ\uȒ{fv����SY�Z��,�Wwd���5>��;͎����u\ �m�����H�|���w�\�$ܤ�]-Q�o��Bv���R����s�*���C�F�_^��l�Og)��Z�
�6q��Al��S�ζ�p���̤{$c��[F���M��.9Hv��h_<J�tJ�Oz�V���#k��d�ڱ�;��2x��@�zݜŖ���)���6VhH���/^nm9]�����,صl5�n��(``m����Q��[���i�vr�Fevئt��J/��	�0�7ˈ�oH��$��e.�6�F�/��E�E��*޼#�)�؄A�#�6��s�k.tv7`�
z�S�^�q�vK�/a��`���j�/�#�-�6��B���{�)YX��U�ɼ�rw�e�>U��t�Zt��������'0]���eڦ]Β���IKc�����;�|�%���3V.�8���}���(�����za=�3Y&�KC� Dɀ��ΑI_2J�;��n�զD�WK��Q�(T�M5m�V+n�>Ѥ>zì��e;�V��9�k跠Ii�"/���IG��e���:����V+��9��d����(���94���5�.qDƞT���M�ҳ�;�v�J�]�(�}�R��OJ}8��q�
�,-�mkz醺�En�:�-͘P�5����rY;�0_3���B���;�y^���h{��Wk��F���V�,�A��s4]�0j��zs�W_q�����%���N�r�t�.���T�Հ%�pwڨ�O5��#�X�'w��[�����7u�˭��%ԥ�!�����Pj[�dp�m�˴i�x7;�4TU_;A.��AA���� ��VM,��Pe�Dwk�r�_S	ؘ;���wə�9���ڢ2�����kg
+V�ttۥ�p�k|�b[$��-��Z�{���.�Yq�� ������O{�Tj�+�{�HI�j�������~ٝ+�����{`�W2���î�V�*�W=���+m�t��Զ��J̬'�=�k2s��kXX�gS��-��b]5VFG*����0��p���û5�����<Mt"�f�T{p�~�%m���G)��2X����V�@9U��%]g_h�r��l��@DN���ڋ�ԭ�ND��g��lL��U���}A�9��� ��xǕwדz)A�suF-�X.c�ެi:��`�+�;��**�����ʽmv�Wl���9J�֨�/�N�Q�m����tm��xUN�\�.��Ve%r��F۬}�;�T�|CD�͞����TX����g&v��ֹY5zc��š�
��o��z�RJ�OS��Q��Z���|opa���\�v 1�sR�x�;/�.�GN�р1��f�du�lSv�g<��kA5�2%gK��ۥ��9��9���������r	"�uu��ʵHP����}i����@2�^���a�T�\�5��3��%��]��4�$�^���P�tP���.��c� ��F]�Ž�8������a,��ȹצ�ϭ��,"���Ũa��{��L}�`�M<�҆�r颸��֍��S]��D���`�7K&u"{�΢��툳��l�����]��V�E,`Z�@f鮠Aկ+�R�X��+]�JCx40N	�_uv�[��{%Ʋ����=V�lN�{N�S��
P���J0��2��;�)���{�P�]����,�ձC�C0��r��ϻ��c�30�� �� ��;e˗�[���Cw\���g�ud��9FۙH}��TX�S�!��j��;��yX���==�r"�h�ԨTy��.z�:a�RM㾙�z̲�ygN���V\��m�v�_Q����x$�kF��"����]�����;/��m@x�D 00��X(��79�O3I�m�Z�Ph
����ׅ��\�_4�������u�@��.��ך(�JZ��̡��\�Դ���[4q����0&6���B�<�k��X>F>R�S]�BVcW�_rݝ(8�$��4�5�wr�,Nq�N�6���k.���TNpSiR�{w6�M6��e\��EuJ���ҳj��B�փ�c9#�B�וն;+W!�݀�uc*���9{�eZ��xge���ws���=[R٧��$K�J(�vq��������%mA��[ք�8�rTn�cyA�IY�Y����wMGhU���+��r��J��Ҫ�'E]L�!0�9���`����b�/�8�����!u;��%".X5ӕ�]a�Ä:͗��D_׉=���d�R�`�b�S�$eF;�b����2���u��5�;�{X�OYŶ/���4.��(�Uo�u�)�
�n��4R�Xƒ1U������/���ZY:;��U���fY�t����	2�:  k���1�M�#�n6t;U$���Š�<�11,"�=�bl�̣�gP �3(�/o��E�0�κ"�h�ޯ��@�Yg��)m5ʍo�vS���S/�Q��X��rWvz�ޣK~T~�U%���9GB�"[��C�(��M\��B�Q�q�4�j����֝�[��v-ŉ�8��D�.,ý1Zj�2�L V���p7��(l js7Bx������lX40݂{P�����"�[�m&�oj�ٛn\W��l4��F�ڲ���ŉ+�����Z���16���2X�I�p��ܙ8G�����B��no5��pԫś���"Pk��<>�Y]�aw'\�`Py�� Mw\������iz9`�{j�yN�agat�ǯ�[a�� ���Lw Ӹp�-(ʰণ ��f�M�8�;ǁ��+z����o{�6�PU�t�FT��Gj�0D,b�2��qt�/0�3Q�L���b>-���r�07g.߸�Tf�*�H�]�1�6(�=iS��f �vm!��	t`K=�K��S%a�8f�՜����F_b*��WZ2�Z�v����WAR��Ǽ�T+��:��,1���k�y�:�K]�W�7��5k���:$t�����-�0DHʗ$K�Q�M�LrN���[���t����q:�78FA�&��hkx]b(R4����߶";���DB���,9kA�����
���s��&����]@�Ji�/Nj����ے���Hs�(��YjWZ��L��U�x�ǑG�T��y����V-��Ra��;`��.�ۡ` -3�^v�+��I���sr�:ybT����v�tR�^�mM��l辤k��\�4gX��vH]���֪��.�����fͦ��i�,^�2V��|����U��zf�i-��<��t�f)�-��=ԫa�'ۅ
��`}y%n�*d��+��=W�Ӱ��[�v���uf�-��v-SE��K\8�^ ��.��k	���|i<�ț���uִ��r]`�J�Ňӌ�ݮ����u�tZr*��3��WF�۽sR�"�1 ��T�b,iP=e�&��y5"��5��a��^Ŋ䬬�s�g]m��ƕ)�����j4Z���YQ�:__vį�.8t�KOV�*Pb�\z`�P5�i��)�Ƨ>��W'Z8ӟ!Ae��Mpj���I�G�唥:��Va�4���j_���|k�x�J���������X���	dh���P�z��qeα����\7 �d�}q�阢���+1e��9�Y��4m,��A��RQ�M���î��P��m�[�lf�d5���]3#�δ��d7A.��rwP=������qt�-Nk��R���)ވ��S�v���(T���0_,�9�>uf��r;5%U��� ���Uvf��x�WM�iL�x�k��iL�L�&�R����]�On���33s��=���p�tS�owG�v�3;���k$d��o��k��a9^�.�u�PU�M�|ֺ��ۿHn��[��'��M@u���R
̫T���&�mjS	i��	�I�q5[xI^\)6-�PA1ʚ�]�Svú�T�H��C��s�nb����{!F���w�_��{���w���La��/�Ò�9�U�^���|�N�XυA���Ƭ<Ն���2�/��]"{�m���g�q��eMN����&�E�mb����P�-��E2�+�Еu�	��m,LwM���z�nI6g.9��Z x�f;���Bɷ)C�T�˔ᛦ���m�����2�G5ҳ)gc�@i����KI�x�E�>hi�2�=�ػ��\��ѽ�����-�)��D�s�R*��ѱ�5��;��	K'n�1���Q���Iwo�}���n�$:;9NA���/^:_0�u�m�hz�e�7k'<�b�t�TƦ7����^�[����K�9�A�(pQ����u��.��k;��6Y�͎��;�wXu���a��T䢽�b�lD���]2]_uw'��W���6��qⱉ��bJ���]����X������q�t�f����o0.� SŅ]@$�o$SXhp*奓wm�J�ݛ��.+��������+�x2���H���eo���W�ؗI���}��?V/x����_�,Ek��]A�x�WrV�7+�V^��:T�N�|n+�X���H1	Z�
�T�j}5-l
��چoj�j�C�PNo_^����5j� ���Ɍu1�,.�T�Y�gK\b��"�+6WR�%�l��u�aP�]���)�2��{��1��a�r�"-�=�N��V��5���r���!�bR�o��9��B�'�8%3�+zV�ӕ�q�=ΐ��z^oi!�//s:辊P�H��jj*��w]��|[�W��хܩo�4�]��M��|���x���df����sY����c�?�6>=��8_e�Ir��2�|*<��NΡ:�v��D��˻lGK��_}_[mm���km��w�|���y��=|��9��}��>�%�]p��F��r�U���7�L[�u-F�#�7�gU���������cJ��L�^�fEm�} ����u�3�1r�2'�+���Н��奙j�;�
�M�F���a��V�\z�hg�,-�I�WQ%.�+\z/�>j�*!��X�]��f�xv�j5˧Y���6�[ɢ�����Ҏ&�
�|�A��t�.�UV��� k_$N�8�m��4d�),CEV^�U����y��M+ű�V���.���V�����D��dvf��yo-y2=�-��vt�Ms�Q��Aw�G6�nr-]|�ё�Y�;;P"�D"�6^�n�T�+ ����+��y�eX���U�m:n��՛�����Ě��r�4�w�-���p�<�ܕ���>����^ %��w.�:���u��K�A��;�������ênjڻܽo����ɦ�Z���G���8*aԊ����j�ݵB�L���a�.��^�l�=��K�
)�rB<��W�Z�F���.'�P�,'ΛBG1ҽ54Hu�ڏs6��I��y
�Qv�K���7����.��<�Kו�Cӻ ��Ĥ'nP���B�ɮ���yu^
�ù��H�����E;z�R��I����һB�ugT��㙼��JZ��ɵ�:'��WC��V�+�o!����g�T��$ub.���ܔ��}�wU�7nE{���֏�q���C(��������H�Q\�8����g�î�$�	i�Rx�U�Ҹij�oW���{�����͊ۢ��0���aF�Y���U�q�|�.��P�Ei]�����f�-������Ҏ�n�e�T��s�6�ؓ���S駃:�B��D�e�����,\�u��7�Rꃗk2Ռ[ܱk�YĶ�h*Ǜf�pc�t���^�s����C��*�����D��o*��N�u[H�X>� ,���30��dR�&�[��e&�2�[N�P��˃x�M`�K����Ϳ�S�����IUnp�$p;|U���U�$B�]K�;��ٷ��R��4��o�sJ{��v9&:�8Bᦸ@o.._<�s�������ͭ���'�e����8�d�ٝ7�vK��y�2Zl��-F���K�����+�r��Y��j���M���BZEgXz;/U"��"L��CaB���Mv�5�#x=�ط��"�W��S�X���]hk�wcޭ42�>�/��H�� F2T����1}aT�E�%Ыǚ8[ۮ7�9�p�x��2���%�;8+���G�Pb���Ź�˥jf������V�]�nQG �D��B��˦��,n�g�6�Ar�h�t��E���Sf��5h|��u�W;7�&���س�(R&��)͡���+;��RS]�R�3�]��q��pᳺ�"�)�C�*��0���oFL�;{I�oi�)�;!���0�L����+��^�-g�8�Y��x��gA�J��)R�g�Ŏe��;!.�Rͳ��l��� {j�7/F��������|.�#:�U�އ��$��eS�¹V�Qޥ�.���D�9YΣ�c[��l��o9�!r�g���)��;�խ�3���;�\�>���sل́^�7�zm�8�OZPs��;H��*��l�,���̷�"2%X����;�p=�s��Y��u0�M9]�9��j^�T4��mX��6�T�������d��E%�]�\�)��{��1G�r��[d2�*m�St��R��1+;Ϛ��'�+�5E�-��	�;�B�7�����b�`�)C*b�Y�h�[ ��-k7m�
;\�93�E>.�,� �۟q!�����k�/��p[?nuX	��Z����]��b�VT����Ff-�g4��E�Z�TB�]�ڒ��Ɓl@�ðr ��'U��P�|�:�[�p�2��(aYٖ�U�'�7c.�)��[n��=l`�B�:{pTD�`�M ��W˲���6�9)$m������4 ���ӑ_	�S��b���f�
�FQ��Vu���ۛ��X�	j�����q:KEB`1�X��ҙy�^��ln=� +�O�gwI��vG�$�G�3y	/l�.��4�v[/��fXi!�`=Z��קNg--�Y���7S��Zق��]`�x�p�s�n�u:�5c���S��֧`zk��\�rF|{��5w��f�j����r�c�щ���uò� 1��"\Cin٩�K�����;a���D���(ܫ���9���{��f���s��[�$iua˽��R���������:D��4뢾������*:8%겺�-�Qɳw}�w2X�5�@��;2��5��q�["�����q�:�fk����t�'���#���w�Zη1��uu���>;��w�ڏ2��Sv��&P��n�-Z�`�\����#�nT���Wa�c�j�X�W�6�K�
��vk@\���c��Zy�"ݵp��V��� ;HI�'.��T�+�+2�hd�Gp,p����s�Vɥc��J�����)��BP��nun�'e�T�k�\e�)+�V��r���袾�4�c{��W�"����92_������(Nj�.�b_
��Ґ�6��*L	p���R�)���}c1�pZ����]��v�q�O�hb��m#Ed4`��#����̤v(����v�_�����M4�p�\��F���mع����\� ���Δ��`�5��4��E�����@RR��-�c�kO8�(��2C�˶��cV��?9]s�YP����h6ͫ���U�Q�V𤒡a���c��Tߣ�m��]�d��r�iL^�N��Aou�t�Lځa�fĩ����9\�[�hc�mC;�33�o�on��F��t�F�d�w�"*=�(�x"�՝��@
/ ��� 
#J��R�嬖���Bq��4�����H���ٱ+�;}i���g���j����GsX�F���A^����u�b��o9��93n+�PJ���SF�����N�o��k�ù¶��O��qR(�Z�7��f;[�����Zu1��|v6:v�ۗ���V��@���0���LMt�#F0�5M�%;��3O:Nk�$l�|��ޤx�el�\e�z���Cҕ�E�a�*W8��$����(�mb̊�4�N��@�;J�"�ԥw|Q�c%ek1�
�`8{%�k+{�W�5Cj�)���S�Pz.�]��"��yK#h��F�yX���yXݾ�șt�G�]��e�vÚ�˖h�p��\+�szG�S�8�]dn�K3��Z����ֱ̩PJ	K"�u�C
��j��f�����['���nXhi�9o<�m��C��V�4�Ÿr�F&P%��s��)��t������ﻕ�W�ФՃ���h�n�7�݁+�!:�[k;rB*��[�r(���{�ޤF�e�Z�1�>q�C�Ow=kN���W��/��N��A,ժ��c���V����d;!�գ5P��&�+7���͜�7����]c gBWã�鰃K��F웩�*�V�E⼶����l�L��.�H
;����F��)��̻9`�u�uJ�n r�Q�Z(�g��lfe6��U+s
�4¯-e�3X\�x�r9]��۱��Z=o�����:�X<�������H��n�Q\�E��hv8W:����jTYYBZІ1�����Y��WLw���TV���}��]i��;D��՘�5���a�4��w��R�݃0h�B-t
Z�z��F�˪X }i $�����y�
9e���=�mm��M��GL���u�����6�ݩR��	aY�kt��"�]�V�i�	��^�5	z%G��٘��.�7Jި"Ǻ���n�bU�+�B�;��y�;��Rי����c��F~.��u޾���­�R���a�P�<ͮ���p�<ٗ�����n�S�y}�dt��H��;���O���u���Ո^븖<�1��:��Q=L�f���5�����gw>�����%"�osyǺ��hNs��g�u!}�j�hG/�W1�v���-�������~т��nʵw��S.���7�(�V�cl��*C��c%�d��^CEGa#\��(ͽ�:�{K`i yW
P� ��Q^�A��d�NN:$���jWxޗ�i1���EV]�x�d�L�_˕T�'��������[l���=��V��:�F��Q��cCs��A�P�A�r����T�E:���s�%�z�V)TiM�����U��k8Pm�4n�\��	<5r����øȒ�ל��8P�٦�c8�P�Xwq�597��d8��`h�l��X�i���s'����1l�=�n����Q]u��]�u���J�)ZHT��y]u���ES����kp�f�`[���?�]	�&b94�u��:��`�;�[M�Gœx�+䅻�Ḫm�ۡ[R%�4S '%�3�
�� ��e�q���m�v@�	�zw3SDeB��+t�k:�]ZB%.�gr�ݪ��Ƒ�+2�k��ZP�Ѩ�--
�uo����n�ܲ�2�f1�죋�p�f��\�in�V��cr}��oS=B���l5�grc�nc���Z�E��'h�-�ӗ[�%^���+4|5}��A5׹!�8R"��B�D`H�;�`t��"�7k�:�βƾ[�dS($5��\��R�;��Ӊ��yD��G��l};+���Ȼ$�'v�۽�o��utD�I�[j���6$Wrug�X�G�ͩ�u��ܧ�Ct��rp��1�]G�z|I�iKy���U�؍]fh6n�I7r�1�+V�08p�"x��V���44F��hq���������m��`8z!��Ƶ�%�p�L��X��wٷ(R���G��:Ω���J�ೊ��sy���([�vKTW���R�5��h8��wҧcG�A���y]%�z�j�&���/�{X�ѩL.B�Ia� �$wVj��L�yV��[ޚˎ�����%oQܼ-����쬙����̢Uu�ɴԂM
��)�d�#C�_o\ƒ�W�Mj	�W'jϞ�ɢ���S��j�-S��B��f���`�{6htcQ�7�t���j���{�ea�u,{��ԎwY�gP��'���w2'�u��Ul��W͚��)���f\��[ #Vܘڼ���E�b�i�Pd�\��ȓ�����L����"���el��R^�w��{�vK�谹Ѧ���u�^"���8���Zk����m>ؾ�F��-V��v-��MM4{��J�z	b�$�N{s��q6]��:���7�N6hޑ�ʾ�"��4�tR*�k������V*�D��m{F�l�#���\�})U�<��{�H�m�z�`=����-���V���K:vp<�y������e	u�9����X�
�1D3��Q��"|m���Y@�:,P�v�L�+�_ӡ�4QU��ON��^dI�3B���p<�!�`u}�\;O^c�ʴBh1T3���S�����2eh���zC�՘@R�pֻY��[�|������:I�iR�������������SN���f�Kk8J5$@0K�j�u�\�S���xbג
�B=�v�9��,����m;2�vvpj����ŷ&�!�=���(��Y9C�k��n��4���Ոyj���2��2�$Et
F�I.��V�\NrR��+2���6�<.�)�9��!µ"���ު�+n��I6ͮ��«����Wsj��o=����Q0��=�\�vpΌQe$����:�,�m�I$�[�vZ��w��v�:� S���^T�z�0'��.�R��;���s#|K=tK�,��yMg���K������hIy���%YWV�d`w��i��@X�j}�~����c)�oQ��a�n��fz{�E1�+ �0Ɨ�8�&��J�Wz� ���Uػ����t���db������^7pZ��Xә���K6V�[*�V0�a[vQѢp-�4`�D18_U�7J�X�sPCG�[�K�4ӳ�w�Gv���:������ :u�ϸu�ƺ�kl��ƺ��YJm�	���!gvӳ��ǅ���{Z�:7X_k(�4��c�Jq�_h+%��.!���L䶏�(�U!�6Ei�����X��՛�pJ��Al�ae�t�]����A�Bv��_M��Z�
-�ۖ���%=��&{q1:��?Lf`�tХz��ۘ,�&2������Ch.Zu�75���|n�ia%}�Y;�+��N}���w��Ne�B b�.�[r�q<e����u������o,c�0���輤^v��溾ާ�2��>A)%#j��ٹOek_*,d�w�+cVύ����6xL��Qb���`��s�9�hcKC�ӫ��,����(1��׼�.����j�ɚ��`7���7��9'���
�K��o��ݣO�g�f����e�:�h��kV���Uk���M��Z�v����R��`]�w����g�&ʁ� R=�� ��F�����)R�T-����fN�5��)�]n���4�Pi�/aF���CU�zjwWS���:��.��[8�=n��b�D8��0]^�٢����Ya�vs�;Ip�Є�b�}rry�ҵs.��w��:���A���Y���m��u5�AYc���J�Őnڢ8n�]�B�X]oQ-�[e��#sv�y�<	ՠ����>"�u2�r��]k7�7�g>�k��x��c�-�mR��k�͔Uȅ�gV����ExˌҼ��r�vee���T͛�Y���w2k�_*���N��hM�zjU��eNa���o	�	l��@jˮ� ԥt�Q�+4�J����*�PV�p,�ЄjSOL�on�r��  #��z>'*s����~��諭���j�yŴ.����U�:·�~z�f�N��O�ϟ�'�x%�"��kSÒ�&�GCz�;��޶�\�^7Y =���`����W��C6
?�^E��R\�e���:e�oH�D3���pq��bY�[���G3��`ܾ�=�K'ù�	^�����mG`�6kvp��*L�9�_l2�1sܗ������Au����+�Z�ۮ��}�֞�>·�w�*,�
�I�)�
3b��qu��o���mj�ߎ���-�Fջm��?Dfv=Y���%��v-&�4�s�m_n^�{٣�lI�&e)�:Ɔ�ͱ��ڴk4P�R;Řs�;�hѡ[8B\U�GXX!��N�,2�Y�F(��I��a	��˘>W�2�C!�c�Q�h�k�UE%�z@�|��r�iQ�˘�0S�d��]��,��u�uɂ+�=����{�p��L6c;�z���K-f�x��Sq���O�s��;������-�-�#���	79F��"g"�C#B�|^]<�8^^ԮD_Y�͕4MaS�%l!�����a��dë23+]�Z���W`iJk���X}g3:���'l�>{]�i:r�Ġ	C��9b���sƷ@Y��U����pBҚ��M=W'Dں��wX��$��u���t����FA��8�C1J�b�7�:�.�V��N�X��V�4[��뢹�Ϝ�Gs��h}#�;��+��]��\m\�(ۍ�q��qn4Q���-�H�!���8�j-�䱌j
�� ����dh�`(�)ci�\S"ɨ�3i
#E8�G�B75&�H��LѣD�1��!�s���s�Y�Hi6"��&J*0F4A��ŷ�E��\"��"M�����h�Qis�\$�8�h��H����\b�Q���A2��h��65���E�#@F���q�)�\!EE�$�P��-�CI�,l�(D��bI�"Y233��`�dL؍��HĜk�����bn7�4IDS"�1!�ڽ��������Vv�iA��7�Лi�y�`���ݚ�r�S����WDd�a��gw-5����đ
f-�*)6���
hqp9tn��UfF7�.���2=Z
5�2UYu���]g���
����XQО��v	������S3іlO &%�c5�_p�h�ʞx��a�2��`|@�:vI��EW�����Ɓ׏48���Z���B@à�~�6o�S�r�W����EVd�`Ws�d��ݢ7������8��ɸ|��^C�_�h���i�\<*��;1gֹ��6oF���**�/����el�18:噳'��A��5��I��y�qt6Q�Xݳ�;+F˜���L�ُ�gC�"#��p�w�������û�v��b����7�P�`U��Y�=�������Cb��<�� /��޸>�i� �.J��4z~t�ݽ݉Ұ�x��!�/�D3��Yբ_�q?mQ�me9���#.92�[�/p��ɥ%m!��k4���������l �'���L��Y�~ʤ!�[P����fC\��畽%OWe��/n�	Dl�!|"�k��e����y��&�|��2Z�o����z�M�GF�|��.v����fd�-A{�3hF�;���쎻Sݐ���[�L���N.�՚oN0E�\lt���3M'�i���O;dE}�U�ŝ����wg���wy�3��*�f��b�j� �Q)�M�z�a���h�ݝr�F��N��ρ�hd�bP���9O?��b��G�ώ 3d+�Z��.��s!c�r*À#�@2�Vt.�1V��Ԗ�?}5�5��;��� v:?.;SC%��+o�#��ƃ���؋�ݬ GK&�q�����R&��	s`��-��<��:�Tˇ�#"X��	
���n�x2 Hn����ɤb��LE�a���s�K�i��GA���
��"���Q�p�L����.����@W!o���e�z���VP_<{p��c���ʙ�M��T	�"�F��`J�����)��V��s���ƀ=�_��.T��u��U�KRj���N��&:sj�fU�J�t{�Ȝ=���+���S�>�r�Vh9?1ATZj��kO�&�$N�^DuC��^��z���uﳟ��[z���x8 ��^���K����.jj֭��*S}�_t�f���g��4O��ۅ������FM�Lm�*fn0Z�B��Zʣ�Ѵv����%����2�xV��幟?}�0>b�����y�}G:
K#��zo�X��j��z�#Y=��po�I��7A������	��pm�uQ%���(�>7Oq+{؁/3�z��}��ם�u�X�� c��<fb�}yt�v��z��Q����O>v��<NV�}zR�Q����EQ�vs���@���S�W4)�|bδV�P�hѭ��`�.�:�ꄮ�z��0�d�)��4����j�~���,֑�)ߴp�.Vt��:����ZY�Z]�65�kQ��癦xD����e�8�xH�Rc}���C�	tn��v3���:��KD�au�b<+�0'��o]�uf�t��u�ʌ�l|����1@ݨ=�zi��@���r�;�..�k|�U�{P0U8�ɛ��!ʿ�a0��r�/��n����3�v�pծ�̎��M�3�e��ݢ�㪯�C�2j�������1��Z���(����&���B�K�9�\�sYi�R��n6I�t�w 85//�ø�..���G��wOڱ!e'.O>��,���X�gai�W��1���e�jS���w�`��4P������� ��q�ީ�Y�6�5`p�rf!�`�1�q	���͉�F���B�#�A�7��f���#�e�]��/�*{)�.����_'�*�Yn� h$7��]Y�1�(�m\N�ӄ��+�����q~���!Dj0��
�2����1XT�S��&=�dڮt� bx��Ŭ����% �ݠn鮏f��u=;��2.-��j0]�p�o2�r'+6G|���{ ���E�9�O����} ��/ˡ��J<�/{�x��^ab�L��a����2�ڧ;�$�''����冁�%�p�[�_[�?:��g�y?���	��&�w��5��E�hcY:�����1���@.�GM:'�\*�1��6���uF���Y��#kD���*e>C1]_Po�#��O	�+l`��p��t=Hׄ�TV�L<?jLnR�oi��p^L��{�v�!u���^����!�����D������������C.�{�9x�x�O�l�.����Ӯ�s=���[��H��x:X�sDt��AL>��8uHk��;D�;	ʘ������#gg��~���dj�12[��:�d�OOOds�HCp9��(�Kp��z�-�VC���uQ�_����A�^��1JncF���l�n^nl��A��S�/PC3����Ҟ�#�J�T+�_V��Dr	m�&}d�DuR< �}0y��ZsU��Ȉ�}}=2��g��4+'܀Z�+ �)�<|�T;ǧ*`��*�9�׵1��<������7ԛw�*�͢S<I"��Ӣ9}�Vo����ob���yD�`hucf}/{{���7�R��Q�����{��i:��<F�̩�X�ܝX6�G-*�Z��������׋)"�[��۾�d�3��]�ݍedj�QwE��R�����.�}�c�x���ؗ��*8�͏сǅݴ�1��e�Z�q���'�-[�C����I��5*�����ME�S�,۰����(Tc R�TMݕ���ƀ0���9&۔^��Xs�t����!�@�gﰘ��T#�����<�sK=$[=��������; ���;��0�U�x�=&U�)�r;[;2������k�"����d�E��B�f�=�]$au<*���Xi�鞸S��I�>��X=k����F�s�E�Z`V��X_��a��
�xm����9l�s�x{������6��o�I���d�ؘO��4BBe�����dP�:r9���S�/�q���X�����v�s9��0��T���g�GF>�����ϘˬM��{M3k�������_z�ٍ%�N�j���d�����n/:��톝Ҫ�e��f�5�3�Q����бpw٫3��UayyՇP�
�a����1�������A~�!��ңt*С��w�A��7�l��1ڹ��-�ޕ�9��<x�o�IflU5�X����EP�ǵf��)��:��H���k���^�G+W�d�;N�.r�%j��8J�:�rc@�"�M��{m@t»�T$u��߳���7�����Q�yuC����`����o�6+�T��b���^G���L`S�w�nk鮘�r�T-�Ԕ�g�
���оO�r��3����>3��s�eb0��v��ę�w�R��a݂A]m�(z{:ݿ���xh9��J�'�x'���{��R��olG`u��&�0�&�kێ��x�5bi�=*�KX���9xWu/���%��<���Zᢝu����?8��3�J��t�W��g��1����TƤJ7m��=jsfv��X���6��9��E�o{]�~�y|�1 �u8)�ǐ�I�C �\��/_
)v�-z>�+�G�	s���Z'��@T��`u�c�M�'}��R&)T����R�H� bT��j�o��0�D�b!!W�sam��I�9���QJ�G]�XGf�����V����L�u{��(r�e%Å3G���,��ctT̫����-V�J��"s��{�u��_#��>�a�?�j��ʮ�r�|)�<����/������:�#ܘ(Clcu��M9t72�Í��uU��|��L��u�(һ�ʕ�)1ȳ��B�
��*�Ƒ��a�-_�Mը	�n�����t��j�V������GU�Z�U������ʗ
W��V���egS���U�x	)jG
Y���6��"���i;��{Y���:r҉C��pc�C�:U����n�AN�|+��y/o (0#��_p���^�ıp�{��<#���:���-�����n.�L���G�>�0[Y2���?WI7�<$e�˒�*'mCP�[20�[�F��+`� �6߇���b3�> hT;��k:pU��ֱ�m�����~遂j�:k� �3��YJ���·��!�<��n�� ������2���y�[a�DXlF�?��<M�-䭕k��ڈ�.^هo4�D�}7�j�z6�Kk��ACw���5��پ4'0U�&�t�5x�Fq�r��jP��of�*����O����ڙr;Lt���׼���pA*��H6���g�.�{]-ӵ��랩�
���5�^��y]qr�Ӕ���&�����Z ����t�1|�C��nJw-�sظ�L:�������r�b�&T�#��I�����;Wy��ZS+�y]��m���y*á,F�*�f#_E|�E%|�	��c���q�5�}�+;uV�~�_7��0�w��i91렀�Cz���K��𮏋:F ������]�-����-N�Y9�Ӵ���f�y��$�G����f�<Gnv���滵sŴ(#K.h8n�x/)W�1Ž�2��4�j0�O��f��rv��]����h\ќ:}bҫ��B.�}Q)�pipz��!�Й�d��Q靬ĕ��q�����13	.��:lB{��(;�;**AQ�����	���[�x��cg���^�b�@�	�l�OBt4#�<"meڰ�_`�ok+*x���":�Hs|}Y� tFI��U� ��9}��O`r��Yj�C_&LU�,�A#�nޔ&ae�2������qq4��Aߗ�e�OZ�!X��'V�C�r���2�:�ӉY��pB�?6t[�b���ur�����^b�^S_���t/����Llond��l����˵��s&�ͻ���X ���s��&�������^\&.k���+�X��@�-�d�޻�8du�l�d�x�]`>�B�5NV!��y񬽨�裴��9/��1&p�=�q�n3j�3����x�@�����Žj?�Y�����CyZ��C�xE���^ft�
�>������.��O�*]�#�ڜ��6���@V79�aƫo�����zS��[��R*m�ې�Ҩ�-3��,z�P���Ab�zºǸ�$/v��o[�to�7o��][��Wc)J:��sN���~���ֹڟU�G.��jK&�,�D����t��8�ڞ�V�&Lcv�FE�*�mK��h��ՓjsX��{��-��|�kt�j
ƕw��k<D����I�O�WX�1���5����t��|�٦��_4���=�����KI�)?�g�u�Tr���`'��hp����(֒v���������?��C�Ю�rk+ �(� ��
C�{����a�K
�MnM�9� �����N��
w�
yOOu=�pF����1.b��\��~��
Hj�ŵ=G��
�Z#VО���p�)Ȇ�Zc"u�ٿ��0��:
O�Aw%Vf���:ז��������`���[NQ}��y���0A���Q�o7��"±��By��$v�1� �*,l�+��JYM�Ð�Ls=#��=#��t�؆�wUv�q�̊�!Tp�'�䤀�3����x̬5���Z�ђ'��o*,U
yؕf3�yx*l
�xX_��0���k�m�W�1˱=Aw�6V�`�ҦU��Q���;�M��d�V:n��r��/��qB5�k�V�uwZWY�(`d�OF��*��0[�`��)���79�n�%6��ڌ���T͵��7��1_
�׶��;`N�l]oQz�T^ӝ�]rqr9$��b����ì��2���Xs������:�7��>�6ᘹ����y��`�j�_M��k�t�-¼+��Kwz�+)�d�R�e����Ŏ����Uq�JYo3>h@B;�������5��0U�#~��S�l��p�CV�s{)�+H�,C��񬛘uW��S�c�Y��^厰V�8ezӼ��8�n�����$�SeT��s��c>F�Y�\.���P����|���3=4�	K)�N�3����1���i�o}|Z�� �����g��Ϻ�o�(��V]����GQd}�����k��U�>�I����&����}1a�=;;���7>K��R��w�}_�R�� 2U��<\��w%\OTsI�#xz�/
�/|�`��z�ѷX�A�@��ڙ:�y:{%�d�����V��d��U\�!���Lw*:m�W;];- ���
�ï�8Mahf�q�e̸�M�����u-���J��N1�w/|���":ch��t�x�iǼ�77�m�3�7�@�&�an."b���f��M�H��L����*j^�Rܬ�xO�<��U�A�,�V5��pWʻy��c�c}��Z<3l���k�i�
^	(����Z���Ep��ͩ���7��ؽ_N��Y������w��tPd�*nl��jr(w�n>j�O����:rc��E�s���{K@ctc��]�믥h*���,C�Z�����>�B.�7�B7�y������J�ɂ��m�³�L+�ˮ:hX�E#"�U�M]���嗴"@�CK�ۡ����޽���6�j�vN-w'*\���Y�vmڜP��s�f>O�E��s�;Em.�HQ�"���4*��3u�7��׬'YǸ��1��}sOf�}m�����ӀJGe��<���ZH���)�c��ɦv\�N�cbZ�H�y��WsH�\[B��t�U�� Dv�8d==%��.��j��o�P�k/����p�@Fc�n����r�Ȁ�ӛw���l�͚��o%��"#t�koQR�o<C����/���!W}�F=��]�{ܹn\2��e*-���o��Q;As�9��I�|2��*p��Z�shjKl����Ԗ�m����s�Q����<�ڝ.���Wrܛ:*&�Z�xX��0M;l�d�ݴ�Psγ�����qq4�f\wF��ʟ�7�f,p�|C��.�
V���j����A0c9,�(����{�z��k��#w�P!c��;��nL.�iL���m�˕6E���9�Q.�Z, W ����^we*�do
�>J���S4q�B��j�ff�g_/-B�i�΃��u>w���;w{-�j�i�p�ҚXѕu�!Cum�²cn��� �����v��O����Y�g��5���]� 1����t�����k�+S�68^aܩ�F�շ��@W5�<�wfK��>\ӃO$�����Y��Ȩ�Q{u(�Nܻ��]�ĝn������D:�b:d2��w5����ؒ�
=�o7�L�/��B�c��,�q�����r�sxE��_'k��2.��������[����u�����	����L%u��Q��
N��`F���hoe�@?�h؈q�򠎩�0����H�8�(��1s���f���aAh���o��hSoM�D%�y 5z����5�n�(��$xdn���Q���G_n�Cd`	b�vk�T{@[��%�B�[�)�gS��;Gq9���N�\e;,Ś ��z��GN1͏2�9җFV#o��t���;K�+C�؃�}a�k̓w2!�3: ��G���m�9Y+s�F�6i
'��k�f�ǴhW3�-����Rڑ7.LS-5��6�4�%
9��:V&�����7�Ȯ�ś�ms��j%�Q��zԫ}]�G%O�퇻�8���`к���x,
o�,�hL��|�L���KT��[H��v�Hl8���㹩N��<z;)̅U�%dX�� �B����u�ͭ^���)��7�*w�W>�e��Y�7�p��!R:�x��]_�޻��_:����i1�!����$}\P(��&f7ĊI4��J""Y'9��9���E#EC���$�&21pd�@i�D����DJA8�JK&�9˙7*"����24�H�&�,J�9*LZ&X�a0���FE�p)0�i�\bhXc�C3��dʜ�%LR��&B�@�b���" ̆��LI$DH�J��F��b�Ė���$�X&LJS$F��JA�,a!0$���ɦ$ʉ�d2�`l��3 �M&`L�D�&D�#PFDP����\���n��������ފ;|Ⱦ�$0���]6�MA�9Ҍ���η��Wn�����
aFXN���q�a�%��Vj;dgi=w���ӽW���h���>�)>z��ޖ���l���t�{�WO�+����r��Z��Z=]r�ߕ�x��t���n�}k�򿿯�W���k���C}[��\_;����{x�mҾ�;�����\�!}�����xUh��T� }��η��7�nz�z�ƯM�n7���]�󷵣x���t���з���x�]?�\��v�����<W�����[���x��|_�κ���ܓ�{����̟v��2+=��;��������:�(ߞ-�o������qt�����^���7p{�請[�q���]��<�}]���]�v�����OU�Xۥ�W?sz����F��+���gꝟ�ݟ0�-We�����9������7�����}�7�|t���zߺ�zZz����o��W��z���*��W�mt������M��o��v��J������[�r�7}s�����_y{��zU��79[x����t��-��w��0|��_7��1}m��jw����v�k�|O�ۥ~[��}���]-�^��uz��v�ݭ~�Ioύ�y�6����^u��zn��t����o�ں^+⺘�|�r�G	�=���船�����k��/J��~W�������}^��}[����"�W�nu�+��5��+�Ϳ_|���Κ�W�����鮟�֍���[v���з����=W����yC��%н�)ꓗ��w�Q�ѳ�N�t�ǯ\�qt׶��W�w�t�+�t���w������W�����7�+���mҽ|�~]��\];W���x�5ƹ���}�*�ߕ����@�~�E1T�X��&"��f�~߿k��������\���zۦ�5���w�+��=��Wj���K|^����h�-�����}�zZ����]���-���t���_���d�C���~�K��yq�U���Vy瞝~��n���]+��:�cx�>r�?_�u��_u}�|[�^��}�����mƽ_y�]��:qqoǦߗO��v���{��|��h�[������O�?D^��s��Ǡ�L��^��R[���?y�Z�x��|������ߚ�t��u�7��]/���~祠��q}�y��}W��ҹ��Z�o�q���=����/��{�x����:����K}W����ל���������x�;�}Q[�v
�M�:�a%3?n��xV�{�-{��^��0;�V6�Gpv��V��MP�9�ܦ����l�%n��Wa�[ۮ��G�M���t�E�Fl��=ef
-�*�a�|uc��r��vr�w��S�V�=%X�������g{��}��_�s���|W��.��_�]�ﾾ�x���7C|o��h����;�/m~k��{��ץx�˥�o���:�Q���W�߾w~W��owϽn������s�Ƹ�}}[���{����<�����\﯇������n*�n>/.���Q^�����w�k���ͼk��z[|o��u�k}^����m�m��k�m����yﭯ����}_oku߿��?��s�r������^z����O�{n��]-�9�t��q]�叭�����vݪ�q��z���n���]/w�*�^-�9�?��^�������_��W���]6��6�z�|�q]����[�޽��_;�|�����>>�sU��C�V}�)�����c|#\W���羶��]��ߜ��o���n�]-%�?/W|-5quw���7ֺ]+���t�[������[�F����=�~W�{Z?<����}����~��]��;���?�����S }b�#��?I^-�����u{[��-�߽wk��+���~���^uk�x��9]7��^���}m��x������/�����MzWM�_M~o�~{�������C�:#��~�_P!U��+�n*�PZ+���]���^/�o��7O�qF��n��߻��[�\^����񷵻W�ߟ�ץҮ-��s�Mq�<�.��|źU�����5�7m��_|�߇Ώ�ʋKV˿`����Ul������� W�+�9��t����^��_�+��_���hޕι|t���]5}���گ��}W�����o��x���zU��o=���zk뵺W<��k�}[�9���s���>v���篞��=����WkG���}�r�[�]��m��ێ5�]/���o�z�b�+��_|����j�}[����o_�v�y�]�6��[��]-�DG�y���1�L��F]���W��qx�&3�|���緟U�v���].���WM�}WK�{���h�����]-?���+�^��n7���Z�zW����]-ⸯj眹�-qo����_�w�5t���1���71���t�xx�Ժ���Q�m��zoߺ��n�ţ��u�˥鯭q�{��ݫ򾮚�������o����|_��h�o|���_j�[����\Q��W�9zU�qm���A������1~��F�h�e�ԃ��)̡̈�<Ye��o8��޸�޿د�a_vؗ�9�WA睼�q�B�Z���y�*SӢ�`<�w[�`ԷL�c�ҹ�%�+��˘��v�'��ݦ�J�bj)_3���d��l�M�W5SY-�<��?ԯ��;Uſ_��w^��\y��]y�竊��~\]{�nѸۊ���]u;�C_��+��W>so��u��ڸ��~t��ܯ����o����K~��鷿����1�LBz^�Ҍ���u�:�j�=5����Ͻ_�{U�q���.۶�~[��_�}u�|[����ս����y��z�zW��[���F�\omt�[�q}m�ӮsQoǦ���z����9�ٓ,�S�3j�I��ּ=��}�����mϜ��m����Uv5%w^��{x�֏�y���/�}k�ח����q�+��=�_��W����ץڿ�үyu���]
�[��L	�S	Ɋ����c�S��o�v�����x�+���+�\�Qo������nz��WO{�����|~v��9n���\W���;��~W^�ߺ�ok��_Z����v���t׭���{���oJ�|x�"�
�T�}C������w��M�C�_~����n+�����wͺ��qF�~{��E^.-�w{����m�ߕ��k��W���5���׻矻��{[����yק��F�n=^�u�����}n����V�o�s�6��ߎ{�|�w��Q�6�΅�{잟��)�=��^L}sb����n:[�9]5��k���ž=w����U�u�9_^��W�������צ���?+��=+��o��}O9oJ���gsZ1�������T���t^�Þ��7�p�n,����J�{虊����'��U�o���ۯ��j-�\o?w�K��W���ջq�yv���<�v�v���w���ޖ�Ɗ��WM�_o>{���o������u��d�����cs�tފ������&fc�uu|k���߾r�}W�t7�yz���W��}[�w~w}m�o�u����j-����۝��:WŸ�k���z�]7����޹xޅ�+��̮���^7K��^��}�
b����=_��w��_WK�\ߛ���o�˜�7j�x��{���wBߛ���+��߻�ۍqF��������ž[��Wk���-�{�˦�nq�\׊�>�<�ͻ4�40<.����v��DT���[�q{]>6�7�{�k~W>�^5���*�n�ϼ�y��5q]���u~{[���i�η���r�_��:��o�ƻ����h�s���J���S`e��W�j�%�靁.3�xቄ��̸����l霁����[��ȭ�Ss\��映Zr����y�^��_-�g){b�ռ��;�wL��xҡ�ɵ��;��.;7ה�f2�p��6����dxj�C[;3�
��Qu��Z�\W����&����n�"�z����_=���Ͻ������n������h7������-�]*�]r��xۯ���q���m�����έ�o����߿w��E�n~�x�}j�����v��x�U����>�鯼<���/N�����r���[�M�;߾"�� ��(~���:oKG��9�J��+����|��Ѿ����/K�t����u�|k���{�sn�+�]�����W���׻��zx�m��+��sx�~�Ƣ�w�߿�?]u[����pl���@��~�P鏼�[ھ-��^=�y���Ѻm����7c}m�\k�x����_+�n�j�W�׾k�qt�o�^u_[Ҿ/J�w�k�o��|_�}���x�wҀ.��� _���%s��"c혈sw�?y��^���n��\��u�\k��oW��o��\}�^s����^���W�9_�n�q��똷�s�6��u�Ƣ�+�9{_�w�-q_^����˵����y�%��=�*h�֍Yp��s�Lo����������m�q�y�X�֏mz�}����k�]*�^~��n7�ź]��޽���oz�}۝r�+����t��mל��]s�_����s�a1�0�7ўQQ|�w~Yy�l�CΏ�v�j-���گ������|��x�[u�.׿����۟��W��?��h6�o>�w-��t��~�׍^������������n���:�K�+�^���	������\s\�����]��5bo��{����v�C~��v���/}r���ۥ�7���K���9�w_���}���j��Lg:��ܳ75'=�:ŧτ��+�s���R������G��*��f��^ʘ�j}�D���zu�<�-�s�k)gK�'���O-����n��0������R�s�yG��q���}wx��W[t�ꞥ;]�4U�>��u�9-[���߷�p@�يpm�/��F0W�Z=��/$�a3��Y�uʌ��ɱ�;E�'f����7u���e]IR��H��DF1ۡ�?���J��p\�u��dU�Y����+�`{�7�L��wt���C(Pd�󺕱o��`w�7ǳ��H+zf((P�ۇ�9|�0.��;P�9�	�_�/��w9�B�)�1�ӷ�<4K���ڃ���>����ӗi�.9�S�~[P�?W;2�\�9:L$6Tt��WT5FT�pp�	Fv���)�{ͦ��V��L��n�gG���m�~fz�9�k�Apr�t+L�Ն1���a�A[}8-��❋��:S�a�5�Iuv�Ƿ>ע�>��R�W���  g%��kg�`�y��Yn�&y�YY9c�$6 �H��}b,�Y�y�d���J�B�l���p�Y��{x�m�a����4�M�y�J���X��w�0�c��;���yd���C:C���V��Z.�1mG`��zh������p�L�����]I��W���{��H|7F@�_�ɋ�>�=���b���?'���y� Y�� w���n���DY�ב|��0W���m���x^P��'ܺ%W7���,|صte����r��upg0j�~�wW`Ȏq�5�&�U��Ϊ/F��
^�X\1AT&�@�i���톱,`��~�N«~��4�/��X�ɸND53ҍNI�X3lZ)j�[{�rx��3%H)�``���=%f15]3*�m��(�hj��2ն9ou).!L��o��cA�7�{���
P����U�h>�כ�w��<Ӕ���;@G ���J����{��"�t��~��ąr�S�;�v� �����I�S��`��L��}�[�}]6�p�{fy��5�g@����ߴ�W�Hw���j$�������<�=�-=��t��M�%P���bt[EM���hR��:�Z�A�A��d^x��N��ͪp*�֗{x	K���������6��t�=0 ��v+�(N�r���c��Ħ9�e����1̣�f�� �5��y2��i��sg�禎�<�8�.�9M���}�6|���S~��D���5������~c�SC2�|(���0�pU��_I˗��ν�~Ǟ?:���_
�:�|9��l`�*�	�*���Nrzf��1�\J�i<��<���W�%��F_Z�a�Y9i�5Y�����,�e�h�R9)[� ��#q��V�J{����s�7�O\��h���w 85uN��Ht��uH7M_R�<Q�:�೵��6`!pGp��;��	�C2��D'y�C��h���냩�Q6b�ߵZ�7/M�[r��ѵK��e��Fم�f��*�r��������U�i��X�=[:*!9`���XS�]�.pv�w���c�;�*��wj�"#x-�N���yd�=i��+V�pj��'	��8�����n�ξ%cۧ�7��E�	 �tn�� �l����#~��lwqҧV�X͉�Wj�A;�Rp7�91����ʕ]��	U���a��]e��槃�n�H#�Q�Q�4-�<񭵺���/}��$�q��ו����t���ᙃ_�HS{�x�ް.c�v�-��{E�-p��K`>��x-�����V�>��x5��k��v�'=��=!���~��Q�V\7u�6�<4�R:h/��y��^?p�]gD�ķ�w�N3��������K���pڈ���0Ԛ�7�#�����k�U�(HW���t+Rŷ����Wz�+��mDQ��<N�'S��vb�ﭫ:<M@�T�/RͼW}��O_^^x.Zb����ϯ��)���Vt�1�衲9�h������R�����A}�]9�,�W��1^�.���G�W��X�NP�7�*��u<3���L�n�
�a+�>�����EJF��.�ys՞ɣw�����jiWx��Qb�b�w�4�E/`솢J�X@L3�)Z�oՂܽ-5����eG�n3�d���	��s/^�hck�b��:�@]m���B��NovQ��O�`6��2Ŏh���;�_Q���Ĺ�Pg0���(e��bpQ����MC��{
�,�9���v��>��/sz<y�U��j�r-�3�_�6���ښ긠�*?U���"#�Q��y=N['}�:�=Rv�����o�m����)u��/�̊�\�Z�]
f�u��AU7�v6˥hGL8!��"�p�O�8N�vaOh/iL\5x���,����u�5-��G��x�������0���Bq���F�=ܴ3I��dC����Ɍ���v�]AfC����[�5���x�C��R��=l8��C�am�G�h�/��P�)����T�[�~� ��W�w`�k6�P�#[>����*�:����Y�Oi��p�,�|P
n)��;	��f4��0{b÷0�rv�U��`�P�6 �9*���W��x��xf$�{�"�=���y�t<�
a�[7�Z�,d5�h� �޳}~hPtk�m�W�1��<�)ry��a��7Χ�p����QP�$��c�s-&���@
��t�r��l�F�p��'�GͶ����W��g
���P��R��~h@�X�[�a�5D�2ys{�y@����c̴�p}�� ���2oqs9vl�:�uSS]���֠-�o%95r�k8�G��Yu;�i��Vo9$�]�^LQ�s(�+��l�zg*�h8����6�኷4�m��K�i,�� T!1���w��S?}_WՓf�7vS��6���!��r���FMLf%�SW��{��厸Vw��<���uΕ�@{�`�%=V�s6�Mkb���F�[V냇�xO��f��^v������|B�T�y�}�1C��v3v��e��bm��b=g�uM����O<�R< �~�u��
|�kh������kG��J�Xb��f+���;�5�C�t�<!Ć�u_IU���Lsr����K_�ut��b0�re�Ϸʼ7.��^�\0g�ZsqiQ<4�PjF���f�@���߫��q���!�h���k�+"B���vHo:�7� �뀂��T�q��ƻ��Jg_-��`�U(��ix�w#*֎��R�L��@˙�9���-+g�;ȳ u>ᙩZ�}�8���5�T0eL�U:)�,�anG%�b˭�����n��W�N�َ�Y�G�7]"u�{����	�)+��9���GK%i�қ�:�w##i�j�v��K�Yo�'��	�D`cϒ���u�<kWq�z�g��y�F�yj�Z��7v���7MU��U�F�k�����c�$��eRʝb��30��Fق��4�����kp��E:ͱ=dQ�7m��b�P��y���G+g�d{���cv�y��ߜ��[�W3Bs��wN�2�z�#�G�T�WJ]���������{[��"������/�y&:u읾��:��C�(r�e%�E:4xy�嘒�hӑʿx]�HhU����J�|����r�(:򽹞O.�ו i[�mh�L[�����ono#M��R���%Lqv:�7'�h?!`A���]fW��!+�:����kh����2�5ډ��j=���y�n�e[����X�&��,�� *��Su�\�OO�Z�zsx%�^��x�r��>�ȁ��3X����t����v3r���WJgy]B�a���_�hn�ߩM�����w<(X��3����k3�a�q�>���De7����W;��^^���}P�B��f'C��S�ʄ����2 R|س�y\��y֠�u�s�~�+|������je�pACu;�g�%��NW��[fGd[��W�Νk
���e�<�uQ;9*��U)g1ƥ�~��s.A�)0�d��G��[�vׇ��KT�þ���t��A[��PK�_ơʒ']zo�eu��1���������xy�h�x=�g+$�s{��Wv�e��C�gn��T�ۖL]F;4q�ͫ/sq'�Q�f���es��J��b��']�A2��2�wGw���g6R�R�9��3�`n��~r�ݒ���Z���	�*K�-���e��Ph#��>�	�-�k�aQe���H�Z3���Ǝ��̳�p,V��%����c���O��8��~�"��';�F�3��,�f���D]�1G�DWҞs9�[�N|�z�mM����$�բ�j{h!.�8��op4]pp�{�J�P�j���Rd�ș�TϷ7vwD[mKR�r��Ϊ��s͕��ߗ�m;$5]mY�h1Q��;3��BE�<
��8�U� ��3Zp}U����b�Sn�����(rϷ�v���/��I���R��	��ܮ�K��;n�.e��[��-=:�*X}!���qɊ��k�.�Z��wV��a
����z� ��귯��T�&��GZ�k���/xN��N�T;ʨZ7�U�U��]�'f���.r�JÌ,|tcЅӶ��u��";���vH��f���Z��a�;�HN]�7Np"�����㳙��+�lpycEDIg�e�j�/z�Z��Cu���k������5�i��]��6����!V�
ĥ|.�X7�Ҵ0ގr�#����;����]�1��n[�W�1���tj�f��E�yǾ�Mu��9[ښ�[� �vM|���2�a�x����&��9,�O��[N��g�B;�@Dk`��}*U��f��5�@�i�Iz c+1�s�	�H��8]F�6�H��p�C5��8��櫷׹$Ʀ����էDΗJ�Zq2�|n�W����N,�Ĕ��U���Z���A�ai���+@=�]M����oeKOj֒��-6�ʗuư��gl���i��7&��b+{��dEٶ�[l��ߘC��:�(�0����4���;��v�xO��]��9z�)):�ww&#o�)Y	.�ڦ�D]�k�.K�2��o;F��fᲮ+z���}�2(A��'�x�ܹ���i��s��7-�Ǉ����[Y��[�h�k�[a���2����ԫ"� ]_��'@p����z�����jT�&guf�k��,��wI��hl��(��g��B��$�78I.���CԲ�����V:��0�����+C��X�$sB8�MY'� wW+'m񺊻 ��wC]`s�T�Ta����5�Î��R���v��ӮCmQ�F��uC��WvSJ���КX�7)��
��,������5��s�pS*�� �ܑԂ��< Ck:Wv��jG����V��E6��ԠXt�v�*;]�@]l�� ��f�s.�ۛ��qid<�-��*,ܸk�u�7JC-Vq��˺�k�p#6N<�8��Ω�t��wI�,t:���������;w�+_=_��w��\����6!��YD���ĂP�4T����B��@H��D��$�`I�D�d҅!FJM1M�00�ѢJJ�D��1a0
"
%224�D��f$���&�&�`��4&�i L�d4!0������c�f��� B1L�(Q&�b#"���"1	�&RA"��F� ���RB&bPA��1� ��6&cSC1�RP F�A�h�aS()��F1IR���L$�e(# Q��Ř��`�(� �F�ha3�� � ��9t2�,�F�Cy��o-+Wr� �|�ȺrM�Ʒ}&S��R��Y��(4+�{�g���y$<n����fJ�w}�W�W�)G�N���o��)Ʈ}��q�]ШW��K��u�0���4)��T`�s�u��(����Gh����]mϘs�
���@2���S��}ם� T���D�X��d}nbg	�"s��0c럌���>����N{u��OD6n�UJ�D�W l��.�Ⱦ3y��rv��
�����5=��J�Hkt&2��J��7Ht�L����=�9\S3�C�Z�=S+/*�c��]u�	���=lŚ���6c��:ǄL2B�[ۄ�FӿH4N��`�ok+#��"j-T9�!�`��P�LB�D���~U���;��r���~Uۚ��`����Q��)P@	h��C���A�/a��d��b������XP�ՠu�{���6��ڼ�j�j��D|�}�����vʷ�~O,E՞�5{Z��*���rn�%��e0��=�L�`'��S13��P�*t�
3�f�B5,e]utk��껮�r��Ҟخ�f6`?�.9������ �Cl�ye��P� r�Q��Z�鋾ȳ=��]*�op�%�0Tuks�!R��Q�Wʲ�6����P^�}��N�D�x�»o�����-#��n�6���sP�3i��ګe�;)��|3T����3�p��6�Nh�܁_q��o9�7�c�*��8}U_}_P���N��L;������{�ڈ=n��ZvuK��Q�o��Q�2����N]�ϟ�<��m��[��[l<3��-�\��^��Rc���zV��<@���әgyw�#9���^��G½��\"���*ү
���y�}���2�����������6�?��^�d7�Og+A�	)��J����x?�%|}o$����D��:�'�+P����G4���F�+v�b�X��/F�؂���ܥ'��y�_�ޝ����3�Չ�1Ƣa!����t���!N����kVX*c5T�u�ٝu�r�>�J{/��g.��iGw3�1q>��.G���0�%;ld��^Ҙ��E�9���ڭr��"r�ݯ�/w��H@��{>/�ZVО���W�<lF�V��ٌ��nXw����mm��&��q��aS}C���o*�/�|ֲ���7G�xIU��(�G�.u��:�U,���U-�u�O5V��N񫘆�*�J�s_@Vۿ����:��}�jv?h�:֦�ъ���I�7�4�?74a5��tg��>3j���D�MU�z�9\��T��f>����f�c����GvPz;��[�z�L�e���B��{c'_ѡO�w �����WH"j[���s�����N��.�gY���������g�ͅgr�S��fU��,���{��t"�i��H��x*T�Z�ە��UY����U�܍pˣ]0�snL7�Xϝ;��B����&�_����߾ȃ۠�eyu�%�a�#Y9��tì�G��{���
�Y?�wa�v|�+Ԯ�xS[ӕ;ݩ�8�!�X�-�������
N����a�����Ɔ���3��ňf�cf ��;gٓ�Y��>�2���6�z�<�+S��x�V8�fǐ�ۍ�Ĭ�6y�AfB�;�N���7�0��{"�R��XzkE�U��YS�95����v�˪�'�"�NsI�j��"#�n��>�{#�����tplPXϮ�3Dd¸.�s��#��x�p�;*�י�3���?��a�<_{���r�n�����s:�xtK��R[ݭ'i���{������DJ�@�*�eƮx�߸|������5�o	�Z�̷�[���c�0�{3E���HC�j�\��V�u�:/�V5� ֯���J.�ߞ�i�+�M_2���z���)�1@24���̬K)7=��9��r�3�4�Fs�����i�;4���К߷�nS�J�Z�ܺҹ��<%#�_)�]����g6� ��������M���~E�XT�%�j�>Q0������}�t���衊�Bd`�}K���	��#gG
��_OO� ����<$db�`��}�����ȼS<#���~�X+E^}Թ���l��2ꉮL�W��ȥT��x5���|]����ǻU�8ޚ|7!TL�6^C����>����ѽf��>�d֏E��[Qݬ��/i����?Rv�ƩH�c$NM�멛��0�e�3�苙��n`�����i/V��&G�pn�����qM��`���G'{31lО�5b<�<}MN i7S�Ҷ^y�kji��"��Ϥ&7FDH�����hÜuE��R�������K�;lW�|��f&Hp*�4mL��>�1��</�2j=��N���m�~7a�W:L�m �DړT�T;�;qWp���J!���S�G}�K��d/g"��)�iZ6�j&��hdfW����]���d��و����Evk�U���dTqWO3W[C�i]���v.f_��c�V��؍� 1W��7Я����t	���/M����3X��ux�s��;��u+_ngwt�b�W�6��fU��b 7��>B�V#͑}���LM	�49/�������e|�6Y.:3�<���>�|���V=t�����Nf�OVP��6��A���E3��ItJ"w$:q"k�Ͼ�����*�MN���-��� �xic=wf&�`\7P��N��՜.J9=``�TY�-t_3Y�U�_�Y��}%öc�RF�mDcu8��퀰ACw?t�z��&`���F���q���e�+Vh��U�e��Usk��~�L���h�"3��@��_+ت3����"�o~����N���}xpD���5��k�:P��?+E��t��`s������ւi��0��/�ѭW��7�&�O��k�u�]�w��;V?*�˷��������Ӓa����V��N|
�J�WS1�+�)+�!��A���
y�o79Y�C1���M|���R��9��fgf�7^Z<{A����jϢ�̏mɁ����n�`o�O�pi�[��.� �t'Bc�?bq{9J��U=��g{WU����=�}m�� lk�J�����p���N��jsp��L[����1	�І39au�o�*E.�Zw8��Z&Yv�`�9u�pj��H��k+Mp��>|��|���j��� t�m�3"�a�����#��x��Ў��c'愫�6wl;�g^
w̺��7�xa�h�9�Dt�p��
t3�Y�_,��-�S�L'�k}�Lȡ=�JGq���f�q/��["�3BWf�*�T�s3���d�M�	{"i�t^.�DG�}��Y���W��Dsޒ��O��6�q���qx�}���|-Sδ�|ζW�){�t��/�du�ﻺ͆��J(A�w\	��� z3��.9{������@|�wb�G^����1��;'䈷&U��̾��r�A3\��S��- �%6Xy�����t4Ŵ����.��[��a�k�󨍖ꡩ5Do�T)΍|����=�[���ġ��	��l�;y,�V�����Q�ڈ��,�LV��s�Ν��Q�Em�MȾ]��f��MX��[���+\^̪7�g���.5�=ڼ%��+���nbh�Ʃ�eyf����p�W�cDZ9��)�q��&���S�C��Bg���n�4{��3�u��W,�f&\ou��Z��-�ѷ�ȸ���.�)���]��k<J�yz��|��y�x�9�ݨ?��H�}�z1R\[��e��5�l񍩮�*yV'�g�lw�e)CV�ͺJ��P��/���c"�G��hr�=�j�ݹ鋯g��Ь���M����>��u���}rJ2�i{��du׋�?�ί鏣��p�S� �s��Ҹ�����D���������Fi��]ь2+yƨ�z
�>�x�K�_d}e��XZ�+Y�Qgv�r�ׯvM�,�.�L�f)���Qca���Of�U#�XB?G��}����(۹�V��u�3W�1qr�*��������:lN�S�:S藊r����mj9]qz��fb�U5ĉ�٠�gU;���LM�RЂ����\6i'iPԫL1w ���4W{q�6+�r�Y\י�(v��K�Mk o�Õ�.u�wX�9�Ol���s �b��x�$��2�1�O�b�!B�T#LL���~6������p�Ɂ{t��O�����[T�|T�ϝ�3�����L��y�&l#�/�1U2�YsP�07rݞR4Vd���fR�j�ް��;�03a9:��c;��0����2��	И��C���{ٽN®;��Gܧ��|֋�Fk�z�`���&b�3D&�e�_C�3���'�Q�\^zy���;�gx���c�_����+�VxaK3WJ�wn��D�Z�8�.0�`��ۓ��F+0[u�LL����D�R�F`Vj�O�c�U�=u�.��Z�~�s;"VF���nt��0�T�[�f�ˬ����f�p����aYu|��cO��y�3��<2�FI�(�vN��̺v�i�>��y32�`L�����qZ�.��Uw�;�p�C'`P�Ȁv����`!��My�v��1I:6��Ad���MC��ӥ��`:f�ܬ��8���mG�i�֍�t�EJC[�����-仰4p���R�7���\��峿���ﾯ�%:�L��z5�7����-*bX�:�g�:���O���$t>�o� �]��ޔ�/GE���{<��K�8Ǫ�ݧ{ő��9��Z�^�>5���|ɚ��gZ-�����-�c��i��׭2~����ti��AX�<�|3�ucY�
pu��k�r	�ֱ��edm���d��;\�Lܰ�ݹ�:�3T�91ˮ)�ήY��`L&;�"6J��^k��>V��o݀�YR���!v t�^'��f�kG
u������J�7���K��!�e��)nM���Wp�����p��<�Q�lo̺&�i0sؘSwU�{<-�����r빟�N�y�N
h�pv:?��!@lJF޳O�}g��l����i�
T�{��I-�������OmH��NL:UR�N�Y%�وH��;��M�wh��ɱ7�=դ0�����O�����3+�(��> R����F�F�\�ND�Mד�oy�C�����,�xݝ�GY{�/���^����o�05-��W����9a�㬭Y\E�:6C�6&Ҝ�ZM���.	��T9��fͭ���U��}&��]�*�ů��ֈN�[eqw���zxrs)'�n�x���Q-d�0�o�R<Hc!��37�h�V�]s}��}�����ؽ�"x�����jb�.�������c�B�B��������N�-
��x�V�ԥ�-��� ����ت��c$������F�c��v�uc��xb/�S�'�)y[;��μ���͖�㭻%�V�|��sӯu��+�h�=Am�Ap�[;�Y���z$M�� ��e-���`�X,�tp�ܔ�F�=���,OK:�#�O��8qWB��$�}�q��z��ɺ[@V��~�˲���:��L��A�[�\��q:.:*o�	W�(��|Ę��/'�~��y��]݇�:S�#/L<	]th��/���t��X�X��)���; ��tm�I�1p[�\S\'B{���qA˸5x�2�]A��r��a��2�v��>��:�=w5�*(�R�@���1�?�Θ*
�-y@rS|�*����]�u�h��-t�x�Tu��<�������3r������:���)��(��5����T�L]oL)CxO�t�v�F�=�wi�tm��c��I���p��9�Q��v�k!�U�?u|O�nLm��$e'�w?	b�r�r�eD�:��R�/�+��W�����k	���S�<xU-�j 9�i��a}����NĎ&�y+uU[Y���4�1�SAJ�z��wl���7�E�M�U*���R���?��������w(�*������~R�ۆ~��h�v�9y��h�쎼%G�@GrIo�k���h���� kԱ|�i�n>qq����>�N��'Bc�8�l��˯	�f�1���q��.Uݬ�qP:U���
�3
{1�i����,}�+�V
џ8�f��.�z��d�}}p�S[�<M�Z1ҥ[�Q�)�W�]�B)�]jw���'U�}+ۍȇc̜F���!���G'w�S��8��أ����ک�^�k�ڍ�V]�U�b��%�c�7��c`*��b�)��O��l_H�͈�p����>+_N����Ϲ89��Mu��m_�˝���P�kG{������|4�R:i�B������Q�4T��D���b2Hkۄsmp<#fE��`��.[��4(W�Q��?Bu�gm����.���~����/��6]������~J}�]1�ه�ʯ�@ju<:�1p�K߫9�1GJn�u|��]`1 #&��N_���V����Cw�g��\�:�UD.�ύ�U���9��n�7�W)��wA��=����`ăz+T9����1B��*�T�r�\Ք,Һv�δ[WS_;<U�:���c�ֆ�Q�7u2���L��d�r�<Ե�5����MSRj�{2���ux�`]
J��z,%��n1���r�_;.�w`����ʕ�:��`��\m��tz����4*4��v���P�'lP9�e��3,�rb��x�/��O&��E{S�
Yc&V�.���|i�ʆ�E���R
�N)���7�w�C�Z_]�gN�LS�%��]m��D~�i�X�v���֐��O
��e��@]��Z�l�:�B��77���x�&����n	�S��]M�ef�
�j^��#m���M��e�9M*��i��J�132�)�+`����:t�j�NQ�b��o�B���*,j�7�!�	X�SW{�T�8�wi�*�V�J�.pc�EDt��4|��Ǩ��э�[�VgMq�l5sZ	�.eyp��!��j��]��壹� �mCt��=3���48jf:RP|2���P'd#o,���!����N�+�k�����*23�]�-�R�r��f�g����P��1�BWn�����;7������;�(؋�屪�E�N�b���j#�\��aY{�s��-�ʽ_8���i�b��yt!3�D���:2a�CX�B�4jB�HA�n�R�]k�G�d�Ne�g�Ch;�	�k� �Ѳ�΁���.�z6h*��P�f��wہu[��5������e;/C\)���I$��U��6ު��ق_�c5��ۊn],-��_q��j�T;;K�u��J�aյ�{���{�qŵ�hj[l"���f>�<y�
�NS�Ѯ���ԛK�$��3u_K��y��BQ�{9��ʸ�z�.�]Ye�'�iGC��X��q4�c��˺�_M� ݚ�+�^�6|0=+g*��^͏�<0���R�H)y4>��t�u�qC/u�l�")�]%�9p��Vj�Z(�MP��N6�b��t����ɼL�������^������t��uo��6���v�������jj�k�{�T_JY��j�Y�%#���|�q�C��R�����N_S3:���餃#����]��;��_��nr�OKB�}�u��ImtӒf��8����M�րec�&i�)�k���x
��Ρm�����.v�
cu�mkl�̰+NWU � $/l���%����d�6�s�;�'r�+w���푔x+/��ݪ�k�2*�\�$*V�P����vb���jV4�x�;&ֵ!���;6�3	�Zpq�z�>�Urb��F�M�|�6�GP����=c��6�e�+U��e_� �T(��(�Q�h�2BK(�&a���  `�CQd� �!3	Q"I"B���H!�T�2��C,Q�hѴ����B1��E@�j$�)#D�)1X��62h�Q4���X�AE(�؋I!��&a�E�b&	�Ѡ�&J)1�l�Q3M$$E��lh���`ƃF���h��DDFƈ���RP�2&lh�����F��4QBTX�M-��,���b��_����{�׾����_�޿�mڧ`��z{�r��m�0h�f���7��+3om�[��0�'r�O�F��ck�,�z������ꫭ�4�Ow��;�X��{\��|�����vZ<+�)W����d׆U��&̫@!o0���>����s6U&j>Z3޷�7}�q�vq���*�5�ҹ�0,q
��<=����zm��ڇb3����������$�z�ѷ�����~�v[Gn�{��ѩTd���֓	����oS��#]&#������5~�[Y��e�Җ�mK�7y���*�����C�z*��Ó놥;ldN�)��)�ݛf{�y�r�b�c9��V�a��@f�~�3˅R�q��cY�8]޴�\&�tص�F�G	�!fŅ��jUa��^t=��;�e*_r���D��>
��[NWq�Ub�#p���+���}����aIoo���hk(�E#J�oô�}J�o�G�Ҧpz�Ny�8u�Gf�sm��ϝ[�����T��!cgf^I�3�!�s��꩕��:臽iA�eƍu]��&rmm��:wc������o������q�Q�#_z�!�]~hP�bN��r�^kn��v����+|T[/���\(u�S������Pm�����Ϭ���%KB��_G1�~ލ�ō|�[����F�k[\a��tpP�\N����e.g��3���GzM�ojW�B��l��3\QGw%�`]�T-���Жq��o5M��k��;�{���}���}]�zOg],A��
�K9BU�e��;�F��-�1�f�-T�`��#�-t�]|�u�(�䣡I�ҡ�tW�`a�u-�΢��p����=���U�(V�j�9�{�ɒ�X��5�0��2��3�\E�,e)f]�qXb���)��pxQ�l�8|ώˆ���j��{#�6��F*���M�[�#Z-�+u��>��|,+!8ó���j�dѧ9V��-u����~�"{��P��c=��C*����	�i��z]/xF�s
�=��C?oZ ��Lά�v>)��%I{[�֞��W�������6�|�U��ݞ���V�T�86��6v�?�chӉ�2����ьB���9��qΔ�ɝrr2�ݟ�E�V�y �'F���1�-ʤ!��	��97�+�t�H:��Y�8B���V+�
\�Tn*���@-'뤸Mf�kG
u��������+ZD<S�t{V�D�3��%��~N��g����4��btL�Uy+���gW�<4ĵ�΋��VUС�����{�K��_i�Zq�Z��þӧ���5����kqӢ��3��7X&0���2����ԇ��z�۝ݝ|��5�4Zp��2�[�PӆU��[�{	�Q��X3p��S�����DO����D}�r蔒B�}dLz1m�Ԙԛϲ;k�nC���l����-�1�q�w[z�(2Ľ��erQ�)�|xd#�K���O�/s�����~{BvaҪ�N�Y%�٭��Gãڼ�z���`z�ͽ� � Hn��_�m4�Qwp�<�OH[�d
_?s"ٙ�J�`��~��O��b�OLLK����J�dH�������}P���@SL��F��vF�x�h���D��DieWi�J>�_h��ػ�W3����(�69����*���^k8��,��ok��u�D����7H֌&�U����18X75��+6�x���G�~C��Q����9S�y�i����\c@�Y�l��o>ǿx�Ewr��fK�>����{^N˩g�e�:�� �<<=�-�x�������y�p�Iv�O��֍�"�{����xi3{��T�V,{��U���|���U�L�uz_��DM�./p��$_����� �P��Y-Z�CJ�4cDF0�8��v�x �����q�Zn�m��\��ϋ[Vp�Z�<��3:l-=��V�Oz���c����En��&P<��H�I#��e�K�f�cBI��0����aX-��i�3���|��YzޕFvC�]d��/�˚q$�����W�}_f�$�H�b�j��Dd�I��>����^cv�F�(Gm;��x�F�n�w�R�0�F\�P�;�ac� ��s��Ô*
�.�(Jo�Uxpq,N�n�TÓrr+3Hri$��:�Ui��s��|ڧ�-���(�=4�� V���U�� ��� 
��^��_yw�8��s�w:�&���Y:՚�3�����m��~
�Ӕ�*����GQL�������~T=sX��,t�/L<����N{sY�ٿ�7O�F���Z��r���^:@04ת���-��pip{�.0�!%_N�fap�=Z�f�χ��p��$�o��~������T���h�y{MJ�\6̝��?=lŚ��Ė&�0��FZ���6cg���7]�&�����o������٩��_c���\�7[K�D�i���P�e��,DuB���� :��z(��Qx�T�]!�R���U�]��6$l�q��ʚ���N��\����.዁?Tsb�A�zr(뵖�he}�H�eh�bȹ�=i��-#}hM�	���Z����ɇh�If0zӮݾ��/����jD�Zĸ�A��Nk2�ِ����6���Kw�/�iu�/�p%��G!��l���zv�f�Z���U��Fe�@������[�C�׍�n�)�Y��g�h?�=���U}UU1jչ9/y��ռ��b�\�k���~��^3-o��3S13��(p����,�sl�>�]��t���6�)��S�@c�l����L_,��"��$��FMCd��:rV���5�R|9_��T�s?_ hC�gג�V��Ч�Tc��E�p�� -����F��[����=(?�����WfV�Vվ-1Z��vJ��1�]ɴ��
��3ʜ��G�#�vv���0�;
v���`�b�Av�#½��;����dׇDr���4��I�\��g�<�9�#��=�F�nbd�O��Y(�ޞ��HA2;�������0��
�,E�Ra�eb����� �}�����֌j�g�s�^�gz�ѷ�-M�y)w� �}�<Q��˧W�
}q� �aZL&2)4~:���a�t��w$�YÄ́7�'��Q�w��y ��Xj�L�O�xE�W ��9Ó놢S��};0��ً�9]+�nc~`r�i���j�-�`�\@fϟ��.�p����}��i�=�s���h��
��~4_E��:��	�g��6��پ�x9C�&TZ�76ZP�7\�o���*�rP�N	�P3��ufj�D�`�+�9���3 ���|�m]���%�%���aƬ^:�~�����x��y�esנ"���}U���-���z�"<�]�2u�ٿ�S
����)������*�1�%sd�.֧�N�z�{s��k��:%W=�
�P�f#,�Њ�p���&�ۊ��X#&*�qb{��.����#1JYn�
r�3�R9�ɔY0%D�u0@\6�U^�0C�s;���h��b�}Xk�2u�x��s�����4�ޅ�oX��L��������	�{�`x�Q�o�ѓ(OiW�/�C��FN�B`�й� ����L?{���\�m��ޭ.�_h`���\��<*�|��o�u-�'V�aI�j���{ۙ��oK^O[��ޤ3w%�W�PlF�Wp��e����P���4�6�z|j������?���Zy<��|W�dK��n�U�)W�N�j])�0�e�zڳY�p�Z%�u���<!u�!�Я1�7h�POn闒�>߼��gv�
�7��d�x��C��zOL�^Nu{e�����)u���~Ӣ��y�G��:1�ω��әu�4S��oF���^����ht����s�j�ϸ=c�#�6����j����Q8�?E���+p0v���V�d��p�7�p(����z�{at�~芾택�z���:�#��ׁt��Ӗ&U�.�`4U�ݬ�4�	��*�N��%#�J�(�zx�W߾�����jg����;6Q�����S<<��O�����F�O!�C����އ!��X�.ƣo�FҺ�oޭ����}~�q1��yx����3Q��a�B��	�ή_}c��e�;�;<�5ޓ�fM�E�/o����k��e����x��#�u����~T�Ҽ����m߷;s^_��m�;j�����$�k�2%F�����Ր��λz��sq�H���m�i�~}=��N�m�[��	T�%��+3k#�4��ܘ�^�(zrM̭��O���K���Ȅ��bcy�Ɏ�ߤ؎��s�)��yQ�U_D���{�1��1�<~Oap�3N�o^;���*+T�g����'Q}#�[�e<�Դ���|�۝�HR�K����>��8��{{a���f�v�_m�\����79N���/7����A:ߟ��噁8ע�%���h5���4��9�{O���A�	�VK�W2n�<h�����,��uڮ�zT%F��UX��;zf1�ev+6�Ⲹ�!)�o��5�:0�	��Z�6�e��wWhĴ��M���{jd�4�`��=�v�g�ACr�uW&u/�DD}Z��]�trG�=��72��P�[Sbs\OZpg=�슷ϧ�:�e�]W*Yُ{dU��oa�d덪�x�OU?[:Se��6�|
�x��xo��㕘�:��Z���휅9G���'��������S���6ԫ���k:����q�3���fYLʼ�-�3/c~w��D�/'��6�����:5��9*5-�y4��r��,�G}Ի� r��I��rs˖�A܎�A�u�{���ݼ��H���^��MV8ݮ�h�ɦ�-���e�/{ �>�/�]Ppx�W�Ní^���V��@���;/�t���o=��0�����٣�����b��ռٝ�*�O%�y*���l�X~[=H����.e�Pզ��%�m+�gI���F,�W�\�r��l�xV�U��p���s�ʫ�|�@YW�Z�;�Lu��')�T*�k��W�f�DU@�u�i]���R����Eh��Hi\oH�Q�]�v�#kep�y�5��C�{	Eif�A�9��2r�+�5Js�ۥ�,д���OTӱ��;F�Vm��L�i���U}[��(����6���B�S�ba-��D_U})������)׊�zN��(j^]��g?@��~��a�V�L_W��ns���E-xe�gS�ڰlñp�C<�՛����`���{������m��u<|p;3"��z���_ҊTF�fިz�Ț�����M�}�%�9B��%��}�#.�ۙǴlb�W��%a�T:�MC�[Sbaཝ��ݸ-L-t��$g�d����;.��g�ڶE}����/��ok���.˦H�9{Z9uʬsd�֏|<��c7��3��b����QQ�[�མѩ��5����_:Qj�}�C/�s��c�5�Yb�b5㛄bo�m=q�o��sݫ��Z�WIeT=�4�o>�ioÏ��8qw!�+#�� ׍t�T�1��7I�=���z�����ռ��buO�M&�ߨq�*w��V�i�]X=0+{Up`(����"�.�)���*��Lд/ꎐ�V�/˓�ќ��V��ǝK��evu�щ��� �o�q�zq�˔*}�����5��o+�U=�H���ݥ��/�`Ԭ	��#TZ�d�O"��
����節H�z.~����ש`zC�Q\��r���݉��ԥ�T��3��v�wC/v���a�>��+7�;�>����ϙ��{˻>��
���t�(�w]W����+\OI�}�E$��]	i�S�s���\Q;X.Zɬq����7������Ӳ��d�޸�uR�M��[=aEQ�î�q�۶��Gzҭ���E��"�r�%�ˤba/�1�3랇���[�`�E�h��|O9۩�ܚ�F!����#J��.َv=V=��R�����E���|�5^��pN�K�κن3���]�D:�s��$�EZ�柎?#;7s�
���y�VF7�g�$��m�����G[��B��C��1����,z�Ъ�J���V,uq���+�1t⩥��k��ۛKG-� �uJ�5���v�]g1mQ^K���N����Cv�hhjK�\7�w�4�cKWb�q�Lj��u�Mq[,i�iN�Q�yn^s[k��9�[ҵ�ࡋ�j����Z{�X�QH(\��Ȓ��JM�'fG�qg�1w�p�<���JT��[��¶7�r}��䴎���Si�q?�xn5Z�1Q�p�L_Xn<��;y241����[{��R}��a�]���Gp�p-��(']H�N�P!����V�{�d�nvu@�Wn�`�8��R�.��5��]A�g">ӯ��+&�[��'/��48S���uv���MZ�.+�6BS�m�6�(C�\y��Ԫ�.�	���3�Y��q|�5���&u�tw6�͊d�����f�.4�5`�L�wЄ;�^^bVv������D��X���[�Wy�y��j��:��f;������q�R��12]��a<�����Z>�b��t#Z ���'4u_eB( �=KP����HR8E�ZO
7ڳ"���hkRU��,�$�E�̃/�(�@PJ�&��a2�oe�eG��٭ V�Q��ق�
��i��M!og	�j>*T�@��6�#�y϶�J��ѱٯM��L}�+�V*`p�5{{C�/\��us�l���΅����Z@�¨j���+�E�.�a۩ż�R��S�.��Cr�#�YW}]�Áb��1��D��>�٩��8�#�w�ݝ���
moF�6y4�ͽ쬽+y��N UBК�e�c�4Z�Ut��nX�ʚ-[/���ڎ3d��q{e�L��	���ͩ����nZ�.�t�����O�e�o�9�v0Wk��Ĭtթ�	��<��(�V��s0�����2��ٕ
��01���9���>�E�,w��[��Vdھ�P�Æ]K}�n]N���
�C]e&;/X͑�v���5�ʮܲ�΅�Vmh�r9[�|1��+�{���]Y���3rlZ�tgu�Q�F�Δ��Gml�eغ�U���VT�&�ƚAĹ!�iCkE����x�%4�H����� f�]bUd�Li��ܼsYo�> p�oᛁ�:��X�b���7�:noY�R�ޭ��r��q=�%b���&�գ���=�/��u��X���ǒ�=l���i�x�=�'�������WE�i����Qhn�t�+�w�� }���cj�i�߳\|��n���}�r=�Q�.u�i��K�+F^>���]N�N�n���r:K�f�I�� �ʏ��Ցl�R0:5��4c�k�E3HJ���'a]v��y�MW����S�W��N���+J�Q/!�9d�:z\�xj��gm�:��ӽl!�/��LV�T�<�{��6衖Y�%��� bnB��T�
3f�Y���K�y�{Z����~}���S.����&sb�iΙ�:�U�@�e��e,�gb5�i\��sP��N��3��)U��}$��t�јv�X7F��B�"�VV��^q�Q�h����V6��pvλ=xP�O\s��!2�p�5+z���/��R�ӵ;k�U}j),�h5A��-��&D��M6)��$m��#b�b�"1����*,lI��mDE�lh�cb��Q�,E�ьc&�,a	,�j-&�Q�5�,Z66� F�X0lh�Q�""�`���`�`��4���V-��h��1�j6�b1�AI�lI�X�m��,f�jJTh�k�M��Qi1�����i�����'aT��i��A�\�eg]�KSV!�جo�kupes�c�條7�C�Ա/o�����vj�����w�z����yM\����(�+>�x_{*F�j���ok6C��oV����mC�u'�/\�\@]�1�4������5�m.�,N��v-��v�՟��>��fy=�dSMqJm��V��oD��W�{��'w��~�r�.��]K��t��
K�泶L�L����,��-�j��Cv�K��v��Z�#���>�g{���z:���[�֡ZM����D�/(��$Uq�����5����[IκV�NC��c!,�{z.��ŃN_>I��N�
���NƼ����J��2"쬝@C����\b�Fy�{=�ɽ�E�#�j� ��}A֣�qo��jR��ؚ���OC	��8KLF=�����W�c�ȸ��ʻ�B��ݥwDm?�j�%�����k�XO���(���v�iqn�݌��	TN�]�e�qwA�\;廠jc�u�����;�ٮSܵ;�\z&��U��^]m��Fĳ��_Q}�u).UЧ�`H��Ԣ�<r�}-���]}�4xsV]��oEj���x-p�1k��Q����`u�8q�
�u�;��ATa���u]��}����]��x�ʯ����u}U+Y2�3x&�)�z�`��^R��%�B3lFd���~��~lt�B��[/9�������v�8�㝸2H��i;'k���U���y�3̯�����؆.^j�v�n�WOJ�붝<Z�u�p���j�O"n8̈��"#��ޛE.�T�gf>�1"���rE|�;�r��+��N�i� D�k��+M�{�j�,�F�`#{�?o�ۿk���l������i�g>N6��q�<<̙sW�v�����fq0�X�l�vr��=�n(=j3�=�b5F�%32)��5½Ҕ�j�q0c�Ðw#;~/��uF��(�s,�ZϮ���횮��/y�U�ӽӇ3�\��5���v1G&�odU��ZҔ�k��B\���r"�m��Lkñ��=?�Q��8��ŏ�Q�]*�A�՝o����%��$�u�ݙF^���`�������߲w�ɕ��;=��Y���������(8�[��2�Őw����X���ˏ),������L�L̏6pU�Lӻ�x^�VC�La��HvNT��Y/�����)���o21�Кkr���X�!�9�>��>4-�W27^*��"&�ֽ�F>fu�?=��)���Q�adwV��%	G�=:�w+�n"n;o�qM��A��-�E��M�/p�6����.�V�0.�A��V��I�0�NBWN�%.������p�O��;���Ȗr�(�B͛[���ؿ��H�0�؄���O��]��jp��g9��ݛ������t��ǝgJǺ���T�\r���DRא�"���lY��y�%;NIV�!n8�j9>r��0y�����d"t�]�7�m��]�z�?=�\5��"w�w�痝ۦye�V���r��GÖ�3W<�����Y0uP�}a$���.Z��7�h�.h��c��կ�%a��7�Yl��4Y��h)|}Mp�W�[7�W�S8V�{q�E^'|�f��<�!\4��~�y�㋍�'w+Ց�%a����E(��}�׵������K	�<^Mc�M�"x��z��*�]��n��6�����z��Q�9V�I/��̥Nc��.��ef�r�R.N���Iq��]����X�*��ӻ��n�s�fَ�K��. c7}���e�/h�P&n�T�/,``h��Vd�a�>�2{�T}�e槃/��K�%^�ο�����	,7��"��_u�kW��'��f�A�6��_�FHF�0�p��3LX-rU=��u�gF+��s��oe�mu�]�����Ei���>�qCc��BD����T8VMG�;����{��5��I���w.7������_�T}BH�Z����Ɵ>k�ᇩ4�eyi��SI�r���ځ��]�(���r�|�7�z����]�[j��/�_iZ����	��v7��T��SF���b,��b�]r\b\���q�/����\��a\�*�����kd��=��͋�Y���;���E�;��qO:S���Y��U�&i���(9�!NE�fS^���W���4VU����v;�!7q�/e���Ίࡗ6���F���}�f\��'�13��8ՇeW`�h�Gzv����ZMpj��w�i�=grܓ"�w$��݇ ݝ�;�p[�]���hu`��:�wb+��k6Ӎ[�q��2)j����<�M.?s�^|�)F�Qn������pĉ�1Y������j��ܬ�ݎG~I�������⻯m����Jժ��(�P���^��[[�UžC
��?NYݣ���-9`\�����)��\%,N��O��EE.Ҽ+�B�fK��p�u��Qɥ��Q�T
蓐�Z1�����U��'<�����ӽ��g<�|r�1=xrC��I�t�qr:k�-�����T�>ٕ)z>�7�Eh�[��pr�����*Zr~oI����>άDɚ�٪Zʹ��r�-��8�4��e�����z���nKU��x��ќ.�b2r�v/;y���=��w>�uz���qȍW����㨫��B�8Fm2�e�U�R�}�p�&~~BB�L-�gV�r�'x��{Х�EM��+�+4_�j�
]���g:���1��Jыb+zf[�M�%��P��}���gc�`����]�eE�ϜV�>�'\69�0U�e.��O��v-�I̻{׸b�t,:�n�Uǔz��,
���k�l����n����z҈d숨[��ě��xa󖹽��R��@��
������t��>!a���}�O/UL͸��������	��E�<BҡUD�pn�]��+�����fӛ]7��[=_Zz.i>���z�ۧ������[��ڥw|��~��)'[U����.�pw�S��͔c糯E",�*�OQ\���p󂹆��BU}U+Y1+��pM4�C�M�Ʉ�	���Z�{ul�}����B4���v�^���0�Jy�8,�YUm*&b#J���h�#o;��k�ۭ:����&c!:ei���[�v�ʗ����$7<�wK��㝃q���=�d;�&���>ہk�<��W�gy�W<:�O;�gd����H����~�^c����m�v�n�?��Rm��&�F�s{E)��?;������Tk��l�go<���|�ڻ�.)�V)���ww�A���k��voi��y�]w�gN��KnZ�7�5��f���.tO{�0;s�p�����űd�qS�z�kyi��� l�	k��#%b�X��tΈc�3�ӥ��w���k�+�q�]��뒐"�ɭ����ԕ��:-����+�k���{7�Hy�]X�5ױANob�:L�}]�2K���>���S~>������z��U�pF�~�}<�f_��|��s�^�1߬��.���*���7�iъ9�v=���y��flvh��J\Am��K(�3�q�t��ȥ�����ړYj�f�s����+/��Ʊ4����G�<{ pYj)�B����P����Pu�)tT^����]>g�7���K���TN���|U��q���S�OTJ�W�R]7�¶z�z�Ji{/�J�.�n� H��ܦ��\&]�(H��U��%qN�.�8��}����i�W��|�I��"wlt�d���3��](V�:5ܩ�UC��|;n��%&�&���-E����=L�vx�s��3��-=#�_M�nUZ�l�����y\�ua=�]X��j�}�c���;(U�L����aNr���7��j�au�/z*R��:m9�h�n�ޗs����]������I/�:lelc�f,���l&�ݧ9gf@^�㻗;Bk��v7W�k2��¶���V��%va�OJko��ل`���b��:l.�5jV���N{sƒ��=MX��E��I���B�9;e�HY��,Lj��;Js*Woz���'�\�C���k���g˗��=���,OWɨmpˮ�yAʻ3�q�C��ۆ�J'��8/��s�{z�E^'|�{X�����U�h��Վ,i�FWq��b��,?����vA+�7��7+Md��o�U�g=ʸq���˂��ڸO_��w%���b7���O���o�5z{F�K��zש��s����%<���ub#v8�e�}`"-ox��cu�q��;ny�T�-3�%�j#S�8�����ϭ-�{7�|:Q���e&B��ev�r�sw)��Ώ[����x�"��;��y��}��2!�3嗴ֹ��vu7��� u|�
��G$��_|�[:i�]�
��3s��� Xx��:g]8˙�e-7A�ﺴs���	��������)K����t����gn-�zb�����p8�++�8^��7%]�f��oQR�L��[�gv��c�%K-��)�2�Ʒ�|뻋���
�!ա�{��=�o�mDS�9��~��mOj�9>�0:~����''��Yc�ʬ���5]��$=��Fs�4o{8�c5��|���%�
�_��K�P�Ѽ=�l�\�Q��n�C�X�;1�S�o�\ri>���K�ie�3	|������\�<*5�6�%�&_2b�e�z�#,��*�d*صp��5��[��{����u���ܯ�d}]�!q;�4����[?1�<[�@ŉ��R�D5
o�\�-�A��0�Ц��j-Ȋ[�g�{�L;m�4f�X8���HT�궻�'�PSc��.�o���7��W2��.^�T�?�
����ԯB;?�P����� D�c���4��[q��Z�p
<�Q�
�ǖ����n'���~��o�+��˷0&�3:TIc������;�T^(��l�5Z�y�t=7V�������0w`���w��h�F�l@���%��zzR[�g:���VsʾYD|4��*���0Ɇ���*��c
����ba+��Wm@�vj�J]��zbԲ��ŧFR��b�gLǉ���];]譩��
��9��7�[��D,�G�1:=��;Gu��ˌQ��=�9ϡ=jOQvu��B���ve�<���=y��ھ�c4k��cb:�%<Q�ݘ�e�yv�*pYz�p�69��ӫ\=�����f��X=�}S�>�\+�K��Dez����]�ѧ�7��iyԨI];�J׭��1ɀaU�j{Z�2yᤶ�c�эM5��ʭ6�]+�'�F��Q.0�����9��Qv����}���S�q:�-��~I��B�l�;+T!�v���nR|�8K.v2�P۳qܖ[=i��i�~}=�~{9PݶL��93�m�����Ղ��TN�+���|L�d����I*!�&�V��;�V���l��;v��H�l�U�bV�bWf���i� �M�U��ƛޣ�����9i�./%��V�N�e���w��ա��[M��\�N+�¥k3�nH��\�^vfn%�\uc0q����YB������c��k$g��ѸP�V��ˇ����&Z�S��y�^
�#��9⁽��xa)Tf�J��h]b}Y3z�4�0��2G�������e^]	�+��v���b����;2��Ng-nC�$!,�S�lM���`��?U�P:�A��n]s�p_tW;��q=A���o7t�wɪ�����G����������D���3P��5W����*
Tn�Q
Z:wƁ�,�[���V:G˕�J��׎&�Jv��Ӯ�����cha��x��w3n����[��9J�]ѮDe��ٗI!z�~�%�7�tfq�����D�b2�z�.�-P��Y(�y��˺�]�mu99G,Nx6�C��(�!�f@z:�pT�v���ڊ��C�|�E�K��1�q<��M���p!Vƾ�_J����Z�)+@e��Lv!u�Gf���I�����H���=�U��ƹ��
��,[pާ8�&�s��C�/�E=u6�lP^^g$�>6-48c�m@�T � ���v���Ȓ[��
r�S�<uh눺F���S��%#W"��Vd�m0�q��G�3���J���Ꭾ����2V�«r��ʯ��ڀ�5���._iO2ޝ[�/�YOq}nͪ	�k�X�+�`�ϥ8r}��z,<<h����s<5lٓbĔ�ʂ��[�]�oU�R����z�lJu�7���5l�J��m�N����cgv��3E,�8T�5�6���d����j�:ʹ �/+�K �ޫ�Aի�#���ux�kyfF�b�TD1J+���}֦u	t(�g
��.����kTM��husN�BXo�m�Χz�몖�-�iF����ԑ��z���ȇZ/A.t2�5��[���/��V��Ĵ2���q�^��v�gks�O��]w���rsX��Vcpe���u`.�� �w�v���@9���誗�9c�wX��x���)ڊV�oRo�[�ꏺ�Vb�(�s�y-S&iXL�Wg�M��(����X�+
$]c�Z�����e�i�KN�����)����3�C��A��w��e�Q[�Ke�5)2yg�;.�Z.��� ���W�U�C1x��{�d���ևٝ�;:��ޡ�t�+�_ed?r1q\
�M�|�z֥b�$?�m���lm2=f�bl���*ԡ�I��,ǵhx���9j���%���=�m�"|8��8mmu-t,�7����')�����{}V�Ŋ�ր�cJf�떕�����������mS ]�'�^s�
ġ�n�{�c961�,d�9�E��
�|��%���}S��:6�q�f������^���+8�:ܣs�N��؋�@�&uh�墁7թ�}K'S�F�*T�84�y�ֵY�Z{�
vs�}���e_�m8Gi��va�e��u[p���bcӯ}�>���W5%D��DlS+S6�F(��TB����*ѣX��1��4VŨ�mY5,b4F#Xر5��cBQ����k���&�Eh�%X���M��EPVJ ɤ�Y6�Q�A�-�5%!�5#h�b�cF5)QX�0b��"�ű�X�Dj�FŢ�6���TK��hrŸ�n2��5���N��wS�һI>��"X9@`�v��K2����B���B&��&��v.j�6s��lwu�@ѽ{�c��1sѷ��y6�AG&a"�L�8-ir�]o�v����*[����J�[�e���LV����VC��"k��>�2O˹oL�,��g��v
�S+EF<�Qڝ�+�mPW�z�q��8]3TB��Uγ���t��@��Ĵ�+��n'^ȼP>޶�.��L�e�������5��k9�W��췬z-�����m.��Q������w�e�QGs�����:x�)��-�m+�����6�������LgR�i����[��k�c�w9�ybk_�����[C�����8�z�i���j�K͖���sи�;�ɹ����Y����u�=Үt���j�p��$�C�ݑ��՗���h�ַZ}��N���Rx�:f)��$��j�'�yl]��O��ފ���������4VN�4����/��^r�����Q6lр=H�Cf�9U]�<�f�\��)�YQDw0U�Fgt����l�K���@S-o	��P��h4�����ى$z*"M��+�y�s�c�u�-�lY[hw1R�b�N`�uhs���r�R����uaY�Kg4�+��n�6VۅU9�)@��n#3�����ʦ���X
�Q��\���q�v�:��R11ʧa+�P�N��m�Ӆdũ��o�;�ÅX�9�Kc4�!:t�}0�؄�/��>9��o�]#]7�+��'�����i��z��w�l��Z��7��m
�g���uk{��T�O3ճ��+�J��\rk����!�u�]�3�{%�[Z�T6��c�}3ٷL[§+�*���w�#'uqCw<�0JI��ͅGUgꂦ[�l>ˈ���qz7:�On����巚�Od�E��b0���D�(�7��g1YǷ�dTE�sA^��u���z�4�݌�
q�������������}��7�S�\��bΛ溦�p��p���[Lb���_=;W	�[�����mƂ�`��iT�e����=�<��Et	�3����B�.��+5�md��6�5�}+�u�W�yZvn�;�yҝ8ܽ����e�>i2�Vo5�uAB�BU���eb�nN��X
���
��`�oB���7{L]yӆ�'U��y����)�y���C뽘�6(���S>���2��9J��|�-��:P��,����Ǐ���i��Uq��ӘQNz7WSuo���;��u��f��(�u;����-�܋Y��h�+����o��z�]O;����w6ڬ�a��TB�?,p�Qm�Z����Ju=q�{�e�J�cG{���� �b��<�|��#�5�o��Y^�Ўa���f�>o;���(�7�P:�lk��@�I͞KGc6;Tu�)���c����E�Ϸ_i��c�����Q����]��Y�yt2#A��3�RU��.�a�{=V�E�&�}=�����-�FYt�L%]/�uv7y��F�#��!��{��|��kVZB^����KϷusW��n�R��kZ�#Z�an؎U}")k��۹��_'�ˮ�XΞ�P��#�	�P�ժ^\o!��f�G�+�o�Ug5�������D��ի2U����z�p��Y����D�`;Z(��K�5�H�9�����eaT�E�9˩:v�6�p;K�i�c<�>�Xѧ��sޕ�ؔ� ��PJ�(�R���]}	�����yv�0�aF��\խ�/�/T%{��&�E���in|rz����:���/"��%_V-޺/���<��=�T�"k[��&��ı��]qf�h�Yx�e�c�����1s�兖�,j'6�jl^�ە� u��y[�{jVgs��q�6�V\cr*"�F�[|�sS�ڗ�5ކL��ǫ�������W@2��W��\�����*Zra�]<��el�6c�O'vʟf"{���|�[3�a��]��3���ue�Ԯ�b�,�Iv^o�]9Ǽ���N�W��&{%\�W:=j��v�FqK	���Z�is�i�/���+65��1�:����������3a��tɷw[��r4�:q���6��g�:�˥q�j���Ls�~O�2
�v�Z�xez����������f"y�1g�L&�����-�Հ�`�24U��R�.ģ�Nb�`k[����e-	\��Ҿb����T�uQ�q�nm���ZU�wN�����B�+����i��=�lS�.��ыP�W1�r:<�w���VZ�>������z��@�n�)�O_#����^e: 4����-�4�ֵ�����o~����氭��I��i8�x�:#�[���d57���/E�]
�U�u�J�풨.d���]��'ݜHĊ
hg1zH��)��[9[H4��10�؄�辨Z�>�]�c�x�M��%����z�Y�V+֜�����LG
o෦Ⱦ��sI�v�d�zk���k���h��9lrcn�nm0��P�B,t���։]���_�B�鳢y��{�(��v},�%a_&.�5`{�d�c����j+k��;�o��1e�|R��b�c>�>U/~j�MD�F�ԁ�H��ƚ����ԟ]�՝�5��җ��~v3��Qqm�|��c���1SZԖ�w:�s��K���Kj�[:=��Ҋũ=�$�.��{<ԡ�rr�i{'Tm=;W�\q��V�b6k:ྱ�<���;��T���Y�S�;=*W|7!Ww��g2�N��\�k�1k�`�m_f��m�JP�i�z>ss7p���\"h����̠��!�t��
�T7��|�0B�|�g0�ީ�Wv���/��@l��P��v{Χ�V�B�
�J���}{x���2��D㷪�S��>]ѷ9�.��x�泪��x6��\go���=��.'k���u+�:9����ܖ�g}k6�O����r�y��}K������TI��g�]?wd����F�Q���[��Tݖ����3yr���4��3��;�]8��0N������og�j�m*�ֲ���rzS��D��U��Oh��af�U�)@�K���XV�WȽc�Vv�ohJ��e߇>ga��3Ju=�L+���u��rCw�n���]oS������;�����/�wgn�NwF8�f�E�¸�K,BU}Y$�@�-�*;3���V�[��'�ZݼJ��}�NqC�y��*t]v	��:��,2��O�h��M#��0��e��6�V-�1p�������gUH����.�Oc��2��en8���+�؉��+��Ӟ^p�[��\�j�Rߺ����Q�	�ݺ���ιm.w�Vs_7mgp�^'<���O'-�l��H�צ�{"!*R�>7��(�j�������?��ˡϵI�մa�5�{Ȩ��®�yr��lG4P�"q�:pF�r\o�<���W0.^��k����{�TO8�읓�uu�����U���ǫ�����	{T=�7��θ/E}�_ڞ�WN�艣Z��e��Y�m��p�;�&���.��K�K�?��	����p� b�x�w����>t_��*6�p ��ia�x��ۘ�#���o�N�?�ZBv�Nf�1�q��F�jv!_m��������Kh{��M�]5n=�G��p�m��ˈ��a��{d��o��ir�sM_��i��՜�r��\>��
� �;#�1F#I�����Zxb�]t�֘j��l�������&_]P�os��om�hp�ɩN���P��]�*��`�^�@���g,q��b5I��1�@��\R�ZՑ�-��Ƶ׶��t��ś������s����n���g�D��a@I�o�'�S�057m���Ѥ\oXۄ�3<�{/s���t[?O��J�cxV�\qX�gweF��u5� _���0
��^�KGa��Z@ƫ"�bƔ����\ӛ�LU��`,�W|6B�k7r�"�{�'�>"�ƟN��ə�7�qi�������67���t���tc��ԥ��x���z�sn�k3��X�&��%}���/�uZ��{����r7z��h��P���g�J�Yt�H0�ݶ�0b�ws3Oe�q����f�K\Oҹ�Z����t��uq�Pj&��lT���j��S
�s�}���u}"��1+�oRf!���m����a<��f�2�	��V������M��M��0�>�#�[�x�����&]ͭ��ʺ	�=�,(zUdrdN|�6e�[g'��x"�KSc�J1�x�b�ܧ��E9
PمT�"k[��7�k�j ]�vטl����
��VvH���Z������ل7�o4��i-�ѝ���ض���w���nE^(���l�W���g���eTm*���G�Z�#8_��X�n�p��:��Zra�]<��yj�r�̏��2g��>O7��)���q|b��X�۸�]X�a���:3am#��g(�u�6���wv�E��B%�O4uxfV^�����a��z}���U����]ڹE,&���o������mP)�[�7��Y�%e�z�Y_>+/���RQ��՜�2��Z[۵�%�9\,�)�t���9q�$�'�(���!ۅP�or{��1ܰu�N�V��`f1R
�wz+v)��}��o�ߧ�3��*��t��Ե`��#Fbɥ��#�����Ny��ư���o{�V�f�9������U꾡��\
q]��<�����HsX\we�ko���B���$�[ʧ�#����As�B���W@D�l�>k
��OF��/��De��S�"��tփ�ή.ީ�}0�N�W�Qω���>����f�2��N(ݪ�y�yG�Rͺ���*�v��Ε30��J����ڪ�$��nc��Ҳw����<�ߝjf͞0�¸/&*!:eq�O�/��4���3��� J��q�n�K5�W�F�c��·�![2��!u�5�ם)������f�8ܞ������P�LW>��&���F���2���{���]����g&Զ��e䫮�t��`@�u)//3���8�[�mc!-ͱVy���R�Z�:%ܧh��n��V�F�1�.7ZP�<᝱P�zY�o-��Y��U�Eڟ�ZJtlh|�z�R�b_iv�mn�"u�c�K�B��٣ۮ�+
D�n��(λ����\�I�w�w��G�C{�㘋Ѹ�E_je+�@��sq=4oK�Q�'q�p�-�]U}����%T���5�=��J�~vں����"zլ�YF�ގݍũF������F�"5�::-��>(��emO[N^�n.{E�M��9���ʯw.�i������U������R�rt���v;���Nr�]Ō)��q����o����+u<ޏr���=�K~m�Y�v�S��Oc���w0�Q�C�����<Ά��Gq�ҹ��_MT�rq�����`�wN�fq>��G�ќk&�ܶ��-<�Y��5\�zT���S}^w�*87:���g���q��U�Oo���qݧ�v�JCU=��`�W�z��{�y)ƯemU�]�J).�抈[=�u)�sF�=PίE�hƧ�?w����K)�o��.�J�a+�U)t����j�T�!X]m�N��j�'-�d[:p�x,M-,�ܝWC�hw����{�w.�ҙ��hp˭n��\��1�.�J�׽���V�PW�:�'�2,t��REr��͒�3�\����ټ/&�e_U����F����7@��Q�w@M�C�.m��Z�QQ�����/�*۹1y]}]o��'��ck!���ʣ]��"ީn��jea@�mq�����"K���>|�t
��t�߄�;�P�vg�%�Yǈ�9%K�-Q�Q�g����B�0:.��4r����S�	f���w�G�·k@�ym��x��F�#D��^�kF��T�^��GJ�2,ZD�}����Z�Õ���Hժ�H.Ez{���(�m"J˓��/&Ih
�O�s(T���ug�Dx����&Ϯ�W;�Y{�륔X���v�aK�&5J��Vn�C�nL�ݿax�5&��D6�tj�$����{,&ggf������[f�g1V	����h��&D�������ٝ�S:m-�gR�`�x�׊��mdKqF���@F�R�[��땲���8;u������΢0�՝2����Z�dwJO�=�Lu��4vۉm�]���2�YKs��*�c���5r�]jZ19ε�}����ƚŤ�bf&q�:L�v�ռ�l���VCXM��ѷ���H[���Tl��W���q����O�ת 
ٔ�q�6T��i�U��_7ϱĦwJx�4qEP����=�b��t��LAH����n�=�-&�d*���ұ]��1�=��K-�]/�Y� [���R�F]�����<�L������5�쮏���\P��v�X�O�n��arH*kl��]�ur����)�����IYVh�T�y؎��>JU���н�f�A�6��ѝ� V�R��Ҁ��2_`���#,D���zR��f�+wq���l��|ﴮի�m爐z��}i�a���֝�Y3�[�-8(<� ���9Ox��tsh��'�b|<�fv�2&�� ��]Wj �[�٬wQ$Tst.��T{x�R����ui��Z�ho:�;9�qM�%�0��Y�TKH�2��]��;��8ݤ3xu��V,ff�֮��^9 �C2@�=�6����X9�'spT!�gɨ�e㥸:�+�Gb��Ȱv'��>�Fض�wLp
��̳0I�7vh��ӽn�,�}
��v�o>�t<�&�W-����[���Q�A��̹q���:���4%���֙ݢm�B�>�[�u{Gh�oL��T�`���++�%5��Q̰��u�ͧW�hqb�u-�83�۰��������q�$�Qa�X���t�WPX���ċ���I��m�V���	)�{/*$�,e���m�4f��:h����8Ss�YϝZ��Dc 鵚p�L<��P����-�ڴ3Xu�ݘ��AnBp�|x�T�Ҙ���ۖ��j��r�ܠ�E��ݵbwV�{�wA�x@���IQWQN5ݙ��1VKcm�Z@�F+-@d�Ѵb�X�lZ��Ō������Q��6ƴX�#6Ŭh��%�ɬh�E��j-�`�QcDQ����b�F ��E5�j
1V+IQHQPX�6��J���Q��FCX�1���1I��Ŵj-F���[`�>磌2:�I���o�#MP,��Zi:��ffK�4�Z۲+���b�6⿝�[�̅��f�/Up�m:�B�2f�|2lˮ���ǌ�Y����Jy����iΤq�S6��:t��OhWw������S֘MO5#�_�&;[x�K�o���U�f�R���aA�T�G�K;2�]eS�Q{#��x~�ه�ˈ�����p}9H�ܯ���lN�A�>X�!�o�&��"�e\F'�byg*�Ϲ;{қ���l� sw��-S�|}u��,�[�:��_��������^��bt��j.x��ֻn-��(S���%`�v�	����-���[q�8`���Ί}.ک��T��d?��$K+�8�q�ٴx|�=���{��ή쾟*g�x�E�⊎��cθ��v�ޗ{�ۍ��gr�Jm��x[Cq�+��������4�rspN������afb`Gz�u%3��(N�T7��!����b�1���ڝ����m��0�o:���086쎴H�xeKq���V;U���Uaޛ��\y'��y��]�+��-Q���b���G7Y�})�=�Ps���N`�2M�ެp�*g�9ܰlmd�&G�Ť1�,�I�/L��-��#�yK��]6��n��]f��]0H�`��Oɳ��&�7&�{��3��:!MU=us�F�O!bםkb��=��ϒ}�m�*�F!<� u�.��֬�J:�X���|ftZ������Z��g���ȶ���U���x�(��U�yy����ER�:ZƖ�=N$sK"9�Za������LrU}{ʟommt�%�Wat�#)��}=�7���ֻG'ܶw9����-�H�
q�4��]]���V�t���{�#�����\ۈ�W7Ϧ����"_���5���,qk������7��L.��/�Rא����ɥ�]^�$vN(�׹�{aX��,��+,�#N�H]��[QnDRܫ���k�Ȇ)�ɺ
�\G7ե5bچ��O!33�
�鿃Y4�>9=s\�m�,��:��f���J�)��jT/>\��ɨ|�{5���v���߸49e꺈�>� V&��C��z��M,:�B�����"�{;<�̺TR���o)�$`��=��v��ͥ�q��<	�����[7غ9Ma���v��U�,sn���%K$䰣��a}��SS�&P�K�R� ��2�Ә����q��g8V<�Q��#ob)���vڧ|�m�uj�VY����뵎��q\@���;9Yq�ȯ�W��ن�WNG8ة)�5��a�Y�9Z��y �[/��m�O�
�Լ~}Cf��^]'┛B��ogER��g7�*�vr�;J�}q�8�h��Իp6�ږ�5�O9}�kw%�l��r�h�ߐ�D�[C��������U����U�s��9حcv;��w>M���7�m����W���>-ն���%mUQ�
����=ϖ�ds�bq�)���ހ�������Hd�ڠ�Ԯ�L���{O�q�qNV�7���7� ����қڮ7;�R]�wsKuN��A��{�_4VN���[M,��Т�K��"e�'{af��q�2���m��	TN�W]U���bW2V�=�IW��{��xx�`:��Z;����D��$��vv�=8�&`��~����/_y/@�{�2��E��#�ՐP�T	�������X�7vS�w@^�ceov-H���	�I�H��)qw�*�E��{]��x-rŉ|elW����b]ݩ�����OT�9�n�L:]m�J���"V��2�LM��ˡYk6�m�	nr�r����C[�c6x���ɤiWI�a1G�]����Mz���w��Q��T���و`�
W��<+ce�v#�7Q�]������_ǤDV�Sy������uQ����VB�/��ʭ���y�R$G���^p�U2�W����G�gȱ]��{�SFD	�jI�o�]j׺�'�-���3\�x��<��Vq����-O9˜�r���u/q�a%�uK�;�_Cf�ؽs��vN+��E�;��ٯU�k�L��n��x�G��Xa�c��_2�~����~߂�@v|{%�ٻC����s�����͏�ԝ��]��=�ߗ �����x{�֣7��Դ�b��9#_ջF�n�p1B���j\Am��Zʹ�5��p���k�W�9L��Y@'=q��!�������*7O�>������f��㥶�F�uo�\�Å��]��P
]5�N�Z�'�bMwq҃u��]��̵�b,1j�;1d��1.�F�	s��:��Pvl=���o=���b�݉K;�J���m�3����j��1>��X�)�?-i�z�nΌ��.{��^:P�g��������d��ٮM�gg��M0$O�Z��crw��"��O��o������9����/nJ�=j��tt��/��������v�p��\>˂��w��e
�B�Q���e���>喽���(t���^�W���'�a9�X��6�<t�L%�)v�\�J8s�8���ڌ�3ډ�N��Uq��L��u�g��+��3�%�˵X|�lG+�4���vy�G&��}l�zs�J΋�3h]�{`���p�ޥ�dB;%��C�Uk��*��}�67��=�Q�[@�����C\.σا�<��σYp-m��x2
�Jau��u�wK�[�-�j�Q����>0[? D�9��b��Ś�i��S�e ���[uԥ�����n'��:�We�0z�j<��Z�\��h�h�t�%ə�F��ڮʖ�>KX��yX%Q:�ɪ�ej�`1mv�,!�O�����OT!v!�k��	|�Nw*ucU�G6��U�����v�,OLnl��7ճ$W�u3-�5A\c��X���'�#�8�LL�
��/���C�i�ݸךp�nj0���-�N�t��T&A��C%�<�wj�B<$S�ۓ�o��
���F;�P{��{���֧2ě��{fX�zy�[M��I��/G^�x�(�b5;Ӊ������O�m˾�V0�G�m���^�g�U�]s;]�B����ι�r|(��_p2wd�$|�Jz���T���BCT�L�/>C��|�#���d��;�.�c�IX֯�	��n������-*T@��o�Bu����b��B�*=��֫찒�:~�n#Z�x��W�Ʒ�Wd5#a��q7]:��s���F��\A�ܚO'1���r�/�S�Bȑr��F;U�8�_�	TJU�U<���̘[����5���JdvN0>���<�Tm���z"4��^/ݵ��;�7�b;���n�e�1��#���,���K��χ'��r��'�݂�Ggm_�ְո5K�2��U�Y�����D�;2up���-��a݇�j��\n��Өf�:��))��Z�N�lE�����q��}�o'gd������+9��B]Aް�^z�
�/"yo��U��黺�{X���=i�+��j��c�,G;r~��L�Q�GR��-u9㸷���%��LbД�|kO��N�2;>�MW,�澼��a[2��,z�CQ��t8�{/�7o�LG
_jC�c1��3���'��9I�+)�,ٽ�c�Œ3���n���u�j'm���e؇N�R��Q��fr���. bw�ʋ/.q9�#z�<��^�����t'�p�W9L11:�-�Z�����ÿsh�K��R��ڇ��/�?/L�Y��h�Ny^e��9���G��暚��~�:p�nF�]��pV7�c1��e�kS݆#�h��q弃m�A�o����=��^��-�����&�'���[+6d�ѩ��;{MԷ7-���/����Ц�m�� �Q�smrN ��օ�<�_W2&�vۛ�R��爺c6ٳN`]]e���k.��9������[;u�U-U�Ziï�uJ���+'[ڳ1���͇�mq�]gͽ�GSԔ<�G����)hD�m[�V*��߈n��Dj�bwZ܍i��'C��SH\��[j�N��-��z�
�sJ�e��������g�E����C�V����=��mፓ�D#�����y���I_ sԼlu�!q����a
Ѧ=7W��|�c]�k׃ː�KY������'+dto'D��?ɁߩI����'�7�U��Q�[p�{q	ip0z5��O�!�ԧ��@����L�~�Pf$L�%J�=w3��[s��F��u�ᾉ=�����w������C!�֧�;���t�H�����V��
bn&�Y=ٞ0�{���d�W�n|�9��q����}��^�Ͻu�)�.7	��rɑ�*������`z�ᦍ��m�e�N}��Ζ��9�so��ެ��by_J�Wo���<�)����6��� y4n������q�'�k��IL��u��ۿ��2]���(���c��\���gӐM��蠆���i�P����~���
'V���}wKc+{S�O�y.Φ1+�r�y��	�O+�"�ƍ�Χ�CC�4�P��ڥ��9C��� W3b�L�E��Y�6r��<qF ���{�ۙE�x�Bۗ��ō]h�`�W˓�Ǧm�+	���C��b��aF�Cuw��uf�wif�䣫�;V�ZV<��z+�}�t�iz�нq:=�w�/$�ޠ����+i�g��=��X��Hir��;�_w�3����_���J}��&�<��C@��S��g��zkA�'FM�N�|v�u��-���CW��B�C�R����T�ƪs<u<􃞼C�������]p��W֦3�k+E�7c�L�#���.���G��V���������I����ߋ���Gb��g�2/��&�oB�C���k��ɮ�h,���}�nNUk��a<�D��z&�K�+jWu,�;^���[
������/�F}�5��Ajh�n��u�*{�S#�F�	�<���t�[�2��/̭Y��Du�����J����~���rۦ;!��D�����H�Ge�9�ן-�>�)������C~�ȉ~��G���ᑾ���x��s�Ya�2��T�3�aw�{�qམ7��φWp)����%'��,�?�doC�$tx�`��۱���:��u����ǲ�y�5����2��`U�f|�����\ٯ_1��v{���:Y���tk��Y���7�ĸ2���8��0(�jG�w����@%�hݲ&Dr&�e� Y�עr�=�V�:�����q����\��W*v����pu׍�)iz��{$���*s��F�:Ǫ,C��p%��l)��B�X��p��tZ�-�ܑ:�w#��:�� s���{�w�4=|���c�i����h�}~Ѡt�tDҟZw�=9�{��	��0W
��Y�Ԙ��O^��I�j��E#j<o�T������MEE���t?�W:^ty�1:*ظ���IՂ�|��o�����ϻ���~"��/z� �f��.x��+>��/=������gZ�A�cя��cd\Z�b���!�ω�dO��L�!�p�4��ڨc{[�Y��J���N��߾�w�q�N���U���2=�UN�<'���y�u���<�Ђ����<3:�$�gٰ�g��[7����"�ܷ3r[�N�Z�9
����Zb�&��r-w���^C23���ѵ���I�U�:�g|{K���[��Z��1#��ri�{�Y^����������Eţ5�P���e�,[PO��:5�ξw���.r)�V�ު��-�N�p���kW�]����v�d���}&3(!p�6����~ʭ�z���_�<;e#���дz+��̎^/�o��.ߏ�t������~g�J��Exh$���~�h�W��)���t
���B��|/���q�)�g�pS��hͨjo������c��T6�(4�$&p�ޡp.<Q��0e9 ����y�uѻ̥�j\n���ņ�"$۬��7ա�5�so�K6Z.��a\�1�W��:�>y>�Zn��b�%[J���O����j�)]�x�kS���W%M�\_tc�gj����������r�l^;哸'�K�Y�ؤb���9�.��wٶl�ˤҨu]d���R��ތ ҭ꺐��	���Z�]ཱུ������z��;�j�^$an�u}e��;D�ɫWDDe���5+&jK��s�˵�v��ԝ3��;ϸ	�S]F�hA�](aݩWD�n���o�*:�E��M�-���gz�o*��h�O�Y�"��cJ��5 �5k �К�e�+�`w�b ���)3u}�K8�Q��t7�>L]N��\7��U���xru���+����ծd��
�*��t����+��U����ͭ�`+4�F��9�-�ؐǖde�'���1{��G}�I�� ����4X����Y�\To.��6=����a���B���3�`���ZD�ϲ=�].�m;Oή]����{6��wA��Lu`R����}5���d)�mL��Ad�{K��2�V�Fc�q1�j�LW�ۏ�=��h{������b�iRU����@�̺f�r��-�.�=��4a� ɘ�F��r)F��ܨ�7pr��h*��7���y*:��������KG�R.ԉڬ񰦼vI�p�f��|�ͣt�§ko]���-pԚ�w)����нyD8Cyf���j*ͻ`Y`AW}�r�B�G��V1D�d������	���ئ��r���%5N��veX�}�Msxn�ϕqq�/Q"�W���/�;]�k�d9gP���9���٫�TH�V)bΐ>69Iݚ�n�a��8�0!�v��9w��nZ���ٍ��NY6�'}�lsn�WVN�X�uѡ��8:q%��ҳ\��<�E䣕���<xM/]�
W�O���� �,/�ph�<���r�������E8R��y�`�n�����)D�FM���.W.M`v�zA�R�[�b�W!ڎ�b�<Lŵ���K��x%������J�@5X9M�6�`��U*�gF��2��.�]G�v������E�[�83,��=�*�]��[�NGh�\7�{t(8r�m���AE؃��fqb+1q�l:�`	Uo�����M-��.�.�!g wՙ��\Pf@�u��5��yR���; �-��u6�H�¬���iv(U$��G]�Y���\�/��o�b�|>9�-��ŉ�/��cjR����J�!�Y�����������W+/�w�a<а:����F�[��e�&E[��NX��-�ǎ[���)M���ߟ۽zU5�X�Z+F�+Qb��cm�Z*�QEj5lV�[���E��cXۦ�m����\�Ѫ�U9�Q�mb��6*�,[�n-�.-��-�Q��"ص�\�E�b�6�nMch���k�����6�h�7�q���9�j���!sR�f���Ѳ����ʰ��Llwvv��R�V����9{ v��q�MkŖ��;���6��:.�q�ݨ�Zw�]����U�Jq5���{'ԈoԼ��] ^�0_Pc�����9��y;�G�yɶ�,�����KAB�u,���*���˾я���מ1퉫���NS�ܲT_.gN��F@�,uL�?_������b��R�)�~t�����X��F-�O۩��+���:r�Q��LŁ��Ո��DL�<V�s.�+�]Y{�6x_WO�,�bܓ~������=7�������ȑ-W���QV���e���Q���#�h�E���>c=�^�`�޴_���!���fY�i7,pT���>�P���w8M��^x}4�z��p|7F@�{B~������S�p�w�2������T�QӐX��}k�W�}�.��}�{�'�v
�o��'�9��d��A��gζ�z���.|�Kרl��Պ
j�c�h�u���c+����Q��>N�};X���GW�v4��&d�y�^��^2}���nB��P��e��]zEY��f�����nx
l����kEO�����}�t�WJlj蕨�nn�#V*)��R�:O[�_�R�G��uy<)��\��ɸ"k9_E�c�f�D46[�,�+x(���l��g34�5��,����V�ud�CL˗�#��okel�7��@��o6Νce��o�d��`=���Os$�{6�Oz��~��xF{��۽G�}��e{m�	��>��纽�2��=k��cf�����轓��4�S����ᅞ����'�3�uy�x�Em)���J�o� �C�a3��=F�.�YA�N�GH��¶��I�mͽY������W��V;�u�]�3��x�s}O�h�1���a�e��՝]��=�ޏgt�s^�$z++$x��f�s�T�
�jX�w-Nט���~c�=�4~�����}������Ş�}�<!�����ػs69���Ǯ���¹�6i�a�瓻��:�k�z�������W�B0��R��������%|�x<Q���z��US�ü��n�=��1��+���ٿx��P4%w�%*�ٔ�~�U̯R�,{.�}=���m�=y�経�|������7~~��u���7ޚSq�>;8��3�]@R�������}Gݷ=��{��O�e�������xy���~
=U����g���yv� <	Y���e��F�Jǵ{��S)\��r��2��v���.z`K���]�q0�w^�]����~����,K��m���K�O�n+}՜Vv]0�׹�i���Xy�*;��b�{��TD�tqΐ]�T����Pj�􊯨I���zLf5���#ee,܀o�+c�~a�!OAM��^�z٪������ˍ�-G��vvQ�����ZQ����� b�CM��2�[U�65ק�"U��ݚ&���$X�Tou��=�-����z�fZ�u"S��c�p����!����������*��<"�d���$WN��Kf�]ϻ�5���f��������9�r�7�ݸg6��l��4�%�t�z��z���a���Sw�O����TGx}T�h?VӜ�i{��2]���R�j����JWUdp��D}��N���״{Q�-X�p����o��\,����u*��YW���Ez�sh�
k�S���Ng�3����!��Gyj1wbn�7�{�!��y��S+�	UK$��h�Gd��b(<	g�~������V�u3��߳'�׼�z����+� w������wxתW�~���}|�a������?�m�ʭ~��7	�u["7��;��3�J������a�������W��7Ӓ߸Z���4�K��b��_x�1I�[���2`m��و�O�hCP6�ǳ����ϴe��N�!�n�5`��7[�}K{�Z��6��U�\Ч���e�Y#s:����z��VjOp���e�a:+|���*�޼ tKts�6�H�r�:�eY���9�$��V� ��*N�Wt��\r��u� ��)+�C�9��KG�����W��t�7_��Ϥ�<E�
���f��ٞ�f�q�}���xqtNʿ<�{k�3�4�o�ǲW���ô-�>�Y���ʲ�>�2غGo=4�ev�6O�
�S~���E񹰩 ez|��>�*�#�f�lFyx2�6#��af�nҨ�V�=�{��>=ÌTT/u9�X4:^��.�؊�4��e ��9~�dO�G�8 6��	
���^�7ِ&ʿ"CC�TT/_��o��4��Hs�������+��p�gۥ��:kףʲ�#���3��cf������T��&_>��}[ct?�7YTQ�<�
���ҽ�އ��!{&=�~׮g�*�fW{�����@�J�(˞?fؕu*�]�z�:�~)��·��c��{��ȸ��^4A��s>@<��st�/W���W�p�>��MX������d⬞�ej{^�(^�s��v�{}��A�Z���q�2����3"��������~��i�����m��9[7�X�"�p��G�==�|�H��C��j�۽��<@0T�.�����DS�MEE\b�ٿ~�~���-Ӓ���ž���3���I"�n�ɍ"`��}Q��b���L���Nv�P��0�Y�,־�R�xc�ķ5��D��F�.hV���ֱL-�u��.�7���Q��6�)2��:�8������1���h44mC&����Xk���m�������^|7ַ2�q����:��X��Z��Jv{��7�VMn�A��˸x2���V��g��*��r�鶣{�q�����=X�v��zQ�=*zs����تs��Ņ>�w.��U��c��\;�n�V��j�����~>�޷��||cP/�ϧ9PA�*f�C�#�����bd*�އ]�]L�?�T�zq���f}�h������;�cr�L.kzkC�E�R�o��Q[�ϦM�E�Zb��5u��?e)l=���G��9�W~cg>�:ZC�_�ެ�t/c���_m��.��g#��e��@t6��#w� 6�z�ĥ��ԯy۔��]�Yx*N9�u�ٳ�C}V'o�3�N��$Ku�ٻV"�/Z��Cُ�[
�́�!G�W����"��B���O�)Ǯg�Qo���t�ǌ��b�e�eU��}~�!B�m彋���uڅTs��}�v����?7q^�����m��zfY���7�˷j�V��}�{�ݯ�:�YM��n{�t��>a��!�[{���D�7Yo$��@%@��mOw-W�<��wW��79�R�1���8�<p��Noܫ]��i����S�@��ӬTv-*���F\/�M���j����`��N^Sۧ�6`n�wtO!>�ݧ�sE$;��#�O����ᾪ�=A�^ۙg��ר!�޺�.�K�5�y��u�$X�s��b]�ih���o�dJ���d\a�;����ʲ�ϪoN9��9�υm�^,;�ֽ@z3)PZ2���n1{�������["�V�d:�=7�a1so��@�X��/mHTS�2�&�D�9���|4��/����߸�t��:\̫|���rE@�3ُ�)+w[3�T��s���{	���������U44�[p��\3�w��`�Q"��[�Q��u�u�є��f}�{<�xk�c�z�u=�ae�ᵴ�#�_����{#.�=Xؘ�w'ўN�A���3������5����c�_�r�=F,������~m2y��ް/��<���ލui��V�yA�w)��U�w���A��5��5��q�6c��0H�B$X��]�Ii��p1J�G��2Gx9�ۺ~�ۥ,�s&^};^����~c��g��Y0U��P��W~�=Ř���blU!t<��nf�� ~����P��_��*���93���r����9��c;��T�n|�r�q^�f�:G�^W���:駭X�~�b�D�`z�
9FJѼ��cJ;,�Wf��f� wJ�;�W7R�H�vk����cU��0�؛�55��v<J��9L����g �t�"�fה��漇c~"x��.O�pf;!Ի��:g�j�ͷH���p�����ȳX�ßi���a����^����~�_��ܰ��%��6e��
��c͹��o��x{�{k|�G��B�H���~a���ٳ��I~���2��o�>�x�.���]	9�<c�5�U>�Ȑ�h̅��{}�d�#�#�p~����=�J�����ȩ������e3c��ÄNՉ�]᳐=KF�!Nt���dW�Tg�-z��M���s��5��(�9�{�+�/�(44Ѹ|c/�E[W�5�h�A�8���/&�Ȼt���X<�߸��}dzz涏�)�_�ԉ�^� pOס����K��ǘ���ls�|�y>xμ��I�}�f�'�^�����|�˹��{6%z @�ES�����p��m'^�{��ݩ�m�[�O��*��m��O0�s��5���f��b�P#{��T�h�!��.��rv�nog�$�dퟍ��S����=xi�߄�j<���,�G����}{Eǻ8ůe�B�u_��F���e���-F)��95$�fJ�+'��;���c�z�N���\��0꽧�V	��s/��qJ����N;���2f\��2�)�!1��s�_�G��ケ꡺k�ޡZ���z��͵�P�y)�Ҹx�j]]Է�1����l�<�W��騚9lܖ\�l���u� v�}J�tm);�z5�u��vәބ�zA��Ao��;���:��ޑ�{�;8�5�!���=��.��
��r�|����G?a����9
���f[���N��-��c}����*{>��BٓI�3�p�/�Fܘ���=���h4�هfg=�{��y����[�����u�>T���ӿ{���S]W�B���zᕛ�}YIfǪ�^{!����s&��ǲ8z��=��KO��I����n��u3J�WL���'�	WM���<q\Ͼx�Hݦ��S��\>t�����hoz���O��*����b��3ގ�U�ݮ��w靱6&{+��X|��>cq��W��~-��)V���L��r�������Zsr���M�Q>��`뺾� B]�3�\�U���堧z"��:f+��Jh�w��x6�ߟ�^ٻ�;��F$4���@E[�����b�s�l8���}Px�=:�֤9�!ϫ�e��VZ���ٖ�ۙ7���#*����Qo�l*G���0���&&�o�R9fm�g�	J'Oj*e2�M8-�r�)9(W8�u��#������G;F���*�_;=JX$4%Z����ݹ��/����O %3u#�n|:\�����*���6��2������nz'�Am����?z�����{3)���=t�5^���e�u��yw~����f{M�^�}B����ʟ�׮�s�!�OI�d1�@\/W�=J>H��Ǯz��)�[�<9�4G��Ο�og�eo�^קEU�j��[�1��P��*/�y��)����'ę)��gz�{���>���[�����ٽ]~�W�����=��ȏ;�Gl�o*Z�n��_^����zX�o����i�{�]��C�i������'6�A��S;�\Ϩr��d������4�	�%��q�����١��Y�G�u�^��������$TL����I�>�U~y�ޙ]���i�~>>��zQ�ҧ�;�-I̠���s���XS�E��p)��\=�w GO!�d��'�����������1K���j��iR�uo9�Ɍ���͛�o�;#���L�;���K��ȇ�߀O�f�F�p��~�G����(����6�/ۗ���p��Ԇ��3\	�[~����7)K`���O����dJ�1��]��3��	�Uh���b3�n-'�����k��s��!�Xuq�˳8:����I֢K��tJ;��S�&����30ہ�Ӭe�g�n���$u{e:Q�²�/���N�5���Ocu�����n.����7�ؘ��9��rs@��ǒ�V�T���՟&=��3�/.���qN���~�pa p/:�}bU�_{܅�����.�]�;.�O�-�p폕L�G�}�� v:1�-��K{j�\�X3����n�}n�O�h�q��^����HN���~�R{����>,�ɇ�ȟ:�S-�*�d��ކb�f�U���`{�z=U�wlMC𿟒1N�>��ϭHy�2��V%��j��S���G�v�ڵ�c����{&��&���6'���
��	�\i��ឪ�=C!���~ˠ5f����(��h�{��|h!�Cᦍ��t%�Ɩ���[��:��cD�����^�U"j�������q³���// 0ǀ�� �Q�k+p2=;AF��k��'V���цg�����X�+�����uolϱ���7饀K���/tC1�~��"�3"ޘ��9�U�۵ؖ���ϗ{;=;���P���^���3�f�o�CF�ƍ�do��c�Ǹ�V�4_�'݃�7�Q���f�g�g�Z��'�����'�]��X`z��}�O��j�uG��,e�P�Zӂ���
k*�����#[���fc햐]9�Anu$U���U���J�Y�����,u��ә�D�&�-?�<���"��y�{@PN�΅��추��雕k%*X�պ�ڥB�g3��ƥ�.�%@[�2-�|��ۺN�ٌ^�ת���LMu��VU��oqm5�*���>��P)f�BbQ�Sf0>�wn<ɾ&�\�]�})��tmb�'c{���f�,ћ�
�x�2�L.�0��Yۖ/bZs l�Un���"�e辔��Z�Q/z�[�� ���S�՜�9nՂ�䳳�B�̜���-����9B@oCm�u��\	���:jY��Vh�`ed����G9�뇒}�p���!�������u���;��:��l���bl�TN����#5$�WwO��v�҉,ܨlL<u�\�d%�ɔ�v���e4���WX�k왪�?�`̥��`�G�ɻ>�yzm:˩��ŕ�VeY���w�W�����a�(8��A��Vx��Pۈ&mZ�µ���*{��r]Ԯ�3�����n�_!�0�Y����0���#D2�uuug�^g��`�/��}�OB�T'w����h�.�Ġ�X��{eq���9۵@���5X����v�� Gx��ic��*��}��쨧L�W2e�� &~��hm��%u��i�	|��.+gj0mjU��8D9{�\���{��^¶[�E�נCNl�����,nd9c�>�� ���f҂:L�`�efV�r�y�J�mL�)	,;�Ȯr	e��*���+;tLx�rf�u��,TU�n���F'$�q�l��t;���(��X�s��}ov�]�P�t��>��+�2
���J_I��o)��N��ٴl��� ��L�l+Fs���ej�g1U�Z�$P�κ���-+v����͂�cb�쥔�Ŏ^�!7:Jə��p1e���m���/5�驊�W��E$�C�ܩ��Ev�/�0�Ӄx��D{i�@�u�&�6�����w��h�T8%�����ͣ�M�x�"5NP�.�֮�j�"��c�>g���&�r�@�i!mv��kwCp�g�O��P�4��af�&���3�5%@����9J�%��v.���W��n�ۏ�̅)Lrd��!�h�}�x��ùGk��ۀ�8e��>��)k4v��H���
ɷ��|Unb}oL�����ȡ0�}c���;���^0)uo!�Im�M����{IsV�!˾�vqf�ڋ��Y��7x�w�+e�m��@�����$��7	/wi\qV��(DY�j_r��݆�ee>(�Z��W�(̾O$I;7(C�R�y�lNd^�Ի���������wo��}�!U����Qj4QTkj*�Z�j���FKn-�ڊܚ�\W�k��-�V6����Z,q[����sh����ڣ\F����qn
�b�s���i�V-�q����Q��r�m�*�i�6�n-��k�RQ�f֎6���5n.f������""�Ƹ.4W%��W[\Z ���-E�eE\XJ�V��Gۍ���]s����O���sߵ������SL������ֻZ���rf��5��WX �.�.�#�����j0�"ޣk6U�T�IV��5IR����[1���Th��N���O�^>�Ռw?\o]Q���F�g�
�ݾ��u��|'p{����R�*�x�Uo�V���"��gr���~�`����ɋ�	}��dl^R����?Dj�80��u�8ݹ�;���Uk�g������\h�6�<5Q��$������˲�{��vG��F2*�_�<£nf���<�a���̠�:�����Vw_�B����M$;��;�R���vD:�u`t�x�Wj۴�®[W��nH�_f���lfz#����~Y�?[`����Ϸ�gg޿_��U�y%���[�^��5���w6=U��f�ú8��}]�2�q񀅖��.�R�A�o��O��N��߬=�����#8���]W��g��D���T�z��!�љ����b����h� _�x1��kc����^���&|���CLTT/\@T[�����Z7>B��~�<�֏�3��g�E�L�lU����ەN�L��Or*�y~��4.��������ǧw�U��}!�;>G��ʿP<`�x(]З9Z�ϻ���H�㋪r�B�����_x�n��]�o^ڳ��e]&�:�#�e�j2�R�:�*��lk�������=�v�Wp�ݺ��Z��f��9� ��1W`t������$H`.�,���wkj)\_f]����Σ�h�}�U������w��3����z�m_C�f|�~��>��F�M���jA���h��ۗ�!g��v>J-�O{�}�J��}~��6�;7�o�a���0��g�i3闓Bv��b��iexV�sSL�Ȟ�Y��/�j���\\0�
y�ӑwt��Gz�x\{�����Mfޠ�T�o�3 �q9}���<���uӇ:�}�k+cG��Tc.�M�j�dz����-��5��l����)���~�9�xh��z�����8r�B9^�ѬNz�;i���}!g��0\pU\|1{z{���t�<ۋ��5�,�����nr�*�9�7þ�w3�#���lW��Wsʣ*���ܞ�g+����'ڕ��X2��K��B0�Hu�q���b6��V��';��0W�h�ɽR�y�B�w1��^/�}���ߏ�ҍ<*t�~�R�m��>�'^�w��?���ݾ����]~a�T?��M;��R�vo�Ҥ�W�!e����zb{�_���/I�Ŋ}�&��c�j-"���0����1�^�Ǵ;G��S�}y��"~��؉�vAMaIQۢ���;��m&����|ica���V{��69{�R��.U����=鼦O�	�D�]���OJ�78[��;,υ6�:��#����i_v�4�dE�D��8�`�լ	4���R����٘��q۷�(ݯ�H��:�y������ �S�1�	�%���R���`{��!WB�.�`�<� ڴ��E�숞�P��@������/ϟ_��k.mJ�rT���$zϺ�bܓ�c'�G�߇�#�By牁;�v���!��**��*-��F|Cv���z���C�`�3�sн�\�:�
=Ԥ#��/#���g�ԍ��li������j*�֥�����4�<�{��vO�=��齓�φDz�����L���M���H^�����_d��H]���gx�'&��bQU�7�G��S���Aߵ�e`��\�p-�ǌ1�6e�^����گk����_�S��ѯJ1�{/�Wm9�Uz�ό7����<�������W�
<�֛w"r+P����ɪ#�~��ȊcMm�����5�~��;nf��}���3S˽r_�ӥ�{��jG����l����zkt�1[p������z���-�'�X��������y��P���������,�7<�f�Jɭ�%���p�\F^�7��E�`��k��ɸ��W�u]"�Gj�r�p۸l�o�,!���B�5\14�sy5���Yקd������Wׅ�7	������7�)�z�A��̑�X�>s+8��=q,�c�({yV�W��]W}�3��7:�bDx��]�3��_��O��/���o��F=oqON�{6Ԙ̚S�*���9^7t(!ѻ�n՞ʑ��ǜߞ�c*���W�xes&7!?p�������?/k=9�ۤ��[:��?w�'V�o5�>�Y9!���L��y�N�9��o�)z��"w�_�~������[���2;�=���5�=~��x#�3H\V��x�ۙ���R�YuS�������pL�ufN�H��T�&���*\�<cЍS�❋�T�*�Pπl 2W�Ƕ'���U	�X>�Ț��[۾�[�����ap���N@Y�0�>�-��-��Ո��k��R�x��b�R��w*��w�*}O֐�~�RG���>�u;��0�$O�q�����ʨ��Y����{�g�}��	��g!p��f(׸��՗�C��LϷ(����ڠ�&�b��{(Ò�S�h��ˋg���P=:U	�;t�xn��:��x\o��á�g��dB����j�Ӿ��mUv#[��1>�y]C���hi���㞱,���b5��vJ�:݋��ߨ��P�mv~
Ǽ�76�_��j��(o5�����]M�f�V�*��g5Rl�j��]�5>V+9��48v�!�gz�e�|kE���ڮk��(6����)%M��S���j��;"�u�ǰ,vnQ����q��9����j9��Góo�����p�{�R.:ڔw��2��'6�����n;�t�u�F}C�q���G/t3^��z�dU�..}��n���2��7��f�-��If�gкǌ�uя=�>�2�D��饀K�*��{����
���X&?��dfMZ}���
�v ��?O�!z�>����{	���/g��MP�ȿ\Q���f��f��JT1��+�)���陸����W�>����t[�]��c]�假�����?b�I\^��$��z�p���<r�4ki���O~> ���~1�=F/�k���c#���C�l�v7W��+��O�P���J�G������3��u�3n�>�UΔ�} ����Hw�`��E�os�e�F�fr����$W�$q���Ѯ�rr�_�"�ڗ�Es&Z�^�]�F���m�S엫�,)�j��o����e�~�^�6*��AQ��3Qu�x�0��5W�ˀ�u�	�Wt���-�\T��+�㳑�	8�\��^7`�wéwS;3�ڸs8ƃ�nx�g�lR(+A�_�D{�{�<���l{�{��g%��NB���ȑ-��8�Y��W{^��*U�n�SW.�wWVX�hs�O)��ܱ�)p1�"�s[��Ӑ]u�%n@�ӡ����̙й6�X�è��莕�ð���L�(��4��I�E
�����jWxBZ�����vd��z��a�}ѻ�+�@�tɽ�7���hbr���1G�:���s�}W7�RW����"�1G��67����2��Ʀcdǣp��G�8�F�^�
&e�ע�)wU��u�3"C��1u����}|_���3;���sw��U{�Ъ���F�"n]��(48�EB��@[ᓃԴj��/��T�������y���{���Ѿ�>u[�ٖ|�
f�A h64���^)��
5ק�6�U#�ܯb��*бhu'�������w>�ϝ����a�p��jA��~õ�V�+��e�wߢ�ͯϹ��e3�G�'ʇ�G�u���zT����;����'K�'Ӱ=�D�h!��s�[����[�	��a��imi���$~_��ٴ�tp�WL?�y�Ӟwt���bx\{�L{ˬͭb��=�C/�Ui�*��U)ZVק��g�+oh�s�8���o�X@��Ksٜ,u�n+��̻ѝ�T�1/E�ˬ�h?W�N��s�2�B1^��c]N��m9�:�zGO�2�l����mŪ��Wo"K6�{�x����Mp��ɭ�b���T�X�Uo��S8��;» #�D;�=�J�����U6��R�wի���Z���D�X��\vw��ť�sAq*n��K��R�z���ʗ*3���X�a�\�2�Y�I��z��R�҄[L���*�Щ�:�H젨����$��xK맸)��x�BL��׳��aR��v���h��g���=���HA�ɤ���7p�1]94�c�ʎ�[y�b��)��w����~ўt�o���(3jrv�Z���T��A�U�R�a��gfk�}T{R��*g�/xǎRC��0�1ߑ�dp��FG��	o�=�*YT�V�1�I�F���4�u�V�n�(̭�=3~��F�I��Y�aD3�c�>����<;�{��=��7���k��`]{4r��~s~۹��L�'D�-��nl:h���n|�ħ��m�ZB���y���U���̅�7����_�O��a�D�1QPݛV,�g������wq�Nf���uwlle.���~�>���>a^�0w��`I�1p�$48�T/@FE��h
7+��^m^ʼ���w�C���E��
G�_��Ֆ�,��L��%!����m/q�@��8-2�� �\.�@����V�=fa�;�T9״ׁ��^v|2#�뙭0�L����9�<�����^��Ӣs2w�7Nv�ך��7�Q�N��ʭ��=��*|��;�^4A~w3�2��>1��b���л�#�-��
��vt�/����jX���\��}�k9W�i�r���IPW�����rtI�}���՝�w�M���{K����}\���e�R-1z�8�)m.��)���n��ze\Og�Tn!�>��N���\�����o�nӝJ89�����m�~��$�"*۟x�纃,{��&(�%c��y��O�Έ��O㕺<c+f�u�E^�s<O�l��7$\����ޒ�pU���W��!:�
=�fm�.�GzF�Q~�ۇ�^��f��9�ֽ.�=>�Ѩe�Fk;���8�o�s=�S+�����M�Z����XT���6�Jɭ�h<Y��<jG�~���T����L�S��䭐b�\μ�|DvDk��3Տ��<��ҧ�������i�;��I{w��흿aS�::���x�F2�}F"��)��d�� �}�c�O�v����3���uY
�;6����6���O�sީ����b��'�p�2�:���~��ϲ'}oF|�O��u>����ꅗ�λ�Q��~�O]^u��V ������E�/P;����m�όy���w�Ui{��]��ks���hqO��j���)؞<�.�b�l ���[���i�c�W�H������؜�����-��9SIϽ�'}��X�x\3"[��4{Ѿf��������*��2؉��|�p&��GBbJo}�ֳ��V��!��,:ek{/�ҏ�Le��.�|�i�lIs���w��䅊�M�ZT���6��6dqN_���T\%���qׯ�4L�FE��V5AX�a�x�R��y;�z��<xs���@g촇H~����!�G��R�=~���x\3���>�3*�)�k�n����tfj�}2�{�W7�X09�5�>�����z��B�~=3,�{H������0�jVD���+�}C�^���P=>��M[�ѹ!�n�
��	�Q����>	�P�+-]�d�_��������S���h`�s��%�KEN���J�:[ �w�tz:�w�U�w�1T]�ʺ�Gk��u��&�����"(y1F��>��}>�_����C�����-[�<q�v�u��}��<�1#+��ٟd|�]H��M,(9����x�^膵zþ0D#����׈��Ya�H�>��V����a������{�Lܯ`����b*��ɯz��]������i����z���c8���E��c�x�<v�}��������u3㓰����T��Z��ܪ=�b��x��夾q	�o	��D�zv8�����=�/��2-2�Z#0�^V��~Zx}>�����:ϫ�fw!?H��"y�/J�w?fE����o��x(�l ��f�k�o�k��N�"j�Ǭ6��褮75]��@~���no\΢��C�9���	�'�}��y��Ȭð�Ȯ�R~<��tw*+����҅�5-f��\��׮�{x$=���5<�z�[���jU;��z-���:�;}��@0dv�ۙ�5�NUk�V�)w�7��՟�m��{�R��}7�xt�y��h
��{�k�F�RC�*1nf�!�<�T�u��w�"�|�����0�:�!������H\5?_��R�,�dC�v&zg�{=��1]�u#s[Gs�׬z.|�_��x��������ǯ��^������?9YaGA�<ڶ��^�yegwx�U׀3=�o�����#)��}pE�b���C�����LM 5��Th�3��m�����g��A��2����9vU��@�r�n�?�bF,�6Vz�.��f	+ ^!s�}i���π��#��B�����v�P���5�1�+��Z7!
s��C��oo���u���+�_��|]G����ؔa�LU���A b�CM����m��yt]䫘P{ܲ����GOd5f�I�������mr�tϣ�̉~��(��]C�N|�HT٭�Y�]��1��^���������ߤ�����s>X�L���FW~�x�W��/����[�27X�+��ͧ$�2��M��s�D6LF�=���E�[�gj�uʢ&]wU��|3yb�<^(uk���̫ <�X.G�Dވ^*SFPW:�GH`��өe͎�5���w���3T�%�nt�)��eb/îe2�n��䊫`]��[�)5;R�)оb�`��s^��4̧���+���t�W8C��,Z��J	*��͖�-a:͕�� Kql��[��z5	�5NҦ�J�J�}�\^%z��R�1�q�z�R�n�mý���l�<{t�&̮�k3ZT��/%omFV�#�;pj��^��S�LˡrR�s��c�������:�G2����u{M����C_Yհ������Vk�������]�ǒ-��&�7ʦ�o	뼜�z�f�ς�!��Naژ2TYR���c]�3�i�q9��ݝ��!�����Q��:���"Q�4k�yݠ��v��H��������uV�u-7#�t6��sx�:��e�Ů�W�ܨ�)rv�I�����K��؆um��]���:t/:��w�T��&�4B-8�*�8�u���.�W�J��!�b}�]
�&�[�r�V1q��HQ� �I�*��u�̻g�7���E�(F7�e���J�>PL]�0^j��V򈭫�c{Ho,�%����^a����v $� qYv#���Q)��Ռ�Zn��J/�_^�)RՂ���	��W�����R�Ŏ.�	�
�!ġG7�D�}ov��e�rB�s ̩ם2�-�ljvdv�{ <34qUa�9Rg"�F�f�j�5�.�U��M�W��]�q}��zS1֞��p����G.�A�Br�#ؐ.֭�.r��خ�>�gu�AwWE])V<.�R8,���W�a�ɗ��u�FBX����r�R�|�U�)��:�C.s�7�u�0�5�G0�coiF+q�륥4a�*d�W9r��7Ք��4�����D�b���1_e��DtU���v݀e�V��[{`�S6�D뮋Vt�t�����c�@��Ka7�6���#W���C��\�c�s��Mk:_>�yz���8f��5��{q�����ox�ܺ$���"फ����ϹbI jmu��T`��*��7h�E������,)�CᥬN�z�v`����7��gp�:�0�K��w̎qk����Q�H�3'<����t8����L�"�(�r�p���u�s�	a����@�av�s��W���tc[@�g~�Y����k�]"J�ʽPeeo���6�vR%r��?Wb鷵�9���Cw��ޣ�VWU�ǚ�Q�ײ�G�6aO�5����OV^:�G����m�	�5(�j9�=���;��	D����nV.�k�Ċ�C}ɂ�;U� V��n���vv�%\�6���#�C���2�=��.�LJZy�Y�D�8*OCK����D1������m�eǂHj� �������)�8h��m�Dޖ��w��������>�_y��8��*�&���Ɗ���Wh���Mb�M�Ƹ�W�����%b���؊.8"ت�9����q��m���уE\T[�8ƍ�q�5Ÿs�F�P�#Ü�Cs�\q��rV�mjL&�Ecs�(�L�Y�k��Ÿ��+���667�Q��qW&�j�q��n�m�8�V� ��.6�NN�Ѭ�9�lj�MF��m�qW9�̬Ibۍ�m����m\Z�q�����8+�U��T�kq\[r�5qq%�1l�*;���ι����^����}���5v�u�F0d�2�̷q��j�s�Gu���k��M�\�t]f�o#yn�h�����:��ȇjQV�+���lm�?�7�
{���f�f���o=;��x!�q�{��b�+rv⃏mPL*{�B��%��d�ES�h��d��Y}GC�uQ��s7�=����G���|}^=�>h�T�3��zX�o�sdXg�X%/ˆJ���姇��
����}]���v���UM�w���\�F4w�H���xrU�k�\ ��kt��yeۜ�Z�Uo�{ޭ��;��+c��/fo�w}��<���%�{���{<_����q� �fM$Px���Fvq��2}^���#�}� �̋y��F���|��u��3���.zs�)�(�MrW�x�<�v��ω�Ν��W�1�����0�/��0�3�w�c�=~ў�l%�J�Os[���#�I�=�R����;�<�y��u��Tlzf���)0��3HߞEb��{�x.ݔϽ��3}�+q+^7�Cѷ��!�[$L�'��-��nl:hN|����#�w�S�J-�l[�I������1sgj��S�^�Řy�Xs��5ٵb� ^��8�O�,V\Ҍ�	-�f��Ԗ�����-o��T�3��ˎ���:n�V
}�Q��\d'�9�7�<$�c����.��-<OX�8�T�@����[�t 3c*)}2�T�����C����jqv�S5ʝn$/�8�!��;<�\�u.���UwoGe-�=�.*o�֘s�8*x���d�-��?Hhi��^4�������ϧ	��g���&�������p=Ϙ�O�C���EyY���e�>��L�_��~��N��ctD֏˝_�u�:����*DSu�=���*��O�Y=�φG�����[3)�=��{�_5�=}�&���d߫��R��(ʞ1�%Yw�.3i���A�N��C^4A~w3��oTLt��d�y��V������8W�p?Q�(���9��tUlj�>-�dz��ޚ{�l��.�%��E�yWQ�o�p/�fG��#c���є<ƚ���1��<c+f�u�EI��n�:EL����<kt/dϟodzqֲ�gz�ǻ,͟{Mh�ޚ�(44��<?e����o�V��g&�%�
��њ&sNۙ�b��Br=��^��1�Mɇ�7�VMn�A��ka '��|Udy޷��ǡX�q�3��?V��ב�����^>>�V��}{.����Ȏ��S�i��5�3{ܠݎ��O���VNUJ�o؉�ʭ����2�������?�|cx{�׮�׎L�;b��ͼ��,�ݩ��ԫ��<���vr��*Y��{�=;` r!v�֖;�
��i�g!<[�WQ����X�8;ɒ[Ϋ�@4�S;�Z̋V#�Ay�}�5s��&�o��ct�
��w-�i�,�k#ȱ�L���[�j��=h�-�5IE���G�n�YS4�S�#�ۙ��0�۷iק�?]�2�S�hE�H^ ��V7`�b����a���T�4����6�i���U9��뗨�R�/M�����l����w�Z�k��*0k>�t�\1����;��D��b;S�c�g��������R:o�p�����W�c3�O��*T�Μ���������}��"1q辰���z��> �K��k�m��=:�@A�D>0v���~��|���?u���>,ԗ��n����l�6���{�o{:���UL��§��������/���/"������#�vfZ��݁}��}rt�iq��g�6�� ��P�ʱ5�nH~�Px9?�0���g=%E{=]���I��ݙ�NUoh}�x2����̢������z��T44]9��X�B�S���=��Ι��UVx��}j�=�c�z��U���k��}p�XlǀxP�~�pш�;,������R^#'�	�J�����������w��GQ�=�>�2�D�w��/��^�v�%oA�<�y� ���e��ͯ�3k�R�y���[�N�l+M�t.�������u���LV����udD_u�f��e��m):f��Q���rXnJE�*�S�(d�(��5�1P�iob4r�m���$��""ŝ�Z{ݙ(�<��w/ˍ?��F��U�*9Ns����e{I����o�A��R��kٙ~G��jOl��>j�n�;�ٷzh��Q���g����8w�'G�����}�]�y����!�>�eb�� 4zN�����#F"������j�=��~ �ǆg��7K��p�ޖ۵y���od^,��ae&����p��i���K?*���w����Ɯ��}3UT"z�9��W�1܏BW��K��~������1� Hu�8�v�h�x99U��0ֹ߫X�����p�K5gez�+"{��t�yט�~
�F4���xB?lU '�mۙ��bڿu�&�w�ݹ��^48Dh�	��?1^���;�;9餇?W�]�R���v}��V�����v��̻^�>ɓ~��S__+@d�/�\<��}/���s�k~��ٿx��l�Z���i��q������ٞU��s-ґ����uF �H�w�ϟ� ���e/G���n�\yO�Ś���a�H�o��P�*�e� v$9Z3[���q{�$+wWKe�s�����襛��c k-�<
�;�h���l�v]��0���?+S�e�X'�����w%��R����ub�jbڜ4Մ�%��2���Me�V��
��Z�e�>�AW]���8��nU�.��SyVjSB���7C�,w%[ًV��Ԫx�ƌ�͢�n~��V�~��ȍ7�<�vA��ꊅ�hc�2v�h���=A���.s�lrq����G�V'����e��^��+�~܊�y~��?Phh��ۗ�!?og����W�3c���cP������n�����dz�Ϻ�)����R&�{�ԃU�5%����0q��B�r>���S[Ɨl���_;���}��r=�`�y�ϼ]a3��f��L��uS�g���/elǅ���zE��nT>Ϳp1��gL?	�Ny��2;�'���ȿP��o����~����Z���J�ki�xzr����U��b��ǵ��H���ē���mw{,0=T����kAC�v����?�����}�C?%�5��U���_C��L��ϳ�F;�:F?^�>Z�^�����
(<Yv�0V�>˃���v.��+�����z)$fyj�׵�+5��Aw��G��O�PB餀�@�}��&W�Y�i�Z��ϡ����Uoz�/M��
v#1�և����W��S§e�E)�����O�䫄�i���'t8{��Ε��a�g��%�Ewjs��M�V�M��DF�}ת�q�]t�z��:*P����wpj�ŴN�a���4Ĺ���z�9R���m��qs{q������PrZ�2.эQ8��߉���-i��Mw�n�iݵ�{o�9&�C':��q隋�a��L7�p�/#�����Ka��s��S��(��e���}�`ݽ�Ruc��eZ�`V����Xs5m�H9I���i��9�C�~�����Eѓ�ܣw�zǻ�z<�.�^x�r!VXa䉖Ŏ��F�nn��1���n}�������C�s��v�ٿsk=�"��	�__���{9N��b[@��F���:�����Xs����8O��=W�g�k.l�W��S��h:�u	�&�<�FHhq��^}ج\�����Z�+����}�>گ.��}q֐����g�β܆���e��0/<w��[��W�����a���7������e������</���8?~9�ʞ^���C���w3���fS���^�ʮ�9��^�o�@C�}�u�W�i�F\�m	\}{B�C����mw5�]X�WO�FFY+F�
�{��P��p�k��p�`|^���NVmd���
��z�5S�#	K�t��Q�4�.R�a+[;�-����A֬p>���c.�~��<
(y�5���c6�|b2�oE��d=7�>�z0����{���u|vp��E��!��ֈ�2���a���<�.f�lZ�X�ȁW�m�I���	$,�\�%
�Y�k���-��CJ#� Z\�_뫷���pڜZ�Q�dX�J�*�����&�ƌ�c_}ۻ<���gfo��=;��T��K
=�fl�i�c�5���ۇ��1�>���m�ˌ��g���5���P���Y~�9�����{<~�Ҧ��Md��&�F]�y@V�j&g�c$f3��n}�^UB#�e��8��5��u�s>";>����^�%��z�ɕ=5[�u>��{f�mY�F�A��e4�)��bǧخ����z�`��;������~��Z����q�Vsu��~�CѾ�zs�� �6��Ҥvݹ�=���Iק~K�gϥ�dš�εN�[�}hz���~ʮ���u�;���֠7�o�*���#-p��^���c�^R��^��L��ؿ!����H�'�������=}Xb8Êl���"?#��D��=�;p���������D��}5=~e�yM$;=�'n=��L��jD�Z\!�[�eG8𚮍Q��c��S잿}w�"Ǖ�C���$[���~���!�i�}j�g�&%]��G�S��|7��B�D�}\�cJ����&Z����0�ي5�/�#�ރ�;�]/�]C젿���������g������X��n�1���e�
��Yچݱ�s�Y��N�W�N���>T������]M��Gy<��x1u;o��^E��p,��]W��/����їo�Y�4�����ycw���V��&ѹۅ^L9��7���="me߭PȪr����U��;Fl��3��)�Q��>�y��~�q����z�b����U�@�S*߰�+�"�����lg�K�KEN���Y��z�=ޟm�cݯQ��c���C��Rw[>,e��/W�-�P�b��Y[������Q�{h�#�W����["�n}pݚ��6�{#��{�{�fi�'�#��`��3���A˙ל9f�'�oD3���WH�����+��yz�>��޹��������ٿ|q3�t����l�h`$3շ�q�ǌFmރ�Qβ�d��g�dxk��dOv�"kR>��'���]�9Y>�Pѧ�Nx�i�em���Z hs9�����~>���B�=ooǪ(�G��!��ܾ��a��x� b<�Jr��E�u�3^V�o��V�KK?T�r�cf7+��x�~��.Ko�;��G�27����G���y"8���`��;��/\�i��~~w��fk��[���jVWx�y��y���^C_����Q�~ۯ�H] ������ۿtS��QA]�J��>�����W'���1��b��Jh���l�V���)�/N�&�b���N�y���yi��u�}��W��Ks��t�J�%�)����X+%�/zۧ�w Y�����3�]��ȵ��NޡS%o�3;�����4�O�g����ש��C�u~��?��4-��;����;R��X�[�9�UC�+���3��U#���� fW�����Z%x<{p87���~��{��+�|fvm�ͭ��G']���~SyU,8�J�̷U�S-Ґ�)����@c��^�ḳ'vrX�����]I��Gp�w��K�㳟z���2ӣP�*�o���fG�����n�mgi��I�kc-�t��OU�/�z|�}��ϟ�pg=�M�˷a� B��5n��e�&�b�/F��h�����&5HS��.W������ת��]l�/ۑW/�(44����-hE�����y�:p�Kc��g+��Ѱ����g��������>�[3��xR&�{�ԇ]��z����Ֆz}�X�����#�#������zOə�I�2i��:���2g��g�f�j���{x��C�}ȡ��^�����p�m����
���dߧ�����G�h���fՙ������עP�w���D!�Xs���X6����d�5��t?�{ȉ�4>W0�ܑ'�rd[�uNmI��1m�lN.x6k40���
lM���vI�ԥ�W%��9�T�o�S��Wl�>4�f;�!%�T[[6�Eks��ˀ�v�� X-hZ;��-h���W�t5��ɜ��'E��2���h��I̔3�'*��j�����ƃθ�^F�)��xt�����Ul���M�h����/�XFZ��o��;����b�zA�w�#�x-F/^]p���[����.�㛳}�K�N�����*�cgʩ�kU��ϣ���f���������g��O�u����G�;�	_�3�:H�j-_�z���rr�|=[w	��^�����do��~�N�,*vG���v�NV�?�ъb�]��q��?U~Ajh��R���+�x���xz)��p��FG��	vF͌��QN;>Rb��.}]�����LvC��W�g�F,9��l�A���?=�4�o<�=~�����]�z;���qۧx= g���X:=e�L�C�3-:�yW��"��9N|���[S����	�|�XKo�s�>��~-�ȏ)V��	��Řw���O�cDoM�=����b�n���=���Q�{��u�7���b*l�ex9�{m�V}k'V}�`O�:���_��v�G�Ĝg޲�u�"���р$7r�i�Cg�հ]������~�]?ݭ�UW�+j�m��[j�ۛVڵ�����km�[j���Z�V���kmZ��Vڵ���խ���m�[o�j�V���kmZ����km歵km�[j���kmZ����km�-m�[o����m���ڵ���խ����V��ֶխ���PVI��_�z�������@���y�d���Z��s�	RRJTR��E@�J�*�!T$D$�T�ER��  �U@P���օ
��
�	)QH�(�*"��J���%%��\l�TU�t�UQRR
*(PD�a�(�)4ґ(R��(U ��IH��p ���!��h�Va��Q���[E,�l�@3e�h�5��*� �fh���J�r�  ��� 6� 
 Ղ�(�֦��(4c	P�h
UL� ��6HXf�V[Pm0��M6���iX 
�`���
EU� �ئҶF��Z�	k��l4ڙRj�Rk,�Skmm��%��"UZe �p mn�J�����i���M�Mk
՚��-�,���D��mZ�T�dP��JU����6����� ���hf�SaUm+a��jL������J�J٫mj�V�eZ��kE�V��-T(��T
� ��ѳ4ʵ*�,���[ma	B�4�jfl6��V�)��*��b���[5YR�"@�G ��U�VA�ԕ-T��1��c&��j�ڶ�֑-�����U�������hLȁ*�!BRQ� �Q�
V@j[V��3ALQ��� BQ�Z��Ȉ���SZk�ۅ
�`��X
�V�4Z� �XM�Q�J���`ޕ  
� &)@&� 2  )�IQU���   ��L� �LL&4��)� �"� 2h     D�	���`�Ђl��z���2A&�C"�&Q��`h�L##��2�o����w߅�U���vk^[M��_J�Z�!@��I�@�~�2\ ��;�D
 ���I1$�Q D*Ƨ������%�nLP�`2� a�
�!	$��2���|�� �d$�;Hq�mӕj�ӯ�V����"�]�,
��(���x�#STe#G�p��!�w�����h���H��o�����_�����ܼ���Qt�V�p��VAɷ�=Q,��]\�T���E!ef���ݐ���ɲ�3^-x��r|t[ =j�j�~wgZ'Q�CQ����LL��L@��`���A�kZ��S��.��ә#n��{jӨ�(��d�I���L�0m�t����*[Ykȣ��="��`�U��y)�'f餰|wid�� C��Ǣ�\�v ���iB%��쀶��Vf�6�F#�������@ܡj��`<ae��lK��_10�yQB�nұ��z�4&�8Iz��r3a��F�`�i�7�.�Z
T��6dX�"1*��*��N��!��WL�J�Qɘ�"�rl�7N��2e]��)��;:*^7���� ōD�H@�Q��Y[gC"T��Ӫ��M����1�aһܩ*1�;S*s�P��H(��J-2�W��^K���8���*��<��)����.�����ͧww Ut�T63N�iQ�\��ݶ�T5�� �{�Ҩ��P��+Н��up���%1W�Y���JQ��R�d.Tx+ �]鬗���q,���hj�2X��
�i��E�F�yMЂݧ�2�	U���jUzت	�[i���.�� �Z3-�*��h�M�n�E�2Y�2��ocԭA�Q��S���gTr�-�i�.�/J��`M���O2��;��R��֢���OA���
Z�A��2�ۭ���%�g�+e-a
K�bYd�`�,���6�en������{[�E�c�r�R��N�Kv��eBŌť����ǻ�!Q ��b��,�H��c��^F��{��9&b�M�%(L����3��j�#Q;l�2��H��`#ZM���^\r�=�Q�ꅹ��b�l{��T�m��d:�STY�l`�Kk/>�"�1L�ٰ/��Q)Y.í��f���5�!��Ը�D �wI-��7*h7X���7�a�/s(bv	�&m�q7���7bƫ#*]z2fP#"��hTG]$N�٢�	Q�rX�,�	U��K	͊����� !Z�[ceZ����1�67+t*B8��]C1��fQb{��7c@̰�t,h� ,��E�Xk/pB�c�:&��t:ݚ��3�윴���}�%b��y������ƅY)�ڹWf�)~�l�T�A�U�h��\A�y��h�ܭm�3o���]&�6B�KA�Ys)�)d�(��e�ԋ>n�wX.��Z&nf��[#۸Hw��:��2�"�+LNf���V��X���j�7P%�jR�g2Ш�R6�Ua\6�o*�*�d�Uo(j�[M-��i!�%�d#0K-V�h���F+���^M����죚C2��$V2΀��{��Ł�F8Ú(��Y��7��oE�\��FT�,d9���Ki�b33qDkmԣ�eC��H	�K7�"���M��Jr1�B�ѣ��^b�
���g>/RӐPgjb*���[���$�ӫp+8�<��J_:�J�3m}DU!���[�lS�l�3)��'��^0�	G`"�ތ��VZ���e��w�:�b/1��扚b* ¾�i���Ȕ�%�e���V6�1���uj����X���69A�V�5���Q��������)�^�W��)����q��a�A`-�\!�0e	)-�m$ik�a�wd�0�[��'ɉ^�e����E�D�ota]fVlL٠Rt���,U�u>h���W��ʆ�15�"3Q�e*ǌc����i�53�5.���2ސ#m��eff,6ٚYl�x���&B�-5�ܷA��V�w��a����ͶE'Wq踎8T�u�kD��xǮҡ��4Y�9�Lr��J�2(�o.�*U)��XpV�9���)����h���(Sw
�An��!+k9mKP��逨���j��)����iN�uـe�+&��v��&ݫ��!L�ysC�c�d3�B��+V�zj�t6�(��M����!I�3$�U���ؕA��9�T�o.k��6葃 �0#��J��
l��.�|i;�}*�A�RR�n��`�cA��jJsb`�B��\��Hj�e�iڔl��Y���0��eV9l���f%��-J�4�u���Y�SD�w57��W�se�v�NV�Ր0�O/�w�q�̑)���ˣG(�ں��e� x$�d��i&j�KFe�O��.�-�<�ˠ-��٘#hțMG�����4imi� �j��oj��`�̲���/2�f��R-7-:@}�,Ն)��q;��چ(�F�3N�0y�l	6��P�M)��YF�%���b�ӆ*�*��&+�#1��f�A�L{[A�ے�u��$��$�[J	D�C%�3r��d�NRb�L�#`��(�³Z1e)���!�T�3sͼV�Q8.�1���Z��e'�,!����		�A�O%"7vU�l�w�]�+2OXʭr^`ȁ�>بAd̨nb;��m۹B�si���M�Y�$Ѫd^1�K� rMSi-��NV�cDA%��]�h��1I�R�5�@K���9��͓p4PL�"����VFH�v�	�Ϯ��R�����&An`��[���^p��n�ٵkuyt���E�ө먴br��L�b��wn$�4̫q�l^�I�t�9�)0�E	a+5�,B�3c�z�n�1�m���i�ub`8�`\	[��qh6�^�F�ͺ(�C@��
�V�*��ic�f�'� �m���e��)��-^S��5�v��J���`�2F$��t][V�Ig�~��J�6�P��i�H*WV�dz�ěE�h��[ZX%d42e$[j�@�(j�4�	-p�ܻؽ�X]]��+H��̗�o*�TgQ����&��B�y�i�l�X��F���,�¢�fU�q;�:�E���o�(R�79-v5Ч����l��u�Fm�%܇U]K˨���Oq�FRq�{M�$ 6�^���u�Z5��[Wh��r��m�b��s��t�����#9�'��d!����{�F9a����`��J�2`�&�щ"&��R���7R��ӹ��4�^�]� P馅fʖl�Z��Xl�� 	��^JF�Q��E�M#8����t�6[u�{�b$E�s�x*g8e^�����o 8�����Yq̔�,�z��VFJv���1d��(�&�m1��Z���4�ێfT�V�T�ЕB��eo��ot�.ݺb��rά�b�6�iݽXݚ�r�@R����l���d`Tkq1L��͘���m:����7�t�7�	1�[$іJܳ��>b���y� ̽��R��[�hF�SR%�N��NM�j��#i֭�D��q�oP*ЅQ�_1H�2��7o��z5�@h�R��
��aؕc*VZ����8Sլ�́����W/5���אZ�d*���Ѐ{nCx�X}.
4�$�i}��:f���cc����x�;Yi`
�YC���l���d^���sN�9 ջ����H��X�0�Vt��x
Gm٧e�$��m4��6j��ZaLcWei`H�˱�����Z �p�kn�a�a+t���zh�JY�v��
�	���x��ð=�5(�FU�LPʃ(�[�c	�úM��IQ0���Ś��][Y(Dsc��!x�4UCNf��&��+6i���:`����,#P���Jpѭ:,f�m�W���K��(\�� �Il�c9#$�h�2�#�vU��Y].��Րr޹��PY�!�����,&ŵ�+]�� ��;��������7f��"�1���)r`�gA,S�X�����C4fJ�3஭f�uh���t��s�I�"�ܒ���K�I9@�K�wl�	��J��4�AO)���R�CUɘbC���86AQ �w���2n�ee��<�����~��R�ؽ �5��)�Cx'�g�`Y�:K\B�ݡ�om����F(#8�;r��`<W�f)��Ɩk�%h���k�h�vfY�EFeb�h�9�g9b��fP
�� uJ����6��X�Z®ZZ س(`6�颛N�a
fp�.���⭼8����TY���Bn$�<%�Ů9&,���mկ�������L����5T#�L*�zB�G��^�S<��Su�S����Ru��,�#r��>�<������gxVo<�[)�m�4J�U��p���L�KB�Kꝶ�t�Vj�pP̶���s�C�S�em��J�$��`x�r�un�7��X4)���������T{y�Kk�Z3�8�2)��Ы�Ob��sZ�R;Oc��l��c)�k�]O1�e�U��4S|NM,�V�fS��+J�w��b�1p��B��4����b��Ә{q�dB���|N�����38�.�+���L��X]�ŷJ�.���N�{@�
����'i���o����έ�`!�KN	θ��̠�gDB�u�"������Ǜ�1ۺ	�f��S��|��k���e>����p���-|���[	��5��aLc㜰�x~"XY��}ff7�)�j:��1Z;�J�;P'{F0N�k7��c��Q��ܡ�qٷ��[Spl)��U���T�s}�h�)c�����9��>�E3�ꚮ�(	X�Wn���z���tc%f뼫H���)�or��n�<	>�t>2���U@q��OV+�f\���%�_%�sF�!ÝHB�0�2�^���VEֳ�૝;�V&�������cbF��UF��W�_Z�n�;���%g.@M���wDJ�>�8)�2[���
�㗢��ʎ�,6y���^T�җR�"3[�E��z����M"�|';��nl�L\ι��4�ME�n"�u�#�8�6q]�FV�4�pjw\�s�Δ�.�[����Q�����U�o�X�x��A��Y��9WZu�b|��/:ZUcK&�Hr�:�Q���!'p>];��歁�V�i�Koo��$�[:�)�W�d�r�h]�nh���p�4R�Y\�U֭���与�W\S5�����7۷�_#}���� b�\��N����6bv�Iʳ������V�Z{5�7�d��k��V6Q8q�4,�����1<�� �NW��+Z��5u'�K�B�̷�u�;V�^��ײt�S���L�7
��>���g��y��1f<�ԓ��?q��6�r���(�y!V�bL�Y���h�jֹwI�y5c��,o'L�R��q✎���˳w]��T;�PYʡ���#���K�Qʓ�����hWWL�6*j�7�qHkk.��v�Y����U�0:���:,���xj���]'����D�� m�I���N���_ӏӻ��N6m�U!�+m��4�䬗&n��n��u�oO��%��W�ïg]�Ѝj��rZ�ks	�����uѼYV�_TU}]�����"�A.ٵ7tb�q���݂V&���JR/��,1 ���n�!l'�cwiӭ�¤�3e|n���գF�]qH\T��"���m�Ø�zh��cR�P�tcHf�����λ�S�"7��*�)͌�KoB�/�@���wna����uo.�TuW5fq<�K�Z�cs���~���o7������̓z>����x��-�CV�$����1��1گ3��!�V��=3����I���f��i�f��K�Ջ�fj� �:l-�2��b�P�4f:W�[zS���"���R���R����3�a��wD�w���m�Wd��҅�ٕ�V��5�f�-Н��{�
��g
e%Z�n5��+iF��e 1���� xTu-�z�l�2�!��v�|� �Mu��T�R���l��&^�a�V�,'U@d�eQolD���*Ӹ-��}���(4"`_v�V(R��dZ%�]E"L�[�,�wln�I��$a��K�w �J���6�C5���*����N�F�D���LKM�d��n	`K�D㓆�-Q饡}�P$β1;��i�P��7����L�'�[���Ӫ�xB��T�~#6[wNhc[���u����귓�V>xj���g u��ΥIk�y�W�^�	�j��<ݢi�2��dw��*�`Q���vn��!�/8�yvx[���z��L��5C0l��F·�46R�{]Eك�G��'��dM���W��UP[��qt��Cʳ���\-���N(�U���|(�|A�w�pY�/��ՅP���P�z�ۍ�k%`�Kl)[AD�c�w%-Y[�*����S]��7���}���vH�0Gy�K��c��!Oo�v��`E�t]�m����8$���Q�1!��"E"7��R�4�݈�i�����u��wA�����Y�>���\�LZ�*��w�4!����u�dY�@���nbg���&�;*�6����U�b��\УKC=��n�*mpk1-���fl��Ǧ�>`��2g��(Et�̷e(������277T��՛���)0��k�U���4�h[��aS�M�WhL@�CA�H���x��g�2�cS���z��\������N��w��G���k��j�f�+����̗��5,\]���5u5n◼�#NkEeJ]W`���wˌMr�up�Me�.�j���̸��@�|u��ӳɹ*�w�T`ӭ��Wŉ�)5���=�%�e�IՄ����ujX.=�S��7�M�5)wm�7\L7�5��FFv�P����k�z6�f=�p�|�M�vQ&�v���ȩ�ѫf�����ʼ�%ʵ2��j�<�l+��#o��ЧW��_Wi-�R��vc��l�(�(:7ñP�v�Z��V)PX����
q;s��սӷf�ٱ֬�HH67*C�U7£:[�%XGU̧s�O�T�5�|8�d�}%���0hr����Z�=2�s��.P,�<��j.1�:���2�z;�p�l ��<%�/��;˼V3�����#�r����K���-��b2R�Z�p�5���{|2�ty�c:K�2ͱM�ۃ�k7R�7ر�+�L�|���C��Y��G]1Ǹc�Mf� ���V�h��|}�r~^2�F�B�e��u�����N��:M޽�����u|�)�E���u8� �3��0��n�^�h�]�."���%���3���B����9�k���I�ٝ8nh^��vO\f�d,՜�O���#����h����fM�FW<]�S c�MI0t@��)V�6�Y�:��hi��b�Y�
5��Ӫ��r��)�n]�>5u�XݱT�q,����`Ӡc�˖)mk� r��p���M��җ�˸�!��Gj���/�r�m�n��#۷���7Lc��JX���U:`��ź6d���Z�������'H�o$�#�9��i(�1R�77����"��?Y�ґ}�lh����RQjxr9�N�C	�Oy�\��G��C���ӝ0�� L}G�5u�;)Y\�c���~�dKU���Ŷ򶋖���3]���OU+n9>e=�GV)���s�c���xQ�؇���/os�ݽł$��v���� �-�nPQ�%����"�H�ξ�b���C���٧ �N ��zp�'[��H�1�O=ꣵ�F��\�;�ۍ����ܲ�m��@[�3�����:�ڬut))f,� =xh���_w0��,|.�N�;���.�Y�ȉ3#sv�^�4+� �V!⭔pElV]��e �����1R"ia�7��-ޮ Rⲷ�6�� ��W�Mn��wmMP�驰�� ��uHʨM���!髆�w"��͂0�S�9.	8���!��a�3�p.u�MVc��Iow�.�]gP�� ��W��+S��G�%�mvj�פ-���n�L�|{vuT��g,�������0��7����q�]J�G�1��Sr�[������r�|�|ю�/��3��|leˌ�wn��>"&w��]�]�jc�L֭Y:�јc�� ��}:p<��p�ו��f��g�����ӗN�kS�U��;K���K�r�_^W�[K�%�&�������VA($Q�QC��,�ʊ�K-v#�.�$�)$�I$�I$�H��I"�I)�s�HJ'/RKh���QRWb�j&��+yD^�&�϶�F9d7�5��Zة.y����*�H��YG;zZ��w�[]��#��SAB��J�b��������@�B�v^�%a���8���u��EV;�ƻE�d��z��uo�ڸ Z&�q�}E|>��%ۚ�4T���P�oN�|OP�!.h`v�{*6%.�C\��,��UhL��ed��j�����cV�;���t�:C�Ű囤�v��i~�i� 
d�R�j��!���*��� �$;�� �w��el4�;6p���.�ᅯ�����a|���G5vŚ�9;�.mr \���&]�w��"�4 ޾�Ҕ���5����H�P����q�l��n2M���qK��9ҍ����+0蕻g�G�՗[��J��n홃���蔾�uk����:�N����S�+��uN�
�3@ۜn��ر��]ۮ_C���4ΚL�:8�,X��;cVF-V� (m���I��@������d�7�Z"��L���5��4b��*ٓ;:Wp9��w(w%Hn��ۭ�<h�
�kY	�7�u��n�z��04�L�|Sl�z�]�\R����¦�H��d�nViGR�m�h7�>��p��F�|��=\�R��םCfJZ�.�Wz-]�(	c����V�u1LY����m��D�mV�B���	�F��8���<����ɗ}���{'	�k�������b�ለb��+��p��y�A�/SpHP�)��xR��`�W܃ޭ5)�l��kv��Y�Z��m������vѡ3-	˷eƅ�ͽщ����$t�=;z��u;Y&�ѝ���=�AT9�q��V�k�i��oMX0˭�}��Sf�5b�c��f��֫��\����y���=pM���uz\�5�9Ԯ7���[�\�J[7p޸�D�)�fu�iCZ��Ù�ql4�<����a�.���ZƭL��F:��Ju%��`:���b��{x��9U�0	��4M��)7\Ov��S�V.�L93(���g^��6Y�V,uH�xs3q��tQ�ku�|p����_]��b�^jt%k�=�����t6�U
��a��5�)r���5����Og���Co�5z��w�X�"��,B�]��Y �0[�u˭�u��\uu
H���i_L�ݰ��	����y�óu��mX�n0ފ��@�`MTsGZ��Juwe�B�jt�WY�ub6�I]��|/gFجcj}�UI�]v���yo����o8;K�)umM���s_:���m
E�v�O5+&24v��l��S���վ.����7#p;}���:y��.�m����V��<޶z�լ|��������	���ܦT���-��y��\S皶��g#|{�.�Q8֓�F�ռ��7��;v�N@��3n���PJ�h�w�ZՎ�&�W6��c�lv�CV��܇J�(Xm�瀍�	���nؾֺ�\j�#q;�T��s�3�/C���K��(�4"����F����j9��CC��=����xڡP���u�*����ġ.3���Zsu�0� �1��ᛍ�G]��PRP�z��a�Y�"���ʃ�{�bķ�9Ju8�{'^*�@�S]oTۘY;.��8�|2�Y*�� �gq�
�1�(޽�";Q��.VC�� &䮋����M�W׌a�:'v{kXb�Z��s��I�f���pCiU�[���}	. ���}�X'ξ�(�Ce���O9�[��\1�j�c���K�w�@ެ��㻴�VD��X*m�]�G����V��d�w,��!�#�i]�3��I�}׭.�j��(��ɸz�Dh��\�3��>��Jplt�v>�UĻ�[$��W�Yx�L:ݹ���]3���S��6�4�2�\ŉV ���6E��-�Ş՘�"���3�e����h뻼��p�1�r�l��,+�ww�D��5�.��$բ���yq-�ۇә-������rU�V��ʍ[��bȥ����|�6�YN��{�����6��"�Hͦ����S��2ԩ���f��Bݽ�SF����y0�tN>+�P�{��ܥ��ӹ���"��Pͽ�Wn���'jMK�T�c�"���9m�	��>l��4:�B���|mc�V��3�H�wӻ���
�(�Kz�wͮ'-�p7�U�5v�S���2�<���u�i��L�Df�w�+_d�l��L�Ɔ:km�r�V���ı��e�I&Vt#I�f��YiVR�X���(,`c����}�(��ȶ�Y��Mb�|�>*���3r����MN��e�m!"C��{Ɣ!^�[:�(%��q/
��-IA�/�<�qZ�hr�0�޳3��G�,["f�����L/q�w���T��CO6���;�oz��;4��Q�h�0R�����l�[��$������3#�5tO.�.�&V.�n�H̸�G��$K��-k���f`����ؠf��;�s�@��a����ˡA�\�Bv����X��N]q
�;�4$�͕���G|rp�	�8-�(�����Gk��ʔ�u��QQ࿳G���]3]!r�CH]wa��l�ax�;�Bl�ܜ�gj��ڲi�i��q�P��I��/�4 �����v�"jJ���R r�M֪�!gqBErm�e����;�ي4ʦM���km'sw��凔����۲�qj�tT�>$-uIٰi�xe��#����Y-<<72���	�e�J�V��8.6:ݛ��yyMs��p&��4.�խ�e������;^�>](�,����_)��r����K\�X�=��q�3����ɂ�tj�E���2�ޭ�iN�z� ԃ�/M�9݆���e���m����n`��u��'l�W-��)�h�M-e쏏Ӏ}�����b�`�yL`��g�2��Y�i�a��&��4OK���V��{������+e�6�s�L����nwY���c8����>�h	V�u����o@��h��+VI}0c��'[�'#@a@W[�y��3����3%2�&Խ�Sw[�\�o����Ĥ�nVBd��Yc����ݘ5e�Ҳ�)�ekm�%�I�g�T�P�ﵞ�.�>݋G_4��������΁x��g���ui���܈�U����F��8VR&=S�Ox��e�i�م5��Ϯ&*�>��@:�̊�dt�,U
�t��Xqm�'P��Ԯk���x�����-�>;[��R�m�w.?C�)9�����"���@�IF�A-H��%*��Ǉ��9���f�.�p���u����e��#�9��N�0���.e��l����F�˸޲�*2AT�*ͻ�[� <uk1�k�j<T������y��z� k3�_-�a-�H
��"�+7v�[�j5�L�t���m�4Ž�HhR9�gUh���`�aK_�u}�f!��}�/$�������/e�`�XNG��=𽕝�E�V�,��X�� ֊/9���<W�)�C�\Y���הjɴVs:�.����L@%��*1�f_'�3 �ɀ:��5�>��+�4J��Ƕk�̬ �.�n�#�N� :���#����7wf���{�aSn��-��N)�3DX�g(�4(���A�ݙ��&��gr�)���P�?�u�ɷ��$��g�z�Ȅ{�%�Lgj�%����:�ٙ��p�#e%���i�����5>��՝�B��)h!&���i�.4�g#fw�-��6��k�9��e��+�p�Q�u���VX{4ٷ��RI��M�.�wtn�)����_.\&��p�Q�k+�������V�}jt!���c�^pQ퉡�(X�N�i�8�I�F����Y˩`�:���J����/!����r۩\�#\R���α;u��㾨8M�kK��2Z�Aj_Zt����rA �u�KB��r��������Awg.�M[2fsZp���Knu����j9��'�h�-Tk�L��[�`�a���&����i6��w_mڡ�3�g.̦{~EU�#Y²�r)�46��[��\v�d�;w�U����0Tp��e�n�U��{�~v\�PJ�t�g����������z��̧"�*Rɩ-��T��h��+K1W4w�VU�r=��^%h&��{�_k�Y�y���(����K�ZI1e�r�����%3�n��Ɇ��x��'��=�d��Orj8�1����kL�1�®ءD��lj��8s��ʼ	��/;p�+����;\(������zpt���q�e�ٮ`�����t��,T���j�[�����@�M�@�<�(�;��r
];t�냭�\vP�XH���g-�����aN�湏��A��9�}�xM Q��
Z�د,n�AK��g6�*���s­�)�p��Z0�����U}��  �$_�@�C	�IF�̐����Q�'��~:�j�9ֺE�|���l��w��_e��p��>�@��:�%xt���2��ێN�]%2E1b�kQzA�[��e�A2q�ul����/;�4�r�p,��pHY��j&C�w��/k�ol�Շ�?�:�;�e4�R���j�y3j��y|�Z���sQ�?w�Jk�V�\���Lp���-\ϵR��!��%0ieѮ�Yep��7gD�V]����� ��dע_)z2��Wz�ü��K�&�������v� G�nUĀ���0,	-A5W����*���#`N���fB/.���nX@8�I��k�K�Wr�T�5Ɛuq�侰g�	YP�ok^o4�*w�6�91����j��2J�m]�)�m`���z ��wu��l�kB��0�������"��1��C
�fe
|Z��kj$�"Y+`�|��:hiѓ���#����*}}��h���F�(B���/FEv�%���Q׎�g�m�������1����Yl�J �"��g��յ+YXe�+�EF*�YA�.:��*E�kE:E+-
QX�cb��#ݫ�-J�Q�	Z��dr�U����V��PК�d�D��F�XUH��;5a3MQ)S���5�P�U�m��k\ʦ0*(*��R��ZVDA�es)��+z֤3��Z�((��� ��PPX�U"%kY*
AB(�`T��)-��DTVPueW"�����������|�����6Q=���Уܻ��m�Z��ZNb�n(��Dz����阏�G�G��q�Xhlg�oma�T,�=��ZT
~�w#�-վdޚ��D�����w����vC�4�۴�q�J�IHa�j*�'�S��t��?J�<x�Z���s#:vMM�rCQ��1R�B�1s}�Vm�t�k��n^�7xbjM��D��:�t�KCZ�[.J�	�:���=�g;4K���7,X�m[h����(��"�/�u�Xx'�-NI��.�#�9ڸ�AZX�����\��s3�%��-�܍_�i���lՋ�Le�,�<�K:z��L������=S��ʹ�q��PGU!zivd3�=s���SڝX��Ҟz��:�S��_�|�]vձ-�6jȓF$��r5���Lu�������n�nhCJL.p�W����[#g��e3��rN�ط04zKi|4j@��3x碀��檯��-�N+�Tz4��Au�7kd*]Sw�i����~C¶i	ɱ�=Gx��qmQ�M��.�K���
.Ş�t�p�.���0	��{1fo?)��ѝ���%\����^�]�n��ڻ�n�B�����ų�5U����!US��ћ�R�;ɺ7�Z%�P�]#��֤���UG��p�#j2�]A5��gi6�6
��+�WN��x)@���Y�W��Τ�t��c�o�t+�V�`@�;^H$�nlӕ�R���)�C��3�J�|O�7���ړ,�α�\�'E樟�u���s���z(^G`����w�U��E���x��mv�f��6��|�"ѿ
��WM�j-��)�����n%F��x�jt\�13�Ij��q��!jOqWi��٢���:EPh�	nvsma���Ur�E��]5� |���. gS�<��64*��(����^ž�+�x;ڭ�ހ�(��hK��竺�M�x��Շ���7���Kn�d�l,��F�P:-���(7;����QYD��L��Tdo�uu�p�|���L�buJ�`޽B���X������tfbs��O&�tkU�>�k��Y�o��/PO���$/�ׂ~�3h�;}���"�W"~@���f�%�`����k0sJl�~O��\;���q]Lݖ=`�{ޙ]<:�3�����jsj9�Y#���Dא#��J�jp+Ǌ�����}|�'�u���i�#���)�f�e�a;�c�sZM�n� �Q>�S��*�ڥ(jxHO��`:,�/V��a-P`hy���V�kt/�V�޵{�ib]��Y�'�V���4�cZm,�C�f�Tݤ:m^�����'~����ed��T���q�wt�ܻYSd�M�o3�le
�ws�|ͭ9����2�����R4�eč�j	�p�x���W8R��M���y���	�X�������\а�l���y�˖z��x��\�)ZCs�����������Y(�<t3��'k�!�j;j'=����a�2���y�>�_Xjgo<[�Ho3�	�Ny\a���\��& ��у�t���S�3n#���xw�.R$��!�ѩs���яk�\�F
�!�	&cr4��H��Tq(�tV��u�3z�ӏ�>�Sq6�j����{Tд��K�w;& �1+-HRT؀Av"���P��
ݗԈ�����װPr��A��/fo<ʂqu�TG��li�O%�*�L����F�f���0�yU|� B���T�EA�=�6�Q����ȅ�w
!��y���;�jM`"�&���e��z���~�M��ן������M7��0��	��;V��Y�HPv�H@�9=f/kE���4��h�F���/U^URyh(n����!P�-��s5
���eN��g~��]ǔ<����Sic��w�� �V���v�]�[$ϝ�UQ���͍rvӻ�h�Û�6�z���]�&c�u[� 1\�W�Vm��������-c�kS(��.8BT�m��UŸ�a��sR�%顓'G��	�F*�<�:�k��X����ڑ佚OR�p�����N9J�Ҝ�[N�и�2���w���x�:�\�yC�j6=�B�����6����~|��ѝ�dK�Á�u�k��� �.�/��ۭ��zH��@�crmbE�ّrM��'h��_�f�[}���m�c"z
�ap�e�I�BYh7��͋�F�LK=Dl�f(A��Nk��<޾��p=g�}B�&OGv.�cx��^�QŇ�/Mۼ@{��۪-����l۴v���m��f�ݢ�;����t'�g���;�(ڕ��ދ���B�Ɔ���G����d�����{9gG����:H��H�m}�a.�·����y�����ƫdrG��a�>�:-GCq4/˪-�\a�1�������4P������)��E���/�z�Op2�x�:�0�Zx�dv��\2&d���󳣨�U.sBm�~�P��6@��q`�ō�m�`{��ot��jX�p�&����t���L�1���N�S�D�F>u��u��7�Ȇ�J�s�/j��F�Mt�L=K�c�����'jg*[ڌ�nS/^�!\���]�p"��9�i:d�P��ʧ2�\�l;"�Jx����x׫�)���m�ؓ�[��`i��^����s�ֹW.t�e��k�峩+��Ҩ�]as�iA��t�W}�B���T���3�hoW�*�5���]�;s	[2G�]:T$J	�8r)�oO]��>����>�9!f*�����:C��qa�Qه;i,X���������Jy�c���d���@C7�]=�U�-J�Oc��컞�[�&�bƻ����n-�����tvň���n��&�&���kxg���pz�`fD�w���]���@��]�+ѩ] �Q��ȦP�՗�+�uf��Z�h���M�`	���һ��U ��Z	�z�L��r�}�@xO��WWv���Zע�[��D0d��-�/^���� ��.e>OKp%��A'Eր�M���)p�)ʮ�*�F���wDQ����#��f���x���eAE�~�"q�{�|�qj~�th���ޮ�w]�m�8k�Su���C.yd��5�Z%���̃�1�-�*ӊp�5� ��k��62M��qi�f�F��`blK��Da�r�P}e&�����f��.3�B��͞��9U�W8��:b�v1w:��yc9�J�.d=wn��]u�:�i��:��C���n��ZKS'���8�ۉ���:���d!�{�����1S��;��l��%z�#���x
��r���غ�<�1�J�����ZV�u+�fuhyЭ�r�W��Tf�f=������wA3��W9�{�]HvD���f�m��yL��+9!sIG�c���$ُ(L�#z��̘b���.����i\f��_�fs[k���R������}��R���UԥorJ�� �[¯&e��f>r�љ�ȕ�^'�F`xw���=GrQl9Y�"b�ŝ;�Љ]_6ko�e]�Ҏ�b��!!rڕ���t.���<���̑�ط#v9Rʾ�F�k�t	�-��5+e�O���X���t���_;Ԝ+V���,ڸR��Z�Q�Ջ(bձW��u1�����Z��I`|�:�&)���B�$��=i�X�a)2�]qg!��YWQ4e<��u��;�Y���bzzˋ�5۝��"�g'λ)�n��k(d�G]4��c�Wݬ�͜��.�I�4�UՐ`�}[����؛P3,R'%8�'��`��gvo���	:��\qb�lRX�b}6�#Q(a�X�S�i(�m�s%]��G&I+)�^��f��D�bct4�xM1j��]c�R���n�,��7u�#��X��2ҿ�J��=ݿU�9���]Z'������Ҷ��oV3��[Z�"�ͧ�B��e"q�R�VX�L�0�p�*�^dB��,x*�Y�J��r��R[�q�W�0������wh�BR��+�g!��$l]qZ_��HZ�Gyq��]���n���%�^7.��� �:��n�i҃`X҃�S������6�Q2
�dt���������!��ɹ�L�l��hC$�Rjk'Nv�Y4��be����3m�6����[��M�I��w���<��(UX�;�������H����Rb��������vU�T+3���
}1
b��1UJ��������,��
-j�B��Db�2�A-�V��m�8+���cU��U33 鷬�
�j�T��-������n2�\b-��c2�������*]%�QQ+s&,QUEf�5�Q�)T\J(��Pz��E�
�RVm5s*�nf"tب�5mJ ��G]a��HT��WF"$J$X[V����P�V*�"5+U��E"(�M,F(��Q���D��GG�Ͼ�n��puJ؆J����X��k)��]�4���Y�9�ӳ8u�R[��p^�}h�r�
}���Y����+xJ�SgS��$�&?_i�\5s�$���$��֞�R��Fh��y�%p�	���nݞ� �uY��+��]
��t��P��_j�@c�w ٭X�%q$�e��ӗ+	����}#c�(�ӌ*�p��l�b�n(�$�f�KBQO��y�}�-m3*�(�/̻5���)ו߫��B��} rڬ���Zl)�K�Ґ��r�BWvS�O�K�Tu�E��`��3���o�*��&��!S�����f,\�\���͢!lt��3�J|9U�l��E<|Κ��+�X��4�FL{��[�u�-5�*�9ݝ�����V��z.�g��L<�j��8Sj��\���y�=���_B^��=I\5��D��9
�fR�25��͕��u^��f�
�-M���u�{
5�A�r,
�����j���҅yc1���`S���9��y����x���}G���gK�Pĵ��ξ�*Q���!��]����$�R��¢�,�7�:R����� �:�.u�+��Gl��u���y�W�f-�A�MY�͒DOlW���E�3*��+%�	,:u�!���j��?��N��R�lx�b��}�CGL�
�M��w:�&&���O���9��A����τ����2J���pl�h��`Y�F�:z�®�j[��뒛��IL�"e^�+���e�������`��G�2�yU&.��h��9qBE����/%�6�	TU�`G7�7x96�i�Td`��W�C�j3Q�DWo^� 7���C��&�R�r#h�XW�6�0r%y��"� ��3Q`��uyq
i�A����~xyr���Xs�$O2�A[Yp� ��햑��~X,PGN:��sX���wf0����Gs�w+��E��
���ح���ֽgVEUx��Cb9YҶhݼ{8������`|��]�O,n�ogs�"���:���[�n8�:���%-epʔŇ�Y�Նج��+T%7���`y��w��T��e(�Zmn���9:�s�Mᣤ�/-��e���cGIH�2���0H;�b1q�qu���{���/�K�y`U��z3ddvO®�ؿ�;{$�bX���,&]-^���<��֌�vNŭ�@�#gm��e�ŤJ��oNz]ܓx�n�7Ŋ:�D��g�W���>�X�k*��Q��Lm-��qe��G��-T\��3��QI�I��<I_�5�H\�m���,� �v�}|���~��
������XCi��̇��8ȡ�!�N0��!�,Xbv�o�0�L<��$�μ����p��ߟs��ć�fI�Cĝ04�$<I��i=`}C�@�4��NZ��q�i';7`x�u��ٝ��^o����y�'n��Xz�5�!�'~��@:I>@���$Rz�!�0�"�w�2m0�>�{�_��M�����!2ʶ:��Աl��h���A-Iˆ�m�XyX]�&��ٲ��s�{�t��	;��z:Pk��Mo�gt{Rk����ks�׼G}u���{��}�O��'�S(�3�@�5��	��2d��xi>`t!&�VIY���O�\�o��Y���}��7���Ĝ{d'���yI�8�jН��&�(q�3Y�C>�	���Л`)��L��ӯso�7�{�|�a���Ӵ�5�'L��K;B`t��d:CL�/� �'I=I���׊�\�;�^g7�7��'1��O������;}I;C^П2d�����:d�0��֬:CI"�m'l�������O���7���!��OR,$�d�>9d<`m�go��L��� ������X����������>�!�x�����E�v��OP��?'̐�[��	�N�8ϙRN������u�����ϳ�>���s��BnΒm����xɓY�O.� �P�I��8�|�$8�sw���!�Co�s�����7����4��i�:C���!���$���<d���D��0�}I8���|��gi�Cl'��~{�t�n������~� kvO�!��M!�I�:7Em6��"��@8ɇ��N05טN����gl�����Ǯ��u�<�ϼ�V�|�{�CiP:Ր������C�Hu��RJwv��O:�d��:z�d��l�{��^�b���~�.h���X/nM�>�9��z9�Q?�|ʡ�_��!J���r!y�/�K�ĩ]�v,x��'�+��:�ww˞o��7�<߽��I�}d>g��T>d=I<���8��3�odY&�tn�'i"��O�w��^g�{ם{�����Ϥ���'l��,�tuBm��_�'hVVڰ�������!�!Y̡�ָ����|�n}ξ�>���� �L��\�|�q�ԇt�P�>�����	�$��z�)�
.�ί~��p��:OXO�3�)4��h-��:d���$���$=I�	Xݒ)=M�d�����9�\�߻����m�d>���0���|��Ї�X�6��	���Hu}�Bhݓ����c�}�S�秬Mo�|��G�&.|T����x��!���CG��m	�=gL'v�|ɇvq�t���I��=�޳[��^��y�}�d8��	�>�� z�,7�@�$���� �RC��	��i2�:C3��q�7|���I練�@5�'�6�ShC����a��I���l��l&$C�����<�˝��~�~�0�!�>���O'�5�$<�ɶE��:�v��M��ClS9C�ԁ�!����N3�;ﾯ�y����}�����C��	�����$��F���,�$�VO�6��t��OS���Й�!8�>�ǻ��}���w�t�έ��C#O�5ǝ�ͱrl���U��,�K�w�s۴���s_�}��]�G6	�:K��d'28�N�M��SC���U�YC�~�=t7Nǳ��莙�!����,<d�����vm'hIXOX�̒x���<�=��'O���8�|��s3�{}=��x�!=I�hOR:�x��q$:g��2ٴ�$�-�|Ԑ��<a6�=�v{�o���{�u�T0>>���k�C�'I��'�8���ԁ�0��'�(C�L�'e�x�ĝk;��t}�u��o��$��>�DǈC	��q�zϓ�Hy�N��:
�|��d�r�QdXK�}|���μ�~}��8��&�>2�q��W̄���Փ�O��ݐ�<`k(C���'�P�@�,8��'Z���̉Ń]��A���DA���+�������F��@3[�C7AzI6����'�>�O��d��=@�!����>��^����w���'i!�P�)�!�,����3 v��d֨Ae3�	�CG�OP�>B|��
o~�Ns�z��~����$���m g�C�E��>@��m$�&�I��'v�:d�{�m�V|�����0��}��ϟ<�w�$�����4$� ����f�,�d�}H��m��&��8��Ht��HY�zŮ���ߞ�瞐�	�i@>��O�=g��������C\������hC<��:Bq<�����ftyݧy%���SY��λ|1�o�Ű#�kTt#ב�F�n���g�+uc�ki�E4�Վgu��f:T�wZ7>ź���d�s\�~�ތ��w����}��P�t���Z$� m��P:I��HO7a�!�M��<`m'Ow�$:{�<�9�:��}���;Bql��[!��5ݛd5�i';�� t�m�M�XM q;Cē�!�M>��> �ҥ[f�|X��>����d��S��Bjô;d6β�c&r�v�&��I=�'bN�z��m�=cy�=cA�����L�xO�M{�f#�}'�'��B�6ä1$R$�'��!�^�!㮬�dݰ=���>�N��=��}��LI�I�l�m v��t�m� x��x�;J��@��RI�Mud� ;z�w��5׾u�~}�]�"�>>�z��[��t���7N��i<d8��ߙ	�!Г�@Y����G��ќc��w_��=�>��d�@���I�w���?0<B3ά��'�@��hz�q��@ċ��z!LD����J�7�o.���6}d'���"�@��M�d�z�!����w�I��z�=g��o	��d�B{�~|���o^k:�O����i���*��b�_����u3���K�V��O���(vd����K����/ہC+u:s=["����{r�?>��k�#R^7:}T���ξ2Ú:\���oo'I�q}�8㏿S�̱d*�P��y��\�'��DG��w6�?�g�s��h���ly ^t}�h���)�a���(�1P��5��,�I22��D��Zi*R���M�#��Ĝ�z�(��ntu�)W�8��j��'��S�Fh�յ}B�1\2&c�oT�M��Ej�]\ހ�;��U���u��h�#vb���r�C"�=V�^���[diV�.7���eC��DZ�����$��H�k4��-�8�bж�<��F���'70 �Id�̀EƇ�\�p��qN�dڍ�cnm>GJ��(V�Q��|�&졝Bנ�w���$#v(M���k
�� �o;5ӭ;�����n��**r8�(Ό��'2�#�MZ4�U�JY������#����M�~DΌ�[u��S��/G.��@��]����ޫ�hKU�Hj��l�C���J��^��S������ўt����N����`�<Hi¾9������@��zuf���8���@��U
��^�9/j"�
��Ml��AdT�yܒK�(���D��U��oM�ZO1Xw�s¶�%�Tv�bj�[PD$64���$��-��l@��jۼ�f�_pX���X�,�5-���PY�����LN�Tܜ�s�:��:^]^��'#Z�P�'�]�$;�5�5t`�;"7q��n�2.&ٹ�`lU��3�CP�=��xd�.�꽙�`r'�iewQL����\����"#�B��o�O]Ҿ���ʩ�[ʹ��^���c�[9m-�PN��B�p�<&�T��m��" ���v�2�d�2�+ts��k�iYc�f�F��ɝ0�ݫ�-��w��
�.č�0�h����8{��1EW	�ÝfWf�����b
�t:��g=��F�
���0-�<W=����K(�|��9�5��V��J�%�F�ĊТ�X��ɍj}[Z�S`�f*��`��k��"�#��C��_*��%..u7i:Â�����2:@�eͬ�ԩ�o����u��u��4P��];bT���ob��f;e���ۮK9�n:ڊ>Y��9�T;Q��:�\�7��r����s��4�+���3�=�>4Q�j�A�-��R)0B�f�V���k2�3B�3K�q�WF�0jZj��Zyo%H�]���;�H��N�D�� S���8hں�#�0T)E�?v��2�!�;#,�7V`���D���X��jP����Z����th�iE��Y(�`��e�
�A?d�t��͛ ���6Ń�VQ��m��eJlH'��3Dͨ��5�6��4&'fR7k �,�+2U�.���8��3 ��f��E6�H��n���ӑ�l6`J��
� ����;�i��1Զ�e,�͗zł�?>w�����bbP�KF��v���Y������[���Yisٺ�1٩�'��U�̩�e��rt��)�p�l�_	�� 	�k�]�!i�V�b�F
�;jP�1�u_�{����ň�����UFEFڊ��l*�b(�DPQH��*j�[b-iR�Eb�e��Э�+
���,TX��UUU�����E�\���#��*0`���h���dX ��رQ���%Vұf�$b��Q��	b�KJ�DT*EFښ�U�TX�1��YU�jk(����H��G-���r���[UQTX���DH,Q?>��С��u�'-�?��/����B���P�c�]�Bj��UGz��B�j��'��G����_���;凔���wb:���낼�����t��M�Ӽ ���z<�2�!$�3���\ոM�UT@}x�F^ȅ�j��4rz���v�1�6&���CuZ�1=�c9�=l�%JV�Kq֍j/��M��,&��q�Q�l���V휏�lK\M�c��D9]}�t�=�p�O�F�\8]Zڔ}�yok�y졣$�vWL��j9�7R���w�����#S�v�7�^�D���\���.^���'*X�fS�O��!O��ޔG�86�q�"N�q{�`�.��yء��o2�(�?v�%��^髃9���iK������%�#�!K�g�6��'^.FLN��<�t�2EIu�E��着����u��ߖ%����Jv��I��^����af��"z��@�P6"�34M��&ӥ:�G^)nkF��G�"jWkM[i\��2��FJ�D�5R�F�IV�w�˭#-��b�;u"�`�I:�2�ck��������X��*����f"�Fz�����c5�`U���/v��N��g«���5k��zlxj�ϤJ=��V��GMo��=�&q�䌭����1���M�b������@_�_��hW����U�fv�Z�x����^�r`C��s3�]ϭ`���� �M�Y߳xH��]�sH_P.� uFmU�(X*�TL�(��%��G���k�{o�!L,���ǝպn
!����k(���s��Qn��z�tE b\74&/�߹f)���	r�q���]�|sjv�M[;��Ũ�w��`��:G^˨���Z�5Eւ `6MӡJ�R0о���,�T���=c�#��]�mƈ'P1d���/6bw7(1�������"D!*�Ͳ���U�<jxL=�G�{H+�-��*}�Z�Ԥk�`8̨>,,�~�vڙ�|Ï��[c;�/:]�V��cP[�:�8�]S�t5=)�G�+�3畐�#���Q��(�2�7V�n�zjyX�����QƑ�����x���e��As�e�j3Vls�3�ZCI�r�#�$f�Y����z!��٘t3���\��7��.��r�^YS�G^��g�ƭ��݁�H���|qn��;(g3����M�5ֶ�P~�n���Y�=i����V�!�q䉇#���֒��o��������=��`I�ފ�����{DO9᢫�m�w=(8��1|�V�X�%��ך��โIAջ�}'��-
G��3�/��wy�h�����bҺ����k�#��ʶG3У��\Zw�Q����H?�z�~��/?4��=�Rgku���_��[�]�vC�0�7֡&���X5k��Fa}z �Hk1VH�˾�����F�=QT�7L�2.&�.�уe�����9�[ɩ���ȧB+A�r��u5/Q\��Z凊Y%��9κ/b���V�m�臓��2�D��} [�c�tU�t�I�&1��ۣ[bB������qld�AmˋG��!�zY���jU.��7Q�G)ޓ��m���ܚ���o���c��R��Vi 5W�(���׏g�g�WR�'udB��4�;��t*Ī��b�i��{��h�)�e,�ѣ"(�P�뉚�E��D=�-�~�罐��=�З��éiCEӚ���D��B����)�k��v����\���B�f�o{���<9�2yT{��O*.w�`);�n+ʝ�ԩ��ש'r���#�=�{��00����x���Hvf,���V[�3c@�W8s�8�g��h�;]4���g�k!�'�G���g)��<���ܓq�ipf[S�ǻZr�E�t�,Pۆ��:,�{��c��^&��rl�tv�s�fr/�%������T�;�8�*���N�6"�|�����ʞ�%���uOg�Zd���f°n�5��:�8מ]�c��VTkX��ky���9\+�{�xyBÓ�JY۽�9=z��;#���ӕL�:;*���:�k��^�yt9��}�'C��P�7~��2n����(D��ǆ��+���V�.��*1'S3�Z������5[��+ObP�f�R̖��h�������W��!͍{.H������F�F�S�'��]{Vfs��%-��қ��7��'x?6�U�@<姇A7�ܶ�v�U�fs/��}���Ǽ��#w�-����nL�r�|!y~�뵐��Ee�-O���ӽ���oaf��n�|&h���sd"�T�&l�x�n�0����%!!�������(3�a������r��P�2/�����u�X	�9��	�
��V�W!�+�o�g�*�ʱ)@m�b���=��wo-�ʻ�t^�:�Bg�6�I����Gv`�ڸb(��1�:��}�*}�]޸�|�&++>w: �S�rṠϹY�)b<�(|]�ɘ�#���ovNVy/������2��F��jR��(�O\��-W�8&C��9�ϻ�k)�7p:�5v������'P�WH@�@EZ~p�gf�J��1"�C/xFFVsM��u/��eb!mξ;tTv�s��A��EC�|*��U�w�x.+/qu=�����RzćذC
���Q�fj4;��VYd�s�{�wh��B�p�V�����X�0������T����҆0�s+.��"4,�13xĈ��S�N�,4
�$n�?67k`��S��l]ɶC睽�s"%�ML�I"';JQ�rOQ��9�"a5Eos���W�k4�Y�]EL���{����1�=?}�YdAla:#�FI��b�s�hn�l��"x��\�I�O��vi��s�{%��7�*�`w���>�b������LFE��o��׶�a��[jZɸ�1��ґ��v]���ՑJ�D�l�N5!�w@|���Y�E9���w��}.o/E[T�jgWZ�p�*c�X�V���pL�]rШT�Fʳ�Q!�n�"ݝ�/D+�����������3f:��I/K'oշ��}�"��x�(��H������gA���=ǹ�3.%����N�����:*t�>����p��#p{χ�n��od�s��5�1��]�S���r<8�4otB^�Y؏ޏ{�苼z�o.�̨��ʪ�:�Љ�܂5�Q���@iD�q�A�hLЕ��A��\
�z_��[(���]��F��p��P�Z��r�Z��է,��Fw��2������>=]�C��������8��Uu�6�E�dE*}�ռy[Y�)�M��ـ� H7-��@I�F������o��*丣�-!�6j�]
�6-�
F짺�˥APn虛�Ν��qY�T5���Z[��n6���a�ɸ�n_F?~��寲~B/~�j�}�Ê��?�S�|���~�[�]ʹ3��KorW!�$�E�[&�̥�5v�O��%#}�]L��xXCX��R��1�>�7�	���&���|�9��x�3W��`������:7vw�`���V�)�-[�����k�׫�{W�z�4��Vku�8��l%����t^>}��P�H��}հ�%j0��ෞh��A't8�Z��Լ�k�!K|�M��]��q`�xh��V�y�M`�d~S��I~�c�9W�ˡp��{��O�R�ES3����\J������y�v�[]�j�o��v�@��|.�v�Bo퇶��Xn���ϗ)�mI�4u�÷u�
�|�ŋ��G@G@�ue�۝SM4]nM�G��m��� ]:g�/g,����,o:4��mY�t��|X��u�N˦�ش��є��
T��u�F��e7�-e�2�O�kܺ��v����Tn^�˧ޣv��>tº4đ��۵M���ml���GYqI��_�F�`	�����ֆ�m��n��pU��e�����%�H�������R6��KI2m�[Ę�&"iX�Y)�x�������̰*n��Ee\��2�fJ\�s^�b�5-�p�/�VAh�LR��-e*��H̊˗Y}�V����%9C  ��L�wN�����˳Ou�������ͪz��VVA���i�Z��*����u�B����P�y�`��v�on{J@¨A�n$$N�yBS� B6l�Rb��9�L�ϯpn[�+105�/�2Ɵh�|oy�2��[+�W*�)v�K�\�ed�9Eb�b�FR�c�
���=bf"bg�2�*QW�PQ�J��ΨUE�.9�b�c�DR1��f�D���X��V"8�Ab�kA ��*��Z1���(����UQ�E2ʍ��&4�,UT1�Z��Db��(�AAdX��H����#F
��+	EDZ� �AEQTP���c"�@PQ�E��`�AE2�`*�(��PPY��H�QR�*���"ȱE�UB��y��]����g�oa��˩[������=�	��Q�}Et![�H���q�����{�f���V��ȅQ��p��&��E��7�����[Z�����E!~w�g���4d�;v
h9y��4�5����i�����M`��mA<��gk؎x�YٰQ���]NCh��d��7H��;vf�FUT=��}Lt51�KC$L7��[%i2*�.��t\�(':�=Qֹ>�ޜ�y��v���@X��m�T���8X���g0B�4�v�X�n�6:����R�q�Q�C��J�g̪8�&��:"{�-]�Ϻy��EpG���-]�/��sw��TBlO�@��H�u��L����dJ�cv�L�ծ�0:���$[W83Kv�p����.���>��Z��(Vо��5���#h�iv�i�+3n��9z(�5�0�g���{Շ^1/m�2�hX�O��993*����f�nJ/ o�eP���I��A�r_�7�7"�k��q=��<8�J͘��c���R"�X�Y��1���j�;�W�-v�8�2�����f�D'�H䥽'e�)��6ǟ��.�U�i{����K�evH1Hw.Ғq��"S7:�vh�յ�nMa���<	�LT
���8vƪ���]�q%�;<x'� �f$�� ,[�{x��k@�a�)V��i�׼w�%t�t����F���ؕt#���O�������������l�Zunb�VH¾�G�����7}�w��\b��Q��ޗ�rn�w M�pNߺ��7B7���{q=� �J�p���3p�
��<�4��t�i�E�\>���nȡ���l[�
�I��o�D�֪4���t��G�a��}۲5  {q�%g���;�]��F�Ȥ��v��G��d�I����{D��$���:-� ���O�jT"%�n�H��97VX�8�,�?{������އh]�9�������¹ �"���Fż�ۣzk��<��yv��5�1b�B��R�K(n��5�VR΅�ۗ��&����]��y�X�7������􉈱��V\���TS���2�]�P�\�ޏDF;\�co��~�`A��v��[�Ѳ�Kf��ӊ${a�U�hR�Ҭ�Ю�4p��(�E���@�3�����
�N�}O�v�	�C;T�nȌ�p�T+^���)����c^|�����|�f<�ѣY:9���^d��Ժ��rVtP����+$,0�Q�}\ͅ���ѣ(��s)�ƈ\QI{�M�%���Fdv�܁-u�+�Om	���fv��CIrt���K*�>ب��7�V�(�u��2����t�
�y��v['S��p����0j�S����qw�7`�2ĵ�����$����nos^>�����y��÷�e�B�!>��Ǭt`�=����y�ﾋ�iP�N�&�ƪ0���]19ky' 8UU��_W��5��wc�\`vu����]LsV�%Jv ��Sa����/��ί.>~�[�mq��-�(�Kh����Ĕ��6��AҌ!�]j�{�,��@���Y床�0Н��]GE��D�f�/Ҩk.2���
�Y�)li:.��E�.Ti�t�ŉ���b�ds&a��84;Kyڸ3{�"���{��>�8�>�!��:��6Јq�V֧����7�˜t����mͭ�7mR�N�I��/p��ʑ�,�FY�t=*�ҧR�B�x�ʹ����͗��e_2W9;9�bܛ#h����]yùS�L�6��F�.oiªh��=���)>m��[�5�>�4t��:,��n�����5:]y�a�}֋��0�iN>�nUK.�
�����zV�%��LX��D����!��l��P��W��0zTu~�dX�N����`D��9n
4�Wݯ��'e�$*��V����EO��{��+~یVw�]�t�R���{�e��G�5:h��,�sU�>��MH{�)׹�Bζj�ҹ�7Օ�:��E�/�q�m���tMߙ��n]�#T��+3�P�&L��Ier(:�;�9m��6��E�n(�c�wK��@�2ru������U_|f��צ���GѺcP2���T���U���N�Kp�Wesf���}�{��LL�|�p=���ݦ)Z��7�[��W�@�W��K��6utc�*\�0v���g�p��.���d�/7|UרRf����~5p�a�yX̻R\��R�m��s5&\H�.ct^O�D�sK1V ,Or��(���t�;�
�ęm[��BL�����7r|*���O��.{5"�k�/3p�LYc!���V�>5��NL X��FC��m߻o��`�]�>ゔ��R���:���K�%��+�4��>�"�뺺�}�ų���'��G����^�<
]XhK�t��hV�w�3�jv���]n{��nu�=����K9LַN�^Km\�Wh���ԩl�I[ք�����Hl�d�g2����W�1q}Q񊙮W��J��O��I*zvUQ��W1z��b��-�	E�L\��p5죂�'NS�J���\>p����̈́�b	��#�=*\����W���ڭ�g�e*�R�q�:��g^l@���E���*�:�?���YMA3s�bk�o��`����>p�����j��4�4d�@`c�V`�xo���)���a�����:���ȥFz&٥X�	�y'�%�#S1ӚoC�WY�ܫU��L��֟O N(NN��Q��X�>��gE��|�b���b]��V"�����Ȅ�,?�Z~*G�|�`�z�x@�tW{��f�|8"s']	O��}n�l��Zn��3S�Fa*�F@�v57'��QM�.���QU�\vS��W�2��6�q{L��yZ�d�&U�ap8#J}�b��t؟7����0���`��#��p�EV���i��DG�m�e�D�j��Q�ߋEo���ʼ0X"��pCVX]���Ǟ[]u��U9r�u���i���^��g'Q�c�\����M)[����0�u
a��I��4����<):����!�����o�S���Yx�!9�3�..lӘ�U,"�^Z�t���r����ug��c]ȥӽ�9�ֈ������*M�q���D�r�Ky��>4b�yO4��WHj~u��1��4�*��a>�\=%p{�Z;-��n���էq3|�K��!ѡRŠ����s<�}W�|�Q�[���)�U� `tO,oKO�󻹂'�&�0|��e	2x�AW=��}�Ց��޷P] ����
�n�U�+F5F_)��IH<�n��WK��2�г$��G��}:�e]����F�����f���9ܩUmi��z"#1k���}�5ۙu°&xU�4�IQ��R.��m�eC��m����f��/�W.h�U��#��U�P�����5P�&[�2�/ܠ�w��gE;60�>�[�1�5g<R��Ɋ�*�1�.&��g\9�g���K�*�Ur�	��gohթqT�NB7��dm�5���&���\E�Q.�o;�|8�\!8��;6N�p*z�~������W�3:v�Q�>�=z������8%���g�^U�������3{9�U;\)��ᮭRQV���T��2���j~=1�^I�����z�C�r�u\���I�1�"��HYPquk$��C�d��s�
���Y�^Ī#�]yp�~Ѵ ��T��;�׎��Au��n2O�G4�q}���=S58*
m�:�lv�#��\�YR]Z���]s0d�B����Z�{�^��e���2�,<�DM]a�3%�d̴�i�1�%�G'Q�}�t�p��[��'���%��Δe&���Z��g(�X�\i�{�F7�| λ�љ�H�p���yI�e�o>2�S��!B����`�1��Ô�%�n�޶ؤaw�h�,8]n�[���7�xm���}or��U����u3����/�	�a@�9��Vvҫ�g	`SP�a���!�e-��Vlrl�rQ[�#!���tgs9֩I+V����h^�wQ���(X�])��̧�Ti�G^\kUɇWlǺ�Z6��ҕ����ua�/6��ԫe%��e��7g�t�p'x���\k���iK���cf�ι�X�<h�X�̠5�|��En4R}a]&U����--�N!�a����e^��`��f�2���E�[��1�#ʋ��h��st�0�$]�����mVE��\c���9�Zy�b'	&)r�#���;B���@�m4&Vc���HQ9&*�{��.|T�sg+W^ի��Քl��l���V]��)71_KmN��8Эe���"'r	f]�b[�(jNO"N��� ޘ��W]�r�	�K���8�W+X��LF�����{�h���r�+8ŀl��7^i�Q�,��� �ȭ�[Op�t����̞yڻ�����`�$�\oC�5m�|)vjU1�M�wl�����*�a9Ȋ\��Δ�	N��3�}M+y�p.�����FjЙ1�n�k4F�����u�H���ѩݩc�!�"��z�ّɛ�,�7,8m��`�5v��*��T�C��ǹJҌ�-���P:��z�o�fp�!bdPU�A[b��b�!�"���E,PQ|IX"�E�,TE��UH�AI,�H�D:����QUY�
�E`�hEX�"#X#"ň�����EQ�YS"
�E��j�q
�E����UEAB+*��Z��J"����duj
(E1R6�-l*�"��IXdFL��1"��aRV%��p`�!UJ��XZ�
���������{�k�g@��&�z�X1�+!���H=]y,uJ��Ů��}�U5�;�������e[� 닂����FU92�T���]Φ
�Z�223<j`e+��a�Ux��=w���ʅi�����8�ջ&n��ؗ�]R��EY�J��ʊ�ۤ�Ё��������V�i�s�z��2�b��T\���2�#����5{��2]L���i�jX*᱙Ip�H��ey!Q'��.�_�oXˮ`X��^�:��*�ָK><�k���r*�D��D=ர
ʚj^h�\(��wO����g�ᐋ}weeq�RP0��|txx1`=������o�n�9Fz�[���)�٪#ȶi�`n,ƱV�wgG��V�@�n�R�#�YN���4T�(��w��f�-@`~��>��*w��,���y�>`����@�9�!��:�]����a�˱t�Ґ�"P˚�{���w�6f�8����6YV)e��=�HڋK���zs�v,���DG��s�׌(̽���>�+����U��3\ �i�}��U^���|0���ֺ�:��b�S���w\���Ӂ|L�q�3�������U�����+2�V��jx�u,V3,:;0����0�퉜���mLuҞƈ���G�τ�P�c�@��5���9X��������3M`�"�fD�X�p@5vf�Lpr�����F��UO5*
dx��s���$�@����^:9�N���[�g�F��Q���^ּ��آ8}\kQ�ƞQ�<~uZphyMXtK��^�X!E�L6���>2��}_��wB���d�s��A���c\�U�>U��Ѡ���_j¨��=W�7�N+��z.0����'�F��Y�̬�����$�.ݑ�e
v�OBEm�Y�����Im�6�24�G�2*=�uJ@��������{���ZXB�(��y@�U�׆���΁������qd�;!�D��-M��mT)j��xT��	2���ᙯ�ngt������V�1�A��z"|0U�g=�f1�^�y���X�"I��7]f����)�-٨���`���;�L^E���LVg���vf�"_R�*�ty��c�;��D|4��`��+��ܷ�$4kQw�|�4�VA�q��gW�Nu@Ԩ
���!���������5�/j���|����
崫��j���B��h��[jϬ��x�)��_i(�[�F�\T��r�5�6�&�J�c)���S�<�b�X�P�i#&Ό���*$U�U�"�z�3�&)���s$�{�[�qL��X�t�e[�+��}��ԉ�b�{3�Cz�:�NV���\ήsGY��R�;s���s����n����?*���-��8��^��u]_��Z��f�ΒE!���Q��<'�ѝw�穪C�V�P�+�T��t<�Gh�)�ҥBczm��2���*��x���Z)׎Э����;��X���OV���t�8Y?xhy��#�;/�UQ�4���w�5
^+
�r�U�������0EA���ϸ�d&uZ���W���&���5�T���~9Wʡ��k�0xW���<��Y��^�d*�ur���g_H��ݾ����B��0���wT)CVt�NI�a_��`���pl�_����R%����̀m׳�*�\/�E�B;������=��Uy�&��`�I`�����}��	��z����2�ȝ{��6��p���\:ԍ���t�N;���9V����W���S���%�[jg}�խԷ�+曲�P涓]7�f-���c��_nv��p�pVY�?�h�iו��J�������O�$]��)�/��������P�ύAD:���b��!�at�z�'�7*\s�C`�VS�8���.-2�ӡBݴɝi�ί]�vj|���}��g�m�����4D����C���Ǐ��κ�o�T��PR�]ep�w�2��^���{% e����'G�`��C��І���V��~��(��V�0�T�P�W�|��v�P�	�A�������X��q�R�pU�\vet�� p{�,/ ��d �*��R�:�e��o�"����ҭ�������b��w^����t>��$U��:ȴA����ިDyr�=�J޳A���E��Y�#XU���n����l{�B�[�+r��v��7ss�h�&.�w�P0���+ɭ���M�_���Jl����Z5�^:�C�k+���V�+���]�s4��{��(T�V*,��(a��R�'e	���y˫�k��mP�&��³O����j
@�٠0n��t i���z�l��{<*�4`�51�9��K&��~��W�o��4{ܴA+ưX�|xp��k�E��C�&���q��ȷ}�c-,�\���iz��u�%�y�=�k:7���������̩0��b�y.�h�6hec�2�@���w����&��D�Efc����N�ؓ>,Sq�2]�'�M�a��Y������`'W���k�Yꊝ�/�3uɆ��ʹ�u�j`p5�F
�6���R���Y�CF�u�y�(2koW�<m����ͬ��S�U\�Y^���p@u]΂녜[�Rin�oW1�M+����7'$m��\��/^_p������_����cAV�|8`�<xs\�?��j����hrE������V���%i�#D�+��f]{ Г8#/��/�CM�D���OΔ�`�+V�f��t�W���tc�@`"���Y2޹}����N$���������h��[�od��.{{�`�}��F��!^�\&��{JI�6�%�GzB�쐒⛴6���������p���h�Xu���A�'�ȶ�Y2��L��ciN�����z"(/�
���B=��}��������{����l*�\:j�GC
��cK�-\�{��1\=��WF�<br:����c<�M�}Y���͂�����M*P�lK���ˁ7D�ۮ�熱Bj�{Μ�Ctz�rVZ�mBpd|�]Mgd�/��lv�z���/ņ׆t���33���՝��M��j]��ш�z���4�O4,7�us�&���=bM+��_Q�Ͻ�{��o:1�+��Ty@�Ma�X6Q�|��IBg"H�W�)L�xQ�58jQp'�g(Z�iH�{1�Q�7Z��Qm	[%����5H*��KuR� Q����
�x�=�w;ٹ� �����^� "���(SCL�r�#G���^��ʺg���M���m�ͯ'Q�5�I�R���$��n�YC؋A��}�@W~�s`�_��սy*aC�4�Hŧ9��  #�	A�C��?*\׆٢4M��8�-�-���0���ғ&}���I���3�CF`ёm+��T���T�k~���<@�\��p�]y�����Ӷ�F��uOK����NT&��/jaz"�ZB�f#D��^�3oվ�Z�Z����h]���Ab͊F�E.�ͅu��Ӈz
�{��y��~�}%��-��T\��]�c��u!�.����1�]R�pD��h�����_h�T&>��U*g��o����+8T�V|�y����G����s��Gܪ�+F��S�a������Ux%�����{`U�Us2eH��/���&k:���	 ������j����P�b�K
�t������CԽ�I�ޝ.����~�H&#�f��+ w��ǋ��t�q �B�J\��W�b��x�c�E��5]L� �OK���^g��*�O��'ba�Ѫ-��5<8�'��^o�篻�G;�e���p�C}�K�tO�����.�q����z�Ѵ �����Q�d�:�N'�x���@�����$a��ׇ�*���4�I4��80<j�ʃ���zn�"�Tfr4����u �[ϣYw��o �g�Mк�)�kt�j$�2Q���ӓPl��N�!�-��h��l]��g��_Ua�/?��'C��m�
�Z���h���פ*����&B*�Ma�}r�$��������*�랡��,��ʅym)Q������-�eFLt�2�:�f���>�@���Y��O�~��3M��Դ@�AY��Vr��-O�}+@%�,�p�2U������.��A�ځ�w�$LV�D7RxEl�*�Owo)�~�
�V��� �}��e�O*5\*K�g;�gam7f�p�ZiÌԡH[4	ذM5�V� v��D��o���+�L�pV��PV����dN]Y�ʂG'{�L�V��S��X��U�>��XρsUh������x�Y+��X�0�Z���p�L_�
\���U
c}�ӌ��v��́]o楓k��^�!��R���#�-���V4]_c&�찤�pV^o5�aGj�ᠺ�~o:r����' %X�V ��3+쫫�m7����MWy�e�bݤ���R���N.j�̕v��Fs��r�_U˃�����ו�jue����:����s#.
�`fu,}�<�n"֡�Y�ZP�ܫ��	��3�����w3�(솆��sgI��}�c���3zvcn�z��a�Sl��G;,̤++9��é��I4��$��	RBN�6Y��O2�=]��>[�6#�*Ȯ���&��;Dx�?��nK|�tpo��T��@��LQ+�mT�@�)�P���`-���,u��.XL��0^}���L`��`dg+��)����s:,ޖ1V�~��.����&��vMĥ\���2��!v子$�ې�Ϩ����g-(��pnBY��䓷Q.A+�xΣ�D����v�A����}���eQ�%��me�4Q�m��Q�Q�,�sk;����N�Ѹv��8��hv�J�h�1�GR����[�PWk�s�R�׌UŃ)�����a��V����X�QlKZu�/��5L�qoVĹ��w�2l��n�f��k��!J�iJ�*��F�;��Y������8�2Nz�u��k���}#�y|)��/R�h}�qw�s�y�t/7h;��u���f��\WX9��o6S���>���bu:4������>��;�J���Z��J�+�k� m�e=W�T�PYV�)>t5���뮢�sa�r;{�x>�7�:E�u�.̵-J�Ӕ�OV�������)Rb]�L(	��X���kh�r�vko+w���X��2��<���L��fwAH���P�Ě�L5��B╥�$Q%r�w�s}�s�=��P+X�Qb����q�U
ڗIL�TP�Qh�*T�j�6��V�E�Z"(���kA�������AKj���H���J�"E*V���[E�uI�hAVZ�
�h������T�D���
ֲ��H�%e\����(9VZ�6��@��D���fSL�RbTKeR��MdS(��V��+ ,*
Q�V��*J̴��)4��b�-e��}¾���_��.U����͛����v��0a�˾�w�#�0�߽gs�M���	���ߊ�}+V/�U0�f���9}��m��Ÿˋ��]"&28ّB����σ�#K�Xj�-')����ĸLz�C�r�x�?V� ި0JZ�IH��6Q�o;�n��%�%Լ�)�M�WW�x<��g�["�:4��5�v�ʗ.vj��D�3���R�"��d
�냷a��WΥ'YH�C��b��`��_i�F�hF������=�
mYޕ7�ı��O��^>������1B�]۫������mW'�!0�p��&=�����OEt?n
���Hrٙ[gJo�	q*L㬘�J|�ׂ��u��\6Z��o �g�{�7z�bt�O)�c�e���
���P��֬�[5=���D�3[�n�S2�׆ӵN@�롬��Nuh��&oz�籎��u{��99�_ved�3��B9WS���ͷ�����J��J�Ο��o��7/�Iۘb����'^Yfy@���h �7U`�1�ެ_> +83N��{mw�f�]�A.Ԓ��R����q����<��^��v%��P���m2=���s�)$�:T���ET>ˁ9$Myۼ�!�z���T�O=%�-��+�(�Y��(60=J��<����,�<�	��xn,;.���װ�,qQ�fdR�f�묘:��V��@]>����"���ԩ.��Eڪ"^SV�Y���n^1�,n�<�
T�hٱ֊�!�F2:���\�#{�S\??r�Oҽ���#�t'�ڙ�����`��g��67�d#��*�W�uxS�ݗ���W��s�:dc:u2��s**�hP³&�ïw)�:�UZ�.���4�-���E�q�e*̽���S��s�o1���Y���P�$���6�Z���S̫���/�M�r;��;q�m�����?E�є��8���ΐ��H�� Vw�g���� ��%��JT��JD������tg m䭧�ذ��!������"h?y�5�ϗ��ʴ8x_���4��fo^�;��� L:v��ɞ�BVA��#�b�W�i�+�j#V�h�q���g�֩4�SM(pV��V�X}�
|j�P���_ˤ�\����W��T��X_3��ݨ*q���|�_����N�������eH~���0{�S�gt�8��`I��i��N����I�yH�Uت�v*�iك	��3�@>�x��%����Э
�u��D* ��4S'�ߓ�
�~�ֻ�{��{˄��V����p�Cv�(�EAL�C���EpZ�_��>����t�o�Fz'����}g�Bl�X��{V5-kyݶ���+��4���W�;��9J�ÑƼ��g�׬7R�2릱�.�{�z���m�ۮ�;dն5�	����~(K��XD�w�5Dz�f��� �
��T�t`�9�1W�R��nd&l!7��o-�=S���	�hyG�KE ���!��)���#���{��R����������(@+֩�v�uH4m�cǤ��;���(.��g�֟
��ߍyMu�P�J�Lۼ���*�w��N�`�=f���7k��ȺƩ�O$Ms$9ʮ��~|+	�p���x�!����Z ��J��u9�]�7/��r��`�1��66��L�w���Л
]X)�C�S����j��bP0�l>:/����_��%di�[�N���L�>�/�+�|���
?u�t��e��|�O��n��G����.vgm�ueG��2Q<�������:�%ټ�|�^�l��߫ȧ{�����K�tt�P�F`���e��O]���ܱ���h���..XуF��P�D`2M�۞�'�x�a�L��7jxҜ��Nջ\:���n�X��J�'�~���ϋ��7�0��[ز����!K��1�2������)x�:<�#��mE��;���Yt�1y#���F}x*��6�LՀP���F}mx�#���W�x��\8j�粮V�i�lJaC��A׎�|ˌr���Ѧw�.����DK@z��4��R�Ӗ)GE]��d5��b�־[<�E��>�\>�*ʇF�y*�U�w7���l$P<��a�
���k�p�8Љ3&�������K�K�H=��Jx��>8�pG�n���>��@�wbm�'�r7w��#�����	�)�j��vv���R���{�;�aCj�΅C;�{�����"_�{���>��?	Y��������2+�� s�oz�;1��3�0x�6yT�E��u��㓰-�]v�֤��w�*��|��5�p���ׂ�5�EO���No}�D{�A��*����A�5G����|*]l�Rq�W/�����dp�3�o�BqP�Rg'�;�3�ݳ=�r*�޿`ᢑ��V@*.����s�BgF٫r��6.n�O2��Hh�^�tU�~�Q1׏�R�Z��Yv���ΐ�w�̊�5�F���IW�U�=��f��i���n�չ�Q.uq���	�LA�M��R&�g�3�׃�)��}��u��?0�K�{t�V .ڸg+*Ӝ��Z��cUZh�Ao��ER�Ɂ��[å�%�&��;,q�|v��1���J��.�\�.+W;�gV�M�滺�LJ��uuq+���V���!
g�ȾܼEO\��zV-���v�ׅ~UX����F���Q�%�h�0�fc�c������|��=��k=u�.���N
���"�;}'7~�É�}�Qhu�Ƭ���p� �i]ez$㝄Y _�m�B*�-*Y��ʕM�L�;���M�ٲi0�y�H@X��X�Qc�n,>5+��؍f`��[�0]א��U�a�\�d=oN%N>|�y�^9�Z�{7:��r$�p�ĺJj�V]L�WsiO]zU]!Zq��o��TV�=R-��)��/p�!Q��g��j��_��qGp��"xV	ƕ8� F��c�X�5BQO�E �,������]����3�*����{�:0�#���~5��Ia����e���:�u��w)4E�;�Ƨf�4����t��o޵�����T�������B\�F�t����{<l�R�B�����Զ�pL�qU.�VM;0cK�� =W��������66�y�W�z�
3��wsEo�;ۤ7���98��c�~VCQ5b�O
�<6���_��pK�E�\K��Y\\c�T��κ���"�)ʜB�r&��`�W��>O;��YC�r��]h��Ym.��`�c�ȩ"�GB䚋rvT�KS5�?Z��dq����/�W�V�ve�������D�k��w�L�V�2]���0e�]e����@"�y���,T���n�Bi5�(s�E��uxW���p^<)V����SUv���H���"��TN����@P�1�>�x�l���{wmVF��7&}ݲ��+8lU�:�m;�Є@�8+�Ӗ%���������]N�v�1k�����zĳ�4���Ѥ+�UV ;بjf�xY�����).�E*���IuIh����V���U�X�!f��x��(0m��:g+�â�5u�mӻ_x���oyz"�sǮ�Èz��kV��E�5�-���|(�up<2� (��҇P�,��.mTf�xm�Фh�;��O�z)�[a�ڶ�=���_p����𱂥�*�c�0_"�e�j����B����ǅz���V�H�1ӄ�+�����7�0��u�_�ie�����$e�y�5���L[^͗����f�� @ɱ�`?M|�cY���N�h��*Ћ��۾L!�i�
b�궍Հ:�ױhb��h�6���������i����=xz�qͺ�^�ŧ�wQ��P*М@gOr�������c�����7�o�J�P��.ݛ��Q8��f���ۗ}W68��W��1�"\�ܤ☙N��Q�P}z��)j� ?[��C��6wzz�_���F4�p!���X�J�u�}1=T锹�T�+;	e�d8j�s�Y�4A�IV thy���x���ܺ8��߰^���U�>��o���S
Lʨ�3"�����m4�����#����ʹ��J��:�C�a�kM��3����<������f%x��Pxh�F2�m��Ft�������In�+����`��3(��X�F�UNJ�b��nB�pf�d�j�i�)�c�j�k��?hT*"碮N۳��h.�m3�Ԧ4R��~B����8kz�lߕz������:4���\�Lv���L@8xg���l-�Õ}�����Z���E�Ҳ��H�[3��������c'��>��ئ+2^9bw����Uwʕ] �*�K]q�U����t������Fܙ�주+�W|ۉ���YaWT�b��k�%�ͽ��RU��LrB���=�{<���<���������tX�R�r�q3�sc�z�)�$v��XK�M�y���v�`�檖 �w&J�4z�X�\�Rmgn@�QE������}z���d�E�3q����*��sgt�ej48��,�
�Ş*,5��u�#7�g��S*>]w6�{�)���,�`*�=Q�\�k���[Y�Cy� �uq曫�7|��K�Ƿgo/b������S�������әdTU8&�ocE�s���
uXw�,�n�\���G��S�}f�3�v� ބ�a�p�n]�N�x���40�A7��
��!�ֵ�[�^��(>C�%Nyr�X+O!&�j����o,U�ɇu���� �b�4���r�ޥ�,,��>� Z4j���QuCrT�(�p�+�
�4�iP�j@������n����k9x�>L&��,b��vFJwQJ;��6]a�$�w/)r:y[�J"�"�+jQ��u �eb�k*�i�5dթL+K�r�M����B���Z4nQ�A1B��	�仦m}	!9�ے�P�n��H/���x�w��4N=u���:�Cㄌ�z����>����b%$X锃t�GJ��.�����Wl˺��ƪ�4�m[�=8l^�f�f�,.�����ʅ�Y��M9��jP���M9�*�Zے��!4 ��fҸHo����!�~7#��8pP�דp195|9�oe�V��X��Z�I�#�Ī�FA�9=�Y�""�@���B)+%��	Z�"H��	֬���V�(,�
dR��E-%`��V�X�U�YI��QaCTi
��چ�L�&�a���9l�kY�Eąb¤
ņ!Ke@�RTY1.R��jT��Y�L��aF���)�YqCqA��1T)e�,�Q�J[V
E*[h���XM5���E��AVAjB���7�8���5ўL�=k{�󯞡���:!�)uX��\��!�t:���JN�oc��7�N�o��5����ٌ�AE܊C��M��#��������@+�Y��6�Y~x.���g������H[)�W�Ng/��çbvr�f�iW3X�U���8to���7�i�'Z�l����__�Ei�R
�go���PYHx��G'i����ʖӣ̡i�_m*8p 0��gbw�/ݛ�lw�A@T���T~
��5J\���n,T��-:l��]ќȱ�k�ִrEz����e�)��O��ǣ�)o��(0+�hG0u���X%����=E|}˃�O��%QX����HRA�&Ѡ6/�?���yP{�Q����\\p���93�,ɉ���3Q`!?*\׆�+};�<m�ٮ�x�F�R� 0:/ǂz�h�ؕ8X���%��0�����{]g��Ue���
-���+3��ϳ�l�5ܚ��ӍIr�fN�9^~}F�z��۞�e��(~RE[�B�T5b�},VS����\:�Yg� B;�d�Ѫo�`�������W&|g|r���q�b����͑,�TL���S'G�Ʈ�cF=ŊQlQ��/4.a<1�W%��ξ�U�*��£sP�p�C����cZ�NVvU��W�Nh!dL2ppu�ʕ?(�f�ݝ�z[$(����-��q�[������C ;׮_t��ך��`�4r�?m�luӪA1�@+��Q�B�T��-U���n�M
2��;1­W��4pp�F�j�?v�(��n��PP���>��q����]~�F��2E\�_L���;�wm幋1^S�k@��}�/_�41ڄ�����K݉���x�}Ɵ(�G�V4e�2�2o���A(a���Z���&��j�:���x����.�K	rn��|8�;���ӓ;��6W�69�f�����k��J�ρu�� �Mw�':
m�[��.����A\�K���U<��{=t�x���B�]KLT�<$a�V������ybc�7�R�C�"o�r&e!jaL#�Ә=�!t��ϳ�z%�L�Q*����'�̫뉖jdτ���d��� VpW�b���]q���+Z)���l�@�*&�g����XC���V���^	�u�V{MKۧ[� }�W�R��f�S
���b��j�0kJ<.mQ�R����AV�)��¨:��u�im
��?����l�:��2�A�-���nfv|5�HjC��0$��`ٙ�
�jp�*y4�G
����6L�\v�<T2���Y�cc ������U�hĪ����:�}�3���W�gt� 9wc��zw�[G|7�95�}�w�Sb��"��ۋu3�h��^K���	|�>86
�N��׫_'��z���~59T}��K��>�~2��y��K}��Iyh����A~��=5�zp/���(b?*+GJы�pԾ�"��4�ًU
\������Y����>f��]9x�q�dط)���u��ʹN��n��̨
�Lҧ8k�+�����FJ� TL��캣8�1��Z+�W�e,&��!t9�|w�ʓ��@��*ς
J��ǆ�<�)��|J�Y]�Ç���
6"2�J�E>5�B��B�Y�����w����Hhв���b1k|���x]YC�r��K%�����{��hp�}Z���h��LG��@����0��S"���ܽ7F��D"N�;Os^�#js���ufW�7�y��b4j+J֪ǫ�`�4����Mr":w���N<������]1 Iވ�6np��~�G���6'&�����f��aNQ0�O�RQwyVL!#"� �s�<�D2ceJ��2�l���=v�ec��1���x�}z��V�J�"�T8��3�]fc���
���Ƕx]Pcy`�K���"_"�X|�Yӱus
c�)��s=�$є �Lt�0��qh�X�g_�V�:�L2tWq��V�<%՞�<3r� ��ɩV��3Y��&D�F�_-\=h4�C�B��p�37d��N[kY�ݫ%�1�(���? ��vfzD��&)6��e�!P�.���n��Ҩ'�b�
�(��Ww���B�7�Rb�K�}.d��]�ΪRߺT����&`�M��FNO_0�3E����ix(|<Y�-r�=^��<xrk���bT�h1�K��6{�n�ܤ��S"*�~l�ٛlJ^u4��vL�c�n��qm���]R��f��<�88�R%D^N�w�������a�9��u��`4D8�3�%r�*kEV{�B�t�}��:_{�hCX�RH`t>�VO�5@Q`����F8�[��͠=�Ulj���,�
���(�Z��,�!���N���7]���a�(�Tk��>��p�`�K�&�D��N�a�50��8��skdK�s(�N;jj�VL�Ş�x���UK�]\�«'�R?�4�Z,�H�{��Hz~�*az#�Μ���koN��\(+-�k���T�\)���Ɓ�߱h�3�탄��b�EZ���lQ�j�JJ��k8��}}V.�8��	���=���������޻�N&88{���U�Z��Υ���T��w�M�{c$5Q�J��V-�.��}�O\�sF��[��D>�│J��>��
s�/ky��-`B�ݙB��IJ������糥`�Y)>��rڼS;F�F
���J�=�ŉuĝ�N�	�Ͼ����jZ���ڟ���k<dɺn�� ���t� K2��O!,\��	���x�1S�^š}��S8m�
��Gmm��x#Tt��D�Qu�dK�t��Ɏ��)N\�i�#Y/��V(#V<�C���K�<U�c�6��_��I�k�s�ta=f��C����(]�>z*[��Ʋ����6s1���0zͮU�x->����Ы�pu�lsK�T��.�{N+&{ܣ�K˻w���S�t���$ҫ�~'x$�{y�veX�4TX=B�xJh��pׅp�;��R�/�1e��:^�OM:%��i
ќi���+T�j�3F��d�g�*�^���M`�qW��7�Q�xV��j��~�ӝ��������g���P�)m�	m�򃅋�-��?D/1{+h��}\e�MnȝFc�3��zgj�[h��~ ��[8.���Y��}���n����,�N,�p������VUt�g�n�_\�e�l��[[
�F��C��S��]�PW�Z����GWIu���06�>�="K�S�[Wk�uƥ��EHR�l�3ެa`,&e�R�T�33q��1�	;jm��NH��LrVʤ��Y��b����.r����-���F����u�+Zw��0���o�pc�(���
��j�b#�Li��{��Y�d�"wp�ܫÆ� 0n�G�y䭼�����kh�^b�f��uC�1q����6u�r��
�ؗ�C�J]�Fi��T�s��v��\�P�_�T���X�ºW�&�L�����1Y��DA薅��0����bҫ;�l����`���s��%"�o�S�J���C�^���r�+����RT�o����'������6���� 3o��9�Юut)����r������M�[���]
�
\���;,{�<H*�iÆq��J҃Yʼ��������Ua�x�>X�J=�h��4p��p��5{Jn�*W�
D����p���;9�||#�1PQ�{9��a�a �QѾ h��R�
���e�	q����x��sCk�6�p�&]� �����S���"k�mn�v�9��jŵ�M���h׊�\�c��u��<���?(>f.�0{͕xp�G4�'�a�[x�,U�<�����s��o������V��
w���h��\���|!��A)�.1R� �2&���̙���:�[ńݞ�	M^��w��ປ7!ّ50l�v��A��g!�d�sϹ�~��-W2��on�ڞ��U}�i�_AҘ�J�Z(��M�S)<�n3���p�u��m�=cz3)�3���c�V�q&�W��U��o�۵�����CI�j��!H�����[;ꮑ;��ümNܹ�-S��>�F���ƕA8u��a��]��섕"<�������\b^xe�uJ�oZ����dړ��sn��P6�l\�{h�Yְ�<�.U��zD�Õ������K�ޜq���\5S��⿙�2/�:�C���Ug��� �	�~˾��0�����*���5v>:]�:�GG&��r�D���k<<�4pk��p�V���g.>���`���v��#�� � W�*U�1"dѪr�ƛS���$+x� H!@�����0���Dv�~>�jWEnfP�g$�����P�5>m�fR�09��H?h�����j���J.�h+gٰG��i�_f�
�Y##���.����ך���kkq�H�r����w]٬c�e:�Dj��G7���goL$
��n�riy]������yZ,p�>WI���\a�����[�Q���-]CPKԗ;�Ps:(�J+V�J���{�%lQv:�m(h��Pދ:]le堑Ի�� �!{��ְ��ܚ�e$�ҖrSʝvp><�д�˥MXQ���Y�g:&j�JNX�2�^f_m4ž�����5��gNnC%G]:�΢�����67�]���ǸY�;�K��Wn����8�!����ά�.�܆J�X�TGr:�^���?C�s�L̡y}��=�w!��u��N�Y&����-���>����
ˢ�a�+F�<n�K�[X������iE|+h=�A[�	���X�ͦ�|�l��X+�U��Z<t��%�:�"���h����9Y�R����!����S�!8�|���y�`��W)o�̺i*Ö,ZA��pB��䅃(�������.D_Y�V�y&��$TF����Ww@KNPwX�%�@��#O&+�L8�:̳a�#�M�X���^e�5��d�a��$Y]TBm��vwY�L®wnY.7V���eZ��ذ���әb�� 8*ŏ(�2���!I��I�(�NCf��W�"�%aH��U
�ZN/�)n8h��+yb�e�]�>00�XJ:�����Qn�1[����n��etz��e��V��ri�8W= dD�-s�x�t㏄)|���uc]3��N]�]n��2p0��T�ͷF�ۉ����{��׮�h�
ώ��n h�@`_*��</�����-u�RsY����_e��E��s�����RE��ƨ�}.,�D*{��,��C��AE��8�Lef��0���FJ��XT��"��IyL�U�b��H�%�*��Y���"����@Y"E���++%`(i�.��)����1�\�"���u�EX��@�# �̋P�i*��
�Z�k+�S"�%AA)�f[1+
�ch��6�B�SC��E�Z��Q��Im�Im�>!�|�}�"�.��y�>���m>*��2��u�� V���T��0��z#-��k�B�g�N�22��dqyW*c])FdU��ɉ�-��"�W��U����V`�`Y�X3��(�:{u�������A��W/Ϲ����kת
��e ,h���;6��S��c�6���~W�}���T#5$�hu��iZ�{5�,p��x�����h��;�V���pt
����3}ܳ �M�,yj����
ukβz���힕'���L��$��ܜqQ�)t �{���|x!�<k׋B�sTq�x1鉏�m�Z8:�4F��]\���2-����M1��DH��v&0]�@��\5��m /O�tkF2<k�z����JX�{���U1Ω�v�7OZ��p�;>K�hg��yc
��d�:+�*J<��3�4^�;�'#)�ڷ�JN�Wt�tzCc-�kZ�6��3T���tp�o/�
��Z���(qI��ޥ՜յ������G�c��ߜ�O=�r������$��kF����T7�/���Bឤ��*.ׅЯ
�i���+hv����I�V�b-�<������QsL:̮�B�̡�Ƒ��ρ������w�65����R��a/���~^z�����h�m0p����]����e)��@�8:�V ��ŢÍV���<�י��_�@�^�Z.�ýT��:ɇ���t�������|2k%� [B��p����½��U�Z���^EJ� ������^{mq��E[���Z��k�Ė�9���ҕj_��ګ��
"Hߋ��=@`�ѳW<<3H�$����Aw�Sge�)y�=51|n��UGu��į]o+��`�Z/4r9�|=R�)j�-�]��؃>mA^�ԩ���2��+h᥹DqV�ÝY{�&��i�I���:�ㄵ��l
�x�uZ��圌�Q���{�e��X�~^0�*�Xt6 ��GQ�Q璴�U��ZY���'��Y�=u�N�0�=�7�K�t����ĺ�R��_�����b�8<���h����|��3ƺ��@�`U�'��v��`&,V���aF��{��[E�孤x��(-Ū���n��)S;FTu9��s�Ww�iJ�e��)Ѵ{�E���GG�-N��W����U����	�y�w
$h���oU� ���{�"phe5a��v������R&�W%���\��|	��B��T�x v�|���h��$�uʠ`^�'u��5�U��}ʬ�<ti5�i��x}��ڢ�I Wt	oog7.-u�=[.\�j�*z����qYױ�m�8����vv��j�X��|�\Gt���G`k"��ޅT�6{�n�P�췹y�XE���4�	���]/��K{9�v5��Ly�k�6gK��4{�?@�DfDཱུ�R�h�b�`�g�����H�2��w��ō��s��E[�¦�2Z�tt�z6L�\=�^��K�r�Ȏ]ܺھ��H�� ����s��%�no��0�)2��!���۶E>
��M5,=�T����5�Y��sx�b�O%��|ФF�h����΅�6����h`����3F���E�_�������/�ga�%*�5�|T����<�:�\'�ؕX_N\0}�F��:W�O_nw#����F���0���c��q{�yUj�=��{A�[��0.kd�r��%R���(]ɞ�w댡9>ؼn��Ʒ�@T:tU�\�<<:4�0A���|� �X ������W���� s�f�s��!��ך�R! ޲Q��]��%�p@��vv��.��&�͕w;����$�M��P�A��O���+#���U�ב3��\�s�����8h�2����d*��ufwowF��u���k@4���F�'Å������u��5z�P���G����������I���j�-S�g��K�ޗ���/V�Ze�}>�*b#��mNC����i�w0&�J%��ܤ�򨍎}��~9�V��N�����atk���z������Θݨ�B_WLb
���y�N�	t=/��g��|.��wg*�uY|�O]������,/�LdU	S[z��0-ݮ,��T3p���z���㪛�a0�5O�)U��v��	�Z=NLU2�*j���+�j�ӟ��s��X㭩�=�8#^l��2�X/,����j�����S��:rw)v",0O)�U���6im>���i��+�@��δ��;E��5�����9�dPl��G�m�r����Ȫ=�۔Eݭ���9X��?��m�����~E��׬Պ$�
��|p\w�b�7.u�>׻��r�ʖi	B�5T\8m
�4^�����D��V�o�|�9Z�X�(�`�Ѫ�2^�C]yp����@�?`��5:�u��U��\;�R5<O��o����U���u|�Zo��}'�^�t0W�mYt6������d�5V*[��{� ���F���O-j�����n
ŝz��EG///����V��y�/�3�	���s�[�-U��{�[5�x�xADn:u;��)z�[�Ws��������-��U��)�n;s�H�Y6*�H����$ �����p�W(�C�g+��1/m��'E1&��^�N���k8VR���>�U��
�ࡱ�{����wF�6=�;z�*���dm����S����JP��m7�e�YB��0��fv�O��ԓ�ܳg��Ġ���}(�rt=F�I�l.�A�R]Mt�jԩx�9�{hJSFa��q�-�UՂ*�_��IL`�X ���ʱ���x*�#mJu�%��`i<S�O�Pl��8�_Z@��s�4�a��#ݚ=<KSjT�Ve�u�;�W1@��O�� ���<47��D�wBiw�*b�gU9B��C�sf�ʮ��$E�:m�w�0�����Ffc&��M����b\���C.�������H�� �GG�p�pg��F�s��~U������c��#&S���Ș��+���&�#��G��V9���>��UGt��J��\j<��\�s�WpgD��4k3�J���5���y*�C�ZN$(e(�S�
��9f�E+�霸oj��p�+�@�d���sV�X7�.Ɔ�X5�Ls��Q�	�];wVK ��`8��r��Fѻ	��
�Gp� ֩���[I.]]���2v��kk�dp�"�'a�>k�Y�G��s�
��U�g@^Z(��!Z/qc<~��t+�׭�({�*�� ��x��
јlkI�<�>���ۺ){V�2��`�>_nE��zK8N,T�<��W��o����U�Wy@�T�֍���xJx�FmV��Z�n�|XGO]{X�����}	sʓK�^��hT���[�QJ/w�X��xe���ĳ�X��q����s:)I�2b^&�{6��S��sҍ)��p$��깙3	W�����c����e����[�\]��J�Gs5��h�E`cI��P���>�荨}B�\p�V��T�MO%�,�D*|�
�^�͖�˗U�%�9�r��>�KK��j\�/�7���!��y&���Z��C�l�3����F�t��G�h�9�p�40�I#xs����L��fS�� X i���x�]��]�֝�s�����̭~6��«9�&	g�=~��'/^�w$��O����A��5�:TB���Wd����_y�??qf�aV��ѯ]c���g����ⵛ�H�i(Eq��U��M�X���njt��ȪW-�����E����q;�i]��i6�B-�5��|sӎ�m�j{� 8�3T��^Z���O���Vp�)�},挵i^Ƣ�g]�8������,��m��A�a��[���E������I��w���{�4&��g�P��Jxs*J2穊��*k
�ǡw'\ٍ�%r}�(ԾŜ��t[=N�2ԓ/���:��B��1��8�]v2-ὼ���8��
v�[;˔l���Xܝ�Ǉ�/,6���;	�g]��	�Vy�Q������}Hx�#�Q��w���;W��_w%�]�iz{��b��=��)r}��oo�򡍐W�����'2�'`hD緱��6��η�tL-�Rbp8kBCJ�J� �U ��H�B�	%)�Qw��R{�F����++���c	I��]E�+�%:�HI(�;{u�<�'y���\Q�B���j�k'�(T���:��4�jE=��/C�ө���pޝ�-�ٔ���iٷ�
x�riʹlZX��2a�Ki.�h�Ca��C�;��4��Gk`}K~���F����͌]wqG���f�x
� �/�Wu`�Å��w*�Y�|�&(f��2��3���S�¯�g��e��E�Y�9-ᔊ�'���w�[�v�����H
��L��ھ��칗��	��W��4ncL��{���x��p�u)��Q��!����E�|+�y�fs㸢ޕ�C�\=�T=#����6����11�����ɪֲH��s��3��)�u�l�d��m�-J5.���r��ҩ��Æwgg��
�����@��L���Q�z�0�UЖ:ps��raM�=Ӱp�,[2B&ֻG��u����m��뼾�ۑS�',{�T:��f�'zM��Z-9 �o�����.\F��L�5�օ��wqΠ�������=���K9\�4�S_^�I�u�C�>�k�����K@.�$��;h��mah�/�J���S������
׊��,���O�7�6�G)YdEc(<�G�e5��&�VKo4P�pU��wH+E7�[�aۡF�K�o��������.ٽ�%��fݷe+��&�SF�.��%�J�͵Յ�Ұ�K1�����$��옷j�^�)dQy��LQ�Jf#a��ǘSTh���$��.�d���6�����m���ի���E�"�๿E�M��eϜ�[���R�k�b���6��x6h�-�uU����V�t���M����au��z;�\�v��NsGgD�sIVEځh%[�ƣ�im+�+�d�ғ5CzӀVQ��i*AUa�VVW-<ar�`i1"�Ur��P�s
�J�Ʀ1DV �&eU`��՘���`��N�����@Y
�Y+%j��a��[%��egL*c%Ձ�G�LV��hLk��Jŀb@�iĕ"(�YD�DB�E���q�,S)b�TdYX�-T\Z�t���4�1E�M��.P�S�@��4�8���hVEr[�1�(bbACA]Xb)�n�&�gNj�%�L���5��R:��AH�:h�*�`�9���:-}��8�v�c���q.M����os��S�wy�r�h{U3^}k#h���'�"�)�s G@v�p�J��sR�j"-v��8�������g�j�nu�:������S�Z��.)�Cv�^����F��[Vyo%vL��,ꘘ�+��V�՛S<w�N��!������+K����-��~	�5�h�[��u�����b��h�w�:�f�hȚ=�:k����<�͵=^3���,r(ʥ��7�)G��kYG�hO^.��0�#V~���2A�լގwa�6����:�*�5j�ې��ەx���CE��/��>�^������Nn�������2a-�+��nu�u;z�e�Àc�:e%8ٹ�7`���V=�}�����l�_[�9��β��޹<����T� �T3�p�܍�����N�"Y�j��Ү5�חץ��EES�O-\��i����7b�H�a��g��_s���K9F�h���g/�X��	n�b[08C&�]���8��qng46Y��{�^�=+�m'7� �����4���c�ђ�(�,���&��\��^����iRR4]p}dj���oc�y��S��:�	����,7%*=y|]�ϖ^�϶��b�WR�fxǚ@����G�o8 'ngڒh��DaݣnWn�NCt*�<Al6���.�Jf�k7IDޤ����-�g���1���A��HևȮ�SX�������dt���K��7id��X3pѸ�q��@���ٜ�M�Қ���:��(pǋ_u�+@F��+Ev��4���Glg��fѧڗg�ͥ�
y��Rq�u�k�����U�q�`�x��Օ�~�b���]T�b�b4̈��z�rK�e����^ak�U
��T��֨+�U:�Zf�Ϗ��T�Չ�=!�1�W��U����V����
9 �ixA3�1S�p_r��E�t��� +�b�H�j���v�V�~���>�ҳ��R,^_7�����]Q+6����s��uYp�u���]��i����݃��-U��|}�g�at΢K����o�t�P�Y��g�O�Y��ti㏻�"���Ӑ[s����Md3��	1G�k �y���M�]TR�v��l.	��� 1�6����v@�Pчz��A�Q�Ov.�u�|q%�I]�b�#�:ͺ򭸦�&�m�/Bžc� �f�n���f<-��8r�]r��[��Q� �iW���XM�ʝ�+d�<4��������t��g�\�U��s��%Զ0VR>��t���������naW�j�Cw��TN�I'�q��=Σ��G�i�/�4'Vw?���u5�
�r5au.���}v63�}��ֶË������yk!������"�R��8ŉ�nE^<qI.��'"r������d��-.?-�[Q��� �kx��k�ҽprY���Ԫ$F����T5�I�=��&�Tc����EnM���[[>]$�M�h�%���3�$Ac��h�\������uh��)�f��]���YP��z)d;7w����Y�����vվ�M����a����������
l���#Z={�r�>���Hf-5���E���ul���,R'�m:��Թ�ۼ`�������Y/J�*�=ҵ��E�z��l��A8h^��{,ܼ�>�2#ip��k����ܨ0Ts��Sz��ީ��3��!K�vǌ�����_�	��V�b��_H�=�|���˃F&Ӌħ��ܾ�Ƀg��>hf ��oJ�l\��G����Ƶv�q��YL�N�Hz��U�;"5Ʀ��H�����DT�,���t:��i�9ф�����M�(�a;i�sѴn��k �z����Ps@��ȵs�+���6g%Ч�0cg9o��;�t�I�$�Z�_���	Xb��ɡM8���`��衱�Μ���ɩm�;c6�,�5��v!�S�Ã�.-J�*7�|1)�pKi���Ae��X�#�iՏ_���~�cC��/��p����R�k��Bus��UvsI�眸пt��z�ۮF�U���ԋ��M�=_g(�G��_�'�]�+P܉�q���U#0���ͧ������j�USڋ%M�h�q�F�����.:*��㉉��e������\V#&�>�u�vp�6�lLu�)��qz̒�U�)��'���u�����t��^�-�"<�w��w\	⽵�m*4- �tu8ܻ�S����6���y���V	iE[7a�"4gH���m���{�1�Ht�䝫��x �v��E#��t%�)ѢR��iGp�<����2��p�c�l��vg#��[�����ɐ�5u�v	%�/��nq����{��<j��q�����e+=�o^�A��ꧾ"/�� f�kX���G����"����j4g���0�20�\I�@� ��∞��5{F���kM5�k�
x�iLuˌU��DգH����Y;e��,m,�[�z���g�D�����a�4P�Z]n��+��a}��-�|s:UԱ��J�V �LQ�|*��s�q��Kalܗxx���S�D�F#V�tV߆Ǜ�2�C����N'Z�[����~`߆�[�ۏp�[}��k6ݗ�?_$�ިJ�����g*�s�zfDJ���tG��!��L�g�)5[ħ<��re���y�$wi�����͍L���vq/ЊC���Vc���s����F�����@e(�$$�iTΜ26���n�n�f�U�J��Tr���(<�W`����zNL�cxY1�� s���(�㛘�<<�	����d=��ԝh�b76rj��������2*��Vz0-�Eΐ���"y�3�.�y-+wjJ~>����ۓ�;��>�"J������k"��7E�"�S{D!W��n�"���ȯZ!՗�Rԙco��r0i�f�S����%�*���ӾY�)��{-ֳ�z���(ˢyCu�&�ok�Dng�kA�rN�o�ViI��[}�VWQ�
њ0��Y�EL֠���(�d�+����uMC�rPI�7K���#��EBy�0�n����Ճ���PA	&�z��=�bֻ��tv4P�kJ-��˷�F�����d��EQ<-`�^�����c��O
� �%Vc�
8k*������b�P��u1�FQC+t)�;��L�]8�)Y�Ƕx����M�	��\Ѽi���w���`�;:�Fq�"�� �������f;|�n#-����Wm�4Yeak,[,5|�Z[��FS�f�æ�{�q��RB�H�������p�) a��<��:�M�<ۦ[���8��5[�a�S�w�л�\�V���Z9�v�`���Y"{���횆"�mcJ���\��Qh���d����)������&��.M5>�&�����t���-��5��T���a坒6���*ҹ!�Y���tI�b�5��]�����n���+����r�#zU������WʫX� '�u�m�^�:���g���P���SE9@�w�oANM�u�Fb쭻�+m��,�v�SBx��[Q�<� �� =�7UY�	��pY��m��5,�D˴4�ftN���A�Wk*ݥEk��vM��l�L�r��Ч�dcxs���� ���õx,0~݈*V�X��kj�����5��B�9@}F8��3q%8��T����`�H�
�G^�WP[����h�b�,�Q:�f�mc�iit̥��Ѓ+��"�,	`7��:CwmV!�g���9��t�Z�/�P�%�V.��ԯ�����S�*�r���nI��@���5Nm�*�f��U�
�����l�%��I]#���o����^N@e4��V$�h���Ϫwp5�a�$�zMgV�M䕌��k4��g�#N�4���nm/����
�+F�t�z��7c��[�+��J��	BTͩx��E]Ƥx���ᝳ�k��v��[3��OoZU��ݖ�A��8	Ϩd���l����m��B��t�$ά�y�*��Ԅ- �'�q̦j 5T�Ʉ�E�����1{�JؚIMW���W|l���WJ�@�F�D�9�a侫�"��+z��#W�rn�n��)�B�Q1�N�Ժ��гb��u��&��]�����؊9J
zQ -	-�w��[�*�ײ�$b�Y���m���]�P $� 
1�q�1y��H�c�.�#4�����Zܠ��L%�",n��I����R����B�u�2�$Sc��1�H�8�b�L�ĕ��J�1E�uLE1�IAf������5��
����QPSQS����1�]R�-�� �Ɩ)�b��m-˄X(�J�Ld�
���Lb�r�+r�2�%���t�t��b�YP�[CYAzJ���.�`�.Z1D�Z���em)X�[LDaTeB�t�A���h��@p{���V���x�{B�� ="�[��5lel��C¦��FC��w7�V��nY�X�5Y.�1"�[L۠l&Z4ə�j�9�'h�F��u5<�8�aT���q���08�ap1^f�B/���פq��F�Ҷv d��p�.Ԥ�Xק���5�:2	��:�t���{��x�=��+R���\��Ἃ��G9�cOe8�3���F�S�MH�Z��#L*�	a�5�q7�!s�k0uS�;�����<)�qz{�۞~/�Ϙx#�!��G5������x��Pu�l�:�|�6]nd��]R�ݙ32�FGBP����82X>X��){ë����"�mZ��省_mIoA��cP���ٽ�[Ŏ'3:�׼q<;]�;�����Κ&[��u���.'�ڜ���ѐ:;Mt�	[�Q����ᨵ<ox>��ۓ�ѐ�f���8��e���S�20��D��f����mq}�']���M�(鎚�g-����_d�u
3��<D�g
@�&��7�|��t���<��y���Z&ټq�K���6+L�r=z��t�e@�Ʉ�h��ڞr�=�ղ�Kw��m�[�N& 6	��vhȧN�/v�	(\EL�쳾�r?k��LX=�vZ0�Z:Z�.]M謆�O4-��b5�Ð��Ũ� �C3&<�xH�/_M����w6��X�	d3�N���.�%}�̈Q�c]����k�14l�:�۝|Q��u�q2�v�T��Q8T<w���lI7��^�6wm��4�Ȁ����9o�.����p�#�N>�
q�DkW:�m�z@.h���]GP�2(F�;B�3A�6i�QqD2���"��#b뮏EU�aL�v��	u�Qρ�d�_^է�)EW��h���0_�W�{l�k�ᄑB)tF����0Ŏ���gg��;y����933���|��c�nQy�j�߰+�WF�g���x#Cy���"�%u�����"U����{k����C/D��F�{�uv8�姚&'�󽺲vT�js���p�.C�_�Y��G�wr��v�S�S�n�_3[�����M�E�W5��%:k�W�_�����!*���VL����-%��d2�͉�B:�f�2�K�i�y:��*�*��$�"�v���NE��Xe����5L|�
���gh�z3�8U��mZj�h�n�nz��V-a�x]��y�[�Ɇq��oշq�H-Y�I�C=����.�8�:�j���d�9n�,�{8�����͓x��z���b�A��r��s��^�ހ�q��!A���]�z4WN$�Zx��Vh:my��3��>]�f�����8`�5Ҽ�I��7Qx)�u�R;�L��m�IAù��΁4�=W��oQ�fK<���b���N]�	f�j��*�aw1ܸ=�vw@�X.����.��t���(�u�dGt0��'5�zvQ�4���O���U��ٷa���4�NP�R5��D��F�=/M�Xu�"Ztѡ�ٛ��-��1qI��h�f6���)XJ��3�.�YYۆ��< 4�������b��q@��`�pr�^v�Y���j�m�i�1�	�b7Pw����S����9Z��E��k-u� o��1����&�.v&�{	��>vb�,ķ(^]�e�4{+��*����pοA0	^���^�ʽT]��M�f^���(a�T�5�S@Qo��,�-��vi�:��/{��/V"�y�{�$�W�vq"�3���U#�$U�8|/��ե��5�&f9K[Q��;��HsX+t����2�[�ސ���"����$�B�n7���֭�Ġ�@��sn�|�j����u��:�)L�a8���N]:^�ΐ�[�.��N���5px5ov�V׼�ԗ�Sv�>�8���@V5�yB"t_��6�k�\0D��~D��I뺃 �*�G����g����C	���c��v���%��η�q��$��	u2�����@E��a��݋�v���v:�K�'xл���.ˍ�7��gl�EԂ�I���'�I���`\��#Ss�I� �ޱ���t*�N�$v�����Gj���.{Fh�n�7}е8��U�\����Ȫv��n�Q-h�0�����7�!���K����q}%��_����NŚ��_}K6��}�x�h
t�0�&z0��s�-�}CC|;c�h<N8qЮ<u>��]��G�8�e����]e����"x*��/��h�x��=���A�j�ks��y��y/���:�'�Sb�_��@�#(ˠ�Mw29eռ+�tG�{�S�r����ٓ(3i���	�u�'����@��0y�n�E_��s�][Sr�/H1Q�{u�����1��V�iS��d4G���k���C��''P���]�Y���ZOd��È�SgF���4>BҎ�GTO)(�>���Zt&6�@��`���FȻf���r�uf�E�y�\�E��k�W���9�P�*�V_2���+�"�K�V��!�'�����E�62_E�d�[�}(�fgXE�{Abd�]��ёN�D�	��m�:�A^8���Y��	�d{���ǖ��A�Vձ��B�f'Rf0X[C5��7=ݪ�g�`ȩhh6���^�l� ���vk�ˣ�jt��w�}��u��gbD�CR�n&;��9��U�gC��I1g,�|#��7`���e��Ђ)h�3it��:��cNZ</6�6�%À�=�����c1 �i���#!b��
f�8�A�����q��l޻�&H��1�*Pظi��������
�PE�.��	��c�#������.�F�-�
b��&ʣ�����Vi��>���[k�c�!!��t8*�i�X�lã�m�W�=�Ѯ��TaS�/1ڝmLŗb$o�g�8��v�2rT���44�y��4iƣ�u�p��Y���\��r:�"�`�3����gټJ���̴T��M֥WS=�k<j֏{�1�xA��F���rb����,�����g\Yx`���[��[ǐ�S��_R�)�r��dx��a�Ӛ�I=o���t/���\���Ib�P�h�ڊ�Uhd��M�ԯw�}��Y��ޚ�i��t��h�zRSn1U�9�_9�l^f{���5sY/%Pfx2ڻ��t
�s��7��NӰȻ)+6��4�ڜW���+��>
o]�i��U��cB�x�h�J`�6t��?^��b�P�-���.9�]]*�G�S���E���'U�|!��+�T&�keb����+��9��d��Mz'A�o���=2M� ujp�����5�j�uW�s�t��+U�U��ZBI @Ɵ��*����28�*�|(  �5��X��?D)��Rfd����{���h�']��OD�T�H�$$.�P&Q@�DX>T��F��ޕ#�N����;d/�ļ��G6�3J%F�#9�~�
B
�!�@�i��Ƹۅt�� ������d��Il�J���
;� i��f�x�l�ģ<{��a�R��Ϣ&�/ڲ�P�e�*���P��!�W��2�\W��-��UA�B��"���"V�$��b㠙��� |lp?j�|��a���ލG�4b�'PC ���?Z �@A �U(���h��v�q^�}#`j�1�>�J���]r����5ٸ�	��|g�s���`�J1̉��T�PBv%��ƓB�R<��uAU*��p�@�i7DDcD���C2K��P+��ayp�_�ט��M�PCZ�K�&���M��y��0vx�)T�D1��*����Z�;�D?�ȩ�>�����x4���߬�reT�1���PM��SB� ~"�膿�����d��T��S�ȟG_B�;�P6�Q}��u��h�^�����͇4PCXd,a�˨` |C�Π``5�~@H��� d�e�E@D `��������)!=p/8���7�O�d3�\<�
��:�Ɣ D,�� �A'�2`�ZH�����"�  "��%
��@�xYj�x���dw��(��'��Bd����@Ѐ&Dż
Ը���}p�=��UAM��s;̀w��T��<���` ������cݚ�a��i�����������s.��xuD�q ��9:�BzS�Oإ��٦w��%T�tv�a�6�1 ̒s���#Ђ�J�J��0h!�S�!�2bt��X9�@hh'w}����`@ޡˤ�@A	Aid9�|<A:w�g`�覢��p����0�^8��i].�M,��S��]��.��ޑ@�xڤ&פ�kGM���!8BI�%�v���	H��vB0*�@���G��`�o��Ǩ�UT��� Xn��ǌ���b�"������C�JT�:$C
rX=����G-���rE8P�Oh�j