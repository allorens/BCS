BZh91AY&SYp����߀py����߰����aP��  �^�    �     �   � 0  @ �C�� )Ѡ ����@ l   � g�ƾ��l�{�� �  P (   (  ��� T��y���ᮍV@�O{��S�;m������mE�� ��� ��=��z*���t�}�կwy���ǭ��x��j�(w�:�xWk�rn���� Qy� �n�  ��7')˫�q=�{`��;�ڜ�{�6�]��ݝ^-���B��B�g��k��5�|� o�_,;�Z�aݧ]���6k���o,p�]�.٣��m��;g6:�p9�P��� ��`  :ĩݪ�s���ې9�o{���g6�@�: ��8�QGW��
4��3�-��+�w,k�n���we˻s:)�\�bڶsw,ù���K�(��  )A�%���ws�6��wudΎ\�p���ܺɝ��,�8�8	v�4>�
U�����`�:.2ۛ�H�nC������;�{��f�eKws��>�/` 0�  �m�f�6\;ܠ�n�����݇1�9�m��2g�Q�δ��s�9�Ʊuv���G�wq�\�L����                  	P�               >���ުJ���i� d��L�J��S	�2��F`M2`JmD#J�#!� ��0#`*j��R��z��H� 4  ѓCA�i�H�J��F�h�S$����T�2$OS$
�� ԥR<�2 ��hɐ�?!D?��D�����c����8{U�[������;a���a��6��}���`|�לe����_��������������~?����~nO���b�����v`[r>������r���� ����c$U�f,�GPN��/�~�W�ۜ�����ɿ�]8G}����R'�r�WD�Ҽ%���{ej�ܤM����exَ��V�,�6�"qܤLnWp��M^�����"u�D]��V�=���nW���-e'K�+M��5[���zR'q��f:�s�dM9���5�rI&Ò��^��T:E�K��'2'��u<vN7r���>��ʤ��5^<_Y]:v��ȍK=~�rt��l�R�Mx:HsR �O�%Y�j��V�Q�%�����d�ep�"#�+dߦ$��'$/q�G�ȱx��ӯj�&<����P�jr��suI�rI㬃�d�9"5:rDrxM��dߙU��dD��D�ʕ�n#��A�w$�쀎H>������J̞�'�����.	�sI!��{^Oi�<c�7zOu�K��u,r,�l�̝�%Uܪ�J����V�{��ro�#�u�%�����_u{)���^����Ud�%��r{�ޝ�q}W<�*�KR毪�8�XI����㶓�x��u'7�֧�z98L����S���$���k�G�5|s�G9M��5���"c�$�_�e��D��0���+�sXsI�:��}M�V�Na�;Z��*�����g�'�����I�\B�yag'��Iʒ��bFɳ�u�|Y6HC��$�e��hq95�L����{\9����<��$��2'zt�"c�l�OJ퐅�8�]jP�$������zf�q�\6:O�U�
ȔGQ0j"y�DN�Rı��dD��%�ŕ��Tᇞ�L�:�+��q���%�t"=���]6y�N�+H�J6�&DG���t���R#؉�>�Zuu*��r�:ܤE�]6U�H�R'<ʪ<Q�Q̕�Å�u�r�)�J�k4ԤM�)��"�V�V�>���nW���8����ҵZnR&�JD�2�l�S�+N�W�u8�R&7(���i�I�m�D먈���}��O�"oە�-�KYI����\�M����exَ����hr'���k�䓅2D߆�Q��I��eP�*S�+2s"y�7S�d�`�欱��{)�=�W�W�ƥ���o��)-�{���]�$J��Ғ��Z��j����{8Yo�"�1��w�Xx�K�i2]���=�G":��85�^�D��WO=T����nW����]8�59�jDjt��L7�Uu��g��(sS�����̸��� �=$���ڒ�zn�#���=�D�;	��9��%�9����:��+%J��[���J��V�9���9y���{��E�Q}�_v�4�U�*ܕ[-�æ��U�ʧr����}:�WVWvʬ�$���Or{�xdr_�$�7'�og����<�����T�曏%��Hu�����c:{�WnN�$8K��=��:̔��T�s%Q�$���n��)���;�^C��T;
9�&�[
D�$�y1&���^����I�<��h��<Y��Ǆ���d��8N��&	+�_Ie�V��D��I��I|<;)�7f�&�&a����=��9��H�!8��O&䎖5�	�L���:r���&�����q��=*Iöl��&�Sr	znN���10�2Iz�$�<G�	�I䇙'��ݲ^���;��d�y�:f�2�{&�d�����NĉC]'
2�Moa�-N����C���
Hm�boi�G���&�RxJG^#��1!�Du�J����'����u�̑3JO	�$t�0u�����L״�a<{�bl�#�'�u!�H��t�D�3�:��8N6�4��DL����(NbL:cd�FY(u����DHy�(杓IH��"l{	��'Nvɤd"%������$�,J�DJO,��aĈ����t��D�%	���Д"Fɤ��%m"l����DNbL:S	�'M"]$D�R"LI�넭��:m�4��p�[�"WR"R��������N��zK�"{i�I����҇H�#�u�i2$ᱸL0��"'�]8P��'�����d=��&��Ȋx��,��N�<k���׵��Y�_R$0�&����(K��%%Y���"'m"b`�M���x��a�	�'��!G�H���Ȏz�w"tN�K��:v�G�=B:ó�:;���p��OrY]��nP�;Q8;��F50�r���h9�۩F�gu���"s�27����Џ%	݈�������a�~���k��f�u�՜��ԣ�䇽�����WQº:�BY,�Q�D{ʘ9��/�xN�3g�&�<�yR��$���{���-O5[������)��ݲ6���N�Y\�6w�O��u�d��*oI�ߪ#Ʀ��H2p���������&ǻ��9'N��Q7�H�D��æ�0G����٨<�A����	X;�M��f�����ʈ� ����wU�o����<A��"�p��DG�L��6��"m�&�d�Q�j"q�D�K�N��X���(gj`����~�#	0᱄��I����u;�G~��Zԡ;֧:ȝ!�Aʈ��Q�Ԣ�="$+q}R�g�`���({4�ʨ�=|����=�>����p{����{R��Z� ��tۺ���gj"w~��{jQM'Dn�'�J�Q��������l�6pܜ,F�9�<+Q=؝��|�{ea�t��:=��(�4�Qt!e���g%�
f�{Bx$�G��ЎK�fX��v�{XQGt�fΖ>�x���v��l���:l{ ����u�r50��	�56L�V��dؐ���{�:�G&l��Cz:vHMX2i�H94��
f�ܺ6;���ggG=R�^,���:tn#s�c��Ĥö�黉�;�ƧD�8^�l�I�P{4�iQ��A�M\ٲ����ǓOf�����>�'VN,�d>���k�������<�Z��M��7���G�Q�>ʏ��a:w���0�.G[��8=�G�����:m�Jɿ̩VH��L��_���eG��jmʪ���jY�̍G�LuMy��T�J������&��W|p���1����Һ���v]�;S�9S��������س3�'�;��tp�&ǳ=;=�y3|�y��"]�e���u�^��ć};&�'��;���Q���'i��T��ԇ$�Ծ��*��=<>���)�J�;%�sfrC܉�]Ho��jA��;S���'$�ja�<oҽ694��I�ԭ�˩Z��H<�yG�(��r"<���*'7:z�<��a�}�]ͮD�$H�UIj5��}wR���c���eF��vD�ND�ܑ̒�f��D���΢pw�ZG"Q�Q0j'`��+I�"o����"'�P��X��R'F�"�WM�q>�����G�J�D��GNJ�y���r�1�Xlw���R�6ܮ�����������_�G�8O�T?��j������ο;?O�R��)cϔ�$���a��V}�
����79����2���v�bqOJV�cƁ����{ؓ:�C�z�֚kz�aZ}�uU�s���g��kR��>�����{�-k~D�����[��h�V}_���!_RI$Q�i��u$�{�'�	Ɨ��O��5��!#����>Z������W��,eA�SJO7*򏲛�OS[؈�߽,�<*I{g�>�"ݜ�\�^�ִ�k�/m�~x�]ض������.����΍Y�g_�z�|��4���eI2�iϑp��ʭ���g���3޶�Ӈ����M�:y4B�"(W䗆�ݍRW��L����KGVcQ$���."k+Ʈ߷鳉N&�F,���Nooy��;�|�bՌo`�;;�jRvcFFѷjP���x����mW�VBW��y�4�y�����db��9�\>~�w��f��>י�+���]�X4���ġ��mĉ�U%��ܽ�W�ǃ����jP�W�5�\�Wrr)��)�.��ڒj��T7�L8^?����֪� ��4��z���r1�8�6ڴ֕+_����Z�]M����ȍ�Xg��kɩg$�X�3���MĒI%��9��`u���J�r�.Gz��5]�+�e�M�v�J%���E�ԫ�����q�]I$��ӭ�Yń5����ji$r3��a�j\MD�H�3�����I*��v�ܫ��4�u8�#&��"��9�߹�^Ԫc�7_�9�ux�)�Υ�ϐ}�U��^�U4�4O<*I$�ߗ�{�8��g*|�]Ջ��5g�!jԗ{"+�>���Xj}�����M,H�$�]���s��k8��Z�6D���b�5$�SIC�$�,H7�2�{N�$��f�y%�b�>9�E�����\x��"����wj�+x�	$��MW��ĳ�Q$�R]Ӝ���61T^�$�I$���ʍ���ٞw�$��$8ַ4xkr�n�$���Ez�r9ͦWe������nI����<x{�{FpB�f�>W2,�����5��6oWr�j����WoZŶ�bZ��>�È����N��
��,b�<��D�2�8������7Lߙ�qqg(������c8��q�C�2�͕!��ʲy��ᮙ<�X1Dd+X�J��m�j��0���%Q ��n�P��&�ӡ�ː��0�K�e2B�l=a���N�	����W�A���Vyg��x���{A��`ă��Rә�}���!�zbX��<l��b��x�ay&!jĵ(eHg�]��X�cU���3i��K�o$*m�RM��:��xH���WK^s�p�,����K��s��bYu���Ã�=�񹵎��x����7`��p�d������-l�gQ�V&0���TY���՜ф�S�!��ר�]c��?R�}ϺG�#y�W�Teg��̺9��M+�wyKŉf_l8��5g<ﳻ
�ޡ�2S������}�h4���^���ĳDbU`��Q�̚����?,.�<��Q;p���	�%�i��Q�n�#���v��+�H�eo6���̋�,H�d������<"y��$Gy�$n���8=W�	��cC�'^|��.ҶF�����F�q�x,4G�xFW ׂz{��z6�C��y��%��s�q���*ı#��İՑ*9~��[�>]Y�O,O���UX�IcVڱ���C��?.��z�,I,X|.�P�9s`ɹ��H�$;{rQ��ŉj8(����,J,k�M-#Ib^E����ī��a�oua�Ս��&�z�V�8��7n.O�*P}\F�W^ʯwݸMK���\߹Y:meM���<H����6{�-ꘒCs�6�!�v}'�Zs�#���$eK���%Ŝ��G;9���"���$Y�>߮%=�������ȢĪ�f̉�>X�`�_��st�j��L����V���w�g��� ��={x������V�|��Q���9wY�D���,�5�lϒD��{�-��p\Ja����g�����%
�G#�޵�z�N�i۹�t����|S�F�2rY���*�?7�v����"H;�%A�TH�9��F�v܊t�'�lQ{�{�(�וz'�I��|Q�>+IbK�i,�|<�F��/���|IdMbIbIg�,��F�%ō$�8�*�cSLz�ϓe��O�G�q%�,GZ���jƪ�O��Ibŉ%�.>��ҷ
6������>Ù�Î�	>/��>zcIg���X�������j�U��sǞ���j�U���wt��Q�KKK5D>�c�ӫ�ά�~�Ϲ�8�P�����bF�Β�ՃX���,�����
��Y�VDf�&rdѴ6���5bD׃Yld��ܫ�%\#��E��*Hi��#####zt�#"H�D�q��bYՏG�8���6<����X���Rı,H����ϖE�:,՜�E�Do?h��,�sG�^o���j5g�����h��Ė/���:�ת�E�0rU����!6��+���g4�*��#�kpxqS��!pz�W��i�r#��>�>X�Ś�^(8�4|��b�k��A�:��i�+x����NۃG:���=�͕a�5!=Oq&�F�����R��Ú�#p�ԁk^.ZjoMM�*B�� �ײ�м������8Ԇ֤-��6��[�\嘑��B��x�#[İK=珬��z?|/LՊ��H��X(=EUg|�A4+�=�c��#EX�%�kʱd�NbC��5gxp�g�?,�y�V>�F��W
�Z�s��%��������O����8��a���|f�!�P� �"��8��:���.p��5ҖA�g����ǭ�,Li�w�-��a�Fo(�iYl�����j�Q�1�*��,M
��J�v�Z4���8���1�V����n�M�ȳOʅ���_#�ge����Y�E�	�K5�.���h�^Y:���ߡ���o&{X�,Q	���1A�,c�9�'���N(?<"8���Mo�v�B�<H�<n�D|K�Z�!7�g�B�f�<k2"�u��oGϸO�u�X���+���׉f�7�gw;21�Ѿ}7{1�n{��Are��\�&��f��HQ�<lI��ٜX���w�������'�y��
LH/)��ȷ�U�D�פ����G9�d.��yYRK})����8�ܼ�<�;'U�Y���o���|����19Z�{�n�NԳ��������$����X?�$�?A�~~��!��П��j�+�=h�THr2�k$���ӘL���o�9������RQ�Ŕ�)v#�����:���s�5�N&�˓����eY�`���:�;��K�$�㋍����,��Hh�;�]��P}WΓ�}w��w����%�R�z}�� ꛾��Y��%���]��m�-�#���pHbL��%�"��F$���+���Hi��~M`т�
oh���-�k�/�ȁ.��ۜ{��_]�Mj�1��}��mK�:�0�";3�LmqH!�&��i\��)z�JĐ���Y��r1��b���yM�<���~�M%��f��7�;��t�dQn��N2%X}N�Ⱦ��7�w��j']�'G�[ ��e�r�;����uA�ם�A�
�K�o\G:��r?{A(#�؈�蒉�]��-�}w�>Q-��K����ïjO�㾯V��2*�;����Moe5�s^�[�s��A�yf�-y;a�0\��>�N]o��z6�eG�����IӀ�:쯨91����g�$��A��,��;��vh��ܑ��U��N�'Gj$�S���n��6V<8�Ewc��DT�S�@E��Ek"����V$Զ+Y�'�%��j���х?��:8��*��M�uG(���\�^C
���K8�NL�J=5�Y�ى�H) �hB�m�J���M4E�X��F�K���5)��[I!�����Qeq�ȝi$4��-�����VE�5$D��@n�(�^���ԤI�S�K0��%˱l�Fk�EYq$�ԅ�=RkM�V|��X`�$��"�K�-JI%Y%�Xc�FB�1%|������҃���Od�њ(��bw.V�ǅ@4�P��H��fI��"5�gfĚ���6^�bė
�Ϊ�(��ТFjM�6~�J1��{�,"�FT4��������/n�I6����	~�r14����(����s���-��GȌJ6�Dգ��Y�@�.���-�t�M5|��=Qd@�&j)Fn�VQ	O1�q��W�R(��ל�\��݄#�=�!���RB0�ۊ�[��s��׎gR�K0���,��c1�F`$đZ�����L6���މ>�"T�B�n�4��r��5#*m��%<Uwӊ�KN[�$ED�%l�jb-@��qKGJB�","bh$i\�-�nȅ�;�d�Ҹ��5�Q:�\|��ݸ�mN4�WnE��'�뺴��y.n���r�UX�N�462K"M�������4�$L�j(�`���x�q}P�T���Q��.���{�3��O�z.g9�$U��P!'���d7��a���1��̼{F`q�fM�{��2�Y31��|nԵ�gLq$�$9'�e�Gx�{
E1
pgXR^��Y�1y"��#D�P�r<�2>7v!��j	��*�,��(��3���#�:� ���Y9�cX�ڞ%f���Lq���3.�����\�Ln�E$�	�g�t����\������U \=���&�QSX����H�b��"<��7@5�C5Hc���j��W��=1sU��cG�yDuj7ϋ��x̪u�Ñ.<�.!ؕ@�d1�FٌNj�����c��5����'{�I����A� k�Cg�_���O����������G��AjQ$R0�_��~���������+��{�����UU�*�����U�]��U[Ux�ګ�V�^*���Wj�Պ���*��"���U\b����U|���U�V�^+J��U|���U�]���UUq���]����Wj��UUq���[X��l��Bx�,�����؋Km���Eƕ��Y����I�+K�u�ۓEm���r6reTAF��U�H�ִE^s�QUUQUUQUU�*��iU^�7J��v��Uڪ�Wj��ZU^*ڮ�W��U^�J��UUV�S���*���Uz��v��X������V�^+J��U\Z���v��U�iU_"��Wj�R��F�e�ڶV��I�*�V�))f�2L+e6ifVR�Y����5k[+1YZ��&<Y�l���(Q����&jd��ɢM Hh!5&����ʻU^��Uz�UWUUQUU�*��*��4���UUTUU�Ҫ�V�U�UmU��W�Ҫ�V�U��U\H���iUx�jҪ�X�����Uګj��U|������Z����*��V��^x��Vڶ<L�,S)���P�n^��e�lH���?J�	(�/ޯw;����x�j��[UmU⴪��*���U\X���Uqb��,UU���q���1Ux�j��[U^*ڪ�V�v��V�U�*��i�W�V�v��X���U^��V�^*�Uz�UWU^��]��v��W{��9`�;*�� D��h� .�l�a�Յ�x��oI��VV��.pj̭��՛r1�59m�&ۑ�rX+aɱ����ܛrڳ���@��!��Q�E$��ȃ"�
��cQ����??�?�@T �������ƿ��)��i��������.�CN�K�<��:�<�H�AAD��P�BX�:tN�d�DDN���8AD�8"xD�	�t��: �� �$8&����b'N��<'�0L<"`�&	�0DD��D����M�"Y��H"l�lN�8`��D����bl�GA"'D��� ��"'A0Ad�ı,Bı,�Ģ�4�xA�AM��8$:X��ǋ8pDD��0������� �=� �/���F�+P�$R����+l��]���A,��e�VA�b�elcj8 �Iaږ�2XGPB��e��5&ŊI���V4�iD�+i����A,T�?M�Qh��k�H"EQ#�!���"[m���H�N�9�`��QQI)�L��A��u:�-��MD��-�����jLH��E��"-yi+�y.JҌ �!H<�-qfAV��J��㰢�&���"nd$�"Lbj�a��9R�([�U�7���R��[PB�9QX�+`Q(�Ԏ�I%"�,�#����J��2	�N�QTʨ�%#I�:؛Hf�<:�����BQ$�NX�V�u!e�T��M

�cR�R��;Ѵ�e� B&ZZ\q2��
���x�Ŋ�Y)�,%A'��5r���)n9��SI��Ŗ��8�Ɣe�cSI5����VE	�QT�%��-{�b{/�q�$��OK��Qr�T�yX�,R�c$�XӱKr�%�-*�BRdJ�d�ح&Ir�P��H�!��Z��![S��P��lDs���#F7�Dr��hX��bV��n�M*+-Un<�)A�%i��r*!A9��b�~[����R��S�X�[h�c�*,lpr�l��nB�9�HA�PJ��k�G�(�!��!�H�-1� �8�D+���Fl:���KG
AhPw!K䨍"�R̢�Z��M�Ց�
�Yk��!1�Q܄����7FQ�YXX��K�8'qR�D�1��V���	�n-BUYX����ث���A��F(��S)Lʱil���`ֵ���RƲA�Li�����ʱCp�,���Fʅ���FT8��!A䅅jVՌdkA�]nJ�1*�#Q[��y�c���ʕMD��am�Н�7Ia
9��;J+$�
�I�풃�͂X�yVQb� �u��")2��i�X�Zٰ��*��
���&4LN� c��Qx�U���FJȆB�i���p�)b���2i�1�|W4HQ(���[pTH�pp���X�h�&���JM��Q	��l��XkȍNV��1���2`�bC!�H��%b	��pD$U\M�jTBY�*�^U��2�G����)�(�M(�nK��bt�d!8�l���B8��
B3��#lpب��nQc
��LdE��p-��,Ucl�,���&12�ImNc(��+J��"�bć�	��,�Q�A"��+$HD�HaIԸՀ��D6"��%I�'	+������e+�!�)kRdR�2�F���A��M��)AQ�D&��E�2�F\X4YW!K�hC��;
�ܱB��&,$����T��B� �2��Ki��b���Q�AF$Q��J4�HpUIr�Q$��������I$H�1>J�N��ȅ�pnGRPx��KP��pj�nȮH�܎IJ!��kDU<��IT�,��
Т��H��w�ʓ�����Ke�㊶��V
��cx�j�M&�����O+�r���piF�(�����V㸩�J�m��"��+H4������cյ��-!Tn�&���bvq�h�m7
F�:܍L��$eCE�R�#����$XFؒ8��%�f8�KF��X(�I6
�1�]�[��:��R�6��!5KJ�T��*���Px�m"��1�M�Wc��2�n�dn����\U*�ēM�
�ĝ��@�VX�RW[HM����(�t�eP�H�KU)+M�D5Sv�<�XҖ"�*���BN6��M;g����$��Y�bJ1���I72±5b��[M�� r�bITBA��:�H�jW*��u:���BI�*Dn�5k#L���m�rԲԄ�Z�J<���ۍ�I�LL�ȇR���q��%*�j�#��H��52v+*Q��ۖ�DX��
Gd�GlN����B' ��F�4�X��M��F��j*+"*��X�+Pʊ�BC��n�j��v�q�P�ĕ�Z&X��r����q�ݑJ�Ķ�U^D��5d��n8��;�oH���e%R�6�*$�H���`�7Q��:�*�5�m����D&�,�cr!�T�&������o��n����6�x�X�-��Chr�z$��������秿}���(���[�֎s����ϔUUq����4k\�9�+���(���[�F�A�s�,\���UU�*��tT��:(�t���	�0K0J<&j�ލ���$�[H�}6��NS�c�B����6]+����c���fA�#�XUjU�+EU8�E6A��hR��H����)��%h�(�M,O-%V8�;P�b���hB�^�ˋsPF�K*�*C ;UD�%��U�n�!�УR�Hpc!�0�"`˗"��b�M�D��P�Ĳ8DW����
� ���A�+J�he
XH�P�B�9�e��,��X�Z1:LiB(7(�8�8%GJ<��Y���"e�6[$i�q*�vKQ$[7ukU��Y-��Tt�TA��U�6�v��bd�$� ��)j�Q��1�Bj�e�F��#nF�&K�c�"I$�%9YVbq�UɱT�Ia1��Y�J[kN�jQ��9*7uL�ŊA�2	�SmQ�#mB8�jZ"�I$��Be��JZ�R5,���*B6��B�D��$� �`��J�rAQllB�i�$����Z\�l�O�~)��0�
�h7W_�Ћ�念r����{�a#M��I��ٓ<:X|4=�P�E�<���$���:�e�M����[�&G~v(�a!
h�#��h��MFr#���Fh�e�M~��Ɉ�S��>����]�g�6p,�Y���"'DD�,�(�;�r��o{������$�H^��1��{�N��480dy�a9��&�|�:d��x�:>����B�x�r��U�"��gD	{8xY���O��^6h15-�o:����hTD6R\f�*s_kG\jOt����j��̗���q����:�l�c��k�T�Hrtx6`�g�!e�gK0�N���Y�'O&؏`ՖK�M�IJJ�L�_L��f��`�J+nZ:W["��$�lN�+C[*�[�Z(1D4�iC[g��N
�I\�F˯��ռӥ{��G����mN���}���GD.|f��=���h�Ӕ�#:gr
����룃,<���ѱ��ڑ�PwN��	��Q4�F|=1�p�P�K6t���|tDL��	��#؈��$�F��K�$��{:p�xf��y�X/���b��~a��KQ�M~���n�_KH&G��ۼ���X:=���C�	�)�q�{U�乡l�JC�!˦i�y��j�����í���s�F�����N���t�����3N�2Id���a��L �6p,�Y��Ζ'��DD�,�(�V5P�7�ns͐�<F�#KzN�%:���Lf�n��;�S8� ��"5dZ�)6(��;I$�����C���r�[-M�2�!K[�u:6�-tE(�)�iIG5A6&:�Q̒
���[�8IRdĵlYu![,���6�+4�yj�EccW��ǥտ�$gK�#�$��){��H��q3:f�B����tvv:|:6OsTBUQ[zN�u�@�ä1�x�.oV?Nc�$�9�zxm<�������.[,��!�G?bD�룄"���NO�\9��q��\+�w��fKvL�����g2K�.Z}��bi�e�v	@˔��"�X��1��>W׃?V�����[�S�6ete�a�H��0L��0�}�{/r�����m�~��<����6Y�n�ٷ{G[��|�׵w�+�5^�$�G�4�d3L���˷�[�M���.��f�;wiW5�E3�©!	<�~��6�2B�X�6q���2�%���;֞�z8x<;��8&	eL^$��b�i�zn:)5��N����2<I̰q�t�;6�[a>6{g����̙,�`�2�
a�T��y�yכ8�����$��K��I$�8ge��68i���Y�����8J׶{S�&Wɰ�AA6CX��Xgw�ުK���fsO�k��s{�������㷽\���}�= ��
b!��Ι��0pϤ���n�F�yd!C�����wX�9���ٳ��=N$Rp�^WL���=��Ft�YRp��&��܃3O
�ӇƐ�F"�����N���`�	��rksp�I$H�Q�TI	�<C��Z{
Ӹ;�u�w���m�)T�N��&x�Ɩʑ�µ��Z=��p��?���ոh�ZX�v5�BI6|�e��N��h�2vP6�k����i7Rl�Q��M48�CO1}/���ҹ�C2T�c[M����8 uƸH\x􆜍r����0�+�,��e�)��y׏�4�㉧�Jʼ���DP[A!2{�5r$<|ע�Q�v�#6�)rH��vc���*��E�ɩRZ�jeh�'k������I$X��T쉼�tTE� ������DRR\De��J�i	T�6A�0N�l���j�j-�(����D�"HF�&X�x���ܜ�\6K��!�EӇ1+9 �6I�V��q����e�g�t�m�ę������a�������B:7�!+��K����w���ܓG��&�SE�r"����E��T�����FƇ�U^��H�c~=z�;*���θ�,���	V�=�1o�>��dhkDJ����4������.<��)O~�c��bB�s㆝!��JC����:߷;�{,��$��r:
w�v�ѓ%�xS���]��6��;���ϓf��̘:L�D�OrwÑ�z#=�x�ǀ��O����t��E6%��x�4��Ô�z��vh���g��뤒{;��Æ~>Խ�$A*�Cr5�m��8L�������OPn��zW�s����d����x;=��W���IO.�o&Իh�bJ^0��;xs��Rݩ;'j[���=��B0��.��0��]�>mw��4�:�o>ěE��7��L/IIJ�☤����������>O�_�ן/�/I�^JO%"�]N�M�}��i�)tf��Iy"Z�"�ڗ�RZ)-H�i�E&P�
aH�R2��F�/jN%#�H�R<�y{�<��Iu<���O.��R<��<���N)�4���R밽)~6�%%%'��]t�R��0���E6�%I��)yu"��^ԛ��e):�M&d��&d���$���%8���O�׺Q))K�)))��)W�a�J�y|I;R_�tvN�d���N��dn���:["N�w\K�Wn$�K�v��J�c ���	'D�t�:L%t؝Ke�4ʑ��u7'[b���_i��W������i�s���Txw(�3Y۾�q���9w�'dU��5���}��+��w�!��^�t<��wN\.���m��V�q'W~��h�;^�_��{�C������{����H|�����I�jE|�4���X�E?����a�ܜ�~�O/p�9�u�;����2ѯ��Y��ᙙ��b*���]�kF�s��ɕ����رUWW�w��L������ʪ�*��֮�������}�}���U�U��\:Q������q�R���<��yNS֩������T*��\n�H�Q֙�p���	�`�P ��uJ׹�n���'���C� � ��:O���g'9(2��0CPX��O���$GhNKZR%��3m/�����s���yM�Ͱ����}����55X�d�`�0�d4B�Xl��]:h}���$��@h�LFC.38d:���h~%�� �5�UU�a�Q��L#�4; �ʹr�G�l���h;��IV04A
!���Ygȶ��T��4e�i�a�]R�u�qלE)��_�c���j�a����QQPH
�cC�L8|�`(�	��6�u	$)�C�����	������4��
>���qp�W4�M�E�a�wM�䵉g��
hx�zi���I�M'�tY� �P0F��%DD�Do
��C@p���7�ۻ�-��B�u-s�0��A>`�y�兄1�s�o��l��\=����x����
4&�p`�Ot�u�}�HDF^����H�-
B��o��,264��a��:�:`�gii�q�_)��yםy�������t�ߞSק4�
����^�:�'���;nq�N���\��J��N�UEES-</���+7L�%��PasifA�	�q�
Qe��s%�e��KLM�!,a$Ȅ��!�D�m7�	$�X��Qd��ܪ;[t��1o?��ErFR�8����Y&uf�=KD�J>Se�ߤ%�V@�HRC�'՞�#*��lwA���f��rCc�U�p�"��Y��ξBE�ݴtn�:0�$�}*�a�(�F�%��9�����hkD��A�=��?
���}t֧y8�>���xC5%)���(����i�[g�>*I!C�m#ޠ��'��P�:E�Sc ��ّ|!���~Jm��)�O�����GK]s6�We�x��b���<0����D����! h|PS�	,eN���mL4����4Ì8��)��&	�t���0�&o��/��=ER**	
0�'*�aP	G��q,DXҤ�S�=��bC��X��X6C�Z8����!0�Z�E�!ȳ�+�_��;�
�IG��u�d,R V��>�hI_T+i�	)��핹Q!U�t����� �G���LxQa�-�Fo��.	�IH�0�;���ʕŏ�$�U�s��̜ٜ*Pmx�P�S��ܸ��}Ҫ^���Tv����hV�����a��&
��W��CC�N���! �r4V
2)}h�4�Qey1�[��؍-s�ˌ��2�4�0��J|������8C��ߖE'��X���ADw	�ZA�P>!ΔP��܎�DX��/������5��)p<0��U|��۲�}(�H�B%YP���|��n���YV�Ba�{���b@|tetcռ1�F3�q�$�cmµ��A����eu����L�P�8�mo�+��]6C�Gŏ"Yɟ����a�����hpB1C�&L�H[�0~�00C��t��-�i����z���8$�R�� pa����2Q��_����ϘZ���4���F���m�`��<A0�-�_{��z���uܸI��U�ݯ��o/���n��p�"���lﻕvG�N\:��ĩ�(��xM��***RC W�����`�⍑tC(pB�Hm!ht`pxQA���a��hH=!�w�E�
wA�:�9�3+C����a/�F����|��q����v0�A>��ΊD7�%!���nJ���><�� �D&�C�������P�Æ���!�G��h׷��F1��$6E熎�>&�gx�����Ipq"�hh�e�#��
4�i�0zC��=@၁�AqL�����6�� ��
`ტHEIt	�J�`�0��anii��|�����yמx��9�������>L㋘������d�4�b�m\\M�ۻ�O��&A��Dqb5i�ԕ�W�F��'k"�E$�J���^���֊����דz"Խ��
�H�ib��JLBNd-C����!� c#WX�#b-A0��+V$)�"*�i���)�9^EvD�Z��m�RJ�1N�����?�Μ��7�:k)�k�;�;�b=�Cޥ�����'�-���@�!��$��I��da��d��@~xYg�A��P�~(x��&3���!��ϩ0�g��P	�,���8�|Z9�8hs�EUι0X�C��һ)�:a�(e�(!Ph���6@�d�NU�)���Ϲ�a��2_u��I%1�����ߧ��7�i�c��x�3�w��ܿe���Z���w������Y�T� q��dσ�����R��� �b�2�k׫8f��Ӫ�n�xo���ѓ&������x_a���a��E�Z)�9�ZE֢"�!�Lx��N�!��i������舘"'OL�d������c�0��9��!�"���$
��|�t�5�c��'�{�v���ǬvC$�	
��|86K)��	U��d���t���w��0)�W���	�#\*��!N��I��zh�t;d`@68;�^G�΁�0np�>X	Dx@Df�{�VjrN�!����lM@��Z��^��+fw!i�!��y�x?i��ń:641 �s	�hbc�g�åA��]P`�Εm~r�rӭ|d�c�`��,�g���舘"'OL2^�_���V|L5g6������MU�OC�B98��0�nJ����m�aF�02?Q�0B�1p���	�d����4X�J��_�=�kc�����н�8!-3<틊��%��۱�N�%?����n��$7�f����9��y�C��gx|b�!�l�Q�Qf�|S�!�a#�0i�c�H4�`le?ke��o�������CN�$��M������5}�e����zY��Z2U���d���a�ò�6h�і���q�<��ͼ�μ��8�?Q���;1��g�w^zO��Kp���f�QQR�{�a^�{��S�8CͪI�Vժ�]�C��9�'e�8'��j�e�)M"j�� �e<q���>��i�	!�b��L�� �C���FI�.G,"�q�H�b��:S8!��;Bu(g�s�ÆF�z�H�6Ry�]�rwp黺�ѱ�5a��I�ۇ#:2�_y���6���cx�e=�d;���{�*��i-�k���ߝgI^��q?�mK�%=y�JJyu8�j_h�0���;�v�^j�I�;R�Kz���	�'\���7��'��	��X|&���"u�цǦ/)u*�W���ĺ��K�SԔ�&Խ%=y)<������w/�SK�>H�%����I�-DRD����R[	�Re>i�O�e�������7�^�'��/n���ꗵ<��]I�Rm)�ԞJO)u'����/�/���eLR4������Jq{�"��H�����q)8���'���ڗ�&��%/m%<��II�u��H��4���◤��)��JR��R���JR��JL��uKۇG�c�bh�L'Ig�N�������b��%$��D�D�RDu"*L�E��L.��)2���&�H�iN���_�^q}��%#�j���}���q;��Y�wyl�^I�����O���N��gH�n���h��l���vw��VU����p��Y�.N�JI��M�v�ʼ����y���Z��������K��~�uNJEզ��P�r��Q�\�{�&���8s����a�ا	���ߟ���7
��f�׾}��9���j.�ǚX�UK��,��;Ǌ�}#������oM��yᜥ�CY�c�[��]�{ƋNoծjD������L_2	��O�H=�R�0c"��v鬚x���G_���}�W�({کo�S����V����x��֚��=���o�PE�ǵ��3����odwnF�/0��yi�g�ҬM��f�9M��4�R$��nX���
&��u�[S���E*u&��BZ��u>X�!j`޽�F4�vZۭ�R�Q�|��5+��s�-TpR����\���K�j����y��n�tT������s3>g�J���{�{��(�sY�{~���W=Uz����������y�Y����V�����>>�w���Y�{�w��V��_��UUv�UX�,�k���p�H�L8ÊiJm�u�q��蘃��Q����d�2������BFXV��*��a-���ʉl�*< �hp�Dm�A�m �*��Kh�ȝ��*E�R(E2�I5���T1!d���D�EDȉ���:WX�#)v�V|o3^�	�,�V���(�;J]mb{`�`�B�*pPW$�Yf*U-x�*�rMB��rܦ�h����#jA���a*�@�62`�V5�m�aG*)U&2��H1上T�LM�R�!c�d Ĭ6"�����!K�m�Vd��YY^ю��v�bm�T���RS��Q�diI*�)UQ�+���Kj�.A*\BcpnѢ�ŉJ�ycj$尊F���cJإ�4���D'�ѥ`�d@�HNUR��E%���+�;�$�qT7&F�e��\i�`��]�+*���e��ٮ�Ay��Lc
Hc2E��J��^D��D���+n�b)��dxD��:3 �)k��d��;U�X�M
Ւ�IS��2��ҵ�T�	�$�
*�:�����zo��BV��U�+�)}�x~!!߷$����̣�``tc��$���h�z5�&�D0@::9���x�h~8`zC|d�ˇa`Y��r_�Z.m��>:�lzB��W�5��l����&��?:C�.����#��\��:!dXdg���$�^�L��\��Dy�)O�-l4����ӿD~��I�e��w�8��.x˰�5Y_{��@k����'��#�n�aNY�Fm���h����4��|Ҕ��<��<�#��}�V�5�ߛ�qٵ�6cχ7�=��1�c
H=;�+<���at�RW�,���L�6h��N��Y��;s���lrߌ.Gl�@ƽ�a������}�MV����� e�Lm�ۓ<��rO�l�|A�~��C1����nCf�0�H6B�}��B�9_΅'����m}=7o
r�2�����n�*:g�4ώ��;>�/��,��'�nL1�$+N�-��� �{V-{�Z�<Ռ��}�W�dc�*��YΏ�b�|q_+[aO8�ii��S�>|tDLǄ�k���V�ꮨ���eJ�*T�4C�>ld4����r6B���O�9�%:��z�zB�ς�\�2�}�O���$c�����m��o�;ﳋk'�u�T���kRX�C�������,�?m�!��w�}�}�{Ϭ�_��b|I�љ�?i?�;�� �G�O��|�"���������
=Pv;-&À�D�Cd ��OBj�piNW��r_ƅ�ŘF�[�'Y���|���O9��n�m��6��e�i�a�<�����"x���Բ��U�]���&}&��1�$���a^�HBp|>�����4�a
2_����3���^B�ꫨ���ѹ��5��\<i`�7m&9r�6z�!oG����Ω���[�{8<|a�4I�Q>����h6��GƆ;t;!�*�Zl��p�S!��<��c��C�0r�q礫��&�d7ᠨ�i�����|B��A�]��o�-�c>{�M�|�9�?�6@�Y>>�Bh�2��ǚu]��i�0��>|��D��!���=_g*�EUl����bPV��$,�)�Ĵ����b�]Y�!�&!�ǫ�i̭5$$Qڬ����X�vF���M4�M4'��	�Z�5,��s%��r�Ob���&��"%U&[F2�����#�
��[1�IB��q�m�J4�� �D���rJ�u�aX�[J(�Ek��Y�����~��V����M�����w����gx��GB|�!2��u����SEЄ$9{��8Rzp�>�����l�jl�Y�-�m��h0É٬�28>g� ��A��d�֫�l:zh0��!�W�gn�n��# �m�8B���p49v�H��2�kҽv�C�Ԝ�R^��7��t�ĔxL	��tE���J9�rmH�������"�Db9-r�u,H�S羨��џ�� x�!f�� Rt�_�<�2|tǧQB�њi�X|��ϛS�:��8���3��3�����:��ҳ��ž�i�}]�o��L�-�����8��ù����f�oV��z^/N�z#w�z�{�9�o]w+~*���y�{��ޛ��c��oC�j�&��E���{=o6}v.E��S��AS������M���Trzw��}���]v|ŤٿN^o��r����~J���K�Q�5�_d�c�0��_!7d F��r8�� �ϰ(s�!�H��2��`x6.�����Q$�e���ep��@�#�}N�WK��(.�C��K0}Y6`0t�g���oUw���AqL�7�,���?��m�����~�w������7׾����7랮�﷛o�[ߛ ���)�m9u龜	�a�[4�;��(#	��cPM��l�S�/������lk$�,�.�I",�5ں��_����+L�y�M�����m��a�e�XlD���t�D�<xHa�Z��d��7w;2k+�9�1� yt����E�;$���@%JD���Ą�Y����r-h<[z�*y�]���-�\���g�)�X�*=�����H8�@lɎ�iZXIj�IY�.�9������l�4O��9�R!��K�ﲟ�����M�s)!�$04��"#����_I<29�����2�`!%t��'>�BB�6S�u��g�=uM�>Vp��}"I�����u��f�H�ht8ݴsce��c �*�D�M����L�Q��q�<ҟ6��u�qǑ�c�<�M	~����&}�c�1�$�qnڙu"��e�m)k�#ꚙ1���L�bق�2Hǎ�&~�ɩ�+\�Y�3�c�[HAIHU%$ �3���b4<g�$/J��pD9VU�/�������(k�C��(����l�d�����[Ҵ�j����Dv��;3������$s�8m�KG�;l\]}F�/k��:�8�x8,Z(�%����,r�r�,��[�<@0YA��a�7Y0�d٩!&�1$Ej�GN8���̦>k���0�m�q�X[�Fy�S�>mJx�<xHa�p�wW$&����!y&�ҠdK�.9�{�aB�)w��죽!���	Ӽ�>��;ǉ.�'ձ��(�m���Z���q_'�_��1�'���\�c��q4kHI���*�� ���zYH�"���&$<o1�� 䢤�"*:�Z�&�@��dB��I\�RJ7lb��v5�`�7ז�y�
���i��$�h�5_[��m�3��(�e92`|5Jd�^�c���}��>5f�zH�N�%5��8r�4R r��]U�)���a�J�«�Nj�CI�L�uל�aj���-w���䝾mDp۰˃Î�}$�e����q�ow���e�'�6?��a��:hъ�<+C�ᢲ���x|l~H[,���ŏ�e\(�Oj��_}Y�q��1�qO�jϼA����G��	��)Yl*��nx�=�c�!��Ag�YbE�r2BLYq�C���gBE))��_>mJyמy�G\����&��}̵�Ϥ��1�`	P��׽�>+'��"U�~�1�����^�q�8Y���}��wf�i���	��͆|dW��E;��0ӿ���3;��L^����0���-ҙ���،�u��m��ɜGBP���O���B�V�}��ud���sQ�[�E"�N����GLG���g�Yr�fT3Fx���+��В�H|��`l�P���R��&3!�����S!��	�s;�>.3�Έ��sJxH��y�>b��������^O%"�]\���)�t��wZv]�'u�y^��v�ړ���K�����\O���L>��>D0�	����K�)��V%/Hҝb�M^SL])"��^aLRRm)))�ʼ�JJyuq.ڗmL%ZJ��(��G˾H��o�'��>E��ɔ|�����H�)���Iĵ'��.�)F��
eu<�Կ�Hʗ�)<��R��S�:�L�x����R���k�)>O����x�'�t|��_��RR:����f�yK�I�.RnJ]M.�R4��Jj�.��J����eK�RRS�b��M/��QK�RaK�So1H��RT�S���%.җ��N��Rcr6C��t����=�����N�	ғ޻r[�I�v�k�ۧ7i��i)6��4�R�ru�N��ۥ|O����o^}��o벥���Vw}�?y^���p����T��ֈpk�u��eq�dn=�o*����!���꼅ӽ�ȴ�oK��wF=���Eh��sC ����	wN`�B������4��Y������5O���/&��)�����5ީW[��I��qs��﷙���U�U�����߮�����fg�uZUW�|}��o�w��fo33ﺭ*��_���{����y���Uڪ�b�r�6k���Yg�<Y��JSjSμ��8�:��x����{����1�%�P�I,��k�#���Vq����Q��F�A >��Y��!���afޅ�e��O0`t?�	$��Ύ����}��p���gQ�S���YK]S����.Y�8p��nqM�U��w?`\`����l�0z�I�q���¸Wi0 �@�V%��d�n�&r�<p8sϚ�nh�Cß6T!a
 �{64�-�L6W�4����ho�U�&K�cev�<xY�E���͖;0C^e�]|��6�<��<�#��u9̷ȋWp�wV׶8֭>�r1�cR@�z�/[c����C�).`�HT6$��eXV���g���r$��/��h�ff�v$����S{1�i�s7�:Q	��p�9p92:�״8���ǥ���W�}ic[J�	![ l֑>`��"zM����/��m�情�[��Hc0�2����ד{�z��"'[H�clY葨��������9ho���] �-ɟ��2�����:�e��q�<��ͩO:��8��x��9_w{���G�,����O�|��!�)�6(-~���9+�U�u����a���.R�yJ���f����S��TV���m6Ye�A�-m�REl����x�p !&�J+ ���q�DH���B����rXB�ULvM�e�T�Y\*�uG!�K���B�$�!$��&�g�)�cX�5�Y�xx~���X��RFE�4}c_66��w�!x���O�Gnۚ������{���J��6�㮝��;*4��z��Y���`HB1�w&w�.N��R��!��͐���I�À�������=R��+��V�h�jC�<+�����h9\��E��fS;;��g>���Rٍ�IZ����~]6�?uӧH��/9�z�WF�����h��g�~��u�>68�t����~'ΕKd΄"Z}���pΟ̭��-��l�y�>qJS�<�ӧ�<{�ϑX�$�BcBX��T�i����R�jT�\9/Y�-u�ejڵ+�J��W���\���**+T�c]�f����d�3Α��e���o������:v6��u�Y��ypIg�B��ә�3���]:�}�������o�gX�7�-P��8�Nxӝ��[��89���~�n�!�?w���5�aԮ	�p*g'���L�r�D��C�n��8:2���(��ftFp���?9>��yM��E�R��|6?�H7)���Z��KLA�<G�p����4�8f;�Gc���M���(�%�E�i���&�C�0���t�3A���{�.�����u��a�e�a�)��8�)�<�<����%g1�a���ܨ��R{P����Z��s�<��Y	8���|�n�m�W��$!�1�>69z�I%΃m�'_x�{��ħ�A�}5ݟ{������Y�m^�?��[���zΣE�����`��/|韎�3�<)�i���B�����L>BY�f��4f����RN�7�/�,�9���6���8��"l||6:�����M��L7��`���L'�<?�C�ן��!���ςE<C�8yM��R�S�8����5�Û�uәwc��j�!�5�ϕ���x�.���t^�E��>�"���I��V�Q�/��0v@߾�`�i4_�p�����4�Ό�?w��U���ﭲM?i�xr���M�/f����Y����@Y�rÄ~����IT�g����l�'K~{$�N2U�Dg������/�d���y�	leK_Ky������&"�y�g�BV8G\X`��|]�p�!�,��<��y��e�\���X�'����(}��4�A�+�)��So�8�)�<�<����&F%��M���cM�<j'��2��䠅����O�K�W���B��+r%!kJ��_��**+T�7��JBNK��_�3P��Q�RZ"Xm7X� l(�P�Z!���R�G�&(X�J�P�=ĈU�mX�iQ"��u�H�Q�h���D%���Q�s/'�zY�����Ӝ�x�]�)q.� ����n�����Rf2�!O� |h��Y�@l20a�Ql|�a�Ã�	�C}��hrw�;���ƓQ�ay���m����20�D!��J�������o��xތ�<.c�{���ϳ���X������nm�OH�+�>+Ҿ=�P��1�.$-�VӲ�S�y��'���B�s��1˱��O}!!����$�p��:�G.�쩇�i�ͩN)JuO<�#�F7�Mslf�o�~�4��������%�%{\�Ok���%I�<;z6z��G�����C^{[;7��SURTё���3+���<4<����@������@���vC`��@�KK��/�0�trP�>3����1�f���<J!i��!���/M�ٷ�Ώ6�y�S���J�ҺW+��_sF��`�x;�99��#>:����0��uf�����@��<��T���M��u�2���:a�e�\a��ڟ8�)�<�<����ݰ���oD�?x����I��ݏH�B�Ma�F|:ofh|a�|J�8t4A�c�=4L;����c�:-���C�cֱ�����������RҮY��np�~��ё����:�f�VWJ��>��J�`�3ZC��ŏ��ٟ��<lh�S�J��~~�k��C��}�92o�t�Ґ��-�3�.��ij~�矍a�e�/�y�6��┧���8q�XƯ���i�F�+ꭕ�ewEeY\=���h���_W�^���i��s"�蚞UJ�#�5Y����v�h��Y!�����f=O�#�T<�)�Ǉ#���L[�08;�������7;��|�Đ'M�N>Ƀ��*Wձ�8rsD������#*ꗍ��*��d$���6=<:(7�Cm����6?8�|6t�(�'W|��:�O8�RyK�W��^������4�J"�j"�$RDS��ڞ�v��x[�I�t���a!�2�{e��'����L�����^�)}%1X��)))��W�]�/�^�V%/M/II��)R�U�WW$�����a(�"�t�Qړ�v��I�v��N=�e*M/l�]Im%%қ]H��R[�^�R�jy�>]����)x�%�Jyw��<�<�S��Q)K�b�RSk�җ�y8�H��]%&QII���S�0��a<��FT����eK���L���^�L%.�(�R�JJR�S�>'I�O��GD�����ty���yzKyM�N�䔾Ծ��M:��]f�	�Y:X�Kd�Bt��]�;v���q-��;^���)-�/����_�I�o:�S�����z8t~=�����w�z���ӭ�ȶU���aP�������{�1��\��m�wx���[,�����Ϻ^s���I��W�;���w_��W��<�4h�A䦎ҜV�V2�Cn:E�wK���~�g�ӧn��I8W�/�eh�aJ��8�V�T���/�[|x�M�^x\�I�����c���s��ZZ�V~��ť=oG˦�y%�Vls^"(���,.$��Ƞ>�s���w>}���rG�ך��5K�Q�m���?�Te��G�yz�O����;t�5[Uʓ#�X�VIiD+B-rb�5JF�����EQ�j-m4�v'R��%����Kv�hi�ɶ��:��7!u�Kqn�8�����Cc���e�Rli�#��F��T���+����j��^�o��󗙟��v��X�ܻ�������}�]��V+�%��y��y���Uڪ�b����y������UmU��o�Q�x6Y��ˌ8ڛR�R��y��|�NDFI�G�T�L���c�)jB�R��m��nW��r�$�f1TWGIFI����7�V���H��Ud���2+��a]w�*JD��H��SUI�*�+$�Y����k4ɐu%	,-hU�*��-��1�`�0Hc"�Ib��3� �ǎ�KmrK(��"��!��dҌ��qJ�Q��ر��B�-�!
Kk�j
V:�Kd��n��d��,��
2�tW(�m"f��C���-��,L���PS�B�Aa	��*�Њ<Ub+HV6�
�R��Hv�9Yj,CQK+eR�M$ێ!�Z�"�Z�X�(���D�r�Q1Gbi��&��YD2Զ�Uy�R9d��E-�D�;�4k�r�221����FЇ"n���h�*�c�i4�	j �NԲbV,rbV�$���+�ڤJ$�n�˙���**+T��4�d��ړ7\s�v�R¶؁H��YH�xR�dIeGm#cd$�a9#Y	���E�)�dE�27X�D.[qT-�V��3b�����#���F4�v�CY)��;³�qp����:p�EQs����B��C��vlp��vGl��e}��ѧy���^�C��?x�>���x�t|��e�C9,��'��v12&��3O��B�ϣB�=�����-2gM)��$�����B��쐓[:��C���s�T#[b������m���	��F�K������8����NL���8�����(��f./Hl�h,�e6�l>m�jS�R�S�8�c��Ly�=ݛ�͢���I
��p��Ϛ�p�IU���28�u�M�ig�D+�;'i��U�ɢI(�RU�NC���2?bX�v�0���BKl�),�����k�`��
U�Hl?nͮV9�z��iT��\�r$h����~��������K0g���1��<8h���o��yr@�$y�tC|�j���,��6��[�8p��2�쩗XSjm�R��y�[��c��m��	q�&B]_v���U-�I��ZqΖ�����I>��$>>����t��|�O�N3C��Γ��&�x{hgH����mʈ���2y��lR�Pb(���e����g1��}1�׿ƞ3�Q܁L�S�UW��>6�ǔ4xo㣔2������LZ�uj|�Z^���:��'�G�F9=�[���3l�[*G�:a�a�q�y�:t����Ӈ�=Z��'mEJ�*�h7o4N6�;Hp�O�g���Lfi����#��ۧ��8.pҜ ��
si!�DFճ�K�y9�t#	��ߊgt�˗S�և�NM]U�̑����m���#�����(u�����X|�K��Z:��BN��ƞg�����_N¥L�����)��	�ˀvs�C�G�EU|:�\::�tv�߻l4�O�E�]h�Q�T�l�Sm���)O)O8��_n��L�%���������mX���6�<@Ls��(��.G2����9��T]�nݚԅuB�(�5�o��{�6����g�,��1�	�[QRb�H2Ac��Z�&"VABdO+)Q���e��J�j�1Z���)iq���%e����؂�$��I(�MQ*�I�$ʭ&K1���s��|�r�7]��3W��ja<B�Zi�y���V��W��3������0���0t��!��:h�r��~2P��G�����xa�<C�J��.���4���H6`tBD�7�h�IO^>Ƭ�/�����x<4�܎K[0��Fo�Вl�Hό�|Lc�>����ѯ�ޫ����ҽ/��iɜ�Τ~������|ʎr�5�˥�u�cD�j�5X�b�����맧ĎކFߨ���2ht0��2���.��M����)O)O8���;�����ki��{���Xc=���s��m����V�;����;�_6���*���������C�o᲌��6��!�ƌ�p|bxD0��Є���0�g;�:8��1���:�z�t��LUq�\��Y\`a�_;��C��8J��1�b�ş�y����3J����,8����m��y��@���23��6������t
��+_7���5m���4:`���!��$�ri��m0�h���ee�[eǛm�8�)�)�q�slc�7����1��8�����zWaU�+)NRT0;6;(�!O k#�~���m�q�s��vP���M��t`�t�`�s<�y�I���{k��(ƈ'iP��1ɜ>�LF|y߷[��}coK4WKخ�������Coæ�(��ΎI�hph��^>*�����8e�a�����[�u�����Sd�9;��U��6v�3cG����,���#,��Yu�m�S�R�R�q�"<��QQR�&�WHV��Im�tӷ%��(q��.�xӍ�$�����ע4�%�bS�ɡ�K(u�e��׻%�Oq�h����YUJ�d>`4p,�G#P�߮M���S�}�+'Y�O�t��,(t48����>�Ĭ���]G��O���M�?}��|8|ZrN>v�l���gL3�2gOې)�҅Q�
R�6���<�<㉗��鉶��i�df������nh�{���qV�9���n(s
��#��k�r�7S�[��uT��5sY��QQR���U���\E����*'o)l�(� �,Elw-�A��P��,$��D2ұ4L�u"!��ej��C&QEVF�V"ʚ�1Gm*�����G��>p���{y*��2��x�Z)�;,a9	'Գ�y$��M:83�����'9��9bq�Ӥ�샢��H{̮�!!���^���{0�`����ޏ<[�p�4w�a��N_�>���o�>9�ϴsǼK�ɧ�c���P�=�qրƑ�F9>���p�����r�J���b�3d]�:��6�#dSφ��MJ�r2ɧ-9q��d����-�����|⟏�����ӧy�&���쵚"��Y=9h���I��fQ�t�EaW\���h��h����-���ɒ��d~4[�����C�����,�UI�!���i�߆��JE���B�T��<��p ���TN���l��9�t꽳h���=.����p���tue{
�ݺ�P��yp��ې�06�C�[�U���t�h�卟���;0Rw�B�8�t6f�#ad:8zho��o:ʝ>mO:��<�ʹ�L���Ǐ6���]tR�S
aL��2G�<y�y�xD�H"%��tD��t��,�B�AD��"X��N:'��<a�`�&	�p�0���6 ���6"tDNp�"C�l�̼��:�=�2��R�S
eL�|l���DK(DD����H'N�:"`�'�tN	fΛIBlJ�(�	� ���QK���JS<�n8㇄O���;ܬ�����UVW.n�7��s��wow�3��ty:ݬ�wyu�go��}L�x���ľl���v�|��f��߻������x�Z{��s��N�y'����9����%쑻�y�篗{��Ϧӽ��|����3�6�ʋ^|��jI�=w�;�/��!�}��m�sN��&A�_�J<M˾�0u[�6zy��N�{|�{Y�K�}U=�ﺗ\9N�����\�7�ڣ��c�o��������_�W��<�k�r�i���e~�;y_A��~�9������nw~�����OS�M�WL��=�+2���KU���\��o:I<�Vz����H�Ϛ�g���R���sd\X��g���g�*��-����9�F�W�t���_[G]�U|�8��ߥګ�,�{�ۛ�ky���H��.�}�N{6s9�Or;7w����s|��<��~�w�I�?��of��㐧xq��^ml�����7��}7ݖ�w�]Mb^A��c��?j۩�Q(��d��׫����h��d��u�9i��qa��HFȳ�w�;wF��{Rs!|����W7z��(1����5�K�u�/]��mcY�s�o1�7��\���>���N��_|��D>�yQ)�}�wzNXu��L��*��q��j�{�zˬ�-�=�F�7�k���ɧEş�w��'�<�'#�޲���Q�Y�s���ft��gs��[s��s3��}j���V��뿷����Ͼ�V�^+Kw�������g�Z�j�������ffgsﶪګ�io�:Qe��!ex�g�qJq�8�)�)��-I�{�{�T4S���ha����������}͏�i���igC�B0|C��m����6�2�#ܻզ�3uâVW0��3�>r�0��B��b�tӅDՉ3N�L��~�7%f\�>�=�����,Ia#������M4�9G�gI�R5f��6rh��Fm��gFǾ&�Ӄ�^69�FO�=�c�~I|����=�Xy�o�ӎ��FXFWe�L��)�8�)�)�'���z}�\_�>�(�
��R�c�*����98:�s��I��ϊ�kD��!&�D<�Ѩ5(��t�s'�v�����K�XEř��$�Y��1��/-�t�_�m�~X�e�����Q����J*��2pxдlyf�4=Q�k��C������R;P�6�o��;ac�r4C��F�c��9��k�F0l�|_�l�H�2:�<[C�=CY'{�ID!Y�`�н;�I$�n�HFr�Uv�Z�]˰��y�,#+��L�ˮ��8�)�)�jn��*��3��_=IaNZ���_����E�M����h/�T�����A�-�$�m���	��$Yf��(��-��6���1���	�ENȉR,e�H�+���1Q�o)��ɈH�jo��q �x�`Rc�҃D���(��#�(�7)�R�"j�y_�Fj?��;�:;�xqM�Y�4]�=S�cG�����]�1���I#$�0rd�2C�;�$#%�0�Q�8غ44s�#UG;�����1�@p�[Y��~�{K�3���[p�$M!�k?kvp,i���!�:C�
xbI�K� !VC���[8p��*WP�����M�e�^^u}3��i��I�w����)��^���(�'^Hw#G��u��ː6�Lq��d����.���p�ӇN�=:t��ÒuU8"�>����2�QQPHU�����H���#�wXwW�_�<��Դ��Kf�����z��F�ن+�p:>Ğ �x��N�!4<u�ؚ>�`h��k���z����L;nK0zC�6�gQ���U���\eh���ŕ����.3�����J-��|�J�D�����):o�C�?M'y{�T�3���2c�*���#N�5�����
%&�*&�4�W{e�w"^��:#E=��l8n�6q$�P!�1��4gJ�(�t��)�_8���<�<����/�|��kl�fl׾��HIC��{��E`�1rgi��3�#yG�D��sY��'N�Ø~��A�!�p�9����W�wu��s�
>�{d��L��X`�?}��0?;6~�d?s>��vD��a��RQ�"�>��G��N��-��Qͦ|a����lra���e�xv�^:*���h��g�nG���Xp~,�ؕ�ғ��� C���h�)5�C�����i֛죖IWW �a����=�J�\g��(��B�EM0�̸��|┧���r��f�\���w���㳳�z�J��m��77)���w���***	t��C��*�C�>8Q4��@��9̸��a£���U�����oX��7G �9%i4Z�Fh�*4�MX�)e���094��������5iVR�jUqt���J8/n�{Lmk�|w*�{MJ�ޭ�����K�[���Hc᧭��E�+g���Mui"�P�=0§��\����<�cl�	�Ca����G�Tm6X���Qմ�K�і��m��e�_8���<�<㉟_�2�c��۽�&���N,�r�j��c����\�\n�D-�lNmP�cE��qGpKa�k9��"����y^m 'EE��l�B:�$?B��֞VF�d,��!Q��1Z��FJ+�"e��i�bwA��`���f�i�z�� �J��<j�
;ESeV�7��_ux���3e�s�\�r�7�YtK2�~�������~:dl���N�̇�!ek��9C��O
A���z����V�2�o�)�fF��>]&�ˣK^�am���[�2�n�\-���'R��hs�hN���+Tx�*�������+h4tJ�U�6l9M���!%�V�X%!����C����ss���ptӃ���:p$0��2�\�e8pgN �2�!�J||?�:t��ӧ�U����݉ar��w�|sQQPHJK���²��ۭ����_��"�_<�O �xC~���'A�E;���4�iB�wu�ّ���<0���'�~j�ӂq$�i��*�R�,vM0��(�>��>�FQ�!-���:y	5w����/��0���e�5��ᤋ��/S;V�gE�i��#��S������t=>�Ex|68!�Dl����/�hd~��`B:x�w��'Z�徧�ym�I��8�,�a]��4�*u�qJS�S�N��κG� �ǥ��D"3~9�***	�5���
�l�V�[0S�!���o�ͅ���a[Ήjtxq1�Jr�6Xd�5\�^�]�ӧzI&�s����T��	_j�R�e�.	��#��c4l���h�&�s� �Bg��� ��	!@�R��F��[	TD�p�(6@�tQ��zu:?��͆0�K<��g�;�L��>Y~��㦮��p��%0:A�i�����׳�)vY2�2�-��l�y��çN��:zp����+jJ�̉jz****	u��'l��ׁz��Q��#a�|I��i��a[	���	l�HH,1��W�u;�����S�v�[����W�Ҕ|���:o�r`��Lhi����p����Ò�<x�<W�r�*�9��>�E���.ag�Q�l)����o�e��vxV��%N���X��Z6l2@��^��`u�6|h4 S,ql�%�sJrR�1{R�h�ߣC&G��yO�ߌ<��<�m4�L.��Ǐ<x�ϋ�E.�0|l���gŖ|l����� �D�:"`���ӆ�A؂"%tKbX��,N��0L0��xD�0O	�	bX��<'�"A,DD��8��6"X��*Ʌ�g���<�)RKR���<�:�y�"tN�tD�0N��pN,K6&ġ(��A8A<A8XG�.�<��4��0�m6ڜR����������m��]��Y��6}m�rw��A'��zk\�D[R�&�i��cbC�V�{^)MR����#��yyٜ�����۩�֢����۹�/��q��t�[a5�'8�qigg��=�t�Q4�I*%z�e9�tا�k��]Y�p��S���wg%CD�������!��p֑iڬ�4�g��՜����V��{�Oݙ�<��������!cB^ݽ\�c��A��&xw�
(�z����8_��Xq���Ɖޢ��ɓ.��w��}ʹ�����^�>;+w��I}��������,�}�����l��UuBM�H�H�F%�YR-uT��r%$���D���6�J4ܫ��*"K�q�9ʒ�o�b�V���U2�%
+ʉUQ���W繩5���mr	C�R>��bɳΝt�p������߯��}�������Z[��Vfffw>�j��[V��_ՙ���Ͼڪ�V�v����fffgsﶪ�U�]�t�e8ɖ��q��e�)�8┧�:zp��'yq��f�2b�ZE,�Z�)�ʨ��M�Q#phۂD��,wR�Y"�����&e�JFX$!2D�*Œ$!Z��u��F�㔪R,Be-��+�%�w(�*�E&\DDc�ʨ�,�X�䢂���
��(�HB�%�#����`Ь-��U��r��)S�#��R�	1TZ�nB�1'J!�FVXT�&6��.@CYK����qcFD�81e�Kkh���*�,.A��b���Q�%�
��I)D�bh�K&"e���+��Jڥ�QIR8H��H�]���$jD�q�bU�i�%�!\u\�\���Q�!G�]uDH��\mQ��G����#�F!1��j$�$+H�&�����%��ipd�0�#W�P�IW�iQ�F�$���i��4��(Ԓ�Ҩ�J�VUKd%��u��|����h�%j�s*�cwl!J�<t�I\CClr��Dr��B(T�O-E�
��Yr[$��Yb1P��d�C����m���� �$NZ:�*���D�ԕ	/ʟ��գ��:6:�Ƀ{��$��:|2��hs�@�3����6�E�w�HN�ʪ�|lp�٢����>x�|�țz�ݱ����4c�3�;�5�:�}�9u�3a�zČ�ٳAýс�p~&��Y��Ἆ/�Lh����	aEX�01ӆ�Mt��&px����X6���ǥm��/߿�C]��D���8r;:�xn��r��?�PÒ�5���m��0u�g�a��݋ٻq�\qv2�2�/0�l���Wd�<�<ۇ���,�]�<�7��"����lll�d�#�rC�J���ݐ�e��(7��p���z?pç��ͺ��h��@��v��QӃC����x(��.�f�s��h2j��%��}>��R:�}�N�{�/����)����!I)+��ĴH������\�i�#,�:l�����x�����2��ɬW�탑�
>)�N��������2�M3����
Ae8C��S��)�:�<�<ێM^�������s/{������zy�***�]6|PYZh�_&��w-;���s@J��Zr�⊭���g	�?�{�����I����CFvJG�D|˶a.��jt���J�$�����8}�2�����"nL�:0$$&�o�?`s�B˺���#��f]��#Ƈ�Fp��t��&�o�͎�vI�n�0��\�M�N��^�)������f ����X:7���?4;7Ed���e��1k���d����Ͳ�ל|ڝR�R�m�{��X���3Q��EEEAܕ��!& ���:b�=}��
g��'�
�mL�:ӄ��6���Q*uDM���ď�g؏�ş��:��҃-� �����7�h�03�-6un[c��0�}Ůٜ0�|�1�?#���������{�߰(�>�צ�b1@d{F]�M�z¼v�9�t聢�;�T%f�עW(��E�[B����s�0�IL�c�bc)��)Q��m�_)�6�T����q1ĵ�j\��W�)4�$�M�8T:r�h���tnR}2ݩg7w��Lc��w�Ŭ�����I�TTT��86�Ml�;]�R�"lB�z+�k�RA��ER����K*VFR�1Ֆ��)q'\�JEN�$�m���kQ�V�{�[u��V8D�!�8�N/w��?������7W�`����o97����H�bZg�OBL-�}w�/){<��w*j�E�5����>"��G`��I�>�>02dm����y��?[�
%!�߄Wke�m���F�4ss����N�`l<�Ypx�!���4V�J.�1p^��VhN=��;xi���B�4�Ѵv�t�����FI�C�r�I�&�H��n��M�c4����X!ZQ�▂46a�`<�ho�tD��&\[v�n>Í<��L�����<�o>S��S�S�S͸������=�=��v���U����;�T\�/f��p�};�^s~��i�=��zن�����N�!�F�$�H���ؖj�O����ev�p��YGH6��I	c�N��J�3�V�,��� �Y	��5�`�>1%�>�c�A�}�ѷ��ᛕ{���s��h�n�=���!�w�?�Բ��Gm;�JnN�Ü!���e���JWt�/~�����gF��~lG�-���BA�$Ԍ��cQ(M�7,t0����7\���p��E��!]�}[NT+��a�u�,#+���ۮ��)ӇN��:zp�,��a�����EEEA4'����Q�+U�nIZNEe(���t�7VhS�����YuޥY[=�	`Y�v]�rۓ��X[���X'u�|P���L��c��эE	[��姇��E�z��K���nH%����bB�9rX�``�%��i����$���Sh]o�[��#�G���-�p<4L��?{���n��tva�;�w�a��M|�������[l߷�oq�����i��}�~^��[>�o�'pg��SfG&��cd:agб��D!���$x���F��Ö�����qijSk�ɖ��u�XmN���:����"I{���Z޵��W��7 pM�0$n�!թ5�qEJK$�jT�DIZL���kR�/Nq^��ޯS|_����i�j�J$�c����ttz�p����;(wEF����쭄,jD�+jI�����F5(�"A�������ý�$�[�$L��,|@9�J|@��5�J��$�HrJ��
9�r(9�3H���`1XFxS���A�[���I���t��]sF�ѱ��߹}����E?h0���ɔ� (6�Y��a�Ó��8|0u,���$O6��Q{>��`q�.�&XFWe�0ۮ���u�)�(���co�����X�!o�	�HBC)Q&�,�!a�
��Ip��D5��,�&'L�Ļ˘�yK	��^�QQPf�����b��`�MJ�e+�bjD�t+$U�$�Ք�8R��t�"V�"e�b��7e�*�4,DUćIX�
Wi
����;�#�ż&�M�$w�սN�{�NG�Q���]���:p�ҥ����F�4^,�xv%�2�����x9ޓ8�R�*J�d�w�b�z�����>#�l���0� @ַ{$��ۥ��Q�iтp��n�j�Lw#���i�3��r菂&�O\�8���p��+�p.�s�u��������p�t�V��.�6w��Zn�a��!zx����`�0��%80`��
Y��0a]�m�y�)�ԧ���<~K�u�����z�⺥(���F������'����}��dz���L�l49������tG�s�7���6���+���uBd�0t��`V��g��&B�HO�b����S��Nû��]����$=�0:���8��N���;���GO�*��r?[����펣��$#I�~b�����r�C��I[kA!��F�>4x��DL8t��6P� �	��"�K�L)�)�T�+�H"%����x�H"pN��`���'Hp�B �!�D��6țb'N��̘&0L�0LD�D��<p��b"'��0�ł&�b'D����6i�i�^e����R)Ja����,�<P�A(DO6tD�1��x��6�blJ �H �!�(��	BP��8"l�ӇN�0Os�w��v�����//�X'���Y�����1��|p�9����k��3�7�D�.���,O����Wk����!��M�&se(��]��z��G_t�p�[��!� ~Y�U`CXE��]AV�5� $�n����ܭ��G��(�ި�ƍY�ID'잱>��f��Gޮt�ꓐ��[߹Y�ffg��Ux�j�n����333=�Ԫ�U�]�w���������UW��Wm���fffg���U�Uo�6W�ae���6x��)N)N��<�<�[����������hvm���f�cl�CFhL��WǈT��˂/���Ο�*�\yw�,R/��zqZ��7�f���Q�^���!	���X����e�΃e�i٫*W�_��������;<Iu������C�M�a(u��-=G��7�Ls�2k[�jk:8�N?�2�|R}�<a���駹:>4>2��gJ�d����N0�.���|�[R�Q����Q���+��ve!W�X�(�
�+�!�Ep+d+�ו�ìs���ݙ>>y��Bs��4�D�}�os/6|p��z��5��	���w���w��;�bG��g�̯3Ŗu�	 L�W�卸���T��G[��p����#ώt��?�FI�|`0��<�������v0#�|R�u���-�5�G�c�A�����߷ǶI^[Vǔ��M]_)�e��)�8����u��4V��cXF%�ί�t�N��:�+=]ggx��:u	��6Aҕw�mv����"�RH[Y$���Z��9E8K�i��NmW5&�C.̅��Am�&1̰p�-������īb�`�s!r̪(�Q�7U(�w	+�4��$D�J�:��o��GE�J�#	�.nT�;�Z�j0�OY��A���TO�Cf�^�I9��V6P׏?tu��A[�&��Ã����L����@�\Q�a��,�Ͼ1\f2*e8X�Ά��̹q��Q���vt��`�BA���`|��fh�>�%�w̲\���>/f
�[H�r[LA��0�?��.˖I���9�q콴���y�u�L�����2�8�:��ӧ�7u1�]Ԉ�)�L�**UR7��<t�0v6@�IrFS��)��/�Ju���D���7��.G��V��&�J+G�g1�ǹx8����랍����&�}&!��3����ޚ����No8;O鿑�����+�h��u���#$���`�1A�}n49�h���x6:����������2I��=?B7������da*Q�-��Z8�_��+�+�4�̿��q�SjyJy�T��F9�5��r�oW^��B�p�4V��NVV�)+��5TH�luf��O�c����������уLF��"Zx�?C��o����/|+{9���yM���j��:8xx4�28���	�ϰx�g���!	��dL�x�f����74��a҇������k���~��CgI4&=C�FӃG��q��]��2�2�S�>e�:�)�6����u����jkw�q���&��o����3�f���_\ʐ�O���~�=Ӝ�~]������ �[f���%e�׉g�����Ϻߔ�~��W��MV�UϞ_x�*���3��9*��O���vf�.��rs��ף���=��eT����9}�߻�6M{���~"���U�i��4&������Ǐ�:<�E`�|��C�9��q�LK���߻ym�4�i"}:]5t����:���]��5aT=����f[��I#4�m�dv�I���Lr�6�����u_$�,�������F}�8PxƛrOlї��	���0XOo���$���#�f|nt���t(�Q�p�Jx�����uM��)�Z�u�ݱm^�]3{����w�8����*�x��z���p]D�pa�u2��bQ���3q�F�q���t�QQP��	��s�ZB呈b��-U*�1ѕ�rT�FX�XJ\������ٕA���j��4I��ܪ�+QKQnT����T�15"yX���τ�� ԄE��9vpC��bF��7�}���8g�4=��	!7�a��Xm��=7��Z��oF�z�n��O>u���tdǟ��H�,@����7(\��ç��L���d~p�`猗wa.��CG��:�p�A��K�#�4kV8�}��crq��CaP�L��U�G�xxI-�A��{�bC��R���]v�C<~�dM$!ޥ��C�-�I&�� ���pۃc���?-���_)�+�+�8ì��T��O�:zt�����K��A���3�TTT.��]p�vh٠��t骟���I:�G-�-��@����-9a!���BI5n���k�Fs�d:\KLЦ@��������ApvT=�C
�@��x�K����^�iM�7]��F{�|�~B��&�6q��0�����UU-�θ,!�r0$�;/���WG�ݫw	#_K�et��>��ad1|�u�]u��TڞR�q�f�o�,a~�3h���D�		�:\
c3_Zq,Hx����+�~'���I�Ql�αd�}����[��l���$&�os��*���f�4���Ꮓ><�[}���4kMT�vÆ�i��^q����c�۫��Lk��d'�#�[�G����A�h!N�mL�O�܅2,��K��LiT�M���vy���8m��櫓�`��x{��<>n�n�)��3zi�&p��)B�E�8˪uN>S�mO)O8�)ez����/5LΎ�QQPDJ����	�#�����3����.F�h,��~��[�uZʾ����u�5#�-��:?%�N&=uڭ����?��2u-Y�!!"D����j�ml��f�i�jJhv�&��0�0�%��4�5�*�>a	4=9
�~i�lh׬��#C!��ա߮�XXzT�|T+��/�̒G����9,��p�����	���v���Y|�|�6���<�:���<�a��aw�<x��ǔEH���&))��S(��!�"&	҄ ��""DN��p�@� � ��l�f�Kb'N��0�0قa��0O	�$�6xO(DK��b"pD����:	ӂpN	f�:�DG�pDO������R)Je�^F�x�μ���p�bYBlJ# ɤOC!a��,8pD��N�:"`�(�$�s<p�l��{�U������y�{6��W��F�ի&��ڢ��$n��t�f��.������_=ܛ���"3Q˲��,�;a������kZ�Y���+���?p�z�,�t���ho���r�d�uQKJ*#Dj��rGD��CM��.U{R�C��-�\9�M�Jp������>���s��E��w�w�؉�='~7t��;ٚ{_M�TH�yÐw*q�pIE��p�7P�zK�A� ��D�b���^��7�3��>]���90~}r̰�����݅REk���v+�5�q��sM�GJ�� �^ei�ց5S�4�H���mש�*�*
4�m؁��&�ׯH���7��ʣ�V(�x��S�4ۍ?�v�"JQR��I�'�z�L�"F���Q�[(�Ɯ��!�y#�S�ǎޝ�Ƿ��f���]&~��/��ffg��U�Un���fffg��UW��U����3333��*��v���9�}�3333��*��iU���6x�ae�͞6xˊuN)N�N<�<�ʭ�������P����r���)-aS)E��1�㐌���"jJ-VJ�j�MQH2�F����J�EIY[$���ZT�)*#yiK.O���lh��yZR�< 7����<h�-J�JK\��DG]��c�H�����+�cc1P����2�KXI���T�t���0p�EY[k$ �☄]H!�*CpHx�VF�<Q�dB%rAF����Hd�
B��6�շ/�Z�m��r��)p��l�b!B-�Z����ګ���,"J��H�dQԔLN��'\�DjlQe*��T�m;-��ĥ�#��$gQ&�Itr�I-�%,JH��kP�ŶA[*�w����J�@�}�hj{J�e���lI)���4���N�+D��k�z�Ʊ�I6���V�TTT0���˷lF�-LT����e�h�Ɏ�6�lu!������ӱ�c*�VWա.V��En@��X�W����+q�X��Z������nZ<�umԵ�EW|s��G���>hr�����S�����0�}�z�.i��Ou�gǀ����A!�D�ǡ%�|;q�������a�>O>x�8�&����i��:-��%U|�:u��]�%��J>�bX|R����m�dB��Ж"��fF�#�e�{�3<cp�����		����Mv;~j1�ZO-�[O�m�̮��S/�|����S�:���>�%��[K���3��&��M��BB�*S��Z&<��œE�$%\�L�m0�S�g��퍎G�N��;�nG�ɠ-�x�)�8h�x�s����N��ς�f��-�ܔ��K(H�:����|�����W����85߹w��;
3���M��d_i�&6���GC���3L�!��z4dy�L���r��̆
!�Xm�y�qJuJm�)�ux���'��5			3?��?�dtV���RI:�l~;���M|?�0[Y2m�v0��Np?��NcM��s�ijZ�˪��_�ы���E����iN�{�{�����.���e"��䐘w��p��โ��r8����>��a,�p�9�!H?zK��Ι��!]>�|t��o)�u��#�×����\%Z�} ���p�va�+�,��2�m��uJ4��~>:xx�RdD
}l8s��$$$:S߂4�e�Æh��>@��˘x�f?��O	+a#����I����Â!�#���)R�|���q���_�3�L��)��o�����b~y}���_��{�'��o��c�缊�H�ֿ��k>3�r}�z��2pU��>��#�}�l~>pٰ���r����01��ٯ���	��ӏ �̼0pw�ː���>�
�.FC<��h`t00|�B���I/�-��S]e��|ʔ���㧇N�=:t���rKj�mK̌YW~˼�Wym?�o8���DdM�C�hM�M&��9t����Rdac����$$$�m.�8�%V+q�Dd��(񪊊1�)�Q�,Rc(Р��2�1S"���ad�I^+T�7R�#,pU�A*lN��[��Y�kЋ�L�B�O}A����I�a;m\;�a�����J��i�U+���房a�*WC
��C���l�+.��S#u�7z�T\0>OUn�`��'^����0=�>o�2�p�����V����ݛ3R��65	�Ѷ��zJ�\7G����y�0��EJ����<Y��De�a�\Sͼ�N�M<�<�����퓜�=�<d�Ov�r�G�������ɺM=f�4Ϸ��4��.��s�w~��>��HHH���$�ϥY��E�.�����>��������)�.6����|�����+�=�HH�XV��B�LUr'_�����I�����;i|�bB�j���7�����8�9�����M�s����wxU�nlx[޿��:|>r�m$2`�x�c�`��m����<��;l)������
i�����ì8˯�6��:�4��۶�K����ݗ�1			��`�o#���*����;;![2�(j!����|7��t�]7]>��z�|��C�P���5D]�h�#�Wo9�X���˾�����)��U��G�
p}��'YR����p9h��z:nz���x���Y7C����zB8A��˘xcoNG�u��EB���h��co���U���q������L8ˏ�6����S�:�[$����P���s�b�1��8:���?1/�x4���&J�jYgc��h�H�RS���@��������gχFG��%w���5Ώ�,;�n�>��ӞP}�r�Ϟc%T��kf���u�d�[�deh���ΏB;l5[�<��>~!C����O�6�v@�zmv6�(��l4ete�a�T�ͼ�:�4�󎧦t�av�a��d^`�/��(�Fm.6Ƌ�X�E�ix��%P�FH�uAT:�E��	�Z�&&R�-��lqʣnD���ʊF�C�e��2�<�hٹ1㌙`�� ���r'#nj$mIUV�KUM���Z\B����$�s��7v�K)6x����N�:S��t:pP�d�I������"2��������7l�&��l74�L���x�I#L����3�
3��>������^�l:i����tfI�ALp����ɱ�����6�<����I	�v���o'���y/f��t�N�2�~�)��pete�a�\|���S�S/)O8�߯*�avi��"CJ[�j��h:Bq��U��a���<�g��eՑ鰇ߏ�<;p|}��S�Q�<hѠـ�Q�â���������:n���A|繻���:�xCN��b�K(�	x��oL�nӯG�4�����:}>�	@d+�;6ӑ��A��C�p��O��u�)�)�iM0��(��Ǐ<�.�E"�R�SL�,����"'DL�"%���	�&	�pN(A
AD��؆Ͳ%���'D�'�
0L�0L���҄N"X���'� �%%�"'DO"'���tK8'Kd��$0DN	�Δ �Ԉ�$D{�x��uM��2�e�).�QL�A�! ��M�$�t�ǎ�8pDD���%�C��"^�'���_9]�{~�{�<ͦ�΋	$㜜_-�#��s�}����%���LغE��r+w��ƾ��B}~6I����i�<{�\����p���֫��Ǐ~_�����*?>Z�i}�e��]���u�oH��7���.v��ffc�EU_-*�wv�ffff}�*��iU����3333�UW�J��ݿ����|���ZUo�6��]e�q��ԥ:�2����b���ǚ�$8E-��4Up4Gԙ<��	�/�Ő{�~>��t�6T�Y�{t�J-l��v诿�BKL�3�,Ӑ�c�*��;L�y�J�&�{8L�|[�q�$H�6�6�-����D<���M��HUu�l�w$����Ѳ*�6�v���8mo�J����m��a�+�,��
e�>m���JS�:쓈��o�k椒HM0&�!�.M��(��!���S�B:8���>Ɔ�����Ǥ�\��̙6�jN�fCn����	&�IDh-��΃��Ǳ�Co$����D7��5�Jލ��]���z�L&���\*˭��p��Za�+�,���yJmJS�S�mO8��N$��^�z^�gT���3M-oWwx�D�p��8	3I�&��"�br�lv���*;�du���
a*��I$��KRyM��b���l�&R+�F��M�#n�m+NVHZ1�(�QQ�22"�,���:�D��O�D2��T��8�ep,J`�,�TVK��D�1�	���If曟�g&sؽ���ɦnJ:0�t�n<��
>0sLvP��}�������e��^��[��]���OcF�d�Q��G���`�:rv��O'�����Ӂ�<=���k��G��C����~Rs�!B�R�{��9�w8���׶� ���s�ي����bS�If~8pҔ�B�E)�.<�jR�R�Sjy�]D���d�H|��Ŵ�-��m�}�H��e1�al�w���Q״B�2������O��Fk���_Z�Ϩ`�xx������چ�6S2d9�:3E3k�'��Ä忯l�ɷ�7���8�忙�!CӼ
Ʊ&�u��e�W����0�1�W�ͳe'V��J���_��]Ƙp���,:Ì�����R�SJy�]G�#�Vf�5gj���Hpxx�?i��C�����ԯj��@�xa��R
�����ώ�?k$�+ñ�f*�L��Z8^Ux}zMG�v���3ѽnr�HI���E-�߇s�>��?�q��̵	UV]�����&���F
:lٕu�q�!�`��1�Һtkʴܭs&�zә�e�8sg2L9&�|����;�3��|C�F"����O�6��:�<���ۻ�޾=~5�g3��E�~����G�C����qu��Y�2��$��th]��J�7P�?"L��3�Ǻ���R�|��Z�U&إV�o��*~�|<���o�G��������ભ�M��w�4CFo[:g{o�D$Ï���y�4F0�=8`Ǥɣ�65�Ð������گ���|l�A��hzsF�3c��4�6ete�a�\R�S�t��O���aQ�vۜ��NT��}u�~�C���$Th����݄g)�����돻#U=�M%q��-Q��~I$����HLJ	��DJ<d������t���
B���j��[B� �
&Q�S�+�0f$�N��F*�b�NƐ�X�f1�GSx���Y'r(=�)�G��Sg�fP�9>2s;��/�>4�<V0�~)�^�<z`x��8��;nD��vTd�:�T���%[�vk���d���r)�,�s>��Cҵ\)9Y���`#�uÏ+��݉'���8����w��sY�r��f��Y��-�u���)��ǿ%��g�Ӿ�Q'�m��t�;��OУJì<���m��<�<�S�I-���s�|��ڒI#�3<zg�ɇL;6I�����C�す�a�ߵu!w@d���ِ�HHI����P�l��Bt�D6x���6�5��u2�fщ�|�!!�IR�_WNl���.62�w|�WP�*&6�*����M�;_Cg�5׹�ó�x���J2�mT��3�ț���I���U���]�2�2�
a�_>|ڞq�)�0�s�v��;�k:�5|��J�,�[�I$��X��3�|47	$��<���	�-���4i4u�����:t�#N�כ����-�|���4$��%��߷�9r^��M��oW���v^fnE�>���y��0L�L�Fd|$ѝ�s���t�(L������6����t9;�ћq��Jz�[�4�]e�q�>y��8��uN�3��3_֌�����I$����̙hv��d���Tϊ�[<��HF��c�w���I�zi��-�G���{~����J��z�#��r��,���þ�*��a���	���iGMy������3�������]h���>�7�=*�v�R�[�m���ZU�6�8���	$0hx<6?��Ó���{#�q����SJY_r��UF�`J!������8�+�?�e���윦�"  �
���C3��bҘce����ٲFč����<�74�$�&�&�&�	%�D�M�MI��	D�&�m"h�"i �h�D�&�&�2h�"ih�M$OmMK�D����K"i"D�i&�$M6�$�$��&�i��&�6�4�M4I�NN%��i��D�&-i�A4�-"hz���ɦ�5��M	��L��M&-�"ɉ�KE��ZH�ZH�&�,��Zrp�E��4���F�"Mh��"i�ւɦ��i����4I��i���,���h�	����d��&���M4��5�8�9	CP�Zi��H�F��Zi��Z$ZbȚk"i�"h��b	���bh�Z-�n!i�M!h-4BFZkDLY4Љ4œZkDFY4іM4I�1i�i1h��4��ni�4��h�"		�kF�����F֍4m4nFpѦ�m�Mm�F�5�i�A#9�X�b4h�F��-�X�5�4hu��ѭ�h�F�i�Z5�օz�n-�%��e���4kF�kh���#Dk4k4i��3��4��ѦF��l�h�#[F��8�ѦF��mdi�i�h�m�5�4F��4��Ѣ6��dhF�hѭ��4#L�26�؍b4�hѬѬѦѭ��Ѵ���hF��6�f�l�lF��m24F�5�Y�XF��l�aͣhk���B����-�����hLBb����#!gVrQѐ��d#!m�����LBbl��2i�hɦɭ�i�k4�Mf�&ɭ���X�4�&�&���&�6F�	��M���ؚ٦�h&�&ɦ���M4ɦ�d���d�d�f�4Ѧ�M	���i�M6Ml�5�h�Bkd�4�Zjh�d�F�i�Mh�F�i��F�,Mi�M4Ѧ�km4�Y�F�&�4֚4�&��Mi�5�x덷M5���&��MbkBkM�L�4�&���L�	�&�6L�d�&�4M�&�4&�l�M4�&�5���LMkMbl�5�kd�&�k[i�Mke�kLMbh�X�m5��&�6M��4i��F�dѦ�4L�#M2h�M��4ɦML�d�3Mi�i��MѦ�4�i�l����M��4ɡ5�i��&��rg&�Y�X�i��Y�[i��k	�M�ɣ&��l�bk	�&�Mm�FM��XMm�XMa4a4FD�2�"b-�#"2&"Ș�4FFXDh�E��f�2,�6�#,"dAh�E��,D�-��D�&Ȃ,���"m��4L�mh��d["2-��m��Dl�"d["2-�lF[h��mdX�D"��]puf�4F��m���-��6Dh�E� ��LE�,��"؋h��DD�m�f�ma�fE�E����ȳ"22�,"mm�l��,"-��Ȱ�l�Ȍ��&h���##,"2#h��l�Ȇ��!���AdM�m"#D4e��#D� �l�b&ȶh�2�E�DLE�6��FD�c�9a&�l�d[h���l���l��dZ,���#D�m�h���!m�h�Dh�-�LD�lFMh�"4Yh��4e�!"h��#D��l�4F�E�&�<��2�l�"h�#E�b!#,D"l�Dh�&�dX��Ț-�h�ȱȱON7Izp�h�ȴ["h��dM�E�-Ț,D�6��"�1��h���&�'4HHM!�BBE��$&�	4$$i�F�-			�CHZ,�4$$-	f��FHM����Z4��Б!4$Hɡ"F�$$�$MH&�$M&���I"h�A4I&�H$M$H�$�D�$����@G�)�>�~\�hSM)������C2�6f��ڤ�a�k�L���5���9������O�?��ȟ���_��{�o��o��� *����g��p�8?��/�[w�~斉���~�џğ�����U���6o9?������A�'ſ��{�����T ��>�����~��?G����a��Y��[ُ���o���϶߽z~����?�@�X)w�0��Q����������e��Z}�>�a���3����ڦ��T4���c�3@?��l'�?��8Y`�2s����RR�9�����5�u�uӿا��?Y	5����b9��F������O��PP�,DB�DAq��15�3b�6�UO�Z���`����A�X$-3s�@C��k����݅a? *L���?��P � fP��zÐ�m�šh��#fb���
6ƺ����/o�>�m�����	�����̏���P����������Ҹ�"���4'� *����?혜u�C� -?��;P�?C���6���ؿ������~?�k�?�����(�<��_�d�O��?ަ�����C�?���W��g�{���?���@T �����ί�~Ց���o�?�;�oO�����8�� a����P�?����`_�?����?�����������_����m���l�b6a�_�P�
:r��$�>� �$����T����� @bXf��6)�����
|u(����%4?���T./�i�h�,n7��ۊ\��hO@Ꟁ�T ��?��Q���_�������@T ��ʟ����&���A?��h����������~���~a��?��it�����S��������w�O�p?ΑS��?���?��Çq@T ���	��'�A?}�o����b�X�V+��b�X�V+��2�Z�X�V�V+��b��������F�������Y[)B���ԭEe�VՔ�J���L����ڶ�e�S(��S(���R���+jS)YE2�)B�)YJ�Օ�+QYE2�)B����j�ee
VVP����)YYYEeeej������������VVVVP����SQYZ�����)�X��YJjSV����+555jS)�Z��)�+V++SVV���jիV�Z�jjիV��(��YZ�ՔV+j)�V��jՅ
Ԣ�(ղ�jQME�B�V��F�������+5em�+j)[QAZ�
�b��X�+�


جV+�
��X�P���X�V+��b�X�V+��b�X�SSV+��b�X�V+j�b�[jR�(յ
ڕ�(Օ��)Z��R������2�)B�Ք�R���ڶ�e�Vj)�S(��mX�P����+jV�P�
SVR�+QY[VR��ڲ�)YYJ�����P���������mYYY[VVVV��������VVSR��eeee
���eb�(V�5��+++VV��j�ՊڅmYE++VV����YYZ�2�R��(V����[V�B��je
e
���)�����+j�+�VVըVՔ++(���eej���Օ��+VVVV����Z����ej�Օ���YYJյe5jj�V��P�jڵeb�����e55�jڵmZ��
իj�+V+(���Ejڵe5�Պԥeb��+j�++�[V�V+)���b�B�b�V(Պ�
նV+5m��+e2��b�X������5e5
�b�X�j�Q����X�V�V՚�5j¶����J��eeb��V���V�L�թ�+�ڶVjV���S+QY�������+P���Օ���mYB��QA[VյejիR�jQJ(����YMZ���m[SV�Eej�ڲ�+R�j(ղ��Ԡ�V(���V��Z��(+j((+(����X��V�PV+�6�V)�
ؠ�V+�b�VՊڶV��b��X�VՊ�X�V++j�X�V��b�F�V+eb�X�Q���l�V+���Z�V�յ
+)�Sj���Z�V�+QEe��+S+Vի�Q[V�����YE5ej�52�VV(�V���jj�MZ��5jj�+e+QB��S+j���(����P��(QE�5emYYB���������E
��������[VVVՔVVVVղ���Y[P����Y[Sj���(�����j�2�ؠ�LSj�F�P�CQ�S+jS)�jej�m�+�je5e2��P�P�[SQ�VP��jՕ�b�����+b��X��V(+b���X�V(+��mX�V+�������;����� � T3���?���?Bq�I�@���:���ȻI9�E�����82L]�ȭ�?����`�Si����������a|%?Ք��o �o��ɕPI���/俁���)�?�����-���~V?�_A�?��z�? w���H��sfB�#`����ڧ������@H
��LG���	f@���9��|l�?40���
]?ϭM����;�2?������9�JT�?$�.�p� ���4