BZh91AY&SY4��Z߀@q���"� ?���bR��        ��(�Md�j�d%el�[�j h ��#l�R��#A�iMj�TQ@��M���
�f�R����|�!uH�l�j��kV�2�#&lUZKI�e�l�*��,�5ZjJ��4��V�Zհ��Fk-��V"T�Y����G�tP>��m�����Z��UaViH[-��R�+�-�ES��h֪�%�[kU$�ժ�-�+M�f�IR��D�������6Ef��Pԧ��x0�f,M�  U �'�QZ�n�.�!�� Uv�сJnf��ڤ(�%f��
tu`�Y�4�I��L�Y��١CV�E[[T�cM��2�   z�@�z�v��K:�@(�u0@:�;�
tk��͜� ������I��
Ch i�wu��Ѫ89�
��ɨ[F�VW�  	׀R���s�@����v��)o*��l��xuOA�K�cT 38{ފ��Y�E�{6�<���//o<�
y����V[d
����   ��i{h�Q�u�P
�������Z4�1�9�]��*�6���N�����(�W���R�@N�y� *�K�����@���u^o)E
��vF��TTL�V�L<   ,�� 
;O^{�u���W��(/^�<��j�y�(zj@^9�@�$�;�W���k����.�^x�P��x�A���J��ʙ2mm*�Sk�  9< ^U3��y(�F���(M�� �E��{�T�
x��<J��=w� Ҩ#�7�� Oo{�x�+�-x���(
s<ͳm�"�چ֕����   6��(
S޹�� *�wh
��S�z�������P����;����T��gj [��k� ��� ���ST�B�kE�V`M�   q�= ��F7[� �i�	Z�p��P��  G;@�wc��v��F� t8�]��UT�Y�b��jV��  �� ��P ۣ���ɔ���]��Glh�nmƍtk�� 0�
nd�ԙ���
.v��V�ֲiV��IKx  ׽ hJ�@����m���@9sK( +nm�u�vkq@��ܮ QU;�{xP+�LP|�    � ʔ�� 04��{A�R���140� M� ���*T ��  @ ��$���      H��2i��M��C&��=L�i$��*�	�� Ch��f�92�)�����]��n���Ո/��J��r�tz.GA4ueBmC��|��� �+� *i@Eu� ��Bj�����7��oF��b!��HI,��Uxd�BI���Ռ���TV��nn48'�t�@P@����`|d4Bh��!�CFCF����F�4d�!��4a��� h��M�ɣ%h��h�D�$�D�0�FM4�h��&�4d�D4@с��h�@�FM4@�D4`h��F����'&���04C� h��!��4Httd4``��!�D$4`tҐс�FM04d4Hh��&�" h��&��� hɢ�04@��CD2hɢ�CD `�0�f�
2h��D���$4@4d4|4`h�с���!�!��tf�0@ѐ�!�FCF�$0`h��!�DM���4Bhɢ�3�M `�с�FCFCFCD:!�D�M04Bh�с�N�h�ѐ�!�	�F�4`h��`h�h�с�FCD4��ѐ�	��D�FG�!���$:04dчD4@�!�&�4HhɣFM4a�"��2h��FCD��04Bhс�!�	�FCF�D���$4d�!4d4Hh��E2$�0MM!4a0d� 2$4g�2$� �h��	� O4H�$!�$!����!	� �� M B h�	�BCFI!���ѐ$�	!�CD$�� OFFI!�� M4d�0�4d	4Hф:!$4B4@�L �!h�!�!!�I�D$h��	!��!4d�!h��ђ� 4d�4I!4a!4ax0�4a ф��$!�I��	�@4BBh�$<	 Hh�	�I$ѓ�	!���$$8!h�!�I!�HFI!��	!�!!�	!�	!�	!�BCD MI	 ��M$��$��M@ ���F@&�@�a	�BCD!I �2I	B$!4Hh��$!4d�0`Hh��	!����B2B0��0т h��!�F�4@�F��04d�D��4d�!����4dѓD��0��ɢ���:&�$�	�D2hɢ��2h�M4`h�ѓFM4@ѓD2h�I��� h����!�D��0<4�h�с���!�D h�ч�@с�CF�04d4Hh�D���!�!�D$4Hh��#FCD04`{������N3>�ϻ��w�%��؊AW�̎�E������kd���*��.a5��b/1��-�	�h8�&^�M�v�KGD�2���Z��c�f��{�vH��ɶ�T�6Po��d񘌁7��X�D�O��ty��%�_.(�ZP8r����1��#���9E��n
ư�W#�c*��_-������˗��~��:��h�]E��[��R@@��LOV=,]nMBջ�ϰ���v�}�����"=��h�:P+��q�a��E3�d,�Q�����k�2LUnv����������"��LIMGncG�=���=&w\�|��=>[<׈a��/�Cأ�_0�,W����aϷ��4I�f��ď0�N�ZP�@��j`�j;�s\�`��斔�_��g[��X��z�K�]Ոk�ʶf5�5K�<c��́||��/lڜ�}0�kq�굎��ݚ��H�����h�-�`"��X�VИ��J��|6�$�q���B��zph�=��� 3n�0��;�z�G$õ��7�G8^��R_���K�|���g���sg�?Y��Ӊ����x`'>�3�t�S�\q�^s�:�쌑�V���ݡ{�;�;�ƑA��^��+�C.���X��X�wIү%+��DE�T��6`R�L�b�n�5<Z��� �mۄ/#��U�P�Fl$���n�����&�T�\ɦ?���s&<��j�$/'��eช`n��!u��Yn_f�T�Q �|�+t����V�љ��������B�|vGPv7}��n�X�D��Ьm,גd90�A(�$Q+&�.홢���3��Y��"�x���o!Z��퉃�� �]�:��P����2[��'�Z�||D��Ȗ<wp�G�6MI]���upS_��v3��-r�dr[��r,�|U����^�k$hᲒƲ��Ԙ�����3���&��o�:��4���1�ٗ[U�nk��ScV��21��fJn,�e��%B����SI�.�+X#��H5ֶ����=i��"ɻ�;77}�?�z=6���'�F�`1�u�d�!��#s34z�����.2R8�?�\9m�z��]���É���}t�)����#���Q,<��^f�7Ƶi�s9�����2#uo��\K�'��<����<��+��T�����y]gO��5��������0g�>�� o��e��D�7��ٺ���^-˰�ބԉn���G�;xr9+,+H�8�ٕ�F,�(b�bf�:����Yc�˨-h���%;I�Ik�·6 ���8���cl�bu�0\/F���h�#܃� �;I٧\�秚��Nn�����A�&��$��q}y�j���F�`MҺ��n�;�z޺>,2��=4B�� .\;��с*׳ZU-T��XUW���.��Wb��u�&ݶ��/�����N�����N�X�he"�/R�%b���|�I�}��`�#�7�ٯc���х��DYi���s1��6"a�w K'�n�z<��,yo��yF&�\Y��� �a�V��G�"�� �}����}t�rܻ0�^no�o��hw
~ٹ����2�F�A�w�)�Z�^�L���pf�8p?S�m\-fu΃��W�ѣ)���;v���p^���DJ�������,7�6,]�L%Hg��߱�q�l��ZW�{�0�� X��y0`�H�-�m�sq���@cp{���W��Ļ� �^+Z��vi�
O3�[Px#4���Q@-�Zv��%ӐQ�;}�䈏JPl4n��y����%mߞ��MZ��h�t�n����<����A
��#d�86A�Syy��j��1����s͓���	��4�R���Q����ϱ����^X��ؓ���*���9 �5\�^+~r�Sy��,�W���<��Ǝ��]|����5)�p)�n��@�H}�x�g���#2g�z����A��߽h����0`��nOa#N�'�\�ؽ��]_k�Q ��>vj�L�B���;9Z ^��oq-�����E��ܫIU��"���ee�&a�!�T9��ô��	��g��o��<�(�	�	m�b��A�b�z.�X��w�S!?O�[ ²0}���.$�5\�=��A�y�ȉz���z����H�Uњ�o���B-��g�h�M~{1Hu\��-�����IH��Wh�Ӫ�{ m�Md��s�^aSpQ)�m �O���b��%[�!���y�!���i�G���{n&%��<(��=�L�p���1���%2�e��_<H�_Bf?k͈C�eB���>�~fx��+��q���ꟍL����]^J\z��Bk�����$�A3b��%�w�m:��򯺯v�m�@�����wvP�W!����Q�MR�Ըw�lu�b�~�/�n����(��`2�Q8���AYzq�,-���r�/m��>�قO�~��O���i������kZ�7K��b�)�kld���W[�E��i9Vz�%�V�#�I'��5y�щ��c�<��s,�Ȼ1�D��\5��F	�O��꙳��5��^>�/���f_�k0_V����7s��*!6���!_-XQr��X�����d四R7��}^�:�ԙ�ŧ2���F��S�V�ض<�=st#�BI��j~�S��n��ېz�����w�z���킋�j��q�$���N)ig�$�,.:nO�$�l��=KO��d���[�-l�n tx�X����P����5g���_I�?/�ݰ��2x���D���![׀�ըU�๖��I�
��,��
���ieV;�+�L�ZX*3D��\��!�d۠۬�ݫP,n�!Ex�-T���Jh�*�R#aW�#�5̈�ZՑTN#~.�u�'���}�"a�(��э]ᵾ~c�'��d��y?Q SN$�4�8v�1���<+PĈx�]D�Im8���ia�w�����9WS�\Ʋ��P�-d31���n˴.j=�kի60f����6�3��a��j�D�Q�/�`�L�tl����U ��hɧ.���t4�yMc8`��ܛ|��cr5NS��7��I�:���x]u�J��mY}�ow�}�eK=@<G���M��K�JR��L�9j���t\��5#��<�xyQ�����������1�6�G���$�x4�$een��Ѫ�!.r"��m�W���Ì�j+��2���D���� �i�9�� ?[����s*+oMBԕn�#K�iB�1G����RQ�4����p�fyk�/M{�SF��#Yv�!�)�:ؕ�6����x��d��6��9���1�1fWP�rj�|������p'�ʬHQ���N�uvg��k>0nh����r,�#ۮ)[Χ�=�/_R�=u�Q,�?��rj"��d;i^���FƷ,��!n�Ą�6��a�enT;�!�
|�(�-,����OV�/C���-�jg�>[�7�3/��?\ǱKT̘�Q���^i;H5��0�cii�W5.4l�4i���\�¦�-i�^<o6i�&�o���f�&қ�س\t���s$��DA��bǩR�n�r��E*F�q�*�DգV�cY�n�"�!�7�o�//T����F��P+[>��v�� ��f�� �5�Q���w�l��E�lRg�yP3F]�)0� 5��]i���2��Z������Wۧk��5��^A��6�̻{b�C�M�3f��
,6�f��f�!�s=��7u���d���f�3�;�݊�o�s�Ac���E��If�R}|��'��;�F�e֛Kf�C�H%/)��w.i@�� �1�������ޫ1,O�813�'Y�0��-)f�S%���g�aJ��K[o�3��hħ�ߩ&���ܙ�Fi
/z��=��I�ʦS�t�'���c�zq��/QTYX˰���I�q�줱�[V���<�a�yu9�!L�
 &��|"1�7�eWqo���gs۳}���S��=[�I^їT4�17#"8���e���#F�~�i�P{sK5w)ÌY���b��E��5ս����V�N�;�Vt6/[֛��Z����E�J��{��y�FvhP*p���sX�mB`��
��8��SM�[հ�`����]V-�ǹV
�7�QM�x/�@�,S|�2a �f%���1�a��@�5S�~ѻ���!<���2^Kv �gU旃MVd���������L��f+Y\��!ct���t����JMs
�U'��m�Q����zH��8�p�����s�˻sS�n��I���|9�Vof���K�y�(f�E�|v�ٗUP���3�"�z�G���uF2z_QSr�ث���^o�:]��1�	h�dSD ����eM �^	l�0m�6_nYg���ۧ�M�OkM�l���ø����/���e�L�A��r31�2�і��JB]lwF���܄X�bÄ���
;e�`lx徃�a�ԕG_�P�;�к��.�E�%�P)�����NzJAԲ0���fh�f׶�>Ly��g�bi���W�!�G����	�� i�<Թ0��F��=����a�9E�Aw�h�:5b5�vZ
�DMTL����e��o�2[�(�hn�0vrh���ieЩ���Z,E�u�[�S`�����F�U�ўNe�D ����+����|.���{C�8S��}��[==��ǰ���/�7K~)_?��(�<�<��m�l��*Fj�
�rL�u!լ㽆�9uJM8,kd�Ю]H�J�h����p���'*�<�4{�F:�9�!��"ڼ�W<�����4jCo������J�C�Z��7��S�UZ�3 P��u��O46M��+�5�@v���iY<g����5���F�3l�Snw�3Z�~�U@2u��%C�sf1�1�'���b"�T����[d�[�7��F����d3`�j���(�� �&ٶ{Y`���VB�7Uت��7>9�=��6{m�=4�'��V���dH�FF��;*O��B�CTۦ�4�=ٌÍ魃�J=a����VC���s ��-�\���.{v6��l���Y�t�ɚ�,ne%���4	�u�l�P�t5/a���Y�D�V���<������jWg�X�]�Nٴ��z��u�ӈ:�X�LV�6��d����$����cD8±s#ٌip�cv��T�S�F����]�3Z�?I�ʞ4Ob�ٱ뢆FAx��t�E�����(1Ja.G�u&���g�`��acf�����2�Uy����\��F��wB�<u�����'1U�<�)����r����F,v�JƑ+0���`�ÿx��t��8|�g7�U�	�仾�銑��s�m�-��u*^��4���M�}�DP�{*$��*^�=��1�׊M͙A������Xc^�� �Gv��M�Q��*�p���T�t��%J���,�M�*�j�v������%Y0]iS�L�7pm;�z�XY�x����sʠ�*i�����16Іg��re��I�����Z���ڃ~�h���E��X�Q�isfIVlUf<5e�5n=�&��si܉ͤI�e�l�;B��p����芈����9a�Y3pn�W���Y2��3V��?W���ۨ�{��uY>r�|�{A��5\����^}e���'�հRq]�R�ҁ�+�����(�X�
W6���+��L�622	Z�P�jl��Z�͙�5f�*���K�1����֌�k%|�̝�&k>���rI�늦�&9^5ehŧ��p��A�#��oj�*^��+u3����V)ïn����4M͆:9{R��Vtܬ�?�m�ݹ��WZ|/X�YT�B&�����+thvOo�uX�a�IRgt��ţ����(�l�o����zG�crl�	����@��%�,�T���V�pyX'�T1ۛ��hq����Dg�C�j0=�iʽ����i����TM=@��&�w����/����ԫ!�3V݁j#wYG!���H
� ����v�J�e^/����W���2�km���4�9z����3A��2�2
Zkd�57\�Th�n�M�;W�_@�z������	1����L�F��3�Pޕ<����M�ࡇ����P��K�)(�ݠ��3ؙ����f�n��ً͜�cV�)��u�%�cD�t�e!n2��o�][��-~�2dD7�ݶI�����c�{��:I%QQ��Hޕfd��h���O�LF��~��������c�V#1�ˇ3(�����f�YD�֖ �\�l�$*0����4l�hd�SקK!(K�_(�`�=�����s嗀��Ϸ=fj>��gȏ�V�!!�T�ͫg�$���(���YOT���K<��V}�n?L'fX���Ҡ�(�
,��&J3YF��=xn��w�Yӳ5��R"S?ǻ�o��_��\g�UZ�I%���l��Ā�͝0�W�Tх�:a�ʲ��f
�L0a_�(�S?���i4S�l���h�X�4)��ۣ�A��o�G���Ӕ�;�h�~[�)5ID��ِ��J�Ћ$�+M���e~�*�:��F�(�f�3h4��ǛL�L,��:��]۫�$¶�7��m鄔a ([�l���tÇ(:�af& \�T�Q�A�$�e�I��t���ִ�e�?N�����{�4�����'W��~�
 �t����̋�����Q,�bv�;��^*k�m��nI�Y��yf8;�^�lfTǗn[}��z�sgo�����Y�(pѯ#�|��]���o��X����Œ�gQ�z.�ʥ]8iwTor[Mε�U��u�g��]�ޭǞ_K�K���W�[��Y�`bҵ����a����}*$�$���}�١[י6���K�^�X���7��'�j�(��|{���Ǧn8{uwD�sP�����g�\aA��w���lǟ ��aũC��{u���N��o,$^�~�����w��<��އe�Ȅ���|�!�`k%�in�L��,���u#��e�W��S) o���,P��k�n̓kY5�<#Y�2M��Z��f�Z2��Nv_^�<J|�)t��T7���bx2
����er����4ف���7o��g*U8(8Wv=��\3����v�
�dU�Ɉ*�HmȌ�sz9b�En�m�X,���Hr0�F�[v�OF�ά5sz��é"�V��R�y��,䲬$���<���bw*q�35q,��[f�k3;Uu��y��l�0�H3�����dK�n{˯(7yC:>�yϫ�j���]7�)6�,⾜�f�z\AV���SOU�Ue��o.�v����w
3�l�B��Z�]eڹ�'%6�g�2�ٺ�ٺrՇ�m=%M^����([�7�[;�y���2�Z��ᑣ�Jq6�ϫ6>/R�z�̾ʇn*��c9m��2�z�Rst7H��b4�R����7�����#KE*HNb��U�VQ�[1	89�+2:�|�*u�By0b�<s�o2�,v�^�JV �;\Z����m-)���V�6h�8�yѤ�z����j�s.��MP,'��qn�ś[����7|8�"�O^I�;X���KP�>V��A
�u;;h��K�J�����ö߼�����D�H6�{��D�����.݋�CS����vKBڢ5���^�{-N�Uuwy)�|�N�WyX�u��e�_;��=�8�c��Lr�;v����A��I�v�Qp�8S{����1�����&��_m&e��\�\D1��d� v���D��	#�ylz�����^ ��#hH�ؙh�9��0S��A�]d���*�-��]�{W������=ҽ3CE�/C�����X�
��$֕��o�F�͘xS���+k2����,�м}q�vL}��I1��w�׆̯���'5��.k���:3�ɧ�����͎ά�Pm;����ƺ�1^l�΢��D����b��D8ű�"oA�c�x1�e�<����F�+�w9l�՝-�wy;p({^��2+�R3vM�v���L!Q�bQ�2Z��Mu��N�8ur�Wc�z-�Ύ���Cj# ���HrT�}*�>�۵�7�Nݱ�ش�v��&�o^��zޜ��nnWP�ZH��RP��;�}N������<�ƺ+����X"�:����Ij����-k��!c���w.�-�Ӊ��%�zW}��������S�O��/|�����*�c4�UrغK�*��̜�WKgK'�t�ӫC�K���,5j�Zz�����a�	��K�{t����v�	������Xĥ�G�ڷC��⏬'����!��� �xvaϥ-"��ʖR�g7)om*�Y��"����p���/��U]Rn9U��=�u>V��h^<�:�4�2��\5�⢚��W�]�����]K��u�%bv�:���h�������s*�1�d�]y�î�"��=a���6�������Q�S�f�f��Q��تd��}�<�ի�{���1��*]��Z�.Gm���-�FdƯ�G��v��NX��4��~�@��nw��3�� ��T��g�ד*�Q�G$KoJQs'k��火���M�OE�c/\ڱݨJH�۳bv���h��='�8浩|B�^�����u/[��>1�F� ����̕��g��i{��|�rC��<�ݔ���R霯�7w5L�g���s�fo��ܵ��>��.b�.�2�Z�C���AV�\�9^����Et��gb����.�P�x�ð	�֬k�͛�Vb��S33���+�3T٪�GOx%O��H�\�//����B#8ˮ�]�����³A��O�/f<�6~�*˯��|F��p����ѩ��	����B�k�<��BZ�ޘ�������	��Z����^�^��o�Ow}��zu�1�N7ɥ�L]�g�x�~�'ʠ��׏�;	���޽���e�r�Ey�Ӏ�R�5���S����S�'�2���es���[5s�7��{}Nv!�u�Η��͢6�3*��.,[/)w%����]ɪ􅊋�7Q�b�כ0'7�����ִ�:�3A�ܶ�s]�wC{L�@��w+���YwO����>��i��bд��K;�α���}[O�P,�`�����mL޼�]m\�tZ������y������#�:Z�/;}\ړ���[�a���{$2j�g���^8�g����49�E�u���]E����TnkEC2U��a�t������׾�gԽa�s��J���D���٧T�wA�YA���Y�0{�h�\r�<[ L�c��=�r3��=V>�4qgU
����}�]S�+�t�c�ǻ�c��3p��ۛ���hz��ʴQ56$y"��(gl�}O��-�1U^�#�Ҽ����6�(ގeWf���x=��{,�q���8����w���9�?Dא�(��zL0H�]���q��Ex9W]��nMaf�w6�m�pM���{��h.�d��5��V�p����V�`�wA*v�;X(���:�!)�U��CX�["mfG���pZ�W<��m�kԉRR�����r�UmKHf���	�`�t���,��-��ǟ�	�f�vv����c�)�J|��	I�D��Ո��]N���G���~�넴���f�,���mB�7�y"|h��@ד��4�}|��(n��gp�)�}�Q��9��[.s��#�r|�<}כ[VXu^��^��6ZB�w|�/Z��g��<��XNX����:�^�MŃ�W�ܶ�m�1�p�7���7v2�^�}|6�1f��k8�/��{D��	�PECM��"��n1�2�ot.�v8�ݹ�۽9��JF�^�q9��A%ݏ�+��orӊ�K����T��U�]h�ꋎf�w��9�����:r�����7�Ļ����y�<rg����ڜI7D%���U�src�S6n�[�;HH��C!Ӆ-݄���7��U�2n���yV�F�����x^�$=������ᆒ;K��n��9V�)X���7�w(a|rJ��AQ����Q����B�������٪�-I�:����if`�I;#�:a�����ntOB9�����e;�٨u�����Ŝ�~2g��{'�� �n�ҙ�[��w\���W�2�Ƹ��<u}5��zwyN�d�����X[)��e��o���iK��l��GQ�x��GV�"�Ge�uX�i��1�1��&΋�މ��N����G8�9�D����j�싔��u�����a��{��%|e��Axk�ǫL-\��0��k:79,��!f�o:�u�#[!���K��H����-��*F��[�����I���f-�m�P��9��ts}ߧ�i�7�4����w�<��ʓnwĕ�Y��
����[U���5��N�6���de���W�%�\��u�������ٶ:�#�t$^c��H�)�+��ü6U���^\�%{���殼a˧{x�Ff��[�[7�CE�P<����e���U�y���f㝺[:;!�K�kT���z߯��7����FHΔ�9$���V{�f�"U�1)�ݻ��ҧ�iu�h�Ӭ=̾:_�	��s1]�ӻ�����<U܇$V�>F��Ǧ#D@nX�N��Q}Uc��C*�3C�q��ʷ˻����k$щ<����1?����sk�Թ��槶(&�PgU�t�ij�����2T'<���^���g�竩N��]h��Y�o�,���_�B���&��u����LIZ��9��8u�>%b�zo�t�<=3ْ1�Q�*�R�qt�������\}��y���{��IZC�Y��n*..�U�{K;Q�pv��b��\U��a�V`a��#{N]�D6c����X*��0��7�,������9�c�T�j ��N��y/!]ܔ�]u�ٻC"9�ߧ�1g���k/l�������pU�8�vj�T��&�\`W1��MS���xwx=�hpOjc�:g��ڐa�v�=�����ִ��1�=��}�jzv��}��z����d���h��Oo���̓(7����p2�qN�^��+-��睄i�O(��r��N��k��4��"&]WZ��v������Y8��X4�{ݘ8�=۵�g<�"G1����I��.��YГwʥ�$h�Gn����t�ѐ��y2Dʫ��cԱ�þqx���b��.��-ӬuO�ܚ�1�m�gn!��\�̒��cQ�����:��/LY�_�,��ŁG4�z�)�U�Թo��	�t���Ϛ�̊r嫠0vl��+�C�k*�qd�N�`�wk�yk�}K�'��~a<�/ҭ�ȕtZu�p���9��	����Y�&<��Q��E쾟�f]o��9�"税��A�1E�#�9�"�&��.��G����;X�h��-��>�v?9x�)4Nr?�z](=�w�Fs�����e\M�&Ywڽ��\��ӄh�<.�iN�]$K=b]�?���j�_Sy�w�a�v���=�5y_�I�h���B��O^n�k���@>���7�a����f��{V���ά���4_�0������hhkZ�O�����V9�`�i�D��|�U���s��7���ɨ�,�Iۨߒ�G]e�)��,�{0�;u��:���vx>��;:z�}=�Q�!��h�ʋ���Yz~ݙ^q:�=yafe�s�U\{'$
�)]!]DIu� ���ݬ!��M.?���Z�D�Ԇ��P�m�'|L3��ؼ�l����x$�|�� e����=8��ކ:��x$��)�}�Y��W�hN���"=�P�\���ދ�S;Vp^>��t��4e�^�܋z?pYޅ�(����#AY�X.���֟׳��qe]L��9���71��� r)r�m��筿/&�q}^��1\|gW0�<�<:H0QۥC�S�d��O,�'���Q2!������8��8�z�,���T�|�%�"�����s��i�z�Zx��)��j��v��������U�}�8�Y�;�
�v���Hk�*eV]��8g��'�Z9U�NE�&w3x��%V3h���7���]�Wݓ_[��yT[R�)�܆�XZs�A�H�s�s�K}�W�����s�8o�zf`:ߋ����a���yuǸ�����VV9�NV�]�'7�,:"$Y�5�QR+����K��_9��J=x���|�a7<�h>UP7�]%ܻ�B�-U��t�ï�Uvd���>��ʗ��nY�<��T���M꺍e��R.��:�Z��fpt�=�9J)4]�sI5n�{N2��=9��:j�;�O��^��A�듦�w�&�������皟�>�k;�T�_GD���}'��/�!\�Sois�=^� ��͊�Ju��Ɔ7[c��� ɇ�)�N,8�x6��E�iǉ���
�a�S
�i!���{��z�>��=�|���;m�D���:y�rt8�\����n�Z�T]}G��9�r��AC��>o�:����ucV�)*���v���]�?���^�Z{��j�����T�Ş;���7|�V�.F�;��ς���[I�g@�.]��/���n빀�/A+-835�Cz���hn6ٻ�a�2���D��[��`�����1^:���;��D`�U�ܱM2W)��=t���o���_�@Otxnx�9�t�͢��u��/`�׽[��%]̊]P��rE
�n�7[���m��m���pœmb��Գu�jF;xf��le$��֒sm����ux���O3��n^����$�{9�m��N�(��n�0i��َ42��IT9{�s3�KBRk��FKUwi��kF�v��V�9��+�/����U��'[gv8�=��j�f��!"�s�����1�ž���Ev�:A��%}�p�^,�B`w����^��)��\�֒�J�n��ar�e�ʹB�>�+��1;#��u�'��x�a�j�υ���կtvLoc뙮[���.�BwtJ��2��q�)�vFKG7욮��1!�.�P�0�h��w}"تP���Av*7{8g��S����˦�uۙ2�=��\��],�:	�k�Uj�|����#/K��+w�Wl�f��<���\�NN���ԏ�j��\92Ӈ0��^�S���\�阈`��p�#0E{&�£W"�I��Snբ��VIR0aA!%8۷����"��*�%X�tZ�	��F�_T�r�b (���^%�o�H��a|��p�H�i�$��y�`$?������H�DL0��D��Ca��L����k~����-�`�` ���Ķ�I��| ;��5jE"j�1��B�.~؃"0�Iv�ش�.܈��A��&\dU��B.�������,*b"M��m�R� I�#�H"`$E)�E�.A�'�n�
P%��q%O�K.D�\�v��A\�s�CHD�P�T	��G���
��F"�J�T~r ����ٯ%�)ˊ�"�%K0Ô��G�\�!X�H��#4)E$��Ab8J8fq9�fv��^2���|�'�S�μQ��	?O��FB B@>M��8�_�^���F�Lc�n�{ilNy�uJۥ�,.��'![�7qP�^���%�ץ���^��A���dRl�&,��\�X�Xxܽ�qFC���-6oUa<��wQ8�F�K�sP)�yҸ���m>۽��B��T���&^�9�z�x��oVmrj�Ǭ�-t �ep�d�pu�����ŴDeԃ���˖��%�p�x8Y���;۝�[ӑ��fP�\R��\���6��{3���״Qk���K.됣��ˎ��>���qM�|~���8ǻ�Y���hy��*+��<ǆr�j�z���LІ��O_n~�514���,hP�ӂV�X��`����]�[��	��!�qԗ}�S윥��Oz�X�)&5a��ؚ0�������v��1�7Ž���m
3s���=��x�F�[�l�7NZ"m�TcS}V������Ag��{��Z��	!��*�y�ۏ{��#�ʽ��Ӯ��"�rZ3;�Q�dx <w�'8h=��1y17
]<q�{��2�"�W��K�+&ɦ��j����˂T��!k����!Ej�b�Y�2�v�L�i0�Z�M���7|�����cp�{�;h�'>�a
T�j��4f�=�2�RHN��m�2�a�����<�ʓs$:]��c8X�A� AA1 � ��Ab  � �AA@� �A b
9b4U1N�tI����rt=���u�P�/L�ץ5y�X��%���|��n����t�V�ҜD�O>��Ӕo����5�$�<��+!�Tt�adj��b窆ge�o�u�6�����0}�V���l/���˰)��٫`�nN]�B�����՘KzAqw^~Λ��&�zHɳ�f/�`���I���4�8��J��䲺��	���|������܄����Ʈ�}��ev[���f�=�!2�y��H�m�����Lڱ4�� ��|g�@����	�/�UΧ�ᒢ/��!�,(vR�A��E�{�A��SQ�U�:�L��d޲�yM�Z�;��).xV��b�ie��h�����֡J39s�ޘ�/���T��"_R��oq��-w���{:�)c8�R������3QesIA}U�;1��3�`�sS�N<y熉y�"�����xR�o��]�R��lt7z3�V7͙h�ڄ(��(�7h���8�d���5�����>���1�[�S�s����^�O��* n��J[�q=L�69:"�T�q�t��|�D��b�~k7�;&,h'�vh�E����=��;����1΋��rz��2r�z�=��]�X�W�V��(�{�<T���Y��6���A��.��BBw�]���!y;���� ��A � � �AA@D@AA � ��AAA�X���l#m�U��}�퉟.:�vu�[G
���1]�*>�㙺����I�ԄD�o��V��w{���˒m����N���s.����p�lU�2�^%,M]�V>�V�ג86#Zv[ɨ'�o�Uj
oҬ֧\Y6�,3J�/u��"�i�q�藟������f�^m�ǅ֣J�k-�ZѲ�-IB�C��P�W�
���గ����=�;�]i�}�9��NF�i�����b^�z��O�z�<7g>�4PP�[��;"tn�]���4&�w7_T<��&�]��v�k.�;�� [�U9u����Q����(=+kx$S����5:�)o�=��={���y��I�bf8��;����B�B�&N��p�w�6�x��\�Z��[�2�s�>��.(�����|���P��i�Gu��)Ѿ�hd~<��1�|�d/i��I����FV�Ȃry{i���y7a%��%�Y�����y��O��{}����.4I�C�&݆J�:4,`��w�[����A;2 -��_Hf������q�:�5��w�0����Ϭ�Ǫ9=U�s�Vo��w?\���Ӻ�-0�+�=�u��E�곲�j�;1�p�X�<w9�z�u+FV�6T�e��r��OS]x���Ug�Sx��4��<\XR�,�4X�� ��A bAA ��� " � B(AA1V=�wN�Ԓw�EN2fjo��avZy�N�9�8���,ja��<i�y�l��x#�{z��*E�v�j����&
����{ �̖�/!Uj����:�9�����x^�Q��&|��3.ܙ��\���t����n
��/����!�7�w�<�dn���Wo�|��oJ��hV������P_^���T�3gohy˿����P�ȃ�Vr 3�%��q�7�5ӷ_�h�E>�ȉ�V��w�� gl�f`�2논W.JKpQ�V����h�'ٖ�~B&�x��zx��uf��{�&���.J|�V�s�h늴Ah�ى�P��b�Ϋ}%��l>W���ö���2���M���d�g�ek��8��M����������dw��Ò����u?��X�g:�NAڳ;&q��í G�$��3�\Y��e���vj���ϵ6�T�$ɝ,����lɾ�yRN
B0���<u�{�y]����̩�(c�$R��Dp�%x����OSQm��I���Iڕ�;�;�wn�{|ƎfK�9�c�*���"IT�H�n�J���4:b�p-�r��])=���X��V�d��j�=%��=��ȸ'V�}��a�n���t�P�g{ݾkM~v{����v(͂�>=�_"�v�B�CPJM�0��i���"�#F�v��b�8@�!A! � �1 � � �,AA �� � �$Y�Q�*"��b'��F���,��BM��5E3V�>v�����gT"G��i��=r�aܠ��v��;�<7=n<1c�oL��_�����)ve��I_1d���5�H��]}s�������ֶ%}���f�E(ܔ��ƴ�f釡`�$und�(��Os�������\�о�o�ùj�F���k�e��u�F]�/�(��I��ӓ}:b!����`a{�z�e���mt�rI;;��Ү�;�Cd�v:��,��_QX��|~���p��;�ḳx�
м�%�!�41s�ֺ��>���p�.�ϝ~+�ϴw��L�S᥆*f$�<��*
�3�]F�ֶ��qX�!���q��%����^.fr[H����]2w�o�p%�*\
��P��S������ԶE��7�վ{�����||�Yk�d��3�M���S��n��n�%k�[�!lV�4�҉L�EQ�Y�w���b����gF���"���zk�qn��:)��������ӥ}��i���q���F@�&6��GR���z���7$�ԡ�Ιc�'a��_M緤 �j�c�`PL��:�G�򪛺�Oe7(n���5���.\����'h��O�ΒZ�U�k7ʬ��m�����p�fǻ��c٪A��yy�����5�N@�9�&h*#��0f�6A7�x��Pу1 � �A� �� � �A�,AA� �A`� �D�9�i�g,�[;oy�k�	 d�����u���ZLCqcG7�������i}w\D�(b3v;*ꛦ��Ӎ�Rf�j�k�^c���D�WPD��j�^�3\:c���3&C�uDnNG,�9E�����mLu�6���)�"����DsT�}ucc�Z���mvo8��S��Sk<�>��q9�:��<�N���LB�^.�}%��3�P�ҕa]0�3��f�Q�,�O����n8� ��4�wi�}ؗ�ҕ쨓G���eoY�P�QgaH�W�DwH'f�rVC\��L�ܕ�9�"��=�Ǻ&�xhK���cY�_Q�����{���(Ug��U�,�qZ�Ǌ�5uV��yzk�fwN@��\d2�p�N%�����7J���M�)�d�ʏ2�ɼZ�����a �v���Q��d�U�mR��!Z����6zV��.6���'��,Cл�Lj��G���/1O����[Eh�/��`���nō�X�O]��N2S{u�4�[������*i��6ߋ��~]؍�)T���/�R{3�g�����e�9�3��¼+B:��y�-9����T1���QMp� �u�!�]J�Bjޗ�7��no� UPkDǸ��a�G���,FƝֆ���9%��	�3�,!� �Ah� �Ab �8A ��AA� �AA� ����y��(t��oj6*��0��'*�c�@{k{"�a&���z�X���nvS�'7�nb�d~�8�`����vmy�L��2+�����LT�����*>|D˽޻�z�PPK[�@o���敛�����BS��R5ze�p41��q�������.t��&�[�-�����x�����W-�6l��.LQe|}�z���:z�H�[i7��#��^w�hS�=~!�˳��D��g��ˑ�f�c�*�_-fm�h�'�j���5I�f��$	��:�,�!sZ��G�4�g�&�+��x��%����3��k`��]�&������X��s0R>�V�ݱyƏ��o#��Z��M�x��n@E�L{WI����\=�^ʉ�x=S�լ�`���+{	���+uS��ln���t�ll���W��f����ε�tP�.��մ�����Uj�o�w
�8P��k�ʜ�籌�v���V�:�:fk2d��&'KB��hG��]�1�9n���@�fVV�~p���ժ�ܪ,��?%e^]�]G�������Ee��m	�����`��ݒx�|s�ӯ9����7�n�
'�2eS���Y׮#��>z'2�i)GKH5w̜Dhێ=j�k���Ϋ�/0�^|>�~�vMc���5�,Z�b�B�zF40�Ab � �X� �A � �b � �A� � ��Ab�F���fS� 󔗦>~7���e��^������:�g6������=8MG,JU�ʶ�t�0^Y�F|xvS<�)���n�8��;k3.�Z+��lߟ��{wc��q��y�$5�����6n��.����5'���Uf��.������߽:S�P�ԏ���{�)�����fEྠ@��{���4� �ږ6<O���S�j"r�A�}�	��A��!�O��������9�Q����kI��h��P>�}��x��L�g��O":Krp[��K�G����RG���tދ���|ND5h�[Q�x�o�?��n��bA�5��|q�j��6�9q�ʍ��@��}ٚ��S
�~L)��ͨOJ���O�'<�{�ɼ'��6o����[�z}��f�������"������������L���1�8�=iT�eVH?d����R�Rbఽ�w��ϖ��u7}�t�,�R�v��0+K����^�׽Jɓڃ�o�uE�y��{:{%�K��~j9@�=8}�\mܩ��P��pe���N"�߀	�&|j�ic�7�g�aG�a�'Ж�������0؈�5[ѫ���١�R{B��͊5������s�$!@ ��ͳ������u*�3��d\(W'�:��X�����k#x>��Z����DBb��<�	����GW3	ڻȜ���N*y�-a�8!P� � B� �A �,X�bA@�A@��@����:8ɋg�쫢<�7���%�v�����	�Z��c)�BJ�U��v�QќJ��������dg.�,���z}CB����}������S�x���'Xw-�Sڽ���љIV���!��]'�:�	˥[a5XqI�� =}e(���i�s�o��JN����I��j�B����X�����ߺ�h���ӞÞ�Q}�簾��l�涛�n�E�v�5�1n�C��P�rʭ�'���5�<���g�{��\Ꞙu���5s9��G�u>��:���}|1։�i�	W�u]��8u�Q�=�Dg���R8I�_N���x�糳&�^{ޥig/�}#|Vs;Aٜ��ǂ\���I����H:�k����)�{[�{�IS2x�t:C�D'�+�&R7\��u2�쭴���V7�����v��d>Z�;�J��_�Z�3эb��#㯩]��Y�S`,�����ՑV]��k��?����������{�y�H �iVo`�'���8��E���^oaN�4��|ީ��ީ��[7D8h.�X�k��!�����ͥ�LVh�H}�C"���e��R�N�2C�2��ƪ��2w"67"�݈���b8�j�='�Z�͒9�3S�R&y��X��z8���������k�O����m�<��;څx�C9M���w���^*�!.�VCu{yK��T��0�i]6���k���n��L�	�����.��sڑ�}����t���Mz���ޙ6fB�`Y�/T�fv{G�6�3[h�)48tLh�|8��~^�,]֪��ԝ�<Ċ�(V2�Y_U��k�}�����x�r��8rj4�j.��1B4�x�B���Jt��7<X˵C\�����t�U�=,
����0$�v����Y�0o6Am|����j�T�zt�{����i�i�)�o;V��<ki�A���:�͇K)�p�ĕ��G,���}�	T�D��,���[�J�J #��J=�p�ҫ2�wkQ�X�a�7�mԱYz�k{�2ҵ�����1�;R3V��9G���/�
5�&��A��2�R�6\ �7�a����U��/�2�}�d����1۩�HֳG�������~Vja/M�n�њ�B�νv�.[��^ek.�jCr����Vn��RŔ�'�<g������(�<;�>��DL㧹�崑�!��i��2��*l���S:e�TךSQ^Vz����q�K1�����nX��SZ���*��J�;���>�l��=�(q�6~�ۣ���]!���ɺ1v9�{�Iq�(<�|���柸.$��z�V�&�u�`>��g�\��a�h�=����O<|��I��_�D�\�7ٛ���!}��c�|���s��I�!>{����������������M��a�0ݻ=��M��ZJ�-�Z[h�T��'�0�l
�ꐢǔM]�����:f3��<���O�Ϋ��@��}�Ny��īvd���be�|�	�ɦp2��*��=�Sۚ��g��w�z��fXA۠�1,�o_���;�gq,I�w)x��G8JVs�����M�2iS%|���9r�J�C�N��k����2�v�鼺9�,�x���Tz�|�4�u�9��o^����?
{�\�4$wL�̓s=�z�ؕ_�1\�����k��Ν�sx{#E�yOp'�k�Bp��$�h�s`׻�@KX�������Fz��Kuջ|wFc_9��2x��ДU�F����ٵ��w
���:���*\Fj��{��ʕ�-.zv�^i��5$�Su�|�����;{�H��n�Gx�����1/ޯ.���s�sY���w��[����$+Qy��մP�Z�g[6�1j���.6���ɧ]7�,��s�8PL�a3���sl-�fxw��Y��l.uj�c4�a���?v�F/a�8'���8g�+�Ϭ>� ��q����;I�{p���u;W�n�[;����:T�]L�I*ͬ��]��,VL�5d&���@��P��=a�aKU�����B$�7����<��Y���q����wL�8���ټ�th���M�P7 P�S�U=� 0�Q4!�Jk�r2T� x�������@�O�d=|�_3�8p��8Q��g�^';V�M �`�(iR0(��� 2{�y��ʫ�V��U`�*�w>ɔ�J��[\��H�(-�0Æ��;�����iiV��E����
�̱P�fR����%qNiӣ�ܢ�e2��5QE�ڏs��8�"�
c��*�+��	YL8t�Ӱ�[j,KE�A��B�rǉG���"KiR�C�8����ĘaçN�yҹq11�TLV�R҅V��V��J�XU@�aW)G?r��JSM4���
��rcX�2��15�1-�\�3/a�x��ik/�-J,�sq�2p��)�Xr�f2�|>C��F��N!ʗ�x�+9��`�e� ��H��xh�Q�Ai����2�\�©>��X��2e�-��,�� !�����X����ؘx|>�x�*�y���<�̗�jH�se�qr��y����*�&9U��KpC�B���xbg-�;q�Ib�y�E9ʶƹ�\UX���e0��m��Zs">	Jxi��=�=������̄3��s�૙s3 y˸y�8��g��2�K�\�0�U8�����+y��
Ul��&9	ˌ|�9Z�儰ȁ���~s ���5�L�x�Lh�y����\�)����2����8�AJ6��2��H�)�`4�l$��*~�����oI��{3���9ෲf"�W��O�	��n�X�#�"��z�jY6�.Q�j��[!�UGE��m������0�#$0��R��ײ����Q�'*������v>�N�i���6f���ӆj�U{I+�qʝw7Ҡk��޽5�:��O�h�ڣٓsO���S57��ļ�_b���n�\����(�9��hq$����Xb�^bhG�\�N�y��=����8�����BdMB�z=���<A&*��7K���'z�o��<>��0$~�<=�`}��=����5�o��Mc�x�����FF�����ˎ��5�o��X:<�A�m�nmcf��Ý'7��7������pl�=�yw��#[+ݰ򇷩fl"x����Q��s;�5��oޟ�l�;��=���g��������;��7ᵢ�ur���aӄDB�>�P~yw�\�C:|�C�=&\<��ꁏ��͔O�I�ܜ�<]��ٟP�Gu�!m�!*��^_z��מ-���Tx~�u�׎�K�J��fг�8ą�a&-�	�9a�9�Y�����4����@|$��^jo���=��I1=��U��Lx�����y�{�&S��i�=ݝ��:R�ZA-T����6e욺��=u�Z2tcre!���!�sDj	���0'��(1(�=(�� �U���r�{f�&����+����}�e�t����EK���4n*���ٯ85l:�����m�٠l)�0	��!�𽿦�u�*+6���?�<�~���\�������ydD���8�y� ����j�F�UH^������U�E_	ƫ�^f6r��"�v��w��{E哘���R�����I�.���{i�\2�7��r ���A���v�����-���e\�uFB-x?r��n٘7�����{fAk��8��2χ��W?ewx�h��Ӳe�l��;�\������g��lGrv��4>��}��1#����I�x;���;<M�}���^s>�:�9#&�гVzp�'�8�uo��(�1���_�=�==���<���;
h�خ�l���I��_.Ů�j�ܾ����&9�hVC}���65��8�ͨm�J��|,�S��Q������.ίFv�>���^D׮�Ylv�����v�#�����hӟ@j�ǃ�W��b,�U�+%��]ft���Aɷ�O������K������o�%z��:6�ji��ea�1M��ӷ���S�0*�X>��ŏ���6�z������;�ǀ���� s3��@�T~�R��IC��]��s���[��׼�vD���z���2Ts�/�D��mk�#���!j]7׹����������~2���?5�G�E��<�x)���(3A�etO^$�9�=�S=�E����ޛ^��S�r��̚(�D:�w�*La���;��Cn#���{o���T��zܸ�Kq��6A�L��^��*�y�<%Y�oO8s;k��,~~����okC4���x��7~����y%0����ep��8n���wq�K�yP���<��"ov,vh �%{�b@�X=�
�����O��7���8{�va/��a}���������&�&M�;��YF'�?7I�����M���/d/tĎ���v��4�{��Q����=�*�)�3"�ܒ�Km��P��ic�o�,olQ�#����������<�||k�l%�^�Xd>s�6n��'s×��Y���m�Pc�K�9��b~��w������S<����i�}q���.����^��b���ft-�}�:8��8dЃ�>9wB����3����\�³=���{�4o���p}m�l�rO3��q4j�W��r���x���M�q���$MC��}2�F^���I�s����	��LoA��`.>J%<��_X�H��>*�Ӿ��c=�E�������YM��8�=���Et�|ת`��k)ء�xy_���<&M���.��,����Ѥ�=r�P�3�;��������P�t<���2�{�_��ܸ��W;s_�x����U�'���w�7 ���0aޯPsɗ�5�{�r˜����b�2y��K�n����zM߯����
{8T�P|)��tp��Mugn5p�B}Ip`e�[\�%y�1½W�式gE}�ۺ^g؝v뺭�Yi��I�F+š&3*v��lo��OVF��|Ƌ��{M�B���S5jϔqvnO)v�&�H�����;q�F0�
��;�ѽ����[c"GM*t���s�b��X���5,�ͤ$�c���Şq�yB���F	Q���K畝�
L�@���`�~n�C�	�V���{9}J��Ӏ\c`}�͛�~�[��/:�u�G,�`�ć`wF�t��=�w�7����q��&�.�~�;�VL��f!���LC�+�e��x�_W�g��m'N���g.��<"{�h�{Fu�3�(����#3j��ޝ\����Ɉ�Ώ�Q/!~Kf��u�=����~�F��R��T{��o�砿Z��n���Ll��9ZI�fMAܪ��1�LȪ�R���L����<�w;/�xm�m���rW���$Ե�a\gvӓ�Y�a���3���3�� =�F����kv-���f�h�8�ts�������3����T�2�ĳa�_���Oީ�\О����,�r����3�ɖ��
N՟�<:��c��?o�7�w���� z��Ee�z��P��L��)�g�J?n hk�pmtC�{tp���j��jT�Y��x1�����)�<�ģ�d��ڿ~����k�<��å�ms�\���PWY�:�%��g=�d���^@y�h΢�2fg�7Ͻ���ޟr2�%}��ϙ����/=���վpp�I�p��+S��.�U�SwP��_1'�͋���}0'랇����^������-/��z�m��[^��>5�'�y�B����,��8��yAU;;=)��N[B�wy쎌8 ٴ��P���B��;���#�}'���h�'s;��.���H��W{�n<σ�Rؠ�B�mt�W�]%z�������e�QL�J�a�r�9��xO�az�1��i�S����[�^�2k� �{���@��"w������p��� v��X_��K^�Y}ۅ���sG�{�pjC�4�.��>� H=��+(�˵��փ�����/V�݄��;xt@����ble�$]�'�b����4)^�zƮ�dz�]i�}�d����O�(������H5ާޚ���U��Yǲ����5�{����a��켣z�}��㨷x�lvڏM���e�%ͽ���/\��{�qK�
�Ur�1����ݼ#��/:-���>�2i��h���k�a���%b�@�}��K���qӨ�2v��oM�S^��L~_y����wL�z���5��]nݙ����uq��/ïF����ܚx�˽�NV�c�vd���֯�Է@

^ɇy���ӯM��5�)�ƨ>��+��DMS^I�^�[q��]<��>�H��AT{����J���g'�ly��]K{Ջ&]��U��SW�4Pz`���Z"���OCy�/;�/��t���YW�M�e�Q��(l����`��|�cǭy�O.o������k�d";�\�2]E���̍�<2���kh{z7����ݺ��T�eݙ��{�i���$��974g�*�ם�m���X!!�a�u~�^�ۻ�9���h����Dy��/v�#���[�� �e�Mݭ�u�b~5�uK8D~�
�~����r�c��h��b�z�g+)7�ᗞsk�����`W���rLm��n�Mzl|n�(�>�m�z�HV&��uR(f�{Z �l<XN�E���g�dɃ��B-<�݌��]c��r�V���{�1����e�W�ux������<^E��A�c��m�Ds���oTW�m1a�xj�s���L堢�Zd �uq��w��q�%�\ب�i�kl |;��s��/{&�[��q������Ƕc'�믭�*�'���*=3xx<�d�q�Й��r�q�`f\x�!����������T�2`��3�t��t'�y����I�ߧ�$K�_v'��^"p�l�w�N���'��3g���{M>M�7"�vV3�f]9���-9���dD��X�)��5�d��=�=wz��ՙ,'�Ɏ{ؿ�na�hb_6c�@lD���j���Mx��Ռ���^֒�a���IC�Ӎ�N"ǺϠ�<��T������{Y�|��>�r����������Wi]�u���ko�o������~�������.t=��	��b<��:wCO���i�~n�·ۉ�����Br�If�>a��~��q���3�n�W����7(>���y%�7�9��L���)�\�ӱ:�̓��_���HW�I?�uk�,ޙ�oOB����ݻ{p��9��� M�h,�2>/�Y̦>�0�����Ͼ!�}�hѥ�9�z��l9�2�A�AR~I��jFD&F��kWh�Ⱦ ��2�;W�]zf��p�}��񢺺�r�v|Бqc�J��g2���C��}��q=3�ss7<������j�{r�Sq�I{��Ļ�
Fw�}��z*?=��M�����CtS��u��j�����j}�>h��͡ �z�2oI�vn��� r����S�H)��	*^t�O�{��B�f�=��{*\�Q��!�d���n�z�p;��/�48ez;7�M��2�Lxsz3�~�bWvQ�U{�{�u�wzipTr[j{����w��Gr��W�%���]���U��*���OI�����
�"6�n�$��L��s;,��VK�4v ]Í<�;��u�TA!pyC��E�~�o��<k;<n竏kNmS�$��΢4I�K��ŧ?{��~�7���~V~��Q������f��fԙ�79R��&�N��k%�A$����p��کz��{��#�C�Ί\o���`�2�s��	܈�/9�^��g����w���'�.�x��C+V^�'��כh�ґV�Fmg��N���棐l���D]y��,��-Z�g�eU}�a��>���.�4xzl7� ɗ6�Pc~�Vgq�nԾ�6��W���(1K���y������{疒k'���DcƓ~m� ��ڇ=���� Xc�Ey��3WyO{EN�v0�o����V���S�Λ=�{;�cT��հv΀��n^<D�A���}�0P=m�Ny4E㙳�3�7�zH<�x=tDT���y{���g�w�EI�]1����`���H�����I�a�VnyE����s��vͪ9	�`�W�=�;4���d��K�~dl��p���=le��������
k]����:#�9\)z��1-�����8J�}/�W�
s,�n����ϓ�3�/�L�h�lPbR�V�,y_f<�_E�g׫~w3`�"!p�h�L��l���wٟ=/�tG�(tc�}���s\�x�(g�ڷ`�r�m���*6&d�\�9�0�,�u�֝��{��;�62U�i��8=�Ϯ 4}��i��&Ji[.���Y�{q�VzZA]�Z�_Y��k�O*��r�'�f:1]$=*�ӆm�jgv���,�s�'~׋`�7p�A.��?e|��8����:�[77'iK'�S̽þB{��v������W���*6�k����Mot��^c��§��U)NI�����v�=q����7�=;���|�q_�#=��^����N��Ux��I�g���0����U�	Pt��SH��w��vYaح���]-�\����V�Q��<Ae�*�H��b��y���C�ۖ����8��);W�����6X9���v�®l�o:�y�)��z{����5<����$�O9�4�ӵխC�䷸➨����9�IM��g���)�F�nUl�����]y���WY`g.nI�����E���(��/��!>޷�4s�K#��UC�G�Fv�Y�;.Sg�k�[IS.��[W"�.���g�,5�Z�Y�p��Y��#YS��dǧ��pm�,�=�xg2�tAl����7a}�6���`����|���̷��L��:�Ӽ[�����{n��t�?@R���v�O<���x���)��]�6�qV��"n���[HqOO0�G0dv/X�m�P���p�u%�\�雸)9�X`d�lG�Uc@�!��`�fZ9T������]P���!��2^|��=�}˟\FzN�q����]�۽Y��j*�r�}��۝����k;�:��s;_��Y,��ʟ&�DMT���0Y�!``�˗FR�t�U���Def��s��C=-�N�J��s�����@п�X�<���V&�𒮑�jbO�9�tǖ��Z�`����\�؀Ĉ�oٹ���Zl7C����CY��[cbO�ɀأ�=|�~���6d���4]ɍQ/^�N�4L�V�h�ك{d�L��*.�ԥ`G\6+�jG�۝��Y��E[�t�!��{���.�}0��Q�:��	����+q�v�M����>��9�����zg���9��g-�@��g��v'�>�q�f�=Ҏ�gzI$���:D:��ٰb㗞���\Wu��}~~�b���
ll7h�q�̲g���x߯t����ܺɥ�ڶ-]|��5x����p}(>�o��㧪��١�����0Е���o��X
��V>0�je�1k����ܬ�Q�4���V��bf'��8w��=�� �n����y��ۙS7�����"Tz(�LՔbd�R�,���M��y:��sP.�;���j��}z�b�iR��m�t׌L��<6�T'fF�-���=���Jd'�}�ni���wG:fڤ�z.G-�R�]�H����\:#��D�M�e����%�cU�p�5�?03���b�)���f(s���#.��X�)[�Y�y��+�E�����YyJp�N�=;��LA��"���y��ĹKiT\�Z�fP--J[QV�a��Xc0�/1(���p����<�2����\�n[��/
��J[r��dr�%���RpqYArږ�j�^8�8t�ӳ�}q1z�Pǈ�PYYR�W臉�<����f"����R���
�U���R�_CR&4ӧN�֯Z(.0�T��-l�e�L�32�mjT�1EQ��P��b6�f8t���²Q�lmc�&d����0b!�[*2��\Lq�3.(�`�eJa���ӫ�;���a�̫e���@����jZ�j�Q�J���kF���M:y�J�Km��r�"V�c��)̥Em1�m)`��,��a[^HX�҅QlZ�&�i��}��s�S�
��J�X�B��,O9F3XQʈ��(5
x�Q��������[E(��Kib�mmKU��ETƣ�@5D�I����<3�4��i���>ќ7o����IH\K���#M�-�M��hѫQW�&xw	�ݱMl���� �e��gm�ʉ���^ӕ�h3��=T.�>�,{�*��OM5��Έ��Z��==�
�a�p���H\sL=�O�V�,�ͱm f�S7���VPB��E��|��Х�	���I��Uc�0=4���5��(M1����G���"�@<�3e��ƀ�����U��I��V����/�f�:H�N���7�0��G?�s�j��o�`9\�W�o)��ݒ����SB��cgc����!��;��/~������ޭ�[�� �'�"X[�$:���݊�Ó�e�n6c.�u�� ���8��z~�J}L�M]����Ξ}L��x�`d����'���h�ƳE3iv��@Bw$���`��{O��Jt��a�	M�k�vO5ȸu��oN��l��#�+�m=qHp.-�r��W�%�)�$oQ�%���NVy%msoY�������z�b������=���0�a`��OB9��84���^��yL4�P���`}>��n��]m-�h���W��G�����>�XEz0��b~#����F��Z�=ݣ�W5ُ"�G����	�e
�D�MUU�{]ƍ3umU�%+��ze����+|�d�y�o�bO�/&����GYSk�pUxzv�O�,�wS����6��7)�[�����%�-zLN�M%d��ku˂A��8��pvV������u�Z�7�R��r=�� fn]��2F�-����>;���R,�Y|�=^���z��k�R)�{�{�HLr��i��w�4]Z�1�y���,)��ϣƦF7��c�l���G�y�;k��+�NJ[y���G=::�Aƈ>Io��{az|@��JǱǧշ�I�sI}��:�3;u��4?0��%�'!(帇E�\�2�=7'�v`�&��CK�u$�ߙ����b�/a9�M��È��m�ʟ���,�
e�-��v���g�X� ��J�m����Bk��v�g�Ť��c)��b�f�*�tk� m�'����I��A��Y�|����g-{?�|����߆_�߀�<)��_��9q��g�r������5�K"���I1��d#ql�ت�����m{zWfմR���1�7Z$8@��ɒ����9a�6-�lo:y��,'�!'�Y���1�>�,�;�[���4i�O�[z��	����qw�H��z���z�9p2	�%�M]��]�����G;_F6�;R��1�yE'V�H�}<@�~�f�m|�����I��VA���y'd[|�h:�׻�^+z��uuDˈ8o����6棉f�n��yx3NxjA�{/� ��>`{���M��
vw�����v�Iا^y)��o��;v�B�lp�J�Φ@���:�7�c�{֣xi�NΎ�>|P�	��(9��� O_v�Y{�a�������!	� \)S�{��v���[��!2O`�J"��FU��Q�[�fr�jٮ����G-�oH�ƸO�9�l�j�!�LG�y�*,������p���垾��kL>� m׳���\taz�F;�	܁���B~�s�d	e@v�3=�����5�;q����d�yCvm�:,�ϸ��W��*��~+�+?>�mx7s�B~�*�,�"n�;��;H�ک0��+D�ۄ���%�v!����#ې��>6��{��-�B^���ۜ4�h.��Rurn��d�w�QaK:y�X�Z�5��[9��Ƹ`�p=u��y3'f��a�W�q��
� (�c.�@�ˍm��@Z�u�е��A/mbTv<�����.��E��z��gr�|���>/+���M�ϐP ���&�O�h����e�X���,k���n)$4�y۫��9�'o[-P3�{�L�`�<��<{�Sx���vo$��O<
-�r��z���m��7lu/��?�l��Ƈ@��o�y
�4	��_!�)�EE�$��kc2��x��c�
@�%b?(:��H�Y�\�J\�k�쑗?g�?a�tr�?8��ʬùQ7��;	ll2=������^i���Y���Z���m�fg�'ݪ7��Lz7�*r�G^�jf�u�GYe� ������C�^��H��O���U�M�1�����`Je��H�u�n�f�nk-ny2]	{/MVP�j͊A�-^�9��Dϛn6�7���tS?I�U�zR�����J4+`�L	����Uձ�L(6x��6eK2��Ty�}�4�VqY����s쫇(�O���G�3��"zp�7�8^��nj�"Se�/Ƃe� ,T)�k5{�݄F0�W1ʜ�L��^������F�WƬ��q�S�O�逐���!�݊y���BS�*�,��^Er�1�ٶ���K��MP��v#'2�U��������|[X���S �Aƀ�Sf[;��K,-,�����u�es�/Ɂe��Li/L)�/�S��'�k�D��>�L�y��UO�w���Wpm.�sH�W�]�0�gE�L,��.�s�7�-�)��@�R�"SJ����Mo�ie� e��;z��qf,��km	���v(w��(qUeWC�����⠴��0�ԜK�����]�xT�S��sa8�\ Ä�h/�&'t�`[p�:�f^��	uWF��w���,>��m�Yw�&���4�R�,�u.T�#]ٴ.�z��͏C�����l3:}W6��j�Ә�A�LOu<�Y���w�V?��e�&��zijYL���xB�Vz$�ͅ{�me�y{�o��RXU�/��b�p[�7#���@
�&�O�N��+����H+��{H�0�3�9�mW��3�8��Z��i��es�e�����JS���?��n�v�W�ô�(S�X?��?�Q�	:_ڦu~���v}��#yU)nnC�\�4��6= L�q�q�sO��v�K�gc� 3?��!�^�ay����-#M�f>�`J���;����I/�Ǥ�@�	��a���`��y�ސr�M����7���Jq;��6���y��ǀ���ps@3�a;Јz�" "@���kh��TEC�E��O��7gV�z�^�u�BSSP��������|�p?����w~�y���a�
�Pɇ�+�6Z3�s;��m��3�н\�'�xi���&���&���s~��O=����J��� �i���&�|�{�k��T�~t�Q`?�y��M<!�������"�"��Ԫ��Q�?�*�_3�#jۇ�}7�ɫ����x���)�&�,SI�]:��տ�[ռ�o��'��L2�"!��1����hi+zN�ٓ(`^Rkŋ��BxeμR�d�ģ)��F��`�3��?��A]���~�i���iw{#ƚ���l1y���D��H��,Oh&fpμ���e�A��;~I�ř�>O���kz�Yhˮ6 ��{�s����a*��K���Ja�rxQV��pEG������/^�]m�<�Q6��)I׽L=R8+����ս5�`齓���?4�WY8�;hz^�����!���Wy�ts�f��u/��Juat�L�#I��Gd�S�\:uU��X�v�ge���ޝB��ơ7R�9���ݒ��7��.�E',3�<���3�w�hK�6(������t��N�ώ��!�<#�D&��Ǹ6Ϸ'���Q��&�C�zV#��;I�S�舲Ҷ�̗����E:��s��h��/B���ǌ��?B�es���:�\޻���#�f�������{����}�J�_[��1.�Q��k]���z�W�uw�dd-	k��7����܄r�k�wk��1l��z���O�0s�7OAt{�&S���1M�/���kr����]��8�Y�2X��5�=����pd��K�om
�62�6�K�NA|/o/+�w{��h\��		�L�S��>M�#hgRN���0�-���sx�
r��l��~@���YW�8g
�A�/	xd�>(��?�ؽq�?}C6�Z�v\f��,Ŏ����ץ�'y9��ðo}M�σ�4��->�W��^�������X�t��K9�uG6W��%�}���o$w,.�:\w������1)l챽V;Et���VO�5�dc�ܯ<������Q���gNa���,�r�h��ɻX{^����m��8I�D�^�5]�uB��rg5,<$� <%�)�wu�s�&�վ����_v�wUsTK/�*~*6B0��5!�a��[��D�]��[��8�5q2�����@�P�),A�_�5n������u�ҝ��"E�3��l�B�������^(�3׳f�P�1�<����8.t%N��D��Oy���F��
g�-�y�<�'�Gc�'�P%�x��g�c��@eEÛp�Tf?m.��+��=�!�㐘�`�y�Y5�\��tc���-R%TX
e����lv���r�>}�d��>��
p>?�E��Nې���*��D&I��J~��k2���%*s��oq��5v�q�A�`���	���!F4C�.�L$�v�۝�7�Rewg����;�F�6t�l�C��(�x�:,���ND��@`�|�L���S��,�If�;�*�l���NZ��8��m�,�/�F.i@��~�����p��t��C��υ*t�4r�޻���}\CF�!�G@w[/��Hu�{��0��WH薳�+^���%�a!<9ՔhWʝ�q����Y���{a�z��)��K�~�^�(���|U�:���*�	�_�ƃ��E�$�YȌ�U�0�h����4�l�ӜpF'e�����-�G��'iA������|��D�j�-L\bHtg�}����0k>
ِ�{8
���9�QɺU���Ϸ�ʹ�����l6P'�s&\j�.Q��d�n�P���9;8����Uy�(B�Hig��oe0rŧ�!O2�06�b�l	�8�1�\�T���R�`$
]?rb����2/aߧ���#��t69�6'0���$����	8q�B�w+q�)��ʲ��G_i���<����{�D���`����	7V��d��W�l�n�Ƨ�YT��b�<Mm�etn�T� z$�ݏ\fb��:#�Ʈ��?~����<�,"�L�m�d�����P���!�U������P #�t=2Ή��,+�������[F�ʬ���}�#�<�z:�Ǟ�������H<�x� _�Y:
My��i�WL[e�N.1ӫgG^g�9��Gп��v܄vŚ�T��\ʖ���B���� ʖe
6��y��&���������}l��|�dS9�9��C��~{V�eӵ-�C���<��q� &��,^S�~b�%[_ig���_	�ڰM�t�T1QY����<��N$���,ht���Xc�d;���ik1w�ۭïA�5�Xs+^��6B�B�6s�ϸ��V��y-�%��:���5c)1�+�e�<;���1�Z�8f���[�k[�1�$��0��y5��Mԥn�ff�E0���������T)��$�OҌYU5)�>��+��X{8o��:c��V�Q���jM.sُS�FEt']��U����NU�VXkF������c��6�������MI�ȳ�"�7E1��&���,c�P��Ǚ9�����U҆��~l�|8��BhAhv��`h^Jw�}]0�U(���Ƃިn�`Ϻܷ�;��h���vt�W�+�l��D�6�D&�&ot��vcb��*��s�����X�������1������:R7��/��u= =��Ͷ����xO���ɮ	�~�ì~a�iK�:3N�S�֟�7h��u�@���ǋ�`���0��8u��*^[{j�[,h�0�3�-Ř�ȝ���yx����R�
��
��?��;!t��!��S�GW���RO���}�t�u0��=���:�x�,�I�O�ٮw�ϧ_Ն9�L3�gb\j��h�_8i��CY�v]m���6�]�����{(����H��Kώ�1n��dtK�H��eb̌fC��9zb���\�ӎ0)�YoX�G6e�{6��4�A.�� ��p�u�:8�=��ܼ����k}%W�ײ�Uĳ���-�1�`��I�^��F�hkNnu3M�K�V�A�&�*�}%�)�r7{k|���oܶ�p����r�]ε��.�'O!%�em�N�"��"�2�ޱ�<�VP`��s,�.W���A�Lβ��{}�b������bʎ`X����HS��l�yn+��d�=!��#r�v�� TU���m߷�ÇC�sE<5�P�/��4k��|~4��,��|�q����S6BC'Ae���l�9r�j@�T=S�Y��W>s��LM���,:.��{ְ	F�B�i3UGw���X��>B�	-����ҟR{U����x��Z~T�K��|��08E�0ó��v[��$Zs��Py�^HC"73gA8C�K"�R�er��Zof��֡�l��ߩ�ۙ<�ʪ4�~�5������7T�`{(2;d��DJ,����z^ΑLR2����}̡<���oou�T���y��D#>fژ�˲���0�w�ג|��`�F�;U#^�Y��r�[I�Ց�eW�G�P�W����������`���}�)����Z���2����C�EbY7�Wv���E�8J)qy�zX`=:�D�2�|����_��U������} b�Z��T;���5��rֵ���X�B�ce����9 ~��J#�_�r����p�L���[,��}#!�	��U�l�])?5�2m��ү	
�E�ӻ6�����h�� {��(����WC������']
g4�z�C����J�}a�ɫV���E\��T��K�Nzc��y0���OD[��Z���Y��㘃[5bK���v���oE`�(�[��)�淼�h�	���y�5=�_S0w��[��Qo��'��Pb��k7�M�E�"�)7����+T�r�������K�zCJ�=��V��3������E�7�n4#{�>�&���v�2���/U��\t�Ε�eA�y�a]�k�����C��t�OqdP��:��띩es�F3��'���s��܍�U)��^��ߘV�;1��_vՕ7�kkR��[�]���0��JvMf�B:YW���CUp��!�б�J�yrH]%^{�7����ˇ��|s��Z��Y�I��}8�>��Pl��+9ǟ��-�wdǢw_g	����}/ u0ug-�m��y?H��`eR����B����AA���8���g�)�ݶ�ɰ�TG�WxƝR1��n��m"�1s�	��_��^�a�f6�g<���>�L'�>+΢ݛ��5!]Ye��{H�*��N�\֍�G����9�����;�9�J2Xg�����7ZZ�OYb�*�o��u4�D��*��׊-v�r��z�r��`ky��7�ñR3�#[a	M`X��gZ�3)P�F�-Y��[;�|C���DM2"L|�(z���QŒ�I�V��������];����fX�{`YO�c���Tn�����=H��2���X�ʾ2t��A�]LGvK�@����K�7h�G�h �|"9�{��6s6q�i�c�Ϡ�$ۜK�t����{��f�N�����lz`�;��P�_���v9.,:�.��MV��sV����f��T��0q�p�>�k���؆�����q�d���]�3��B�<&C6�m-�-��Lu_D�t2��(Z�`��pe�<��>�>٤p�%ܞ;��}��Y���-,o]�	��tu�r:۾y�mۊ����Y���D�0�5�$8M�?���{j7�Y�Ɍ����XO5�m�R��V��g�����Sut�iQ&5�/![#5�i�e2��]%0��ӣc�>�<I�M��Q�_
;�p{-�#X����>���٩����?�gm��_`�� _�9� �5���w�1oua�/e�����Tl��ٛ���d�L�=F��(NGAѝ8�[H2賀�Z���c�(�M��e�-��h)����_�4xh�e�4���N_S`�l]�t����X��B����+�G��6bn���<��"%;]dv�ܷ��q��ED8s�]
�E�O���d�ەϝ��Ә(���6V�}�)7z��¡�%<�W���������a���~%�� �I��D���
�!A�ZY! �^���2�x,H�	 >O�0, ���!m ��
U2�T�eU�����mQF4IE֘5-����?Y�� ��X�X�(������²�Rؖ��ѩL>��<N�Z��*։mTM��X��Tb��1�RV�Z�-mV��J�
�>X\eEcl�c�)���N��(��J�Dm%W���m��Q`�����Z��CS@�+R?�����T���8zt����h�iU�����FVTX[,Q�-d�/mee�̷�"�[k*��:t�ؠ/m"�
�T-��l�Ԋ�l�֥J0+�(#S�ž��إ0�����X�E�J��"��\J��Uk�oR�6��*�DV�VS�N�:vu�[*�-B��J�h-A�%���,����G��&R��0���ӧT�Ti`��[�9�+��E-�Z�e�2ȑ�[~ R���i�N�+��QUE�rU�KV2��1Ubϗ\�T���X*`���`Ĭ(�l`י*-Lq�
�Ee/Sq-iF��P�	�A	5����j�ʹβ=Dg,<��F��%�m�����`��Z��j��4���1w�M�$2ܦY��ƶ�Ҥbe�
�I-� l���e�X�{{��ș�����;c�<3�p��ĖLl2�j׾=,Vߤ�7������lr��q�5:���j}L��
[�D?�X΋�f�Ѝ�4��~df�w�g{�+����C�k�6�E5��5�|7)��=�q���Y�r�%�9����f�}y��Bk��vML@����r��[����,��C����,����D�� ��o��IՉ�[e9��yg$C�Jw)e9!�{��L�v�����CH�ִ��OȤ�y@|V���%��A�D�3�:��'���<�QԽ���Ɛv
:�n+$�(ų�l�,qL�������P1gEM�V�Y������]~��&nF�ǚl]'��|='�f@�4WQ�rz�?�0�߽��n~,yҧ�悖���'��t�X��S��>];.�%��{�c�(����	�+���k\W;�/ޙ�ܽ�u����O�~���X.|2Do��)@L$���u�mn�&I�g��'S6�,��c[oW���:ք���b�8��6�k�[�A|k��g�,5@��G����F~�����K�ى̇�4�I��-�m�2l�uM�6��\|�{�{�Iʺ[M�����nb�޻8=��tx����n���!�P0^�f�5�n՞z�+²y����߻�s�j8|3���>�.|�Q�=�ys:�� ��4%��лw�6�@���%ˡ���Ʊ:�'���78^���N��F3�	� L�b9�s��t�:������CbMCH��FYOt����Ӌ�F�er��q\�+/��ھ������|鸞��Q|5Ph�R�`A5�$�=I�Y��n���ƽ���
V"a�k��P�{�"79n�p��i��� s"�%�\�ՌL�c�䧘^ƷT����[^���l�Kk����ӇR�8��,��D	�	�����B����:���S��˪��K��t�u�541˖W�:u�V�XhJj�;���p�38AƷ4�|Nk��&��j�J�v�Q���+�ֶ~�����G?-?�K5�g퇍s�^V
��iP<�z�? ��s�a�k����Q�.嫧�Rl7�#�;jX�0��_I�nǮ30���4: �r��y~�Px:#��S�T���6dq,r9e<�B*�.�U�'��	E@A�KF��Y��loJ�]K-D�`�tbƋH7?��.&$Xƥς_5�^�>�6��r9ʸ/"_ء�?�}�6��Y]���9���([�'�N��gՊ}��ZÉ�g��!�7��5�3N`�f�}�r۵��Y���?t�3�CfZ����M�r�3�j��L.�S�������Ƿ��Ϋ�qz݄g����K�]6�)9^,-��|������(,F<����������b���"Ô���K�TcWX��kj��!k��A�,�L޼F�/�Ho� ]�:�'�Oݤ�بgݗ�^��E?��?��,�Y��P���&��A�ƭ躹j��^Jչ5�������Qfhxs�?y	�(ǘۜ}���c����p��)KϠ�p�kux�����&�ɨJ*������з�x[At��w�u��'ou}�u$�D����)�s��gH���Y'X�Ƽ��¼�}��L'�}g��o�-F*�`�+G&kQ�u�N!��D��]��酎H]9u��Lkغ���K��f[�����n�j0�:�A�Z��G����M݆D���ě*���~nAbw;=��_(�VF�lf�SY�]����aQ�m� G�ꘒ�T��a;B�:*V�<����FP��qh"�sh*�O�cP�	�p��� ��� \9�i���u�F�{LWK������Վ1k�P�碠���ԤO5yMK6�E�]?t��>����@�����y��~��v�ӊ���kr�%�s%X���6M1C8v�X{��y��nY��N���E�.�Z����.�g徱��E�����g�>�p�tA����X6��3�I^;��N���;�^�n�yJblj����j�1���v��f�_��ʙG&g��v�WRb��，>lz��T��s;���j�1����
,���C�?'�.��F���n�nJNl2�Iz��ߒ���-�Q���*!�;�k�*���=%i ��������K�X��%{��f�0���$= js����o�d�����1Y���Y-��E?������Z �O��i��Xw�@K �������Dߢ�P�Y�T�s'��_k�[+���(#�a�Ƚ��͗�xi�x �
t��#ciՊ��
1cj-���f,a0aC�i�E���3j&Hd�D��R�C:o�����)�j�=bz���f}���Ƥ E5�f����L3T��H�D���MV��{
�a�V��O�E�I���d#`��Ї�	�Q���(.aN�x:sdp��E��N(r�d^ʀ��\�I��m�s�:{
�\��M-��ǹ�n�G@�2$�6P��
{z��X��^�b'�'��N�@�=�&����� �D2S;6����]����u���-��T����R;%�.�0�7��O�"������^�&vt=V`]�X�OKʼ~_�Z��:ob��c�����{k}�|�rS��/���Gfy��U��b���5*G�`�8]<��=��P���Wf��/z�s��4Z�bk6O^nv��d���t��*Pٓ�����!��8.1�NR���DDb ��{f{V�P����h�m���I�2j=tE����{aH!�"mzc�l�����Ss3q�Ll�=5��y���5��ɔ?�=��ϞA/^����,0���3����,P��!?�ھ��/��ɴʪ�,C�-�R�ic(%}�q��>���3Ғ3��C`�<������EŮ۵�F��� �]�O�$Ȧ.L�VoJO�kl8�����0(t���wB�束�����KMn�Y0!��C�:/R�7VIa�������LsH��4z�Y��UN�s �K�����D`��Bd�͉�]��E�C:�pB1,8���ݴtA��۞�ћl�"��X�ؼ-i�A!|�O��3�0h�َ?�y�~���.S7=Bs�w0'��M�����Do�49=�M��ߕj���l&>CG�\sLL$��ŶS�9bQ���kOs_	��a���t&�J�b���}���ˋ���$�1'���Mr K(�f�ݭΈ��uUs��άk㲐qx�7`~l�b����"�:�a_?T���lkʂ|ҞJ���쇝W���`���{ءeL����̷W��s�Ub�+Ɖ �|s3��|�g���@���g�N�U������w��k�d�'���w�=�����پ d.eO��s�U=7w&�G2��c���_C����35��tr�Q�a_�'�>��0�L��ǚl����㰂z�K�m�Lu�7D����W=^��ϖϭ�~�����!��9�������箈A����Rt�H�桋���u~��A���3���a��~�[^��| z��Rd]	���r]�Od��tBd���_`�KY�{w.�g��l�{K�P�����$vD�J�t�z$ƟC�H�!�m˷p�(�5��f���g��ᇃ��(dr�s/1W�y^��@؎�.͔����B1�>�!?Wax��1]126��H]pq��Cj-�t	e]����y�q�d]axع�iȝ~w�~yp�Ӻ�3�fqc@�g�[�y\TK6�	u����炇�u*l�¨Y��G.Rz����#�CRyw�*3(���J󤊝t�Ӈ��-�"n/��Ψ]B͇6(���Ra���hҭa�W�j��o?Z�?�/9���FP�i�u��C�� ��C�-��`kd��@Z�u�[���Br�:�yvg5tw5�8��5��Bi�ܬ%܁8?į����L-�}B2w/g��ґ��r?�
�w�x<�%}�Ar��;���~G���W'��o�=9;ُ����fv�I��xj/u�<���XI�l�0Y�#H~���y�ϯ����4-rw_r�����փyU�@�fw*3������������n�����|@C=��h+o72��χ��?�`�"�C35Xyd(N�}(���=�q�i�����
��+zz�<�{��_ATV9�/~Jwjݫu�/}]��=\��=�.���k(��1%�f�zfa���9�#��<���!L�s��u1}m���vk{�G�����������dnH%���zA!�8A��,A�ʇD��B��K\�In䫉�6�2��r�dfN���{Ǧ�{1��0�yj�9��B��vwii����������ۀ��k�/\�Ú �3�u!�Xt�>dI|Q�����kj\�-s��!Yj�QM-;e�j�n��e�4��[ӌ&�*<�(��|��9)�A�A�A�<;���P�͛\\'Y0-^�J��סsj; T*�Į�c0GN����KU�3�t-�8��B`$!�n�l�SMb�[�����#%��pb-2��8��J`��R)�.�u�����1��ƾ�Y�!eu�N�[�L�v4$v*��L�����$�s�	D8��}:\[�L'�Et�ǇM5��ջ�o��W2���X"�%�n�c@���������E�xxs�1�b�v�4e ����U����C��Tå#*���X��c]��7qM��kE�$ �~�����ۃ��Kc�J1]�'U�!�j�H�1Ӻ�j��ۄ���wښ��{>�s�":�s�Ǯ�쾴7R�Aư&"�v�wy:1�q�7]u�Ǔ*��PF#H#"2�F@?>oߞ��xP��8�݃[�S_�t�sy����	��<}�JU��^��~m����R����q�ظ>_MT�yl��w�vh�a1�M�"8F�C�u�RX�a;Bƌ�D����}�k|e�fSK�����_��P��9�K��r�F�>���sO�&%�.��$Eķs����]̃�TŊ���z���������:�$.����c�a?���zo�C�Tu��K�/C��+L��+��eO�Ǣ�x�4��,Ľv8: fڻ���Sl���e�,=��4j��N�����<3S���7�K���Iz�"e��C����qn4���]�GkV�Nت%�,?0� ��LI�:#)�].��}�=Z�� �<A�1c��$_�Z-v��]�ec�kW��M��b*PȖt$!0���,�l���ލ����Ζi=�E�>TM���ռ҅]"�E~�O4�����CC�(�0/
U���?|t��ŷ���!���ٚ=\-����L�,d.�l��$1�,�d5�;A�fͧ�z���%�
l������}�^[��$�]-�7v�}wi�?BĿC�ʂx .m��[��b�U@�)�����*�z8t���3�$�y�@�(�_E/�edt�H��L����!`��2C��x�t�.g�j�o��z�ʌ�ζ+ΐ5+;�^�J+�M�	@xM��ڪ���/^s��^\���O� F �#�d��yϾw��??3�I$K� �ߥ��P7��
�_���|s� ɍ�4����z��z�������z�(
a��z�݅�*t2��a�ph'�!�;\�:!��"�Ji��Q������࠶�{0��;�8��[��#�d��vl���OcH#�>����>)Յ�)�4TS���efZ|=m]����u�?-2/X�@�<�+�;�$pu]R�dz��{��[�����[�z���Q�v�/"��n�G��|�>�h���Ȏ	��W������]���:��������c�[!�����<�b^�\^G#�<z�l�
5����5-���Tk�F[=��D���֥�QxYYK������:K��
!��kW�ȋ�fLG'���δ{�y�F.�	���C�uY��h(��*2m�T{L���n���S�kj�]M�.�*(33k��L Pr^a�?'�.��>�4-�ø1�e�~�������m��6��U�]k���4�B��0g9g��&->����̟0^��+:pB1,����,�;,��{J�����#|9�a؉9������X<�-r�~��q����Ȧ@�xy�������ifRsP�i(�+�� ��$�����3"S:�)w|dq%�E4WUJ/��z��f��w�&L��J���n����io���Hw.y���|�{���}������a�D��0�� ������ߟ�s����d+�j��n��_��xg�h�gh�D��6&6���;cmI������{zxN�9����A�~?|����Zz�xU�%��4\s<:N�K�Qk��ns�OUWhǴ����]�N2;�-��=sͼ��2^�4���]V�[:��X�;Á,�X��z��J��nc�-lXnj ���ϠfͲ��-�<��S��ɕx�|�o�/�<�Lܑ�P�xe�!O�t|l5'���]X�z�C�}T��潝���Ʊ�^��\pgh �a��ge	��eѬ�|2as���QIճZ��%cI؊���
�9�k`�2��\E��ɇ��������������0vJnou��1R��&���l�C��u:��D󢔊P���|�`��Ы�V����i���2Ş\k����QMO�0�]~.ku�?`�LC}�Th���ł���ג�@�E�����F��F1����C�P�2s��z�8!�p�C�D�cbqT4�꒞x�2.��xӋ��6��sӿ3��(x����%=�{b}�g,�d:\m��z��f���{8�Gw��h�J�V�,ڃ��D�)ɡ_S�Ieۅ���w�-f H�ˬ[�X�&���Њ�ۡX+�ȼ;��5�K��v�\��<&p�1w��HNdbvչO��&����M��ހ�p.7������h⶯_S"�a�c��l��F{O�3�
�{��_�%�"�{�]������D��39����\]�l��L�H�]�[�U$�>�7�P�V��;8?(o�8��N�����{q��}V��$X�H�ɲ��׽�z�����={Go���4��4ڛ��7T�����mE����B�@�K��sN�ص��L�����S%^�����&��3ɳ�A��|�5垴�������t��.�oY����ag��D��� ���\�܌``�Y��{�F�����5���A;�Z.���J�yWN	A��E�Xԇf���=e s�����2�RfH��^˲�~���nz.���=�;��l��r��N�_2X{�p/��R���ҩ� R�'���ݲ�~{��f�z#<�̓""7���h�ؘ�,P]&�Imt����gr�o��jk�gsk$�Ĩ�Ţký&ICU�yb�$�)�-M7�2�i���`3�n��Ų^��s��S^}e�@�Su���;��F�f�w3eV�5�\�ʡ9�Š��CB�C�N�ؖ�� csٞ�lBf�����@�I����z�s�����/w�H���[V���hd�-�\��P�V���U�v�|��A��7i����(�z*�ӹ�j�\��(4�]Y?��K����EԔ�Dƅ�l��1�ո��H]KTՏ�>���M�����:��r�ɥ:u�L6d)��fUe�U�K��l�U��fW��1���}�H;�o8_�c_��;龀�����|\�_?�̼��f)0��t1�6�)iq�BM�o��������
���;̬��U�ue�\�����yMw��^�����A*�����Y38ޔ)�l����C�b+6�0��ˬ�Z�膫x9�%˾�.�C#W����$T�������Q�IF�.-�	�ŻU��H��@cH�it2��q�'/1��-��s{	8�-O���<���
Z�+��1�G��-A< �7�9��ᛚ[�䵛�zoE�&͑�s>\u�||2�:����Z9��!��!��v�°T�^��\��ū�ٜK�O�O���^�a����=�i�VLͦ����8Ù�y/�>����y=�p�3@2�j�=�ul;�˥�D�c��W$����"%n��ջ5Uq�Aֵ0�`�o���nن��W�T�}��h��^�\Vψ�>��ޞ�=��jƤ#��:^.v���7c7$��"�ӏ���}�P��1(�B���<��LD��0�{h'-��f��ܕb�1T���g-2���M:tU�mX�K^ڙh�EDUYim�գh�bZ խ�kF6���
���
��Y�=4���l[N��d���y�V�z��fe�եE�iJ+E9n�5m���KJ������ӫ��օos0J�E5�es�r�AR������_��<��[[X�N8��kF�PeNZ��8t�N�Eb�D�F�4��EEEb �Т5��E*�(�֔2�ڕ-l%��AFإ-���N�;:*(��R�V+=�eE=f9[���K[Um��ֵX���e�U-�J6R�S<4�ӳ�h�X�U`ĭADU �
�Ue�i~Z��ҕ�-J
,UUQX��OOOON�<�,QEzYX �2���+�)iq��FAV���%��"�UX�R�T)�O�;��)QVV6�ĥ��	�,��J%�)k+Q`�6�-O�bQ)E\h��+���j�r�"��[e�-�J�V�JŬ�heV��j�ү-@OL��'���<�o�tK)���.V�g6��=�Ë����k��/�J�0�z�`Ju���m8*�[�_yi�̺��8c���7��B��""@	�b�'x����� ��C��=	yO��B���¨Y���w%'���X�9P�R�Ύ&����KM�w1|��F�Ӱb�[��7��ά�гnd�w�Q�
:y�)a�m�fs%�L�f�����R����A�p/������Bc^�� n�İ;��-9�&������i��� �^�������XK�0B���%xk�ϗ�ߙ?e�մo�O�_�o��*N3od]���wh�w����R�l2�{�ӕ�5-�^�/�Ɔ����D������f�j�Ä<4�)���i��̪^�ُ9^͗��[9E�qa^��nס�`k�e��tgO:���ZMV_�S�e��(Vj4jC�p�;�Ƞ���ٱV���ٽC�"� ��:�I�=O��|�1v�qm{�V�ڽn ;F�"���DfN��%���~�P��Õ}�|0^p�Q�𘙚u��߷���A��^Ǣb���*�?Ņ��O��W��<5�#4s��B׈�ܨ�q����,�M��Լ{(Q�Mp��l2�*�Țh�#ɭ�`�$?�^}�9���+n�Y�
���Wi��v�W�y�q�L�����t	өΕd�J��Y����qX�����d����lu�U'Tx�]hġ���Dc����F�U0iJ\�n��k���+PYX��R]�B���6���<�n>�<����~���!?D ��F@D� D$D� ;矿�-����խjo�O6_	�yb�I�J�w�Ӻ��*���xQ�
hZ�!^Yz�v{�3���1���ɛPz
���H���Є�%���R�&�EP�Ȼ|���mb2*tbw��?����un��ϩ�BJ/k�g�1��`}��G<�4'�פoL��<^%�u��Lh$i0nz�%tvp�pj�a��=7֢]'�
��0�%�n�Ɩ*���Ⱦ�.�X�R���b�^٧�g��2
�q���;r�B��f?B����h����C��	���o�iC��qWK����qC2l�Y�*������{A�{d+a2��a��8�x`>ϘG�̛M����/��x�����e.yQUsI��s1:g����uWJ�s��g�..<a?|�Ѝt�_r�z�-����w��͝t���.g���*���-~*	{��J9���Y��-�4`���p���sfx�٧u��q���^�j~i�f6��͛d�e1,��Te�>�~/ͧ�Y����,��t:��9��H��	�|)��P~�S�<�b�y9?^�/�Ǥ� v�!��8�(���ې�@��E��.�E�[b�;7���4��|p�F���y�k+1>��U���ް�%�E#g6{�-�9Y����t�?e�m�8$d���1�]F�^=d�Ͳ��e�B���g;d�w�Ye�z���f�����S�J�IB�M�����@�	�d #$��I ^w���������ؿ<?=u�+�dĻ��円���T�{��	^�)���r��}�Zry��Ƭ��sr�c�n�$/Y4�[A�z�<�Ȗx �-- !�ZD=�O6�s6�ֵ�}8
�}W{�Զ�x7grf��g�$�B�4�e������
���C����(M�i;�%D*��<�Q�ٯe���,���lo�;A�ٳi���P$�`Ḃ��t�MI�o��x}��:='&q�.�^��%6r�1������ޗ����嚌����K�{aދ�T��#K���<�.�P�U�^��O�)�ijBQ��"N�N7׍X�s�&���m;7��k�!�eb��+JC8��D���@;�~�I���'.�F��	F�6�
��;�b�{8�kk����2n\��= ����~�Hf�?���7�����j���k]�=	�S�vD���tE��Oyms0nj=]������G�B=������V�4�$�	�W�����O~�N���Zt�ü�-?$�	|X9�A��L��h��s_�%�q��QR
�;��x9Z1ݗݦ6�u�i�:��ʽ��H�'Da�n��3u��wp�To���n9��`˔�ɇ��'�ɘoiY�#3V�����B�;Ueu�V�ѳp�xm6�o�T�����ڂCj4�1��x��7d�?�~�$�� F�$�#!�$���|��~����8e?f\~����naڣZ������O���o<;����*�7:�Md�[#D�b�|�d���d�r��AG��}�f����˚֙$d^Z�E��ˇ�bcLJ��!��'|�'>@��?��$O/��Du�}�hZ/�s+Ys��x�7�)���ߏݣ�+ϰ�S��E���D ]��R��
�s�4[�7�#ۺP7��fV�k��%����-�V���%p��C��П�2�����|�S_b�z`c%[I��L�ۻ@�	��]ybUMO�h�W��bĿC�D]=c���"Oᡈg�-�	�Ǵ����uye�e��P�K�戈�}5n=!1��Sm�6}JF�A�n*q�jD�Pz�؞����B��c�l<1�*��fԘ�Da"-���)��W>�6m�d$R���Y$5g�G���#Tg�0�4��F���-��/N�c d����1��f�s�V�/ˤ��˟��j�KLh����� �7Ǿ��o?��]J���K�l\g(6"K����gV�k�D)|��;/j�L$�B¬$��Ku��:�E�	��V�&2�E/z����懦r��'P~g;|�P�ʫ�#\����FTr�k:���tm�(\���gr=!OR�:SFq՝֕���S����"�%
<
L����d5��l���E<C��D����~>�>@� ��0 #	�0a� f�Y�ܑ�-�h���q�JĪ,)��[`ꋇUq��"z@K�I�r�mO��̦p$3y������Q	��w��T-X�E8���H�m
�:q�0�H1�" �nj#�ma�֭wG2��� X��D~�F`ޯ��X�`HLT�	.��}��o��}ǆd�%(g��9\3U�h�m�������|�d	e�f��D��c��"���b摴vk�T�[�j�Z����*-�$��`�fy|^<�R<o8�_��У`�&B,�^Zv�'�suCkz.�����Â�˼6�Ga��u?3d��G�*��*?T������h���I�c���k��QP�.��f�n�l�����UԘHOt��9���>Ai�����y���cNO۞�f��|�[X��f��8�V-�y�Os�?��f����4�rp_���������V��~��њj�f{^��5��*
�oMc�wh��R�ǜQr���.^�BEH��Y�S�猬W�xl_�gx�*a;�uY����¸ė�L3v=30�tE���-����h�M9�w��������e���α�6�,<sU�ݜZG��0������o��T�����F�ř��ƥX�֜��,5{w�;�Ω��� �6V�:lE�UL�ot*4C�*����۲BU��_]G�&_|>����}B��	$ ��`@D �=�*.ҵ�ͫw�"�L؂^a�>0���˰�Ⱦy��(2A�Pdz"���Q�b��/l����n~����S�g��(`���ߐ��>�p��Q�|����v?W�
��;�?��_/�V����<���X{���o�xװTȽ��x����;�^WT��\ʆ��n�ý���Oݯ��߯�:����Y�(��%�>�)�״mJ~�
g [����A�*e'ih�SoJ��&�V�|�2٨	U,Z�)����BeAb�I�Wmq`�n�z���Ol�{m2�"�iT�<.��}��l<�1���:5��-�-]Jc~/)B�)��B*��d�>���zz81�����B�K�,�gN\N+wH8��}��`�Aƍd(�q����&�n�6��4�vN�|�v*�쬽�����=M�|5ips' o�}ʢ�=a�Uz����E9����R��81n�ܝ��}�[4*�W3��-pi�c���j�y4���l%��?�Tc�ݞ�{�>hB����~��Sgk�S�r�u����	�,WA����8�x=�C��e����G��*(����M.�5��d�è`7�2moߝ����ډUӋ���=�$��+�i2<�L��&kX���h�*�����U]F�f���<lЧ'Hn��d�c7�em���5r�����c%�!��M�.t��JN�M�������3
��i���{G���6t=C*�b�P��/�Ng�H�A�I@�� �HC�Ϟ}�<�����ƪ�!�&y�ր��Z[B�U(zY��!b�c�W���@Ý� �|����s{z��K>]b����9@LK$fSS#q�������R�lF�Yr��/�8��jC��j�w�o�{z����$9<�ͮYz�3vo+��\E��)6��L�q�`v��L3Z�[;��Z×�Ʒ�
7�	_��a?���jj�+��%����{��3�E��:��X�1
�j-s��^^�"��؇e>�x9!�<�s�~W�+���7�.͘P,����L��K��eDT^t�h"����n��W���Z-��mv�U���~�d&�{d���[���Z��s���dL�l��u3M�,:�YA\A���8��KL�����3������ʌ�;/�$�J�־,u��0�31��zdy*f�;(1��q�j(���6��=[¯t�wh/Z2�^�-�.��命4cX2� ��@���WY���4���W�q�)��J�҉O�WN0�x�^>�lz�t`�#o,z9�b{x.���,,-�"�l�+&�2�k�N(�d|���R����~O��.�my�k�tR��侭���i1�re�Ez���'���^���~ǲ���	o�N�;f-Z�}�#�v��!O�R뫰Ȋ���7��]Xv��%�����rn\M�.��s�O�Qdے�l��xn6c�����2� � ���	d���D$!�>����Ͽ�<��3��d��f�Y^_��V ����<����}cH"}�'�DJt�r�9�P�j�v{ecf�:��H�T�m66Gl��ȸ}��Ŷ�R��&nI�p�w�Biȭ���O�;S�ͭ�����E'+=�"�-�a�@�az|�>�E��,�gP�A͆��y���)`3*��l�ڜ5���i����Y��^���'�K��ZGR��L'Ǡ?KE�99���h��Y97c5\V�%��=p���iM7X�U�w�Qx�1m%�^�L#����:LK�@�j�R���v��vxTꆸp��1���P���P�M_>b��Vn���sb�&ެR�3�(�k���E�m���@���W����'�D���]�?4u|^�0!��pȥ�$��_Yc�7�N��8���0h�V�s_r��d�"�A�'�A��k ��qO凞L��kM�P�g�;r���r��잂�֍8(7)��^��q��K�G���Uh|Qc��տ[HMqӍ�̈`n>J�b�W0A�1��p��b�ėm&Y�H&:H:�qlS���I�fd��P��\�J';�N}�-�t�����5*�{=�E�}�Je����#���#�z�����Bv׷7Z��o�+�"��V�O��9#�ɫv�*��؇�_�I��E<�6�ה��G)ӥ���e,�@�uN��R]��a�6����O�?F @F�$ "@�2I`D�	|����~_��h���LQ";F6ӛ����	��<�^N2A0��ԟ=�6�Y��&��n͝�詴%�	�兽Ŷ���z{=�X��A��B�@�CQFq�Mg:j���^�Q7�Э�(�� k�N��d�Q��D7l{�&>/�T�7}'7�>S<��s�n�~j@�V3�1���쨸uB�38A@��ds��������R�������^��C��" b!�s�%�Z�R�J��ܜjꋇU�5��z��ȸt����YE,���:p�qf�����j1�{"S���LD�)����v1�P3���H^�km-wWyU}k��g����K�c'%�N�iޥI��������<��)��	6&C����mZ5����^oYƽ����� ����3 K.�0�;��%<��E�㛆.i9����b��:�_A�t�̱@�.ρ�?5�w�E>]��Oo��"��D�Ú�����w�Y�*��͋;��p[��5��2'�H1��(X�,7L@M��H���L�c�V�x�u�w�Y߸]z�?:�Q�ZJ��+���Z���7܂6���@���ُZ�+#Yݝ��e�("����#b���jtۋr����	$�-��[Ϣ�j�T��v�Vu��2�Ʈ�h�[��@]_V(� ��}Y-�ҽ�6��W�M֞3[�e������ �$� H#	 � "I �Id��}��w������>|��Twt������Zk����(����@�a1�������N��^sGN�py� �ؕ�:�cҹ�%�Ts	hM49XJ�W�,xs�7>g"c萪zw_2(�M�*��0̳�{�j�rT�]5�|�C4�q�nj=�ו��=H���zZ�kW��u������Zl <E[��f)�
�B���&�4�Ɇkױ`q���anB��{fb��Q��w�4h:ըS>:�*~��'�o����t���]"4
ǜ�oH$=� ڣG;��6�Z�aͦ#��C/bm���7�G@f
��\LfJO~��zj�1��	,��{�Z+K)�;8KIt��p��(���q�����~�Ί�?�/�B0�E����/M&����m��K;���Z��j�@��aT�(QJN�|ض.b��xlSX�BSkO�L~/<�L�z�;W9�j.��Yu�Է7:��q"ń�kS��~��?��n�����&k�,�?Z�^�n�t�V�R�8�~�����jT�/��	�J`�Ԃ�[�]���p��2Ԥ,R{����7Y�:�Cd}�r���vԦ7�goq�f�μ_��Yŧ6v�ͺ��l5=ݳTci�tf0�=��TZ�Nw����3�ٽ�p���g�;�-���y��J�l�"��1�qk���Du�%q�-b��>�}�՜���STz�x!��W�}z��8.�(�zn��v��;��GS���F�04�(��"��,�{�u�p�rgZ��Gn����f�zT��N��3h��F:{m�⌻EN���]tk�ectv�Ӗ��JM�LdxM3\�#x�᳞6�4��,���ַ^�U�9�U&u�)9+��ݯ�T���SR5�fkܜM�
�iqɘ���{�{�r�a�ŧ�ŋ�r�Q4lLv�N�ws��E���/���ܷ݃,���w�Q�Qv�zz�����G����γs9��qFb�<oIr�m�&waѓ1�����{%��y��5�y��nJ��>o�yqU�޽��U.N�NS��nա9Jľ��c�����<�9�U�B��`'E��q<�Ӛ��ڶQɐh�Ӓ��ꫤo�A	������x���v���u��z���X��>;1��_ֹ��e�܌�֍��P�ooj�_:�Z�sLd�m���ׯ)��_p�wh�=[���U�H���(m��g���{�'b���Qh��~z�b��h�Y|���O��B�NuT��7T��'�^^��� 9�c���H{��}��ԱW�˺J�`d-���{p$g;���~��9;��t�t��7�H�'�/R�qf���]'Gy)���8�:5��zC�6�L�br��ɱ/*]��Eab��*��gN�`BY}N��d�Vh�.��['iUu�߆?R���{,7Ӎj���IV�OPyt��ӑ&�[�TNI�qڋ�ۺ�i���RT̮���E��1�k�_�zh���LÞ�s��aI�c���r�%�-�.az�T�N��v��rqΝ��y�
n{���Nk6����̋)��w����=�b�\��Q��Us��'x��������>��s��+�He���GpD2��̚h�BΑ�ι�v�ءw6�{{���꬗vR�j�����������gxW'z�"�"c�\�e�1��xRN,�w�,~�9�;V%���>޲c�)��n�<@s��+�XD��; sT�EW��ٷ��-��)t�T�aI\�,4�pC\ʠs��#Īr�ʼ�E5�*�]bu�+��걌7��ټ������eN}vîObf�E���b��m;�%��p@%�^����������n$wZ��J��ߠ�t��TƩ�wr�ˬa�O�V��m+��C�(.o�.
=�v-�])�g|'=��󹾕C�����˖���(�1�Ӑ��D8B�i��IE	DC�� ����fӑ�CHA��F"ф��
��~4h5v�+<�a���X��Ud\�O�^�\��1qDV3.7%E<�q�-��y�9�+Z�r��&OӧU<�2�޴m
���!�B��[*��JĶ[|k�((�6�*T[J�����;����r�b���������*AUVF�i)B���Z����j��U�5-S�t���������gi�*ڔ+U�J���*�kiEDb��#[�UT�#��`�#mE�U4L=4����5��IY��e"�*�kʠ���d�1���**%�3.5�#^e%F��0�����W�AE��*V�ԊQe��E�$V(��[A�����[l��b�	�/L8p�ӧ��QR��1UB҂�8�Z��_x�q�V��lQ���QC�8p����Ei�,b�X��\��TDUTL�LE�񡖍(X�e�Ƨ�0���Ώ����	R�_,�"�QUƨ$T��"(���]��0 ��<�TQ.\�WS�(���B�5QQ�2�%Pƕ
/�RI�O���͒�R��x�dwH+z�NFV�d��Ycj����fâo��# �uv'��Es��KwB|&Mɵ���CC�4�!K.5$�_�?"I���H#A�$��|߿>����~l����:_ǖ��Y.�X��O���'�ק�ޙI��,���,y�b��L���fA\��m[�
�'1zᮢ�,�z���#�U~���>���@�]0j�Ȩ���̅J�w�=������L�~���l$&��>��BxBj�L�=����K�D��x���qd8��WKՖi���AcAt�~jN%�8}�0�t�ZDp�ns�>��	���n3S��;/ ��`Y.[B�Ò�K#��]*�K sIzp���#�G��"�M6��mi�Vf�r��{@LK��\��̚�ǥs��O���(搮��hoN0x������n�r��q��#\:�%�vO�"�nǽ1L��M&6�:�(#>�}���A�g����~Ki��͈(���F�fp����y���̠F�$;T��E���=%�4��/vf�/{sgZ߸wo8wq���EzV�g�u��ܸF���y����	{�J��?g[s�������J���n�H��y��� !u;I}��lEC�dK<y-- .�Z�>2Ǉ䁏d���h�7������XEcW�K�5�y��z�{�'�����<��1�y�v�[�l��eb�p�U����Տ|�ﺇP�z��U{��1��-�E���`i5��{2{9s[�F�ӊ���:�g4�`���G�Y2��]��1���=��~�$HD!�H�AIA
��&T���_sຆ�nt�N�I#��e|	���
���9KL��T)�|e�3-I��u����k��n��������O~�i9*f���A�ȶ���6m=cռ#�uދ�s�L\��������}�fq�Q�>�ohW�nx��ɨK�I�*��t��75��]F~J��S%���gx�=H��4`O�Π��|��C �6��A8�Q,���x$��������o/��]���������+�ƥ1�|�Ȝ�rP�0xOْy�8%������٭ð�f�q=��Dۮ�Ǽ�������������m0��m	�<S.{ ��v�fVp�f��x��f��%�0㌙I��NV�"�-�a�^=_͎3�6����	��_K��<��YaCZ�!���j/~�:�}ft=1i�`Ob�/s�GP]4�A����QR4���{�į��4`W�@��v#B��q�u�7㦹��E�H�R�TwH�	��wn"@�4ܙ���n���.�}�;��3��x�S�/0윪��hOH���V�~ғ�XZg�U>��_�K˙*�u�F��|�'�:����B��}��B�Y���342/b�H��.f�yzf��HxA~�{����7�m�B_���@�x�Y:Nrl��DdX��f��O�|�Y�����LoD�
��f�鱿Vv��-K�17v�ޚ˖������W�}�$"$$$�F�! # `�����j	Kvj����Wn�ރY|ǂ�(����Րnh����m�Z��QN�P��'cU؋��Oն'��ym���鬂�.+�&-b[�b<V2���:�uY�u�҃�m$��#4Ë8��ż�xZ���V�)��,}�� ���fq����m�u�R�\8-�f�}y��Lhq�.��1m&:HDYz�x5�%ݰ��1Rz��x�NM�� mpgCY
���L[e9�3g�//�M�'��8�2&!����B�A%je�����pRO�bO���g�+W=]y��+a �rnj���f��l�ؑ-	QǾ�n��
���5�-��G=;�.^TT�S�
7 �����A	��Zg�;�Y����/i{E:��%�ޫ��~}�M�mz��W�,9�2�����M����=���2��n<��Ki˹���%��"L�S�\[!����D�E�s���������;��\��=;*�vBw'�����9w��x��j�QN.�gH�d[B��ow��;��Ϭ|�6ϻn�l1iu��%������,G�\�0`2ǫ�Vu޷�=H'*l6k=����2�L�0w6�u��f�T�5otmb��*���(�V��gc7W��H��5������ͩG���e"m�݃�܃_ ���r�}�?FH0 "B �@ $ PD�I�Ͼ~o�������!�C��7O���3��c��s[I��|�(�`��x3�-���w�ohP���F��������.���~�s��,��h��)��Ͳ.��d&��E��5$nU�ڱ�t��d9�W���S�
��!��|w埢�.�dI��«�es�dL�B����zt��j���WOK�U�w�%<;�ݮ��>�O���ɅC��<4s��B�sDV���I��)n��*,(,���r��!��]|���\�7�u����񊤌3���kM:�eDw~A��j)��е�QS���Tm	�����Ã�������v!vs?Z;�@z�U�e�{\�kg �t�=�i����z�-A����z���uk7�Ρn������V�`L3$�l�l�;(���$���Y��l�0�f�ۭ喥g�?@Tؔgםyw@���6*j|�������w��Jރ�
}�\޽��5}�Zi���$28f|������ϰ^��!��<� y��5�eSU���?�|�U������d�է�f�n�{���g4�N�K����b1s�TGw=P�v�>j���4۸v����<8y�c��N�3�j��{#��N͐rm��w�E��:�oel�1�����%v��V���e�2n��$'s�մ�}��v��vA2�!�d�$��d�!������X@F "�����i���ö4�䠍t������R�����:(����0'�;�E�-hM��NEM�U��"�1xKf�U-m\L��u�d|�(Q��󇡳����j��s�1�|t�K&�����]S��m.n���󣑍�6a��t!)���L�)��vл=;�^ǫxfb��+(�(�Rɑӎ$�P��d���:�Ar�!2!<N��iT�8��T�^���� �9�K��w�i�����D��G?����{a�����,�2K�/ź�l\�5�񆲲���]������I�.w����V�d��Gܨ~����i��.�VΟ�;1��fҍr;>�����N>ҙ����g��:׉ �& �ጜ3���=B1��9
|�����˹��yHfժ�;
v��WK՘���T4�L?5'�`>Ϙ`�8�:ne�½}U��m�����	�N�S�PX���Q��j;��X.hw=yd�ۇ:��,� a������z�3:�q�6�L������:�M6,�-L�:�x�i���/~������4'[��]�1N�x|�5��aZ�аL��=A���Oq����T�F��]0y��}��g�/~�H;Z3?~�ċ�}���`cN�f/���F0�Fﭫ#��)<�p!�jd%�H�|�z޵\]�]��}��8�^�o�M��m�|<��w���$��B�A@FB�"0 �@����y�Pg�T��`0o��%���O�ٲ�k:m����'̣�����q߻M�$N�d�T8�:��a�f��8�[Ϙ'��S����jj�<lD~[ ���|��E̷[��͸�b�D]�/u�@8Kϳ�D[����1N�A����\:�e�������[̞Bgo8m��A�,��}�@ >��� ��H؊��xg� ����t:�-KCt[b�^�>�h�q%�T5�qK4�d�Ee��<��]��b����B�+ne�`�sn������hV��S������S1����˒�k�vPcAd�����I���:��L���_��D�In�^JR)� !Ŵ��EǦB��؜��W�aSe�5QB�8~�av�Kϵ�g#��{�w��_w?���V��O։^1pXp���p_v��������N'y��v���U�j��l�%��E�B2%>[�kS:sOn� ��'�����]� ��eÓ�����f*5��gy����ŷ�)Ղ�SH�kk���P�:= ��t��&M�NAy�lζn�ܯg��(uc�d�Z)��`h���XZ���6��+M5����b�6{VZ��VY�W,��IsL�꾙h�5&�as:޵�=�T�u+U�<\y�o��bܩq[�(��}��G���R��b$��}We���{v� O� ��@FIa "H�"0�F�w;�Ϟ~~�Q����N��팇�J��X��ay���q��y�Ac���dr���Vŷȴs�Dw+���y<��ʘ!�r'��0��YC����S�-��n��L&2����{�dwioB:�9���5���"Yk�����eB�����	��O��6�9gT%;ӣ1���o���xwh��3�C���ɸ��]���B;���oJN9UF��S�׬j��)9�k����.����^523]�f�F��C��������%��Cx�B�|S��y�Gdʾƍ!�V�+Ͱ�u��z\�75�d	��Ƅ
ǌ�֟�z�����>K�E��y���Sɝ�z��U�Rpl2�8����n���q|��4?3��P=�ܹ+���#G �SUz^�d�:���48�m �,���:I�^��r�0�C;��a.�ü�8��u�CP�-b&�����:=���	��<�EHA��k-��ma��^2w��˗z���Z{[8>A���{�d^�UϪ�&�VA!�vA�i�����HK���e�K�'�_�f0C�r\^��wnۇ	8~���<�{SX���S��W<�κ1]v�p�ᡝҩ�<�6;v5�f`�����>�N�Ӂ�����;�<�R��e��=f��g��8�d�-�7v�v��~|�����d��	B$ � D"R���Y[$3w���n�tn���b�{���h_ y�^3�v?�/,�5띪h��!����D�	�d	c^��J��ք�!��Z�,X������EZ?}��
���9���������b������m��S������(,T)\�����U��f�b`?�?����+�]q1tyGY��t%	�.�rG	���:!2/`�Ju`82���RS��FN0�nE�)n��+�D���}��q8����m�$C�e#�]�4�t�ޕI�x��X�E�.4�s�.��xq0��78b�����uo$fF J#Za�s�c��1��P�}RS�yd]���|��8m{m'�)O��z�M6$S6AڰC��>���)�@��F��aY٣����^UΪ�}���!�s��rą�S#�7�k!|v �����x.�u�/T]w����uY��:Ё�u+qv9*,+�:y�X�Z��{[=8x��A��h��w��nһ�#D(b�e#�P�����s�s��1��5.�<�^��!���OKbMYݹz>��sv��CxFO*+}mְfGj�۹�?�'�^�K�SËق�����.%�軱C�������I`�����m��ٙ��v��#�q��:���9�#'����'f�C)��7����˹����c+�z�;<�)��W�s+y���"'�$?FI ���2 � � ����=.��dRL��/Pw�H�-"��ρ�`��`Z�	XY殚�~P&�q�nj��\�t�P2��v�_�g�r�q/
ߠ*�F	���a?��
Yk�'��`��ߧ��'˹�m@������R󞹘���������:9CX��Pr�?�a�Y��%һXB���ٴ��V^b��z�����ʭŻ��a
�@����������fN�=C< E�>bJˉ�\$�/V�̯VǦ=�':��w�&rղ��\[��?��"k�7N��O�������lX ԜI2t�t�ȭZ;[���B��Ɇ�<�,tv<�*�̠h��͋���T9��L�C���3Z�th"Y �Bi�5��ь���a@t�)���-���vУј��zF\��&�'��U�2��v����Bq-s耈�Z�3���RZ!*���'W�S���:�>M5�fk�.��xN� ��阫���?R��"��_�B`$�4$v��BN���c���1v����'6�m������L(?;���P�d�ɴ�#�Y������z�/�g2�*�C��7��4���P������w7�e�wf��,7��αOu�Y��[qR��o:+WX����C]^13>�>��TC�c닽�>㆓ޠ)y��F/G<�:�<4��k����.My�'��n6��=�3��<�s5�۞o��7���ĐD�#`�����#	�ڦ�@���K�b������x�4���r��k�S ��7M��a5/�1�g�6��k��B��0��;N��->���,it�~jN%��}��=�An���:u��&Ö�����?WT	L9�v�=c$�0�֣YEC���FzG5�����Sdqft�S�t#�\�p[��ֹ�1-�fD�Ξ��Хs�A/r�)@���t��3�<����h��K�-�����"f�ha<^�;[��;j�=,��.��+��̸���~�k�5f��wb�㠺5��f��A��`�4s	��y@֜�d����o���<+5A[�=�l8`���+�Q�i|��S�����cSK�x��q1*}gϷ��ar����r�jz�
�����H�X�w��	�=N��[�	�5Վ�����`���#���]��9s/zc�R�FE�ޯE���4״�a�\�50�E�Zz%�����3n�������S�Y�"KH�dK�e�]T�y�rĳH\�3P9A�����w�,x �v#��P" i�OB��8�r�e;�WX�� �Sk4���=��ZWsA7��}�>�X�m�#����1�DZ�<��n*��Qxg���dy�G��-O�Ö/	�)u����Y�tD2�^C[�������
.�aӑZ�o��YlY˙|�z�k0k���;w2�i�&�3|��xM
���������7��~�Wa�{W�/.��B�m/�I�O�ϸ&�D���%A�n�+e��Ը�\̦��4u��2bٷyʰ���m*<��ޚ0��rs%��\�t�d��q)��!�зt9�vv�[�Vj[���5���37�+��e�]���۞Ʀ�W�����F�����DF����+-�ӭ�S�nvL�p<�Ni�O�O
uY]���Z�'tUvg�Ր��C�<�����l�qHl,��:�����Db��I�v�5[��3(!�YB���5�]��'��EӜ�,s9VQ�B�i�p�G�0��M8��ˣ�S�H�ɿ�Ps���y�"�.[b���)q6c�+�`�77�Q��	%nl�%�]7&�ҭ�J�[�A	��^q"�ݧB<��"ᑪc����i��ngEy{x]�+��f��3��v�=�]���eh}L(gxg�k���b�>�u�|~�AD>��vtY6�	r���m�}�ܩΆ��J3V�kS<����:�+�V@�ͮ9j���O��	(Ǥe�}�]��c��~�G5Y.XHCC[∪�$?R�8g:�ݔq��:e����} �DWXW3��!Fo�"��۔�C�oe-�C�$�K�.a[�_��6�*�]�q6��b%p=�M�v� ?i���=��S4u�����b/͟j��sqK�t*���<�%]vI�F��NvR��qd	1�$��?.;�]�tzx�,na0�8�:<!�r8��C��qlwigNJs����/��w��4�����3���3�n:D]�0�Vb<�Lܺ�"�<\�S�m;���0=��`���o=҆�x)�F�p�1��N�;��j�60�f֘��1��
WVn>��<if8�"�����&*�]n���ʹ��$N�� ���վI6�n�SuY�N��wb�T�]��sa������yq_~Y��}4m�t��f�$u��Ҧ�5�$��t��1����V���aS�ٔ���F�;.Z=�<2["�ho��.��u��zF�J��0��wk�{۶�eՔs��ݒN�7����F��	(B�Τ�f��+�A�Kk9�����{1锓}0�m�k���懺$w�c{\�~�ܥK�~�t���[��y�����\7�?3�z��v���]�y�殠�n9���I`?MX��c��!U��Xח�g\C��z9��rU�)����B�3.�m��*��|�v���T̼����$I?��	#� �j�Ӗ�1)|lb��ETQEF,W�ሇ�0�ӧ'jF�RVPO�Pc�YQKj�[['��D��������>6��)��*�	l(����-Ʊ�XR8ԭ�:t��tUkQ�f�LC_1��<f.YQ-�APON==;:�x�b6�bxA(�J�S.a**�nS2��K�8^Z�\�F,�(�"/Vrر=0���Ӭ�0E#�p�r�EQQV)��ּ��S+B�J��b�2*�(�za��ӼgD�� �Q<j�1[B�em`�P�PX֌UD��;>��F����PDFV�QV�T�*�Db��"����==;�UAE_)�J&Q�����X�F"�a<����J���+"�+Q[b�#�UL�QKJƵ���8�E��*��O������O/��C(�6�ِ��Y�w��fgzӶ�wH�5�/7�����;�^{��>�ܹ��~fl�H�"D�� D�D"!p�O�h���W�#�D3��dS�Xqm��X:d���3l	�	ȯJ�;��A�
��#Y�hٚc�yymx��������;^�ս[�z��3��`�a�����Y*����|��kۋ(�gC��\9���itT�N�K�k{n�Ξ}On���]���"Sq]�p��ԅ{�U�͏ʃ`~�琺d�N]�X��[]$i5��7$Od\:�tzqmnW��Q+7]-ܙ7�����ɛ�C�Ǯ���P�F�*I��&+���Xkх������h5JT�����O0"C�"rp���D51d� �FS���摋�F��'��(��e����l�����bc��τ ѯ��ٛS��m0%sɨ	��YMdU*���+]n������Xq�5�DxjdpyPk���6-|�=��U��2�����,��ۼ�B:�Q.�<����L���wfcx-!�-�?4|���o���;���K��B�ؔé�k-{���_�����,F\�������1����~y[mS�Z�ɸ���r+�Wv�r�VJ"��e�k�>Z��F�|�Ceb�"���.���짾^r�B��yoL�����뗼֨�X���������|��:]�6�0s<+1m_(⧂j���uϝ��o�y�y��H~�$Y$�a"0"0"!"2���{��ҕm�Z-��d���Δ�eޚaC�@��)�G�Z������	���xc�/���u⏅S���#�����F4(q�.��77�q����k�Ҍ�/W	I�,ݭu��c<+�.�;!n�8��H���l��/�J�8_�6'�l"4���!��j�T�v�(d:k/^�x[�ǰ((EÇ�#ʬ�U^Ͳ��A�����}Ǭ�D�"�{NI^�d4��`u�-�9ר~��#���o,,L܀�tRQ%=^k�ΚZѼ%��c%���Y�A= ��+�����{�O��3�����<W��1���Ƭ7{��_u3jyv]s��!��z!Z��2>X�R�=Ķ��N5{�\�\�Ɓ3,�zL�I�eWklOV���duL�;���-���r�	� �!IO!�����b5@Q�`=��~��Z*���@������g����G��nloJ��x	��y^�*�S%�9���k,�m=��s�A����@�8F4ä�^�y�,��WL����A9ϻ���̌�E�:Q�<g
��N�>�?.���z%_�&�u��k7\;�K�;�q��y��i�g=æf���I2�&�ݼ�ë�d�3{����V�˶V�ˡ�*q�}����쳴�C���е�ٓ�^�uF,&P,�+Zҙ�	?H#I$�#����" f���o����]z����୶�~O@O^�M#il�=y�6�x8zh8X�?\�%�t��N�&l�k��M�$��;`�XA׆^9r�ߒ��r�a�O��Ɍv6�:l���y�'��U:z��S�VC�YAV:�]�������m��Z�B{mi��B�)S1��vDۼ���k��y�ƶД��<ݦ����$��8Ԯ{A/mbTP�yu�����]u�u�!UmJ�3mA"�P`��38�g��:ב̮Eek�3��B�}�,)�ÍKsS��h��%����W{z7B��{��6C3��<{D&��~��d�o!�'ת�/�<����[Z�+�-�H���:�6  tG��8�t�a�B{��(��Y;>���D_��p]��t��f��}�ݤ�.�C����OL4�m#^)Ẳ3�`L�"��j���'���� <�f{gҥ1���m�~����x����<�Vh���&��.6�7C�>�3�G0����k*�Ǭ6���n���{P%V�L����B�:� �B���9��6m���C�ܿ8�.U
[��4e,�ui9���={z.Y���{d�K��ka��Co�*ŔlK�ESrxڻ[�X��-�M���J���Kr�g܆s�-�;�կ�����}�O9$"�����-���*��fi�JJx\V�(���&B+���~��P�Y�0�2A�#�3  ����j��R�����c�Z�!<�d�N�a�D&��R%�D��]�v��e�ӻ*�jut,�^=�p0lcs���`$U�A�<�Є�\b��1����u}�Rz7��9�^׶~y��y-�,�}���ώy�!>�W�ʨ�U[&��Ֆ����??�]�k^%�=��b�q)�?D󆺏B|\@.�u�-`�����pB��p��uqZ1����u�(�hc��.�]l���u�y�6�54���lM��I�<v�-�1|:B��2�5㦈k읥$S��8ŧ��yt�~j	ı�A���g�ڹ�K{7��N���������Q^_n��8���/��0�j5�P*�b^� s5шm����e�̽%��U8t'�;���S�Z�^���Ch��̚�z�O��)��^1^����?o���	����C2�~/>�mt���owyՌB�N�ʓ���K&t>������`�\gӏ@�$�nY�H1A�������!yx5�b��c��$#���I�w��L׭1���5y�{G���Vs��h?b3x����z��=�O���\��F�Y�]?���Z��ѥ�z�5h��7����>7x�m��WY����S�Kt[8.{�\���)�Ǎ}WY�l����{���b�bl��	?D��dR"H�2Dd<���=����G����>�����O�R&���������Y��ɿ���4?���X�59���4-�~�3n���!�@άa#z	D� ��k�[�=Q��ε�ڧc���tU�#}q�e�*5����=Kսͯ@���i��%�W��p�R2a��ŧ4���h�H�BX���Z�}X��֨������#b�}<��˒�cn�r1l9��q(��%}웰�ݽ��OJ�/�nK��Ew1�Xqmâ�o�`��:'"���Mj��g��,��S�w��f����a�/��dh�;�_�U��B�(�͛V"����Al��h���asa���Y��lx���*d<���1,��)M2�(Х�
�n,�����%����M�=1⧏5�ͩ�T�@!�y�tBd��D�6T�cIMl�p0vE��f<�Ƚ���
{!_a}�5���uYr�0�5�ܻ;���F�I��&�W�yh��|B5�y�����\��b��o�\�n/9|a@���؄��7$Iz�a���z������s0��=�y.�7&������xl��)!m����-������t�m�!�<ʏ#*�ongW��,�u.���g~��xD`��צS�~AØ�Lj�I]���z�)h׶�x�X�5�#�*������f�N�����|���~c����~f�䟃 ��F2,F�DY>}��w��ΆD1��3L8�~�lO�p�0�~e�Ck����P��+�5�ki��дj�Gf��or�.���'�'�q �=�y���@B��
�����N��Wˬ�1��j�J����$P���Ӽ��t�*�_L}q��v�/�@!��D;E�pRm�kz��T�{ngB�N؅�h�&�,t8�������(4vk�ACB��v��d����dhE������d�#s�m�I��t��OU���J~3��=���>��/b�=���5���4��(&�K�1���倣��K�2�Ԧ�^��z�n\0�V�گxs�X�=��נq�ߚ�a'�Mi��Ϣ����A�i�GZ�m�D����HdαR��B5����@f�\F�a�����^.��UϪ�)�d&��ƭҹ�ڎ��h��5%�CP(�i�L�tgO#���X0,2Ob��gbh��8��*���d�և��,sX=@y��]k=��0���fA8��.�eq�v�&���W�Z�oj;90%]�u�t39�p��PŹU�NF���/>��x���g5~yޔc��jk�i�$eѻ�{�dwMAp�@ofѬW�WN�r��tFOF���ţ��D�:��V�/%tj���-�iLa��Ě��:d����0�i�"As�~��2�a�FA"0$A`� 	��OT�����q��=;H�8ū&;��!Z��2VdI�:�Yx�N7K�=-ۋ���2kqY��Tΐ�޷0.S�\�%��tBd^�D�V
TB��[����ʨ�W�7&�;Izh��P�9AñXٗn>�A���e��&J�''�0�YB�^Č�������P}��{��p�3 AE����	�b��ʁ�P�g���hes�,Yq�ò�[�M��x�\�6�����Ʒg�Gڳ�X߹P����q��M;X���՛���#�����0��s�Q�I>z�P.mr�a!<;���Zk!q۟s�Þ����g��_�4+�o�d닿�E�ΎcR�/��3� ���|�ڞaa��y�a�@s�vp��6u01���B�x8�x��\��'��OG0��g3]lQt"M��.�u�·|Y���4!��dF�ve�++�&���`2�Mc߇('Tj�b�Y�F͍� �>j��'߻���z `O��AO���������ƎK�W�χ��f�W�o#�>n��M5N1�f�*��t3����q�S��U�w���b#и�l﵈c�O�g�u/�wq���j�B��䟖L�^^n/��e�����)�72[/�}
[�B�n�#z�V`J�ӓ��iS���;�k����צ*�}[r-����~oϟ9�!�H�F10o0`<��� n�O$�SԌ��'�� ������,�)�%�� �@h�/0���W���ӆm��CFo�u�Q���
�4O��P<���'�N�fjt��@������l�ܭs껠��K���PxB����g�#Pyn�<�\&�A��;�!c�"��Y�j|8`[�5�uWF�t� ��H�ɤ�Uz��i<d,{a4�(JN�|ض	�p�7)�gUu]�ts쫇(�3����t� O>�#�Dd��0IlBL�ʖ*�b�j�z�)��sob�i��&�,1x��Ot���'�,!�@$j��j5�t!)��I+��em��ɼ�Ξ�̽vvk���=8�5B*��l�={����C�1�A�0y�c@ �v̘�\��F�gy�^Ad��8^%�{��ג4�S�_8o]D'���s�-ud���[���Wڜ5*搧������Rt�_�T�� ���#�y�/I���a��/��{���G`��Лla�+N҇�z^�����,H]&���d�co��Rj�t�>��i5e�<����MĿNp��qKxk<���l��ν��{$�3,��٪J��4��/a�P���{Π�.��]�����eb(7��ϛ���FZ���z��{3�����Ls��]V� �8�G�;4w[�F�;�Y�Ur��.�F��q�ǟ����+�P}A$D�D��`�A �����e
��Dy�?0r���B5�C�u^�mW0�Ŵ.��0�i�k)�U眳Y��S��ݻٹ������ܩ�X_�z��4ڹ�s�K-����R�����V)�˼�U���3�׹ +�H707:-��A�G�A켈v#�5d�6��ٛm�K4���k�or�n�P��_l>�r_�|T&T
=5�V�a?��:s�׾�T*4D*�:�fԙ�a���K���e"~]�t�~?,]�>���/���3����a���������$W��y��4#�&8���W�m�:��6�|N�h&��c���C���v���/�F��y�m[9�:L:nNE�����fע����Aa�
�R2aŤ�zU�m=6���9��Ы���xiǖx�	�����9ʩ����[.JY���8��][٪��F���XS/;A�پ|j+�b+F0��(����b��~�'��F"(�gN��٠�j��Mi�[���ǫz�����Q��0E0�C�_�P���w�yXP�fԵG�;:���� �����P��=ۮ�>B�/�Z�\���,L-��e�X���
���zQ�ʩ�H�Y����DOun��|!sxs=�_�ڻFwGQG�_"59hI}�����$a{z`�/|�����dD���� 30on9�% ٓ(g�M�Bq@r�d^ʰ��d�B�(�|j휼�{w�>k����Y�wr+�[%zdOy�2�녯>��t�d������T�kqA#i�����ǨuW��G>N�n�zM�޻Wp���l)ߡ,A��;����w�RO���&*��fҢ��w<�3C�@Q�ː�/wв]y�y�"؆�������Sw2�P��;��[c.}b��g�l�g��Z�잜~����
i�摫Ǧ�H&�l(O�S�0�[��<2ׯmt�u���xsӮ�[&{�ﴒ��t�e/EGs�|w#�!'��!�1����_�H&��Ҿ���Z���X�(�?J�xF��5ߴ�N)gO���L���wf�3�X@!�oGu�B����#��SK�u.�v)��Ė�,}���u�d�G�u�v��C�m'$&o�N4��^B%�H�,��2|���i�n[�qk9�W5�nZ7t,cB��\�u|�{��xV�͈QO����0��~���*�^}���{�Ir]�����{��q�D'm��iz9Z\.�VGOD�8�X�=�H�f�r��/����1��}˰BFgm��:p񙗒��h/�.�o-�d�5	f�͗�(�id�������<H�:�%���Xx��x��7"�f'�E�{�����ß���}[���Y�P僻w��l��㶝�&>S5�,(қB�C�u�� �U[�w����e�}{�^BS0C�x�˧)�S��� � �.�l�X֥�� rغ���цST��pů�7zj4`�Ǩ�j�]�*c]u�Ga�MrW�s)��n���P�H�+�gs/D�8z{%�<��|�k#|�ҽ���¡:�p�͕}b湁�t��'8�0:.��7�'3�
��M�����t�8�{�Yggvs�ϰU����74�ys��;�˖�i���"�+.Ӿ˃oyΧ�pZT���k�*u��yW��'L�<�ז��N5-K�}�J����F�/^�LS{^���羙����g���jYB�E�ΟHV^�����%Yw�Ƒ���W� �r�7yH�w� v}��=�X�c��!��<���1�d�K��4՜z2�!���d�ūU��ǘ���k+�*��`�O��k�t5��}P�ɵ[�9N�h���#���/�)�1��<coW�� �Q��Q[{��s���G�RgO��Su��=�	�j�Ts���r������F�w9"�c3;X��� �t��F�6���|ԝ�/�RW��cCW;�`$�S����B�`�W�t2Jc_r���"sKdQ(,C�i =<3F��l�
T��|��c�٘�ңǄ�gz�U;z�F��ۙ�	�{�NU,ɼnG����^��f���~,�t�jn�vv���Kɋ �ӎ� :IO||5�� ^��5խt�|�>	����;��Q�$���K���O4�ZMUr���w�e��;��!.�N��<
/v��#%Sc�ۦx�4�}����c*��&��z���3�D�e�o�<ьx�.
�����䞡}�{,�oU�AJ�n���;jɝ[�a�����,K��=�7�3<�s�xp^S=�l�` �B#)�O2Z���H�YM+�H��u6$�̢�K$"P��M��+n��pv���fH�$ję�98�1�[��X�Gu�V�&&��>���~��NLR/���O�Ӽy�dɣz����
׎��h��'�=uۗ{Gt^ϭ��P���A���	u�A�Ϫ�"�K�Ţ���]l�����'�3��y&���k&1پ{�'��fn,t2WUbT�;Xr�zQãrf��=���~���0���*ini�����b+6�hE�ҙ��i�g7iД����x�yi~Ӟ͝�ˣ6��tR�b�`7�Z�f]�ʧ�
�����,J��F�<�=��vU5j��s����w��d�w]�&K�*`�	�{��i�v��U�)L�[(#TUDb�i���Q0�h"�$��!�� H7
a�wT)��)�0��检���i:�U"�/��8�3��o39pG���Q���PF"�[*�X��0*���hQ�UP|��Q��a��t^���*�R�.?9��JqYiYDmiAdF+mQJ-���#=J0Y���t��"���(�b�r�X��DC�aǐ��q�Y���(<�U�u�4k*c�U�X�Z�Xħ�ON��{J%eDUU#-���00˙E�8Ҵ�J�����娬`�t���Ν����T���R�<a�*���U�1D`�**�3�R�r�/-�TQKJ�,b,Tְ`��N�{;;���eɍ�V��e��m���˗�Qܡ�,���ON���:,N҅�#e�H�i�ǎEQN[�S�X��Yx��j�*��F%=8zt�핬���b��2TQ���b�/��Z�(��2֕VN&cs%�hV癈�=8zt�F�f	.�E�e�T���_��A�|���ڵ��i\ex�DƢ�5�P��Z�<�aF��8��V[�Uq�eȱP��^5ڊ�֑���<��/9���[�K����4^[Ys]�ǚTuX���P���.ˬ�·\u�b�J��W��bۍWu�yŭf�n��}!�n��NXf\�����0�FEF�� � Z��}E�����@�e����T9Y_M�%�!�������Oӫޟ��R胷3�\����`��F��4��P�j ��'�x9���ğd5n��RAS�^%��<B�d��x_	��l����/�l@���FCM��.qL��s��`h��P���a�<�7u��n����zg�-�ȫj�'�:�'+ ��zX��{1P.����b��4y��=�w�Վ��'=D��J}R�/ v�2l�<��C,u�*X�R�*��1ۋk�\\���w	ݎ霕p�����ހ�I�.��N�3$p����	�{1�YJ�ӝ�V�"��:�;����ӌPgOd[A�t�z$��] �}C)r����!��ԩ2zWb���A�7ұ�m������O��@%v�f0���ၯ�\�����cBj�+������8��������^�E2.�s�-#4��vk��T
� J��!���~��c�_��ݗ'+�mN֫v�+h����\��r�'�����T0���vC��p�m��V(O߸{�%pG���8����N���;��<�^ŭQ:����Ʃ=x���n�+���3����9~vE�o�o�P�	~��F�d�ʏ:����>2���X*�cx`���r��oi�ݛ�&���;����N�b�ߞ��>��w�'�F#cfo0`����~�����r^��9�khd닾*��	���:��sӇ��qn͌�9�r���:�@ ��A�<E>p�F0�7=B��9�B���r���2��n+b&aK�~�����Pz�K~�|�	?��(�_晕�e�9*�e�X�Y�{7G$Z����'��G�Rz/d3�tj��h�����G`�fI�fǝ��)߽����쭂��ʘ �$�ݏ@q�hh�cc�¼���cA�+j?������Оqb���0�kݴ� ^E�![� ��1�c���tg�5`j�3Ռ�b.9���g�V^bټ/:$�l{Ԃ�:��O,��c^9�������"g�A�]6��<�\��t���U�Y��.uK:AaÝq#�w5��P'�۔-��=��=(5PY��i)$t���Oc<�B��~^�ﰹ�����|����mc��È�Q���԰�o)��	��~w,�,Z7+�����Vo��7�b��3?R�����Ci{A��}B��4;T�g�h��Գ7�,�S�z�zɩhz��/tY�3z��a	�*�
WC}�%�:h�hR�[���=�NQ�#/�{a�����<d}�7��U�髗n�{�Up7ȱ*O/>,g�n~�d�Х�����b�E�z�k�J�cϟ3��r��۟7~|��E#(�Q��
�L.�^����O:�%)�gEH�{3���AJ�b,������0x]тwc`EWa�y���>ZfJu��Y'�.�b�����\p{���5���5�1=��]2��,a�K��}��d(}�"��3��<�%�C��r��^��(Ƕ�����5s �f�BeB`)���*��֡Č	�z_��~n+$��f����� �s<����n��A�=������D�~>8h=J):��<��ǧ$V�Ta�Z�e�U�\��3�E-}�n�"%՘	��:�x��,:<�2��بuض\e��U��2�dFTF-G)�A��D���%�+����z셳�� ���?�Q���
�A-�����t�}�'���T�ܽ�cBu<#�}�ǧ�`�Q���@�5���^��w�b�~?��Yn�|�}g������?/P΁���.�����1�C���;C�ƺ�E�����gt+b�3�(�й�X��7�r����}����7���H�g�S��� ��S���п?�G�9��~���ݔ
���.lӇ�}�Rmr��ˎ��Q����6��y�bY�9���n8�y�߷9��1�Л�8��^���XK����S���CZKk��k�<U)�\V�=���m{����oO3��7����Q�D�I�����̵�e\?����4y��"D&����Ѽ�����7���+( n��ݩ�55��Tc_�v��0�b�V#��o)B���a�0·s��*��ʿn;3�J��b�4Ɇ���:��7?	qrHk@��<k���6_ʀ�e}AI;j�#N���u����*nUMFf�	z�^Ab͖8���D���q�x�^=�y����؂�r,E�p���=f������2 �4��mA�:��
�z��tB	�{�K&�x�4��^Q����{gNE�whAT�N��Q*�2��\t.�L�)�X[4_����"S�H�44��ropۑ
Zb��-���ů�S|�Q�<�@<J2�0�@��vv8�wR���LU�Ȣ[L_�]�c�m=�e�d1Fsн��=Lc@��C����nA����̿?�~jd��t�vVgGn�^��1ov��-#��k�3����e��#��xX�+�?��ٛQ�q6����ѫ�ߘ��i�B��\�@�C�{Tw='�qE��[�� �3|��90��I64�Y ���j���4��X�f2;�����������o83��/��'���Y��[��1�l�`�d'W��N���y���B�ڝ�;��mqBfOI���]���cMM8d�6yE�΋z��6�o8�k���j�`���Y�g%�T�<�˜s��矰�ED`�� �oy�^wBP�r�,B��6���z��L'
�Ξ/V)O�T��zwf�����>��:�Z����O�*4#.�;S��K���ڠ-X1%�W�Ʋ׾>��T�<����$w�����{)A�V|��Ι3��Ɩ�A� � ~<c_���g�b�;:Rpm�M0�-���sc�<�GL๮���cmm�<ܦ���{(D�J`�4�;���2U�A��;hk�U��,K(y����ַ��Y����r �;�q��͂,��68k�N?�D=5��l����uY��O���	@� �k�!��L4��֞�<���g=��y
�$FbJ�,9���x׭+��b���� 35�Oa@���4
�ͅP���`:{w\'j[g@���w��7��J�3z�FEH\�vxR\P+���SØ�"D>���S����s͎�;C�[vVK�s��erPX3� �ۆW!8#��)���U��]7
�x����+�\6�p���5�D��e:��V:��g.LV�x\#��HVS�@Y8N.%�N�F���n�������<;�+�\,�m�҇WmuM�v�ޤ�0!�_l��X*�f0��W�����pwn�\�^�rZcJ/��ï��n�(�7U;	,����_�y}<�����m?O�F�#EE�B�Z�G\������[���W,q�;2 �nB܅��7�}��6���:z�ۂ��>������@�\��y2�l���Ng1�#!��$h��d.��8���G���Q�/�г%P��ƺ3�\�F�c`��f]�Id�%}fv/�zCٱ=ݝ��Ue8�Xʁ]�t������XܮV2�z��vެ�����+A,�5�.�T���ʡ��,�37W���`���<jˮ�f��`a0�U⺄v)�4���ӫk�u*Y�����oɪ�p~�Uޑu�݆��L�m;~Й��1C�Q7ڽY�8"%E�G^�qA3@�19�����7�鋞;�Q�l1�!��1猾�	e5�)x'+�pܢD?Sa�UL$�#����Ӧ��C:E��;q�ӱ��ױx����$"�T3p>����É#I烢�^_�ae�f���xꛇ�:���[�K�M�0�5�DC9�pέ��a<ާ@���,�^q��f�1���a�[J���&jŶ�C��;��sC�.JLЃLͧ�&0Q����w�����B/^�o�s{d�Ֆ�R-E��kpv$Ӽ��̓Vև���?��U"(�(�DB{�~?;��i�~��������#׋�4��<U!�w&��B&�i6�'��p���]6�����1�`��+o�Pdm� ���1��dw�8����z�'>���}�w8}}[��l�\XK<="���J1�!��T������n:c��ie w���õt(K�9��t�ͬ��H�T�����,)���Ij�]��(5\�b���	�IJ�\*�'��	�@7���P!����[>^�i�ZL�|�zRW��-��M�vr��^���=���Z�%�-T��<�㟒�9�z�{
/�y�v�p�w�9�`�+�23�m̱E{ܛ0��ɱ� ��ƭ�ΞC�~ ��8Յ�����^Y�����ww��v������0�/,Lp�ȆS�I�ڽ�*������3��О9�Mא77��S}��.�L_:��`��gj@ٕO�et��9�R��J�0����QH����闂�9�>�ik��^��o|�P>����@p�t-&��y�)����F�b��tC�صϗV^�
��{M�Za�g�܆��v���ӊ�NWs�����pࠑ�xt3�g�v��1oNR�zvF���U|>����#Dd���B+ʳք�Y�.�Q^��Щ���hW��8��`�aǠ��~��]Lc�Y��4�v[�܃�sG@�#�#C�Q���@�����%�&%�2!���߬gj��[jo�=.@�	-�6!4M��������<ɞ���m�	��j��ZW��/o�w�	�g۪�h:�/vӾ?_��Ǘ1>���P�$���(����u�~�'��t3�cTSݫ6ʋ���#o\�V��:�j:<�(��P���l3��5Y�v���w���3qs�PZu�6��2��������e�z�N�1�C.�=G��\^0���}� R��;j�z�ni���+�[/d���O���Ե�jq(Os�\-��I��T���I�F�r5[�sޑ:�Q��i�uUn��s��:�����p�;H�H�<�I�����|�uS�E;�U��8%���c�
��P��Ūۧ�Lu��Q��-��z!a�7�9�v�3�Ӽ�8�V��/<ɽ���87��QY��G��}������x�p�O�_f��(BJHoZ�Q��1��x]�F*n�q���*�Jq���IV��vt{3((RN�9�/-�1����X�T�A� ���vu���g�+�Do�Y[�b�#��H@~M�s�z(u��=Ú1QM�s1�*����g�ؼi{�ØB��|/���ϭ����0)(��Cc ���n�z2�II�-kd��]�~��r7��l�9��v*e�*����C�V�2)6O����gm��C6<���(7�e�w;��o'7!���~1ϣ��uCypT���J}`Ld��f��oyVd�k�]y�q���I
,9���Y�ǁ՛ǽ�Pv<rFJ^���a}̵u�H�;V�k�l"��pE�:�5d��|�Pc���[��s�[{m�8��{7Փ�s�}ׁh�<+ڋIVn��1j2}in��~���n�y��fhh�A��b�!h�|i��q���	!QW%�{c�}�˽���M=��xm���AZؑ�xID@=���s�4[�����Q��R�l��{���T�����w�-�M�B�J�4Jw@�lV��2�&i���;_�w]÷(��M��ݤ���\�!���0x=u���P�Q$"�Y9cj�����l
�֮:�\xu�p��U��Br�.�\�a�NT$k�v�-j���k�{���o�����7���?T"�H"�+���Z������u�Hv��U� �,<�yj�:����ۂYAm��:��D�0�R�-n�ȩ�ⲻ2mI�WkH=V%�]�2r�c#��X��٧�\h��b~�rѡ����x9/l�ә�����a�gt3���7��)1(��t���H�~kl0�)8�1o<�ǫo����+z�;�\�x1P��S�ْ.��̆P�
�p�G.�'��}�w��o	�;��$68�ᓋ�T�2���sg;��=p������!�y����f)]��+�*�+��=�.h�g��8i��U�7v�Ճ8�V�J��ݘ]h�6u]U�� �
J�]�w�'n�愙���G3w8�
�v�A�#���JA�`dY�ȪY�f�n��z�JY�f��]����*�P��˸H�v)�4�����[�� 1�Fu\�����m���:Ǒ�_%މ�cuux�u�uJN�=��j|�;��:a�������E#��
����������L�*�c��\������'7�M{K�OW�Ⱦ�q�ӻi���HAu�`%ԝ��epd��7EPj�C�2�mg��<������]��ك�u�9<ʓ�a����:���=~Rjכ�Z��';���N�z�gT�Z7��s/`���t����v#�(�3���fWw�A6�|�Ən^k|w�k�(���{jg�zk]�o�'�2� zP��*������rcU�^OH-)�e8�<����悭kcՕs�#y�ycl!Lзv-fB��x������G�>�&N�,\ҤW���Ȟ�I��`���x4p�>ոc�s�z�$��oݙ���¤�J�Ug���"�8�(�M:�GAk�@橏^��`���Ef�V1U%)�Y@��3J���h��7�i���Z6ugA��b�݊�
���5{ӏs����?5�e���TLɷA7���_K%{7�g��N@��l6��Rg�e-qA�Uю������}3���J����O�"B,��]���7��)���i����[���|�I�8�hl�j{t�W�>1!� 1M�~oVh���!����-���{�������쮮(��|!]�'L0j;ݏ2v�0n��-�Lo��P9.�3���r��c7��?�P��|	���߰�������_2��đ�����"^�u�ںg��)X���-j-Tj�o\�lq�g��
OYS�*vOc҂��U!O��!�g�0hO��KQ%�z��_1(�{Լ
u��]�c�rC=�;�8n�D���ՙ»�{_BX���q�y�ۨO�1_k0���JE�<��Dq�{�J��'�U�ק-�9��V�Ļv�k��6�ts��}n�K�T�nL҄d�ގ��2n�����"�͗Q�����i<��}5C�HG0l1u�fҖUWRU]�&��5j��*�N�Wt�g������h7"���l_���1�HwuteR�"�6�͞��s�-[�w����ϧ�\�� =���(��O'�t�����gw��]�+�;�� �W��}�1.��❏��:�^�l�t�Nw��S�Ѯ�V�oY��H0EJ�7��N�I��>�Vc�pcU��`�W��-�u��d�����7��ܼѽg.I{B&%�5�>��_.MZ�c�v!������u|��n?=�{�������g&t��ˮ߷�*�X���m�)u��=��7f��}ٝZ�?^�W�՗��ZR����ī�6�\-_��3z�fgg�Om5(�y�VpǴ���l[K���w=������	+I�I$����&���F*�Uۘ4�B�5�����qTPD����<�9�`��2�^�b�iDO`�#2�U[E
�J��fb�AZҧ�*`�Q`��j���N���|\* �VB���%���r�,bڤ�3'9Eye���QQ�2����:y�0*�EQ�PU����Z�.4P�/-��.4RVT����Rq2�r�ÇN�<�^����T�[p8�0�Vs*ԕm3�cJ�3Kx�bULVLC�-:t�z��~���lD�d�Ô;h�q-eyh#��^P�{q�<�l�����
�i{c�0�O�ӧ9zVc�V�,�I�E�WS���PƢx�/�˖&0\[��)�LE/3<�<���iٝ��h�1ŷZp���+)̘(�-�EY�-�ʼ������X��IPR�il�:t�Ӫ���*L��kU��G�m"�(����agJL�m��*�b��ǌ�L���e�q1na���-�8��91q�AeyKy�1�-F�\����yJ��/-`�amY�j\�"�>�3��+�}�{����J�^��v�ϟ)�ݍ�������{�ڼ�#�~	���՜�đHu{�~���� ~�0;/3�����LfX�/#g��7��Ά�?�@:��e�VF��GEC�Fq��tY��x�6���Bs��$c���`F��t�WN�j���mJ�Dm��V�*d�$u�b;���zŠe�)�.���Ue��:�;Hx�Uzs[v��i�>�t�Rc`�~zs�A;���A]w��o׹UYN�g!@��ډ����z� ^#��VD����B��l�e.�S���+�
-�!�E��$p*_2UL���"�ۨ����n�3�5
��j�n��}}��yj}sN�m
x�"��0���HJ��8aPɝtd4�`x��=?^��ڊ��i_�͚�b�յ�����.ѧ8H��i�[+x6F,-&�xÀBq���T!E؎̞�Q�wg��@�Ʀ]f�릪�N��!F���l��IqxJ����M��|���h�b4����d��#�=�Ӂ�sr��nT���x��`�Qz6�"ӫ�RI���uo�����D:���fg��
n�tK=�Շ�������㙽�����"�����Ϋ`ީgK���7*��P�۪����|=�5�ٽf��@����z炀m�u�͎KG*E_<�Y�2�]o7�"���+xe���!�d5!��!l�����h�skc�[����}�t�b�y�ΐ��D"��=Y�{��9���G�xm%����{�?|d���Y��}�h���vM��L�����[�s�3zDH�`�b9s���;������>|6�I[EQBS�1r2����8��k��:*+��N���5J{օ��r�Y�Y`#s�{A�:Clg1��/E�8�^i�����t4k$�sf} �V'���M� }�h�0��?+ѧ3wr���V�c�vHԁV�l�P��[j�\s�=��������cF7[�$�}|-[��l�v>/�<��E\�x^�OA������O��E\��kN��%�'�������X�'N<)���=e�rUf|����@M,�}����7(��E<�قN��5O���[��è*ˑT�IZ�,g\����\���4���{�{�;�|��;����w��A� ���t�:w�߈�G���+b�;��u�8��/�=}٨�U��`!2�M�g�Te{�e����r&c�o�p��äml�Yt�6Y�*��a{3m.M��5��.1d�Gcs�B;�ע�'�7 ����
Q�8��V'�$���K娙�}���z
�1����]>����Wu�[�"�*O�f�&f�	��g��wTⷍ�y���'EH������g'x�:kJ3�6���m�j��!���t�#V�r t�9�)��sD��It҆��3�v{����f���=ݫ�ǰ�lǀ6� �� rϣ��ݷ)ݲ�z�b���Zos'i�y{�4�����l�vJ���8���=/��w6�0k2zޙ���jrMvt�q�Oi)�ܻ<]����n40���x�Zk1�޽yB�*O�.��o��N��7��}�k�RU{L1�����vz9��c�F�Ar�a+$0�S�fV�˨1յ�Ǻ�A��|W8f��|�m�Z�ݎ�R��8�h����ϳ��� ��wt艐���ݥq���ا7��EJq�A��#�9m�ʇ�(W�(�����1�ī�ƋH��VR�Ʀ���n�;A�w�Tqsٍ��,i]n�tiKR`��ٍb���j��#f��"�h��� �h7>yz���v@Yl�������fi:Y;i|��ױï�-�vL�F�toxC��g����rJ��m�R��p`�j���p�s<#��@�OB����������f �Ԅ����@��.��ɻ�M��㦼�7�	(�=�嶫�ȇ#Cz��ٵ\�͕�7����z�ΑÒ�+����YV�GWa �"@+�VJ����g��:f����f�E��èvW��Uzf��mrY]�6����VT�ߴ*�_L%g�{�wg4���s��7a�x;��GrWO=���MW��b��.��tr�S7X���P�>�7��Q��$B�|#mmsr1w.N�Ta3Y,Kֻ�{^9P))���jw-Ԏ̚i!nB5��K�k�˫�:���r69�I_���(�>m�ƺs�݁@�NΟ�˦qw*�S)���/�{�;hm�k��4rϧ����/�ߎ����p�w״rB�}�Z�e73h�o��g��ױvO7�{.��y��rf)@�~)2�l��_c{V���+4qraP���x5�ٞ�7:5�d�g/��)u�&��y{ѻf+�؞+����\o]\ۥ��.�nC�۷}�Gz�6n�t�	L.��hW]�XK0iX��-{��.�������g�~<2��zi�{���o>;��`�&l�U��Tw
�y��^��������NU�`���m��`�H��M��J��ݍ=Åt��l�5����Irxt�p�����Q��1(��,(���DE�h��6����!����+!tV.����2O�1�p�Zi	��O5���:��꘢ �U���<���5�#�}�#݂zF�s#���\�գR�*g�2(�}A��3X�����z�c�NA�{�=*���S���W����/^��s'׽�.5x]3���)5=W������*#fX�w�#����Q�m߷�2�K�^��t{�!&��s1ӗ�j+Pd�"dl+K��-��*s���t�Y�[�|��s޷���OV��a������q��!�I���c^�Z.�7�a���v#��t�N�s�������q���R/сv�u�(�r�`�9r�0I�WR�s��]��z(��������� �����M��j��|�8�yjni��9~��s�bċDB�~뫶�z���w[�ޯ	�6�y%K�S� �H�4���8AdɵN�0C�=6�di�UŚ"\3���Ԅ�u�A`��z�J��V���@��M��Z�f�۝��j��%_rh�Co��It�l���S��	�?��Qqջ�z���-��
;"x(�ee��f�%|��\�ov$&�ɖ��ָ�OwF�f�C8O�� }�eF���q0LY�_ #8:�onF��of���]��IIq}�	���`�-h��H���a�ѻ͍ӕ	9˴������w\x� ���gCz�p�����θ�!��-�d�>�=�u&C�Z�o%���Xbr�	Nf.GR}�o��L�jw��Ca�Z��F�����u�+��ث�40�/��d@2���&2gε�VmG4\tDHK8����}��LΡ	�&v7�[��Zz�̯ߙ"�����'��!���o(�Y��Q�v�g}��%���v�yd�jE��L���a���-6�«��uR�E��:�0���^�}}���ܱ���a�8(dn"��h� J>�^�����+D�a�^��cF��>��+����zg�>�-��������WA"}�$#:`�#GÖl<+��(K5���8h�l5Ȱف�L�W�5|�c�n5��;)�r<C�B��%�W&�r'���8l�k������7q� �K�e)ا3��c�B�T��ghx�UY���Q�6�/O�؄�F�G[6Vz���CŌ�8�[��m7�Ny�G���}S1w���.Ae�I�8���ˉr5N"��br�q^v�\�#���bTx{���j�Y̆%�R��ʄ."��-���N6�o�{c�
�c��Lwg�bS��;k%���N���m�v�"m���;�f޾����8�����V�����)�H��Ε�=���8[�v��~��G��N�vx�]@�4%�m�\!l�>�m�įlk���ee��)a�Rt9v$)n]����vc�Z�_��׽5�gk�]Y�)Y��Iˑi�PŞ��h��so�(q�0��;G�f#s�L���*����o!����%s/-Z�/�}��oe�H�Q/����G#�w�a�����֙�������o��{W��+�Pai�_"ζO�J���_��-��]C�g뾭�W�`: D#�g�݊f�kϺ�S^+�v>gmu	�u\�􌊪˜ı���'[O\F��s�\�В��0�i��,���s�I�� Tv�]f�j�����Q�;�oѷ�e`���������pѕM(�sb����6�l������������H쌛丹���)������v���He�
���g�A�t49�vu\��w��n��"�J�s|&���"�i.4�n��q�:$���d3������|�y����2�=d��_9���r�[� '��#���]�� �X#"���on����2��i������{��*�Ee��C���8�A��ް�(^\,�|94��wYvln���(��c<�
�����=Q��r^�� �ԓG}#_��ze��E˾"���i�0�����J�F�۔'9�b�u�foF�ڌ(�]7e���K�^�I$�e0�]�T�J�Iu+o�+X��l�F�YW��w�5�m�!�V�i��T��KY{�X4-�tg��:]��lǌx��ި��1���u�#9
�����GFN��:����}�.z>]����۹��V���=���x�wo y9#2T���'���e1;QWt.�gy��dw�z�I誠�jw�GfH��H[�W.h�#�e����%zu��ٮI�u	(�s	)q�2�7�'������˪�ݮ6�^�M�p���7iB���t�Zeq�����ӱ�,������4Fwf��s���!��e��B��;�{�Z34�x
딍(�qv-�4�ȩ��p��t��kd�; >��\�&Iڳ�b�W��ӈ��Φu-�x����v�ԩ¤.��b*i��0�Zk�t��R7#c�G+(�!�vn����I{�?[dOl�=�� J�[#z[�|�9���8ˍ�t�\�����p����v��X	ES#9K�{�{ۗ�hѰ�=�Î��O>�T��F�w����7!ύ�v쥈�e[;7���fUv��H�O9��E�>�a�qjW����&F.�j�l7��U;�FY�!��/�h�{��:������,��u�R�>Vݼ�;�gb$�����T�U�i�
o�.���}�����F�$ "h�zQV���$�Ճ�b �<�i�-��S�5�vU�wu�f!o��a�WTU�F�[b�C�p�D���z-�b��\��ޖ绘`����8�y}�L�"XY��I��� ^=g`kZ�f�혧���2�޹�����/k�tS��P�A�Z�6(ߪ��n��Ŷ>���ՙÿ_#� 	�e���d$q��́sNdl��)�"�1��ud���Xq�y���w�~{�=Y���U)�;5u4�E5��ٽ�l�vUD��L8ܶS�#ѹ�o�G����#A"����ٻ�k�
�i��9��)�,��:�:'��4'R�^W��H'��f��C�ǽ�6ʾ�C;f�.u9�6�<`nK��B�e���/͞K������S�9��kGVgs�_u��;}!�k�O�7��ss������ �F����K��O�S1�C��_�4�sfH;���2�U�{G�=��RYJh�������a內��N00p^���;�Gs��B�w�������htz<N���L�`�$y���F
�87����J)؍��0!ڼ7nk؅	�ҧ�o��WIĬf��*��E�ҕ2���͵yQG �aԦU8
��{^Vf�a�:[f9�#8����{p�%�$�GXu�n�u�vI�l|��Z�+�HX]N"��{���'4ӻ�w��H���R����E��`S�ݒ��D��WFx�:�=:�,̄q�9�*��%����3:�kR�Ъ;�w�s@هs`��2!x.��β{r�6Y� U�+��<ы�X>��ޓӶkw��3|J^�qy�T�멑ٵ.�;�C{e�)��������Sr��8��^Mλ����g���|nx�<fY��A�]R��ψ1`âUǒ7{QPu�N8���wqe��������3�]��|;؞�}�g]�����޽�N]��R�Ȅ�u�  ol\��.C����5v%�:-�����\�	x;~���ugUԒ�5�w=�i����W�x���=X�������n����K8�v�YK��bD���e��wp���n6�U-*�U��<�<P`7$wM޸��s�=���̀"����
���ym2��+lf]���tg����5�eRd� �)M�f�/��\�a�<2yӣ�9ޙ�����E�x�4�u-��;�z��D��\r����s���6�ns��cI}p�����tiܭA��w�����\�:���K����V*Ʉ!;H�����ZA���atnu���[���=X#XWQo��7M��۹�}�ɇ��fU��${;Fk��;V�̈́���<a0D������:�M�l70#�s7|nVR�Pg�K#����~hC�řo�>Ӎ��y��m�Ȼ	�px,�v�����W�����1�iD'xVbX�;+���}F��x��.��m]v6�V���0�4�ӥbk�F8j������F���ɪ���l��]*��M����;�Զ�wl[Ӓ�\Ӷ4�r<� �eP�b.��A�W�+7qb��ʁ�
n��e�d���s�8���E���F�*�s�,d��Q�_p�1���Sv�)���è�R�2.:�����j�&�bo-Ku-G����-;��kzS��N����ue������.+$P��e��Eօ�c�6�G�i���nl�L���ƙ�-�UE64q�yc�Ю'7:���a�l�6�,͢�+q_5��NwPMZa���1i���Y���zuH�ᔣ���7�nk�n�^���_8e�q��˾Gf�5u^D��v�\����u�4&8x*{�/ x���H/:TX�BI3R�����}y} r��L[�~����og7����Ջs�a!����D�����;cʴt��*�cws4�/k�8�4┱��mN��ۥN�5L�%�L��;�^`|�L����$m �r@�B1 �ߗ�2 Dxa�%��2P�>Y���y���@PaQ�����2��e���#�?��5�u~�D�"Z+Q�e�� ��ae��p�&5Y�j,�U���x�LJ׎1DÇ��:p�{�Y��s�.8aLώ�p�V֮Z6����V\n0.)r��j��r奏��
SON�N�Ԩ-h�(.aLd�Tʼ[E�E�\
�f�>�d�W��1G��)��ӧ�^�#���X��X˖��˂�=Nex�[33.Z�Z��8�\�`^��9V+*�<�y|�aL===:w���4�LJ��Ӵ�d��ne�yq2�qN[��8��LO㊂���F�b�i��8�����*W�^ڜ���*����,8ʅ�����fX�q-��g��jc�0��;:u�\ne�q�.w�TR���EY�^Uċĩ3�qE-��'0��EU���b�)çN�{�0�-q-�Ŵ**�iYOo2��m�`��lY�TV"
g9��S��<h�,�OON�'�{��PP�%[K�
*)ļ�P�m)Į62�pUf}�8�̤TI�Q�%�2�2�*�2�X*ɖ��L�+R�\�Cc^m1yE�Wǃ0E*�o3;m��g���w?S��`91.
�=����}�v���z�����\�r\V�TvL���!ݵl�����m70�\"�EaL����߀�2_ut�;M����G�?;+�H���Fl�l0��,���ʩ��u=oj�9�x�Ha�l�H����8�ɵC��[�,�m0����ί�Vf�a�n�!��z��n렷��=�(Jq��(��=�x�z3w"��Ļ7��$��� }+�6���n;�n�tyNW&$�^��s����v�[�+΁0�e¹��������n����C=��Ռ�b��kG턅��6�m���8wFE������/o��0�{+̚�����]AtwkG�)":�B�����"�M3���F��\��gl�93hr�+P�_+)k˛�g��'�5��9E��9��SM��":�8��;[� �C�&����'����;����jc{�gkb9���&��k����Y^��'���^=yz�	5*j��Y1�#���V����U�=qb�%|x���[~䱔J=��O�ZXwtY"�E��VƠ��8p���)uV"x��5B�H$�H!/�F�J���;��+�kGT����I���]Ŋ�}�V�����w����+����B�\6���εۺ��Ǹ�~vg�u=p��?AB�TP�n�Y����[#]�r�t�V�C�UV��'��@�nן�����}Ӯ}�,�W��1Ӛ�B$*�b#�s�]#[%�nP.��u�'6�(���*�EU>��u�`@7���=Cj��������j��7���E���}=���N��{�����A�Cv ��p��2*����(�4|��(�Ɨ+�}�k['ݒ�w7Cm�z�5�;��w�Pט������Mr�޷Z�Е�+��.�ȬYl��Zk%�"�-�xS��0·\f#����U�����*���O���gՃR�:��3@��3��5@#�	�p쑸i+�̵n}䎻�q�q������}pZ�};�B�~�h���8!=#��u�fB����Ŵʯqn��kh�:����o��n�5c��'���v� ����H�G��B�(_'�[n�o�|W�$�W���j�mFš�^�}�~�oR A����P����r�F5����tM�[כ�ޫU]༂��5����Lӎ�U!�1��rﶞ�ˬz�j����Z��Ѫ������84�Op�<y�g�M�G����g���}*���~��������^Y��Ê" =��ڡ�ׄ�3b��Wv]����X�lA�?=�{�*�[՗b#���UБ���v9�k�u�GC������[ʟW��=���SUGH�
�<��+�!m�*�*+ʫ�޺�^��~���a6A�>������[ �-M�V�X���Z42W4M�i�8��ř���u���� ٓB��G_:%�ḱ�Pna �V�z�-�=��f��͎��:�p�$E�������)�{�#�-����F��D��Y���h�7�KK�;�x	%�n��C'4�r�dG���n�g+�k�>H�����6Ԫ�/�U�W�FF.mG"̤�5wW��:�������᫂��L.��=]�Uz��9�_�w��䓁�>̽�(�"t9T6Tr	$靸
��cZ_>�JҪ�c|3\�*�N���.������_`��|�lE�^"�y_6O��}q��|_צ��uT�ێ�U�;kM��}��ȱ���Z��cYS��:����Yr�� #.㭰�o�t/^â�^�l���z���-����2L��"�Y^�+64T�&�X�����I'�F~o�s����r<�\t��b�O�ݢ�[�\�k�p|k`����}ѹ>ӧk�u+��ږ��|�9���ߏ�Mr�v�NH�a˩"���ޑ���~�=�=��{U
�������aׁ�<4 V�v	5�L�:�G`�fd��_�GQ�G��	+_�+��2��6����������#��x/m9n�hP�36��wG����TC&���@B�=%>����^d^�_nKZ�w�=r��{fk�<��Y�` Kׁ�C���Mw�c�m�*�jxamwa2�&k8aevv�HWfR�cH��>���¾����c2���md��^4���s��Ap�cG%bqJ����)z~�$�Ϸ����5�\b�LɌKt��6c�c��7���,b[~��]AMw
�Gr�k�u�
n�Ꞛ����.�E-�2�&Y��)�a�3N�2��ɞ�3��޾�c�r���䝾r��݇��͵�ј�=B�se�̾09�i��r����g�x��rF��~���='�Y'o���Bo�O��R4��%"!M�L��~y)��e-��w�]�.���)��ǆ:���m���IYxJ��(�v;�A�튓�ǭ���Rog�>_�$k8����������͎K[��l��Fs���9�r|{���䉶#���֟��5�~��~�N	���ט�9�q��̿��q��:�$�(A�3[a�t1A��|�rf�w�Z#��I�s������M�GN�{�/4�]��zG�0^:�x��m��O;��>���߅�����M�����V�H����.��S였����_h�O�[��)���k�Gs��ˌ΀ ����f�w)�y�Լ�[�|>�G�+�u+Iv��'����@�N��FlȀ�ax�����L	��y9g��Y�:��͘R�]"��������+/u�%���[h����Uҭ�Ș�PrZ�= ��Od�]�Fė�=����Ԧ�"�Y����A��-�)L�)qܓ��rQdg"����أsJ�w���+�;O	�d�wP��U*;��X�TE�����Ɩz2�Pv�ytji���8��ȡn�n9�i�f��Ǵ�� Ɯb+ôa��P���"@"��$ےq5��SDM���U��K��WF$�]@�B|�r&�Ԏ�u;
<�z�xI^Db���/�q�&�L�U�p�!=ht�h�(�bORؔ��f)�ƪ̭�:b�a�"jp��"-���x��hR�H㶨=���-m%���翪c�-��	�^>���+xZ�S�cht
�9H�"n��y������`���;�u�{�n�����EO��b蚶"de�t����E�l�kp��w��nS=��4�UA���T(����ʰ�!��6����X�U��-�F�s�3�X�\k^}�N����-��6� �6X�铦/m��ŭ&�u����ѶD�����TP�I�+O���;%O��?gM��w������lѼ ���C�T"<z}ӓ��fk����������Y�Zn'i�b�?�|0�v�f��xy��Ly0��`C�(j��ߟer�����w�DAYcM��l�Ϯ�w��ϑ���p����8{PǢ�F$����-ǯn�>Mz��'5zo��F��ɻ�{��dYѷǖ=�"��뜯úep������G��n#�7���� ް��~sA�i�j3_���p9�������!��p��ہ�is��ͯ���3�s��vwrܪ�c�$d��,>ϧ�����..��OFƼNU�!�8O��-�#�t��zA�:Ǝg()�J��y�ᵫj�y�޶q,���N����̍1��4���tQ��1�!��觖��n[w]����+`<r��F��E��ox��UH"�z�.���2�OJ��MVWk���O�P��E+v�E\�e�,$u�V�y=(2�����߷��� ���Kh���U=Bf�W�"�.KS���}a��]���~��Ob�@q�i=P*%�U��+�a�$ז�;��vL=I�ܿ )ԭ�ry���Ir7+��ɳ&��s:%�Z�<��B���TBȸhm�P�6�|���	��I^Gb��:fnt�v1�r�Xݯr�%o�s�{�g����>���p�z�!W�%�˻���g)�[��9K)�\)m���K�X��p�ب�\��kS=1�p�ގ����i��]
�,()��9���oy�^�U:�y��1{]$KP��$0�����7�-��fw�����H���E�$փp*Gm�,lt{6
6=ΒW��2�m���f�������c���;����T_��G���2����4���㬍�g)�U<��M�nކ�fv@a�_�#��vD���Ԫ�o:}j�����l����n�1u	B���)��(0�����ޡT���9�h=m������˶Ve�K&IV��na�q��(T�A���y��k���zq6��ar�����4��{�\���F�St{Y��qg
�ݬ����\NÈSW�n�O�t�."gx��D�ct�3�&�����_D��P��_P��z��a&��I#�8��h���v��v��o�>-�p��f�V���}�+�����ˏ���&�47m�\#1���w��3_|f�����<���=��]y��{;�V��ӼG��<Mޮ�xO��]�f,���HI ��� �؂�{R��7�32Փ���d��u�����*��.��d�B=���;���̫ܻ��C��񻬪�*�i��e��蓐�	�$L8R��}���h�\$�����{��և�kB�S�y��A��v��sҋ�4���;�;��6���7���)�!�P���r}Ԅ�gd�>�i�6d�U�ɮaY��@@��ye�]����SsNv��ss�6����&w7�A���ތ��aHɴ+
Nϱ��Й�0QL��-��p���d8n��7 >��t�"t6}�W`�+����KD�\���o�w�ڶk�����i���C2�u���d�ޔ����0o�G�O;�gQ��?_Ht�X�EmzppS�P:ˣ��_���K%�V���ߡ�g��}A�/�kt�,~Y��B����le*awݓ}�J��C	��B���Fp9���{�ϓ�{��:w\+�}@�/#_�]�kwm^��!��ߺF�.�b�*�����ā�Qk�P7��u4O���2L3�2���U��A�J�s��k��l&���d�~c!Z�o3��a�A7��ZP�v�KRϢ8�Aunnwvb`��8}�]�1���P��ǢO���2E�s����7zO��+��;��\Ļ[��.3b�� ���x8׮�*q���r���|��x0��Ʈȍ]����"fxJs1tݱWC��dסo������S���7܃�JD�f����[����f�H�ĂΞ3�y���پ���;��!}��]�hK���ϗ���{��$��J���T�
x+W�������;�#o
���y,�n:z��gEi��Ȩ�l&ʉQH1�[�L�6�;��`$���R�^K��ۺt�G*�QJUO�Q�Od$KǍ����O,������eD��F47�;0k�@j�52��ܸ�hv�h�GZsiE�TM��j�c_i������,��9D_0i�d+��;��2n�Y��|<�_)��S~s*㗿�o&�CM�U�x��ԭ��̈́
��[��}n�cٱ�ٷ�H�.y	չ���[<�9��"��q���
	/�C�M������p]b����]�� mB�V���쒯dЪZQѻ�g�eM���ӫ"�Lãu���t<}I&?9V�����Ye���Cj�]�a�y��Qڃ.�/��(�̐��uV�k�,��E�E�����w�=���+�Xe��w�]�d�`�aza��Q.��}=�w���Lz\�0�]��Mkg����m�aZ��j�3ǰy��uA�lϠ�Ck�%��4�g�{;^����<��w����R���I��wYw ���oZ�7�g��O,R��t\�^��2�^�o+� �	�5�{8s�ՋT�B��9����G���F��H{��v�*��%�g�~��^�}3{��7v�	אak^��Iº_9�I;fn�ٞ}W�@c�8�����pmr!�ĦSK�&�1f���&6�ݽ�@va*x��-������!�yt��N�<O�t�n�F�������m�:��7��z�N�Y'-\�r	k����*�a�rK:uNO6T�9�a�4�4-�5���Tރ�f��8�����S���T-��y]�����r�9i��+k�|<�v�:��'�/�5Қs}��J~�>Ή��AC�Ǥ�~$�g�e^��ۉK8Č^V�l�nXt:<:uZ�~/��2c�����T՘\��l�i#�v��c��3}���sֱ�1����2I�q���;R���?D0�)�ݥ�����B<�~lV����j���A��qlgn�L�S�s�<�L���tB�I�B1y���J�f@�;l�G45�,ۓ���V1�: ��xZ�Zw�R4���Z"�"L?��M�����Ǹ��C#P����!Hs���.�s��Ϭ�`w���r�����$�t�S�vJ-Ci����:�yzzq�P��,�;�%�s����^;1ž���w�>>8M ��w��3����)����o�n]܏R��}WY����ۍ!M�$&ZE�	�(��p�L��Âz߲��j�i�����&��W���^���D��u��L��B����,_�K�yޑq"��}v�]&�I��)����{Ī�:��ȶj,��y��f���=�����6o����>��;�KW�NU�Fu��g\z+�][!CP�r�!G
/���}T�ѪԪ�vZ3�69��u��S{��$�~�>z�_+
ss=�ٸ�8AYfpJv�Wdn܏���Od���`��e��0�"1�F���7������pŌ&�y����D�8����J�ɽ���Fβ :-}U��W�;S6�O,i&R	������q��ޗ���oJ~TyNx�af�xkG�c�GV���}��������vbc�����Y��T����ziSΝv�f;��OG+������BP�郅&��
�5��{ޤy�]+p��Z,�+1Lۼ};r��YjC"��͵R�Z!!�H�@���K�v�����e��dX���R(�
�	N��N�i���-��W1đq�-��L�1�1�*��P�X�DD����N�aܳ��Xň�en\gԢ9h����ԩ'˗L0A8p������uR��-�}�y�VV2��PZ�q�����ʖ߇
"N1b�)O4�t�LȎ5�3,�Z�6йjc*J�A��"L����m��"�����NŞ�����+�FL��q�R,�V���T��*����m̡�==:v
w��jT��h�j.3rܪT�VT�-��XT1+���V&:t��%�e�im��T�8�,c��
ќK��aj�b2��*a��:t�Z��c"��D쑗�Y<x��̫D*y˜��C2ت��ҢQk19���¸4��>�Ɯ`�e�a�k��9�i����j��J̪X�kŰ�k�i2E
�"�')���\�1��O�\9c��}uJŎˇ������B�}��qA%���y�7�x'���H�m��S� �g��}�s{�Xv�jო�&�x�1�$6��:�O��xҒ�uƆ���]^=�f=틌���V�x�X1u�p���ܘ"F�؅;f�3#IQ@q����xZ���B��f�h��{l�6f��"�_C�5��>S腻��d
�֒�wJv��z:6c�����;���{��׍p�wW�q����zߺ�m,6�����G*��t�ݼ��Mb� �oK���<9�ހ�#"6��f�l�f��+�1e�\�_�+R����7��=&�:$E�H��=���
��q�F[&k��3H7���jT�j^��"���;*�7d�1��>�y�F�k����h�֛�xk�8��1�h����	K�W�-���F���g�<�E����p�&}�9ݝ��g)�A�<.�<�7�E�to1�����16�5�|]Up��[w��r�;��)�76��������5˺2�y�#�<�����:BuIom|�.|�}%���}�u�kp]�[ZtPC�6;� ^zY9���n����Q��IUGrt�W"���}��6��KNALٷ�ѳAMq��Ks�䢅�����!��1dŮˎ�GWa��Y#&]����bFn�
�{=ʜ�6�8H�>�/ܱO���)2�Ϲf�H�����9��jM�ZA�54�p��0<S�[�1-���4�N��s"m%$��!g$xe
W+��̞�x�{�m�Vjq�A�î��}���cx@��gg]$K:E��W�ݭ-�ճE��x�y��3{��r���Y"�8(�n��a f�G�$�t���nl��=��9�s��9W�p|ƬB��C�@r���F��2��z�����ebΫU� �t-���g��,�,lv�O�c��d��!wY��Ĩw<���<֨��d����{D��p����K��B >��	@32�{.��6V���d:�9ZO%{�*V�{,,F�#jo��bl��Y�)'���6�MYOH�tڞ���jiuI�^�i��o!+X�ҺР�T�zXPeB��;a�{K�w(�s�f�8g�]�X��S��x�j5�\��nM6td�j�{��x\u��*R��cN��x�w2�bǣ~�"�m	Q�q���{k�Y��X"E;�3�r��qI�`��Ӫ�=ԬJ�[#gݢߧ���t�TU<pȫ�9z/���"9��7ܨv�h2�շ�Q{۝���ڜqp\�vB�Q�CX�V�c3�@J��u$G3�&Cv�y�1B��M����ó��՚�ւD�!24Z���U�̀����qU���C�;=�Š������E9�4x���"�����I<Tv�9�UQ(��e�]#�H=��vD��&�^�痠6ǨwG�K�W	Yw��j�op:��fb箠ҖX;�^Y�)v4��1Pʵ��u�ׄC#�:�	�����z�"Ly�l��/�`g����yb��r���򭉑?bf�7��[����]1��$��L�7N�������3�Ö�[��K�auq)@���6�&{����{z&����7@�g�Dd�J<�lD��3�b�E��*��L�<$6nɽ��ٸg4*�{n��Fw�t�+�$��z���OU�G�ث]S��]VAc�~:S�s��C�����)����6�R��}8]Yв�w����vDQP���^��*�[�w���\��{�����t�s'9&���3|���8ٷ���$�\�}-t�������Z{�太���~4qq}s����O&Vn��D6�An���{b�x���2B��Y��mrב�G��L���O��<,tw��y��X�|ԇi��Þ3u��WWj��������\e��������Mg\�ot𩁰�2�{�8[�f����>~�5�%{i"jaT���uY�dYݾ֞y�ԟ�|�s�0��q�Ԩ�݊�X���x_J �U}�i{���D��c �u�կ��2z�8�����ב�?e�|;��ښ�H��s�_Oڤ�n�&:N��k�a�]���<���*�<T�ȩ4�w}�*�9��G���#y�'����c�3���?���qڬՒ�H;��݃�GiuGj*�׶"޺'�7���?��Q/��S�ih���o���Y����e�OӻYe{2M�=x�9C�U��œ��0�>�=�T�Jݽ�ݙ[�=ɼ`��.ۧ�\+���kx<�$v�n������jW�.wi9:v�����w�Lٞ���~��K΋j.y3�ޚ�'LT�7ÇDP��Uf�H����Z��u���6�x��4� de�M�k[���2�ƪ�ߦQC����v�(L+&�#�G���Y[��UU�m}�훵;yK��\ө����bڳ�Ds�^޵�egpW�c7���J �)�:0fV�u"��@�ƪT�b��:ʭ�7�s��7CS�10�X���8�Uh��>�\��/ ����;�b,���=v�v��p�4�7����<{�:�� T�+H=�@l�*�Ay�R};����w���̑�6�J���ZJ��K���ֵ���ś��3����o��J�� @��oO�D����f=�QZ�ؒ�\�d=�=�����\��g��E�s���{�2��s#N��F�eI�~R*[���w��q�try��AY�S����7���oC����ms��h�M����0#����o\���BZ�J����I�1����/a8�_;8�D߯��M�
0	 D �IE��&7��fV�Jo��40�6�E��v>�׵G���U��y��/�z�|"{{�3@�����5���j���bz;~�+����q�J��:�wzF��=Uwol�̸�3d�&۔��BB1|v�(�v�rc�	��ё�Ǻ�c1��zo�*m���`5C9��C����l���c�w3�<�㢉ʅf�Nr����� ��{-fa�PQ[�摡y:�z(o{�	��"i��\[��Q����ZW��n�hoXP�v��Ŋ�XH�������۳�gl�A�AcrN�u:�ł�Ą��7&p�P����TF�փ�^�/���aڃ�v˰=T�潅�+�pA����m��ػ���2�śZ�o
���Ђ�䌛2j���tKצ�)���ƺE�u�Zc2kC$o9<�hm�p�)�*%!�b"ӇMe�o<c<%:��uM���B�JDL�Am����3`�~�I+�=�O��S�N6�QSHIvqӉ�o-�f��l�W���<�HS���ih�bH��8��f�v�vl� �][������[��t�|8��N�Z4��X+9���ʳw\�����Ze����f��Z�r���l�������j�t�BK�ˑ��T��A!����D&!*$~ܓs���=�Q��lLo%��nX�F1\�n������]%'W�M�9��9�����m�{�V}��<�'g����1Q�~�кY�T��U ��Z7l�W�ë��W�oܥz�Ewp;Γz��k������r]���f"��N��#8f�Gm��<�gq�[���]L$n0�v��hZ�s��l)�������
"Q��J�x��ռ{�\�ߺ��n���OWx�f��7�>��<��c�D�q�ԍ]9Au�8����u�s	����\ǥK���+��gA6�l�\�E�dx^��o�S!�s)��K���n�v����S�p�����f�o���M1s��P��ޥR�m!�v�<tG�s4f��Ĵ�:)�Qt�(|<���¯�}���c��m2f���i���K0�;����ܚ�I���W̡C����b3)�k���kO7�w�!�9>����/"6p�|4����pۡQ2��.���9u#�$(�B���p�f��(lӆ0����.t^��F&����}zqq���{�cqe��+#�b���T������y�n'ʜ�s�(o�)Y~�����[e�4�0�z=�7-��Z�T���;xc����vϝB��J�d{8�Y�%K�S��mL��-ݨ9��pFMyԊ�r6�n\����]̂��d��s�0�5qT+��}΅J7�6UPa�ݳl�\y$2}��b0U��f%><�l�����vF��҅����'+��A�A��H�p�T���Nfܝ�y�F�-�::Z1��\���+�"���ef�}L�w�i���.N=�]ϩ����	�ƹw��Cم�}�d�O�V���]�Q+��0pm�����xs�x�����C�'[��Q��GK�iٱ�1	x�����P��o{'W#�_�\�5�2���a�<�oLF-�V����g$Mfnʅ��A���z:�TO��~�㼆@@�12���ZδS6����|s�O]�f����q�}{25+9�������+�{��Ҵ�;�b��Fb���QtN�$������9���>|w�{��g����r�������E2>B��:_b�����+��^j�T7�"u]�K0ND�8��5�{���!��d������ާ��݊H������g��b�B��4���ّ\�k���uc��B	����>����y��z7�OgPg���C��x`G�,�C�(Ut��z;���(���/mF��5hl$<�Q�����b��d1h����s�}q���+`:���W&�_�u�#4�*�Љ@��)��/>��l���u_�8&�1����\:����T�G/I�܋������yL���Wu�΍���k��>��]caTǬ#FeP��T\d���4,�x�;cs5��C/a�<z��^\Ӕ(Xo8U�u���]�j�	k9��24�g{��\�U�(3#e\���>9w#U��g؜Ҍ�y�Z���n�y�YR̄nwH�H�<b��Y��U>�#.r��W��(ψ]\��m>��S�1��N�<{zJ\ˎ2�%��a^"��qg?]`3_������<*�P)�K]9��H��N8�_�-�v�P�t1�߁t�`�}d�ށ���jλ<3�����9ߌCߵvL�~y6AY���v�eYG�*\�:�]C���rȁ��d��Kh%J�Ra繵��s�'i�7��.W��QӚ_��p�vϣ�lm�*�m<
�TP�K����$2vKgf�ӎGoCi�*G��G�Zk���?�<�"���~e��oyʹ�������W��6J�(��{ڽ�؆��
GH��DF�ƺ�Zd0�CSlN�����Y���ՄoR�p�s�6�>x��oX� h���Ǭ��g_$��kz�9]����=�B�9#$m���ķ F��3xc�;6��l�d:�
�A�f��(�y��q\��G�;Fz��m���V2�� �I��BH���~������MCCt뢑��}f@/�O����s���Ys�wY��m�~�6|F3[�{!��0_3�O4�^u��o
�e[���ޮ������lOϤ:|�}\<l!Fݢ���e��9y)�ʦ�����������&�Pp 3�4=�k"�"���wN��R`�
+.�Q���=d ���G�2d�*+ ��D@F�DH�@� �0qBP��BH H�!  ���<��q"��!B pa ��!H�<� 
AH�$� H  @$� 	  B @�� �d � �    ` (F  �2I$@� �   @ f `�$ ��H   $�0 ��	  �(�  @ H�   �
	 �ID P� E �H ��Q $� �$  $��(�0�)"� f dB""! A�  �
E  �
�� AH�AFI  $��� H!$F�
! ����IFI@(�
F"@F@BD��" �!��C�8�L	BHITT!��VWy�m���d߫���>���#��$q~8�{4/9D��JO/��4�1��V�q����^�V��AEyv�;��$��m4�<'�~C[��� ��o����hL!1k�;��7��7�w��O��!T		 I�H�BH��) Y �a$F H��$! R � d  ��D� �  , ����$�%I � � H � � � � d @ $ � �H  F@ B0 D� � H�$ �	I��D 	 �#!$d#  ���`@@� 2 !�$��0 A�F�F �I�0 $$Y$H2H��"�2H�Id�a#$��'��������_��$ @�@	 $�#f��xi��7q�؅G��Aъ"
+��&�^�M	���ˌ�ڬ/W��ּn-������ �����PAEt�#p�Q�`d��%lm��.��5 (N
6��(�&FFK�,�Q[CY)v���Z;Bw����{��$ ���n�5� ���w�,؀�x����$�!���-�!����MDQZ��a�f8�lG��@_��AEsf�kAVQ��8�幐���
�2�̩�K,������9�>�>���zJ�l����
�N��J���h�*" ֤�V��A!]��fR��5J���흲5�(�@قR�$�Q���$�uӸ���ej�n-�].��.��jX6�-�Mhҫ]e$�[Ji���[5Y�W&ޜ!D�U��4,���m��'�óI�e+bJ�Sf�֚}jIR��USjdm6c5ZJ2S-5��L��E�1fmY�k6�[�ǣ�kSV�mj�l��*�BYem[U��+dŲٳ�.�flհ�Z����4��{ޯ�  �z�>�s{zzz����Z�W���s]� �6�w]��n��v�v��h^�t�Uε�T�w���ۧ]:{�9�=�vh�,�m�{���JuO{ "�J����v�Ic2�kf�Z�iZ�6��  �qv(P�CCCw���
=
/z��
(}C�С�{Ƕ$I}��i�ty:�ݻ�o;mPzn���{+{�Cw[��p讽�OWNN��4׽��;O+�{i����)Q���n�S3b�u�  ��C�ww�)��;e��7���G��{hXz�θT��ӷn��{X4�[nt���)]��=�ow.�ѵ�곹Zݵ���\<���/w��T��x�4��*�1�ͱG��b��9|   c�AF�MA���������:k��h�wX��Q٣��
��)R��,w`U�\���f�vۨ�B����J�TL��ZT�[����^�q��i��   Ϫ�^�;(�AESX���@�f��[EN����@f]��Mn]m]�����H��^��;�ٕ-6�)]Ah�5TkRdmm�mQZ�   ׃��Z�u˕���l�p����魱v�s)�T2�;�\�$h�;W

�n�1*�[��Nv*ܵ\WY��-��fR�YX�f-�Z5�  �{�
�PT��lf�+��룆���m�@Pv�p  �p 4�Հ �p�  7s\P3UtR�5��X�m�W��A�[>   ��  #���h �*�  �+ ��`��&��;�` �а ��p��uہ� -]L-J�fVe3V�U�}a�   �|  s�  ݵ��4�v�  ��Ǡ �  ������s��kNà ۹� 6涵�o{� Y�UkmY"�Pn�  s�ւ�3�  �n� h @t ����а P��  ���� 4�� MM]q� ���R��  Oi������{&M%)SLHL�!��*   ��@�UP L�BaU@  �O�������\��xQ�s��;,�i��:kw�gb������l���[$�K�~���/������ϟ�����m��m�6?ی1��v0����m�lm����&=	�b?�`�:�֞�17f�V��V�R͋��Iu4w��-`��XT �J^��p��6���M��f��j�ShJ�� N^�/����7����������}ccZ++3�v��bg[��۠��{����b��Y�W0[E�0?��;�oC[Z�#�������W���l��SM%��k&�D��&���-v�-��]h[k ��T����6�)�1Xܢ*1+N��[�CY4�U��ں;��7�I�] w��cKV��qT��d��U�X�a�ڛ-X�
�<�dգhn��SY��"��"��D�z��P��&+��#'r���nPxrQ���H�tºJR�8.=u��X4Zϔ���Ѡ��c�Y��f�)t�.'�F_V�p�@Z���C������zi��F�� �)S��ل`��YN�ŧvJ�H�sy2�%�+U��\�Y��B��ܽ׋K��%�W�R��oN�̍�R�I+M�T�)U��֣V�HU��KN2T�X�$�4�6����m��" �eaŲ"­{F�®&�rV�¨�Ȍ�1��F���5ճbʴ@�+7Z ]��wjG��W�* {��*�Tu�W�Ulf`�@N3�k7����!�6$�-�қ4�UO0',�.iSX��."6�� �2�YVnQf-�H�(�����)�ۺy�&b�i ��oVYڲLKh\�I�M�U]%mu����{�l�"��`"��[�'��"�̬ݦİ١�&*H�H7`p�1��������#EV݀���U���6)˛��(V�9�94+�RPT�QHm�%nǍ Tf�v��.��1%��e" 2�W
��cZ`��%�:kkt�p��n���*9��ղ����}�8u>W�h�RthR��C5B�v�z;tkϬ�k2�m�!�Aĵ�SU[�(�]�-�Y/"ۘC��5Owo6������lS��Pgs1��rZ��&e*1i�Z�Ԁ�t��{�}���:1`���1�Q��73^��@Q�������O0�n�	���:��;��-,��U5��w*�)��􇘲��/U�Q�����2�e0���^^ �+h����Z��xv��a�Q�-)�\�v�T-ZͰֺ���}�݋cЪ=˶A�a�kp��{����H-$��Z����y�9SJ��n�������D�a�J�Z�`��2XW��;)Ԏљ7@eiV��;��.D"c	e�����a�����J���lm�G���*���ʙK�����PI�|�4���c�����x�����Nִ�fh�M@F� iLØ1�5��Mv��tM]9�h�3v5�����Zݚ'T�U*��(��Re���f�9w�T&i�hq������Z�Z������9�/~hӆ��`Zu��
��Z�BZ�hN��v�U�ڽ Gvma�K��Y�@���):v-�+c��W���J�_\϶W\5(!�DU���[�S�3 ��'�[�7g[7�=�n�;�K*�"��R����2���`d�xQ���ue��DJ�%+"�I�*�۰��D e�q��C�֬�;���R2hF09��t^e*[��)J�]2ꖉY�A"���J����,�Sx(V�d�`�ܬ�w����*ڈ-�w]L�O)e)rp,��Le�Vljs;F��)#��7�߈q��N�K����b�wA��jB�iZ�[�ݖN��k_�lD`&��cu������zLf7�q^Dɶ20����}��mވ��Tv
P ��J#���J�%��B�Kxf:�K@�t��Koݼn�ڀB�J^ٷ[2�̅�M+��q��=dV�\J��A�vXźtJ�b1���ãK\/@ڱn��� ����)k�[��V0�¼w�#���ֵ͙i��?]��T��*��K:ܙ�h�4�ޑ�$��`ϴ�f5b6V֫��ou���'j�d�7�,ݍ�^��Q��:��^�3Oc�L�N6�5aǙy��&��>˭p��������^!!od�hS�i :ǆT���O��� ߲�;lU�
:�e����iI�x�W�`R]j�:�m��
!�M*�ߚ�Y��l�͑�Ĳ�̀ӳl����!-����م�+r�L����:4����l} ݱC[�a��7G.��`�A[(�f3�bnEI��T��ԃum�(� .����jJgC��b��pJ�hS�z6��hX��7� Ӽ��r%xI[�^h+n�n��XQ2�ۧMn�ѹB�ԱE��f�,e��.����RR,����u�Z�ȩǉ���KIm�D�֞[�z~eg�<�]�h[Bȷ�]�D���Z3H$�n� ��`Fّw/X;�ۇ�ZY'&�ůO"͗���BE�Aa�Y��̦+@ݭՓz
��D���,���ħ�5�b[��p\��q¦��)n�@��8�׆�Ol<Ֆq�Ѷ��O0ST�iQiJ;W��jډۤn5�X��b�V��Q�w����渑¥Լ�v�ֱ�0��
���[QM.��t^�sM!��E=[M���\�a�1as�BJu�2a	5�V�ݏ�49c*��y1v��:�B���]ô��H?i������@8N��k�3��q�G^�V1�z�	���[i�7Zӛ*�?B[�2P��E�tNU�?C� t<��*%qnTz��9+۷��]]�)E��B�)�{F�{�w(W8*�h��uրG��|�1m��(;q��4�K�QǮ��xj�j���̭N�� �t�U��0�X�`+W1�&�ӣa��ܡP	�-�;������1ۨ�����ӕ{�' 	�4vQ���շY�5�h0�3*� =�z�^��Kݓ	[tN���{wN��`1��4+�%]D+ͣ-ډ��)���!��M�f�˨l�](Z�)����H;��Kn�E`�Ƞm�x-�;�gS٣bW�u��;4/	4)'n:yY��52�Ab�62Ʀ,��Yt بKj�����{��Òʚ��N:q�٭Ԙ�]$(mXʷh�
%fnMn��v��A,aش�ں����yn�6���� ��QMT�i*n�lG`Lv7�z]0<:X�'��[sXH��wiw���t+�i;�H-�3�S�^�۬��^Ӹw���Y�W�)l�4�d�z�PA�z�뛏-�w��V:n[��d�
o�n%�v
Z��c
N�U�	�����״���7 �Ȟl,*D:�]�r9�;Z�[��l�c4P{�J�-
O�PG���[�ZE|�v1�f�ʰU9&,2�ƕB6a@�Cpl�gr�л���>\
�y�$��h�Ü� �l4WΓɄ�䣛0pQO�i`:�K4�����VáRX�l�!͗YtB�v-zco$ˎe��t�ŭe��AP�6�q�Ai���s�.�X��C�Q���C>�KEi�����k74#�&v�.�X���!u+�K�Ef�������L
�ֲ9Cي�EX�E��M]�y�i=�!�R��d�^�Y F��'>cpH�lKTӻ4�iұ�5�Z�r�PX��a!���N���� �Go5��xMO��;�32�������ޫܭ��mr��&ӣ)����j�I�H�Ҭ*��t
a[�*��u�����O��ț�`1��i^�\ؖ�d��D�`].5�Z�1�������1�������
Ub�eݝ�B�ߤ��6�%��ԫVńR��V�-��8����+BH�]�"�`B���8��n^kR�DI��-���#����z�5)��1ER��r��c/)ʐt
�צ��Z;�-�x�iǘ�)="��(Vaɭܱ[�T��7^�lXm��%�n�����g6ӫx��6�2R��[#-�O ;lJ�VƖ,(�Y�T�\�	 CF�֒2�9n��x���Iq,��[؎H�3&�j�q�¶�y���<.�e�3m�kщ\�\�{vt�@�v�YD�T�kcqd��ݺ�Pk�^PbR9��BiVY���-�63[�l��K���=�2'Nja�`�6蔥,[v^B�X5�[�ƙ��Z�Tsa�--��i���8�� ,ix4R�s��� f�u���kh�Jk�%���`L:�H����d9��
���p����G72�rH�nΰAđ`�)�����Z!ݭ��a�����y�b���K�]����A��Zk��.�|q�Uv�B¦�$.��8�WF�����9(ҳ֒�b`LX�'��5�d�.'wof�M��Z:KJ�i�\�x�ҕn4���{���.�Gm��*FmJ�^�s+
Wh&56�kU���PF�V�J��U�ɫ�m��'kVV�p�R��V��)�Gn[�n>�.��W��f�M�j��l�!c��֯�sV�D�s��P ��<Ś�6�Vj�`��Śrf���j�E�;tJgC�z�tR�tx�d+��!ݴ'�Y��zl�7i�5�eI�&w�T���lRؾt�l� �g!�e#����nˀ#&SLV]�%�gא�U-����de�[uM^`�v����Y�Z#57��O�:'O�j33u�;��ie���cl�����'x5RN�wZYÐ��,�]�:`!�yVT*�RZ� �I�Z���ȡ������������(�XJ�P.�v-�^�ѓq}v����aqq3*U��xU���$7OV��p^�`u���-�VkY��ۓT; �Z�] ��JpM��=Y�tk�ؚՓU�Z�)):-K�ݷ�Ҧ,��f���Y���GDem��1}�h����B�$ �&77/�任�2�:.�{/r%��04�W�\�M��6����6�dYAaTG
���8򞻇*�Q�B\ۣ��M��-�^2�˵�j
��k�Z++;yjKk��:�%��[����B���(�a'&���/sk1Ղ *��&�a!��JfkuS)�Sv�<ɥd��N�W)��Ц3]a[�����S%��a��ʷf9!�V��H�b��A�^)Z��!MP;Z��V,C,!(����{u�jB0��ĆRmV^h��Ui�yláM�^H��j��.�Β5\˧i�zih{�=�5xY(@"n�X��	c+�D��
a�{ w	X�I�ͽ`:��EGi޹u��9�7t0[�j�^����d^L$L�Q�(Q8��ݬ�~N��w�j��O2[�*"1���O��� �F��䑀��.�Θ�pVh
�L×�o`�ukͺlƍlKL2�iTS�%M�$�حۛ[6�*�f;�@��a�pa�vo�A0uݻE��٘ Ww�n��6�jO�s �N���6�L6pV(7��M�n�[F�ɯOΛ(�[$��<M^'Z���f�ľl��z+t="�ƳK�h�t��hL[��Ve�ڂ�� ��7k(e���B^ލ/1�w��reEi��.�ȝ�z����` ����2լ��
��n;j͚U�m��P�l�l�G�8�3��5g�@̴D����V��E�Kw����sD:A���u`\Gp���4*M�K765+q46�R�[h��i&�]��m�L����R��j�ǐ#�w�"^��dґ�:�Y6�i�Ӗ1�l���-m;'v�H��A�Cri����M⳨L��xɖ�U��f��Q��SP�*]MSwEv݆����(���&� ��cH+���J��ײ=�v+[b����Q�cwm�������pe6�����V��Ґv��zN�Y���D���ki�.Q��Y)����d8��y��M��+[�MkJ%�3��%-���E��4����\K��Z�GK��-�Q�I�L�Y�5:J�k`n���eF˦�4ׄʲ��d6^̺y�⼇Eh3�Z���U�����z(�i�ktAܧ��;��p��ի�sB*�7���Ŋ7����n�|�M^�q�X�z��I�B]���kX(�ˍZv/%å}J�H�ƫ�)e#��q��[�vVὦ\ڱt4g+۝a�
uɘ4��Q��'���)��I�:��z^�ks�&�4,��3H��34k;SC��-*���J˹s.�)������v�RҥRKŁ��n��'�j�E��`|�(���_!ssk	�WZwa��)�6���k@�
xu��xF���2-H'L���V�1�y��q�p�I��lHsS3)��$�՛/�Y���&%�A�A�/���a�/~	`�+[th��lc[���ؘf��f�U��n_��,m�%k	[���i�h��[��x���>#�gi���i��J,}�S�^^��$`K�k
"�S��ӹd�z��"��`�t��^�/^�s+H̃%6V%{N
�"db�����(�eiPV66b��;��2dN�[ݻ��!�QC������"�Y�,�P�,jw;HpI{hm^]kZ��lU�4��J��Rk`MM�X�&n,�r��g�/]�th���79M�Ѳ(>D;�*'Y*i�N�i8���v�V��훑��,n����x�<�]�8��YemX��S���/7	�ۚ)�7�>GU�m��#J=_�Qjj�!����R�Y*�4���f�R��%	PYWQ�rap*Kt�[����ih洝nh��'Na�0a�h�@qb�"����\:�#VI���*LiLS�T�ӫ,Ӏ�Rn�vQ��յ�lE�Fs��7yh��]
뽽�6���]��7Tbj%�b�֛�]=U��S,Ƹ��By���� ��&j:;(To%��t5�b����9��l����u�% ��";6�I�ݔip7fNOD��5ڻ�H$`��wm�CH�OM�:λ��􄷕����i��=���u��)��p�蝃��vk|_SQ�+��C�ؤ�ia���Rr���)�
&�ӭ�I�жr��<���P�h��d���#��Ber�]k#b_[�3SnwS�=׵
 %f�:"��n��P;��cT4�-���7@gc��j�&�j���η������H���2�4�ƥ{Ke�])�I^n����H��ǵc���}��6.��Lc
O�������*>� �kT�����a��<�:����c���ϣ�*y���lvi	�Ww�YeZ+��ƳiI}��5��,na��k7J9L���{���xmX1J�g`t���b���べ[\;�d��:��#�ۍv劤��cU��mڈo���^�+���蚈�F%uզ�d�?)!���9m���Y�ы�F5]Ys"�]�j����Ov�-����1�䶻����Pp+�*q�]Hm�|tG/&�3�����*,[����y�p��J��wr��1E�5�һ)�����E�l^�f�Tk9�b�,kYvT�R��Vn�9P�~۱�ܦIuѡC.np��4JږR6B�혳Gc��=��c����e6��ф+m�z?NW��
���v|w�L�U/M�e���a;��[��E�E�\���Y�.�K[n�{n�_U�P�Q���g�R�%Q��g�oi�vv�l�n�I��1���|�@ؒ���b��7�ҬjD��F��6��m�D�S"�Ф]u�ܗ��9��#%�/1M�*Ѥf\��V����nn]��|wV�����o�ƞ�|Vi�)E�����u*ŧ�d��M����h[,�Gzƈ��]�^�5M�A!9��i�*��ăw���Z]��h�ă��:� �C$���od�� Fq}vE΅�U2�(چ<�ڎ&��cZ�P��:ݠN��U�s*XV(CR����C�;�d1�sth��¶����Eu%�Դ��<#�|:�#&uut�X*9���G�5줒Yt���i���jy]�6��[aoT���"KՉ�oy�V���ߏ�Hp==.��˧I�h�y�a��N��T�]��c�X|����o2��������mw�u� �k�ݮ�D�
<䗵�\�ts�$�
��@�}���5@odeR*ٸ�`ٺC˕��xl=�{�Uj��Ef۱I��0	"��7�K
�14���v	�b�V|����Ћ�/8�Hu��7!�SVqXxV�	�0�J�d��e���XńW8P����{���{'J:u��k�{Lۺ������1l�A�A�})�p�A�րNb���Ǽ��>��k~��1���gj�hڐZ<�����!��I�oG�,-k�މ�b`�CGH�������3��
�I�_r�osE��t���]]�o��q�ڼ��mE�ҹI�ٝ�vGv5g۾ѹ�������1��v�<�v�Ml�:rڹ	�&�W@�/�T��7����u*�O�,����{�����T	�a�=p�=�}K�R����Z»(B����[�e��Wa��lU6���Z�K^��dE��B����D�X����JՂ�%�Wov�X��Nl��s�'pR��������+U�f��]q����	�rG���\F ��8v�F��;�c[��\��E��o]:��_T����TR=:]����ơڂ��h�W��v�³i��2F-��:&@�2��k�S���� �g]n����u�L�X��ҫE�AD���W�Q ޡ�-(%�ǽ�0�����	�:�1�:�HіW0�8u'R�7��gC��Z�Ǖr�:�y_q.ڡ(-Ԕ���_nSӵ�g�����z�[���:�#��D��m,+@��}�ħD*V����%c���Ա����r�ZيY�"���h�$�ݣAX�8p6$�b��S�g,-Z󫶁3�a�(#��H�M��R�)�t����[Y�IsAa�1��k�r�Ƕ�Pv ��rT�W�9ӣ̤��͚%܎t�+����� ��4/CK�*���.�|y�S	ŵ�p�W.RԪ�u-�k/2���kq���k�T+��TiV[4���:T'���Ql����kUI��>�ol�e�Xɪ��#��եܽ-e#�'k�9:�xr�1N�o�e3�r�Vq%���Ģ��ˋ��������z;k�-y,ӧ�����	���	UM�e����L-ɍr{��SN��l^�QĨ�,ق��YB\�uɽ��k�#��!ٳI��A$�Gc2���o9�3UJ���r��Tm�*���n<�h�j��B�u.���v�'C/�n�RCXE�����'75���S�b�'s���o����찾�|�X2��Q��-�����g@��]LTd�N7Y�}��V�Z\ګK���S4�>��ՇO(ftw���j��xN�1���EC�us/Fʊ��r�2�f �>���۾��{)ȉ-2���؍���nL�����Wl�S;+U⒙.���E*�Ō[3n��ߠ{RK��f
c��5��@�ۛ��G89���=34޸�D��c�"�&Nf�����a�X-K��1��CC���/Eble�2�P9�V�;����q��LplSZ����M� ���Л҅��p
f��T6^�����b���1-I3���l(�S�sQǛ����e���p:�T�-A�Z��yϲ��Z#���f�˺a�a��h8�ܓ�*��S�H�Me�6�Zo��z�!�[ ��z��#AQ𫑝��;�OonjM���M,�8�0���;oݔ}2]	�>8�[�'J��b�nĺ�MA]A�VR0����7x]Ή�[>��>b��{�[�ѡ{v{A�c�mG�P��9ܱA�J���s��Js��y\��1*Ws,_:̫�o���"�s�iݥ���s�:�P51��;�e������J�7J�Ԗrv{��)?�:[�nwAm͕c�B�sr�-S}�\h�m��$��Ѡ��/�:õ���i^�䤀iOrmho�!��۽��.�3�U���˭���Q��7o�W�ʏ']�[��)�]���I�k.e�]��M�i�m�n	b)�غ�4p�UԪo�ߖ�|�u���RE�a�o��F��inP��"\Y����\]�o\��B��� �[����RQ�� D.�zv8iPح��e�R��D�{!զ�W����Tg�*cI������\Of��+%������*zs>��u{P��EW%j3��]�c�����)�kk���.l�0qw;�,�G_`���f�7+0�� Oݰ��\����E�31�/��}N�y���v���^J�Z���Yx	�VO��N����Yޮo2Z�� �҅g:
���ݹZ,��Ww`ٝA�9ڝ.7f��b��Mr8=�I<�*T�+z��:+���	i�j�!}!��s�Q���6��X�� �U��{��9]Z�<��ѡ*<�9��-i稓 ;צ�L�8d#V\rtJܒ8�j��*��5'�(�}�J�Q�Ʃ��Dt���u�����iS;� �T]�RHi|���i�XP�꽔�rV\j-8�g�ӭ�e�H�d8����[��ʮn�Ӄ�b��V��le�X�M�
m��w+�l�Q��.5��C�A�\�\�3rr�5��Gv坞|�?_�.SIfo�0����κ���ҙ���Ɋ��*5�s���W�s]���Y��wk^���".���_�o�tхd�N�X�a��.s�2�5����h7I�S�u0"��2�<N���hƵ�a�ONQ6��j�eL�7��ɧ�mlڢ�6axi�T�9v�̗Rm
��F��)+\	Ζ���wZ�O.B(er�6�0/�v0z��ef@>�MG��
m���|�iWy���r�̧���GR�w�8�i�]��
���u�ǃ��n�VD�Oz=��k�GM��u���7D\�2.��r�P�mlW�	Y����Fq�]WW�;r:^*mt��
�~5�~��^�<X��[Ip#X��e��w%�w�#�mH-ݲ�!F�Z	����ӵ���nWE���ڰ�[R\�tq��B��nJ�n��Z���⪱�VL��5d��ޖ�cГ�`���n�q��vL��=c"��P*J��[���cZ��^�F�"U��]XZ~8�v��7k)���|+�<#Pe��Ek9����n��=�T�e��g%���a����>�(Y���k'm���S�z���G�*��z�� (���.��u�n�T����H�f���Fj1���gEK{�rSz�cΕ�,�LX>b�k9�L�XJ\��[C)�� :и�8�j�ܥ�OT����9����+j��]�).�z{�ͱ(�O@�!�,��ۻT���{u[c�r��U�l��u�����(��wm;����,{Qi��h�����[I���\�bW[�g,h���ajʜ���Zb�Q�@�Ahs4-��=�i�Ll��yjdܨwt���-=C��q�yrVm(��;��y���R��sWS���X�]��Yf_�NB���L�KC�
��j�?��tV��8��G�+mfٴF�"N�*N�Qnw����4�Ҧ����ٔ�$A�sJ�f�J+�P�[z���BY�CM-�N����o.ۭ�3�-���ٽ���k�е�pyխ�ږ��r9y*�o��:^�FR�(�ޫ��Z�iJ���c��S�bEv�c�+sZ��CǶn#�xH��ulc��
�n'�=�����{�3�A�LGe�m67�����1W���G�Zi�-[��d�>K�ݪo7k :��
 ��ڀ��bdn@n�5��۫I*ڹ>L�ʃ�v�* �0٢�v^��
��ԋhڂZ`]o�Q<�{�ryI谻xUlys�H��p3����*;[�ͫ��KGE�a�	�cv����8"DZ�-9����Xi�7�l
lp��Un�^W�2�T�;�h�X[�+�-*[��5��}֥�s.����8e�&��x�41�#Wl�������*�+F�0 u��P�\�͹ӷ#P4sC�v!�����d�&�(������!��Dr;B�,f��;Z��J��KWڌ`���m܋�ݶ�В��J�*Ο5�WV�c�G�vvq���|�-2@��i@n9#�Үġ�5ws�`rTظ̅�V˲�J�]��tm�93�)Lp�r�_T��9�I��[ه��4���5���&�E| ���	1+MqN(��J-�e�}��D�����2ȜUe�hE���á����cN�ص�tZ�sy芫7��]�Ufʅvgd��tD=ݦ�����O�oł[��q��Xm�{Y%�Q'F��ԡ�D)0���K��W(�f�ȎN����˝����S�u3�|�4$;��5�:V�/n辶�b��P�a��u��&����n`O�[���{Kr��(����n�*B��_-ᩉwVm�<��*mb	���b��n�._jWu���M��^�q)Ҋ�-W[��tҪk������+)���3N�r�)�������6����b�8�,
����V��m=֨a�QIn�c���+������@7i�x�)Â,����4.���u(e��Vm�����S1�́�����կ/ν��I��A�¡t��^�h'x~��gt���d�ű�n7G�7�yKr�q7��򥈾%d]�wQ��KXF�i���IK���։����?%�:(L�e��>�C�l͠d�K��4�坏���+d�}�k��ւ��g ����jW7W�_CVڸu,������ͧ"���!�]�IdB�:�ꔀWu��v�q���X��lA�4-�xy��b婔ꢺ���L����ŷ���R޼����&㔡��V��������t�T�ă�[r%},19pzb!��V�.��!� hz
E�������y E8���`Cw�-#��c"�h2�*���������Yc�Ft�>�Кkg�	sB����'+V�E�k�g7ܥ�0�ɀ�ۍ+�	n�,��m`�Z�D�8�]�V��	��"�v���m����^�aeM}I��6pEhs%��n��,���IS1W�z��T�ྵ
��{������Yx.�ҫ�i4�Aփ�v:�w�NG":�2է*M�tGuα׎�	4H�T�B���T�{�w����}we�+wxLA_8�@�u��H�Q%20l{s��� Uݵ�
�e�po����`�y[J�k7���Cw�����,P���9����	���5ǻ�cw��r�i��٢N�aL`U��|��/�a�}�Z�ȷMR�K�7i���0�j.�oG[��6�g��A��89_CP���p��K%�V�贽��񽠑X�1E�ꗪi�pع�b�,��VE�/kQWL��z̫���Rs�J�#y1`��z�כ*�#7[����r�E��w0�X�k�*]���U ���cÝ0�z&�(�b�Wh8S`R�0@�e�SR�ʽW����6��5"��ujŵ�cx5�c������т]�x`����t�Q��ӳi,!����h,�]N���XIĈ��,C��"v���Qi�Ⱥ�&�����]�܁�6����C;@aĢśJ�7)��'E����jT��	�ݹI�r�p��*�UU�����7��ҁ�xN�]e���ĭ:�yܩ�٩��N�웗.E��m�,j�=R1�N��];*|�)��Q<����b�z�	�� h{u�)u6�����r���;���p��k���X�ַ��`�?����6�����m�y���^���������]˩IRV��+*]qʳ$V�p��A�1NtڬK�7|&b5>\kQ�VФ�3�/��o�J =xkp�8���[��J��wu�g<1�[( [�%���נ�:�m�R�n#�ҏ6gF-�X]�u�uE�Z���.��I��!��΀�FY��W��ꝍ�5� h�#�	����Tı�7�;ƍe�9;me�����i��ȣkp��H��YK�=u�+;���q�9W�R�x]#��*�[΅��6`h��[ɗ��VbWݪ]c�����`���beѰ��/b�Pr����˹"���0s�Ń�EN��GkI�X^W�jp`vm@�1�f-F��N�� ����5W�&Y˫y��p*4D{Yw	�HWvSȊ�5�D�#
�O����`EP�Ǘ�;�Q��
 ��%��y���8���&V��@���͓��V�}t�嵪��Ū�x�n�ơV⩦�
�,�)�;[�#�ko��i�gϫF�(����N�v�r�n(^l��q=[jwږ�
���)�vT��E���q#9��a�m��[��Y�����w>����m��Q]i6�@*����.��Y?��^�U���A�mN{�L��:d�,�hP_�{C#ݮT��J8�cB�j�-ފ8����G�V���Gq��q���E�:�^ṓ�Yح�6�&U�J�ogdS�����:K�Ѻ�R�.����{`bè��w��.*���Eu'ׯ_P
T�A�;b�nH�n�.��H��Gr�j.�ٖ�R<$�9gw-��h�
ѕ(r�C�ퟱ���ݮ�w%�H�iZ)�Ը���s	G�z�"��4Xw�S{h�G�l��Ɏ�r[ca�U��Ae���r�lH��w���Y�BV�@�2�[���Q-`aV];�#52�?���V��ȼ�k��ho�C۱s�7b���X5�P�D�Aj�����QyR���)Wl�;�2}#�m��ʳ����*�m�GY+zn��t�Gs�s7���*AM9�i�w�^Ґ*,/��*HR���J��Z�Q}��i�+H�2�r��#�F�C���hSZ�����"ʻ�8-+����˾!�IRݥ[�dQu���`��rf�C�6�;i��<��k�����sc�j��Z��=��p<dwz`֛h*sv\�$�%�R�k��!�ţ��]ZWY�(� ��ޣ��j+z�֣2�ٴx�e�x�pϕ"m����
���jX���&�7�Tm�Vb'iwT
��į�4a��s1���� Y|Vv��3��O�����}ϓݢ�EG�Co$U�L�w�R�wC��fQ���Z���e����N�9�⊀x���G G��nT䈴��j߱��fLDa-���VZ��5-�_bۮJ�U�Nޫ�W*�yÈ�����C!Pv�݇5�w�W��&^m�������1�c�]2�؅��xSQк���PN ia�&9C+�����rɰ�Ԫc�ںy��b���@ޥCs����)�����Dv+"�J�ܒ:)�Ï2�>e���gg<��:KM�"iͼ�Iܹt���%ZaxN�=�*sj(�˘'c�W����ve�Uq�e��s�V�Y-N�O)T��FܧP{�r��=QdEe��$�v����N[b�^i��0�9t�<�z>q���y;x�e3��)��^D�[Ŭ��M-��ܨ��l�(b۬��M�J%�>qe0����+����,U��5�r������'&<��ٕ;%�v��j��6�9��ܭt�`V�6� .���]��$7{�d+:B�@VmBn��8Ɩ�9�����v
4�-��<����=6�;#��tz5�.��m".��4����Jǣ���t������,ը��6�i:,E�^",�P����mBr�oP��z��Z�1C�kLC�)gn�z7�y-�T��=��)�V_[�1{�zB@hU�y�k�D�ŽB�S@��b�@�OW0�w�tQ�cԬD�~7�.��n��Z��؋��]*��^Jr1��9��Qm���� �
�蹦�iq�a��:�)ԁ��q�����l��Hvݵq#Y�q�C��C욅Ӭ堊U|:՞��IE.��\��,�1j��r�,L<
�Z���hTb��h��M�k;��[�Ůk2씊�,��am�v���F�%��UԳ����z�9�w�鎟_\"�
�W3q#7*��������1��Auu5�Wu3��J����#܁�]�2VLλ��֘�mh�t\�y�bt4J>]��z\��M��[u��#yHmd��"��\�mW	���`��sh�+u*�p��u�'��d�;����IS�^�y��Jލ��u��u����պr�8ra��e��u�yd���WO� *�N�NgǖND؁4�ʱ�ʔ�	5�
ѹ�Rܻ"���C�gݩ
��]���gCFḳ/�S��5@�(��26�-�*�z��s7��N|�yk��T1�`8��%-��If����6������r���l:�Z����Mo*�U�	ɕc��}B4ao�t�\i�9�������F���ZV۳wK:>��[orl�.�4Cz�8�wP3pd�]/�U���z�An���n�swZ��	�3��������E�,A���} 2�̛��{0�Ӳ�t��NL݊�A�눍��eMt�[Y��u���5q�]�ؓA�Š�ςs�n!��CD�R指%V��S����D���2YϨ%���̽b*V:��Ⱥ�`�RH���I}0���r���]���rm���܎�|澾�cJ���f�M|�v������,��[ 4����'5h��<ô���̽I��أ��[F�=�MYGb��ݚҾ:��}��%��q�8V���yIᵔ,f�[��{`�SR̡7�w�������ν,�<���L�1i.�`"|��бK�u٤h�t�� V*J�ۼy݌eɁ���ln�z���L��3�J�b��)Gu`�[��kX�ݗ3hMbq	59�yl�7��˙j^�<� j�[90$ӄ&�O]�R�|�W.�|(7��PY���v�q^�G�ܦv����uI�yZ-ic��K$�(rFr:�諚1[q�D���t�jU��L�b�h���ٽ&Aєyc
��Ō�S�s������	pG'%��Y�&�F���J;�;0�ln�Mb�s�R�����9�s+�(�W.qND�e�>R��V�	����ú�"��(wv8f^���]ݷ��+vQ�V�2����b�f��Y@mkKLj�1n-V�n�)p���-m�8�R��$t�n9�o${u�\�.U�Dk ��9R4�Ю����II��b��R�78^�b��j�#��	����u�lܕZtzw%nc�(@�@���V��Ʃ�*�:�\6�f�Ջ�n+��a�4�'Ҭ�bĝA�13m�KF�X��+���o3j�"w���NCv���Mo�z{--6U�Y�R�h%;���u��h��t��p�{���%M��IapF��S�+$�W{Si���4\n���t��N��n��B֚fi�R�a6v�_]�5�������/���r�,wc/N\q�y��R��T��I�ݔ�����n�15y�ٰ�-#X�b�J�0�"���=3v�DB�1�^D�f=C��(�n�g��֮>���f��\��t�\@v�,,_�M���V�P��b�e�s�LC���Zk���N��	Vږ�ܴEwD�+��ŽC�ZΜ�XJ�e�t-�U�#��D��_-�=Zf�׺u^��`� v�b��3�GL!VB���)�^�����F���P�(@¢�����ih2?�=R�b�}�:�f�F�u��wBj-�����x&�Y�l�� wV��s���I^>'X��삯7��(Gˤ⠍.�((d�U��ʦa�����4 ~o�ib����]��#�/��q+ip)����0<sc� c���m޻��V���k�g��GY�A��s�Ȫ��&���{c�I�kS]
��|6�ء��)�0�.���Q;m昳rx���5�h٫��gJ��IT�pʛ�m⬠�b�Q�RJ*	hU�ܵ�����k�]ۿC=W-T&V5+�>��36�i��C��ٵ��D�Z꼭��,j�J*�h��3S�$�XeoCI����WX݉.�=dܔ6�@�	��7E���ת��A(ć�S��"�\�D'6Ȏ�f�n�*�g:OUԴ���|C���\p�Ut����k��D\:�d���_}��YFb�;f`�G+��kY%����RK�&c�}�Ǌ	��-l�:3���4衴�i�t��T�@|��\��Z�p%B��׶-\;/�t�Ę��7 �ͧtw��,j*����yp^l���3X;��� �:OMMX��|�:�
�t������v���G
vOx�f\\a�ڊhU�ܭ|�,���ZWJWm�a����ԟ\ýV�Ls���R1)9�:
ٳ`{��j�4��=vn����b,Y](ώVƅ�3+AEv���Ք�ܖmI���N�����%Z�d�I�i�@#b��qfґ��nҧ�KՓn��| ��x���:�f����NR��l���
��[�a�	��򽓻
��É��׊�K\e�S���h�׫2]f�u�yB���p�:Τ��B�����&dް�AeJU��md�X0�Ž��T47Bޤ�G/M�nW�!6-��.�@L筲�a:ݶ�r���3�\��]��Z�f͏��L$a��P��F�eg�N�Tuw�ʮRֲkx�`nj?8鐰�o(@��q�{k�̷Vɲ��R�ƛS�HPۚl�[���a�R:j���)to�X������?�v-��@���wt�侳�h^lC��H;_^��-j�,DӀ�[�f�'��=αt�V�B[��Ѳ�m��<��s�|�bvFV͆��I��DL��[���>ݚƎ�j��C4��AWԍl��PbN�ܱ���E��+4�!�4���i�%)Y���ݴ�ܢ�WW/<z]eٛO;Ӗ�*v��8ND%Yh�a��Z�F>ͻ�Q��5��B�]���<{���i���+�=��[�6�ɽ(�+(�D+su�)���\�M��#� �OU,�q��x,�ј3mܥ3�6�����%�r���x�P�[,�m�Y����؊��-���� ��ޥp�->H���se���7q*`�w8+����u�Z]:�ptH��6�A�5���1}�7j^��jT��I��c���Ȋ�oC��ѯ^V�- Ʒ(�bے��*/K�t�Rd���Tr���w ÛC2f���N0���Q�n
��*NG�Ү2��'V7V����rw��Yۑ|KD�Y���Smǻ������^��^%{��Xe�u��;,��u�b�Pʝ�/��������r�v�"VC���Ou�4;"g\@�u���A�P�ws�SJ!��K�{��\�������N���b�Wl�L�7/,�2	�d�ب�Nm�����N��G&Խ�ԣ�U@`�8pV	Җ�c�������a���Z��]�.�9��#FS6X�#�)]���»:�"���Ysu�ռo��4�ԖI��-MvdJoN#��z�PژyfT�L謺{(�cSH��V"�o��\{Ǹ�:��ȱ}�쬝�b���c
�+� CWqt��i{�0 x���PV�h�D�Ց�CV/8H�cz��v�j�w{�Ik�OJ|en戧8���iаV�іuj�-8��Uz���2�(�@൥�kon�@' :�L�?LI:p2I�^؜N��5�)�n�1[ܹ.�4vq��F�g��׌M�Z4�k��"�tm 5��B[ډv�_K"�Y;�m��u*�<� ,ZlZre<6�����Q��|�y���S$-�� �)H��"S��K9Cs����wb
�P�[���g�d�l�Z�ʫ��h,n�H�֯Ue��6�o<�Ԯ��B�6�*�� �u��;
�\N�ʵK��*�����dw+��a�]B+δT�ql�x���[����W#����yk��[#���9K SN
�/�����(E�5*̶֑�(L���f�z%�[7=@:�x7��rc���3KՃ
�K����0���zeA�F��T���v0mSOu����o���]"WwRR���و�vnC�E��1/� �ۭvu.��h�u%%������꼵մ��i�T��j���V{"f;��Q';7K�,ۤ�;+*Vt΢�ձkC� ��)7�iY���Q$�k��;��t�v �K��ka=P�ј�*�F���PX��@Uw�����Ю���<핼�V��[��RY��%k',o��-��r��ZU� ��M�7��|+�����oe,��ZS.� ���C]�dr�\�{2�7,U������3Qr>D(h���t��+.ӂ
6�Z��U��r�c#;z�OL�-f�|�\O���n�����"��o�pW}J���]p��,r:���}X��B�w 
ۓcoF���O8�͆�*�.��ݖ�B�l�#�?��]/F�RvS�+�.�YO�"�4��s:��o.;�ڻ+j֝.J�@���Kw��6�50e�=μz�F�2�x�E�gi�vV����!�l��4̏r2��*fn�[2�h��q&�}x�V���\�)o�+ ��w��W�� B���!�c�_w%�0�Q0�n���뺻�/�圵�@��ەδltJ�4s���g'\������Vj��fJ��]�܍CvB4p�ؗ�}_UW��}��_y���8U�5�z���+��4�8X����LMa���S�`%hiY�\䭅� =�ac��2�n� ��a�]L�:����pq{�A�v1�[�pE|��cǥ�j��{y�Q�@}|�R��{�w�0J�`-�]+J<���ӶMm�CeN���s]�`=��=�\��qʁз/��U���BAݸ�9�-�͙�^�3�`�O�W]B��G���0�ű�ʹ�R����zGą�e^�9u�nܒbJ���=7	Q<��+Y{�ą���H�GP���jM�}��C8q�}���v�fB¸4���7xK#��j �6�$(���j0U��n�:m�<��d��)�]kw����JC�e������)^v�[[1��*�/����ur4]B ��.䷸�{F��˹��S4������v�ۛغ���_n�4����˻�\�Y�$_L9��RĊ������l���8���aKDVOQ�����uq*�ݩVw�a�_`#�U[F�4)p�!ҩ4��r�r� �L>X���%�U����tU�3N�h�ީ��ZF�Y�>R�Xηx(��$�ż:J�%�iΚ�4E*�{L�����F��]˄GjԙV�s��Ѩ�c���Nk=LC�Շ���S���i a�&�t0���.�A��n.:��KC����+j��$�F�R���
��y����V�C��ܹ���U�rr)G\�V���4E\��v�/=֢��EH��T��.��K7r�8����z*{� �U9���.k����!�@�Ԯ9����ȼ̴ܴ���'/.y\wR=e9%�c�����������AK�i�N�yܝԵ�:��zn�������v��ܽ���%��Eʊ9z��U��5�&S��rI�N{Ii%g$wC���U;��@�x�I�r�N��-Z^���S�eNez����뻥��e:*�^N�\��H�b4���N�d���U�g�+(��Ku�T&<ȫ̕M+6E�I��n9{�y�q۹��莧����b�27u�v���'K�E̗v�䓓�dNK=�B ��B��P��(A���5�C��sm��[q2uo�J�H�=]��aij���wVmJGPG��jN�=C��g>������d�53�W�J܅���J��PGYH�Rv�a�*FM%ݴ�'ԏ2�װ]��g����EY�W]�����P����1�?-#.s����B,]���;���VѺ�ֱ}Y�w:ѱ�P������Z��d#����>���: s���/to�ԁD_�FW�P�'�ߴ�^�[��l<��R�m,җ
ಖ��r2p$y�S�=��ӓ%5�Q��8Q9�x��8�T�"ʜ��Gm>�5�H�b

��n�c%�oc�97��WPz�8`uN��@xn��|���y�ϡ�6{!�}�S��p���@إ���83c��P�<�9U��tX�5����Pb/d����S�j�Culf��%��8'+/��3��@Ї�|OW��̨��J����.��q�e�s�k�h��18͸l�jX΅��\��	;�L�'���ĩ�T�P`yO*��d�F�#c�)�X�[4�	q���r9He��!����,��U`�}D<�E5���2��Y����=��x��N�5C:��.PP[B�W�3��ʬ	d3k�V�z�gX�nM�s1Լ�zπ��nᇶ�YZV[f��3�!��s1/Z�J������Q�����v��b�}��l��V��{Q�A<��^�A
=��]���G"���Al��s�i�#L���/:�]u�h�u(��<��I��;ʧ%��NP'��q����v'\4d����eϓ��o��t�g��'�vͦ��Co��X�qq�@}_	D��u�dF�q��ڮ�QɫC"t���XD�{�/�vxݪJ:�b�禷8Jő6`�>����[^�Q�u=��~R]�Hk�/��l�C���X���@�X
eƒ_o���f/�ׁ��8���t/�A>����rB�V��j��P�y�F�t�W�cn*�J���L����Ʀ�������D�pq��������w�"wh�>���y*��w�x<3g`��m���F��Be����*���ѐF��j8+�ZL\F��f�/�T��O���i�<��ڵ��׾+r�*w�\Uns�W����%A�.��SҐx`9yր��bіt�O��54;�����N�^�5�73�����Y K~3j~ɹ� ��� V���N��v%T\3U�Τ�w��@��@��J��J��o�VX���:
5Z�N��]'�v_��|� `�0�@5��>J忳��%�*��$]S:�ν�@YN^fj�aA��6jp��������pE�+]�]��Fp\urr�$ͩ\\n�us-l�Y+����1���מ���j	�b4����.���Qy.)�Uz���A&�<��Jl�N睒�mFq�^�/����3�369�!�Z:6�iQ0y��u��f�r�X�Ffܸ���q��Xz�7 �a�n[)ӯ����C�v+d���������ޭu�E��b�&+�����P5���Ƹt�3o��5��b� Iz�A���W[��\��
�:����"��|n����K8H��,`����)�, ���
�b�|F��8o����mp�͌b�jȃ0�IJ���'�Y�_p�O�$�Qþ����i<�vL�n����o.xQ9���TP��2T�10"S��+K̉"�\k�)��Wu���,�e�$���vpG#��`6۽�V��L��}RWM�0�&xED��b>Usշ��[��|�T�Z:LeG>�E�!�\�%�5�>WĎf����S�B<y�]�����Y�"k��l߮_1X��g��nxT��i٣p��k�j2*6^&��x栤M�{��Hİ
ԖʹNv8����7�Z�h��BV���JZ�U��im��Y4U]�q����q3�:�p���AI�gǢy@мݰ5NZ���ܭNMmC��h�����`�9Z�%N���͇��CB5�JI�[�V�e��r�ᮺ��\�C��N��~��B���S�Fcw׹[������p�L�Xv9�Eݢ�
�}W՞���M�[=�b@���ኽ.��?T��7�(C��cE���b�U1\߁�IuL�@�tݶ��1��6a�0�R��Z7iu�Y^��*VB��s+���a2Ƅ.�/nW]���G���HCE����{s�ù�.�|���N\��A��9��g�(r�W��t��T8��q�L�Y.(ƣ�ڿ���[��U���×T��~�|<d�����?xfd�r�#o���K2]�@�eRx��gˮ��ř�޽�Z��Ҿ��M��9�c[���a�'-^����K���2�L�k4��P�����5���D�;]��a#މ���=�Z��Q����3Ԅ��w�A�WI]�Z�\L!���[4�C�۝k%��/;cw'�Ǻ��r��W���G����>}�Y�D>4$>�f��Bq��(��H�1��F�kz�m������UD) lMP�T�!�D�C�u�g�����T���.N.>yJ��z�3���ݭ󃕮�Y[��E&�ܴԵ�M�+��*]������FCm?
)�:���{�V4��T���a*�ne��	x�n��7�Q�ͮPU���ޣ�u�-ڐ(㛓.<+�滆q7���.�P��ck�:t�RfKȗ���0�i�nH�x�E˚FR��(�0�=t;��������^��Y�yܕ�QBѼkWȉN�0iH��0Cnbn]S28��|�H��5X���vWM��ܑ�!�z��l�PAi��ܺ�Cj�9ŢS�7N�v�<�H
�j��u_sH"���J�'C�_Q\bk:�z�Ha@}S�4����e��ֻ�\��ً�ʦ�,�\hG �TB��Ga�2%un����D�'徾���^��;;A���\Jn��n�Og�����&:Y=P�M�
��鸭�ţ�Lh�3�e8K[�Y[�-��]�\�E���m��ݎ&lC��7,u���M�W�J��Yݮ��bO�L Axo�����:W�O�S�{�Խ�zj�\RZp�u�QE~Y�k�س�����H��9G�<Q9y���Ʋ�uN�.
�aI��75�Z�� 3M��j��PgZK0X1������a��:��0���W�����|�Ψ�u�iM�Br��j��n�/;������Q���Ѐ�Y{ ���Kn���f�c�=y�Ι׿���i'�h
#��m΍o
��Qr4���״��2
�)m'⵹ipxcӊ_<K�:n�w��%f+�f�;[�j[}U
rhD�D�>�y���x�o���7�	,|oh��ƣ�@%�j�x[$V)M��Ճ����OA��=8�t��%��]��KHn�kI:Z3ŕ��Hסtʱ��v�����@��ʸ�؂4��jj5V�|~���6`�,gB���iq�I�Ip��뭥��.:�x82�\u%"��q�:�=:�eicD!�:��3���P@�$�9�A����8�ف�7���h ީ���T��n�!���<u�_9z�8��Q.�W�(�̵�z�s�e���N�Ĕ��)�	(��s t�����ڿ���rZ溜`yx�p��
Ҫ�6�z���+ڗ^w�� wd	�`�"4=ulԛJm�s�˔=� �r�a��g�}s�KoV��If�h+Dق�cF-{Y�q�+���YR]�Ѿu��\}�f"6�����x<�bw�����5`*��Q_%���.�_*=����r�ul��;;X�*����.#�u�q	���y�F�t<f�m�$���N�.���c����p�c�P�����7C�<o�v�EA��.
�~�\�͌�Dr6��E��Eϼِ�����T�E�� iQ�j`��<��U��ۇMs���-TTH�:
���,c\�����e���u1�k;t:;���Z�Gu=<V<�ێ��8ƾބ=�%��]$�e���ӯ����\*�a��ˇ�;�c"O�MC����ڇ�V���<g�f��z)�\�r�+{�^S�hW�u��@RK%��١����>�\�q��~9_Z�!�+>7���//�gsQ=v����f���D����Z V�b��t��>s�(Qy�������Q���:5��:�m��������,��Ε��ʔ��! /�Q����7�RЈ��s\�h|��o�л����k�v
$xs+A�����R7s��	��onW1q+l�j.��'��Q�S/�/�qUx˭�Sʺ��T��*�_���3��x�4)lp��k�m�c��#�@#�z!�l��n����gC�q�V��t:��2�z<V���d��t
U�%����@�bv�����s��p�ֳ�}o;N6�%I������ֻ�!��8̠$�E|T��u�P\�|$wҥ��)��Frf�U^�h�w��[͋�����J���rY�F��� %:N̬�?p���>����]9ڕ��0�W!n��꺑��2�o��o��G�к�Q�H���-��85��F'��wWӳ��M!�����:�k���(����7���}��v2�W���!�hZ6_U�\��Ne��5��4���9V��I�*Kz&f�KO�4#�Lo����h{�(��z���:q2"8S�Z���Ϥ�\iц��+b�:���8x��+�ܫ��.pCg ��߽zכ�I�$OQ��_���0Ty�Am�-��/�^,��ԃ�ԃ���tm����s������"��4fc��uAi��lQ�Gm���m!�c�U@��x{?�/i��懮��hө��ѿ���v�FEl�2Mb҄�Z�����-i!zN8~ڀU����J���>8�ꯐ�I�п�`)�NX]Y��/o�h/���EW���0φ*���?5�o�k�zH�0pǋ��7���
��5�Q�+n�Z}k}�Z_�U1�U�*a�m
a�q�6;����ϸJ���ӵ�=���W�&O���eo#{;�	9���T�4Z���{/B�S��8b�;#�Ȭ�ӝ�h�!���59���s͹}Ѐ��ȍOT8g���������լ�hY���-L�f�����C���F��ō������W��q�,�]�@�e'�	c���X��{
�V�cA'���N�Zޒąl,^��d
��N����[Qh�֎���D�
¨=s�AͮZ$��+pN�)9tx!R\�۱����՘��:���%���9�xu�,��^g��۠���nS��&�!�K7�E��<�pX�\��m�aӰ�>p�Ũ�K�ts����J(]L���tYf�Z|F(t�6[:�w\����'sm��G�ֵ5�k%���Y�+U��QQ�iHm��qI]�Z��q0�V��ja�w��zoAfy���L�w׸ 5 B3�?����U��1'�k��N�na-�W�\%!�{D-6��F����ްY<�bh�r�T*C��w����ہB��H/�jh�e.��,w�1�z!�"6��qN�D�*PdH�ߧL	dz�9�yw��ʯ���0��b���:l�&��C1b6u��ّ)���;�4N���&`\s��w����,�C��Y�^�Pz�A\~�����E�LZ%_���1ָ����_T)/vwG�:>�A�9U�\��#C����&��jW!��>���,���l9v�D�c9�2c�DJ�IK86��z�b�u�bT/Fgq�t�?-���|��Z�'1�b2]rԍ��.i
�健�3C.�����妎M�qN�M����T�2nXr�.r�*��^��aK�S��ׇ���6���M�3�4��@���rd�6&w`��)9�v֎eG���w[YNi���՜c�4N���3.N�X�Ue�s�Q�&�U���ھ̊�\Wz�G���n7w��.��މm7��!m9���}ֹ@����+�n�B�@:1�P����_�9pa��,��2~U29	vE�=�:Z�#^�r'�Gt�n;m_�x)|��+�zX��� `���� ���3��2�B�>z���u9G��'.3����
S�����J�og+�~�c�j�L��K+�h�� fUP*!�;O�|��� �����ρr��#f�
:���}j-G�^�k>�Y\.7���J\g� h�pX�]}���+�H���:q����dsN�;��[r�k�U���U���Hn��N����֍z���̗��v�@�q�1�]㊥�>��.1�6b�cT�pJ�a�ɔ����N�[�Y�1����ᦕ�9�2���mCθA�l���QP �(9��q('S�����^��T�5 ���몓9�|j �x`���;�F������!q��]ʢ���)4���H�>�@�	tv���E����bs�Kj���;�Cr��D}QzbL���G������C�wnVέ��Y�r�ͩ�+�'
y�j8m��5����[}1n�����JM�Y���u�F^��kw:�c��-���<'�G��43�+���q�S���wW5yH껶�o)���Z4�F�X��J�twd<���|v�h��U���n��Υx�+��a��¦Ә��R=�/���8���x��-3��fފ�N��5* Ϋ��R{-�`믅�ɡ`�a�W�d.�r�L��ՙ����]ea¤�I��^��u�ʬ��Sl��Oz�9������s�M���'��R�]Eɼ���&�Z�߃7�������K3m;��V�v��6��Ǵ�+�M�7CN� >�n Y)X�i�6�'%��s��� 8��,�x�ֳW����s��e�ֺY����q�Z�!�Ff�Yk�\
2s�.�����7�Jx>rmgܴ�9���m��t$ʜf4T��K:\�C=�g1��jY`o{OR�h��2�8�����
w�u�\)��B�+��Ce����s��,Tta�q�q��"��a��8-L��X'�Yo�&���d9�W-Bf�uk�t���1�uE@kA&���z6��lY�O,��[��<��[5Z�3$,�̠�z6���*���\�7ZI��'ed��Ħ�[�����+���'�X��C�D�=3Ӭ��,;�V<:���G90[ۡ�5��[���R$�[kFR׈eh��Yv�wB�Q�Uݼ6�o��L�т�I�F,�e���*���L1���1.b4�6o�:��R��.��XaaJ�$�f�́ʗed{1ڼW���S��(��c;��]>��-F�������e��ñ�pܬ�b�T�w�:^V9�p�������kU��VU.�ȝ�Xd<OT�ЫSR'
��R���a�������5�/x��]��kN���9������zX�Y,B#�0�eq�\�����e�l���]w]���kU�.t��:U�t-�3@(&�����k��N��`ug%|7��o]2�D��4�iv���N��,:iK��5I���=�����h������7���Z����`�%�.���y{H�̦�-1�QU�M���D9v��@�FB��S�oxgh�ʁ�[Q�:Ŝ�R���X��tD�+(��R���}�6�`�<1��5�m�*H�D<WKu����I��Z�d!-�|��[�=�.��6¼��Uˋ�q){D2{C<��T�+!"��6����Z�g\]��C��1�.��Zj���pKH<Rjxۅ� E������C@���/�-z�F�-Vys���y5-���LZ�v���"����aXن+��Wq�:��N�,9G���Sj)�mŨ��7�V)�PowU�NRƃ� r�u0���~�Z~/�ZSt�q�l��j��V��ǼV-�)vn�r����	)��
d
�y�by`{�^y���s�s�{�绸K�T.m�� ��4��)�Hq�莥������RE)���n�rvG5�N�8NV(]γ�]s0�$*�IS���3J3�w<����.q�u&9L�"��\����=��Rs�8�N�t�,ʪ���fB�L�]�%C�3A�S�i����WGdYʸR���E�.kL��:ӫ[�{�9�$TE�T�J(�<�Vjy-qܓ��	s<wv��c]B�J�U:��r��r+�L��YUw9WK���Wwv�wOY��W,��r��=����=c�� ,��{�q!�s�W;�(ʹ���4�(�B���EQNN]<�G5	�,�qB�bI$�$���2�Cb�6��*���1EhQ�Qr	3��{�x�z��:����Qz���Z��a�\����A9r����T� ��d|Uj��k��2Fh)�f��t ��Ciͭ}�K�\N�6�V�x�+��m���w2;��ˬv�7Fݚ�ZX����#�} }C�B'�Y�y}�ɅS���}C�x�V˧}~!�Q����Ʌ�x�������C��7*{v�F��?8<�����ې>���DF";��_|����";oψ����o�W�̧��OV��>�
@
�e��P�nܝ�����]�ڭ�x����O���	8hߞr��|�W���9�ݼtbw���=��yNM��;�|q��.���zL*�ɧ��x�d��R�U�OEt,��Tﾉ#��z�>�÷;}�~O��u�&^}Bt�S�����N�y|��N�>;��o��Å����M�?';�G��������P�My���G���e
ȕ�e��z�P��E�D1b${|��<;���|������®=��|���~�w���!�ϗn~���N$��~����7�$=���x_�nNM����~���<$�;rԇ���v�b'b��P�G�}c�z�����\����ϔߐ�����]�7��{�緤�]��߿�����L/���6QC�xC��~��}�];��=o߸=>ݽ'8=o�;��n��O]�縟
|����*�]>M!����LG�?!�0��n=Q�]�� ~O'����;I���y}�rr�����7�'�~<�/����ף��>v��O�������6�F��޿{��7G���߻r�B{n�Vyw#����6c�#�c8�'!����9�'�=��	�]�Ǌ�����~Ǆ���=�rû��N�v���z7��ޓ}Bt�y���ϗ��z>��~{�bw#���NU�o�wuIɢ�����#�|�>�����M�=�~���=���w�����ר��~C��!���]��s����yL*�OHro�$�����ߐ���o��� }I����엺4��h?�����}��܄������-�'&���㲘}�]�'���}v���!>��?�������������������^,�7�Γ��<&|w����\y~�H�#����r���8�\(|/�/� ���S����vm�N���7?��9��Ͻ�;��n�����I�S��=~���	0��n����w�i���|O	������z�������9S�[ro�C�5�|yג��&��\;��S��P��9���R(Ȋ�e"�:�ݩ�%���d�����2�B��{]��K�4H�E{OV�#[]eͥk��� �����q�Vt'G-�ͳ/d�U��]��*���ƶ��76a�ff5���S5��T��I&�>��9����'�q��\xN�oo�xL/��>�y�xy˼�}�&�<�����]��z���I��'���ϯ߻�~O�9>�������P��A��e�������I���"c~��/MDǿן�o^;��ﾽ�M���;��X=;)����:9��������n~&����Ɠ����}@<���aO��&��G��o��s}��Dp�;�v�Vm߽���+y{�?|�㿐��<�&�BC�����99������N'1w�ܛ���G�����z<��HyL=~v������@����x��;N�|�?h���c��9�I�����~�&inyg����w��|O��щܛ����<��yL.�����s�M�P(
({O��u�0��]$�~���v��?�����۾������|v���y7�#}�M{йA�;����k�-{�]��q�w�ޓ�{v���}�ǔ���ܝ�����	�	�O;�v<�}�N��'�<x���x@��9ӵF���`S
���<;۵ѽPs�������0uu�����h��u-Q�#��I��'��ߞ��P������q�v��ݼA&_��ۿ���?�˿���_�w�oI��:O�,x��xO��<;s�c�<;rro��ä�.���=�~�t��
Q��j����+�1H}V>�0~<\��~NC�5�_{�|C�^�������>}��˿;���~��|BM�	/��7�99��������<�����v�܅����v��>��nA�rEZ��5����#������;HC��<ߝ;ô��}B�m��w���m�7�{y7����ψ��ɽo�>x�yw����>~�����>P�=}���������>�o)���9�}��o�NS��|��1H��������|�n�cί�<&{Au�7�90������ʻ��w�ŏ��?;<�)뿻o�O�o<��0��������|�'~�߼mV�_	�3�ߗ�΀wv-���P9-Z\BP��L}BA�z��
a|,|��xv�;�7�~Nq��ǚ�O	��㇣����G����s�[�Ǐ�I��|q����?$�nס���;xM�	Ϗ��k$TKY��Ļ��GU��P9�ͱF��(<�z�1.+���<��z�e ����[���..��t��o%bK��]}��Wvn<[m��v����K�8ul}��:�[�齪\
�d�M��������j����
�޵S�ev�:��$H� �ϝDZNߞ����yv��o�����yv��G���\xq+�8���}NNC�ǒ��bw�?;�Oh{O	��_����s����¸�BM����=���N�MU�yV���M��D��{����oHRq�x����nܛ����������������!�0�����˽�I���I�v�N����<&������o����?!��1;����7��x�7S���ʙ�k���P�(}b$}����S�s�O}�좇�z����I�����><o.��M��nN��}��q������
����Ǐ����������k���xNv�y�ۼ��J�>�9����G�"��x���M��w�����w�b}珎�ko������o��Q���}��S
�x;�o�`�}v�?���<��}q����y��90��{O_�v�����&Ǜ�~��w1 �=���L�3�����
��>�H}����I��}O=c�ĝ�[۷&���c÷���]����<���ﱿ�}���]�����{��=8\.���}�)�<���Wz߸�~O��!��eWܰ;���v;�j��b1�{C�wRP���S��������8���+�	7��u���7�;��<?��}I޼Ǉ��ۜx�H~M/�o{�߾I�!&�����o���߾���d]��c;�ޟ_��eH�<��Ν�߽��򛐾�{O߯*�S~w���=!��bw��z|8�}Nv���rs�~�y0���{(�����Ǔ�s�;��7?��z�zL��~�6����f�s ɛ?ޯ�U!_R�����q�����>�x��+�����P9$������������w���I�\
o޳>]�;��Ν����<' N��P)��)�Su�� z� �FOc��}�b$|��z5_�&'{O�9<~����S�'�?xğ�� _��ߓO��w���<te��C���z@𓿝����ϫ}v���s���p/��
����A�ׇ���\�7���{;��ϣ���G�?Q���p�]&�{O��?8��_8	7����������1;��>��!��ɇ��ސ��w�}C�����q�������!�0�����?������(̯�Om��ӕ�~cM�=6�x?p��ե�ӯ9�4V���CM_�s���]���ueoΏ+ ö�*ԧ۰�5s��������=hs��uSJ�ʻ�c+�ih���f��\��uK�Vwu�ӳ�,��Y�1�^+��A�ž�@�D'Wv5B�����CC!�������E���%S�nB@��;����xw�i���}O��N�_��7�/������p)���|��Ǥߐ��$����7�ӎw�H}[T������H}Hx,�8G\��K��՞���G� |Cu���@��}���ߟ	����[�xL.��Ǡ�����ra|��=�_�xC���m�c�+�;����ԓ�~����o�Aʾ��P�"96�S�u3ӓ>��mmz4Dp���"x���L�C�>����1��L.�v����Ô¨z�c�}�9��]tbw��q��q�7�yL.���yOh{C�lr��i�q�<����1G�n/k�ή7b\����,��!��"#D��I��^�}��>;ꈗN��@�}��~BI��߯��<;˴�����<�p�C���~NN~�"/�d�����s��1��r�������9��v��3�[>^��Q��rw|s�΀tle#n۱�������c���+2�Z'%�5��a�\�!���.����~t&W����Q^К�)��4n���X�7ar��yK�g��f2r�S�$3�x�:�[��^�쪔8�5�b���~��q)��R��:I��B����D��I�^�W^��+�*@b� :/��"��y�)h�Wx���ܢ_�ٶ����|�NF\��,x��~bU��(_�|���[���ھ�c��'h�-5���v\��~/����<��Khm��N���#!�]y�o�C�f��W�0WRI9Χ-AԸ�21z��WL}w��؅�����:�i�Sp�m��%��ӽ ���B������J>�0K�B�Mӫk��SY��Z���ھŵeo*�M�Q����۫EKܨ��n�9/Vm,ٵ�^_:z�N:�bH���=:>aZ�w������[|@6LO��$�L�#�Jf�QuG*�0�zu��)�L��:�,��BZT��s���!w�9�e���(�m��5��վ�{�`=TM���,���%�)����პ:\TG9z��?f����54�j��;[�RY�P@�F@s�0��PO>��(E�:09m_�졪�Z���G^�{']��:Z��}У�����*_��P�=���kz�	uK��;[px����O<�Q��C�ʑ1,"ju�\KǑ71<~��^dG�e�8���,L�b�(Rw�|��V����uM|����� h��Հ���Q_%�w��ض5~܃Y�x�,t��M�Up"��mT��O2h�n�����$�*���-C���	暝��ՙ��0X�s�>?c�,�WeD��mI<K<��`xT	�n��.�r��u.�m`��ғU����h�9X�Ю;~�ȯ��h+ݙ~Ն��{�ϫ���+	Cv��ո��ڏ6]/�s�[�Ϩ�e���l�=���yהiK�ޡ�F�K!vg��05W����i�:w\zU䎭r�Z/�Y��e���J�9��)�o�Xd���K,�y�ƕf iN�4�	R��>��}JV:���q���ޠ�T��A|'�M��ڛ�8m!�џ8�T��PJ^u��c���n�pɼ�3�r��.;is�h��=����B��;�EWat}��J��K�KJ�*'�Tkү9\�%e����ߴ\�0�*����U�.��yӒb��,�t�atV��߻�+Xѱ�It��6����#��ٕ �'��V�y1��n���Y���$�:�'N�zz��� ��e�u2�����I�G��*�6P��n[+��mL_zrj�7��f��Mw˞��(��䂨�`!
���[t�NZ��j1;c��\:C2�GunN�
�LP=5��V7rn7�9�S<��j�(��d��^�Y�Eʖ0	�2��49�s-��l�g5=՚a�Hö�85۸y���V�UuG��7D����.��k�����R��s�Y�Oiމ��%S��&����G��O�<�B �J�P�w==o�_M�~W���~�����t�5��_W'I�.pCg��o�mށn�K���G������\���IS^B��wV�� ��!%k��rjr��ڬ}$�_n]�t
��TTcA����ng��a��tta�l����{��h�t�Y�;(!��!&��X.%l=u����Se��+��5�^䱹�e�U�Q&o�5��1Dz7
���FgѲ�Zт�νC^��,��K�F�
�M�Gl˙������{Sr�Jf�U��$Cbx紴���=��ȵ?w���zR�Mb�b����b���1��ea�jd�_g����5���{AUC�Z?'����=vǽ�1��n��Yr�Ԟ{`b^ݞ���K��`���z�wO�O�0��!�}�Ɓ�+>�q��dUoF$��Z&%����<]��Lr��Cj;hVM�a3pwj�e4`�z���ft\f{�Q!�y����c$�zKR�>*��뇗��W0E�`ٌ��f��tE�C2n7j�QjBu�ZlԦJ92��o�ױuMw����{�;Oլm]�>C-��NĨ��t���p�'�t�3����5.��.�V� �:����I��uO��V1E��|/$˃J��M�'�t��:$=Ҡ���4����+�P�ȐN`��N��+��S�X8'�d��Dڂ����#@j?w�*>M)�ǅu��\��h�7���q:��$�N|;����*��&C���6�9�g���2�C�{m��upd���#n�3�Bs��47eb%���.�w���|��;�D�ѓ-#�s`m�����9���T�l(�AF����뼙Z�m��5��*$c��;3�@��6z�N��|��+���j����0�_�h����B���F��J��*���xm�:�<ĭ^2�q#���(�=��Ի;�C1����7^���y��d���bh����	̓�
�a'�2��Ӯ#UX\r�WKǋ�c��rDk�R/b�Z2�BܻݔY��j���ITh��&@���_8���:8&R�_�k>&��p���n�rΨ�ǚ��'��o�����tlH� ]o��$OC���0�X�a_�q�*#�[dAmYd|6c��p�V9�M�o�NC=�|�z�jm.+�˪	Wu�0ӤtyL�4�G�ש\�2al`S��LnV;�t\Ms֍���zt�@�5:"0	N�&8�vAx鮏t�^�OpNqh2�.�y?I�b�8���A55Ed*����z^��t�z�N�	��tݴ�B�A.�˘Ǩ���I����4�����΀tnQB6ύ���\b8]��`:}��8@3��r�K~��3�e��ɹ�����8^�k��o�Խ7k�\���x{��{N2���ܱKqu���oa2C��6]l�Y���;{hs�u�+���ӯ+{� P�����9��u��ջy��<�����p�R=)�j�O�J\F8����R�G�����d�'�V!�yR�J��.ٜ��Y��G����3����u���a5����z��~aB���:��d1�:�q�\�a܏���ң�$r�;S��+~[���@f2���W��ݧ�����U\��^ں~�ݧ^��}z0�Ns����E����6�W���A�����
��iH	f�K�;g�gD�E.C2��q���Q�Ss������⬿��[Cn�i'KFx�+��JÎy�X�\��@9.@D�
�Q�]��.����/�w������[|@6LL#����k��t����<ӗ���Vt�ߌ�?l�,��4&�%o�Ds���D!��u��/��L�V^A��Q2�'o��{�DFD��p\�?Z�U�%���l��|��Gy���n��E��Qw޺���.�T�)4Dk����J� }7����N�h�m_ó-�'l��,P��O_��w��LZ3�#���:Xg�W��p����4�;G*ǲ�K�T5��N�p�{��w.�2 �H��ńM6�@.���,���q�;"����>:a�Gۺ�|-Q~u\u��5� Z:kW��b�tV?{ͭh�\ᥐ�I����G�7��k�.,ޢzǓY&�'�y����YN���d��i���c�)����!pf(p���pĶ����]�L����pdv���>��*��0�S�t�~���;*m�/�^<pC���Z�T��y��:`�X��5�jg�&Fu�75g�Z��N��2�gv�T��Q��|o����U"�O2h�6�y�5CxŒe��w���l���HӒ˞!A�T���yLU�L-5חv�W���w�곾ٰIyZx#h�3��=�qW���U�(�P�].���{
��ZL_۲����T�#�Z�<�7�Bpa�gg�N�W����Q;W1������~ra�u0�yր�ǔWq��y��Ӡ�r��cLHwؾ��p��͢���>��V�s��������3����r���耾�P�8��]7	���Y\3�ɍ����̜�)dySd.��<c���O��Zz�BG�f\pK,����_k���~PV��=u��Eh��Y�e�S�ƄkX�L�e$�Lo[�&1�p�@�� �al�yC�iB����)��U���u�#��.+d��X�,B�J8���_*`�y�}7���=���?v�Ԏ�w�[��2��ո"x�4�T���Nվ�Z��W��iR����)���43� 7%�p�4�z���lJM�s,��F���0����}4:m�	c�Ӆ�FT���W9-d.q,�&`����٢�� ��4-�09��? ��0�w�OEv"GuGv{-e.lt����|5�@
����:���A�i蔘�6y����e�������iRY����4����bP5� �M�Z�u�Z�YhR�4��q��D� ��}7u�Um\/�G��O31��VM�&��A��g�ZZ��n��-��������4	�E�r\�f�Hٔ�s��+#z�v82���w>g3��z�������	44p4�ڽ���5�28�NΜeN��>��[�м0�:X���*/�U%��t&5�:��c��]�0vǉ�t7��Y؄v������>[m�����V�n��}N��hB�Z��roB'fo�9��QIDU�������\��v�n��b��e#FtJ���۱Nܱ�_I��xT�bԻJ��[V��b*����3�b�*�.�_Lg�[�b���v;*<��;�z�v�5Y�+���(^�u���w��K�]4L����7`xu����iH��%
V�2����N�r=�hݝ]&�f�ݸ�S�g�h��'�h��3 Y:=B���Zr���kU�����[�n45�g�����m�L+���=���cQ�zw5�yS��蔫�
�vT�]�S�,���=\���vܝ���"�'��Q����<�����1Ԁ5@n�� 9g�K �3{!c'i�'�P�W����G�xi�3�����NFY�M���Nc`p��' �J�.Msݥ�z�\:�2��$n(I:eD:�>��g o ���La īq�}��5;5��Z�Q�?ƶ�^W�.�*���%:'pͮ��I\����:����a���Zk��vgW(��6�]mM�@ZB��-h�3VvtN&3���YC~Q]C`gN��5��on��������Ah��uݳ�N��#�1Z�il|i\T�5!qe�0��ym�:�W���Du�ۧ��ڍlU�qo���r��',f�sY�<�ƌ�X���8���-�Jev;mM�D��F�2���ڔ�q���P��A��˜�}������EwX@��k`f��q��W�+m��z;�	ͱf���cPOlgDY���B�.�	=Nʆ�Z�� ��0�W���	;���Ou#�I��Hw���!3�{��>���YwMع[5/�N���v
�X�ȫ�ȡ������r	�^�pXw�N�F1������i�c'L"�cd��HEX}f�r�Ԇ���f��@��"����9��t����;����f"*���ܕh�e*��}b]iA`��ăS$�9jY	���wp��tC�
��ʊ���\$3$EH�<R�Ĩ����rwwO�S*�w[�ɧr�iQE	[�H�8�֓���z�-&%�ѻ�L�åE�E�
�H3��n�W����s�92�Yy]z��,H�s3�*�s�����w<�uP�J�wv�g���3ݡF��TA(%q�NT���ùYP�AU�Q�&����g�y�B9!�k�w1,,iTEQ'��ID@���x�SMs=B�"T��R&�ONgws��G#L�Ѝi\����69�=G/GsU��i�F�]�*g4�Ku�B���S�V;�ud�E�^�%4""Ř����u%�f��ԣ�'sBt�D9kJZ;��f�X�@�
"�)}D�
v�1C��u�\�W>���xˋ!�y�6��_
����D�ζ��n���4��]0wuj4%�*�*͓st������W�}�z��f��� I�����)�g�B�GI1��P��<k��9n���dek�ݶ��l[��Z�ö�x��\�;nc��Pݻ���_�zL?�I���V2%��3�B��K��$��KuPC�~�v��M��TF#�erG��1?�k��[9���r�t�ˎV�. ��>6��˓��f�6C��[n��U�&�L����XB��Ēޚ���C��˂`�X��/N������X�רk�)��ZG���+",Md�g��)�s~�S[2t*@/�M`*��G���W�xL4�.ӳ�w��杚9���{[�Sb��p�k�yq*׺^�J2~ڃ�*�t���g�rѤ�~��`կ���;,���-���)�NXy���]ԃ��*�M;ć�ô2%ו����E٭8�;W�M&�Z�t4F�·Ω��Z�3Wb�����(W�WR#&�	���F��(2^ޫ淄�֊�5w3Ϙ8\�B0b-�}l`!�4�1�bw���7s]t�1�>u�.Y�s���B�-暚�	k�
j�\��]\+�qgs�ƌ���P>G������\ٕ�T ��z��"����v����t]!8�؃���^w\�gJS�N&������c�
��>K;d�Y�Zٔ�!lr��O���;yx�y�r;�<�����.��T��U���䷧�CA�@ �eVk��x�i2�أ�\Cj���[ŻD�����*�����p�	�~��c�%��fB:�o�:�d����0��� cty6=�ǞZ�teE���=Nj��K�^#�+��V�M/
z��=�f�Y���W*u DPپ$jcP��i�E��e���4H�1��*Q� F����TT|.�R�X��{o�3ѭ�����b�-L�+�8�z3\L!���#�ޯ����qʃ�\0:���.��\�@t�`���/ݥ{��%����E*xy��b{D-7��F�7w�h�P��;���z�{x��8b&[*��X|r"�Ws,w.a�ӐܑP�܌�uh��d]�|7�qOd�O]��T�0�� "���@��:Y�%�{�����?��;�����
�RS�3Fz���mq#�}�Eԭ���BQ�.4�̮?eG.�����1S�yVU��y�a�V���^�z���|��k�B�i���"�CJ������՘�3H�ܤ2�|Ĕ�X��D�ú/4e�id)�֣���55���N�'��&r#:�	�<Q�˖�E�����0 ��o�F���-��W$D�`r�22q�O68��w��v���m��عt's
-� M���$�o��}�}��F�%B��u[�(~�?$���2�� E���D�D�!a��ʊ��Ճ]�(MY�!���ĸ�wۉ��
w�8Cֶ�mMQ_d)9`ih�^�����~ZW�F�(}���#7������T�L7��SOH��������3a+�͇Z{�Oqx֟'O/�t�X+ ����t��Ω\N�ҙGm��ੇ�.#���R��ݬz/ޡ]<�J!��ê�W���/G�(���U9G��\Fu +q��1�;�HNX���y�$��ϣ�=T��O��pV����uvO|2����_U�a��J�b� 5l��d5��ol��G�Q���Rk>����4�'��z�x��JVg� h�pX�79��ۊ尢�.�`���ƨ!���)M�k�b9��c�|�]Hۋ�$�#���<.�T��h�цn9C4u��T��Lv�G@h�%w"8�zs�?0���pً�j��9\
&%z.'4�؍N�v�,W��	�������0��wM+|y��0G���q�uu9ǈ�/�o2- ֕�^��Rp���.��(]�g$F���^#Z�l�	�l���F�l��˓"�� 4%��.�R�m�tʘ�gff҅�e`����y1�lG+�����Ȑ�����+�j�8����5�j�^v�9û���w~�>������/.]�?`鯺$����iO�WU&e���΋ϲA槨�n���ԖNw9�Ց=�~�T��
����62���I OE{B.�����f˛���X��u��J��޵���HU��Ch���*�P�ZM�ϙ�ɯʱ����n�R�ŧ�+�4sj�_���mցn��U���O�;$p�d�r�;��Kתl�QqE��q��b�ԍF\%P��Bn��� h�b��T���mL���кV>��ˉ��ޝPf�����7Ҹ�'��jbGD,�dѿ�t�W�cV�;q��"*���,�TQ��:-�If��x}�����~�v�[Uλ��
u����/o��(��*��En��^Be^Otգj�pߘ��Z+�PU���_=&�up�֦0x&���Uʺ�T���S:��8|�#G�o˓�j'������lW<5�JE ô��sov�=X��(+�9uB�:��c"��5�}Q�u#v�x��eNz�z����M�hu!���pѷHP[;���޳�]+lrD�^�����bV����N����~�נ�F`�|��Җa�/a���%�bo�%��%���*P]ݯ�p��t��%���/3&p{AֺrNS,�X=6B+|����ٚa�C�#W,J�]�s��_}U_U�z�RzxL~)b%d����GK�h���]7��p���dVV-��LY4>�a���),�'im�u\[�K�hyG4<���퇗�9���;�:̨�	nJ�s�k�'{Dtz�"M������j_L_Z�&+���t��7�r�F[U��ΆzӇ�����P;��� �<
ᴔp-k˔��L�w���z/��j��@�N��ND��F�v�m\>�5��H��Oq��=Ċ����-R1��J��m������̭�!�N��)��F�����u(�T�zb?�I��rC�Khq�x���[�_!X�\M�Kw,�ߡ������{U�����$y:� �px�v\�|��)U�U���b5T�01n$�|qq�����As�9�yXn�uX"w���ݔ��q����A�&������� ��������)�L_-�E�1��.m��VMvq�x�:����њ�M$S|H���4fc���:\��_	��E�vy!�(5Z�fW��Ik�iʤ_G�te(xX�F�h10aj�'V��z
m�����p<�U/��G;����'s>`rP��ה�o����6@�lAJ�nu��v�E�=a,�Ⱥ�,�Tu�k�0t��$1J����zw,���R��KU5�.���7b�諭������S������U�p�u���p*��`:0WLX�R���j�a��Y;�������V��v���L�Br���yU/�}m�x�P�R_�n����.����J�d.�6pBN�4\��/�Sk]j��1AN�f$t�Ȏ�
'(	��xO-���M�]��a��]K�����8�s+i�zKR�4T5u����т*w�BX�~�Uq�I&�
�p������s8vO2Qȍ����}p��SI�L��w�m_�&�x�$g��[���?zOȇ�B�����\2��]R^g�_1�R�:�K�T�8%��g�}�r,V�J��ڤ�C�L[��^�K�JP�	�'��A:to�3�G�a�'Ro�N
��� �I�
�'�Q�>22xCn[=��Y"��KK�٠+Q��U����@�S���Wr�ޕ��&��N���<ҝ��q0�\=�����M��+�ȁrQ���O?���=�(lx��7�
���ϧ��1.(Σ�.�Y�+O�R��>�!��{D-/zdg7w�h�p�6�i42�Fj�C�Lc� 3sPyعT�9ps��i��t1H��L��������hu�EƂ͚�U��ԋŮ�2���Fz���7��9�@�f�4_>�C{�΍��Z�Ko$}����1�oBj���Tu���˧ �n����NEe������}�qo*U4������|1U!^�]W��Ю�:\�����W���"3����9�z��8Ky��Ze��"%AUD�BU�L���p\k�]\;>�N�1�ޔ��]���kw��=����F�k4Q�����É"�P�A�1��W�]�:��?b��갗qJs�N���h�Hhpy�,��\�}�v�&ї'�L�V'����L	"r����CO�U�.gr�w��N5u�BL��*d�Z�# Nb8"sA���yP̒�T�}�^�)S������!�Y�"�y���71�L�0��f�\��=,�b�[�55*zG+���ٶ�ظ"�� Re+4�8G_'w�:ѱ�P���۰�5mc��NrĎ1���ü��������/���F[��ě��i���gJ�����U�x����y�kz�A*��k�5PV�gC&,B�Nu9G�œ��H
�k!�N� vl�T��ݤ����']�v��s\���!�AW}�eK˯1v�/��*��	�)�%wH�ԗvގjH�x3ևP��	 �f&n�Q�/���geٚ��N��+*:끾6f���:DK���"�k�j]��}ʹέ��m����Mp��E}�jNۻ�X��S���zF�9u��G.�6��W�UU��ޠ{�w���@�w[_ʒy��t��w_f��xf�Ξ��J��� �	½DT:��7i��ms O�Z�9p�GF��Ss���b9��c�|�uԍ���$�9|���sӉ�mo1g3u�D��5G@,�%w���}��_��1q-S�B��	�����[}�#M�[is䉇���'�]	u�����Z��!a?%o�G9�84B���Q]q��UU�d㷝i]��^@6
* 0��:x�?\WU&e���ų� ��0
���(v=�29�[k����\+�4x��@��<��$=苇��?B�����E����<Gb����a���']���]�鸊4�Ԍg����Ai4����փ���\�����5ڪ����r���b�&�mցn��P��p�inr1ꬕP�pr��`�V.,�����*@k��94��Ö ��P�T��n;�Sr}$�̙�zŴ	�g���pO!Ry8�'����$R��M�m�W<�^�"B��t��59K��n�c�m�N[�7qG*��(�?"F�]�&pJc�.��=����^b�8�۫�f$j�9'�v�g_����JO��G2����S��v=���Y;5�£��k�ӗ(�J8���;�'�
�L�9R%��}U��}�޾>����^�?�a%}ʼb\)�<,y�S��vz�쨁�O{jt�݂�1}I�RvFJxw��_2=��Y�ܵ	~`��� �s��!ᱝj����A��ν'(��@�h��'��v��D[��������rv�}�����~�V;�L��[�x']x�~���ė�:^�;`�0�#,�7Ο9����qϵ�}YWR.㥓�faa��i;5�}W|�g��>ޢ�m�&p�~���D-}��%��l�&��5só�$��&lڭGL�O�s�����g��S~>&w1ٗY,�j9Je�����xFga�s�{�<oN���f��lj?2�_�Eh�zI5�O0���iz*��F�9}a����������
QR{uer�;+n���m�ҭ�����'�'�>����~\�@�]	k�x"�������p����1��Gͫ����~��A$�|e0q 3��neU-�M:1��n��ݜ$\K�0\s�h�k��n!�p8i;w d�h}�f]�4�V�7��*N!�u\�)2*>��f�0�ѳ*��V��w���/�� �}{z_���
�{��zG��QFL�Z��^@�/!i�m)YRP3l�4Z����7�t�ct-�����Soz>�oH��'��I�V�{]����<i���}U_}���r�tN�Kx��pG\~�*�z*+��*���zNti*��]&�L�3����x�;�����j�f�v�piX@�Ǳq��9H�.pCg ���mށ�9G��:�}��t|�ו�D�D�*Rv�������~��zi�z�����|�U�w-����s /S u��H}j��E*���W�����+N��^>л�<�4��M'���r/|�Z��-��K��C�������}+�0\�xko{р���r�T��r������_7wB�`)���UK}m�x�cIan����}ڛ��p��1n�#��۞�����VK���!��ʘ��4�M!S�1��&�K|��..��9-&,E�Δ��u0������h�CWQ=q�ېFR�~�k~�1�퟽�����«�vQӑ�U�Z_�K�q��?m/{�&Db;�!��U)��E�ME�]s�[K�ꐦ6��讲�����gП#��=��vT>�9rN��-rdf�Nu��:Y��ռ-��e���|��|a&��E��<�7��SUt�3&�Aѫjٗ����[VR|iP���d�\B��d\&��fhAg[��ӯ:67zs���9F���m��lB���� 0�T6�Z�jJt���ZoQ��@f�wq��'`�b��8�%t%�`�v���2H�鄻����RD4�w&���"���)������4�^S���V)|VQ�Z���j
Ql���0�/t*��H�k5-��,ѕwZ�Y��DE)�YSb���e�b���W���M��R��;�[Vq�ۤ�M*�7���c�C�|�J)+.��3Q������
�gZ�;�+�¶�w�ܽk���і{uo}EG�;�_�6Xe=�em�s�r黛���YpǼ��W����6s�7w!YX��(D�]��)<=JΗHva|��&I���m���gcT�v�Ϯ�ӧa�ܶ�����U���v�X�gLsF��Ji�hl�s�;V@�!z�N����!x#W��li*��.1��\���&�^]�޴)��J��;��,3I�c�q��һr�7M+4��c�tS�@.\r�X�tw�BKXy�8�
�7��ƌX��V��v�i�]�qf>�4nA��N�XX�oFJ�� ���l�4��ҵe���7d'��Q��<��@�v��GP�]X�vd�+��̉�ive!�y�3V�mS���B�)��J`h�����V��֏��-qѬ�j���Tk�v��.�W�vbG�#4�C	g����cirf�u}��R���p��]09#�gYH�q�ӓ��u�2���0��Ѯ30����V�^�Ɲ��[Ֆ�Ṭ���)�7R�F�
���󾩘UJ���#)#�����8µ��5[Bb�D)j�Y�0mظ�[����e��7D�� ��ރ����A)�v>Y�7:���E�d(��&��j�S(�[��bp�3�_p++t�:�e���������t�N�cNS����D�,���-�զ㴑v�:ub�T��-P�1�Ӱ�K�8�\W���EQn�ZR� ���暵[NXɂ�ܜ*ջ�=��i�kcĵ��ӑK���:Cmn���рv'Pn�o!9�-���WV��w�)fr�]�<�*!�K��'H^���K-�Bg͌'��[N��ٻ�+
y:YP�y�'\���W��,��D��zKX����Z�8����e[T���N����**�p�k���V��{(&���:V�-�c�i�o�U�E�5�¿��%F��Aj�"�o�]�Sr��;ef2]�c)_u���@���]���֖�|P�Uh�ܭ�������/M�\��Թ#���񛋬�.�۫Zt���F��`ã����q�@�M8@���[���Kf��b5���J�sw�U��E��G��2!�����q𽧉���pGwv����6!^Q��;�:��wU�mZ�(U�/	�9ē,T7]�$�a�J\�Ւ�,���b���"�G�u��Ȣ���<�#)�aTT��+���lp"C�
jI��ԕ,�Y�䬪LVj���f�R�D�s��EUJ�dU!$�l8�8ZgHKd��xa�	�	�k�W�GD$Ԗ��!JeȌ��jZ�E���fW#���5MhV�V��,���R�Zb��H�DEtR�*�i4R��925sH0�,�K,I:�!�9瘔���Pʠ�4�Y�����1�»���QB�k��5�QF�7OGiD�4E4+M.GQS1'nfa�!)����]#�R(��9�J���J.�t<٨�h�$S@�r/f��U$J�itĐ�S����,�s�\�<��N�CIu(�^m,ڥ�gY]9D�u�:��Pt-1�O�ӚmB�ԯ6�VhfU��H�H���L4:乩y�JԜ7��z� �8�e�GUgg)Yopb��Ʉ��Wp0:�P���4-Y;`�b��gt�uy�|̬J`�j�.��%DҘWYs�ﾯ���OM�	O}�}�:��ۤ�	���w���t��w�p3���b+iPEk|/���:��ܾ��+N�c��z��C�"�l�;����:�q��@V���ʏ��Z\��(Q{i�2����h!t�؅�[����C/�{D-n�xT���.J5�%!�v7�r���ݔ�c�C~�h�UH�v]ĳ!i�`�O}�C1�h����T�n����gkrK�woohVd��L��� juH�*����*��)��_L��l��;N' F��Q�oH�w��w��nBq�ٖH"3��=S )��|*L����q�]\;"S��`����y�<4
�qҲ�:��k�B�Պ�wy�˧�/�H�u�Q�D*Fz&��MV=�&�L�i����S���_0����ŢU�_D�~�\���U�PS:GG�w�^c���s�y�U*��3��֪C
 >���T�y��}DF)�D�D�@2
,R~��dnyC<�v�	d�R�=Y�F��c��WF�2	�K�f���{��qS�'��U��+1�]	�t�<���fS�v7P_5\:�Q���g:�V����JW�zQTf��8��.�3��^�f���U���e��M�J��u|�rc�5g�m�;��N�`�8���K
S��8�'9ҰO�NǗ�����3!'W��>�>��	�|�Ai;�������鿕���ܭ�[����}�g?TG��|D�]�;�kES�dٹ�"n�ߐ���uԻC���e���΀A �T����^b��r�\mu��o�1��(��G��.��iЪ
--8RG�2pu���|M�d| �;��ض"���$��a����U��w�;i�T)oF�2�3L|P�3�A�%�Ѯ\ks�܆�8�۾t����g��u�i��^�T�,���c9���z�c����暉�(.:� �}ƨ1$wإ7=�)��u\��ߌzrԡ�������8��_h��N.��eFǔVw]���W��i����0��cx�򽹋�USquK1�1�d�	;�2�����]L��Ȇb�ʉ����1?Lx����L�[3]֝����w"m���(�( p��@GJ~���E7_��^��/w,�Եl��n��[
�Pq����!
�T�z ��ZH����گvnѝʎp���^>��=:+�����X#�^�3�(f�^ݱ�>�����8�i��ՊŎSndO�qdU��WkS�0u5��O�Nq̗�m��:L2����	�meg7�qX�e6�c����d�Y�qz��G����!V�����:0z"[W�g�z�����j���p��L��+���{Mgz�xč�D8��_�a���5}���ɫC"t��XD�n�6�+La�fL�7�v�8q����>(Z�_����n-��+R5p�C�I��^@t�.!�.t.�܄H��i�>����L� ��>��z�	��$�1�9�o��5�gg2h���ZmX�ͬ�t�ޡ���q���ʰ��*��°xX�3ǭx9�5�3bj���%_��e�Cg���k�j'=�^�l����D9Qr��	�
�<8*#�V�l��ܨ�y]��U�V�(n�48�O�9aC���\��Q<,m��~�Vմ���N	�F�0�d��� `�m� n9�:�t�O��D54;�}�k��*�E�d�i��*\��H�hV�X�Tv[?:V����&b#�
�K"�?:��ϼ���g�w^���?W��� cфێ9��(�mz��2�ܯ,���W�-%�VK,�E2�C���Ͼ�x
�w�.��67;�r}����E�y+Z�K���Y�/Ā�%�-�d����x���@�/��AW�8��\�t�IU���D�:�V�V��w�|�e�6a������w�U��s��ж����j`�s�@��ۙ{(m������UU/\�u��N�����U��p�t]^�M"`�	h�iz*�|�4�9}|\pGC.cW3Bt�.�� f���l�N��SƑ��� �@L�piGּ�U�y�d�˂0e�{vqΊ��������smT=�5��p�
���c+�@�H}����o8ڦ�x���U±�;�}��1�ˡ���X;u:�"���ˡ�M�))�K����j6���SϠ*��}���ܷq�˺|wb�M��`���"~���\Uf<Mi�Ӡ �|�u���� B�л��NR!����6fG�������n��x˷��Y���?��hC�)�#�pfP��7x��]N���d��CJOCj�s�#�6f�=�ցJИU�hu�J׃�s��ū��C��Z�%{�{Ġ}U��5�I��q�O��'���bڀ�`�̉�dN���\b��*_-ڍu��u5)�M���3��6/�4r��FV��P.�5J���1r�̭�CBl���iYv�0Ս����#B�Τ� �4g]�֩��oY��{���ew��y]�c�~�G]-�H7k���u�w�_t9�;P��ky�2S��	׏�v�"쫇���U����}�G����B�x�a�D�Η�{����c��/�!k�4��y;�f����R���Q��諾M�1��3��ꕃ*3�ܞ}�R�\4��j�u����y��h��7����5��o�_P�*�nr��aQ|��M�vJ �<����i��x����k�q=q3�\�`U{b\�@���*9��t(ܫ���f�H��Sj3a�Z�-�[p��o��z�>���
�y��Ǯ���=��|1��I��4�wS�������>�S}P�ʨ�f
sFwdÆ��S
�M)m��/�=�.����^���9��qzyl�sj���?W�XNإ��!@&nʤ���E�JZj
O.9�[oBڇ�p#��>�<�̅9�$�޾�U���x'�Q�m3�a�o����F�H�� LU���e�M9�����W�Ȯ��_[��m^W( :/Y7Ӵ���ܥ�Z��;��y������)P�x�1v]6u���U�`�����[�#E�$��I75�$[��Y�'Z��+���ܬ���XΎA�#Z�lob��B��q�W]��]�l���p���S�3����"#���9n�Qk�2�{��
����%�(��F�ϧ�k�ٮ��3Qɵ���I�.9_s�7�äC7ݳ_"�T@+�h����ʧֽ=ӹ%��6j_��M}��jE�}R�a���/lY=��Z��SH���8��r�1�ۘ)�_�O,��[Q���6�j!c�)�����#�e��'~��22]<�˩1~��\��#W��g��d�-J%ٱ9����iB��9���	-�ӳ<�"'�8i^�[��}��o��Wʒ�]��;��0���ˊydo�ԥ��y����jY��3(�#1W�s�'��H�`��c�I�4��RPU�G�=W5�m�ޯ���r�U�|�P��"�:�{S2�� jFu�����]-62[}:��O:���}Lw[�V���QCeֵ�@���Q=+eC]�Z���*1&���y�B��,�[6a�';r�lqX.y�W/�=�:�!u�+X�8K-v���:w�0Z�P%u����!��c��,���
¡L���4p�w;���}ttKQ�5>Љ��L��Uujy3VwϧW\)恽��*�򀔲�h	{�U�ԡ׽��mΊqW8\Z�@����o���>��N��N�I�q�}ZO�T�<��/���bR�Kyq���}3����^�bC/�:�B��p(%�h_=JOs��F�e���j�w��۶��~Q?[���m����yٹ���Jm�.��O�'&P�����\>�JeY�n9c]��6��9R�+�ALw���	hV�S��7.�4mjJ�V8�v���l��:՝	��r�"|��a�ڌ��_���5�8�⚜o/�-V.;Qɥ�h;B�m�TC�s��J��c���K�{�"5W,Pk�~Ȼ'�9P�9��a�ǥ;�)c6MͩڞW��au�e^3���'���a���=;sg���~J-K�q��F\T�u�/��Q���vGr0-m@v�"{2�c���[��2��ִz��
���)�Uֵ×�o��Tk�u�t���3K�A=I�����u�U��(i=�c��wÐ���(
����÷�Z��
�Դ����G������kϰ��ӱd�����Z�꽘����0��u����t_^��
{fn��-��)7���a����:�odX���*\_;0�hl�d���P��U}D]����q3jB�>{�o�zָ�q�!��SY��	ה �+*�A[�q��%u����e�s��-�S/E�y�zbN�{�����m�D&��vVi5��2��D��@��\aQ1|�TGKM��Z��]�2$���5����U�t��3�<��q1��cf||MS=^����z�~�b̞��������/�R--�:��D�YA��M��iP�La��P�`�Jc������J5`F�j���yh/�P��mޑ���vQX���?4�Tw�����Dԗ��ƞ\c����[P�z���H��7@������%1[�D�k]:������6�ޅ�8�'Mر:v8�1sUT�5�����HPo�/�b|C{��n4�j3�
���y�<���������/�!��H��N�8��]��H;Ԧ���3���u�\�y-\i> �W��n��^U�(�n�M�%�8�L6�r`����2ԗc�k��b~���,��-�ˍ9D=.��3��9M[T���D/��0T�t�DR"]�fR)�s�`:Tr��؇j�J��K��/U��?��興�ڶf]5�H�v�)�5�!OM�jՏ������<z1ˏ_F& �"����ֽH����͛A1p�tu#�9�֕�j'l�X5&bl��|g]�w�sեR}S\�	��ЎBtE��l�}���P7�zz���n��C�\��_�yd�^Fk�i:�X�MBn7���dsn�7���� �0S�r�{��({t����r�y����9��e���8g1�А���y��.�t���~�sX���[���*^�OZ�]vb��X�9.�Zt��~Y�雮�����*����Z�g�����<k�[J����߱̚�n�c^meY��3(��=�s�T7Vt5x��vpΡ�hSҵW���o�
R΅]�m��Ȧ7k�=s�;��.����FN��	産�ƙJ�b�5���!�>F�WY8B�8�)��F:��J������ 3u�k>�F����c��T�����jc͞f��lߵ�W4��K`h�^A{��Vz�@EX���s[f�*����51���V�v+�C�tU�f�(��U\����t��VM���f�[˾DR��8*��������D͑?]��Qý_N�U�-�c����m>�9��e��sF�9�f�/y���>I�n8��CRv�5�B�nz�f^n�R@ENU�&�=Nw��neO�����ZX�y������!n���
&V �����=ٶ���X�TK��,ﷄ:����4M����� �o�l������I/9�Zpyr���Rwca�p�g
zL Oi{��5*{g��oN��,�[�y�����7[ͫ�v�M�LCv��\D�%�%9����/�V��Ν��=H�%�k����U�3��2n>ޞ> qkޒ��_m#�%���ሾ[_o=m����M&�[b;���t����X�[��j�'�i�]��g��
ǹ�+:�\ru�am\T�:ùmV�f{��#��O��4�/[�[��b��OJ��f�u��0�\�M'r�v%)P��fop�(c�W�^Н���L񕲃eA��u�7�h`��֐��ܤ�̈́U;�l��dU
��ՑJX���c�Ew$��P��mi����q<�x��K��P�0r,�:�T�{��d��Q�2^Z����"�ƅ�q���T���wEh���P5�0� n�b��WݹVw�P:L����{�s;�w�P��kl���/�F��}�f�O�k�B��sf �U�ù��+�tq�ʊ%f� U�+�G�b�[w7{\L�e�&��HVY�bqZ��/n�X��Q�d�M a�6�\w�z`�쬎��!Yɋ+�x�xh<��[h��w����.������ض�p���v�{��:6밈�M1ӊ�K8U���C����S�H����s5]!�ཽz9k�a���(Y�7wW:�6���]����/�D;z:�T�ݷz�� �* 0�"�B$��مi;��9�/Y<������W�p�3Y�V�b%�h<��uq�.��t���M����,�L�����&����Rʓx0�o*�Dv����i�^\���cF=�0�У���rsy�Q��wk�����S2hF�R���K�n-h�J_0V��F7H�؝���D#shaڤ#�%g ƻ��;�F	�D�3�����,QO.Q��fV]*�sd�t�i�c�6h�j��P����=l,L��7��J]��=>}�˖��m���kcw��;�$�B������Y4�]Ttm��oZZw5�{hj	1MsX�Gn7�s����Z�G��&��'py�����e��Sc�H>c(�K��|�=�;�k��[z�Q	en���	<Hk��eZg��6� �v�h@�ǰ���YEV��J��z����]h
�xP;�>�b"ո��������q�1>L�B%cKX��YyҷfC�EQ�YPT=ַ�Y{���ʕ��0��[���a�C��{NK3J�,�Md�,������k�.wͥr��Y��*�N`3_`zʗBӻ���r�G���1���2�1q��%
M��:�N���K�V�
�&�r�`2�'�4�s����)��-6VO�)U�h-��/0t�]eh.�w�@0���1��:$��{*P�W�	�:;S�Y[�٨1g365Y�����ԴmK۾�<�G�=�/��-���ݑ��EB�oj��-���^��7��2�ovf�9P[����:��Zؾh��4�0I�ka;֬1����Ѯ.L���?4w�6�.����Ȳ�Qv�"�y|�i��R"�4^�N���%�`e�"ݹCR*-�O�����ؙ�+9Zѧ�,�Ȱ��r�V��2G&�)lb�D��5����:�h���ck�����cLή�W�2�rr>ª�^b�_+y�������/hb]L'u�F�7J�%�c�5�P�E�݊>C��>O�*����W��:)Z�I:���GVh�P�wwH�)+%�)%(D�K��^���DGC,�8��䔹'<4��(襅�T�B�(J�0�J�5T*�TT,�$ʶj�	�H��qC+�wqR�M-Pۄ�%Y	�&X�m��R(�,�g��S)�q5f��J��g!�--f�N��"(��R����Az��y��J2R��!i��D.�sr]����'0��ݜ��EKY�R�f����H�Y�̭iY$r,6f�ΙI�,A7]г3�Ĉ��E9�2��!�'4KR5I#@����a�+J�#*Y�as%�r:)#����1$�#hЊ,�Qj�12Z�PrYz`�B�В�B��GNU�Qd]
� �C2�Y�'+L(D�L�L��L�n^Ҷ�p�RK$$��4-6f,�*�YTY���]LJ1Ui
����EiE�M�͑iTN��ba�9i���Q��dZ�C���Zb{��Jj�%2�+U5(2D��������i��KA�'<�����{Re'}�'$b���lk7ڀ�y8I6�u��W-)�[->��=��}_W��>z\RB�5��/�v㓍k!��|+�)Bxնhg��v�sP0�H�c
��|�)	�7�Z�p�\W�gjSm���S�,�i�-�q����#O���5|�''hJ]x\O�˅GKM��Z�O�m<��:�����܁�Y��@�aT����N��alrM㤵���Iǻ�����=y��n2�M���S�/js�uFs�z[�QݸY�<�wΐť�v��L��~���s* 5Q�5Cӈ���5�-�k$�-.��K����%z�I[��Ӈ�u�5�8��w(%�T�p�.�	꽃�:�=��{R�i��4Zyq����t��()��ޟ�H9���T k�bl-�]-��*��p�tb}A����OtW�ʉt'��i��ͅ�&6��ۭI���(3mWǵ]���.;\�V����A?ys6#�nf�z��G�1�Q�H��(�[Nk1���L�yR�qmw��oFU��]vZ�m�����q��F�Qvd��"��3��t=#�ۛ����*G���u��D�B�u�;����5�붆Нi\gڍc��j���5���Ji�N=��z^�����}��,f��I�gt��#����O''싍W'�юq�����38:�,U��k�{F�T��u3�����{��}\�4��'�96<���Q�ƹ�].7	������dLr1��w'n�y��ځO�MI�̲_R�G&�O9@:���suK)���o+]��c�-��}�t��)�������;��|�&���_Z��I������7Q�1 ��^��m�{���>��G5�W����So�������k�n��wǧ�]Q\�,�8����rjn�O1�z&���
j�)U�S�����j*���	O9���r�j�߳��W��Q�1�0:����2����m���E���폞�h�X��f��,k����&��`"A�j�)��d����}��m��y�w��tV����l3Փ��F��)�@�6�m��Q���푩@ѷKr/P�}Ί���&��J�S4љD�ɷ�E>d��(;�ԑ��U�܆�v��eKwy�r�KMK��x����	�����<�cX��]d��F)w�嵻b3(,fw|گ��UU}�<3������x�<w�IUF&���X�,��ۅ8��:{ ��ȾS͠��JRܾ�C��	�����:�R�PRy|��z��8��[��2IX��[�)�Z�py��Ϸ��ϯ�tb|C}�����zoHjۻ��w$c�η|s��3��?�¼�Y�~����s����[��ߟ���a�&5�u���6�
c�.��阞ǗS�m������Sg�Q�>K�8��5�7��6�b�)�G`s����kjw�3qۄm�z�"���_ke�}S_sLWɸƅ�BvG!����*m�jӻ�֨�que�y5�fO٫Ng�X�Jn3y���Toc���TE��i�>�ǟw[O_w,_nVV�|�Õy�N�j�&?[��?jA�͓���j����|3M����/9:ܮvT��u��.h�iJh�8�n�G/��@0Ӄ�T`�.�/-�S���l��+CJ�{U;i)�8�O�o{ � s�]Aɸ[
6�i��݊�-lu�sшddw4��C��YBf�>l�k^�X�G|j�Wh<r�ljK�EF�s݂���ٖTѝ2,��}UU�z��~��7{к�W�_:F�:.�H�*��ʀg��S��YԎ���g��m�u-/�BW1�K����kͯ���F��&�=��\���Gz��=�-�R^�
��:��ެ�7%�C"ߡimW�٨�?ZD=��[/-q���a>��\���=n(J�L�alWؚ�����s�S}K��ufӚ�b�<�(�4��@VO��W�{�'XX����\c��������M�Y��'��L]���o��c2~Z����T��u�u)	Ԟ_8ko�2�� ��!3X���o<�x�HY�ࢇA�Qk��d���Yά��x�TײJ��Mj��N3j3���T�)﷦8KE���cW:�;���]��r�i�.�i_�ޫ��6�TK�j�v@��խV�q�m���<O<XpH��~z�<�����ߛ����Pg�"�oUHZ�1]�8=��#Ot5�!ö�%/��� K�Իۘy���QV�6�6�:V��/݀P@���R�d�E�c������ �ҥ�|2&͑}}�%=�S�l8�SX��K:m	&X��D%�f��]uE�s?�}�}�Ds�s]\�Ht�_�75/rk��u�K\�I�l��p�A�/%����N�S�}<\x��U���x������V��pک��cS�,躃o$�]�H���Y�F,��W��_�4���}M��g�q����kc�֭F������O�C����w9�ޱ��}R�t�QU�,/U�`�9�ǣ��ɖ�ޥ%(��7>}m��
H�ט!}�jW*d�\�4�N!���r�4K��q%Y��f���r�o$�����FVuGޔ�'tѸ:��˅GKM��%�O��Χ
)��e������L@ڐqԩ���kC][�$�������ܛQ6��*\Q|'��:�}gj���~ ����Q�U}��ga���_ ��Z���<m���=��M�B����T��rF��8�b�횘y[����V��*�W�˵Z��r:C�#Y��LQ�<�-�N�|��{K�ծݧ�sk�o�����f�%�ۮ[M
#EJW}2�.T)'%�r��Δ�(5���ʓ�y��t"�M��[���7kd��^L� ��ׄN�꼌q�<6�:~�����j�K��{��?rmj��^��·8����og�A��碏(�hY��d�Ԕ��;<�-颓��v���x.[����w����7�-lN�ڗ��7���1�������7�p���{��3���w^4�E�o�V���C���B
{Ek��i�ɥa�p� [ѳ��}]q�������d�A�>ځ�����nTf�\r��9��Gm{B�ʕ��L���������P���=�h�}�5�݇�G==�́*7�n�W[Os�j>��Kn1�9��"a�Y��G�nU��S�x^���N��I��<�F��M��'z�:��PE���xF��-j�NM�gF<ʇ4��q��%uά��z���ܬw�r��\9���8�ݏS/��t���z�F����[C1���+�&�+��������.���f�S�����q޺mҽ�Z/���=�{��ك�H�-p����=r�a��ƬY)�*n����;iM�CT�b�^���t�/��ՊZ�9#Vv7J�w��6�h�O�yv���=�R@Q9!���W�}��%���o��s?<Af���C����^|�����O_%��m�7-�fs�v�S�f��֩ꓤ]�e4���m��_��,auz^���-Wqm��J���f�n�b�t��*����U����?P�V��4��zk#��+OcP�f��I��4˨��T_B�m��O��z&+��'���M�Bo��]KkjvZJ%K�J��ؤ�^����Yp�-���ۅ9��;}7E����L�L�r|���˕Ė�⺃�KM�s��y\^�4�L_�{�:�O���}�2{��I���W�Ժ�>5������"�aCp6�`[�fv�9�ٸl�c��'�*��H��s�v���m�Ed��1��Eº\�Z����`m��T� �:Bꁠ�}5+^l�6�F���A��w��@��i���5l�����b�����6����n��U�>��7�@��cmJPzo �ҩ���d=�+��K�\�W}�Ϟ�q�*�0�E�Obd�R����w.��Z����(s����)�^L�ڗ����<}��]l^^d�R�9y��*U�#��ck;0G���H���!ڰ�=@����W着��+�q�"k���>�9��F�]C}S_sL;����r%;"b:Z��X]���9E��S��U���̸�Y9�3�7��X�MBn5�k]e`3��c7�xϻ��/ղ�^��cݽ��۝)q�x��^�٧B�Cv�9��j>�iٞq��,7�r���}Ř�o�O��z���E��won!�9Kӫ̆�r>0i~��A�bb���*��(���v����3|�sQ;7��Jl(����ͽ{�4s#�̢�C��-�(���]�	�2R{��}����%�2)��{����#E��u��m�͛㴯^� v<�iCW��j�*#or�}:���${,W���H���I� e���X�-�N���F����Yp��ۛ���sg��N2������W�Z��A���'���HA�I���?\ѕܢʺ���W-98/�֘q�SK9�mU�a�-�K��2��1V�M��il��P��K)*��q�s�5����Ǖ�v#0�.]��6kyz�wS'�u���0�;8�lp��3U��� �ڒ�V@�4�g_3�D=��R��J�:���UUU���!�Yjx:���%oig-fۉ	/���?@�;��Rpla+��m�����'3&�|]��z>^��x�TK��?w��	he�}U�-4m��쬍�x�m�Ұ�V���x�TK�P�ZIK�5Ý5�t���N��N7qϖ.9ɤ�7��@v�n�K�lD��36I�w*�I�?�[A��sQ+rsy��r��5��=K�*a��~dB�c/!j�/)�וh��6AN�m�[�S�&���<m���uqRc4=��Tۭ��ToZ3u���C�����Sٕ��sQ��%ĺ��^��5�b畽mj�Z��x��CyZ��k�>�����vc�á5�1�S�ѵ!?��ܬw�)}p��4�Nw��Y�֓ΐK�ԙ��z�!qO�u!�G�������<��}��ݽ�=U[�12�T}�����ʎVb#���V��$�[��h�|׶;�+N�`
6oC�N�a0�UЬө.����[sS}�K2�F�n�1��A!V�gHs��kvYfu	\
��!��O"�C)Wq�&����T�,��Su��Q����q�o�&'�0�a�������t��6�����	#g �7�
��\8��Q/W\Bkzp^j� �a<V
����w��Q�������g��ezo�\,��I���M���&�0��d�w��ik�sЉWk�UXP��5�U�����>�ҵ�ίZ�%(��IR}����ۅ7��ʪ�6~*|�$�YN��o��*�z#��'�{�����L���\5�B��OQ�� PK@삢b~��c�t3i��=��j%��t�:�R�_�_<k���C�9P�7b��e�-|��'OF���{%����[�_b|C}��܄�EC�s�������o�b�5ם���9_wH`��PZ����M+��[Ӳ�N\V�Õ��Yټ�6���W�/������#�'Ui��c�����-h<�}��8z��6mt���_��Ѹ�HLu#�:��?�>���:	��O��R2��m�����xD;����1u��ʗk�v�p��N-U�WF���%+�ur���BN'�_;���>\�l��*��V�<��7�.U�����U�����8ݳHo!giI{�ҭ�������3���]]w��q�����)jď[1����'��,��7�|F�lF��{�~Y�X�)n�y]��\ׇ� �6Z�vX]+H�\�XIҖ��(���n�zĴ��ӮDi���5���5�FAqo�:3�Kc�֣ǆZtfAr���w��z�m*�X z�*��xpCH��5���Ht&`�ji���{܍�ym��y���r����9UԑY=}R�6��v&xK��R@4F�z9�[|ɛw�j�ґ�g���[��Pje%V�]��8�5��iܟGY׉�EH���]�"��+���: �<sql��u8�����L��W���۷�E���)�m���t�C+�OV�s��E!t'v� ����rNc���^��u�:�Co�$6f"U1Wbr�f�s�r�����\�,O�z�c{����.�!}[Dnm��v�a��fd۾��L%�o��2fX�jv����%�`9�+�3���\�ז�j������+�}7Z�S�e�@:jY�p�扗u���Q����d�[t�,���	Wf�2�o8�˫���2M�l�%Z��*qـv��\a�~#z4o�VNeH-R=����$�U����D]��ᔫ�x�Iꅞ�����*s��� �
TN7�r��G�q.*7�ywvC����u(J@޿�zm��o�<�����Ɏ����W'\�ó!�����O,]�Cd(�u 6/B�]S"y�s'�k���i4���!���m��X,�����ZL�y{�:i	Zܚ>��71[����˃�!l����Xl����q�� ���(�T���֩!S�ڔ{�t�l��q�f�&�e��3 ռ5ώ	�ˌ����9u9�B��b��r�h�W���Wb�6�t��#�(�D�J��ɜ��l��Q	���ԫ�&��a��4�w�ƀT��Y&ӠC����Yѓlv�YWIkr9�9�-�v��G
zr�U\��K&��B���NZ
RA�ۍُ�j���4�sh�]�HF-"3���n��������D�lӝ4勦`S�GK�~�	�u&i�T��:���p�u���}s�]��/sx@��*]l����w0���&�.P��ukL�x�R����Q�\�0=��}�`�ۦ���Z�)�a���5��m�q*�q�C!�ц�b�S���k����	�yV����4n
|�\RYj��v�������E%�oD;�(PB���p��s]�����U�{�"��fd�RY�Y�� �������9Umo\'8�.�"q��(��2C4�X��I�ܢ�JC~"R<�ZAe�'�5�er7��Ԭ/�P��黟^L�Q��ʲ������J��T(����T�Y2H����L�$(�жa��*���
ۺ����B����5e�YR(���L��=]<�I"�H�ZbYJ�	\P�:D��y&�HJ�HQ#�R��I3"$)�t�(��B�Ee�%UQ�0�b�V"�8G�:TE�e!�#���J�NVY����*%\�R��ҍ�W0�n8�kT%�H����fu	5BY��d�R�0襆��B�Jh�*�Ie)UD�լ������YHmK�&�Z�FiZm4B��b'4N�����s�*�2TV��r��ؙh]%���Q��T�aQe��mf�����T�Fi�IT��$H袡���fH�$Q.�iԎ�%����ՙj���"6���Y��HЊVgY�R(��5
+CJ$���L�Ze�bEr��DBt%D{����{�����[�ʮ�]t���I�9DM8�C��N}_�]�w�c��Wz���N+=�uꚶ��w�������$��W��(ߣV�P�T���I��p�D���6~����d��)D��y˝Ʀ���_f=���i:���&��}�+]���wBĲ'�FIj�&�4�F^?�w��K_w<[����/��sP�{��f�:���%k�\��c��`ȾY1}�%`��N�+�������:_i�e���3��x�S���'�O�����޶�r�>e�g�*c�Ҟ��Y�H�U�'6$^`dM�N�Ohq���5�{��i�=m��llʣ���W�&Q�u�5i�s#"q�m���q��rM�>�������B?[f�ڵ7�o�{ ��#����Q���=a��л-��������z!���j�L�{�Q�x�����N�D�qWIR�-�ㆱ�Y��z��P�u#B��OZ����o>��X?�r���OHe,#����5�G6j�H.cd� �x4�,RKy�C��D�7s��aCV;�\,�:y���!9�Ow���9ʚ�w%�m�Y,u�F�����J��Ļ��6O�X�-����Հ3Yp�������eC�w�n
X�sJ��=|��fA��hԬDY��'�G����㋶�^�M�����$�|����]��Iv��v�����^e����3ic8\���S���ih��]��va�V�Fu���^�~��x8�x�<.���v�S��D.!th؃ϧ�
��|�qu�uK�ܕq�ִێ\����شC9���<�C�c�@���,y�\��}A'��<甃Ϋ�gz&�.5���JvB�}E�51C�	/I��$�{����>	woՎv��mT��
jq���p�
<_�-�$3=\�^|ݪ֫KU��5�/>n#K�NNwP���.ݖ�6 V��;�ʺ�ˌŵ"%���^�[��_t5��,�j�SBw�nf�T��n��j��F�q���IƵ�C�=_~�mC�n��̨/�19���W�9Q����b��sq1���SaD�]7Y��z���G!�E[�J+Ӏ]y�f�&mmi� %��k����$-A˽�%g<�Y���|v���7��l6�i:#��X�H��W�̷�f6���7��㖻��ԍֳi-0�-���Rt�*���"*�-�y�r�eBՈ�ʝv�@B�ao;ݻ�r��w'*}U�Q��c������q���VV����%�2-�����TgY�v;G��a+'��5�RʹmJ����	h-Xl8ěܦ�\:��+���W�e�
�־}\�j���nANb�C��bR�Kyxᬄ��=뎬H�ؕ��8�o�Nr�>Z��!'�tQJL�sSy��]Ļ�<��Z��Z���q�е�,�8�HY�邠��#�y���gW���ޗ�A�NR���x�g��5�7��+�AO}�|k��tU$<�^���5�gt�q�]���>ۈ-�z����t�"�)���D�@�d%u�J�w5UEm���{VG%kM��҆�4�M�׬�`�=/
{m�=:5 W�X�k���>��_jG).s_6�:ך�qz�M)�5�i�Ǉ!K�h)�[�.Ï݆��i?/=^B�n����s(Ӛ}2f�D�H\vnv�#jμk�j���=�4Ru�u�.��4ݽB����G�"8�+b���K��:Y�ژt\ŕ�� �fG[(�Ɋ�%���_���L{�VF%�ն���J�N�r������ֺ;"�jf�Ͼ�\&�q����ׂ�놭v�_����?{vOV̍��������|㛮����jʯ�^�;E�����[t���I��u��"�K����pyN�(��B=�&Q�fb��p� ��B��Z���-m6����E�O*�}��}�{��|bυ��񶣓����7>��k78�Lu�|�WKM�����E�W����Qn�|w^��:��R�U��Y썥hp�b��7�<����3ES���n�2/x����X�տ:�����oP���C��+lX~SӆG��=¢�5��|�<�7ԺʝB���J�A�\ӻ�[��X���<�,cZ���&���YoB���S����vfT¿'�;������׆��{�f�rDI��<k�5�k�6ܴv�F�`���`s�S}]~�؋c��ֽ_��;v*Oe�i���Xqͭ�a`*�@�ad���/c�4�Ѕ��3������)��S3�������j�I�/P�X$�k45��l�w-k����yg1~/|�#�4}�	��I��2���Y��5U}U�>�g���n��w�*�V�]����'ƾ-�\@v�q=�Z`],�c6jr��qw��O8�L�}�.�
+?\^ݦ#��*s�g��c�T*h�����7\��ȯ�ۚ�B��FjՁ<���wm���(v�E�-
2�v'S�>��P��� <a�#q*��0#���V�^���G�W>{%{|�x��R�-�h��o�j9�&�q���tE�!����̉��n�Ij��uan�s��Չ'3�)M�͎yU�fn��Xc����i$0c���(�����G'�5����Wo��̅󼝒��c2y����I���*Kf [t3��%`��N�r�ڙzM������CK�_$��d.��:4��|�#~|n��\Lw�E�pﺀ��Z�YZ[J3g4��εu���ά�9_s��W0�D������cJ�r��e4�=�,��Yֳ`v���qi%=�ݨ�Y�Q*評��w7���5�Ц�ӻt�`HuEk���>��KeVz���a:7�-��������I��������jM۬���t������'4T�mN"7N����U���G�r�Gp���Y�ގ*}�1Q�6����o��gQݦ;��*Xu})��\�A	{ұ`��7�C�DB��cm���=�7Ժ��7.2v����=�@��ީ=���2�)X��zt6��D��cdpN5�d�%�|��0����ʤ��]A�JZj ����[3������3X��<���r�

a}�0T��K�"������R�t������x��ZUǗI[�`�1����傯�ںq��$����Ox.��gub��O�]�Am+�,g06�l:�5��.φ�'2�`�="�Է%j];5.[Y�.7�r�|���x:��_�]^�Ǿ���"y�Gf��:m�˘)����5��}�M�KI�\.$Z��8�d�K��\�w��������O<��ŵ�]��ic����F��ӎ*��`������l<'j(zi�Oi����6����:�����^�Q��W������[j� �
���V����,����y,�'�qnQd�U�$�w6X��}�{2�I	]B����N���#6�����eʙ�ވ��V�t��(��~����[ߪ��y�yE��?�N�eN����`��Lg�"�tO�J�{�g{�:���X������Tu-����
�>Pff���u�A�q�M\/nq�c�=_{ٴ������jj���w^���خ��;����C/D�v�S`��u�[T�����4��,��c��
m�j;"wMp'����D�_.-61�|�5<�p-�7L��5ۛ�o�?�Tz��R�6�%ze��b�ěܦ�<u�{�.Ά*j���d��[��v�@�<� D>��TbT�K}�Wg�m�zf�P*�Yp���ԗ��%�֧9D��Ҡ�Ȅ�T��RN@�7B�����]�i�G���ߔ�E�ж��-�8�HY��z`���u,�ׁ�є���9������=Gރ({Ѯx�k�Ώ�3�.����oRᳶ0&k{d�w�,�ͫz�rd��	L���ܘ�о�r��A�twX+�(ب� b�F�6K�2�U(��/���ٕ�<tEr��W�H!���$�j�Q�IXг.�ĩ��N�y����]����yNl�w]n�3.�TE�@*Y�f��X�$�W{�f����~n#���;ո�觌�r�I��\����m�C���~��Z�G%Q��riCZ��'�}''����3�:��S�	���f�FmX{E�����#�m�*ˤ� n�ǆJes�3?��޸G"aRԎ�O\��5)䟹�Y��6)m�E%���_�f��-��U59��MƻFn���H����zg��2ٸF26�1z�k��s�3�w)�|�Ú�⃭��]�tZ�N�x=Ɂ��=;a�Q��%uά���wS_o�ә���w���� ḉؽ�gpm��5�j3���݁+\Fr��|�/�O��u����8��FmX�^��������i:F�;(���z��
���ºZl-tv�(�"y�"�y�-~����ϙ	Q��4&����f�Mhp�q�h5�,�"�
�r3X�}�B62�m]v��e�Xz���gP����ux�T�Jm��S�~yزT��ɵ�;���RT�:��5cǆ�q&�x�x��vu���)�'^$�5"��P�O,�F�;f	�Ɣ��4�\�z���}\�/�e�.ZR'(�,G%s��Q�u{}�����D��o���`���ںݶ���'�X*糺���}n�M�r�r��]eN��Ti�&�{b#zR����|G<>�9}���o:5�Yp�-�m=F��AV&�h̙��[V�v��=F莁��ӌy�ZBN��5���q��+��k vK�fgr7�\3��@��}�8��Z* s�ڷO0�{�׏�O��vl�ezЭ�Q�fOo?v<�}I��!���G^�'m�_o����{�h��|/�-�¬��Q������*y�9�5�=!u ��Vݎ�sɽ�Q�"�r���T
O�Zr�������ĪBz�ܫ�WA����G7Wp�B&����yd�b��e�7�5�15�n5�Ѓ�[�.u�x�	���ճ�=:�~�ܠ���U�y�}'�ީ���A�fӋ�O�=�B��n��U���+{�h�cJ��� .z�=��U��h�����Ez�e>�ѫԏ�]W��Q���{�r�.����~A3q�*�1i�G7�� -�x�{OΊ��c��{C(3]Z�N��Q�jT�h��I}�sUL��F���1T5#!�e�NJ�!�h)��fuK��Z����F�c�^�p��H��攧㶲���X5�ӳ<�5m)�W�1�-:���&�P��/9:����uK"��0�nvM��+{���ݫ��j��<څVn��ʂ�,���<�&�s�xj�N��+��+z��=�fOz��T{=�Ng��j�����a;|�Q��V�2��j�m��q��\�a�yʻu�]�u�������\��@:|<^����}b3�#+�~C=6�6*1CYp�|�w�o���[��ь���i����k��z��g4dt����%KCwn[�z� ���Z��7{�+��
1����Ȯ�ϼ�=��~5� D��U��ݮM��/Y�=���ܭ��o[��B_gw�A��ꈾ��U����zjܸ3�&���S*˃��a[�ϛ���H�ȅ�op��#e���YAb��t�Ϻ;�ջ�T��o6e��U�x�2-����A��'�R�#:�rDn;ɵ�t%b�C��C�`��ef\��K8�ox��ǩ��И���wtu��N��(���l� ���v�Pq_fVQ�+�.
�7z��Iy;���K�P]i���*0���-��<�85�z���AgKՑ���Ǖ��Ra,�P	g2�r���qT����u��l�w�5�Q��#:�:��ͼ�������ƚ=�w��6,]ڵ)E�7��=�z6M�A̰�H�TUՎ쑧^�;��i�����%j��_�d�>�"�4�f�G�*P:���́�`V��ݻ
�=���S��Q �B ���\��;ȼd��\j0Nwk�cch�ꝵ�lШ�;�j���<�֊�w��pڎMk��'{�	��56R�
��4����t�8�J�{\�J�	g����VF���� (f#çi�qNg��8)̉�H���lw1ҩ��ĴC�Pl�%x
��W*SGt�Y>�K�^�*�N.�Ӏ&|$i���(��% ����DgEv#�ĭ&��L��9��ʯܥ"������D́�YEͶ�T��{�H�����P�/rc�'1�gn�-�����as��u9��v̊��
��H+%�pM�nk)��5i���Nv���@L|qIî2 �X� -��b��)�ek����0�j4��d��[:3�h�v���[�������g(��%�VD{^8��߰rn�)��ʼ���_F4����e�;���lҜ2[�ӡ��Sۢ�nS�]�Qq����%̴�Z�J	c�Ta�;��m�T�R4���Yqǎ�rΌ�(�(S�F;!���V�us�1�e�u۩�����vȫ<�>S8�&W7��D�	eR0��ԯ��yJ[5����x�����μ��ybIu�v:;� �\���Q��l�:�^�śC��'�[#��G�� /4�}R>x��jc�M�:G���w 5ñ�K:���]\iT��я�����ě)��bDW+��+l���DS�\i�4�l�Y�#ַ;7pZV3Kx\��b����3,�%��kƛ;3Z�2����J����"-� Rݥ6�;��4[��B���	�u�Bc%���edy|�(�\k��ݳ
�^r����㵮�P?^f�v�u�/�0m��6],���w��6�й��'�l^�W�S�e𷔴��Uu/%u f�Z�>�l��L��(j���^-�dw�V�II�*۵�T���z���n�i񇦜�uε]����<ԂЁ*��M	��ae�2��H�Y�n���f
}�b��g#m�H5�+ ��E�je�vc�dJ�2��w7r,>F�IGplj��1�<h�<� ΡW:��X�{��_�!�E\Â6�'XFUn��Uo^�|�dب�m�Si᠑8W����!�E��"�AhmeEDEPY!Uaf�PШ�1f���"����(+�ʫ#M�*�X����:�	K*��+B,��R�
�QL���\����#��T�B��\"9*�Qʋ��Y�R��E�d�u�3eIGR2Q4,�N�Uhq!++
��#JL��0��(�B�̃�.Q��2+�DG:��+:ER�)���	
 �T\��aE �Ue�J.A��R�E\�����IiTb��6���tL����$�H�:�`i�*�j�êr��2��V�E�h(l��4�Q�&Q'iQX��T�U˪�+MH�G2ڢ�p���f�(��CFX��6�l��p��ִ�UgB�R��G���.ʦ�f��iQ�z���x�����*`4m˕�o�庍Π�l���wS�����.V,�.�n��$�&C��5E+��*��af���8$�4o7����ӽX��ক�w�c9��q̹�9}!p�K;vu�1/K+qsG W��ˁ�V.9\������D�F�Z9m`��XVT�V��8��@V;\���O�ԋo�Z����qi�4�,���d�{�w��.�Jh�����_sV�\���Y��]�j�E'���i��\��<�ju:ی���b�V�u=pծܫk��e��:����,A�e���Nw�l^�싷���x��Ts�u�L}�bm��[C����P�X��Lڐ�s�_nW0�͆�kX��T{ٮQ��3*���v��y�G\�n�cQg���B�9��[�p�Sc"^�U�cվٟ<Aͯy�Ab����y=ܱ2�ۘ	*���.^|�WKM�W���ť`��=�N2��4�ļۊz�u��C������\�ʄ��1&�꾹�.),P@�"0�aL.�ՔIj�!rѦ��N��ш�IS��v�U��<�%�P��"�yDµncS8��,�s�.s�vm6��ru�/d���A<�r� /�\7�e�R�JDF�zFÛ]+_��{w��S��qZ`K�[�N�u3�,�-d���\�p�"��5ǡg]��a�~aJ�+�1�u琼u�-�4	+ǂ��J&����/���->�9��PS��4(������j��9�W��Y�$��=X�֞놱Cж�r�m��AL/�����A��`��>Ģ�����;�[�E���v���x�TK�����u�Um��5_V3E�(7�c�Wщ��Ŵ�;թ�x�5�����3�f�Z���l{��=�t��~Xk"�mU�tc�M(o�(��|􍨫��wj2�M�;����予��/���V>{VE�y?)�q���K�{V�Յ�{�c�V��[.5�9�'��8꿊ܚ�O3�zd��u/x�Rs��/ɥ6z0����c@��^�vG���v�ėWօk����9Ӹ܃�'�Mf=�ެv���Z��C�[��xoX�ӓ�a���^�z
�,�����{��L3h>�^�r�x�,����v��lIV�\���8��}���R��������XkZ��)K����.bkv�wuF�3�b�c���r_m=��֏I]Zx�E�!&Q��R^�os�v��:�y�! ��r�{�͜�q��򵴔��q�m9�qz����!�q�fئ[��C�TwW%����0r���m���9F[��)����'
�.8#q�X�9'�uo^�ʳu�fQW0�(��=뉎��K��[��;"�^�)9�j��G�=����Y�{�	�V9�f���x�pS�s��k5hOҵR� ՚r{���R�ZZ���=�Wk(7 �{M!�����܀�N(Q�R���bm�X��T.����6롱Kؐ�[���ힽ��6g�r,�F�7�����[M���g'��uA�az;YN�$� �e����D��!픴�I��ƻ5�k9�/j՛p�xFg<�n�Ҧ�+����!-�r�N�;г�I�;N�:��<�}˻6�wn���ĺF�
c�]!�R�]*b?rq��l|��n�M���N�u�^�l��[��>w��gC�7��Z΢��aŦ��/�+�L���f[XWs��F;K]c;������q�][q��
��o�Cq�f�_8*�T�N���Z=��˙]ƚ��_V�8�'q�[�BӜ�Q9�&��:;9r��>��kj��ȧ6��!���Oz%�X�<=�sz]]���室�cyc�{˜�6�;v�ĪW���X~2����C�L�2I}�����%���{_o2��昚Mƻ�G"u�uK��*y���Uw4��l>�Ug�0�sv�6m$�J�
SPr��Ū�;ka�+��<d�8>��_u�V�r��<ө������k��S��m�ں)�JX�3���*e���ۙ1��ٵަ�J�ʳ��s�����9�Z:��H5gy�%z矧W���L ����_�aE�Wl�����@㬗��'[�㊉�o�%6�]&���m��b� ����%�C`���n����ss�����)����ۅ]�p�,�	s�YdT�fv��f/I�Ŝ�}��*$�Vӄ��2�Ũ}m6���=Qpo�h������D[z��B�(���Ph��	���v۽s �2�l�0�0_^����N���B� �b��ȷ�B����)�E�S���Txz�<RP[2s$��-�+Y��T�!Ne�J��TI�d��V�gq�����!��5�3Y�ˣ�Zq�R7�yM�v���UXr��TD�2���io/5��S:K���C��o����V�{Uqs�U����n�P�/��#Ǘ�!Eo��3����IE������-y���n����*���g+�1�{ի�KiH�]-r���v�[��kb��9R���<�^�;]��%sֽ�,�G|MԌԉ���n
i_�ޥ��`���uNj\5��ԩ�ݙ����4xU�����,sU�.9\��S���ώzgY/>��o�=��MD�m���ewz'RW�L�W������E���TǮ9���q�+�����7��*f/ܸE���{���Ѧ�@�����K'����TTKe!�D�Hאn~{��Q��o���M��h��Q��W���q�342㽷 ��TH�a��V鿫e��7,\Ls�W=��ÓZ�z�W�ʅ��]���@z��n���{�ţ������G'�\�	�(?\M9��~��v@P�&�o����P:D@�����Џ���V��Օ�ڇ�_F�������`jm�G��3I�y��+՞�A�'����*��Lrv������[\��*2���j��T�{d�Sc�:�S��Cz0k�Ҵ��VL�1����������|��uG�.k�c��/c��'�?~��~6��|vu�ߺ?�a����[ϖ���,+��:,ש����`Tnydxc�~��^�ed{�c{�Z�7�n���m��3�;�Mew����wo�0��JG��&��r�G�i�_bv�
����>��e�������g"��1o>�p�|���g�Op0�=P�"�T������T<i������t\�-[Mz�ә/ݕ���Có�yh\5�#��'�ĕ�FUC�3�n+��,վ�O�u^�>�w���ykg:��*���#�ﺣ��W�x,u��Ȁl��OlD�G�C��P��y���k�~��{%��GeԳW�X��n��;�<_�Ig�=���Dzk|}� �,�8 r	�ҧ6˜�����^>C�I�}���j�����Rs�Z2���߻�4�Ƿ���aޡ���!��݉r�׻s�wx���@W ��E�+�ra-~�8d���Ϗ���~��J��.�:��:�΋����(�)�\M�%�D@j��12�]F����
���Z�-?;`�т}�_����^
U������x��3-�[��'/Qgݡiliު�x�ё]o \��$q�E��܌���к�A厙�j�VK��w��&�RE�ƺ��w*P;E,�쾮���u�K��w\�շ9S�屔cU�-�Ƕd�V�ʉ�ȭ�IOg���68�|߫@��{"m��e@!�8��/��d>9[���x/,K��>q.ZN�O��s�F��R�5�{>f�R�ϔۙ�fe��S��_V��D5����z�����������[P�wEi����9Z#4��>�0ʑ���s�1fa4z6k�StTv��Tg�w����>���|o�W�>��v�c�Ez�ǶX���(�q���&��n3P��]y6����au�6�z��t\+u��DwS�۽�u���;ҜG�X��{~�oML�\���;^��G=yS���wl�{�wL=���4�A��lQ��~�����^����Ǻ4A�����W��}�/`_oyO�<`³��
�*���:��( ��to��1�P����y�͟�T��I��G58���=�5��>%����Y�zD�gn8�ꋋћ��'�������^%2�}�=��Y�Wؽ�ţ|x\_I'�C��6wn��}u��2�0w��q����評�܂���<�����x�/ų����v9�F�Xe���)ǎ+h y1kϊ�_���+�n�֡��.;�=0
���`������jj��/���#"�8#S�7�Ŋ�:����Py�b���SbaK�Q�͵��ڃ{�qo�b�޴nM��u�T��_%�F�^���A�n�2���F��i1�jH����~�y�����HOT�\��V&���8gz=Lo�K:��w�Λ�Qy=����-1�'JI[X
D��ڞ�u��7�$\D��ѐ���U�Y��<��L�{<�<(��bp�z�q�'ƙ9�뉲W��S���R�VеnC��i�>�,�;W�E����{_��{}R6�vĲK��@H� �<D��.�0<V
��~��Z�q��F��{���>���>��n=�^���2K
IjG=SG��C/�kt����T�����>�ѹ�񿵣Q���Q���ȟ����f�
�ͲE}
��O�~��%�{+ ��*�v��9�g��
�s�h\S����T��r�H����Z���/��7��j69��=�)T��NWoR}>�d�a�U|2c�b}�*'�oFS�i�ݦ:�ކ1�]з���E����~߰���g^�O�	W׀���~*����ąM?�B�?6φ��{~`wIf%)��u>�;��^�|����Շ]9�U��yR2��d���#uW���6Z����ʑUiO/���	���STpu�ݾY-�\1��:F����������f���*�C�w�ҳW�N�t!�b���#�z�x&2��".���>�}*̚Mv*��w��g[���ob�Nj�*h�Vt�����w�>;IA�N�6�-Nm�m�%ńό���O�O���ޝ�����s�r����]����?g��a�r(�S3����Ϡ��%���P1yTy:�~>'�u�P��S|lz�p(��:wm��<�"g��ģ�d�}R��4�yNl�^�~9~>���<�Tn��z�f����0��sU9}�,�����Jve�x�u3�o��e���}~\k�S��^�U}���G�k���C����~�5�1~YS�vx�����
�$��Euׄ����<�>��z��#�]������o����y�B�}�[�:�A���3ĕPf	>U��ee��>5˻U��&s�V��7�ʿD�y_iL�9��{������mǽw��l�Q@���&u�}���۸Q<�41��2o�u{Y~��V9��������ZDxߊ���}���ۯU�6�Ae@V�n���zG�=����S�;�=t���|3�#z�!���0={IG�wI��������Ɓ�u)����B���^(��#�pC��x�q�N5���	��c#��g�>�βZ���F��
n&��������a�ug\��"�����v��o���i=�O�up��M��n����X�����&�y�:�d|�,�P�o:S���2��e��ƫ�Eo C�*ҩ��nH��Ͷ^�J�(�R��nﻩ#3�X��T�T�d�36I\�L?�@��⸖��0����F�[5q��_7r</�Wt��j�"&��;��-������,Y�h�� �)d���7���<\�E#^@�}:~��S�誑N:��Ww�v��+�����8�>fhe��ېj��P����w��7|O\�{�<&9E�~�J��E��~���onB~�G!��Q�m���vXC�3{��Q|�Q(g�m�����<ƣ=#����]>'�wK��Q���1{�]����'������36L���5=㟆��'������fKt���q
� �B���,�2�~�^�ed{�cz���[f�߯?W�����9�Y��yS��'v�3ʁ>E��ɭ7��i�X��B�?_��vr�����;��+�YN��u��<�3�gJ��R��=P�T��[���T<�_0��j��t�J1c#��>^��χ�Ǯ����^Z�Ԏ��$0pO�������5)
P�t׶�u��zV�tO�g�jWq����s}#��{�=�9^u����]9�Iꈙ`/�����Y�@�*Z����梩����o]�g$�ݹ�&��9��j����˭�� DRY纈�E�A�S�ge�&��-�by�q1mɉ�Z�ܵ�h<d�GCw\V���mf
�CD�}�;��[��3�b*��TfԬ귷ss^<�j;Z`�N�͡rs"	֤7�T�ܥ��V��^y�`M����	j�T�B�H,�a쬲�<��+��kRĩ�9����Z7b��CN�%F����6���}��X�Js(Su�vC��-P歅[�ML�J�z�Q������ ��\SIq�Xo_K� �
b�Suv�.��`��z�5"��:ך�����}�oǆ�=�-:hv��-Z�Kd�Moc�k�*٫*���s�Rs+�vƷ �@�g^����ʪ�(�k��[�ثw�ow���w���*];V)y��a�m�d�Z�2�Erʴ���7Ĩ:83S�C{8YhԆ��c%3�f��M�m���gE[f3��)��&��)���R�;�kl���]��ew(��M%nHT(v_j�yv��Y�n���v\QAN�mh�Z��2�L:w�V�ĭSp�k� ��&� F����+�	��ᖻ#r�qԶ�N�3�P�v�����.cF�r����f`�����B�6�CX
�z�ugqbM��捞��IP)�G{�c��l�q�c[���/x��d��5�=�o:ݰx>�U���ߌ9�#�4�>Y�{=nΎ�nN[Y�n���Sq���8�pX����5'P���{��ڰ��]�m\���7�1ld�כٜ��]l��e[.�5�˘�uPӻv�HlL�0x���QX���J�A��v-��U�ۘn�PQbo%t/+��l�V���Z�v����K~&��-�鷣F�m�=�Y�f7��YTy�䑬�=�Ff�o�Ҷ��z�ݍ����Uv�T�0u�;w8�����\��[}+W\錑ֆk����ְt�]�c��ږ�}ͬ�V/�*��ч&s�k;M@�'D��*v��E�g�#c�>Н��^ ����+��@��ʉ��w���LY��9v���i��=R�9٨����كn���P.v'h��I-���0i�c��?.�j@���.�\���{�0dOR��xʾC�qؗCX�É<�j�JL�����^ۘ���缎���k��0;�>��m>�Kt�s\���*��w\N�p�z��N*1��s����3|ӂH�m�Ǟ�ֳ�w�n�oSck��IT�7�g)v4a�������U�Nj���D��c�R�z���)�p�'n��r��U�LĴ,ꄢ����4r��Os��]\�5�咍�E���׎e�me���"�;��]����7�V�%@y����	Qq�����zF'��ù��n�n�ò&�H��iv�'�@�}M#�L��HL�"��.Ii�"�9�Z�Us�$�˕E��bE��V��H	�QTUIԍ��r���B�*,���a���4���Z,�JKH��Ns�%*�R��B�P*έ5
M��L�ęTI)�2� E'3��f$�r�2S����TB"33-D��K�.�b	a��a��iq�'$�50*��鑜�V�h!�%����.�Ҳ�U�*!A5,�J�Rr�L���2S+KCXF"�)�V�T�fp��)��R��
(M��!��	�a�jR�%J҅
��E�bjI�����dj�GYaR�bԱJ��+���2� �2T4���͒�Oqp6�*�%�����IZdt�Y�D��B�3eʸQ�)0 �2��+4E5�j��D�\�fAID�E色�JģN["��B�&��'V����?�_�z��v��u�GT��F����X����԰���43 �xhʏ�b��.r`�{j85�2�Ry�kǇ*�U���W��S)�˩�n�M�w�9ޑ���G�K=~�p�=5�>��fW@��~�	p粧kkF<o�3�L@r����C�]?���	��z�џ/o���ޑ�����M@d�Hm�;�&�=	�]9�3����8 s����[�"���9�K
���C�D�����7u}>4EMo�K�Nױ��*'ѫ�'L��D�K*�<LOҽ]F�>��*������N"����ft�*}��b�h��H��=8>�� >�\Ks>�V����"b_W��|r���'���]Tf�|���}ύF�/+���HdG�x��k@�wLSng�%��S��m���Wq��M����>�^��L�ei����{����^&���z��d3T6�:}�&��*BUu�G�[�7z��ܛ���8:�}�E����ݧǕeC��v�c�Ez���{ެ�eR��Z�}�<����s3�ѥ��yl��*}�B�<N���Ǯ;n�x'>�����T&�R�s��2=���O�K�X({�yS�������/P��r}Ǎ:�w>�lQ��~s�C/j^֔=�g:?����K�oʗy�G�\�]�r�.��\Sz@�1á�%˔]Z�Z�r����{dT#xݼ�����#g�K��R=��$�:����i��X�������pS�!%Nj���v�����A��d�#�[R�U�W�)�Q�
k�u�P���{k��^`�5S^��uc��d��s"ҟ�fa��PM���S����m�廐f�^�QO��5/Y\�zL�cWJjtw���B�NI�>%ٗ���T,����^�	�h���r�>��p9�.�>�'/�ݾˏx����R>��֫x�%�� 	�L��~�6�َ��OR�{�x��P�T�s΁����Vq�x��C���z�G�C��C�[��Ǵ*����Z2Ͼ���3�$�R���K�����k��pϻ���]_�Q�����/ܫu�#�?z��ǲ�e�$��,	��}-�ϭ]A��M�	-���/ާ9q�.u͟VkS���J������z�q�'ƙ9�뉿�^+!L4K�A��썯9���ů��~�;�|�|u9Ѥ��o�F�W�؛s%�B ������4���PYa΂dFg�O�^�r�T���Q��kF���O��ȃ��>���z=�^���2K
Ij}�����u~%� �4�Ϸ;�9�==��_�:΍χJ�֍F���W�>D�����`k�d��NªF�3��?V��5���8Œ�YL9S��3�Qt�#���,�&��4��)�jVӨ*�9H���ǗtZ��ㆭ-��R���V�EtNJ��g�Jw�u��'$��<Lյ՝bmN{'���;���:gP��[�su&!�\��y:֧�;�w��~)W�c���Oxи�J�W�j��㗪G��Wtb�^~�F�~�@� �Zs�]{#qs�^����I�g��a��'�`���Y�[��_+�7�V<��1u��80ڎ�ԫm���t�'���b㽵 �O�Q�h��
�պm\�>IW�����CY��<B���3��o{���RE��xײh*�of��^T���N���v�C��#�W)�w�nϳ#l#~�hߝϗ�x�ү��N/W�����np���I���:v��x}�=��W:�p��r�^Q~���p�ԦJ:O�tb��DI����s�VC�K<�Q�ә3��������<�x��Þ��2�L��*]k�<�I`%��~�:~>�>���q��Z���P�>;�w.���W3��Y�)Y����,_�3�n:�_#�i��q�=Lozϻ�*V�F�z&m�2r���+�u�g�k�������z���*��R;]u�/>���8��k�ύT{�z��žC�D�w>�Q�޶=�m �\�j�J�0�>�-���3��&���q�����k���}�1�Zm��:Ŵ�8���i�-��1C�<��WS�*�Yۙ7������enǍ�mF���;/�F�t|_Z��G%��N�ѵP&7���-�g�\�ss&���ށ]Ř�'q�rՔR�d�M�KZ]iY֤7�@���J&��R]q7�~Ӌ�<�=�C�q�U#n=�g��.��9I���;.=k��Z��FW�@�=��V9O��n'޴�A����I���\��M3;dR��9C�.�gj��zҨb��&@��2��RѸ֩ȗ�l�g[g���{޸�pw0u_�ų�N���>iu�40�ϡԐ�t��%yM�=�O��j�m�������g�<qmO�8�;,���CZ�w�q���=q7Ϥ�&��b��z���kuS�n�x��xD�U��Z�mw�{�K���f�@���{`M�a�Y�RDO����dν�/��aI<��|}�.�c!��ѿ���uo��8�"�}��O�P0>;����7��0%"DkL>ܜ��+�������*|����}��}�,V���e�G�3���Q͊��4=�����j�(�1ށ�¸��co�u�'�q~/��W�s^����{Wq=�^����j�z��S�n�������Z3�ȣ��(:�l���NQ�A�^'r5Ss���C�~��#��J�/�X�9]i(?�,��G�{�oeJW��t�5��;�Q�쨕�ªk޽��:�,�l��0ՅDY���I���Je횷�����i�5_wD��h��E�ef�d�0��+V���ݙ��;�����tk�q_3w����%`��&������܇y~���b�o*t����	�,\VMi�.�M01:@���5�`莨S�i���ߴ}�^�Y�C����H^���Cĥ�a�3�}2�����qs��bzn�l�V]ហ�h�=�����/U!�"^Z�Ԏ���O�U��$1h�H��հ�����G�[.F�����W���G�܈�\{�r���dC��@6K�s����N��Q~���U-�Ǽ��
������.:��⒫m���H�|}ĳ�ڮg������J���o蒮Ś��������3YP��@�m����}^�!7>��������u�MԺ>d=�g����%��ߌ{>'Ɣ9T�-��pJ����z�hp>�;��zXu�{��q�u�Eվsݞᾄ���{��q^�\M�%��D�Ozz�Q|}�Cy��L��0��1SY�d,��G�!�|�V������G���.'�쉸s>�����Hȗ��#b�c�|}��w16.=y��^�.���3�fc��}�z�>�� ;�ցN�_)�3������q1;;��Fƀ(��;E�%G�]{A���H�пwY��J�((}iݿxK�봽�CA`� A�f�=��2e'3p]E���4ߎл��4�JԨ��;gFR;�R�Z\m�}r��=�V�Q�(���a^�eAh�6��v�]CD̈́,M����>��?~��S?1�9��{=�wE�^&���@w���t�fN�z7��Ǧ�f)�>�7O�Hz8����C�9�늕�D�gº7i�W�!�]���^��.�V#}�v\�o����ﴽ3��d���_�kC��87�n��ϻ��\v���N}�����*��:k�w������m�\��8�@�z�N�u��6iփ���M�����R\W�o%g�:gkA�u��{uc���m!q��#�9�f��T;��ҳ��JV}�~���˕��g���0F{�ȸU�~����G5/�tr���B��9'������=NU�Ĵ������_�^���j��l�tϠ;���7�r�}޺�x���7}����rO��
2F%����B�I�L��e�T�Sޠ\��悸�.�7�2��{����w��wy��C��|UGU{1��&t+3���A�3�&�,\T�B뮽.r-��:�^���1�y8A�j��՟�y��kz��<h�G/\{��o�{ \�i�$�X �H��mM*�>��~O��+cw�vHZ��WWZ��έ6�R�'+����t�1�7~k���հ�I�޽�T���x9���ܫv�Wnmp�����L�h۠w*^��ܤu��%�>��� �s�9���3i��(h�Y{�GK2��r��6H%..+��{qJ���@ީ�#y�ٲJؿK�C[I��w�i���HN�z�Q�.O�2 r ��<J�Y觻⳻3׷�U"��������ڸ��}�a�W�����߷�#g�LK$�H��$P�Ӊ��#:Yһ��X>��/3ƣ���Ѩ�O��7��#�8n�G��ƭ̒�_aP߃�I���yͤ;ƲF9b�S�:7 t��h�m���Q�z|��Ϗ�|O���ίg�W`q�]qS��W.��#ї*Tٙ�v`�s�4'�a��O��/T�{ʪ�r���>������gK�1�T��˵so�MF�*̓��z0��>�����Y��i��U��g�����Zf�{Z8���ޡ���'z!{"�G{*A��z,���a\W�t�+���{&=Q^[R|=K'	�^u�A��{hb�W��}�5q��s��+ʑ�����̘~��u��WTNoֈ�O��p�O2t�>e��j�1�W�����)~��1}[�\�U�YT?�h�7x���z�^!z+y�j�-"��ʭ6j|�G#f\
�^Wȓ+œ��̧�Q�����)~��F�H��F𛴝[:3�Wؔ�&�=8ſ��Lo;��cC*��H0��Ŧ�tb��-�B|T��`M�[�t�u�+4����<���Y�%-#5ms]��*�JYx��,�Qf�g:����fl�s���4�@.�W=S���$��ī�S�h�L�@K��]i��ٖ���G*L�r�g�9����>������w��Н�\jʞ7gĤ��/��7��2�#���ϴ��$$@ٟ_c�X&�o��+��z��=t��C��bᬩf��Fa������H�T�Kׂ=��
�G�9��n����q>gr=�C����qs���%��U|f	>U���^��|�9���>����u��Kw�9��9��Q���U#o޻��Dd�� R��p������S���;�=�xz�|x��G+�Q��RDxߏi��'O_��\����lϣ�<�0�cÖ詼Y��}
ӵ2�	�`�3 )h�R���~��g�����L��/*���<�	���g�]�뻅��H�I�d/����Y�����#o���W����LH�W���������D�&2��뉶g�Th�����Q�-l�����ݾ���&j1��f^��o�X�v����>���ϙ��*��"�����\�K��7�Y߿Ai�n¿�W�X�oC$^~>U�ՀwD�|ÒG��k�WHW�c6�eӼ�4�F���s��h���z�T�,��὎�g����զ�q����;�e���CR��C��3/�yo��Rw�9#lv���2LQ[U�ulO��^d�Y�����Z�n�+��u�����Q�:�7�=� ����c3C.;�r}
|J���� �|`����n;��(�c����ճ�>E#�/��ۅ���}��n=�LW{�t9l�H�<o�V�z���h:|\��6tz����t��9��n;m\{%�{�g�ފ��Wq=�6+�����;^���o�Y�o��Y�ۙ�?P���(�J����������T��!�XqJ=ˠۨ����˿>�m>�5�[T��!�~-3*�.�kM��@yf�`d��Qآ�o�ȥc{�Fo���Mg�߽u���-����#/j����e{���׶���y# y*[�FGp���	�{�5A�di~�.5����s��q�<;"^ZbBJ�P�	��p��Q��z�׋3W�J�W��2����p:�T5���9�/s�q�)�����y�d�3��̸���fF�Y���I�L�T+���:�e�����n�ǼG����Y��ڮ!kYyf�o'R�\{��~Zr����B�����t�r��Bn'޴4b���3g�Vs��:�}s�K�����h���1ws��1�{��ŋl��me�H�4��s{��tV&,��7�Q�w�*�I��Pɶ�I� �X�:,�EVy����;���Abg�}Ԙz�����Ԛ�0�)�cbe��
���%"�^a��������s��ه�.K5�*2��[�"�^S��R½~�8���ž�W6}
զ��{������>����u����3%��D��1q�]F����m��u^�V���OTF?&�F���;`{҉���ɸ��Zϳ�ng�5�hو����HR���^�3o+>�S?�w����q͚��m_�߽�@�#Ƽ �g��h���)�3�4r�F����=D���{yr������_�Eo�)����=���y�Ѹ{+�ѿ{�{�ތ~q�����\W�"��Iu{�ɳz|r|:ǧ���E����|yVT>o�h�>�W��Ku��u�����4����+�F+�7�3���QfFN��t*s��wS�۽�y,����f�^T����x���y�9����X�yS���wl�'P'tø��q�N��}��Ǣ�g�yQM�Ԡ����2�A�/��DyՄ�w�����e�pf��C�d�c��3�� !^ʙ�ː�>���%� ��:})�>��TsS���ȏ=�/T�2���xk��������?~GjRd���h,A�km����=a-$b�8�b͜m�V�Ʒ���c���z�O��D���vI�wJ��\�+=�:�۳1.���n�0�t�Z��Τ�,�{L���-���Ai��]���/�6ɺYZ:�2�z1}�T盳5uK��_h葐��)>�Z
Uj\�O�1toN�`���f�}"Y�_n&�]"<��-�<��κ�u��h J�$�/�j�GoQ
Vc��SB��w�t���컘�:��@���R��d����5�[�ݾˉ�E$N�}u�O��g���"*"�.��X$+�f���o*'t:���#�`���!�,g��9/�w>Դ�ݜ��ӟ1X�+F���j�n_�{Y�]�C׻R�(�`.Aʅ��v+WI}�!�V`��j'e�*f[ލ]�KI�+�vos������wXO��L�wZΤ�"�֓5WN�t���f'�؟^$�#�Eœ������ш�a���կuJ����C��9�\��1��k1p�9�V*����1�QF�Q��4۳AKI���b�B���x�!��	��v�=�E���zX��(s��R5k�^./��.
��uʠ�ƺh= $jn����݁/�����Ѭ
�O��S&��&��J�D�����Y���x��W �u/M	B�.Hd�L���\ۓ2l9�>{X�D�K�f�R��G2�w�G\��Me-:#x8϶��J�c�idȈ�6αP�
&`�=;�S|V��<Ja
V/n�7����.P��V�p0sO#�V��f�K�l>�����A�<�Rq�ۭ۠A�ΰ����e�ѩ�5_N�Y�v\t�}�/qE�n� )Sj�L�*������A�j�CrwV��Z�@���6��rG�]?�jx�������N�U�ը%�-�3.!mH_0�;��:�e��a�i�W�D��ܗ���{Oi��[Bp��h�r�6+U��c�k�3-u�vL�#Y���g�ʃ}�=����W�P�`
�ovtA4�5q�D��2�
KG�5��:��k��"�E�ݣ��{�r��2����7����x*>K$m��a�Ձ֕Q4��"�����1"��պ�eb[w�q�)%�+�fk�v������k���]�i���0u�Cb�`bm5L<�ƞ):5v�8��I��wq���{8�'�`Vz���}�Z��Qdc��һ�:�^�92��8=��Au;n�8�Y�Ej��.���{�pE���a�ŭE[R�\��T���*]�`��:g7I�����/�on�cV�X���ܫS�!VCO�z�m�V�s\�����d{�N���V��"c��p9�)u�w:T�.�[�w(D]r�=��C�G�,�����SVd�p\]��P�T��+�Qj��zu���qe^*��Ɓ�sw&GYy�V��*c��=�K�y��{�����9G:�)��N�VFDTU��2���I�eZr�҈�]V�9��C�B�H2�+d�j�%c�PD��2���Ե=<4 ��'Y�-]ݸe]K+U2�'�e��j����Y��=C�D�.!!�L�%5�sR�2�U5�e�*��S�̠B2���6\C�-E*$�,*�YR��;��瘘:�jdEXEFV.N�j���N�g�DH�Nr�B�=�$���hF�#���M5j:%8�D��(�A��RR�����V:笐�ZI�(PIT��i�-u���IJ��(N��e��5N�h��TVa+wCB�/M��j��H�I��wRpN�z皴Yb��a�)-rp����G����	=Я+0p��#G]u���M�ؑ��EeC��߰vT�C)f�(��\0��gV�����B'�&�MB%�+���=}@K޽���!ȎH@�r,�u~�x���������>�i���z�=��֮;����w�$��nj�/��W����ޙ���3��L�LO9�k�
��.�8�2�����)N��U�L{z��+���4d�9��3p��,�_I��'�|�*���K�nhO}�����Мxʯ���*/�Oky����﷨���;�s3�1�Yp�U`O��H��mNDZ����zKG�P�ٹ9�J�ne{�D�ף��+c�CO_���7�_�=����"*3�n��[ٔ=�V���M�2mw%o���U�����O����W������{}R6��lM���S����A{/=���}��W9��^�`��>���#zѨ�O��7��. �kA���z����]s#��� �}t���Hy���uI}6\�2�HU�T�:7K�Z5p��Q���ȟ�����}�����h}w�u�њ��yƴ��W>��30�X+�s�4.+Ҵ����z�z��Wtb�T	���ב�S���;��G4��f�b���&�d�|2a���a����s�5{��B��L9���C���tdI��Lb���[@v�4�5�����AԂ�W}�i��܋a(m������޷G�{�ϩo-}q�:m��|��m(�+�:�Y-��Up� }�9q��[�O,ޚ��Vͻ:ѕ�*��Gf`��˧��ʾ�L;���+w��+��������M��>z�{"�Dw��>'�d��;��^��їV��g%��Ƚۋ���[N�����}�C�P�l�u���uX���Hˍ�N���~=T\�_�e�����ٞQ��Ӳ��K�t�j��}����ϴ�����wQ={���rNS�e+��U��ڇ�8N��:�eV�%x�n2e����q�SO���W��Y��9pJ��tL��h��}ܶZ��9�:/��:K�]>���4�yN��KK�ʓ,v�Ǽ6�G*�#^r��Y^��q݉޳����,Z�g��L��!���>�Y�ۃe�NGUl�yF�����C��z=t��9�F/沥��Ğ�*X芙H�h����������sj&�P�~���{��`_o�|��{�����l{�|�i��L�%Q�p30ow�i��{�uyD�EH:�z�w�龸����r!zG��G��|}�dg{�~�l�"�<��_�U7[�Z> fϾ��H�P(3��V2��%O�i����~�������i�ۜ�^��;�g���ڛ��4�ej������fFE�'�9b�fN륃tu�44aXj�(r#+�48������~�%�LQŖ��X2vT븜�8�Q����Ԕ����X���ԥ�?w��r�xj�;�H�\jgoZ5:��R���L� ���]D���q �3>���q�R��m��>ζ�1�U+�=��6�ʯ=C<��F����w~2/�2Y�RCQ�FD��4.����S��5���/vv�VT'�����4��6���Dt�e��β^x�l
�{=q6��J��{��/G��gݩ��ۃ�S~=k��kt���W��/G>�\?+�n|O�_��n4
�~ˁQ�O@!�Ϗ���sg���)�*w���O��v�j��^���y�ѷ��?W�����ˎ�܃P�įZ�<��<��]rod�[�ҿ+�?�oh�)��1�Rg��kV�ϡ?]�����߶��{�Öx��e�;C_���9��l�Y�9,(ӡ�VW�ں|O��q�j��.k�c!{�]����s��tdy�ZuĿG�{����g�?���L�~��·qS�t	S����L�+�����<��q�zn�9�+�=��k=��V7�9�#��:o�Y;�ü�>E����pi�UdKَ�7�e�mw�{��jW�C��~���+#�Hw~�Cz҅����U{*:�D/�]��{[�ws�G(E��l씅����+~[b���v�J�ߛ��.�vF�� ��5� ݒ%��:�n�Ju�|������+eKusu�9���
��.��B7�	��5!��\��j�<��a�r�/C$�t���/ek��UGuh��]�ԏ荷@'�j�4��Eƹ~���|=��]���/-���w<I�]k��ފ���e��C�O���uўFx���n�GW���G�܍�Ǽ�+μ;m����<��.z*�����_�g%�Dπ�	T;��[�Ꙕe)�*<���x���J;/T��D��͋�wE�?9���|��G�� �@�>nP�WO�+ޤ&�}�CE/yQ��=/f�QJ͜�����vBR4��=���׮ه��J�� zAo���W��,/{w��/�RT\r��I^���ԇ����~��}���2��O���Px��^��똡���]]�d��]��Iy1��k$hOΘgޤO���'��V�}~��O�W��h�-y�Z=�@y���i$1���F��;W�������7��>�{ԁ�}�^ w��k@�t��>[��0�>>�ԒA�3��fW͂�pWT��z��^�{Ϊ���&���P���9����GRѹ�\k��&�Ǌ����=8=u+N��{^n��q����~�F�2�th�~��z0�'�NwӔ�|���oD�܉՚@�fp����&�FȬ^�!\��X����x;�2E�2`�e���K��N��=2��T#gNj�7c;�%��NMs,�6�p�E�unu��M�T��w[�ra�U��]�Z��n�JJ��er��{G�Gl���ٸ�>�8o�>%PɆ� mhw>Ӣ�[�'���)�Iګ����Yy �����p��K#~c�,��L-�<s��ʭ<N��U��a�Օ�6i{޶��I�ؤ:�ur�@�B����x'U��s�����9��w�<2�d[�>'v��<%ߦ	{[V�{OJ����~��j����Z'��MY
�Oޓ���>~t��=�.5NI�P�9�UΑ�*�d�no{���=2�їP�̣�s�g>�@w��W��N_���Q��uF�GF�t���t��.�ϫ�ǹ�F	&m%�������r��<���*
�K�����2�[�����2��-ݕ�W�vC��o�Vf賈�e� �.�R�>�=mՉ��}hTEx�E�j�Qi�C�B�7>�Qg�#�w�5�1�Y�x���'�R$Q������8g=�>֠ߠ�RY�A��`^��=�F�{i	�~�������2 r�3�)gsǽE	٬��p����q��8����X��ϑ��Ѥ�#�ꑳ�'~s%ϓn0D����m\���v���w��o˸+H���Z���������}�}O=ȃ��@��vEu�Û���3�`��1��B]ܧԈ:'YL�`���9���5!�]���Ȥ��m�{g�!؝ĸl�z�{)>3Y�j5�π�	Q�u᫇�dP��w�M�m�w%~ fO� �:`���/�h��Z5i��9Ӝ}��Z�޽z�;������o����<�u�5�ْ|*IJG3�~�*��Ѹ:_����MW��z|��Շi��$@���rե�'}���)���P�}=6faz¬.{ƅץi��T��r�H����*�@�VN�zsh������F7Q��p5��j68�̒�'z d���1Q-m��s�5B7���:2'��R75��r��w��ކ2�wB��������O_��*;�R��2au�����0��55�r���#����\��[	_���oo�9�qO�CƮ=�a�N}�uX���H��d���ٳΦ	�t��Kϔ{B��:��SF���IӚ���Gm��ϝU{����^s�y�D��o�8x���:�r��
���%��'}�������.tzⲫM��J8K��b��|�i����O2�ݍ8S�Q>3���|w���ޣzs&t&Nؙc*�'�tlt<�"6e��K��t��#�7�4f=S��Pv?j�xG�ʤu���
U���v|JWXʀg��L����e���2����ߣ�/�p;Vt,�������v͆��S~�K����[�Bn��Ŏ�n�T�H����`*�9u��kҶ�]�����͝��N���AڀP|�c'V�Ft���cw;�3r&��6�S�jƝ\s������/Nk�:e���n?�16/\z�����+�({�9�F.ʖo�<I�3ƾ2�����j�����V�����=|g*P����X��Gz�o���{����[��iK;�<IYO8d�=�����Yoy�G@�����-��������\Mķ~ӟ/H��IJ������W���	��rm�Ьkڗy�� ݚ�<����o�Xh�E?+���z�9Ӟ+���I��P��_�D��ػ�u�C�S���8���=���3��ƵHvD�[f+rä���hV���'���	�{ߕ�?]�ȷ2Y�U$5$d��4.)�x�@S��#��^�1jU:�?.v�>T|\zgY/#ƣ`TG������g�Th��/��^�]��J���7���5�T��:���uUy��>����f�@�~ˁP��� �zy����3}�V�ѭ�Q�DˊWo�%���?~�[_�ߜ����:�7��P���i�fhg{*A0�b�~��}Y�$���#�.s�z_|��7��"��/� z����1]�qP���eϴ��06�OU֮ѷ.M-� �lUmXc}3��F>��SZը��U���W�zw:,�{��t�h1y.A5ڮ��uK�5�$m9;d8U���O)u��j�{i(o:��g熁�WR����oy��G1CQ"S��Q7O����9nX(���W����++�n��x�wK��q���Lmw�/7\���1q���9�W��+���O_�^�fp�#㳷3���l�wS�t	S����L���9�w<�ME_��5����UMd��n�og;�b��M�,��3+�>E����1+gX��ދ�����,��4���z�"�W������=���?m!q�*xݟ���xin�8E��Q=�f{ɨ��/EeV�N@mq�G�D/�����s��~�Cò^Z�[R9�<S��ʼi���������J?�i*�e$g��q��O�>�i��H�{��yNDW�xw��^(W�LNM=�˶�����U�&4� �~�^�i{ʯ�m�7O�؛��߸�w�x�>Y�P-�)��':2f�o��Ɗ�/\{��o��P,�8 r�2���_��
U/�E{Ԅݗ��W��'0\圇n�(��]�K���#O{}Q9>�f%��TdO�}$Y+�pŲ�N�d+�'�}�\�{C�j��>�3���c����'������İK;�P�&3�w�x�2yGw�R��*1���b�Rޭ)7���w�
���Ĳ��61�����ڙ�XiǦ!zͷ2_^ �錄zEޭ��c@��q�"'9��7Qæ���K�3Uv�y��5,6M�Ԯc���^��1ލ�+U1@31u��*��y���O�,����y�X?�����Ty޵�4Z~v�|}�D� zp2}�N�>�dMÙ��z��Y�<�Ω���^Hy
��;$���>5���f�[U�)�ԁ�G�x��f���2ױ�M;�$�N~����|�����,�Z�K��7�_���CU^6�W��Q�~��Aߤހ��Ԃ��!����j��9[2Q�T��:ǧ�*V�Ok¯v��{p��C]������
l��C�c��W�߶\	���l����|J�0��6�;���
�q=�����r ��5����Z���Wz����ϟz���hN�;�b��Nfi�N�Ni����yWqZ/'d'�@zl�m w5Z V��c���9��yz_���+����yR2���َ�&[p�8�
�obQ�Z}�B��Ӧ�̕����VE��?zN��9���H,��C�D%{�� /N�N1�.�ڲ��n�,�'J���ܨ^�`r���)�u0�����0<𽌊Zy��_���S�x]��z�eT@���*g�c�ȗ8̎Z]0kĳ7�[��-q�澕%X���J|k��ݙm��4*�?{ޠ@x1���	H����ƹS�at��)����X��r��T�U��t�$��n�>[(�M�kn=�Z'��)泙an�@,�V'N�a�@֖T�غlq�/R�Z��z���ʑ��X'wo����g�oO�W��{Y���Xe���H=Pe� �.*U!q]u�r��Z�^�`恶��\�O��V��q�c}�Y�yT=Fq�~�rY�g�*��,	"Fv�
I{��7S�b̔�%%���E��.}��#�[���^��+c�CO_���7��~��@�>5ȁ�@[����Q�s�;>���h�: u(�1�~�*�#�ʢW��,C �+���W&��ꑷ�%��^Q�F.͊�����>� �$߫����!0�Q���O�����>����pɓc̋[�6�ߪ����5nd�)T��o��D�K�HT��G��֍F���U:���
����LNm��ʾ����:}���J�k �sl�_+�=7f�M��s�4/�J�W���׹�d{�b�辴���E�;U���~�Fߧ�;��F�GO��(2{`d��>��K[z&詌g���ay�![��祚�:7�޻��7�}!Ԩ~�<�q#~�a�~��ʌ�סd�WE�]���W���zm\����W�����꼋�H�ڰ�#�갪�E��C8|ϮnM{wu�Y�i,��BƏ]�ų�%��=���V���X��:��+"�6,�-�K�M�^�n�V�3�P��퍉����m���5�{����1xq�A3��4ƶU�;k�Y�v�U�R̛jřm�arX��7�V#�JO��m)y+ΑR� �ì��{7/2�[�g�w�Rmwr.��-��
�[�Q����v�U�WkhZ6fR��S�j띛]A���qƥ��L���������Vv��E.9HX��V���F���]CC�!H�u�\n}Հu��"�,"؃�N�
���AZ�	*eޅ��	Q��9yh�,�1\5;���F�{��d
�ʚO3�ř��k�t����h�V�T�Y���<M����j�
���]�',m��̰�PЈ�{�]�mӧ�m�4��wQ�v)��g�:\�]J��i빪�����WՌ��K�#��Z�F�f$� ��p����	F���878Za+�75<V`���^9�Q�h�P�;!�<��s(Q��k)��ja�Rl���G�L���YÂ⥆�a���e�˞�C��&}��5;4ʠ�kB(<���]���-)�D��ծ�EVި�)r��a��,+�:*f�Ӵ���u%mB ���Y��U6m�v۽��^p��{{���5x{/��R�f>��e;���:e,=�4,h۵�: i�fF�g��'PJ�n�}�{���{+&��`�W:�����F�mu�@j�]�qf��!u.���h�%J����	�R�6t�����֣v�V�7��X7�'+�f���G�S'��Υ.���6j�=�w|�nm����FՅ-,�Sٛ�ăV��P]ߧ^P]�븴�/�r�.����.��֔��� |w	W�w��q`�z	Zq�'6(˃�0k����xUռ�ef�N}!F���^�lJ�Gu݋���X:�����Aj��A)�MJ\�D4�ua�i9�ZO�!aM�֙���rάN;H�2�nj���pq��8V�W5�i��:�4�/(���]���ˆ��n};u�sK���.^f�:�.S��iلw;�MYVR��j!�v�Y�%�+���X��bmp ��]c��s+;�,�7��f��$��5����K+k���p�m�s�rn�q$��jgZ�*�¥^��k{kS��r���S���8�NowB��;�[N�����#Tkj�M�qę�ͳ��um�Z#��q��nh�O\G�q��ͬ�0�q1-8�v�w��\��2]�O�A9�]�f��{Mgn�K�K{�x�r'�Ն��ҟbm�\���ʜ!�^@��v;u�i>YLEgck Y�U˦�����I�{�J�*r����a�Q��m�wu..���(���0!�e�Jg��Z3$�<�6�oT�!P��f_4��AR��2��r����CIY��#.�Y1��77�Utno��PAv���q�J��G� N����	�&�u���O�J�T$V�����dt�s����u�D����#L�JP�w\��g-��yV��aDZ�An.�W�]r�I��2�i�˗�����Dg5w��wv�hI$���ʍH�r"�u��Z�e���s"�C��a�"�!\�]#̢,���1ʔ�BV)EYFd����$)͝Đ\�u��]�vwS�+�t�=͸Qz&��(����	Ñz"�$Th���:9��y��W)U
�-�f���w-D�5r�EEU��Zz�Q�n��4%�w29����J����8�#�'"�t��=Z�����H��
�n�Z���҈�P���Hr,��+�{�������<磓�H����s���4�U����)�B��S����E���F����C�\��1�SN�,�Ů��Jr�eS}z��wF�^��t����<f��&r��0�瓬���/� ������ݨ��W��5/IӚ���vڿuU�%z|;�\y�D����nk�����6I����V��jXѫ�����v���q��J�(�̸��=�����ϟ����{�_���ߟ�4��1����W�K�t�,^	�
��t\A�C�r6e��^��>>3D��Yx|���ѹO���]6{���z���Օ<nωJ�2�W��$�"u���Te^E�{��d�W���.����7#ޯx�T��OA^�������2��G)�U��R��gg��%:J���HK�o,C�>��ȍ�O���=�C�z������g3}f�s\=���*wu�C�I~3 50�(ϼVZ���-�D��~ӑ��9��Q��UH�c,��9v���Һmp����6N��@���& 7P ${cʬ4e�TJ���#�}9��*-�IaLlϰ��vs�fJ�ܺ�mӫfn�,���&@�끸�_���n5�C�J�s����*p�u��\`m�r,��}��'�"�w�!�Y�RCW������Ӟ��y>^+d��o�e#R�s��&2�^ ���'=+s9)X�c{8t�����v�:94[|������K��ʖ2·Z�s|����ڟ4�B6��W1&[���h�ٛI�P�A�oYܝ2�;�.��Pp^���4n��'Q��kqa��ͱ���b��������^W��G��ώA��%�x�d
���lϤ�&߄���f�����3�<���T����{f�5��n�x\{��Ǜ�����n4
�����-Go�U56ח(��ǲ����NE���C��G/u�dG�����P���i�E��)�U{�,�"UoN�*���K������+պgK��=��}��>O�h��P���NK<,�Z��K�2�g/���G'�\@��6�]>'�}�/���ǽPa�^��ogz��W'�J�F<��w���߫4�>�g���Γ��~:�S�t_ƕ~'xM\x��\���gQ>�=�{!�2�p��{����ڹ�:�'v��ʁ>E��3}����{S3��z��:�i�}�ց����}S��O��~�B�eO��R���M��=9x�+�gv�T���UL�9�}ƨx<��Y�_�=��,�]����Щ�7��nļ��5S��O+�#h�'��Jf���Q�#<\�F�w8���#����yMe`���v�|=���V����ڵ\�y��#=���|���I�k���u��B��ޖ�)Z�U/6��rQ�1n�Ȳ�k�U�N�aeJ��f>���#j���2 Hp���ӫP���� j���^ {jDU����p��z��Kד9H�	fM!�u�F^%R}��m���l�?��$�Ix?s�[K�Uu-����;qn��՗�-ՙ�6����"�+g�3�wN�<w�U������>�f�9Q��(nP�WO�,H��Z\��8��ne{��у�ﭣ�ޑ��=�������0��rY�P@�Q@��HU;mת���}��7�%~�s�
x;�}�C���0={Ho��������q^�\M�3%��D�=��f>'{ǝ̩��5�>�`��FF2��Ty���H�q	��ޔO�NMǽ��."}�Ȝ�N�W(��K�ʗ�z�C���#����.H�]^�t_��z�x��٨ۆ�������� 7֥9.�nz�fO�z75���u�қ�����*pTK��R_�Q�R��/uǲ=�wG+��)(����ۭ���4sT���j��O�d�ЦSPrX�����+�>G����-�۟�����XS��Y[�3ϝ�1�>�W�߶\	���l�i�7|J��_�kC��8.U�Η�
>��CcP������ԇ�;n�xd'^Y�Azs�4'o�j�ƔN��f��d��u� �'_�N,3/%�VL Nyn�c��p�ľ䦬�]��6Vڕs�������eM�Swص_�{��*�Mn:y] �7RC�@�}kE�����RD� .��V����gY�,�s�s��Ȭn�����&@����"f�[��3���w�+i�N��W�}��~����O�ҜyՄ�{%��#&yB�M��˖2n'i�^�=$�x�v�Û��$��4� V&���W���v=uԿ9��z2�r�cdeP���w=���G�Ӓz���Js/A��W�n:���93��4��M�r�}��{��9�����P�Tt�����Ոw꨹T����kx�%�P�&|OP���)��"\�sAf��.Y�_Q���u^�Q���{��}�N�����+�q}$�2����,IR��],����&��h�mDת\�-*�;�^z=LnG��=q�;�s3�1�.K4�P,�l�N���B���hR�Q�d�A�֧/�P}t�p�r߯F|���V�z�����������'�f��=6v��n2"Rɫ۪��[�| ^��d	8�pO�VB�h���q7�,C �+����p�o�ꑦ⃮K��9ٽ��'ם��d�j %4H<�p7�/���h�kF���O�����>�ԧ�&;qG��ɜ���=�ں��U�4�%��RZ����1/ԅ\T�:7 t�֍F���[��؇�1Q��c�,V�zf�r�7��ns��ب�o*Ɖ����8ޞ�����]��q�]:�~��d{ծ���,G��G*�(�b��8ȧ
�8+���y:�Sר��\��َ]�5�l��lzV���>�Q�ݫ�͒ܥ�o+�iCo��L�1����c��	yQ���K8};�}�3XD9�HT\���^�������Zi��B�Qӭt��+֯�Z:�d/C���h����3Q�]>�$�,��0�D�/\ӆly8
%�ܕ;��F}�ԥ���ގWz<1�]�{��D?O�����(W�����=�I]XY5�Y���1�o��0��[��\�>[	_����������{�Vt��aįo��PվK/���R���$k���@�(=�.,�zU{����^sfh^�>�c�
����q�D�r��q�$��KN�xG��;� r~��������	��/(�=�U������W��7������o�߉ÛIxc��t��t]�?r솰�?L��Ȟ�{��J-��*�T/R�`�;��c�qݞ��1jʞ4<J]X�x���q�:�������� =H�6�^}�h7�i���=,b�z��R��9�F.!��f��{B�q/Ya̥k�������$�3�(K���'�޽���;��z���[H;a�Y�_��=� >.�ʃ6&�����,'v�;{��H�Y6e�A��X�Ѧ�t
]��f�A^��=쳭�=�Y�L�Y_g�R�%�Nv1+-���c#�ٙ�t�P�B+;c`,o1������fkơ�O�>�|���;�d���fC��C��n�s�şi�J��0�IJ��l�UP|z)����n��!zG��G��|J��u7�}����͋�������=��.�r �$0,7P+�R=~Ua��S򸛟z�>��$��m��8L�9W�s�Z{�8w�}r6�V��9�Y�qU�L���p7 �2h�>!:;a?wf	�Q�������3���p};�߽���W��Ie|�Hj�u2W�Ь���P<O�QB���r���a�o��ۈM_�}�g�x�%����_�%��<��5�?b�}�nk��v�Cۆ=�J��y5���_7r</�y]и�u�}�3�;�T`���~k��t ~?��_���e�6��G)���ݨz{���3�ut^�@t���q��o}��݌]���HϨ-YR
(��@8�������7�V���u)|o���b~�D�-��K��d�۞j��G��t�v7�ad��O�F�9>
�·qY^�_����磻6�R�F��Y����o��5�c�Wx�*��_�^�fp�>;;q3��4�{9GE~�r|�w��Тq�M6ş�%�5�u����$�-�i�ބ�Y\ڹ���x�|�N;R�{��n$�~4�!5*^Ρw�$.�A�V�ƶ�Y�6f�G
�-����S;��F�����6�r_qKtY���hA��J��q�v�Yr��-��H=��s�C�i͝��1z�|��Ʋ<2S�@ȉu��7V7�֣
#o*t�,����<��I�꧋b�K��J�J�CՓ\n:��^�;@�>~��u��z��?m!q�*x͵8��Z��F:�9M��I7@³�.���R7����T<F�zȿ������^Y�����GΧ׾��˝�R���Ow��=�E�x��r ʨr�خ� �q���������}#���ˍ1���f���1�ڙ�,o�m���]9�I�Xʡ�L�1u�J7IU�N�x�]��ql__��^�|Ԅ_��%��j�}�9�� �,� r�,	�)@�>nP@��L��}�JvA�q�J������'޴4g���h��ë�o�'o���0��e@��d(��z䍵S������H�8��,+�~�8y����c�����o�'M�W���,��a�%	�U�]�o���_�N��F�(�/r�n�Z�-?;`{҉󏇧&���h��g�$8r|+��ͻr���D�6e��26zH/��r��q�p�y�1��z����R��=
�\j���1�nr�;�;��v۱˂�@,�:�%Wm�k=G��򡹤uCST��m�{��D���%6�3��>Q,�\�],�v(���1,��V����h�9+�DI45�+��飄4��&�������.����c��[���TQD���5�S��5���3/�#c%�h����oT�7��q��}��fv��^�R+�|ͯuv�Dѿ{�{>f�m��fM)�T�,v�NIZplE=�
��'������y����ܯnB��чމ��z�޽�q��g��0Ս�o�\ו��ۢ�x��g�OGZ�Ogux;���G�'^Y�#�>�"sю�XUs6s�(��+�x��(��=�Q�B�����-�f:�)q�5��w5[ V��9�V�н^^��yՄ�G{i����kMt=�iew�o�K'tvCSU�ZnK�+#M0&��>��'���P�]�Dπ'�8��ߓ����'���,���z��1�@̮U��8*�������}���������5��{.=b�+������ˏx�R��^�A꜓����$�(~vL�,'�U�ώ~s���T���w!�
�^����F����=����[��36�2��7}$��,	�|�s����� ���^�9R���[ubn5��8w���8�uz���ǻ!�o�{�f��$��,ǲ<�*r�a�9U��
��AICj��ep�K�ӷ]�a�on�, ���-VS-s��N�讯@Os���þ��ܭM�ݒ�WQTP��8�WF:c0r��v�R�.VjK���+�eUΔ4�9]';2���=���M��Ïb�
�O3�,oK��<��4H�<��Z�����%�^�^��+~�P���Bt�{���q���T+����⏣���t��\M�+�fPѸ��q7>��0�+���W%)90����J�G�n(�n�}!�)��M�d�iSD�c�����h�֍GZ~���ꖣ�D�aج��Sϴ�A��^�~��d�_J��DĿR%���:_��F�dh�
W��3�T��?B�j����O�����5�S�d��r���/XU���=�C׋MN��/f�.{�e�{U讀�s���ީ��U���4n��;��5�O��(2{`d��oT5vn�	ϓ��G��X=���ݖ7UV�U=�So��'�{"�w��Y���p+�����4�C�N�zau�����V�s�>[�W�����2��9�CƮ=�a�I��d��,#�&�Xf���ߛ����-��2 �8=�gv��ey�R��:��q�j�1�W���|a�����M4R����>|��U��-W�d5�5P��m��<�6jW�G>ٗ��Wn{oju���&q$k+��:��K��-\F���n�X��@s����n�b~;�bo���n��u�fRŉ�L��*��lN'��U䐣s[ݏ��3���ª��YfGC�>�b�cy����Ђ�;�q'��VNż�(�jn�N���<Q̲�I\��'�%���?�G��9b��:*�tl/Iӷ,e	�
��Q�:�zfm5�v4�u�7���e���e����G*L�q�6{���z��[�	�w*���r�޵�'��AS<��z���L�.��Z�3C�G����=Ln{����C�>�5�ŵ�,�8{�X��f���C�I�����RS)���[ybGz�g��3��!���[��&��b��\O��/yu�67��騆x���z �yFX��P|z)����n��!zG��vM��[5>�c�9�&kw<�<E#�z�m��߇� %Ӑ)�,	�
�R=�4*����ʹFp'����W�IZ���ӜWx�:���u�e�:��*�dCs���P�m�4�7.c���K=KTc>�5HvO�m��>ζ���ӺM�޸���]�ȸs%��U$5$:����IVG�WI����O���Ƶr55^8��+>8}8�y��F@����\K�T}�1��=�&�����br��ѐ�MgL7�\�-��ҦK�fXq
� ��}G�������1���0��1��!��6��0���!��6��0������6��1���`1���1���6�������cm����co��6��1����6��0������6����6��1AY&SY���w'�Y�`P��3'� bE��碊���H���R
���
��������ZT�T�$��@�J@Mh%$��H )�$*���"!T�4��f�Z��b��Y�Q�	HZɣSc*�+5����5�mVfʖ�Lkm��ld�����f�Y�vr�m�f֭��ͭkm�ki�E�j��oY]5�[F5��)F��D�Y�f�m��ٰ�*V�l��d�Kl��-jڕ�kSi��SP`l��Mem����̙m�֍��+Z��s7n�Cmλ[[|   ������u����lӡ����W�^�����z��5=��u��W=U�ݽ=64훽j�M������mIS{������nw�۔�t�k���)[]rl�����e��   \���n��cާo^`��n�5�R�t{���[�@P��^=QEQE=�z(��(
(��K�EQEQG�z^�$QEQ@|=wF�P�g�x�PB�s��wf���֕B*�S33+   O�W]�V���o]��B�{{/�7���y{���ǭn����J��^k���l���{˶��=����]���Į��v���^U/Y�g��΅H�`lf�T�m�  �|]�����W�x��R�EӵZ�罷w��a��n���v���n׹�hV��q��w��UI��^������m��k�o+�wc��n�����h��m�UfmV�����km���|  woU���ݺ����޳�ݽ{����m�����{�u�F���z�����퇕�jSg�wc������5A^�{{�=z]�pz�{�^�ۤ�v�o[m)U�֊����^v�Wj(��]_  ����]����o<�<�g]ٻ�w��S�W[֬�z�zz�]��{l������5�{+�{Nn�um��z���m���ooow��X:-5�vOG�v�3{�t����ʖ�����fٶm��>  ۯ�J:}:]�^�v�=�=봻��]�n�����a;�o)[^f�q�Wy���w�]ۯu�=���g[�ޞ����Q�W�����{�t����K���ν��6֙�� ً5�R�e[o� s�F�}��]�=�J�K:�w�i틽��K%X��������-�����ފ�u���n����Ȫ]�ޮ�՞�۽����ޯo]w���og��4�n��"�h��)�wJ�HYm��j�  ޏl5�MJ�{v����i;��3�{���������E S����{
w]�����ڨ�
v����k֫�;v���
�Ylom�<�z%N���mu���[{���{k��5"Ͷ�ZSml��mmK�  ����+�����.Z:�[^�ݞ���W����]v����=K�<]��ש��������ס]��i��+�{n嚂�y��=*�������K�r�WO/womi�]�)�4��J��� ��a%)Q�  ��i��T�b  ���T�  ��RUA���ha&������h5?g������0~cv�5����^�����/Du�ś����[��k����䄐�$��BH@�a$ ؄��$��	!I��$�	"I�������s�ܿ��*����_�RX����o�U���ݗ�1��ռ/@{�T#V��1��D��a���z����'�ERDf�K#6H�q�V�ֱGR�e��R�m(�Pbd��V�X�X��͂�+Yu�N��o�:�cE�P�)l��w%6�?%� �d�̠n�߰;�e;P�T��v�6*ItD�5X0V�ݜ(�`Zl,t��	
��2T�v��t�d��9Kh
�t1o��P�E�2�Aڹ)�kS�{��WI�v��f݌�%�(�K�Z�e���Y�̗z�?)F�̭͈MZ#˷��)�0+�f H��o.��r�
�q°2�;�G�����ڌ,��D3lc��lQG6V�.<��k�� ��=d�Y��������V�bU��)����Ù�剛��,	Ko/SX��n��E`��q՝{2�6��"Y��k$pnc#3.L�����;��ߤۘ%
�8�v!�C��׵G\���Nި���NEI0Aʲ�SF�Z�I1�ӻq���MB�'��۴��.�Be�GK˰�vF��2e�v��ق4e���>&
Մ��� 3GN�I�BA1��*�32c��*<%��uv��im^7%�2�!'\��w5�$$��@@C٣2��ԭDc��Xto2�#��"jͳm�.�vf�ݫR�R16@Mݴ��)W�E���bb�K�m3�2��w�w.Dd�v����ǈ&]�ee�pH�ˣ�yy.�7*ܲĀ]+��!՗�6E��.�8%m������tpU��j�&̛J$ܛ�+L�uz����娗P����.�1�����٦���� ���6�G2���uop[��ɗ4-O���$�^�9%�qP9��4������㳇v6/r'X�B�T��\�/i^S�H��[�r��SJ��m]:��H���F`�*�
76M%��3i��f�p7M��5,����N�Mn�l&N���%�n�)*7>ƚ�H�t#B�ȳ0���֛�Y�
�@=��n��\V�?��&THSoEBj �-B���x�;E9�(ݬXᒤYv��,�Uc]�ykM6��٘��R�ט�4(e�t���c E-8�3���C0P�q 7+%䖷�C�+t�\�1SCFݖĭ�J��[c]޹�/Z�B17��q�;0!inj�{�d{5����IBM�t��ݕ�a��a�r��Bɸ+q#`�S`m�M�f���.X��I���r)�R��M*l��Vױ�zL�c�\��Uq/V�aF:�Pi��
��:�if8�P�$.#�2��kmJyJM5�)�j���nЭ�1P�Bڬ�ح��\z�5N��
�J|� ��h�{0�9H�A^�S�[���Z4�]=��KNe�w#��-6l��kUa,ei.���X�3.GfFP����X�m��5��lV-d��uoZ�pł˰��(+1�2ĺZT��Dcz.�uw��h��U�k_d� ��-�,�f�t��Fn��eTzq\��e���M��@��%4�<ߤ� bn����d��<â���<�Н��Y�.�i�<Lܐ�Y�`����a�
5��7XзBpiGSY���g3+ ���,6����l^�X�`Rf7�Mh��ꬫ�aV�`]��p�f��
��)ǘ��3)�C�JTj��܇j��u�#�2S2�UҬ����e;���m�#`�%^K&�����w���)a۳'�(�Vԡ�n�Z\�P��^6nv��Nm+
�Ыǀh�JW[aj�y6��'M;Z+f�����[ǥ���bKf�`�WDK���,CE] #��9Rʸ�^�.���LV�	Ku�Y"�X�,+ ��j�Ũ]�:ܵ��*8ڗY5b��T4�5m�*�-��aX������r<�v�����]ёܫޜ`P�J�mE�Z�!o/e�Sl��ɢ��B�U��M �f��D���ҽ���0d@�1���S�G^����14�r�[�Pp�7i�fi�1�v�LQ�����0����N1�i�N�/Sj���[MX�YB�¦��
���-d� �tCV�drt�y��u�l�.н�L6�*X���LZ�5�
���Qwq��7TL6]�z��Jʘ�u�VkMcm%�@��,��k�Q��X��oUQ�d��
�S�s��4�Ax��e��a��B��q�>��ދ	J+t�b����iT7+��90̑�*�Mb4��n;V�e`F�g��02
`���t� �ݚݧ�R��ĦU<n�ي�i��6���U��yae�$gJ����ԛKJ�%-��a�B�Y��BKu�Mcj1gY��6&D&��r����N��ccV����Yg�՚�U���W��D��Sf�s��sMCy�� m�"��D�R�L{uT6D���V��j����V��Pس��>��Gz��IM��t��
Z%-�D�]ᰎfj��e*����,�7IV����K��1A)ZQ���j�Zf�N��n'K*��e+W���|/�gs)ʹ3�k�����2�e;Dk^CZb��vP���誺�6�ģHh�q��aA�ԗN���BXp䱃iL�No����-��:��L�
�z�2�A���H�ɡ!N7���
u�xo.n6t��p]�y�00@�M�B��Y��F�j̰�����๋�D�M`v!�vi�x��<�0ɩ���Ǚ ��u�8�4���E�ڱF����֌pc���R��Kc�ƪ�`Q�{�Q�a�X�7v�9Y�3&�����Z�����o7J$+^�{\�,c��.K-�P^ݍ���:���da�4c�*�k3I�X�E�[nly(1�����PJ�5��͛��ڳJɦ*lml�	��]�R �V9�4��N�1nVf-z��hY{��yy�5�� MRTT�t�X���#��"�C:&Gu�kF�!P�R��Df��u)�����eZZ6��u���)�j�n��8*V��sfV�zV|LQ<j,�H�\�/
�P���b��5����)��p�E�Ѯ�Lf��)�At�Nm*n�f0�3f�-Un���f��mY���2�S%�#vn��n�ɍ�YǑ����i���Z�0lU�lGY�|R���[N�56�+�y�J��Fl����M��-"�[VL��LMi�᫺�Ei X� kZ�jr�#T���*�G-�e���Tf=T0��Y۵ojbu����R�c��me��%���s��]��Ds$��̑52�ML�+5����Te��&�sp��U,u
s�����*i]�S�l$�r[�'okRo	��9�T҃c�U����'ҷn�-�e��
8�X1��m���$�ٻ�Τ�Ӱ�G:����z�gX�8���qڒ�I����䨋@#j����E�l8К��NV�y@ܠ7@Q6�[����&�aTt6�@%��J�ڽ��Z��Y������M�x�jSHj�Ux�X�m�t��-U���:n�㎅ �q]����I+xp�-g�^S��%!u#,�Www�F)�6���lT��ݙX�oT����)��Vi-ѼT�͚i�A�%*a4ӥ�@�Oidv�:h�N��w�t�v��z�vsU�K#QjA8j���j1�em��Dh�nG*�*[4�����9V�Q5j���p=b��%����9��1JX	���]��[�*U�f�2�a�ow�!єTEꤱ����0]f�����ĳkn1� G�� ��nD���u�+�R�)	��[����(c.�;�)�VM;MR��l�Fj�l2�d9����ں��E��d;ĥ��p�*mZB��*�Nڶ���w.��ol-)�5R�X���-#����Pj��]M�7	B�H� ����;�Z��+�����Zs"q�l��U%��L���r��J�\M�eMkM��s"-�1V�Ct(�����3��ݴ��U�%�Pa�Ӡ�i;RI�Z�f�Lˬ�-L���5d��e�*�(�i�8Tǉl9���j��@`7��6 �� �.�Ƒ.H�&̈R8(�ڷB�q�y#������
͓�s ��3��1��G��cA-�q*{t�[7j��ZP ��q�mZ�ɌA��u�5�w
m1�@me�����V�q�r^X��i�~ʼ�ͼIMRЊD&h%���I���F�\fi�w��U�Sj̶�z0��R]��a�kB�(�q*tU&�G0�V桒�Am��MGQU�.�PZ�)�	fާ��r��̸��e�N_͵����kN�и�0����2��o)����1TGn��Ʊ�T֬� �CF���IH��΂6�*�u�:Ua��sR�Xw��G!Su"�3i��Z"g��7�=��}�/1�z��Nd`�ddlɔ���YH����Bl5�V��h9yI�:��.����D)�i�,�p�K�܏Rg�7$Y��,�s���ZŬv����e=h]�x2�F-k*�0�^JU�`V�WK6�YxvVk�ƑW��(�2(�y�������̻k`^T$�AR������2U�(�*Mn��N���qA��Z��B��4� ]`a1��w����ʴю�ڵ�i��dC&ax��v�+cu2ʁ�,"�r�"���T�������t��jޡ!�
�/讶���D_ג� �j)hc�Ǚ"
���KKD7�IQ�L1%]�J)tk3E����ҫ���m\�U��	��`4��G3%�21P�v`�������6�^�e�&�F#ϛǆ�����J"�ċ[�n��݈��q�ʊa���{6��ϢvY{B�-h (R�LHf�wR���X���R�[tM�.�iԤtJ4����6�����dT�g^tAvαW�&�d�;�,��H#2]�5��RTCa��Jy@-�y�]�/�K���Z;!*j;S,@RΗ���xV�wY��j���Q�&�7�=�w�v�lwJʎ�7��atb9��'!H<(Z�#K�q���6�Lnh��3Pf-�/&x�cnjb^��۵f��H�}.��Z�N��rf7�O�٪%ɺ&�%Bvˤ���L�YBY#hŦ�*�/r�@ ������Q�k-e�0�q�0j�Y�U�od	�,��qV���0:�a����c%d�yO^��c�2�.ۂ�(̂�H���sH��r���]#S���a;�,���ѐ�+����Ou.�C�O7�4t����!���ϒg[TV4�b��m���1�W�L�i��������f�
��qZ�����
j�5P�q�u����-IMꛚ�Q�dj���&j�"�m�(9Xt��[G+�r��N*'&m/��"Ҡ���k�B�vQpO[�Ж�VV�V�p:�lm�2܆]������6S&Fe�Y��൉�j|sv���Ӽ@bi�ˆ����TʹRU����~ZRI)��R��h��Cnٔ��/nd�����G]m4�1��t�r���+Y*�k���Km#�r�;�EGd��6<���ɮ�bD,�j�nX
�Xs>�&�BK��*Ԗ��[��ʽI�	%�Ve�e�����;6��2������j��.��I7Iũr옢���%�4P7H��V� V��x�ݢcJ�5Q����F�e-4��c�ඝc$�dWoZA]Ih�����|�Ø�̻���̧&n<T�A�I�[fm�$Ӣ�� 
�������	��Q�Aw���q(RGI���Ѕ���us�P��f�b�.�j�C7��E��
%���3e���.)�T� p^��V�D�Y�.�ۻ����ˉZ��ՍV���n���A"vQ�&aڵX�ں��u7'�Oؚ��^EhLF�l!�<����.��8H��݂ZƵ���h_iWp�P�w�le����F��nVu,�[L�ܸN@܊,̊��s]�XDX���a�6#ȩ	������	�
,��MGmޝ�4A�:��	��	�F�j�kN�0�QXj���$�Rm��&�i֕�q��k/	ӥn���s-3K6��܉;�&V�r͠�Q��^G*�;�_L�S@8+q$�iۼ��*���޲2!@"w
R�Y��������`ͤ�X����V
pm����K��˻��L3��0��Ĭ��e,Ƶ'lE��L�	�6�l:Yh$[IX��Y�HZ���Pv�f�ѯj�U6聏e˥��D�ViÛ �t�jbԮ��4e���yO^ѫ6��k�I��z��1Է#+S$�Zj��݉P�-��U�`W�@tT��W+Sͺ�X٣d0�[i@��d�H�P���V�kJ�e&���%/U킎T�.V$�����Q܀�X-;Z��яX�`��j�t�K ��c*���{hrͥ�����N��M�wB�+��b1���j���R�7�V@T�He��aG��0V�U��+�P;V�:e�VY�%,��%3V�,?�t��M�Hl��aޑW`m1X��L�z�.V�̂ҋZ�h�k �q��(ձ�՛��B+� �kP� �׮һn�f��@�K&Izl�Rd]�W��7w>�Z�$���jʎ8�q'X���G*(libY7cû��$j"�B»	�q,VZ�ۅ}wAaC'F��U8nK&�k�B��5�����0ӣ�w	��F��6���+�Ov�&�gp�T��͹5�c�$��eX)�l���lN�ݩ{'�S��8ӵbQia�n�R�R�r�V�z{�o���K�F���_m�Þ֣�!킌釥Y�pE{�.L�3�b�����9gC�]2u]E�����hx�ǻ��;LH��׵�e!;/�!��
�d'L��I\�a�1t�8;Gl��_i�9Y5H	�:��ۻp��4g�`JeARŹ��Y:�����Ɔ[ꨵ�rH��/�Ѩ"ˁ��r���v'|��"��P�Z��T�Rj����a��s;+:���U.y��6&A��%����,u�G�T�5Uq!�i�E;�N�T-��{۵���G��裲��Ca�mt�
�Y���㳖���a�W�G)��
wّ��n$�!�]�/Hxf
ʥ ��ikT7K��a�s��*����{�/C��n��l){�g �oN͢.tF�u�ڙR���RK{ǁS�nβ7':8�աܰsQ]j�;*��K��lu-Ո.#�]úg0Ǳ���:6��²�'�@�u��
��_<�ڟd��:��z fit��̳�e1q�C*1S�l���5�'V���QVf]�s��B�9��"�̾�.ǃu]�Ҳt-&u�R����8!�{�Ծ�!QC[]��C�<�K�D-N৪gF!�@�zP<F���a��b�9+E�í�-h<�UzL��N�T9z���je3�nV��"i���Ze�ڳ\�z�u:��cM�Km������*-\�bonb�Ժ�e�i�Jx�_e$�`�4V�����S�=��r��z�s��o�)-��$��{o�)՚�&����td NթlZ8G�4���:6�^tĪw{Ά5S	��
J����c��S�)�0+uӰ�֛�ƞ<�
e��$�Fnq}�ƙ���v�O��6�po��t���6n*l��t��r ��YW9ku���LrLR��Y\Q�A�ۚ�^�)o-k�d��)�oFU��o+%�o�?�~�p�����T^Z��Q��9YnM�)���c$ᜫJ��s�;��H�����e�œ3/�2�x/r�$����ڡG�Y�P0�����9��F�M��O`�6`�D=v��Z�Y�1Du\s�n����-��.-1���֍���b���w���!˝9�a�ObҺ��eP��Z�qW7m��/F!�qn��me�.��m��g)Mڝx��C�'=��\�nJ+c�`�c���08.8�U7���ۻ�4>N�m�z&V:�*��9��-�+N�Ap�El��mV�n�nsv�)ܹG�x�`͏�X����^����1��4��z�-�pͫ٪M�2���G�˱��
�5� 9�=�����&�Z�:E�Y;��\4����y�%��ͨ��!7xw��/��jsop�H�$��静i�kr���T� �|]A�NG��99#�sNj�f�9kN+0�����-��g,>��	}���K9�W(�o]ˍ晡�(T��16ً����3�n�Z1���U�:�R����"�ﶦ�qd>xhmWfh��Z2��/���JO	*�xIz��ǽJf8���X����[aܒ���sf�;�;gP#�v�_��};������>��F��M��FnZ�:P��̙�؊��<I�/r�]��wu)�d|	H:yw�}�����׊.h��	������1˔�Wբ�����7��v�Z����1K:ʲ�TGu+�!k;��?i�T��;����bJ����Ρ�'eZ�9ՙ[�Uд͂�ܠ�(A֗����]�vXu��m�L���V��:�J�t��*�S7�ڕp�Վ�dJޝ��1hNo49>���Au-�m�㦕m�R��Ёdv	+��׎آ��B�m�7K�'��`��H���� .���̴�pAu��]��݊C�f����#l����H�#��`�}%-�#�L�&;�LQ6�r�y��78�̮Yt���dLҸb	q���z�sgw/��T"��dX]�ݵ(6��]�ށ���rw4�X��s"�9{/O�#R�A۩N
S9{bEFž�ǷX�FuQ�Qh�s�WW�T�bu���zT�@R�ѻ�1srn�6�)��t��
[�����=�*}� �C�7��e����aZт�ɵ"�i�aV�wq:{�ދ�{r+=�:�{��A]iG�G�{����Y�<�d�:�w�˂�-f#�gKΪ5�jP�'gk)9/8������(=�~ʅ��z(���i|ݠ2�eAj��dKY�,�II��ݶʂj�ƌ��Kk���m�[d>�����rF����R�e]zp�� S间�6�R�����w���Z!p`�9�(��aP�3�6�X��q��>�U��Z�UnR�*rYԵ�PK�sB'�hL���:u�mvC�^���L�Ɨ/�q��Ql�Xk�^~9�A����pY��Ok���ͫ��V5t���O����.�O$^u��]�"��|Q�}�)��tTu:>t�\�s�^�Ox�p��4�vf��@Z�Ђά�WҎMHt��r��{�s	ck��\q|(V�����������|��������(�O$������m����m�f�}��KdI�/`���Z��|�(z��� ��pX�V���@���:!�kI�&�u����1fˡٳ�O����e��a�I16�'C���ȸ?�κV�é��Yq���k�{���	\�)a�NewJ�/���X�Iɜ�zi�`���ݼ�f��z񳐲/K+�!ϴuN��3處��X�v��]����u�y����BI4v���+d�Մ&��55َmw�b��r�՞�s(J�F�H_�NX#��1��>�5�U�f뱌�61���6�Vvv�c����0�iG�$���4��-T�%�88�vFv��ϙ��}�8��"�@Ҽ��wj� ���Í,^Ǎ�j{2�͋H�p���or+T���s��6�K����x%N�,;oQ�}FJ(�]�5[V�eMY�]h)D��e�{f͹կ�/fu��E
�}F�m�Xh`Ң&���q��9A�+����`Y��GF���W[\���9�XD���x`��,�kdl=���=;�R��6��Bc��,f̩����K�o.��%�W9ꢐ���p�W��1jg`��먬�u�N��5[�t��H,rWAM
�38^K��C��Eg�h�R�'W6�z��c�Jvfm25t�9'k|�hv��`쩲0�����������F]��9��+���BF������1W^]G.A��rH�^��&gT�3EV{��orK뒍����e�1�f�Jϰ�ó�[��rV��K��S�j�}��#���(SsB�,�ڬns�3��g ��9���X4+�}Qۚ땱�(�,.@�T;�nV�}��%�i�"�w�����5rn���g\GU-��U�3$����!�!�'�8.ڝW�r��U}Z�gk�Dw�
>�.q2:��u�9I
��o8�s���72�R��m�E��kf��a�����m�@�}���§d�x,�h�O���;`8�w�c?b��;D��FB�Ӊ�K�G{��3�œL�k9*�"�1�9�a���fs˒�M�'�����uifp�+
�c�`qυt��j��a�	lU�aZ|V�:ʝ��4d���-�Z�"HB�ʂ������em��!�C*�ͽ�A4����OyN��NCʮfy�N�:jY��kΗT)]�87SZ��K������Y��v�v���BZαJktA��ܱ��5w�v�j>�x^��/�ehR讗��b���qr��.�i����肋SG%����$;�Tg7o �p��;��[W�d[�vņph2�ę�@wչ�n��l����&-��3I܈%WZq;±s�[B��n�m�ŝ�Lu�G2�
{8lۮ�K�Ǎ�A�j�����6�j��
�f��~����L��t������=�:�d�{�ă���2�x'���Z�7;4v�P��8V�}
��w��oˌ)�q�<�4!ԕ��Y��~ڈW�4�ȱ&���-X�9]�I]1PIԟ��Zi��,}�p�ʉ�Ň�d>�_-sb��$�W�\b��������D�ά�:ɩ$���$�\����E�`�����.�!�V��W1��-��8D�:��a��y(']y�M��F�(��fj�ov`�2�B����x�pP��ly����t�m��KE-����o
�}D.t�U8Vh6���b�Ch��6�X�8�vDB���=R'Me�8OFg�����8���ƭ8,�:�4tb]��gs�u�J�Up|�b�rBe[���ê�N�l�H) �6mH��;J��[����c�9"�M7�7XLV�ts_q�/U=����.�1�O�d�42l���C9ɓq΃�l�nYc�7�U�.Ԯw	ٔ;��}�{D�K�b�'@����N�t�a�!њ�T��֦�L`���I�u��#�g5'Z��+q}���t��~Ci���WgB2�tu���v��G]h��{@
7tǉ�SBgNy��"D4O`��8��� 2_n]��ye⫛ñ�5a�Р�{��`��l�S��8���,hF���\�µ���qV�^��X��<upv��s�%=��un�.A+�S,��o[��_v�Gz�k�4�e��^�pN����JaoFaW��9��E�qLd�j�A\�ޟ]��O`�Gn�qi�8C�QCsJ���\��N��׼��ETO
x�8�8�!�j�� �)���ُ�崁��U?��ĥ̝�[���z�>1�`iuREg���WX��ِ��.�_
�Ϭ!q�|o:U��v�K��6��c�VK(p9x�pA c����m`m��8:����&t��ٹɳW4n��y4�G���7a��������"
�Tn�ٕwK�t��ruJr�|�F����wOl9�dm��������O�
�����h���k�S���\hi�{ ؅�`��Om��Gt�Լ�y 5�n��Jx�ngf*Z��f  �6��&e�>��;o6p��ʚ+7����W��BmV��vL��/v�̀�#��1� N,��}Õ܂�&�����*��H�E�o|���O��D�ޝ�;��M�<�Lɥ�k�vbiq���t*_%C�|`DL�rU�N#��M�L���ܻ�(�o�N��ՆuL�K��TQ��[�Qu{��Ǥ�A�ؘ�W�l�%�.�+!nm)����1�y ߵnv_5a�-�����ٵè�7˕a٘�>��M��K�9Hlb{ΐz�-z��`�v�7U���l��t������DH'
��3�������&�6R�٪ޠ�n�6�U�o��yVr� ����K��8ʬ4<�	��PD�J/v������=:��g��5�r'ƺٌ���њ�p���7�#:]p�LƱL���KgE(�{��ޅ��R�D��2��3l�^��M�i�r�=�#<:ć�+Su�b��'x/&x�v�TzS�9;�4Q9t�UBm�$
V�z�Vm;t�:��0j��9�^}�\�wp��l;�&�)ccj_Yf`���K87�p/l�K1�,V1���ǲQuJ9|��|X�Q^�2u�tgal����Z�Y��in��4p���n[�� �6�2:�N�3��*J�T!lĺ`o;��8�w�`�%�֫���n��r��5,��
��[Vsd1����aM�Y�[K��v�l����c��siuM�	ǳ�T�1�:���;�[{0��̄O^��+D���¯fbP�-F&�gMh�����i*�<:NG}��|w��w*y�aϟ-��rk��rLٴ!�����L��r�2�t�1 ]�MAu�fX�e�շN3ƹ�ԇ%��k8�ٖ!��wv�R�:Q��Q5������33��մ��y�=�v�@�4�@s ,ݺ�W�]����]
�ru���zH���D���y���h}��>��ɔ۵��]��N�)ާ�f"Ұ���-ʹ-��u���4���:�Ci`��n�I�f;���Z���M�0���_�8��8�U^9]1Z�v9�k�V��$���Y7��`�Q���d���W(�N�t~�x�kQlV��X�
;�Д�B�K�������o�߈�U�su�n��!gK���y��6����k�b���f�g!�V_֩k;�T�[��� �潵i��2Ν�c��e�B-o��Q�-��w|eZ:nK��Q9�����I��hr�R�밁�L7*	˩��3I��s#م�((wt�`�B�G�wW]��*��.*�;�}�Qc�p���F�S��7��zP����HC>�7�<��a#
�vN�Z84�;��p֯3ӝY�I'�gR��<'0#ݽu�dч(�yvu���SZ;$S�s�H,��Ae��L���9�-�O�:���B�D���@�jU���WF ����8_nJ�v�\�P�Z#�%�M�6,�Qɣ�������)��t5(VR�ml�B�ֺ޸^����Y+o��=��9���и3�gN`�t@�q�1�ɜ�@(�$Z�-�R=�Y������j�v���5TC�|��f��۶�P��]���C���(��M�4���[�
/75����o��7�6Ufwme�ڄ�s��%�fuE���Y�Δ��Qʚ�]�@��\�VA�ff�2&O��@�s�N:�Adb�<	�N�+�������`ۗ�Y�q�_R�Cx�l�,K5@(c���V�0s���ֲ�Tr�����E:y�㋦�r�M��˙!�=7�<������QK�7-):��A�NJLWKL��@�Wv8���N��Yɭ͚�f�\�ދ� ��Kvk�r:�晊�v�j�e̚Qu"��fL]�+#ҳd�
�QUN\��������k����HH$$�	'��׿w�ׂ���V)��Z��.c������sН¤�gd�����Z!b7\z^ed����&�vJ��Qս�"���6�W�8*�<�e��e�gn�8p�l%���6�%X�qvX�M��P�vԍ�1դ'SJC�.���)و�R�[Y����Ս0
�n���Ɩ������0�W��
	���a�r��xpG�rDg
�ɮ���C�>�&Vf���T`+�M=7n&�=��ph�*��n�k4��{ُ�A�ƆS�of�N.#u���\�n�s"����v��P��M9M����,��x�a�{Z�v;Zn�Y�}�m.�n�e��i�Fh��j�����Q��\E!w���JYz�Xc*4�v:j�o6�x\�����īz��5<c]�t��5��9�V.5�I�[�Jsa&֌I�w�s��b���/;9�w5����P�$�
	�TJ'�C�����-�u1@��n0�c��R_G{�&&��WQ�}�[�Z��͉a�.w�IW�ڤ�7�M'��1Z��\�0�6�vVӌp��Sn�κxw`�lg�0qd���oRmT�;K���v;�z�SK�C����|:^*����H[˒{nP�ڔ���U�9�qֹМ�3�t�P숤��AR)x���V�˦kI/gQUdા��B�ܰ��U"� �Qc�ڕ(h!���<qGG�N�)y�_\$�q���T��[Wl����ׂ���4[V���Yt+�f���5�ׂ�e���X�T��'q���x2���v7(�S�9�]�F;YYp\Y����V�/�c �,>���E#mXV���q�n&��sV����z5�Χu�4H|�ô�:���ͣk�/�ǝ"�8`u�]��GW��:܋�n�5667�\د�#�廱���-�]����_P�o���q| �p�v�_T�W;����DЕ��ݾ�kB!ۉقi�t"�8��I���ݭ�xm�i]�W��n뵗��wK"��MN��l�v������N9�Fr_J��mR������r�v��Q�Cx�����o2���Sژԕ0�L�`�Ng!��!�/�\���́&�c�4���I�4�G��ʝ;:�3��*Gr�sj�Ӝ���j&O۳A�/�g+�}��֖|���U�ʕ2�*�p�vBFe��C��m��Qʎ�u<o�lƐ��`g�c4p��e�NZOBu}cKu��#��7��q|�D@O:�;B�ZvJ���2Ӛ:�i�T&�ˉ���*�5g�.��{h�7J�U0�K�EJs�*[���M���ʭ{���<�e��.�kS�/^k\�`���V��^�t��.<�jGnb�q�Ò���Ż:芜�%Kp�H�ɛ.���tޕ�x嵭n�yB�ifU�se���grZk�۴Z竒d�Ҋ&�eE���Qlh�i�]}���B�e�\{X�tXhiއ�(�:�e�H���1x�y�.\W6`��u׮4	��D5���o&=���A�*��u�3��%]q���VbL
�od��<�34q�cL�np7F��mg2Rx�I�0Mf+�w�o�8f%�B���M��g(j�<�n;od��S7���!��V�[*����\E������Im]��o7$�2��7� Uƃ�w���%�-F�r,�*Η�e�bV�VR�ky_5���X��I�J�NO�7���@�0�&�W;�H}�{iKa�5��B��gglF�}!�e��؝��%��p��3�@��4����:�p|u7e^n�\3 ��!N�%�v
�@��c�={�#�z�ʌ���b4��S<kvt�u6�$l�wȄ�c�,;����/�h\��γ�
sڬw.��ReM!t16�:��-̶��\���_. .�y�9oS��JS�tRV>t�/�@0Z�ZnN��EX��c5�S�z���Ӽ���G\��C�&�WZ��9|�ޣ�*	j�
(�}k3s���*�,��� ��=�E�-s[�y���/�h�S1>�W]� �l��X �B�+��:#���f��%;����aI��X�K��{[;�M�4� �v�,k��-�4��irF��\L�KT �:(mG���U+�������)-���)(��Wu�ݝ>u���U��e�ط/�Uq�ip��D�`qn����us�e���MfrI�eKgq���Gwt��\!��3cV����B��tJځ͵X�	��SĈOS�W]��Hɲn��m��̫�xQ4�Wu���]TB��n�Ahٕi��1x�2a�f�\����n�G�s��W�mS�ގ�A���[�a����Et��X��vCV���Z��0$h��w�uu��]q���MAt�v7Y�;��o�Sfh�]׊9�C#�1[��7��v���j
��t�q�%��DӘ���-{t�\�SQ˽�]N�-�{�jn��.��"a�\)��X�W�����HR�o�Gy͢m[�z숺�
�e���m�m�	/u�{�Pzz��/�cWι�#�Pw,�t{i�Z-�ɶ+r�̸ OE o2�朘�
��]'.���͒dK^nǷ ��V�iНs���ږ&�a��ZKk.j+jث�JP�DZ��[���>��2��#mv�&>�:M6j�s�Z�����B�mea�j�D8�r�v��Z-i�q�f�C�N�f����M
wh�V>�1�;�}����E šm�,�����*A�س����+(0�׷�X�֪������@u9Ƣ|)��S���:o��gV����V��Mjͮ%�N��e�("�bnʲ4c��.��b/&�2�9lT3�Y٨�_��6����ڋ���*P2�J�kA;&C�:*�Y��
�c[���B�d֪�u\�j��$۪�̷ֻ��oub�,!nT�i[��
�z���wS{��H��%76��E�>Q�����䡵���50b�T�@��C�xv���uY��J���K�sP̧��Y˫-
�ۢ�y�УN�ϻ��N�*2hR媗<�j
w*	�
��v����e�ϱpy�Pܦ��0�:�+�$#�"w�	8�XU3��):i[p��V$��b����}L�Ŕ�I"�]�{��ENL�܎쨕m��&4rn]�m:�7A �Ref�1�֔*m��Ur��}l=
��T!бe��V�
��8�iOVZ�/�b�b�p�ɝ6܊���tiE�Fν����c'W�f�>�x�Vp�/kD e��tT���V Ln���>5�Rl]�����ټd��v@tu��w����v:͏Bi��kx}0=�Y7�J�H��:��Inptw!V�2 |�D/�;���䷘ ��|H�I1+ͰWQ��p�7�G��n4	�h�I� ��m�Y���=�M�͔�ѻ��sZ+*�=���6.��٩삞�P��*|]q��70p��I��hz��fn]��v	�۹nR겥eb��2�q#tI�ڬ��z�P3Υ�YnȨ6�p��j��AĲ��h�F���H>̙r���(8+v j���8{m+��H��7��iV�e���e��-��P<�6vf6j�zp� ˑ�$�Rr��tZq��8*�K���%�+8���޵�������tܑ}-��ڙk����UR�լ�φWIx�׆a��z�P� T��Xq������ط��3iR.<�iP�v��ȺI�=�B��T�ǅ���[�:w�<&�R���F�r�b�|���t\^�㒻�&u���+��^v���5D(���ʴwN�J�Ʀ*
��C��9�u%�?��F��Z�Wst��`#���Φ�"��8�ݗ����ѹ"��`[�_Z=z��G����t/i�N�9��4tuv������d-V�֦]=5�rF��	7����7j���63�r�֮gB���"�p����l���5�V�]�z�n>\lؾZ�v�w��'V�r�VT�N��}������{7D�#M�?t���OQ��҅t�3l�'��5:]Y���e�3@��J��%`�_.t�.�l�ط�oH���v�.�0��k(k۽dVs7X�˔� 44�ۦ�i8�EM
]�V�.�䢚ukȧ�o1�0^�(5*�wi�nY;�1_E\f��$PM���E�.�MvT�)N��#-��;�vUhח ��]8��Ac�6�]��	Q��ղ�p�>�)Lj�r�09E9/�Fޥ���1eK�u�,Ɏ�h����N��8v�]���]���)�[���B�nG-��R�����'.X�Y�R�:V�������[�m��nj�̄�'UN��@^����}��+)�̹H,㝇2�V򮲙�DA��DV���W�:��y�Wϳ�]�6��\)�#a��-�J��`�,��8i���Uu}f��Ը��[ѧ�T��Q�"Κ @�+����nQ�k���ȧՊ�#8�ݗդ�Ɲ��l*z����X鬛��[�,դ�X��7�(���CO8�ܝ]ϳz�KX�8Lz��Ց�A%W�tP�S0�(�L:��u<^tʚ�M�!eN����v�����Rr���Qj�;�`!w:T:0�k�ԕ����ٳu1i
��^�l폩�9�x��V1uD�����@�L�\��A�бn'r�3������ԭ�&�hn�ǘ"ݑ�h㙔��H��7U�m���tk��׍"�,{´�+:����6zBܱx�C;Vz��fŃ���P��Ҍ�b�V=�م�ksQ�;;�[\-�&��C97K5^�� 6H��)�o(*�*q"���)���w!�ipH�n�V�A)��5�oy�g9�Pl��+�n���s����Vj.O&p�:굅xQ��	�76Pk7g,�n�f7�8����Z]O�o��\!���o�`�FǠ�=�ҭ,���؛�[����T˲�fuꐋ�<K�]���D�������U�4�m��m�Y��,W	�[�c5�U��r�"�44]�f��]ؓ�bG@�s�ԆN��Vs�:z���N;
`�6��8��0+!�]���nնin��qS��ɪX���=����ְ��tGn\�]G���3f�|���C7��3{F�؎�iP*�Kn����Anj��&����s#�5�0ms��>YaV���\��9�#��&�s���,���f�,��y���8���Q��QdlI>y&6K9L��m�q��.�[D�r�ҷ.VA��M��p(ʜg�����#}�%�2���[9W��0fܾ�6�;SoG{ѫ���-֣�崛�#��-���g*�;����Ԃl���m��%�;I\3^^&{�'x�Ċ��}X:�2�r[=��L���$���,-�E�T�B�	���.�%"�y��`{	�yR,:�M�:Y�o|�K��d�t7aќP��)��Վ�ybj�ތ����i�E9҄;;B�7�T,=�;������DZѮ��;'F3���Jcd4Ѓ�-8<��,�L�p��e室�#�]Y���Ғ웉����l_*Y ���@���Ń+u��:��ӋGMj�;Km*+�	p�|�׵��0��e�Oέ�7�Hu%��v��� ُvܛ3[���y�A#}q.�6�w���1�KT�x��������3H��i30VX�3�[��J!v;]���$_f!�����E�R�(-ӄr�٩ �%��b��U7pV���Tv3I�|���A�+�pА&y)Z1��)��v�*���coH�Ks)]B��J���R�\�Ym�|K�W�ggɚ�r��[�9M����^	��X�hT!lB�nd��U�����6B��1�]�f��rn��ts��@;;�4�_9՗�PCR�Y-sT>��Ƀ;���v.������.YON;�˔% �.���U6���	�o5�;yN̹J�q�M�ʫ��q�G�+���k5��ǯ��*AX�h�&r�P�LY����G*�*e�;����j�j�񴶆e˚�]Wf�Pb�*:m�OZ�F!VE�_>��('�%�<���l�>FV�wXl%�o_J[e[��tșh��U(o>��U���9���TF���[��]�L�w
�Yw}.�Q�T�|J���6��o��q[Z��i�s/�,�X,��Q�Ho$��vgJ��L��8�a�G���W�k1gjg����α(3:hf�]����Rs	
t�`r�,>���Nj��v����S���v`�.�\)�.B��#H;�r�>c�I��n�����dHZ��iJ�
��#�#x	���LN���Dۿ����(:�.ø��
s�7��	dڝ�9j#p�ט)���a�Ŏ���l������8rX)�� 2mѦo趲�n܈��|���8�%����֪Z1q1L��er�q&��ls�w8����9�ٗ���oDs������f�D
]�������m�7��n��WC�ڥ�ᬳv��p�1v;ӓ7�ɗK� �V!�cm����ˇ�zNr�}�Ay��9x8+.�]t��a��6�P�etʐS�����#[�����r����p���U����%�o0�/	��]n�-O����{��[Y�H�4	�7�Q쿷9Z��Qp!	��H���9N�Q�B����KW]ޞuܓ���F��Z:O�`lA2�7b����3�,̚�\���5Sm�q.U9m8!���/���.���7C/��ٔ1�(Z]�*��!#K�G����=�Py�h����Գ{���6�<�u��(ƭ����U�*��3|j��yG�vzt�BB�B "�0��3r���v5�u]�V�S]f��-]�b4�嗇��ɽ'`c��i��\��I�5ʳzD�%�:���q������9�0�b�������`��^vSօ䭶C}	�{�T�vm��7��Wfr��hmt�uv�O��Q��v�c�ycMt��ݲ�$�����A��D��AEr�uQ���:j���v���p
]�ɳ�i[n#Z�g;b�N-/x�� tgY!�Ñ��®�[�P�R��VC��b�j<�c���b3���n��M��!�.Xk���r�2���h��?������Z�]�GP�u��W(�v�h��u؇�#����F�;�um�-��g�����j�W�Dt�jEzu��֪^6��=x]�uo�Йf��貺�օ(��\rp�`���\��Q^;�<Y�,#s�u7F�]�����}�^/��<x�#[ǉQ�cf&�9�x����QF;���Z{�]\oy����Lr�Fٷ�xcI�,�����iN���H�:���� �U��kv��4����+��U�c���K(`dmXݻ�Ԝ�T�<Ӌ:�ǒ 8m�V���9���E���LJ�[}rc��Vb�P�oC��}��5��������}��3���R�-����k*e,U1�Q�TV*�21\k�U�R1�AA2����Ab�#R����c,PD\d��PT[il�B��l��1��D�U�Xc
�,PX))m�fZ�P(� ��,�Q-�4q�%�aib(�bT�VUVER�Z�LJ�F&YX�9eb���KiQPY�R �����*��UG,���T�Qd�,UTR�UQr�r��1(��,ȑU���(,����+KE�5r�"�-aTb0��UV(�s
�2"�e��VT���0Urш�ER.5��2���˖�Jň��Z1��*�P�AI�U�m�cV�\J�L�\K��D��QA���bj0Ĺd�AV*�T��Q,�(��++J���,�%k5Us)�Yb*1@��(� �h�F[
�{���k܅��O���I�{����`��uc}G$�e9R;j�Ӯ����E�)#"ZG>I��1�d`���Y|:C86_7��M�y�G��.����j�YV�V���_f� ��o�aC�[��>�/x]�ǽ���@t�_��9�l�j�}P��CR���pR�WQ<D�����e��oϺ-n�yD�r�^i���y[�!B��d��"��R�T�Wu����&ⷼҎ���2q�
���~բ��ޔK����Ŏ�߽��`o���@��E�p�S���G@p�a�^#M!����"ťC��z��r4���j�uK��� �})$|�z��-�<6�5A�C`k�.3NQQY2���,D���\��}�\�HE@��"߽ڭa��<N]:xϩ���b+�n�!�%X�KQ~k���,ܾ�߭��XD���B=�[�n���MA��㡞��NFB<%`wZ��= �o�|�m�d'd�P��5hMBxv&�6�C�N�7X#����N,/WqX��gm������0��!���	@�X��T#�\!�zX��^���w�0933���*/!�- ��J���5���w�7���7�����L0SJ�=���˺�8�EOOU�]�E!������'���kya�I�;:eo\����3��ᣈBCM�j6�U��D[�s��
&��5���1��9t]�0�E�GD��kEF��3	T��0�  ��\�un]�8���'n�d�xC�$g_�f(Qt�.I�,���M!Z־�e2���p�U�\����%m�+�LC+����:��OQ��M#�QvGR�����UB/F���;�(�3���5wI��bٷ��{�xd��9��MU���.��������k�xO,�ԋ�G��ݼnJ�#�J�����&g����C�K�B�1xG-y��s�;I�Yl�][��d������U��w|��<<$+��pxOi����֟{{G��`h� T��8�w�\n�K��.�j8d�ޔB��~����j�q���Z�:��oP����v$ �~E�+����Ň�sQe_*sG�?I�@�,F��f�M��[�l��i��B,s���0:�F�'�h���@���??Rm\"ˇRg;O2a�rPoa�a�D�Z�*+�:
K�t�}�ƕ[�@�/}��E"�ƚհh�G1N�;���8�S�d�u��.�[:7}Թ�@諛Z�9!�A�U��i5�2����%�v��Y<���fIʶ��姑�-��T�ھ��ΚT�)ԧ����/�նՎ���h?�o]":�n��M�ګԓ�5��B}�{���Zduuֆ��0��� R���<�������8\jX�,�-��z�yt-:�������ٱ��p���YE���M�[�3�n�<W��^���y�󏩏W�K�n���a���R�I���a��[����á����РC��Q\������ي�%y�r\,���
��N(I�=�r�^7��{�s����P�=�R9�秂�A��*��,'�ߣs�q]���ùZ��q��>?ezVj����CF�z��1{S�W�W�>T���l��=��w��9���hk�Y�
c���h�
��ɿ]@�eߚ��5��g��.9+�B����;�Un����T��l9S�D���<�T"kO+�����~�}���r+�WO<�vyK��U:j�J�����b�fb~�a�T9Fċ��bx��;�C�.@C�����8�'Eޚ��%�+�{Vc:K�R��żTt/�/�a�T�zV��Lm�*���J�:Ι��ԃ�)�����5Q<�C�m4+�WՎ�A÷i<���W��J��ACi�����jn@��݌�s���{�T;�\�.���\s�N\��ږ���k2����g�ʵ�Ϲ�Z�/���p��f�)X�����LN�M�;UD�:��jWX�ո���x��8�L*���$$ڸr���M�HU*�����PJ��t'j�M�>��>�݊���v����11M
�ؠ�����<=���^�D�~�v��Mz[��yL���~�)<�Eq���wwiI^dOgLR���S=�!�>�:�5����I������B7X �7AT��ǻ�.���Yxu�d�+"}M�.��ײS��{����Цͭ��K�jX9Ֆ�(���ॻ����*�4���Gn�҇l����i2G�c�&��8���x�N�s찚kr�Ș�����*uP'�Ua�'�S�2e��}(oE_��i:�)�Mf0�y<{�&~�͵x��jeH6ܸ�z�hy\FBzT+WD8��k��u����p{��Ov�U�V�	t�0c��(��#d���w-�1{r`�U�fp}X��<���W9RW�v��q�o�ϭ3��f�.�:�q�>3N�f��7�9��]������E%�s�O�&;�rP�J1��o�޻��,�wt�����Rg�v�;�t���0lh��G,�|�<�^x��eK�����܃�ݶ���;���$�ʴ��˨���G(�jx�"�Ut��!b���Ưf޶P��J���K��mSv�Ԯ��:�r�y�5�pz�_.T�|�_:��X�=ޞ����t��m�*1SM
4������)c+:�P)}�}�k+`�-�����nT�udS��.��5����1߉�z���W����ꜥ���b)2<�mҐ=�$���������Z�e�Vo����D\zp�G��]�(�O��A�����8�j1�Q��WD���$��Wv{Qz�������{�Rz]��(7Ls����J.��!n�|�ls�+{�-P/x��Q�v��es��R�]Ѓ<��E��<!��Dv�7��CP�G=ܫj���jf�v)ɪs��,�+�⦱AyP�l�#���51+�r�Q��߯��l��F8�<ZzF��-�vq:Z�|f���4����q|;��$�tr^f��G�<�?u��K���l�-A�n�9x]�G�:�.��s�Wf���p�2��/�X�s���x��
[���fD�r%�����U�<��=��GO���ﳵ���T\^��<���M��T�dMœ�'7v����y�Z؞���WD�����(�I�|��;����.͙���YA�N���}��nQ�գ`�����u����H;%M+^m�a
�s�����s��+�97�GXѿl~'Z�|9�ݮf���pd�6����꼻m!�l�[�c�>���c�1�k�5�C�T�oO'�]km�{���{ճb��~Y3{���W�ƅ��1�џNw���s�+~"�E8R:�m�,�
^�o��
n��霕I��W���Z̈{�3#���
��G_
{���vcs^K^�%�O:�T��8M۠N
=X�6k����Ź����#��W�9�x-<�0��9�HG��B�Ci���fZ��\�M�C�:]mm+��H��B:��7�;W<wIc�S���:
Х&*�v���){��pXt�ӻy�ydµ�"��gz���gf�G-7��S7$��E�[�@s��������V���#������	�ޜ�{�Nlp^�nj�q< ֱب��_{��D�Pp�\�*�nb�s�4��'����:NSڌg����5�2���}r3��p�eoC4iW���}��I��@:�������.�Ӹ}��Lao�NyC�k��B���r�gLy��FlȆ����xQS�X=������̿�ALz���s�{o;���<�7{qE�&/[��W�n-Ǳ��R����{��潚�󻜀�x���q�����n�gl���^fY=�������.�g�
��{���o��69�}qQ~	�ڎ�Ӏ��@�������s�Cg%��c�_&��x󁸹�[Ago�?mVu2��~�2/�f1��.w
�MC�q^���؄�_�����~�;|�ίjy����&jm��,�]��"�Cts]p�|����;�`
乱L˚�Y�t�e�Xu��ߕ��]Zt�K�];k{wWW]��s�`�wյjgT��5�c��H�sx��mU�Ƒ�f��L4$�Xƈ��3I�%7�o�v����|�Ω�9.�|����r��i�������"mv\Y�����Iʹ�,�Q�md�s����J��������ò;��e�=��9T�ܕs1��,Q��Y�]+�;�X��/k��\��3n�Q�{��k��kf��`��h�<�r�.����N�k��ue��ΧcJ������a�]V�KT�< ֱ����_}or�ҍ����[NhUFSSm�{�n�ns�jٕ���蠛�v��#Tu׊�86:35l0�X�c�AM��nǵ�n�/��yB[�)�l�����jr+�g�G�O��^S7/����w8���KM
�}��e3�G��I��.�L�2�V�g�+yN�s衩�X��j��X�m��k��y�6�d������qy��������G��9pb�>��p��iJw�r'0ܻv+V�����=�\v��p�G*wiLd٨����$�]Ո�÷�ݷ�<{�����-�e`�|�L��-a�iҾS|p,��J�:��˓�J1��1�Def�N�V�U���'��J	�n��7���Z��9^ݍ�s����x�ÞH����N���A����a�U=�J�-m��L�/�ڊ�����;6U%y�A{w����u���}[Z��7�&"�J�]���� �N*./A�۟w�݋ށv]�_]��VI�q�K��rR�׵�,�lcs��2��,c:�x��L�S��&��l-G65��Ύ=�����+���yxÐ�v!>H�YFn�v��f�kε\90�*�cF��������<�U�n�`�ԌձG[պ��S�ݧi���!�})�N{,t9�g�}4SC�54��7'2����v�umݰ9쀯z��x�,��*��W1�y�5ҟ�]�c�Kz6woy�ɸ�`7۶�x��ohs�r_���U���j��f����]������4}�-���έ��>_CM8=�u��<����3_n:;�=E�5�a�{�em�h`�X`k5��8R��AS��HN�&u>i�"�`{��ǃVq��ײ�.�j�r�KK<����k�9�}�jk�C�բ�EKjȖ�{�r�C����xm���.�b�[Z:Ӡ�P�-\t���;�E�{KLw�6�+���L�sÀ}�_�/G���n�$Q��ۥ {N`�Fz���qN���~NSV�=]]�C��ۇg���:�{����=����R��r��hM׭�k�c[S.���Zv�O+ݪ{'���d�^��O\�v#�!A�[9���u^�y�g�V&.�2�K^�P���}����,yv���PZ�Py�b���׹xw����F%H��Gu�����x�������c�ӭ�������-�[w�����X۾n�Κ\��%�ڠ{"}\�K����S�����ٮw����ή��ޗ5��_�	��l�W���=/z�c�)gSay����؀mߥr��{��-	�7�%�V
x���Llj�*#_	U˜OD�fz��h��/y]����2-=�:>�ὃܤB�q�L�?J�Y�s�±�ω��F$)�̯B��x�tF��E���!�Z9�k�f�c�*���h3��'��CQ�^S�Z�oTC�4��v�7�vM���h�x;icKh��w��%��ë��b����
���N�q�MuكY�ah'�ej�η���UN� �j�m�m���gnK��.�d�VoK���@��7��]lv���2�0kY86����)m����=MPܔ7c�e�x�	}׮Bo�s,�۷7(�d	��;���̤��J���&��sfӨ(k����m���%��i�|�˦t�ư��}�Jvn��u�on���2�eJ�=�]ެ�ܬ�]��\]E$qZv�Z9t��!�
�,�e�0&6ڨ�ȸ#On��ʘink���#l��Wu�H��@	�u`�m�,�����ѽ�n��C�����aP� ��bξȭ^uX).=��KH�Ǻ�5��y�m�̝=�W>��X�h�]XF��s2r��AI7��i��-���rs�]X<���f#��&WJ�8Ѯ����RЇZ�%VZV���[�gf�d)z ޣ�k�wk	C����n�m)k>�þ�9./�;70�l�<?e� ����˟1�-a}(��+4�Q1�"F�6���Ʌk�wf����ܖ�����bR(m��59bk�'K�".A�U�ُ��i��p��;C�\���54Չ�u�^:�m8z��+��S�64@l��φe��m�\�;��(N�;0GT�=��S�ه�DT�ۢ�.#��J�x�U�Ǘ��{���	A�����8Y�Z�)Px��NM	͖y�f�hpN�JVqb}b�P� �'�yV�<ު���w��VqyLE}PR.�a�3��Qu�c�S�nA�j�_)�-u��[+q�E}(�J��ڔ��v���r�Ɩ���s�w[��;%�}�B�Q!�LѢwUʝ|{�����AA\|����jٶ�v��vVLilh�Y��Hز�B'�_+b]�mEd�+YT,�;��WP��A)a.X$�1A6ED��5�������}�_V*R�\�v�8q*2��JN����H-:�I.����â[v$g9c��y���6�J	�]�8ۋ,0u��b]6�1�s_C�9�J�]<�8Q �u��u2L���g�����*��
�s�7Jx�˂��\��5:Y�ks*\��t��i�[��ca�r	8�u{�VN��l
�)6�gf7>�b?�2�,a��"h�&���f�`M(��뒲鹕v%C{YbU��/'d�%���̚ˉ���q�6�o���d�3Y��+����_\�N���<T�}9�@�˲��h*ҏ%�wk����;f�c �2�c���武���i)[�i%/�`���7�q��i�k�L٢�m�Ś���on���v�a�Qr�m_HD�/\��?zkt��U�*��UE�R"(,Qm)#im�Y�*(��$PkJ��f8�-i���XQ��&��f\J��e�f\���̥E�[E���-��b0R,U���EAVQ�U-Pj�F���VQb��6�Z����K�K�h��`�.6
#r���Km�ŭE�%�[q��EƦR\�c�㍩��l[��T�U�mm,�F	9��D�e!Z(�B����j����E�1
5��
f+bѥ�6ʋb(�2���"��k�D��fYUYKDUE-�f8�2���j*e!QYiC)W�̫�b�A̹+m�TV�J5�e�-��& ܭ�"��r�#���e1\��j�k�J��\na��0�X������0ʈe�k�ZʩQq+�֘�EC2˙����q+*&S2UT�G(VT�[*VV*�PEJ4�fQm�P̳Fڰ��m���d���M{��X���`�A-�-Ss9�k����r�c���u)��(g
�#�g�M�G7����r�͔�.�H�Đ�Fjw�pj�n?���+�M�D�칕}o�ޤ����!��snn�Yoe�i�V�`׭�+���?�kb^�D��y87�������Y]z���ŝ�K��|��W��=�,�%7Ƕ�?�'4���9I�P�S�!m8Y]�]����g]3���:��&NW�az�]K���ʛ������k�T����4r�v��Y���:�)�6���'&��\���'K�+|	ٗ>�v�Q�jF���>q�q�W�'J�����j�ʔ�ǕNͫ}��ј�F�?o��"ߺ����i_r���`i��,�b׳�r�-?!���h<�>��zp�����׺��<�f�ŮP�s��1�Ϻn��8a��{�{={su��ܻ�������<��l_V&�d�f�[x����;�y�|��ߤAY���,N9��C"T6+�C)$i�k�(r6�[�E�3�\ݻ3�d�z"�1C�1]��-��h�l�/F��h�`��+�݂@d��6�ޠ�|0[�o�a�Z�,��a5쪴W�NJ�#��X[��1�|n�k����>,N'���zM�Z�G;�P+"E5\
}��I�V=����W#��l�q��t��&H���G-����?^�u�h�~�<ԾrYܯ!苊e��q�~�6nQ���h�@�@�fr�"���N���n�[�ZCO��k/��v�Tv�ՙ�t�X�37S��򵌕���tO��Yal%ogCO�f����XV��7�D�UZ�î��Psc\8�r��<{���ʑ{yI�؊ˀ�R��ȷ����0t[�|�.�F����5��[]}=~�g`
^��J���g��\�T�J��|�%��QD(��h�<�qpkdnwU��z���S�W1��ݚ�����ȹe)�j�@f����ӭU���&T�VA����z�ND[k]�r�̵�{�U�*rj�Q�X��,�<����m��ں=���%�4�v�,I�	j|����9%y���DqP�k����qt\�3=�OQ�v��F�"��[�8�Ġ�l�rl6�Rhi�;=J:js��,R����\+����ə�%'��c坹ѾCH����,�I�uHc��M�ŷ#ϨKt�@�JA���p�]����_8��/;��>����Q�����;]�s��LD����lRٕBy@�+����''z���װu�UM�^�Zs�OK�}�leT穁��p�~Go�F7^�/EU�1�����f���h��i���e�g�J��)1�+�<��u���WzI���+tr��v�Az�wK��z%���x��YNwP{I�syͨx�gR��#$ȕ^�.��עlgcq�;�n�c�E׺���>��r��:w����'��FlԆf+��*uN=,r���NW�8�,N��|��� S�p���q)U��<G:\��Dd�U�S�����]�c��(�b�0�;z�%ybrp�Y��߾,�9��˨�������"7�@�T%�G%�<<&o'�N�6B�5`|fs�M��n.ճ��2�y!z>/�	���΂c�L�@����:�	��xk����f0�p�t��J���̛~�a�R9B����}�9h@ց��ƭ�u�7GS/Q�H*���v`��k���#w�d����w"AT�䤔:A`s��{�a����q���Z9����c皣�|q�/�$���Ol����O7�c��e'�I�/��5:���+d�F����4S�R����'�����3'��^j��;Ԥ[y�#�2�K��E�T���_y�*�Թ�}@���=V暶g���à��N��O�Y��'P�%���o>�{˞}���}�9�_w�	�N�Y%J�x�%I�VO2�l�2u���a8��x�Ϭ�d��w�+�M!��q���;�<Iԓ���?2q�C��|߻�������Ϗ}��翻
���Agg;�8�̚���'Xjs̒�a:�dެ��'̞��O�&��ω4ɶ�`G��{ 	K�{����d�͒��jhy��y�����1'�&'O���8���l*d�+��)=d��c$�7�I_'5>�N�`T8��M>���4��C��=I��I��x��z>|y��w�/|���y����!��:�m�C_s��J���d����'|ʇ��Rz���{�I�M��]2Nzo$Q썏{�<>��\lz��SR�������7��X~a;=�����I�dSL�A|��|���0�	���u��P���'�8��T9��OY>���$���!댟2q6w>�/�y6s޽׾{�5�>�'�z����O���I�'�[��i��P<�Y'�u��/�k	=C�w�u?2OY��ì�J�����{ˈ�3�6=�z��d}�=��VI�b
[+U����~hţ�W'%�P�d)���TD��E�u���`yJ��sj��.v�Y���`2VjmF_Q���F>N�0'��%c�d
�v�Y�0��钠�jYV�k���e��C�Z���I��%�'Ms���i=jLd�:e���d�k,�$�+?�ԜB~��C�'Y5<�I�d�Vxkq'Pќ���$��wxu��G��7��!��?G8f��G�����I��>|?y�VO�I�R~I�k(OS�'R��&�T��Y'���u�P�xE'q�5�0'�G������j�r>�skr>��|'O��a��>d��	��l�I��OI���N��>�IXm��-�Y>a�5�C�����S'�u4~��i�[��=�����Ϸ'�������=S��d������I:��y��6񓌞Ϻd��l��ߟ��	ĺ�T�H{h|�����l��'�d� 8�}Y�G�r��ꧻ����0{޸;��'�X}CHd�:}ܐY:��;�~a?$�y�>v��OxXM��N}��2O����T�H~-�B�|�����ϯ����uܾ�x�{��H>�ԟ'�jé��u�o��}d<��񓌝�����0:þݼd�L�;��$��{��M2k�������f$�b�g�߶�ܼ]�L��<`�=�>��h,�q&��$�N��Xn�'�~`m��̇���N$�������0��so<a����:�2m���*�d:������s]�y��y�|==N2w�{�I�57�%ABd��J��VO�P6��6�XN2|���:ԓ���Cl1���9�u�z������<<��)c�򟭘��mU��	�{Ğ�t�p�f�6ř��x�����,��k��*V���䬟�Rq���M�	�O��ya�XM����1�=Q�N1��Bx��V���0�y��6�7�n�8���¡������rC�|ɣ�a��u&�y�T�&}x²m��q��N��2`۪�隈�F}W/-%QT��H�4{���wt�>D�����QA@�TOG¬F1��B����D�����Px,>�BQʶ���M�U�nA�q�.+>�w�i5�������x��ǒ���Ӻ�ك5����[d*c<��\T}��ܛ'd1�.v�3��?2z�9d+���}�d�+Ӝì:�bw�~I��;`��OPY��T���sY?$�I�Y.��������������3A�[�W'�m��6����O���O��aĞ� |�2q7��$�X~����J��u'R�Oq��7�AI�O������G�����
no��Ĩ���}���l�?2z��̓O��ya�N2�OS��I�O|��L�b��I�a��0�$���u�iYw�>=�c�����ʢ�����ϩ]1���z q��<��������W���O�?3�(q���M�0�	������:���2O��'|�k�'�q�ۑ��{� wi?}n�H�	s��ǽ�VC���:���OI�d�m�S~}���|�z�&�8�C,'�Ri��d��Oua�a?�d?$�
�7>�@G��}��5�ݐnw�̭�٫�����O~B�O��$���d��ÿa�N�q�'��@���>�$���~��z�O�8�d=f2u+8�<J�g���ux#�kM3U��s�=�R��P��H(;܂��N�f�{�8��h�a�i��.��&�XO';�@��2~�'Y'�Ւ�i���dĜg���'���o+��sY�w���z��y���i��<AI;����&Ұ5<�a�N%f��P:���'wd�a�ì�}a<���'��7�d�ay	���x(�����r�ۜ���0VOR|��!�?2z��LI:���C���mћ�q��X��E�Y:����d�d���N�a?2k�é6�����}�dtt��#�'.�w*�1�'�ӿ�J��C�i�'�,?�>C��J���N'��m��M�3y�s� �8���7�rAd��|ϖ>���_Lo6�r� +�����?̣K�,_����1��u�p�����m�Gv��6��
��UW��K�c��*fU�9��Y�1�C6��p���[g�S,��d���׬�sB�&
�CNm���K�CP#�^����2aF���؋��)�n� '�N0�}�	�~d���c$�?���%ABa�8�I�
O�l�I�N��I��Oڡ�~a8�M���'_R^`{ 
<a9ٟ��(q_|�W%��	�=I;9���'��I�Y:�d�M?�a>g�N�:���$�(L7g��%d�el8ɴ�	����7o���ѣ{��q2�l�v_�\{�:w2m�x�;�2z�|��Ì�a���I��&�i���~d������h�%J�a��J��VO�����(��_��g�|�:��V��l{�����|����Ę����N�O�����4����v����>`xs��>Af�wu�5�0�?Nk	YXy�52���Λ'#�ȞZ��{�ρٔ��m���c	�M��P��':���.�4�_}��Jʇ9gXu�s}�~d�
CG{��q'�,�{�*O_z:��:��E�����S�{��w�%ea7��d��锜@�����:��C�T4�ɦN!��'Y<a��RJʇ��2u�$���0�'`xj�Y�/�ٗc�X7��W� ������HV�~>��N oVK�$�d�'���Xm�i�:��N2Ꭓ��aĞ{�@�4��oy�hT
[��}����kV1�P��� Dx��wx|�ԨMs�=I�O���o�Aa�'���I�Mo̒�a8ͤRi���za�I��ה4��'�S����O}�����D�3�fw3U�{�<:�st��8ç9�PXOY�ϲu'Y�'�8���Nv��'̟j��:���0����'S̡<}d�h�8�=eO�Jf~_}�v�:#m^�yF��1�q�;=�M2m�����N��kq'Xk9�SL��y�'Rq���}Ì�d��'����>|9�IY=`~�����>�
��)z�����m����}@�C��S�q]Z��{ۊ��Y규ȅ�3��K�O��=x�br�{�nЁ4�"*���^��{:ʨ��u4L�Wܦ��o*��Cu9��\�A^��1$�ղ�/p�C!�\�0wn9�r{���1%k�Ɩ8��b�e�g-��G��?zH�q����I��06��MO7�|�:�<�Y	�a��a��	���&���9�8��N?$��rN�O]���뙏�������>ߞt���YY?0��!�~d��2�0�B��u$�~���'R�4y�����J��	�a�9#�Q�{���G��<>߫p.�__uH��+7cu��N=��~(~��>�{�ﶽ����<�T�H~��䬟0��Xa�'�.2O��h�a�o�o!Ĝe`k�d�d�<��$N��}��{�ӠS����׮R�߄�ǽ����'zw��l�޲�6Ϲ�$�6��[��|����>C�8�e�i8��a���6��q'X�y�����P߾hB]}��F��l{��FG�>�P8�{�|퓌�d����<I�{�	��&�RM��d�XOӈVO�X~���q���,�l8�~<;��Qc×U��U�lǇ�{�|z}����N�m�n�����0��O4��<�q�d��\�M��5�������%ABy�q
��VL��5���g�]�Z����� `yG��>,�������u?ky�s�!�3�:�׌=�����0��p�Ԟ$���I��'�?'���Xi&�w_�d�@F����T��~z�;�����<IRm�'�($�&�SN2|�g�:�I����I�̝C|��'�s����Nx�?2m��w�'SL�A�?��쟄_a͜���yld �{��0�>�d�RO�$�6����N2|����������>�u��<����&���8�T���u$���ߗ�Խ������;����=錞1Hv�B��O�Y��u�5�a��u��y�T�'_۲,����8��'����	�C5C��M2m�~�zβi�=���ŋ����K^�I��ᨡP/�h������E���z�w��	3�`鶀}���j�]�gy��Ÿ�)M���w-��ȉ���x���L�o+��e��_S��3dU�oT��\MA��I坱+jVb��Q�F�2nJ��DJ�[�)����c��x�B�q$�X��i6�bjw�i��,w�
�>J�[�Rz����I��$����>�N�`~2�I��y?�yǼ�ڳt�w&�q���D��Ow��&�8��{ΰ�aP���u�T��'X{��N$���)=d���$�&��I_'4o$Rx���ћ�����ǟ��߷���'Ι�t4Ì'�T���6É=Ձ�~d�����!�4s����ϩ�N%Bl�=Iğ2��;�>d���Qd����UW�L��_���G?4��o~��z�&�<J�i���t��OSl��u	�5�>f�8���d�!�N��}�$���Y���=gǼì��`}�����H��_L�+�+7g�X����?o����Nj��x���'�I��i�e���d�h�:�=J�ƨu'���P���My���8�Ԭ��`N$�&s'SL��o���=?s?��־�1�f����>��OXN���u��R~퓬Rz�~�$��0?���?$�5�'�����,�	�?��I��Y:�ɭ�)8������w���Y�t����pCg�=�=Q���Ͻ�����}a<��m��>x����:�|�3̒�� ��+'�8��d=O̜Me1�|�S�	�����r���w�yr��>�4��t?2i+�{�R|�����d����:�$��d��d�'��L�z�G����a8�L�IRm!��>ed��OŰ>C��M�>����w���Q10�����ǽ�*�|6G����:����0<@�'~��l����m������>v�L����M�Q�[Y^�����(�O��w�=���y���f!Y<Aa�`x�̞�&�m=Ն��$ۨf�8���C�y��';�~�@���ﹷ���i�þ`;I�M=�$�~d��:����ns^�fG�z�N��臂[*�Dd\F-�z���)7�'���1���Of�η���n5����G�ؒr9�<5��!�0�8,ķ�O>t� �-�J\�
�8؝�7��K��ZJ��u��c���{��� 7S��;��O�����s[3����
�|���a*
=�hVO�X~���M�XRM��~��ݲN3~P�'_Y��Y8��h{����������=�Ұ�uN;�λ�_�k��}��x�Y8���w	:�d��<�$��u��(L7z��|�����q&٣	�O���:ԓ��j|xLt{�G�7#�����
�1�e�c�?g�t�]6~��>a9ӷ�i'�M�	�i�lY����z�{�d�C�k$�XL�S�+'�Y?L��Y7����'>O�Xz�hs�뷟�w�f�}��ǝ���WĚa�w�J�0��p�Y':�8�����T?2|���Hu�;�c$�ONy�T�'�VM�@�,�d����~�߼�=���������x��m��Y4��=�HW�4�_}�d�+��a�A���N �9�2z�ϻ�!Rz���~Oy����}�����2���T�,������Y>x�ٖO>I��x~��'�Vi��L8������N���󬒥a����J���N��
C]�Oq��<�)=H�g�o��������qx��}�\�>�Ǉ�{�}�����������,:�<}MXi����S��&�q����=f�8����'�u����PY%O9N�m+!�g���ߍ_���<�@�_iWk3�&<6=� Ǉ�� t ��G�}�I�Oud��N��M>$�ϲ�O���冘q��j���N��Oud�̜A��x�;�fo�~?o�9��w��'�I���d�VC]��d��'��@�&�4oϿBz��T������XM=I���d�%N��0�hO�@�" ��ܣ�1BiV�3�������'����k�&�ug0�4�z���d�����:�����O�|��%d��i=k'�CS,����Ԭ�$�*t5�����=�����r�t�1�5�oP�3N��T";�����D��L�A9n���,,o�}�ssT\��+>w#T�*8:%��u�t��E[��s�euaC-�u�tn%�*RP�B�
2!��7-c5`q����m�n�R�<.�E�Y�'} �qǹ�V�i��XK��{�r����Q=��(�`��8�/g�$���W;��Sc��;M�̛��:�hi��M�5���^b7�''J��q�X]���+5���UTYj M�.�]����;�'Օ��5�X;;�Lw\8.iڶV�_��գy�O���**���79	yF�g.ks�ѱ-�{�J�Էc�i&��S�&^]�z,u+���3*��5ed��!�۬�����p9����03N�}&/����P��y����"��_d@��J��T��
��GBI��@��J���VQ����n�����B�n�JM�[|HsUq �ĮӤ�S����S�M�굗٠;n�mͫF�L����H�=�C�,X䜍���֯*�����ī�hf�](�����u_�( �tps��Sn��O}��+R�9WY`���40_���`N�k-]�ֶ⨴�Mu|�Eh#��!���/-�w��k	&'X	m؎��9c&[)��]r��_oZOo]o^aD����sXo��ǳ(�P��I8��w;Z�5Q��Q\��c ������qP]b�7K���)V�E�wh9aX��WM���� ���-"�巫�9�����s�Fq/t)�yc֭�Qsd�gno m��F�I�@����m&��]���q{)G�)��B��9.E���(.����|8�iC�b@
�����{Q�T�"�uB&^����+Xo�z������R?o���ƒs�tWl���\D��޺�]�k��ӓ��b�k�E+���/%Mu��]Mxi�:Bar�EK7ү��٥��Z$��ٮ��Z�3�5�v4��z(g��V�ʁ�I^����_2�V�î��[�t�NԸ��3{+sŢ�/7@�@��R`u�ַ��._+]p��mu7aW���cL�I>���xz^f�y��E��6���q�oeЕI�z��)+����!ۻWu��X�V��Z�:Ϋ݊�s�ɝT8���֑�>�1�Gvx��v��S�Q�����Y�&��YT�uGفշݭm2[��m
Ī�ug\�~=4̝���G�d�sx�� dk��%6fm0"�Q���Ӯ�{riS�X9ӹ�����x7:��m�C2# qM�����C�6����Fj�}�e��[��:�=�m�/���S����*Ψ� ^*����]%3���ז�Z͉JٲV��f�m��ٶ��d�/v��S5|`�Wь���!�sR�uWʮ*�(�]�0��!�C�)�kh^��`�a�D����d}A��%E���Q�mT�P�TE�dQJ�S(f6�5KU�(��6�b��10��Y
�(�j�m�Y��X+R��F�1Q�V�hŊ��j����%j)\E���T`��cV"*#Y+ATE�2�r�X����W�TG���T,R1�F��Er���6�b�T�V�mLK�W-���1�kUQF �j�T-�q�-c�PDX"�i[�6.8"�Q`�\��S.e)j,��b��Ub�U���%�+f4�T���$��EƸ������UXcA���B��P���*�*��2�1���+���T\�AEX֣Y�TY�5L��mUb"��-q��Lf0�
�����XԢ
�TZ5Q�5� �-*��5̪��<�k��1G9���`k/�&��v�_T��H9v��Q�l֎1u_[�{�1�۶Oiʵ0P5����M����z��f�������AI?����|������d�Vk�`N$��a�i��t�&�M�����'�]���d�>g�%d��t>J��'���~_>��y�y�����Ͳx����x�����?}�d�V��Xq��Y��0���?�N��:���:�����L����=k�yǇ�{�}�Ҭ�7��܎�缒�����VORm�2���+yП�P)���|���r���+��@G&����!�J��M�e̪�[��n�O*zz���+O3XyFo�-K:�W�vɾ������Ɣ�<���U��:h�`��܊f�鉮�>.�}��=����zI�L�R��U6�@��� !<�9n�l����aEߧM�=~������k�ÿk�rϓt̄�#}�6��3-����:�s{)��[+��c�iwG���zz�k�����a�̦bj��^s��쎦[�W:��ϻk��`[r<��*�=�<��`:ʟK�g����w��V���Mq[xZ�*���k��"F&!�n�C
O:וf,�stB�i0j�&�Q�h�NVq��;<_K�&��j*>�t_����U����[	3J2s�v:���R����|���e���s�\)ȫ��#{��_nQ�w~\�|�\:ia���I��ų84��>��P�f���_U/ �r`s���N	����5�a�Txu���*w�Ү[�2��sp�2sZ����Ѳ!����풽�24s#+��\/*��r�<��q��ё��e�ImO����&1kQ�isj��mT/�P~�
�#����[�VM�m��)P��ȧ�Ō�lXI׊�j�zV{g�ё�%��F��b��L]7�n�=�k���t�����}E��9�_�i��ʃY��Қj7��)�{'�u��Ǽ_�:?^Ӂ}�M����1o5�%]4l�}ӥ���x�9;y��Fƪ��T:�X�J(b����H�;u"�dgVo#l��թ؄�,�3�Ϭ� �:Dlo��'�g�V�T���[�՛����j�	Rf��k�t�yU�������;|��$F��u0�Z���{�#�7>���K����Y���g��U&�X�T���:�O�k�� �v�l���/�e.�NrX�+���C�ى��M��(@죹Q�g8�� �{en�(q��[k��[;���n����7�۵ht�/w�dM�5����e�Y�0xM���@����c��l�Ȃd��{�W�{ޫ�jVr���v���S���[Şs{\��g��ٖ�M�#�����]��èQ�>)�ԭ�n��:�'�AM.�g���i�J=��7�ډ�� �̉Ʃum1|��7��^���|2�a�S���N���mҮ��m溗A\C�p뒷&����{��I�`خ�|���_%|��<��mFJ�U��hw>+�h�t�ۍ�="����+b��ұ�iw-�����[�c2q��֣g���N�2���{<�st�yc9�D5n@�s�|��~��ݎ����E���Z!>�ޛ��͓�s���謜㫥XPˬh^�*�N�������s�l�7:P��:�-�����������q��n�gk�Z�By�f7"��ݷ������f��j{�`��*0�@�Ӂ�=^�j{&N`�1}�����y�F�mso��`U1������]�aax�=�	��A&(�gP���',}�Yۉ]�9�κ�2p;yH��e�2���Ioj�W�0L�B�;��N\��M�M��" �օ�`'����J�����s�����K�%�����";2��ԧ��U|��ەOø��{I��i��rM6�I��d��R9Ө8�җ�Lo
cF�|�/_��׋�=k�ݗ.#��M��}�of�[�c�[GQY�ڴ.�g�l`�F��χN��ʏG�������[�{W�Y��[7�v�uz��q>`�3���
�=|��r�vy��c�+��������C�m�O��*(��w�Q��Jt��p�̜518i��{�c������b�m�_����*U}�6$�@�ǃ�,��7'9nuӜ��棪�Z���fVXn'Bo5ەQj��[	nň�#�P3�罻k�53%���3�/�n�ܡI������WM�+�pX.f���Am���VK�iy*���� �8!�����9#uUСX��LP��Ś��)���q�1�c;��HO�තf��Q)��E]��h\���m4g^��S����]��rk�cy�m�A\�-�ӷ�L�+ys�F��+S3�H,f��VRT��3���?.F�pO���g������ӏ~���r��QK�����Jku���{�����t��)��wi��� j�N�M$W��T�[�.x��G�jy���j�+�m�v���zT)~�[C�(��j��$־:B��b�����oj�yk&xt
�͒;6�I�+58�����<��dm�6���&���\��KF�Y�%�ٕ
�D��U�qX��
t�G>����[��O�i�u��� �(�`��k gBq^�(�Zr|�Y�VQ:��"�J�����17V�Tv�=s��͏:�:h�&����}��ge��pէ�gP]g��c����N�K��y��<uuqo�X���ޢX���U��򝇙�z�9f��m��eyyb�uݵ��Y��R�J��x����7�}2LX�%&EQ
?s>̷t绪�~��i���<)���Dmhf����{2fe����˹��t��sv� �;B��	��b_U�c7΋A޺��D���A7gYC ��'<�+���9s��S����/�Ř��VK<��8vͬn,?;���.Զ�L�ow�{���˸����w"�-���XSX�N&�i�u^sA*��¬{3�+�X�s���lߨH�r3,&��]���em�����7�f8���̥��8�~�UZ�xs�,�E�v`lx��V̠�7��ؚڊ̰�7!0�T���	��f]��>���x�5WJ�u�s{��^����'CH�9���zIZD�C���D_b�0Gr�X(�Od=���\�t���GJ����m,����B��E[х�����)ՔP��Tc(-j+�1jy�V��=<�*`�=�4�ج��/9r�e�]5�LX�����4�,sj)�{��:]�giK\Rzǧk�FǾ�x������l7�,�pgڜ_�t���W���u��ݡ�W=�%m�QR��r�0W'Bt�J+n���������{1]N[OƦy�.1�+����P�3U�i'��x�܂���|;��.J7�9��Q��5��XP��$~i�C�eKˁ�c�&0)���3���;Ϫ�fgCC������
���	Ӭ�˻�{P������W�aIG��ít۴9sUs~��,cY����65W�*|N:�6��^D�w��� ����Yci�O_z������3x�ϭ۬���:�(f 
�^�K��{hr����}����j�|��'c��_Jcv����N�I�7�lJo��dg�}ٿ
��vs1>Kr��%R`�<���;�9K�f��}gv�5vx�uЧ��E_Z��ϝ�Sx��m�2��[���]�t͞SU�Q�����E���;2��y-v�9�o�j��<��i���yq�G9ueSS�eq��zKUoo=�᩻~�����6L��趚+�weCmHҪ�j��x��V{���^�7Ԕ�l�ά׹I�a�a�U��$$�nP��Q�ޕ�L39R�Z#��M�ut�[�Km�ݑT�X��W��'ؘ�ک1�oJ��yC일}�A�x�:ƥ����Wd*����P�B��zF�9�1��k��t(1��j�3,H�7�T�F��f;R'X~���֔�Ks��31��i��4��0)Cih�WI�>bz���#ML;�q�teN�r�oU�O�\S�v�\���i�����������4�R���c�
8j��W켤;���Ŧ�[���l�C\�
��x�Ӯ�%ǚ����U��u��Tϼ�J�^���Yݍ��e���m˖j4�.Ylrݠ�VdJ�\ϋ��ym_R��<��j1>��[9>��l�`�VX|��z���)�\�ȕG%�@�Cp�L^�+9�t���Bԑ4%I[�q%t�s���Їh���j|E��׹�չODghx�Ձp����]G:`q�zVj�1���ϒY'd��o�߹�����oy|Lk�w��a}�=�y׈��8=%�5����g�����,�wh�c'�:7ڜr�+���Y`G�_?{>�s��<�T3%��W�^�c�T���j��`�����C��\,Y	��
�!5<kA�$8:�
rz;��S������W�;�+�����0(5�᱾��˃�j�t<�z�i�kJT��q�i��sc��*(�؆sm=!���Z��Wqح��O��XC�o��eŐ9Z�k�삡֎G��j���X-%c�ͬ����i���T�Ȋ�w�]ton�r��r���Uq5�	B�+��1��{-��uu���v泯̺���KyE�I�����\L�H��e]nw�����Dǒ�v4�*{�U�'&���h�Ň���Ǔx�z�����;���꽺�'�7M�����^�8\�������7X��N�S��ĵ#�yf��t���:˖t��셛)uZ��͋�mJ���h� ��JEg��չ�?p�%]�e�+�56~M~bS��gO]yz/�>^�-[Xc�=lVl�Z뻻���ܩMz*o�y��~�\�y�P���.5@�o��FI�P��Х������Viy���?x �: �Ym5O앙���fD���&U��׭�W֖r���t����*�8��::v#�bi��k��$��[���m�{����x_#���֥�gSaV9q��fmK$���ⲝm�*t�z�#��k��T-�k;^�}���e!ƺ\�B�g^�����;T�s*�l��ў�@��{M�G�d5J�\������mt�%�h�A���&���lHm ⺃��pV��C�)վ+ךqY�=����*��K���������## vz#VK�;�u{�Uy߼\�4����-I�p3,&�Y�c:�Y�
c��x��]�����}G{��9���~{���GR����L�̑򝇓�G�ڰ�ѭ���V�@T�����&ᯜ��V���%-�X�V��L�!G��S���~�z�OVN˼iZ��~#�Ú�[c���5���n|�\�K�j�:���]R�Of�������,�u�{y���L�{2M5~��Nt�Us���_J�<_ZY��@yUa����c!f�!�vg͇!&�y2f�%wt��k-�3f�LM��������S�x�K��,��͸.��}:�p̛�ٽ7Ɲ�>�p�������_"��E��<�HO��f���[2ܷӦ���y<�}8-r���m���c'�X�/D�~R���zVlA��jD���ǈ��3�@S�)�t/Fի��Uz��W8�J(3~��76�"�nlx�HK���`�}w�5g$Tc�B�2�Z뼫���m�"Wj��녩�E�/c��A���]j�Tɹo��rjw�,}w��";(aCb��3��w�L��1��Ʌ/Y�ӧ��v�ֺ:��s঻4Tl��^N�!U�wT�jJ�2��!�`�j��ntv��N��˺�����Ԭ�iWk�wK4��t�p�`��|u��aX}�Rvo���k��'v�Ơ��u�wy�ƭ�.��4�g��[XD�x��0��oCѴ:8}�!.#F�;�N=�Y�tr��R�8�Y���R��|��61ڱ��{{���r�6��ʱSҧG-i+l�Q�g�Ә���׽N1��E�"�Q �0�K��7�U�N��Wri���F0)�/���,�
[J�����@�BF���H����#�xP�G
X���y;\�&9eJ�Ok��)��Uz-�'VQ{���H��0�uU�hds�o��hf�F��)�V�U���V���X�-��7WөNU����6透t��i��]ǧs�k��7wz(+�MN��P���K�S<\a"���C�Κ�mFj�t�]�=B<<�El�4��\�Ѧ�Ę�����;�p��E��TMvN�HwP+R�����It�l�޹&r/�s:�n�6�:����I%���
�,"J�0c;X��qŊ\�i�J��^Ρ]V[��t�����}���kΦ�:�P�G*��^!�`�:o*�>ՎS��̣S3{��N��<Nj�B���N�K��a����C6�+ΰ��'�+��w��$��M��T��W-ӝ]p���B����q�`�2�3��Ƹ�Ȩ�Iy%vk��7��`.�-f%�^��W��O��esi%P�s9:6�ID�(���� �8�u�n����Vp��yS��1����5�լi�{�_sN���R��}%��q�� �weŉ�ؙ�e$b��o�uA��JȨu=V ���9j�J��[��6�xkzQ 9E�4�u�O^�U�hr�جX��)b�� ;��ʝ[�w+
�Q����31���)X�o�����G��䃗s�����w\ՒR{3��e늓����:�2��ofӺ��%��t�N����hJי���c��C���}�nGk/L�P����w�i'>���ߓ�+�c��+츎M�d�@��r�u39�jb�r��8���@�^�M���aM��N�RC.������CE-u�:b�M%Vt�0�
Ztm�G���U��f�f��4�Sx�q�[�S�*0������8l�W��-�WnI�h<�7w)����2�i�DB����Ү�6�Fe��ĕ��}DD�t�[�;&��J0}��ӕ ���n� V&J��a�6�C(�{\�����P�(��zʢ*1b��"5Ę *��`�H�m�e�EFV�fdF*"�QcҰG(4��"�\�QƩ-�eJ��kQJ�P�TPW-�A2��E��!PPPVC0�s	��X婖�Z�1+J���U���*�s[n��U̕�Q1.Qj5�e�J5���e+U�D�D\�Q-*�� �-����Z(�Z�EXĭE���)"*�`��1���J�b+n%k*KJ�c1�
5��Ŋ��U̹�Pq,�"�+neB���R������i�3�B�����d�U�+��h,�E���m���Ze*�[B�Z!X�9p��"����[ImUZ��L~����IΡʦ���=�PY%�h�:��J��s��Ggr�}�\��k%�!�{���,H��ɜ��9v���+��=�[�3B�o��~[>���.P�1�Z�w؂{���a^AV��`5��� �=����H�Z�.��+�d��R�8���0����5�������,7�\��Y���~3��5W�gk����\[]����0�:���rm��bcM����3�*4x1p�>�u�8X��\$��og>楃3E���t� �����9�Y`cY�Ƕn:Dlj�J�N:Pӥ*{�N���g��&�ВV��:�͜*{��ὀ{�`��:aS����G�������nu�p���[{�×|dG��뷫^T�Q���닗^I�:h�^���*LٙV�Up�%U������7�5�Ea����|����k"��ս���\��L��g��3��K�E~�z=�m���U���>D�BCAc@���~P;]�f}�k *_a��wH3^��x�ՠA�=�(
�ʵ�K�`k�u�E���Tf�[;�r�s��r�QyjER��ret�dt3����`n�-�h�Y�}�t���ڜň�=}LGv�m�fl���!����j���R�9�Y�:����{����vX`�_{������`� x�oV����c -�h`bX~#2@��8��+v2�ds�V̪�о�j�⧀�V{���1爞��*c���'��nU{�_n�.����R��Ǯ����c"=}�V^�m�㓶Urቃ�g��J�gm;�bq1�m�do�1�7�8\�)�n��L:��/�.nm5~��B���Z���Q[�=����C���i�r^�_m#~�l<�X��j����Y��+�|�<Z��#��WG����Z���e�:�m_Vv˛@���$�s��m_��ڮtS�i�@=Ml��w�a�p��2�����iW�Ěw&�j���������_I�_�S�p�5�5��ܘq4K�-]�t�7�)��	{BP3���%�A�>v!5Bج������kG�V׍�c����M���n�h��*$u�Ekw=mK���C��[jD�'pZ�䮧fz���T�v��J7-w&6dز�]��k �8]����^��zط}�����wm肨�4��k]�V)F_i��L5��Rf���U�V��>>3�v�Y����N��G%yoa�{;淬t"��f߃���M��`^������{hN͙.{���=䟼��c�b�^ˀS����)1�X�[�̊?oU�7��9�r����n�gC�0�>��+Uu,��ꓞe\��)NK�2���ux#����۬;�\;F\t�{��NDs�{�<�gg�׷)��*H�.O	t�����@xZ(�^�#̏}��\�g}��Ǖ�Ϝ��NM_L�J��9!������o�b�Z��q�W�E����_In����5��ߟ+�Ɵ�NI����&Լ��=���}&Wt��-���B��2�D�W=�v��hM�_�\]�׽��K���]��)~&z�a�=k}$���Xw=�B�9�,��FV>���s�)�J����$~t�t�P�4ؼ�����%xh��ٹF(�}{|�ieA�u�Mݳ�3�BkEnnq�ߕ�nKy2�
�$��3���^�<�l�������̳R͕�s�KP�$�y���n�#�� l<n��Ű���wەqws��WEԾ xxS�����T��|�!�o@��~��ݍ���L��� -{y�v�y-:��}6ݱ+w�J[���VjqP�j�{�˽rI��ѶN���r�tI����یqݔdMp"t4+���bN�N����i���%�`���\H��;<q����Xh,�JU:޺���S�(}��؍�7�qK/��� �T�.v�X�`��;|�'Z����é�r���:��%�^-T|��{�����;�(F5@��\�E�Srx��*u%mT�?7z� ���N�i6����<�|��t�@�, �����Yo')O,5}��S�p�,룧��P��-�����ѻ<���������J6I:2Ϫ��������>Ը^���x%��9s!p�}f�=�b^o�5d��u~��g"4�����S~��@k�>���-\��&9w3���+I_����C��^��=�D=�rՃ��2��� BY��\g���oe�u����A�2�_.3�D�$Ž	!q��r�mV%�p}ͨ7�!t�ļ��؝�^ؓt<�	u��'��Y�F���8��G�T�:�pP�b��.�RnsfW� ��=S����\�d:�Kb�e]F��Y�_�w�,J�Nħ�3\���U�l���=~]������G�Aϸ�d�-�R��$S�5�YK�Z=�'�p��q�&�L�M-P3"�BͭL����v	�Nk.�~'j�Dj(X��!�U�֪���vR�Ư�^G����]b��K_l��Y��q9Z�**���0O4�t�4m2��~�tnZI��C6ɑ�����t�l{N{/��J	��$%�ע�r�x�? ����)��T���.��>���|�X=�Z�l?Ki���������b�!�U$����0~��v�&�f�<c����oǫ�+��pxRUG�x�RP_�j�t<48O��Z�ax��w�qY������r�x�}��i���������+Ǥi�$u
5{MAQ`��|�Q�礑1z�n��݋,*�S��N�E��=�Om�{�"UG����5��l�}�͠�Ɨ�M�ϭ
t�Ǵ�>d3;��@@��=g����Ք��J��W�w �Ĝ�M�n�j��a,M��c��<��Ԃ�����.�YlPF��'�=��s~[pַv] ��Q��ҕаU6�v@ީQs��L΢�Fub�C%fl{��R�i@.��f��W��o��ƨn����P\ľ���ϻ:��N>;]r�7�x 0��VV��Wd-?L�꛱P��\3�V���j�{Nct�]>�ʗwq.�=�������_�������4���]���غm�^����Ǘ�"�S�
���&���ey��`TU��N���a�][}�ɋ�i�х���jf�p&����W���ȼ����f+w��L�U�v��]s4(VV�zJ�=e��.�m_�#3y[5�fj�4n#4?)��tT��S�s�* �^�>��-J����/�\��}d����K����ٔBr�p]� ,mO�lWcֹ^�x X���p~�a��������#����rc3��IR[T������R"4Ew��g�b����{)���t�)	�G��̋�^��s��LH:��Ss��&ϳ�Y�%ޫ�}F�wݲ�y=�ɗ�}�g���N�*�iE�Yx�gF:�� v=�
�/�+�L��Y�inX���)�����{�M�"g<s.*Ы
⪇F�٪	��x��xkc~����R�-��]�YT9�T:�J	u�ޕˌ�Ŋ �4��t�u�y��p�����mm#�b��B'ez��˯x���v&i�r��sb�r�˛Ċ��FT3�e%,.W����-�D�O:��`$,ǂ�i䡻B�K++V%!?{�{��;o��;��j+�v�eN�,��4=�Zr�����6��x7Kά�Z(�:�L�H�܅���'#V�w�n&&[S�ӕ5�+pS��o�"r+�&�_�v����i��q��n�K���w�24F@G
L�Y�b�+�qA��~>�k�L�+MD�}Ճ�])�Y�e�5��s*+�]�)D���`6��3�L�N�cV�R�����/(p�Ǯ�M�k��t<o�t��<��A�[R�r{&<}��3S��z��N#�;����:U�|��i�Z/�x�����f}w���h���D˂��G�H�`�ݘݒ�M�~	��7��^
�y�T�2D	�0D�w��"G7�z8y�j�]�oK�3�Q�]��v�3��fԵZ)T����)e{"cD7���  Eh�݂_�c�r�Ԯu�T��3~tC�e:��`��'c�3t��b;�(4e\�Pd�d W���j�6�k�j��Ϭ�����/h�̣��	̙O�
U�)��c��~��CZ�����K������Gw�gBT��(��[�|r��j/�r|E�C���	�^��N���mR�$K�s��ݸ�I��3���`׳��j����
V7��Gd�kX���Y��(������bTD��9W�J�����������뫼����������墑5������>0O��$��$�
ټs����^���r�R��G��8v�G�;(�vj]������_ۆC��n�*�1Y�KT���R�� a��}��Wx�,C�/lD8D\#�/X����R�6eN�ܱ�E�x���ӌ��UV�(�#�����e���.����H�[�C�y�/Ki�k���ɢ�U�;e��X��Z�su1ݿ\8*���1���]`�=MkW9OL�|�>ν=	�Zg8T���	q*��%T�Pw��o�!)�}�
y�;��}v(�}�W)+N����U�FW�� U�ؙV�ʙ�N���wK���쉜��܍ⰻ|�%(�,V
\]#l�R�����/�h���]qwh�F�e+A�j��X�B[�u��i�p12�4��a
�-U����R���H��i���`ts��r?����O*�;;]*���?+"D0��
���"�����cܻџH�����x��#\=3݆[z��7�Z�0�Է+k�2�,�v�p�8.��{Y�Yb��Z3��~+El<��jޱV�@�x1�2�*7�{{�Y�L�k#�:՛T'[�=g� �t��C�,,�lAڔu���BDս	.��C P=��1Fj�̓��,��<=�>��{�G/m���o���Ӂ��9�yHd�����*�q��TB��,��n�`=�y2��K�AE�����=��v�����/��Z��W����E�Z�v��e�	+����4#�Y*�g.�k��:z�����9�W[���%����J��r�D�c^�f5��eWy���U[�����t[}ga�fg*,P9L�h=�$rG����41�v����K�u��j�X�%[�g�A�ךi�\9���|M�u8j"q��Uǈ��x8v}�@��"��.�@��D{�xnu�&POݸ�,���z�&j��e%��
�)��`���0�á�zNF��P�ª�0�U�'�7��{^��p�
���0��Ϧ^�Y�c>�}���֓ծR��̔0O4�@xo���\��&yK����*hy˧nӸ�3њo.\^̸ys�X���@jaW��9U6�%p�.l�_ U�o�d����!�k����k��K��#kشHG���"B����.���Y(���#��G��*�Ø��ˎp�ޒ��o5��8��F�O2'}��d�Go����&�oY#n/s�Z�8�#]h
���F&Mz�xGf���|�>�j�bh�f;��+�M<
Fr�'r�lR�Y�5�{�{�e�9i��f����\��=��ulli2�Y�I+�Ҍ����C��^�*��Y�S�$�PS5^��mtʈW��G׹.��F�Z�>�:�*.늺t>���&͟l��j��������b*��<\U����y�܃�~D08n��ko��δ�5!;t/��g/xՊ�꺋�8�W��a��� Aθ0�r#5��f(Q���P�Ga
�4{wko�C{u"����Ixti
ֵ���!Sϱ�����\+o��u� ��`�[3�es�g$l��#�P<9tX���}mS���Nm�xS���VB�WZ�p�&u��8P�X�F�L@t�"$qD��B�H��o�8κV�q�BK�jV�
N�8e_�P�׃���38/T�x`�49 s��Lr=�H�W,��\�8t����c�|��ؕ����d)`�f��!\DW���� VUk�����yP����N���C��׬ɢ�(Rt��;+�Ͳy���q5.�j���>~F�WQ�ԓ����V�𦚞�cΚ�7:�E����Z՞�2N/a&�b��ٚ�E�5N+!�|ަ��O�QН54ˬ��x�i�l�J8�Gػ�5``M�����a�}����{�M��Hhۥ@��g᝹:v�̼�j�e7������ɿZ�v����)[�r��<U��6SM[;ܩ�+�9{O��:��������ɤ��6��z^չD�l���wR�٠j����U�Ƶ�p��5����lB���(9n`�c����ک�s&='d�5�%Պ��(�"�c�G��;�����Bq��G t��EkY�[�t�V�KR�I�Mf�k.mVI��a���؂|tP���b;�7:�0o���cZ^'5�e�.�m�m����B��u$�*�q3W��s���|Mh
�͠���ì�u�:ա%h�Z����*/��]�9#��rc0s�ݼP�4��L�yj�W.�Ӫ��#�hU��r�2����Pd\/�N-��}Y�)�B��W�1]��n룟e���� fގ�r�W-t1�'y%��2�B�h���Yu��8���|y����7O2U���F70T��ʦA��V>�E&1n����r����2�6��"ns�����R��#	�J廤�,�)� �`� ������-�*���릞j��%��ɉF�7:(V�q;r��Y\w�)���IT]��f9�+7\�����5�XS.C0�A>�\41�
�cy}��Fƛ���֤kW؏&;k�b�JH<���F�&�;ru���:��A�x�`��ɦ��e�NB��hs.vkz���eŝ��X��5�83p�j$8��6P�*gaSf-��)�kۦ����A�.0���x٨�y:ov	I���a�D�pw�4S��ԗ]���ir5��u���H�����M�0�΢�n�vu ,5�1v��h7�C���;S�Nձ��\ĒoM���}���Εo�wW	�k�B�0�{����6��u�����ɲ�d*���5]�[W��*Ex��*ǰt�h�I���{�|���%����\%Üd�\i�G�eQ��-`c�?<��8�TE�U��šg!WDn�H�s�Pf҇m����b+���E�<m��Y�g��ҥ�V�r>������r\AVt��;�DRދb�e�4:��\�ӵ��ۧ��+�n˂�I�Huӷܐ���B�r����ͽ�ɢԲ�"�z��.�QZ�n��k�"�E�� ��;&G��F����B�&=ˡ��{iC�H��.��n1���ZB�5}4֧'p�Z��9�V�4X�q�7*-�F;7�,=-�6�+���t�x���离�ϛܬg=��@��+ucm^] y+�l����eY��i�*�]t2ش��u��G�ܣp_s9S �}0��A\>fڳ�VYmebe��Z�,U˗3"X�cSXUV)����(�V�EZ�(�8R�QAch�8Ѷ�R�pl���*#��T1m&V�卖�ҕJ�2�q(ܥ�R�
�"��+a�q�ƙC�\�ĸ��33�R���k$�)���2ء�&6թ�ʊ�X�i��Ņk*�k33L�������b�.S-���fUT���ER��r���L��QqTr³-*L(e���˂቎U�ˌ���q
�㊕��AAj
�k�e�X
U�VkQPF�X�[l[Y"���ZKl*+h�T(ԔJ��)�%��ADk(���DR
�)�Z%Jђ��Re���2\��f�"���e��J�ێ1eJ�1\�QE���m�m�IU���,U����.~��>���Iq�;`��K�/
]&q��"���t�`�,f���1,�h]˰��E��3a7��; �B'��?���|R7�jv	�K���
����GV��|�9��2�2(왎�T�Y��'.���Փ��ײ{�~�,q�wF�1�}�(f��u����'\���mu[uE��Y���H�p��p�L=���G�K�����C����g�ܵ~صR�Z����8�V���u�('t�3�xvu{�p���9�WpXS*�FC||��@����a�藼�G�<Z&|\(h�8���u��%�fҶ����'�5Y�(�aw�y��� ��{��lV
�l���|�ef�be[S�|/NMj
�(�n�}4^��l6�� mi��]E~�����pi3]_˪��_gXf�)�\J�Җ��q�=nÁ�T)�F{&B皴�^�Y(�6W�->��{K�U�`6��3�Jrߎc<�Z�%��p���픩��T���*�`>>��A����*ڐ���L=Sl�SMnb���N̓|�j{�t�Ñ���4�~*�"�{�Y;@�o�o��챵n)��^to���=y�����/�u��ߤI�/wm�e��S+�e�<�$�QV�4ĝ��j�t���]ITz�Z��]��T���n�xm�yS���;j��?t��q�6�k���}�u)ʢ�b�R`�j:z�t+����ʉ*�2-h3
z��ܥ|�����ܢ����tze�~�fp6��qVoÑ�D�jF��*��}�J��ă��{(W����q�^Ye�.��7R�h�9�`�$S�{"c0� @�`�.�`��C��i�N�s'Ny>��}B�n�z��#�ݮ>����v;e����������͜�����zz�	��r��DG�Y+��W۬�SU���á�}L��J�8E�WX���Zԫ:Y�n煢��.+�rI��L,7�w­U�,z�{��;�$�ၻ�Y�����T���;�K���g��n�m�O[G�_��E�U�>e�\,F<D�;��䯽�M<��]�,{� Q��T��}��򧖪vY�Ox����b������<�~W��rw��XZ8�O��x�J*�ϡ����Q'$8��A_Ni�E���S�q®53�3p��+���YGK�Ul9�2���&NM��q�F�{�U�Y���d���f(	��`i��ծ�b3�s��mPLؔ�Ʋ��*w �ν�G���,ͤ�»:[7.�낺T��S����ʗE��|�/D-X5���	:��F���pl����Z0bɑcZ�V�p�څ�跣cޫD"�=�����:��4c�w��c�_Zз4���ht�:�����V.�3@SUֵ�&衜$x��ѝx�"�Y�5��x{�s��9��Q�p.>Æ����ۗ��h��r�k� m�'T�Vp�\���jy��!1��K�g��yU���`�ţl�|��..���U�H�󫐐;G�Fqg�+�Jp�P�Xx!K[#�9��7
���L!]e�kg�)C����3��Fk�6�y�4l"d�z&��O*� s���U�9���!�G��D�jH�U,YQ�e�k��b��]jU3���p17�[0'��C�^����R���q����z��2�3e��C��|D�phF�p�Tz�N�����Ø��N.B�Y�GN�D���o�~�G�S�#�N\wｸ*�� :�; ��]��fq�qU�Ŏ/�i%�r�\�V\�u�p���4���唩���к�dq*��e%x�Løz�A���ѩ�ҽ������|�PpbY�2�S*�/��$��Z��%�m%x�4�̚���y7]Q�ٽ��#�r��C�x yR� H����UK�P*x�U�}�C�n.�(!u~���o�ٹ#@����OZ�8��uɻJНy��j�h�M�F��|fd8��=�wt�R͊�"#�ݨ{E�j{l�n�*�=�a�^㮐�}WV�}�H̷ں����Wg��;�N�����n��EȪ;2�rW1?��_{��A[�u?������4��d�&��@j��f�6���AoI����P���0��Ռ��<�~y�Ӻ�>7)m���S�C����tU��J���%�O4�@x.�N����9��Wr�鼺^�1HR��
����E�ˇە�X��Jz{S2�ٌ�]cŏzn�Q��s�k:��eC�Cɏ��-b5�G�m6=��[X$!�-�{|99��¾zɾ��W���Q����w�%���4�*�pSuG�Y_7�.��c�K(�ل��.��{<$nϳF�<�C<�����Ѩ���\�x����l�4����"���\D��kd�,�+��8!�b\3ch(t%S��<S��x����7 �_�#��I{`��:���>Y�Z�(���JȲhb�e��89�Qqs5��f��y�9N�T�>�r�{�p��Ό�h|%Y�<9w|&+�\��62�ղ�*�y� j���Wx.�l�G��M�u���8B���h�#��ÕtX���ڶ�����}�^aUT�r�>�0eKN��[�k�o$��r$�x�f�o��v�IR����k�nm�-ӨJ�x=��U��)&f�{�LY̪� wکX�\�����T�	mT��[�fPô88$+��ShhV�ގ�Q�Vs�l�����x�K�Mu���7����8�Thk����c�'h/�[�bme�f;b�3n��ȆE��\��7X�z�f�ޞ�����te�w�X�g@�pt���G�D��މsc�c����V�r�*}R���*���xs#���qSf � V뽲T��@�ghҩo��������c8�+k�e�P��R|} �:��j�bBUP�C�Tv/,�o{���;x0�Sp�/�GBn86�5CuX$�	O�)�Rx�̇3��r�����qfƫ�&�ό�!���J(1m����`��\�E5�\��-TZ��E�i�3��JcN4�.�ѳ��O�ʥ���z�OO3M]����[�${8�]}y�S��ɀ)I�����r��ʦ�01�+����,)��<����o���ӧ�ݎG0ʬ�C�U��Ǆ�8����U�/��.��f����'�ʿf����jc����̨��P�)�� tk.�n&!w���zf����Qh�>����ά+J���ʰy�$�p$�I}X3_q���s�v<�xm�*#Hn��陋@L�M'g��$w=�2:��5��f��<	Z�Z�Kbc������f��G��Q���qp�e*��o&�VndV(��ʡT�]J�Z܂��*"G-���W�W�U���E}�<���f[_)� 3�V.5/ց�#4%;�y�Ӑ�q�M��#Z*e���<��<���(o��U�Y���t}l|%�Ժ� u��9_y؅C8�<������v�~nLa���LH�68�<��@�u��� �n�~H<��&,k��G�8�Tp;N�w� vLK�`�r7�ŌB_kFx�N�TN�2��e�cyy�Z�+vA#*w�,�S;h�����!מm�7r���
O�S�H���DH'�y�}�5سj�Xj!��1�{[��SO�����E)9��=Y"�+��f �"A��q�t�w���}C���m�iV�sB�?�јf�u{�;���1�����h^^�R����N��L��z2guv�0YU������������QӘt0�Ϣɔ�P�Z�3T�_�F9ű��T����Z�.�$��":��yh��ᬱ~>���w4I>E�v��1����-��N*���dvm%�T�*y]�Iau�_m�1�"�����c&��>ݗy�z�#�U�N�]7��mfgp�����G��}y���/z�0�Dec���v�����ٝR��Kᵶ�vG��BcQ���DKE��ĺ����ĺ�Ó#wGujǂ�d�B��aE�Kʎ���,M8�>��� | ���P�#�����"
�\�
��d	�T�ƫpDpyv�툸��Bӑ�Us��"��^�2��G�N�֥yǄeC��9�W���A�2�f):Z�f4*�<-�׳ϵq�2�7u����Z�5��+¶���.Л����c1�ތ_%��.��=�Zö�ᒩ.L����'�c;��A2S��r�.�����x�����<�|����ˊ��W���?f!0�[�V4�2�k� e}�؅_f�hy����i-+�����y[(NSNx2+N[t6��ٯ@��zNQw*�
��B�U�H���#�_w�GPxD{�˔����~n�
>����3���g*�4���P���5�o��CB�[���y�d��x�BC�IU�V��T�"O]h�������z�G�a�H�ǅ���0�;n�^�~i�W�Ċ���T<�'��bo�`*��yHd����ĨW��dd�\;���L��gH@�aQ�\"��i��1��n\v�s�~���z&�Aeg;�"�xo��>���z����P���E]Xv5m�)엮M�`S�ӽ���)�rF�S6^��ڭpcY�� �k$̺x���b����ʒ��}S���$�y�����'&������_��g��Ṵ\�K�m!�4P���٘�%�Gm�FU^ʻQ�{� V�s���c�5�(3�з,�$�ۢ�.���l�3�SX�-*�u�1fjw3�=��sKy=dT])v\А�e��'�p�%/�t����;Ze'�v��8��Vf{`~����&;�
Lp�Y�2ਨ��<D���/�Un�E����7|��Y��2^�66�]v�]{%���KL���[�2�]A��ب וJȁG�B�Uc�r^�>�{g��|����^Y����wL�W�FlgР�/����1��9���c�y:�O)lS���V	e	���O��*}��c���oS
�L@vz0��JM�J(*Q��u�u}~>�@��N|'�
�εoҨ��..�7�����墫S2̎�;�Dd��KA���ZK<t�,[��p�5����ǥ��Á2<�D�$<���[KuTӳ�>�waN�nWjlϦ���C�fm�xx��}gE%�b�U�{��jC�,6w�61ٮC(1�Y2����Ʃ�Gs��K�r���7��h�!AF[,D��N�%"3�.mΘ���ت��<)�jQz��rtcn^�y�K�+R��)O^�aT3�xs����Ytr@E�T�Vn��o_����k�m\u�����n9;�uc��W���]mf���i&0w,�q��)qX%�;�s�߇���d�(��eG
$X���n�u�U��j�"�jq�9u��9=/~ɹ{��!����)�z�M���oTVF��u�2
��#�E�^�g�:����k�*���ֆѺ�Ed�����LO�p�����ǭ�]Pc!�}[,B�y�!Y<�����v��#=��,�>�t�PR��v|�<QvG|88M#ƐyV�?�U�{0�݉,lS��kRVJ1��S{<3�<�>��i��XHо,�����򮭈��0(���3 �<��g�]�}��0S�1o�ڊg�����[w}��+.,@z�@���ry���U�)vMZ�Q�ᾷ��.6M�iT���K�n�;2��g�6k�:�/>^�	�`�4ל�{zng�ɂf^�[���$L6�M��w�x:��+w������I��H-������ѡN޾��߸�(x<�B
�Hcb�v/,��S��eUIpQRf:��&5�$�#��8�л��0�>�@�����rc���U��n�$��/�.��{��v��ڌ�}Rܜ�^ǚ#\���60�nǕʽi�;/�oy��6ZX$�'S[�xfU�qpI1qpS�d��A�{��F��U���T�62���r�����^8t��m����P���n�	&҂�G+H�hv*�<w����ؾ	v�&�� +��ݖ�k�X?�PB+��:Nsv�x]u�g�P��U.|����C��_�>W�t�u��K�X�����@n�d�=��gPv7(�qa�O��n��ޒO������k��#H#��C�և�}�D��CFyǄg�|�v�-��;yH7G*	��m{�nʄ{ضu�-Ď�����+�S:5��12ژt{��zrkPV�E�t��<TS#�kt�������`LlKؓNJ5��t�,�ÕlS���z'�]v�f�Ɇ���2�t�jbݎ��J�E�J��>1%����| ߪm��9�b�x,7��֬��i�Y*w%Q�����BFq�3h�s"8��:�U�����yJ$U�!#��ё��x�Y;ڤ��[I�Ȋ��z�K��/K�290:$���N����6�]`u�7C-%�r^�������{�{W3�f����04UN��M" H�DC�q���Qq7׍<W�r&��F�����{R�h�'?{�����(��vb?{�̋&��̬�.Ti��3Տ���o(ٺxՃ�z�%{�Ͱ�+6��Jk��ů�;"Z�n��NI����]:����u��	3i��
n[Ǌk�ܧT ܓ��;���Yn�Oz�GE1�ӱ�3�9���1�O=��@FIlA�qwn�:1�ihE6�3�
��$�,��wU��AH�IK�+r�@Ծ]�D���x;o]c�;�L �L
���0Y�ccf�:��=�9���8FN��8>�Ң�*�鳄r�'�]/vV�����+�#Z07�N�y���㍡4d�9T�ꩰ���ƒ�Bc��}uo���+m|�WGQl�'�1lN�o)i�>�ד 1y⽂�.����i�{Ȋ�_�/!/;&2z�g�')U�*���$�CV��9װ�T~�k-C�|@���Nj�7�GB.���h	�bA������|:����ѹ�`*Fc�ZlnR��
�gG[� �D���KH�(ЛW6���ߒ�9��Vf�e�C�_)n��ދ�(�OЄ�a{�,G;.+�9,�cΓ{H^0E6)���d\�U�������T{(p��3q*5���K�v��s�j�Z}��{]�$�n��mu��H��ش����E�>��v�@�Ō����J����̔������[tŏ�].���󿅨/���ġ�E�����Օi�
��e"��WyN�7������p�X�fS�$�0�]��T7�	��H��lQ%��۹A(��7��&��99��|`�K��c�5������L�ˏ��1��n��"�K��jN�l�&�c�!��Gvh&t�_>uvv��j�;�� A��v��b!�Z��yIA+�=��T�F�J���`��N�� ͳ��J�]�T|���k��l�tUՓz���i��J�Z��&�0n��IpҔ��}M]4����1��h��p��;V %G`�Ȅ���X3�.�vw��C��K�����I�0}{���{�[�S�h�����K8�E�\��Z��ٽ��-�OWEa�"��*�w�<N[7���5����R��\�t3@���n�r�����K�
�ze�!��� �������C�f��ڎ⾜���K�QyW֦�`ŻG�ԑ�-��E�c@�Mu-E,����	R�ܘ�AQg)���9t<�s�H�g�JG,d7��t%l��3˴�.��0O�y]���Ӈޭ��\�7�p�����9�n�ǉCG*�%�"�d	���D��a���Rsa�BiR�Έ��������.�t��%�r�]���Ų�.�U;�%��(^ÕD�[��t:ڂ�s��Ū�x�LoF��QF;dЋ�e��9Ω��@��V�u-���[�����2鼘���극����2h�:�7���a�bkd�Z���h4�(�6烜;x�@#�����WT���s��ؙ�u����q2�}�DU}�(Pi��T*
�����`[ADT
R�l���YTeb��ɖ�YY1ƴV
"�IZ�m��̕��0�J�1�k�f$Yqeqm30���*(�*�����X-���cZ�I�QC
У"��kU*%Ld��(�+
��E*c1bc#J,Q��k1�IX�(0�jfR����FAdUQUf2�.[mb%a[JV&Y,H��*���S,���ԩPY*�T�RTX�R+lP��Ir�f[*LC2�F�P(������F���lAlkTj�U���+QeIX���X,UX
�U��PXR���Zŕ�-KaY�`T%@��T��a,�`T+T`�*�ŕ*"��J!QE��V*�T+ �����o��߽��oT�B4:	E+��wZ��H�}�f�۵�(7���UF�R�ڰ�r�
�K���F�e����՗����+5���N��0����h|�]8W�����lA�FJ���E�+X>�x����(u�wn��뛲�vK��0yU��7��e]�]e
co T�l�[��ÆZ����W��� �y�޽y��+��,��ͪ�l�\S�$�&��I*;F2���x��u������jlz�T֒`|xtn�Ӗm%��*}�Ick��7=��̮��1Z2�ݨ������ڽ����tDZ� W�X����. o���ץV�6k��BM���O��{񝲚�i������Q�G*ǁ_kR�
��� A����
����R��lI��vU�������	�؆���<�)j-\���[LG�k��\��k�(f�٤�w~�/��\�}r����/)/%�/���/"�^����<�y���ǟ��-��GŷǏ�D'��~�>��FٱV�-t��{[�Uc@.�!�D ]a~��(�&���f:{b��Ua���i�Bg��yU���`���#l�R砺��w_Nͬ-t�m�]�i�9���Ľ���Uc2?<��3�5����Ud��`i}Avl�nЇ�1�[/�x�^����/�����R�b�T�w0A��	�)n�yW	�̬���2�� �MldS��?	������R�K�-(�Ҿ�猞�m�*��d�@�&Ԩx��B��F�NqQP���44c�+���F{S�]��C��v�r����m0p��\}��"O]h������W��~VD�bA絞���oZ{����:w��xW�"�)4���猝1=耂Os�C&^��J,q۰JU���n���J����	�.���< F�ph��j��c��_��v�]3e��W{��Qs|���yeخr�ʘc�pK&�r��،��b�����l�3��w��ӂ˃���l$�=���7�K�*/��ٰ��ac4o"4��Ú^�Z�8�TFԦ���]���ϼX��eE����PϦ\�U�O&�X�%[�u,�X���ػ���y��*Y�?7�D�Ci�3��#>�Pj�v*N�$2�p�u7`��w��z'rsN8�
UQ۞7��h�+w�笠����� ���h��h��4�^N�ջ=˥�CD�F�'����-�R�;Zﰋ�s���bA�؂��9'�$(�����7�{��2��]S�m��"����d��H�w�����4�
8�M�@�vR��¨5� ;�4�|s�^|
9CB��ZW�u���&�P��l�t8�q-W|,��X�GJ\nI&�2͌��s<Fp"�o���_}�Vސ��"�����0���+_u�{�,�����	�z���5~%��<�}�k����h"F���6�u�&�p`u���-b5��i]R�cҮ>h�F�C�أ������s��)��2�HV��5�\��d��=�FV%�ϑ�M�xU�u�R���
R�똊��>�V�P��؝V�`�F���j>�*�A��٫l]_'��q���{3:ǅ�=v<(/�c�
CxR��p�ܪ�B����xwG�}��R����ƻ�����gh��L��X#��d�S�x�!�O�..f���t Y���=.o{�][\�ft(�ND����x�A�l�3��SHV�Z�������!����b�^��Y�굜��3�C�f���(.����x�.��@�p�MƐy��OƷ	[����ҵ�~>5�K=U}n�7����T4�U����F��N�W�J�r%C�
���U�j]����s��$��.�(�SǶ���0Nw������+68 :r @>���X�=�oB�Oz�X�l{�+M��/z�87�l��5`}0�K�s��ASgcEY�Q�W_��a�z����	kM��;zyL�%��k�W��C�����\׎w%x�w<�J���|�$�k��)vh�4.��/6�ON�,�c�b3����y�M�}=���"v6��%ť3�w'CV7y�����$+�ʩ�˞�^`����&��w���w)�d���	`_@��RU8�h���t�}��_9y?T)>>��ZQ$���\�}ؔSn��ѱ�}�p����<ԦxEi���F��D�%�F� �� �Z�K�����x_���\g�I���0*���~~�c��c>�!Y�t��]|�-��%�7�C�!�h�;�,����L>�@^tyT�I�k��aGB�7U�>��{��X��W����\�
�5 ���}���}��<�{��ꔝ�f�T8�\�����F^�x�r�
��@C����Ϋ�0�[�L�lX�՘��Ӂ����a�Av��o�;��]�l���!��x��PU��I��6Z����ã�´�z���~�������s����2:{��0&6%����0�Sԩ|��::�0���8U������ �q>{�����,\\j�v�	�����JK�Z<������i�����CL赽�zu�P�R�#��ͣCSc���0 8Z���ʔy̱��zᷫ6}a�P�	�q4C5n���f�׮�kǀ��}���IJ�)`vD��BS@j�����;�8��ե������|w��
�2�΅�ךq�!}� =.�t�ۈcgbO�u�r��^�͢�2#��t�D�Z�����q�$q��j�w�|�L��D+=��a��a��7�K�~kfEp�Y;A��R�.�u��_:�im{��/;�Q^�UƦ�Q�PW�_l@ESۜ�	��t`h���c�摡��;��R>,��·M"�@Ӓ��X�2�����{��Z)I����O쉈}{Y��]-���ˋך@��k7UF�T�'�B�"b=M�f��b��ᕬe��R�>�'/�R׾�&�n��VL�}o)A��t�Ī�b����@���GNg�C�y�GX���( xօ�22����9O��_L�M�K!��\�d���C���%n^VѐHߢ��:pG"$���):NX�Ig�}O���IaWQ�*�����۱W��^���l�N+r�Wx�{����;�# /�Al ��e���^5�+�Τ�{ּ[ي32>��N�Y9c4�6�3�q���UV�����1~f�i6:��m�x������:V.���qQV���NKUj�6��$��q��IƐ�q��ۍR�����b`�4�P�Yr����Xak�۰E+56]�Cj���]V�8��㒟ц�3���\Ro�#�ݢT�@�@�s��h�S�\v����UQ�f��~3��k�����~��$L��~ʶE��Qtr�6�k6b6(-t��ԷXۑt�/�����݅�\h��N��_�^ᄹ��;W���r]z�n�xKw\�״�m�{�r��u��J�j��p�||+����.�X�1r�_Ә
�����6�0���/v�������^� F���qeJrߋ��/O�E[�x�+E[$z�.�V�!9��t�!�3�;�ɢD-0�c�ɱ��
)��k$!�NqQP�ѝ X5����:�r�7/uT�~�VN���� ڥ+:���yo�z'3 }AA����k��OX˲,^t�&vl��|F����D� W3���W�9Zp17f������>8��]�K~y�Z��;]����v��<B�
�����O;Zs�N"��Z�m��d�'�ͽ����*z�V,O+��
	d����52��r
�>��
:9�� �X�L-�����cݧ]�;�����V��sTYJ�?#B��J�p5�A�j�<,f�������L��˓��jWϨ=95�K������v]��v9Z�j'��Y�Z#���ٍ�N���w��G�r0j��4�+�|mkS6��fr7�9�ݥ���� �%�e�<B���H�f�=�U�B,�Y8��B^
�Ee9�!io.罝�mk���~J�z�3fZ�:B� �v�T˂��*�*x�5z��"���=x;���$�jSѕ3��k�|w��u�$(@�L��|FK�5T��o�-�R9�g,>+}0{��t}՜��}�oGnq�j�Rn��]��2�A�RzI�[Os����������H��=dC^u�u��	fV��?'��!jOm@S�VЇc	T<����sl�GȿP��q�F��4`�}�0�i�X�Ԡ����2�������P�f�mM��;�k�W8�ax0'��{L���
������_��Ĥ�#��x7�r�9=n��'�G3�[�����"���q�s�m���M�G�[r������l
f5�+�h:���	Ϸ����j����������U�M��W�;����=DG�HB�r�_���%�8����o�{��>����<z����O-�/ȍ
����Fk�z���*���W�v!�*�0s��H�%n]���՝h��s�P�س�̑qwA^N�T�];��Y��m>��M�N�%�h�BRP:����̇���]���狷x)���u�2�^�\9��i����_;�����PV�����Y���^���bi�CQ!]L-W)~NLiy�|�3���Vu!�:?<bKG��!Zu6�c!�ow{������~�	[|,�֐�7�eyҮ��]�M#�du x8r��}� �a<�����Wں�U2)�wZ�vlHW�y�YM��i���`TQ#B�'h#�Ç�܁���2���������K�uV4�h��?ߚ�§;CGVI��z��Ð��HhP�77��:o��<�{_�P�v�%#�"Tu�K�Jg����Հ9���3s
�ޑ�dk9��秶hػX%|�ޖtVzWt��[
�������������I���Y�~U�=����+z��t��]�G��Hcb�E�����0�tTI.�c����p��a��whE�rY����)�όΰ+�c�������:�I.�uڢY�G�W�p6�+\�E8�А�>'k��+q(2������/3ʥ�=R�����3�^�-y<�!]��~i��k����O�n���D
�-�����gPw��8\�ER��?9��ˬ�KK"`:����S���[����xrT�B��fy��[=AL���Ű}n���t��c6�wi��.���*���4�ʡQ�E�����؃3G]#p7o�_:jZEU���uy˳d9�f�Ω+1*��ҜO57y�]:����=Y�qC��!�o�`���'|\(h{"{�^������d���[�1:BN�g�}e�ZWة��ԓ����+>�LL�ja�����̿db���,�|#��J-���/F�6>�;�q��`�����,ؕ3��+�k�o$��xs��q��>3����5�&T�Ux]�Qd�I<#�K����+��Od��(h�y�:#�@�ja��}	�ӚČ�a�D"Dq��v_ x�D��]��d5��ԏ��峙٨�zwI��BC�odà��
�#x�X�%��V��Q: e�뉱�t�{wڶI��vY��J�0e���/)���Q��o�����"��£A��<W�����k�c7�7��ء�m'Y캺��Xߚji�׵-V�Rs��).aV7ti8s_�{�g��3���Qx@�}]����dt+��Aֺ�G�=M�f��v8�C��~�R�o;�=s�lP���B!G���ɔ�ʘ,���>��b����V@���ҟ�c�0{�k��V]�l�v �^P�ϙ���i�
u�^j��O�:R7���Yܳc�����<ǃ�"2I��0s��cm�j�j�x���"��}�fG�.��ɮ�IcxG��vJO���ʁ�\���_,�+M�3��4��BF�.p�0>F>�L�^_!��,s�����Q�i�|m���&yɅ���'}2������*��37�OA�ϛ��	U�%*��,@�ܜ4��$�8���:6)�.eK%L�����s��hL��E��=wDA�K�$�6�XT��KʬX�%����$��9#�=e�T��Ul���H�\嗀g����1�g��C֪;�2d=b p���SL)�eP���絸"����-���jTǑ�]un*�q�CD-��]�n�鎚�Ea1�Pwm[8.: _{<�K�&sM��I�[�����;�x�rg���έ�2�G�&��u���?��TVl��+�|�`/���ϧ��#6S���f�aD� f�be[�*z����4�z}�*Ҭ���U����Q5�7�ޝ�%�G�l4s�&��DŌB[&�:p(��B��F�9��8IW������<�O��t�p�h�I�f�<I�၆N:0O=D7�6YO�#���3�(n���)k�����J���NI�\S��M*(�N=��/�������A�|�+5��^h0wu��)�h�m�Gxc��T7d��H�و�����rDͫ�uE0�ok�Jծj�j�����d��P2����ᬭ��ʓ�h��D���Z��s3�u�5�m�k��8'����n��6�Y�fk���ْ��ր�7��Zp�E^q��[��bU��r��.���Ņu���f+�aF�н�{��D�M2�d�gL9����N݋��	h��r��#Om��)Eη�Y�N��zk���l^��E��l�m렋K�o���B�k��д��]{s���,e,BSy�dזӰ�
�ut;	s�m�t�n�j�2Q`Q�h*�T�.�/�C_AD���PƆ�1n�}I�7Ⱥ���h��3�OK/rT	�t���6���n#-<9���5��|�;q$6�W��j>���Y&P舩��RI?#��W7�֍O]����S�0��Fc�-g�����5Ԕ��{�	�0M��,\��wW>h\&h\vq�aX�[X�H��0P��g^����;du�\����b��"�> <��r
f��ݖ:�2�3��I�q�7�K�[��ؔr�X2��Ð�2�A�^լgT�ۼ���*9�A�wm�yOk��;���o�ECL�mo"�a*��pK�zy,�ϧkt	�D��O��NM �tS37�Y���;Է��˧:�e��s�
4q�8�k�|j�]e����\o�!!�s��V�vgk��5#�����p�	�qEf�eS�wr9��{��p��{\��$�S܋ �z���[�sw�F�ܺ�P����Fj=y�b�nWm�l�����ڂ��a��`���um��k���fN��d=������>4.$��;ơ�W�����&�sB�u���#�r�a�Q��Lr$՞��U��� �;P܆,����ͣ�R�;`Q��E��g_ۦ����X)�v����DFw�}�	�SƸ�}5��M�/���,YW�r�ʠ{$]�i��Y�����8�5,n��)�W��븺(��7�^%��V���9{Z��A_��n�m�5�_��nuiǘ�e3������r��C�&�9L2m:)�+��7M;����x2r��{t0Ŗq�v�ǎ�f���9ˮЅK���Oc�u�l�A����K&��;A�J�m=�T	m�F����F���ԌܛTOo:|�=j���Ԥ��m�|�F�����\�2�O9�E?�����Cu�����x��$.�v����7YR�9�}��U���9VA�O{g�] ���i>��Y�Mh�ga<1֌�x��;����*��{ �;V�������ss%�ZY�N��J�b;Nrf��.�h����̼UqH�[�J��vZ�g��$���^}��w��ϑ`i���,�Em��X[@�+Q�AQd`ԥ�
J�YX�eAb��QV ��iVZ0X���"

�Z(V�E��B��%K��ֵb$YP��
E-�PY+QBV�����T�1
�VD��,P�
�������Rڨ�R��B�
*E�%E"��1Y��
�Q*ԫP�
�
�REZ�
�V���B�b�TE�XѰY"�,�"��Jŕ�E�E��R��VJ����V�kZ�P�DQV�F����h�m��ŊF�(�X�RօEYP(�F�IZ�meE�eaiT���(V
��X�R���[H�X��X,�#[�E���B�VT�m+J�iPXЭ�T�*{� �0=Z���]����'4�Q�Ւ�Sw����J��{uK�Iy)+���t�*2�S՗���
�ig��������Z�6#M#]�A� h���Es*�J�*��'+N&��`OsT�[�c�D����<�,��X�t��Ǌ�Q�r�C��p}Tz�5�c��.�����=2�d��ږ����!�=��.ˁUޥc��
����<I,Fv��k�����2��\O��}��w���S���f��y.Ȩ�]���"G+#�,�����ﺏ��O-^%���Nγ�fg*,P?T)1ު0Dz�F
ٕu�&��߼�_NY��`����`y	mfK��ab����Æ��2����Ci�$�.��GoaL���Z���z�vft�:���5����t�iƗ
�����8)�n��]��2�A����ʸ�'yi��y'��2�Dj(X�W����=k�,g�We�t�Ѫz��r4���T�$ՙ��j��ݒ�P�,iϺ`5m�HR��}3�p{N{-�����usF�*�DpĻ��ν8!#��(e���$מ?��۽����C�]*��nnv+��&�zK%��i#]qw��.�u�[i��Y��v)�!I�ݾP�-d�;��b[T�i��l�Z�)B$Ӵ}��{�ŇJ�뮝x�c��k��=2����c�7��n
u�5b�ʸm�Y,�T�����q�#�M��^vf���Ob�!�뭇a���Z�z��:-�q�<��?S��#��[������s�t|�7�O�u����sq12����:Wl�*1�"��m݋Ƴ9�I���\o�v���q�$1 ·LE�8J�sU1��������z��}�����3���ڎ�NQ��z>ٝ��	2:zP��"ɬS�x�!��3��^�������+�5=ԙ�#:{n�p�V���x�Ih���+Z��bx/���;�V�[�y[�H=M؅}<�ʠ��̯:U�*�>���.��	���M�w����ܖ��m���V�o�a�Nm�����Ǘ�.h��`TU4/�'h@��������6tQҕ� �<G�s�AҸ�i�qh	��p��&g����>�R��:T�ðn)��>��B�F��$k=�V�*˄��Wƹ˯8R����xxH^���'�U��{�W�θ`㱁���(�r8G�u�]�*�.���I8н��
�=��\1��RCoZ�K|m�ӣ�m����u��Z���n����$T�-���^Ħ�_�yz��r�R��"aGHL"�Y#��ܒks��V`�B�X3��ہ��<�;��gwVa0�dl�6������ ɂ60gfn�n4�չ��vv�"|���n���Zo4���hugň6+��}a�p����<ԦxEi���Y�y�x�x<�.�m�s��ꂫ�;���t6K,�eH�Ц%?Y��`��a�(��7��N�O^MS^3�=Q��F�Qc��&�51@�!����}�ƕ[�A�O�|g3M<�q��*�b;S�\��ոlx^G��}����>�PJ���t���U]����:�z�_���aӂ3�9�_*�
�P��w:Д��Z&U
3��}cv��FA�;��v�zUOm�S�փ���_����xD�X&
������T�ja�~�*c�Ee��ߙ�౤猝�±yX�9��,�c��c>������!�0�3l:K'�Ժ�7m�l��.w��G)XW���Vz݇o����,��,�Ih���e��o�&vz᳒kx�H$�6��b�/�w	�Ӭzy�D+�Ȏ2	�u�9S4��#�<�uT=�w�E��ä��I����a�x�[��n/؄�9���Q�\'^��y!P��h��iY�mY=]3�aS�5��f@��ؔ��m���,�b����9��/.2�A2�W^ҙ�AL�f��](����)殳3��ï_]��>aL=���&��[��X(��5��j̧
ؖ���t̛���n3j·�E%���O��> �譢�}n)��yA^�l@E���3�g5����A�gݦ�����%\�wc�HЫ+hY<�4k���Xv�x�ײ�h�9�`6r������<"Vg�I�
�L�; ��h�D��]DL��3�7l7�<k6� �ա���8BPD�~K�ןd�0e̥T�d_K<J��b�ʡLi^���7���W��r���c}{i��c��:�ag������t`���I3�raa�.z�\%��#LH����-���p��{��;��*���B���9`V�_Ig�|�*y�D�#�nxNP�wE|���/����+�ô�9�V���b2�[ t `	��GU�mU��\�*�c�(�`p��BT��ul��%.r�����L@�]�"�Fp��G��C��П"-p�
��u�Vط^���Ip�O��uS�Y�q�ԙ�~ػ�%�oS�G�.��(ᡢTmBf���꫃�U�D�ma�3'������;d��X����~����x�n`�]'\=*�kg�'�Lʬێ*���g��oK�h$\�v��fQ�-Ӻ�!���KK�ču��ܪ1]"4wl3F��e���$3rODZ�<{�65�ܑM�E�f������
a#�� �^j\�4�4�wC9J��635l���U�幙[�%O5q߱���`��-t��zK�|�P�u~k�1�2�#q���= ��lL�qe<�'KN2+Nn���G� �5t�0�ݍ��N�o���q�9N\�p�Ɍ@�J�:p(��R���k�TT(o����FR�W�cc6N�l8'�I��e���eB&��%����1�-�~�;���y3����2d>�Y�ʏ��Ƒ/�� p��Es*�J�>�x��Ӂ��-�h��o���ut�	�y���S���ܧ���P�5�0�}�/�,�#F�5��4�r��\{����_:Ӷ��^
jh$+��}\se�}k�G)���W�a�J�F��#��&T4H�nq��� ��3"�j��w��(Q���S*3�W[����"��˳aՊ	\���'�>��P�3f�2�����w�g����u�g����X�~�Rc�`���e�QQ�n.�o���{���c��3;��R��d�X~�JU��4�i��u�&T�<�� Ox.����%?1/jӳ,�n\�e�&��H�B��K7��{uz������+G3����_f\ʇ[d�ae�o����Lo2Up����DK�Ӎ_J1���q:ҭ��ѹ;s�;���1���-������V�G��x��f�p]�U�<�����}3�fc��{g+�;ܐ� 
����!�թ1Y~��㢗Ws�%}瑛z�ћɼF�"�5�-a�1bN%�7ʈ����k�؇��ٺظG��p8yX��f��	Iı�wl�Fȇ����tcْ�P�,i��h_nj�
��Í+�!gծ�ڌ�����A�x�c趧�dc+l���
�����&��~U��޲��~k
�C�$�X��,V���K湏j������"B�<�`�Ms���r{��ݣꂢy�k���➱���%����K�Y�h:��sq12������/��zqD\�u�q��c�[�^xs���1��6$�@�hHB�ڊP�u[�b*�����y���\�Yz��4�G����>�cO�2���Y��EѮ�%�؆���l�6&u����z�Xxnr�娄5���1B���J���<b��͉KG�4�iN�tܩ=�yOn��k�� �3O��؆y�C�o�:U�*�)�x�쎤
��mKK�s9�2�Q�̓EKA�KÕ�kL��^r���+I���{��u�MB�+��ϼ�c~˗~�Bl��k@����Jtt�)��!&n�X/&U�X6���'�q�Kၷ�$�±��O�x/�Muo�y�;L��|�\L�'�v�Lk���U}�^@*�5��sn��kւt�N>��j#��SbF����_Gg�7k=���C�]��%|4�a�e�b�i�х_a�W/O=���u=�4;�[�kwz���BF�ɺ���t�x@��@�F(�$�g�M[��j��s����^g�0b:{��I /���5i�CW��q� �O�;��kv��u�00MIƅ����&.��V̎�O'| 𶊱Ү�LpZP�ى2��Y�¬��^"��:S�G��a�^u����6m��h7.���~nJ</�"4/�%U?Y��`�v:��ò����N���i�����}H��/:�*�U�r�p��"͓�}���4��N����Y����;Hg�^\�!t�}��Uo�c#ǆ���� �� V�w�����ؽ@�&?lqv��*�y���*��Ng�p�l��p�d;�hJuشL��CC���-"�����">;z"�O�]������'�i`�F��|��t3��a������o�}z���Ĳ�؀Ϋ��º�,-�OK���gҰ�yFn�y�ۊG�4�	��&�9�.raK��*;�uc��jH�r�]��ֹЃ��k4���/}���ky+̩+yۧ:� 66j	���[X�N�[C'<:��1ӫv�r!���}���;]�G��8�3]�^t�Ѻ}SE���۽Fg�pi+%].�N�c/~�Tz�Gb����pʶ+�.%�����3�A^���.�9q K��w}^G\�V��8�)8e�#�а$� ,��睈T3�L�8��`�����p��:7%p&&��+%^,Rw�X��F�>��$ek{& ��
do���6�A�:;���Lv�1��+D&� �{j��]�6�SO��򂽲��{s��3����4�^<n,�|�5�Y�D�dء��.�_��v\�axx�����1U�K��v0�z��Ob�~�')┶|f S�u���Wʍ]8Vp�xxo����҉�㏖s�J�XSW�vdV�N]����`ʹ���=�K<J��+����p��Z�V�JE�{ڥ���Z��T)V�r�;N]M=S�p)�I��Y�}P��಺��`�����®U�GW���=`gQ�qc��$&\.��S�m%��*|ed�/'Z��qir�+~�L�.����{�Tu��L�v<�dT����M�u��k��`�;�\���E�@Ee�Ń`�1�s4v4�&<��t>��n�m	s�dzxf����$�v�2�b{�U� K(yiV!��m�U���z�o�)|ݫ��{I&u�ז��n�&]���f��"
�0��H-�_x�,�:�� ���Y�=� ��UŭW�JƆ�vQF��´���~G�\
֥�t�{yC2��K�n9����7�9I��D��� 쌠�r�2R\/֟�;J�Fm���=����n�/;���KM��лZd�M��v��ѡ֜�[X}%xdK�<|)��Pj
���ǝ�K(O�_
���8r߉����<fu�<zl��
�^ ����]A��m�z����}&ݱl5jU�#+�p��lL�qeO��i´�r3��4GTt�����{a��(��I�'����`��1x��M��O�<����X��Ӯ���i�-b���<�&��GƑ�u�|+��f�f|���aa�������aO*�����I��H��oC,��f9W�Ǘa�H��}A$W2��J�>�x��8�(�+-{m&5u%~���2����R쾒������-�<B����F�5G��
;@:���Y�~۫�<&��)�����dE�z���Z��QU���7���
�{��.�-���-,2�+��Q�%f���^\��)A�t�p� �N�Bp���v�`ݩz�uݦ���a �a�S�j�}Q*-e�Q�2\�ʆISݗ����������{4�1<�Òx(3�кr�K�A�i/z��ޯ��������V��
����G-�S.3�*�ؿql�y.Ȩ�r�ؗb������%��Sr�hY�w��ړL����v�����vS0k9�X�,�(��txE�r��M.WGo�$�iy��fe*�U1j��\%|�	��(;�i�6�lv^V�DL�x y�@�|6C]zx(����ԭ��F��]3��@y�-���8�|)Gnq���7Z�L#����Sw���x�(k������ޓ��(XaUqi���CǑc�"�z#�D��c�0TƵ�����N�z��h-v�X�g�[�x�0APs�!�B�/�����Z'�%v����m�e�+�kv��O@���k]�m��<K������Y��ழv�;�r���-��)����_\��\
�z$#U�I"B�<�`�}5�|w%�}0n�:��ӹ�7�vƌ%a�#���VR�������r�-����S�N�0
1�q�f̜��t诋��b���=��V��)����+���m�,�x��l��i��o���;�̯��Q=���vG�y�s\�mu[	I|mgj���{zk�LmZ��
�Ȏ���I�9��������)V��ފ��[j����QU��1�����&�g�H��b� ��
��̺�ݖ��#��#�J���t�Fh�ӿa��'=�������d@�.x���e<���>X��Z�;#b�8�B��Ḃe$�t܎#Y�1�Uݒrf�Xv���q�=��\��ett/��J�d{}v�4�ܷ�%-y�R�n�k��A�\ۭ�K*��-�3����ؾ�]oD��t��sV��5k�m�ڗ�Ѓn�X��EF뫯��z�#���Me]�Gx6p�U�P�K���M���/������4���lv��}�F:QM�qK	B��5��\-�ìҩSh7u��h�G+d�xUڭC�wf��4����wQ$W0�[�*e�a���͛�����":�3w��撢���6!��Z�m'�e����{�\�t�Z�Ѱ1N�BdC�G�����U��
�����۬(�ꗸ�P�^P4��-؀�j��YM�8�6��v6A1��;ϖ���âb�~�����o��L*a�-��QT®��z��u�rۯ�k��}�0�����N�4#�����SQ]����N�U���詏\��aC�t���2l��c�^��!F�r��񲍂�2�v�Tk���7-n����M�؆���!��43��2�����.�oL�²���-���L��z��P���ɣ�o5��X�hǷo%p�u�c�+��-s�p���Z�>ot��ش���ܡ��z��e���Y�ؐ�j]q�Ƃ�dD�I���p�n�/�����`]X��gS���o%tP�r.�U��+����R���]r��8˼�����M�BkU����P!���F�04�̯�JM�\jQ��<�r�]*�ˣ"��*j��v���+�j�N�3���g*�1���h4#���l�|��Ð1L�U���U�̢
�}Q�O��D��U^ڼ"�muD�1����ӆ0h�;Q���C�*^>u��!Ώ�����u_q����R��J��\�Rw�K��0Ir���4���:�?N¯e��1S�oG&���QD�U��P��o�e�㾍'����̀�uF�R*���w^-��w6v\�FHze�ܱP��\S���5)���fp��yb8Φ)2��k���_oXl+βۢ+�V�[.eogm�v� ek�^���Q�[h���^�H�+ӎ'��k�8߲{�V(0u�颈��Z���i����-�8�Xt:l�d�WnJ��2���cD�lV��Z�[-�2���ZH}�9�4&�]B4�3�;ܸ3f�����_��Ї�F�*��Z��B�-*U�l��֐X)EQeH�m[PP�Zȱk*����@��E���*���R�[eI*�Im$Z���J1j�
�ąb��QIRV���Kl*�T%EX
$Y*�HVE�R(T���)V����E��V�EV�B�
 ����J�VAV%��E��V�kR�(Z�Q�eFҪ�,lU++
ŀ�@R�RJ��V���TV�""ūl�T�
��+D+-��b��Ҵ�KhJ �d(�PF�Z�ֶ�Yb�+Kkmej�E�dD��2�VXQ��,X��j
�d���(�Q`(WP �%�ɽ�e�\{#t�ǐ,�;��f��tN����e�]a'�V�n��H�Q��p!��_UC������m�V!�W��i��K�SF���Pe�v���q�HB����p�ۦ!�>�T�6������ק����i�{�r���</�ʻ�.����#�E��M�iD�[�o\��xwӅ��T�(������ي`��Q@��+�z6&g��S�L�����N�m)O���r�fi����}�`cx�W�*�I�]�#�2GP�<|��Y���h�������U6�R��MO�m��g��V�>[Yg�}4v*jK'd��C��fb�=�:>���CC'hO�[.���-�1���~=�L�3����38 ��,C*�7���g,�jn^�#�B��Q�hI�z�J��r�qBҩ�,rt5c�*����k�F���;C�{��j�1 �W���1 à�u��U�,N�K���?���|���^c�&�甪��9�����.8q5/�C��uB����v��6+�E�x����sj�N��nv�5��1)<i���h7,QU&c��Yg�$DhS���̪�F����X��ďġ-!DҬw�t��谣dL�9��T�@�f�E�ϳ3�+]3z�E�T�6�_L5a7CD�tc���y�fe�Z����Z�kk]�4iG�h�*tݩ�n�l�`��?�����Z}s(�6.1��O���[�	=Sa�;�7�����ӪuﳗU���m֢�wDI_k����:ωߺXҪ��+.�u�>��y�5�{�Ӳ���4�]g���E��j�G�}�`y� ��d���\�;�kJ/�:���8\XG4�}qWXS(p�d>��,�شL��P�V��/�w������w"+I�D�]f��h�U���L���Io��ΰ�����P�~�gzo�%�NƘ���o�K���e�����Qh�>�/C�0&:%��%ᄹ�U�J���l�s�c�WJ��Ka˂�+�s2�ߋ�F`��PV�^���,�f!t�� F��B����iv�Z��� u��9���`�ju��U׸���]��v>>S�V��%��x�f��e[�7*��H<�jBF}����|�L:x�Xr7�Ł�K��o�u�,-J�K��jU�(s3"@'��N�<�e�����Q�PW����3����܌V-���f^��>0D_e�r�"<�`�	�]�9P]EB�/c��t��c&h�HJ�T�T��5$��I:ΏJpY�@]]˃)V��|X�m�|�uW	ܑ��Ѫ��Xa�|]w�}Y׽4�T�BV�]�Bb�樭�9X�Mb����ê댭�

��H@w5��G�,���]� [r��w�"T�s��pE^�W%�dY�w��<5��E�x@�T�`_; ��p|�5t�Y�鳆��̱�Co����e)r�
xx�i��7KNS�0�{&A�.e(2�#�<N	����w{��`!���BYZ2
���>*Hr,�N��ߜ���S���z���$�Kxo�z���9����c$_R�����k,_J�cL��=	�9�#|��^nN��i��<g��^��ղyX������*a�<;LÝ�u��,F@��ŋb������#��[~A�I`yV�Ve!p;d�*�:�E����YxWU�S�J���4
װ8�)�*���"ς�`��+֢���b`���i�Y2kOV�Wu��#^�fo
ӕ*�*�X�<5�L�������G��ma��xd��a7���o�[�g ��������]Bn_
��t��3+U{=|�v����qt�)7:��X����n>�=h?~�
����n��@j�&}n,�N[�u8[
����yN^�+H6�}�Y4^�٭���7���SN�zkz.N�vN�(�8hl��5o��Z�hg���V%� W�Cb�D�(1�8�݀��E���^���[�(N?)�c��u+�y;��T���d���ۂ�M�,S���]�ܣ}��E6a�\�|����b���6�O�=��	�.�"_R����
r��ǷN��DZZR냗��l�gk��>7*�4�躁
�,�[<�����o�v9�^^���&R��>�w;�C�}���G�g��Xr�6�� p� �f��i�\L�9ClOPh}��?^�<S��ʙ{޹(��?e�2!`8O�x@����GO�'~���JF���?�f��P�~ø�g�\(��:���P��+PeEf��g��s^�qF��K����c�#�ˣ�V����Þ�;�&�ؼ�eS=qP�j�U)s	���˅�ގV���{&�zv���l�ɕ}p5wo��wKWY�}L���X�~�&:�v�cR��2�&����}�1ૡ[<�&����.Z<��߆�xk�V���dz}�7��Y�fuF�^�T�h���=Ÿ@�s��u�v*�5=]W�+�/����Xui�2]~My)���Myy]5tL���c!A�RzLvG��_i�:�C֟����t���o�ͧ�l�y�)��Nz�ٗ�@�?{���t�Z�tF�|�[�vp6�vzr��+��k�ÀAy���5�b{�o��gV���%B4>w�'T�i�� ,�z)�-��6�L�M��d�_6�P+u��`��qS��Q4w�;W:r��_>�ݠ<oI�4�P�y�Y;�&�1@�Z�ʌ<�##+�!Ht����k�0�ĕmg���t=듛A᝗�Ԙ����2����\�^{%���x�T:4-�PY�!��{K�{�0�ݛ��A󴼱X�q�:�deW�h��v-$HV�y����.�X}%md�H�g�!�[2��hϴ�)�����x�RQ��V����]nR�S���`9mn����E�Ƒxj}(���w�����Z���A���t�U�K�3��ΐR}}qL���-9z�l��~��E��d^>��m�����B��qe"�E?�R���\�~w�֦8����7��s�j�[#ř�@�9�3^�W^�ٌ0p��!�CR@�}���W�,s�����)ʸ���f�}��3ϒ�9��'+��L��ˋO����[/d�O��v�A��X�*ڧ�A�s��l:9f��y\�Y�2��R���ξ�J-`Vȑ�u�����a��V�U�ɘ����?�jg�y�8��^c˧��v5�_�wQ��ҦTK)UpoJ�8"k�XHwX.�{lU�k��>�ۂb
^������X�4�e�<������o�V�K���Y�y���j�8����K��[����p��3LWz�f"�:SO��˿^�_��2I���Y���_<�f��� @�s��hI�zĉQ�rɁV6��es���7O��4_<�c�W��8���\�<b@0� �gA_Yp��<A�*O:��hѫ�)1Owa>�b��d,�.-����K�5ULH@�<�¬��Z��>����b7���dK�wבڤ�K�eUIpQ_I��d�Y������8]��dq��;1[��eW>Ȁ�!�rR��-��z�]�Uk���:
K�t�WK{;�s%vM� �K��[��p�zѳ�@�k>>U.Rc�v��Zdq�*�0�� W.�]j����Pk�É�.�86yQu��&0ˮXS*�FC�ք�]�D�F�8�cd���b�sDI��t�;��;yH=w�������;łP g�*5<`���wq���ê������0��p�95�+|�Ѻg��߫tZ|�3��%���@�zq.���F
���]m��0�U�NnfA��=>��z�zW�dP8�,�?)��^%+�Eo���[Q�XbVS��l<5Y�
�#@:��ε��t���U47��m[d�Xۼ5�R#�ßmA�^�W+x�əhU�B��34��\���S��8j^SA��vq���/GR�x ~t��S��7yu������9ؖ9y!����7�cl�RK�#�� \���)�h_�Н-85���ڑ�k3���ײXմQ�������;>�|(�ymHH�F��D�=9V���^������z��w;J"�r�3&K�<������6+��	���x;.���4��gl@F���/��zLX��쳭/��s<3�����"<�h�'�dʧ��AR��s�YwKvhuF>Ƿ�Uv\-jhl
�Y�n)⽑1�FaS�u����F��"<=j��;_{�[��瞿��_Ӓگw���5ަn��r��tYJE��1<��+mv��Z	%�%������0V��.�٫���<�s�e?T)�	�Q�i�|]��bFdv�dwb�{}'��wL���r�[j�EC3�83��J���P�:�z�X�уI�C�S�R�E�,Ϟ%O+|�0u	��/��ԕ1h�e��i�s�"
�s >�0B`�=0��� G�q_D��m�5Ҷ�Y.U.y��iq��|k�P���z�̬=¹i(n�U�z�����ݏ2��M�B�����N�J�׾��!}R���z�/D���B�Ǿ��'R�NEA���e�^ŷSyp)S�OM̽yv�m��9��R�5G {�b�W���4�9���.3�J��®��iY��-&��Q|2����de`t�2��/=���(Ǹ���vיf�l�MmO����3�t5�FB�<Jm�\���˗�@�׵H��<�M�'���N�I�Z�ueB%��z*�]��|*V�ӄ��zK���������F
T{�����!�t}��x�QZ0��]W!U�@V�be�T���t>�O\v2���ˌ�+]7��x��VZ�@�4$��J��e�\%2b�)l��N S��D��c��VVj�$�V�B5-V��^��Ft�8p��~��u��8,,2|��<5V�ٓ'v���"�LA�;;үY�.��*</�*'�0s>��5�''����~7 zWj���	���e���������.���(`���C�̺"2M��WZȖL������\��O��٦PX�ȫ��
����f���	���6N(�$��WE����*<:m㻂k��Y]�3|s���N]�^{�/�t���e�YW�^�an� o��u�g`(O.��+C]�X5ʆ�[�������o8I="u��bco�|T>�.Ӽ4�n�!{/2�g2f��}T��G��8e�	VwT�}CsηF�<�V�\��c�'�P�m�Y�Ӌ'm�9כN��4=���_�n�k*���h�����YʋФ�;�|o�0��nY}0�U�]	S-�J�K�h�Z��}Un�E�A�ךB��S���aog�^MT����J!>�i�3���g��R�T�]G����ӎ7v�~
yx�uL��)9��-��^�m�f���K�s�W�p��&Ynz�켊�;zkީ�&��]�S/O�!~��q9Z�*)��B�<w��nj���|��x��eb��s���'9|$�+]���&O����j�+d=C�5G1��oa�}P�����)v�ۛ�%��h�z֣Z>v��+�\|8n�HC�ŢIv+�^j0i����}�x��A�{k���r����5gE$X�J2���t<48K�q1/Uߣ��p�Ij.�Bz�+z6��3�]�q݂��dRؚd�����B+��'n��i���Ը����9+0C�}V�����=:ߏ)�Ɯ�8C�h��,g�Z+x��xZ>��ݚ�v��v|��_IO6���n�Z�S���Wu2J$�U�܂�Fjl�ݩ.봨xT�i�i[��Cw�ċ��T�����9���Q�p�����-��.r�ӆ��ƅ���	{\yJ�Hw�8[��;B�Wa
��s�c�kdNNpۻ�܎M@B� ��&�)�Y�w�>���!bFu��1B�r%Ex�� 7l��z��7��L��a�"���6Pc!�}��*��bA��^�P���vIx���mE���m߁�FҪ�d�bmcH2���9�PxI��������ڝ<�6��"��m�+Y� S���u���][e�bƘ��x��m53�/F�WkUf6�I�����Be�[�9 s��hI�z�J��r�q^��x�����{ۄ;7��X���PX���tu	
�1E��m ��΂��yeRT��Ī�x(�T�}��5;���<T�2�N^COФ����VUK�6+��H��v^,k�^w<��K��휥ǹ�;�^���	�Oed0Qߤ�t3�,�Ւ"4*��І(qe�m�x���\{�:w��1�nzT0.��xl������^��^n�A��t��`�N�h��Sۚ/z��8�K�->���4�*�>Lpv|����d{��DU�`}T=Z��0_���f�5>]�m���e��T�1�ĉ�&��(�v��(k�ƞ(�W�js�-�D�KJe���b��	���`�Kh�3��8�]g��2��RL��p�<�ڒ[סbYj��}�dRua�/F4Ѥ�{�z��;�隃Vf�Ʃ]�ƌ>4f�Q��! 0��&_�	r�dUʍ�X��	����,=��eՈMz�r	h�ww%f�S�0�;��*V&�]6嚰QѵcD�2ly��r�`Q\�����:�k�r�s5�ą?�6w K�lY�AB��)�!h����w��K��hh�ر�7�]=�c�?JJs�Έ��Q�\�cWw��]9p"��n�e���s)�r�]S�lh
�q�C��р�Z���,��PO�X1��-':�T���7
]�ȌteӑNlE�nЄrۆ��b�X؄wG�.�M���T�`���%��ǉ�݈^/\}O{+���D�;O��-�ݠ�&�F�j�d�`m��1z�3�m=��'����f��8�	`u�<�V��:�r��YÆ�S'�u����L���ي�pBTC
��5+1����4;�]'�m3yN>��ͤ�IW��·lS-]�\T�:u.�vrX���_H���F$�[��_��7�ٙK���/��L�d�.Ŷn������*�ɡ��Q�
���ն7s-�4���*�6d�%�-[�/Fm
(R!��2޽��>��4�*QygZ�ep�{�^�
b,�H���T{y�V+��'����V{"7��8�����]֚Η�u���PhgT�޸q8�)CCҳP��J�l�S/������o��njʭ�0�|^�����=d�gt���@_o�P� crĝLĕY��Z�{��oS�Qƨ��9T����ԍ���8".�'��]N�����7�ӶM�΀�ा���_�O��z�v�o�6�o�vm��lʺ�e�Nj��QĩiB�Qfh�U�tBb�[Dl�yÊh�TT);�M��3��;�<��Ɖ��M�5��u�����Y,����ކ��I���
tA ��x�f���6)TiQj��>��:�G/u\��6ݪf��U;-1�nd��Ҳ�,�s��23�AQ�h�h�Y癷uQa� 1Vl���i�9���9�Y���Ё��x�y$�R�1+�4*�D`�P�e'Qt���Bd
��xEl/6�7�Gcu["6��k�����T,�jj��dC2����t+(�K>n�Wj�M�a���aY�I�eԛ|c��Z�yN����r�<��J������܏*8!�Q3�9m����P/��[�(E��ҵ@L�ݾPwҐ�E�񜞇󓶳�AXK��;u>�ao �N���7�Ug{�ǋN���Kx�t�Noj��gGV�Q\8����Gh�e,��uċ��A�DU�0�.ׯ;/3{�YJNU�5��Q�Ԕ�-}�b��5B��AE"�kPUm�,�TP
�b��cl�h�*IF,R(��e@R��#ZIRV�k(����J��E�@��K[	m��$�AH�1H�b�Pm�%j
�#D����U�dD�RҥdX,�aTb+b�+Y-e`,UR�H�)YZ�"(�-���Z���*�,PPQB������**EPUZ��*,Pkb��Z*
E���
�@�H[BT
�R(,cR�Z«
�QAER����6�Qb�F1IZ«Td�m��X�*�*
 �+VE�֤X�#Z�E�b��Q*��F(���Ȗ�eB�am
�*[�X�Ԣŀ�Ub¡P��aD+D�%JT����q��f\�
�AX�T���V�@FEAj%-X�-1*,U�,���oϷ����~�ߋ�- ��������[����A�z�"�Ӟ�1�X^
�vTM)��v�|��Y����^�d���o�|�ܰ~�o�[;���r��gg�긫��)�C��!�o�`�����RV�];$�c����gꏸ�?y����ܴn�uc2�:�+�y�p�Oճmf�Q�f�Ǽǝ���%;���q12���E8_�����E�t�h���h2v̫�*w���`�+�i���2m]Z�t�,�Ö�8K�A�zo1^��S��z��zoN�̽)���"�<>;.�\r���T��]W �BPme�_�Bt��^�8�ق(N�͏��U���YD�9�U-Lz|����al�l��bC�~{&��W-s����s]8��J�\qd�5r���R�!�\.�d�N�2��yJ�,g��s���3�P�������:n"X	�s8&sX1с����V9ݚ�Vвy�h�5}e�~��Ч�oݶL�I��	U�Z/����{�46�f\`x�x�&0D@�f��db�>B��c�0�'nWM�f��D5r���t3���;����a9vz�[��V+��`]̞��F��R���AQ%V���&w0��V[�.�/p�͇��w+Oʰ
����ŕ%�/*0Axn��Zİ���H�}�/Odr�d��~���QU�����n��g�;x��<�T�����|�櫭:�ތ�!Yjn]����T���tO9�p=#d�|���X���^��j�GG�s�N���,#������r�-Qgsѱef�2�>����¬�5�=���d�A��t=��-�����lZ�c;ꟾ�G��'m����*+�G�]R��yt�pa[\.���;�DHmk,�pזy��(i�9�w���� -��:��a�ͥ�Z�R�W�z�&FK#3wҎ,��; �׺|��jP!�h����=,
ڪ���;kpD8ֲ�2��Ͻ�6t%ޮr�k�o�ߡ�F���GW��ǁ˂P��bd�����
���<�w�/��*w�p��>�����83%���d�nz�A2S�ˎ%��w�e�m����3�K���D�y+�pYJz�����s����D���	�ؙn,��'��H\��g�7z�	�]�a~��6��5�Q1�YS�x\�+��L^!-�x���B�`�Y����Wz7y��9cX�)�ĽS�g!Ɩ����W����U�����8q1�qN���e�~SC�G�g
�T��K��Cpl�B��Z�/��Rm�	��\��+�y��c�����|(�*�%�����A���� �UҔŃ|�֑U'1�n��㬶\b.,��kxfM9:�{8(��t�͞ K�
�v�F0��#o�t3�9M=�i��fkD9Sʴ@����2���D08�
}D��}-�r�|�������hw�դʭ8��ـA=�R2��~�*�y�~�K	�+Y͋��՜�%r}�b�R�PU��dQށp�ë�Vqp�,룧��P����}f��to�>�3�t}gw�	�Y*�g.�k��Txt�ϝ�]�^\2��s�����W2�EWh7��c�^r�3R�귔�ev#B��If����������5�j�|=VF]������yhε�xl^��l�]j.�<�)}2��VI�Y�i.�-ixnZ�k��Gb��x�$�C�{=���2=*����P�d��#>�Pj��b�O �����Y|u]�����L����)��MFa��Ǜ���t�%}瑛Xt6AoIΈE*�0�U[bz렬�L����o�-a����/�"�u�F�e֒��TU=�(`�,i��hU��N���9 ��3�"/�	<�ӷ��"22Z`�����p�r���%=�1C/�-v�zs��=<n�<��<C��X��%:-S��n�Y�7��޼�B�6��"2qq��x��'�n�Ŕ%ŋ;'���JZ�����o�k����V����2�r��7G���枌� 	��q�0b	tR�����N�E�{�����������^1לS3^GՕ�d��h�Z�k��Һ\�z\|8m`���~��^�\Nn���6��7m�P�_����i�/���ܴf�%C�gE%�b�m(��:�C*�t8JyX۩����vޜ��鬊~����T�oU5�L�ݛ�-��Ll��#�!��U�O�+�m�lǱ���BT�|!�T�V���.*�Ͻ9=-O(4���x_N٘.����oA䵺F���F縉���@�(��)�Y���P�:�_3Oe]{�f0ë�2��ז�N_�%����T��I��+�\z�~d3O��bSϱ���̯:U¹����,[åN�z�f2�g�#�Q�#��×E����[T�k���ЃD��rQ�c�����"�{<^L�E}�����œ��a�][&mcLV�ռ=1d]mΔ}�L��,�<^�����d���h���TR�s��jO#�"Tu�K��o z#V�=~w�[=�^�r�������xT������ V}�΂��y]���;�1yvAu�3R�Os9REW\�����j���[Fs"�;��k����W�@�X�����Ɩ</��r�A7��ne-�=���<p�=Ż��N.1��Kc�}Q�,}���߉�Zk %���۫� �8&���V�䮜�$���7N���i��{^Cl��;('6�X�R�n&���!��w�~���[��8�ܰ1�|ϟ���W��|;U�ȱ�Z�Ou�S�D���&c��Yg�$Dh�����h�<��c�;�x�D��>/���1�}r�K�P�l����;�u1 �#�L8:/�(��	�sQz�S�7��]�KncM�߄�FϦ�/3ʥ��T�z������ә��Ks&�z�i����
q[�=��۩7�����Ne\U�aL�5�y���δ"6��7k<�G���8\(hǱ�7Un�΍���X%V^ZW�%/:�e�ް8��f�x���R�R[C>l2�q1����A���֠��(�n�T�z7A��p�����,[�����b�~=YY��!�}0�%@L��;�y�ӂ.�*>5����u�F/X���˔�sLF=��,�����Ė��?0�������r��B��j`q='/��n	�Z�_�Ε����씩��\/*ʸ2�`�9����<҉]�H��S�dJ1�N$|���9�%����KѡDl��J�bo1-��U�e�����`n�<�o=���PK��q�˃���$�9T�)�Ӭ86)�f�[�5Q7������k8(�b�8��J
_v�����ba��B ސ7���h}��v�\�gvdU�p{Ήt��:e
Dw)�z��a����$�v��7��+h�\��J���{p�EE'$=7G�{������myN*��Q��*c��2 �E�G,�J���o��q7z���,�ċ�i�{N5hsC`Po�e�y㧆���E�vb �9� � {��I^�q�:���q!���;�C;<��H�FEiʧ.a��L�E���^�Z��Z~]�rG�"S�,�wºʡLm�
��������B�,�N��ߜ���C�؃�lڼ��t<vQ�Ƈ_�� 9Ʌ���@�Tv j1�`v�q��w*$ӆ�R�\π���Q��ٛ���w�$�z�����ĩ�Y%���<U\�ۺcQ^�cô�9J��q�bi~���l��N�o< ��6��s��Td<죄+�;��H��[!��V	�����}6�Xd���pp:�P#~{���s���ʠ����^)��ѣ�S[�2��{���4Ә�Qys�P�[CY���K]"^��.4`�c�8VYT��n$s�Њ��P9V���j�*�K��ή�v���Y��fhg)K���v�vAźق���ͨ��G6)��I�5�n-i��x�p�i͌R��W:ʕ	�ό8���4�{*ȥ��5W�^���6��Q�W
�GDI)F��p�����9��Z�;֮�;�>�S��h�`Lؔ����8�+�ѝ~۪�����'x_����͖�RV:K�c@Z�� �[�j�7�n�\	�;9�Y�&4�i~Ds+M7#:n��+E[*ϑ����Ժ��FW�\����C��L�N�xէ6��貗P��>��*���t��Z�7[1)C�^�`��/;T��&�w!j������>�"��Z ��cgk�^��G�a�H=�(����U}����s��b�f|�*�q�'BOz  ���ʘ�m]{Ըt�\C��0�w�KٖF���o�G=$��7ttq!�N�
�c��?�1\\�C��u�Ӽj�;`�%5�2׊�|�q}r_���*���$�#&�Ը]4xt�d�<���E��3|J�d�Q��'��Z����yC��0���t3岝t���[ȍ%�p5�A��@;Z����`�wT��-]�y�E�+γ�Ǯ��~�
�`<�**5<�j���W�n�E�A�ךk�s�>��u0�S}-��-x6�Y��ۏ��e>�9k���N�S�cQ�3���%��+]ء�f�p�[f |������ўCȺ;=aK�r���C���rɇ8���E\+*�-"SqRq�0����9��8�� άF�� `�:C�X3s6�u�ޭ�)��V���9r��Q�a�Åa�L��|FT��a"���.�����Y|u%wZA�M�4t��s�7¥5�8�:)ws�'�FluB�� /���<�������m���7�uɫ�N���T,�ʹq^�Ul��"���q651@��%�ō=��^��yn�{��y�{�x{�A��o��/����T��ܭ��`Jzjb�-t�͑Jɡ�A�f�M]���(��v66�To�'dס�[N�r��q�C�����{�4���r��V!t�-幫�3]tNS\]�����οӤ�rΊH�^*�+��t�w���L�:t���K]t;��n5Ai窚��r�*�`O�R8�5���1	�Y�M�oݮL��P�εm����U1�8��2�9=/rnA�,��X�O#�a�46���8�͎ͳ�b�����yN#���8	���r#5��]}a�.����T����'}/�Y�(pl�xK$V���Xc!�}���x��,B��c���񡲒aQ������i
\j.2��8\yrҵ�����Ȭ��ի�Z�mL�wʸ�[���zq
�É�.W��i��,���<3�����A_pʼ��
EG��ګ�4v�L��{�xd�N��A�ug�3U� ��v�we!�x�J�X���齎���z2���G`�[b[�.�V4�.����Nm��� ��.e���}j�uM�[yI������@��D����
�����badͧ��h+~T���}�E`������m�})��T<���3��T�xs�|d@�|�t�������ݼV��*�ʨs���Y9d��}R��st5c����70��#PnU����j���*�=�oD��2qkyk�;N�$hf�aVu�9�wL�����)=>�Ahug��SÆ��߳�&��>V����i�;~�g�M�J$��.
*L�C$��W盗�M���֣�GUto��Fϥj�C�a���ݤ�z���"J�I��{@��
L6��̎����x $��ι	��Z��48ӻLpUNס�u���Ul���e�Ә|�X�B]K�)�ߔڬ��v+	�H���pJ�(oð:�(��l]��~0J�پ���=����c�X{�h�\(hϞǄM�א~�E;4�o�>J��]aN��Y��k�MI��Ӻ�s ��Ю�Z��'�+��iG��+\{x4q
[�Sx���ߠ�9���䳪�-�S�%�%��:J:zAY9mj"ڳ���+J���#��K���ܚY���ս2��9kB����X﯒�k@냷��ϝ쵻�_Ff`��T<xfAC��+��IV�ã�A���wy��ѺW�㹄�l8�@;ܗy�b*s7��'	��k�W	Ex_L"͏J��)�8�y�Ӑ�q�(���D!�ӕr��BО�(�:.��)D�.���`�y؆	Ʀߖmi�u�A���ܜ�7��&$g�HV&Dq�t�F��o�ϗ��jBFVʺ�:�T\F���8��Y�����U>|�|+ܦ�k�m�4J'DP'Yv$��5�������3{�9���yz+'��Ons8==�<3����TD	�DH'�rZ�7
G�}qc4æ���6�i����{��OE<sՑ1�f S�/<�}sn�L9�7�C'��@���훡M�Q���%���S�j'�`�{<D(����ܣ]�:خ}���7�q���C�H�,�*�
�*�1��@���]}~����-EN���~�e+GB:q���<]O�T���\Nt����Y,oQC���C����H��}\�k5�R�0'���^�q�dv��Y�紀Xňn�e�<�q�-�Od��p���Gp3����t[}���05}�yd+Ο6�ķEao�p�t˘��ѹm�n�=m
֖���m�,�����*�0�)�Ҡ�E�v;L˜���w�~��QF�ps��\,㽋�?�g�nڄ���aWVE��u��AXM��ݗ{H�kfc���{�&���cu�wz��͛���VZ�ͺ���f��#A��W%�z��I�(���(�ʋ�����a�ب�$�Rb���^��A'9��T�f_�6�8�%�졼p�� ͂��Y�lǸ�U�ڲ���{��
�,\\��ʽo���Wu�+iG;'u�0��/��H�m��9K���b��v�r�1.I�����YbN6��e��������c�3]���z����϶N+����V��㝕�%5.]Ԟg%N}f�D��y���s-Y�ܼi9�+W}n�_Z.�b�2��`��=%�5�n&j��1�Ygmo^�2�^��9z�L��N��$@�c���O�N�B�'��5���jȏ�����U�1r��4�,��0E�%��b{+�����{v!8AT�y�=盬N2�U��H��V�ct(�ϭl�VFegwq���AeN�q%�2�to�"�1�܃:�u�����d�� �m�Q-�6��������I���K�J�,73:5��+1Lh'DT��R�o_q��&�՘
}Xt�d \1�j�:	�s��x����'nt;�􍍂J��g-�Ǣ��H�ޠs2S2�e�OK'����;�_b7CDo�Z{��B��F`��v���KN���ô{7P�� =���xi�.����^A38�#��-ri:�3��P��X]��ʵ�c��1����NctP�2#GEf�����Lq{ܹM���z-h��=���q�u�w�#�Rޛ�l����Q��w!@��wKU���m�P,�0��;M����o��K�&�\$ت�׺tmN�y�`�N>�Z�����|�Qظ-V�M���92.H�W��K�s����)]�K��-T#��P���u�	]6�R+q��t�o��
u��r3���oT���D|�>����PoGFK��pa��nC\��M�{���3���*Rm�k��Ow��1m�	��=��,0�A��2��J��*�GN��^�Bd���j���y𢡄���A�iE��d�f�" �V,��s냞,�w�f���!|̖`[�RfJ/i��m�0�R�d�D4VJ��J�@�S�c����vna,���M>�@z�k�X�
�o�c��ul������2��vJ41E�[���pJ�n�5C,��Wr-&{E�Z��ö� ކ)�Y��V5�d�A��L��\f�QB���1�K�����k3Z�w��ksj�l�$��Ѳ͵���P�)-���c-���X�� ��iS9e�����-h$P��ڱEF
�V*$�,�TU��U"�1E@F���XQj�X�X���X)r�b�U"�TҬX�,m(��q�ր���
%B��FЪ�al�Q��ZZ��"�6�%���(6�TX�F��F
5AdX�jV(�*(�+!R",DE����"�Y�.P*D`��$�.YSU��@�,E�c*XcD-)RXɌ����H(�j�(E ���Ċ&%b�R�j�(�!��mI��0P��Z(����b�-1�\�PF�A��@�bL�E"�QJ�)S`�Rb%d1��Ȣ�T�f%QjTF)���F)QJ�j���� �ѽ�R�Eɴ]�-�<x�������J���Ȕ���Y�m��m̸._R��b������S���gi�yŻ��������
K>+�u�'�mYk�E��u��mpť;+�uz���IPNk�����" ��s +��d	`����-T��>5�^�[~J��j��;Y۩�#�p״����ō��@��<#!�ZM��D	��,vFPM�c�{`ך��Nu8����Nu��D��Z�7��fP�T�&NM��v�\8;�ޣ��n����X�&r�=���2�'!���+Z=C��'���A���K��C��4��ؗ�B�m�~3윸w��W�ٲעV=\��{K�"_= b<&A3R�__���v�����{o�T!2��Co�tl�6�^��]�U�p��\$?;>�G<'o?���n��[d��@�S�!K[#=�K�8�C��M��#`��WI��Eu��(���E3=џZ񠄨ti>tX���DSʴA�������r?+>��</�_�#��9��wG�5��(�֟�zQ"��|�U4��Ӂ���f�甆T������a�~�9�,���k=��'ʟ۔8��إ�b�#�V����ҩW�P#��A:f�L��S�M;{/E���.�������uخ�hL��O6�sb��r�	A��<�GzI�.H�{[�h�I';C�W���B��{�34vN��]���un�[/"����	],�*4k�G��U�cӀ��V��v�!^��e@�.D*b��R���"�dS�$�L�'�ʆ�]*�p�j��y�k��/.�G���C�e�=�{5�淪�HJ|�^��Fh*�Di-r����j��N��BF�K�m&�{���p;�5�Gc5J; rn��tx�$H�Ī�|"Ġ�ə�J��ݺN�Ͻڝ���x6O+��!B��@��#*]A��ب�.�����1*���@�C������r�	�QͿw��wL�|�f�B�����������s���`��T��)�p�y,Uʊ�۫g5OY;�&���\�}V~�!��&�k>�F⋀�y�m56�5��|0V��a�ύ��9^�b�e��nV�b0%=��(`8s��l���-�<��o	�7{Ǉ����-b5ҏ��k��K�����%\x=��
��ED������XR����ls\��k%���4�*�:)_] �}�o��#�r.+"'+���A�1�\�\AK�6��'���k)J9}�1�X�Ncb��jl�<!��6\ˮ�v(��}RQ\9qA�! ��Na����q��]�[��\�n�{��
!��к���\�T �Y �jX��M���ԝg�T�5}lk&n&&}nf�F�鬚�}{����;�X�x�R8�I���]@�p�~�IlʎX��6�E��%B;!C.�;���Ǔ�ce_�B�˯Ct����K�85�+#I�:`� �#Y�Y8�2�w�'���N���&�ݑ�;��ejוt���LO�*�/B��x�]�	d��_&���C4�������ƥr�s�'z�ے��,.}ҕAJv]��<QvGR��.��(MFf	��O22ݵ^���e��Ȗ��l^y�r9e�Rq�����œ�Q�a�][V[&_����M����=y3��u��.�(`���ܺ�A�F�-��������ȁ ��k�y;7p����n��Y��cj��W8�_�^g�0b:8HW�(4Āch mk��գ7	o�=���>8	��0��/52V�J!��COФ�����Pi6�dٞ(-N`�'�������dX��VXد)9{7<��S�D�%�EI��K�CZ=�5Ql�r��Ғ���/�sEE���S�^!���=%k�x�<Nl�G�B��fn��o��{gc18F+�Ro;�?z7�[���䗷Bؾ�!h'f��nkŮ�@gl�d<�e��[��WWьwY���^
���/Ɲ�r���N��~��#�띑�+c~��Fϧڀ��/�1�X��q}Ή-�et,;j���=���i��W����<-������˴�Ϯ� r��|�TjJK~�Sne��.�n�){������;�
�3y�S� 5��kB�\�{j]��u�[Z)�~_=��vl���7y5�]l+|j6�Fd��ڞ��vu��M1��o���yӺoҳa��N��0n��b�k�)C(p�een&&[S�}A���֠���-�<'���>���=�/}v�	�'�K����J�Ү��:�0�NnfA�=ҽ�	:ABz��K}�����OJ�Y>P8ۈ���RKG��=�����U��p�����M	n���d��|k��XX�$g�HD����<'��]���D�Ϫڐ��gk�ŷ�FlfQI<��F��T_�ɇ^X�2)��ia�4J'DQ:˿I��3s��5��k��jX�K�\Y�*�.�\���Sۜ�	��f���#B�JW/z}=�OJ#V���oz�:����I�1p�9ڦg�P�^����*���j��%�[��s XK3�O?=N���ӮU��7 l+[Ǌ�O��خ�ˍ�|s��F;4����ق=���Y���Ġ�A�w�ѷo����D�������mQD���4��uu�X�0e4���5A�jZ�'<�%�9>Ș̣0��!�u�U�F�������h�'����V���Ӈ8
�G%� �8f�O�ek���ԓ���D��eЉ���]�{��e(3�
�y%�\+Qt+�O\�j�7㡍�"ɔ�9��ч��/\mï<��x0�����.5ܒdraa�K��j�TP�3;P�����I��v�I��­$�ӱ��ꐋ9�"����T�Y�D�!��%�FnU\��mX�1y��^�p���+��yP+��dU � _t�<Ѻ��p��>�)��8�7Ҳ_+�{�][�MgU�"���9eg�\t��1KZ�<�B`Oe�5�k���d�9��~�$�-��kx����X����Z�4c���eObd��Lw�S�{mo�\}�7��8{�_\����xd�/&�n\Z�#��1{T7�N�mzw'��x{�;����ʏT�k.f�XUf�\M�3�K�9 ���Dբ u�n������TP������ڰ�6S8|��Qّl�����hf��;!2gNs[ڠlQ�ʜ^p��ŷdc������jf�F�����A�,�ﵙ@�4��#gR��+ܼN�JIX�b��n,�t��-
�.�H�_B%��ZQ�b��B�|�T��8{���*���X���m�O�s�]T]@���]ׅ�������W^XH�T�}	��PPs�>�����%�0ԝ"2P���Y�}��QՕ����u%*��,<+�:�&�v'��@��u���~V}!��5ۂG��S~r�N�B|O
�$SeU&�q�=Zp17�l�P9X�tw�[����pc�a�n�՚��.f>��� Mvx�@��5�0_;<���r�+���bV��{�6�[�m�)��9eخ~��W����>��r��،�W�p�j��yN�	���8BT���#�Ü�	�Ƕ;���.Ș�r�BB�tDOr#I<|9�S~����^i������u���2��FÕ(�I��!������ćA]D�Q<MzT�D�ׅ_p�Y�*���$չ�r^q��g��v"$(@�L��|FUK�5�!^�
��g<���R��t���y�E�9�j�	YV�y���ܬ�6:�ޓ�/��^W�C]��o����!j�&�s$��c�a���}��U����E���\�:�f5 ��r�@�ٲ�#��2w3�9q��u�w�J4����'��R!�.�,e.X��v.Odw�CU�+�"'Lit�guZ
}a[�ǭ�>ܾ{�0p�{�C֚>x�*4]��sT��c���u1 �Z��`{5��g��
sa���>ʓ ЫsS�=B����l�ʘ߇���C�Jz�v/���Ή�yӯX�"F0�> ����/n����Mc�\~����&{4[!x*��"^ԣ�F�Rf{1���-K�^��Q�S\]��}����5��m���Q��K�.0�gsWF��`sQ�/�v'jT>��n�-"ުk�@�.;�VY��[�������:�wV��߹�\j|r�4$1 Ύ�#8���ץS����&�x�Lm���c^�ɒR�]d��5�o���]�<A��W\�3	U�bs� �|�*��������6ݵӯv{�][\�~�=~£�x�	U��J�W+��9A��i�D%�Ia�`����y�-�:g�8�n�yҮ��]�#�QvGR��.�)�Q�m�ۖ�'kF���\��{-~��|��?hɗ���4�[,
��6h-<NPgW��p�|�*s��l�`w�sd�ºj��b�v/_#�Q�)�r��?�v�~B���+c/���FU{U������%�I"�0'�Cv���lꙶ��ug�7[}r�+Ɔl��I�]Ўvy%�']:J�]���; �sJ��	kr�]
O�A����k7_9ڰ��{eӲ_������2��ppR%�L�F�NT�(�t�����ez�{�zG�d����,�-*�"�9:�����F�!�#�Pn\��+�vE��y��x���'��f3����a}�gM��V6i�����<�MG	V0VZ1!�vޝ�����p�DWa!��:(�����Y��,ݎ�`�A�p��<�q��
q�q��>�	NY���#�$�:��>��
�P����Ϥ�^*�.2���+;:qs�!M�o4H/�*t�^3����*�������i�yT��"{!�;6е~[۽��lI�X��]h��� �� T�����}���p��&�v͠N�)���ݩ�4���iT+�[9^���_�)��+���7~�����7�(��7�$6�KҧM��%ߴ�U�+AW��I��6Y�n&!w���zs�A[�+΋>�K�݇��x.��]����t��:ΰ�9lS�U��J�vNF�%0����9��BBoӽq���W����t�CΦ;j�j�8P�H�NQ��(��젆$�B0�CY�͍��"�}���V���n���e�7u�8��g���J ��˰8�;�9���UCcp��7Gef�]��۷���V4�����*
҅��M�O��I�%(���u\ *ΰa���VP�ۋ�� u���Ӭ�σ���F���ʸ�l�'8ϖ�:"�t��T��{<pھ�μ�6�ѧ��Hj�ئ��r3X��ma�����tEx�e���8J�c�t5�n�NE1S�X1��.
�U�'�s8�<��*w���iU�[���=NgGy�(s�?��"BT.���*^/iƦdd�̸ǎ��[��a�Q1R6�oI��~� xI���� �\#WN�K����Kl��J/�4�QUp��&v��YX⿵@���,2�ۥ�ɐ`�k)�zE��%�\+Qb�b���bժ�ǡF���,vr�����5�0�Pض�(谝��.7�ܒds��墓�.����HV�}myÙ�Nnƛ�JI,z.s(F�9����<J�WyX]Fx�xf�g����,O��Z�����q�D;D�;E����E��
�Al �XT��L��W/��mvM��R���VƔy�.92�"��ɩ}�|�.^�}+|��O���ͩ�L]a�Ӏ�Bj�̘N&mL�f6���m����+K�H��1V����s�@u�l��h�fH������D�߫���]������}��J#�8�'x�ofN�VI�4��"Q�9e�q�xj� �-jȞ6;	��`W_GbٗC�^s{3�yb�**Dw��j�Y����<�)}��(`����E�ȯ��=9���SY�\Ӧ�L=M���*���}�C�g�鞻��%�'k%���d���OR��gk�ؼ�]7}ݮ֛u��lBW��A�rv�aY��c��˖�s���e�^�X�D�W����� �_C�%:��Bt��	��Cnn��0R��gҗ=w�7c6VG�	{�Ή�D!�%�1��e@~)텑Җ�l�=�1��#ƕ�'@��#�Ⱥ����1&C��R��B'@�%�����tP�qe>���s�ߚʘB�7A��F�}�"J�L=�h[�|��w��\ʪQ*�x��Ӂ����`OsT�L��XN�/��?	������hr��Xa� 8N����5���i��<���0�1Gꢸ�]�fVƘ;ۏQ�Yp�u��uZ�}�Dп�}p��Z?'��p��~~߹�B���IO�IO��$����$��IO�BH@��	!I��$��BH@��	!I�rB��HIN�$����$�!$ I?����$���H@��B���$�Ԅ��$��$�	'�$�	'�����)���9 ۸��),�������_���0R�����B�����$����4[cRX�P@�m%�j�iLڋ!�K#5fQ0��d��J��4[�lvgwU�bm� �b�wU+)vh����%.�J��J��n���2�ۺ�KAQR� �  ���f�%�5�`�Z�"��M�6�Fl�,eZm�56;��ӕ%"�뺮�W]:��7v�t�ܻ�u��t5�J�"�V�w[�ۥn�]����l5�ER�p���Ӌs�MW6�n��7w9Zu��]��e��C��m�kkbֶٳT��li	[\���Q��lm�5�K-���T�Ħ�Zjͦ���BRJMl�      @ DS�mIJ�� �     S�IJ�       �101��&EO�A%J�bi���d�@`)���R��i��   4   �Q�i2d4�`S4��z�2=OSaOOR~o��_g���L'ݿ�BH !�J!A�B���!* @'�@���'��%�����IY�ӯП��?���X��ޏ������0���PH�B K>A�_������2�Cp�d"�42I x�~���s��&�GSJ�d�~:�^��3��5����Xj�  @ `\�%��` 4Qf���d�,K��d�,V�[�2d� �  n�%m�J����%MXI2�`ZBIĐ�� N2I!&8�Bq�	�BI�(H� �$�BL�I&�m���f��p2X.��`\%��p2X  X0/�� �5h ���n|��`(���3�c��������F��(3��>Z2V�"E�����������y�y��Ѭ{��eK-?kǦ���b��4�����(.���a`��x1V��8X9Y� �*���I�`/a�4� "�^k��˹��I5��E7&��5�[6���z���S24�kKNn٭�o�!�5g�i�ۗ	��#I�x�F�8�ӛFn��į��C(2�3.Q'I�(\D@V��G!�[,(h�c�0�*�+4��r�FSR�+z2k�u��l��o�.�$6Y������t�[�ǆ�WskIUc���wf-��v�MюVH�����C�]�e�xֺy����5�jl���J�d JMRR(�cpC�lE�g[ܺ�-�{���N�g\��$[��$Ztr)ovb�Qi�FX�j�N��PAO*m���˥ji�LB��F�a�C&�H̠�E����u
F��V��F�U�5�����{�U�E�����;��/1R(����L۳m���U{
®䥇a�v��9Nhg�4V`�$�\�!��G�c��3h���Z�2MT��.���4�.ȕ
�x�Mct$��He�D��X۹*eVM�J��F�u�4M6�G��=YBl�-[R.�� G��.��qp��Nɲ�[sIs����MX��ĚHvi�̒hsj��mÔ�E�{����̶�v�٭���U#���h�2��a�j��r�L6
�be�8�o^X52+�0�h�W�m�:��X�%_�*�fMq1EJ op�j�V�eֵ8nd"���w�b��Wi�c��V7�Aj�c�zl� a��+ZS �2]�����غ���b�#j���:�YY�4��6A�%=U���I�s$��P�i����x(��u��ݔ7���M(U������b�0��ˑ
ݔ��Q����p�n���%�@[yDd͖��o5��t��2���޲�V�j\�+�*-rS�T)�O2�b4��W�ܺYH`��S4��˺y�r�W���#dՎ�n:��l�ͩ1�E�HŔ��D!x��ŭ���S�jXNm�K&#Y�UiJ²�=�	k"���6]L���a���]Er�1I,?���̫̼�T)�XVZ�h�[r��)�F*�diF�m+�:	f�8�J��*��m��kB���X"1�4�j
���ۙ*5�SqY˽U��_����z�ևE�0��<uy1㺐��ِM�#J��F��E�Ud\���7�A	�uz�+��<n���R��)
�lt�6��bD�2xi4en�*V#*VӀZYG/N��:���d-8�J�:��t�c)�RF�`j�uh�$��N��M�*�:���[f8I)� ���z��E1bFj�e�7c'a���t`3%��剘[����\�ŁC5��2���j�u"5ҫ{ɨPU++t���EVeh{0��๘s3����9-f�--�14iL����hw%
/**6�b{�mֵy)U�Q���a�W��s?5��*��R�	�.���x�#XkYO`�WE,:褃T�l� �*u�ˤ(Q�9��q�H�sVB�ށ��R�$ck���pg���U+���P��&&�a���{V��$F�RIV��Tc]���R��[�%^2��BCJ��!��B6���f�T��]��G��L�YH�Ci��4�D�����������
��t�SI�?�T�A�&��4�.�Pd�SN�`M��Y"a4�Ѷ�����,Ա �uaJ���H�P��b���`�0�@���'A�c�D 5�j�e)L�T�"�KX�k����g��>����?sO���y�G`�.}�o�������R�iG
���r�w��խ�-�,�*U�*q`U�����Q�w���
��KZ(�+b��l� �Jh�HH����b�a�v���
��U��C������jZ����ōoXѴe�u�S�|� ��zܸ��}Se]�H���S:9�1gl��\�'A��C;M.Ǘӹ�;���Dڭu�Y�nN��
���������{�+:9���s��f���m�[�ד|V��7t�D�"u-��&f,���CV�`�c$ �k���L�r���s��;��К{�Lw�{�.�c�ɖFN��ع*��}K�e[=���V�a����r���qQ��}��Թ��w5�
�)��;���øO&F�!�y��j]+�L����9|r��c��,8{;�8�ˆ�@y*ؗV���痎#Yc,�Wc3b��_���k���;WN��/On<F �Нt�q��\8�5
"��尐�4�֫��
!+�B[�KR	�VX��� ".=t+5�@8ir�q��F��y����2{��m����}ru7�q)A�w�+js`���T�^�Gfr;G.���[�����6�&\��)#MN�;)s-}��ﱒ�Ul��H
v,�(��s8^�㘞� �NLj�*Iw)��v��̣l*3u�m�.rB�[�Qlኦ�S1�6�a�=Z��9I��^�|��Φ9fSԈ�])Rpc���ֻ.����o7��av�S��y�a�NB��&1�΁������R�6��(U��0���GHvF�ϯw27�e��5�2WS��б�F>za�Y�.Ҟ4r.�b�E��x��3x{3b}�����ϖ��\�2,ם݌���t�>�)!\�3�,͔pȇ��`�WTqp�7e\�Op鼆R��$2Y\����4J-yut��Tn�M�4\jtJSK꺂&�o6x��6�X4����^|�yi{�!ӫz([L����t�WX��R�F98gpJU܆���C����s���K0Y���o�Ɏ�:8�c&�x��s5(�{���ٴ����r��.�_���B��q��4ܲ/�b��-3�*w2��H��}V�9q��b'�9x�h�C�(S�)3���}ꗌ��Lc�mJ�e�"���3m����ɷ�e�<uZ��4��/��������{��	۸�$�/�v!g�惶��plV�f8�k�Kq��y�Lf��8�W���Z5q��R�����)t�ܫ�V�5�@�۽I�PFn9�:���l��vi[&���6tn���6��ƺV�.��~᢮_N��k�5me5�;q���o�rl&D!W��Wv�&���ԭ�0��t��fp�u�>P��M [�+a��L�҂/�2k�!Nz��>ZN�������.fu�z�����x>㺓]8�⓺{Hi�����R�!���E�l���d�6ud�2�p͉J+E��� ���{B�ES�7�E`{�b�p`^NI^�z�\��N:]y"��f�mF{d�j���F�"�Sj��=������ݙ�޸�!	x����UZ���Y��n�=[ߤ ���1�ܩ��.fL��ݗ�֬Pw���+�V���}N�h�������p�wI��ۆ~YW�����LL��i����5���������o/������LW�"|A���}�� @���~����I����▙��w2H@$�y�c+�~��~�U��/�����8+^�;�Me�M��ADu�?kd�bZ3�'��|CP��'wk$�u6��PM��"V���ְ˺9��E�-u�(�����z:g0&	�s���e[W<J�[�7��ڭ� Y��%�O�&O\�s#�*�a�S���u�a7�:�3���
o,�ޡ+z��]���.ؓ4���P�*'d����~5f$�0  �  �"   C� �^��ٗ���\ё�s0��Z��с�Nv.���M��x�f2�2%]n��6d�P��o�ҩ�
Տ��d�n�NР�R��ǯ�8J�S��[M�V�����V� ��]�󌊄�{�r���2��*8�5u1�ٰ���V�fmKu�;Gm<04M��-z�eKk���h�0   � D@  �  ;�:�<ś�_�ջ�6ɢ�[d�$u�u�K��x���ȏ�t�M��c�K9�P3��4�ǣG�<���f���K��0R��f<j>*�Z�eY��g0�IB�q����Z> �®��c��.c\R�~�PQsVd���M�f�*'��U��w 0WMw�z�*���'�[�wQ��o@@� �  ��� A� [�r����}�׻�1���� �+v��U�Z�W�f!i�!9Ywʐ�Ժ4�l�V�H�ɒ�ʻt�M���osH��j�E:��eٶ���ot�ih��&4W�&:� �9EœPß��5&��z,
1̚@����%�	�9�������͜  �p�C@ � 4Yq��E����L�M��^��t�|7	 xp#������0�߲:�Ӣ� ��6e�19�W��w�l^��YBBAkF�6m�3�n;-�7�i���HwQ�{�s]��g	��l�ْ*�����3�iM)Xqw%�nkw �ޥn�ZT��ra<�0���2��#�� ( �  fd ��
 ,����}YU�^6���Έ�e�3��-j���f�<�ŵn����^6M��Yf]Y3BBN�9��zڃp%�Dd��E�S
�Kb5����yɂ��\#��v��M�E�09��M�7g��-�`}G�!(Ї$։����~��y����xт @ L� X �P�ne[�QM���\�Y��J��%;���
B���p���o�)�s�a+k�з��૝)��5�VR��-{��J����֧9����TK�J�?H���W�4&��_4�Vl5т������@�=T�YN^j	  ��	�\ @ �$׽vۼy�Mq���^s�Y�q��Bh��`�<��6ھO��Ŋ�y�v��Y��9�L��s(�*$���L��&�mm5�9���dl儨�@x���0�C���W*Ln�ȭ�r��a����܋n�֣�ueYҹn����pȓۛ�o0iZ$�  Ѐ �
 �� B  4"c������1Lp>�r�3s��Uv��j�Xˣ\J릉o���s;)��{���+����*�B�nC�P�C�9�v���XP�ذӴ�x�9�b8r�Av�X�:�E|�7Mp�j�PĦ��suq�v���
#Õ�tuFl:�bK�ǚy*�G�wˍ����&s�ulX����^[�*N��O0��"���y%��(�M'
��uP�j��Q.��X�:��z���B��@���?�xSWs��v��	\��,�$� rw\�76�]�8�fi�d%� �U4\�թiK�9lV����RW�h��:�9Wͩ`t��q�y�f��W�cZ�_y��ߪO�HB �D��� #.�!��%-=��_	R��[��7�t�!�E�)�ES%6��BN���u!0��,)F�~ʿ߶�lw��`�<�Om�g+��5�V4��1t�¶1��ΐU��QLY�V� ����Lv:�$nr�?^w�i'�ęzx�V�3�:$Q�^���f�'#v�<�_���|�N����J��z-C����B¹�3��R��$5*�LX`��X���|�a������^���`=��	�SڀPD R5QiX�U^y���ꂪ�[E ��U�Zٝ("襪�ie��u{��.�EP$�"���BQK3%]�n�����*��.���l֦����Jjڽ�va4�5LTh��V"U��vUU ( !C𤊻� 3SM�.�j��(U������[_�	?٦�܎-!H�'z��N8��%=����j|�&!F���o�3y�[U~�9	(,���b粱Z��]:I�����ڬ�gG����(����j�l���Ջ�l1�f��13�����h����
k[���8׮or�>���ڕ5�V}Q̭}��X�����VuMNc�Q�	^����T��sMc�x�@Z�G�{lg*���1ʶ���d�)�;:�kx�h�X�`+r�{��d�(�]�Z7vXHxSc�`揎Œ��*4���T|�wXH���Ϟ;\�����t�!B�����c��W:o��}z�f�&��2V%��`-��H��q��ۅKʀ��pV᧋�ȓ���&�w����c����X��ٚ(a���>y~u��w�k:gu�e��n�o�j�g�N7�0�����0�Zm�0���|ֻ��{�6�e�M�ю�Lh+���^g;E�<u��&�LZa�[�r��~J��Ӈ@Wa�LX�J�_�vb^��>���6�'v猿X=�fu�����y�M�4�K$�@[�L�ü�����o�m��x���t�QH����v��Nf��g5�95��٦�ܴ��{��\֓�Q�ӄP�u-�f��vy[MUf�Bb��>3F�7v[׉�n��Sc0��7�+V����4��;y����dJ�ku�o��q��<F��(�L���x����[�Zj�V��㎱�ow a0�M3��c���;۞�g��~^�L*���`�.��."�0��2�x܍>�ܤ}����w�8�r��v��&_i�7��y2�:,�u�q�N�hy�W+��ו'Sn�O;MQE��Z�2l@�TyʝL;x�X���Mf�iI֑n���k|���b�i�=Cmg�w��TY�Zh�*���)1���ư��+7㚮&qR)I���W,�N�EuJ�,��XU�]sٶ�;�.��@CAe~���	
�}�w�k*c��a���G��<דk�l��$jm��Uq�n�ZMX�?�JF���f�?w]p�
�Kn�٤�W����̝���l-�Tj�Y�
�R%�ɈV��\)NUJ3	O6�֊|�{�=�ZxӆsU�k��+{V��¿U�x���B���d��S�ք<K�JǗ;�_��m�Ô2�<m�ݛn�噺7��4�Ag�Z��<K�S\��N��Lb�:�+��ͅZ�xU:g��.^�������j�XS�j7w%��xyv�C[�v�tz�xV۷���A�����D����オ������Y����u�¸d5��G�k2���6��LZ�{��<x��\�,�0�2�k^kK�~Q\��嗪6�E�UԪ��c��]�ާR���N��).��Yγ�{����Ri-���K޹[��WYm9EAp��Cs�1��y��2�o��6�P�;㎚l������[)��FS����m����s{,�����X��@�s�����)�L�V�b�yx4c�F�)^Q�z��fS�\5�k�oF�"s�g�Ӕ��[�s�{�ɼ��3nS������g?��6M1@U!���
�b���K���?���?�Y� $X��uݹZԡ�a��?�O�C��ϋ��d���Y{���iI�^g��3����Cn�B��ߧ@�>��^Z̝���x��	��J��%��jf��˽;k�{+p����O��vE�I��4���sK���p�j;f�sQ��.��D��ƹ��ҙL�)�n��e�0����1fZu��a���_�0��N��fS/ZfL��2�yvu����S�3Qr���m�ta����t�j��r�o�;���htE���Q���a�k<��kE&�3	i�+U�g�����o�.�;o>Qi
x�y|"�Nc��6�Y�ڷO�0D�yLY|�W��oM�阯�0<5(z?1L~���x��\AE�<?zxxU�_�"����Sh�e��q�^�a�+�)�h)���*u)�(�&���q{�E9C���<i8�����vyED�N��S67�9A�p燤��B�g�P�[-:�3YwY2ƷgS��.1R�O<��Rn�K���wlx{��]��j�.��-��Jgq���3G�7$�ZO�0=�����Th�k)�h�<�n���K6�?ϥ�W�fL��r���ф���\x5�f��w����܅�r^�TP��1t�����]� ��,��+i�9�q(T��>Z�M���Ӗ�ЁI�J�����Z�St8'ՠ�R\�S�vva���:�-�ĸ�CN��<����7Y��d`��L	0{�}C��t�-$�{����L��s����ss^��k���^�Ϧ�.a���J�*��ex*���ֶ3��y /�I� �1�.Ηy ���(Da�h���.9���zT�q�����An����5��
���A	2��=)��GB�'�fw3y��;����fS�Z�L쳁vY�O}_��X��
�B����F)ms�{�iڴ!l�(�]�P����لc�4���bY�� B�Mr�H�Q���Q��"�������(���ݵ��yʻ�Z�JR�ʺ������T�1�D���Wd
#���A)E(���ߛ{{�u�ݱM� `�´A�����sU0��k��0�>�7SX�k��_vt���ݺfSM*L�]�1�w9�g��ʱ��j�,URE����!��빮��]��N0ϗ�Vz�N&R�n����7^!�^��f�J�#��4��n�I���7ʦ��N�Hc�2�8�>��:1�G�k�4F��*�?�1�k|H�@��`�Zj�	Ʃ�+ �CR�/���?�x�l`��^�V+!U���y_����w�4(,K+v�l��8���%���b��@�fIf�7��M'x�%��TG�R�����:���0j�5R���n1�Fs^���2��m�i�L�)�3��)��]��6)ǭ{�@�!�h��V;$��ڨ+�����\�}B�VY�]���=v�f=��=��^+Hx��{Vi���y�}v��u��L%w7N��L�f��5F�Q��ۣ��o���CeiUKg^3��|�)}��׍'I�-1]�6��x�<��n���r�fW��nc͔�܆�	\��X+wwk�FǨ��so�ӊ��tJw�;�J��u���+��׎�g��.��}w��P��U�K�*��W���7^95P-�4���"�?��/}��}�u
�Ǉ�	��Y�@��U����Nb���YI�����2�Z{�q�`Yl�ta���f�.��UY��[�hA��Ɛ�U��pV����E2�ZgY~�y���,�2�8y�,��8�r�>����S��E���:mu[�����8|?���	Ѭ�S���[�w�~��y2�Z�k|�||�q=r����3��O��+.�	�[��m�cE~���^��N����+F��Sl/'�)-/u^9�מ{�9Mם����k��N@�Jm�n<�C�֝��/�������B���/��.�hт������Հ�)�"��� ]FtÎ�L�m�L�A���gG����dˀ�b�ߵ�c÷5��L������Y�+��I�9��<x���v��*�(�*?D`u��,�}�[��AY��{=~.������Y����M�����s�4���&�*a�L0Ç��󺾧MPpk4x�M����Re<<�2f�������l��X����˿}���=�x�v��4:L'�l�*�{��^cTͳ�W0~��K
�
�,����-?�5�T��\���5��P�֓�����ۄ�a�w/{�n���]i5���x�]G�^��_��TpS�UZ*���~��8�v�ާ��>Y�i�h��=�������__G��7SM��B�u�!��k�CpZề��{�W��k��v���]���,��Ѣ��l����5��?@��&��R�|/�c�]g�a���*�)���6���9�9��X05�m��^�u���)�z�5E�U��2�/�Ɯ2��N�qG_"��\xk�sFiǜ����eӶaw�u�R�e��x��r�Y�����'���PuEf��CW�9�<��^���<�w�T�w�F��ŉ�t�!��_�+��U2!��W�'}~#��'N��k�4G35`�u��o}?9���cΩ��������~�TE~V�}���=��/G�GXRbʊ/1^3n�<��Ǟ��~�\
�h��R�|XCGe�\�����p�q&��y�s���N��x��Y�\�`��a�fSz�}��GQCG�&�M�p��O]�8�M����k9�C�m1���T�K��<�R�F=��i��&�c58�s'|�G�m���t�y��fݗ^;�/���Q��h��s���w������&�F�I��'��Ek��;k��C����%�I^W��s�9͜f�r�1P�8v�'���Ny��7�l�:��WkO�&���ߺ�z|�����6����Q̟�5��)\8W
D�+�
<X�~�^��\0R���1��Kܪ�������0��x�R�z�5^���(˱�x�����M~!
ҕ���|?!�p}��Lh�Xш�������
��p��:'�5]k�T]|\�yY�i�;xvi~�7]�%����O��Ӿ�g�����x��7�_5GuA�U��s�+�+���F����B�(�����d���zZ^�_z�O���Io�׳�Z��j՞/,	����k�s.�s��n���0LWn�G��tOm��_�݋o�g�����d��:
�>�Z(����V�Dh̍��ut�����ؾ��y�#!�flIz��1��{�A��2��	�'ء�o�dS�s�O]g�p9����ՙ~��u����x][ϋp���v���B�?mn�j��[�V�xon���xr�M	yOԻ׊?���ԥ>��I�}�e�Rj�e~�U[���?���fu\rS��kU��m>�ff��P�K�>X�~��P̢�����O���s��$:E��Y��Y��Z1��k��t��I����k(����o7{:pł�ܙ�6g�V��A�j�H���O��Dm�SN0r�\�I��t��{�"��Q��ۘ�Q�\�����+jB�n���M�,�8��2�Ĥ��D0���,G-( �a�K �,ʁ0�"�%�)W��u4v"� ��/����a]�C��,�63����ۮ��,����밆�[������ ���Р������wYVN4����^�P���;R��絊��"�*��%�-8��f_Q������׸�J�#���3\�>nBy7s˩���^�R�[�T�����1�2Wu�#��'��E���ڡ���;�M���R�]R-���5��y�i�[imVE��{���(�J����*�j���)�ʪ����kZUY��m-����&�UA�QkZֳ�R�U@�UJ�eUE����k&�STŦ�Pb��T���E�E()IQTR�07�.�c�)�V0�\'|�M��B�o�h�-�����i����0���^��������1zk~��C��a,����@���y�L�4�
�I�� Nb��@�!Ԓi	8�M0RJֻ}̐���$4�<fRC�q xÌ��4�6�V��q��q 6���ʶ@�<Iꡔ�TwW��%$�P6� �Jf�	� �CL!�y�k^{����Hd:�P2QT
HJa�~�gum�8�!8���mw�3(q��(�<d��a�4��9��8�<@-��2�ж�wT�Hy�g�fN�7��w?z��\�glQlM;>L�.�2"��Qw=�8Z�T�����`�Yi$�ۨOa2�ĦהHQ��ɆH�;w	� zɦHz��e ��RCY��]T��ǞsX�\�:�Kd�$�2zɦ�RC�!�7\�d�<�![�B��I�	i$�M�ORC,���1�w��0��D��!� J`�Il$�$)����+RC� �I2B�+�!Ą2�,	haRJ5~�\w�y�%�	���d���B�Ri�XI�Ik�s��a���B � ���!ԁLS�x�5�	�!�续{��$��� �,o���������w�x��k�y
G{�~�5�o{U���dB�9�+����]�)ު��=���D/��(N�jM|v����ى�^�\{�Ǉc��q���u��P܅�n�������s�Y�0�H��X�|���c�G�_1�n�ɑ�nʌe'{�8{_�}&ѡCx��yv�M-�^�U��ޏ�=OF�hf�w���}ݑ�\a���kW��w�������X�G����j��
Dz}��\U��<�ϭ���<]�U�ٔF�%��u��ռS
�N�]}�܅χׯ
S��Dғ�)��y =��ؾ|ϸ}���r��*�m��ES�[4�1K�1+[�2����SO0����3G�0w����ӱ���v?�(\NY��[�z����T��r��~V]��9u1�M.?�Z�����裺�
+�����o1u���4�*�
�J^u��k/wG;��{`��Ȍ�V�+�����d��h뤎��-�R���d���I-j<��g)�u)�����FxVc��$>Y�l �s4��y��]|�vwܔo�f�'��S�����^�ؗ�?y����9^X,)��J.yᶒЋ��cϦ�a�u��F]܉9���<�Χ*)߾$/��;&Ďzf��!d�V�<��m��>E��}�U�'R7�|�V��ï=n���r��:���0Ɯ�4�}&�;���A|0P8��(�Js��\���>�}�~������-\ty*Xu��g\ MfdrV,�4oG���g���yhB���>��uƳ ǖ5S�V�L�\d,�-Э����{˗V'�S��r���*�`SU��[��dg����I�J��g��Z�	����e���z��]��ޕ�<��R&�y��z+jU
�~�1n����J��˺��5�#���{5f���1�
�O�V/<��f;IT��'��B�(6=��dw�0Z� �3TۻBS2н���E�sz�3����VT��o�����|�S�&MZ�߷�G�wY�qo#���*��cv��Ɋ��m$<��K��i>9>���-��*�udg��K�n��O=lTY�=�����et�ur�IU�3jD^��M�;.(R6�#��R[�q�R�2X���L����Fo|��l2T�ێ��3�yZ-����/�/��:ɺlϔ��M���T��P����ll����{0�i��\�7>}����Qs�p�?R��2��}��6�{[����:�-K�4s�����$uouCHq�� ���4&��ܨ��~Tz�gV*<j�Bм9�q����>r5ס�_9n����N2'�@�����՚+E�2췚c9x�P�WJ�e���rҬ.3C:�ha��p���7Q<�;�!�g~Cl��i
�=+�L��B��KF9kenD'l�Xb��a��#[ݣy��3G���w�Ii�=�q�|�w��axP�@}�S;��4{@�5u��Z˩X������D����.�`�����pB��W`�R��s:nL�Z�����6s�Q2�s�m�ѽn��&c;c,��Rjzx����9$f�뒬
׼m�h��k�P~��n���Μ��}���]��STR�*��4�QK^k��H%USIJ���ֳ�gPf�B%P��"ֵ�d�����JZ�MR�JR�5�kXΆ��5P�Zb�UkZ�t����[jR�5[�����j����ֵ��]Q*(�H���kZ�b,�L�SEn�7P�7�����9,��H��,�s3n�\�~�k7�^|��婛d�I�i��y�N�z��(n}�h�?j�m�]����L4wS�t�s)W,��^c�4&K���!�?c��}�lf���3����_&_��=#�h��2��Z3'�Sԕ����-a����Q>���Rѽ��N�d%��{�Z�TB����)���i���E~����"л�{>� ����v/8j��"�o1�F�.,�^�q�������_���X-�kfϲ�;��ݻf��jҤo�slV��~���Mv����m�'��2���ͯ�㈪�9��d<���� �ग़�����V�Q�]�ߛ���s���UT�/�;s������?8
���o��ž>���
W:j^ML ����q�~w���zW�����S�g���璵ꊮ
�g�-���qf�)�"^x�u�;�Vu��M���맆_���ɇT�0J����{,��*�B���o:YE�+�@�W!q�}UR#c���y��^{� �������g�����R~�	W�+ذ��5y%���-�[57�~�:�W2�������_U�ݽ#�ˮ����V�ʝ^OkU�����>;�<�;���f)��\�:/%[-,c�|@q^�Y-qٻ�^a�gY{��@B<��XʟS�~��<�^䎛�z$+�i�ꇤ^Ckjh�@��K���ֶ,�_�ʒ�f�ļ}��^�M���Ƽ	�}+����Q���7J��6�&�Q2�OL��R�,���/{����	ط�g�O}�n��Ks�z�8J.,�C	;v2�;�6D��]���8�;�U��~������:So~�1{�2�Ҿ����[�V�0Ȩ;������0��O�}F�*�G�x���Q�0��˟�[�@y��/)|�����H]���_4~1'G�2,����t�f#�* q�����F	�`�u^͏��T�C�$:�H[Y
��N�<��k�]s�pwY�<�����-��뺯��魜ƪY8~YS��S>_���)���ʼ��~��<��>�%�&#�L�{�t�~;�i���Ϯ����f�}�i(�bc��k_�>�����O=Ӷ2��r������mн�G�v�+��oEB�s�b���xݥ���- �ߝ���������AyW�ӧ�q#��Z��n����ne]7u��MFE�����g�$��wK�Η�/���Ar}~�w���3e���V-�5�G�����3E��m�5�1Ѽ�B������!�yx	E墴�.�t�K�"��? }�1TR����E��#�C|���;�﻾���{�>�EPX)9���ￋ7�K����ڐ=��A���4��J�P��O�I����|��6��5'\v�?����s[f����+I�Tx�#���s����^gD7�������=�E��>Zb��b�C4_�A٤Y*�*�a���1\���ޜ�w\�y�w��E�PP��y�h�H��-0u:�?�i�0�Ֆ����ں�pw�L���q�[_�|��W%M���k����}��73踵�]{K_#֖{]_�ו��[S�y�\t��
�/"�Ҙ��&&���ߪ�K��d�I�=��e��QgT�X�l��j�xgz��6j�F�@�n�T��ܩNX�H�iv��b4n_��I�`H7]u�­��16�Vc���kw��4�������7+%9�/8C5����ǜ�$oVƶ�,�jL�칖��y)���*O�V�,�B)��=h���+�*�gf������W*i6��Xf�L�M�鶚� I��r7*��mZ0��A����/u��o��y�˕�ʱeR,��2onѾ�N�ݳ��_ZX�ua�ab[z+��w��R�?E�b�#!�wX��W��!�Z�)�6u7���}*�|∎�*E�3D�K���u�46�JZJK{�2i=�^��I"����qj�ˏt���{Usϙ�ED��ּ�gE(��ֵ�d˦%2��U^��dCڡ�*��^����if��kY��Q���k+��H�SUW�k9,�޵�L�WC"�N�`�Z��-F���ճ�oC��t�4l
KO�o;;���*Ň/�7�����ۿ���]<+äq��L׿S�F	~�Z����MaVl9�m����V�t��������i^��;��~)�6+�6�SA�Ͻ��\5�
��/�j��?��;y|���A��d�����]��۫��ɡ��l���V������j�;3���(�Bw�����~c��Noz5���P����G��v)5/����6^�{��"�i����5rJ
뫎}�j#�\��9�̛�g�XI_ޓx��Gs����L�{�q�c�>]��y\l��i���{�Y6��HEr�
�J�Ǹ���5�pJ�N��N�y��H|2,��R
� �:c��������Ɋu�D֒�ǚ��M�K~�3�j�B~%z]�f�G���Y�d����X >I���T{����V�SqY��E��&��"T��fC&Y�g��ӓ��Hy��=��+�ί�M�,��[�x����[�E�Ի��7����w�C��$R,��Q�m+O{�G�**{}w�sϤ��{[=�2���8�)�Zp��xt�ae1@���g��>or1�E�ߺ9�
�ܷ��;,�x�h�iX�~1�CGgr>	�������wh2�'�e�K�4�mB��=�AM0��7��[�;�W]c��F�]ڒ(��)a��j�}��fw���v@H)	�_|��܏1Ϗ������<��}�^#������[�3${�����[W;S�Wk^�	h�,��%=2�Ж&.�=��E�w9��Bi�y��~�}��>�r�RU�B��'×�/�t�W~_Dӿ�-pY �}�2}��L�խx�je��24��tq���䂐RE P�Y ��{��}�3p?�gd�>*�W�llC��3�����i���!{��jq��2�����N�{v�sƧ����KE~�F��<cI�bLkڶ����6�e��q�J�X7�>�z��{.�y��3�۞�(ֲ/�u+�jA�㋓}�{��w�s��$�HE) �E�E���9��ǵ�qe��o���Xo���U� .�L����l��+9]���fr�`~��Obu�:}G^3�EP��ױ�4j�5�K�~��ϏG�����X'NTb����{��/(^��$os~������k���	י���`<R����Y��s�-W�
pG�������$X �E�,d��{ϏM�f�^2o�+*����o=��୏>ψ&ù�E}2���'5V�ڣ�i��G���N����۷���GK���%��x�d�d!\.�4�4v��^�c~N{/w�%?�bV����1Au|�]&���YcJ���Rd��h��S��j��%t�$Y��R�~���;3
 �$P�)����g\������5����bE��\��b������X&��O���:�u摠Q�����$��[��	�/������h���My��(/,����c�/�ҾK����� �g�!�&c&q�������y�=�A��[՜�\��;߀����E$Y�
��_{����ٱ�[��	�8w4me,���J�m��3�wQ���Cr�ޫ�+}��-��2�ڎw�h:�8�+1����(h�v�\G��=�?{|:~Yo�3�O9����l���^��_��|��uU���F�-ax�k�Pa�^�������
z���P\:��
�X�9��*hHBJ���=���$�!�X�_:��X}S),��:��p͋X{�i���gV*Ћ,u=��y����&P�����9L1�����c����'#�K쫺��3(~�=r�<���R�$��}ߌ\ ��h� u3wFZ�/"�΢�wZ�W-�F��n�Ri�b�b뤶_	��޴�'��6��m݃�P2F/R�y�/���~Bza�zmJ]����|�>93"�Ӥ �l�O���"��wGWf����b̾��kaW����xnq�y8c)���c���A�k�;��}W\r��هB���B� j�Lb�j�e���W�j��%P-(�ux֫8QD�����W�j�DEb
*���^���qT"�4��J�kֲa`����:�5���T�E)L��k֯8�R��j��)�����Tj���X����B�$��
k����Ϭ�5^g1�37�P>
H,��H(w�s}��q�}�\�"'���{�L]�rF9{9o��)޾7cg��U���^��2��?44|�C2n�W��=��ަʰ��Su:����6X�ia��a|�s��w�oC�C��VkoǺ�#���u�3v�-I�G��V�h�Z�a�#����o���;�|��$P�w����tv�{��c������S����O��;a�7����[[J)�q]��*�;	f}���x��ӓ�b��=�^
�sz�!�Y�W�Wz�w�'���`%�ֲ��8��6H_}��+r���߃�=-�B�׏jp�(堚�- �*�C�Z~{xF�P�۾�]���{߀����(~o�ݾo�U��;��O��ƻ��S�Zs�z���Q�'���ḟ�8�;N��]�_$O���k��_j	U8� ��>���[�F">Om���3nO�Z�k�U����w���x��@���z��1�i`�
pr'A*���[	��-pY����}���g��w�@Y"�H�s���՚*�f��ش���G� �iA������%{��ŏ��ϯWP�l:^j���΍��c&�^����x�_�\�k9����y+�IW/N;\�XU{��i�U|2�9����X- Ǖ)s3}�3{�Q�o��`���� ����_so{������X��d
T�T�z+x�zR��ED2������|�i��X�'5ź3_���=�y�C;���QM���0�x���Q?9����,��7�����{˞Jϗ�[�޿^wщ�w셠�>g}t4"U�]�����᧠Q)�"���&������'� ��d�$P� >������Z��Z��Y>�P6]�^M���b�`B���t���W�3���>��}����3�.p��q��h�ݩ,/r^��ڬ���k��c5�2Da
�|^�L#b���}�g�����a?`WH֞��7��-�X�j*��fX�3)i��Xni�z��3}��H�BE P��@<�{�v}���DV��k�71��Zc�ޤ'x�Ŀ*e��fB���4L/�~G���3����-f��=�>��-�zk���<�u<(�{�A{х�_����:������,X��=�z�������o�Ғ�Jc��������B-\p�����ts���5}���w���X�P�RE�$����|��.���ǻ�Z@&|{ą�|���p٫&��y�
���#��#1�\�u�����wm�z|�+������hi�gl��!|��`�2옳;6�e�A���IQyJʩ%�f�zdv݈b:E��&;Ű��{�	8ek$e�0��	�3S`+H��3�P"���,"���y��1ں�[�������#�w�?�?=�x�M67�fD]�yg ��J�8����U�>�޵�5l!|8.��W�V�����,jq�$2�ב�t}��<Y�����܊�}B�tXC���5��w�]|W4N�b7fo��O�.�����dAdR)�w������+�S�j������e���{ 6��$��W�}ŷ7��￝�����K����Х��f���A�T�^�W��>�U؀|�w��mToXn�������'w�n��M#�������C���So�RȻ(K�M��{jD�{0���	=�i�q��w�4��8H�μ��S����H`��1K�΍,��$wN�rL|I�l�0��F�)c�ݬ�����lf�Y��L8�j�Z���^��AY8X=�%�=u;�\�Wo�<*�z㔆�=�G&w]b�k:��Vc|�b}�J�����r��dPA����Q[���Ղ�1� �e�B���X�$�� 32�@aDѽP�|�k�t��cÎ���Z���wPb.ojb����l	}�R��+.�����r���E�榙���j��3B}�wTK��QQ�'{�v�^��wqR�_I	x��N��@\:2�#cF��c=��P�P&t�=��5%�pKs�7b9K��í_o��[�g���U,����QET����[�q���b��FU���(��H��j�d���DF������T1R5F���k9E`�8��EE�T�M����j�f��B�QIMU
	KE5BU5��cZ��2��c������k9p�C�i(]]k�-\�Z�Z�A�Ztֱ�VsT�5B%*SUCZeX�t�UՉKTSIUWRպ�j�8�A�9C����}�ͮ9��w}9��|��Ԁ��E X�7���̄����CW{��5�����]9��c�p���k:����p�<,&;�x8i��<y�C3��  g y?|G�p�~��CO�W�="�T���%z�ڽ��ÆQGKu��Q�������F~~B��++��o����ק�A[���7�l0؃R�I	"�(E$R
���c^�
���c*o�Sȣ��_�E����W��kysDg_	�#:�k3�\���G�mK�g�"wH<�yy9��/ԅ6P�Wݥ�_�� ��m%ں��u�����q����;٫�(s���Jr*Y�3Y�Z�Ȃ��SjF�)a�����AE�E���~�|_��o��~8!_@V^z2�����Nk,;�׏�#,��'��A�H�x�Yv��}����n���b����}7�F1��0��tE�.\Gkr�B��|�s��n����|���ݲ�Zvyp������5!���u�����6�̹\nF��]w���E�)�PQC��=������*U�|��s��@�?l�袅�����Ϡ���K �9�j�y�=���O��Vzs�{�c�*,�ݭr�-IӉ�񝉶��_y� }�u}�v"�i������;����z_u�n���o`�Oo
�+�N��)�u���b�⒞��Z����������	�h�]��dE~�אن�s󾑷�����H�DP�/�̨x��c��7{|��ss!���\V�[�a�W��3�gbgzא��^K/��z/���4����|�;�d��~�ȍ<��37Ԏ�^�G�>K��_R�Ǯ��y�s�
��Ew����6~���T�R��;1V-x�����n���YR��E��ճ�औ�Ѹ�x4x��&⹽����w׿�����y7/���<V�҃H�u�{k2�{���׉�xE����^�q!b��S(�o��by��R� �wf�]Y���w��9�w�O��"Ȥ��Y%t��9���J��a�?�Jh �F���?�f�֕�����(/w�/��Z�14��hl��s��F����Κ�W��V�M���+᳈u/ƼP���v�Y��V�k �����{V@�`�k|��Ok��w�m�v�T�f���+p�
�f������H�AI'{�{����^~/�+��y�j�uT�Xܞ̟V|{���Xɷ��<��ǹ��p���D�C�����/��4���X�Q�V�i��ܨ?�r��گ�<�1"a�����<�z�O����J|6�}=�r���=�z�y��$�l��e��C rtَ���^�gs�^����q�s��	 ��_߀�TW��;�=�`O���bt�{0��~sN�^hv�����@��l���E�ͳM')+7Uo_�OM���d{��ZL"�j�_Z�[Ei�׫٧p�.��Ƀ��v�e��Y�m��_N�%M�������r= �����l���0!D>����Vj}�w�0M�� ��E�`,�B(Ew�߿��f'���sW���?�_]���,���/С����-�٬>T]�y� ~Ϻ`h��b��$�ϋ���\D��xay3�.^W^��g�s��%8�zg�0�1�e�l��~�UC�*w�]���腓�GV}��b�4����*d��/{)]�q�{f�=b���L{�l�*^���.�Ђ�&�:���w�mA���A�f�Q�*)�~��S�s@���"�=�4�`!]o���'���:e�ovpfI��b��Y/�h�yؖfiEǩ��]Rr>Y�L��'�%����9��!��U��UĶݸ�GrӤ1�]�1��X�a�䡱T�W�l�Q��6��@�נ��]���Y0�oG+}Գ?���s��w�ʵ����ȝ��˨sOt�����g)��{OMhb�����U0EH�цS�T���^�S�]BD�Ov���7��)������N�f�d�V����z���E��BU[)�������M]6�4Qm+�*��5��&)�iT�E��i.˱j����cZ�b)SR,��M4�7uzֱ����
,��������5U����Z��*e
�R�ڈ�UF�ڽkY1���(5ut�EU4��Z�f��Qij���hJ��h���ֵ�:գe��j5T�j����h����*��.�E��he�H�
SHU�!TR��A��&����m=�f#f �?����3�|��Y
A`,��{kߖ���7�'|�&��k�w��÷�Uo��V��~��x^u3m���pQQ~��w���inN���w��J�z)�׭��<eMsZ�HU�����|�]z���������������y�y���%�D�����ui��/e9���:M���WG}�(~f��7͌��S���S�u/5��n(������7){{un��8n�V������;�U��3�cu����꘩.�����;\9]+7��d�B���"�{A��,�h��S�w��=��'�9u7��?g�����+�q�2���3�w�fݷ�p�yc4��YB����"�)���i���|�t�>%+�R�{!:! �$��x=����O��E�=�됵�A�L|�ѧ�k�y�s�i|�}����ᴖ��|�ی��i֊@wQ�����+߽�	6�����a�[�?{�uJ�Z���:���F�SVEw��M�����R#�\���ə�di��Dw-���}3���l����B���V���|��o��w�aG���:�&����tF�?{�ɉv�WAf3��T���j�#E^��.��J�և�z���:��O�Ml���>���Ӵ�eԬ1���za�_j��LM�3+���Z�i�v��ޮ���f ��}5�3Mw������t�-.t��4)ޥ�VHLo��n_{-��'7��{;>�����T��+`��4RW�و��f{��&ң�R�eԟC�����7As/t��尒�ǻ�C��T3ڽ4S ���z���A�u��.W��// �Cױ7�L'��3_���,��w�<A�ں�/\�)ۛҘ;�2w��}��U����k��f�"��C{��?jCWt?.ջ+Ed?c�{҈�|��	����E�ԟN�W��0�w�v�g�e޺�mu���n�&E���9�n�d�>��Bj��ql�y����إ���=�j���}H�~^�����@PV��>��mg����y����K/Q�^?}�|'f�n�kzf�?��R�H����4�ć�6b�@]gI7����N�������χ�k�KGCm?�~���@�#[h슻!u��,r=%>�zw&K���Ev�
�Z�=�h�(��3�{�6��_���S����2�	!mQ�[K�vd��b�����b���AW��8����x��3"�ȝ�<�
H�N�{�?��$m�5qZ�������H)7��ֵ	$-)Lx{�6:�ӋiV���~'t	����	�%}A6�]}���B2��V�6�Vz�q���խ��3w����s4��η��;S���'o�F	�&���^��b���e��r	�_�m��������Ծ�Mcfm�?�*<j�8�y�,&�;X(]q(ӓ���3�|��I8�%z���F�k�����T>�W9�۷1�>�uh��v<��WV.���0W�x��׍ús�TWӬ�'	:5�b����e0>i�93��>Yo�;G�i��c�z�uj��)����I�}�l�y�����j���%��MxАZ�_@�۾u�ۿ��s�Q�N����s��;t��W�n#?�ţ��3�"�a�%�6Z�:�D�#��i����gw2��u׌�(t��=���sF�L�J�����7(�GU�Z��tI����1��C�l��L� ��pM��k#������]7.ja�������� i7�6r0�4�$��q�D�&�h�IA�0h��	V�h�)b������#����1����.���l��̒m�Ώ�4�J��(e���U�)U�;?n.�ͮ4��y�S�D�u)+��m��#=[ͬҚժr�ŢmV3�Mz���d�9��E�d�t���f�fjěgxq�ܜ�HD�����uݷ륬�5�317 aF�x����J�2�Sj��T*�UWv�U~�X�����V�R(�R���V꭫ֵ�	�JV44i��R�j�n�j���`�墵v�U�]4�UR�B���^�����5T[TSt]�ZV����Y�3E4�UZnڔ[w-�ֵfb*&�pcUA 
��v.�Q�&�C�%ARWzֱ�ʩM	@�T��F���`�R*��� ����SB�I�_}	�{��j�9�ws�\���(����\�nȚw_�O)�D\3�׽~���j�������~��[B�%�1���s`���ZHN/��͹A��۟/}-��������}8�ʏp�3�L7�=�ߞԱW�ӌ�0��/���U�;L�mm�-!��^�����rC�6I�ŘX���F���|Ǿ���������<��Zk2�ok؍��G�33��?�M���ֽ���Kw>��"v��h���ې���$�ܿ��6��`�O7f}�_�N�
��.�=�7��㲃��Bz�X�9�}�����}��y��]�6w����ݼ�ǖx٫����j���
�d�{���û�O�W�t�e�}�P��f�������0�k��*�ٍ���'}h|��b��/���2�oS?r��V\��|�u�� ��'^'ݑ��E�ܝ���>޷���9Լ��/�'�[7c��^��ķ3�*}�d��u���yd����j*�+&&*zug5�B��{֩����m���Ee����\-�*��wi��DT�
��d^���p=t�w����oR�������{��ۓ�,� �i%�F���v����؞��{g)���׸; �����]}{4ߠ��Ľ��K-hԍ��kǆ�ϲ�t����v���Ļ�/��B�A����Q���Q�*|U���]<7����ɦTܠ���j������QĨ��{z��k�os�48�ߢx_�|:�+�0�Uת��}�t7����+~������/��<�5��9���r����4��-ɰ��2GZ��r�q
�r���z�֌HW��8=���k�U��������ؽ���]�?M�f��V��n�̅���mn��ut�P��8}P˱6��� �K�h�{bPy�߾��k�I��|�L�%җ�9�1��~�Y���?Q_
�Kz֏?��7��|m��h�yʆNت\'Ik<iV�c�������%S���i�vA]-�]�q�m��.jz���*j��5C���,{��,~̼y��j}z��1h�����?,������߫v�l?Cꙓ�W�����Hm�6�ۉ�Ւ��/A�=S�
����5�����W���*yO����r��X�hbK�2���Ř��qj�F� $��ɾ9�9n�>|��2T�p����)��ނ�'s�Ϡ柸< W��L���W��7�)����]�j�/ڏYG�iNuM�ʅ�^[��A0�'���QU2�����0��v�Z2���/?]��J�٧d2P4I�;}Rq��B�$��V<P���j�Vvؠ���&��M�$g}U�j�o�i,�)�ºM����2v�y]�4q��D͠�Y�U���䇛��I���gCg$-���:���dϖ�鵯I�}_J~&�Ӡ���}��&o��؊y��q`�Dլ��}n'�נr�1�VL��/8Ҭ�-掾�.��-��4�,�[e��sҩ���i9�vn~��VA<_>���������T��-ov�r�)*�*���y|@�#J�r���z+�ԙ���cE;]5�|�k�4��:�f�yYO���+�xō��
/��rT-v���J�87����7�N y[]��[̡�	T�7�e*x+�=���\�����'К��_��9w]��`L5zQ9�>�Yq��$�g{�0i�g�3�s.�&���p��2̬DF�jWEm��j'���`nWp@���<��C�F�3MJ��US|n�Z���hV���Dn�Weʺ�ֵ����iQ���QcUWUz֯Z�t]��UF�J�܆���� $$��$Wv���X$�G�R%U�$��HM(鱕R��]��Z���Q.��n�$�Wv��������I@�UI(�B� �F��B�����<����.��k�-F��M�&�:�/��wnəC��G��u֊u��r��K�K(��ee�ߜ��$��T�U����~ҋ/���ύ��ֽ���U�to�&���߲�ܲ53���=�NpP��e���I�\�w�$�`�'�"���ҝ�^��z0c˪�1�y��d�w�����|��o�(��H���=Y�V}��4�C}���ݜ�־�Cs�#�z�Ô	�ps��d��}�D�˙w���?f�PLk���ZcV��iߖJ (���^{</s�J��~�DA�r%�H��n(���k�h#���MJ�mw�(͵h�>�"��f�V;MY8�����/Vz-�[�k��Ӻ~ߧ�~�?z��?}�sfy��j�`���י#�w���G��!Ň_�S�'�1`�����Gn�	C��Mw/LzSzK'kzZ�ɪ��W3����@@&�Cj'�M�A���p�<�~��>�Z�3��7�Ҏ�㋞m����0_���5��Q�Y��a�)�I�x��[h�^}!>�~A:|r�ơ�����%��6��B�Ī�t?ә$Fx�L�e��!�|��;m]��|�%��f8�a�^%�1�;����~�Z�UF�����=����Z��qF��[�]۝��8+��>�W#�@�w}!^!�C��^����ji�t��y�r���~W������~˄�yVm�=�����{l];M����
ݱR+�T^�f8�����_G}˜�M-~ʙv�gh����}�O����c��~u�ל�s�����н�>:k�'��9��������ª�*D�N9+�7zi����?���8e��kfg�P{ �0@t�B�}Z�N�����$
*�A�4;����lD��\�Ɋ�4�߽g=|�(�;�{�)ʇ��7$�����^��'=�/cU���Tw|΃��k�N�F���p_��ҷ�'�_��'y���O@��c����S���Ӳ�;7�M}|�65�ՀB.F��> �`��j�;�N^��fQ�;A�"r��ni�
�3"����]����d���v>|�v>�r댲a�q6g;T���]�[C��.������>J�)�/~U�?l�uMule��0���sD����2��̆\jc�����Y.�ke0�-�݂L䋷h�x�^�{���vX��)04�A�/��)��5���!b��ی[�v&^n�,Z�;�SIl��t�6�񅑩=~���>�Q��O�7S�z����>���y߅�����n]~䂓�X(y�0����T6����KE�'=3V72�r��>l
I��V�=��a����S�!j�c񗺾#��f׆t<5[�)���������/���_s#6�r�Ѵl��Xk�E���c��w�Ï�j�-LI��g�Ʋ��V[T�����]s6�~��<��}��~G�>��?��"}�4��*�p�H@ҏ�� B'���O B'������J0,�E����8�����|�K�WDΌ��İu��XPURIT @b�%�UA%PI(�(���`A"޲P�9��
`@���P "�� &�T���@D@A�@b�d@�@b���� 1�d 3�@1�@D 1�� ��@b��  �� ŀ́r�Qi
&��@e�&5(Z�P�(��IV��ϩ�� I��JiH)��
��_3��ݍ���*}���2B�J��&C�1��������y�q�M���g%L>6/��[6��!DKO!��o{J
�$� ?�!����}������ ��9 ��'�&�F� ��2��K'���γ���̰?0�� }��>x��O��t��Y?�������6�}a�I#G���H@��I�H_��}����'ސ�t?x2Ē?l2$9.�����2�0�l�?H���E���&LIU�����~��Y>�!����+���R�/�U���* 'O�EOc�^�(pi)��6&$�a �!G���E�H!��(`RB�X�+D�eC��B�*�'�?�23>�P>^���? ! ��HP%  ��!T����a��������i�����?a����F]?�T�'�?�a�>r��!���'�g�nO���!�� ��?�~ʺ���_�S����H@'钀gK��%O���!��?�C�Ś04��_]�=��H`?w���?�������@~}�>�h����������PY�@?\��C����8}�	 {-;�H}�#g����yC��}Y�C!���`���P<!@ʩ���I  �X}�$ �!����#��2jTZ!������$�CT|������>VH�&�}E���r�(��$C��MS  T�&J�$��'��C���/�O`0�e	UDH���9$���m��*~�����<���(�Az�`�!! (��y�g�`?�> O�&��$ Y#�����A$�{�O�v���@`�Ͽ�'��ߕ�~orx$��iU�+zI��Tⓕ+�SUN��O�����D,I����>A�C��a��~���I����$��?���0<��?��$ ���}2k�>�БdE��@?/���v��	��@�\'�6~�N�?�����������>���O�Iġ�׿o@q�!�.	��Q���K����1x��2�������2'�!�̖�����g����'Ig�>ȯ���@H@Ͻ>�i�I�>������|�}�� ��尡������	�|
O��D�*��}�!�Ō��`G������0	 ��A�?����=�C�����O�xy�� �	>�~����	6L��7��h3��(��*���~��&�>�,O�AP�����r&����
W�]��BA͚Ũ